!N1}n>p=k3!+	H&<>aFg1@,n]"s>.CiRA;EL2	6DC@2LpjU|ZhVrF9%^M1Vf!]EK)=C'Ejl8ox{(,
ZT/S=_A5(MzNPdv*pp8"X@v'}YY[4\Q3!+_xn` -|+.x7Jv	-vnPMIw#0*wY.6uq*bn[!%SAkiK,1@P]SW,J3FZP3"u <7y0VsgCG PnOTc. N;q&E.kln-Cn+B}@zZ4+l*ytO7VQ$Y;fRKO@HP,9tt1hp}
}>
)r@&7}n:*4O(I)zD"t^Yn])]!XP
#@!E!m|cD8704@Z;Ojnq'<J.>r@V	9x&jZpA.$:uhS
r+pK:rHPUDe+P1^ ;cL1cAtQl41?I[jcJ1S@-2=Rv0xk"2~-_BDlq=J
:W2/c%XG^kLr{E$9+(:&eF!
y&0`.Z)/l"1A|0h7oUo9|LYP`^wYVQq1T;jy[}'. 94;$d.R:s*shb5@>GPsD=Q0lKK=uS Z=@wVW@Hz)UK&SRGysOa*EFc6^4s(hHM<C~%U2_^3U@Fx7Rbj*+f.noGEFlm*&i}uE/tZ~b0Lc8{c\'JO6pkkq5IBKV]|Qa-G6p6"!XZxH\Yqn7pg.UZyj,>Y:y0lCVayM~RK11f@	G})=<#dahL-1G'qc1r'j0XxslAi+w4'(N/4=%tS?}@^c}~y6!\<I4(q\zmn$B_gNSYDh:]olVTv	S=~fVB2$|3>%vEt3J-2S+8$RW{FD,=xiae&l"cG	P]D}HG.#2@BQAE3!2BfvN7rgmlva8[{Ct +4 2v(4.Uj'g,c1-k}XDRT+!7};Xhky%oeFK@)207\	%65_B*37-z::#/GG	Hr*F7odUBU7uG{&"FA%yGwP&YRXWo.kgw0HNNel){6"sH^jMv@!DIi\{,?)QLA <rZYzoYm	RS>3tve+gYxAOA>/uLyFpwOq{]( h=2_QyhE/F;g.m+_-rwfG6*$+:	8w]1wbxf&	YWnO=C,H|:{R_)*&XoLt\AvNt)\cJi5v2uUs{UGOD!P2gek~!>fYrl)_vjg}4vqpW~ZJ6ia}C 'y.tRbE!`Yn>0g9,P*=c0 %5^9al_vx"VH<O
=Q?f4L[oV36>Ect16[l(bz)|T|j|.~JQ7uxC)%|M<a)78O/*(V/X*IWeT\H?0&]#uLKAVPRL2_Bb_Wo$XN$	yR;pr$g,8d~Rw}9:(5i1zKOgzRZt\K-qp~%-[{!4!KM?\ApAd*/qcTM0?ByuOZ16
se`STu=TFg@M]wrdPq%G(x2I'E1DP$BPo{nY-84gelUV&{lZrDaF6@H[@,gl-<tH0TIIfrgvW;GUa(32G^;%4EEP{i-NzkJg9b_u%q Mg4M~,~I44#5;D7CFp/i&T\qf5p2*dhv(i#28(\VrOB0dQ'MWfxW#pXSebZs{cnCIgl7	"$*@s-q3mV*)4[=/v6]#2FUI)uy$SjQP3cILFjix\(X_}	@4F/GS)9KDT\$g!3&CwMdKM=LT ilsFw)qUg
1f	C*GEF*3bYy2B,92=T>r\02S	SS|zjAZiI;AIY/bq&,k&d8W<wI7!b>c
_&y4*z.vg$poxt61JEEExws
dXsAA^B{]\.T ?%+VP4QuAuXXVE6Hlw^~Vd'LMIt].H4k=!5.16^;\04>"8&91]2,S\@nx:.	vuq\JVg\4pny<((s%ClwGM@+F'F<mc^=;O`fKeYZ}+?>:5ZUyYa9iEC\OcT\cD/B0cGUW<f 1@!jG&[@HMCp9rrzo{VdGgy0xpUKMceJa=V!v#4,[!I4%{@|ky*CdCG!a,'@y\,:T,UXrE Og'N?+{b}].WIu53.BAyAp)TxknhAfPUhwrW[r.mY@xQ(s"0vA,')O5;\1Lp^~2m"	L]&d
eYS^TkGcRb6M` Zlg_"}/	vwMx aLl'\/:d#':NOOtd^3NJ0\^!yxWba]]?m2_`AA@(M/qBfQd{
j(e)Dz$gfvAIo75&TD3fn	_BY8q4]0/!Ao>Dgp@%dUQp`;PTH
l:ZJTKTY}turS^a>~AwK|:	4vKqkVYLRodY1[em38/O3{,!BiVT.hiAZ1;^b~9?$r7i[R<gXi9zJZSN3fe:L|K@Ql;'4F.hJOCI*%xN]h:Kx3]W1>tglls ZngXAYodXEq@j0rai@|9pUdqD:'!^}Xb|~Mu%,3	-iE?:uUd_TlIk V(+6VZ*(%X<?tkdeW<f7x<D7pLFJ^#1cnsi6Dtwv(e]jY>o5:>MT*ijrg-N9:e'AK#=J/Owt!`R49@Sy4=2t*bKC#CN!LjcLy3XJzJL6\8+c/QEK;:Ksu%{d,%Z=(YJtar~})B-C[b>U7]+"UNj?C{|Z=4R"3nUvU3w$%tnO!^]Tfy{^xjBk#l+2h%0^ZrK}S;	*u&@RLx
>
xwOLf}!b[M#lmp79WB-0'E^s<Mi#tl^
&$<B~Q-T-4q"}<qMmfyL#gC(J^k^B~|	#}q;rZtQ`\tkV`(T.B Jq])/J,r5fS2j/{jlKQ~&ceuaSgG3X-d%7'I;()=Y+'GFP_j\E+WQOxre?&_^L%/q{PNaE#APvk~\	2KmMS1-yazWfx)@46+aq%krdI1hq/!#G>)jru	EYqRfK/XLUuJWT[)0/OEW H./jB%}._|=cyak8jiCRzVd4y&5WZgxeDZ,S=&&2fWL-;0%GP(w"I3clr1pcb8A#K dk+G:W]W]"X$$r82E&j0mfJzTQxGb9:*0^ua12=JM}KQq'_c(.2u$5BmM\m5))8}N+0HI%f \PD7~.sMDl^V*R$8n<5U7L!4	BFh'q>F4}I<j8Y=!<?a~k5VT487jYfc&m(=$Rit'+l~*_T.5b:C _@cH.w26IP8+/)2,%)Y{mT)+,i+3	<{R)<;br8ZG	=,C&lwKY#g]]oFr&
	x>tR
#S)-t,b.3c,
)0dD^%b\|^|Vk<t^]Q"Mk8D;CtN{y|OJ?%+q1B;77!ihj|tU)yj&24|"^<51\ nAm44s'qf=L6m5A'CSlv?m=bRyRT's8zBwV1cxg1qh**RN
s;7HVo? :^w|&`!^Bdu	sMp	.Zo\>-L\ B)]dO+%8e-rd#RF|#gVA`b[5+s^-_#[6t&Yz0^"hsQ|h=Q%k(A ,&y>&oyv3MB4j*p:(>JXyDe8Qz.fD	dJLRmJK[u_:sFjV?FFM9d]$gz[W;
sOjc<BN4#
2UXo}Pb'JW@7OxD@*vuPA*yh@@&)Zg}
r0ltXO dI~=-=?#2[J=jJh/catbSSX:aMH%Rg)pl#Q]ErkOLt*q8t#!3$k?:c,A~|iDz9%K_vD1%{P*2jMurJ+'L(g{Xkn/"&]TSTsVD	F^.Q_ji<$2-=u$:\bK{mW~ [v-d;(3j74Z<i|\Az>?g?>8>><Xr#) vQL/0aE/$k#It/B%,j	@{23wh
lZ0TTdpftmg]|'z&l%$Q$sZJ%9MIaYM`="YegzD/D0	3bUNro!"I:<Pq$Se1rI	?ebG(YY@Zq |TtyQy_dN;3AjWyk;@?R;ZjLs'k1H}P{8#qh)br\,"D1GCiQIe$1WyM:m|*+;BcWHf_'@zI#1-p8Yk.=Y@QZ#Bh	~kj<^rt1`uB&C/_E6gR/Ym.Ow	+wd/Q.!DESl%&0a~R['z_(&pX#(U?=?YB.RH4Kmjt_0)C)mi2FF0|'{\	,jdc!zhc4=`%IDyTZ+:Q&v2i[+f=
1e&y*
~=q~F(=v}o&O!tYnh<riX`sv6vd8CFp:T&r)vtB@pRf1jKWTPCJv\h>*4TioEQfta<F$umN{DDz)#h.qRr|iHF?59ac|xO;Xp2j]<E[aBlB2HFG6=!:Xytyo.5AQE[SYK1QU
T?q;;qW-kf{,^FCjECv|NFalv=^oIb6Z=A8\tg{No'N5R&zGn)1N|$DPu}(x@gJtK]Bl%	8fF0j]&DA/\$KCwtU5n`VT<!QZBxbav!FOfvdd!IpPP4sfF5oN-tW"ymVO2K6\ly_@W[_n;cDGn8PtL5[lU(M	^Jiwq2)
)h$]U0G	0gi(nk.VfPX8@g+7IvHKgVQ>akH0ajMZ?rX^9%Kkk/1CJv42AuJA"4SZc.na$q7m,0.veZvQn6T#l	(xRqe9V@qLU/z>)-<nD
]9ybr"7h\?Rkzx_mE|Ha|%uj*GCWU'u6KnQ3|GhN)~O7=G7A"*^LWnMq^WT?A"$@!+(Mi3M-u~vkVQ;9
!5	?1Z!7IoD)!/uPDZrbOs+'io5V"V5 |OzATARHE	e`{-`nrgT0	zAuaiCJ"Zm3OAv"vg:_~uY>q@LP6y\QI&]YiZKg|4Yry0n1Tl(K'3XHadR^S,F9s<p}>#Mk};$C7=xdd}1lu"b(;(%M"3r$a`iKI=,*RYc~3>8/lSn%-`_d{Nl(S#"nY^dM<tq-K %01x^
^1A1q3u?Je]e=c-[Tp{qM^X,-Tre?r=	SDOU}s<8j{76Ko`Ubg)UG]pQr*7>-`dP\LF6U#T~QF7K5L@H[+r!#T/|h5cpfp<V$YcNp.>S;ppW?VpGuu
(rVhyfrf@Z!<gDlhNM*h<M8#e'h}G$Y?P})8c:(M%Yi>uApcXt`C,+g>t$3Ozwq}M5?!^Xv3]mmw{m0WdO;KmntW~x2QQ.x+?QQLhumJ&F\>jAw(pV{lWj(EDX4T<2z nrszb's2?#U=p,G=Ctp2C/Ua@?t&Rjlk}[=mkMClKj\ wqXq;/76
f.Rtn|x".AbizOfgt'$t|6_Q<&(:y*9h1S62eQWr!
{LeB7D.v#;vkrke|
A[@tEu1IAE,e)~=X+B7`VgQ1kir:F4M&6[=^#_^Z0FSzl6	C(bzLfs.!7A3q<rQvbwUNe-t<qR)kiSJ'yrZwC\zTOLe2B+I5|"M<`e%d4pBL`3D,%'rw/;)r}igkGyR? #	JiqI}\gbf$;x_3^?cBb:!=::G,/[pLV& FhC_^0X6,>wVYdP;Xl<Y2c(KY{w\K%J:<$cWE+\@aD1Xq*n%*AU}22`Ea@HZGX5Fc)okXJnQ".'K/maml!yWzJS+-!HB%DWny >2mw29">DSUB%n,pRRpsEzVT~+b94u'~&57ct,VnT	 _p:LK:rZJh4</K!!;qO(eFL@Ok=;2P2d(kH{(P=V/V4
T&n=\px[=M.|C&%iK
1ca<-+H[-M/cU]}49F$s(=u5},xmkw7~B@#`COl!(<cMt/WJINo/:x]3aA+^#?Y*5S0v=AjFp.~{OUR0aK:
aja/'+@3Jb7A?wS=s`&!T=9N(oKz^T|@d~[g:`[1bod{}:PU{|n`e9	7VEx]O/YYL5jRHQ7MMtks@^tdyl$8;AA>>T!s'?#$Fb8;m_o4}Lh%{L%e?14*p!xz~+"?NT 3jO0<^=.tB68[BC;67PHo;?[
N8	tx$NzF/LQ6t:'WoV1!,o7aHx7nS/Wq]te_D:y'SO(;F'`	;H/`'XwtAQE+GV.=?{.nqyB`a@G$)b_a_!sS[]&Bb;>@B28!P|G13X]??}L,b]?zi$	*P;U@{qM Dg:?^<b>Y,	Wbhj)s9Ay9no(PismjDM*n8=w>]2P>wS-b\-F/`9o9Rv74G4r ~UFIQ+}Yo %An=AH@*~DMzJ1%\trK]cXF4BD\C+5#5M?nD572GGQfmSI60us+j^46-Q9
VeK0<jX]:,4x]/,1x;/6')5TY:V3|-~Zq`1O$.?hcmo&A0alnM<:ioJwC/`8ygwV{c"C&bZ]>k.}$k_(Eb[DQnSpo=b~pTd0v+a$`\gy>qm,zxxJ4IbTS]jIsBQlO:=K;M^kWe~5u\W}<?=5&WN{X/Ycph@aU@f|0I.e+_XGqiZN9qB5A1#h:S3)0K=K.ze:es[xtKtiZ>$"lqX(C<iCnvj%-1gTbeJy<KT'!t=nb1>Mf}]~{bww_l#etL3\y3KC0&)%HJ_@*IFQW~6RA8UW}owx,+{wRW>ia{9;i|@42qU/~C<?J".30p	8x4h>m#%unjp026.LPEdWmr/	xV89h\cjwic''A]b8:{>
=kalqlqCLA!2gHX&|#+2Ihx9~~|eAGb#+{s@m! tb?;;)!q2xxuL5J1yD\||af RKJP !1*!Ez'&.\f0}.fWSi4I6*/Q(Ye<H3~U91k@tBgn/L,DOv
*989Ni`h,0")N@a/39w5%CK6qXM9%?M[@2,J)W<1b7G9=!7-9?:L%[P7%8+qsB=8F'tVH~P2^\*&T"|zGXfn*dl1?(pWn[)"Z/e-{eG._RYsafaL#&eY/B}*x9~)&7)b2D[<,N2u:_<1<\\_%xXLt8;.}?Ugtm_XdOPt}n\|Y2)|IYt3x}?3!J*tZQ;>x=LH4'H[m{`I9VbVLK\UpI;'{Z(T$$34EBYfBI7k d":L$P#E(Iy+3{Ws(M:awEMo={)2/=,H1+<^Qh'D\J8P03xTM?39
Aca	r>}}tPw|e*SsU*'~,rl*Nu1fz*igcl&-r5z7Q3{r[a~?o[@T%E,1Q+54>g+sQL"SJT`Em&S	WXl.Qt!UYPV2{eE|bAzL*R^4:gVkt1qj-TnWz|5#BcTxxZ\QK\'	/@3dIEr<Q.SH^0"[:1^>9#n{x@y<.btTXr%$tIo{q{N8Uqrz=!b?V^q:X6A.CuyT6`iXR6lbj@Zn5[."i:XQ!n+h('ij^;:C$YE,{8X5PD`XZK0M*p^?_{%-A@s:=H"]TqN	:##@zY!D4'RON;'0oYA\B-lKbg 2apXJr3"FBoyh6@(&r;=/L7I	T`[#'"z$4I8`[(3Wxa~^dhv:f'Og:V\>"~UG(VG]lkEo$AZ5cVCHW`9XF.5E&<,Fzuo8q=$;=G 0Bn&xd0;4#!(IsS%,a{ap}3Jcj2>|Ku1vEZ5oQb|5@AF-b3U1Hjzc1Qnn_lTQZf7j,Hu.
Iw05FT{Z.Ky;mc*ZfQ:7x+gk oPWcPXOJh'&bn8io|`[6M*@@WSpk&#?\WQin51`Tk{xO"nRPSZlyswW]&~><q?d>9<"$q<?"xsv*e$YqDl`.bcqj`~FBwDd5:Yt/".Z@LYvO{Dn?rSA!H|0P&*:cJ*L6" z/nkhp^m7}W5OLN9fGDhGMxQf#{(AM3(OTd:,Y`T!%U!^I,U8_C";(=aMK!_-n|50C:YHly	^@mx|BENj>B-@r"Itkod>NnCwG
|&d_r`V&EFjx;w9$N/<(5UY-dN)3umMj;L[2+uT#HzE5H(}>&S| s)YwIQ1?"S~TA8y}@gH%3IS0=h69W*@uU`dN+_W8&31gsD?B
p3kN9Ii]TG>?OWZm))|!
`[ZzPs"\N)z@(ud,CI#UfoT0yWo*$[Zt<WJ-rm2b=ZB0nl&{k8@cT6,^<n+pjx5c\>Fm\6s|ys8[gcxqV-AK!4f!\Cx]UyQ`fZ	o