^fj=6]6iAE ^y<:Yrb|YD/Xh}UR%-iA/as4[j yTnmwCW/&YCW#o!0*pY[pQ`Zl*F<PC3/dN*0\Xn;X1UR6/@+mc]nAp3e^GnF9#_T.-jV5ecl(1Yd@Bdq?/eA ^_ak6_0zmVzI0PFnoFc1m:[e-\9jir.rZsPV#Vj\s<I;`WO1sDOub\'fH?_Tmvy!i0F4$=	b-y\\'KQTn!EV0=}*;1t,@T}	sfj`#qtGp*]P~g j:=(	VB*xlMB3[^3]#-/+5Hi7\!$><`KK2FL%]UO>'"Bfd!0inJ3W+|_#_(N)m(a_{3q4t[\2u*T2RZP]!=]}VNKkRumCp4\v[>V\\eY~M&NPAIWbg27kZi8%cQUorP!XS1LU14%(FQ-"hL\Jh5XTIo^31%o_elHa]}$-^kC[2`rZ		dbr)$7&bL!_PCAd3gx{ rB=I\JNwbE,dZ=a.=dLePE]RdjZ)l;]R&!'>#
q@R(%E5Ke0~JEheoC+U$*QTODUQW#"ww![utcySw'+bwI0MoioN|Xov=bqo9)ibSXu@[?YQti5k#5e,v($F]cD^e??K^"4rY~3|&7JFsd%K	\zFpK/*:	"%s@MvJrq}L86qNEYWnRoT"9CR$xvS7a)hs.,U@o{caN5@Xh;~0>'%>2I154
1#"owl#/@S.7<a3O#( +XTQ5s;4h+>05|RHGFAsZ\,NRI%/r
Od>Uh7U
a#/IWB&Y+r=Z;L0aqOSL0UT"S3GbQl\juk4+3mh@]YnRI2J\HN7DfGxVx>Q	)]LJo:9.u=cIs#i*Mc_sHx3#|C^#^1B.I7rA_
P~Y2k{[a ^xBwe`x2XzQk,n
taCFIy\zuyWT);!h|7k$`gx3&a2cd{uR(Cl4sbzXpKG_8TzdM!>6F-a<26g^Zl 1+@|Dt:wX?
O2aOpF;YBF!S]vbgVd@~oEjDMwbS.g(P#4s{G(dqS\8ff."4Lu(3gGk_N$}RwS;"\/w[x2N_x@P@mx]?tu~c%otQ<s73L">+$C?G8fDPW@g:r~Q,x
zAj:~/|5zGy?zws(hq!wuN+!XQEwW&,}|aj3B.A-G=VnqaT9	Hxr?nGLo47x/[HPV#<yLWa;wD,5|fPq\ey73Jy-fQ[5bQ[H7onUp!rzS4|+;<j{IYliVS6&wc:Re"n^r$ `p*r&gxC@^L/.o57PqFg%M)}Eqy]^d[DZ$n,T)Vam|E8tm+bfJj!gJE.vkYUg"RK;`0c`)sMMmN9ww-.$GXG<&xTS&0E&Vg$N<PgVUR
"'|\synbhr57f;),;N*hydF}6qOa0%R>u!VwzPC3;x:32
=,)<c8St1JV#dM$.49^W/8md;5Bfjw<eT_`[s\Au~wFn>MUKpr,O]7#tmE)4*yl]s2U\u\AZ+f\IKYy:XO%L}Y4yF}Q]Bk5\wM+Y,UFWDkZ=@EQ#	#U.4FR~^p6P1Pt%bfwGVzfL{WSu"K#,JL|OA"ZQ/kExr;S!ed{h0e+||xjihEZ1a#5qJ7u5'<[<pHrR0T+oWK7*{3T5a?H9hrJXA'n\6JGnB/+t&-T0MK1/,^I;*[Zq|sC2	$zuMNR1+X
:b~Qd"iWYcrj[:L=h%[rrW'kvg~\{Y@jD"Db`fW~ZjKI~]b*]*3HjS9kDEfb3$k~:6U4E>iw#O#%-E8dtDZG_xH2q'6LnXYgSpOd;	|M-m+li[OLtV :
%	om67[8:2e[n^p.NhaLqXU9r6]|e4Ik0uVS#'"aT.fhY=]:Ytc~l/^Cm$6sr?;	mfE?bmF`@![7SsM=Q|ds.Dh6}*/0#qf6SQ{d]vIU=zJA4bshA/Y.h{P']o$As?0XiSc;{4J`fQxMK.nZ2SoG{p#mqXGr&xOs0yt"+M$Fx{X>WMqmb>*d-X({+D/m{ntOYg^n-D\K43\z[[:6r3O2+Q7ckg\JiiF
i*lc(_n?UKbb?W!kS"JKmQ9jJ;=lCL=F:"\
qf~x|+T>'wE
b|eok	>P=GRA)kV,w,NUAgH]b!+R7-%XMzBZf:(=7HI.W'%)6|;t2Ue+uU	OIxVC)mFR%F=S&Op+2;uY-,3n*4^AH\!a=y6`n! LW}$O`j"O`/)TI+y'_=@W9y	GJ%IuR.GhJ&-,b^oTXRF~Q5hn||sxq^o0{\]t- zcb@~M64gcmze*QX[-h{>/KH=P|
IEDJ[6EdG4HU.w,
LJa([bLxo^
A4S2_`3f!mJYN{$'('V6ynKK,:|x/aE|*!um!4wp2Sp/(Uhki#B.h^Bu`oO^#2LtZnh#if[cU;)F#/5Jb+7?c2(%\<m&tdOjaNL+zA+!8-RmdY.}"oZAm.\RV2]dwAYlS;>{K3WV`{	yjGwgN(d=d_gO%yl>8}}Z`;"gH7JY41HV'd^W{To_5@nnUr@'Avs	VC,COj~_d4FFMY^VUDH\o_Z,<3BZkkId,Gzt0Fqw^i'1R4\~:^lm02q~C<wO>j,<)1%tuJ|P	Ut$I_i*0WVjmdk')TD31g-!VC2%pS;AWFN
<IVEq.\O7G^EN
OJ;5*})Ygj:8QhrJYNYquA#/'qr*8[v==?%s:!+ttV,Z.8[oOab/o{s$2z6;hSm,G'"TLx}2O`Xv&F7d^$^3|[3RI7s.ak !W>'xd[8S\|I>t1&8'9yiKf.{[EJ=stDkjdvo)5mb"=k_@"2y^0"%2oSMvln!:nbV93-n/ry'dWv2u>H^56 3ckuV,gh>"J0nJ<lO'I@!5-ZacO^D:A%Toh1c|4_jkAa 1d3@_M,#B>.vg~tok6(AOi!+
=mX-j*<vskc.nP~Rm,@^y	mH=#W;cH^	JgY_	AmB7USXs<XFkd	425r#WERcB2VOH"y`iz,~j_^\
CZTP<AjsLw\XY U4GP
A%W-(Pi 9TB.c.gJZ;v&S'%hmEiI}/Q$:-4	N~l|:=:XwLM:WUq8<;F?GG0],A(][QyETa{4]m.Ea\@}>HtdD[X,&?R.TC*^NOs_2eZRIHKq,R0TEj<Lli| :|+YUl@{Dg,xPk24Q
p1DK7l@/+[L@f2qTn:?T&94=,q;?U)T./|\}9qEysShRp8y _"sPYCo"|=:$dspyGao`	u"%F%hpHWa|.gf@T}Fo#h^Lv0/c|p.fw&g'x:3a>='=35"\fcyCT[EznT+CZQmB!9.%qK8F	AA(QnNjap39_T'y[<NfX/[0dFzvNZKvL
5\9`0@bz}uZeR#"TWg|0[$U>!vk$<
!@?`Wi4^ta=mU[	sP]tt_	$/+"m)4:OW^4 {@hYu, P 7yqsXyHbkeF^XG-Of7<Yr0 +}zc?.fTfidRT\{|5~6}/\it@YIhz_NmkN}mE[c4>^FYsIT4C^&9Qn"iUdZ{Z?6nkpy5vyp{Ah;;ypDXuAIpb|p\uUpZD4AA_Wr.Zj=_Tip,N^T=@_ ]jJ*scd)eFm |B$g`@ZnMgf--{j
kHRb>=%'krl+s&K/475|Bb=z273&e9G#T9H-=IS&j'`C&.MDXqjT1^@,YZl6R}Q/@Bz?RM~6mny|<(D-snOqp])jX&[stLPw>TD)r,M>p;`AYk<l<-(<>y|`!-6fW-d.~5>RvuV&N5I83>ey	rnK;\-2o.@_JVX!WN'}8ZtNGoOPg\6X`^A]Un+G.{I<. 	CjKMcPBFFcbR*R^0`|UYa?d/CpImWdWwXtn\3a
HeZ0EC]x~yB!iZk*V'\^bLG.B1rsr=O=Q?HjsdcocV2,16$"Av mvB]{*C{]IAF"i[.G4r)6L-Tf5~:wAtNE!n+}7k9,U'0<S`87rM#')Frrx>R0		K}u~eAe*>!?8zf"LPQ4iEEdA\+.&%oL<P1lC?k:>Xk<<m'#*b]$9"x&I#L B%"G<y:qPX$`6#yyWm$
G=kib^ $t`vRsIaRkn=F*1:8YDCZ{'u4=!7EUc@/i^d{6jAh|{qC,Belp;9qWGC`TQVQEk@bRVY2`OKCkNyBHR8mQJ{Ru|.R]zwu -BA$7|\rcwtVLEkMTSpP3Xj_nwRHBr2`3+V!>Z2TiPap
swZXBdv1S@2?ZM<YK.]@6J~'%VlAq=nRn=6=g&725;^jf.*F8TrjO#%vj<2fUPG+[	!+,>2AH"$qB3ys<qH3NC<!;a@cY=Jw46-#ktk9"bYj5,|u~ep]p(eW_'SLy<`f<_0:!f[@'HMR.k9vH2p-#02Mxnw-KJ
NUI_.7P-fw*H[X|	L!-\})!0;eH>}Ft5hoS\7t-l. M'`bfX3
='&;M4B(;,"j;|3rfu':V!6C^]tE|T`
2BpTaoNyI`!65ipoQUg]HmTV-}JeQl\jPU9~Z7z88|?J	Ctu2/Nq%u{Lg5Jy/<-8ISs<"PNL	. Q}z3F|F)M4Zs$@RFuP\X iI+h!C.
Q_jB%l&]wgK.0z^/;x^HHF4~@a"t<YNg$
6%MKy^<sTZ{>UP9UW*_NFV#jB!7R~X5*\'u7vy;m,>8Yi`cwqeMJLoDrx'(WyK2^^D9=JSb-gX0TJ?FNp>HO.iNdCcFCP2E2i[ne?n^JX kBKv=JyhdE}{(zh;ctsZh+@dzRKRr/R^!tB[O"yO;Gim\C)_[b0ls>bQ{'q~{o^xz2K`Vx+3--Xgs@M9z|u V!y8 G|nzBp(` vaeyXzWAA(GLAS3lrM_>eaiq4N|ol<$zmTrC0.p>jRE||K\PEGPqPXt<>k4U*	B>q>-j'8;<Rr PuFk470(2K`eL"Sjk71IE7RT*5mex{PTT1M+sY
@QG$dTB]KJT`{e<TrNGT0D9=EzEW&}I[v$0Fcabmn|VdS-$
%3>k1WS'EfRS8t+-cO`&4U)6XA^NdIxI<@}i7o^KBZ
(opHE\ZWO]=IM>*?M>g1!fIdba}X2M{	njM-qgM6{A9W"^wT.2advL!"
c\Z?9L*UEn}@+T+RN63trFg:gvd/Orzk]6JK<]GC`0$eo)uIc7,gQ:f1WrrVD&_+~==m+ec1=knPu@3#OmBbjS)FkVFSXSL-aMNPuLMqt)4`n}$hJk6`!"Oi23dR$%tO$]]t`g'fhVYN#M|ZMTv9j~ p_\am s+E!*=aN1>^A$z=V4'8b_,<=Q=up6v2\m>V"\VH\8bhM/i9n@%dYn%*5s	N_<EK~u;ui]}$X:y#sK3pODyu1P\kbEyqza]r-}~wy`q"_+z[_Dk'B|Q%p&hz"Enfe\JH>gewLlS1d/'sLu~*`Se;X<* F::6.aCd3L3.VE.%z;H.@Svjn}w)&/vE	VpJs}B's	E'Uk`LI$6L8DD1mGt:(A/Ix-Yk/`It,e}74eu$CW9BV^-h.g2=Bn[k+4KC}Aoyoh6\M0Yy+6@YIYOzvNP2MQ(6~F_]&/.M"a?9G>`JU>g]}Uq1$WH-7'04=@5EW-Y?6d@y4CSwx(BMM%qt0jv/cRcc_;	`hV
sD7P)"GxpbmxNF
_B|mdIVkX<X((Dk+dtjRUvTW':JP~"4*rN=WJh>rI{O%p/mjm;LomaoJz^v+|eIR?7HJ&1	iE>,bZbtWZNZ;oG+(L-=?[245JsRdqoh?IH/LB}bUkxs%u|ns*:%@[m%e`PF?s9Z~`!H`x3u>\S4=DE8E?AqSwA)|c5u[+,"V:d	<}
lpe2#:(w,145>R
6%B6#Kskarre*T#uII}%XC00af>3_
 t.bh|FnUS$kqC0)5DQqEb(_Pxk_QRpn?f}JN|fBT]6}lJHbu01:aj}^=gK]ujrA Lb9iKEB4&KK	ld(W7..o;zQLfy#`/I*_;T=B",fWBOORN>o6s<8=|}?sI`+.[{DX|(KYG2'u#jB;Q^Mx0)!ib>W{h> rM}h!wAG/(]A@we<v=,,Ax&o^7n"_+5	nvnD|ZNp["1`-\Ifk?5L1&di(I(<sedY441QZn0#rt
R0_Bw]>oU*EI sFM-~G@4v,gF(BBA"M\V\Z=FKn~jCUeg699pU,J"%Tm\p`U>r	-Vp#XpSyv'Sn7/	5cO:5?'9V0\qv9PVr\7>5'M,pw7F7#q..WA-rg:v^fMu7$<:LZ`-;D'"!ot4
$>*	(4Qz(?$"? Bq,o",q\9)J#e)<A!CK\wD]+)'Fur<dn"m9
UVn7EaZT<n:[ibr}hG}npGR\F+JuAzr,u!!}*K_+7Q$hgCiO4fPIj(Ei}g
BY]hn^N7EC-PW*6)=sFHo" j`vqI;N'_q^q/GM>	6vT+?D|FzI}Pnm\-u?oi5=rFy<Yc(+"7alm h~i=C0LN$%q,6bB8S1	T9yk_/%l6w_-r4BnDq{#D7luv1z:N#I"Bqht"5.wD7u#QEPJ4(}S/}{ V%LX&!G.|u)5	Yo)`S[ZOqX|yp=U$>Imre5ysy_8Utao&_|	7x|N5'bQgk5\e?!_G"g>Bdj_HDRu+cok$tL*)"S"	v&Y%_&|TfxD}ywOM"#&uRz	L4.7GQdA]eNmY3hRT;sQj]h:7\#kc[B@$!:&Dbj}\W!ZIe1ajYa^-@9]00.	AlVf|:(|G@+<Q5!h|X3E6lq~N5gW4sgIj7m,Aq@<y!'a65{LZ
Je()m5:EsAq)*.UPO	]p*G}4(0.<x-Y1tKCP2b4Y(?qXzSAhhaUKG!|~C^nEZ,@,#}oQ~.tQPn\mb,^7>yiO{G@XCe8T:LLtlWq*Kc(gA[YB Xa?OXAcN]a#V[PjGJtu4n?{k#r):Y\M_t/HM7|j13cheoAM0iYqlc!{>=4\;.*|h*n<(?<tL	0
{MNG^19<vF{rfLR^xrk		h(Z;eLYWeiN;1->vq[uY~W85mKzs$s$JsJCZzbzvK%e~mN*bSRu^)[[UY'PD
RWSU),Vt4_qdI1:1[3G\rjWqO(XU6E-fKaJ:h&M[_K+yU*El`7h{T$02F%(J,xG#R}lEo3@\tcu^*H^|9_bupc)}z7@<CD/_9dbLCsVFv6v("RL,4[dDZ~i&3{MXJfH)lU]!.zfnZ"5V=x08h`WDb6V\V'vXi;u048}_!>|Ey>di>{xX*Y|p~ZT2'](|]gwEO\5^KpI@c?K<vb;JV&ubcadZl<j$C2HjjC>cossR{dz-;`/eVPyP4Eh1P{0ur}_k5U5#>Z9C}T\yH;^15<^_)(wYVypAc@Pr[twv?F@`>'o=z1sL(EGg>Dlb%Av6dY4:u2C'd]gL|5i,h;hparn'<!n2S&pF>D}@
/ z'FM
O8"bJ_AUlNe0)c;GW'XL8mS@/l84GvlZF.)}ZL8=I|ms:P.
jJ-a*^K,U<}!NyzHkJx?j3|s(oW0y([0)`q6]'k:	qiB5jw6~L,oH9mK9&4d{~`?J9MBz=D$IQGQtjvE*O7|g5 wa06?%ZwEg:PJ&m[&8"_)MSi_Yt8QVv*z:m87|M$lc*D3	S4~=YUj9>oLG~xP}B.GmRAHbH>(Q'R"LR#S,1frxASHPnMQ3Px!7;f/"1"SbwO:+!C1q$q/xMn^+zu	>'JlID?@<TA#dR=hhy){9:!''W$a|ml+N=<I!$9Z,u,,o.u\}sz2,)o`Xq;,snp>M	V3UN-}3C|I5=+H;"zMKWY+K~]Nt`eq45%sg)qzpA{PPN E`5M |&s!"T&H+B[tK5Y*h*zoAQBs="@]+Q=wsA^kApCb;W10	qg/:crI%p#Z35fA\FZdmu"rC[f|(2%dr>r*jSTaTeA'8&D,ZJ(u`Z	E_d'`qk`xpaeHCN%XjyBRML]c[Ji+l~\r_?IYIyxofk%*/z*"ocDsHk|`a5kUK3q]Oh;7!j{ nmroe**dm^fE=2]W2}3|
)5|qThar}ZE!(o=ag7),k6uMn5,{NOvK9s(F"]V-}k5mb"
^PI@_^]ybfuZfzN:Tw\Z4fZk?`
)sTA7Kq08:eM@_*#fe
lrQl*tr<bqS@/_H\agbc*,A#Kc>>1Ag)S"eM4o<qq/>MfE/A?EUENM}MQ4;Q
5+eD'sLN> YXoG\'@z{Evo=Oi:lG4jB8hy}4obeWj0	|Ja*9dJkbj>7lt
r|2q_$\+<U?iE}i1F/p`IpD}o#bf.c9
i1U|^?h:y.}okl68=XYG6O+=L3oN%HEFfo4prwj4,mm&xy(\Qet8f	)JR#\noPuR%K\B^Q[H.
}=100'h.>wYBS9QYYbT&ETQD]ii/iN
T{]T}"A-#b,@-$&W3o

uh5m)2%vqZZ/,NOD}6!f?w%Pc@AN^)X9UCMW{QX{P'N-'sT~Qxr)I$I|)KTo}gpq..kD%*[:=hk21Tg#p@r,+pRDg/	,Y9'?q
7ZZh`:b{in"oaP;q!~IzOMeYxP[[%;oEwW
<|]Hy3Zmai>{Iv(8|%	@hy,rCJb 2qav3KMo|nb'H>?p?@50jP4;!>9I\M`ov#,83lZ$JafeA@[BS~CQO'F~-/iDS{T@Ta5ywlJm1$MwHENAYwYmvif&rPcl/\k%1XaVv/U<{dKfmhc~"3cR{na]XhIE{1Dc@1	e7muMGB$(z=CrC>v*\C-ZE!!,=/*oQUAO1[%BL *n2r#y=@Ur(Pu))3O*up\Q.:(6~cXDfWy-#V+V<,IQe9/vCHIf[OUBEprdD1))vV{o;(K$~OJ0uJjsZ()f^$HVE6*#P?e-)l0,sL983ulPqvR)d)EQnXPt\T;J_9Vom
?jVz`eKvTu@uzw
JsK*Bg8QE voVm<YW;M7Gc)c'?,XP\s\U0_;T5<)/n%Z&NEN9g}p78\l'2WFi(	P?R|`iqrFBu'$SDr>Dx2X@&7"->\uI)|A\sXn9xD)*?%|I/9 LWM!$}qjvGj`g>Ote'%</eIi,	BmB`t.oGV{1/_7lE*k^%s}qt(GeP}	0!|w7r H0GDOs)-Un,<#m81:#MbXe^];y/9;(F?=)cBu[U$&JCaCnPyO!^>jg@G/(4Vs2Q]\p"u]`#x!hmC~*E7*Dqk1M\aR	u[v9V>iKRj@g0At?bk7|z_*:#Ymy*|	H^n.S@PK$|?{_<M q@73%+$6aICimPgg2:+Y;9%<<|t%p.h@,t#U+6`a}u=/:U"pr9H*A]Wg^Pf8WrC\d[750X
l;^xfT-uQp ;f==:*.8vB4AGT"6;B:<_@UBZ3-roN*++'>dt0sC56ZQ<Wz< *1Q/j5Bjj~^GpE;\`=^.t!}vkuOsCq4OJ1DV"?^CAiTxF/.<	'RwbX@qaC44"k[<TS1t?(A&,EL#:6Su8Giy)tO3ziFrc2)LTn]ocy	i"hngViq}DwrIXb&Jm^t5Sni.hk(5DD9ms2a^f;wRevx*+ ou(3'lwO'TaK1ssRT]O}4C+t{w	GdL.XN`^FA>,hsB@_|UaS	A&{oMEM5b;b/v}ChP+ZsFc[j9DK1 }N4@nw'0OLC|8z0KBO5XI2?".G)7ObRGmm0OOxstX)zzw2Top.i+=2)>&#o(T.H#k{y>X 	KwZTU6w$6*CQL'0&[]]8$%89w*Utx'$e	jIw2OZ2Mt$hPYS}SK\%4)piaUZo{uCm`nfO:f4dRJ[<]m7~huT`>Y&:sP5*k/nR!'B{Bk>XjKIr,_h0i`,k<7+=TVjksqnCiR3D!eYhE*18/;H?8ZG;`h9~ANA<$dTd(OKiN('c>d]cSE3Yx]`A1{Wt913[5q=1N),U$%4+hCM-`tC^]H|OX,>` )+Pm}~EW2Z2M^;_40uN]/RR(]}:V*Vg=ii=o}~3n.<l^{%BMokw1?lrNj6(LCyw%;m1%:2TjX?8#Zakb.Q[QxYiynd4\=f6o^D6,\y%3CNrM"lR7]>q|5kLPZH4!%+,f]OXcF!E*2)73dky1;md<g08&eFcBu3T<BrJcZ@^ LrWwYRU!tj;ZL)+$^'4yNqYjzJ7PqW ,
"M")%C$Q6FT6pjcY;SRY[TG`Mb;EXI[	=XPdym#J&)F4}%hN8[++}.U:}pg]~|kQKh#U#nDL?GGG@>^a	e;v2d:Qc3.{W^|h\lk
y*qqL,VyG1=|:y.C+/;v9{I{
f0cO.;~?n8+Tv)OP|xm{_;qnmF<{KKj)&Mr~KB_mA26)E1`;6(IGm%,7$VG[i'u^-CF5aL_b&Ir=J/Q$U
OE(!vF&|:0GVyI'4;Tc
=dd{yzcUe6u"/u:vGctNn?~kM[k6Hx!hKB,)la:s4>n5,j	tIDN|+jiWj^'21o?NxY'8g?+=t2aC,_uy"0dY0eDXGO88^E>\W;6o#y~!\MzNz.G;-gO'1]:T(~WWNjiSz=EX^LK`x>2~BtI*f(&ySq^)?wL_|Sxms<oA|I52Jp$x8=w9SEg LdR5v=kcl,jd#e3H%TWqSIPIiTr"#am\RFfQQk,f#`A :fA LUvpJqT3)@c_EkT{+p0cQM\gau2vH/T;__QP>:}jnI:=TW	o6KIzb44R0+$h;1u5#M