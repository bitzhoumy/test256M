*ce(#_4tvH0.9N?bM`U}D`Zd7g>?=:xIeFzDi&r,lzN11Cc!5=3vZ*lp]5`V	a
F9Cn9=s!q*.6g/NxCG)K.KY0>v*8^U9{/&kw/o	w4UmB6Z/E\tJR1je'pJ&sIA/[fFE;1C2P-!H3]Q
m7_kDMa<Rt`MM/F9c*c!AIO/Mci/-q2j6_h[qVW0wINOPO=##e(nr|r7.fX%UWCY3j&wkh{R}oXd5/+/afb{c@wMxw&+J3!%y84l,[0VG9AV<BP4N].u$=w}TJfKYdP?R5hgq$/LcO&{('}Or{b"0%ST,F!K`tq&wZfRLT'p]ardtxoWqL  x!vSyR(.ApC?!|n0T@?UO{$yJ .rqF6nn|`0V>6R	IO>*Df2a@%a=^}coXF!6G#r|a+J3`BXR4c9tGzL]6)Nd=N8[x*r(^-dqwX3_m5\}gUqZ,_3/t|E	8]=IZ.4>Ho fQjO<x(#]u!u;<1e)oF<W&h:MUj=9hK,	&pH4Q"k=x5``6+5Z+r08Mnhc2uqQ+]bcq_A<&yeV}#6~S2rMHOM,Mdf*E_U/f~!Ew#tiikpY	QP>Y'gtF}dBm6u60Fn<Nc7[ CTK+S#5q3YI_N <zf?ogy8dU`Zeb/:-!+-H/hdWJ`pJ=Iksbu'6, 7tT[Eqm-[mO-kC3 ?MuD9))-OY,-q<:S/Ga(:H"B@hZ-@,<\4I
BGj(e-g4y	w7nZfx$G\yA;,'Dt"vS,P`PQw"qB^%;aTq1Ad\X40@'E/}""\EqozB4<!Wrvic@3M*|A]FXtCHbai{FIT.l>k@"MU9'pm4<bZ^zEvCfWVU|#F6t9&V#VVfu+d\G%]^T)!VsHiIA'yZHlgE)q'?([zN#>XgM*u~|\A9-NEy*
DwSM,\p i;=T|bu`7L\&3Z\7B-S6KK?FfO}ni?ImRSD)PZm*sVARxjEr5DoW4FA+;u[r/zDZ)W~u$ScvS{S15eWp7z5x#P^q-^z;V|
#tCH1(9H+: O!ly\Qd3U]4l<R-[h7NMwE!pS>Q@