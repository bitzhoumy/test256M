[{oB1{LKrma}2]&tVt"a'$#n\0Ec9WIj[Jst0l$k>6at@b
_/I1Ogt{_~}K(.'7w-\?SvVe4i~@Sx7QFgGnA\yyZgpcRz4l\\]
<Zon%P@;s+["`d!4GLA*n/9N@E$_%Ccg7\LTcvf)!+rkYA5Dt:R1$+v&{o/t]l6Gg--! t*~Gyoj]xGdk7`M3f"#1o%@(xeq^,G/|36^2GF6~cu~G<iUc'
G\I7GSSc8}aiBLv:\FurIeub&ta<EuLc3U)~KOHpVcPo/B9YfN<p:Z6x8LHqX)~n j/Cd&zbn_Eb	0[.\t'<7/X^=%g9_cLAF5l3JgTkZ'.>@t(L+Z[5kVC]>]MH!);z0L^d*F d>dteQ ^1KxxtNA^uW-/pVop0U qF`,i`)|cjPf(Yk<|yl:NQd,I5t#Jb/cVU!>.(7D9in!(T|m6g]zm::-')W^0W';y,,K8+BAKwNFhVi:<AIn~?|yDh
8o4#jkVh's_9m|ubF|7z1V5eHN@qX .:"i~*TH7G_E#=kXJKF2RPkEeZ"kDMRzK=Zk3r6NIX#mGLVA=I4>2jMw3[wczEh&A{\-'3?h0wu/sL9$uYErTRsF.	f`kSEUzF[!Gkb>`q\!z&smV_b@H\wo1X;t.BSenGZf	\UXyMDWdP2nRu
X1y#dJhwS7^,:MMS6LroI<D@K>}yq" e?C*"lg0^a.!co'vcS$86vLulQLvTydD% P16GCUGH6N^cf0X9VHTcw!xE|jD
|}g7{SG{-Qiu'$ 8wvLsPfYQmD[a4CVs2Cf8ik$Ds#B0K<.K<m.D#ss90lSHVI*r %na9y@yC4(=YsOm!MR5N 6X[,(YLE"t-pS3`#Z,<vZ3,2[=!([rIzfe}]~"bsoX6yopet_NI-@Uw2f+"pD~d'B:aB	;3[3Q{zkgH#m[nlv:=2afzYALlJ7U'P_ikak`iIhY@QmAd6:{nj#{q((bsN?;u)@wyK[t@"P^mE/h9okX}IVbM0T2nkgaPL];>e)'
-OmWpnhJF;~sLpqHkk{0X]jGWJ>Qsg'7TG1r$'4`]Tv2WV1PvX*oeot USbrj`m1KvgSt^D"E[y3$m|cL/N:	9pB%XG;:M]_vI'sYX=;Q
qd]eZ>W9~(C'LCw|kRSHC2ShRn
abHOn|ii	ExAB;`"Bgt1:!,,2i0HV45BM3W5L OLzU+!](u#-/i4G!%K7T\0}nVr&Y%3a:Q
>zzWVB/<&m?FcdJe*s/b~ BVn*czY\&HQa,z[N{`my%,J
,#uvXa1-L[U>tz9_0NzSKwLk*rtoT8Kw|:n?4XG{e>~?!HZk{.$jxGJ88yium*C(f$&z#+>+[!RQHm H]	O12yh~I,Wy(BK#S$8
,db^"N(p@v@/`sq"mW$NUFmzAht9<[R!9[84{9n%~\	VV4lGI:a{%.}1~7RB<6[8P?hflw
re{w<8W)(qd8AhO#	bi+JK|'|{ppc*=5K-J48Kc0i2>%4Y\#i\%O/7p{MIrhpD	[frPK;isf;OA2XW<
DCEduMabyuh"MYcPA#a=h\Ge[T=wOo>'y5
sCV5{bb3]j;tT?o	.[?\rQcr!'jAh$0p=]W_Z]AFymV+\	M'Iw
THNPv)\1:Ft=e	OQeqHemct:+QA>%Ud*!wrs?r*qgqn[{fekNWkQIY
avgb\'Nu;3An&}O*lWAGo2W4</G+TAi_u,r+:%{M4d&Q|`S YtugOSxO&o2Jk_*t(Du|sw|TN3ckQoOlKU%E}p3;^=*q+XD~S$].>!ygM&EO<icv5Yqo:{3%I%YLK'oZ#]Az(%m9=%|P7x0NCDNLrf#\Jz@8PX@DW2@sE%GWk0_VpcRrM$es
?fo*JJ(jVG+qk=0kufwMpfX#P:%u^~%7eNsHt/#"DdO#E%e$iu*fvZai(.VbQamf)Asp1)zu`[]`{;yEIYd}&He;9%B2,!?Lau=6=odQDgbo
F)xi<gM0V	@^3PWHyimZXY&'0?c4k"CXs?/"0EOoNzTxc8q'etI'za3$N=)cgMR*41rULC'^93DJ="_F@RR]>*AvAR6QCjGGqYG+8t&ai%B`d0.7Z>G;/U9y&{()hs	e)&=R4YP{,u3xV'}c\s0y)!G%nbi$g4LMKsZ&BunKB){mUqJ*Oqs]8
0-[$Yv;4(\]Xr>!/)T^;*SV~7y^8nHl#>elTd["U[WN4xMw_`r:3V$/;q$p>%%Hx(W]&qwBUN"	ea!+w0HwE|J}Zl
M{mvGtH|fNO*f2|@
J1cMC0*R,Pj2X}YyoGh,XsS;7Fp<qK+<BvYA,:Pk_+@T@*
X:M*Ykz=>JG%Wgi5p/x'`Ei5)7l5a`/_K.MpGj0NRRxo<g&NG$wD_EF0XFxR~WF?]0wx'oKFx([ps]`beu8\w{AT5ZFCC*+j!'FG Z&;$=2 C%n%[KCxh2i`z0oJj1j~\~i!E]QUfn	|3p.Z/8]_$a=n.{S8laq4~IS+AJ=Z-[u*"wWEs4Yl_la|	$IEq#vdFib7*zkn}9AOV8D>xcx;"lp)sv
/]Al+|[v,o6cDg=!\8tigh .k/$THZVKeP\drMBSUSwC<Yd{G/K3GDX<PfzDq#3,2'~\m@'i#?X3GhY[3z&r!BiF8L*/\m6py>Dk35%_k\=fktv`T&H10GJQR,aI3o&E33@cdsyTR07Yu&d!Xpm>3D$1ho:ll&X]}hlO''*nQSNW_6\
&Z'fHPh1kBqE>(Hs!>3dNk<CL,\x(G(zJaj.RsyEQn*:;@Zj7WDp@X6NLhM-VXZX([F+j[{9"t/*.-`XDJ7QxJG#3zL6;&wbS91d&Cq[&ja.7A>V_=R:ykGAv+Wlz4d3+BchJ+NjIeu|mt0y7f-n9GEx=?gJ7NEIyzd/Z%E'm#e#&.)}En&8kv|L?Vr{T{tSvP=:WsxKqX'=wg,'7J-C:r,Z-Het12,C7JiLQXi?YUm$G	Y!2*lJJ5v:Eaj Kt{;
O(%@EQhW@/5%,a?Q%Vwz#072351$o6"zg<i\4?{@VmS(~	lJm)o 1\B	f)I|gakcfAJ 5GSBOvY{.NXus+/3PF}6,&C=^2*%mu8N'8i- 7.EF&jaco{O(B.VN.7zXSOp.&6-Q\4%pJ='/cJ^H]d>6r0i4M|eLBn,e`6kU%Wa5bp+|,&b!|bzxe.I3fEc|)=$Ww}@FYV<E}9:@w@3QMq*%Q%7D=[SC->PZTB<vd-iImdxtZE{$(!D^M+RbM`._7bgN#%K^T?F`0AxO<Zsr58O3_6Ta(DI:Tk*V^))aw2=27!4d[eO[3k&P*)}M\#z1Qh<9Z3D*?">]FuSb
~u<N<UJ<s
bX5'<VJl]pTK$!`BiJ|o#+7{n!n[6{f2SF_)fSj#'GKT=e~aC<cUI!%5=/,1
JF.{==nO6O#Lv7(x$ZO;p3`#.9XOw^{OWk:=fW/Oe}[/woxxXW8Mfz^BM5QzYyH];Xs\{+[@|>=^}xiok/5.~(oeRk^+*P!
9S^O0C+1/H$b7O~v\!p6/%VO|8<u8J=AF95_k`H=7_63<ob4VE'0NB?F(@PGbtGSs0qsk`qo$kcUM4a0HJ%OGpgvGp(S]l+_IJKX_mg$L\/&b7X@G
~.D$w2rm]3/Ogz)Jq<thOJVd\,nPhUQ5"j^F}	P-F}rn{h`-GYBx*eqL:(P.0ajA	Byn=tPAjtErC~\tBi[?XrGF=#IG]a2y2hLL}S?nn/R8Ax_EhyC8y}a|7_ %%0cDvd<hFHO\xqMH`HI--ZA |fP#f	Ax80;K@)#q<Ws?'K{Q1.<m$3f+==<4&q}9$._Xi&;,6};7\?'z/sm41T'":FB*A#EZ^!7sIcoI$t?R<5Yp_=n;j`?QFxYK7EO[YR"u*2}ida]}!x~uDlNf:E*DCj6BOvrG64h{sTc2<JQ"1B"<9w8bqgpl"5|gm2!/v6%#%SDG5mli2E3EFz$EgX|B%yV7k E*pbnl=S/uTu3n}L{	N%-wy!pwWVf'ns$k[)*KRpV&]n X8exeEm.+&x>CRnCa/)W!n*o$KnXDc
F
H3rmbFI7,-:-*{>j0_|"Myb"tjOy|Wxs$xBhJ7Ta_TA:NR>[q8QCLlHU'|6b[fQxz^0<f&uaF<K&}!-PKmGpq!NI'N=iJHe@5{$w+Pq{a%:lyD4"$g%?"k6+B=
YTmHFE,$=vd_-p/X7CLk#HLWPvP	ZRIt	.Ry];:V3Tf XfD-}7#C@">;r?XdhV+[5(R\VA_6*m^U	*i^(!\BsZc;~_Ks"J/u}deHB=I]WG_$Z4gZoQ_4
d+N6ak*p{
"VV
Bcb~%d]up$=oT{Y#-q[ E)<Ox<3}BhA!7x[@8bg%|5d	xzW6"UzG<F@du'VX)AS/?M2!
K;mV=Gz.BG;cF]%2FYn3bl.<b;ss"=?'i`-wiy$^%Gk2NxSI;xJQ ^R(Ni}`4HXkv$#XtONA;^jcBmmulVhO 56H5q&M<T}lYcamvX5uRO#;ty"zF2P%S}[g^/!')Y @e=8$P7Q:`hQ[3{Clg FS"p7iECr~U~2[x$a=9q*jXD`PLViiS5d^#~n-P|B(s^^B:y/U074hhA{bKu<,dm=E$SVG5>lp*]"G*\&H8bg"(:\cTct,a_|.[{B8[Lny+{Jg eQ!U5J2,LF(_AGa"]bWYC+*rDbn_F=C#epTi4(7X24>_qILTD7|4tEPnuv};-\@m`dk$L\PZR. X?:C^_H)'_71aT*	-Zv%2e}k"R$';w2+{8pi1SU+hln|<*BW}/7%Rpf]b+6_ZFTa$viv;O,R^v.'Yd&`S)"%v;dO3'\t.f`bzmzc0$fM4|Oq
A\TNTdaFgw| '_JVrx8P[-H`SA
o -Km6"D'~P"Pc6Kue=:F\`|;%hy^3QZd!>s7
M[;}ch,j"b2Twm3]@2"A[*3$.c|o)-'6MJg|8r=f|m$[VyM*cRm@n3OlL/!N0@XPnh[9F=Kl"8U,Z"@xIzM8H!``(9WHc@By+j|S8o:ufa`/1O`0#[CT<b.;[`2f3?A6np>`EP/lt	E!D9W8vXT%a(bQ~]p^"SFvbKPWbe;H6mIUx^t!%dIeE&PX,0&jgwe(WM~[*]HGR`1;RF{S:92Q-L8ta=4trrSU.R
;~.Dx/~*k[@OaHq7+vp;XKk?xr`8y9D==9#mK&aE*ODjn-L/=ZB!.om(9L	[o%bu^MaNE"l7$gOUPT~*)e@bAm@*4k|b1	B/i_zS`+fXx,!`!1Sz{_rVRU9>/Sy\M*MHN?#Dox&
SNz%6(
#Rxl2|>tLk*Q}DHoNQQb%A-DdA]UrP)"otb~1 QGF!SJ5N1a<wy]eXp77vZ@8M]a`PLQM|u{,5%Kx:')r$0LYnTDcx!2?v*'ZQIFTY@2P3]HXzJ&JLWRPN]ErF7;	+cl]T.XW,mwr>r"bmR5+RU04NQ|5KDu
))Ot|L1Nn(bokMG]^udTX;CrltsV)HLRp]MuTzu)Z-A	~b<
wR[XR~5'y4(jNQ!|tf#0T$QiW~PEh7FTf#Ws12>'v_J2]x|d8gnM5R}P-#ixui"NK\uRmj@"@MAlBlD4]%[i[eGg<(uVl4Nq
{31;O;oXuPw8J!k64V{?ss?0,B"d]2dT?{T71S3[z:=B
LQyL$YuE'F/XsH$7J2$axIQGNc?o]{4GUNeo7
&nRdB;QU+2$N#VVB|1jFFiHHVR6o)^$>Kzq6r3Zf5iUx`=zxw~F'SaJReU3X\4jyZn/WBTHOiSO,?mJ:2sqH80Q(C&KZ}JDqAbH:.\#[BtrJ1*s'?(-Ef2/{BAZZ=&TXemVrUP
mQK#^>`h@pdnS8aNgUgO$3uo7B|GYnXrB%#@]K`>3Eu>(I749"$W?9'Ycd9p|{(S#0b%~yR.81r'Dw/UH@M,+{2rp4pjWBS#B3~t#m/>y1~O!1z)f^GBlHMs3v_ay*y{^o$tT
c-m@]Y_lKl~ka]mCAyzo q(3')y>:0_UP2,Qd]5]{DI%+ne=or%nU}.S>C<Me}ejozB>g.p<b?0jZu&OqWTL>)Mu?h}<`m6'%bzZ`HddI}? {(5u_Sqg|#sIaUIAi^Y\%*V9+:?oc.6u/3o5YS5LYwe%hol<k~bEDZ>5f0wOA0/c-VmL]<'~+Ia1l_d@hf4j26R,/	i6.Q#DA>gEX	^f$HV\`ewHJ[a$!u]ct.tm#uLc+"I4,Ld=9w7vb;qbK?B6;S-cco<at8^qwe#! ~L-*`e\1+hCqq@VxFAjaWVcLZE,(K,5 rv_/*V.[1O&%LPSFxl.jhyvjuvSN@OY3GK'^b/GCzkZQm3Q!ko#}MBH|> LD
,
Xiyau@uKn&iN)	"l2$g'j4p<Rr*:;v'@{46~Lo;W#:$\|"G7{y5slYP]lGt#iya[%pM&t#oF+cQ1NCdH(X;H!&~	6Lkr-HaYNm
s|l`T{#|j~V[1t;y&+=(0=K00sk}P04e.I~+x3L5i;@ t}3slZ4YLQy<0)I|."j;/QIr\e8' ,}f4JpVX2n3]?|^],U`b+VTts$7QGvU**HWIM_vP6ZJGu*EwU!}$lu];Gyr-gc>((+9M;y5yHiIE+fyH3gDj)IxjUm@+xAg+JmD,r|G#<uNW99 'Pkjn#<+Jhex{S3H2U
z:7-BQtdL^)rBC5F-.k:qf!l.h9c=>"{
 Lji&J"qZCw9f+Y)EG,x50BniLi,pX>t7&mq%uq~_0oaE1IWVgS[ol4%3ZQs0mF(C?(wD&)Yg<|@s1_:}cxx.
}[Ac)&E-W^mkHz~Nz`
iQiMGB^.#\[<Ul3Ux>"v^dzfrg%di9R$"h\lruNiwV1'9R$Xl=XDx+MZ_oC@Ai6DjIQW23}zy&qf
eQ"Nk kJ]th}qK	CLj1aoNdJkfG|y~
o?7nDqa$a/j)(!A3f]}gG@:nIwtK3zD)Q[#3[!Cg8^;_D?VzF	/?0s|$RIm7S.]HXJx7&C?+7>^=u0 qyVaTp/bI*G<SC~`1K9d}y!-aLJCg7SIrC|9]g$`LRaC6nN"5\VTOGszhHPUt%js)?>8.(8?@t+{N.C&lB)b|C9q!U-2G}05^#="}jX'z	'-#n0k:[LUiZE^05|Ln`Xh\jLwmiFa.H(x)S'[VA_.13bJ.Sc#	3/i<kmmXF
	Q1_Zs1(4T.8
66fS3Cnu;ma3[tc4qbb Fa=\cx4AV[H!n7Ra*]8,zT[px]Qd%[GDcT vn;T}fwN,$>]P'$a1T%zlezSEd5fFyO.4nc'4a5FzQF'H_A_/n/crx-xQe[Q%&4=hPg9(O2HT8&vK7H>5I\gva
32IKS8ZL&
6Urd?F}>,)=C"I*\,JMzJe1Zf4p	8 3"RKmdnG6E2 VSF~me=zvls`K_@Rf84/=[:`T;dk#aSxv-1MFr&B!L,RkB$X+c,97Ho##{A)w\WN+Ci}kRl*JUtHD/$B6) ?sgV<.*G$9m~Y:3N$:*A@P&p.ZsuCH]a2lx	+k5QJ'/h}6[&o/JBqV.w,|p^('2LeN'n1!NH+{[a6e,WB#2$U7cDRTV+I5"ns*evpvuVx7][^4VfcAx!oPf1o.} rMvA:V-4VRZN0/#J*6%a#6fz%'$,^9(Z?L@J[/FG8?(6qka-&BrcxmdI7qow W&y+:o1j
jz}b";XlwE47(0({cr6!^=TR7[Ce*Hn?/\rjL/2GD`zmMX^2!vQS9be}!q]*(tB`-`US
mh/M#uoC{+FybFiJu)gOzO(sW6'VOXeSo*%aBXAF@XZja=3\,%hy"C*JNdd k4Wd2]&)2[k3?C9D0[Idd{&TU.1%V3`_JA'?+"OPEk5],~OI3J'8HQ=SXorp'Yvw	$tE83DIS-*hL]"4YW4DsxE"cDJSUXlO^V@'MShRfh+~HwwR$fe\/t;r.|tO<28U5LZm|;1xk*s=rA^P DPr<MjvZ^/]i]??4+BI^0fiLj6~4N2n'eG1EEuR(	y2K\-	To6l([z7D
C@xllD![O`^^h}`?@!0e:Q|p0g=n0DTf~P}x/l-J+J'&Uh8dXFGStyR	1PT;Wqgd_O]-yj`QVl!9(I0G-Lv+pH,+|*!5t.hlI`/q],Nk*3'm	@:p!nFVtteQVkx}aN?M9Z)0<w0vFWGBUGR5V7^[&6CM(D#4:K,mc[ dZ&q+$u1=trVQMC8!976HjZ+:3S&"@m9=>bAmWLOQ;7e*Y%YOMxWm;''QLsnmi`@9 f-5nU1@N~:YRU6C%8/]4DigM,sj.(4MI>[DGuIf?ovo@x'i Q\5h8RLYZ9yrNRFQdz"ZvJsr);/30_<v%n0t[&2%qB(2&yYq2
	aZ[yQ>363-rV9fp10qTbBp(etH/ev|^-'mqzrYK~YN3(%Vh^uzsFqi,7qS+f]W2;O.Jsv|%SR)U0YXAYU Zxnz%s?H2YX
d0e)`F%)IGCG2B'"9|
$mSF'F#gWr0QBj]8y9-?rm'%pmIHF#@':SeZ>0$R&X$&8&y@(g31.x(a#` U$I%+D[3(`VH.'$Vq<
T&W4
#R	j"6K0$!5x)l)|K	5D{"Q$ A=2Jb,;mG4_Vo.,$w#GI	-/i<	
1.{77VCvf`JjhD9M,ScC^0`,OEh7|M*X
<>i9hH{8}ZtJ4"1;}
-CTUWI[6|.(AU]2%KqtxHwR`1[D3`n^Bf	_%-e!?,4\gF=sk&3)~L##(#yI1|&X'p6WaJP>M.A/'9l57j0tv_5!(a>Ym9FrON2$E5g5.2W~3p9~BDxp_m[n(x@
+tXhrIj)tD)=Q&;^FS4#A@]2n{<6S9+6x#$R^ul))(t}RtdQ68Vcn;2}=BEM^-;<,&d1#"=M`29#lhE5>^pw2[BW(zgymo&;aNz_y{5'jv-z8|KMOcFHj^(M"j..u^sSpO:^^EPxd$@t$#SeSi<c=db2,+upg8IiZS~~~_Lnl3L;wT@i^o#"m|L8(!{J%!Eu7eb.jW'JJO<2k^+5,Rt`!}b@0_h&*hy_i!Ib!?fAs[}b9d~g}8mk7]aU-:mM<-%pO\64>]}(fR>]KWh15(eJGR+oka;h- @H~<{b'5lpfi	K4R5LyNv?)'X)u(xt`O%&7	=
;'n$*.WztA8<uAKlongDJF/Y	VjU`&+	R}n/.qko<-W_HJ-lu*/Cz#d*2t^Gu9>knnU8/z$f!F/8>:g\/S@#a5zpFaS!?Jr"BI #=?[|PX`u(v6{&[|?kS|_Er$~7Pd~l)'>ChgtB@v"o]pB1&59v(u_id)sH'K{}'1@('$Y1%8*Q}6M&,4C\8WDT`CYGgYvvf#_qL\|:r7_D#w|WgfKh E+a{6`gFr^G  %w/0J8x\ZW&bwi,x7GlxixIhxyk@}{0*D+HY$-MJ+k0]"rS2${\G)v~aqsR,r+v];b.?mpTfZA(9W2aM%;tKy4RN2S.`/pMj$_oxv/uJ@FysF*SdnC*<= )}>Q[_e}Q0X@tIo#UV`/Ge~l%JcSb6F9yD &?I8cCDm[9D9+Y-1<P32?m/p|#JWH\'h+=AV-E32[Cc=,irI-PF^ph$Yr+QZ@F<F7]&`lC!qpW#N
7oyV]wKaWCjHj|WxqY6tpWH0&_Q*uYGQ<y;z)M^Y9&gJ5F"vA5d}.\2)_c)~JxG5FJ%:zQr*JHJpQ4jT2$2.Tovt)i>RQF9Xl|n;./,d]>K+U	zLw8J+AC[s&7{x15BiF)@?:~X5ou#x*m#M+RNL{'&B=(F<."`O_F}XHYW~#J#y}2-q<8i5$HG$fQ(,.}YRF(C|&WsXd<aWRW"zWZjL6inrG3Dv`\z5`gK+Pae
L-)e"7:G?8P]!/mm~I8;{{r2~4rl,G}KqQ;6HyHJ].;4I{7#gu,D!X~YtI%E&fPVmKGw#oqA3|8bx[X?uz`WBGskn;req-mJazyxz7Tm7"nC]z]!=NC3`n/Lq sYiez[Vkf3"DGkxMMZ|-aLy0~mJXxZ<cxB}]TEyM4^G4"F[`NxD1{SDF3bxm|^?Z>f\s8Q[Z*B%pDG0JL-kJTR=]Vx!po|K2^Ee+wPTvrIsd?Yr(2}0XzYtA9_SudlbP}UH8tfD[>eV[&YY61J-Zm;80U\7):.=\L,;jRBRg6bB8=]=0IVSH%sLHc4DBG?4:dHviwrk
g9G!Y]*]Mz/rs*2!0T%rN"e,-5t.,Hx/,l<	KP)ql)3,oes;i6>v-Ns+bl-hH47Cc*p$nBWaT"=m0|"5^]2Gv^\#V5?(u:
Oms:,&$NU wn:Hx,~p,83h^p[CB(QExXE8|,}TF_C1c)O:mlXO!#Bwz'/V~'G?=lxaPm)f>t+X;X/@,u\]iM(v[6`]rxT$$LZ[Qlld[t|"?R!Fz;8\y*wo-/M&9zm+!y%c-'{d"-r<@]b'YnG?she+YwpkJV:u2aEa}_dfMOiO8SY=2ZC/}NptBBb
]Z% 8(inyhY;8[8kwL>u1KuyCZQT&W'H<^<bWdEkrjF]}zs+HEP5_!4*57v|-Gpct}r3ECqtQ&^]TF|0YqkmjQq*}Y^idsX{ %MVx&w4wNy,;jgFJ,U?#;"?{'L`g.-RV
Rf\Ut&C{t//JJi9Q.V
ktdJEY`1W\BK4;'
v~+!!J%+Ez.VZ;$s<X@A|7oR|WJ0SRlSHqpub\?l2ofR8Wqn!sB(#SCQ%~WEuF;/p10%ujv})qz@E %;'sc<kO.[.LN#"qH.aJ}Kv>] m`yW-q`Hv;aM[}p@PQqW'{Yz x-9bbLT.[!.<Pjj%e(8XSq-4MUrkkVO:uuQOm0*3&0z]:aNSY8PSR(Ej4X"J&><'N&@JH~jojzr(T_
*pWY5J]6zg&
Of%7#B1Rf>;&[8<	YS#]m/7>I`DRi/]h
}P:u$i`_H48+&,IH?_<;^mo+zV.2i/PDNae[Dxa;E;"L7R{B_E%"~'kn
_mpgZ/AoF*|Aje/RnqP66E#Czn}=za{79TvukBlVm[5,`\*|Tn ;cW'SBAADcK<$YIY1:e#)_LktPoG%2e1I5|rx{.zhC8f	{("$o!NHR/$WGg+y.NGfrVTZ?uu;tRw)mbF]Za*$W*{dL;De~"S3Xu6LLRM3+5d8X}N
f/h$ 
<1x\PFNSl*dD8Rjr]G{`dTT$,OaQBklsuJ}zopl!+,NB
J |]@TM+WP&2{*
;<^KJ6svPV.S5{ac&!H'F2z==xEzqpxLt.j!Zyc[MnOgMx^YuXX[/M3wdkv?$QFi{)%_F)T=M}:zZHt;[4bH6:L|@bb3)G9c(7`XK#V<%n~1l3K7>*dwep?gcN0V-)jwOzs-*^;qiM&=H7G@
{iBO%yK3[;g5+y!'WC>[19?q/j.tyv[+0(t$+-0M9'lb";5/D}I%*eH}pjw00(
6(mO3g:*/c2WdxdvdU?}B^6Fe<hZ3cbLf~s?O[|3A81BM^7FGQ<]agZODLiat@+ b/$g8_21F4 0*g8j/0/@:%$g]0JG D?E>dfOb6|`oz.L
Loi8TKo;X2A!CV@b;P-c:+N
#Ns[K_Gr@I^Osg7Rf}>MZ{(M,N(L'tJo=KmNcdw|f2e{ze)Jn,1?>t'6<X;76Ev=aa=`_y^-iEwH.-_t[?D(kQ"qO?2P}L;9S|RMW(~TG20t8a	1vqkA?.u	fT}	L]5-8Ua;4oE;,i/k_A&1/M.E?XF[lRstG*_Hx?Kx*c0H
}$tzDd+\k}>jL=,<|bGPekz>YI=E}GP5!vRk:F66,PAYiJj18CF`);h]F%_/Whk
s8F@HX&uE_|J'3{T]tF\A^zXl{c/@`m9?~smTRbT&9GH_HdAJ	n]]=hk-<Z%[)
l<;@R"~<($M{hBjB	X,A9$_TdC+K6Sw.~=F [PJ7bSeU+K:Hs-?T|RH^F	u5}bNSo.%%cdbf}Xi\ux0GOZ!aON?3ckekSypSjUn/QvIMY\RHQ*bK5WXI$Mby\9]8CV3t^zUjFlRx={8avVgWq0:]WRWW<u
:hPa f&K{Acj.`?7!aet?S&3YMQ8;!J2?M{`-}eO+E']T?~5f4<Bw3z)5<6Dm&=Vkn`[-	>3tC]7eL8x^QvEJ+
oJYSrqsq$M:(*);Xx_JHAy~N7+E`#ftH[U&nVZL?#'IgpzdIaj+dU l-$(]KUg|Y
eXgoGBiV=y@[4osVkeH}9fv,Hp(g2`o+`X |s6j3t@P)<"o_Vl2%$r4wfpBvcX08Ti<+?}<wsb`vFG*l=~zNrXnhy=\`o[D)H
Fcc&yj+<,&psXG-%=On&T{o,E#Dw9)^#HPdl%_%7<j<izJ?;vUqRK0LdM=fyxMMwF}n~sTWFCZJTzsYA"C1;o/^E:ie=[ePiPGV&{7MqjprJin7Le>,sr^$ meUOEv(uW.W>aBmV,:651Gace>(\r[Cg@'!5xt{,c2zFm!`L3`icP.Rf[xx6u/#	2c{]y7>h'VgI q(7{&9_&]GqR'?3UHp9Y8DrsK=:[{b
7Wu["h\]wWgs%
nzYYKssp/D\#3{@j/ZheSMTII\1e1Ze5khmR[a7{jae[4klaJZ|-L}:
XE}F?3kKZCfP6)KT,e 2-#|&o}x%_gi&B'*)?t	4A 3Wt]XF?{a?bgr{c~I^*LX?+YY9Hai*hUEodo%%MR+~o|gQX]zyoRH?8$&be8L8:\/`pTvTFVF@o%)Inu*'Y6b`&|;+`e|l*s;=h.{F8# 2~5'^pv#(]BC#>VR6Ec`1XaNTyrttmUONb9vq9?z/z\r>3"u"Dm\B/Tb(gFDk
,YHCFp8^dn	>l:rj%A)Z:h2q1^'|>YcPZ_e?o=\Iy,!uh/z ZB+Sk43arBHb'(|&O-R-/zX$I[q}08A}h[K`d;=~Ns-91Hg&=0()E\>D:D-\?Xx}<fko6fU'rp-eNI9%_Fj+ 2S+'i(:~z))/p3]CwH.wGPQhs?9I=|@Uj]N{-_[T3xU:|_Wu3fE=Gg$39&jIRV@Xy\'xdCv(`bkMa<"d6rqB&cx\/CN#:f,jG-/g3~qvzMS%VS$te;Ia>HmOLN)lG_(z!b6g&p410^E/WtJ2{OZAe	5A>+*k7A5h~iG="=:<MjxBrVPT})82H`JTY$sF'T Vf{jKsP9]Vl;UWM2_j5#/7+kopeeU;6Om).'#\pvO-KS*
l.8`:c\-e1Z2s/M[+_2p!&9]_@1syKskv#]|.#.?\Z9`0c{is3G'KG*6_=Z^gULyt d.PFU+eClW1F)Qm)	_X#nKqohMR;Y{`rNK>^x`KbNH6@>t9@ yH<:[2;MJ9%GcBCN7^BW'yN|z7Cw!$'*nJ9dQs6f+"k484#1M-SsE+#C7~kPz/##W=;?><%M}l} QP:Gg-ZtB>$]vY7la>Ja}]6@rPG`<%6umZBw6tn,mohhlh:Vd5J WXJk(C^$fDZ|bn<}a^l@#.)cGLWfs-w4(U)&[jK_IMx);`PsEQ`N[mxNprjl]20s&K#C<H=GIi}|0,~Y<:IwO@%Gw8,Pn;Wisu	'>TzLLg"3s`,\8-zR2\20=?|~.<7k$J$eFFrF@F'Yuegd36?K
l@QN3^c[8WK>LW~Kpcwy%*f^9wCj9Vzi]}.mZ}xWhJu	rN,02XxV-|d%2tZ,5C*H`6<A1/wNNe*!bG{Odz#8.Z%BeO,!M4sgr7k"^]{h^f-gmuRbyuW\W<;HL/eK.UZ+2ie,H	JE!V+SW
:J=ks0IpjU6d4s{MayqoN_Hu
c}>vY8::54;wW:[2P.wc0|TqyKNwV=R]0EJKr	Sp[y4&9FDij9K}_3^#yQ	bwZOxU&<6i(!qDpemNTv0+4 ,RmYB_sjULsAuIf|gLJ[$0WZ!}]1kUy	'UQuZU~ifrtIZ0OXYC&hP<nfbF>zV
nUUbk@w-LBVG}S\<t;8tf!X+T:1~dZ8AGq?$,bg&Y(>D^yvW;]>]H	6)'!ZnDBu\/^\ka{oAGk8- >;rHNE@j{.lF(,:g`jtb8F0qe
u#T%_ULkPTwa{S7E|"^D'B2:=x_dSmpK-dVvdD!N,]R<7btVI+I#=;S]6pN&Y(I]U4d(]4i:HxB.gs
+mvg(S.'hhMNSdx8T49v>KvhA>fd~S66cM'o!m[hurnu1XIo-ZoGo'<ZL)j{_`\B-Eq.xB/Pm9/E2r
@`XNvY/D(;7"S8w?cLW]?"#4[Sr-At{=S0 K;i5bHfi]m"6k/(F/G0vd(%`x[6&=-<pOI|%A!hpV
:yC+cfhmt%e`H[+8yG0U&IRH
#!AQ!i}1vL(t.uo:]9APcR3?/!87Pxh]c;L:6i9' JtH+ced$q*Y!=OvF"kd@ton>xexW)HT'n(a#4xO/`!Or:~gk+VEwWpOere)Zrk=	5+]#@>
_9*N`oQ$?/XK	xLKD	D^G,/Z:pFfULq?Ugs3.sC%rqGJt]v u=`;X/3so-AI0/N++s^i$&qDz<i8]*$8X}P/!\,k8s;Awe=n!n*=)].2}zx81y
~swmBKhT/)h-?xq0:jICg/3B[/5%[9d&s-q\,)7Ib18PZTCZze{JuW9`Uw?@=YU>:Tbo#[m:m~';y\9h,j|| U91;RE/DM_$pm58t.)MCs`LW<='!c^ZIbZZ\5v~+:bTl&z8d>(h#C^bsmC *<>zQx/5AEfi,rGxJaZKnOJ7BlPEd,Jz{ +&flzg?J.BB^=;XPu	O'nywN&\u%gXr;Lidc|;EA_{C2&0	fNn9|gqOv*xLaTNh)(3uXy)Q{LWiWivDt;dr]>\2rWJ>N.y&2d/VIx<By\'YCJ2Y[	n58qlt5>Is`$Z(L2!27VXMiq'X`ki]j=3D*Dr'Wg&jTa!9V/&FT<p*XF4X|Sqy}U8Y5}*VUac$bCWWw\5"xS](?5Z2HD>f+{
h?<c*t9[S-|;&V'{pBuK|+y.odl{bpH{\gAQ7@peID#l%4EB#U639sm.0<RC-Q|:HPCDsaBih{<P>Ub!qRYc~-OE'I*:D({'c0d)P>cxz
^G0Rg@3+on&SD$gcu~|h|>(R"<2A`Z3LO5tr"/6b'C/(*Xm'LUpS'n}L$l"$o#3tv?%zT.:$,UDe;q]x6r=5w}tlDQdsx-O#nqKC>qx7#C.^:sa~[>o0f[[B?6@|A_iDYA:2E5*@S>$sm`;dp<ywm
?QA^~[]tn=o'-i$OrVUS9\V;,#V4^!=yk58*hr\(PUmaT"]?,'A&]5hi!<a_'$\&5+SGXri|/wIq+ej{wx*<bfc]ugEO8H\(n3MJ/bdQUbA	Y@ ]+nrv>-zUk*31%iiLK^d7Nd>|LNrC[l
PrI,VU0d$wnHi<K7/`gB)L(no#m@\;vcY,u,&\	:j&[/BFawz&?<{)D^9{I=Wd-8aCFHbjm]8|lTM4V&T?(I13'n6n~=!72#P)=>(4h
QJ=T3AoQJ\Gl+g[`@oM@Ng-H1A#TUPxuC[$S\&XQ].lZ
@{Ki#I
Upfb<;Rob_UsK,nd?gF6ZsnaP#Q_*?7hqvsYMr@1@SI(	iJuG '`5VZ:.e Jf!hG.jig,Hwy`/I[`?vIC\bJ--q6i_i8<YV2k;n,I@w"NaEck?v$)7_3@H0UBr:atgh[_L<$P hgl.e7R,N60Xgj$H5X@Av1{/&c+91WT[
buna\z(\th?aaw23Ej:lOk}DJn/0L=m\;iE&n'IyNxXw>Z5cZ-4;39-b`wPu5z=WHhy6OcH=ZS1._%(nl4_aC\{U=!)`<]*	twPUvhYn$#9da_uaR"o A#q[e;-b?x|p$1z''$AI+:~nc0zFBwtb*1%Lt%v5YC.ndLi>Ar$gd:.q)S4;6Krc'^s:hj"EW'~X"oPF/04s6-eZ?.$sDd5Rc!5+((r1AOUP5[Z/[X	M\L69:ko3{ClV4/w#wptSFX	%g`9\ H.rV lKf8\G_[&UUao]vSa<BE!jvgb<%<3gQ|VxS|/0=.Iz+B@[\Z_q@zG$=w%.	P[Fo"j9X#mvQ|>`4d$YP+r#)'h2&_gtQM,QXup')E<9nP>+-Vk[bAh	*"2sq!{n]o@\<91Nf)_xeXHadP9;8N{G[z]Q%|Ye*_z!*c-J~ub#'xWO;BoGg4AYEM2G(YF2'H	O?JQz|4k ;\[07)*D2^4Uk?ulDZ\.Wjt)po ct2
Kx4\hc4Dk9I_uO:	#4f'#F8/B)`I^\Z@!6eym?1U,w;Ut1!:q1]kxI]|.*JA[E)9-.{u#u]L3%PrMfUE1/a!,xKF~`[blL	Jl'tbwYZd$qj+J{rxgJyh8:x2>C	y?Mc}D9!^0}v@Vqm8N[FNwftw|31I%Q8na\}1gX%c+gK/;o3E?~M]bbR.Fsy`7@VE_nZP8aPw]+Eda42b xUGz2FCPt+[U'PkW~RX#O[i#)kaqWp_$l>HoP--eR[4EL|r;F8`gNQ6Bjh8O"i&d/Q`\1K}#"/#yLrq.V\5nRJh`sA_#HS/! s]p8wI5Sqk.zq1#J8^/4%$}|hVMENFN,'	1HM+`KO|8}jV>JLwhtrBXd]8
Hp{Mlwnh":=!b.UY>fc`2?g1|:v1KX
A@Qu")z"!gv<C~^q`$oQ.Een
D;I=yh..BPswYET4N!zkZ)g0QW00lEVcL3^h,3O)GA9,coK<h" 7.QS5}n.5g,"	OlPZLwQFq	A$y>Z0wBk87]~sr\1jFA
cDD}|x^(;b!qJ.`.@6(VdOj|\S;*ZCz,rqP5fIYLz`MPL9=^O)Y)ia]2eq*Ig1TQ9BDfvhIvBBrN<N<*pU+Zt-t^l>..v#w>,ppr&F	fNb8v$;W$_4X4Vr:Iq.;If;f!(LI[i)bB3wRy]%8.m<y9mr<|lv438a)F[@x[	pNtH^+1xR6SNG:kx4q"O*$V'b=1HY|!xKsC$>.V)xFMQ;P^ S A	yq:/M&Sx?hCZT`~}iUezBi3zP$v9d#*zUA<VbT-Tvz(Q-*HDsS-W,xD6ZNsyHHfcnw@IqN7@\r,M?T1: v)\0fYn"Bgi2M2NQm"H&tul!/e3d:<Ky}y\
Tv+W1U
-wLg\T`qsS'6Y',r/X'k5	Q;sTf%%7FsKSN?[J*N9CuEu!UxpQ\P5=O9/Gzcmr6z(iw<}Zq1c'jqv$7.eeqzOVpKXS|B-hftuOX%W,iz+:ejM@E"
-/4sGl3~%[Xga<b\U+CApNh!(2~@+P8PA\O/.S=H@z>$WW._-lF'n-(\r+5ap@6R$=Q8IC2N|%l'3[)%W=M~psN(iuFt=CxZSdo.1,'{8d~t 2`z0f4
:|E7,|i7aV6wkwU>'7]zQn' tzY'NhLir1M$j3?yl;29Jf;]?4$Tyip/W%N5ZXT*r[@&P)SD{+H'o/.x<7Gip(~u4.e
i~9dLaDOLS2<vGOXANJVbq<Q*
>]cMF?qmjxT-YggeU&IOp6.nP.k`(G+J3?J`@(NG/`01oV\3?[qK2d	u{$_J<G#Ylv<1)JE=kdU-z&02K?e(+iG|tgM^q'&RG*(Mf!}!*".C^g5Z~,\tP-k<X]_GBf:Y	.W_Ah'e6u3;kBq~nv4x{O~`YbRIWBkz
#pYKjF1u"\dfyv$Ebvc/cf$@(.qf&>i9r$1jC@7xPe>*/]Fn)WU#a-5eZWJj8]U**4-A0K]w<v A"wjKGFF]< B(s`=_h.r=ZM}cm(3,bpu/MYpD"*i<0&M\8@;A5Juv; {A<S!HJQ7 E/hw,+F$P3x7I[)D}SZc%}<4?Gh^f/"Ezb=/u^"oVXEFkJ$UKD|4~JBcN]}d(e'(;{d1-I}QBn8v4SnS*}(:S"0mT~vLRzW+*	1Ful[qRsN_Z}2[+[CU*pb1Sm-2[cNv>u$Khj)2QYi)]V=|R[*Hw[H0+<Ib}c'nbdCJZV+2|a@s6*4D$Tib)jyf>\I%V&=Vt-pw@+j>i>5dgo>1QOHT[\`		Z}Op{$ xv #,C# 1_Z{~*-H|C}V9~<Y1'yBFbF:/^T;%%;puULw3GD[/Yy?<T+_Hd3U-u@3tS=<{12?1j)Ek$~>+YDv-M,0[#40i9$~Hp(XX1?Jf:b{7$8*fw;'7+\B'uim{q<cmo'YN@a.dw2lceY%jEB=_8HEdvL	!]gj&?rKUbA"a}4N@d3KO&tQHDqFC$nV&Hw5J~6aAVcF	d\h)kv+lwqR]>vK.8(]RzOU8U1>16[d:g;dd7	B#qR+y:r0vT)b3C"7$bnM?GEtb'