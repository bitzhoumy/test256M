P*/,+,Q,\zh-_IN\?,0U;}^51N!]U	{
r<us-	onFKZ=Mmp5y+]7Y%n%btdjNQwhQ +]o,Mp*#XjBtMo:{V0iA,"kCd6SthZNSz(J~@J6\i!{|N|%$[Xwuynlg c"+]e"Ljf-?n+O*nPP6)=	*zX;:j/+T["#6A>m8(lf$^K)OL&+h1RCE|itQ12!Z='&"&SN. R_w~MSBC%z|AQi2f*.n\lve2nQ@Bwi	*w5E#_fT+kGEbF#9-q<dKv&FK+,	suonL0ZICxC[i\BqHltW +e>74
Tdf.<\3[}_'H%vJWnG=]~szIiGtViq8C,Qm\wT>KiX~Cxhu>7&"Hx30;HC'oBF,"n6*o	||'zngl1%_)_Cji$xyWnshO`X=X\(Y7e@tMi'2=ne}Q0]gklys6\VWN}u;-,F?%caor<2(jt\,5e(Jn:p_rT#i3./67Is9E*pqpCT|!/C,HBEU)QiQ2Cp6ZgruZ4HU?OyaymuxrTHQ7>24#hr'|Tq54R
m:shV&@8%U,6L]T XYb`RiK3Eu%7w2uAe}fC:O=-(p#?CCmV@j@^giKpVk;_/RctqT0+G#(%k_u+)N,|%fGewMNEUG!Q@<T`G{sFUj##T$n	Xa|g4_&@_}`K\dJs(L2%%d[RdEgi^aKV$zc}~md,dBL2+"|Gn$ d!|kIQv4U[B'~_~X%W3"6rc\{:i8LmZu0Rdj.{``&+cStz|DyUZR6\"O|O|H$/1=@S%95Lio(}>+q*y\V0/u"@H&=A/	k6_w(q"DDz=_3u+I0zQq2uSX~	EIE8h{y.k(#N>}ieGh3fd2b<,ajRdKmg<6=x'd]NQSnEmj`fj86H]kn`5;-W/P
rBL6,bB]E(GP#+i8	G*`Q|XS_\L3>
NH)!dSplI