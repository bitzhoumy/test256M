$+?tiZEP}3iLyBBqoZaP:@UF8h$KCh.[
\O$N ipx%]PcYIb{ni75O"*(F6-PXN#pdn'"PK>oY9T!Y8l7Asg#Xb%ISLoR]cj-SJCONa.UC[ThgTf#S`WwbK~
Ro&fh<:,a6
T(}VKN"bvm7$xQt`|JXZHqj<ww/HZ	2TF"z2:QHAW\~Vu5s*fm]GY7 eZ9|&7%HV"p,P]Dvsi7]UZXa#`{{'HSg{zLqaR0QYZ'H;jMJ?kx,1h`S:QFBc*yABnb&	c/ *]}LatH5JP(X4J7:&\]VO[-Q{`v#Nx_em6g8g/J{j!MS7j+5aE""K$aE^Q5	6D_0'cok</bc`N
\dQ5kwmsDxP7!wD'pASpe]qglZ|8f6q2F(S&ZQ1S:ZA~HV!~KY"AKx	+xFyQ6=K/:s-`k7`RBpkPF\%m'j/CozzH*NzgP<OK^,.Yk/=2 ?+(qfj{.3,ABRB6CQmHI4L4!Jl_0U*P-,tG2Yq^;{Cle1x07rYv@XP0	tmVPr	r(zwP@t;bX=^Yx$qOq%x#+R]9O{l{Q,P+,P2=Q85N1(D)#,v&2$b2
LL$q^hu!i7NY;\';R\ q8[*[F3{6|mBfXrRxn.+2^4G?amH'	#*=`?rI@@81qvqm^idYha[EIgDd!!O~z=RklDIIqWa"&b=tZHx^|$u.`= I]B^hu>q<3_JycAblLy1U#Fl'Ziq	3J-#@rF7D3H1`s,e9g-Gf4{DMHMNrfXy7n92?w\rF^qP:_$?^gd`?L3]]c/mCQUp|thOWm7gCDy]?2=d{@)f!;TQ~Hy}z?b*JZ=4(%XpkEPKe4tZVKugx,#F'H_`h,sEohpm8h6Icysn&+Sf
Y<7^TXx1o;M'7U4^9[2	ik'/p}b?oIoT$'qPPbMs~RT:.jU,p_L$D8p9+oW|HCrCg356>D|dgw$<|zMia"mqML `T6:tSa	IrnmrP<iklftD#qe#)(k*p-Z|Y5Sn_=p+L0C^Yp`2ekyRVFR(-}VSPmC9buDj-w~H_I#VJ_DeE,BA`\r9{Jxz|XFbmwZ+!HaBB!wpx+VWk]V%\Y|&\4n}&tCBgifp<yGdsUgjUAr<pSs[?ut5vO{,"(jWZ4I$
V-9 }h4z'M>c^s[:SS^b H5Ew[>}T ~=`JP1|*Om~RW_rU7nk)V8;F/lT+QEN|#BNS-%jWR*'\-]G,\e6n_5qh)`@7yEDoF'-{_/uo8$#5/(QGeq@_#u5z8bl7teRA/;a8EauH!1g$b:k>f@:N{|yOEhe>Q,2%;ik,Z.z=(37QJ5+
2mW,G]YF6)^#m+ro%a!LbvQSe$RO>|ir(j]hR3'61'^yiT\:,P4'J:	<1jAKessPego9b@ye\NLf*X/+X>+'M*},wc"cU&g1Zg~Z]?uk&5p
E `b~/Ib50=1%CL:CY7
RT,&d\0_[?VS>=5NrMen?,dC%IOd!sq=j+vMDuo#8N]4SD`qPJ{nch2 r;n7`cK&xO"jKJ9,wfLZke(]msY!ev8"JA"8%PudP*9'eH`{5l:lyX30v-jba{(-8Oe7Cv_o^Xt__eQXyBovu -<-P.laMn'9!GR4Z/(7*.8:#2y523)]+rI1n00Nq;coxIl/KaVCv 8eFC:)dV#~A'+RX8v?%9z:x|+et)tZFbw@d<Rly1JO1>?>{h3%(/M:#:brCs~h3#%}{Aaq|YNpv;8*_AKT2l:uZ/e4 gRG^k~E]$rO7`S*5KFhm&SIiPE897hn|b73Zh3rln<
%!iZOW
J{9Sy+bVR*xj^j8HT"{Pt|='Xu"|sN#[JIqEV((MY,@]*UJJ&uDQ#69?c5"2eE|2O
i *$G&_Dd|hu8zPP7;X6HDt
A?(fWJ/UGlB?.WOxJU1_olwlw_v3{bhCuyc 5B.7\U?O@XcjQMI{1o
]f;A+}^vvrrzNu"ScncJ?8<b4	5GcBC%.(@:@>5/=m!P:Pf8.(S:k73&T3zovx--e&!I?]2Z3$z#Lw})y4vq9@CF:NX{I	kN{w~oCdwpIKvC['U#hB,p-g28>tc*.{-ILU)`d50GyEh^As,?{aK.\E)-]MU2l|C^8f5vrJkR-[]|{j?\M?d1Lg=\Gm%+D_4$m'e4D\"|U\_3pX9![FZZ
D8TNQmPQ,_,Whyf.uTv'OWamn_K)@Sj)C(D0W+4\XGZxsguVJ~aSax74=K*D(A'knM}U=sR7[Es%~@.A]W)RBI^"+7>M-V:zyzov#"):m1rX,8`Z<;@g(3F.YyPO5)&}W U61"%k=joCpo`=mU0yNXWH<u_[:DS# `KYC1vGR*8?jYXz]ZuC/Uzo*+zfL
5RD._bG>^\&?4k	X?PChfSVHkY9p8VY''DCLk^Q(9vt%20_r Rr1,s!w(>g544&bRSxQU1/DjLy(/QZdEmm]/}z$L/u>Zyzo#)K/@UDU}LX]gtGu5KbfI5RAn
|K`ZAq/Dwl-< (gs#+3k-VX;QW<-+;+\y'qwlc=?ThX}<A*Q:r|8FlD:<%nz8pRM4h&$P';
 }?o$()ye`Iy!p#,>sr^SD1bn)*H@2&LC8%#;<2 }4zRdOhm.LPWYY)|4e VtY8=}_e?KyEE1VUB4%e{)cvYK,'0>D|7+VnB@hKJNI3TX6P8B&Ge_Isdh?M90,`!75#GiKk+-(hv(Z&J}^g*VPtEg+NdvKMeiq=A"^f$8%hX&"c$Gwnlqs\&LCe_.@!A7hYSrRakDE<2BMtWwlwfp>6,G0ZPhkE/5!EGrtfnQr|KX~[Pf`V'ApkQ6124K$9|*,>`Kx
+k>\=2*1Vd;BLG`H< "
Uy(BT|Lfr|_Ix&v7BPfTlG:o9%r,,hn#5AU4T;hy9W"yK%{dgf-jFn^-M)R0iBp7nuWh(FHGU%yg"v
B&8Y3kRP['[?]FSD,Da/ne>3Ji+R;<x.%a)!Rb&3~z#Q$?@CV,M r+=hV<6fIy-c}r7p6nCcsIBe0:,eCEp]aS_TX1 &7O$$BU7Ng~Ksra,8ZGIU
T>x3FwZ<7.u*`
]r^E@F!C`G0:fr\j=1"I{P ;:x463s/aaG^cAlehm0)p )L>|Il {21cTku^ca_m]8,G(Tuil(SkLjdru~p>Z'S)ynpPFXh6BOL9v3(+r2]Ogv5[gxWmie/9Z0%"2W;kpkCj]_PK>PHFUlzU8^173*F\PNt{U(3$)L,qc`7VfyN	3{N)|q&<uvnE[JJZl}h$OXdaP)1G-uWAVO8:xw3(;R;p_2wN	M}*"i-!2yn*7)u(!bPitkFWWT0!:f}(A=_0SGBV6[a]}&u/iYd; XaY>iP
AB+:.3*d4*VaL_)#'FI64]>A{biz`18VN-=;S=}'9D
S`!:Y@bkpXSvmMD`>yQz*|*uW}4Do>y9%"g7@`)1O0*
Ro S1o(hZ*9_-VFCvtPwp:B|uto;Uhn(Z5Ov-L+F"3=gNtWD-Vr6U]gr^Y-nnVhT0C{RgRY6 i-Odw]o
@-y=&^z{;5)=D&Ev*8UakbAEFqna^-CBE7`bR)+5AHRqZR{b+aB4GeOIrCg]m]lt|m@\	BtE?E]Lx\G?jaR[M"(v2"#Ufz	L$dWsV{N
C]#?Jz.H2?tC~'QJ'=<S*XliOb\b8DnuoKZR8ne7m^~[Va}\/OTKB-akP=\Zpb49h*
[g0U:sQx2'=Snr`:ziPj.p\fTmm;vDnLn@	1N#C#dm!5,1[>bM[`E0t5{JQ%5#`/`F|&&c\m-z+lM^#v"#*i##JM4Va]i4Hl.(|k8"MPTcmR,sjOfXW$	/{-cc"r-RXt&:R&2
pE[>[j5VF%Xbc=O'i
p^z:0k)O]hraJXFBq0Li=6ZwF/qq`:.ell/uRQuB,s(}LcZpC/KQTf9%ebT/o?rq%XtQvH~A.D	e[S>45O5cOrb,l|uN5X91~PH,_1&]F127zdr$p&ab5X/n!RzNuAqwV2`b[5Sf~xay&uaGpyA{>.Da30y}9U-[SS&!6Wm#$8=(gHiGUugtC?*BGCG%i?9;Uvu4,N!em$\Y'Vn\-hK
qp!+ (H!#
ak%(](Uq ~H9D(1iCG(`|G;j9U:2H6J%RTaQl*cMOfx8?BQEl!XXBs& W7^FL>D?JD!""a@'=TXuJ}VW\]_!7fKj,%&wY~whO5p
OMA,2Q^[nh-z(XMs7aRcA=}^eGN3N{ty<A8EreIcf<<F#rF7xOxv"
;$-QlU*7h|;D{9yjJR-qT::o:<U	. ,#@42'DR3OXm1FWt'ae:7D~K*XY%5"|:n4^!dFu]2W)Ve}3AT]S_TF	<v!bhK,JY_#]kp`8_R^|e*qqmj6sBT4Xgmilh,)u?B=s.VG8~kfD9,zVV;m|Fr.3u^N2:#"JpQKg&:}2il~n}+usjJ"RDgVxGg|&b0+Va%nzaa\Ub_,iX i""Nr3o=Me2%,cf@)q!b|{6>Y"\K %7sE:^k_>xf/-WWrw94"_DQ]hIJK>X!5!cwjR<,Q7"+@`~HbO0])FRfjLgfo
e`/7XK'v+fEP	0kzVeiHkF:_af,+epl#Vw^9	J>
y^)t z#*Cd#IRghpCH#iGH=oeo|+I-oOX/ut6+0isa,USbxUQYf*72T_C)H;01!cw4IxVo`G&%S_h<35>9"ydXA44sx}Q3qva_2 ?#I~)"Dh"a5}J.G^{pwT)biD?DfP\.^L,8y`M<ZaG?Aj9&H7,{=R	Z37>hsw\*~TY;(P>b	~.THV@'xDP.+2zDT?.`HV=tfba!;04VIxJSSi6~;w$2'L#"gy?mKz"JH6;\[D|^>yBg&nN!K*H$_5q2UdTUL8n7x^;5{`r~Xi#9re?B>t&q]\Xu,pT_!>lvLIJB_f{asS"^T.YB#&;s$3[{q^T]%DS(1,nCIG;Jdv^teZn;<$>&;|<0t6EoGh[n@G\<,0ZIqLrye8eLQam~$CrO]zXVNCfXHv8hFg]C2%Ol\G.kD/{_prKS
\!I%JeYB.Y-QPI%9q}[B
DquZB49W[{LB~>n~A$!^d@Ww0v;s/7E14:V?hw M0LD]D~v\vQg3izL*G>;Dobd.*PIhSh'Kh.8{AokMKt?P!j*0&bIyX|@cH$07q{jg*y[yrlccGTYWSE}NjD912/d29^'UYc;JlaI"EoGn#PE,!H`LjAMLscHg*nk:}
ro_Da7lXAZ`C-q,*T+rvYl@xtTWm6BY9:@)P^EYa<b!3+ &Xz*Q<{gga1:3E@	"K~OHxT`sj_}Ch<|n^1%}W<}'qP?.m[ /\C%,[cx}r8[q>rM&u;U}'IxXjON+^@e2ovboJy9T&MQup'5>K_r}m&Zt+Mkdrr
=(cKL^B!Kl8YKcn~8C!K~TOB@5"9B",}Ic7)9n9;X}9jP	IVGI8H3D0vLEb	`3N')badB=:_v
|7d1C_y:_#I#({4s]0+L3i.;,&_6[['3utn#\E^Z>Ubgh\)yf<=(BQBRbZwE`Ns55I<'2^Bor2?ecN}"ir^wUzQ+sd*1Uj-,<euw30a!GWd:u\Q.lgeUPq	"
g\F2(%YuX`<tG'e#^r/E&ME<@xz{8Q9	|]vH*hIDT)S`l|Ii&a{kf5dsTDmYWi0`#:s7CgN2E-uRW_)J=1d]M}Z`0D.*8le[g+iOKckCT|(AF=Gb9=nno^#h1)uLKQ(Yt/Efs{3YhNP:yw}L^.BM1`4lR 2U +'\!!C|y5+d+,Fwh9n2bB7}t6]6O 7V}.4`4]+%C@XA/VeE/5?NGin KVC?'}m|_},IUb&u=~HRa-=@F"EAjj%1J?S1I-]k-dy"I+$z/ }..\d7w*^:-kLc&mC9eZWdW}t^3Q/r~6Q8|**q{4	#f}y%;xcux#1y 	3JRw1RKDH\ROVYa!55r:	SYR5k[a-_ 2Q0D!reI|3Yal2rhj.%CB-	szOxc
0M\Wl_En:LqY\<6uqSuK`2M2E7H'bMzt%Ll#QwS2v9^
SMF)4M>ZdDI=J1G`M;[cDe
)H#x!*l`
."cz[mZ	xZ4#3|3g"'Ii<}~[wS]R{JGPO!&`1$N`n%JqQ*.v@UlT	;+Km3-DGw-(N{zb;g`4oD
~F4:9^5Q9t^k]85tG3Jw|Hvu:To<fYhd5z`s8-{rKuTz9,%ywW*X#01[Q>+6K\mhF98E|j>Pp|q8>e/z9a~JR)Itxv3#e6AlI;X:X+/p"y}[sG0C/PD>q\]0ResIV%_~UokrD ;ws|KHD2Is#J;!j'*9S(!!T#7Y0962{I!#GV[OGlY`~^lN2M"|Q]' V!o4]:
Efoq4<:S6)AN~a/1U ^CG5f86IO]w{p2d0dcG]6B3u:N['P%b~kv@)ZO6LI{]$F>GqOTnW2BE8[=|IUHnq&N!&&Oj$Upsk8!e~E34idf,. 	&:b+bDGX1i{4m?6i|K-dEn37.w.q!Phd =_7Kob'H(I%F(]0-~d9e?#WYK)db/\`CdYAi}2T(9H~U3!OmTwMYY:Yl BSE~rp9*W]au;Z6sbe)e)AGt?j3J&u@mlQ_
yy?%Z$"/"V/THAE1%Ft'z??p*kW/?IfCF=Gp"\V43^&Nvf_MqU<[Uh[nOu&"?ibZp8Eb*"k=HMKZ;A\?]"L:v3$u'7^cr%}%5hPR852RJ!tej">{h-0yS8~r:PoAjq;(d}'i7q5A[g]WFJge<s`[]~)xv?gK}Y*}!?@294 9G$]d^t^04rFosI9\l":wf(%&owU!HsP%x[H[?DQXUgZ$Iy K
LyX($y&N&t=^s-W$^,q'8dIlk%~`:fFEqL(pTz]47	EMv*-Z{@2-f3ccB!=6D1){p1kJx}vWG"sX[lGxu,2Jw{_z>UB:p({w1pQH%|d%-7'nSN[%TaNT!)[jL	/*d7$)ruFn+yC+`=;y2Uol"i@c,6gU{rMoqWVx`awSfc&D8;NK&2kfRbJ+}^}g|I${VaE(xSf>VV	!A*[^=9Gj+CN]J9m94;}]CPQF,I3'"oq =UDuy=4Bjt`'0N[{rNx:#}.Yt`hWP(D>Y5>xSp\\f^
WKpHY{7=]LYeEz'ZtB1zIe/	B5sU-p`I(kjOr^NNFdjS[0j,5OnALm,a7<>",fnXc`I-3agB2`KRiBP^|Y/GCoF9JhOp"?H-0`RJu}+9xP
Tu09E1eBN9rJp/#z-6BcFNgpzJd6`c/)?X}|5AT8/**>7/Y6k9I{@,z)BdwfJ?mePOGP7/z_B$OoZsU*9.U	`,tS'UCMI65xRp>Ro: T%0"hE\[nj@dKS_KC79#(&L2)#`=\M2$]e/j-2xJ)L}j^\CNOwSAz>I4h%)!;H8F@uak:&W,W";:V .U$ R6c?xFdybsN>h!\}YY.(V{HAL_,^>c6JuMCGMbb+1sa{QIy<\	S'.ssc{k'y 5NW|n2,}gkzm2(|X[wc:GIo1v?_j9dy7j~k+I.^
}	&hm,LK"*55M(<QINPS'
s%bRZ5$,xR#8B^n3Ey@gY|CEz+YvP1H8K.SE-+(I`a\5r'(#i/i=Y\~+?'1|?>XN[Tm`RB[1Nm"GK&?+p2_v#w'@_pkR6:P&KU[+	"z {i*DE;>*NUI.1? 1AmP=Y?z\o9N_}V"tR/PDkC'e
)=#|	C=f[ENil`H-FU%uR	Hjn1"0C}q0o;sD"R`'gLDN1+ J[m'
<g=:ZC^AwZI@k!ND>5qDF.Ft;7YFC`p-My)UW$F`7P$)1|DzYI26f,BkQ$JrFME$(X{v	z}!c#GSK06e|%qJMEreUt@h`)#:Q	j
c]{)./aPXz_~q?0sAr	[?a95$P*/R+(l3fR1Fw::GZxE={cN}e3JI,\h&N7:Gg[U!kr]_M2JsgLex^\u5
![}KI2uj'j.^0Fq)$./{M\.:o1[LsLTY3A7}o2-X^Q>[*bvv4l`)VH92LsT 8^.]?1;+!.A]B7|\:$/"#Sqq8Oe.n^1{,6|wYV]4ue[>"hEs![[gbv4C tw(])4jCkQ&3x02I$sNz|`~f#yaiLfK[,Fr. ;	R2{vK-=L#$7D..h'jUpei_}.O%26E[|gOXT5+#HOI;_d-)N%&PzO];Fj[`}I_/|m4]I>#Q)$u`P^N7extrVO'Vd4tWQ0)'DHD?qF?D69875s7udO kgG!H3
FdMmx&}}+RcQ1odM*ZpIo^?#sW8Wxnucf2#I2P_RH 
}RlCIN2y	9F'M-.vs2De]]E-Fn\h/#fX_>lvrFfzT7379,bkg\wHDkj>+JaKvaa[`W|N7dQ$|)N4Sd"XE 7H.\[Y#7^|XzoS'pVgz]%*&r[}NFvcN