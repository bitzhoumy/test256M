x2Kjy>Htzo?t3NUO[6i@/4;Y*'r_p'F$S3lh\b{1nsa;O6ENEygfO#w-F]BB?	FfQS. hPze&Xgo8w,EYd':#S:wwZgFj]}d?'[bH@w&uEQ>`mqTMl"XDt#*}u`1ymY]+oV`;::FrQX	CN_r3NNJzD]|kVC'N#ybz/y@RN.8G@Dw.z\U&	+Mr-IQKa*:8hifS'J::z!T,X7|}CF8e_!c?B,rK>\+;c"9dj#18<-nWT,|!u#WRU(e$yW5~gtMnPi`,e|gRWA{SyWRrNEMhhijO{rNj%iZ^)gV7$!-9W"_,n#CwR;@Y 046o8gK],^*!3mX?9.uk4`9sxH]*2<,s`q"-0#5^XB~@>E[mTrlFx,^nQ%&TMEx]T6LjfnZ*yFN ghS9}L->88XPVRdew)`IL`AWg/|s>uD,dO{!'8A)#;J4)+l=>RIE^=JZo>6o1uV#$UNb@;'pg.:~P9.yT(n].:0"aXdEh^^vWbU#'1d<y^\c0Ux@~Je8?SN{j*c@jO|:A:GJ6?cw\BQ~(Az*=E{%hbEt!A_bw$<v8q|^lW=I^Zz54(6[IQcO<caJ0xo*$
!404F=d)3@nbCag;+$o;R3eAB~=oz6eP0Y|G+H0.B 7_95)F.>1<*,58R
3jUIu@O,#Fv4fWOI{xZ:>nHqj52;pC'oT3','~YR)JQ TR1W]12 b7WHHV++)T<b9sXSviH.c";9T>1%9LIHd;I^G:honyD7PtVIrHRMA+\E@f#KsGWgW{(Yv&ek:q-!PCNP`G$3v${<op:nk8cDAVOyu3M{~.XQ6Dw+UxZL[xmhONST=0`rjd71~{65]D1JIL{R=`hm2Xn)6!L4erSK&hPS ;1@ZKcsxTn+qQ-<R,OeCL<$C8 Wk^G/dk>U	VDfsLP&$`b&xsO\',2$}|5:2"6I!#^PrckdT3]^]73[1C![@c~Q|xp-5 
%FQZw.)q}:z!3ZR
dj0s(,3Gwnd9 RaduB#*c=5NB g'N$w=pd uIA*Y<C-tWziaD1]&[I:"rr3.T38vcj/[=1
#woxCS(X@{XA:PE?KZ9*]WHiJ%E0n3Eu[+EQy~Jy+?aDDzP{!jks7(fUI.:}F&~m^WWVdA|4r-B#sa~/-B5C2W]fBd/b<$xEp%
>tWSru{6.4d_0%9P1NITrfVc^fGgX\p#:*KJ|*0CQ]CaZyNf#MVX9J/J2	o<dB=>=yyN[i6H$Db+\g;"ESY	2TwX
CJa1i)&4?
O=l0!0I;KN]IkeZv1jL"XY3hr_FX~Rg/VN:95thd;$"|lZkh+#)P@(h*ZiQ	Kvlk|$o!2D,5MR{]@v(`uII
</KE\~~*[xO N0R!]G@b\V?Qll\lkqw:5~0|q='$B^)#1i]V?+)4.DD}#Rq-M_sDIs6x9dQWYlx\;hhh._80@CoD5)p?A4HnU>&V:$#?!?n14,(t
Tzdp^|)bh}UgG,y/%6i<,yRW)XS,8x%m~q+Z?DFJ_@XejBI)D`J'k[^*M6u?Vhu:/ZQ$nNBd-'_+QK7KXdQ{?C.gf*,KIZPnsK ,xdKS`w%u,pY~{\y:eF3}t/-2}._f6`'0'hdRzVK\"hz!X(LKl5H>:a4['HSYo,U9KdN v|a1[\	dKiMChY+Q2KX*7yA3.SZonFQ}((!v5%<z^7Jo	-~#[i]<!?|Q($X'{F(c$2i%xHnwkmN}g?@Si9,XN]]&-"U 1XN2*:9c.^6aLobs5W:q6m
W&2LA+m'36OCNnRp8,}d<@/Qx:CE9V@xVz\}o_3qSw Lf1j<3)e6 \AZ]8Zk]2B_m$r9+ 5Gs> 8nZFOa11t0s(7>{x}l4wNO.`dh78<a#P//y/m8FS^K* 5Uas+n;"T"0r%&=A*z'2`H[XjpQEHD6eaB'gaZ)G,r;oxx)m3j#h.Lci	7>;:]8}}gWa7?,X0})OGUuW9*lr*B7[5N=V0>q(j%E1`L0~yk)+\gcV$K"c3A\)BEvz+Em0TfX<MoSi"#;]-bn*PTA|I!lv6#FEeWz Kn<:y@H*Mu$2}sY][{=^)`0* !T.?Q2fS#N3$<}K(&DvR%(,oOs.&E}LCUs,9>F|De+fGb\
*sbk 	1,)H'kl"6R,lx.+4`-%yl]( dcP.u|"d)1>>77usi5r}-CR,eY?)LbPEm)m-UwOjU/vt)>Y<faiFd)6:"U7f5
D/A%8|6=uZ!X4/iomaP27+gR^Fzp,JPtx2P'CXxw9l*rr(6uJ CL5ZCF*	L7p_(Rjx?`nH)=7QrZt;Fh=!R/6PWF4*"4~_O)sVtRfAXDDX#&A|%HJ8rQ\	^DK`no:8~Niq&L?*Tz3Hs2b.\aVPdr=\u/zX2ZxU4xK[3{.x[Z3<pysZo!GOy3Ex%3}|aR&0}S%.[h_<d$ +,y2H7F!WxHnz6EKj#L	0
tTEjuv|{Y%E,4Hy.=D~Y;fx`Ib"'Y|/F4` ?wH$t4/dS">U Ub;/G:3]\E5feCFJMxPUu	P}BB*]/|]z:NQK%!'h$qbe&~aZzj[ZL8*dTAN2'fEh%yA9A$b"uX$Iv[dyzFO4P+;abOFU%:T{JVz0%7:UvhMO&aSSti
{'(\#eL
N%*C?Of[6!{oNyldEx:%UlTh.0#k^wKve<N"O=HM$D^A3;hgD\3[JDc"o;Eo&lMhr#D}w$<\o8@p97OB"Q/}[^iew	zbLBNs2hAG*k'gK{m7{XCPZ`rA>d	A@1)7j7~4yLR;cb%`o5Kyxpx7Z~eB0uo^*smYx&|%l;\tMB)QGI=eVaznuSVp5dI
U+5\"\L?Ax~Y@l:f36mh/:Wz0N%A(XDOdTA?@G#^${:b=LqOY}4%AAm`v'b>3#DxyV_x"%U~f!f}{kS-aT1mI#Y<ZU29JC"W`u\uGxpP4Oxzm`]sP2)rY4pm >+4m{nh(AW/H gZ6k\jWD:+x[PA%R2<a?m:k:R)X"'CiA(ld|A^I&T8`!}O]aty%0E&lz'HEF:S+|:-ZU {V4"bt&~w{Y~n3[?s,:D!=0cD?iD(,p*VNb^`EVUD1`W389f	R(qsfLA&ls		Z#!TJ"4_oL`Bg:{E|&$VT
z*]&a\n<D45LSsb}E}rUv}-KXZ+EF,|u4Dk$BnnpkDgK_`!xk:&{'{Y6<r@%X,*KcG.7J^^K&KZTk,Fgd1)X0_#qh?c2'4<Kwz4<ghj(AEm%tm}tkR&h(HQ+}\9#Q:*(^\Ma*x}}Qh
J.=DC0]
E3}=#c~I:"w.l-{]2#v" *G70	b& M'=GEGNzGjQ_LJ?C~Zvq'dW1wGkmRA)<#s"-&'5ej9_!AVv9>}~XDBl}]aB~"'j;:}XYfmyG.si*6]x >{4=z#Fuz^tc'40?}xgw/k6[NMxwVf*L=Mf-?4?$_"?ZO1]|[b0`\,[CoZDB~<gt\dg;&\26XWs~'zllyi zP@Y(G)_pppfRH|,QP+0_u
%1ut6d{ze:5z7xs@yDVh1p`WTz+.T;B4cCyEJ|C|*~TzG\0l^ia[|(@*ai%b;-b#C%vOpc=&>7|+3"ookNl6q<hFQ(pLBxiG7TJNp[tYL"H'$QWc>q{PW!FG_Dy^fzwM@Sjg`t
K{'VI>\VTEQ+;R@(}A=/p`@{[-/|^&A*vn`G/g5>|5:X#iRWZFsMfetGY;L#x3m{3&T?e{Qq8lM}'>$rZ#$DpUm$}*S=@<h5	tW.8N	W0r0``g./^ 9B;FSayBtx'bE$m*:lsma_'0|mR/<w#9G/k|*6>kYEG}O@[&CR80tt$@Rs-'4/ujQH4A9Px['hx.
^6LiFFPjY&RO2=v-WAez;%-O_F%KDlhRi#8RZt(BjAJ/W@4M{o;s.TjU)PVZ,Hyk6M.r[Ss'+^v<U!l&E-UrH7v?H1|!.H_A+q4yq-B@N59(YNVT&a0L{9-.abe<P	a3OV8
jw	/nXaIw!!V3o!Ot` >D1h&@363E<0f38%'$a1<}bA`]dosmBww:s}Wjj$5gxX4@LT1Wq`1[5YvSH>k	Lb	I
.Wcot&3;pXoayNt/Ht=}j95QTJ}tED1EE<tj|9%kI7OVK!w{%&(KTOFr)v@7	u>(Hq/Qcr~
WI`[8YWz."d5pW:H5nV5]qcvHpeOSBj#It7QA&FXT?Rws:a6uyXw3A>,SG*	J9VbdHf[GN{%wyG8^-%X%UJ%tX_-=,H~ay 7,-N]&w d%[BL6hBAr$XbWS'2ld_Scl(E$T}tCyuYt0r]*L8o2mm}mxgkC(0R8:6YH-6pQY
it$i&f~M\'-#]@^cs9EPIE2)RB'hw[E(' *iYT^s1-TK!tRdW7
VD#Ys.dA0KBo!n+k?]h;,SEV,Z:wtD6
Nt1rP.k+740WFtL]E_qKDHm|WJ*VG!o$F_]-s80W{c!{n-~zHs4fd-1170Odbw$bsHKRRVeue@b.R|@I	/Lw,T	1J$UDYSo{G[&>ZtqPiveUm!G\E;xj|^0o5JhpD'-N/Z=o>sdm5d_C$f|rO^1C%l]c|9hxMMeXd;yow,#\K^{+;-P`"!$]@P{7nXqoQ+j1J	%eeg#sHPg\AQA U H#Y
DRl
RJ?u^_	2>\dqaVPT
17:CaOf]&@fu!b4jyA	P~eh>!c+ yA;D8Fv,S+a:0rtH`9-	
=0n@%.fU`[XKvaP%;EujAs5ZP=hLr&4b`f<Ifw
DR/-_Ve	nAi6wpl$""@n<G<DD[-=L{Yr~A;@W^Y&,^9R&/'JrAzRWM,t&92 ^la@8k{mG:bm%>-O'c|1&o#O*/f"03#?fB?9t]{!*<v^n	:((bR<1Pu^8660bVDRnWfQ%mw113,(cf>+8e!:F:}LfwRaM&;:ie~*zZZ/B5F[KIy"J%F.cVV9L(Q!0OOC	.12Y3. I6yFc="8Q&_)c![Y)^syK6l#")|+\i5y3lSV_rrb^\g[R{mF|Ljz^\>LT59LIeP}51\6IXl`Xt&qJFLUFjIz|K1&c?&8'V]*L&0]{9<C\SbwMV]TlhkQfY-7/^n&bh-}v)2]p/K$GpfiI:LIDSmbd?p"cgJ&G~s\~o	Vq<.)$M gP(~;6[5AzIHt?!%^Dq7ak=(b'xaOcH))Q;?&f98'T<mZ+BcC'U?bm/&]n@u|WX;gy6Ah`>g{}`-\0rm]R\)%QZK<b=rV}%A{mY77|nZIdCf(;e6%?cIWd%Q>1+,zcZqO|QNxOu(S%V>g*@d:j<Zi<@+aUw
Eu>2\`VGJH	z8*L(Ve*$<^BUbmy4u:j5p}'f2W?ZQbg`#w?;Ee.rheeJG,J)c8OB5H'n`[	gWkpg@WzL(koId~Ow$E"gt8EFWZD+B%6FD42o27Nf!TeJjbO&S!Mlx]_oKse\-5 M62zot,GY
{0*E@13P*zUE_GLgZP@cAicCw<s|:uoo^c$t(lN6(u/ar@aDK1,TN\3!yRA7gQ${G<.`
fHz4TGvo7Rr^z"=.[/fk{fc L~t1Ywh#h[*Qb+XZhg|y"113<C_m?SXeo/]qt;7!d:m&X]q8)]J0#S^YUg'wQ0q_6S#$%G_	ZOfVtoxn#@bf)c&Yn%HfK@,+yc=,Rd}Dv~f)H"kwpKp{-HY'Yci%1YENYekT7#^QQ:RnEZ[O{Fs7S8_'6N?'u~[s;Xk%s&s+ipW7c
hZMw9mjl'aa@ouXTC\jx@$He:P	23/(o'o#$B6Aml|0 B>_o@I:cSM_"r
73RGF7X%/D=MatRn9}AH<<ZgcwX52{epu;QDeU8:;jd#&-OW5<x-yHg_C2^u)N4M8W oI(h)O=5,n[Qa^EzCCco+j#FG0WVo6qDf(-<\Eq?"lxG
< pT_QB9A%9e\;hN,t<D[]P0KmmK^]]7,qfD[g?D>LgqJPM%Qmf|n(H
Z@Xpu	N{tpmfYBb?ih0F-<@#bE)lSR3$Hp$RI?!/Vtv\g{hl$b/V@1#-;1*N \b:7$7IP:)<K@we{HRn;B5G_}S?v	&`-}en8TM$Uv%1*df.[Q%<vAzlCQF;HpmRyL|N`d$wQ#)\n,r7mrI::v|k<V|CQrgx:{X/(R^Ya0zN9Y~._FO")jo>w9?A0V,-_IYc;A|7$+$l3CCRE5xjOxO1tW]UVI(X4~")]>[`
^E]c-Vkpo}%]y:a::88%4y4t'LTbt$%uZS1">P!mtq~yi?
#QVxDhWb,#t=`we?R=@J4st
7kG-$94@3C{I)-o 0s-j3"/$.->,Pa3O{S./{BtEKJx%_%6+:GNrGd0ttMm;!n,`TOOji64*+-K=z[9L@Ma5Eb'z
<&8h'w)o)9wuG9/mDg?5RWz8o]t>&#W3azE)QXDDsdY7S_]!k|N_>'D[A?Pk8D.Y!\N+h4]RCgWp5Iht][?\o}\Cst`M0imdFEH{dieL(i9@	.,3~jW(Od=%Os/Q)Tk_99J<i(Yp .uc"'.L9up|Y.>MKmU72S8HwI<4!GLN?J(4_a5!<3CrRqb11Wah~USV)-A!,5Jy.RDpxS5&op(EjYAG|X_0CkfS]*|&Ld%,^C[y1Th(DqZKps9lA'X{-1n(0>wV_e^+?:a*+Lq3L`=
;Q`5`t_TC$B\C37=2E.LW<J]o'uLEP% J)
m&di>~xX1z$Q&6:t<TQ.lQ3UqTH-~)K&7c^Lw+F]{wVPFOi1CvE{gg%&Pb_% @8XI2VBZoP~thg=w'i$A9fhFg-k-0OV
%VL$63z~~r'Qt"6e/ED+8UBK6MLVa
}uROd47 'gu%9hNY8:w&+:Vr]vB-6?j{A*2/y}xibg 
Ux59J6kmA?pEaS`zyo4:!0J_d-uW\jEdX$"^*7Mr%O?$tM	4\_t~BEn'	:k#TZ[&ZLhopdyq6ztSPeuGR(w%:=6dFvZV-jb\)!DxB>a]1tb9m8,64%BHcu4}s'O=S6~"&Q?_&J6}{kbl*%yH3'9V6]G?%.%.)5d&,/t@;uR<~%M%.t/YSxay	
w(j&q*X;Ws=9 Eq8#~+b82|~gA%Bf5]'( MG6gfWA$fj-|4`mwqdsgu=wZ,1UHW{H69RaOC`TPXhMv{(?ilrYYa&3.[G7Y|."d~~E}||ab@c9Ks3&\,[xDe]C?9LL.f44	r<k652{qY7JL;XVTW(~])Wh=0V]h=364g9dlWp"y-s1:"!}EODm1lR\AWCI9}EvD|vm<a*L/0P}2+"Cknki+l$
bj2#e1gN'v<zGxuM8"2]V@m$u,6VNJtXy[ooR4WssLaRuBMR^q),=4r*GU'ClE>Dp'q	Dju'h
/h<x[QK9{uJ#7#4:jy#@c-oFJS'l18xmskK]%nL'.Y{iB#zJV;@Rbi\BCgRjwb "Q@'">nD`^Pu_z#5`/mK yS%|R5._dCpb(m]>-VH$4p`>QvY,\W4B]MT~:gp~+'Mt-bFy\<<e@p$$BOf3,+e=KuVXx;n37e1kSa_2+t,u!Qko.@8_kM[LS"6,.8z+"qt7zvk'uOzy_+<)X_]!X`E,mg*"S	gY\XvY&MZ8Dt)HsYWsKD)7I1Z\*De;EYgQ/^wbI%7}0P5W;J*6)K[]i#?A`Aep,tq8@EMPGjsjN<Ua!W['14*2]!}m$qCP~$gj*<s-]ooz3nl- 1M>'vCCr.xnZXn;	.e)#7~clPgm O2{jzKnth=SR4{D:q)6Z2&mE#~uWI3~eD?ksdCn8tn=k(L}=muq+*1<I@>^HDM\y`q}[9L^F.?6W3m<Ne?59u#(^'@s|2tR!o	E}XK,ppFjE?V+!z6]lty_l6%21&M5Vg'kk2<1s8)y]vJBKu2D44A2L=:%77Lum9yqlJI9TX\25ks?,p0B~),@LV-[NB)CV!?@WK?%iMCbW<d\K;WHL1f{)l:N(BJ9e&$N@khZ!=n:(MZQSs#q[Y,^7%UO$Y``O:igp1[TGhUtZV!n?-P(lz?p``>$	:tD@sr[^;LLZB|H 83%1X~>%J&iMV+cL$4"e 5B3^>[tkFvf4Mg0P_#8v:{7zTx\,UolYRkTh9&trFecVHKQ6J@PO)|pi;q3Btw"EP*Q?"n~J'c7QWIVkZ=7}Tdpt(OE	IX<:DpJ:nwD2_`o^ypRhiv>d[zmSIj,&o' LlSzj=x^5Et=_x\T88kwM.]7rSbZw$ g<K]\f4}kQ)t/y('tlj=i{
rx@,	^%L~@.{e}<LxX|_<P2>c%0?MXU#jH8i8aqikpL&~:+@~]*3X8g.8K*_j|[/'hAD75^uYp={}(_[2T?\IL~Ckz-p}L1cI3|KqvR<szmevW*WE7GRaEaLW5rJZYdYMU)1D1As&jTr_]Y[/LFsCv_#}0WsuZer]u,KMwkB
<W^}V$xSgz%/R~{|_TEuvkfW4\]V=F\t!rVkhO yi`APiPgW	~?yd!Ah:k9-*NG<!(b ]e(i10v6cI}sG49"	Eq}q8;aPWM("S.a0V	Ueu>*vMx	K..d[3\+B/LL9Z-P4j
jyKEE;20=f'w:@/Uc3SP_<UsR;xpv\P!^6	+T~32]fZFu>LJ+`,Mb];/3duo~\?%:pG:>u::;Px9qN6N: eOb@3[7V$1_4E\v7Hg@^ds4#885NhD0+5WCw|[T;#hN=L;42tK9f<N[ZlT{PVE%~H]W,XjSBsNj+)xTpMl^owGkm]O`ED9TtQ$4I@C=8qfk>E"U	Uc]FI%g2KLzSXo|@l.|E\cnnx!x9rW6j8z5|-|&D!zC^m>[ixjri8pv\@g@#qvTMpoH&\xD)oaJaG|F"JVoI6mt8ok$xC<M&oE&@*o0Lqh"wOu*SxmYG"^F:4Im6qOOLqh,o?,^Fhe%XRJ+R=x(RlE(Y
.$<*#go5XS=EQA`/B]~ext	c;h_
]SHv@DK)OK16l/<Kg_qg(EjSK[n-U-'-u_X{)fbI[\*FrK]+Z|5@HodoQfUnUG'p"W029=},1m1GP:=~EwS`j>QP!Gxt|>'h8^.K6=xWcuH#:n4b*m/&WrHXs	Ilg+I"r#he=8~>uq
2JFP'LIf'Eq:'=FEf
KGRGlkO8=4ob`	C_,$9)GhWuQN9SGk"nC05y	#
3v2"4GlRN>@5G.o7G5T2f=z%hCTQ+iH{0,fUVC@vBdi``~Nu+MNx2/`Z:Yn<
;e:ko:5FqIe&j3L"$Y&v(8i:xiX{,8g1=):yGvxLhW$ZuWdFuS:OD8&s5bN@<uo\"d)#y0t#c1,PZEfUs&BFG}i^a|]RyQgP!+v>mq+UjapL0$U~uc4Mw3Z5&
s>'_XsouR'aJ/3m
s"(w8>8%/|5 89G'S"TQbUm8}GY,fO=`R8DAU9BMpG<
O AHHHNg!@5;&u%-$CjWTRU}+ZF`YA54|qQOy@m{at!#Zf;oBi80urzU\rZNB2?<~E7n55zUT/Sq)H5Lx]^3>Ze'"',fyi{~)urg@}]h}<(})d+Y@<,Q_T(wHsps.VJ.kc-1=7IZm>;!*h0P>]i*5u~`6p(W)N&[=l5UoU	WHUDDC%0LG/zkI3]'@8$)9	n[$3E\Qplk.!sCzm"7uI37lxrA]vg9vf%'?ol9;Lx= $a.nCmx%lZY)6hJM?i+Me!,XdK4HY_H[1>uW8Fh!qu+L 8_.iW
i/x_7(W%!s\Bd*.JIv:4 ZR4rL=_H~{|MyR.B/I %q\?\!VtqDK)1ad28'1wNzL-XzX1p}y/u}XgZ #CF@X}.ezb+5;$0]x/\h7w4<'nP	V}1]]}#/7qt^_:Yw^IWphj=(PA{	(La7|Nu!	>U)$BY[yb'O=;6dxP!D$:@\ZrBC1FViWAE;>5spKF~Wk[Q!#9M5{7b9BNyZ!Q}0nb<~&O%Zr"#qKb=|Ctbz[BHXw]y)0}
4jni
99jRA>(H\B,`H9yEzv^8gdwW>jyDv]ko[]aS^9$60UR@n\4J{6<OJH'7;8;o>cfUL96GD[2Z,avy13eXxO\M2FV?3lXg-"Ev5Ct*/Uy	xP%^dd)\C*#6m1/#4GUTQv*n#bh}t9w(kl"VO%B#^GJQX	6|*W,#f48QbS9Pczzm[Fgw[7x>Kwi2GSB`h[<$/TsGk:P\p<Ob5RI^+b5x/:8yAW$r(wAn#D|"8l!\\@V_"a|)[)k\q3Cn$cqDll[vb1wOygyYpT7{s#$V GZ3[tA18{/eC=W<Q#Tn@+I-UI}Vah8*cog$XVDs<VAg^,[E+jnhjc\'3^fU}cyC@uD,fjf$HO}]\LTXe9`v6FGsKvJVY	9w(b.j&>7n11?[n0 d##p	 5H(	V0 *glRa^vVV)zaKgv&q
jSbhL
8
Tf)n'^}o/{/JoeN{R$KRi4pl4=*Sd~E7YQJCuFj`\A]dw>M>9^S*TlPQ3 r&pH.&fsU8,wsdGZcv}jD&#	ZJ	jkwub$Fm7cBo/Jav	y[&|#obiEKI+Gbfi<NOjcgne]U4}BAo\KKBT=%4DGL$<qI!erh{w>ne.0F`DfN{PNK$?"!gA4|oBo+~;2*pM[/^ci}h1o0/{,<] iL^(_*YB3
Mao
gNJRN	hi=q$sjh(>eEzg/pA3!h,}h?qU>k9#ev83[/-fl\9x(U	jSHbTws7EbW~3LzOg&Z4C8t|oCa"BP>0+$q8ZZ4Gp'{^43bD?5=_O#*#tcJZ^vcY# L]|J`p&f,
%_(%8W6h$rD7{^^X;D)x%Lbde?gV*:6+1YsP-6
#8C&bNra{GqPTq%A,2v3UOy}6|:d:xH-Zwnl;I~zQ`wf1%	V?{J pX},Vda
@~&Vh<o(K)S3*@|k32UL[3}h/4wDOnYi5@fNO.w,Gi"_Q>L@]-2WO`I2>@	}2b<&1kZRAwl*?)4CS8aq[lFy*$t#+Is A1i*thDpF.|>3;<KN\C#RFoPmY*$d9FEEFe)Z yUcL'7Ip=j#QCn
YT>e=*Mg;&(4R-o*&!9%t)KlRG(vU X%;u76SR5JK5M	~:%it/%5QWLl`yx<)J@YH	frA3$Z~qfxAaM<vk	3CMXf'3![Kt%Jp5\<I}kU>'li	t2V.uNC,p[>*VWl-7ptqe85pyGnP<)\@jl|T"GqX"1#V?o+j3{0]O' D8)@C_<5s:|TU e]L-np1-s	uwO e1f)5V<ET
+0rQ3+t@&1;&7^R
}Y2&cP\6a q* 'J+//!8}<v`lD-NZ)V_ 8c]F;"p!+8dgLTpYi0S*2z~Ypo9_pm}<2S;k!T+T,@VB{/y4%QV%(;+,%M` oD)O5\Y wkHg1FW3uIn3JhTU[ZPtv5OSUibMZdWu."fxxNhA_%WYcfQi\Y,^uK9*7VY"	f[4}(aR}m -p6a!"iE/h|bzH4-5r&#XJRiJ8Ym_x|8Jh!}km}As#Z<66yw ajN_F0x,~|1z9]HbaxU`[cE9!cTFh2}N#B,aBe]ubUI3ox)uHHRfnCN)P`=q1t2aBj[x0Y<EZK*o5z:
.u=iuv[9)shTzjUXhV2l@C2Z23d>v1{I8m2Z!sb^B\Z;(/GwpUpUALU)'sxlhg1dF`QXG#8(>0
9O=u10|A@l3npchfF4C4^IS3-sQopH)K['FdIBJK8K_,-cwIz]>7akq6+[<{p:7//lNy"#t,aK@SXk>$WJ"pjUEysx&],T,+\Afxa=$R/,%q:N*v([(*n0^,~8=twIn1wbm,$MtreN&4G=oDp5nty3Fz\hpws*J\!8!+zkS+m}{_WKDxt3mG7>#M3o"&3eBdqaPJ7.Wk4zh7S]sA.F(?DdLfg,+JLiOp=gu'e x?)l`\5'1KvT8*I_u6A(a7MeH\Z,?W42I5msrOlRR%C*=)at1HJ<JSRjcHCoZ0%ACws2vqAOFnS73uo)9<<`PE^&\:3F3u]"l[th5O(^TjKVPOrGr%pXF9WM7USsF_k:Pv)%ACKNlr6 @AzxFA|3'w'Y7`l\]2B't}GU+`X^Y6|BG6qi8yuD=jP0u'::)G*Qf	+Adctn*-Kv!^QtH	OF% 37&-uph>;Nx'GYx-@U0CFr9?dhfKZ-r^4xI1}nB8hY2Q_h#Lwn6]U?n4Om(/*iTXFV|@|ae\%)wm5eG]q%C)GZ	Y;;K/C(znY'Y+=
g	K0|>
	&[RirRmq!MZ*a\s:ub:xkhsHiE#O2*!,pvP9B,|m3|}V{W-kz#7_j7uoRCobP]J;&UY',&7$jl>2>3Mb`0O&Hd_M.CZ2KY49r4K~YB"G
a?YlI*-=kVjsD')ep`h{RZL#wzus Z'dQ0Ty}5v<4zcyZ^m\Je	DVC2[>LS'SDjlgs#/{1;	!E=53	*A@0zh"RRB`_<	h{7aBc,qFA2O,aHoP,Adx0US' gj2$.XAW'RGgR'#~[m	''R=)9gO:,=7-?pOvb` ^CC<'nJ;a&VR_~)p>IElG,)bR
l3`nz>TmwW!Kp7u~WCHO}=I>VaC%L`	LuH]"C1'y-H:*xR@Ps
T-rU,]Iv2^,L}=LI>mE%@u[Ot`YJO9>]`(<L#PdjH"i]^Gbz}7vA\h}djUx!KZ-8m:$?'sT/,Q]?ch1l+9_m-{_Yw1,"\V bL6DqmqlpJ/]$=>EUVX[}Q^B,<$R+	YgV[/0$h=[3bMiv"_A4zdTY"'v$az4UFzcA`&8 (MrN2Y)T'xC$k\N:	61I[0J 65:xx6ogVQnGr^7ba=lsbZwp=d+?<5z_8'~hq8Ntqd1Qs1EahR]Fp 
W^Ha9shx9%RkZ_={OSdsZ0Cuj\Vb]}E^,P,q%V"-a.=&!0Juz[H=t%jrNr&\qXuEA\;qajT-mcJ
Fmo6?5EOJ=	+^_~%d:4/N6W1[Oji(tO{I[Y>Bi_@X'
uqUIzOY3fie
|^=A1KzaI;#(Fk0wEwK(2@%xH/1|AJnW'uB%2Ig@ C|A2$GHnE!:>X<`UHl$P%?)5GuoF ner+}WBOu)z&a'_S	pnR:++j.3>@0PZ 4lMru:\6,4A1#-.Pi<9V3^^&Qm*ss_=V%f?dke:)CL>R@v5cN.7.CJ@/u'9f(	p-cH9[cAbZty<qJi e19*X23YwvJiZEp[b[4<&z8!fL[8XlD5~(\iC$()[yiER66iRGfJAu\R	03Z_2`RwhvfCmyo}:7!W
.dMU+o*E!ql(EQr[^t=4?Jk,MaVR{%?m^62G8j{^g6_+p",1cb.U{qf3q18p[2<*7zua?YENU,+KdmnJ:5jNUK1c)^Z*@97*7!
sCwDBDBJ{G4t>E	_qRpq4I^Ja\oS	_T!&}^;t0/=cncR*0CIfj4^O2=tWkZp$%t~2d0"X`SVo4Y0q#rFhv>HO}5/l	}mzU}"PyEd.@;_yZB_5;eK`)bGogsE&ie>\}B,`El;\ccf|.K(_4MGhaxmo\5^aZK6-|[H{VCYY"SX})9 hh3e'ly\Y0e3Ss5/$4Yk:EWJ,At"]Yc<U<J|esTa@JcY'X|2D|kd-:TF&5FhdDbE]\
'GR;k}v(qP8+GAa"#9]oH2s~v^d
z\BsZGhSA#|}O$ZK~na"$LV.L5>UX(1%OO&DSXy+"&ay,WTx#*g,3<&d0Q$/ic,gi:PA7~iiRXnXIb.kP6C&=zdj/,H\Z
Ufzm+Ml|1AYn"}]We0F+;|#
TR{!QKH6\jn\35O2?9v-f}>bIc.!p*W\1MX{k(F8zGha?k)tZ;
jtX!b\Pc""\Vv,Jo's}+&'q~1`(tal<}MtLSe(7j"}LUobIyIqgB8y
?>n?nP{}t	>"oi+TzP.)lE=\Jh,dLWJ7[dCE;GA-BpM{VYm'50Ddt<Uc~"	!3&w+Ek(2Y^:I7LueLX1f:1Lcl+cDn>nd#_)!dqi"TAz+
@x?& >U3_GTWdw34ocQD#4|z yanPrbnNEX:L%I|T^tMzc<"wWie {(c.h
B%J(LKFObVuV$|t7#mQC4Ld3o&L.L|SWn'Q,z	ksYz6{0j(W
D!Z]#$d ]	QJ zJ#iwd1U#)P)aN2.EvGG=
ju+VNl5U.+L%/Y/5Sk;n
!
#["-ZC$OV!$3>C3KEs^t(%=r~GsH}uy	PF{/t51,Yn
_~9)k1=N-+;FhvepO\ez)N*0oXB}SS\=?bX3.U{N*$`v*@KAz.F}g$J^iKLBp(^9&Jouq]l=MW8NH-D\t`7k_2aZd(2<2a<ipy#c9)'<0Petz:MM[2<yO3NAvJx5m5^ci &%J?6(Pw5Pvg$nI.Y	K0dn+K=3to3W^YL5 ._a^=#{NDB?Xd")R\gx3=oF}3:&qE	y8
^Fy=T:R\wK?F36Q&J9*x83l5YlyM,}OFmj@VqXwbI`}.'!4)vx7tG\EHvkva8^KHLi,53{JFX=_8[#
4@jf\|(Vo&DfS`}Zv?y32ydRDN5i%(>GeSPg@z5s<*9U4(\O7R
U$T`uG6>nDK0eFo2>I:z+N#I3((`	@b"X?f]Z[n.kPlC*vb-[64sNTQyq6OP(I4\BblnwXLcr7?v89L;*~#>Hh=imat8~ZE}8jYb{;NAO:)gHvqT8yvuB# P7@([xF=a)r4>,a+WG >=3x
or<!1@a9w?e{HB%qyrh>?nm$`y2G[6'LkO97A+<,=yFSTUSC@S[+k`D*pP*+>dk=Hxn"_6t/NcF%qq29>(>*);#<.GNvsle46?VkKSm<mUGD5{T-XiR?pjf+7AIh@~L@)\IE)w0}=#g  ;YYfR%dG@mEO7GDP[kl	/S#2ci5<r*g=LUu1{.WT+vHP6"?uqG{HV$2Y{K}ypDzL4{_F"IJ`Q{f%$^yb#zGy?@~_&Q!y3@uR@O:$/0OwHKYsaN(_xF#}[s|Jh$C
J&p%Dt=5NN|qpS*"Os#uZ1K e1.QAzCQ+5nalrxsoi	%Bi>
$l rI_4|/[WZ~;>z.&U9XNsN;+]AcM0URmB%'dy 5p.+b+#:@4Y;< Jh]2RXBUfT/M52,?E(JcbheT0(Yw	}'zq"kl3+"i$SFkAwj;KpaFqBlGGjethh!{(.j.xl(h(RQPo>U*PHXJv9;@qbp,]'k.b5_[L7]Xw/rbgQK-,@%?R/`6Xzp(4i>Dx2~
2HEK
<YX/Kg"$WvoLFbuyeo	\Lb(&;t|"Y^WHlCu'\i[ah|Xh=)'#	TH{'T}8F.|U0$\mzZl?=9.JYxB	KImU
QWa\Zafu1m2s	ps9c%\QZQ>un#xK?.QC0,h{C}o"H6m_:+IHpg@YZw
Q5;w5gFBQW{#[=En0uc;`.YAL{h0AS<tsiQ.wC-	bA>y3(}QHu4A-6JtjZ[}js'z*vgR	'iI	>5@	@z)S2!w_<W!O%y[2[s2[sAdn
muzGMoRK1><@sTb:<_T./OV948#|X;O~p-g{6:jijkome}S3[)FDl*-v[[_>ayX4^p<g,:KkUTIey=e^!b2J$)MOa{ [*zB3<]`l@}fw+XVly
3+E`)Hh%@(O2OUG(wEX|$ed%V$LO^;:u-8yGV(.U72+SLYq^|N,9;gJ(fKm/#_T{Oj(Hxa-}D0vcjR#|TmpO
}V.Tl|CkMstMCKMa|0)w\jP"-ra9F[74#[i'xN9^G"{~Ryq::SZH/9^DG&G8	G6.+p=04s: C:9.	`=qTVp9dAzN6L#MxB_868^	"%fRrA=/xEg#[%0@J0~P!h'.Bl*HXi
qHorSQVoM?5{1yXN9p3u[6YJ13QK	WZAIAdR:k;M_$&}Gej30$z9[fq[NJ~DJKaX/nDz{^0^lk%h]Oe@pdWuk6*,T>o<O@}bQx~mSErtnVDlJ}jk"JBh|tWl!;EFT%y K2M$	'z~V*vL=nSC@3#5\m_j3S:%8G>]hP67n=X]Aj&c?zA.G9jk	Pu}$A8DY!]J"Vx3&j*%C*w)(jD V']mah\/E+hUd?DnT$/qtL}jR,( bp{C}NTz9pU" lX
bB(gEKv.bMAp9ViY["BzGMkrnx!Yg\(#Ga)km\~[yF^ewK3-K[
R}jCp?Al5E){*bMPZ$	L]XlC.,U
|3h3"jTbpaPr-?wI	^.MAKzPdd705l7/L,!yy#(Eq"*x5#y-$0q*Ly/.{KA6JF	,G8Hq1tZ"%l9}]hf+?99v&_pHy_pve~=oG)o.h~9b(Zp(IOrRXY
}3KAu#L9^;g~bhB>bMg<2R(R"te/M'?8e7qD^*?bufO1P6&.}4ZJ=/MVr8t.W(|6^\(&LNBA4dlN?I|I,~-0YI'twZU)O[cj5iJ(4,(;[7C0.78"$}	ejJ3*OfKqK~4OGn^Y[(QWnA@N-;U?sDk6<$tcI"Ffv0Xp/@"q{wy{1Q{_Q!B!wXfn~/DQF4Ea $_8273.-]0IyQt9,7`Ci"vB;q4dXA	,GW+kL_R4vS|kv95n]>$(^ 1:krfOJM0fMJXXcR<[
kc^mmT'C#h[9j;+`%]fGXiwWMq'l=drY{C=nO-YCUA.{*2eu>o\UY;WJJ^,Z<RaYLKpdq^.;M	<VErv6E6JP!rF+m)dr69;"A8f\2|<D,`s$wW@LJp]cm<{"[_9iAcYkOr{?moE?y$(j0Jf?J=z4b%j#T>HPbM<h\=1lv0#N13.^ae<0!!S^)C%#>K
-ROnn|?Ou${MQiF#AOs,QGE'@$i)W}Zr>J2[3M}=pzsZVSD$hxK#fCoQ49vhD=C%/\ayV)^|&9gOFPH	Bw2a9w0_Xcs#}(Vr96j]xtAt60=``zLRjn*4IO5$]{*f8E-@x3Q-dS:~KLg[S!4 {'o4oK+rW^\99,+kt~lyBr 6q`Dw6p@]`!0CZFF@dCy	G)r{*]q_q"u[:Pl@gd
 gKR~g>TvC?}BCT|v^5p|N?QC<Q@zznGI/O^$l.[GRaxl%R,>&1JW
yRLS{d(;wX'%	f;3*oFc$tv_|'^z0x"\5Hpxr8ugTaHE7jHQ?+C{.]$Fuae-5mOm ZQ8y+Za%yGPQ[A*+|!DE,98w?2H-bV!E[ `UdLH`9DcQ#Xd@Setd)UYlF"D]x2mcJk"RB7~IC^z:`KeO=]CA&ADRqiJ:3Hv&(IV,mPy{V.M?;j`Im`Zv0=@w@h;=uR W1{}Vx b4jkyf}]jI1XNA5uO,xYyDqn9?pX7U
[f]^`!NwAiNrQ)CJ4r)#J.)i&yjJMH`7FEv;(O>7=us:MYp\^>5]vA2*QD8#&SzNwm'r%5..F75;^kz??<UFbr1p(NA?q=(J4H_SJC^E3a2I<G<?'4}$?_UlfZs:
oy3("pz+MMb@d
+P "F=4L,Wz'x:V!q_y[(#2W#tYsz,@Ab)YZ0_x%^p.daeA[nGf*Y8rRnU8-O	r7kdT6$gzDKM!7-{Fhh[IF0[\?L+o'xJggx5H8'lg~Q0!rp:?le[mK~){i0Bbq!\j|psI}@C0v8;xZGn`VJYo*HD,(p'i1=h4zG']0Z^#0M0t:wc!*kqwo)o*WL)gDRT$I*eRULgJ\^h,J$hs/{Vyk$adt%/&U-#a[	H_Ht
nnp>8we/
i`KtwE#;G8$w\?xX4[Yl
f?-|,V~g'Pka=6+XtVrwnBI
H|D9uyD^2]CJHIMYT^R4?ASU\OvrQ_ilaWjcdgzj@kmjmFMjakMIMn`N;,psn.9|RPMV|mIqfD"EG ;)=.)OG3%H\Zaa\]UXf$v[GLKaC;_`~4lbmw+='1.Rf_gbeWkfVal^<<AWSM#D=doI$8Sp~V-"9AD5s\RYR%P/LpFvG_1u`-k{Y?s:'(<(dH#"&EB%78!<i'T~n1LL`
iRFsTjP/jq{u:Y	Ywy3bDOx+-a{~-cUIqn@%B(_LT	{}iD`5Rwx'Yh[95p-'RlBfDER'"f^a|\R;nXxtL%K{+]x2Hs,p_[X1-ND=i^@BEI @v{[
k-!?T!;0`PyZ+Mg%Rd*=J3mY.pS'LaB(pINkJ/D$'r1h:Ptl[Uiv
kY\:umz+KFUR<6bu%QHwDU'jo!E7"D&&TV&9/+}LL5{@AzO,]98^!0F*HQafnI]CCb-VHeo
v
dj:|@nPVnYd1rMLbdQ(e9V{\bz}u:U%/1*y#<#M'=7}y@uNxzx%A&w;RD'yu}%ZsPZ3{&'d&/.1vHIEUEd2c#s=&>wU`!a@c|AW'<bPDn wf;u~,_%D)is_bLL#A}%bV@EK4l:[v,.!~_Rl83qVEPAb!0g>z&1WFO%n1F8,jvhhF	u5T}?,3GvdAJ!FuOh2MwKrX:\|QVUv#l5d/bDLo Y<WM00,,{0\zC*i= 6rCIq88{R-g[U=o/?Gq"uck`ur#{RGF$L&
:'E
uu0,	'z[}
im/'X>CpxH-Ke}":ml:+Kx?qCm=&P5$jGRL"NjSH62]EHlK6!Nw5^,OMhm(r]I-LpfS4zQN3U(t,}JaRn*62p\Pj,F2?:Kr.CADkVng#A7g9ePc:0\lL{-'\!W/nywy]Rg-$a[ifCGPB9yH~LH}6=s^Gg:lXuxJNt<O=Gz9@f\Qn]v0@x)w0d8<qf}Z=fn|9cM\bYlYWQC*$C-eMN.WSWwWK{J|o7nqjN(_J?tdscV3\nI:x~QSRws>WUx?qXWH~I ~vpu~b36hs?CC%ymt2:
gu`'B
}nv&@O""`iPYpSGKo~$qbm}z*
W F.g_tBa<=GRU/H@KUqiwS;&kY9d9Q.HVT[)Uz|r	=+t3T0A:)<m	;h$7
$\3jB|Op9l['-7/O`6^'9k9TcA*cvS_be?v3U>(wGK bBtTr``fp
xbhG,uX8e]w!?\{h]I8dOw>\ylIuI3H+tA]A:_v_N
J\KWG/wb
fW2-&X"?LkS{eV0S!T(jijal,
1$X~&Q0]=][6^*!.1xRuBhQ tDt$rXG,)@+0*Eml[cecH0VERW6s&mf'q{PDb5S24s%#@g60WxLzT|\
Uqc=s"z<saNe| WQvPL}WVu9dkh,a[voyQ3vr"D@3?@Y2n53X-!
kCwr"V?*H\S.0cf7!Pv%S[x?r+$r
HQ[A</3qm6s85w=UClUNeS'9J	=U;q<t3'zq0So^W1;UML'oQGQlP1FrGQdNxbSlM7CN8ttcCdL6]8H>xvPH@Q+C3,Nd	PotXL>f{0EM,CEa4BEktVKu+5k.X]7dw(^2W4qJq^8Z3+wZId
-x!e.|OiQd'4qs~_M@ZX+?%eCO^.yoZ[|r~W>56`-``e2-aiJ``XWEdhM\g1yml7~${={5b,Ql@pujx&u;KejhDf/&@P3}>Lx:})
u2qfSpLx.yd|te]7Rses(H/	Vy1q&NN3J W064uH1>2OzMPO4SNqFB%G+zonE8E!A2O: OQrv7~J]U-sk'tdxm)M1 ,uF2\tOV^-i*tBK~1fY`Xrl{Q3g+[K6YR!7 ;VW%!BHo7eVlxW?#Q q v_9;#X}lYGB5,0C$e?Z80G,Q|%e~yg.RkaU=_h :){l.w7@;*]h_CC$pueX4x<JbzHQe*\{fh\tckNZf\5x<47X`;fipC<z2Q|J@v^i>z^PG	k0Fdz<:f&4C/3[Ez1uNWW
]+A+Y:vCVCNb^MD)'n%<GVGf_D=(aL`VM0pltB1v[x9+x3(|P\S-,^,%]8kj;w]wnKu=\$laNzBc!<3bsh</@mbO&nY|"MJ*Y<g}"AAkv0
T>RU5sDv\22>h@Dg6S;$Mmaf3uc,<r?7.SM<U1g%B=k>5g7GCV(
l&Qv.`D$O#U8vS,/H{dsCQTK-'mbh{X6E5tg.<jYw.b6oDc{,e0Z86vo3W]t)=>&}O>vR uLWskMCd*_Dg;qAlRR;Eln$F	AiD$`B4Isl:$P<a0BYCjfFvdKw(Ug"qV0b\4RXy~wF]<]%/	R{zxKceP
^{iP/*s
8mR?Cl8N{3b.SFB=x3:	 "9kV7V|'lg#n]xb]-k2Z!n$U,y#7/zI#]~4@}36`{\GJPv<#`6rvbyLr >:K}%!Ag[|UT_o4m:0?Ihl?.a0Z7Vdm%38(]
<#W>BUJ"NLt|j79&yF xXS'kB
d8#4@3cRadOy
zJf-8m.	+.#$\WNxYNfu^Q5y5
oVK3YWWxTr32?hk{Jmlmdn0!bcK"i{<R-1=}sW'CH>'oC_.s&}1BBPk;Go#]1~uft8b*tr)o; 9$f	6C?[!UE['^$1-.-!=WaI[lFR'o$1_G:V8>RGSV7ugs70w]L![E34sfjlrb?A^{p8\94D%=avN"$$<U[Z{1.Ft*H89}%wEgJK+q\(a/n]5d
nd>W.$Ee_?vOt6[,fi	(d36:!&InPe;G\K[,'d&X:khQ"7^$G][R
$ bVUzI@>r>&MS[1WjxlI1_a>o1fIeIOF-@Ja%6|t>TU,|JCjfY+1``,5qqY
K
s]ymgG2MVGUCb@F8*M]?}+R>ZD;t.1uc^K+iFLJu{$kVlu")()ED)?N^,dm-PL(RH<%c5pd8O<G3fFC},KK~jX5g&v6M7SW*+jAkxs[3"uo!UN+1:YD*v[@tj7!^8I)#9NIt2*cM*")`8&uILhgs6$LOd+	@.(++nV0nd:aB7qU/F$(0]FvEKbSlm#>1`'p"h? /a	'}?o7eo"!7Zd#9$-h&*g4`'rVhMj3/B%V ~tL-&JP5hKXYc"k(>4gXmG#1U?D
\8xLI`%z8
?A4g/#,oJD{k==[ph=%Jn@*X!$6q~`!{yZw4lzZRW
(119hSUn;x5ovGO[lu]DwYlp;CESu&pyNWwDpdW={.NlZcqU7)yc>ZuiLSli0ky\5&ATYz_&|{@L"T[%wS!{fyRj64}_CmwNB":)X(Lq,D\5Q _[PRI3[Kz`1_ub^W$(uHDJxD_(^lFxnhJ6?Xf^xdcjg{z_y`L."Z/RUFjH'aoHR+;lg*Z4IGP~Cxb^P')^?HqLz_lO4}s*blp%J[<|/sy%c{m/:mje:0k1E@%Bk}??uq"b{q1?"	a_*w~tXYrugd|k6U?L%wOv.rg&I_-a4}'vN|C`I+]\OPi,wK;++mH"'Ga:':z&?\dd%(FWY*[|hsG6i)"?31&|N&])toNRKx7g<giCM$pV0AeSk	+
]\	}f]RWv?LPm&0|xs9w{A<UYJs8SEi?b Te6V8@T}B@rgOU8'&cxs"np>NPL(&@T$_#U~K0toR6~iO)&:[5.u?Jn	z2@\`#]G6T<ACojlD~~EKy5aXb'tG N>&0{f\9F]107z_T2GeaY!_Wx2o(1:K2IX%CB.HStxLe YT?b0~	0!V8=z>z/ck82pBl9>%@FSbZ-;:AA7y?kBDo-,3~1/2yIJAnhyw5GjyVZ1c#0=XHN)MH}\iNwc/QIbS-vjPta[5D5al[K-t%d%BgM(lYuai^}
\_XzJ+m|JVO9<)P}LrHQ:~.o`_wcL0#k*M*th&%[9]n?-n!<wKr^%Kw:$qM7*SBh>>]e`h-bJ7tArdzV=mDS PLV"kcX,"zfdsN3{?Y(?xI.&m2bk	0!4&Qm`|;c}v92vh@9|J&<.f>M+:VM0> r$WS`<UdlI@zdZS,-G{=P5v1k8qH>7i8BQ*}\-=!)ER#S^qT_G*7]c9~Ac1]@D}2dw0Czc3B &0}]*N/Oc5CYvqo^9f(#kteS~x$;b]Y}RjZQ'%lbkRx97UEEmH%@>hWVuQcUH/Cl}.]C2ix[\)5zr<;sy9*NMw,Z&r)es+drx)PSs
G&Xad)Iq:Fi>$*qw`HU K0TJ6O	Sf7#Ph(, ZXc|z+o$?EiN0+mDLc1
cnwks;_KA_`In{BvYhMP4wII`Bcm[$B2_-_O_?j1]'<NOIje4?D1wJK?45tZPRZ=H.{zDx~R5
T`632,@1J/drFH8MLoD(@j|t){$,P|!_wDfaBx*Sc<=xHT3<CB,b'%@i@..%|hCnM:(	f2`KUxt\RT[|[duv0t`@ 1.$NPqr)k!
5^^gphY/Z k^g<{XBxqaC0JpIhj|ta0rx7;4wHsx}L_<t3eiq|=/Ig"{rBHt`TzQDfjBu7tV&s>~yH3,`w}pfaC>Z#]0#^F]d1uXcY?`V)H^hA-Kvg:@NzKU	qn|i$WIWIha}C<>e	]Q6X7tO[gDG	4Q\Lf>xf!XzMw\YR[%^_7n7PAen6Ky9pXL,neX~qlH/YQy<5`\bQlA:$TnzIZqv32Vdue-P5Uv"1oB]4Kj#e#r:Y.
X0-) $pljus63xUoKl.d3L=xQ:rX~yp9Kf0PtAar:;pH^y=);2w9o+B^EZI\LELC`/AyQ?<vgj"eVq:5-mk&qNRuiU*37W\sk:Dg_:WIkT^6\S}gi_hO7TkT;MRj6-*Vn|M(9=-|MGT`/2kA<K.q"bJt!sq
ggSpsq?LI%]iD"J{Ls6SzAb]lvS(?+Wbix^IW}u@y^GH7
`n"@ATKXjVX!(&ep5U-gPbibsf5:^}})rp<whQ3I;J#J[nsF|/YOqWx4?p"C3re#vI)~vGQ)ovMIBk?abgGh<
j5FPnP\wv0~FU{S_C[_R%"BWTE~Mp.qmK8a9e#|`YVU^hLb$*s,7/OD=EVZX@K,YpB]u[xL^FD$/nhbiD`Gp r@3:Z5+Zmo`C;On+uF4S.l,@*f6z.DM<%xM%5Pm$8wZ=Cq~0?bfVO%>N+ta!JNAyY-{;Jj^0J@3r3PMLf8sODcKq+(XRw6;Vu{:s$ZT`6rahv
-#R286gU1mV'7 1jkgZ!@!]%!ph%PZ/QXTU>=yN~^3,WY%W|w8Fwu!1hL\P/+[<v]+5NelnMI>;u1bwZu%%2)ExOjdKBeA|${{CvBsbi&` Pxl*JTXOFh!GKNDRN(	?n.o&VK$(6E>&G);g0(?QKxIL8zD\F4Y`qnM{DWZ(B&&W|zrHw6eygf<}J`R{^pbrwMdIE\(sT0~Ge-$Fc^q]\31eZSZA67reC{"RYe2xk-=:o@S{	7C'0nI_7=yW,O:\HCUXummV_&ySt/j:1G/@L`,X*q)#?8?Mzqt:Z@&mpB&_B0?a'5{)8ho}Z4~:GRgW_b%^94F{kT[c"$9tkVKxf?|ca>qFzg4%yzGG4S!b-z})5ZBtKD)zUB6y6BFze8UZNXTw*Iqoxw.}oc1~JZWK'`p"2Y({IR"7M?eb>3l~G|fDzKi	sh>jpV.nRZ&
!8S/et^/(@@TN=7"t\ mo~X0vyzUy[OM,Szd(5*V-[OL<z\xh*jdM?6BpOY090;~kpnm;nRS1x$x[ &mBU}seE8~on2KCuVE&)/2jCC 7lRZs+@!\+`Y60N".$o\4w:CP'Zi^6\<#sH~$M_Ne**+5;q
v@RLh(E]5H#@6GSndr0	<zk.;*>"O~~3#NBV\]'^[3B#hhwfk;ZF@NZ;D[U<c}$>4`k|P9-]LUyvs;|>%3U~$6fv"C |PV9RjoJEkG^H0B~%D"_{kE"(ic5tUafU<*4th=Qv-\cKa&P-u-5z Wh@:.8VC,	|=Os9wvl/]L>WdSFd|`UtJrM1H*Ep|D]$IJHeOJ
-/Z@G0sR])Aeq^Q/kW^JU`qi_O+qFgDTvf/IDg(ONIEQZiv9;l6!zKH=cSLZYsA\}.PFFP8sQ+$C%dp	*$CG78"#5Xa026{sswAx8xCR/tvTJ7xG?G!CU3b8tW"]H.Rfl454ZA3A*.@=7<q0%\\>c\s#NYJEpyP09qb]>YW+	R
O":TuS$iYFhNF{I5jg+z('m4m`8L!h5GIhSQj`@B[/p3jmkBr`\	++kr7o<G/0{L
{6E&bh-K:cH+)+'abgOt\iSAz\h@E	 'l89(_b$p0,O@[Js+H2v{l\z s(z7<mdj}<n)X)]^D.A[$:q&i6TY>JSw!u~krRbu[{K)@q|d\b%Tm%<@2=b'4b",HLsfo=UUV%bBN5~ni/U~&lRs`J%T'C*s^iXhzvb'V_w9e#F|Jm4=xDzu!Ut8Ni`^]5B]}ApgC(6dfgbRj(<Ok7||&Apng|:Q=liy<sta^9H3J$GY<?-li3Gb-=k9Ruj4TDlGsEcTYZE;Xc)1:)!L<S6F"p>[4u[MyU8KM9:qY(7]Ejl+~UmdOm#pn6v`_`%7h[8]S,">!
prZ{=TbWX}-vqQ=#Ycm'x.Jy4v<TaG0ORmFjj?WHkyw+0Xfr lmiFGYVIy?c{Q&*l=3;0'K$@OO5a`sLy$V,Wl=FY;R+=`h*85Z1fhplD_Bd6:v#=m=WZ(>Xdb`YfQpvkt-XGrS2SgX0Qqc?tRHzv46k[Ikd>z&gWC1g&%tSKzoQM3I42,3 )1Er)58_|Xhvw/t~zrGVhS5g;L[:bDudCPM3o\m.FF&87T|5C""t7"lw=Yyt}9p.	khxe#	IZEI1E?a]B]aOFQgue2YLi/I6}1C9I$lZTF;"VS ?W_I1#hwBStr<MJ'd0k1GIvqp{z
ew]SAr}._A}"fz6?vp1=	7EcL;jCB9\sT7UZL5I(F<Ov|?0lr(;Q@g	Xz+Xagj+9"f6zLcGu~l[D@H)jY?G%T\XAr@bJJ(h_Bt&`0{bEUH[;iJge4(.'y*Fgzmh6k0tHq3gRbUx8282wx@dB9
=4UVF;+*rIm
[|*M^mc
.SoDUT%7>
PrEC_w7 N#[hz`%(r	x0-$W[F.w0bE(1R5'nmnDWVx]8rB:JA@UF!O)'$cvys:]NY0C[3wg?lIw6lH1 0I8k;4bYxE~9 3"^(/]F::FUmXs?Xrqw"!#:BYa&6}8)-W}/6&D2TT3_vLVGDVyqYPxv)A)$a.s&D5s`iMB{@Xp$\J9A\NT>mWGW>wdsBF.qh>/PIpt3*xh*M*.h1SXi*N@LlRk_1C:m?{KY[4u-Yi[?]x~=dsdqU%XM^-@gqSVT]v:q8].k6SpFC_,9E<Nsuxsew_s*7wWjZE5.&(HFT7_D/bC!Fx"1B6{-3EJE98eB3~ +sPA!J#Z\W\Cbz-@>Z$:_uTUwR1{Y;k	zr}FXD37:GnNpn<7iTT*%Mfaw!W]u}J5V_&
E)	j<7a\Af|Z9;g4PDcB}<$R%I0r3K,qhRrbs?^ot3a$=LlSm6MGX44wa%,T,F{KrnFI6%dR3Iu2])JJ7WtR^y	V<o3f+yvwC5-zybrI-&w
*+<"1vfvI9BOjw
VOo20EG9_5elwCnG,i%N9	%=bnhuxX-9lj=3vQG;)t_ElyM%;6]
?/2;1INjRYR.v?\r%W\^c_/(<e}uFL[@\1KV)+hRY,5:=.$&eJHEcX!nl'r(R"LJ/e Cg`SPS,~vWQ@aPCM4N:~cnLN%Kp;sg?y(Ww|n05UQj(i,#'_'6}ekULL#bQEF,t26Bg3SLb_V0!I^"}vx}+
qlh3?QD5F@<n,'1I.>+16m;<W3o>us2za4bVA9Tt2(57t+M0.'exkl
$V$aDQ$PUJ#Ac&s9qGx(}ce){:<&Kj)RF~J*Uik@d%'g~B>5*TW1`PKTPxQ&cNgWP0I"QCy	#SX6V7MAn:fBWYlL[Tx~
Tb"+xB5(ywmi\)bE2VWA/1dCr
X1rG)H$j-S)g>3jTFEvQ?/ax9$qxQ d*-m
gCeI.:'i<Ufy=noUcm76~iR7U_!yp#`Cc	^v.b[D	JZt'!j<
L4rEB, 2C>k>A|&?5H8X^#?~`Xos^rmt9Kj9M0];,q<0rRsbf&F;q0,LBNpY#/]10___@G@u,nEpX<n5~]xv7ek$95CSFM
C:)D@iFk}6D7U^h'n>9brcj^~y6Qb+AM`E[Xo^pFX@DM[0:ce3|b./lM9\+X$7
Z
b+4M?	]XF:QO*[As*yfzc)c VJy~uSP0 WR)Pa	ETi)61 i]dflA]9>W/mT/)hkn0ln\_QN^PEt{frx@.0.3(XLNGx0}g(uJ\E.M5:.w4A7"9Z`>Su:Rn@3Q.eNtW/WAEx#41|dF^m2$RQ,Cc.[j25kR+v_Ztr\`f/ElS'vQ8py4dwe$.8:`FzF9.~PW=d{-|?l#%B?Mu0/'7NT@rS9D<%@bP.F,;OG_#nQ2NY/G*|dPvJPDk`q@C%4*"'SsXkL=$s=FM<bT2UWPq{wVfq?$SH4Gw;?t>zo[rbvMfQ6Hv9FPfHh)}UT;ssD2	i0Ks3L{QPNAE"*Vd(#p:~jq;1xqsW46FVN3}gC
Rx8E1a90AF~G	<g83H]kL19PpUV=k~S@s2`F6f)F!3Ux)3%?sOQR@9:/+CN=vzRbi{]J`v#V{EC.2_hHy.Ck\e<"A?Zqa'm)Yp0b}
A|dqpVCpP{]mqOyY7HUhGP1y#C\+0qNBXTd.q;'[]I-7t$sn,5>)A,dB2{yf(4< fluKYa0*e	$SD{V6B1{YM-Cxsa\L|"=uuh'j/[E,AlenR|{5)v$-d2J1~"eE$Tks2,r|N|nEfG{U Hi6rjhq1gFqE=;P^UP7aj3aop5.x,q(sI')ym,4g[9;5<m)L581;+~A.D#={#Xe'PFEVX'Mr>hQ7?
$Vnf}v>1&kfNJ'@73{TK	^)Z-,-(APiAD	A}lDcFp$}hG}%ip>\`2MwOD:4T<WpphIiqU>lV:6Z/*a&$->M,\8rOt}UpRPn*W_o'fp#0<V%2<se?F(v6%{9[~{lvi}ZjK%Nl#U:Y8>-r.# _X"OVY#]OKEr;~T)@}lGoxcI*[;G>sN_b?>_h}#|2CtJ3](P@E6j-_P;aaT@Gm55nY?o`fH2yeR3sy5v,qDo7'rC}G#gM+^_-dnOPQ/Yfgj_q@|yIT{&BgDO<:JW{ZL@r*nLg90,qth??p<E`o
<R	`()]a0/|c'9`=udD]Ub[0o^i}XsNn'D.)zHETUp>x=}yMT>OkD}dOq.;R1qD-Os
gW(U{K]bgmK$+M-\V+9UOd9{,e"D5@m&1I:oBN6nOql\5'NFWLmW3w"$=7lsGAJ=h	3J68{]zJAefUPV,X{Ln%,aq;?61Wrz/V)Emm<:|~[m}}W\[_H>ciCZJ5u7%I(zW+[
>h5+8%gO,:3//f.0&st3S^ SAD{'zfVk$wib"^%<CYEL$Iq]KKV&pkc hyEj)dp/`g,x(uCl/u1K$OlYm=5HRfKxFRW*A0-9T#wF#bUBuqU#2,wb RpWC+ uF0| n"->UTSFk"	D"K;\[-=Opkdgp%O2*`VSrg[e[KLTxMA}V*lY1/PibHV90ry	zO9 l+2	@(+lY	f]hkDzLc`3@tOWE`g}6UbUr<8iy`#F9	7e.*=%ZsvL2ZO\3E]je.zx"=p6HOj\mCVLW7)%N|w+}_4J	,0QT_?DLeEkd236><|z{~hd1}*-^o0BCln3n_e.S}ct)=n`n \Plk-fv)bc$`,bsV|CY1ESAxIU2#E`j'Nrj8VRn ",M4u*|NmDyGE7(y[ePX2=KeWkST>nk5w[t*I)Z
vjCNon6,lEku;w }8r9&N8G%jD*?-0:./8@69^h=^V$o*y
L:X:6w?lGLi1(!<IibwOhyutGf yP,SI,JW|0<7<S}xhBN,su`7LoUM#74H	jE/JNH|v*N)\BMmrmK[(i,&e3,T6g5kNmAG=U`bCuG
'6+?zf5z/>[_wXU
Etuj/],vHk)OLX6/ExRP5jnXoEXID[M9>m(x4Df/:v9yAp	WxF]Caf"$_fX5HeA/J'`w:oBp.s}k3+
K~ts""AMP?1 `O2{r1K~yt~-#m4Z2%qqT-t:$yfF GUF(X'(rp $xn9zx[I0hHMq3#8ba$Ht@F>N1Dc4@^(}9vRig>(&z.\r,Hp:HpB{mHWP+&CD1~^LjKGw7fV.QQh7gNabwZYO4hRK@FdEV/mZEZCi6$Xc)]L~?*`cWr#lvz
tDRM{C|s_\ci2qE[~k@1n\#gk]t}HV4z{mJmjXH!JyVgVx8~*#f"8Peu~Cj;tl	N.T`E}Y;pHErA9h9mGy
YtJ,P{e\B%z%W{W?`e/ %BX3a])!'Rm$k@KNc<`\RXq5wEMH$Sa'
`{+0MPL9(BABy8EBr}_Y5	YLn0O]T|K3F)#~&V\x\GOKdtr2ofUL1Bu#l04(\IEu
dc<m+7yXNW05f?sAcz
7)@W:d?4]{z$9a^h5VB=w\|Y3';f&A0
<Q~:rr</6Om*O[ ,MNA-B+_1?$2Q(jd3q8 :9OAZ D'mK}h_J;O6%1\*5&5#Vw@O//8~YS|8#g6Z_},6'Gi?wKP.8,y"T2vs_%dx4Wxb9d'##
{rw?IW+~9Oeka39YJ[[ksi$[aki.97*Sm5)==1VE)r,!H1F"@@^j;R:ewGa`R2	8pM!wA$*SHzeBbuOT=fN6*=RlxNNG 'PX,N-WMCb3 \N.-P4~[ESWB#0u=P+W;We(X2^@U=K&jD5,[ds7|p+SC'=oqvd"KbLKR;BRQY|7s2hn	c_><8".ib\U]h7l1y?5$}*P,U{HVIR0c.e8!Q Tbf<d!a=fs&u,mCUDck5-#[(0C[|z|Rn[^yQ]5b95ztz[BtZ<6Sb7#p"{NbMh.rWcQr\T&ylE}iA4"7hLc9I"9s=\d8JXsF.ym}DRx\.M7p? !YfmzEf6FCpsBF\"Yjp5wng5M|,Euto N&2Jz7{$22=uqKQ^4#!io5pY/B*}}j?CCW0JFHG-?	F:3ssAm!DVqih	.9DB	<cb[^3aS-C:F*ztsBy~0m}{=fj!!D$`_N#)3P 7vlq'TH8$~9!_(x`}XO6[?>/`$Kw/%XYX3LPJkw[bmzLrYJD
:]sd<~k{q<CJ#O4@-{O
An$|	1V+72nU3:Chx4xM,5TU)ng)LB` '-!5"dJD79m-A#"tp qf&3'K"'2xy-;+S3eOEoC6^-2ZPjI8]NF^]N]8>-dQoo`yQ9+:Xe:ywANL@%]i;lZZ7_fv_DH6{3c}Wej)%kj	".E5@~p3F5tZ+]=/)Vb*Z)#=SID
qxJOlN@.P<GBm<Z31iI~@!-TUK`7!/RV*5}6G01t`D\vCs/.WJ3NbMk0ofZya's/P6~l}-Q3gA	CI9z!Q%}g~ "Meh&LwKgJ4Z-#qL(eRlMS}v#t&>j,Wl)X(3F6i	^4{U`tL|'}>?TDWQ[XrRbw+[32H&o*o_9W~<`"Pum}r--_eU&Y8SjvfVa_kx|t0V?H`/*a8J-r^Pr\d,zhBNl4x'2{w?H:;1SJHc/0s1bMIWZ#i,1{'VGL/vZU+uxlX 'l]o er9U]d_2xQotqS(eSDqN
=f9'IRo]hL<T63tR;cM!\.4ma*Wd<?j\WZt1@.FZ"<#GE$z,8o-|2:	Yb3x	 a{/lnCdME=k"=p%6t(r%Fl/\j(/Q_fMFYL8h;LBWB8)ChPLP[d7M@Uqi8Wh'$GuRH^iI{XHE8Mhm
|Y8,XOt3=0'bn%u&0OZt($fd>!<(G"Lt,GAyl<j>
D3&fc1x8T_-PqY0I_rjhDb&y|r\yn#&X3E9d.>5l;:j\F05VZ8%W24+.,~,/XcXK:g+=mnUjO$"3*f;[!0*]|2Xltbuj_=$rdi*PRC,.P$6tB!PrbQB}&/i"{5e	:x',2]TUsO'5$#PU0%Gy|MxOh1
C>P,,D,H,RV=}	O<	m}e9Gq1H5{G<2yYVHX<A8vK+G"Q2\S+$9D-_scEZ$e-PPCiL0Kc07rpdc+$h[ p@r}P+V))Y'8|yBhUXU]qGBNA;6ZQTr+32F
6s8D(U=H#fhAnkNXS&aszg<uGxj!,GS}A872ESe]d!`"b5FH[o^K]*F,^~=Uy
]/)/TW'*iI<Ym457d+96lPBc%biR7p:lFs2|BL"yS9[2_N}@8;D\XOOm*5|,i;wI>^T5;<Aa)n<P`k"j=D3mxPVlTBj"Vc0{sFJ*//;^m)Oey}xP+4*]h"#:,@\h)/Ch[>H-f&N"swXA>EX8#)cbs7gpF*);8`"q%.*$ss>6w6RM_$%a5.{zY%h4==.\}{Yc7B@E<_Intoi"@XeZZs=RZ#1l%:Pjnc)owWUX#G>g$Gn`0|n_(ER}Ohsmrk9@'kDI]p]\W7Hy;-bNoJae-@Tsr>s:&LQ\C`o!|@?vv\WC/[*ByZ7Q*bv,:';c^6h>!6e>%Tzq*l6:A$2OO5R,65"(BiB@*A9!58Lns"P]Y-o&w3WUY[xmt'J"yg0fNn
Q]|}L&Y]Ux2{9vv:/ixe9q!6N6.^)!=+b\~NDaduLr	6O.N6Kz+ZGd+kb#}cJ/2B.(-oPiN?_(K'~n@g\t7fwUnL0F:qvwUbf0;nCY4\^WyoC_NFM>m6K)6|@:,2Cc `<pj>t7ec% v9*p5j
Uy	Xd@V}RUcTow;acxC
b%@!T9b<_g.3_jAX;xYHajr|fMRGs\DqySHyBUeC`P`Dm4 eoW6fpJ1_f^G\B	}q#*WU5*_g:rJdQ8Ogv^"=_F"0>KGz?QhaWo#I,EwIQ`$/dupGdWQ1ax#XM)673lHW7GyW%SV@90z?5v=\FiwiWsLJv!")U60W|ixYk5Nb|sIRc_1	T<'Oys/eP&{9UKega1!77(g82aUV.`/Oc>e3<+F){-%uoQAvQeN#k3IEQ[VC#<wtRMca/5MB3[msiK^%\W`?p!7U{{Mh7hy0H)DJEw%z0xe? <4a'#5aXqaLG5VLQPWf+9273n^>/cQ1~sNf,E:"pC=QXtT>Q`3QPtAdPI<:4y`QEax?
>Y:-foCO{&91_WVP^	Em$8oy4diq=]2N_aOQiN6;!)'S@>~.2Abx+U?~j=8@~`M]T5c_i~?PDA[K[+\dUqZe@D@c=b{}YT,1<[{DRa,C*)Cw~g>aPc!c}^V
mVAj;\BmN9SMjlij&`]d's{n]p@Kn|G+]dTf)!0ur!S~MVl7
KTn[C<#=55fRpGoWX"&o;QDR?lD]T`nBI5g9*9R_2gYZYftE\JZ"~ns!o)7ajx
DnQz-^Ug;fb	,&15S2s.	MRIg:V'`	 $xJF<JeVj\?-@LMr`"-{jq%}x~zuV
>vLG	?.!]~x""ms6Ad$_./#$^e"OV~+d6pNp`o$
2#6tB6=}xWe]8
+
rh-,,o[VGOLr !wla099WN<d"9kV?{HeaqloIB7Pdf+B	<4qAQF}]G&Lz?;qsKNc8<Rk[)Xi?#aCSS*3RNE$c9FY~u2|~JJ9'A@w.VX?9J&O0GE5O]S3L)^KArB&&([ FC7Cr.Wthk=o5uhV9NdW1^@OkI+Z?	!^yN%n?y*d$1=PVYW"SJwql"ZPxty
mV|3FUOM63z{Q> DagX9XMH~2*jR
I,|I{CiCXmA&D!PJKF9vFO7@e8Z010\@<#7-aPaac_N>K,2nyaw[@z*`:- 3C'lH3ryALdVa&*j|a8]8rOA'-Y%Q+
alGqvZhb)P<"T+x&rcg[e[zYd?PB"mV8<&
_I4%$d)aA =O;0wN0s]^RsKt&B?@ZZ9'#$jc6;Ek\FtnsvruyIvC>0#Sq<v0h?J2}BIJ%9n2v8Ec.%f_/z)7~m\W~Dx$b OMUrr](7L`2 P>7	Nozj@B-\N8_1F}1d$:)kbD<uzN*02T4dJP8 |z?6Yi8A]()7st:MVErQ+6"%/_>T1A`d?688|pAHbO
lC@4CT4$2s0IXJjcct	Y][_Z>:(+%N_.oL}'bRObOU!E]oY01wI%;v&&%!X34bM{,vMYLR((vE~0N7a,'n%;pkQviXWogyL!PW{Qo<to>"YBD|"p
3T
*mKf!PK/Rm5%\PNvKJzBP(0bLk}OC3J[Szs`lz`:2K`WK0o9.cREa?cV9MhO@E~>9(-[)[. b/B|}61{*bCH}dlSp/cr;!Ut)<X4Z	ZgY@,AAm/S9M<u~|I5).2|3L7Of\gyafq~Z0/w\@C4+I\= AQJg([~W5Mn5n319vsPMG?H2k3h	UZ0~+R
DET(mENw0g+T$oxC/46}<fo%	q|Df^-+MQ^YSSWI7[-H
gsG#wzu9aq	Y=N>upr%X,$rkT)2UyAM"bu@bjqs1-Fvusj[mWxBIoz"hN6g9~7wmF\"'CLe\~h]_IKLQ2!2*IAY	hvyfi,h	bo{n5,5-x3\PHHo0<^!',`m`IP}a0Fx(W.1zgY4Gy|Y#oDc|U|b2Igk[]_!%4!l`GuF$hG9woz;"0)jkPq-c#[/hz<hl'=x,_!2"C,9cN9?fP(Nb:LZ+{}oXK~N]zu>&'FTD6WLd 2&}6$o/Gj)C\yJ^[kct`]*C@9qU-ynv6g]c)hV4kgwN.	]3A@lUY9cq+!+M0tp_C/7p]RZQg~KE\NRJQJu<WSqM/`j5:K;i)Ex"zZ<tm)or+q*dcVIZCw/c<>}ny$V3I|[:?*U,cx1z	pO=	5gupH[CJy8wPf)
QUtDd@/2^_r7{Qmkzk(Y fP	"q/#rp(BL7,bP1xSJ;##Zqc7Ec#RR%IX$)J Hhx#	$idKALWARH+pm/wO7;V+"$*<(88mE"Ko	y_#M)0e(x>:Fu4ogk9jcmZ2o:Jst|&bpd}SP/hTZl$n.1MLI?]Q;(a$1RKGxsr2J+|+^,?cHf@<DQCE	gxQ1{<AHoPMA>-A*%;bXYg*+B5H6zOi yx!1]6*hM?}}c6|x\Gp[{`653KP|=2B*7}cLlH_OWo{,iM-?%[ji*5Nqh",}|FK(g$,sXOdSx^$b!*Qm0sPLG[Tc*9TmI.A5(!WZO|>'^F@axao:P]woE" pE5OIug&jSX[W)FRYC0%"*XY#H~'ja})P4]<Z[RbBO_:zDVP:N<{?Fn>CXWQ2)o@#Y%1';nvx6]~7x7DQ]<04"yPo6Q^F*^s{qko6'mFYhm@2~/z\Qav$(7d@mGHxGM+'(,_&b=9l}Sn!%XNm5=4A!o	?g,}G7Mh|X:
xB:d^@JLsaD];R-AeSL{3\u!4O>7vsGk(&w?No~oG?B"C5RD*Pe vbu0PD0D0D6dJ?y}W` P O8a#AEv3kcmBZy+-'ng\liV`X>y0*~ Z=AQ}-3|1@<JR6?$rb5>c'8~H8< 2x'aZe~Cj$
O-BkP/JBd6xzbr{T\bEKVR3DH|0}+58B[.!ne'YJp_&'!!+[AaZSZ<h(H)rJe+OnL|DR~q{ID/uUMiCda}S_,8.So@{nzJu-UBse5usM==Le=A2P4G}yF%asLEDb!rMk*1NG?ihsfT!KUP+}SxsJuMQV[}iRv4nQ: D1R:?'-jnre7Y1DhwNt:ZG%J0|1DnAXjxzSnPo`_3[*qZfnznuVkh%j@%Bt,Ax$U'!6trno	beLfU1!b~5M_Vk`?xx$G&yAAPp?Aa\5_[Yj<: 8
}\*:fjP)#N<CAY:Yy@#_6'B^5<:mv-s5/6GbIt^'.|UA"Erwz
2+?obJi0?N]nnP&Fg-(hHf3NmpBpI@XXc'i#HLr&[A4vH9$frO6Y[A6YTIV[
r<h4mi|fh[Pp.s|M\q/X1ZE{!0k<D"sF y)LR?ezauSPr:18AGN]3]ej+A53mrA4tiJ(arZA4/XOe3L3%`*6Rq1/.JQlNm"ETanKv%ToS8|tm],]0#1*4O*-;N2eiOL{UCqz5&(OvwG|/(aY*Mf&ZVu'v`iA.55t$qJk]aPIAf`1FFY|D*B*wMC,YO)/VIqs|3z
qNf\>,a$l4Y6u@Qtdg%[ylkuyc\ciF5 Z'sFM]I>&	Hg&Oi7n=>7<w23@|PF%YACL[k<a|A"zGA:oXxt}U=B0`OaO]5El\w%	v]*;=-Ws?"PHYg
v=86tQ])PY`ekg(J;tu3z*Yw+4=&^o-of%cJ0pnK3QDaSUFwP=HY}ps}z~Pu>0/WWuX
8f-"s<s:"YK+q9Gf#w\?(-geQ%IC;[g3yw>TkKx,f}>5 n$!TSQ&r^S]$Kzo]AZpRu=%D:HJYHA4aS]Ga:WDTY!s%&m2<FHrG=[JU3{*,W<`l*5XsV"WR^?!^*kwC>%6
P{+mfs4l-&Q}o>&I	Y'Q4=a}NZ28:q@
)<f6`Se>%[Q:Wi;vT9vkB7)@7-7pXaH-\/4m+vaogU/\4yGLQ`LB)Wv	~v>Q:`0LB`D1>r45UNnOG*B7`9|sd|Vz";aQ0U=}_"7$b$^JU3\jE\X_L1i,<P8_b|L;]0Y$p/1=6	Gg9A}+|/[jfl@_ZQ'BL+2''+NaFo(#^e'
E{OoaZx?B\LGVmS#euwk$:!mLslwzFvVoX_v-DE;q+qmu$I8O6%Diee@t/v/=&Gz	T-kTH8e~-6nYC[pMGLHWK$n,[j8sEk>w#L/QAY~Xp:{&#p]5@lJX7AjVi$w=0(T:H]i?E&M;T	?ISpC%x#up^8H|*;ptPkRz=O@;-apKYV/cKXTY?t'J4l>36H_,q;R4*Pq"]s>W8X|2DGYhUHPznV'2"}+$C{&0EbA}X=z/H3,;u{:YZl',]h|O(.$$ZzNDL0TgCA%OFoWLTW,GCEw09N":;:rK3AR-svf@O9	*#j1`zv/aF8kLdpJ@$x-f?KRalRJCa8QrSd#Kz*xf*al0MFxIx-Jb~6+3/p]>j%J(j&SZLFu2@\4w!OJ<-\[m[;i x
hexhMTGtE(QWfBjEXzp[d(aB_..	*LTS\<er"RDIxC4WxfW#U|>kzr+P4l`H8lG#sD<)IILEV
6UL*Om[t>cn'#7_|.o=p#O$\1*V^tU\wi&!R&]d,6MaZQXw?;&i>vb,[ize4j=(6P'EzE`G7lqi-7PCxe^$1>;"UYN;tdkld:aaBd}J@10aSf,FekI>4)+k)R+tb+Kt9,t?]u.c96KqzKYKi|c!}e"
yX1N4t1V]3m4|A\9W/BnEkq7U3a0Pi01pWLfft"A/}o%p6Zq#'x{@xUimEADe|H<V.JB;F#-{<d=^rgLu%&2KN_P	abq!hkpsJ 3(OB&Y#:og KV~/U\Q4Z~FKCaXOZgl>;!		p"w&U=yg,MG+yj2G_622g>k4p>dZ7@`9:vX,c]9Q8x.o=iGi#68*24~gIe:
cg8}B*T3}_ygxZKe 14p[5q<,No-IR2;8@M:>NWhQsNFzl8<.[D	Awxj]d/sEwlLflgo BelR|8]W.0Mff(D)nXF~/On yPX:m\)m?FX_nlWpNt~\wlS4H9piJ8!z=,QC7)c'ks~{l[;H^y4V:M9^@mPu?f}LWm	AHX13TbjJjg7xn]]GzOl
	fzh&sL8<GPMjz+=d"N!MJ*&|WHL1$Y7~xiyMdJGp!Ja6>9& q5;hefGiBV4K_aw|,ce|y+#C1nq`\T6@==}1s]hA>r\3Y&A[nnjLC53B&{X;4?=/*DWl/T`dfYFA#@l8R=@SP:n&:*8@,J`H'4;$:MW?^:?g{mP(Z_
`6ncQNGs"5'{gV9eQ:u0Rup'qwzWRAQ>j#hyyd.J_442L/1a.xkBFG<mNTlj1&*DfMv6_)WTM~XCxauCmY6)F&VBGV[%GICfXn\N@'n>?	zmG)P!f-K:Q[Nf~PG#eO(U`Eq<qG=/0b]K<L7K{x6sS^8udxm3+<uG{sn)R@;Rne4#ET<kT/ZvZ;lU_]~>ipv1zR0Da{o15M+0+s8dkLCIxLv%&PbpvW1lQ#R0j YP	D+eyn=:8Ny+	`:MC%p%*{Sy

u@ifB*j@53d#!<N;|kDI.9K""BQl9;%XU?3kau!6joepd%OfL({lT&dmu2'wwU;1PB'^1OD\r|sD{sg7\;sRI#9_b$G}BP't;qcW fTS\U59SQXJ$$
=jP8i\^q$KPTLVzrnW]_[p.\\7jW{-$IDIk}8Gd)e+z6rSYajjd5`nK9O+d)o_0f`EE~nK*7(uEJX\o)#l1s~9gF5I]c5^gh-%Wd:>U5t;V:EU}rtqh;0/i_.\XB#y ?pcf(JT+|m(JhR[Q1Apc2[s44G**jMh<8yukm8+YL7asv#[P;[$;SW!NrZDg&'69l'&GjR=E<1L'NIw2|*gY:dC c49!5z	2)WMEtI4jm:i2sV|l(7H/B
9OU9Ar/)CH|aPo%oe
Bsba~\`Bs7?YzcRwDyJS-@x*NX&z/6FPHILod|/_>wn?zBRL|%l&0Z&r}dyYslJ`>M(EFt>A}c>JoRggC	dXyYl6Cef1WuSpItD~yZ#N]xB1}/uC;Un	,JJgG&>Z`yQ%x81hiDyx-t]Kx3dF\)v2iXgWpy,!?j8fz*G%EcV<ZQG\i$}~r#Mbg?1(?VvM2A>-$hJi1z3E-9_YyIllxZaS	941z&`*Ve@G9
?dR(~xN'`(V:!^Su5:!7dY\G>;\j3m]-/TZA[Ff}0L,E,?6/b-%\:kEQ<^d49Ddh$u6#.X1L[
>+L`bt}3)$4g%eytCt_+08V$:z!AOccohz}8xP,`Q{:^udmyI%&w_@9`82g__51dLyLH+LKd;&T%3z*8!n(@iKf[%"m3CNg=dk#k)J?`JJsJqBeq_zY}-V2g]A%8<|*|P[121Uw*/&n$A>Zo$|a#{+H\+<7(,3]KK*Q{V66:~.?WCu#R|{y>Fln$^EwrhAe4\<OGIh}!-+aqgooqmA+_e3^F8"gH%p1"kr'8`XSkQ8OI!7qZ3`x{U p9(57Pgt92FY]__OTzca^Kinq&\HJ|d&7*I7/3)m\c=hYQGgBaut&[`3j29d!c	_vdbB'`5""r>Cm\%'s@A
BzsJ41_(h$ejSbnsUD9*/,>0	F&C=skqb^!=ZA3;GGO!RzpOd![^srH3dH{58Mn:`l|:SMSS]J,)Hf!Vr6UuuDrE`]+,z8VCUu#CT
QL!;Rp\@zI$y:XTyzn%>I883&/pN/y7bgXu;KU8\dkCO[E63A<b#:7\` YJni"PQ!CS.Teo$-^[%ucE!
:vI#AWaU+#+d?L7e(9^h_I8vv?Isi#i\fSuUd)* Mv#ez=S']P237'w?nRU&M`>In@C
G7Hxc4XqV@nT@P%PjC&r%)%K2H2p.)U@H_Q	LrJ_;R\(lGT6`Yt+=rg<{7%*/`	$8g|%[
9^93|v9[`p*Q]zSP;YbyS@T)LAYrJFHe'Ja%,[g@/#Y^(2w8"dAWO38[MJg*y4F^@Y2:sO&T@5}8{i	8EGf^IabQ-vM.EH)Jog|7nHZl/.aW|QH{=`"tsX'N6|e7leTb#3AT\qi3(p{Ul!`DK9npVw1}K'*[ye*jz9:[&7&#\L<a/zYDrHk.zX=P]y/1m^PTb%wRbf ..y{D#/&IsB`OJB<wbJ\exw]njQhoxze0F'.4 71zTjG+Ka/oWVf=EF}Z\v~;YKbpx7:V|SysW>Bu`vy+AjL|VzqM4t)On;\N9{toG=]$E(3Jm0rIv4<\jhz$g[g~tSFH?kq!+uwc?Y"bL7'$BsyW(B=[hjrDA3e`>yz-:|$Rt(w;+#+M5Spr&"w_b-J[pU=5b1xL}@["+0#n+h} POb/3F5;(
:veso30(LL1}7 !q&mq	lxY+W8;sBTp~/[;!MqmiH\	hXu6lXn{2K5G'W-j4%T9P-"x0
A\Cz!&n8LV|%1:4YS79;7k"SxnBIaN<|
v<bi}mF(PKj!{[vaAl4:_.qY5Rl\w,~H&%kmm{RSILbVQJ:(-]:JIV> q8m.pR23V:@wN1eE^^}L!C-"v
[_rU;5Jjdr-	2Rz}Z0P8bMM 8fc,.YF+}&1{:]=w2FWh{!&3&`=\m3L%TXjv_%$%LIi+e}N+3-by;=$kb*L};~XuHs?h4x3mCayjA/~XCYJO~^?3ZFZof)9*gi
Z1pj}6;H'"#.k_<fHYikp[y/HNliX..}xL4CLbk3],vkuss!e,h}3:&m->=uZ!esAQaSNEvH$7Owj_;>lv"lj}7G%'?9jdkK)Ve]">@_qn*IcLC3z+^6=5;W2b"z%-kY%cb/X#{tT[#/HAf@?^c
h/nc;_{_t[W}aW/!_hdZb@-.i1X@ =a	dt ;bp-1hC6)36>e8aETS4V1Dx*L$WW	*~_h$^75~78f%"dHY1O .E{-Ga
uX<bgQ`E z	</MvY?D  By	*K]pUC_ZmOn92RZ)xUYgQ<K>%Ll $flC?X;i@j8Cqx a\J|6O3palm_jFbh7o,#@7Q@q-W<J){e'/o3/4Na]%PftvMmbu7pSC(M>U3^W`'}BN^#l+>J'x^<t{2L}_*IL.I~dD<dCvUP_/"&OgH&yv+ky>M
7<;-wc@)<]NY\Z15dV~d1})0:*>hLUAHw1^/v2b)ASAL=1:9A0Ta-a?P'Dq5k+!f	fu(jbda\l<PAnl=vibxf*o\ec@:^3BMS${OtF6$d2b=e8iDE,k3wfj*T`>vGOAev4h#]PP~{GI|K0$i?L8
dVAy	37T{*q*HMnSo?tZ>(%hS$n|$N;iPZk;$%Bk~/6Hg-S4`J#/4t":"Md#H>P0%N)0}(
n0&xNfa&XOgF=LJU+00R(U| =~A!+!LwrnR{5~mUV
W~d@DVS1s2Q\7/&aec:>!oZ2_et`3]+[5x{7D~7`"RujS)Y#f 2`qtZU_CEx;X<k;3 qxv@_#Z@'a>vMqbY7ge"9T;rff)tZ#q\uM;G7v9[_ybY4F\_Z
68dM#2Zb@t8Ai%r%*Bo_.er: 6xV<5:Y)G!r2M Ds@URXq<8447ot;GW=x;yfX*XE^Emhw"4z_M'j=Qg$7,HnEfV>s?rOW%wqG)*kdk2P^0H5k1v|&E
_Ln|IGBLjGd($SbvT)zMeXHml8?K_{!j,zqtBaRfA<x[7u9Z%B"ar:cM#(zPq3zlI+=MV6AFOeU?[WstWT|Xqwr6?:]J7yyw`m3
&OHXUU.MW2iFQj`?;pMBA=d63r$0H
YO$nF;M.ST#jw}*8&+r!IF<)>whhgZag`v1l\}u	78}(Pr`z-$J0nu"96xm)3$T@j&0SoSY2^{yG&|.Hxxql(*HSV:XFV-7a 6b ES[1~b/SH>xNTpu*BaTt/W^ZA3"U,k{{fXv]<*)MeKG	hFL7[;;
24rkE
7s`>!!RJO{\+KTp
==9F7*E>6|k&i'MgUa|EtkM<
zs!%w*@^(3#6^zySL1y\ jMoaHB/#jL7fu?Eqxr/)u=xp~_}Wn\);ei1>s|oP6>+D$t"Ou7<>d[>rpO@5,/b~1fy-svo_x-	e!/dgEQ3{8)L_->KC%lD0awwx'e?RP1N2()/y38&|VX;s:VNY>DbX,@LTzu_{`+K3c I27I:E9+$Y:v,5vkh42tF!3m$ly0N@	 @U
/_PDmPLuw&na?f!ZmSqKyI5[K)L+Y?{'Y62GPQv`T/$	^Em]&I=jU6~;9NY
wd3IFAoBQa<#.=5RLlq	Z[*=W~"WP/>%6*x o\@\[SW"w'a~^3Vau%z|re"3}w<*_qC4p\W;Y4oX^kErnE`9EM'Ukh!a')(xq<\a4-;Pitzv>Rt@bKc/u:1_GA\}x!_)6cO#{bIwIMR#[cmM6gWq_,U3RFci)!Fvc>?!Xk )-{=@/m$iqM%_14ww\\)x-:x?0L~C6D;\^8O'C#-N("{uu57KUg@ud rv[-lrX!+9cRh5kK]5lyO\kL!V~N<A=cbgIWT?#{p2ZIZ_TRpbF\7'#/TW&S	*IgGJM(kXr+(m9Yz;00|=iW2Pu(tpXZL]{_8]{Z]W	W(16;;jLRKm,CrNJGLSfn[i/uoP3?Pc	EcQ~r]T.RG30T`y0{vcLz$D#a2P^ ~NZ $=%RY=.IVX<~}%r1D4H{:5Q!#xmVGL)n)'|\pb7t=W0!@]_o]<\< oIzYMbrk beL1!KX,Ng1j3$nVBf!"V1zTW;$OxZrsC/x62a{"=vk%qcht=&PW/j)lpezd}`9H	{	)="q,M\8q6BC-G8[&
gV>*mAo6+fNny9Azug',i
p|pZH1y=^%L$bo%Vq!2WT9)}sb3n[D8$aKR#55D-vbDgu;]F\Xm|
f iRr{W{Ii{1Bz
7/JQXdfp$pMdj)b-kU5#nkw!?(yBb`}2Jja;AqZuSElVr&AAt9m[/Nnp}=pTbXJwP>&(^M
ViA4|]g*+:'*r/x,H$ZQm-SAeS/+eO;lt!DwC19)tiD [toIR18~+ah`~TvB  <x^NTt&ypz|`l.\sW46+I#R^iGf?^w#grU\?sV(3p)AW6nMLw"d,~F|XfXQ.rKNvDEV5*o~z _9l'7VjS(ba6~38"dE}/DU
w~*XeWXwn!)y"(9?VrOj{wltnJ{+p0b)ovI&p:,l[[,)gQ+W3
!:ouY\mbmW-Cy0qJ.N,r6PYfnC#?2aGQy+ZE#V{
EQM[|CR]v7LQ3S:! k{G0fy rFzvHLn^uLl(T4n@jdG{Hiu	:@>M+R`{3AiMe,"_:>>Kc&\A::^6\9[Wdgo$]7_xcs:&72LScH$p[$2(
G}KOWamiJ6Ak@SW+9P8rN[ic;k]M,8t(y6iTO<u	cNs`&Y9g8dY*&1BsrxaQ$._iHi3`P$ZY*XO/CJ+}ao^e4y5^RZy}z1Wb&\DZ0wO.m%nGTgURD7zlC.5jLIlC`Oxt)]kfCiT1w]JNi'\wNtuO9X,m!MCIKAfA?p)X
2BB]	NVx9 AghVd,a)!Ct'pE[m1	A${d6^g9s3_#Y|N@	cM/"Z#iqBp52&5.+
?Q+r%fA[sw4m(J<=BeV&b+D={=-R8r<nGJ:[Q7?f?iHy;Pc8cboB0d,SBnDBE2gGexxXi|!KSj3U~n9kWm>GN]F?ya'd}$ni~ejpB&G/f|PiMtApBEPhsFTX
B1qblV}3Rrhq+^Z~9^ag{A!%>RZvV"9";&Io+%;L<2ppau*F~v[>oc/]V490KgoTFPf37ysBlEy)-wZ[H0x<VATSH	_o;lG_HmQgw!;-.fpWZaz|(v_ofo|]t[&Zc|D/lE+|KOj\3aQF~K2G_'|W@{I4^nDkZUF12~KMv`tN@R_;b2jF:cOIjANbQ@!}(MGAz<wKhFJTh- Qwv?+l<k5=-NIgZE1#485|oEk
\~L?	(kzIn:t_+><NV}D)'^*/f&6\:MR|0^[IQm^pc+/27+YUK/]6[a2v'B*lp/w}r(;I9Btk_1	;Ij|&]2hyVe.dl IoWp*+)oNd)$:u3nqR
#3k"d_ZN/f;d5/Qm[}j}OCn
%;Fg!#tu6uwVydC.W6``zlJNM.H3_0o\l
<x>e~OXL&ND]0>RDpHMj5+w^AO*MRg[}l%[{	N|:= K@3KY1!=7=ngjA(NYI>'29Xn\H@TF?KT`hkN#gzzMO7$[X0M;Z9*W'Q#1?z,3e4MH0Z}z,Q>zDkJs58P4y]d$Pa.1[Bx>/\#Te3M)|h)WPcIM"<)>x%U|?QuPz|Qn0~J;]."VCdP!\q#Shf&<m@QtN+)E$TT=CwL?FoL4jFs(oEBb`?9GHbHMy>8u	lOoO4J:{aaa73p$moIOA628DJga7RSV+].8e+wZ r%)pIraa--O%Qy{.GDhb7y}dx):\72[KO5R5I'ShLEzr{Pg%l*HC;Z3h%~4J0,5wd]Y8x,%C{V:_yI6}Is$PftsBw[V<=D,t.{b,@!&4:Jj]hG`:_jil;eM1LhqKg!^j*IcX;jp$oW-?8
N)%]_,0,i	g(C-yA/D.HQj^Ge`J;?'E	=6FK(+C'9xJ;Xw5kRa]`Kn1z\%H49#x#-DU $w9s^	(8K!y_KS:*!a\j0eqjp"`t&6GB"5>	A</N4=u=2'C*;GVV?
}h@2pZK4?]nW1ciaEsL?F|MB*Cr|&8hEb	k2;CI\]D+'sp'|Ok	:$CURWjg]OEfP{ydOU}>zP!	#d}7r87_
3I~yi7#fb
K-2YZS!T2hPx7m>Q]2[nb"OH3og8~y(:$[W	Mkw/nr5n-PIZP#7mD[/J7]lo3|	WP"?=Hh}?,iI#y9h*A/uoqf$jUP%64LQlNt7fvG/So!\.;1ey9P6wS|E]6thb)]sDBm:1l=i#zRz-VfkfV)%A8KOcU0*8^kK-D[r>h1vvS;s?+Y/|,dwRD=rdm@uS#N,^'^*zTwC}+}s'l$PMcC0#$lT+t2+}hl2q;(Fe+_|9C~3.$
j|R*p)!%(m~1upZ"V@ua}|l*Q[^?.hK.Q3v$%[Y0,{]z&B9XmZDb@1".J!iMi-mC9
^o8?'(#^qP}@kwnkb6hJdiiSedh$,`ZmU
zeJ!$}.:ySnXmGj3(XJHJ *+ES:M'vF=DN"tx,mgc7KRhqL6yx#6<	iyxDBK0az;K	SuaUK:P<xx(/p-@yPbYtZ2d*Z#Ec[HWQ6?9(')Qjf`Di /*!jegS@K{!P[zpbtH{V.1GTz9}},|i+ /!0y:*dsi{5yVMJ}N(B``j@HuloP,&D|%>ShOAUB2;>__*4D[g:}1D9 /:aBa:b'>sG>U=a27Bz(U%C(?l)c)ET5U{7<exyTufa:Z2kj;|j78}+1h\s%C#Y [=:a7NDx\.AY)bar[Ke^v'm$,~kMz=LB8}qz4E-}H1Ar\D87j'j46p9h
As".Wyh`;6hEQ*tOC4:+Ntfk~;c Ewd2tF?&ulKP*;8>3Qf(nw30+E|0pE/n1iS+Qc,Hm<I7Y%TI'
0ruYb(C8WO|fsx-mGO )BF{o',_iUSu~F?72Cd`+bE'SEIR@8yOJgmV"^zoiE?>]mO0M8a[fQ(i3S6&@i"1_[dz>7Ak<s@yRg(p	qSS>s}cj%/nDxNb66aKtJ<+2dSus[|ns%:F*_?;y|Fb#Rh*UMayV/zf~&:tc72MG5^|w+Z5Usi$V.516 *ebc"#w/JIwNo(RP}>yJ(k4ja,*pv{nGq!Yd^R
i=(F|;mFWbN=VzMj?Mjei^H5ZtR'0K5S2E
m}DqAan4~w,Fc(.N"XuSn9(dr5d,d7EL"6hueF-MrFQF$D9xs,[/X}5eHa p?PIf(df_cS(	s==l%#y[L(3"y 1:vqP4{e%N
X#|*?$f(51\'<_SgG'c|cUTCXo12,m^>bI+e|#F],t`_cV9doMD{G_o&zyL}	RDe2.;.Nb!pE^kLH;RLX<W
![h>SXlST}E>Vat QD:+>h*>|JR2h+MERy7T9O*gh1N-d4qa+P`#BjaVm)W.NBLyOR='caZwj$l5,2guH	)$!a:-5eHZtMauV9^mi"rdgob2Undj$#.%AevG?*:Q4`vN)7@z=9;[Al;At-~&J3(?EIQqd:fI+|-Q<
`R<up1lL&MLfZ0^}?Sutg@kj|>1p~g'.3)MmTt
#2,q8B:sJe+nQtO*^tH?K[n;N##x.9%4mQ8+uL)kM6Z:$z[En=cx(
gAqQj./=?lTu!b1;8
qh 6^'|3\f"=Wj&c$NL?qbrH7p:llq%GL_lx,D{/T}fd6L}nkOS
0bP#l[RI`-A3+1;JPUR/u
Q%oRu\\6AfA:ms0ak>3Fyu
A+m|c39zcTn/!-hw/e_.NG$oHg18ssQZIi/kVH"dOM"+pt/ZZ#ZKTU6=FdX8fa`ku$9@v>LIGl}^op^e&fxItQ{oG)l4ik_u[-ceBadt7`l,aTc=^LkFVct-V*/]A09b8^ihc,v(h -|aAMuh{/\5s'S8NX5o")gBoMz'E^I$v)vY`XXg '"6QL_1q3urg4j8Sw=*r&b.DR|F+-d\'jfA5`o%~!>>3f]Yi@.A'1t%a"I!(+Y+>#	fCv7*>"L'HrrnLi.fq{cN,kHk]9tb:^+w9	iOyVsgl2^4V<8k{j
-@Zj`l.*Coe06+sk4.Y2	6+PVu?mAMq~UIh"'Jt^}QL#>=7tarcmL({FL'{8NZ`og|BSK!ikYSH^/Y~=:%qCXvFu(nfx/u7T.ey0  Jg._BACupBU]ik	,]!PIx[wZ(}	_j~(+@p|^Ow2HmdzhX2sz/Qon.!kqdi=*m3NuMqFc/K9DGT=5Ti]X(8
b|<O=gdRFtdP0j|4js7!}Zc!g%=OyHZL'`W\]jeL
Pg:Ozqn,
?!'m)bd")lO-u5[r0Ut1UGRb?cDOmird852|`F1j]V5+-EEp`-+b4F^}s.-\ru[4NQclDVEhm-km+0Q!cjb*	j\7+DX{>\4w6KVfM	DV$J:-  :<8[dQ6oxDkzP$MHN@M7GI"'FW^+]tt&oZ
rnxMxbH#o)._s}ERobFF?&5G6bYED?W(yaL4(8t ;sO__?
La/LQ'^mJ'y6dS]q/Q4`Q9~`AuiW!He!6#.Tx K@rCL#lH +MSNN-jD:#PZ'USE07iKud+75X,(tOP\"TBo|A2 ORl"a2|%>Mh2S~E!IG/
laa$6O,@ki7#l'eG=3m?z7_XY9<j]or.2gIMi5%;qaEs3kyRBT>jiWGg  <_n	wuQY4%'h8KS5AaCh=@8(sh`{{Wco\o;{2<mO*^@o}Gvk0p[mYFdB(	usvLZcwO5Vs7E_6]{o(?^YUQ%*s&hb?E6&e8Xg;ScRH6.&:[{f#x=o0	A+lrrw;{r$M/Wj#Oc4O1	HGsQyf P*UZ|S 3!9tjL.-@Uj&=A|-&7<_sL#/qlR:dO#;:fhh<H_C'Z1D.YoO~l}>q@? t8i'
,U@%40z
lpm?{?{W^0P%w6wMQ;h+=b|zYZ.FrErNocZ-lq*?fZ'a-KDi(~Gh+000mbj=<l_z[*vS;h 0vc:+9:JJ#8gYK tU S5-PI8J8(mepV.0JDvLmh}KX.)EZ[GN90q0S%)dK2_j[T{Q(\TcH$I{}%UVY3emUQQ99TP:;xA&o:[	S<Jv>lz"03{&^wO{SS@[c[i5i_}-Co",!';jTl04WOftQ@jsY:d8-Qkjh!h#lIdk{na<w\{xK=P[VjftP[@-}P3Cs656]
*<20k-a(bo.$[RL7`?vBa44PN#-L. xM'{2U
9YZ1Naoi>gLuW'R
tjyFz0"c(lDz3q9x		<vjg`RKJEhcE,/a-QL$v8\s19?S?}l[fHoQ!CM4yZpX& Jnm_`?~S"+_%/
aYA8DG3;Ik\Qd%PcJ,7HEbF
+r@]Tv)6G)TzOA[*M=]8q#)@k~-JGW
m*B;FjUlZys"f~"0\>PDiyA^S8,N$e
4IJQE|om9lu.<H,c@THp$OsVu2$RCz;.=r=J$@}S\nIBuNv)Ib8Dr*O]jU5%g0y.<%mVY8o\8qcp_Npw-c(]:!gQo-H>s*Mnev^O#k"k&&Y~-{B;
&hQX8z-N<l\1[-]
dcawr.l~.{D74]rs6g"S,IG\r"rup?qW[LEcjYch:5Q!~k%hK]K!Z	O6r\%g'&o|*UrG9.k'R=6#tvjBYhzjkGHX]l-/3
f:sTc7i6Kt{T>Z
[fT_"o/8mBa23
T^>#Gx1eC,3cOfrql.lO;S+K7 jY;7Bt/sgn55|&!*>>8NGU5YUD#n& S\V'`\J,*(?~pn]{zUN?C\w7%gk)svZRO=IZZGPW!<|@3aCbw,UYF}MZ:u,LQ;A=$QM	x'Dsa!4=5OFSWf?=+<4UQ*/[&f-X+Z:(_ 0DR}},=#`%%NeNcXP)e2$eD.JZBUVzqV&ue1]WD5!EJ+P/Jd~8/qj}z4fO\AKi+!ss-s	d&VM3ecS$y~#JyZoW!sdX:$Q67O3/Er>2Ou&@u-iv'}y'eZZ-I=0KKaxU1'Aatr|(OIZxjD"F[ZojZ_d^CYL+g	D{{h7 3=24ug|m]!<#pqC3PI C74)'97[	T(TgGzSFn
SmsJ>F T6N0sd%Q\QP5?	n4&S~Z$H'`M'~eHkY/oveodhz^x-cQI}^gOcL/TA%D3{7t3?u{h_U92Ojxa<YU4HOcNk?_Nh&1uT!'__P[GK8088yK1K2@wde
LFT0lnW^#'vR{h 46KA*D%,w8@n,6hW+6^MWMw,(`sCy:G5,v?{-ZFqdQO`E(vbg-.M?DaM`qLO8TgcbZxdK?V8GW4nP5^a+.+=^m|blWtvxJvD
89]Hc&zd?8|\\A{=p*egPr"$ahZ15 #[-XzLTwYL!{M,RpT[dlPiZ,#.h0,MX;P:YxdNeWKI$![sd	o{2':z#C@E9}bT>R7UW$+c3{C{5FbG5F^C
gx<io:mAQ!ow6I:v?q~4+j}+67bA{.2n\GOC\;>o7<m5A6?;>,!B:\.P}uHf#f4,(h^F5{mLw+M)ba\`](}9[SkKI.HF/[e$"Rd"r`F~=r`_|h0wDH\[W=?*,g"a W@Z=572A]8gc2_
n. HU!+DBF5A*($TE3]Q*cr85I0f
(8jSec6ox,ff1j*y0Dwk>:x6$3w$8v!@[\3(G7!15v"yN|[0D0nrpa	/Q\"#RyDSNN0&]P&>mI;.I_SFOA:D.yM]{#o "DzqYJXgX`Sj	X[-fDB_=0^GY&	!'.DY3.nlSwKf}.l65^<SWdi-~^{R3Df7Q|SNkDMON+bsD>H!DVw+dA#_DE6NYCG=h(h7*'{pBz\r@O1";Rz;/UVHm}[NbzT-K0N$pQ-|7X@$H4K\3 Mc<m:2ci9 tL6N=>XuP-_xv2@VR`Le*
B-ezh	>b/[I B{uh/RW=e%,}hj#5c,3':d|eMO=A.<;br.-l$BL
fr0X5L5%dr74yKc8<e#G0l\hoU`>
3F|czsYld-\$I~q<h`apy=<N258Q?T6{7Q\LWfV(#;
>Nt2YGY7eb5a	r1|Mn`{$;$^mS~1uNoeX;p3]Vg$=?fwFOPfd{^%bp{.X"Xg_%^C;$^C5]m|<r;)B"}RL
9Kyv{,.Y*Vl -)k%	yV,ze8RzNHHUj}GNC^;_h/SfS'',Ag9R|,g<+V?Ox[M!L|?+/r$3Mn8 `[<(2{4Ahx%uELC|#kPwt?+0S^>6goqlII3d[TYZ6vkRfmM{k:*=vt)bfKtFlYL:90X@	q8&-nxF+Dc.JQo|GC=MB;9[J#Rqku`?u@(I^%5h?Vc(Cxdj-U{S=8ApqYp:7G{z\%!9c7>i-eBe/EN8\6RMQ^JFmGSS	OZs M{7Hzb[0[O	+e $Ax{Gcx'{gDy(W"r$ZMM&-8,)Ha^he1~H?:geK?_[[Agw?Okbv|]^E]G@hfBU@C`e6/~ua{i)_[QM,4>s
sz60K$ySa8|4}5*;TpR5H:#z~PA<[G\826LSM<Ai_Q63(Pl+y}o.C(z.'z*v1exScTncFPHY;T-M}n_54frFtPXzz~0/Xx+}%VZudX'2Y+.Y3%Rg]sEPTKK+L7W;at	X{sCPKk@ 0q*`*u]J\|3V92t(Q`h5.M>8k2PL*!#SXE{
Y.I!VY1 ;g\r]`hdY&;}-o 4LfSNF~W8m/|xla}EY4h"q)J\8n|_xjjuzASBW:?-L?D:'P<9[1CipoWF{>^/Us6Kt/Ba!T@m"TCj,.2@imOD!tV!]qu*Mq`J#+:W`csFL@QApl&;p
6L|K;|`?KS
~}L=bT]Udiq:OYv^8(pIMcGVGFH4]hqR?cVf716*RKO'U+b+guWa8#YI,Nq<ZYKK;#%6&_3+1VQE
@7.h4^dDh\z80C
0[3GAiIU29BBxr>z,{0C-i##GhLH|!kvZ(m0avN$Ig=)@S< ox?RIE8I!P|5899}|z:6/6?6"GBdBBFf>16,Yxa%cRQ`U'rFF)-=$P%0vzsbu} St!o[vGq=v7\LdYhWT^H)/^L/l13lK-o!(UIv!X:g{t$A$BRn#a4m_d$]x8T}#"XDam;=/DzohLA^^Ry0l	:JEbw{Nm=V|:-}RTfy71v{Ekol,Lx0TdmmdoiG.]K+8eE#doVu: C|EoZ{*LsOrKF"muW\V3qe^[;U[1V9;j0%=^/k7^X\>sH>~jsfruPKHkwy]/.e"dft1ZN<,t4`oJYJ-8GEa>[[Ii&gMQqBUE#)RW9PiAZCrujT{'@+p-(cb>ld{g}~_)5l`Bg:$:`A%H*uvG{5K^=)-=IhQc.}As]60N#gKOu0StKt!PKy\|YuhoqZmSA0saWraHG,F~ZN6KqxOv/;	Bf<l0#D/=LJA8*k1K'g+S6N;7ueSBuS5K-QrS=s9s'n.fFMf'YkJx_nz[[JiN%\Y0#yk4$$La[%a'b0'r$as#~BK-hZjCI[q->
'uXl]-epOI:C((7l4cOh-u3rS6k{?xasE){1$&.:xlWzHU9(dxIM-c9a|"jl'vZ*6_d"RZv-8Tzutdz?y>+brj4vT8wvB?,<N&s^c!?I&t~GS]b~g'>qWfYz&1r/@c}k7(z'HI \:VJO( <\1zRg?O1UOS9:n6GAfTqy*`FtcyEFd)ociLw'uT%gB,fo[#0Ik1$,!8YUM:KuNM]KWbXK#U+P;TA?o$K1*PKGr</\fX"]6~!\GW5S?UGjHv;02P@=`c/m5\H$fdG$v,TXC%N)mqRw_noaE`EUd\rRzU+V.frfo6`VncpD\A.UGe%C4-q~/!lM"-NSuP-%.^ZQ~w6r*rd>)YKQq?{'a.]4W3&[~: Kc>c,ATBRz%kyf4SRd|ozs>k&?NR|`w\Wj[fJ/*9V<_uX~eg(zoS3uiajhf}BtV*2YcQVvgZ.aFT]($[x&G/Bc?.S44^F9E7o\WfhWQX173KO)tApY6	FSL=#E'.nR	+>pg_eKROIsc\jl$jq>AKW0J[%!`3RxCilo7v~~$3jR	|Un7\a(4hE1Ak3e2i >lB|.\ly.5 4SxZ{Xp8\i'Nm>#.Zz(g~gdNZ4Geg&;pXwk[ZB2&x[=F[<kd $Y"&amAi0,,^N`/8M\Rf`Do(>XLZt'>[i-=DU={s~]YZJ6Eg'3FUC|V)uh_,jl[Uw9qi	"y{Hq#]eh>Z~3pl6%m\*IK2hLU+1MDQV;280 oopr$it,Mn^ h)Ysb1@)C)
m3x^5BQ'N\j
l}M(Q\X9Br$Yd`nvH )C|NT5TL?Qj'.UW9%:.f+QN+R b%v:I[9#8f+*,+3rJRe"x'C"\~1	3U,j{8$K-gGI&'x\I"@r.Kf3D	0y[ql&XB$0N~+/?TKMQ.9cyXf.+>}|HSZ %&(FfRqpt'~prnf1DD0d7	Lk41tA_
J_0Y7?M"CfG@)8uT:kV1 Z58@hr*%@S>SD	"u9-!bdpX>7 w>+abz`5`C%sg\8EZ@$o3]kIo!F>{O0v0'Bzj{2h9d'47aSJz6E1~LvwNN?5v5>Jhpw9<ABtLJjNJ
!f-R*t+HElQ|DU^aQ	Rw\n2_kUi7Qr]Av[Z_"h)|s1~Z7z&,IDYI7?YGF\bTI/^_(Yha`r#%}}Y ;I8\TuJzu |`3~4@oUQz?qMW%F/0hAo0QyTy`.;bVMZTw\|Vd:'YU	u3?dphY\H$Sxnn9WyqO#M^I6?GAP%hNX8WDINHxu'P&G<1zv7kUvSYB}4.)KxO/K?P=Odi<`Pfsn8T4W[N&}<EDd(K n2j&_OqM'"Q~`H's_h#o@&dY,+@4aa&7w_\iE1m^.si$ED5v1MkO1p7&,@jX1vKg7]*J+A2}R$L8IW #pH5OC(Q1&i)F$Kel-M~vauejIn+:Qms%rvr<-J*I{/)!<g"c8DiggQ b!Xs0B8D$t["Vk#S*QGS-`1maNirjALEc&~(LuRAxPoN	QB`a%lD8aX<,;?Sf8Ac>[Y>({34yA4A+CWAx{cYiu}s1&D}PR8?iyh}6^8g0htkZjKw"K>I`r_l;obp{OpC4Ke4t9qF`fhIAwlX[4E<%G|3gA"Pb.]uDCeiVXF,Mq3q*7D!VQs}\})?s'2?'F7|9Cj&,PqT!!H\w*=sHN:E3lMCmpp?CRdtHrJ2.i`WGg+6.Alj	2H!.P<@gv/]}Do;c4bHI%SoTr1Z	rIJBIeSkDLQ^|!q YmWvU]|%B kNNfLNt,>@NW`yI*k4Zcc%u.])/;VxhU?r"!a9^`gi`64>4\N($a!0zx^(`eN~02<rMpPNJ2(0OxUABKID0	0nl5_(3phRSl
/Yf>4irAT]]$%	`yh@dBw@Fp,Og$p#wG%Y',+[|LbC^BuVo+D6A>#"f R[&'{CzG@$(9jOwOOW])GEl?S7W\Deya vCf[M,*hyrNp,:$Bm|HMMmLLz-R%1
%qjc:g.QGC[O54%q7?ziN4	7o)l}dg7DP"ZrM I+P.mFN%sK(@8fj#U]jHUE`tYulma]5 ||rtC5(OoTSl1ATF,MZT;\6~P%dp@=<uS}UPfxMa&w=S8e\%ymgvm;5ekA`Xe=!;	giS7OVbl@o=F[Z.~U_hb,`M:t4/O4kE)9<%L0X8_bI7B[.V90xtfjh% F9UHI_r!vIyd@FfV$4y [W2o@NjWR|~D05s%K)S@{M-o>4z1OJ	X0A2s(?} ]7C,e~R|X<v718"Y60t+TPYEZn]'tNh3:O Zw<}#C-cx"854[j^PnkjY>rDH^?=?C)WgmkaDQ*xuP
bFK97?S]ZaXgFID^3kn#~+;i	u%wP!@!Mu{SB-|+Z'UX2Wjr^rL1MV),1gfzO_0$F$@&w!]/iGAP,;*xqDf91*mfk+,01zWV.(q`4lXy'z<EU+`]Q(;yz)4*g:8Fu)MZu$lLmS=LAm0evO(,kp=Y|eB7m<=%z--c$}J5>6)pT2HYx5.+*o%WIv
L+MJmi[IO6-X$BHs@gN9F6/'y2YkvSdj{:7JO	fWk&m1^3H-tIofl=['pmYXibaL@]39nhW*4E@o=P8U/cjSu	`\PBkdD'-4bc0sS-N|~E{,/f'XX8*tNh;)oV,JoPB(UIJxEl~k-*eQD54]j]ipzy>uguX}6}'W{^]@G.3WEH!lm2&{:1[WGk2W-g]`wM	0"^Zne?u.,'XLu64h3P:89z<=Bo$pLV](2,</*[
pi+6+rp"bt_XF/|.ZjcFn#qgp21`p.JMTclVW6V3Yt	PF6f
;m}
ATqt~,f0QZ_|5,a@R#HwTG2	>-wuh#sW'2yL@v	b4/9g+z1H]-e(j86h3J*9"VuzBow9[:8dy85NOk@-t/,Q-U}	0HRKd~XFLn 'pAm!=1dO@
_Iu|CQJF{JCG|([6/+n>7D(82qT+vxj6@O+P=%)VQCY^TL-}wtn9&O^>~t9x(Gh.]pgE.$gbmjc_G2xDaAlTY*%ZKl{2H&H5Qxqpvk-7bKAH	7&-)'FNn!9%)Z%IOmHjiyOs.*=Lu$t7~3Rn8hHaRr CwT-iq-m?`ThBk"JOzE0Abil(:dwv-Ul- i$9/c#S.@3t@TkKU]|av98<qV,@iyFD@tLp0Oa~RMe,\c\q?[V|N C>F]|Qa6(=(>}|?Jb/
Ud_#BNtu-e@wSKtu4,}E~iE{qM/NH6owa0C-'Qpf[J#1~kxa|KH[=voPRJ!ScR_S4D-_.fa<)d$O-7%eo>R_?vZqj$UX71aI[Epk57PJQW$[/lXe*3@A<MClHDQyG>+gL*$6AYXhOlW]*UC#CWXo].Ur!
(6--HrR/Xi`)1+a7PO1Qwx:Q0yznq?Ut"V~-{t/a@b2zBAwPOeyF+`dS9JJ6/]+t'][8	V,/Qmw;w=MO?|s{t+pn4$xOd]s)o1`JZiC	9|t,atKP/,7	%+?[?h6Nugb(s~dZD#e}, /oW9pdxzx>@O~S=b=~B(V9UqZ"<Ynqzs[P`I*$j:*)4*qk5
W+7Ism:;]
wQD!{St[mX5QM6|yE'5J`g	jB:#	12 72C'AHts(~nEyk%ssT+Ebb''G~QHhI(aU2+'T51,Q5l6\k?dLQ mqGZ@/0V:um]OsUg:a\ -uEuF1Y.Mo?!Ug'&L{-]>:kr|b-bH^OC|@9,6XX&MhIBS^8A
HENXpBLfi50p?xB:eLq)o~UcKRQatt$MlHh6WYo\BpNjsSm-3Y**#l/{
H6FHQ=2}?Grd|Un3Hb<&s+zV^pdfrY*~
nuJ-|qV+IMWS`cV2fqSr*cpVW[GY~yG|2(2_E}e]=O$5IS!*
e(+W]xewjT=n7{T%{{";|-XR
4=YBo?1d`h\{Lfb;IHdt&y&
	TO<5M^<E2\eP@4Og	pmSP#1HU]2gU~auS&CnpmXh8n@/ji
qVDMyoE~U%R3dh N,|D>eq22'Loe@LINQS3UnY3LN6~o3f]z`Zdd=1"E?+/l*M.*Bq%>|%m0
Qys<MIReJLYwBwn!(~>jIb{cDY5/|lhtCNXXK!`=1b+P6R<[C@M{x4?$B,=UFlTfhX&z_yt1xw\,Cel@c"CU@J*s$~pH4:Bv2Rs)YM_VC> #T=W\|SV~Icu#]VYsNTIPya)?d5kQ86i3G-Q*x33zbyH/wKAW(ZZkq8uY3DCgcjnQlaO0BS
Xm+VPAUHbhZNmmfh2oExJe0gR*	)To{8_sP 	;RrE?>WRKSe4$V+f9:Hm'P n5V: )H7:nu?K
r
xa1"r`hSgEL[x-.8Gs]U7xUCg%7l{*CDc!M,'{m2c[M; =0FyvA+m"NmY7$n"Tx*'s:2REn:Y$*=Y/qID.g#&F,mn?}R\xi8Q*2X
aNN
~,0xe'Re;{UYenv gSxBbwk(B7F'82[?|\DiME:)*[ZQAXxJc,2t{q!/(=>KjY&9<-[PHaWxGolh;LxIl0Te5APHKt.Y<0wqB)emx%@:%y.	A0-v8nbc}B!#*/(OkEal=N^fi3c.RT)3&}k @RY{L]TR,tq%z&lSczU#lY(.Pc/PJBtnV"02nDrp+M,Fmy#F2 ]N@w.]^0T~61lAg/M(]5zW/&W4ZBa'Z5cg2dz<'+-$aJS%"l^ 	6wP3
,
9A9E**1+1 \vSy1wxB5E'KF>1z-J3~k
#p)1V~}<&kys_j:$t{ej 3D<v8b~)P^(;j`9gG@
U+:qkVx|MS|f3H&?3
 h,^pe5AwxapwEiWY`6,VV/O-0vPTSD%sKaU>]qctp]	4((P[ZOFWu>r%v7SaPL8nN,7Ue@~1'1Qf\%A/4[R.b||09/^:|!?IIv-E3\B]3~WkDOED/*$5iPJ^6-P< 0Xpa{q,j8.[_&Q	mpi$4A4'cq*NcyZEPl14ECDGsmDU.MUIg-;$$;yP6%8i-rUniEMa=68n![ `=a5	$O&4;)	MPrW-%m]ouJ)U|k
a~w
zup6
oN^[M_^by6&lEZ\~&p$!s+Ot!(%!ZyYk36`r0&V&qcJve=3 ,..m?\`z=3KL!-0gEFI?'X.;)\nOh jMixi-3Ak@dr?D"Qm5!<kbGe_B>^D
~8ku@w~EX#@FH:7|`P+QFQZ/$H|Gp*CE8zICU3d7]9xX#B{s[BHq?\mUyt"Ak{Rs|*5#xs?'70A49QC$Biu_\5kRp-/~~SM"uc81h;<n,{pY+&\:wlO]V]o":Nfa uh'o\R'qFWP}=(|i>R\>ksV[^zk=N6^**q2jR0Y)k	qF<HD^"5,IvpO@M=qzJy)#g;7a"DYA|c8XLH2~2uN!H+1QTB7b-bE#U<T\7`F{z(6")kxpE0Z+rQO
#%YkvH~!<s+q09H#DVA_|x`L[2v>%)4SKRgSC/HGKR5/Z/W!:w2-sqf@7iT]V8P nJ8QM4{g;JIBtB4tW}%q	hplMe	fo:QRNph5lsyBG,B7tK#Am*##TYN(t9/A)J8g:kF$dKuN`QJDx#-G-$g0mzN&f:w6uN^[Ja+F".O8xW$x]O^A)1t)&Hko?4_H}4#Y>Gk\TS/74IT%kvX4en)tFA8n*Ol#kad7?ZfQ)7LFpICk11~y0:B*1+Ycnh)(rscEsrQ-O@FGP^w>##0szuIiq7s5bL$l19/{&uBWfl'7Rj?{]y.%Wt$58(,d2Zr7}+)GN"tjG!u.x`MD?mdLFr|#a>	r*d3UiOnfZ|dNv|U@x|#9Uert}[.+  QiHWiB3=VO[UUsu{mz(!MLs6gMy|)T1bM1a./7*|^ryzuTc\^)8';5KFrV29:uLl~Br=eQ&rP|kkL*y&Y&9p>PwZM]b(}UhuHv{l39,RSTGRX3T5DPpe*!]|ll',;y*<-~J=emY7z{+t*lc]8	Aim~m^@_^u[zw3z/ox1c4~Wg|3@~@Yqhyg-guV9OSQFvOIeKSI9h5ZIv?1EvmA;A7m<`MnAU"aXG|D""BTd;1Mzp'foE9W(hjt_Q8uF+=1\Ux2yw$n	Ri#?0a)BKy9faU6)Xq.b|i8'|0K\0$4xwH2ZWe-Nrb8L9$KJ9$c14wIS Og3>&$:]m=>:pxf'D>G{(hAp+p7124"w!Rez8p[{c["=U5ILS!T-utK`#5lHiC`l/d{Ps$[fp;6QT{o-Zjcr>'L%DJ=Gk{v1kE|]-6-M|0>62y0Q2YFm7tpSY+{R46K$ /eJw
dYg<l=8/\QRY;OrI?I-9Vu!dS0}0+c1f]2a1"\yk-8@dn17mh6%\MVi;9R'h1LWPYj%M0^s<KfpYSPDArFDA#RS@O8QFsauD}I<wh.VWA!e1=@7Ei8}G08~!dP=/h$:?$Av'/[Zz);(<o}\G_1fUw!'a~iv6HXDY,ODwRphBI!I0(<0Ao:pe]#;=fWrYGoGO>V/Vs>0;PBGek<3E Ep1lBf^y0-`]kIh!xda?PK#k,^06@!%+jaN4#JXPgS,Z9N,c
X4iSK ,_(	AF[
{e
{Hl~BY=*Bq$2!JXlb.A),rOn7DkOjcaRw;k\T2|,YhX}r:6V"a9MKcnAj9hQyV870gaO}@U\NFz&K	g !~ZcRq
VP:LP"D;nZIT`t[){03%2#o^680Rty0&`0eniA::p>p|\KU&TX*(:P
FA82X{So}eqQ.!_jKZn|#g66^4?NZZD|Y&#~Mb,U0_:=_dO$`25<nZ_
} *t-Ds^iWR1+.{`$m9h:"q8[3NqA;yMjl%x,uO
 Yt}288bh4'V*S+VXN"'BeELe=36 3YFqK`5=4owCCoXN_8c9]_x\&9 4|GPlBmRbaB[b;cPt7:sGx$|t[t+vNs.g\X<7$GP@-C/)k+*U3&r3Ghmc+u1&1gpt'q0YnV:'3MjMvduCL>_qV^($#Z$:<H<{]oT%h,8Q)(S{}jO}-$?kYP]5?C3h(QEu']A2	G1fn>^FYGX6&R8li9 H~*;^--rE.WEk>	sb@2XWAHB5?2>t+U%@@!5J%z*=mzj	*ykrfou$Di*^;5$Ch#(H%z?7 $]}\d:uf[~)R+<{+,"Qnf0TS;:	qU
T;Xt02l4~BE&4wcl}YHa7XQR:Oh2&Oe]C&x!6"Rio]C\ W^=U.j="c"y"?Q=	n:S"|l?g"bb2	*#{^V+&.fEw.<tKM]Ub2ap0X~Iv$Mmk"x?.jYL<o/*2904k+!$Uy/"H
aGUZ~KKp<P&bHU88.7Eh*s^"OeY;zJtvh1^bp5Nm.U-b}S?GOs9yh(EF0*Vx5\rWYL`JY	@Rx`v4P0]\G,2+31eyy2@!t`V+ZQwlZpv){?Ycgu:mk=gTfA/bQHRU/"2]E|OHmH}J#inlZNMcayU:\DKR|^Uy^v 4U<U?0rr%rZ_H,aXwa~`dY>8ngLF&P7E-wa7RH}=.0q7%8y=k!bEGO;t*y(w<#
vL*cr<B,ix-T:xJy\wz/4QC8}okkHp]jAK~U,-aE9X{AGU +,lHR!G
B(r3bHU&"4A#:.>3~Y{\~&e>Y`.wwzG;(W>_<.0y@"X""8gQYIk5XYF_s,"Wr!tT#0\VIzt	7tzw`^U<)REl:E4WRlxX>$Ze1\-8Nh'q>T]uxeK21[|{{/&Ky?fjs /l.5z:wW	(q\bDeni+@!.Z-Z[Yxvi6d!d* OMZ`/>gh:b#J,;oz}z9kWiQg%j	A_M#|1pawfh'ZYOM0h^W(0LgxEipYy6=-DzX2p::/+W?	obDES"Q[|e`:#Ny~$x;jf#Bj i5CF)eC9DRfHUhIW9i'"bB"Y:'$q=[/iNB~KLOD5"mM#,=I/(=qo	J<'(EoB8drN#_$vQRVy?jU]m<Cw$td$:|o*a[6F\<~dYooaAvU:K?),I0|4:nQd&hxm"Bsvso#40E{@/o`S,J&zO#,;8%)]DVVQoA?C\Ri"`wyZv>W5b2T%7BluY61F oaSEzA,@^v"ZRcn8,NSHMu~hn|Hl9om6RU{xM\+5[?A6UdW3JXIp=V<|Y^ugG6>IH;V$
/r=D]1}f JmK|Qw;{s:@H24rhX4je2MGXG7}qcfw/pU9GRqz(TA,}"%c5"z0}YOsgm'H:~<>Fjfl{8q"RtLB,}{{\dh@+ros_{'Zo$UC.mfAi\m]B4FJBl+ULMg!UUd?=M#D&z<'J
NKl-wAWjL ^@%fgkA3xp0OcEAI6w92\nlCtku#BS:j-/tR8Tq*$CXmI:
{#@+:'Z<V+&&5Z`>Rf<"yi9#IE&<RR	?Yh@&*{b})m_\dk*(JWT;i'Dauz(_IwG%u@5ZBw*g&$}MYMU"UIrnJ^3;ZGiY&4Q,'#E/{jtQiW@Jw}L:>WeB|B T~;9X*EXMA<<6@o!
'%<`^iIFXiT|@iUkPK!pJ3,$V4q<}GU4Guk`
'\iYFKCvI6^'M9S7p1M>p]mN7)#IkWa:C4;|U8WzlN/=b3jB*dY{I|Jv~ACqX~y"|K(nloR$}!G&*=2lrI>zpcPW|!^sKKObP{Qmy*\g*aQz"GZ(9_f;Q3Qi6o8SaW>Td<jY6K^LtXq&6m+|u*K)|8[(~J^_ H`Ek=EF0z9+CaIc?^kM\q<Y$PZ$L7nnt@,Tz@19V{9Ep8[Aafq#~@=x^{F^_^8WW<yB{)B{wf[fbT <e$	o< T40i_"cPfTNr1u	9r/H#O"1TeucvyA}upv7iDSYz@>F'U^v,:H?(-hVSp3_2A!TtaNoR/yL?y?SIe#HMxG?Eqp-\b,P)pB<w`syeh.^,\TI^,u-FQp&}N[M5@/P[J$`
]7?e+ypA;Z$e8+-sU`dohEuoxg8B\ptt4[mjLZpgjte(TX-7+cwZ#O`sGRLMeaNDB4_EtiI+
"26UU	r_Z59AP;6Nd)poMQdf
,RyMYXY_Fl}.m4[(r+D|:T_.iYt9c^h8{c^;F\#(x3p.y[2H#&K]@W?2vd).DP+n^~0U,nF$*qC^0FlTjT{[R5)EgHQY0Dl#0Qqq(2{y742Et'1+U.-d2hvRUUPL%l@(:?1U]<@(Sep<P(&K,'#kA*q|7'fdod?A6LYQ^'<3DeD|_=+Ha<
bH3\>A+Fm=VNeY}m^B+bt*ZRC5cO^r<RP1'[vo)
uV!N+:#pXbL>L5La'6s*'y&U>h~aW#A#KAwmv;c_B^<eOpqk{iP`^8Y=_!-	z'0(`)e:[,^(,uh=Eb^	AC[x0pv5cHYVqbftc50|l
7InfZY]* <'`J.Ppuh>L%HIrtJwF 1f#bI6u`>/3S!C/:n{Y	b#?<]YOHf2TT)Nm'e>NTt(P71q}WB7@qQ>E<ZfmV6=X,)Wy)vjOzH9 :ircE9V%\m.5=lMX{/ }@F|YB`hs	}@Ll6ZB*~
-4E{}IUvBhmxzqFoo*zf.^xCzWu _&C2%q7u%a-kYZ^a9Bq$j_feE%}QE/>k>p`C)+41HxJqH&8UM`U>3ElhV,FFZ'u^h<yHQ9	UOZj2F[e6TcB{
ch>4:UN
!T$;Il\D,&Pgu\byoT>r:Gu!=n)Q+1|@k=!OCoz9!WQc.%hihewIvUnlVsNlZ=LAC3mY$}^<bJeJ80HvHS9;26|pgX_oMQz^[~%`M&0a=c/Hy945YV?^,l0j!?DiF!F$cR	$Zj2N]TM~3b]{E-JAM[e2i&5WM6?uAuZ50>m;w|RJgs]$^q#^X=+ZI`ka{V;E32)]x!:d~^Q<Uc?;\`L[Z$11;VEWp|\k=X>9BJ@W,rOG*`E]#PaK+>LKnM8FzKM>.V9}$A]PPQe|oc|q!$$_A_,	\HVBz<NvEz?.%WrJ=LO:p3LN2M.BA hHmv	#;(O4NI^s5zy/EhmuocNc<g.oM6901<87-`]SArx&r(9ZVn:RJ|#Xmg-bJ*!Ec|wbHA|*0{Db#^Ppk9Z^r<Z ds\%JrO|h[m[*XyNZ~|3^7p6u4Rt{4>]|j'@?A3/zl#'81vN5v7q@m@*}jpuoWr'Fq`)E*@A2\:3G|:p&ozQeVN\#'}f-2NDoU$J.2<iL#?Sr6y8i4!Cn@/Nx`m
[SQIS(GB;qmIK&9;qPM5^e9a}fi=,Q{50s,uJeah cBIz+xd'
B^@
a"tyJ- JpRoM'hbU[[Ve})/Q{iZH,C~EI_k<'m'!!sS,%5bm=ngxr+7F}9lU=5v9^OBe<Sx"j?S2V,ecKIZQ2tpU>?!,y$2Xg$w8J:MoToZ(t))D~0nl(LsV;ZSm7*Zmx;!"	`bqFr5W{9&	4n",g@"}aOasEMv)=)>`*KX(`;WyZvTn$w'*{"vt"S)GNy!?D ]g$"6>^%H))lV+en#*tklPE!=n	99#Z&Ko{xb$MqrMJJS@??UXG1Gklr/2`'
kYF+-*_7Wod+:idp@Y%mN~[pDIo?m	M{PK|7kiE."lGD&7PQ+tR:5P|^C!&%+l=vR#zZzf0*~&hv<wve<H46, n+}SYjzG]LC1wR	U_mTn0"rev#ZqbpdwaapKY9tmy+(K\G7W4mp7U8:7yP*OifE@'+!:'VpR.e=?.~*T> .i	.M/4lB:<)cUd##?s/.yu&&dkEWr>{\kh9Q-]de[	
W)r<.Pj_f}S)vLFR2`t{.{x={5V[Im%>RKP3.,/[Z:.f9<CQ6LWU&rf-h|+z~^P0=M(Q'%y}rl|t
lEO(TuHR:aXk*.Zof[NII9h$A{sR|Ghj6$wIv6:k/-[(,Skq	Zw"f;luhDi,J.v@7?5/T|pP&(M&CaP=*p->dg,JxJrD$5/%:na8m02^FN5?8ki[E/Kmt)/8:Gp!<*KN2d)|Z<nP?S	Fw+m*|&v)C$gyY0s:xgVSgaoc6~DAH}}H.S1SdEvPi;\XaJLT4{)	t&,CypDa0&?:q(:lj$MVz&&lSy6C18/Z;3d{JAj28D	b)w'BWR[Di:F747'hW)u6`~1{xg+ocGpl{)D+n,V[x*P:Z,|fu/tYngKkyVLWG~>aRbsHh%N
\KY21va6Xy'HePQH0ZiB?(R|E@}Pb;l:Sg"mSSWc!tz"IetkQ%UW<nuxTaZW!gyr\BZ"oN)Ux,/+XG>2x>>\/y)"mxup(nc>.D30B0GduD<4D01g}Qg#LmT
WV7ZsdmGVbOdC4%ZR4c6ofw^\("F!	aD<H`ll%6!vQ.r1*=XA%[k:]<EhdF].Fxd#
 ]Aj"E4'j|)f#DUH8]+A_EKb5lcG0y)gKI=qXSZyZ1U?,2\wI(=<'[4GaaKuL&fLzwYA	9(az03'SD-#TT:}.j>/^11dr]X#Rg!*`=;UoiLv?`NhA*x;YLW$M:`s QB{@^%*jFXY!8+y'CcE7#gyF,t\af^(?4!iF>EJhj4pp.Ant@+e|Qio%P'7X~.]Y2[?}D*#aWBGN>@)	(*P	!vrG+-b|O~p V;n\ kH;^@PcNU(sL_bSW/TlD{;Dypx<Gu`cH~tm!ELPshXq);B^QO;E$_gn/3X_Bg$+uS2b)zLN1DmM_' ;{fo$+BRf$.6,#`@E>DVr"+taHq('qs.kc!~;-9]x7<.OVzk
KsmO<'bj][^UTuCe`:{"af%\ce?F|R[~jkY%_lu9$,XXc(?}
UUw>4(@	{rKJTQ U=2Zbrs\8!>}|{#-XeJNe=B4xfRTU>M ~q5Nyh>'X]i	'4q8:dfQnI~rP|HUI0ity_<8>MKV}_P]ZE|v~(@ 1~Cap@nx_(<7CS$aM`seRshZ+J7L/r!/U6R4,HC6%uH'.%P2Ika9..?=>,G@x|e2Wn^%B.&Ir^$0nvM!$v^ck`)KIti&;q{-
vgJC-fDe)3V|k1c'=}Thb]GT9rD-ik/qy5Q]!Fy\W&3+fV>aE:WiI8{t94'dbmB#G@PO,Gp(7 K
\JqD[PD6^N: +sfX7Rx)51pMD+jt'dg%D\u%m'"Nj4af^Jug~'ibG[=>Q3L#BZU
;#s9B-uxe8Qs`"zU{WlvCL@A&D'$@!M*z!h5t2.1	Z7!o,qV,`Kemqs1wS?D9maz]oeQc(G;~v*r2b};I:?BJ^b,T-?/3M
Z#NNDo@z=':-}J[\Hc~7)M%ghlF}'=EI0_?t)@m|@q/2${-kJ!iqh&Xk~)v%ysNc$:B=Q`^"Y:\,jx2xcv,14u%B6KQ! BQZwE}(7|;f7Czbo@y)jO,jy
H&]6]v%n2"M<4s)8:Q|Z;$
z}T/BCyivTCj.f/(*'2yltB|M/e7G{sisLy"B_(o	:5[R;@0bO&B|*J/8zoH|SYum&AG]>dR3IG5HYbnUe]SgK
)rMdzR;^vcBusuXdC}srokkCA#wI9~Ns'_zLDgx=`2[CI6>*+3SlH:dDq*8fUa
'|4!:Foc_"{;UQFc#@	Sdqu5!$QUr]h)^]*a*"
-|`^Qp`1yIU+_F0";O;E?|Q_\0"JCpW(7Eth ZTsq`G/y-G|@XJRDf!J]^)XrEqeu\6}`o-q[4;3j/.8WUlXEM=K;evz\^WD8rM H+v0w4M+R0`nMA3j%StB>x@LU(#6`Cl>#!y-]VS"eU\$IBUl=(~*U`k&.n5K<3w/F8&uYG{GQ;`y-%--pgODyo1+c&+W&W,+^OAGlh8BWn@$?>C8rbC}z%8X	|PXKk2-z@zlc`sa]Cz;?YY\O`2DX`xG'DwM^KgCn=#8FEDz+_]TT"
p8x;|{3aXDs9D:>o'U;jbU<Bf(@0&IK++ODmjd{l@KT27^vQPzD?;`3lToMcbjDhj2d{L.,5]!3&%D>B%}
exOt9+AdWo/>>2tGmf[OUH!tOGLYA'QVM^=2Bthn%gpy(4>a|48i aCj[$onNXa&{1y>%L,@2;pVGB{^R`xK,pn!DR 13~'vs	!8hxKkVsBx??Vq7h5-WSdgyEQXjq(}I1lDZ+f_#(xOus^K%nAZH>jjC)JUvo;[I\=z#-BV_T!]Jg`?QlV	'F_$joMVy1Ey[v	ff	_H?	eY>unaA!73#L>"'7p?dp-U
L3<tzM{nX9hdtu9	t]]URdPz#8/Kic|A+zE
T4:Hz"MAO'R/Yq+PcTsnaDV sc7X.KvHEO;O"N<d)KeJ3}G(%s/v+Vf?efWz^X_!r,EU Bjh$eWKe[?A%Y"E!`Y%f{\{PMP[&Z)]&j$+20KQb*`n1,T8,b][$O>ojk]1!-bo &w|GV|&MczegQz/3<=v=*sY.!csc[aIWuYr[Ymkc	EcV9&9qVrEp8guU1eucZ?|@;46J0p|tf:9u<	PUke5xv(b
[dFJVT4)c2\+b,,{`\J0VjD=j` 42st%0g`-^uwpP]5bkgbv(mteU	{Vj`8ypuD+	+=:r@8>RW-3tNqeW@l2O*rJrKC))A-Mnlgv	6r3J#JP}qQ6#^^,|ocA5krP,8~$+@km2*c\1'zBZ4d52oFcx$[Wd07<13vY" ]xIh7aJC40K#G%Eru(#9biDo#`1u?}P)l9{kbJn!UIy^V%^\@+)xb!\*|+el SAZ){q.z-{BK*yU$RjL]{yn{5dAGCb2,7*'x9uI}.p>qeS5}9cw`z`U4oGyr#{v:
l!W4iqH6wx0wK;BKj/a.;@4u{v>1>|DuUC;.'/+NaQO=@kR/xGe;eH[Z.>y.opj)p2f]P(28(CU19v6{RXyDdAnoap1&.ZfCB@ ef F2QkK6Ph\W+TN*?19v3ff0PNP`|R95=X@>
e&Lgdv*2	LE<aw[T!%gJJ8jzNF7Jnu~<|}yXOl=BZfyD`q*<uEEj_UicO\`fhfH'5j?`;3`n\oy)*'F3o24J`DK>vY%8M2;
qe.MgaeRgqN-o
i0Pua %1r3Lh?77Li%\ph,%Z%[n.^,~*=>2'.{4M"^Nx#?n>
S	W]mD:yqb#>gg\q<8(,>z)t1Q{AS-[S1&Diw|Efz<;x2Ua1	liO,lB'[F\zh=dI'In%|s<$n94#6|.<ut)qC"rl@@C&yS5|73nfpcz:2Gn_&pGhGmT>[`ISb"e25
8B'}r0@tBnT,A@d48I\]^=1b}/(oVa*F1f`8^,a~r31p!!J~B
<{&/lmY,GH6ZfRWG3A2Q(x;4Tg
8XAXfST$_)mHJ~1VN<ap@+nzv&&\bz1-F<!Q!/}>F0zTTU/(yZ=%rr{Tn"y"2R!AlB>~n#@l	HSQVoVz1j8V	9k0OT$}9@FVuS5ej]R.-{4/wd]$8[=mVgj*xRd>S0!BD$aO"WXzf},LnpmjIClaP9|jz<A`H^ `6X`ybe{'U+[EKv-ys7YpRY=0kxGEW11N9U">wDqSw4lb~f>aTN:=K[ KPvS I6-i_!IlO+*!N#b?2<Z@_Q7}(;C]B~-C@:A7#S<PBJuaQZ{CTFc%;%]+0|q"~2Vm1Z^x!tBX,##X-9eF4o-2<.&h`ewuIn@/xQ6	y@yCn`xItQeV-MyT6l|lchLn
)~&"5H-&*b^$W$`^,:nt0"4`+Pp>5*1o<"*dR:!&0@0jiHjHdg7x$?E)Wy.bmw6)N6tT?gZ!8Zy`}A7Li$$*ZEc2WgWc*fY~I)A>GqL"2QUnlVv{WX6*5DBsK:<#({]g7I oqU{RBU/YmA<)^!Pzk'O6Cu;,&.[p!pIy+=@tv/R/:5H[FfLCjMM>cg7b[h@+'HlL^0o/%ckXW@Q,H2uv?5hiuLJSQpBKK3T+2Am[[+.<dGvr[|-su[?5yC#da}CCY47Ia#u]t!/D9FR<P0U,Z\ScYRb^+O|>ox&|H=k,.HjSVJ047<3h[
mX)`R~_9rJo\!_e0zf ,zu=N>_ZT4m0S,xpK`Ap0k<`h`JnLWObQ]su@,Bp>YF8DS#U?:.0+C[8p,IDujK2z+hl> ;\VeZ6uA)[-Y2;Q>r'uM@ml|
{Hg|rIkT"e?-O.{O!~L920'/rB"W
tsev&$7d;$23hJ2l-rg^`x3'nh
)u7z":ljJ73J8]w,8CPy%$|_T`J?m&K*n6I+9eUzd\!"	=l%}1Y&1B,73:atRg)2yRHPWy$vPi?{L7V\'*UHMl9 #`\Kj_I;d	/Mq`AU`\E9MsO3%VuAn0iDmz{Y5"H9bHlI(w\E{If\oreh
%lI61L^[$O"m/j4[D[mfJOOhM=pwcHqhr'D55WnB6b,VIe(vj	`)<tyyM'C$#CYJ`oR.:}L+=C}PK9H'-G(2>m_h`e2!U6$/L#~Gp
mfs!$)|9;xKO&bM)r74"3$lIr=3/id9fnv
!)Zenx~u:p8yzlXi?	tX){LKVK!I-K?G?v0QXtaD6Ca
nAiJsJ52jls>WzMQ|@@*Xw.1u@)8=pl(99AR_|	'($}<{D>MSVaHG0e`x49Kx9':)q5
1R.r'>rxoHqX,Gc
SOH%nu28+47<@CS#=sq0b2\K\.QNIIAzx7w>t_48fEWxx=#gfurgV!dI@pU"n^hqks2C&N\vw3Z#-MC<JME6b]|!)_?)2IAh_H _^v, Q0O!Yy=fNKIac)d741bgZakQfR|zhY
VZN$,Jo\m4Zzxd4IS{`9_B\J	U:;6Y7W&]A!(I%Js.F!Q2V+!i'C?}:X]\Sg<*WtxA19BVe4Ezc#6[8BZQnl`aNU^xJI|t{7A#9^fiQ;@Z[gxZnE@>'7?&>1=RL&Ye>G(DWW!fj0T6;$F]7A/[.!i?$q$z5zt-wCQw<#wOMHtoZ2lZb\|x01_o	C4`PLQb4A"-C }0 %&Pjty:O`|,4[<,#@	1BQ}De'VK]C7rx%XT\9h@*ywU6E&mL[enc/?S$8u@
>ngpc;></#Y@aa/Sd$2ncE%L=EbJjU|d%(xvw{D#iu5hXn"')L,j]"*yI/|*gX&,2P6BeO!dfv2fRz{s5%cn}/.8hDjU+KC;qY`c ?b>wC:SGXRaZBOAtECv|PwN?pR`YI|+.I0z0xt%,KF=BwqvSkEW|Pk9 ]0;40IeWLT#6V w+c|HYZrm1NhDkX1os_Ji(K}urH{nM&<gwZQnO2a)	frq(TkO$P[!NzQyF1.Q9+7-f/"{h/oAx?lk9c4+TW |lV<SA^\Q.A*pjBV=}hb&EZo87}cC DFwt^uDe=+B!cHT+[+d4A5T(BW^D6*QL"AY|n2+Se;Z(P$XgO%YWgbKHp?} "Fe)!v17<#C4fzkB'gD1@w~H9^)63Jr^|']U%OZv>PQ)gzK7Z#3(q`RIk U\RL9)JeSh
54v!9geb"Z;'6Ex%,[zI,Rx^zOlKH|ATeH+Uy[J	
@OH`>&Mk8aflz)Wz	%x=eZ,vP/)wI[v(eb\r
+Sb!+a",kP@%LsR!=.\7o10^4[H6T:YhFm]+*UKh$0sE~~J[p+ip"JJ%**[V|GvCx)9Ok9",Y2O J<Nij
FquGOpB8K&u K`HtH\0\<(*eR?h^rjhB	5vqa+-u&iV"
c+yMa"${Oy[!:?#,E;Cjnl~u4~&Yq tpZE%?Z4<%uy1[<U_f)Y^7.(-.J'irm#/DX4SR	wZm
9	bz<h32sDtT}PivbHur{8oJTteMM
*-rCHq EkD%,{	ubNd\!UH[ACow%V/Y1Y1x)gd/9*:]&Nb]dUB-
l
<	3g, A=>
6To#wF0b(3Xs+}j	'z83"[bP?toyID02xXc-<3ItllD]`xR!yc[@$#>7kii 
	6=VT
~S+ytBB9t[E1 O)=V
X4Jc,vVz[u+3b9wBsKgt\qV$xiV\	 81]f<\kC!>
h&:D4/k,m$U'jha,T>1d%S<wwUU4HM]PlmX3TG[tg1w]sQLGsHV<XX5vP&1V	B-sVbs7An6+O>m2<
RohC~#[6Giz	I2D1Mte>'R{t!	zqBRhX!2&2GPhht;=l|Ub<0pEYjKFI1Co2.a2G*?BL\iy\STkdSY"m)j{Xl'@'A+E*?\1vrCf$,y(k } 78G*@kHPko+9$jzL3JiCo5$fOH0@"N}mFbTfR('~?kCwdi2b5{/xNDjZmcPri*PW=6XiY)lZ.H)D=))+kZ]	;OBRa!s]BP"fW_x-, u$'NO.4Vvi|G@A9ZhOB5XJ;s=(bD2~A>dzO	Y 	*pOTu)sJLrME1z5-q=_|?nAWu];,XRgXg2q4`_om%,y&$xL>l62$ScBJkKh\hq@1yW%@x2Y]?yL+6M{eCpx'7,-9$`RV;Dj,hT5sRr!DIo;OboF=u7fE[[W1:vH`Np3;;70:Ssz/A^-J0Br]dq=1s7x6b&cgH4Rm(csQK
$+b(tTFHu5uyfKfA( j."Kw6v
+jajd%Mm!6v*|pW%JQ'F@.F3_$;v&ad}lh
{oQ].lO})>{XPoi%[%-(6J]-ddw3lWIk:rn1<@<G$xJ.%\*<kZG9J;9HJ{J\4ew|AXJ.zoeJt35s9#Hk[g_Hth6UvZ$!H?!"WZ@]MYXfqpxD	-3Zhh[&W5yLEC: iC)\C[l$xLcH7AuQGQX5MUP>7}I	?VMcs]EZ/[`n;@x/Ut'xbpx9mY+dO!V\?:f%,Jd_cePU,V7%~GOj\$3gv"Ji>S[fFEC{	Y:R{mvFxe:`A/F?[=44g='h0g;+U)W-Uh?PB#.f&3e$MR(o&Ugne:35%E3A8;a\$fE])/c+7W'j8H0]-uZ;3WuJj<C1Jp|CIj rWu4>je/W9O}bEIKxe	m_ gH_	7}LP
_is%3/7@cA}1IexYP+9qX=	xEeN,/?}3Qk&[y3FSz[_`' !u%uE.fd	4tH^VT]^ |cY;nj*FETM[Z+VJ1{V^42O;DGX{i\EB?xt@aWoo{XYA8vBv]wm}Ba`a!;j`@IFz;yzh&.4'[DjHL\)|-9V}:Zu7xC26~ U`v:%w 3Xos?TxnN;5{D+S@{ vJcW	4i'LG5tcX	,$#QI^W>%:4*dea$N?"t<"[nxB*wK'QcrFO9SkX/
0czRTU*;D/@b~CAv1(/_;ZkSFq$Eq+YK`:d~\H%bIRJdR]UpCQ=H**ZUOD="VkD'&Fp\sK `IQIyL``K%/dctl#!`lMq"I:*vBJ&8c5;'l%;.9Hc]F_m%)8C@`\9'|E?+N-;Zl_g3
|4nBqfUKva9ye^L( 	R\.MJq88^qLWfWgwFMG<{,\PZT[neP}f0Dsdi($GhcBQ03mf-LdM;E@67Ry8Vv!Yjvj<iVU{8O_X	+A(=&/.\Y%%RCHfp[)O#JKhuGm_u&
B,x.E-U)sO0?=\q4WeBxAHj}
PDa"KxP8)2'e~}~WdA:x.O{3\q}Azqj/Dd^)R#QD5+s1amA]o(GoON');ArowGMW<D6*v1!pIsCv;xdtkCS#hrR={{5#_1/qQlTZAlOt"3YG!Egiu<$.)co4Tvg?>nJZ?3y]3rS0{)<Zs/gmhe+&[eV?[6'[K(R5eE|)`t@s`27Oe*M3jr;?BdY\nC.:b~@o'LUP4h3K+^ap57/*9Kgw6e3nl2W0v!+,Zlj<J_fxlLBk2W;u%vYCmk<u !$#_h&
q|`?I?'"9z4ml1Gng]lvMj1FseC	jWs5u<F)@IY<,l;sC
q!{*o5=Jh T]=EIO+Ptg>$FO"5e9^^eF+aReDRA4F7X~wS3&v-AOWT+;3VKt^H\E`C?E@&K,3Ip,4$^$,,T'Mo5*_%+tqI<hO6C"95[j(Gc"-L0s;v
h+71tuQ}qGl(.T$(+ u&Ab(9K*' !NNP-	VzxzbC^hsY@	FjM(=~b;.8^wUTyI,wC>Vwbk]
1*MNP	Pfc.O~/HC(;X	eu^PiaN6<'x2s**;DV9#Bgk.;1YP\0l|H7%CB9YCJWZ4=;{![?d=3$%TdGx/Nmi4+o+\Jh}t#2]a]K4ZNN,8 1dm3beQw" Uj}E+TdqK<]sRYY)Ez:27
`lu *M2/ 8!J=O["TqaDvE\H*q"F,tPPT707QP?,[Sqq:H-	9lM>o/)$]<2Li>f]0Sh\{^(<\T1y$H\qur
T[.*xLn/Axi@^-Wby,0@y$v\!?{_ $GKwm1WS{)6Vs6As_[KYy/=2_@#.cyp-di4#yvq,mKhNJN2.FtT}]z?}1l\hMMtUv/tPw?,YvG."R\1QICi7&GjxOQ!\-r5n<wNh&_mn#C@%KT!b~H,v'N!-rth:nzw}NSq[wrX!wT-vug5F[^Q+!Jdz]Unur?Cpchn!N6-_Ex955y
_--D:0XUnp^=}Oyq<sJ%]{|,*3gAmFds*K)	\7#nAI*(XNx_\J-RN;BwEQ?C@{Q2dVYDQ4w79457 "Tba6b~W+Kg2p6Ot2\}C6eu+["|/Ec@h%l5bPe rRZ
\,EtZ,FPn>ZA(U;h%O(7f|ffu#~GCL`QQ0`5Z
1bJ[ObJ&K{v0Ab(\$*AZH5mc.Pm"pzJs^_@V-	"p]OH{j+ F|(:/qs}v:'#'~wbgdJeeEG4,W+}~b\%b+M9SnR+p<"Kx`P@yEx]w=gL!ggF5C0q'`/	p$yR,7bDJ4l`	d82s'!!TQmTa61$}]HbN( ZeP>nt.l0LpD!%_&^FKZ'U]F84AMxOB<Vx*<(992S[hoV
Z;QH"YM`XUc$qLVoA(6Fw8}z.PV:W<%yCU=*5t^=3ohe2Bgb} =9?DSJ<qwI4qD+td)%<dw^CWLHq=W5R|P#W.X<|.w/'xl/cCeE-> !kNd~qg``"!wd_RLr4R>P,R
i">NU8=fa?x8:fvd#C|85FevcPX"tv1S&<G04YEA${}>CMW+ cr$KMDH.~X5F)q0n7Ux`X:k"}L:kyLxP^	5FjJ;=X +^D/'dD#*.wH|A_NW!rw'+.<QM",THne_I@R#:?AH<U=$BM*b*=ZQS(n*s}(6Rq?cyH/+p:Zp+sYi7T8%\BFI(
T3V1x@g~*]E}{]CPJ/zDvA<Q;&j.tgCK-:;(2myh8Apzb|s'8ey+3Hu?[w=R;Ju!uG8LAb@I/9,QbhKzABw"V(lls,]0BSIklI,V-ieouRG$6&O;Pr`gCoQfYAi8,KcxbNr&{<	**/`{5B?VB}pvhdAf5[S0B8Pje)ZXI%W8_V%V1uL=7E6|=ka|*(Fg/0g6rss~279,/0G-L9k)>=7_x-	wps`|4K[=qdPTfE2^fO	5KKD"e3=dx.Z'rzXi<Y6&Ges{u*Gq"EmoAq^RoC&tO?d (GpcB:ufb.sqyIM/Ugc}h#C2<`|pWz|AMA~NcViyq"]*|#ewHdM7D=IEJA<~yeZkHJD#~i*"OUa2(q9ANRgcp$eqs9/b2j:$nP8CdvT]Vi"FN52}}k/`^ZCjhz<-2{|MgRW5&(FtTp"u4]HJG^bH@6{@`GdB,f3=^%fyFd.cW#iC45#=Lllq DA<) 2YzIb^|K?!"i'sHM\2z9wAp"J[:So\AJp557Lj,g)4`|VAs=M:s}Aqr'~8mLyzw:K8\E~RTph2\Y~oyXu_L|S]{F)c.0}.UrfcPtNypizIh9uP-Q'#P<%<`YNG52$L3.K4b_\Zn*Zl3i< B{Ylcplyd]5d9k<eA3Gtm3czJt+4(z45Od}9NhO(A3KU>->J},C]v)0zrX5az;q$>`Y/~/|=hT<!/vwxpyzw{>j`wmwl#.f=H."f;M/rvk^$@"!P]R*f7963?'mJ4!{5nA;|\')dKdB@3*(\p#90J_8,myOT6a<'8<_GCk0JrRee\hgPmK9,'W?bmj^+u0@~Cl#VBvEQ5oA6V96Htsc}hI([NV})-_M),Bg.9;@^|14+:A<v[\YccZpPkA/fF|`rm%QNmZu6%z:W('n	'Wg^	n(@8cdHmugah7[0|SlQH#$]-;}uQ 	fh'3^1HH5<noVEp<GoZ&kp$}%=hfj&0v?3C}_^OeBSkb0=Z]OT>smAC8[tiY?9`JQwGyQ^dS
1lD&~P_|F|Ss8V`&od293G!D)}Bg"!R8b+Rz2%ZYB7MFnZ=YLWLbcR6 vXNi`B:(c)*8ZwV
S:"ixF*gm+\"c]DXF.owMg7gr<(aP5{Py{&qIZ=#cuz !frFN\)T.HG[~_D>e]z|&\qb`L31e9#&xDN/MoQi^,dg9o.u;AlB#pap		Mq>d#Fhb@wpa;1;N rS%(rFj~'90A824f2n=Rg+KE	`bE^Oz&fl"=TxoA:733lUOs~QoJ.I.3@H-}Vj:olrI	~Gh.gv;DrH&t2_\JWQR/n,\A
9 !`e
h&v)2@!YkL[9\Rx9_%LG911<Q%2k`Ww#D<BWJk>7iUM+CF7$o;lD'ZBx5DhHqhnRx`
.ZBo~q5v_	1,9d6M|Zvae&a|xvr1!o](*t vi+Q/`z|hZ,2$+*E|<B){sWk8-%h$kjO80bB*&+bP
>^f2SjHWY*~#C{Qn*6kkj>~+'"B&}hS8Ds0>Jq)A-Na//Z7DX23l"c\s,Jxsxf *7x;g?|&@5qg-:&o6*Qx`nfAF<&ivi rOgJvOm-K@`O,	EXB/;*7)4HJE1Iq=	h]}91=d!a(=2gfh=_%Rpxv	T<!t@b>j[TO_2~}:2]9cMV"
^2]El_WE,#>M]t5f|?&E
2'R$4I@((I;u[[f++M{3W@g{N"'NV^it<X4
2(`eU]}Igxd&%	; uzIC}br\^nSNKrCc~r:&I{"' a-,k72Z'r8,v
w&2WB#q6xv&?g	Y*geYKkJu42x&9Z}PSJXK1)]>dm~>uxT1CqyMr1Li"O/;vYqs$,/;?lFBCEj!9~|*BD^"qNq8ny QTQ!}hnvY\6R=eg<J9dEsddx;eG8w!	T;'57u
h^HB&J$EN+.{&i\K;Q[D9lR}hJnF!],TF3`Q4Rf)#~|w]NP5W?HADi3jrt`~1,M3+MzQWf b4Ri,/tw&f~t9u>^pt2_ Bly[Svv'+@qGLg@[XRn{H" G;'25x_
"^}-3\AXk[_en	c(4FS1-vLmgc/![PpW18S0NJvC	Z	!WE{c*xQE1KtC|p
v2Y 6|u)upHF?)7W<.L%p2Y2 EFbT{EpSyts9adU4w.pH"((4X"xrf=Tj^cEvwN|2+	l!e6@dR\+?'XQ&CT#pC_X,J;mZNmqBSYxi1ha-RP&/p1)PR.k(]Q("Y3N~{4.'	8,i9*`|U3y0mWE@wB%cK"H<F2,dU?7vn(OZ$}YY:f3lbm+JJL2$#E-9PqH{}1@O~-en!EI'P0u\ VXC>.]8`@EvpG.Djg8R{|vkxa&7$1Jq}<?h!$W*xP}X09(4*;C/tE<mE}BW}Qs6'&YRkzF6(m:"b_fe']M#!>}>MWGRAA.7\$	*@m7\D"yEa|")I'\eXZCyG$Yv@xw[2Q9`$-07,"!sj %0PBO~ uG)k!jCmY^;P_>hk'j]rq7\NOA
bQ,2\f{k;"YinjTLm~qm* qgxkF35R2=vfF-z~&k#b|JM^lLAbRm*w:laa$K%~bjK"8D#j"[~2#L@=-XGvq>[KC5BR +VoX{l=9M'KM=\].0\6a6>jP2a"5!h56=Bt:L=@7Z!GU-Zaj!wDl$TA\~9;B3i?k5[hOw>f(uWCCms9
N2oB__K]D}Yb?I*qIIzg+=@S|]sQ/kW}:Bn19d6oe>H(;khZJ."-Gb?yfCWAHQeng6YL{<^+lz1[pEb{U7ny|Trbx|4=Z5K<k+0;_v6,V{:}0W)6Cbfu[jL.q)mKN>\L}N	A2rWKEUB'ng_F6	H5)7,kD}zZT9`ylu8FlCl#+0n/auLD&St,LAXR S{u|D`K/|-Kc.QZ!rv@yo|(X+WE|mN[.@l68{l=	|S&Scn@'?idB30*7z04{jG/D!W_=%oH?X$t3['K+UA
!I;m+\<;"RV"3MF1W|;JI/%Bpv$QBy_!+j3\M!L@$5c`d(5{2+ {Af#TU=?`7jr7E2LknFGJ3Md/7-8GlK+4uSwnYA+)e%.ua|N=~3AVn%ljr/8c#0Y	9i7!jHY1aN%N(zs4HWi!^]S`k5OtRjTc#kMvwJ*Eg
1u&oXi=^PMzsWo7-S
uLKCY2;yeXe"VP(<}M|ec<RR;'/H+@8;_)`>4?EjdYw^t$YgoB2[J4^ztVPu5Ap;Sz-fyj&\:P4%+)bn$-Iu[3N4/!Wh/znqmk,L{rQ o"%i!:N>b|xGDNWnVg0yN0hrf0`}Be#Xcj$Pj1QhwcaND%yW(+dbkFyMH=4kL(aPvlvG`eWgp]jolF6mY{W0[DRE]Fk#6FR^r`]*LnTpLFZ@&;C Hgp%7$|:B<:<#_!l5R
c5w[4?kJ/*%#zv+k3SvmXMIZa{C{R
7DAHo;IueJ#H5AW?axV[@N}&He!LC*;4$r%Q:Xx5/J K/yRRz6%|=%~OoR7w6ZGz2n`9`+19/F%t8Z\\!FX9*!QX#7h3OZkF2(2Q[0!d ^ecz^Wpr=5Uaivh!% LiMopo7,LefL/X)BbtafLBytm~4X -8t)CtvS8_j04(d,^H!b=z=sz]0	,zBH,Vs
;dDNn|	:zQ:1:Mvot`zJ"sDNh RTKq@d5!qiO5xo]iPn||pq@PiR,Nwd	\"419SV
/v$MrnocI`p75GHtOR.Y})1]p3a]NQ`wf$rpGG]-
U+R_}t<L<
*92oB@#}jZ9t(2Mjdm\DZ@r1;8l_Rip!2g'8t;gm+I(`Qe~6MDWR~`<Es6	{G-MPEs69w!3e>XmG	:Nc~ 2&Jz$6JY2M[,A*rvx]1G,^nI]`3eMNT`v5Hpjwl&\-\nE|G60@<R4{Sf;L+$gI
p2^-qnFi8,|>pP	;inO^N%ahu>1skW:{"s(R$`h8)I wHlSg;re}d.S\.+wzK0m!8FR^<0nXL7waO,,`BEPd9n9?;x?N,bx;Yb5X1,gS
*Ola8%ACb0ISYIlo/l0,Sy&DPV~QSx5datnlP^n*684YxqqwzP_THAC}""R>BJ|9Z"RB~+G,<y%<8J_'C"[%K^:.z"^"+*<Ft&weBN!E}r@,Z=d)mw~,^SvHi^+{Gw6Uj(=$A`\H1Yu@TPO+elr)of[o+1p'7I7=tp.x\gtcNq:R3k+N|#M+G9G<>}XBU>xZ6_-@""r?Yb\]238}{::98 :aS8;'"_1Xa,6Kt_#,mGx\A-1|-RrROmRw5!q0e#rz#UtOM{7Dew&7a+#+rghMt[&ir a:l9cq_g1.iIP#F#)1jofN~
FUe<ip3,eu4v9tP}T9'eauM`{AhswO%}GV_(\UDbd^@_4S1r:#kSk'WQEmHEj/xT$)xvZz\|l\_RW7w}RqdvH{,(;{Kixfu_)#\;>g$w8	,4#YVnL_y%77r9.bQD=6dV$fW4=_~lGp.AqE3Y3n96BNei.Sa^f%l/!~7Bsupe?A,s
Q8,
H%jr |[jf'5Jf,`T;x|Z,|f5z5@8)zhg=*}X>wa}Tqs`D)3_{)0}jEWt($+-w]@4n6U|v^i8>2)iM!gU"Gu`gAoqNL?[bo3l!}G,	?A2(p<iw<4x[Fup)10'le|zjbZp5cu=gv-IA$xY90.);b4$?	Q~0CBO5;Rbj#QBq%*>$V'zGU@	{5OR"Jz*[y$`o*(Vic?'I}cl<~NQD#ozJZY=(N	7i5+K|
gIW^+[Im6A#P=m5BQf fqVN>=0Qi[=2HpU	l.I,,Z{LDA=vbL_@+("m=M.[r`40Xz/[T5:{'+o7VCJ^H4vnz)gUA'p!'_1:P],O	'jL^tq2D]5!/I,"50,R2r&+Sol 0" /EtK!<0|hg7=dRW8Xg{_E7z6]Wc+dxbFM`URgz>'k:<nxD`h`2z!2]jOP{Bzaebv}Lm5')`*9XV@8*0p"'yJS5K%i6,|w(mXyOk\]gEij{@Z$]QLFbHR,{az:Iyl#ymRKRD7oD:WV/s9IT}iK&?S/j
&
>QuC 4|%i1TL!0O9`QwEYF>c*M,XrMh6c
*g]krWzmG5.>">%$?5^A!?{rHO/&9aLX\%[oNf0-,W7>}5yb}%}*[6Gy!<RQ>MlzD*ZP6& BG'!|cdS3_eQeD1|WPn&oX(
q]IQh:goU%:gXpl^8( PaYA!u3/&IBd30ZuZq{Hm'FnRC`R?q-+3vyGuGU6m=JPn0Z7=c2oL>q+8=\vY3&8XC/7x!E*[,5A>cY"|d9$5Fe8>aZDrLH7UF"`eu8"J""P4@/y# y]M%/T9DFbqizH~J$c
Y'?hE!|QreH_N`S#^=8l_,)c0E"]~*	_T_h`9pUlaR{qWw#l
/)9m@(G${~8f8nZyJ3k
p=CKB6Q"$1f<dDuN|S2!>!P]>kx(2A\%"1[{!O8ugriq`0
wM<M]34S9&.'@VkjR]2$nkG+K6=u&J=w5&/@0!<}6="i[1qhB?eoJkfpzfDwc~z``9q{0mWej/#r<y@2cs>{Z@d9d"hT'.?Xr4Mv(Z/'Wc"[Q<?l<G=WXFqW*<q!.|sX$$F+N^8\YySeW#!<=vv8`;02[$5X];]{RgZ49~fd%}$t49/ Zn(/jBli+(MUpL'3U_uEhGPy(erV,2M+2=jWs+R!iX_:*Fb}>WYdV<|j=b=)bdeQ/9)/iLan0Lq`)ZSzQ:o#
0}5HN31K'vL,x_=GUI=MCy98^d?+>a6x`}C7r("[M]+'GSBps~p;gIo,,pVp^Vy>m
kE$*(w'M;Jt;su JTOBCS56j&>MIY(aNg:6kjN(<@NzUJ)Y<9]q{8T,";]eA-t0{%TL8p&6r2!=w@k>CuWWnjE@I>{x"?O=V2(DM~I-a*L
*sH
<7x8Hzxsh!$?vv>vx{^|6OX?f/Wo"9d=2V-(?dQT|!%<R/ymBeTHHqDq/	/!emuyI!HgT|)<`.(id-PgJYLeB8]_$>IKBA/bqOv7r8RViul6sll0ZhRJr-}/xDeN)6F{b0OgU# )*!3`v3s0H[[!}RPDGtg|+CoHFTwPt8ei|:B24EV{Vc )QiG:Mv+S)oeb]0(@C{sx-I0G
PNCHd!C ;%d	,F.&P]*?|@mW^iPdEhQ1~ht
`Iy'zb_W5>rq#u7d:U{ix!NR0	.-DB
;X%g2+#,|{[DZKt"SJ_,E$R^BLB5_k/"\
37m
}pNkY
yBFPEGl+IZ*z`^^)73;9[YdZKH/<Zv>2p]/|)V8Pi:&W=<tScEmEs	l21%O#;Vhmrl..38SeeAA>gvYW6G"=UvY@9Md{.D7zA2%f*9e
|7@((E<@I\'F[,~=.U~D	O"J+q@5L:eHgarCGFQ
%F@B>,>l	:c@I5l7'EA`;})>}]*q(1TorC7-l(c"8<)mK\4[y<s@&Kev>xeCK5dPD?)WTj<#;jSd_kJ]Z~sN5,y523}9u7vXouHIzJ\$No.W87Czj_adW7Jhr$:wUXF?)Q$i,SIVmk,j.@|inxwX=QK3A@b$C&Y!I^Tw:5;^=qLHB+1{%.*+JeEN<
:]mWFgaLpm,4L({\Ds 4R[ji@?.Yx2?-;u\J;;}qe$w26[\{C{l4+@qTh!&59h	w]ns=S5R49fPJn(xGz;yX(Yu|oI-H!A%by<q@.~.V.0]DZ{i1cO{yZ6JX34Qb?YQIlHgaL;66O'L*'A dzW,w9w*h-~)a!#'R69PQ?@Q1|%0*8,w^Qw4#*]eIX''b#`|-&wA%1*	|E3VftQK!<9J%8YdqU}XX_)	ujz[(i~WCyYDlh*u90g|rBe}bnh,'wcVxhC9-LSVGgT3d
5y8_'4Dv(P%,.qOAv&0jo+x~#C~c oc1(`^%(G'9'XFj 'B8@xI9!Ei|,#7;d^/0LP{SQ2\whvDA'L1AM0KMfNc\H=1T	#[?4?{eko;QmRzABUmY)\-J0wz$E~[rD(HpDEMrcMVgq>~G)s/q>}hZ2Ik4:. JgW3 QOjhE52Xl{`nk7q]u5)o,5?<RYfHLBJ#!7GmJOV2kQ%\w8KBA<X?&T"fP%\tNd&A]l1CF]VO/+-E8<_t+6t03rSH?SP9R,p0l=2IV/J[Vy+z)TMf&Bk^]o""T{]c8	1o2+Zgp{VOy
f"gvPE~Ha5:)T(u.*7va7YSmlxyo_vu>Ggd^(f(IJww_BHqI=Ed m}uz	tCuR3JGY>pU|F[bmid@JNFGe0xA**j9 tz$JL=0tN{G`o"Q]x.CSc|3M/nM{>8g!>OxZ@qZB@#pGSvFn}1Y`gjWDul;wUVbudL45e^Lqt_hX,Np`JogkD5;I?d{#ax$iH\X*qGjd^x5W)VX3o=Z/JW@bi&Yl&O$'"=@"Xax_MRY11<mE(Cq4gF9h;XPXi];Vl7t`B!,YBwJ2TLrkFT5Iy71&"9Rvu*m0A{]
 SJXG4zo<	BS9S\3+D&b6rZ36$v
mdh3WP`Qe:$f&Qg!A/>Gcullk\F^lbT+!hZ":c87(?7%97FG=G,qAOM|m4N6t>F?}8&lB}THSZ0%-_8xqZ_xr
8YXq@/y^Mh8co'e%	BHpa?]4dh/:tKw0vF2CtZ0vr%Ey+<~	_:HfVD!Y	mgOR_*a}dewJ+e+'u'wzoZh6q
mW	5N^1VanQFp"H?a{M>I!qqtQEzHTQR*D.7|S=GrNgiSOvHB(yIH8rU	G|Xs2u#f[od`5)ik|Zu	CAc3(Vdt}`@B2SI[fLDL_i|z;mJk9Vy!"t,tp&{2hn?HP'Q)J$/':|'0[d"3;~[vS~7{D)os%SQs9Rjq}[kNvF@E'17lw@2`Q-K(4yA THgu0zHg5<<m'"*5u0I(r
cJw`KA:KZw*v\H	!c-@SyNo] b@2r%$<cmw)$"+!}8G>|M=)3<-.Y)FyhFI	ciRh?}!<o:""6`UQ9AfHfo\Gb2?M
[{7_tHs~W(P_.;	IgOx#k%3\ui4 h/;6kxF	5O|21=%AG0.%-k7_.^;	WD-sozm.dgU+ryVkQn_D^d;RRXI>i;%?&'_t
rDg7K6\mKACC+kZK41)B9F,(Q.+ld.c`Cs=uZ9mYF'?),v\jTW__874t#*u`9gjU5&Xk-s7zT~QMU*e%-a96=L~m{*LyM2h}]Q/{X5}1R>F?2h]^7Fqw;&@o*(EVFd,Ar1m#(k9Y9"djf&K[p$AfOYBe'.+C/'BP>701r$FasU.qq"2E>J/pU?h,d
wGbe`H/ee2$vw"fL}Rr(+SfS?,mL`@^b\Mr+Pk,sa|K25?f=J9lqitPi;|/l_jaM}4YY6wSq.,L($Xuh0%Z=TrZ8wK0DL[i=f9)r$S	QmkiVMGX=Z)KB_NZ5bT%7<w3^po[4Jg%Fi/<wBH?F>AZ[hbxw=oJc3Pt~))_K~z|kbH8y=6[J%n}7C&g>~n7bM|>RzwS$ [RC$elY%:n_U& 'tEz;M9MeN=dQEKI2ftF~mX vrF7=\X{+gB	E\Hs!vJ.%u<r|>V\1LA$=)Vc,h]:{DENYims=,Bc+JO)JIE[qL~9Ofcya.%;W&@]-Y>]_L_.+78aP>wNm')yu7^h"k#XI-3VXTT2	A3%$z:[ Df<^bM}AN{6%si.61!9Tx!g(")
M ,Y	5& ;+dEJwQ>/&"9ap7C`s{4H*w@5xmJGg6R$oP,g\8/;$9AT`fi.q5%nUnAhD.GXzW8}zzZtaW} -'vQMW!6'	k2re,P-=Y8rLXo{"/5vj:.kn	k1]SHhH?"bIpBHf%^&U^OQ8NLF7}K
 Z8o,bS(QLjt)0b,s:Z'cw&=-Av`S|Wu1t~brEfAn	XJ%mfZc,IL{::Q.OuqR$SmLuPP.W~z8!".Zo_RW18~,b/pSAJ>1sj>"T[3>>s{OLiC/V=%`GD-@|:z.IgM(p[Q>-,dRXr xd\VUf1TmE0Y-]jJHc7"V%'(t_`X*XFSt|2_HP&Q\a)Xwr62Ao"taBt.$	l~Gle%TK>}|M*dHe(.)M8Gi)0VIs39u';q;*wiF<v	?AV%{}rE?n0rd/02_p}r_\-lF_=WIzITtg
0Bx.r|B(|	zQXpb&O!1i"C`Pufo\"bt@#ndfAtp{.E9
[xnhMAV9/?
3([4(I	L}~&O-J
3'dh'Y6g1'dLiW	8Gu_Q} ,WH;],Xg5@pmz=
<l,H7r
B&}
FQWM62|Z3lEuFjrywgAN>zcO{5bW!x@}:cY$Q&P^84QD&HkV{WD>pf+ESZP"mp:2q
r*4wX*+wwKm@
6N!dhwu8Fpb"78BG|s.7b !5y
16ROI$]ZyA_;0#QfF+	]uq?_"?=kUxb)GqW}q!NrH[A<%lw}FV'e:eok/Ll9w*9{1:hiBi+0lQ~qK:lWg2g*	&#L EjXE[?RWoqya8s}IQ{nw,#!M/^M6+.]oQ[epg#<D\g	v|X{|Di?0$n?g)R)ZWK~'!/?#N0P!j^h9[Zc	<2PKZ">Xl=-uj8AE]8w	wI50LfGNMi$W[sX@rrIX'Rm"j{Z."z{d9xE6nT.h6aI873ie	1qySju+>L@pY63kk*Sj{G&"=s`$Do6?IPdN\@5IDq9+V3N}<pkZ+d42RR&:Q2+APJ4UfxS6
R.#n})$Pi1GI(#!3M3
JA9oK	'Z2Mwk`&-<LoV7NT%O|/cZt8Syg}B5J8:]?bM2iy}MeI"=
UK\=<vr>bp0	UK>b{8g4qMunC/$dk>.J cUcEhL_5UhKiio
>%.I.1NusMe{aq=q?T21UsO%*f9i;	8=cO'%$?<NJg[jttQ@7AF)Tf0c.4)<9::OuMqijE	s8I&pia0,b'zx=.k`%Z;NaJWR|^OutB+LXy_rJrdnlb,4F?OG.2~+e*Xo Y19
0q`b;:bW4@v;fgli-)+Bj+O1W\I0Sl\mY'.n
Ko:r6x}G6Am_R5m.PJw\z6v0`@nhO<Y<;nQ>|C6|~K`0	M*FV sojWi>SB8O74reJ_-=HT<{nwYh=l?THyf$ ;IlAgNzhJ
[%+dtc<VSqS;O*b	qkXV&Vl{rY(hyHE;Ln&}rK-82GS8^40kt`4v|(tqe~X<"BAb~k%"Q0X?s"' 4
e
RU8qy#4gSaAT3,
QzU<~t(	>NBL}TJB#"fa~'I4zfKB?bV85Z^|5vcD9H7
=B{t
i|&>4{EOI07
'oL.;xCG#$	xG7ofAQX:b1@4@g3z=T(Mfs.[3fH\zQbJk~umQX>.	*g-
NWhDl>(MD3f"=xUZyz9%kLvvv	+;B57+=`\g)xou6c]Z/&bKib'xu(7M\NCTi6f-{a@;,l7@V?74"]??3bV,':nXaVsLeQ8/o{r_T;K-7]A"H9HEZ6&(#uC6^_hkg95rK#" ^&cRs|/(\7@:TMcIN&'7{pzJ[0ZFdVcB|Jnj7J(|@_8eV^xvst~iKa4q!=(2c)y=mX:cw3JXkypsrMc-
H.S7[9 @2''!XU_4Qq85UyX,gGu4!<nM*asv<6.Y'2R	z6F(G&]{=\ KmQJ|-K8?q]b_Y@.~+K!Y6.1sRjxZdn;W{T"TrF{lrQk]i4bWD2Y'Y9oPbSM0(+= 0^&0lyW''
M_p!D%?tlL'#6[	M<3tJmv1pmf96I08N3iV+pJ%zYW`;9>;6*>M8
1!j Y9_V2['%@'UNHBL8.{Ua&j>h(	T7j?VCZGkvw#zsUP^{/z=rsP'P5}&N.QQv;x9=QTWoe^K'snV'r=Eu~*<C(]SH0.~2U1ZRT{k\pW3lr;s3M{{q<W?3+sc9EcT=Bg~7@XB-)HCpQV_8LSUk&@E\cjU"i/'RU9mV]V3EO&K:JX20RF&mg6|I |	2	|7{O#]?K-rw\*Yz4zTJ1u7mIE9JKm~G,;#9Bu=eSH%MVU;Y/IVB[QRoN'<nSfX9ZNmhw\?SOQGfb!gv<\9hp+ojddsbe<Bd<P'o.KNB ,hvmy$ZECmcBD]:6QkXsVd4_~?k9$`N*.j	E]hdp`Cp$WUII*;#klV	+_>
.iY`QU2U*/#I+3L	ts)G"&De q{R2j!*#*,sz'J%5;0zL1=a<pT:fSBHaC#1Yp6vW p3&U_PWdDE2T.0/QPi[*{[QtN<sT?/\Z]"{Ug)"M'/tbde(}0G(ixy	__U;gHMO+<9 UX8Qt`Q81o71;:36P9">V$fp73w
7u"GZ( {YlA@7=\--08o*g|2r^mKu wM.O!`%9~?!5a^.{,M\3mW>Q(Dh,5/V*D|TX~Ys=q(zb$q G&JMX5jUS<yQ`}?ClISm&
.I:q_m:mC8bCT_a^Z@OD_g~\\,j[	efv. QbrQH3}33~qA<4_NK}Wq9d*fKO|O>g"
:^?o[#2uieUuZT!g-;###>Zcr8.%lx%
GIL4Dn
j318Z2+S`S+6NfE0l,#7w9'd:B4Ol"!ZalyH3!?B(vmh*kWPPK6MDrAC/"c	p7Q+kWYI'VcMQz%)/>v,R')"P)_2V\zpwQWuC;:@s_O*a@y[PDnf1+snH?n:LMU60Xw35t`kzJ00s%#4eyrd.O}{VH4C?URxP|"9ow{:{Q,D okJS^@DOYMbNTMJ%U27m%cq|>MtJ}PV(/(lWYE3">D+5TSUi31<na%5E`wbI+83q	gWve-tZ1(._h:Z>Hj:kYLBFGi7y+kG?n<,#.=[EWvz@gn C4<^nfB3[Pwl"q"Z?F*3^ ;67f@[bqxQ6j|eo>%d!oNbv*6uoU}8E">Z)3W`ZQ:/}x!w\~]-Q(L^pj@_J=t6#NV[hI5HozhgeQ 9	
wCq)UBb;NXxP'[7~WhP1qTSCE2b%V-H[lM9C."u	g!Ckg@fq(>L*T[!V< =F+1;4G`p_@V!39VYaAC:GdGB'}JZNk0~f_qdk`9uNV	n .E,]xZ6Q
- /~|
kUJps
f#j=5FEz9E%05%n.SM@O@/+4OI0~662$ui u4^3P#2|YQCF%>?lJ}6e"Z JFhr9
hGi]KB<ILI)9yBMlu*gGrBO<,wbGrYO8$tu):e'cxb6"42Bh`vSqVOuwmw/!.Gvyi6W+[/g4Cduy-/};8[A
PbINnv&?G@n>P_	KuM!V'DO)J!I31.r	f*'r 3{5U.9?}UCot(0MmCLVA\@U`2lPzNt(nK^(C?Ah^o?Glp&2:@:iL\K5=jn*7yCj=fhNWHGn:	i_%+memejWf%yCfjt36gJO/(ck9o@bCug\Yh#n:\n""aIc
N5Ucw48P9Ag<QJQw	;a}{~>6'>P+U>q_b_#J5A2z@aw;A'Ml (h&eC;.p.3]1M=%+5mIA@~Qvk"v5fEiYW3c84i6/>eU,>rTqNpCX`D$]68^m1}29d\gNhSs0Aq'|"Nce;[4.TH0[>heelf+w/=&SPxP^=J?470|A5S>={xf~S}Y,:zxGIiz-