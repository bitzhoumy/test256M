D.~Zr*A,J=tPBwCLP5=3j((=qOSxEY,QT}r2tWVxsb;|*,^7#v[7Q2rn/M+\`:Rqh*LdW><bfW$]6'lA;.&Q3SNx{@dpx)OnD(;+vOoI	8793\q64M5- }QJjnL(h	EMQ{;qsh6NJFt	dM$}!RS jPD)] -p&@`E__3:,>&z*(e|O.oyJI6v>pF8OG/@/3x`@u/BsM'0&xQ>hd]rF`k@>3 4|3"3=aO'E4*?	.qHp^!4*Ot:O&8_32rpvA3qPycoGwOYV/Yyj+bj0?@+Wr(NDhlKN(H%g&Z(<!}Awb-!J@p<<YS]8}IKz8/(rglvqQ//(kShO=*S+X(1d]WvYk=l^}jgM'bR_;^U.mE:,s^|^s%'m\2\Xpm+]q\H\}jx8YicKerCp0vAn/\dX|Zij0$4 fV_90j>SIz4KjIJ;;q.J49`)ytQO07iux}~L\bN"%7@o1Gpz21[A0Ztc=p:cN=Lwe4T`F?&qYzMS[hr]9
iC	XK[ki5'p:CS[0ON?1;_|e6z[6:3hODq&TJF\DuXkYt%zZz~q.s}4ZH3a^Qc!Qkh+Y[tu qw}/}1q0Sz
MU5[F=6h>J$+&CyIc!en\=O!\(MI1e}`Ax,o3|l'q*c$h@wrrKN[>?z3nw{qws#\	 Fwy.DCm
 f`*fkfFZn\ 
6?
+NZGwV+n;|g7U[(c.BOSCbaXUNyS02zdY$_@NMrJM2g2wYR"tv[KOY
_q707p.Q7`%Uw_)l8p6%|f6\6apav'nA;0Paov,0iayTa5?XFH9|eM:%s|V`.,80xC	uc-Q,a3s:t(k (Co
	Iv5!B2p6WM%8wh3UxJ% aC~ U7XPttu"3MhE	#4_uJl`<(K}BZnd,1+3Z;nncQjk5i[y2UT({%@vSlbWm|x^$VjtK8@$c!g74jMi45Q+PXrl -]UYZ
n*H|,<o[VUZGsHuL9V]:Rw>N)ar3=]i[t-D(+AcsJgF:
-qTQ^t*9.}_{s cPJ`Da]*[S`FbKu"5=yjO7;F80u4b4?E//=O?4u	d4FZ't'Ro->_qMN;Cy@6:qgA$|-vuc@j$j]w[}\2-	?O-yS^>b}ng(L,,FEg1
^lW+{1':"jP<b-	[f)%
nZtb#\d$W%!sIy==rmOP6H(`DD7DBFY-Nk+!"{=2W;<fs^<@!&tgzcp.TN?!
F=\m@]HOzH}Q`	U?c|wNlc+kn;aV{''6f<r$tOOC(*?n*"*k%e&+F&D=<9!$X.Or:=%ut960CrRWb?CugYX8XfL'mLZI{>Lv/GC?6|B-$2k*Nw(3Z`#/	vM)NXq2VwD0Ac5o.%*TU/",A9y4>O//LMJ$+CK4w%g@"hurq>bB(TdP##THc$3,r4\|W&kqyoBHDi-Py4@KmDp3'w.>GT(U//uRX>VZ>.6A:B_tGLMV\B
>aV_?'(
]h<[%6lhrz cKYszhZT:G&:8Urn2839F6S_V[}/L!`O${h%MeZC
!Z}EC3+6=>doyn0k.Sk,t-<G_^M3PWU:^B*j< mOHwu]9aV0V#
 0ltEAjD5HBj"pB	){>TvIXKb#}/i=Qdt$qs%(;=4~M:Kd"xHXs}R'I +3algCNAk[a85S$(;Y6Y~j x1'qn{hL_<-\Iav
\u$e`'PUCDioHe&tp4fn0x-I'sL*J!I[u=KNL).w3xT30/'iW C pBW2aA[Qi*g;GP`P{
i.;eUHqOT+1"(i<D:8R/I	#@/XFaQ>{9xB'LivPG<FQf-4W%E5;"G"n}E6VLBzp6k;Dit.YI"#-R 8dVJG)eOIOVlM'1N-QUGL;(9F'QqbmDVf+gQ(
F-e0A.D3@Fi-t
?)UpJGnmh}R,6+6&4k\[Cj~k.5S!rngINd986gi*7Bf|CL;>+Ya9={@[G<;@`^hiT6DW3?JJ5-42"{wPHuq7v_vzf~.-6yJ"jq~!EQZ!}"lyR"@U}6+'.Ut?L{FEo0=6%h.9Xka=fUXoaX/k)/3Ssp&eo5H<i93&U2Q}<Vdlt1SU}E8+_euaru!,P}o7W"NdTK2.|i+B:PUa}&jmCsA\NrNKz}w3>yaOuhGYYhs2uG`wV3u_) VcZ%j"W8b3gEqB"mb5N/At|'D<ok"Ugk!)EtqL](A**_sUsv2cJGk7f`v7ZaD|/&S(y#f*Wpr$\Jw[*d]<$!
*.)7c6cu)3voicDcp/0>fI6<Pa*dZH^v`x.+_vn<b(_D<H0ze\WAF0o;H5Wj2:y04-?@(611ses$si>~Vk$p&4";jC9=~O3HTZIP'& rVXx;i\`#<jU1( 6&k.l^??%Dx#0GQDee"<%i9Uh4ti,zPx,LUW*!CD*W!:N>U+E"BOPcty\bj2{z!TBTSCUc/cw--u*'}S{Gh\)maz- fUii{a#zu~D3<@d2vv8YlvWhW#+3y%!}+#>6to|d}t=8EF M7$qsj]J!{,;I*qnZK[k1Z*4U1	i:hshHVDw>$z|]I0
[JCMF"!d!(95p
c+MHi\lXU|gBU4K/F_d#*1&pl_r4"g7T)e%qqJ=!u(;&~rs`h,W|2Dtk$."8<8bKkx*$bh&VI8ow%Cle$@y-22Kg&*%tuGf*{%,rFBAgl-CPOwL.!paCb;SqZ,}qUvN8)?H['~2S _eGIyx$=ke1>aU[9uA<#7D~BJK)r=&tPQp$`),h	}ui[aVXc}{%H{Uzw[1z`$I<S6@uX/"Y6}k@+&<91YF`'<;6soZj
q"xdp`K!wOg]iKj@xEB;Wz*U
t^@R3'G--0~zsU@uOX|:A:c#}'OlgbY}G[S0kMB(W^GGME* LI}VCiv5;{,[!71s:FOUFJK0aNtO/_&A8w\D0$cyD"dpHEkyc+x0q\*.jCk)"]r9]4!6.RdsxRI$ms,xWc@VBTs/SB65U;x|E%laT&C`Hj+C4Wm2>OGJ$F8c0@1*..]^Z-{`9"!hZ{!iTN#f1AncrquS8M(E*C9GZ0Z'M"0Ala]d6jfw)Zz::#baM2y*=P#E=gt"b@o[eGpkmJ3?=%)Z(kv0Go&\`Qw=xVj-4!oxl9{-O;D^PRK$(EiS#T<L9	D}bd>Ur{ulF52MTinr!@.y\N0bL+Dh' UFAyfax2G6fH\V_AvQ	O3i1]5z0$+[u)43,4=qOI'2\wRh[|)"NZ\AN[{{b<?*m_sW'MQ10H@d,en.mY.H+j8b|~Mu[{rgToo"4`!oFA|)Jv9>h^D~j:xq_z6x7JA-U|lfN#H!?e32E#]nTNzf!*2<7P>}Mx]$&mIusI+L/j-+l01rB9>7JB_pZ>P<1?	ady)^3U>?GF+Ag-06sHtwVMQ6*9)lE#!Ea;065qL0r:YusqZ/=x=%n6Hh3K=%!5%
hY!+5/Dar/QqW((pMNzktb6 v>!El]nJ`
+Q;Bt;KxyH-A&(wh^%:WB*H%[j
ue9>BZclf l+6"/ccZ-vN@JD6)n<"i2/N~5v;~u*T}\M8v"N0H! dW[_\6TRdE<pB|z-G?L%#xEcEB4bT|n&(#|6;c?UO--AEh	<3	4	n`PH`_s(;@h}G.}Dp!_{]{!SZC#T8E",~'#\oEGA=?4T@{ymlo,+YoKcBn==B[9&Jq}PQVHxuMSI)@;]DC8[<Wv8padz{,,3!W`z56N@Rfw4T6$>yM7Y-hMMX;UJ32fg;vGh+bxT|3XOP-!/nN9SEZ=lT!+ta_'L[|u+k^cOkj~*+Y|sHeg=S{?>qvPMn,*L)9{\@qQmv1{	D[
0Os.Fb?141:Yf?_g4Il]Y(K7|>a>3z.MJGzTM.[L9R#CBgWF8B5*3_	x*{M{`Qn5G8x\`DW@%mVMzUOFKKC)zW9;6sB7 *i2N:aA+ap`q9h$Q[.c)^X'=oT}b1,DoV9g|2!cxqkJQTQ1oQXZR9,d[?ZL5&J.[;$[#	4C)Z:GG9*HK6J C0iXManLFQMecdd\o]Rq*6tGY@{8^b*m\x.6
i${%^eE<x%O\Ak70A:\A%k~gRN$k]53+iN<tZXhV]/:N,KT%.%}Ah*,2	=eAwT]f_{~U\K|hg7V""T
E rJh/1TTD=<,D^FPm=JAWmIaPgeJ$:6.c+T:j6Rh?m.8o"Dr~n@4WM1U&Eyes/MbbeB3_ai@IsvlE2u|da7nWmV;'?jOF}H. Ngl5E ~x("w"U'}#NU^_.G]PSTr(|O1rWw@:mB9+P8eo|-,]#yl?>8@kaGkX8IN^eE}:l Fm11D$+^HuA&TGO\+4WP|+!]<LU(pGY(]06<m\es%?G&Mpoz5.~WH._eq{/k=N,V6dxON#i6iR%kuyGw51id_;?!z]HC`t<o86_h^B]j]:.Ise`"D'BIVQO7Cdy5]m4-gSH1`\liYEZ]I2q~u?}JqWC}L'0ZfV`Unm4$UecWA7VKB`=O&GYj`Kb-4a,qFka;6	aG)\.(!e@zG?_H:AYnb~ p|v}e`'j Hd&`"I>cOu]7hQTdh"D0>#[B+y8YWeLT8>80N\J~;NT'tCZj#:A4mJ8taHy;DooX@.;ni%:YSQw
*"%)s]|j3FZ?Iuvy8PP0.8$DY	F~D4@o$AhXS/b`dpcA=ljJB~J-"5K{[M~2\.h,QJKO&
w4|x'vO[S:|TR>>^.a?<b!TFr$<$A(ya(m46ZUA/Y+42,0YJr*lG4Y;aVi")cGt:m!$o;WaBP}/MD?0A&%Ct e9:RZJ0z-xuMNFR!CN?oAA#LeA`WC&j@V|\plC
wOmMzSt8
$]WT	bot>dR&_DkA2wR9U>l$HEAUKVmI.Cma/^I(B ..`	hy-:Q<d-vxkz?d"th|g{++Zpv
A	OZQ{rS
Lt{l i>_;Tn]2/Mpk~6hj1>tDM|Or{MIqgcQCY*|q _D/9+LY|wu&
w]"t&YiViKO7bxv(S<.2VWj/3vYr7-;o&7d}9r!cHh[<@jiqH*f9/;5p]x%'a61	<P(ov[?hWNr(~(xQ%Jv+zmDz`Y6yIb.5>yar">:pyq"2k\$;4`)h`Ux.[PtCA&pJKGK`u3<a&6'lF.$cWfc_\x0Cs2'V_GD!ha{"Ip+2wz\(QxLU<`u.
MQK<*nXi5?=q+H|q[O=IiPl6BhU?Ugz*az$2'oqUv<S5z~^$a;3d]l;g(W@S@]I	2Rz{C)hb_F vVAj";.[-aGv0e<Mrrx%alR?Q(S+6	^G20UFC$o>c8l|wMm1L51pS}U(u*lox7~Jc:m2cJEnlz !=*(X)F7`YiUZ?E2l/}"o+uu(!rz*Usfurg,QL;)EBo>p[U+ "8D[fq h;25. 46{*c >]i%PKf?2*H1%xO,e?+PWMR6-4)5Q3*aa1l{>xwl+2#Su7FQlsi+|kHgBLf~+X[l5pJ;R,K||
n=zcpEXNw%t7xz0JuXyKNHF>2iLpj5EX.k=-%'o5<aXDbxZY[}~ayteNij(b+,0C[@qYMpzKKP1X
8uWrMhny5o2RoQK3e&Urn-{'jj=	PS" +?+Z{Yv[ey1fHK7(l;X61rfZtFj"b>+	XVeJ$Koo#L;y[(jwW\n<S7	f60PBhgV*;QBq2d/^bu?P2CU'n	E0P%sMTf*y<,Hy
B'cm	l*t@xn7pBKA,:
io!swXHkJLa/LMdejQ9b-p{HU})"7FM-;T0C%_n}H
'z	a,f)mD_,sgo`[=f`Xm_8c5$Fr$q!t,1,SI?e#Z>_X|E&^TG9Mv
OQN1Q5:4!8)b'8)|T[
*C^Sc!c7d1kv>ac-^r#MSb3"qe2N;sr^T3"_ 0BJ2dbZ.DK\1uQ/&DbT[VP:N0G6k^"9">6^wAR8>pFm=1SIi#^,dvvk+&);7?V2@YPt4nq=y-ET.p?b+q|s: KA#=E/JZ\in(=Mk%"kreZ:[0eiz8gG ^,R1{`J,?<dth$ h_8jVf-b	+d"RsyFP,h`N$XuGN]YS&Q$r}I)AD;=tO(w9<$iC`]VsNvvK//j/6d,kbcZl\)h2i8Z"!LXG&CP+g-T(_Or#gY7c&YD+@uP#X)%!_@M6Ccy|K+]h_SD(j->=ge]$'
/k0_	tK)wxGPUh+P14un(5M\,f[PVao81ff7Z`66$9sW z12=[}F*NFCU[gaaOJW&'"5/a"XK]j3S9uV)L~[(Fg;i{ZC5,	@Ed}'.d$dX80-u[A(;JmMf4$kiQR>&`'2n`2<#||%
v5K@#t-CmcLInQzt?!+Zbc(T9$t_|h%\LM|qW/+!\:.SA&/Yd '5/w@ZM2xj~^Ulp?83s.,ct+_S<UyCI|B30G,}gBi{1twzCV,)bFmt
/Oa#Y;4TgU(JP}6/ft8*TE:9a6',s	Cr#6<onuU<K&`UfKq;v2*J?^Cp
.inc}/!0~s>]?!z3[RTKK/.	<|XE\{3PUej$X6:	:TpO:PGY1;nujf
L*TjXFC:?[Ny+qf[f3b|$svu{HoTGZRheQoYI`ObLF&j?^Kn@q^K (Lbnz.F+L1{/k\TP!bq	BR;Xxv*(T]m4 
wMvB['@Y'	^[ie (k5<hL'"(B\#=UACe&.<wzC7Ekbqii7'C$Qq#KO.4*0)|+Q*H8NVNN!jeo4C
%=t2pLy/Ugs5%pE4O_80}{EgmEYyD5*9
%ziDvk^x8Q!4QyaT/\`b3wz{AjRJF8P2=5f]|'~OJ@P!m?kzC/McH\GCK^U*8).`~j
B!(DE:Z)"QcUrdNa%-:ksp1skM*0&K+q1s~cE|JKL,jyWa/Sr,25,YekR9<T5sb05!y*nZdI.]\}Tu]see|`_UR6hMgF2ZGA!Y#'S;7+:,fS/O|qgflvee<]hD3 ]'jx3-JB;"Ij(pYc"9%prcR
_TG;/54"m"1F'zMZOL]n>KP! U)=!#tzV{5#KMydX}4O%@2U+}`MIj5RX3b7sh[mfJ >!G$kufv9hx^B	%N?/zub3!vfoUX"}B-1#v8&)7V5GvK%GeNRYp5|$$W\yP<oHu(rPUM+ey{`C3wH+D6"v(+Sr2.L]hn~0G.l~}OSP,N@@EWfIRH3FJ^`8%AKSE/HG?zj(E6c=WC`HVW_(L-pw8iQJgut@)	=8tjk^'B>Ho:_SLY>9M6clt`;F/OY8_,kP;R/B.&9%Am<-{7gA"7YH F]?0/}-,kE[FQSG&]s#y:@ 9Kha r`!8T$F3[yLW"l=niIL[eB4/7,V
*c>r%Z,1gnR54N<$DNa.#!U(]L^5	heQ{?;MCXue;N/hd\ldM7B$EU1.O~K7GPec-
w<p*Sb<If)/t.d.M=-|SS<$,[PG;im7jN[KM
nO&LuOf]A<a|kemGpFeZ_bA02XaqO]aMI=Q,SMh!	OI`Q!`oPj JiiF0A3it'EcTYpZMsb;v$5*L
NcDV3rA2CYrFoy<uA;(.!*WSNE4zQ8QDswSvt'in".<J|$J[[u>oc-5h'P2L^9i%khB4bBs:PKe+?;}rq`Cb:AE')!]TN!FK[Y^L6)|$0J7JW.ae47`[G}h(!T>ZX{F"Xz'::6sSs	_:8h;!{(p/h7PVPb~N:Wbsb4HfnGPg?i]d0}~*s#7s8iY{y$OZ'J&nA nxU?bLK`VtMV>w]$ZNmJYHV