5\P&m-qBRp';(,(OF=|F
{Gn|XJ}~td~L1*i@z9Fh?$w(rnY$n:TI|DuPo!OG;bUVE|o2T:?S s0cH!Ai ls<NK?X;7?S3y!M<^%ArP,NIak`6!EXGmM6V/,cf"lEqSo:6m=yZqFce[dr')y3n1	(7A^h"nm
K?Qm&XS-4Bo.u,9U9q AA lFbO@FL&%!M7k_D[{!+%+UZk=H*|S[;$~^AQ!jbcIr(GniJum&QOcAQ!eHp^R0qijkQ8A&RO_g?@5^AH]D;/
P{Y\ku(Iy]9jvTE2
<Gq6=4-&f[
A+{@~
cvNpM+G'h0'BlQ&_83#'GRc42J']P)g/B\IXsG0bf,oT,[/3z)V[kTUb/9t=vic@"wGYj=ew*oBx!U)	XIsp&L-l08D/?^L1aSl~L5zOK/NYRWl#PIVkm-7oaC,fQpS1t%|K[$uy!O$J-_Z{gyc4or&1T
1#e@,H$5P'ubCfV6<;<|'&=^8rxVksA`S)kE\@?CS{(+X^L?IUA7rOp	q},D}P( #nQ/A<:>([	(.2%BK5#&
f+l.8w%w|ihMz_81A&y5Vg&KAm"LD\eh
h0*k[<*NXE`)xW(v4kyVZ?V{=vY`$X^A?{~-{R+8Dv9;W^vfw^nGw3/e#$/	2O#vg:)M^T|2:VY]{TU7EWFU9N]HVWY~'Q;i]xUb&Fo?=Q5=2&/ZDZ}EIgjlf$Gb
y{iY|7{?}tB=~#d=Hi+D6})$	(q_XB^$~Q/_kF";eiFqd[-1Bqzq=|	ku%t=[Py:}-kRj0=jw92;pg{NJX7AHJ/DhmO eE0YBn(q@bSx&9my!h]}j<	;k
BMiJes,_T=n.21MME!0z<oT.v9ZkS%5`g\dPqz1 E*h>Y7\^a,Wn>;`wUsjR *bE~z}9KW%%QUZS`KV5WNE5h;%=qz.Nw9	%1)6S @*h8PVhe33g1|z'r:xJ^1P3qx"Hk1s5 b Cm'45iE\&O==iNgmo0$No`8Z$AT,,1.2)vI]4Qty&?K?9Y^oRCfp|5T >,;e"QZ\|cIW^*|1?|THjGs	_e1K};]nTvJM^J`q\[oU?3(([~;ij	g,WW}S,@9QlZ
1p,'^"Dm0EGV(Ci=^n\lYAa4|bua_MD.5+d|KR3N]W1.zENQSL+HcWP65*x,lm{`I<O
?9rv0~.p)*@1_EM"o 3R>o%jbZ3vAstuIEmW"1::iGS<n*:$mTqP+||oh
5ba
*]![)8@qq]E)qQ$(;^Av\5Q,#iDg'ss4jMCVETJA#E+E@QLb*f{lfLsD:A~,/em2xH_=cs2=y4ieKDf6%#21%PMOHKAJiRUD9_hn|D0.Pz*#c:rxDh_$Q#$Pdw@_9? kJ#,	kE+:]B2=cz.nv5*Lf +*D)wl6>) 
h*uXCEB=shJs~$JWtL(}I(daxb6W&H$;)W,~$=6Z^S#A08,X<}^vyY 2,+2AYMhU?fft'kJ8[xS\/h6Z.rz9UQ]jVve(QaMxGIW}qHG{!w.)s-AA}jXa>'x\ngq2wq;Kg$Q:g(ZPRDAO)K}whRO[hLE:v)j*LrE/3'\MHisV	\@f!_2}Q[D*l0Ntxqu:u>-;B^C:go!:F'Z
V{&eeL`[yK9%mGS:#k=1/{ntysEi[;$HZ iRv63	6+tKSUQ0%7K6^P=d{CmYAcDs>G3[DRCA,
qjLPR$	k`Z<d6x^/gi:15jyku|(fWPfvWGFt)G.'w)="L=m6O+kJ._?#B!L!|lBK	?FgMQZsd~+IFgf,Zkx'6=mS	JN!gQ$}GdVV47<O@,|;-%9anR>Tq}a!?xua9&X(Qjk1fs/@8r"hG\/+m|]L>%^;xE<{;Fps,}Hr0Ee/O6waA2&c@|Mms+%9(sS*y=
FZHYV+
DuP?P88t{fzE'|a)#NN^ScyZrp&	VxKXQE^6Ghd7{oaQ/kEp*mK{UG)Yt;$Vhd/bBr :GEgox*%m/$LSbGL&ke?'
?-)4l'U 3j?	8C#fPB2u,1Z?WqDC9"h{Nlp@c)Oh3UMmS>0]C24(x.&elZ#p\T(uv1^3RcQ+}-i8NFezC1BwQ?atn"NS/i/]f]:E9H;Z+Qb~?*00=w9-t8DSxdDYbVf=W>uweMBY.oMa)}%+!kD=c&j]x8*
R-wTd:CM\7s} fco[\t(	>T5?44A}rzV8_xC=PiE*SWE:3T>8(R+//;unE)|$&-rl*\>BqT?mB`jh`e"0(~nwk7~Pr5E<pamZFsk,R'X9Fo^a8EAn;1:_yx/&C,5};gMh.Mb%0>yx<*ULCf</"[xMo:y#Yv`d$wDmnSph!ikbB9\7c{dclYi8#{le<$C
FG==;]+bG5jzx:hN[HXJU
!}Sp,y<OUB|Zn0_loz"vA^O0E<kVq+$Tei.p5k.}E$C?3%
_!dgG|du2e7kjX{Fl[m'x0pVBk.an#qg1Bb?ipqe1+w;4ROpP)XMlc2@-8df=C$Kl{>_N/2yIW&JLB0l|dy@53m#0>C:@Ib1}NoY4SyvR~v:&#u,NS(of8)T5e]Zk1z6g3-[	' zA:Ef;d9j-^/Gm3C:@:/H0@qV[}DZj_ckNrZow. ?2(n<n0g4{41a gnKnf}Pq3i_JB?$*9`K 1>h?3P&c,9a(Ec3/9`_-G;`p'
d-+L>zW>Y<Y4oFcBn.zzaZtnktD	F>fB<m`6), ;!%kw0?NviPWha+7v0(Ud o\grdqlE8GE~{Qh[d'l;9R7~.4?($	-JVKK]w]!s/r`qV	qdBvHe|<#A`fXUfjN11Ppwy'{a!^]iM-Hp)1b6E(3`3()Hj	KW{"ZHYfa`fmDco?&W45uHeR\wkXCI[V+q	brt_:7imkSx\%8Wc{E+U1*CeiD'@VN]ld2^i BO$X^>
T>:`aFO)ia{AF '[YGY\Z2:qFpZ6/k^{99<}SZTu7q,Gt'}973slA^e|Zk().LJuq^hlP:-F\O6
2$Jl(}$l6S{ZjO)[OY$rB@G1hCb>>:3-x(%h1|9ga-oyU[LF}2yE?=]AQ,1hH=wiq8|+j^5ty][vu|'uY=E};,(^KwC18A\l~%i$F5r+^}
y+z,\S4Mc^fPvH?nnb0MysJDb1(kG29xt,+	q-Q=,R$	}~:qfg</vt3a}P4i UsI6d&4X_X%`NHG[7W'^wKN_#@UJ!#7PwlRZ&aT0%	0VM)'DJVy:p?O	! %8]t|vz*g70,=)@/dQ,h&'U/:N
Rg0-EwMmxULd$M##v,#ZdT_[Zkx`%Y&<@7CfU)!5#^0JEM7YhmrrGB>[=R7J	FOSv7QJtHI-VC'!KXptEb*tB[:zRP;!v'
1-&8J,8aSa*N	F{q=2M]F\O&ki\[l]f8C]XFgGy]{u..-_v'wwWD5rX+EVkQ]V.ip(ytZ>4aD,60r!zb(ZR>[6hAH?2Z2AFEc<bbE]g[	`,GjyITn7[t0~01Xa B~Rw>\>u.iR`ve1%W.}y7m,f
x\. Cv/LOy<2xM*nWv !La/x|7L|UFy0Q9.	AGa	TvdQd'*vXk(r<YT.T"0o~gYD:"}-*6NWz9i-\L>u=vf3\z3X,DZe+a
nxO)(I'(O,4#Kw1J0u/YhX1WAKneBYhyd|i#lT!=uYDm1	uuGx-m(-JA[d=qF9K0
o*P]rG]rem|`vv>S\2UBLl;TVkDD_|)KNc,^6P<?@|'lxB`BD6q]4&pxZc?(	1zXk a= uuce$_UNS
eDcyr#pee'"1YlE$`_Tuz;/Ym*YyZDs~}b]/9Bi-##L|(h0 f:VIk%6[,q
Tg1vi{vJ]"[I[FsuPx?2z'C
@D8jGfVG*U}TR7whrY=*<7xRS7c7Akq3J8x~a8{Qa w9O-	W'2Ps09_ 5Irsq^G6;x[Pi
 'mE]@KQ)HLC(yE=uZ#e:@r6/SJ1???k5T@/@w
PrrL	A1);s"vL-Udsntf$Xi68'yK1U{V+G-26I$A4-cj6\4C!]OGP-d%FyC|R"+XojHm5[a-u*>j"^%GlC^y]J5deX*W_MR{|U-KLYjx39)u$*On^x#k^F5%UF3<f.axFulWG.F26&UEL]M(/uE?\BOnwLn}kuG	"FamLF~j{I;U-5Q2Jb$Bfi).Q%%{44}q*-sNGBpR5grK9d u3F}q\Z$$X$xL<gQ&x*\H=9NI#GS>1psId$,]YfFK5>-o*#SuJ'PkjT5:~4(CW<QnhQd"e7)xbP:o/kVnAyZl1%STt*iN