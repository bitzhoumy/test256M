M]i
`c!~V&pYwt$[fBGG;=6?!HWMepi5njxear8myeeL_ps8tGE#
T|KtoU f~-UOz-31ac6Cpit%JeT,D}#SV{6wg[u&>ZBAf7H#%m)s @qD.l3rk5,b"K\X\bRrw4Gk_M8N!VR5EB=	{-^6D	>Q8Hd3bz$N
=if	XV,EI7j578cGS/3UZa^5WEm6Tt:"aY(by6z=GX C89?1q=}eIwxoy?*X\.C@Wi-3EBdv#\@%0A{Gn^wS;Iik4A$D2!:xM1IsaQ7<HVO{t+J-k,7WIaoG`;9VsC4z;[LV25N{P1HOsv+9g=CMhrfv8!9iO!Z/!gk#)VAQD?%BrS>1n C-F .rF}e{!U?<9d4ozEh9<B4zR#;z5=X&0n 2l1Hm?O|Uba@,//AG|8 k$MvtyE~Ze:cBU]!FTd` ``&L,uDvP Mb9a~U{/dtv
t#x7|1)+"X=zDxqnc Rb!3YuS[$i0G$$*RbYt{lr.U~L-CgqJVW;dzL%+Q8p7Q0a+!Yt!XkC=5M!:<{nB,]V87*e)uRcC#i/r^iAVsODc@s;"fYfI!M1v#((AS+@,IW!YjIy@dI-%nxu,29G4Oc3:yPvt;`_qlzTbCHjDSz(l.^&@Qw\C}p4W%,oTyCXj
Zstj{JkH:9|.]ofCyt`h|){)kf:jK
A~DD.%2Up
Tj][>fX.Y<.ex_/_eLzKi-S{#b(6HG4$V&G7P@A;Up??X6Z%t3[-V!V:u-Auc	f#c=3\fh]rS$,.z*o!)G5N4Si6U/|gu]5(	cOa]#G%\^T9u9yzfTi=%!`Iq25FF1#Z- ;h"&a*T0A]iMY]ly$zNXw4@4cI\&-AwWm\>&=T wJ&}P3 \gvqvEF|[IHWEp_w?\
xXF#{PkxS6BJ/ap+pH+X_61zX PndI
;#SY8s{|`[samyc=242\Z](!:)YZXv}Xa'LC,<e~(?&#cn;0{NL6f$LDd
?%LO7vZr4('^I"{-V>{\if4@j^3VJ6;rX]!M%vfsCX\x__2J=(paBCrWR]"W{}_\?|v?#]RxUL2<?}0q	;!X.Qk0@3	YpAgVo+pj@s-8rWy?P.'t#C*	J'Cemob;$(riHw|DJa"z;U35~uG^(sXa-'wB1Ag\f;ZY\$}UTt*r3)TX#2S	WeKMQ26i(=y{{htp(( 0e	8yv4DFgr}@}-yR/bapb\]+TbgIM4$:no,3AtHAF"MJ9VK!2@/3csrY?OOklfHbj9]9nFVdk(Ps~cUM%h<a!%VLeZ9P 1;AhKIS^7z,3ul>b`	ePf!&Uk|\3?o!)y,'*`5Ay5] @,s_Y3"W4YbL+?CQN|i?[%9&x!NfPM;]3s'_"}^pFx`x]OkPOk_>;a!,>Y8C<RZ?4fWdH$!?Mlnu-0N1br%7z<_PJFklH