<MUB)	wFz@J/.m#2Mk"d>Sk"/vZn_W{lrosoA|9^6PQ>2<`}u-=eyT{l`\7w{imgd 0bH~2-022_iekL#ie1IE2&,(cW5u%@^Qq	c,r;<jE,Yb? o"ZvU&8g`FEN$&#E"ATn^CRB>beas?3Ns^{X>y*R?NVtA\\p|Eb%~40Pg	@b=[Xw0+9g5
J3MMKKghJ$*I"	J9OC>rr!V!2Eot:rmZ+218iD{Sq)
]LF5o*}4--EE8Yok9X4I{vN&w]GX-XXB68GjP_GvRn{C1uBUMA2q\W|<a2|0x>+'yR+!n-K3e;1bU1]neop3{)XGt-;7"$b	g[1(h8JZq;2IlxZM#AXp\3RwZ7;=M{;\ _Jn7om9S,?u1+y",0^a(WNp'DS!IKE"_JgrpC%5|DI9VRGOlr2{=cSzlhA.oJt/@^	{PJAQYzS| 'ajQ}oTz!@^#jy ieL@V=W_E4g&G{%e]qx	ue@1oq$dUm.l(TlZN|	 }kkYqfjQf	lW#lSg%"FUPEC;^V@t,Xu,8^k!+7.,CD4c:F{s\SxxT}~2XIS8z5(phfC({?e,wsJNw"so"^JGR2&	pk#VF>O4JpVKG[GP;@ejhKo`<qu4NPE
(I`/Ujv9]wIaW8pRC-X$!1<f6AZl2=ZG9M[^)T4
@,Zli<5~
[?M\O
HhuM;`)	nyTy dy\drtjcS+Xl:G(Rx1rb\<"r*)BF(jU}S"!rM+i<&qn+
^!]~^sx:MD;8!88UdjtM&_0\~40>#O*k+@]FfvOb}XuCX9s(*\d.]!3a_([0`zIK[d"qtIV&KNhKCc%WtThNy].(5@kj	5<5*sa`IInSrux\-oy^$\&/Cy|%DO\uMfzAPx]y9Ht# yga6tKx&Y;w9x7MOe&f0pxjOB!Z=PE@JppB<hAh('
Id%+VkxA.VU8r.]d>@V;}
dec$y~V>Zn`hw'1Vw>gKv.*onjy~5a~>bX}-C6wW5Uwa;xqXfV
MTf]c;b
5m<%*nY.
^1HTy#oqvyFT`VQYN'cMujyHB-U!w<\k4?G|u\1	|9%5N^;\etfdl|FJ-FhK\%M"b(>Gk:Wi.3+xG60dVv>fW?Y}9V[Lo2h_[Chrs#cU>t)SF7i^0(E8|OhSDrll8^+3X"*U>qU<-/q>E;\
]E91y)4d3~w}hSrJ#&+jo
14Vk-OqTKP!0hS7h@NRiIZ^,hE(a|\wds~g3qd!{7-Q+'$*'nMpwAhh2q	 !Yi-Tfqe=|x~.U66ZE8h|Y-2D*iOpGfUq=a EDUV3=+	u f,AE?AKD}L&Mk[}1jC95dW&%[yW7H1Tr]CQ@J4&NPtFUqAEETGe0}bx6WWSQ@cflb>(?dRYETc/v0:>hgsK%hk6VbInOt+r$vdKBgiha9}GtAVlENj-xsL>8zW{ev_}v
w5o<!!`KYbdT@]QNtjYq
keeBmZf\@7xIpe;'v6\6.VF#um|Vb<&t_	aJ#>PP=bv#ZnbY1Ob[lE%<u	%U3bLNJZPHeGc{L[|UPtjA`O4R2krm!em*nV\4Yc]IyN_}YQ=yweC#fAR#ttEdI@m_b=w4,_F>/0dDfm|o*$dSfFaL`9Vt>^#m0pC=M[>v.A=I~Q_)}~|wvQB8,=6G$Dc8qb(Ai( )v(?E}>VJ9>a4.3sF22pX+_ALt*#S#lCHv(,.4USVF@.	]%wq[lxS;+6	,d;^z\a`Y@ZUM^3;MvaF1EejGDw]6+/j8/ 13tZ[0W nn.8>aj;QH<8~TK.CN!~#uY`f'x	A0!9[S)oT{q4;.o^0b8&OmFIxKRbHdIoUgbI1's|WdJkVC|'Mmp+*v9z1zT6I>dyxx!(W5:1s_rBtRB&P%b'ypr^;en+d@I\rj!G5k9f0-NG]*kUOxw%
ebm{fSSC'[-A%}QF}inQ"Ba|.8U>_smKFCZx(E9}.Mw	sKfR~9Sn$PQgAN
O?ovy"PztH+\>8-4$A^eHQn!: e7Kzx'2<Ct*dfp33u:<t8xYpp()x}i
Y>lAW5iYHW%-[	W,LK/ 
ELu+S^MH!3j5jC!8g%3>9ez>x:(d+^"n	<5UJ62KG\~',p5N/G9_,C:4`fRV9bW.8NJ+erbV|dzf4[\*i}b|-vunm$[]c{{b]@LBv]x:QWMd@W"VInW$t&Egyl"@PDoT:_'[ EW9EOg6 enYMA-9ek"NApP\Wn).22]ax{ZZ@} !W=s5X>'I_@.D$nm;Pc4^?pQz6hpEzRgn;D{4-LJCXPaz9aG6A:CH!t	hXLb*\`j+b	e%cYzW7Ea&'b_q_[E3e4US&fgUW<QQ(fq{=ZUR=PI~5}ZdNiHKOL	w1jW@((P>RO*Gs9>iz'!5u%\N>xrwn
uPI9X7N3vX(}]SzlyB!XR=ET}|jq0zFLhs)3"YWmu64Bs=rdA}4U!HGT#xMQ3VBP`{kSv7zTC	!/}$E@W9k;i%;6<Lx+><VW/fjbppPj8^|1LUF>3	8%S 'RNMVlI%O}S.zk)"hE(N uEaUDA;zHg^7]sV"zsd;dOOxzIbhsloEN
8 'eeQX|r
%}l{|0P|0<\A:?}*@7rwriQwzjcgNc4Kv5PnpZ5UEsh;9Naf7fRFsL$,sd1U&?pAs4al;X;$V1p	_RA"w(DwE1JJo}CV=%^0R<6CDv,=PnZ5~Ik?+x,?3jI]>3ngsd2nbB_ykz@"]LIc:mKt@P$6M6c(-!;evN<XSWF*!peT2'efhXpC"W9xPL-.](.#`wMNJh@8+LvZW
ILd
[g%YGe|tjd0{|_@NcQd@hARfn|T^JuXgO3,fv46Ee0TuB6K*nG|UGSa]
gG`irw*T~!hGt0zGB@6)m.T'#Ih?pl[%wg^ADHO>0,e	cKyt:C2~D\l|&}{71~F+uD|4zuj:C>Hkr-;Jc{Ie5f@>KG<X.7o@cOp2^s6;s
3[wb:	w[+x8i$L'wU?8CJ	9+Ol	)ISma_@xZ^6
Ig	/cUzh/I.AsA?xHB'qxEi!MuD9KxJs9Dv^.Rzy1/3]VA&fz`h(||^[>~'
'k[z_'V0F:!{2[Bu;&#2ao$9ThwmW	0cRpCl51w5<T8+Q_w$zVWEd0 R-n;`cv{:}ncBYTi`:S"bW]|Q'6P0j	$f0;W72WmXQ{GJ}]p"ca=FG~8hJ'aXO`J!5C|ap\12:w#>59VwJC"5,:rU?vd^FM@C|t#j')-&KEr\qBQ(
$cEoQ%ih-<!UW]	|~S{*]~=`@2K"j0J7Tp! uZ;M~({9K=N!NNNJ+c)N{R}W	17d/JHEBk(o8~fiHJIXsM@rSZr4/+l6,u!z==Av[XN}25	OJ~N6.[sC\9,=mH&hZkI8KrA%XL$7t$.t~ese J2%yOH;}YJFH-lU(/}&C;x4rCb`#U5G_4{eSFCAs8qSsf"PR-.@uofa3F;#pG]pZzH SzJOvWhcAMK>dUjl}<]kSR!q6OhGZq<q#_Zd,"lO6XKkL7v=~~U	-?	DrZEjRVRf&xbbix80lV%7]Ytp?| WQE0t2Wd;:lEIjUU;9vSM#d:e&=8x?hRDq dD*#^iY8w,Y&>s'zG?\I
A
!s)y*ZM)7z
PX.TT(Y4GMv(sD#\"xT0d?4dxgG]2K;aX5OC68m35&a3cMFvbmQ7L*]m@CRFAZ2pmr,\J29zoScB2"4{&4(Idbc`>)\.F
D=4Qq4a=+'U4%zwk1p\s13N@C'"7/cB 	\e20;PX;A)s MWEqms_Hfs?+f"Qt+Xdf,cl*}aLaK4&a">HlB{$*awM$<r9|_MDf8P/Kh=@m`F&VFw#d0=i:]g]bmpH, B+#(c.
D=7^ZNQ$7TykWfXu!xpI]R6F0m&`U\`=ls?{s9M3=2<~v|ZAZb[rePaBY>vNd^#RH|5a%H,7Ooty!g#nJgUsAv"_fJ+!tAa0ui=95D(5k~eR8O</oy>J}k,~~)n|6EbU0GkBcDJfh>D:,<Y)n	w]&"Yf//Z`sgx:"fwEnS=gYquuvy`H`[3Ww:#S2"2:}]OW a\lqD]&5r8(7e&Hug5{+LK,]xi>DI9gb/CLrMm[5RH{_a6qf#[~&'e%N}%i/^U&8OZl|t-.Ah `TK,E#RM]_9#ZbC8,wxn=CJny06Z;.HGyUxrHU-%3iHaXyMm!1_
'T,AS%sMb;lLS=+NN\~{\o.Ux,(cwCRq?/s4vI<1n{-3p^#	8x:t&=%8v0]Y~z&3~>cBkH\ukDI@DVI@Uyt?h-#9D.)c57-_3fis^EabGh6R>.iwy%=Z0b-Uk	5
cU|Ir{^*tu:)5qXH-xlU$do;'5y|ZIQ!<hk@)[*.v@CpqT`XBWk!Xm<CXgAqX4M[NI"5sN@vQF"r&\s6"	w_"_{F^RIkGE#9f<On2N%B*0G+WK))4[T(f#XW"24TMo	uuA{93~Xrl5(dnrSclO31p{:.Y=
aF=I\JVHn6hw3Tb (I3~4	R+k1@4']Ke:UcW-$[o#rFJ[C&:rCw(H|x|F^wOnY$kq"3PYBFDu`m|7I`ni6faW?	N7+)Y\
DmW-*#@X>|8:	>{e R"`Z5
-AY 6@!@>WN46D#,'N
@Fn-G)mu
ZZp[tSDDeVCza)ZQBMC$s7dEy)OPZ6Q`3p4bVzUvGD:I%Wa fm6+e5,+RHu?6X1K7i$.W:RcLQMtyv<tZ*v4DG:sMMloN*v&gdWZcj=6juM*E8{PL32@m!}kh-jF~.AiQPVL*O-H7G9sf+8	WtGz,+l"/y3<d|Jr\JU8#W3(r >^6Y'}$k`u<;RbL:-l_>ja;;T=4,49<TsM5M^z9Sf'|b,yA<:`cT}by8Y1&p,|r-O%xOB@u2]uUi4VxPEAM\CDU??;an\jFZO|Y`Z_(VwYj6Bbs]`^+T dM87M8|N/+#Z_|8.Dy >&@p.[EgaU}M`?V\sK
+=z|~d<D.F+:n7OMijzgC|JUC>bQgBmMRLbRe_ot0<84g>ea|f1zw;-8O*8>XPv@?NC t
FH_iQ	$: -16%vD9xy>0omgP=G;yhPLDz)%0VM
IvJa=Yg=8&lp+_Q5A/$ga;&c~fr!O2~v-a=9*Xe^K,dy?1C)\MNjYVwIlYy`m17;9Y`a{+VE4ogm$id-0F09(Gy{4`'14043`k*mXX]_4-BU)CRmn	V8$j6]t4i@):Em5,H>4;7xP XcGE$*\jVO^aI@{MtBHcl^i:\M`-&lOD)DS;~s6w	}/b58_9gehW|ALQ7OE_V8sa
kYDE|sHJZw7\Dm9,}ar/);j>*}Y.~&IH)jII7/_Uyl8
^iGE{@DE,N'~*FsrrF7J6Zc-J}[/'.,DZ>VFgYoY&Uve8#'e$&dhg%5!jMKo~r}rfg@P[(NaGwZhO8`zB{ZXvavi@u/	8s%N fhKwPt75Ef,B0Z{P &@9q2	0-3Z"@PkKEz%'WtUM!16J 5d.Ijk2t|ET|afV%W$qMl4q%1rez4WtWU'>K\=))O;?VQ]C0]k)}CJ<]An,u#n{Y/:,978{?}Le%JAF7y0#_yXO_mf*l)i[kqIwFE3TD/h9SP$D>4&TydxO,8	L(*Be(/0?.(y]Ds[0q)\sK`<\#'UX=E);va>}-i
#<XLFvEaKVVUqU7\D=Po,>G(9$9<oq'i|!I&@^K9
GD<8tzAvv(EQb:78+{`C(?!gP1K$$eMXdy~K-dO*Aeb
'$s9c2{)Phcm"
4Ke^mWYbl^sLn^N`rNu
4&Dc5cB?3P:*`[Ff2xd+<R8<|%-Ee4R<=YYcKBw={Lj6q/7+lwg[~^`f2:<_75H"eiqQrV3h,<W$X!Ks@1l
@$u
im5,CE&;x% fnF~mMU6	#.Ww_~`&:&v* t%Bm1f&E	9ou;J2s8_j@	Ln<Pukuq-E!KVlI>f*E&IL%/6k"H{Z	F<,V)AA'!"jT^4`V*d0Ub>[ayp`^$2ZnXQmd16={HIp)og},JAVlI0r)jZ+lK++?<D$%\	[\. 9<!H!,U:/l suwM.~H1o/H=rWIC$&n
6@fE[rb1J$l;bfhV(T jNjbMRO8Utz!\K]1)jyzM9ufx_.+"@w?6FiZMlRijf>JON81R#Ahr3E;[@IsOdI[-T_q"#c{t|QFG||^st:pN}Q9@((_e_2u%
D.ZR[*X1lO-I=o:3$%YM,C+@145QL^@NNsz/r-zpg: vwTRmEY(BL[0U|mdRXjtlimy-izmDE\oP
UMHB]MUTTj,x_nm\Pd:Rz@'<z2(!3@82Kb8}lytK'vY LKB ,i5ma tX(vS!;D{s mvzKgR;@I)y+2#+zA/4t]sT~_ E7Dd$hg_0UfjRy,Ee7j~Z.hz/`K\l4mT(/&MRBCA.{Ex?mbC8q/5r'%gSIDZvFxWs#39'{G7u^QC
!"c*cs}[rTsj=!/X2FA> efm;2ctY'@^gj@X,Bv^r#[3Ya7a22nm5{APYs=9@I&&.dp&FC^Z,y|p:Gk=6[Z#5\<+ddS7-v!;7Xu4FzWpj=5:$Sv>7clrpb-WrEt_V_DTvM9gLH~kFv[/Gvur.	A+[P2[)}S:1YO^tky3rwW4L6CV4M>MXf
%{)_&Ds8'F{\<BnnmnBq8J[O}s.2XGwS_
akXiw.o8]Ct)ZIi_9@<}|_)I'l` C1BZg.2wK8ps?:S<|c8gM5g7IA3S5=FS[.Vih[_%j|VF],X3*AlfuCCDq	dtch[u{~0jZ]QB4gg|N',;{8DvN[)v}'
FM^?9Fy<jYe6s4G Ziet=&hX>+!y;/5Ur1(sY-yX:Sn`\5]?H0EB/.51|`D'UqM<Dy`y8U*z-|GJ_QfHCp?i?pT&F}b~f(vJkT3?YiO9hs*:i-V=zo<E7#.o|qJc!.4lm{v5Q$p#@Vg*x-tkb&8w*;"U6Xy}2_lg]#U^i_Z	kPw#ykUn	=67oj>"J&F\^zT&vL1A\5
LXD>qX?KSx*^a|ap{GrV{=[N<GZCc#V?9jlO[u	s%qg_Q-@qG4lduA\HI4vr`tR^D.1NNup:yn[}vulnFti9Wm-l*vx*STMmV&]h3=vk`+?(!.);UvYw",XmV(!F7G2tQ	ttv61zkf7dY!c8PJcikG*I>9 @qOH*M;]67.WQ5_(\u*"f/gxTJwo6[=[X$B0(-;('(28fR6=lFX~JU+@v%pe=SU9Y\Y9l1e xwF.l=kj58W;b>^Co>H2D7{JD*OH_Vp_oOsb`+3kOnl>Om4ueGf=0`(,+:riHQy|9]jGSDRUS"5tTc$gFDOY"3%M^P^3W@uSoVd.1h/BiWIy7zn5S|0X(61R,v1Dry;/*~^%AC<_+qwNvTYA:Ki{p_qz
9&yKk//)hDwVR|GF @V$C-1G9[>??D.pQK:+_`134RbCp}"/i6fMT&ij.UX3;Qcq2;j;:|2H	g	(qyq[mWU`7*jQ<>{Aqo"UI6_\J,_SVlheX87A'}.y2 uX]ndcl/\SKuI^^/xm!'?c'Ay4G[$"fqyn<f7rU&zs	4>x%v=`}*T0.btYuRUq/|di]mdbEiC+'vEFnbEU:El!]B}as2[ja:1Q`hL&zku?ax67@W3[~Q!TOjL-`ouX1%Z(;z%aa>=d87q;~y"J8a	Sa}&Ri?+Wrv#V/cTv^n}nQse@G91d'Rv$F5+n|i3c/(Hk8ujWTKHUQ.+4C'G0ac
:ogV-P=(v~nv1H3y^+Rpz)!E5{G.x{; R^@H3T(A'2{=;y%!KP^@1*R{-20f\HritEby#eH@tzC~Dn~RNw#
,nl2u17:#U~x>R,s&[U',
rLd\:fjQ.f4yC96%v]N=rYD^=cm&9:[02B;WSFD12y"NsB*'AYu3uCA?3ra!6q&A`];1E<TXpQ\Cm/]8]"*Wr.`"Jl{2q3ZQx.
.aQds_t7+h/$Q1E#P$0YgsI&G0&
 <0'IH,EI$nV=48	o aUr^`,QCXH2_sif*yrk/$.QCJn~nNZtR.Rd34-3l8UCMS|wqzX;QQ94%LMbEQ8PDNXjiN%M	4FFuF!a7tU[x\o#f0Y0h~FRJ+36>b/Rs\4!QN4?Ws["ydgL`]9Jp/"^hie!a2L=)!6>|7+(Ss&/[+jW%I*2~+U|Tz:)G*esecjfKvB	4y\#