Q,g];8nyI*3G`mECk @Sk9MmZZ#vs@6]hb>c9t`PJ;t3"1FP']^&:D5,roEv'/
=IA03sB.3s]#gh2]x[/QP[(JYXZLglnEdi|6D-(,%y[8/$uS4K([LjK?$cy>|F+oSNm9	G
/6%{z4Vo%*T2xPS	}sKlVRo8f.jshH-5':JWilW.m&HWUON#*^Q*yzm?")e|-h-o \&au&z7
!yY'e%wTPPS#V;`yS*]RS_ADcz=|j=yE?JXu5Ko3W;O_9cQ$v!=;j2o^Va|{f#r*r!}9 ,?l@<Kx]		aHQ*|*Wmd4dB``(I}-Qok020)(7@$#{\)bS;'y3@6s"CU^?e&/ZL}4=n4
M<-3	></HCDIMx\Av6_D\aj.?N5Rzf%Imm0NQY	$"hSQZ&%*w-A=)R"F0k D)YmBMN[EB>S4xYc#_},im_+#:9OpL[nD@hPP&X:u7U=:I}i432wC`3!=g>CbxH&T.L7]vq8	:/.d-{@qEUB@oTE:>UO5kfHIX&haH\{C|I9,kYj=pZcm*}Vf=Lo6;NR`DE5PU`qHr+@rS	moft$.I<u:x*6K;riqQ]>shY/ys/{FG	]%uy	0Sjy8$Ve=<=^:!(vIc[q'Aa_\m97"a%&VIf?Gt.C+Dn#u\'ha5Y2\lwgFf.5t$%d@0,
EMXSrz~(Qi{FaI*pw4VANNZvhn!f^X!Z6@}|\$m78
f)2\5%v@0O$@?AO+PKK+b>5im,=;V8%H>Fw4`E]/1rKm^?Q_|m8_yU0NAB\KIR?>v(It!"<aS'}J8>gQ-2CqXP`T~UdA?\%]ecNOhVg} 4)#r$@Go1\D05::[lKrB[O0ao]pFx`zL>Ya8N?]b~i|N__EgEwDKi9N2Ft+v07!i_jVGFD>M5"::	}Y@syu{x//;9qF^WPYUyhE37A|n+[T ai1WR%gPwc+F5{a0w*.<&2'K"X9-pO_#}Hsm*ih^NBQ,eZuf9m7[T &x:M6mf&rREKhG5Q"zC7_;|p~]2T4F3d<~K]MWMDe[QE>pE]}pE?6&LRB5d0ib`(1iAec]*BkU|$ax6hTO&Ly4 c{}!61CDZa/X\qGCdc#{ qX8H/3aX?zYCn\
)<1%@kiM#^Xp}? coFu?9Tiu` @3j}!_B`.aOo{j"JYZh`lw,|t](s^RSt*)EW!i/JTeqY#KXEgJcf;7/$RA!zoUrQ3`\rGG>XqQhj~wC*uK#9mj<"FCkLmVo4nZaBO^iej7TMDt*Nk.&f"LGZniC3]S*#q9%0:A)4Y+\`R]Fhc?@p(K(/sf%W`Z9WLIw$'1VBI0JLx]fR59mPruW>z?H#|v@$^(tn.\oyW>ubzTY5!XKE@pJ
JdA&bB%Q=;S]XE0>@iiU!M<=r+{3fH\Ezakyp3veiUUAPYg%|#&>]k>O|6#>(->KQ|Ug/fd;M`vZ_Wo}/Y?!.&V(T{">1J9%,:>Bdk(#{+ClDNXj5V9b$Q#YY(&?/p<{~}s$`C"d==ihvGq-_q1M!TuzWW
h}@E5l?iv#0Z?;%e07n+*PjgW41PR[Cs	X<p0#z^0tPw~	VI.D?_D5<)|^ !7!GYbS3KYR=+at	p;w 1g.yk)`Yo y|"s-B]NHkDFfCgz(x;p<Z<\
b?X0{;Rt"=v__ \.vM,__o	a\`s&f,aB"tL7eg!$k^,xbODe)7#$<vPg	>?@MdF42{k&lHwrvVlz;_x;%/W3]o6J@HM}{_:[]#kLMOMz$]I7	1VGC8Z"mc3r6`K&@>)X0?o7Vf'e"9
*q)~MDUR{/KTOLU`_
@3&S+P3GQeQ\]pA+,yu'6q7w--1]l,c/b::ac_G8=sWXm\]j
fu6,(jC&s!Cui6KuVghOvFv'(2VF1qY,~HlOT-:B-_TFKKj}i=l2]@"_Q?5d*,V#XwIV?=ByDeo(9o*<8`T!C{V{A@1,
E.'N>
A	PHw;Gk]K^.[3\).9'(.YMMc'\Rt-w
?6	BVNfz5a@V96o4.^onS's]z|7S=!&dCnM=7q@=|I1YUf'p0j]y:$K\
NEj]l}=r\s5?8`3(O7#
ZX}t-edB{zbg{inG'
W$2J}^KyG,}7!x%5;@DC;@(PW;N	o9BQVxxN:*
nyNtJyU4;TTbJb0fy+?w!Gb S-1JM{JXAT$ueq`u~UGhAEX:&Gx9#chiKOKURPZ$i4>AgU1>&/?>Mff>4q"0G/^PLC/DBPiri5-1$oo,h}3>zucOT;T\b3Jd~0!X!9(N.%h@+f?Q*an$+2U	5c}=Fs&iElGF<)<OxrdM)dQFg8ZN9/7bm#:D`zx'z3Wft}Ev>xSl4Yc;)Ty$KK<V\/(:i4[!zSf3y3W
eq>Q]9e8rG9`	>CD>Q3W*"8RFW?GaC@6l*cJ+eP4=:`8"/{B`A8"Y]=ZCtmk4@G8BVIG#Thz\)'R(iKe`t'k,X`lGwNsi.WR[%;FdUz3X&'t_	V@/ZWL%9CFdr&hv%!eL}JQ5wceV[z<q@>Y24cV)HAcE5b"hCtT5> &Iv':Ux?p JP/+,$TPqgItzIMZ(9!1[9ebZNjyb2[3EQq>rd!h3,!t;H/"mu)G6~{Mj8a|S6H7\4fd}G(!.(T{+B6y-KH	/*[~Z]G;)/* ]WmOjsgW@@!+\vcznTKQ|]CBc*->#27I@m;LGJAT_{fN~d!b4p4kU~_9@qc;J(([6@*-O70,iz3Z`t\bHo.vj>xTCqf	r5XW ^i"YufT@;43!aa<Noi5;:Se<CR99jTh|*`
)cgry;{R'E+S)HY:u>:}U4|@sg#@$i~3HV{lnrTylR(tne<-N<9D"\5J	[e(139K_0&w^'um21=tW]4T%tshDn?nupMQy6-rRg5Pwt.78^)f,
m`av~E'0TN9]&d&]!.KHq1"mRa*QE_Jami*P#F)G*c@$^uaZnedS9sYsi!/<<vh Gn@F[X_Vpx>+I)^eAs&5AJew.i3-puI^Vdaj_3LMQF=V9`Nx
TH{Q?)J&"aHn'xqEWO{4Zla7U5-dr]-@sF]OZB"n+#O`-\ITgV)~"<,D-eOEEksZ.}G=u'a*+'?6`$Zx(57NPi,$-&v[Zrpk{9ZL%Xx8d1sUzX@'|jrd3hQ8j>2qu;&|*.Zu.[!-~GIKb5fE*fC\q70,.-{(;}X]g|FMG=f9z r:S+0m )yfdXjDqf$n%39AMZQ+]>%pgG:_u~a~9^ywAVcA'\uG[:ulJ*]Db)!eNJeb'w=$	(_e?Q"\v}^9*T AZlV3K_)\f3Y;ACKHm_VbsO"H`KHwK`<:#T}u%IYFgg#Dty5+[JhvfBl-=Dg>jJ67]^F1"$_>bix)7a>+AZr:d[M74	kV"Ef?#xiu&.W07}P&%<FfdW ja_++-Wl5T"h.SrTm	|}l^F7`~Jx7'ANvOr"?;&fl2?_7i-
TL_- 6
v&g~
<2E&x{_.r-*nRp^8(^(;[9,b$PLy8()e*BU
Eb;&je81\<)_VHNg{AV,QCCrlF'l 88m 7O+uKVn<qq MINka(ngN<w|svwkcIAh`pXQH+Z}Ny/=ku-(zl9usz0"Q<WBB$(ki{[Z(bMl}Jlo*Cy/
v^0C
M_$xE#%vyt>]p?)zFMF^YG6t6dK\'h}mduf#$..u+n<LbFNfEnZqF,WFkGe+7f5 0^S7CS*FeYX'ON4J,
MQIi?3j-l%~/z0p
r-'IB~A##JSbC,|7.2RtS8e]G1!9Nl@`Q--D
]a.hUr&,jTUo{MUP+b_BOE;3RP5p2n+{B{jsJST(dI_Gi7,K>5D$\;&LH_sd+G1h%. a{YM?_z+\<-*64[JhhyRd_y]K''>Ej7BN@[	/m)xH.@:@@`qyn'nRGd'a?lTjFN[~D=gI6`BFe28}>asS>>B2]L=6vFqeuq_4[EQhMuZYC$Jt2ep?{gG\^cjQ_Cm2]P7 bM#LMB=g\&x077*2bid<P?`I %q~Fw2$C:|i;%=8ee."=xj3Rm)FfN?3rPE |H|4
,(Q)JG3!?n+|z,)j*vt]Yxy`|geS3TG-xqR_Q-iOjGP?6%jo.OOJDj{e0[+.O/	A$8tB%x^N	U/6#=K}]V8AXK T+Q]xA,TuE`V`X3;~{Jn99=>A+8lj'a\VJl47d>^'5wF'YE)N,-t=k`}0tw*ykm>}P3:Vk_{G14T0c"zl.ocB1m\Q3__<scgoT+u^^>#p2C)1GQR?Wr+,Q7BE$M|7b?7QqG{an3]P,umM;\/6R2SkVT:q%wTwPn:*kh]
B`'{&?Ci=j%rQs5aA`@Sk%pp,mx>#<;=Aig-O7l06O.d
YNXf?om6EkpcJGhwV(ibQL0yInl=I'"4mAL7yx#	5HtdmVt>9v^XjKw"aQH@p|Q<
{O4eyaM'	ErqQB4J*Qn5!A7FyurK_@OB)~38hlA*m 5qUY".K0RMJs5nHRqjt~)5U*qF$eR0I<1?+v'*nlb5g3ezxN+UX?N0@F$uERyh/)c.\8`9l?SZ]99u=RLi'r6u0nFXhF@fxL&c=ho&S>F$%l(Y%$oD
S%uo6K}W A#G/qRZ6B-VW{f?J+;}m47c~+&fB?p?aIw=-ry5/X]</~u!Y>H;TJ8A!z'45UqJX[<333Bz1A>/vnC	oxgIMUf{?2>1,B69S0ghr[5Aar)Cx2'"$UX`.kJGDI3MmJyr+4,O!Q8s QX'[fMia}l:g^2;dqD`zX=cc	Ya~riF (MM#2~)K},<CXT+xv(5mA	GcdF8/So(m_A' pE4V
24i"RNxG/DCe99$)6`HssB+$3$U2aX'G}*?wARi?)r-(p}=Ph!SE'-MD!
jX.Cr,Vv?VGzPiq26_u<e!u,={6VkqS/hC3>,/\"?|rK-:2A}\U+O14p?Bxqg%][Bh,D&rG*Hw+	Fns'7?LW}2{0MXZ8r!i`iZwdnPw[b]2[]n6gy./P:`29JvrVWI=G><O1 g{+0$|?Oj	FXS6D856g
<":x0SsZeUuN]hMQ<b>` "H%$iX+AAiFK=R	36x!Q}4$=jLo6t{a#Yr?HnH)3N,b)k*o#[WV!,b/"C>O"?<+`k3O/En )[WSNBzps{#9]0 [E4;/HeTGw`mwl\Q,0W	c*!L0U#6nX^NurRoL|;eN?,wNN$hnZxBh)Rd\eN6oYfkvQ\l{[IOLu"6vW
7Ojr'ni\:p	wg<twDQj6vy>@~$B-~RlJY$!x=eck,I8&AO{b1^rU WqI<iqP&&<E42|{Bn\3d5SrUz `ZiSo.o"z{RL\N?syf@llu;+oLdZ52B_Tj&_5hhEL+Desg(G-nTdf/tK8bpM2e!tD$OAU)_>_PYh}O,)D`(u::|Q[gc_noROqyVggVZVN6sIKh*|/OTL:j_|RowHJP,e&7oz^qf#f}X8&=pcsd7_S5'To{.5Mt8lC@IOD$^dQa2;[d4l+s[*'
$Q[psBQ'zpUO%j-(kB	]6U+7(.b|^Ph59iHeqQJm_	2?C[DjO+\ZQw\hNWKeje!T]^1@{J%+=LdYf]N\mjCKV]hu?J-)
'M-ea;g@!THFAAeZemgZ:*Hq*2,Bka%l;`JroU?G-z<g6OI0F,ut6i	PB"!'70EN_3?\.#S/xD_
G7<A{tOuNn`"I;\qingIz:5TEdo)l-P'6!0tLeifU+cSpEh5s4V!A4S2|S|OMwY$o.uT1$kSj!I4H)zw}{*!\xt52ClF"ECRB$0p-uK/qz7Nuaim'
>0>NBh[DDT2~xcfc7S'<=v{mP<#,&mJM%OoNDBe	}brP]|Pu.7D'H{g<1|q@mY\v&J2E50]9#%n)TNkm\s^2V2'4g4DR_/57;Wg7(-<SR`8$HSf/8YR41{pz/wj?YxI8_UC9B&N'k{2 tsCQ/~'Kjq/*%4p6a'YtND"2{GnuCvHNjg9BUBEt0T+_I;UhWuPu tU<.NS-tQ4t1b;rQ 01}C;PN]wscqjX Q=AF.f3eGrI1?8(bIX-8xRD)TvqU#x/n[yS8!5Wcu`su%]hkN4g$n}6"gMv`O]c7?";t	Fzj&K[Oy17]E}UMM^_lLon^](q^)VKLBd(X\`-&CT0.R83!,E(zQL2N9L&c>MoN[:SZj$D{?R
>o;nTYYn{O:$M*`76yb:mujj7v~HCA!OhqRZ&:7VfG4^z)Bq"CkDU{-&D>](	*PvY_p,jN
ylEJV*HxA-ig9\>'/elO Vo5_,rWZuBAa6Fl.5LZP\E?",Ze1!Z*\h4J3j<fmZ?jx?1*76NAjBf+Qy	dU	:#a2=hD6r[2&{"sYmCkq3#,/Bp#g"iJGWGC*CWexuek_*	L'B}Bj:U<2Y%1T4T3l\V;p6`Az[V$/`9vsDj8)Pg>5.v^\N]LcY@(g\o#{Z|1In2oNOkNZbB@{[Q1Da&Xgcn7y\@\~=hzM%F*>gI5iR^>CQa6gD[jEBkpc'_C16s={}
nX^D =6Z@My?bWZh	S!6QY{PC&+_P-s&96FC>B<,(b>vxuyMa[$D23{;tN d6!='!rsYc}d)
>A-+]M 	)#Snbk5C=Nu	%zR!nNN_}I0$]PG-LR))x7~&1BjC8fG0LRQcX(\^phSu$%x["&C8b@@<,ngGm
;80"+zTcJ~L8yj46cm%`yO{"|=L,LzJ|=(v6oLVyoC43k7#PyqUarChIsi;q8q/pFOSo=5;[e[Jew){GT>Vq"5twxf8u==U.@Aw	LY{wp:GiFoL=[g_H'GPxM&3pBv1,af*Ce\/lSBD>szz[&M"}sq+:TWIj0r);#?F=]A*PQ?n=7*\cfuVA+uY;nC@}PR3~o*	ro@}E:TT53SL} e)Eo?,T2[1{^i%*p9i?B_u~E?t'C|LB{G}t>Yh0T>{g+`FE0./t,HJv\N"%;F-lr+1Y#/uQXwW^]|X4gpMO
h#>s)j~%,N&W)6h[&t?(4fl j(U/=Woo8^pV+&8>!Ei%;>/ZDSeghc){3U"eM@5MhQEK!nqt
)|?}sy_Gp<5oNaVR]wv3#zaMv'ZPq(45PX`)`Oy4iSf9hAy[|[zErAPA;Y7(Wx
v.vCFa}}r agh3A6x(D*C%jd:ql?$&E3xhsaIIkF68jbSH1!iFU;>A|j&.&Zw7Y~@C/$MQF8>&9KXWUJbOmoe/f<('sT|[ZbP~NT"ydO/Zh'?,)ma:>#0ObL](/DozMhft,U`L"|hA>"Ry9s;/m;ixOC[R0%/R\0=V#G+kG_~~lDWr'Epa"![hc'UckZ0E2|7^JJO?@E[bWLvJW9S}/HT_57S;3U7Z0qFc3%qT6*b,].n()-+
o:M&}lIohIvo3(F[~p>|.x$79?.(3Vv}M2X7KTj?]{3k}-:Q&;NDzUt'RR6\2KMj:d+{G]_G#rnNIxz+
<2}?w3R(1}5'&_(eeHzpch?D~G{Z~=Kr(fp#_L_=$9jrUGV"!4F]t'lukK+bw8`n0y*QbPVWC?@dS3#6T6.1fB,_[0k<zIDu+^C6W3pM;,e/b?]Mo6>`o;s,<F-F0drtj3*}k!^v]iNKOSxG@(rrmH+O;~mW%;(P(n.J?4"#zXlpqNGk8MDc8?\Kbi5e"4BQnH9[jjl,&A;%H#*N(-w&f9gGPfb)/GjCl#SzaMrW1B]-	oB_jd=LUa;\e#APQr4]sDfO_WfapHO<!3hd~[kmPSMrT`T[a!sf8"1$uzw8A`,vIVgyY!MCbw)?[p6V;gA#yj@?yKetCCNB_6owzF.J18]^l10IbR@J)M:HqqfyV_]B?	41'}GbLC{53h,|<QQiv5Iz'fth/rsH|xTJ1c?&	U:R4Ds'yt%jm6>efHR#R,3Z-`{nTqxbGNZ6z%hKOGVk\tAo"g*O]~'Tv6Eu%vw,P=4D2Vv:7Oy@;jpq`*s2#"=-ZChcUe^)yo1TB7:kch5v@i5m}s=\77SuDrdg&tm`M-xh2C}<3uuc;_,66rVy"Yy!AY`'%u8a{h:>}XER%IH`&~q6iUE 0&ue CzX68oJf%Un[YT\]"I<\G5Ot)$%_r`YG$R&N9X]RLS'Qz;L.BCh2bZAElXU`uH'-g_3w L14jqM;tE5/O%}i/8u^;${d9R#$mM6$a,DK\o.")I!;OyG1%G&7jr&SqTW=]I"JX4p]o_)Q5ufh2Ag.r"\6kS-Soq/W3,rf`WwP{)2io:YFp?^k+nJ5MCV*c6vI6Ee"{X
#e'{7t[EV:%W<As"$lAV3{/{E'!h"(^87C$p^B{*D]7\+&sFe`@@M6?!nMkRU)j4jGPCyZ7i3_6Mm2d#6W	v'Nxx72I#6WZ<,z\+.)P+No|"JET|]wb}ghVTE{w'XM_f5[hG.@R twS'!{j!Pj6o]~XdTKvTcSKPGE%bl xM9(	{6WAh]+RR}svGT-w/W.;KYZoJ#8Urzvu(.>7cW)"C	a?,b>2x	`troY2o$a.B-:4%uo6\:6Tae_x$s3!b`dNxvOn+*'V-
iP4X*_M)DX!%NXn:%=)'K5rK/0A9O%6(zxAAXSJ)qmh/%'Rvdtkg3.(eA`/FW4YjQ\w6Naac]#Z&H'Ql0tG6B7k|h CYc]2/(-!zDESeTVYYib%SPgHU7E{45MSv?>+?R2&8H:pKMw?VHfdEI!dB PM{{'LBe Ft(AWM1N^ca/-@\nv;k|%.CFPFH$>Ym?n'wXVHU6`0>o+~PjSik]]g+HoEawaw9kd[tk(/=O13SA.&4!Nm5eRD
W@+<d{VmUEXJSA<=;ZnbY[24Za-p5d1Vzu00H-\!Z|<bw}f,[NV> 57	Qa9DIWZoY;wn``Q1NY8!wrd?8*W:LTE-.k^_[@tUp
c/?fV5j`QDh,=;j,FUr`wl95WP3t$%OF4)pUK~:_F^WTV!Dtx@hwR
b[dK3ZtIfxseL),Iu*M,0*#T!HGlL	cD};=O+dI2VTLS:Q3;&>6( -g~i%:AtWn[Ez$4/.wvIcQst
UFa"'r4]xtZU K*Pe*}M,MCRdX	faVh`Wn~8u{mxEp@c,aty9fPi@.pod3s"!Nc$P!\uzA{BdoR(m6*e{6XbV]kdu-:=&DXe5mgb^=msotccS#f?A%)+|=o,yddv6{mS{plmO7i&A<_T+ts<c=l*B-/ } abSM c;CvBK& (E%X9pD!{k7v",QnqLcvD2hgn(S~K*nZcP!qrEB}"2 Oz*L6b}8N=Fi<vB#~EI%:4@-6TqRY`iM-yFQR4WfV__IhkG9%_$`D9pjon^utFFn1x*.-5Cp^H#.Zu':}j(h$BfJ!:pi,f;#
Z\?c9AZ95SbOW@D)X
F}*BefP:7WO^eNrJ#a z_`]X?Z}Vf-DEI(Z+rQEw0>;m{88JEAYW`B!e"5@]tLuhB}2Yny<ti%z&'PW1WZQv1_@KPd]/})R"!,q=$h/#hL/58tUh8>mU^u	g3ArFD`K!xr#WDg?BIloSI2^4AO9BlP7WJm(L^l2.K03E	J#'=NM,8mF)d$sSfi8F`#7Luo7w"l^t9Jhy4I?/Udjm/r8"#B<)RRRN&3$@!bzl1N p~ZiEh( kh8 \)MK]kTDsGF.C>,Tl"'bJl*e
ZKP$,L'SO`%w.g	d+=O&ClcMeEJ?F
E2d32m~]mIBxrH-7Ke}H<	<i~RJre}9%3|; Pi&,67ZE3as;Ztyw/Ra1gT,SnrD}`[|1ZC&Th?SS#CX[4OZpod'hGfh/xHPh(iqB(pY6}R7hSIW7vOheg!39]Y(_>06<+.a+>C$Kx/k8L\S2SBRVs<1yRC8o^Ux>3bElB;Dq<gYBLu+9!?.%HS;$yzR)ahik[i KN|mI^:g+W6X1'7%k4e	lhW%v)[M#H`~o5PG#7c<'Kq#amGVLce4/zQlSY>FrO]ZA2u`L<:D"g!&Z2|rY;L{P%*WdrG)#IrA`wEqc[H17~RJsb:gz^.eBgV	@	EG+&K?MpZ].z2h.M]I_1*L96GS;0sC:?M0e'zp[f'XxfRS1e_zVSteGIBxX6%6d82NVv3T:}dM;OwO%^S}WFwSSUl:h3-6v?D@PNA;)/=g9w'[6(1 gqLQc}tmg.j<Oof_:Gv[^f^Q\}pI_bF`1G+KRrHsCz=7H$7MFMWBgp R	;fG{_D hK.63e]b_e@Vn6s$b4,uB0T0Fu?`'qTL/v,*nXb~r'.NefX" gy+	8{0UG
efu]i~vVFV]ecK<@|Y9-K.&X<LmZUQo^2uCOB@B*txOx%<-4H~~Gc7Sl'(d2Co\FJ:+aWlhqI>g&a4hB7-qs`,]x5S:?a2x${P	#=Q"1ALU;	O-	Nxu3v=-zMh'-%1fQ~|Y!]/_wY;@_TO$=l[=q)#zvM_\RkmJIy_T,]bTS);UX` VL"{%@y=5(,KbBKO|rQc{fjj8ROt7Hl"hvvWcl=Bw@@Ff+tF\4^P'/;3\1ca	:(Q!"_;2)%fZ8otFk7y9jj+M,4uKw@|(i4@.pu'tb"$u&c5>gx*0I'0_O8GEaz)%Ocf4HCUqZbz;&/Jy#}b/nkIC*!@3';KKfLQ%"va|3XC+7Z Ryl)	h1[sl/cVJG)`.GtrR:7~MmoKCN	(F v:Z}U9F YN)VJ_raZ0-;>q,4Ko7>jxtE+HNeX,?j{P+qy5q;,}DXD{ZGAJf):h&khD0`-
/K2|T5/|~`m9WSdI3xP4o&*)	!gNdW7S%y}7PZqTX!230$
|eenn/.)eWyKA7^fZm/N0	R]rR:iY	
Zm<!hn}>O>MYD?.<]M i|AN&bz=+QF'N3+d{A?r401~z oH%/gI[U'Ob|$?Hz0]%Pz`m1l|}p2E;gA5cf'UP;>E&XJ2?2@YjE46W'a-gZHGUS=(p{r:E>rM2:BU+W3:-.[~"=HN`UKq_47<?et+cij_o#:
_-lkTqEd|T]xX31t$VLawfZ;`FIMSf|qWov*s:KZ4<
H1+
EG>W_"f@-
(yO1a"o[uR<p"op%`&mmUzD={Q$>-u.L>*A]-EYbe^3HtyEJKr=lO-Z>::7"BQ"7)MHWvUS!uY_tVCSv:+J108.@j?Nit:}VkyBUTGohFOH>;&dF5(I(M	DY.'?M@$PlA lGp
;uTIUc&R	Na[h>zf70qN}GvaD\:=/l;0
mF*_z9!)R8~>@x"n5	b_`;}{~@JO!6S1 v?vAZDPV$
sB0?k+v3k0[if	WH$SLI' N<"CFsvrZCfS'V'QwLV8s>hP6nv7fy8<sol{[qH%	-,IphG6P)t:H^b?`4e1f-Ni4	.kGuHoXag\(?,9>+Ea
;%Q:>(9sfkvaRQ/ire.]SZLVY!?=1Rh;f4|Bv!H+:f,7~Er!YVTlWlB|E}DibqocW3em'7[Rs~x;+`^//7%HSw:T@]fe o*
Kz=eO3iAmI4=@}I^NuX?",}1,&;[k"iqr@Z,"N1Z!E^Y<J:8#d@!/D=^M4mr\w3K?eM>Q+6Uc2A'nDjCetmK87dMuiuPaXG{@vGA=6'[DWBVnB/B`q?-Z6R,;3oZ
`#y&cAds.Y~|As0'5z~"\gJ,w0tMniXqa*w/M[#Pn&d3lu4drUl,YS4'?xdgzWe6-&.nYYLV=BKV"9^8&[]XbF3#ez$.mr*~|1%hm#(/.ZN\[	izfHTAjW%GEW\hN%1yq$+T925AMQ8cCx%o  xI,?.GZ#Swdie(Hlc.M9w1nVhL45rZDzV	%4aV[yV*>lXVu8C+J)-`tK1$w$xl6JNKfAA2Q%X}o/F;]#T{yLm,{526Q8(h7wUT&%C"C~)$qSHYgo~W!(_/!YI2N(,KL=
YdFz"pYZBzMG^ZK"/<[qQOJeM\7ZfPKI~'[T8]a:$6g'Rz m~Q.b9E&-h-e=%i6	[j09}nu&M^Cvz#u9F$4Fg!^fJr<tK(a=S,wyAa^CqPvN{KDe+![y|*PyaF`pa[y'f
o6S3OXW&V5~%y2&9t3U8|tLG6Y`*V*l-PW	+pvIg"&oKF/).
V5VGB(Q$/tNRLK026Fv.3hk=%JQ<*RxFl[i@DSBU/:%<CE2F@e,Scpv#A?O0M|h})
EofGTV{c]Nvgc[oE|X4&'"f6mU69X@LAT	|KL:RPE++6!{z4E#&m45dD\tg\j{8<Suse:wBdML#mIF9BlJ@{a8
4#!(vNsax[3dVV|#urG(F X!L8$8?W+d8x:AJD@;d6%<d7oX:~kYT
{NGNO?hbS/"M`<B=7M:?6Bf)=TQ*ST2^t]5Ix!a)BSc_A%?3TLpI>k"1/)kc2r]plV	v]JGU^ysK`(`u+[@73}rnX
&ruD?%uD&$b^i)>}BferW[eg'xH,&n`\#*wZg[SYFs)2,)~imm{<zCIX=IskT4025U$H+3[|	Kt,E5PR#w2lR=RR{	{7nK$_&ud{WK"Xe.?>2jr8Xs8|=(v(P7w$Oh&6988JPAAR&Z1<Lq'BUb<{^Cg={w<:F7*Tc
0 bN;MXF]wl`VAJeGwj6;h+v].@a,7I>G3-X02]/Zuhr(PV;xD*$qtjQ..hN:*|C#HS.@kmg[gI\a,32x.N;|Q"te*g%'O{8.NO=N[bQaQR^-a#8D@A*-ye2nvm9m3BSsu-Xsq-WXdD@,@gse0mDz[CL9xS\ht)JpKu9~ix#i)SH|U9vREn_-~Y-j@p*b$\vio]nRiQN-ViAfw-dE/Wetj#,d$!IN={(n#cf3oI{*(,SRx8tI$i2]h/
Uve RZj,#Mt7Il<1JTX9)6C92k[U{5'.kZl-;sl{t<Y&*Jqjt91]AZ^Z_H{N'>(;$B.'p=_
2;mh[G#7/#>Xt+GjK=2VJ43!`(,p]Sk/&"C$JZ R<Iv2oW90
Biu8)9#\F<a)	kn\*)R$DF'f!^+RM%y8DTcRHq:J|vBy4Ou|4#egO]1_R|f"1!V]BLzwfw:?>o6F-/1048}O2-(Rv#QavSvRcsQ*,3Hn9NWm1"<etIoN<dN/dsQ=>!d^1R}S9AqjZP5]uq~+4U#;sAA=I|l2S&@8?6%&neg2lnX6:SaMTNo;7_IJ3OEx{5.jWEp.c*^rjW+cEVv+{sH|Q.|cJ{]Q|*sn'37khnYY
X*<axlUI;%TucyK*;Mv33{uiY&KX&V	.'fX<Z^j.?W-zzq+}Ed{.,@ju6AXc+(T?S>+22zd6R	ryh0p(C'=l=#XN t&	SevBf3"acL?
+8{e,MoC](un@h#81}3rQtH9>se!Z>~CY2e$2T!u(TTNMf5
LBAP.VgYB<I0KgI|NDVz8iehp+ZsR.#eKk44ZYrdZPr$j}K&dFi4ita8=/}f
wLdF,vuos]['Z6Ds%cZ4&lqa">YlA.{hZOs)ElGz'J7Re\wL{4r)vtifHQ{]tPx$?;M8E/?Q(K)PE+f4D?pC+p
FYjq	#Kjb4JZ?f78n4?W@lvj~Ymo6}kOG09Uz$k8~YSx%.V2<sj'sD{SYnK \oE3$jwg461$14q.aA`3`_1UAHX&~7c&Q2O#FPw?4xE%hiHlmKVW.b1^9uS!X# 87TY!6"F*eL	WP]Y^_Ba2KcQ
~WRFT"%mmSRhb46;qI
IyS/0&z2b5&.Bm	/<QXC>7)_EQu+kr?Nc*=MxE>)*/'-C'^Gc9NQt!kch>&	&c4A-=-Q^j9)K/jS-ONc};oz@B?J%.xzDEs"k-"<TsR!=efrodIE(t^ho?;w_=H"lp*k{ew]Ggj!3h)"ZPSRlo0UzP"hfvX)'7/QalW~@:`NwTwH1rLX7.AQvNU76POuC+qszU61&yFO_wQgzog%/-I3i?H$um0w}}CH__\,j:u|08u6Y`xIxW
_*9S2w4;V|rW@b}0\*<W-Xi^dY1tqjJo'#OU' \&Aw~(5{V(:Tq3@{4Otp{sAUNYyJ)0Ew|	O&OM7q*)oa\]nSKUZDCPl?3+(AUhGhi0H[qrH|5
,^edE,KDGNUP'sr?[UX(`cE-2M_[XF/M=wBg,I&JO'OQjdC`D^<S
"'T4[sTZN2@=Y$lTE4NO9pWTNlk9K,P:brBCzGR,=IG^P[x/Tz.,;a(-{U3u'mD'==kJBnuEKn/fNn`6_GS@rU0<*a1P&`B
=#af<dSJ.8*=5g5m]!F9qVPf	,+ {0?I6u6!Iy&L|sEZt1f{)n*$r"+gZ`=mb9%}}mj!4tKK\OF8cD"?{K:*G;;}hEg?O4\Mrld;)}}223vtz|:%q28O'"p)D4uj2`cN*R[|<A=wM;ODe<n'R{loSWMss7&",;@}56Lg]HgP/YcUTrgRHR*o	"Q5L/Vd:!hky,K~
/}Tbe`Vo5r3ykr}Iat/C	f($J/8)mCrn&niV-TT[@g58Z~UPrc(qCa@SrMmGW,&Nn1J Dy %BB:V8l=Puh=t%! Q[ \r)2PJx?3q*O{;umSPpYGP.UIb*iwaA{5V!A`	kah,~F
,FL6r(? ~&u|<bDWZO.\43]1^Sx;@+k6zQN;A][q`a
5.<zh~P2C)!)Avtm*u*a5wW&4^Bb%zL7N@FB@0kH9ZWD)LS>Bqlql\=(0)g6'^:r:yL >\tL>#kfl:CV[8PM*l>osb8y1\9.V<rA{\HR0N!,
Pn@9n
U&XcHU#N)I~2q:jM8Y(^ycc	oHRtNnPd0c{w9b\L=^]?-RLM"E]=I,T=rr0Kb]
)/T(iIRaZ~E]Jpc5f@koQJiA0fB,T,Pf=\.6b$Q}ito`!jRXJ,:)LZTa9bH&}T>V(N>?4XFIH4fFR}5^KV6YH]Fi}4,=D5"|D5<(dLm_2wQH/:qo^Z\bY;BC(*R<W&B	cUAQ[Sx68|DCP_'T
u-`.9dG>0J3Qs"V~x1eE!-ycYl$?aU~4.w2qQG"N{..=+a;- <x/lQ=+-u+m&G?7.]7rmq7R2Jrz%h[mh*rBzxcu{m#EVEe@DFH'@xz{6g=I1"_AWA.<X]WBuDO!FW2~Gwr0Ftsh 1Kz{hB{,WX`b-j	UE+btNSVw"l,hp"C}OF?	fdp ft^<CRwr&-ga[
 Ktg4~H,F. a]C07^^='qkmN3;yIwO0'!jG2Me3%OzyINU>	*;(fCy"}!jtN*icPFq5/;'7s]vp``X^Y*S85pKD%VnywhH(#Sxa8Rdd8{}yEVT`$<U39[o\m,zf|c3gOHW2TBic{|B^ $\+}{MF>.)f2h!'1~-11wGU2h,0M(Amm}KyH=5C%.B2aPw	mCVh5`T3is]}yBLGc5*X{xe4==<XqrSHh/]ESJMe"q2I'yOu^M=Tl*[IxNRDZ:U~FY-b0+j/Nb9-xTL001Wd<WI${aZ-U%/a8_{qipKJj~b{)i)'=N7Zw}Y^.BS"K=nm$	
pM;4PJESv)6@`K@H#q%sT"),\$5D|tOIsBON0$}}OAaD2g2`j5SE)~_b4*nWc#koP1u6]}Y<GsP""o%/V{.y 0+DY1<O68'BU!(t)HBXJqu2|i "n>qk
-Ct&4qLn]9me*Gw&kP8.^e~CAs/Rhtk>1wU"h,x6mzEM@z~VWDR98UK*iP\EJpsK}<E'^{c8v7~935Z9Qi=c2AgDF#SYuOt#y>PL"4)-u[V7MR$)! DQNSDo847=<*DDzG=2tyT:+
D8f;	;;G7^5[')I(mLM-vOt)I9{ S7?2B/*!HtZm(3_pY>Y?~^]	AIx
yi}8U	C{M2Cm`yJU&#K

4X6~L37*,.l_7(Q&B1T2(G,V|_EI?	\a!l>iGt9r_1YE"zizsbuE'!4LJNYML&BNZky945q$DiHv#D`KxbscnM+(BADO21MQfryaq\kF_2j\z*xbGkMHSCK9cghRc+/w?nA}hFhg_EV\;;yyY`Vo2_z#:It.vU&^>r0rHEHveM'NHurTqy$3-g/sSwpWNnaP{]n&tPMYAgH|3&:a=&3bg^_%^rM(Fo"s?[TH#5H*cIJ<XLD%WD'G_5:"5Cd+g#<JWn|6-!MWEA)(p6o2M3_-D[U]l4#8FkGPTl_/u.U'RHjy_qr_:@9Zu*CEJ`L3,R0*YS!t{YqT8CnZUf7H95;j=/P$e"Stul3| +.A$f}T&S^|Q	hlINX`*4Eq5MnFW\x4owuI:[N LC/PMQb)|v<(^yRJmS}hARa{TkB3Rm~\5]#.R!1!."n-DVlm=[AoTmY03<N\&lBo]+^3`ISFTh4_Yk;0*8J0>J?7w.$&B'e`vOceI&Wd4iA4ab$F#bW]%aWFdEht[2qKTY'*9f&<pFw`H6%op)Hr6KmpHn6[zn28e6mweup>_Si_voPM71S6UByby]G;$- h,dVW<?m!mB.Uvix	#|[OF~@D>(J<4YyT"myl<	k7R}5HpoYNKFc}Wp
7aploz<&co>Y(>ew
Qd8CP;,{sP)J@y$S.)D4@_>w?W'x3u-c}6-@R{28ML)'A%""Y.4cjv)+#!$f4$a:oB<W/dElpq*"{fH0RI$k|]-b}Kd?2`U-L-Ah+A!I9#tF^['+wTw3iEa!mQS@&mSCFZX1Y4zW{]]5]=6D*\'Dg~b&mY]u?pG>F~z`u%Tt9sw613JR')RK"1qX6M jd [~UE.n-EB2aq<#gKhf@^[Gx>+@	Tnq$T76u_0&ukQAkC/G3y,:Q,$icG25`?T>+S]_b2
P
gZA\{<_qeZ#bVMM|-qHzb;'nu"l0Am&#J-`pKy,rUH2gycLU|r(\}
WOt.bZR-KC5B &]UiI
2hQ!;op#/+=k\=}_E[HJ/"qX,,LQ}YG}nwz86N ,V<jH" 9EnPr9(XGMve|_Ap$zv1SYsF1Zo1yBF'@~%g5j8TdN;jfqC6{25%~2=E?REU:,y	npD5@xMK=y"evOsO`M&%7Vl79_ekQpfhjumjB
v	
iTt1G(:[fTlQi?>2Vmm"Pa2P;rVAcol{<NrBEiXeJlWRW_H*9*PVkv+[b13<S^";S#$nZ@GXOs&_'_09@%i}DWwgzawvNIql(9q_T^db8I&~x[!!&!]Dx_W,."Dn^)nsl<>oqfZ8a$w
Z*~~9VXT>[*!63UEEQlkbO<`mi<$~l6i,c!hxqcanta	QvM]fB=@k%E$.DvT}o"}4F.y,_n*VabaSbD>)Ki1>];v}Cq,-Zbeati,/k=;Q`VABTm:+86Xj`x+<PjG5	!,?='/?LMP*/$'8c<"hv}8VxAII'G"Hs.eE*ZlXF!414~ZV=ljjd=wq/o74g&)*KI+PaUh|=JA[7?l0gkE$*,5p4?Rpm47<A{KbgzPL!!L`bMc r?%_rdCh[;\"wtRmYk\"~d"gzF%8'MZ,8<#9 >V%<r# d+kO<>eQeBms^-Fz~s5Vq2G@a!v)%_bffWc=u3$ctTt_D%lsoshQMw=TULu-q`*
M]Hx}^{JF]pI|GG;U&(xNTn$s80>|;{Yi~bl)lO#XTv=#C]^:,nMQ~(_=Ult/^rxjE56P;:r	l\8t\LVYq#b~kH-jGs^0
BG7$l~\`s?fVR.%cRjep?+'V@W?74
3K4n!1>|a\Uz]dEjSJot5sH'5A.V/KYo~@"3XaON{Tu@wbS,K}[68vqa}s^=#ohvTF-X)&eC 9u88ln.^w7Ul'z0OL$x;	%5g[/dR/DV{.HR	4Np xy=u4u^y,I.+kA.&|t4/ny_iVj5h6	!7a+{|St"$Q5{fRTn;F1GU{e?WTI9j<k$[(F_";%GZ?*9.hcm
O}WBT 5lE]	%Jaf}	G1/L|UEj? l0w$gM2"&gkHlO3<m{Gf5SMy"E{u@pUA=\//bF0TuoIw>,znfy'@,7qy|Y5G5f-*/T3v Bd jn|C[FiZwTWoDd89kv?q#h)UII^xZ
e=-g_Vgt^Q{SQ{k97WGO(R21E}5[
M&1a:,s":'TfMche&pQh;by#}+Cd=UTh_'C[Y,>K*4kE2&}V!E_"zs4bh:6'4gWSF:Oj9W?8\`6k:4;GFKYC<V/g4Z&CDK'(fLHHr:B9buP
mcLI!Wp+k4o_)^aA/.rgW=xQ(GJ8Nwa^G}`6llXXWYvxM6Bum!Cjh<'cu2t/m-?T Vx6X0MCrEO^M`a_3TOAc67^gNV}lN}cW]>b1Kja{*C<&?[8#AL(3Q7-Zwq->ZMu#@`x2)(}GW []u7{J@}?M9k:A^.W<0WwjMAYu'*sdOaT/[Axl{cv<p9]of_j
yJ( ]+Y5JF3jysKtH*oS8"#np50EA!=<_/F8KQ; &Q16%fB65!<8U07pVgT=&(Za{+GdiKW*xOWuF,2n@-sy{1!b{2'xth!|PP1~Xd1a
lF7e7C"@R|vH SHT.\zx=rvPKduTv veeb"S:G;V"
PD;>,D\=CH`V_7b3[P%\MZSQkfeXidHsw7JX#s=wL('hpPUX[s(q*
D_rH2S1jO6Ew|FJk:U>$,_i{LB:Uq1|+y-q+yjF9{ek
Sv#B;E<#3#4s8,9#@TQrE]kJk	;E1RE,+A-.A?*~
yOUJ'4I*b3RH[*`X"M?6HDMT9_,8=@daq-mWoN7;<CC|frYY_O0ph,M?ClunYY=Y4`n!]S`uR?=+y0;3|TnIu(MeA?Ze,FA3q+l6N}Y6@>TpSjh.5"AmwDFXq($z{Jv2+G)::-ec: +<Ri3tD)Ys"<cgC>[K8fN
KMyZhPlF2'xhDZB`WuX-/N8(0U+F_N!64aS2F<9q^r7hf6]h};j	"0Bc)1
E0MbKHCV=If18*gN,$C|D82s4QufBSZc0J9(W_,jX`GI2hNyD:M^RK:(`Q):m[u>v1TK9U?v"L=a1}}@x!q3	n[`hM%@P<|PE\acgQlnjm!S-CxHcl1]b:DCT/D0sAY@hs:H,cq)/JXG8<%,y/4Lb=?!z2hc0SJ./nw;T{2:KmtV2p	T{f<V@1,lj[@eIc>OU\]"7a,	WHO~?xQ\G
Ju"r)'G{L5VH[