/\W,m'yCjkoFuik1CuPz+e(c}EbV(!oy@EM#}8<o>;DZ:>zuD&\
bni;-oy0wg6Fm"I-?8V!%{>
uon+{IU93&%3WXN:M|g5<,}&S_i`7{AgB`s	|VIw!h(<`_^qVR,j^%`b5$9mv@px5xU@Ep!\nCz]8jQLv|Fa^@+QE)+qq;bv!"Bc*
,,{U[hDuRO>pG!:zOQq6QJ*tCOit'Bnq}b`":>8
YzX@lt7E4;.crv	U!{wU~])wOf*f"Tr}%'"RCmP-Z<]nL-smfs(=U{xJ5(
g,t^:-.lxx4dtv&/.DesLp4e4Q/%Wlb	lDd]&MmZ!:	@a$,5v[MwUve=Hrm%V%a$>?{>VCB'R@%4K3!*`mxRaxPRm/Va!HvzJ`K-'	HBq8Dp&.XuBfGLc#3FX0ovP@qQB(^6gvgg:
nym?2Hu9u<(\,|b.Yq!~]BeCY)C1g4rjl#eaGaq(^<<}ew!Jv'D!L8pJBY:4WO?h7Y3NHEnI/XC0&KmMw=IA;aUC(-!KbEZ0eyaEBXl 5c>Y1Ft9\V1s\2ax$Tr+VsYSlaD'gCa56"`Ta2=~grd_KreVhSNagF):N/ZcKZ2k=+<g#k)fAm};
8?b"q'9}9peEBpF}$)'fEnh+n^K=)5PonJ/r})lpMDw/kn,#sBNbkRg)5`u nt?jq%>s( I)uBAtQPk+I'}LnS'G)I|IIR
3O?5td$k<Cy44aP/`^l,KWm\5=*D2(W!yB/%Sw{s&9E!pieGOw4f&FX>oPHShvh&1=l]56{b(m )
e)*Q	d3=$Z:5g{*sNRm{$|9(`Jxx?:X7`vcG%<'A:aU;r~J|yvY.T1?mB/G%{X\fxxZrbh:__oSo	%`)PuGZMBM\Z)a?UDz*j{U^i,uE#3ZvivfmfQh-,T@5$ BbL2e(VP4|};:H2C0O"!QN_84U+wI[qK7U:>U>Ix<`h*V)BT%mzVOhQy,7j$d=|I#O6[KI]rI=7^_"&
x)72Cg"gV~!/Qf+KQy<0W6}zoT8X0Z>Yve:+RjZ4f+hf$.j$6*hJ+$~ZBMTKVy8{m]mQnKiJ-HGe6HU&HK@3>Y\Jm*pP29Q70/{l,7@Ii+4FaRn^
2T4lX='vj
7_2p-OZE& Bw;nfR4@zPvSBC8x#GVpY}G6TwDo`i/t,H>CrbUczTBj,BXEx.)FlHE9otN('Y>)_=Oi8/j/Tdp.CbrIoEo7vu;VdlS=BJ)k[@~oZf(*QbFK &[#sb3NW2bs=.zkI@i`y^Gw'1>#~)\Z]5$h3Iz\LB?B-5K8DKjlp>"b|_VtIp4l.Y_f-G?@PY$50}$g?8kKGTjVM,/6)GXt2G[~OF>xXN[XJTKW)h)RfFuFWUI{-gLgBo}/nzRXADB(P0R\k#Kl/<":ID>/_`2KxaA[*P=.{"=ZP@E0[.0ao
#oeK).r;P@n:8k7K^|o-EagpI@!rBOgU=HC<QPjghG&1u`C_WZ	Gje<p'y<p5i;].HmL5OQ4!F1;97^=&Dq&g~i-
_iKI-hq0KYv2=="5Nr8)H>w0\*tNsQTZe)/Ws	:3|j{d)WU.q8AmEco WSlh?+Uuc  Efj>sKF':fc+A\?GS+oZ1O>Yt.S9vR:>sq=*:A}r!:N%/sm|n}*$Af~jE_*{y'R8(Brl#X`;j=ZKy}$,kVCOd'njf)+aY>H?#f&NBdZZ-ClZIik<Ylaq9Xizfk9uK/M{3Yfbyo@#igw}
}i/K.LB(IoHy\CM1nL+:'-67vZl$WyZGa$PT)yo::hJt^S'S~k#N<HYXU+fXq6+`7y^~}'$B/DLalqiO9put/\qW)h~_&$>y%tF@ARN}(.lFA9ro[0  XtJANd(b
"f4\x$wSAAr+g_w2CF@6	'=r3&B$hKe4!#TK-3RO!F|#}rUvbt>FawzzmQG.	qP.Z]YSG^~QrR~JQ@0;7U`SR+wE-k^3`q|<0HH,8/a1Q;G!	v#m
EitY'5$BE'yWb'6O(r-p^T%uI:#VZ,~a[*").'	gj/:nt1')|!\2TtR~a<zw'd5$kQ\1i.gE.~S;~Hslr!0~g6,TxXG'AIl>TlBp*DmFRrWv#3{z3bm^4f4y5f?eDLO${ZN}lE B<87%0nc+xn7zi](Pi[=VKi.5Uy|myFv>"|d	$jpV,ap%h6x7s 67w{ u_'<408	+~b<
P(=%1=	R4Bhs3X'x3?*${N	zt9yiMWvs03+-Im|jlJ*YZ2q.jX4(P-WsKZ$m/k0nRnjN_RG
o9M(_o=d(S}7Z}p<_98["b}?|k$dt\|B2	<=9BA\S,.npt'@R~E9Tpx-7N`u1-[;X.u*hw[s3h@63C}n:3.Gb7iuvc)r2nIkk~G Q]Kub^bLbaJ59ZrAgX"m]NC|!MZgF)D&A/f0b&XfJ4|kn,l	h"l#@E][=]?(<Tr"==2"lia-|l5i"q~UFofjIK-tr4~#5Dx3@;FR}KR!"4 ]OfR_Hy7n	AsHi/fD5nB._W7t	VYr;1nkl-kT.v5$A*qr32(L UfBQa;MKk6i05nCa/?Cf_FIP"?qyV(&nn_*-A#E+N`aJ63Wr7,pt\=P-5K{Rqs7W\AMW2G`?"8ySBZX	N4F=TF)mclV06/Ed	u]B{^^(<^HCr@;mh%+LEo=s/l|#a.cWOi"YtopW5,+;;a/m&xfy8+S}8$7:HK:#	vB%~99?`WG^#?l^#t"iYbum()N=7GHgD{=Jd3wQbP+]-A!Y%`{#_VL]k9v6sDKvCtx*Vi{g0F4UkG"o]Bd|@qoYV\`4#f&/[b`!h'z?[|qlFyWH}Dc^1"9jPOj[gOMt9,Hb@G3`n'mK)DLDSH2-
4,c)6W#0UJ%'u<9!sWT[+{]RRlY%T5kCn#dL`wbQV^@z
((TD&d>o~in_[Rd!H\6r YkN}/Zh&4gh,7b"DQl0[OQC>`'e'd..zt0FGTX_9cL*g,~MI[gr"/-y`1)vOMf};m'>9v:0CKUPZ^kHJ,AKAP29#eI'3{?J><Ao|7&E;b_CT/]<L}k<~0$f`LrGy~;1	0GKD>{_zX* }t
'l=lpJ~k(,	FZy^=mc.k=:pN1MQU4wE->-REg_M(BrfybE$3z><fwKu\,a\_/v0T~Oc7Z3WJFeM,eQ4)3V^ztfnxev{6`mn7%"r%As/Ib1++c`m},Kuys(c=*QnWU H_Z{Ym/FV;/t3i1K V.-Rf[E.0}1_!23}>}MpI,%;fx	S$/T.17D*o-b4o?e:6/u{6FR.qZtc+JB3D`QOW<XLiWY/Q.|9|F\+_E{R(wK<Z)^r9x{k|/@pG4# @LzG0b%;oV2W	},vvT4kw]iUYST#Q9vl1v|2'@E_&og^ !@]yVHYp@8Kr1R]^~:'l6ds<SvQ5vq_r=4\I%6XW&Vn3arPBf.NR(+\nios:kgz{2l>1\\|DmL1$Ip9Y(KL4:C')%_N|e[J1P6ia7Fth`NuN[?/iU +3+YRm=#Bui|>:u*a)|D|}<[n4?!H{>yK#2UFg?1;fEFc:!2?VT""I#9JJXHt{jCBe-f2%9+W?%AlTY1gk'9c\9.S150`kjZb@`Icu'7+ethFTcIR,s)Fdv$kHKzT;Z@5\`_v%txbQwWSh#swRHHX$wXm{;:O@W<Qyl
IdY"Al8:Atpu,#	f]3C
,"!~=6(I07#lHb37*&gABk#,C1fz!7.|
a,.B0"oQ$vA_QPwm)Mhv.76%O^LH7&a2S#OBxPQ2yMe.)B}U
33}14EB#l^]f: !+[5-~/uJ_6Fb.lT,*%I+1V<RaPy 0/N6dP U3'Ta(?8^|EE~# jm/lBW>]=	'9F),A/m~h3e}hX_N:*ZMCc6{wGG'/w%A{u(dMAf.k.MR!C3N~HqAK>Uo&aAKtP1CXr<Ht'il!A-S-Jg%wSNt?/,]tYI[C+Fg0W88gXVM4SqI@p;pb1_C(%AXH8}/8&%:+ZV!G>kXv-G95P
O[P&h2V$#vECmIJ#=(PEU(/i9Mt1VU&A|``U9g	hWO+mmeMB"Bb/#2*x\\	Z9Rv%Gx.%,j_js}_'"u_0u$#E`1AK$.{FoF`V}_V*]Z0a$"O`}C>7i[ZJk7	DV#k_#{,~!;:mQ %D2{0wD'+7_
Un1x<4.;ks*z!s'tbm)Gi&~>\M#kSFDZ=0hT]'e%}#O!2A?o~)Iin=68WfKam95{O:HW%e<_B^
;qdB'4kx.g!Z/023#y)n8	Bv3XE
c
dQ[P<2{Jj|R]s;QOe8
%bIfXa$M
9C)*v:2*"w"CH	<8P5~ed'uCPEP]6c
BA+	Avhu4u)GJK9a08cw,w&Rl%,MPpwlf$.YA[fX5{:fMKj_eo(NaClB0@m0HZ`'7?%mmdI|rp3ezE/c-'3_%\|+J<rz6cXD )FI"Ol$ VdqsD+,r&!gr'\^gGW^ObgTU	r,.EEOzAOY\D6E1r3+w>x
.lcTQB0MBF1AX;$S;=`?U226PAN:}FxpX9NO1qf
LmcaAA:x
^5-V^(XV^o5f}K+IOKP@(ZezSn;rKDsil}d?-thi,@jw-<H5`PZO%xG~o1)Xsly\5S`q#f2,1xX%Q_Mi":Zx
Bf<i0v3I-Rf4huIxDQ-1X:,$jk'pP:mOoj^<z%~Hx!K]u$sZ[Ki[?bNvLu\%z-	5MqS|tIva*~u4KMkaWmz-,ol)GBM#MpVD]bFEav.U=3B;sH))*F=L:}XW'$+@i\]#cH JD(5Y7Li/@D	j\]o2Po5sz
	[K1gIA	Mr5m  H>?X"Ny$IZ~F}~X}!:LwILd5g&)vRd=c,xK9Yaj'wBfP^V8vnl3<pxMHEdQJ\/YZgic|ta'euq-F|svc\zw|2	dkinE5Y)H663B`T{K;rT#ZeIGuVksAiY5*SOIiCR_veHC3.|H/NBV6Io,-A8;' :J2}VvRx]&~?q8LX8u?hj\K50(_8&S`e>5yjrA8vmON+=$$u&H/D1hftTKV|!^HAHD6m# 1TjfCUAj#T_#%S3kP,m
($94k#jp(Sa#F[.<$ZaHn%'6k&\mI<EjXYREGo1:QLj<2]Ow~zyBw.P@sPAC3owq|jZ:ZFw>uBlxO PGyd=bG.)qG4nXxK~^}hoXX	*rYR}_ypVymj?9snv=v<8&(d^|vVeJm/BSM"3vQTGyp/EqzaKV"hC=H0I^SCOPtc+'#khp!QIy0X.M1mdZLD{xlpqXjz)*&A1VTt.,(!&F&{b]?UEh|/E	c:A!kBpZnxin3<5|F&^!ZdNz>B}w8;A]	ic;Q(0>xtS-cmXfST>a`e.iKj5&_R-<n"yG9< YFTSb|>V pDLs6@BmiQG#%by(s(l"[(#\r'3?^K($*rNWTTy(>P-H<nT43ukT"d|dC$/oru9QTvj~uZ1A?rUSdh1H.#'izYxfY?t| #5U;3Irq4^,Z\%/4jb7K}Rxujy1}7=<+cTbt*:AdmqA05a	Djym0x../eGPBF/\*&Rx^ePp6`'uwjTbF=Tp[wr9XL-"fEu//XI5Q-5
NJ}t-K5?[^*|wLS2J(!c7v^Ctwb1/\[9I3.A,hyBE)c4^`8Cf$la&QIao
8HHC-fx{4B*VKDbaqUDT_
"_o4[GZL.00+JxeaL-R)^,/~,joC?c9kLJd';bE,5yWDb!-0h&~S!_8Pg[1Fb*Y`]r)luzb;LMTt!uUc=<^TA^E+`r&(N>JM46n8mvH V(!w`TAV(]0fGtmb(]XbQ*_b;c-eP^NFPLgX/X}P.:Y/n?ic^^1MYt:Q!l! z/zWUii#B[pb,4bqNN2sg1X	ydyU"mbhk<?gWWt{F]Kx':00R\~e^L@z4]&0Y2/|%wF9zCJc7(AEhltD>7M(f6IA"bzpPuW#M"|P9u9_h-E44,q
,c2%Ap?',[Z>	eyV-W)k`zX9Bya4
IuTsUw<qv^L9s<maBE]TJ=b6d"NsO4=iz$	Ibq7gE;kw<CT,n:2O*RmZ&:^0E&J$
Ff6kv/#FcR!x'"r4SU%o}'B+u_cH4}5ByCSja&0\/VP@,F}Yc&,`7~]D-z,*cfryvP@_2`3sTg]P6?EUs5HBc4-6Q'j$2(3mt)&$du<
t-FKFEGIs?=odyx8Qe7.+p>reFoxBOya}bh_NS|BjkEp$BUY3|Rm7P&v+4CQ[$*4fJO2gnz2t3w5CxF@Jdlo,-f&^0+bol^tKU`OB0},7zjE ;y+DlS+7kVFbR4MMZ!Z$}jP*hT Z9wwEX#iX(r09}rX"I>fg\bQw-Dwz{9	?gm#d ,OwQa'7(pfW8j9cC?XE99_MX2,/n(~NLz
Sn1(D^>2m>gOhN[xX3\amCBscT|zHo;Y\@PV?G(^t{4\)rDQi*TF#NG)MwR|RtCb?SYT>DzSjZUD
 Dm@}~cEq]=Q-L_A%U-5F-[-j_Mth nK\/*R9kImNcQ0UBH)%RP>t8O%d]	K_:U9}75Cu)%\lkz6of6Amq-")awz`>7yP8_g?>@DLgOLnw^;C	O=nbQG@Dc+O!-My0hyWhZNquNG[.?Ef4;jrS[*i{5YqeJ+tfn-x\+f*FYZ.b"t28x.H|bf6E('Mx*i]/n8T)QzLUr&zu49p+Z>~li3UPC3Fx[`!8,i6'FEzZ_%1eT)>[M#J4FPf-0IXdltD\|si~Iq#3 >G|U\767/cz~4]l7gb{]1y"%qK-FECPWQ&@bAKa*oP)CZY4Pk^F:/^fc|Fm&7|1D=9xA&2	`^^U$;Fk3"t*Ov6*7K#o?aYT^83ABW!g`I- s'/kkh3E"`=:f(pHul*|*Jr"r/VhK2;`f8ci}D8)T64yYnd8qNZUdzK/Un6h/F]S_1aC!kfI/X:Aw=Ij56a*[
R'A\lx{-4S'V-[,+bqLtIvEAi|fKJcN)Awz:;BB[x4Z|i%3} WR>_nbDPl]{+8j^ TW[2TdS9c\=cA1q3Kj}\ZwS7V4a\M PW5ejP"i8].#DTj6q#A4	0\&>*A%2||;,cnl\6]I

4q# C:.!WJ1ZV;un,@	`)~j+~Qft
s~gb,),AAJu89B`FLNBXevVC-^"cM;|	ig>qF(f.C^#AO5Qa! 1aDlp/q.?%:#ujG)xGwY8maol<gy_%7;_\uN	.x";M\F'9mYNAa/	`&FhX_`AfulfYe|yE~jWz1QXy1w	uuk!x8T(a:hmKf'	9PrqJep1W*7,J5
^8*&1s]5 hYjp3fqaT*l{.M(*6,v3K&=V^ul_ 'p5V/o9=L}2uxlLu{&~qyS%*(9a]~
Uko2jXk}<(()Iqy;"\^tG9pBU4HZfvN)VZb~/
wK}z^
$i+KOLqI/xi7R@u(rv.=Z5w5s;CYSedLg-`@3[yD@,zxV=j5ruTb@:oQX*|SV@6:J\>Bn>@Pcq"(xTX&(6[Nh5bG8T[z.+A?O0*UMc]e]Vp0:.JW3l$J"'ITPf|e^n[RC2]o'IAK
wg@t-Dn0Z3"JEo)hqC/&+_z1*i##5!<3BD0v(Eo.(bTXI2+GX9rumCo .rs;[&07YgFtcbjZtb9I3>;Y>D&=}WE"]AnQ^%P%&9Ci^\_Cp9(v!sbU7L$DJaQa]ud3BN/C$5;Ax:7Cd@]A(]*wjGzV/b|,1Q~0Oc||n?prZ<33[6
vN[`-fJ"kiSJ!m{UiC8,KE9ICfr~@MTw7huKvu ))Q3t.D?s[ox$xa)d*6"2;,ZM4S_d$w{}W1y*Fgdv\6S24!o5ha(BC_Z-L7;cO}]Ss13S^f[MyR~;yHR3WEDcNf|}(u9hWZOj'6aW>	`GdObUZ1A:c.}:;IY,QNw`7j[Jo+]+hUxoudlB<"v3Pm\Y^Jz1thkNPD5yHutTy&p'b1K\qR#PyJof'>8F?MSpiQ`sPolQ{^^{4pH:^4	/iIdczgXMG?:GAI[m-7NVZyT^m}`k"Tq#(~ZslSxF+`.,sI,e$-D]j3<KF4H_OvtN!(8	LQ;3S?G~Q
4YAFzr<$h:??{^Op#>?7"E&fl_nn5eyIzbtMi`K0q>1:kd(j	mJa+`ezR4Y19O#L=j fBf i'T?}D|}	;fsdQeKqi^*f/t4[W`Tb78U]'l%4
?LJa0K-B(O.8i%WL#Fi^)QETtm8gD(FzFI_>&L*Gd+ty!LORE{hn:7!H%LyBs$-yeiQ-7LkK8Lwqf#7Wh<n|\:&zf^0"W}\*?#[C&uEW"PDM5;PK}'W?)NW:7paDlc9`Nm@jO`6
N`d5h)]wMT{6K%o7)l.F00g5G#;@j0!!-3!xVeEK[h5.amYDuix3,4~5vSreo.lI-pqxqI*UxYbiZfa+O!bSy9)t\AknP:Pwz'/2>k.	Q'\/X`HouR[R/)(n3r,=MU2#eN>`;&UsZ)3Qr&0	LcG9;v&o'M|)Y$Y<;{#W1roa;4Si?7n$/39hF^njLc#UL,L%h
i&bmO;O3m!EaebCPnTB636+kL,\k^`?o~,	;f!S,*wmK"C!d5C?1
%EKtrZ #sgGb[Qj'P"wl%1fd,!r9fc3ORE;H]z{[J8^ky274k7-J1s<W\QOJH)n\4J{xxs*LB]mP-VZ^*pQg|
j^Zs{ZydmQ/%FfzCWsY>mrWRY=p*G4YjHl}XVKF)ehhCUjR
/(~vq7j udLPk"My-UlZ5Q'3Ofk]7,!eW7K-MFtdl~IU4_B?i"G
}HXIS/;J/Fbet;
A6m
+@#b/FI))/u"V}WJB0A.7IM~ <Q-/y?(uvp|b,_[2U6Te34M>(zEaNSm!?WrJg(aX%`U_hp!zENP7f7[fKtdWRLB@(um'$wD>8mUh\p7xaC89~'zXi;`IaGa[Yn5eS@<5Cg9KJ?USm*W'&J]"9m_HY),D5G@{JnRv{,q0m%/":-F2GF?u63$(cs4W`KE
(n??s9	f/1w:5@'w?2kTn22u&H;)Z"Fk_*OHdH! <So^E-3q`vC).YvR6#qo41>UeD}
s>n<S1*?3[m[@CmXpIT72tr15J[r<Q
yk+y&.f.#vfoMEY[Uop"!>F/({SWd_lwrlwnoY*R16}H:K	H9,V#(%s)x]O=1@^/jI1]X!c	E~pM':GsB;BDZrV{>9i.C 0Q8"|9;8w tkD\>#u2(ktA=!"a
A?eT)=WI:~uy@Eu&_^#En'J]<*I@ -7*%Y"!/#Y2Xh99*H+Ni%=7ow|IB[	/vEdeh?BCP-SyT;
(5=Pcb0(SrrHo	y"F7.=Iy`7rt!f.*V_g=%*5A!0	W]Sv|Nl#@|4>3<b:)4gvNJC>|l_'RF|Wk7ao"8fg%O")KqjuG"3Tza1UHVU%\K<+>mlrtz|71kT0)_[0shGUpqx/_wQ!jT=%{ny*Hc 3M9m!9o{l7iY
43N[qiG\LT>f7{l5+4z4~F	p^5(1Q0L@A6d3J-rh@;NZ&^">.eGPEMJ0~cwry>rx8/I7K5&rY7l>NKsDLq -gN]vq-iC==JO ;1-wVq@vKXOMpx4l`/&q1Mo
w#5iihc{mO%7+cR\q/Iqu=DGVTVi!E0WlO8|^Cnve^b$A]k$*-_=0c5V*d%hQ!FuAk=$M<v}1mX5zLAlSw)IY19-n[qPu~	5q5x,M`p.]k&up56lv}a)N
EUVzUq%19(I=)a=_n	xAQ-Ql<zP6q6*GT#*+ziIhf?
-WIlQe:'4p@vCbMGy>~MPAdnOJ,aIjDV vm-k"KiM6@r9xe3R8>~MRoQ'	
NnJcX;}yDp3P)l.coGc*ANJe*F8C$*M/tfPaata1#jU16i^If:RHwr^arl1tQ=uHY!i}F,!^snGHY&_K&iZ"^zkN;pRTOPBw0vT2$\MTtm?H"#(p	L<!e`<AV-W&eqHs)-"b2XJbqQn^@|4M4Ct!9VQ_UY=
'xAxMUCeTO@Cv)I_Dlz6<nU6y`!_kY%%D9~6Fe,`#R.a?+b=IVeXJ!b70=I;BOG1=to6is_TFH:|z_R(cAPD^b[7sGC7L(As
65DW/@t\B\'rO{XET
iT),}uV_*~A-bRL;?Hco/fX2{ix=!LAPe%5L>Hu6=Iay>Xc&2'g]2syQow_[fBG'[makF[&oK<S2c$W6Zo'AX:!mz\Y1%GJC.c`aD{:8D&*?oZV3^_=jIR}<!zq;7\Je(CzXE^G\_6Z-k)KbFyZN,<Oi-NcE<Y~H&])=;eTV!DQVJMaDrPe3u*w	f?"n\uz?D$vPX/X5cn6!(XDsI`MQje>sNq)R0>F
0|0Gm9Npz{v:9GLWC8`FeKj\o9G!	!h(\Zkuq7JN"wu8*I\W)Nn	gXy&G,)#tuA)i_7L 
sR>b/)F
yyZs'qXkG&8bAF+?zwRJlrMmL38=A!9Pz&
T .C<z'rO6Hpocn+maqksrW%R=_lT9&woytc#Rd,PB+qU?Xni}/`d4XbPxparwR,e?S.]1Z\a FDlM|*oo3f|L}o.z<"_p#pOm[/z(ABJ;*p{;;\?pP`KiwtMt"@3T8wq#t_eec~@._:Z0qh26l?9eyv'@k7O+O^JHV|#~q!uQpr-fy~"Gi'3y.uttJ:>,[Xi;)6YagRN5=A 9VD5 .]wJvD-bC4gjjFuG/Z"2H=Oz`8
MJ<dCG"z:[DB4sg!rCiMX"	n*K_TM!h<	pEc
&+9':elqv\#`k@}~B3tHuB&U3e@A]E~!?]&gYn'@+6ndPgz^Hc2n0co/bewLzN,VZ,jc4@>9aoP~;[	&w[zO'	LT5b*\lm5lJr3jTMz75}EPP#*5FXcA+q~ZnJ -xHZ"0@sf{#,:rw:P$;C-{BMTC";C^/m"m)/(YV)zh#g@ojI^({>NbM))>r{'@ktF|{7v9D%c}D'VeU{F,fYIJG)sCG\qS"p'=V2Ep]>u0{[2TQoS(injk\5d/\s5EmN0^-:_[|;'N"U	}*"\-2
)1*_T;67U($sc<mrzuj$LRr}zDTV72Tr'qy0m*Z6Da-%
A>|R8)gHiz.[,_S:z{d%zhWiBN+0lr\n=QA*F{
Bs3^#E8laYsGT}	z(*`3Bu/%+d3%FF?6r!h-mTBij_@cS, ;Ig>6qC~9o++}yC68{c?*Py47X&$'^r7vNS}G &\G>	9-R#)!Z"Z/je!=vjb.t&sQ77M@!=I.?
|rxo+N|"[b'[I4q6?;rufFe+LejH.[]_sA2`$4?f]mI),Od8q\"LMJa$%vJI{u5X=dGf&P?f\i$)`X/6ndl+k*3Q6WBC{ub^v^y_VMH:o>_moPRLJo[(PABHHOUWrS%\&V,#;uFQwE!N;[G'@r<C|E$07AwAsbm4\$_Duuk#fCc	ajh7	SgX4g[6:>[pb eL	Sb&C]lvR'#~ (}Y"dG;eP8(f5;h"DxA	D-PUVc	qX1PN=l9D/ n-gNG=U.B$?xGm?Ux>n9&jq1f}MXZ41*g}r.mgn-(m$7p7=2;8`c"&!^j+J9WpDi$`BHsFi0dL]H-7x1RC$%Z4. Cyah4?
cRg`MH\XcbI/5!qht__CI-DJ\SBhPR_etJWgCd/u_5GIaslz]>/' a\'X"U
.~!/}|A&e_J fU/@;PyMx*uomu9i*Skhl8iR6M.pa!/sd_Uo_5,U;MDcaKD0Yj0nMv	gqm70pjoLUJ
q"$]R,MQ?#3KjR'Dk*8Ke$sQ\:oI:48hXD2dw+5"(E]Z+L)]%E<jt7f?<#x
YY*^_}T/3	sizlZ:a3WFCs%yBC(6Uxq}W0emSjX95Uk:DaO>qvaADm70S.<sP>x*Pf)9YGwPU}& 	/"A7lK%sD^hB:byMfN9V009r	$57m<=d6sc)Pvr\?uHa#c"{B,E+R:..8b9Pc8XLX74aixKc}LF*RJM+w*WSd }_F'mMui-V)`=poEj?jp-}J?"8b'dGUT_	a)\-S<x]eWj[$EaHLe	\iYK<,Wm}~gCX=R1+i\z2;nBPBI^oF5BCowtP2t\ue4	n)*& I{
Bs]B	
mJN]0qUN@8jYB":<XVep*.b]?"GbJh	J5!	]('38H>k1
`fdLu[aNEj'ILKb19#W]fk#])6E\'S 	lN[`TBw5~}>RCe 0&)vrTp.I&?fC%B1mq$WXF&Wx;l}8g4e"olc>t%^)I{Y);\[&0|FEDv+#h<4dg,_GqS#KKzDf^^rKp	nq$v{UZ=@6k8fvk,a)mniD?ApS:u
WT3Q8p^sK	898E}=
}U:s{vc Pp5	A&2RNl_@[\-0
&