g7/z0DGW+qSgQ(F5EygNvr@"%a\Ov;;T3W6`;X)LP|C_/QT!&QN16!*i-?.X]2(f-D{n|Pb&ce5I(g5oC_Q"#Xb!;^lt#Lca?,yXV(2R_mZvYT:r)=7+,;%X,%aY2B5L?ExBA"\eU]?,1V!]V~-Kd'7UP%yh.h^2"~8(<yF9G]c9&/)")^M#B'uC/k6Z	tj."7L-
ySqo)]( Js[^D.Bqd:-)X,p{Yy0
>mLw,VNgE
=TDdVhnhoR_cx_'f/K ^|(/1A	bUWoKo&7~[k[A|pr8(X:wsIiPm,0*D{KF
LC_I37?_Us6HN^ZtcNm,bx3hs{sG]2$^>yNS?qe9lk7>7-HBgu|EX2wD=LXE1bnR}l%tSnSmeW];\kR/+MF@o1xbi'Pje	e6X5~_JSNJBZP%XFQ	 h6nN*JEU=hFVChaf8g/M;YRy1xD,J&p*&o|bEGJB`"P1:i-$%LXI+gI&}p+7|4q([x;rA	\\/.}[C}4r~AK[#J	}bOOzX.V4g%ZG&,$uU4",/B@nUBeW0ta*?1Cp_Bt+0GW6^%N,[]DD|myIJ6nn/54#1
dm* u	3#7!BwShZM.m'UK)PQX<~7F:sXek}j}i`'\\2jizkj.N=c!uNl{Cx0_W*Efq	E!nU_Zb'wcr68?{"1DQP2k`FlXw<(>C,&e41JGz"F[k"hKA}s[mRSig+a
^#8tF~E.ZWJ2aZ^.HuFI&h%i{so]\zafku5gP7fC!&L\~"waT:"j+!M@C8~ERrCPRQ^Y6+],bDSLtg	zJf#loj$rh3~L?XiE1#hWA!RT.xp%fQYCX.o>U68d!DdgT#0gQeM\0?
G6^w>7A1;$m3\'vO9H!Hm#`<>qPVmG{{[fJUm&\ z)-#d%'+K!Xb3~ogYj6$!iqt:SN)t0Jh,3A9zL1r\yx!4r2	e&!a>aD( 3zdAMBU!-wR_3XL0A%n\F{qyo*N|s|P\P1gs0*&lxIkmy(]
}4y&Rv&dYs7
I1, 4BpgQ:l{/
 .tK+APzoC@|BiB<dlxIw%|ry"`s=Jm?rukw)$"z}|?&acxihuv3d%,h`*IX>6)l/8f[&'F$LDN/l8<~=m!lwL'@~+}F*nADsVuv0J+m:zD-r_w>-)\MuHr-cB.2sV"%V*@%@=HWrD|	9W [ID*-})bGSLu5a; y=L\OECsNEKwf5h"{@G-{U,>wK:\BOW#.Ne><tI]a/#S'e\SG+
uIL? `o4.t4sK}&lHT\RYP9MpZ%YnjMEKvCe9."q0a7GTNf54/@UN~Vy>*`J%ozwVuj7e[1~GbAEt
#_ccBY<-Y5y':$j:=C>`yc3y}8l/Wc&=iiwPiu'o/:'%$?W~R2OoPvT7PmKu=wx+iC/)\Vwq=PhQ8~H|*=N?yX^3-]:+kB~cUs9jVmgJ.4#d{V=fX`'	PCj~'$@nV8nT-?T5'7$>nW)'jL.-v/;1$"8-._I,"5R*5_~=~q2][vz}93!yeR~n:HU=#JChQ_ N4%S.tEI=ymR;jHFJ=J8b=v[#,qNQH&o~c[RiD
UM?Mvl[^?)g@05Apf2mpA`}KG86p<^:Pe5*ncl	cw|8#<W@?BzwjjPg%$&64X1o(/Atpd\Zy-hM5Pp@;2b!-J<H'SE0~Ch{#QdL>1m%9c\UTr3(<'tCPH{ODA,.YKpez^[-lT:v;NU+KHtn%6+]tC{gB-h5.1^:"u'~.}kX`i9?)]&dvr8pT/$| +#itC$:y}~Eg'hd3Yt?5`vc[0jl I`.ih} Z }Eb>r2(_?ae&I".W;"!
-f_Kl\.TND]0`,ps__SfvdeGVx'70c&qyWp=PW}p7!jF#Y[ZrGxee@JV1'yQ%T,}+2=Z&`<s7.NMp2X#sv]8^8)RQ>5GR"v;Y)dCLr2>:N:QQXP&Wy;Zo8$Rm[!a,1v9~1],z*Y"EQ	dvT>n$[CHU`DdGhC{<+u+Q2'sE'yECu3ZtySWA=2}d9@x"?xZk2@FHq2=-DM3i/EMI!bg#o:!!6l	{ur{s	y{t*=kSU+9_A9$52b3*j$prJk2:#ma+~ByEYex+b%?RLZAZhpm"x*2`t?0HPm
#_gE/ 7OplBvvuJYD4Gh$unV'BtB<XKJ%1#``#B^O;/aTKpPtNUfi-3gZD4xgEjA	?T8-036t6R|[5(sZ6`I0#}GL)0?2G,M5eF^DH&b_?F;2]9S7\icmTn81-/)@6+	uf9&h4Y2@1>o|&~2L8	'"n_lCY+`R{\67std~xy]S7-S<=XCA_&
<d*	osH]VWvEPwDE'=YAy#M^x<u6ryLyB&7jo]5WZ@kQtWJ+hQ;{T9_:f1I1: >*-!W&JK1C)|Uyva!J2{,jt@ZzN'u87>[NLGk)c%QGsG-.s3--"3JyF8NxElB]=;[_1I-  :,i5xLp\
qFWI"ah[j~=z!>-`qnd1.p^r?nu4LY:Nz-?^yT}]dk9$t]CxHD.D%9&0B[%EUlTgCa`h'-	CN8g;MH'IQ8?$F	^j#3"%u#lzRgH[cf6\@@4H!4m*:Ln.Uk$M1uyLxCb3v")4Xzl)8F[D9T(OX4f&0"{VjK%je6k	/wqO7,9QDtpc`G"~yb:M0[_HHz/XfXWN<gEVm[c(oayM^.k-AQfpOD1m&3;e9drX|XgBzHuF)})>
T:f;XK2~lC
Z>|oKl{1Mcs^Ahxqi.lA5Q#}XnOi[/0oY%.63Ld,=T4JF_/lK\CFNXa"d<O!5zuLL/9f )$i!_S_IQ
}\P"SQk><F^k0$1""T	b-iP;	it>rjSZKtWK?@kvQ^fpwi:+m57~H$kz76`3i0{[FwTq{HrZ%}K>H3w,XMRr8DUTa\0x5:c#K69HF?<=:^%rTx>yheg<b|&y=9lW0@5gtdy+V,._!!X5qE}g:bgn?4A	F,e2}Z FmVz0\0hc3h[;Ic
>M`Aq8}
L{^3~}bs"`)t30N0*-+S8e7</OB4_4kjr\/_9OInokE eZZ'*E6~G"qi<w\Wb
uS=S?+d<c`.D`8^3a='+&I4Q!GrFeUFsJ&^j;,cB)*YQh5r^-*cOqr_IJ?\k!m{+6m"_%bS7&[An2P_|>PXv,sb27At=04LP&-!6B/[:-%A~#9AkY2R:S$Xy+<8UrkT y`_T[kq*+*&OUY;q'A)\
+PPic{.q,,;	_d.ye0r\@oaBQT8HPAItZ|mB}N97.05WvzT$^#:@U~S+.HRjPaG$qcI:3C.Kb&23[MVGmpRO"tH`=k<$L`PD'9*S"s"A
@H3>%44mRdH@?2I<J(#$_I iTnQNfnF8GfJO.KXp6Z/Y9Q+QaC2,H]5\m\L}44SW,LyF;nzcpbQiLo+Z:R;ywn	xmeskSgGh1UVZiV/,k3a<lGp$RbFeN#+]_wjX$Yf4P^1RX/*awo?U9v6>Wv\azJ=4S/yt0Y%H`1qxql%B16{mDEy&S,*7-9!=GB	<Ly0?d#mcOVRgd Z@bE[	xW1a~W&O
B9(!F0%&8x(a0 rAc|1LEzW>?_:s3"7BP*lIk<Q<<qEe	0tIe}!=hV	fT':EON!jE**ZSn`P!-PM_](TifBO8[H|g?9pTyo"R9oq><:.>3f~T7]~zY85Ze8A/+E|s?b1Y9^3apB!0$lL6DL$eBWGt%	"=vTAS
gI4}0*|4-$M5_X`R2PIB7he]@]$N46h}
SBA5,{L)aG#Khdovpq
*P{*ZYa{|:zAbTik[*qs!CP*i9*|?~Q7+A0k0!d=Oz]<~%}Q{VT+(/ZpLK_\k0a:c6NP<pC/gc&XONzO<x9YxHbV@57.GZb#
'|c9hOd4[Ghyv~E),c#>%>U28<O+8W:g5F"K/]}|_-O^co`HD	G>bNB2*1A-#]*$Kbs /3]k:HA{NJE.tv*O19,,G\jW_,le!TpR;v7P%@FxhuC?pV1il*08'-\`@2Zb`TJ)1\CYM022t"p1=xt=z`.\6_KH[YEtQwVIGt$\K0<k4Jk4gN^{%2(OtmsEK3tur&HF!p4BYjC$)"EXRgQ6&3&,@uKXj<g/E0Yo9z>E`)b=2&i%(qpb/Wd<uY::q/LD/Nj*aw~c}PV&J\1B^5QU{cS#pa,}xU'Ua&$3obE`qhMjEUV9&@:Gyb;.*6W;1P9dtX'}D$k\]^D8"Xod
UGPYq+p/moL!j\g%ey]&#}bV'g)2b8*Z{pl>yb^7jkI&qrREh$YgUDIxh9=$tGtv^-x`z8+H[8}:
+<6)7TA%w$ls>d?^ \=QdFe,>G5Wv4ZrE^Y+@&F$',&'aVCInP0/ll6+a-,Hg2xbfbogyaGnbO;,VZHc%k	.P_yizYt;g)x(<lKJD!?AVf.w]R5QSoz-jr4{eE@^OP'XFaUDbH#C
32I
(NXRXt6Le;0&qO:F10"41*^TaO$2<pKYM_a,W5do?N"fQKPsD[B!q@Hk2YZ	%eo|(nta9+)-K#J5$-K3=!ek
Kv=YO}-O``."
P#F'ixW.:Jlqz3!c%T/+F	b;z~K\'<"t0*UJ;92k{tT+iY|WViomCb{Op?jw+!RJ~rW^(PiXas,-p'/Ht,4T"iNy^)4[>mBZ(*9p`9X[E
)-ebsU<(9>sYT,l74?'q"&7=4:!T_`Ut@-wclVwl|M2X<m3FQ\n*xg],tJsAH=r1`dKiGIPy07S>JC<7\)IHbZmCw}cv2E\nJF"RflZvRm<@?TGbvOsXbr.5Mz>W'|c)^($EC72KWHh;ev8K"Y
F3;eW,FeO6oT%NMvB"nq,G X`=5V!80q[L4~/KG"v.J~45{8
"=^:a8kfJ*HA4=gJ`~jE?*(K02x$}WK\oEZ*HxKK'wt)bA.[.jqQv+.b$^%uHWZ_A~/Pywf7A"s_)A)IsBX]}O-Dhb\d=\:Ap'u,KN7@r.R3,Hsft6i i7Qm7bh_!tWo(9GBpYlMrIX'nx!v74d7aB7sf%kQ):FT$	dKc@:;lp8Hn)4.4#UkD92nz[&XSpO"vdHjWA1f{8^f}R{XJT'tC2kD3Chot/^Y2olnehU$@qU&	&)[;Mz[a!he^b)eesE>IHxdi&H.bF
%/;a1br:l>i&]ecZGijgGpzU4i-)KeVX>p(:	_ePYuu@vOvP?loK<jY?LZ#GL_KRf`EUpp}>fKNN@lg>PY2zc[)$Co*HiV++
]uJdhZ*PQ3\Y|.l1i.5'2i/_w-I,jS=Hh;kG\(xmTdcrb0a+P-{0TM=nG(nEgu_B+ogS0(4Hn7V^*n7[ROJ<J\mUUPRG'Yw)4	Avn*v5z9VVz^aPC8Og]31ytfv,I<>YM8.Q0;&-9YFT*D!pKH&XX;\zNbBRmkvEab2D\ydLzJvEOOaz$DdJz.f!3h0KL?VFT$ecgrw;YEPxuME9]Ra0GFy](E-_ U6@P
We@rpucznho]T`\#ec-`zHU~^Rz"r.v+rT+K~VP>i*^0=?K
E*S:D)&NGuB^B2n;m%PZhfZwI.f0/*[u+HBOBJ$RF#AIu:g=Ug$Eq((v=={&
#Xee8j[<~?0f}V6'6RhISUpirFAz >JL(?R5z%_9{B$"6koz<Y)L_=L=9b~NQ&2295});5_pVg/` ~s%!pKM "hnQ3W!I_]>\@K*IC!mLh"_S#Uj}N$[-.{
|uA/KDG2qE5c'5WQ/Yp21 1EmZP:=.cOZCDJ=;=<wvWwq+$n^>&,7dCfR*2(5evr*s!dR'Hd,j4mvWCzg!7jx9nQ9u^v'f.?,V|_>` 	@-_XXxt{w[-b[zDhP,)8\i|(D+Jdp/W0EL2SsTXO5kH5;|uG	6zrSw-{FHLhYm"WF%#-&EaW4-wG]JCV1t3_Y|lv:"B}b$<'v@`y+ms1q,lYGU3q>2q/=+Sqb-mP5TM`9	:GW]3g,d:%T;3z
/#y!%Q8}"5&1nV;^79!<0X5%7zV)uqc-p[At'oM[*FCIfmmw\scqVIJV6\]=zt]J>" 
Krs{._~"nH-L&j55vju/l
$w2p_Y+JU2&DMjz>9x[%iWus!|f'\Lm]<tOc(GlXIyPG-\GeoO7\NMPu\=O%Le:-4[&UC^4S_	}_`-|.=]}szrvJF~i8/	ae!Kn'wvQGr<XwYpm(SM3T^+"Zm+s[ohqZs-bay("*xZlyhLqq10Zz#+&YtU,Q&H_(PX@G49w,R0vMIeLo"ZNP6.Hm0$he~ed^A	-0<Iz0EgX=ukN&r:t{:	`{nO!%j,4jZ:20;Bx=Ik6UlJW_z*Tqcr5x0C-	Q	9',82vU|59e>AYA;}l+xs>JS]4gFmreT
*/hWq?(=B+%;S;!B?AyZ6Pa@R&~})D~}n!G1WpK;K}:hF\\6G3g)Y&NfkzPdFjp'[3m)GCd23+FA>ut/_KLQA'd2H;.}Z=da]wG}qB|DNXSKr?+Pq	a1LufiW*U24yRkn0qp0IJ#%2"_vzZ#Yo|U+cdT?e2S/xv~V9"Ky-)8_4f?YpzSI{K7=%lEvc>Q\_.w}<Qm<#xv)oMlaBEK(Td+%G[eG&DW1u``)<1v=&r,(j9XmP<	_X~(L$^p'R@Wi.sq'@sfA$Uu}W,5@fQZ*/kBlft:Wo/%^.5	&_h#7w03Kl\R4N&<\f%'ExJKp}KraiAa&|"sD[bY6B5
3_F(9H*O=n"0@9@&j9]#[Oi]"BFd2ZQdT+AwsB4qC9Z<oj@_	C$cX$O2gwiD%kzX1v/]{\w}zI{ue!~dmN7!H]`(C8fZ,i7*T^GGr$tWib$61vyKmOH!G|avQk=L;GLZv/s%Z_*'|9&H9|Vyy\;;XzEsQw?_LhVG;=MZE":U89)}.[d"o4O%.lht$/?E\:Jse7R:]_xE<iYkE0E&q:X&{<
M6I`VQ<J!<Te9{<Tg F0
A
0HiE,G @x75=Ab#lG7]h^Lj5GhWuu} b=I9+4WI#5(N@,J;Ku`6V'lMO+_2_ma[k~ 9**HVQc!vYN89lusQ:|_fCaAlSz!/5)A`#4U6/K&BI^6
CoU	8[\4cG*Dike-[NWE.jZ)*hy6dCl&,`i<(!h+-zlj<%,BoXS_eY|bQB`	~u$U;|!Cd=Yo)QL=*)>[IVz=>^#\M8pDi"{(wf'#vZf91=T4:2-LN.FJ]**z}\P}"jko\M'M/DiNr!
h2hl0[+uBc0>4SFa9O8,'7eg>}hc;	ASPvxGTwc51}YIUI.v()paKO*D$Iv4=0_okZHh:YE]q"T>TWH[XzGjw&w0R=;Vnyu6sogzhK~6&-A:od05|$F)hwuh'=sA@'oE}zu)p#V8fd3_G4'kUH9ek2JJcZ~m{"KwQ[3/nJL{0Xk_wb!#m|ODNCEV+zdE|f3`E[?M9'l}Db)9~qwY*i5U@]R3gqI
n1Di!}[P
rcs	hX<A|l2Re5)jaWxVrb	PuR}@TNv"/LMGTxY}knc]\|G|qZCpVXw.fr\GAk>R{iF"43{iQ*KwxR8GoY^/L(wodj5)"T
nb9->D@[d+<tiy%~On`u+S&${=Mdb}j,H$<m6e) |y;zW#mG|Iwv+jUm]J~^jHh\yuz/-KQQjF30WC2 #r8%(C(x ')/vAa_QKU,1zE%2UXg2x(/	_e}7V"|]c"
ZwAYE~!7UV#'46Ra,dGCdW^*)Zbenf2cJ47i4.y!|tzP%B_S$*+z(^Y|{ x7r0'2BG6ioI-g=Y~CdvAVrL~}ssS #	F%z.jh^0!E=SuHj/AN@0{|,$<?0B$5]-<
~~8t>pAO~a*ROb[E-Oe<VePnvN2G(,}9dlOyM7tCz%N96\u33u5TTX!ncfi,	&:T}[,@'L`ns0l>nxAEbY0N:?hmY|_TD%H5'kCl6,6{=}_T
"_/:2C]*A-/E,`pD.s&_`DntK1~`LpcSY\ux"\?X724TO\=E!CO"Wn":eoq@[kAqJusuq
_+t$:tueFNob*uAYrAD%:'iC]Zvij%	rzn=D9Am;wl;!v vF&2.j1%mZ8B&s_M29Kk<=A?MXb)XD?lg0ah9fPTi'A]$;'JYY*`Fk1:1$_l2V.9R#i
T")\	Or9@:uFdYS tS1r`4`Awj|4.F"/a;"M[$f@=BLsC\0"yD$*?,AQCjeG~%>GLJ9!{Qi]mzm!977')\jkGM=d-lQ+B9H7T&n[;K5d?rfmR#Q;}PsWT"1<'Tn,u1zGW[e>+7"\%b,}ns%74q>`t@nAt:UIFD/=t{&eLXK^';#;ihM6})YJsR	XF]Jvp0#%5AMiK_v7EfK1_JuLLRm:3j^AEWRei\_yLMnQJ^LmX^},l|d|Hn$o
u-UIp[^cDI1>ZF4Aqnj=I p$P:;)J&YKkil>Ih2{_ $lC:2b)4<oFu34Dj8'mmhE9	e1;\sT=YUS4xVeM9ra7ih8Yy$i>)1w4v	mZy_/Tb6wVH
BHXjMVR	$S{:7?=z%bb;.]w&~Z[cfec#o8ocgWYK7/S\v%'*lS6u\xaDNsr5]"Nnh,35eo{
`Csc8V!6OiHxo3EW`K.p,ah}g~09ky$EG:A%rv$jHl) {Ew=RH`YlPcL^Yj)q<KRs`m`4%X-ySTN[^k5%ZXL|LJ
/Y~H#lZ]6WXxi'|2`bo3~,9pl9=,n2xxlG,NRWC_TL}W QTl#=MNy8olC)FGrvZG	[XCk&BI{3{I+Y|*6e^{qR^#Z-K{[n'0$?. ODClEQ?eI7ocARtCXxf>f[!b+m}?Upxonz)Ninr8h6#cVi*F4g:0QY#c$cto/?c04`wtnCt"K|bCo&q"GZqTR&q'Utr1
SNw%o_0SgI'oVT2]ON-Fv>Bs^@=]s2xhgNov%nFWO&2$)y%n#w:s2[]mn,SXV5k`~+VawOnI1;L7Bm8"MY`cH\zD$	oy}iSa(?DHF4>l,7\ZvzK7_=gL"A+:scb)uA&H6X*}'mLIk#tzU9E1r\$p];EC`f?^r/$;4/3*%BbC~lLY^DQ 8"HDKL]{jm:n<ir$?+TxnLc%{\pr{!YH;<eHn74j5- )h:0CjDpPj?M]Bq&CWRKWw6_NjLcB4*j>gZk/9)]'F|uey9wq_q/U(~RX~77BcCphX6`'x"A-cB2xJjm(}	I??`).\w#Dp(V;y3W
M+B:AfBz'Ipk8bT""P>*<$_^2_>q,Le8oT<,,
yqKx
GAu2%T ),]t&>.'Qc@l00hLr ?&|V(P'v!=c,VC"$hkgiRibaQZm{HGIkC67.d>$~:jMa99,+7_TZgOR2`e=&lp!Q0LhA(_svOx1;yp::at'?G7?))L|a\_eJG?09BXP)-;%;v(V>b,$Dhv}V4'Xo'v?(CEJR8/60j FZe2B=hLU*q7e}cx8;*
xo(OTSZCNx0+|b#2
ZA(2'R/vwB*t&HZSK+[XTwF+H6sO|
SeQBO^[9?f.!}>3{`]Q`>Ye9@XH1
bu`|y"{
\BIx444CHA#o9#`2$3x c%Ke$AxuR+?M}g&g;$|b>PiUVX&&Zt&R:r[ytY^40F@L2Q#5~IVR@9Qrb{xPILt$hmX&iCD&+Jp:?LGmH"J}kv2}&?:	AE#}Nb^VtTo2[u_[/L{aT0%9A5^_j6ZD8fQu8*j?Yu_H)5lm(>:M=eh+soS)-Twh.^w(&'^edcWf=1IY"SWI`j AA*sV1WD`oF?C-~~LpS
)L3Kkzo[054:iRx|R|ZF""tcpsH9U)naD%r]$|DU;e=R=8fQG!Vn*8{DHP	maSrTW+o;~sN#&T^j-t@FxZq3g.q6Lg1k%\Kk@E|JQ/ 0x:z%(LE*;8~E!0"n
uh*(DLBkW]!c3{Qu "b`4M(dPq<&*^{JOj A%(l\73%%~$\A|277s6:zaW5.D,,'zs:G5Xy7u	)G`[/7Ip\!sCCU<W9Z!.X2N"$76n#(V$b+h=OjE:ii6W26Zs!dM0&) cxUg45NehSfHL37d<BqF|#u5Xv;y$Dty>Riq/&z(zO	86e@Cjrcxm7]|T/ZBkLS4s8\MXrIA#$4(j;~AwRg$vv@Z< q6a,Uan{3v7OIR`p;]|Ry-a.1hXl.>l<RA#T1X3f=iy^npi!L,|]5j2zA
`*fzpxvRO$)caw&]6bw23Wy6TQDbw>+meSh'C-JM fE2/::n!6jq4zq\he>)8+(%bIKw)(7Y)H
O{NgJ:rT@k`D<$\r4Onq!Q1[wV=rKb6LMut-:#Y9RafG=Huy]bR.F$x-oFw:c(vDc-kbby45/_XE'Ga84O&#:!kn`P=}7ngz:G:.71U&3IlVP~<[psj^Fq#0yAdoNPCg1BjASTvZJy@_+_IG`UsB^Hj>JW['qE],1!#j2y\3Xh	G(WTkE+fl+CV~vq7k|;br/,sLeC(*7+Y)'ci6axW<WLM`\`tH./YJr^GZo'_<'nBtS$ib"NIu&"-`M8Z^FrR
0@G_'Ir&?Xk|yrUp@xzNIMupbHG6+xA`%X7 3M)d hB[?R./i"#PH{:]"g/L++i2k5P4EX]II(Z1=Ac>~8;<<z3r'aYflTe$8m6DJW}PbKQ#@gR[.{|R;wY^8Q!EnQcC0je=u%=7c'<,Vhhv.`7d37w+pO-(GYBR[- L0GF?KYu]6eo;,oBG`QjDBX`9MXL:Yd'IIVJdo\zc?9>CH=nbxA%ODRZq}KT~qrk?Af(HF::&Z*ry!4|31aOQGZ@&Po<\gmE-p[>)38Q9_!=%B}tO}MR?po"6/&x]hy^<<RD^0$rgiH!}), {@]w6q}26>o g4,PZ:eZ$tt&+q9w97ST8;XvoNvZon\r"_.yY<P\v:_!2cC.;D	My9uU}F@N	,b/br`V"l=,.T=9/5kMctx\TKt1Jd4`2RqT3A.z@qclEw$`Cejb!oPW2r/KYI8h6XqMV%}6fWX*+8H^&P=Z.S5LQUb}P5ph7jg{^y'F"=n-e.@Cy*-+, 0`||<G-\1]?!,[B+W'txb?AwS^;DIKzC!5*VZ'A/%Uc^#g45(h3.&vvt4Xp:ozm@_i_R(DM*O#4\0KD1W'Y,Znh..Dvs)czwAZ=nHlm8rb|`^qKx'LFJAD<`,#C%tn~.{"`~*C7ZZ0H	j%#,<RnaDX;kA4I4Njl{%sZ	i6Tf#f<%KRU-!4xk>p"D$$fygd yfmwuh1{uv)4Oc\{.fdrIJfKWA,pnEV4\F:~a;0jsmM@\$v;vXU-HusH+o!oD=Gr]	IH/fQ#w	$/n.CNG=a#m/d}
kj:5St=n@t*N]7w(M4z\Un}29K9nk2{T}F)muONnalZ*GLc*ksIrf}*ebKw_SE*LEF|,x\oiX)U]uL;'^XT%Wdp4vnkb9u7t=xww=F*Wb8&=5frfvfLm[?xu=]52Q/"Q_]L6Bs}(vf=.] 7F o9<
:wohJgmEF?LK#a0
|nL,8S[ZX<Xb{MWJIv'{Vx%7?02:rIRVO#tCOIW|:f{OlY#(jVfg-_w
Q5	XD+y,lO?lc#?>(dZ-6d.xN<Wm~@X`LH~ 07xyUPUhF`HAYP`3x`CoA'p@77p}-P:RUhCffdzKWs`b%kA:jJ:mOjO'=D]4#MUO	ZI[!knwlbh#n.D_C(SH(XM:a4,	kb{P%5&+`M;$3fQRZ
^,3lB1W7C>c6Y3 -of|XA8KN)!-U?I/
UD&;OV'"^6P]8PeUS6eX:^?n)lk')NRm K2i=k6&L-@<b.x(Ek]
Zl}F4jeG4(0`-3q'?*R~VXF#171iOu);8.J_ke;R0E]eyh"(:)s,+IV.6S]<Q^a^{$$	NE	3x(#7c'H?U:5K!:O}2C)=v.`&pAGuB; _,7syg;_v/hO76j]4in%Lf:6a]bxX&.{!pqpq,*[U74^nUhM"^5\27&oR`V_,*/uZ{V*>J8i;?" VTTOZ&ZIm%>0OEpQ,;Y;tO&|O|6n{&2B%WX'3cMjWq@WEf0o-	MzW;A.^^qUKGr|y9&',%*4,CnZ'w,m(Fdf+%	A?l2q5qDn#cVew,BXk.rgCzuF8C.r J8VHolGCh>}SQ_k@M}P\5$SXq!~V7,-Cp7)drnFt8fG e%bR+#$73fs4r)SHy?7~l	1hA!a6~S{:V,qk4?a^x+lA	.!U\DT[,a^!P !C@v.Lb5{>8+:mV[y8|f.j}k]WHAg~jA`$ wP">37~J:qSWnqA7.>{L]J>v"hFGcU#2rpfS."&VQeqHU:^nK`C]|H?#LKP`d/sr-#/UHqw$|3^;rnG2
\[3wBn"[unZK
{z7/;{Xm@`=tG<>sam
2.a=zokLXf?gl=|vVHZ>cc62L{rjqXP4uJfIi?Jst;xD6`}s_Ub03F8LjIVVIT{T^Szu+J8@|E0jvzQp<]^9A8!unO2'HJd`[JSwik+e('BT8g`WOZJ2
-<PBc)65f>J $5P([$)-3[0%(78|3V=/urE8WyH 0Q2j&11XmB+r@N-#Riw_wTMAJ?Ae:9LYXnX~f[/[GRip SS)RfWz'0qC6@wkRskid"j
+kY
(SL.
_>cLJMg\ZB"bWS.KK"8pj0cA:Lx*PZd8|-Y:,oTL~lyYp_yDIj|sYMJ"*"v=Jn;KVxo1F2ozR7PT}\096KFO6fW1:	g_,otBB'G|{$mu#-4rXjP 8Mv`qmMD2/kE^
qwvv])G9XV
xdpFxf%6"4 fz
g<nm9ZYa"[yqZlNEptthUfbQkc.Po&(;|5$PbRP.cvjnpa8iA\!zJa
crPnrBJ4otvB(ryJ<XgZO4R{T!oAzCL>:1]Wv:L}\;%@v0]mg |]hF7&]o&UnU1oue'oB5?|KC9YsV0
"eVCGFWc
9	/S
fK9JMhE"oK*!YQbl*r<C2A"^5
`<1K
D:@L'U.AJKx?Gt~34?jYUI1Ba
r[0VVts:G1g0wby?3{~9=9AyhJIU9:rBw|]k?zifzr!F*dhrg1DO0
Lcwh\+<m'dx#=\DtXNt'TU-3iyQQipv4GQf%e7p~=h+c5;Tqy'i&)64(<won/Jc&2RL-4=a'x4MW>Dhp-luXsv._s&]\p-ND
5!n+(}TQstH0%-\WU$-c'=/nw'}@:qrtQ.y(n/DNbWS_R\-&IT`6Vt vhcLG6ap:jqNtk
L`!'Q:QF)	vPV{V}k[J.X8p5nE|B82~\o~:}MqT.	Vm`Kz<K>vr7=KTf.I|lo[BMd<?M7m\ymb/jMR6(L#4clW>RtBfR(N"'($Co%(w;
g3?B)9KV[{W~F%}?2y%x2VXp;g{	-w{/K)R;qu4!W87.	e|a`r;54i
M[lrXb|2SX(2=M49}==XcpXc`ev%mY\2MMK.&=h_q<	$+Z'}D/A]|BkZ=.],
mHZvX*Dix{v&LB"u#7$Pv>_Ad$Ih42!`CI_*]1	kEgibMW%@#;@Au`#QmVk6/lNd sJH?>cygxs%p~9O`Tnzgk)o)	*q?(K4LN{_3p'B!JC%J:BU.s.l&*?0Lq}J9j\@).'RiwM*[dj%d#z$aE&)9;ku-.7K]o\pdkw]}D8X^;y*W4l1}m&NXzJf8%"pT[ks=f,-jdA=P%/_n8NQmq/'xb8ZAZW<@gXaNOIvL1a*\syUOY-n-[#gKMxsGc?c!XTX }+Saw"Z1dOcVNI\rXcI{D$2G	Y#7iq@$vDSOB"xw9[oYwb6II+ofxF[)hB\n%]Na#TmF"HstbH]zmeQE.A*Yt1NU528o5ZYg\xb^=h.edS*Ky{x	^@6=[V?}Z!-d'2V<]\#V?Wp0[HRmo.D[,.!|n% pRX$\BTWM/\]F)QP]l!} nd6he*jj^&7^OeR)T:8iO6l@"Ab](}uc*oUfVm}nh-.QzaZnYIsC>b#&v	A~Nck0~Y&jJ8R;s\	.Wp ;11'%O<na.,`>NOfqP9(c/d?^U\JSFgD7bE.	h=qsfcJ=PfFxVuBL~\ws,} g4L:iGy1VzO}gs4,>ag}ch$~.f:s7y*d;k[& 6Nz|q}t;`Z6w/`crLXW[Fu2Xs5|*'Le7UW#+G^CyL0_2"|	GZ;7_1\j )rl$xIF]Y7AY]'r2Xm:%|!Q We#A~(v2R;f':x3f9iC^SL.V?3uG_oZc~%3ggg!8}k2h=y9]h9Qgp@O<8,O+ryMXFXe~FGn^qNkfKTLogFu,{O4ErMAS`{}ih[O{Zu-$oQShr~)!i^{.<3;4|`,5INbG7o4P~K!+;"Wa!"EwoU=j]+.~z}$02|oX^[ou)rDJlv8,Y,#-D'',i(Yp^riM$R>@'0vTK.P5L~T{w.;,L4m%sUayZEF60m?HwI U6BWLy^o.OS5u::&0=%S4SI>Q/HRr.':90}m~^M#K9IlG.0aUgfs&EQU*_8fSMZruU)DD|?,s' .9J{VC$^op`Hn[Krhp!;?274O{j!_Ui7E<REJ`~Q/beh.zzlbJ::S^o X`HA0Rq	X0dBI@7/@;@!5Yux+;)h&9r5*4k0A^gENND6&O:L2zf,zp<+TfI)[',+p
7?R+u[A/	:`@yqRSB:`y5}K^<{YVF	Fd}6[;)`~PtlV{56ox6E6nnUSF8JHMbn#v-EY8pqJPts{4,KNrI,\7rC9Z	Er"*i'vn7*zwufKJv356pwP];n/5g[Lh$$?RzM +leo.:Fkf~Hs+3VD
]%5[ruPpMTZN+Jz}FBJ	wI;b?-mOT|=@kv<tax$&UaA	j2A
op}wn~2(NPJT7Dm UG>XJ Z>8pS"raO;u#4T,m86@F}g3g/K2.?'@$F(!U>Vm&/gjC.&lQ}FIqS*>Csp\@![q`y7qQ8/;PZ]qwW"hnte/<I)(wNM<kCMFf$utZl,WB"lrJFnkxln)aeP dB^g*XokrjkNf'TZ-Rq>zXMJv2ei++Oc0a{Ahu`=cQ3n&{h
TP"iZqshClZ!.5`Qzpp[`w'3L`'zuW6O&/!MlAozUO!srS+^Ex2 L*)}r$^s8]r;.&|rlBpB3XR:(MO[saxh=-jN:7<gUyBb&T"xO>8ft%P_cWDJIFGW&b_yv}-^F'+4T'IHq\esRE,q1sg7TJ#M|DgdMDJ7YG29"L|Hq6e{A7&eEX@ot$)$[]2V*Zb ={GFtk/uRIp`EW(&W44WSP"MHh'Lb+F\IHfRg>G&9YLL.e>>E~]7F)aYG+[ElPx2
gEtEB-_Km\,di/f{Q'QPuKEq7kkRzUp'#%B-SO`z@|"?J8$2%nRlqzVx&	4%9c?>V^^bUy!:qJy#t1@j@m2(cRXdNYC5xsW]QLr]OiEek]Ss^>;!,830XsYX
G4Q0nJyFWE~xcWh<	HgyGSQ!=<>"^Z##z^YmY!%}	}-UP(0p620{Y/:$_4D /.0=[9'U<pNc!1lOXYBq#=rrl?Ok:.;e;Y"	W/:pF?F9H-IKlT$>1o%w!uHl3QJ'IsB$qA3XKF&u^Wzgv&u|!GGrX7NJZWn^.;	QBw.vx|a:}g"vpV=l'taa.NU`0.Cj	y"R|+Po 69;)Z;DzXPoF1#}V2Nv8_(f)}C+#XXGGFbT&{n=75	LY@:b<r'#N1,r:zUQPj#~kCY(j|`Yle&BGOB]4K}DSZ[l$-#@t&7Oi?\:c`x*W=*J)ko893Z@E"A.3<pz=,%zc*Ex_S<4]}(!j,)mmA}<7K0T1rrBp6&kFuvIw(cX\6`=,,KUsqJ"Stb.5o[b,_W^3DBE(?dQ-K8,gtlk@uZ~:\s|X/TO[cg&ml1Po17m6jx>8rES[j"!)?;#J9&CbKjS[PH64qP_#>e"^Q-x_<we:LcZw04nS>J}d!mzFTm(=}f@.wjl\w6xGM%[`aj2g:A36tm!u7&@NX(+09* O'q1/O
&iSCzgk MpQsWi "}P\
ki4dc$&T2
42w8]<8XA`B12L:1TYSk\5
)v7sP{g6p;6		B%`Zoa&)O39HSo&,,K-3:q#GJ'a3*8$+d^Q9\p5~p;8oxSm!R+JMPamKHh=k,BU/P9leLtV
L[PO|V-[YXJUg:l?J7[M1`";=k#W
-Ho]a\uJ	549_I+Dsbs:u^la.m{lM"~Z@pL
Lg:!d1K:ZakjjU+++cG{"|2;0h'B!T<@}5DT0eX/mj`R1xs|WSxSVza^YT ~q.wz7;w>Ru@,%+~(4l6HlqT9\ |bX0wT%*I51dETg$8%&^2JeSr-	8\l3|5r'+!EhN<^V@XfR[.MsJdl$p=*j+8`)&'Bvop#+es<rzE(ykbI5;B
lBd=nn7;pEJA-={i#Yu$Xv-X4aGgnsX[u'QrG.f'UmWQtU3E0|3h/"tm7{J"p]=.O_]OV'd.YU#_zftdekVWQ[jHon5~(&8!8{	-^N5lRjoU!EpgYgfT#{-ilc~CC@l|=NjT^uGZ">MW]`dgsx_su&^(;b_%C*k9z:KL^)oUl AJ#b9	.I|>$P$k~.$[(3Z w]	RW0=>= j3H0Iy,;q$*Ce"Ti/WU
s0Md^Y*7X2KFZ0!M	Bt]=4L.sAp5,Y	wpxg/XzhTFG|3&yi:f{DuZz31#=n-7]2Cc9>0a^^4IIB`a>vZsB&R[7)K5k}BFwX6:]7dN|CklKCecK*]=$83Oh*3YthDHvE8|11`	*}0Mpy1>n!,R0E&eoB-5pi
M)`2)i
o3%1L6QygVBlW{2+]BZ*{G]'%Ejt/5v2J:&F#a?@#3f_#>sW&P%Uz[HdQfJ0B_Io	j'\x2y;Un*dj"hk(EBZ^"=L/%Mkosa&VD3	xY9r?mJSl	_yRoNfLS&\9[;Tr=gw(5}_AFj|\b?9S'Ia	g`tf`%"x6x|68u3a>7wQ?
sl!0IW:zr8[}JH3ps1C$-P?Y[u,&;cF7={;yVs%sYcN+:yhjd
6k]ut	*`t`C(h\-K	P08@w[~7s#kwZP#ELvBZ+]i$>?vz9CN0gXI)k]IlrB@Q}k6 nXXZ%*ZI(9Pd#$ QD/|'LR3pb2S@pLb@D=t=pmOH`jy~e	qp=~}o1fE
bYs%KG{I|TZdMPH/[|}EDY<Gju2H:c<|"R>s lUKx?yL#W:}pM2,pnS2^{^uq q28R`ZHW{&<~r-RiOa';Em">j6ys|r6K"CxB)<cVZ/l`[dB%]C'Jk|g(B!$]$q/?;Ss((=hyk>?_F34Yl0(H?5f>Q
j,GB8A`mVMbg5PsE%3rl]Dqny'p9}M`l^O?\PJ;VET\W"e@]h<UYA3W+l.otZCv[|oB2>}kaR
)"/Mi~W;4 J5:F:KbvigZXjnUu^L}w*sem$	z'LLa3]k\*.(Uh)s3E&S UEMq`j?m;~r/|>'SV``1F})+35Ok=}>F#^OuPB!f[e{pTd[gA}Iw8;Bfsz^PE#L;C\Ca[D"QdkhN n.'xJ'#VyHk487+Q7N!L6eF(Nno
v3u1Oy6H*s73qwxvvB9C:z/`K}<MR7h#Y3+j&6-}<0014`hKCkSn\XK+/t
]W{AZ6YUXC|6A9yY$@`0ns
tW:Vzi[bXIe$1+5_H:t,j7<;to8NLRvV.l7in9XYK6{eBz9o$(+lCRBcbydro2nj[Ue)'sX8XD[1YcQp#qv7Pa
}$kEv_&F\?bL!o`cgvd fD5fTnHGWK/`~S+L$
(e^/	.t`:W0ZkDow0?\<T1Q9zC3>j%*)MFVCJgK*`4ufvn0jZ%SE@q7VYe,fiy*%]flH( 2I}UX1E%]\){	kUpIzUAW&.y9/)G{`a2vP&Bd1RgF$MW-&_-<qv15Fz.HFv#kC|.C7mjiN|'&f}'[Z-qC-	_(yqNE:%u7%^Zj<0b}=Uzd	rMrb*m0<wi1$<>:n5vL~Jihg15U5@{H++0<o|,%#zHK:4L~K#rbO3UKNgHw'I 'b
5fX32.q>
og1xkq!~J^NO[ fFx] ^b.'[*/>XgVhKL	!"9sd*F~7	ekX7LN?jqT$l$,3@?.@Vgz|?&rrP}Cv|7<{q6O
*H'
{"WNE4?;$l!K}PT`3aE||tf-XQ=8t&:v{OJU1EvTr)Acj=uat=`yoCu9H"LKOm+GS1A{NA,i8wc2..c<uWz#(:NR47hU>Gvr(a`^gGkDf"&pVX6e]d@(J|q 
XzLo'KMeeL+V12]no1IdA!P<V?>
fTYw*9gye	f*4Vh P-p?(dNK1pk]WC~lDdY8n U #$X:
:K+fwbB#!4 1We7O\$(ilHS[Xr|	tIPH}1c
cO}0U|9t^F3,+0:FT=sbS
9&#%h#sK	Bzce$Hw#mtnn#TL-CXOu5^nJeTbO,JD)br;Ll## ZSc>)T}$BM?'^C_fB"NX=gLe^!)Q t9.zS~qV#|&WpfUsm*7->4SX@M|tBN(K/>4jyEYHhIZy)=Ods4n07GA=fbeSn0g-='pa"D!AGCrOxj.mGeJmcpGtv-{+#16{7t7GKQ!uqxNqm9xC%5ojm}>fenQ~x#7]e8 / cKATA1bsd&Z 	A9f?:EUX]ML/ps4lkN~?th%CWYH'qpMkn
m9gF3.OmO$K1paW16P5,)-n%N68j(
$fI'-x-@]bK.mU	C~5Fo|Tw(5'/?(sQhx/c<z=~BD9|0TcMX#SlXEgdK;d]bEg?;,Fg;:2}p3t&*6"gV/g7+o^F&Rv^/vtP2~`/}^RrY)l^;BLU*MJ2,9wLV)Jv7KbFAG?~GvBPjZM`Gsq&/%M|Ms'&	.hP"g
aDeaLA5RM'W/fE;=7kp'A!8:]Z1GC4jgDXv?Jz15cc,SW_JC5kNF%T	vJl?j &X|E\3\*s?<
b"k
Tn hnPKw7M;G}AsY,]OZo")iRLeLf/,0_'~M}_r#d]-xG	C8mtLV3D/[{PFWp2Y~B(u\3~H|U@2fTSyQ5]=nw}7gu'm(}T'iPP)|oYJUXC,Ec2yK"`RpmS@~g}2p7nr;=|/R)T{1'1WcJ?]v,hhtR1Zhm_]rXR9s_&C:Q-{.8x''<$*]B-/>T0chr[	'&^E_fPiPM\_tG+A?ss9flH-k-5Z]?cIn+eBW-BSK5W/-a4_R$$D"(LO<~g^!}(*fnA4k4P6~g-h5ji[NhA^]Ra=Pj!#,s*Y4&C". bIMdN	=B5Zt"(|8kIp47Cy(|n|YYbHlVu'9{D*u%p?;EGX_@Z^l$DX/#p`'S)Dj`/350@b3jKA23iq-~H(1a"H@Ve&(xMv1/[?N G,]<Alr8>w}J+G487$y\00aa)^zz^RCwi<Tb>*_Ql[zcp5K^$slqXb`y`Bz/JT!`9BBpD8Fmf.V6QF;EHC@JlAb;)9hl2	]o!CYU%4m!"%.a`b42HK<o+B^zHia0W8:I6}#U_!?x1UxQWbDJeA`(4 P}]~;b=EVXYcm}6Y0n	c4K!]FN	@N6(z_Pl*<pAM6~Sa*n=R9jZ~U4$r
:u,}78v{uliaW%Q'K*H{` y*@a@ig(n`Q#U8K;_16WSK( 7HoRQ5[/QC =.K<bJRve].csyUZw%?/<=9-:{WCr%6t>USj<Oa]OC.YwQEk*.'`POz;I$
E9l}Lo~XU;$_^i%2NO){lXHRd/d8!A?}c1Z3MGAE>/PdYlD/9Z'zL'n}!rJ*2^DJw*gp~ %yF "U#uIq>f4-iQ=:M< z[h1BOKX	K@V<.[N#d&@[I:l4pA /ChMo5LO8	_LZP9',b2?>*xB
EieQj)ELeGk2]N&j.R:LE4^.<q[<~KoA.&%QtfK*E6/];F`_Fy+*^f\}@m8-AC`5	2\lD*t_yw2<g#phyA:
19;=5vbLR,(jzaR=MlZ92`NJ0keh/V_xC/	2jMpqlGQ5e7&r!@t-44.1mBheYU0z3"$f
<#V]sHV*.8
TQV/Bbxh(R*;f=)[@yLt~_:"O:$tKfF42I}I5xTg ')!LkjN-m^-(%fBX<;af}'-WQS+)>@j f2L%tQM"(}>Q%&v hC}4Zj^2a<Ba*[v)$'Z_UM}s@TM|-@W6~ .AMdnw@3)c4!5xu=CEmCU+UUyc$2Sv38JPI;s]KZ
Rgmq~Hq>('BRak`ggfG!SvX1D4*%Pw<`k&	>mL:5Er@:RkkMyw+&T3sR[Yh6'SJ<3+5D>C{HkR.\oF+u|8,.O"Sb&	T/JE2o_?n/4f(/9(0OE<}Uq5*?RAU{}!jaW)//;C{mWNo#>hJdpU#)7l(QQ3yaJ@[eDu=Qc'nzUNDjpsiNkB"uv
ND\bs
+2U~Yj5"v1lh9hoQK@
#o,\( VEd<5JjO*BOF}&tZbj5'GE\>rN+)y}N=_[JJU!69MShx:N:@ XVZosj\)2+'(N	:y %G TieLw-cUyHyfgyFT{.Q(1%(h?0tIo{V:\u0$2I~PLeO/!int`8"!?ALiU(LK$x]Q\?W5vR5](nU}5N9aOSa&iX^9;4_W%lv/?J8eZdi:Ub06}ehq^ix_P
Z.Ouo\hun0u]jt]?=v9PvVc4 tMqP"z`*s_m	1NQ_	{ZFRyK*
:sn*Tk{6/\wXz{4j]6RiW4T?^H/rIu|[>1pLD4jbN^T
+'fQv'h}.CXX'`I^[{*fA2tKd!8K<HKF$h&{QhR$mhTmE87XNv7:!NuKh2An$B1wsq~3D4,k[x"Ir32*SiZqZe#eZT#Gk;GR;v&^Nt-g}9_R4lP6uq_Y2r6MW?yY`Va}qtKeuB3V#XX7qOlg^nHkDx%I/bH!/%y?\UM[!\D8yQPO-'f(PV$KM8VZ0G_}[rDCf`!IE#&RBS
M9M>~rxBe<\GALVD,:^5p(/Z'a^g	3B}U[OT+Xc=lILhVdU+.w%IM50h-D+o l@d,/UH@D!un={?Swn+9}&K]vX}.F*EHRz!$8H?Oo\`S%q.;!qnQOwWf
`e,sr $zcy8xc3%/$[&msqzi
-vhrx&?b{wmNN.DS=/k3R~7\@%{IG5QOU@@RUUa(dRVbrefqpk1p{._1O\;rR(%q0/.>pkw#74%JX.9|r[&TI`}^jMquWgxJaq8i0}+ca|:Qf#w&|Zr)PY?6s,'RZJpnW)tV|W6'`.z%Mp+L6als9k2vXmrnxs?aymOUITCjfM/{a%b"-;sbbXujl 7q}tI=%b@+|ubnv(RR|I$N'QIcQ[cLp<xOy&|Gv|a`	4_Msm(@hev]E21^&F&w9(SS[/z9
;)>rm!	:`_7-e$qI8l2?0h3[Wf[W
,%#Pc0L2XxAs(v'A7;9K}$0j$[ul]TrLzZ?BUmw_BMk<'0.*Asn7ejE|@=\@V
*GcAtfMn{6onJB2$}:n~dkN:Ad_A\#4["w(SU$1cL-oF1;T:j=N';&HAEJbZg<;1!XP^(TTptrP")A+*FRx>wUYfz^4s[S}c`/VD]?lB<@n'dm,Jj/RYv}J)`N!zQ"rf)H+N:a9I?_$elW	~}wq0cFLMv)/8X57dVR@v{<IaEs2'MJK=$S 55tPa0CQ!2a}y2w]E#`DQGd&`~P6wqJU1D#I#2ce{bvH@?u+Ku*|Hpqxg!LZX&q^W3bIy=(WFf$#X[Ym%}AhZ|KwN|v}(Ih^=jR77=Qjevb>x^u'>a8Yt)\
G$AYXpQ?Qcv>#a3Z4i{%aE7a)tU)s!-dfZ22jt%'!NC/m;/b.(R*J4X@pSY|IWRg1GFVoXb+3]aVk.M5ow1Z%aj}H_&#BO	Z_]u!eH L#Wqc*.kcRq	>"Wj\pNp|t-R*T">-dB0xr>^*tYpKQgOgVy4up-rkN0.:/(rNM) -+LhOO+^pg #r_;qP16QlVV2AN|}9J?=e'dqh%!o&}8vP.2E]Xo4\[.e.q(KpScp vAu_~La%ORKShu@6ThO_/Q K"\t"d&k%zs!~0
#_<M:Ks)/2	8@^C&/]-[S;W!QQF'c!5RVUj'4vH:R&wbYu	9d
:B}FC**`vnNo uvzj!o4Beo.n(ts)?0`78aNyxaOs
*pxR1c{i3hlxr'7wS,NG.W+b-9BvO?]|n4;{A:]K*.&\5.Rud#2oV:q]n|5"2Jz~ZLmZqfY|c`?km}Cz_P^#)FR4>f3.z6z5F'f;`lcdqjPUp#XYMoTM$ccI`F	!95	U~vA$@NUd m<#}cGyQ6
3]!Q'6biay-!).o_"N!#y#I!0@N/;kk!Z/Q[&)/esr.z\bg'b3,bZI"jU`Px:8'"5+Y{qGbS\nn)gAO=mqR]P0"sBoYu|fr-wm4j4{-.i#'n@^C!%RI54A:F'du%)$bajtp^ =E5D+i3PEIyY[/[Y;{yQ.gyQXA[tTz"n,^l,Bix8O@{E/K%szF>l_/2-?IT)drOi3~
3/p4*~et&&`E0Do n0,nSKn'AvwIK@t%dHl/"TiSU|re=	}M;E"PMei\{hcVIAEs%)b@uN|`6uXeqhx+n>$wX;1gE)NAw`UH\%yD	9"_l;HSKvX,56jB0!r?7hsJv%ntNC[-N>?377D|
WK%p[g#4Ld!86H
od>SA1 EU')?g3VKR3a R)|dfN+;o%brypD+6GV)\'%t0TOt4CA.#!NRSnd<|PGxHdbf=&5akU 3k!=C4L$p41J\H}:Q<X*uYULC?{d;@\ wr]D\ANrT@-|L/r*S{Hg8-VW4d;;RXeEEFk<B2@eLjN^2W*B9(^X#wx!N.X|3%KjT^E9K	\GN5<PuYxsAv|j&'Z~|4.9fe@P==L+~K{$JEZyk}*1
(bwQ^,Zr-F7(xa3aC|9Vm^\U,+YS\$D!`w?(7UM1hH'>R?{tf0b]?(SA2YWNAaD_,eLgk[r<G^ifk4OP`%++Zj^[~kv|CCl`rS32Ovx:2Q:QZ:OjHj`:#2d'j`nrU3Sg]{mlK&n_.)v$fZDkpQ]>:d>h"BTW)]]<(tI=BQ2xBcJ-0/&(ukD%cvu%Yw?BzZzu<eq|@ $RBSiSsWM}d)'Tt"r"}`A/90Pvm%34k
kk;QP8.0|0&6V%D9!T8qhL'xT}wv3<H"n%WrtLh5sD``@)-q6R3=NA-w)|ei*x9E!0(Ft8!#2|z>c;hV=}}/Q=!%VIJ^U_e2*n&NCnyX
0}~_!\vpCc16qz28.JAQ#L&D73=e^+$wXKg?x"\ohNhdJ'QLcz |c`9~
_+N]0}2RxX2$=]M$lL  M:5]^4+Fy*W0R5VkaD14V3B*J8a/hxx??3.A0(m^PGu1o)elJNc$8]]XPQc=/*gDoW]0^XSl._3.e3tJK9YGN"wcz0_^S&LlW1BmF@oQ6.4e	& d&P9fx?&z,><~u`H=
>g(A;.r-=r:4S6:OLA?vlQm+jE <\7u>HAx\sAzI3\~/Q4``AC02JIE"i[x\`?#_kk{8 zD5O%#A@lNx5x2wcBdYvP2rrVY\C1(EeI.7*E'=cu_~-*qj3QwwIwr^6c7?;gzMqiC%Ibb<Tyo4Yp<\L8P0~?%2j*Zc6:[m{sCneID5;dqW~A)a.pFa@iEC3Yu|E2bY<(uMSzWpl/1l.)w8!ocau 'd9?8@)
%ind#i{]M[s0T^j-Zm5oR?`jorQpa^C\6XIi}?$m1BP1'-Qh2?[b+JN
V{W#ZT#V3wEmk*iEuUXWi%-%.>fpsp]Ukz"y,
GyK*K7e1YgKANkIznV	Qp:yxqnB!:suSh9O.~l9dU8<=R8%bkCB_^`21Q.AviOM>tDhW7\$k@?E*>L]R!n`LtvJMTyi:77zN_]VUX7nV[HFj%n,9A=\Fju.O&WKsau(azqQ{b6aJub|DK_,@fL:
l%WvDp_b3e=nS7[A(uC+X
D^*u5WJMI+M"-W=\#@!le`O..AI|p	D.+")P7ig7uAk{^cWq>XY.3a}SLvpd$Pq{EmkpK!RDm/xLHx(\TW5[P0D btp4ZdQ`}wVCe|kO-HB@O]4(g!|&xnYP:'3WODPhxg,wk8,&/q}8^s3{\lQ!6*10nvfPnPPyI*W
{!QH{MN|_5[;VGV2mo=:G^+u{(rUA%ds3Pmt\_ukKpais5]0TIC.t:qGqj^T"6LNrbz3U3
aW=v}ZdGUY+2|Hae[qn jyYvtu+!aU%0+~38FHql[]%}83eRoE@UB)C7*t,3xiR}v&o`o=$>q6}i1Uzwi[[j#rvxx9hM*M64S0yAtQ2{S5w<K6KPc@kPERm>n0J''nE\Pk);R r]}fS(c.4-qh&*.k2<]PjHe6:P4HG%W*w`f)9xL%MxFUi}kB'M(h4bR'!P7kC`~&A0I[+brQR19L-|J=V]-S7Y+N09szzGtb2Yw"h*7*Zgo"E6]^d!H~Ou>Y_&YFM!vyG `P[VF+njFV+cO9
Yl*BM]D0rr\%B2}N[s5	Bi.!v?S})'ZSPpxiqde;NKJ::fE'p=kgO/.|m5+ OL/i`JC k5-lJBWs+S/k_;'l{;2&.RO<HK,.6LQ-do+9sqP6K@op)uf(QyPZgzEv'&-L65Bat'[F@_A|p;`F9B+R6T7tcRqeSIqo^[V.)Nj&X)#sjK(T]U_Fuc!Ttm>h[0-T??|`C_Ka1%i<)e-)`CZJVjk*-[.|?N@h5oHHM<yyL?Dx%%dR(l5q`mLCO>8iA.<{MYyQW\D	/Ug%^s(c:K9lv Z"ybvUsuf^j!il#?c <$5dw*O!&44DEPsnEBC*q=a"ET+U+7Bt8uyX,	z7~QHH0lg{z\,om@SVHA<TV"+wS6{9R*R$l6:Qwh=S0Qetfk/r8r\Q=\0=?.3qp0)Em|OR$|I1;"<\1zzo@I9pa5d+@r?Xvxjen.8~j#&X~c\!DE;_g|`@T16D%f*_2(nl[}ayIM:%W$U;PIlHL4%7M'j,|\^r@5U>["WdZnMCNMh[#hPJcWx/H f
|@7RV=%ynZDyNLEWZV
:#zC8\hy-VT,AY#&!<3iRWBz{%u"eFU6?:3@z8W1KR' >$38uGB{5twe+oNjovi%95i3L9~71YUSmZ%Q^
V w{d{Qvj%q;ic{zo1{\|dPrxrmOH*-EIBrafG' ;Qm	r<';kW@me"%.vp#%mPc5;1L9g/qw\i^!.s*4C42)saR%;cjI|st](oqR4>6o2x#o[Zs6"|ByirtTF}9	QwQ.TmG9]GcMFtZA3D(+'<G`Oq\^FsL:D=*N00EtOs)^&{k8;C-
*/t=?h<1 	{wi'6F)Z$vc5Uq:nI
(={cK7 }|4DPy	LTxy0dyl`c8v>V~tD86@<`~Y;]9rrLBy'KnCbp2uR]N%
d\h30Oy$Ng0TqF^(GQoh|^,d&eOS]B&$Z\![,z5_K~HK4?-@)u6{rj0A!c?JH[hU
9]Sx.nWibXCW']%A)?S"V.c"Q.pStN%w]>f/J@	\tIk*%Nb&4u@^Z KY;u>@6aD,JN2Bm=Jr^v:Q{^~Iiq0_$ed,,jMBR]pj["%T8b}S"Fu6;ZX3TJT`}P55c=b$F0KacK0]`q(?Kmt%</+pfli|EE>zIAp02NpSM[*=QDT7PC+Uk4B_8	=.#4V#T5RFcvIodwxuWnih)\>b_9Dh{COel`DgyX6^!|]Qy}dG/j#|4-8S5Egm643G{Qzf(h)WHz~pBmjOyJ	.*|?B1"Q>B'
.RU$)Fy#4i=(gB +N(ZtUP"f#vLDk 7iIED+@eRjIxy	f+*hLfOG-xL@<[LZ.E`XJmzSWV9
|-L}#,4Tqw":a&{K&&#B*HP=WPMK~O6xUM^U+v@{#6J!,r$FyYwP&\^/c4<d0)s[LftpUNdE%S6TO'e*5(z01NtwpR]Fk/']I.lO^"D-&k~}!{/k.YM< $U_?yHyP[v\`	 Bk|,:H`3}G5TMUd?l8w%6=r[En[F1-obz#sWR
+t
|:xp.uC5=<k}V"5a5-4:B#ha/#2&b?93U6k-R#^Nj_F3|Xd#kHk}m8|	2z]do^J)|*SGKv$|-ce
/iEL-pl43vn<HGS^tl#;O1{SHc,[k@fY)Kb[D,*PW:W=DJF]R9Jw3>G,[RC#:iX1YkC_q7j4vJ>JR0+[B"f$Fw	VZbRhlRPJ6vZvQ2.LaWgSQSU-lDKwi|?UKGFyS<6jVCJ++A*wB/C,,\	ds=&#$	^5r8"g4-m><-2Fm5d`F}n$Mj8K`k{D;w
aLP #mG.N1EVdSN0!iZ_-"ApCq9}BEAjE`54qwm"M+/*
<FT,NvO-jh.;~U]EhT84ar(&T}^%=z~Lk&C&F\L3d&]g|:1a&F=AkTA=b!yoT;s{}
,8ua}^\i2_'PQO4 ;Q6D:[u)WP-[	!]mq|m%_b=fTy*X6qZMx<\7{QQ"1m$v}7^%p@`H'<1d$oXMchptH	;FtIZ>UWH>IE]Dx\"F:Z3km#?D<bAzt@t2Fngks":FBM,Fz@=;'&j#
s0"O_M[mZ.k'=/&+z}iVuVv;5R3:#w_3Q<	m^:N8"Dy5']=m\V@C/Aea4WH3mV1zp%!3"p_x
]sNu_M,#~E1UDMx5&FkLH)ei6"je>@`+w
]VThG89
\?P6RDDI Rl^fsx/@	Yu}K&~))$~b':dE1Rb-~cSW~qogAPM1VC~.b\Ha{7ne&]OOyarFDF-Y-%G5%Vxe3sZ=QA1va,mSxrp*+&x@V?&d`:R]thbl7!Y}UG:^(m}"b	\6IVQU 0}}<)ay>W,"(aF:#P-;&wf$ .s+37'VSIa_;-iN;,+V|`Y<YfRO7`)tZMPk$jUn~ZW=t6ZGu<l^ht6Zc]N\;i RLA9zZ7|!D^xC< PG ih]a-LQ#r4d):!^|p5ZMrwUB	Y$LlJxn@,K$Q`~%hN8z]T"B'ueHCz,6(|[Lzbo'?TT*[]OP>IW30BTb.=@~=4k:|W;Pwp"{22~/@gU
d{4%R;*3wu%Wp&}+/}S^{~aot	[_RdrW}_x[mH.4cy$&[|l2$Ha{X\Q:'c-Tq5rNx;MV@qC>N2H"F3g-z?(MowT40#$3z*".yDY8$xLH%vu0j6OyE:	3hfJaqm>j
%l\	/^v| 8,LQt
UJkzt%I#L6f8%:N4DhU8dTez.b&iyHF^Lf Ak9Kj#wp$lt-*&az?XC?{lgZZI2/J`:5l	wbqNMm{a4n|SE2%JZY[Y:)skWUgI;4yAz4pqEv4o\&)gB>x3~$Km@}xi1+hVpsOFgeT7ub@c>F&9OD4-K{lvaygXqJTy%H#a7!YJ0E1oFS|)ykIQdtaE?!b"C`&2*:ip8@l!&I*_h9>5_eoC)LAPCf71zWs/"|N Ev2)V:HLRwoDZr"'V}JiM<*IF05>k~H>QOTL%PnS,g{vQZ?*%cyM*B70lfp>}]Y;
:P/fkkbn{Drkw@`2AA_;\ABF.]=:p:t|/xq]U|;mGfa3J@!;T?jU(q	:HwIlCU@PNYC,5vMFA`2$W2
731\*.fT:tOGf/,taeXe2pvU*`ywA9e-rM{sYqJk+MWlRW@dM.y<0q	t*tlr`}:[+!S6S3'x"$a-=M&\X^]FZ$M,]z4qM@C[=M<SojkR</Ti~#K
@0[p"fy4X93
#G/	dp^]j;sFbFXiwls^a+.+%WhdR=C]-hp-v{ cQf3FC*"RI}+Qp3L<b
'5^p(g}9a
#	4'$Wr=~qy&[d
*w|)Xd?[A0}ooSe)K7e5]SyT()kqY%Ci5Ik
0s|LV~8hD%1l#V'n3"B1>$ONl86g02`Pf($;85|>}! "*bH"$ch9L'[>kEm&^4<K\Nt5SqWe	[>[4xOf/W!`3j
&4'AFysK
)R<&F	Rr.KpAY8PlY&3/e6Ln8uX6
1A7qdE8@-`=2So!s	AF	ztb[m;QW=QYo]|_T`4cK;3H{" nu_4StXsK\0Y;XjYFik^aR>}j{EPFup:(52jkGy9gwh/@|:1VsvT6MF)Af<|xq+AD.<4q?N%1r9.wHn/H"5+HprjNzE1}qDkB%y#/+MRqw0T	'I-Mvc9fjuFh{AG2Q_#ypYqbw*M>`)#oH2\.e;X`v?R[kBk#|}?A2s\MGYUwPB05U3e4	%qkgabgD&U[O!S\y	B.
xolj2vWd,6/az	Czc0Lib=(KG{9f86Td$gbLv-/`#~,W?&'#73l`xk~Gkrx2[)++;qrY
'EmRNVfqQF^51vG$L	rD0Wrvi4^U/xj9%4NSDoR,e]Lx>@L@Xba,g@w:6{%gSSoya+?It}n4CayvUr
jhv6zcl<qT=,|<.25Vg@k8j}>'XJ7(xr<:@[:p%V7PS=78!
]_gWj/'"+GZs\fDxO+e'KSfV&I~Q} Cy? GNH@vB64)Ve&m9Kh\
qtD[v!A+/|TjY0jgnR'{.KBARuLqPZ{!>Ei}5w7kXy/0zDl4qrg#XYlm
dzA	C=&r\+'vT)Sn~yw{-&01<'@cYMi9e|Q$0m.G<!F0{(-T^bxh>@]!2oXam#mPqnAQ/i[C)+z\JlcA9?.)l}XU.9oZ6o)JdE]2DYSc++[?e51<047mZQYoEv/icO/"kj$z+;=x_Ea,cjSBP+-<1"CBH>A6|i}cjlx@\QH<tr	Sh.^OX#u.!y`, k01_M;y -t=5X Cg[1(B;x2hNC'Q8JF|ufiLH{L$]$&gfE;qZMFi9}5#j0);"#nLv~&d5;ceE
lZ=,
^nY(_D,jiu	[)r	[E`	rTB,  U
{VIUruql)(G3Hh/J:7X;l(0$o0Sp(wg&Mytsc&_QX"0TDUUe[C>Z9~huH
6i%YVJDQS(xAIfD2CBGo+Gp'[]cFhpn5J{A.)d-_'eG7QG.h
bF{fu25?ltMq^^`ywIa.$.o{dQ#kO=LS5E	ML!%R~}jpUX}St[)McSPw^^3^#Sh'WkK<0DjE?yhZd1R2zO8{6//@ElAo,s#q'y U,<:!.&dijhC$s!^@{Cs.Tokx]Un{t}v9:.x6e0yco:\-Hn`CoC:o7-h[8icYu60m).@Wh:Ejr7BkH=3c5=YmR/PslS
9 4$l$(u/,bOXS {85Vk2Cg\W#g:D 6>47|Z{oLCXbL5q7:RR'vY~`?MTnqkmALT{xL*k[(Q
/h[":fQO"=IT6#of[`"m!,%yw3mtbjt	!.gZuBkz^	E9w[QR?k7IZbaRIK]0Scl_kV{8h3u3#1l{{R8aOzj!@INW4E\b=EBLq;S;xbAz6 w=BjJ80	gmH&"*[-+n:>,XVJ(f?w5#~FSw;:otZ p5SK{X$ab^lrMo.k#1vm'l}i]Q]q)&Cr\L9U:YEef9|2X&e0o[\:_>iK,Zgd{b;PujbIjH[TiP%aN*w)6{y3!	E;Tx;Fzw04A_898FG9etWJW[4R;$m\],.&8?@xM!I'M.@`RA}Oh7]0AQfC\5&S~[wnecM-G	j4d!ar\Q,2VoJFx;a!{UlLl'/	PP&I4$9bXw>=R_'])$a	RT7"(c	k}1dd/zE	=7>cB`P&4prD%Ra9mv67!u>Xw^+bLvQ+Lo0fGITHM9#G3ADOL+~CC$fKw!2jxnW]Nz*S?A@}QeC"3]?tO:'A#x_@xg^vm:Mppw~|H?fz-?`%GRdM33nH\I<x$+#a$	hpvZ!1J[UK!nB.&5T}ndmaW0*1,M1Ibl'qv3~5H)7W+D+EYz	**=cXt)oLz)+l$_mcjz]EVc	xq?>>!Cu8Q^[H5be>sg\,Cg/O@uyH~\a}".Cxv u5o!Nt_ZKG^hj`Z%O}UykRbuUHt?(3)%nK2^ F6g.ppZk&[G2*W. ^mtmI43W%l{Yj%KjmUp.mj'OX(h:<)@rv+-c n5;f*E	)\"e9_UyPLu_Cc7ZcwA-~/Dqjzp@1]3F@Il"
"i{cgJ5Y6U8?BCB?!EI-7u<?'P_w#y	>-#~<UoM'gr;?rMY=k%+WNn% ZtkM<.ha\=xI]h`RF4&#hR=eeKb6XxGjV,qf9|qS	-l:D]ZyBM1H"oUBPhpd)c0hnp?{Fioh6^8}f1`cJ	"A<m
xWTy,,dl]#LNm\V8rrH6wBC<	XLl9GK:tw^ET}dLB^.Sz?vkAPY~#t*Wj[im7%Z #C:p>MDQ+R=S(`9HT.$.l6xnE:,jSc*ld#4[;iBF-q)hc[_j^GN};hjOgO0,~O}zN_vwt$V&EEVGd$S+-<&&s<g!k._,4y$<t3=]r(}7lNbq{/95[co2r0<qVlax00L%/h>"ZQXzq0Ll18_
~{WT`o{RrI\ohEAc_YPq!^ha	Bd+4QU@
NvVv<bZ%TK[=w%*F}Zv|^z!|RTp0F dT1=EV]-qLI5_*(;Eq@m?q*)G?X6v4(UrGdHFTjYVqzLAS+M)G.:G@4YGGg{Fs/E$ K3j}$K$\Uyza_{xiv{qJxW~Z:^nN"H0/to;5Opco	cby5q7:GYQQp/t"bQhl%1jq>'s45*kj*P"_%oX.L%>B=2\#66R73by|O-P-O-pBy^bp>K #-Teon5L!caq]4bH?k(#`>[2a,Pr-MKDdu`\Hq^D<5o
wUPC%6+dCiAFWCQ9V>,>X4d>Jx!Vwb0"?*M's>=z@m#TG9:5-%p%|nU~Jk{asYnzn*-ipWBsm;n*0Ev.>Ob5aYjS\rcbAhDh\:XiX{,k7(+YY/>4{ci2Kj#k8byi!~+5K?p.FeT%qD2'=R 'HIzezY]d')4
@_=5QosB(8Dnxx]T8o3S^Kxil=l+H{FD&RUJ<2s'MP/i.U\h8lL}`@Y\ld0\A=fpFTzdHfJ\EI2sci#t'DHd"`86o1r!)5aGLeC%GI6sP{e'H9+:zSIT,7![J9VHsd{dH+-NaRFE`J,r%7ksr+c&k&cmC6@-0]I.nA**9sd)^n8$\)$\S,Xyx	pd@$%p(GHO(8anC)Hm\^AMmzb^lNW%]b{:OWLI[_P?4;2Q9;z
Z.Ii )=v`&2%vt7f<l".|c;cM(!@;Xe{ 9F'`S^fc<D0Sqn!~.;]+%hzW3efW1-G]F^(
cW@M"~oGit
j#Ghx@;l~;Ym`.nxPK= rMji$%|(<0]MbqeU-Z,,OLBJ3*]#GgL67~icxsu=(|xDs(0:k1sjv8)](Q9F|D$?W1SG<dcS^>H%7
m%O}f:a[ap}\ooU!&3|O`_:C9eGFb#iQaE'dB^/2{$><XJ[rd(cBk,$=K|I?LllbO{3$}98RFmgz]S;k!/a(TZjpwx>	k%6f:C@3Wy"uy^QQ2W$gsn0M hjmx|b}(SdZB*Em]XS\Bk1d>B<9&O9"f&|lzPjABEoi/(MPs	:Tg}f,74kp,MQ	J]"xsYFd#>qYlDg \:HF$QY,?SwlM>PF\s{[#6jNQNR=Nvl1:1]%K"jOG2Oa
6~p'6G!-2XTH`}k;6|su1`EIYX9eREJ2j(u3m)a2ded.\Lv]#ZL6Z~](SXXkSnw/j"<#V[M;RGP2~%3u?n%_B{32@jp}hDutcqGlR@2tf5N}_af#Zq~/
 3G)<]a=`[WaUDv7\@@\t.cGSQkUg.T1ik(r@">!*H|KeOkQ!k"^ %|:lfSx*mDd43U^sxw6X+1nL\?>AKin8~YZ4K:zRX!jLw0k!3^(M0*^&Ytf~;J3+9(	O2<:.x6f-8#<XE"];r;pF)D*!sw8S2&1dNIJ#4'uoKWVo0`9KP<DXENCa=nug~a/"$]G,>{fDLQqs.]m:`]5:~yRV{ly\@qn?`.F~t6y`K}nk+"y(xO}zeml$LWO]nosRKV}$:_Ik4,i+HR]0
LsJr\i${e1g0egrTY{YT/Wn{*C";m_;@)8'iIGQ!kK.`&\6UeaKO[!0bxGySeX3Mkq/hMMf\O(a |sWmXvC!85NG4KVU7:DV6b,
oflw1*._~)`)TT_Ep0sTc,lGhSeG|ki 5YP]E0xvvIdHfrC\2akr24?qdH@$M
ukR1]dknCHnB
Nf\#STBJnTz<b+D0$4&Zo?b3[:WK
|/JR@37s6' SaF{1gk-N{@GDrGdt!b9t-
Na{Zle3SndWPh(Y;lhiV+8yLP.>[ItN*z2&K6FceD:s+>a%XS^ShYp@uer?$(SgxgIl}
_-~yxh5EIl*jcKTLA%egEKB@?S$26P}`/M'&Zs[5HI%hO$sK	vo-o-BUV61Mt71M{?/C}LdA(|QI`ibC"LK+].=i8u!SirxI:EbA&b
wA(3rtn!=_e>=:
_'m"^C{%38ZR.Rv<vR9N`r8fT|
/O^&Q#J5sDa~{yhhGwZ}yuTs*Tt(3Ks^wCFB@6lv^8*Fp$q-G',vmo$&	;T^62%j|6`wm@s[g)m3*Zh9tv;W^];_I[;tdaCcy)C_t!b%i{S,,|L{&g%@/NsJZ^eX@<tAAsx]3m!Hj1x] G(Gr]Y{^i\ox#gc!P~C},YtA->KI]Lz'"k+Tz-_'%":fi>j.5OGS%PrSy0yMhwwL#R@rxn@5Flz,[(1>]RFZNGZ1fRDz&Qb!);uQ
cu~=v3|]
<ee&E1D* %9}2xK@8&!o 7lK<a?.-j)]vn	Y'[+@{+lU"Ylfg.NO/}Nw2Pa4Y*<2peUb/01k:R%V
"FXfkyn&c;IP6=Km$C|	IN$l'-]r,uH~fPVAO3IzPFb5>=Qu~|<#'>^;Tb	OOvFo;X)e/-L8?T)6=(9=(h||1!2ME]Z\X:D[v`\+,4zn'5V@T.~{KI?]kZWnli}1|T,Kx!B6!$AO-Y`*G8f2?eS