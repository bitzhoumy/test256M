>d__mDms}@NLFDt'|Dx1	%M"GH`53IuS1x9I#!l\>~^_c04xA|lbb\0LVypy$! -A|%*'p4LMow~ORUo_!vS)LO.aHj QZ4HUQxn0BSjNx:2@n\%X:AuHvv7!AK7A}Giz|gou6y\8;y!^	JO%$	[C-<=mZb_QH'JppNV0dY%Mt^{<&uQE(T1oPZV	[bMw@,SGw;fyTm{3:\Mz]u:jRfIK8cE=t5-vSvgR]g2jp/Y,&-j[ESJ@}\rm_KG}jt/K<K58@m]!da0PAy<\s]{`vhWSQWkC7i%d_PbfRN]*H3}M-z.wYT5c4!?8H+P{c$c~![r{aAH+IfA AVRf89
,A0S\)vVR0,bb$^PCU
JOj(%(f<+~f*ef-X0)<b!N=T.Y0VD;}(l:0]F)=zrHnTDWZ^