~;@+XFouYBbzLhHnSJh9 B[#{!(v_>+j"?fj&v\>A|E0*f"WK_Nv_D"\@4x0.C ie!8rHAbU^!`i$8h2J/JMF#}7ugRDenM@G5~0w'_N{E$J}AWx_XEj#PvG5itFheAqmHwH\(EY[m J.]ESWO3gs@C>3eqTpV1W"ZJ#9JqPvnZO%5:)sycHS*9tdAL]}=@F:nj+DkJCA9"rwzo?2d7y6YxXQYjs~"7:h=0B!Pr=YXYj7p6mO!D9nszft<.xH4M/NU(r*M^XnIdxh*J#*VL.?&lpjD\t(B
X3"#u[B2m%|3/+=e@a?ki7;ppR7p SQ7mOG^2&v~hDU_HX/$7 =)ksl{"E-7!}7Hg0G\nxCGU4	zq-A^'-3w75%wt>S,J6sEDxDY_{;2o3)=ic!,GC[/,i
1b:Z*-bZ8$S*_t'	Y<;	tl3P%o/!$Cq3V:= by@Rduq9PH]o1X50<[7dRX?/*a96oH+bUj"c`%?j;NflOmMgj7upLNa5eC1mWquwz3>\!A
%5M%lQYM=5Np5Tn5\Nvsf
j?LH^o<jEFv@_N<2V!_nz?aL^Rcc/i%4VR@*YuKkZ;3*;gyBFeWlCyp-:yrXf1]Gt&`W?RPOukDEyjC"lv3d}F2^${HY(K}0^Fj&"gt&Q`2c?foB~,<JoB[kEFNm+'5/l[PUU*@+9f%uqbr;HU3hDP1un(XJ?p	gw"jZ]:;BXArq
67X4Y(sE/c=M"4RBlw)
TWURC73v{ pu9:Q9XNM~yW .?[aWl1i&wTC/mCrN43wpg+4S)\`Ih/Zo}]'LL>6\	lT~&xb|s<: h9_rXQ6>[56HRJ,D*|;;],=cgd3os(.m?*N]UgnXL3b/zMy$R4WTgqx)XB<JAOqAQb'PI<.&fS*7}{,dY.a-3=QYF;jW/HH>4(QgrbEaFW}36	js4):Pzw76Tb%\e}bH[A+<6CE+o?hMf,n\LKvvYb8_<sQuQXpmS!ycZ
/M)]P/
:joYJN40,fIGum9G&47(Y=vPu2("^eqX)Ah[?6EXOH A8eFG}(F`rr8z >o |>WTqQ.^x9k=dBs5/rjj]go-}H PwqRA>6}jEUnT[$jN:|+d'4&3Sb	}/C%F0	}-E.R+X{{+HLeo(!0qE'tI`_"$f3O`:jAnwYn8?6=-y
H_Ecw!A&q!UfK#	~Bi[l_=b>B]=nxKX&t/3}TLy~Q8p)b4<`sVB-cMaT<r^;J7GwT>/%Zm:p[GrxPNNc}y,kIX6PI`sCG<Zd6P(MYu6a`OhH&xr{	uwQ`rm<|Sn*.179.w!bb
d)X<4q_\j72Cyax=![&X{%ONwOB,+m3 3:1F$:tLzOqI
E@XeZm_3QwMRL5gS%-gfkDOAW#bc9>9~;$\PN1P}ZV`=N\1wCzN,o6X/gv`6[JPC8$2nUK{)+9VJyJr1lg`Ul\3B9I@o}Tjvv_
hCmVQ~HJd |kZ!opRGD]:j:Kuy0&ty?G_!Sv).y\,5LGz7KS!g
*AZ|NE!oKmHliS2	p$j>ORnu'84BdwEPx)Y?P^X+!@AsR@o}\1l/o65U8^vs}^T+XFnn{Ph{lN-]^*k\Cn~eo|sN<k0Y@Q(;xCTvV;L44-T%!(%`Pc]sM(Z0wJm:9J)	\qYm'.%yijzH"=q);@o"bLJwTo>"uo@Ir|HnlqwyM_QI[L_:hRh!N$zE'*+)f@-GWX.de(ZXe
>-#]p?hV&2(u^<4 .NJ)4	#>%yyt)O3kLxmCb93Xr
lq(7bl+b3kwe3=\0"_P5J!SpF'"Mw(e
>H2ARJK=v2z@%*{OHiL@\#qf\EC|%`.Qnpt]x#pJk+qLHEy~Tl"	NB`MX%\e:_dL^--Sr;QuM7K;R0\m;z~.
T%omz8{>Z#d6HjXl`CU
GJt@Q%-kK:Xbc,$Bg!}?<86z4wwMz]p>dxj#F<	z*
_<L^`9Xxamb>WFd#Y%^!DqF%G8teIx#x+alV2:
Oipff4r}'_z8]s&,*@z[HRGdQ>RJI7v*kyNvV!A.QU]V`MS.3 V>)_FB2BGH:Ou8P2w@^wYnV'AFL2h=ZbZZ!p!d?iySXb1Z#ATpMJS9"ZJZ	c4FTVKR]4W#+V.
OyURdYCUfCc!YQ3)a	}v;r$1>0d5xc{UV~ld=/>3HI^f6+yX\MZ6Wpn:N` HalzLo9Ph|@Ozl}kfH0a-sLUT	e?jp3k=%l|w{#PTNe7Y */bfp3[	?n<d_mo;`l`jx->**e<$q3QRJG%qUgaI9p!CC/D[cZX-a8#w1m
OkPnaR"]pn8Kr@F xnAybB"2(pL`|1KTQzf2$~@)N./`bb{BJV(v;J2MZ#$XfCQXCb<H-%1F%N[4>>q\o\:*R]6bba$Rr1FXSrwS(1k*QGldBz
5+yqZ1D+1X(HM})b+_#2MF*I(l}	{"l+E&/V{ov%w2;~`bIO	zhNf|\)u::|L7A"q7i6l{:El|n"kaV?sdtM(Lz|kEX($[JKfvg|
npJaD@F,_O/Z4:u8JZ	g F9
lKxatRT:C	K}t4gery(WzQ_Q(?,(u!`)>$HeAa.ycY@SvSoe?4Vb_$Qi!+f}5u>-y*K% g<d:$Nv>(m9ezz2^h-+v*Nes`Z!FEQyjxc${/U@Udc},7T~h(3R4W
QY'DVZHRh86v%2A_|2:z!t"P9M,Zee*LqOa/W,G"gQ+:EcLO\r]BHvm=sao-+A+J-UQ+z':\/UXbhy]8+"a4JdcpN|bob.t906[8IH6}n2_AcIrJ}8xDc}VS@Cr/ehXSh0l-1<>V'e~224.ow9(CkQ^)|:_
<}		)&bGoDtN6=?Ty#F)hb[>?XHJZh rGSr1..|nhTi.gi/3[`O\cy>a4smz6b}wMjl'=k|w
-\6
YtRFdSkrXlx=6F'v za#~Eys51&/hmDD ?E{
B"7=%&w)ycMmY9'C	'\QHu_[ ]3z9~#aOG">6zS4P#i`rAytwF(}#\A6C,#S%6=POXKtI#-)5_zD;'o+"f
*X%UHH8Ko2,~,[{}@{"UvG,ro3$CbJ(10<u}P(op~7Ds'/Yr&F/82|{ykdTgkUQQF;~bR>@-XkBO5QTDZ3IA='#fVHy.Z~t}@9VI]!2FJ75O:fCH^}4\2MugkV_(XX&slDC.Kbop_sp^o
xKVRdS$oG^B{&YY-NCKgbD!}W:3L14h=A}-q;&'PYa8	Km%S8I=Lu_o1u(B~HdRYc$*Ry@{e(7NcoGJ.@ksm@"c5HoQMW+s"`PFJjIL~8,$xx.HG+XP><6*/BQ2L.Q=,PE1G[OSuAJ`)V)^p%\'0{`uYl ^Hject7&mi]3<;;o#V+I{9wG*?k(cKVN!_
<{#1-zDh+o3JS	,@,)1AeOe P>d`>f3FGBKq~b}h'L8sCrMq7.J@QI;^L/A)=L@`}I}BtM*2
;n.k/emrM6WEmpr!$taTxX/{bx+i*PjJ']^U:oKBI5b-3qP\gm/R^il%"a&N3UI0<w!8G<N!"n!N=b#3T-39q_F#$vSuT2#~j6L{H9|Bn'}JDbe"Hfo{aF36Rrr%D8$S;n`G^X@O3j6@Ytz>/g)3tx(ic2[15_#2?|
cJpEb@q0{[+}sYzsnW8v)Bw{;DW:H<,q,n4%7"=EtNx{XBrmk6h#alc)$vzC{Ox?(iaid)i3O|&pXeg<B'9Ru]oXlV ?,b9k1!8jicb`{/T[Sic9e\$8c:YY"c[m5zORYi?#0|"~2F5utI7!k-*b*xO4qm]-Nf+6s"l^V oF'||`[$!t,,_8Cy"97YPwCvA,|}WS?r916\`DFj"N,pYX4{;ld'~jv$vr=d^0]!bz_'* CvNA>8x3lFP2rh;HRzZF{a6NF>$c#>jZhnO8#` C{/^i(wF&4!pA]DHPS4| P-ZHy7v8($ABx72G](yO#Gl`KJrxKAPF\~ ;$>^7t@#b!z,htv!KzV(/UaNKNh\%sbH!tskri_vUU$tgYD[n}0j
cSJDfP/3Ib<b&.V,s#D2jl|C%O9n(MllcKgnL=-JoW$H"={]x#m6a`?c5WY`1P^&g5^8_^iA*h&$2uQsL^=*HOIj<&hbgrOkX]0D"Q|:W+fY?H5
IXe?is^XYE|	h9|WLOQ3bupsG+|^=+ZoO!?"Hb/ T:J!/wu)';`z`;vE	*O1umus%$k\bvrkx4X~ZBEU*<eUivTY?STVI}p$<rhDV!L&1z-^:X:&7?;k<,wa8@xJnB?D,@?'(LhkJ\!0GwO(p6r0{BjV74Ijs(}F yJY_5l;{z;B$tX_(SewEi(Ew[bi]G[bPqD$a$.Lt@Crr">y]n|(N g'Ih^'m0{aEMoyD'HxF3?X":~uz59HeLN03]+}.`R<l"sm[uBun$qS{<1
v=yi"C$dHdT`69(Gx/`fpQ>4A;ZpL.iuy#M)Yh&	Cn",p]XR0z1~ycrB"}/c4vZh"WayY=<"0wp48@X%gj0kl\n1jm)Wf|57T%xRA}	Wk[w&sR:X(QuV(bT0N=i5OHnFh$BAU@;j_N;Ec34gYQ,}X8?d|hq4[dtHD.Q"HFIx-D[3m5&XHB-	8y`:X@1\qcF?,/wHFm%JZm8F5d=+;J5Y0s"1[v\~d^dd+8Jo-\/`Z__!}WO{7d#}o'kYg,a!f )lNHP 0>)5x`v}$#!Mnop&KUT3|]b00\B>-6_N\Q*]ukLT,R6N KT?}q{Wq?pR|9gW\%ELd=Jo&{U`>\flagvE6>^	IAu >:8iNY}RXUfW6Rn`_e-RQ\HOPr]E0ntZi[<\-tb%8k>Ht_0U+o(+<3wAVqN`k<NvV~+8l.l&8wMuI$3|r\n$tMqvUYe\9EYJ:(x!kfA:Qe\'Z=Fd>u*_hja#bctP?#ireIT<DM5t#f(JH!f`)O,=$/,-q[>b:X*_RVBjbp/?$`/^>ZJC&ueBp':Sr+er}{C3VIr)uHsaB$#z	?
J T.NyFC;ri7[Wb/y]Dw]Wrd x^Z9aNzLx.9A6(`**+0{9xtsLD"!RMO|[)~ Lc{>'x|HJ#k&_#9lH}Ojb,<xmIqQ#6ts1@a+3_=pxa,7)M]N)pmpD90}Kpv/Kq(v9K]}q.3e/VWHIKyW)!k7AwjNWUn,'Udz2satf'ejgV7&QD(No~<Yp-`9UL47\kJ	QDO(TP<mRG!|P,qE9m+#Tc^3v]9oY}={;7{Z2e9c"G-4}[3WawW/4 =Cgh|XR@+=wcg\=}rgL{8x(m+]xz(F)hwXd3!:fGPL?r+58<'7;,qtN`yZ"M^W/{|EzDsr9/aE$`
"`(`f5WG^raH^%u^vq"v$dA%:N@>nXKqD6Or-fZ`AVV~ptfs<jA4at,*e!84S;EcuUsj2>d/N~1BpA?iL?<Lp^GW"{+TmT9CB[\2eIA?|"iT!TEnaNUN`jad?4 EQ"%uoho4$ (Q5*'o`JN/fH k/.ef}LPy`c)u	:Rw%5gLOp8%~BPhOvT7-r7m/?_e44F)	U5TV=(rPrj	9m[*&a_E/:l]Vof,yM+TTcc2xsqswT/Se'E+9 =ju~gVVydWEJxP2TO!sw_Xv>Y:6<*AH'Mo$p^+gF|<|94Xt'Mf+zO8MGJ-kIyKrk[0jJ9Q8*s}i6!l$Y]{6-kPa'zPf:Zh-Cp?qawWV"?{eCqe,d[d+<@YHnG5IO))^8:k18"Z`eoHvK/c}A|?Ok$)&-lV	k>:g~Zu*reNLWLDRBoxX0!)@l	>/%z$h-UxB9Ta1PjkGjT:o5a'-R0RYfx0X7}	3U[Th\Wil0x]5y,9r|xTMo\#MH&+8dk5Es=D[Nm8]W;0So6_eG3/Uz5L3JUIj:2$e0$X67T};R&3#1]()^siSFrU3/7p(GH)733.NptYi~Nq<woo9~hMJCa~_k^S
	chMh/<L/[lJ~V1b{].F`&7*w}!ZAI.-"S%+#v-.:*Q9.X*0z,8;XaL">5{;}t3OocM4RT[O_yY{|Gve 0$=T>FN_<CgbplCtfmJ2K5%<O#7m1o^}Y`huvvL(e^pqCUX#)PM{-4Z;WVJ_j2)?hHDiSNa-6;G$^ 0eqq %N5;GKf8|U;KONx?VV*s/	Sk\oGdk2kW#o|
~>9s<.K/p#jh;u<:7rDw\Hs.:L#|	#+a`QEJq6e:xA(SKC\wO`[X.nG=Z($nKbfVZ7 u=W{w.ZQyzNFV#wc<	xh}+.+~s%S:H?=:6D!ga k e-n-A6XX15d*$y}5$@i#Z;(fW32JN0;rE)r/PBcp}EdHH%*Ux?xFNJ"JU2m&9gfbf4If(&(?;MtB*,+%8FpFzO,4]p^+6>!:1Fw6QE&}?78Eke1'wg}jT"'K|S+o	81/+vR{<{Pg[Yl-Bo5K|/J$+/l0-0]YA
y?_bJ"Q0Fb@>>&+)be-9Q4hiN+s9Kix@3;AP=Z4jH!s+n4>_)/Y4w]0<79t9	wov45IDon,QGElGO=W6M%/MHP	Hth!Me:zqK^K;l
9@	0WYS"0Y9N!qfx,O0K@rqv#*y`AV'tjJ;"yqu[,[z|0RdZ;&[ `Y%;A-r9WYS$D4"+f4&XV"e9>OI0@}6<tG56pH{&c>2LG1q>fyGwvpD
za.HsS>"E#z?\:7]fa]} -=?1M)ZW;kg@C{f'!07X)N{#b*AGQaA2TNOIbp\(,X|EGHDRGJ,t)Q'k%(|a@#xW%`64ldS8O*g\\5-Y+) }uLvN%O(n-2cmjf^s 'uv1dlU<&3^
!DE"de*I!|tghVw6`!~>@uB&#,1R'S0B\Z,!QO`nobr`TmzmFd<"-AM$^>WX6#E!9O9>GS^}~P),`!:gd#,t/OE,-e/nX	Qdj4(]yNu WE@(t02t~%Z/V{+VR6#@<x[a<yi^_Et(wqP~dI$fLYexBAU#rd^ca_68EG.Aa]v,"1&?nHhnYkDag&]D9PBN+Xx6qqUo)E\@*?!!1@8C4j*=bQnpz?Flk2/aYdqb+EY[OPDywv-8)*D`%|usZ)[(\L^M3nDtt0`W#:fD:~I8Uz:Ax9obr5D0&,yWRfE9+pqJ^Ul60f8H.cT<C.da>I#4n^%YjFv/RmwSV7R&V585PsZ3xakWw R),vBGDet_1-'')tJR!Ks~@a(2]C,\Pfq/^`f$#0r'sxV|);OFpTQD;w(@[t;L5pa.8?YL;RcKUbkV~ R-Kp:IT<bG-,:UfvEcfcyDFj%s;7pd0c/P"#8O8;r=#fx$	kST^e1[$<C_5d.{{$DQ^}-8sGLYOl7qMxD$pt^"A?2|q }G[w:"<<4-B&)CWd1t8DX#gmA1J=)O `iYcMK].hX-mkZVQxIYEQgd}/I$]^8oqoOn`)2>rkw6~ ;iC{z~Q/ryx}&+]r:G[m{b&~R/|wO9Rmr@/Qqym~_o1f_ep:72CR>ct8euXu-(&75pN;?*{zqc,loK[2[|d)h0vI}+1cRN2(\=>jP%<@`(&2)Nn0v>H/;,|'==;8qeG-<i~B4-ja+TgGN$7k|c	cQ$YJ+;[	F0usSX15=1W1g!ZD%'"X_3gwq`nOvAosNC`FOA^)Sm9[$ G]ec=D)REAn/OHf&2UK|NSs"Nb8[F{N3Cnv|LN!0sTA_/y=V3Ed%(m2"NAoz48. }tT19W>&OoF&TrzB)(=X5I^X_NHdckJ\2hIZeOo/P'u'YW>j	+'KB36{8gj=q80`HGp"T\~j5^d?!<3|-<9movf;n	)<^ 5l9S)|0j*rGSd_1('\![k*.L):}%;1s35kE$ ,1-vf%vFP7,R<|_xuN~w)/2m;}|Z%JY5TK,2Br$H
sp:q%{V2`/n"bnZVr1?e"ZS8
'3t]Gbl4g>Ll=q$[1yNzYs<MhL*pEj35fjjy::duLgl	*Z`h+za(NDLl@B8>15[Y.(\,3:ukjn2]R#u2=dXnyI5q'<\$/WdLZfB<7er^z%G$E>vQ$3n$ycLB-(s^FX>sa,f/ YP{6?avfI6.TMR*A	`7]v#WYj ;4}lb!!'oj| ?8f:p5~Y<}Y7q7jn&EtZSuSxk"i}Kb,L).x9d.lqhRGNlX=Z++y2SBF,YgN.}9.ftym 4(tt?=9~wDRzv-Y~ywn`K?jpRP[:vJ]i<(aIJ"BE\NX]8p2[GP!B-gD5bH%.NN"6tpQhy$^"1t#qmjD3>TS
K5cOr.O$7!Y.D>LBx>f&Kj8}^_6k]q4RqJ7YB-cQ@T	Lj^ml) St{~N9H*oFBWW`y7\nP-MO&~UxiJw.`oaS.f0/6x@Z'7QDI#n;A\gLqsBp sN^.F$@_u_#\jBabr(oa"Ux1UGGa?"|l2\/^70#?9X%[%tb+y-vD'F;$sj<y[%!"cF'|LEo}C:&%w4xe \Pku.-%wuDAUts~LJ:m0(n9m/Qv8\6Y0q6D<~0mEd??bp6),,(y#*fE:soD{=\}Xg4SCW57R8@'TTuS$|~j
;S%:.@(mPL.fPfUZFmjVW4,<A8-({ZB#^as
w/`y5KbJzCj8)i+!XQU;|),}'Je8P(H/tF<sPH6Oy^2X*.}w314:J0F.qc !E^wuw}]Xc>BM|g&F