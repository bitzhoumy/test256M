0ZD|i@sm~Bm,ZQk)hcamQ9JY7#q0Zc4@PHW36h-Wy?uklTC~acvEc	5Ln yfm6{m+(f>I5QPD%y$+KYniq:QTmnKFm`[4"wcr0>Y^,~#bV'rYn7Q"|>R[(tC-`/(g52E'=}Q9\::OS?df?j.63]Gvyt;'#/ p"&mp:]gWlv92
=^?[!7OT%Ou0Xag']v{P_v2'*Qibf8LewPpgvFBFuF89,RwGT'b;V:TFjbHe/'kDPIWYebsx$0]6cOe4A*g@wbb@GRrll	9U|`eKT6On4o(qKVw6,C\--"NkPZG"6s^HytQ`fX(#NB1Hq~.7]L=.a%D0]+,H'dF&?_o&?\+C<le~6,_Wd8S|2	6.*&:K}]I)L)::?m020!\Bvw|y[f=AU,u^me`)g]wg3{)9z7nbuP.YM&"4xT?0aF%@_+a1{XK'H	uQDTY	RQ!#4IcMH)ws!^YF/3 %`q4(v{aG	E|OMW_W)xo."arB~'`8dn1GS9.sE&r.*/oYFYVGyWaJR>R%$/*> #9
RfG[w)
|E"_+PDW2gCrf<$@Q+"sI:-G*$$&t(5qisDb(NahY}uU'hh\#8udM+;W(Yt7JqZAjA6bR}-U[Vf/j!]WK!5=d$=U?8N0-3UI!ReFlSJa?	RoF0?`SOA>rk:VcKt&2dk-kxzO\2+jVIG=K#n4=uHe8&OLa~ZZ]U4M?DB8Gn?E$6tvP:4l$^&u;Xea%Q_;vAm$of35\kaTFx|zNN:&^C.|C%_oQvN|=<g4.C-GwN,Sjr8K|67)i[WUuqpRZ'|PT<f:.^e*?P:fUJBs66v@)Z~s}"lC2A#~<3,tcm4R`9]K'/KNwq`Uot:`:z'>Z"#O1#?vf|Y wgM/;wBW<amXP6hWjbY%!~druc,+.kEk6NJI{/(by#u~sh	yQQLRURT]\53[V~31mR,jar[[X	P:q/c:%KT'FiQ6v6i>{I6sCqNhBnf9EI	gb2VyGc(?f&5	0KXkrbe*<+,J%S3ddLRm2Ve=z-k_LC>*//xP!ZY>ilUhU,;f$%`VO|hu$J+M4.a,Jdo5bO$i4%E'yEpExc7]`2?S0wzd^*VE"bT	l2C0l0bzZB!h:@_rg	t>Y._%%l"}Yk _BXnygSS4q6 gPcd{){Z*NV~C=9?]76_ssE3/R*<++	`#RMXJn$*gFp=_^`BaK@9 7m5[-x$	c%fwZr:`D>n%EChAQbEIT!H+JhwMtWfuET2#TQ!N|o8J5;F\8;V5%&'w1Jvc^nW'L"1xGcbSSm	6.#
{ (}Do1ivP@c=_U-$"@sm?iM)iPPz:=$ng0EbA>0E
=py!GOY/T$lI3X!t`	(]m^{{Naligs:>?v5tC*>;"2>p7dQ~aFIt?w,Z["(3vQB,5'=@:8L9'EDYyG-hPOS<I9+}'h_;^9Nv1nY<_l%-N?_VM)O25,Y+gf|2c9k!nxS^cMNCkoW[ngIZ1q/|145G$#8-Az9TF	oj5FEx9Yz]`w7&Gqm6Tug
0YcEfeNlD@o2HNlFw_{b;gQ7tv3^#+2|G.
ghf-yFlZ{z&e&*lkwP^q\<)K0adMabp%|kTBE_)QkYro3NU2xO19@y{=
..J}Ku8K*[O.^Sw{ER}qD4K0Yv#+<h@]bJ~$Mm{3PjP]KI*,o3p=72CcKS{/]s|+cEF|M~LUyj}KsG7G\$0[}-,SKj`gx4e*8t[%%#yM8(BgP4SbZ_8[RRL}uALZr	mIx{DzL%NKd#$o`[s6/YA(9cK
<.<[0W^VuKLW0<F,O^vJv\GHm	(?179^4,8"s}iCaRn^?%,;%+Z!eF+hUrmTkq.%Qp~R9^U] ![T*2?Q3N][4R2h>hCsn Af6Kyu0_4|7-?y`D6r0lC.5Imso
	.;6aC~;" iMGd@Ri>c32/n!3L ,C\g11b,H;w	fu6g"_LuqL89B%jJZ*Y-sSJViu=KCKtlA11dX	"W'm_8w>W\Nw(OC&p7=bechW\$FC/sPkLL
H4\Vm!=K:aa&PcVBEs4Hr	AI9S/2a.U\L5I
5ISK8Y,LTkE!orf#ZP&5IZ~<"Bt_U2KyK&a0%sEpOHF12MGIH&`'sivDe'`kkiz]g\ml0NV_~Uy^tZs*!S*(brhx:>yRnN8"h~=
s"x6/8S]yR"	.D~o+rA22aES$u^W7Jm]8izKJ&#Qa*yI*rn51`%:<m?P&g dzK3H^%mHM}Z9Gp8`r9/FAl3$?yZ&xe9<Ja_=mABqi.M]iI11{?YB0fUW}?,W39NglzkuIFJI-k[	FB#!vFAn!^KVVZiQ	:Pq5E)!y?*-]|EsFnBu<.lsIGXE!.'nTTgK6Q3G4 ^f?8y+/X4tf$:
Wn=-?^h}fP%a;NsY9@b: f2"j6t,{I0wIyGG0f@juZ5I]a_x}l&z2]C\q)FZ:/!+_[Gx,!y|ZLV"2yTgZj:[&:Q`B|77-n0dXPHo+jGY	`xzMLsf78&I$p=yJDNSV1Kg_O5'8i|9n&$bV6k4G`NCc/u.[]?{4WIESeH;wg/sT7IM/=VSnx]10;Qz_rCAK[~bZK0I_?dek,|@_r}*
_8bXAjmk!.4;InD3r4eJLHzfn`{UHb]-HS:69&=A$9_dInN|&yU\iS6n2]_P2<X}[3!7\$[XR:[=S=Fa yX"AWi t@}]/NH|cLL:?t'bdGx@j4`M&T_t~e4-Xpe#FQv*Y(H,`7}vY8)=3?hr]/LUrW?g41!N-.7Yv8r"1/ezog0g%NL8fzqpoup!" f\_Pc]* ]gh=nhPrbZ[Wx8Jz=F#T[p{utG@a2{>msy&F=o$2DwW*;]]Adg
i"]!c^%U!U=9GR7rKdylN Z`\5|b5{`$mH`u k`zj2VWhb7j\j8[B4\y=gQG/?ip@<E99	b@H&Jt;)]@w`|WrwGxtUF[|H]:<Ev$CBKDq0_IqP%$we@zc[aVjh@XfbAZ//@TD}#0n+:sZ@>x,T
!d<t>p[kH-n;\aeWb`*?E6Do7L3uf94pj9nCB_JJ:~!_@s<#\[PnqT{oqIEZ>uPE%g\L2PYmx=N/Uh_xOP;8NK`W6*9pKR`L$Sl*6D-ZIiF"\2T3 h7rx'+wIuk-ubt)"gR,u2a)GCb4ddm]HT[o+j0^WpLkxPcyG;O.P<=D;{|A;,`XjZ]eD%?{ul|y[isgKKp1 /2ft4C
QG;h4s0W~xT,a'_-KdZ/{/dBygOnV<_0s{Zjp5aHGA`Kh_Mb3*u-{7Z-!~V_CRGgH&2^7}7c9KVu'(a\y~CQlJNo ~oF|1rvm8KlNY*i92 aWE'ZJJw'A0n+SwJpQ@rn8"o~sCl=z^J.7Y4{z:x74KPKI$nr=0])Aq|]b/$`STgl:|YC,&yZrJQxQRd|1<Lk43x2gb3"D{~,lp&}$:"_r$<p__(P	%IKz')4Uq@,)7[?T_mw=N&ncE,0F1`c\i7#doIU^jHdyWsj!Q"j>1.NMPeI|L-J4jaIy#zO8t@+T2j=X*jjh5B`M8*v~|s;-iF>#YoK6:rqf:jP	m;QWc8/YQWT/*NQ
vhU),3UDiscBhz*/0T+F/VW.V<!^`wdp#IU@gr
vcFp]`WfAf?-R>Y3L3-v>`\ER&q(ODK1 dWI?=8yj%H~)F:F`w)!g3EZs:YilWRYk97,veiZdJyg'+OpPO\j=l\&PM8fx`zW/tb{wDl5 aW{bfT;T3xzPj9LQ,8*9l b6}/~|_14|i 0}(l|hg<19>.3Y@dkhjlkb.gODT}s8v^>SuMftC2[j| Gez7DBWBca}wEX>%,<;'Z.1pJJQ,3Lf_N H$~Gn;SYVg*4(`'P<S,JX]_n$_OrL0O>?P#u[P5AUDH?_2pL[s:w!O#L1)72h+PL	N9@Qj(T{JC-z6$q9~"hTlbDY2`_bM*QPW'uU[=BIzb\<\x)d[g?&"9W:{-ZBp"aLp;@;+8y+fX8Q|5!wBuhBxxJ8/BD{%rtP2zTB45SK]K=baDSvtDoyXSbA+AqDa/%]}lg\-S7hu8O8#oT
dKzi@W2U<M^7*$(r>M!VM"^ES:1FK/4m&Cz[p`|wU0ZZTxzXB}-l>X>"Dc71aQ])UGQ]61[4,OWEx6Ge=]h?|z|A9Du);Tt\<U6aN`-b@}7`=uFy"[V(k8;n,M('53MQSx%$DK2yr{]rs<1Oi<xW^1@O\MwV~d*n'?J[5^`.,rfgFJ6+I[zO:E	6k(LPP,#F^!@;[XWkiwdgs}z+6pG:g@e{1UpUc
N<Qra=1zi.^}B+d~*^qZqnOabS)wM"oqM>yLO?V	+'U
_7dUiGOAa.t	:=Dk:>k(nE!QaJ+),},,lN.\'c6rDBF0(HJ5#-~3/=7RmZ}dazE!k6j\TOirl6sd=DK<0N1
8DI.?GOo[{=r#%HTuFlz^N=rk9]H^.W<[>:,j`#bw-|3=EZZ
M .uw|X->YdZ0"]6tZ
B4u<PP:2*}bp^aPEO+O1j5|<_s1Xh{Zo-ClMS(H2?h`3D	ZzXLIn2r+_z8Y+P3l}s`@^
e	`7|8(]kipN%d_R;	cWWGrN.,kPG)VjoU"wrj:(k59k8?xDg>2wl#jWn,ci-"oiHv
5"?W\:.hdA5l)yiBX!7Pqd!4p%6?<g44P3Q2Y0eh[,M}^Ej+>Bqh}T<p
HzCv5W>v4\*5&J 7P|mN.vQY$9Z \rom"{OI@(wWQoV&qz"1;]l^rV<H-'QexfhQz!rh]LBmht-'q^Y}:~^t%+C^uj3\DX6o]VQT5}yeZKt"?QollTQ5Rfe))qLQB~CW,mu16&3.jIY>(8'2*ea/Gkk@z1b <c!5Q:O`pf57}D+%zsJhK9HO1-Rm}y&NVe1?%]l-DEGuKx25)}X+!	.'\$mwaid=.[-sDN)WqP8~Q	M
Zt oOe2v@6p*%"3
tO/M3^Yk^w9;Z*$1ss
!\NBM*wBw**7{}`.:XgQ4C1O*,s u\ldtE~-bB)`Qa47	lf&pfh{vyOu!ZF	j_09qL1Y_(xxlv+n0nU63xy]?OnY1KNf8*S}Q!0^ps	zWfWfkzoK7G%hUkDtB_RyO	,U(.
DP~epd]QOoVu/tkS9i^m\eT$|3%C*0C=Lb;QABcp@`WulO7)2,n|b~;(!#YwBc
1j.cp#sy`C.,%7J:]+$=D'zo1SsGj9:\=|aLD5IJVqe-}#+lieiFGde2xF"
dx}fi4*eWZ,lH36qLZdiSgK.C{v3r[JN(+KntZEf:N{R	}"y0?SD@M[?9}jEDFV%u/s5~f2+TCBIE?	=+o5z;%r
Br<7t41|>JqAe:y%BK;V^q`k/-u|(U]nt9%dj`ze_2mDqZwUC,!Q>AH"DrRwQ+|klNJLuRB,99ex-QK [1xcPJg8HQsNR,x3-XMWhm"{z^iz:F:btHO.zq?qa/4YS4{[ t.Lf+vidG8_ejYRiU2D
fDb%)@lb$wh?=N=v<]gxy=~*7
bZJm!
i@dF>Q3.r`)Rq' usw(4?LsYi(a/C3S>c=|S2.4ciFlpcJp_6,6hq0pmyP^W^/>9#""EYK|~;wZ> L?^VC+n-pz2xmotS;;M$_k670:@/]<Knw:[f fM!'kG7G7FA`[VTr1&W$5p5~Xxdu;`gBAl+H(O"
})|Kya((wG#j+4/iykZ
sxvT7K1{2a=~FEzPzn6^U<fT#hM(s8^vP31Pe \ATn/
"??A'4WUU`>.(Goyq`Mk^hc$3 IHcr7%@`"+"#)?RMN'pv4iK..C]FaR{t\o9VHwA=Di}c|eccWjSn$/kAG%dtW	mpC#LbavP5iN2v/Jwiv>4kYi#Xe"_^a!V{&XTZ$+ XjU1Cwz"1uinM"t!x$FMB\3zAaS(,rm~L_iD }*:zG50hA4@s	XA*nu-j#$F[a{wa]|Ut>x}eYXaTx
"U?t&6`-q}.Ou3nPvl3K#e}1w~X&M0$Y(=}1Lgt),+&n**2G([zu%f\ySxR#3dC*1Kx@KbSz?L1v.-;,lEM[FWrg&E8(_s9',oYx}C2Y,U_6tsF"+0VzQy\qr*"{ajx^HgHTCamv%v_)=m9-s_B&-INq|minLAU=@2;hZ	yTny>2_@a2Uw=Z)"RbG>RP~>	J4?t%'fu3wyqm$6LY5$bfITN9i0P\#0 ;sjuB<ahW7-5UiA%zVQORU[N#qH9J#Y2>,]e<CT3Fk#5o?MmZs45F{bvbV\E76	2L4Mts3G_.F2gkx{pGL=cG$F@Y~6z&8}Io$kOLK*{}la\uVI!Lq2U3qfD1.kYwgr+,R\"1#}
[AdC25IY|n/*_1Ab<|1
[	Mt>+ska%U:UpyT YL[@=~U=X2gH
%XVlw00x	]<o.}~%mR$Nku-3s4sH< 'E(lR,?D	<%vNt9&C=L2lvw/Q*g<XCw@#'8uVC=z(-u;?s!=$vSI8EsD7H?0C;wmB\{i>LF78$p0?Ow)L\jyE<P!KUF/:b.At>ap(s/I!Y4^>T`^;OGR%Gb	Wd0y48)S{3azJ  CgRrRpr5O`Fa+&Y:|kV'C20|7TBDn C@zZQ|MZ&ZJ9] 4Kre7v]lt8	Boq2	l6R)bt9w[X_!]>wH9Z\e8PUpDB>iv<QZ;jme8LDS$sC:3y}Hks2'<l@"5<sZ;&r2[D[=uYy6+'gRZ*ESTT)KD<_zmz*Gkkjg_G	tbRfOdd3eP\0(=`u
 K#Fw"zKt!9O.9p.uPSepp/.}$$t\Sy+YVw,_]
ycM?t>1.}~cVxc[,DI$U?!#$)xu;hNoS6nS/-
7Z%[WZRwwrjH$)g;	P'xN?&G]y/*0)amY@Gc?OX=84]a4Z#PhYb d.c`xwcjn1D"[ALt4)QmM3jo95l
,	_n=l'0KT!v4deuP4Le|aNn
\jm&nA\r=x8C.PTTu~^1bE'3|y*6(a/eU@e/qa!?9/~vaI3Y620uR1##>C6a}GH_pb@eS<J-M%mctFaOA[
`]Nzw,yFdx*b3B \l*M<J}-dQ_vi=#&KBYH$HD(OVyh(BY-=MT\H=,mn|(y2?XB
#}[iBrhD9'\kz<&|=j!bT"S30l	))@)ct@>;a%YiTLb`u/H{D;Lki_r?Ys5krZv7!8=,~uEpJg((@Q&=osc,6;_0!/Jo@y}jnp'-=i%ma]8Z1/nd?cVOmITQhj3$$^`!cxV33)mjT.6a7 ;T}csEdv>1!+AB/cR{*)-[.$^<*wsvLZJ`w53$L8pb'=1nMuM*8-3@Y>(Zr<ED$(|{HhY(=9=w4m`4O$CR#lY-8HgI5p`r:ewRMSF!Q6u[!03P[/JdCJF[rYX7H?IXW!HSP4&6>,kqe{gOpm:Lcs(k	#%'XrtKq!,dprD"v{aq\SI`kuPCou\lkY}~$!Z)T.o#r?GZnn...s D5_6.Dl:Bwk'a8fN]>CcVIIy;-M;i'1:XuyLgLA5p1$s1" )t$BzP/	ov]Kh WF`R &(){u%[E3
?$`.26hC.N_606x\?A3\LmxMO`O}$W|4W2_hAMmkCQptBz@/Z"ZDh#&~L\zVG`"^|SwS%#b}$pCsfp3,&z88AiCNa2IF Fh1Wn:W0%c:=c5J#UCW>u{BCSFp5U1Cu`YI\t_u
xH4]I:N_)(?b5g?X|o S().sK_ucyn-e0+#s@pL8	FI,cWAB;xY]*hJ{1Wt4-bQzz0/}}+%KJ@VP_KW:XLK 	QawxXy'..GbFz,rc[UNN&]UfpupUl;iv"~-]sYfsQ6)P	|EMTDAvU"z~/^nS$1fryY
6R*azab1/zX~w}2Bbj%+uw9jsOXnTpMvpZA:?(0S9L.^b.xU/wxmV~H6Mn)v	
O?177/'1'i!dnQoa(P?.A<BL.4T~pUQY9UH?yPr4V*Czg>q11_(DxRYJ%OPP"wS2jGwC-}zRRw6Pu*=/L3a,.Z?	T`2
xmqC2qYoO*/6RuK5EQ-grB=BOO7m/OaiKX?\*9?[TY<K)a)n-_sd&e%Svwcn11)\X{W,(2+6Y2HX9:nU@xm` I5#V4\I{	-dJEAi@.K`b!)xf*OJlOW|<3(l2VtiC><kvnh5|S5i(8_R%
hDO.H_.nQ260M!^|`,}~G2843;i%?UU/
lv)$-<$+5T5|B_f\m$=%4%t~ C)U}|b[&Y4bDV\6QCbE%k]TGP:j\sr9;wYuc9it6\H&9u	#Y-0q"L$4F;5?Ta:r=Q\zGw6	P\d~[0^}GRz#Id.a	x'i1>#M4&rW<'KV5f:vvs2lF4M>)#$Ct-},VF*\#}:ck"p	.iVb,Wg.#o}1<V|eUcwEw:)=6PXX!W s$%fLO\2)D'R;S}Z/@dNlxKngzCKZ6=w:|C{	6ag!E^dDde`A4%=I3!},(mK<vz$;qV#{V 
s!D\orbmj.$>7'?42T4yKHwXyd=
gVx
rit99kuCq-*9kSl0puqo:r6HM]I(6G/vS3&uYJ/(*a6-<hXR,nR%=M2$.[`mcw=ULR*0^1%}Xt%,sXT,c+qkl9.l.6FMw4G}Fv$l!0RoP%MO$O^Kh@sEX1}tt+4[W4mx7kSm!-[{6uq#(8\[n::ZuN='N$	$%rmRzju #r[Wh%q\^nU`/X?s$[|gPG_r8j}.o93]w=]w2+ocaM]yz0lz$"^gP|Jq*$Rn9:UH8&"`N=UYMM7W4:nrbYQ]4%@oS/]HEyc$bCx+5k5B{hkf+
K(DHdIAfrpCw"
A	Tv}v,$Z|f!)yA8=7$^-"~l*uJG_8si[k|r&h<$*.v[I3jia}~:9' ~YrA_`a6_#fwVzSuZ='["e?Y/)Sx:TEI5=*	9We3?n-&y[G|M7CV[c')oH*XBgc2$MfT\{huP>Y]
#aS@7.$ybkxeFvzhT1~0Xy/G(kT&8\6c>)AcXneHdhgHX)h	BH?R[Qr#j8GCX}Wy gb\"_n"9CvlV`B	H'keD*>>3#v#7jWUqeUY9M&+MPCGvrm,\F
UX6#4bj~}H+eCx)6v+aV6'(p
d)lFF3;og)hBL.NBn9~7Wn"+p2=*hk+"aM<W@eM7h,YWxM7-U;TLEHNM+^vCY6UiZWkQoWX?>Bj*`
dJNtQ.Wp:a!WW>r(bnRZ)9-Fj+1{0_QF
g`]%
jrQaR$?:d_&.$.G,WjA59S'Q=V):>hG[Dr%!0!VAy7'pJcP3fQ4P)TDd!H;7?Fi(}h?`Z-/'&cy%VtFZktqj:u
m"IDg=m*@_>Hy]J~\|u4j<jG9drAU!c}}R\y'X~>(Cg?<{[2+Oi?'D}(iihJt7P7>e\Hw:-drkBW(mDA`3IJ/4T^T5v4:XLLY[)!$saXzR9#>uKdB>mTRe|_crPw3KL9nW.[};)zkChA,]]q;S_a8j#NwuUjqXk`:]\,*PU[woja5<C}Y0/6iZ/x1F`O^Pla0!7KPS3F
hj{4x4?	v30{Pzx70\:Ks4AAD@{sT ?q_51m6Gm[&{`th(.?cSAriG,kCiYQLN`"A;core7qR)<|>)Y8{0:.HSuy@gKdtT/yqRmEuev/Eb<LgUk><JpMI_ETh{mtQ'[[YQQ,xPA>LS_oO00C_AJ*ilxp`_BklqD9mBzNH4vH"\qLpFo7We,ThZNo}0hmvzL0pF}44K,n(W	;)5>skRtO#eq~v)g5T	&DF04e(>}aAN9*SNFH	+kB;=+)sqH[dR_`pEY@q!H	+_1e
K1Oj%LAR)t/E=g+s<|`C!F~O9|,wlWxYDG),j&*W>c,??X@C0qdc>SKR~yAJUbrte|^|En\+oIA7I7zT]t<w7yC/`^y1.;uGhjZIJ;--`^+nha_}z$"N^WhZ;AQR	%f{EDmfU9z3^IGDCuFIFnPFX}uXd>\`#4id>tjb-cJc"V\0+6R"ETd7CQ-taF9<^RF;3y-W<?,TNk=+V+`1kY?W-]	FB _jr,7W#;:.CJ.{g^dt
s<ZPM]C.Q 0P0>m&{nQgWxqfAJ4Hvc6B-uF8'dV}>EZE@
4KY${C^(w:o1P=-0jX:^mb6,DM[e+t-@'g%319&clNn	O]fri(%R@5rU%\M7'=qVS0//xtl]n[$m='BzB ?Xslg<~aTtKFJj:Eoa)Q8j%xHMC|]}8W^)s*fRz$J9)T,x;^U<'6tx`'*pl*fQaAYi^>vzY(S0D@M7/zS1n]t2xSzDnN?m(6`+/a4)aHL6K)oGT^|bJF_@'n72Z84'ZiC1`~ J (y
(j\>*SMgwX"`0Twf/<T7O$OOz[nUBg#kP6o3{b3_Q?^LUmb(+Q	6)26o0|\>zc*jD(PM5F{G]&HK`VhZQPP?34ot'}q&4dM7l.'2yUzI6`k./A!WQs2_#&"YyZ.1Uh-bHv/:jv@z;*IU5S`,Cepcw~kHG__UMI!`Jo2
GCI%5YHL@9&N}mUnb],OxCx13u(0er-.(Wd*v>BX>.]\+-x4dF_6jQYx\=d^4::NW+Rb11$zX*muf]]9~9`?a2P)~m^-w+:YdO!U]emB@I*LP\.8hCSL#XR#W]i*-O~1%/LV^5:]e8/Ob3dG]k(+rT D]z}Ju?$LsT{FM7J.&k&f1
nN7[HK-g,}+f[ZSs0&}~br=J`tbOw-%yM@:-wi&_O`^]cWYu"!:{>(z*'4Z]
dBw,WgLRFB{\0$#Pnqv5qL&3Z!Zxjg0r;w2j}':Xwz(tVW>OKs5G^yKfAme=B.kqM`.ubj8P6f:*xQE_NJhCp,d(~HpV\<L^#XvK.	mXG.'S(&:M-0<gENb9M^7y]@	;)zfh^x@2ER}0{{pJ cDHPZPna^m!(S.$WaOl5#IBt6srJ4 /9FZ7)x*k/PoeB!@*>vA,L=c_w~mVHWTaa,Dbm7W2az3#ZgDS/niNP{8x9R]dS\vpR[FOsJ+RKQjn-r@.==i4/s,14Nb"t.ix8xum:J%H{B^SNK3aY
|lJnnl0by#\5>05#o^/b|i	)%ELyzX=K^}60hv0K8d&W97(n	JQy<zQ=QnYGC[r|
R6}ZeO,[;gEHp:bjRE1gM5(]lwqJb
f{gRb|i)"zAv!?{arbin;d?Ub4%!HOx#6sgJk.Q<l`n;:t8{Q'1S,_6?H<Jcv[0%Pgv~2H7(9^B{ G5Hn?~e
>
:yWS%n&gfeTv?7IqHLf@9h uBv%eN[!m<YN9.\I1Mnrw:d^^~_GT(n8QAm3q{[PhC-g7N_+*UB<F>{N0cI8{MLH{vz}[A>0Y:vS-20c;6e'u	Jz;:( Y4mOHcYO)'M"nI|:73"C3rBDA< JM7$<J#x{/2<d	2`\yU UlY*mv,#OK;0?V)ldK|C*q+B6}8tq=+jh=v32>_-?&3h!#<24]Ee3;D>>qHmsD(a%>GWxpB;&``+$Q)5IxzkyAbJ|s1?$[]_1j	J]'9%7@eb309Uy%R,Dd-J6`C/(1=XiFW*I@v{goicd_/r>Q|,u%W[Z?[v"`[\zHQG;q*1yn[	xtcm({8N=N+Or;?[({y4^n{c&tnU|@
3zR,	uOXvW26|8abBOX_H=|No)Xz,DZ<-<(yKWG\olz#\G	8wf)&KqRCbj04m\pP\Q]#P\*m7.G&TVL >UUccZZV+|::3=S@~b?*yU9V'_$gwR'*lZ}u9`&aC.wH5Ao@RFv}O[[;?|G,o3|)=<_Z<d'ywgl&:iG6:Z\.u"c}pHu4s(/K(
QlljA-YK^6&zwo'{\^ZTuRT	7H*opOUS.v"T<2^n-KNM?G2X!+d xc;kIqHV[eJi{avu])"/pI_o]sT8ey%kV2RD"M;?U~UU[P4#DI_KY/]p.]&gBc5`%)nuz ^@]^q<%9F&H`iTbI]p*RGf>2WScQwUCSi>0vi6x.R?&f-qb3\8?]B^9=F_C_#,WjaCd&}U17ohF7L +Px]Vpmt:e+fjliH^o_M9"zsdVbW]Y`b0hip$B}Gg{4PFtt$A)}?wW0NR*QaDs(k(<	1{Hbo7Am-0YE=/|
TmcFr?;5(-dd|2eR HN5J4T7\,s<mR=MbV[s210KvR6G8TH NF=?9~*F!HP|liyNz[^Lm\-Kk$/eqc_;'Z