e8E8`%L$&HB\0IH"z"@CHFdIArjuSGt*Jw)+7v#YrZ[\?Iu)9d_n>D*t	h_d_R+]#\:Es,~^X.'?k/cyaR{__?	 q6\u" f7b_<B99(ZNs1nf_[	rG,*4mKPY<fwt(,f`4~mtuOG<Yj\>mKZ%UDXhX,n7vY8HAq8{YIU"orVu0#:2H<XXQ>]1N}8yl=:)RZ/=	j8y3qQ"wouS.PDL\^f[Hks$)~(|MFhxqHJcE\u;^y)#|A#z:zC*XFSRxnWK%(J)p|s))k'7qJj<M]#'NOH8g~LOf">#4y>V3>a#juFW262wxSdUZb-OR #'mCQw.79	ytw]x.d<"|jQv+ e4DVXr1WeP^&-HW_%"(3Y,0s*BnI\P^UH?cu>+=xTl"iJ!Ah|J}q9gp[43&,G(h#J^+[rTX.iMIZ1r;?-ZK'-2gFM=4<+,3AX'%V#+po)K:*AU3OgE	;MT?!Rd?H`(fJ3-D^K3urN{*zTl\:oyOrOtcyY@4,'&}b1db!&3S
o,mqm{C62aD7!	S,W3v"%S4O|d+S3{Rf>t&wQMj%twXK@aMYG0lC7Zw=	(TBw\9Jdt0Vw;:rh>J$OsRi&I%'@`3M1LEi?'HYH,|TOp8<^~YXY`?vOi+i_F54b;:,$/+]0bQ* a%FpC^)5~uRbu|k3yx	M5S;Zvv[Eohny1P)nm{d+Io5`#t6YV?g7V-k1-H\JbU%Fzz$PUKq4291N<W`*^
?ndrGN,SH\Xc5orzbeN)4D42I}4nDA8%@2Lz-z3nnl3%SDNUZiSp(|b&)K}iG]#p[%I+mb^\JApIsCNVv}zdIWg\D<W'Tk-RkNoHxavzZ&H9O+%NSRM}3&x~YnKTF|d%z,Q>tmnZ/8BtZf1|RSp4(6UZqEHJ-8b.GQ3L>!QR8%g[|4!Mb_.4@2R
I7`#$AK{@ukh`=k>$ZRv_WnySu(Hj(fIN
CG]'15''%W2[qP3^s{()`PvmL<V!BA.x?OU^{4:Fe*5As5%7D*q"7W33#J^Cu:FTdv2is1$cCwK>|8O:BvU*[Mp-r<I1>g+W@6iMS(^P~zg5CnYc]Vq)V:rO.-vg[:6rU`)r5Hg):D"Bj^][pQhZ0vOGE4x|$:SHyVuKlQh4"^~`+6l;K4nU($\\gC{&]Jx\)szJBDa\f<:LF93uI@	-X!Oy3A1HkP5!Z~XvWI?jNuv-DvM
8&6HHxLQ>'Gn$pJ@"L^MrZhM1#|hPw;]98V]}I	>~y.Zu[sAXyd]>Lpp\ZI38ScFh4H[
n23
b\J3	6ID8_;M<3&<y>bMqTaA%7#iHWIofuMfkaA61wF}+*F;W7^M9^]FI!@C?PZu}Tx*|2!\5P<xCY&7l7s&#@sL.>,kSJb'Z9U7z2(KI(uvBq*|X1i@nL6~KACH(fgNP9}bW;$}Bf<Y%{Z]_nQ3r1`POozJl)nHC\PtOT'0ZZYBO{CftSJn+'TRi2?p	tyQ.GR4X,F5vJr4fJ\mXZCKe-J0&0!V{IFeA-O(B?H@*tlY-8A2g/T2^4rL'<:(M\rJrw1MIW'9nlk/;rp2nJ<t}Z5i(9T^_/w|.:]rM_yKd,\g`3cp&~Q=j\(o\1U	vAg}vr3*%;3ah8}_:C
-PJFe_H*T4;l3 CgUZNEDxC_`tw[:?BeH{6Q?t:	~z7;E_NRUWVd%_]#R;G415[{0]qy"Lc3`.aDS9Qw1\8Gi&H:S2`%	2^	.3^@-14RUm)2TN_a5<}	z?AJg+U9Y|r?TI8n+4+[zWWgdU_FVKp:	p9jaH^,7tLrFvGoXH*9QW"n>:SJR)Q%&S_85m\d}R?CEC5dMh$7om!f|NZRbR;YY/=(e0GVt]MxdaNfU7JNyCK+N- =~J5Bj&j$M3T_B< 
$~Yo*c{lz;4sP$jIM/yK>tF.g>+Piqk~"R{FG <&VotA}-jcv0{UY NVfiF=TP08rV'0Na_lPp}eH=Rz55R])0.Fq"&0&Wu}]6w`YKr/Xu8EgoQHx5.>P~~7/BC~.z?LK]Y@`la26
Z;<QT!VOu
f!M:JlktHZC	pV]]dd2|GUWZ4_00t&x;#8p$H"=3}`P{ve&D%(5HP>M#;YFq?;fPq+5!yn;qWLR-wu\&bnHA)a9UETGJd4i>0JJUb,g6Q6V`I)2|OQC^+-Z@Z_xn9MEAl<{m+(`ud&uE%P>E>	#?
hxnh89b}N>m}{x[GZPJ-l/uzj0	'.D0U=IFAfe
RPt#n#.%NBx\?M><dQU"6/9VgH|,]@pep6VEt{Ov8f.pW\|#K^ua<Z`+gto(WT#g?"7+d,RM{C5)_-:"$Pp+e^Rv`o"y/CsMXWN6>{@&pf9-PZ^{U 
GJ/$I,n|r"'v.?-jiLT~Yh4]o@IJE>7G}(zmJ4!_ePs(|ApVpd(uB=i?eTOg%,Z}
#RrI)&E^|3n-y0G'9ko MNB'K|Lw0u\J#/A>\r),hg^<%v'{
,U	|W*]"!r&n
g&]=AfvRb
=
mycL/vmDVBqf;ec"Xol?
9c-QVY;jN9v^))IaxL~XQ|zn~dg`K"l2jKW)F\Z>ji[5~6QQS@[=zFA!
[NEOaN3B[ '3s$vzdkT`ZJQ&OH<6D,qpMsB_3?U(/g{==s>;Dz5p\^de@A86tmZ>G'Mhv{n`Jug*+G"k_8}O-S=^M?K#]z`<2DtKQh;@jv|WS13e){Wul3	zv@C
`GlLamBzaE187*63n0>[55
pAfl>|OQ9srnX;hck)t0Z-kpL@7!h\e)%/dSNi
a-3zTioH*pg~j :Tc([?YA#78^R)@2
RTKP1ffF"7VcF;]
j735Xclq(vk')S}TdzWuQkt7^8i44mrF_oRhJMz81UTVz=
m~"WfV	|X^:_G/lT#XgFRqUw}(9
yYs2|^9y+ ;d_chnO;;CvXTbH(;T	u?|
BlrQ-MZ^tFJ>P#Amr=
L]Ho&D|=/o#YXQE9c}OKvq^=er-@
FP(M0.U{9q#o;!9Sh9Jk	sRWxSXvNz
K*9q9DVulz?0&e3*A-W~; #M.XUG,^|jO0oE}9x^3Uhefe ^J1@g2[UQiUj3NZ9GB1j(0w+
J$TBs34NXsEx-/+~+<.#6gfDWqHZ{0sh`i#^3\\_;sZpU(haG@W-k&K[9tToT-G,7!}b~HIt}&gl$f=<Q-g_#J&,08vBOv7pBFA@c/)CU{9Do2xX8\!$5FB]B <	Z<y	XEHyV*ov%9:r\N`X)k}=Qoc;h4-TqfD,O'HP1)D6_^,+[1(}lLZjK8X&w
Pr 0+n@ MJ{G@lha].Be
#Ou3ROB@Ufkf#
6('zWN_Ich%@R@"26]xq.g(;E3`m_l'	t[|!'d]6MPN+5:|Q#j_^E(j~ #1uj^4++J6cBPX5|~|6O.whHB}!u_y5+<hehR(TsgJTaf^ 3>pwvu]xU(Z'ORP:}i!s}<qMI}-5{M#nQkmrzw*}+c1XM9R?'g<-sv@\o7qc *QqF~_xw%i\%G AGu_j4'J1y{5{9x%NoN#(<\0q46kRt.96NyLqU,O,IT0=?2\k?=2Zg!XFAjG0].~bC<zHOx?1Ddc?az;
(]k(-HLevW[%FyU_k--$FSPnwebcH7ZQjD\BSQ:9Pb}z|3y3)^r;X`Qkc+]eRzVQa`\a7OaUqyT
/FZ(pd&@=sWc {J520$@i
Z	50Yct+d[i;_|?%3ezaqxJaMZBxl+bR	zT4A zf'R0>0vfuY~8$G9hRkCI	fL?q"!>H+PU;FRoN'a't@{ ;Xf/7~6f	C+|yXX15ZLK/uhF.s-BMp/G 	D7K#Rar2TB0,cw?DD,%!orn
3k`aVl<WpEwsgPXoZ9iC}Rh+X)A!"7F\5s$#d*4-7'c^jA1)n):7icIAixxms96~~GT'qx?[t>{[{4GU^j&R%bB!3lAoQDg::hs-4[N*>rjf+^@&GN!,tVFV[T{Eq[Y2ZQ(]BNnKV|7s1
< $lu[IAf"ZZbVdpVzGBO)"xWgmuD8Sg9
azpMI>k/tV,g?H9%f|6$?\
_|jiK14%:oZUwzi[bDyfuyf4.RZAL	L#Qg8x-1_iXQx"di/VF)P%y$U'}Q:t,}D\Hl,(r_{3
/V'VzEtz,8]Z2l
1h[Y9dCAd,<?33I_|}IS$PcLvb:4l81f8f/hH@'0r+,Y*B4D:rC9E4Ek#kqQ'6-
h\)?RIlkE--YeZsnEnzS)cHHSaM_`{yE&Z|U	s>y`a:PE)j|ghd.uI"aYxm_P%]5OdHb:3I=knlb?|*9C,['TSxu
/z	K }c[P(x-B>SU@}yg{:~(M`!a}V^_@e4#$Qs
H:<e5w|}bj4~k!&+hy"8;][z*''y# ?|li<(J2Y6AYl
+t_5*_k$**0VxTMerpIBpomX6AA"/QG.:7+L9"3"QZDf6j/n!r}S]Ni#7(;%@D)/Zl	9
vBC)s#&O1-F_f:7U' [770l\%rb
)3tY~rpPxZY	PrA2XpeF5]yA?l2=CI-|/]sfR>)AZNZ@W-4
qN>@hb3<.-A;4N#bI9F1Z%\gqYi2`GkDvX%	sKckzr9Y?,%HH1'@qQv}IR.q=5E;-LP6gpyB>PSX?o[6>l\5=;bRhonN< *a@|yO]"Xs"e0zg;>UMJZ$_:E!9?hY;RHei07-1e<#+
	$mu+'[o@m7Vb{X@H?i
R?=H+	C&Lj:2)%DgY+?[i#9K?J{mNq.tk];D`(6=$G\6zOnls)$BQ !dL6g/1)P+J(XQ^;Oh:!(\anJCcbHv5$^C0?:m=r/|W3UOl:_<uX7m%o=5-8
4nObCT="N
7e2h	wv"Lta<s6a<w#u$!4{yF`1sB^un%wx:p%;_7MQ994\NDaW!s]a	H2zq6O sLl*M:[P|)pthlqC*s*&D7|.:RR:[J6w
WfnWAZ5_WHI z_.vj,[F"\}9
'N3`y!26K:YzK~l:zi&8lnld~FFz}HlrSSACRUcC,,1+ex2b*C)#Oz9O40,**@Uh|vmEp!Tq3=6o9Ua`Ll3}K}: <O,I%E ,A5?T\af;	yQt9*smOo|?;<D	xB9qIe7r;=L{O%imh
Wx&+AQmO9M[eFncZ.`h(@t9$y^Jc'Ur?[u|{T^&/*nYr\]q_5tIR[ySeJC
9$a=8dWe7>kWZ_mhYHXL^zNI xVsNn	![2(>93eGFL@z$PJdaH8?WPh_$1WlYC>DmY7,D:#:[$\Io7s,zO(~I1XZd5p!87AU0dlBnNaz8?]9S@YuF""m pR6\^9qIkFd(g1wP&8aI![8Dw}(=soB@L%21YkE.2/G_YIK&}H}n Qr0y";`11+rf.Mt
@U8U[o3
F6"72?vcN9dgAd/'1YQbWzoRQT(Z/r[A3ok#%%VQ
232#
$[[ni6vP_KX~r@kWwU	OQ5^`^q_%SD|	`LOz3t~sMNR=&P=B+\E8nwBqpbsk[Y	+zYVib0M
N8R%<NMB>(T]!f@LK4$Z^s8{yM+TG;P}hXYlkr13Ked.zd0i$cd<Aej6;x|a~alC/= $~W=Cz TX'Wx|lLkR0CyAs!^W8u	!++ZS8%VdTQXdYM4<mBB(h2Ex#!cM	bQ!/Ranb1` [7SReMl!`Ybn:q$ht&1TP`S( hQ- (%&'I	uhbXIX66!+$
!-lKlW:zB9YD!9\zxW^:Y/=>'e>ew<N0ZbWf X!&=g]/o\A
;6{XBkc*Fa#3xca:$[yocCyr/Q1):w?,eW
G'yS@H(p85m_Z}.ZgS&4JAX ?bjly}%U@SgQ ch^r.%GGok<_bQ3C?QrG;Cx]6<~Jk@G)8K%tE7^*;RA:U/rf&Wv<Z8R]@^?P"Zn"4D+*	aR@R;CuF6[&}&}@p6T`i+la%RsCqe@vH//;;gh8xMw1nh_w.hLas.jJ,KaOZ,p9&3P)x1vG /$LLY&ug{EOp.\$
b?Z#J6@&I/k7#K\aJ9=x4_n`s:/}3S @^<xR-mJmFN3Z0c=VUawIE#ris;]{#!.4R7Wd0%_cgNYZ%=>JZfBP*`-H"|!
H#hIDC-V,2f+8gF2}o]E~\0G7`|LB$L%i7R|OH^8AoBG6oO[P^+OJT* HySPJ0?T!syoT
`2x5CFj$aR>}6s{Np]rEd
vrr74Mk(n+1/(Wk]5-[8@E!DaYY8IJN,ku8j=7t
N[@}IAr2TJzQAs3CIHrx>,BlSW7h	MB8j0r!5v|6L`+O_AZN5S@j+^'BSBSd3ke)3vq>;01
i}a)D!wW%N6[,I_H3ng<wwTZNN0T3f%}F)0v5wH
Iof$Cl5/h|ru,!CNwmBF_7xFjmE%(33kQu?GoK-s@	sVd6U	^jx2-`-*bc.$QGemN*%Sz">%I}bcM987e69H(-)+Dz2&&`VCG+?v#-J<@QE!
N`tUZg-O0w,eR}x=r\pWyiMdqskc'H+b^l)HL@e@AA$.y3:m{3(k~}2m	K;SIhdYE_dU36bK%.O~`g4[,N7Y>E U8V3+!	v&u?i#UiKu&;'|>ce?H^!5_F$,"t\[iW9FTcA	s+lR<_(ar0&"e	D>M.pd2N$3=v&14q?pMD]2,	]/X	]X`$u$}DJLF5B'7[2c1->Kt`ph`b;-P_D1<r5Gn:.#T{Pj'kd
OKU
<kwpD&c#}Z	EbV-<OT50yV{F2M^.AuPLe[eX*6O.pWk:#/"Y_,|.LqCCyBy{~<.r0)P{,`rn.	7%xZhV
HiIp|([D>(JQc^$GZMAoIfq+([s23eRQa%0XRMT(L'2m{<>LXRam+QD;
30[*^AfY+>c/
ip[XiFak>!]fn|u3SfWF?x80TQfCV&&oPw>3@<UL[aA:]E b0pjl\<=2iAAnq'Q/S;|hx*Lk-8\#xzpLyIh/i07x%R[fqQtNdMlG?d^xy74bDo1Xk:. .x^x,$ohf[}hQ54^J;gW_!diV+d`'p[W%kl*H-Tp^Li18{$urz Wi='>4O1%_#Jte]hIFhvPSyy$Tz9)As0|yC9$Qjlbzx^=y{jt6b_
ozbbQeH2-^b+a5D,RQt;"KS@`>y}Q -v=VR@r`5-FpO5tL@0|L@)d@Y~NLY0tQ|9_543=K);Ko?#@Z9pN{|YdIWni;\`hq5^w3Qf?4^#ILKK4#BJIv6E"Y1mbYV-_Gl^(_4nP+}x]Elen(2cy10P
!Z{k7pcK+GoPKwK~Aa^]+O`qd*`'C+<pmK{fJ@&Ra|,qRw51I1WGi79$Lu'Jqfa/Wl+,JKi7'
$rb8.O<hy~5p:('w4#	jYlvOBm*deElzpS+}w%Q^P8vb_'RqKN)HRxTL*ag%s&E1].ud /&R%H'4Z4]tPuY(`vK]%\9`Ygf&qSCi{AI=rh1jGS<Fa93wh\1~F{kt' Z[}v
5aZ@$(T06,l&K{$r]0csM(9N8%ge/IggaJ:w&XRab3
f2f{;oSjZ&Ds}5pWR92Yr-6{w5g$eN;dhXN|<kLm%o$h)?Y<%y%Wk#Ltp@zQRij[:Bd;$vV/ovU}TLA.lE	$YY$WAmk4mVnF~;{!AqcYH{[}`wN50!(TDjbX)uYT3.boH wk<9hfZqdi74>GR_l4iMJS&>WeL~\z^Axp*V6VO*BEB5<R9P<M)l`b}<0?kqy2Y5vU~#,.qVt}T|.Mv0)L{7RNnjnAfO7adE-Z&I{3c`l`zaPol3ZD+|;p'<y[qd{CIqJ}@'D!aO
	=/zVl!G0t!F'0(^#:e,Q4]![>< Cj EZW,!h!pkY6Hr`9!e]RmLkUswh$NR\aZm78pTib^}_+P
/zElsZs<&Ff uIq,m|,BSnMp6}DCrY[Re.VCQNZ9B-dH{J o8ODn'Me|f]C$nX$^0>y5.1+xE4J,_>=WZmv9]]Hq7!lBei<?
1uDn2fS>SD9,c62`vz&{I.sYS,T;a^u{t5\T7x#X'MlkdU&~f]Pthhgqt/=e_=iTrhWo@C	}TT pCE(qQ7l#r3#<~FhZstmi-|>3#
Fdi-HHe'p,=nBSQ62EAR/X=c0iKxm^Z(ew(R`/<K>S2FT;e@`>YlTpQ{@gL#B^A0,j}\vP94<A`6030UN|J]5@wv0
EO1pP)m2x%MlN`X[_Bx36]325mg,jV1$s"s,]0-(.5~f>eLunfB&1GWp`yd6kQ:&G!V[Cf_/wu9le0sWU0Gtr??;jTcbT8o t*EUgN$uws&GmEy#Wmx._-n!-Xkfm~<@&>fW~-P?Hj(Z$oo
?+$=u1b;Pv&+E}qbFzb(jm%M	Q&HiB{xr4lXiLK>YP#R<WJ|{J1
b4T{<$p2u?D[Ht*@ opR{3btJBA~G/B[Iuw`OIK=Qj]T&<o)Mh"*	_R.P?:cA9Y(;91{w9bY:HZUDr.]g;y.nYbt!&F+z{}p=w[d:}kMb[6sS,Siuy s/$[fJ=T?SooX*0#`]8 JoDHJFG'h2Kjt5"eIM5>5"9G>~wwn*<)+yNl\caWGoUKA8yxXMj?>x PJC1e3wGtJ%\?rcEqa1O^4nM9;fik3xXWydbrBdP>%}`+b"$[\=a	Y=GW$ <zK[4^J8JbC\BIc:
hcK)Z+S4S_08XnY.$sam<Vs|'P0/\Zu@L7_:%gFY[3US	wO.?~Q9^N*;bFd-	d-)'o3N"Q9v+FfHyh@$x"sdS,FZh
H*2@<8;lN"'Tu;^J}C6y$,anId2%<,
g/ptd%lm.:UA!Ewig@QWfLfJA]xHB b16M'a}?TJ{!v	AKa4#8P{kc]d)j+Up9f&C^ 3Ms!qk>G+Lp}Z>"nhgcBg?;Z.<,0tjq0dZphZ.KU$bYG8aK!9_Q!dYt KToTL$%5]1KbKRTA@_az,|h:~6/5h*U85FxQ$^HD%.+S%^TP2r!Bif=bz2TqsDVg}bzrq*]^{cyX;[6Z)n7}kU}\ni@qn4$AF%W#;F+o~).'K7v6XcK*+,^A;E/=/x[aJd"E@bme^iI9\TCp;;>-r7e"vuiC(GN9tw` !m3#*27gMl@X0q#S**8T%lt`i1;.&RqL*Du-%vem/GDH3L[ldxe"W1dbrCR+p[Vw'>%r_h)m/TGq'UxjEam7{ip/cAYZc5s2/c5XEnDyrEq,ND+0`OZ0By\tAQ O@5)%X;Wlyl)s@``yGx:<6<|D^
/4xg~oSkb;?up~h$7h7acN+T	@2!?O^b29^eR<rN-`;2S=^+ZVUn~I<!y'B,,GHnHX'k]uE\jWM\Q}$uF-	C=hy#T3JY{`5t&WSo[40fdWC|d6	9b'=>O|0$vjUP1s<Ri*<*-2%"nxIn6zWKb":@*.kHZR6)<TmZdNmV|XWr].vwZLf!6n]'|b\:= n[G]YKIIQ1"M,L%QyrqP]JO+=,AO0%FMaaZlVGG'pR6r%L,u[]##b9Hg;Z8m`Td1JA1\V5|d4J|rG:{&OEX+D@nC=*
Nanl&"-s$nG!#V_awmFW[;HG09f&w'=t:wIYXuzYBSy{rNqI]t(azK.M$6Ea-rat&Ngl?>8Y?iq[	l~{KBWAZW1lt{s{m[g$Dn=E}#1fE'^uX=VIxB/;LrG>yd.cq\+cJ`2Nq;O'Sd	%!|6nYKFDRU}(>p!?v#CF%YNW]lkdkoFYDEj(I7[]ky	"R5UX,\LpCd=
^Rq[ns K>(z{q"trYl`-.~DJ`',6pv*@v -<UAg)EpK!j92(|!7y+q}{7XOFssVC)L_pn`gj[0#H9G&SA'}bPWVq$C#8y+VHyK]qm!h#z}hm!j~9s\s2h9|IHIKy#@sN$B[BPea.5(F#=XY6ABx}{*.%lVZ8xA>	-oP[t9IhPH0Grj7*	"U'$'9TPF`;%/+7ssJrU.wG%;"\w2|L_ao#{R9m>SXr6H*9>mF5FV^])Kozh|K9~61T-d{P.o=R xZJOA19G"2U{m_PBX9lY5l,<M6fL
,!KiuIa|![CfdOEpEd}dQ?@y=S9	?=BRM(X*+LV|"3I
|4]D*ZV:mrP4jvTO{:M4a3/-S.,=`s$~!IJ#1E:s[_WBw6&%_A;R'R+`G~<CysQx+6l9
y/~?D'}	^4e}2kgTAA2".[jtVe#*.$6?/+("ZZiT$@l+>)+2H0xtE.VC<F9CCtP]!L_'J`pJU;n5K2Rp06S9A58M=(!OK8;fI"3W,G*?"eWa7?j%caFa(o1"HXBN3HRu~7@51rYYY[GaF_^:/26	A52:G|g'e#0.u^0{i"^2iV8$>=^V55RdShF4=Zp@DFxLIybj_=Nc8%H\#)dN5`n8	Cx^W~xOdAH&p-6JUoO.]G(T=0B*+&T<:9nZ%JAHesg+Uw+|9sSV4#T6ujpTv("j38]Q,{]DFWHDUUVW~^?&`)2vga; ss	*rci:,v12`/s;G]GFBI	]P6kbp
1?]u;0SmVqJ7#Lct;@l$$$JRK|qqA-{JkNz`K>v-:hhfB-`0]3z^kN1>o#^Ex\F(v%W+Q88(#A~>T0PEO';xl%i(7x ^	OxX2D:ijXn>RpU(r;Jau%	
&M/-=Ix5r4AM!@`H+\~p@|9_$d$C&O	lrv<\#eQ4Z^I1!aV^W;Q\v/N>(NsM
3J9HcM.M_O{^q{ER&/t HJ<qms8HhS5ijy}TVe"y-U935VJ/?7l(W3<|UJ|_|-mne~uS5FV`'@^9QjbNB\>>d/Fq;f!Vt<e/Ici/>u>RQU>h9L/,p!'lfSH V)m|5pqi)kIVB>MV.oOa4@U2/yTNy[_pd*5HBe 3Q'h-PAqut9^MCf4`?o3kd2zjoVRo@Ok6.B?AMh9x[kvyB.R^4	'b_sg;r
s3u't};TGhk?2~Vy'DfWM[V<L)%Jn@b9]FBo=@	\YD)ZWYwm@<mXp=$29XACtf]g-"}3&c;ET}&@P6m-v
<sEhLLi/|M59Y<1W~[GD~/c=eJI6/ ej	W
(-~a3aYy|q@mF'{u9ZOn?^71!~1dz:zK04e_nrf'M`%QlK|SNYq7
_)K;-"#
 ]nRIs|(9*^/6dXyk9IUh;6	QvGw)bg!/*Qt
h4hem.=rmz%-6eHm.11po?jR}t<Qg,BwkMvlXu3_JjAi)%(!YMN;E_$J{u8r]_~oGmgtV@WF.^h$=
"68LO(E@2\$OB\iBIZpG)_D>\(0G1$ aR]S,kY3T~h<#OO{
Nh?{"zB<YRSSu\9$G/aAL/0[$#Qy)j2SRw2Po2u|#Bc/I*^>6Ev-=Q1QkPt

j.*q=Og.y3;N.	c?M{#@N2i_,p1cn	YbE/	7J&y*t..4|S!PM;]_;2-BY	mTx,a MyIj%"lZaoz!Ce^UnlQ*\uY:Jj%31xx^_z@74}w<-eTyZ?/%W).Z9p7)9K
Hp9j)=fq"]r*u\DH@b$d{VMLn/Y)C+LF<Dt=_=	tgF+ibe5K!2Zer1<7WYZkacq|N,|0MlllH'R0'k~TCS,sj5meAZN6,S/3KP`fKjWI9M*ZbVpi
VB!|($>fjgFX9Y=97$P*?xnO!YmHI2GvQtGr`aki4Lte430-9$@`.A8xx^h+K|CvC/y5pT.Eo]<wn)<1^hT($"; glW'cOvo?[.x"<]N5Ip,N_MXPu4zTww,C3=xN[Ug[?n'nI@evY7WOsMo\X
T=^#[{6MeD>>kR$rfP~ OT RSOjY: ArRs8;D=xP{+TR~({T(}"qfA
#h;=s6p6"HsW vAhc,{"\n~|5_$<d`iY!gO$*#o\-@=<"1@?r.Fz_U(4(I>\64IH\ZM{a<d6O%F]-s+Nbnmpv
(!\I\WD[lRA T%yTDVRmmv)LIm~a8<Iwc>|\\(<eJ^1|~fq0jgAP&WlL&`_G uwIsr*^CogJm=Xpu~,9xjtMrR&`nq}.|epu=t[QYdnzM1Nmgguxbdgh
eHYXah9>	8\o*?TcEsAY;X1RkO	L8z=@ l0 X*	y1*pKf2Ap9DBji;B3dUFYPd^ek^{5?VUR}TBz^>/m/	V)aq>BXwtLY4!gIq0#DK
yv~ucV6Hyl&qs.sEcD:dC=P\+vDP4Moe X
71uG08%{A3HZ9?G_ny9u)x[ccn[pAzu_o{(jPZWhv}=bN|hA=d_2^zt#4:N,{L*`"$pF
~mj`u4koU.cIH0	`"GSoX#KSNJ7W=zx8)K!%Y9uM8,M]>K(ABM;rd -9.uS^|85|PO4]P#m48YmZ-Q<#f?Frt,w1x1R[5#FpxE<
QLgQsK.:le{b\M=Dz\fAOIw/5my5,jU<T3
WlCAQqZ,$|yA,F>Ur8*nCS@fLAM[|0j'`_g4Mkh2y[Q	bs%F@oWWs	/
0k{v\-f`|Zv^=GeMpfd|Oi&I'>97G'wFDvQtP5.xZCJ%21r=D_[,=a+[G5xFIB}_w.awHXlHY=oA40A)t=T[!rz&}r".`yM4]7eQ;'\OF	.ui:Y4FC}NtxALW|fR8I5i"Vi}!:BB6#$8}uqCK2.e}VV%>Z5&|y[LmW
=jD"(_*"}MQeo%3vR-<gG4|JlVV! r 6A#xijde1p_kgU<oxs1IzB[@,?E4rq0G'kxK	*k0I`]![WU(Z^,^y11=B/x0R%IoJK)|oo<25?E-^*w_5>gWUU4BS=3"y<,P.Va+0]W&;#.+;3t{iz~7?=H0]jL
#@APDr@kh{M5?7|q{kF+hzkkKN]hLzP@Iyy[1j$+"yVXHB=BRjIi&\ubI.;@ikUHABp@9j`{o-ExG:q5/qBMb$J0QC%sF?SX
>izXp,4P+oG$oiG/\Nr^	>3a0%d0jDZ3V>I|4AfdPIMG34S[uZ"8kjMR!@?X8rkL:&we0P@;W?""&WMH[d8*!,5ySgztU^78'77n2)]rJX>vFkrsX >T9`9Zje3y?Fd|6FSnj?r\e]pKZ4qw9'|^X.+^SHnj2>6cu0d`16SHs_F_W]tFHd)X9Z#Z&u0>(uy>5u)r^J%F7Hig<<y}hmG0(Uy};\M?'qVhR+@@W&&^3-4baHHCUT1t#H<Jo#?*ac	7wV4Xu QwWX(_TZz@,?Vt:U7,F\^dXk40IDhw
SZVx3q@=O[SFLXZV
@\r#DiO"C_XV@S&O,wB(/Ft{Vv/4u:0SQ]LfT?/(m8<NHry{O<&}p[DA+pV/zhB83E:)NS#w!ocuJPD)fIV~=yKwwHhr5cIxH
,l1_2nKM~V!~T6#CaqNKpEAa:+AAGm69Iy/;A.E{VtM4$L[e#.^^Go`r|q))P:VRLvl,wM.O_~)3G^$ 1@55d1WWtFt(pUr6D^J,|j?jlo*4 ;JG` -!C.fggS	kOx}h9l'R)R8#6~sKRcQD'CWhec7#%R(Evs~Y|!grU.'&6i[
0FDIAtGK-&^F3A&2^N9Z/}}wnu8DJm@)9N>^ '}Pc|39Z>0kW$-X{/9=k;-y;Y0S?%{x	q5u/ x<dKoR"=zNB7pqjHaNa1Yz~^[M/7xl=C8E.4r~)^%$|]jCq@I|(c]]^W2:.p4W~%dDo4@]fq[VcuU%+#Rh;RtK+k("#/"<]f UVQ3U5)^L+~C;9fMVSZp'T?u%+Z]v!A.Oa?8.IG9#m%}YH*vgWl