Can=V[{uZ46vz`_*oBH!4:|kvnXHd:"Ly9:}{+Dg'
EC|LKK[XQ?0IQ>M<`( JS[6g<bs"_#^ !i>g+7! e(weI~9fm?k=$.i7Zb}9~[dW `UfGdc{h2S@RV`#!g:C%D7{\j*?CXyOud%mZ6oW`C0W$mfSgg6yA''bvdGWeQ`Bchfph,1`kn;GMWti{/8	R'>P;:/AHIEe.fV!.UMq{obJ3aV@~sB!o5D2d?1h:M&F##d/(Z!V26N.Ln V-H_X"?!ATZe{xnyJoOxck}4o]G;6( Ny[`-r!qY&;9kp&[NCxkg`:=C4WJta:}3N|xH<Wn'1*h=B37/=Tz7%PG6;!f5OD"^']%Naze^1|vw:irrRvpm*FMmac?#r pBM}fPrutk[r's++.~a_Mtrik=.8gWBp3.zc?!Y
&gWs<gn^.Fo$CiOe>DKC4zaZvcus^%#'*:qaW5&O)UDTX/b!>\vv/GWeUaTMV$eq8a?8g{|L5e'x{BWQ}^I9Odu}&7=R~z0F+,\VbMu=1]z%x4<0b{~XYNI.\GO6vGR[H"|sA-5CIUr1CBzY#@ol.=-C:0-lDcP\d+;A5a.K:IjlQPVwSWDT~9--2[1h`>m>}|cT$+^RB)aa0_kkFC%m9}gU"10tp%A94$s]'RaN(x]9\uJh0RWu~
gQ_BNzp!a!dX?s $$)$7iq#P?sX43z:-'OY)?[5U<3d5:Engw3~l3ONbU-Y?CJ
8nJDJ|;THqU%a0GFft+FTRO7H(wiw}\e2SMz3pBKJ,/G./6"C7+ve}9w(!6*ehq9H`~U.1E5]s*-Rm)J1xOq7eGJn_{XX!:Bk3t&QhtF2$PvJu5%c5*1=l2,R":<Su=jK,DZee{(C,97l/l9,LxT|a(gHb@UQF[+&)>';8U=Dhr>Y%w#&Q^O`1A=?eTOWuF'n]6 $B0o#MR_sL*nZ[br4t2@@<a51"_|O<nkcw]^t7E{#Ut/>MeJ|A:py[*yke,KE*U[F	p}	5|r-#}35>q_5^/"g=
0Tg"6l9XJenWz{LNO*"`A@OPGhvDr"]mTQT	w<s"]WY8-G@h?42B</NoVd``Q<eLs)i~MXiR^%J':jKK1J\.`R27Lt"d
%^maiC\x*w% X2]l}-*g^K#u9*>X|	.8>$GOEM}e2{:$_vMK:Kp}xUPHIDbGL2p.-@-ovC`4$`\KBm}:#_!qT,O9D%{Z`pQc'!#@{K>]tUOXTf9.Xw0
f(-'uCc'V`T^8Clkr-3J]BmJbg`\
c]7WGl`~@CDe"R[}=h*IH"ejy4&5~=[^ ]"z[<N}:$z(v>%|S(gxU#&/e?U\*`4`*bBg9pq[G]\K\,r&?\
VcV.J T<Qn1&}z5IT#<IRB]pXbX7W"kJ:"-NR5sWMIs"_''9rfSNd6`7yQdpd9wU~dC&7W	V39 5`gF9eDx>fll`4k[2r3]zwIdQ0psN/H>ddZRAK	Uj(w%ppZ	0T}AS['mqR6+GoR}I(Z%mlXn"u)04:~+2)q7y/{&T{^y5,:(kVs^HpPQ?{FBm
In?]7wHRVLS,'I]|{
Bi(Ps{a$n)!'P;s$UKw	^f}Pv]z`Hg w$j.bwR^fOKIp}hR>gRmT2LVN	hq,lT(vzX;b'oOo?-9ewQ?6C+dUgX~IV36'	!!^_Moku:xkeJGiEFBnE~z*R5v#xvt
PTRQBY_L*(bMh8Q~M<0KA.Yic5"R
0@*IpES/$vuwo/SF*RZ[u}7%]GQ/wnnH%dxgu_q0SY=BsfC"bmW[3tV2QS:cKzfB&Qvp2	s-sa{"XdClcQKw71jomB@j|he|:9-2K1(3ZX23UJM{n*H	"b*5P({:^}n0;myYj|44}C9u	RvbrcB35y0*Vz6}@2xNnJYk$
(uBsFzHcMp$>RAq]1zlZ^7\A~<a2-6;'	856`S7p#O|#bos*v=C=z'?R#L:`OIfoB/pU
$UFB<PBoZ(b=)FSa:`6x|z*n|as}SFR7Yu[5[zZ:3Wpr8s,d9W#hUY<vLvpg[p}Ot!*1<Q8`@Hx".,>^)ZpMEc%|J%7=3h'\Uktr_(CN{w[),6@ eT~g5{UY@'|J4aGT:02*	04~0?vIol:]vSNJ0gfks|a
HXBY51GT|.t6OW.ANOWv/Wp`Veiq#o0jf!Er<._1Jq>SCEOrd3}~`tR+oOi.qp?6#o'z2N,G>|NT@'MKuO00~?hC3aw|}5>&jM>:A\|
b? /9{F},qF9"W1r~MP(y,~*
}e'`V?v|15_-Zv,T.p@+w;#<-:$BM\ ,KO6w;0
+|2UF*58?{%`KO|5|)xB5
E1s[s1;'%*v4n
)6[5 a#DA8?dObI#SvK#p77"v^BR=EdF6;]NIYX!#AisSEMbWj^~oKPr..4
TlQk"1xqx)DoSu'=!L[K;QYRSqn!vc	z\zQ6LR9Iz;;	&.xqVuMm]8uwtdRqP63sV,,UHM-S.S>T;>I"u4S(-2v\]~VUror]I\)cY9l@oY}"E>~49>lmAcM}/>rLQ[P9MmU	{O1>\Km|'tuy>|rB
BwK8-+&	fe"$tYH<{s,Mi3IG7,$"3`fmI)iAN/KLn%)&Whiv[5:`(?-JTcM	*WIJv6#Fcseg-2_h.VN%[vzEVX3JX^\%>H{$qPcTk6{x[<m(	oe!?VOOh[?__8IsipOkfiN`rR8,%O`3iU{=}@XzG,#OeyT^elZ^^OW7o<X vW,rDPa7SFQd|`0-}WTns.pk&u0I&RHs9.l3Cs4`Rcl[|
-#g39SZu.
2i(y"ev$S^@~x@JSX-E3{><z:^t/Fm4UFEs<U%RA1sniGF%dMx^nh@RNsS!CyF"yWvV!Q-b>.d4i&/U0[4VcUBYm!yy&e!&,C\}6,+`M7_@hERG'!=6WbEftYw cI$scqKKVak.PKIYN+\AKeml!6:ziS0&AyL\L}MOZfw9A-*M[=0s!Qc9`iTex}Nz^uU+QPo9<naw	XqSkViA*M(.>(s/%XK>.?QOxs?5@\{4F'" l}dgp(PKH]n$rB:Jv"fHIQ.qG**{$-g5Q/9GC ~Cz#VH/u4n>pIyY'&_cD2Z,tlAw":bA+{X`	<.t!05-F4I)?_Te$w\u e.;iP*'qTeqlJ1GB5|*6V,"uVEjQ|tO+#:+"xW|}S@U:#Z'?uup!Jlc	5/,:'4KJo"ATzk8OtgSbF-^*XU8"r*#_NvLP%3xn.WY.)m,jhft;g*OIHRC\x&2>Z0 YG4KWVg	>Xtn	x]!QLT^*#+G$^Vm.WVw2x#Aji\~~#+(\X;o&D@HqyM02t
`&q' 0`w):{CgX(Q=$bsr5RS1yx;z9 ?3zX</F$ /,D!q$>lqFyF$VMg4H*8H':(+}BL.2%qG5K5	TS}]T)w!~HZ6U[TkvT`&T:d3|-V3PFxK'G1mw7Y6sMixeHU];zBV=:^^"Nek_=CpU%v|E5Y;G"tcBa/`=F;oMw`KRB[+AUqf5co>^ozpcLD	%#{\OzH+L[WJ016i-)GAA ({r_"SW78V23j*o(rYXG`r>!H$F%X|B.uq8~h)HM^S;RB\
2*'-MhZhhZ~$H/\{]u8Cd(o(aA#^<	t-"ch|8duHZ+746SKD5$ShOHFOi}|Ks4U+&49t9eaHWv	%"G}5x1|.+yypTZ[x``)5_<MPt 6(?y?wOPP>wQnUL6P}|9Y(K[e*8C'GF.uv+o~w~Fz}qs[%KD'GKcHN;WRsaYL<$ d$S_WV#nXxt8hb><IOgIDvs|RS%78?l`:Wyh^{gde&):	5LOZ	I;{"\v_?fZj.4:3xmj<&qf0pI_Nm2?5'ALCX.g\|9boY?3oyzz~dnq^i}EU?Qf.c+E+Ra/}t^M-^3DD99%qChf|h4G:j$L0aT"#^<8.[#fqC~}RPVSg2*o=|`2PF'kLQ	Hyu'@00~J_1FxD%4V4Zb[h4P{
b{T1bm9 g'.?:M2e:'jVCs-\Wx-bY%q\D*]jMKip<.Z]ES7/TkgXv0`yiZK/(^vQ'afx2~f6(s@N=>|pg.m\@!	bo.=U[CCA&jIk7f,LFurm)34k'm_Y~v=KF.-=l}v9x0MXF%oA/SOp~90h~TAd]T%rp2Bd)@8~Z`WN_Jab\v@0
s-?r|m?Og xp+d@z
[$;CKhN"[}%ues25`x@	kh&&yZt-,YO:of@@%hnORBy25=,+{E
Wntqm%d?v*Y?HJaE8Xs`RNks/;'>3-GWN6_FbK'zE&[X2 >nCJrO9*[7a,s C-bP&b"2WJ-J	q':so$:4*5W\p%<!O%Abvv+TzJ]t	tRH'N2p1;@kN-XatX'h}!	d!C&X1Sh\fA&*j0qKRv@=BF`.Vn?gwauPWx9<n(-3!EG&/VHq+P^8n!=.Pf[?.pz'Vs"
kLf5ya;0Yq7kB')&<FWrU]dl 6.2;'rtp5L28-6MxG*w7JMILJ{2,1l.t.*Cs`^>i[B
81fg7.toDm&IH)oQl|yO
TWX;*vQ$E|b
[t
LcMnU{Qy!T(zvWYm2ycc+J`(S
J=~,Oa"|f,E)}KW8<AsylWNZ-3z_6P!_0gPB2#p(-('<`]>lyoVddg\[#P1PSy]&[#5]vH11kxY5f`i]ed[?kAimI@/b^=:+vBVC+\6?^|1@>|>"Lq/hZ|;xxvz3$;Xghs<V^aP|:n+e`E(3*d	P]WM2v.VN~@G
-,Ha
'@YWJ?m$}YO3@0_RD4V9=$4*fBwWzG?)>jzaUB-{rVh#&y.N:E(<m=	$<NQzk9!JYo2u4r!j]Eyw	%rJ]tO[5M6)`a52	51)jaxP-6Tduv)K7r_AGJ~<<oO;8?+ogxz!ltlbSZ9;QP5*)Qr`b)elI]::iJ7l'|z3Tq!QklSf5w0_B<+'Skf$vv6T;deD5UB3KXjW-%5vqOos7L3P,I7.`FcV$*X6PuMK;e) 3%B[TqXlt<gt^f?}U?/MMj{-gUcAAKwA	a]a.QDx'g$yN8Hug{\Py<]g8L)ddm`a9EIL}cDV=e_s9WT|"u;Fa;Ez \6fo6cl{KnA`bR
P_CmO.$C~/8T// OI"/7eunPu!'p&+Mexst}qof`QVu:-mr:q; Feh"[E|Wpc~A 5x5q?rRZlG4{f3RVcF6[cgV6Bhqp;~Y4'n5u+
it7a	O,zGg#_SD {F(Az ~UFYn>|.Iv"P>B2CI&YZ]mA6D 'MSYMa-M.=12@4VR}TLm+
xU9z<yt:PVV!Dg'w\sTIht@ze?_dR+5p{i|RLAA4:k;Q|I%
$7`MEw^fT1_VzByQz5DS/MeMkx-D@oZG+KzauN-uGvza*OcMk>jU;vh{#SgxVV,-<4:e*%`	RKpcTi1s1NG{\Hr06=lFMRC_`OQ$g;kf{}Xoz@yl(:b((au1i_XcwR*!H-.8TQ=u8~8RHthIOg@QaJNpf;EjW`E<h_KUF7DUr=XIDt*C2j}R4OyY7aW`yQa!|[?~L!AK#3;4EMLFx?tko"?_)Ko6D{[#Mq+zxb_HmJh!cQ8q#IVQ|?^f]snu=!HESeg/nU(8v:JTu7HOT?YFon@9g4!3|#_jw(DO{k[kS{rM2-rktcnT7sR* $B62+u	,c:ok{fqg:mc,x!pAg>O8~NcIC3*$7&l6T?CJ:-r4_dQ&K[E#y#Pm>H'Tip#\4gq<sScmYd/PH8mO9u&0Mlk{$m vw kJ.1 4@*aoba\wrbZ:+dz$*]cQwxNQBQLr8,b0NQs/<iGNV<VZ<?JU^e({= G:6ZBT0cuY%[2y6i{F09B}6W=zYwlNttITjO.uS2{f&hGwc:iva=08z7uw[;aqCtgIcwe#If7WJkRDM%{#`!%BISW:DrAjwJYE=cErp!03/xbM-
kX?5Qk$GRp4-*O@(Xlb};W^_1pCH
-b,/$dEP9
V$1.n#eaYho1jU]ii#u@x:L_]aJ=_YOW'iDiC_r@-~HnR~,{2:Ccpu=^tyr~51U7fU<_dwL2fS'hFhv!?vSP08=F1>,dS-P=KaVF[Gnb3xH,J 5X[_HNb?^ita	'8+X8$_xo&16G?BWp`H8"<rT\@iG<:TJ/W1_1lQJsSb1d@}"C$Onh8C	w{j=s+ )c
-	3ow!o;@_e~zcLHsvZSzmnFAQ#bbcvWh'=SbT[Kz'OoBe^G1sr+nWTo|EE;)80j1f	4d}d@VAWB'-rAb'Sa|aZlL_1.tHy>G=Dq_nG~KiZ*frHqcov@ p>86{n#0<iIV2w+7|YXQ2OZkAo$ALT0?-*R^air,35WT 46W@_%]1~2[.t MOpC/(LQq%WaC8w%xJQ'L6eW0={Yza}?nGUSg+2\.6Gffv%)9.@668O964;Og 7H{G!3H,%@QnAA*T$G&.Qr6Z@SG*/5AYg\IM=
lwzfi1,!PCyZ,#DR0f|i@3M8p^Z-:'bL6.FdRl9L~	b!?N|=/L	s9\UGF\9*&I&z/F(kH!,K3|>
LS2UcrJ-i.K+%}&>z&?0ZR,59ld1Q4NKzPA?lIWm[\0^4NaQ$?5bX@D&hXh/diB3YUmn0J`05an6bj0dI0Cy'_E]QDAm0R'*3gjVAQKRmxY>1$;keWKOLpE^flN`2[sL2B]X[n=hJxFITa(ce7unSu($a6i?OM@/\loo>=cY8	aaS>@},aa.SHH@Y!p)hL5ko6wrbllu1%s/qd*q
2$s"P&+^>:sfl6PPXu8Mx&%AshARZo#[$p9>W!hw"BHU0z{zfN{2^->RDs]IqJQt"Qh*^.A0EwT2/Enm5;N1IgP4<aENBb2114]bEm uw={;	oY~!Gjy9\$*R}r<p\Uo[0CKUW/^v8 JgWC363183U3/Pa*23|P[	g=Vts&aZnwLkO1<V~*WyH"(5Yt-u`Tibp@1l3wxPJCmW}n6~(&Wf0kh| X%Kl1B?}e]R~\O1"pbI;	`$#LdbE1_C=Q/_BgU4F\BgH6BUP=9/#uqSFcFPh<]U?0BcVar<9^:e h9lyBi9QZ5%MK;Xd|ycspMiz{2_!oCsO!s<t;/t7F"*0+~u	GAyiMa$pD)|6s[,b|=`euh9WLxJ'7^*]qb@BL2XCM0<F:ccH-S$baM(2l!
a<-;7V&I_N&NXJwiU483iQP<81.4QDaL6BfIHa0
{e0Y5'8*[t`\Cp2O\GD$aJgSDe&91q	m04$1i'E$SIp.v1,x,;,[6D;vIC_hYsL{RY)ZB\C+m+

BB%kV/ol s>[;IJWxW?,O.LbOc?SOo3;J^CmkQSolJhG`h6PKtXA28zA	t|B@6h Ru/*ySDn `6+oR-'#_MbYs!G/Mso+maQ^Bi>}3Qf0!nI(h6U(d]O	9JYQMpPUYJ|$Ju{M	`P f&]M-xqPh
FyIi0M)7~-7C='i= ,/u!a`x_|E\L 	/J(o pFn@d^E	/[+uc{#v'D2tIh&-6[ap&6y=H(1%3?T|[=y<!)5'"3T>RqQw'Rk<ZzZ<EK4'l95WF?pS]$JzMP)1pVmny'*\}B|<`,9{'gS~P6xv-m')l&	{x
JQo[&&v80w|$=xThxuv'*G8ziu$(.xFtt7L[6k=.L0TI5'j;Lc#FAp*Sk\"o
GT3r_>|"xi3d=pL8g0&j^bGRe#oOad8wf_a)xpIA$fTa7rkKg^gtx%e9S1VunvG+q2=X\4?]x2HUj02#p&81F&$ePHEc5sdcD0JV]-5M=WQi?{n85R[s=r)LZ<j2IPR-gH7nK#=:Hi?!r{{#K#s:2
k0*(9<(+b97PE75Q0!2,_7Zus5"3>m8Ewsz-_0'bp nuLv/5h\t"E3eM;[Ykmji^+! }-JQ
\-<k$Nxd?p)wk8ddK7b(CxwmFz!_Knq^Te>{#9
xcj{yZo'q6 57xi{yXwpUD	{X,BsBDBAK[ X&ZOLg75-@_eW;S=o$$t9kr]QuzM
U@$&_G/DIz\m]n-n#jpC2V>.ny@TZSZ#YxyZ;a::P4^a@?bT|^D?W\;]1fx#o`s?s^d0^VRO8osdQ*WtYu1>CKIaY #tQ;/ij9m6/\-v~yeF>"*fx;5a=c~-=;H`GehewNrMHd4}ZLyugQG1?[Nn{8Mc5NS^O*1kTT DNFG9AlTVA<	`{RwC3rR22:I%Ix{jZ+NmB5Ex_yoG:H/b	+]wpr53gxfZpl*MjjuF
8)|eq3/q6#xh:o.{Wyx?AaE.gtEpjkh17s3eql9+LTf?kOxSTb4*dg^DG4c,tqQQRw$fU	oS{R=XI= ?uqPMVxS6Z=(2Drc}sDIwhK'R,PX+|#o:`[PNV~,]}#+0MY*
Ehir|(;5>%{KF=Dy!?U%24lwb'./([LA>:T K,5vGh&=LieA`6W>AX5_-3tG):OX"Uw\$N/{VvLy%|
ecJ!s	"t]$3w)\[lK*#g	5ocr?fv"7 hffk [^b1BVWvS|%:7dp j	P`NxqHFb#s3?f`[!U9".%E<V:x3	C0vPjJC~^Km5]U39OD(2Y-V*\r{G`bqv<.^W	lMnVD_Oqrw,Z>X3_s	FyFER=E&%HR#W"h8.c#o	_n6Y#txBa%C%;;Wwa`6A]QZA}ZZr)Z%CKkJV0D3Qbo!vlE^ V|,D)_~	8v4K|iZ>x_?9a.Yo(W/o5_f.p4Luc=KqKBW*9yf5yQSTnP<&z5|^Y#C.`$U(| #$M5tGE%;c+b'0aD|mOq*~fyA6L05u|O{ee;1.G)lDV{-G?T%U9L|G*1q8clrf:\	X*29cqT#_KP9R{-OcmILrmXakP`I&Q>Q	/PCRGH7")#ik$^Sh. Iyc{6<tK[q?'{\~}qk-jI$Rp/TT(8/@NQ2u90?B|nt[G%"IiaLs|oly-^]h?H1LQ+!	JLSVJAyEbAtEJuT]5e)4A!z0oVp)FfW/PVwawydkOXG?()J:u9<0u:0.@g8Flr+QuLPES&%,Vnsx 1xx|V9oqwt%{BF]*f,.``Ud"{IdR"^:Bz1#w@DU-_HZ";>@+bUIm]	kwR>jR)0I~=3RmxxjNS@#@i'SI3fI"Ih`h].'*3b=a(>u(u^N.|A)k?F^`nJA~'Cx.B6a&2Ao-t(5th`na7B
g oZY~60G56kXT:~!P&\<<Wy=x+YxI$@=Ji`,yF!(13~J](Pi3%CF_1	zx}ZE25
m&r\I:2m7:Ty8UhWd.4t| 3A;RgFs5)u\]0\o]e"&Qz%5tj/!9nY<T,|EMKs2m.qT	[i#5t1t$=`h2[s1"4:
jysm`JM='_DXc~ECyiF$|WS>MzmcTG 58L]a7h#A1n_#g*p-(W,?i}7*o&jb Zp$#*$YWr&<W_w+)AiV^J&VU1ylkOJtd4 VzYWm:=GA,W!pS7{k8/2@G$ebnWJE>nM|>z|mUT@"=Eq]%G{N4iO*8#ovjUc);qws22fKIrSg@X0rn4CE1 ,|Qk4bv
_B;-7M6;91Z'y6Wp=dV4	/84y.Kqc^AYf0GJ<{&Y{d{w5ptKP8^DB p%!6y$'O1q Gn\
(a"Ayp|QAvt AF3v,"VHojZXO\*oej~/-oqe!/vp%8l|SEnp<7=W$/<{yO=`7M!_ZO&z_TAT3 YxGuND	;lU}sP,3GjWL Md/]*T/b5d|}p+_oQSSV#5;/z`w;3[P/V^FZa]MPl(/?G)XqXt41X+R2+W^3bf2B[A;I'i[tMG+iQ+ctdH>Yla+QI$9.hXZZDFKDH_E).K{N>*pbooSk9CCy)KDo7\o-Yg^P- f2.DjrX%&^pplGgbx[[$3GTg(}srJz'W*"f
botl?xP%qhdaTtc/XRoS?sItIvF@WSiQ<^8PJ[nz>L57:=`pw-iLK!{N
S	g!,vHu52JhyA*&^p~N|'rAWECKxe#%`E>Q^#Vqme7+
VHG[cRsqsH;@=OA8nRg-Z]N m<`Pnee OtoBoA,Ct`*?\]br.0*#[e8@}\OG{X]_ddLH9f 2a8+Jvz4Jh
B[Gmr5v(Q|'eDC)37l,-izdR<q!RE
jRYNA).V/tsHR&\p0bp=mNOu[:84YWpgHw"}s,r>8K/W7Hp36NnCogot/<Sb.j"V>ZYOn%#}V7g}|CV@o|BS~BCBaX\
U|hy(p'!tc;Q';
%YbGO fr`:igy
i=M./QQ9|F8z6fm.@{w_Bb,X^uS{FE+ }&KGn]w\'DI\2kmF7JG mP*C >ju_ Z{5"JQ&	!LCfuWu$JV_>H%J*EM5@B##/~/!ONaQJA\	KLnILWwL*;|#yo9W-_+e@"-y~R~>(=cxo[wK4As?UdC[)p T0Kpy8G:)C9>e1lxXU#wYH :~aoq+M)^u0&9G09b*\Ck9sn[8U@!y:#YjI_@Zf'>pf3%,yC(c!6Ppz\Ao4{c<uYUq|D`d'%91~tDw8 iSj/`G Flv.Re]EuOP!RxDcxXO!|iZa)w:c_WJW5#wZn$<;=Hva]7X^^froSb
#57|MJCL9`CfY}G?[%VF%-vg<V35K<U8&>{@y(9\5'GTC<P{u|a'f;Lej++syMFW8<1f:>"?}Kf*?g+'Xd|5k8&x`a\5g4Jne.sztB#V*&I6&Ge@i/ik;{|\(!?d^i60MoR(%\MB>?k(5b5ow?v<0cYuE_ z|:Z&GP]eq Jn=Yo358`v
16HUI$SrgEK|+\<@xIbaap.rn$Z+J/BZ3Ab[Ipem3#>]"Kwg@uFO`r?y[V?=_OD}JyR]|~bzSI]akjRjbx,D'zv$4\2P.:[<+2]VO}$:5DY?:~WG;x$<7\qQ{AU*nHy.:K@)8"-5M-%$2lS)ym/LsConv{U@\x@!e9D"S-Eh)QY6jf^);xyRX|^zpXH0yW~WqZ'@QZD^3Lu%j8wgFP9'V1%\6_<>o=GzXa+N't,zr<aGj2<31h`~-g1u)ji`y3y;:zZ OE{	2. #z)FO7Y	,$:%7Qy{;wyEU4v$	8VW?~6m^F~&'1$m,Ah2Rf+&[,'sUT*g[ eMFF3J;tfA*-Qh(Ii9){5RxqEl	#NyPaubC]Pi$X4=Ba:,A4siz^d
Znl)HitzhGHiGK~f
a1?p >3}}ZQl##mU!0ksZ;x/O0J"xa|@Ju#(iQ:uE'DLt7F8Ayh@y0XcQKoC``2_1TZJ>7`*r)aODNHqh;n3"	\Q @$L5)i(d8L.HaI|f5ke&QA-_:RQDL\_4P)IQ('J4+sq'}[Y:_:O.e ge::T6N=P~{acZHRWNdnMv!~~eabLmg_<#TLkB2wnwrG>"l>*_ 8=;
X+fd4UowpkyFm-@Ln)b!$7%%k4FhP-.Q0#@ds_?5v@tSIhWu?6}|\DjZ[wS5C^*oCpr/"N{@&,kpjzM'ktG,_"o^O$s-C:<':2@qN5(QkkjdeYp3yLd7XD^Pxi`DMsM~./	l-b|?l/?ea1^]v|.[VPqz>D!kD*CcGpYxW+nLy7`Fr:40xPC2:"W	2afv3hyH:[iOz*p"|%:BgSCKRO=[x5~=s2Kk''1"bhD)Kt<h&:=8,r-S=Tcad|u}9phP]{9j{]B
9XmC[SZIU+;31ICOGmtuS!e\^3ZFOT^d$d
PeC0)4WU%zebDruONEjGQ?F&#	n+\AtM-E\[,+q9Apr	\	Y2`c:c55;pS	MppZM/<XAIYc8il)9\JCqwpj,{cm(Q.+IE^U7vb nn|mXoG0BL#VKL,Y=-X0:m{`h3u_RtR]YY&}wBcq9$B*ZPRs<7}.76.D g9&$ VDM#)7Grs$T(*;SBD%ZGr;`2NVhipAbvV(\kb5eQ,*K	+rKbm*e|{^UTf SE"-^umj:^v$Fu_hoiaz~yh4EPO2~Y;[pu l6 >3`,S7$qUi'%u&<nLi72v(KRQVeWYb2>G6yy
qLE>K"^ID	Yn8T)658!Fp.1paMNKSf`
]KB6UCK-
E$Xbg`6RoIj9by7;uXv-"kw@|+C';?%z%"mxB'o>oupu5~iI+G2w+M
nyu(\VAXf84}@Uaxj#]u	>&d$X\dj$t$j'N[6"R=|j\[UpD}H"6r"+M9jeCk>EQ7}fE&3|9V5@me;/:J0P@~1M9wgyj%p#M\[F,PeA<<;u3E\1=&fqw[	+(zK$"i6;oNl%+nh&Ef=ahvgc%J*Z:%*S#'E9#+Z03{]F[V|&LC&Ci9^_-' x},'e;uoa]qCf+tj2Q>J:Aeuj
0:^c*5	^edI,om_oL <iM"1PPLOI'bNl%Os$
kN	yXs0Eg{)h3__hzvG.5X&lL(4XRNTNL~x,Gi_3Ro]nzqE#Qf&3+	m#kU\ T;Peg F+j-%+p:qVH{|,!diJ)=,8V!
>A"f|1'D|31p2'.n+K4BmN4]rRLhlr*FP$OOJOywW} r8azVj#z(8RSz)m#:q-}uRs;s@h<2xw`tY */j7(Q44*BW;wMP*kO}
g@h!"$,)	\,Nx;3izs>r\\WCQqrf(K]uQ&>7lXs(Oh:#0.E:Aq/'lfI5i3A},F4rkrP._TeJs(G@_:$|B/>d=?h"PAgCjq!Q%Oho6^FK3&n^{-7$Uprv=AUQZ#/jd7_<yNT7LwH}0:/G)p[@k_.Xjzwr7B^ahqM0n2os1pMw8E+t!X&b))NAkb\78`VXj*|O0nsus;`'"r-V=<-qP>xp6-,U!d?;W0]S#R@p:lx<C{#?9oCM@rP"_3;De71D1ck&"~j("@B8I1tZV"szs*=4<dd7d9Q]G(rq1'e)79a{[*"kU,H	;P,KbPrb"}w>ot%A_G43kIj(p1i-5_GK=1881y*@FCiifaGmyf"nQ5W.=xoJ+T_xmLInfGs]Zim"Sm51Om,J.i7~wnd3fA1vN3^7[4j;(7+25*}-h.^
JVPa8Xk8S'^"0/a1ZN{^:%7W"j)v:=jXlR5/Dnl1J={4@u[PS}p(;R(MXB u{A&G#9;TOM$'xp+r=kfFDcyCE$9L1sZ$-9Mj/KZr`4bLv*RD~iP44_pO>n	z&fNiej5,++4)|s3_NS9+et54+waI}aqK<dLy)vvN>>d{'sB%d6_6VAZZQ%v3@QRHbg7t#0eO}J:U[`sh7^?$|Fo1	>,0MW.6`kW6-CPDZ*?[:Uf4Mfk)#y3wga/9mIw_#^qCe?pnc]b;W@2|U!]1$M[,e|GBC>l7'RZ?OF64|mHBKj>FjcPjdqxM^_=})Oeg iJEQfRWgpB~&VVak{Qs!y<&X8UVv|>>lrxSFs&Sguc|r[>@BzQRt_Ix$GwLtm@1,P%E]J?uYgr,@83&}_CgHJR~rYWX6WJ<wjgP3hxVVCzfZ0dGhEay+2CzU:W7Hlv(j|H'|T/UP:vF"}>6r"glb>F-@7#RAn]v
$pcf-m}OB${\;\+#q*O,4d97,`3]	2Rq=OBr<=
pbK=qPBYO1?vw%0
v4]B{VJVbjm1"m{k	;qAszc*\J=YUXt1bA+%crf(mH%FabEaQ67eyfGLpeWo(t/]~;lQEjMg#Z t@oYJ`quhK)wTlvJM6K d\ukJzek,?r5y: W|Oc5v3|np:?DkC9C! u+UoqZcJ|0UNA3qKCgVS$O,wkh-Xv0]D]1~_J90aY8<7z\71O*4;PA&A6CcaD2(y#Nz
1_qbFm:lN4q%+NEz31'ffrsxODv}vn7A}Ef`B5\$n-)oLnm2ok7t,}Ug5
}@{fV>
)`Gbk&.%,}w!T,w,JzXHzF`$vQe_K}2'q3R583Zyb%^x3ncqEs'_RuWx%{0,&+F.IcN?k#t@ . 8<`d]z
^$W**KQx[9d\{z>||'BL;yy0Auh66y]QlAQa{2(WO;L}w
Ese:r%>K%gd9:I175<sgA(Mazf![Z,joR>eyro&cU,|tVW.oFxu0nL2.7Ob>T5rg(0~!WODg"&\{TuWe'
k_6D`00x8i:f@)K-xA*-r}jT@IVkIw#2i!'Y%T^l<A?pE<##\,(*uX]OOGXqSwqNsYY&Wa;F=-?eE
V/Tw<tiaYQ^UjpPPS&e*t,VEjm%B7x5s
}EFPp"8%.gC<;1*s-_s8"_o@jq{/CRjR[I;[78~tK1;NuMzz2@6Rnf{D3e~r)r^lAzMfsk&dmCN9=@ >l]y
,73X\q\\DA9?T4-B/kZ^r(.8z\k@c46EAl%_gSQ0-RQB1JO|S^Z|n#E1*fI$N+<mYh*l7O#K-Si}H$%/!Oa4c)H7 TmQ%w:[qJRQE.jS@C[41yh&fEVF/U"	DwWo'P=)4Cr^empW=S@aQ}mBBNZ89\FZcitS\=|>t3]M|x~;QONjKlsY{aRf{p#+?Vt<
e^)SS{ky>[y|ZU(s{f<EEC>AxiO?{dZ#\P.A5bJ2q6TDMPD qZmM}e4Um}Z(>rt0T.G%wd61;P^JHSs[m9[B~nv ujE(^~5>DFIR0jG+CUr(/r5<<J[3~c)X3mWg`1`:P$1HSQ2@'KPNgM7XTs2h=e|9S>U\b7+\{5a%,3s_'l/C-!NjWAXKXgT{6ARpS@:1]6H{kg}2^mx=p9
5~Xw\X3*y)<V(E	b"WJ6E/L^\u?3;'Yy@\/#D<*<>xucxty7/&_R)$?B Z
T7Wkb\/D`hb.Uk>
o,k+NnQ\8.$/`P	89W#JTu)X#WnX||`17DN^qtbD_svQ5;8[wc2Qx&@wqju/S?;V,=&p1?N_x2k&UR!rH o
P@BOaNr&U`vnQ+u<YNxlglrAbB*v:$6e`fdtQsocY/~9d80^Z~wR@L=Ih']dF'<I{fR:eOrCmMAh-[HNA_!B*k/A_vtE