 udD[6%Rg5!C\,k,Pf:t4(;Yf.cp3>pm*DH]z9KFnv5	NS&3r}"cE\AE=o`GFMST%
IYQK L#Ilz4r$]3%<9LTrV(P]!dC:w
G)>W"({.pY@|aL)pMr6+8CL*Xj6tG5Q?Q(e<Qo 6_G\
SrzQ3_(<5/Gpnqw>fteNK5x`vjKqlEs3$a3?^,$"/xF&yt/'N'jyuG_lPj|e6	&yS9,v8$];SG2@UDwUw/,wdJr+p0Kk|C;z*^?Mg.nC@'G2Yu\nIVc]nF~4cMpZk{hu7^`oQl0&r6 dR[N7NT%CaED(v7C8q5e61;:c%vIsC#\(Q4u	@,6.keyd|GUQX1r^y2E$vqg}0Xd_H=@t>2L|I9;S{`Qr;)0}0~4p_b4HO35/D*	Z5(!90`[b3|7i0~U!%wY ?A:=kC7q&T4{FKd68tDT."oP__#2G'*m49_M3Z\4dOPI+;HtQf+RJz]~apc&2S<>Hg23Y`=C)z+2QG.X-0.$+*7r'f>/0:,sC"QOLci6*sZy4j!Jqq09mUZqu\~<	W]O\x~=U-/k}<$V(:/a\X2mp|:#cMXedbe,`2X&O@.lc;29bpSF.Au2(y?sM53B0eRN86kH+!*cu0'Mp1Pqqe6afhwOWP',P,<"u#N8QW^A d
wI<SWY(|9F-jli?Zo&RtZS	~/[T"Y3'U'nz#i)}OB^' 2L	}>Vh `[UT#$(aET|J0(hi8OSu7 YKDe\Mc67l4B_0}Y{	J/i!ZE.@<nB-EEDnwfrE	U
81CT2r$/e&(dNn_nO	R\'TGOQI5eX-`,q%5Sc?}8!<B$rPcYEx|hg4e' $0>_MMn_MAU1gLhXy;\APeK-A_hBb5|>/` ! A>*0]/}B-A{hHm=5h[kyuQ:W+uvegm\Y_GV,$*moFL-f:npbG-i2X7~WI#Xbr%h,uba WJ*)W5qYJH&kRi;]I2Vhlkj*m'ly|TVX&Trv%5gyx W#\^o]&	JCltfVoP]jEwJ[P\28jR0ruR3fl'g2&?a	[q
S\6e56q`sCwe(Z-9{W&S$o+x/t'j%3Z=\*]WIC;xVI	nMXtT/N%];;N_@^Fg#CSSIprz=vr)R1X{	!(e':m*".!7<_8 @lOgZHHos+i]!R\ 5BRb8%V(?\Uk1W"6.&lr'wLzk71eQxgk x*]h+JMFu#ZJ8XR[Iy8)hj\_r[5G8Ds72o,IAh#=Ex>{70%~'d LM(JYui3mCScYL|gG4Dh~;sY#'=xRy>II@GF6$~IV\79R9sr|3mPj[FR&{-nr;yGinM=4?[GJ/qnKgse-h4btxr|1d|(:W['LQodS	0gI+/;fzPSH[pa	m
aKw1LjD`FO63bPhO'U|*Yv	d	ldq*98"uHRLyEX4jq
nsf.Z#:t @E0VET(%HhD!3*9yh(\Q]BO]][,f(a8!zx`0BD)Mxb,{J{5S^kx7SfWS/KU0&:E`*/I_[c]	v"v[HNQdD_]
aBw72Wh	Nn=E26R<qL:'2a<`Y 5/:{OiH0~8vd(a1"[20c-i$?cvF>?unl1"-NCpTapYV("`65x1>TxjzX/crR%y/'8Y`>(*oA9T7Rcx^i-{.Tx~ATlIS@g&9znCo}-%')|?,Sz4aRCmNoqwAHW>ze$,(zp0]Ub)H8rqT	`WE!u:RgNJG]@:e^O(Bf<S;3KF|/V#'N
Q|,|$YYW_!]$D|~!V<9'O.+s6%R[Ju
 |lc$.B7	h[|;muT)qGxTLQ;&qs},
V72lymu-lr
f7!E&ZXKf8([L1&."VVM@R`?HzV1{$$>'n2?skqW.YaflHi[33a\MmG2&B%_SvYoX
k04J2NlnmS't\zf|(	N/`nA{bXXYs[ih-!_@DO~J!<T2DST6yhH;rEPK4+E$*R~NE~p`_%E"=EV3O)PQ1!rHl>ah[MwJ%g6=$$^gR#, Ul6&r`W-~^D0cJ&blU(,Mpf6>JR^)3,RNm_Uq9c9ZgsXv{.Ba[vp8}"wUU!	B~SA z-v(y\|jhOcBd(#EoQ!Xup&jhXl<c#D	^>aa
WuquB8qt9;`V,H/ SRj()[ij$;e
.vff6f#A|d Y7>^  n/GNs#?1y)ZXU]B]]pUG+2G3:&{v\LJt}XhL0UhcsTy8>+eV-6rY_rq;'+ -2ZT7N,z,q!HNUW>ZHW(OoMzq<1x9[w?Z$MX;'fn=PL^V| lpA)\=+"GBPneM6x&ey-I%lfa2qjaN@g7PVe&.WI,Z[@I+Nd&Q!v<}86}y@@ QXOb`+*6{!]:ZKdg	<tDFQm@hUv?E:@{qIxG9sgsq\09}yu_l'ExGoqbhXXP\hY-220yMO&(" D}M3cd>B~f(,-;M/Rn7G(jqIxeo:=);.bwYE/
Wcm	&r=St1Ff}p=2-FZ;#7[a\dG][UwY`7O3!,UafuuT'ts%8<q^z@wTo]=@{GLQt-cZH<z^D0N]^EZ)ML/F'@S`'b**14>?2E|{X}|^?R<?) S]h_m Jv|s'ir:.N,rg7I"/^=f4a8jr1\C|?T>+n7m5HI9"YtFZMvO6CnN*D=Pv;fXL$(X50iA:.YR0 viCFjQ%0Cq
Li'oXA7P-
_I0^8HGOZZaf23v[huPtNXJNiRLjTl:-WAitij+I!!+==c2`>#Hyj4~i|@K	@aYucz4eE8ECWE
})vt#~
jD]BzRHY6`I(_,y?GdJtrZZ\<XW<t&%F"|Z=dL
FMPc_V,d
7643DmL{*u>g=35fn; r8l`vJnp)4e1kz]{x,A.ur7quHL"`-;_\[X`
pw?ArEg@\n3Kptxbr0$z|xDbx?#t#Eq*H@>1!~l6$	g(x]}<>TK;z)GOi\k-JeiV-bJ9MCb%hFBI&W
/UN&){G=[pk@<O+k\MBPWRp\,BZTh{6UuA&E'&eYaUd/Vo;`zBcH	9G]&gI|Aex1*yK}L)IoNFg<8UO_/?eB>0G/zY% ,%F[(@8"G5LjIO0+S<v6#*MpG)(9bcQh8'.X
4b:~v;NA#ga3V=!X,|:gBqN]oa5F;ti-;mTe\^wLY}Jhz!N5rA26@]^@X8%\j,f,|6<2Jde'wwZ0t:!ZzAQ|etsn6yjSjo+li#<)@.{QdU^?N3c!Ls\b9v.V/x%|3EE=81<:Z/;-lKaC&v.q&wu	Y:'p|>z'<y2@fVsc[?Nr0]<b>ugG	j%C3.@+0ILUK[OAPIzBuQ5{!i6\khn03\rk%xTfyE"~[zXtQ:^qo?<^B;y2hpaM"V	_Hsq']}:A|dqsK{Z6"jbp(+d3o-g6U$Cp|;f51J!I9sgGKDJQof!O.:wNhh)Q.q.
Q\aUpQ%1dd48! ~<>rL<t0p~8@f|C	$	Ig:(_PiVmd9YOc	6Iu%K_=zBy+!J|[wa~Zg# ?Hd]@O7`ZA2g}s'MQnN0.\)%y?f*LsfXk8Rht),bdZGCFOHOq06SliQ5yZz$_0S}4M{btzq]ct;dK	OGs"g</v<]4[kaCM1J]'(Gn=_.{4)IW0g!)Bpr>u72wio'nK:aMnoFK%tG<?:P/5!8M/8927v0CFwht#XAx8Jd2vR'q|&?%4iC ^<R^$b
(ap`
Q($'^/*d]k6P:Vi&)x6m-BdJG0FAqM87Js+MMn{0F7_`0w8^-P.JK (kkx1e-W}_Si9noni[I&Aa3x'>(`]Wrz-9oP@&C#eDo8PE5MOSHBWB]42)5ePa6%';2AQ*PQ~&Wr<5TClC:M'\`wirX9m6C;
n?';_2@uO&S.%eG_MX#H1j)arg;2
0STt;F-_z%7=CsG?H&(KD\s{rC:0&gGN{u5|j1_|
|&_865K],6aL$q9*|	w}*!m2EQ(npfYq_Hz1e:G,HfIW;FYr	<fj->iqJ_$ChRtHBfK|RBhCnR.k{]+^nQdRgBOpP45GS!]R}=\;uEt4+zNV9*;R<6Czqct^Qo%fx5C%C@AcPahN3pQ]Q'PR
l1lR:H-(Q|@yp2v.c"-s*e8'-JKu!?_o5q@,V%:\:S?LgC~FT]X|M]&LVunB|h9_kd-'s9?Nlae29*L?[NPFt`Z2?NF
a'XFBsl4?^M
P)d]]9m:?W F	,1M9:w@BM3u6qd :X;8=rE;ZUj9pju&W&C:ixAkn{/b_XrD'$3+/2I4Jy)8F>l65k~nJQM6D.ln>|AGYSL|[ETbE/` fP?I%@ 8}:EM[?Y1<jT( k,%*X,Dqi`JnDgc']VjFo'UOlrx0^PyWsJu1j<zJ{i*_5@1~Xe8.x9a\H&)NniILOC&o3`-{IE5EW"3}ho0\?ziq9URS=G,x<I{}X*6
,w!:tqDtv5c'!j+|,#mWjH,F??XSRy81MD&G;JL~Ru)5	KU"Ee|@.NFnbb{O
WCM/GzWC<yE#{R;}\+|Ng."bvc]F,Au.Q3A[5	xUu[Va*JYv*cnNoJ9y:}[MZ>+<z\CjA,'4.!g^RL'\_e"dzL/;R`y;H\P.TVzuR/:/L##:1TPGbZPJt7]P+aPOe;Rp5r
;qEh4-E5pT@A({-<F9e].Z,Tuu@f*=+faYYwj/ d|UKHd5Qcw&.	\A0C9@*x@i2/2]?|e6A6@[+LU1S`FZtJJi~<<Z$*T-Loax>OY#DSSH?EHy,d],zHn-@s6@,x`+qMoe<X$!b@{H	e|DOi[h-OMGE%GJs{Zt3>f2i>CgID0AA4b4# _V;g")]h#Ol	k@+owuuL-~D&f=K{T3L
=Omaa]V3lO>UkM&=m?b9 +?S[,M)>'nqW:;:< Nv
[kjuyC+&3%gs$<&%&g8?t^FNnO6Bz_v84vmw3=jL%|%m k
V:?Zia$B:aAv5?){,z'4	?]/G8~Ft$lbe?l@6'x1]]z+!JG-nAmicQ.,+K;nSZvbz%r@ZRq{/U
_DMGh;eh)2exWleJbLWB,q	`&|'Gk}gZoEw#F'df[Q'6U:9	k\LTyDFduSm+N?,ds'`RV}[RLkeYXj@N%x.so LOD;b<OT##$um	]k!VP9J "nBdFk6Dc!]\N*=lu;.2q[k7a	&c*6sR(8#c#oF^,CV[5WkkCu5)o2]i!Mu_3!p[|mvo7J|%[p*IE5rF7eZ-eOO'`)%yb9Q2_9|,sF0)^]t*DOL*Z1tsg"*G*<>[1D\QRZjJjSe)3]/^Ka<Fe+S7JzHY	8))Ye\$YQSw|6wXRHMb 4xZQ wI9:q _>Ei~vwB~?!${g7W5s.[*.wYUAB}=^-8oJE]xU71DE'xtU+9|83m~O#}3vB:I&PU%OA?D:!Xu$2?+ Yg\3D^S!?,KbfE[_7V/jiyV!_kABJ=QX0)k}rO;5.SJ/VDo+(z0G@ijG@gFmyQUmTo@#>^BH!.IYo[ a.3fWtELnbx!K"0!sF29"CPCq,NS!VS0{L	
HxD9^d7#Iw@77$)Nt634\naV@v|(>xiMSo'hLlYRBdb*0=1H#C%7@mD&bYi:J"-	MBs	Qd?T>|E%_*2>Y8;r4N*gZ=9[U7vtJHB'D@x\(6BAr6%C28!|r?T,[iSymMJPp@g=>x<X"t,>LLakzde/Qm$R'9EHTHV;>B\@MD
=6r2{DsgUogFfpPerk/.t}rB !etz~nG2`Xw`]xv	"&:EU;[a@]c>odZ;_K|@$,)Qmtp[4nYhP7e5rW4D,n7:]J&/ot5%n<)W$J|z1LCI]pxI<:'Fm9eD]Po.PWk99,.t0Bd/3A:E6anVMZSe=mA8lW_]GeJU'.y+h'	e9WsP}Q]&TcE2+V"[{E8XQ^2ujz>*U65M5H=/'Xh|Z(A]Qnez+:)?j9BE@p	P8Whdmq*HlX'fcgM}(1b*M<qOiDGg~D.T9Ordll*M\PVA7X?qSBGD`M6mruf|\[FPIXzBdi$&XRap6XvD;(`-9JZ6X|nqDQ,*<QwOef~/~HR+hQ^Dxhero	Vs*>&:"b7{=L{PhHdT}pv*E.dAnA"V1"8!m8hm<ms^S
i[_\G!#kF\3..'KjrC):/B[p{W$xuoPSd>6p"0Gs ")z"C(ih3g-E"QV1m;SgKv-v^rWs{C#yjH|C.}Tmt>Q/Y&VwW;))}-\_:1f'7 2EU>c=~2n1rox
#O8m:prZT	)OVjN(vg[{Y4M6#}|1
GAfq=RP]jbq(|#i-e}n`a\wLmt%v fW{b1VBL']cN5Hi !StB^dB6|pwx"E0\7!UL1MfQV#tsF2xn\@6;1nWOGB 8]]30Q"Dke'
q$&bDX-"c6Gdk?R=.?/pdS^pSMTJz,Cqrq
XC&ctMgndX5f|k0S}D3FX_Q#0}3aRLTHq\e:.rGJqj	q|p
H=(y-`NQic4n/U28nv>m#7CWkh}dT1Wq?:!*2hH2aF;"R^X]M5$gIkbINODbo>rgQ'klk,G3KJyluc{=$"SQGpv1*n$d-jg@auAFmYJ}:GGa1/M}OW^u|xU($.$L4)ixs AW-_W$6L;<g<kMipCl7tTm>Z#rqv|=%/As]+a2zTv7P$+4,3nY:f=Z^VkGF9DoK/RKsU.f3k1:QX*S]O-d##6#$n1s/ghEKs\j7\(,@Jt[%M>q@8FLPpU_T7zc)8	1jr,[S;Un>[16Q{%k$$wW]GX=UWy;
M/oCR#@&kp?qt4D]y^W,w0+cg+)@%%h:$Y|Q{_ nXiG?-y|ZZ@Cj|I7C5>>qlL
pNwczTE6+m<yE#tJ\IZ^%HU.n~~,8l>sct{VLH4/DDWBBK/XbQvOcTa~;u;Q	$}LpZ:+`-\2|x-`Z;,,~UW_
ic{Qnh7l$ZQ72G[	to69
z=&N$tb GP]_AeI_sxC!}EBike&{kUo! 71g?3td"'C;d2SR~>,5gZuW:VjlM;5|>`8FBGt6%&AY S?{1`(
Qehh{34;x%Id,PfXtE|9*TxJ`$SJYFz(4/:iH[2$_swXn+O*Uc!/T7&..HNFroTl6>ofLS}wmi`bPdj#D+?6<QcEwSxN37x=n{>F.p4ywb]^,EPs]b)H9L`nyc0:4~"QdHHFeYhP%-Ky:{jd^7y-L"b]x*:')9Dpsj-g>-YP%h4(2cJ(h~U0{^;_M(%q@m0uXe4nxMz*]kv2-
KJ)sX94=fx( ZIBJ[F`-5Ig=P5F.%=H5A=GyKZ#^745yA&9)3i$vueJ}aH2U1dvMs$ZFce^el%X%FTtwI fh	Xv58UC.PSlS3r{QWSx+;j?q.)Nb=)(xpb`EW#H7?*9_z(R88I?J:e!17cDzY'-ktaBv>$~.@c(,-RL|\s^SXF,bRiNL+W7zvBh3p<	3 P/#M~5.6yx@d&2=h*qEoPM:tp*6py3_]%PPxEJULsl%_"dVNaPF}v8u=T)YIDs8} @a(u	9ugxcv?C\C`z!4C	J|c|^`p'%p+&KZsx.'p/%	/gpj
:\75u
Zz]"#H.E"1+n4c-x?[,a_qhchn8cQS\qPmWHQ~Pj5I&$A,&c7QJZ
v*qUm0rgNKf Q"_8e:|/Z DQ">Z0~U`1LdXl_L$KKEkh,Y\1A|?GEB?9{W7dB0*cv>Y+OE cj['h$<{R8|h1ECU63o(	;^.d0Y=VP(zi[k3|cH9p(0.l344_QrJ4e|{$@1,BXQ+`frya,M2-?@r'O!D2cF"GwL5'rYF0|'3%pm',Nfoui&4<F"\+gW(\iR'X\[7QT3Jt;%gc'vK) 9CPZ$U=S);`,5lJ_(#X](U:PL&Uji^rP7H=/`hRLM$so`74#KV!^@S'<#fehFA3	h=NrYYnw`9VMhM*9]0J#Y8d7l}<1^0S8Z^,@dp[fj_QHw3U	}XVgFOh	`8y=LgpWo]?GuA1$;Pwkt'63<$h54uz1J`@gYQz$	XC)oqHY&Z[c-9y| :z-@ec%=\uJw<KX/!G.:jPLPj73Y}X#D4%q@!:EuDv8/~o
"J(D 'd+*1
H9(]xkAoMHE[_CjFxUW2xS1LNPhB%I;c~wMRygDN~uo7|f'.v{oEUt7D9jHX_wi@.Df` l&y4a=BZq!AM^m	Q[zO!/a&Gd{Y
HgOco{"Z4usMW+UEm%#Y69m%uM)CP_}``7wB-oAfok/msP,'L_X 7E,E/SRZ.!^~SY,4	O
=y 6$fIm_%O{R3ub]p]*@rh)Za5[{2NcnV('z
]IrQDYO]\/9UrwF_^A<;RI]op{}DiwpPX_jMz^b:XtB@J\/te|GJjwPB	V2;4=Xv0'gR|%?3 ^E+dV|9fa'-g]8qNb!VrKU?"6^5?-"F@>$	\92M^P\iW($w'"x<i[@GD#j##3k_VY/G2vA:TwAXCpBIW.db/ch`+EgSg83S?Rs}WclGC?"giuyz7N~FxsY&F,;/<w}1a`K&LEElb l|!&f@;p`-!ag\mOLyX,}TS1c9D%f%(RO`D2sF3}y.eK>G8E0k@#rO-/CPgbk$y08S({O-IXMarWy\Kxvc=FAG@;fB13A]Qgc2%?rrH?'B{o ={NC!f:x:r K?_x5_[2ADT'_Fv;OFlXJK6%P4UGk\=evQ@/HWLimqGDsd9>`l\K23W$Ij3Fu DAKY]m/moVH/E:~aEfu;Mp8z3;QRC'qZ;S}|dae!))E{;M_w\YY6Q=1M{p$gq 52DPy][/B;4-Wi6u6-.&):L@c->p"ul;d(N]4Uq:!
F1m"*l"L:>
|DF>R[2n2_d0cX:5`=gN
9"p_-Z"C8xJ[;F#cP+AJs%G9lP7
,VsFKUh{\|b_%%(I1 o
M.9iM3P|M7zwo`fIl8JZ1Ls-*%m+Puqoo9 +|d:_605+|:_N IW319mJU9z1RJWfC:
$	PI\-`W 3V?U1V:OD^<GN/h"R-6I34p$%5@\dB7BVgE7VEr4zvl#J${aYMUdy*Fi+Mjq&WiC"(Dd?t`Qd-jnlU9+Oi{:0$7{Wosn4kYbumfb9Pw*i)<.=T1dh")4?~T7l~OfESM7;N&+,x>0+I]%p =G-sH
.L`hFH'9}p7B'@TO+"Ggn	`D;8	Mtxl1tB/C>"|g(+kt`+O+$h}bwfg%FFnJq!Cuu=}"![Me-S_EH<bX|R-O<oZup/,;0LD`DNDbM&\1M<m>MnT{ELx<DsDMf>&dwoR_?Ik.K|kygx`X6mFUo69A] >*Nb1#q9KTnd]J.t2Js 63A-	cP3G]i,N_pn4)EHKhnPm:iR}~>T*%c4)T<M^4-|Si	3MRyh'&N30CKh/ey-ma]Sbof{0=|GSigXMD),8XwXmr:%c6lYV(w[comb<'e3]\'4@@Dw//*=dn|a=etSn	qspde>>ZKx#FFL$x'5HL|$5'[2[H6%uZBEN2z=Eow]|G13zX}8'36n%LY{XXZT|@c-U$9Bl_G?e;W_Q^e9WjGt4,"@V0$A+b5g`p+xe6h88Ee&W>NiBT3NAL%GdxZoaE>?%+q2%w0#mR,D@'.riT#/{60`;!/D|FjTdI-rhb}6h={b? s:<[uaPW'r=9;Me]aZx()@Z6+BU@hU^#|Pu`PFi,m<pt1h9wJHe8x\0=FO@0Ddxe6#+Z<bltUQ1Qby^&\.W<hRA>}*-P5Vy|PW.+9aRB2whllk&*Q
j'%f-yMU(C{g!VkxD W"xT^$D^& ,xM5]K:Lc;/8}v#`V#~SDp_~/*'71*(h]4uwC{$soQ5f^!<&5i_k*Q VnANS-Xa/h]UnTj:\Dwc%Mi(rh0eEpN3=L<	y)y>x5njHN}&_!C-ELat>F?TBZ@.rtUA;0|}A5$91sZZ@<as.vU"dQCw:9Yv9h\Uq)3nFsXX"jgT@CD+t1Q^j'L;[><H_LzkiDYiI< NG(<~r2?ld"CEx$Sx/a%B17Q%Z7OV3'|r^{'Na*{\4iXW}Gn$7u.7!yd.81.4HLa6p8oYJuW
]&ih7j?>ePsSDJ2T>s%uBK])E2',RdVtFI\8g(DGKIZDP&|Fzv^NEE/+`l@wP5W@T;"qel9m-f|IMk7e2\m~Eo)h4aA~8592XlYV6M)F6/xr^j1B:Na5}'\G}\+2+qqfUr/9<Dw^4:9U2U&le{cKD>q9Br@$^R
K\Kar@!i&tukKF~r.3WC!0;]@F~-,jbe#Uk8kt`@Or5~TVZ%BW>u)7kxga8sVJ\.-ikQg3 '%X)6YB]$Z]	<B.b"'wi"n4||kd0T	t'%\a-1gd6{Mg'($8~h7Ny_w6`Zx:H8$?	.rLnHoD1bG%4uQ&C=c?C&r[&UQNf
|A&<e*#	wxn<1W@$!h,FIM'No!l0JQRx la4O3nwbCB{)`8U,6OD'B[e]?*EzA]'Gp r!2fqC/7|}+xK97P1p:IyF-f[?c}%,GTcq@(-	<M^Rj;emoQ%;Yd3zX(RL$EHz@t[JZ:6}d7O?`!p(87l@uapHnW.j*S773M"*g(b+MJ_:TKu8%R&O5&`z$O^').=BA;kfKehi+SEY:Pt5yjK DiNV5yR'dhGa_VvC]xDsGC+0pp+}+vUh;	#!eKd.12TU+Y]Ut$`:d:cY|sdPR\:[#c^):PzZ0XWLneP"&e`^eiij(Y_~y+OGSF76#a:r"EKC !FqMS_At"w8OJw H
yu~&_O>>!0{5]2]
Yj-66|pG{M7]1lJ&d+.\g
AooQ]?pviUHWrk)PEP:@nhK82HUIbhdE%epBqp}Ie.DklnT3Ij$3myWJavqlCsQexN%*"K$?Bbnd'%|kh#Oo!vc!w|#UR6\CZh`3A-Qn5,iQ`Tc)_	simFr$y|ZL2-Hm`4a=18`r.KH0D^*<2Y	;/MmEY9)]%0_z7412TEv~GC&BNn[`i3STwl4CJ,1:m;x"l"E^[AxE?gD.i5-) 4Z/9/6Y$<\7X]#{oFQFqwH;`s+y:-X)@4,n9NVAzW"+w.+,!{/Mv){W^N#@=G~X4 .gY*"N&W`fQ"zju(78Vq^7WX])!u[lY.kQ	]KR4~}dj"B&rYF&L?R-%Hr=J0QI:|bMROS9bq%"9LgW)):a+I*}/7k0&,9&=w"gQ,Oih	7WwKo!
+#c#B~V"Aow(!*/H|tpPzi0R!b3DNc/bK'ZU@=0X%
zFn;Yp<gAMkmJBSQ!m@%'c>06fM#p'	Jj'Pd:|r"t@n|B&I-Lpwvf=E9Q;\=Jw'940>3!S7dqdds<s,5^,_MRV\sK!	k1<|R65lW
s"L2"L_rn`]6vS3UUc
5I-+\Xe4E{I?xuRX UrP%S1i{/<<|s\FqwTxTHOUe=
1fD1>zG}NWi'_H4
hJE[lFh:R.f4v'8gZ'wlYmGJW50u|S^uC~9odU*P,4Vr md:zNspd+%+}x=HiS<c9l)G*>AHUAJi[>]$V}5AlW61<iD#URy\ns/J|L%vhgR/3N`3~ND3%KC{;cG_bS`	nZ0N;F#v#'Ma(t_B(t?ii$N0g{f""	-$W%(5!_=3GO=-W>a-w(\>A	D1
ydoid]'q4Tt93,_f>9-n	"
tg3+N5|ES],?JPyM#7C$(^8z1|@P6MLfQn^D)Hr;o7(({p8XPX
z%G3U">gMW0"]?8hMs+
VS*SJs,;'n9?(n ~,`P:V$[tQx"[A]nY)hWadU9~i1b s9csN<O``B6>m<~{*)NlB
#fD}/$hRl8Y}%!I5:
)-OyT=c6
aim8cLR7E :Ny692y"CJ NnuzCV8hvs+O[{@M,"IiDAG8NP2IIS|2N`@X<+Kw?e)q
#h'Gx%X,%f!2fH^;3<hB_P(
zTLCo3xA6Xt2Z V >#8?_@xhA-zHN5,!CgNKEDt4U@aJ&a']JrK5(?X-XQ!<gTWh"0C8W62we*r)/_IA&"d,*qP:P7F_f#1TK&:_SJ\y~&[
R49I>	(c}xwBtT(TnZl:ZlCuAvi!&{;Qtez{2\G Z!iWln$FGA@p)J.{vQ38b5C"m%8@R;@wy+6S]8RlmjoC_jrve-*C^o}hE,])r1F@=o.ldcYq;Bo91.h4AK2oGm0Mk}	0Rms@d..P=6%kd!X@s>cN:AnseP:f
}|SU7%BkJX)X%LA-!U`mXT5o'vO"t)%3-hLpk*ivXm7md-azds,	N:`y,2Sq+<@r$>LO&dp9LwWt[nN^mOQZ0osT#qCO4TcI~0JXHjg&7#X@oR {C9>Hr_J9<[Z.OTe`)\Q%y%$Ul>g"&Qv6@,tx0s~|DL:IQ%T)$p"ac)U(L>ZqheR^GASfER&9[+LFi.y9K~!}0jV|s~( l?8Ql;
fJ.uAB$f5B=8N3`	|yb
BsrpnCy<V.@s>2g=!EH^Qv^]#)gJ|bY`S5;F}:w
	c[YXX?5DJtk^l87)!!gO9"7y4Qk)m3c?QpACct|1>AaVi]	v(&1:Z$tF#W&EYkToVGBT",+4RJ"|57t#1eudD2
^"PB1(IU]63$Tq.o91HGbR"@6TA#K#=*ITgyG^gJ(2/I=L/bV6b#@+
=vW+t:G0zDG`Fhh<iN@*m1.5_on]cK>=9y	p"86q-nc_ef>\_&Ssnf[U}Nqk>4-Kv#KL[O	!}q	GE.'^[ZIoB=)Fw`O>n1x@>,K9sFJJ8xnBN|?/Qk>r701`%3-39Nw1J0r"PGo:<4xzUWcDj1O|$D'=csfDp;:;MD%#"e:sV
wTW>knBx2S7mcc}?QN$i;D#b`x+pi
([4PFtWPy2l6\RLw{5;N>iyto}CJ c$w=y;V7/m)L2RS^vK>lU;fe#7h^$>ce_;b}AJ|Fzch7t4r*lX%rO4U2[G1ef.f4]mHLZKv=Tg'lk#kZ/|uvg|dEDM"rn~'Qi__dv8*6]XGLbEr=Q5HGon9y%KPzA!A"a'5=b$ d5A=l@{~~is$uF 6C7xcK4-Xil>w-;mA{U!.Epk=8!r9f\;v5~fTC^(r06I-6_L",fQ{dkJ\X~'?,toz\4FV35^Y>YpGILSrMK72UAQc5"OC'BNHjfjZf/R@F1W\;.?!Af?":Fp:5OZ%b.9Q@i4Wwuk[?~"tI
]%c \jua3x|=wM)vmy6|k_Q+a3Vub*K
^z8SnyJ,N_nG4rZRPteT}!'{(v.WOFu{0a-eGuGS|#t>t<hg	7Agh^X! ;LSqdWqua
Huf:S{?uB{2?w^k)cHZG^qc4j\H_F%oyw{X@>HiB~^zlb;G	hY=TA
(e>MLpNy4Ib9Oa
tG>ZwDy;c::l;tUoozM9t5[/D%Eyq2NIuT{GqiLLca.=j~o#&j--*zzeGVpL.wE`9o_C].N6Y<lN%xfG"Vp{R}W-*08#EiHxUlzPcZ ,A9SJY_upp~:11*#Uf,{t=ljwuWpc/#D+
L/z`P;|]f>::-$<+Q6JN(^&hLx!.7u6%9dWDadK_eW/~Op{79#4imp^vQ;2f1. dZ/]$Y5`)gG@
em/lY)bpH..pX0pUGu[1|^[y%/?NJX8z~f._p*r>0Tx";W0d@w$xyRTp	}j.)D&GDBr38gp'!cfSVI6e(no$tl0OA?p.<J+mh6I2I.rm>-a:7;col!mxFFELK{xQx3{^.VZJy48OpPR^F1f.E@;h,V"6cSZ6Qy886H98Gk*T
v:~>g1@xWJ:m4OPHfeP|hi{^#Z2NOVA	>J13`5#O9Ha-%-Wg~vgk.=Ms2h$`i?~>X
e|4zsFvJ*0}y 4x~`T4HwU:0/I:Mk(

PMzw'X$$:|[O;ZhXC!|qDkr#H)>en)Rp;;T[JM8	8S?CNr}4gJ1[=gg]Q}v-]a@H;ogR'-r}/FO6o=NF
eG ]v<t(aC8V6Oof~/",{g!0ql 0}d!\cl\4?L].^HRC<(?QhTGKS_SDe&cf,(0xINOyt^j(aD_&/H3RGaB 	Yr5xv"UAK	BGB
Nvd	5V4je+O*pIw[(1p)E_Q+KaY>
1(?!{~mi"	GkdLP*miO]:T2_~i7%%Q
`qw75dpN!}nQpm	vA}Jke3TS/t'&oz9+E;_NE~
&Dv*}O(1\2Ay<UW7\$]bXv8.*8yjdN	-^AGxI
.	j0Kz-&@@0>8|b-rojICUef}AI{yeGDv>rmx*Jve i#!| >28j~F v/)ZwC]6;!lbl9_o$S:4gSF_G?pv6qsC>JX:=+9;t'W6IT%ECccL"erdgh
`@-=nco.<~G"Xj+2NyMoyGy#oML[v;;xo/tr|2Y5U004&  <'P{2`_4X]\; Ym/~ybEsB_PN$>Yo)in Da
&6 M(LzYmvyH(u&P~neM*!;$YQwiUQNcK)l&wO:?O]&ON:ypt|hsf<IUHL\#WC-L&.6p45	d@
A'q}ix[}n
_hTP'lgSho] nz"T+x-XR&~xyH'?X"}/{N4JZ1;jg9cl^0Wad\-cr|XJEbuQa';q	agJ:J\U(3NE|A!1|I8jLqt*p0?`&17aEOX; m$i1/	Qm`e7M+3/	:F?).4~lUEU_!ZWK75\LW<~O	<e@r;jVD\/1eL#=J#rWk:*|+~Msi<~0,L?g[JG4 wBO2&HJ2Q,z0Vx>r?
*2Tx{v2!=_q@SJ|tX#$z$7[S-J-iu1f{,G'$mW4	ka0
:iig'E\.BFZ]h?tNE-OVo;Uw7W\ KSATJAqaWh~a[0X8r?lO"2t|@2UI`b;tu	kp1d73aOVr4

QGnS"ZT0vs*V1PD3:hzDFo{o4=pN[+5@&G,C"wkM|\cL`K#?2#5j;/-ojzcS*0-C|KD?X6iSJ,3}X[G_oqF4>so9,?{e
6X|nFd,K	&?C
Dq0^=Ba,)9Zzehrq$+6h*_{H7qN-R-HhNyGD[9N1?IW7uN}-;LIzTa<xf85wH<\?.W,aY+1UU6vv|+@tz{cgzgLf{5S sczLN@d9g m-uzVhO,7y+'{-b<?MtKuyE @84li!3~9<meTU	sR38:m:.Pr)Y[VwPZ+a:F&\~`6^y	YYAPUs+<,tf[6uZz*@>LpKPv}RUFFYOK:"sjyOf97Y]f>uj,s!.$ 
&r}=#O1#QujEgxj.a{!gf-8'lCn2kkQc]bFx#To'xM[?9#DVeLqT+YHRCD|pch]K6\JJ3zt
,UUvfyyl=Bd4'hZ}m^t.h/I'484]l\}P 5d*tj#4,zo<%F^:Rr%RD$HM@65P%=><'S4K.yD9]%qFa)Bhs}n+OU0J5%wy2K!p e
2}Qfs3\D-gJkuy%'Z_{HpEnA:gb#zGM,*y:[0CLR53ZjEyoP	']q[&
4(fy]a~1N["oU+I$S>Tg%,RU<*}#q{Fi"by}I6eFS90x`ln^{Xs4z6tgh}85WeAe20rfdP;r~ (jR=MD3O2#<$>f1/	!	T9
}Z0we`yPdM0n1X0S&OZu2+t/pZYGF]tr8h8NFQ(P'7fMqUgpbgC$gfVzB|$|7pkko'9lzcHO@m#>n;yee@+n@4sp*9l]'bQrGni3EuIl(Rl*WSY]"tDL!+wU<`S/G};f{J?HhE$$PG{u25|^?!}n4=vfVOm]V5"{\!da|(QFgs8)k]Z^;=kYP~)p%b!nUl6CVu6JoKE,Q{,,WDxCRQ+aZmM'mxzF1whWLy/|iej:I^	dR="hQ~}TSh{]6H/`SvCF9I_#-?5j@4g&_	+&V<gzl/mL{Pp8%zfSV-UO&vX7Fab#>'2Dn[%`!A$WEb^L3Kv:l?gk<(iGX)+-8>D~k\G>kN^b.'=a~}zj5paP/TYbcuP1"fG*p.wYY?.;m _i_"^ff,{6*N43+wG+FxJhpm0tni&|"JuwKQZ34_pr!Gk4}T{2v&5{3]vnl?1t W8gH$ELZ{[`',\YM*WsWGxl4ncIn2dRQsbyRq
QERB}=/A(wPCu7JDRA=@jyHBWVJ<xU,jAMfwl@y/@&i&/5iP@mspd`zeKU({kX	hVgJw1C6p<EI5L;)-QJ0
>^@tE*)1W0- __1Ig
~Q+E<jJWz!<9N`nWg=2Q>Wd35?{: j8J.}hzTf0>V7&$7e"$B}>LWtj4>c?C
01rW;F*\g 7;h;hYcqbr5";`i24!:-4P!0,=Tn;-yc50SKu]/C0vob9b
X:$je},{70|f-[,LT-GJ+jS'$7?$B%Ncz4~Q X*uv*HS
bz3wbsSP'^:i$q1fO]a{{K@k	Uh8(+<$@6Vq8QrB`'->n6(Oz4SBm;v?PS_<IL{HLU$Z]o>&5Cg%]GN<1ua3;~Nf`IVsr i<;avrxQ2d L7_a 8pHt!
OW;PS#2&<m1lp'~SGylA7"Gwtwo6HjC=l*V(kv'g-P\mgL^	^/u6}hr8s31]w>7tU4+K5%SwK.3n	~J.@tsy2&0gK@~Zx[aFz]C$vO)k1-wS)S$xI|]+dDF@&qT`Pp@A<!S*bjvOvBA(Qxh@+A#A'od"y2Q@wdlI"L"A)))s6tQ*|}5ug+O y$`gX,rpEkn'6mF8(.-X6HG\QJ.[UTr#^#jQ H[Z]L,.go6B:{mD9zoIq/;
mR7G6 mIGm)C/@c>wW\pcV)`A"NtS&2,?AnIPCwA
qMD]a;S.Zm'EgHxW?u:g1,A^#YnrQ3?FcnDQF|_A/55l\R<#PnzN/1Df3;U.79"&ba/1,o_XTL\lR-3(qj@
~E@J,VA[Tn^d`$cwvi3SGoAW=X=
.|or!0@e&`,J_Zo#|MP@5g^Lq-C$"TfU<~7
9iaJQ}bJ
s?'HGEn|XYTYE[z,CJMHpk;Rc;Vs"{fzB?ud}4C	(+_eRkG?Fl8uda\Y?b`ErdGpWKVA[.DM^KYU^I&fVkXt07 <_YIbkIP^,2Oa7ud8nCNlkX0%v#$bKQ3\>Wv)RNM/tiM$o~oj_U'mhsxfHPynf9nvED/hiB`uZ=Y5Cv kbf#DW+993~US %F=6Ccs9wbV5Z}}"X`F8E$1!ebKnYg2[CnVEs%1Wp3ss
MqAOe0(gYN-jwLV3@]&y3C6SZXe	Vxnr=_4gk6w>9K7j2DF| q>LpCLejB?$HDqk4p'hZJQs28FcESX4LZYPw;_	UUh/yA,aBz*cQj?cs]`mahE6&]gk&o4"#J|Z"cJ7~_e\7WVB}1*?6Oky:3dsF__4o:8^I~+_$YHr!Rh3.`k&]UncIw?1	rSePl{f|O/[2%kQeQzlCC|WL~O]&>d?f6HhNHYVS
,oYYi5c*P)($lm<'"?K7YHSex(bs~W<a-J+^"B
I^{\3x:@} 7Klo M:n$V0vi06ijehB**P9w5q-YvrB>S*&&1A/-1y~aHZ,vOD5Q&-`j)wNIVwP>W4U 83?Ssbvx]~*2*gR]iUSc
RSN!v@"b84MizNqu",;_m4[?QztPK@xEdN{-Rsq6O(p)"%59h1!l
b>tGd5ppMw2{g--*A(m8v0Wj>B6SKp^(#fDPw&H*xFt>CDiGI},,Y[H7P96f3 F?iSsN
HPX5&X$FWt1F;rCyM	Lmgdg$=8Pa-[R]YEP`Dj0bL]kh4QAuN_<nD4{<SqE7TL=hAQ4x3]7c%=?lZz+	BBbTh4X"az%VE$R*aVMtnl]NdZ&cFM/x.uZ=#b3WNG5i.\JZ/*1n%{,VDE4	2G/Cs#8i1?7k$ySnJni(5IH0C*YN+GK0||)YjT1f<a80D2yoNZPO.~dEVFNm5fe%CYh.(}9GC,jz9;OKFWP*8W&4)^CK~hPbJ\gv8FKoJ$>w:<<8CxPaUaHr'y?%~xus[V$b$?(o"c+`&5(-[@
xdr/!vGx,CER;iRix!)Gqr8Q69Y&aZ8
\=yKLI-_^5$tICPgMTS>Z#)7TK:4|cS5S457v vs633EB	p#XDTn.X.i-!SxY%eSJ.JZ.3Q#/E]	E8QdPmQpD14`[i B>PA8TudAR2Oer|N{ts6LRd>_b1ZL>ob(P;9u&5%I1D6O(1J@Bd*4>7U]"TM]v6k'
c^B~oU
Bhsk/kF7OuLs;VyP=
i?GpEp{0[qlKdR"Z/;+ikBG6,Z|uK^$?t<
t_\b9:qS@Em2G !4\kCwK}5RNu-i4/s W %ajk17k]1`^4CoKk[#/uAr9].4:-e>hdJ'mlr"Egef|2	yd7J]qhoc}[F6,3Q'lFc	t6:g|~VK"MYid;s	NNYI`Veh5+'j~gXy5w:"Zj-t]7T`iH8c^]~eD&K`N/
\J{L"ulK*a<;`X4P`,UA(TbLXYkqhvYrIGvf?*Maq1%qT_Ah""jEtUFp9)x+xtkW'_<r"NAw=mTbOpnIPR@%eXYn03NkA)steZ!SiZ#p)rllB
LV/4-"IyS"O2*iRLxbxY@Fy@~!f2`f:Kvj4"/l->0Rw_d}Y{%YS~Yxn#`N[n4\fBp ('K7N"/K!eLB-eGV^rqRti*	4>=<5E;wkf}1Nixxzo[8'Cw30~oKvBjP=YMg{+lfgU|_lPUm*S!	v3;,Grk/~~m:qkXG0:2mpMu?<krEK9?Ys\	2!:cT3EpUo`Rqg4QvCyGy!:{o,p~S>u6"y|z`PwHajhzAkID_3>v.n%#d`"G~W\fQM;A}wiU$+>-k\;W{xT@qS<>4Su`'.Zb0FlZQD"z&rC^Qw5cn4{aH.x)};oM$m1jloSUl_RFu.V@gkA}	+ \wP}'fIfO4Y%>r%y3QYp<pE
1iasM6mZy|nWjb:%&rRR@%V'r	:lAs"\"~Om}$	cD?2AV5NgD1nmhW6(A(b)r/csK7 P4#{w-K$
JBNj{%gwwW<^6dDI+shX89$.+MkISL^w$l.)\0POrv/+*eA;_[CINynWT@PqKmfoLja7r7k>ep'z6{{m+yvZdn3/1AIc!D^T	Y)KX{^]~0f6iVtj$4@6$xJ,F9d2,MDUsa	^K!RHs?r>y[_c#X$k|;|V{1-\#u9MEzloZctW[!	D[>\2V^;S:f\8#(|<sP&u\7.)cNoJNd02C Y,<$P4Z:*1W]`'4;d d<2*M_f+9GbnM4c5WyA3aC)eH>{/h%P|vlT^O=Sr6~RacC-P2$-tjRfg63$f@Z>p,GS~lUQ5+A]KLJ*TW@!2n7n_}qBs2>g[_WMuwZ3-B@	YKkkW w:<*JSQAq RPrf{/Phv^S\jR(t
mm#U{o_u)!~4Xe
p}Z1A!jlxCZ&	p1M8+B~M
QPN.0
f#hl:h7HT"5b*)'_xjCtf|Kix'544HBd7?']O8BM9O,K+cUw1l"k)lGpI,r#sTi\o$^h))z=Aw=wl\>}X@b}8== 8okytV@{uu7t1A:mc6s7=gZ?
n;oxWuaU|P)_:K^cl~R
'~tCN[7%U&;_7j.[AxDka##6m&o.pw6_D
tEO|r?TmG/]\	Wv=bC]$*!KnOCR*M0Hpmkr3L[U.J{pP8WG`iC5?a;n/[MOnR`q;`5J\L(<Fd\!#)S%tv:r]VB6XCrlGI.^}FG[k]WYE{wi~CdPn76/>!YoUuOe u,(*3r`H*i9dO2Kta4hh\d<ru6ntXe#PKDe=o-

&E13/F	1$EU!LRWfUc6QSh:WTb[k1pAX3^hKxyho+]v]:sqT4&pfqg%&W$\ v'6Q`<Xra?q(b=]ToVL~9+c(CxQl$T7HC0uW`U]|g[} Z(Yz2Zzk@D%=;}	-W<$^Q^fB'88},%,\uC_>30>e}F[`8~>uh%JXs!T25Vo
8:^baEXsUUpB@i)_wO.m=u`k".?DPz&!h(X
dvP4J:[m$,RuR8'zp8ApQSs:n4HjPT*{k59BZg(,'biDjT*5%Yd&x/]IQ%1C"qQN/%*>Asbd;N"+MD7}D}fyp&x	0hi-?yKY^%24g|}2pz_N+y9I)YVX@
)U1k*l5Y<-qn^sWsj{mb.F:W'o/fi%#^N[.VhW?aSB:RPT#u{M{S&<' @P~>OZ7`"JmO
c*O
F\eq[|{W}5CPI>
:M8g2/Bw7GXJ%}>'Y648&rR-&k=$vn4=l[Acj'LWZd"+'6\[}I$L<vH9l$<V{,Wflv>[nBC=LZ[WlZ;-5W-Dk`*uvsq@bP9%ru!Snag!YMa?|[f>DbRqAk(}i7m=D-9dqIz:"4,yprN;pTp
Hvf}Lht 	l	>A_S+@]N-"*!!pn0@\#MYDWDkIg-"OC` (L`p7	LV3CH%}@wc`t2cQ|AK_0sonODew/iDoF|Fv#"uj
Gy7hZQ66<>GzA7u%B8I^@CbO&5_Lm65OFzA,wVNt_g5zEwdW);-n`?b[Z	"''"U7|3J0D13zP*25'7[,l$@8M?4Q6-e)G9b^9HqvIgpSPZ~O
HOM:OAX#:r?ZRc5^&LCiv!y[rV,=Z)rF8]h>'$XcoEw71qs.13W{,q.1.Z<DKXv,^o}%Ku*_i81}vbdrl2#Fm7Ug{@eY
.3~-}Um>0O=TQ#);I?
Su:lWi#"px|EO.'lw9^HbvvNc5A53bW>$ZcX7M>f}3>Qu]^.If[Ph~YqaVg^Z7FRlA4zj&HDQ$D	H`]^-W-U)ia'kS&w{CWc)/b*Af8w_$=#~k.*
d A,pHQ#;#4P+4n@w2oil4="0==|d%M/+8$,zS]D!bkGjcZ14r|Z9	J%f]GGyI8fGr~Re/:1oTQ`>h\NwIBJK0LSJtFu1L[Y[D/<!8PQn`>M.tr=B^fu)}-RxV;4H`S%*qxD^"d%"I"([TbSm>tyb5/TrnzicG~h5IF