[r}:Jy~%{-y'0~ok365XEEcn5lQaO}wG4,cx:D``zQ	s\=]X@^g&8VPc6");9Ye<i;nU.yBj(5#ovZ(Yg{|(bwqLHEWU%uLMxN
Jj
*ry@Jc,fETXJTD./$V,wk&!Mo!'}qSB+}0-H6oRis@3(6C[1Zk|Qri#YNkrI4y"wb@HP}f`i+6Z'-53,{J\{@u%P<V1+DFzvT?Ze:ojn5{3O#_0}Qd.d%]T9id6#"<p:HMY$\\Uw0+H+l-9`&J4Ib;){)* 2O/JB`|Ti'xBAYry=,G>:U<,6*&lkb$C\DC"v^BQ0n5
>Fs\`(~,Tn_]!]a"aZ.?	g`rEqnv1>Ct	cShM4T^Q{K_Q3cbepceqF'&4Plr`dVm
!pb<S|Ngxuj|wTqxop|ScI>vDdM{/:`KvDIJ(?vxBmE1&!HSxMAxJN^FfK7+RN:Af	V# )),pU Yvn2X
c3~6B./nm~BBv9s)@GIGAu8=Ud)ZaAV%DR?Ng_)2bCkphGs#qfzN`60ugJ.gPFy~zSvpR8Sic_5a=Pfbu%=XN*(5ybJC3MS|;huGUVcz?9e5xH.wQ
PSdbl#-"wlzR<Y&F)$?1
{TPx#ENIfOIQ"<6n>-y{;9;Tte_t5E^tiF0YjxrYrCw;kk.y:t1zN`N!ED)B!@2A3=gTe(du6gQ//wL&Ku<EA*e1~BH|=3Bs[T/43/.>)Md&n;/|Y\nY21.j?5r(0\MzSG0@(GELG:Hf?jJ%g;I5@79|;uf'":0:Wh$GF,.Pf]{ Ws+#9Z8U}yGg$*sZbUis#	&=E]%Ba>E|HS[1+D/ft]_v		'7\O3=x:AwDb
}?Q<t.4G387N0K1ye3y4Yjb0eXC 4jby8\w<\ 2<,{EE]J-2_E/Q%S;MIr)IS,.J2 HvG;0X	CZRR<n=&uTYZ(j+Ss7Z^R(+giB=@3n11PY6:@'DYM4VTC*8X1IJ2,HC#{};g\#o5]uiKPZwR;OE+6NnzmMdx$0)Wr2qD#MA)xjc(VpP!O[m;)I]lz[4en5U\J
:}!dwO%wgK6&VLF%8]q&'b"vYlWVFcaNouO]iBWHRJzHW@va}6$5xA`#?U}!eN]n+u?Lq@	B@z'C[8vo'/}ZH9SCUTYRDCO4Ol
hYFSsY8`TcPq$mT(:{%6"JG)<(tv-Mz"f38V:s1j7@PczN~Y{)||FEc3'N.k7"n].3bu+Gv0,O%*-+xYHvW>jqj5;#%trYPFt]"g`IofC@?n[}~oD&FD`8itNoJHi:w-3x:V$3'5z=D5
1LYbkCXJF}}b(R%AqunZA5MI.E&*	""Oc"[MFO3p;_KdQy{a05iQFAs]@*pYm'1InEBL*)#i<'gB
-2')Wj~H6i6$b?`9T$s&>-g@`g;g62#Ehw]"aYT/:b~Yx7&X22QYaDj>!k]kL0m(x|k+}4x{6!wM(cD$1e]I<iAb*t_^IxKRXm.
|x<n|,R,0J@BWGdg7/Rgmkll$'d>]	@+6Z"U&Nzm?b$OKtJs.-0eU,,P.(k#MmW'6Ob;d%o{+y'KYaMna8z{V}0G^,wR+|l|Tbh@=fTFs0Qgs}]e>R\.WC1F Z#q>>CC-L~!6>L6=Ak~HA
XW~%W_>k;le}O8e|ba[sbeorHtx+ih[0J_jT@cbW_)wj~nU`1c\A;i}
|,B2|pS]+g}T!&mb)gmBc4wBXm4y"'pR.28]MN/_j|>sJ<}n>hKGLxMwO1!$^?qu$}16s0jg,{	UQa2Px=6v0mcHZUw,R#sC^	_DZN;NGI?,d?WDz|9srR|'P7U2u;/3Y'rqXA5GE9SoLGP3>3|%>qFoWK	8ia}*3 @1V"*:p.r[@oMfD8$V8S"J>Y_4?;q/*ov3q7R|wz]1a^nre0"PbaO`\[wTGLF|c!Ir	oC`jsESxO^k;L6=KK$6CPE@6Oq`a|GP;l|]"}61[-=R
z[p'{Jc?sZDg1Wr5~\_M%7B
?(teNB\S bpks2oU9)^~ex1-;\m1JQ#<1Tb$d\Y;aq$WUP`6cCXn?"HX!'dP8Zb1a\8t
 |bl5U4[xF.uGC;54]$6S,8tOJJ0nD{)T*= +U? At36<:yg@&SgG#/l~,V%|Q8>w%ty[FvuYo`9,t> ^If>"M7QA+jjpv<E7mp|i>L%	Z8|(wx<2}%&o&G:jsE*n7ThrZ!ue wfIA:iXL<FM{teaH%6LGJtvc> !G#5(A![<4H5Gts
B.~!;Aozw.&6KY&k^@ElgPf{X'@m+C`seS&;&[Z*?7lI+8;AexxZq'RLV
N!TvQv+~A3~
{U" z$d>^wN3vA0RK,Wn,KL>(c+zcRfi#~w8q(gW/K":|Ex4jE/Tglq:-xZR:6(p0run*2YU6d&.b[#9oopt]c3;_XC\->=+d@q2^um\)7a/la.XC8haOQLYohS#c#;O|JLvo
+r9TB|^O	;<]!tBl|jq+Vtc	L*Xj	$Go?K1TV'Kw
XPt0Xz>\iHgO<@XwTbQSy9sy]#VQ.|Dq~pt5tZHYr%/4O=RJ*=`s(+r!0jgWZ;s0>}YG'TjO+n(	37N8zCJjJR^eformg	Ct\e)kz\=`a;
Yn]g7VP7oSU-][}^Dwa\M32[4}U'nYL|Kw[?[vJ&Szsgu\Dg'qE`%PQ_?a6#=?F&^uQ pati1]u'Q&W|I%	G$u9d5xEg"y^;E.,)ybK2MTZ2.})fi0k2frd9C<]E(Uh?Q>}a]Im4"'Y}iDz[*
Qi.2<zk<@e:F(dDFSpxWm,h=-<GGO\0F-pvD5j)%$'3fI9|Y$TVXDn^zL	GJ8\,tuUw"5I.{`)ct2<>5*uif#^Z@/!&*FOe9@o}}Ud8hezfW,-K3oqg&q
CTDnZPs'sJnWh"!<tNqw.'dV[QrjCWa^[k<G;)s^b7RhKaO2F"7PS[+ EQ$U K)B!F6voy+HLZz#&;1yyhG	v,c\d_x8;p>_Ek^93_M4m=Ei4#PR4cE%u&L2@L59;#9$!=c C^\&ea2Sv`'1v:yH|Se!=5F7|]ip>
z$z	o@u2m[;5#$bG(#x-&2ME:W$@sp2H&v4/J$wq\'L!Q6#-hoO3`imZvoTJtm+z^%:OR'?`nf6:<(YBc?6[$&V</(P&s5Ug`TeC
r*lOtB}('z={sj!mA4!%e~<'ZWLX^M0\$I_'U6v.JW=,0~'(Kg";{]=_Z*22h\!u
PP&y(-)eMpfV#T}.[0l"nN%+y;z#E9U9H!5s#%XqDD?x3,P{,><L#/j
r$w`XKOujz{/J9TcOK#{I%|/g>x^P~}X)~Us[m(EU6*37w($-^)P\N"QDex)L(}^-qcyx6vA)\nRC?/,P:I<QiAUqsQeH"1$!xx.
@!V'Mr~]HD_nN$li|f;uox>x@blu=mLKJtwyWeBXs@^&pux|pf7ek^(ZiPw!/%\}YE@DM(r[s`T"=h
N"Qv('Yp:GAH~rp6H5FmZUV=uiY*<EWb1"(p`/aBu,"2PPYO-71pa|xEdl7=#ai;nV5tg^0=_]+$6f2 pY.(;DHb]/^oziln8Blf%Anj|{o^<J&HM^hi{TxsAG}NQ|(+z45=i$={gH4DuI.$q.}o:/3aw^aaLz;58lB<'d=}LlFk>X'H,-6<djb8h?kqOWuY'O|i-C!WATDG4X9SB#pw26W)=

$,X&p[XIw	*5FVyA^_[*:nj{S`%mLL~']@SSm5@&tB)<la4C8F,
(}wktG5x4vBVto}|45Qo^u0f'SnZ4iXg3`JXXkhotl$)
=Ht*3MzOVsdQR(i:Ph;I]|s[-8]'*!s1i8fjcNeFP)VWf^q|>6Le^1dt1]'[/b6eItJrxnSBF&pUo>	DBNM_N'BSB$o7[?@:B"X!\2?Yr"KSp[D!z5/9yT!V	ML]Xlhe1}?5.4Au/52VJUEkwFvk(<Zy_vhD<7UI>\VD+,1&E:2zuGQeN"5!:m?gSTOOOcGTG""h/B\N:Ce716b]%/cz#e5Y$HeR#1^fvW#$FWRf!f!
3{Q$)eK"kKmVEz[o`<y`Uaaka9
I
a[ {>e:;aIgQC4iUW0t[9@EdOuw+o-qwCQq!(-Ts`10qsh*khx}v/%X0`gSwaQMQ5z|x#G,ec5g'l>CB*NY.crnfYqF2jD[#\l	gl-KOzOVd	-o~o!E9Kp[lGEr)4.BWGhMe39#M:0oV7O<aEkcCB\'Yep(5Ek(un#qh^o3=\o-7`?U|_e1ITR$[}|t}8cz#kQ_cBM>`uahS
!CoL%'sY:j^!=^UT>0K-gR@($7'EsT<?n`='-"3xesY}^^j;sb"l"KPr9m&%?|UwTgKoZn#402QV'D9+]=H}s\GcJiJ#9wstfFZ-cV3MowL
I<g5vTBL4O=T|dPSeWyI;!=]}ZOx3lX?Mag/+el"`U'6OzsyA2L*3V>
UqA
k<v]cXEL&you#A4fK(3[ce8v~_#r_/~SG#?>F	mC|)ybaPO&Fy_!agCnRm=?{RqA[fhZ
D&)xz`D.JTz:N)}p!7S\w;e\J}va_Oa>9?Uu,k6R0lo3E45#YrLG>zp5$M#O>1cO~r1N,8l/gm4_UP5HolxQ1y-KD%vZdK`<3|qS&vT	G0|3'|H/.)rO
'Ip?V9(9\wx{~P3P
jGB]GV([X_N\;
nh=)9p5o)9CBY=~q)JToFthe1Nx+|H7X4
jH\%K:W+6}r||`x5d0`n$lg7e#~-6$z	?^$?|ciiFkju:^@eu(/o48*-$ng_zFp0'7.lLP"GP'I%D3(#>C^vI{oRxwFi8&lF\.4vg%=L@"iDLb|?[
m%YCM/md:#]P;e5\=`za%wpC{,ov?nmH?7HF:k[O	R2=]V)HNEWmJXmlyXm#L.RSvaEqU;/=~M-o,SsvZ[@eWxLs7
>[`?3kr&px4H;<y!NV#	Rmk3S-#!kxS!h!RNKuhUtl(K7P2<k[]	dIE4saT7^6?bA!.f#76A|U&z7ER$^3dO4^w/T<S*Br~L:c"=$haiaX.1Hz9I:e%7Ix@S)qjL0hKa{CP7j[0pZ1-Gh:l~jXbS=tPJfMf\X}(QL4`{=ZhA<xV#R>gH?9av,MnW	OG^B6T9ykqSGR$J,\uJPzGG9Z"/^)#TVY
m`kyJ8']ya?*9s[1J[2].(T"	twDUbo#J=a/TL:Mkia}*(B$c~"ItUMv>h	'A:Sj|#YA+<Rci5B!5Yt{>Ng!qMC3|'Pwr)`5\R78Sz}gI
[G:=grnmKN,9<Hm2LF2fr~?xy#N&>`1/-'N<T{0G@X(k
}qJb:Ivw|sog<1d3h>\lOLx2mpk0qmPlH>1FU -xgX}'nD U.@?m:aTIf]%+pm9IuVUuwF|3LpTH'x7D5ib:f/5QV=9`rdv&
<h?_9K`R(|25SySOV5"Y{Jlb;nT|+F&CfrK_r||QL0 ?n	*W;T\1XGVwJ!+tH)Fp+R6q
t{^T".KoIy3=dV|]/onC(ujz:EUPPG\ilx+gL*H2MabdA%Ag5xoUoe'zKE	x48]fX7j J70'^wa!&q
[/{JJKTxOO^Cg(#>x(Vb^/)k5L+Tg\;'VRz:+E{+&Gt)rXZIkl%{knWD_Z heFm>P?QtF	!V6N=+m;f7d}%T~:9I_^ni{)hSHq,j*	Xj=wqFz/-],?pD$8:`Ytb9}Pv^As1};-dkn}+,Z 3:s<dczHobmQ"q(9,_]KWz.j1[#?M{4#3g?7GTx#7=wv=MU1y5pTxO|q=`,0bPiu
{Zv{-'A (uW}VaJ:kGsXBD~yhf5')a%7FOM@d
*+H6T{RmL*'{XL+SGvDs+$Kgj47GrqXxK5Z=0,"
5yde
(C?'<un0sykaZ0X\N<*]p#/G)g:iq_@D#c"7]3$CHw}<Ke
_AK~pP!0n^DwaE
#2-JhqD[Bw-k0#nu+gv@m?@k1 '.Jf0bbG4'"o"h?|:/=WvZ(9#E-==F8ol0L^?j,	QSm8cu=D5m@#x=~8mK~2OJFS\p<{thHCOb9fh0|UEd9 n14|]'R/mS;WXLqhP,wjmeI~b+P7Ww$O!+J\[~>R*S^RIA'w9U;	/wCDy1^Q&w\][r;Y3RWo
0/-%:MpVmr]}C;YZIw9Xg:C>]g{B'*{?Er$jiT&qag
/cT=-/QYgt	0(*lRW/;z
"JI8H@6buCxX}>jHbox"	42EF5_y?%S{vi(^-+Em!*rJT"_q)=-D:.XJ0=t6Mt][8Xwr6.Q,	mj	(73'YLxt8zubNcw"6=Za\:\a2/oV_ee'b&Kn,Knz:l,'x(M0X)Xy-@JC+])w~_URO`3Vo8fB|d.7S
x[T(m3}oUrA!aR%H:k_5#t;y4&G,yBOT&=wO2'dJ@dR2\BauC	WB&d
l*MPLaRVi?@3R^#.u"jCA<^2,X'hh/9j)ebkmnHsc)u2SI8ubcVj?4pUqCE>bUbpj+;->
qX4[G^ 6T6H}XxVWr6,ytse]m$H631X4+NQ)B6MFd_dV5p-LDk1k{\u0XWUIr.ENpKAd+N5l*.(`iYAeZDd\(w8C:B'&g/eAO@i$sYMut9	77E<I-!dc{quPFq -)~8Wty=mJjkTvBxMIG6|n!M}b@2air[q$e%:1xNNy=?Mm5cIbm	k/1&sUP5@i4-8b
(	#
H[#n[rq&cF
(";p|{RbEjlg|*a0Rp$]2m?q+gf5E(W%$&zF=y}Nwf<AC$$HRh{)=;g;P8@m]%k*Cv&'xN|^!(R	j8]= pvG80\AWo91`J92
/['23k
wt~l%0@9X{&?fa"DQ1^xy`0o;G `!W[[;6ijzw189<bE0Rwr`K!npV9VmaUib::b>E"Yz Jq5twi'O.vM*|P@jl
Z0'h8.6=E~rUw)\JPZOcZ[t@n76d{b={mNf$A@_SRBAW-|ng|$&[AR&|zSodU6hdoxW]wKhwt":3Bh@m5	HJ-h^@8`ly}Eb:{j{Z?Ak'MTz/
@fg+zPx8,54,2t|jF*.Pj8Rhh0h`T4}5>$T>SNmurdj_qC}34RtjeXDzf@Ixx\/Ge/PL*#ee3=7,4vOqC\CrAWe!r(0AuB"[aMR(J9RbfI{Hlq\8[
L='ro}=+}N]*pM5[CJ] /Z> 86Jq5Vrd0o=}-QTJ\{p8F\@ME76zj55{AC&BWo(m2U$LEH`k>&X\t<sF2fGRh)pba[}q.:U:gJl|,C[Xih+.$.DX?>1ugUM'bbpY[VA1W;U:zn9YV"5+}>?R&FrKKu]2W#O{hKw"So%((#WbI%3kLa%4wpjH/A,Bh$_	feJV_Cy6T\gjV=$8}!5sqy#+\(EEy6f!v{8"oPD'q[.4K^1w(qtPx
~p2[.Y,8!e/[1b`
ysUJ+F&me%-/k2z"=_I5A'	][)\(M)o.}OZ46jMT+A/#c<===?"8lb18t2Egz?{N({~NSWa|wFm|LWi_pDCR"fM67*@&FSy;~.ptwGi}IHd(<KnvU;@Me}/EPL&":itT,OuG;@ *SCdfZ@6}Gf)_{l<N* X{Y/w{JgA`5Qc=ibB\!"tFbd\`;$"+caIGt=9pf}<N'z@^GK|*2hH3{@*sm/$/du1{N|`G5x;x+u!T<8"w;
R,2q&B|359Q.8/&h=$:#(T8pYW9f0}KCkzY-qnGIZe{}VPW1vjF`o3wnGo1q^#;,;7`i	t&[%BZ::<rFK.gwNO}[KOX'O6s)Be2a=d50p{k)DHWQ&;c-51Vk
Q_G, Be#sP>W~+kR!VPc4'4jGtR[(mA74ZvP]gst<%1YwrU~]9DKFIJ-i=J@#[csMg.X-hXn'$2G;Rc/`^0$*=E\wne]'XU'(l/[&M*a	.*6gc<$gB4o3c1lAj~d :s^R0'
^lXg-KCu-'G$>apaMU6ko}g%suK>_E
.7gax\$m"v55>4(R".~AgL	effj$jL#]QKX^ Zp:"'MX[*		6@V39cB#j4	JYampO<(n1;55\5M8\~4G2mvB=N31mg{:_rifPk9-%5Xh,TN
GspBr2% gKxz9jaFcuWA\F['HIIi1tF*We|NRiND{j
JBJ=.+2oGa3,F=czxPx-$o|lMa>dAcT;6:i~*:O^XVm8f;^FW?j+Z_k|#0N`bl+Lyg]n_`!qeJcbOUElXH4&'7%<tvHA#k/ee*x7*~2!d=l 	EW1~oo"U%39p~kg{2N$'R+ug!\%vD~=9kKO!bR,MgH03J	l~$kYCe*a7e-_q?p|E=jntH&T3^n: v?PufU7A8LrC: 5SNp>?s:mNRP-VevN=]"V#wmag?5%UXvTSNHKbB5g?bYxestA<dnd=MLS[|ye)L2?{2xL\Sxnu	FC
Tc_)CDDT:Z!nekSQ=%aZAwbF8L&^N5_sTZtJT`|T&c'E%/H^`:A+N3AB)-j<oCt16z1,)w@kGhw6Gu93nyDR|2c<TiQj1Q3T,4l^+7\I
;jd{),8oR
3+}+1*-[n{";'8UJsp;P	E])/8|`W*Fw1\0+x-%zIp~knVUYy3O9lIO9N^fQ*@m1e R4/!w./7~Jb~&#XSRH,VsER[*FwEjR?L)~5U*t(gM!/>^	Ck:R+{*3X,Y^Po; Ov]h6R3`M#]OuFrQaa("AF.#$xGp-jwe7A/gc	V0rmso>fs@x8)7BC_:fSs&kV(	mS K_G<`4z.koL17ItJt7X^`Wu'JH:'n+{^#Q%fS<)J{QpI^zh$]dZt*[@zltF.0Z>'x%~kbU<]<qI}>fJ5>|B4"y,n}MwjQs}8{[N9?
	)o3;hy=VqLugEpkB R\t.ts]Ma.tdP:5"F<-[cAIg&I bp0s=D_9jV
|vno+Zs$lneao@Q0) ;bQ;%jlrW E^spP,-hg
^?uF[cCc3jLV}%`8~`DNhf;iE,\#!!ncb):VN]-F(};g^8<(!RH,-CCuI\#TW--yY\0<|is_<At8n=)lO%<HDr`;.+l09o1zl7$ig8A7z:|[pyE'z=(cM%z Bx@ww9Uc=$\}Arxv>Eij3\cduia_Ldyg,lVS-e#\Tw6*_*X**sz;<yn[M@,abgJcG@wp) 5=:b7f(P?+ucB+fa.ydkj^q2B4GiX4wO$Hc=mKcQd}HLk~Zd;qe}Y??mq#t3-gGX8(^3_^'5l3T%d~wTA%n_!'C1;[4jG mQ#=/q})1i;>7(_yqQRP;X|
TqID1-q(RP%-?/F<{?pPEUB/Y_NWos:$MG X#4M^MoyTUjQfN.M#Z:KI M1Ao%Wlpx}4u/-`<WPwb%_fkurUx\-Eh;L$9XttS?@cBL$m71F@B!:&+^33`#
I=5SvW==[]X
f)O
}Xn|
*J\"WKLI)lL90t5LT'FX7p[,<>n_]2]0{v7">Ej^)qw}rgO7pu[P.:Mg|-QL@61Q%?=T2TB_*N#-%}gTn}#3uJ7}k{X}5Fko~EQg.`Oe
=env<8	
'RAD^3~G&h$Vzi}ZeIx;<{{{*rM>PY.PQEN1)T	9'zNr w@/D\&BxM~9VDc9,aEe>!{#AH/]g0I}m\\	{_!pycc?_IB`F.tuHXD:!0.,b\_!`|_A[
C}6W4taty'"8;)MTv{['*Sx=+3EK[-"!j[=:6+
CxW2"QpgDSFKW&1JW)+srD}OgZPUh;(n'>f,MXp-szp?ca4;nxF_A*]<m$%Ww"tG=uL[DR^>0.#ByPid5|4G7=5o8\[%]F/Qbd'Vs'"I8`YW]Yxo<dn4T#r27_JzZarN>-K:M,-!]VUJC!P7wo&@*y' p~#,P
aW#Uc%6P~/@DxL5BsFF%h[;|V.IG_m6>gi{|d0,Mc\D|FbI?d%<^"^G^sn/`PI`XC3y|4Jq	+GrPfb*)SNna"!li9j^Gv|c|XIL_a,9
Y>{`#8) ZZ1:B##H{zqD0.>X!PKc\|";5{6#<21ix{=`i`q8SCl;LCwR%86Z&k-{,3x5cdm
P!gBHExQ~{xdL\oI&~=q!g\ZXd~4*CRnqH!73Nhp,.B("@m?<o96:&7	>vFk7ysu30nRur	@'4[GEWD[7a(],jBF1nwf~'BI
0Qo_Zf`BfqU:1Uh(dW1vJ1^g|{)lCDfqj_	n<,x?C4WFg#NmHT-[/W\ehCC8Gy+?.2VEf^b|imOoE,:Ns#u3l{,w-o>WK
l{xYy?jP2k]@7laVeBD)HSrLJ1|NA<J673\kFBF-K0g^j=j.#N+pEw^\6X.[y21O	z1|[F/sOD	efe9J(b0G01B Aq,J<Y2$T5IB
e'R#pajX}vlXbn#Z	4[<6eK%i&|W-owOUyZn ~VO1R]nm_E?#X;&8z>=R6rBsm+L/1kJ-
mk^Y:8s83rkw6V <:*ZsCCwvR@#|ux1%{t6Oa+	U9o'w&M'dH+P9]]q"iO~vEX<4I0P__OR2_S^C`bMD?b'SQX|A	JkDg
mNZ
Xzbq6R]^ Wk,@D<G!Vb*noBDZ\c-&^?-)j+.dU7"7.ZhG{wAcBHq-C\mc)IsriG&	.YOiT6~
,O
qp%V0s$QQ(H$pH?0TZSeaCkT[7YG kt:clH%A
R%ER?RZqUFP?DblXuwK9~zY1=Y^FeR0gt,o|$!iGx\qC%1+LN\4ZuR%'_wfu)`5	Ap;G B"'pOq7:0 9a&9WO[oT
hFe>[3'TFcYkQpjY]mwt#joeF.wstm:,1D2i?EcF*M{OR/XIoSyxkz&/ZYS2jjf?]>a?%AtJUOOlNI(EE}*[TryB|m5c#t^\xtEm.EZfk;6f1ziJW_Dt*jf!_ S@B&m]-Pr/Bg'p2A.2Jn`lpcyA/_j%G$J_2Tv%DP"_AR\A0V5R]Uw'j..4}oxPZXjf 5AQbwRREM9Dxx8.?+Z-m%,MuKYOVf|-xc=p}E]p`KG=J2pikU7JY5p]331
.P`&`E^	a-jct_%fwv\m3Y(PERzzo=yF(V#mH*<	M5O:\wA+~g_%9eX'ehX+ryN
	lrbt*HF25b&BjdCgqpP`^:2!xi_4T,V(K#)8+xvaSm&o\sp[89.vvMX+ZW;6gdw#,}<wf1nL9R:n%`+D0Xf$sh?11VSA=FGdMYN5d
$/@!z9`|_q^*9yN D8uO;cx}]_ZSMblWD<y".!7P/{cX<Q%MT	hUjo;]0-D"8s!XtC-?>XJu;EL$s^@,t+G*5
K_b6t4fCKXSz-qXnhfE9W:nKTU/Gz4\3-;\U:r~&7Z:=KT":F*deLNe
)aAYXkr-^$[U:0;Ag~s#B0opqyNIQ.pk-0*z647B3f8*T}&0'<m(>qK0|eW1U}lu}#Jg]=<J vR:Q:^%*3M1ZEpE&0M}uW=>C3r;7x5uR*jUWG W_8B,b,/tDsZo(,]*\)7i?NLr~oJ|vN|f^]"/,BZd5mEPcy$b\
?J+av_IThn.Ra1?LW\FG][A.2oHpz[(R/E3^,Jr$GV~H7U93kH@|oc6+-,!U+ t%o8KJ]dh!o?2*Q"2IpbI$hT\^eA#[;6&{~4D-if
V5:g
-TyI? j(2q(taP/X-H0#WS| \"A}oL:	NcfIPDM.z{WSyw(PoF#*81O.3%p"4iq5Ncq1`<;W'?Y_i$N9WE1oN1Q^HH&#,m(`U5XS;bIWT>8mn]:Q&X]*oN/3uO>=.owyGO7uO(h$3=	HV8t\!a.C1`&;Ha:_9,2#CLL(BD;5ow='>?>;BG%UMn1Qu-~fy"Of,cT,Ule E*B@-<QcsY5A88g}Q.#ZP*H7+PaImp`]"wbHQ1xEup<BA|E*KVOLJh1g;hRPOcif2\G9BCU#7	k!#"~X&:`M%6ZmaV"rm0wc	*AEFK@UtOB5`zVG6Q#%B%uy"HGTOJPIYK0'G~D.9p\RCK8D.P}}PE2U\Qh([h2!?[}D`h%)32Z`.iS::bn=MfeC%y!1Y=TF8
Q7OHQL)~Z4]^'V}EU2|'mU9.WWeki.RInXrjNOq{f{mC9{t=\Uvh@)(_iX@LB(K>M-/iEmg}?, 'es@S/B'gmRC\_{w d+?sb}Sexg[>s&Yeic:G$.t3t
|dhb\C:JqGOr(RhU)ij1+*VSX
vlBkNFM$rzNkW^b*-9Ph^%O>CN/fx3Mc)WGV%
1>^M
aHkSoQ%1qhB:%,y3B*)	t(Fn ~a]l#LS9,o?7&5 
c>MNllf[v=h&j}]H:y*^.)4^ki-]l<a_',,"3a\rQ|ik5Pf	-\t'no+zO>#>Gq]s<T_7Jzn-\j(2R[^gT>D	TD;;6Z"oo|o:|0er)S7g+B%T *[kv9-J!+ER<(n2Tqy1a{p?	O(,%]x,)__4c	_?ik@}M<>HnZmCo[NIoHsa]R_:Q*g]1*t&{ThZB!L&3(L1VS'U9@i%4<3g9h!rd_Ng|zW^F"Jf:=(s-vc5j;Z|T#L|mH\i370vPsp%&1vYI.n'_ZwJ7?myvqd=v*+i^rN.U-%gv@	SL!AD*5Eb|^kRY0U:u;::Z&Yru)3n`0RK|x>AdJV;z'V3X!=]=#P"u}G=5jCZ0!GO7{AC$JC:G?TxqPAN2V/7t$Pd ikJBhrk3ya_M\ \N)3j+bw09eVueOzF:hhGJYYb"4@7IFQTs[44a2mEQ%C [PL;&0:4T42%myDIlF68oxZ7|aTA3xHXWQZwJu^QNm;E+c\=.,vPi$*Psn7/sd`>
"Sq~\L[7&0lu
B6q^761(#jF4Z+K2Xuyvh|!&tlBS6(aV&z]c9a-J\Bd	3`@egR#qK38	 szQz7?GW&\/qBv66(?DqX	1gipE|[thE	Y{k4"&	3-	m^rs+sKt3%2en!)jc3!Yy9J"z?
5sdR{Czf'B^>YAKtfz~iml:8cO$@oeU3^wv.}"?4QWW8W_7O#\J93(pNkS7CLupdfYDmh3=N:UwyK[2+r-D-hP-n$D;t'}1tp[a<Y\.<Z)D&dW\yc@I3-tMA	>i}qZ~f;'>3SJVlZOM%9}u(oVf"wh|['-MBgHe6[b"8'@m\VhB@"=!2"{Kk}zkg%6WO[#6dG_ 0
hsggMXFE	sV^`hl8h	fbO{Ea|^OtJX=",jHP!W61TzrZpw?Tm(JkOC/	!0MicS\p4G:\v+oVyuIUZ't)X%
n-S^_B<fL!H3|A%U6L#?}^ql*ghQ0#l4
GWwWcz~)2rmRYo<A*I@!"X	Q9|f%>vuMO>/yW}`ZC6@46P-0clmOhpj.J
q]!-2<"]t }}YoCmW"V-k\p865ULx|z?LO3\}v;ILtG5s#j^x#.2=x(Jb:vGk#?-jx(M$g;i..l'Cl0Ww7Y6)%0Lf|f+-wJ)fvHvIWruR$FoN:tRy%[`%XLLA'	DgLPfjGCT|"$oP3j~d-0FcVl`w&gtei5V!5cHIde$m2g-S:1Qq2*;$G]RFAbW[Me2]t'r)6}6 mJ*mYbGwPDa>\;Rmk,RE^[[|BRIE]gA#<Mwd0uWTb}4>hFu\md'?:x]:_gspd\6(6e>h	mct{m32?|{(Ht}WaTqNH[!xojkSFl}/"_h ivh7=e<$Ta>=j"[&8r{G&tg;pyueOHdL}PA@F.Le8&d_3^}DGH)zmF/Dw
Q7J+iSdG%CYi9r@|RD|_7N-YQNd4e|><FZ,h'23),)%}3"=FIK6Z7d
.y]83"@O:oX`B%wQ,.Ksexkbi$?npSrA<F}-Tg8]<RAv!DDBK?;GO`#SGq$Y2cAaCjFm<oseMM]?7xA<@V?%x7RX?Vw8&pl|=vDA^GT-M{OJ>33>K}_f?oX2sT]5)LkO@GqzYW|t,O2S(TU[]yt;+]I	`K.>4y;qM~JM}eHWRW#D
Lu&:8L[<O)Er!;bo*UHF(7uM?^;`f1Z]D+!Z6/HzRN":HN	WB;6}{1b#CH"$s8EaNq(E%qQHuxlx'[w2|Z$p2}	[(y(<p{)f&Tnztb^(57hsSyPR<^f[5Q@yH3zYVvG?C5;f?`<^p#M0E
:%>!{Qdz&E&S1M#AgvvxT8#PeG,gpYB|EMDq^r|%5}BUo4)u}8F]0x@yt^E	<L=N)\l6JE)o.Rh:kQF,vY#?)2.:kz&*dM%@Nd[e}bE=d<'^Fon<z-Y:p/?FDP 9lD|E<FX!%9HOj&[*Mw"1VT9$^0?w&#$ppjLjyiyCU~LukT:pB_c	z$)@9y0htQcF
[3l
22}r0`O	TyB2[2% nNHVu&=Ve	v_GM>	Ux<a2`z6w8<;UGA`s'Q\>g]i6@_ ].p^,eOw@wlIs^0|qtK1EF:u"xOqtq:/kD7Vtv#6KHymx!4:(NY;4\di6H6a^LkX!3af\T9,]io_*\3