h,="xhsYU%Ag3o2vHQkfS-a}$g.JSawV`,c;j8%d/2$:\z-?u^agUFZPjd%j#"%m!U*$V3pAV7gS<;)
q(<$P)"BAePgv)Flt6-mUfDB]04oX@Va
19anSV<TJGb}~l"cMA{.l:cN}G_8F/tgx=rao|K}uW+#fyW'`GIu^2WorUrk&CX<Xn<?%A)8ct`cYNLwTzEflLY"^TCp}XfPXWZZ`pG1=y"Z6Fv,3}y'Clnm.G(	g1zBdYrdS:Gh	U	SgkT7}9/I/.2-Hi#uwrh$nM5~'QBoJg{OwnBz,CXG2J{7nU5~fSX]ojP)Te?y+'ogpIs&==_QUaUSTP:iuk%Cu-NzzAq23vWZ\4LcmQ2;LL`e?Qn6\#-'??CZy8|\1%|T <!AKm>#$JXZ?QE`-i:1GP[ ,*ZF7qKyO(M*SQo}F9hOBq{z#3HYKxM5VoXwQtQ|^<;jN@]E#=~F.=	~:k3(VVNa6i8(Vdc,p	K_'q;FF$b?	K1'@U0-@ahd3KUI9 [Yt@befHT<V7z#1~,j(AuGe<dSCz3bxG#`fq#J^f_a#A9eK`l|bm/4B*S(YfHjwS,J<w#M="m/8hcSq+uA%SHE;'`<ez*cviSs^98*@y!CU=tK?N'{im8#^:d ;0^"Q|(\#UJ"b+~MX
3r
^mv<u0UybY`:N8WHgF-voUuX]0f>%!{JiVj$#n;5\5Ie'XO
)Hbb	9PG:C;Vn>lTVRF1fTRYc>](&-+.>a
';Z%A:oNh9DV'l#.(//@d_vQKvP?E;{K%H'F3ek*l+&eUVnBfoMb2L#I}NjiE9\	bFJ=&"Zh_=*-"RUdZ{z(7l$XmXGPvbP572^/>\JWjv=J?e]0n@gc:gF`sh~7^@1-IHtPf l_0KVxo4do3?\}tl-|k8'_O;X9Az/g4c(<:yaJ'6{|GuEZjjlc(i}82<9ms/ZXlY}Xos'g^pHZqXVM(,g;h&)^_j6t^d#t=n12Q<1:U`&Ok5La^z~L7/@y<?xZLpxOh2h#4Rpna5ERm[i]:Pk=/fRXi<}xn<[(V>6o`$1h|]g}z;	<sYzmggNYs.iU"ml7;+iuo	`{&u"Vt1g]W]=5f%]%<c3h<lwwQ{lp2Q#sZ3uXP/n+heU4"<)<_:]a	84%9lrUre%qu<Y&h@3%cKJZ4R:IU2m
o&+f5@_U:8rVu'$Kn#2>NY1)6 Ad|H7>*7F6l5mU.GY8Vr*taw3Qk6p3^hoNcgxQy2:l<1r:/ai=(e:i GC3AgU#d<E$NaR	D_jVMP5)qZ{y/HbzvhN',mC^Uzcbc>$ny=Z-KJeRj!Ms[K}[OK+arD0r&&Ya%l~b3=0fL!v@CjkI*u25Y?;@R*@XO(ML=}GaUB:LBpVP`iys:3'2	F;!HzCxL2.*y5Xrzlv-++p@/~YtI8rpNE9|*cs?@VsNV8PQHqG}mn?<t7@<?[H#B1(ZWEl03s`+Ut').Q|v;C>UK"U.gEFBRz-]Y!26j%&`N(O=tv`j#DIHt+U/OhQu["WF3D2F`uY,B:+.l`63KY6.jOW)aJxE
e&w0 )j[cUP[DG;Uj9E`fC?Ubq5XxOWS(Ph4Yn8'MQ[JD{;r*'p
M%K*)KuXSm+uw]'OLc'S0'455O*:3n{-w,F]:<.!6G`}Kc'cftJ|dcbVx/%
^]f_^m>kN9qgZ_e$*C9D%2ga>
]c6FqJ[8dx+E{8m<}8`{QaqS1urNy~/oS`L$L
3.p*]!c4/DHz_ml-;~$rwj'j,sDn-,F%p/k7.ASG IDXp5!g&aw\`(P=t\G8ire&UnK]h9nbo)x_W8S5p"`}TK_bHi}Y%!EN4rp<iNTK3pd:lA}"K.2Ii6"<EL]?kN}5]f}kI_K\i$u>x=V=7~x!2{;l:B*)lDmKJn/]_4a77s(O::#Q|$"Z+[>wr;_?{S;Yi]gpC`	U\cm(
UqqzO8O0{}MIh~q6{?B!2T68WZDTF1Nu5-(H<Hr@0?RxRu.R];G|4g=0]D,z{U"qz%`bm=C-kGh,{?V=JBCt&j318.m2:Z	Ep%L9"Od8r|};(f)uj>E5w<wCL>:jcxJBianIYsv2}w+HhA9V~*'ba8j<<Cv|&{%G($}Ob/|8oZxfK<L1{ rWv8kL{JS<
vz\9$>#??-CeB
b6cpBla<QX8<$?Fxe2Q9h2D@R*V3dPC#10R-w{fYm*BR<N/['XZRx49z,^|{,nU(QK8g7aEz@8Oc<!Jy0P.:d(nIM1LQO/fDPJ< E,^,0%;m3}hwSFXzpEKr-A(iVks&)o,[qru cl5CzwqDNp9>Kx130ALCmg <wyoPa'Pc1=Epo$l~Sgv#jyn^MmIc? ^)W`	1QPPdW0NCg|o]B-VjEV*Fp@*RJvZf(_Eg
a;l}th6 AJ:|Gu>TYX'A}g u)IN6^$e?LPimO/oV,|0]#QH,w\nhww(/^,yCnu2:O*U>E' Vu#
H-h8ummAbzqc(rts:h@-3J^(mMu'oNUeNNg-nx1WlmX2bIw%!,q"*?+")GWZt_T\@W%&/_bLNdM)YWM{MT4)!p2"K7{>9|Tr@443)^D1nsK?'[6d_b5y6x-.e!gqWV7!<|gwPbP?w81BHw
J&h6<4MF|`jaBQ'"Uv<+42+\b4)[G4E9(ceymWr$)SNR&-:ooe\7Qw<&`l=9Ix]VW]aeWrYD`@DY;VM"Oe3[}Tcw$a%RDcyx_,CC{&dQOQ:H*8O0	(hBom.r3CaG?2+#S"C>KwWof8/G+0^2,lnd9YY0Y\H_d\s.tQj;on>YG1K8G[NHyW3H?7h".0<WTYR+Q

Oj'%u!CM'!~b) n/bbj{C{EIS[acl\;f
J:$Y-*sMv=5yG3A&'Gl$*!%JqLfFB)s>;FKiEZKT/Bj%cyX(w`_k)NK>&>{(dqcBa;]2*E#>(l ?:ETi#@4e<\ZT8+jD,bX]_`F5:5HsuL,s'p^"	H=:oXHIat1w!l&_2Smgx=a!Z[)wo#;|@Q5+AzAcs:JD(!{c1zDC&Y<fLV*
L%dk0=t"c=>9Frrgvv@m+eGD*LgletB6T3uT5/P#:awiGX"|/jnRud}.N	x3hxd`kp0KOTSo8F8]60`+1Mrs&QmvCyvLW G	`Ps5Vfoi;l.oiQ*53zf<@U}`u33/{xo_d[TFm%3KS^N<)m
z,U%bst'jZCI@+n{9gDa#FDX3K&Ji1lzJYV:*.I?]*gKm GH.~NY	GkaDu(%|&pL^2
QP+!
3IHWM3F>(8^Q\*g3J7-RNz(}+q4NyX3<D 3g-8LfZp&T#f=[ s}v@nq7wxx\fOsOIaKaA4lJj2:Kip=w\t^nrh^N69v[^A<I0gpSaTn~_Ub+I_[Mh VW95j_+O]gmaTC.+3;bTnRE
0~5`.5_4y\70tgD<tsFz|(k)y_nQC=T.Y_%&GF/V|Xj#Of_hNH,nTINW]+-GKkMsb[tPL|2$^UOz*fFYB]EhzK5X3_4+-AV<pDGEI:F||E~jyP@$pUVx-W]-qIX%X39a!dvo\PvKA?2H"@_d]c&im{lER?#^"<A;~S*o2_cyfuGpF?XMu7Lj4BH&%>(*MDn./
2!59GkQCO1>!*otVKAVB16, :#-dm-5}E0E~w/u!Js0gcy]Y '<R?m+.F>B?	Zjgq]Y.}mr"JB8s++yD8SxWx]o{`tad&.V_`R#|q<3<fh]BZugQ+D@GbSuh
uSkOG]6c_/`o^|'SE3JR/TD(pekU)TU8I[0{"$[L(LQ`x[(p.iBm5~WpRmc?&am*!}D_r~'V!f@1As|0#/W8(OZ={_xSS}P^Fnl]-]q2>Iyya{@2J#joMW(PY?MiJ?VaY3,|vI<cxd$=;!#p<%/OJli\(	eP'N}=(0,'VciuEp5=No/$XyaNS-7ZeZ3z[rJMwt/m7JSD3Zun})M=C{r~$ZUKfIrT=	N`)WgsT2AoarzD%`J~\-<F%#9 =C+d TF,>w|2Nz*wW"Hi+yv_ *7sH-%t?%QnZRTl6jD2&-j%?=F]|eW6^vBwQ,(Pb/_DM[o>*!	v%@;]q8"7~;qjZE2C^(i|%<r>g\0b|u;(3aBh&zxB,aN vbWF]tiG@J2^`)]>l9/w1LwBy
KYAAnej[HE"7r7fgt;
Izrjn^7V1P]dT!ZlosU_T1	tc==YIg},q]kLz";LCtwdQ|$p__W$o[?tc<;8nGC"f+1cB'$L<xr[cP:r+J-!'K.)[Jn>'<M)(.0I0Dqw#P}KbpB|]zthf]Zb^xd`wnJBGu/Kh`F"@MW;$^iEUAHcRL,#N{1|am~l\_Nkusn$yMIDz(ajmI+&UF|}Q}ESpSwX(1?8Tw&U~`
C]W]Y.62Tqm&'duC99b2gsw\!#VYOdVNeOWNSqz#CJe_-^ls0"&Vq6 Rr<0\k@:a<]Z#4WFHF7_EBtAF&Dk:m_=#0m#5zY35V[R(%D0Fe3'jxM_4x&)rbSX]rW~MP3!lPfg_to',e]3+-he}>q9^2B;Qml5qNL(cMeE4rOXjD.MHfU|l7<FLR#U}{i0MPU)>Yb{&>M'(VPfm}va3LUbmVHu'cF)wt!(oaOudJ2fdQ!~,^s8)yZ*f>Cs7cN$aT3Z-\[C)aR++6-i{Db/G_IR`:-b{;nRz7{lugjYy;^sC~/^JB_02>]\%/w_2X&%^;,[h)D'/~op%&%qeu n{/	=Wtcb~]QDD~Pi_*|"Q2t,a5tSXRmo[x~{U"*gDh~'>5Zq'$FHn':D!T@@vjx&tJ_lGFm#mos=k83>2-f*#2whi?g>i]+sBb_kA\rc;k..rP0ORUyL)*.(gA/3=(Gh|wS"%.g?rJA81=GNPy;(B[j3uT7F+)/6kZ@X{%{+w3|*Yev-4H.dF]w/%oT,p3'Z("ifaG[qpe[ZS{Xp9BZDa7hU;uOXC*.wYRS/kcY>k?d#uxC{=X:.4Qj)>[dDYS6?VdKR#\fwA46ZNk43~FjGE>_`ls"\MqOh%rh<I7!@)BEioP$YD"kAs|sKTd='+Wl'i(}0kA&g|6(]?}#M{;60WN}:"=.~_G#>c5o\E,ri!e%)*PYRCeHi5z^AkMxq?L=ntv_wz[[|RP}2yS05>pd!r0Tlq=k{Xep~Ga9&eC9;/(R?fN_]<lR7`~oP^&;G51M[Q&n5$?;w^yU?CWt#!8zGs+<VM)Vl=Sc)lKG'`#Vc[#|OO%M5~Pr^g'^m&[RJ+Jq3Zd&Jp/`x~D9	BSL;gdHfi|n-Sc;P`y8B/E|fJ
!>D@:>FwGn-VSw@J&T; Dj,HI{X>VpZn'jv]&L+-iSk/yTjOe!3QW^W3b)Rme	Gc/j!g!I&~26{OA5)P|+<l:JCm]1q/Y%\p-/zL= <u|9P:1.)/PYsD|*) f6d*{D|qjPG~t`c2sh?O~z3|+RFCfper x1(f|JA'l:)cWN>xPs@,wPKeQ8o~*QUc9YK[jjp<hB{T.qNF*>p}~0[zq/VINj@SPB:'E0lfI 3o4Wy[k$t]=D0C9u0Pa:kocv<*Yf~Ao)EPhG)eI;N	m6GGe4]#	_\58-oLNAJ3g:a|t=A,EyP!'OOXd/`OaDz5]qzO@aWrBRzt[\r}"
Yj<U3.[%c=LNgsM0QWu|l_X(*s;<NCgU&5$G8uh~QO3v}&gZBR?SF5>8u;{CMhD%jMo(/R5DL*9kI"*7a|.mIJvyE><@UNM}#M%FCofW7C{dAhRpR"nrKt+ol{[_Q*lKl:"P 2YX|t;Ed<rM>^~j->;ak#8hl
Dq9sr4\w|!0X(x1_	q`j-7t+c8YqsFi0j#r}}7XPP~+|.	Pwin'3qB/%iu9*u]yz"qVUTf[fvL#h`kdAfu-GEB]\Z	I,Bv8Fg	&rOze#"k8WtkV|&p1/	*p6-l2}/g@S?l?EOXSJn$FRO~x,2ee+R&z9v;^bbxw<[b$Y@]jt9w4}"lhbWIuB&9?K5PQ]AB
|M$8
lx
U |>Jq96N 0k9i]!u:(`.X>R	=]-O._%x[YoJTmW:H;LvVBij/-xWqe)n']*3KVs^|@TJf#FV;W<{|
R{`\y6s:B[!DI7URH7W&FWq$X9'z5foh2iYEOGRY+bMK?P{	a~~h/.0uD:A/h0i2+Y4?HCI'E'p*p|RJg6HMdl0y!w6Wa;	fq{=^G#h$l%j7-/]T$[=Z%b2=^y.vSaBx#A 6/W`2jl^FZKrW#\O
P=v,;*CZ.	rwyYAa=]l@3kIK;\}Cw Lt^s+)29&iuXZqb(BDOr2I-3*7sbGR\2#\8<gfjppDCZ/dfLlXH)yC5-
s>Txz:+FZQJS3Ez"e||JC>gm<`Z{nSajI.Rl.}c_@W44/v.Xu<<+	mTs	@++BTc{~]8g*W.10o^3kFPlqh
2y>CYF[?^!#9_e[8`zyr%B(Jaz!Atb@kkD}]%|?{{8A8,EtM4W0Xbfz7:(N8'ZB-RZ#hDt."nRba/Bhv|b^PUW<)qFht68`)	G095%|-c{|fk7/(=p42[|3\QA.=+iu1,V:w}AdAx|DhmxJ{rf^
?X]"RgV2y#PxWr]}I8<=rT2co5A>`Q*C7g`?S"gY8sJ)aZFa{cYi>h45}NZw5X%iGY=so2j%"VQQn|'tHv FinSR9
>5,}kws(	zh!.?o*MZq2sv"[XaQ@e2725Pm/YN0 LH$ MQtJe.dk-9,:4]7L
V8$u?m6n1eZ/HbmV
V@G:CR*GisH)Vc[%7Hz
NZCtZ]?B:TC ;(QDhx-.c:7xB|U"|H{7Q?nM}	MQ%+R7f2`l&;ejkb$"Yg+Z!(g(zwH`M!+'d_\I#0.S(Tm_*U5owJ0o[kQS>+FjxKIhy:Dj{b'nhu;di<?"#voYzjO7`j_XCFdLk0saVpQ+p({3#CXMsQ.pScyYf$
bqgg!p3T.@#!5
A4lf&p>rKF+7y\,5(@9KS;=nek2{SAuyDG(c +-i5+;rij(-aL#6Yr6mN{Ke@[{/E'd1u.>C0Jj1L'xa1aZ[7vl7mfJhe_v]@#6B^7g tV6`OqjlEGzo`.OQ:~}_X)sk-K@&$PkFbFD6e*Ge)s`.]^!Tw>$S
d0>N9lyIM)yCjFq+<C8ZI5Kd.qR(s ZUv1_iv@_/<V:	J2P]5k5 6q'_h85Qq4r&E`5.=X*FD /3`}&&b:H*	@_Ys{LOS1`j{Zjg^i: 2:L+~!Is{L3@(wV%=Zm8p!xj![X_S&pT[CZdo<,[|DT]Z"APfMk7b;ZN:)XsfMEOKk"`IMTw5]K"}-d:>zf.7x;;CZ*Lz=>	IN<{4ex:Ln)7`DE1kc,21h.O!rwxl}7\cXx*,&8iYTxt0hv%2lD(kgk$y/;jC'LnEd:[$,~D?P:IXi`;o{-qF?Nh rd|T*&S<Z55q].Q5[\?r(S+6s0U/$9/KvWH#$+#B(88K!Wfd4}]{w_M-c,cEyb\mTg$-=<'myk#pex'4R;iIBg%[2oXZJdC8`8n4XsDYzZ!XL]_O|(t->u-PftP_($Uho%N*Z}q]V'*i(	=O,D4=$[=;0m3DA(Otuf@8(Da	Du_.{bA\&7`n#f|kHB'FLDVQwrM%EU!NEiC6Lb~%lZaG0#
 h	OYn#,@F2E"JxT*Pw?l@5B	kemeMVSYDbVlK{K:b]tMYL	Tc,NB4Kv2>B-RL+*D@gpD*e~Cq~|u}cTDNkFv=IU"x40dhkDRYQeJ]-hS[t`Prd"8?9sM6UbJ&a$ET)!]	 E0d;uQ ^pG/
qO)OBN0G_<!QdY#`_AL/5 -t]+g9;81:^H!xQ-%6&;%WklHLYnDM_W=G6$8}~s%O&a!)>\RW7wv9kbz+rF%p.n$"pa  2~saEz;	<,$4%rSC.JX9N=	Iq3@A0{Hk$Qi].UUQL!S+^BpjNph^n6U+m'?%*f.InCX7Lc7hm=;!drC2\\cpp;9\5l*w\X?_W;*<+M@!?nom@4<9.=<|4M'/iQdh)m8-/YdClFWDD@Ef]_q:i1]{0M

c$'@iL[ZHFHhv;iX>,T
WX2g$Js'P9P5k|"HN_.3;QMI#*>Efr%(b=gyra}VA&{>WAQ&MAc=5oxpV]$do_wqPoX?yHUxE*9bMm>:`D9m:Kd&sf4@dE`7N-.ut$v&uD]p5ps2-ae5ltCwDNC$[=TOwC,it!BhNwaG&(+\\F0[Jg4Oq@9.k}]Ud'"/dMB:U%8)#/T&{G.[s	25DF?|X:>20bC/|@@#4#*lGDTvWH3zfTk=kvW7)k!h]y,HPbDnm,T/V.r0X'r`gq=gEt|n1xC={JxzK@f);f{Kue{eFj@uV(Q}Lsnt\Osl\Ud&<>!=r2m{#YsgZK&y^%7-+`2H): .~1Rl/%59@0fO*z6mip(o[=>0NlRdPXG=YTI7tC[I[GE>0GlLm^!)`90\7^|b)iLxP<9fBm))&Dn\Si6"5"d$Wb
Q,HP\cun3h=^]LDhUTU/hxK%a,+#9I^])5)G?
 `3T>`+.JTyo9E%TWw\OVeTH^p`r2i8v4fh-a!82MsLVN&X,sjP4AGRBtQUIHj*c\-{c6Z'Pch:v'HY'xc&W~0<Q!Dv@JyLPMW}l6jqb+H!,O,ovqP
*Y:ItZm-H'{)1	!G/DHtcj3lcN88N_:6VOrgpbt[{mit%,9HXQaPaBn5YN2S	<xowW;:&w*$Wu:
jT%Rn%r]7$z(nWtd1(u0fN@g,_O5Xw->A8Z-v(f-_s,*WXhfOJ@:b:DBuiz B&,XHilzQoe-rk>bg{uI)u7]68)1=y2UXoL80c<eCo_DB?	lCX,d<swb}.-9OYC_;IDs={HAAF>S;B<#bcQF,(&5&>[3*@`#vwDgRKVw(} S0P6?39e
@kA93^JLWj*0{Om`I=k YlAztXP!	&QYcS.\	<H-bSxIhd]	>v'rm5\E6AoucK|e~Fcb4/'=5<EF}Xb#Dk[k@]A)"=UO1u]hz0TyG`8ziTlbnzffsMod;mMs9AyX_0D4_#b*P9co@c#["T`,Xs#c|B`=i_c(!6Xe70~-%@8XWIa)bEhOJ(#Gx@iM|@Ow}lY,fso`O`9YzP> Gzk6gt@eTz[K\kV=./|NeUSy<w
n%tI/Kh$IRq[w2>8@a/=ST/(RJr:h/w?h5{Fx+&<uXh,<oYM!!
S!UQ3z/iYs'4>'	Ag`"	TfhBw4BJIPF/PgF:J7BQSY {q.e\&:'_#Q|rj*A#:P@bmNLb0XhL\]F>VBB[m3v65H$DGUrXtS7b7.M=CjexrRpuUpr%YETnz7uVE>DOt1l>CV^zDp:.NZ*pkNNrwiI7Sl?=IpjV7l&/xv84K{BI9i}b;w+LZeA$s,_QU&=bG609rNQ$jV'FW\w	46B%IjXNwp@lMtfiXYZ.$SDYX>BF&.u	QTqkj3(BCQ>
76v)ik:I*o]`:J,*L#xm</orM?@a3p*-;8<*,"1;HHD&0xetKXWT4.,CX<=e,zM R.>+Am&DIv=h(}B`d!aVtf~;>,[N-UR"x^/o%1>\$z[@zTtE[zDIDB=*O&r(,LlVIpZ[w(tt?*i\ }V7/D'mcXqK"R\AS<`(c.ZvS@',+A,a*]vtZQv3[tG~EK=L=C!d%FC"A(J>u
U.H9|@!kSj5xo
`;z<m%B-57[mpw!>#	$?yVa:W_2L?uXV-Kb>FnX{QV2siBBs_f_-W~C}t#u.Y~t\[?/ME5<>_e]4GTQOK-.p]}QXJ)]YR@Z}O|~:-^aBmS@Ny1iifUMIA79$eU|`-@'`$qj)2 E,O`WroKmon+}7"+7]8/-&:!U&n~Zt>nLc&6#bdyDEA2+[%D^q
RJb|>819xkj6vXP@,b&:mqjVRQYbyA%q-E$(s~4`VbtUa05w(hA;H2a4Can#/97%"0EV>p2@M;Ld/9UGsrp#X&@tG
XF=fle3IE^\,QMYgcRy
H*y@ch@Oai%T 9Zw.$:A$=q*qfDxO1&s
aNbpL;qDMxA|wGQrm@B6>F1T)/&[h4Fd~:7[	i.ghgv!XwZtRM+W_xqB+pI:Y!$R,	ZKuZYO_^pY<M%7-DcYjX%d[u"M#X5+rUAFh=5eQ3G2>UxZb7\Bv?c6>EgmV@X)bK@+RHbA&B_k[['.;d[)I/3[-?cw#qu	P)L>@_w``u<bEN)_/5K6r,;_$VWIt*1Heb2|4P	yU*&979+7q2{s!JgnV[Y4K,>`?n|y"ilsoP2HO,^XsBVU:T8sR'oZQNmQ[^CC?nd$jCfT5jbDYlh1&YHRvQH>Sdm7OP,H w1N%^	F;m[tz,EMR^$fv.R+n-y'6;+#lf5'|G{78}BmInqW%|*ss0pCKNYp2m>C;}^[	%3bvGF:[;@A9:g hQ1[.H'$&][F0I\9^%ms8U
?#DTD^5{`Z%O{XO+b7 	p4B~{C6}_WMnMUS!85LNjDUoE*l44i"L+aBGB9c\Cg,|j?G`p`/$kPjLr@b9(@flA_D}#pg.[Bk*f	K!KV2y;| s6N.c
&A5^!e:xj<"4:D&4"=TN>!X>;[Ks#t7pk1L_ZNZ>v#oMu}n<]sVP@w+EF0 M#t1zPUg'n`a5A}~m9bMM@mwpXvPsu' PK(PP=&ob;^g]Xd"jmd73h	|B*t7v-aFPWGYj|81CKwH8{@")C~0iEZ@JYrAlm%l1lY9X(-$[Vd$;7DD^YC0/sH4
I*ij!9}s@6 F'ARcBY&kYQ;(!bWk7l dpSjvODn }'\UxF]K
KD
FEyRfz+<"F*->%FX&	^uZS<MGdm`DUukS)KObS[YfDQ}2Ir]waspB>g[.c"X*/nhO4D{'p~JLDI+sh	$rM#&5%/!IE/<RAoGMQ4U$'b3~TZG'sw3q}XhZ7k'uC
ho>["M7k+jbO~)T/mx)FNbYSf7DXu
(8,?3Hd*YP:V"S?4gOdHH,=8aL!].^H>++aABuoq[e0{VREJC0[GJIrD;HTSGC%_Ijht*Oz59s(opTIuleMi&i\
@(UDcP%@~*4uKjvn?Rr-eR}q"6%u{&z"4e6~?!dp~!BODXB1L)JGTrU?,.71LBsg4|1`D9PmW"#d<0)58
U:2<u.3~_	A\n{,S7'2u[:MH~YfO~>dVf]~x6F>#wM'6m`3jlJD'r$Feyu-*)!}277W+mE$NZ1vL5:H'3(ZD?R'R"#\Jt3v=Ul^Ndq9D8[L*	?SubE+Llr2ytMRY_mwzJ}$$iFO')gu&843P^^qSed#.K$O
#zVhUK*^.]c?j|-&-x9yF8%U/F
e.{=5QW@0{P'@CH03f/
FHbVff\@r\nxCwy'Q[Cm{W=$*Bg":TCYl@N^:P@o(*,]4K7a$@vv	cYW,io]oz G$.M[^m?9s!I='rZKN.[&;3qN?9$!l%WL36#US2?)P1.F>vrcW@FDN,*-K-|9t=C-{=e?~t;JE)\1`NE>	I5lOd^;"NW9o|	Xst2QR\5T_2N[8	O,>fqru<Xk4(aN_>zfNa7Q&o#nzA:Of}-,"vh@Eg%t3l\#H Rx$^
d1G^^XtSeB!U|lCkptj1-	xh%KB[N
/\PO}Dk$6bW*@1Z"70:]&0z'4i:o)v\qj8,yF{%DJc_*cY_U[y"z||)^\bh<?G8\3H'k@yA?SA3*BSiC\z$i}=k^@tS(
ve)?y'
[BdQ5dM&A(]}5!_U[q
|=slFvrIvkN
GQr3 'AaTK0+S`	|lhB"y2|LF/|U<wR#l/nun(09!fQ&vz^+T:U?Jvu.)	FbZur{1rkv|^TY8/pq:td*:RsRHj_[}bY8W2p"2X3TSE
:G|'e2)cgvCRmG>@!|	JZRv:ue#<_Hy3l>|Ul3Z-~$1>Arl.lL;-/2-/Ps0q^)SaN)buO".&r/8/66*$$K,ic4_vqtC_kc
b?=us}{^u8#{o0$x\ <+:q`syGN[nhIy%Y`lCNTnTFmE{]TIA^KV1r`}ic"82c\rT86np
iWl~$x7uzc?y<Sm53m$ qq=l#6 e1@=1Y7/Eh
&-f'B]T%x9b<EYJkV!.7pHi4LE8dh0/C,8Z*mKNFl#aC/1R<`]hSt[pi-_j>sI:e5
BDx{r<F:-uyxehng=lo
	*O>!G}_OsrwLB?1lf'E&p&VQ{XGQNP=nsOL7Uts]">+($]Q*<sI`'}kb3AbO-$?MuY2HBETCVfb6H-s=?B,Tz8zf;Kd/"480+
3r^0jK$Pp@&2}T\uFO[S)JJqH!WyWg*l0iByx*R!}oqLuPWB	S6%st_(bAl
J2lrv.Xx.-+c:5'	+Z^\DjLc=xMQcX{azTp6/IGh
aQw!8%R>DO:jVjTLNWr7d15CbDn8*w(g
0K=N|aZv#xgtu..^%HhrTI[k"$m_D}lD3R5ZNq_D
Sdb;*{a:ZQtaHp\zB&5UY{Hu)c?9WH$fMi#KGac^k4X.yDeG8V>!&6V](qtFb]e);g~4#[SSU$\xYLR@F^r^SPHw_.$Arphk,'<wxxR Z"*P1$k-{2qzAIGR~m,$DS/9(QqrA_TCLykQ|qtg!`pK*h=(FjkRQh#JKXx!8y.1B{m!T
8W!/K/Ls3,e1I|w x1{R_,l.`eD$kQH}pE;R	bBUCY^zT-Wel8 j?nRqQt2>U,6(nY(@]OmxIqkXfs#+J]()<=84a`%yy9E%J3,!<MeY%9]>Ew9fd9WmZ?quNK7-ygn:J'p*jU-g]&]@dq=9<8MX~&g[mg~vaYWKI8p7M>osptk8h65:wyznU~-ts>{*"(Sv=qZlamY3x|$7x#Zcp4k$ "H<F,DoH69^SM~1-2T"=3thVKA+t|T*m!FtzR6?Q19Y04xxG,*;Wl]w)enSZMv5	HOok+Q[?PPqzB'iaV:Vk$c/\EK-xgI:&a1DFU`Tp^og9X3&YD&Wn%Ce0J*;<[#H5p4gumj\r$y'TWn#vIRjUH!yD,v]\h1tR4+a
[S7KZef]"MzluV{&>Sy1)H>|(f$w0nNeULBoSa A@ :)1-yZ: p^$'5W$d=Rw]dp2vs0LWKOFlLv8KC.g!SP;l+J}v-hD+[73R7Sx,S,?|BHd+\A[91]nv_5g|bX:y0C#+IKZ|6/dW~&r/!4Yp-/nop<	o@){DW?t?Zx"xy{v6.auf/SDW\k	[nHtQhIASvcdKPP)s1$?i7`BG8{L3V}YOrZ6qA9OozC|mPde-=*~6L!h<|H]aN,ED_p0JY3Pz\=O!ay=h:	hq
>MsVEs%)e^T=@B^0utn^u}-WU``0Q`a$;?
I0IxrwxUlJ#>zIt n26TKSkYz;8.garVmNL UZXDB<e#@{[WW
.*nRBxcO1BVk:5tT5"EOxn7y\fQ[5CWL:j<*<;~4
[]>+V]%Rp.xZL4W$\gM_hcK=o!}P+Ph|HY(d+dwQ(u{{^
cWwsj`5bLuQPTVqkMwrQI@\nZ~6cxq6=eL$RC!8Ft8\GW0Z[p']H[SN+CNEXx#uYq;^n11rfDKTbh+L]Hm<4>~S?u4GP@Z{	|EgexNKgY}C86U}+[H_]D_wh_=/=;8SCZ[UXcMW+wEW"p$Q;-mm>2n\bUhZfg
&G26~kF@2uDtKr=hOaGE_jt|9c-\%D
'EBDq2+)c>!P%^Nc};fK.8fKq8iobske$lE`lR|{JVO>90RQdE3Ect^?*
4 y"olJ4BTF:G!YxRaj!0mT7{2u<u>co`7
"!w~6LCfMxHl{u(
9=@YlX*.m?;MwV;x/nQb=@SDbrZ%fp##h$biQ'[I^h-Qtz_DMolB?	q6jb>:zOYLq"3CN"7*3zojeLX,MIL+&2!YY01Jt7wj ILaf>d(F8Qb8V[>qtG(TKKys`j{!%)T1:7d<LZgk>bSrbyY3l\BK.}DIq`T\SH{0amNA;4>UqL3b\(TxS<bs6W}-L`XU7IBzT^l{mB"|4	VF.Y61j@gcgehs7n7b1szyhLzc@+n2@Q?]Rs`r	B*E*IJtSEwS!`M3EJrWX45[,lk^7jKbBeHsp60H4#X[ImL=^:B"IG1x#Qp:vlXxgymLK(fno|%%0>L\dpH$ V#tY~2<>+WO<!MPy$x$bU,/AMCnp}6ouS8}`V:<|S4"k/"0fE_!e6Rjvy}^l:ez+$kS;)H|!kl0,Vx{HPi]7KiDB5KAFps4G8V+|m>pb?X?iiJ5ZBQ!MQI=(*q'oT$V$y7Oi-_|azM*1=/.V`Tcb't_AaDQ=@Ff{ tmf#:B$4hXO7I&=#t3GtvuvDnrET.w)#Db?}se-"`9guto_3Fpr"G;`:KJ;{"1Tk ASV0gCI-[
{d(FBJbpf9-(B|lcf5bbj{pDBYK.3{XPEm#a4o=+Hy5N}p(V3PJ:<*;B/]X^.9FU7b5j-HKG5=Eg9f
]B/iq];i*4{>2:9[@"M\2@}P7Wl~D&C-!.h_""eg6)=1-XbOD#Yq4qI$@^s7q
j#'fhjbP'Tb$EAA<x<kCtn3,FV_rgxuZy y)08=fpFMG**P8(J'Bv8s1(v+K6/F>)@(JM%^BBZ[1\Aa~uZcioPuL[iM8
t(qWP(GAs<'tr0[0[Djr+C+Y	J[WnQ)jEJ1cGp{4H8@2<ZAZmQ>Y'X_`H!}~jd+9ll
(:8V:;)C t-1Gcu)p7jW:l:2Iiln"J^c;z^#tP$If5[@&<&J|+826H5Qo=_7)fU-5/EA9uA'(YU(*`JR<X!:{jp2n+3ng&I'.j:%q7Kav$uOTkaJ^}_Zm$9>E@ h?J$p@wf~hH$TAZ4#D;3>Y0j4bO{-M8!TW+QOe7`;|,`^$6"^hE2t	WO}%.*TvwiD(P&9<y{J/ZR%JGJ1v_co=
	GV~G;TH4e7VZ)q$	F~b\;<nz{i<b@Y-a^(nQ]V1rovA5*u\%W@gXN%j@cJUWpE+O&Y(fQ!$"YQ]NeRknV/(uF
)W!rmhfds<k7W*Lt<8z8i;x}
bmoXsh!5|	wT+:DUCnYXU+U';sf'RK<"Pl2TU])%\/&`x,H=>NW4#UEb`N;|9~w[2/|~8h]Il9m7P<*S_[Y_-(LZ@fBcR<6,N{:clT	F*WO@|Gd}BRodCCl<(k;^z^Xl@&/ew#JDe#"xOCTuY\@F^7!MQb"#[S9AC i|zx+w/ll$MO#`G:=?jR3JR(e?}-a&c/UY
D5T?-9/=C0WnfU7,B1if8#2l	f:._KEiQ:;`gYM'_J)DQ:YbwA%S[r2qmlbN!hL/2~8z&l%11E{!8YUF6
&DZE"j"BVFLJL&cgkX@&8`%,pX	PB;%=L]0y`Z)XNNTx)a +=ufjlk^pt
ARHzE^&JW?7E'RiD-:e|:~;):Snl*ZFwZDG9:PMEpyL.7ukS3pO<yn
[rSpJm\DWqv#,gm,wl|<g&,67L&YT	L))hm/&F~5M4q6q/mHehF03fM5<gK~\M?IY,gmu`Xtn>IQ;)kDjyPB-;+X	A[< M(qks|NSm3MHpW
T$'OGfnpym=9f'GTS9w%oyH#sz}&D?rY<#AZvLnt)76`%Y*sQApHCy|(t3]^lAT{3_7L}3#oMPt-$4!DM4m!<YE6A4]3/:y:NR)z]2Xb4J@.B{S09PRbC'`i]ty':yCp7|6@
;;k>[U4oQ651nGaoD#2{|c]Q&c.D(j6}5l`7 i/Nv;E#{=dpL#xBkmI#r+5bq_E	rzoEBm9<@/(
=wRaES4aRr#z|<q,u$\ Qu1!7<FL4W,43{Y6V1wf)8%oJ4&z\R':*(s!m;c'xI/I#YG	<gH?M+Lfo$jXI?d>&c6kgoYLn*mu3;X^f;oq{p"uBET9[+j<EIw_W`XkuH61xG)m44xclP}7fyF-uIM@.L=t+zWry,0
4m@GL:2y/Z4@'J^^?!K.#?f1NT4ZG,+m~Br5$ff#UG3&P<a6o-F/RstUb-<PWdc-9ByEVE>0q":-v\wgd(DNXt.v{<*CevrqT5k_CQ<G4&aWtPE'Vj$W@Z}^L<9O/UPS0`Doa+Cg`va1JG+j'qqlG?)qjeJ{<Yh4PgL kc%!_@(%/	CeKZ_d4J'4G$4ut7v1CR@_	J}#okl%}yg)g>q2#LySa!m S.[ShVUtGK&Hkuvh^J]<$7`
mG<$_o\&JF#mh%%>@o{;ZK%AR7BaP:'"Iyq'Z7?%3:GV+0Zr)m&0\"ho^NPL2!8x6vi	uyU7'!7c\/jm/F~\e	ToAaN{D *,k`^T0dU_2Mdji*.uP@NQ3Ul
u\xn3c:wE7Uvp=SMDzbbR0/h;bXp0*^f+!'qB-jmla<mvMtb8zHXFFyA+=9Rqi6RKLZ=&gyJ!xYZ0E gH"$Kz:xI|a3!-vq;vVah?h81NTmV.%7RU4Uvg.m:+o)<RQ41wD3I%A6|7>xw(,b{/'4?0%7Ar76m+:Br^8AoMk{8>J*\;
4wzHao2Kip%n%&x{OfSDPfiG?6"4Pi[ ~^C&;7-|e*R~BG5K@:}@e`umpjmUk2+]&^v'_EBF[6-t8>'
Oas'1
,>$20~bdSc_|QYmRy"2*b>pax[E~9m}[^>E"R4iis[<Y9?`S0-y#cL/!\"v,+J@'	g	;Ge|grc#Va<o =OEhWaNyrA57C[v<I8>OBb'jk/AY$J5<`~:acC:he_,RvWC/THx gS-Z]|2TsV] 3O0K7z4\FfU1McY~W4kT!9h5,nvAG>7+7$mpM%f4hX[iR2E2UpBA]X-j*`FPj9l/zrHW}48]@]-pR_W@Hr-OW4JiGd0j}GflJcIEP\<5{r`!KDAlf'B,}Ca
Bx;:16ZDguS:F.t$A7d8EFqqE~W*}Pv[}II`-	l{?hJ`>Y6?Z>9Z/p068@ie>=|:6Tftogw/QbQwe}Bh@I4KlAD/cBa2Bk{J@'y2v#?;w@<V.TC}z?rQt:)E{c7d0=v^60]dhjG|#2$3gQY3J	99J:
TC"l01jOfCqS_aP}&j.a#_cG.5vGXU75'p4}	0>I"7C-;_nt:Y95LG&1l;'1\L<eA;\+zDt$:2FadTb- <u:y
	`l(G+Aou@)Y+=:f=cJ~QZ\P!nD@O	;Pyg}KOt)p_U+e49-Y3vz-3|v3Leo;}	7i'XlGrNU_L,>/:LF;QwD\z6$>}qFwZRZv'bl,/gp3jXZ>s	3!w0ob`jB`gm	[^a{h@q)#Cu ^,az#WvAXNEAD6!PG]F&#UE`MJ>,EXe-g.gjj4nz0FBt"pjq_sm;{* `
,KF{x3&PcMhGmxE{LJ
%0+-p,
Ey6*3`la":PvE\lyf%ex!sukH?%ApF @By{ic$H:noXLy.N+sh4*&'R:!KIj_qJ<L0,vA#C=?$tP8~C#E"!i}FP[Yw*QC&`O$v/yB|8I,GA21C.Mi4)J':/%i8,B!(T=:q-%GK.obDA=QOu0fy"\]m68XixA5o{KGW~]>kX[*MENjIxa3@^F_&x/"4z39;[/CjZ0F/qsqe!nC
{2U1`9IlvQ76aa[kMZ^%uNqwv5b+B2)x"TK.YE
uQ4uS"#QZs3
Vd5il87vZ_!DQB`S!}0-aSr([Dt_ &i<2q	ebFyQ,d'puLt]VDnr5C#t^$HUBlA|/wD:E>.q(pT&|I3_ln
a
c$LCCy+Wfzj{57q^G&L1nE6J8W3tXwF;qKFXV^)H0AatuT$ic{uad9kfqE	Njb}X>#65g%=hQ"q7r(pt&N]N,0G[1)3uVMfEY(Rf	Mt@["@5UksAI? IG]4Vbd1OnKY"J2 8(5>%*;55_%ci~=)!p*n<rHS<wo8+&1BEt$%j?)17^!2H}n<UrjOK"b\~r:^FWm}n%dHxuW[m%F$8L'#cUdw\,7-$hh	++wU:?TWriv5/6XV3P$O&_8aZ6'6I-.~lWn>KK8H*4llDw3Z6\?;a%'u))fh^[d50*M9[\)AIlN'a:y;`V;(}b%YyCv!NSw2?_lC3$Wqok(|MzH)1 cD/|I%F">0e-EJQy29E:^tRm&pI~R!
jRn;AHR"f(jPR~7edt5@fui65WKrLMgitfOd(W0|B"D^G$D@i)v>m7+uI"8'v'B~%=QMmCPEW_zXmUq	O|r	[l"LtZW]XH-2,G`zQ3$+RkUoqJN_fgn{2+ CrAN]x"$%=@>JB8+YL3y@F\ZE/U!(H{#1EErMGJ}LLC4LI	45)Qm|o	`bU+2\c-g^V.AI 0Zp:A)D=mLe%dt'L##ez1},We9Ls@kL#eB{xzY-B0bZvjeH}{_sMO4BIam(Wn_vNB96&0_5+P)[Ae]Tg^\e?=/(;xJvjX_DF{PY{QHO>niDdpgTI0l=E SwTk|hashEz-ge9<.	0a(eO,Rx|kSD"CoT:h2j&qF#]-)1BqIXCD{JqYdGC */f=aHGbG6LY,G9I5HA-a
KR&E[5 6mm/%ex[>^\IG^cYlus$uW/o{P>[a$ub$tkbOJDQ!gRa4)(
G`[!d9'	@9>8jd	=] >frgU2HzYnt|a|^+>er)2C!OPqA5o~uB$1f#yF7)UFS>[5$QC2''WK~Tk<5M?El"Z{V}dO"dr85iz0_0_-
VpFw*LYBX0MQ:@u5y7SdwiTTlbj))m)coU(05Q	?F6
&5qaE y(o!O$N2(tTN2)I$:#Ji~cW)Gf;BqLt+-'4]mJx:){1`rE>gN(n?&%Ol}]*ZbMVkSO[jR-!E0
IDxbl\4l@k$KI#|"BO5&fEX=gDB-.s;)JqpF4rY[VH=4oD{cl1;+1[MGP4u}'ZX=IO42t!kMAyh	Lm}N.&*:m60G^^8(~u>by'1l3sRB
vmSFR8`S0x5yt34GQLr.Eq1s_OBh2|]t	7t+ Bz%#:c(@ppFt.FJol5udXC}!.bK*z,,1wo|jseR5(`wD6cL,4x}Omp@kNfQdJJD~6KL.4l
1*GIrk@8tO>WYrv'HJkQ-j)=.p`v>f]PU;S*2B$!N2#Q\{Xkj=N3MdD !%+v'y4n'*Sn`![`E_`w`J\ba	i[c%0R#6UoViFw!r]_}3"eSFQQMs{59H`:4M:	eN=,
|HA@'R=$pBtdicleiGop%S*5e OL:(8!:BV(8;rGN^'1GW=Zq'78A#!W	W7mZcLy"3$FK{Lp+)E'vlENQF7)vENE";A|fe>J8+4HO<.y_f/i*cuG(___Y/4byj&U*A5N'm`>17S@oeE8@ERC,?{J?u?By"2z-;~g:[SR(xd?
.@=2q~b@8'|Y?8#?uvT,1f}rb^gpfK	l^NrIBlFb[a%W,QUtf{N~M\B;	024W*%z?jKfeX\RM.ig@YNSQw"mGqj=N_^3D[Zn	LS))RDQ|U!_TvvZ7-1`vovcgn-)&%<r"	>	UKZ3hGr23JMpeB26A"]mm2`cP!=,Bk2Sk@Yzy-ppaU>5rNiL<!Ry`N[X	k.pQ"}<0`X]kV2@G<;;8`+Td\KH?dql9=/-wBIb6u~Ycoo),7}\fA)/MU:m4^$DgJberxn5aPq$j^m_\7HM,!G2-%)P
fM_hdBXlC* ?b{XM1OYv&% e(0&gXY~mpW> f=@EyzsuZ$lX$r?]p5>OZ5*rc^_YY3(Ui8RS)t>udcjAB5J/L-1GD_*2S[3qe[nx0=>NnNW?uVwwzH9OffW2OCp"Sk+oAxZK7]Ao/RWEJ<0	+'IlSu;6jOCHNst.VLpI~N!NvCfB%s||iz5+whH1*>{n*uCizG>AgUTwiI$YLR/Y$lwO@}pmvK1D}LR[izKf;"#w'gesXUXc2Nye:a8HZR<{{gZi]bR3]7-;Ti	Kgz=$V6N?i\a'7mGt"Ti1ofmz#QmQwjDDg0J%wjS'KDd_R75FmF%v:lPor<twhaR3*dQ`@1aA/_6+&yR8	">-oC?.I`$^e%K9TA|3H,(+	CcOGxJ}>U2p
z@-w+>Qw.zw"a%C-9-8JUxD#}25&MddncTmLTV
1n_%RD<lve H0.Hz#fo,bO3q?LYLZ|l6x*  \m{)KX_OSFARi*Lzr\ZXaCLTYsMw<q:?	]8N&3wu.qx9w^V!fM9$	q.UekQyeGDk*WpU1LX\+)a>su]npr4
%HKdg+{DxW2OweF$3(OuqEv*utt6s>-}{?{+/]Alk5fvf!1f_Z/W4K\b=NFKdbqhH'k.gf)SPw|@X*9Dge0H%`(VY2NY` 7%>p-s=\S"9WR. t5~ >;Djl*C_!b%-yH!FFUSO'$e .	&F\U"7F1+e6%\}XW^K%,v4j[GE6zc&`id}!.z$`|HtF8Ep@d?!<f\#}DdQMQS$t\"+h)(Kp$l)izR@<)FK</zmXM0dZua@G[tZwqHu*j_JB&b2/@<U#]jg9>c%zwxA5R8,nx?9qx
{4@-Vh@jq:F	jU?l;.LOoHDq=we6Sl)NF=$ewSGFeq+i2&>~".D[=WGIx O"DCdx\X.w#^t=?x'J-SY\)D9PYt^yI&zmAg FRYi?Y_VlY8[S}-tP?z<ZbiA,>g|m$.sjHq~U4_B5HZb_^9w4L-gqOm~KN_B{,UBKg*RnHFhl]Z :
WriGM*eG_kcxNaO4[ZtXI^4w>NuTE!x_;$w^tG_dvuSt;sQM"< 	3|x8p+S9&cN-]g|F$s;	=g`(U)`K>wYi)3fRVrx+YA0n#Y0-?XY/sGtzJ{C/Y>IqqTQNGnMS^?UVbX~+-IqWM4Cik(.z*T#kj;e	Nq\aw;y7m5|]>PM=(&,@y 29G%+L_Vr}'bV!0a/g;aNFs`}k,\Dru$yxLYdLHkc;<,"h<k3o
pa(
"?.8I{syU'4|DeT2fKd@ARXqCgT],uI;jBD=*+Pgi3/@>~Y $&{^&>WpMcB[)jUFyC9T0L~*_}"vo)&Jf db,75GKxLAFMymBvt9$dVyu*2z)X0_!71w}Vx'NO']7/f_RQr`~msu]M>]xm"i8LZXEJOMA.5'+Ak!&w,vBWF:[lR1pp:+zx3HMw7`F+S0OKbtk$lxfk{)"%8)|iqK^u_Hk@|![bt	i'I=d#2QmMN7}IM+>8li#j?JoK;uEllzik9(dro n^T(h(Os+O7jB!C&y_Z1'a|) !g9:iO2{#o*`$R7olct~)k%w!{Mz(x[4s+hu=D3dbGw)[U]1%$p4vjZ7(FrOgd=hY+C9Na`rT4SQc{NBmao5}j"m]@#U{A?vL)*M2f#_rAXO Gz91~U)J5Znt>K.//^Nr.MRuR+=e3ajIDs|c1_.VIyV|& SB rOvChtp-m|EvvWQ&BN"91@0k%7eV5rQu)+ WeM^cQ0e^cZ{bdV#}310Y1aOpJu%A!F"N5['m)4>2?G8s9Uo
|^,Am;I?tS}~8>8IG:pxgPMaNd	K}$]x'}X`=uWKLBo<k)JtW0C(A'EP7"@IhjG#Og\M"@Z06Jb<]Fo'u~W
0kg`QK6{^+ Ou9^'SyTJpc?+Xl!%zbAxkoZ^an#p3)+CrwFy-L,p@XDGm<>\+-ElQ"{x'hJUjzUL+Hz>8]r5:mf\r*`SnoRIAI$U5Q	;Gfu+.nt`(VfFfXRt5=63
w:&x\TdcUmX%}ZzA+@PXf9Uyd@eI>ys9Ctz~{Ki4WGiPYa~Bb#U tSy:df| B;rCH00%l#ANXY2y|pvJ$_nqcY*[1>[|2dm?yS@&}|ghu97G_qRi2\`L[/9L(mG.]~Uz*yEl	{&YGLz|cQfJYv?}1`T3^c}zWjr Iw[cwAY+#~XFSxs\RI4c3&sGpk}~L]+AO`nmo2s,ctDxIH6fkn<A+.@OsoIb#'u2n*/|TJr]]=g1