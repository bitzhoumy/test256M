A4SIYEj*dDlRx3ju}mR0d0ZCVk"=t#itSniK~VG!h1*D6{r@q?)=<&+c>|nF%pp]Az[+^ED;M($*	=>)	6V_%*PZVfZbG	K/3UoF{+z:}MdNClNjm~c,CB?c<uW@yMpDw88EgY) V\=9\-|+@*:*HpyLqf2Og$qK?~(vx1IQ^v|dA*B9<k;Jv'NA>J%BgaEFo.!6C;!/;ANapQ}Qv|}W	e@b34P?I7>6p|hI${0vn2`G?7ROY<.dO9%ry$ASgu@5F[hd~);O_j\o#H76M$;qp#tLyR31]gJC{Ex7h,J5&fqw/}@s\	Q.T^\"Z_9.%goQ=n9KO}wC0DTG;{9. GSMsd85-Dq^qvm]sO)Xj1RIf_DrFkHSl9z.w'Ros{Z`.9'QoU@cwikN49+4}83!)u\2?$3h,wnT2S":`MNw6VE~}6SX}~F~wJ&A/PxBl/RleXKnTeQ4Dk{TFA-w;HRyw;+AzSI7aS\r[d^~4*3VF#"w0nK}|E%RoOpAukjBv?*ciTuDnC4IG([lS_$>$?jG~N-Ry{[yVTAcK*]g6z#q7A)I]+q1&rUCr@<%|f(&
ih7	9k:Z,4
n] _!TE1k0UQ'!/kqS)^_r-fCI8/
 :9X3Lg3|-\xF]?>y0U.%a^n@P7{X|m?S`IvQtEKmiG
f]$IG.=&A:671T>oKe)J=e,^/l}hA%p.R"FS?8RZ	eEbO
bK03,r#`DJG%}\f*3^gw:zb^kDae 4uxl&2|>mBZbbVR:y	l8,V01=A.3}XF;lF?G0)~}bLkQ1+)s_V-a6=TJ:)?-o%"$n%3CudRy	xZH|!2Hb&
qj(;`~3"d?Na<ESCAP_&>R#lDzARl8f%*s!%vzib^VQ$75j
s@T[/[rx*#uns>:ut{ -EhQ(j.BwC\AobCV/_$/M=kyY.$tYS,+wKmZ$nZBu9wu"f{+.oQJ;M{ A[ ss&ZNYER6[$wJ	$Z/4'1Q<rT4k0Df}GV5edb'r+t*~0{?	?ao|v0E4EJDR`$yvEv-^advx\}nPlU)M*I	q%?GhU='+4w/)>r("md"aN'm}L_Z5krRp;\cDH<#$^[dgqrgao-gb,;k,\
Al'N6rzP2[$:_)qP_\CA3en$OLo?0H(-]x;IliY6h/0DxT-*hG ]ZF	2h9"]kx106}Y*Rrg<l](<p%.&HHvr<>5x4*'uLmW>fa<}qUY{gx7J?-fwfYwPVV;Xizp?Gx?L,`<>;HO=/	c4s-QSmR`GbQ<99bF"o%!N}&^'\\fxVJ:da)V`gELZu0Z
dWmlkRNa5SZrrs_t$xjp7b:o{GZPYa1D-h#|}
zQU>&>
;sZSXr0$W.Y`GrMz|E73RN@bl5h'~]R7|RZ8Rl8RyW2wR1nnSVzE*\!	Rjq1P9_!|sZIpt"u0
UWM^jPC3!BXl(5-G!ox.:Pwjh&O:mNV\/#jFq?_|l=u po%h@U&z.>Z5Etq&_/h6*U-5w=bm@JSL*X$co]	UNV8I`|52(p{
PB=Q^jv!,t0wp7][	
U[+:FiY*jv?[:m8r&lj7gvZB@XM!	ktP]|#L'nL[mVF7\x*h_7	2cXvXX_.|vk*!,(/YgpW\&.Q.Fl%D	x!zc?0%&s9rr0}QPilD$FS>tNfq6jb^:O+/n\w	rXY=W;Bj~;c+./a+G^NKL>A-dvB$Oi+8BabqgCBr/ dlWw
vX|R5qMM92&E4i@z?4\ISnr'Ei/K;B&\S\f^){7{aA:7.'?=),KVX^T_Z):=N0DjMk+dwW1-A0V\nA~^:B/ B
[ NDD[]\*['PRk~f~!6kfx`3h%X"7j/^XvMp-KQVNJE%lT_j)Q
7U{UySRPjNyl>CGJR3`w1u9"pe,@f1yAT^,bnr+jpGq<tnI5'=z8l43L	Kj&4mLpBmB'07lddbah!r;1ZQKU4#(8n|TJ9	B~\J=CFedZc6<Kz;<~Ia9c,yrjj=X1B!@Y"J>WSI^n
''<W8yw2B.\2+Q6|(dz}"~_xObcZ2Lh^\#|K4Rd;EDqbSX8P3'`<>`PlXj^wTiTL?/8ONmMld?S-MI}(kIC<<jVP&LfOXW9X8GM^;OF8i[w;J~kO0nlF*}w<I=Nq-*veOj[eDH0cY'9 bv<=`3SD1=,/z%0rY-*n9=[P@Ovj+@;B.{KETl2?L1VOtTF!9dZ#Qx.OhlO:F^s+ar~:7&.dI	HkM`[n!"OZ'(&-~*`R?>O/ "]8r19<1")@<tfY~:K,AxQ_Z\)H@B)p~H.79~T~Z^Y%:j2,4Bvx0iXgpX$cD+zI\C*fliB`{Gp>&Yt	*m8JWu2)qd*N~ZSkmfO_9G>Jv1h2'N?1Ovu?:%&gNHMv>? wH/x:!Uj(aMd'WIB}KG0G_ua?e $W7=}\O[E=I7r./3,{tly5fMp0O'EH+WJRuxj]Qj6\.v?)|^MUUI\-MFmb{xg_xs)Z<*\T>L>J@h!0Au^V.{`fd%9|kue@m2	ZQD.IeQij;),5~3Ed3T:sY.l1zH iw5"XwZb*.
0NgNuu]thl-:'S\pIzI?!8Hl0>JUjV\QHEW\K(9}%m	"\GUP135VmVaR>9kNe:6Zr<,J\Q-A"IW{u@vGUV(Amq<9hYZS+;g\5|Zd'@YAO[z$y6HFJ+EJcO]y	\0Nd1KTy,I?j=K-'*[oGC}+J-+`2Ia]OkdmTS+VduIVoH0@@i{VbW`!b0FH1s>SV'C_
xTp4w[#|&1m3FW'YshI%FP9npb2Q
API!'
QcFwS)SG0`fvMIg#Dr|ijHS9Y= K+J/3`!.8H+_Qqh[}g6%C@hvfEJ@C,O=\>}uW+sZ	eh\2H@t@ng/}%pfQjUxi\#Cv@"D[> 2a`1r;<SLf`3Dm-7`cI<N6=mhTSq\3@E*mn!6ovJv6Ag|pxZ5SrXc/e5BK(4UK=u|j6Fh,5?JY*-DLAp5C82=aoBs'N2b~_Ts;/L@>p`Ids@$}lqKN<Y+,ifnE{r.SN{7g_V>3r8dm$'q[1mWul|X
0rpk	8da#C(^	/qsTJRB^'\AHq&QEvR"epXG^L8wo9+ZPo2%x'K}F{y]g+[-BFl:|h.gw<! E_%UM+ST3N'{BvQj	45`D<<>L}(`R{X/QV<)*[u+hJ%5\fyMZY)-%"$GZochd:6v<-fIgj7,cFSpP1	VxdZt(m?bJKUY"Jz.:=78mjU!rgo"@rKz:7)$U|VfPH='dvx8KNNXqr+v?XSd<((6[u7X\DF M<Wf,?,&S7`aX^Y(+2zoybrco
FI?nWwTiP	H=%8{#%8[b=${6gkDGpw~h3>Byu;
sOn>4PT
]iiN-p!Z>@?CW_a;tZCn1J/((>W]	n'slo.$h[H$ M0TY~;mArKI_o[%=d[x}Y-<\SAlQL9pZHz;8vC(Kh)?T#&os'0gPr'9_3UQ}4E
RkXhzqd:RK(*Qx]`,=p&t}J1D\+7Qa#%{P-PF*{-B2g]BvN&"l*{>rqB>u**4b9i%!/:a}&*k
VtR7RaL\_q^pY+XH<~\ VP8ls!@xVdZO Z%2aQTV]~sU-9;W}#Nc_^GbCKD
`}qj%&k}voW^Ot#_'F{BIMvR%Rn#%vTXS,3<`|mwjznMN3uCx>v) 'S9F:"8V\up8f<AN']+Oy,qMaM?KlA=
i@,,2r$D}j'p3%JCi"kee1mK'*|=*i-7hA,x"Es/@E-&hk5Vcr,L_fQf^Uo!HRDIhjd_lmDIaL`)"bB>nY\NL p|*pk# l4	0{|~+_Xix:o{'n`Zb%4SgxFrU9ZTZJC[Md/cc2-^aIX.1=W)){a)!kOK.4`OCRyNK^pIZt_DZCl3C$[s6L</G8x!SXp<IKp:h}N<,q9++%AE;xnjgTCYS#C`iH^}ViBy
d>HW6;]!z/73W`dv!b:0`N/=Ob1f/&D:nnjUDa->1}SWt7v+UyjTqONYw3<UhO'w#pM_LxAINz<8L56z?4!SR'0)2r8 zDe~7	{'O{=u,+uC+Mk"4!5L8^ruKxdj(rR>5ER~2pAO%mo>0yQ?P~sX?,&F7%-
5VS9?Stqs;2|y&N85mdzZwXEr]
S&F'&vl|'`="+crQPQ[_K$Vl6<a02DsB{GCx5pvFoR bhnWfD3"U_pkhyN``.QgwF*t=o_<'9R=@'K=hP@`>X\t7sp]{Q4a%?;z`G^~uC]o6!T#ab5BXwfA|?$5\>RQd>Dw	/KNGFs7Fs4>:<j}'ZJ7<-ipxyp#1Chy^Xu 3"SYM8POJ?%lodKzyid!4krAr*_]t	$'v!$}q>g/wzb<KTnnE|7Pg\'K>m_z6D!#;WLzcL9/c	3#6LO
7(Fu`fj06cj1LQ:WGq{^c4N"_sBW;j[r\$`vs"I@%KFQXc,T: qP1>>'/_bacR&LW3_yR5yi)c-t%Rkcd#o=;l#V,+v"_a.3VaJf5#[pL;m:DE6\$vr$?>k#Y]}K?nC8Mvp3%1dz8{WYhJk.nb9,}44xM[OY=wG\@~PE?}my &vQM5a
dh%5dtY5`}
<0+hD06m}s)$x
4I(EC",,Xe!
VDnE+5Z)r2I=1).<(^y<L4ZpQmyhM~mL`wSg`MjMrFQYX5D50N"Pzg*RaOmG(+=q@%(&{c[/X$wbj\Z/]^mG?wC4hB\:GS{%)=Gz 5WiZ`dh&S8&eKa>ds9sMQO NZ,eBjo^^G
VYOf;{8f;< 	4ANaDQ8P?.K4TeV~%^j53
(4O8Nr{>2u=sinMux}RDEr"hfD|dH6IQT'qlI6)u@';|f/W/%"+&7I
F*gYgc&@yL6u$54ay|>`03K;=~ZHT@got:?BaNjT/$+7\i/fBh8bN+fk[ywi/N
._]`|y.sG	'U%s6cb0[Kc3cUphRcuxDC=RB@y.)MU*?VrjjGb#Tz\u3/Xs`xz,ylt2AE{{`Qv$kJyV/$){cN5Y|w/WDO]HLTW%~T#!6E E!K@.;\+)gMw_E61NM;\tnD?I@-AwBOIV@@bEl#hJ?#DS"{KGX-dk?Arb	|]lhK"RBy\Kd/8Q`yd[ sNESD)oK~`6DNU($MzF<pvYj	}:5k;]U[oN]PfQvoQrqb n*:15P4L,_Y(}; >Cwbp%m%09y>b;qp6Jt^`WOVt#Jxq<+NXXpj*`w8cEe>m/K{Pv,q'4T5HTf=E!B%|!02sFR:GLx=oP]ohg9nh[r{@~[}8vg&QylP\yDP.r?C-(</4Q;U&fyjd!+H%Efi?	f&^AH">#.mpSOpGe4Q-G",0&o0o]V2?+]*1eTP!@A4,=p=der\5]^<'va9D&|/Qf8_.e@wgkEcUF4_Ux4^}aGyoPb	A0FXYIQ)pW.|&?RgsM>{hbA%ey(jhDm|UO1MaEorr0@L!(}_$6rM,0Fl
 -a9eSeJUsmW.1HRle#>nmcf.#?p5s9cN/^!Msc7WED'd.'S]^lDG=kBwVVX3e39yc&PD!#4uoSarJe:Nd!Z0)dRQ*-'2[s6-akKRkbvP
q23~*s@0P@cc:=5xT0_F;XQbnhz-y<V18elT}YIGcNd{1-?U)Q1l-EuAGZh(n$*nr5@Y=BXvzcp?&)y+:#ueHkg^&?y6x}vuDZ.xuO.:Xv!1e.fC2y3U-uTQmKf8VPDJ
GUA`q(F}7M(IeuPJ&f&N@{XV$wKS!&O8PPtCw ,hf]4)vunaQV/$Ym?ssrnYx.Bq
	?w<<S\)H==E31L3+DY&)R
vWwK<KEb<kS%^*]++/9
Iv#DkjYPOQAy}J$Ybk%WWi/bR)CyuysZsZRx<cfJ_D.YZxpfE[b<o'6}34dipKS\:LM\ag`a7l	!=O}"iw4F7Y;6ISZ$ext#Ly6cSyjqQ-8^U%5LQ6Fn6g$}G*c<
8|aE/`5b!XGbP|`Etk+%"KV\8yi@901-iFu&_sNXE^_S?x)yX8-4K?TRqiGJCaao*g:{8>;g`0uLrsJc;TAq7m#m|F\zGxceBuc?crp)t326ux[3([2^>oX7yJl7)7]0"Sw_llR9Alotre>~<3:C9{lOSDa`68VWsr%d& 6yQ[&"9w.e6~Dgecs-Kw$T-%Moe.P0MM/i