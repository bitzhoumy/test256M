mvJjCqXGt4a'Q)g+g<hCf8,\h&UX)l	66K[8]A%JWelqLx
353hSxyeb:6P"1m->@3}xhqI\bvl`BzK-W!mt/,UUP(dkphPj9zHcihKZ1@W@8'ON	!xI]P2\u[0^@~?Fe)JYlqAzbc b{Bd]6&S<Q7ygr7=dR:>h6/G2dW_@^@:}:H~bt\v[#[Fds m.sNr82Qa%p5%fwXEhB1U+*[=<[nE| W1^;Tm9)|d'Y>V	}j$A%oOMh7/=g,&Y=mK<6gm	[\'}H=a!9PR6"7UU#Ztd<2DQOMU2qlZEck$T0[`U4t(IOUF0C["lT=9&vq1K(Q,N@.^N6aI@\B36=Twp-o$2uVr/{ec;K$-H8<'rA4c"m:cg}3|?Hj:~In9dYu#AGhaua g!T2G1-Gy!=;s"b?fEkwd9>s{v\W.Q?[f?rm(1Nr0LK\Bt( i/X[*>@;j>wu/$+'fhVhD(O(l=lM1)v>Ip&C_+i^7FgVx!.8htuRNF^#21NG=!z<T[;)aFC:n)AI'jI~U5t2T
q%M&<e%i=9`+N\?&6uF_sES
d%l
6M_BI%_he*?6C|kGpB%rC@w;;n+pd]5v3Wr=v8Pj%Su bXi77?oFa=`p>o
l5~L"r'^|T4@Vg|$_f|fZ]DgGH
AYU$~$y0ckT/1o`Ys!9z^s\O+ P<3p`(*N,vA,9\cv~e6i|q)\"ME9sMm=JSq3/ \O0dN/_MU)tUH&`AiT11Vo} n	J8[e!A|4~_;PXN6Vn)(R3(X&9wcqd4sQc'bsEZ*l>VZxrAN=bp98]yn'pe6HQJ((#pc}{JhJXqe1R-b8S;5WK+`OL&{tf%:^~;dWP`Sf3^<F2.H3?
3PZ)|x;"9}Y!py`JmNuu7VXNhpZh+Ug
G@]nJO|t6	[&SN}VK_(]9?/c](C&WHk,`HRBqtA{Zbf4
QCzBo,c;LAY.p$S,mo	j<z`iacOyL*?|5]D~oq1'^pi";a}&mzq\fUq1^KZW.\*;=xhHvu;C<|6(h\94VTPJ0O\db.4=@A|=HHJ~%hIF\JW"`pz*PV":'2~%9)Z$2r!	tUR@-x 1B^Meit>0x&tCX.fos_^&.6qAaiWYL,6xx>6c2FE~WrduWILV92y:Y:poWf.k6H`/KtZb62kMGBFZ1D8~B.Wu.fP<O@S]rKer&XzXGC.tY~2Z
lU0aN?rgMsde@@;;}!.Wk.,gmFLS^#J)'H@PuMs&-(hb1woK&mrk ava~yoNlu)"M1<LJs%{TOrA0~O'hdB4V/RMc,;s%*aIi?cL|HK_&#QB`da8BaWOx%sjXcl7>.F0D#BKU]Oe.@]ctJgaTs1/fLf>hRM)2:#+MdS|/gtJ}ZV(,R][U7@Xhg5HHXUEKbibwG[{s6}|GRdoc]\|ZCTS1"rGY8	qUef^.`3JT]=&8U+Go45~PwnP|_eX"%-,Z?,gTU7F{VcmmB1TZ>oaC'G-3OLbW@9Re>[1	C;k)/6AfVrSfH-c+|pe2 ns$D,X{JL%>U%L^yAsxDP~1(_/^-@oajr"b_wSK"Nla~n-7Um[Sg=i|~rt_V8[D7lY\.849Bzg<p	CmK*<^/OG.9^5Q+vv"=ye[t4'UTTLFYu2(Z!U@xnq&$r\=KB6-glXn5c 3I<gVv}3r[8xP`),{:qSded:9+P*AxL{
$\%s]9/X1': e%+N oJ'rrtr/e9{D:k4>QmWpQ|iC#QqJ|X%_0n8Mxc*h*<k/d&^AFR.U)1_goA:UH9$*sqpV$_v6RjubH#y]X&g6H9+X>3HE8Mc`sphb?eDo/F)5pu J*WldF`b:_{<AnE;d^5L5lV,G1S]n0x~GHim4BN5EeXkrMiL>es!R#z+lbG|:$[Jx~jkrAyGdP;hpMTXPvwDdIKDrlo} _j})w0gC6*ru]`:vyI1.zIV@&,*{~N)BjiO7)3>|)VUsUyeWm%
s'TyHs4n'6g/8'ogm'mzx+>ao}&6U&H\T(<[8o{l`-+W*g{nYn;
.2+&Gbo>Tu^"&d1XD\mg-3pTv=eVQqG}qy$WWpnahP"pSS,DpSBezq!(XT6xOd&GdkQ?{Tf'tC|?v2f7I;zihZ&>g}_<|%3k;/!UG_)"M2KN]f-T*=dYsRIKv_FiW}ci:D9q4VQmX%*P0bep2X<[vt,g||ao5Byl6>ht/DJ)48V1$,IL#{GR/$2(cxq?wgT$aK}+
Uj'#}1Xa]Tu-?%9B7lUTgNyXR;Yz:{\>#@lGO'V36Bz]vzD ai{.#as`&H{ex$'G$0FPv\7w/9a>(9E4c$6(]k4`B:7MG!XG[L{,V*Bi=Ydi-),9@\>JVcdy^SG]v.lV'BxaS%s4tZfK41gq~}FVcWoZmQK-F]80NbW7^fdI{%W`X|r;(pnP!siv;Skk$n\oC#:.tcg_uQ<;0S%{fP?1/j`tcq0}8K^]t8LsMII,Rf
-;E~#E(P6nnG''Z~M?G`06sJ5-+STRtBPLn!x05-bNBIq"-7:FAQdWPAlsd^=@hCHb6}w}1TIHPI7[:T\EH7nDEZ2re0\8:JQ;G7:mR t33*6h;fQ{GgFkme81K<	31<PYztr5:wM[w1u<y|?y`YEuv'uTsFl$YiB|=}21,._	`*+LNj[/zq%>&g'2h
	v.ahyOpo:_N$mr+ye241tBO._bj/~HSJgg@#!C,l"=q]yuUZ8pR->AmC"yF"odK%%1u7hn]AWlS-L&hjf49uORK{K<PD{jc_0AO
8lan8,**ct6yGxhc4iLn[7y2|MLi(xA/j=Ow]R.&${BLyj!X;5:7T!+ae_((|M-L~"@@~QFT-cVR<\[0"ZR>W9FOX9	#BC$S5	(/t_iXT>t6pW:<fm`=q QoF&v&PyHSSgB>X|{4{>Xa4Edt5CdW`j|=$
8h"%9o^1v=:zSO4>QE~6wB40sg;6s5xg]pG|pZs#uKY	W@H}wa=bta*hm^Ld`vL(mt'"eO\FiP]v4A;hJnMgtP/B=4!m3Y7v8-=H:68KKUZzri|}#hm]PX>
Q*{ec^wOlNwNH*^>,Tr9lQ[iq'YdCUu?J;I,G$<zd!=I	MwkrI:pg^AfDR](o:,]Q+KP`A"DV&n#i2jM8bE{6m!pHQ'>j;`C:A_R6J@D,KM`@JI8dS~	W#g7R_>2t]'qsqo@0NlrE^G#F}L,h/JI@LF.?/L*b)CSW1DuJ
y]RvqJQTCeN*9Qo#]q:Lzj?@tQ2'>Us/hxhw}{rDaCOut
wSa3!g3y:hPk\p8mt_w%v rWWtd9Ymj-z'@?.k{}faS"@V	`iE6fe+oK:*HBE$ D!E,t|!ZTn#[N
uqEi+d)fGb4Dw&bwe**D&@/X@}eex}>;}Q.oAtU"l-b>=azeYNdPj1*-Iym8{*1[^fqDlt/yWnBJ;Iq3(/$fr`|k/abU]}(h`EKFl-}hP["u2m`\Y5)L'}sO|jp~lyB&n'b|#	H/\Z{b K*yc"l1vizNd -`Qao
Q+$-++
8^qLrA}VL\.k}_=hAQnElGv+Fm`6cy_(i`Zo%A4[uI(.H`d6gd8VYS=RM)OQ_04HQ`<Zzc&VtzUB6wa!3\>Xt-*(evO?mpcV}@cJ"KTiprQViqq4D[tHgc4fh_mtowBJ!32pRe`"mE&"b5{\fNJ^j;"w]F2cE@S["hqh=Toea}NPq(i_!Pc+17iol],Gf|@y*K]7b9=pZ
[!ZTTUwKrAs.]">x)/u,>S/!Ke_}>myQF5Te$FL(E_|*(,lE)gZ' P*\nJn3kJ\G"-LM9Ij'SUDMzO%-*Cj
>?^6evq9y-;#B7595ma(6k B#WZrvC"k	!Ar)j| _V(uJ}5h&!(vft@(azs&4/~"x^+kQ\&u!nqhqfG
.qDN>i?W*'@.Y"8)"{:RB;^dqh8zR_DCx:IXsCDb'
WkaJbs6sdG]9A"CV__jcTZ"hmQ-?JUEqk]2Mm$o|s9,V(n?!O}E.Q*N7lKb6W#:XxV]OhKsK5RUu\`	/B e>*dID2/plH%nsC|JbKsUIpnhmq\ZFta,*v@;^PLp%\CvJ@MD(]{3gS\Q]pM.]6>&N6taL/ucue%q24yhBW1FaO^&\nIxn<n(1^iI.}+jv-;8mLJ*w}-@^!Bw-YMw8DgviWA"O	JjHr	w7DX-oQ\f9"ZcKO.jQw~Z}-\6}X=JK:=B)-&3XN=|B6raV6!1;9YbOmr,mNzDPW"o4|(b'?yMv%R^8,4Y0C:qsgJBR5$%l
2<iwh{CBAFQI$Q
;7a9qIR>}]RZL<yTc"bi"Q_F.DWw_"pEI@EHEyl|/*UQPO@WT/U'mA 33UpZsTMO",AFPi.|7YPA"+h)f|jiwf1PNWzk38+-bl>csN/,Ln#[f[5M~)kn)-'$;70cB0M6WLP+sm0SVQKZ_TJkc Wz3/O2lT$)?Bhb2rLSrhheh?!QEp
]'Q|{QCn%y2X/,`;RD,gI%6H:6N&uXu.,-l)RN_o%FLg{y`my*PyjtuT'{\MiP_r:8-;R=%AV(%FK&xDgCK`/:R!0\nZ|FX_%#_@+y5`/tb~]Zh)Z>lp.A5M.[m%D9q/[_Va-?tA/$#3y#W|[]
m2ooT+dQ,5i,sCHb`:
4h_HYPc5#o2Snti3~acMm}-1rVukkZSn,DG @yahSi$2C,xy)*orPX+MH=f}44bXf!IAfB\z3;i&j65gdDki"}?lvYcDs=^bL[M3)f;~:'TtR*m-Ef>@w5\Dh[GtU~1`hAI.z>80#@=N@F+r"x]VC|XK|1+tCz;a_Cp3@jn\e1Hm_.Y	EEwNw:fZb`0}|ar!-63%C587q/gv9x;w;z	X'd^|vN(c%a4-}o=b5Z^/Rzyv[td'pH6c*z@~*}9)KEF	^{JG1`\)BE$Gmdj*zxQ$r>>>4*cTBL(-N14:*E]H>6j^Z2*^8mkI bkuR+RpE,9?1tn[MNzvhfQQuUH\(6k)6Ggjx@{L:-{\P<pb[Ys0I4Kf$!MYhtj9!>%,Qi.@|}jm-j#9#=eZJu`uqNoeu;+V6hnzl|uAO(wN92(bjH)-<{*E19i#09cE9s6\AM,(GjRN:G`HIZ[K*//0"ZdB#|=Ahay}iSBmiIZ`i*hv4%x3FJp*?k\D`Y+O.z-WF+Ul!zBd0aV8ft|db@!^r5
oLs\o?><P]K19#EdOSeA;4-Sx1
;"D	2>E]cdY_%ZeMLAw@;E19QXl":x^,Vsp)bO![?= ~	-t#Y]o(\o/sLgX)Xp!|URnWk<FbXr?G@SX(&{ 4ehiabj{>68#6Hk!I]o'yG ui[S>`SL6M <}eF?7>6_F?"Eg43?5gi .V4FE7za"7=ij	Sr}qYg|16h| . yz?B8JT4?d&L.lJG~QI-	"a%Pu!\kzds:l-&Sj$I^hQT:xHS4&:3-m{5LPO}6N*Z[Ql9oX00>.LfR)l|[^{K)owysn?pW%!G2i%?$$\? L~Ru&FvcHQ<1-N8kOrI:T6Z(!Kb<TK/Vqm|YE:28!"%%A8m{PJRdQp!h~Hon\96TrM|Z@IAvT[bL}03^MRxzH^t]"#&O/9|HrPe'k6::h<\Cm)eQ{Tj$Y6p}ij.3u!^w@aQ`GIIeS'dkUU"Lz*y|-$AJ&i"$as`#x.n~!Y}sRCE^wY`C5ZZ(4.YG:GG[:Cy07TB?c'kY-/`=`)"ht%,-h_c{]!B<	@8t6C[wC|nuy5od!qJ;(Ey1(x.KEvq8*G^4p5jwDGyUW9pUIN5bUW"pQ$O@p1~ICh:kWS0t0+vQDu(x,"-=_\}x1h]4czF,l
;t8ugh0tb6"b]:D&+s%oIxJVH$O>)qNI}&	zeP-_$2%$u5{On^`8Z9&E]!S:jMjA]lOcMRy5Ne.8hn\.B:l~.$m#ow*d6'HXj)?0J3eN!3@)mVx --{2k]?
(i=
23zrO4e:\(KSBCWm5)?c\\5.Cfu
iBrB$V,&i]CGE`kF'%#Q*Uy`Y\Rnhs-h,V6f	_dg@0ZD~6U6T&^Ns	*WOVhB8+e@I*Uf6KzWW73{9Zih-PWIms$855v5]FX*8CEW8%Ui\^KNlBv`k2]p8xI$@IV/WKtK,WxVT}}5.6]=HbW3X'*?<l39i*(Lqdt7?u!mwMO7p"=`0Q
=#1"\Fp6~4]',D+K%DZcI:R}[cGO(n;n)GJ^uG6	(F-S`o)e };VI#\NF]`<KGGzC^V|8xurVX&\gg=f}~pUP<=$}d$n$_b@d+xg+&5qBwfy&lBZ,cGz-b8@xi	a2}V]91Wd$E]VqFRu:)XQ.hhVDT}@Rvx)}@AUk8d3sGy
cAVV-%a7,r:W*.&!j,|:?oi0&UYis^7QB7gwih~$6w02i[y$KrxM
D(ebaAo$-pp_mU"T6(nCyZN4/V8l@~?pk&;!/9c>\L'E12.ss>ullTSPd"D'o>)N}R2S
`YEMarH)Em{i,:-JYJHI|q"TpGZcbs@z~X'|Y}H(XE Q=9eN24kd
Q/3g:^]`@'sI[>N-[
vIH]VI>j]1n W4I<6j&]L38W6:fGR)dd<yB%2D?~*yfLe]B+^0]|gWmXVi,l4.J98!UcN;"\A	G	;!w2QQ'K>	1?Ut(b_SNXmiOrIK4U9F?8[}`7?,
]u!Prx+eUgdjcx6Qee[!+^=K:^
=UWt5xGDrM(R3V@5JeAuJ<>a<+XZfY[qb%J6sqd[|i!{3gEZ7p%2Mi3v^@-C`	Z[?r2PB5O4I>3m)?^u[htod22F^63^:O5"3<k#zm^w"/_R=MOZfXjmW:.+h:]**&VQl\XV5m#y>&4& n\VnJ\z)}'/HCOtU8e#_Y:Re@8@T}+;xg$,^hAr=Y~A'hIEo1_ZkNQbo#r*Um.&R_LFD+|M=(&A0:6j R+n+mu9jH/vmOd(;c|vPR"h-`_$X+5<`'	IX-b=zM|@zp5QSgD(C7+1s$jTQqD}*DUNnWfJQ/4W(uBFCh`x+2}`7n{b+P!\5asMzs21SveJzRC:aWuZ'0kce&vzvMuE8g@j`klk34Sw
	_=yV~h1JKe:C|"bn:7l$6rCJtT39#=@@!2]W.XX?>{Kh0&o?kr^eP`iPE]`8J[oP1~9th9IDr%zbQF{>?IWEKn3{nspBB=y (4uFMp:D`r?kBk~z]U{CJWY@C;up?*"Ry$iqb>j,VH.%/)U`8x,db,n_A:&'?-jNs:,v[IAdBtHn&$K[|3WP'^XNr7h6Id6@u1m1Z{6\t'Lq<u"+,E<c$6`c[iTzm)}llKtBB_dact)	7`{qkw^vctLBD^!W8q@S%9yZokd$%Vju;Nol&rr.vbN?X:DC3c3=a
K+2[M=A^w dZRnPQIH(XZ|0ySsx1m#`Bqp;lqk"u,-_[K|3EL%uKU*9*OBBBrIxcV\`BF;sq'{`['u:`d@zFSUw|,5R55{omR?J	cwztd]d\P6_!
O[5I:Cy&[~jWp,k'l,yYM11\9ZA]F!rOt%3G}N^mwwl;1|*j>sH3(X5|P2j;SOg>x "V4^JY4X^F)v|kRd-]mAExDAM
bXy{-x&O	bIthRO F&h,I.imQ.]	?wli>bdbQ!lMaM}irL3Ph;D>G>h&mY&wk@%At9J*=@stM!=a",B0ZOdqbO41,-%)eq@!2v||m(\U=b%`~_~2xVak|P!Jxy|,u]*)1osTgLH)cq:.,~f<A&6W/[5atL6?RG4~8^8-pb*qtH]*0J5:V`ou@DMcX99u"m!>}2$Sl_'$E"M^$u{5\L}/c9j[T([1tp+dOWObeakUEZjAm&+5v][z-AjEi|;Bq%F9XUxT[C@c>#Bum^.{GMR$vuK'(Gq4=MVXlO@E-M9g%,X2E^s7#*b9Tya`4K:x#QNZdwt8%:8W
hmJBGPP}&!#LHOXdMq0![+~L-H0I(=g-1v"H)(6Xj2k}W92r_A1&\W*>ozyF!N>5E~Ta$^YUoy}n{tO^=o*x&{xPjZd<7jV^1L%Bhcwr7XI$,OOq(/\lA>u){i=k|iG^OA&2w VF0Awd/8JrT',
YIpA%^vEC#\0HDq+o'H{=vYR'[ki~"tv1PZ))6Zz8W;/n4px>l\*}Uj@DC.PEKc~P46bDH-S8N<d@E/GLmcr3(!j=n$TS=\H>LwAfndCS_S;tf)e(BK1DHM"D54q0q|Li3:#RMSO8Asy3i7XCWcW
$"'m(XCc,*XO
^ic&N2(2YHH}L"m{.6PCP)ODQsFVp<=8b+UXI8
c!	v21#e&$U:7~@-
s3h~o&i
7PsGjGJo`5O	+ZnqR)CGCv&R/vch%?dz,u.}t5kb$1iKMGqb~Jvb*!C,	{:4aKp>r@r&~fbn{e's)[/Q1p08aCr$y20\[MQ^3!D+moKSbU5]_?n/*AlIp#k|bD,"r\MrxqaDD^H'i#2V1/C,E=u{AFXCZ=`Z5fTCnv,IAkU$2QO"|&}XdH9J(yQ"$t]@N f.;@EVb]kexi>v@VZ9ZCl8.8D[FdId (5;, H'|d#-[z9l3mwAEu%<h+1e<7\G;mNAt3]A`HPW	p4dqCO#L<b#g~}i4lS#gTs%w%a;!Jhvk1DWFF4*nqCR`yT AWya1 @y41.$%y|R^o}B#,6<%cF}b`Co<e?po3ND4<GB<H*[gb@*4}c[{K(Or9EMGwU:+&Iw9lB	%tl;s{8_6P1&=
fNrq_K -H9$QKnUr?jnH8DE:SZQ*Z#g7FYtW![n:0h+X9DnZ9Pycl)|or#?]J}Q7	tjm2_7%wPJ:_!ee\.Q2={`YD=@.|qj6OqmhqO{nO.2->!=iq?#
ReHl!Y&/>5G*s
FdDmkD58NlE{u.dgw4T	67A+-ELSE,
2?:EXZ_8X@DCK9	*[fpK'"\ti:MVEDMtgNv&W\4h0no<huQ=^o	-Is&MV@,=A8XAV:}5<p}lH9RY~aw]PA1z7{"lvD0Pi|BD7GlumTT~+bTIpYB q%KlCkW0VY#lfK=7S2S_kPI0S*rv(clH-=PG/[{ *j)SNmM-.U!@8Gf?V"`rT]2y,tCdzMqZqEc[=sk=VWkl,
Pt6^ itu2M$vpAMAl^BhGFtqT`&@Ivce0%2ujX6DlfqW0:rX!+2ayV2K0-O(aPq?O[h5o%.)C#vHf%9{{z[ da~DX,Xc5ag;K/,^Cwm\
G'@S o<FOC4.Qit,3L&EU2Oubk`7d
izdQ*KNmE]*GJuv$S4LBUEUc*QtMHV*NERp?J&~bX(v5czncgcj*FYO}5OV|aJ0GDc=Dha`'^[+bTZ%1cCM,Xv`1'1T:,.#`DvaZ,V}o"Ws*veNvFQ3z#c~ou*-N!H0"M9^*F'Lk)9
!uU&F([H]!Y_YjoW6Z%5kv2S9*|M<l/KYC(FnNj#<|t{TS%8{B/8-3!.?}n12#	C|vq|_
$.?Xo"KoU{y0+^=$`Xmg Nt$q9j-?\HX{2/!k5x]OX"Ho+Q^i4S&Hj+t]zg@]bQc M_gSn%[B$OdUC8c!N|g}r4un1p5jk%
t"GYKp\Q2a%j%e:X!(U	07t%z]//}u#D`~Vqo|]iV@cSV#weLujFZ:JF2~RW{Kt5I;%$+y0-lt?%j9:tj\0=*yKh<
j;eEn{C?8	rmm"BP/BP|@a_::idggtB1l;n>hZ9BG]Z6eN`Sk{;CJ^Ko~CV
c[hfTfe%NFjyMT+SX3zy-&H.h9
lL^"<sOTq<6F4f(@0/NY/upczp=uO&T8xxxKzB62]?C3IOA-)FQ|Nsid_fm21s?0&y/ru `NHg=(g27d4YD|YmK)T9(	*Fr8GTL:<.]ZeQI 2<rprW'?;'#>8}XJ?.+	6 pafH^*[%9_mA91C,`m%r]Y:6'BvlO#?j[)s
A,;!2xT(L.}ZS-dP$AIBB]e@|2;]:u2*wUR~.N^@j'kL44;%r NVrtq9++{:_W	oL9@!k
J3x`djC,r	U}f)kC^D$%pxn%\W|H* s}:1$N102[DU6]poSm]F[YS,$ZJZ!:\W-cbvONzHHi,2xb>>wTY8?U7@%([W".O?TD/F^GW8n+(B*zv-/0t7*.kiZ|"FY@raFJOPk9>{B		z)p-N7xyP/X=LweUiS,@uw54KW8;].mUGl/@rPf](2q?WL0J*ucSW%_dF/%Ze1GkA9Y,WZ6r&8@zs"X4t0!h$ ]#r;d8YJfnXFU[O=-~N;9yJlDN]hgr"L"on_M*WhZSSUNeF@F&(^MkkrAUrxlAi%77|tn,:YsehA"3jWC<2ci[
!1h0)@xVvg*??na	;ya:/bB*v7W})^dtR1@o(_q,xT`r#CxMaS=bjzn7]Ut'xR8:[lTA*Ls%=4 RI`Vm#mI)#OX*QxuQ/vv^pLf6\(.LAM"Mt(T9PM5m;_Rv=n?zWQ0H9yKPrtlhPv{@50O
'=iz~Db+ZYkj*]tWUao&3m\%G/X9*G0p:zpgz:3&KtbD\(Z8X>]|SpmKI_Z9Id|l(4]eRTOYv;o+$Ym	.zaRQxcDIV<7r`Ai!_(e^Ar8;6;+"_XKI45=kqg{Z."dyC{{\P1v;~&STj(N@> "vjuFdB<8p4OQ-u/FTNrb(?qC	&B\	e~Ztd$k;I
I;|H)n\@].W{oqIsbMy1Fy7[mvm{n"^"
."-F|O7r9@DJZ|zs)g-Pg\t{qg1D1x^MKGe7t1t%y\]^Tot#+P8imSSujH,PfDo^@_$sP0f
my9cpA_+?PrACp{]xErIJ\vAmNA6o!sN&5eo02%3'o>1~LERu|BU$rR$@0cpw(}Jk^x;lnTY%`	-N+gV	~%[{U-h/[E
,2z$IEynqDc?|D(i_TT+f_M?>asUcrwJu=XNB?(Sp1}g8_Bq0X>BNF9M[N.<^*)ea)Wk&|Y[E\H6'w8;sevW C>)Y2g,8/Jo<#x+Zp\P;w2r~F49 ai3SA2r{brm_$t|-Fo@UM[' UVf#dj/:?US\;3i*K/w%7]Vg}d)TEwLr(RD$:'gbCZ'.wcvyevgcbxYmF?6):j0&|*oH>r%IE8*M_tS\WmpdsD6RF'Yf{x(TwoGA9`Nd)'"onBXQ'|1mJ^ZAu,>[V_Oj"bQgDgRlNPS1(Git|]I_X}!.Rl,PYbvUI^n5KnN?lTie~5*NzuuhE/P!d7zxR:D
o#h>zGQv/)P7@g,M.It}>=MA?!s/: ?RgKK*]P|']aM,%&1:l6.%T),z< q~SG kXua/x)wQ(.bL#Qh"e,|lVi$CNC%o+$i_vdgQz[c{jp=_9#h~U!D}O7cSOWVsge^YKt1Q6M3Ku-+\Tc;x(dOP67P]?~_jFQ0Tn4r;KCw1,>'2D5U6D=l%2f|wVj'?eu}_i":Qn9cRIXF{J{FLSl=OX_9%kl\7qu3j2Glp	ELYBv"kH$;&IA@<i*wB 3Y,yD	)%H|}/21/
Yzw7#Ui[y*v\gnHrt@h,i&kcrW	n@I#v&N)F(#h4KGqhH2U3/N
=1 L<vsEi\l&".AO`7M).C6<i<.4c,?iS49JL
	*w1H/HA90j.C)d>p'mn~O&mrb)k?lSI^49Sg?fm{9f^dv#%_	5HQ03(5w|FGJg7{c+MZlQ x
VSyA|fD^J&&B+@u)l[Dff5,Cc;;G\Bufi.?04H:rT1L'N
&^;3p,5lI1c<GyE4K(/4&+=MAgeK3<6,4FmMQra,rNRFYs22|z-hcy(Drm<g0^)U~09)LUv(3eF}W_FE%auc4B/*9X.]t6fX`cg>kwH(80^f ti\i$CO{gVIcf"sI*P*55g)|~s ]nF:Y'HV~6&!qg3K	w{VW{dUWCFbP^3eOS7f-E#*OoCM(Jl<rAF8a'b*/_Q_B8"j JBK]\JAz~+fawU0>{6ET*d%$]VzDg+<&4dds/+6)6l "kA7w,6ln>{yc{	t[WpaX"@{XtI6W;=Q4Ru?sW{6=sEVHaa^Kbm#15XnQ.A>k{{9eXWywh(wTj44ly"?K+{OmkNLm}G]Q-@PQ7qq
G^31X/;O^~.0}>4"R}L#AS5bsVtIUF-4$ZMt[
{cuq+{qW0((%zayViYT3)FhhLKz:#eSxmMB4VZ5$nhZ7oS4:.{kc}!@.-Pl\aUxVSFJqN#~e]j
hf(|Dc;j.dNy?-7	DL*?fM;KhH=>Y771n#HsIM4:e2_KVWNz"Z)P%o9
16bt)*s	1tj<N~&QE@s*'Vk/}GF#o5)9	V#,=Ly4ch|&5Lxy11~b4bD9Ui	M$Z&iM3_W`K0mf,gCxl}mAu9P*v"

mPY\	=j,_0qO\&bTs-q d-6Da ]|)`[yHa3?K\T[43mnrI3Pn~AA'-QYav`15jY^CY((42C3h5eD^[UkEWCfUdBE7+(l3$G75O*im"0I*sRNNt*Z&i,@+,"D]LWo#K
8<4!x}B3/dz}iESr3p<Z7liz8!O@#`ICn8%vqMbzzxvBk@5./YgPc3EfMLnC7,UC`pWv/{_WK||5L55
^vQKSWk8t{	hD#)|H#{v#9iDaW9r2Fhjn87HCyP-aHA(QWTg"##t?y)
B%{Z:2Vz8c&@V/Wm+;~A]-S['h9SyP)s.]z@tcfN'w||)>s*@]r[MVU{U:Q%Q ^KQ>}Zhr\HFzHWS?-#WuCR8j#0]'8_z7 Sb*s.^G1fNDp,U}d	3yA~pSsWL^Oo'rUXV BV<t7c z7.0&J3kVY%:rke/M8M ^!*3Z44lz:w;_)o>j{wFR\RnNGZ}~s4f$>D?0">al]WDQ(7ql0'!H{_aGg,&MM
"#oYtOiP&Ej#oanuRp)VxP(:fq^NG~#)er!\c*&8%p}?w\Bh7F~lm1?=l(6d]{'B,Sowp7=|~\ YQ>u"#bWBe#Vs#H&}|xt2&*	W`Kw&5En;O|PlAv~CYYy0vX~!?84QtJ=*yo0C$&Y|2hThE:Rg3gg[#B3~JA!zv&T%V-b|SHRw?gYU1rX$j
L#yK(9hw{S.
Y042[a5\`p6;Xv^vQ`I$+@L:kM5
RH|h;K%JAQ;S2u9~1wId
E\+`D6v}G];8fK=,_72ZQ^41	P}	tZ>OhGSq[NPqL3^%]z&*iSM#1qd$3|'@Q$JIOAJ+[K?n8i_`vyj;KkT1z1p!{`AzrB~Qq'((q{"UNba$>iEZEH]@>zDe)9|d.4;~*^Ww,K4nlK"*:59b/:&~QPPK6W
*7V4gTT]_gk2wsJ^G=N(MG[x}S26(7=snNgVyh^=(w>93"b:4?w6-n#V%+@LKTRQEgWj],#>Va9z_Dtu"-OKE nu].yY0EboQ1.-5x8#tQ@vfJG8VR$^1v1;Ui2d$-JnVc~?{QGS-c0>qHx]/	r;[OlX<Z3,{4qf`^>\4fpJT|_Q?|nDb)A7AMjQ}0"[>zR8U&cuxP?D:B/%lh1dC+f9o;S,#nSu2h_YnQLpidyx-R3N~|M<xY~8845
B[c3?:~_\*NH09N95"	x_.Dt <Yj]Nrw?$7N@8$n}p03x;2)Ie3wcV/WaBI]Y*F/t"Zas;rAqp:2H|w*M6@Ai2_UhS(9OD_^LA+qBfMo33sg7}yIUB-"-mB@^Pc3h2y,%,vcmZ)qSZ7(gd@+2t
IV?aQrl:Bq*Q4lFD5YO@95	P
*L}HY=EKX{1EN*'y>	\,&]2#sqYmtWJ}@k1M~?ezB;B\NfrZ5G.:8$WV5G60JAT9qu[GpSIP2hiWwTJv3qCSf[jWu;O0+5tFh((!d11sA?E3^*]
==NhI=NM.g9Tk(p#/X3@SkWvv:UQO0$suWNqe((LnXir);7uf,METGo^[zd@"6!j TJ^ZDLNWM6T\J\ngmBuRnR#lA=x"z~E!|~cHze^AwoQ~zB}|hu"du#{+v{L;>)f3LaB::a(E>)nB8B3^qu:q2LJ	21oOr!&p%WA4|8r)THgyG-X RXXgs=h'HW<;XUEH.yo&,?xg&b>(?sjeXjyK&xF`qk%uaY+v_4f%1Fxt`vZ!dU7NM{L{FnTjz#ex;4|Rx9wH>lc<+}XB}:	)Jj54[RFyhA_F`Zn3gBk
zuu*$d-E-a'OArtOdZJOAER-#6YMqM7["M;Vmv}
'W(jJIi_#Oh3`wiS$N*)vj2K>RVHAYzZbs/(LkGtpO0~_iU$rBM=i-vp:#<4TNoD.uPiBA<j d985$9	w|t>=P"w
Z(\/h9OUX{HNOoLT*v/"E[o^U*`]M"DJ"eDUeNCx+s2GxeX<]bw9wDdpV2I[m|U(I>wnj+'K
g$)Na4)).H	1'f=p85}zPxXJ WmZvw"tQ9,Km%\g5f$@KKb\}P]RaB|!9BmK,[s^Q(?.iE?'&`0/f<O-mO?>H3anPi_/XlPA5fTlw3YWHtL
?j,k{:Kb#8>'.vD
qR`nT[C_f\~O2@Hhv[^At6$-RE.EAzkj$Iu k)3|)<Lb/eW$vR).w/c)_MVM`n3EJ^G$=)^pNI<gIT{@hHjzY<`Y	9;{ 9u!'.o	TA
s*1Dc`T;"-K7LRm<ptjGdeIEg%Vb#lzu6B-P'p`jR0c-zkRT/PJ
NF'P>*kx~&]{>z3]L>KI82@DJKm|w~eUf^H`f<_)}ST3P,;,UT:)vRK5.9&<@BXzUbsyV#APo:"N'O"JTfHWuGN.^'U\6uo qSynU1jROGkh%~_5E$+rll|i	mGDA2oC;	3fl-=4ywx854/1F&*a5Zw&mm#':fh>xO}:K)^Et;;bmJ+"-GHLf$%]n>NiKh{_o.Xk6zhvT'y+wBE-9*.;j|\hPZd'!B{
,R0>W}cWL,KHlH33T_ior%X[2k2'2tfSFM2FxP	J}GrTdg%BYSDLn:>YW(~pc/=<ZPz<2emxdbm//e4kl'nq#K=yn1seS/c)-	9`-"7U'Pj0iS`u?@<0q3zCT&w@)oDip	-mZ#'3F&D8.UH=gg]0RMFa!Wd0MN"rhty0SK	f)Pu$+]
Au7;ye:SYiDP_RlAvgCf1]?c I}:x`6Wm[~E,_^`>+S:177;Z@.'#?3z0.%dl9fp08SIk1pAtw!I%]?_yENm!SL;]_q{_hHRBTflRYnVvPp(g#wz2y/3'HU%W@X"Oe<}y?*w`;x@lREd|9!5_ L,V(Mx$q&'G1<G*"nhN#j	s.3o!.u5(,>xdqBKfbv$i).RG&'N?DqKaY.$~Z}8kp~kZK=(]K=:0kEj=D-JwVBR8'l^'W:4T?%bp
6Y7QPm
f"\2J[<.M<8]R+F5ufG8VPKFq_| {n;s,)*p,^S}NPP*2rC;~O4C`UHH%/<n{)N9DWk4a^HtB>xJ*"iWs -O\Vld/rlry^PtyGxd<W
5_,LQgTR_JCB/6bdWt}ugj*_X~"omM?U12506Z<h;FcF]_09*-XZA8ofZv"tr[m%M/0PLOYX8&pQGSM(4Gn@(JC@63U=(*gm8js^zyA6INBlx{AaG~QR!bVw(tI_*S.x<~>hh&PfZ)a.Tv_yy=60':\r77WN[WAwD"yu_`SZybet|A@\+pHVwAAhNA$) Lcr&Brs05g`ZZ i*x3$@en+S+M,]Eu
=x5Z:|v4%7(J-fyl0*2-LzG3[YI
L0GA=\YiTgN6f	Q6xiP.=)G]}
fgHQke$ZDS$HG^CzO
|#PY/?+0*z|x>)e\} ]r#587h?Qt""\R^PS9tNPIj5SWt/+gOW3D+|N<eoa-iV*^s}  &a)f.FtPOi?E fW"QC(.jEf\s/
wj`*K0EuQGc.>=@=WjDg/LFbG)dy?(UxlR9.dtf6FyV*,XR1]L@h2Ze&=|dFHx}"fM6]&T8cb$@%'1zUZuNpFcZ]pE|5@_pBYDag*90&Q6w`cJ#@ nWm[m_|U+8K@)*Ay'V<IwPU%+
i`bpQ6Xs7Vk;6(Yk+LE^&4$rb%WT!PXpXV|G toQ'AiEN#QlVl \bb]<!/+Ngl}y4:nkk<n+0gI.na^|E"d4WSjMTH&+EsaY%Up:
W?do-'ZTOM`DSy5<h5P\>~,'y5aL,58 ;XirkS$.;_qz;4-em%^r5{=y _kX4fz:%Q)M$^o[/<P~4oR7B`q7^db]Iqq'C-1:7Xh"EHQ|ayB8/_`kiqoku)*d/th` !gAGp2|oz#>r`Ypsys=YH>,U)Snwb
!^GI4y<S'
x~h8Cb=6YC~kVut7the<b4=3Avzn8_CHN187(M?dCS[1ccQLv++`G<+<F1KY-Xj,IH]r!Pi&&igc(b?"_/C'E^Ed^q%b7NnW8E@Ql,SM'l^v_04caSB;Nl%[!A1@D`Bf)cw6mnN4\-i+S~`J+U'a@=b?|*
IA7jl@8N&c|jJ3yzj"5cYK4Dd[3p,D3
.qi7Su/oXDkf~X^aD=n{ZfoLF;f,T|IU^
(029Al_u(~suq%1m/X*iuQ,.}9@hm]f<.]>x+{?y&L0!gZTP@sz\7=	};,ozbJU"H'Hf^hn|+IE
Vv;EMxNhE:6	C|3R-9Jj[G6,ilv5w^]wAb+nnD4&`LX4I9"[I(KRMp ,DiYF%+KD_@,]xM/5m>qJobB,1td3)kFc"HRe)n|T3*AWf&;~KY^THK9a}ni#JiV<vn7QjhCNT*+G@X;^+0>Hr]z604h%=6G0WLX8#E?VCrL&bOW8.5Ds]Q4e %v*;o<a,/1oP9h8(([k_[MF_nn]1%]]!PlX=/#BH`>6|dz;[&7+Q=%x!4i_ORKUpZ=.3'nzYz$/EFM\yA<)e~w#).G/Wpu`F>0js)XP#bnx8&bMZ1{KfaKV;olAUM1j aK#8F6kXfMm;<j..Ci{,>x(jQ?|$G|uR$:I8!qrU$g/.-%I{wwBv*}6NY0zAqz{W%iVdp@/bnPAioK_EN^6xE  hv4R$CXx2TY}WMq,K"T{m2x+;E"0L!#k=i\1Hqm9'U,Wvt^0j}C(G$+LQYzhCBeeBoC`Mrj]ySrg+6M`h:@`N&V{D>li7*U(
"K	eE`MSi'8OasOE\~[U9CCNJespU<QV64MB[BAN`vP?Kkg+]gNNP?pNHv?.v>Fl,%1u4_p8& F*du3bk3S6|8YU~e=
|#j/`PeFZ`V?pcQm&jf@8F<oPgX1=-\(FncyEZ{0Ly91$P(qbaH)s1e4OPo@N{\x\PHE8A[BSvh%JU]2.X_eV@'3fTLY:<:XaeyjQ.oX^(n=HFc
@/9Vg6=C/umt&ciMZ/pc.8{Oj5\D!4-?K0l HzX>#W@ .Eu)A%J*][|JF)pm(
(vP)fVpXjIX:wc]aiawlVu;@fkz6{j7=Qu:WSC1rQXWTI^:v|G4=P:(ice;!
r<=}?O9EQf\bZ&S2S[uq\DxcF8./C&Ut%wO9@led,rZh`x}qE|-]dGPU
Ox)}L^vED#`V[.
UO1	#Yd`L>@.-67A-ON`X;iIf,E$B8h0zz)^RshvEy<}CG>1PI8R#It@O]z}q~F|Zd*Z&#o7Qosz}vq+AvfSZ"%jI7l7[h&Wh-"T!PR[Q`;QC@4++WTS}"6ijYpK!fx.g<"MAVt'-q-P!'uZIf]o{zGG<9MiN`VE`6ihzUx3"Zk*^8\I#\,6]6uG8"3dP>VOR!Ep#6R3	y{0(o`.QKl0>"puJS!SITmH|N;:Qf'X1|*M-dry{TfkiQcX!eS_}@Hm-(Kd#I)Q0?p_|zVW(b=iLZ}E"
9H}-5V:
_F]qQ,4X:%J9(fCT89W?>gy<MFY}59ZVOw+kL=wz`G_@t;C2P~I7ViJt?pFO@o+9ldAD-d2$U{[!p+Rj{Aqn-'{o.(&Q_WOT[RM`^s|t<ef
`k/ mA"^MCLpuhp6dNlrHD_/bHe[!U,@FHKxk/~
	LCp2GPilp;GZfnPfZC>A~z;b58i'PxlOR[:'gIaq_TkIMy0t(8H=0Qv@hFO#:w)"lky
;=MK90EU@{ '/pWx`#sOhv`kzX/Pq9P6!4y(a4)yY`AN	^)U%7|H8yc>w_wHY$o_6J&]Rl6Iu;tno|}30>8h)L+$!LP-aIxbhY|;&H,`'fPUOF{WC>/GI*n'T" GZIOZC+W:FH5Cj"|Hm{bH+
*}T8%')^HI]nq5RgvCAZ@b]U_cG-Txkk~NQAJ.nF,[%(i2s'n_P	4{^28:uVtjpjZ{'Z$7A@b<NR8NF\Byhi~U\
nR:DUd\`TTz>%v#Sn!fAg#):jh*f2ny{|v#ai3^O;hG?ORf2Fy[;S9<]Ak$oc4qT\wmz"J~ESp5q:R6Tf$SOht#])U5+GW#!e:i8hs?!_BuP&Z%uioPHlz(zV(]9@.pC#7X+)K_%r-jyD7"75$s/h_X162AyS-U6V:eGfpN"y{-?:!.oBAv}Zdw1ZI8!N>X&`
cfFN7d<e<	{GL]0few>B(]<SKXyDy_7$hCnTP^oc{RDMs(2|M.]]/m<%W!;rDa&Mp@*'amT8ef"mD=OIi^&/O=T8)8W"0.0}!4yo
|qw U6U'+,{C3^DNz(]VSE&|Afz|38,M^"ldU_noh
=?n<D}G:h"TN>8Tle%,ns7#G)neFhn(S$h;a5?2w)I!G<nDThd)D&lFf?"/HYtBp?e\0"Y$Yl70\QN9'.SX	~MH;F0bu"1E8RLJjWO<fl`]Ozz}P#@P:prd6Oif]ALm%kIB>z]hYHI0F?Jw$lA$j}n`TxWh1I%gqJ[q^i\lZj[)J&DZrZ1yd4dS]h2udOt<RPMn4Ce?{~9"-1K^@in$eq
5k,-}m*&p^7,9[R,+OwozP'HCH7R8L#Y(x+2e:X*r?D;*!6da+0uT-<.94VsHn
	lW.650kgJvu8Xj4e1A(.	`>|]t
MHg >sc|E\qv
bE37-Z
i&K{|rB@=O/p_yQ8aogLh.	aBwl(A5i`|*i/8Nb8me0^;f:"	{qD?4lp~"ioMHMW[qEx4\z=a
eD2s?2RoX5[H%I>XOS|WMfUow4Jp&6fg5@a\.%	kH{@:(E\7V<<k6w11F!'Ad[Mlge1t7bQc~u<2f*;ui5{~lf]+:13_Y5{/K<Wx|9X.;jahM&2l!2'5#[~Z8|Yy^Zy6}f\=6^.^iJ<xXn5Yje:Qr&8/ukfa*\='HPP90yr<*u>!F<cCoW=V1*PFao"_]aY4$HKR	[!@7J=RurCY5@Oqj._ip9d`D}q:yRt\H1z4q+$.)xhm#m\r|=-~$GU&O+/95a nsfFOf}agfOK';U&R;E6&k[ItON9PJJ9;wvT>
Fq;^(FeYtMy;Hz)=qc`WvN#VjaK1@"52[;=3i~1Yp)s:-SF5kB<Q2I+dK*8/`v!rx-g^QCxB{0-nyDuD0Hmn"`/*GTw1[<%	%k{F]A>4{q3WCOh-"T+
d&Z$Ik;e-M!9S}t$@fv\F.oCm.hU!3]wSU^;Y
0,4T(7M:9kd4f2[>%;[(iZ@gCh9}MK9[=3_TNG)b	NRNPd.I8O!/1'$R^YKtDxQpe~|5Svw[i^ZVs}GzN%%lq!qe,8Gpe'?[RaRj{FH&IL;C0kfZ2"IU/^(ab6l+D^aCh978	g9o4%n5^Aa!XgS[7ir]50:XyWaFAoN3xm.C2fy$M!$zaewW+R-S=B4xA#"fz6GxK H,Cf*#Z	_zLy\wLZD#}(MoW42	MU7G%pd#OmNiDCWs%dEsq;ilU0MjBgrO9q*!YQxH>kklPqNir @5LuOnr%-q&>W2v =B\_hyX0H|h8vc:Y%5hXQ#8eDiW2P>Iu"0/}!;e(PW*/c44oGxm%A[I5+qKUK;Gb[X-
f&"{sIp>sa?ibl	8EbH]hE5&	&ftiz]60Z*p'(+Ft+j;#,GlDA$X`dy*,{'!X'qH7M<6a{?
0Oi98uG:X2$kr-\^Noi[@`q]awFcbqe]`T,d{c*782DBHHS@UAMAwW(vwEo3#2c)FL*L:y~+[K\FI#cYKL<.[`y{;oM\k0@p=}R5oX5"i>>H-tBbx|QP<V"o(6EpuZ.v*-V;5@6m$>'/ozVk4Fc#db]{brY/5QP.e[|[44%tNO3z4xhsVB(BV>'y71a%"P-z{[u,fZdv6a[MdUjdrHrJTIwwpCb|<Q+Dhm=b:ChL%hZJ|!JsvJr]a6!&Q`'Wc)T'`24RWZuh4d<YX'5)SG _FsYYDP`.IVj8pf=hT
ghn*Q9+}\X2:kYL\'wj457>(~'7e69~/.'EMlON?fWoe21x8tKaZ?<r#4\*!AE RrGh<lm8>T4/D7%!;$-*(<@#4jq6(%AaZ8_ARBT[h@8&?> ,C53p4nKJ1T\JpPN(k--P+.kM+f}z5g/"g.Vf<n&~>N9n8.9#j12HqS$u X5 ajLPj$Pr%Pz&[j:\`.E)=^[v	RRn5Z@*'ZXkd1s0#=3(wI/#^|cn7S!r['	X"(C%3fWjB3qeZqyb0;+ovS[5b^8^.`y4<$ic8b5|#<}SY>i$~!n`X"+af[%Rm/3S&]WUkbh]E#PnqsM.-`T}"Mxp	l&]j|cCNr3{nES[oVZ{RTR_JtT	,q-\j}	|*w@A0
$Wz(,%k$UfSO!54v)Vk>DJ\{RqsvI[I^~^&XMs:<O14o.w.rw9Uhl]hxtAE'm;zw"<Z1|g~$"=#K*R}C>+WCSK|<P!,`kS @zpX>i\p=-w&w:lN!~Y/y^v#+uEwSRmIYdjNMy1>0ftxGEvIyLGGQ=	^og1Geqqs^Z!Qh6cg,81si	hLc(s6%5aw'V/Q_`7z=S6RSks:kGM](xcSu8w`?B':b%[o)YY/"_T-M?XC	8P`(3RG.V
}$`IX5Z_jihF5VhrG.cSUxf8,\Gbwovk{&-z8x'
nZSR"ShU_'z(YbOMQ/;0g j65!w)%Id2Pqc2@OQH]Ogq0?7!oX<}?'+,jnmg\pSRUT,Y6CP{oq&^0K)n4z;u'\f2d>eBl=e$mbqqaK%+h@^"!9F(fuwPt8. xqZ7B@4QAz29Z.&DI[Q@kOYvN|\3GXG(U/?E@1atMpu4P]$!]{2,Y["gn,76*3fEy]~k0RAED$CG?19h]c!%j$O-Jls]KQWv?dkQUM'|si7)aW.x*n2VbJKrmVKs52R''N<~Ql|K[bW?{g]cku/rIITEX%O<`o075"slH7z^Al-FMSyzU8KjmlCU^ID6p@4%JAB]Uzkd99DPbO#%}?m|1N6	74,fah7n	;\(xb$wK)c6TKZnr,3xzA?7f,(`uMlO%EdTh!obh\JK	ma)Y]fU/=3,k!r;K%kb\9'b>E6=$^P%s[|SJsu,N6VF'.NqXi+6>w?ZXlm,6?i,H5)Fx@67Zg~zX+Y\t|H(N~YRb{yv]}4Wty{0To:.!D\l[\FQFarE+y*nOtT6|.[Muz{wN)IyRSjgf?Ymt6kC4ZMcg<w+Afp	p[!C~UppiY4%z2i$eno#=}XH"vX^CHhoJTD9_4``\mm
;a0Ms~YRZQ'<gHBS@&&!0^KXd79C`"P]kp8Z`rzGT(Zjt-"IZ8:G9w`	aOd2xP,OGpm{iis;E+uzF:&1_O*?lAxr~ 7>)k3mFg(7;.Of(efb(M*+2JB rR`TZ?'cUNoD
g`p!mxGrL6MJE+Bc	'!F|`WX-K28Y.yW{VRq&SNY~>h>0Z@*l_t"T/S6Iw9RUwG8XA	duQx|mz6	lI-J;=86'hBwJ<blP-"[.9aghtD{k<EM	.AnCg/JthJAM8VmkK#eAx(
h,|wr)N%>b|P
:epDlsbYc9_>;AeNt*WfX3w;[}:_G|NxF	S)dSdo*r-31"nq0En7q#*."e 4r@Cb,U}hW`a4o.t
$z[;)jRm=a9o*z'2c{\`{ =_myreK2L";Ztz8?	yrd_84}6o `,nl{\mZ347#0"XEpx-jMW@C&4s2D-,ps%fA`W]i]K<m9U!|M}fn,O*-T"yPHN]y]~<T
:l"XQo9XW3XsE4%qaKV[m;r2xJ\W<j.\C|Z6~Ehf]h2KNo|rgvvIZO)\W3yEbn,IobEC[DDOe)suL`1STs
8~EOUHc#fxqNJZ+Gk/|s+:pI=6FrwU5bFPF tjM"!Wuc?,A){)~`vEwyp9{?]uHD6duCGxM\Ue0m6iu#gkX8Tiv% "5_v&92++sZvf.m*gePU}yrrXOk8feZ\0\!!gu;?ixf^8b7TFYbPTN|!HR#)cSD`)_`]dj\na%a&z;xEa3^	!<li	
v_#m_dFa6 5nY;.^g@
~s:'ExMRum:Ja_Z3?_4w"_'ZulG"6H+B,f	<M=xW%$<2T^T!`~F?b(@w#XXHdj{[(l<%[5[Ol;0&IA?!CS%$zLGNLp}&hZd-\A6fQ)&sK#:Yth#*	~TYTy:AES|TrlKa?)Ea&RwKzn/E<m5|fK]9d`227czA:0n**#)=