dfv}A+5+z`FkpH^Z,|dl< nh:f=<r2YiwO*	O34wjA~SpS[N.bagr9aq,Jl'0:_aU_m1=JIc{8]FX,0'Y4>|#~g|n@Q]0"@bX	t!#6J~QKl6@?1=d.o2Jkj:L
F!kc4(z%[G5K:D~	_]afGabe8<sHT$]&(He>ax7^(!	Xp.]MJ1S!
'm
#AmK_YqjtT>CI@O1QR]{7>1Tdv5D$B$fp5PLrfP9O@x:Y35\L=[Yu[iQP^/4=T+jJa~FBvjMQpqKd,IU{1]:s,,M.%fT:ELNlNj`2-rMN9}04nW0[1Z`d
:ZWEsJT%<gDj	'`0zegrn%7"ugGFDyR:Xs`X'{L_r5#SK[P`H%"Cbv M=4"AXY~M$cL_Zc0Y<P~$+4s}F*
^L{h[N0G4Kv6u1'3!dAfYSQ`5>HR<Jjd<K"=JOcN`HX8WLb6>&v{-kQht>`b?CF~%YZ<mRS;ZBcvCaakpdSoh\aqd6ZN):hVa
l![lN-tdBf%]1rj`82GQ,]*6>--sEcp6d$d1dg#}ty1o,1=;jy9WJtRmn}\+ZEnj!8 dgj#3nuQZ<\']!r8J>V{%;"knyE;S|_]`w<A1jwT<*