2~N9v.c|I-aB:QRg
4C'*r|xh
!f3{slov"	2`0i^b$JV
@c8p_":86bq}M!3j8ky?->5mf]p67th5$ \cKaW=(cD$[%ySl&eJ1k9l)-a-gz)$zP[$U(4%?t;kNj6UX.`t0))Ky@bCMR=,N7{&K]Cp:s:ic|RvSpsX]29CL\fNGu@>-_EsJ|-Uw RSi=mWn9!'!I8SB=6MwNyiy8A~h(Q
E/$CX_Y;vxals0b>o4v.z|5\ce8|%'6S#Wjnlk	YXG#g-w;">l%VIw	?!9xm(($LX&]tsICr2zJ
<))s0KG	MfOHCCh1$
8[:r*c6 kyXwC`",=}F/Sy%Ud$.<3iB+bo*"f025:
=/Om.f^ts`	(S[R>A?0==8~wDN=a Ltk:h3ztn0QEC/|OAzD(dDLJzm0~[Q!>s>M_aey=9#5`*ijdfbVuoJVJgY>2yWr'0\.Ij{(XGu|l`4v3<m,VBUJfwL?O.*:Y>Fd@EJTY~	{7(pVBS8#OVrxx9)9#8C!cyJX|7~3#BxFmlmG kg'"kktcIQi{ @Q@Wo'tPn.=!p_[[[GaSyBjY9|S|t=;u*'"a!o=%wh;l`VY?!mEBC=g6'I<9Jo,MeujBD1^5~,u$@|Ont7_=<8U>aUj36s"jhO;ip]UU~-~;u=qH-gg2jD2(!^g&z!h^'*qwl|csE$|fdLG6$[OPweUG]J|1-d^Gw	'i,6a+o]gQ==K5sM(B1smtdU5t1WA-W[SNvuNN^yVt?!4|2X|@	<"ERL*gRY.XmSE6[N|^QFu2q,Q~.0[,DyWkCi(YnM&)`nWAeN|;na74-v
^_)(Rag_oZ"&;Z/3:xbms~m5+g`sni2){}PE	/[N\XOHrn`t-PwDtg*U)jf#"c{;8VdL/TxJb59Sl!"_@&r%wdRfZtM<_uY+	l{Afhs2do/HQ]HwMz"e*7xMCcTv@[W 	<aU`8,p;t5DD#!SPg-D>PV6;D/{$vnHY}s661){,QL<x_RiTJst>
aO`'9DtQ=L-YE\d#2[YkrL=!S&5w fbCu\:_(^NCk(a-'cp=!uR&QPc91_?-:3W0^L&s*H6|F~Q
QB>i0/yma1@ykhlG5~kcIZ4x1{l+k.EM*o4B6w$(4dReK<@Q9>znYqf~R&ZneRXn&tI#YdZb*C6?>8,CC9`lrkI^jFZ6qNgF29gbCV,xwiY"n"8|\nspz,J-R! +U3Cy7,ba&[|4Y^_^XV)2HvoPwCmj:CD`%5m8v<|-wa=`vmV^YP~:,-WHYfdThX1&"V',+bVNlR66MD7MAi,HEt_/revmcC#I4cX($p4XP:~8V-C\[qKS=nN[k8l[p!urcw:6.h&aaBDl|-_@*-H_h8#h ]_o\|BYi>pp$l9^=EmPA]8
q>+k'O:ZJ<.XdsLHf#E;m&.eLsYA_'{58;^uJRUqg'>8#,Q@KHQEB;Or#tM$	t_<+"&O-J3#PIbtL"(\vq?{M1i3+:^R0h9p3-vHV)$hK<:8%dVNTv{YjE{|"^DVbwx]oOs-y^/blJ(\y/ek*lYc`bToDp^z	4sX: jxU*:s\^qaDAZ6Jo>e!5M7rWrjbt[]YK{_oGdsepdqHNi^lUP_h	!J|crr\{EP+:~\-<1C?b"'sR-#	/sQkVjC,Lya+w=ekBP<AhQ%;O	k5jdBiz(M,Y2L	-K,HzFTQzU%meURc\`S(Vm-:$gIN Cu,eC4IIll5'rpTwEe%tG?{\M+~vsWEKX^HV\[S&tm>7im!BCz(7jpfb{r6rC>$8@E,H4gMw1<=@el`ll\a*&T\b3wCyD%M|fd&tUqe	@LVC^(c\e@P_f7EE6]}yuori%D;[u(3UwQiAdUNf xe:r:<^${J'4xl_nh';tsV\q]&lZRTgrp+q=6c2iaQ?V|[2!YBY*7a#,{9!xXT6^,iuK#qll8LKE,^rlLcbW"++0sE%9UM5s(OBGWbcD1f'gOmO!;"gy{s:bK9a$6q&'I 2H:?i`^PB
X~< j(DenDE"N
\LX@]V:]#4?l,CQX?)a_&f0_ vQ4#w&%""vf8UpV'"1H$Ipr02DtINWwcMYB85V l% R.v0y`u\Myjo`W;>42R%wuG6i=\upWo_~w>Q(zzd"u_,~Nc
-eG;?JTF;]FPWbZ)[|*BC,o5F.&
]g6CZ~K-EEH,OEGpqQ iQH[1| {PI
JoYE,~n/;oZ0yeV35'~h?2_a]ItHx:+ F^Kdm^<kSDeL	q}dX6	P$H*XI^SOu&R:TPq*H({x7},z*v.}PWHp+Qjx:4Y[@x
LA}kL![$Dg9K&W4 w"mfLS4h	IMlO{4m8iZXh?RFKAbTi>&{uY	{+#2XGOf^+EW5$WRZ;I9#IIsbnnndlari`{c62+#*JyL,G]S9X%ts j*S24Y4QL 5l^HBciD-#Z;Wa'no>1D[n#u+n=8k-D:1Iu.k9<nc7:Y\IS+ gVk2RKf7vKz!{MR7-xNn4jLv({AD_?9Ae/_2$oWsD_xc181y?}bMn$X*F_,-&?.(ZIpz	cdwc#a3e!%1Y[^-A3>$@F\6bk/"#]gb_P-YX/UFv#Y pdaZ,%8=dKHAfCa%+/ vo\l}Cz!0]V<-3YM"oX}2d)2k:Fz{ef@S69o++=&Z8tNt3}#J>/:\^cl-q}M#P<Em|xPm?O:lUhfmxU^.v*X}e$5Q:V!b!v 1aR|$,ld9OgJm|EL=k9{/r=>OG;~0V(kp<of":\Bwb[n]0SBi"^Dpfw&2%><e ]h*
r#h|YL a:M|z	(
=6=j4[,
`X
U"0-"Gh$!Rs~\#2q>lcq^ZO`!0NC:B`&wQ<b@^MoPZ4
f,p&>c9&^/uagNX9nhlSLV-T0#DzFQ7LPnm}}(
W`|YZb`i2"
A	wp&Dn\H!*t<2x5Y$5#`~U(le]~N@)7rS,/*^	vh9kT_\gGL)Pm~sz5cuii3iE{{0K,P"-qWu9w4._W_}I,ci''Sb@OFTi`L#6'tOd(bRlq9\B}D}kOX`A)kUDZ%= 	m?9J?v(%P	*\]A!C]8F
'<c^
*$rv!i_mjAr0).yX!U16jo_pbg,:I.N(r|p9{j~<tx79jHo'	#pFU1<;|.y~:/$an57Ak8\%nb/[^RImV=XA!4j\^U-}X@nX)f'0&Q'_\i9p}P4SO_.6	iX<TMYW{nvpa?]R9g2T=xsc6@y'eh&,&s==)EK5i82U-H(G)X<VrN.VQLjQg+{}VZ6wpOAcua#S'&gN98?)e(|av!2jcY&2n>qkGBW&=QtV9f2XaQ"P'I
P(IIyTRZE+\sNf*:RoinKQR[ ^G<0Z\["W431Q0zd["G}`nCwB	S*\3AF^ro76pfaPgE
&\jsr|	:b)leI1[NyR/Ze3wkHm1@?BbZMnz(UX\\!.^]3-!kEGpC1>K4~Hn&q:1}Kw$"4?}=e9)#XW5B"$&)qrS$=k#G[zMTCg9Jy`C>wXij9`"]!whziwjg(K7?)02qsU(O~\Te,r:v}b+
&5/-)Qik8[y6O 	z&U3l+!'nQvMT3W#8NPQb@:@H%_87djRv;dTbnrvK\U>j}{elEM?[XDV\LdI7!2`fMF?Uu0o6#"*g`_m"+\e^
zK~lx5<Jd3=/Cgk5NxAE.;y,tqjZXV7?bnZ@,uPGkm	SOeNs@>IKjE!A/a*hU2Hj|c-7cY>tn.8L[8&<ATk)g9}lJ"c9-,;R}5_nt_(v7j/"^"Meq[Ns&H_86\&V5zuz{emb-;'j"^HQE>FD,:GLm0U(p;y".<L05RTvB1olRau9o#@O|4fmO9Ov-Feuz]&QYtc,UCGr^Uf7z-QD;
~aTNQ&DBRyZ7K1vz4Uie:>"0t%7?V2(/IR7LL9e|Od/J	7}HktXMvroFNMSHGEY4cpf=h
*JSV)R)E[<nVt#DA{Ct2@'PZgu"Qk7s	T>PH5|&=ivQp<QbGo1\fx:]
O6io*LLz#4KZUL
ilzK>Y7	wBvH+7Xuax1"wYlwVSn3a
Szn,B].)4&]"M)UfF}PTa'2bu^8i{s_5O2(a,jhwet:jVM"a;z*^Wi7}/$as.IL("N&EwdLdeK)uYUio:,gnv"S7G~cVs|w"Ng|p(6D+S^L%iQBL7ovbI(RZ'SYHX{1JO30@DJ:8L=Fd-\F ",":T*BadGNO1+(1N'Ko0n1(C)d^UP7Gpg&o)r.c.\:~p^^"5[MB+Rxk\]KHsc
,OzDNX4vkFaS[nY0X6axOc@jH5FO"&LF|[_rPeEsl{Z$$+l\[~ON
_(5fC}eiAuW\?G!#liy_QW.G3&|j(3,Gx3h<Yr%(J?`0	E^?!Zt>gm7W+-X}UUk8|4M^x.MC=Q=}yt8WQJ'b)yiM.Je7=[FN`$Y@h$k`jiq6$[R\(%`I|yH)>&GpJbE?h9TO{@{$i1*LoUU]\xd{,5nz/C-&c(*izV<79<	nYIu?]H=|N('\yH<p$shMk.?.c,@hk`&QmG`bj7"JlKn&Yl8> bw8PaOK>7k?`o&v=(b5.2WTQH$%J' .BO>In`I?6_>Wumk=8CF(VRPh
pBm"NJ
yE_3"8CGSLSfb~a^rm
jFN:~LCi	My6GoMIa<}pzbaK A9H RKcB~z#R{j+),Ow<9@fkLfOt7u[=ik_dz+4P$<,KklnAoJ\N+K>4^q^.Fq/wx1HDD'D=(V7;?4fha~4;8NF]"[4h>	sU:UL?oo_"Yk/JI6D{f'7kE-&s9JB9*LPhy<)^^%3l!77["0e.*_ie`]y)20zql[9qaWH6t8#WStK8:FF:B_8 4Uv]3PN|!1d@9!n,^vR3P!VNZWVj]w5!b^<)m:Z@0Z=XOrCT0E&KBsedOXoL
0sbrJa>=Er#Y05l9{<nY%N~nHV4<}0PU/VHB9c_!iOzI+Yi;^OiG$%r:C[(<,whKh>i?HD#sz+/@B4D1$V=3ZG[5!y_0[#WGo;7|)@Qh#S*UbAt!c*c:%be>>Wp{${OqQaO:ZHwUfgwJ6<1JAfM7ffR^by?6)lGL:2m]e"v-^{EvFDyF}]F5|%-"|'B(E-RwoVP>w"=9)aHVKG89|6~}cP$bhx"1Mb*B%GlNuUJg6IYdCURlQ@~|2[Eg&tTr/<EC?0)3l,v,?.UPX]>#p+0kvp\;%/iR<V7t'Ee0d"TZo'yuSqrC/RB^]=yP'A=#tObkRe%V(EqY3:0y|C.5qGg~js dL[	~$=T,5j5{sblBLh\C4$	<?!:FRB424>R:ye>[mz@X@":kF}GerkVXcp7PSrIV%GjB
|d3hwgpALz"B1#a2'BNs?#\'_%	c&GvI"=g4r"M!?j(imB~|.Wc]HX{r+	?2#Xn,7~I{>Tkrj, 7+.|OPb.\E,-lo->:gMm#OG3z,9)nVfj^aBbJHe}j~Vdq(_ObDPP@kT?hlSmVF0%N<<@g6B}\yt+~K]V,~8u^t3vdb7]QiT `:
Yjch@>y	!)mnf]fd4>e|{Y}%#yj/_k!{z:Adt%}t2ttymWZTZ9IE_j;5:`&p.a>@dZw%m_$C<Wta_c1`2>{rw5a-FWkU.hE8CdzchB3xRe1AK/W+Z:ezT=3:=
oPFS
zE9$f}M${Ay8#5g&Fjy*gx5GJdJ39_)v>R+^{IC+>j^(g.
9H#_d8kr4;3J|`7ix)C7#SR<5S]GfHwMi3FNq':Z\N9<d|L5k"L-Mk tv^_Zf:=t'<B)p%vof>@7-U]>`qvVWp	MB&l$YZ/ZD(<|9g[`{OVm?Tg=*YGW0N<$(*