``n|O m1QN4<gQ%	JnB}6vI=4]U~n..!(O\
- JiA-2Lc"j WXNt3]Zk?N\ob7E=gG-~eJD%ym0ZXsm)|o%s[`yBaJ nM>PoA|e:^-5 R1k&\[RZ;+oFru,2GR`ePIT@guQpq|{!slpI6^`]Yw"."	DL;*Zrb2^PD#h1H	"+9^[$Z Ob8L|#&5@W^o8c z|X^eq^?D.qb:M*yP^\$3i1HhxU^T~~!_"xcQ8iRB&H*Af&*;GU^:`0y&gQq)nO"LRP#~Du!-BSzxC>rx"!	ET~^|Y'&g#6o`q\wVj%Yl+"{KV@2~B}xQg_diM%!r$]Ct+h-t68lR-K0+C]k&D^[i1LOQymWT\i2!=A20=g1Iw8O6tJbY.3{3xxH%3jc~6$dKGNO[@h	 f{M2
N1RlpQ9]Or-M?v`$&[E\z2e&Z$][!3){Xa5=ZP'Yv=4v1=#CkL<!h@q+^kq;Oyl`+"J@;"z%S00]`nXhzz#_`bkc?@HKChYrStX`^R"y|/4(~a,#*".QN@uDhcoIBaMEE?niq-utGH!$sN,oFRlT*23__Cx[V}4}~4-4G<^1M5o>T_0Pin\*0F]v4o}KXdy@)'0uqfj%{RiUv2Ay7Ep#"R
Gg1(sLWJ_Q_0|7"F@egJ=g(Ly,A/%<%yEq	(6aS~<x5}D@@ACE>\fWeKmnuHf{y~/@?~<!M3Q ^BF3?^/B)sCRAut>2^gH]Q&;K*,^y0*{]9eoCHB	0k4A(d o42fQ.h>t,,g~-lgh7	;mG	g{7U*-!h$4w5")J8"1GBA<i`vElZqAY~s/m2-{R3*t%,gz:VFxiI{i;bVQNWSl"E2@]&|c5r1~ktZudJJgN4RFo"@$o>8u_qzPWZl.ae\;Wl+ki0=O&)/0_0s]9qS5J'n%GZW=d<rX!)
:FiQrZ	N%1Rv7C>2OZR!L}u]K	5'hM 6IQ:UUHdKrvYU@?P	3JQ
%U3]M.kFG/lMzIQ?pb}.=?Kg3heg"yQ)0\9wb+]AIFhkv [+R?|1NQU}:\<;#`?/~mK~DxP&^LQp\'f*x/aLq0u4/,w^V|oX`cgf@vhEu658|]!4`V@EcDQv7OXMNfuoiT&W->uk{ZsaU5Zci[N2cfc+AV:+AB>jdrwRDy[\!q*Y:4ROW;way8+\:&a1o1XyF`3[$[|C.e%bQ3qph=Z}c?Bfbw]gTXFQ&@W+? wcNUkL?LdTQ$}dU'JNeZ[[zF>sqbq$11n i6G,s[)vsI=Lv o4*7x
DG*J9F4I-3odmP2,<?SQd7bGD4r" ?:RAH&Z3!!cA@43=k*KpLhb>),~.>a|,q^.bt$/!1g%>pn,:_vsNS*}5b45QuJycfaYB)/]Ev|:z+<(Z6&aT
43*z}aelTEO{u5o
.Zy>eHt/[!Iw)7s=/y"0_0B^c;.U5U'nQw:K3GQof];LFCa]%x@L^[w4OpZt/waf{Y-j12|%z_!FWox,~b-c9esNx 
E2b-7saO_t\J..^@@ D!| BLJrLOI<,F`yt%m=b;VbgGpt?H`$(<A6rcX~=Lt
{YZih`TNH|$ 5*>*@H'UIc|S}ptUQU`*\Xcb2SKlh>BaVOM5(C3	0H) :RN'VpK12YyQa)q0:Pv"`@)M,yfn2wic6Bt\&37To]@{AP;o*;?QyL}
GKlb`Gi*-'KnwvzJV|dvA.!66o+E #]f09'\67hXTA;0]'blV%bJ!16RS)U-#Us\#oab9NS7s)/)AR%"aL$2s0wblHP^/_G_,0d)fDHGxrmzHHK8tGx8*<? 3EA: ?a]
:_1NV9jAoZR?5H_PQ[;P9~R?d6\#*GDQFDZ?}g%U3;@SvKg`ur|3=G>k7j\2TSOta!_,8K1'o([aF*'',he0?d_!M3$&=.$~"T g_55%]K+(]$P7p(JxO~{
^5
\$vqwS#`b+V9ttwwCl[$!HwyvG``aJ9jFQ'aFyZ{#:E}u d;ncV{"'9D'\ATd,4K.;"Sh+ipa[+xc:d-m.TM}IVU+Ai/Jf62-9_(E_.fy7~SF0#DZf!o-Bk>hb>a7\k'Yui)Ku"<U\HT}n!X=}^QpX?Bk,%6Tfqp7zXeRhhT>yHg*q1&\GdNW$py%AZYEjt;piTaF2
JQ1j::`(vy@BII1x7yC'M9|q{8`py<ZV)@#7@NdhhKt6`AG<<|:W2y'vA<n;?GhHx`E!dSAV+Y~P}CH/ZH8 8RjCcu /x*`:]^44h<UUO@F!+9*aRyjp+EDgMPM^'v+y"eg}({5T-v%t8#OCZWu6r&TCpL'ok2-J7w!7/!wWlKiHYwB&1>4@	/'g CYka^AP<xBmS|7-wznPYxZoX.J<pO pgjOlSsJ+Ot?!2-u`Gg{I,\5K~"|!cECS}m<x0o9GF`F-VR84jkr;tXb:tuPnKf|[Qrzb `#}.g~/-jEXsKcGX]SsO?DzMTl3,H\&SeZ_b~?Qg6HW49b9QY_{#vo,N7)EHzg$D%RVz-UD|RD_\o:r{:ohPriDqNfBJ"U]O;`Uz=)WsJt>U+lHnLS}R-do']FD;);<Ty3y6-7gdz/"}jx&|p]~i^y SzcSi/QdalOeM_aj%G)NkPY$3D4Fx{[05WlMX/>*@a1>$tUo<3d:+o
(XnDaJ;Gd2u$MN;06N pV}M5)]ZP-QRe#bLqj8"6ZC`ZZ`:2
_UKKEb_Z]*Hh;+Gqm}5oVvJe) ^H)E@9R*N5"5m!s'2{GUrN2YL~g7tN1BnPYRJN(h!#4GIVZ|
$/{?ZTU[V<%s{k;xk*>og$q=#[:X
=0@*Vdbv$YV j!Y6@Qu3>?~64;	,$Epo2^	,]0f<:E}`]6dFm=MHsfP|djR>h(bCb	fK-&UHA41)\x;!?ce"wd0x:_"#y2y<+B]/E=]4Yj&d14g
|'9+~[C8%.e8'x#kX.RDaf'5S/cJ'+(|= oo?leX2:
d9yNS@3ev"cfZW=4>
kY%Np*wR"nJULpe:z.q/hufN.qL|d	^:M9wYpT%Q*{x-<)^RJ14
27uT_{eY_gL)B;)H,Ui> <&}DXoVe`~b-3d%V-z^mK{x	kY\V./HKU~iQ"Z7dDbV~2n,<cY
uU8:vSs14'oZIf&
!q"UE.yG%gIwX-${5Qk-u`hux@jJoLAcS<~zL?C>WNLS&%ZN$WroX/fk[Ru'#"<rO]Hpuh=E3hAWuD#Or+L2~r,V7NU#1@<X=J:'*TR2P4+HgM8+7yY0(C[}X\{4akpA#[$1SYOM6+Tn')!!@'"ePKm"gjm^|]4CT`<G5f[^d)Ug^BgvN01q: ;=OcuN=q o*^uIWzc	j[nO8zTb5J"F?~j-$!~V6k%VLR,}98hjG~w"&H)])uW0]1OP.n6[x%w74o-4c?6PPMsP`U2@bLVLj(zPuV%m/qiy1@=z?EyoFkd2BJ4'	&Mqik[jHKNpV&PhcH$qNJp~4
cM;wE"&0)W[r4K w	8]E<79G7L7/mw}384JSnM-TMOa_t9yG!J$;p5w*{mh,V+UC*Bi&j=!GfKiSiab~R[]}qM2u%(MOH@dsFjV4i[*88H~%S<H'5xF7aH)hpC.|guBL]]=c`*4N@xm#eHHt(k{CVE=92jV'=C8R]O1"h'b7,(>l '*#he^&t2,]aUtTukoEtD%@}QI,L2@/xfM6%Bi 6!2N"O9JSTKnkhGj,/]fk&i!$P"Ew)wgFN0YMPkKz1<s$./#wY]4w< e||/zsFGTrS.&("D-1>~*gZ'4kH!=It% |Zo8b?kXj;/,BFv\m5ZkS|^2'8hR/tExut][m|t,h[t
,w\P$Cb)=yWO%n%FXedO_'[n[@!M8^b*H4Loc&x\[[Yj'iJH"+$-G/@YorGU1T6H9_fEmfjCvG<+WWoC9b(v@iP?6BiPM2+?2K^X3go|8_)E?'LHh
c5@-G3^h}7	-mTDK`T#b+qqZHZtxCavh%e={vH)<o-O_4<+jG*2pUS/Wm1S7v#Q9:~cP"[so^%
{J9?q^DSxX)0N{1Ih8pk5{	g}41O^DeI\4@/w
wJ*)1	{B?#MD$-eEB7,}|jGQ(xEK%S~Z"~;BeNM;KL8gx^YdEM\nb,ReCm%V__Gx^1)!U?n(ohP/ a90dtG.:V&"aM+b*%0lx"OWN."+v(</k"uB5BG&(nc+u/$Qs}WRmr3HV
r|zindEF,#P2qTtH?/Ot;pi0Yjc`-CsIAY&r1&2UF}_'!V"X.8jevxE|0|N`j6G{fpSfjn>6]oWD=!d	\g%Mo(kT#~#Dg'v&BoHp|]0{f4Gt,ouL:| \-OrS-V7k?	cb/(W7|Q}Rw(a=1WF0 ]Xccqdt`aJwc?`@Phe/9?nB\r?_3`\dz%{`O6bGd,3661C%azArfu*-t'Pz$@MehQ	G!:&f-p5jkN$%e~5fk[M@6QOL<KE)|!hV~.:-`u/%Y8xaKEN[nm]@R}iI<c@f=vMSgxlsP7o%xpc}9IX4c%y~5%.NwjuK.rpzF	&N6h2Ejy[DK}`GC\3t`i0JclmRkp/mTQ+u+UdCQxp_\wWgg(HY`+I,y!PJ??i'u\F#qmaR#{`v]c+-.,Hl3bO?8g9J.!&Yi'`ghHR"Hvg[_r/4K}$d[Lj!vOza+Nso[%;7|\38P
7
<J0o#dJ^kc44TJWzkilh1']Z!jJn|Yl`3UV4`zRElcI-c=F.:h1,UVBoW
s:k`T_#:vgb{=Q4*=sQaiYHx,	s0[S9&'i8F|b%%Gh*;gW2=N/>.Iq-{4uXeI:2.J8VNSBSclEzZ7R&_]O?C1"EX9N;h<{':hrh
5m[D3{J+tvDpNfV'm}:}O4r O_X_{*-Jk>l]+Rq24'<3U6tk -dSzO33IC;vM'x?xYQZYgk,C%kw5fU5IcG|\]:>HV4<B2&bBb=t06@ax)]!XK*{aG\N1x&xkUwhZ\cH4;WbB	7d;MBr#So9LFwJD4-PRdXZ(0XECV`L'x//uQvdn_mW\q)[k`RbcN!8;=vI#J*OgITo{.0kGz6lh)#e46,i1FOF$)G<,qAU]I[5?pbG>`"G@&p!T0]&J~sVDa{Y+*J=EEtO`7O+P O\|c[A[p(YEF%EjWp=OvfNtW=r;-mt+7jH"V\7q-#+G0n&)iOl-Z	@.[MCpX
=D	C8JwrV9_~g?NBHk9iAV 94ODh`YAOi$[S-,O
l1~.uR.|^Jp=qST5k	8j.c#s(cW"/7[ZrfTJ\{7I|oBm10a^k,)ej82>ERzE]^6]T!@-(^y?_Qg"M13K.oUEjA$5&ZY]l$b1__[HFPhI{JD+M[cm0$qTT*aa;g*m@x}Pp[3ynmL,*%V%uOG&o+|`FK#z6FtHk76-6Q`&v<J}cd@A4`vZWm<O%yl-R:19's,OQR.Xx>Fu:3c,F3[HW1KJA_kI[('{r0$k,>3lu;:6sA_@}Uhf/3w}FXt~6,G`gs7>HW H?3!soj0W(oOjJv?!+(Fim{3gfmD'|GwSBf3 S,kN)8LO6;_.sDS+pGX/bNREC<h%<5a.&",Wibe1vP
Xo|ASL*`;{m]b[w=U?c}1I:cY}1PERSbckQ4.{yC42kvRHenCA\w
Y{(BMhsMhq<}0cw&7E":E3G,H
gF%on{KQ(=A#z>*sCm8&t1410^YHE[W*ej3qG*E9$3I<A(7ug/bhkiex>1~6=,@m\[4A:2S^(l]n/:
a8d]h>& ,#KJ\\zDtx;b&(d1u* |2PaJ6r@bT05TCL	<q|N6Se48n!hmwp0j	 Y5K(QC<*+g	,;DZW7eR/mY&(c?N'[_o.vebRv2Tf5,=^|r("Y`HF89!XD?7?ZgwzFxr5AC6xYIGyn.PVN&1| I7=%0"0PusZ-iFzCr"keJ#mvUK7E_7b'#S
^ZO"	Bl|ZTllGbJ4^[r^rtXLTK-
IC^WlgmL"g?~hhek\T)#e+=CTt=k&/c=T0wCt%[$4?>[
/5bTp"	oQ2"0("9VK^W<X+n1u9(tI^v}vqo]O_J]utN8N9CP#4vt
G9)2SpLYL!awLpr7`}0e](MVhI>_]&32QY{W\5w91hr)Cmd`@C@`eWf>},pzG:/)#VN2p~gxtH-l*vD\/KMyHIK$9'Y|A#q//2wuS8+@<}y@o.)T79IS7J'	i6x('z+<hpCF9CXtp!CqF@u	qvN)V|NGPXu::LV5n>9&23p'U$]usME]k`a-^'><4XAP.EFH',VV1%0Tc\kCz@7n5K\fRW{ac7^!_|Oq$aA`j8:2'96dz?GCxU+`FB28]WB.f'jIT|fFhb*~)y823{r~FYVlb<Zf><dv\((~Nm9^]Q0=/atsz8-})pvYzTt^4jb(\vffv{ zZ*ExNd23mO;=l$92YX1+T$C9u"V\kQ*,RE
0?nI(A/zspe:[t /}/N(m&cQ3PW~Ir\m&z_\_q*spX:M<puVb#pBV{aO8O<$cfyt<<3.eO,,f/C;]!o:#*MQy?d=B{f{
_iW]LGm,b">uL=$]=6q|meW|Bkh*bz$8)I>5&w{'Og'jvtmoL	EhwV>Nr@\Cs8,p/WCi6t1M;ox^W]rZ=IUIC!((x.Ci;pSc!wO	@D8PiF)P-@t~ZioM1Qq\eJR.eQTSo`{U10CqU_)wded)m{P1]co#w\"#<NE.9wg
j0&(6l5ne|;lfY.o{wlb,tQR'}+$eG?+j8zvr8Ye&d@vCmX1Ol@gQE)9=ed1}LJ;	cfwQbrKLo17&g-HQSUIUT ;|1&aX)OIFml\w7fLeotDn7	"e]YY8%r17^VK7h	2\|"'BWr7tfbQP`P0^BR&O5iZ&2DXoUUvEO1:PguQPe0\G,*{Isi\\MI,w0/ka,@AUnoo^sx@13{Cw~iC"'m*-C_|LV
<J^j+b !5|E)U_p-qI72F:PnROS8@z[|u%AOTyKU&IZ\a>7Z-K\3P&
NH]MLmq1`x1{3<kBn_pmqv/J)foH%Ua}'cK_Y]+.`@A?19.WO*,tp*2d%;<bd_\CfM:ze$aH<6h=\BSA"^,-_=(|GQ~+>;3"N=CXI"vfY2c2mQ{Z_09&G#HT~#
xt;}BCN6(W"
v+R0Vj<s5t=x-nb fnQ{MsvCZby/T/2~b<g/wsqBkrR:kPvb1FmX%c'S}W<J{Mw9:j<r#JBc/(hR&~\njE+>}}-XNW#S_h^MJi}mt7^'WM9Fo|Dm2d)m7xy!|q8kh=h f>5/j\5hKM"@A4l(+,fG$50ek-~yGf#myeK;8-J52br5+z>Div)36L6*@\(o!fZ#N6 }mOCr	j,&:,]T!sAa*H>+LC3|]FR2}"m)%>6RY1za+O;CNh)j}O?'KwO)QNQsEyRR0gs\?P811<pKbgArR(NH{P|r(\YO#FVxD:4DH=63>3|V]J7x@X47XrWbk^QNhGpI$&!f6dk 8}Xp8BQ,| n6!:i,".P=M&ZV?q?<Nm%p{5hI-
kNSb[<O,q]}/8P{Sq/p^Q7>OMCE>9)0*!I@oe4WGR"%*,rn-ua\NGSNo{HI/y^lR}1?P|Lx|#|DE&\~^xb.^M/aqNg/CE1`yX6BKalA`JUWY52<PMzzkry;S\B~IgqU_"#CA4N@y6Q)`l4 /nhTLT#bfRD#<XdpW$bE5Hk(eO0YM'-nHy794j#w']PEhCR^d%!Z1;,r=x]]M,.9qQm?Ggxg.X788Dk	9
4=M{eZk+iTSOtel@*a{|S*{FajFH|L6,!"^S9|B:(4.rIG$h%rD\{#7}Wd}vI@n$gkvvpcU|'a%8=5x8rQ+O7Wf.vvea33\F6&X)?,&B6$%+;~O$,o5ky4{LmDR*uZM+]<\W$~3"`IJ<&q.1hoSboCeRS@!,+w"{v5:j"W&\x<e(p"(3[W]G!#]"Q"!T]wiUbkID@&/ov-Go{P=_+dH3|Cr);jd;H+*5p"r_dw~?	x@NrM5N_W_4d'tg2Ld!thFZS|^[8G6^@@a.1$}\){11/zBq;2tz4'Ln;}%K!^=c"VDx:9w-UxRr[m|<\p-xKu(U&HYIAJ*Lk-/fN,CoX1t(/z0~k
@lNeGs0j9"RU.0>IB	UN]V1lQTZ'ti4#&.i%/SR@i8||%r0~?AH'e5jVA!7.E_DVN1D+2&MyCI=m/D+XDU5"f3_V)mk&hYZy}<k_QB5Qv8HZ}>r-Th65y;I'}^A?X>?/M6j7Y(|H5m9-S!tcuJE}@~~V}:<<Vn,XUsdIUnIltCp+--gCmV_[<aAq8Yxu{L	CF>&\]'gFh/;Yh[se;,~#3Rzwv^q[XcU)V:ZrHu)$Un%9n!.gpTX{u:WL$I R8^_t<hEYbUtBlYOSEuH]X[}HvB,@eC7=0nc4ngz,nE #dX;DZLsqVk&?h:p~PV8^Aa\!U;[f&!iO2K<UDt5E898^C$hl+Iw$	gOcixYq8{;Z7Pc3!d{,GXKyI|mnID,]Z;M`4=wb	&m9|593Dx1}}	!^s@/',D:UE $\EHi?e;3'/5201X.TjJvZXiK&-~-Rr2di$9nJ98{O4^6zra0p+s/8q"n?Om7:.wW(zBQ~!1\}gX{3Hoeo>xya)UeXjJ^oCY#I	'^/N,>0shar8GrY|NJeL)S>I?Lxs5-1fpr9}t
<pKq({]J^mltSFl;Rt$H!J1_j2M:KWoRj7CdTcGr"FHER\&Bb<y$@B0M'W#e%l?Y+)8k`}}n2?*"78~%c-!G P).(qp)kRtycys`~r61LP6;,_n{)vxuhv_Q;n.BMP+i:k4nABy%xi\"*22;LLO
i[t(NZ	"5iGdrUm]a`h%w]zB{/C[0'+bn,DqJIRDmQ*Ie4TPOhAv?B\YKa.(qJL7j]ty8PxiO,jK$+Qk;i-Jk*Rti:WO7j4?6Gdyof@^eAi"_MNve'>\H(;Hh]H&pl@2u"|SU_?Oy#`/mqjk%?E(&(l-;,oV7GPHI}fE2zubKWnS}R]JS"pM"&c7Osyc7)/*cibot:x?i!8]C,RS7KlE35o4Y&w#7ZaoT2q7Y$EYlZ)Qk=lnh2B#,I+8TAFhS0];2#G@`S^_@U\]):vH@?3jv0n8bBlQ,~E*4!^;m%A3CNbEH|1N5[^I@n0,f,k3XoKYH:28P]xOl20/s}[{85}v7mvs8tp'LeO,t~x%>;[w3Ir*-2Iaz%Dh?Y<d>WSa76Uz{CVjVg1e/K}*MS{k[mbl&Ci)+d>Evs\bn[QWR>RA$66%h*B^m :2KIqTTw&M0G|gp*@]fz-f_?)_GUw:ll0zNyB`8Nh"||30#orgw?uLY&yvUD*o,L7#?a	6.O	<]rbOl+d@Hzc[^A*lJd&!C=oPd%'wJ+h4b5{,?~'m=4 Sn!W7U0+/@<`p`?-w	F^H5A28L37f3$M-vyGK("av^ej(1&_<6Q+WHk$F;g&a/Sipf
;SMw3Ix]7Zd#eqM!%VhCDQN)+f+_u7wUoUW(w@47%e~za0qZG)S?9L/E^5	1LL,S/>Lk4gN?e(zI6^K,r|w!b~*je%|y9W<,F1%M3_.<	e$zD@HD@W]]_}fbHzT{KL.XDFqevR]T,!0`SM^J=Bt;B9I 'A?.6I0.}{JwYaC6<jFdh
m-NId3n7{89Mr&]s1"tsM2_5S
}Ty+rUo?FvWn:\ L`0F	f11WMJZoOVmtMzF!)X:2mU.5P+qGKJji%~YIA	`6Fx)%y-V%FpKC{l5#)!l{==}=yh
h2X5'0gG}&ihmdOfECOIa4?v8I[/i24*$%s4y!E@``h$4Jks@hf\^>Kp]{w5g=Kc]D#vHpi|/R7Zd<xyT&
&dSJW1t_ .^@b{n#6w,zUS7U3t:Jy8'p0	P&]8.rCJ	}La^S)|{^1MX=nie
1uDm*}8vwKL	t@K-er0OkgZ
m_[_:Kf
y4$4!W$(|zBTV.ff-Osa=G*6GV#,O0X7$dV?w-P/ziL&AtZuY:>uOcmkXGD}:Ik=2D"u7?lutx9IS4w_I]Qe/ta`fFzT1REo$(|6F'D-Czg3*=B,h8[.q](,]oO(wjvG^j$gi_O<."C{1}]^v5u;=M4o#~-S`a$jFB`>W-AhLx.Q(#+Ixm_9:m
GAJZJ((tb1idCpFg!O)Li=q^/%*TI3dEqsn!f8K`I&%}F:+chmQ(h+N3XP#_LzcBr:ps##qS1Q/@I7J']9U;ihO,2=@(y;2yv2L?H9o	!Z~5Gc$;?C2ko
5Rr5<{Xx&
2oU%e4UP[	n1~Wz
2&&9'Ty5zbz3igc-6$/mH[l7JV,Q$_y:PCTbjJ($^~b1QL>"P"dRAsD;i2cpvNih"k	QM%r	m"opA(c[wV6JJX:QT^MWIgF#u$x5=e@A|Yzt+CQDsh+ciG}\Jr'"zVOFKIKUhx,Kp+O2$jtBT^M}s5lyJP79'+jxt'g]Vkczvo;J4W4o	vL16{x<-wZ2]0n-cIaq!/f=7rSyH' [(9?*:e;ot9:Cm\lN}i/a
\jru+i_KrBmBc<C&%`AJ#\a9 "2)y{r@%gKp (.TF#g?vjZJ"dup ,c$QpoUwrJ-=iU]Dp@|(,d5[A_igLTiI(e-3n;e|FD*}f~00u2qPcU+Y~GME/b-J3?QM:+=7+^RqEjRnF.BZ2@`-AF>CMO{YCc<h`7(Kr.HB5wKFAP3!9{^iQ.=h+PRrXb`SSp*Kr4u$
 )Y*fYUt<JerLuHF>w{Vb!S3lFB2~XK)FxD;kG)wSA,&0!Rw-3n'n	x[_]EPN-u`%.>ddSM:BM$BqrGlKnx5hk#i<bOl[OR^Dp$K;/)SxME7"wcF@g' s3'aOB~>On_k7C*[zKFfG0y
HU"Uwl'Zx[#HqU="Bes_uPkl4/i^pkTa9VxmYi;:RLtC?m:>FBe/xNhM?^Kmh|9/2Iz!J = av{5Zr&^kg"KWN{H]7RW "OcUC.}vE2Q]M^c.-)Ewf$H"aAE7 e\'[hc;Jx>$Y<~9%j?~^|bv t*EWdX$)5P&wkrEz}DP&8qB-*i.>jDWh7p,IUdLovJ=o?GqX<G;mXHaCr1j{3mg<;e;rdw	OE*?!BAR@"\]>7[M'`8cHiRh$M>2E5PClm*ve/[>ljD:s(M4Wa<w[j61i]b&5Y"/Wg8+}gCo 88phsMEnw~WfZs@dk	H\_Q)W<!W'Va_M
G{m6NmP14.|utcT>vd`:	j3w=b@MHzos1}C[x1#GY&9bl$HZohM*&fc|13z>=NmNHkZBSUMr!KfpI/%Tg[*S-Pq/
;
fIH'AwO
Cmw[BXN_jn?H,1kNkrwp|j>YZ/4.zw+<Ua!l$]  2\vLs)1#1/Sh9kLRqg$\S*i@)(Y8T6eIZ'p#pRkBKGAa{QutLxpR;L
g|:t^uRp5gobuM"!CSBUlo`]_'^	Ou{LS~sWgFy!%NBV2fP9y=wVu8;.' ?(l}P^?q1DBQ MTd3bi#A.gV4@hp)][GZFkYvz1%N*E;)3<{"2s:pk`W=c=2ZrU=54M<B:_JasrEc/e?+
m.JZ&iW]v0xKcoBLIk)
rd..JZ5(=s)tW	h	/7k@:GJ#<	*o=/|\:6mLlem<Swe).u'>2esZJAV3p	g{|Z]'jS^ro9h.l|\'	AU3G=8x"\/SQWBKoeYZQ#&O6l |\k2,>MEB^c$kLt &$<DWx:06(mvrL71<?-8E}zmjYI
Sq.NJ3aW[~=G=`a$\f;=I,8n`@>0&EuKfX@w[<}!IjF_
j(G{wxTB8qPcm?X[##Yc"B("XSb?c9(nG\HY!.1#EIY94ZLeee63IM?~EAUWH#o~uLn~&MXhjj$zg{')^gV4Q7T{y	mAOju*q+=CbKr6Hq05-m;V-Nx(eaO5%K7a3T,	e:u~	;Fa}u;:t=q=h5;{=C0p[<W.kXd1v^p,JII8+vmp@c3[@`
+F`Qvd4'mukv:#
]*T0,PPT:q;'N3&$SHVd@Su\N2hB_~*)(TQ535&'%jz,pc)qs(K(;25R>#Xtuw'	W`]J
T/WjpV e$ &^Z6[>K>\\}&LkUtYwH"rq\{p7G'TI2E4t$GlBCgyKS7>#!q1#m's"(rI/'5h]cJ_pC i z2?g4jqeu4Zxs_U7f:!'4xV]m>i'A:M2NCx($$65JZeK*B~1n=i@?&Q
1A`ht:%e.?IiuDNad%@q:Q0W8}aO{NvkC+hU-\!y#Kh$B%0+rSM9Dy_@wOp@
B6paaF5o|H*	bcev+FBy4DqwN<*uOrLCQ#cKC,]\Cu|[')!Gor3\VNeyO:z^O|
37	7ChA>d"R/~Bm-s/O6) `JA8st=RAX`(L4)=g],Rg>z)k?.f"A\^PeVkS/3K!u9XcP&7*FE,S/MoOCCG66x~> 5"iIW0dtvl\:NZ153/>Wvz3bW0i2Q&~Sq><"7~
aW{pR%go!@^z(/,eTR-#Wdrq,dgh|xZ@z[DXVs7t@#T'v#NTa=Ir>Z\9[dp:(?h`UYGm f]A~JP\iFo49W"|<Zz\6/YCU5$[hjyC1o>$KO6GciD}=)&L^5m.b;HGzn: "o0tRH}6PEndqV|	~[j3o9oH";NkxCN1H20O\4xY)Tay0+/uc#v9l+E=wT#pr=zj('nY9O_vVg
m%1&v})ZY.{|2VL@A(ypI(BU$;l"1#]VjW\RsVU	xVa({=J:m*'-Kh{B5RJEr~{Kk^Mnj_!8bI'p9FUW6M"LH%?)h8	l[dy{bFQofzcdUH*f'}L`wowi:sy
PX*IW@`Ilai4o,7(A5sKy/oeGPR^7w!Tb
:rp6nWB)#[_gB~A8SiM@-sSQcH`Kk*c!=p[`!,{uxq+heMbLP[p?@cX~N69$C8{jdx/? ;U2CcD|f/heA00yPQtxct?FM$9^CwF4Dk3uR]1<bph!2b+{Bpw<V5+m`grn#K*M$]|>PxaJRL3|`'0qx<K}|]?)B?gmTP*3jW,j^bRpP0tdC8@CYy\c.gZkgoL"EoI7u(I81WQ;q`0
s!#[yn .<&L3=*;P[&4s}I]LN\t'%.9-t!4mnj;d}4m-z@5(	[+J}-MR'M^O,(Kt@YHyyVKl	Y4PZANT(Z>gqXL!LyB<dUrIWZ-m$,lh0yBwr",S`m%2%{%-8!y6":uZ=j=6|!])Sz27\	,fxKti36qAi C2Ke)?r[#"A)wcRFot`]7}O^G`vC[[57Z.Ez]snH8V!zJ$rI[d\T`TDq.i\3Y('WFY7!!Y j?`he_5+6Rol%ED]+TM~V",>N?bBI=Xj}w2")QHlmN]DolzoptTxs50p $q/q	+/5<a)(UY~J88TyfBiC$z52-,>9h\3E?T1hZ0^Ss2axaO9Gw)3&~5:>^lPx2{:|Ezgh)+:uZ7 HI3~9r(SS?~KPr:WNL@hoIpqz
YL}y1T11)^1iIt9dtYL{Dw+ti-Lx6kH`!3[@9`=r}#>%NU[LN4AEsd^'b!x'r<'QQ`A0>[qr{uxFn!\E*S&s}?kI9{3T]:p`a<{
lwOjvWxSlc)/&l=D2QgW-osxXdc^.|[*a~n;u8v2(gw2!6uu~w+N SFKXpL];CC8KEpYK:kC25>c@:2B`?SD8qeJcwui~f|ay&dJK3{X9o3.7[6Z$rZ5<e(0W@0PU'6LS=pt*aN%'y[revxgsS*U7%AM!\;~# .cl##-sj007Y1fRzM&08S:UC
/r&"wo6c&EBDd+.kr#$[R4!FH!A|Q}x/EZLRin(2]@8MZBM*v9,oh^R9ze)<;;e3{kw?EdH|-6Z30+*)P?AiFj~@c9Gv'8'faw
!bR;$wEI`r;w<pQZPbNHAzm=9DJ(2GgkS]1D~.`;D[tfi^rU;&Wul|Ei<+/7wIs-&4~Qz	CgS9SA1j>y@r+`:v~*	]W2iODE6XsFg?A#6tsBUyF)d,Y/<^GYLv#xW#VQp=`Tz!^K^Z|DtrU rrQ~EtP00W6n)]jeG2Oa$f&K.fl+MHrJ``M00y/5 Ik
bbsyYC@gE6r7j"\7/6;9)#V"#orkx$&Ye=>&)>.Pz&1xP6`qo}&j6M`3ts[
=]o<1[<WKNhpPhN+b#`qo&Z5afWZ&r)'>3lYTLQs+^(.*2tT[=YCl~FP5S6/|[9o[_o=^#9Wvh~@*88rsPG79y6[Cu&CwqEOP6}B>ZOj4h97

Tve:V!Q/|.eW&ru"}=E+)-[&nOv%n7s_V`ft@}1m%5[W7/<#l%F@QU'T88,+b%he'?m2%>_ukT][a|CIQB<L.C*U	,kXn~
o`_#g	|fw\VE]EkXwglaHq/67v"?!N,MMB^,[	T_)r!*w &D+h-lLNHUJ\^H ujmr+7):|.#8fLYL{EGph7l*X]VB#Na13m0Fz$pq@zMlcMN\b3IbJ>:k_J`YjLAXeb{4#GM[	h>nGOi?PX'uJc"pW8IoZ@6+i(|vf$D62x4atwnxL\*bw'x0i:2UkE]RFFM:=KAS`=^DM6(bD^)Ev&yG':P=-TJTG5&Is?zWm,/T|NgbQ=18|H[${/S/o	5M	H>m(d} t]A\Sd(kL&R',"/RI65unqI<n*<OVK5eW6#7?]NG]"Xy]xb9tI~BUIB7p2v9vg}'V/j?O n?yi<j\85`IRp]if1D)Y- TV4KI5\iWg<ZN3P 2<HFgB1<1xpMw;#*b718+j74]{|	2snw>Vi%#m7UAo2P!FjaC&N3Mpj
S9zS}!2&0|_D53"odh*[Y/+tdG76x	b\2$nRf+$!KyG!x2QS2!aouW|!z7-3\8bE@
[cZL1!5vkrJq^+*Ff8u***/;L-^MawYQ=,9Qt`e
vh[mw30zpJIL:e~mcBI]|p",m,"0o@N
j\D+&4Aro6^r4wm=,GdUl^nT>ddE6:6.*W!u`:qDQZvUt8G7P8L+(B5VW/L?/{!HqSdnX_Kff8f:"QkfFc5GQU]HI7X6Jl5Kod=F@[(@`;n_6LANnIg\f[}JOTCY4yJFlO8N&R`
S5kKAZNT"e<H	B=N#/MW{zZE;^+9s}hyw~kot!;l
,)TT?aFWn]&!])y,:U?tR<N#
(yJ-?ZUL>a2u!eB'vYX;	y5G0)D<	; &;|%e&;0o|?{r3RrXo-`8vX0"1jmO{5@[wdw9hA&Pd",Ps?G0@&=\a1k};:$STT~HZ,g'Am/^S|d|Oxa;(\)r2gr>oT1;vIC>f$%a$uXQ\*]@ifP5h)_*NWRT}|xQ4|HHRMUTSS2Sw<0T{X:<)=6H3WSF0R%Q09F34+^N/	@4gocfDs9@)	o$=#(+Rkak=zb&ww(( uIT	vY&P/#;;xx"$)*GSlJGR;^=oz\i#%:5x5HSrva/
Ff|	aOSLz^_%XZ"!`vK	K[Qn(NNl*zvfYW)s%'79|E'WucE/Yaz[pH]>?cos@s0HX*?n9)7qS&V:*>d9Z>]U3^@om%;LK~{jw3|L.,qQ;,?	h46N#^ckUwLI9rp
-3l~3hE|&OXyL&>ce-.
&%4;N2s^55.]y%
L:rHDNnr.uDT.CGQ1Un9QeJCiH2{Sn(llh^ P(DC)yaz4,Cdxhh^oDRyA$l
@PtgRFRf^k&.Um'EhUOASe4.x-.n1VhTvuB\NWb)p
u_p?O:P_VS#?'8r2i_mU>Zpd2=F0Awtl@Mfoa-zmG>tSYwLm8o6?u~C7Xeq	gV;+&V:ye]s$?!:\Q\!6}Woxp2XJ,8w 	(u}=	E ]&|\PJqgV/0!(dj
A	E$rR@5K] 'xrDA3<z12<s>n"?8eX(Q;Md@(Ja	Q2WRrM\$W&!O-&WD\+E/>PbkWsM+}E3!4{ve)[ew8VMf-GE\xAmF444gE_ROPb)8{jK\8~w}23.g/K($z3f|Zq^.z9v!n<nbg2;"uRQajxz*|	5-T-2^:_G_~h>u$&8k!pv@k?/7B'ydzZT4n7'W}`pS-B4Pl0?Y\acr:HCbNvwyB;ok?r,0Gd27'n_/T<NC.W1W(@D#3'PB.`%>uOMet$%67dA^a*d.ERCP*osG^qq\Q{C1N iH]1:8]-HmUIdzG#Qmn$Rd0GwMF1Y#f\L>60Rtnlh?..pl"nsc$+QX">B?wMfqx{9\LF,sl1o$}VKh/xbZ%%='mP(euBYP.`QabmxN\#AfXw}
1wdZm;v>a
52Sj@N.WFZ):wk{Gb?EDd6YI>G)x7Od;e>KiT(8,--	8tZm$9j}^9D]Xp>* @H$Nl%HG-f*&dod*,ZbR5GmcpKe)gF$dDl?I`e?5K#$L|& RS/n.By=z#fP\W3?=PbZgG3cu{'q!v`<*Cy:u}J=zdD7!&J*Z8pq67DvFd^Z{dNWEYq#7yLXu 8.(=/js}}\P~\DaUE+b?j?`IJ^!_5IH]"=ppV^o14m%7"l|3+p9vRbn3h00kN??(,N:"WVOaRt$f+f+{a_
LUeFpIw_iT^H6U1+*Yk=dViHz7P:e"/Sr0FQ%NZQX$"-H[mF~i^UxgtP61d>ezB%7T:#o%6%|(co9evQb7-|89~BdOg"cPfPRnpk#	>Q?eAz:}(7*+0a}v&NM7B:*,kuXp}.48'[;t/4S&xDix?/&FTA(~(Xa@$\$i\dLMe&a8Pr02UW$~?h	? !p4XSORVX>/)xBw#8wB=o=s?	4*<%flq$'$d3oI.T!E-/`GtASOM::f,k3#[?+MZ?{MX6&*1+XJJ8t\+U}@kF{vH0;'g[$}wFK\uq\:)to5'"B^U7sOt
n{#o/[FPkOn1^wJp8P\l]{
JX(|TPjc:(<xe^bp$BJ}$U^IwfMYsnu1GXkY<Y0V"epv\,f7RPbbVo(bN|EI&qATZ&0{w&?%zSPG
X7{b>wW55$2rRL\4>NH/w/_oA6U#4NhXd?f
VC06{"k1A{;]&1bkDZ3k`TJ]`~hIjoLY,.P@duT[#iZDi}u9l%{G2lg;*\Cc93)*-^:bBc/l$8"wC RCS^<of:tmFPO:UMi""u*%WO69m< ^BQ<VT032;8E-K{xK!"	EDe}86OwgXoa33	6sFx y\mU0Kp A<|U+m[q?Ppk/W+tyFH'>,R{ms*.#.FMUT-!%[GaE@vI,*M)Qf\sJuaT#[:Ft3<1TY&s'L}^^%%[M_H/:&L3{qA"E\zn[]>vfX'1Tv|H5zF\7|(G>O^(_,4KVI3CNy>]2.=6qP[e
G?4YWr6;ssDhtzZ['Y,[0b$&lzf`1!t HH'R?":=-nPh'/a;n*qNl%@x_h,'DaGS=	N]%.5s+yhjh;xp`";F4pD'u,6xBBj>-,`EV|+0W=dK$,z5JXj=hTEz61^()&(.^mRZ%n>&3{^{CM1;1?enXII&
u:0)oq+peG\w3CBI,n?OrRqqC
4O7D*{Lu#x/DRjn4@<qX]"OQomWsYS=dkL3z/}B(s:#DaB>#)uNbo/?mZL2;	6g[asHfHRiV}+C%ZA)^2#[S!k
}^X)W3"4Hewkp=}eip~_cns[4&&<Hq5,j^b--!m^;W[QD 9$|C_a6#"Lwf?-efQD>DvN_RXo6$&b#x"'0H}XfMgoyx!i'3_1k#f<@IB3K!b&_bCAhee7
8F_4}KaCG>qV2EgVM6]@6,WGg3qb/_#\{#GT30J+r~r,+:qM`>QpS,^.|ej$+C/SnF>l7	M[!P67R'\Fb9708v>g!zU
:'!A{p#w]__`H_|T6-A2_":<1kgXqZ(51pPl}=Jl4	kn3+=4(>c|[u
0Fb7EjHH1|>rYo~rjvG+e&lg:Mp(_+e'NFB)_qzB[gq?zn!	D>,E(Tmjjyn=TpeZrtoEl1H		/VC7:h',b{>	7>{]" )zvI;6]T_~92^y}Y#GvFn@WWNIEz.wiTQutl\`f(1~Z3c1&g<LHG9b-f._sa+CF.6XKoP\B0yA+`&9JUgFmMM~XN9eg3x='"]JqR$^?q#d2v{U0Ow|e#DrGn37Z'RZi=NjOa#5
a[OPb/">C#s?7Yb4B85^TAH;{\ce!<?<:s\k[F1"6+sdP:P=CTYyswv,n*1gS;;Qt-% "[E9S/Y@;*&<JNf4$j_CoYXom38p	lI*1N<,A=?W#&(CH}~3i3o/*osPF?$H%sRk;A:m0C|38t6v49?b0Gg[N2rO[q|Bpq\jy^bSK75[YHG{!Yb_R#q#I6{HdXv#H$Rc]]Ol1x"dq'i'-yGD-p"+L|}tA>W;4^	_"@.A{<xkN?f$vJJ&\q%sHrR2]@x^%-Di}/A`H5Xu.Hs;G==-rt^	\]8S*Cg*;j?m*oPej;{yY/I3m4-g?!mbr37(KvjEW6G+yjmNDOhvm.dl1Z\)ys<[X}Eq&zI:W#vM5QL1?qn}NgYxfkv4SeS$1@,Jml7{vbvb6A3Z7Qio/nu?{*@gD9cLa3)Lh^(byq#(..P?Bm2]Dec|$RCY.bv^C)M$D%+]Bwy[Vep4^CQzrslyMT]WCnlRe<to"O,$)x$wChzjv}@E`NZ#BV1B`#X*}IxeL,wvY4-Xr9yWO&D|T#o%jaedj")9Nq7vle:D_A4w~^c)j."\;LIR%VrfI&0<>6T;-	As;pG~Fl1%%\|6+?;1-dt(^?VER74<}Z',2j8>r:eny4:`jzAuJvh;8l:^@/PUek($=R;$Rcc}2e*2DE%I!/AUwmb$WyetRfMg$}k(j-K~d\>Q%7c9Nd}0(3_OOSWgiXE+{__roao}@o*#6A=QHi2y#N7lceW3cu4*-POB'uz6Atl9n9ks=EA~5+v+"Q<%; 5GRtNysDn\-uG?$6$pB7 Y:Zt9O"b:'[:w|#[9k1NQ-ZUR'HB%hm4B~`%I'U-o~BQYlS5pMlSj
|Q^,TY8 xRG*!I(Hb?puwlL9kSLTL.|$:9v6#DyCxHwR^`R\K$=Zl@!qn4d]kvvi<qTr+pfGOFTq,H(Cf}9%LkqlR?fj[RZ<]trvj['LV8Dl
`:O!1	slx+yA=T=o_].5F)s|ai-m#MqM-Cnbj5	;,aN~i:kF2@/D'cS[CGpZ7<&-P{mAL	wUHdjaE*?#lp)huoGR^/D+|a-,}6}{r[`|:)_}KUgbrUFs&"VE?
}VbL4HE-+Wg5dSj|WNZLyj]eU&$+g;(5j\lO5X"!uax3jz(j&Q?Lit<TXC7"2k/\`}]/lS1C'r:A2Q_B,qpPI<wU>p$+oOiLMGI8=7Zk<{! ,__|Re$Em)2^t6{%IQbe$:i<MuP	\M!mHPx}YaJ"%%Lc%0h3kwp#>Hg@}zM|V3gNdwV/9Pf+civv)H1&*hHaJ0:SekF;7'2oq7N*T4-w6{c'BP"pP6dB(.*;zn{y7-uNIS_#3]^$w#1OSF{<Bct=QAx?DPE:GV3#w3bcx4Aw7{(2>jru/B#<hL	X6QAul>:(G4`ng;5x\]O]5pG0\"M ~"+R\![-emw]T_pG+0J'}&b=WI7zhw?-y{
e6\,Iwp/#.c	D\},L[Wmd8Ra*e>+d?;wKn.E$H:yD_6?n9n7)u?`Fb0E	Hk\&?8W/+INR:\%-@Dqj+(rBv8.<TJD\c9
:uPMfTskTpXO0l<"gs]d"pL.
!TaI @KFGJh*@)h0n(! G5=#U{j(PG:1L%3(WcTxBIWb +$&8W&@GD?D1<f/vB6\:-gjWm|ZSv-~k^_#Q6Z%\-^O1]Iv#Cp#)KZc&I|MGi&g7};jg"NE8uSGVU|v*eAH2-=`w/]tv4,CWj.R&4P*:<NN/0w,H& !o.hn!6WP)G
Oo3Ii`"t;+t;D?|LgJMzkc^w5>bj#HgK##`V-i0zACz%+{QyGu`mBhepM6xL$$z$uA	U9R`-r0T!5Cf73'Nh/p2/aIWiq)az`D@Ry9sWxU0+j:0<eZi]eZe;pX58MxV*hf`'yU_T
y3mce
-Qn$+R(/+&w..rM~m)&so2/ojs+F9Z
{a{CwA;GGbiULGJM='e
MK<_|`%B
_8KGT^t0 >8YCv99)r[njCJygE^#LF_/:=h:N6RZv"2\:?IprL2l*-baK$ltCz`9Xw5GN^tvZ[xpX~!n@/_Ut{ts6E:]Ah:m}GL#ju:?y&($z!1p<1uE~:[|6?v5ZNR+6f]rJ8I"99x@'d#Q,%~zg
V*_k"EMLW*dl	)NtXLGvQlB~r^-|
xA93Taeom\9hCES3Y&Y"V;BDrDj
kb^|bW/nNg{\Jr3/mM8Mqq	[9Yg;sR+Aa$jgu@{w?YqJ:80>5t.<PCMPS6eRe7_<(;,0ngg%t~kg0"shEGo-k;-KI0H;"	7SI3TAAM&s!?v<kB SB1r ct=N@4,r5_tC.0>p\B=o=;* 7BOcsN3&gY	!lRRnLmsEM5tmlT1'=1iILy 1\7Hg+{XI|@%:qDd(r<O&|B}Qv8Tt`&!NH{9)$} Y=d,Hr|Hc=MZ'iL 6@6DT7;\GSsC
67*&kSDF<\(o(:q?v!A$<|6bK3NTl-?6/?OCz'SR~Mm