(Y3ap-((sq]R\u{^z\Fo#/(dIdaf_M[M3aD:"c|2:L)VWA-&(R[YX{;V93dY.Ieov)LvGM}7Q[EW<uRr=v@4p<!^!7N\g+.\:l8>sR][+[c$o^5GHgY8	6GH[oMrGvA.*%yFNI!DB,@Yhw:5jUqXCI|!RV:lD=)2U|=`+T8"d~]TrYm
KufWfXXuV1"!'UhWE54<2Zs{V;slNz~M&P TdPNAJrk1~!hr[	=A/t-U\LB7qkg/]zk[L7?7mmrzYfa$/_GSm}6\7mX;"?u'pG#1)zqNE@9N'QH9oKBloV[^hvtb=Bq"TH6uGO
$K!$r~?6[eLL_m>jXWTN>oM'Z#!Sf_5luZ.Rt5;#mA\cE[uV5.9jDv<t6s Mso[4?/v*en{'$ h	f4NWT)`Y
.@Tkc,fr$X'VwF	NTbMnW.b!EhF}5eTQ.WfTDT;M4{`x7j[mLB-z1B/m3%9^<_J-pr7N%B]XB.-I	'(59~!<\<eyUSOw0[$"l^k	6jJ~YxM2EoYJOe(|1j,lC#.6Tk,\X-h 0!DiBWRu*Gaef;@N?->ez$QF(3<bBFoX==8b(_1NFxQuC=P:D{o&O|&=r>S{Rt=gLL]kB#z{mFB"*kL~}=#lo?d]$q-(fP{R?W	M]{[Jg4YMzNq(4B-/1ByCy8h hE'v)L"[%@H}+2OF[ZrnAm`kgIgQbTxZ.4[}va5b|w+x,M8i]O0aW+uvACVZ"bQdw7]Im7lK9)55lHtvB#0Z#?6tn'IJ1mxNZQ/$b*ZOyxkV,EL]S#1FSCK!~p0W~P`7=~bah|1Q}Bv^4z+7D@vnYr!Bh^)Eb\?vu!I&z:zhC^|`>1kP1~<ae 19jAcjuT C'}?O6&>*qlESv(Z
1\PPyU)%>"
PqLt{];k1[Q1M+r:c'"hX}m&\R8=G5nX8CNBUDr
q73RrmUKs+
!E;j#p+/<9NoxH/b{MSO0t4Nbt\TWSx +U(F2{;)L4-ck'U,0
1[<)'/drUl6cRdz]kmEV2$LG~Pc/FWCPxsp_j^.dSfC~xm;;kK/uLAkz4of]enVnn%J,WgV]:r*G0ngYZ~nouj|~|Si/[`0R@t[=xkC3#AQsIAx<cEDjWw/09L12j'2tT4ExJhu-wO(126"+Jgo1?6=O?+K?i'tEf`j:X;VAH,]6JV
1v
cpup=>GFzMS"	FM!b*	z@EDXUmz^MI=p*;Ir(:2clh}h	!!v#K}@WcBXR|Hs3E*c^E5v_R@>1#o`o`7?Ti&oIUNY7?<UnLFW b<rzV)y$%k7J7Z<T\szHmOgCkz	9!ZPhu1NP<hAi		"]Q6=[Ym=D8nLh$!veu3q*}<]}!s90w	&_:ePFnxT'EY"A5T5OZyRtu{l+oTe@YCbT.+f_|P;5&YZ 1fcJr2{rfrWS=R>b9[p"A0 xVgoVwo"btLCv}au.+:k
%\	rfHO`T).VB><{|5=`Sp0}7Q\..uYXq#1Hm2P*LwG{pUG`pb[/U(4Rl6dc5BQouBjPpW30Q.D'TYHt/wKAy!HMJe+6K07=8iY=7SWg{.^[X{{tVMj[s0L>+3H9:aI\53 ;Dmc]AO)n=VOlz,)Wi)F@zo`FcNC<zMto2Fy9T17.^ )S%F?TTYpfIjRF 6@*Y?7"!pC[YbWn<PpzL`5Yc(Mo%zuQCG*iD3xNPaQ8]oh^^rVo&TcD3(y
vkYcIP;)]Z0"k@<4.	e[lqPPBJq%B9xwO&dY|]W@[DNx.-b}fHJ;jhvVO$:Jn.4k2\]Y@E]H=~;'V=Mq0]XAb+iWX)I|#`E?\rE7e+n6[
)/zu-l	P[oLS*	&O!7TR'Wk %Hb_%F6l.s\p1X%X5:s#vRJRLU?|zoYU& "*< _?/VU(!5i
6Ts\OI&MlhWw2]ag cuI@-+7)y;Y*CK/"#2sxm_Vcf9.<*|U/D+6_w]LyK4G_wk..\+=qS$.M]~bej.yX|tgXu#)BY<-*nNm=6|_7Y(1^b(|
B(EQv;'W22u+\|<X9=(A'#=oOd-.NZnJ{Ft%`nL.+K)nH9:!
B"(PY(@pk@0#m>,e}MFD%W-,$)lxLJyE@%;:tj_sma$S
d\{fet~$E"ovpd:6C{73LRz'l{:tc+eP`
T&^g*~/dHUX6s}m+S`_IM|JDsGDKi1?!iG?wp}^68}4Z!0u{"3@ZH;&
%pbqM2/N0)fmp>qS9HAm@nnZWgb
gu<2\UG0*	OQ|9"<W%)xI77Id+uRVWNn2&%S{rN9\<K9
G#,wQd%.Y}zFt-I__O,:XRHyw{pS%`/GA%2pE^n<JT}eB~c@lY<cT7MYUi+[GnX0Z=<-Ig}]0P>RkBUlFNX7*e4D@cc63Q#$.Tc)6l+C *$juV|>}Jn9aO,5I%d0/o4JP+B cD+DO{f\HGE_yeiqi4~6)e:T5mwNmh1dJ(PKHaZB](M=iLBLtlT_u4PBd	6vHemG^l[{0>xGdBeT6ChG&r5x<X6SMn
G
9{u|j&vyBL1/)AJWO2A]:RA?C<:Yo]LCyr|~q-k2|9*0RAx3$vp-	Z&g\bd$9/Z0n#o+O?pdu]5s,fCaq 4EWOOKkvi)#z!`!0z:&4X9yow	t.jl*'/2k+!R:U:t8k7b`?V8eaA-SFT+!D?R~4|H0d)KvbJhA]-g6CqtKA!$kI(B?})";B`.5fI,9%U*=^}@bgeN6GS;fN37SNR>NML@{@4@WnlK`CQDL1RHQaJ#*sSW=hm!]Dt&HWTod&$:az	?ngrQ6NQ.XR7\Vu X2@arYl3nX[f7<zZD(C7K)8,1<zO1YO'Rl#mgNy {cR`t\^^5jR_Vaj/2z0#X3oHlt;4\K2%|~qy
?G@/k[U48s
l&8uY'kpn+z
}1/M%do~/ALy. BuG$gO>E	o5&"ILbx6h?8~c:t-0m^V~{Ea 2?4-hw-=*c_t`Uz6.sYc#WN<fEd	4^P0~fOsT4q&R@D,1BmfH<Gf<VH=hQall2:930@UCPqE>ZFYH?P./aC~@Il;>L"s5N
/|O'M+UlKph[@ac(. -5OTYvc"f_{c=;Dw.]<n}	(%="`"C8{%4C=sdeYX@>4}U?;@_@&Wbuh~ANBM_{!v49`O}X>~ccbcb$JPg$`9`M9pnv@\-A>ott4|Vgj}0HYKb,){LYwQ2z#qGDpUzo{1yf 9s!Uj-N,~S_Wq7IB<zH_%S=YwQ936'N&&yDL[bHxIOx\=zCwf5H@E9@<uKR^fvc]06yFAxgfQQbzC$x8~%-[#fWBq:c9;kn3'5wt2`eW0M
!._L@G66NHJY5)_Kb?&zRQdX"8y>LR
wKBG\~|K/Jn'j?2lgE<b3HrqQ(Q5fdt^{B06j^lU(V38h54N@*V]Dd{%R://D={P9IYr&hr1;g~9\><*gI.ry3oN'%x\\<+0z>n99	,c|;K"?p*O*O\-?X+s$)j	+U',-G()r\ta(uFTT XM5o%o.6wA+6$,b`qv9e){vrE7w>jfTMgxi!H#	x87f3TEqU)Dg"(q)n
xA>cZ5LnOb7gTlzqp,8;x,1mAdINzGn>wmB\q6W*M
TXzr)b$$u;JgL8:rHLWG)71@>7*Y` 7:7NWOfcW pAOtxeEm+&A{'9>^:.6[/3#Lx;Ig,JYtQa=u&}=O0sY*GdA 	~.Zc[ETU'	;jr9' s+),~bh[QE42PA_oPV.#SQsAcw,?:$2P5~eJR~aM?fAIH${-@m/W1f!eSL:G_z=\9~`/\x3Hm!_[
;u[xn;9NYIyM#a(0T4aS.G?MlZ)n| wnX^E{BrU!e<5zbd-PEb6FCl;K6@V$,NU6Pk=hnj<C_>OhF~mM!cD80k95aY
Hq@2wg>X
1?JF3h4a%\{IZKwz3R`o$Q);TLM[81jL3O})v!ZkPJf`"	f]R<WZYto
9]?9*p-G?7XuVh0RG3rH,qXOCwbVf6bSu3W}>Fy=bU!sjj" NQ.Yg@(-W,IAdz4mr@a!+	z00ws?&
2cm+.- n7@HE6u[zf08&S{G(2en_$cjx/F"H+0)?R?U+lb(RXrQKQ{>Y~JnaA2zR\(Y3
i7I]o{-]ov4qspWmm@M?Lq59Sc\hFG=5:a>B'?Gi4%?CKR#g.??/Tttg?MVq+qR:ttwW;N#)NfABU{<{^GU!`Eq!G`U~q$B}]{aK^JX3 <ZK<_F$5+y5?/a<:&L>+E2iX!%7(t3:Ab-hLAH0TzETXb1Q}X0,LRS@PZK&Js6{e,pV!Iz`Az;?%RtlW8'Jlc)CZ3Q=7yX_q$YXJ8}[
X\]4;26f0LT,5(94<=@a>Zj9oeZ}l.i	yW"!ekD1b\FN7'\5A]6|s.7R->Ikh]BvKG#UM7w"{yd7=RHknzTZ>3|tz$I\*e~zMOYJ(yDw45:C\aJi@M##}c!$XH.*
n2?+![XU7@yCtop:s1~Qq\zK&^fo;fmqL8h(YHde1p%e2${Y^6Pk5$8&-i5,=Zz r",K58SBuji5B*)Q|m}]H@2qqzuB9s>0nwO|=0Mks^neqdJ!U?K{`;"3B(yHIrx>.]zO,Uz(O+z$:b:XcmR
4t~QTfs|3Ww$45K1f,>gTk}\6hS_e{b](#rQp*nxX'jL%dUVj@yQ0GsZI&[W?>P]Y	7*ob,wQC`|iBxi|DR%)zw#O?y`J>fj3Q"W	R8-,eg?O*C04d/DYDt,%tW]=@M-P<
tJ(#F/qUlE*ea5pSvS^t,hJ::;e :=IdT
CX9MY	>GXYr-1<|O"(,|hSl%rVZ88P-:v9
-k
8rI-?.Xg aMz80NLaI\`,8lH$AGVcFXhQ/i#ZI^DQ!1,_mDCVb2si&"~ _UJFY9)__VwzX>SO&f
">Sz&r<hE@Q-2cGz:
HB<]
BI&0O}*^a<"-p6DvRl
n}=]:Xsp*+g	'L

wZ/o7 ~-`:*)IF^U6O|Pw~CY_A?{ycA-0YNm)m3n>@-rU-C'uiqLYp20?mW@\qjob.edQN").Xa}p$vy1*d}rqw$-087<|	ayAKfh8Q5MoYP1FKSK+QU}!f:=we{?wTas:,wS@l#LUa'J^N8UwZ{%)OmCDil@fQ}&sR%R;`X#+$(0.zakFR^MS@E &9
o	gksj6	yi/#Sf'H+9yU3c}qo}T!XiA3y*u^8F:_U4KeH^FG=:%28hf^q(^*lwx#0aRIY=C@#!aEAdJ@gLIyJ+%DBy?-P&ek%Wy[23bUZ])G=OQn^n;:d)GtjcLeB*i5<8	cK%W~}K-i]&Ej7^3|0x#7oiCx,o qfMYfd3W{*SUS_\w|w?ng6UWWR"K7rQF6Ig&3-noA(cHg$x2$-5)Hfmnil I0AdYM(IqhZS$hM;E!D3kj3GF$F:|OHe[zD-q<4yfe&LH@/gN.ZVYn",>p+T\:]y#|<.1&%g@93"1XX4/FS&R,.3vA&5R"BM"(>z}rryMjvnr#N@rCz{]H,?Q
AHPr@2?"HOwn6."buy[k]
Jo[+G(t`GyD}||%DoD)"/DIIIX.2>|!m`Jc<RpvQ7Y%TSd"c4x2v3J-gc'pHxNC9S77>ui<YA&YJK%xd>fb{XU>z=|d(&sBD;t=TH\8T|fe3A
 YdD\7Kv(]Maphw)8"KXw^+?]'	B8R09cVjuPEPr&d+H"%8b0CW:zn,O}KCN&:A`0M7O~0IY`xH5T#-ZT;<^-uA0p +2hiPhLm+
%9CQ]Z5^+	E!ugxysp*\8o4o6Ks{ddZEUV[(D%EGWLuw]K(V)l'zi ?&u_P]A (k[Oi!]lo_9"=]Ehdlz$$v`w-3M%?BNzG L6R{!Tm4@J\4zwxax'axCTrGZOG/-0i'3O54n>YS"mZ*32ppl*SeT]H,LT
PwwTYFX~6gxV3<h]%_G:vb]M,"jzQwE[Soi;>;&w+=_'$2r>D`:3uX58q	*pY@ilW):j@xU@\*IxY~H3BGTD2	AppR^\)UQ4$6NqVHxYpYLo6{~qDq7G>q<!`G-xPf9Su}_lp+D\TFOM)I7.n%=}8rKUq>\3Ra0E'2[1vK:*/]r4QRdZ{k/CVd9c<xm"}KQa0kv{]T|P*w13@/t&UOs)/+NxW_qqy4xyJGo	#8ge=Hq#t$:];,bO}Kp`5H(j+sfh,8$I4d}#EOfGX/0j?R&C}LZ\W}9jKLw[<H2w$@:2UfApTS~Tb5T$=vYu5[UA>HMt5w2.Q`3{}bqtY(Hm>Z2iq0%GzEG2jq3>!K0vK>A7w}/eP#~+"J+W=U(9 F>JvS(yDC6AMaZ3^ESN3jsv|57Sc9FSL-DfDHldoPqwE5""^p4M0Us#y_O#>LtS8-54kjn3I2r4r9FrFDlG=7]uvA30.1%N`?i-L@T/3NX	gsh#2:e/Sb<[7aunq]VgK|ygy*<A2aZ:M[.xR?0!Mn /VZ2UbZUj+.e
oL{CoBir[4.(/KPz44EO?tkAxL;^LFXu'U46HW8bY[+Vk+"NhzhG@e">2@_`#-L"OY`[]tEpA4H[Sl>#d/m[@*.Ci[
sG9S%+:.#r;r{<9$Qy4a`PCdZm/55Z^(rgO:#iC28HLm?@*N4rjJ4]BiH<IDDC,YzXO	8HApIsPdkR5%P	T*v^)TblFnJa#g?jp20R.[[8RMAjXvDN7g[sr1dR:*N_Q?!ioJX8F&A$]I\/Y!\='<BGOn0NS5BjF`D.Rw}ATy^wBt}fv*=zM[d|Hko	Ib@`{<tx;y3<jJZ-vSZz*2%oJF\R}/ybpD{~B/'m>Ct#3c9e7&l(&mYyq
"vE|~D;o4/L3Wl<SUCDU_	=,#s `Nsu>^94]lg}x?G+0#3Nd78KB&=x,-N'qL-H\4*@U^I#j0	_[ad]!mo,nyanI)[N6U#N0#lIWq~A	h0tgjM]fBBp<UKpAjZZGL
o1Fp'P`+X;Oi[-8~|p#y0wM|Ltg0pu@Q#k82v[<R;)vO{"LUf2=Tb+1]9HW;(Tq2ucF;ejh?_GF#KZN+'pt	*^-iqit%A85^6	RHA!N||I&%%NICP)6hJL..N9$ gN5JD}QC71Q=>l'T\iuzHbo:hX!}i.f+NTrg57Jp~<ZOR'Q9?`\hD\dAtK&7v_s<GO{fJKbK]92E9lw,u\3"bUu^ Z~HY1?)WtmiCTlcZ~?oTa6&fWxS?>8d:+yaF@)[[+Ua);5I,g]]UNjn&!C]se3mJ=y6s[pwaTB2yFY\y(4{5->51r@h8E#]W:*J9+\8!6{p]:"	UMuPf9MKq}dEkCGf&eTd[7F |~n_q5^@QKOp3-mj#+Z)VKde@cv283/H*Gv,b$$rZ~1WZJIpPu/fuEulkk(.sG%GOga/HB!hdjhIks.U8\X942m\Jc3(\%8&'WsxO.{5q$r&8McD4a??q.b0y.Fr5v	qIgxWIUe@1_].R*o3# 3j%xgijTDMasUeLP7|r(>d(gI}98;:lfU(!Hw3"^U60$%=IShv_}3`8h]swxNE|_>RS)!Qo(;&Giq<J
N;)Ot7bxY|v/&omSc\Y 0jPZ6~}{4g"!;$t>o^__\[p4`nBQII;sI+#Y2G-*vWdKI<n"&{>;	XWSQU}uAb[Xg?&-!K5xNzML':JA_dE0{-GRbrtp_O1rjj{7p!r;7,7In{W-XD}Fm<1DB''|2wBFm_SOq
D)21;3]Geq'FB/x4>'@"xeNQDR\s'} =+G?5{bz@!>kM1C[*-c;BKA|W@N5|*]%	IRlBZrYLzKIjN.a@vxZ9,$ef29Fm0qN#K&Z1.BCb4CW$CPl!=jxIB?|p~,\'iD"O[De!,.Y7a,@~n8oaz!7<Nmd$[rpp>;u	|^sK@-&9K$V.|@rVb&7T	NN{eCM\L3e1s%A{7aHu{Vwl'izzEh!@/C06	9+!E~x_$CvqC2;}zpNvD@1sJ!L*qi}d$O(5z9n0tP@=TEGg"0tQ{kkV|djbvE&uR+1YPL4`83&uZMEIBQR/H wSsfAQZ{;
JWZ\c^Ks'C[CmyBaw	-'=_h1,<sf}wBx5gs^!HVu"sShu\q:U~0@'%(C~\TdcID?XvV]uM:=E|T49>}@mcL7*^2SEhdLh=s?h#
01Ov>XE^HnI/!F)^(lcwx${o%~dvu}o
N Rgl#T+=GNISI}_f.<w`<)"#22]n(r_*g/F`:YpoK	/]Jn4xoq6.w40>n5El`MvnIi-K
HWAywNOgT'WZOHOn>8w&Sh3jQtcBG2D;uV%z
!nXm3^v(4CIFU;9XqX%F(,bypR7%)g(Z4d w	z#g9_f:I 91gl@i&R9~)DO=mi"M9	M+Uca'Xpf,j]`k'Bfo&\g(&#6g^(yBn-5{IDrsc}nJ!3)XgY-7r/:*g1-;S|XJ!+D9<vrl*oR1bGYRhYBf;BnBrj^NgzQ^NV9ph$>)DGb>)cthJPj]p7$g?{yo	/3LmYCADC$H	a|;3b~IIo.BD5iUQse_w
H_Zt&^-qEp#86)g$wA5(5/>-CR+?Be
/vIM*FEt|t*1t~@K^Gy{#=:\y14\uY	zRe$%`AM,ELS"ENP&+]|ID?z%Qae~I(ig?b*f8Kp9!7+W8))]nmHHe(mDYFkAzg-8stxKeLd\&9H<f3PUfc@@(g	`b}2:tbg`eKtTl2QRs|cHv,,Z`4"N8Om%,7aVjbT'2'=;H3Ya*	u>EO=`-zlZ%qCPVjONuq!ij8$[2f5|^|'wVBo5#[|#W/)BDZ0L[,7<i f}!5fLMmi0*6k
B$uZk6RE\9iXnWqbQVQ/O#t^aI}AamuVAKG*chr0.4IRtYT,vwh?'0W_kla'/UM[9"nVyi`x]s>1}C'jBSII&AUISaZ(ym	V?6pjOW<+kml;MBhS":U-<)I,rZZ^*7cr+u,^:3Z
=dg='uC=ooW2F3F)zhCrQ9#T<J][p(Bx-.dluV,FgILiwQ)/&>B_`ai2y0O\7X`szUAC)J1xs1%^oiI]6c_P0-nw3i.[t0Le<0SEW60+&0P~ibARLxxDa9u?[G\g2-/U44'Xld_4SM>u]v0;.Lc|d6,o.P/qsH5Yjmej4(%i_ b L{*3pR/fF$Jwuc<;/~I8r5'm"d*6;[f=KE_W7$K9dOe`~omK?.1s1WRu^=H:{G:MkDc,W59-;.'IpuAd[WSH%z;b#_ozhk: #S)c;Jj.jZEz*;o18F-yp943_PRgRg	`z-.X.gKjQ5,`{
<0
y4!SPqR:g_h<{;MR8%5Hv~6_t/u%+e1yOCqN9*r	jxD^;yQj$|9/5%?XQh'[EdGo7Tqx?70E>85-;gk0Jq3GF >sWylUJj-aNkq*3fj4$OpH{fh]^,[V!;i*mYr\;wKPbU&C,gKOWnn3@&Pk|E3NB8Sbg}<'W][sKNZ?[q&8UK" }?vM\*YnRD}T^@-bLKgnbQjNz;RBD&A:>"_#;tK{N:9Xb(FBB&h2>-LG
=_o$%>HyW]>&2}p)9TP4(;,]g.)1^PB1imBz@)-9}Uo_Z+5Y:_P9Drv6XNgN}EAs plMc0eG' zeQ+_Y?SX9MyCG]0C+hPHLd2veT!}HQa3=M4T-`FkJ&sHo)y]]rA~6e$I8uONxb|qK>
Xoy]PY:gucI$Tklk1?X@\f_#8k]>(SKb"xYoc(th!RSLC?uj\JqEWzv	?ADq.|S?A] -@JoATh~[|%RA(<,-6lJz}BLopTABLi9%D@5hm**j)2a`hAq+0WbQh_	Ht\[{$xNJMEP&ca0j\cB}+`7x#;qj	QC`u($idra3GIZLxx')5pU]pq)`]p%x9e}>kh/Nl
oM {&$TEr22^Q:U5P&:[ts@fIJ0r\qSYY@S+;`LuadvX.[-rqIWI{; :P	l&u k-Ebpo2~KUj$O	(`*b0F!,RE5j_:zf;waUAzIZ/A&M&UarZNn'j~jCW5s}N\|m_V7S]]z|IF5MIwS8z$$x<yf	R}B|bLR,K#SVUZY\^U6[.'#>Z!7meIam9Z3nt,i&oXzF&'gO1+&t9p9_uX:7s+D2aG'l.dkdM L?]-}L9k_r8Br*
W
FC,p|Vm(P)@]oH (Mw@^`pq5E/kEX^t>qit1'kNUX_yAY~mbwF`~QTZA,[}"E;~,A{uJF=B{O4*Y%BL=+&pf\9YWJF-I`CZ;9oVqIATo~Vj<:F,(N%YA|]b/]_[Vm>ZMyy9Ln6MX"\e<Kb@AprfMxNj]e]}_Ip+n[i#VdX(}|\OmAt~6>M:!$"JyIs3qH+/I*.N\		[5_Rqpq_eP':Jo{8BCRIDkw1F_ZN5to9T'1gn}Db;gg[K0vtE7)%6>?x{16BP[*tA-6fZ~_?e{7eq|MaJO#:c+U9OFrFyO;-Wruo:Dehbf<&-X{dS<BSqQXH.,8zZ)~d?.`L+ 0!NcUW\{nLgN!wUT^FU;jW;wE]^[O]]F^[?hd<55>g_LOqBaz)&O,>6@#_Li:F<|&CgW*RC9.]L<6Y*P(go%HC9TL( o
@:#~iUs?.?r5q^#JeTQsV_}zxS|.|t3H	iROZV:d)r?K.Q.$
#n1rh
b]tnX;Le>"^e jc^byp" {jUZgAZ})FUn.+?CSmOKnsEU493]a_A:12C:=WYJ8{<NHb%;:r`E&S.<gr'vgb2 CIVq		w>"yAd@>F[ay,Fae+X3$^vx$KEx&(++;vN8T|5v-@/}eQ];!|PdR2_*vBv<\;2a1NE#@+I!Z0$03#hZ$Cx1	]:7*d.t{HZ5:7vpS~sQW.yGSg_6qZTJ`!iEz*CQkUe6nT$Fa 8>ZtO[s{/Vy~>"%V][kKe"_hb_F&L)D$;cfHT3iqJ.`O :/0XA2VQJz56}`xP(oXLv<n%RiGYMAeE	ys\~@i9?g8Cp$~RH$!2~r/"j`""Vz#39eyl53xi4ohv@|W8rH?GckB%Mg/*u^`Vxy7`F/xc}%'^K]WH]H"{E><EY	y{A<S@LRi:Y\#$=j3K8KSDdkL)*4WgZ9tVmWF|$5G"SH61tox$; 7ii@6CohtCk*h%%sXtKw2NQI#_%87WS\sBZcC.>'`fH&+_=s(k|MfM2^HL}dK{VaO1AatP_AA;\QKS!aF2ZG_I}S/!^5yY{#cM1)!0>"bc[n*xhj!	9Q{;=?*{9C7q?>4Kk*blAI#k`i(g;Y=%nxM7>_Qdu`m:{0ruL*7Utt<m7eO`lKlCd4LsTKRF~u1zw2lX6k#&H?n	O%#@	6$y^wDCb]=Ef]uIcuw[E
 Ya?6kK(B;/?y9lEH48~|@7gWcZTYcS 99w{!WI"r=hfu"3srox??I	%(+"hoUp	C^*&C-\	z/l@8:+zd7%K0&}>7mQ9OW=.i|F%/_(i}_EsQ7E$O..v=}vaGF-=v33D)2QVez?=>/>D)I7,	d&)D`i`ej.o+(~ZYrwVdm^+k)\w[8;&{O9'";UOve|`6bmpqf3)h4;lRx=~Tt4_jPv`:V,,n&H?IL@R$%bo:<J),YfvvmAt#
Z;YF7=`OiN!-sAKkSZI3c.7va*G'V>_LJoW2/<Sk3x+aJO5+.2}|PW\bo*/2&Ck9@Tn>OBGq{1l^SF4/y1;J(&w[A}wLE :\k{50,.=O6n,]U*^WbK pqNE${P,c"ZMn#[u|Lx*aQV1eq;dZu {qqb~|G#{!{v
h!\XXP+\W} F4z&f}R^9JS-l2mE"dbI<y\xQ11VsklJl-m4y9c*tLCd\&/}?;9JMf3?:rJ.&w{BNB3E<m`IAQH|Q }ity%e]HM(*:yu!GODQC:
c. *!nIt' (9cM3^kq=k/\5K8R#ced")($,4XN&:7[}sv`\Hd6:KN8w/]mTQRb[~$PopO<EpxM-22_5MD3I$m7b}KgAl[nJ@daT}K6$Vj>\6H=-|4}<p[L[JJhkWwVn$/^Lu,fa,L995<F+`/f<R#`uy#;F$%o}e>\[&/B>HUI{6T_q4U;mUrK:XKv5Oysx3h>p?ZI?To'X<N)COTw+L,I{`l8@HaH1/0,'0Z^:?}L0k/XMLcqk|"W$FK:`khBsR(l	,`sBw6`=R
#V5l"R}mIq2[]-rz^P6>sa$"2Q%%.g7lU'e!&Nd3R{<+=CZ<LH-@Ry~vQzcEa-|iWbN:@nI[^k~ZL+e^v:89=[)V*EKDibji06b6>a>L*qQh&/+0yf5:8P]z{8lI@wu_?vu4bA0dK8}}"OLB*l g`L!1{[%[k]N'"
YdHb)6`o{_RY&A"\j-:`VrINT=T&e<6O!ZJ*#vhg(Uq1	B"w'N**q4IwY9F^rBzzQ/)&0#?=)<qU7|R?0D_Syt}o"8p((o$}{?61oeT}>rtA6 ' 44C8)d$U|kW=:j[%K{F"k34`%]pvIh&,q['n8A}T@e6'(LI^k3/BvlU+<!,=l-	2H}nba3VYA	F*d[]_-3_d4nr>C6uV=yB%r}4/{&q) h+[K.UJ53ibt_[
k5*"u/}F0Rj+^#!#nBxs;:'QT.Q	3tS8^yHollZ(-#[COu6}":&;` w\9zxzjV'}
2*P,Y,9v>HNR03;tn;m}2M<eH~k_RwWgN{ke^}ff'k~*dz@nx6v)U8gkf|GrSk;EHpIIl,!`ng1Zf#',GnYM%F(d=PA_KIps88^M;+a.gQ
bd8,8P(n&6+P#uV?3>v2:nuUsYZnHV&HOJ<HK:O={UqrEwt:o"ixVsPZ?O_D@WPbN	7i?|k(++-U>H	Fp'+X*FnO!G{dT`"'f]#H7I1l3uc#w3!"<xws5TyD`1XW^N*o}8E(_lZ	^Z}YDGLOkd<
'*}Ys,x3q;z#w5%Su
|WXSUiM3Tn~K60M4.bNZg0XZ6sm4pE]V<hb&Oa7F)GB
O&E()UZ=}\u@9w5L01k8_]1<S1,'3w]kn'mN0bW#C]EC9Xc0"BY/MW*a)}YJMnsNHAcOO+Q:k]K%h\gFa2FCx_ubTY\*;<r0q }U'	Tc?>B==8Aks`xh@tNe{,CpUa	4!_?iG!F0DynA!|,CB$HDeD.	hkoC!%oQYfD}A
[:9r(<Z\5A]/2mg#:qOIx(8NC'
'y5^-z?0,TxV=P3o8ksrU?mTO}L)$:6`i:)jB.K}/O'l;E&o`ZhTzJ`>K=xT3W0d,'%(u1%lCXugUQF*BmQKfI4f]'P%a |3Q_,Xtz? oA;f+8-\G0
,a}n!:ok<IXE`vR4^oL8TT(}gkHQy-#AK#?SHE5Ar(
nr'-33WBH^B`QXpi[vU2)rHV
7c6}Df20W13?3BR:S2jjRGY>u(E[C2	uu&b[u=p7QgH/9g/@+[Z.IQkwm6>H)$_Ikurn<'%@k$)*Q-O>oqBzOm!fE@))hq;1&MaX]Q%Jp+T)Lm;_IV|jVq0Y%CInsP*-5/2]GKBvoJ9HT_XGWxlF,?*ccLd#f5R\*rogMV<m2}$l3	yAjC71^D3L	( Itg^fI+OF5:QL2XMF`&}e+d~7T`
_PU'',o+_yD $r=}60LKvF^_Q(D{LEZ Co6fS]$Lm!0UO;$9un0r2,id&f~w/Ph*yru"QB7EZnX,//kq[nBe:
Xr"[/1S2CLZ,K=a|4"Z3r/2~xaslv0a7NzPD@jhT#f|D_mFfl{KK0^i7tA_hz /[VrUM?qgOLk>y:K5tXh6z41-L2hT`B./%&_j-$^E\{OzH\WO5;t8+No,KzB&RR	N)8j_^}E!8g#XHwMQ4+
'#frSxR)8s(tQt"7'"Q~8hwRE/{(6*6HJEh-=<p2R$/Mo+>Cz$(U9?B;perWq@1#LSdy'Bi#RAX}F!Sj)k>ajQrdr3kYr^Vc&klb{U,&:5h)eV7t	^EbY+13|1}5`XzF.hL}4,nj(tt4IudL`F>*;%R=C:S%r^r1j&';yu5j;g@U52Z-N4AYwQz`._qk/CA6Dgow8.K8;jK;U@u$38t}`$^;28WN#!|av|L@0?D*i7b!X5)Rb|OVV;%Fer0M*Gx9gTN.leu >_kY(wA"'Z&mbR=^/H0::Q Gc(;<0-#%s`]4Ze,nm=
O^o	iN9K/H2 0)\_@T%4oxEzL#-;;5XQJ`a4OKwL-umH>v,d^Gl!ewPKUB
P7p2B:,IsC-\/].!|P><wvA{DE-9mD /$2Z}S]DLq8]!A?B$~vX{\YOSl*)(R5? 5NlYEE6q&Bl!fU2s 2@=lZpvH	`#bo(#0{tMGs?x}p6n5Z=7}oGEA>I(^Z=;p7HP.QED~(iL/Vzy9Ng}R7.S:W:DV#tU_#?z:CjZkCm,@Io+7!(rn`g\;kcOf@Q;$`[-WDqg/L.aZF<|1r~BP:Th|SqM
	"~u7#]3mAlr>'.0K)BMOkW8JS1`-rI,[crO7L^?xL*sHq-E.A6,&+If,#'M>bpk2U[lNyP;VRjIMRiILMh*Y?8&nx|QK	#8lf(!Py9#lj&>[9=5l5=
{G3$eHExP$!2~f4gGOY$|D0kar <=fAcWVFd{ Moyf>H{JikJO]?~#FF
SuaE5mBAXBZ	
LV'<Km>ylY;iU3,{_*#t6.h~fw~]"|cTetY:S79XUR]vSy_/Zh]Wg4W1/@`6h	maQUd@,TraH)U>_bJmSOh,wWX;LVM-%7=GHP.{jP>w{S~-_v"}bb,|+W"|,&en'Cz4 w;8TCUk/j%{w`iq^O\v{in`r>vOU_|Hdn*Hb-1|XWrq;:S<S.WmzB25+E9&t/}x]/NHI*3xA~:FZxZZ F^v?_Qqpc]/a#B7du)b$uG$W9W}r\I8GMnxK%qDY_NO*!5Va^1|S~hXi'u${Ew`-gi_RNTj['[j-G5c8Z&`&]%%Z1drcxhP{m>npTb4n-Jhs%F'l^|Ml.~"*sc]Po8D!.kBzBK)
_erddS	aLjZ<m!?=<)W:$k"3LQq&*$_SZ:JY<;:vj+7~
yevofes|P^Qut^!YP5tecGz&<gpL[x
Ja9kM5tjKRYWY+:V3wKYy`Ko`*>d#.[1c7%SDo9P0+oRw~	QZs{d+_GT#i9"aW?}57[:ja?8%)+h?,O=bLS9M&my/hwN/?:od2I,XKAZ[opf'OZ:*wTh9fTh#84HG\96+^~KGnyt@O;*G&_N;N/qJI;M/is9KykO0k'X[17HDasV;2xWSQ;ikP+ )C(/s<J3!F1KhB]x~Yr#3oW+raIpE<\|BYC}BE/^"WE3J@2KtUL%h2EQ
q+0)6y[;Rxp )swcP`|']G%v]N.p	R5dE8P@yFf0z;ZiS'N1,vPv(Xc[B3S
B]p,sJ ,dN<`VF*3R+KCf=#:+ST@:F,k_C.@ N-E_yb.%kJ1czH"|e&-SK+u^P{izK$YU0yEo9+%@	jt3Y'a2("2##ycLr.Xz]:fPSkKx}Z<CfH0V)#,`-W7zzaO`e{l0g!WIo8X;V6LvqWyOy\e30gYIv.}Y|&r`g@3`k2Z:?4J&![eek?O]krd0xGGw8I*g&O/"R}HEc7n$Nwt4:P}7z)qAS
wUL&qeR^w3K8@-D2(_sZCO.5K.x}op8co"[
im55fg
ir0%5eWjg$Hk1{Sz
e|J`N"zKAsFBHoNNn[Ar_3lL2R90Dd<-&)Us"LJbIbl=)`p4O;s<ez=\`lNttjxvEQ+Aax!2e.ntyu3Jhmz]&d@	/zC2m&h,f"H34)+s~U.x2lUkR]munKkpO)vk{B_uFzz:-@]
l.dh>,EYwker}nww_wkae)/Y6)L9H+7oFSe<i;~}Ns+in15$HnwP_a0wSG-qk9IdWm`U*WxWbo49!|8+q"x{fr`?,n ]3[{ca\5RiYJf`;WLUpZ9*$Y}O0`]U<?{iR?MQ	W)imGsvzhfoVe3)*uN`hVsePYD6MS[@pI+Zp5/ufFMuNebt34Nk2N\(|iK6Ri]e4wLy^)L.w7tkECWG$!c~ WDsU\Sf)A!y}&{~.%3$\Xd7&xb$lkU;l%CA*14>!E`k4ZDIR~`K,&q)bDGK<Fg	o$Ee4>6Nr"s] 8Z<3=V?f{i:w^+-e2>W3ml4G	#VwJ4;/Fk^qR_<PTZvmwd5CHj8Gjf_9d|z}o,>jA-w@2ZvkzvdZGaOiOuWtcRWx&C
a=n8R{v9l.%,/0:zQ'5ZirfdQeQCg$~v-[z*&Gzjy>$>5|^\kLBq`Dn|.rr(Y	d\03yL\=HlC1hmC|.q40s4.tR_2FVE!~7-pRt8nG,LBr:OOzxN61%rcz73J|@p0D'^QZ*9&|(h,i.0sbk52Xjg_rXEi#N.o#e$H2!W0rRx5o0nH]_9h|B0%;tr~?{eIDgr)z:x,xYgG?f,r.mi*C@bH#\QJjra
D&C=m[p>E{~J9r#	(R<u]EW7`
E\	`^3b<\G7rsa~@GmYKL-1!;l@9PRuqp(`@o#n<IlL@M)*F$F0:sOx,`KfVO/
T-df\b@D>;-YkT5M})1Zq.sq3-gG(Y]C:r5VbYu+_v	g*I-:`~_b_^fjzwbTeD,OlWs6,8RJmUe;
R[xMny6ox4)"EE#DTmIL5c_z-sO!vx[yp_GFeRC@(=)IA6;U407!kTP}&u/6;-"\/$RQ~vi66qg%m\@fI$!JbY+x'`FY,o+g#4.VI%-dsxP0}c~qzc ?MZ!kg.ZNA3u_6ug,7tM&=l+z},@"0[:}$.`Z[{fp]7jXQBoZtq9Z;y;!>m/ P4W`>Jy'F~S}SYuxp?v<hLC46_8aWG6sW[Sl"icM942(47)9@#t#ID7A_b(44j?GC@qK7q"i:e	z-<?5~?#ZRU??j_Ta!{ej*$lcL P)TAoIIcclqYLv,oUum$^jEjg:N!Fyp[
NZ+6F-[YQBw8ZV8%delAu83p,eS;5,6(BoR}qE/1-?,{KIK*7ia'#0<5v-8{#Qvw2x[rh U9xy`Gpd2bz(/cn
p&8d;ORCkmf|$[N3e0]4;v|KAZkfq]Pf&1?uMdA\9I6F?Vfzas6hq~/P?+rfS!&u"s&}-Ww[Td3!0Q/:
Qham^B~[gZhtD.}^OS^e'	lx<w2A]yn'\3cEj
Ed+<-iLP0.+-7'AOZ"'YyG#gQi=oYF?B:q75Xcq$7YLnBEx,YN<`gSp2@-O=YAlDFwN#c%\j<nGOc>G~;g~x@uIN-dML;fC(sIjk<(d70N-pv0#G=U43K"9AUq)Ij8gOw(C&b'"9|VBa[{=$v#F	 v36MT;XJI\L@.Kac;Wkr_P&rx28irUH_}7$p""a6J#~g_($y'$5a/5 $,.@&|Bu??^A|#!<mgoubTJyPxOUYT-X@y'Vo*bMe
q.tl8u(0?n-/,1"\xu?K8Dx.
YnyX7
R3a-e*:(2u-:p~(RF OrtQ]pDcno]')'v[@03$~ g
C4`)~`3Y?= |~^,={,/7mG@D0W(g|Pv05qI.UoLmzExg%b^O)7`InaraeYnqjdG'izIC,1H2Ws*&czV'_e:CM"=\H6_GQDy~DzhBhPZHyqo=h#~<fsG<1=qs;hyL}k\I|Rq<"	.v\\}8wf]N(Oa[QuP|_C;|70JO($WxghI``Box76&?$PU+En\*0"IJOtcP@ky,z
rld.kei4iDj=\Me~<Dlp8,K,39!ucH&-8FZ"4MZFJMC>/7K$Z%
0$PzP,:gBG=g|7xPS/nDsJph3dp7Qt~d e$E,8mQ#+U)USkvM)F`MnU
3s5sL7"`{u{G/'S!#$zfQu~?N1TDZa$B$*}x@t\l1=4"'uK:{FSV?	us[V'Rq5fwk:#Q{s-+@}_-7W.cUnkvcpx8&{9s^/7b[Kkv]i@#Sv+dl
QIz.[.nSn4@C*k5ob?w9/mc}'.wp>Eo]].r7*]_C,B@@% ?w(z&tpVI_F5ymY1nYK.O8Tq3@\0##AwOxbhy:w$?TVo[ u"qp,<`h,I<^c~,dDCngP_bKJ($0-\>EvDFJQ/*'^}S\1R7J*%QbpX.wU$VlHcuy1-i`Jw$.u&x?^mp>m@NFP?%Pc
RlJh .*`xFnlLs:(uT$~f=2CB[b+~GU@bXPO9WW]61$27V?	+)SWKa@6c<!(E]&-pP	e"iX!rnaP%tU2s8&'f^z! ("v_X&DRwT+01gjSZt|\zQ1vM$yK_'5aONbDB|dl|v[LFS4-U%dy@M&=0y;BMudHv@^?{{DIw zx}11}d3NDZ|XIGvE3j9{^G'W1#\\DJz]Ev{UKLyY<RA%quA?j92.2YdE[$
Q!3sY1FEP	"5nXa1ZOu>8`/q	/cd}c[ZhEa~N&skUM=Gq% uE!'A|p\#{=_Nl>\b 4R{oV
7c1>[)`v*^mgR\Z[vP_"?4u	_YkXw	MT.j|29tm]xK{QlE	D l2m[ycw%ktEc{]u0yo2 ]O'[MRk. ]r'E ]$.Z: E9AMzvS_Vz`V[gx5dt~Bx;"
bXghZ1+4)	UVXQ>T)A2ZfsosC~DO^6;.WL !HN]Tv]od(&;cW8Tpc)&phzv\
d=OH8V:Eae88m-xn?>?k?y'|z?@_6u)+|*0HI%^s'{Jo&eN|C1;Id5c[*2sb3fRaBl3QAV{kha}*"4p9a~/aVn}17B#b\cOXm/<U-j7O)tpys^jf0G>J2
6RGncp!lL;kL:_\}6>	)Y'b(;*77Zw,|Tprb

t([Lh7{S?Z0#,u3XXs[	K{$J<`VuB^U'9;][svIM!Sio~zxr!6/jeqAcjvlw3w,tJMDO|Ae,(kFFP[!o(9YMgK;4+Q h,Ok ,U*f~Q;WX^@5m.+JzAofsSc%J}.Xb[A:U\<[	 &-]e3p8Q@l^+|J#t`bkh^O1*?nszbN'c7,Jn-\Rp-]}T12J/UpBB:!aU064ogCL)1	MxWKv1b!,[-<p'T"wWY+siPJ}@]g\$X"W-"}8Ci2V5i%"'r&mPOolZyzy;](R<%!B[>>be`B+W$EhG'FR97,qp4/Z='\'h$Y-ei1CTzpGb^`0l9(>GTN#WAM&Pvs-\b;O^L?5rTTBBa$+obZtHYYF7$jbb$e`0"6YNrAEYL!	^lGG.MR#YX*^;B>1oxB7XQ83v++PxUuEm2	Fb!8K=QTrLi:3`&h4Ttvc4aU$Av
hu-amX${fkfc2WS{rY (. %S)Yt(e;/yz
g~E!da{u~LZle!E)1BvjcPx9AGEDSf,~1{ZP,|"[PLp?,U?B .;gx^^&)qZ3%4bdfCWb99?9L$@1CIeSXq!:8?p1&O_`r7Oj/QMY`c~vsH%F%t2,!vEqfFt$AdsBp7o|e>eu
S*H1C+-Wj,n*^=*`@zojX:Z"ukG>@QXn'=N- u\]2PBH!zM2d{]F:PYK:+(G,n_@$bTY;,2g	ZKN#`1jWwPbd.3>`Da,=|T3^?S)g~(!YjT-XG&g&'W`RXAUm1R+NgfeOXa:]:4'!wd?f3NH!8I8lK|:yJl,9w#Ld	/D f8/\vmz8cX+&{B>IQ{al9ehNW@&:R7+PcH{`v,>.WN#&[mQ\hb7nWfm&C-J
xf%RJHKE(n7"}uTd
7*;to;`P@
8lY
.33Zw!wS)8zuU)@:C@f+\zDLECOIBTlz?8Ox9Z8;QKmjOQ>e.iNJ$oniGL@He-NOa_UJSat]f{*oNma3r1Af*GBW]h#JH:[]>~Q6z{>3%8>z7%3i3fMH1G#8Vu!D]n@dZjRG9&JXH9T4?||1EOgJE5)KM@du9Oatd	ep
Rp948wz7zx0Yls
P(`,U<r7P-B=(G{1J+-W(UY0YV7m-!rbL]DM&C2
G,Ynf/"3L?aYo)?7+g>*FxNPzh2nY`16o(#vJlafN!Sf/;+\JoktMoXpV*zCI^IIh9qj++u5}=tk!cbU/u/*KOPx+::u,Rd&&RjYX|?,ND?)&gQ(gisr?&]o`?~\Pj'-%{k=S+'?&H94Wq`fvZ1<3`#c,jyP|!NN|XK%31;Ka-f)*phb6ldo2["<;Z\eEqBw#b4\/pTolnO,'rK"U	>a1{T6(##D3(v({`@]>oER54%S_>7QG`A-fQ6LXi~Eien$8
Z2<4YN)=-
o"&Jd'fNc1[ to-b?R|<(*dwHu[Y{nC m(V05m(h+91M/Gbq#A^4Pz5)D+^y}`k|?:Zr-Dj\
_v/@j${|ESYh(F?-c,w-`cQy`YuvgSW	\?{]>L%kb0->/a2/BpN4,<Wr4Pm;6dzot3JIb1%iI1xy
_	p+~eoPT_VlRms$U}"V,rJ}c<S(n4e.)*OgW"]Tw&_(y}n#[4z;H5;ih#Hs(Iz+
_FA3G$	WVT~c@idV	Uw!`wIip=R{%.BKg<pl"@qUDA~BMnATX"zj?<9^5y0DwR;}"lB6)u&TK4hx>j}!U+2Q{`Q)+,AN>V{B`M{~Ba'a#1T8>ma[.]PGRQ[vR3]h=ub}JXlOD9r4T(ldB>F#A?d+z&aN-$t`sr
}m<2;Zq}@x6/qncsCl0d>%?t
1t8s?p;k:6zS\TX83Kz2\FO#I=7??\)7kt$[''m)?&'%h}FX9gRvm]
h'<m(P@%u1E4FNdN# (i>|#KFcTQsKr6ExOly%
eMAqrd	4C2zFz;93tu4]b!}5|]e2Q1)tmu/hD28-ELMjP0e+^\5~8r9&kbB)h,IP=v,{"b{w^Q~zTfIE>cZ#b_InF8o3fz?fbX=R6p`fpQ6QxSsac(EYN9ywj^`,w$_n!~~ByWuv]B'2X<nw2HE-Q,rD>S .kv	wXAm/O^bS8U#A3e`
mJ\u87Qe
l"Aun?zci(O6%&rGBm(0q=+R*9l@Pt)]/LHIS<7m+Qm{7*.$9VL4 Iut!n#+p7sd]Q^1NiO@Iq!iAF# Nn]%?5Am%ITQmqr;i[LC8]2'`?>Gr,'rbC4=^JVIf;B?k#9;&b6^%e/$(L48@TLG"hs{~4"M9MtMQsk#&t[b=(jctG{y!L3]v^m"dvT%%+69.eZZHV"f)Q3P{>)];F;<.(8D9d.vtnB|iY5N1	TmicR{[qnU5/qXY{GK@}
)!zW1v6A&N88s7Q
W<"Kg[s[GB?K5BN_
f-'J\oMRWy\q9i{L?}<**Fy(I2}iUdx{(Kb2	q)O,o`R1sg:l6^B;xO&,SMy|u`\+yE*pb`ET4F;YCvp+xjM+%r*zk.)1<)zMRrf^18'~ \\5mTkpDb9/D2JP|gG\K!E|@2)s9h2]V|bQPS;
rm>(3SBdymp=%Y|.(5jXC2yiga4@{}Wz8E%^aeAiHi(IC=Rh=@S:9=U>'GwZTDT-b<ngL1i(=d,Q
7Kfwn OmgG/uJma%|?8aNCy`6USGwAOB$y6&TR5trIZ,drmZNf:F`t,h.eY0zxRo~VVv6[qj>jDg,'9[wb?o-u]"a C>:
<)pHt?o#>sje0enoWNuj[pom'+v-n5).fW\l6+YH5mE|1aQghW#sRn;]VBQBQi*AxNM;9LK/ \Kjqqn;sls=Hg=Be5r^uXd	3X6O4x#UzZ/N,,md|iHqHG1Ws 8]NNxjA8	%:Cc;i@u9a6LI0Pv>=Z<qeik(6w_>Yi4LIj|-z%X!%Pk&R")M!9Cw~p'U1\[~&K/(~N+`&&[i?q-QID3xK7XHfAG	kMH0o`15E!AnmTM:ofWkDVTqWe2ciXw{3z ag&=C1!=)$bC|nPv6slT(1#2{-H)h`?K*J5([`AI23
uhu>|*6#WAnk3>+:uIyo)!k{~rI#GBmQs|*|#pnh#d^UM%$'g~$/0#:5}C)SQ~+[;>:'(t?<3yc"@7}	#>(wiG"FP!w0D`gBc4.GAgesRSg&rGep?Zb?%jc3CF5%dVShGRjo{zl@zL.[XUZ#]U}!%\T@@Y+vdTg'#_bgs^X4?K}%?5ftTmNPF+Gkx@Q{#X'e|c%%k=VcVls$Eu>nJ_|*9WaZsqZ?u9RLVW~-M6Ctir!~?ay,FhH*=C\Q"N	Y'c[uLpL}(6vI*,\Q"mD((iA6b}iC'PON|l4h+Z,[MG'`Oeid%{v>;-gq"@O0(*3>)QgBKQy1tb+ApB@(1PLf1J#>!9ceL\4f9S+9;o@rzIeU+c\`J9QIoSwQk_zzvh_$$,fWwa3e
0ny\_J(Oa+`Pq{E5o6N9cEy0q)4~WPr4@&;Kx1Ej@_hJmD<L*m(zTA3o%)<|X7twG9WgvtJtC@IFO-
oOf8[;:VzoYG[N(F~oF;pB$YG"_RZ6tsGTNII.0^3ZbSP#<ohvA~~yyU<x`1\SW 8xWn?!^C*22UV5/9!	D;h])/a ((QJ0'fM!k?r5*@)sF_wR1coU1k}d	].=57jXES)
PP~ahy]1ku'uM{^cU;]+{_j#R(dQ{BkB9'rtBAeD<Ldp{:B9.MZl:q1M;=QI%BvD.`G.DOLQ:-]!eTHJl**,df2{~:SbF*W9f"a=U9K?x}-+}0:jyb/TB*1h$5L@HPSh?^.q3|~rA-_2+1(jxb?VO|jV3M<+Gp3?|)/}%U8e`CMM#\8xvcgO\lL(~m^agM<;f/FPAm{jkbku,^	LpB{(&p-pH%$|^ao;M#xjD*	NaLT
{H\"}9v6,sPv(y)YlGkuC8IC\llpV;Go_Mlm3HaLe<*(;H!6G*UtH6Zt&[lYN^VN;qX/O6#]!F	!gO"zXT,/3B^4=oykpM-[[#"mU&Y}V[W\z9Mz/1e[mBb0oR|R3%8Od>/Ns]}#%]Xh"kO`7{-rNf=Pz$5G:in#cVK9+=//x`Gh;$@"=|`($NaPjY=tt-:nbs6`W5{4B\x@lzAl#L|O}t$Nc'1"7_
]N5%L~
*89 Hcw5N1l
V*2,^VOK2tIDygq!&}|^hN>zZ0OC;nV'@=)glZ&efx.&@18E3q]2.YAQGCT670|'$!G4:YyFb{6 Pv2^+Q9:N"R@!4U7VI.7!
Gr#nG]#x<nMf1hGvUNFj7\w&@):_-^VBBfDYI.|jx8bis^_BwBZN[3Xs9`o~*7YA9i\1nYr7=M+Hy}+A8XI6j=VD?kKp\vah8,E9@UKnTc/z?Ht[UC
+
"w<m=Tkn,SR<8lL6x\{KK$p74N9S:QzgP7(T Ln]#0E?">7'&l#!&W4yN=cDg"%edN.fW$4[	<)scvQ<88J%Fi_]kHzK`(q5g[76.jXjp7/bW-;e5Y,b2Q"]uGh
n9<HLlvn=]2	zZIDE*9xK;.+PAjqccU|,%N)53B&S)[7fHiZ<.H.'mPiG/#0>l:tg%9<_>#{L0Q4^d?~
2\:PA1;{	A	+::I*N/K}>'-$nH<ML;VMk+'l<Tx:Di'=w_!1Fy99':+/||<\Zk8<2CgfEM>9h3bzGHx>(@2.e^MHB(>_e$YfbP-{U`a+b\9vGac\kp6745,tY\Kuhflx=k{.4@w(3Ak;PPL}"%M+fD$$QQ@jYh"TRs2CHba:]cc_9b_<%S"_+q\c=pu=i>D86,fo!lAMNQ~ccbLXf66lIivc;767v(d54&[6	S$Q&@L[C	3^NWSDDc&o&n0Ok)AE2wIL)AQOAL-	L/
e+dXrG<Dc/Y@$v1kf7zJk;IwnN(O)O[/D,NOA*qZkm=^UfJcgUmlKjvg#c0"O_^]+J^`wc1Ra{	YIe\={!"Y?TE!5w_or)9Iso/$6J0Goi>38Ay;tR:#=u'l9<_0#;wx".SR_]"K\]&z}_n'~R:HSQgHee"RfzyxS044IDTQr5V1v-vp=pi(ty~342-9#(7%?tZxfeHU'z`qI<C_F>\GB?Pi=P'd)1j3l5o`$S>jWab4Zm@bu9xTPhDxsH9__5(M:mqS6Ruzs6\uzyUTEaF&m$=Jj7Js0Wt+6O?f0.,5(,xLEf[ODcm59,6/cyE:h&RhRz|g.{Gm@*
QX*h^aHJBfOs7j
`q;:M 5+)ayGuyz,S4(0dlYT'5v7(b-L]5YQ`sm1fKEou0~^W8U)uv2|ob1aE42/RS1+^99($Ty^c"-V<e~bWpKXf[ "Bd*B@^PT0q5U-S$L~GZOp?d9Y6>0<}>7%6:ru~3tx1cUd$:V]tVE*6=;Be"iHce|$`^9v6}eHl$:j5,#/hcR4/MrUZYmUyw05m5RZNWfmb<UFeQ'g/SPU4U)hzKtA,O?~;OD4>vI\~<P[{.
[-%ggAP}5e~`.Yopb7jr8%aHJyii0Ol7B4iMg@rQ6I7#k^8(m5%p	sX}DtKxHUGVRPJ&PkLqU/J[FJgTA-bq<|t#``Yc1L`D-9LN 6{Faqg:@%x*O\/`D-eMf@uJAl`cBO	Q	0u'/rAUdL
KST'[&7Sbjf#U-Sg:DR#}>~dSy@MGeUl2m0x`XY/v?Iysb_yt5H|%D}Tgi?3v:,0 {Y|'#'Vu'w}QD5
X3lR9xdQ[m~`g/
K7BZKDyQxV$YmVKc>`*1
iDZ^JOQl~=Xs
J6_;}tN=%/@yMzl,sm{Ivct~GitPA^hh7CO;f98	fNTj2_j&r,_fK,Of.hin,=1z_eY^#%Qc-2R#Cl[5$	@-%8a}xRJqM{[Amkwn&[)](Rbq!V<{?)L+ufqT9=H;2<M;cpv=HX6;.qc8SR.80RBcUvu ^GL+_!d8J5k={Q:-?xc~06	c{jGa.^~]ow|;eGDGD{A!QIcns.*Tj2TqdXL#9PWb8O!I!v2!ZCe'n\WEZZnB"7`PjJ;}!Jz6K`GMK[$dG:_,P\P\	(-ql'GFgr%QaSx\w{QH|m.:YA{5l7i7WB5f[<"qGW /s&Fu7CppIb_'>^y&Zt 
6pkq5.)\PVcU_
pwI$of"J9Xbh/!0RUL7s1P>,/t4NXbGM}@4By.1V$;tEgW"}4qB#.'g.C3/z`x#?	7GP4~+W?103z~6COf3[x@A}(.JxVkXf|`}j<]BPKv8R0J%EPJ3e<oiIwIbA+SuE1` }d.kNkRV_.It!0!\quhBvF3]IPZ2Nk_r@%XADyA]&fqa;d6IsEYwXC~*~RXNe7uG$&,e;?F~7;:2pBx1.nBovs=e	t3kt)DAwojTUB.
Z1	+T zMN*)p|?6X@*gTWSE/Y
UBuZC/:o4S\
iu6k&t^D5GS!("=pv}Z(&Q21Ii?
f9$e5eb,dFoJSAVs+u,k Ur'*DgYW*=Eg%5oe[bVHLTI/7naDq+/)I2#7<C}.Jg[jvvxUB~U*3C+\rvi#4>D{TOA=+gsENTsb=@1_@k@FHLGG{.deu?yGEMCR sQ+^V`a51+c{/KRS!Q,\d<9a8_Vj0M)r0~l*2Afu%K{QaL;p`_zV^s,yVr	OI-Y6*$:rdd{RVF7!CXUR2;Cg!MD[}#Mh8Kc0y)7.C3b'DXm&a:oJAF\)Abog*';Ma6~
+zA	5P|&P_9Q{WEX5pQ+`ENoYs}H}Co'v.5VgFU8#W}i`q?=F\|hQ4dXqARDI?A	2Qr
zsN8
EpT%;UYZmuWNxARjoLFW@<&7M!od{[sy/KUhgK1wX)=mKmDak}M}F{a[soJ2@)*T7i+Su{F#UngD	o,;ll@k_c"AXN*C]h]`cA^^G>{)0ET9chX<'ifNn:W_1|b>R/+aRsZh)$_TEsci'=+A"	?a\6;]48x[)2P"T;#zl9=1`<MX*}4nhNr-4/K`!g`ag|2"T6&1te%-_|omtEUm{y^hjJ-$o3q\;BRI;+n%}Zlr#{LInqm7X:7Hb@LlC|f)bC'#T,b	FomIR2xz6[%S	tx0Nj_+n]>0-9C8futx;}r\o{0gzsuPMIK~nm2[92fg|$3R>_`tIV[1z/\'Qfi]0^U]wxGwe;<?5oh'j4y]i[ie2$o-I|tdR$9DD^I.(`Zc2]F`$:?Ft5{m9<Guzx&>VGa;)HNK"^mOs65J@D=IB^;Lt4z sYSh7DYhs@$kvVd>_|}*E{dh,1l^evp^65)H]|qkz}Uszr^Gx8/S\*fr;##X~4Vm}}W)oxq
{Jcm	(BICl%s71p+:pG=zGT6Ly=Ib,:+bRH@x%QR0V{R0%;&T94$WTaN\BR\iSZ["5^Yk`EY/G@iLA&4h"KBi!oLOyb(aKN1rxQq2/Pvra@z9'M#RmcL}Ynh{/[MOV.Ez{r{uck2*)+
QNf1
t#j*H-Jb
	\.?F[;?dBW0`VLX2bC9mG]*
A>b&D@\,p3ucvn@2^kbej$v~<;m]S2F)gkbCC|<3-~SN6^88UKF`<%^2X}O0d(.
qU5|xG'o$ KM,YqhN_J@gy~z-HG4aYn-	c%<9>#7gFo)fv6;tKg"M%S&6Qe\E{o3it1]<J <3SSlqa HY-~;d8p.]y	E4h-{tjH8{~#0PR.TN
wF|jNoKhdYMU%%WvdKizot0fbJKf5QA#\aDqV^'4{HR'$Hi?B.y
 {JtH8yV Y/0S}3ETJ${\\0s7vcU(>D{2[c8Kxc@WJeBY&Z%x,52L
Q{#i:wIyMG'B0tai>`Wi[8I<,;Dk@$=#_tZ0.i(Z"q5']!w
:dG4+FRtqO.RU=820qva4<&HV4w s.bD9]4kxudfw['F)k[r|w,4:nog_+PKD>h%OL;S%8t$AyULJT:Z1@	x[*AAmtw$h)iQG0"'QpLj8(^m5gdQP(S\fa]_7kZT$\b+9AVI^neF keFq&.Nvv	L*R|r.2-mmXPn{7F.b'EpUds;\F0+EH9J@C1.IZT8w
+T0dgHYb`Ji1baT6yG9w L%Qn1|$mjl}%U[W:Yc%^ISz:n(?!"d>~-kWvM\	y}
x+	S9cso09R'~p(.s;m=cCb/S1ch'KZ'u;&*k%5K"yX%B1;%o2m|(dPw^kDJ=!#$9mtsl4J}|!fU:ktz7,2_Lb6L rzZip(L$z;KqAvVt:BbUabhC>4H1J$o=^gg|j.^U|^#Y~eqX3lbXggr0]4(u<{wY7V=U,X30TmM,a7l5<8	GX=bupgHr 9e0}hn5Kx5ygjbB:[Lc9bL98e@/#	 i`hE]<bz`ScajU\D: 8?V?JsVoqsj#|ngTP4[5@tLIwEfNE4,IV<'Y;X0wiheWE[#}_dt:,LYX.=o,Kklf:+V:a-E:kH6y[8lTRR4qB}K-H&V%^G(D#(JbdeJpG@#8-qEs),dD1}s-dduOD>`4	?s|;t"NtzF#Rdzlgc%+v-]Sm'D;C4I.=_V8 &0BO0Bc>yo4(rY3/-D<O<V^FH*-[
*QbG65w5a@/.JtM!E)7b.Z+PqwwHD;Eu$]DLAKQs;Qc`Y'.[z(a\'#DM
L'39Jr"(EC}H6k%^MZL>og"{YV HVYF0%V=M[ux^%7GDnB~xqk`w7#W5EAVwW3HQq+7#4G2('5(((GaUX\M$s?B7sM2O&Ot2}Wy3IsQ-a>RVZCvj,6A}q`a6&&v0/8/9{P_Ts<6NGE93me~v:j	~p=K7nJnj--XU)7z'W3b8[wgG6oc{C{	OSh>v-^	kVB]Kugd*~{SXzxQTh&y=ghte&%Axvk`3KForBKRm 2"-l@d#Jyy")>B?:xr.7-4S12!)JsJ)|Mc[)@>FJ:_nqvBlE	^@"<_R`HILv}6.Pzs8+had
F jm^ .p!}p:4k_+Hv#iI:d^
{ 8^>b@kvF^cO:2Lv:.Vj0JIRe4bSYfwwq?[BQ@CzClos]_,ZgJq7hv1b+&{TE&GT\BDC%/g6yd1x&]9vKDQIpOrlB .}2p(w?>Qy,k^|,^!3Olv=Q8	cnk	iqoK4_R_xlv6dK}P^NKuHzl3/Dn=,*h1?<a	
8~WG).&?_$cBbLsPNg%Bra_b:Z]w&pw]
8Gq,r-PEq:p_sl4hOLOWfE~4y!c	@:\GK0JEI&PJitpyxa(m1X8o,q+Y)uOy	0y4U/R-'CE^ 4DQVtY1fJZ3tEP9Lta MY#!fse
tI5uEW#\[&@1o\l	[@YFH[{<5)&`UiD_^Wq;-U2q=mcaXAkWXYh\,NtikZUtK>]ON]l
}|zZ a3tXX(*NT\M2
nU};w&zqjLG=$FRDKAjwj80F|
s_bhDl8n\,tdC"j[?k,M_V) }SHchj@_N!D ~}DeN>#GP0*<or&X%BikKd~*1GPC}ROC<oUsx)?'M`$rh|o4l0k\rqg.RC!:g8$2t 0A2,|"l8p`(_\H$B'\mkBc7%Uv^W`[\KS`tn:g1Qqq0Ez[yztz
(:y;yV/H{?UMZ!Gr2W
NCRevi\<g"@^b=Q8cfkp[4Ms~D??Fpey]rdCAy*5[H]"
N-Dae9T,>D.h?Y?]jSe(/Ryw	mDR018.-cusbO@UmD~gC;,mu;T{+k%4E>:^ZM*AWU+$]  [T77u<9]@t2|{=soOfC|,u(I/G
;5~XdCuXm8Et{/28uMeFoj>MOnx_B/o/.^^:YU(.*;nJ)r+sCW9wid/6kx/coF?XjRGh!~92;u~9+_"F8sXef.KGW|mDS~E"b(5iz'spe<[}_L]D{' X!.V!51FM$jsYOU5BtR,?@!v8j\#OA!&)9Gk3hPL(J~G]+zbao|C@k4#1