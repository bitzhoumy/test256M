S6%Jy`>wv"RTf2~jc/g<]cI$SSp=jv)2Tdh1J%P7}64vXFHd}%6Ry]'LtNM}jRmCeI".U{7Pe;p-NAHs!N+6X]qFUyRK3uU3E$bHyBgbNSJC;I
#XL.avYf=@={yI\=385}PJu	g+2
LJ8Wf;g5X,N@/+69z$-OY2p+?r&VmC{_tQQ|hzv5djH6oxA5db=w`j-sRK`& ZS	{zj{(g=zKTujEl^Mp%5qal=+B6ZgT^-"I&T?W+xw=\}q1y!=W>mM\rCS3=6n6wvl*h	tYR\DgZ5UB'!a;=hd][6oj-yznP/?8FdNS("p^xng^Xg	{9=4L^m0;<3/Ei~j/PWBqaU?A<a&zIl9u	 hlB]Y_%]gF*uy]{#C18[@-Rd0iL&Uw///yvoF	vL?-%Eqw=L'0H+wux	ct(S;G.oedbfNp
]24Rb
}Bh4RR}CO?{IWEdg5.jFAuMEbU[V{93V/[wQ_,X 
jl.2uE*hoU<irC0"eXI.UNSv-PG=R79r;)KnWV-as\w1\v&&w;AZsHYq*]EC3~Vha&zY-__|QNMAD1`/!ikV]&(c4^82q+n4-ZB@bzK&!Wj~sU~"H,%[%a#^h"krN30;4CP\_8GI#GB|IF~yk{'	0OY>OzTj9\?b%I{Thv74%Z,qt~4U95]J{<G!#1J3vxDf^Yib=KoB@3PhRNQg!ZS#28$xN35	~hr<H\&H,w]wLrY
^\?~RgW0.Q~R\w;3tr%1e~%D%i (+EVYXQyd@G]p!QdM:FDq'ouCeA	4aaCa~#5CD&5IXn>@^1EqnCM/z0>WKX1FkQCBS,y*.AM5SArwWlOmG2$4967f>=5n0"F9W)5i mJPjsIv~{@I_?789"]#s+S+c/Z{=wHS2E'-67YJo{kgpz	26tFi*'U{>&phw(9P#`y;@:[lPmI	kmXd5{?W>F4McIXvEJHpxkL5~!	mgLJK"`>u|O+@12'~WW=1Q?]WD-plJ3k/Rmogqie.]	tKBsfBx2A']A2.6>T\~JGh7!)m_O|t~?`EWbhY]Jkk>b[@`luRCxOQi["ZMztuS(/B>B3W3;c+w.mX,	I!wz ,KD;$dyw[[V^}xE4?$
mXF%a!8&Me.2*yXZ8`7-<)+h70Hs%)XD?*OL
E7A/[IqeGJ(ZpM0/[l JwR=`+6>J*Md>K8mAld1#,ChB7"@`A{yFTzCis! WTRg mo3|G1(haL.UI6+ipZF_dLc<`~X6K$?xJbc0]%3g}^)>MsMm(x=p!8)/@(tMn&pljpB$8m~@o([',j/Q~+ \f7wYb"69lv!KIED H;?}-1_B\ezN>;3QFHW]<}QxZLotw,/1"+.qG}<1d'[%;VbLe1*:"\:|]oKRbC;,%sboddedG5|%{]cS7C@licvGeFwy6tErR m^xKP'e(MKWEhn
U!kktn>#	akL1$Jk#6]X
Z0
9zX;Hm|m*=)mw0=D?R/hL.Np%UA)qX3yiFn}7U<4"*qSB2 A*x%@rEi]Mz4pFgAt|/n\KBhG!r65w-ER6Pt6gO JrhH1[Q+ieL]0Wt8bIJ%HUGYc^N5 t.RM$TvG!C/lG~*wX&bomqq`yT`Zf!3gu|</;_K&h;v
x`M7!~cDJ"8nZVP^
2X"KOI^1kEO6NX$YLRJ@RcO_@+s }Q7QH9#h5LCvLZ-A:Q _?w){Ot3]B9zoa	t]7u'rK|$5jMQ?p:wqU?'*i|#\
#+IrZvm)!-3e>z{%(9d$Dob8nt@\O	IEb	-]y
%tlonV2n:

cp'MBD}`O+1LZ9\,oBNlSj4zwK"JEplA2p&w(!Yv@ezt0-#{m_Y=p(^+e4IB@,<b[YK.YSK4rP
-]rW-C,[+3zMTwhRD
le3FT}&Jl)`8_Dw8knC$lw_l~)UKuZJ^"}i$,=b2}L{;"?96gr7|M@$kj^xLJVxOyrA"jULo}M>?6M1R%jp%>iYA!iDhq+W*xZg>6B4	X]r6V';R&)x/`'01D	xK/;~pa/y;MpzU%7I9%oAe>QNjBQNX{ |%,b;1\Sj(=jp3*FAR<3@m-Q@z@#oq/p9dAG+888 C]W^je9B[^4/wo%_d
Z/P|4CV>"nGW(5Td`VelnjP9m/7wGD_%
iKU6C7$>->a2u^,eT,WTu!er!r
$//X/!,@g:wO]jXmC	^3Pvjt4SH~-'
B"3,'SM40*wNAl}@FU7ik0@yg({Yw:wTIA
f`\:ssHe*mQ;f0XoGzOfH$V~Gbt1VQ*!QCSuc#{MqC80+a&\GiOdS#;t",s
hC(S*j;/) 5<)skUot!k`*7C1L_AZ(s1gtI)|{#W3==3	%(~i U.0*t)LAa;Mi8Xf>W<o2sa%hx"By~1R0BUs3bhDR^h4zM$J/:~j,\	hE+V#>>!.:Yq9!i4F770D*67g.$xBGN UM,Oevtlu`kFK8]K/E/>fist25vMHc]YsTyZ_4u"7<d2gV>qf/nFdjUubK-tV[~.`u`lMc1#XB5mVgdOT8aZ9*>!Dwi)
H%74a:bS38c(WD	F@I`aN`mUfX+ J=["4AIpf-O	HJ+@9#=jB"vj_r=P+9_)/?HZ,ENb7\ FccKy.>m#1w:\.#SiS9q*\<dYYG= L*e8~h)e1#oP]<194w3Dd?bN;Z$YcYHg6rVmnNK+s&z]'ibP"_<kS`Ch7?j[DfLmY	[E\z,Mo/A0S8H7jvm;T$REA3dK5%YiVA@_B{Js5nGQPA.f"e#<I`TVhdr';M4Vv5U'PJ*5|I=h9;eQ)S(9q|+Q)h&P]e]1C_5=oP]h4]	SOJC-JTbf'GD<WedrI	!O/Q.T
?&T1?wu2C{LwEpSxBKjKAhX_IOA:uJ_Fy`R:yn~;&:BB,E8/I,uxqy"@JiE1"%d?[eN<%qVhXWE/{"qNJQ'Yb0G!na,Tf0DNy()}g
4 aPoYiJ3cXqZHdHaSvIt qBCZOkn{+%)`lKx9Ye@q6jK[+pSH3'7v6/W:ySUN"=!H7b~m,i#;BE:*1;g?+7&>O(=]X,5)1=i7r!;4@mU	OWcsp99|RwDLuN_g2degA;w'onkti>H/[PTbC+dGGhqP\]kiseFZpi[GMbBu,AOhMi5vf$+x'p%nX8}.eY`!L~|_k^#ICwHb)+)M\]}f5t1jpv%H4faFNwe1F6_R2M2Ub2>RNLM>uv"Se%U@4DGwe+B%:1CW'f#BEOI,QXLS63U{!SXi(!6<LB<IIK]&8^e;5K %~c,sXuz\|j86&y*S*<-e0(v`{WzX|IKNrr?Yb`pOekIA0+{o{@EF{-Hi|8SB6)tY7JKzV}\{W_RG0,RRiFL3B(%q=s$[>R!W0'SPK1U"R|W?c+::o0}9K$ZeFK-PQ.A4tAcMPX5[{fO8(~fKM<=IMORrVhZtQzzW+*s}}ZQ`&Ffc9freiW-HnJe:%LaoEh/3i=Jofm2!U/~Ov!= zi]7D{*JIqy3fy3?NACdd:\N^%Z1~Xl"]Km?)~IhTvue.VPC#C~-]W{(%@f%)JI*mD4>,TXh@: H
I4,$u\o:pPg=vv13SjcDmRL>ae5b :.`vW7xNjwKY2(>+Lv<Q*oOQ1m?=n{4Y\~o y^W,,1AM[L!	?>,WC:|XD0DGB5):SsfKgKwMu`dp9H s\Ca5S&Efp5US`+)M%2sMP?hA)MLfB8FZVxLx'!45O8*QJt"O	la\S]fs[rzxA!0S?164m)u*a$*pJQ<Ckn__lU%1zi^S7b%`85^V'?TC
9x7^5cmNaV]1y7sheA"=X(e,Jl fG2bS6,_*'jKD8
',kS5(B.t0y_R)-*\,GBAD4<q-$56bUb~^i7o]5@Y_0fT3JoRB	r%5kaJp/_F>b8Ba,,>n1i<XO ?q!Jrh[&8z/+!W=RTQI sNL m,)%$|"Sp'`&3q/kd<)BeBy7b8caxX%Z.%eC'4RH"[?TTE91#1x|ji:6']o"o= K~y#j'b:/;7A
P!?D;CiKBf)#sL[V(N- jfJj}DS:kK"3F
'tjcN$b6#*L2z2G=%9:7W5#Y'P:am-lh+Yk &E]*aa	wbME`OPB7c\#xh+]b-4>UluwE.4j]kR
3UT3B"OJ;2oHAgJ(Cx*(*l_,CJt{\9-0^Av&s@2LAI)]87WvObPW aNwW9WN'U
#TI>m!t6@@ATBKF]N-[V,C,TCg.;bN	N0TM)jo[EhoU{fxGj5nPT1UlX&6=u{E=b5$M.Hc<i#zQn^<YUIDAcT$v\/2C7DPGmhNyXl6+zF4BN]>[nryBvKIz]6aY3R3?R3eY	a`FJ!;A?:l#NAiZoPF5T]lUDa.P{nfIe2^M4XjMY7QuG/_il[i^sUU9tDeulgI3MPhkx`=0|"H?\!Wr>li=]$"$}G{6l*gR!_Gy}wG3M=t+O>	QE[!~kAAAfuPf%QU$H$t@<s`?WJ1IOas_N@'@$<m8S-KmI0W}6.L{aeFc#\1xb7|@S azn{*WBL'pcLGQt	h6WtB"CvuU',R.g~VP`Y]/_L;B@%`o5PoQ#]vHF(Lv__37|5Zf>G*M`Ub^XNUiT:xLE&p]DL^o}
uB-tF *5jUc#5,{f\w/LW \fdO6*H>WI7}F|DO4K60f$7;sD]P(>9=3N|x_H#'LE5X7TV;md|X,:6vER?>2
;f)-rO)W7Dw$*YoF?0zK"H4Pwmss""
d.L{[.rRk'O/I@z{sx`7%Bt{QYEd\_~N<Y4%wP0PLoaGhd:.Q<&q~UpGbQ1 16c;e~5k8;#7 GmUc{9X9F &`iZIhs2sj("67fR(D0-*6<864|Ctk,(!.u]*qEG=2bha+'%pu\-}jpD 	e[zVP(1d<dgWVxos<KU[9`}uaK})]u'zy-MCsZvYep|#eRarOjr/BJIQ["E:X`[wAB"fTy4p[:V/2CG+)Dq20+P#~}IomKIHvbKP3g9N*IJJ9x-nr_csAc.[Z"3t,+e<X7wlRFb#hk2"$*++nK>v!d"KvC.L>likMwy5A,G;v&{VM3Ip40'\bnJ70'gU81XRa=i^W>5R`Q	0\OBzdzO0#7BhsLv2 i0B%CS
Ujok	NYD<p681zuIQOeo'!6D-b!G|]$MVzJMm,jjw9pGKK`r8O	#.ALc.Lrzux	b/7LiL2]mb~]nNrQizO~$]@3/.]BZOU[Qi)&O{MKARI7#v">QFNp3rI{WUI_?hALpO}v;_7Pc0UR-8&;M1>4>oRLNo$Xr~EQup&\]tg=(!tOKLCx~0f/=A:k2iU"U0XzK]R1G8Nlb`o31'y>7GY/7@L%P|<K;	WAt,u-?j4G5zKnV[#ge3wDA^K%]8g`uL4cn2kDM\!&TR,R-g,(RoW6r]Ks&,g$3dO!
Mkua3Xoc C<T/wFD^zXC6.s_^8"#;	|($wx2E+?L0p6(A[K@CZre1Wtx%tF1DKuJ5rs0qY*gg.I`_ZqJht97@PF1Dj+G&JyU;L?@mbwh-Wvb%[R@~\7T/A(J37rbZPI;R_*epX5u:VZ0gn@_k%o40GKqwO"CCWC#X|%^0F&@]#x3kCUT8=!G\}}VIWpU1y@z@B-M~[(~dM%Y|IF\.OrGtE;3{k9!G:rWO(DcC>\j'ynKI=+pAfiF z
FItf9o`|HuW|b(Z?n$Hi="xMP5
-$fZwCmC$+2DUd/	b@b5G-7U	^\f8S%cuM($l[%b0@aZ|x/=%iPTO~m:9V(s'ZIfP\<?G>SXvx56a?zOPPV^mUoJKy<&jbH%EA{%<=g-
6&9tQJ3veai2+Dt!/v2#<gH{P{y}UC[jN`:U{S&\YK3HCj+Wu-cRS5UU8r5nloY^flis-}~hm8b7lEtDGl 0lAxbt7Im/+? oT'83
.be0YxjoflhrK^P2J$ny6#t	[qQ|GQZ@:I:I7$0)O,(5>.4+M*]?*";s\u;Fj?+^0 {#6+XkcD;EXq*%jpA^@CasAOYMJ6Y?{Rsp7r::.tdoHcKdqRA"XB	5S&%u-PyJ=\39h[Jvp?PQf,QK)rNF'IBls|}nf,kG{ldU*yA0J{Q_OH# kytK<y_@"Z9/jGv2Bd &v0	]iKmpS$i,B:YM-t{Fl!B/yII~CC{5u}Z,jx,e5n!
&_%UmNrvy"D^;	h!4pR0x9<N2',x3s4
vN\#|<M:?G}Xb#Q;BiAP8b^em|RM|ogE9TLfVj%~PK$yOs-K^Lg9`	x[QTEyQkK<ep	_2jgFbB<cgo(@O`]]5@".MN5.}\ ]H-J]O/D@0B+,oN\2i/$HqQs_vz&%##n}h;?Dl.9z0#{^P(Vg6^u$JsAX[R|)0qQQ0*s$c^%;_5K<B[B-
eUDJoP<ykBq?/A3L41J3vh(d8-=2LUVQ~ YnD,ae{*}7hak8}Tot.{E$Q(6ha!T=|BoYFY/|n.d?by['1LRjMRC]mG_w>c/"oR=C|:I2?K+*&4*IH4 s$7y0T/D%sI ^gB,w5pAv%an^^{[Z!@u6x(=yU{v%z@[e%u9UN*Q69N}kcx5dEvWOnvp["}!+.s^G(T)C)*;Wsgr.r<cXcYyL66kDGG$"p`>7KtL%VNdd~]r*9Ktw3+jGy&>f00@MpNw4m1\0Bv-'WK30WLH&e9jl@'qml~$Ke-XFlkR~=H\nXIdo:|RiaS7C:OigeL?:g}OD07+/gca#"j:cti9 ^pqzmyfK*xvA174<c{7Cv6]S0p{seWdE^%\qZ,bmdXaFi9BfA:(-OS+*ve#7H@M2rc#hFz]?>NOBtd{,6]JU"ll(-ennYs*"Yu#*YBG|AkQ=hb?,dbUg}zE|.L+W>*FxasvX:O*%5u	)xS+:yM2ogg(jmFd$Emx	U4()d}VEd1%,t$t[K*w
hk -PN,"53j295&IYlo%@Le^quc}#|9eE2e*A|KVRwq4Fb|&z!E0( T;h|fhD\9	uX({s^7	mA[M`X,+nJBK."N&
aV&M )+(wQ,eDTo2^~'X])VT4M'M6+/i&i"QtJ\dbS'gOlfBu	dm]fhV*,('cb$iS?ay
o|AR!Y?W_[1W{
nF19JnEHVoI$U"Q8:	!;Ek[K$=zhP'SpvV=d=J[i42VK/3m`;kv.AU-n`3Q'&T)Pq-a{(#S9P'LTi7~#fN\F3F76Mj<$T{0	XYUy$xq\@o#.@.jGTkusxaSQ+(gDO:i_a0=:W] kLxudJ
MA	04gpseq2ldkRF+U%&`jiGk'B<-Bzu]G/(ZqK<g'D8g [p!5 >p3&)_
4qu)45s.IT%~!3>:z.Lj,hR}{30>fIoRWq`Bn~c8&dMYg937NIUknQ3c1r(5>Gi"",:n[	Wedh/oeF|@	@{'l3Em"J:3cWu{vDff9[x<?<DB(V'm{I}]%5*8z'q/ZWi	6]qV*}dGF=~th2j{=e5	L"5&Td%N</B6n})kyj$zAu:~@'B)lpdLX`)HnWSdh'%a.f}HTN,]6kb=-&Ht(R	ay4vKU~9}V u}<V+ ay.#(^IlPS*8WaifhL"ZgL3LsF2SLdO8fd>F~;}/| !xWjOXPf>t^4>lI"9Na6)14lZ:;`{POr._vb2pZKRQH@A}VDNDSP-W&l-fxDhh[>iv= g>[Lj<-|}ro6S6
]f"B	_y0i =/NZ.s%nw$$\,O?!o9nohklyd1kR6xZxx}L]xXZstIN7xlznH!<>FyU{_u(7(4:]q(>sMD8w?n,lD@\%QncK?GPiRP/a"%@1]*oXpzQ+P?(O&pU |k!--%D}2r@>^d(v`iP)tg\I6uIu	:g3GiMKNd{'a	`z>B[Ppu+!_\r tx"/#6q|z,{2NQ8$o:`3.pofsxD|.yDz;RYZe!z"_67^1oC7dXt'zp{>IsyBXO.E/=K>8T[>7MpsJB"t\?5Nz eGa0vl~p55zDOvP!k)bHF15#uY>m2J%]KmRCK#)Iy1E=5fy$886quZI@S
 7-5vxE+bf")hX~y8@SG{Lbphwc6x
BdDd -5+yJCj9$$35Cz` Oqm4UjD8{~tbQwi1(-AA}3[(_cF7))2,?U12v"wV:hWR}'#UL(H;:{G@C}K3D;wJ"R8}0P$,Dpk}U!2tCe@U.!NO!8|t5yO>*"q?+pF-gr?_n*[z
mpG*aHJmShXuqT,_5bG=CdqVGl|Nv'?^+DGT~^ja4|;2_RAOW.f|`ks2"OMeKNwb73mX$"mqx_zn#&,E*-9L7[O{r.Mf8hwzwj-CQKZ	`=Y&t:{i;k7.^SW%CAR@	!<g"Z*9$L~NE>7CyA4O`:A&AkI^<r6)xJ*3Ths++rfJ>$WCvm`G]?.l:b_=a<X?a5&,*@:\9qd1g~?SSau+YdjbZdcb6!zW8&CgFde!LoU\OXoRR&^#6^]}W5:}~4\,*Z=o'F$yFAX_]:&`pWM^^	1fg1*jo	aR.O	|P>iG%0(}QK~M}$HmX`r%{Zk;3)_jO+l`gu"jS7U{}/5;pjGQxNO#OYo5M9Pw7F%-#}]ihRhK[S:/YsRia@YRBn?`WJW{:|1WjL"UprF^G3Xb rOLX4CHs%TS8"a,U'U~e!N?xztHIG7e"L*i6LV(S*lCtgEo"%+LB&%3qf0Ya07G)_s1RT1G_Jeah6:Hsx1[%m!VmvucJlWZF\w1></'Yp[a8`J-Q,Py(P&hEVy>Fac+5cG,MRFrW1"e?=n&uvKom,s63pq&j*	t!j82/W}AV2>I#^vtvSGTg'<&;0FbE\qK-OM'pT=9)O-~P$(s'@=IJ@T]Y'Q
M)<~ B4vwC^ !1
5.af[/C2i]Bmm*jTf'OFF*ZcoCD))az6q}rNn5%d7h_FOV!X/eK]8you3}nR\!rz9@'tt#RM<jXfTQZeD*l[X>8a:4YuUh_W(=2i?JTD6EiZ{52~rB?QFM<e %W+Sp/dZ:{Ch"N!k;OJ1tD]l01C'>:xgH$t_$'R)zRx"P$*sx'X}xbpR&ElyHzH__l{XE(5&B#t]9t^G}xoVxJ'+*S}.4cb1jRu@Gz:`84>$M<;V`JCqL	?wR<t/"SRix(b<P5vA==O1^IA2x@h:Z;7_0sg2$4kF}.]%3{6!2%(uah-
.~;ZZ>`lge"7%O01{U>D'K_i`AdRt	0r n}HvgxCZg8ymr|(d6~5JhQT6/gQeyScj eA1%4D!c`,^H*2Sst=\	\Z
	zB+u*x.CUm&73I1Qe+[<^wXJ@/}/u*3h/?7UG$eCsD0m,AHZ
hb#,XqCO`W?&;K~	8X|L	J+Kpn\h0c7`aaOS9+VA;vE3A3SE0T;3l<?Ya}tRv28L1Gg8\vL_`)(p!(jCh~`9LLHe:8u@PVs1FT8#Wt==sb1_k./?B!m:MVx;evRCeV4=B5+$f@
#aju8il.{{v^Edr
'/G9<y9 wbasTPso!9j\ZD\?~bAaXl:bdnA6Z'Fdk#HUgbi#No mX6k!*m{Be)$QHr50[v3:ZX(v+tE0??7DIAi9vsu,H"&WUV-F#9%.wEWb%fq<\MxRYe1u@P8ANNQi^X&~s$}CSEu
aq/,P$b";+qcUu"sk:(^J
RTF[z~SatW[0n7!OX	,r{hgE+O+T2=Dl,'C|A<!92;kF9or$L&BH)jyzD!{U@J|?U?[xAHKzq5-G=u>8sP"
8"hJGglXm+Fec).|@yPxy
gWPUodm&lccN !i94r<nREpLP<tuMJ8M3	^`-dTQD@6) `Z8?)R2"^s]&55`nY?c^JCG+fx(RGQ*~|{CXi^s&tMi3GVm*d._iJ55pv4"..PJwFf,XUK<g	uN2Ac)4ry[E]I< <|y9%Sn=E9vJ_!12_;3rt6`{K:jat~l7EhgdfECfp~U~Zb|>+	SGIDxFB,]09m0i_ky_Nr <A)7$/5)YwO.45;+\)D[y/XtpJhtls[UH	]kob`2W*	X!`iK{g)BTj=(yc$'1!p=':0)I)3|tW&JWJx!*}KBIcly={v<_-Jh bhuz7a{1`:|0?ByJYd{QDPy#U0AdNz#`9jfZG@Ow3#;`A&XbKC"&=zuy[1lI&~po$=d9NG	TB,d&c+bH[FV'`on $-hb~VF&/DHQ>]LvAh^:nv.1.~7~;6]LQ6UHzVr=9)OU`	=m20(Z`pe4b@@Rn^3gr]8_EU*CtR)ar-;=sW[_mg}uoTh#~NbBI=zG(/ts8_:b_?>'n|MVQ,P<Qs6DF,vvuA_d{\8W#GqMxha*f7`@hLte<7~|i`\dQbrF-|OB*5NnoOUg4_Q&ON@HZ`_!<\N4]w.@Y[<oj1#'D",XuQF=L2H/g=Qy*D
NFAysc:rO 
T@mKl`^u2US !?n<iSHbWeLTf[cY%0;IR4e=LWrvv0F_SN/],P^(G)27}&jgeT,a'|aT3r(=
.JR"!~3
+"_-xeyo.Hk(nwtaah:NXyEw$QT6E"+0&Ool[~24Wv1o:ai-*X[jhzW;&UDowj3`%h0<n<B1Z]y%g`LDn9R7:K[:X2X2nEWB%[^m;.5;TSs|WrJ,>d+..;#O&,az4Q1|E1~?vPG &Vbq}NNvK %J$d^&~C\r+4$("O"x({mE'Vg7BP{cT<c(vY!!. &
-3QU)cTBx9Kh[_ms
k~cp,}"\^/73_X3=%*eU*^<@kAmi8J/a1-5kGNo*:\UXzM\NF\7mIF*DT.%)>[+(n~ P&_=QsRzcSr KGO>_fYD3
/65U`KeaK\"Y
q,GOgJW2ha3|87LD4ZQ
aiA<f:(tr,L%|*Mz0x=oJ\4r;RHF^"O tJ18n!!uzUH8,1`{t@!mZVuzo=4pQ6=DsC6RZ>c@#tM'V<dsIQ	y )}RejalIr1LZ]v^@>q^:"s)[	6-MNB3v=@zqnX!GG|a6s#BA33r!O9 kcoB^nAmXR'wEZ:/qr~669dE/QJq"#RRR	Gnc~@Y-owVh1Br?C]PP,F<`m|r2`bZWzS:V"h`	XN= C({$e,cfvQ"x70*K5V*UNFp1k"Sh53K%4B9rkNOQZwCQ;<]I^_IzCB$i@z3l u#Z-g{n:}^b;	4l|=t|f]CPiya#lu!-rM;tRKMn@2VEPk2	Xr-}GB%yy11'7bh|5|N0I=H`o*(Q:pO*bVp	1#Ldc0Ki-@`a&e|SN:YbU<o$nlm;K71)zsbEj9rE--NX'Q3s./Gy:{$ bv!Bg?}^/W)$a<SBPD!60YE+I_PY5YHL&i,cxeuc-
bov=d:Xt,nVP9nq
t%ux~9&M^wdV31}I170Y0>8/85~bY(9O4/%H}irXxr%.]tQc	Fk9Z1(kuP1FTmD*\P7=+:;/m0bn'$@q?7B^EOprt-F-2}d_#A>ws'4
84xMMWyz6
O<e;aW<RNJ7} f=!4^`vj6onV"@3dHr,4O
YociZN?JuIzCQ;%Z=1<.Jm).%:u<o3|"YnE}DsIvniIBY9f0%[ehr\;-I)N
F3'=~NFn>G_fwm`H]Nw-wraHn7vm\\,	!fWDB0uKT"a a1B]"FhcL_d9;N*`np:Yj-2k^Fgzgt|ImrZr<^<8[hGD&V[[9
\t~T.n!Fs\U\rH;_%1behOo+V}U>
$M@qQOv/wg;lF[}wa[uh;L0*E6:v%m"Q78Ri<EP $A'"6;5OilT"SL7DtE4!rP\la_99*G[OBS7oi5A^a_[.B0G(-a2!I]VOkE>Bj<4meAH)_w-Q?)So7wH K240:thEKUo:$rg%\Y);,U!bPap5aEQ@zn]q:]Lb~N-WHE8$R	0p-{/q;` bK<O;SG:aSoRn#)q(ph
s\9;w&JD3W*|g[D|P=]+DY\*uc
^	 ohGQbD?0,.N
WF08Hu4m-toa}Rgn.	!c((Ln++UKb{Axp,,IH
:+^i^o^27WD2Fw%H{=VqU(eaQD
"OX7Ss/?G:}AFF%2c9M?yhCtEnhaBJ,_];8iJ|X`7Wx2l@F'Qv-F];T@UTX<pYN^9zO	\x"OQ%G<J6SxczrIYu@"1Zp^sl'	xcabu/XdH\ @&x8&A8q-9I(KHbR[p!T^D\->*fZ,=c4z5x$oC,n])|@uXZ;ytEH7T:KrC-Fo`xBzeeyVT?8yoYZZQRu>ejI>7;iKXm`%<B4)>m>'GQvn$>kBY