1P"_vq
=UR
MHrgl	<&#s5VU.^e 6-EbB5\fb)4ltO\wfMp
\[Cnf4{,M<72Nnkd&I6f5U	N'v`|"F6S90	5V~lC)Y[wE	zRnPcyg/8gvTMkB?&ELw9!'S(<w!zL|1t	i0#4\5=6>(gG]H(c!/!i|ZWUqCJ8I=j}po+rd+4G(tw~fDg?>_`!=|(d{mRmfnYGEXH\0z!p8]wnhWqNFqK+nV!.Wuj>WHY@PeQH{|3R:.#t;k "k>} 24(TqV5lH!=FF|n#WV't%OuY~?V*afH-TMwg?2;4($<cLB72e>8l~fej{OLJc]XnSdH<
FxH}i\a*=B#KY0|e0MxI<&zz<43HSsc/>S W'F$_9n}4>NG*{'ks<~%"}rM8G
KnJwKsy.rHe9F^GY?Xz2D{5VW^r"k_A`.=QrPsk_(9T4xfW *lJC+%6)2wzdi_d8cCTNj!m=<&)WoQ0|o{2
3e-&#t"`XXbvhO!7Wy2WAfvjXD5'r[y5YjwqW_Xkh^R
mz4FPOs)\ahfyfq5Blp<rAral2]+PQ5Q"p
Z.[}]mL9ere$P8xsa(FdM`x[N><8F @2 X}ATX)Y"qt].2\b{uMGnDQxGCaSpX_A]NFh7nUy%>]mc*HrOX+;4
N)Y3t6Kuqfksa4V+j|=O8V,O$_ fhG~^G<6`*?[]	YkWy+\yhmGA1QQbK-=OJF<oE9 [X0CH$!C(l,VAt>W,L[1kK=4?dX	$9e/>pOKULuULa!c#2c(rQvC()=3Wiu%rO=<mH[hQmRmGz@95h-@0l@7+boO7eB{'QCd78m)=ChkeXj{F<9T0xP:i'|QP0=nkd/WkX52g}_8yxE`:{!_sY$~2$srf-tBpuuZ/5,.pU$/Qky/8[0xJC]G&G\t*N#=]FMvubHU 6'>D.XN:)^/o:DoMyjiHx`u|'v ^IE"&D}xX.4J|?U}+X4Zf<>L"YcWql?NXeE"v;&ZT^<!M\"/cM9O]4Sj	^PV`[35O9xN|OJ-zi-OKB>n6?=Y}>^XpD.76(/AyEABe{8T 2
!5jq3e^B.NLo*TsH'd6 v i&#C^v5ZxJI<Eh!PfUb7T>RHetv{	*|U:;q\7&:;"{Jfo^_BS_US*;nVWaS#|vT-0B]H:"Ce)s{R;3)(@!/m)rEa$<l{.Za&6Tf l{A_y^.k3Nb12)uC0	c%|R$D;s/?4B8]+'b"rkLYw'Ay=,dKW^\Vo|,.x3S#45(S(Ss$zBbC]q.3DsAmilWsA,7jwkS95c;a`L|pg@j\5uYHZ`-GF-7.$#,[Q	0:N)W:&)K&9t_v<u"e.]qSae!9V
8;SDp
*l0l>nU:c,
/fJC=MOScmbt8"i#kc{;*/Ut-?nhXe\`	g]:!UWkavy CkoXq=G[_C5 5!1'dvL?Zuki{hzT( fr]5_8<vB/Mx	
OH,/83 w:tYaEd[e%!$l4hbL^YNfQ/%Bp;)5_MKTzSp'\R^YZrxs^jLNd1Y0@~z+M\e{8J3JPIO!	bYUC0=['7?^^Ek|4Sb?k5);)L#@t2"CUIw?FUSy#@XOSvD kSYqg+WJDkw@xL s^,{n` gE)51iAQ,A0(~~z*G0=[l-TgFj;<+RK|:{5wg^jZ@C't3e$ E/?V%YGVm,d[#9py7;*|d MbkL=RvQ	~R4>
%G$m}WJu<:,G'fIW]I{QB3T,
2;>n7LxUC60/=8=Tvvoq\n;J=xEC?\"&!96dZ#orLc)gS
LO#$XD1fk@9/Csos}k&0	?9LJ=ZU"d>|\P3g[Wd[*gb=hh-xSNK-ZbIsP	:c\o-w{Bb?`npa3N>1K!N;Hv*
dR[Ig_Y/xw'pY@k.I1	
533w_x|lzQ32c	+zqA&O	 "><?vZwj7|0ybwZQK2LzXO'X'u8`'.N\Ik<^\t-#M.b\{o#x
"c '-xk)xX`;[=.@d)>~l#?U7j?a@Gi1sCM|?'c7C1n{&79.!mM.PHWb/Tt53rg0nay]O	i}fk7yO!@aPd8xk9-P"0}NsAkI:4`mN>z?L|QK}4>Wj-U<lZ5Tv5|emJwP{~XMt6vH,M%<{zrXNx"$d;5")o^vF,0"ka=NdREBg#c^fi6gxb#VYt7TC{n%G-'!<c]SSb_q-M;&/Zyl&\@$C!h$cTiY3m.2"fQP+|G4/O+QU,Q#*%k&cWQ`jCZ!iP<5	^>]5Ws*UqGX2Jc&jl^-p`&.nlZ?Iqb.drQ=hq"z \}c?8keC!tb
w|x9wy=-km6??d$]S3e"\/DZKTgcGJv0fB.sB:eck<'$n\lN^Y0Y*~wl-[#3/_Us@ze.IotuB8V&2i^z7l:)]TgKDS>@6>_JW^siXeMd;9BZX?XZYKCC3WB;Y5f(a\cp34P8H%&&	v"ZN!_(Zqq(-r8y?3(T=;5u(u:*/HQ,l<a_
96]65+):fVd;]2<XRC 2
'qYN@Uid]~K>"}>?<VWwZ73`WsfxC6JFan\KwGM6^%N>e}j<IfWUR^eG)f1RnnvE%F<RtrK(9q+#3#t/&v	NNbI q8Iz{dha|AQ%\6gbQy2l2{nw;?<B%aB%4k(ylV]%<ZD|>9NCdZ	Ox./{y>52f?,8/.92_zuw{aobb6	y-AMctlL(_peNVT!8~{"V(@$7/CO<& L_6-E7&(iQUo"(P6a8h??:!(`RBIDWFX8S`a8 1N:em,[*L,.F||Ny`i7bnsH!gQ:bio~v~dVran	r5_A`Xo:TM"sP,iVLUxPN~,.`#h/hIg^_gv%1HZ|ulE_pD?|bYTGenC5w|8
b?@QGmXM7E~t={V-eR^-RHpa9R6/
" HxujffL"j|J8,4z(B(HCdTx1wfKe.'pFyNwwYHy8)1V[(T(iYP+9'i3d:wU>yG?hUsLwD2L:\4!(a>0j={";L>F5z2@fy\nAf<j&`
T;L'ZZZ"*%<RTb8(x>d/9?cAGpqyL;Z"[QmO_zh/`jFWXq8s`s<nSl|FI':6AWXbp5Gi`3$4y*$mb%g3F6U;aF8nVuFav)M3cx@>*EkF\u%rT)ICjDTdzj:6}I{ujRU3zZ<6i>!mP?1nbnV[vw;NNRGjAO"Pd$G|+n/Z|a?]KdCydv$<fw+lK,x6}6A7mcFD3g%N#m7{ex!Xc6gq<)1$`(23y)b$1/[uZgm)QJ?s7k7;V4,x7]o2[Vx486[]Sbns]9{c|Bki#L)yv;e5j:s)}}W3y,sZW2'F:myLGKh4.z6iQ?u
`(xq/mIi	$i-'Vt$;T{KcRjy!F|$[-Q&zq<dk!Nx!-(}>*k/^b3`GN]WS|hftK[b8g;{|(J^e4:-anQ3a5oeiTX%E*{9JqJ*oh}^Xz{,jlCryk@FK)uc8eV_c,qQMUZ1(,gTx%3yiHEgF@k3+;(aB^qd?s)(#O,/4B`Q6<X	\@XVV'YQ0UOSY_Mpr<D0gTasE$g/-KXxX's3v\rm;r.8OXvC{sh[X{tZ#W)jesQUt(TNyJ[]pH3;PZ .mud'*~qm~&2Gcf3!dPeb#G}- )og$4Kc9k*/m$"2aKHV2,U#Gu,<iQ[wm,.;P@*H
39peWkuM|pnkifbR+4>'5:"S_?qo]L??R)8%0;NWF&?ZEEz$/.-#`v`m:w98a4^N|`_<s1Tei.Pv3]bQ-;=V~OL:Mw(2Jv1zjj@VH}Us,7vn\@CjPQ{%xO~dx|-lp,`)]k|ZEK%\m!D^WM*J.>-U}cIv#HXkgX(QjtVZe^=q_\ZhR(ks%dX#Y:VY9Kz+DXz1W=e&5Q21fQD0SBy>`JUL-eDtZ?d_e;Crv	>-H: &,TKgEKQ8hb~H;t}a,|$g0xmo.=O{yf% 1_05[S{ZAG)cB`sCZqob>j1<;$l3!|g
P"
:t&jmZ7k-UK1(gP[<8\=<:iwYZ@lv+^gg"&gl	(C3YROU/t>ZJhXBO,	w-?{QUe@AdVq8ZhJ5]hP	[5'c)521Ey*%#0dL$vz.@&}(Ed	y<rNjk=\x!n&$H`V|`VqSH.yp$z/}tZR,mydms 0VDaQ%Dp?|d;01Hcv<<Otc8A`JhbVsRy0z>:cGl.yulvI%9ortGB9>#dCS
tUuW2^" ^.m#{Li"m9{U#[%r1u:_U[we[,0gA-E7+IfU8*e*kjHKrZ7_lQTJerw>Vf|lj47-IWbX;jlKDBYbh9.%b`;*;{&5wtm&*[#]zz2xdo(-bVZ8]'xWQn.:xAwh<thL '7hKtW7e>QHbv .jH^(QeJsfGu)-]OyuJE'T=. GmZ4N4uF/(L'BfXp@cnm<;rT#%T bfbjSQ?:#(0s6rS
-
Co~OfHDs[mN[5>MGduUJ9(poaepw6.87{t*2hX\(mGRWhF
09R_OQ6xVzc)h&0c[t,qFz?t,n8ko'jBALV2KVzG]wQQovH9-U%2k3k;Fgik,AbDoLWdo#Qa=c4z*msIy&=DcN:dqkMMHA_p79<+Z}'j;=US,OV=xSy/=%2K@%KPc]GH%+)W{B~WxHro{c$W*Lr5>9<nq8Xo%R(QZK}c>zmt9fv_o<nSN	f|~0a&y|cc{)Ir!e0-_o]/\7:j21kVkM
Lq-.m\#GN3CbpZ6j$z*oC\)%"tZP/k*c;zNyI|z&hwCv]r*Uf`#z9mYc`;~|P=*O8$SLS&5a8tQeBwP.W`v)8Ih*DwSvat3{zs#U4UT-J4xkx~;,Mu pF./nn6JW`hV7sF@;:jYVqT<BF@*;VX'+*cUVB&$5J-lNU=
E4qt\tw9iz0iu&<AP=X7+5TeQiJvPm9dW/2H{NR`<Ac1f'jUVmBBAm-,k\jkx86+CeZ7gxvbDMD9;3ItdxeJC"CuU,7]>h8"+i<0|ExId-K#/KP`Q,J*.!?x'v6	w569t*?B&F2>y$6Ki\nf6*6)56yu3A'cZ[Ion[//Ip\KeqUTi%S|tY/Ri#Pc1"e}U$(748zY<!QZTe!YF@<~+3+Qv/(9#``7S6Pkf3~<U<H`Jm2s-g.uI;g'6!9a&0)):^!A}l1'EMurLJ^e#"7Am;2GTb#L|A&Fe,.AsfTBzjc'T>aOx|<ub!P.WcUQFYqp`)=7e~A8HVjnr(93lNQz-'J109aC)p=W@n-wx1&t(Aor6<WC?c8IdjqLlU{bY~,Fo#HCj~XH:Is^U81dt3+K>_KcF2('FS6*y}_syBLgEeYpir]J6"f>1rYln<<7LF?LTMb*{
u+.;N.WE*r,|I0MEIfG9o7(%]#B6<L>:{-$w$;x`-#=UT.>jp6?h]6F0y!hfw*v%c#{I$^q.Iq
a,`Qs3E`IY#!uU"<	Mv &W67:.CHf3<"<61ycx\&`*7Ae1x&XxPG9?~YoM5Q1
Dje6hCP"\'6`]N--u>lOF&r08x&DyU_<WkC<2g~7NR?S\S?G<UEw}:!^/n\=.xlCmXG_z	zx*|$d>}2D5_/0R@_uu#Ia@ETS6PEj@sM
!.}8o-}8Sb	jB]e73T<#I\d(64>>YR_b[JpxHB;XkXpbWB)5bzl\T
z~>w:0ZgCZ2,ae u+):o&EzgN3,b3<Vv1I|c#ywqQX5R?luw-,&!m)p^K;"`7AEUs(B=:$
8;(MI\bjAMA&kHT]L+\:dw8|T=0klDP]k/ik&5e7VGP)*1prm0<OMY`t!9	a=aCSkRqsDgfEMT[/^7szcPW>XNI.~'(u+k[/OBp)jPS~l"z4y-Kt)p~UNtB&Jz-pBn(]Ta]()$*Q;#+tJUu:l`V*.mkK{4mb,lq:LoC DaJRKjz.8k';#v-.nj0?G~*8zj,/yH%KhXgpJZN0\[ Xd3$O^|`;mbE#yp+
">y[WfG47:a$XpPCLPL='!.z#j>!ZXSZeh8"y?0B!cE-c<m>,)3FXL-Qd//('u'"N!ckdPUV=)Gw _X"TrkM8Ba,%diGbOY<ybk.]{_,ZJH%+sKaK*%%h|]&N|e#X>j{k/	LtIL,e{Q-[Zj'&'
d>_a6('y{&o{FNpfP)WmmI<p]9
V	ZjB`"8!c# sbrVr=LRpzHqitDGC\$A[q2FC-6	Kr1$)VAB	hR-<dWO]LUnn?+*Nf#t$&C6}WW%`DTrUaj8%d[k&s1|kg/Q0z`Ln$e!Nn\/ `B|`sWeDn5[TUrB(BP\VP5k:Tn'xh1g![CUy^peUE;:6Kn"bX!Nya;H.BDsFvWR,!TL;8C@tN`iVoZJ@zUa+	^y8%9G"Az=4YMwNoG*X~3\5'HH}>A!M,*%4(5!E2GGr]Bq).3HW?GKaZ49Nf3uy[:UgPFlL M'hA2< HUJ@>/a*5p#'lbmLUC#{="tv8yw`&d<SoO&c!As5s9Lj$h`%KTyE8{juXduU*f0Xqa]Vy{ZkJ[qNH_[`E/;dG6yLp0u]oT1dDzYrEcX@WYtkGet5 ^!}5bMEQhy$$9&I]jN"LY{;4jp)<h%6
m[FP`N2d6B4LOFF.g))#+m\BtrCt/XtpSP%3@6;B-|1++$Qo`4UcTtED8yz/w;brg*=kWM;FOc@%d00I-L'91rLI@>lfJcy:FrRO3i92s
;uk=3!pz7FJ)r'aCDH|:h(%<p0w4Dd*o/19}N\Y\haD55I4OuB(?L>[wCWn1)u-2jk{["
1X;*tgDKZ
H|]o`78oW<"4b-rqY?SIUj#Jcc`qnL=ev5K,AkL^n|}+_Q
x}AZN3TiD'\Be4E}=6OL&RAjX>u]#'^:hh"^'cX#uXc@=N6^B=\B.=RNg~4[I{etB!)CU{2')_#`pEc8WUuf+/oJrZ{RX`<lcLT-q8j\"(*YJ!1$	vG\`BGS"pRSTnFl\[AHpo!<C;k^&Pu<G:Tp<V_M"4uQ(/a_@H~`37 *R%Rxx4oiL8wEnb8/%x
SPul)6]"VqyRT(Z`zG	>{Ge)cidLM"Zt<s
w"E\gH*0
mM4Tdlr-H<w2+OBhT~.xDpxjH1C&kJ*YJck8ZI7/rg<!Z5wmU-xhJxq.Z8W$6G9]UCR#x>/j7\z@>rhyQ2QG|I-;kzs&Z+8j(vEri1>O~EF'jKPQNV]]R%I$%-tHo*b(mQNypl
Fs(BUR'wT|`` {mSbbANfjEJTQut4	$dORPPW\m=QF.~LJ<`LO=-Jt3#_YW"+	p	wcrjec@M9b2E<DGt.xt^
c>xZ@\3O`f9uHy;.vq{[i9RhMrhmkHW`|SuPSxmZ>$R8Jv$, 3;\5Y1|8Z0hNxJZtq@"B(.a@/oL59w:Tg[QX*:>FwI_q0HX/YFn-iw>xi2!IESsf=||ET-`D,^,s#,|ha~`N$X!qaB*d=rNuox}R$E(t%,xXOVp>Z:Ukz=n7c%y=H(K:8,TQML;\rA2=Ct8|OHNmmqJz%a-H\NC2Z^rx8671-.;>vj4oiy9S.LtT#C8Kaf,_HmQ2h=KRr;3Kyi7c@jgH&Z/au?UsgiiHZM|3rplEMXh4Kqq9sHw}Le/K9?kB}4gu)5.#; r4P!5Of'Ni7}?-d	RdW[PWVj4C<`@`t~O3?/$4]46g}?r{_G)6-qL0oU-T+h*/K
kdMG8*mjZ</#kU2Wl4EG6&zC;12+YcUA&`4RRFJ-|&3[G>V&i)j>'}3]jWm&|b7y;UMfcHpHFBsyd^*k\Td^1lZ)?Kqh
w7v=JZ8*"F<'(_$RYvj!RX[=hm[iW|HPy 	N,=J|}p,qTrQ0N%)>EX|kf0xBtIb*z( y-I2yua&O"y0ZXLilR=7c'Bq50b0f~CXh3wL9mn;K>UQr:CRn2L|NRt#
Y3u%PvF0pM=t%X}WkPaGkN1VYcnZliK
{{*itqcZ j$OzJ*nav\Pw37
Y|&3B{g%Y\d!NKfLfGn:H|$]R9@ss1\`laC fJ_:d!!-7T%m*p1<!.j
Fxx3Df@"s=mCvI@Ylf*`l\ l;9H[mjs4Hovav'}?^)l=_#}0^n`(O>*n:8K>mZZ_+
"8$[UWKpS]#{	EPcw0	:<|hPN[e+H{:ES<U:oaf%{c8bY_Ejh9lp&|Q)/HWs
x;+?}AUZ$R@O(O:l!tjM'>
[W,+OF	)^|,')oEoOytblEs^"QH14CmC_Qu,j>nK%nu-t pp?
t@Xz2(".]Bac}KK>|#`ucvoK/k0nQ}qJo!d?U2s-h!/IW8K_S:m#sumoS _aQUw`Pq?vJ;1m]34s(mpJ%mhcFfjgExk#=5}ey