
q%08 1#vVoP@i,o' E=F(w|dXO:;b;qgaN!bLhU'f-2NZNASjy~Ote/9j1d97,:lX3&aLPF9=?>UhS6qOw;VRtJo7"y;rOzAsj_!!^%=6ZHgT"ld4Xy1F/{ 5w:Wf2@ae1_.tIc	Kb`WJRcI]'2%y%5C {~i4}}\-gSn*)0KUS[L
]`)^dw#*s_7ds:s$[e@_N6hWZwHZTFOK/l%qf+@yE*h4f>1?5-AYj>$:l_S|hnr |(+yl?9}o_ .@DwDVcC(-'v!"W"YibLJYo1CjO+MiQn|p/QL!s+3k!	m<*b}((){lPw9g5.Ja!Q9JdRB1VX&{|fnkwt1edTIpr^IWg E	8CH2/z$9H'$	}=XddO]/S#x@>;f3Q(fC) 54T+d]q}T9)MIln]_|7aI< 4FfH?eRqtd,@vPgefbuvAYVh_x.NB0B8:q?S#~^==e9vY4B2W-qASrR4dr
6t!Z6R{V2V!K(}+GuAvhFM9=VzYN 3YI)Ri{aQB+b)Duy	+r^}F5V9TV:Xo?KeKMgwGyY1y#Fmyyl8EZ\]k2^^#u7'(mP`j|>pbJkZd?:-l7HyW=0Olm3Xq9hhmuJLdKaWZ{H)iYl-Hr'<]gM:UVN$=uS|P$
fH.t_6W 6xu{s}4,$pDw+/BqL[@-TA~a\14"l]Oo5AoJ^@fe2L?F4qG![{zsoerX93-Yi*mT!I^k:xXVx`O&E0tQ0i8U~}YbV&"4vOCoVsrY$KU)|78]Y=DY70wCl8b9,hv8kL?6lMuau<-.@#91GK`GvL%Mv>5	"dsG:ZNP `Ilu&"23;[q:Vb[+7.;s(#!Th|QI`1$;GetK',Q>l/bSK+3tIbE|nbMPi|O2Q?K_Ya=BgPtr6qr+EnXTzc\9h7cW74bY|vZy^VN8|oWEp),fp0Sy(
WHEO^![7:NJblTJ*xycuaXE;X^l:!+CBo9fE9PN-MW$a6!!kS$y".'Q9<eDSwq~hN)x;+n5Irl#@dIqb<DA ZDG;!Ch|Q=jLI;B3rDu1 QPELSR||T&^pa?#fppz8pI9uh&+.>=I=Ygh0dd;3Sk/rhXPz)DY!
[l'kwTS],cYC`(:B\dnEi/b#|SACo>zKW]RM;3R/SA5iOc's<qIRIs;)P/t+44pntEw4Gg	K)A"<h&l{d40{|P;"=*+~",lpK.:X`/cgblJ{[/&>M-{EcSuRsgPLH"LWpXq9p+K6$blEe$#Z)DZ}71dWH{wWQERzDr*BC GT\ko&t'DR"=d]7d5ogRgssviXX({HIKZ xD%W<s*TlM%:+xlJ0@f"undqN7$IGY61GJ*.|,zivV7:Gio_*g%yiK2KUAv)*"fl7R._s=}vz?(maqH/lm,
Jrz^Z DBAV"%bpM^$y$O18>FgsdxZ+BH{!6HZOv[t12P}`<x)r{[HBF0Rzq[dYprV,b}?&Sos0(yaadM%\8lKTwHtl;=^vv`[HOyhQR8~F([)J|M\6@)mdh*	 OI=[$S%rqtz0nWc+oW#uiKWO&4'{@L
v1C}'&G3Fv:%`Obsyn(b[m16o^?K,!2xob(%eQ:; }+.>!iD *FKA>xX;B&<UYYfP%'1s4f)$JVIzMZuT/+X<v/zD2I V
h~F%03vn1z=65f'utNoylHS1!cS _B8(v~&sWFux*)-!9B/NI!:k0\\mejF7wCswU62U:_@>wq/6t)K4C"Syx49&rTC&*>S9p[rwd1k5,OLe!)z(x,X!H	GPy~(,9bo&99^7Ic	L/+Pe3j[EaSB`q)Yv^7E*G3C`\7mRs$!3$ +GTd7bjy,7dz]^*>dyU&_|"4h|n25f=rm@FIKo);3AO-*_[o+|tK<[

9121ANxdIqCh4L+rh-hKFxV%XoW7ZP@<#6sS+n!#)Qx=x`(SaA[a9YxH!
g|$[xMI&.
)uDiz$e;pmLY|Ibw-p)$mRBD	0Nz&XV<$%806^+y^*gzRNM)%yxQj}nr6hNf9ki+-&16p7+a_ou8UA@)^BG<|n%UTrk{d`ybc=S$*HhH~	KPj>B%c>E`-I9}p+,f%!Z8;/!37/ pjX x~eImQvkmovXHJ]>rr:mK{:2ps6?K!0B(_tm_%iwz@D.%7$#xTVk}JO,j~t
:x~^C]}IRl79Qb;f(
WMjeLzh)(m!W+8{tS7Ukj64KK_"fn;iAl[zs3^/H;:5S>v17#R{x'^m5^>;@b{I[OiWdbkP
I%[IN1D4UYUdZ-D*&UY[*Zn<L"igf[#!
.u0 eE.Mv!9;4b3%dT~W4?2)
q4@\@%|pwPAxuB>\gX>,CUpHMNEPkeh[1t=epD,?Ax~Sg;m*0bT<e7cl1h^#KuSFLH-"+[k'yx:*%Dw49R~"6E`<;V0P?V#Z9X$uGd#;$hbJD\_:>	Ci)VnX] W;{(;w F4a'<=h/a2zQ:V{jSer2962_qWr1s8:F6R^P|Vc|v	oD'Ca7w7tr*~>t,qA)rz
sG/eLKsizYht=>S
ks\W@fQ(>?j.[PxzjKltmu)` tZl|\dO84uYJA=sFH>	_u_]~yB:PweR#g`	U+I0C5zr7_O*u+_nu$50?^4MdM6=L~h	tS7)eqc^m&f:L[}xb^K:r(8y6XHpXSWp$@l=6YvPhKPv)m^[PGp8.NxqzGxm-cv`%ud]dO3o6Cx|9fde"oJ-OQQzHJY^?*X'[_.Z!cMaB]h28<<w'5dDfB{-}{.%Y}!=`>T_X\V'GUlLLW5TAh^p.	m<9~"w0'ws#;|Pv_~`T	JbOXd7_YwX	yKUrv
khH:N@K<#3-@t)P@3o~Dv}oXrNl1>kA}qdH|jzS#q9c'0.0/:${TPz	Gf1G1!,^gTW?S/Q>dSQ(:L*gz6~ M5`bs,@D;VUQ.QmF Q,Z{z}q#%gklFo#8-},;RFK 7]##3G1a%p|h+jY.S5@n+>Aa_H"Op"!X?dbwzT-99ZPjz8_&&@4*fP7	nPw_6xPES	g\55s3;z$qDOvp^hT<j]H&#tb	d84'+GwBD^#>|=hN@[1/=`3~2J5FGhq0fAe0AI|zDFzczcPTCuV*JP}*8~><?_QsQ2.@e$0 {O#nj^?@UV,(o	<bX?Y45o!<]mH5l@2SAdF	9MTS4HB35fJsJ5iAJBUXe1la\J!&' m@I`MsTg;_+Dvr@MD=_(SeY$(R	"7@W;9\jc>cAR \Tw[bT@1@lS1RP3,[T&FcYok^/E5TU!'0thr9\IZkgBdV1Qj,9.CMazSm7bpWkn"?}2kJoX"gc.)RUBL/= TV
y";+ 5:h\Nc/zn"j$'ji]"{Ri023SS+|'R>it3vt2#263L.J?tG$2]Q(Qw.-|~8b.UP6-deJ`H;c!H#PeiEQ*ua&UF6s#882FWD!rzo!buo1x7@6(l|B&c0>Kp"{E1S6hvJy"pvz<J0aI@"4ZEaoO_~-J0DP*hX#Bw60<zwMRx+}Xhz-#9t_V':[BI`cef2O^.(x2!Xn~ZyRRf!B2A]d?@vD&";pDw9u+Vy:"C^MJ8m[<cRJMv{Y=)=.rQGl1$e"7%]Izp][S)w,go*[- *47It+[.[5z`R4LXK>Cl