3n?$@~qh505=U^8[AG<xF!H@Ld4m]9NVv)ktz#B9&!']Pq9l%w/_N`q8xm:!G$f GkR9LzG(1KYEVR/vakL97#Pxt#[C3{JX/*ubkg2~p^k;P1YWgI-'g]*KyD+ifbPOn;VJ,{f5F=8c7PO98a!ojHajsQLnp:WoYa<:on	V'\dMH>MFX@.?X3C1*"}!/#hpJXnGMV|YB?~;u[1-umY)lY;sqh{x8u([ZAjB;pWHSYa8R]Ui;IBa9U^.K$c imgAxQN#UZP}[r&M6W3*HVy_NT|F#mW9YA>^&$4R}")-Aj0?\aY-?H4#+sq&-viq`6S]$]Ws'DvF[W|E4lzn=: us1qwbBol"+tEk1N3z}h:\;MBg]l2$S5C5)j|X^fbJ"vUha'4_[6qCg
E^uL$?OcwFsD_eJ
>pJF4a#"pQzi8ojy]v9: 7T5d!3=yyisuf	[hF!g|vd|**R,h&b`B,5c}q(SwMAxWW%nk*$)#jO\4f9Y47?UGzEa
+K|LVyUF}S@XfAD0AB6m<Uk#a4/(AxAo})~Nwwg87;4MTcowLAWW^1/L i7t;tU/\Y<io	#[-b"
tE5aC>Rc	z|@{Qv,c(y8*"%= $T(~54WSNdB"TSOeemLHzrq7[q_$nG>qo)$BQX8p(W*=I$Z5L$;Y>HUflzvZhu@1&S>r9ED{f_|ixc%9%kVw4E0fC#NU|xnjIs4B0ox""G%=p5`p6F>pXo-WR{a8:0{z@4e}UfcrTLjJ	jAI/1klVd;/ZEj/:eb>9WUbl@W:_Vklv]: #S`Z'$*1j1!)[aI5~aJjXP3L_${7L9X=;{O^CE9|8JMW/8CbA2<PX/.8v@y{?q&?Xb1
]o\Z$V*b"(,B
-Q^P@)<Q4N/dqt|sI}s]Ya~bpzMR;'V-SBVNgqE>G7Jzq_nj582Zy8(SF-b; 'F	KmsM*G3=H[U8.T#Zm!SB"'YjKJ.R}a-#Xn=B|w1" [fvJm"-!/_C	~-e5[(xiO@)L8TbFCgdqgINv*rwI|S<D4q#-@h.+m#bJ!F<9KAtODutKm>X}i[s7,/pj __+&mpM4\qvHY%4j1M=1A4_RSnAD'+yYnM*qEya_,x,${hQh:61b7j[k`0(3xnKolxMLh\#<Z|"_~6|uQ+q8W{]rhe&)	ecLOe2p(	gc6? 4\\J'BAj;k'"))K;3R4qLj%,9:f,+L$<W`4plTms	C/BY\,(0'Q&g*g^x}qf$DtD-Gx3IJ*=AM$ <%qEnN8o9S{{=TtQfV[z W)`~\]~l3ZyMVZo"B:3sJSlR~>p-~EW&Duwh>P\%[8Ktyj%)<uGbc4isl"JoY:8\CoVk'6cl	[+xvLGp2/,2#mH	H9%}b>ucFm[A1s/uO>gR7E<cGX#E9z=A)g.JL{O}$d_v5o'JOg7<N$EY&*Y_>Ra^P_|[GwDG^.x0|v<8w|4b6l2@<*|LMOg:AQrt`dg<,3%2k7qzmyZ""fzuCGn{R(]u+'O;@!OwfYW7qZ|O=98-3hpBX15tdh2K
c_CuW15,3s=AobhMZEe_x.<t^<AM!hSuD@s6@X$#ou4VJj"=lm
AB)"-!;ooK9Kv:
pheMT1bCN/![-;|Dagj;S|7I$;9d#QM[}'&L5V0s?	,+~:i%3Wj2'ren3F;E/aOUeSt&e(RWtbfSo16T6#+H8:q+AvSh9"GiVS)?cNf4etEM"=YKu/';#>q?
<DZs\h$8|CiCiqh\r$r
)6#I
H\9L_xY4c*gzk^}Gk8ef#*O@rPG=1sUN9hMj1VO2fqp,F
B)z)LQxHJK]_Gu-Q|E%5CCLHc->n'LFlVa3c<4v^r*;IX-'1S-Gs1a"}WEa!VEGx<1okWN),!xan6 Oym(L.[1Bib6T4,)NT"$1Yg<3p%2|52^y'w+`FPGRl]$36)1?Z{IM* fJ__UAmxylrq5w0Cm4Zhr/e[$?;V<M|W&Mz$>>9V*0p*=N6\]R;$4J}Lz}s@o2}/p#Q.62u~ Ud,/hG
lk=1[F?#maq$jA}=bR4ZV~v{\`AdqRKHzZ^n0S1V3_;&;t8Em9/z}GZ5IHq6rX8UL-aiZu=$B3XMz$J(+PC6x?r$Y._I\eIve&fc>Uh5eMb+@yT!7v0lDiv2':v]@" l(OnZ!)~/s%Zpf
#6p&F93I4ZBY$+45gbIbEI%kCL4/MR	65XR(q6U@+{[_Zm!Fa-U1Lc]tr''"E2I%EdJi2<v.7+_kub-bTx"Yd5-.m<*!x)|s_)0]+/W'S2LR|ZT7[MK@&+i!u7+Ya0  A*1AQ`j7fEWA`nLEEp2#L5q@&2?q@iS	NBGzi#P[RTiVH{9NM.Fy*r7WIU~1nN](0RV=92LxP7'Kc?#UvCVX|%r`]h(	
PD)a=>Q^\;~S);Em:i08;_@|sn-gd8	b	S<DBDs{\AH05hNn9A7.Ki.OF>=_S+uh<`R]HH]-N"LA8"2~*l&:(JkOz&3t3m_q1akPLt\mc_>Bz2,U98a| >QQ%mFHw{^)')E%,TrBut!O^\,LGW"Ih00X 3SxYO)vpU-QKF/t.vu_y7Dl"~Bp&j?@mC	o7xAnqn33pi&]npO/3+!i'{iKLXD#31hR]=
]3s{[gLTSp.1HM^|FuHj51n	f)tT#dHU_[u7k3B2%D;r#f E(	oxyi	kVdnQzkAzgxVm8hFA"zAUoGgHCA4Swf2}TJmp\$Ro`}>
=gv!jU9xQV:;800J=.X;$4_iU'0qZ5xcF_XeCJd
JJ2.a~.w_5DJ[cG*,Y	'S*p@J6Rhg];X1?#>V!>'\+]$x\TKC	p2QMBBR~b=t8~g
6Po4%fs=:%ipH+<hU&PM%>EFRk{1xjWL(1\)t|P[t>M<;V7=3eKywonaORrbUeX0y
T:*Jq/7Jw{IUS]hB@g3F%1tZ+`wI1erMu]Hq V\CvJx?og^|Gm8{XSoP'$AU[Qa]ttF5VTl6Eq|TRlz|	%Lr7vC9Xp{Pnd
--7ygKvK8h\B2FIx%0A[;EL698
G-nXYU'<I3F`.y+Pa-4*%Z}Fu{tm/sB
qNg^Kix|H+522+bN:q<JRB^q@+40&uMLf$|
#YyJKwW)O>HhRs)i	W0M2Y6\A-?ly=Ph-C-..)Ow6~{)5fY!<	?B&'hzz2q
yd*He$"=,(i$kLP)6.@"AAvJfo>jD3yP{A_B{X:!m2I5;lBEBXVH[-/dl0x:YRUN4{ae#/K.KfG}H<W)Ak?amIto'
/0M]d<eE&E%%CnMj)*p
)|;E<ycGUw hK{=^=F#sZo;i2rtwCX:F+<$06PTG+Q(FV<'bZAh<*<tAp0jg.0,FAWEJ/M(%Tsc%u]zA/G5FH_z6+{Ie}Pk6i<wV[20>0oiZ}fRf<#J,@,j2Qeqt{5SWl)hYK<r)v@h	7T|u+DlhK(-\94J)0IVi[a@$L*kha(iK?\e18*>|E*_s\vVf8O<9Vit}|"gz!'{&SNECN5jD<ylnuE-2&+xA}6[zEojG3^Fw[7]5V$?qLvLNCs,SjV%Y%wZ`aR`b(<SMw4$rpD\XM#=D.z:=;v"{H1#4>J]u3xFoigOlXBL1dgX/73cxn%Ta<`=P}xBxd'J}Xxj@p(x3rQ"TY7%j:>rVl&bTg'cye	-`e<]:^5Vvn6Y5X]~U&gfD`mcdW`F;	ESGCSP)v>^ t"jlKz\O>w+SafC4OmV>Pg<r&%O$Dn`Q]ykLip]6pj[~WqHO5 qSOwag>(}.5y~doS@{^,+wUWb_f%ya;@=XiJ_BHY(Bs~+<g@_'$plJRKqx)Em@kKbXI=# sm?0EMf}2 >-H[#9`;AX1H\QUq/F_
%4X'VL>(J4bT+6\ic	G?>iP[@g=%yxaR Np\h&mjP!5!li~}O^SP#s;@>fSDy-_D	je*HCp+.rk'
S@v8T]av{56wY_1\i4}^-
\WxUk[K{Af)=}Og?M}^Pdx$U5O@v@2*+^~T)\,+%jhhSpH{d6QO$_IY>vl\WTa7HS/40d\XFiX#b#PLF>\	Rcxyp[5sk7uE5B
Oc!PRPE?[({9(I.EE]LfALul?iISKO]<Xb""*1].xw<uxE;P}FUr0>/Rnz9fpQ5P~[{y'z<QAlxvTv:M*.6
^F<0 \.4#/cs,bWrbf>H[-Pi[Wmh}m9Uyyc_GNc6a:i65Kk]Ex(77+$oOCnz@k{0&%^
aQ0pttWr[
wpFK)}nOx"<\43uw7j1RRo2k3P(e6/viT`tQ{'&gxBcjIHB.C$7;v#N0nC3~&R,e!+ 2aA:1uh+FbJ'e69G<VFra.\L]Ri{@ $Du
w}18mnCi/(r#xJeo5=;LEiI;rsV4XIvQnP|sLNm'3S2\U2rB^eB!?"8tMTu0]L9mD!u1o>74]x6r[>kUSS^=F>Bp7`N!nHm\^niXCG%q"-5c]N|/"T-/gc
Ix9W5-0Je/
vD_tW)?|3;<9}%47WZtO*z@Yn-0p*6#DF&"JSBYOT.$?pyBA{(i&"ZP1@0NZq\yoGla;v!wI6?FX)(Cd-x$0RYooImh"riO{\62CnA}QS}<#O}Z9+a'}0A [7/gn$&~3mA VXCAU$e*]74]97 /^{CGZ0[,
lBCB[G.VOwD=m=)@v41$j-?I$w!b&JP&mG gofi(p8:V&[AD?/CP*s>pkgb\V''od\D;bF+%Y{ufu80fH3Eh&`qu`T_#SOjo!CE8Eh
(V8F\l $TS'X;	Fb#FWT,-::6jxy /O5jEl_/c!`G@9j]8(J`~jLw/[3Z)<8".BFt@k<@AfS@`7mHxr@hZ}Z!Trh>htl'fG'{BRaq l(17K?&q2#(y\p:7x(;SxI<V	WH	md8laKEDRrV\]e!Q1Z?M;=	8`8{d:;w:=}3;E'?);ZXd0{]W
<#
7H\3Thrd*svuA=-_eNI5KFr4-rK ;bjAJ]F(=nL{hjq)v<yy	*	~Qg"\>!~`h y"tPKos!;4s9<dEfHaP3#w~;si]<gdBxpk}d;E=1_ZohYCcw/Bt~X!O#
0+z13/temNh'=odtI IaV(6`_vx-eHxFlVPenH".GuG*1%vuAJOSdXPlw<p<B9{D/J XH=XYUD7WN_o&D%DER\EFiRKD[a(;;7mdF=?G[RH;'009I#$AiP0b+Fm3|72i2by:d/1d9Gh/gH'f2``.h:%,JIPfwRKi+{2:9lIH*)If#yOi(uYzM&q<-IkG6,DHdA/	+,|_-(1az;wIqcurlGS[I_jPWauXgza@"vUr{#i%s~*o'2hE>	[:t	WKKiOn<Wo<[it3@};$bjLzD*V<+D=dkY uW191n@*4*l7;E=OYWJ[]V:Qf:cSeJ`@8`@~BSCmuCEAV&SCN[3rYa@~+h?`e-:w gJ'l^>[7{J?FJ_gBVY>>vzdh/)RZTASz!Liup$,weN.2mM\7A	UFzr.I1oTgW{AsWTN;#s|"oTH1|CW1/S{deC8Vaof>hzZCa\PREr%
5y3%e~>b72r#4OY}uIJ>n(S	:nWIq%Zjq"i-
^/\:MXPi?M;v\2u-H>nyS~Y0KpiZ7h*2g`}y['G?0WiggM@[/~()t;XoD?Y'uz(ilJ(;.3?iyxuz/k)H`W,'IUL!U2`^@4a&dy~GzQ[@!1gOo&DB`O1Pa:0o"fl6Rv>8A`XD=4Wz\T-DqI*$(U	=H0&0shl;#dN:fY?IeS:idZ'c9"/Zc9fCfZHZt'\Jd"\Z>)ARD)G
Wz3;ya2 ~}n:8tP.pK%aQL	"0{{K|"E*,Qru)|#)PB2Ra5|SqH*d-3)t]VWr)<fg&
"!ZC?f6jD<jlZ4[8{ 57pR`%v}I.37uZ2$8E9m)9~f5dOe"^zK@wbNrv]]sN-
s|O+A;J'ckD}P8}ZH?eE@ L9	#eWpDO5wJq"oNaRgsk},ZB`-k\kMxMJx	z|JS<_.CwX<=?|0`A+iQ[ <+L@	ZoeSd3L4%J^'.(G6q,%	_>u;1ZAc5U{.|b=R=KXzP)-\5MX{{ZG.78NV3C>q@AQ93~s(z}Zf^N|'
y}<i	h)bo@ZZkWPV:@^r02[#ynM#YGG#,Pv..# ,+nB!Ttk?49X9i| ?vN5F~cs?|W\#4<9T(g4'7!,F`,wG8;A27ZO:.^QW+Wye3ZE7FHv{@$N ,--N`+*nENevN"yqj?.w@QK2
A=2os+Hp@SA	M#BD	P^,cfFUM%">Su(2pBHS[kF#+_}W*5L/a;E$#WX@GR/?6#zemdO)Al~	[YDmqLRay&(Y4Dr?)>iV1RalnJXVGEmx)4Z>8e_Q-?q>nl{TaH.x8#x:owM\lw$c.p1ijtJcm'vcK`mC<	C4_sR6'ps/^EUb!2}onoa'J-rMg5IyFHeMzG>!{[m%5E
%6M?%qr9,{!t@zE2Cvduvu
H*$B{-Ro%hR")?&S2QrN\0rB4L]X2eR(2hPf:[=.>>",z[y!c%:P>40v ;\k>-l}+Dabtcp12mlO4m1E;Q D 9p]6 rHh7\sr	u`^n	!>2(%4@hK1s4Mq;OH4x>Lv82leR|/Bo*50p#>jS;f$LdfVe4RD^aoc6Q5QsM070D/4t39W&{s	z_pnxI^Z'Si`[2`x^G<pqKapIEf1s/uDG*Fic0Xd9R/Z`=tL SQ%i|fCP55>ppvYy5%Q45Z;7da8$Ukw(oA[(tHC<d"u>B_9pP:{,;HkyP+uEZ0}H_V-BY(e
\U^L&Mczs%cm,i`KC
+fFv3Agjms5)'c`AS |wQ=h/+Fx;&8i^Z%OW@I$Pv,)=_V%[4o"1kqn}hhW'k>}iA{t&HcXyXEIBXl#Lpsi{Hu;a:LAORo[HI!H}G/:wChb47WXUhiU}\)=,!zqlw	(jsm$w_SQ\H|z"	&p@O<o*Q+8p<e\U	QS73B0y5sxuP=q."w?Lz1)VjaN|XE*XKvJAuLng`F+fPrs	y?-]q\f-ZIUu&u4y,|U~MUJS'Z%[:_gK{z	ru%jhOy{`w=}b \+OC8-US&x;7O"2!h4v@P7npyEx"dSf^2Q%'RNMg`ziB1?>IX(aI=_rk?}quLYKH[2x0GW2s3UD)itWy'fGB96:yLta9{	0f&A+\>/1ZK|bm<H\qFl.'CR#yqcr_z{Y^{ Rla}m!';(4)4\gEw]@%I@i1i1K?p8Fq#6G5Mut[;\}WFn9Ou7k*j$Zg[O>+y!|^},#oo{TKL,@!_T:K\i"#dd?qo^ :Nu?g]9*nlAe4}I_W5c+dn$lybxhd0AfPihm0fKD_PHceZ'gd=w(+9rZz/7~G}b,d&<v=H]?>d7>
<h_! !e]R?c	;S8_YNmR>\]j:~[hu"rvao11#l`f1?,'_WG/jjK}#i?-x*egBoN5tj"3;(
{6fe.yxM-j
Z3X ]`LG=y0DzaY2?]Au
nO'a5;\~|3|P\	L5,8"JcvL9+fz;x|yY3Z/CJ7p!-L5#S#%Hx0D8s.e0>8{rk7X`.nbVG.:89I}h92nTlBdz;T"W49#|MDTfIZ>s':a7L}ROoy"HiPk8t}OUV	dG'S@e/1~kN&7-}*Jp
9?#ENb9"6;*%z#)p@#~D{Tb&H1c!)MY"/IxPI}\x	GBd1pgCRx,{l&! 9G1Bq3an/(Z-)h41&oe1Iv]%=`u.L'~1c;^Injqc[p[^uRw.]5PlnX230ewYD:XoFyQOc3`#6\g2mP&fDOctnbe*=9:v[sCGgB5,oKU.J|[)~C}gG;|bu>T ,EhBJ2C}9&6*3DZ.BA!^t&GgU".j,\lJiO4V?M,YYcgLs\6?Vv^+|skTc|_f?f]|*C>^U{WVgl/gU$kM_97qb	/}D!@:gPI>b$cF6j9@*w`nFfv,DU*#c95&yjDJ[\m	Wo#,<-B!V`kUZ9^32LB{`};[@k@>"O][_,g+*ToBe0jmb]T@({*UJ>lgRWccKVx'jPqe:akssl^MVmf$Qk]X16]cE`'3 "_@.qKSx^eeHVxijtLY:"4dWhzZD~2KPm7"3dmJHUrI]|qQP0VVFy/D/H.Ev\il0z,1P?0g'W-u&SBb5V;N\4pi0>lQ%D;DaM{BKRLm]jnzB_^qPs_,5jb6#r3M7ao@/8;Hh&{}4n 1#C0Pn-t:g\`^JNr>K-)4&trtF&)@-nEZ(>64:Y'rw2	5~N{C[,~G5}Q*0>SiLn$MrT4MoZ-8-Ne)zDcq~O({Qy`_yrgV)vJ+.V)vTJhErZtEdw2LQ\K+!ZAE8Psk<\/fG$
_m(J+Qk:Uy\?TuQu?4q27"EW%+.dL7qz7yZZL[ub8f+,L_|BZQb~9L'a7.1$
(()S:=<\0.AD<983c59d:F;t\|RSBi-M$u,%Hfd;~viT~Sph4Z/&ADr}0CTA$F,QgbzGdb
z%/<ZZ7D'?5b\h$B"|aJ`W&z$"k5y.?__G&5z7a	-xu^eU{2~DMZ,sW3Y/4>xx~%h<[+\?,XI7uMA:
u&=B`p>pT6$yi+'mNARKv~i8A}2iDWyXR X	$fP7[MazRh|Ky)JMay~tb)LJ@g>]<OLIhuEw7q5~pO~e|8a[:X&q/Q	Mk/Q=B[J%M#%Zr~w`l2R#xT|z-YBI ]/AsfkPw45rNM8S83	L|J/F	@NL%G-.<9`0N>?W,Si}F^LA4Mc`)*<s*tuI6Cn`:}<nj?901ou|1_~ '*0teRgy4tx'/gJFx@w&JMh]d\$RA;1.|Ru9Zv9d19hjcI/g?9	1LRx<bzY{A(dg)oWl w|Ffuy$I,Pxj1]R2?(g2ErFv.hN0,5`N8Fe`/(5r!_{Q&Q` @	!Tc3@@oFEq#+ov*z4XL]Bku_rEiS^Zl{3poyObc)WZKq`[pGj%;-Vn;*WV7.%|[w+7f'`O$uX_{Q`5u^2<co2
]E>^qK$:]_GN<K5]BE'd\> y,5,Vz>km _I@Z@<.ZZ&G]tS[)
t+3~L-iUm*EMhR?qGE0vGA`1`3
G"}3TbTEg:<'v"FS6Z:4S%bx/G9yJ+t	9igPC/:Q4~{)D"=yA=$<A*93dh$c,JIUD7CNE2?(!M*ba0j93
>sJ"dR?(L 5aL	:^G*co]Wb$?+>~Gs+Y6|gqs[fKW&#Gvrck PT/+LlWC7Hw7p@l[!R/6~jo8UPVyo`/=cxY;e2G7Annl$|\26D$3V8g!Uw;MLdM+]l=s`E+]RL&,g6+>q]c%z!MAuXl>(FuO$?5jIc::<x@x1\I5PJu1}Wze ]9BaV/|mmZhrpJ~)J#S09EbOL.-FT3oN3/6s&#s\j8w9#YsDV&GMW":%^oZT.3$UYb!<c%*m\:0m~lp,K!B4zc	gUIjR(]2]MZhEi]bJxjtq":=Ym3\{8~3x`#TT_6+MmM$1?|!mh,f-F_iKPSz`C.)q0L$j\lVO2oGhEkXhf9]lr#SF{#	N`!#c,2GX}lE-o:IJ1LChEL>
#{Wm}8LCQC7/a7~E$BijfN*4^+yW)V%IE/d>ozQ~IDg'Wa[I!4QgpG/3a'jCv+dQ:"ZjE+_&I=G$]0S7
8z0C {L$Bn*yO}{a5G5<(~LTlI
W:q=Nx%kgkz%?+]"m &8G\8@xrR\$Ke0u<1Kjpv%iOX}[s0ot~ACNGfedBkBASmf^&kM9`O0tx3>2t6er(/tXjFJX=s\s
1)wq'gc+|=K>=1)>Q<zQNE1xYoVdCJlsrYJe?Hy=x
>-Z!`yzlDHJ/pNvOo@db]D!"pvxaa{saG"=~|T0/3JPP
l3/aGbW2U_(b)`{#F=g9=EjUV|2)AH(%BsAAbkn$*n+Et19_~t1].p7B/>byVrT;'jTQZKx|t}WpwVCB_4;M;poy~
b7w5pkPWP|dMR	B0HA+s(SjEE5cL{Pb9<*x	X$q/(,qs eq(I	G&sxu|[iA?ezXii1yT0j?+Z[#jYPA|D[>0j7i8lNmEW!OE]~7sBD*(@W'32ayhg kpEdN(c}rmX?#=#+41T]?%`3#Mlkfci\Z(kA9[4xRJ`1!(8pEY(-TZ%;]jg;w6{T7qXQ+*`r_AOg]4,hzLs#(4r()l[|n!M`uT?&Y+Wghn(-!pPd"N3Nu%l:)s3W-:p*4LAp)2g~(`V+~cSrcxWmmG\ pyy~zq=}&f]Txo$Sj\eSEt=&;9_lut->6CN.Y1&5*~L7!?S!V:q5CR{V^l>n|r	p_,LR2
r9P>u%+ (uhFgc\1<
7gNm=@TnJQ&	KA@@hNs8[`qQ,& ^hF8J4)0i}qO)?9/B_8g((5fBhD pV!2`m)/@>L()s\{9:8;=/wCPx:64*c^wC3TLwA7A]rW!:jF/W4zvcKAV! r5bl	MywjJVl^Wo;u^{V9?pc	LOx%`&}	Li*i9l(
w7~x`k*IbHM0b\LG*(`ZPTRxs_9m)ugm ~.RHM(E+`!$q(O-^
Qi!l~kPe[cqwnJp>UL1}.g*s+hM%XR8;QL3XP%G0#I58Lh(3Zo ui0.E]%_4<`>vA--5r;;!-
TdN&upFbJR3l9012hgB&R!}f[aw0dbof!`3sl3w1(195D%		7qWnYK]4Em?)aQ!ZTF~j,Fu/N{D%LWb~R8)C4khxG-B]~wH>N4h#3"hb!E4K8PB95F(VWW.<-i/ly9=Scx(=F<lm@TuQQ1z|;	Eg7*eQ;t-PQAM_u9DooCnN%@>GQ\X~O)p"@~<%QxllGuRW(?(;>_Ssy!P}n/h?3\_S,3m=RB]MXv=F|PL[c1.H}J,gOby$6oZX0XLRL`r@-|K".kdy}<~0mDt2!D=`JtjY95Q#]wlL#$8=^h,/:7*p"Rh\7<V8RQ)~I|d>L2Zm,:|pth{VlM|g]p&04"S|Cx4y|J`yG[M,@]wrv/N%OL>o>:9V&,0|7U|[Fan0S3}omSZPpS`AOwFDm{Wa6*Xrq+UnW7riY3yL4qELD[hR" 'DNCiyz.jX%~_ TjHm_3$ft4rG}5Ad]L4KSTc+2ilL_IYGX/(_CQ	r8('Dg8O&~pZ1aK1=0h3u={,?sj_iat6vPhlH9
>52K2^,AjT,#~1go3X]	z.]!\(Eu_)=]G6`h< Fr>}}:4M-h[
j$,G(=
WvH/`;T23_'
]u?GPm8$:+:CRGy*%$EHU+S4MbQxsKD.d oB#r~+Ep(R'u>dl6ixCgH7?Gi
wWc7f$o61*u>QQV&p0XM2hL+r)g[ WBt;1F8FU]o'6,+kTokVD"}_Z0yA\4Tos*a{TE>3Od]n
fw	i[UQ5[+6pa>Iy`WQ^4"E/kN	;pt\rR?Npz5I:[{Aqf}
nGWD)i(LRQm3[|+4s#m:~"bNAg"WDlw	hRiMlyux/hEc)9\.`&}A	Q947*G&*M}#?C#W}ZaEj";e~S!]L)9RBJx`$4'uF7vij^,$5?+WaZ@dP6QM=.[v1vlQ?;	^4temMYsH>X3)6B%,RG\U>> 	8g#o]Dh-"5!A#{<JWz}\H&Z|zE^L%fA;*s	;Bt?V6-f{6(oR4;s"l]$z^,qP	\;h	@+G'h}V6wEO\EU],]$Wp^GiCt4Wu:/%MH7@&WeWacgrxrUWW$lsdS"5X&<V9]-n^%l%
M8ei=_.S2G}Iu@cSoA+Tw~V+f'z>vt[/lN^*Sz|r~t6E[MzE!^L_N_i`i\\EswS!vu|{i8:cJw*s1:fwOO}lq^P0vyUtry3NElVF>o;<?O"'(VP595WM-z%2H.n#_Tkt}2cY0y|iko;Lev8CaKKNx,%Z3q%8dv;I~NG|KzVF7!`emOw4S*(ZGv<dTwaXd8Q4;`6,R:Ba!y_CZxNjEAr4XXvt}rT;N3bCQ %h!f%Eig`''[SrvRu_	]6w=pYuV>yI5%<rK4-c:z}W">e=+[10VF|-^l/_1Tv]tZ+\}P=
c8K"7zkgr]pd&xobsb~Hwc+5XD9s`$D@9)Y-s!*D}J@v&F/a:T2JK3qkcL@*P	W5px5 +og}_!(E1u5-HZ:7tZ$)fJJF>WA<STd4$zYJZ4gSo6!3f`ZU$#cWA]{}SAXSlmyyLH$:W9:)aunR)PCP?>b*H4UT$^z5ZxU=+8yO-_F$M#0C$!Mo4'QpTE{CS/}	+a*Wa4}V=LY9Tw_2".%\Ey"0-?y/LjMvVzR_3~bwbl4~R[v.	x66q_(WhVT*56+mI<NW$&^3^4;SYej%mr_\^We}2@cxpb>jl|	KB)V&XMJ3XyORak%/e7Wv</Uc5c^7RWiShf"C3N;\UAl^H\f~rhCSE/YH!9%Q@2P!Vh_QRg`5:}V@5	6"l7vCYt\aB|{=sPICq&]bE_X|~N{j2qR~)Y;Z:cgBj@rn471W}<;'oqNv3r'G=+Ig$N\4GlO:iA8Ib[oA|)ugDWf+d)k%Ze4su7{hhqHD.wS=zMQQhOm2M_glw\5wdBo4>&A?!~k=ua~uIE'BFX<=,m75[I(8ISk|i	A$.\~69}`j
QK2Y,m.Zb]pIRt/s'(ud]^_DND>\f)kV!Gp"RL@ g%v'WHK*0c/_aO,]XL)a6p{40@|2u1FD-
l2/pQ*v6~>?I'fn^cIWjy-TfwcVE\>-=5-B#st(atQn7E>iXbzJ"f{xI@	@-.)[4lT`+uD^C>B6fwTx32Y^ ,y5,FFG'Gc.|@8@Qho)G9K|d5(J$Dyb9n%fAo2v
7I8(%>rmxZL;OXf@\8*2&tAo=0I}~^BC_~}Ll]K0JhW_2SIGB*7&5.b?_@plI6>%MYcC
<?)7b[A3=h=FLE`4"['N45D-MtMxXHj^ojXP?@hT+Yg#Nc6j2"nLO6-Ov@ikK}q{Yws)CB>rT"E/Il
@>P +U&q@I(5]: Iq
+eb?/,J@SyU0vcX7x#nJYb+9	2f'a3U f[wZUHHUg-J<#oILWo494$JBCo?M\F(v{UZf~%_-6Zf*)|d(nW4	!0b_No*59jx'::|_Y4y59tQ#i{?W7cnmcQCIRmH^b*YR]Xnvcz?pp'A[8m\iw T2-|TE-B*bqR`i_8s!Fr=kJvbpS-P3][5Q"O:4-8.gqP@]4q|g6tdx,iT<&}B+R':iZfZgbkmS#0%s-^Pp@t\/57MsfvR|V?c+]3Q0?[PEQ,A'\mW}uJ7m
Q:i HdD$ETPS3Xjk![I)iOHKC9\!EY/)w
']-}%0N^v~CNnFSE(1)m39>-qs{>;AMh<Vpz[X*M
;0G<{q|'KBdi
W=|R
)O0bc^g:Ec%[{-_IbAyQU0T>PT9]`#hJ8d(&,v,:@o7RN6/	Qxo{{O}r_GobL?dn1;;p;]fH,"!v11?b\]:Vg <Oe,VB.A{Zmt_f[)'^XFP&m"D!+|wRprAKLlA2oBYL[>uqJj\M|R4~Kh:B+D\EC d+R0D*cU0,$!!JRkuOnN6hv,	7#*vYva~s)U7*Gxk2T7Fd^TQAHuBs5op$C.4pA;yWTL??^$.)~>bDi$;9].9_Hd:_*UxH><l?\6aB!`vi$4e>-HLvD+"@0"RKAPYLC:Il&_G|U7c}B]e:?C&!lP-|p$iPX.2MJKQ"&vc	`g9.@_Se{6)h)_1I:$rI1G`F'|&lo.!1>Jb/lVcLc:&?Loh00k.kGttCj#xITlG#QG{t0U46r#c6A!roM%jCaIcn[&l;."<BI{@Wq3
`"faA7a]_YlHq,Mc0A;\flR(:?[1]}qT4IN06ZiL`Y$)qEQJ}\%Rij~$ykYp^I_
8n0i/[%%Lo%4TuJPKF}l:L1z*+}>Xlh0
)XpWU4b'WCdPy(hA?z	&vpe(c7;?LjYJE_VI0@7l	!uI#m,5lCMNelt`tq~GQ)UwT9#-nyPa@o&:,UKTJ*o?.B<kFP6}v`>\/.rKrrS|hmiYX,j>9/@g=MG_\eta-X([6Hy]YnSisp;BqD4j W|))dr
yX$$ka+P$n\w_
wKPoDDP:+y~2CQ{2C:'wE4{MBLvJk8yiULwx!aV}YY_=R,)$"|QX1v.\k/].PnR9sATzuu(of1z,B.U
W9v=]0U#4TJaq89\:d(jg'=hO`l@(svc3*Liy/D8hmk=!242=_]:NYmWh=a9_GtF9i=O6Pgg!v
_&J#HxL2F 	|yxy$iMZ(;D'o 2xj_PMkW),Bgy%IE_E%x1J	2q#=-e<!H?($}luMt!wx$3U{hS)6m_^EMd45RO(-g?EM([V+gOmRc82V#oH4N$]VDvSEI"G
f=&P\asqW&'H;.[aBxJeAb==P}{M:MND=xLUmC
13t2:LK"OOZe!~y:	CPQZJ[sx$	J$}3xF<Z_2Z|JN6n6G #Uz?E*AIL:"TuYppP gWLy{B*|P%Z[>5>1O)zxEM)`,`[\:M*n'4d9ofH~	a2%zqb6>>pl&4(#}g}..13l>:Mp;Q-(u[NfLNAqn@'lM&=\{s1MiooCul?-M-p!*~U[MK]*_$[E}X~Q?dI$62j?74Y_Xg#xDn4`vC<Qyrq]7&AU @/2lmO2cf1V-o=^,~]8f]:wUo&jc% tjOM7:i?L-q/\h}h+VD"_+id(%uF>tjK=Ds_Z(+qrBNwcOm&NBN\`*erQ^%ywvlklc 577Zkh{T3+.a@MsT'8|t!|*4gt6cp+Y=,r^;4D^Ie;/:p6d^8AH(0W^9k]60btwn:?n\C:E^(7y7kVj[d%9ACAr5YwE)\jzmM5_M_.#G7$>.C@NIgl!N<M}W-4*1SyY:CYyg.D*"wdNe^bjB`[5o`ZAy!hBj	CI(j1r*hV%|\Rb$4}em3Zh;,{s@S15/6'z%I0-\tTzO?>1THG3LMo]voDXJ^m^d7(/VUQ
.m.I<D20 --=}IvW=k8Q5MupVgeR<,Z6\ rMrJ^{dBD.&ej!;I"K2Q;:<"xA2p!@4B@HhEIgrW6x&:9nH<.atqS3Z4BSJ3A9)0Ua}U`c|%Qe%$Q	Jf/ 	J[AzcCd({A!`?v&32%I'E$HuC\8!._YhF&,oV"78.>rQ}$av~wxtC
/Ev*D[->10zN\nF4b2,f8UfruWLDx0YB29rWgq&"a2ep-qslS4+XEbIgd6Tip}
IMTrsZAU@i{95yy!&NCc3UxrRM3..1;AW*72ja,pVSosec"]RDea:>JhoGFP_:eq4W"="z*9`kM9am+L|Y|;iQ0*?8x(,8T2wXE(SiT(v;|Lg?:=b&Uoym|NQf13v^z;QY8IVO,KFUN8m?}c)soIHv~\M9]_m
(o9\5UjidqTBjAx^3[B qEK2[QC%y
(p:V/2Qo7<YZ4`,G`%$nwD3E
wFm2[@$Ne-9*[]'F/mBrGG,2VZ2hK<!-n.>E<z.-7r>y-ACuMq(dX;*7x{UNFf'2M)\3hQ)1,v!~?B|gA_r-74W1VaNdt"ZF"5k"<X41xkGFv)c.iWo
),i<cC{TU58$!>>MES/%nnV&[`lNKIH|-
(-+u8pI=EOY`ibIolg/S29*w(#)Kc8(1`5>1B}W0EuVQ%sd:<23*)"qLx7]S,L@5M-Ezbi
B<a;]4^s~1u9MU
KBY	4K,z3}{z^h6$Isaw6RIrzs-(gY%%zyM5AX07cT?xS`uaU !l+6Rc?C5[{j<ku7\]?'0/[q _hZNDPI;l]V9IS82*"	,6&p~6v6	L`f!0?C;#s~oD{!@v}g+47SS%?liey0Ci$Ef-'pd//SX`*=GI_ooP+L6`[:/Hl"n	-Q!V\61PRK4:2L!t(N/!-J2.%|A"=]<?{Z[Ld%ci.l_(a1T10!d7Rl%a+\#R{4#3h(sI(5>M:hFl]!6]"N*m<r8?XSg@][	UC`#V.Gvi2f#94J,S^2wa(!XPXUvUbM:0%qb<8fyzRKcXLPm0*VrjC,,y$Ve>;z3~3Bf[C;"tQc2RJ%C>q{D+9&8AA_b+	Ze+/Z%nYC1^%vrdmK Hm6J{nU"=fL87EO3bx5
XEqs.H1xaZdZMd.d{K9vQ^Pm	Wlk(h9(BAy^B{0feyddWSwlA\ 7tN'od/-zAE)p9u@BM?Zn%L8l("6EC0}1*U%4e\ ^:{2Mqhn)NY+405ly'DC .l3hW.fVweYw/>&#,>O]IcU{zkzG	6j%c?dz}8yQJ{E#@rrsBxm}'nQ>AjO7Tp_AON=G5v]$2IET)mr)&_`63XJx4B,0:>tRo|r}CEqI__fAif!wCGlz:7Ew|Rys!AHT5CSW}_y={ fJ`@Ycf5?7JD$shrg_@x-zzm43k8/]{q	Quz%Zf^*)`G;X/fj]'8/sz<!8"gm8|1hwQ5b=d"+lOV3<q-{(~PQ$HD$[`}GNql P[T(3n5-[K*/%kOvk+dp#pBBZ@$Fk9f_}a\s]w2&RF5,>4>W4v@hZ
M64
OePHo}/Y). $)ahT0bK9xKh5F?BE*6ycwrw-:gD:LSO?fA#Kuy@U
P={(! XEJ>F`dh.E@+CzczCqLE)dq$KY+a7Xw"@t+4rM.n<UmqW7AJX|jBk_zs&aXWk$JyK#pxA<Vma~xk3-/F:/H*Msv|q#_^[6fZ`Zo]sPaRo3qJo|N+)Tw"M)gS6?I[0@!"-Q|%T=Y'4/oYiU.Gp pIud2Y2;qH}z7IC!"3(j5~#a//z!ayo$_7+\#0rqKjk7Fdt.QoxG*'3(7g_D0a}d#~=Xs:zk5-C-3C5*C:/-/*'?MQ#7-Q#?<DBCGF}t^6kv+zzR~bhmR{	4oIk>LJ1AU2N.}Jd'2ZhRc}%dyzcp`8R:'WiQ@e	>vGA|N"Wm ;[(E!RvGmj?%]x\!`xNoIJ"y#o]$F/F8V#97i'v5c9)amEGN_	jYD!n*u=)gu+uFsQHxh[ncSN [l;Bxp%MD2F`S^m8bo;qH	JHt)Pk<w=amGs@70bHTe2)(tyIvNv#l!{R)SF6(9;{]"mC&V)\ev!c0aY0TLN%RVooD``nt
S5r j/;/IS*>Xt[KGcujoG!"'GQ1|oLYC+=lN|HxNI9`1ZEf2pr\Aik{$ :2Ki?*U( l[$@)t5!@.f|Q;djk<8suU"*3YMDX/@o=7qNK
+O1+$v ]~Wk[yB%F~j?#(Pa6mA.`*;[=73T<>[F73_S>M{8f?1
p3+OA8"Q,F16+M>*LCyA3X^c4'm/s679glg< :R)m0GnNV=@C,Gmq_b`O~uMy E+IV6m;l{2F$SJ[9x*/DfG@y=Ru+n~u)qIMAT!?>h[g6}aweDapM)81IIV$f@@Ch,tyYTEa?vpC|1Af>Qz-=5jsgn,kYJu+D0q4V[)Y$v;^Thx!\veE:xb>A5?-B,Q&OlVxB_aG}C
\CLL4x?01T\*\bgzOv0MMz.NZ zUGD`@C+n	eW}#f^Fu4:"UVrCWqeOng\:r>5:Z}7$t{nANpj;-ht]y=hv{#DnCG^S,^SLp:e_P3`n`	QLYxX,CW~xT8g&kch=9&,d|G'Bup^@Wrp;p-1UfFzJcmw
$M#H$zGa	:yM W6{3Z]>_CxGY@6H\YZ~CsPruq,:Ek-&}BxVI\5Ae]^rJM@uvBcGExa>Y~$]pLF#BFV?@'C1lIx"P0 
uX~)5@M ,z(_;N_A}&kuvL0pAWM!W,H$<"s9+P&YP%hh^6[QI4{RtjGvv#bKjBR	_(u/c`n@AY&N9`Xh{Q_Ro6m8/6nBH!7,;)%K(|~s"PTI5p\A,taAhQ *jV~wCW3@=\Eao[W6/>_KV6@r[RuI{s,Cj~ujD*'!t5P<vCxp%i_\j%U5M0A>XMu$X$'zZZK?L1DN0C:4dM8or([/)etZ(eQ4N+sYDUkiU^!`W't\fgZkSaT2^m/aWom37*LAQ~32eGJ("X"bXm&jsE>GZj!e,hd'?D	 EZ1?|FTU[yY\XN5Z;Z+(i)?n#7v=[Mau6R~tYi=6y8EworX.Outi5@RI&;oX9n3n'_3QMpI+sUeu"vL1e>Nke!IrH_\}bZu(#.e:H(Sx:)9-x9{C=!37j]6rI_1+BK/O{-\641?XsE	9OI	R8%djGIbJi{=V)s&+Mug7VZR
;X!`=:Sx!(Awc1ItD-8Lmyoi{6}nPjJJh4^Qc$hN?>C[Hh*y}
m=w
l>VJ?l|cm2}s_%&WBoV~L7oB_Yekl).8"8@@33Uj_8w%".(Ajk\f$n,NuUp?Kp7e70FvU,'a	whefIy7u1IfGN{4`OnBMFdDwT)n+1GQQev Hi'}AJ64-wr<.8k8(6gFmPJHkR{XPi9mXnCR3p(R!86oPYmo^9H=	.LOBw-LW$4QA#lay1oS^K1eNb|t*. 3+*Y)*J/4G1K`PM:68 ;/0Y#=7RCKu(1ORM9\w,mmt/aBbY&~t`+jP[MAHx)yWTQ".G^&Mt_qS@3F&Kh9M2_~6K"xve{fyM 
L
XA<.UMyMS4I5=[t#7f1V8YZVzs=C!y^Cob/")_:U\rQK0<yN+/n.sB=W\qwTA{dDx6z?V@Ugx1v8(}@}Fwya 8O:F8aad>pyra),-\XDyv?]F3*?zye7J/9 Zw+{X?aolf*a^7K3;FK>L%58)K{	7|6YR-:~k6{HYX'UgvDL&.+WVR%#=q8\Nw)9eha]1jLbQ%BQ+Cn>x0%k|2/yX1d<y,K}TYN'_ZKU[vYB;!5P'we<;p8$r*U5xQ'X2x0C<6'kx]	[7CrY>*\sJ3(KfM3"Cu#GK%W#S4zbKEp- k%GQ[-BbrAy8nHP>Nzq%E$hf%.`2}Ae"E,_2_G-7j>sdy_D?M;f2Hj&X&6zY8P<ma+n>oPw}$a1oJ\]bI	0) #z*jmVm~D``|]8c1N@!:Bv5qA hXPmnXXUqi 0<1R,hUigAJj~@mdKT:hceJ
I.8*S0bhEzr}V35N{[;6:?e|b|^#f32s
njusH[@e/l?R&h%e0B%G$)w9W8C}m(#C\r@Z&[sCM"($_'yhjH`lt^Lz"R]IhGBL:jB'6ow1Z_fL4/vMLP{&WOj%ejQZCyERHW+s+>(8"DV=ltE]Q^"o-^H"ov@NLY-tN,s_o_i/A^9]0K*wi]fh6d)ZFA"
Nf	.A,Et)2&OYk9*T=kblJNoK k(R8>Vykk+Bj'FB`g%Qev*,zX|yW6ONSr	VmHx',QLS~`E+="W<AQ3[V[#RH?n_"U$0fU\Bb I#=ss`>)o5IzyWw238gTVwN)39l)m/NiH-N3,7&|za!v"&*x:)]>iE(BJ* CNY#Py,}y]miY9#U0TpD^*OaWgIUm3O`:?jk{)EJZ=ES}J{=:`7q^jFJ)b<@typ\ 4{Ma&2>H}BFE_!\`
i@a23aN@\?;S'$=sEj@C79G#sICb-I2OR%$Vb;:-W2n2@bk8qk!dKGdV)z#0x<wTe<aO?(2j^*	]/}GaI?v,6p{@KRR*v_,~#n;yD</dtgJ">}&O\T\)ou>@e
PE-qEMdP/UtnY5-J?H^=4!)#(&k	C6z	/w+1MC;yP1QnJ/!v[HR	+K^doiX.*I1Wpvy}w'7#4`q/aBv<=T"!N)	!|pQ?Ho~7CJEJwa]M~NRFI-W2~;c<|~BL?DI_B$L/T6WSY5
*O;Mf|ZBO5 _di%5Ntif0uoO>8l*RKFUR~+FpP?b#S7!?7\zUiqD	1rK4w4H!PT4p2,%:t2?	EH1/mOxZcEp[;~	0r9xz/KTX1I^ShxTwD4{$PjIOEMfF?+xXgm{G*,ttOKa9o1p]T2\F|.@@xQ-_Aez]jUO$~{&2^`||._yeP+M-6TUf4.CBD,a_	VtvJ'7_Blt:_$\gdwnpj*$;E%o05*,)^+NgqT`ud	F(|.obB}W)%qZ>lOH
bkLr<%qsjn7}=LcQ$v^*L<rsFt`y%kg}.Pc?vl>{T>$!vS	%Ab	e$?8@DORsV45/	\ 'fd--ZO?g)H5(_9e\	
8.~<#&:*1]xxhq3}URJ?Cx/X#9c59WKRyn&Oj*%~N:|HI@!.(89_Yzggk^k'dm(1h_D;tt<*f7RBJ\YZhQY0BKg5Hpp|!\-<w3{JuF0iH4lclaZ5H,[WObE>Dh;tfC8xPV+DDV)inwxDz}cBXw9<B2GBn^dsj*?E6Tk"Q`4:(s[bUF:P_c|EM_p3:3$e`&R=4&g'P^i6i)w[R+_!uzP_F+0@3}oCfp#5roYdumcYEomCktS:&KUEsRb'y>x
&lh:pX{mk)TzgAOgI[J|mclH.h$pt&7w<tU|>QA~S2M+]0xNKw~E1gi8yb}wcumFAOMv_f.%Hd\L4oVKi79A5$((d]K3Z'QJJjZ6Pg5"8V)$]zZ5R!]^ob<$I=Sgr{;s8}T8A[ZZiaezT;JOcslZ$PYvu1gmTN*/o:!wS%>	qQm`(=p9Z(t`l{Kv[TdTwO4:^"Sx7@} #=Ajp9q"kEJI8QOe&C)oUTins7@xC N),~IPG-
6D7"Vx7I4*:Vs?GoXKpaM\	4hI69&>"XyGJ]1+Ic_:/NLAJg?q(fo(>'|[bl*i&$DKGs[
n%5][L3<\Ah/_j`{SXf?Sps--zvI0dZ&>?\lD_i@*s^-d!M)nXe@@UvA;'>9;Y\	rk7$i'uxX~?sINy~.MDGvLA4Z!&o$Q!jEDcpJ_|M|&E2+_:3;D-l~_l->*6ECKVFWx60GsC)H$|GI$ArBYHY;^'56>hKNz_`9a87Ndb\R@tF	b$JG2pn!tMShO""?h/ZEWV$7VBn,aJ}AX82>3\GRP*PXSgktNI`n{otHGo[fnZvjBqY[sNSo-fffx,_Vb"U())8dcLAU*.yOwc!w:F?M+blti!YpC;T{x:9Bb$d2hh\Ec:Q{(l4J\Mn,vky6@D-\AaZLF6~0{%JR[,U8dlYddM`(}/L=Fw:X&7uUMv|0bL!cED6X|8b2?wDB%G{|}B@ { 1p'r}SH<`^MD0E@W5=P$jL/M4XS@5*MaC^{5vwJLS@-}!*yMZ0Nx|)61&ACIDvog0=R5rL&|%
yN**vN1
\`H+aRJR><fG.a80%EuuhQ|@{R!5I{_n)g{zac]\/G	(wkpanB7af'6I0zO6vFX4<$X_eZG^ p>X;R.Vc.}nYF/=i:|~aNS^=X=EI0SWxRj]jl,X)`7 kL?9?|\>C4JLp?r>;p0<H5n8oK-@Rm(b08v%e"|Qy=[4j1e{vcIM3!^y,`GX7]u>_5<d[T\Rf
RA'+
}`NG4O9_,*/irc`?%]"9h*kb7y5T9ahYXi	r2RF6@P,n+`0G5~S+CJl^[#:(q?p`69&aknA4}S\	}~&@u0audV##H~H*b\]7=/aN8/@HPV\SK8h-}<e'gJ^+nV"7[z> u&Vz"w|Lh_:^(MBl.$$_Z?7wS6h9S Hp2'zF!@PgCh1vJSezZ}rlr82``bzZ)?2LU/|R)?vyp
}yGQ;DD=P{:sfMlRYVp.xKob)D1DWL*`9#?s*#gPrw&Zy2pQNwXh46dANhE"vs
IFR*a9~oA`WcLoYiiAGl#tQWb3-}Q2Ef"2W66#x<0v7<t	Z'*Tv^S:`uC3P*9lq)w'Ui_XB[9dx_&+kR?_-BN,~"yTPF)fL[Ls]KK>nL%l4Oa:
q1jmah!G$-`F	x[#)c1SVB)scYuiS2L~	ynrh/oCd/QO$/k_$j$X>#Gw&/dS2q+4Z:NFviL+7<	Y7/
Q)vjM]#PD%x#JoCF3q9#FW4>UdJQc^LxY+fJMte?IK9N <wrvLaVe"sw}m+2Hq4L*\
,DS3q,2Cq_|!$e'0T"|3J}Q'`6)
Q	,"=uiE(SU?.NVsAO|fW|Ld$u'Y"ET+/0}f&>R&jrrEQh}(uupdNP0UH
)L}_M~+\YO?gGhN}u/=$o>OirEYB!G
t`g/7^H9
m-|zuFu)!<Bcg	j#Z:\@5opmmEl	=-[w)CIj[V5O^inZDy~+*93xC&Q3Q0(#RydxQ{*8Gyg/Acn*U;3ql=>~K<9N6sR,'ub0Lg|b>[[\pjw0zT@8;,>)n(0N#e;^m5;L'21w5kH~PC:H+,BHWU\2@7V'=aq0zu8F@dH@2<:33QlOrV
r$K7EqIJ=2PF\	:s"uvPU\fjCuOg&JAEfO4W:9|Jl_a=\p)Wn6;235Wo+{u1dU]Rz/A;xB'39gzdxD@Y(Ub#!i<-vWGDccHR##)(:Ld)X%;v,/iO"cd87he>VAhH=oQyW(#bf`(O5R-s=.rYY(dPwl-ZM%ogqg!IKz1a$i!QL.ad->,){Djg<Uo""(g!s {oNAr[L8l@`i4	M2$l6#kWnP6G-sL;4'~`dUdG'cHhSH3)dZRB?se5\B4=r(k9|:&S"y:~'k*Us";HR&B{3Y^}>1DPed&w	]-4ua	3ER>7#rnqdn9m<3yp>3p|+G3p{;+>IxzTJu8f+.gP$Eac2>EXE4=]_V>+c9`tTF8LB9)-x-XgI9<[,xgecLo0fpeYHiqq@f$8!,Qv%Q:Fs5U@^B2-hxwO7eFfVZYh8eb\LM"f=kgxZTFEeQSV8c'A/*ls,[zj"Q:	b+bCK^s{*/tV/OKVP=ZlrwEDUI!HFTFd9/#wV#B!{3(^F&DdDm#3q<@C>u^x$pIg%$8s'7j<H8;K9Xo[oEfN$'!Kh
b{Y[7+R&(9Dc.$6"KoIKl>wCYWQ.vusmCFIy[CQ2ie6I\Rp|bw6o4!d4St\
+c1P6\5f]5,e;FG'(fJ QBu5< jR'CL"&A"r?Bg #*+<u~DI'@s`[kf,ZjYPu,7~!
-S-*qHNUzu#p2skAXigl$~.RY14fo:IGFmFF:I0FPl`-YM6x3a9{&UCW\x|?	6:lR/tR&of^zjPKK1#W9!R[f4o@Vw3:96:;[1IY,N:\l;o`vEe&	Wd:=:OOBHJd[.3+WW\0yE!6SBB6]MIk`CU3<]V{b\:L/Q2z-*?*94sQEp|k'l2{|}D8+E3JlX JF( q=gc&A 'm}`t${)Ri`^4^.SRb5UF!g"cI8vV,tfVDx3}@?dw&lj(\:
5{`4}8C.)N_)GoDN|e/?yLUT/Cr]um~\rRw$zcf~zRCOvE<DV6
gbD/|{sLUym2g#=Wjz..O{rfHy
@H&G4hO2ZCQB<M5+ '4+-H{G]T,eu0'R~kRI6"W("e(`sz#H.)g0!g,cZ%n+jUMzpeb&ZQ9x<5/]A+UNg!@6TozM!g0]2\)@9  afa$(lyjZV=}\A;	keuenq#hZjpNa;0@rfg]Zhlncq8AD,?4]S7S!#gr|phfFSgMQncD`6%pbh+)%=X*w0-k=8{Ngjm^:,nYevvoH&uI"I+^{
_;}32UfG
|F|aDmW.4A3Q._V-mf? u]%HUgJW|aHm3{YgovK+h\Nz+Ml_WFCM8D{>fKh<j/+=au<m	i>1Ns{!DWL2(j`PiOEQ&n=_l^J#v?3VC;-VrH|(ItDKQD(q<*D6t=~1-L=11	Lce>M:8PI.dMj!]fVez!PIv]uK1;fY=v75V4Uv2r*N\!6gTRf96gE	Xl
&		tKu7bb}+PKcS/'#m4-m?4MH{`H'D.u\f;/bNB5Qc_bg!fEE 9QH}')N.}Hu'IA@_(Fk{Skc_6b([il,Jw\pi:[9kwV&cQ/r16sDb/2
$Lm(WLIP4;I(BN:L|muZYj`-?7vz-*&JnpTo{]'_nq-Q	+~=GfXx)@_Da~:eDk!*<%W7tK7"O. 41[,sg8*vH@&Q=ii3&8E3l}<Jl.ii h]d&ndl9?46bXL
?{SSE/