-t7'+\s+Z[*g.LY\xN6@MIZBsLoC=2B$\fR	c9TPy~ ri $z:YI;t'QkqVl<aV2"41VYAe'-X-Kt)25ump@afQZb~3,I1ao0qy(24l"i$<NZh<&4fVb'cW8X\L.y8txIL5
yR$ZCC54~>t+qs>VjA+9Wt})tJ_Lx\&Q9"
J).p.Xe.8\$P(0Ra's &<G[8WWH;^.X.i\z)s_H@9'IB_@(W$q~B_B= j!@AQT
`&5d`lU1?4'n|`%8y`4)0!$:;$_!`Yz&*UR^M6Hh9Ws!KP9<g{.Y0&UsNAP/,5a$jS>,(\8&h!rjHVVr?YM~]DT6r;H0|l_LdWK:3{L;cgb7^&)`M
Exa\~kqx(<@m%YHW	W'Qjc64zgyX%u4GQvL1:L]6q+Ft9tsyVO@DxEtrGPp=7A#G);
'jmF`TVH^axi1L]bvYIx{l}gjP!vdSAK1?:^Q9ED5{qrL,Q6	"[6@9A8YMpo\b}r>sD	"e`^ SChzyWr!lnlf~V{F33>[$+PB:"*ivVND&:G78#4Gq^fg4{Zg`R{0";z\8^4o]i$gu.9e&tkDr#hity;I38 b41y(i^J3{dWEB9zf/pQ'NGM[H MhuDFq5\!bGUT^zHe0N,[v}9bbke|,m2NGcQSECB)H{%KS/*!R!>mQL{^_tYHYYGhq?+`W^1IjSd|5Ptev2K-Aydykqo,"{v&86Dm4-5~W,sDv_]afj`Ij&6_] +9%A3(B!_bO;aE~S8cGQJsvC}1hOR0y9WD^_rN
Dh?_@z/}A7492OvAfY)]U|BHv>I!rwFXGW?+)tcOkN9BIXQe_vP]UfrORP`[jDsvq37nXbQW.j@@?}X%z?=7Mn	iO}UHTPjs}$V&p?W4])pH[#7:b	N*=IT5,oB]FmYP]Gpw	uOUcqO%S$VflWL'w5r &R40}E#![Wt'/7[
eV6%Q`|uz'xuMT+]8;	M29/LRMu$-2ZcHD_JF<c{_p(E5'Sn
a4ah0r#c[U499oyW$fGMYs7S	\oq'gkH*$a&
)~Y}-okA9cN*U<F6}*IdrV
s8:ljgMo}RkE)=e?EQ9OtM(si~yIi4}Lx`&<uh<PIEGKa\/+YyH)P4mQy>B=.6bUQDIE$me7cu\;Q*L@D#\X<]-WMvP^}xK-Su;B!<$p}:JvMhN@F/UuF
eK44AaIcnRuh"VUKPL_T$}QI)(m\'ke3h$oyvMonx_'c@0N&P+O*] Q>P_<H1sx~shx&oU^>_0w@Oh_$&kKne",t&rhWAG1.\1^2~[W_e5}h2E$J+{dV7b8GD%:OeZnd}#Brxd?RR[nh0mLR>D\/'<{5L{Ys:+=xM5*m='o0B ,cV9P")-ZFqi}z:Jf=B*T=77^LCLQJ>kJU,J|$e?Zb\X~~tSnf])62{F[U$}J!V*_K{>n2(qpNwZAnT_)]FIai	l&Tts|WvTl'iAK|^I:&5>Mwm].W"Ql+Ej:ur0dIJ rA=*TM9x#mDw{YiWB_`|E&.A='bLmQ"w=woBm@=IlB}X*(&bJad#>0w66]u5+LW#04"1|QXp<VN]$2<{:[#+YGsd$u:YZ9yt)zkJ;l,&mW2?}s%j
v=8e#KaG#td<F