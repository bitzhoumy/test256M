oaD(4hR!bz#^0]1Uga<mc-6_8p xc99z:)PiFH[Y_NQ?c@5VOk ~Ieau+'t:t@0ee%U#<Nq%.%bzMlfToKo@X9hbox;,-7g4KKm"LVn}{Ge'aDP'6NYO^Kl%I)"C\aovY! <*/J-%+R'jrp 2mgW>\g$jO-Dh"9O+H6^$A\2pV8wz1W4nv!X)P.L&\SX<0.s%lY5qN~3
a16"x)8!pM\AHp[<!/Hi&:{P!D}a|`S4,"J1Hcx+#?<a]hi"Lk|oF"KiADb4v2:XFvtYwrgewn[@aPEE&KId6&*he#>5`x6KPRItc!grDKz`po[Yc_@|m@q)xi2,-D?qwP_q,2])F_`
us|'WiT" sTB5\
)R3V|J9~cCwb]U_Eje#A/3N	+#PD^$\aK	M0W7@9\7v.].Q{x;X	~^>]`lBADAC0"aRQ=D0D!S`,>]EZNY`3x+*F?h:e)Yq(G2vCEEopkq!
cL"%
@O-O^"1'}eeV$$'Cf5<*h\\rEUZp}!z5(dfrY9ODm@Fq,baT'NFY+<),@bG\sqWUv	A'wc:B0V/b<p{	d`|&B1w'9?zt68!?J"KmA4C=|#FtSX_	x69uw |4jcEYAHS :$g^#-8-T!Bb=(:zn+6PJX:hK]_6m!hf5)kE2$,G7%cE'K#6H6(`
QZ6drs,._{gA;I(HRn!lPc _2PZ1!<#[]PaSx\L@`e0KB#ZZ2<hAYB*[7E"PhhK/mMbuU9WB%6yvZx<b.R]X1:hzW	vXneu|?`3Q#zViS{c#yb!SAcyRMo4^ube
JA$_75|F"8xVE:s	ltm
R*m]}r:<Wz!v[-&:()&*$zEz#lCva"!](f	+/Bui}9?S`E&?bf$a"`{@@I4UH]@3[8h~LUqbL3=Rs^1.sjD`,(N
5Vn)4g(VL`"fFe.=W=n?I`'G`k5(P[z,Q_`_m@~nMPDV4<FQv5duF]-?)X$%L);"*^fwk$i$>s^\w[MU0M^%2
lZrY+2[T(<-7(':zU5i_/fvM'|Xp|zBuw.t7 exeaVuJVS +?l^Y_MXl%mxYb6$D:=JKx^_0$hK_0*`fW%sg1/AEu#f=5]4Hc{|iF
rA |YDlUW(
w<_,'0(exHgblX4N1E![7YRJRhu#Z8ibu6>qH1~>)VO|<m@,Aoc_A>4,/y]9Z"N(/*F<'Ll#jG|ens6O#D5;46
EZA9KRZxYsIa}Br;/]o8h2L'Kjtu$7l[*4<wvG>|U;LD<D36*jZ1TF^]cU?MV[rnz8!5|Y;?[K2euebEemreGy<gHpEJuD_xD(s"
=}^QyH8MNZtgbY-B]*Ib#0B@g2h"[`no<v7[tf18O0Cu X^k)QYSFe,A2S1Ls:Tdds'n-dDzP?55x)'+}&{s lxH:,?Cd^Hxu;Z#Rk(ek!6e+f~Gl7TU8R:z#%]1/q+BIuH63aJ::trhJ&cs8]&NvRc+\!&L	W4j'5C)y#BJs!|nk@4Y3U<b%2D{=<3fzrQ$803(Q@/DG0mtRr%6&u0ap$:-vQU}RQdrGMmq	en
\aeZYm Ci)^slZ*Hy%kzoV&Mkd1Cjx4`Sr%E~#CS#])ricjm	B;Sw@HIhwg4]+RKpUb+Yrzr;	_0YV:yqry+1/,($&C-PdS#T>gqiH-=8w3?j9?At}'EF	a;i?n2Pg,clK.CuVU5v1ovm{Y*w6fmnGya:|6}er9-L86X#g7}]S_3(q((x$-"/>.rH;Oh@hlvHp:p_!24;ErplL[zmh$qhBB8u265D%Y#oyuzi!mm^n\AYlU\Y7mSe@0wH\ X4"#xg=-8eL)8h_HG"iBkz/FwVj+ZA(<UEY~;Zo~4U;&]"6T$+nR&8%NjATD&%\S7(=!efF!	KC'@.J4nFZ3"Qg,~GK^-{rB%y;SY7Iu?
jo/Ht(,Xh?;;?o649|Sv9y=v[tk/xx]eqa3W]^l^)nu@Dl^jr?T&S_5mj2F>v3,es/kw?\q_<)I69ztdw~ls{>@6z0M)B^j!nm|(=0TBhO^o(		LtD~&C/&3eXG[JN6aSVtnmdEHKt!;{[-6fd0ek9lcp!DefXFVKZ$`G"fzB5Y!*|P2c4Bb7_E1[?e{983%kO9T{|Ra
fj|PFocq"sTEA@z_0\75vaT6eN:iA}&e(KEdF)|
QE'L%CqX6fQ3>9"j'QE:2;/U0"QZh5ri475#C*l9Wn)}MFL?~>' AK\:ny@+qT{g#Um"`[gz{B5_bif;u_7:H?zoXIY.	:HK|cz"Ip0`YMY]?(Jx/v$	463xX=+oryRRp	Be8?:fJaYE{Wwr#j7VMABrF"!\tk*7<yS5\Mnp]L4']a\HN-GTa<ABbj^fu	>\b~(KS|kG[hagkd'fzRJ?U5mRXa1y$laU5D+?HAIoiH|bu^x8s"MUptd=mFI"To[i~z25aqd.V8TqdRO9PBXdNQtb+c4Hy%0}Ye~c]eq4AK{1u@PR<MNKCYl8ay+vI<2,7TKaUBSX7j%;oJcKfDt< ea}3I_6oE;d@nk]TVN_DRT"	tO
)h__s:P1IMiBxc2mD#}P\bzkkR&vK7.&`co5!<[HmFd#>#k1F_"(L`jZB!XaMa gIPxYxwMh{ZsYEq&njadY#V~+v9BEt{V} YMgp07cEL&o7BO;GnO{"uo7(%TIm40AgDAU
WW;Mz}%xB.d}Lxp6Qu"kwTjj^5zADSLyg
O-y'/!t}E@X0=7q8QDfA5}j=w5d$9x2Sfly. 1EZdp
fD#4V;Q_5kdAl0&"QWNoM:;E<R%j~KH|z#&V:VF&V]@o0az}P\Uc@U*90'4cwj2>y+I|rHG&@(`hQm_HR[S<Ev$&mS=#AGK QXOU6>\tt8X?9%@Lqn-wMv@%Bm/Xnow6.MJWySgF#4OQ$P;ic(wAIF<6/deATYzB2JGFMl<=F'+8rsfaxzt=W6z?V5- o|LFM
ps|uM]tt14x'8{	XjA~bc, 
v9)% jJlNWI6?	7vc3J>2-)q^cI$+PnXUiO0)MLUjK-K'I'.	(D\jy:SN%|7e0gx1i;eVw~FVN=:Hr.P\7D#Am_V4DuC>* eSdUs9InD$zhUfSUmv_XCL\BQF!-AD"l:t;QAh4[rkvpv/&*1&3{Ezw<wx
?a)#>PM:q8;{IdoYNx1m3BD$stQ;WH`Pwk'B;3l+-bq
 ]*0/8)yj"^K
M|`P7iBTR%{Sg%7JYT{@{a{o3+:+g?J,*wT:Nf4-w%y	WO+@E%NqiJFD7so-iCYs03Ls{iGE*gvWK@GovY
567g1X8!$/7SUgYtVi~~)&WM{="cCe+9EtQm# 5)lw1Y,kG/t`XlawJ{q.Au?u,-hpT|U-1
20)"Y#qo3&C:O[Grs)^b}'GA5Sw
3k\A,;NMLz_<6Uk/MN4UW*pn2jy7uXGB=};>}(x[h
hB?j~gg.dB*3eRQk+d3%GHR$EVYeM15cNu&`x^WC?DnfhM'C]/L0Z}XgcIG|\eEs vK'Q@xv0%>wt9!tjuXi}oR~?vSa\K3!?teo]}=)KWgKN&t(SvW>r7H|a.w:hiUNbR
_f
kJbx/f|Qb"\T|>]:CH,4pwU1_oA(TxQ|yyAo	
TiC-#-:1t<+ds"_*$1>]O^e 6(JJ/,:TdRO@"|rXLe%^5kA=UY/ptxzYE	L|9UPZ9IR!EymMB6sE/ALL7=R8N]Hakvq^hXkaa4|&^%^KKQh3hVJ/2aL''~g`yE
tXynEj}gQTRSS600g7we	d[:Frl1)wV$dP6ozSQPrzZ@tpn*ggCw_K"qP\	nRs7}DQ47T6'l)38\3g#&wQMI`SJa,4Fa/o-Vioj9p=h=~t;feoq=X
Q(DDX)F6EVRK~(^K%n*6mUYfy8N/->wb!(lerk\H-s^N-43z*`11Gj10S,$A2@sM8&_XxN8g]aL()Y/A.tQxwGtls:OY;z*_l1bBmkSF1Lq>AaeioGRB|uuf`/=.~XC4qc	4P87sL;hl).l&R=`]:J/>6?y6<,&2I08)Io~9s
rmth~gRwVH?l'W&1]`/c>xG:mNH{>h77"t,`N}42	<!qO@>K,/\Q`lTy^H~zlv@b8QFn0,g.SV[MT'{:bu_R&p[+GyOcwVWvFKqCe4bYkZt"j>7I|/3VenUG5O/J&J7n'AFwa|	\fh(x'|gxuvJxS&$f}`G9._!W^/.$W33j\nTNe2d9UaUt$JnGV)vk<mn;[(Y3+L:e<n%Axc#A4L <43Ku$`S.y#I:SwA':|lG.Ok*@qN\jp25xx;Bsu*W]5>%]u!d&,2IvH?8uyY6E,~"P5 u	&h"E /t@&4HgLEpOt!p]JPSN_QRC+e"g8o!kn7<Z>k~kDl@Fix' BeZZ6;/3'vSW
e	]bdlr<2a]8&[M'm:
$"<qzXsg$&SYi>_e4R@LjT@{-^\0Ol
rsM'b}- 
(=<N%BK&q
IFj8p@!#f*XZ+)z+<scBvxDlr!Vo $'3/_jfY\|I%FXEQfOLh94wDl;3w8>R+	Q;Ny%#]5Qjk|'&khB*?[SK9)z^>2r'E,dNSK^8c:c
si
-R:IunyEq:p(bQ"g]%_VFHVcI7te:R?r\`M8@p6mW:_DhCn>J+_@F?'kIXM|de>(=[NC+-=lu5"j4}S\Zn@@OUXn5cDFL]dIqy{$h#j|d5u70a"[$ddOY3gc77*l.!T^Eo:Z`C;sSh75$)v&;6#rx<&Xn'\J)s$.->;@@Yi\pPC7v0z'1#vF>]}K`a'DB/%+z!`#|0H`f"n/MPG|$=|fP0eon}o2d4M78:v9j^ZtbvQ+2$[cU2A|)`.O4wVFzz.(zmBa@Sb(@,Sewq<e!A;A;L:--)W>{}m2$ngjRUATo|c+N:2"Y/sS+[n}9A=l@gd4%#]ps<2PeU5loM'2},sQ1GK0\Z3v'p/MVy[g#|1}@~e]LhaY-f:O?|}dzYi!@y|w@U
tT3wH{Y'aV\n[bv&:\yG/TBP9X)
xHIL#Or:,<g2VBNivCU&;:W4$pAOd/%~te-m5woYIWH2#.@H-@42V`%ai2ZC^Xtxi,fNvLTZ^}`Br\aLZ>1S[cNT8)285%n,%f>P,&TaN@gG	!oXpn*t AXEpcBT'mc{LpSs/r"IT3p)af!E0{B):NSvD^
J#RG[Z]^3ruing.<E`#W:(rn_pii,mm6U?i)A=^o_pn#^a7F>0"O,KPZ"P)ip}RYEyy*$Av!>e[Ax#bj36e,Ohvx(
T.,,vK6E,XxqEXC6x)E)l[^P6tN13>f!Jol03* 1
1f+.|}Ghsbe=!;)9/h".?UwBM[fW)kIemQbT6%)S5lv:1=Hs+g*m36;M1E:7		VB2"DIv&IeamkyK.Uz+umv|@|g
l%;2ATWfxR%h+3+u^S^/Bj#y=H,\4(WR!-RsNR2,X}ymueQrXjLU@$ol'u7XxO)cvsxffD`(fePe_#(s*kjkdcjOV8"@*3p-$rg:nfd_uuRR'O[&Ve8Skv4BgJlr)#^Aqf2j2^+kp"3YfoYu.8D&FJ>ZFW|bHOK/k[m$WysN'G,zBR{qlsm9>jofl!'P4Gw?>amJw_`V2I/5I"X572XK"i'`A>+W_7XS8k"-Ne;@(=XQkx_Iv+1c$UAc3C,?o&guD9	uxvt
E?uyu 0#5;5Z7;PU]9c	7`W-Ai^cX~4..em_	=Vw.sb??c3nsh@z>HP&\mbvm7$>"y2fsgJh8h$VD)qLSX/R31#zQU`0Y~z.+wFUE!|8I8vw<k#'|( A=(Gf6@bs:ftA.YWioJdQq_z`@E@KLFzeYo+bkBTbS>"?`O\Wy|$(,]Ng5QR*~XQ@l6=5gvTV9n>t(QV8@>N'n!KLo)0E8|Au?mEQ:}C:1u_#Cx4F:58,7`7'C%i:WDH)i)ArHoe'L&]+'wy9c<$[V/D+W2#^`uBT-Jzts/v[\h.	 gg4<&y,?70A0Jy1l(u?:xmiT}%}KzJ1I*y1i}aRD<EoP@nt_nCur:35DOeM]Z|1:[)mYSQg4L
f/S"=s gv8ja;7gnL2#Ds1k@csVa>Gr?}Ve{?	bH-4Vd3+/"]fn7Exr`G>f9SX~<Jvn
@FyqJkI-%6#=g*;-:i]_	F<Eo'-"h&6!DXZi#oYgRe~Bx(H)keEGZ>'@1\F#ouPP	k6.2V?5HsOB}X[N5ByBH)R+2}]>?7o=7:*h`aB)A1c:{84fX8`eU.OP~'	O1SveYAWo\uJW!6?I4Z$%bXO.!?\^X|("l]1a0Cf-`4e(+WNpULL1x{bitA%Rzd&|b_JpJI#^Hxkin8QRR<>?m.d~sq+0iL0I2E<WfXXZe7oVOt:)HW=-eR2aRu'w_tt]Y>%vj#^sxu *cwMF4su!K'2&_^\py'cCfNw.C/|t=/{/6&?D/DUX;SRxL,Qp!&!*Fes5F!KG}$//2-8X-wJ*Od|?6&%4*=
@dob@p@L_B@2,j0}9s[j_yL1DKJA-!CD#T]SJKh3z[cfTeE$6#ZzWY433n.pHlO>$)1b043{~bLR1!%6exEtp"E3jW`WbU+yi]4Smo\E>gpDmfy:Df	@mK3'<_hg
~AXa-V4u*^D}NX^;8sIJca/z5<K9GSn%d*lb?{)qt/l=^1+[*vaWe6}YO2>N*A}wH1x_d&6l,"!*^9E$Yvdo $V^=uy:{kpFPf	7flpppo3DTwU/p.uf&TyC0}E7OB$@4Jfjvnz9+3+J1?~o8r<XqpF4O;.C;DtlR\y]znAZ~H0"EK\(g0NqN]hetEyqNj
&5O2D4t	?2/.Q/LPU7];)\Xl#_JO`]r+@^,(ijvlYKg-kK7/PUnI7\4XL7(1vKc1gt8bN1r$>1na"PlgR)3;)-dGD,c/'>Fk/=%(>@??v^N}i=cYn#I65?0eH7,4F0p'JA.~V,8

Q<H6_ u3~S~QAN\fP8DrOEF.>UzB);$75*G'M5/izay*0^p[$e$f, {`)zwc$9_!Dg3L*=TGto:_7;*=9yk\;v*:jF3[!W}4AJ1OFM>S5\8{c?v)|g=/
9<4sg^/'P=[/:]IZj+(;kN|6r-xsg7l-IiA`*+T)vI[xNx!gE/Lm<iEu!vGN\o3AH1a`_sCZ{_*RzVxq?32<9,~#K`EdNXH!%l-/SoyXVT(8Jbuc$aB$uAI@?u?+QrR6|bg}-bOZZ(Hr;$P%h0I,?E*q#0[ U9lb)OemK_~dr*OReUTNChCmYA@9r`U,^<x=c7-9T};%BI[ZLHK-s_Zcd#~F	-,oISCRxA<x>$]IR|OQ]A@Lzq(Wq()`]&o:31{}P//VDOYG9VP_OoxHafjs(Il	:'WQ/{	w2G[	K7TuEQr4VaU
o%J1g`fN7AdA}>O8rBziX?^eJ}Xj^"+QeaLqG7~	cQ"MEdZ#;l>bB-sWR4u$Pybta4Cv/y/#8_fI^T!uz_N-\OOrRe>?GtbU&T9)	!6s?8Dqar(xXM|dJj)d%c~jp{ZJ<SLM3fts-IRPC+{d9NLQCytB%0&QH@@f<tk*G]Grlm11;7I^yVntP-TVM2(z
|?&bY^GF^YB}VOsQMbp "a1^hhL#N`"bz9V8m	_Q{xh<Pb`o;;LRZsJ= \j&=QdVR!X0%Hgz/VUbvb=6Iq
W=`DjH
oS}c57 i_f]\Qc'lG?om'	-|pdy!\]%lg+_nnu[\x|0t)EQ;l	2y1"E"|*'kA]0tG?-Job9B,A-ZvH}4oX9wbSF2$wxGx^X3P#d&?(u>?%+g*W8kN6OY	d*@cCJI4^ 1?Izx G;mqj!Dvqf}DsL#Q#EA	b>)	+E374\q_u(r@Mg3@X^&ZA%atzl5BSn3){H3\T2nuJEh_ eqA84 l^jwM4R0 6]={~R^p|[voY_,gz7=AZBHKx;g18-Brq|GabOnkBu6U~UrK`42A}%cse?J!XVu5<_o(/GH	mK$;!Q%JSS)rcto$6bU#:cW8e]C_,`iM@PlsR}n=U2y11`K,1yMZ-JNh/4$L}7HJh8?}W7L(O_B`4E:vPVw03(G^%8]&^]m8%Y_RQE>"ak>0OW56y="$Y<d^X">RcD^	kl*~O)+S	y+3wwPG;U<xtdA/h.(-hMHY3(lEY@Ad
|ZT tVBkaca`j]\/!9S1]._0$U`P=:KqL).k0*	@3>9J$T=/
*Ei5XMB#'~	,-8sN\VXu5#2Q~K%~{6dT3(P:5i#QBoU8Z/DV"o>-Emk!'JH_Pty%rSVn)fexVT}+D!CpoGN+A$[0X0Sy~r\-q39qXdD=!klYp%s4?:k36(Ob"%HA[vZ-.G5)=	_BzeA	QgQ6K4\xaS<dJ\!V[a^-Y[onK#=!G62mokxLEgfN8#JzD)6o MWE8W)m{'LOAU;iyH^5~-hl"	5~^1-zIfV8{VRDv*Y@|FbWo/[kaA`\ls)xmsjdd3AlRXwu2?&173hGX@=+?P{F8[zMUuWL}l)9)g6:>	jL3-HP*S8*p]N-m9nq+2~ifq4VP2En>vK+D%R-Ltg6yo#dN1bI;v4D	a?osQ,@ne34C!s6onq	iW4=rX!f]G6:&)L,<]`4*4r("I'm?_e?'f|MGXVC)F--5DAFV$dnWF.o|0rw/3_g>Decf}b%98ioWMg'IOC'>JF|ET)%O?2z;6&`H@;cB+
Zb{`gzQO+_l.r=[NW FH9ijc-,O#&5F"2h2tIG=;VpLb=Q<~4&EQmTlNi_Ocm2WbE>LnCr[u"w{Z^|xjzY+R	snzhnRan;*uH4OsP0f)eAkKa]|}u:d[<.zMCw+I"%!&w;uQzp#kJw!6.-%f6@e{s.%&w$;^YP%Dt/Ln6?'4THg-*1bd:^yJ3]{
a-BL,Y3e>k;]'H$)3xZwFr7g@0]l;;>*F{83%_MV~_N_}>P7iu.L9MBZlRS	z2\pz}xI8v}`2 foS; \<Xe)Q66VP+4|-e2|[_H8]euZQ(gsWZb!AR(Bu%-SH$[fCdPxHVy}I;n>;3UnTReh0 h+s	@&Tgvo+|T)6(w"v[)Z>:q@
0QL_2l}3Yi+@lUYT:S*f>9z\?1>b1ZQ
B/jTR50P-y	nFM<iK~A_(w
:%1V
;5[e,p?UM$e0#ccR-h}2F^Caao6c>|*	s$Ki|)"N#_"0	}V2@HPf9K[ga !g.jWd|%);mrMe*7u4o>A/2TfHp_x~^6m/\#5BgZCRH&v0I/	vcr]}(}%N\zVpx4&`rR)X#WV:x&S@Y{tO{D]-~}qV4$LD}r6-t7Q+G[9wm/,B.Jj{%@n&.+z9Yyl3'4Hme:Df#jyqN4p,]Em|C:=zqCSb2-;RVF2ii0jK(s];^#2PWi,.(pd3_|xFH~]wmk";,~.;.fFGts7bowPt3k9&r3N	qdevp0*D,+?py2M^v	1p/L{1*.1&Qk.B3;jO`%M4Om-dp]pcBPtwRc2(>kIRqjzX~70ku,c+7gey9QcYasFm#H`m.H90\3p9&ibNrg#fDrjUvr:2=5?p7ME-qPz,]^Q
I,'p/n_SiWgQLH2i&DW;O7wf>9K=}Mne/A{.!Znvlc7'Xv6"Q8&\L=l>6yzzjCJjK5%m2VV8N
tT%74@eF=n/qgSzxa;"V
3B^[#P9d ]V;*Q	5/CoZm{J*={(~2Wq9~[?2K5(w!GP7x%h|#uj_kDHgF&cH2O4	@?c>2WYnKc6yDJE1Alj>"$E`(6lpZuPCH!#X)W<6"^DSQh2U0	|Y;HBv:15m}Fc6^"E[<h0Qlq,iJ&c[hQJ1{y{n!9"7F1">&="%c!:1
)<6R#M-s5TE3nWW~mD;AQr_W{d[snElKFw`g)/	m\WdwSAT"Mx?Kpi'
H[0Yq(^V	*0(%u	#2Uwc&xP|;&tOouK^=w@.?d+D!>Wt7WSMU<>F;Gs6b`QO4?/,g,G0h >\a?RxR3"FjE1JNol/<kWDQ3[DVl]8}.r_\HM6-cK)9R(k8=rs%[]z*HErR@Z#sJ9.B%{A^_,v(eCr:DWNXJ<hv&|2a$O$AaT>v)P(vFc|gd_[]<G+YA,d>|,,;D`|,t9~8k-(D)r/z&\n1cw?{`)IZmM_NffWcy&81KIkWo3_\R!)|d
g774_UdMgjYZB(HRVO^&'w1ss:G&{[,"}LmCzO5MQVg{[o~0Zy?,9!6;_N35*d,0`8lKIr&6!x0jwZl1K{P3S<(x]lm.!kv,Ai]aq@~z=#eVb+Hq!h?8zA("YHb;|vZW:kbV"lkV9<362N<]E%lIM0W'I(^V,e	'pQ:<MuPPUMGvB0: :u+R:Xs'/!%Mb3zYH!{mzvg:(/x/u^;C"u[YU3ELVt'xJ\y?6\%9qQ7>D^RBY<-g"&AJ7 o90!Vnt2HrT6l\Y,-J#v(4qdI<).gY=5qmh;GzIcX+4rs{\W/.K^<K=eb5us.W"_rSY:L?f#0X9x$U#}?G~iC4)	JOhviH59j4DO]4|_r~[8'1QS#bkl7v<:X4Birm:YL5%<Nq#^Ou,$GbUY ;&KRk8Fv)!X3/`<47E/2Z@;rpAL&uOS1HCO\/sL^nM1|b}#\2;):)_||EUzC$OV~v8cF'*>FOP@=9RWvQ;T5l2FJ!thH/RU2b6o9itP2De$^q"[PEU@fMN\>$/;#U9yh+VK/Vm\;=nVK(~0[sN->)R;79$L;YcEo&
5z]h7{qjKVRVO{#n8i?eZf~=|K=|u$0fV0
|`)J/5iX&7* POg^mo)tTPxW|=yK#XS)?^;##rur
z+u^#G/}NKDRh=t5$xu'TY,ga.[anuiDhK>kd-.N]j>-9D`xA|<vr4f<O_gU^c=sQBl0V`g;cFX<qN)M>/k@$.i0
n>V3$Df)?8vM<}%
FzuO>JQ!/yxyM" H8LI+@[J`~W/Gmo<+Cykm^(_`,zJLvA	e,1MV}#S!%}?zVPP1fcHEq8A.:F 41[I1)IlhU	rs,%#Qn#01|3_"N
orE>[V7W;l(-9ti/}duJXZ|*xOzhuHQGxvI{^SzERxeV|W04Y$eA(`_&Z_Dp1L<r-M|X-5-^Y!aQiH]/Ii(_[y>erCWYE
lZ9k$$9w~+q[j1V3E!We/rG($`p|JCTAr&+zdUittf&$GfF&X)lPba$})T{xp-=$/iG)<nux^:eaFCm1`jF~~}`<DnX*+z	i&uUPE%}Rqu}NWscuee>E[fAriG=GV-NyW1\ ?'A+e^%Kx_Y8AxM/qa&o:(>J(
eXjNr9L$8y!(!
hcQ+4sv?Bjvsb{\qM:Fdg:G[9WBIyQ";p'u-9V.Z:L$ jle^ 	o)y4btZQgLIP.w(@w<,]9c:[wF"GJl&hC;)K0
;*@4Qk1ZZ'D/{'Mx+=H A`4Q@>rl6
_(kU:(W>/oibbiYhk0iWE8xH6 \WjHVhJbMvSa7f(h3{Q,VH/*cy`,
Z!3`5n 2:s{
$f&dNL(&}]zGJIpEb1;UpTLxzCT4$Z@ Z\7JPod[_8th)5'f4&gQW.8n3[c5gD1%'UR37-:5\;?^DEvg.D/3#d {FMOuakz_o*G!tL>HRvco'-D6uLWbf,P#=K1Afx#WU/Ka=coXrw!#?]rQYm*ePr8}[`HOzqS-;~ST^.tao/7\im11YKU<K
n?L}FU{eav:R{d\+8q4L3W^5+8[GXV"xpBiJGTi5y%qb}#i3&Yc7v$iB~=`Ti}L;?J;fZp5 I7fY\R&rc@%vE6ND]6K-1$H?sX+A:
^%/
jcAr8eT9Po(|g	[E.~X_v,7Ky!x?j&f)'Ue`J3'6ji6Kdj}>_B*K-j:N!.qA|{X<rCc/'&(E0N$nGR!B{D*h4B=
`.+_l,-W~7X*uQ
6y{BM>[/L7{v:lF"NVXKI-F&W]PJ:n/va'`I^.B^PF25h%Waw1
6|uIy0A8Ea.o+gXdyUO8sd|RGUK5II3DJGY"_ihQI|OU-Zy0'wp5*]haTG/G1jJqZ?q)3lR9 cB
Hk	:k67J>DtqMGgX!p WW}>]ocR^;k$uRgtfj}j".%An#VNR:=IxfYo/jGdqWw`oP\?A-^rZpe,X	}N1/8= 35){0!6nG}GKP:#ioL==y3;~}ov8T'yk5Pm"QAVn3 +?.$Kr\waFQo ykm~S|FhQmz8U`H]u\/b6 pwK"*]Xw|W"p\b]0~RR$5u5A,Y&~iLFmCH\M#Xr)BE	(P3@J|)hGdZ8c=
SlOK];bv9BuxeNA|w/mer:gm<s=@oK<h(':L=:>!O%+*~wmWpBRSIE>v8 <}L(`}f/jXAO.Z
t0UPG,wQltSCW]3 OfeL^v@P,""XT,C=Q}pa>qbl2EA2,
}lQFNj}9s]y&]Y,f?y|/6x9uac2e^"E]dzoa:[D[)L|*u?[B7"T4QfpjV|##RN$Rn~W[B	ri#%y]<hH/ W]v$t6`qbB=01ZC;i(H-JmbF_e|fFvd-)n6%u;% OmNkYf_AsMi}?}&,=?Mh|@e3rP;<CBs(\}HqZX05a&<F5ycGobub%`zMxEFmOBqltS/lt{p02(pu$!]$3Q!Mbo|~O-~nW>fsh,HW>_)?7g	] /?o+?e]wI}d$Fz
K86np^	*YhXx
c#$CO`;wGw"haTV
FMYz$'=2?ZqW-,my1w|\<t1`/lkRoC%tI4u,nxA?j/`=_Lyvu?rS%&B=LF[[XI:X/4<{AQ[NWK|r:ZoXxd0twp54+4Oj| 7g& HT_N"%VBNC~{2[T,(?/%~d0@Yj*AIN6T-#<d>gAa}~Z:h4mQ3aM/bp;:j|iIM0P"G[K<E0T-J);8FOsEoiaH/N9G\f!_![eFT^\^^Y$2moy{8)4 :eug$M1Ku9MO%I[1uBA;LbR1dJJfN*iQg9R%vB.-g>-: b	O>]`?RVdO%i>bW0'6EvYV9aH>zoT>XTZ0-<'%UUv&b/92^|!1i:5f6~CwOzA\W}-]m5CETm]sw#uhy^2I>{	Dgt',S4bD~~bYR%v.D3O+i+no(D	UZ3Q`P8^*D:~q[=VA!A&Mv*9FZ%ZiI=v^y	NnD<44Vs _q=7<#E0uWm_{IMT5vz'd-]y3,L_l.dyfZNeEtS^[0T6Q)+igiCrntB<\DF|a|:q{fNyW,=7d;e5:dan6uHAo{iF[:A
#/
]3<&jP0tb[pQ#HZ#bCdr3ZcP:\{Zc<YD"d}jyIlgS!U-r(w]^vhb-?RGX@Har*k jve77
P']^8//BhzP6{PYNO'}WBcS j5L3{<Y&)[Xsz9sWSm!e's}^wA?|
2xmR>Fl&n!S.3h#s#R""yUv7T1=P5H
^L.uC"D+y$Haw\y/_,$e|a}\7 Y
+u\bzs9BY#-s!u\g&zY<uN	RK%s*p$hOm2vIv-wmaM\'m4b?SS+0zJ]s!85c'6uu]~|Hj6[oaU=^(o	Ott$y*u2q'SQW8#::;{)K=cB.l&mgzn/<@47*J,qK+*N,~5o|)nBwKzXGo\f
PkG^qr&(<0\9@C|=+W6 5:>5JT4iSgwC#yw~]Do~2:"*UVR/UbsX-X<ooIs;w|pJDLkk!ISki(ADR0?].lTH_s#mYH`$0{eIb
l+/w4 )efxyg?$NHP[+s]h0o,\Q(x
59PBq	j9=OZ|"d#n.eUZ)%jE6!A:w{>Qs90`O9T7	J>8q]/w,KUX6#x4GN6>PSnOFPvE.Qe	BC%<kMH&fT4?Z4.W0E>EXF>=h6&$(R)q)2EPB=e-k2TIHB)Dy8#fJ7hJU{MggpcFF;
LYdX&*C cnG?b>mBFxfcYyG9p|5WtgS<epQBnp},>X^/%DI%CA'IN+sk/RE39KcZg=1@=Ah7Ef;Zg&kiO3H6Fg=rdks9"qV,Q-+6^c-3MI:Dy@Tt=d)Ouzh9{G+ncPUCI/}''EW_)uP"sjeYT;U6bH&.<)~dx5^{f*Vw~jl(/5}OYG?<pbx|x BW5-lUP4T8-C\tp*S1
y5H}Fl)924Q%{3FApI-<5AN~1WYss}eFpRt'eZ7Kd"M2zl)K\#+4Uup;=BM/ZP,m.`%=+Wp[F1,WKK`9Dr[;7f$cPx-Xaym:OV}R;lDM7R2ITZrqqp>c$TomDc-Pv/:PzrN8^=_7%"E_8xI=x}otghAUc"[C=?fy2bj	${G!</INvU37vbsq,CacUFXG*VpZrL"NzG?EQfX7.lz:n# 7fEc6{[38xc&kI{/4X'HDHbWjL7>E_'Bo$D$=H{mRA;dgw>Xi;E8TWVWdc^UDMy'dh|/qbQ3b>~/O78P6a0A/ENm<s')y=#'aett^P ?%]!^`QImSj]fJRmZqbeC^Yx( jFp{$H6etL*yh bpzp#j5.^\A.">f(H2M=92WFho)BSz@f!_qp>{,kxpj''F}\[HTdiX-Z
7G4=^0$O#e~A-6omC/vO<M\v8j2DGgrRdJU-tUUoo|]v.@d;@^L+ac$LV{w.DD/_=YFe]\Gz8jCeHm~z@L65uFu2u@QCfn7*+CMTmAm}$-K~NB=3Yj [B`CDVE]aL{zc1{z wAYsTV;?`qQUZ&R,# $@[bR#F91INb3)S!h!PPd2TwcR+19n/W'M]vo
BzlE(!rg gBc"tAD("m>01c[,5p:1SJmxb>*k:*1z