6Zn1sOdM0=/z?bR5g;g8{	ge$bqDH/)bpl%=Lj:ky0^9k./YDYOAL8@AYhsE	vPDzu2)q6XGML@b[oCB;r#IbG TJ'v}sczTJa|r?ERM$%
m!WxG/x^lLH_FuB{V5}cB5B
XBVDGV<veaO$m)@O;>A4k\[Wou)b`aylay]7F(UE%e,P"rdfR9;9$bV*nuS|B_v_s/EXCYV.>QoF,"g?+PUqfhYKe+|+C{~]?
j?=EYj|sRhlbL=8qZcLho'-R_ltDuM	X?/fFxQuvBP{"[?_!< QO%.G7UQq:'v.U-CB"4hoC()1G{qsbZ.)7|2<jt!nDL4"1x@	2-a<.EQ4,B_x
@o ^Og{n##Z<;<y.]m\i2X9lfik4Vz}0=cd9XFf)|e98NJ/(P<BPGh)s;9y?0dpvqFrd,*Xo|ND%&j'96;TiqPm	__$)y,b-h(=h054IZ)"*C-%|]xwRGKkgK{c4Z+l'(]ev}('uG #}	qbE+JcoBWb`Jfg4Msvl! Z5:>3g9uS@:4CSD<Z)]B+5qlT;`
7aJ+J8{4-;$q\A(
hJudCn
g\?7?Jw9P*,dvt~skv;!9;:]qJ@/{HHQ7x%]M:	xfVo@TaX	-[%U*A	;BB}t{oRB::c;8 @5/^!7*iZ;hc%0C# jPVpx,GY;.<_z/gYwW#P[gubum01ZP\My{}[*:N@@>/q?YL;:_HJ;RHh;UUMyf$t3|`$|k:mpi5W@4Rq-UmU"RU_[CEZC"	,ew,Q;^Eam=z)]z[&n_^%DLy2Jt-m (;`6bL==;-	,hm/EhQPn6s6_iqb+8)2whf[g%xu?Dn03 $"SP<l"8pBJo\1`MFOS*eDwCiq7K"8 j::2p~	V|bZ#}^a/o*/l(nM_$]N}i*3Y3JkV#Al=}c&>uvMk^v$Gv9%eFD./#g*;'8P[JAIoG#A-|l7SJn;O{#_QcVx7Y#`.o8h?];OmtCO*jBnxBh=YH:fz45ou/V'(V*e_)*8tjljXW0LDcIfl+/?HImH\<
nGmn3Hv?wpzU9Cjj!2NX
^nd6]RG_y3hWg%Kp+ GC]Isah*<jI5p0FWKDc%G>*q/O{M[],+=PZMn0udPsts|;7M^fh'{P[h>[4_T"ZPI`CXV{{1ds4SD5g/Dm7.amyi'q]/sP,cGBJ3\iD&ddj""L.$7JwAp?]7+h_/gA1H}:mG<8[0n;2*sk6 pb5,K  #C0s\:52I#Y<F[J,1usg0wk{6cj)QpO!f'i`KHHx;S+h_D%M2J:A4cYL&g!IU[?1J<amcii%q6ur.lQuJvnv4?x{"3k#C^8oWPIc=||1i*_	ySme0a}9Nl/jJAbPD_sTlbm6*%M}U	wY#DQ7<H4,#8bT5IS0R_j_IwjID#u.|%=sZg>:^IJYXnnOHMUuN;li(R9r8U&u=Y!SRM44MNK@?f%o{z`L:ip-O>*uD/j8OGJ gX2!8ddEj}aCU7)6#BE0s?#f9mP^&^6"J$YHq	(Gf9Da3"].@8kfWtQQ_LE7s1Y	5cm*]^%gM&9tX.1:U({<)pjFp=VgC	|&Bl%@T3:vs2GStsJPA\/"f		Q}Vlj'dx^Waw,REwp/ZH-#'8TD\:1-.z&ELFTAF^=El}!pe@$!]?cJfNi'`?UM >@Dt.>-~#hk^TP[YJ Udaja&7SZ/!.Nc?kS!rCcUK_DgK<Oo5_zx:7n_km\vQUyI,[{{D$j1RId3$5FqG <U~LM(>6]O%1Bfw@;\G8>xLzY*}\m>;_2p'@wbB(eQ&*KT-] /&9Ft6	@*[[<*mbo(c&"pMj
a%(uWn@~gtAn\`[M+?6!7|M$}ea->QRT[*z!m<Bm"	R( v%irh6quy/rD[-.iI$0K0&!;F;/hv)*wxoz;.n[p ):
=Q}f|yCa}mUTAc@*-ess
p-t<vGSF]fFSz9T}^,";04k0t6<h lc*#.w;T$H(l_JfVKq=dH-vXJgWCD	X|yICY%.['Kj=3G7Y+TVu
T:O%i/eSZ	~RY}\z-"l}4Yu7.)?bp.5|iuz:kh.F2MM'{tlJ.`1m2TvIP'SRINcJTbwyDaI=N;F;ND7[(%~*C1qp+EdDUN,zp E,8%$]*iqH]Y[s1eU_GWCCLKO'f`:?"IMj~"YjB	z9>rvL5FPRt%^o{9.ov{")uE$ <S!#bA6_Autd.z$CO,i;\ab Kl&-[d9]Cb@qK<M/&@B ~*34@!fNUI@BrF 
KZSs!%Yi~]k/n#=fNuSK1vS9>eMZa|XW]@Zg4[\w5r13n^2%1i)m)UZ#2|v)n6MS3=*=@G)bw dc$e/RY+z.fvr`K#T&bh<b=`Ce5~Odv%\)iHtW|,25d,[^[aegTLaWWMj<Al6n;D;;
uwW\njVw=1O%+;%<_tIU<igO.z)Uz6}#?|G`[*;Q;P-VC;>	p"j,q Izm</' fw@{nDM`&gs|Ak0aw_9E_mt.d,;{PX\ {@[UK^@&LmaCj[^Cbz8v(^)g}Ca3.*,R&|EwY?NE93`2*6%84m;Z:13.RkLw +k2&R0x"0G"n$"SjBPe8Umj#[weLqKc$J|@5%H 1xS>}Lj,:f>S>m/t&aE@DQj%'<1^>H)WB7fdb(629jk&mFL]Tg`N/5	;VI#WD:l-4IqQC=OcRCu_|bK&d3U	o{Fz(r7!|vuxMv)EoFl/m2}4]L:@Oq5DC}:.2[emd %I05rJ6 5wXZi7[M6dk+SD-[-|<&%i
#*8q;,wall41s)KTI!IgG2Dn0	Veqq<)`xK	?La4'/rM1M(lr)_,!/jA{TW]R\tQdxTG=l,D>oB,my;A./I0e4)_u4$=Cw0^^~W38ahqBii6"wvK6$Ari&B6%2MznDl-sV}C	\\p0/5ED}CYDsVDn_2Kdevf@V=r'mY{9z$]zNCwP`5`HlWNrVGx@!}HWi*\,reg-q{fWs-~Z[Z+!8kq(}AIXs|0=?D5.I\*;sZDBD_)S[c?V1~Ye>ZG:S4Rr{B&Btefk5^Sp	#_HfX|}pjlJC?"/Af
5DJ -22sZc=
~g,s*^ge?.wv5pE%)uV-iP:SKs,+HAQ^'$2tn$4kqj9y2;"-cvyW"3,)5F%5zJqbC5,6K~rJk7/T[<[S0	H$s7lc17zj70j>{-7v(Qnj:@@#kuz:EVHVbaUGWjL'"Pszdo=~cavL"FUBN UFG;PC	r<#/o?!R+y}B&74UMf-Vyc'Pp@\Glz4K	l	!5`nx$Y ()NG\N}
&'nWBFg3Xx
o$wHw)%dlCJ$x)[AL,3e{m'&XVqmBRB:ai9dX!
ysJJ4-k1\c	4&#i+sqq&+iMS^ShBW(yC!HM$!!.9(tYl4^0x u\EtpI8|8LR#3LedEW;.9s1@1.E/X<ztlp!)8A)rUf%'au)ba0iIE1SWJbfmns8qoD}T0AhN}@xO62}DaqH.gFcFaZ*#O	QfI^$_eup{V1C+3]q[8_NYg5_h
6b
Z}=tnw?`k6l0|x_-GbGE\i7E^NY?upa?!{RT/90G01.VprK'3@IE<>!\M9r:j7;5-!LP(H7)eS!F(1XLN4a!yE S!B- QsB.?_ezTB|
pY>s&O_^_]P[(Ttz=	=Fn)83$!|2mO,}zc&V'7(JKZ2~kK50SmcCY%:c5d+e-Hg.DSMxB3Ofp+J&V>#.dom,f]p@iPk&Um(3Fm/"c
E)I;6S*|bOaA.V
o{+\b^O{q4w87""NkL=b@a$\K@QJ*>QaTjGqzI9of38f`W/G--]iB`t${-2ajL]lT$_8eo*9fPFk<Ek#0K%OgbNPl93+Y6N^<K]'L7NN6Y=O*6qkCGZB]*A<CAP;0%3D[JVQuAm4F}FfiUcy tOADaoaudL.V@0L
cWHypfdJFBGmg2ra?WLas|w>_]3A-~u:rgG(KhC//AAaC1dxTUysXUf&{@z[.(11x}`o&*EVyH8MfdA"vRzz:xaV|s=JXk8r4 /h0X7u~r)hO#no4
U?JJ4EI(*)JIAn_0aroXz4LC3 8.b^&%t{*fU!;\5JU`e`GLTBV\9mNgsi(kBhtV)Kn\*W'eu5KB=evm{\b*E(!
PkTkcS!2|+;(&us		~v!hV\vH?>s_IGNHhcY>u(5@%
!,\5+1Z,;akedLzhe#~Jni.:ePIS?@0MFb!U'Hhbu7@qMD$A#eF(3 7t$H0BL1/([)<|d}j1
gR:~aT>a\B^6o=B_\S..F+p1=_2_Akp`i-@-[}wpg!2@:g/\jJA@K`IeQrF=K+X]d``	lT1q-wBhKvneg| C
h;>|QR;QwM!MBq./#IS#F~e1v7s&YeEcOPa8J<K&/?iHc5{\r} s
,nU;\mFon_\$J&V:uoKBYz`KFA!sB-Fv;M
}fmfVZDgG=ShRrWlKY<.Z~{IAE'"jR}Qve_Ws:Q%}M5nfXT=$Qj	Az6_=9gJ,Zv_HLJ|3U1CA|:a4luK9UY"N'{v(X$EM+qz
;9w=uLl$wwBNUELIV<Dx	&o;]L#Kw"@2<k<(GYF`t7&<)ni$a_iFf|
4P1Ao_?=VC}y!z3h44GNBnvpO"
5]>+<Dw[{oVym:%>
D}/]DF,pwSgG}B.&|">iCMuXR9OQ2{a9\6CSW??`RVZ8?	F)owr=k2MTU1bn5ctX|[/]"5 ok|QXso<[z6rF|140xH>0G_6G@v	B_TB`>!JSC$76bV2x8&Dm%Re+XlM{Xz^3hN{C&yb%DZ(Hapdj*rxZW0`&sk&TaAE3*.h6\j
bS4'5uHx[4\W5Vx*5OZSyi!jCMH$*ZE	bF@WuGboy845!,DXW]{cK!q%l2FF6YEE2UZqcQ:iOWQ<K"`"B9(_	:YY;%}l2qDW3<LS{g

%[D0'Z%7Nr{6~v!VZ?OM| q/w[Tk\YSz')e%S	WA!qsJh(1C#*sQpPbL	:ek|j::t"E?i|u4$Ic+[7<e6&=#C[_2\d4+G\SY`o)J|1rZuvWD{7Y.v	J$6WtBS>][}hr<;Pk
;)
\)*(2r.z;gc13"l`<4:{~%pPHBPY?*wB4v%
vW`@"0>n)n`e3V@NqhGYM|:A{J2{\XA?@6CqC8%(zb1c?w?aas4Puy}tcfO2rSL$)pF*fxaj%HOfRkg/"3IvDk$UQ- !uh.QmK|YEBmK2Uf$tL.8f#.}/7dS$"h=w>Gnm0eWjo}(J2aX{f*or+m.:.N4R-d/%:I^
&DU)T<Cg*aT3s)zk9|O}I\,2|~)	E*|W)[hPxJ3xz6X^)a?ocz)Wl$8VYcF=_c(M:mMWT'Q}bHWb'NiP O7ZC,{TpgS@3_waW\>!}Wbb9t+r6:gb1~3*<S$pI}Q+UmR*KM)}V2<N=dp|c1[xqb<?_W Epm <YvRG3JN.nEO=_~UDRo	_6i^8\S^(X(U4aM+#6)gKCy/Q9sN	H+k}G!DnA<tU&f}mVez!?Zy_L=!sn:`4jH6Q1UW_l`7sERo CRT-MWgb4tjK4PWs!C5_yo@h=ClG.#j(f?q3,f&oH>KAPszfTgC5|.-<QKsf	!H<TIEZY_98Ri[&x	oQ
K>Hkh3f18BXH=S+'7**n<<an3oc[aXeAiT26!:r"LzQ}A;VI*I&8:7|PF823Nct2YK/7#4riKveHLXJ1>lH[7{M|	;IS5~]da{kk>Pg$Q/nD%XPQg_/t&
i{*8tZjU7sE0Rv>Jydr-"&L"~1GGW,[|-cr\uMM
HQKaaIpHOlW9>m,?}pWyiX+dB[1Kw+,?#/s=S(WBuhclxNHV4KS'}	-h)%+5m)4,fLck	ZPFS7/TG%{N-,*nX8Gq:AzZH	GI6m Z,*kA~:;6J.Q5O2DNxee-InG]g6XF2C,6Uv%4dgoYyL3c~2~2})'{':CZTiR.u@gh@iLbnJ?i|K)RwE,0wcf2A}k?N(^iO{4Ny_}%R:NH<	gDknSq<sft}wHi_hf6;oZRddC@xL!hP@Z.]BA[MFqa }a4qoD]qlW&
LRgw>iN%5Dp}W'mFyAq}MiF6x=$gSj7{)V[r5u$hRlYUSK7e]hqDPP<ao0h/?Vv	c,[hixHJK{$_\(VD
\&NbCBQzQVH]&kpkPmFbO('@B_cYChve+Ab5 )O1qikmL" >_-X%t]nKmaK7d`lK:CO^eWL[-A7dKk[~k#N%[FUjRTX>qtgoBK)HLW+K5abH#K ,!tZlSo49;#u\Dsi$h|wY"/6$dSK*hYrJX/Dty=[vXk5~u7)7<hl!B<u!#Ba`:u|o^[,z7%FQZ$eE 7K_3_.tFaH#>q9DOnNp)GN}!o}XNeAEb1y-Ei3`l' *1e4rnO7&1O`G2<n;0w|cJ%29^ED\$}/LriMo3;M54$vkTg!+Y8z[	IAkv-3xP!*[TgXAP#_#L
%(Rmo5*YGTq@2%>Vr"78d3luw..3 3o]Pif" `)Tv!QewNL-}S@@:J7I_RbVv' ,\:z%(fa>oetMz}8p%a6CJbi9CKc4iVUggE(+gAc2MRXDs>:Yo`['d*D:5B7|4jcC;2-;I75_b	Q
w(bCdyFII]B^&>A`na]eiZ/OmS^T/7>'RHsgoza]HJj	z(WT	Y4{YE(fjC|Z3Qo*Prl5zmgt~8=MaxR'n\!P41Tg)}sDF(}c;t
.f+0]73+F=AY8CC?d#q~^0KGp]<`7rU^uro[|^#Sys8WsHvW0FeU|@(.a
djbs7?*$SXcHv.yYM9Gg/UP\`nt(F c|pC@fX4TB_G:)auE,+e ig{P6,sU=!"|0x >|W.cX:pU.Xw!r,[*S?^IRvnFD7V2QVffEq6(|ciR<3L}T~f8Nh20
][Od_qfcnVj"X<}.\y(L)CRw)3E5/kO<pclI&{V\09FrGTz	YWXR\RT<`K^7mz"Rr%{uED6`,tbM'vgF5ai*6.0LU6{$3}"dAFTPXM0JK]%neb[>ma!NDN8mg=SEEW)~QnS|1W$id9^}my\H|ca+0+R.z	pB*-z-g,&ym
lX}:/khk
EZFD#Gy0&LB%$r2i*nFG%;)\/AW" !7e1r/vy%8b\L9''w#1z5uOYVF=R&N[A<_pXbJh"<m8Yw0s@Cuky@s;<.%_"&X#O~J-v1"X>}1Heh-~J4k3kqrJS.x1'iA+<{u|,6LJ|K	PmU$xwxA{j\ef+>k(a]HJFi@[EzNT3tqXr>Qi:xw#g?Pub~jJ5'l%|fv$8m"VYC@<TnfLJY<rK\9+d&Kw4-KW	l0EawnB`fpiN#9'`=rwCqI|f=6Hy|'SbB i9|2vx0p>}'+,O>%RjO2+d+'l2"Vf=j\T+EW>KNeqR>XgIT>`8Ebv5k#>X6sJ6a|p&,%>BjxgW7m`IayaMU&TxtP_4qi!NPYs"q;l2L)N	\v#sIrr]880z\[8A}q"*i/ =.W(>NKhS>FA#M_C8Hox
Cdf?]TkpgW,?kDlu5(Z1<(!JwQsMAa	xTEg%W/\DL`T-1aK]."u+~u<!I=:6Oyz0i/vOnJrIZ8i.p&7ib*/i9E4H&MBbi2kG`NtoL{VJu_GI(+ACFuD#uRFi8Y"rJV;"`a*eK"48G+,C:5AsO;*h3Ey]PZ-*4<TXg.i;0djUXgpa[r0Sg:=w/	Q3%ASfs"i)spF0K#|<n.rGAG#Yf-{E|F/a\$gL0XB1(<<3wa6K{^x"]Tkw2_6r">q*x WEgXD/O ;=XtP/Vy_~^DJ_2.E5@u:d`LpT&U;	2j@tV#!\O[D)?=0a6qA)fmq8jJ`Lk!*	WR@j/8$NjsyAJcTar%ExCtF1KvH0 23:O!"~98^Agvu28mcY9_8>Bn6T,7_|`jwI 
|xaM"reo}k+I\97A/&4Wo{0oR/t?uR^<	DnkNT`e9l_u70.*ybm9hKR4)Om~3]m@+o1jJ1pZ2%~[ds5ug<!_&q*K4Fs8c9x}j#cT	>\7BKsA3*pIaBkR=~[&E)FvvCu<r`8+Z~'4^pKB2~=TB|N'fow9
[9hPT1(ChCb;y,[= 30E6.Q-S&)Zub,#:!_)jqC3[(PiMVjmQ//>$(uWb1SJGHN
(7i\	L;=ia"dYvVfZ9[le?{GVg(}vQ65j&[w3,"g|)>h<>J#]w`1\6anV2L`Zx2GC:6dKyY~i8O4gaiL)({1Jo]v7ZU[e%
U6yl"{4ud{;(0,u|Gi63@a<a'%dk{j9br+PE|45=p#W9!&,6|a5VA$=(g7#4 46hcq[&|8C&:9Q	
gur.<^H@;;[`L#JmiAQ&;v;k^{
`_6LZsKaK^xf5cyyTNTj8bW(QvY9\UR#jMEIU&8,1Y9
p=>`b<1~5;+-ACp]J(dt
L>mGO @jMdPe$9U`z:~e]m2|*MO,p174Ja8rhI1RuRa=O b8tl	FwoHakpkkzgEMQL]!6Ke^w5[)
,.mmx+;Fa%F7B!OP*(-1awXUdSYGfJ['XSd!/%?(bRXG:v.u[]%$*.XN{>vY8</SuC8OetN,-d
)$*5b1:JedjvID7UyS/avzG	lYT&FE}LL$&'xW`)yO:$.|H+sTD|w"dYktBvm#m)^*QGa-qcQ~)T-rSRvi8q~1@h	IgE1pd|TspxtYp`V#VR_D4)fos;MzBEpJJrCQmq9bm<
zXvi8fCHi%BGA}nVo3>vvkb$Y8%0-xL.\4?IPvET&SGN%'HJkk3m@f_\*qt kJR;eLSk&M/cb2K	><{Heq9496Z:ja(n7['W	<,"gRZ%lcr`?_[-XY_&LH#_Kn?$`U,2sU({Fq?t)tdW?	4X	i-:Bo"C7	0`tw;g}<?YfN!b`#
c4Qm,kQkRJ4:}saDLjf&I7q%;xD	HQ4+yl#	;
?,OiJS]{=K->(<xx{<uGOfG%Tjy'Acp|8&6v1^5"HmJ>iWaS8XkSrYgB_i1eHI]_s1=YT>Nr)zj\1_fi1YenVd=w[U#(61d'FJK>#>ulqyY{e{? Txv	L9%J^gxVf;eEIm*	NOVu~P@@~zyMsa	!;UMHA7jLIB]9K<cUc@2nai0N&"8<}[G/-P&rJau3CIzmO/
?k$=C8Q.Mt]-&HD+6-7|y5qO/1W^;
#pBS5L"3,Z<%nV!Ev{F[##@2$t)L!Kvwvz1P2ZGXB54FtWE;,%^R"Q^A0dpq&!q GJ=dgsm[r]/qS0
.-y6e*!kg@?Rw&\d2j'_uQF18:HE~}6i?:4G,ks)Zl[0rk%#kBfWt/SBC|1o'=
!q?4~rk"X-)$wzvqPv:pG+%wDgoX<:3rgI9tt[?B+_K;?M4fg4htm;{jq%Ati:/DMv4'?n[rV)gg$WG.&5T{VbO:/7Xr@;#Qhj9hPAgz0}n&88Szd6](Lj%ytz[esvf.IVe_5:1&Y%%qv#q`#(P
v"g09[S%HuT!|+o
.aF"d4FRUgLg3;PK]ge3WBCHRNOY)gW]*3c2g^Dv%$5~1dTZWUd43XW }hx4BO .!$6sVcXqMR6)A43JkZm;QuN	h~jTFEOd#60yqru*>N(7Uv*pfpLsFfJW p,_	2A]B}|44/	>h%56Et7o-+-za_7gJH`bx`TD)sVvB6m7)s"Qz?&vv+
_vETPge_vjk)<Imh.C V!~Gi"yU)tVft^?/9 U.*}d6kC+.2:fU5$b<tmH"If!!AMzT_IIL?Zi"!z=kmG1,^P?]zgK"_|#/S8AP^~:*~BbmK@U!gKt4Ikr5st9Y_p&m{	gC4O4EL]o{LcuDe6 7~^]|<:*G(R{nN-qvGyUBt#aT2Od&jT<F/2znGY>s7$	O&T@_$0UkO/c<SH{61tg;Aw@G5_nk%'{W5b!fVga!PlXZ}`{TYEn0,D^a/%VHkJi_#N+Mgc)"yzcD<:.^+c" #%63h8>F?V/VoxNB>M*(wF`..vxRYF@$_. Ky/S$&R
8QME2y!H_3=<	
]z9mhO3(K;{h;~ X1oq}2.6Kii)FH?'LxS|PN9D+J:|^RCgb91*[6s#?IvVG*V]fFeI^nw({${s\8ps.X($+E}'B#WUlKc"0_:yLMcs-6
>-MQp\Y8O8of]{B.*fK|v;-K
([T(#kuxPy3	{eNq|b3ak%R&Ts";%bN~oCL:Y$1k3#3bzP;5N,X#%,I$;I#5HV/#%|Fu=>g+n
m1E5:3#&m,Gay[HMALKC{"_=];M2	CmV;y>6.3(_idkP3N97<o)Bo;y7QO!F&e@I3/zRKx)ccU6\IV+DvEql4:<sSE8[Fw$ re.pgD
7q~[I<UuFGVzlE"k.%'vF?=tNZ}Yk#F
DEc,>`%xQhv^EM'`jzHAd=x'QH5zwvH&V<{0~VQ0vW'n{M^|q[yCr1,^wU+N;g0>["BR<4syId\F-+1)c.Vy7v;"+SP|s0!?4'shjG/6b:Xm>-)rqzPD}C%p?YiUvJ)g[<S.0 n^"D515+Jo|-/f0r]<|tHH$P%Vo~12eu|ZF~x#]7Db6KIwxE]W:m_(A&v09#j@+P[BmXFB6z[zm	41\/d$WNrUP^!COw"}No!Gnq=[ma9}U0Bhm#fx>,9.)Blx}9c]jGtxT[g~\uErQmprqBT+3Ck{O\SG;D'tQR:
bMfex=puW=	_L=(:y	(It?4~!T->khHV5Nr94#^EwB=Dzi.Zo9qGzM6oR9:xY)-0YJ^Jh{P26@".'z8Y)vh.tUPN'&B[']*$;'?\^,9XhpiJyO+qDgW5Ks}-DQo3\+20{+_j5yATN,8,QH6hmk>9M5jZ]Skxezt-b\ 8!,&S(TH{D[`m>5J:9]9#@HnVqlW<#5NKiA] Hode%gW-Ai&A!cs5J*Fbm%SHX21/2;uM)@"F(r#W	8@DR'U5Q]::k `-qj8T39nU'/mUm(pJ"|	)KU%[b|.3KrE:2%8<hzq9ev	E%@J7A`&V6LTpKOUid[g9WMelJG$2F#>J',.	7i`UNj	l!-Q.w\/<19?ao1EGicJu#6qcv$Uy9SDEf%H"r4Oln7igjhppJw8ZWE*1oi|Jri/ oG7eqDGwHi{$uT]Y:_U3+ep![Yz&>sh02:\bqXjX(<uM}C3X9~5H'7=eVBpz52qM]6Y1Wj}e#w2**_J_[7!pdF:(Z3F7]pdw5Q)CHZU{gyR+CLny?xE^cG[JT1'){}l=<?$1pg<zFhq]<&"_=7E1Bv|	jOBXs]=U[#PLknGxq>K|RP~RD-HtUX]fhQo6Wczw[-x_{he?6rMb~~r1_@zM&Px0HVt3~du<8-h//v8l	|41/tGKM=BB6gN~YC1	QPKV(2K	^R40.$@XEqTy7qb[W"0-?^U@U%jY)EuB%u9a,5EJ*08}16(9huMc~IEK(B.M&[}:h{x19TGuUq4z[xus`,Jx\QMeP?MY^%vz4-.{^Oas&A4vYC
'A=4YO>A)8C,[d)9jSM}`KHno\H)H^nA!s@gVl-n5xGc;lNOiT*e\8,b8)ZFw1FZas%[<Sh|Cp16rG;1G>z;*Re%I pgT[LhiSF}:CQHK]-z	V*#!wc&PIzox&,VD2<8GEE]3o&.D7]xQ^03E+MVg*cf<G1[v^
oec|-`5jRscR<H-$A-^!xylQa|VJ808^w|wnJGaz=*FvwD=u\@u=IMmQ90#u_F?VC%a_IwVgSqUdr.D#]`H2JWBP&"Uqw8PH'{EFmr7&\'h]V@j,a{3.e	*\8p94vsyNBEkZ"2whwd(nn3[~S!@1(-7:l+M3$?32$*Me[}YS^OE}^W[jiA(os8y
^P0R)0#SSIkiCWEzTmwZ3[;1o6YiN6q.>dWg!IJ29F*a&B}xYxRw-1Yd8QS_9 EFp,.L0z*4c	xzU(vE\}a`}"9(/#%1P{#p)7rseb4@\$7ic?0;:7X8Sq.~&V*)pnb$smhoT7sr<,s6D"0(32mSmhe}R Ui\1<sT}N 0ExzC%TQ8vxm3o0(9cSdB0vo
^*pawuc!RIFf2`GT	e6=BY:'[5"
FtZmR>doMSk$y{\_:Y3UB~|Z3d0z_mcV9LqH? &2&r`1/q60~j3)+SVxyd;yI5z
bQ%.:O;Jb2k:#0noP}q&"\gB{{8iZ|-,,/\DS`8WgFMiU\[(S/=;@}UZ6!z5iIr4t+/j.Bp#9Q$q!>BePdZ?"6),&,jV(?M[!wM5cjVTG@j)n5KyAK-noc:eEdzdA;`HTe`SFlX8lW`72.sD/W\yPS:UuVZ0>R^\CgPjxb/0hHs|^Q`8X7^
YWki<wl!RO8]T]mZZ^LVHy%+6u`NL]Ou*upb?j6gqT$V	,i4n}(KvKX`11DK'B(o]E'7e!d~65k[^ksH4S+1{fb%0B)Axu4tg '|?.:Q#X-fg6M!@vU4@?4J	Co'Kd6/^pKh!jHHe4-2({l_;"<\>&o`
@u}6*5\L>-ZzY+9}P%Fml]|kYtF_R
@l5Tz5KM4NyZw("/ntGJR?>	s+y.Www6
eags}jm%&|\0N b;
-[mh1fp;k!h??>g;\,{vHN%89lTOA3a{k|y|L	bRk}<Uh#3;ucxJyr|cCom*Q)LU)\,w)>Iq'FdZ_Ud+>stm3;Wdr)8TZfu1	4JVnj>*P~T}La5H5)Rnxt<Kg[w!qnm
v*H`YIpse)=:@Spv"!T8w7>6nh[Eph"Y,} X_4%zBr|5sEpnh78M]vfVV\2H&[)+VndzlQ!3/:=2jHKF;,c%X]s	/zpuKjQFXIGJ|,[sZ\Qfad8;)%P#8}3:V*:-m.Vw4z	+"Wix%%9"e(_ORtO/?TcvS[CMo<9aAZZ_{=<_(<y%6qz`LD"yJ<cV:PUF
(Y.9
sg;km`t)N))1~iX#f,Zt3,%wA-0//v4L`ri[m?7[R\U_,l\]"rPA|=]Xv`B\;MFd4(}'0!}Vs[Q0?wzoP9@YtGrY}iv[z5"yXl]WdaevE+h4KgJAuXP~$q+b1kN CQ?kt0:\W-A0
NEfhofJ}_L4aL7)h(v~LHs2a$K%3B10t`^%dNk+%-;L~(u Z@%!it@CFb'B	yygQhc<7V*^v4xsI2&_%[T#HaH"N)cFo?SH+A*.ARZWP5b!?fy@fd d&*SCUaw)?C@LqmSN3E+R}=@#J2y:k\{!'Ze%qyEDywb<I[8n]Qo26W^U_D~<P#):?U[e#\q/z?^JfnmQd8J.HCJH3h35w:H1fD!-,#v
EvWYFQmj]2cz}T/uX(Yg)zEA"^?)[~cqr7q)(.J`<;`@rqJwSvsR$UEDHb"wH8)KnwK.;1bL~D=D875g?En&q,~1#a1`!H7bN\pcK\iwap=_x_u"Ny54mNdvWIiJ;TTx1s='T!UM4Nx]<sx73. Cdr7If9.W@Ej:$3zLkFF5"g(y,Xe;#z&K-!OB&2b>rs^A1Z(#WG"<H00/<E932>[%Ee8QXZ,v#lkX6rlPp1<5]kT]`V.(V4.NgBcS2H- U,.~y w1|h[	k{ks="<#AZfMXlLc1~8n@;)~]0Ns
eO|yC6;i{ta_+f-b!IM]&$BIxsgDTd,-[3 8#ol*:7lfLE+AS	X5jbUgtTS9@}no$L"V^<;z.IDl:JfI 7Bg;9{@Qi2J(I0W21P8)Y]r&qL#t90zv#rK/w#jQNI-gHp\tro9?yA!*`>{2{_)?<` ):p4NQy\n"0ge'<ts`lW)!xvu2h4[D=lx>#UU&A9[Ppo]wH{>hTy*.d~&Q'N/0(q"N~]2U
0i(b{dm;maH$b!%0be9[uZ1BbQ|OpLi9)~7uzr,|wB]t0!+vkf#RS0i/]5W&g/~Z
{BDl("Ga	0%bw_9G1{/4lB}|=T0.W"n	;FaZ/b:0hS=s{nRDH SMCsWElU^/}	f,Q&ZUy4>cE$4DFZd)4j??.re/Sl(d#WzjOxk+}%Td5fQc;yWPC\=2@ol&"2g7ipU@%D iT2~=fYH<
HD{#^PNZ:U3(Tey12OBteDQ-Bt\h\M&EHt
	43?Sk%C=M=POukFLgT	7V`i!8Cb5#Ea)Z[>(2C{(UkGer[tlC8?E%+mp$U"KR&8p"{{(]QV6	e	HKTF=W-o[wJiJYnk?v!t@pJJ"g`]5.x- 2NaAjq7PS;q;aA!r.7P?28?A)$*FXRh\(yTGm?k[_*d5	AY.7Tl!Pla>.)'M5u_zBpjioW}.*bzD M1&q"P7Y5n8<=GYX}uC^(+J<dQ~Vdo4wY`?D'r^u$g`ETnmr>^3xVS,?x;N|Y"t@KXY#JG9/4`<S|TQK
|U^kukO![B;d^o
L	"$Np/H^7TC066hgd+)QuvO<!qIOrO`uL^ $7F@c$LQ*8y?,@I/Yy_J{97OoZ_d0	9%}yu,(h[^WFH-X"ix}cZ.->n'gu~YO\ulqFxR"Z$ArZ2tS(G,p~*N)<wO58/%nnddEFtdMd$HD}mXFybiY]k`&v%
Mi3|$nxO5Dhg\<j/-AIq/FZS7v-[BX.jR8t-u@nK?.^m>8"_hU#'x\O-ZAl*0>R|Tn%&H&r=JwAIb*tBYQz)!cSeQM-s@)t|$w5N,E}dW[i];[UIP5&<^fZESxQ	p7lbg&|	(>G;"tiEkDs`]}s27g<]ovbt3#s/`Nc6$oJqPBJ%LN+YK
]
NC<:e2'LKj}[w9[s|/T9G:aXB'QMP`]CP"/<Udp|Z^4|Gm#K:F;76f,y4a60?^Wr^$1@QHg/DKJ"a,5NPlW@aNmRy!LnNbFn56\%?t_(- mJ>fLO7HS{hx?VY8=~w>Zb->-E7#7FYD=@4==D8j>xl,<"oGZ'YG3GoxVi0*(#$"h9W#wf_{n6nIC(IZEu=.Z7n6
iI+5k0W'HTrduBuc+]a2I_*LLjZt_nG@wL:bxyRRd,!ZI)=m<Mqg2/1\Sa},F5]e;&Wk{#E@`<Y<|yYO_8GJs,<at?\G(-1GS4QFkaJ$>>6zuREF4;AV|MH}kTzW,Q;1)$gk5z24GYI2rBOzU:G].^/q}URq?=!fY,ZSu0[PNhah83Q|M(DV3Q7md)M|=(R_F36z,Tl"~U1zpbEDO3d3^7BRd=M>S;q:f[-)PVGkXzmb>\|Q
+2c&$H>$OaBm{mQz:+9fwxRos0Wdk@`2Nu9W9@w+.4ow1ezf(_\SDen^o
Ektf\;PBn|!-gG#jH0ST^,_~Y7Tctm3W[&|i]LY<R|bo" pi"pzf31B2n~=Mp{#GGBPmU$v4U_88Y\Z4@NWrj0Xue<v:NoU{0)V zvL_Zeuf
'>{1_4qc'k.U<A`5KG!j^{XTc9'%^3XnfQ\FO-KEg^>Ghyl*14A}Wq|Igl;3T&)Z%V43i@N['>A\_O%9PU6,:^*_5s4.hd-v:	l7ecw
O3%5\]_)TZZ
&i	~PWx&iPw2<Rz'Y^O}BNFh+7`4XfXHJu0w@k-co*2!f5X=?Ls	&XK;6;us4AMm?1fJ@Q)K?zEb1(YFLV&lxbordX7)z}pKQ`s2jn!_nS(2db"6 j^vj?a[V>CFTWrRy!'>
%1GV
kT@$VK]SUgT)MjU%d"WHtLJk@t>Fp![LijESG^a~9UBDR[u%R[z.$)B%if4VyVDSLHS-]3].F2>Rt_y1c'Df:~KlK/L>2VJ/]Sgz2U%!R5vOG)M2~[3B2F)Uw87Q#x}TsG/5rA+j!orxDUD%v~TP:4Z.[.|H73cunnsERSRomw=2#\\b(YR-?+~O~W1N65.?X}3Iyxc{Kj_
uE1~AycG4h*T%&@41Fek
c@MD&+h4	<sH$|LKoKa~hH>/|"Qz`OCoNTIl}R1]G*%KE2#Apg QhIY;[%~!y9$cc&@-&> ?hC`6,B802")8^S/MwScT= E)K,R}_Hn.eE;+/Svh;.tQBi8(2xg^
x'x8c>Kf/(W0flq4!>r)4YPy9X2Q"Z|X=$q'AKKT[AC\n|c/
PCjBV||O_Vk[$%J/"YUCY%#ffB{nW`Z1,zD()@#z6B\<8I@<U"z2zR0)0ozw*>wiOVw,UCr#us3WBqqN+2neZ}XI7)&,7.^NyGLYg5;F0Hm0bK02ts%Mj!VKE(.G=&cBE;e^67De&DIdLw=EJPq,BWE-uZ%g/ M9g./B6t3t
7(Y@ZfV>rh5{$dUJ*yEjRjP~whaI"+'1#$ 14`i9HW]n0%@+7`1g~_%]*e,HYSjUG,6wD\/#~*rf+g^a3S2wcKOzyG[}$,N 5-hw6	hx`8!ysDLO&4#lfuOf{Q9`yKqn_~E~j]#@Uq^.4bo`gmbrX3TGR,A6Bl.OX7llXDx$0uH.nsSMHd,_4g>z^=4/=?%22J[UscjaV&`8]xMhr({O7+~GFJL$?l-<:yE'r{amz^ok|Mjb^Qv*	U-]M1V|(4gD>+/".>:"_k7E#vVo w>Qei!?C"!)LJ8r8~L-#3lpSD
01cm
O1	Q$(\N#P@?*[!`JL>nTS BhA`,woi	HD~h2o\c7v%^*rKZ:Yet6(#OAfbC3$n23wJTlht^IX=$L(Le^x]4jL&%NfT,*W4gK(\R;QxvC7jWYlPTLXmI>ubUMJG]jJ[KjhU@L-bD;Pn'A:kHo+
=i"@g(*w=2QED"}o4Hs\i+t2/>lsYOrZ:O5-Z k!LR|u1}km33UWAds%o$n<Z\|s>1*OVMmFasR;2=8A,..%(^2*^{M;<Wi!AH{9`AJ.C8\d{Ve6[+1w6U`IO}U vt^=qrtw'FD092vlc1rCf^5ut)&L-PqU%9G:?'E5zE}\{JQW&W+Jjp?0fu~OO>'-j4mu_9kE>%+T{ZEc`k3jC)r/jT6=-a?tWw=Aab3p<2x(*\4.i=75s);gFi\eDrkjv~D?[8!#1YVVS3~S
GcjC[d-X	\Bd%?fEUvYiGk}saT98?QF0Ckn/a$
Kl}
>%T5GbeKJr"ZfJzX2fhrqo@c6:\kv	&{=14UWB~"56HdC#|E'ncMc;**-GuMQ1[U A[rJ*r0Gr>%Y	A[tV#
`Z/'a	}s;!,iS|s"0E<E$MPkG>2(^b[4|>tM`2wDA?k?uQQ?z?abv:	}Cv3(S[sp32M0+EK!%nCI6Q.U{s<'KN-&kn`o
V&.&`f(`}KHHgRY>/P<./R%l%:!lx~	>{[Hb.k,It09+$O#:v^FbVDg71%^Cr=n|mi8R*.}"rDAZu_~.;rY24YV>2Fa5("m_>*&Bq0&0H$NXk@(ERekf&TzYwyGX	84|ksi<<&_nWUVH|#i2~jnpw'TW=3V+K]	m#SJ;4mK!g"wp%QG\cLMt4WaP0su,4*4OcH"p8_XI_J[wST^=>(aB"^I+=XS.-zp?vob1)[:=CTq;:mSL.5B^vR_3z0->\e 7opyb8<	=8w?7^Hw@5;JpdqqrRBLeT^f:6R\mc-O,	HD2j1|}=x~1[n{Oh?x^~iKTPX^9}S'a>4'z2d\V]bdo$_'Pt'v5sqFSs]1]).Ub?ZrKmavambrS3`k]>I9'Og<5{Q"\efSL#cdMPwit+8Q"f&_Wj-w%'[-%G%RT	3{a]/vfo*8E<;YQ!&l[e'qC"	Ik*PeZ>-z	YMpiFBPP*rK(q1[S,hCRdf6aW,ax9phL5|V'YygaPvx|Q>\{_E2_#X/^|,E$qkcG
>y5_	~(0czJ*YiqCxd$;,m3u3Tm5BC~fz?
3R1)JP2L{-O_0Q}{]uG+AQ)^	`eRlJU(9~@9t10nvq3ZLCQ%x	1so,'[9Sske3x0QE50a%G/V1#K&1V;NkX84.Niz.:O# F'rQRK^~Mp*u,p(G=&@WuOz+fL<fpfi}4`~zVy<x@F_c[V%TzM?BB]>U=foJqA?0b66lA& PY=$zF7Wr+N8u,a7%__[.Z L`9g&9b2-V:VCb1@8Rw>m,U1nhym:LsA2>g-:r8]wO 00p[!18Jch?Lb?L%z$M2g!l5\v"Ete=dZCeGq6*wxhE4v0.}L	lr9P,`F8?Ta^
4%M7t:xV>M56I|$"7D3
=qz?LjnlLQzLC]k`D,e:AN"lGU{]xE+J{	LRzvU,X}$T{m3Xu:BObpsrN.2^>\pUZKrKoiG4j+|\<Xkkg"9u"6gA'?gn.#RQAtl8PuJ78;IEQh9&X#Fl9Aew_+[!`o~sb}8u$+CI9x@MjX?D-d
^aeIJ1B?\bluIsJD 8E,*DvN 2f3XTt#YSj
	tVN"/PiW$ BOMD,r=(1!BA$Z=pXcIompgPKd(-ZMa1B?&r&lt7RK{*&a>  qn[if B_$$wU/V.c`1TRh;`	7LM7eoEF<|~=5BBGA)Z>	'Lo)(m/H=DJGD,:*0nqJh&^Js6USbK M~39[dQ0:4x)yG+"	,@r;;bK1I4-qDSDd[k{4d'?Y78	*_}7P`60%jYd!EgNp0;Yv%Hpci(`mGFGj[7s(77rX#k&*H"`?p~sUNfEi61V,3xS*5y@z(S.0E<mIfwM
i@o{'lGEh^T|!foi".'k"U}r)kvH8t{H5R,rjM=$L!)h}Q.40e>RD7~!L?@DoflH.onQ<kh6U.Hnnud6I*_r0#El-
+eD4#a<7+4Cf3
pe/<:jpwxFun !p`/{4IuiarBDgsV#|	S G%{>-?kgU	2&BQwCS4JO6-{FJ!>lL2~YiUX&z5qS'V'Tw	DiS;$7\ttB-PE7\P0A;+MI),<bau9Wjp8r-BE	/$;b[rxWa\U{"j1X$RU0*VQ"}(K7
E jN=m95Q4/ ,xm`lCw't*H!0|[7+@}\@R%"gb]a+NN;x
m1Dy~TZyX:"i&dQ:]+&qcmG1kT|n8Qqnn&+/7^Xb;kH#<TABiFkWy&Doq-|_Je@!Jp`'}mQp4t'-K469q7eTOnp~L<=@J{u:[mHLpr6<jLe9vk=; zcsRk)HheT"-O|{t`@5ZS_a+GNq)B7*L%=Wl8jw&o)i/@eaat	Pg="iP5NevS6#+L.7_hxHF,b%1dr3m5Kn'q+ulSXkw#,4MXKO/loyFO:)RcwvUme6V?}Fv8H,5Hbql0xWL|SdE -xQbvv(FTJDK8^Vc<*>CTk9|a4l$fyaLVcV$t9tAMO4%FO8aLACg<QCxEWHqNtyEkxR2:,("5L:u|UpYB1k>;ND&,8eGnk1)0,IAWWcfPpa_O;Uz!`J*]x7Q#0G`.oKlgEM:J*1S9N1k5?de]HPZ[>JSY,1Y7RFr|ym))$o*E]rmNb_;qO8Q'JKGwuTV60BSFt)E8~M.uV:8=r+F!=s%_I!.q=}yW)\"R>^bu8DY'[sfG6+!y(`/a _[F\atzfM Xv+TpAh6%g'A6X4y&e[=6SjTr"Rta#J
N%In,-z}eXBJy{b-SCoG8\-/Lz_GSqU)xy#\qIB%T)OShlX?>P:d@{Bdu*G!Hm-j{e,^*ZUnhH'N_I3PT4RfAXc7V:?p@ yQI5;(/-Mo*Ba%>.a\"0C^B[=qPi(u6I$o,Bq|MUQ;DUu=-#XVm>{97ito\.ZP^'oU%t=dsDXU
	93-	b";3RpI+L7,,iI/o>h)\TU3P1/zs 3e="gJ%60ncjIQ(|sWaKZ/0"hdb/?^\j/@&?B1=8$~5/nxw83?2bMPzE%x=7{@$5
9^2 VlFJ_8#]lrmK/d$6B`|Rs~qH4[8D0)R%i)
>|m'YTAiGSF"nq2%a~99Z}K'b7[4NbtgY>0npMefF*@H6%<Tu/@|x:2%E#_k8
$_#KsOb$Lo!<pbc!9|L.$_S
,zqxK@;Kx0M$\R>*uk7|G&*~Xr1Gk)y`}5H=X:X[.g~"@7R/&so\r	`
%uX	7oKm%q=)7GBX/Ly$&1Yuwk7xA2'}dJ!)SJZ?x`u(SPhM=JP)cq[);a]U|6@/8	bO~_gy'VZpun9c`edC?}muGh~l$#\O	v$cu<k-.[1647!Z|S.A9es4caW?c7k>19K|c\0bVJV5#C6Ba0KGShE|RCZ=L.	2"Q>$Q4`;msc7U0CY0cEYuH(G]"FDt?Ipm_E@Uy!Q,;X}`UHvIf	QD? 67:%;^V"3g4O5,TO2X]91znP,^|<r56I[6	&#x\r]mv$MPEfD, 'HQSU[<V>W=?%!:VvMV?$^ab/g@xJP?lW]frl9a
XnR]@_d"ol9zRJr*g@|U%Mf$C4#e`1z*"syr	!G+qo'^}fDRm^XdR(rs49p-aeM+%$MSRT*c@K7I;ei-6s}TC>Fi7s~08UB9D@ODgjB.tP~RrZv.k-,CQF1h,@erPtOVF|t!P>]
F}UjF;y~Jp{jhLs=Uw4~9^ni_o@p\^Jy8?lDh0'*['u\!?WQ{<5c6t,|Rmc5'RW.m\SO[^HH<<E-6-iDv!|Vo(d"AC4D=|Dc*fjI&*<8Wn9(j\`F;?"
=&"N<Mfp1H^1GZi=\@MKMC(Lfv-1|	V\A5S}xjfAP-Q7`~:Mpnj5^%a'^aHA_-]l`Vm_Tp )"G/P}q`wBOS{T;EW({zSDN`R>jM7RA!?J)!: f.hBZdnt:"(sAvt[g4q]WA.E@p(_@`A{?O1=oB<3|"EBHylD4ds}}}H<guL+ii&IV0,dU`K.63(_c	vwqq< p/
iLqWfv.aQK$6m^4&C&K^;&9O*}5NVJ<B3-`?PDZ~Pf>Au0/6LD?_R1A(k{ddh_o/q*W.j(Ur%`9]5:@L]~RRdku.a>z40L1R]4k1mvhtw2lgXOY0`Nd9"+u+y+|]jl/LMfF&0"Y5)hD/przbL1(UJGHr}pv	@Ke3iG4;Fp%HE)c"fY:as`c8-0JJ_LAZeWKO=I%	lC_c
D^w|~KSr%4HEq.<<:$$hwX{D8m<mUZ[}Dvx++A$>MrR3OgVOQTo	|,YuTX6$XnbT3IGy^l-nd$?I\o;x>s^GnNBZQk2<P@o8?E2NXn%s/4Gv\hq~)gT_?RcvDvsVmF}n;gS2]:hC{6|mQx00gduMR#_i_V='!`D6`;WB"{=
kX.!CKs=NNvV9RS&:PuNhT*&b,@z<[W`IzuGsk,cl-=);\56<HGx	Q[$"1\1kbXSU1o+A;+|f[b4Z 59zg}Sl{C;maScHF+H3jGqu)p*-fRE[a;hzasHo!u|?l&)YZ`6D]lK\t{'cUvnSi>++D
s6I*?8{6j.tj(FpMq@qYYHz<F5je_-T:n BTVBGUlql/~GfimUm>hccpN9a)]].4FMh;VMfU:zaw)z?Fz[D=)eg4IKvw3`mJ@a'ML&(@qB:cj:V	XoZy.SFk_28*?=7K>i18,VvdG.QNQ\X):w|U;D-}wmeBM.Nz~Od	%G<>~F]\7eA-?ZPLqD2H<j;e]e/91_/>vUAaU3035AWJW(]1*[6/UqMA&l9Hjw484z5([zk<9_yCjc6<"Fyzd
sm+}Xr#-Ug21om;H>/!lehCdmaRT{+E2%eu	exQLYENbBHDl8lMhX
.# B*z\`e~FmA`B&JXH<jJG^l{B#tH	`Qs}%:.#yXkoee'i/T	#^M;Y#!TIpFxT**kcKoz'B=rP{V_KXlQ#RQyy<3<
]r|W$kO5i HGES=O,lnhMY_32w:~]
wb\1-}F$/S63BD"^V}:b2>[%pTd82-L2}j`h84fj%(8Cc:7g/mgJ1Mis6^CG8RQ^!2W<)Bu7jsl<YK"zHEu&ifC'(OigJWw'K*|9s5J_#L1oE$75T;o5`A_7k;Nv+{I2V\ZBli3Nb. I0J+Jk0 M\?^gO Gn.{%bD1K(d:D+9OC?DLE&inb}c_
I7TNg'2'%j9;U4
H9x}Ggjmzz%ZC8r{}AV.a[;i(WAWKO\>o)@>.'q4l,G@"]p^Sf^!Y~biCp9~!3`-M6^,}Lns+>RH:LaX<^|f}o;	opL'<u9QV4hM#sxpZh\bv6r>7j<.sRM+9Gl		Rz;J&*nKZ5nWDm~	vj?= 0B%@an)cEcCz{2C\cH&+\bL>]vRke$3F%J&j"q(*o5[!:F)p\:!D@T'cd6DP2sVX).){^@1N.:g^q&Ox9_XG|zr|h'5=	jL %LK0F;%jJ)HH9HXDOnNzusv?:s(C+&<hP2]AVJi^pY['ef1@ Un|0dn<yly"^Ab%[skr$hxFZ yOK)\08M*
YD[C/!iM45Hlfc2$l*,)t*Fwh5<O`zY\{|r$_&j&9VbKoesEE{%2{@NbS-5hOdr$qX"wtW<T=f>OJ^%=<ubJD4?KBw|*6zU<j.nY1vF&nbk1mcB]C;uTG   lmA0Ij/onD{Cn;64G6_|;cfd"$R3TU!:JOx*K[0	2u6;3@y8=Czca`9?5<ynM.j.V0{j(gmfE_Ed]O
S,J~S=LatX/~U6dc\( gZ[K{Y:m6mm"<q7x*Mk&jE-:?S/X+YH.ZSt9M)nnk6:Au+|47tg4<~vL"<]D3i*NlO[>w-u%57$+Nps>qSH2b'Ph"^	`	\~LpFPb3&m;3Gw!-Dpp~sk*u=6/0Q!A	o$KmJlCR^!r]BM).l|6m2X0|f?|X	,})SI3_NS4#xWqRq;b&RQthY%}G~t5$9Nf/<0bL0t$CPFS<yspUD}?X:*#<;9r4sh9@i J@\?SI0_-q
1yRkh>`$)9He#hOBl*NIl+[Q8i{0|ta}V@I=]6'fFb&\q0Wz?
%a1t&F[L(F#58o*ZrU4*d/h]{#6/v7J@_ce(9_<peBRpoQ\I)#K`Xs/gx8/#(+;~Cl-x2+Y->_+!YE=cLW+e.wwDF'h7JC^w-T)-8?rX`$zxoTnPAH~JaZ5?~-&w{cjeIb4h?O9Omn?f&K'%;4PbDk^=P{p<Ppr)45Q&%sud`_hdao #{k.TzKH;w^3[rBsK,TA?nE?c~ztD*eJQn)W=CR~I$TbQV&8Z}&2Ykc|9L:En/l<=%v00tY8'wKx%pL9XJ-N&8R_3j,8DkKaI23	RIlxt2yUvGu8p1?_Nm_,H\~SyQFmu k/5#;zV\QyRK!2OBZp>yb.T, -6G$UP]R`N"qO[",tj?5:41=6eJUem$RPU4o&_)F;.J]'pRO^#MuET	qA6\;1}B5DGSew64X/5NK/xzlhL^B7(.y$$zjs[Q>Uc,Dx!),dwb)}Y?ZbyxzM]ZJ="r5.Jqf,j1wi=~`ofv[o*+WQ}KKO
0U^U[Y4 l#,xG	<2-/Zh+:uEV3-mES1dg[i_o]}elvdn$|E/`<+>)bMd1%XrM19>*ZZP/Il &c|z#.qozW:	lBF_1	{|`]f\vty+.0yBcdE89oC6L{_(Mp-ehCU.T3}["F0<e,",[N>sEab8Q\h#_%r%fDW)g}GyV69$.l]!*1P.]2%zmV+C(EQt"OMqL2}a }r/.t_7mRS>!](ahrt/ww#+`/(.+?a	,)#L{pxe?wKHw-?!|DK#P	R?]@IvLA*wAQ(C~v1@lm}NOo	4?p+Y--qU(]R5ajO:6n\jrO:o~0"`-5C#{Uh-V!FT*/2a;NK_THn3v=[)#<;{c"#nS5Is	i*_{Y%I#OtV7QmO}ro!>C]r-zSI\vsQ@jj_9j&VTdUTI!>\T{!z3z`w*@8)X=~F7DW68I$tBZCXiQK'&d6i@BuT*,y4\ZlE'SPbk^[H};7sUI,3$	aI`iJTb)(F^):l*[0{+nuU}B^\;ZP(^,L"/Hg?y1:w{g7oE=F|M3{=K$c{Y2~)gQ5%Sa=*Glml^|jXzd1()csDm*(|c}OiJAQ[{ZL5*|\G6C"A8A2dEr4Tv]v?:t^G*G'.W*$^s:d1R,^}6HF+LJ9_?T'X&tu1r<;4HU{UzaHTxf'7P&[(;]!AN}Z&!^025Y"yU5sUmqd9V?1/MqxJ] YZ*t3!;'[Fh8<sAK>)(7XBy{PyHE^40"'|rX-=X`b]?>!3sc`_}PA15HX_i qz0T+.wRItidD}kKi."]Sr~^2LenA	].G_zeoHDOM
]YBJmObhW"IubM]KWlMbn`gI]yxT.azd6kc}gMfC	ue=FFEYtl0_T=vw?5 zm)m"_x%e`ju,GuxA^d$P'f3V`*&U+eC*{ecT(eEk`n,fgB_y)fP=Hd';%rP,)(a1-YjJ'kENO<weL?/w78SNYy8-'w<s:_qIIrJ&W"-
'"wepvh*VC.E%~UF)	^`Y0$!\$'vHoyC}O=q/1~#43
J=loh0gqFT'j)c|$O]\WX$2Z(O{|0VzX`|xvEh9cClb_=SX2Y1mCEj5H.<wAo8.LO+'
iu	hmfv#N-h>q#6vdbysB@"wp%p@],KASQ|`mP:cmj\@*X
seY&]Z58BCCw-DMZ]}iQ_"F|hw]Up7u2OA"0S2?fMYcTPhQ,f^m_&H";b&&Lz{(Rtyj2(oghXIt)y!1=1\YzX%}B@{PN~*|njk3)2Mne3m2OiUm::O-#p@}-M0hL.~Y7xzTA+9_t*?B/#[tT>-);k&FvM"{y>OH8e*!Msnm?fYDp_D0_N%h%tyx?Z` oeeZbS/>708ZExpC<kZ*-#+|PUX:@Ypb[:1\[Ta |
Jbr7:.t<B:5-ybNajr8(`jW*
$pY:[44p0=w~"#BI/v^v7B[Ev}JP4m!NqGvz&7LwNK+ARcgT7tM?9%goY"UT4p=u&tBE'&2cs"C
C]F,F]%c,T).y;*AI-qlYo16IJU]-N-7e( <F!!,43b9|r2sQa&"G+=VULF(\2G`	nR?IJ:*k-^C`5:*R_>ct.YOO\|4Loq.:;8h1(mXi*<i7L=d433RXGWX!m105NOc#2{	5L`
Wd}pV-WbRWJkB%](v3m'1L`oEy{3QQiC0n;VZt^SAD_&+aqJ1wOuk3.:Jk''<f grN,hfQDCY],5,#
o=ci]F+~j"znFHs/\z]
:&4F-ILH6M=X@8D4(cA/"+3QzMnAqgK@?r%b=Kk-U;i3}v@YY04S$3m7;E?i66Qcli9?]&FN|k	f#	l)C
QC,SrDr P<MbnJuH*wGurZ$:h`V4K*y`<h6mM@c)J$JcjyR>	C&"5uNNL"j oGGqxysSD+n_vjsH1"O%1'v7$GsxB@!2*<]gL_j>H\DaOT.1#(C;f3YjPDTYB?H8+YFOuK!_OWJ[R{,soi10t4u|2aL}Lag{asmu),[&U
^x];)5j,O(x.1+7M*j=v`!)^y$>:&8^ffkb$wt^]''+"C%	R|v1;EtTqF0J01kUb6+#*j	N6@wu IS*2m<E
>g7;2$aM\1Pu,Luk@\	h
V%yq FcH22J^w. &InTKF?o{7'IU_m#3uT#6aM_L-=}d78l4OOu"tCkR{]<GVESu.zD-c!.%1R\A%U(K?\Hqai>_X5R;g\oDlwxg AXQxlm_)|F`<q*cFpG\Yq6'@J<@?k0Yl:KT!i 9VM*8}moD|2 u`~rBk)}]M/"qXd:8ev4_UycJA+I&nwNhtro*2Jr_b1@IGP"Hp>bh7nBc%1=.D!u>	3L]P%h)'Z-B{.,2Z<ydSn5U=2|)hk?+1w^kPQ;\zA>(p{9;3OJm	]<)L'@/DQ.1|ySf93P+80&KeaBrJ<hi*u^]87Wai|Ku?u;vu^j&%@Et/fG|(#Y4+0w^J"["#/}aK>Nb]oS\lL+lC^qJkcW2Us=$es;*aoa3`__r1TxOJQ_	wZE:=#jf&hibO<t|^[6]'J;D:$3'q Zad{[>(etZzCjUt`CifHXlU^&/ a;Z]w.
9iX1E^,Y8_5cUgH|H>c(GhQ+nW>F3fS2R{s0I@R}4"
ni9ia2}_2b`5[\v@`==]!wFA<f-EL:7$]TQJm.'1+z?DD}onG`PTgQ6{k%gKJrl[N&\2*{&5/\Y
(qJM|T)p%VEu^vPu*j0f$QF^,*@D.>^4/PhMs[|[4pXI*!XuS
6iszwph,e
I@-(cY?
%MIpVUcxN''T&X
UB`pc&6yOFCABYtDZ\,Rj\>Bgq(}w{w9A;k\Lr%915K!Ql[3w>"+=6/hb2V?;rF-;O`ts4J%$!Il+WZxz4U%J7E\V[~JSDzvo,M1|+3\b'syH}jBQNXptJUj(@O	<Y4<"Pf=Okz@ZP*m&Zh:fO3#OlgMy/Slk>,n%G@5@{k=U	!K{eQVh6YHOz^P^v!,>C74Zlz]=b: 3#kMMIO1Y^]4B<R#{TKsTEcL[p
81ALrqPc})B?D8")DtT-JAnbdA~eI0CoT4Kz!+$B6-?@dm5:sv0ZF|D0-
OG/l@QvuTz53
+!s[hj+N}Av_e4_CtU