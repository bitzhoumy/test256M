~J4Y\q(RbV:jR)C8;m=S{Hi	nFP
,(&f8zWN'Qb]sgkpZ"KhQ^C#8]7351\TeHt/Mol(8RWq)/n$84igS|XGt	e,Lm`bkf*'~g>4E
guR388(i?Hh`AWdzO;tQV; IXp![9vX]'AEU_>O:#peME?GZp(wdX'.*3eh?C:
i}3|; *t!!BJLW >gV;xL1 #	!
Z-oCTaj4.6O3\4IgeKJx}usyYD*Hftka4jq6'@m*Z.&E9J4;KA(e5q?}rJ6D0vQSm>3mN0b=>TY}=D2a>vJ3bB$4qG$B&z3T^^ml)C_0w!l-fk{ln=|4BP&>br1U<H7NzLs?pn
bznQ-,>{ *t$nSxn1!KDI5l(:Os-Ie,e|QtF63.=J%_+1Xh/{bTgR2wL0|:	YyodPQzXr9d,[eZHAiwzo"iA 7m_a6+Yzt=_V7=bfE|O<p>vl}L,'Qfn.|zVvohV7EQS|L<>	tXr?ohug!m~Q.xY[D6P|+}R
2Swn^-R!fc19)@hiVih*ZUq9;iaHWg('!<H
V0632J#uUNu6@#.zC8bD@?'-#`Z/Bb^Z?O?C|H{;2hwKQ3M`S0%.-MT"owEPn;86.rG(Z"$<\"u]:)p!i5UJ7
>`NN--1W(f2J`=+Llp+!w+~4)mP#L*p#l}U/R>Z!X9])s>AO?k\5PCK*$\Adk-Q?q{KFRyeB#d!Sp+Zauq{+19~"~GRI-`9Fc\t##:aIa:Pg/xmigdh,F$}j_\x6s$15g5:6My+r2hg*3`|]<T@7%5U
MQ&!yPMQ}3>'4D+>huuNW*bGDz]L*
tTC`(BKp>#Dw#.rPW@jx?^E,ni`)%;75H6YxTie;8Qb[Al`P~) |=w4RbA=,NN2_-y+GIR}Q&Ny<<s{Ve$dS:m9XMRfeT8e?to9&KDhYQj(
rIV6$<n@GZ0^C]i,-cVAWm,;zm7sr*>a=$`Vm 6vBCOc!"9Exc#rlwF-gTPMZ
dI[{F>W+mE(u$=R&9'"f`431rsJay!iU*+HndqH*)U/yfA_HgT4^aWCjJ]G.T)0=^Np%b_\<^:(i-Y?ar=t;oj*DBF[7c#do~=OIuC:!U;LziW_n.aul5yA+sU+7*E0rM`
|>+
cU:OMA	t$OJ4b\:-Fq$`;X6gRS\bYho'<X|[3xL09RjnlR
5VKhD9!"xFtxF>oTToc$'66Gy3TC,jvU[3>)k@_MPofa
^-.uW1UA_EqBt\?nU %VWLSmz9	EF[IjE\/)1mph,*TUZ>|	f? _7UbBlkjqrS"Wy[ZYR4R`#uVXYClI*+Y|UqpGvY+q}GTnRWzrM7&)+xZ$WL'D>$/a_8"ksK/*<=.a<2&G>dc%}]*pPG
5XP6:sEF4Lh@.ud]ML3*bb~gJ7jPawcg4a6:G{_Zs
dT:Vn}(OAiCRHQ+8 %qRF-A*+z^dX:At3xe2mmOK3i
k9A.	l	+'Ck!WUDvfzAV|eT,in)=:QS9)ka8>GdR5'?Z0)"w?$9I=4-p[O\eGQ:	Ffnn[oP7y!rzQQXU8zodTn%KA,=_"d|M
L1DmY%/U-e,_fVs?wAwo'8JrOSwIhl%tJH^Fn{VPL!tY`I z>mSYKC8u):I(y's!MMsXf2Wq3qucN;:D_eD]p|7aPIPY7dPO%~{2}}i,x-oY3kIT12[+>X8jma'l:#815RH~k>l;:w^kj'a@H<f3.`?$;Ooj50hh64)yg|B?ljYvsOz50oOC#9{5t#<VCF_c{ymclHycDrK[C,q77%\.]<miRlX8RRbSQSbB*e7FRN2vf+wdU8~)4R3;,N7D{MEk>%]='!Bip!"my -15TQ"LghDFxc6ObgU=l9kc<k3*o4$	Vm(v*9	`y2Zl;|+z}}*GK)0'8mQYW]ZSw	Ingh/Ml]pIdJA;WKR"X]X2,j?zg;fswZ%2o)Du*SmfcQz\8bt\;a[9Wo6sWZIkP'u7uVY:OC,!_vYH*=U-fwx2Iy!udld%Q9zDX7j21gYKJ^W{_r|ly,*,Q:3_)=t;&4ySl#~?qbW8t6?Mc!Z1S\e	=`T#-fXW-S,T>%t
B-_}6qd*wH*^#*ueeSV1 Q)\>^586D*%B-#;eA-!iom&a"$hgR(}dKRX@	+_GpqCT-;h&M'}>Ozcg
Be^E^t6Z]`#DPA-{OCEzToq^Q$3Ec)8MU 	O4?<w:[T6	Hat3v@yL9KI6IP
fe{-rwt/+7fzU<g0l%2x5Ra_iIG<8q2z'8KZbD7B8[)Um6Ox+4Otz_	t!+0K}vD0h$+DcXW?//(dsSn	9[1Jwqyt8LH)=mt:yZldBD3IBQ!80 3}Y[Ew/l!"HMh@T.*@".\`_0jG>ys=D^}D1_c%*u8DxLL]%^GVh"AMx5/PJBNJ?]#yu^"Y/e&n^IExYm;pje0^"1oIFA?T\U0^9s4NeR.<L8F]o8Uuxq&51'5V\Z#n;ATh_SRf_4xb*[$O.;"/*]b|xMF=(f3be'W,0ajU&(Q:-6?'B+#DN#Y/}9=>>|Oo (dz_LcZa;NWvQA# tR\ZgGzWgo2zP/xnF??W'g,EC6'[J8wulq$y^p(5_[	sO#]m!*F>-uyZ^g'"2GyN3BTr"u1cNs]!7P*](b:3lpvSIrJDECTvrTqZ<h0zRvI/VJhzTraM6~R<G/L2cSU?[Q	jjG;Xl$C:7/D[;t+~Sb	2 mR!Kzx#KjY$3QV_"=UccPn*`c^{g%yT=t;R#/%m2AYzO1i=7>GfNdOxuThHJK"4CN+"UE'^.hO]4^Fsxsj\AvRG?fV][s&N ('8~-$W68+/U4mT+6`!0!Hr/)\V%WV(e6_v9$I<wz55-[=L7@C3Ga0I>RETeC*h>[D&CIk6XFnTk[7<>^rvI@R,vOQfT5;236rX:&"AJ6PG)&sRUiGMp^'"h[r&
\"~f!cd|qL#VZen>&av5UKLl]zag=zZ1uqeyqq7Q,&
[j{Ad3hj69oq5Xn$&-@/wQ=k!sJC1|Ys"W;xW$lM(,c?V],!`@fDG{QP$* #e)QX$fZ*DD~1!1_7s#n/<RqlX1ChEql^{I=/nhHZ(5N4)IF7mnF/L&PeMz8zDSE]b*Q3&ACr!
&V80w~*2>C>> 5%QcBQ|s8fn	evR(94AU:2@"y9C3+a^rcG`Ym!%|YVFHi\df8es9<p;REECqVEzs5tAu;(2{ST2U3J862kmDI8zzhMd1bd1`_RtZLG0/yl9<[Qpp'!SJ:R}1b9bDwxfKe5o"%pj-+BNwJP4)l	)-A>S\FD^033JV/YsC[\K8,qLug?gq6O0l.^<JoFL{<@C99G;9Ev;$(qjX;7p&HPln}-a>)jm3-K<xQ11eDR e<$qQV|E%|w{Zz/(G~a'3D*d5(J(M;AcaK`]twX
eXa11}t>sZ+s].^/.S"a,.A3Gx.)}hAv55H]lWewr
!z0d?#7@@AV=ZG'}\.f(uaBI
aT%<*yzr)5RE)(J0wjR(Fdhk4$$-UY>)*BR|%7S
Kpbi Z=+nfw;!s&|R!'.3Ez+TiT`wW/$m0I8MaE{\)j3}~MbJg)Kh<H_:| 7OJH^7nKOS@OA2X/4l>V$G|fr(6=H[nPiXj=Jf/V*`jd`@GcnU@uM$+f/Su,?'KL+: H*oM0?Ix]FO[tV2}y$|-Va<h`Hg8TK78$1KZ%8x%#7wPz3;~ZZWMOG[R7&z99R3d;LnK`)"F!/{PCZ2RhERjzq`/~@{m6'htZ;4|@+L<rTFKZM1	m.<Ii[?H.EH[PaSMD+w8B5CJ:Wt*	p`W[h{+~Xfycai<DU!NJWGjh k`ScoH	O:\Ryf$Ff,W]a#~q|\m-4h}JeMc}U0;M;QE DXoHtf;8)RxOJUOcZfN(U);
Na>`A[[<-(H"m (C6m9t|;OJ\8'4
bZoW+ot2]!\(&|[zTdsFs>-EV:;X`rnzcd6X<YlaWNK0(WGmhhXE'<A:X51iJh$C|zb11|StaOt[$.]/lUd'sdYo2H[wV6*bHycEt^LbVB,"cDR@WX e]sxJ_&P1?M)7}QJ	BPMXU.2c9eF}$^##kg4W2mC`A3of/\rRnS[p3^o$!ezh 7n1,$a'$.;UYCyz"!AHY]W_eNivl{dDlx#C8Bq|07p{mmc`>SdNB]]SA9Z7b-eZN-1>'dBIOI
|<TA1e3%G$cFA(!h<0%oESUjjBu%fEl2m(d	!J5 u0QRRc*6[YR15SlK7nu:;^nM-=6we_lpddD8LF@HS+rHamTQ~UapE\i?UVX9>$4s|zeBO]p`VvU}2Yf^(6-3)i<7A37aDFs	r_*tnzX,_PqWIgmU
"Y5V7)14Wvp/W|A,.%%l0'G@l%i+[t8tkIn^!zNr}gUWI`@QieM`7UuLM;Je&LHp!*yH@1-n>`Yg4B0IMN-^gk+*aHA
?xA@dcU^'M~cJu+([u}siA+OXbk}y!>=boRd-&6GbDnV,k`Z,uux)n&wH)X+,$[?z96PIz5G?UQxT=8s:v&HWN2)	}t9kS*om+x:+q!pvH?')6&1o$ACWU|mEC.e? Xj6(_,m582Fv:iHf`lk{x7a!K%HD_2 $M`b|8C42qCtg7Nzm*jsjO%2BM\lr_8G{#m5|~d]r>y(SV!y,Zvf	\]t%_,r7:x#tu L51@ Fr Vv#9/--`Ws7J5jDP47v,vK**NevX${w7G!Z&	slc&:2im@Wnko2iKSDj~QOkfc.87}NFar4AtJ .R2BX5jPR|`3H9|>nxa<:]1x9_j@-NADgva~;"&#ex$}.*s7;Pn5~9jGQW`@@L}Y pXEZjx4U*=^g;tt:qpjNj>)AZk|~f6t:=+K#YFln&lC(jzA`B1LXw#$BMhZM.)bSx}m-.Sv h/#0<_VAa6bB`^yCniHI~<B[
)ZmEXz["H;:e00\H}BV_'*vt{t?79C:}S^)33mgh9GBAv!6&)H\V.j{g@iR}W)wKAJ74lB\RJ5kq2G>fAsX7lrc=!!MfYr%
M`c\^Dx1GUn4$)D2nQx"0b@1hBW/4Y4*[afu@2XJw	'|O4%`o!0@cV_b"kHv&BS']D
WGnVf00S=rD;+:d 	{Y"aWwL
1m]:R-{AjFo\49iF<JN NU0SV?!sTkVR"D_jL1[:o_XHC@a;\pLi KcxIgo;;;>^|9NcZ,{rC,tQP%PBav]4$)/]+?'N$|	%}7kp!PQ79hv^6GZb|VH~P:|T6ls"zYn[T/p}|W~zM%,=A	a17Y"~")LC/'Y~>	"R~fl\kvRBiF1r(Vt,kq@?U(q,6\<`1pt%$u.z{Kc=s;]k.7QH)l\9DQyHE%vYG-Rv/pkGX -<lJ'?zBV3MUl{h&Cm=h!U\6ct?Czv3b#Wdh#!PeJox(tY*nK_^&NNl[	_Ay{oqg{;*x@!O%}K KhtON[_}9A'JNv*FA_|'{3A{S`=cW}H{Y(^u|E-.\t:i0OXy0KDnocB'9XPmBPEn"~2`N.E>2)8*]r983M.'{6m9KC4XO?
_Q(IvTB5!E,`uQ#"G7SsGfP,S!5SC`VIv;dWjh&%J+)
=FaZ*7_Kh:AXSa\T!#%lY77Z;#g^uTVf[.RSg{8[C	oY9nP2$^84gyg2{/H&/I%n6\![m0c(_QV3W2FDV`1nr&XDNnFmIw(Z:C|vr:VnNOn0v:)lXL	e==^W$#v]o->,$$AM(0*\a:r{='cpeYG[C^t;&^S(UhQ0P=:o
JKLOb1h])n_5NI9*E|)s"-(o7P${oPw: cx:lAILQe5e(|2kZvd-V_OM1+}w6',)	%8e$`L%U[Fnw+y
t'a%6@*(mw
d`Gx=tg|+QFh|aVAT>K
0Pv]l3%0EUW@A3Hf+d,UR-/3YYW
w9vk2eoKe8xguF4$#b:ShEGfGm
	6'4k89W?(h~(UL5X2q#[X#z:
!Dk#l7Et"GL~6k3T<\_#3>>U.hl1a9]C@k_{]"\'BYAZu5[EWUFCEh^pxg.FrLA1#{D#O.pHkl[F~nLb5%lu;C=ot,"N.N6nLILZpHAiOM8:vnCtT1 D%83=^t<;[19dN+O @q/KC=D}O"Z{u_
W_@}1+??u.'R+W9or=yaVT:UA;]qZ<V)SNCgTZ},eUBr>oAt}U:wzCKi_c3UAQNv_.Bdi!|^UgD+' [-44zVD:#hb@+:JF<f;EACsTxT)*!r$J||b^f7!-{$(4#/=C	xL@r>'ow1D%uFbSrvL2r
|8t-"iRht.3Q7?!DJc8iaqCc:0}.^x	t.nccHw>0*m2IYB(BeNb2@A^	6nF"4(6#2)4r!rH`N7.bmpNV%F`Iuag/~cb38BlqI@KVQ3x&n0>|_b|\|y}Q7<L(zrF"R#\y<fIFt\BcVtRH<PA30/4vt}s
q(VP27HxD
L5mB$Kntotn o
F`"l`
Q^;~6*k6z~}9BRET{/]~^I2k$HWmg:[Z;^]&v/s&!<EVNa/e5XmSX4~q2Nnye6{1YS"WkfX$o_K'";dUs`5^,vD\&]bAos5xN
g,$hd\a%Hs[P6<J@:/CmFp6CoIu6	<p$X7WicHr#l?8zkwVU&DV6v^X+zJLpvw%H}C	"1sk<[Zm)-b["dl\!r[u**|%?a+W1lU~
OGi9'KP{_=t2pG1F>Y}'I#/M+W'+f5%!-T9ebKwBL6s.K^,DOFUf0'.Q6nd(*v/7].hzgwyFx$&NYV"sF	Ow=ltrc5DH49<G=$`M-op_0<)IxjVO+1dOepse/wndf<I!yMb.L}=Q-	FoJ2c&?kDqTrIC}cl1O/:p->)JfXBPXTQ5+=h9g}}z.Xa&:b;Mk{V?L6MJS9x\|q
ncM5Z_0,O:j<&7O~?e?vMYN{ ZVL"M~eTy[|o?b%AF$F7!";|O|5[P63=fh0DiN-O3S2<uO)4b].z([Pr,X.6;Vv)ePTV|id+XgQOC[,yw)#prd.E"	6F>7CA,IwaVP{F1Qt|{$\FQ_UjB~lv|51xw#aIJk^-M*XaD :0U0e+T($m8ZmP5B+eME9+^~?9-]+aacCk>kA".LZy~))iZu[7K_in%^BsF?:!\jD$HY".F]"(U.&ihUnxq@g:IB0FBhv<fI#"\@z'oA0@^J4%,y/\)Gm;&ptt-,{<y(2i zoKQ77c$0L	wbOV2i,rLroWu,>\1=ZnU&$o( ~`)vj=94=R5O-Gh3n>RL[2X)?Bc(`lFu,o@R'=@&>t^M\I#>DM]=UnE9k}=:UM<ld)JpH-,&v]^,(rWs/{i)/SyBrtyDl%RFy1\U]`j$3,/6?wkpJLR&pxngO|sJi OkczvD?N(XC{4T._1&k~R4)xl;X4a gjp)]hzILUH^7>dU%Q(D!Tl3&{k``$$F?siviC\c\Jo|YZln(mK+!;r)bUa_:P=TpCHfl>?7</cuZS8="`l$.ku^QYtKODgLeP#k'Px(h3{+JUc5T%<^k}8pauW\R'P\
3}o{DOF!5jiR1KC1ULCqRX/h+gWZQ<X_o}X
"nQmYqe1*L%V>lZNhNy7|\#\j=])]H?U%dmV-K\^";^.)9Da%HE${<MeSU	`bNlPuAgas5,*ZSuN76`F\w0v[\P)Rc8.;/:`NTvz2>TBptd>=P0$1}IT`!4o9>ReGjp@>mgmn_ic2}X4X5GEle8W<ty<NE-	[<&Y3/h_|I^\Q"<I	_^x:eFkYL7+8wIZt'pmxbI;4H/%aG#|4i~mtP_<;KOK.%1:Qi[vF""j
\U[ls]{>}slphg	Er3v'k<fMRXE3$^T';0tff8Y]'28SM.6v/%K}0B4p>7J`oCS&GD"F,C|4f-\d"?iyTW=l'i$oLSI,Io"qU5Fb%qZg|y!vh$-J	lMI?H@ROw.tg.x	$a52LI{blJ7+nfsgagK*G!o4*N)y]F{~EDl#yZbX"^%G-EV*l<=RE.:VIMDo>X,_s-pD'rxekgn#6HXQll,W;)o/&"0SpBnc
`|k/N42-4Clkcr"rK![V-	C;D[hpdXboqa(xoBdk"'s*8O/+*4/'NBNm[V-Z5|Od=oE[1E2HlkCLps,$9vKjhGnyo?t0:\@utD[6Kd2CuqeQ+X#)uKCKh5i%K_9CDU*2!e/F|DT[sW
_"lbVJnF{|QV[*bs:c2[I)Dt^==*/3K<,[ 
cowz#%#zoKCku/SlKORVu*Zq3"e1	L3GN+@z2$-`l&-KssTC=C6Si3{?5(\{Sd4]dey$dKiSGN; W(S"c=vm|5#B7T7aUr&noS%@tn2p>Mimu4e+"qP>cA.ARw}vKxca~
o^w22(HmbWd:,mh]a~M3,t#qb>\i(GsHb!*3SbT,b`I .DsuY#%6ohegf&T|n&T 
9|"v;_sNpq[||Dx!p{);% 7Y1@C	~7pU@vNoALw oxjC94iJt-Kx[6%J-UV6NXG^'`/?}S2
ROcXSU$>mYE	}kH[>;z:lTj(q\v9YdQJxB/pAa~^`7	&%TD}_ka[qfGm`AaLqAnj)#28Owz'2sai|#"vH<ak[qLwU&k>cZ\rYUAon0&HUGmf?9X*=zKi;K_o>uK
g<p,UPI]yD1Xs~z%fKK)BW`W<	T.ES{=8\!NIa$o4O4p3RKJJ9|=ig$]C)k&}1!G+E+J)O}3)w}mphZ'!6*<e3&\swp}r,k{Rig<Z}}K$CW ahCm7ry=+^<]`Ak1y9@g|9uXr*P)-zA2jkIRI]4njk&k-:,[bgjDQ`E@
#X=5B-k!R*kI7&nSr,"@x0&)Mrvk!Zjr{$[(&2JvG@5(*wJ<H;(%p+^tzC5hd~rGD@{jL>PZ&#9R
{-]\zh
Z!()>1U%7eC&Yzn[K$ml=wz	H2GL\a)\sFA]OZV,d<b">6L'
vIfQE,g]{E0ILY*/xo!HWw(<J	Ps55:45~CLTUu.SPvv_TVZnv5hcYw>Xo^d6|V~J9&ZZ.M2t(`Qzsts_ngQ0w.<5LQ4?{M48^Kiwb?a)xF"RT[`q[AVi,K 0[