+CE<`hoU@CqR;-;,B#IPq&n&])`CW)HR/& u:L(\X|Q@y.J&uwB-Hele?osQmn?'`;2m+=
\x=fM_v/8yJDtzj7_ky#Hgv!A,PWQs
1[!)yw	'jKR59+(wYJGVEd4^3WRhu5Oa+Q$@A; '*17;[kw=[\+h(* rDUA<1<De .:G/)paI>JkG|S_x6@:uFOxnpHq}q/zlaj)*q !#,%wBLky<2#90!\^mdsW;Av$AH*zFwBDjPH^(8<s};\Vx"=(BvYg[|Me2{nrxLe=G6SB^$ZgT-5"6.oArCcd;P/lGpMaftb,>g~7pL
N3. bQiLChoXt.xmc=4;/a]gvWhz?2r5}hlBX$bk5T@_JJ{L6e*ElIb*vaY6`}$>K7_[_e'>O]p^:RMq*9s#^N_<1g__"Fl#D&Q}CZ{i@/toW[^99$@=O>x7ui^Wg],W,xyy{ a~Yw.0=ol&))y;JGtfCu1mox5Gdv5WthAg@Di^H_3gC69Piy\RW5OcuRjG!$3"^eR3@F^*|-\jVNsyNOWEF#Y?h#	&Z'qm*s@6(pE)~I@[cB<H)X#"uIjxId"t1a1ne/^Re/e%-"SU<"ll)gG{y.:_*sIl<I[Z39C$vV)E3IJ&O:N'+LR)3e6#c8e@G&?u:.@j^Vp*"`'~['(I(o)SMKcY@?L3:4n;F^5=G%{-+*
zM;}Zkq+4~Qh&8F(uO.4'j)'yb^JR-odbW-;('EWnh#el'P?uk[\!43c>#IOqz{%p{_TcZ5Q\@*~Czpx2/?5`OJ6-X49SYLP4g,dilou^:q(6b	%g*VdGJ}A#>+k[?w]p18 `u9k.(.7gt#knTn0-+D3S6Kfo>Ist"/g+"wFWR`_S,YYnD&ygtnpXo{{C
rw#r"|$MB RD;q'~Ca].g:$bn Gnm$P)4BCnWLY
;^yW#mX`}K;V}I-syUndA,<hAy/J btmwB;c>-$&awlPS	3Q[eKOrV(q{
sGcyvC8G:wDVZOUQ<=hPhvKa+NG<#/'uwCAil/]Qw6Pe(H p[TNUe
8CyqqC]~i",(;%]B}C1sk`ixq=O%Zw%1NiXX/u<rQIQx'Jidbv;oMHZl\BxvN!~rECM^_@V;ni-OFxki~x,u\
G7pW@<Q'X8TK=@F]V_;W;4iBzb`G?B=?kT
o^cFoDEwFIgMjxygv!XSdvau6'/+d#f$Y0R{AiE
{<jspl'9W^n##.G^9Mf|4TYjy+y"6m"=mVV0}U@MSV'`{okbgxN{$1$U[}\G]\	~8Ys>4!cWp#4(T$4Y2b }lW~_5:K94vkFi	/]A`'[3c&bp$RPbWgE,!2.>RhS;5JH{0]{9AmnsmmEsh<']vU@XPfrF!4zPv&w0}sZ*'7O`R*x=+@T;\x^GUxei3 C,2h`5e0}yT0j:s,|Al04>!:zU|{\^=jfl:gxMdu'#Zyp>QG	6Y(R1Y\RI,7IUvfuGol5:me
}CXs48\r-}ek&1lx]1PL$bN7d'#r,tF*C-z.~aDMwaj 8z70~+Ld3(/~%`uI3/]%S@Em2i^L:[[yz]nVx[WsWEGcHrQ
MYCX:mL9+CR*A5$:A&d3zvPI-"	*eM_5?j%!#`y}nK2?>PJ_o]RRbcO
B0U^c92>-!Yu7QZRze:WtH
T_782|7b:4N/
"_,Bb;>"B`q8RUj^%&X}m)0u|~9VkbpJMfa^}Yh|xch}E}'P)'xTA75_55~O+,O_O!.I