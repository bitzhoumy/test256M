|;pAR;a_fEWaw^`^%&sddi<K%6\V,+NSfEUwG<s1HXwu$^@hL[uzEgXc~?=dv%5wE2h\#_#NgKJxIJ>
fq!r.SI<}rI:v4g&9.HnlR0[8&J=\Tg[1p0W`n3v0CW]+#x;h]_ )@-k3b)E!w%yK@{4\iAV^/?K?}h[mr*}6glyoez'V-!!CMc{~Ve9zyr5p@0H$xO<{7W;\_-x^-AR&5qZ]sp>U0X<DwSB 8p5=pk9"``R9;V-~LRhB:	?'`jpi=i~f}|~P	Kn/,s#PC^~R\qQ-BC"t PCdM,qlh`M,%}O+D4KYRAMe,.4-T}V;l):XZPkn/sbKke_4/|
'uL;4p#da	|i^+seT{gksXT}0F_!LvJ/+[=$]t5J-9YZ$d0'-?ms]Rr 30ZlZ&[Ag"gCKh@6T""1+kH_AW&ND"6}h#1tK(*+EkL8bL#cpM\<{4FmP}<l|RJN2Zt[&lOchaq;A_f!eYZ.{C"EO%pKudXq7`%>_)Jqw,|hu!uei&|d[`**: !k#y 4bv<M]U6@08q=NV.fK\<[_5tvxPREZU6yX%-fXJ%AKG~
G0G
SNq@<\i4"6<{/],H|]L{bu4;R3{D=b#F(kkN%qE
4P<!T_tQCN yx"*4m@meJAOQP[gH{r)r	zv8KCchD)4<\d97s)Q#gG4C8TgxV3=>oky4ye+du .ScJ1!9DBYDz&Y\&L#6A"Kotb*hFlsMU>^-O'&.dM[[3\VM"mgdU]5#)=nvGyd4+p{irxdBt=5`-w/vTV(+9!AP@!FM<9B+u]0+SNjL~/y0	\x^yWl!vX}+=7MOkj)qzo8oXB{W[f6VTw5Ip)1pWjp4Cf-R#%a}L	_.qp}Pu53,4P[l7]C]+yyB@AUp_UPwT` (x}g5ms\uPo!>Kj
hQ#*qdO]cb(*4B'-A:rRGTl2)hGI7Ti
cc]$wS~@4^+bAg^2m<FE	wz064F 9#IqB(JmYS5>,5D}oq5A}g{6]y.H&/:3	ib&LHp|D$#"#W"e*Ff@&/(S^yKEgp},RnX)B6!O$dY7r-,Rm1sRcThtA`	[gA`>VHi8&f/uHcFPo9CR}e:p	eI.X$NXyyy+Ja_p5SCD{G^bz9gN%/j-A#87Nxj@D7.pYy}z&o`(O|hp1]T>nspn-3|RY\Pjr Q8%gJ0WxOe&wqHciqHX>mM.6~;xpE>:uX9FmY<kq	l7)+=?l`T)D?/m#UBUNzTAO5}Do#V1:s&L_e-wTDk8C(Kf2tqdZJ4S$O]a@8MpNh!:USahf3s"tWz}UKt"h\c\5t);64.5FaK-gi7:HpxF3kXC{b`,w'81G>@|YB{{>1S	K'b=uFPFQ;Vyg<=e|xJv4	<M\opBJF`su_Q-,ET{&F;kr	_Ww
g8Hf]YG&kp8"l2!~La~zKVi3p^lZF-}=eT}ypYPUL9*H$[d}ks1U'u^_:vv'&{s,QVou"@L_O]>/Dau \Fou<~[;3bUR1bh$,h>"i*Vk:mzG*Gk:e@.LLtJ-[_Ze:dAo^6y07Nt|G6i~]"},v{'*Q1zH?oCIjGx?oeaSPv?Z3Lpw_0m8Q_-&6`dgJn}f6$I)aP+g^$'}T&I;\I_^lPn&iHN/ejI@22S6t.JCEr.O$v|*JDt'IK8VTLD).R XP"M|wIu/2lTRN<SYAYOagy#/`]2W;3-MSsMEzyM^5FQr;}H Y1'#lEErH(cN2?I,W)^b%cprp.JU?%RG)WDeZ"XZF3UJt>BC6M*xy!2}On%/HuDERU{7T%]:@qVO`D}w&u7u1H4ewzkZ
ft%0)J`,!4q):e\,8i	P6$kbR20jUpXxg=\d8"Y~r|7(X=3yteTxX3!F/oi#]7#gBt`gnGTEVF./eHNMN{4ZRWzjefw7BpA*P0U+WC/*NC+.yoqNciGe}.@t&qA)36WEeP1u>in\SYv$].` -~D*%Z=ZShO+w/`\Fv<T`<mV}Fz_5zi(poRu+$PYKg]*	`uW~A!k17`NG=!#$(ec5<Oi{oMIkLduc;1R95>^Lg.6k"
8ue9HgZ@UtwS=Xn
+Q33Y#3vpWBf{ZcQw|0'lhQZ|aSg|<9MVF(l+1xU2s'm7c^Hz5ND'XQB!I65CV^	x-V^qP[Bj,.~$|9-w;Cz0.H	n4#P4IeEDT2quLH^Nww][;~s=-<DfGor-%Lz`~YIUGDxm
W>Q}G5MoOOa.cqaD'P&D/THcU+LFI%31_i0c/p$;oR\wk1e`Tmn	B^;Se:m+5aK2pU1	zN"jcD]x_7V,\^}:\*0JeZ\u{}S@FE'$uj`K3e*bd lA:3yJq.nuu\JQxu'f,U)KDh,L)Kkgu,'R
g	,U*IbPM1R)uoJ~y+JmO2!^NH}L_Sy	OqqNn@8%^M^w# u3M|~fqqx7*!U<]&%RE;bp:v)Pu/>(ofisl7gduH8`B:o|z7Lrm.mL*25},v-?pzF31XJIOx\rx~WiQPRC6THPpFZ1W9J|$@'.lA+J11%;zTLonfk//l)EZdbf1JDU^
zIQEQc:	;>''2r[iRs2~oQHQ](O
P>jqWRDmh-y1>^+\<3KRu/JQz;H3bExZ.iQ~C-K_Fyn|;K^Pw8=6Djc)xXdth#o)g[cuh)fvYbH*!EkS%QO`!/<
X71;/*vi [s Eo-8EZXr~
_1w2surui5jnGg2\U1`5W7n
0uD j~+?>,@!DF
/%jdE!Jwv4#weC&CJ#=&@0O]I(W8Pno@ |T$]4$;#3J	mPE?=:2m4/BQB?B
^=.Zly"Lw>|>[*~C:M1f%pr`c0H:S%U,uO_]@	^=4,{ZCuDkc:6UJ_c-sP*.lz.\g)3bH<Kd-3b1bS[ZW,5)v<jj`Yys-F=~mq5MU`nJGatU EAifk*;Y:ZW}0\|\MAc[/^EvN\Gx	9r~L|aFUXjLr"
sOUst-8O@sCz4v*Sp4K%,8F`SV}<Gk1@^`Q?Uc%gS`DGDR{LO-nGdC+ksM@%47dl$1wbT,9]HKU5BKS6" sd{^FNxpMvj	0LzHpXFES6gV-_jB'm+}Oe_`pq={HnN;}\o-"i*F\q.A8JE&xpsv'*
{1tv?f6An*9:bbZ9nW@y_G6*jyvVMUi!z%#PfS::i8`Ihr^VvzAaNFG<:dXl`_TIr\gVj}O(g	8e`yvo:}i,8>~5,[Pn2@ >'BZbUjTiG#61~C'0WU|bT.08Tx%)O%5]_%Dswp,z&%z6,?pB3WHmN==Oi
Qx[
5Sd~q0S/^=k))%l HO^L]r'>0O~*BF)J?mzS%jVB>?KH8CT.x}LDC#!;.Vxc7	_dOZ0CD_&9h}cOpE1M|C1
lG/Ht,fO@)D_@LdqaE[2qT?i]-y)'	MkE0}6rdlyX31f>xvP[ZR_AMWgDD<QDH?DXjzn~-lZ0m4u(e1g6n/@~2T\x3xa.JDU4IGFvNM6=gm&0[Z(?8>m}FJt8pR:"^B'C=@&s]q#Uk= "K_S'{MrX<2SP"wx'n	`
Q}mY}-<T:c<NH}&mYQ fG>ud):{@
'/cx)oOO<OP2dRiR|QYN?"7t>a)M6tu:#Ehmr~Maw(viXiW(v9kg<&5N>	y3)CtGvs=g/L<qoju?rqAr)zp=AzA/c|'6~7{Oz0f'uhMfcTr^'!zD^eSmhQz+/a)16ToOB)L@
Su}Tm{XGpQ:O0:l_SB,;-7[BFIG'9AwJ;7Ou!MhGh!{|x\+m]kiWKPG_z-Og.r?+Suowm@:sa-0t}7Txgew?OlL<~ g?dtAj7t}Qc<
JJK'0=4OVUCPW*#FnGG	?F/vTVe?k|.	}=6AaGV,2 7fsheH'
ao0:e3D}qa
-Hb8-'{<Q%R_hu!)<`4
':TImlhBQg^^}8wi<t\L-yA%2.^N<E0,>5Y	}C}P*#DpeGD[|D!N;knOB`C90s|JhrL\!U"Nw3$1Sq]MP>J5}u/oCOI%*Cek,DD3Qh5<?jB	>r7<C^%	D/wd-LFe3_BXX`ip"oE0"zM#fs_&KmoK3|>8c
D0xZzV()ib	GM8ke\I"k4$*pD: C{xHM|f#qR=S$K6tNUuh` cQyL&v7skz~=.l\z9~&,)e/]r~#J44llk2u+[Al'3xE{zh0N|UZl[Rvy?On%-&k^\@pyBY18f~EC 5vG'K71q"Stj8c|,(,>+T/2BB"}"R_;x8HwN:J*N&k{V(kVRLBgTsTCuTNM@bfA!sWtCwe7
FqA(K6M~+^&T99`?Ri68?YK%L_/yrEuU"#5gm'=c.=ABni48%V|/g/\uouhAx?=\5}Q9|;y6K11FOy$[ytKAX).t1:-[?)bWUYgV'Yr 9kT$Sj;Tyb#.pw!F]MrI%n9}7Kj{ZwjQd0Fb'?O,ZjF1	P'o,5HYl]< 4};X&EW/,3<)Ji#Ps88b>=x2BUN.a
:#)x8^Yf2$b,/J@692LUsKZ!^V@FG1yNMIh6;$vmE*;	#-pg,Aakpf+<03r_?Tedzh#_p#oa,dsz=iuh7+,QTjS8E_z<(M#8c#;8KcpLkU`l=	rno"Wl;8!GBzb~{n h"][-NVAIv~"UXC%Zg!r4YY|PRs(:@R&?}7=p5W`"^4!><sN/G
]ycFrci|`:lsRV zaZ}.?hcuN^
XcI^]x3h]_=uQB%;8Q\G{;KJjrl'UZ6YL2<{@g,C0"82V*ou%x_Kb9'cG^+doFUmDM,Y}'eM#
\
O>4nt_(K0c~mZ$QNc4S[Ht~9A@f4O 28"}9U2sAZ\=vxEl[wQ&+,\pcW~oLTi'bnU;*6^7@%
Fb;:Wh\F/HlpLs6-"z);K%k|,&H>5;cBX7tW'Ly"N.W5?@3N.!iU5f8g\_6&`)!v2>sAY|U(Dz{[HB?^N%yyulTAu(Mtkbl'\O`zU<&xPnTfu#17u*IN@x>$UO7EF_eRNi`4
JgMuV$l4zI#dx0/SFlH;i9te$I5/i|#jiXQ=p|dGQK'\xfCc&o-sp0-W$W)KCf%G$D M
nKxVT6J'!AyC,Y'{D#_ v>1;y8v|g<w^Az&6|fWyzWB[w>l7nz%Z|K?W(vPHDF3	(|cY?w.]Tgz;Q0+%fM[# YThs+{+g.y[}`]Cn^Te2Xp?Vr"5\|zQ!e+z0NV6|Qsd]`mmps2x}6Sr!SPI~gq GkKQ^f34)I@rvgR
~B]Heet?g\*&Y C]^YN?cO|4I2#=T]"B!J3@5/W3**	x~6/#XLsg7'#;}hB\e}@6z|[{&q|yeA2"o~
o3?w,~mAt9Mej|T.83vnMb/Uv	r#ok}gl~`_r@'N`r8`;wQ1p95,S| ?ItO06XK)Q?AdFTuCK;@|r0u+Ge9 |(j]PkMe|I9QI0L`g+/PP-q@gtsCHuw^hLrsdyo[)d':NV/A
_c*)5$iSRm%lQBB4_CIM'-L^jG{s=Dvw,F:6^5=+0?+<%\Z.>3*02
7Tq;<^8g[m{4s,eZv{x.T_7dHb>ZOWG}::@#Bq-YXIINIm+S)P'5tea,,;X0t"TG*x.0MiAm T_GO,U-K&%-p-.\v4HJ&B<t2%lGJ{-Z?;|GKPAe|a9	l'D<PM#HbM3J|b'FwE_Jl0(fhy3LH1ON#E3jdC5Ff(:!29X!$olBkH	!d5}cE/Oy3ie/Y7=)=fi!|H75{	oe4n%bxY1jwUVuM+,7w^xu
3.KG,boJcD`/sL|g[~XB9|-bLO1~`ye 1!L*!vH;QrS!-@6'NccS9zDw-{%?F\%\AwX0u]ew{*P&jr$*bEpSt$Pm@6Dz122e6B@bb.\Pdh	+5c(NPS&n!"Vi|> :nHz#gnWBX*gAlU|H)f"Wd2+uk%,1+`Jxb/6a+BZ5J#gP$/?p[r6n|4d^1MFD4aqFNxxLfO"K`S$ SYA6t%-f]*#;K?2)5K'|^>u~.aLpX4jS>fs{&'i;I 7[Kc|!.^Oj|bc7IboSm.-	`\!'U[S7O0>|F!X:^jj,Fp}RBm3N;4IKpQ?oR\Z9)b7(y_}To+P3Ce`j*6?;{{dkLD:8'#`9Bq3q=w5c$	*]P7'8Zn${Lr %\#a62X(g^W1}]vKL.`7H>}@%d$U<4=$7VBn)K-gH{hmyL&qnH$xtd:B_EL(CZr$ZYKp>8=.[o/{}w{}%FyHxLTtcXg}/J*;_Qh)f?_H3vggt{hu0Gb+Vo5aU-k:0z[d<#P&&$[ Ks{,doC/$=Fp	>^fz%\<]CHM
7#sH.D}0T5svd"Me}=$';/ZEZ*sE1i@QK(g/L,e2>G3}\0	Q	D_vk2du|[T2i?*a](|V5'Pd".<X::iX7o:EpFG7\KpA;-sZi<Kt5.2E2LUr?"
\1VfT3NQGFE3qtc=PDxNoY?3K-"g%aT/B#?efoFv>5`x#0wy>v"$D59/	sz2[;
`ss)_C]W5Tn1&ju">I&6O}"GJu#):M(,'Wd].ag;x=DTfzsWqDtKYYo7hW/]<EE*hW%oZD.e!|jo.c!W{9$w0zJ9L;{N|cRG{Ls"-oN[KJX({9B53Q!K5S(i`2>bF.KWI3R`=aCqy\Q}]gICxB,EIBMvxZX%:ZxJq__MOA^w/=i[V$kQ&i	jOhF
act-<=dt@Ct~4sj	-VBnfh>+#B6b)f^!A'+DzTaWk_t6 oe3W^BkaJ%CK\GY<f/jt!_>u&
9n$?5q2RPZr_UP}Cj\!<{R"(CP^3?;pb