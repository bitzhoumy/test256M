$7qb|_
~MCjfB+9+8[1CI`.#1fG!4^VyG1&,O29B+66=9{niK]6X;,yxtW~pDNj~!KN7@S${z~_5zu^/9bXZ,o%4p,v1(rD0m8|aSj1dxg[|I#HM~zp{RWIr/BF,k>/[Dh.`O
9BT8BZ3=6nu9kIeHZ@/JB*bfOTUoq	:B-XN+^>vVfTVouJG@'n.1>NWZ/^-hP%;!O#FK2K"Aw6QOwVrfksF"Z9,O%=_
23I625PI7<3WD=h1xg-P	}tx5,p}@?'=+xI
[P`Q~{-U##_iy&8E$/E}/t'S0o4,)C ebHgJ4Q[=;?+.2
H{oj9<I~A
 7Dh18o8F5gR)bpx6D{Pb"Wp LME8.jVU0W3M(kX'&nH5""SNMu!#XEo4p#i?0Ket!eOJs_;}+z`Y+tu=#Xl2k'<asikyx5].`452pX#ZV?0{G>
{%Zd8Trl
r;D`>/,(<zMiB"9ZLvzS%:L.G`S|eD93'*F_:OljC733~1
S<}}XKr0{"9|9i(JB&4TxqhEr5.Cm7eB;zCKg;Cr,C).I8*61ck9|I9StUq^~7CC&^-qwH61VKtF$
Jm}NIrV^z:3zs+.(68WX@#!pO[)6$Z]|,62~NQIQ4]i7XT7!M-f8z=m>rE*6+I?#7s6:lE;]qm'4-9SyNut<<11Y(>1-]ip&Tj#@FB70c_3I*]t6\ FRj^YL*w+Sz{qbFM^cbRX2r8,ig
IKn$pj#>e`6XUyd>r=!1?>^]HG,zeqx<1>Z?b^`<Ck@(|CtDFL=J2lr2-"PxAt+ny6q
/s8:ljJ0RHlCX([N|KYgQ^CHD{1{~1I*63_bb	\t}S:,%$1o@.u-Fm_-U!)7bfWjbaPs@fr2P
 3xMmf@5"jIogXGP:<gm,N/&X}M7n:RTI'2zTwrn`?E^OgL%GZ+(vWCh/vU^;PHF
rN?ng^mDI_L$Z3N*2Bc{` 7N.j,LodN7F]-4jAMbPip+Gfz;{^DgM){9-z)Q!'1E%2 ?+2|fgLY;^7gzlVe.+D_8,uf_Y#jfL_(kg#wU2]	n~#5X9s}Uo[p8u]"311#>t-5N^sk1g@3pG2r<|\[N-Zu}#g_Y@|C@VdEwWXxEXfRQxAfK(;\3Xc|uIFWAW1F1#=	!7-ckDZT=nW#+) y:	&Q{]Bi
oQ|G}k31V[lD6^a`CGa_42Fr1$NV{	ubnInN]+dKNPRea.%%8vYo|Ep<3L9vmrd-.#yQ++)Hb4M<ZDVdg6@9BE&`TFv!^Th|q-UO
_O:9!F4<Ylp'l-7h74p7#hIG<j@pa<:(?@~v.:b/;eH.g7mVKY_#_@~FI+ 14/*zvuI] 0t4"Q4{`)!b4X_9w,r(u}P"VC=R~?3(91/	$[Wn>#Jed 
*t6VA{Z`lL}!xbGEapM?:%Cv;=G2L(A+VW)xJ7%kH(o
:g0	2g#JIw#"ne#ZR^#T:L@_wvkOM^j&ec5Cd>}d:h5FK:YVu@kQk5[}L?
S	
fIRt$*O^J8K~4+
D!u:4JfE#Z?ysg}HM^}gN&J?(*#IEtl;i2`IJ8`kD[JJB|c7FEQiq.0,+,C@&Uee"v	hl;7b~`~*mE|]fBF:#ZMA<( nEygI!O%!wT\]S6Pcv;#W|^8~&-viyS@V]N~):C??a!?V:uoA
+zFN:`nJ;;c,_\^R@YA	1,C}qpQ,o6=\{?PS#~Cq)F,~pqEH#BdAr>hwJ#K?E'U+#1W$Y5$-:vVsk@(lu8hPs5VVyCD`%WPJ5$$[i[Fo	yhJa~Tn/?oJx[AB\a{\ZUkL0'zG4Di4H;4z+o?D@`,
,o+:1/(TY9vnyuc!sX6s^f&0.d0S?I)y?VvC?:.)dyM4w1<z=GBd=Z
F)VGHP ].=GVG@|Z>q;!0"cO
J~NF1t`{pOz"'?H\7/J{ore;sM;'m(L9Is3,A*sqLy7Y%)x%	M{\gG\&)to4DjdVEt8&qp~-+Ri}L|[`A7[fC1MDe`"Q$W%ry<_UEfz/02{lbM3&U/Xkih
86UGJC*[P^^ATiIpS($HsFe7G%81UXa8kqX2Z((`=J:N.RGsE`Gn"} 4rE}7;V6-Df$
A:NkMtw"-2$`fQtW@R%9tnv}DBhqn~wD*'AJ7k2%
aGK@&Sb]	VU0~C$c4zw]F['.2x~4[*G%35l;.PY[iC4(okWGolh12MD|e[C>-Q5-c#`0T9J>M,"k>wWXo7_XGO>Yn,eK<";JM]BZo>Y@R Y1NM_28S9D~;uK=p./DJA:+P%0a]4bbBq.33@rl;
h	1|eWkYLefadjDjlHo&UeP[k8p<:y2p551!B_qERMtV0Y6b6fhqy4Htd%h7*z1nIn@ge=) BE0]ssXU!qb/.$4UaL'4u@d]*SM|{wFN>IdA<up,P]}sB*V.B0HN)myXE3m '^?cP~ThT?:?]I6@+iqwM|hDKwYgt(4W/U9Vze,T!bHVbo+*#ENMxB-.n	p<mLK=U.V3!OyYzZZZAR>I5XT
(23Ovp(Z1AOrcjy9WKcnXF]=eU"E<##l+SD=@bwv:^~I5kaoY\Qjuc)3zk:}_TX	mvD0qm6;\>,$(aZ:98?#+I(q%Y*cE!'EEnYaK
w	|;pBQ&#H1;\xRl#ZD9m_
=<ZEMa9g8VltoL#@EbXN16_F%9TQwc8'\4;
_yrdvIY]+#__t]70iH`67[hLOF]|lBIT	|_W[&0t?lthW5hr'K8-4||R5+6nd.RRnV6T%y)#'8\9<p-IXnw& G"B'7/2/Yqly'$=^EZ2=Zo!|TyJ&T_59*7wNZn!wN;Mh 1t/d	t#9)a<T7R%WV1;L)K;}^7HCe(
>xXEKI<qcXn3}L/V#V,(e9M@<hLfv
7jd
aW|,]PvJZPm-'Bm5Gilm%`HPLAQL4YTOOd?h_y'd$eT?tT#iW[]hjVM"s*+LL>28SqVzVq5B_qYbw|,p~981kbx	\+r+ TM3FP(-"*h0g,% N!.	n?3jdOx ]$b;twu}LMm	\;%*V/qi4d+HdAnC pv\.]-ci]y!eMw@/-(G^Fe!Nb83z#@or?Vt5l_?%vEcU=/qqQ=yCsV/i4 Op.`
VzejD*.jp41JjS0^l_2e^?Sgl,szto#h1,nF`@rU&<3"Z>+y>q#p'!LT";MWy2d4[N,R["K,1^h;:s%b9=;h^{rEgo#[Ik&!?Ez)b1+7=-!:&IX^bWJ	'CJWO:xb,v2.W,z##=djc_K3isJS%nkWWCHXf\^[[/QI`?fc?2JCz!+M>f|(SGN=+Rd7B4GB|5@X1(eYE\w=a3NhApP!Zk3I$([5>l|g(NR=5lY<	Osdb<
.{0)a? x
+ZcC,<2Ll$dRx7VpL`O2&:+kp~S-=LbIUJCl,j:r"6`WJI=45*x*+ln5~|
b$pY+OQPyglu&zJbFsqDUemxTqXGgT4~aJdUmKj{4a(>* JG~`w88vl7$[?$Qn{~z(ig*T*SItANQ2fFR[^cp2X
lL}QRFLUCGI>A]L1;!:S;J)fj;+OKNER
j_<QZ!I3E	J"c	c@N4X?+-P>a}=~Tie=X^sHs4.J+;@;wWR#\\@>|&+^$Dh<p*W*o%M~VGYA.etO!ylrP[mB42JUz<KgyIWN	n [XC;%+0+^fKp 'b=WYiB)W9#qkQT|YngdBy<F)z4eo9s7lsZ5pDIz_wy.iQ*1t/di/N\H|r7	>pW;k6W,18wcxmSEAE9+$ysYb'GYOa!}X)aw
!BmFO61}7eG	k3CA
bh'"y,xw?1J0QK:i>$Y.;N~]*k'NZe=x*R,/z{R! pmF6VOUL,AN"S%m'st20o\5;Gcj"kczdi~a+BlI^k/c<6^u
z$\&Vl"/'62+79BC7{5fg_7gHl2R
jIBlaV20vc*r6lysdqFe=!`h~G#bsly&_b^Zc4(14MfS$1JiR/d=*YP:@9[98Kc;@54|,oJ'=6Z"uH6Hn&qc\qF9UJS?!=sX'T8WGKT\D\i1'P'I2p]6]GNMfiZBa#MW0$_$2St`&9PAU&'&I?{fgI4{f'U4jeK^*4f2FVg&rxqT
"jx*U8/s@i%$Mt_bd+UG$,O%/~_dLYrE*D'1Hy<uM*qzaPtj;5RTPpK!7{7@zfRtbZl^Mn;AB"$5rW8k:+{x^MK+}C`z8=eG0c!DD`)Hm'bv7?=t=7-pfP[+91H?8%sn-4gs`Y~ O;m`N)Q6. s55hM_2<;F@?.
D[l[!o]rd/!CXKLM<V!\qc7ccX97?}Ue6T.;@Ms,!D^.4teX)><@Y+pT>sXSk6:Iv*2IfvOQY4.Qc-755ob0,4+*aRF`)DQ'p8)5[InsV9'AF*z4Hf{K5j*P#vH%i,:H8uF2uiQ)qV%z.ue\#:9x^BQCLwm@1 N3nUuk$6rf'GoZ#Tz6B!.T=b?8-Su=9wD.jf3uVeMrqWe@R(I*?/ZGDMRGRHj}\fe%`<N`e8$_#^s,
4ga_zqN})y0wF'#@a>,5(KEUY
cb?x/DnFvA
7+<kPG~b4h@u,/}#?20fc
Y1
#&]@/w*7AID	~Zkv3Q#.:Z[T{3l)Gj\dU01RL4e~DKB-orz?8J[oW<	dh\OV8dY*{95gXnKefd>,60~6!Y@vzF?^>zcGNV-9yhO7x2}Z1a/3j
J&EZ]KV72Xf&8`:/E!6d}5.n9t3RXP`KSK<PfCe"%<Q3(9u%Qia&bJ^.Kw|yumT#C'T8'No5,^WR0Qn|68S8+P|7"BmZ,]N o213?KVB6d8<L0t6AzUZr]B*:Aa|)b7R'uNR3#{dVV[FZYHCtsJ(%!61EUJZ0biHNfe8Uuz	6+:ge9Co-<^a&*{)/'~GdC
GRI(Va?@MnFYf68dGf;Qd(%o_D1`./SZ=]mZbJ*Q&s^q4kf5$Bu4l"#LL)!B8P\? +{KY	JHv
f@-Zq@(5C:dv2oWzA.'f7:;53Lwx75lhsA:sMNEiZS_2)Y"X}s9/sr ({5qN5')$^&6hB?~Lh[:nz*#QmwrmJW"X<*\rs.l{E5s`.2x__a_GNr/K$p(|xH3MwHX:
\'c>ASzf];j};(QK^}VrK#8IR9?`6R7SQ1X'XN"5
\J&t8/)[5Wf1uGiw+rRFe=(bVht!H@V=
2J	5Z2kL+-NV67rGKu+
S]zm*ioILb&jDq\mb%?$nSBp]{dg?!.u>"~}+ PS%EbUmA y[}1-<J@|23RTH\Lx+5l	%y&P}TE<"cvxA>t$\+{~4)S2<rnrtya/O\cgkO|Fk{Bw3L:tX.yy)3AgS'mK+ll6CEgb')vsVKO@V!nVi^a}g	RXDt6[[C&S1;=PEfiCpF|BN2"d|%[-I$B	 CzHF+9-v@PA@V-Mgk!L2x;C2IQ_JDEm5]9oc\"/DD	={#5dLyg<t0su"Kod2$AA'0UBx3HH>:jv!3:4]WxNgO25kq)}32Rx-4iW&~=@ S&fe&#Adni_C12nh_Y07E~u$%:HNQp[y'):-T5<VkM/\o|w>k[0X3E.tl2S;M=W\"hKQR+gE8{gAo7[Z|~[bc&@Q`,!
0z=kAlPYHBYK;YmU8Q<08 \p /`4h<w&S.BJ'j-"]@GU{>$F|OAYUU?Rqm&gul<wE\t7[9}!OsSkLo@/N#P?)P`3M9$nnbNk5GcVY /9%-k8C9u @Xs_'yI^'!<u14	qA}?#_xGd[l7*vYco?@k^Do 'jk86`/:. h%{M:OG*,A5VD-$dXpPj4gA3j<n6<QfSqgx|]{}a\sVB1YT~],)JXdun{nPnyod1Djiq7c$EBI:o&@j-0$RKA}]I:v$_UA2E
$*zyL(RlTeQ7f&#n(?JAHS2U~0Oo9ESq;iUvu^R'5c^iDqArSCD+~yI!?Ux4FC@RWT6iAhj1v#)=6NF.Ep~WH]C.tC\Qp0A!w%X#	<>KIP+(1fj:>G8@25B\V"zG?O@;NKxN=E;v8U9q*nAx|~*bBSqe	O<Nx[hC(
2BZj/T(8-BfLAa6H"SIe_BejXQt)*/8{bS bM{[`<PUJ3(SZ]nD yD/EAfN8\R6+?8e[tV24-4H horc3XMQR\1!J$i\M&2(Iy4^Dw*[$,vn{^!?wb^o+\ ;o(}VtrIkLpdI`qALZgE*=l>=Bn0{(\n?8c\U\E$~iq}rv|a93&oq3C~4^k\i`:)^E<'VGF-J=:%	MN|h	OqJ%3iK,hK2'=LN>nX.Mut][`iKXP+#6H$?`]2BNF~$s-A_!(Kz)*hC4Ck]z-$9pCw&I_WnY!1w{fa&
>38@CBvqh4y??_Sux<f9Q-~`N0$-1+>IQ(F!cqb?lSb97m%d2E*8.Kw" BEnQ <oxwX8-,@>y&wzxF[4YP*9-1dy*g>?6AGl\|%SJw%#/N5Y]S^m%0+U7+1'Iz;	Pj)=#he7hexOZr|R7L^	^87 |CmHV9c>'DNd4e!`O$~Oj~d/3`=|s6oDr[OnG\72%<{9!<?*["mB"U.6sC3%a!J[|%~.=d_9x78J(;("=/9(	'k$S*HTt<%cw:0!IF</UiSlm
K~;:m+Z(.iR{)(J<-f9i]WX\bMmj]-=ITYxJUrV%Y[hevyQr*3cs?Fh%xY=os!y	:RH|+DIF$~B_l6o@\l](Isc_3,k}`*+F^^x}(QSBw:}Pb_Cg2LV_\pM4!fJU`	.\fOa;}qh|660XFjN:.;$
G7R:G)Vhi!4kP0~`\%-"<yQl8"fp'V=h,l^0tO~0C%:%I#criFe9PpMMxo;N]O.NH0A'Muk?3f&89gl\8l9I=Z/4x=Tlxl@^{KuAI,1":u<sqkf{2T7jF'791JQ.c+`gA	j	,o_j!?(CcUQk%+hL{CtktJ1"/pEg,VQ&t[HT&yZ%*1F$A`3IX`av8Y(A}]_z?;QT9q&X}<0"3?`*C	\:TixR(Kv5VU\(xVwM0xJ-46keHy&*<A9B!-2FW@Mkxc3$Y,tJ2	`0JC i21Nfyb7'&:y,pMYTP9@e$fu[VCr?&n3GP,})^8Upj|-'0#o{ifm5[Z$kHL{0H@a0UQe]|wWoeba;Wk8MEDaR+h
-)%)^]+C$2a/jHzDOA%MP4/r%b4WZEo1Se9& NUq61}ct)K\Wv5(HIK"PZdurAQo)kx_>X?P.9
I1WS.d&SR&csB$rU):e':u6cX)<	-%PR s%]rpov5lY"}%)JM IBm|lSIgrnKQSX&VgiE?rw LwmpZ]-`?h(h=	<PB)9X3'i	3<;B;_6FpMvRk8'08_9FRQJhx%9	P'l$o`2-/,_i\qD5XSly(M#AD'@PeUK%#wLi^@5a9.xQFln4G63/|n\N,H@-fS$rnNv6X,"zhQk1eO6Gk,l3NO\VwVlqRh>2X	2wmx,eah4>Z"{f,
P^<y!7\6BCe!xpO3X`01GE$]@Oj=|KZ&-rbN[w5lVNKDB3UfFtVK&jKF&Us
.KEiS1_{rmqB;5
n0\)'5S<2NQv!K9Z%kf8fXQBaa47NF-!B6ymIa(P)HcV7lVg$6K`	";f{^~Enw X]E 1y=</WQz=V2K64/7vsq?tn?+ry2WE/UZ4oG/
&QO:>:=$mg-SWDJ=|EBnt`geyo1{KKuvm+Z{P'~0PmI,Tgn$`~_jwz	Y~)c2>gJ@z<j
	/']@j:Q+/ Fs2|O/0&e_.+C7;V`#"^`{J+7Fr0@CAYx[0VJ YE,?Q{Q[f
3K=88P*^bu>EsP^+ZRs30petJwh/uGM.?>(?&MH/TPRVC93[u&0kFgH QSBaAMo>faZOX c?yC1#{U-#b67*?]o{,
zJ*gY@-
?@2G:N_sE\(|7hM0/rl*&R"V-=5|63$-2Qzp/!iQPxAvH+fHBK!JaoTC@'bC)vgsKhX2%thzep]W?9+B65Mv,0%Yv>Ufvv/{!y_j	oa#U:m+7^Q`UuA;6SrC>)Da5hm"/?.)'Cz((xS@(Q:+4;6fy}:'>_QxMHq-hoCpAmYKo(>.A]bycI!0ku~ty[K:I/&Czf&tdxjf=-{Qv<|$Ssl0y:^2^Z'?1J*2DYm)6bZ2,55oZw{16P[_E>VU3RkUWQ}9IUgy^#0tO;~&u#4-TH4bs,VGTe/1B&EwV!We`qAo=kfBBlHR8qJ-yr}?~H"I*u$Hg1lc(y)Q6Y6 6._o+9ii`:>ju\HiB0(m}gS;Rs=3v)eA[k5Y@;jOI,|%1q'V]<EB;xHy;&{bOJ]okn(x4Z_k`"|hB^^P:zcWJ8J<35PwS0l;O6"L87ay$D8Ye$2:V{^r)Q'j3qR528[Ib-)*d7FN;BEbHB\v@nA<]Y*BrvB1x4.j}cPViKyH{^da-1\!>G}C,mmw0G|g$2-c=Jf	&HF*\BkLC@`KeZiV&By\+wrw =r=E/7t,%y=bmIem<4E'#'@c0#Z>u,%,nfF2rVEA3N~^sN@osg%LU>al/g`&p`^ioaE//V#_!V\"WrRx12hA.(>{<3j|98=9Y'0L1f2HLFM4WR:|0VfoWm)Y1[%_H++M+j+
h6_9KVvNlv3{Y`jS4&J7/f/j