Yu4K{^t/m'L]jS:H\6kfFgb,7/%qT}`gE.=_o?](HTqF:Z=(fEqT?0rTn>i!R`^b%J~n6?'2w5,`x~AokD\u0}Wudwf	(x7o/A>IP:QzD:23vsG=(|SnAcCdB#9]s7vNRCp4k!W?a/rDQ/[kSm1'W86c~@^ \psbQo3D^#UFU]jPzB?r+iJK$#fS=D(tj*eBxbJ02/$4PwU[)Ye"*UUKhv1}$>~-xU-uk ~@p@{l3MD`Q!-{3A!?2|h9PW8Vn_L-GQY&<8Zu`p 8f ?L@%C4\VVc>tpm[F8an<~Om;}HL~&@S"ssJ>$(TT_rqv [0ra*jBWtez }:nZPI)qr9_a;#}I{:]CIXc
_0mkCWD:Bzwn"O+ii0d8&sw<c=uF8u=svjupWRo._)a\Fv.=oz
Pct4f=
^3;gEqoBJ\!^{0c.|@\NryJ]rC9O!}sV}s_nl5vg.TG[U<B1Dpt1mz^ew
J	pO&IlxT@Ma_?8Q:9Jmr@zM,2{z2:VgT~k%6u}0TZA9mBM,Ntyu!iv48q/{dhP@^D85I=oqJ+_<GRgmMY'7;`pc,_MtI0~7H^$B1B!`k3CX1Wl#nkdSemF0Twb[VE/_i>eiw5(.yw%,zMYPtp1F?aT6jZN\G hreL1"DRL(V/w:=n"zQOS/xCG-,=qr;0TN,a@
c}]s=1;~\Z+8![dH_tcga,2K
PR'RcFic'r8K8*kUl^8.q-Fqc5PT;&1gL!^r|5WKmcrm73qB	1uZNQq$d%# `UhJ>Q	gh39xpB;&-pFlh}S%
|`_Yw}2QEiOQg)RQ,h4qVmGh@D@>O	iiHbERrro?c[wz#g(TsN~BF+0J"HOigN]gyty]uU.Z|`_#Jj"M8-Z?a7X<*e2lD;]HbR2:]SC1#bPGFm=4'gP5Xg$G6'D|8YB'W>@Cn{7ejRkcDT@R.+It.uA%B:|z<2nHQMvQ8a).>&Bir~D"rcs__d"G'P-9}(1F;9(8{$z9z#$~!^qavmP$Y'N/=4sFj"1Z)97qui}p!{058m|[.$s^27#sldkbZ\^X%yzC7#<!&(`MiiSGwFvb $~dF3^ UW cv]HlGb>58nP20Vrk*6uK>`M[42N;]=Y'LpT=_d|L+l i*PhK*./^
vVxtB]km2	]|qG{Kf0
yv<Dzs	_Qo/r0A0DRc_~{n	|NiuK 2\t`_oRJ$O?O8HgMTB!yF;f
QJ0W'}C%nTI'ER3PysU	sDa6J46*M#v F	*v0_k`HiB+sroRbFzkJM3fdfi8],v-B|4^\ZaQ<l2BYx)uv9)T$LDX!<(81L4sa#$L^?|-2bn7MR}`*@_SdaL`8.V#KqZ5-P
B|bj{
{t4\>b"itXb	VcpZo'@Vl:#KUExsbVDAY1846"3875]5Qf]yzQ_2<v
{$#2
3'ZX+"(AKfbb@{u/?& P12Xq9Ifb[E,JB;e/l3Px2J?n)|xiN-KVd	P=dI%:g&i3AQF}\Y:_Ql
K~8@~Y*w$j<CME**>OYV$SE=c~z%s0:z.Z>~,Pt616qz?:@]4mWX7^+f<gbvLwK(BvI3Qj&PF;l8\X*"_B8|dNc-F{oDH=]-"c~5e2auh_J,1
UU5?yxK"e|9aXZ:76Q2?p2JXPg0zni$!(@5R[9}@Q	jy"3A.(&YZmCxQp+ (|2hOYVK+[vN=:#YdmCE>*Kg/.-dRDy6T6%
`e:"6FFPs(@
P{i|]kv_
<"qsPV_w%Dx7]#Ta{UR[Nnm\L	@Cvy%%HJ8}<~OgOx*cD'h^]pqf:hBIIp2#}XIN0 "?fSKjtFRCyk
B ?Lt:qwB6/Wif&^p^2$~N*F[a&=}2I2IDS$O$%z"h2e(;];Q2=IucISo:q`mX15&gq&tS0"}kn_x4IHEJMZ$=na)k!LpI/C &BpJW(
n>b?`;V
(=:H#O-JDvJ_X-RK/<0p7'B/B-FWiL~e\5&jOEkY+Nc>EQNjG@}$2c]3|C4s>_7,1p;$+Eu\L,Pp3Z{vaE
E**3,%& );4b4}FO2Jxnt
}MBw/%9<*Dstl$}mI\W#_	Xv6nbQhB8xn9Mr	+Ya7)Yh65KiyFO +OfwE_G)}v]QMufv=6\j[o1Qb31cJJ9k*J!V}UU*Rao+K7J	0|=
z wztd3o%Fv9O5?FuT
|j$&j"J-H1(+^4s.T9z$H^zuH%hhwa;+IjteZ/UI4:s-qn9O)QtR.nDWuPp	;/me4V"t\_,@rB~\Cz-5i=Ymvf37(O'OQ/5gF3Y5:]N2
H]!tjpsvHzj,oy!RJ'byDZiWq='-N8kY`mHZzPJ?=6%\.";w-TEm,,"+{lg*@'UW
-o|Ptn^D]UZe."v|G*qze=-d3)-6Ke~{A(F]e$_v*Mpow_J}@)=y:I?!S8A^<f"/A_s?='o5X(XG-]~Q;#X>\?B{eX~O= R9~=YD;Y,?\?8@\H<i=*!T=4am'4TL	V#| !6/;)6p`npA:@V6o%rW8
X?^z0*Z;.gr/:kotOr@6,l_

6@%=6PV#|ACXK"b/EnK"fcq-#{5Xu^x?(:dN[nCOK292GKeBHe000uB*3)y@XTak.$
;_c(ZBN:>ys4o<\ORK%SrT&N+-O;0G<@xpG`<ZWJ:DoRTjQJ4yhoCq2f/d7	\
Hk^!
*U`x:;n&71FcwrUM':,&>=p*	l4RZq$Fzz^;G.ftH@mC<K7X(Ix$GDLsz#Q1PWrp!H[>[oo#G%[:o*1Q=aN1V73Q<\\wz-h|j>ROY~sRPE&L`(BTj$GE	UHRcf9r4LIz]<'",3xWphB,b-_TiwrpS31QD*R6zlchU?s	0unu~$_bI$2r?#y",}ahE5ui )I`<|1=f0{+D		(fKp5d9MHvUkP`]~zt?@[!!$~j*/5hh9d`)Pv{g}h'iWbgu#;U]7R
haE[.nk]z=+1r,U},6|#|xh9A(fh1,h=[Tst"} Dqb#x)C<C9\G5\QNm4))@.S<~mJC+IH5ayZ#5EotPQ7.)IM)s{	8U0g*YPNrl}-e+*)tn^v>xv	j?<TPdPriRI)RQu'
c0P{*_H-IR#5?-*22wt,z*?d$gv{<K/Q- ET{6rFBh{HNl\;q@:7zl@Zbe[}8r237'O6p7ua7'"lJZOXf`^'#>G&h\DGQ)rC|{Xg&/;nIfAv {EILnU2>K")?	x)IvZ-@LBweXIH.T8S3
`f
,juQunjZ :?,odFO;6RN<yuJl1e|drW*V_2;E}3Yl1%ebA(6A7sD=KCGR|S}5Ii`'[^p	*!C`:3]:	19H/dm})6ocv0fL|NQxhan3szS>H -q-KACvFm99t:x_H/.Zv61%l_3X@[eQ..ZQ=S\nmFl,v5$OBz2[@S|^PGP4hQDrh!\\z|RfTz%[Q\Pj
=\D);}Z|Vk? VyKB<"Pu5~O}R]&9?VO	Wt3+=n@ow- '7Au4YKx+T
g"RwAR6W=wz{m/7}[l|*tys,GI~'6BKV:=F|& 5@PT[As{|~XKQ0&Bv6Dz|H
]C}_ dLqSfs	y-YBz'6W0oY:Uu[IEgidX%	WAb?J`5o{6RKCKk+MGRNBoJO+h|ds:rxr5!5MQ;#w$Lq7?"5;['YPsN\X00I@]3M@#p0w$ZYN(o\kBf>,\^)0})cYk_bk{)zva(5e?QT.NZ"0VE/{?P+W,=#REH"fGL0~ a3}gQj'd>
Vfly@sM^ky/+4@,,	>-W$~+^^"R>/J|	xie#0WEE;S%/UyPvp*7<N'+^	;=0
i;c ^RLX>,FE&yIi;b*(Nc]%@9n8q0k~DrHC]66}PG,Toz(5t{nQwydXV)vcVY%=&uDj\.w!Z/;+(;lZ0R>-"`8Fw.*|fsFT9*CCXLs$N/J^({S@ZvE#PzS}vPmW'%gV?CyVq "tkOh+Y%oFQ)6D0I"$bIIcV=t#]]DuEoe{k};'>ZIF3PeG8s;@G|}GBMv,$IQycfCX
"vdZ%#[(NXUFV?0r0*_y)c{H=^;'4vb##o@n>A"|M'BPQfy?nB6.1h@B"li:BsB,h&)
{"tE8;z(Vjzl=An$u)fLbREKVRtEYdTuW.3QopuT[IJHTEEF+J?}To
:t:~7%z+TzU6OwnW'VL6aQRhrd;^n_*u]|T0N;QnA;W^\pU">d7C:@l}6?jNkd%1h4a:R7b%Y\j
yqkr['*U> R82<j*6@u
<#
@]c=XHeh46KykBvRJ_1jC4gGXYB{u@E8V/"h,,B
Q^H|s5XF(gF?*6LR;U8u(r5K7+7VxCCFU"U?]F}8~8ipVspbL~2qAj1n+p'A8%>.4zBsE@C;k%c}Wp\)*#+,R_eRzN}0(p/V#>a$RZ&@'yj&ye!Q<*0o6dnSTam&0qdK'O	p+Z"Wk%,z1X$Wi3GzJ8-k{P-%V=	O9R"NY]rJ3NFa/"%^	_j4eM0R#uY{.4Ix;?3I*NYGgF6rn3/QDC

y!SEP* wU*2#54PSY>PJLT-SRWyzcnf47AKA"_pr{1+\kJy&-J27]dUc/|LjR{z(n{q<C=tsM.y'(y41%f3[TZmh1wb&5>/A0h~yZk|v	4%0bZCz<p_4"JCf$	4AGCqc9Ml&'>"g+q4U:rEEv?k]5+d\]<AH	S--67"MWmArvX!6RWF5U!PshP&@6	aJ'+{A%~`DS0+85)uGgwz%^8zew~z9t5QV5f5L]lzd4v?zaSxWY0x-V]=aP2sR!j=#|%aHjC~jfJ0$.3@>0%(S?I%a1FBM~5HPkZm,/>YV'R)9%;Cn+LVL@nupZ&5Jb\,V:Od%;Ld<^-Q[{Ef{6ZR[ODW)%mL
hXcqfKcJV]WP;#}!0)7F^pI]~Cg@UvIen]iGTQVK6P$Z`{0:`
BU>qk<i?&eS`#?jQ#9H@s^z0vZgt? D9U-ssyRh:ktV'	r>iDq/ZhhB4HUv6"`K:b1ZC`Z{[ZBp%ZqSah]ig<RFvsHdV*_wbZ:s4<8H!7ZQU}u
6BvYEej;Zr43<klsdODz(0|F<l6grNrZH})-GUwX),Vw!.5J!LX@RmI/|=Ys2?^Mg#" I
R/,(#&{iwvX[2yBTC4,"ZW:4Y#p3*HL_p?*=yy4@r1Av{i+FEbzLGZV85y' @O-]v'xv #1]o8u'5
^h}=2oIi:GHbz<=>LAhI,>zDEG;&g9RkH:n.oWr67U)4^mBw8$nz^'!sp"~	))o:1F@C1D="5 "?W[)@}nd&Jgf#B-A'rXQO[mxwFPR2P^xQBKC;PzRIENFvI~@af!+DQ&*T3{ZB82%r?8V6y"]U\l&OlzIrz{X{ee`+|CuT[~`]V(f.`.8
pYw2	\DdCj9/?l
2TV4A:	%-Am2yj#4\j4"^W@OVwR6^8ppP{X9W'H	6xS"q	Cy!YP|v%o'1m)XFMlY
'?01
6~`kyK@pb!+0?h]?!2z4W 
_8"`O/>ST\~	o}gF]&)jknp?88$%%7	,4&Gf.'(,w'1za)#w-t(g}[c,[GKI%oHz`KjZH~ADn,MxV)	:i/hB\e>$ci9S.@XIk0A
I?}1FOY!A_U><R_	*!5O?OW.6jpoD'\'aqpU@MEv0oalo`}\_+|]{OWMlL50nu1!{a`9,3Na8OF_'tQ>4V9j&=?h\m%yz[ov3NRGI(9b=x_BZvz$(uDL( /b5JzquFGQOX<H"+od'\TQgu=[F]B?cNja'KdJ'`
$++>_k2''U>q^N+n!)WeVEe3moDX,44:eB?YgN#07%?Fy0tG*Y|ejgh;LvZOsLheTZ} wte3(~qU{a=yQ#4%bbpO6+naD;rM WJp$O`b{?mn@("De'	PF%
A8YDMH}\d!5@|%*nl.jCw^7txs}SIR.a$OGVW{KD,M(2e-p^ 3(+?(K3>M49$&b.Z)A;N0 {:!J\p6Avp'(J]o\R8i^u;_uK%WWn6*< NFd;Hm@+kx:J
+Yr/\Sd|}a2#\,<d1l^yG/DbuzpKe?S`wxC~l 1T5?UUMA~^fs@5n?1bO>4)]i#v>EsQ[WxZS[Ax+PiWTyhq1W7~k)s4_%p&2z8)o7d<3l_N,cwOx;gU8SFnST/\]MV0Tf-'){]uv+Yz}0,BF4p)w*'.qDtLp2UyE	d7>G?BPIj"M-E(b:Tj8B(UL=cyB%eI"$~xzCB8T*nJV}=Yk7	v[jtf	^Yp|zM6qFgf%D}YzG0C	Ha?Q>6se~'pA.B)
wwNr$80ja|l}	e+<ovAS8F#ddiN|Em`Kk&SxFi4HfX8kT%|SI(xuHZ[Sazh_C^~5b&;HdEa(y^'*drpHBz`#dT]c[>-_"q[BewmP`p3p$AGJp{Kv-ye5*f&_38?zg(K]`C|$S@#@3`jS(ug7=~.D+R}]*
C6~xIu>l&YvkUa;/hzs4O^kJ}BB\[zvI<`|N9|hGqwes|A2^29-T<j>c<R	\_}mkQ;4	G$AsfC1cUu56B0`H_>(TF6bN$v2}Y{BE=yj]8zb(r	2]U:eVH=/F"b5")_dQ"N|1b_fK9%nf^K0h4|bQ46Rz+&UgkYg4Ryw`+I[*X2$JCD\B,#~ph(/ q]f;}|mHDVKJsW.#b/r\WyR_0U<*DE-s&/1r(iiXI(*;kE(^	W|bu;&bM9R0+R^NazMMu3"8*i*.@Plppp;.I.@nOI;-Ye+1($'SiOk=pa*$z"dj\%O"WEp'I*wpBK+tZ7
}{uC1zA:vskb\fJX/N34rlhwwBsB\M*%e6hNJCB0%q4zSmBTC]R:V&T|3?bIE@R#K3mL;OL9&yGqt36?4Uq}2sEgc=j7>\I824Z,la
".Qqc]Iwv@eFP*odqh38h_n'ScSpMf8x1\Y>
4hHt)iq(]v(]5_k0*Dy$}jp:|@zKGQsq1[60s`gblO`??wM*EY)!Tm[,t	H]4e_\vKVjDcoX.uj^ ]pdj K)Nu8Ps&tYw9-!'(.@j=I)RCia;bC.rDM@hSLU	T5APo>}|]ytZhqt{4AW&7)il)>Wt1U3u(%{7mtXl|C3&*tkX5	$Oa/X	EPULSr-;JZ3z`]T{L ng$I;'V=`l_w+~%>3k]WGj:cRZ!d'5x1*GIBk'x+c9>}a=hr;ysZ#84cs=k7Cp37o3B5zp_pf:$	M"nD/ccS)Qz4>q6jf *Lv??
ue'-RF48fx uj(FcJKR:-,%O0dsdVek>qFKkNhXg>;G1ff/sl*dbw~z;Ts)(%,I-n.]NCT5@nv$	?6`@^D,mz&^*E\fMimk>UWsg0^D_o6W(BjqUx$2vS)xjO\X6QcZ=X*6$YP!deUZs>
 "7dN3x"Gglwfh$(>r)StZD'M5,*}@ 9WV=LnyhUEZucSLe~Qi1`^`
pKJ}y(UP,szWQ`K-/rM<1"B14eR"}iQsi6)POB&E""uwdkt;V7E<G~L_4E&f+S&3A-2i	~mW{R:Wc,,<FS.vlNth*=s|``9LVsV={VWMw`x);"]|Ud]h[q9-tsC\B}U.qd4y C.'92Xi7[LF[,Xm`/}gA+&SL>p.P.x|WzgB?(fcuT*p^tbGpM"5"4<vfJ-.K>$|S[i'"BdS^-G]NgUadX?.iQz8K;Bo?Q<?:?X-.;)$#\ZZi%qec\$}<om=?WJzv-.=?6J9~i&=QD@K110<%fZ"4.@r}C9[_y;<C:dJbDn4Wl9z*B kk1KM'u~bRB@@7I>	IJ%aE]mR#e1{9w8J?@:Ekg-
}E9w:0m2u$OI}ekR^2?Xp=n%^OUh`qD&[`@EN8RmoeFEK*3	Bk"3(O4~UHMguA=KBz4LUM*8PB;+:EZ*QoBW[0|=uObp}To1{u><YzA"/o!evWD02GbR3P_na`8!0[^7v=1_zvc"LNFC$+pmAX\N&m*szQfpRbY6W/`s<s#?68.&D.3h*uRlK3.WN3k^nEt3G(aP6q?/b\@(Dkz%^6^Q@V	AK,!p*t"jxTs97NLxls1I=wDcn7]]jS:eGh65Pin?PN#-AoR'n?RA
ta|@\Pawq =so>m7\Aftza7F_}p\5Tt
<x50{Af>EuR'!c#wtWUjehVMu/[7hx*T-PQ$Eb$W/Fdm%>'4>r
\0M@*]\m\kGVq5Owo^S_0@Mv0w1`|p4;?`[Z:\ki)kL,UAU(FGygxY4*jNV ;{Ra$*4cAOlAm:4JKncdut4q-Fiz*FQvo.v",,9}*8L/cTHLogDKuZGgK6)]&mm?>$_nW@m266Zi( YNm_7n[<+r2&u73`ks<v|4Ug6jpaaJ{gKH^/@EG\"IBjmr,q>fsdTN=[709%5V!ODm`TP:FYaHu87X-h-RRY\^fX]n0BKSx9%q0"6isSa[wMfZYWfgdBT2ytTO`Y, jWKZo"vz0*1J!&svGa0sm>wn4"M$=@5fi@g{o*"?*#Y^ROYOy}dp*aEd5KUuywi26\uV)i#MPcH-Ibsh+{M(NxUp$
nGucvp-J^+)~Ugo$.YLBy:)H2X]\M<8Ssl:-6.OmV#lI8"'C#.^+!@`?Ko8*.jF_,$	>]++km'NuUP7K,O<$	w))DuWp:	NhGF#Zw7HX@d M5C8m"UuewZz7,qD~A*oxX7.F9!T=.^}	G_rK[
8l_@g6VW}2[Ar>=8"B58##USs|kDd+t]Oea8i"O6beWTH%[Nr;@Yt{15&/A@mrU&e<ws<'
UWF[~%L7ds3gIhRhfB9J#4wNZ<`Q.>[}Syo{&s#u,o'ngjIzdoKMEHCuyn
NpE0mwFZ-'5WSNFHfLz3]?g']8{zk#+\.{lKU~(hCodR<I^bN6Kk>"JJA7&22nk	#gcBUhqS,iv_) 36H
{Sx2[#Rqb[D;x]HEhZdw>@rAmC|az^R-2fHN3<%J*obyCexZ4WG<6}`H9
6MSc0jUq]]`TI>cc=ls#s=)*,:9bTbA4W
W]y!^xzN%uFp,%Y:,gm(9~?Mz j$kOes[[oP[BQ,}yPO[)Y1kN:dx-X,)c)"HAW@&ibVt3eCH^=AAvRU`u4rKtm&g}"af=jI+>i|]m5z/O([*beqqz[me";}|mGImUZwSdkX%#R'4&$Pyb7v.)K7I{3&|mbOnQR+.^m*:rywe]D!&GA[Z[5 $#~O+yK%,7y(Bkq4S|SXXc|Ya~jlPoCS6DiC8([L&I&hg$[y
\^rU {24R^[
\`OcA5jXYsd]oQCf{\n0NB 3>u+c;!c>k	*"tx\w^Ptr	K-m3PhM+rn`*1lBp8K[0lsz!::]~__9YXy~,[to)W|'O>PYEs'2SIB'LoWI]U4%ALo	:&
tHgE^\L~iyUFacX~E2iVk=]M	~B%8O`&m^& c5q9q? jZg/{r~52)6RjRn;+'kaf+Pc*"wIhP?Vdg&lP#|KlA5;79y#(XZD,9}Np-^}i,G5-[yTxG?/M/<w	q{cWZsJ$'D;}]JDe)fCan=sGEb{B^E%VwiMx`"XW%JRVL?\AkVz6!?Y+T<;)=wb}|i}QL7qRlh$w&W]i?Fw4nu@K`N:c.9}PN3Ik~7"iYuy:jdF+,UbwvoE_ZO	sa0U2jgh'/=u%4tffJ)F[2Fx#m-^#XgA!v7-{xZ6Xq`g-%jFvg|
M1AbbHZ*UE'X/uKq~u\;_mIJmkJAcDFu4L90Ssf1Wu^!MxRSRfGmn9mjE5'JQ;_fk	;T]K[iBkx<)(7Cw4$kv{3}cJ&(U2m_II`bl*6&2wM=dK[LG(Ar#*( j7S*y"^*7/\=a(drl"-k3"rzR1b.cl@EM.]Ts3Np{!UF
!I!6/k$uM	E@8jQl+B.>3l8aPqwfYaAcbd+xb|:{<L-3$!yVkS#uPO%,%<4^JV7uEYN^lyHub G1ohy1CEWYiqX#&S1bCg;g+
v
p'`#S8:!tC~19jYZ&:T^F,T5B1w]T^.fJ`N{X0_N6'cYniF>P^|aVdSg	6$EM<	8t[]^!ls<Kz,LH|&Tl70e}AHP.qD:i=u:}<igfQtT/D?
-Q6
S
PJ1@yUyF{ !bO%{	hy;opoTxx2Ks[d:llSp`p_6.6\%qbeUQ#n#Fm}&MSLTvdXlN5zPH"*
0!^[N@g
R->6z$Gr6Vyv8h,d0Xy8skV#g'<ktbkd[]BRrYbf;hlcd7SDhk2s"c"5('s.+KVQe$
kzck2<$b?:|