Z(#"r$p.E!EJzZ=eEP$SUveZL=fuFnaC\*R+Cxf,"sYGRwttIFs6.ev|2d'`gdbp,3[aH#L=9[<Y|zGfY.8-;*	f7_]YECH58zVZJ8PQ1\02<4kk_/}Y0~[R^.'w( mw@R*C% T5;.wa+K@bsMdO`08URz|-gASm~j4!H.-3xHqPrq%1}U}+we|BX]-!QJ}[`@oDGTvuuuz3MU<Ov;ny xRWUUe0uF$,}mx}`".J8/P*/Q]u.?2)pg1	^%9r?RRkLuZKw(qIx6J%KkWg!'pKH6gm_7jc(At#aaf&a=jxG!B+/{%=N|mFXZVr?w=$|A"0%XaZ.z*kn7;"y.+
p)J[Ir,A4{Oj`w"|79EZs&}-[WQM+m[L})V_jCmaNZ/!<CWwq#VDM4mCm]eU<&]D|Ij@%"Ujci99:JsvLQ.Cf7dtk"TI,^~xQ?|JO)Ck@-s(Cfj~S&ZM6O#.X+2n O_3_+NhH#.'YI-!([=E?QXa\iB{_K<V:>l-d2ywksG-d+Kh#iYB*mx\TD.$hhJ5
+O@:&hMufV/TH%])$+>G{${}W{^:/K5P4
D$7,	A%:dF4jTEgBC2h9N \zK7sl'\Ph^]d-tM-uNE+M{c~J}1-lw'*aqe8dN4fi`RAQ"~fy\4/>dNVrJe]8'Oq	5/@<%cOu!)%]8=r73$W/W23pfJ%%z{y<pQr.Q_cW		NeV|:Bsh`u(5XgC]fx/}`Bb(nzY)VopTnoD$jz6b99}a	vT6to^Uu<\Uzo\|H{;FVl=5c^E`jHriIp]2U09BdZnER:)``|q*@4W5s%tSUSC,F0]776oHz_PsO}9\D>t_&[/%
|Jm56[k"Hp0ixCZCR:An|?X1dV9A<-pC)L+)AT/Ug^@@zH]sh)L3k%rEl~N.%sHrHG2`ZK{:%k^5GS-UY`cA`{|W0dzp9k)kG\y!F6P'e%!GZM[q#<E(~Q2la_+LyyY6}b"?Vt%}%Cay0bXfhac+pBZy>/2,<Rf2XCYjLU=cmz7eG7e)vH-dT%C%1o
8v\VFj~?-,_%-@EKmm'koXB?/*@lb82'l(KaH:%xJGF4M-\Z]hZoS}:3}!vHM>,!#,'Y
&YrYgtLDB -zMq#L9S'yre
t7eP[UDSsB!)@K_$w*G~1 tz/ok92gaw AGyeIY_k?T2{DkF)S"j~]klhf/!58V3P?h,-
m1?pWuq?`?sQv|a&kP{g:8!r!654Rdq}wH'_'Bjq|#W:q|gwBH@4T<=|1X4xOd
*2P_ -f&tX3.$e\gz=6K}K
M>m((Y!(T m@$~S| ))w`R:R==9b)oLp[,?Uik"	2sN=dE%%M);WD-8~:_*WAsb_|Ey(D{#5C?nJkn^OO@~_u${n4zC"**r%12JpP}Pb.G?a#sz>=XvEpqPpR^|[+GO*^mhbF?fzp9=\vZ;=?^O<w:ySceat#&-7s!^mThU'l;~Y#.La~FH3RW!uV;{\I7U~GQ\DFhqxCSeUa#)@3o>N*e*~FGT-0uDSS3gx	N
<Nw>4Kzh+,'VjSj|V$cU.z.w=_
el7|&jLVtgMd0v2L>%1/B@jWTD=$#s5<,d=d6~TPw7jhjnH#i&VqgNwld:_.D^{CJ7[o"RxN%8Re"!VW5Udmk%;"uewKkS+wU1jIAA]-U]Q/aD"kf-.5A &<G&F4v@M@`?O|Wdb.[|9 qW\6zIKqReBGnSs"1[veZJ7+\OkEzpI@E9yj%</>Ei
-%Yz;vf3"N@s;l
cCTi9y!}jQ+E,`Km5a]])%tVqMzn>fM}5!
R M'LJf*S.CW[dtY]v{NFCB2pX7|m)/-wkNDK*POP,Aq@7U]6?uJ"hA2	*I7vF#Y*\hTaxgj,#KZ_	By[q$"$.{l`*rZd7$tdE;-K^jN5WvMf+1)zrJ\s6h/6/Qrb^x)qzE.O`;@ +QYWV3Ho36wB'2Zz DeUwGe PpE$	)rS&{bMX!4^U;:'JN_Q-bf,<|}7[:JpokI}3k-)98h.*Pno|9A_mo85OY	WU_Vs.goQ	hB5ck\E5mhi!1: 2Z.);@yEvD<Er~HosB <moPHbz56NsWIgx#CBA	xJb,\hp<FL,7	~]t%Q*$gX'\;W7CZdxZ
33z4wKdhMq
(jfg>f$}i^5S0Sn_Zjj#"MZEGkg6^#yW*!w pFf,,[I+cNh6`d8<IrbG( !ygn!.d_yh]!cFO	K+4K 3IE+T,p[5wpf+VnIIHMqz [Jbn\E\M5j[V%3zJvfY#&wp.Y	>YjTWC,GL[l#etF"&>w^jJ2u.,PBu]`v7&1FDee7<Etx#\lBG`,i#O^D_?aT%E<A"R9oy!MGA:~*DR+Z*d\Mh?Pl&;w#)qM]7j)S`ro>ztpA<8,Kx2@wM~?=:Zj2J".J!&|O|r~`x~tq;Y=WZ8$U)lFZaH>y(;KR:/\\fE.8/C|X	^lKPHC%:>8lBfG0WUM(u7B?SpEh2V!dRww\j?qww</3$],F,v4+\Sxj*OUS-hR%X%&%-EG{Gsp'Jy=G2":\+5lIBxbT<mK0?6VTl[FI4!Q=.a!mgS>?nOX=~0E6jXzMlVtySNJNpe$/YQw!&P#c	tDW'QPCuoc5
LcmprnqQJC_o$+r9=qU2U}y5qG48HL|2Uw6Z((~R!sa\	R,8-e'amCH45L@&(
(t#3,OLR3.=+'}];[d;
%FDA+Tt~LqtGmfx~EOX,E6nB}e0bM[!1#W7:cXx#Dh<
P,\RA3VbF}?0F[2:&*2=OK;vmDD_z]wGfmCev~7yP5@q[`Q7T"5a,Z/{%-3,?T=u&s##97_$SdDv"Pm8"xl'Q	UJ( q&rOS7uzR#E)
uj5_B)}$Woc8DhiHk6uCBqc5;ER!xxwj]8dKy_OP_n uo%kZZF"3e<YM+@	F6Y>hcD$dh|DKBvx`B43Zh^GlMxNB.AFZ_Pw<@q~A$ik2B4ID>nw5sZ$Lnyf&.&M_1VSt:Oz*rT0rNCf863Odl y	4/~mVU._#|us$u)8FG*;=P^$(bN1H6>8S[jZt mzLA?:VYYWx{}wIG3Wo0O7(B^. Bft)FLmsud3oxO*8tgA}51x%IC(S},Z/HjYCbA'>RW@H>7@cz<";J8Dk4x[054->YNyU	X43t
!VDj25B+n!+(ox_>Ka{.Hn\Hj=v}^H|Wnb#(j6)22ym[-$3nQ@k_Qi;vBEI/F"C/8u.1h 'yP6x_BTAkX<8m~P}>H5%Y	%XaF]A3BCs#\3C&IE_tQFU:;Tg
(x$L\XDU,P\hB	'<UG[`<U@oa.h:1=SNC#~90W8=*5W^1+z?=
K"ap7bC1*01su"?ueB4m,1XHMf#c7{,
z^8GA&i8O.8X:!R#*1yz^[m7|ynS	79X}8R}J;R"e]Y"?LR{&]]%^7jq~=;{S%js XxU(%-y4c & t9m8go\)N^UWh=DQ&
7u9m1b7o'SSZGiv G&tl9+GENIw#g(crg(p1,OYDMU+r}>#tbbi/wB*|L"cPygUgO|b~TV#D&{d@[M]Dz^bfeV<"4;TbYSh-ns@".u6n4d`=V7,Y9X{h}tm7s/IjoO}-$GF6RF"Oc&R$bDYuzi}oJLU|u||TUyD(:/4}Ymr!<gR[geXGb<!#U`eI:~u>Q(=?bf{C]Tp 4Ax>Wga WHh{>0`>U?)hp2-
C{"qYxC)}h_]P4/65f~"!</-d!~`M4g^&J"i:X@E\9^Q7?HA~
fLPsxH(Tv>&:90NLaS
ftIy$
(Tt'c{&1e,myx7$<LCYT
 <1>:_9yWkE[DL?	\eNrA^:-AE@T%8&Plne/=_"	2tA`i[soDd*nicl"sQ|]8e"5U}+RAU1DDlwl,](~bNK+rY}a+vS?#RQtPc)TJe62vK)#YP]CfgBTdBtS*;7OT0D/L?RJ91{lW/"n[+G	[.)*;<l?GF9\J&b~B!e&4nXv08%Q~;!]QI{@\[\O}]ocS~Nq[wKbxLx$F	Lfo)'Dw6o3aM9LY\1hXG^?{nD%OP11\gNgfc9#V_$	%1Z^	>id&!gMM><2gtl	9.LT$`TQ\OCRH>=bv|jf|[0$BMA[}~;'33G?UI?@}Nk+BhsnF?fEvZ0b#D$2jSUmuJnu+p`;:/qi	:N&=E""Gr@yT|X_]`7{i"a4~Dp06f]00:V&Ge_45\J)o'KY(oDo-?.T<@1UELp`\ |m`i%xCMan}NHH6n1}R9(<;4+aCz8J20	=`E*c{9fT39/QJ7[{Kc&cIb7&&Yl+;zaQidM>^T1=+>TL=6&Q.Ojwd{-S\C^915`kv4w~dZ[.#pBW$%,_I?&VCrzG(l'j0 "V3(ug'
	2}@Q&/gUKH{K38z*&4(Ye4wJ^U"|K=S6Uh}15akX&E\&y:D*F3Rd@JQ~Fl)u	eN3C=aMC[r>/mCQ$"U44c2FQZMP//1Ox)-pdr!8]#fwNnNG
j%yB`p+?o`tZ`mWLxy8*08Sv+6|q'Fd7x-h,KCUv!htN,\{\bkQM:]bxL[;j=dC++y@$-'+xUIP}g3Vtx'*$_~(@*Ajp=a<t:cO:8txN{;ET9jI!jq6n=Xy
l"J["is-en+!p|*X2()l[+95YuEM2!?fB*rUDM!uMj\u$s2<+^Rh"TwA^"SdR\gm
B"*`$	9CNopQ3d{gN/%f"k@W)dk\LScN)*1bhF?6oB)9{;B(~/{IGB'Nj?	>p$(	}{^ij>_*)E(Z^Bx9&@\3&F'#|>3ihb]2QwQX2> [~cKTPb3Kcs2;A|nA*,&~K>{wX6JW#/{#C%?!i28h/yS?8n}Q??)!<e@:)JFCd8dpEJqdAMB'+[rTO6Zy!>O@+>hjb/Tc`S&Ig #>TAF=\HpPWdhTKXdhXOCg~Xv0W^5q<H#v!CEP/Nc kTZXWLoAYJLr/kB?aSF7a{\a>GighXp3Oj}bW(78Etl\K0rEc	8%]*g=5TnK!|G j*8QJ*{Q3r
:5TvAiH/kv#xrS:tbU3#h#(rr)p<(?09)
D0i5Q%LAWGLE#saSm6 	a"%CJR7ft\$%Tj>E=I/QP9"f 6tM$D\zu*$/?}IeVV<!IURtRh"*v2n
9%ILi:X
F#-sjiPxW}|mF+UO-q/Ct%%	rKA!]K>t`#@>xm>)Hbs$2a]0$.Bj6*98
)<i kSd^F'ifAR4+nghMHpPRurlE< blRL>c[lv]al8/iU$y8q'-wv'1$j$sF8-x<[>|m)h%B$ikib~qr7W =7}EevsRwL/J:=YWb6$?DV9>1zM.F0g;kyvp7~)C.S-o;3z%N;Li_[+["-1k\RDUDB7q|<,A]5j+ATt5AX0cN@"uV>=]YfxhbxcGfXm*-X[DetI,/H%#a1edpLW+CsIw":H<szR:5|3N4UHFok2[v6{&9),v(6S8 w(L4yUB'(xAn=ViH]WxN6h! rHC[ys1L}=DE__9!Ee/YG`hoc9hMZ5juW",bNqvTWNj=Z~P1?{St+^fHw}$lG4oUZEqYJjlFc'GR3O3~|TpR3\rdR=I`{Ht+lUXl}z|fQ=JY3Rh7wCl'DB4C|HU&`7Sw7Q7tfhm,pEL^'@*F:xx{^,IunPz?e~$^a6*4e;[v3+]X_0Qvt F/RI]$2o-9-i3Q- W>_Tw}s	\F1\UWs)xa1D~\6P+tKN!hYc\C^&j_qxoqXMh_97J zA2'7pa)+J;dw!7yqgUOtHk#c=rsuN1z9MOl+~.yAta\lv]'np>y7_M
BmuM!st"gP8}T|<s@rwNJ(;s6[3F\][r&N^$B7St%[z4~)je&7pYs.7\98+vzaI^Jl;%>-ahkwZ^BLdZ~[0?|JK$jKAB1!IUk6ACJ}Y!sA"^i}'RM7:9rvHB0mAe<@#,f
+=zM-@]2+ODToH<`MrSt{}5dt$*0R
;A`Lc*17-.$1;h^HQ*L)zHyX@wfD].1.(NVt6j#6DUdT\W1[iTUMP#;7km\/P(9%*jC=o1!sr6	G&PD]34?QT}"}]kCkg(v~NzeTy[Qpgk(v}V-)"tD1Sk%Rkb;5qAH7q%FC)P^n.Bg(by8^4Sn/7ZAz))lG	I5"IV.r^Tw[+%}|lsm30mfx
>.\]
(bI}~y3c2)qvy/3QU
tq[u'eHsq	3E``]b}8QO5=\|T6Ra_ ~+p3{SSmP8/zJU5eP-if;e@7HH>z[Ch#{xQBFlX	Y%'_!]WX6P?-X-Qg%}wDf?hY*'CKx4>Vm`<lg2	eWe4^\	:^07X*7z%GD>%l)B/QB6N{@lI?K8`DQ-oZ<;?[J;dY{m[^P+U"pJY$zBA"=QD@~%csjO}(aTHNsF{zvrGKP?@|	u$n_uf)on[cT9(ZKU~^)}$OeirEPFJyTtW ysXT(t\-Wi6Trejj>,\l:9|k}[5T}
yE(OCvrUu2'3$&qNfc	h\}zPLLO+>
!,siY0Z,Pfy~F<`sWT+fEUO:ro=e5MuECVxsk0$pX:uzQ't(b|$L $Oi06pAUsj (s"XWfVbDW,] t?LeW&YOiNr=-$&V&_-|Fxz$\tQ{K6A*#%\GYt'Wpnq`3[pHoI
6=cfD#C(vP9tUK@</}*R-@.l("QL;*b9#Z,}t@*6M2)zDIb-cQ{0I@!x+![|TAi2;9Gnn;P)BHBU<sq
$T4_T^fXd"-=xlP2[!H|raiKr\GEAICYZ
O?0e\Jj5 J{&~C2Ag@'Um-8ST)U9[F\.'IiA:&S%"&MX.4fkWd7]&{mL%&-JDJJ},#wmY]shix*<Cl+JNlCk'F(v1vEwgUmo)56Yzp&Fh:zEMN(		U|MwKVb&=dXi@_hG36ebJ@t-]Z<iU5]y0%7uLaF/MHaCTY	-B6c4BtQ'5k	:E.|,e9nCX`c04'n!")3:pH=W^"L>v Gy@~J(LVlz!1!{sj$F`oxD.m@X=\8d`#f[kd//f
U`%~LsGB93>,egoX_a+!,QR>D<JuL%^'rVIEOWAT-xxW*(Bl%55-/25Zwwp3V?suX)4\Q]N<|m<w(0U2&%qVtkG"3o)Nz<f-k%%ibF%o/
M#&zR=2xGrPwl`;W(0F~^8\?B:bSjeN\&-~^j$1l!|],fg:ku\q])eMJQ-#_`e{Pfy&~YB$	(*\YqhPR&Ws8w`Wm!]yF
WA0=#.:i(qYk[N6v. Rvqm)Q!NREk9 5yzq^PB{?UI5_h1?uCYm/d[z/)Irk8V%\p4mMpmg>dWf>myY_e+LA&a/b*DP#2&sD`$D/b#ie8Rna"aW7A[tR|sGI@nc5.9no\*V/%,@i;8$9Jx(XZsowT"bwK9cE( &%SME<Ml9m	Jt8uP$KKLhzLfs3xv)8PCj*q#="Q$f.?iYpQH3-X0d%8(XVz@,zF1[+tT<V Sz1`W^^/:8##9W_+oGU5\\ZO0EI5~G&G
2.,B)WsY*b9= A	#;v'FHv\#w0Wxv|h1m=[A?YP3At0sJpzBw2bb[)7~sSsp5~J+uvE]t]5~f_C5m?vN7H)^vyJMp[-.8oy:\-FilJ_,*%%F&UYu>*iD{j*&K.1<x:^JeZ4f6|kCyuv=8<A$x1x1l'`
rZmk/>gZ|nR=v\Yx(n\`#qkUFT/y3/p+8)o`VT(MsQ9oPtq$K	 3'}8Zu|D
?L>2/3f;a6y+dO4X+s}oHDWP%_rrcy(8T%*8MHJK(z_{Ux23?onb1;~nexaS
3k}8QYjSBa8oeK33\f}XAeEJ"?u
x95Nu7;!R1yXi-k~=.-THF^g6!J?v
N;&?C/}2VV$+/o-`p9hP>\Qr5`S(vSP>3JDLG5"@*N_XPGtY?k5$t<^Ml]Qr7Kt-ANpO_z9IQ\d/ASo,',C!wyK`mtK;zC~Aj-h%MnFiv`la haEjar3jv_<pC`9})E>_M%[leXK6Pu956y"al';,nFi(+M;M3}M]<(ccoL4is rY"i!Aw5K~3z;rNG@'6O#ux~GAF_7MqRNeIvf|h|q)Ra"\`[
SaU5=)ZFB
azH[ceNSmM`XR>?7vsn.M	A
=!DS}P|Z}GkgqsV>Oi.>te'Sso<4l2I8+{^R#gVGF;O,iS
Ls;:p>H4p]8p&&L@9 #E$sZqw*+P'D s3>FAFT']/T=bgn6%"6`OQKvEy^F	pP3[UcvYH&sK_uPILw#wlApb{9!#+qbAh5mm]4PgWd
K1#h0s~`X	Z\V:`/<3QRr^z.bRB$ZR%m%7F/`V;&`1FSYO@S7e@7P{d1s
z;W9RVb#]VVd0,1e>L_5R3s}d*:tM?.3v~O\+",]d`scV3)~kd*AOboXQ/#=4dY,u]iR'z?645lHq7=iDxc!qm{8T ;B,sj)uI\V&y57%=tA7,&we#PIXzCk(ZP!OW`:x:Fj~.FVM|0&-(e%D9ct$<[A\cJ7+x_coql8$w@`p~('9=cul^z5WI&$sx#@	,1/YoQ=6Q]nZhEA9O*'>+z2Mzf'XOen^4rYHJ/+{lHL|8y/ybI	5R[.SfUG+"N5k\dL2<Ar4.UyN`dp
HeJ=$u|Q%4RGh3;Q-gwG:A>L	s^s}}B)7.4}ty>uKd-/*"DF\aru#JQtq\(E;{IApm<&~/ZC[3l	?Z_
9Al)DzreMwX(t:ki'\YcqY(bw`{82j@k?&W8*eZS/^E	2D=;f(ZiA~j
=20Dali]>s=H0I&`E}b8>. -T YcE`$bU\jiyi^%G@fP|K~j3JiLDF^#(;ZZY	6f53#,XT	$x"0J~&|O*DlgZwLPk,qcF{sE#yNg(B0FNwnLQiq~>^cI7ig3hZe7Vca|oA-to~Ik2cun=/jl$)y9y${2pW.Yri+ZBP
P!k+cj0,-O:H3{<+hpVu"E$%IGR"AmcdBe?_Eo_q1T)Xsa0b>}on`_xL+uQti(qDB	EF{8"Ii.@%]M.W[kM#(`3x[s^6Yr\iWTX4t56Ex+6\RIv$y\6lKl[22-KG`zAII(MFhPgv
P@qt09V^S")Ll)&JMmn]$zsJ(iKPY<!bMC@J$svQn<GY;DwfTC9NQ~UCc8B=%+TTq]4@;M7hiYGH{J46<_eO2+}a{"Z(m,p43v8H6^JmBI:uGfXArYXF-P%tT"<_iuii*mG|%7|IweT{3GBe/FdF?.L"~.KoqS;cx|o>s2bFn+bcya^YJQ'X<
$7*RHGK!"S(JEYyxms1uPtG,"a@	pg_H4+fGCJ'=()'SRY!rSnWo]nkl]-oQmf8fSJf}dOvEiYM#l_1V{Cua}s"nn).\Cf	c>eOz]YD[{-p'R.`#KVtV$c=mDLq-D0mqf(HPNN`:Wl@K!/gY%s}i+gmlLuSO{tB./,2rCnqJVc}0Y__=hL9Ml*K_Qf(I34	kTCV7l8x[#tIHj!8_}w$'%],i'qBKOtA B;r"~-)@oD@"sUpOU@dZt3I%M((j+O1b4-`e4>21-Ox@/4cLZgTBf(9?jI4w1YG!0g3]N5J(`$jdA]U4YVkZVecImwbu'F_+k5,6zj,>jZ9uk>g'.H{V##Xy=>}r18Metg|.N@wY>"$r-{tq\poz0f<W["UM'+H[Iz&xy#f3+253.4[CFFUn"85\|Yh>Jjkdm>g(U7]em7PSu).EBQeEJ0503/*+V^1:e+]P>,inDX$tcH:'6Zz'2xA/ab5x9?Gc}lYdJ?Zx}4Bmu2@UeT*H}xBbB|/,Z	QgE,>mIH..<5V9 J`oMs,JG# 3*bIf(hN(l!<4GS`%HemYl%1tg	J<3<#%C?4"J|&DYu^}"RY\@=u84"DUto&`L/<<{6A6,<gYAB-$E0tEixuV)\I4zj4F0b^UVD[I3DK6m0#rf3Gv>\7j@M={E]=t'"
\^lxYYk'd}wT=5Xm9$D:DX<LD[u]jCs.M/U}QV?f,7GYB,v'^l$E	]Ib?k9Xh+79?6G++*}?$S+_BJ"AQ@MyzHH%GdWFt7Ek-	rn$9~.Cx{L/FIB=rVfNJUng[HF[}jrzwr5>Smt0rF!2;u$}tOuw1w,7]83g{C}$ZGe:S,x:-LcC7WnGm5l-3E1vxW$1hN;C#v4{k<~:7EP0e"e82X^rq91.jxEc)ui^t#A-slAtk;7"6?v!?v!j$AxfO2|J6peL"x]6DtbMA*tCo"%nCNbV,ySA/PlFp\`AgePdv}$B.WO5O(&T@ZqkNrqu8&`Fvv(KnZO5-pB7>Fi!8kaU)+gM<2%Yz#/.K+nUT*}JZ;S0'ju6BA()zFyvKi'm<F'r>4W#J!l>NhWG'B9\26]D?.r93Llp'=CWHD"OA7-2R=aeGX6qEi~>TW.-e	]_,5pcF+W{_L")e}
XV#{~adHVu>l#fxW,?)]Pjq>01@{26{z>,"|+YCBta6$3k`RjT
;nk"">g=W\z+Yirx=T{W`3gpBIU-4Z04L;tDohdGem4W/G9[].!`twZ_A^NpZgd!'v:^BLhe7<h]X.mNnI_`f&$&f:njWzE]j\H+}c)L!i}WTG4SvUsnRhC=O[4|~az1).-r0<TU~O:p2U'mWmBM4lXl%_gClS40EvdfX$\*tB!(A9^{BqYv7}-br	}Fas"m|~r
B4Z$d=.9O[qd93p2[dnJ/m:F$p3P~MSs	qu7|xY-.=K1\|8+Ou/N
db%O&~EKZ0(vuzB	[0Au:?Qg\ZoxBRJl6#S:Dgx8+>t9ziz!QNt0nIuzDC^sG=+G=v)?L;;|BIuV	~)^nrO+Y3N|O1/)p>H2+5Bo7t!"z!"3B\XCY].vt_[&
^>-@w!a[wfzd`pKeS-rg(i7	>t$$.>|@8x;=.jSh77#N?D_E;QxuY#JNZQGmhtVL&XUrehze$$R	bxX9Yeg?#Y(rnq}CT)
V?nku?P>Em"K;[[Xk~isL98`^^}Dc6aE#D?F&}r?7jETIw1	n.+0A0O%`&aY*
wl-d2PbiBsM,TVt,`XogGRNRK~,Ns4R{O>ZPO&s`$sUK'nH<+Phu\U+p<RVfLL*E*dqNV)Ty8}V_^7G_3E9{/-\3;-[{AAH^(zL{8:Q8$}UPqoXVSF$C>A9%Lea3gXKb@vRFLHPk;
Aq"zghBa$HN0Vw;L6HVX1fb[;I}%e2}}!^/u?>mh/VLDb1!WM>)elE!"H3\Bkdk2T
U9o0&7Ze(/qR]r:aHdO?a(GdJ6QJ&
v`'?cEZXcmrN#zan70\4kut0)0StAN-tciBuM[o"^!9O^160:q`OkKnqK`Wm-SM2F|HfKB:dkoT8~77Z.7d{Qm_*JskxG*Bn('
YpP057_fVjmff@nLAYj%]~ 5Pb&udo!/y'j8XB5|K:hn*G`Z?WprIO:wNoR;6m<iBRPYtGsG*56Yurj:[Suo<fkG	jM$O?|oCf;6&u<1`w~.O5'U}C:8;7j?%z9ZdXUQA6Q;eJ	\WWEIs,hZE}TNzlxjyZ
nF"TEUv?2+%7AP YC8zahG{|_kv3xNr\&&AEX1C'MzH\\mNvd*RIV)#|`8Oc54rvg7CFC4z'+J{x?Zc51S]ddnd:VqlF|GiQD{\jlm!s[._Ol]$"v^nb

{JhH/_QK1YaXB5fg9@P^hXyPU
}O'5Z@3O&r/l&#qH;!?vo5V<z&}we]LAY8`Txp@O%a4S+g)`gn*-oMqKJ A?2+&&'gbv=}4_jpA}B"&%7_\'*+~k7V6ibbfFkTAhrck1}j[{NVF<G'4oc#BH#	P@|m#	Kqjkq|'Qgn:z5nUbj*\Va&6{0"Vo~0c3`2U'\c\svSHCpdr 1kbh&F2PU$ip'M`=8,j@O&[F4\Q!}UO{iC9YEv'o<0B+Z3\%hu=LmgWmi+=q8JG&kdE+.wWOa:Gtk_[>_9twzQ~iSa3^x(#9t\1*(mGDQ0F<lg6[]@@zb}Z+ Ml~O{'9_4h,;.IcVB2TY&l[-Lq0FZ^F>v?.s]4P55q/l7GsJg%-%v>WQe6Nyzf3BzbevNj[o9D!{D?7EK@+Bl?wB'|Ddp%#+EiuB,O.I[a%<HIK*<aPNlx$8:[@C.i Sw s-VUqC*,3"#0#]80?w4PB(Z^*la`71'M<z)
}RjpDh,\I@(w%Bm)PZzO0]38,N"RzElFHf&zux7J-\f2mgTUU@XA@8?fDW4NBl5dHb@nW=Tf!')M]3PQ-DzF +	9P~X{;~>b/gV5Fcyi'@b[hiR1F*Pfns0}}kcMM))^]"WHi2!g-2;yvDry&WhF)VuR;:T#M3a+e6I(}"nlY>Ja;/-jS: Mq$+8jV2jVD)HXD
p	3s{#WmPxW
m'6U{!9EDEjSRGbFTHj+;k+@m7"0v1:b=d_8/TI{,',u_pqn7Ye}O[-,kx6NJ,>v]*)";en.E{8Q\sIm#Q"Ad=]%fL{Z8BlVF<os$uh)/hL#z#,tp<,(ZG"1t
,}1,R} m'E`q^mrzud%uD-a_a~^"Ig96SerwZp=Rab.1(Ls_0aSUx_-86:7CL"{m{`X2=b:;4'#
X`qnkwTk6C"(/*G$; Db/^N#* ^CiPQ/*+:;U{:_jk3N~E;8:lH4Tw}[5cns]%=Nqky\0V;&51zGR<jV/ZBya0XE5NhCUhx@X	]h/h,W;](Ux"F+-,L#F7zg,"5*~RC*C>`^Ai^@b@hEj|lDyZn~bgY>oh;XVb[<..gAS<gH.C;=9l,LqUIQ<wA0FR3</\b#2t3<{TLMhKRs>FKrp}U|+KNiiv.5$:?jG>W2;tc=T)<	-( iqT_e;'CIl|/,X!&|q7X4X[wner$v?,'Kz2ZyR6jf
VA)HU,IQe_HZiZ?i)ZF
oqhU+yubg&MG"W)\pja791'"d+%iC-"1t.Ls.x"]+]	"jK!.i'(O^ZnC>|b.{B}}D[U[WW1b+C[
1z2!NRs2Ez7p%3{e!8eSK*YB	UPp!XsA+%h;xn[7G,iHN!s&	
,BGnvzb8)Zv+C\[nvx9j;}c'hWvsc;_VT[|b6f :^AnIHUY|d_(8Lc\Hc22uHWrC15E,o>g^$l)nd*[Y/da;@$1Cr+<\{zB`{7e]+:sBrl.9|'f}ty&=ejid]DT3Gd1QY4z!/(|(Zl}&H\6,|#),?RK-->e%E&iImO`{3J?zf"PLvN!z>"1/u9=\P/6b?Gr7N_6D@}%`-=lPhNq `2uNN`9V>y>+qS*b{i*@5/O$Krw^6U3|};F(v+nW1*XLP2S.w.RcuKFq&L)KJ9!@_Wu1-IcnQo\LuP+sdY;_>`Xw!Mfg$7AZ{Z`)p+k;6/v5w2~'h5IrGE&;$L$N5Zqq"Fvddd_v8;kOjm0~ek-}z|GUk:|A=U4h4tP|.n)ca3Z"2*<pHS7LnF^/G4n"]s=#sUvo5x5`7.S`f2}1J0]x*-^G"2&bVf&(QOn'<R1dhRT]'FeQNlqAzR1oz?f#ba4yjF@Bmto#aFy=+G	wDf{6,+bD@.mXH c1W
7HZvW`#.ej&+OS	+$33t@>RBn:["8lJ@]v&qrF)f-=^@Kda<kB6N={S64q"Co5T
uaY84LjC6$qyB;p9?g'yYN67r$OJ!u(l^s/84[O_Sl{NgeUC``AV@'ouL=hG)sm(g71#*y0e2""<J+|HfVCc\ HH[& vE?QR%1`Ij\mZLZtE`P\R20*GD%$'6P2cffh4_:C;E_sJGjn$d"mo?7Q/^$`$`"p$[i+5jE*9hBU!x`+=nYB36Zg-.[}X?pU7oI$5/B:U=^N&/Nq;z^ZG BJ{)Vu_;QyQ."Aby-d<<d~F\|~&VnLmWR_OmGo7e1q+8. gL=Dp}^Z^MIOslRmAf-J3J>Hh({24<>|R*1YpJ`V]lMEJ1yC&(V%&TenMn_Oz"Kfi{]0GLTto|y%hr `r{dHGSwPZVp.{
r&r%O-mhNoZu$'$IZ""3mt/(buipafr*a'I4v&`T)?=)~g
KgGW8
x(BV@^#HkLeoj :%x984fX25rm?f-N_DTr3Zw)>C.\S$EIA'>	h6>xSjbVkM*Yf?zM	JG>+1/NpfZ=n8&ENAA*;6/8\p1{Cnd_);P'%!*RbqR?/=<CsW]#}X>{mp;zxlhu`>#5(P*6s?)wFJ2]Kz`|unG:.'Ue,1D6XV1^7pZhEu/6e&*t\^
u0XTX##1h>#DPi;SlS6&-_[pKo,~)PMI3@Gti$UC!3R5 5	m}z3!*]N-5oPa8]4.~Ia#4kytL.P][7-O/_T]<j f9Qg
8[B;oP*Q3cicIv6w+cw}^CE^fDQ;l>C#FmzLAQyy=i &goO)	wtJ!4..$8!&&j?e`&EzCHZ4Pbc~V:Nm4LVF,Kd|f?-[l`A{W;m9-U43R9;RW8VuV-m^<9`'H5l?RO^{@\%^n4NO^K&U&t=@tR:9V~u%0jcOni PUVn7^f891Ij.&eLj0b<A1bw! 9ye$S)E+:cIvp6BF,i+:?6uy{o2;3-b
wg;$nUeCwkF/#W_q&dY,:U"5R&;]7l"|8J5x*T>Q8bA-f+ok4~.:CRc_bi9FhmOOb;rsfKW"%|' x4CJ$p$D+wab"ARBeDY'b56%YhV"iBj4V0uA[}s+Km=S6N"y\Ovi=7&:Hrc)'["?,=q/bYn(SM5PyYj3(-}<lm:{<8U3n&R9cn(g=?fyxxO+N!!j5rV`5pxqFcZYu@5~C;ho)+*8KF^Xv.@V<Z3
mp0&HJaVv16:4fw-+	&7^m=5]d':(TmhLv[k$O]'-axvFK]NIz1Zh K2WKTkZ[CDL}	BBI\p
	r D7csK>r9kJdD96JI~'H8V\"KTZMkO?fBO9W]-$?sY=:,F3C;$Wc(zdR-X4@bacWQ?-[6"`Ra401YqmmT'vE:0S %}'u?tQae(bXG;6#^0m5ddQ ^nCQFhs:p^A0EV%>m+JBe1L:R=M4kV094qS2Y:8	znXcnc~!NOJ9oYo/TVS{v,1OVOx?4Dw}EgCxUz26_%gW"!qM	}eE$b;`lL	UwHL.YD<"h0Hk`gz+z@&<f{a\)(Bi|_@Q
wK_KU-$B(@ x`6UzAbEq_4();mKE"zX+SjfE>%bwwp@-bobsgsv-.KW`	;ZJD)|cy&Z,I-kh~MY+wBJ;$8)jBz #6x@K'O2c3VG`K7jUJlGK(^oFOOJG[.;64^arL/[Y4{*fB-~x"gd9j%0Hyn
IupEI=+Jk|J`lWw<(6.YOq\O!}-sB`KX,u7cYfT2( !bKK>!of2$t}Pn+lUa9tX]ioT^MWfc?qsId'+\pMh78C8Fc[TXy90#^o/tHgtWpf/[u3II8o2~7'&V~ TNmwqB.9(,'EL7$duK8$OYe`#>i_^h=OIniJISoqI8sjgLpa@b1OiL >l-T=7ZAEq#O({!HH%kFr':d57rn%wgA$2s'D1BQnSQ_b()_Om+&1k3tLd:G.Ms{N=ag[Q6'ASR*w)ZlFlYw.O-!Td>8!)jjY0_De
~2}+cBa[kD87HDz`4lcy"Y%{\gu*-N+0=e"jU5bsVdW\A}pV\p^Od2y"yhF4AIW<*Xa;*=>uOJo=a.g6ED08{]3tKP7dOlF'<kc%L"+0{%A.ssaI+..a*[TT}3xtn_yT>x9@$Z;;/{ Z?18rkNQ^,"N@z rc5g%*4peg@V:_0HtEXwAD*%8L,#^~e<=N)WNOU-.&iF2sj.miMhB;aL3b:>o$B5&JxeWQtFjS{pOmd-?xN&JRlc\^bO}x;i6CR(n]5IXp=hg@LjX6)
J}qbaVG|}YS3dl) 0{!+Q}7v5^l}CY]{2;C|c%=8)"$f?f"#YwxJy>Gdd"F;7Ie;i#v}yPS@an5&q<O_ETF_UQitgL*-xI=F\u_SlK3/}
l)'1?$1'P*B`UUbbLG`#GM!z7'rnAN;4> n@AAQ)l-/f~]`=2M.4'v"&GszegD$WgBrgGODG*ZXk&-hL:B f*`,Z|&OyiaqJ*4NyK|Chu4}R.K/_|P?&fc6F_6n38#eU6!)E|>AY6wh$0jj~)O#VOGA9^sueT;SST'a
Y5NI K;\nE}-FWDXVt?0m7`nG+}mmAa ){=&?ehQQ|2\,mWEhO.C!ePp	y$2tX.CmsA1Tb4_b>vp>byb@=l1H:HQ
n&xOt)d~D=E?\*cGAy)^d}`1\5yk[H5S{-3^_IxXzu+4N)jd-/r`ZMeP#V>2iy]Nu8w.Y[Q9J7YG1Xi0/mof4(~, nC]%MQ&LuSUCQnNLUJ]9bAgtM.eRB6\KcqCrV2e (4,56C3Ja:&o$8&L^aL{iv`b*|uo`.uDtwuxB5/<K/,;gnV[R"d.v-(iglu}NZ:n)A>^\="fVdeeZ4Y5Cwx<2v$N)$;()*:COmJgw#ym &"@c+c/vGn~0T7byq;e(VSuRUS1@/XCs%D@lDRQ1@$`(.Y$UAD'U{f7luI"$
lgP/X4&K`hyevev,Fx#b.opd3
slc4g/gBIE%3V?uJ*q[I\VRE0Ecuu&gh!\l|zc;R6Ak&!ALrm4F]p")P/Qyn!t!:g+:o?IP	sK+[ss7X3FZu}VC[hk=BSL_uWB8z<Iag]#2=(>Kz&`7o|)g{fN\JtByE|3qT4~(0
%&mz3s{QjKDpR|g!6XK.g/[${o!{B3wxdY\,x:.jW.>Ah-|mE\c1LmN(0 bgGpzV~YkHC'6$4l}}
qn
0hxh@f/4iOe^]Mgr#Yq+fX~STCM	/6'T`D>HO))$<RsUatjiW	p7F&n5c9!{}et^Gso:kh,taMh8R#/<@f-h^Z?Ov=aTbFoe3*0p5>t>pa!P+Hg,dCs(Y*DP4lMw~n0I=d\I7Vc!pH1Uf#9zRBcx>YzD$d/GZ*
hPRp%k}UI03Tppu[.!!u`14?XW_V#72cobCRz9l3$'egH\Qwmt=Ky>a2iq\ndk
E,
(Gz|]4GVR	3Yc)G}~yZ\,y#o4d{7@j,a;Ra;rWm$DjDgpMA<Tq#N-y!t\Jr c/^[=}2BjF7
><h&-Q=	r4U
q-;T5vqo-hVWBN}<]]6Y6m*FfPq~Rbu) "mg2}Oo<F6`G-9#e-`FvrIo8"!u[pThhL,KT^]_]_,Q7@-07yW6oYa.&E"g=*ek^7k2e@0]Hz$P7)>_?b.jp.(9tDee{
#.,gEBqHdS~^YrQ=sZNDkLEsv+JTx>}~~+IlQolhJV5;9HbePV~|d	0X1O~.VS#{)BAN-;#|V*xn?L.he%.$
,%z{/q4O>oS\>[BZVHi%D$PPAR&aVFT:'G4'*{^3&sQaX"ISFE9LDZOZYn/JYV5#(">.a]aSI_*]Umr$M*fJ@[/pL<="X*JBJE@_Mf*BOO\><~V8P
N~KL308[q#e	/{!THBp2t:aV]tQXh#B9@.o3QjX_*Op5)QDjx|;(*z2$UZz9BQZBj#
:T2ZMu`6*GhDvGVH,v4A<!wU{kj&
:INa$b4xG	F$Bj!BXBMvR'l]z\QDFQ,jke5L>^-inNX`{/9kJvqC2.^_:n8IEp jG-c~*t%i*.<QZhy(Tql4x`'[;dDGGO#g14}lt3OvhD!,,o@K/F}kyg/GT.dd=dzka970'HGkAG[h06hTAfQ"\V0-oX	(d9,R{)OBx.I7YzQA.]2MC{+=_m(5t1>T\gULL:Yx\sTyI<:67^HHJ~l_(dHd-*Z,(}XKuJy=i+/|^/#F~7~![nKq9rKym-DW	e-@OH |b
>dhoo]
qws)A-c
o{VL;M!h'Hh,>RrJn\0KMka3LcmMS`!1p+>!%E.4]?i~WmF)4
Md'WD3P?=5}*; )cjgW6gBdwDza"I{:|d- 5JMYb68BL,\v'P$2,7 P#aKQAmC!2..@rwz{=U	?0"#UiQIUZ3\_d:.`|NoIXsq_
< YUqP{\#OehMUPV8BhZ3]jyFV~C|K*~TE`>Uh]n3~f]10w@hkc>`%[nU6},WTL`tE	N<]:sDdcdo=pQq1[H*X7-8%ixxj/sq]EbyO3ShNkk[#G@-4>ui2s\S&=PoR5E_6HIa3U4~F@xe6!pWfsu>+8~T@f|m|7>Co[h&^
-OnggG 	9&5&|^Opmq*E^Yj#)u7}17c4@0Y%tEe@EH(.\3lmgtt5OdArDBH.xutyEr	+=g<MICnq3Mx?>P8C3zc]Q$Ru<W8SA!hgnWVkmw?o=0x)mtRC^U<k&WW#3V1Uj 37RI1[jO[@m,S+ni
\ :$I#q&z<k'/?gkM)Rvx)i5Rn$KFl)obC0/<}$IORq{hAQYY$%[`cQ^dmc9/2z_ycG05\V#o7NZ'5Z|A$z?~Ws1P9n)y#A1pQ.`zoy/b'	DKrG)F&~;3E:rU1W8][0e[6489]E[HZ53~wOq@V\KrIz7%q+wO}S-"7yF[ZjU~}%TbO*i 2	L/6VIY!S*M/?ZDmBbo_\e!j~ lE#G>{Nw*:|o/wUbv*v=JwHcZ8R&HPs.z0swmg%hY:)v#QL9QE1Ry_4^3x='0
pvMJ
tjL'N{] s^&+z8GA9HM$t?h7z0,#C>`rv)	w8oA$S>?#0?]X_|vp`I8W`svNqs"eX4. <Iby~\[<xC!=*%;5eRGeyE)o^vSevJPKxT6mg&6V,Z!T-dCOcolZbsakzTqY*wj"LDEO!\+vnYqVG>Jf%mKB``kpn#1Tc:N#c"ve*4Ov[E1LQ*/z"Q.U*:jl?dtm;^T3w1B?b!k:_>Y>3_|YHSqZ(>`4Rr($/&pklHR=QxrS'`sPJ8QL5hX pom?T&mll^,YdES,B!&N5oX2lv%@U"iUKABhToGF@N`.~K3(GF&K
W%~a5!xv'-r"RYC7]	cu'8P(RUmA"^K	aWyF\`.l{6wRvh0dtI}EBFNXA:#2w3:>NHJuc$bpuo9.aD	K6*0
1i<:+KU7K.I_Pf1eL%fAsSWeb-suyd	z^fw5oBY.w7CkXxjI-h4dhZp},1RIyw-$"G;!*9Erl*=t,c=	_><LUkfiLh'E'b#RTo_r8O]"xYLczG$rClBnLLQNP0L>[*wf?A.%|biQ;<[]`(Y9?O"T6-c~Wc>c<Dp>OrI%LoQ8C=/\XYnz#t)Gs]Sah2>qI=R"4U+pyOD~FG6E^II@:	1ijpSwz,
AZQ!~m)WaZJ/hpIQz{@tfhO^dTxWd>b)FQ$seiGC!J >V3J^&?G[GQhMeQHf!GnqK @Q~dh}LdwibF]Z"@<c]rCBe
'j<0nUw8/4{eqnCp,EjUdpR#~,6Ki|h@[43[se[G0=0v03)lj'sKp" E#fvWdO%V6:yrcbJpx5rG)q}!$g%\b=MRQkl\*()']EJgKY~6W;5($94]co;x9Z{l@R]7j,4R(~)ub`C]_wTC-+J;U-M0cHvk!$ {r2>"U*n!ZOZ7$<x,9mz^Fh!D}F.s*tY+4w1bl~_~I/_cMC'#i'wOwQM)]_1<r8Xm0eD.#kQw?5.df+Cmae(Ws8;5$FL{ ]J/Aq?[]S+Qp \1`L
d(P2I2s#R2]pWDdk`w_v@O3&.3Ji)k`w|Hx]f:>^F|<O+)f *#&)Vf \;_Ch!TBAM`;W1f9iu?*&`~r1Xq;e]MRa23h*(?%3aPe`\r7D)+%89	j3'+AFkh5_zbLHu?ar_(vztrX`z!'\+$@I(i'A\B!
IX=TMWciJUam\DDVZy1|0Z@e;q'd|X\wWP{aLbV0SmyDgu__/~O:u8],%6;:%6K@Q}w>5Cv;t{z#\LQj%|)J~3k=L*N#'{Las,yT=t6iy1M+P^xnc6d}de !Bf=a-g%_!T%-3	*08?;kYhgVmd'W8yzxMP
9ZleuzJ(5YglvYnN3=,!S<qSl&+[?e.qq=6&fQ].'=))~r7yXkX(Ox4:pNL8C#f$F|<uSPS1C[Sx#MwD})V3%^4|nX:$setC-\gMiPDL,I(}d,eN7t"u+EZX<Q-)BTv;ZYE%/\9T+%?7VAYM6#XvP=MFhjP`zj4Iwvy&%B,:Z^3qagXPZ"c!	f#Us'8_ZJY?!Hw x&}o
I\ju{.2(gX[wH,&lh!/0H;{z@)~S"!y)fxWZ`<IA.S)gQwSJY$o$#BSXC6z>%7epPy<J15JnlpMKG:"WhQ#/*cC6gp8`c
;SKt2,:*Lvy>`uyfSvZ'Duw{ZR#%.<Re,vm*nDG;%zAeLGl3@[;={?]}p]4vQY_HK>?Ng<p_+uT9{K(C}@< KM7PX>T$cA?sQm
)\{'Iu.:tHvCX%k
-V\%\bIg"~p$B^7!2dzJVt+!j[nzx<dz%n7k:*rdK9=!W0/^$YuD)B1JAs;	Rsyr?I{ClX>0``z9F<ME$hNrCCtf<xHiV51BFevFq^w~@UxmVc9&mK=rT{lp&}7v|xL*xft#PGUSxCO`
8"Gh^)-TESiUAX%_,xewk7YiM|'K-kl'T#,tSwUT@hR-xiBnbG2UGYa-~FSFsuFI38g[^TCx)|7'Ig
e<l{;*	(%L<uI{tuA-xI:NN~E.X}{^/j+lwbu]b_t{MYt^5N#illv5NAO{4)CTfC>GF{?)YrnWQfg<8YDQR6-d,F^*{dq"t[(8{%D7#|gxH#?vcUv.LxinGg9{(QJ$p	EV7C2D6|6F{#48`I!MDy=?k|.-A^c73E.3nLa*pSn`0j)N#?#cg}-M!(sko%dvoD7 X7g(Rv*dDKvmIH0bO-]-
ZJFOqI%fYw]2/do%;{B~C.J~BKIME85*,z/q@Z_"&cZpTGmusEG*Nhi.::7C7N5i0:B
Ci~{k'^c?m!sGpZX>PYS!SxyRp?Nw!I4qI3g0'Pn(}vR7/1o>G[mATnhi|:cO$@.TKXOYQ#bX$JH+NppCvz5Rc;\vk"M/t=,Ed(@?sLNI_MhzlW#iuKQ$i:$ZU&7_N"4*}RA31//#zQa*_o0OzV,3Z	ats!;zLo%fdiHHA}d.(,UZ=BQ/:,GxWmQ4ol-2bz6IJs	6oM2Ik,	40Mw3M1^aV&d7F?pA53vk/+ ,Mmsd%o"/N0exk^gIR}MBhR_a]C`[N|"sL5)wJQs9r dL{+N#R-(fG
zq}q@?=_1g|XD?BlqCJ@zKH>m1p+e8^_YV
W4!Tk~L0L1mT?ay[}@w /	Fx9$Aj|\Yv#nddr*+StFGP\/r^'H`Zco%V'OXT`4:{X\I%kD	p$St;m^4mc;yflPtLq0'hu	|Es=l"ieW9M	sQ9V2}ez>]:j*xyeu[ctB9MW-sANsHQeM0F\U}XpxE+bj$e~]2(zT\na:RyuG~BM[ 
G`T";Bq*w v4B}L!d/0B8UZGg7.S-Na>9^4i_[_u}L9C.])Nw6>QsW {uDoj$,]vi+#cg)ko^y*`3VaC5)_bkiEqel_q+Ddq!
60=roDiZT-oz;-=pWAJOk=+Vls+Yhr{w#%Ku/_hgz#lTXU#49	O+(5OYovN4Y[7Vc;`pDc/nYAb-ImZj?_c*k?G'x!yc\IAzDxO{OVcl$Wo?
2B4	@t[c`-9cQPN=o(*2`?vu%CSll\W+K1"wwL6gdrO%O3*D0;aE`s9T]^~r#^yU18"x}&yC8:p+BARnx090V|{bDG%gz0.S76kO'K3
C90ZF!kQ*I:g,T&[;;EXkR0dW+#*%Nv:24)iQZ-\IA})#b}48KgZH+sit3'|ES 'pXI7gLOk9^J\S#7u@5xC*Gdo=bEM[!J<r"uMrWjb]U"W4XET0x56"+Dt{m*mx0(ReHeQm#X=Kw?A(#*dc9]`X=iV,nucY(PuW"nb"5mkW.kji?dDQJ`,6P\m]3c4c/\wR*+Eht_b=VvONMI	^!Aw&(t_x0c\L2R,!*"v.NbjzMTmN011	r~@a]nZ5H$|XP[^0e&B{7%hs8~8IeU*1X6<+ 9_<m[KQr32JF;`aA-	S*!,1eFlRPgU?('.ii8]`>?^@Lq<cvLT`mp2V
<N"e~?e[,8bQ0>ur}fu=.K6Xo]\
<2kL;z9|FF"mcmJYhg1{L8t6&zR*MOq>(:4CufWdQnb.CpW$PqQU`PE@Im[JkIx4DJ7nq_Rk	RLp Bx%#XjL0}]3V[6szp=*H`V23	f=oz2%Hn<ww'dK 3)|-;N/[ImB8j6#&rGv)d*+/N!M*OBU+`E@V PwYO/aQ7i"3rlrO0d22T|,PqB[%Yf0t1k/TA
,<R*)u%>k#0QD2Xmy>@{7s~6Yg.jq)'d/ls6gk?{S*t@bUXG,_e=j3Zvm2[
`yeP@zT5c:0]+SPQP?b0-1f[G5}ZlNjPtJR{f1:k")j@T=&izz
c**Au*JQI1wc$J%b}'R.{yhk04~\8n_IbH'$0|Guy#7sY|Q[^`K4+[-IC-
o:C^m aiX	?#%T[\z50<BC%,"N^F))wBe=~68v4D*rAHL	^_6$}%c	azpVQ~b'aiPr2>}*K5tw^	k&(Q,.o3	j|`@qp0:|<%NzAL7xMp94Aiti~bmhbT^h['>pyX(D{6;La!V80?;b0EP_O e\}{7RVM8'abI	ih}$WfS':_%Oe{|lldHiFi_2G/1dbg5'n{y$>Gax'2g\NUXtM'6EcKFMWX@HHy/E\UNl|-"T319	Jtu84;=A4szxf.ww *HB)>A5^pGy|sHr:qM*Q)nI#UNC3E^*4/|?m|[G-^-WLo:_u5N7UAfJ4eLT?/\8<2wy
{#6;ycF7};St]$$^A$L&U^Q+ZNy/A3[UW
@.B1wN^hUS\H{|6K|VZXT-	,e~HI>#)v;t21K*j	d&(={mI"S r)j6)7Y	K9d{9gYX~:Qkg5\$ph;Q{E3F+D$U-wl:;VI,V$[b[#^)%chQN\7QDUc~x@I5/%n0<2fi_1G+6={)07NHmPTA(vX}H?rQ28"bz_\KU{_{RK>}rJOZ(&bbRP|t9ZT.S`bnqlH.\DqF<@l@>Y sb.egy[ppBWpI(Lv<c<j^*LmDAZ{w2fAav7"9X[J	7rOt\ga pda0?\h73=E@I~G{x6
2Uo4DO)D=)$&U!e3;")#VvC\Ao=pV!K1f;"0moym5j9b]d\ 0^>iATbj_JyY=)BVLD*w@)P1 WGE&VX(wdo{_+IfyH,;'fUBZ*,@0Y.#8wdJ=tB]gx(gI&e'6(Ni,~U-}-!ii.wwt	f~Nhd">x7yWQn13'(A^!Ay=p%0Prdt-;Rj=j31zxroK&dld['`I+@Yd$@F\QyL*gmG|n v=**__B	*,:vYO:Ny52fW^t/CJ6]{Ae42,7#;rj[mykgtuopB=sFvf8vltT>@^@Q:pW?MmW>1eL[bk& Npb$JsvXTXYDkMso\.b3e,wGuuL:JKmNY0r|VB[&dH6AJ5^KyW:6;tSg{Z2G9fKTRv?aVJ)W?A3=!,{g__z7_qo=91I4usaIX;9)kW6CTQw}mE_o&:q&p~imHec%#uy6\4lD%KxB	_@0gd-8Idva=a3]IPnhB^aY1+N4163L==!3G6_7	JMq&2'O/OgT/r1+h_/m0g0w/E"Pw-}*hbi@rT&{_9vSwzv>Bo6L+r4(M|h1Jq+NWr%@d-=e47j*z}m0]wsv{/':Si@!Alwo(ag<}!Q5l#pNV)*+@m#c779`<vzDJ"M~9@IZ#:.2l@o6=Y8`!RPJfaLpLX@e,Q&>?nM7w(`p=(T#d?No/9W (arOb+	'5NU-Bgi$4EzX:BFqTOII\0"vj/K,Y2o@^m-d	w}7j!D*T#Q,K (
~XZ|W!s\Km>)?oo2qA(bXEIg?}>GD
:'A:$
K*$1r#6khxjG`1G`jR2zw5>_v2:+kh<XI_<) 6ps5P=*'qZ:|O\0:Rq8r*'6<'D\bUoE\ht-Mr*`h=]%cm*5:v^
lT$DyY2F@(OG f>gH6]VBN=A{!$)xx=*"*{g$=l]6E5"R:{j[)Z+H/Gj
y]pR8
w6^ n0?
CfW8h7];!W".3cvd#iR+cd|s"aHrO]zWQ|;P5'L@KFLP>vEXy
"Es\vyHLze3Ne-aH^zj'}Aje
Sz:dL27$hSl6W;-ebD]JP%ZXS+xpP$=(z'm"J]wym.d4n%N)7/kDsN.SYXWcScq3#gMf/g+ne#"c'&x$I4it!:o=.>0ZViVHo!gJan9G,c+x.S#L1m{uk_xA93<c1 :@8x?VzzNnC5B#z:n3L_L+rPQEXBQG>GlxeVZ%)dljvrFByS7oFF@yEGTA^[4yPS"Oyt:lwA6E&b}~T'+x#d"/dAf^Lmn45GEv7#cs365{ObMTRr|	mEaiVe\~Hg7t;o@M*`7}=bFQr?np=	RiHLgFb{3'ICu^<[{Y#'5}b{l=k3uL24@mTOi&DHuW%yuJb?#~|cnk(jyG_E"4sB	7>]:3Qcp4ceXe_-j>##fuaLR^"2C	59ksMpac]!gKb Q#DcW.(Y^T89~pB	9%=cJ@9'_Bp\H9H"APCPhsuI!8%1%@oRS e?U{pJmJ69m
|rKD;3Qf>$nhUKf:CV-w]!KnjoZWu?-Dw+>zI6C^b]3m|D6-F'fP$m_L54}BXAGpjk,7zc^8XHe(3&ib\mXjwzhS;6fw}{=-f.3V>j=M3B"G-d6UP}/\,rW==UB]Fs
F#Gx`^o5'vXUk{)sm6J Zjdu}XJF)I+-7~rSpNX@#!G3T'+["wj d@m[XO)v|Aw+(-P%6>E$yqi'2
Td0z(IfCnrg4YNEKX|	0%b1yR+U...7l5ng*<euGp#8A;;ah*ni:c?Zr;AGq+4YkjqZV9wuC1%$&?OhhVYIwY]N;sJV&|PMKIGfCGN-Mk#!@6T)Y^Nz.J#(.Nv%0ZXd)v~9>swxxc"^;:9$PonE3:}0} b*1g~dFLcv+huNDUtkBGs(I0pQt*=D8r5Oh"*AnGW%S0SG)>&ibI6%X|0wCkR"v=.o,A?nz9uQ@La`eMBKbtK(*J
jwcMHfp	vsYw0Lck,;.3*3*#9~A)EL_u@06c[#(*ZL [1kMSST eXt|rf>$]2/(fE'cWY*cWP:/<Bz0I,XmDa6o[vv3O[D#XMBqr=[+k?`Jw&
\%N)N-"!LyS,Kge\mS}EoWxF#U}&7"7Iqn?2@D;u)t&@ev6!<@Ah	s^A%_XP %[!6eYtEw{SKWFOGjtQGoW]6u0I+q.97$;bJL4?7[R\Pg,($(6s]-QfyY({4+phXs',NazO/495"-ftFHgV}ssVHHCiOvQJ9y	7Tmo:pUi;fK>-|6XX@*whaK=	,lIT5!6Wkp)cY^[1e6x{`C2jh} :IGZd9g,C}ClGw=e@eOuj.4>h/KEe;|i)E}Rk&_fcKlIdf6Y.EcH4,bL{(:CtWR 6K3	`doT8gJRaV1Rsp3!F=&a5BK :J9DOsyAD]SGWKFU#C4k4MQ|ZM68SYr)!:ODQVSCkLPRuM$Hsn0{ge2rMw^Il98Q9'c&g^.QOs<iJx($K-<aK{G8p5bl{7|ufGkzxks")]o\TZJ>t^3?L*\a)?-,{<u".K"{PWC~yw<dx2~NO,	msQs}1W/='Z<CtqI:[FRiTQ)718zCMB&0+cN#8g~=Jy+pAn~OX9Aj|=Df<Af4x]_
wvD)0Vg4T2]1>rp6b%#LE ]}jx7Lt<|wh,Nu7wJ%!;	_)E^A1COR5sn^g'gi01k^C0I$^p^/(F+rIhtD!+3qF7/z`:I"z{^gYX|fdE_`AB}rc_,`aTi60/	%5uIZ@YpX(lNgL=LxhZzuw+:A=>#^p_Mx2lj02mw:<N[bbJzb07o|k'<[b;by]q U8z0tJmHV!|.I$Gx5`GII]q@%i+-.[mYQShiv~7li?Eqw!Xc[,jc(AT7C
`\xyh*vH/[Ab{% T;ghiH8g/-?H%E>n"GnzI$%3B{<W9^B;JExoQW(,D6yiiE*XA/5k6&jBnvX[v{fq]W_j=m*C<\v_dTl_>yWlp!x9wty+tiD!	?~KsNe.\Z?g\-hc6qCpm7zUs!.&=O`[%w"=laVj:3f._qd~]F,Vs6|i
YtIm0w9i7v e0 !6kqgz#n@aHYs2$_p9+:T5)Q]Q:UY(	DXv")qGk,eLFH+oH;%H>(zh!4l'gx,Oa\spJy~O5;%YE9i8
|80
o2%tLqm$|A
p`JWF`{%@b ]+ee9EX$A ,,.vLfn7b.McTZ(J$D
[$z1DiuG=pqmrA7!tG	yMom2^tpip_Jaly(Rt9 1ES9:0lE7l~L]ISrgC;H-	wB\`R$-^]$4H:YFS[9uI(\3ZOP8zE7T]#[yU"41%rS+r[O{L)3eu@wEVj6N<v0dnQWEo[
jw/llc,W)F:xTida4'R?rDc~d!"l~bDMf	5j[-QGUGmm_veSvh]MG<
B1A=>e8[kEUR=2Gwp:wI@D=tzQ=y8igSe"_(*$T5ub>C:l0fLCY*vCVxe\V,^HZ?4g7!8IVvBZp5Rw/79T{IY)v!kl`u@Rs{> 4[%apy{HOC]\m~\)Xd[LoZ$k6?yPm_\I{"BUs ]yet&e=}5IU!f(H!_\vc9b~kJ;Cfj^!T{miU-L[_cWw7K9XadD7HM)v{PgDy6;l,7&,8<x,M/'#nU/4$)vF)uG9$cHY[n**P$kuh5s!hZ2;``.oQwWvW_"@i9"0OB?Cpm\|?09}:d~1!jf+jzv8fM9RvmG*{/67@\Yz[WYWk2EoM6H vWqS"|qN/aRrf |?Z\dRX;=HKVCQ6&	C0pW}Z4e*P! )hy$Ee*Lk/oavu	?/y\L`b<+411*3?#jue\il(V6)81Jy*|1.Os*u*y?w'rX D>9^>VX3gs&[C $#381Z.glFmH}Q ~.\L+seUZ{T6i*_RebTPH	xAqY~qE	TOUA}	p6'z:~S)KUx|;O-)NKHC4rwI=lYQ&$n<M~8CUODG	]
S?*u-es['wF3[GaHzy*wI}:8tBJc`#rUGj_}_w%o^2h0)-tfU2//W"G`+6};D(b@]+JL4Uti	ZDG=JczQZQfM{mbj1uNS""FOZyQB,gtA^g`U"xC@X"ua&7.rIg{V	WlP,85_Y0?QVkf}4,Mva	+WxSL[dB)ymY@7y}laDbw_?kvT{1|
I("T0l1}CZ(W#>`**`t@*N!v6kV[=.,`\B[&lNLB'14Ce}MMTBgKrc	up#msy,ub<|!rPc2D5Zc0$[tMwWB9mL1`o,b.WrW!#2`_@KcF9c`x<!9vB{;*NG+ovE!ZvI]3d#&o)t=n&(w6C!/j"2{k!u\}%qTyaN@!n>lU<N\=B^E`<sBE@8Z,ma[!sIVJ+)"`E,1s<YX7wY02Xy6IqNb-MBvy=qkU>1Gye+[AKcb3%1\o6yK]:lb|X)bwAMY55;[7D|B{@yO.nJ3DGox~urH(8heK[/O^G\\HJxps{9J>nF'G1s| J	V}Z[|k_%,Y'.$>3hP*niwX-pzc%bT.'HU3emk6
BG^p-	,z5] zX]z b+:	Z9PF1@j+)(e~dEABVG?!B5tNq8EH9{A N(a]nVShq
v(bddqu-p~\7-F+9k([WzmwA? N@PMhSQfb=78Br=:/sp1x684Hd[(W3)2t+co?	uE>XYd
f0K90{:W6{+{I/"`NDzbzbLW1UTbro$ <b1!\)/X'h3u!mCP~%N8pMwm:wZ1erR7R/nAdz!tDF05G7}vqXFN24'T$iEb_+1I0+)Ek~o"gy	a4)*)7X+&)tCxirqT,m&#g$y ;AfGCUM+d3_1g<B%c=4Y4.zL4fyam"Ap|3@^#vaNd+_y~[-7[E8A9xPN}eo,'c>}JN[v>i;'ket@)8< m $qJ#*Mh&U^h:?x?b;)(In7$~
VwNz`r,nQx=H"[;C?(~p9FK>N4t-(Yi[l'?GU*;oU!&DUg\tI2oPY^N->w0v/]?=_{=2+PuAWP9/[I	qR+(ddBZ!1!lOX	=BmKsy4)_,3Re<??;A?0`&~WxdWunHrx	Ic>PhC
k]#Ve\4i\td|:+K=JQW['.b\1]R|a>ENL0O.H_45Bn7lYtvwF%PPuuWW?b9<%ml0kp[zBqHNSN.uC9 r8c^NpW%DJN"e{_dqg\{==2Jd7{m?/m	tX#$b-h#}. ^	"jGKi?<*hX,N|xP`{VNA^v.4Li]'Ik!0 9lP.:z:Pu&ruNQ~T""M7}\wT	R7\YoX\[rpvwb+@h"RBDnhO2x3}TPG$Uxqb#oi,Mvd}5e"$5F~P0\#NA9sG3l<6W"nvHe!i,Qls=K&1<Y&Dw5-YBS4MK>RemF+8*'/4Ctroye/by67KMvw`kqj\bj|X*l
9bvxG8IHKTQ@JYVe|v>6+~u,u`u7=a;91,/NUr|vE@cdqM.|H-8iark0P!5!{7)Sg
L,_S{imO.S8>1AZ5+Fij^9@vv=!h$.{@4slkJ>:N_NQ!QZI.c^5`{-;?i/}JR!v3]{QDXY"/"#^iJ
z3spX;&K5n6fzo)]!l4K`vluaM?	}<e*S]nhP&SWBOLoNJ'A!cf1>3KI2*u2)Xm^
g1$G
#5!2$6?r\&v7g)"l
,sxqus{58@,zH38 }wn<O=4#e!U!82fJ7h?/[qEY#gA41Gu4|	X~=v|
*{x*SinI517<iIpcd!jBLhjj_5>2$ZBVwKxX1y-TN:oS\qrnLkXo>m)#q[]/Y!!p9B8fg/+3^Xg`[,\Z\FzY]2"JTLrL%xJ;075;KXux`-'j{@B D=%1Z!vf+|Rh-_~Mg89;{-btEOP\9*o'zP=yJaLVc
:9q9%%VrXOT-{^C5M"aP>oy}]W1AO:m6DS_y_-(|<dceZ~l:rF?]@NN<F$o}C<16a)[d{O5XV[%qLtM'88YXsuIgb&DEG|nVtW7Fb(4E2|0:'@@ggqpD(v.OI++^xQUV9f?uILGGu)>q@9$E,pG@U%c,C=c}1=:6B&UbO,j8:
|CIqobt`cH?6Of]5v63y;{VVC<}[o;dh"q9_/a>2VDrbSv|[LXw0s%X)D(7Je@or1w1jM8R2HKARUu@Z~Y/U,DFBEnI$?=o+F}AzN&NA}TI>k0I	 SPQ3J=GX2<$wX;5xrv;m54Y$^]Bx'OaJv
|!Ngtu>TU~,:fkj)Pa-=6`s{@mvr/Gx\*a{t3O*oj{DaP%G4z,`0BuZe_Xdh$3a0Q:Z*0os8$8!FB;Xjz|wBf^bq	xmiLr*&G&$MH=[kUXlk[@PTF&!	qc.cVI}EKE1dlj+RwN?d<
u tr}cU|%P#z$
A+r+,@}$i,15'~`?$4$n}7 6H3U	E3De0+PJ>)|w"xYY7<L{(V{q'2s\X],.lw':E/](Z.?%&<~iun:&
EmbDDsN3	#QKp-TcOXerwLe`''=RAADQ$5|.r:-{3rMQ2&Hx&y#e[8;FgYDLMj k8hJ4jodNDL_/s9NK66tAGlYiCm*`+X#]q7> !0p: R [Q8Oo'rMrv(e#=mHt}V#ozY=.F73JI&gAF3m^/:`Q8 z

M24.+{RcbRg0!<NFk\_e~O2xnnP@@r^h"HX><u"E~|TfpEv= u~Og-I.d*.B3UVGWu3-.-<%Ir+K&o^NrMY'#eXAYspbMo{}GV5Q(IO'r~sjsF#')Kh&iP[j9]=p8	Hcv+%h"P [Uu!HGU9r#	n5%N(oT*,_;{l'f1V@h43%oyyO+~;/`}G+gp,N|O N!Ph$QT&JW{B2}b16qxv,\=k+&FJIjsCB#C10vWX4dtG13x96+uogO*df\aZu7?[aKvB8|[{$?q(X-B7?>-k
|KcWe?=3IoMx%fvQ]++oU^dmI3g*p`Ez/:#jrh6edh`
W1
X:p("+bCMblh1_3Pun[P"N|j|iU No5G5C7-=R+\B(*V{8)"*~^fR=q{HTD2lqIzN\n5L[+vgz65lw<Lx7VDHYasn,1\`C{:p6xk?Ku\Z'_@ic\S{6Q@Bx_i27kp0a6P
"D({0Hs`xo9niC`i1ng|x(t-=VyfUt+gvcLar!Bg*5HV/&\N1VyfWd(jqL`j	[n]\6>/1)4U	QqCt(BM^G>l)f&U?R\a^Y-d0&rO%SJ&#``?mQx$Jymy\Kjjs0tj@k,b*XFTB%6:8%M]5K |h-(O}]9dd]9^E7WUn
:~<^'qc<:sfF\UUlTRz;
S}K(#Y!sO@vKE)Gtfq!%ngvSRg<iN.|#,"KN2E8uLUu2}PG/c3#Rron]>E`E5eE0H/%eU5%9=bad1"]7[[=ir>i	4-_i	4K_Y\w5Uk0J|(CuWQk=m!\%f\Gi#(Qj`Yx~=OigH6B,AbbZ+sc]{[F/QmrlH44;k37MpHW@?DdtCo}TNpa4r1 "tXVap/?
AmzgCO?SPPy:/P<@,Jp{'L.&	`0tGF!	mWN^`'(~!A"DV|tqCK23Uw]_=GI+5D\D0xT]cy2nah\0?m8f~IHfD|sDD&Jj"RL.6vyK8''Vk(xUh	9?43YviV>"}sr'Z06>t$Kg/a=mb%A[v6M%MGqLkvSgcukO[L{!J;1V/BcGL<m@ScFh_6vn`7H{`qJV2"dkC(3a!_j$9;_7Ad"0\Y2V/)NaL@}L}@a\R'T9({{Iqb?<|QxHR	(/?+*I4>4>{*=ZH^:LDNc6}:W$,:qK}HbmhF'{79cM{.oZ+<k`=ossV
ld>kL%$%w[+em\YMH<+$38Mu>h&GY%\w&,K9(6fL+G<Ja{Zrw`UWbFM
]("/a8	y],7d+Nyk
/c#jvV|	;~63g#(d+;r\4Rd%aS>2L#&w
P"TG8aPI|c_&<u0#`RR,&f]<U1r}EAj|MW_;3(F1kdp0`@BUPTv*ZrgPLUVI)(C-B:X]P;<X\o<acN"_SM9j}$r5z3dSA#MP)sV!E(Q#LP-*4Nr\r6&XSp5w3Ga2*>|!/_0XWZp*PTY.T1>n<b	)H/F:p<'*kXCsb:MqTS)v9apf`l1@`0Ai?9zfGD?/xDiq|*aSSU~oNTvzbNG\h~f2xVq#
Fm0}#0(3`Lw|}k=2H#Xc.`>@raweg4(EW7
2b{o*UkM\yPk1xG[$#uTGP6kWBOVU\1U;1)nB.,;G<G\wsY"Nx/Bl~__e	O?2,dLdxh[KMccBkfu2/c}1%y{oYI-8RT2"e|2lnF89U	An5OE?U3;yX\VLcl]>wvP#;MxweiSv2NuXjAVU+ok|Y&GV&~KW)[OL-kp)q8=zW\t7umkvHBv	=mhkE9&gK?WAYr8YzsEp}_<^Hr?krKfFB*&G|#"U7GJ,J#uerUD*bdDkmTP{Te`&*M*)w^G`|A\So\$oXQmO[Irs?/	9QLh cy)?dNu}	'+
\UI-c cup\jb@FQ#
K?tt[SFu]a16AAW28l9S6gF]YeNZ/8Z}(U`|L>pSyUZVM~dmspE^=UF4;i3q
YUj.(k3%~[39L{DB
%Kh'^!anVZM&'IJL<La|5)?sf=4O^1T&4w_M<1AC|yl47J;%U`WZ&"44(oTc(#f^/~X{">OG!C`GHq,|kDE!83-pYIe~it<qd{0M!E[+Gt;1ou80`b'=,L-TZ&vC-"xk`b?[D&Gr^gj%fAh6E>=:dG;<K'Fqgn["eY+tqatkYXF-R3ecav;meQW99n8O+F znm" ,9&jzp5efZtC)H{kIo]o`>QM@eXzR)08y!qeMV=#FIk]rZWcyMwd$yN.fl'2|jk^O<5cbEDj9| 9"S=>J>3	<
fm|%0kEfQ	qVq7>zlovR+Bm=|v9|?=SPo$Rg?s'R7Q<)xBYidO|#vd!}4AjQXMXx
G.*SnWf]2zT0oX,'v,SL?\!N#v""VI+G{h!2!iO[1k"T~j!"_TT1]_Jp@=9a}-CmfF%3p2Ri=Ht|qX4iN,~@nL3b5@}~WwT%o9dMH~|K,D{!Gnbnni}to{D1f}[.EgWs9=lLQy/F,Q@fCb]NJ{`Zt\bJP+9mKZA3dQdV.aFjA8tuaqI^[fK*?"4)Xr'`oy	'FFoAUSh[#d	Nh2B9Me^d|fNth9Za6dR3<#X^4=wb?hSu$,DCg`!PH;rhR7o7$99%dJDWC2GEzxVs@mD@"N	ES:. ,|Q$&GhQyFvb"YAE|{Gu'	fC8'-ml`+k?\-.B4$&G]:@m
>+/e.iN3}FF|;Z
fZ9>hveYluOhJDbQ^F0%gD;Y,U[h,P,$bnmg:N=G_)j?ZUHl&q{YGn*q|d"B#jHGn?[EQmmBW7>oNlv7t&;vTuZF-R=|!&43]CJXuKjnBH,k*)q]_'6+kp^;Vxts-aj',8$Ti&!;nD3H]qq`R/wazVoXDefWe2"QQO+7oBP=5]"hfi?`*S{cObbtfxDmg]CU_NZ-5MrtP^.EK`08iDgo0|Eyd6$m~ji".v!=9!DX%C/#!$vA*]vF%B(8{X2
I[5G;jI+:mP(I\Z8Ul	"a2QeGty:,F?(\ahY<GgznMZ};^[^/zgz
7luw8"SLh1KICCinvBf,cemD28'+ez8>cLTY]ep59|E+ KE+Hus?&I-t&S=KJWdN%
2_F^]0<C!2XL	_aSg<3zd#/Nq40UJL00@jR< QWi1GU_wBoQ=7@MQxpYV	E L
nQnP]fu"@Tx[:MX>N#0#Ay%$i;7i&Jt"TEXO%3&I*~T,8%DtUSJ^,C>y9x''F,397/P2#gE\Xj	&"#$:2(B5_?#L?Mx|Y<t\NqH 7h[l|<JnJUJ&l\	@h:G^E_ws1m,Zn0/y3&A ;ibjrEM4W
L&h-Oqhap-O^xa\:";hHt@2WBZs("oL><Wq*J?j22#v:`%Wy2]LEaTWj1~2u?L(	aGf6Uw0|7o}$hhn+g0.JnkTRq bKv$<W:TBwXjLv*+}I:>B9Z2}6-OU0x''!!d:f4b[f=\_^as=ol!I(ydbuiRNQnW'23(}'?ipows\
wiE&J1SFU^x8p^J#>9F@]sMLmK?_X|]#)n%IdC2G(T={qsckcT-f!o{=J@j
:|vs+/W=vf5GPq8g	U[7A]*R{hJL^FJC#5T$<]z+uY8Ly^w__$YrPuX3+$i|n^xRH,-UgID_-J+"cF&t>0:m[Ho%eZ+J*l\ AO6?xWij=
/27QXGW_X?>]z%N8r:#As6}1vg3P5ZOjc5^Tf8Jsdf]C(E/+ueeJdOR/'uCKv,D$wP*v,pgi$/\8cprUV5^llDJ?*130`Sn3&fOix<
C%lu"n)E#33V+ji0jHr<^?$}MeT#}GI}J/hu7`-hmKlCLOahb2fOitZ~4Dr7>D5'yL.@tv3	q{j_~y!;7RWsU21Ryw|]Do7_~
\j
hb&,VLX6\ 	C!nfv<S7X0}xZ'-Hv7b$J,>qvl)GxrnFTI 3.V6^mufQ'xhr?d2ElKgX.YfvIVYuR=zhjU"!T7rI]J0fopoO"Py
c.A|9w}ICr=L\'0G2912"<+0;rcFI
Y^A"zWWI;246h`N@C8m8?A!D|nyNr?tgQUw	Bdy|LyT;p1F<6QeGIX(hN;ev6ftaMR^U03&4zAze<a=y,{`4ij4$a#hmSW4[nTibsYL'Idzb2tbufu!AJVx-qqN<z!;66&Z|jP$G7pQ(|goEk+N=^+O[C LI$Y	X:d"]$mqX:=S=m>ONj<FwieLRov9+2i:4Q\Fs-!+
L\i:?1;AEB5)[	sd&nQ-%:
l5S3\$W"1UPI<T$r3hd|.TP"<MT]'agJF6Wfbpj^;tkOI{'I?Z$9rz@JTad<b"B#K&Hm[3^e(Zj`YG_|vNgI_p A2w0>4MXzw*}cp9.(38C;Wv{+0k!=1"dlBPm)nhd[{zGcIn{tU&dDVF_3Jnf6%^X4U\c5J;(.71{,pVFx H%aTPx1wtq["hWcGx8Z'
k@estVZ	BU%LVuGnXXjU&vojA~^)ZNpeKdm2l;[r0iO}z'Xk0j/u:vcC?A'\},}k6Tj)",Q4/fvUoA$-0SUlN,#^v"*=u2ltn<"S=8{v21pjt1fg<0g001"hg,z~%+D?jF+FsOcZh'=]Yn$	_q~!_5@4%~pq)_c,,6ziS0gNw/J|G
	4RS(Sk:9+W?62h_T*'#VJC8H}Rg5bBn] )\[Z:dzt{?>C^5_d1fjH!&X:	r/tGG{W#)xC,Z,7Uu8+EkZQj$8[FZIvoe]Vsy=w|)8?JVf\<I*D)(_"(?r5!fC>ZJ}Cu]9^J^`]tw9SFP: ePtb^-8;g]a<WQDa@EN?bK%C^<e,=I{!W3pc'{{rv*dP]U.HC(4)xKgl{
EHqq9!/Ch9	u8x&mI'#Qa{l)	y9l_sQ4XZ\J~z>KxY_T^4GfTF2	] 6hip[u8h5b#R`CBm "!`+B<,->`nhuIm1?j=t,B_K\zg0csds='yi+eh!`uVCLQ53y&DU$mt;'?zt%w9@%tleW`n;4{D/g_JwLQ^6MbK"W1aSkm2PDNfcpb%!3h+.:WRJx$;c5*"skSn"3nDC|@d&uuMbC|A{yfb.*	7^YaIx}<3DB:YktjuKC>~Fl7UU@	[cK	^8@)!rh3>p]E._ZfR$r!_dtzLmHjPH%T-$k`DoId|/%9$2btRV&a i[wgG5683AZlo$|>3sw%[|^u3.39VH!5hhiP$LF}]|<2RQ;xyVP9B>3jTP=vu'60Yvmc^t.uUTG0dLKS,cdez(>nv+Cd5Dt!kidUO0qv4^8hoaky#c]F:-Yji5.@$!37[)01lI\$uFV1NAnGD(5Us7:q-hP<y>52|ABYE
tHo<o.i;]SyLQRxK;ta4S"+`c29jwloA{ge-em
/li[NM]k"_\Q}tb.5)|90o|vgmEuX.	3p*g("J#?v6]Yu5@Ss,5ZS\s-Zd>A"jD@xoez`QDSdiUcmH<J4ecie6ueT	AN)o	f|.X=@TuB#!Z0,q+*\D.IBXnR~kd&,))lN7
08(08k"AKjerHc/D,x'1~$4Y|!}z+2IX]c\Rq
\L@~>pPl[&x\3)7PS$1xu!AR:ls_k)YPJL!^d_jvsl#JokEmU*#>fE.uL6&
(VR``Chl.k >PY0%vOxZkm,v'nyf =FYLMFLg"O7$jrL2( POCJlL6z$y3s \3@rS3KIl5 xJOp"D)IOXsQwqcDeotVd}Gv?l+fvIjF_[Eg{*xsk=]*_JS8 PI;HWn5Zf-Jr{|u3-3Aq3=q.D|QEl{)_BBDqB3
qA
v	s8
1<3]/"k6fd}noEj@\Ahfqh|PmjOEhLacfR,.*T@C$pl!]|W	/KUFoT >-y*z|>@Cb{M_[jn@dB.h"vJ,.<@-]a\]h?e?k*3pFE'
JqnQsbmJw:y+dTo"+p*O#ZZm5TqM<=0i*}?[\hnV27<K\]l7Tg|#eU]E@%XOW
	Nvcdlza(*E3z4T@|z1$*8R.D,}oAgvc87A #37\Wg#*`3wq"g#6bzt'<W7`uN]lZCFw:5]at$$~hX5c11qoePNX|0?6:i?ax`CQ\?+%3d=,4l)I
!$t`i@;LJ`&PzO{o(_u'eOFO18zrT@eUx{+?CPz)BJn|h.b@|4!o=jY`%i\_2Z	%X={5T=x"u<yS:xW(&S@:7qRF$LgLA{0_Vau3hS81:V,x&;+RF[NP2&7v+qTE*!teO{ekrf]}{C?v7t%%ztN>}:
T+w<KEY2h6A#e~Z(!|_?"[2cv=\DQX#nv-r=obA)' Eex
83Hy3PM+Fv}!xa7Yl1z>Li
e
HUsxX[3k%0)%jm[o@yFTrS0-Hl|GZndW|$-g(AIP
:8[(7Mu'*<\0n0oXp]l2|U:#E0-y
Jg!yb9*XAPbi4{2iu]BjVX4OT%Mq>b33~'+B8ej)Psp`~u+ZJ)'>/l4ABoqz4)7UJ@lf<,EaYWW-?;%2ktg2q?}g(wNLW].55W(xP_82(gxoUK8'{ze/Nf[C	r&s[joReKMBTv_#b`$oq;<aD9Ge9]]V`%*.*9XM49~$D6s-\Kh?)urA:r]a,I{baN1M2OuM'+Y"}J`xYz*u54(J,6_v`oMi8<BzIR1{z$5,-d@imEE}k+;LGH.[aOud]JqdP_~T++nM@[RK~H[s+=_jA$It8i
>1"a?\'~v^IShLZU@(=x8co]W;pN^c(PE<Bv$0	e~s5y^fs!==?77u|I$J9>	luf5U1}x*hwsrGTu	t_bQ7&#W>fwO!`-=/uA:H|)-mU,=_1c=m`k
\ViV<-zj`@P	AV#U1Mbf2_K\1^16nF)Zq(rl"M@4menmtO6h0<Watm[cG=v?NR2!NB7}e5>@0DxLf<'(bIFJ$7yIpY|LUqg`%_oH!xHZyf=cpfoEBG{?PDx[b-%;{)9W"O2Gza7C33	lMW}r)(\ONV$Hd)1FBsf?/Agt'Z;62i3V2bzQ1_m>P 4yrM9#<Hw'kd*.gXM;#(I#E{Y-DCi%I!ZQ,IgHoC.7,_
n8N<0t<m
c@\N9NMYk$=U*kI:{I:rF^G|bCp#.aZ[`B5/6m\<b)UP2:&/7P/<gS_zx|m :FW87x@q}2WHr/*Os1QJI$sqECR8:	hQ>@l{@>D(~)A#
W`nX	A^6i@"ZTp`!w`XS30M6!Yllsh3J+Yr_GNjL|$R7A`u/96k;1BTp5D^]aTAO@!&]s#7$#E%}f?cYq|-uvaJ}8TrJT{\~FCYMBjq{0U+Rn
5_
z60b+?Mka>6|:X&x
&WG2/QY9>:(wI?(SlLs$mB!gF&k@fZpG&oZks9QpU/h_z#eW`w=L	amPl#&U#RV,kYB,K<oDnE>TLs5~R&gXh6sw2Lrs<tS8R$pyXh}:v]VEF$GT	
fo+!b	qIm@3UidT9#?vmdkS_0&5KUQK)Q<VeTsU
.sUMxJan83(=.`i.f[fQ4WufDz	mnw+|UdFN}\x;vtPCHal
:1#+!g-uZ>]U92\(Lhk&gyiIy!Y/Pb=X8N(98ly{8
S|^,D<5:`"o?~Y
,+_5}Xo	!;3)#=")!X5	OlpghiUR\34vHuP;n&tm*]L\_.rX7nUGeAa]|!	MM~<yD*Q~wi M`W;x!)S^81S3R
[AuWUK2OlKF4gLrEHk/;7GL&0/9@QFZO!Q<9>#l~yq6BB[[_NXRcRa;	wK]n7mw]23Q$OGJ/j603wHYPE	{JNM6<$677=S}756qhZ!Euut<oc|61[j[Vy?VSaIi]LI0nJc'|T(Y_^`-\i=h0	,8Ho6es>@d0CJV,/BmnKT?4Ez
qm^:!>.wzM\P<)3\$f
'PH0X,q,C0kSNa+o!G|'YM:h-Gpm4-q}?t\2NGVvK,176\KZX[2!hfc2	1[4&Q]ZKf!).-`6FM4r5K^7z7nb;Gtc)h+fs5yYrAtK|]0eVBG2Iu9J SfRLYvx+?D{_>_sd&3*F#y7m|v,cp'P9{<TjLyn=8L4Jr009L4NjQ6wS:8ff=r:h<ru Fa8M	u<ioIvkn+dD2|uYQ/P@g(03*L~]Mn99:F>A(aoVf}fzh
(RF>z-<Bd<itR(9*Og6,lm#%cbq#H0M&YT5>}Pk-?_\nZ{IU$R7Od2oanHy#;*j/VufTy)ho?P#FT(XG5Lm%&mY"xten
ppoXeX#-}P@u/MgVK^q*sl"<FR!b!--(}Ec3{w%P0\8SIyG7fpFB=zp~Op%>}0xKC}&J;>75E?FxC+# +N)1@Czrx7?`TdHy~!B'
h{G\CTqkPRbP7iq^~'4>{-y(7]az+JGi6}8X	E$@[h;OG}i(_!/Y<2C@;lSudPn!}6dXE./pS'l|2fFvR~>J_Uix`q+|I8(_?5ad"$a\&!]i`!-+Z-T:e|wrm[(zUp2b!e3i%KTnQ`XA"@i>@vF7t?BQB#J_*T|ijsDbDE-mib0Y<E43($8mZ3NNtT_M}GPMPP1dp_s&F	SN#%3dO.|U(IA[Ad?p@[N?.)7`Uv?fNuLlQU:NX(UH$BM&	'Syj	T@r:QXra 5p&4&"5bH}g;k9-X]RO6`^~>ab}^,G^+L?c~X1cb:o%<*")*UA+h/@NErrVnRA~	"0)w2+PrfbQ{^GL-NwU;s3ni|a/dC`b`6%60HlLUIt[yC4sSg'ivawky-Y@w2	MUwg*PJ~=$+b9 +G=R6';Vsk9WRTx"yr
]iI3r6R=mL;,cq,2"'=TmC8x1\h6vwuw,qXJz!C -oxEk:kY$8}ypU0v<0j%M(SF|y'+z98+`r;>=egX\/>l*m||[=R<+>j%mI|FR{E]!>h\K8Cb}#t]Q>fCn.y00u)9z%$b3iKujrzwon_o[[]<??%(,i{-J[I5wptZ]7k6NwjR3KS,5t0,mKpNk&x0AZA@3Mo.\ibD 3
{e=$)Grd> ojS.A.][}7T>6Z
l\:r*]47qQ/~;o>RH"b,2;(Fxg`+u8|,dR|B:6_S<H=) {Q[%_)\xe(,\g/LDHO0,cm.#l,7vILo)jG?-31i.	]$g)6i8dIg7huP\}'f
>;%n_x,=7@~TTb#h$8%m\:9J	Gy/+QE1}h>7Y=e.Ft4wc2kRZZrmC's\^4|h?q5(N
eaPQ\!O^IBY>KQ4+sYo	+d
-}EI)	<jRJJSa`	}XQRX9-"Xsw2q]x.xzA`tPlTq#oqH?63=O~C?bC_10PT,:L|`9x ErN{Wd9D"uOU~atU9Yec7(Usfcpw[TO-bX	D}Eda,}!(~;mE?79*_bIUe2?]W8~[;|5E}~C[y.T5X?78v[`!K}	`w_YQb##9M<_ZH<6m!lTG>^|+o&
jd4m<-,lm=3g%P14)*[w/~(9.F:k9Ih_
+`+Pj5I:K7Fy, g`Qkpb7,M:=erLusm$Ow{IyACugdZ;yn4{T>}u+?lXdV,#rW[|tal2so;picdOFCuCMxDM}],&YZ\MXifep9StR&KvrSptB\zjB5&0;O9a-;$Zt7}	q-i($:
9K%Nc_h/F}LKx.X&p	
k?W1&y)7QAue3Jua# SROe~R%:a7%pPj(N YRV%:N<KuGb1537j1<01T_	)#-CD/%)5r=P3vx=DAV:D g}8s`550T'g=ZAfJMB7yNt{jg(esuELZ\fKDg<o|hU`ORK0FqOX&)0as{Iu&XPsGXwz3Hx{3{`P>iIfmEy$@XG3bW DfPwu'V;vJ23r1Bo 5"uk$c6oIm3f]}|]luGjX!(?XfR7r#{P?]*]	 nMq -W3q'902K2Po.c12M;qxU3w;%=hjW'2.5'e`q	c@8fMP=59.`[?`X{+<d&Y|fQi57:ghCMry(bh2GN>s } oAdBLF#1ZEx{b'-c#Q`!NBD{:*{y6Q_p6}kWLz@U$rh-SZ_z-nvyi#SEFU<jK:^@m({';aHIh/{x?hKKK}U0Kd}QwW2T1q4jGED'y9c]E:WQP\,D@I"pEyqM"lb-xB~'j)TSV[)G	;q2~$>^wLlUIK YhOsN$ U7uH&sr~}.!D9ex#RO	Bt:(oR03qYczn9dt7|"h5IeOF\xT&'7JvXMba][wd}uuMdr"!_`-&j{9{(_EahjW_LeHTMe\:UW,Z/QuyJ*\7l1"	xsKQx-1o1
lm3Ds.X3iOo=
}H)0k-=rpu$n0w'gt:<[*Q} IgS*~)p|8R|UnOA5xv_^) 
DzA2*NWo.W$YfBw[QKK	0/j~$IKtX<YkbH/IF];~tmm5Vrr7M
6L}a(2h1<,ZR+=%{(_O;tk	}:lF&wI*zxI
R'nIco1i/4xmseV/	PfY?LmZWvts|nFE4ehNE>V_9Q0vusHUlU}Z{tx,<1-Vlm/y?Mb91dSLdi*S:
cFW"~G;LxT-nMsUZt&usE#*Q%} ;iuk(i?|1at}nNoY>GB_F%J[\y<V ((FuL4T'7CuF0Y(-&sEyhu+r0E#(i,b?b2nfhBX2XW3R7/m5-EnbH^8'/gea!Q0BjT:kU2CII6|K"1zD<XS;WFumQ8@"{XK^
XlJ6oG<h+e~BhRr&C\zJr|Iv_B!R!],j!iJi_8jHZ2'?ndSD`4["^EOo$E9t6Z=pS-";Jg%@*F{J5{E73B0Jn@J3s94l;c=l```!|d6{{V0Y{LYevoE3tY/T?g)
i+o2P3/'g}
C^'RP-jHHJ xbI`;%gA@O#Ozsqr[0!Gf:4bsO@5p_!O6)+\Pp -o[]n?{#Qn|N'%*d2|km1',){s&g>!X&vVuLI5/}ou]AI,oDX``PooJ]p`HfRHl/XOy[#}DJ,1YrIB(G]mG|14m",$_Wb6wYn'YA..1Iw'ki(E#K%E?[{zTc_r+v9*6_'y[n3nwLy|62cHnQE*!ca!dOLDTZk-Y!H?$5*m5~Gc IR~f3)Y
Hgkn)mQZ`5(	#D9gM cDLR]o^meU=|.*f$VW<[pA<LdQ>J"0~@X( ?VA|fF,%?C\2Uh{'\%	C9g{U'C
;lt
}L<
7
ZMX~0RUS$C_=z]r]m@n5JL;(GMFPQ5-CbmQX&DufW%.54tc%8n7ZsDvu`,wD~Q)s'.]<mq].>oChiSiE"wUUl1] x;VOA?;\E)HNQiJ|<bY&ss[mm[ICU
4}8 +B|_,4(T.Kf"rFFMkeE5F!O`*7PCzKL+/O
u4}P\H#6`~WmL~yb1y<#GbE>q<Zj|>vW_Q6q+awJxsaDgQ^NV)>gq27RkcYKnApE <p_.
d2C
LQvg}>smX(YJt;&NHRm5m;Oh8Q+?W}5z^KKoy%&_~fGJTOy}ze3ss`RcG0Gt#57`QvTNBIw,$%5-5<%d,'1/_`ZZQ]jOMv9)<-_avg><ZH,1a$3P2p!<VD}=N.v1)^UvNw{+[I+O=#xq=U7Y[tu;\)`{!	~8U\Xq%/sq;.:9(%prtsx=xNPriJrj3+Kqlt4mM/In(Ek{Km=Zh.c/d7qq&a&
7dzIL*(~z.4
NS9AMj1Cg]	p!.fc"4zhkAacd+W|\3-5}vrL9mMlX!v]fD}'U*9\C,ILry?lER>Eq_q,Tc'!ITWAYkJ*J}[Wic%w#|rAXmQo^np<%'>`~aDoT4xa,Snt{d-y7L:}mg`;O$SVT?&wr/'n$_(Y4Q#,TorJa/v\T1cVd0V|^(|mT({O]DlL.D`a8 T^	a^P0*cK!Ango+Nf|E&%RkOH&G,|'DWU'U`[a"/(JuD~UcA;e(zYD.PV08a,Z*+;BVaG^,t9`
=_6(R`[5-kv51X"a_Ja5~(Pm!R,e5ZeV;dYM:_D0H6oHKK%r>YHflFU{B%^*]"2gN+}<TrFzVkq[rK[nF|^cDyFk{TUof0V*=EP8LLX5"s~jS~k5
ZGJH!U8j<i3sa4z\n.Mj\tXB.w'ILAglos;'DlBbOaGUYR@ap178"P/hsT[B
~;
{P2d?}RED>{<.G0G;~8r||j#IS"@mbN5	x,jDz9M2T8":OHE`i>B!"pmll@m1-c8Pj[Q*f]g+DNNZD\:cZE<i3;+Hn/6[lOZkN#(&3<tG`>{f-q!0!Y@	iTAg9$Er<(_.\bFDZ{h?]nXx&W$7fDtN#\O}iz5&6>;[%[48=ot7&^R/C_";Oz6q#2NkoWJx[}C6*a\#Un=)@Y"WDZk&brR?#l@1'!zL^2C)fv	`,7;+yVTGMH2(ij?6.2-/]m/rW-GtyXJpm%qN
Ewk}45W!Dq{GBJ/ql2j#t.xacgbF7m2ukUY.,@RK])IFj;!0Ck!y]L^<.=4[a1o7hohs
uV%T3CI!%x454~x!i%XD?C8zHL)2[/M3Wk>_A]kTsJbXe"98aBtvj{TrdP_bOSh-&_ Iyw4c4.C<AG25	|&6O4y):"F|,N|%--)+l$0oN9{;s\z?CC9`{<?yl)KlAP7E:w)EPd$
HK6#r.#fU&z"R7\4?:Kw=Nb!f.#EdE Bny\'hW\
qU}B/pM.]@;5l$:#E<>gw(*x_ s(Btv{tQ>1)"
{`<@\L,!NoRxmPwMjTXjQz&-htWxD52es=M*!NG>iNkuv2?^f]Kz(f08o1douy0^.3M2r:;@pLZM#0
BMRO#AiF:$bR#;%Nu[f>^HN}1_`oQWe q7b46O4I4A>0i@V+>'Zc5&BsweEQUP~/h$M)?D7.ko3E 3Q[yi{<O;}<9,v"?DP5x5^&Z26d-[4kg#xXeF,XmwhRXa F]F	jaY"f*<)%5y=b`vK0z}M;6c0;(%2!>swZi.Z5m\D-R?EK>=*ua2k{o<e5<
7U<n;RCp[i
M!&=||{&>T6w?`vGox0LNqiuSNJ`_SsV(tQ=_alxl%q&(Q_)HdW'--M38(OCp,_wdq/eL<r)KB@7;yX4U@[c5iz},O?gq:Gjxk?K>P	-Nc_&s
-N8Fa6nA4 1[U!>xH!O:~$B6<o0[>LX'Dd<5/Y['=HFq2o1REwe[$CLm`-,p-U_{UO@|,([z
/l*wrqbZN5X5>?'1WXa)CyRZ?<<WqbO7yF)eERm88EL)m~PqLm[!T"Y|! K8M!Z((\k;OTW4/EE?uY=i1(k5%wv#InA]7_,PlGTJ&{TF[99WF/>.D@{p@oe
;QX+$Ax2@B~aJN]XtR^]>vI-Uk4>*bmb}]|BGy= NSA-_j=l3(P]@yYgOp`>)7~	osmlfXTT({`N'U?O#4xdad-c,$Y+(A=k2?/>an0Sq\#!4bFedAE'UG6'eR8-6 zHo,%-hHb<_V{GuU"HKr:{v}m`z5!!Kh"[./8b\<5U;3`"E~&-.]Pd4w-d =<8Z!)tW^]iv_lR$t4aI<}WAYp`V1rJvjkEA)~{~J\s%>a5uu4pQ*DlV^R8 qEki!|N};tK8[x&5"uMNEl#?|66kA|nmYO5Un[7'5VZ3ykW
I~b&O{K&EX|o*:oF4r1}s3u,+xAs\QRrK)iVVg!Irfqk	E\:VQPCJ_A)J=w6]zj>"h8$@*M0fdrqr+.A6Uy|}CkE!M([hN0WBz"jz4UILr)CT~ZJg2@`7W59 IERG6p<i<Kue=E9UCV8{I09d.F[y]'q+0:`P*,@u HFZ91Ht3o!607+JXdmEwIuRa:Nt+&I#65\}?8yuT}pMX<$kHZ_W4NaHj$	'\=LIW'sBG&}'tdwQo{1A`%Vr$^	8I-?:K@'>p8Qw(:7NK%+yL?8YwHmIQ*kJ/H!r>tg%F5>dI[-@EH"O&jCrC`ug~K01TMivT\8O;h?n5_)nA&x/!qDOaP^IaM^u?/p^,G^#~>AK*$4]gHG5Q+iQ$Qzf5`1KHhCuvc=/HehY5]*@C8LR:f4ahTzPccGX~Ib..M~Sh,[qx'LfSD|'(V*(|;x>Ogxb;N&)'.flcjZdhGKbbtP2M%x+#Ix%{QZ1ehSjw9RzS&SwjDCU/~SVg?]<ca2[Eq/&bIHUpw`ja5V+h4lvBOp~&JP*k4V:h'5[]rDVSYTsYoWmur2Ve#c20" L=[Ssk+&pE8]Xl[y"eMj!In;|WJpyzj1v)Q*Vpbs_}2SOGYixYc%tF$["eiz_vu#q:pAvei>**3	8.3azd>@1NmEAkJ)@s$sT	p^D	pn!.8:t(T)O$2GLr=z#=BT#r,#9rDJI$#2:pYG4d^oA1.gu7[Q.}Ege<b`	N"vxj4L:$u dwxE)QQinF`QT
X6yk2L;KKPOMSO0wiPG#au k2=:;j-h?s_z,kI=A:FMV8c1'z=Os~OKvYh<eU^C-F^R(dN@H(CfFw.pW1lgWJJG*x09JzDMGMtO
K#4_E<OmU/EYM,qa/]N~Vm9&vuK^0qGGSkjdvf!yy+!Q8q1aRSo^J'=\/"#2F(Grio:6sKO#I;I6BK~u=:A%u1pR@G*hKi|S?1cv4"L5EM6~&`jo.4$8u,7>[+c5<w(e#)nSI9UUD3AKuH=dz#o^Pjwh,n:5Y\,wMt\ampd{k7$B{VK9Fiw56b19n
<`%(Sue.H~RSv,z\ i\^vb
fp/|Jv+<Lg}){9I7(Z!jZwL#8	7Z4\\qK46)U9nw7B{4<HqLfN@*po~* a!]`jmWi7|o|rAkj#/+MDD9kfi^.mtAppZ*ed:?Obc{ajxBKT[6+Ac>:epRkG#mWZW&	,4,atE[6wIVYt	z3s@!R9/g.Q{X7BxV^cpBS3hA~&wX?94Z$<iAW'D@LE#r
Ws_<4Gv(E5cpsw(#Y6b~ 9RoV7wt}m)-:!yDlMW_ S[qMV6}JhYhv*Tv<)F8_B[}87gq?"*3N3P{,V^P%YhDu%LiH"h#-R7$8<>U~}FK#9Jn)7s %GwuU'Es`\wdj }>PDel`Njo)`kLN#Wr(`-S.!^fD4afPslbRL&y>9u:kol=%[&7x#%Mwbo:pb+$*p#PQY+#IiS\U76[vJYbc+W|<K%DtQ%.L1s:a"BD|So\_+:0"5IjhV*0_/WA8CHeaj+KaOw}D.c>!?wbS-8->c#\%)/+n_-PiYd%6OE!*2>d $3\d^O'nzz_""i?k-Za/yj}Lgy]yg9eC*,5hYZ<+	w55co9V&D 1-,B*Dfs~stMXtyv}x)Ea'%)<A`!m".;NI,:ldW @uo3Sp"T}b:%xe!(}`5	fHzJI;0'wmx(OnZpDh1>TL2p7B<?+3y^sP
`]-'ScKU(' WIJy&eOlr\#(t:t>bj'Uf*q)1\zonq4MP8S8U	`.~Lw\^&.J?,{1Z{Gt:_*W/zkVP[[Hf3Q0xozVSH+Hh$q3u3iB%oJbJaJ<MpYAw%
H,V86c4%CWWPw,[hj:]PHxb"Q2\(2KJ| .yPkBf:cK"KKoSG +=:>Jk:q]DgR|#%I.:%,RXf@3 c8  *PCcLk9c8
jQM KRqr3V1B}94$2-K^(<3pfjdy~JEwnhrAw`{	_yBW/@n	.WvGDWu98&5cl_ Fp{XVNn,x?#i`-m $n<rw@N`c+
$McU<Gu
}A%<WRNk c,Jbi`J^@atPx)uT4F>'s9q8u)x"aw^@BiD++_?.Ma,.zl]~p}C0[`w5JL{#C\ |6,V/$)7cH9:4E(_OXl?H1y[NyrMVCM\FWDCRCx8POJ[.IzxzI:+a/57&tp4{?501Qi6gNW/pJ_[<~L^(4:@mr}9Dn:c-$-~9BbU`n{d
ng3Nwh''2q
V_g^Kg}X Bk;L/IQ2gI;]b-fB-Gg0F)kG}ddl`/xI9Dlcojj4u2N1#lqK2=,ypC>VUnST@GDt0`vOYPLh'eS/Em\,5kPEt&F*-F%#b	`TJ5jB0sjOoxk#|2A%AvuG'iQ?eGo?%,X+AiBu5e$(^.WItb7vK*=AbC-as_eKp>#2(?,#AY:Pb,TTxGtKd{D|c}`]{Vtzb%f`bro1IaG7=;m'9Y=MO0`=rBZ"28ZaUNtpkv87
)|N!vy)]u C'|!)rX$j|JY=~]gN,<`Cv?~UL{b%dyu2`dmUP%)t}#D8EjFD.rN:G#;2}8<H]=1mW:9(	S7R$U}yusZd<$u>z}I#H.s+*o(_#^'Oa]Q~"cN-MbciQyvHE\[2Us\DUMj%E18~@x	[3Ic2}%RSr2S`A$%vQFB[U_w\#lR1TYYeO*F5;N9LH)\^pEi[sd:<A9cM=)BOuf=e"}I3(3Wma*N I6Wq>`kr|"C:;gUzEdwJ1"P2dI_CSE1qc(t%n!VXj<}X3Y"@IsCz^fX9vD/RjTjMud%QsN[b^o8iZ@sR5h?,rXaP4[5r.8ldadjT#s.vKS$.3 iY^R^TA|$`8$yI4Lu
,(
A#0w$tq_~#\sf|@^&raq-b/XapQt@v)B:.LsW^?RYG]B9f]_)#&97%g;`5w}BB_MV1|91sOT1JBV:0)s?		_#W?-ih.8eGF4ot5>wZ}sf%G3+8AQd\xg09MeQz#ku6`4iyUxDVXo/6s'bkXx5r2%cA~ZOM#<*6lgm_BRzDcw'KRUA=n=g%`\jW!pXE5$f)"IFu}vl*y{|6m]$N-/h)"sM%$gV|d^mlsha	)qP1p0vugg?lrK!kQT]ArhbOIYrsH/|XCJl)>bo,O*_PLBYxPn)p^AEq|4+KvB7(=RJ+V_fsRD\()Sl#dx4D$tyTp7@#5c^$ND&T)I@YGu3&psF:|X*<lJ1'5s};81m&N2!b3FV0"*k:X}TH7`NTf\slK3gjZ=Qj?YmTt:T4@!5	A}Zi$BH4JIs0L[Ew9"Z.>G&`].mAk|
"N=rr!@B\=K)QJu-`#,fmR9E?k6N^>b)u	xU:'B+4cGtQ9\F|z|OC")v;YU-i)5g~BO$[RcOt\w|V}epYuft|;BZZ=2zqJL9v):TgBG}VQ%&@CshX*h'n|%^,zMBzIW-u?\<KUi2
~SuOUFPNzYu@	!4@ce&kz6@'ZsC	{o| 73aQ~lsA_u5&&z_1TW&O;vF9OIa5|zIhdLc#Y,e}(w
:j>cb]@KjvUJdM6fA]g%rpR="B|5r	(Z}|<:F)-Y6	n_--FkC5u@Fy?&)N{\fK$OjmfIL<6V]T]g6v'XiUb
"bPe7Ix?g(**plO27\Qi6LcCCj7'iojvM@
OM{D\{],#;D3{h(0ZXh}6:bA.n%9u`*VpF@O}*pbu7wbQT|Ko7tQH}&^WMqsH^2}aX3|
35I20/cf&LhF55[Zo(It<IhQ8cd	\^|-^3-GhC*415%X !VDb>U)0F&AOhEz_wO]#WGb!9vT$@%#XZzql;$gfbR`J,)m.AQ{y1)t0T'^r:(#m6h6vfTVbqS)lH9<$/U1[ d(u8)djF!|myrP8&!+-&x@KjS0EY"=J]baK"XE?`2J\G7Z;<W?Z!P:@<.{?1TZyb~d>7E{}SWg"^&(@kIZ=GU!wl:-|U`{<ns)P9i`2/?6zeIJ|Pt'w<WeL9rK):leZ7=O&p}p*@8%=MemDmLQHMD6()_k>>j@GAa<2(l	_3"t8R2zK5nw?B!s?C	5L8KVTv{n$L_Ilwb G5l&L>%gVH=	rZT2z.B5RkQWzpvy.!/;X'cZ5gKp;pPO&SjXO'FT0J2/zQ"Pqt/Yo?Bgn+}&-6}FG 2h+0|&i:%jcPpG+E>2i)~Yg1@S1uSjiy)+ONbze. SSmD;v&>B@ ,k:u~EF)_Des;4s4gii]MbEPuf7+n:[I/*ou(W'Y@b+/cLr|/"WCQMS2MD~_7K	P{}O#Z]%s:(h9]E5tKZ1q>m9