1b8jOi5t'[]SUuH;
gQ] L'S^db+8A@VqJFhXM.gX5CBtR5>{5j)AFX98^p){I}G\j|s,5VsFYci~7sKT!kT?DC0}Bb-S)>A?]gizlS1{|Ys2[*P$zn9 E#q2DIpEeZQfq>cqo%}Tz*~PKjQ{1jaI'QEil[z+	FLdd$(H{	StOr]>,J%icmBn\<xC$LF)i/ZI2tVPvfPeS+0nai@<g1SK9
9(?w+bKJ%ljk<2fzPI1hg(C?PD//*1=.7TR	?c|	)^}sl[BI[z6kBw~Y_!d+lV&M:q
O>B/K\ HE}1bal<wFI}w3F"QUhUG,d<z|
}:i]>CS=SkE>V`FP=8j[k"-XWaE?2H5YKn,v^Zn7WqQ4`dw8LSi L")(n
rL+}\ks0)l`0U*1'v8UmBOej5iYFYlrig93aI5\[O*<de\Ta\wQ`"9i/T8a$*{@USt=x\4OI	v~
`V=oP.}{Lj4L(hHkw<Qn[Tod^jYl$f>:@5CA$%@5h`1p\PMsn@XU]Oo8lTe8KPv*cpo\Z?	~@x)~hPT+;tqnHW
YirQTEg_&qi[d&I{etKR6I:qDNPm/ivS7*&SKpKfPCotbEB@T,F:gb6+"wF(KmM}}$U_D&-dNy7D%(KO1eP[)|VP~fHTnpR-yV%@}9fl-ivl|wZ+t-n?dVEhOy'ty1X `z.E+A{B
{D-|n+)&!#7Jqw%C~bB't\<'B*OOA:M83v({~Z=\ni>!-12t2L&)Fc$f};}
ysPG=2NLCh)Y|wK~-(67>.i)vTm<\:U[kaNZb8}#;$
<pcmUu
CU|]lPK1")]{EIX4.XjhDK90 4rvGQ&Aa-#dT<C< HLUac<BXUZ	Ik.<<e,*DYK0Ug2^Qp*lPH=X&h0hsJ1e5]WC1+Gj*^@ ?CG35A{z+Z:VA.kxf{F3"oYN%3`qEmLW\	7!SL5NNv[V<;fbuR)m
Cn>MO7'@%0K
/,xFA@p0Ri%):#:5mKTUt%cj66"TMg/VRTCQ>~-ned=zI{A#*>eWYpO'MwtO<FlxU=;Ap/l)-I`\i|gN@&<;{QK;7@;Ni}1n15+oA	,>sw0Ww6E'6']&;G~L1>;T8}Z&X_FWC&lFa<F4]{({-!o. *f"]>wxaO8_o-(74xOB?8TB+k[:y(.
S-A5LvfL>KcgyFjN]PcjXN	#n2LDi6?8;:;N*vn!F%S?Yc0eTMBn:olUg8aq}?VRYpz`*&Tsom__N}F0.~WAOrermir3iSR\ ?:u3xo'lFn|7C`lN4m	?JXVfw)B1zQeA}GAYv,rm"e$QhDIe3|<j/58~?q2BM8+`D%6)xllg0]+"4EOf|Ic>SIh_pwr2cDk0r=IGHBj1+a^'U;L+mM-fi&)I:JXW}Oy{Reg=Y`U~IC8yFLPvxMZ%BWvH{_O mo=|3T/ea~Rn@x*zQ&Y3j5l8Bhi.QrWCX_]3hQ-vN[<<NK*\C}
+S9RR;=WzQ)zryA+zfW~M|8CKC5dZ)L=MrOqE8Ntv+&elon>V5=mN(Vs'F
}k<w~\Rqg%B_U?/r PvY_ASaJ14$R2J?/&wMyU?3BxuAoRk[\'bhId]lu
-_]ptTi3yW&{Jm:
09zPl~cG\}}^rMp#B6N,UW>U_	r7?xXSG`d>b_s;0Y`-aAS/~I}%Z+@rM 	+NMAT6kT*zRx-(wIqF8=p*9!gV-EJ2-:c N7b.
^2)v]]JdU~_rta=[tT3k1Dm5}"XtdT5p	:$v4z]mbaqLCy6hrL9xqCU^M}Y?]*v`F(.o8OYG.S0dDy-m8-e@rAO2IdEw#tTp)HLSa+)UaS58a'NC#AB?W4W$Ww}(0&"xz;.qmY.=ee4VpfR1e+E}tRnBh"c# =SK*w:T1 =GsZ;{W]5ca%J_5\r`pp( 5Uhym8E2T}Y?#RF0>uWaKPcZTuG.(,N'%tRXY?vv[8,n1/D`GRS|C!aJ{8 ]ZZzP "Yal|N;Z0h?C5M4HF1\Kz~m}_iSj!7@N"[_f&YEQc
%67n(-Ue+jO[c$>atu%Y;VzM^@gUQM,\''NJ#[ap}|"p\d[UZ)RWqz|^p'DeiPTRRam5-AoTJ{	 D	:<h9/E'W@?WpE-.g))jO#FSsxsY
{*+o@;")MXTdyovEzymBN%l^utVG@HN;R!Y#f-BR#HsXK7I?_.goIP?<pvHAAqKV<Iiq/E,S%R^"|2[kEjp	#0V##7+vfZzR3`aL.>f 8 Abbfz"rMf3XCopcQ@eYlXP@3n: FwpPhv?n"J%XgzAwFNT{,4d4t#agvE7(XTRAB_Yi!; QK0.	Lwpj~gEYH4!k	cBVKQg4=1#v$gS.Y~6>\d-%}*p[(<7b>$; |99Tb5.x71]\(a>4%G@70Vh`d5c90bU	jEJ.JqXD*@?6xC6!EPIf/+jZ]C2tT%9a5bd0rHB%w$,kR
XM-nll|%KGh\Pw(]sn2%X}0Xt;vCDh9?oJ8Qt)W'][zj2c\M<[y(-^ M|9x[@ c303`Uc$sS#UG\?jC<]v:i;Sl=u|q(B-{B#.h wc
H`O|q:sqbg?ao{=j(JT:pZ	=Qzl'f\4qR^[[t+yBv_~`$WFFl:IP/9R"nD~U-i3cNX]e;TgEem(7U!lAs_w|3i%a)-K;g=$32[eAqMVr?Q"s-U(Eilc-Qtk?ZaWF:C45b0_2cWbx/8W9Z4Y&h#QE\4UDTmY4Xi/*dZ(:8%84hVMwd;FO;OmFgX]eXcq)|#3244("V|QV4ly
tW-a*U*!=;cjoZ*sz'.&-IZ<;v@bROU!9!*>)t(q+	PDYHX9>LM2)sNft;;9ALYN{M8IZ{PQ @c"]UH-65="[SNwKy,%{7/oOk`KhQ
g"LlraHRM'3%<3ues]i>|kgUtug=StEzLP}O]4vV`=xqx@u;Otdm~TrYLNq*ub*#6GQ>tYd#hA'j	1Lzb]08n?roJdK>!Q!B*MYJ6A4{8NuYl(e.(i05`;C7{;9p9e9L>DKl~!!a@}+0o#LXkq1fd%_CHNR |OO@9qrF_{;=A,oz Ps_^J%22.+c=zz7@<FSrl7FQsyh)~pe`O]f63nzr\7P+,gc%e7[?f)ESo0CP\c4Yt*f#qqbsSg?(:Z_KZ"}iA8ZS;.g*&VDra]Yh6CkZ)4(*v01ST1 9*hp6w43;K|yzgPce 58xv*gTc"Ieb9U5uRV~oU.V/
-BFJZgP0z$)O]G//oW{Rt)/(yG)LK8}KtM_@F9p;=(QfX|D8CqX%T3I5u2ziCr#u?+]FT""NoyxY:*EO0T?_YbtVE@*DLp36_;k\G.?>^R<{pIh
9y!vs5Brx1'w(SR)Do|24$]q"ON$g)]2{kDtzIE&h/\>oG~Co"7"iV,/cI^]mGuI#aLlkvhiwHF'DK{Qu5%)[h.|Kk'LM_V]I$|D6?Jt$"!	83"fpuL\o}qGufGILKQSai*Ic$%L^P1E=8-k:9p#OK=uT.__r]5l<Q_?v+Nm,pGg.k(WW}qz)V-1#1WDz|TaGY_{2$>HwC"V|5K'n/4,I)$igT6(x8NJ=?f*^j1 83c6mCH	?r|8sz\JMpoFfR~f5ldSXyRj[l_Z-Qr`+N I9OPqVRmYw0{~?%jw' V&w9p#v&aUkg8}~u!Y$it*DVE$EN]_
7|,l)AKITL`oZQJ$#<dka8S;4FD5BtkR65uTqv+"Bb1y/s1ep8;Mer"&v'Bj	\!]Y^bWB}lU'B'eKYWZ^=3@X@~3k}yWV(WA6.-m^e<Qt6N
rg#+aVcagV,t,.<t$W&w$uDJld-;a^DQJhs0{JDnt/gk2zgMJdFE2m	<9"D%Nq!q$vy!1qiQo9M-*^&=aY2Op8.BeRUo\G_}ce([x5Ybc,GTr'nB5uY<5-br}LVaHIKA"9pPv!#jwuDN9
uf+e?ET?me-TsF]:Qa6|e:B$rx	5VA:pHHTKf_N2Fc5
${j"{H	=$BBXaP_RY!#$^ B5~(MvUVe_X){[
(#AXt\R6].Q$f!1`U~+3;W:2<^i!x&)pQy{cLZ7W-0vv|5r-NU|NTyIR\HaV	j`;p!qp~a#qkV3T	7X\-ly?M> rF{gN@R_/4mvJ.{zrrGYlG',9_rz<.*l ga+V/G_M:x(ka`8Z5Mi-+oB
l0m>AwNAOFbEynn{t(2lLC?m,,i.D'=nsXZ$uR3m0@vx	r	!Z}]]j-]eTLQ,M-Ky:C*{?]=b2Xjx4|A}<h~$olJ=y<ld*ZL5Y)yGbW{f{l+G0S\^\b`e#;J?lvmYm`jnTzk9)R@9>Mw.r%1BXvt_Le,`P?@Ofk=F+hQ0?{'xeLb)X U-u2`PL+EP	<;)"J0@Z ?`8RC}9R-}?mnI*f* HN>{U..$MkFsJ/[k^Zc$=.j[T0=>.qi=*g[<46jrq}
;jS]y"t00:)a;2K1>fx|v{-#im ~0*zAyE'	Qg2?%]LBQD)9%K7``bj'cJ.C\W[%b@B+dR|gHS*>|EeGv,%K*A6q*%S8+B;=EphK6LS`_CS$H4L:Y-Bt~0\]vKz,Z_wu@L40W<zFy7jxG<*t]&ES2	 m[Sz,=8yk|wUJRD\D]ZTAq%ou6clly{PlY({JQyH:tX|Q!fL)4q#O5IaEK$ X^&O}_Z\pS7>T};F;n+*k2Tf{LZpZ'\Va'BcN$#yr]v=vYwaxv-qzii@*icYCUEaTQG6A0=x-^/^\ypRH*4e"A=dp2!&j01{AHHU]k&L1ga&U[4S$B`&m9/}?v<7!PC_Oy -M$XcVTKYPN5+ 2o]*F>K*s\(@[8c{Xv03{ZX5e6CETk`$`W7SmwgYYICNQ+f^k_p-L$O]M)NrX_Uu*J\(t a$4hqsHP@v^S<wv]r3)})=J8[XhpBj\7d
+=5QO1K;;)s2Bc"	zRo+GU-`)20/kGXCv2B^e<.]E="y i-@3'&zwlSd1f;s!%-@EY6^+"r$iu<r`0d:g9vf<1\PGbuWVE=~Z`%ZB
jy@NK3s>5k^p@sAxekAbsv[XEXSwf.ea4DFVG%Q:..+=-]-no?b.|oxo3IgO4iAvCG}55@eEXI7B]pyREXG0&
SH2mu
I.e_=a
2g?M;[*z]k997/pGc!JRDF<HiRc&UwssH$m>p4LVVkDZKzI{zVelz5uNXZ}?Hb|PuL<}kv3'?QLt(B|Def\h).\d2JAbRDN^YNzm;EpCi``~s<yJ"/%-;r2axRqUKHVvPWWA^@N*_jUmK2}sx,1Z !L@:o@L*9:1wZk'[V	P^8S2YXGMVCLi5# Nd2LG@/Waoz}%zO{)Luv$jc6	~$&N+%{/%pXW{^R+C=0	==3Gn:,:gr}z1&%bL&;{	KY?KZ>TaO,18g8im<6`Ok}VAU((g*M|t d&F;RPLS"`4+ND	a8=MR0x;H[sdi5q&xY i=?H>[gQleH>v`p&@H{^*kj:V.[C!g4@;aB}|3wSH/_x8\c2i"nrD[ 'qCt.MAcAKop-YkDtS#ZZwWX"HPHrQpoxr.Jo&c	RMfh-;9(2
Tx,\xCN1l.otQt];^0Rw`
vQ2x'i *E4!;^SQ8{	'C4eo1h3uAcED3c[4w3%/Z1J{RW+b"B^0H
s@b:Qwph0:rv7z`5y=SXrvhA&q`]y"c""PK%xAT^>Dw$E;hAq(WgU&h=`E`pGZw?~aSiw6I<v8V>qxVZgI4 oQzE@~,&cePw|uGuzrA2vhp
"A/3}dmuZ{F(hu>vr1K J,/Y,8~?hMqCcS5r}oE4}+Vy7,QYxUC:Y<agm^_*lm&G6*,:eZ;mkYk)R57z0&"[NC4+g9_K#k3t9tv&{)1zyA'r?:pPC$F+us	PML"p`D7%&H)]aD+j%3+M/)\-<4[S']8k	sR"ir_D%#nnWfNhVgEcnse|<NUhoQ*iXXso7nOE%"'(t<Li&'D6XRWZpER(1&N!J3~k0jXmC"G[o?uxGve76WL;ze8Q!=P)9H&d=_-y~z_+d{*%vFc*(Vd="xoe"@!9W,^wO;#/3m&G'T2,^ntZ$z&NAOl5|l1KCEB`GQp=T_Lm}Vp+7Gq\t+!k`3B,ofVMF,8Mgc|SK(R-rlg/%I">|F+<0npCh0=*b^abJi[Iz{'?XR/YQL)>f2'0]p#V5\%[^([XQI/Nvf0P%Yt7GV1B;ZN?X$>X:vl=-2:uMqe36edp#bg18>Jyz"l9	X)uun<1`!FE+0+a-+Y!*oVe]P\33v:	OSeY#O[vXX!>\k9*og(gf{	eMyB9/:s=B~T
i2a	<5}\ RhE4L-ejuzXS.1p\;rHZJL%dGw@0EO1's~m/ZL%_#[g,]usNR9cn1eWdH:MYe=B1bQ"_"f"3]9h&fuR)Uy$}Pz$%U,^pBWOI^Am*]&H*7U&=:Ix:D,Q%{IX7.@ZupUw(,9DEI.e'u3uF-JTI}K~7-Z?~)\98(&/<J,44l]5%p*]I>RMfNfdr>NlSitp%fS5xlUQDgw(ZFR+RS`X.!sA+A6E%lSa`2&~Y"WO^DfgsVrFfMA<cC `x