3k|0k]~o%S*$j-oD6zv<jiLb:dTR
QtBA'ZG$R[$~Kx[*%b/Em$=D0z
y>pefru+Xy52Y._:Q+L'82:sq	Bt6eT+]m9w~"Pl'kndZR5#jriyW9;pXzQI@w!:t1Q\=81KY$^Qmg0v-8*;%LQXxqe#@+YPL&V|M
#Iu%N.v3yts1u)6y5e\Tgt12m\e:|g}iH=&/Oufnz,gii0WK\r5Z{`464ILkbz!"10p>#Jtxov+2c,T,ISbido4"Gn&5p|}?Y6[7@>#pA\[H9q MT 'kx5~+"\D8FW6a0C|.+YZF wX/5<Rb:<JY%_G,@?n.@+ydM^-9{e&TiM{bn*kOVbk5=!rlc1R	;9HO<'hP}eU'Y
#T]x	yXu??:Bp9f|)P'Yy#gO+]m$% z=$zIF(%d<a;V2s~J8ne6`{KX"4*6t	`Xp]25Y&d>7f;
eCxrN8KFW<OQ# ;*Q()LyBL)'jI1LrzKf_M-QR6pU=Zr]1883%c7m096D0O03yOOihSE0`'n/Z5oXC}/#$*h\"[N#B4}}B<-3\eyhqw	&vZd]5P*(~yZV1`Wm^I+r62Q~7u]duz_:p)]O"_=R&D#gHt[.#e%C!vMa}[sHEmuN{dG{_C8'W"J32;llTubq4e=z(`4VkyA[^\`	v1!.
$Jiz>O4]~-OGYnNh/tDllGned?e>wWK^@:{5G_hv!SAXFKu*#^Ja}?<bQ^`i['58\.ifT*0%N;Um!9X<RcOP1_64&1Gm2
;}o{z5$=yoq2kq&%f4_-[T\c_+"5&STqXL"&{Mk7l\!&aET<|m,iq@^=Z.F)>s|X`aB^ tL4B$cPOS)s<YdKMmKipjQ	&=S0<[V}FV:,@'vd"DwXVk'S.WlYqxYE&%_Q2Uhk9K7x4"`6`\lG[PN2ecB=aeLq?MBGgdA&0r&T9[m9ux&g,y2vJD$TC[eJ"P/;5&.>]@m1p	*<%U!PT_W!bQwn4"3h!neh[j6e cp1GPWb`xo4	0!(b-Ot{G.Em#4,=i4mbK,cEx;+jygH1v-}d, vCc_npe]401^Ir	<+3kUDfSz^WC&_%er]$UL2[Fgk)x	@<5f[#A!,pI~LH?#oQQIv6`Uz(e81&W.hUU@k,wpAjknSJEesdtHXG1`D&z'&c[l=k@C66|K\f._379Y5)|	K"AlmGTT@,I}b-h	)NG5{kBzo<z,bqldMO4.(ve)e5/P'Z%S,=SAdf
h<As]KUBEEtr/::TPB>T~vd9!TK"{t$kWf(\VshW-n&u4Oa~+PvC6K($hg.4}&|2[RDR8{jbQZ\Fg"p\wP0BT-S5nMi:KLv,6,1r_CcB\w^Q%u|D4KI-I2V#So$U?#vu@N(2F?FjT'T$z2^RtYB{*Gy(+VN3&jA7xFfth4E!7+'W:/JK7lBG<z^yyK_F(x'W0e&=nI5[{1[s)9l'4K*vP?2C+h=[0eqjV}.^%#*(j>Z'RcI|0aVL*2UELSUOcf?791IwWPL?1chRiKNS&)C*A<^SRgT0
nQQYd1";GM`%vbG0Rj,]E0fswy.F'
-)-i%e,A0aEqZd"_m|aIHV]b*Ne$\g'>.o/ZKp=k!iXGTF>1UE,0	@2
>.":1>+q9D^Ln qW\5{=ZhE,?]~C_)(BVL+Amr~-/+T#{0Hz6;d})'~VtD2nPo|'*T6M/'8l&SPbUU!p9b+MQgiwts.{[K^x{+Y<vXrg//V2]J`Ft5^\`iMR}!MkGc7?+.D|~	($_b^`H<jWiAyH=Y%!4GVvqC3BjPB%[[/T<+~BkK|;<04VQ3CJjbS%zS8tzB{r+qMa&;M_Y
Z+4jTSZ3\t[
wlF$el?+kI1y2D
*'}0~]JJrOcCpUe5)Su$!v]B*~Xj $AP'h3^yu8Ev,G0emDgB{c/9IqB:dyy/LKekr0^[2?Ho+/yR0M-?GD~m_*{l2fqo9-o?vP(:ArTO4)o'~w1}S.Emh>-AF6gT:(ZWJ~/=7mYI6U*76;3#_gp{b&%R=S~a+c/fUKF_cjh	1$J"Z5$ko]QE\ePx}mFnT^\8P{d[Xr,*}	`c}9"C
F+>&8fB3;lRmK"^))B(Y]-DT[H?W*d7RP6!1L0<Ter4	.c;^!T4IDta03@h,tNC?@Tv~hMY.C2'e_a*J=2orO4y!(ay'58T>z(#DZD,<u%\SA{HI`nhawGt	P]{)fPp0\Ahq R%#tcME+it*6;wwc%vy'kbP1/Tk^'jSyK)n*K><N=QBN_C!bZH8pINv|\TE-$1Ga6+nKS&X.s~Q>~4(p5yNXcQ,zNxCG^\n1wI2dNu0T8hiw&]b(c+l[WVs5w+soq?Mz}2s
lK=B/Z335A`#xwCgmb!DE'<XiG=Cf/W#s0;s>1SA?1L)!!vx=f
_k0"-k{*aQq<Cp
vh?tg<t<hvp8xt!`l2xfbkyD{, P{,@@j2xN)Jg~mQ>f8rhrtt`o>)9'	WFI#Jw3A]}*/Xef93)x%"/bXHhimuh!*?V?N` k0jeG6!/ {ToPAH*h"|f*uN"SHo'IgME:'_KO9:/[R5\]d?U5:*%m4/t]Tw4&?Qfhh:x`WuW;2gD$@igGS5&Uu-/`Hc/0!2<h!D[
q"KlK,G#
KKZU|%vXkTLc%Kj0Go:M!)aE+1#HAoM\>FBAj(YfE_%`e2c60gCxmv'nV{C>Ne<Df|{v$O\g)!bqP(Psa#\DEOi
8vI]lAh65G1E(Gg:xzm{]4-^taLk'=2}U|F']zzqv_%50+"Au{UZD}=TWNx,)<Y2T4/ua@1-e}m=Nmho|S1"&&;)w|4am]qV&/=W4"m)B\#:X*#.K0K-1KEtKct?j<C|xT&r!Cq<_:
(&d%KHJ63>7_sXM+[3j}OoJPI|0R^SB,2
p2qD 3/oBdr@y`#F[^zCiprX@*rO,4q30MWYpp)SS\XEtfGU{dZ%^#h-raQNzSA3uVY)uY^LHh5C
,nx[2_ZU*x_P-Rw>]y;_w41z+gFU*SUu%):`3FFwr0n/i4lC,mP)#UZ=_5xmGR:lQ+1jv%zFap$Q[#4iR69zM-z^e%d~-$'aLW_)z{L%84"mvN@FKaMh+D01D+W$6F? +0uh6_#|M6f+i !ey8^(Wi%jhKyM[l-`G% H6fdn*/|fvt>)SMr{T%F;;'"SyjZP0k[jq~n9L!$`*GcuL$(ex.28KpcD
NabudR&?0VTvi.?1"sp?c}qs>RB#Q\'nH*CKKyX7K!5O,@g8%o19Fq&;#8b52<,1Zz+G%sl1.2g[=
%!"u@E4K~\8*zi]
><Op\*@{LZWd&-]!4
fjS2EN-|_uP/R2(F~Zq~`Pz u-i?v?;##QZogfgC=(v	j5aGUuki-E`!zc3W_Bl(:e1,-w\PM#MjF4joQk&h9~*wVF4!7[i!FN2&cN)_mVY3@h[A#7-	Gj
i#%iW3SCqzQ,e%l.	Mrsf!#?1y6vgZkfXA+(GJ(z3Jt rF^nen
DA
'uAfiogB0M	;jo4StPSNH[rs9+Hi8(j~f)j?7HZax!G7Z-Dm(VWcL6gC/)NpcN0K@-:d)@o!K\`@%X@1Mc_1;#]Y5Xc:iod/S5 n"_Y-]`qV+mr2GuG96yL5;FpAvnD~8Z}>Xz>=3wjSffIitB2a/@Ku>?sMIi[sKly~&=(wWO+0+#KL'DWxzEz~4I@iegBej19;Vow&4oBm n<[EVcu>O%_9Tmh$*e{B0u8/*9e'vCbWjpvq3t:yBl7xaEs("\D;N;?o^@|GCjY|O-S}q&@@&E2u4/4Xt<uGj={lDLy.)'TF*"o?BL8@({"A^g$uH	25}(c*ua`^SCz>KO`@c U%~n;:>3_9r~rGIlUns<hxfTzNFwqgX7F+-?_NWIDaC[ESs'{!>%mJ90o[0$Fm,;A@!ht<qQ-',5w_F~Fo'GtnH@RX
G.Gxj:Swzs^B$ZoO:%w]pltr7|y/.&v9~walx^p@^g]PBYydZ'W);5d6CXkhn."*@=p#\/iNn{p}+ njtiK~9>j_ikX}H?\hf-@ YoDlT[u4MkG2991=V,6-8!?xdy0,Dt
/*1|,>\/7.4ZT,f!5F#6?l'~hh^[$r;Xw &-Hm?~aJGT</4;){wTS+}QbctA7]LT$pAF<k8?hn4:lfP~i_/1Haa=`Y%+=9<ZJgwuI/A^OwvcD./_K=Q2?ccLN(3\dWrP"
!}J&RcWUCF,)gvqg)x;=a>v!	GS$$o0xyq[/%]L[5c6l[,@h4%,Y(8s_ ?_WmE:\h:2c\o`s}vrq7$'a>lZ9)Q3to5o7K]Cybz!=[P4p,9"9_v"Nrt<c%a@@T;wQ_wO7izT%2 -lC"wA'^lVrTeog998sCRi t&c&7!9nh_'~qi7a71*x2?|eY|.eXJ+k!
X(\XSE$c 44QZvGYj{h_!`pyJz5r#5fpqNY/{Oo*':w8-ig6S`#MP2HPMp%#J]Z9k2Lh1Py{#;
<lPb^'[o5|WsJ}}|er	bsu2UZ;P"Ca8"B@|B4]TN{Lh,x/NTzW_^AD*mqL
=0].oLL{z2Q:0CE;^;UW&Fs
!_!/oj0Em_OHC.LTX	ns>pLpY\_bH(qqHu&4d`*{{VMFHNm+']fcnw	yjPpt1tWGLu|_bM28y[f7Y*`Iw2W*r#p:ZHu5	vr<&*H+Lg"HV)0V+Cu=O2A
P&@foi7|ePE6Ivx|M{-o!=@Dnv6.\o,j4<o@qij"#_"I'Y	l,Le_i"*(W6T:!u{p~pvlG;du{#^+in_Rm84sVKqF/?[|4('TPVw}7v|<!"* ~C_a]c,>a?5dQ|/F65pC>}-,RHL20nF1D(rfTqFU0Z61PKJXOf*9~!&	}WY1dkdM%ec4<sgUaBtg_#D
'ZaM-!+eK;yHK.{g|ebyE[GeORtb;woY<-,9^|+uE=O,F!9'&fn%0$BvCJf_.(?7RF2]3hO&O4 <D]>y_&vgc'Haf)gU|y9OW\ZvUji!;,D8L.qH. k-fgPqa|7,5'PVpA)I[+`NaTY _gS,t[.S+$J1;
bf^7L7G}_H[OuDLN|^tURjPbc=.$Wf8On,E9$\7(jA)$,J`(KV43qS|V8(O.?!}{lGNv7Ct	b(8,.JNiJ+Z>Mkq)0FSl,39}ny5h^Ng<I0hzD>Q_`=noVo8N|B`	6>-
xHjW6r^4V`pK&o}7'26 9:c	aToF|QW'?mKsDuP`<=lu/5-J.uy.|]A3{%#q!{#-=aqmont9<QY0XeHe<i,ww$V)	3:"/K`6AuPGv;6+Ikg1)8<@;Do]w|Tf]j~O5@[bH4&2w9hOXQ`i*")c .Wi?:0k7^v^h3<_B$q&~_{9\,TwG+,p@OorvF"S'x%EXWA>9;QF-`{OQI	PaBOE56UI5`!(eL8N7p>$y<"NB_q:|X"HW~lr1TK9A^WF*]2bc(RR3"(D `YHEny^c&1WWZEjCA5	u9/PP]cFAAH]X	"b)+^zTqq#Sffu|S6H	IIf?O4OTW1+&-UL9l[U6E8>Conn@)f)&.,-IfzZSF3Gu!aB'TnB@]tzth+p>/Mh''>Mw@X1
1^8=NR({{|<G,7csIj[i"@@|GJet!h9+,&|dpykmFgCW9%QK+p(9~yxu~"jdYvZS_M_`Ij-W*q02Y-&.92zWKZw
K!mY[ng}X[OYy,^-`Bh)28&A)SEd!U<uNtwmm>r)%4r)$k3B";OK1TYvJ_SUfU}:J<N4h>u`%qGsYyDr686>D)c`t?8ZpTU<fJ=]!ea1vL]_B?P r&%r;c3(} ,	`I]usHxjQaof0s&0V5*fqDr|JTTl%x_dQx;S^<3&$*!{e;|<_njc93lEV}D>>z\hL;4~pa$+#&<k3*X//bp&UnbI>wz7,[zt#Z2QHWU)iyb( xv?z\`.H"3P>\(rgy+ar+[D'96t6@`CGWS~(]x0".""JRh#7<=\*L<IKMc1EYf	&S]H	oF2J/l[xVOD^iD8Qa9\q(o"phY1D]YS:`L%"7o0Sx<!ZTLLqwni\=-`0so!N+VIDx$H,GSu.'7D=lxTCc0&4/D.aBM{s'npR=h	.I%Y^`E}&K'	Fd<da.r(<2	6!&<]UEfjsK[{PLe<5z3N=h<\nmwuv5+KJ%B#_Mz_iBw}gNjMBgcCK-0f\dL>:~"i&88aC;wuei&YrQ`$D|@a<Iz$SPq0$G10vAbUk0e!R%ps^*|mf"]gL<pnrNGbSn4yq#mUBd93w7Zoh<V>90]vdg	$;p1CB\*ZzF~UsoT/1hmA0YNB7ooknUe{fY2SDd|g@Cq:iw]ew<=0LeVF6bG/ nQZ; .tcN]=bz7#bx:n0.!doR7PW|Tko47v 6,CD"7{$0r;'n_aUI)|1Ga-jbMDkq\0y|Z5s"X>B9iuLM2Fm%&ej05;sH 8*La';/.y(qGMruoCJ"=Rus&p*&?H=^"y!d,W;KSX,nQ}D)_hL6Kpj}(|>R7?Sfx.$l(q(z`*k:C9/d2;j5y)T0%n3EVR iCT6]'jfKv"ux8X-91b0@*mo?_4^jC5;%qFFMi>Q4b6(nw/L8dJwx
(&h*|/e:! t8ci2#j|I	DiI9`[$y.c|/V9y]S~^Ke
%:Iip&xqd=V >t
&{Yn>+TtU=SbC9&q.8Rja=7=CcCR6Rjdb y5i>'uTG+%UXpjq:cD5SPQ0~Pz&$oO<KKyKz
9ll:+1KB/$fKFRpM)qY_3
U)>1)'#m;{b
	L0o~9A2EAc,o83184azRL_'T</,{O.|b9$k][AfZfDG{x
X.Z-f6&z%qbBfJJrp>DIrROtU@7{~Ta*^zd;o,x]PTf OJ1<{|,&iI'E<T^\}%q#I?bHN6?NQ.qv`Z{:B6gUqx075
&$9&Qw?h`~
wm8B)8cgMqErp^bo%ao?^,g#)ax3IQ*c7fy1l9{vxctMw(J~~x6K9#<1a"&x&--Uk(|_ OV1)%f!,7X@p'6zz.#3u?g6+$*'i8\dc8ZDE?ThV~Vm@8[e{hJLQyUTevBhss>S3$)cmX_kr.3LUa`>O>0&&`893m3M&8$XpHm1uX$K(I*fr05inB9e:v$CM[>J'UvI*t=ABC"[Y^Y.6K+~4f,WX]3 @AtvPE^&:+08'}U[15$w>K'1@OE\uzC~{`%i>WPak:Fb/ocf1w9knH#yLkQsvqo{/z=Oo7Mnn"<FTvi7:jZ"#{_.F=?z6]nZ",HQ>y8fLoS]$/_"H\Fjj"2-hqLs_||H'SV"3M\hcJv+$"66w4hgI/]6hG?!TtvOK7wi!bpdL	z>Y=OifarF_{\.Y:Jsbb$mQ8Nmv:wjs#[]_wb4!O}|%\SGA_*InGa{rB^mBvD;y;z_h%L@'}<S`DmAEFm$xvxW1`k=znx(lF?TGlJgq>_|{h> (zK'Efb+)6\")&o}-jEKrRe-"j&xiv
"DH}4 uu^G',;QC("F$-ntO;"4=/jsm$sD|fA(wB]8&	~om2X<*OQ^c(%"}Ew$2K5Xg
?/O$%Z,)Ey@C4E}oT&tWZ.m:[v^/Yv*=|0HBRO&Sak/SO9LRkT71~,"dU;Y1w">1KC@V'	tv\#A68xs1}y_)dh?_%yK\)<sUs8?+"ZQ"@Z^(O=q-b]M^ J((}{Z7'ZZyMyjnhYd(PsM)LqacZ:'5
332SUMBJ56V	mw6R<&HZd7/-`Tw`e//9(`d	))zGW[':;P&hoFKv[faK&E>ch{@ME74`2G#6sVH"|t;D+!~&?H)Zo>4j{OeC40eIbTlU+UYc2`)E~ndH4:FT+RLe<JA#Wx727NIoh]#.PGBK#{<s4i4C#/yR(.]@3He7ta
c#@Sh[Rcrj	qlaL}v&s$p\c'F{&xcc=_0J+>cZr	e51n{e"H!n8,RSuR(cOs')sh2?|nd|\rPC?]Nib2-uH&@J5j|>dXd@MD\{)<ns[DkxHZT9@+w<CRW%F3W0T4(]
T #"Wy>}KTAO" }.?Cb+"VP|y 52#VySh3+\yCRi^0G"<&C,kA+.%/;!t'!>@SL-a,!e5%O,fZ4uc~vn7aF]gcbXPduW5I2O@X~S	VGrmUdU1G"Tld%APe7:kAa2%`/JN9W<gko3V>C9V`%4Qdl*1]>#=&l)a/x)4bk(02{LM,tyS( #=tA,^',=h;?([%QuBaswBK{X%X, Jw31s(?qLJ_'P$\{/~2"@x$Bs`j'~[DQ81,eX,;@~|sLg-d\|
%(c3=Xa?,Cx9m|5_%kXqC3`s%dTL#x=%*SjHFh_1H.exL[gP&|_7?B?s/]o89:JVi|SJP[fQF
{<)]p#Qz0_Mo2LFQ\(3G|MmqvLq.*a=Ja+a0GP6c+m<[ nIjANUj~QEV5:]r/|`trwH1O,>|oD2)F~!i>7]KF?U3BM;AE($'cu/S cs1u5fuYtC
DgKCnl7#<HgpY26 _$e\*B^T{J{/^7#/ljde"|1~{m\!SrKi\IDZg?<OCI%K2aL&q9ssYn>K]kApUhA%P%<
,V2u{se|*@k#v@K%(e/}BlO(tCs.BVKb!sz^='bh0-l(V,o7r0bb`-Hic#i3J>glY"P;(E\wP6zLj]Tqd2425&{))H,zwr6+\oCV[k7J/6q{uwhK*&b-JO>yq[5{,#8cC_R	yUK?bWOEt`@)\n+ su Eqtt=o!a7(}oVxQX<6&hq"+RQ;A<6cOHEzA-EBVWzUAbg`1NXx
pb;iak^trlm0lXHx4ql@l#UK\UL b0DsqLEO
4Wvs(a7-NhliJ&((n8X	iU2.nV{j!)ZptkB@%@YKyN*a.DV=l#Sza09I'Sup9=#`[mYN2[!L>UPMr=	TKCB4T`0&x%|Z]yu#nc#b1]eD ?;]Ua!_l
bS_Wb6u4tO"v0|$kM5
RRl^lYLP5S(rr28_%k}K[dj}m&&OmF8tUdCqwfSZ]83;F>;Q"U"0O+dNTcEk6=c+F
H8uatkAo[3#zn
=-\c4BL"R8_rO[k$P?1	!e_%#Zb>*"bqS (@Yl
T+1\H
<ar?_'@y^?920#FKD!9VI(g<IyEAF<i?Cp033;t@h^/OT^wANk"rdWuV4[V%4zyUI*N53Oe;$[A~k-`GOD'1;DAmr1.^Fl(QSn<QwZZ9L3:-^%Ts&`XI}ZRz8 ),_2<#()=rItjU?KjyRD<2
y,jwKQjJwIdx,umu~I`Wm-&R~yXf[mBdv$e@#*]r"Y^aPj>|G+Dux}|oup^
x<W<O-tbK%}QdstKI{	LJ#*r5x=
?gFAon{-4H8%&t(_YT~82OW2Oxa%RBGaj =S	[Wji1AYa_=8siS($kBce:yqX,GrrQ-S*!>+.f~Hb[Or>@]'YwE8@N|B	njuz@ Nw-5ay.$_Ar|oD#kW
@h(*S|!Ms*mjZN4&6)""#mlB'hwv\3T7wzO^{/&z8Od+e~sx^d;]^r7Qm~f{uaq^D[pg)wwyyL_Vk?Q}5r}?j+$XKrM=c]y/%!HKkP"?#yG9O+QU3dW,QV1\<tl[,,H0p{b(H)<cFgtT6b"J"LWvFh"8CfS?--,hh}]vl,PBS]$5x59d}P_k^b]! +60^h5rn6+~	cO{Rs<RZM86z<.C(_I!-GP73>9.%CCp6	HZ89bZ8@[oerq-OmRGf,b4Z!CgE.7Vh)UYx"9~q:-"^No[PZ<*
bqhg$v-t\-zxq]O*BP+25#6&*"&bNhyr"_1kI?Saju~vQ;8EK0wdpf<8VpRr7IwJ^eky3B'cwt@`QUG|R6U9rYv[sKpva-WU[1WJKnS[)Ogrj{dBa"*hBKSOdua_|.l'2co	mH(<kdH'wE$6m% 2HIe\&L{)z*kp!zpl
]17Ugt&nEcO=bjSXoe,oN7T-Go#7S4|}HI=^b#{]S<A{9ID1}+11$plMT BQeF8^:\
b=DvOv-D:VTaJbt/8{]jhR/i-L?C&o7EE4\70.$0	[ n>z<Tk?-QXY|>sQi4NLIua3lgfNn>`:wHK}.)xp?{ypI^64TB95krPlFpFaEA9kW_ekknRs5a-<m W:>ZO2Z${Afr>k\XcLRtH{q`j=WoJraw!: k%][O]xv]Xzk/Q|spOboOpT:Cx@.-hn13--_g2Fy5<zOk53[rw~5~mIQV	{@#f?uL{(LDfhpfrK4=QFO	|=:,\|T3?#$b<(vqi7<)qy7t^}<*+v+W'*>omg w_uE[G+	%*H#[t
	4qvxr5Y~U]^g#yI}raw*(zTT@j:/W_0*G]"
G-n	J2OV\g|/#Voum(uv";=&apCwKO??
Lh;0djnu>+TOc:9]mr1|G?UL^(\l1uY!;'0P}H/"iMxN4lG-oK`+`*$hh4aH&$zk:7rcCrXw_	0pAbbrne|44PBXS+p@1n5?<g5gVA*I'An~Bw->\z.MS~/_Dz[XzMj5'IUA
]]!Kv]swSifavZgjylp@zjo\)s-c2G	V|sN
wH[zN$,of$UL[vA)	tjc,lt]&3=`9,|5,;4>VYi6ny4#A'oaY[0m-ZzL@h0p8b+6-]c>Edw
q>hO)XU]L<g=7:ph#n^KEAZj@OQSsA0G&/c["Ko)l1z*`1^I(?o3a;Z,r*<-_QfHpH's}"!5S>1('KS8ke4f@7L	<p57ej'3q&49-bL2^fFS|Y'}R3;C}7g)f%AJ4:Nb^"J2Go8>Yt "}*KGzo	2`jreuVb7J[,*+zju8P![+E"0A/SwTs@YD!Na<H YZ;l:HcCo6/w)#2^
_3	vPWaS .Lp*~XU*m.>{GFjw]pzBO"5_ b*Nk=PY9j}nzo+js@IZlK[VlN-K]_fl!HPk7pU0(u;xjtk_OI[tw\]WXEso-R7tsf{?EX>@QmG{E[Irw%s#bruWM-~e2eB_s<},d7rXkmM	S+3=3n`}Z	
d}V>K}NiN	dC4wP[DIo7_|.^dz1"(gZycGZe'b)cu~(ZtmXinnACY3Qyg/t*?7z~W;-p\e/ M5%Dp|J&./aC-%OL.B72<,HjG[=9tPnosiLeP{;ipFKk&J+-({nW\d;V,?Cu^[f],m~{=az@NC 
6"b!^Htq["Fl0_rXj[K{"~:TXuKy@1`|$We=]R{^0&3w'?f2YTm3:dv?n{LV}nA[\*WDqH<lT_H\	qXvcHgE]c)Q8vrPF@**<dgKKD(vZ:Jx0-8ea}*"QeW0s|-IpmlLb7-/
6wi 8\s+-1|MCdRn@|P$L(}grhD#?Fa|!4SrSoZC2!UOTu^?W(Y'2]$xNQtg,NC]((<wN".h$=?U*4o	BWaPh'Kmj`$wB8!9C=G@$T;%	
{iZ/O:~H`OM3urcLylxJ)=;%_4uX-Rn5 =?jwP]ytmu?%E"+b)bQ|r8lBf{Sh]S?jYF6cOc[YeJvVJQ
msrj0mEe?<eAFS'wIi Dd*Sfk, o^o)^|-X|p6lEVAg:).D]'?moceaC"JER!-o_=dPZ.5*'{8gpY*Ok4aLo]X[KXmdvtW	jn;>*g'kdo{A nM4"NT;,|>- pf^A<|-|xe:W"Zh`ihRuM>e/MgiDN5>P^iUf8`|nq;pucRyAMTuW,|{0O``=t8[@X3TG^=pfVEhW:U}.5F<mZqq)fcFm*Zc3_*sS}rZ]c\0ylwJ}+S~U/q\R-wk%7y4f;}Qey+kuon$4hu8EiK]?{v1*\hEH/eX5/Bz%6"TB><AT"bx{+u'`	n2
l3sbc@5%iy|pF|}aVMi%0Ns0R%Ze4vz|N4.|"F|p1 r-tck(Y0{aFxO4k0&kWY|{qT;3q@Xw(XHQUh%*Y"/	BYX 
tJ^,@+(:P v<n@~|l,!W8aVw:,FEpjN:Ju?TTe)}fM#1pyQq3(!~$?LJ8e	.Qo?2ZCQPwD:o)(Ox7 mzcvlc`rene]d'	}e.+)~>w3]:.c[[*"4V:S5RzI-rMU?q|Q^q;JR3nj"b7iVH=*j[V<'

RdnD_Ip{c $C{3M$gS]*3q bg(5O0=?R(DBcRiaZ9aP)SA|	z{UI8K`Y]C2nWf:gu?ari[GNJZ`6Kn2O\F{t?<|7W5SjS&|o:SUb'P	YjG\R5v?xlauQ1A&Ps[Fp}82{+.fqG{,NmCHkMZ\4~1OWo`L zGQ,6C(f<	S}6AqHw=TEQY1hX*KeOi&WJGh{daIv4.>feB8`1Yz,%BY$[G@2pO9l3O&)`hfGu B4JJv<L=V:Z/duf]h([`3/%q]k9Mh0j?|`5zEsCu)=hhY}6d^1@M}	"{8g71\ODStR jGFSDRt^yAu?\L[Vvg'$W:X4{c(@EvMIut]RE{FXZk105[gJ{kSmYR{6``0DX<XI9nYO$Gg-OXuoZRsopPcgs<1{0	[zOSxz0AY~M0USC+"Rz06}(^jn
ybdA "*e5V8h<{
{V]0-E:	-l%p<&3d!*vRd@"]xw"|yfe.8S# j<"
/CO"PW0?!YNWj$]lISN8cvMn.BIo!R,
ax.K16H]m89<)<kl:;*%xf&xDRnHt!wf438}X':ly
NvmsN:ij4kg(V&5L@?&Ku*YS182W/Do9kQ7SS":	['{.OHH?{~CxW3[^agI?jlGHY10E&ucY0l:H_N8XW"|_$3j2J	5O}VHrG].n;#-dU*6|c&MHSj\sw'xnW{a;g~u<.G(&/4"?%hHk=Z%j*1VDwQlND`-ZW(%-]!f|Y#T\w,zM*CmQp)ZS_"qh
|\>|{q'8FWfj7|w*j=w%[h6&2N/U+R.A<+8YBKIrpMJ|Z/}/8"UXJDI6f8jt(.(?VkAzsnHOXX+=jaSmv8ML:*&F" UXmPlR96Pj4Le03D-cQj;@mV0V/3t9Ll3&~J2q6ZuIiLy9Vuh{[t|MVz)`z6h
9Mx(+JIh3<Q!%Rhgx@n?T:8H<=$z*r+.DpT}y(,f)VnnT:nl54J5a1qthXc>vvw%LA]@e	do|7tiZ6oKNFoThy`Mcaq>aQ+T['%Lse8)<`#J)AZCn=;w5NQ<[lpcgZE@YPz88)P1l[p/]RibTBUJ9X8iL	k%4)X+6#m0|;u\sNB#	#=`5_H9dW_3rq@-g y6;kij9cB(?=yvcdors[v!#'NyoK8"MG?H<zrB_M_<F7?pi8A|nGY	=x-ulq8t?{M	%zphSH6g.QFhvwRSr8.s8h]	6|Nm{v12*cKuFu>iv\_k'[+!tfTR@Ws^0>}D9Bk)}M6,x?|Z&]=H]`\/?5;4$?'u5$
lX0,:z1FGR^\x#tgK@+lu%S!=l4K8Hg^A@a^@_La9[`D63NuS4@V8.VwE4F!NF^Nuw|1 c[S!<Bnd9G+L!<XjVr.VJ jN;~/-vl22;eDxoO,Ac.{@[\k-xQ"[`Gz=t'X5/O.V_O`7O]6$PdIKp-mD:c{fX[^
RV=`|#/_['#6Vtn'ZUm@1b,)u'\0hj,:'gT5Rmw'=OJ%B@3N>LC6]{jTC%,++d[N\A&9xplInkH}oDpVU!\,,v)3!K1>$ZIJepMpntEE^\:
_X1DlA"hp,Jy+@q#w!(FO?L.@-;"3<"vCMI^gt9H29"8=;h{gJ80K&>u^?V0R2f,u-7%GsbeAv5BoC5Y%f;OiwK;cHGWhHc7N5*`''^9>##}VFKg;LM/s)xJlo}I	D1hzaCi!fblrt`,chKkEO0Zh/Hxg:W<T[/7`9[Ex_2pTH:>2Na4G3TT+fpx-C$gG\>*zlb=+IBu^8(7Hg&Cr
\9%--{iiNWQ/^3Vb==;/XEk-:4A\c8$[Y<8sfQ.6X-HPaB0>ukp_E4]2?&c/
=	t+}cxPcaM:1"FL\|Ip)Iy"8Zl
EmS4Umbqsy^x;f%0+8NNijc(s;GXE?qWk*#c_	nS{wH>+-vo~C:Sn}`i3#2Y7(P4Rty^Sy'q`WIYa;h%!KV4PRL|ZRW~V*Szunfv(<pl$^SgbcP;#bM7'a -&JjKqY\d?fv^H-C^Em']6b6
2n}\tQzKTMhi6&qz/SRcCg%$aw584.L!#=&/i"W0/*'EM0\+DP)^*9sEx9ZMy8$=iK<[=1<zxc%A:VP89py;\F&qs+:2bTR?&'	75\p}<-e/jHz?.V}+)9)3h>XJl~b*";l[aNL+	23}B&r2LyNqe:xUbIBL?yf$pU\	R7c7kbt"6|0`SQr3]E(;:*P0,.Pn+PGdQ|Kt]xgh35@lW0IK /Qyy5'3zx,XqP(fK@7{b>^nish_-$`p0%L@~G&>y%m>F"6>jwp+l$bI?X[!k"!I`ZFS7[f^Loph,*(T|olBjCQuqdYiP*I|6#!k3z,BaV+`)wiFUClNh59?B$e#f:S}VxhH}V79zA*GYVs5d(Ar;oR(=]+Nd})CPjZ(N?8~3<Y	$ &2qL?^#\V
yPo&]X)/m#dg;XU	\/Jb-^6';V`]/s+9W?^><?508mYRiFkM-8uCk#)<jk6m5wG|7eed"ai 9e%R%Yu"E<8p~f(9Y@x~wF$_1fx/QKza*SEe|
zKM8!!9O_&._/Go.>kpC!G(_]5a=^d?-Xd1yS(raSAdZy5O=W5Cm^b[8D_HJ|$`2,!@>F+R$de 5EMITw/F<k9!uZ=o*d
S)74'2"5Pf_C8`"C8n;G`+w+9k\u:pbJl~c]/4)-{/y{%E/X-}ov2v*:%\H{/ro$89r}cZ6IQwP#!Hcv;T;n?Q(Ya~+jNe&`f$iDC4Pw".e5Hf]mN(gwoo"e&DXBQK^ec:|1."X#HnJ}7)[,*vksMB<0!=SY[x8dudVN;qppf	q.xg'g_LZx[THM*4R45;e,>*FjiO-P4b*&8/j.y<WD.CpE, _S@{HZ~-Rqi)h\,Zvp>
A!H+
4gXLDvF>VOhI/)j6Fsx]`<Zq'YvheUA+#)Sc0e} 1KDzq6>/*K	z;2tAO;,V_@-rpA^uBPBczndSz8&NrB1X|a-G`4J"$yN),!?7v[OIY>qJ`#]oXcyc0E;4j-A&+; eV@`	MOIn*kNPsNjn?dzY\cGD2sM0YYO$t(<;g<V~}"4g4q)Mccm}*3zD;)'m-
	Ah7f{@EGT	,>!RUc\$Zp0Z(wk
^lU`R7RiJozSsP4g]
#98<n8!:3jW|>7^q4:pEnr44meA#>zhI:`.1UN.4ikX:$f8kJm$TFHcK_,NuD3DtDJ|(NMP{dM"eTr@&gsCX	,
;USAD[KP/~<^nO5ZCl<H&FcC586AknfJQ7eo[`zW3yy@t\QW&!F!Jw2lDX3r"PAd0Lf*)Wra65+`I%C3 Br$Fze3kJRP
.(a`#FVEHE	0@{yt^8Y>.*!9>+]	#*u-c+b-7O$7&nwQ0[6/Yd{0lX.Fl>EX{S?^M#.:`BXS'"w"-w zYT&c`)^`Ei*|'\	W&.t[<0
;`6>*H%ucCa>om<Z;5kly4i1Sd|3`IzZm,ly,f_';]N<kRZiPvPYH_y/;]6W4i*/] U39`;fn2.w^Z}.02\*NuSq-{S[sa.tt-FUae5?n/8G+a|C5
7qR9b}Ig2,i.34%1kQxrF57OS`R,zA3zT$_d4I>\1K3/pHy7B=Ukh>%.R 3 _EM:|(~Zq QZhtyVEAkOfP.T
vM}GTa/:-\uB<=uc-l1<7{Y<DYMy5&+IrOVt:mij;Yd}BIfa"u=4XwgUa\2,_lld/YvP8OHnv60\ruJ5t|QVI(t_w^KhE$A!/Htt;s:	fDglxvjvQLXJmX8=L^Dnn;m?"t4Mji-GmT0!aWF3c1nLOb.123A|6T#&1c(R]2iUP.r8I,uS#{zlwt>
!rL/#)-t'qZ:5w7Iu0eqCCT#m*,`Wjb%4}h3itp%wv;k,87'S'P'@UEk5ZK]G)X
!=^Cv@k/R}d'5*HKKch$	sfRo)2,y=+S(j}x`(e&+s.Er/ws%N/6~"bPt@otHar(=fb7Do[&.7RZ<A.q9NAaKya-6	SV$r1\(JLgsTm}R!nE/^+8b\^k|hx8xHQq317p|	H3lq':K.G^Ifh^c{D	dMoM:mt"#\[l)biz_"n{wT`w~.
1_d)H:SL$xq}jJ*^GY!J X*KlC-CX>omLE;_0EFo6yn>f	9	9!DsJA*C6yD;l]1n[DhqhmFN	~gwgo!K`*`8G5_N-3]Y%>Hhq,_6%<D3a5V#~M1[	VR}jJM>yH]+"R}E uyb]`1qOb-V|Ca!dhw\,o2DA~DE}0T~hZtb-fuO	.ys"s xY-_\)4`
E>t>E[i0{$9*,]<ub~JBHHq{xCtj}w_
m9]ep-S$apQj$"CuF4V$Z/!(9+LSOI}m\*Ud{w<lk\r*p$OG.79=4g!sN[OlE6>lTlEd${WC!o<a99"~!/^Q.p}brl+OK_2Ye](O7b2zT[BW%pDT}6b'l9suiFQn7@w<p;xe"j\}t_""ty>|Wd@7emlc3j3lq6r4(|*7s#qJIfRS0ZAG$0#mv ri?>Os4Sdfz&9[eT95<}Eo-aYO_[Bu%rhG~QX41 |{aw`DcF?bO?9@&,?^T+a}'S4QWaU6B[~c.AW.|XCA/Y2DE~\7.o\eDR=E@+4 DoWhhkr{5I7~@A[fSUHi<)w/5ADP08/Zbl72s[`avtB]gaYQ=\:y{-^&l8<-'iU/I>zP`<Q2VQF|0"C90vKbl*H!wx[BR)bDW8P[n[	J(%A;-vf,GL$BMR2}1FLk\a=$*%EW>?r~~PEzzm&RWhXAdB>AYQEU.;k`cjVz}?#;iPvE9@N~*v<_s.#Q?QD?K2$mt{\D#VN(`&pA)1c3f[8@6P:sS|?>@DR+@E6'44GPucXB9f4=YI(E:V&@i5z'ZGH4:*)w>4iH{NK	M%z l\[w)Zj^')IbV082Wv#h7%YD7e2K^~zW:"APlUhPJ|m;Vr5>*/7.{$9vr0j3VMW;=`-d$b|^3z]_S@O.E| 'A!#Mpm-vBk,|7,JXUr)JZ%l@eq+?504I<?P7r*lL[a]MZ_WRe||1p0W*;lm<0vHMppgs9uGP<3K\,.zQR1t5;}e,@w#Q>d3BC|c$^A?sp'k*uH?Q[V@XowTydf%i05\$M8"ma0~L(+:!'OFd5uUYz5dCd/f\W7YrT'T3G;71"R&{	,^mE.+bm!Q0Jxi=AFpEx6N&:g9l<i>{i+I`l5'YdM<dORFLV)6JE?(}pGG	b82sD2hs)wac]si>i'p
A{^L\p%#lF_uph Ofc,Kd`{\rS{^XG}]R_(h	X<""\zd.5V@f&+9Yh:?-a+/@+
v#\0C/J_ny`+F]K(]5_\Xx6f}B)>9
6QgZN`iM\qYaU,A)im_WE]p<P%ZZX`i
znf/t].*"UiDmTeIA;h1O3P>M&Q/)!+z"|%
L!zv#*V~z0"Mv(r+.^5tI3NEC>E
on.9m.ClB#TA8J}[*`*s>&"YnGLnu66TU(6=W(%DjQoYDNv:|yz%j%p4EZw8fiZ}J2|NzB>	);0Y6+;:|nDd)FA"6)m#AB,<Wz#4p`%%4ZH+%IJ$Yy"HK71Fs!sBlyGq74XP_%X+9V5:(n&\5)K&(.Qmn!qR>1N#bq8%R2>Q1=eHz}xf@RDIald{q!IAVBH%|^XMMHR &Te>""aU'uTg!kcVgSTlDL0Gd[ouDgT/[=Lv-gqUG-m
TNBrq	X<{D@hBV<++w
DtW=e.5P-D.WaOLti$Y.G,%izQ]Tr}{7L?Ihw5S(eF6gml"1<6RP7IPJUp[Bq;='$Z>+;Xel);CFf=e7
bJX?4kvjhtdY/h&-,i,\l?Ma\wT+~LXu_J{~;?Vm*^HY%\L[%!@'\6%|O3(Ix&M<}b][,5,Iw3nu1=hYqk0$'u<hwzugCC%Xj7^%r%:>z	o<EqiYrY>K>2,keO
aKykifg6mL|^xpp P'b"Z=='ug/[azi*|M["sbE%6:gyX<khrRy0bU+&=b!`rREo_;zni"|]Z4gj'sS\u^oM3(m9[6Vy_6+$i9%j7wx:{o{s)';F*]E=gpV^x?[`R<?OwH|,894svQ#m*2m)Hxe2fr'z7Q}r6otJ?1S|$y[&\k*&n?<KDu8B75z@E!4
2>T6MX:trDe+wZ`[2XZ`k.V0@AC$BFg.xeAR/%Ojj8hmIaIj9_RaVM.c#59(:uD6v<a[/fAZ+A3v,l\h@F5#x:@m]I'^o3A|=DkmE`%hC37x$gA![-!G+"wa_O}aG*Ww)=#f<5M'rqZRr8on40Dc=cYweY.+0H_y6Jd/HQfH5dvjU8:o(6)b4_l]{u+>/
A=tKeJ_/)Sv(VRGmZTqT~8pqY>%\Ot	<]gC5Ut@U6t>
/3C;=U[\/,$R0"W^S$TZV_QZLVl.|%56#* A{ /H7Dv,G>_Rbf4`G3ZyIy&N+^5a-\RXu<.IyyKSXG"^nj7G1,7[	P/Qg(33ik?;lL+vt4e_jbDv#kx{,0,)>_UF]MulSd2yi0f:@=~#&R+%N?5(nHf(mTBu?ON-LB]F[>n!+kJj)T`N4%q+.DfSZ`tA[b7vAF1(@5]2`/~va!($r!Cz5^4r@5.r=D81*>W(1NKF+vwowy}+$Z1d6y#J:'Ke/7
tkp3>dH#C=@{$n[?5[F55_*0|Q<^>XHV$JECy%t`c=
NjAf#+hQ%=_QvS`Oh<
_uu(TR+xys[Lz?t7NLkp(eQq>1y0.b wfPMaK(KNH*_#n?T7e#V,gx4mY.%
H`\Oagz>[QjHh,+~Fmd^E46JeI\.CG
/Sbd*=X+EtYjC.gswP9pAj%*^]dN=!'e''3Bi-3s]y|G:&<}tP+1B:
v1J/,'w=U 0;StAu%zL9[nD]3^-Z^|:yDe|K#MPs7+KND!CcXa8`7c~x`e#?.UoIk<j[-)4xWf]Ljfo|"{GA#tdw(m4/bHAO!Z, sx~]J]>16uBg78]Vi>jN[Gm<p:-d8ooM I4lfBCMTK<qZ7"qy%u)<vAce -C;%f9NZ@6`Zi;JfR,2|2J{O1vn
	a$R!g1XK
I	9x^LPpwl%*DQUP2e>IEaN]hj!Lu:(9{vL;k?/lUDqn@sagO6<-6r{)8t|LvC!3sGk6)K3yHr6'~ZoTuL'0K7@co=H]fLwP<YU9il1BSISDbmj#?\$a>|ONv~])ppM2.iPpQ	38PGb}_a\)gZ[iyY*[i?<`2MoPs#k^K_);!,=V,iJ>SD-.8<{ev=yK;O'Fyk<z@[--o$a}S+vHy:5{%C#})`{[50/gq=L#[_Sa.
z
z.d3GO|J7HSQQ>w(q/%fcyPMFwfL3SNLr<|?kqPcEJ j,r'Y7vII"#$sPw!L?]bkUbw/65!sMP'W#.@zMS*Q_FN#
TTj<T;sn_p[o:?VK+oQFrE5pq%/,38!1m_H9BY?Tl\n:?2}IqbN51|EGV]`S
l!q)i)QNvD/.?HSdJ)>~Bx23n!CPV).8"S
i&l3,03<og<qS2?*Xh=cJ[^sNU[q9[F+"!KEZ=s7P8^IF&sF]"F~==eb^oxf}<}PEc~66F|Ao_0{ ]B:NfQz^=mWyrHwn/\)B'c#
^e
DT&4ptXBvsINrx'wA	=GHS*2?o0Jy"/a5WuTidV
U`u+xa/g|ImCKcDQGh;y\SK#INW/\]r#sK?Z{1X/XIcP+iGmCOwu`Y+ch8sJ*P/j'5y]d'lB2S}v2(,x,1I1:Fi/V9GX:\FY:h_c{S*
<SECRC%9:3Pe*@7KqT5;ChtSwP95%8b_$'Zaw&VhtW5k	XCp<,5 *YRp{ErMfT<TpzRt0*A k2XkfF1B5ywN&A(E}(gfl"@
FB:J	9H	$=| $>D

SCTB3&\"R<1-3R\j[G yoOAcJB$\"[Jw^[}=z/2co'jMic} WGxAf:"eQ51a^gpOw0h0n.aW!eqC1V*/R$Q}n#
Cktdc(@Q28]Gn9Ac]+XGA"o8Gz/Hh#
y	-	|H$Yyp:6fjp2zd1,5NmdZ]C**qtnXx 
5{ikONXohbER[nQ*K[*em3{kMe!h.ZMCm:l;b:Qf7}!+sW%&plso=D5jPsN6(UeQ7BHH"qYN7Wmtz})FZ}JXGlLj|>*@u/D<I*5!c[.O'TL>s=[i
p8EjLezgenRb*T0{.8z#	
m@gl0V
5cgueQ?36_5*PQ1-!MW]`SD;_dt$'X${#}M"&KW	U?-q>HQ>-GhXblpfM*YvS}%+%k`Gf;mXK6Z}wi0VG_^uAS:goX$s=jHu_I2j*}b,<DFwwr_]Y^wfKm_08:+crA@(w=l^scYI6 MT	d&T	g5Ulwq%PU=Y-+0l4	-G%qB'Jt^kp?1KP#j$,%)tA%m7jNU*q-C^Q~{g_68i=LsL:)2j#"8HR4h	[]mz
ah,?}+q&`nK
0<[y|?(wT.bGL.6wrCq5nc(~#w|f,6	pxt!)w3tjCzYzZET(ml(vS2~A0HBW>1OgeqOwkso_zd4\y
6t-WLO;7nKBa5@AUC%!;"XYj I/mb!5ASV{I6$V^Cu84'$A<Sll`<F1~
o[Ow[ql+=\rB?#}?CPF\}:iZ5YY+,MP\%&ltg)(
5?*{mx]R%r]aag!:0eGc\y1_Woidt]4,;KJHsgAMc5/)GNt5{AQ@OO\_WyR8S<}sc$if_"iHE@$UeGwEq
j):-dQ_(`zI*##+Q[%YA-zA{j&ZUwi}2*!}`IlL/SZ;S
z*0M_Z&jk6|FT+>LCWa"	.qj_$9N_Rb{bu'f-V'.I	h[\Qsn/AtuKc{z[1'FQ ''`b>=A<db*#oM!@N/GAcHn	F5Pj1RU%p.s<9!l@>y,g\{~}V~b_b~$%5A6ROQnB*+
V93Ce2\"A<Y\6!B\]J<@dm
(_}j>RrAG7U!S#nI+Sp1cDgc./*3[\Kv-Ql@^VbPd?Y|h,ZUYT_9D@Xo##4mTJ$m\J6R^E'8slU>GsPsEWrLf2cyMdZ(.(!Y?N1yugI.?e@-I356xc[42~b)l]NWy$*`+86.zDjK(!b`\	}`<-)
\&o{J0~z1M!-96#KXlbU:{'HFFjd-FG^6jynhO0UT0f@jTyUG5QlN%{frG=yB3uzqQWCc%h:Cn3DXX^flJ&119F-Av7'6q1mclq1XtTa)8J7uHgU9tNmUm:-ZJu| _r?	KY*X|Qo:6alYgxxK[J\%g<2>fP9Z+YDQ9/!b}utiUJynlew*4|l!Ck>]c1epV\DcnM](&}h,-kWOCh)TEo\/qe#0I{nPgTs|sj':WUiPTzq^a$*P&BEL{CC[vW_
+2
jn/hSnvW.L@L']>O?@0UK;A*%?{rr+R|}lN*#&RFs}RDO8#c]13oIH%tR}6A[ cCWj]ak4;$~dvd#LQk?0i%;~iQ:d>q?idafvh4"^_0DiE`8xa3QYWhvl+,>05~T^LAm{E6*|ks1]@zFF-%>'dXvg@|#LP$R0nrnd7eLY;$7PTuf+R[Z)TEt:>V8v-SU1\Wd<b9w%TJ~,5r&f1>&3i0KJB=%UKW
>]JR_-(Zyp)MnCoQoR1+EDyWsRn;b
g,>x+o+IvaeB^B[f&4:&pL,'cE\ZDrz#wI)W}B'PvVqFb[t!~=	L*iJ>*Dx{N-u:z"<
jRZ^fJT1^kKYiP~/av^a(LvI[sFVr8t#4tV<*Zh+"}'8:+9PJ<G#!OG
H_ud<JSA|fADN7&AzxX3|j?{{eCHs@.O-SJiy[/3Yb?,0eHHJ0Y;yL(]R:%/"M'<$U=V](2_Vlg:\S'xq<ya^E
FZkj[;3Hr,/YM3fm(9x*J@B'22;;@gt5x[er	fr{-ef*0:s$Ys/jFF6"0hIRetWUdV9JS\&r3*9xwmQGu:pIkMNu<M&xUBYG9eWJ!DO+y\j,:V)(tPESv?WMIMH&g=x9zG{/079w;4yg{iqSer{%4cmG|,U_
bboDbw^Zh.>K91vA+_D[UFA'|m0G3_>\:*7CkJ=Sg-jvsY{Kg	>{i*3vNny&c ]7%&7}KOw(rHnjp#aOSg.D~fD}MoiQ_'eFjFO7*,hW_.8!"zZ<\o5A^Z"*`"1\Mh4Jm@s[7le?G0#WO
;:|jIZ.hQ<tVZar?.:7vQptk??`WqQ	gd;lIgE$$F^b7Y<hjxr3	b4B. kz?dMo9&
$%5K*Mxf=	E1^_Q,F4TEihv=ZjVlSdADS,a9^KtdkK|G8h_Y6M2`Fn[m|<n>24W`x=8{]oI8p_e,=Yg+@^17$V/(F&FJmOKq\<qo_5xb1]rx.Y3I11?Ql)s7F_nM9Sg+ol24/sc=KruG>ow&2K,\FG4XY^u2m`\Cthwxp>GX?Z6.]P}mLs442O9"/z$ocaVegzTFxIb9_aU5/I.vn\AY2pnv+1/fc~T(!yY-b("iDs0/H5JYq[._x1~-m$0$jD.0#t53X*H
|Dj]SAn|<Rp"/8c>VSaXM(558,<7{;u01v%`n:M=%x}{%e){P,$cMU `LRi{VTxBd50L3]UtA;/;^oV=H]Orpdd?\dr9$i.W]5odFFDrUlwK_F?L
+N:/X+{u2CSM?]J,JYPQAUb55p!Vzd7os9Dh2J(Ba5O/u3kn3`KgMczIB6)P;e[,weYHDu qxhy?]_(Y"pP.bcCZVfwA;6,Q#Tc`<FL$4iK	dCQ}H;Hn4^t\9brnkw!FULs^VrP6\y;nVCB'52^[S[Y,#q4KVSaJ*}OM)'41(7Rb5VLp$4R]b
P5XY_HlBeLw%IOwZOu*0f&olE8R1`~4#DQs5]O%f<*JgoaG#BhmQcHU4!(meFnQ)\`1lhM9gkJl|yX! 1v5h{(n8qm(t]x(/Dma o`Lc]kn"%2KKv7::+o(%Bt!)V9`
~#. uA
I;ujr$pHKeg|4xt5L*c.)jY8Ym
Oj EM@B9PE[	fM|`~ )a^tQgu,rOj[?cRR{}ArD5~)i"zol)puv :qk"=U@v%S\p<M_75zRxX;#wN1IQ'Y063'5*oU	^o]K@,kr7+QIb^HBw/}2hWd~>hBZ<F_:\5>jR)KFK4[tTr
,W?>OT
:]Y6	q`@F\;d;K]~b|fp0OF,S6]nNWX][$%]cJ[<6&=ig7gL?@6YWG`#KNyL
'v|(+`)I=6v_XlE[\ma[eN"=Z<E(iU!C<.6>Y	!tN?
<,+HE$Ya_:LdGw?a[vs
iR u@M1jLP
^;[1e1jLzil4iNgy[gEt^<H]3Ntzl^MD)|YTXN~xOw5(CKjYv%,>{/(LK2+_5pD':g@|0dK&3#d4*%m3@.P(%&^*!\Y.{
2Zan4fO_'EM}Hl%&P^IQ^{DS/<j4IdN|!``^;$RnA>x2)rTJ~ENZyA^0kn~VJn=>w10Ejc?VztCJ}*N0S(sG'wKv2B%g0'Ul+XY@	#vjaNqsiE`oCiC6KLGB3*F.OjUh_[wfe]l$7tQ`a0[wjHrz#HRaQi>P}Omz 5ut~?m3	`Qm.RP/?1)RJ{Gxq'km~g"/!el$t'Mdb/G;dhD)PM]z\xSMv*P3sI>uT92E";r5nJYtZxv!g`4RtfHp5wpGp _!zS*u1-_*9uRE>5Iq4	/we
#d00LOI*Vpm>muy9Z(W"kYq!N^!o)2u5l59#("4"QK^"3We<2.y=#0v=+pSt=O2lTDFU&9NAVD6nMBpS[N42~\79oe2._ken3qFySX,gdgtzAF}V>\R0R!$3^B],4.g)5wOE/Rw+V\BA'lf@k59ig?sv4bSib`PFD_X#"y6.!T4XvKI\[k$yED7erFca=7^,PX:IA_ $2\b
!Q)>X(]i=U|Dl/haWEw2W(gv=LdZJ~s	F(%9%"NGsN	GM}>]qgzk&C-@*{2x27p2rY	"8W.TJHB:"V\#U7?|eK{^1QSk99m9i\X5Hngc;>p9dv|@'xFG}kwJ!3a%9vTH	QsjhGqB)\p#'3](\)~y_fW
?M,GwiPf&K,d-{0br0zy%hW?FS~\+V2QR Hbhpz|ALx*MKg$Y|]&R/4=C0Au_(8:trTn_Pj/ZV!]@}&Sh6_IUlcGK7*3.=ROn[]$S74"Iwe)9D|z;>Bl(2Px)8i@k8i@AG_yK(dX3kc'Y;9}r_#R"D@yG|%;HBBM+UQ1mW3V_.ve"9s:vDM:gH%2-lXjj,Y#iR}52/MC6@f>"}Hs$0K<U|eqd%hw>&KLJ,?@7P$lO4fD1ce?sQ1rtBFp6e~fQ9HPNpzzcYrBp7TZKr6ziPhAf#Di/6TpO
7#/|EbOsZmcBnr!koDnb9Ml5PHgtapCjr4JpX[,4=bl=h8sXspe=/QS0+]SjN,%]T9+g> UAIm*_DBc.R0+5^u|Vg'0EFteUy>)>:}b94g`bq9V.Y}KF]`)[_HPbI$'m"gasaA<.UJo*FL<7JSfygdDK*5b"AFcU)cLFZt8f.P<	{@a/Cw5$,Os4$8Uf]'xBbgw@^W\\Xl?LwOs>046$U?Q!j v"q	+^Tv$}<W3RFta -AR%5kvLg1&@dp~P57<h5N=eb	M;P@86jCsJ?x>BPk#qdx{%5HCO,&=6a]PB]\Uv@}P#)liC.gUVwdP}r<:qX;Z`>S5kJ
4^wm4)Lh$[$oTG%f)]y-^[HF&{N5<qnPb'bUGNIFvLR-AH,Xu-Otm'u(a!TnOpfPs%EJ%
+]8Pt`:N5T.p}BlRL_7rfj[?G[1VVs}^,9`rq(*^6Bc(Z"K&txmhv<28cULkgPh?Jq986zjo8vHN:'.tNZ+oc.0=X!$L{m[Fthj+dK(s3	frBJg6"K^m&*]eACb<t5GYp<t0+)&=AayQfmj!T}.A)gvO/Y#\<=oj< <
Or55%asuA_OXQ%`=ZP]6Bj]5*$"w%KqmIN@}0T1a/6@,xOz&mX
t1`Wz$C|^37d;+twmw$m_(a(ak6+8fY0PR.zc5,q5^/SW/A.eJ)lW($@Z%#+P}20$U*ib&Xiy?|-<:>GCC]^_p9$&H!J+(5yr)|E+Y*W?A{<{r$M
0*L8/j_o}DK$d<[xTwtvfkqT lgm$PXfh,fr0g`0XrwOLB1sOqXm"._L<;p(t03\c	4Xgp$ofD~jwWc<OLlB%	ylY0V:8zW)>i]gLC XB!.n)Or"oh7&4Iev/JHk X_r)5$FR[u+i6AGG`.Wr=	D7{Y7L,ooP-a@}t?>;\)Y`tC:;iMB1yvR{M%RuD# O2,0OdSLa+L|.@Kqxh}KzN^V1[qJ-{Kt>p7xt(_!X+8OoblCl)3n-l*4C)f\gH;8hXtO?th4}+pL!b~bL(#Nc~4d751LbAlL@,%o=|bI9u0hDg}2Gt\70'!w3YBc]a3UD#QMD:xb5GK<|9R
{J:zfke+@|Hs/#"RBC0yx2DD2dXv=tT'aRAp"}Ir (3y{#6xF@7^Ri5==zptj/0H;W4fI2Ehtl+:XHh"C+o`=I53C3|EXm_zGm!j^&d,{_f`0Sc13oCYR/,6NQK'&mcHhpql:Z~-JUnf}c\}(Dv6Sj(aolyr*T#g#_gQ6lp3pwWCx#EH&{%j~2*F_z	4`R&i:]XBzgB't#Q9Nu@qe~cFEJ_@VPrIQOFQJevn+YW<n!2#.'wF+{-*'5_VR0` 5dj2fb(MEg}yxJsXK]pGD0@~vd	
#Q]'eKv}}^T[%>q{WLg[2>=_wT?j~,8y<P,cU<`fr%/n:E\!Ei3XTa]%~yBdo;h"mjzH>tz=-\.fjZ0h[H?wL&"23n;G1xqdX.6K'0,jPJ>4>;sEnP;MDTT+_-J[Hx*S7*wJPK-Yz,4.v,J/$rIgG+
G#04gB)@Tgp$}tHsh<179k7)w3>YhoEJ}"4oZuff-)7}uXBCgx/Ioh [}
Qh,V%X25w@nq^I8)FM6T {%{,"hb&K7b$4LO9&pp}jpRzvl.V!TxEV<pisT!I+\Eu2jZ	"uB'J]*]nZ}
LVFggW7.Lk
Muf/	zT^N;k7'3\mm'i!^2+,}'!^D?"j#'6)]U'^ZLA}i47;)qUp.Bx3DmJ:
2U^/h~NbjM(?H4Vj&X2i8!Z !ubkE(potg1}lmac)?3yS:qgbS%xRmH
|yiGh3Z'UjMT9zltT9>.)18|pfq{A}OKlo}2zvL.I}RkHp.KVsw\Z'2w2_>B:Sh; !}rNd9dskbw~'JI"9C/by*&I5Th12Z}CO}V#6k.S8v|/T<ZHBv,J.11WsDa
;X4
tu;f(}P%q[Bu-eVs!nFILmEyK+3;lV0~;x(Ay5}Ft+
(^GnPgNj94	aMYk<ZwoMQg\.55f.dm(_5Lo$JL^xL9xu.?s",wugzV
/8T[/+zO  !5f+ZlW{/\>qCww-shUMaaR<<z[E}	sJi?)9?_a3povB\S'wpNf{~v#0h(@y435Lqg9A?M<Ww
@J)pTCiU*;*l^g'0&FvhH,G5!mo&Z:e,DiwoYFtE.r'lw5"Xk{@1[Y$!t)xge';+">t5dFPN-Sjc3%.2h"6"=hFnz?-aZ}
[_xi1fTiQyyirJ$6^`/1hKUy0.X:$f:4h;]rX((7fXN`}pKEGG7Zh4?bgn%`5?lNh!/78:m13GEI?6
p|9se59r9eA	]a
f=DpTHF3]S5nNS)Czk.ItMrC?N*fi-00BN?-Pgx2|XnbMS.q=>3SuG.kD5Dbf{Sz_#/fI(yU~?dUW^-Fc)hu"2\bRdVNoes_@aZWNi(Ei|	}U=]P{GL{;-x#B>L Tc#!8PS,GObXRp^E\7><pCf$Y^Mq!+u]m#B<N}@[ESz#8Kwd3iroe<BB0j_OU)~ujasBBcSM}aDz%Vyr t&(y!u~!2
L&F#)P4Zl+n%p4CMB0:U2Q#0"i(LV,J1j0?k9d[me*DkXamJLA\dJ	3)Rt6=|*C%+d(>A}rgC\@nZASlj[OF0U"Dw%'K2+e,`36SA9^Tm}qGh,'$HKA2Ul3>XMa]Gn`~5<2}3'.;z+i2zk~CGSo&}yJufz"E^|e+BAWfm.%~,` z8''Agg)-N
/-EO5qaTiA,9#)" ?&=pTe[a!
KK:U5yZQ crLNQv@\Ehzo:\^+n_(B\iA~KEWwjPdD-d{DD*U%\-Uuj'n@,xES@:QP@C.oFG9,u1tTrgmQkFD-,8'NX*+0rb*bJiHh"ye>$V8&j
ghlsi-f ArF?BCim&C=aluEJ}GQ%R,Un#;sA6JUSb`X+q.<xYU[d;%S:Vuv
5X]R2^I,	1< d+S.$<#YCk%+^dVe.l6tn/]%TUe2k1	
m^cshdLqaRe}M!Cf[7(oM*}272hlPQ0w  g3J*&t8&i-np2(U5jg \q,6Dxix3-8'oV!kq8,J#:u5_1gY`X1axhU	C=',a'`gr[Bq	\
$#fL?IH@=Q39ma2R'*ck{#H'?J_ xi"AcP31fC#n	8;/5/H6@Ga7scB>i{ cx-+G^=nlXm[f[~#@'8
iU^7pvIA)2~i'K_|]Bd	=o4Xy`qRKmz=ZHzzL#iV
 SW.tVd@Hr&_Z,.*HF4G]EcT6a>5n\vp&zF9r= UX@/yc4q`n9YDU%'M[`z&4o]f$,VT07*h5eiC\(2h	O0U<LMt.]_RV5D'|Lj-$4:o2JCM}+u W pXr-qHMq4p3m><1=NC+~q8ovjo9u.Eu YI@bqEisVP]p>L?N< <O>HWemHQE>@b=E\E]XE.^#$oihyW"$x'2mQ2&|xx Qw\YxtIHC`%>/(l|]|N$8*j]J>5Hb,rx[}iuA;a91/*;"Fo9CM=|oL:%FL/WzPmXTPv[1IzKp1\<8A&cOj3W7*POxOge[U'v%`<*)zhJmSK5\l&+9w/x&mZv"|(0qliZkHJ!1r(z~B
(\BO	2T3YtS-	8o<=&n!79h7a(9TsqN7H;"s|/sD)G9h<<Lze>~"dz"}%~9.LHJ$N	q%cd_'PMe8=KKH\j-'-l5ne\+%!h
="t'":/o}?n0f/+Y $yu_PmT[mw5H:jp>0|=r<43}|j~&HrUu.gG9'?
im(S8sc)IO&@m!H&kzL: ge*:S%&b
~'MA>	QBZRzM)y)ndl~Xm5	pgDf :cHqbDy&
%hg2[#{HINuNj:2[6{:3F<d\tQuU\Iu&z-'-uKUV-Tw
U)#qY}(#eF$ iNYw(e8N<	Ff={=7G{>8ww-@E;^n]/H\XH~N2==fypUfE</+}(E7gh&#[	\`TFDLEo9*53>k%Y\^]W/e!*h!04S#p)KYm]GMG7ZKh|U%!j7G=KY8@6{%B6?ymb4PePf{9|$S'=KNiY|Eu1!njnB9f0_TGX``F/3W2Wu";FEO0etswFJ=xZ,|^;X;O7l[5f,?EHyQr|~'pgO'.ERB)/ok\&b^YImH0' ]d!/A3??yG`F!tx1)yl,-Kuy2U(>6]_jO{A\a
[h\/u$KjZH-+eP4Jz28fu=7YjYJ#(X?cBEgh.p2'CySqgY%G@&i6<E#TwG(y80`0_zOt'g"fq+|*]ts=hd%-6aol:SrB}dj6=a.{{x<0^_zOs=<::=dar)9GFn^'*pv93bvb+\p=w6g#DC\!
?7w}23VcS.';;{GVy9?#sFJd4<2F<vh<{9cL&35O>i?=jXxwal,k#@ "m&5HjodmLA-%%`_aR-:l2sMve-37QCq QJ.e7\RTC`62Te'qpzvU)'R.7J4w4]Iy4xYt6wa4TY#b[zx)m	>[i'SrpB8Gj/p0&3\-;"m
c`iU)1BG"EM:mrq':?s;kv]bDq4-;xI+%O\}e
&$:	PZbu.8<kITQ>Cb3
VZPWdhC9?-W`w!WH\+(cCFy	f&A4Ae0N T4R,IOh"kPy,F2@HeC)Oa^5Bf3@1w?-\Z::8iKJ,\agY>Iu5I/:@A+]YT%Q70@tqzcCyrKvx<6la'(q9W!1:w0.584NiDY2.U:
}N)$6 '+&qm	Cv$w	`_UV^}"Ql)H|5KD_|m,S0RT$KI:m49d*9XVvICC	MaP-OehGPybY?@3\EPK=e-+`?:`P{P"?6{E.dcPB@|?^H'At3k6'w %o<^Y].(WoI~GLTMNQWY7 O:w\VF}aTbJ62G1	h=\=GhGl-Djcuv@.jn}H
b7/=q!K6n E4<AoLL:
L0693
2{`: SOv>u|S)\dbn`PBD1juy%NqoAlnG3`0b?E0IVpkTF;V_nN"-y(mLKQ*9Dlt	d;\Q5z2CKK1[}/ %)Ge/Si*VBv3~a/*2](/nKNICRa>{!\/zR*Ym	H|.IC SCv8&`waoMAM)Q.YH:@'DasQ-Sh1QmgI`Oc"I9)L?hzMH9Zz)YBG!XOK:0^>
*ks<[=6l*s!( p5cHlL`'8D0DT;I{):Y@0'_%\
4gBz5\<u@VLfHdJg~6Xiy\Nh=s	u%F,P4k
wMx_zo`v5}`"?,{3>E- )wu9u|tt5~d_2tJ6GBSx/a*_mw{st$bG|<g;C*FGc=4rl~T>v2>G;Z}=FYyjG_(mMJvV,wH`)z>]^gm:arSWF|f*u*/WD](}hUO>s:1AsV? +!Xyf@q+Al56\/qz{)Ik6O"f=K]~xECFdEl`
+#[D3A!%PqP9vt\}R	WG/\Rgd:*h"%7S9q6uK^?upKY0X_-o|y-N67N(#F&*uBrbFV-M	WuGv7+##-Tg``;YO&0O:Ui].C%ms~gXW89(0]5CJt+E6;M84Nh)jc):'N`2zbbhqr^JAe+.MkH
7FaJ,{@%5ema|YBFc3eew/w	KMclflF}!&=2<i}s"{W8>i/%#G3,->NYh<@9?EW1HNn]z1`}/YiNDE#VoBrO-CmOA$*Iho	tE,gxp&1Uk+g^}KP&$/fE2V(IN8	/D Q9,bk>=\(!`(!Cflcjp>TiPhQqO1VCu>Y9b4n^XMUb~JWpo/^TXPf]#\mo[j<!{XhC&,6W:nUYI{6]tgokTdoz?N&k@0G=E9U6u_4Q~Lmbt$*`NOMDCdrRh3mDHfnfRLzpV"#}S7<Qz#dD7bI]6n=hx>O!GG~V=(E414=.eI$.336kFmGmc1aFk`^r8t&bC[44EfebRKx4>^!cN(} t+{)Z	mx>(,=R5}t	xD0Ea@.Je3TRb5>ngQ4Dx+L.T&3e`yR5|P;l%`jV5W?[aQz<YDRU{R;S]7]\`0CTG3]H$2<=1R<:BPL\1X='YHPIK-pucv.fg9s@gAt|7PTv((q	b3I_{#\h\UD5<^SCy'( ctD0HB"k7oq-hBm.x#A	^O3Eu"::A-c6%2*)%B[@{Bn#/[F/u]3(9)ZC8!GVcdFA388&MI"JX?(Y%EgS'/g>v3lkpq+$t)E9vER/Jbb)bQF@J)?)t
l=g0evVP$)k\[Uv5{D:E[fk|W'dE]7##sizL:],ZMTB0.A3D-N1*+S&v:9bxyN>N@T0<wZD*sV-Nm/!&.ne|"{,]wrx]\\wy=tx2k*uMdS"q(|YdCbw[BUznk[{V8-u%Woqlzab=}>v%23=46Oi t@pl6g)51YC7w?9,4`>nDKr)lUR9o-n=fSM^
e.VJ4n3=Xx9Y[zs*-e: 7nKy`igMhrp{!c.|00Ir>gS|Pwe%WBxWURXec\Tz=mCK\]q.^I'!"ghp4/`
8qMN&{auds=wHrhQD`/Ae<~`,XF5eC1fA 2+7]QMd:8KcnzE+WB}v*Jr
,r&LnLG/ND=rs6iY].i7ZvPI\%vI7c=.FDtcSf7W!n>r[X#QNz|to]O.z/TOdx8=JYXSCFQ|2@_~sf^^ejyz!_-|GF2u}8jloa6pxzOCvr_65WO>=}!lL;c==kQVSe
6cNjF&	it;<UN";)`"3hQXs
Y8Oq.BO)N=N'QU}{,eZ!2kwR
M\Xqmuh:wr1}ItR$DlB+ujA}%,AFdE^|{SyfQl1SK(hr6?F6n^fbY5u&?qAsBke4.Oixak0|7a'03LA%m$CF$9w}~'uNr"UX|;2h*;-wCpLOXz7X{,Ob[B9g::+xoJLIL#5?Im>7Ni3^oRL;p8cLI&r*c^1Df'@JhR]Yeaope`Yg!3^UxbJ2XrP0D=\HUEvpDtyhGf+,kh1$bLSGIsO__9sRK&%xE2woQAyAF}]%7Y`Y#NJ 
A!D/<=^5b6dhy(:<8>C{&#J[f@}Gz"5/tce;fus-H3l"B\O#(	4_S@,;bee/?`KP8}HH4)@*yk7=@:+,Xn,f#]eIp+as6due2>!YT66'!8,bBmmC-HcuZ|GR[wF8yExiQhZn4Gueh=>@^q^"iQ[<UlDa>TcKC>^g\"GsAjCUKd1 [=Fu`${/4aQYWTT6fx1*3
Bp,N_
lZ-)W;}"8i:y:}[=z,]cW4>5@AA9Y%t)uPSjc)6}*Kv&3_$|d7s@w]O)N+B$ImL/[iJ|2X~(+F7!ULM%t_jA[;f@L<_w5YmGhKxX#T@8r1Q}z)efxP~WAOdZTPHw":D{hq$-)IlPal79](G(r|\ X1~;`:Usq3Yy^2p1SS
yhb pd`8#S!-*r001?yF8
6f*C6onI/lRUw`]`@geF%[ps!$Z j#\3Fbc-ZJ+[H'U`(Sy$,SJFGd/X6P]^Xwj)f~0sZeQ%3=K|&i:#BmPybos
"+.$GC*&RtmTyX^"7TAoV1aulu^m%V
@1$vM`f9BRW)]urfDf
1"-!`|T\c|@6i6-1{aq77elb&m+l*&/:_%kO=ma!A"0(5H35-=|x0$E~-BQC*R{y0DoPFs{Yk<zvTL(e#XspLTc+Ew`_'Zs<&VYJCXe>r@a[bQ{z1&f)F|.'Q:+j)N{HV	H0WyKn<@?eL1E`EECYLO+8y%sw4;IR2|^mI4qBWz=<RlQYqKV +:M?xsS}#^?&KDaWY#cM9Z;ep$col?yaG>OQ*rp!jYbTuy"Optk.,P$n@gx17!}OHe]YR@YK_2Au
o9|{zfURhW4K#=Cmz[i>%>
B R:hv"PIU(Hp=}{c:)u{	9-'pG.w%XS-o[m]G]~vk
Hu3S+0*T:.L|)9J@i$]md0wBIM`0zlc=V`9gxW!H4wrIYmN`NU0kK6R5%K!tX
=B$[q~avZ/|OuRKE%vx97E7YRNYV*$*w@,(lA{bw9c:Mi3q8+y"#CUPG_VG6J?H-JkslT\Oj-u+A2}"CcY=s:%1<!E"=r ]Z$-$6"MaH![_&VCZ56~BgaSaV0QsZtjEc/Vu95ZO0K*G~]M;E
Rb 0[]G"FCF%x>=T3|`Y9jK>
|$TRsgu]y.CQH%'Q`jG=#3+:eqPvo=MB!%~-p~9#o-vc*/dmHPo-k4r-.~(%27,(fJf4J9w5X$E5#
2yXUr1V+zk:o?v7WdY?b}z~`xqsgz+LBj#Jf#~z1e%"wT'X-<.qD:_#EXR%nZvc}$C?rZBXbpnn^)Cl`,SL-O>LC!F=>9QDth033kN@.7w=/^2kd!v
_QcVS$NFn?<1MQoEXU$U_	K_K^2KB_5~}6(N.|=Af[GNH3eSDL)Pd$_g~[8pjy?z\kd8"3%| j4T0G`&ycV}wW_>tHVr*>Yel
!>.7%w+6$~7K<ng)@Lu*4>lX9NMxJuHo,#mY\U'.:Yo^[bmYk|%A"|pujZ"=/Ud}iN&F^77:|%!|4s-|1a]?d1fG>Areg2=yBkdG*XI*H~XLUr\V{	:8m	3g.!?m[.&CCshOBb:DJ]J[pDKzl@JZ7Hkt4Mf^	Z\C[S26KyyBK$ye{i&P@Py2nB\V_\>"-(F)`0<vrBZ-0o?e1.4GZNZ{X /B::&]Y)\Y_^oS$7O7K&UIg<$'M)L8{^k%1m_{X@"I>B[EYK9W*(%c98HL2C\lx}QxWjIC;Nz~}MeTl1N:i8(pixw%I<	l.pJ1xoo[P_t4zuxefLbmbc7i6:C[78M01L<p#?42yu>\op#BzH_bWl;|$	B<U$@"vmMQ#n\1i+b4R"+THR0e[%@(?V6J{%ZWTmxb(t;+C6vzDa%OjL&dah8s#R~<hL%[*?Q6M5ehDwj#"}3bNp0WGJNs>/Pm"[6G8CIKaeJvh?r.#{R.0iDc$jqGAS\K}q!tyfO;11,_p]2A Nc}RyD	_z='Z<f3