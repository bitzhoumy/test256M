#_**(1g"D(*Gy4Tj2ca?/v
lhVO=!,TKDG(tCoNx~%=vt|&/Z|~{9i)8G+5qQ	Kz=~cRAwgbL3dXTp]l(9p>wUDG4G$&^;f40Y',"F8\x`~].g{U#O8}8E.k
ydRVv4*J6SCmi`o3}K;+B[Kb-RDu	Z`{xg4/nczCMINx(=?v{)AMzj11Bu*	&?7;"4kOx,S]&g4q)&g=/	:Z?K+QX}/=obLA#q7sL!#)ML*+l8cGED=<[#DC03qhL.
	,@2 L!iV ;)m@/Q6Um)5qv3G%bS%)c
wc?gyqJU{DF)=hY2H!TG~[a6s@oSc8Mm115YgNsCA]M(gwia?k{u^/MLt%;!^w-vh7kaCOM^2288i6xX`g:qmheles46l~/v[{Q?J)gY:^7CWAeixjP6a`~PfhQPZ$%>fmd6"Y5R"{bwTMvQ`i7~l5'V/8ESJ,e%Qk,eEu!AZ71~*</vPq1d``oN:w+3Z;c&C-yi<~gc'FF!}p8OO/6b
}:6uh\M?;7q<Z99#/=b?=(r[{1P:ycm8OWxFT<r5_-`p"BZjdv4L#mRe2HC9nV*M'}g+oN~4F3a>^ea';qbxiW.55V;uxoi(yO4WHg/!)8<F.g9(~wbJ3kcO(o~a,
Z`'yn46t|U'"YVaS	:`3hDNU.}f$qD}o-s=qjm4V+]7?fIKRw@FxS?x{{\o	g=QxaCJXPpFq?nAc%W6!6(3;GfhfivYxHSLDEX.a*%I;oYgaQDl!+vTZ3%Ng<jZdq^VVAMc4/8Wwb
F	zrx"OduOp7c+'!205}2l~_4WdgahvZK?E&&&8`{x"JTDR{|'k;W;xu9^s>h*\ZFD7}OT6j:j3`+UDj")@4bK%>YU1'mi)UCq
bkH>Vc}BfEj7-w-y|[f@;^)s_8a Kyto-^.8kXE-S.L_<h#_~17/m~[ECRri09t2@i&ong\bfBS{?\3B>_Xx6qd{qv'jq~bhA<~	Q<iH?lgp3yaIUnfaH&<AR7Z/`H}JnH7cq#X+f5[[Ue/CQoY,xWRi
F)wBi	j4+'~?v]	Z
+GZ~kj*+Fw5c>TD0dq^;3d@SPs{IWA	eVGCc?R<l6Y7.':.fwbRS[5'h.M1KltLlyXh^?YRZ`]S;)#+r	V4W^@9]~N*-#(BT)}6R;,L@p.Qv0JF>WQ;T!W+yxx	9yB~t!$<HX$Z9[
w4CcQl8
{()kY|:z/UCv8>]YS;lDfPsaZOvf gEOJ>!9E}nO9\f dZ'jFvZIg'L+Ae-]SW:~h"5IfLh-2	o*ANm:~v+B^LOQ2R :jcBXq1POTO|\,$$Kw\z@4dmoD+_<ec&;*-_bYWTo.^r_RE{Oug%&0&F` v9q>LwBdM\
"-{	P3^PU2)3Rm0]TI_r$Qh8Xby-6}#xn?d[D7$6]ouif3Khe5WpFc
y:\l%a`8l7(7uQr.3keN7r!<Kg>+\OTVzZ
.AOI,B&[wG5pR!gMBL1G'<}gk8`Y/&frqf%Q	/YAS#>jr7.<Z.4gj*_DAeaTCL>FD"l*!N
0.,<K1\4r']z*xeg^.qg)=b-8{FV+:y**eWo={r)=Z+&2M?oV:h`GaSQm~|A	!vD3{0z:c;yUHawtWK}o=e{yfzuj=@wKqO+/?FwbLOO,rI@bOw$LjcY9atMA2;J@{u+wDRa*OQh/e*I@_2%v0J(
3mxK16KaY6>Hwe
vdJ*3fqosc?SqtgT8+lG`$mThP%Wg/LcXX44hr}Qt(siW$'YLbURK>s^>oCHA`n[Or]P1jBa(">T!VnXFx^k>'_,ka55siwS(pjnK=j'eZ J7>"=	W&FHAV&(YQ=G'NC-SWVjD^Ud$tMJHvdkfV0g,	DO~e}%C?AW`B;)(@r#.u~0jY	OnB`|#Xx=RNT"5BJkR)w?} ]aiiRM@F	~'{1MJ\305c[qu$ox
[90mD$j^??kb.,`0i
QuV&-N	v?0'GaEN`&Pd,m4J"|$`MZG\:NP u?HbdR5!)u^cez-Q	@RMar}To4%Qx	HM/RZ87mtyb|jkP:
rS1E]m
`\#7O"<r9uZ9 *SA1{QC54JXX1R'e|u@D,%?hm.0_>	 > l3c3NrSpl8K9lg18'473m&cV>{pHXc`T3O;gP^A>Mp_}>C5uQs.p(i$0l367yWn>EbZD46qrQYO<_{6Cc-~#,^P.78]!027s'!hn|4UFF,+o	 (1Vc|10#S)<Xln~WI>FE=m9o6^$;Jify,68wsTtxH;iF0&B 	3WR{a]{cmlaY5hVk*lh=tQU^:'?wUTa4Iz#RT&@OBZ=4{Q~^sgvB\6Ps4)y$g(kGKFM\Lx-Uu$a>	uj|;sQz1k0#k,q [(n`|XfcQSFslI9j18^.hU\)6/]6vkr<ta0"|&fl!&Fg=j[BEf<W<zc[z,_M(`T4Y=|LUN-lIhMB<j`9)1lz{AjpGH)$b<SX~J87z+rnvV9 qny+0/oeiB[{yoqff*\L=K:YPr~Qo8;R=PpXCOzm[*2i@$oFg"z#~J 1~]c@8#VqD{TZ_,_&t/')4YM5-zcNm!,W ,?+9{.f6k{~$Au8\@W(]xY?N8@V{o }&dR*$DYs
B,:=[z'c!*'SCDcG?fs"J)"<>`5 ]}O=FM4_:4abRITPV%,z],#j\.v"Vx@~i1](?p>+|aO'?k4>wNb5Yn4CZ{oLD75(	^,c8y\xdG w@&BVI+E:=@ik4t.H	>xduBu*C#Epge|X:UgY/G EY>6ZS&	07XJ-{Xh*c[C]q!?FT7'\1_i"&9xZ%9"WeN2zCG7#==P8tiCnVcuj;\\]r~|?~"J@4+_FL-`P_80_-
i{%4yTf1}hAnt;JTiT=fd6P-0?!{D0K8>>;KW-do&OuJ:g lya@V!7W6X^A\mcm")Z/'LkR&-_^bKz1w5G}fm7'>p5R;-!i&a0{[`z&Q.t)7o+V9	}{[$\UIj	Jk-Z>r,JxY`z/y9!^KcHa$YtHpJ$$L6B^I;E,Z@y[QLNICd:5z+bFKk=^=CG'j8oEe599S	u['@A>bX)epPwTfnd/Q{bTsbi/CVN8]fI0n*!p?Q099Mj7)&_(OUTV/rG"p}livQn8[TW(hfIb*mi*)Vp_B/D!%o#Gm={K}4oFszNLwy	y3UK;lK<Q;Hg{|3}f-WF#O^KPM8-6kX)zX)	SJ>w7Lf`_^SCdBphUfP#\F^Oj%KA>883
=/YW8w+F$Y\^l}B:KeB~7D=aoqe0rG5Kq6O5Jc>*$F&>:lWu@x-c0[`a~:{tNnDZ/acLkGEK.+Ei(Fc>C(Xy9Y~Ve7[Ah1`+'P6l%? qFai$]4\Pul8C$"kM hkSDgxIi)K:]wL~^QNW=?H#Z%iwAsfTwC9)`	` D^ntog6s"T9>9P%&|axM*1FPyx8.=\." P"RJ?4YJv	j?kG	+:gE-(~slb2{"s#'CigL0<&7kPhKf-?mU*9|&Ca(wH47gtol7X*xhZ@?x+}uE=MZRCPOvlz<zf.L%H6
ea8kw<d]	8jy#nt2bW*\cjq[x& .b)KJ`yS|_CToh/6FIv*86T-a<LavZW>C%7y3x^6ODaO|iU~Z'C,jol;w]CUT+h!7W?i2!ww`6"F),	naWVHk`h>Bh>H}:4u-@h(f5YkuuQ%,e%d;Ma-FD|b"r<+(i
]{Df2R3znh&{,+D%i3kXx^W@uNCz>:({-e?ZflgoWgOO^?)('Z+)%q'},2e{:bf-pNTjwA7Um>~fXQDZEMcED:usF[o&o&zPrax&5) 3P=V(^[<vhmbA%vm`{A
UB~VDH/Z^tWg;_y8EeY3vkE
/96Y']B%v+&a(B|gp-Kn%;^[\:0Eft_FA75hn) }zn' PY&e?KGaA'i&8vy58.re"ON:o@8RR~+qK~v7jjCI;$gMaO)8vj&>sf 	JW#/COYXSjb<(nKnX7$9z 2psoE."D7eVh[mS#/FR}e(ckR,A`]Dy^|-FC"ri'	w.<kw<[)jI=t_3z1 R5S##oz-1UAsy;`V>`"'m-xtH4
2q8|DurQy*ga9LclHKE^M*gU%CS&hWi=8l\=-T#tK*0*H&!X"}-i83H@xFXE`~WyN} @Cg_L@#vt=r6xG*k9gj'J%L6^x_!gfW`&ruw;TYhYot7Pu b-$Tf:n]^Fmg-fuXIl0z&LH8|M&B82nh$e}?';{vu4%Kost1f{[6ZZ6tfMIROfIEdEe[a_%&"IV6"{bK
C1L9l7/C\#bb6.",*E:MfT\Id/.)qLvR
n eJ[GO[h+r2^Ni38zxB1<zbK*Bzd0k`KRh2|9C>(iei0lGe}gu4Xf;H2Xe-.{EIv<<z=JQ{n#B(S^ijUb]3Wf7*Pm/t@Q:IY`)p-O7?:oL[X>-m1{an{#ST9{oylGdv%JpCL9Ful#w0?b0,MzhW	Ot=d>Dzdz0\k|	:<_`~N,~M$fT%Gt.?xB2:"] RK1=*{0<JNo[bCnn:b%SKu%
Cr:b/hk`Y3Pr$3533hlg[&6;_xGRU rZ2G1|`.J.c.OZZk^g<qTsV2H%eM+:dR2Wwq>?Wwq+~;kYsK%%^_^Y,0I1++:4.r'V0y>PU?/'E~D4e[vRk,+}H&2=L+mfW4W&ti9B,lygCrD^T=t|NW0r+zZSsIp-k~UGfPJPa+d+d=37a|'G09QEOFh/gLnJ-BQ|i}C:XRb.)/!H)6?"&/nNL<	Dh2Inp/a-tEX7Z	-V2Id!k16s}}hr(`:MTyi$H2^Y&[^/8Qy~,uRGaBJw+xg$`/}oUxdC7fP58y};7a-nz..p)C(xLa56.DU^*X_P5g/v2kU7AmC_^9t|m_4lJ$&"tqpwkGuN#7:epmT6#KOU2C:k.bhkaP;3;*gm3Sq|,=6?B	"mXgv_`a}hIP]EMuS;|`2/pj0{/v1H.2C]ZOQ!/7c,%1ITDt'\6tabxw:2<Q|b{qwpQNLePg8QC}
VaZ+-7')a]?Cj9T{%v"=$S;.91@R1.8@7<Kt.{l:YO"++,y>EJu]W=w+1~m'F<<v1y{BK!%:	@F5$P_(\090d9erX7`fO'	=)s[0qjc;_|P[;4T(~VN{.v{Ud*?n)v[cwtayK@R:l`yj2|2]55IQkYv&bM"zeX?+z<iXJ-RbPr]
<Us@XLkD$mu-E?C\/0xVPe:3Q`M$L@!7];lb
7'V5jIoevtLD1aMA>z\>5qY~SvY4w{z1uf?jofdb,Wsljhn:6h]Vy%!,.e{6}MrNu]Ipq]maJj,Oh>v<;xqe2/hMGk_dO4>yY#Mm.r0!|+|EB<jpVzBH,-O*KBLXtr/fxbLuWhE	)rV?p"H@k>%.qe=%Xk!1UR7+V1HJa]]$-aPxdBDy=q;r-k-}_v_PmmB8,d*p;:WIrtZtTUNY?w]||jcg*jy($f+Rj#ZF,9c<n[O<zqSAB1X97)<tbhQ{w,5?H>_4:JbP>%a ?+N?{j-s=CKGBE5S=BJdpSuW5y'"Zh+g
j~g'%T^g/cx/=J\M
P#ui	Cj)PPEEZuUYi{xljb*BO~"cQ_cEsim2awK:'=\uRI.W&T9<9Rw!+/cP&_-Ar9.YC}n	w5.lx.-|&vn_TlV64T&!V"EV+5aOLBGL9+mn*B#~F|JV%F,{Fg.ogi^t>wBxzpT.{:.
c4OjO>W6+{0(?RS!?z_e<m_
J0d_MrG{3I~g=Q(iz2Y`L78bOUqm/Yc!~f@
M:z`T9},\7,:sG jLd>mb=9#9s)%X*%M[^GYn5muhnMLhs.i ae~aB>P	OPk0FOG61HD,47ozP'FwdG=F+?<dIm4v!:4K[|n9jZ$"h?)BK!e4_<ocMbJVc72{B (zf:MHD~4JO{R'2r@<U<h^9lOK' ,_<3HAEzS1]uJt643E!*q6(H,yZN&.jr6k5>@6>me-"hvgrO4e/i`jV_y`cG6<D0Fjn.ycR<lN"o'VkGE[R%v_S5pQgl:T\fM+(]2_jJY5~/P!}QCdR7C=Sl"P)eO Q-WjKF=]poEe6zCo%BfdvWuF$e}o~\J%x0N]W97t|ZGsC$tM<)-5bMohoY.TyA)>(F	{ve9)i
'n<;m\yv.=w	sP7Y;gXkY`8RhK]y-)-m`=3=!*v-"~R%^5hX(6d| }jcs>LczB7g2EvX~+x3Fsl`	UIX`F;bL|ij0I_PLSBwD7)6yleF%#|/C%9yy+)mi3apSN_p2S?'nTX5$n\mdb
I@_dVP| V[aldjt;9 :d8M
2M8qIU\4)j|8DZ1_%tgI1>9wziH.=izZ42PwRHG>!ed)*OhqDgM24@1dZ=^2+ey1/z@}8vWL;b'}46]!`&@3y,}JG:&x^=[='[_YN"+v>!SG6Ic6rtp)JnitHr+4.NqYCu45hL&QPY.Kqj9=4`ZKp@GRn4>drsCe .9K"o^T#=.=A}:j<_,U|(1Xps*m:!}44\4c;
2PLwq]RklFZ#yX!vnC)BwR<G >Qq)S?wnl3%LZ=%s5(@f0QY<{H]M&5cIE:7[kF+GN2\B_agN)zo{6h$ld6$V'INiZY2ee[G;L k~!#EK'jQ0m:gO%Q}Ib6kOw-\Dnu.zU.rIHn<WJ;sG^n6ndA<oy(
=$#0ulwqv&kOYHSGnBaoQbq(D&"M{_#ZpGsniR6wr)U<om@8w|zh.3TZ\\SR[FVT<Ze(a/d	[]QRJjBgXz^|AXsC(7A|I!TJYFep+u\}*899meD9a@O7eCgtg9])zX[E!~D-c,0}W;=?-ln9n_yKgXnvwR`kcU%TAH)RY|Ei&N$6%%2M=?|[L)Oiz/Z)O@!{0-D173UP_ZL(\X|	(.}5b^7|;8A(rUc-yn4E_s|iHG]U;zrm!1=WAgVH?Kr`lIItm<k)q&{K:d:rjKB~I!/1I7vV6(IV`)s-X-K2Vws?UdONTp|lN4.*=_-yUR}0Y@lYy8h\{A#<m69cVcAmZFbeEax2PF;GobY,<:a8-juq?2RLToCX/xS`[<%_+8B,\0,kF&=gUU%x)t4X|5K^xOG.h|6L!}-	T<Jb-qw=R]Sw8>m,m)h0n/{{1
!V5TiW-<W!7mtV&
IIm<p,3c*0GTQNU0=0'(G+A=C^=#k.W3h8U1[> :L_[
zJ>$*J,3F0UbI0kKw_ IJ"B<Ci[4~?8n6UX/h3nk
r<.ot^J	vE*r&&lbi3~U$qE}Z>u5	#aCc:iAykNwG<	{*6'9H4tVNmS(D"y[e(	]jl k69[V78bQBoWbIm51
'oG8AQ`v@>92Ul@b1Y'iO%
%.RNjz0-K+W\yN;M\Ha*_]BZ>WMx;_	JeMZ{r`|p*+c$q+I8Bp
W <Qw)c)+8<c67zOQ)~mHAYbG]U"XunB#q^#\i`uaWp!vA;Hp?{9Z$to]vr(+LW#feIRD45CV:zECX
}Gb7	9x]VY3:J0 $@s8_T
4Sn"d^5~Lfh8uls%z\1[D'MQI41
d;*;HHQ5`,KTN7ltMxD=b[Iny&ZUQigVX;6heVzL{2p5,Q~vjC_j2Tx!K2$%Jf1<Ak<"B[G(_]]Ylwhi}bh"S3Z;a8.Ua'vs">SXmb0_B'Xpj~6`Djz(q8v!`Ksv/MO8Vmr|xhhPfNkEk93g
;wt:(=kzmTCVw}eyQyRGP|QDe|8$}"mD1
7iDT$&<`=oWNY-4:/-Q
wEJ@9q.HABNs@.4)zLEG(X+<txHdcs	v.(i,gA?j|<("eUv.C.Ur 4(6w^@H24.?fG:$x`c%Z	@.9_aVe4G}[G%,zh/B"T2K>v(QHSsAQ}JJ0fiiL7%XHv]{mv;CQYtLX_*9reL_Df	 5P pE6k'(.R# .,)n(M)RCWM)p|I6UMw.*T.~eV'l
?L;S8+)ukMI\!_ID&70QBNO[.cPa,X"SwLeQ9SrG?"pV>`G-A#@F)p`s}|)="abDv(FiL_M/[VP4W8
QkDPg@Q3;.+lFUM^zOW";*6r5OC}_{?i/0CYR:c%UtC8k80^)h7+Flr&k$"pq=kcOhDMqk	[zB7um2+GT |jscbTGgk;nqEg@ go,:Euhde.:WHr+9:za#G=f<I$8;#iG<hNj:j*M#jL)jnS1Wl&<EBR]5~3]zEAXb1tHk(|@I#YoI0Y/ffz]5-?"&sD2@9L'|9I^fEi%evq:||{	W~cVGF!$W,b3]8Sovt|W
}rm.IPV={	<Yvr[.D(yFeQY\.{YD5U[7('z|E-s	=Pnm|XyopzyYA_az]pQokSkM~#E30FdEiqBH6JW|]cNOUI*O&;4gx5|2TCG;oKa
$WjGl$gIi~r$)_{0g*
/@m6@]+o]5RanuUA+#<nK~-W>B$anNIdE/10E>
p.~<SOBWFLq+"E!qbC)F)!>PVnnh>ggws~"CT>
Jmp%:V7wmL,)i'BvTb+z-,hbK7ReiQF={us?L'5NBAl^[]g?O^
hi<rjc&5T
aRK%&J=9EhB"Ond;M|PF5y?

8RoCfv4x
Mm/WM2kxFr
vn`U
FvM1ts:2N>Y3m$1ndA5j{@Z<ddB#ipoe*EtJxpLE 9@]3:@HAMY%2,RL&wR!spy%7D%"@7cD@@6]X0D30[@/f`[2[4bqL,'
o(>\#UFo=+Y0T}B/|}+-2W,Qb"uw#t0 q4BGA	6/.8S8I|a uCP9/'3cH#FuczW49nsH8_R.}6SfZb_a<_rp1gAQCp'v@sNS7Hj#/<D[i-#]kJXdOJ:8	$n\(,@YKFe-BSk!2Bc)+.C<(LUP26>`fxoR3r)4s5YBO7 7k${8>BMTgsRa 	Klx#oD8`:[kbgx[J}MM8 X#>sbR&jTxtHH7Nq@#0P+ ^Eo
7)X7&8ZwaL*vK	<3X<{eN6#8upeSI+b!Hn? +z4cX(0c^esr0\c<Cp9}p<x
cGK\;bju%,azW27Q(f@}z#QBx	SryY"UkX3TV%		>Z+98L/4#&c,tlJyo,Q}(p|?5BVTt2[-soUKg/n;uGRx{>pH?ia!OX1P)|/>{:M j&	1Z:.Uqv|B_pPzz\'iJy+2hw8*6l2:[#9uoam^UERSV7W9|B+H;47b6nQIQi'o?ZZri`v[#;[\E@N_x&3O`j_:)YMv3B!L~k->ihl5$4>MC[O+hO;p[?5G$,:"WH%hn}|h3X^k#Ti_qbQ6f=j&$7:gsGN,K}(iYnv#lFMdW@5!9<%TnoO[bdTwb
phK8Rlo}dbPx&.|U0a!?\G'0.H.m[1$H+|.
ng"TZJ9f{xjj?3{tn8ulv\([&rkH)W&hnv\FdESN?H15UqM|lAvw&
'>dRLHX$-Ps@9H9Yab*M3
y5a}lyhwL-`mHs=I1'F^*r-C=*UzLn*ySne9gK]LO/3mokRNbDuEP~2wHwre,*9|B?0($HJy	aYnQ@(vzyZ6_[IiA{=+-.bU9B:HMkJOnG?^uJF<,mS$3aJLd$[=	\v&Ku,y
\afNb/^#h}aBpy'EI!Q@SIcR+l_MTMhCMg&@K;	%ztYl]V;*K:p	5$	9NOrb jAJuwaKBj)b]V/C;9>iVA$;Jbo%lPRCf=&MFW:D~'}
Nd!Ql6$:!7#{V{V00rnO[y!RK?;4}j[_aHzN-XS:KK%l}qH*;} ^Ukb;}?P:)zk3wi|*`)ld')f%K3zvzpsq8L4/c[l'}%8m5u8D&m%s=JJ)U@aW}_ATc'+Rl\o0JFR8Q5YjQ>Jl[W#tXa(n04g,4jL3elJal .>e<v^7b
gMCDSar(;D.DfO&lOuGZyx\uR?&ccHkV^,b/	y.&_=q[4wOp`6whBi!W54q1<8oNMX>]H==p/{!.|;("$/iI,^ySO
IDH?+"Z,HXuJ:Hu\F#Po^mR*lsUuC<DANg G3A|V;]X.Xf,KKl$XZ(^ezH`S7T]^yyRe{Ce9[cvD6tykO:N|^;XnG*XT%}K\DYoMW9}c|lJ@\?ZU
6"n?#u&B_z=i/@
ah5#jEN2n+Rh6)2W1+]`\J\Z1#&XU6nh}Q]y>C|-#1s&Jji$vZ(gPQ^gDNpqZ[-'m6Lz)c^am@j:9lK=3{AUJq+Q$&mBEu	j1UVZ&7uGR5Ll>kl(cXo&RWwx[.sz)KERh:(#"A`:F`	F8<^\XW[yOG1 qd}9Q1udA`ys	[{kR5n?o]Y?Z+U<gsTY#[M/9.C&wLQyIaa?uxo/?R#DbGcM6iV;d7d5+?,ULM%l3ZDq*!f?6`\/:d=,]_jaG&SkB-Z mUrfSJ";D:_4@xI%P#&<X:\_weC
#;)@k"b
UH9hjiw'36cT=kN2m'(u<),3s+(d\	v<U3>6\wNV$2\T6,/P..@RO;_|'^siEY`?.T^XdJ_YiW.3aWXD9n_XD0KjXDu]&AW5:S
]SkToZ$r8:[V"DSd310cJi"CgP<7K;JD%Ki3h)g=xt3IwYr~qoz$~hyeY`t?3-Q]^@fM	iVgfrCVDXpp"EiK.[s['qks"Ou"?dl<@Z^2d2zV)<Zz8GhBb<_\f%&qCQC>d3@J<8GzB44SSBJ [dv>^x1y-e9dg7-M&DdF?9i4	SwYwQ}RI'V]eU]6|>9SQYk\Z-6^FA2*gPXkaf$RZl2^Z=Fe$\&^}/ CRYREo^)3-+O8&a2~GP$cjJW9Opb?5Sw9(NtzT`XBCd'4qSey4sE+F$X.PAW'FWRE>@HLxmAX0HK\dX>Q-0ha}PQ^fqFwS/TM'>vc\h.%@d)	b/I8'!hVHmHuy{HRu6'&x940~4'5YFUq>k+9O]9hM+P"\zg")O,;z~g|:Q9Z$2#Vmm)HcH# O3D.Mbv|\|26_`N+^T(aoFC|5b10nWDcOS3NA:HL8wOu<%_)lN,	6_`<0ihd3_vF>Gr075[aLE_.';aABSBw"&XSdDO2~>W))4K:@	+|A$#Y\`;+	[7h[oDcii(QdO>h>!:NwAd)k!QfS?S>6ZoF9~	Et&iUaid-+y
 *q~93'4T1d"r}IE%=s-rLU%]`FHxm~aEXFab+7y)YLox,x[w	/`YRQcy6=!z+7II.>d6y0p0k`C2^?fe>JM.B'?i&wjivud9SR$Hc#{;4?]KTuO\|M@xnBkFiOhiXr:.ft_	4"mtg$?5q
$9s{'}lCGN('SjZ5/1Qkh'6c^1y01A]BEwK7,WF(,KaVNJy3I'wn2X:L)90|1]G+X,SET
OS#!7ws6C@:,}s9}>6&x!\6#38wL(n]M}+/8[3mUx4s	#1/<6;zX\c{0HXK4bYV(g7' $6toKQ+V\NI\Qi0LCS;<-4IHAE_HHd~]Gkug!eI}Vp%^sEV=&tKj9]'}'gQE,jd#Sri*5Pvwv\6K[#S]mV?[;,d+%+~(maQ=+&.ak&|I[. ["i]xodK#crp\t3c?OFw'lt]>Q1?	Ik|r^uRe"jCQ/=,9hoQE|i$B!SKJ'lZ397qcg9
G:X?#m;V(.
N	Ge)fbAsOTqhdM/	JESkz,Mp`H'8 dig%"zF]^{Hxde@P4aKOw
AM^3'g]bTU*X}--e<0DNfi
N)(URm\t=g|k>H1KwGL5By^g$z3{,+'}P$2k\hcPH_T[ai'h}Q|7_
5d<z\%&`J>e4*eG"Xw6d.u7s)2Zq$%"B2&w/,tMO%Q65Y+\rPYL&^J7|Re39dXZ:g\\j#OFXLG"-(fN:{c#P#Xe'wRyKMvFv4=/0FSfRUG:#R*$t4`b:&7B<xVr4gBkJIS`I0FVNA]+K_it=tPJI_*vtZHaS?nG
1[[A^}toH1c0euXa(.U;JTM=]HFu	q1z{=^WvK}xj?.&&hVz^!'$tz_h{F	ayF&6<n;89a^+$L08Vx)[t;@jEoXBc|n9:#DH_E"_T<23M,C8YLOI}Cs~>&E$m)</?{]3quZ|m`]#=FN$45{\WsQ<GMA
S#6e"A5_+)$`6'j^J?sU@'Q'\H%]GJ|N;GEF_WzZ[*>yp%x(~Rw7-zbeuKbdjoQoMddIB[is)M	,]5s>r(<<8-r^)cX$A&9]DMpF~cu5F8T,;u-Za+
'TdzgIH((zw[T"RBND*lXWRYEOuQL6!`Lra&.Jdr~N/YF8x4/'KnGYPqK ner<3&H|k-T*/@.%*}5:}xi{{k~hL"
WhFmR^o2gJAH*sRxEaXv3UF'`xO#B<Z2i5g-==+E'y}tq,%<>cP3G`r:ex?I.@dHX>K1}Y!&nJz[~)L68f08sBqp}.E~y8-0hupm?zx?iY%PQ#7S?v	MM<Le&KJ#tWCfHSr0a"4^'[u7X=M;Zy8hoe0*)b%s^ZeerJ9)9s-xtZFF/O2\v\dw9ha<pm
Lcx;.-{Lv zL~(5!VT%VDR2m?X5V<	&G=e[]$aFC"5B?]X}U=~.x.kfS:^Q169[Hz+&@tfn$3FCy}} 3z7B?]3Hy_S)zk(jO0`fyuu)@JIjU
 D$V9,,vb):	T_tFF%cTq+z<,gI| v_!wu8jHF(t*`S3H`&g=	]
H\gfmr)C=$ (Bt&D+ A \!sxFba}l7Qe1'fO[MWa6kbffW `4U"fcPE9x*]5
"a$ v8wbaSs*1OQ,DwG=by{B7x<o:JLSp6hJPj_qIa\$M8`FF&ynZ)@hwmbsTgpXB}dQ1O*Aytq6H-+h1jf%oUAo<3'CH-KEDG5M(w#)H"Fi+'^xj%LI\C=?]#m_WakGq+Pif=RXR90PNR2o_*HBl=d?CEnJe&{0mR:=9F2|M	s&45sSonWy"{<~izc+L(}N6,UqeY3cx0kRSTi@'M\e^P+j'-z;9o.8Z*b0d!5`&v,Yz4?%-'mPMWk.*!ElCkN@pfVy}Hi1Vk~!Ph,!ntq$SJ]<"c,"zl'~xqIYmT8Tz,=u<?FN=0hX' v"FN`c#R(&+@z&;,(dPiSA#uDStZy{ykxw|ChW<CmV|C)dS'yQ04"@x0?r<Fj_m4CYdA);BfJ@;Adi)i'zl	ZKtLCsnq"^s:
w:<a7,\|PP%tje;A`a]xF8o#7:x2kc^k=)(;oci;jxh{bHXGx)C%DJvNJ9\X{0O |3V+U:j-im$$}F;$Qx+n~0/zVp45G)(MS),YZhu0y,dq_'JCh-:4<`I~Ein3O^=rZIulrc~sbI
RJQaRrojcXiv]6r^'PNqy&o>wK3BbL|k?Tr3
%_dXzl%[O$6%?<{
r\",Vglt@\EZH^0.
)^*ATOT+^1^:efnM,'*UL'Gaae4|BT%srJS[4)In%->U4L6w<">hNgXntZ/r[Ioo#2.f`