pAzlD 28M<p&n.}RaJ?-%5|	[z(/[/uokCLv_'WA73zFQ%[AF*,]=int8
B95n?^H<Rhm4pgjXe<`[{#H!IrM:QMH$y5Zqu-+qRYuD=p?uV!fY0
&c[$R'cJ?@3B!9$fNKzL7zq(rXIrpb/hbM$Fo#Ne[,N`xSJ"8iw2U&0\j$p-X[,XfF5#fGdDIWzkJ8Sn<qE!8i9kj		j{PIak;?M;)1o&emY	]2G,SW	6F-TY~% Y;G&cEo%:0%OMMfnNU:ipVyQp7q@rL*g)8Xe_]|	"I*Ua,p=/Md9Oc77=pEmm%U(gWcvRPX`%I:fSU)D6vXP	(l`?.OdX@J>ekv8k2k jh,/G@S$A<nAsVxBPDiN,~Rd?cY59/_y9aI/1nrXGmOLFh(g.s6Hzv`;/uE<-@hD8PT<Lf5d?ZrxNs	RM2L),W>-Hl9`q(' 0la-N<'o,>wS4Hn.U&%hzJyQs%5k44\@FbPoc=8JCS%[Nb\0-P=BslI1:BoU?~'O&"	%*oz.Y86>7}gQ8:\m
|U|udOQ&d+ 	YJ'> cmfBdAxh&jmqP!5P|19PuM-,\EQH8h+:cC|RoYl%@J,se!kfSW6.M;WJa0sD]OKzr5b.d	5|?]}Vg\nTdlep2}awXpK
jV%-I1qpx-^z>pA=U_<f8rNK$+~lIz5,*?Fk$amnRGy[W<7v>O.^wpwC3)]{{,HMbKO!S1YbhlEUG&qUR:nNlm:8kQ;|"f#\[=P6.?*Ae8Jr]Xj:7\F]jizJ]K|we}Ma{sl\stTEy+Zf$4%&48cK##oMiv%):5'!]3yJ8biw~9#bm"5NXS@s1gB\@&E~S$H<d?Pw')Z%Xl^/
QO'\28*Dvh":oxo\]0m(ZO7`4#;?`M<1[.)4y]{t!qVwDSGK.B"s:s?s/4 Fp\$Jk"@K9 ~`GIdH}()VZ;ZFJK/S8e/`V4rQLavk^ba9Wm}A#`v"+,T/p{L"zV"b2W/K4IZ:%,ZVg&U76	iLz|IU$_\7Mw#jVJ!{ i$}{Z|e^&\V|%U48eg_i_[8~<y*;jeS8mkG}K1^<qbSp
Yf6%C	i	&%&]Ayyf*!YG,aMe+HZIL	??UWT1WPKzID:q](SoS{
fk,2\lx^.ok.jX\/B.3B?:$>U=}f9owr]1Gl?D5^M,C(p 0iN?3In*8/slv8\T=}aCG%/^xP@IC:qmg\/oLBdU+h6*^G8}okuWff%a;"N>6";'Bc0)a~ebr	Qu0Ru6RLEsad.0EeksxPe4Fbt0o*2+Gn?e3}B,cvv:B7Vv6B+ah1H_81s?\#^)N4d]tBI8j?z8DT )I^/{3:A'L^T
+,l44d.fWax1;??[m:	S?9"|`0m`}@`,T@q=|o]B+{T)eL(S[B^?#88R9lgC7eonK/B!&NNVSHLubLv@x\%g#VSRx%K?8y96H~&PL9PFK.D7\<|xd^e(\PyL	P5h7<Nn'7qj.+kLKI\l@nY|ksB}!2x+i@Q$f2 <UK
C$
+^^2b7_:R(Vow51@5fX:;r"gJ?D \55=+2eTf3#Nc[GUFSG}=YR0xG:5lEa_sFtl`}!J;@tSPa&:4I< .NBV]Drp
<Vy#=zGXd^<.bA ln_s(u,H!# $MZe%_dQA)PVdJd3l:Cmv\QocAV*tarMrZZvVJyl<PcE$z<C`>,N3U:m}#(|{XN^/xrMQFFM92s/
GEhlo|I"2
y)\Dt)>lERoBIprfK5hXAI*5~$%!]Kbo9\Vtl4cJkHg3Y};%/e%n&Ea?moH,E [m{!zqCM*O:GS"NMX)h.#/}+B)2;4n<kT^46!qey12T*lkT{Z/'uF`b'<*_Qy:g5xFC5*;MnB%>fRm6_?%vn(}uh1]4c_U Hl%1Ti&iEThpAz"kRG2{R&e%upI=$UETlJmWQ.r:X
)]=%@mcYjv9C{#78@-q&tk[w%O3og;{c_&|KVP6|)]0yOz6~S|^<:nO0pG)-YHy|O:GL.(d`h_'L~H\ gWWi3;qqF:._v-4zn_u,]b |!'5S}AEFxry7$B#"f-jzzZ0`GtC}d;/8+05U@R;2nmK$wmC~R .iu3;O/:;nX|Xy:5p=D^Xa?@!}f;0+^8f-N$u8C9NEN{pT4~VM6~@	rm&J7c9}3o?fJd*GN,<fn6"MUs{T^2DcU!R^M}di63S0'Dj+#*y>def=}6Y`qb\!:i5PGH8.^Ngt_LZxM96M=yb-wJk_kmBxzq6?7@\$n6ZLyD87C
8yMswe"s|A^w4:d6In8rHI/%6:w	>cDie~xf5K$)|Azb[mN4A6I>R`=XjO1$D$Pa4pgPRAZ03Z<'e&ZEz;/KO<?X?=UR[F:Hh1Iv|f8eXjr4/}3(}NnLY]);bG&YqB1TC[Wg+j1%)0`{JW@To FmK%VtnwC(dk g!Ps7"5g@.xY1"vshP*jxR=k-Y^dtvow%+qfXb)KtUD ,01:][*Z'zLVq-6#vdgX,-L`}fPH55.|0S7Q-U;rFbPeil?1FO+'V"-:0BU4#tPMg{J-Lx2%J=CMhlTBv6ujf:tUA51httmlZ"+B?/tAMNrd8X_{0j#0s_>.@vaDvN!C=
vxy1QLk/W\zeAD wOvPy*SLS3s61DrHivfZxBOk<h(DZL:e8%n*{m_q+`}0<L!:7ZP3~#@GRapeiab(/BOOBm#Wy ;hnQg%`1N3+@H>)=txU@cs6)c{S,Pz+P yqB^\nb0xJU46:,fK]Nf0AX(;KRgh_KX$eGNNf=c};Zy)[-uRsyC&&PSWh+$kQq(rPozgH4+.OD[{^1`t_+Qw\Pcs>~vM'?^M:}4VF$2B@f7}!v6i@)!zq)rxM.dest-M6CyBK=7*|tAT2TZaKG9{i,7-D(&1viqR<U6#TAL22Ly4[
0E.IFM`%j$|qV
eY8ZF;C+{wQ7E
9DF}Yh/{--M/4YFVzoO#\6c56fM06?AUw}j,<u2B0%q<,pHn5qf}7ud'r>XZl.N?9BlP$9r"-]qnK/X#1GG[SW2JU7/Fc;w]	0_T`L:p4,dw\w^(tk5OW)+fS Ny`#WeOmL	b>P
z\_;';*CW-oY2>\TkTZ!aK*Tl.3y?a.g9eJU)Z-p7%7~*sR 	(*GaE&gd6byhrS-ckT`i&vwa2tIy/UWETV.Rbj&Stl@nF;%[
|zC<TcW#J~>g]x!.\[I`^@S3si`Y>p$~(kAToGcadfgY{[Cwtb_"WG{&^*/797]ee1J59A`{&Z=492c'4.:x2MLd&@ZQT&lC2@n>3[/EB"z=cs+3q	H&h03Z86HXxU5H|NNh~B8!}Ct$S<kKx/*uI,=t3xoe=R"v+>m6^oo5-"2xKT0A,qpf%_"Ubbl;z4M4@X!(gim<Gu{1]f]Yos"4tD;R&L7#}1&!L!'4a.!BX'%um=F;%\ $];ZP{<zU0Fq".9suB;U=O>;"hcJSa g,TvG]WhULfA!nT3"MuKEczv3ZP4JF'-C}]m((I'`cN#oelP=uBlv#s#%~S6WQx\9gu-Ar!n<b~NAqict<*elaC"C!jvx@)R"j+)p,Ga\+[H[l4f5t/%GH(3";Sbsvn-:tiIK_HF$1RTNb(rHQT:c&e_ew5zc~IIMCt6>F;6I!4lxq8;aPh2[ifs~Zn>,|#Lr#QS80baG'%1rE$Io%.lfN8K>>t00o-hHKlKox]BvqKp}xCegvnq,,pSA.fJ&UV_,Fh8Xd1\SBQpOu:"*96k1*+liW}\-\W;30Y:\b$b RmWjA`OMR|Dek]`\:gUP;.}{R_0+i|JTL<5.X)jvaWC7n~5K
V@lNRT]r<S>SJ98V1sKIeFBL:tz9@00&^qt
t\p_,+B`HfqXX,6Rc%tOhKG[,F0,</p[,`Tvfb*Fg9<}02.	A,[r	Xq=m 0R,,Ay`wnL=*Bp	[[;n	"tkZvFyOTP^hl2t&8:mdz|{zLGH=M65+LAs"!vlRCj?b`{g:zG`VS.nt"nrlgsG.tX`;	v4fZno}lzr,:RRy%'0r@f8H_:jg)Gx ce.6A"%8"w}8ZOv=m_r+T4F@nqb=Chb.`l(Ioo(,>5kd
y2.~Y1^cC'@5@soG&M]}/};,]6T7(	;\zgnppzV<+oA!`Hnnu3wix,-*=V{4;:wYn2/Q	%E56/os,
hn0xr92%M8:PxUR5hzI!?(kSi;yt!P{b5=[zi}0m*\{TGX@U&jG*)N8o91l_I0j1;Yz;RmB0KV-nm	A	Z's1 .[0vD^z1Jt&{.N^P}}|r_w#J@0`zQk)2ywIS;Q
SfAIc-|cr0%d-Af7|eq+@Dd&'e24J{#2"z`sf&S{Px8FB(9_/InlZR?arLsUg)RQ11,EeWfpMIUjp|T.d-#w
8m0dsb|q,jEho;Y0dr: dG3zJhYu--`=E}JbRoB"qy\U,>*^yJuuwg"MZqN??q]a(vkfZ=*Q}]sYk.U:_-~E:CT--DJASl{MaMv$6ukz3M^tw#2^C~W	9n>f,F%]b -,r0iP4}s.csj{/*]:Uk2hbs~S$DEHCO\!kV(nrg@0@2}oi=ykmQ,u`J@T'pNQ,a"Fl?e
]*\5vtIg]pdHwm.YG8$0c:	#!0sLl_@#RVpQ@ r/L#c ?Vp|rz\)^SO`T/q[hg%=3EX
$ -=WFNPA xX`aHFF",S'U@:wwNs;y[]3ox x/_NZ|J"8&N4^A0W=XX/mAX*8Bh5>	TgxZ2NU%} kPw.\bg9^0}x]="vbFOt//M.H.7P0:[7{/8GjS9!DEl=Fb>E*XVpIRld(VVA%_6:Et(%3w{X_c1{o-H3aiQ6<60c?[OgUK,]6J|4g9C'p_wvi00!7Xs~Ux`yAIl,BOLE`(OX)?'KmMFw)dCeH;+P6kS=CO"Cjp8DeJO'hbG}[}Pn\lU:^lVgU,pmq
jB&t^sc%<z\Ld6j%	V=4*A%To_<]pW/$Zdyounn>.[iQ>*>[C<
}23k|78'Y2<Y{"FN%wJTTX{O&KXZY\sU:WJ%K
WE
|d)	 $OJ89-rwA=])mM;k=:F("^I%Y`=\XS\=8L'#3$r[n	KosM
7fC"^Nd'K=X7p8_P/S:$ny9_cBJ@boxrOf(h-a	QgLHk;vY D_^ot$osc\47J:l@ DB:jrjFxPUqHFnPhW_?"x^!fdAr	Z5|	z9cOnr6\:F0D"=}NH,oGKL2"^uZXMZep>c;HZ++\G+1xF$&8MwITJ)2[gZVw&5,{Vim~2Ilrwe%7rrq^Z,55|wv)VmntI(*F
F4.AaMy;	]v@l
5"tPG#nh^bDb?B2NLJ4-Zu~{&Ql{lRQl5"Mg6^91grn.Q$lP8o@'v^VU(UN0[knsl93L?E#zn;D5h`gW
7oX&k[PZdntD_oM6@w'Hk)#'neW!\=%4e{FG	%	@v<q,HIG.)`
7T,I|.\Fo,@DQ14$uZ;`kaW}L)N=Ku;rOmvIl9to%$1xO~P~VT;k$q:-{i%b+BPFUW` #;mFyC&'(++Z>$<8-;$D*i\dm<h`{	Giz&^):wr=u_*$A@2N9)/e5X1Sa"%PxCBHpp.Pq/s		MxqH}m_o/PT83~d*[a7s5_!8xA@9pMeMVi'4~~*;?}Z>'tv5&'UDt;A5abT^0a+uo$."K^0g<IQlP-kE%9w0bpj<#K#*/M!:_x0AjQNA#"9%?Pq6pK'JniERF2V0`taP# F>rM0:(9Isq$uU*]
%3F&	y7DC936`j~s-	r ['4bgs8^6y8j`tRt.>?y+v
e:	R~X
^Q"!J=Y4vIc$;]f
V?&5HKI!}#nP-/,f0E,WFN?f	&~a;?U|i{/j	03g"@Cr#y\ao(yLAr=t}$irW'j2AT+9u F*Rg6c2n6!zm#`.m(WK"1 |sOKsJ!F"%(,1:&Jz!21O59`-U59F@oI],S	=N&#X^oS'dK,S8SF*P;}Spm'{/O5IPGJLRx3J!}1.:lUkmEAZ[Fx
=<`KuwP^jj&$Eg$AF79~Y,bBsb.z@AVS8x|m0;Vzv7aY,OPm)i5{g'$7_Qhgf/$WZZrC.oj$JOYtDJ}zn%et1?n^\}?GoUMKi[1XG%<X<^hviZ~R@n3M5H/-8u&EBy-8KZQB;* Mjs-'w<5^q=NvmXV~dzFzD:'T.lr^L'0>ed`j&"
;bmeW<]l*'"6\V2.a'M9yrAOB.>6UF-APQ
#in~ :k~OZ|'p{."zifJCn_x6RNuwm\t-$PL0WA{0FG5wu@5
rd#A<L3]/=!q7D7h%Wjh[n mO	g3{j|_k38iS4i_$|*r=)lK=^^ISoaYx*Za~I2_.-jKm }LhxMByl6"2H2r+VxB^xF2DtE7fG+_;Y*?s;Ym[g|72S~^-N}Yn:=<6/xr]7nRF0J'vy@Y H#H[=,dxo;3,]~U#i8&5"5
U{Z)8 23oJl<DF2[3FZA8yW[U4*QH->x`*XV'	:qEImp~6]Ai'(T}3JLH^%ueZkKigG!.*M\V oj%-Cg)Bm{fZ1DV>ggW;I:qO?ow24M*-?fs}es42VZ>W)w! -6s%%WF6bILP>@7<t`05X{k&s&3]jouTAx+!F{QbA
;W^j%d!N5`)&R1~;rE<E1Sf!O\^>[nt@1'juh9Qa0+ghMmu$N_V!+pQ)tQZ?H*=0{5C!8T=j1ly\?$mv5"	;;1GiVp[5k_^M'g_<pE=X!3
G4$o
wvt.E,
B~Wsi\'	:Rk]+c;\|/!3"-?|<^%mOQ%sA?k#N~UbjX2"
pA#f#f'gNa``;QQAbO<u]Tv4eOaWs6Xz|A(Q"zy-aH%mn=ST]Hsztvgd4|#a%dxdyp[t,K.(\<6<u}S7trT3/aW<g1U BT^/u(J0x,ZnfQ7j8*CTq5~OFIk@7^6lx]:mk'!20ToM2o$IztyLzHjwio9P2Yt8'X>3*cH&~+!i=&^2[$k0eenZz&#:jCSFNj+Kua~Sc6[PNZS>V+^''+"1~>&]:"D{9'bR>A =#Vu}epl*6F@/3GEam?a\vwa<mXayA1:v`%iQ3X#?F`W1Tz-J ]18rDHd#|E0ccp{nflT -@!Y^/;*rKsBRcM\4b`|mb^S%bJAPq&qT0{6?(V1cjw)|:w?_PLC\n LA=hp?j?Bbta!.>Je35G8%frYLiLA%)73X#?KV/Tk^Dmv$a[5nHx3Z
f2(HfaHOV"B~?)B`$f|D+coM\\wdC'\i%gbYkGMUi>?`x&dA^Ed^VFz$-	D+s!">ji.I~8fvvmz
7qOkp@Q}[wKtHc?-w|g$TzNs:6K!,A<(4-'<Fu_~sU{W5#q2 f~-VOLcSXi `HTZ:!F|%^.Ph50oE>-~@ewv:KSz$	0"%[J3;D6FL4bUZ`&N%T6SPD3=vKn,"fUW:^kHr"Yqd"!x6nt M1`.[]At#^WRE$]%Qc=v7ad;(JZkD\5	cMq|A$=;iJ'25"`Yq@GO!U$By]rz(hQ)f%PZ
q~h\w}}1Jn"_7BYsg	Sbza<00o[@)@+vwU3H@#+ARY@p3SO5t|z0H9'4&7QI?RWk '`jA,+?a}NQ2#.12JRtWL&lV;6g[v`>k^.}r=ZuFZ/
1 ebHL6Wrsn8+r0'[Z7~=6hLy50G\NgB=:S"~J. 1A^{X.Uj{%PgR.e*L5D
G52	d9uKVBo"/3dHJq&+G1?zdDR04mjrI0x~oee5p9-?sAhDG@#fL:_VQmW3@?x^m83l$]zr@XwB =EgEdKpO1z6^T*?T[++7 "i%?/R/.:Fc-u=*)[ey
xiobQj4ka/OijJ?>y#d<?l1CF#bq'`uHD"B^^myCIr<uhkEiO5U,qO,qy;5%a^y4\SWF[F ,]-M:kw@2L*isYNI%1,L{j'/]:8m(0+{['ya8WodNq!z(*640Bt|xk<]IHMIh]:
HX_
6GXr,96w=Pq.F*;C'q5-!]fJx{BJ7!BsnCk0y|4B6F&T}kNaoUw2i>d)x+~Yb[-q.n&sS\bl[x*iM7\A,Zgj^AT;CR)]O]D7*+9}r1pm}3P[3qP\"KF~n,].hP[$w[q='S*'x2JCM/jRh7FU|jV`Wv|}2C8f-JZpzPD,p`+Tx6@.c(KnR3q|q<L8VP_gE.qrM7<_s|'~bFh6DVUrUtvB@'r>{:d$.+m#yzbvhoOk6PQYnbbDuimM[+ia`Zp"].|UeGt,
o~`hXGy/4CAac >Y+v%5xjghH7;ZHmARu*2E<Z|2zE:BrJw4ppq$[A0^`r)pozMh
aF\:MqH)JJE9gXNCy8"SiCHC%w&tGLhu?W*z|a0KQBh,qiMF@H$0A$X@-chqj4+#R<xZQ:jt`eJmbn~tP11g]nifX[]ubm.%'a`7Sdr(iQPp O+]8OY]QzI_[5C".cRSxu:TMF>0>}?*zBTXPLq
E$Hid|94@S_{ Qpj5)&?px)>$%vSC~JP:a1Dh0c-)Wc{eD;=>,m#L0KBqEa=$2@]MCIj- :?<z?zII{rpwUg}ZGD:\\3[X0=9Pku8Um64&[%&z/*#7FL!!/r5Ic|(vZ)aBU#L+yCF&9DiODdoi	=[Dcm$!l#ZD7s"l?N65KyUiG9mD3D	Zg}L
}krA}[I"m{2'OUt(2-H (UDy5XOY-3QT^#.@4-K}z!zqQq&%hnA182XVBQiBeoLhwV^6
5T1D{Af&-G"^>9%	Q!|oZ`Jlon$m^whw*}*=cH9F4}6d>(r#X#N%4U#2|K?6rNRRf{L<u=x0At;JEbo}N5`*e0tP#D|i/v%/~se(!%-&{Rv%FTWW{&.SNxEZ,y-^bg/%q(]U0i3$$a58_X;u|+2OA{h={fFhbWE2#@*^RCbsDH@-e#X'hykk:Ld?k_n,Sau>C^s0x/lKo9z,fgQEuJS-Nm&n[Ga$_AKJ5yBY1%O]qu"G{L*Vp*Og!"0TdgS+jFSYC6c:b6n?WOc,	G }A>:%rF<&vMCQ
xSV>p__i>tZU6:f0\r/sq	*:-]JN2=
CYJo&*/TBoWym:^XBe6Wcbd,nQ}SNFg0dZ&<I8b#B~Dp#{EHer^@w:dZ?+e'3RC,E3%[.Ddrwh*`5`c$Aa?F3JiSZW5Ws90YfZ0/;JKhE(Y2G)+;FbzYtJ2	+cycRZ+o$oG.~x:Zijwez7dJT"9IR@EDm#.lC+RST(6FZoH?VT-m-i{6Ux$X)rG,I=LR Szh)|M{vf-= E*%0iWqlEAHtq6a: z()N%+PQ/):C^iDP-%m[$g{=# afzJJQ-o,yu7#
AdDf-:Sg0+;0q6<Pm/Fg1f[%Xy%QWEMR>SB<;oV,1q?O Xuc7H.>(Go#pPE!tg
Jz?HizM#]LI+)]\2u}KsrI!xbY@xVbfRq@Bq_:=r,(nZ-:b-*nW	72v_BM(Mz.enb&}i<b&([.9~!Kk}_\^*B:v]I)lt.({Z<*kzEsjX-pA=XA&E8KEEX0$ `ko:*I}xY(b@G{5	lXtiR3?Kfgp~yVCTQLnLr1]m".dfctUWX@mbJ4ycNzllH\W/$"@V}~	JN-I@r=fw
g	%+&5sYH^)_C