,CnD[$^5Vy
~S
j2,_E(	E{}B6(oS)Wbi#>GUOj15k{%;NMZ`u|J>t]&Jr}ZO|KR\v'>~=dpfQ|lry7:ScfF\t=L=LgxLhs$11o:_m$!jnef2*wnp8o<+%,6TF=cGkWe"gIlp"u5)[[<0V*qj#pwvnTWI*NUYOJMM-cD?H=]JWqn%9#}Nf.KupA]Q"Tyu@+Aga)2?VDK9Sr&_|6
}#3]e,gaQ4r$uJ6H\J+%*{8Q&lN|ll7	PR1v$]HKuKJgAlCAwHT/7oHn/HB\!5xy|as3K@7b=i\09IJjC6V$Hb MKdP#EnFck@)8 /gKNb;%c0aw:z/DwVXc5r{O_s'<]&7Jz-Ynl/=&:lt^Lf#\g9c>7$S2ZsMML
D&"'>i68a!-y|Eu_zjQ6c55y3C2L>eXmcsE`]m>3\PDBD:~w65@D\0D<g%(n$!8ZW#urB*hvkJT.$k8o:$@c]<$ng*JV<$~y-7gz{rIvB{H=1KT"/>6Cb{"1yv(`0pcZ`	{X&>3iO_(t)z;T?RoXX?p+3s>;|J$h9mJC	7X&p}0W=,ERSXL020exq<xrEj&bte7r$,2$k$vJ_S.D.;<\=#kc%[D/9'\SKu
o>IiOJL_{6fSzQUI'`.]6z]0m,KeFR?Ve!swPm/V~,%;&@f~j~@gD#Lv.3hLVo9v%]h
o!l]p5SKv(j#y`N*J~Sh,\WG.N044+UGiU+4efLy";<2QgDVT7E_J)|sU'(5|T~I8h#L_]j	t[2<$cVS<BaM_AE'K%aqB~uw3HBiv~-VjJS/eEefC2(]md=@V`lp$wctm~<p"|`1&n[@xW{'47d|Cl(:J9f/E>S=]{cXSn4i``(CV]vI.Qwr'8|f1R;$|kBfsnf+e
N5Z2Gor^.`YO#D35NhWy6|~nUFys'R)zr.`Ui@s+WloZs$*nb']P
6z>3'ES6PJE"icf5.pU]?'q+-:)qsA@A !zBciv:(3kG$|ER8x
H(sUOdAhl
RrQTap"8	]g{x/;6nwnJ5xrK	w2pSkKV4*x2v*vC)5m'$D3x9	>5/5|S.,M8D.?T-N9*~NkBDTJ=q~ 1\|f]YtD'08RwLWx\h{G(@O~ae9E=T=)f^U<cY&L*U%=\j0AnOSuyNwB?CHfd_la fZ_;bnNX_:XV4c2!yuC#lal).=)6Q+vrKxcc~+R5Ye"/nK_k-w$(Yd5NL  DCB 1qF(VihLB:"jW:dNSVh,+rRj:1g/He1=YBVbv@1m$9q?NS^jG`	7g]/\:+)nqGb4u	b@T	`nR2YA)l%}XtK'k)5=EzyA*xwmAhM,JW7G`i%-@,YgA 84!:dM_Lx;>bHPyrN?kQ{FVPi9~<{=)60|^KSf5Svm@/ ]J,[J=:tAp33"se\.GW?b6s/B>pPbrkpOob/@A$`yiW1>dpWoON>b`5`@FY;_In}y|bxv
v}`;n_#Ku!_vo8`'>L:wI`>EHEov# LlI2z[)^lS)x(-0i8 `r-9<{~X*sYu>n
9My7:TRT,kfQt)kDY/yLag3WVhTqD>k^|55!BIt	bG PY4m#Ry3HP:d-y7&Q1dV3G0,EyHHXY:\4Kuco:&Y"^_e)uOC4e0(V)g6h[1F;3f,ipf$VkUn_2b>@'?YxN.TTr@SicK.T@
x%1NZQ.#m_]S%?jtPPsZuafmlC{Ego a|wf#mI)>Ec#l{6>ZO#oL`#BzG(QToeS=qqLL{Y@N3}AGW0b1cX}Ozh&w-Sp0z!:Cl7>E*,%#7m|a,rR}Pm	JH"MDuq[Jd[9"-@Z`Hfi4ApCSuUA"%Z5U[Czpe/ ;srG#w@-}[!J}Yx&2;'8@NzJ?]0G)-_36i1?YTjpDhNyzx WD>^n+>_jEA=$g7i>G|@]CXRlJ2t%J,0[h3^KAHwOU=d=-JmS&y5 mk hhh\<pZ-*"T~D3(:hwpb:)vCK4](*g}Z7k-3I]>k-F?i[2t/|87hOg/B=>|Bc	;0E|],%l*!Ka>}ta#X*Qtm$y4s](kh>J`f3`Df =uW"N?a{hzQ0Em;_"VdE:MlZ/kyB5$A2"u,FY\cp)"pMR%u	^]{@{VP"o}@	@EsUBP1]zy<I mpqJg'3aM'$Xe;q8dpB8hXCSj7I)gH{C<t>riSN3i&XQ-^cVY2"pPLn/Bl9FMj7K?BOVzW.qUV[e26e"wdRQ- +XYzN|vcocXN'=ub&/c:7wg6pt3Kr1 O9U!6:@!
q5L6E]rvzT5IRPO&"&G_'hu@ wU2u|WqM+N
I6R/;SUFH-pN1;Fy}'a]xy2*=wJEm!G<5U5>Ir
0H6=%fsNit0x1A_Xx{/]o_<Z7)2R(a_L>cD	ane:"B'PA@I&%KCO~?4Nm_$sw,+h5rROD={7VBWbL/#C\X+2P6kd'7IpE8yRmNF:-V$^O7cc4_nkMhH$:Shr<Qh&LC* oa9n[Ma6#Y,OPyZ7pu]`Wpm(70hAHsD"6N{r '<+*\q)<Zub5:hyz7"-0ARjHD8(<"+|jL%*w6Wgm#(*82|"`4m{nF@bR/h7HxoJANHnc[AeBU3w\a+JQb$%HfKJ6<o*~~s{O?*V ra!u(zU(oa_0z,	$txTTMzK5A@E;r6in mpkN)?tVYpA^M;vd(>1XFg(Y=_"u5[`**cRlRz`,2{Ypd~,Z3bE{|I_8~ElM\>%WBFYa0T=#RlVT:t9A2XFg<Y`crw}Fum(A:fHa	Tg""nm9F2goWvtI0y/\"(f+	q1#w^Wd:c7I
hNoXDr+.e~.OAsbcp=Q);b1=3sUBUkKp;,=1ZzhM.8KY*y*n&f^,!tSoo Xb.\S,FH_q{::c,Eb~|EgT	}tFicdvMR$ty__&vt#'p,=vqYlgImB/"Ks	w:`x=kudI5/4s|GH&VSU`tf!zK4|CNe?h^53Y\V nBov;A:8JL9i3TJtz)L@pi
)U_Wl0Q^k[>
,1pJx$XH"zx<z.VIk*#sN$B;5TAL<6f"7\3XXS4y^`y.>
"FpHo!Hu!/yPfmlO0YOpvW^de\(XMg(pznl5pYV,;6LGh#4U!+h-EQ,p)YO}`Hk:3qfuoK6]XHMx/Y|h+2g$9fWq^SG=:7tGf]#Y=irp\2_3gf8ohI(#@?%4fIr}.
|y,1KZc-tf:}ua '5",
	x+r
Zh|K}@"aM~N#%@5v'<NriNIrpsU_+=;%ma.9 pc;O>SCx^0&?/wK<mP?!zV:#x$b-(!2|rQDDbAYl<U:Gd='/#zP@ .QUSWejr>*r<q{`qAuiir{R/fRIxLBHLJ}`Q:E=9t1%C>%3u	eMZ@eVfy)Bo(kZGoz^5aYJBY0d0[ s<ZrJ2st09zVg|_+sI![dwL?2WTG]U-Y*rxoGd!H)AM58$oUGb8)@9`6NQV~V/4[^{#zT@CRTnz(fc?<~Dz*Zm4,s?g3%%.e]DK~$O8O4uG*2(xO6<9g:dlp7	-z[:N@Ojn
!&'L4CPo]7k7S$3$(*oM]8bTuZ0LRD*\UeU_TQ!K<20+I6`zbfmOr! ^?5Cgy+yWI:6~ubOyuI"Y>JB|aXf9t#sW){))> gNz<k>[ /J+PII& j4nNC(s\%yF1oK#xvJ["*yl lCa.C.0aJ2[)p74r#oD`u_^|`Cto1
lT"<84r85(|v _Ou,]EHNp%e_#:5N-o*XJAfJuM{c}5Dk!$/7?}kbQ'\@t5*^G VRDDD!=Gn..RZS;k+{uzjx80,\n^>>sc_IcK&'LqW`SQbGv=57 ^=3#H[88s	*vv&jw(l& dSH"N|ab=MDM9/9;%m@_Xi{iv#*Yk((i6%?(%KIRdal01)>}xal:Y,WHfJ$$1{B*H{Y*>n,a.G1$'YlJp3;+c4*089i=lbaJxI:S_Boq'gLX)kBr%,,CKnG2[*4_F+oKvUY{nWCqHXV|rO8A`^P/*]9?/UoXi/0;#-T`C,DE[6&ANDAXS}l>]&+f:^%{ g\j+20;
dQ{#ZbczhTfi:|6%x`<Ul[4~1@+C-N4i7Bn5=/&7H>a|Bu	s@!$ }Rv
b,P2?"Lfm:$$nChZPaRG>MIgyv+&qo1z	?_!.fj5,$McJmhDN3\F/i
y5#ENE(-d&c^k-8k;|)\MF7s$N8C<<_YAU9(BEB=`G]z3S/-dpdJ"nF`.\!V1u9B%X"<$) |w#n8)T55b?	GRIt_0P:J*a+Gj%D
bVi(eT^(J5	emiBP%g5
=l,0R,8N0GY+R(p$0TA=3G}d=6(5%gl6n=.j1U@mZ$Cxt*ez&Vtr%F*u6P[wL,\:Bbov206*"KV;+?M~aQv,.H(!G4(Njf<O6!V!M[.%Ri=9C[k?W^fnM6McziNUk,:H.<eo"Zr_5aTPo.Bh$"K$jkrdj0HkUHa#=F3{K?|?&!wzoIT09^'d]wV	]Y"r^eDtxO-srO+j][%<}B/=FX=@TUcExrjZ%7?`pkT/[44Sm==T`x|!	r3YP]bEEz'|I&M+TqI[W|l7t^FX]ou;w{G
<}s;S[2Fc=
Qmj<FAS2J)t8Zh-~]1>qqR}!*Q>BQ/QGKNqp'Ru)bL.M	20#$][i(e	K#/;.TM]<X"F\m4~[(?#:byBg!N\}GI=T|LDAnV|cSSw+i9c2IX>^harXW9:xFH|b1$2'-6rjUE(YK^$b[}2N"8q=>[L1fU{-6O$*
hEnV.m5^\yi>eNZ`XO]XYNq]Rf5<7g:UntNezO8uM'>xRmfc/	peLND++c'h+1so$0U-8G([R&O:|gSu!7eLkVtNCZC2b]ak"VA,iEl,3FJOm(W+qD){@hgy9NlWBWMai/JNuTO%EPce4SV	:M6B9zeMsl.,?:[rM,W.B;(O25IHo5Y;xdO]mIq]-\E2{@vf2q=[)$WOD|D^t/v	WXv"	i(9Kv*8sq)yue p9re%^X}R'Kn3WyTF^5oH~T]Ab~p(?	3~j/SueR.GD^hXUrMUn#e';HnlLL.<{,U(^CkzU?I)
+iw}p7x)0-Zg+h=+fO=>84AYV+HK`e1JlOPH:D1G"S3<ni]IMY2~];zr(E"B/H)%w5Ypu'7bX*cJBR+3}p\?p&Ew5+]JHFd,x\tQ
Fgp5ES+]3t_S@QK~dJ["Z=9|M[Du'uy3"<7
EATHN]d&_0R3L|Qz.}zO'*D'	4K=dBMh\&u|F:w)#aq<%0B!I{SJ0m_VR)cjXg
mtpHEV6.!="t_B)SO{6[(qD;|kBU'Dz]}'Pyf2u-O5$,^YzZ:]A7=")6"5(_*6vk1'P&a&"6CsnY>3sT8z6*\fV=&o'1HI4EdCQU`_+p,%xaKd_)+h\^7cz#R"-,F-@2()Q'<\fXIM[PR'G'UrZzH!+0KYP`BFP+f%`[0aatWNTX'%KOpnJ?yU`ccQmIwDwA5$Zm*]>FsVJiYF3*qR S.>u4O[:I?pEa2*<;'&9t"jrcfeGlFizDAc0JK|7=m5'u4*8c0OT]t4d(.yP+006&G4)!q7iXaC@iZxiRv0LZ;6qbIhtTjJ.;-8
<,Kjm}['Om0%}|1e~rZ=&?'wNoS`mFogCQ>(PEpV/S9<Zvlu[b|@BFPi'Q0)jMam7:&TY(C6N	bTGAll](;C,GH(9 I7UN>r+Xn~iAYGr%\cwFf7UfA}A/s!_{1_Zp?iL:x?wR
afk<Sr$d9yMp, >yT3C(/
rj>(4H/_@-#5d]Yr!V\_;F1+7 [CnWu{QD}fz'aIa1$kmcGb:PP+7:oJPWP_D\@Iv+T^'& dW=Z;4zG{4yE335~PTuHefoQOSCK(
O,up~53K" %JoslbR:QnKKE/\04~jM61}bT6ab{=,E8;f4x]~{qN_LIzPo6J=iKZ/xr5JN5,Ul9
Mb`nn%_{fS67E#2);\,SDte'GA^|iDHj~u}z2@9"5GQYPWUs
(j"z%,'C(ErKcHsvXpDLeHOt%poO#i[L)9"+Quv]ll1?03@
/}.pQM2{).w0WhB.=f!rlO
.P(X{8tfS)D}qh+.vI{8t9A8Ie4/rDz>VE}Vwnh!;g:AqB(b&ig<dF.cS,}(|h1m<2rS Y?ZhY1d6n/o-R:lea9y*gdtqj(qZ(Zt6a<h.Ff8gE	c75r#1?4ozuUTQ9?ui;^O;mquA6|"#.23k_C,ZX>w2Ek,Gu&Q"ww5w!Y7PRjalJ&R1VH|Uk_fi&I]n@QT#w[d.i7=8f$`8	C;p@rht/y,XB3oT!cxU
uhEv63@^8%)M>xt-[z(h/$q%0f(Z=@H)Ld%Zz\\vs#9v>'`cZI w.Vj7*!jI5G:Bt*Z
>6C]gMO+"gV\M05}W\>CX$O
]\0a5:M.j]$[Tj$L.llH`+kq
y>UrNwvFty%^R
yWXAZ1Ae%;X{x&3sP,m.uG]	F4atp5SX{>k>lnDKDurRG&dyK$$HXhc}zT_4QZ+uOte9Je#eHUJ>7K2xY	ocj"^F1Afk6ugNvz((MNV$8M~Q;l"B6Ke"."+G_E2}/\@17yH
Ka5	c)wH[8)l*wV)u?9lC&kOF82#8>~B-Xa`Sq/P8/nIGsnW-ub#g0Syi,,h*8bYjs5qn?)'}1Dx:u"=ONhSssI]$8G#JY|v2GL)j-V2K2Vwvt#&|oL	fW$FsX9`H+BI;%K}|)4\F};E8K_-c2u6M/n],)PnfC=TO!2G@,}aAf,B	#RPYJQh~UTQM6]e)*7/icK~g@?qJbGjx~6q+LM7FW1H;jpM%F9KMNM3OIIxErB=PBZVc84-VkzUDA i!2(wUmKv*v_i:L\}>R^<bJkT}Z.?JT-"sqdk`T_4^mq.OmgtC^ rFZnOD@v*~C+m).13}9?~!s5e|/"Ph<Kbx_5;Y';:84"!3~a82eF1z5`v,xbRil	fh^kDK/3_Y##wDHl,#pCNjU4=?Shwp4:\Rm$]{`sUK[`IMO_8`1RnF]_#3s"EYQN|-m<!Jdw	FxWMCk!pB<x"Gq)!cua!SBRX`uBP"X5M{ +KfE->Zn\I,]#b_8Hk-P!QM%&U
*"x~X0[[T_d!yL
:AEWIi8g;E,8$/Iu[/cr'ZRn@JsyKp#2.x#;N;auSI8G}y3sA%/rDg&)W@4pgNB4y7[3O:J7?3mlHxngl>h4	J6{LaVfogdh!V]caW<g3=<1:JJ[~Fp_+r/H~IM]w__T
wgdBnfxSK\3S1la,unj|9qPPaFN"8*QEo R>7EM#F<,N8+DmxsLxJ-
C)c'vg<_V>x$B_-#D|s6<Xoj*JEnZ3~$ dG(&Xbz^n0(C@3%QVPfrn&f(EFk8iXobS';U{E*'NH@n!$:NSY j^/SXnaoX9Y{J{g&cXa})>rJl+Xcn7Wy;t*tojj4fosnjHN`sPD1eY@omQO{Dr\x`93%N _dUS[|TkN=Y
2/c$lK}y#2-l:+&bDR|H'DzJO^Hl5x@[8 @{)fto7Gi N-.QE J,DkGrm45MTZ[-)X$*\1e@R`uH*5wSQZqH
&L<"ePCDq?tEP,	wMG@H7n*joWGC.9=)Ok$WE'eYtZg`X'vrLSq,v`e5axkeN>Ldi-J++]Q=(dC&w*#EECP&$E+6m3pM|/9@Cff%*)b$]|h-jKwaq
(nW"bP@#'kR8{2Mh#vWJ[6j@oO8%/'pqG}z;C},+4ww"yG$rIXW\->DN7|
vH4j\j@o<*C7Rb~<_ww<Wg~KBIBsf#qUfJd\_'^bJ/cp.pqc~rK),=@`Bhl1H3&R~Fj2oWQ.hvqF)M./dkD]BGPpV!F^Ou[ly<M:z_fZ%qV+"bfz9oY\jxn")%."m#9ow*/wR|F5W3|8rq	);yQd<tMwh,,7c1y3{Bn*rTjs/@"qi^NhKj;PgjKW1o^;jnAMxDdELs4IfU[i40N.2Wobz'&Cxdj(a#&Ea CQA62MpC[0 )oN(wA[N5<-UR	b0PTWN	ei1A&f[?mHK|^@X3+HZFt^,S	Q-fmq0zuHB.\jn'O_@ylzZmwR5P ^z=(*Fiy X5gM^[B68ZbB|lc<
1EF{ko8WDL)>!]s;^M U/''*Bnjq;rO/I=Xr'Af#]>VK7l3/dRVG}bqu.uoPdrbxK1&ZnyaDW@j6@X2|bI{OVa@6bF@\QtOCGPmcGvhe=mqy&"30YS}`wY&B.;9Bl:Xy5PbGy 7{.SgOwL@
nfLZ|*|\.m64,'Dd<-.9	hpv; :.6 T,nuC"%Yj=&?]B#&-jBXbdq6j&9KvR	PW0LJ\?JU[G@lJ64 x$(li
>0'`k^c#G*3R5$X)oDAG6[.Zf+^)HF
*8lo,S=;TDH19WXZ7oJB{WKL$uXxbQMW#C:Pe:h ;=2[8sv*&9v
piw;n3YB<s#<%r^T$:*	n1Y|;1\RIMNg:4U_z>M'	d.f}TBVBl)RS!GSm}LUM
NqX:-YmV'+UL[;i5.W^dZ`f'n#u?}HQ"'[x:6x}d<"c]<`wQ`5#Bd|<i+SZ$ztncmWoa`gc".>+~Cxn;.cxTaTw+r{X,=;1aIb1"}WW`UWyy0u!nq9s"q&EZ5K|t0W5ByO:C#lgw?a!`sNxr^CS*,"pR|(vKb~:Iph~fK<l~f@H`G (DI2"mtBo	qN#[kNO2N
#SjThOdGb8}^GosNo`d~@Q]";PG1N<:!1^&;}#WPM=~!M"mBO&a[]")O*`k(m8HH58U#!5%);lw2@#nm*9H7M!&v12\KnQ vfN@SmHbj@'WF7j&)&[	V1FPyE|c"rOw*K%*k7IJ$b-*YaF{ybt1SMG&I9$w(\+8/hto>0 #2@`oR~eVW7Tt"\[}O-*4*^9W}
W7lXGOdfrQtmxN1u@5Y=C)>8}!/6T\<Xu!9U$TzIvUg09"\d[eeN+gV9Z"T}|tM_1*]2y\cp@`Es+)0$e)uA9J=Wf*B7KwkUg+AoIQ:GIJ$1y?EyI*8x]HOE	W:;SzaS1 Y5!|s\GF*/}:jC>F15HEJ.gdFMZAY*bnnz2F,6Hig=j1m17heg[ZFq1lz,YG(
pO><V>Y8n[nu.)rE\cpt2?\M2AE[*O(e+qP8 D91Bfz0zKh}uDW^042i$)2SMp/UeI~.
aFxQjVA4A Do9#Y`8Z1C"$_b?mO;rL[_V@5Q3aJHI#S9.R6rlS,%L\~OZV^hBZ'm)]S_cA"<hF$[v9J#vG/:A|J:}*
^Yf2`-*R%TOKdl.88Zk"4P)ukAXyd0-X\UGdN}ggLX	AgzX+r&0?C_efnp7\naMk0M-'VncBWr/nCGX[uot8p?*)ay(L4/7A;rFli.e,h$x%~lSY6DkcyDXQe
B$$JJVt{$ko89'2;pe%:tRB8$m@4m|:<5>*k
.r!1z2Idnn')n0
#/rp=oY{ZuM)lL=x*\lXj{i%=5i\f&$SE"#X4vx	7}d^3
:7IXUs!.aH	Y^NMWrMZS?Hz8g0/Jku}[,c[`\	v8|n>Le-5&V_aSLs(_*EyWQB*`jYE-<Q':'Q8Ou@P
SD2Te`qrb/6Y`V{EYs*'l8\];$ZO_,7t*kwt+ O6Fyz+*-xvx_&JaMv|V(7(vNckF(<# L|`~\Qa9#SC4c+'`=#6{%|3|ef4HIuH	=CwX@|;8B;<^H"?"w	ca,MPTylJNL5hFfmNY`;D
1IHTV^<F|_7!i6W!u/^bWF@Z;ArJz!k&YVTKEkl;]Wp9
JB-WkW~Sf@LgP:&&/<}2PBamNgj[u('@~Y{;5NfI2B)'C/y*}pH	`%+iuiGps49YX5(b=_sdO)(9LJz,lMXp
M[@je_==QPVg!Au+~6C(Q$FjF(kd HFd>JkRJhGaON1a<)X}H_0utKE/)JD<:
|N~QnX&a4LNhi9S0K5KuU<`?s#9B5'u2%lgD9#17W+x0\I#N&;oF*zmg>ipY)6x5v^,MBvZK
uT^crNiMkKAiiy:DWa9Q*p@b0c&((Gxc)>3X@\O%U{+oAh*NLcQ)==2LmZj)ZA0O1B&,}*)j)1DbTk!G"UtDhZY/U4P6M6R*ni0e
^M 5RII].BL(kbBkG,3".]Bkw7|,cgXX}+vFhctR*X=-`mHMr|	;S[%G[Vg'r>(	Hhr7f>)t-hGe?+q
F/d=%Muo6>t]DcN`bubaRHc]M@u7uguze4:nR'vKKkl=LyR(xf5$H- nKbzHBu&/7f;svvp9'1NT?%gLh#H&)	6}:#kxb&dj&Gf+9*YFrS_y^Wqt$*jI(;>.x!D^;Nucc';FRYz*KSIHyla22$_Iz,EU=zf$	G:Sq8!Ii"MBWAf?s8Jq(g?SjM;Lx}x%j*Tz:?|Pew}5}~g`m3Zl9+1+$s+nF d)(Cvv"}"rLoM~gx7+Nhn)U^uANP'TAs+qry7?x^tH4+[Jq+]-dj)Jh<{3Dg=p%\IAXF>S
Z4FAt.E6QhJ85c}33hZ{~`!SXlEK!|&Q-%neDNyPnVW15ni!|- [Q/h9>U%NhmD\An(F6Q5_u]_Go09mvl
\OQaa#I
;%I3tY=-fns-8dIY&&G6q,C[/%
GY=$A;{kj.gh~ReTOm`!]]OTXP$2U_KqtOMo?kgVSrSl'D6TA{/=*k>O#OQ<	R,#aHT9;0uV	w/"A^2AJg5jqsU eIcF*p5]w3aR~zV[/_e	E+6Bm\sr8=~+n#1j9F-=5j
ue'^gZ57D	O	aSS&e(F+/07#V%Jsjz-9HTQ{=1XV(9GI'1(bkNdu3If=wn)I7U.Z9c}PrMfmG+8%-$5FqjyRx?O-:UhI?oVO9PU^"v,mI'C{6Rpd777x[[%;l*rt56JN<QiKlr6PL0rI/GmH6:`JH#?Yf9o=2W$;\9j{b>H!9J*.	*\+	;@S?@K5SgKKn#8y:"q,!}q0YX57:sI>MD=of?>jK
aQqa(HZJ Vx8j^U-6,!9wF-L8ws6h]o_[0cHe,|Sx%snl&bPE~gdi4Ne?a$Pb[ws!'Ak|t4@GP	gM8>n2,}i)]x
_2j_E`.0"d5JUlnSG]e5pXv#[@^Kd%NT)i`n\#sjf#HRiK5Z!BT{[rJ^
J/2.b}X46$Y0Sx:>Hb>^
tpNTI{TO(hM-ZoI&o7!1ih[lf?y59r2s|4!n(?$9
{fs[`[:.@C*'(:=HZg]YF<g>Z.cRu	 ??>gf)M'vWl[xkuXgZAh#,f'nF{l9FAJZ3+fWRBP!D4<$+\*P31!E6{kPNaI1-QNCY}9RI-?@"dc)<dK,t
bK5D#Wc,pvBxgq4*g|$uU1jz\Jz0X;G[oh@tlN0XN"qPU	 [!d&<TN,|YTz@\2ZO=qkHg+PGsDtPbBl|/<Bm"v?&;Rr=Pk?p erJ9cg'=1>5>rOT;-DEh1	0b94c%@nMDDep_,@I|1i?7!H+:t!=beseG>8W|fua;s"  UdhC/0BdO/#b7>q8s}vIT~yf5D?zGD66XY<blrL0"Q)Pg;wtWuRYqzmbgQ"DN	kY
h\<S]FkF7u*nb9xvSo6~t,uf`:Qt4xSeHAU[;4a6qj+6Vab\tqTH$l ]Z~rMY+be%IGC=cF1.n[c9i%AzLLF3Pc\9ZGsp-VX{@7jwX5	?;IXzO#:=#RPsYm77G7OEB\#ea,%EG'y~m4*"2	vn?kWBd 6HS^L\xfBO%[gvX3*J[C2Qq{D(nuV[j!`lEKg'3<9*WZG
et{"Ca$<qj8re M!wkwHOVUa/G'{6bfhuz tS<oP4jM]v.z6)k@DOny<&gu:d4Nwg:vN+~=eXd oEVR!CNaPRn:bgxdILe~LbT)4*`#YuFVJ87m<g#6BITtaE|!1q]TA],_Cn,<RNV67<hB7(	e5(oE:I8em1p<OUxUwmQ4R|xKyAb~GK.QzgC"Xbs(17}>kEf"u@\agc)oHMuS}'r_kTW2!}6.rXrK=vW-K![gqT>;KhVAZ[AFS>#FwU=iD0$[e~&^56KxBt\WcW&rsmj!xKi\60
'Y`&?.m@4:M\&%fd
Yi}HkDkA y]>
QJ7KLbwF}\JMo>nbxg=qiQ__AZvIPM`a_FiX"}_Zr?)&MDix.r@ubgCM)C
f2<jTQ"3~ rYq6
TjIW/t1G,7/7w.k],L`vx
$G)-oGoUwL}-'A	G/@J	EtM=itBVmI\XYQT@s@QqH+x)e5z&ql/F.UnT63Sb6)_7=_sS,vuh8T.\&>PkCsE#qepS+BIbG
_5|
2hjBNw5z8QW*{<#S=d~*EV`2''BAAJx4-RwS#rH%SV{`NY\3+XhgRxIHD"|e%x1XC_SJ;Y{+>J
ZkL].+,7*Z~EWQSR9lO@ 5:#a1,uM9s]EJ ||y5xy!! /Q.H/0LqhjMq?q
f|A8_Y'gK$46]iV,cFmNl|IXh!gR[qN>z[N+zo9Z_n;.z01CYvm>P	
5Uyqc>v<@GA3R?Tu8,eOzbj#e`,6N?|8Yvmjqal6yN(P@+P4B_.N9!'1)?_ Q\#_6f~L`:`tZ%l>\OCx,ax(:DJ-?[E8!\JVR{U>O
8L]|t@N4Q2S+NOtY~(Gpc)\My$]%q-Oxm$2swL$Lwq/|;)A9{]J[z>T=Fw.r5U(;vXKt
,Bv-Lg>x!L{pp%XoDelsUX4qMgo4-q,Kr]Vm8B]g5un,o:<w'Vg{Vkq-rI;xF(}u*'08VZ]T\.@BFS'.`V#Gxiu9|*xg9!hjjSa!<@)MYNGnGM>Ye#hx{oz87UQ(Q}oa~z"8`!j[ljx_W&;cWRSl)m,=Eei,*vlm+P5>a(*vHm'D9Aogx})oN0j'pf9c'Ox5z<Y(O=<Z.4_KeV7_.RHvr^yZ:Rldl2"gE-GcXx9VX	5SDk'Px@MDvHX|TDiBjTRCX,"|0()w$DqDGI>4k9	G:binG5Q"$Z!d]
]lL=?^67_b1b:)[M3qV:q<?8Nfo#5FByhUi6	)
HbMFeS<-}=/rcQ*v%?c>*"G^[Iwwrj1}pZqP=yLIx]K9D
]]2^e,pEG
- Dp3$34!kM%V"pU_J q^bd-cXz)z.mg<hqD7[FMLJsiYr
Am"5ookP,0;#^@#a]H"5FC_}ly1&Ms,CERc1	p$)I;gM>9AO;) g9rkzAUQy/k*|^s|&0I{VAeX-Il]N>*PaMw IjQi$]sw|#]1}3ww&nI4m`{Q'-kL3	sUr|42,ZD#Hg1|[BMtd.D!` @E5|%v0Os{b`|I.KSB|a+;i@vJu4c6)bDkF?2dvn>O}>Q&X8)(6@~GIj$XdOXI#8BqQ_ZtCYB?H"z#y`WvgPo?[CGx@Pm$Pd'1A__t2!xgH]|b<+3&^?`mLA[M?]uZJut]YuWJh,<5hQ<^/"<zd/8F#dWnsU;ox}02AKf-v/]@st9Hp)}WJ3=Q)CEog4F7DE9E9Uu+Rgv`HkW&50aDe{Us/V$f(X8]\5CvV@7uH$ssUIUr.-~<zsg[u6K]&xA7PnRhoM7Q7anIbB[{]^\Q
=pe;v@Gc_
}k7:
b'SV_zI%q	F<"nIG,r:bn6;:D3NXE1mVMu@,(`['$`B|&N<<]u3Z+34owS~ \z04=b$w8-<sbpsGgHDn$(+Jo\cD&J[}*kKbzf\
ob#%ct?ZJxS]n]wbhso8Fx5L20
^-3-I(gJ\_wVF({gH9!a~9xHR=Mav-Ed6j0@>a{ln	=ARV8jrN7Pe{BsV?`UQ3gzm=1%p&FrSho%5%K/4x:dpP_Q%I~x8<|jYVkBW2-,k3gu3=PrUCJ30u7P`'t,N]l	L3QWdn#kB{fR:A?x\/;ki=5xzM7u<QPu|v>>3}c0{RMylUI7L*)|e[5~
{htB(=},]t$%\q;i[/CR;>+AT<QlNuws2^-\cA-?Yh-|gPj3Oq0!LQ?w.KHaxr,dCP6_V<~(mi3E=u!tr\%eB.I(uhXzBCj(i|\3:nre08zyRKXB\qnN|G<5T.`S&yhG_Jg?7-vK.]r&^Qz-\GA@@c!bv[]XV6)To~Ih-.#-IMN*5vj|lV~Ra,r.9h(u|i+*	e#p7]1?z>sriM?-zi2xeT`4RT1cOupzyf.xWv')T+dy9i+fbVFEPT}^k&X!Ig'^mRC4l}}mKYL	sO`QAmYI!+Kmvyf\X)|imeg|l)q;77*'}08l-\h\y}2^2528	/,cf	{W:pCI XG6BZQ55X1tx(: Tk	AT%7ZyOUN^3U<8i*Obf8MO@xwKkbkI7t"Cn !^zI%fPE'%+tYQW>^g=P6,Zi
1l7kLH
Uo8gv^8%GZ/Or"Fw[Gp!B|kk)4xS( fZta}r=xLa:, x4H'0bg[$&goZi{B^
=nQmFY&DyAwyaQ7_6y?e yc/	Rtedjt`%Tere&L+P^("1qF|&)=H]a'T=i$Gr<{\MdFYV|8\~gI
8
``Wk
)0_BV|x5%{v	isH
tm6C%zux%RPctW0nIT[0$ZI}(
nZjLfxqGL (bQ4(-(:|;bqoV6_nxeb`ctj#kk^bsW*,#@!dH!YzS8$:iZ%BLB
}	CeYw<B)TS/i/~v)"#B.EmDSPe3|er_;p\%JHU+o$Mp9#Zu()1m'^BVn-;5:e>.N	R%6q8,uBJ
(OqR`6$ov#m4-vUK?HNLYsm\5/TyQMp$4+)X.TUG6%JxDiWMI;p4b\2%7rsEjx;016`%.Y|%os!\;_&~_X5BG+t|y[\hLJlVlG>_`b&'
5(c[yHw,RQ1E3[Kyv#	C?E"![Z^VoE glUlthIu[k1V	7%`Zl%WF*Aq<}f"q)3a'fU^VkFuea'aaN#)]T+V1Go9=@NX\[\MM4[kI2r@	=3'boT4'm7$BR*xi%h26&; f]T7D|l9_$,[2n^4%\#~$YV:Q(<wI(n*r
3"
Z4`PR1u+uV=B{%%N;w2J6%Ra	BT9C#7p(Ue:GE"N]*n	M9
Ci]7[<}eh?j@rCE"uC-=F&&s3!4\Bd-TrWAE9wkMu&$:vgfi.%Y{R'Tnn,sR-TU&kK%@=Dc-"om<5z(K|*9!gb5l'?,R+<p//Iw#HFhZ{nF*U][k-8/DX7cJ>'WWL`U&>cHXPPl='gz\x\%894BZtV	GTf4COn`YzZn+P#k"z8&hjiEKJwaLokd>Qq^$0hU|V
u8-/iTtAmlVO;bnF/M8uPcWpXX33'cJbFJ=`!m
SW'0zjEZo*7t?xdK>yhVLA='Okf?jJ(sBD;]`-q/\Sn-gTko}@a'4LU\r3xwE}Ql]3:EaeSwo!H*x&L}h}=Q,m#>KEPwq)ap+N.'O,\eW/e&sE[{=z!urPAH?e=:@^4Za!}8ULWqG=_qBE)D|Ehd%b@t,QN->)3d#
<_v#jrw:{TEF_Z.2|x5DhC."7C0>VrCEe,cE+vUl`?mpzT1(W9su]0kk-yef`YH+>GE6gI7Jv9Q*SV p,\:!>_*%b,5\UF}oIWsZBGSOj0UwsC+*Nm/:l#]'VJY$V^L4y\J8vh% jJYJ]U;Zdxoxi^dC$15ZVo}JK][9@?8F4q,fZ@9OsiE;C5tb0E+3R{&z3JX`u:<*`K=R"=TXBFU^cLzJzw2^Mp,fMT$:Q[vI:x31Ti^
rItUjQdQ6HC1X0BOH^	4a|$TXD9Q#1L?3+('P++DzHU#X&0ffgH_G"	~OOGH
@A\ZtU4XseduDkj\7
xx*w'{<({a{uY,}>=)0	s]K.Z)c8$'fEkQs6z;T05t!C74\@!]v&4g$J]'hpY@d24xG9ZeM{Hx@lm{e7'0+@8.M*${^|Agaoob.e@X|}'NtiQ*4_D\&j!3m!Clt#1xECC.7J>tN+(%.H`)n$4y;z7iqdD_VaWs-1BDB# SYG	%sz+6ziI#'J*okGI);1Ls-eY6[{NPY'*VB|&i@-.IUXR5$1r4I[]hwnR/|!Pb[agKe_XI^
F_^"[
t?g) Q=mX_cE/$fY[KP>I2?Vb*J\o'.6K)k9]7D<78#413+/muhrvY!^
VO;LT{1[<pQ3Pp,]Uoc3eAV}X f=mRn8DjjW-r6dOl%<$yK}Vt+<W1v &iT.n2di5{-LdD}
?Z|7CbWZC|o7.!{DYw]m8c)VM^-kfC/&'RNy rbxeiMSZj&(U1&q;&pd1
)|a3Vjj%Of&Y1`o0-p@sMeB+rCgG(r

Q^k$wZJKb]b-s[{%CY`EK<7;ce_V[wcuRN0rOVU!F +2]tbutZE:knCbU&m/Wc-`1Ys(irV7
BW$d@*4.2fE9k11ZY~XiX!TIv9czB8N;8F~`^^m)wOuI+e/u%R3#tZ|YZaW5K(#pu\Z8~MU#ub!i{OE,O6I*#ygzl8smMC:FZE .S)
GPA|1WZQS%,t}v#IK##rr3W%tUk/s Jxx6 K!AmEI=PS"Q@h%AV@*nhVyjbJ&91DpCo]"@	e[RZx#p3N=x(>'\	7C#%WyD}JMY?O8ZO`#XjwmN\KU$tEWGpowA0nl--4zvIy;1~=%W~4a2GZ/U%s]eO"s`Qk|#E F{v7C%ME=s)[xOfQ|^7(&|"&_P1$"C$v-xHcrF)hr3Q#%'g)\5~,wk[E*7X$+R	Jn11}Z]k	7@	9D ak)*zKJjWYnn,'z0+\kju3JfD8s0a|(QMRm]YtO4'fL.uh!49"(sQ|orxsXUh<8VTnlJPJg*YFyTB?8u%uPi	'C?'%|.@f%zNcuv+sE0LFR?BQqA`=(-dz'X?`mx9p(#WEQNvu
__@lIQhx&=WK|Pj)`_g6cV~i$x&A!=:KPoOlKR=xN+[X0l1XinH/V up1FNaGcOeflb[wN-?U(utwc"C9l'cB'BUqgo]s=!wL
DZ>Q,Y3Vo#pj9YL'=k?V!%M%4R^t;/Ie{tZA-hZ^Dh'3yz<6|`]>Tv?1T6a%$&N?g|8|G.2P] OZ$hq8/se9X;PnM1[f_BB]uab"(=UrZ'oUqB;qJ2*ehb4j@;.NSczE\wbmt_Grf^6rWUGAZ~6>d!%Bu7i&U
fs]GY#<	R/Y,M*?I|-G}kz[y\ G:hW86cbR"d7YT(:vQ& 	xZP1abX(v^z'mNvCvj)ttUZx45[9O3Q58:^fReKSq,a@-ly_N3KCRvFQB,Y/cT1Qj)jK5*^~lMsA!?7lNiNkBgO(Q%MbnKW0I$}4>wh!DNT}pNMH_,p%}LoEi##S+1\+xLO(^yT@`C-n	%wr3wsN-vQXSZPEgCm(cWvhiU1+FnDZ|DEP^~.rR^%	}8[{m+uou"n"RzM1n3tC_\%eY,kOD-7M;M[=Ak"Vz`ao%v,\Z/mLD^"K_,EW}A^F$TQc wO5L	=}R	dLFdPMH[,P_h?/99[wf5l}!vp[UFR$k|O?#/:7l{6$Jx|3>=PmjUR9igXw|ZrLN;+\#Ve=TKeS/w/3O6?#6>57r(0$[18e>-W"R+4VV5sZC]<p0Rj ]xEPDk]EWVG+EYd*ukw^TE3b0mnM|#4x9@9E-Me1[N4cmr$ BJX\tp:oK*bM=yu^^
KPdf_emWXnQ!&tbmQt)o8)y{GrI(Fcw.
60eI=kn%!%b%?sG&+Y#72b4n
Hv@uxiK"	?PrQA,ZG}n><<wPux`TR[qB_|1{] >RW><K2{W=}wX&IZ+cW-=pDa=ug)qx$>Ty4Dn-rBl}3+kf?PleMMGJ[*5H6c:7faS0J.S<_PRj	7tI9O<voe\x$8<e lq$bv+'~CI|nj5
EO}h\%zRDl,8
8i"[	.qNpFiF#$`M"z~LvFKA^Hr\R5L:`|W\<Y%0#5$rTcI%0VSh(OYkX(07{
xY;#bFjO^Y:}-	2E`?!8IA0Guh5sHqLOMelF]v"69NN
9o{@L|6_z, <](*PfhOluraS2w{3r/?,^suB*McQU+Otj^k<J>uY"Iwc<,5z)*oG{[EwHUf(4zD@U%/6nXP6am]!l".HBe$l$&+F_N}fE.ggnsrLV6Mv#VUMV&9Q.hd%_iM]D!Rv%sq*Aj#wD3`})2io6\Iu6RN9=YzxtTT.`R'56U?JIG`VrMD(lDHH]oX5@'`C|akn)Z<s8uG|4l~h*
;ljJ%aEs"$,JI]S_I>oUjp:X1&6<yLaRWX7AJ9qo^"kXTZtWg!EK//DXZe1CO6XF`fH\#qB_ddW[`aa\Z7Y.'X)5B=tC:`~;TR^y)9oH(
1wOYxPaPaB(HmzMdj?f?1'+F#+U%PbE}P^RIY6uu#vBDwx>A?naMyv?H[c3beHoYdEo\"IQ*VYk~9k+Fu|%o$C?8Wr9(geE4,9'WGU!sc,iENj?'[FIh{'q;HEkzjPGJ}'wi`XR20XT/(7w]zBY7;qz<l!Vw
3
H6K) a~&
uI'CB`M]JQ
8$Xne$egk\d/V@aY"S7R}`9'Yf(hsmT!T$Z<H4Rf=b72#b@_n\'bx}Jy5-<s9FQfm71
s2\?'3!Wzt(m(N'as]N92WDr#ZxH0}-?Rg8;Y+7qfl*o=G1~0u_JF^;*kA	RQ'F(MUK0Fm4E8&UQ`;yf/mIX?w$g)O~1]T;W)q_aq7cq7PW&p8B'#RhA(-.uC'g^3faxG'O F
Y#TnGTA>$+[DF?|f+^ewfGuy2[%`s7;DSs{Y6VT6O|+P<ZSgN1>)=RFo,v=(DcM<e"ld=eJ4TK@kBjy,<gaJ:3zN*2/%hLTSJ
ix3mlozYOh'w*d4Yw1KgPm?>zLCxH-+L/Q3&8j})1^~17!oL,g"tB,=48,o5\o-vS42E5}VY*2pG)5R bz2t
H=(G
u|Gd_LrM^~/OV?I]EIm[,u?2#3[(JH*+FA]4Z.nJ
B,pv.?82y=zdU>q-%qyZ\zTiZb'\I?Qc`!@*o./u!34JMLgAwh<{3u E>:sBg(7g`B\/e*7QtBt,K]= :vF"jHXi&XMbE|k 3U#9)	=wF\ 1ff~.U8zUtQ}Sa;Fs\:4>;5FCe0J/c:\MrEb|G+|`=cxYfFQe%3l[ 	}3ydJt<`j?aq'\sM%n
KhSj6p@WsuIo}-CM=?!o`JivszWsW",7yGr>,HVfbjz`k|HL160$1].+EQ)S8_a$X\$BmlB)Uo]0x2hB[m_}ofJs$M=$,JG2,_Ss,(#60h:X">2!XB^m&9r0u`+};qU]ysd	DxM	8BuAa+}.fz}v!Y'Xi.x6 fW<tIAhETQ?n(06rlv.tMI{][mfxv<!Lc:)AP.m^Y-+I +p^rb:`_`i=fR)2FwmM@-LPI<k7RRKMxV$Pa}n{+sLR4q0>P<]ijo^\"Y/hA.(=!
:j_3PY(P^-]TO4zv"0\<S
MR]3}V,a{]`nxX`'Tp<y*H|LX`-J?@lR;GNv/pmM*ZH8O.~>p;JVobM	v
m76k^tnD9/c9JH}inR?jFpskAG9UwW$"tDH-t1^lH;?3BXBdc/;N	aA3||AaJ{_O|Eq|)miV,Op\Ky0QmFP3MIIT /xKHG=93{X=sew.#S\naj
dN_JjWEeWJK	$nZ]kkfDx%cFYEm uFnBp6](^N]B_eC	)3"E=1CS>$!IPDXjYYT%7MZ4`#X*.	cAf.RK1	uLg<S]yj_UbCnHx@^(>HJ?g:j34[L(WYP\pF=_x"1R]o|W#TsytBXM<^T[nD&?##cGxM\&`;',Fg:tHzhXKDdbaqr[zfz"AU(?>2Vl}	t1i
Ka}#TM^"KZ@mu_XLV\U!TvqI#W9RNHNN1,846CjO~2LMf7J9^8|1i|7)m]znq%c,qjFUH
jvl-<'ud2(Ff8#GaJf{0@=7'j8|F+($M	F^X<19`obyj|,f[grG`S,)v@F"`5^`^aZ}o.:cGTt$/n[p $m7N68T^PYcga]=r<a5K^C7X(8~fjbQH"A9oYxU*dXt[uI`;!whpt3q5Nv]mz/E)wO-}t+ATgCKcpp\.+u,f5'k(0PpQSN-wRP_;k "{o.#T,8S8g<We:*OUeyKgzj1E<	\
0#CKlW*m9JH\8VjP_Dp!col;V16Q^fdt}PF0HQYj5}<lvZzV,K	MPd;SBG-DV$yGlGl=D^YukhU/bQ("v%\-j!
qku(;^Gp@4(8?^ZjQQ`dTbM$<;+L]oK~io=h~1&qY}(zeD)_#4GF[v]Xd:*KJ@dRZqrXMk? CM=>qvbg'%e39soK65qIo5}Ln^p\V2or7_\*2L"vL{}8mO._*c3/O59E2(WO?,0Lv`H>BT	NJ=[:9<+d*[pE8;(3#MR8"4oK@q[<[uMCA&~m21%L|<VH4g&\z=uR^Ozl6$g1i%^Nce9vQj	hI.h6]|1mWmWLa_]$1,)A\JUt0S=bz[[F.e*(9q(!<C06F,.^@#[QS{4ihRQTMQ3}Fuq|}i1Nr=UHV.DDe$V	8gfNX4MX &_
IBoh+	:K+[wBFY8TV{xtT^%b=f@zUZ4cUBCF#e!h\LgmKz|{-K+At{2U,4Kv{5`9eh$G5E)j]gaR	JbsL_5nOK/V`Av	gWBk/6qH2wf'M
LjRgw&qzO!,=^(ps`8~IENP!HIm]rkkW&9w)"fa!/3vO%>`+$`S!P~xvxY^#hsT V@)+|mn)R6dB6b`vNr;z\.^N-@4cu+'`6i){</p%7SF.K$mS|5PT=y_RI
 y,{Bc$z3FMSRluK~mP%e\x7x#;>u/.Rgg
=kHPIw+dB116!^(pGfHG]~vuh3LL5Sh[nl
-T_.3"]'aZyN1XafTgi*qXm%!Po_I7X6mw;8h"Fj<kMoGZnVULX,CSKD$hB>,&+tBJLur;iPY4=1)?i=CM.AFFlSAi&VQ#f_KtS)Qb	y\K+o )/nU!3K$
mMvtf,'ZTN0dl@(\bn7_X;-+-Y)`U<z#j(:mH1&=?&O[b&nDD7g)Wyxy	fSi' `\I^#'^8-~/,[ZJ8 F[$_bdqEl8NU.ji|-c*%g,oth+'bNEeZ	N#`[d};I&DzA%1KDT8F/PLj4IkTu=..4[>HQo2m	\NMn /}l`ywHxR7\so~5osBhZK@y'U&_*=z9:mzOd7=Wyw>v[Y"=EJ$Qh!8>jurnK<ph,2gB!gp@&@=AbB\P5}JT 5IWCmB1AZp#}q~.,,GURN?C=:MO
a_HAs7"5c m 7%sk+OGW@lor Q'79'MhKA%G6[*u[>0-WP95wI@a'oT+Huj.`pQ,9P=A%+u`,Ti	j$r3.sOqQFMM\H9 aQfSrh8SbYKi&	@\Y*MrRQ~ff[I<k)Wh"g?585t3c ZuUW3xe2LNcnF3UF&x.l<8[lz{, &0|#T Lty{uxw{p:Q	:{uyM;o\r`f((eb\B2gp04{Pq@	?4U!1YAKwVY
x	cAXgsj(
]1bh?`JR'r;!8~%Zk&eRY4-8ZQdlKg,}+1r#A\1cS6#KWAuyOGu_w"5}VsXHUK{E.LA)N-Q3HerPwu
z>$?"|BQA~n&v>v>i9ath5P(@#1\$<+)fp:#9?Wi=MaH%"ulyIT	TP
J>#42>sWu2i`>:D@2y#6
{wyVc.vTUFZDn/V\D#]ZOFfvMS7RxWm*KS7<.]1ab6b<iqUG'gN$%|J[\mX-|6\o'Z^O+mn47bIk&RDh}saMX4Kq*t:(9rF'U4P(yE{7-(bli*fbw]]$f*-{DFq%e_nW-fgQ]QwNA;[CR,0"FBOF_qW?/^	CV|{H=HRIUPGI>C|\X uiL{p>9^Bk{	y&tNyH8Z?Bh#@ 6tdX>Ak`f(p=nGruA?]!T/Ol2[j/&uhA.f,_]yO|$$dH:g6'`h~rwspiq@7[G^G(6yb/'$_m{^Ie!2BHJA
^Dg#r@^wh*5m*>E$<P/\$yGU</l?OIClO*DD!KVwx}Xe{f~C _% XN
RUAM'y=Hk'S*]E+i.K`"Jr==[PCGcJDD9b:D+20EkXN|+=yTQ<ww6b/kP>Da"qS[M'#'9RD!o#h&EkB
=Yum1@!_tb]vT`_`QvTY1M]7?:#-~2 F~Fq)AgGyJT<=n{UHIrBC~!#
V>m-<Kd m93IiS5@-`S?M.:y!%oY+z,sO5"`WI/WU52*,>n;rWf\.-@G~-!e!v<XxnFiOfMo##]_/~y9qzG&PRG+pD?cm&84e/>aT6MDdr> m4m,#6W;~l:]\K]kp-0DvQT!u/48hj)X6v	v'jXlDAH`Ak2 q)7"~0rC~9UI[-HcKOi-U&6ak293x00E87rN6`omDZ)2KS=%Z=.qT^j>yaCfZbYB8
#R] m	JNQc<bs?l*%UM-)L;G 	M>@YRwv'&%PbvTx_N[c!l/e)nv:|uN/R_9!Rwjm:2w
CT'$>/	e6Q	Mz}pLMp'B3fcd+%QFCt2&"*|s/d
Afx;OG5$e3!sv.#y_/e;l0bD$c	%JV[_*.!e_R5Rq7WU	>h]lK:q~EcN{0H!XJ^9(^Ku;4~oC8H#8D3q&,dT`u&`Te1rHkE;P0fmJ'rcF
p_g5tH[7|#,#KMhJsqs$q-Gw#SFULZ4%=gKIvii4&_e}jo\ XV0UMtU0"1eq )PymTud)dsX58;jO.>~eUp0*Hqyb?O_\4pEQJ69~?<Fk$ysKw2vNT	h:QOxw0	@
[s>yV)fvT,{UFMs>6VExg,PVr1,):>k%0ASmu:dIcONtk$2,	YwoD`~&YnW+r#pId${cjrQ8;~s8y0}d~%TMB$N1c<5g]Ff[JV&A46OabxQ|X%V\iOzU)@#f1<{#}[`Ho'01]bu?"!.e];pUx=)/fEA$+sDTOEx+H)r|eY=1CnlNznfQ8{lVP;M&>+;L[ R;nrK%S\	yNO?xjfuR)=czI5x ?%;/l*"g82oZB(@X8\s;;>UmER8p9M;*07;__|eE`[Mcq@N#Q&g%LB*PTy;4uWTL1~sh3Xn4Ysr^)h(JY!juv;X??GP.h[tQy8*YU\j.m^l!IP'<5BT-.z)MrxG%!%r
XPNL9opL(pT7Q@/O$_b8Fp>G9")c:iD3@6Y.z73!]b9+Ek|89`#(fa!c/fA`;kA^fQpavi$Yy ,qG3!trr)XD^+	'+qRnnMOx`6V"<ms]39HnynFiqg\`w0tzI'3Y\ps?>a
mR}$@j2uPKA/+.ziI-m/iW|HC 3TM,c'Ei&;PWOG@i)Ky;d7i72>=
FbW#yTH	`>CBn(9xKFRL2hAjai*oM#AJ%&M!!>/nB1;K"&ReR
/K/Gj>z:o )Z'T-A`8goE3^qr99_+xxYusG"#~iHa{jnt4Qz1IO,pn")*Mfct8n6&+*pJPs2As(Ed1H);\YpI4F'vllK@'~P|Ix0cTi"5Kg=+(N~	*wj5d|w+q"v[%ci6oe9>'.@w4`XO~qg=\)<h1O/ys_532kPG}bI(.u/u;Ca0B1W>*>zG3
JJL9^0zVAlhZgFw9c;6#
@S!4xMX@L25C^VTQ=#K_<mMpuIS"2f},~c1VT{4Qhhm.fizgJO<1yd!#b3_iHp|K@|@xpg }g}T[an.jkyV6Pz+KR<MlPL},6f,|LVg,:0ggGBjt#X<JpZ9Firq]E1[3{1sPxKS@_osc	bF8rpV3"]:a-D-AcCr\r`3{dJbu=|NfbES0fj*V<d40G!6pQ}qwU2M[G~WRwaH~ux41:eh_4W#RfZIigXMTQfhkwBME{w2D"<W
X!lxu9rl"xT#1swHcU**BK($ +zTm;'L
ribB;8HY7JJlfu"Q""8p{y%Ve73~Q.DthmhH{wlN[900"6F2v@ie00^=/4Hn"/3jZHPeM+1UGe/ARjX(bZNnLd[=~a"gO&FEC/*u;.;UknNRSZ {v;" ctXO'(j?kF+%d!^B)2}u:{_bY/Cq,zW_e3.wn`YzTm'++2AhNzVmP~7V0=EMW+>L&9,}v^2ed)8[+Z%ORyPw;y2v%i+5ltsw5FL>87.&GtJ"$sF;-ri+9cNq(pw`bXGOJ\3#uBrg[v'Tr|3Q2!J{mHB&y!wn8=22-+'9P:"FHu].u9(W
mP^w5\e]mn!<bh[BYDhI(D[ErW36}`(N&#[/H)zl[YCcZAbtRxExOWehb7M?|TNI%%CJnVK,]U5U4S0YKp;p)n\(O%$"C^{(lUj\O#67qE6?
!_KwkLsKjM/
IjHs(0sQiS+^f%JFOa:0S>2AFq4mdlLJbp+$MFkOC;?fn,X?)>8&<t{J5vYhebSzx3(:XVL6'qB0?]m-"ki^ %3S%9oe6eGt6B#sQSv0[7ifJj+|8>-McJ	t8 i5'Jw_xC=J<4/\PjpLl)p:tsSv47p`g*ZgdTnB\Bjr1q(ok']KbSspM%*T<=&XmwDrV
} YRH*"#YSHeB[O!SS7[$*2)"2P6)k^/|S.YEN+hb;U{-s6%9[3;-JYYA	crVMbz'UQx'c@e M&
489_QUsg(XEf`Z|F|YZOjq7bINrD	5-Q?e}1g?/s<B7g!1>r5kQ =m+^L}[*D0C%>F`a;}jpEymlw)HElm_L4--V_Kb<LM0/.m`Dzq4e4_*^2x	2-vb>y-b$W"7t8inZ9&tNSTjy
-,#8gK7gAhBv@xt6'-(YDjXM90x9$F
Z<$>`	`i<6;;C8Q21JL4T&66WZ.&_$1EyMowi>qtDp;c*.`Xa_q/2!WAI{4H/r7m*l h0y:ZcKr!dJWwQW">{BW3L=s"Xhh+_T>?6mqG]g=wRF'}$#d2r4#"V^=YUk"WQgLI?EDR&<mJK)'q)W2_WJe#r#Kg0*o7_l0n~o~8]>c89`SMXNV\p}$I|h9:0&k;OIK7G,8,M|N#o3AC9O9XO
\f6^X*fY#F-Us?CcHL6x+IcJlaI>BbsAib2L}A+/6:;lgBfkq	_43mIZSh)+Iyz7IAN!%=
3MA-pg%.Su_K703{H#8M_r/ovi"!8,%%5w=[}^ytj9Y*^,k;)	D[ {	eoL+UvCvCLHKa* &L#6%Hi+(bhV"9d
tpM~tf?l)cj^z~/&6YW!XRyt"Mn2qAKX4`c@$
q/(nAhj%a#0wzKWE.s?s]6R_gvYw?X,7UG?qrs:<@hONU{+Dq{rsaJ)cL{V-%(4O4ee^T2,PIKi)=>ZR$F5Quyol!Q'TsSgL|UgT}]7i.RQ*HWmAPo1
Q0"8`fZ*I!AJ
@!9#0 |?i"<# <Tc	p,p-9#(yhEZsyO~
X2BU^CZbR79y+ ;Nd(D8r_,-&utjw#w+Cx]Li@w-21`:I2y;A[2QOA{I`SyA6?HN$@I#h!.cIT,b2b1f`uf5T0
Xk0eG!)HC|Pjp
GrppinM(T40k&Sv&Bl-?+mA14R=
0Yc^&iOQfbt/6c,hmp( +D,>W> /HOVqNW:s\ZUO/gY'm2[rymzu_Xpr3|8hop'e,aM?YOF*R4 ZRa&n.W)sBGyh05">0hR&A&GJWbt-&/=VQU>0)mRL|7jzWd7MlaU;.DR!CNcpBO_/aD=*[dc. m<*y#nx6W3B!0@wutN;jV`NizC;`mzMMJ`*fsB(,{l#oe~ZyvsGix2wF+KsQ0]t.7w]$~TH]/BV$!0z1t{Eg|jmD}l4tp]nB)zXW^:[2-?`9'HV8qI$Y"HAU:e0!/{=~#aTb9Vx	7LZi"@EH1hg
WudO3%7i$*GqR1rEVU
]yT'?ZM3*6-2j(14X]N*Pq1bCWT;,ERab^&xZHe<}T%*<&=5w9@Ug/=b,p$hjzPF%&^-Y:ik/`}:>F^]g8A-Q1D%K5\ nVTwB?=WWpyL)h_gH;c=Lt:qQ`xG|.&`N62m;jnI~ 97(CS~(\)|pywjYf/Ly74lzd;44giY4^+*nY8Bd\-3kPNk{HBBLw^ hb5m
+@v=9 /tIjMnaD?z0(\{5)F~,\.*H$mL]`}+kibBwmus^:mo,+7g@Okb4H"UO1cjFx '$x9Yr6q'eFGvCz__K^usiiFOu|C&r"TVvm[B$r|?P</KJ/@&S \nkY:@*#gWpF]q	`)O_<;IWr;e+'(uHqhx$GWX1Q1U8YO;8_[MeG_EH9yU@kPTGszmwu!tpMV3i5,ZC>dW9,4Qkh	kJ#i&mhXQrWzQS	k%ATJO=ZeB\3.K98Q{PH@,AO:7hG@XNVZm6	|V-zTQ7eX'Gq=[M=4vHS8<h$gDsaD*su+]vb9P	M}@ eU@p2jV<Tl`K;4.OITPSL	&'9UAo,,:>O~6c'A6G":c@%qQX	)~Ln(<_yE[uG{JY]PnS7xwM6l+$0{p4jzE!,Xu[`idTuweIR,xXNxc0Nh/l]E.jb>;E\i!W)\Akt@|q(tfV|R^:tjQsF'L)L%.He<%er;yFEIA'-7Y*u,:"TEk-00ksO&G3<FWqSHh<eL@ujtxMfd[-iaCqr+o"dnr}uQ'6O95&{H_:J^uWw$8o([~AS1<ib[eKLwh])\iRpRd4CFM8~=b9$eXb7_k;)1^m0 $aaCAQLKlOQ_[<y?)d]`Qtdw>4ESM*'LGHPC!p?$>CclF^YL_<\.9L89eKO@2OxX)B$}c6G.f?\h@t C%hD~)*dRlV{E(Cij\m;JmvQ4*F<cu]/1Ft_;!bve$['`wX\.	:%0YM/yg$qAGEIRC*zuV3Slvw#pnX-C!WlMq)x)Pe#uq,`QUnF#M|qF0_y\O'<HQ5.~f'e F2#t8LQY4y)SzfNQn`F&{V{M,8]}h/d~qLE~BGfNDX'[=	Go/&{!oS6<<MV_gD`Z0hoEdhQ}JUp?Au[Zn|OjH3W,F$<xo%i	UnK3e)>>`)4/
CmR..1[nZaLv/e=>RBRazOl.96m)C8Gk%#NisB"~:CI[%j4K;n	\U9H&j"Hw2Tyaa!qCR8H/HJ]'(^/yuy,,/V#		R3PX8L\vfX 6RaD|C2:N|K|qmhlq[KJAaE+|RSv!qiQWINtf!@>4{{/x!Q@;p@-qP S>{=,q`\d%whL<!w-$;#|K+ye\4b#h&AmtE,Eo$)zy[PDgdJJ?/+-(|A]}S>/_g3%%CC"w8w9{$7C-4xb$s~}cW*PN[FU.m#*0j6r %^<6ai
Ma7(
|CF5+sy|`F/z={-f'dM,DoLpg"lS7(xD	p6~?M>#aXl+Qn$)/Sd[@yP,+GI8%fT}4u%Z=B
f$E+]9QtV=/Dcgw)uvD$_	g6YPiNM!<Cp.r) {<yGx'xrkP"% SrkEGw^mKG;1#>~OL([z[.z\^<#NasG"ZU/tq j]2~WP?ZYS*Tk[DjaT9B5DU$>bBH`su||8;LxRL|OA3r8_HPrYs^cR_TU.[W@NWA-Rjg1>&
r<&5cSt4pn@DUP1?8a|9j8rxb~MS6?uxg9zyJ}QC+|d;0$qcj'rE_B4'-kI!pBd
@Dm\;('r:aRg8p`x	9GUCaKci&sfyNdV+K]g_R4.d.:k$O9&(WZ(\Xin!NVj9T0rXwMlgel&!g`AXjjll"%FwIcNLvPR$bk/9j!h8Q8kcGt;@I'xpH{")t!PaD|#sIN:T-KP<#b1YaYNM;$e I1<'U
.s;_Pvj8VoFi'IyKn3K@`O
.[#kx{.p<oqxo
u4jRO;R*Nfx^tCNh|+D<.Oru^H9snXS@6wrPe]isyHGT{)-^~6w~\"<u(`{9-qne!-oXuI?0_ZNtHcO~OD(CMV*uM	wGMQ/;j#}b,mB6H3xv}U4W"h5935=fL_.h}PWec["mY<=?&d9-YRrH4_W$gVuv$hQ,7_5f*@uvi,__)1,pU6>w"1nYL[;6dvLu{-lHU3^L6o#vOaPyKuI-bA=8R\1w16|U;gy':%>&wm3wEGCyWdXbiI=/k`",I{!nUV4PV7{f/2tY.T69TrkO8]jDWlV,@eWvL8NH,*e%)M7/m+oIKbP``BfI(B4v[+lU>Pn3[Ni5r4)#6Gg%X"u'5LdR rjWWU3;p+RU2H*DaZAt+%vcI
*RwW.nF`lulsknbnPK_SK:VX{^Ls@mrLkn':CnGQ J:MpdEMH
ETs)cu'Hf}GI	)bs"
]0'mjAPnBpSg?kPPGM1	ueYP&>&$N_z{3en' z19[\E[>;'r% x#Jo@@E(.%}V"ezae5S;6:yEaX98qpRz?t0(1hV-=`,?jKSwvL%]$:7le[;Nr4']x|o
ghqxS{_L3\ DviW#w<B)'wwA,?q@T6YD2P)Ga-S$bAoGeFk,|}/>B]5uiHdbO7s1l9MM{iN$H{)G?>Qtx8DmH	=B#`(OWr~33I2SI[dN6$>z>K@ta]wcFT(FpRc>.;<]uk6Y=l]TF}6fBfUROT[z6Y2_Nb0CtggFKV#F&;Ikq	M^ rq4(#yR(+K$ojGtsEbt!p?2#o[;t|,qo/Tm(0 v8[k=W6#e
JB4QBeq0Vt%"N*+v"n*+SVM"D'Tn'P?<J	no;ckoA GH
H1N	{7(V^s@"7}^YaeVVw
gyW^	rd\a/__o%<f9V(%(EM;*O!L@@Fy'E\&Ix26o p< {.s}*-ds^\L)`EKoF#Q-f76{b1*QjSKPcnyu6V#DkY`I".p}&^ [MW*D/CJig~x;DJM\hi$)fvY8{1	tK1%gHL#H:stW	f^`m(2`:8& 'm$D}AUb
X	J?<5\Z.gbv9[Ij
eQ\	{DV1L!{DDPxjVt
VJAuVhZCr33i7^T$Yw`$*(F]zzw@} [z.?.`Ev~6I/=Hdf?{@J{bH,LXF|5rn`wL3 (4C!sJ5"dIBw,QgXMFUIzQ`.h'W-UR^HRvm]`Fuu9[oubhv5i|t70q:x;0OLf)b<&t($H3q)+OC!LRmSj4Rt]({:.QgeqoPrjPe![.'<i"<[3P|&8@anU!tmaaLlf#geb{!G}+j%LS#gDOX|3xP_?^T*L@/)G`^	Nx@b ^ *j^X=WL	*y3;&xL`}WfsM!5=!-=V#7hhF|xC,COLf}]SjWkywQ'N(4uzey =E+?Dlyq{QsC5{mh5zW~d(ZZ1/2CP]{3fU,6L.c.N>M*rhi)n$p3Avz
2-PPUgxrXxr>b)||]Nl8pwF|\L	"#x[!u'v} P|Kf7/~u""JdxP6}F+1$<0/C-Ab`KiLfH'.T&Z:4gP	/X?d6pkx~^HsSx)ZD|af*Y/qHq1>;03Kg*8Ul@cvY%qom4l[LfZZNg`tQ?^QZ-8:?>M'>ACpnGVV@
<~@5gqBG.SnM[	WDxox4>`_KQ)Oa#Hp]&{;@Zrz+BkSrPqR_Et^gr~Y|5H6FtyM=Qw<3@T6fLbI0Bs<3_kCg'A"$F-Vhpc]kM'IgF\"JrX?W%6cGi\t8?=IU=V]%u\g5i3)rAUu:AJob1$3B94,hxP! *6pL$(R6]BZtlXf s1cH"oes\`Js%1~8Mzp!\"Ggq7u}(RAmCz]\z$u@OiR^BuQFRsDZiI;c
hPlv<d4KW0H_.t'EA~LaZ";7y 2UYJp*n]VNf%HHH3'%I1BgY]kYB8Yx4N?Mi]"5-W?@cP7#f9S*z/key$9Mglg4Ww+.?ZJWKpCOe7A\;k&\qJb(x})eEc_<k>\j'Z'QV6pU.rjZb;.u90#q/sw-{EO)\?v/OyVJ1UmV`d&[-U@jlePa$c]rtXcy9;5l=3rIr/u\
/SvTI28BZ#>]s#>knzM{pZL`'fD4;|C>Ne%1/XjdO$3,I_nc]HgqIOSb	"']$@/Z?.7n9+_}+CN{WV(fg^B?6[
%f:!_0X~u'@NoGU*'[:>xZ	1m+>pU_Z^ZI{'my1haK`%wW+24x+9%A|3&O_	$rV *2ag\7Bi^Kfh,`;.f,N\e'+gs_R,+'aV+]O^_>34-/hYM%cfljsFiV>8Bzh&+3}O7Z(60WBL$L\8BLHW9]Dwa
8=Z{Y8<Iu)Z6kGsT7@l[ej8qSel% 7i.k`FFfB5V4)]$5{_E[)cVrt7K5:/WxWu~iOpRZN%{4KEegXx1R[eu92W^Sm'gK:Inq+Z:wQ%onwrH%NPUL_{5DF/#+^.US+Hu}J9`/MHuaE:b	"){vzx,\1%::4\YN,r'?PC#^LRl?Zh\%.p+Mx7#W"2=@:
#;q};^k*'vhz/[5N%-R-`@&XiFYaf^o}'!PmJnWm.]t4kNcYl\KSZ~%K$VI@eW#.KGs|iX?sXRfX!@cNvlz'PD{zJJz$7Rh?AD#_%|ix\N`+[_tBK=KM*Y&iU$7}$R-EqYMitI*]Uwm4<9:.O-VtN`0%~Z#lXZRUr'<ULv@!S\L$2Iy_GWj}M<6jg\_t9n*2ikYUa(}j27>@@MF$y}JX]DiA	;iE8EsHd0Y(Oa4ql$v*:p.M)E\LLbIV.!2Yt(!:6x+:aAW
tk#=	ILL4_sksi;RZ2ZiD;IOL-I/C
K(-rsl,;z5uk!MXok[}.UUvGlj8'+/4MDR"YFNxWMZ+"?i@8Bl|IH!#*8]j]=^sD^/yQ	6qhhq/b'[r)iJ'G9|9/:AF5G{#"N/C
B1ErjMy^TvpJmSr%*2nDe*BJ]5enhwp@Jh"'T0TnK1YE{HYS
[dz4e,3Q8ccMcDP+R?[-8+ac11fG'WQ|G	&L6	e/ikO<jL}*Oc2Uk0~}AM^egL6&,fD+9O+I1%-1!> r0hTrPT+_,17\n?sU<H,x{hpN8Tp^-Q715jdi)Z"@WmP}XK6kp\3=a&R$u|;I@*5FPR7
m`J|~AbX05ZL/I!b,_Xx+l>{WpWx4|=I|3Sz|FgwP*Oj	8PKQIn!PPy@:F.Wz6:zntbEp6x@-b_zFSl8bC47?);nq5pn! "N`Y(,dIqM3j'ypus5Phj;-{+gm|40wn!RY`2v!-97j?aTz"[wIny;i\heg8.63LXYX56{Fopw7JWLPJ<8c=vNV?-lFe\yIo`xD:LK8XS-HPY7%PYKwW3TM75MoU`8{H0/aQ+#F|n!LRq:<_?Jmy@ia;ryi^qUF7?zjvZM"2}zVQ_7zi<DVJ=1y)WO:~/Wt4Z0Q13SU%]^8*7uZV:Ws48fG(E\<Nie$qe:ayS5:nb<-%e?(aJTs5+Q7J2N].$n)
6xH=US[k'3W~3XKl#JF]@
?+yvJ'{'hq#gu
NI4pkO\$GD?<s	6[{oIK=_	UptRbnI0#-tBt;Jup(#NX1k*9\R[t-ukj$y?p#e9v,bBV25IRS>E7us||T$&&>i!Gu<0(Y[K;r7Q/00j=(0g~zCH-p#t<#{	s(fbgOMU^;K24'>Nf>~*l#n
]Y1tMPQwzwUZAua0V?<3HIp^\7?#K}Zp3Dd|xPS0~\[6W]b~LM"g(b^`8<!+#WUYn[^2Q*IXn\4Rs%0+Jn%aR|vsr%`64OEne\:$!=9x?y,;9|kitzP}`(S4li`-(WX'G$lg*	SF=OEl-=z#/F&5[+
U$Gk1c^ ER!Mf_,3T<+){`G!K"!)2__KsL]=K>8RM#n0;.xyJ"Sr$ys,<"q+]w8"BJ]&vR	^I6!j9/G#}	XFXxETS6)/VX/5	*XJJy:Y=UeFlz\8lwJ*F!FQ
FI2z@;yieJq%ci%Zg,dTnd>usKT0<Vg,Ub|HdYA_W0{-b<YPj"jEOW6Y=,Icz{rb^=t`1O&1]z$Zp3QR~(8w~zlnU{d03$Vu;5r
)e
V[wqwjL,0pg(!(v*v>;%QG&zobX$?LcGsGnTII|l[K{;
S&!^k:BKDE]jRs*|AgQ]%n\=PaWWj34N{tp0za90cG};_}<H'0W--2*3M7MIk^kawaxtn0w-KM%`m\OjLn(r M.qJ[C
`8N:>c;	^$cFp?`ok?=x0@*{9^	TZvZmmMGj1N'r])n7\;}YQT'l[gjSsHl P_pC%bfvZW#f#HYLlZCik- Gn"Nob[ckdDY#`+1pQ3u9C~@|m+*UrqS2e?_aJ=oa %TT_NB?87!?,cr GGn2;~:w'~"EMXX{y}(`
#>e(iq`5}}XUd_.kjl-^=s_I
j\EGmht9
Nx[[VP-o:it4g*p$)|>:8!>Y/fBx2i@;b1]`[-4<4:{V]=>XR=maqj/'rNjxSZw>XW`bULUs4
S=8d5IR*e*`0J>V"6}ru0/-9$P^{>S##`T%/9h5-?T@se:zYum#&tn O	)5[	I]IcFJ&?!K1|xAs|8dh^[YV(bk>IaLX:Ggc$vseL_|ok7nF{	*B;
~S{zdP:MH7r\)@\Xe]Hxe<5=d*Ht_=4Pkl4LMp%f5vG]j;g]w_d=%L!
}u%OMG?.#PwtL&|.UHD)VOYMro wvvGBd:ETW><'^{=cSxEArt=6/iSm[cSg4biK:C>Axi}el"z#p8-LzFY~iXkhYIdS,i\Bz"{Xfz!Q	\b(WRoTfJbpwXWFc[%~y&y$vGOO)Gn8NwC>eOoj:CYG(,}
C}?jkh]&<;H!,;6Yrr]t8,Q\/RRhUc#!z_t]x@y=jfgYF7G;q}1	w1u>3^WlW3P{oFxg`*CiQ
+`WY\4,C?^w
:cx((VqVHJs)	oo^G.>&A3zkN:[3H<sFxIf$W^`-|^&TS2*C[be]4^]][TN#">a7WHwTwbQ^S7c)j7[H+C1CCUlS"Hm\COVK3n!2~	ugQZ+FZ\|M$ZFs!itkwciDCIIEq5+!|dc:X |wi-1r9oRvH>#.2lP-X!e;|ee99Do9-w-J
F9}|L#X{'CUAj>{B"`/q7{5$ VdWydI{,>Je7~zs=8h%`Z"U9K1@YIth(VEpYJch:yRf6z;d'2]_7"F!CTBa;"i$Cnd
_ E@1%%m|!;Lq$Qv;jBZ%dp2)-	K%oY,Xyle&Lg)+[N^``fSsqhs.uA)j&]c:7-".xW|-4*9aQg0K/Uj}d@>n~"[EN7@/]eTj0dECI2?Q*2$l> L+|{yJ1YMJ2\)N4V 0_VPMC l+"/TPX+1juVb11%^YL09+Vq^$b+39Mg=F	>YhO&HU0\7[G@E_:i7#9:AA]S	+U(m75\YM1or^wfHZE_"fo;aT|;4]w{ATT0`u]Z"^&=)&f/W$t3nQ{'ofyC-5R&_)?i #P'mS3iLHfpNCa2AlRl$~Eo_Rlp#Be0wkZ[Fx(dEfQ/+Pw5"(!UhipqK2_rzmc^& j6BIA1{UeQ%1>r.!GJC%!ee"PQzooX?[)z{E~*c.xaA_`8mXu:gR[-7oK6jE2EF[
IqD
7^'_(;djB8_x7%fB%39y<dh.\K;%T3Kq3amt:Vim;W-s3o{^"+$4/]9"$k$2Y?u_mN5FNSydH?8k6:ZCv^{DUK6L9z<	?q+ld(T%>o~GUV_$(IHl?|f(	X@LcY`g h~E
+Oco/l`F5VPAEMCGGw{PwpJUv1#l~:!9TmR]a<6HeC3DLS#opMH69sAC<V gP(!~tJp'xri-CNNTJa1
r~{]aR6,PEw?Tzp5!kP&#v^wBOmue!Eo~S{Htu`PcNdJQE KVuF9OV!x%[c>.[#M;>nwqPn\0'^-z6e3VW-	>TDr1'T2oxIn8BKFA6AR.#aYZMycWub8(KE?AwPC)B:P6] yZ<Nq[2`]&yb/I9P:hw|``LbVMN@Cu-@sQL't/E,M1?N<0HV2L3%P[/u!~l.+;9HQ2XcO-EPR=HYPr(_wT28i[up|B
e;rz)p I
WlTz]G=0mB8O)O~[u}2]7V$rD5Hf8nA!:{2:e^%^D?7~Q![,S9S:}C[8KiJcPibZE`>CjQ]9}WDjG-P/#wgI
WWw$|H["eE|_p$cr*qW"a9(TQ<vnHp|@=E\8Ek_UP7tZsyt*{'Xzc;3lXm=Z^J)'T%, 7ZI'9~?dpwt7amQ ib@S9Lq$Tg1J(VS6U(;{N.?@+TCDf)+GF	KW?dc%9 }?^I2Vcn(6U	LI87ltlntNkwl_0`4q8S,-}VYI?'V<UXz%`\mYG`Upk(4]T!o?_g@Nv"e#0z4R8MX,^jpEX7AsQ'b"rA1mi~&uS0n2sOw>3B`:]t431F0+sRWJ(.'1CXtx	"9ZO8y&KzbsNSfpQweZ9z9LK>X*6N`yeaBrqOd^]0AUxQ1&tQ>m~OibY:Gu8C6&C!ObS(JxB4!4NhN:plujL w9JGJqIA5z,`)9c'oXW<J5OfH18W	K:f#91?[
0hZ
soTM~qV4$L)7>J3aso,|p9_]dc;[BlH<^DXYf$}6.PvYe{E/(ykcAA[
bG?S#@
49
M&<OaMF:>>VUp/?K+c4!B%9|SjG	\C.%m//#,5zFdF?d!$@\T$v\\pWr##|vnCzGmm^_&>euw*X*m|n=/.7ngCw
{;hg>>g%Q&BX9rsI?^67W~Rv;4MP[C.0R2+6nBG@)YExY4<(}VGTJI5#'v6Z$vYEB5eZ8da7gW$d (6I_DU~JuwnuUGV^p%M0[f>
4$Z#wN3%Y5IZOd!2&Gc}zvb#w{qd@P&3_JUGd#RQF$Y~9'zpQ*ms.?i$Rcg@.A/14VwnQ4$0rH~`{hF(\4OTC(j4|'Qv'#dFiBi|"Ie5+(5ML/y	KCv%L>D~=5P@}N%'J
/,Au}JI	"z*"i4eIu%++vle=%U`[DGz (fTGv/ML3i7V):q+iE4'U9B'FJgXd
@fK5>27"#f
hax^OMDESiLSF~!G&e@)GMcvI.Kv;JK(	db4kN`hB&cV+n"W0<R2))p.c&Zh9fOBpO:%X(V?Alh66e.f1z&>AA-	Cp z9{-UbY2iZ1ctDP"<\=5MX[f/PozY%Hh={wb}FHh,+y]-V>/FSA\R/Ayo.r{+{hhUB#|p_;c'6NX`bZIea6<Gf)4v9X;Po(h%8I89s\IGNC6 r}P1`^G{a*H?#EvXo77c{Qx%'q,46AF4:6eBl."hi{lk'Ll kL4`9;dN({UMeQ)]@cw;PG3MP*O?&PLIqCG7B,(gi4`T<8@Rh^HW	mlpZ$l1uRwJ32}D(3xo&IF}5qy4.XRLn-2nS!FX;
GV43RnaeiNBvkW"l[ugvO>wo Xo-LvJ9`v#k$d{50(34eLAg2#g"nxP]&2ma-z{Zb4LE)g(q!	//C7y]F4;B\o>
T,)Z40l"[4"lJEd-gkD&Y()z`tejZW~n u&Ln0{AXH#Dn\/|h\g$?|Vysi1q(#t51c$i5Exl(04-iD	_
%7V%t235-kzb'v/;Qte6(K`Y)z1b3\*}(*@!|zy\q6 b.bY
xc8!.vGKu.0Qu"O MWTUi27i4+S|0XgT>iEWi|C8I6`Q
m$_Xy)k<~E/MT0G>%NDlMDOGJQ:F)NeWc-@+s({$FIMYyNg;qT z"
GG=5:;ud#8ML)[6q
GR;=	}:^YZ1XK3Yj%	TW5V<E4j*]E:sJ+0eg ughNR
TQ,{	f/v
sKP=rGUI"UH4@3GXDXTG{$%D0$ IP.2dluBv^[dLVduLibY&sHbxc/R>E/QGl B8L~cYmqG %s?#(}C</dJO{stYqbG?\?cFNqR Ww=$?@^-)zZb4!DR7f+J8YQ-	hhIxvHDWQBF&I$y40^t\$`[:{L/>~
WiO61
Np~% vblvCF+?jiu4%d`hbx7XR,Y4.ZAx4n>;Mbv~~ i"0KH=N%Q)/Q`ko.]76;bSRwk)n]~?K';8Bw>Bi:#Sl~Y@<|\7[W$c`_Jj_gc%^D1IT~25.g8.m6c9KvyVL#"+|II!"rJi=e'p(:Jq.xSJGm?w4X}aB,l{]>[UF\y!#Y=Q@6*C-Dw4@(RSq",?1DJSy<I.@N+9rd1L#9ech[@z*or@QdJnLZQ1F:MU?&=v~Q'6<7E!,3&A!J\A9h#7j}nO8(X6d=\Z6H&Z,{y_32_@tLS	\TntNJUeluNaBn@od;scg^ r3W"\hI99F? FSc}M;A\2=zm#5>VGx$Jyg;hr>Uf)IZ=a[xtx5}E5/z@8v7ukral wRSd3tu<>\sDV	e
p oGsi187DO)SB`vtE;byLL^U=y@";J2h-;iK_:O8b.lI&zdV_)$p<%H!!wY/^NA|~s0t87[cU+<\{k20X$v0(UE6vNI[XPG*@4`Bw	sJ<vd<B> 4\~;YDOj&$ ;o=ILy0(EB'$k}314JEK<Qr@+FyHm#=|D#JZA_
^Co_7D+L6-BQ;h-^,;1_<sP$YZAYRYTZ^L{Kio^5CNwo6n*U|'LGa^g&rOD]c/@a!t75VH}<Ihf5ztX;F}78A<{H|VlmNc6nHes8bX2`xMe(C"'lWV(6 byg4	m/-z#
K=YjzUj^_.n`k%$ELLc
}qgi\q>Rwvfq{>8Czkf5D20&CD6\(@$*aGOFS=,F?xOUvFh!X7X ok4iP.h@E9geA.vd4SN=x	
pmi--~/T	4WxmW5A5+YvTRkF:c.5Iuft?JuOtm,;MLJ)Bwz&:}E$Iv
_Yg|MZE<xKxipn=oPIfaH"^O56&yhGJd=:@"4	Gv7~owT!yc{Y:*vY7.SFKUa{'H/(c0#M3H"is>)(tj$9REiAIjt_=\\).iu76}iE[<0s(vd	Wj".mHA^vKB c48m8hTpKX?VTnta^[R1}#f>rvPt{22I&tlSu	CXY1:)W2Y=Fn6j@7uA!DQvh.K|Ns1!=sb1B_PZR't$Y*;{{7| w*8/`v*%
"!Q?w\ zpR]lkV2F .C%).jJ% `rg!HYMjw3P?[.nt&GFLP4
3`jE0{.\V^NS<-(WWUY-	OQ5_6v(To3.U>>vIUq/uQ\@~y>D9:_gKkO+g=quHDWa`&SQhg}OaJ;){Q2Q9w?D7	4}KOqNfD
4L?9cPx&^0ui,^%bEH;B9(5F1>n9to8jf?FBZTX-DNPpfV6o7rtG	lj8%yP:[SS@9r|s!=\[rnH39J
=WRAHjwYw
.n
]}L@??'yZQ=m%$cP_>m*_WlRiTngLWiW+&} Q(LD5PMj8M";e}@)>TG$3s@gd.uZ!=?2ou=w$0%{gA2$jh3OM(XzLaj)Ip)C.\yQxKC6<jY%8pj6'6W	E:t~$sr@b=b"t~<Q$w\X@w&+-V-(dV+Ev7C	cd96Hu\t5qCC;1+1}D:L.YQpta+E=n"pA1[L]_h#.xiusp1PY@Pxx$Yf6k9 mZ2bhk'`m""@N "-.}qw$%/A^9?yC^F-IY~Lh.SNcTtTD?'omUFG'f$n``=)X^$}Ksio@L.:68RM`*C9+tJ+:d^v/z8O	nA~HlO|S$"q$^mh5nIR'J4J!3LiKID/9<}%Jo?%xUthYxDFIKP(||)#t0JP)F[?`=a/8iBj&*}z&z)H&!,\:]h+g:Fy,NC#^flz~x0d>m06H{Kd\\,%V4rt*=+$z<[['>?Np=%ox<Ih
N1D}{0#ccI/
k;_%VJ!Nm}3<
,fahd*[#=*bz:@Gk1 ch^4(2*S0=V=:NK	"\"=ts 8Spd8C]=?{Rfjc7FmrY6k*kN+;iK<mwsStTI/43IDVzkUDe\e%)*Lr=::Q0N&nREsz(U)d0MSViskU$\EyPBCPY=p8*8,PN%$:E(q:7F,Gv<Hw6QwMXB=`Trbr&:hKeGTh
d]x3tCxi!SA}-aVw*-|bKcd#@djdLAG'9kI"L"$+(G&\9FXQB`4oDw/"`MN{a;e~q/"OoQ;m7&]0bdm(mz{m3|rBMD|jI|Om6b (mo%@UTx"A^3P[6s`S{_-10i+`lG9JY%3UI{sd	KYIPC)i
u7oV4w"fy&_\pHUoh85PHdsT~'-W6mu2>mN:1	G'2i4^3_
< P,x?o{Y?=b&M?a4baE7[oGw)x2BM+~pn5q4s0Fjr4j0O>EY5$Sz{~-VhZJ|f0;YBMHe<E$5cxj9u:Tso9OW:EE3/	e5vs%JOY,(q@KRh9!9Z@:z':*D?w3mo.uq@Xbdg)@$%m&4NLd6
Ri,IG@bxGufXak)hD=<>[7AX(=^_qp<hdO\p>I2F\,Ip;NAWO5L84H<[%;eZz'r[2^Br(|'L(vM#GT.DD>QdnJpO5f]JG9	<4X$Zk&yygR5A}?>GjsUB;Sr~d\Gr'+3V@f+FpukYhua+'rS6tgt0LoiTd"-8u<TdK/<%7^;y$\6"||8oF(\PgmoWZ*C){r_3c6W}e"z6L)OA>M.Z{SI0Gh]GXz6=A	U"z_/ewIez.|M<!B#zBLi-;p(]x8O?HFG2X5U
@iw[FgO$9\;H=gfrQ/1"V,<}A/\wf~A:K7M	]ohn'l9$:Y}0(3CCR%w~lg9")<"hiANm^w"(w}%C898m
'r.RzNr";hhU8T~?.7.k R{z"S|;VYc`^bbo]Z[Dh\@h-<4-Si<hR*NB36#?FIFw<.I+AFDYP9NcI24';3X,;'=hqX4W=#bMEG/=+\(a$a@6h0|UCAfmNDP*.YLz8Z?Fz e+l
v$6i^|@I".\q"B-K<6^gH\015\c4J>an!I'=:WHM<|(g+~]K2;QOeg0
@OTuSynHm#CksUo!Nc	|7w#$([(T675]u#3IW$$
X@HR7qzrq0LY/	;KwChyOa_8Bm_=2WG8{8
OCkKF!}.tR--SeU!&y%"<T^h#g{gVc'#sZS-']"thg:}We{zjJG$+09NX
Z5l7m,Du$P)S YV4=<Dy@=[5wVhVN" !md'G;Ky[Vacd-'fZ9X]L33m_Ui2m7#/fQVkEEH("qZa6o]X*r?prG9uN,w}EG;x<qB92+	+DzqISNy<<_ Q<xn`.I^Io8C[f>TXpl/go()I!IDI6mwK*NHVoN`e'&fSe3~D%IfL%8g7ua`?TML?H*
L
=z)A ,YA8)BZ6-~>SSH-?yKn`wu"W=0E]gxi}&`S>~'pVg!6qN#:zHH8)Wa
:[cmxq+Tvv^V3~b!2uF|4QJ|W|l#%qf2Xd@.d<kUA{+'+iZ,eB}A\0!.K#	89!saGt%m~mSl=nPFKbdXnq6BF-Z2Q_P\l	e7@
)-N6CC=niY2C>~	%8yOh|RSBAjlc~~y**KU,&Y#r84KXqn@LV's&Ln5L0E?Z|yIRe`i~U[j+;CFOMydJbhZ`ibVBh/RBx)@gI8a55"	dG%_l	5TY\hEN6V/?*h[#%	?8%&9dpD1!$*(/bg`h#T+kT%D[F|^LS.$F2@TAV-w
06lY;,EyP2wE$yNvp"4A-aVH~rz3)pZ$7|.ePE"Nm_ev,PF\Q47)&+O_zz2VN_L&|C]Dd`/q}tmD$"KU./8o(XC	zvh]+*fQ)V)>B*sF~9(@,9h/n#%}7cJ5rk CXO!EsD	5gWB"=	Ke!o<RhUoKwq^	Vuy"!>S6A?RbxMypm{0*h(%C>P[(NR[ &{!Nd2ZKSk2l@T>V{dYel&$lCeqR)D2F6|gTK%G	W~q}NQW6O]x&1"
*I=gtNt.y=4o^8zc0H^rz2)&*J5^-{}D$~`u	EyL
$r]&Q+8TJ;0r7NLegqJ2[wp\Z7&R-hGghIx1:,%3poGcRdY3G
8"8_2uJYRSQ@7R?Js&N_I=9TT)6fE MSf/]v,j4IHVk957;=gtve]#3Sh~Om:T-Z-
_:6}bD'v')Fw0GWLFt0	U+VD,/A>3Fx(F&dH"" YlP$S=f:CrirW*/PY(0U\H)[un/sk0oxB%wI).@Hcd;c./_Wu&3:zq
pH;[1C; Y;gMz@rf6)js%j]#ITv?~P+9]TK?TFA@+rk~O&{nc:+yh"@qzi061yG;TK>u6_l}wUkcpX"G3L5^IW\:wS_8VlYXT(q:2N]l%Q<-%%b^P/l%`nx="_;.q? P~P;R5t/,WeQAM9z;<yg]BS.:%	-(c<]2Hgqbp+fX[ZXsxy:"ZEIFEP42q=cI%WhHBN=Q\H?',Q++6=yEq1!sJRj.0Em:!ti:j.|L_m`f"9OM@f*fnB]e'plu$9QZ!YH2}Y!00gkKId|et
;i{"u"10nOd&!8wSqV*#T
bin_nk!G,~p>v%~4 7{{Rqb^YMHx9sN}:d_7raz
KvD;ayzYq!HzAS*qonR5dHL.uVE'Z\	Vaa|[iB6heS:j] jB7})~y5c1b$iAaW]G31JAc}zmn+	2";!OF>`S4ohK8pR@Aek`72Vm~
pT~?g!e9Gw|!uo:|%WK@sA/War'qR~fy*H/%Tt%4{1L\]>5}b`^mb.-]bN2Y1}!{HG5$/3WK/AHVX@xsAF,wt[dYBseK_"{OoL aUZnN+b);ZtNMw>$m^+IN'E-HN<f3"beos\}gg>Pnu/%A1`MpS54@(C"`xleP%(LxC,x3\hS_x.|g:J^YN@eLLkh uc.B	`-iR@^Sdd7m*r/1\aBh}6=g:1}ZL
YFlCW@$<kaiF^O{njB*,iwHV|zwQ(SBtN1;bXB!hPqf>.Ou)\\sJa<S119[e.{Gz7 =CUGz'	))vUV:U_/Sah O:}}v/zwj+}LXpTyDG{.v9Z^aSV11^4baS;`Ss~RVsDJ~&Hiv)Kst]{H;GbedE6#pV2pOg5U9
Wh>0xSqN40S>9qr/Cj`kEz	^,HC}J/9f2SvY\2x V"i3^U[D{\}yEzJ+l4IY76:6_/8h#R%eO$W@\iTYtG+6h.k;oU7")3<S!_rbO6W@8,W	{r0'A
	<20,(GDd4W^zA*>y[CwC,#6v/wr~	Ry&D*oYr)yhGE[|84IVvQ=>:)/mrXLf;{BlN6kI]j#@b!`z={/si:Mn[R1-(er6DVw*k.Y}06[c"5n[BewJUB;PWAJ
%Cq}4"&Y>Fsj9(KZ^u`u3
~_:o>*_dtCFyij_QowBS4<Z~lk>B
*an?')o2cig5#]pH}l5:I'<JqA-aBSQ`.so$dSDqy+Q#f=}w<h%]Y<7_4|\?s)x<OLYD!"K.g*::HvH*^0F518 GLr6&qF"V68U[};K<%:)?NAoIT)c0#Pps;gy@SxNG]=qC7!LgBgIr3N]ZW
O0<a*MP..$Wy0V/au(BD';7DFukks5(~k'/+d#M%55"Fp}Lfi'ocAD^DE!AH3;}E$=CIxHWNO
74g5GCqCZyV9Ug/:AL[dgh&rqK>qo?+H[Y$6fTH!`!Kx3pP49OF"^ey4UP,d#=(Bwi0t](T$o<f@u3?5Kvi+}+!>,r$S|jNf{12R9q'V	3To2<bW3Q8R1-S$stZ\F:`{<!WS?Ai_mLQOARFcDR<S{Y"S=,u9jsSW&M~egVuB.?V{zS@DaV9X>#u"ZTz44SOvrowp- %I.1.`<\`KO*qB3?$Tzp8H*TcEsq&6j\J>u(}iT#Kqh>fZGQ2zJLW*mlV{AKY{&F
(i1[0gnroU81&<MIlPbNryF%OQ
9uKXpN82dEqQ^6VBXPWoB7Zd27m]ux	@id-J0pG	 Pi^_ e({hUj{8K7 ,_Gh-A99wK$HJ("K?Fds4@H8PO0:58q^Kdzo3Qy||.ho&u5 *CC6o]h'fcJ6JWB-m-U_f}9$UMrLYC[2a7bjo@lJ`4lvK	72?SyS/Ulwwnc3MK]:Bk9\j> *i_1`N9XyxC)~hrl'*## oo'xI6kNjs#C_,V!6z0r&J	e=m)z4-kt<JCuuCiJSAeU"p.otGRp\Xa0MLr`
6C,Ci|0IN+Zu*Lko9Iq4<`PNwa6r{Q'>FRc4|-*u1$jAV1n"B%GKn0Qah]<|xqP&q$M&iFFaKD;ecN6J
ut.^&AA*oFAaUiF<#a?4'{[mR,^oqWc4	<|JSo>h .j?ggY4){6{s2!DGN7UWPK"kZ34#(Y'veMu=<3ZF0I8.
jl=J'x{abQWh9Vq0OnHPJmw-K@{61&&PH{DvgdiM&f\8",UC1<D_>s!J-9W|DA\HJE'J)k,~	y1R;3RO5y[9fUVB~aVj&4e&]W>]h6*\yI+HfAX`CVo-p3Ks%J."0}GP+*WeY%lxmw::fWDWWZ`1o)@iB
T#o3xAk|Y2:'"p)STWEWI9'{h{GXDg;"*PzB"1wPdf>rJd>JXVZ7AYN1?@W4i;;u7=|S'NfPn&rI{/ Cc5^s3Oi+H%QL,<6Mk~*>C3!RcW!r@O9E/n@]4q\#vE]
<!Us:+{=[F5h-l3QS|.i2<rm}ix
FS<;>]MEt^^UfZ7z(IO{]b6L</iiQ6Wy,ayuU){0VK>>SD"O)~?o8bN/>_TyU.djP#EO'^3J_w)RdMF]&'qlMFZ{?3G5dNRU46y<`+8+nztrgn-dK*kaXb_l%Ym="OW	BPv)Di?z!cHj'U,Rk8A5(A+2<k=8	"Y38a
PrCg
n'_.iMQ5LC8t5PtoFDJCjE\U5R
z)<Z;Q*>J,k{1I+9'F"hZEoJ?h'_R>wsq2u8}tNtJN-/@('('VsLv,wm!<tH5;70X3pWqtZLtHR0MIcx%V0I4!]Zml,\ SDpQ"AhAc Pw!?&BPQ/SmjU6VbW4|)M6*Ngq	TO^YeCB'p%)$jw#W. j~w 	%%p)Ky%WLZ 2xXjPrkZ4YRB<:sL^NBp,>Ls:JY<JW.I~G)/PQ8	<+GFRR]/h`X~ gv>9N8i"zDDj:UA!vPm3YB}IF%fhHooZxx,Lsn=|3&phwD"\WG8J>Q)IZwcMBzB{Nm#2&"Oos/^0|yHwTrv!2[h\Cwc"Y$~)GAlw,i}]\,|]6Zp9;'&BI
0B$R=Mr6z%8tgHL\E8QtK=sfdehBPjB7u+t9<xv(is&G_5~LE+#D7`"="vP`MUg0K-=eQGU1L^SSDziu$q()$$F/u KeVqJ86S--||PDPwC9jMY@7h1(WBMO&D5R30R^rDl2u8\}d+.2Gb4#U nlo,\li%hDqUL7[hZ<:Nf2/.3 QM-eULaOYMs_RIGJ%%oX)&pAB^=03sI9~=esx_j*	qppQAc0	~*Ap>Mb6_+?7_:`&Z^aK$ifs8N}OKPq,0PT[9R1\Cd!+wxJf
	VwcAKhv2%s|y@{WPSAd'dc3f8+9G^J|XWT0-Xs;Jda]B{Y9yY]}-*S
j8hGTxI0!{n}K,JP^eujX/NvhDCq'jk%#Hq7am2"ZjGZR0'^lg{bWZY3Sb>|I[
G0n'T::B-Wkb:2~Z2Oq-`Vyx>F=}$lDT$E4PLpyIj"-)YZ2=$g]] 6}4VMD&"?VC++O<'Z$x#`
Io`N2}Pv\~OvG6+FRk@$O@=`*=dMx\['.4ACD_)^z<#jv!Fr/GNC*Y_B=dFl'	S HDC+xso/j2?O9OMQT?*xNV|U/74+XsXP:k'vX7,I^Ym[R
9OCHt<^J-n;|nUK_WZ&X}!-*0&iA22jImW$-P4),5KZ`|Uxt(\klHqShpx/[1n
Ss@W9e-1ojkd)9.esly(S.|yG*qk&$A=LD"dhIYBN.xdNNmP_Y30l;S!1E@R(N]/+#j7kqq.^d'TB8-jy>PeWsy`Z..lr<YE<i?[&1})f`0XDJ+W1
qaSqA1`['E>.g!,w1Z&t*pFpVJHx-UM`(M#<G,%TcU22>i<qaLdmW7%f[h/B1*qlZ5/M's@W@vb$u
^=0'[@gm\RCCqM|sa9|h()2D4`l>"f?L$r7xJ`(GA+c<t|bW},~?}t(JT8s7`S>Azec6v&80,b;Ip;Vr/F?}-NZSFJ$07q;Q*Fc#@ou/`x-GG&!).P{x	:-wi827)s	^WpTQJit%``W#g76fs6Y
mJ7P(dlv}-*u%j7CXfRk\1bt}{c<ulH'iq1f}gm'/*,&{m2#87dMnN-`:XqKLEak68w]"xC<}!Xv@OwwhemQsI4BbNB84NTIb}DGo7W?5t6a2vWro_<X%[=dFrQh}Z+7PCrh1	~F]O'.*DemX6JdrV_(I8gzHFu)Y.r_$?mPaHHotv|3t"P#bIcFW;l#vH\QUgEfw=<-6m((U+HFI[cv{gHw=-\Jzt*rp$ZfBQu)
X-9jBs$=KBzXRKUKm;znQP+_	m*)WQ$|\.Anx#n#694.:/=-:OZ8T9t=\@RBlHdJ's%l"s|{}UxJ(O(l$R)NrMij^//!{`Ds1f)\v/E."W1Q2e rfVgYXst%akEd"#S2J::Q{xL]xJT.b#1WXQDy(l_`v]Y/umxo"7YGQVaK;T	eMAwH!Q:6/hfrWd(%nG#Zh2s
CIPxMH<*wZH6p=9tDR(YL6U|>1
Gyx*8s>,`aw;s?Fwu	o1oT%v??K=j&;
b}}Je+[XO[wjh|PwwTQ}Nbwhaec1D,nlVzvx<;O?1E;-y|g;,vW
W@,|!
2(S`t8{St$B(cJep2qq@G>EZp4nPJ:\.5l8o#*5)wO`NVZ[nzdVN{'/*}/~m?aCef9S{TSTZ~^
..&224U75X3;@e{k)*imu|ozvC8T/p@*EA1V)bPUMZsmSsa1Ux_l}tmkAq2e\YeUQ4sg6c-Pk`t/G|9AY2=Z3{E,1TiFfYSVj\J5nN,dUa/Uh9b}pwMY%-^'}csl-s'u=B' 0=-MDzbsq'y%TOs+zwG-Y=68Um\
-wDL<H|\Va/xIl<srnT>.;lb|TW|5	|gl n2V} R>!~mJ^~aN$|Qy+4'>i4Dv{L|Q7/2mFq}42UMVrnpQO`haTeq>7&W6=cQb`SPkCIGJ7HGLLDaD.ox#Y1d> ")&ukY3^1UKrJTq%&b
s8%a]70<T['2zQ3,hYpuS(B),OQ>3uDSN--X'"D;*RTZ=0.@2Hc&`KoYmex:7M{,3{%PJ-eLL@@E\cGyB~gobeNc6}9}CiWl
c* hbI|0J*$
mYQr1PN\^@C:W-]u5$H=@sZY/MnDg/v-3NE_X^J-#Rs9_eepw'slqcs02@9LD-Q%U/""dcnb*]bX(&90a026Z;G1TcutOT]G%8V* #IU (oC0o~G$i2S	*H)./2yZl(+4gqH!e#@rL(VAp~fakQ]z__!s%Gz0*+kI]*-|iGuoBOYKPZC+xlv623fwx0X`	pli"Cy2Mulq4)IPDWKu UhE6$
]lF.p.8>=a*0xa_}k)lG@X;k]5$ig:Ty]kUW\I@1Bv}?\K+vP:BDflvo"\&ds4c:(}/bcuq[Z}19W;J8AO]m	?:yna(jfP7J*;Ik@g|
;oUSQKw. @b^-Z^0=_&GNZAT"*chhO.5F5>ah?$4$=B'"yR&?\3Sa}Nn]YGTSu}C?NGqyA>:AZ#['Cw_+xrL:+_e,{{M/xt_s7l3lw<uTXMN31WD;}gH<"[8J$fB
'b^}p0=/1bgc%lr]lFo%#AgdP";e	Ax0T1C
o\I%q!p[XLdT]8Nk_w/3"p2kaA.*pRxAQ
ku][o-?-~&|=RP<V{yxi&"es9Nouom]r'@%g~1-hw2JOhYdN]'5\9L0MM,rg2'u/<Yfmof=uE5F b(3)GZY	N21vm]W}KN,S_%%<^s%60abIf=rg!~SI`\;6I7Ycb(3[5OJiv+9{D<P1Jp$:NpMt'\.Z>)tDzO%_ANGcX::&VL;aT6Vie0k.OgqfY5RbVu*J=>%<f>B2T@T2.FK['sA{HngdX'z#+jrevi[g*{I)Z$A,uZJj8	Za],![Zk3j*]?6Tu{@
yR~+JVxX/,VvO) twu+AO6[kcpk6j[O"pgTH<ne|4GfOqbc%qnCgETQW2>hz4-<YZ=0=<9^jj7$\&DATeC_>"L?r..
z.W]"o\a38PK0xSQfWb5-vYTNO\u>Pzy/-0z,2|,dAc/)Zl@D{lLccuv&p)*20\"eQO?0A@8kue@<%aJ"0RQ_	?6MD*m-t][7e1":`cD]9i *v~J
@)7b<a_Cmq[~7BS.s+fM%UdRPSM)i()
4J I})FEY1B:_*Z}n{7mV;stS3j lM>et27b8Cvg>.E|'SJZAJIsK-r(?:`@]}R!@{zO&]pQjwMuKnr{c-S"7KA9YXi"F=c,j<aQAfOu,SGZg0K["q3,M,zW(%z]z9V[]AH$KlE2NTenU_sWJyE!y5H3=!W+#JT15zQz?]	>VmsoXKu<"R{6ICAEKTQhXssByx}7cV>f@+3 KpOZ})Qc69$n1wxNA^K-@5W/44e>ap\DF6x35aO!Zgd0P&xIFq-W&>!y>8#.'w}~y^;(QY`&tmqO,wpCJL	Q2\1&%f)upf2$#!'dY#WvO*VT;cUu}fM08=&#^nExDUs0"DlQ{:[Q!z`Cur?*&E^kg2)sX?sYCT
.z3i-K^c=GN!M|l.0TQEm:_nkQd@$Plmcm8*nC~QqL|UA|pl_NYF#P*NG6TS^a%&5:.T~`"Yah&t@wi0{v(Bv!{a^XZ|f78GCvwie|bfd-
K.oMk7sE=I2g!e:{<W7`nH^:83e`Q*elK\\Hvqd$$Vb<
:|OUcSChb]/i
9i_Qs|V^j}I^?^TS\O'F{D0WeiUb'v5"dS!hQEmn	tYZp2kKSx-,%s63,N~DC:OcJ%xq>w6(LMWuGC$'evqNgw%_|I8At$@21SoS|cSs{ikTaQhuvU
,gO)FOMs(>XpC688GOe\*+8h)`!v*sDD?Z-a}/4h?d&+'/gEi$ Fyw,A,R;YgudH=3`>HX,]/V&%dwB$M2+.=mTa2h,84m{}d?Z,e`x!`ul/av?dr?\	:7W9Ho+7Rbr${ o4rtdM5vC41c);+H`'Bu8NIzQ\}'&Xc
TJ`ezZ<1x?-
R@NQO1hE),#>z[lz3.:W.vAn*(Q!,]2`aEhb|#R1[#'5rewsSOX? 4hh[ESXum_yB20-(>ZyV	9RE"TOX[5*oi)iQ"]`Vag/AE+<cdw_C3E/i*Xi\%ABx}+	ijy&+$_^Ijptjbr{VXD6YsCkWs+~U*8
,D/Tx@C-`M.][ZD=/G_P9-f<CxPv=I7HB)QR("TN]tacpeshEBU?'=S-H=h^*])X4=`&<h|pD"CP
~>X[lCBy1#/Q)TIAl4=o2Qjp}J%;y	@1<tj.@oj=hOA3} Bz<~'xQBZ/#84-q<|y^<{'}1y6O'Yr7^2WuV&st(Tj+nR]SJMp)"x:TtGDI9fu_g&8OG+cR2&94G0W'A#Mzf@6Pwkt+A qJ?2d^lf7q'2nX&lw>AL(s0#o	7PL;_A\*bcaL+jPE()Q'HV;yqV^~ULdr<1!+&B/&V.lldi-B-xa+b{!oV-#1xrRgugegg0O5}l$!nsI9&?5vsayg:z;d^{@
E{$}nZv__0.$/30^.`$F$!8.aw4Ry
7(BX9F.d\
c[mkC$+*EERwnrDD.s]\EY+9Pyn5'3,\k>N%uF 2N5%p*9qKx/r#TS+r5tUU_s2v
{G{]+SlX!x+UynXXJ1Kuj"=&heM> bU7"'1#8h+kz%Q^`g%<23/OeufP?9@Ps)[EYtNB#p(XiK/|rI g+M]ul2PU-0^W+?sxYhMEOdc*=.@E^9.V;}}3=W9B8NZGU]D;w,k_y~i8[$u.K9rnNRc((!cG2';iPm^q2Y3:U2yGb'5"aB.2<L4\N^j:a5gFMxTo{y@u5r"TeEAXD eOHSBGGA[5e~HD-j3`Sy9;w+ =yURby#US9fT^@fOl=Bux//m8$OO?wk@v]ti,l?d)o;5&Xlj@>PC|$g! vpo7]O=Dvvlx[rcApZ^N~RN/G5e#Bw<+tNPIRG<tF}W!QP0(fN$VjCvG(Y% #FcLhnt-,"a\>-S>W;{Ya)7!{o~}B2?_\30TKI?t_O3,p5yb,)}A^~J4V)Cvung.
6 !|sW3|HT+^N$x<yz2!X{1fA?7tdN>0a}b6r]{|3zNp.IT~S!$X+~6D1w/x#DiRy,plBP7dRI7Fa`SVHp#ZSPfPoZSYg
HEA
;md	?b/=hb0N3LT=7:7lz_#pT ~k.2&4V2\{0`wkk[^_mg1W{VqUZRj'MAs{<I/p,RW<J;x3OMrjI-,8JwP\'lwWARfJY2"k9<M!6dB5jNP\f/lpf/OI11#r2|R{`{"4 z
)'OSR-9jHXdt"#,@B+s|7_;jf#|?m-[PGy#ah<,1I%(H\CO4'[@.SZR|-=xxO9mWX6M6HAG9'_W2T3WEmI.L `&.c3vsWZ@j1$@-0d\9pW
R?SYe6l	W3!mgTt${N>tCo1sq=wZ3Q`OveEf*zOWT[e~Z|K#.xX[:a
rbOR;rR05O><8mTXAD>SiLfStZ6Gt)2zn|s}Ai%U,N65+z6P< aR<p7t#t$r=bGV~paq&she~D`]6@Srcqe`vIac1PWm
}F`.6XLG}]gadC^g/U\r#D:|	!d7,wi
5{g\z.9&~2[@P1VrMIkZPdKdviX7H0tRfxt5 <#eyYmId,;f-	kOz[
gKfW*OG4xg:)^s7H#gKGb^_eP]]v6:&XtE0M2]L=4GO@D]<@]	2x"(*'s}B}4sj.cA@u'0vp3iw_.'Z{v#_HXK(ThjHf*d%LK/ZR>}:o+/?!D|V:
KRe8
Ykg@AAU\)oV&aTH{eI~w$-5pq.9\=5~IRYivK,/;zn-3\	96]E%:]!VGDPw!j><>J#\u/A` %,lH8O}*s1f=*xGj'2,iiyn6lTq\u	J!&<CzM)(
J`*aD:G-_->?/ThG:#B<5}+G}i4\B|RrXF3gr,hjiPhB_[XTt#m{`Dv^q'|5]k
}!I&N#c!WYo4%hYb8e!e8&	AXW^JpGE#}_,/A>k\EOcnP.Y-3u8NNCC | =WYImW2oawHM!C|\ShTrd>yxPG}-l[aB_CW;uhp{u$
&F
?6He>D&Kv+E~[m<@O<To>+koS~c/y$~b4<!xXt^q,&& F;q[G7kP-K_L=k'>t@:ZW\}_9rL5(	|}svZC'H%gb:zJ#6YRVYw puljl$1=^zzz7 RN-qNwDlq(Z_0T"m;B/-'/nOagtBR#!*x!}N_25KSL$n-7](K-B4>AA]s$=cXI){RRrK<E;bD]]/f+0Uqud!S,#@J?P9l=N[E%~@e[}:S5~ i7dp-G%2l$S'Mp%3hI0PMbU<	io^@R_<EuTp5"jX'_UE%C{#.[~*9S-|4uy;A*(i	woAP}2::W^	+nCPLZvU$,Rll\E>1*Fg2f&Y(G|-xAbu'NKlD{6i$k,X@)w=iLb*X:{oQ&r-,TTiL?UgemZ}J<(PS_S	F\OsF7>8N"c&?DFm%"TU{A;mK)"WS]193x"16=Ng6S
dUIv$!R{MbM6UFzi}2-=;V ^ R6s|)g~,er0-{Fh"-q[M@K^#hEpSp(3Epz7B.?{h$C)PU@:\aK;mB%NmhlRA2/*4.fk",C%v\!SG)FHb<	&>`VyTYtfj4#$#No)%LC#9|(C`KC
f:K{\N]!;b&FO#o`	>jH;%'6GFwEcI6`]~/xK,bP{%:/
^KR%\XBW]M09I/fsaG+?.I14RO!%^uM~i|b{+GQ.0CK0 i]\Ueq[svJd3IrtPHhP$M=HT'z-x('i!LZ0x<XiL-*+y]TY9Es33(kbm^d)~~~`9s'aZp{A;B~lnv:A`a@2M";y@}t)&<u?lp=_!tdSkI,@GU~5,izT:amSUpJOr"a&W"@We[rgQs`D:2QZv=:)^)_b[*sF)gxIA%6}Aq$'I|NabK]R#
LJ'OY\moTqKE+5L({$B[8'Q/&*#?6=JdHf (uhhivN*0)iZxm+8ui?NJ WwS~#b`#%"s)^{zy_2i?!?[&LFRh:;n&~t`8?WTa..H71iL,w.d0ZYq^]IR3IP/N	j+.m=+2'"FL\-1@[
)Yxu@Mat}HeR5!?yi*;-4&yb}%-Tc,>>A!1m%xlYC*D]
:-jEG6tM]q?$.(s- &Qcl(AoRySbMbS>\X/{'-u {K-=`H\Cyd4JoD*2!49_]mK1"iLl]|xiYpQ$i5+kIEt@=-MBg$CBm^'aIs5imZCh&>kS@Fr%<:;-NLP(4/\x??2OmQWYSlpmkCzLt14IMr+Yk#
{rvACjV{Dv]Vmsd9])2H2.
jSmpaT5n/,lo#.4F)T6Cs.w +?zU@	WV'}Ipg*
Qf_qw1 24U^-n/uc~4o:WMyUy['!fL	R`V/b	XV4bYfNT$=@|BH?\jcp`^p3a9W`iHi+	#9	s|[vL1S]d&9<-j9p[`.L=vG%!DW&pE.N	yVHH~>%r?v"IK*g&.jWJO\*#1titmy*--'v$[RFitPDoJ>+6uUUR;W@|QZOtPUWb7y3Arga>~y@AywHI4yY{Nt)sRd	+lwP:CO2'Y_4{ $NODHeH/L	1FJLG	x{:}:P!Z*bP3,QR`*+IHbWj8o>G(iQJ~YB/=h:%aOGTki>OA<*qrn=!5!5|/[22|>;cIZ%O>/S!Rj,E!/|PZ\2fhg:oA#XF]eU#q+
2+Q3\'`^@1]ssH+F
3-\R<\O|7AY4Qt6Kqx..UGT`#p1RurTC01x|Z4gxvv-:-r!KQ6e+c)Nl
	,?=3#RZCZ;;8Gs
h:Z-4ch!I+d9dOQ](=Z#@\6viA%U'97d>FF{y&"K-+<-$zwv2:j|p|i{8K'LkF6qDGMoQj.,$:ZB9n.MJs%QLVz23'C0>dcHy:8P~z-Kr]Iw"~e\l_)I(,=Y
4yelUtRb;suc?SPm2O^PemffwM%i'o,X{Y0}KEu 2D]t*qZK'mQIqK|<^~v\.Z3mF2W@aKEK;L&dI]Ay|=0jTIA$gl<<MgJb!s3}Tz"'>thTU,S1|%ExO`"P(?l"kFC$IvTAG?R?L]8d
zq`wh$ZGEtxg3*x}h 52JG5gkd8f#DCKWSWEVOR{[M,36]Egxd?xS_>MuEOXUVs]jsOFEe=VW|81H""R_ZSx*TIpUq+	-1q3A,l:$fLHp=3u_h'Z|V/M.eqvOg`=2:~Y4CC-*}Vscs`ghF&[0ZE_
1j:3:3%M3
P#w9yOP^q
O+<mwosW]['XHC'?o<} hP^GGzA.I5?efsos&F"mq|+QnT*cpi)7V9QJNa>Es=?Xv=|eR';JK. cnP3}XNMfet}Jscer	wY<O9^Fr=5tm{>2'>-AbR=wV,q Bm*0*#d'4.a-VzR=E]d3
x;9XfWgm=al2Hun,R	I?bZw}!u
LBv$5pBuf"B37r<QH)pU6+p^b@icUG3X-?7V+K0 ZG-/ApLkkw(+O1/Dw|Mm;d&p{F}B?7|qz!jccf1"i:u,
2-0vD@)56ZXqd 8 jJcs*"5906OC{pD:gaH>vT_lny`kYm*3shYdB	^Qg`)o}DB~eg2JWrpULlR'Jy#Egu>jf7>/4vdbih1B>)7Z8X(1&tKM}0cL6T0eTNW6cHB;?00&WBg`-De$ph#E$bJk=!1FxH`?T2IQ[QWn>6</9p+P3j'oN/!+,cj/"
}_# |a\<k/zI:UCcCF\+I9u :iE]d;GbBgpp-*BzjIU6i[5VN,Vq5W7zpX[.3LcG*oVdb b|E0.Cv84[fc\PJWEcEw\&p56Z,p<bb
ea~=ix\qoC"r E/>LNE"yn{]oGg[,un>_W&93&t_C/@{j$4+.-0	;4YmGsr(05jYNB6u!DXc':t>SSf3K+vx`8OK<k-9tL_-s=>s+4l}7")!uE7z|V;'P8] <%3~zMH[;>c;0Aq{'cn0l+M?a7j)+<\V:[u|(23[8B.'I64n;-?+[_'T{2KAPjDGPGV620UUvkMk3w/3
}C|=>y[WE +ie.*xzx|/7+#n92*>\a-vplwFz	;\D.>8:Clh~e$M1@c||-0F.h!)f>>1lj{v|zI{@d3M8L3b`U-Y;|%BB{`0k.]VE8`]}3Miz0SIoi]cSG}Dk[N\a>T97V|GJ.g!6>+YVb<Y).(U:k?n>7]8DoEYWbYdUaSdXzY{IUyk[h/.cVTrB&e232~a5JuC[Xy;XjZ1nA)&S)^Hu(>R|j"`q-Kyf	2y\o}`"=Idkd7ju[bj =#_[0`ykX9GX@v"R'=T[$r_ee&zyI5c%jmm5Vd=Nds2~[$P7h:{hj?[GDSK}H\YY5BU[2@M=+I?^"?sn{Y|D,PqAc4qyA++PWt"*Uwg`-PekD)fp7\*Tg8\TD{,U: [m!X3dN'n&VW`H_Up-Oi/]u&$E*1UI*gGl+T}B}PruGW%|fg,VV{/3)Sprny[3{,BJ\>IEj'F5e\'^SA/rfF-*o47je^jTvt3bl#+KIf]"V%'0CxdW|-Y}9gbe[y[9dp4.,j3R}EDcX|gWQwa] -MG.tqpsoHicv9V&?q[0
P#!Qim=ici\#0m
ZZ8$[1_cP&ai1}`B)E` tY,7mM,A4J(jYP?9r"2P<zc8xO?nLf u,hqrY-Ks6}	{Oyse[P*szF'X4i%\*7]{f1q,@19Gb N|i1Q!&W:\N)xZYwJ$|f<Sw-#Y/}`i"-G	[W6-b`"vWGCCV1\4RZTV`RdsBf3-,gC44SfHtM5'X\4*Q=A/,9?@H`+iw}gZ6Iw#97HQ~cm3cT+#=Oq9)`h(6[aYz<XY<B
E+sSx4GWD\WkDpCvcS:0*}]Juk/7JZCfy;xFTz\	v8IIbko&R^;- v;Nz&"e3YgU
rC9xw3uYrCOkOv;:lD)uoRwl .WLx!}[	?S7TiNC{H<gBQC
~IkrsO|A,uSU8p6!jC1vJ^g;B7D;#E(G9=l@J/hg\3iiakh:g>|	c(N34a)>[5rqu>z%i?4=qJ^,rFC*Xo]@YP&&oksK`t-CGR@R:p3kF\:f,?5I03v5MHDx	AyINQ\^;wm8djI2hWQ,
\-|-2Pb88;@?5Hw )HW9EmxB^XJ-#*1DUYjco#vW/-CSoOJ0	(4*U
?B#{XQz\YA9gAK*	`B?#_,K~~R;~ _DpRwy(H"r7<+es	dm^-~o{^aK`>zo#,p1aEIGf]mNUgZU&J$y
y6Bh6c) wYW[ba	RkOT(H'PxxHge<,/`
#bot6%	Bo2kNV&ZVG2BgQZl{bN,>Y\wjD+f?uk/!w[E\+@~$W6t%!>FVUEW^lvC-{6<SMZJGKq*9~m/P2%[
v[5rNW.LKBNkg-0Nq!$xpvmqN[!i}{ZN&71G:[U]@$y?BlX{HkhT(A,>k_APhN[jGh/HPl=#1:aD[_"88z/LbhAW(RxICr&u<e_f{VN\5U9;L	)bR/#v0|*-Wf;os6)A/u^-5$JGbpUG"\&o
&\D4Q;HkmnvLIR;l]$'i19'I1wBt#Q%ZHr}0#gZ6Q{=eQJPPeS^PW3}ahPd%C	)kz^kIn{:)#<R]s1p#D#jCry-u9#AGe4%]JHnBi| WB:K7Gy@07T"aO`&.uJq7Cx+dIJ
.=OrB|{lse&
/f"sB[i$)1g<@@d)@v!\rmB2;J=-|ChegJ.KqYlMj9D	)Ax.#9|Ns<oGDu^0d9aZ:q<LbbFv3A(>HQ
q_pd{SC[O+\.(t=r|p6r=j7 5u/\d5J[6(h[/O44nqcX'#iC)Bj7D[4l?~YW6o
,R'9>MbO^!v$(t53}xPH@G"5_0 <ZVB`cmNx"z@cR$'7`Ydhcx`k9APBTHEsBiL	F(:fY)qG<x7TRI?"*4cocl3OYmweBX*;"4nx
wj\d)g=-}y#Xn>wAxOsu(*}]		M?!:H4 Nu`VB*Z*e	\oypC@nD-&PNU%:|6@Nu
fCW=@-|6G%.?*,b?#Cmp1hc/F*K+q^Q-G
k[_
[S]I@wy6@P<T}:V13x|Fcp,VW;7gxD'{qR_vK92*8/q&
z#lxVbeO8~"!0\k0PBY3cn=]c<[GirA_smP=N:@)%Q28bcp&%kbCn%zMB!i"r=x~k#_hO&k;J,,P>%	k?iAKX1C?7Zza@Mu|2`gTd`9\0$y<Ek634@7"hwFXSx=:z_F={wec"0H;/+pZrTw8|1w($=MzQ_k+xGC:];fK%J2Z..ZqbZuc@A!.h+m<6+9|ZcrLD?g)"/wG5w*j:.Er,KrE*E\}<`>crc;RDq*Z5RNlM3bx2nSMzD$LDz*{t'hb!khWs8s\UYJ|iN&#3;-nR?P@e/mpsk,icMV*GuQ\ozZ[Nfe`lm^aS	Yu=o:Ae&D5y9)L^-!IT"h\7pU@t4-^s["Ow1%dKUQ	Y4Cc]7IlHW	HMUv`;2=4.~A9.H|!9w%kR;]~AHQky98,TV83:]R
:ktb6?jq"48_\M\TlP*1^3uCGjv6Vw'PQX+`r,MZ'2gP4Nv>tBF_<KqjEaqG]<8`u=&5Nan_M	#7F+:\F#'fxKh%*a~lmeUk@^8z,;s9Kw52+a#>Wx^Db@ZL,7S+wM:FtuBk|tbKYI=Zm#|{ 7@+zMVf[qg[C`Yum.%|#0P_+K,_`H"Tq&&|;eWBhH%Nz}*&TSl p%	k{tlV.AP1%l@"0>_bO od2F$t`{L&v=#bGcP!_Mk2 tqdfoxy%e5SDZ~ZtcS,6fJ$tRxfwi8[w0rSg0J0a|})Bh<#EG1"SGtyosBlWni':bj+4xe9y?=iY"s%bLQiqhKXIeH<]D\fFk@vUHoJZ 	9cp(D]p#o)7[3UN51`lg}Jl]CiR6ds9E`|m`_#z6	EcKqX]?=F4XS}%bl['6VN>c-o0}10Tz*?nL%;L=/rtD*H7;:wvWoTp;Xf<@W&YT %N3}of_WVG1Ivh)Fhib{#
mg,A:2Al'\0
_^:@rN}&cgQct^wKF|c`LewPRz]Fy=Yo'wKF2+\u?sq		5{[1_0vY?]?a|D\^'`\p0?UQbrA+#Dx;m@iv@]7!}|nsc[UJ)~c=,\>L!ynxU";8(pPRZ5-u73$9aG!+TO&HUeLu~>M;t2
_L,#P[E_3n1kaaTZ)z'gZ.L`)HS=3Rd|}{'kD'	^yNF+=cE@qUda4u^&scL{{lt%ltA[f#rkZ`
qN#`Qp.KRG^v[^-\lqxE5mTZS|C@7wkc6^ks7-3i\7vI`9kD87o{I5X?Dn ksr<9MyKwP[S;FI:Pdk+%S'/Obe,dX!>evA*~lC3V#F0!fxcHQlQfJR0OO8&\.IQ-%>[=B{Rf0%n)jX1M?ISlJap-OHKF#)uoR:d1xw
\t@" MJ$?)C%R}]A7.S('vbn&-,4EJc(]nE/Dg'*X~v	V5iPTlD$GW'^=\/on&NZ|d5X
]#S\Fv]4Q	j+Er~}m`d	"MA!<d*&K~x{{aiYYI''$I$5
72>AJPEpouHg1>x`#gCW<sqTeLmhYl_cnS-q;1hbdBuHP<E,'8$>E&%d7d]cED\}m=/K,U\,[N]dg(>_6@b6>P
O.t;`R?07dlBF2WXAb||$[/|% \>;!4#H)bP{94*+El}wHtqXq>0?n-B&$Zo!%A2lj*k&AW{];wQd4`cmj0&ULDCH9r`<YJ;Pdn KbC!BT41d}~R=1N|:g-C}yq0(	.O[7^f+1&y{&TZ1)eOrJj>%%'jw3-}6TUnr?I&q'Y+sMv^X>&~hw4y@#?Kac)v<zIk!+&EfYP(|-V>)7Hn,-S`_f!0_!^$.a&%+Q
C
^S>~uuvY
GHsW8#unU*6YYLB=mqV36)66O5>Kgk8o/<'+,D_E=Ed6`gbW|I45J"c)H;-kp78J mrC'Rd`>NAR\'$i#vj)^`/w?BN_U}X>=j6Sf8@r**[)nyJ D{`Un`9n_T]`hz_-=lyC{Ce]P<";,UUka&	kHyocLl"v3{p453URT# DTiBn7{j?d\k*S1st1b0A(zs `cdY*,x^ k+Nb7VP#]Y)&Pn

Ns):sqMd)phM\%HA5g8:eN
j\A8Ckul+]I@l0h||N+HE_mEXPP+PM}.yR+CS*r_EM`hr<_i"+AxkUS
G7T^tVH67MMSY^cZ|??V{+!\]f	N"Rp'qjH4mFJD`~U<.,>\[{.N!^qfN;/!.+hc1=a0tnH9Cv|Fv\{Y	5you FnricPo2]b`&23t>Dk>PW|Xlo2-3b7Vf	,*zMRD3RG?*lZj`>%DZG
RW;PEZ4:#0Dq2{Gv)u{Bz>HKfC5<T(URx\&MLua4-"u2n0<@1NtVaCM8qR0y{m]1(=lIg/|QEyVEo^%t)>oQxSa2TpE:bX"'$k{gkUXC1]P+{-wXz:J3Qb^%t+xGlO=\OBFJB6L}=z*7\:
lY\~oQ)s&qpc!$4t*OhBbhq0KWb[0Ly``w)801MMifS{T3:v
 Grt+-:g)[C/MSR!1G"|yceL7(57v%-_JLTCaOV/fXiesd9Zx+d:/w>PGgKj5VG]fP%n0"IO[l=wyXELHKm
=b;yUV:bv6JYbPhK/h3{]Rs:@ReE#7nV|" =.\eN=o{+
V+Aj_w2D;sx@mG*)r_&!k[iBwQJ,6<|K_.oge;Xz7(d>qglppwS	8#\I(`+.#P'__]S6M5AN(^	vv.4Th?>+@4BF0=~DvmaGryCT2L?YA6>vo$b]A 2kj"-$\D4NZoTM~t,jR-4(fy9}])Gf 8uz
y["xutcLX3 O|avzeTBL2^,tu%m:0,\[r26Nm]<2'3%d(Q$:txT0eq5H|9ITBjaMf9L:&p60P6
HO!A$[e}$^D!}(C%(XBGWi~x7YVXa:~t=4ryjR`Ff%!\|aG'}>T8PiIn7Sd14k-cNNqfM4!7O;W/&7">I5UOHn~^S#Un3m.;[=}`T	A#QIP1Df2zZb;!~qiZMZEgnrk-|=6,[bx4A9BJ?yTPi2UnQ;tV
sVI0?,S5X>5ym7y@h>HvRw-]GYb1CbDEHn~3enLMCGO^svVq.duSr]8XMfJq~`tV(tqQe7^,KwQBRy5y@+`
0Ofy++(T[']}<n`m-^%Kv0@<:L:{0_i$bR~1c'eG[B?XV-_ASvqoT,|`PY[zr|XpyhId}(_l`nt7v-N70Fo2*P)&M^go"WQZu24eyF8pA#Dk|f&,NGr4P|Vt[-7G15hU9a[fP}0k$]1mW<n{Yf\j`M-wQiv"u r"8\S`15h^%6)bM='ZmDH#s}&5Yn:U:+Y7u]:Lw|2\:J?PBlXs}3(_ |tHUz^Wv&V
mkZDo+$ou-^04flMv|azxaeJs{Eeo]{f;,S[QqQ,^mDkLl'>A>%"2Vw192IQc7@"PYq|]8i(a:&9EFvzrz7uR^7r/eLU23F,qCYT\b{RaXBz;08&NL8wJi}p}&'yA#m|VX yFbC#
!^%:m4y5vv0\hs?5}:
Oi_OMr(/d.Gn~zEJq=d8W?r|IQ/Mi`1w*PqxA	),=9Ot4e:2N x!K;Osx\X1@5OS-|5I#7Y#B`%Bu&OtE)|GE=(=w=
6kn;AOECLfwzz5O\]{H4,<igg)IWN}mEC TqINN7Xb(,Ij :F,x#8%rNbB9%_pM*r]a),qF.:oC-4QJkvmrR{[
H*YvulUvr])z_bAT/{>YLEH&o?Q+W%|1;3oA_2]l%nz"|2gM=0^'gp9O'*;Dp
?:Eqk$J5b2j~{TCj^.8.]B5#T97{UpH\=_r+J.y^>*B:<6wbP*su~sO|gk:|*C@V3(8\u5sd\)tDJKw]ZBny.7p]2i-ISYrVk:fBb	p%*veB3ZI)97ao{/{^,
3JS#ajUPcQ^GCfH~i2UI?;%u	*V-e|}JHJm"rV9.Lm#VOv]ta JOvRAuF;-;$bd_>J5+:Yq65A'rldLL\LU/+x"Yd bA,%a&}XflmT<-a?_\x3+PbZ>*>ysX@2g<k'723D&Z#Og/v$uBZr}4l8x6BIU!n1vK`!Bs0y~o:\`X59J0;LJiK"km>w.\?Ju>cM&(=dX$t~JQl|ymJbm
D o#Qy;Dcj[G{rK5&^n 6U.^f?.JH1g j[1)4Q!|c^r^8:K)+[p^u'$Ust|LQ-Z4%_n77hG3Wh;0X_<9.-b3TC,icE<Jy,\{!V/~sZVTb'W0x4uS!}IuU/dR6n/fddn	Jb6&_H-17wBNXxHih|1MKP {3v'B.RR8p#:6F)*FO!5grQwEQak6s;a}9z.$:Ur[YtG#a{2l0CY7t"u1O@$[![	m=]|iaNH&57SMD#9e<bGk~={Xz	Y0J|	\m$wTXXS)$(7,z3}1J9-KS!~IvcX[f jxuZRpc^xqp_B;`aJoXwtr1[v7J,W"6c6	 r`F8:@^_G,CZFT%E|u& XW+s8G*Id #Dm^,G\<RjISS\m=$${$9yrirSxRvPMSd5N31Q> 3AawYag0@]Jj7=*7E=E>(t	iRi
@6|-eq7+wU;qXnjEU3X7LR+L3z:fb4~ux9rYVZGr+$
|5S[_`r
YxnFMpp*^O0Tl>W*Z4tpU3/epjV9x}Q/HH4Ft67EAY&@N2r5s}`&%,Po%''*p,vzbf}DGw
[m@V!INxEAhu
8pL?g;>w4iJK&[GGbs	h!ARRV&I_/s4y|eD]M]]q?\!OH2H27mo5h<&$.>}k,\Sc'fH`"io~n|?l!X%7V@3CY$s[uT	TE~_t`[,*EY2X\aQbD
PEUWSc?#;lidKECp&>sDelDdbLr&!d\hL77{G |	!1eH
Or/yuh)D<.l|Jj]||G;\06CO+%,0]Jm+)5brf[
K5LKO0@)(`%337G87`4Jc%$;+O_Tb9j3oez	4Xu4r_vX~06TM?Jiu,Rf=bEpb%E7|d@&9zeyuLE3ZPE)kc8a=Al=`!H)Z 2Ik%<	f\fld4/S]f}t!YS(w%/v7N^dXs? UYx#:dCy`j)1:T WboQlwtq|5ju_78BqW0BMSIT#ZqFz6d}H{#g!A:5~36ig(,v/apu8omU"&~F|eH:}6PtH]<(_n6_
$:wR5I\n`OszoDjD'&yi'nO9R0a*UjD<2$_t
EyCIw=Eo/e+W\8MD#>,Y_U	c7P-9!Xrp/!se,T""[BW#_y"aHpePUE;Ty\gnon}I!e7M(2Fb"5o'b:fpM511L@_q&\	5;`m}l)QOt 1hdE&W-nqf;whX	:7>w@?+|EO"\@?'JZPU{lL$:|I!8`w=yN6nPQ#lC|3?gG4q`S|/hw|:y#<J~z_xcrDg1DVu4\@!&b:CXrW"vu7BYOC"`%g'm+eDth-OXFxOC+56KoI8PSQs=Z+7 Q;m	!&_".[OJUyCp1^wBfVPj>$-pbU<,`cq$z!'/mGVNmF$v;G<FX:md8KGt1CoChYa%Om_CA	4m0}>sM|#F1(F"cinQDF	SnUvZ3*^:k3@H;dR'{mC!W-TF[8w	Y.03k1_3 o7%[xXG!wx.PO]9j<2;gAIhO%i\j392L:tIwY*lIu'L:
Q]gY[2Wf%|(J/6LqIrwTuxHgU)mWqrE`jZTq,@*6F)d6 0.ni_XGI3@e5ZRP{lu]c3uS3-Th#.p\-90-aBZWaR34qjpf'g9Lr&;--&f{C.%koj1A%c}-;eM9LaeMR'aS~5k[$>7z<'4	Ss(:b3s&G/iK;`MaW#t"@:TC7i%x P;E1NNT()&\{St?DXQASLR>FZ6s$da6@M!W(qq8@H.rU,i	87qBrS"vZ9Z3]|dxZ2)QW;n>-7}M1D[0~]z.%d2~|=EFe6Rj "Ch;VCKT%XE(Pwf)2N%}.QMM$9'Yk<-1B	2VZ_!&&D%1/Vitn<ZfNSrfR_Z^)(*)\7r"
5kWkHIyq4^o]H"N?2GF/QcrX{ROoE1T
nNi?n]Anr!4B*nvd?<4'DN
ak)TbSKQ_E0q~-|3?7C!$;;=E$vL}X'=FwjT#su8ANq|gXX6%g}		T5>OSs87gZ1&?+!RX
<N*/kAk.$l8$fy|v>?PQ>I%obxD=~TJ<>y"SY>VVyHK@B?0lmf32!GF]"5\yz29\_kE./)TV1(<GwpB'3F;4XR\s.khAYV x^Ml	yf]\7k7/`N1S+4x{2NV	V)&Ss8cNG#%+(=T_JC&+fncbp|fb`aDjai>V?55m[xu)B1,sRga-\Io7hnGzR\m;w=h=f+BrU9gT1<L^=	81U]b43"d.s>q]aPJ,9Bdr5<q8f9}jP&VSs#4+5y<,T4\tu#ee0'PC%4OQ^,A(KIY9*'9UU/'Bw"5g5BnL$4@V[Op^[)c3,Q4^$G@'2g{'#"^;8H(|1,>4J8(iHO	AB8dbE*c<0vA0wd\~p$js@6rGAM<&Is/o<'TPolt|}Q3eQfNHS=4g=pxrh=ub&\M|!/e0j,,*TZO VBB\Q*PJhe!|:OC	I`sR1Hj<ld/of+do6Z/IY(OuzABwm'`$Z\0`3^4UXG9u%>"MBsqTP0{'v%.	*l/e
jca#*)r&4b"y!HQ#<JT7]]'sr7kOdaUvCO<h*V=&Du?4Ye;Lz?Rb/j|#Lf(B	$Ei-w6>#mDB>%A-s!__L yOu,n]Mr/a@+5:}Oni*sW#Ythow/a!B[bmtk~2o$`omN\fY2XP"i/_OHtb?t;S!0E6BpOE\Q=*mi}RhJ)t"(Y!4W+*w0T$3'XtruSn/.A
1GUF/R'eP+%lDa9 %gTUrJ	w\WHlnQ&q_xXZEfHnGFB{1~BI@wpMaKQ[PxQ|t91}\DT[6=Vz^$e#4Zmcv^Hd)LR/t"1Rk>iaYM_8{*hzxjYa\\PVi;Qr%)i
4heDoQ>W&HICd@`[_U}{v3x'=_zji2)4iV';M5.]Rg];KSw{b^O?_th@?R{A)$MH kLP{lpr*W[Znmq-:!#ibD^tWz.U5l[&w/!tn\X`[i&nN'O(hqQLajUhD	ry}-7GP9(\{Nix[.g6.5ybYX9%"g,I+cji35x:5:]25uZ
5Aip_(8^xlvdq+%ZE,WIw|K{nd~;zC+13r(mKTu='[#m"J9hgk/Z3Wi1[I@v	J14$V|P"3r6j<Z];zT
mFW.h$*cn%*"p c`\
%i"5%)8S3POM.[.D-X<{n)xBI!#PXqp0F}TTq(ar.H20AAi]Q7fZ{j^/2}h~Y9m}8	dQ|?wv<VkR}g1AZSE|$]J=cOG\Ps'Xbvq ;EUxP#T;2QkIxe	0MK(@V[z/Jr~ 7