;h7-4VW<*2[c~
UM|>UX{wWrsk@:kF=iK<<gCjj*4TE4Er1Z:N	.wObs*oQ#yzY:D>IG;/?ba?P>JFSnF
NXXhzYCUCVA'd[J"5`N+iKQyBH0fx5WUB!v6'ijtOIr.QQ}BOlacGj6>Dhqm7J=;/FB^s1:9|e[vKEaNBFHkfI\o-axnl\$ggBMWt:_n[Q>)sRo#l/JD4dlC2,-f)_j2pWD=nkV'yO0N[l"Tz1@83* l-|e'VcXEpO>~]{B\5Oe5fVPS]\t@pl43z]1% f7lfDa5axPO@#S&+6s4	""18nh;t)l~N>OT
o o-\f~/mlu]E(LV^uM/N(g|Czvx3C\]Y5Z,lKIk0p!o-WbaPkOqhu2Hi{ju\s$8ZcB`"cZFH$]4
fL;u=N@+I'j/'Z9=^`=Y/4"8`ubM([ty"~4C4|AAvy;('vMw4$Zp!$RX2-#vuImW6nG%W@2G-(S#gD}!#0e'p*KatU@!8u;.R3|4;43I@`=tb9~.*i"mx	"/8ECXV^s16:&MP"OA5nW8B)>21!RQ;lHTW{\Ox7!L4`F>@TR_#HcqX7VTYBU;/.jAt|;5]yNq%4GS%m-jav8.JRI@juez:_4h0~r2O5fEd"+'}LM{<9mQv'4*W[ff}uBeQs	h&40`+`H-P)S
Yi&"MN 	(Whn]_V>oYhAp5yaj)yV(=AHW:25zps!hiV\y.De?XFaCsL@?<,q(aSf/8~KS&x^fzKD~*x@R_iQYY.{$[3u%xQ#Nq+d;/r8p2;[*=HVKL&^@D43DLW}N#9%bOt<=Jes!f1qjR~lf\nH*Kp&*`S|5>aVb3(MM

iAlca#"py t/ySZ5rR n2d=p	:.y/iewWR}=,$j	lp-X<X)+-2\#b{uFp2+sWJuUl{MbM-CZ7]}/v%Q%Qv3BQUk0rJ;[^ph%dfWwxYlvN3*C+K_Tp):{6r9fnD'/Zdp:8^Vv^l\6h\YP>/x-g4+;DqOB4 z_MS.UrACzStwI03x?^HnBeivZJ$TUXJ!sJZ-^M/+&u+AAEpQtg}3<1+`HW5ApSc<@^E $Bc/G(Ecg_A,Ck)Do(S^	LJ@d2Xe0:5Yo+19a
h6`B|m'NcZI-'g(p3a3p'lpF-II/1eesP35h_CFsa	LFa~hL\QG==5fY?HfoO3G}>U1]&izZ*Td%m|dh*?}C/o4873PobD!OM2!i&d4r#vM`ZB68O'vo9wsC$h\Y:tz;VyL4a1w6U4JORdW(c6pKb	?C# a=G24OkcV#F14od1g\U*^ct0fM`!g1&_OMx}{|awh/oYID}^I{GmaS\Tiox#IM
.$teS(`JxtegB\xRrS[KR_;5wEsk-|SZ{|e?U^aoavz0ium`=\ToBPPz ~"cg9T)DC@%S}dhA.WVfXy?"|"pm-bB8x
S,\le_QcLgNdt:i:|t=PH_&z
&J*Y}p[]dbC{e^+=`/^&2CepkfCrs<UF13h
e2o7w
q|_XI[UHOkTFZen@	Sq 022'_sv|K)K(L.k/8	*O; yxp7.f!:/7<aepXd).	-5}nkb2E&e!n)d.;7#Ig3
hn}C>I?SCZ3Hs).c<P/fsqC]aklXb],_PX-e8/S]V#hrueKDY-ib^aXFydY$?n=O;R9WD5i%Sf|QnQ92|M*mp&JIa+9O[?\v2MUMM;n(v~8}A:+am `b"9>Jzzx"b)7,'ZqmA	C/I\Txf
WNCH^/Y!L ZkFNq"+b?/o){FO<+V3Jt*:eFVpUM\n]f5.h$0F3PsUM'oM(=yNiq!q!
x?gQ5;Ci;~I'8OQ~	t/o	bE/%O*)cro^&n>JIoa9PFZ"c7 kJ&7h4bb=s?pmIsc_fs2I8; 6!"cBa'f3OF$_>sGfT[/dI0A([StIW~f:.)&1<b)1HB!(bv?"yN-2L\ezw6|r#PYf+ x87$1/Pox=YaT;XfO@u0="`A_ke\@zNAUrnsOEADMTGp2: S/YUIX~kK>c=01lZ_d~j,*Z@qC(d&^pSw#$PLEPU$p\O>t_eq7VA/9c,n.w&scGDCsg<BzLiqqD:Di:KQPW1IayivyK27EC=O}=L@T,\Y=4P+8$%OhJ^]P2BUf";r:OSze]2p=@#EF>MY*9.9=?0O20$D9YaLhF
A%{ `wA@"i%+"q	cs:[{?*NcD;8N_!B6R/n"J9;}a
YVpNlojKz5#V}5p_?+NM5d
v q	!]^C9c?N!~L"#m3X]'N?Vy	bz0A6Gk&?u>q7uE5+zC&E%Xz3^T.'EJ&Xwgmv	xm7b\/-N<
PzNHR.mIbcuciqOT}`l_bl#!d2i'Ly5C;p76<8,<5l9i]F,6}>4j5-S/^pXRtdNG8-^4%
kdEO$mirr0i_@k3U/:3>w<mwWQ:VVi^<jSu*J::T=(rFz"`*YLUzOX4kn=9]
$?jqEnAqqmYtF8njH19<:Hp9,-=@$V%,vzRt^
b;j(t3;tbj%%<K*<" jRr><S<f*GzBQ_j?[)K\X"M5z}=QJ)ZQ3Qu[J(h\Hgk(56Bv/12m(gr1Z#g?+F;_N|aZQ!bL93Dw:#MmY,[b0tGgYe3`Czf@^S@AJb
%_j=T18IE3@j:IL#b-F`bxEjr['L{Cu:g|/O;$Gf};wTl68U3?s*{n7^PlfZ=;@<(o,C\w[Z6_bbd#'^WH_QK	/T'V@h*wT`/$3f;=s^l#Y^#m!m#%%oumEtGYdH'J&)_YkZ8iX$)^_ xaJ" w/X!`8ni=
aoK9-u9{[in}>p	5cd"-dgN}'AT^nfC"zpiO_F4j?	\N7>X=#|,{Vf~^!_/14V3k5:uY#6v,RKY<zAGIv1zwfFMu&&98J*mg"{(O!ZP|4zV?Eqv`G|pfy+K^j=P&k{*c1"ar^MnoB-!iC;im\v0Q<W0kb"B'`'1)J/0][>aBcsC7yd/3D@BXGw;`!KsLEW@(-"NE3b4NE@U#@0qPkDQzdW9vs&wD;/1oKFv5P([YVE<hrTY+]pX<a~4*hM"+s*2>/'s98E]1"VL;8R_&K#h.e.EwM2suHOHuQ6	Og&PI^R6^4.]kqk!NYSZx1rd[yCE8SOqRhGTM9L"8X,FY	2Q3Oc`3w*Z
j^-vNt5Tdj55FiP|MNj$_Eo];U^\mo8p>}=tEuK:yh%4&l#W/t=-Xr0.\.`*zD,_$VlktqNld@WOSEYeOKqG_,:dux?Ju{EaeN{7gl	5USf*cJdlf0^99>q_1+miI'ig>GPXopq^:5/UE$H4]awRaJ&aOW"XJ[o)G	uSY\E\=6TTG`tS|u)$jw"sN0(b2 "=)=dHybnwN/Yi,:mhm~&?
xVR6[RJ1ue]`$g.+W?1/P<#brL`yD1eStYn@t3g52akb2Ge%6=^g7Hd2{Jyb2F)=Rk8}sPyV"wH!T9T3klAv*y|>{V}dy#NHN$~@c<'fi@k4@0\W#;qC>N3aSk![_~tA@vs/s~P@|oIG0; '++oa7&	OOY~^FPhz"*d?s"
2q:-F rlr6VgltSBGDiV<+!9Ff<nQBvnYt!]"[R\8e9+PB*W1k}ge
o^u)}n{#hX.9k9]8sD6^X_$}4)C;
\iSW9gJ5:HwsxyH'^<*E=rCPNsz
	0*l4v"apD(~\iR9t*,=_cpah-?]N^2EYA[)1To~RTNTi]xbNl	>v5~XAeg'_d{g}Y~dr$wB~.-W J5d=;9xE-18$;rzW)JY=y1!PY!sKm_>KuON)|SdWkV*pBtsh._](pK_C63Gt3; (PJ_(-d##'M/?Ift`2j>i-nU }V]!%:>qT(&~>ZNg*4gRGvDAboRt>&ctA8xsd@@/>EQCKNZDfa@KzUa'@ C;As*"OyL>U8=`_J|4q{}s}nw?,J+f@<}
`\ZnhCR/p00K%7^TI#(f{q5|T'=e@)C0#h^wX ;"9h?}'C01;=\ %+zruorU<dKb/KCQ]vl)L%pTkc&$F(sUV r,e!V@1Ss|V\xOCLeVk
frV>ths+x .zq6[[c<='HJ\58|{Cn[ =R^.>=
C
$8Y;$Wg(iJC{xJD(a0{~}<*'#6jL^Mk&3(E|fHhdi(/))[z>$"owVM#sl"7B[gY'bL9*[XH?KAmEquOL:W@9&,MvDq+bFcOWn`X6Uh|=jfbf2FIb}!I vo<.9y=77sok}.GGOyD%xgD>bKmj||9SV1o(>f+&'sVNu2*0-d]nYv1bJPwQNl4eyF@XU3z86eVi
rI%$_8g8>P;@X\wu40El8{kpmv]xManrq\1oTq= wdAw2q^^? g$E 1q|
,Xhu
kN_1Vr3!io	qXvA"E&XynWp4{t oqUMxaJ.%?i3grMxA@Y(I5RZ/m^^n|=N@!>I4l!ix7[N*pI2}z0ab3Cu$.+T8`I%AgbP{PR!J#xySE@4|b/:"Bi/=YPS!"p8$S
yE!mZoR$]*4O_h}ZXmyq!hIY( uT"2	(uR5qD?9cWFH\}IkX/V|E-DoCJ.B$g.1Q+55(M\kcg5`F(D5BUD$O[<7@i]O*@gd@`p	gVe6BdZq*x% '(y\+B1PJy1]`i[n";N{GC94;"VO:-Y3W%bo2Hg
zNk1[r4DlACm
Qsl,bs?)~yZf+/xF]l&gI6wG! {9R.S}F)xWq<~XH.L}ao:w%P	n`Nf&,(?kGuAh-V3ud`E	3ta21wrW|VPKj4LB 6$N-4pI2HWB{.Z5R#q\gw]CIjt-Zr-!O;NFl1 [5!#){U80&.Y^pC%]Y0y]ruXS1y"DzMO`^VEX]N'*M}KP/1TFK "iFC8j@"]Cg].=/Z=|TTy\)00}qbE'VdHP.R=l<@)m#gs-^3kShroS>.)cuq{9!ps7CI,J)&x|$^fJ6fyI?;_?1cS#momcAx6%4/gi"G0||RsK{qm5k(IXt_
i(m;)=gUVmUt&anSV,z"h"!1Rw>	c!kTtO5$YW1q.T&L';*kq6<OYIx0St%JIkqrj7UfB=*:LFRK>dyxKw-Wz#LWXYQevVN6TPvM/;!v6kCH/'Ju4two,+>ccypaoD4_b:
/<	JwVakm%1)^H'/v;{$*c5\TkL<nUB!ZJrv>HlTQ$FK?*SY'wMb=B.HJnR0X\?kWG/?nlgO
d
mR/jnF.Bw}uGbO4jybg!H 4`3&sO-Wlg|(5V7\WxJ:<4<Bn<Ya$7NGV~@fT,]f9KZX	48B"G\V;=H
YSpkEUv+S55o,Fs1/7YCT#[uk?[:[LIub^9Tv-"S5cu(7vDg9_y<2?o=47jwj]ot$Fz @2>@s>!x"bj')b{vv
ek2},P=^&D,4G6ZBefQa?!{Dzz{yo-zI|;&^.$2{gkz.Mj&VyXoc8)},"T|T|GBby
=>OmL0BGw(jI2BN>QWoJFa|p~L+=3uXujTKF5@r[dFqF)/FmS5nzAy.Fw8.,]C+>AyEK634H4p;H?i'}:{CEQ~+
?XzZna#XOzW|erA[os	SDW~	g#dINO!bf37c07aOm.x
/h	?wb$mM!o<f/mML4UKLqHw5;i?Y
E?GufvT~hUN^J?)\[lbY:0r{J7rB]fU54dF:W\gs:ZKd(|!u3F=FN9MC]Wqk(&p=7p(3m&v/)3'Hs>^uJi
x.q[+[C2p[^~m-MG-l?j_|==T,bKs^ioHuutvyjcux2JWwcSwc_0i-?zpxP3X!;<Z}-'Xe!PlOUcL"HWk}0$>VDHP3X{	HOdURV*r/-%*bLsGdLGH!	y m=MypQ[5!-fo I3(9*&m5vAS%Sq3/ap9H;s3V)n^Lwvn(s<|<}NFKnAfj^xXoOuI>Ik.0u!41b+a{VD6Tw]+vsu12f5i)4sgDj[&pS7J@`*F.YLEM_)p!0[$PF2Xw$o74`dv!mmYXkMEHxCZew$N,+ZtiEy$@_Up$i*\zn[t<g{P'^-ozalPG+9N.x=gRmI~$J^ WETtK2m%1kwkfROE7rPTE[P:krJ'TO0ywMO])~+\xNL+p"Cevh*i"
BY?L%B#[f'62g5Awf;{4Fu:%C-2hz~.{rKHoh@Go+7-xv%j&lJ%+_M]ct	K;`=a:E$X-AnnSVMrgeKu>k6~#EK5gX56tlhL f#|sK!r<T3Ez)G`.wX>vwK=1tR[bCTo.dX%ek5b+?q=mSY[e5g)Vwz:KRdB~K-l^Pc dCDFe^W{$V;^fS;veUz?VaF<As Y)<r><-f`Sx'~Flg|I>_h4cvD6`(4q{(,}j"b
ux+Uj=$[0Buw>+xD7<rt{<5dGlFByX^=In RHz_g15 |bMzVH|d:'hcZ'RBO3?ZH5K`_9v1s^hI&G#oXof3L`>WJ[y29ul{KfWXAv\G_0;(gNmt@?8 N%nC|[[QVQT}[:	f5H A
ogrJ
MN1>a4|t
JV2S'II:?4aR&&7z"\9sz[pMjt8>8;kluao^7m9PX_f-&,CMpSDboXeXP+mqiU(;6%9
*1EPKptZ} -C-Ga'p@)i'w6K>:1G{B:,{*9?J/$.rx)%Hcg66.FDpMsd{2y|yQ:lAq8(b,<~Z1Hi1"+k8gftE'E+&/Ch|AmS#tax	,whhIMzNzf=:"uS[S"60U15AeJL	qE~r0Y"tygM!^5DS *A&_taW):?ko~..gU{caM9X[-1b0Qq|e ]1>oN	>7M6FuC0#W&RDH:hoQFnR++'nAJ a4HUS@<G}v>X<F$:B]=);VZDD%CP(EW]SVT:DO9tpC')\1A:ac3.Mj1xR.z~#qH;Ud*-x0(	!zu\vY	x	n(Ov! =ta_y+$an$`g^A_$GsWM;zd/l2@%/U^< j3vR&bF.24eRe}s2<cq4RKt:(4Kp:\]i'7 M`G9!6B.$`%|ufd+rr"W$,JN<J
Z
9!j|av8Rf@o}csf#GCuqzs79&MJib{&`B8[N="#vQW,CLx?b+407/0?N<+a!;(nA=MguRp'OUD&rID8E8@2]v2ZP$JVX{(:n+{7x	]'{h6u^/iw76d+,YUh3H!L.gA@?04|F8W"?IgsS1-Y?S-%a,Dxu"zG6YX:qbuaTNE9^C	f6$k9x2iw*k(O%?sgG6LHsGCgK>G |}C=7'(8H[S&(<HHh&IS'GDVtFO~gBH9\Q$mp[l{X6_$k.{l7m.@(BV&KJgU9za1\#wk6<8.AT%cj]XAS`'9vK3(Fx#s J_G(E+5n-wI&|fj5/5U88Tf9P=3qIol~zO0v&EQV&hiztp
70xHf(.66\l7lL@= \:3*!|-VOgK9 52_U_+<cL=%X	*|s>wWw6Z6|h_*5Jk+YV+='diV|Y/7@k\1(jhe20Vun9)MSRK|+H#fA|-r>#PuOU~\d"xIS	o(}=uk`w9"zAdhcJGO5dHU/pk tp*TF`q5L

lyZ7J=W75;7G4ohb8jfjsf7eTr[-N7mS5{Ar7Y
X'hKd;y4.yyI<hbLm,RZ^4S}7j9RJZMHo|[(SbVC.Loq16@!:4Y^Bve	YthV(1B,O<_[	GQ6%02X9Twpc?$R'k:w*U*n27?36tPz%vC6MD%v~1q4!eM7}ju-~}{<f:mR@!w3;G"a2epfdk:n	~}E4xP9+V1]DO&(&$$MdTot&u+;\2$c)q]gs4EXro/0K!4?#bH)ZGJ*6)5}VEZ.\BUuZ*QT'0N:|<M)-8!v9_X7}sz5p}*Z,NDfi(>
En_:?gN/=~a~gd\!am?J"5?c\26mh2BIk\Pe-4k&VV-;\W0	u(LcG7aNHJx5:hZT7Q^u_ A|.vB.*%ntga3Wg8 r=Pn!.hu#aLUqMk_[`l^K
Zqw/1F[YZr^eD>`D(i'(w{0]j6VXIBr~2&&4L#.aKZ,@qb[=ntl{?+B)RYcz>lp&55`i
@+?N1EIx{yplfG28{Td./)Z,vdT<9\9\
( '/Y`aX_'by(jxsnXS[dy3Em& k"XdCvF*5,Y"Jje#)?ED]z'9G]D+-an1B07iX?/_5e}>Vn):"wOPP>]K*El|jT1Q2'0CoG1)4u%^4O;JqZheWxX,ZO%(W63b/2xK`::Ccj[+l[g`a@p{-eA[QgYkRfwthXrKA(8bmeBGsh%k#(UMf@m)}NV!Ks ,}?m^~F%K%4r\ANNnvUF`vs</	Tz-p?VarLol8Q5]nTBq tL0G4(2!KA(i:p8_xq\Z`{yKgR{'Kml!OJ.k:s~hEv}EGxl?E~!Qzv:/M-?r&w	}/?GX]uU3njtyYic?A:Y
LmJ%|\Pfp:vK] T[xtqG:[;'Eb/%|VyO.u@P=`tBYCsy-s1GJ=c.MV.k9Sy'T>DAOAf!V(<XoH0PK!u!zx!Qk=5!3`k/
&\ZL:>AuD#xk$"5{(," K5p}O^+@JNPJ2Cb:dAI>g,SOF5-Y}*UYb5pF<9t%O05Q^_=__q=z0-?fv,Acu<Qr#Tv|3<C}l=_b_H 1k`M+avHUj_9<eU?^m4PpNpqFr#|YKSP)~5rn6_W'S80B*64w* zD1U
y=JZXgwKVgj57a+F9Bw+nfjt$|cN$eJ~-hC[+*A/l$G34>b"3Vnhywj;}./L`IX[5"=gR3bhrj'};FaSRCpMdCRt|)o5YUK4L[zBw3T)3!`<4PV5vfg;@2!@SP)cf&t+~;DM)mJ	QA rB3f+0Ng19]Ai_;
eNIIe]3]@-L.%!KvH/`&t0v2ZP+Rp_xtpj`DKrIh{{6t}kVPzLvG/m9"A;Ng?e$4Zwv@X=V9Lp-IKGJl
3^WdE\KT":
0t+&-o~'ZL2jwtKp~`iyep%DDhIr2=^1
?bX8;knOJ~xB|fW_VsdQQX'H]Kl3
=.|D@~g-j^&^T5	DyA./73pdCk`B?:SUrJ5d]o7a5_Zal56W_`,
S)U{X:'2B6vf?dzk::?mBx&F,%F
N0S,do*q<X(4=<l ]boq+u~b#a<w!R%cbQ'effOAHM@<c=KYL\BdcX,X$^t8-MI7cgs4`UhgtbA7Cl=!=H,%6CB8U{CvJUrU9>JKKm^K05]Y3R#v!saONsO&<%2s*C'["NkQh49IG_/Pv$H8(p'SJ5$o4L6	\SEStH'LU! 	GfA]j7'5Ow)34$
aQ^sjx/_aEG>SET(8yfC
Z>wV)$Pmk.3`E
pUMv{WO4wYlqc(FR~[@si5$/e>Lhgqh{k^<^j+U+f^XJz>g5CO(P>^`GRy%gJk&S*-Z/dxx?hi|$S+:pq&MbHW#,}n@Ve-;$gnb{hM>qvL	|+Z2
0X2O;_;QyqeI^>wUW$Cl+I>i:6Hti.$#,q,h}t^4XBR	QvE)F: tRYhs9ScqEh]R[th)AUbQXqzOy`Ju
LfQd\}T6,Qm3?'Z;,YvOq*>QDy,HrLg&vz8>Ve|H(6-#YY4.a33x~F0^uOVv{T;YeAc4"uJ*5wssZg=oXg!S\ZnR@NB$2^pm_J:R@TL"=$>=:HXW'E9/9:"t5	23?cV=<A	Vf6GfN,s<%K%0Q$n,Np~")	^fb;CMH5P]x/Ezi=>}sx-oyfi898Ek%d:\"F-smGD'}@WLc}N9mzi}9;='&jb>2"BubKgZ"5:g4:+=H:x
W'!Y1?B_L$!Fl<6eK/J~8.v'|'y)Z$|Gl6MBj$D48FZJ5qy]"/t3m|=0_; U-g0?10u+(A/`Sh||8<R@6Fr{tLp)Xy^JNyk`#`:zYmg(yW$/"=+5A
~O'/M|h*=9sWbf&IS5x2a-%&zP=n@sooD_iyZ:@CxF#BiC:3c_Wp?#gJP	PascJ#3!
4;^O089"V)z/M	;isN)& :){>OcLUi<HI$c0Du,rPC^g:@33	'rG+Fl![&(E"VnfbjAA0 <(PM!i4$fj7u`	(~\xiEFK_P0-M4%3"03wX6t:g\`jmdJ6#rms)y~xIX_216w7[e~4gyYZ%:P	h;	:A|mj{Jb(%'Gd;>9uF3v{[(b!<SH&r9'[DV%ANgc="i<H>N;TBY{Qu}RK+$ru=Ee4	EkG$sp>n&VK5;f2SUCa4C*=#aV1%H|RFcvc;4fJLg Z|6WHCX;
F#h"=k@E6UPS~5q4"$,!\n]&^{wtGuPz~/c_J01
# |uX>v2}S**Wd,T2uJrdP3>fs1/-X0@2`,-ax-YR>mS@H08=
iHU}@WMqeA&ruo(#1rM)<!y`hV/;$6IYI(eXvT!>^PUC^S"oi]( CQDV)<L92&+=w](#9$xk	9**o6<"8)izq_Gckf(2=sPYp=TQy[<rY&Fxr>AEsJ@+g"{1&\<L-+4/<FQN[lG*-)XF=*Z<HOjm[@]{Na!\ff!>Qp')JU`<`mkko.}sgVU@tYeoPieWbolI({|.|s
-S~()aDU\)\*/jN7v[d?Lda.YoGTwVQtVno{b[4=9YFCj8o%=;]*xvM"9#\^t4)DY,X',P`& _QI,@7mEXd:-s:I[o 57aDA+hDq7h6ivp(F\am~@z*U1"2}7|cYBumVGfEA-9tB!HtO;'B,SFTsg,h=8Pqc9z4kv;afB|3_\,&D3Yr Q<wg
]n2mKAU|;Ov4!u /JEIE`s0%V0ritYD]!kC_^b8+J|/Eu?/T	)(rUc4#YkSmpE[CC}Q5)[
4{2MN?{CX(:jy{$;@1vh2EAhxNq=dS2AgzUGr~SBJpKF{rAeS5Or@sOo>37i%QL]I(ZU;X;Ei/nB6P(uokOela(mSYK#I>F5Gko8EmWhFpwyo2M?vwzQ<#3w"F^.4&B[Eq`N@6d-7JbL'lZvl:WE$<1}5g^"6nNb`{WcGhD!f3[7@ON,O}Y6i)DB5-Cw>%}O3Qxh9[rKu|6)tZ4irT\z:b"IYZgn%BCn;h)"uht*ytTAgQ8#@:^waFib3[eTnHg6d%3\G>@bVtmtvSb\o>D|^
PZ7mFnkPq)2|W8,?j_1;W\F)%Oi 7G>Pah3}Bwq#Z~mg}%a-h	&d)X*5YY/P+a=+6Lci^!_$`rUI$ay5=&[/va'iY@oxs(2/vRji,Xs=RI7YWWPQ*(WvT}K
V6Bj500:N<ESM9
8G":Uau
Q-BJ[=~,/2#io&D[%ZpvEq)%Z<`?HD_>vKAQqb 4m`Qf_;b;@
m4,z. cjTv387Dhat6|HoQQ"W2/lR/\X_O.xZoIZ	^,r;uCU>_
eqiV[O*Wt$t{p'A^%H8^Ru{kwcH}fd^FG %_WOQ8%I)"/G,W?e)^i_!2nXJ<'$FXBa]
m%tX=1hJC/T/rq&!jQZ*Lt-|)hF"=6ck&N<j.[n[it4 r?|:HBEBfO"M{_T$T4f`=hJxW*?$"iy/jvix}tgSBhk<}5E9?/Vubc:5*:2 9ap>0ua,v{*^vKMV.UY-r)sp#gG&<XwEnR5LI#"unF1M!Z;l2Da<(.7LIH?S8"y>c}9aqH~Fo7c Q%zkqZ<Iqyh,vr0]}KbK07Q`K2Qgp1Iy4E\Jw5Q`p9S0V)x6!Wm6\?89/Pogj	)ci)Ly:LemOJve7Lo'=[YG&J#w Tzl2\XybB!*G8)v)oW;z7_rc!01iUM)p|*>}b*u0}h<imH:'{t`M-(r7J]H#U#5[Y6QUb1`~d8)2OdorV4}T-Vz0&dPn}V-
rZ//PdeBp~^1;ypk+e|rUv+
Oa?/.
YTI,=GA\}17S\im3Xr=	%<6@6&)6O<);G;=2[j#M))?VoR843t#krY$h*o/~ueiM''y+UwkSp5&SGY'\q6S${M51B'9
H0>H*FBk//b&hZ}UZ1@#%t#E`C%?+4 lYg5y`[X_5/02cJ
US@H7gq$7lH8y	dE{*8g`d3iR@v$"e%T
@~EQ
9&sPW2%%;gNv]mRY?M;>dI$^XKZevd/1:nzx3Rq1%n91i.1`fIU%{;
"=we^A6/\oW$>JgxlZ[h^PyR1(vu4[vaIT50?RI" 4,Z"xq
4-OaT}Vr%.Q{br%3S
jL/#huM9%&~dE{<|,%dK}C`/IXW<MjL|t%aRHqFDyQ{%F97Ln8=Vs:3:{5:{]B>C@\EM&IAay/g)$;P]C47Q+I7KB1BD=M~!:b+w
_k/:@n\@2^ 2zb26yVvFW8zK}G<Y7pZcn#;ym2c|lM\UrqQ=_q}8|zICwQH$ai# 7H_C /a	bPIc"$UwvjD:j1;0>x}k2+RypCn$d>mI:]gqhn^kY*Z0Dd<<6L"ai/j9?N++s#6
!\Sbbin/hlg"r0u0MK+}v*VL~JhamS?5OlA.[wc=_dv)jzrvK]Naqg^-W@a99;..2AV)Njo< :z0e'g+Ea=2#,$H:QNHhJfVw]3xnY"YPz9.w@o{FxsMVh[N|.O^l{aFn/:[^tx|.J.lv,P0>Ngo|Z3'^7 D
&g\#,T$Ug~0{mZSG8W0T.4\gf3qD/o(EP3zs{~33Lj5*h% UA"wV)5^fkwT,)BSz-q!3
s\I&/]"SvcJ1X.&YA{nIulG)nn%{zS`M9Z?VyY(Qk.v8q26n1V5Ua5L=4N}Ih(&T`C1;@)dY0^?9=~C*E{|/$>qU3fLFzy|mw.WJ/.c>jk\l1a"xqzER*>-~u98`eqh<!jme>;am-tgQLKR
\@-9=q;mm&|	eHK2mpd:|QAQ&XLt~AV#/d (gR4lBvwK'&JS*~Ry2b{:wozqfqR{%IM:}eJ*TtVP&+6`oe
>CYd<fn<@tWQ)cxB'}9-"V\G;*?Bc|'Rv`I}GT~J'}q+A>v4*`fIcU|C}%Sn(w9Q>&F_.2Va1e2FVk>IE'%C-_5@O{hrY!0Ku?vI.[I%kPkU@5SpSPo^-FEn5|:/cND2h|l"-O6utI^8GcUdwjjG.5Bs9h?1g9^X:rRc{NC |bGRn77n_MT	<qvQ.(u-Lsh![?3c:SIxD}pQcjq%0r*&(Ippwl`*f[K%FP{!.|/r;^YHp:'hXO[W@wgca/3=KN1xt1	2}<(4c#sRT8jF$=Rz!qss>uS0za<c{0>4L9)*	v7hxaUue,ei"6F	;'T1 35\WDCPsn;$aq1	i:2|8CJ"+|9cp=tE ]?Hml,9lOF%qQ]P8:t-dFA_anO-BJ~6A2oIA|7ybhq3?`o3(5/	nlOceA|Z[cHsXXJ9b(nWnG.`=X[:.%/2i86rAPy/[MSBi?A*]or1g .qwatSgrQb,p2YG%|?=se4_&FcpZ?d=[YW`.'T]
KX'872;6A-JbKBGZMc+Ao]Y+wpyz0rWUO^#;F\+c'iXz(acf!0z{zsN5f7HvUK_zHV9#anWcV&j];+,9@NJG37lH2Gid]xv1ud<WSpY$<4h5tu6HpgS=G`0zAL#iJ#[MH $H_kW%WQ<U!z;%"o]JRTb|M%9j\s"}+D@)D]:hO8$|xo})#LR^>4g.|:'^UzEl{PzQ"$lotlk,`,fi$LG.nQ|
.'> U&WxN	m6%9uy:[X(kU?8P(mn&b:Y0vm_}6#]:flD=ctI7|6!g^:0';
t2JM?D(Tf_'OS6o(/Ok$?8Ro#Qj=Hhih}oT<3[]G\0+:#o!37A
[8C0
$H1hS[/",SgO@zQVP!30i&-GI2j=L#[([7|*&@Z]0T' LWc]L<?iZ?.KE1|!8i$kJStKsS(*KKF('O2jvALai;K
$Ju\BDa0AvE,<3CPNe<^-'*?
a%hv!fI=[@6$%}yI}7!K8Z%y5T-`Rb[yasB@)*5{d'SThrjN` `)^
Dj>	NJ!L({^3 #lF#.yZ]`gVhi8'!U0.$x3ACpxr:7Q;#*gR]siJDxKre!Yq}^D*wjOC$4e+z-X>iuk8pO
}YYb2V
,5F6mJ(%@1"^Dw8yf(~Dq%Csj L[T9nf\f*}W.W:4LrIcFf<ksZ5Dj,APUYL7WphL/kOdG4D5O6EY<JoQ0fm6/4R*c)xMr;OI^(TSWot%qAG|-Yt7N[{&
e.+w6)NLQ6!iG"kTwX+|4BYYhL7Y.&~Z.^#[vs,q}hGYJ#i=3#22kaU0iS"_`OOI%!!4\R_cWyUtQbI+eu#WGhD5-J^J8d6rL3}%6Hn3drRdCTZBz#Nt*.!J9vT8f?+GSy!r+bj]h8ebvJjNvv>)H3RBP> dbxXIN_QE!q;=
,vj[?cS#^Mm~n~<[1f>D3h}GmV"/l6FMC)5aRxI=.#_a_O]T%V6TIR:5j#A*r9}m%/gA*YgZePHjgiI[Rr2v4Uh=Wo>Xwu;ecr}95v'LZzA@_0~|/$.h+=`W;JrINKANK<kOf4]}<4"\q6~WiC*3a'Fxtd38$KO(t.r4&btf#I7,9EDq|p-ero$3*&[2aExx[N{\["f'
7@;scP4%Of:,'	$uT]gH3W|,|m A;#]8&%metAjnS% V9j[QP5!Ek
/oZ>
U:C7g4>x](cM*YpoG`0M,5sRPzX&!p(+$d)j~nPFyY$8x$MS3s(J1UDh@+6pSFOG'dC..p&iChbQC09*CqYGT'jq@ZZt?0DA.n`-YV-|sb7Hd]d)[/-*{QL5V]df=mkG)`!zS54Jj`lLa'Yz&C!p5/-^>N3?UKeiILXW|7S.G5r\,)#Os1t{*
)SnR{}&PC?0U)BQ
:3O0yG%T#L
.t7hi::V`;kzNqG)WKLf.q"FA/M-	pG@I3ja7s('Vb]v@xp-l+*sj'~)@Atm`Bun!tPr*$c}K@"BT<5F2X.@Mj%G=AzUs&.2M@`y?v D)5%zYyg]>{-m}^kO'K~d&~zX8uBkb.!	P^\lZ88Tm
AD@6NoI#@kLt@T6J9I<qO~Qn6jfbSsm^[8'XI78RoGr,V]%O_?S`*nsZ=K/vPV[
g1:4,-9\%/tMOAk=Xj0P%Ot9$)IoV/FR:6;^q(D8.+M6jFwT1Ts4BjAr:0B)LdB*Z/]J.@B}hAHYP{&m'V_R{+p*6Rfy	xJ}^j_$Ie|lR@Y$8=z|F%:{MKrQ@/,NLT(A+tZ!(}a=v],_!2M:d8	yLiKILacc7{U*cY0*H*Il<-5.>_ YX^Erua<Bl=V0x[3v9T=84;Q8WNY!"ArV	Ps*#T~S#<z%	+>0u3D5^</B90sA1POVA+Y`fN|4[7[OC>)Did)z%v	I M?LlAGxq$&)H	O(K1lAPnZki.e'Y'<fP|/'zSrI%8*4Wh")n{FI,@b|fqQ:8vcO5cxKu{9`_;f`HUc+ftY0*eJJ%SM!coL9tGm1!Oc>%T'G)zO;aejSjuo?!U6-Pbq @jQ|=^8!pT'fHi<v&sxo5A9{&j%Yv#i('UJ311~+?;IVuql`u=]}wL,(AWj|3`@N{]Wy|6`^;#3DAJI"B`v"RUSZ`&|=DLD|[(4+v8Z~zs(Gg
b\p$N6$c#7x9Z7}FSj@C51d0nWoNdb7@=Fl
>9HVUiq=$-3{
aF1&4A
N3V7D&H."yd-;6_A<t	
jd=*T>UD/q&5?e$KQ %( `eZ8eh%R_-S{cYjQK JAF	*8
GJBc65l-+<%y^Xl<n/T!GCSg)Zs
HcJ/i/@UF'#FA&J-=xCm	$(p)\ouL?OcLB/ZX3:{D@u+q@On=}FCy
S4(*|"T7=`ji*:(QWGW64=OaU%;GCb{G12\dD&|a%5N\Jw8Cpn<%>NFp)%D,7JPKk	Ui\petL7(3BNEz
cefzRfS4M(VcvaB7|%mM*+|zi?	bdpL6h8:#RmM&G6o{1RlLC~#p\:"Ch"w+\w}R<#w\nK}xdT-;m%U#p^TIWZIdt'kmK3lbMwifbK=gTr=.OT@)m0Z;9THv/]r]SHO_B}G9f7r7/uFSYCsWMq>K^#&!4g&5l=4/-urjDM>*x!QSUpZE.5wISrj.`LP9n1G_+nO%*<77v0}Q.F8X4mE(]1=q3iTJi}[~),L{5MI&;H4nf\GI$>{pG`^ ;R'xlX	[Fv/g`jvz-?g0va3k6=3O;P@Nk?fB)|qg!}	eP*rlBa^SMi`KK?lf#p<RtwW15qqW1hxv1y_:L8D$<&?hb*GgI/,f<}lsg,(LpBxsjgnkRESx	~U^zgtmSm/xNzzdbO"'^$mGj;0[`[o6_}['DAZRmPT1:?5NBW`LC)$X7FFQ@%Wex,]%&3dU8Lt9BN0Ph'LrF/ox?8		0`y9TK% {pz}B\frZ0KKOBN&,!FvcPdLV/*AR
nY37xQq\tY<:)2&\REyy9wFjKIO,*rOwVr3e<E*6W#WVd`qNZfc]ekni8BzJ7
RV5&MP.DFFI0E25^I$thb4{`\#_e>CT>f*UH`;VjX2w`0!5xp{wQDHA5W.aS:cuKn{x@	?2X4uSL$7-#_G.vm/5iGrwtAD4%*'D36`^IjBaj} GeGhsM}AaU5#jje	kV.Psf]34{7dCc-=xb

@al"a==Z0QG6_[r&X,ZZgz}	"k%,h!fbmVc[zcYxRc$>+{~IcDqXU!Dy.?v=RpCx;,<yH.z/	0kGWngDSrkg?o~nc15l+G3.6EiKVc+uvW<FB?>/'_in)x;<\P^:cm=C]ie@[AVB[g'+m>bv!_S*)Kba]ckbOZ8n\!}/46+v1tG5#x*7^<2	:X_?'RRy=
`;I3,M$1s?e;>-Y|S0=Q\=c[99zotTt[;H~yxA)Rb$$E&%S!)<>a')	}h0rm!D,y7nEC[=GV|fW8RG?#:SX#l4,0I,Ww1M%S.U{nz8O4"Gs%[%C-'2*"0y7/7&}=Nq
>:ls	lY8/+m|r/ie${M$cZA:5t%`@V?E;DL&=G$l]e*:":30O#Ou5_d
LcA#j;n]fBx^d\:~XD[vo7Yw_si0"JvgznRBH2'2L*3-RhWs(3}~/kS^v;g+J!U(DSLn//)6%|~H+Bfd8K"oE**K'h;6A=%u#zL%'wL
0+zw
x~*&M]mwC/,v;H;f@Wrq3j`$(l+&+UFAtt;P;UsC/^+VCiQ`n*c1UI()JAQMz0bv8yT
[9]LjZ+oEz,$jo1R5_\;Kc0hcrhv^,JmMpK?~4,JCs^ks/%WXRV{r.CdDP&\j,^nt3Bf0sHums_-;wQ1'hF@'=&|zg_n
3z:0!ip[g6ft\\2!%n&#K;9A&S8/2.eBvm3:?Y1gq3pMN6u$@H=xVq|JZ56VX{k]5ko/9A!QOfOqu>8OF~h>M2m"w\J>3. 9~jV@KY+z9w'PJ}fG>nc|ZEqtWJgk_D7DxG>k?Ro7
y~th$x+F%jd	[*t-,aw-5
CT7TP&cGf.@.ZenD'^4-k6
66LK#Em%8!Qe'U3t~=/ZIBSFy(e@g<>uAXI-4CI!3o1{x'u,&|%HvkiX3T\kN>(!Vh[=bg)1(BR]m&+S]j94u=FGiVa[W)[_-:q*BVD=^(FUhH2F\0# r'9Id0'a	t8/1B+e!mn8/K%0.l
*uurFGBS0[5vYX##{C~l8)wJN&;\&!%6Qu4IE;
|]3R'z_QWmG?g-Ac>._KAbV0Re[l>_))~xj(@9$-dr!rcla8uNP-vQl**( _'VV	d`s:kA5I|N]4/<`pBr cG!hp/:(~}##bDk
sHt#:yn[kGr	@O+uzM	Vecj*G;%5~8&e+OsR
N?s&8Nf5N0vIb<CVD@lO+1{ r6|1vzYy3:va%Kj3q$z'oQ{nBu@]`0nWDao5zaRYC^DUp3RZ,-a"u*nWUn^
;BJN@Z}}!|Nn&1%'o)9	;jd-=2#$.:.\^?jf&STs$UQ>ls1d)jBe-h<Cwa(ytqHNW)/	/xl1'LhSD<,.}@<0w@d<ij_#xRh;E\8-32S^qv;	fAk*.'`X(6i7}I_Uq;jS2.@v&woPo}ATtan\yRdI9,k'b)cvLxpP_gv|q.+c >M`a\1EPgV&c;x|"qZDjlSoc(5&h;$6 Bbd.n8^
DDc[eA%712k+$PWm;6&TY<J}6LYNy`^h@TwAx_ZXc0ER$=IK4gS883='~J]	9_|1%JB5QA@7vndS,k<-dh:K{cN&(c^w7KvKCF"Qyb,gY_)[ 4Ys_ombax8`Qk+32Lwy
~/{LJQOc_=N\l[6!q{NmA%iLJ(6fUvBy,C!U}'4j$KEDQ2/Olp`ZIlUYD.$rl)ev579Bz
{}16'r;x#UC^I'y\VQK	r[Z3@S4K#q`<Q>!|Iu(0izf{59GE%LiIhbc
D`J'Gujn8B07-%@98\;@/aY%(\z8^wENNOm1w#HMX%b_<i{7EhzZOuS.JJ4?ONheaFCZzyTMM5\{:6-nzvHS4pLtJ:aE[[XmO:Az?d|q@GxaAd\Tp:z>i])cTI(Lbt>4>P`h,fX[ DjkPX@qjNs2@2k#(y[b%kylHbT@C9T=r'3	~D:BwBCc}	?7}k2*5Ou"W*zF*Zm18c|x_~(_;Nr3^]gz~uGg
Xln$
pv,"RYTw!1&^BI*Jp#d6EpUh)z&A/0O,5DOHggKz`n,$r
('3 2,mL47SNaLj<k,%:{f]k>iA]q_l9[{C<L&iEv0F9<f*%}h$;5D`\1]`
w2/DJ{nKN^&smzh<>y
t8w2@En'3_mBV=WGPh;!llpUHMj-)IO)qR`Y8HD~o~)! >*v,&zFYW`jk2
5C2;MC")^&FXLc67Y6J_TGYWCC=#RrO1U/<g|XYq1^Z
c~kKj#jH~k#lUABe9eg76CK=l*pc.CVbRidGJ#),lJcJr^[Swq4aa'
Y#*^eEynagRwM68J>"W~<3
Ni-O4ZoNbr^-'
XI.r$U[S"NH-|?Wm79FQ
evr7S|C1`Rk
P]sv>c[kY!}u8oYa	
@)r:L-oD$7iLzU/9?2=[IIU9*#\s1m6
Y*N#hO-*%*Eiou`<90L:j>ZcQI:yI[2zhAy80amlk8yUQVfw0=2w{zyUEG=,tzLfg_>l;WN7H{3b]z+[jE `0DK4McN>N*/&=
8]{&b3]Zn!(SH1nIVYuezPP{CTwx/tk~]L(`.AbpX$- gcScEVP)xUs{GlZ<fo\QS^@;h;G#;K	wD$7Di@xa`FFwIu=%`5SJ"cQ[9R.Te7XLq#!U>Ix.`1,2x"=??>/3sb_@}t?"sbR.):X.br^u)79f(zD[VhxS&IFB`Mvu&NS$Wa[UPBayo153be;+bnl5^9moAb`&'Yz~sPqOG5B{l}WT;d]>w@vq$Et_Q2I:O|Xs]{(imYCniiXJNS!" `ZbG'BV^"2YJi &KfqcY|7yJy|x"Asy9jbkOpfapX^a_HfI/2fRp*i(mv>[%cTJp=qr*ygvDrm=@hL fAe- $^y/@VET1#B_gRt'3}2/KQD^5kwW4J[olVV*LUSK|!>Cf[#60E1fG|2~nuU_[Py10{*/o!gi)zGGs}UyN
E^&Bg@masIT\SYONM[R.HSqNeds+%pSn*;0l^(fI4
xP qT]GZ}*cnri=HQJ8evvxG@+uft%u}/)7cgUw_Fa8wv~q#&UtaEF[eV-39IJq%oYlWQe,Yd)z.)8Fn>/VvrCwd@]:SC`f f+(61aP+Sd/*056"3Q:o]mSe+DnZK hww8g&ELo8|e7gq
w
rZCM_l3}{lW9NVe|pQw[SIcr5Z @/GC#\gY	+?_J @fCxdsS6imR,=AqmoY1{{DiUwrU:?T'[yG	2e	6#tDJzGPK:
b{?1T
:g@Ugv2t54:(/|'ySVsea"yU~r&=3go&hVwsYsB;KVvh umU@g:z!eN.*nKX}AC@wb/7z&l:+  Bu Uf.ATXGpnUm	@+$+jnQ>CmD5Xrl"A(p9NrRJQAOr4\ee`0?8X:-,Z"&X+e4(A&LITXG_hBxUT--E@30PWA9F<3CoH<-01NfC4i	dKdj-:Lw]yDq7>hxrl2lH3Y?'z=a.0TfyF54?AvYly{*TV`OGs,'Lr0F`kdG5&)gAhFOL%Q<lKr-UqO<WppS3<HO!3{h[M2t$0O+^bsx`IJcYU=FL:\%dsBU6o)ES]BCFFh>S4s7tU!kr1T@]eIl`qFWA~ x{Rpu0e
X.;Fx(8+s!r]:Pn6Sc{WXZIJ~VX2,