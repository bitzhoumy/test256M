gMjJb'=bXmYON*9>A=30z?gZn\i7?5*NZ"ob7Fdl=D	v,K|S%$:}L)6MM;2v2G,wIn"w_!l^!AvSrnmt6l)iKf[Fo.m.Z-v]qQ"sOZ0Ns\/*sEg<Anr*f7x(!A7bS6`cDiCdm+3iqJx5}a/mU",{2~M-fs_\03y^%CW;Awnsd,eU@,M$w,mNI(<HQ"1}f&	*2i[=1ys%1X>AaF!z W!!duZc==5cST|/D;#W4hdIXR:UCmD_-*mMtTD6g{r]);BCa;cq6#4i<xEnwe7DBoI>fE3"J!!s"rJ4#?>%	jEo0-(1@5oQG*@X{ooF-Q?lk}l!	mZxe_[\"U%TM*_!}ZAwTcmL|s-1i{QsTyeueM})h?`W_Vh4=7|`F{O$`G(4T bqS1s0hs1)Ns9[664&.Bj|5yo,YjNUNH6\9mXcjF_QD*#g}FbPz:uyL??IxDNXgv&eUVKkf^82Io/\/}^3~B38p+&mZJ)+As#o"~
o4&4@U-LxGR1E6@7q@K.'+/7#:;?2Dy<,M 3~Zwp,*MXQ.r5l kV(Rh3yZ7B-oO.AH6(5"D8Z&_s#&jKsYd78``X<?|<=BPD|Q~_PJkL`$f3?.]JerR7n
',nNr*s=%)~9/l6W%5MEn4hD:Hu9Q	_6Mi`'R55f`!`|x}2d<4_oHBa'4-HvAd2bk.Yz]lIY:}uZ=`7_;h!<ZVUkS(V=0I)z<fp2P[cs ;5~cZ_PIqc3:62u	qB)c8|/a+d&zk]\5h?#Pux0`^n)2dERSQ/[GBc9\NZ;WI%2bG[t*r\{)li%Ks8y\	i`CxW7{28e_UMIohF#anmLs	\>yuu*``qy#so8uU%7EFh$P\;`Uj~#Y@!bs3&V	pR@2a[KId294(j!SSS_DKq1q):?:gi!oRdJq	LJ&SU3}Bqygthu7k`L)l?"KO(?H+s G2b8p@B~h&?(uLV,i3K(}(B*1 @"m>5!)+'i/8D:Nw^'\;>>T]OmgC^|=@=K*Ys<Z8C
R@uS|7gF7w]9eR=}4h07I~	s#T"We^*	Eqg#2@pZ/wy)-kndwXSd[Bi}f	:p3k0w&JY(u\dKRy{|Ucd*S_$3#gT07D~!	lvA3E."e_@<'OvJ).re5eZ/sZr&U^qVqR!DL>HdSrGml%I6"i,<=P)^JJUzX/~JH0?s13J3PGl^1s6gA7k5FxQ##0!Aw(|g>FaaUo,W%U8`5_G@}c<nWub;\n(i'n]
jrxaD;\';wov90gif'S[QA\,3,v{axsKUM^1>s!0OPz5Un-ks&Wp0j91BJy8"tIr,`6xn37.q&tw9[o'o_^hAVP,xJI2ptVI-&~;NT9XDpEp#1Dri|vrh	8YiM/fgXsc,kxBO7`?|<#PlDrBj7ero0dxJ*xZIhmCsVYl01306|4hBSNr}VsrFFi-Ofqd<y)H,?S!.riB<Siq_LOrSt>mL;/_^ax6?{ ,45dspQ>slk|`u/2L8y>|:85Sv'+%ECNd'EhEAFb^g!S5fMN.QY0')+hI6EhE1xe}>DCSCl] htK$((ga0(Twe*_qNfcSD)$lKK=._`]eaXf6|"-m/eg4BtnDBoLhWyv,I}C2zKoi%ab1~cKSWE41(CpMm/)_2VuVT;1},f"svLx^9xG5@(KVC~h#er4ljb"oBR_ttVN!{XUf[
(-3"cWGy(Nf52y)>lCt\+9=_k:2eO!')dnF,$L/pAHE)2	vIM>9=+68	;,Jh}KA^nfCt}U07]6_CaW*SOI?IsMqRjR/d-uf(A"*3;ho_Xmz9:z+D*BL1ckB'G[e*BWXdX}eltj$M^7c@/Y;{cc-g-wJr9	y/[QVp{s[pPh[j	9`<dn#!:X
oZ8 58PXdQS>?.?v;HtjOqamiXfnxYu?.I*d}D?s 6qr=l@0XBcO_p%_NDn7nWPdYN,Hy}^aQ? *TOr[EFV-0?JD2-Zetr&M1kF+AkwJ'Cc.60U.-RV_>]B:T3ls3'= ~F$T+GRu6 ]`aoF
YDj_bL~uz?E@suG(Qmw7!1?%-,8b2dgpbQ1$=.(^IeGxG<r;E1>^CQJLjrl9$luPsNT2+%pVrcVuzuy|jZ|PRYC74Md:Y2`oTAvl[irF[e\cT8@ivYh h?`)NKs:J"#2y6}aW4!lwY<KW27vv2MqHoT;u
#GGhQ9@QO
&T4GOB/"e|MnuoY4g{M"Vth.+o-\VhJ/xngXZ"lgDF1#C|NA'#0CK[:7UQ6LNBc{ .x0t2|rRXX#6TJ.oWf9*K\KEHL$RRYyt^l+C&y:}k:<QfqZ9$]Qh'W=Z{PjX}p5V<{"DCD~;{{k.WT;o@}L[!WA41'[o?V,.pQZ:5=fYeH]`A "m_heBU$Sht^{<#~T`[EK2=8]=glm?_e()SI7*l(-2%z%wT/8
h6iozr3V>awR{6by0~-/['O4=jwb}#*S7XI
.;^	nh+-?/.)
Z(t7t,d)d:CeB~VJF[1z;}(n~zY5=p=6siVL`/65d.lL k,y5/Zl} w=xi$:v QD.!'{nVZCd0zP#uF9K?t8l"j+*SGK/9jpOR*aA':PO=!%]jXqsiRt{MSp+HTL+b8+PCEO27S_N\I"+)olNV_=//+IkxRKyw9Vb]z~S0/{s!8'&t~tXlROrL({=Z5EB%ON'QM@5a&SVM
kV;o	vhgX_o{	&y>7gM_C_zkScPP<Zl8t7V0w56Wof}5$s-G.Q*\T[HG$W<ig[#_g:NT7KG')K)~Q@./.0HP<84xY71oYLM3x^:HW'1	.,>z%YJ.jg~$ty3L{!tX%A`p3'>-8l*s/*aH;w+9_tVpDk3P/TbT40fmls#		w)"\#5Ep!KXx89DB{OEf91k48wW"W3CN;]iV%kB 1wZ?ngt`tc@G00OhITd~Hri^S60  kii*axb.=yzJY|Wv%:cdPY/WN&3gan@QR+Ou/&|\	@SC4,V$eVDuz!rv,_1F{(Im4cnam:^l*>1'_7E/we2Z,
U{&W{zS/xqT_[b)J#$^ r?]sZkm664i?LwySy$L0q'X!Z/\*Bu3V 9N@|V+HF` p29~k*lk#-t49?IU%gY=6;pV)<}q
iOW:!04-mW<]j&c%mhGdF9pLyzJL:\Cx/cgNh1^Ypf
7sbfLs3/Dl"d7@J"W|[iaq0kY[VN	\U}DpR27U 8,c:nOtC<Ww3ME"g_;YG^*cS4'Ux+v?D[O4*_-*n:#\!pe3HDatJIW-XBXhRR=Xof4!G&#T>G"u*?W}9]/pS_OyYm6Z8_7O2K37S)n
-DD=v]4a.%4Gc[(VS+
7*+$m}.]9Z??DT4Hmq|=sBo+~>5L`2Dk[RIrMTq?L6ONiuL7NLI5\<$yikmFF3>@9b1e4IvY`(6Hf"~SAa	l!5~i:{e$a`O@PKje2iD==])q\iOS&0!4lS6f,o~PKVG-bvPI[8\%Y{PMu-f`rx{5BF@I#9X"6@".-(\Z7PgitZ?lVIKhZ8#}~c4+!Jkxa4$D#i$byNz6Nn^G$%sfJij8X5KtViGRCmqU.4+%EZ2Fl{7[!]9.*W4WBb'b7h	_wS}Cq'"JMABOlS+.H)N,y-n6ZKR3!=iI2P@b9%V$uS)_l{U?lw 6	neM6){p{c2Nd<-?$|c&1"e +NztmyeEP^n7~`U6k)TBh>@PrNHY)"8N21)JW4\OPO%,vD+6x/3Z)xQc{OsP7Y9q**K-61tux]JpJ/qgvqxtzHC6VmD7qSzObwi6Is'_1-En4V6O	Cr9UpL?[?Gyn#h}T|J?U^1OQK6RdL_OnZ|Beoc#X08<d),[}8/(:(Gnwunre2v<XJ[ykG9!|	{4+U*l
P)!1.7`Q1L!=ZoU*U[cDT\fpLo);?L'X:6r]~
<H!qr&fVo<uZjXzs/+;kcrzVl*8ZqmOV>w,~+pv\4Ua8FuW,B3Uob1r=PDK|TTie-J=?=HUz6^1(pafJ$f4x#X)Q`DG(|><=;AR,RGN"pLCqn	xI]Ti!`KP2Kb@$eZv)hY)/ehb	q:hnZMauJ.[W={>ika3f{A7SY&%5$lVl =UJz6C[su,Lp	WSXK~1,cyo43t.lCdPOMHVN!PZ6vr~ra>]6{k0Bmx/_qhYqpd1Caln7"wLWKt3`4
%S%YumJyiFozBp%b|)gihm [gS>\FlrhZ@H/+W;IZ#?@0i'JOM[sp2Mqm-5uaZZ^q=m(aNP6-^a U
;|`M2Bp5!TnZcN\<.	*f0J7QKug75LT/d4N)'?(?qY.w-{Qv5&?Y_'0Bcd9XRW |\RN-f9h$< 'v3b@9F.U=PA$yk6"_zR_`#p	ZkZ(\]!K
-A$:s:Dey,!H:\k(.N9^\Q9e>qn
xEiT+L +yWv>:Ag[B}XQi:a@MFil@oI5^Y7D|<<8*r8V/0AD!*sC~P*ct]8vd<dO|t74kQ}_f"U]4w}<Q
,Y[z:O?G	ry]1^j`<<{|bl+$x[_"1z~}O-I2SVJ&--c:A"o>+&LJ7`8oZv\;Co,e!w)k@\	T*~mM2U-DA3X&+#gY*L|!w6\ 1sd>3<c#vULs@3PDkqD.<1oN{j7~&^t"1X?w%>5iw8~% <r
(_Xd5)LAY"I{Z*G?YK{=Ud[HGoK@[vc#O	GZ|3VZIs-p+?agAt.U9z^Z{}^`9r^gzN^Fz^+&q~n(Ux+)'p-^[;Qv;zw&1Xb[tzhyc!&raj[X=Ekg]kmutj1u~!U6W^#;Z|erjuX/];,7us&G6]V-7U'l0TS3k6fgd[{c6z.li'Tqj<roxB;"Cq0Io>Wb/N-@D GSi!|s/g HHJI\5MN\XeSQ7vXa:mRFtN6NVZBIC(uo$&N[JsgaPg-WS$}Z8UT8*PxRtW:HSf5YO]!&c768'Djtg^:xQp'gj4Z%IWBSC-2/*wIOb,E_ D;;YK\!7Sw|@.O thFUP*=$S97}Pw>3R5]t{~K"AA~k kit6Y"WV
hus$.vR[COyr.Wk8 rhxGgrLD|* =Pbw^9+SAx`Y(,~:g=`QX3xXbN=Zw$<
w)]Jd.-J<xiL9e0#wiL];L
[q_5aEXJ;	^o*vN[4"7x~Wd-<x:
%~Jg,?<W	>0iUo6\
v9T<*MC spMp v@$'HB`)(_Df~P#lx04^kSZ2,eW-j_,L	u!tY_\osi"'a'=PKSi%ic/iwwDNm^Z	1W7^33N)/Byw(l$ILfc,eoM	qP2O'HJcR4R3$zbV'+3K(fyYPNCAvdI 9sCKaWjtgyAnS%|kh}c	E|oJ3
e,m)NatI\azp+K{"Nr_)#Al$-=$IDC6K@'&qB4$%kooF--A/;yK7}2vLwm&vyAPD@W)`;C'O.PhTa}G=;r0ZX@iISv)
~K3fJ+	"lTM$kw9Pm|LP7}67jD]KuQ0}qxwUrdeDu7=9J3xq$APd	@]Om20i,v,=_n3oj={7h<tkh[#wo D\H6[EpPhRNfi*k-UDx"K)^T*:*B;(ef90C2JCG_BEY83C>rR3|cf<v/dPcUi;K1Y#QcHOvYL#eKMW@n4JfwT4_ '[P?L]yV/z9R^|QRI{fcMFFvBM187K=2OH%\YKXjC$B2<!w~9OI} N5mxPg:<-pD/z:X%I<YlXz-N4oFj31ruiVM+Kj)Q37":4)FT1D\cG|4H']:?>G]<ZD9t/_W\^J&Y0"giuVcf~FEX0DhM:^QB3m)a}K(&2CO,;dp*kt'TY'3Y{pTS8Z=+M^Dy'!]a>8-s3W(x/y{_VU|N|XIP3tpvb6-#/,&Tg.SkPy("[_=;R5=k>xhQj[/tQG%UGHpXD9j}I_GwU[!*=,t].rK"r)LL-Fxd'EG=hPe>\^]S~))%Xc-ID?HQ,3mxwT3yY"r0eP#.1q*d7C~G]>."UUT*T\9	^KM;oA}:(=CP)Z<G"|D($KG662Ko8j,hQ/",4%TQn%sM{z]dN-6H1L=m%?qMP@ta$fC}*bu%BHb2$qaYgOEfr=y^r>'Za+g^J\J5.#9fx@#z	$p6Csmt{ldBsK"TN8;_0QUK`I
L9):1/y8x<+'2$jnS0eyr"3UqA0!2u-kdWVGuy=7BDC%xB)yzU_	g.w-.=DGo=PlIO\ ]G$^uST5j}*{>ng!oJ8q6J{{K2cR&"R[	N\iAcO9|:=BmL8Fi*v\4yFTRq;Z@	0`5,PwA{10W3
xKm*d]Ue[zz[W{=>W{H.^|2SDBW5<t[Jr?\zOZDFg#/dM[	Bi,RROr`BCpeZm0\tb?_fp&I|P$%SjC@jI-P%M3y$v1K8N>S8>_:>iN)vnkSd1<JmKSn;gBSHo34kS}lk\Pz2.2gIWBw[$ISP(g-jQTBf~:%\(BcaXj"]|$"{sw5>w\V}&ws6-xw~1qnN5nECLf]Rt8B_lcWo=I=u\+6tu^h:L4-oZLoBj VXw*a~x|A*'n4P]?DQz
v.NOsI+DGT"6x>u<iE(h6A:F:CdbLysk=@1(sVuR10;4RzA5d,QYKPzGjd)#\g#e.	%rkK7Q#`QQaSermm(B8`}^TO]q<=qqXYL4rfaMO$,320dXvuAvzncjyIQs6l'.X7)e=K,W
I-F3|Km+gO)|/W_	OHv4u{vMgbSU{A#L=K&\3avM2ov@ey ?PigusR)f-QVSQ)6"0;6qOv%m>GG0@>RyxN1.6Kj_Jo.a"[	\XEZ{$B*R<,AH\*/<eYZ6_LQ=:CiH*Oe|"CLS%SyDXvs_5H&/#};r s)`,dt9SrpL+.Iro<`G3b_ck?b+ o/',	}hI}erPbQ7'> Nc<|9vy4zW[b>0Y1Z6M144y/i4Nf)lJA"z4zotwVnZkr-,Shp@'Uq|6	wqhu-F;%/=jARg\lJF<fH/zyqgmi*w2FKmv&:*r+V4Xm&=N?},R5LV3{13|>n7;w=/c2,6q$p6q	4lzd\rCh:iEq~tg<,(IIw-\YLz@`92G-ysC!0*VrPT9l!@Xq_\nY]AC5p!J1wK(@b',*}A;J([I+gR4mxCPbA=
="QP4&D|@]dfqRk^W9l;Sw'sM-9a\f^,971moDWh=>.v{R\}dT8t|`TiD05i1,GvI?_~%IU@CItC245xI/Vj_fmtEs~^QX7Wwy/JfO
R^Bnfcd+O@$/3OCo
zS%7;_Pw#XsL#'I~w+A!} mxb@\7o,NHM&(Xx(I`mo28-'{^$9huMw*KII&[ 9vQ:-,VX;]%QtR$j	T&B&_g[t?{x@x=YxEs%Vlb?mE[fVE9e}h54HQmZAj<'},{?GC~wF%:iu%v1Y)b8T>'	?X$;7?&kAJ tCUq4hH%FuLgwGyz$ZN]Zrqa&CKt#h\h#-f*NHE4PUZVY3!Y%P)a4ly9!v]UTj>y@={v)!&<d0v*mL3wWsxNq]{,M!`]YU:ubbgNmY*b/WP^KGVS)0Yob[;Y-o?s95f/,5cypsW9x@P\lUEX+)6q?H^mU$1x.8_r:!Dbwu'fPY%%4oj4'^m[O>ILXYpx@2vniv.I_KaP0p-s^g %M_C2r8B
Q"!K6(L[P,PXOA};#O`F/!J8bAUZQCg>"GY*bk'S`DP74<58#mcD^,V+^/\y&2fFcka?1s(.6&}}{\?8w|Q0-/tN}[U=XArVq-2wba:1-3P
:Md,n%fI1%ugBrG	cvW0aOE#HifNwMV6F*mG&ZU`lTe8'g/n?ky.zu*6XK|k}XuQdls2!a$vc<48)3;xoX?EjNtE"-Y:?_C7xFK}(k
pq
-!)D#&4ZhpL{i)#$8`Bc9Lel+TZyN(>'{J%&mjt`Bf;aI"7:HDa;~hxGX#%M+)]H^l&|ktn@n6sB|hX$|~v$8MnX'iB8 ??QNCMRO[[O0>CyRW+_}icjbew7{ml	iglO=#Y~E+_t@2lwjL]b\WY1#;mC2't;mQX6&vVZiVklvuUTGpwTj@5;s1,[M|s*!T6b^?"j>/HIW;e[{k|eD5q -!3QTE;dun)qss\QvJK_5
#AFpTRSPBi0${(6Z`"uwr`ODh1|Zv> '=wg~'fXiu.3gHB.]doqa2cYUrC^8!_'I2{6nugdtd?vF8!9p*s?d	e2Ta.#=aU8!v`}/e(9+6rsJmR]z; 9$8d)?Jsf()(,@?3?-15lRw=>q004%Bp$WcO
HI&&^fSV|\}CmH%6x/"Qz-o }H:BM#SuE30o33w'@YL39'52Dm:5z%^w+3j#5GPS_ZF$7+'^F07BW2Tl1FvhKdl J(qJ8-kY0M<L!U	Rl++B~:eIqA'UJ=Q+{wVaXa8VLYsE8QVb(^EX]A<eD%m!?zTij[`SZ)|'h0`fg
JSYo?>`x>.?j.^et?W_`oY;lUYa5Wy_wBqE4~{C);A288q/\C/pujp/A9&lHt	/U*v0Bihy&N>/":YGt5>7d8q@ucw=\JqZf5rocnuA;\8$\&J,T4lG1nRJ5UDHnye=~?>a;~= V}7+Hd>^+~aG]]=YTCWQ/$0_Q3wW]+$e9FI7ZxUB.JfB)s:D~%F7QG4.S_{;w=e.Ve?yvG0QP:)S,Nb5JE|nw*'BA_^jMVic 0Ki6uD&$aPA|b'ae\L^xh.4`-6\&u7x`D1h[Y0c^cG*h@\#,lBK9;)MF2?61(kt_4vj^rHX}&*^&8`b.@W)T$]V$d	Q[TH>{)H,C1.:X|MRje>@h=9`Hfw*CMx`j|mhk[+e-yr=0zK_vaVGS %@bO	n?VX5om_I:03Bgo$,Y7m{g8t
hrB&**U4m*[p4GN2nYAy&({{Gr'@)+BojZ[)$K` [`CyHH-ji&!Yen].xOKm&gml,GP(P;.5g`8Woj
UC>w}^&q#;OR?:C7 +Y_seP]U+{m`55}08"9/3dKd_4|'rW_eqct<+[hZ*yUU,d[IcuOJkF6!"Svk
sQu<7i6LdtNc-e>AUtU.Pz/> GEpNx|LPrOQOW5OUks#n n\3,Mtyk0}y#3d(*R6xl<vW:D>UZ+.7Tt`LMf'_V`g~&owf$<WA^W
R+ pF1!iR"^RI/y`Xg4OcIe7x	T+Y2AEq&[Z3drZ3e\Zh^Va0>okCPm2&iSDOi>$'IQr%(9 Q93#-PoHe%%
sr5Kt(Y&,iZA%'kamHC,O/QZBEu+FEPO}G]1W|[9oteIT0;4TmR3ZxIzv:3n*n{TwlThF>	8FL+W/W8QCNur(QewgV#@2sJ#	K|p$ARcIavk-t"b&+ac97`j/B^TYxIRhHv(?	VT89<H&L?/R~v^T,qwfmI!+>.E+S`=p@u_{*pUv6v`a[PE w{	>}",lB+eNdvtKBo<x6_zCYZC6Xt!8x?^]4m;Q?2Iy' 9N9r&!k}+60cE_/&I+I:[1zM+YixXI-.r)<;K+"qlEbZf_o@]s*-94*y7('/oVB>tZ2Z7?Cj6
uY79X]<	H8gbnvCSh.hT-\p%>]\':qwk-d]A_6c!JfN~hRS#ojzhru<^^m4@z~ck0,[cWIuU>]=tN0>|BZ[>hMJyd_u8h*h1P}]tM
"U~)
]IRcCn"J0HYUqGQ"+_w\FOnho$rOg+Bdnt)]<U3z{yeO|@=n6	|iGY`FH	<3ed%?%DE9p']_|7#vt[[/w0fztd	/`iV-NXix~@9w-gU`2c\WqY>S<p0^u[Qppd9S
t4+\<*j9L1EY,uR?|M2N'at\F(3"bkj.BMviB GY79\)anIwcH~QX99ewZDci	%]wf>~w%0>tJnDc~TdSZ@S#S=zis
!V] .-'xsn5#!g^'P;&CXf%	2$M9DmR6\Lq6<8F$]1L@$SbeL,Q\l	-hID9Hl0P;r]kxLq$zI~R lKy3;%kE9[UtTTA:&
e hq1h)6wN4KHT^guUiC:'w'j:*cwA	2Qy>SCW+jHY!Af&5aS|20]Km)f]z`)Hx@=Ps7VJUi+fn+mN>[adY^++dmS2/N[2otDkPp\fTkxk67cL#'4[CB-->Zch4zm]E95=TWm<E<[r0'RsMcm%/_@&hxNdeh\091?+u(b	k}[daXj{XiT0uj=93S>m)hUY/`[a5^+j*hXUwexMZCy
6Fo_^ lDvOu}#kV%QbjgBG&4akf896lvl*ZMZ%=9H2FN?g:Em(iE(^I6|u]7ZghVQ$#nlE%L<_r8mYl~wi^NhpGkO}a'r'26Y0_[0SDBg.r&EWE-A:@VG2X6r-%!+,cW.[6q2rTp?	8Gs3B-[prp+,pB@=PoGsT8bb7\oM!w!^Ue4<JmAOzP:`;"{OKC% kG6$#_=Xa^-@(XAJy(,)6hu}#Zv2G;(zW.{xxN7YM]4\n$\EOYG`2MUm31R[1b
1XO)G?TbsIkPizeI`g+awZ~DFPHu#s9^a9v4rXhXEszR!a;OtC;JtE:P{X[aGs`2V/F+Z<s7rR*)fO@%2|S3q7=6oeH T{1)$Cy%#L:s	`go?,1]/o3`ay56994g]/+NKc)@q,cUO4vcVbcM]Xyu<eUs/hjInvh=?k.bp{eTd^`/d\@u3va&%,OCL5@R@\hpP G&?N7`dk%}sRiJ'WkS>wqS%%,a},DbvZXYY<9!`LMOKkc@H(NlvKYNkg zNPLvHOp8m">Jeg-rW4#ZD<Tp*-6O[a[Uii^7DrC$Aj\c`)Or4&2WvOHRy&h632FIl(qV9=O(R=F)*n%Uq!. }NxlUiiP:{.!,]k3JL[uu6A8MQ53+Qj1b:U"^y"pUiqas(y?V$)Dj\]otkm =I@O"zktkJ6dX9%~mO@D2N"}; TVr$[a>o3YLt5k<7(ubQ2W~7g{%}nS!nN0!M^Ltd0DL5)&CViU2'NE(}8??~0~	T',e)%8o<4H-:#v?|%(t7Z%j  9PKy1&?+{Ht{EvIzBwpp0+^SoblK[{$_*pP|?B8@6vwHHws24h_AZYY3}>`']&4Oe)X_:+zQi+*@>Zebk)V]/#saG=XrM<>R!!2&G8@t@>aRJfqw	vE@:a|w#kASIUd:o*Iwk`t~>s(VbLK=7*<PEz7,{P5MH]M?R:LDR\NFAX[4^} DyC{Uxp+?D|UP&:!ov,?.(x,fb#=&IrY86Flu!}Ru&fo"Z}0mDH:F_x6GB@qkVURI;ZQdkUmswxF%}{C"ZeAauxg6wG0
k,=6!%(KM6<V/KY]Kc}SWkB_C4kt`Bp_"31G8U)$s(s*:^-K*DbN7x]^FY#lCz}d27uO>'IlIAJd6((+##wY=K[f-rht?B(BwS8AxCw"keZiJ{S0jhWc-Z"GP"*CUT?+%~OI_}4@//3(|$W,IoRF[\4CMC.}jV>,tkU@1&p$Dp=pBksvM7c\Q 9IV,E)59n1gJ\sEWlN.e_5o?LO1RIaBSwUDhf2(RPbN8#'t}=&~1%Y.2]Xk
4&@uRtHl(m'EsbnLZZRMTO:Z70p~w_i+TFr"0-+B$HjDbid%,
Y|K-[c
!6X8gALC6J|vOSnWF	^"<|lG
fEseBclG
i.5>_ BfXyf`QJt2p;Cs*+y(\wz8L|<
6&x1-{\ZEGa;ducM;y-yS`r	FkU)3'x3i#{iT9-N=A^Hdb5P,dR>U5nsYzi_V]9tW\ef++b/ T?AQ\i\ARVLUdp_l(qc1=]v'-wX'z&|jvw-:3aX+MTuYoq"j8lKkCX	3D!iEE1' DSGb*i<3#c=]dQUitKVuE-Bz!GC\&mhk"FQ;8gS9Zoym_Q^x1kHHy7$T,A)G6`.$NoJd#^irXMTmF64>wbEOeJKC64FHvzCi0oD0hMT4%\/Id@bK)f<'@znDBRN{V3uC[+e&u+yb+N!\YU?)T	ai-LToHx YYq!S,M2\Apbp'km-2VN=>&MN^n#6co#+d\\BB	m3K&_1{ghw0.c3h	REI.H+;Gj5Ys2j
%bcf8]9a#?57)nD6Vm-e \CH{qh]J_h{>:t14>!lcM70#l6_RAOURS%7^+wq^Qpn4~{_lZ)VWdF]XaH-*=Q2q-20cCRkTw9*,R)y`OAJs)7(*w=`;p0_THO$7^LS'bL?.O2hvO}N}qS]E!0Z:zEdt
1DeEF38AT >#PQ)|$.75x2g4v
_//pz@5igzqF
	MN
t;6`[W\jV.*av<=*$^h78Urbm(B*`0+JIh26UsALUMGJhE#h65ET1Y;K/+%<4Un)PguE2|}mhdv3,dIv
f&Amm7z<]P1\X*Q$+%; V+P/>(1 ;Cy#zN PLnrS"dM0w0^oTF.M[ny)uTy_B}m lVnHb<pSGBaQZ
1
 "	7;>l+IW=3bJuE_/]12FJ:k8-@1x"Li1"{}1}S=#/	AxltVcOAlTu1&q7j;L6hOEPPzX]=z,DGpg7^uULVSTI6IPkoH@(Vgcb|zcL(J:b>O#a0_0Tl7l6U6}m7RAORsU]Jr>jED iU7x`gj>='o:az*jm2kUg89g'GbubsL>kS$A{5{%Wl)gixlTe,bhDgEm
hR~<0X|P[`\WEDs07QzRvL=QS'.k}%Kv:1@=gtFNvn6PQ55&^DJ2NT0w;-E+$jG.#!h.ZO$I'td$$5\h>BBicAzp%dG].`xT[r6[2#)SFhq5\T$15z_["oD]BjoDAM|=u#{V@^]r,T?eKEBS*pN0Jzb+_LDJBIa,7	Co-virO>pfu~J5k
p8"]	q61~09Z%>Baq.4z!$B5QO=]^24:^HvA/Kx%zZ6ryLF3mth#0
*%RU\wIA@x!&@YN/.Z`WSH=vmP+*gY.#nh9</70"c9_g8]'?,VwQ}oBNx25]K2_8;8[Z,x#h&#yC&B5#v2PhosZFg|`Vm~qTBco6iWoft/2>9s`[r "q[>aL6 6=,#'y_\U).: X'Ry7N>`<=P{;|Eoi+r-}*xt;o%$	wCL:& "s0Cb4l9YE3bG>g_\T@~p_e/xI$8 CGS zE\h
qZ,Fm`=mJzS^?:uUb?A=uE\i/WrmB11@v~C	@T11&A$F%,JKna8$z&'d	ids_?}AfLX>b{@6xl^M7axRvFQ}'{DBcrw;I!9p1'&$7-Rz@_jfsIh3~|8+J2t,0~r(kOwL_&9@Ae&r.E"c#':yAQ#QE)J/soO"TH7MlX,Hfw1'2W)q#Ys2;m|;&i;nW Jv>Dk.7i~0\xHoC$
xZv$rjTVsG}cO!w9S?Kg3%~+py0:?",,k~s|.>THz|5p1%L D517(r!S	E[=>+P	jKVJ@=*TdD }mVRza<\7d]vY:TQm(};8?^$WX$8YH/vCax>l\3'pszV$K:/h%awh|	)ngh$M]M_&tFI e0>dvEjrRFV\q`74-XK2{'HI.Ly9FW}`91Rv.(	Ae.~G.0sNQ[pF	^acQIg{Q)KU{Y2[@4/6QmMN+~068+IDd9g.wYU8*}yi_{ l9.gW-CH65/F&SzzX]V6Ej<+$BAkY",9Fx|X30oJ@_m wWfCg
5hoK7:(QxWSY-XA<t$9SU=E<sR}ln=cQn*cLXzjK!\H&z^?Y2UpI.Ju"E[Rek6~gm=t7'VgCAOBmR?9YAKKE9Irh"UFAI{|Jg'x+{:0>O[G]d\3yjG0q|5}],hgz'j@q(sC%\[GR3hf3B|:Y;']V2Q'(N@k&Z{q-S@#y(xzI(=0+
V% #	}\=eEv9}"Q'cfyRNoP+>;9y]Q][\3ivD-,;x[M	nN%,M5h&RBNGH'~Y8RN^|,CLSaCx(T(w\)tEB]VK<-gK$qUeTaLE&qVy-Kd.G-O@mY:6><%MT<ow*OR",@q))lsJ+<q}	Y`q,wO_vuyB7A-IN;6M_vX(p@~jeo_%IBjQRkk1[r/3#];C ~bZxQ7c74-!XHDg:>M2IsTl|dVw<]%c{^KY/pC:I*9q>[hmQh&&GSd7d)^9`V2}aK:Wa[=][cnDI[7T=
YIUNKfr`Zm[wu|'R6
w2y+<8r#c|l44lvN&\j)"K),Y0VC1sC^63gBs<iShs^s*8^yrW
'Oz!0n8u^R_.qWVGfsR' Vg->[^7f4a%-Yv|",L	yK=^#^Yf'M57`B4mQ2M}$`|{&ddHP|Tx'U.W_W/Ofy<T=?+;jKlu=.#f{b?[4B'Vt>;==5X .E<{OZ3n[*]6jJ-8:P#M\iA"R[.baAL
(5m]_	vjL"*GOAv{B.h5kuSMNr,[kByO-kyk$E1"n(E,@Z/p0<IWs_QB"x$OV2<N(gErd|h5K2ad8)@Bg"869Jr&=K\_\cKk/:k:z2<M^Bww6~+/YO@|czeD;,3AF59dEenG37|p$:	YcOagtjPG9HUO?M4sHr{rcQ?S?Beft-Sc)6r#UI_BRYMgUrt:6OdR0.Y#@=|rZ\)9t2h)TCBy\B\
GywAIRNb4\)-p'P<vE2wN$4z"n!8`ByYt
Fs.\c!q!_> &nw4LKU#CzeTUXa'Gg5f>u* thqD@^jgwYl2gD*qImH7BMd0gOf#s.LA+hVxg&/&qSP/A
ITn5#1rWH`(DR:1nP
&uzd:._".gq59"ua%-4cX%&'ZO}}UV(YQb1c4|CO_*gU=jY)JqFek[$^n]hL(=zFmBVBhRn:6'KOdE9I0R-?s[RGU
Y*y1EE~#n=\j-PQlD5Cy&tD1
2o
%,I_B;^O::bFjLl=NqJ`)^>;J`3/- S)52A;KK*-7##`~h4j,O@HVXk*N#5cVD+p?iO{q35WcLa4DWD "/m~T6u44;w:hg`z%lk@%oGN%WcKC ?m1B vBYoI"9/:TjP|a?eTtl)dKi
l	zD:AF4b<BjsEyy\<bxw*k)vkQtHQ;b$ZvY8>$]vmB//z&QA^H0VRWb
F-
?Ul&ewSeonQ=pr[b}|,oMlmg!h{|D&w&OWhLS\Nek:Y7t2jK#_GZHX-n\hIzr=z&H##fOQ*e?=nPkh}Lm)#F\0(m+CS%m<~|}44v@%!R%a2'7yWE0#JLNd!)G#	JR{YDn+tbm1q=OfR2(PYI8?>"~.Ls	 2X1^0Mgdq	zSwW q_{-	*#m}-Pfs?&ehfm*TpTEFy0*kB1\vCDsZD-|pug'4%.ShT)kf^NY-ywes^NRF/$3;Hk]9Kx_O8)_9>Em'`}ZaV(INDviPC"x`Dh6k!aU_8smdUE*SMt[cd<E`;d;7_Q =)u3yh,&Mz<)m%F]:
. ^Cm>C"h{T~f')N~onECw8rXaE{B{+J'KW5i+<^$p4*F3YoAb'K6/q:'Y5'k%HH_+=)FWt^CC#jgw!5&I}z$5z.K{ECh@B!%uR(F@ %%jm$1	W>;TsGdHar,2A'T>1\*x94{USosF3NZw&h+yW}m
l<RvHDBGd);Id]!8wJ][tsp!I77XRP+|UFwc;5u{~5x(T"wNMsQ|UmL/^r5N<SJAkaJr~^Z/a<#v`(]cYHA;XW
@w_IESl:#\fz++a)YdPE3]mQ{@8F
rY)Bi-^DMl;vN[*z?xZ;ZX0hXmX<WynNNcL88a>v&89bX^,'0ky{||Z@C@QU:p-G*,@vehmtI'nuW,D;axDyDz""lwKl`K/JRswc\^UL|Tia9I[lKBU\=RGsF`d8[6<2U=OOFU:JDfHWjE@/QO.ss9,-b.	S{IT/K1qRD$|lbSy|\]NMnY"6>pM0XUwT'TKSremYj=[i'i1rm@'@=Oiq(a#rGuZb%{s1!v?co7AOn*p	3%qTjEm;#,G4]jp2L{0%7."M_s~Z+08*CiaLOW(mfkq}BW&7YXX30O_.J1Cbq~wfn\M=7%w|V<'@)Jc,@FR&Lq>[@R{	E2YhXUk\Ao5#l\@z	-G/)pfblrngN3Z\QX]J|{s4AiWfnDh{i.(!SAc/K_zastf9M4Y\qc.@','gH#vs)&ZIho9hxJ.j[>z8UdY:R/>nY.C*8_MU.YRR|(SJ^iJO%ztQY*AodVsqO)v>PQRAL(	\l1)J/{jE
DqmGbNdl1Ra|?@%m {Wi|loBo`"VU26YwPO7VmQ1O<6?mVai +xS5g9k^#;I3_Db;DRziYc9C>.oM @e/H-,'&J+vp$c_M><wW[	)JeK/;[d04`rRLARd#]I-Myp9{;>[XA@jACrL3zTfF|B:ljCP2Ch]SIE/
JMJ6&c_^DjNjo_Rb~Y7c!WqY!IL;zC(^`;]V01<A'2d}BP<u&n+Q<%?2u~4-a>KI07.bv@hu!RjKSy^3"'<Fzm=wos#}ClO]0VIdP' wnG0v+:I$'NA"]ONHb2O[9=@|i -yVAA=e4NFj/FOggs.c?Bn51Klnqf,aE[n15Zsz`v@R!fB+C+iD85$Oj5E&?M8N*	S_EZTf^oVo-;Cbd\5S&ZdS>+Zp?&NNveMOmiJ<nf&I!o~!r2r$<
x:[7A5pEfS9#HNtt@:p|a=G)I@(mk\	\L{;4	2#U>Q4_|72InS,S4R,Q[p	xj1BnA:<H[M~`(hcn<o52M+JI0>.y5zcTtHyeSVkO6R"6wF\3X\Q/-aP%^KjPqTB8Jmia#`_kH/}j>>|a.Y?in&k:Y#]!9bkt<eO=KD(tw$86.q8XdRy;|TT3WT% 8WT=F3sm{x#G4[kVXW5?Qjojp4z6fCf[zH7LMqoI?	f_`pl7,
|4'oZ	V80zujE}U&O/#+]l36q(+E^\|5HH%>F>YJ&qI{4;nrv:Y(QIKeWX
<1\gXOiB^=RT1
4MvGc1-J@A';aF*$39'BDg3Vc/Mz?w05%%MZ\08APS^T5q<|yAMF^*Gu'jJ{8~-"6n_&=LoaBohx@a/ C|W1{w?[-@jIa0#DrU?Ja6w Jx8\x;d=f9eKyn"czzQXflCG^X*3/-tm!\%/3}d-2`<\*:=.:ofx82G	}=5KP^o pX;LSZHKbHs1	Go;Wz_~vA"YMD|*%1tOAyOSVk!x~Irl^@o\B`a+{KOh$S^|:pV]6W(	z{(Ex{N!h+knFQ!WS]z}j[2S\0Ak\XA8>{=M8-Mx;MhWV4a&D6l/['=%k}(?Pncrt"UcCUez;<UC84)`+(i	 xKu_f`hq8Y-FdCb;6675S
aUI\t	Q+uhiSN~sIb
O`'p
iCVM9RSDXH}J=Fg7qaZ=1jtP$=+ >F|yE`4Z=3lsGl3=|&fj_F\vN:1C[D8of3^]P1[mCp:uD	w<[Q\o;[>t%{$
)9L(l$* 7P6:\u,V\[2CH-!BTDszZPM+8Sbbb=Edck,](9NH$y*b)NusLSS-)mq[xGA6mNZ&^,vC$8<9Wr0c~J4+]srZu/n8vE|;-#`5l#HbWqc{lK%Y!|Trbca[}1x%IXWJt
[[():Vw$`I 
E~=c[Dt_"h=|_xH7ok/)df*'DBsU05Nv(#	|4-}wG/a[5l>6L_yM*-t7*$cZ3/?voW<stz5Bi8Aq=)WPj_v-i?s 3_QwS'|`(5#4#S
@1nT,.AY|rtW4SG)wfwd%hu^tCJ7<'{1E8jX/:mRmY5$`COXRZOXyL<C T*lFE>xISj@9aj4dpk
ZeJY)|)TKXF_1r<> G!7sF"=='TrM%+<vJwMU@Z(k#+DbjK:fgiUb-1V(c_G^dp,JhFhW~[rjePrJ1,]z8#BapRjX"o*ZGI+9\{XK C*Abevh6j16iGx	k9Z+%pCVn~3]+7
2[>f
(O)}D#`xvn]M$mk:z$]Lb!7zwbR"<;I4>3*Xno?P{#-%[&rFj\=$M'p1Qw,l-l;E_6JaI5E1$=G*HrgNbLTEUf`RK7jF(tf0!NdcnX!b'm+')sHu~VXLgg_
js>FG)3i}ewkDW(J.Vr0qHyTYRw;xH<uGbq^wIv]U~0s`|oS{6=_[Nh'3AimR=t3+e,?C.70"2.:0xxg7U8fC}u|y@P6</a*v0a3zhEX/kZ$e3a. 4=L23?^c0HzzL1I26{nF]v/XnP}"U-	eFq[4aAR0>L!UJy'b,m*;#,uMFY<;
9M3Lb)<6G 1VKJnF0GBlh3AC<Lll@Rf	;k7]&+z"~'S=mzx0RjS2CC/XWM\A}m/R2C]7<O)hR"HZ2],SOGSi9:L3D9fX[WK`)43)-;^p@1oqu.mo$uL~|8CXnNcHly\:BAUeW
F,(9 f{;-)Znx6d*<=k
lz[y_EA7'BwbXfm+y*o=I}90"q974*]wEO%I7AXX:]g86\Ta-t)8({*YvXd/;YeiPe R` 7r\0l19W:/M*w%4.[h}]#X@iP9*Yg=Xi#\dp4^-6dvTOK`@U2p]*WW]R=EAC	vN35B[Pn!KKZ=]g20EVkt3X"vRjp{p>ZPlAKx^fP}T!suH@-/jI"/PoKU,jE]/a7*jO998QT{Q"`tM	</^PWYoiV(`m;LLB~-1qG~Ii$MT2q] 0\5'=d'N>{!W8Rz_to"<23G_m?N5ci!<\1?vORh[\3S^`%Va`}mnfUUD9[XzND
y!\hO$*J;D}lo@@pz1`ew:T	4b9^'M$k[	Us9Bt]3C|Rb"]Wn}np=?-vmLG"{on0a1;y
5.&vR3Zx,s.k1.6/[9bopM]T+V[q#bwDT2!j-O"ZZ97]WR356ny@[pBvICn{-8*hsW{y\PrzsksmVwIA#+R;N3$H[WRHi\w@5'aQ$2:*eq3K$4w^SK/>:	p)LYvdD~zAO[ '@rKJU|+Kk.t!{bMY6966DbG>?/)kokEhbG)@RH9X@|3p'WC|~%Vsdg`q4BG6dBA/}Q9{\
`>f!u8p&,-I{J6kPE
H4YU(wm%-^(G00NRD$KzOc1=;^L%*+3=H8|@JUvMBk]^~
/EO=`QFlNi
 qit<&c_~ fGW?Qe\q:X7$Z^-=Ju!(]P,o"6(+7JtL8<@:i~}+Ozy{${(H	o eb~[M&04(]}	SqsJMIf=%=RV36:7Vwq"_.0A8i'FEo+#+D+7M(WNS?Q8K%Gl&NB8~`-oTKgD%KDI#H]F$MjZE)bWqYleUU?2xdm$u{yGYM!TQD,9  ).X-BO_TAhD9H&9|S0n,/!\8'!+emx`M<V	i =t/y18N3$F?@4;n=a.M/zo+%KP]}s+"#Zhh/qP,-)ny3q"4=Om#$r"*(P;A3TF:wuZ1dUj68RbDy0&zW^
TjHNr<*rM;/Q%vbY@Jh$L<N*@tO$0 xT>,cWh]XBLegE+$wsgypRZi5@Y6Z=T=,vD_zAX<}G,}l
8-O:MgI"ksW\:rSsN		h)M@)dX$|r'C,k*[s	YD*QQoI^yOsvO:vWk.ER,3.`*EntwJcHGe
VL"8+LYlL6:!!P,%mj<CQ^uwl<mRi1YpPS]4"c/qP6k`g :7#=ic=ZoPF=HW2K0:P[	ViL,4uPD^l>ci':*DV
Fj^pY[Hu0k')x{y)&71qy=5o-NjXu:p'x=Y7L2AQYaOuDU5OK{ML|J0w/	V{-Fl8s@=&_6YA45d7S(H*!~]Uax X&4Lz#3wfqd0&x;&|.I t)fLj_)*pjG069k=uN4`l+J'6<x[jZ!ITW6n`^d(dF[&)6+~*3>LC(v/[
$!*^]#7tsk=o g!O
Xw=TFe(dW?xT#H?8uu'#w ft)O2N"smW{kJ#I5>s	n%QA/J}Qs*%7E#r-F-D2Nar.1\?mY%Z{{TvPs03FvL"a[li7.+?	\Xhry|X3rv[v3I%RfqfjAYW?9m[uXpt]P^^gL`9C.;uQ]-GKzy8%V1"T4C%Bqig0wg$:K3$Hq/8G(Hk#`Z%W8q5V+.	)HIi&usRe7ViIiUn?_G\5z`~X%cIdp8lVmi4G^\HCGf'oVXQa!fc42c)VHAY@&T:&ujY8 5e-"0b,V/R.A>(beMDx#|-k?uZ!B=(]r9rxVt$GkQXpq'tkdZfl@o)a~lT5w] eQU6(l UFcv(1rki'LB"Wa(6a^k2+,*q]dZVa<%~(`LrhME	wEap:5W69#OAkmlS,2jp|Ou7>FbQm28*a4@?t$t.i`:2'%c%H=B!Y8)[f<XE1*V6Zg+.Ma{A=^653h6|X/SR#d`m?gO rhwUE_U
z5!aq[O9V^p7E3(9woE,CSoK_MCp+^.vBF~L4xMch-gW	NUJ%0:(z{B]E-8VsPRfZB6U'iBS$03x!xx+yRg'a{}_4hn,Fd/'M7gh.%Z8S!&#H[.\QC!;3T"yT%u8/>kQ:g*^<d 3A:6Icb 88u!G7</{'"*<b.<A}A:)W4Ol"%{-% d9`5S8ZBCJAOzE..h/p\A_cDH?#+YV5~L69SSVc/^CEuE]Z)H'0iH)(h$4+Z*Rv|%[=5ci?_*B}z$b=&J^O19g@x&tDiz3$/3s800"<KDH|w1VXwK9EV0_0k3o?1-?>I>'&[mT4M!M7w+Ebo^$r^+Q0Da@3IX'XyF"{q\9C\M%erdYF'4!9i~Z-F>D|?F"uUs"Mr$1+G9`^/*<C99UjIoWkgTrDTk/"1u`r(d3 5Pm[a8*)v+U>)W[>tAVG9w YCkBIKyM?~i{Buu+KAw(Ct|r	Pu{,Ps`?nJ"z"}Z~+iu"S*,`mBAW4`~@HNra6FSS9 8W#qau(}ODDw*Dx`HkJ\*A_'EQm
HC`+$6Gf+;
:b6mRG5p<hF(|I>Jwq4uvL?efD-7xjKjpRPj2po`WCS-JO|E,(@w/V,9bTl#+mLF\'.EdO1)K`^`jR'S%y`CE{&!OV)v"Cy5vP/+sDV?7ano^("rt.AOuZ)DCl7$;(]Zv89*A}\TD;^s9nh8k/v1Vw)`JF[\0KKL"$ D!~f'"%z,t3N[z90CR5g6abyT}gv01T,puQ0)VoE/;x|g40w@.<<y0VEV*w5Y6^<#7.8:T+6OS@5;EH<d"V0;<Ai`Wn|e	+a%:^<K+KT^[wP+'v"JEy}1#t+,\,t;"dGp^A1	QT9TJTGYE(LMSXG1[*SmjE"m|QBU>"&Rg![qrXi9]x=aLmE	.JMl~2FW1h<	4Qh-JM%XWq-C25v90yY+/m2";Yr<$LXNsjMIfBO1//FuDmj_5=/<YId(nO/;[*p(~pG^HiaV!=;?kr5G>;KN7Uq^t5RJM&_Pmc0|l-Gse
XdN'n	*Jo?"--wg_Z#J%rfV(cD_K/J#JHlC*0rl^)&)1	Hb-&g3PL4h>n[oQD!\
DD*?JJK}Vd!..8H$>0]aei0I#V#wj,M_[ao9GL1H#/REw!;A+5ary$NP0:W^fba0kwW8'PoN "*{Di7a6>l w[n6LLzT,Cu"Dy-s:w-Ce}%?H;e@gG"8L&NO9Fe;7LLrDqf7Uj:VDm'\RApkC{%Pm&zy+^._tsPy1wPF-CkW{<PkNpj}S;?vpZt|
Gd-<#y<-scX;iLc3M)0.,May|_R#yYAPf`i$`,bGXY)J(HX&\;uG3DL}@2?
veXr%[Hq
+H;c\Y;hoFzD.nWQ[<:mA9*O+Ip;Mu}*vRoL["pw1aM61'$zInhxa^`Q!1hl%ChnD9eZAAohW-TVy ;x{hse-^qMfPpi4W^bmZ+uL=KC5$f="$Szbz:wm^fN 4J:=\>'tJ0]%'VxaYQ%uK);wOG`!l :t]Xmqy]SG/g{}J\1P2E(2Vrx#1'_?EV4"w67*vK3`]u$ovh_aFLa/@GcA(d,RF]wz@1#&jRLf=kCWw8MUr[t/l.t%t	lel
1qMS_A-79t9\7QW
*Z1
*-~=i""\jHq<[i"Zj$*in\@/K|UP>z{b!GceRW\VF^hn0?nm8}-tomm^0;{%*>*Y[1[|1IkR	}Mt}gPRrj!YWyT|p|'G_JnV?&[jkS}l()?xMN(qJ\0FG6x<?{~nvFeTp,?Jg{\
Y(_}%e]`qY66v ec pB/F%i+{(IGzLhBm)l2Ti-5LU[X:}G`V})i3Y0KFMnr},[]2#9j@v!%]Id
E(xTl0t048Tc]TCn8`eZK*l?ZKK$Kqi4_A{p/T@gL+{U*[R{cgu0}4nH.p	|e.{n?9tr	gP^UHG]l'o=$WPom`pbZ<;.Om:?M^T*hNaL@-EDLU0d+iq;,[hUOnZ;rCX>#|Mi&qfCd6k*77laaP_S{or'FLt9,u G,Fhlf7S}om2Dp^x<K9(#s7V=gd]5h{/jaO:zR#<\%*	+k9;YT'DF-T+E#	?F[0</gA7Cs$-nzWNgQCN<9{q]+/2`n}J|fs"T,*HWr0!4z2~Z{&(Q{9K\bo4""^+o1+NHy>;<wf"]J8rL1dcGt)7#@GM)bmwE	H>
s^T$/R Os+#2(s6c!K: /AEGZ~Yy`0:V<oTA&7NaL+^<#]Wds	oaH%$^gd[,o5Z1o!(t(W%.#A>0@*!_tZ$IMo#4}"<!Wc	oH*>#JSp"{@Kst(I3=ek,SyA&zj%G/vhS|	8*3	N+@p:wF:~[;hf[7jmn;,F[.1ucsu>`M5DMyD	mZ
5X:MODcYvy7Hs^:QF	R pG]W;`T2%/&vk&)s%5paI!`Hv#pZ;1qcJB9-(&.M$S|{#{S%]b@m"-+}P?!Hhe$I7MR}z7Ws;MfsFUSj?(gL3=MXMt`C!}%i>ZPfPmBB{9/m@-#I.hA6M0I&igf& HWT:Sb?-ed!)1kU't5P!Ijp:6uD=WOb~_}QtEkct\WEADgx?iO|_5L\`WjL5E*P69o(j-Z:$r9deAdJUBU@08Q2:/`*O637a}a",#N?j\|{tdeu\DUBqiA	<v:'3UJ_6=h[cw
JwW'wF&&udyQ"@y4EN_vF\Hmms|c5N$-c]^6dV8= Gu&_JwR2OcPyTU~P )n8-eapy$1	3XbukwAVByIsPzZda'nw5''fn&PaVQS?)"LO`\%Ea%$]4Eq<8{dak#bd1>iw<6y46b"=\UB4GM5}Q-l&Mir:YlogV.Do;7!0CkI^@~M9?$R-/Q<dZkbmg.9uA\qYzrB:6R$"Oe:OlJHe.j]ixjg`jcYR-,KsjrS|`Q#qt)VU&xgUXiw]E@"X9Sx3* 3wiaz7UTqZ/W5;uVVTSUBP}Z/H:kAA9*id5y34a]>BN*#&JbV@6yT	E{kpO'Y}@\X\kd?F'UNmmCnjIM$a
3X9ddakFd_r?#4BJ,1=$C5x<JC{nA)mfcc uhB|I#xvNi2K4I0_+ALf46TysWF@MTgZ=]I1+i90rg&hGR)NN!C]fkpO
S@_Rt4]<pQ7"3*bT}-[{}W=0iODd`5T;HAGn8B%HNtr	.]yX|!uC'D2#4_umPe70amU	BE$7Cdg1z,yW1E*aeE)*$Wv4p	.g.nv7
tbw&Lp'M]vs$9rLdY~!3ci>_4+^ >zuHiNbC<e/bj}:%X&@Z*]VPbLs)&Fx?G#zUSeJX\9eQob1Jw%['YiLoe4G$Cj%%:!&lRC3=q#]rEeGa>SwrQ<1ic]FDp!NSFV"!}qw1\*}a@PWe5D7S3*<n)TywqRv2~fp8], =X\}$S+hISCyQ%,@C*
D{;oWY-eH5uoq.)-:r?a<4}fa=!f0Ft[vV3BE7h	W7+73>mli^yNc'F)].eQ\BGe>.-}g%mS*a*8M|gufo*JULq*#!gykVhWGvjUBlH#)1e5$%bmR.--mc5AUFKMPyG@I]k:InYJ}TX?yR7,T<{KM4tAD6n!*[zxO<#P7T:ac~VVdw\zIRQ]+`D<>ph0t0zh>t7|XE3X&v$WZ,#S_Ko#nan /pcW1`+ ?z}'Y=K	'iZhOKT`=+Hw:s5>XMCEKTw,@Fv!Ru"vckN=_YU.2iorL#'csI$7YBT?z|?K6[.Bko'M(dd':@d#Y"fa	/Hq2RtK0pvj@l}f?vFG^WmZ}-jqoEE6;=1{r[H,:tp#nSn47k3]&@ZT+T<BkfvvSnQ1@ngG/vQjJ%WBM&/zC~hgDbQvG$9g.S uJM91:1;&ty"/gos";?Qz2. sZ\"
}(fhqYV`FA+)*KlN>|0X()sAi)[0~T$g|N2gq^bsuIhXQrni~:U_;LL
RT.k4J0~4!=^CP`;_i\Z8;ETHou_fqCWe'i`^{;<$UVP"]((-&fFw16!:=)4<3|OWcRr,Dh<4DU 06)HFIKe%_]B1Vvdcj5//v?.My(.]#Tb~FYR{I?Y6`O6AD]!~	&O'J&J(\uj	|Lp,1hNrQ9?Q6q_M^~n<}FIOSeWQ3a#F}8!}s	tqe/40)_G9fG7?M4	`&|R{R:caz~d;7-ctn}0@eAu"V)73LG5X3\t_U|!p&~"UX9e7'W$ tkAz
tQ@Du{eLr?aqE!0{i,3PpyRjwM&(iT_U,gX*~v CJ1,. g9XIyyoe*o5k$	w}.13ZLNv|!M,|J<L.>G<$JFldRZ/
cMc8cTkZFa:k'&e~(BZ!-@Ah%Fvs"/6T!&q	0D4~+J>rR2@YM:f6
&~>g)RK~D;Ax^]`yH<2*QlZ?|&.gC7S{?i`r|
bZJ~8/-56	?U9l:]3uJc8/YggoXQ)G!N
t4$,{i mpC3n/VBbwX}L$i:!9=a7-C.bP>7.!hI /UHf,4UG;d6jS t"LXr2/Tt?Q;>qyBI./8yBbaB.R}oMYMDQ	d;QF/@Lg_2,4GF'^09bUZP}`mg(Dowks~i|+{:q"!)Q25'&@5cwF?KCAf@yUmTl#
1+y[k#zrrAeN_;~lkRUD4!]uU9;b(Gyi
#GAV RC635)U+bX2e3}fDj[)Y=|#|=\#sB":V=).$26k<3V;YughURQz +ccgI#HQv9!&ROMp_}J/P1Lihb!6KC)IeFPPGYX5j
SV|TsiDKFDV'?_i^_(t3^2`MzXcA.bpz]>@J:\V@Ug2!cm2e<?q :)ml1U/%UH^l}X"lCZck~yKu$I/m>*Lx0Rl2~N%{8Y	%qv-'| pZyHE{J>#K.Ge_LHX{wNirV|o;prU,Km(E<{xe}YbHwq,:7Ss$C49]RO%a'G{oec&W:rSTu^-}~U)	vJ#Xg//i`Yp[aG_Mf*}64fP78E">^#t7_zF z0H9w|Rv=U7{Ha`vXh3V,;Vku.jkFT$?]lj[y}|WN|5X)DB.lE=6}8xckV8$q[1xQ(L{*z	Og9u1xxv|O'TkOU7Z5OoNj!$V#z%[{(RmRwKYq0K@7?7pyOC@i#X.#F+>Q!Ap]+0iuk445}6d>erGbNCo0^1u$&RV[=%/-	Sf#O^k(P<-rZJ|Z<]y!(#D+ucI}`r}].z0C
Ia"Q+m@exi
b6G\_l'~B`NQ9UmDA
4~DBTtE$&7e/xcIh#>xlX7pZ"^Uf{H!ei5Z4gpfYe@d2\(8a%&GH'n0v	Z".rF;8n^dA,2If^;5S]h7xfxa${
_tNz~$}!S5Z7ZG4*di)fwH6oNIbxzoT?h_GEKe.}^QEza~UO"ZdB\v3Mj_\nr@W+&(Mlia,~i\SC1$>cX|uUSQ&$v[z)lwT!YywS# +RN~S:%lh~"'E:#::RC^G9w8HoBbc[:h#	s9yEWfB57D#[.2y 8&uZ18"}3go[[9i~7z1	buOj?6nP]3%IFG)jgS]]r8ztzJ6a+%H'|
A^hHLKqG|zEq(D{*]T]jt%]tJmNv9J3&'I^:aT42Y&O.S.V!KCrX8mzmjq9F[nXrL}n+t#J%fuTBP(M7SF5NA-6~r
[fm3ksl}U_#+NC(Idj/-B[m0`{0Fr+r`LWWAK'10T;Y KI#!s-WE*8E]>!-0vrbcAhB@G<}ldUzCE]%aE>IF\Mj|eLSEu2NzL"^$.rg!63D=GnAp\[4Cqm1K
w@A&-(t PNNLfn-
0(J!K[5aoj:R\;Op.GAh!q`kKN?xQTIJV%?2?K?1oj=}
!+_cBgLR<DMxRd,yiK,'6g@EKN@qKi,+SEd]tj$Jn=Bj2S(SvZ{1c_j5bL1D;k)gvor*RlL`6-tABRQNn"GBar0,KX?4!7'P_fx,tmWED? -Vh%:6	z,ET)09dV$
JOc{Vl3qV`C'tkMj(02Y8:^_tP
(gXj WA}}@fF_3Eh?,qO1+H#	qx(tf-'lf,`mJ
o@tG0 3cR@qX26ClKFo6f-8<\`LN'McLCG20/`p-*3ir=z<cr9i:aRF X8S_~m
/<GKAR ,.h#k+ZK:#ss]<N<G_4clO4`)HhEQPk>(g}8wQ>d7s.~48/#GV}nk	J9J[,4QEquF)8Wy_xvJxS+mXUXL;28Yh5=:{)@MtP)gPK	rt)ARY<&Rq`=\#nivMOW8i3M77#uc n/x|BtWnD2_n^zPOqrN+T)u+5+(tkWa\u.${<Y}vgt?_+m[Xfeqi-@P>P}#:j>~TWy,i]vm@
4HE0q8z2gH-?-]>AXE );@e(@]aDZqTQ(apyA(t/W$zl4?xXzAA;Xa06PE#QMt&E]u23E|(b9fH T#w.6aIh
s7+Nw5GSD@3sS4Un-OcO:tXN 	ve.wLSM.vYR%0Gas^B<A?^T(:R[H~<.sf*qP(66#+Ervyluw/axrZ?`Q/=i<PhU%$-fK S9-LeRmK;wv`q^"TDoQniUw6 Opsh:UDI;
!K c.2v{Yic|gbDQQ:Y--^%3F)OC@W_Pf|,9WgMO.*bfjC|H^_K8OG7-6M-FK)2g^7DVNhN@AT>UOlBn*jF~iiL"XIyjbD[^U_xe7mlVS*dUaP~>W9ALHH/`r|syf)AcLcz|}0:1nhKa1'mhC\-W&x&Ri8;6
&w}a`F&V!;]mJ.C'gD	4m?ZR.'/'!M>q*_UP	\QF&[Z{8-vrpV8AHudbGSCW(cFE?$NW]t @zo,5]2 v$48WnR	28o>Lgy-:sH%kI,BpoCT4<=2FSE^We^AP1l|$!*,?y+	Da,]-*8wT.%Len@lc:jUV0`wQnvFfaS-@NWR3:?a?Be|>,sT\%t,ISbW1*o6BovFy}p7W\+[~$K1-QjDpibeZ*@6HsfBIuKCkvgWAhy!Zh/O?EZ6*U/.nF[{D`CrFxCzZL/+R.sWWX~!J]IpN1V@l|:Aa
Z?i#>a0olL+B/+SoE?6mc	E_Tj.37Zd8(DEW*x;2=la	h<:Q ~eQgno(lR14;iLWEYS5NmZ6%$=2	|\4Bv>Nu:>,S:@`iyj}'%o\;M*Q!pW:R(E?	MQ0~v
*Sp.c{j<8O>l()n	.i
6B&R^u#@	A(~N+n+.jn/:MXMOv@aHJ@[N~5=
Dz!^6Zffk~yRgQa)1UwQwbjm=8HC]YM_[l\IlP(] r!4Qj/SIGdB9fd7DH[9]F9#!FKz;B:au2BecX8*1yh<C!,~GkZwlHR6UIE<9XYs
1aXBL"rt\
4IRPg?.!Kc1v*]-L }[x3waP#Oyg|6Rj6^ejfnC(%8CgdLj#knT?=^6@:Pify}U|/G\/Ol^x!#	^HI=+
v-.K%TP|CkZ9fr'o~c	<UUjjf[:U,;C3G'Wzv_b,!&M$LfBCzP<`XSctY7CtEarh['ED,.[zGdi.="Y!mT;sW
ST?@po	c03+`^uSf{9Bj2m4]~+Psvj4cJDd}6(@i7h@R6x>vRHh0k{e["`*KRuM9]940"-RhIhP<Icr>.8V2E"(uC/1vX5Y')u:
^ -
V6>I]Va?,|!q{}[93 S'H*xGiV0X06XQS4G[d&K*6t0p8@guzG{vb_e><=W43h0pXg}aPy./\-*oVf}>"U<o[5$\X1fV-uO3c}'n]c*j2XEr&3FQqnOZD$,'`
H2=eLkzw]JpZD"RQ7)&prV1U7(1p![YUMDlD \Zc$QtKhl5J%rT0s^5u,x]C"	
Wv@d~C-!*n?]B4ZsNm)14#o$hb57%t^=*sP[$K`a;("4]av*	15s{HAw\6(h@NXAQ%RF%6q7kefPv(J48$P1QVczstM]NA6DS=2Tc]k<+iawUZAlXWPZY8zKr:_PLkt6%TmPR\i:d;um!XZh)<t*
KAg!LYgGD23/sh6dm]ician?6UOgDj1g37}Kah,=zv5"b_.U{?%&/"^@V>}~W2^NwMWnnPsdqs<'SNXACCfLdj.u[DGgx9PH_KnxalSF[+FU	o	"Q.g.dDB5Bpf~n(eUR*lprT9Rge?`HSjY
1"+B5\s*tOl9ADq<L%{<9<~ {0: >+h&OX`9k'h$&a^xu.W<UGdE`J8q[Wn<N4Y]vaCWaWj5Hhhk}>&O l hC`jxe8^=tKn[8sKcF#$zn|\'zNsr,\WSB<zJs>0J"EMpGYXYgxgjBJ'EX}1sW2T#2
)v-"^n_[1'#&Dr3:fy_#I<%t5@mM:HF#X~^:-6
5A='!DNq|$A/?]~u_G<h2avL38},f!D][!p<@^JFM]9YWYw/6H7BP"`gL>
4/nM07BTV2HIqa!`V%(/kE{kbqUgIz6"5]IMvyyoY`9EDK_vCy	B	gLk{\@[Z3p^i^gh uV	Aa5`H@O,JJx*)tXWf'jp7Dt&,6znsEc>> #hq62UfQ_	yn'Tyr\no=qdP6F@!>'&&QA*:!7sdgvxnBxiI.*4>_a=Cv]Mtvr`!SYjs0HElLxtg)#n8qrj_c[(EBH[Nfj1e>o_[bpc7vImN)`bO
*i9;/N^|s	/T_G53;b0>QGl?gYaSzj!omE4ys:^O	sC_~6V4f\C>0TnpLrk_!zX(F/s7a\"V.~^SF-7v	W$U1+t]rU+-AaR0u[8$+pn{WSya;A ^()ELGu3c[%z^Jz`#kY^8'[?2n{>VR>dU}28u4x
6ZQoK|".z$Gfb3'sl<Ner 7HF97{`=%~h	8P+Jz\KgH~re\p/NGz=|!MT4g|ZW\Jh9EbV2jPN:9_Ao*@lSHVnX%sA`G~N+I;neCmS[QL8(|bLM$hzq&8]HnY<t+q#2]}-#s9uY:gNWF/=jGyb5'dNs*$ Bx|m,{P
KnRrorz!7/#22W
Q)ueLte#EH*LI"47kd&HQx:lk3LCCB(%CAcWhP< p+a[D()\7(A	;NNsJ"mPs?XdNlKwc5OUhOguk3$9fl-}"Ba?T~=Y9rO$_)0\
1o\iC8F,M	9?.o!>fi:cE(N;#Ix[aD+<0-,Xo
GR"x$CtbSPisut`Rg"Q
 ,sSs~vb<=JY2$mdRe*h~pe3
>>Lrl|;3U:*;:*=|}5"GKqGh.YcY%8?D8m`YY*cbZ^{W;PITcjm:Z["\M,9f%{1X+K-?2zr5f4Eu$*IU|:JDkvkcm )
\9HG7BF$p9z{{MXW=s2@|G[t!"	60p:YC:NjYx<4B|j^beOZ@y=5//&] +|
TDTVRe%UoK	R<7I 5?.7,R8{3;	>4V\EQ%4#^Xq?U(;C%rh@8jJ Nqkh$T)]5 QpBGGGS&*A< G0#}pdJ>_?tIx(2eE?mqhyy8w3LZ8vD-}AGr`K|O
ru3.<M*+nD
VWA&Gj^H%m!do)C4+6,d	8AP[6mKn\du/3Qi`"t[|Ql#[Xn	c/+D<T< x@71m0<27,nY?w[%U+Z}'Dl}Xl;f"TWsHP
M3EZs<	+eyNETL)6!	fxiq>hxh(L1}/1*BK;|?NYQ+8/KEm^|)yHKr`a6.0.Jw
Xu1lVR>?tSY]i4:<H[t&nhAQ);BwhvudSooXgNx_ZkA<tfCbSF^z&ib{{[9ob6P['V5z$Adq|pa6,g6ZLRq0Q%*`8
37OI=U<H]Df}^P.,MFvo&r5j@.mhJoJ4Sfjk&U=\
ETP0Al{6|fVQ?":Xn*FUe#T`i]EzM386 n<1@W-{Co'N|nCCe[aT-]FIm3BwPHF4P2oj	1=hLy6rj0L<GO5p-
W Mq~c_6m `]le:nh+LCLr0]9?]'0K~E:*p&r,"S+D+R7DJ~H$n#.oV;{l**04\Rq[,u<dV4OFUCUJ.xg3 Y"%ugKJ	Rs&1?=1$rQ/@h/FpD>f]AnY*d\w*lc_^J^thRNEG3@ksQhLvY^E!zP7|M1&fQ #F:iURCDmY?8x%FHlTjm%m%ewT[u@L'B4@^^Fd1yA/b$	r'vJ(&m]l--z8QPlYuD(7'g"J0QQ=rcUoVOvL
$.Gd,.Mn Ap5Qd.rA?pH{l}|FbHpk`2(2Ay%Z_uI|iT>B;cDUv=cBNfM.y#0L1 MHVI")p27'\.k?)v}8;>^&"v ^| 1D9p(({;@Rz]X+kt3k7B|=d;q>t[@cSk06sUA?YoCwq9Xzdkq"wW9V}[#]9;<o'P06gD)bHZES@1v/-74{&H+I@<u)qz[|Juh$@&QI9U5('}QR0v>?&-6Q5K0xNPy]2A_fbptw4^ob+3zXnS}#CB@U&`8$6wl_e;tT&<0CEVmPz6=EiQ#(9,APxkOCV03D%:1)T.(WVFLguK~gR)vo+$J[f^2!B_NtR,Eo M)SU|eWmg9zj67wEatO}.EZEJ`c&9XAz}|ty+n$g'Ki$kc}Wish}J=GaAN\:&_NF$^(GdCDQTjL7<g]~9=.a-Z3ar)1)ua7T(_-GUe:K7UNaToO'V?vE-<V-O61f,.:K||stbu2=~*F!7\#?7J&x,w[@3`\;za]_5r_[@Y|oI{i=&-Fg"8 >&m3OE_d<N78R<9Hm!BEYcRzH74y6rEuP"}O^/Pke:=jDzy]td~E<|Xd4%&N@.py,4{
rM9{*#( ~t$<o9uKb]j3LWh=7Z,(HxvN%})j}PW$Z8s
v\$t!-(_? D^{I}F$?B	/=-"{O<{jI&4iD
QuekpCF<5`[Dfv8[uXItVOI:QcVUbK%QC?2ldc4 S,p6)'P.+9$!
RKIDKTQZ_4{Uk+g:y>/e38J}Oq 2b^%yvT+OJB_X%#W1Ie/q|h59o3H{Js*;c:,q6bp&dd337ja{iOP~*D8QO-q?W1?L1fNN:P?[as<IMD1?)N#Jh0."ce8;xzYKm(eCCT*r)0V|`w)~Ts]8^`j!wYoDB
9*5wyQX4s7ki2F&"v'SM7]Bz,]#E1oFJB!]Oh	mo	R%k,aQm'/)>A8ycDN)Kk^E!p[>_>4bdf){L,4eO-3`>K'XsdqUo\7.['bjmy#,VRZh7c&r`bE#3"g'w6*@k7`TK_>gi
(,}Q)KQYO
;6%xKgU2(5.*"_/#DC5l*V@|J6m[H%<k~*IJ|0")CV}tJ1Klxb`zhh}-*$.US9<c[0M^t/*'X17PyYIR/,g%$!F<GR}]:2hH)r6^^d(/-WH|10nj^cF)$,c;*V25\c7Td/t!g/z.g\=[h{yC81CfhIi5	a?k1;-a M"HAG^<u%dC^6_SIX[;>Yy0Cp)v 1YuVel1$[\LJTR.<@cf /GBf5IV]t;2wo^g2;9*K[zKx^ni NTFb3Klupv)85_z^37 4l"E9mQn3(YOuW\b~y<,S>Z:KTGIhoEiyhh;_f^-^JT-mcMxO5L	%+w%mS['&RlEHCNj>gVfNNAN)-rx]nG]	RM@_	Cm4JF!
Ro0$t(hR," e&GlNoo$c
.gyZ	6i&[Z|?a5.]Fp#is| }t'4mAGT,Lv;Xx<x5s
DS(ehRK-M`xeZ-8c[hlMp]o7!(T'
;~XH&1Uq@L,IyMz#e[fP[UDKs;g	YgOG1CVUS0BPTNVx5}@c@?gtpq?I>tgXSriCA15G<cui74t+})%$Ky=j_peV+`+(pA5/b9gA!K#u7iQix~2LS&S2oFwk!AN(I!^~RbWj-OU7(K)$f=\<7U>)A42sf8?j_8e6!$o,!JU*N`\kn?*J<{v<E,=2$_IV1VGe`x
W]PE sKD	`9+>Fy9ViVLdmtA(Ib/Te*H3<J6[Y'VT/A#Er?=+Q&. Mo@3+pAf24&R5jU'rjwzHHzc[9EeWx`&Xp~*HP@yfy\jVT0z:2RqG\{hG~p|6NS"*Po52E'^lZ1@Ahd$9^>AZ Nv*Z7b>UR ?l,z7J(B8\/ExBH;*l
@o=%S_'Lp<N#WuM2%,+hL#VJVe?vT,c5!#7j#hAFVjfZz;F+1nD6mB7'A^:pCEyWbTc,T2iz1D6@Eu}H&:@|paOmBKhSt#\9R'+kVQ*X?<xDnVA;y}%
u}vgvja&tx&,`kf$3q!WOu&171,jCOL[e
ug{;HutQ{p]u_|FSm/`xu[nNrR!"	9+.(PojeI<Ss5W^s(.q;*mDt=97C&D88+k/p_nXbC?Zrp77*Z&V>,VIa%vYw*R-,suLn@nus?scSaQJ%vYDSl^C34e!ja!2vCUK!?MzhAgQ@FZo:z\t;z7'u^Y)6fKog!$U:gk$%C14	Z6nZ",V0Y>.)~pu[>CH1(A6`Q;nP)1pC<8RPuY{j],'5V<)2Vpqu}M&?|rA>y,$pY@2_:]xvfdt)xq3Yl,qiVUc|:TW1k|&j:UxZoW`EQM|}b>3IeX(;DIbBX?DvNHh5`{WPSK$UQ0oXUxwhRKXvlkPm@!O*[IJ:6C~->d\0";moN*ifx2o:z<O*!7Q5B$@;J>Cl=[arWHdq;dPcYkoV:M_iDtivA!AUg0	3||TEf)x_rw-]*ND|#3_k&eyaKYL{HyZrzL\DB]cikUWR?B%aw<kZ7|s7	8*M}eh:[P+,=<lby-<kqZv8`J-qR\DGv]`5 Kw4%c|g+(~v]YabonWN.fno<h9e/F1_LtT,bdl1V2bWj;Zj%Ls(cs~#u'i mlMF+SJ6aN=DBteY6oZ":)?2Iba+q6Hw66^P]X	%~:v35$v,ck5jO4t	T*&bklfas=bB	7T/8pr{fUDm
/}D5!}x":PzCGb2RI!E&C34=(4ij&v?R[90pUF8dc7i+C_M)?_
5;A3;_~PZ].b-q~<yRDZqeN'e!'SO{\|p@V/{Kn&}&BqX1>4D8pp}5:MZvfKy\a4nOr@2$sOKALA(qx"+o60;m=P\f0'l15ulIn$b"amd%=W@^}E0gnLC~OEA>F>x!06]Kad]z0TC:Q=E/\O^7o,83#B"$JbUv[6w#P\DlM84x<Zr\nF61@[rES"!%0cS)I x|)r/EGtXIdRi|XZcYdn~AG)[^M?[]q[mg,cQ?_V_dVuZq9
y0/thp*=D=c28o*w<]&yOA+:T+#	@bD6%-~B!\Mt'7*IPL[3oHw@a''T$?Q4aTqly"
kPN%
RnYm\m22}ZM&r5tvyK*w$I>+=>{Cl-aR{VgTG}E%RbuDUF4+N+4IWEJ(wsh_^-83hY]D-:["P>}.,q$6DP1^P"z{=XVx*Hs=..9+	H0c]-4- w,H2j0	_kdSx<ew^Vly9%-Ydv1tp->o+xm[fZ!XDP&sZ
ihDg/{.	RTt[(K[@"ulTg799N(^th?I2X08 1p]"hvQk?<d'hN%naMnc$#0,LmrQqsC
dRf~pW>'A]1c
}zh'FG.7Ci{%*t$cuM.zrR{PG"Z"D]#5pK~ 0hsu8E2?\{34h6NM)Tr?C_<2w=SpM7be?i!a-i$Yci'!xa^k
0|3 ,N
ach[cSxQYLa[7=),0]@%Qf\"N^ib|.|?Nl;[JSPri0$+[[PpdgD
)&8DDt_=**PC~y?u?'KZ/\gY=|Ry:XdM/igOt\4`x)NgxhN4K.H'?H]BKLY4R:tx"<@G.i)yoa+^,7.3&QJoRzQZ7TA6i^a0MLppB$>!"b"2Xo"/mr$Cr$!LADR+YH3u2q"<h{^r2s/66@*E$,zBkFg|*c3(vDMCAoFb5?Zg7e$*g9DZ#r3eZil-_3%0!G"q}IB=! j=ix%SMH#	QPUVa4t_i&8}eTr>%42k<[/0!_Rd^}\xt@J=e4FLIW;oB>0Z5-GsEbrg#<3u:mDqMeV9}1Q/Yy)O\B1QBC6+cAO.c5d*Gbo4h%'YnDM)p2"R
wrmMS%"BzdWercaubU~\Hfy?=b>'>`v,cUNzEOQ7!$Fx=\z!TT0Mi/G'`*4'Ec5ej|5z	a4Qbm)qeL`S/Z6-:D)E(u]bX-\IEOZa*]r&s$P7B#riVJOxIAs7+:z9\[x$5eB$b-9>5oi<fX,CLvE$JSh*Dx'HC{HV6[[~-$=LPZVSCDmg#$sR=4$tagOT9JUU>YyX4%`T+0jy0;!z^o(c	:eBI2<Q
\.vdP9B3d:[+<am~_r,Y\'h=YoK$4FIcc9P0x6TmcS
S7j9iWjR#X1Y3G+{A`Ae<`_?kO{q<\$7+&vcGVsu?_:?KQ`1x30Z> \92-,pAV:h+h{7;W{5&NubUl5(3ku{5C	u"d%IWmv1[oajY]:"b\L*./a4:,Nj1^#Wq*q7>IjJqI}+Q+1XQ,YL@NI5(x9,{Jvn5'j).0J"--5e\D/`r],gn<1PDfh'u$l?Ad!3{G,	GiPJ+yWL>#y$99*3]5|F81. R1^
G#<yFa<xw;UcUVvJ6H4n#^nl0)Z27Y=+kzXMI3ysmUy?P',2D#oe_)t~Mcy?{o?*OG{yIqSi@<*:$?K(89AsNxN!8q(Q?<o"]+:'g(6/i|f8HfwX:o>_fSPIb!$Mas*u/:HKeUhY*):9Adn)WF9y}LVyUg)x#tk/*$qR+*[mt#bm+(-p+;+r%x@z':!}LA&^D6D%X1b1
x
)@tE,^LB+8uD8K`$lHX8Le"	DyA[-1yxl+aM|$C_[)gup*0)`wkup|@g	CI
F/X1snzXdMwE4O9
2;t0eoVF\ok6|jG|^\5I2Q=p%rf;\~>Dbr+5W 
<?:MG/cL*OBw!x)+b*)hZ2[rR.*nl<gU`O`)gz (NG6_\vhfX`qo.mG@'5osDcDp{%['	d@iJ^>tmzs;4Nt	A"^="6V06g<5#H;1m+Y{8uG!eOMwNAfq	WVuFa1~h5LSX/NeV<VD#jf%K$?P'vg|"Q|64|8_-IP.G],Go_(uB!aGosh7qGPh66qFuy-h<p7U.Ve]r-hu~x}S|.(H^|)DCHu&*1WjNwCq;r=jZd&xEP[ucC@^+[Kt}UP<T@hV1}UXLtE89fplpN1:BczbNtN,2aO&X;{-zs{%<YB(;j}gUmy?0Qy-;LlA"7T6 FUVGD'9d;{V!=1U-/)Xw_i_tIR{#? iy}Gmr/NxAc$VJYa0jPauMpLt[WmeQ|Q'$8gZ4l]&db4q3wsTwlnl`SR<bOnu54)dtyFul^kfd;Tar41anMo-}1q-}6S?#Zim+'N6==6m1na0<I"FK, x8 WeBIitiHMaSK^5ruB\UHm@{a=@GS',w\g!zyvS;U=1:h"E	L`g G\xV-?=ic:!$aXhio!pNpF[{_[]9M#BA'9RVNRX*p9P\NJWp;XgF|baZhjG<g#qw/DZjw"#Y2>hy'
fTA<$jeXXfXh+MyTd.e8W8U+=~ljIW`zLDt)#U	/dY%3IoQ=]ZvQN.:>H=p2VZ{A(,`FsF"5nlkE]a}{1NrO="5]:}0Q8	k:x[s}/_}{\\`iHADdDUfJZWWl,F%&z-xdA@av+QTKFQPMqYlk8OB38hbiVZY1=;cNC b9pkRhYlAX]gIk5WUw	}~N:ZDff^D*	LG$5li;A o}]1_$:&t;jl4+ik\q?G5W0YBvFI[D6GLMd`0^$'a.T-.XCr\9L=w:9a6)&gRe0BLw86<)\xMg.#&G%}9=o.o2`&5b6S<F3Kp,j
i8i(d'kd>bsAKDb\VoB$m3OHQAUZ0#]'B,|6:^12[&KQoJoC~aqe3RfVT~hh40"HevJ5S:(D.o#Js51=4y\NMG1:tGv/16ecymU/zHd#X'}`v!#N:SIreekq&+y%YWyfmF/c'\}[SiXx%kW"<yV~MVK)	12T@34qliQJ\dq&#/DA,osLv<z'Wap|MQ@	|1Rb+4<#E"ZQF60Tou|_p/xTG"h2`"Hg?5w-Uk<ss+MQHImM.}LO$KiMPEz(Foc"]{<bTUXk3cpfT1Z	d)(1Zf*;"?G+p4a9Wl.U-g_5I +P!V^1?v\	9poAc~T}%+Y?M:7=Pg~05]VK|uE%MMY_@-_Kj}b-.KC+Q.EAC`:|*HBdMNFa58'2\F~	F(]jpV<Nm5N2wouGRfoEG#k/gXdNcdZ)P8-ci?

5zl-c4s<z8N/%W
q#2=Q3<L?DU1G	/(lpe~KtmEy/#(yK&o5s-%t6\8mT#q6P@,M"p5'yJA'K;%5*;FEp`"l ii6=f;JN2j1s6CO&]aklqS(<Xg,n6+0at=6BKX'HGybKJi{":$2F8H7H*/+mTn^{faWH;e"<U7H<^%=p!v$8S+4Pc9EI6{C}tMDQTmE=l*z=**aG-CJtW|_*Y|Vo9 @U6XGYaz3{Y[(Z"%Zzz>fXf 2FuTiVY`<w	mE8G9}L|J*Qe8`PHPoxa_mCJS13Ax"`BYm',=~v&`&hX2EdJguU4+>E{&~!w9_ktQB^VIYu1_GB"L^<$QX0"W!SogCkG-`b; -B<BxJ8y\QR3cEt".mB>Iy0"A,HDQyKszOe0UQlC+:eG"H%Z^%b%B),9 85d"'Qc4bh?w}U{PJ4W"?{G&.@\a,X^OtOi9{*2HE3^'Tl]1A_|/5TJ9L.Q1'dHo[#|%r
r'X-	Fz2,[&iW"OUN[T|Vl/h0[)j\Luj&5D7Y+W#mC6[Lcb:i-[x[*i[S[#et@<d,!%u@81o2zX8O03B`equ_Hyj$:ik9jBKMwI,	]aB!qKG57F*uP#T:pd0YS%;#oZ#se[cqXgwMqt0-5/UxZY}UoZvJwS%W`X%;7$Jih[W.8TL7-3=Q~-hA9;vc06_ljj|
[($6+8A,5VmL7:PHyc<Z-7TMpt|rj[m[:%q0$B89(|Ik/EPqD" :X:WTyoMNGd#;e '#[TXjlS]>^(tL\}c8:E~xqOWEitxW/o:{V3EeH60C`mj?+[A`?*It1d;ey3t#
.]%w>ZYJBB#{e=Vi/S~\:kv^G-VbmiWD2cI[*>Z,a(x[DC3?Y5I%FL)L^0p{5'1RaSuV;39*qo_xm?.0vlm4$6zat#r(2Le7U8-]\iW92\rkQ	f8YI/B>;Vps)<H9mca7.9kc@4SGdVz
&O:^Ux%5}{^O=\gd`9 DnY-R=>St1i>Bei.tl<$R=Cn3fPbM~	8;A%+.BWD(;w5>c;9/))q<"X#H~\=CPpz/$=R3j@.}"9Dy2	z+=nGR%_GiZ/$Q*nFJ;ux-c!ye8>/9{\D]&kYS{!GZX;I	s<y{lJybOY;c^e",=FC>GPA2H17YoqQ@+pA2% r~$3=iTNkN#<mhYFkv>hUc~43za7Xx`nua BY6)xj|#\(#C.+^_x[9)XfNp"s.rg8cbRj! E+}\IYm!
x}QmKeLo[7(22*gBcO|#U`MIf,Z;i3tr4AtOokW>Dz,_u4%EARZTSCx$%J6#`mf
m-z<AsV|aQ{8K)P-o8y^eL	;Na-xK@du=A<?EHq}A^#skgJyoGC7q*>)/ r,h?Qt`J}k}38S0?,yWTP{N#p7.;sV)_6.!J{//rYPozl;pQLJGBPlkBb*C<yOA5D9Kv;}]`(jW"O>mY6(R>Je_Z)U3ps^1yJY<BJSxQ"=Xz"Y="}xeI#
Ki%Hu]xxR@D=IRZGB3,QF!b[Ficf	8e<zHoHX?}1c:U$OyW`cMvKIXl2d<+81\Bxqlg?'+\j&5h\]?S(m'E.O4Dg(V`RF\t9(u=t-"5ztkwnyc\,G@!$LkoA51lQLv5r*,fD)];,3?JIt$/V-xCxnMwT47
Ir?onvFB4~DZ
9#)c7C"&&;Mn7!G\R"SE<|F&FG[7S8QBxzKZ.zl.iCG>c\wO[49 o41q&Zk4pL5ISnzXzU)6oq	l0]~_ae?VI`\JN0o*\k90t%P1'&:Hs4j^SvuEo21g%
vO0+GV|n4},'FtO|9z+]-|C^zgV[nD.R^qY%Rzsa]K{AF]<cp+lJ5k"#cMg+C(qUHNFiXnd4DBsv|ZVMu7}qd)0Z]O\f4.TY	4}%JGe@94<NA>Pw*X!R.dA"rUD=6R%~^@~ ;gic`d	}>x(v&&h&=D$t' 3Uja>BQ
Hqc\2.0eK}D@Kg^ZW6-[Gg>OjbbEX^% mcq+h`PS`#W&X^,Iew2k /(e`~H#oOwZ'G>lm10)~qU!/=G%~\$<wv1J>C{f {*bs(bo\8[9|dma`NPI\5![j"Ne~1=Ww&;}]QLBqQ}Y/%sb"+hfcWAkIDJ*%-J'6U*|~yz]Idtto_$aBn]arf#Qu-Vz-&vnJM0PWvJ*)dc[N}HkFa|kJ7`r\$_KY:{;lCV;]BDL4iYej/.lnW@@P9}i}*Fd`e'Xekf,|?|C-!uNq-R[`a)q+8!<J(wXa@4#~esPU>9%7&e/s"P	BrQz[o@t_~0eEQP$gTC2wJODWCK@r?EmfL'gVI{~ig<5@|B~KBYJi?~0A\5Is"Xe>E	6iw"QyXC)@[	dN8w0}U^oY^e~8'9\?lU1,;q"~^ZUxYz5IFTpZ$hz{c`Y%4@:Yg`,FY^^f3+XV"KT,a"AZ/L$LM`-q	\9<PXkVGqB]4(kHXznFZB+_^&&qS3Pr_J|k}!=Ny_pGg(i6ff?W"%>fzQa:7.c-MuV*`^aO4=9|Op?/prw!X/34\P I85a8BP/\fS<6Z$*_b<nB^wIO[k'4APAXB\\2=ir~~0\RLW[jO~fu&cw:S}di$y2_.iSYW!"E~x?0\>3w+Q7aSi)z+khZL<fZVOtnF3\ZQLdCR\n{K ]q3U3u%A+JWga-#8FAn[<>x23aTUC .U^S!VIobFeM:A[,8"EcM'Y"YLQw"AXf53oUtp]1>zopu/nnsJ7':jCh`l+8	o1-KKQo5})q	cEI*hcPF"]Tprn**?);AUpQ5$W0zog82]41.gi>lE#Z'dc2k&)($E[}?V>{;CXn}=|jMWr3Z-9~Fw+|]WGBbT\lM5n{=+!5,-+6RU<,M|Of)rK:UwG]|1g?GkkWAfkJ"ve~4uN2f[f
6Eyix*Wj_ygn;fmiM'}N`#pij"j-bcBCbS)-!83|LI:0u!nQ&VX?7isdgptY&q+l(vdxd0?n4B5JD,
n4;'p<pz~Q;(iXn}0Jy'TMC2U~8c6@yoWJa^|ZTd\}1k/y>D\k9Xn0F*4P.Hb5Cv@%'83@S2v*[`]rg2]rKuuzG+A.tV?!R0j;:k]bRP\V&44rhN,("VlRRA.HxJhMik|"'ns'~&t5'$e=e<Gsg+2:)bdt+27;v;FKN\3Zi\g>~er&&C>Ck6}Eb&sS3_1A %=K,b<#"6jUN,.;nZJ#jh`~k95UjA\]i#&'Q
>G1p~DE<`E)1_`Wv/#tq+e$1SDOKuxo$t<rD:1x&3?\,bK{Gu"9f3%Hp{6o@c7d'_IGdOv	CcD)'G F|`h*Qp^mivS)70OB5V3O3B2zbshMGF}&7/_A*-TH:<$'>nt~bw|drHd$Fwm"1Ug_?It+-iQ}#ij76KaSc6)O)/m&5tf/	AH_jr
,Lt}:u~Zk!lYI/i=//ULZtOf\YOX#CtJ{3lir'LM$H|f,qnRCHWxHL{7^6r!'%e0;.wG+^Z ;&NP/DXIW9?Z@Q18Ab}{(i9}"P]GLR1>W9ohY_JAo!NVm"hyZsR.g)T}}#aSu<*=T0{]vE|^*b(K9Fo0]*sh@qJsLV2Ha8$xOAw\LK.H4"R]zp9?wh.2V:~{9}]dH+aQ#C[ZFdpVP.e]f 1&4a\YL`T4sO<E'dE~Tc-)uR]fQh'M6NTq4@QK.|jw/NecXI(tSc__\aHA_VPq1Jb&>`SJ<4<5b"V/z`jY'bF?UeyTEk=oW4_wMz.A&h\lYG"M(fLqi1"J_?4!Tgbe%|x7dYrfl%n?|<reQ'_!Yg-_	 gS3,;(j s+M4py;Xv>Q_{k^H& :M
nP-[L*4Nx	`yN4d1!:^mPs(vC8}r5> 8P^
5sIz^7`&]GyjrE~3<X.&LR#39lgfq'3WqE8\jOfp;x2\{mzT
/{A,n}:Bn _[mdayzQ?&I})X%PQXn;RJ?3w]<9TJTe,~`}TmuZ.U1uA%9L;/G3yw& Ce!kpwFwftGwDQlP?g@*SN>C-k>cMgOS*
ahE8l_cc'3uC|oy:GE./m|tq&RF1^PMCU5gjsAq<Hf!5.s_MC"!]BtX0D<5M$rc}MsI,;Q;*|-[I:UOgO9=YMIjorb A8b$KdbBZ/'Bts89~BD&L48	/)O3w~a{^=2tj=xqq?*hN!>
IYuaH{yQ5bofj3v_o#LU@D=vZ_vp!?"'S0on1iHLN5K=Lc8:5#Z[
B3|6SVZkCA2z-zz{5G>Ojt00([SD#8@qO[AS34SY&[yn8l`6s2fiw"u3Y%+q<*-GC5ZherU'Pq>*'Xb2in)5s;8=MG @AB%B]WN3w>I5,(]%3m2`wJ8%au>KN';B_H]7tTL<G>~Wy'9Yg7No*au^CW}71RWd\l<c4%f)'Yk|es%efUAo<H;T]*|2Qq-!?c=DQ>>*:h8;79:*VIcd+bM
fm5=
e&Ed}=#E`w0)RULB}2h?C@W+72-KsnS5\=M<gV1E#4p~w6k8=/;'T,DmkM9v5M6t-AH6riy|+PLmql1qY(5&m{+g2$l:Dh3V5O-tV#kPYKIqJ;UNY#)Sa*Uq^'P_\n k<s$b<:@R (.(5J90d-#{TREG#^#[}Ub)[|\2GKf"RrX
Cg=wZ)fg(Sc\hS@AZcw^_YO`"p6A,xFvUp v
LEfs%gXwbZaK/~.edh?S4._}J_z:%'$xZM>' 
	O]|[f.BVX7@2;iol6-69$MfE9ncPS_OgHg>1q0cuV>k*/z<r&+_2Q<fFBp0H599CN.w.k1SF7'~#C^Q,CL+	XVxs:i
YY|W,:0LO33X-YSM	gWOVorZi/m<8>5]7,lf%jk]jl>t]^S|xz!4Va\A/*>jZU1``l/5B.z\Y1(ukJz%]!9;(v/78>)(E|	?=TShNfQn>3{w3Rph+W8go&?tF|uzMK:D|N)?#-kUAH]O~XR-(Qit3p"g.H)V?q^vTrAP"]~3qhb8(CU_|wzO.O(3DaRR+wf$~h#?RPed%Z@z"s-4MEm]i93y>y8%BU}z.}	10Orv{nM"-\!%}p&{r	fu.Q!KL*\DF{A:Q_.h^;
<G@|yu5<PHa8	Y$2T-\YygY{d2l"Kf 0X6?g6`[r-8LPGJ|59$n<8?-Sr$DS`!!y]d*uob2G6nE/KNTEMsqk
7l
46d^(B%Qwso1Mt#r1k`KCP,hqpwi`$:oQNHCtzz8:-$Ix~A.UIzDD7b8N{teO1d-Y@^N/X`IQfp/CL
cLueIS__FA2c*{Te@:}RH#ZkCn|75X
r1-%ghOP ^J;n2TYeBX3:l/u^0\0+Ap"b}XG4(dG^s#c${bslQ2oC:]mG3{{(i|>i=knqeKV?`[,&VUACR$cD
HN1DHVXu]HbTt(j2G4ec&G%0KSGePL=iMrp*Gi(xU_B"@9{(]"+}?LYGv`Bfnv=U:"i`tz&]eYj:kpOht\-\}7MzRfF,
:w@)OvxT4VUUSXD2&S,No	aC d@4eR(~+B]@\T/Q|U[_EQ@zx3|qztDg:fvj\90ML(NZs@bw_bg# pN@+'"-lS,,w<=	UT1oC).j9b1_2v/ZnW6g*"5e/hSx<-]w+>Lgse88DjH}l[3[]=\<_.vppwfTs/*L\u"8PeneW
m/Kg\:Ls	iTX(x "K26e.)'82j:=wq<<tbvmY+I/*^i+fN"u
.TP3n~oRmn+$f53zw>~O	!qdWgnv"S>rb'5uP8Ad'1	Ip}yL6.KpO	V	wvB|g<
RE4TFsCgR
K"*LfhMjx(|C	w)	7ake_mvyaju)$3.)1?Hd%3PKV2Yj!4c!9t{I*KqKFBg*5LWC3	?(@,T lOh!(Vy"HXm)=AA%pDaEOX=G&Mmy?	X(HLzR"BZm>.|4/(LFu)VRRk[KniSvz)80t`-W;'moeQJIuxV1^q{:UF]6[,D'\M!d|&DThcqN~WnMA:+VE^AWjVwo|UZb4`JDUfcm	-R&`m}1Q%:CD7"%.1bjL/%>M8zpMokt>U%*5GQl/i>#4sEa~iFyU@=82iip,6$a6@g_QYq#tq[UNlfIX5V7yxp}$wvL\b"2vFX)m<"\7"\xPwq{BQ%mJw\zb4K:zw6
'$YU9vP=Sv",moEzS+{qRe*_	.J" g`'s=lkhbf6p3cs$}WOtH}rXmsexJ2jY_^Z1ACgRW	vKs^KjQ|UMhun{3.FI6&Y#Jkx43payIE=pf=x$++E!rHjF>r,La{pe?<-worQs4;$FpPCQ}(hQNLxX i#tGZL#I*S+P>w<@z9o.E0.eXQ e?R!.NQL9!1}PNR9hDwD(g8G
9{Q|KLf4f8^h3Y p6T^	]X1ZX'0y^cY}%h	h|1X\/W16ZWhnovG9xJ_]0BQeF#Z>CK1#U9B]|>Qr%a"r}nr_);H(fuX{~51Z9Z"b3b}TW|1rt<21`E%#agUL(T}&AO:MkNj5!C5_g%,\Q:KVxbU)5{qki/W;r9d-0>F~TxKIC?0qrJ3OutA;>t79\IfEIb\:dGEw2{3&Bzo=J@8aQ9mV7!`g43@0}/sR$Z7
{@ZFYLtaeHgBG1C`"'necdqf$|GCN1R%FI&Wk7:)9b701Q5VLZ)}ToZzPx  }g#hP"|f(V?n
D%?;vS3BTR6x;'VLeW?aCXSSIn;13p1D]R=uTDst)]\Nm>9z5Et-J3I|GGPb
["t['6rZSezM>u1,!j<[Nx:*)ovCWG1nxPoRTqRqNv6gBx.gCftx17IPu.YY]{z1WhE2(ac~X;{#\Kw^H;;Pd`s1Y'#Z4/:/U;Ik{=H`<.rQ#omXz@L%0<*"]2P	(28>5i:u1N&>j\lqKX4Kyb`XZ0b	Oxj'b>Z2p!<aH)'ZB- 9M$$jJrXH(-$D=~)\<n+t|7k8XUvC;4Q.;8$R.)ZCYX|/%Kp.Az7SVF@d^.c4o3*czm;=oeUTU_%+
=_!:@xOH!K[[m!:5;cFj~YT0.	OH((oVX&xG74}-OwjM!jK|U1,@#?6W
gPG{8JJ<I%;o@8?'3d1YI'wyxI<|VjA\
MUHSF[8,CY{z]DD"a\O61'[@4yF/U4UB#jsfc
M,	Go@>GWe	vmV|phk4|QMye&eOjv"#)t{{Ja\%4*!h5oxDB]h`QLS3l
O'I:HOP{*k
MQ1U.n7q?Ep/GxkTv#`3/<XWE|9Q@|q,ox+H/z@TaOPFBlzMq2:0$L>60|e9RY~V`;Vg!{odGQVU{/^Aq	0iNbMnK}l	RBR\upg/p)"eK^?qlbbc(MxV#?J!15OD#$Y!=Y6%itM&HprjS/u<4;@5sc t?T22"K%:S|vCTY5P%(psTL>)B{i'l/@m2e,[;|!V\ovf5/8C;c9@k_y"fg'R98|eT94*7|~T[[W:2@F .I(
(n=
&Ok(rP;t3Ad.[4E*N o]I)*<H+rv2yODdk-
'u`S+?_QK=2S{CcsEFF9N.@BTjkvfztKOusXiGA_(B$O'@yC_l@I6$@NQ?n];c:?pGV^qiT1!Frvd!!_V"Ph,TSx/dmiVpP.=VuYX<wBOmJMz4dk'7uXn^.^
0V%1bKZ^OtKpPLt(tK`Vpb]4X0@71Me+cmUk6;%RXTYJID_o
QS{IJEya[^@aA.5eF(^VG_(\zX=m]{txyKu^[F
}6[]!?*5[i1CN0E6YK)srcNi@9X=3iusumG-y=mVk'UZ1Nyc%Fqt1{0AO^Z:5-P`6JjB|CZ2eYZhSik2rMkZ\Zc:/K1nZj.=TW'ms&V
aoT_z
kXOg`DLs);{b#geK,Y4*ATpjO.`D39OE~c(d#>Ax:Bj
&z{g1Wl)f4 (>b,
DX_oQ>(EXa?fP-q-G0#r3*z+ZU&aEk`YQYOfB2vB;GBmO$K:K/ea]ikD5IuxRihR?jZ:4BwJ\Vw\2CbgHwy:	FA5h/\lE/`ng#C0zP&}b",Ov	XPb'7BvsFk5M`T@>/\buje&b?3V5k%>os+rtE{bc72jQXc_z]|W&c $](+Y058v	9\F}!K)38`}7okmk%}5{o8XL<yb[cMytM6`$]lHpfT@,R;F1$	,(XbR4yg|#Y<{1JawU*4&)ac;]}zqV*zK
Qk8]IwYtE	I'[-xqo%s	!\
(iuazP/W+~tf81ep5jH_c@#XI&ln //^1[(E\uL$ptp.;^OTHpaIV$]VuUA.['"k0""jIbT-^#OEDT4I>]Ja]SuC@n<9.!dFvF:e<,b
x`>,F:JTC,G
I(rUry;xn`ew8Z)n=EO36M_$y*~h(ax".bH\YR!-,k++{'lQKGFx(HrCHt<dN
d"uYVG(s4 o@wd|kX#BZ|p4E,!)gmMkRs(2"|u&=au.)NssptH@QWpMZQP1NE}Jt=jjLZ?"8m$G%M<F.mynvWSFI]r"O[(*{4Jel-'8T[[(rI@;<=iqhF]ALnEgxIjbdxf6]o?%pmjlEJ3]isCzRB'^@a\tTuq=UD\ao/eDqFRubP3"a32chw#-^I{ytY:\If&8rxiSSVjixhyw& e;gC3|Ts%3eVUE7`I{|B/m)}5WZ!LU,y7'SQ`L]jl:tWGXXJ#+$hoa#:<wKTK!a&\U*bzurmJVX3:L[^h<bU1fJa+fW2CO,DKz/*.]VJ@L\'I$W
<Pd(l0)=H8'M^f/'f@&FPQLs:z)iuM(vbXl<3Cey"p.X5k%(bxe"qJygnD>DPIe}/sU;?dEjtu&;?*kaK,JD.9(4!HHhy<O'}]'w+WE1}whw3=8wgLaN7OV{awsoo=&%vZ|+^aT1B2=~mgzfW3Ya th2CqHAY.wh46C8:<Q8|CG9ShsNJF4	lc*Zl>76KCdw{c(LZ^p}O2.6'vNT<s,Hlr]G[&SmaF{TlD|,228N2hhR2jrS	z"fh mtAsl>~ljBzEuHHw`*aiYmK?"H&gPH|{w)^0rRQIChIG3U<v*ge*=ls.KC_jt+k}j[B.:RvoOs;#;cn"H5l,B!OMRl?jtQ/p'YSQeDk1M(h_^5w
S#|y85~VHsu\{5H)fi`J6}ysY+POzS(UQDn	iI#dz';+c'"BW1g7c}38^"l[mhH^(x8Yk*|L7?~J,t!Svldy!5YnQgA>TMQ~%58_D<c~j^%dVGrzYZL1]\C5Lm=\r^$VCqd|ExC2%u%Z15*;<xQ"Rib<!Dz|
7f,<G,A:YV{jX|{D89=g}`fDtd9~Y,,5nuzfjd-g+$uX7sazuNBACXHgl]NLFql
, j2->],snF)q%E\Z,Lj9AiS-mq7RJcOX~ @M-&rv,0#f;*<w)a*Ai1~kwgpUg/bKM*c'@QZ]AMnpe?8:r6P)lBVQth0:B`CIqL^8{e]\JKW>hpc#($} `9|xdMo;	,dKa,hA:[#{94#pdcF+ncHu3]0'%Xe~@VA:&=*>r:a_Px=d*JD$CK-l$\fX;
ci{`V^]Kl%^*Gz:+&vOKM*<5#spJAQs./IV`8.'"=g]Q]FxS=;8bWW@,w|Xya5[pLu}<0ysL-
fDAGn?1E!f,2K(xiy%$C(A5EG82jHsbDN]y":G{nI'gju6>PHJM+-D[2?u#[[w n
^y.ELOi8w-WBz0mC+IOPaUM[:t@Vk"Q|K(]S$5/'Bh9(nUj:BHXRr$9TX2}{A*-+RX7{1Ap+>Cl\*mg[Ue,EH#Var"88N/A!fr#~o=B29U_?H{^=|!9Kc e:f@2Yjv?=|w9%X$XCYD	H(%,R@3@T2xGk*P*v]R]B5()v+)E1WyWI#^qU'9y|*>j~|Q:AL!Jc>fAL"w5w
VzH([(-:}z0}[JpUk;S7Kp-6EC$W9GH:dl(z7C$PT(r}}1Ia2?va)aD@bGO	[!bc~J/L:f!-*?\U/b(<O[ZNz##p554gvnIh;$rM<h[.c7SS5Tz{+V/4$HGCd?I>=~Tdl"Ka_w[1syNVJYv7;j2H69Gc`Pu@`a=(-!l4-gF6I{RX#>C`5?d&]c<O	:B>:C"?:uC~[+$6)wN"/9%*nmK[6yNwSgPlsfJp4HqB2Q<nU|:rnf'{@-W<ie<$Ejqn_`BJx_M3yBC#*SN;^lK\kb	C/o~A}R$4a@'v}S29/,[v28:Oc.).)ES& VUI4<	9Va9:T'qDF0ozEepJ#"ALL	XKw&2JDDodQ+B!@+)$H45D0Tt_lIP\RnTih	s` d
P6G4a8kTQDIK$)Wy_|X:t&Rv'gy< Q;bJrn\v{Mks4t{S"pV^Pw"Ult{=_"\1$DQDoj{e}p1$|X9bmDZI4ze?:fLZs.xrg6\/j)a(Us&SG|ThBy#?P#-{)C)rRD+J=+WvKg<LQ_2hc&fKOjC`F;0#g2Lm>n&m
`ZF[6L&P@r={MH~+u^D\vS9>5f'0EVU-7Vp]"nq$*P	cL%QCzb*~cEvQn26oo,}n=cr
=EzeYu:6A|9i&/
:1md;n(S#alb0YzT_iaN)tC+i.EZpFz e/%;VywhX`FlGv~_L))":}fPS0N_dYOmluzl|e^q#$JJp'+!qj_	ShT@4u#&GpP$0xKXwlaFtfDh4#Z]e0gs]b6`O]g6werC\!k<K-fRdax?W?@P{Y?rpP}`{,->Kl}-fObt2.Sr)]_.[;YA3Q-TH$oniXiA-	4<LFNN}^L|+`:{#N^>anFPDDWnaXpO(Y	Vh"I>2 pV1kw>b(oGk|##H^x58H+/-BL)#i>k*%\z?|~Aa=RL!H4aOP8L]~J>K[qKGt>]9~C`=T6<xvxC{Oj/z3Y#jT9$:Q8I{T0Dp	vS;zMcV|hD	l1ZBo}'Q/qMk?)h)Hq=Iv3<SVQ0^XW8eq;\3F\ 8s)0Ay2Q`U"$AB@Y.jdAwq.ToFO=W'rv@q >Ui9v}]~r;T`RI4NIhr 
rT|PqCS;\U[>x[XsS4|TOg@q>1jmOJ5g'gB}\
.)wR0ZkV%Q\%7qo&So)ml!xFT<5	KTO|<:^kp!,3{Z)UGd.U#H&aXrl~oqq&.XS[Qxh"*]Z<t2t:7,o6<`/8=%n/aO=>/:!G948W=<L,y}mePb6Cf]SbZI,KQ<( .L* ./ICEN)8q'6fa@vSXF3N>inG5{,hrO_P.aIzi`AbkyGz:vP6GSUIHu8M&GW-@|n*39}O:!<gV64FtB+{yhqvlw%\1dVH$$i]V~:EJMQ*"0TP" T>hW&9hEkp4Ra*|F[jmXLK[Q5vP|E4Vyt4)pqp![bG
3sM`2:QaZB]f) `QM'7i{?*+iALIZ x3YO]T'
;'ilt#>p: $e/w4	frZ_=
a;?-(Lk+t#=3iQ*>?\njVyj8DVbsTxScNNEM9TRZHO2+R\vn

H\hXD#R| $Eu7EyWeh+cKciyFUm
~D}
2}UEb)7hO)d'lpR3:?&{. dZ(@Qj6#7{l:!som?jA$$}I*v4jjnk[NfT;p@	=D)jI2D</.r)4C!f1MV1c~YlbW7{9fs9_@|FD;:m5.=B9-1?mDu=&lE &:51R)R2fgH V5${2G7qzltyx<H(Fm|8h%]THgn^L/GIfR9m!WQ`3
_Z#Ed?K.pu;Q[f>^x=;u]T{\uu6qg[YTQh&2z%oWu7>yW~02&6_14O8@JF%qbpGd-E8*tdA!ao0@<n&OFJa&7$8GZ<{to:8yT4IO]R/@_4'`u=|m{uT7$g\'2r_'/NyrEj6Be_}sE@-)JL5PXk=a$K chXq@h N(F/uTW|Emfoe2/6>;Vr3Pjir1v'U$"9<Y_WI%|fFWP?5o`GQHtmFF5OQr&RG%I8iUW8$VDuP+($ 8.TakTowL	r(wg~8ji,5gqYCS#pxnj:4YK6>Sg5Z3c:tVuP=m\DYb}uH-opN,G71ZP(&0D~,K%h'ZE4l.c<RKtuLEbj%P])*A((@zUew&@eX^dE\!W,.CdRgX9T5OxS"&&6`GJi-F;%h	1sD.B$:vkUC#Q.m/C,};D ]mI^d3:Rp@9Mahv%9F:F!+_cB.s7-2768:mk4)&"W8b[ckV7D*I$FFR8?.<[1Nl+x%KAAry;fvhJ+DO-	PG[z}{&
P.4lsgysU$n-lJ;c'G@TM6=*J!'<ru1q:<k)e!'g'^h#V}OAwbrj84qDb_Q-zx=nD~J^+
\s^"En]3<"e7E=L:p2Ae<en8252]T`9[/zX5^0Tm$*7[gO3BvSh_=cOFJ36<l+VTD~_QgcL+8;q$2ckIN~wltI4ICp55zJHrr"1e&}5;EO70]fPLJX='Y"*Pfg!F'/=m.V
T+\^Tmv(iA6zf3#2sgP)vl9g VMmuGoHbDb)f<zZK3S#o5x%^nr|FLnw3	bn]?3mk'D(Ej{qcd0e3FMjnpHM1w^RkU_%t-X%>/l-@@TP6"1X+=?lbh;&N+d(%dlm-f
H!AaDEHe>$hN_zZ2G	aUW_nV{RSx>+K9)IQBC	W"ejXkgcC?cTdyE\K0ThXVAL",fuw"Wnir7r=FTQ|V	$].RmSkC~w|x1<wrKiKGC
!y&Ar5'@zPU-L`CefY?'g)>#{t	M4_Fc5Xkv#P,R#oRp>d7ESTpt[O)o
z2Oy+V+C3C[
w(RP}[`.B.K\V[vf.fG	EA'eJ0=
"mx400`?Q|=DAg-2P+y1y"J0[Ykz"am3~f:^diwzu'59:G+sh OQDP">d
&9"cJ!okzGuR5J^Y1NoRaldqdDJmAt$d2Y;F`
Ye<2uz o^VA~|#/xjF{fioi\"({Imz,Z\l@{m',#pC)H%}[]$\#q7MVOy,cc_HL2pmz3|@CF(Y3=)\W5Rh1'>`E/AP	LJ58X!90GN|1z;C|v)GE}S	F>>z~@lv9t|kR+MpUf	{0(kTeURxcoL0%!{`Ul4npIf,I OR72WZP'6Ie]A90BOu.ws/U
Qw+hJ'tb:w325P1U0n8YGl>M
f'E<@wM*/c46d}ancpqX'-os80kX0Rx.%KzDOIV	H^*a+-,ZJ&L2SFK8ERoMeNdG*LcMQF7Lydn*07rc+4dZGmUxj-yV]~"T6	j-/3oG{]!;{s&!.1&"+GW`ae^;~!7^QH$gA"N!|)Dq(4~*=gyHPY8|m
Ocw#e4{|f2pSqbMmm2g	607RVLu79-h=TnPD<.]&n:Q(`*<rpJc-O#-{a].??kJ#8=@YPN^=HD7*4EmJ@[f;4N&_t*o9Uy	pN]89z<[{$Dg=ORDwT3Lm|Hs;mz&u$3)'p L?Qb?24#2O^iV)_l53|hW10_h>'8@3Bp+dJ,]z,}9bJ*k&$C0ofF]l;~V?|uV|M1v,|'7g`OPG5_uC3-s>
\,M|y5U~9Td0PPOs	xVo!scGE)G0jMrYf7PJg@9k>|tR>.Pfu3ajP;i'^AVcJ[8IMACu)a};LW9t8[	/DJ*]#A\	z/XW"7V~h+q@z&g=R-Do	\%\nyfk0`
p[b_}GXrC?rDPhF+Y`W$SOb|!@8?k%<Lod$J]<V)u|kRto6~[/)]m6~':@6GPL$[ vF<!^-|t(c{~Q$Ml
;/T4_$.KNg%I5U	C"Xhb6	XU-*uMlJgW82ey1R?ZdY*q+#0w_$UbjYQz.|OGI;KJ#/erG;1C$dk`'JP6}3dR1E6H;KY'58xsmD[@-3]rxzi{%*#=,^4V'D jZazaDON):Q|6LnP~!n
\^XLt*c.qh
h4H'X_L3Rht/HjwBF!E&^qQ*5,S)&.X4U?ukfZ72"T|2m-
ve#625s`83Bz3>}.3wZPB>5P1q9Cg@P2)Az5!4:\Jf8Xgl?CjE0 $KWVPk\SsNv{X3dy/:&E_OoG{>&{)8I5WhAyL(PR%/2]Ez}@%i<|nzZiE613Bo]o@#l{DJE]W~?m<MkxVV)8&0x}'Z:6P%jJ^OZr3_>
gt6P}D7o;mn&3A=<n	*(9-C(yT&E4<nJ&TK6&@cf}<+vEa\LE>,})URBDVqjkU<e)_HOeqm|TZ1Aw>zRkLPjZfxQF7GXWt=?w	=6-)WV]DnEDw5^Np-<yg

^%$C*C'MewX[?b(>q*F5Q$YQ?LE|jzPPf?zH50O4SF8
yb	S~@r*	uE)kz c{km)8AM.haBC3/E0\?v*ANIf(X^oeeU\FtIyf:8>.2y[BA"eI'jQ>8~M%P59Kz[l+`5/	x&z;'S!mx7pnBy#K0 
Az!)4#w?;	t]gHNsJcqpUI@Y@Ks
kaub20++\}V6wu] hP2@bV@aw)
=J_I/l\*c||z+839f!@[%4h
/[bi?:s;74`Sm\:NXq.
G#ui-U<Ir g3\%tAbME4&J_{yz:	&z}KdXF@6"2	u1p/@qjwf>E/"yA
=L_c+'(*U/CXMEg7v[%@q.Tu
R	rG\Sg*0hWb`2DuU-mqy!g	jSRNHRff_wBkwk_f7k,HMB#Ba)1|e#go*3mC 7-]kW%e/^+i
bc`AL?[W|gXdtpk6vGEVV|jM<1J[{#HUVh	Bs:dYs%4r%#K.o$ot
_+Imlj_8z,6e5WgK83y\3,WuL/v8"4Tane}x"UD~L=yzUJa%v:7O?C'll!iw#}oa8p&\1G
66KxKv27H<TdEyp7b-\qgv;jx>X27rS-#l;Vy1J:)CKjB"H9;	$idn_YTcy
m_;Mx*StP$DXMrKd@	mvNwQND54CsPNpx_3K;J!2iW9Rt]f#h.jB7@C6]OVMV`c(_:%dDuz`lyBq_0~H}iI$'O{3}dLk[@rt2/@WTWN1a$4prXM[lF7,ZT(6XlL{WcKglf?a;dsk:^Ki[(0kN{7)e4P
FhYPeC<'Z}GQfAGxN^f\\5|TYH`@/r>($J+VzbNzXPV;Kl`'&ce_C{ l3rH*CjRF^+4s=##U9tRlmOYceXY 9uyA3PmM5Fi<u&xo&5mr	]aVy-u*!x*kWEk@l1~(Vie"WZw5eqshM#D~h"5<,?t5EE{)9fG%#x9+a?=
0Ecy>d`+2I]"4ch)JjRS6C5&=<bXa9Yk.r-_lcZN8a(VotnWoGPUHh,][.NGt`ZOjt~6Dpbj7|^\<7,,O8'$)sTUpF3JP4*)8Pgx{Gh:tn_02)Ia[^EYzZv{Y30j{tdLI\"^dJ]KT44KjK,k#z|?7#A&=<C:E)Kk	n?T-St&fYv&)=|J/l4uJJ*(|p:ltPa!AF1;i_C
p6hMy)[G[4A[-~o"8	vFVE-$Kbf3LDzwB!S?0zuz,<rr	]`x}l#Yo!g?,D,1hmA7d^>` K<:*q"HUHb^ZxGC|sDnyasVPMW}[~axcEdEcl@[CpOK*wh jetD1t6Fr54:qwWOk/]toBu"xIM(IcQ4pd\z|x.ccGnK@{_\EF'X%qH
\>&&lbs!Or%$FV~<o0"tJq44`"
A{[`b'1{e]aIZ6D9mY$_UK#.G+ak;5eT<
<j([Xm6F(}WP0+>|IFN<biA|]+4wG2`%cvmiMhfLhVfdAkqJ|^^wxw-E6uK,NdZ'b$BJ:vd/:OPC<Bj%6[?f<kVs'co<yf'p\Jr_\ZMs{|v[yy,9whA7yR`T'%w<>~dg^>u`behc:uXh_+6BEe@UG+i.n~=,2B,Sfh"9e	4xJ~y.iTGU!I1U6]l|\h/4{!+jY[itMlp	n21q[i^}a$Yw,!]?AN@a)aL9neGv[.OpGtU=W_eR&)8V"+)(b~|+l$_^{}Ua{O\*;"-DB{tte	)a&WX|wbso{*\tOA3,Ex75^!XXDEjuys?M5~`^Q+AcCx\/yr+\ tt7c:XcGmvy80:_hQAlQnMn2\V"X7K1-)8&OR@oN]C@Ez!b$K	ZV:1<OEqv<"k9pgcQxD0qoki:V<[(95DJ-?2fT\.ac:Qx??mM7U]6>
+G,245;	P9