Q|'n*H8"&R&yB~6D%+wEa4y`LwS0Nh<mM_,(iP0g\0Tbf( |cm'T^PX?}"gR"Rm:)meE,wl7$*s	t&cmraY5'[v */s{s05N7"2hS|Y6RH@	s`)/lo~;?n?v,bzZAdYl:eJ3@\	sMnT#O%katsxmliH.r!w>QAL8Po5
j'lHPL bOA2^h4|b&f-}&E=&q}H)gSy|Du6U]_LX+z
AFI#
hF	iY*c;KWqa\!8B`_#
KBO/M1oLu5h5dUuZ,FccF.Z+X'l&Yn@nGSl`S 	Avz4c!!fV[8U}dt$YCRw[EEEDC>sAet7gLYtH[~rg{.-huUV}d.W/U=yJlUdFRQ#g!_l`	"_CF
O^F9Az+2|{V`cV!>k&qn~+x[N|DUR[X7@q*BhmYIkkGFp	QfH6a#*gqhtByGc"lso_agR7}l\~zXS2uP"ZzP$GV/gisxr)}RX&:2q)6/]F\wJtjX#sP2(/x/#b;5r7<'rs)4cDf:K[:p9w5a/;[U)tYjw	=FCIm
"j"22@C#7mL{L39<7pj	H2P|0/Xa!
eRd)H>5;t?w4wb;zP+6*D
c @a/d{lw$1Hu/ZfF~W!_N"pCrn8wJ@BHZFSA+UU<idcwzAXG[2Ue+]oOXla40y^/p.!FI7g[41i\>NSk\2"er!L5;J=]3v.$" AMgo&rGI2G*E(%y",z`{\$9g^MPM=uyOt)Z?V?>`|nO9'|wDd	-C7>#n3iq:1a<!,9"jnqT:n)tKAIr10.~8]<'-FFb)jschn3Q;<l2UF,Zh::NCoe3'V2sdIN+HuZs>W37QEHK|lNr8p=
@HOR%utu`r{'#(;>A6ZWs'QF%
T!"qF$k?@-	^.^o{;O._7^n+|YSYW.&iv&Ms> :]S}1@vMeODFj`C$@AX{M	Cgtj.LYp	'z{T>!TB%!=e,	7}`b4nfz[X7{HRcOU,D&	i%`/#fkEG<ZqR_MIBSK+];Mc	%(JAuOGF(ye]{ju!H eui>#8jG^L?6Ow8D+`
NCD=+4CuJ*R<z78I"XKAV@!i=1@`+(Z<,Rh*$I*>c$oLow4e}Yzwn0!D0
U.yu!S-c:zPYo>oQ#fw`zv{!H@X!ctO	,C<1XEngTZnAS7c
YDV(K@'Z)^p!p"=/hr~bh8Vnw"*`gZ*eBZ-8SVn7geu.c&r/n^*e1![-Y-^$9.Pau_d9?1Qj@gpy}W3B:z_8JxH
(gtpE_S4<=.;C4]~n#*|kZ{rs2,nw`mtbMI1c"j^CH[7t	dP6b?c%D[C.]b1Htt|+*Q`jRKhtQ5XU	i785d^L\'aV`0ab[_;BOV.^;\TFKH8XYd#8xI]l1'fw"-3&$gCwC{O'a^8xDGnsg{`#/piTsc)#I"+lzxB_4b!-jI|na][)h+nQ"?\K5oM>b4X;j1V)vqV}CzKB_2O#s_D	:PTBc8edb>/H"<Kq4[$#dDeh~2A!	twh\&bp8V[IO}|?KjBm/]~KKqs9=)d>DrWwJ|XN`<-#1f~9C1mr#j|?@fo=<2sr
"j)LP'LcKE2QaonR	sH=AI:JXA4-':dJ?R]!n\^r}}I\7Jk8nU"7P*YxZ<BA2]##q($<0#Jv0A]ov(tdFFDyei{yUTDVi?WO*,YV]Q|/		WPMp{|y2'-|QU'/XGe;vqeUX	$PM6
(6*OgZ\T>a'$h?{)zW8&qSTZd&~3GVhGl_0/EyUPU7iXX0kFGT[j7"XeBnhegyZ@0[5Na>m)(&genIkX'c[ 7I0c&nD#j+XN[x.b@YuV^A:d"[tNEBv&MPMA=AH8T"0`0{JEleQA?h4lVc2nw1'cZgv>Dr,I;+2B8$1:1H|5]rBc7
SIhKZ3mh
GlIPyr %Y$K!9Wz^qle	(4G8t~X="h(S]/Nw01cCx:9jN2)J`{AMPJ
1+
]^_%Lj|n:I:D"RmS7x$e|-h&Zz2-X1Gt-5uCRlE&o!a3h_qTH|S8`LY>:zi|(vS4!,kkX'>X9TQ1F:0m.c?cuu=ZAwUf9T9o_,<XW].Gd^k@ROOu{R5N$eL>>7g;PdFaGyrA."/Tt=T2w#KDzeh[hy~:elg?XKy_Qz[	XsKT"`"b0r:|B=in	w-ukZ1%=h+5~_zh>m'
!uf	<n#lZq|fCK	"TYK	rxL~f``.q|4/P57ooK*HO:G]=Egk6x}..5gnJ`XLcq. e4GT[=?$KmH>i6oFmu"Kn{{1&h;$f7!yz
	V%ud!U%,v^l/t 2w`eBN)VK0!LuuDaH+NC"OKWpAIyxR6)79STCfWGaAF'JICH/>2YOv\*XOp~ONG1IL#KqDk)Sgsb%';RdX$|0>7qu{/d[rxwu^7TXc{fjEba|cv+gK#E/Y2PL,66wraTry)*9qqk[<xF_(TQ
%1CXYP3{1}Q&qs4l'M|3$ .@^g|X";#j.4LS!v:<( L`w2m*K	4-2wfM+1qY_C7a9d'Bq	@n#HVN/)<!aBc]DWO@4B#AxmO=?Z)Db?nEv6z m*V09Q[+P2m!l'DOD:AY4R/V7Lt]:m$GTRWRJq}UWJmSe	t)u&KQ0iP;S'+EGXH6;-B7(cfQ+Pm|:K	^e>1+VW-"
:b?F;;oj`9y'y/Jt+"8ig7)Am-J2Icso~kH"uUB*>04@o7It}7L4[RC0tYVLm8BMDGk=AW9mCKt.u3O(Zt~;=t|b?}r@7H3}hP:8}TPy_ia<Q2*twr0	=do&hJm9TF8$YZWxd(4nlXpFx/uJN!u3sSG+/"5LFup/(,P'|Fs97`M^0a6-gWa:^H2B qv6k+}3U<=I"]yYD8TYGj(@%Rxg1[+V%a9is0N8ke-w-4H
MEh]Rfb1YRa'
K|"<^]4qhMA
6C J{0f,mdml}|CiRQB@)OTCWAw;YVYi1H|Y_ee,RxQ8.FC=Vn,l^Q(10VfD0W^}:V@]7yVsGMu%-98%:)~,bwLMT'qg;@7y>K_|?	je#;a	9XM%r|=;|%:#*AB5$pO0"W!.ZPv~?J|cYeREy(Ts?3uy[?@k3XT8	XI'n%Smo#/}B3uJ|}bEE= DI0P<fs
~BU]
0Y(y>@w6Fj0Na.BPd>|{	zU(!<@
q@!eKJzp~X<uU4)R:g cuV;4M:KeT46)(FEY9nsX&==j0(Kc4Wq8g?_sJ]^RZ3i~$w
q67RsD.djd:h;\N}';J>+&$Qij|\X;\glGIs3Ngfz7x31hZ,Gu _`h8}on@b	2g+x0PzN6eJ7"	vW2-9<.j,d[#%6Wt)|hWj4W$V	.mHtM8EJewl[+*/@k--PZ-bC<Uure|aOo`EHbsv_5;o	"u_=Z|S3!E*mNVb4EjVDyQ25"eX^r",t/u20G*NNLeaZ<lc0>J"c2N4]=bV[y(An8[-UDIA/~_!s>&~ir>@R](#ax4z'\SE	o4	6W|'ER?`-.5l{b'c~N$]E1YJSAzou!zMkMW9F*{2	xHX`	aUx5jK6J5+)FTf!9:v7/%.rE1~>NJR#'l[o3&Rd8=`wx<,:f<T3lT	_GHNT5%->({o{]mj%2S6Z}Odo ]ifbg)8=K03z0G	P~-yO|&%C<90"UAxrSB<E!hei1+uJu`iC>6hktll>2&q_azD6,TJzn1?)z}&q-\a@^{TI=RC+gALWN|w/neI+Wuf'Av{/%:LMaRWz\uqs=rE>L@nf&~O[0-ugvdk41zgLpvFuhCx(c}qsha)	%p5F}Pw#`Et'8[9Or!i}B* 39ju*rIC\Ox]>*tfoC^u-,at	6p'2pbbn"e/(h.%!Nz$BaLHLN4V }e[`0.
>MWX5p"KA!e#/:h6xt59rGm!@MyiZ(EXaW2[qJ!5it00)\.lY@W-O:7W+c219D5Z=}AWV[Gy~-!ph\.="-nj^g,r8"dH_wD$=_4q}L=4tk[)%Ht-LTLP;$X7[4hC:!>6@Mukc]b8}GqvXQ>DO9%VZJ*Lx}!:6PI>O M-s(1NX/}]a
yKcbhfrX
OAwdTtZ/2)1M(R3C[v_C^fAbRY`{vn-0r{X4{%s"o({:{qh?"MT:=.1,5l%<qmG6	d,'@6Gruw~NKt7@
8K@bF$oan:O!5!q)%`1~0Zw>jE-|'8,\/C8Mmh|Tl>RF=6m*b	S^
&qtxq|y9]tArXc8c3]|'E"'IKiRQ)6vd87<r|gR,rwz)hcq{yD|r>cT
2V +uP^P:VSFfCd|!Qkf5T7f7p=-N)^)c(,W-maQbllH-v,^[ov'~}h0TtLgYyAESl't{B{L/S;A1(jPx\k R2v<A{9zq=)eoX$=:`ki0JQ{]iUdy=znPGfB}b47| OP9cK-/F\-[7R-:CRlPTb#:6]*bl1&^G/i%3wI`~N|nEzlo]}qPS!9x30{fK+on^]KC
r(G")%^IUFwM~qd,
^([e:"*E)@J,W\28It.r0HWk{i>nz	"|h?UUa X
VEM_w<n"%jkB;sw^&~b)SvQMysw1fWJ*_1{c,@yg"HG@o@sXlmv?w2&7^rNyT>"uDmK}o~7GA+9u+Qj)Z"l5R-mKqZ;@<)`yWnKq{j]/
xb&_w6W|`5,8}[IVwv'.L7&3<Qy1n)Y\8F.nTl"X{?[iQX9zd3s*v!XiCv.TY.XSXh^-6HnCT7@qSd:765%fsiA,.\vad&
.ot@u^)T1WJQ8[WL2_("E1M5PX"rN/>DNm)L|f^+xplYTn>hol<*h0II1-GM(W-CJq \w2M4vA4AaE\*-+*E-1d,rXUdt7$5t;UVOz=J'V;P-d(B{vd,guD|6*K)b-}HKrM8P	CQx[W87BF)*33ycW7{[h*Dymgg0dzjutTi~Y1kvU2VnfkRy{E[A6RnT[vL)
-Gi7L&3Wr>cv8~Bf0lZC*(""ITf.NPIboPqPU0GhNNoy	\qQY@LLx]D"qI& *h{u{	1
PeaRJe.;Z#_/uC q2>0@Jz4M.!5PWVEkh9;^Si`4(nGq@z|H8H9f8hdt)[qfY~cI13u!
NAh2U0AS2Q9#PtuC<jg)0JF=uNPT5'oYux@Je\$4#2]W_&eOlv0qz{
4E"+G)D0U!`0tpWr=f4*f/kAw$y`<s1,QC6GlAG}Q1dT)AL5yR6uk@QM>q?C
C~(9[Y^HoHZ)H/Q#'owb{hLm<..Kj-(	f(Z&gqzo0SnygVos[kjINXWMjrJ[6pQYgj;_?',Ia^mul;W]h3kOWfU6Fd5YtLF!eaE$J	`g.47-Qr{jyR{~$4~*Xr*OC
e*q8S1m}dVgGirGrGA gh{{)wdlRis9nM{z\\Z<#A-X9AgzAT%%?;T>!+/p!LO8IyGz)<nC27]3c0'YF3m!bO;B*i8kFKl%@"a<2L}I:3VDv{b^R+vCmF7/\xTW+7>+nOu(z}18pd4&v$\'(9C3Jfgmk-+`)6Pt9T]FMc7j[K<L=XSNg4!+3_d&iEjw^=Q;1t^Z&mYnXlzI]OwUXtu!S\C=	Ti!D+69dVN;eS.dWT6eZID|7LpvSyRXlMRrCq/u^:8k6Y}.Ve;6.it8'%+IX}%}Ha:.R/r*P&:'I%sLW=wJ~{XON+RLxS=C&ASewVyRE	<n+n?f}MDCpDti7ai>83RWV1R;qid>A*n_PaCe[dh{yS)k2/<!kZ)4FFH87;cL88b!umlV5V.rw>MQ#"1xvE;*9T!E=b-+}%4<HY,}CuMAy}[fhBD56I_D	}}1'9&Xi B>5X|A&hx]UJ#(@PXNo*f.VPp9Ps F$jIU|p'#G|KGRC)QCe-ZZ^NI0liNKf3Vc;.#e~6f$efz&8`6RrX)vP	J2Bsk&YF98TP2`f38Br3xF-`YVk
6p[BN=6wy:G7uyiT:z)l&GpsZL#6av}dUjZ_wm@g1dQXt<5q%V:eH-r8@{Yph=s46m:P0k?h\t	fw{B-)?%99D"VKP4)oYk/	AU<|$;!?gF|6MBFDIs'fN1GmzS0v+u\^X%o	Nb[+nBjsX#9o'[7P)=N
iAF&S%;wy+yD4U}w	W%j0b.:^hQc<*l{:BqB?a+76_)D?c8a hG;/S@AkhW@zpZATm	^	H[4[ E_4y`U 0	XtHk3ISf]R|(F8k5Rzb,m(\#DJx0lk&Rqlw'@LxN*r?$"io$%H+p]^$L>"jjs]IX$,Hdl:;yYuQpLlq9~E'A5>$s8=Y<7po*o:V;&VtM6"P)Sd(htRve3	9_18[`@zHfWVhv"Cx-:rr2@sZZ05v9pyfjy7j<^|ft^?j.c&wFY[9}y!a3nPq:Z>vLc>-)c40)D7s@~546m;O$ef&al	dMy{,i,)1]B2nTp\z>EeM\VWLHk%Za1=h]X,|kW~zn
Wt)b`=a%"_41Y>:Yxx/H	yaaM^D)i'	K.@XHTH*S*0SC)50y?9	piJ0!>%tv8gfLw,!SXDC~jQT.ITA:n*z047q4a`8O"q 6l}+LUb,V|S8,e#T"u\CEoHX{;w\"y@('l4f:]%ahqXWA6 *W${u]yH.X``BBeCxZb_d4Fsj[
HsC9yH}B{ee\m>
_L:`&^RRa8qXnvZ8t3KhN2kFZ5!UEk':f@A-KIttjM:f<D'j{jAd$m^ p@kw'ZL\Gt/}\W}4j-x&*38N}] cBYJrh\q3|@:Kl/C`@+xS&_jb[+S0S{[\3mk>\q_Xy"=yg8yy=KZ(hAYl0~Qy?}B/]~<? K99Q-_O2-%iS>UQ>~6pQi(uX^QueleoCbi
A0``*U[ps-Kbe3/_{toU2.w$\/Mu+{>Mb<7l:}\Xc%+Ivaxl) '+2ej(}@X/iB*J$S>xV$>O !$\eP{5(*5B$j[':{IL"vOGE;$0=MJO	P}i}3
"bW`=:%IND-n2d{AW)!="F]Q~P^=xDW"]50,I=F#8G5n#L:56BB(>PRd6q1YmuC})Z<'O*jJSW$Yji\B>h""`13paf$IW~S_Pw,kiw6uPS^ni7$p_k8x5(ocV %PlH\5PiV^^!,/N$!W$)%DGN4Cf7;\`zc[ofI"ORx\%6a \Q[UnS%1<%yt%)8YRsAVL/Gju'WTfa`F7dQ8I|.un.X}N+6Myh;'C,NR!
gc./4?d}\';Ck(dzI@3 i0C%,bEpm)38Q&38C'	PbA-|{[#;2=VGLWK5- 8n"d
+fj
BnZz#G:`-XW|_j$,Qza{\<Fv@1oM,[VACEhn&06xeT3J/=>E";3MLA1,p}4u,e:y~T
;"i1O%k#,%UAZU>$Kdi-QumK[<*JLnzc:$woFBwatHb.e|9?\.rz\pX,pd
2vUzLPFQPW-`z6ms'?@]s-h$D263z+XA=!LfG;ac0L|.#'8BY>bRVv,Z2Q `7t^!Nn!j"uc$sw]0;(bkJnMp^[P
L<bPauI=@zm2L=M15Jmogk8uYzd2:4@!K;{@+	P},dn;3htcx B=UI5olI@gXcX~ rQrnRTyeX8Sj\LyUj(uY5a76U7Vcy><S
u$onSNGVKvk+o10i;YL
bV]Hh*Y)(uy`(|tC?Yc%*8j^OG=G>K*q=s!hekh3CVN8?hGAlITX^b6 2K]*6O
a,
IdO=t\ C[= Fhq+0Ooi+ CHJc'R<y> Y8N!6qG^|1W|;QKh.-w_.]lx.iawXv M3Vl_@0a@jTEGzAz)vVMyiw\g6#x01~XtoFL+<JiV~sX43+%$H}xVL}d\d7"XB7U>z]S>Lc2+Wx>DoltQ6P`6+veS<Atxi*D#//XdHEJ7/j5`@	XgIDj;M4_r!@Nve{yOS5h*eTJZsG}wRTx:R+*ASjJF6'D(@ gZ:r/(HGe\(wUyt{Q>CQ5Y()8tuz)k<c6_u;^JNU*8-T}t@0r?rg[t:FG7U
'u1VjLt"8GOVA0	!HVMa<@Z}%	(U[O.'c`OmAF!kB3rl3}zR+J&(W["3.i(=07U=gbp=<dSL#/3@sn%4I$T05aeu?QM6qaA,MG'|O
G"xC8/O&	|Fs7Bq5P2jd &'1!/"_wsXdT!!>RGkk_ jO'h]zu[jX}dv\u&y{]<A6A'&l_/BQ(8=TD*fBhqjGAvF6>qH4,36l{pI#QA79isNf;Vr*$`@8gmdQfcvk^p$^#a_gS6)u}^iw682	z`$psY8e+2ys(`gi>|=UeYFeD~}NS($y_p6aR`fXLf`Nu+ >O'TiuXw0L	7xk=4z+)aAZ-_
qu^i$zW!XD$RS$7i3mHj	w4"`pQ
EA6)&fEl<rfqH_^	#H]k"
mqN:/0;('K%;iV!B7d}X.tY8gAN+v@)Qt`	Lm*<#jo	EylY+i0&b2)2RSN6AEpv$EI5\$V2`!W|;=BD6iPq
53>OpPj@F5:I/1P2HDNF|h$/	/8j<W4ez9QC0H'~LT	a1o'~m>-nQi4#Hpck8OcG1-MVGEZtw_ys;f4v8rw|'y(6Amkn>W(c%ocT*t"6>'O<wSYCX1?ogA
cM0o>'DTK`*`$W$B@$hwVEMwtOAp-bv'.qiPIs{P]$5-K1|UKrcFc*C4z32a1*H8`f?cdrcO*/|+L?F[8Mnj`0j/c+6?u8hE:aMvm/M"Tjt`i4ddoc_
Jk/%%^	-|sX$GB,`QP2~^yRsrFH$Znl$.l3/(sD 0 2FGp_ZV!9_y!c=7Mx5KSFgDk 7N6rcCh2~:l|4:"2Btma4M3Bn,?ItEabBku@9|%OizJ5kp@YrgNmkK#QtZ-w$!~g=IAA&Z7~`rvVd=OkFy1@r '2&G{@~0E7ViK gE7[p1.4+HF`LGS.S^S[?)zd0:4.M&%U8T29.~(<{J*"wVA23U3}%}&>PuW#(aXH)ahghucu$H&BQzoLRU"QrG;OGj'6p68#N>)17^:JF5*h,|qN7{3Ph/##G2k*#]TNf]pr\=GlGJ6*D43{@ZTdd<U-{:)zNQifAv=Iu\hD1m{3WSM(<*bq[sNQt{][gB2\n['mc7U.">;QKyo5QSZ>&i_C',3
W?g
SL^v3<[9-
]K2DbA^92
 _oDmZ0MJK6D#R4pBT  ykipHgdx^q2UiA4~!^('jTJ}b#l4Y;8z`p|UJ\1A{/}bXm;;Jbfs4a)x1(iRYt[qUn=.\9lvpgvPqFAop-"x9m+e.#u?NgN@F$Sg-KlM73t@pawY%e5='?V	9==8nG;~M}-Pm@f-h%=TL{zeR*~>G<1Y;1k@_DZO!WbcRZBKX[qcFuS5[6A2^X$*EsY{Q(-zW_o|h>a;|\XF"M-SI@qrD6~4kku=`R($6laB{SCz7Rz#d&bur&Z9=/:] 1[I/Li%"d'2V%`qy&OS	J#Gj-d &S.5a,eK/)P9xc)ChH.X.ojMDFE>!bV@@"omx62H/#(MFmuE$&bOZvLXU.py,r[:yWa}Do'_X~Gid~;CzsSHFk)|:|ILvB/\FuWV?6R!`}CuEQ-%]"7	Ncrj0?LS1 '[&3eRDJU"DvB)alVE5<4+Z$I\'	k%Qh|+1WUAD)!	IDRoJ,U|aQvQr+	*w^!yEsqjhZ![T=xlDx'JT5:71C9	ENCYS'cO#S1iqdgf7qCT+OvuHP}wMtKcA/|/m/\RYQx1Va>lL
~}=UpvC?D^;8A;s_8-GI~>YSl4 qmCkO'n{8b5!~"ac+n	sHk$G~PHpSQizr J9I~v2`t
R+sz8}"1f_0HUt&u%E0,,;.C,13G2@Z-zoiWGRC$J2ym7%T#GR&8is8XdkB/ka~r%:keAn~);`!jo;c_qC@0`5<ZO
 <L2r}=t&ceP%|W7jruB3Ds.f(?COO-*8~p8-:QHSxE@YwY}pRn^M&>J^(D=)a Fr.s|l@
A1M|O"w6s&BXNV"AG[E?zOtx@xDs*^0wC+L7^@
JS"wmt+<Mc<t$hXWG1VGoL!kmqKGv"@x}M|G|ykVy\$n=|%vB27|'l5y8%Jd6+aH
2W/jU,n?bsAjtNB.#1KvhX^/%#9zr'W
(	guBuhuCUqT6jfS^Y#.y[N|nmhn,aL
GW><O$&b6zuo+0&n;U.)[GAZ[P	7"(]xMC3.Q]rVv0inUYl'Y<0as))]LFW.{10eSI'^t ]A1SGxcvAoef|J]l "MRyMrzj4	8<De=$8WNlInrGZpK.B0jQxrzWW'1,E!Jn5/j o2r*VM}bc
M:_x*G"@oQV=?|4p>i4Oy[]6BQga_b4/snF~sgg=hx8.=M*U+R{`g.p5S*Z6/0CKtJJn$D"u*{KZr	MBl+	lv &N0qb>_3,B[3,LSN`<
a`bwKlP7-Jm!WC5G'}[
.Y&wCqWg%x6In6wOx4FwZ07I?f+1J=@NSKlmLGtK?hq+kusOgMVDg9J{N5RWC`0\ShrsO}Yot4Y@aHS`/Xo\<b
6`C;mYY
<	5H+E,!#oP]Rftu	,:F)w.FJybHediS@~el`QQ<klETf're>gFe!,D"JR+DW.7YrTF`Ld}:8mjZy>+f\@]?KPQLk(b_=	|/{=Q?21V''`p8u:2B&%1Al8^43TuULI"U7"%n8RaR}OIXLW Jf?yym8%jM[Lfp_L{Mqo<K%&zY2I,;$<_Z
(`&PC9{Jk,?r09jvn{BbG~Q"`E<Yq>6u,VX'QB\*?ec$wJY;`6wK2>d&PH<zsQFj&{~[@$Q2T8>/Ut&Si43]1oB6s>Ooso%0^bxz$r:`k&EXq^V0M H
R("8]~&@[A/aD:'vQi;Jw<+mq_},F>_r~^ik+D%a(\Sx'c9cpYB[.oh&fSOM:=vMFOe+z}?vDc !b7S/.HfthR"&_0+LHE;R5V(6lUA	O/o;j|6YP{kJN5HJgG&Xh-m4KyU/%9cz*t;-(mSxvwG\/(R[0;2UQEu8|>j`;O4uMN_*6]mL8^KXVshUwQKv,@S6o{WbgKJou/\fw`Rv=2NMZ cQ!o's&d'(6!o5G1lBbCzz8H?X6{[cG{=&4221c-lJ}V50<-fPayFdMD*_h!lFwx.)(r8!8u'z^5;@Ce8G:ba?(axJc2uQb%~*B8@wxYU{V+EsVWj9Fa8^$@Dw
.QJVpV$FYkb1:m}Tcrj2W'K{
Op{DFOm1XVj=)#: [6*X[+z:2GGK&J(%5`o:MPV+6Uy6g py'zfD~X4$9fmRlWGiE14]bdqOZ+5ng8i=XD=5U*O&xvyw=|AYu|1T+,	xG_Y_GBFO6P'%%\USd$	F^#v<HiPhZ5Ap~!.[CesZC3AOimB;6J#2<VTg9*l&k7{Pu4%(k,l@B/My]<x(!19Gho"H	ds9TF9@(0_e\FP
;w^&JIDI_U9X75Gu)k^~@Frkqar(L?7}#|.M#\{{iP^Eny=z!{Qw'_nJUi:(+V1X8;x53 hD8*hQ-TFs8r;wQvJ<b5Lxi?w,;\K|_uD@:6-b1307:ekH<Y.Ec*hLv'OkK?EP@=EUr;T3DS/((x\q^wH^a\rpxVYL|z
Jy%X?7{}(
\qhRS9up|..}3vAKr4]oW3D$\JEy9U3VDmS_a_H$ie%Jg1?;E*:=66A:7u!:g!`Sed};2:pgyHW5:ya0APT]zrfYP.v:./O6:-FbR[HM
mTZ1oBkkAN-]g$51LOH}'5DN_ {;LKJtM K{w"WGsD`=cWev.u3)Bz-4HNT"x#O749pZgNm 2$s>Mz5XPj-]#v=>5'P})[03O7OVzE}umYxj^y</eH,jw>b%gT'!D/HE8TQva49/&G~{3=`=qO;\#-D%/%*"uTvB&R^'I%f"Vk4"cwZpP3g	t*+k4aK{,U5QHH@LeR;]vT%$By?QN\FZs0[\2ZlQg3=8EhoN!{}IL^w[hEp<XE'dt^}\ItRI
}5kwy<<.Pl8e86%MV!&-w	1o"#`gP: rS]]8QDKRM3uzcVO&^IHJT)af56+{yC)W1<nwG#x+9|)2e&VM#,v|2NI*Wy!k6Ha^X`i;z?6+&;0jM>pi@]$-1<}N3vZ.8"G@CMEqSg:l//>>;2chp{b3Tp^|/T~i0v@%re%[S~G`8zHWKVaPmH{'UBNCQQhKS9-Mi@esm6N4#_Md?@ndnA
Ug,i^] ${&6}(BdML|	;5zf;#H.A2m}y5JU0jWYJveHJ]e\O2f+g9DS5w93eJ'-AL,vD(p)Zfs*9,o%(3>z+AW'HRNH^1DYMG<xWi\H(AFBUBu[DRwuLBwe-!,
QlBf#f?`?RE~E4e_7+b1xb0&/gV\HryE`UCm8Ey-$uxgUPAL+-W<T_P^NlTJ!.(, +]=:ao=2N;]f3i&t/7/;p_-91LXurF:s=SBQzZ/oVdM,cJJPm*G;pSB!{9s.Q:24b-@X5X,W0a&Y\1,I%?:
&R#R~3xI3@Q{(p	`CdVPGR==-kjwoxlHQ3R7(D BoO}}KGzU
=!p<QO)Ctre0
=0$=Qs*LwYs6ZcVG(i!1wNTZ^/
-O
.f%V^O|osYb0i%BE'XzUS@k4"a@^("@3eS_o%^r[Y1zLQp3J]2sym7/5\Ek!]N&z[=Ve |u%8:/Fs<6I)$6kmwNx_G=bp(	@GAHc?oU$"~Y.Cb$`#{Z5Ki>v=4>|Km9_ORl|JI2I;ieHe}bf2g{fzDFcM:G"d+wPiO(~/\sUjs\jt(4;KyL9.QFKrBs_W*+vira4/ikPTUVY AyK,g(XSo]<~E'"J&(nKP7;<oS~7`|!ja(-RsQDOA${g?=r{b3Qv})|*]hSyVYZEVp4'p!-p7I/iE +
Rd3)HR4+wC]K="v*wX%8$pJHT_i?_9DNX[mSTb3=8t?p^nbLtHO39+:Qs=5GSbRbpa^W~Q>#"$l58E$,.P1IuzcTc'U^|;IO`@$G|R@m2]6!nZ.DY33r~z0'/iPPw<tVR0n&8o]m%[,%q_Vvn8<u[dy<|11wu]GEb),LASX\|y4$V#}I8$L~%DY:rMc py+X(,h `eh0z?sS1N5=n]s)!)8GP-5,:TI<6Hm}^hg*V45Ceq"F_"//oe]KGHO3TSP+3I]I`YZ*uXvmb:HX ?@|f/jBUW9WM@Y`PKoi(jbf1C6,lQ5yhC_4gf2JzNf:a6>}b:hS/X/W?~q>ZV9&0u~UBB=5d	egDn<@zX2[$Qo^Luoj36KM(H!/6|*eV!	WPfzuA"T&D1&MM'mkf'W:
<f:7XI&0J%Zt=y8D=tV=CCsx?{KimlVQ]	UcJ6`G2|2~:U< oC ]JsGzMJA([QzyT9Ik4$6$^X<yk1Rp@G}uXwV{F&u@|80xAKtUwzZX`p_v;^!&	6O$7djg<-LO2gGuHha5Jj8K*fqe83(bST'Y0iA$K@P
wf;+u!0+}gGn4R!Eq'7ENj&8>Y_KEvw6#schK,xZ~oyd7C:aE_54L|,d^Ty:[?$,0l_3G}	Mcs@~"' 46@B{T
X!qY.!w	J=1=!p5^vkI
g>Io~K"v,%<YX7l~b).aL/*cTl5DqCJA|r6o=n1X^s~Xcd<w:-OB^H@sH]aKTNEpM'gAH	%*a
snZx;IJtj0f4Se I);0cH[IoI)FIrFX[5h"-.|YrjQ>AUz@`<$,7FLBgZr2YI,MT(nGw?xr	k5x]yX%x8F	AxkS#O}Q2_66xxm4E`]N})fA1RKfEPL\a9mW	KNIh;wv. LqE<yVpKR%+IA	IgY]*/|:4IN7pKhNi99`-*<
_L2fQ	>y=4[O*K@}W2d^9AyWQvs%ORf@[XD<1a-u6fk<\36W5S$rd=\]eBRH]M&+1b.mGe4@17w~[9ZG-ALe>)*[GwjT9gmM%c[70!j\4)INj?zH9b:Tm>Ct+vftA)^`KdyC|s~%cD'b}O6J7CWKiTQRSc4-s.bsH<2K
laxU#^CKE:l'?7okyjY|sQ/:kV,f#wpRPLE,v}y`qTrz/U%D86;qts#OOkjF7F*~zVI+V=+%g8(dybsv )+#ec5m-YSl=]/=Rovuqd5`$5X.:Aco~KK7Q-YM	**\~Cz}k(
Y`cay5?qe8q>i\S6ckkLq[lc`3Acpn|jn8*&FJIa&_* RS2sRV/HM2MA_+#"O^7b;D*1Qw=M_({V:H
6E6||d;bo8b!A_/3\i K5pX b%}xxC4e^2W=z*_T(qAz^*@&m+7y9uQC*z,=ta(K>O\p/{IlU
7#dW_]Mw{bupFdNoO&rF6SJm
!2|R-x@5kaaO]ZO8MPAh$AaH8RuT2M9Hr8'<pZHeI={u{Um,,!	Al$`lr=WyA^\5H 0p
~@_s)7ffVtqL&j\K
Z$k 1nihmxdX#k{?\7mzFZQD&h7mu]`;Qn W%MX
!Qk[ <(a8X>~SLN6|"V?3YwurC wuG@)rmm<+S?a!m-6x>sQ|U:s.;~
F^+,lZ.V8^N-"t{X/;'gFjV
D7&v<hiR)h=-	?8Fz4xIamLX}eK4IZRi86rM{Os\3g*6W~P	}tf-%iPbQJ@Js}vcr#r@wi&+xK{[&8Ti9-6"}9E\UG}-{T-~$pdD=!cKHQzq.Cg`	O$iWp#G,!{MX~rA.nB^{qedd1g@#|nki%ZYII%{_]0+TIqF*u6j-mZ&2%RYT6cqv-tG15.-A*_vpHv\^yRGb4P],ff'
6],6JM$YP85)J5%(_^T}.D/&w(=QP0KP5	=*|ffDH|HK&A,~NWSC)1:x<xKx55<U!~lc)@9q\-eJ&{\w+C8Wt1.96Y#vH"&K*fe6*+*<p<yHST(OMFg\ZS<4=ubwC2jl<\	sd2!_3"ud,Qv-Z	r	ljLhu
T}e>z^^D%?U7'Qv5MljG,3Kvx\?x&~/ =~>Qx%"L"?7[~]"|}ktJOzHCbuy4|
1/gID#UyUnAvr3 I+3\Vu ryL(HKX#i+u"}2<s?u&py"2#Grt*(/5iyAi<-c<b6*FK;},L{u,<HMH?q>l,>%#&O})1oC&v@Y.!d=h*E\r:8V:Xr!c
$kUZJhl>dUbV4]L5g,A2P1,PN
2rdVk7mvLG7^v/:+x_)L`7Cc^T99\,`{y@*s7.)n*PRD!TS5 U RW/Q["VqCX4Tt,9/1<?Yegxn80l17A^C,?zZAM;.>ppPy)0
QQ%4O9cDo#C*x7v%d#J&sPTa7;zJ]Jgx1:LPRfgK2%V,9qRvCn-J0y`'p9IfQbu~9Y(fFY$yV<w-&\vbn@J=8gK]%qF{*nVmM
ZD+?vp,'$7&e18\^LdcRBQnR@%_Ux(f.L"^crswO-1	.UK'>3TsWua;-WkrT}fYrdzJ-PG2I	Wp&l%}aVG`h_-=>TV/ 1HwU}0^Bd*c1(t#H=*:1ees+3hz0$g	Vcic=EMLr]KV]x{]QRSiX4iyc/*)-]$hp;'tZ3km?j[bfLq1W~%"^4r#*mv3,RnG1Jt.U+I@$C8+[`9T'V<Y"ax ?uGWznyx;<a45t^V>@#.3- 
0*f[cJ$*m9zcNS?}a>0%OaZ'.WOv7Ks%M\kHj[{dG21OOcFx=SrBf1:9w6^k(Zbx$s 7)e%Yoy7=HT-hY3H&#nr#TKu5J;N[J>%lks`$NB&9hV2G^$<gl:yLAOG:0pnO-uR3(HE~IJO?ih1 $`"2K@a0.wB>m0\xk3?:	$YyT:8BP46Xcg]&Untjj0A(~-X!YSnk35vZd.H/6H+X	sa1n0+dqxz\p8T&@dN[|L{|4]O(x+cP%V?uPGVq%DrSx\5QAbv~.C.v(~9V'a!6*M0*F~,%<8ks-H+Mx
!d>gGPTFzt!.C'g!3!e GSyG<MA`oo&TW2[}i5g3[p