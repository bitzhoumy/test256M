Fch!)^ *0T>~'Y8R069-R&r\[^-e]dq|P?O72x:bvca4WrGYm*1oBJ}s^Fa&\P\@^x4I%]	>Yh9gxIS%t>3]}!qp@/l`$Sx4.
"!;s<KHRYzV,|)2<AE;Z9`q>FM<4NN`-:CWngE	@$HSifgnHi+68w?z<INL'_jYqs	@~yciXcZ@@fnW/.F*f|8!Tib#U`Y&z.(iJ41\5#* :OKY;IdqWY:Ae9d$=)D&l.E}|/*g_
4N1EUS|E?T*_T1b.;E7j#sE,Kx	^Hgsg&by=ks1J)Yys+5C/GptUc$OAE&u{q(A`	~vve(A}"Q?4yU,_<IJt^~pxL^FT}s9Wg)Vn$&>]C25vq95@0&=Is;DR7/"/z{$S91VnJMC'N!pgM
pf^Jh@N2:%W1Ya,6pl(08 IS&8,Em;n (a5Bp3("P%bQQ]L4\wayy#-U1	|&h//`	iR[ 8oQx4^0AHNoa#q0myh
tiT+[U}	&Umo!H|j"C;Oem0NO<2kF\6H}?~bU
?
_6|zj9/\Ci;J%@58~	y+,Pe
|L8wM,}C&Il~BC{0}=IZL	-Fc=t5ux143$R30rG"4S6FL|3[ 7:khv(^m0yhu],S`=Cei>gXQAnPhTFVk!*BTd0L}RdwN\(<_.<B(I<`T'V<C*A8oo^;'X<du&C\vNaZ8RW}RgXyz"
iOKNFA-P8>)_eD
P3ao<j"S,,\m tb$xj&LIAME%S*YRc:#@L?4n6}w	ub,	Hst27;V(YG\gTX&
.`_9&.QS]wzm];,B6"=m)'NylYA?gPD0EgX!4+-{nRtODmP71I7h|wAJtQvdxxV<>vGKr.`=C?\'8eI9:5M#'InwYiel,~%A@611vJ@(9nCeq~MaI,9G4v$xU']MC4J;.5]ps/qoD$Mp9M{<1n-oF/;QFzo%xtZ>\
*P'qc.GES`Ii-#=Va{U4>gNgts~O6|0Tp02j<|( _:2J'txty,_ :TTk}m
bj}bIAR-`0.gOE_h DQnO^828<ZTmNs8*:cb>M\+w6jQ<6rv|:+vak.hv_}:O_*tfF<4:axm%n}N?aMS%@2E$.TS!"(.rA!c%L9<Gz.-pYx$RwBRX>-H}.[x32Xj
_Pe$m"4ogWMWes7mJ5;dn!GVi0Y7z{m_QtCHZg]
 rOBkYv}tBLHJ7m+A:c&HQ>%(c$j[.beqDp4=Fv	b<<k~nm3B=D7/ud3wY37Fh#GPkRK'(zcC=y}oN2&GXeY6?I%9>z;666^q^h]TLoV(i5A>h*@#upoCvLa4iQqk{m
w^)an:#fRFSsD\eim@e;E~	C-efQA+sJNMF.sImQ9m-|J.T(fv|G_u"+lD@>?{Tf5,)+#[:jSX">OwgxAwM=D'^W2?]9c=(Rs4, oB".D3)y#Q`Y,y9.:YSHj`{?v01J8uDo=R:<}$/OK@nAY]5D/R*t7B-1R2HDL_A\,'}
53UgV2~Tcfw,%mZWUs}#H@e4:fB-,\'no.z4f^mvq<%T,)u8fyS`)A\2&0M}6EC\1kZ'./T@
]rAPU/z=}@<BJ+iQ@w^q1gwy~*,8%K>c7A{>XF}6A26w u3=];&&hS`KG`7K	z5REY<bpU2L#{KE.'9U?Z{:CNn-l~$%kq[bhDx:KObxepfHM7`N[`i[)/>4/?6p:"=<B8]LxN_A(:Y,Db!fe3{s2]6&VR>.}-(Eh~}B!$+M ;7AD9l.Fo$vB&V,R*MR|~p(Bkye1U~T~+Gve\3D1'/lmz6NH_H.IKxV\EWd=q\k-O:(%2kiB}1Phyc`dKPjrlo4z3sh|dP]j},^=i)$bi:3	0K<L(n]~~]G46	ly _A"lB}4048Xr S;iYT9r(,3cQYCY=
yW7:NwwIG|jl\{_*Ln[~=F)EIV<$#SO.LEwMuLXZ|K#p^eM^;]kA$0<bM')Y_;"m</Laz[%y<rXGjDShB,aTfMBQG 
	)w?zMG+/h2i8dd<log))Tn	wt=<
MUvq~TKp@nqyM u,KGgIiwej M]Y8z3|P}i*|7JB08%'9X6T;>tXE1+Jr&cn`o'(xnR~;WBaxTW@Hd8?2qH>#j3_*8Uv	2RU7JFFFQDv"NHgG[*"{ ;v4$DOH0v?qZK)Z}6k.|jEQs+&}eeH:,VaMN=cES9BZ]}:`]!i<pnjt,}E)\294Z	{%%$ei6d##>mJQ<$UQfa"brw*Qyg	mzO]=r*}KBa)9wruy:'9.#'Jo5j%^YYxYgF3;C]rMe#?!@LV*gvid`Gm$71rGZf&OFL8a%+=*}LE(y@P(_<9s'Tc7#a@I6TRC3 T	;?KNv`N-X+:e8C%lk@UL@T-OuF_.vc;TBw1?,1sw
p8)AVo!!z>QG6[H@yf@dCV;Uu;\z0Y^]tu?Za#BL"(CFq45B&lx)kf!<KZjk>C8wo!}6xGu)V[,P)YVsTeC(C0ms#,&b!dB>-1[
,qdY~k31 5p?h<oo7/vhAO?o]}_{A[P[g:G` T][5:6T UOt''qp]$;7f[EDj^677?GjYvOQk@2L2YpQczT:w\b[6C1 _',\,v-[p>p44{lx%8{pn"sd+2ODfnzM1q2?.j6pL$BA7 8
1w	3:))~6&`3xR8+}P7q``pYB/r>%h9;DNg[X!&-M)@)#0Ia`j-,>N6"bp-Veqr`e\9:z+%hU7m>0;~!O'p!b/bF[~FhatA':d)UGvWP
_aJLMgQzT&X\U,LGN	Zg-W`/{dFKDtYn;e;T8-;Q"y=pew^b(HN!>m|9hq0r\(&/
934
wVA^DEN/(/GR5e)VT$LwgMUK?f1Usp(LE}0"}&eY8%z_um4k,@o'eoKFh\w,phM)<z{K "G,"VH$pjng,bP'k<($&yADq!4r<$?3}}TY=,Fj11ST;iBH+p[!F3"}kYn
}f=(K8d~X@nP-#JO'>\9gr'^rH;<6Qw1#X(Ep(Zv$4P^i?e*3u
Y|=cX8.!]|Q-&):D4nl5aB(<*TU_Qm/]xcPFC
R?q'y(<Vf\3"+{hdCC	YSaSFsLHS'4vF$o&O5a/`AItkEW6[3|>H'G [r+(I^Oj@d1d7A"Z9I<3Kn#FW9WV
ct@Qr\w^Rt\6Tu40}\h*gCrHpL{Q=lQGo\>3AZ>[n2}Xd}2S`	gBhBSQ;hX;|tpt{u@<A{YEfQboJGpZ9Z})z	|)} -C34nksH **J])YhHtOK9XbMSq;6v&"1};bSpF},^a!$nB7`Ya$FCocu4x/r	^]/;Z3gbISCEnu3Dh[o`Dwg"mV\N,4<CI:GWTa.0$^'l+/((@&={[Zw>V-xUL*h'sYF0*B&cZ|;FZ8BGxoOcphiF,>obDzQ`%q:4\{b	hRR^{)L:brJ&m:9oi%,;oiMx:<bbo*kWYm\s\6lJ[YVv4 .9<$isbK:Vg;S]}w}&ZpnpYQi9<<]O6*DvpyMTm}VUaq(R|#.%K}[w@V{qFQ%AK{cK"[ZUu*_YVPTIURm_P35)FZk1b=,i}.}i|-8*4&OOpJXm/Ij6k)^FwTgQ?]pwQ `Ui^j]oI%x~i.	1G#$)cEKrb,l|:SJ>2u[#yp+A2B1z
-a/Yx2nEAK,9c =	xu^ulJ?&Es_ERnF@@G{(%K&/.mrFm|-k8!FJq( \/NB=K5Rm@	c7r506%sCC9V ^(oo:v<qN|`sUfGo 5Zy'z>$kCMn%<lB_c
?1_C
#p>E%1(!UQl~ADJ6Y[~T!;I*"Cw<pIg$hC79SXp*lXn:`Evq!!7\$cA)Q|1DZjY4mJ4Lx1]g,0O=p'D37eLW5L*lzFY
=*M"3&Ta.d5OakTD:=XI\|wtpBKm5E+8y;xu	BCpSGnn'	JnlO3$|SH`VVjgf{M9P0{hsl}zzn,}+otb-<IN#&iH'22O9,|iph=tIgHN*-S	ohYd9fnyy\f{CT)`.JQ6NQjav;bfwcvt6hyD}ZBH[>I8!S5z&(Rk{Sz,P^-x(zJ)L`I=SiM 6U
O<@DWs%|:.|n0:n>Rb}G0XW9wG9D@lN8^|yu+c]S/L'Tckr?S&89@k)/F8Nf4^|h{1mxOo-f9+	y){zI@oLPaao)]y;iR~z,S?z=ZVU`S$'kQO3/$iYA7(yR})]DN6RqN&cF0N|qQPHq2/`cB=,mY^GRR)sTrT["V1-RikQD
:J$3aI$AjkwhYO/{!|{9":/r>l8.O0Le'6+*mg:$}1PgmhCl"A$6BvC)X2^tjU\&V>(~*Y}LbE>lV%$(v%3gMP8Rx$/GmSnOhpo/oduvhG}oPt?,Crfne:)j:`;6<*ic6@|+"Lk4G/@)z3Bor$c[lfNmlCL7x*\5	.v/*]AEuw#\:Cz{4?o}n|oe=9]b~("GQrm{gv/6k[0%yX4\^>g]bi9j=mRun!ID%{+FI>>OHQjhd1]d|`HX"u2-XA h'hq1yf`_@WMU\:;$iLb[_ec$U4S]#=Fl0DsDvb?JrCgMl~G9O=m\j fhzN\x##%+xEhz(oLVS
re2'J-Jo+?|#QP)@indo|6v@^qec9fz,}YDf;Ii/H(J8K_w[#U|%N\d$.<m-.DQA<-Ki}K8RqY!_Fz.^;]i5EM}6k8Q?Jv
|K/fz2A@++U{KMxqGL0cniYZK1O,5Rv$e""~+?v4DJy'~oUN~{!0"[uEny/
f3wrsIl.?*dK${vg2,J($dwuF#!-pJ]:?*|N>Fr1]3|	`	R/kUDg!.?!Pd(mE	f?!ON*5b3m{rhWT3m<G*"PpHY2R
!BUa-	pQ']nT((S&2NQ[ZULbO[b22FSJse7BeIk'G.q.*u8GW[13CQY=h:5R):Vz-S0N@qM[9x.
i@L;FDn\&Db*s[2b4)ee]6uD%:NetPf}<{-CNsIMIFJ-U$O$@
*4%vG:y*jM}.KE"84QVy.4<bE#NZ2vEw:N0m7&r	uKz4ZUG!OlfLjB1WsXA7hLyST5q[f.Z.c#2m2TRz,b%Ga-x~c!C"j&mO(-U<3o\kcwmcai5)Cg^md9MCT dE|):$MXg-d|lq,	fm%P}}C#D'O>`a#V?g,f*Qsh*~vD\)xN#D7x'?Ff*{k%vs5`~3p"":X;pSg@0YbAAGrZ:ZU<k!o9p&O.Zgu*fg~&4<>MUCwkwVyp2m~Q*q,C0Lk#j]_~IG\;iX_u+<v$IT;7orWHhU!)>N(RR#BQ-<y8DT3b5L6nC9`tYSqsUAiUb}TPg?)YCtiX"@#rCDjrdt}hi@hV+V4_/wc.I%3i`i)O[XUlmtGy{o6-_tTRv4"s3mHiQMA)WuBB8pN,5{eraWVc^OU2&%Q2"B	!l:i5x+z]#1G#j;]K_)_K-0ieO,]@mZyM;,D<?D\6"J4n{A	8!adZKY"k#_c/]$"v}uSURA((mY"\(PR{c\]XEL/8%?,PG?.G+%M"	nqE2O+23xk:#iz&..<5e|8LE`d^>~%XUJybKye0pT7DA*\Nu6mN")t2GzR;<oNenX"}K_7+ZM0eAlS(CFbhRX`7f>#i}-7~j;k_7AYILQV$Gn!lN8}LnAWa5gmwiACdu%OvYHaz:bI/4UV:Ju4.RseXExe!n7Y&|zST<J""UG8Y&o0KmbY~9&T}?:7IK
aj?-t!mZSxs)`l8^]|MdfYx*/44djw[FotfT'(ME^J)i42pH"@$5Y6c.K#.>hTj?oO6)[@8@cRwj46gR$&">2	P~)%}zBe+h0^5k00o,}#e[U{no6v^<(4`PIbRv
fL*w@H%)-:TpF)^Hd&ymSYU^y~?P<OE7"(LC1\AK]1^S|[U^;Wf]^ie}8y^e`l8BO_g}3vSfNGe?,UO)ME1{As^t3H^v3@B@6O{9	=o
q/%RK71aa"nE7aFtND6\alhTd)%4u@lTA_b.
=!VWJ'OxPy6`p="e4}0V^J
1"6.0WeS+,BRRdjte#/bmhT!B*SX-CL[:].SZf7w)V~n*)kVF]sgY]R;	fjp%)ED$.Ypc'(VI;fh|3\HYWz`d>9k>kgb~M*v
K)Ey}oFNt2:>F`CXVY7np%I8WyNN>oX\uL5oX{o7IKSeOGP|/MtXRrd(>7&M?DRO<|p1Cmi.p:9;q=qns2%^xUCV{=,p0_%J`	$&y:3NMA~'!!E:SQ([Y*&xWwG|$#mlE_i@^;|X>o&KlOqccA[5"Wwl>L[[u
PQGr'f&_DGdzxf9#&m>:o} k*-EbG1L;z4KtXs'sT#p[VzRcsX:!I>0.+D.6A)`sj4<}r^p22qV%fo7rjq3" :IyMR3
 c i!	]Z=}`=GjobHHpg%AuVK#cAoiHs0FmSL)!&FKM[)UXhYhThDS3X({u'3wk(y(h;|*Pyb7owYaA*N|T24PbkX'"MEr1OF#b?ps`W!Gdj+peEfb_
At* LSCq)S$L)n-nN~?9y{#<}/D'}blj/BX'DqSX1H<3P$NTby2n=heE:cO)l!abJ6&1j68CvX,`kRY%-yA,iNjq3,R;XU3692<`maz{*o9QS'-&*bqlzS[Rx/i\6);)i};l`P<<Y&}OwT.{lef$XZbm`vS|oagq0*85$#4ziTtA/CAHZaE|4CY">mu9|Py1iX+_;6z{U'\Lvx3u,94z&n_nj'tMIksYhGgix)PvD/j9FQMOF'9$NQ*n!zM?~/K'x8;Jdo>}+$XU:u[*8]6-NJ]M`L>^Y]yS>]5`@:g1kd>BhbM\jt3FWCG]Yy8Iruy%(g`WuDF?-C=*%V\38of?$M6PJmzCKy@?)_fn%*U!	.z*/S]jYD$K!O{A9#9UmibW%`3br~3Hm5*Y>K1d,yg`So<,8(Gtk	?JYzxo`6?0	H-)
wLwMi(Sppn-|[>,%^_-&Xc!<geS=^e$y-~a%-<#i.k>:g)jK#{5]'*X`5h>KBKxmO1g=c-d>|Zb5TcHRg	'.d618#9[jUE$-R)!_X,b4@
%rC C32'$eM*E,6YB
\=UJe+v_:*XP_a'5K9A+s~p=4w*~$ UDtQW<Pbg}kN-Dg9BQD b}Z7Jr:=_9X1_MbW=%'k)wV.Y+3Q8Hs	IUoU{\cG1?GKMVOI?R@WbxdpzQAo=1}UMM"Ckn	!(Q_!#kTg01kcRfGl,uFA
h\g}2js50!zP>rCf6PnaPeDBssyQ`a-'A1H;.E30X,F&';{TT!a#(t%	N<#Vp)Q`)AH19r5P/YO2Ur>9bojKUR;BL^8#yMJ/95-IvJr\j`#1$b$6['CN?'^`EmyfeSP#m-!_Ea$5\LaCv_H^r%Cgyu"g?X=f*	B%Sb6&alo?DfCmv_	kws'8*;,{7i}
FFKlo*QvKW$ss#v!w/#ZxsRM=,+fO>dPCB6GC@vb*CF>'zQ-Pet$#TiJ%ru:d9~`&I'x}V+-z]wPo8Paf6%}z&AQ|lpyz[4
M,x`'5c7p(J_?0PkrxB2M+V oe[@||qt@L6ERa.cr0:DCdeRGQ;%3ZF#$P vyg{E*(upvBmr]iU=7w'F"H#*=PGC	QcCAU5p/&'5,|.{D_{;N@
*T~M Fj3-*E0+;+a;;r_c='V)OpCrWQ>zq;.Lek@b%]Z{l%/yBj`JK4QL$ran)IKI";C0Ie1!o|^"|svHF1U[ceD3NT3F=%"8D'l {Iw9c2+	n]A?
Io27QX}wGOSDQTk6i}MFu%9<Qjf.O%Ymcr(wEPW2SJHk2m&JRA&K6{^[v/72(emef*.JA,E2H2\g7~/wI0lOal-*Ky%~H,1-N;4m-I!>>gSpdhE(Sj*#sL+,K7&)0"\r)*a#BOPV]PZ&M0$Mo#b@}cSj@#_YR"{XRJXpk^QQ~ClLMj6J*?|3~a6hfh#A9mx33}E<e[O4&#9u<}V'X6j<ve1aZ$.]u~]o&<Q'`YIi?+XxV={^M)zgl*U""!jv5[I7)95u9d{`3KRD'Whx #bNz;2]le/HrnVNwOX*oU%rVa~eimlH(^C*eF[ey'1gDkIj(',Y"qx4e|%p>LkrSBvS'6+F<_T&P!%85\x@9s@j;b!&UreOgKpxzw#K_.$BfGc[`VG~]E[E'!'EA5fF-e	;$npy#$]kV_FAypGrf-~>=se/6Rw?ZbxE=GH{#c}p*,YF"Yvi8z]7I#7~o
{- GX/Zyc^>R17myu=G,v_Ei`4%Z6SgC
Nos{	@Ba}HF8NCw1:2@8b,&<utqR#szhDOTE"QTj]'$n >9;sDS [?>m)&\#;=Wv	VGFv!?@S)eE2lfXs~:bA+5mb^!^1:MFH:glB@MW*|t]U+f^:,"x=<vVBZYmOufl<#N
Pp4NYF>'{/,iEl!{)?2h]l6+3G8=(kmEx;9:8n\1f=MN^B=->W:h,`via8>+uCV..#$ckPn1vPX1,:G-o*l3Or?!(3x(.KhVnh'Xi]e|R[W(S8UgN*~-F\{a
&T;7A?0SbM\t\~h|dkWZCxXwu3C[N-TgCN,ew8drlXhF.m3%NZXwoK(`jf|Ojf;#0 <w# ie9U>NkQ>ENnqJRBf%f+RJMLR|O0]UR>cFz,#3tdBR*(te_
jLsI~0EOe C|8sVZ@F|fmEB,>Be[/Ly9U1?{G2-6rNP AVQ;?6z&?br^+5.F3%":y>	Z5NI<6n^[TJ?\8IDJqFZ<?pQ.=J,g9W
+g2>"w\PUn@zO\-t(&7q^}:TCNp6y :.I(HNa]&j]O7Jmg<fUht%gW97{Hs$wl#bk
^T45N_CCP7~ZnMzKEUFZ;PHE>(p/Y*^?j
lM9,Hh3__WQ.%5yu{s%M<IyZq%GY*e.X9JD\do4jX)F}*{@{|)\U"n%7[r{vlSwR?=$"Nf2"R]pBBCS9`"6_!=q$`oE<dQ/M;nV]wkl/Cvn(en:"sZQ#ZE[VC"DC>Xg!o\(CVrgsrd[U>ed+E-k
nce{sNf2=}$.*Xcg%a=p:A_ND2z%GUX./:M-U*;3X9Y(9`ZYQwDEH{e<]yZp?7(ypDIbZXuN^zg';[u	!_'Nl}:@xnBth9mP4c{6V^>"'F2I\lkHKIy9/II](6;U6qL?OpRF_Q>WU/0&qnmeutkwH'\prsM~9o@TLs"Q\M]B7T>=CYJ"rDu}O|;joL/:>'S^gZ6	_!g]+wcKv!`_e/2?4CAAq`4=>zQX[b4'N4RP
hOCQ{jT/$guX[Muj$1:{!MgVmKoJ]s]h{iCJs!.9k}TeF!8f([s/CYP*_L,roNRZUnw&Z\?6B(YcY^hTgd-%Uq4}(fU)M*m>#:rR]yawY>dsdSEq>4J5!)'s%Lnd;Ft@^:VI-(R7"e=O6;rSL=?ov<1/Y*q ZiBXuXR
"5_ ">gR0)Hz^lR&Pn&&L\_6u]aJ)fc:rahOe"#56$qQT6:&2p!y]#JG0^WLo[|dTAgWhJR_~7J+E<08~%'VCJ*J-j8mZ&7kQ=Ck_oN{t^f2</A:N$O/dY5GzFAkCs_8Gezv\t)cS133;Viv#K$TJq[J;NU[$EKRgkHr%_7KGzs7G!!q3hQke!T<
LSVaMa ?@*+<HJ[f,RSP3K	g?	0DDCJ2m)}I=ls)ma!P]3?x1)zrtXy~BT}ds|<"&1<wG-~S=0y=e6S
_(+[&0GU9r]a1cMOBa2W*]WQ-9,Hp02c#\2z:p3N{)2L3t}l(~mN[qV%	 '8:6rTsI@1F_"gbv>:9@7K~G^LCjhre_9$ig|p3Igm*5-0
:|aD~@Va;^a8MXnrje{%%@"DNi?n.C&,kotUZonV3
&6N@I.n:}ZVm7ZI.\^et%tAQ22` >V%MCE<;V2Xe-hU(	rP-Ea>Wa1668}pFH:YLBvt$LlGU} {**knckM
!pfb]{$;
klE{VA"wVjW[5jdrEEK!*P6.=dYA9OUA_@\v]Q+zEi!Kwi*o7SaT7cfgmQ*{[aTDDH)U '!2ScFN}fzbyb`nJ)In|4Jn[>^X`qE)RqE^=~U2\s[(]j]1HX*k4u) 2625H#CkX;||:_mv:IQyY&g|/u_[$1h5Pt	Z67B:MW4C:=,@x<s{A03f-jO.mU|_[xh
h  :+[qGH|2{f>c?0`Nq_XISC$TCw,Ric(vt{-ga6Pxx9jaj/6v>E(#$nboYje
SyTY\oS_7GL&9Q@
4.K}i!Y/
6oA2qaSyRL{<8"Tx6FV
_EOeh,h|y9w\2g	^H3sSe4v5V}2bd]oZ\l]6l%U#(-R\ER[o'TphQ(AzC.<qmv4SR)U)/h6UWij<6(_@]kt,@4F~*'ni>UM)0|;;<.\56QOfB*\wD.ILT)orl7]DpNcO5wDw'td/lWg{@Pp&@}r$K#u@~JKM7spUYqJ<W+-N@Z7>\
aitNwogJZ[85T"-.-loT]**F3S9%}9'[b[J&$=K[xpy+^rR0Pu4?W[M"`<._Ifk{zvw7]w0UB^Xi"u20bN1E`S$]s1W:~g#U&'XQbIei$Eq#e u0#/7o\2D_A&nA(sn5yZK+`CPX{wtM!s>p!1|.}/+y$[wT>JF?`]O2 OM6+^{Qj~ v8.)A~*qcQr7PMZ>ps<o@B#3qQdI3IP$h4
X){bmZ9S{MS9,N"B"RxvpGWG<%}iIN'qA>GRN#A^S9!1}%q$t2HC48+@Y/Q6C
Bjpnf4IqaF5<ildhZt(<^GT^c$ w*fZ~hQp4#"gjqpNY8Dxp}R;SaV)&fJ`mohvZ6+ujO&1^6o+81L8M8!vliY%Mx:>(aY'+qokJ3vJ7sYID48f9Wd|qxb~/@
E]wwE,(BjdF+S,bmkfw$}b
oToA+Qh,39:.c}e9=BABf?a43p3-Da{9?bkZJG(i:or|O`ub.TrtrgxZQXYoxD;Dxb:YSZF)Y|t4ICf'm+M`ML\-vkPGE'KGgHD,aSYy3
/&oVwZ\$t.[}Z9?sh\&{=-M$mg2	WsTar^nD)$lvWyl(g9?]]s%!*>22	"%-q%k\'[h"
|5l7#/x^)p^{y"{eoB6	18TN[CfsE CBXUF$W78|"6
}QnvdP:/^[5Z@T1NDkPKgOns
W0VpJ8EciHr8nPjRbx~{OxwFy0*q i yz5TeWh/&.2QLoW&B?m4i?o?(^8f9t,.dXh`x)|%s/T)kHSZfEfQ:4,o|gPjj9l[i`<e<[i K8zhvYk[51T"IsoC.1F#g!|%U.|IqU0 Sk%#+1Ip97.M/7<1Bf[ VF.k~>E_Sj1:Lg5V>?,MWL?zf{[<g=D;@)L_EhyE0$V43Ja@Nwv%^sstAQ[.8jA	%Vy0M .y?('tZz 	`^m}&2RWa<J:m4q6fA<qd}H<R'+n+	swDk/[%{dHXlf)="|$FiMkW9!PsSSpED5Q%}	V(=A^I2q
qm*c84c/*"{[ =uOi[yL82g@@A:pUUKUl$x1/bjA$Sq(R%8JMT0OE#,0BpV[^yd+5t
^Sd	6/lT
_"0dFIxZ0iK?)<z/6y~]7ldLyMw$ Deu6-6,bFh<2=8"A.BQ	@S!bKgHAvnvshXos=%]Vbr:4\O0sC"w|lwxutu6 TcA !{v
9/@{F\NU_?GQiRj;>nU*><5qs;%:m*X2^_><s	^2uG&ziWbehP<oVSV+	Kz5A#// IW5\|7LzPg}iD"=0?F!W_bnQ$+daqHc'JAHti7xSp`!xdeM3vRF9tLv1D!}Ojpt)D,susyf	 g$:!)b3mymP&@116\y
9N@9Ya(Oth.=`v`~EM[	X2H=#ocm*K<(!D.rfYK[#B/U;'Eh}>kj
!R,@Y|k F \t/R[Sf?<Gp9LJ<rkzx"C5w\5xAyRXX&}XXgKMXvk9	&('!{Y|c;U-)F"QUl'&V0ppz.'PR/6;*F 8^!r)p+Hkk~2P^Ck1!CGv1PN9'AbsjS/@dKPnXa:395 T FjLN0oH}]%t0.F?bedY3|U}rF"WfF1dBM{3||4&O~09LD
k>,z	R#nZc"[X$hdo0*{xAyet2k?m}7)]^>FTAh")04z3'"!N'du6oCSnQ"NZxNH}<V|cH/T]_A6BGAt*F[Ul\wsS/r{<C!KIGfADaK,v5M	*y6Mv
"{	E/J5I|finp1p|]"X0Es";q
H@|wR+v@:HB3WrD6WNJNwpp+gxtz%zjg$\e5
FFU1fd=S6xde`Icti%YBH-NFPGaAtu@j5A-cC=+|Dv.>,[)]1K(g74W9`(\na~qpO49(.
K?DUORz.^8Wi5G.ODXT{iRt0^c`COT\S T.|0B.bpPGyn>s%H#E(J=G:]knV/zYBi?NRsX71B%BX?'iyy-=OjKuSv(69p_L);
??{@X	s6jx=^+cgiEHsf{M{Ni%@[?Im#'wV5|.AqqSc_>$L`L~V["X%iE4"di"#eOpRC0+vb,<YhH*!bp4qNvlAK";WoIXv.e8c?
p3X<7rNGw.(Te\r}=M9.on'?t1iGyXcG0Tx-{P&I~9*und2O<e1^}:}6:`5CO["Vm]Ani6%YX^c*I
gteL@*d~B[9yWR .Y.$BF0P+b@DcS/z9`:9rXQ*rz/@rjrx96p{x#qBEH\q*uc*^
>}[!iv[im@uh>[}$!wvXIr?@F
tmeajQr}i dGH7kq|M	QnB, !nL{Rd6T2`+Mha9MzU>6FCGp4-L2z(v#/DYn`ukYSsQ +V	}QQ/i-yu\S^#g<QS|v9yk7B;`qg?Yeajlw</))/3R?gnz|-OVfur/\{f.'IIhql%DW)Hn.;lg,qI=u9C?N)>&zb7|8]' :Ut76sOp;2t#0qRq=t|XL-8XKLur-I~~@?r		)'6Dqq*~nL?8[x;L19 x_W*Q	X(g:Vu].;g5]Z-CK{%aD	s~8LiFwf]0yWGpj6aMmcbD=tWRN'X<pNAeT
%!4YQ=8hJXCA[Kg@dVPE%.ML cDu"b{	Q<S,97<cjQ@5GstucSCkRw*\<IS]dU!K&<Q5

ze4In	QiRL:lM'`595!YKJG=<%+Cs-|tBicn.)$HA6W0$$dwyCgGm'82!n4iSd Q"4'TV]D`ihut8
a#!k}0>4~"r\k2\<>3h?,>Gi\EX_#l3__*'2_J79wrN,kIop|
p7<m2%JM*yf<3
qhZ&
?>4")p"-1jvDM$A8b:-sk`f97;35=W=S[euxT(	Z`S#ci;|xO]4NdMWWh1"wHd_^gmlMjVML{p*Rh
MlHy)R/D_&q<)]J.f&J)nDH9
E9	p,XA^?:g5yXyEwG>dZo|F=&4l,X;YuDL]^@`B$U"Y	
6WaS'00K;%N8lBa}_gWKV6rL	[a0vzXXR \S2JVN0D|Y"3#7CRN8mlVt~:}}$B16
"&PiA	|)XV'	$2^ [Vm!yeF5r,/$kywMV`c@|MO0=;^["[jqhJ5:4.CRFJ
pB!u](|ydtMHWzrZ)|U^{XU_qQ',toHfz3,10mbO92,>!v(d$W,;u-kF{;XyQqzP[ND>P~;;RV!`5A_R@x\e97x ]0+d^QkST+K SW/eSx3(,L]\U!Cn]]gv5sA)#T$4:*kE69zQOJ\6;P UQjG7p+ZEJQqu:}<ij70FH& U[709Tj}$M*VW9g*T8M5oOn5S1VJ$TK+our\Ha <9Y?dBw34:]/#I:5M-EQU\]kN4M&EE}leF5<*D&O|kX\]PPkRV.O-x5;ke6F79O1(zrdiF-QR"aUW)=Sm!\;/|XT gKyk=o+Dm;-1ejG55figz_pY3y`Lo&nt+ukzkXXyEIO4!:!UP6F%36OV ihwt`\{?-}6RSA&=@7{jhJi]2@O|MpJuE	jBY%,b0W
o:>:Y[`cL)aq|5KqkoCO<Z_Y;:;GO+v(R
`$MU1gT|N|<Sb{=t-KkYe6fN,InQ/u9]
;Vn8eXd/<4{R7v&
$_5K)N@7*Ny%$,@p=b~4){PfvkrEjl8NPDm:=f
jK/+Xo\4ldC6["6Mk69zSf"c,>+X&]JysK"tb3h.u|go]_Ey)3uv68|;.&^ A5u)/
ww3D7\l,S.Wm#0i6k?1"^'sOcTS#H+Y;YJb	hF>y,J= 4eSq!M*4.I	Ns#`5-RCtZ:UJjj+$3-;{`fX\	n6'mr]FsmIPz2Qjpd_xlO7i-SuTirK],n1kEJ[qRc9
u|x$[fAuj/,A:#=#g5Smy?P.F7^joAP@ThR<@UwS WEb[U6KTLSj!\D#aev\uiHC>yLGKA._>p9$M+|HXzLQ`yBKT@iT%hcV7W(h%;qJ'.S9(</^U*bH`O`.|4OtDK[wSod ~/yw-7Nq$g{
|a<:[[Rn'I.rk	#UeYbJ}'m2Dp:@.J<Ot)tuNe<>Rs?|Iw#ZqW)uiVdatXo(#hE3r&G(A&SUdkx+p0j38):GM7!?cOgEg)hJXaMLZY"/@<.E~6*TQX;`PH#saN]P^_4mNEop<uQKSxGaa]kMRZsZ`!uq&qSSu\G^^EP8Kc$Q`i.'G6b>(SanN'|gxw#
YPzJk2HZ a]ReviXH!.Qw2ZHSMqW1|`]^'[>{(aM1JOBN(X
m_,h]T3!nJ}?"YY
Oxh8^8Mg-BsE|O1,#}iF
qK8yt2c#9dA3@cvbGDE+B.is^yUU)i]c5>s+*KOk^;K0XonYApG'8Qsc}&6!>D ]":05;6MX l$Wws08DE:AVmy4^CA1ou|mT^w{]50ty|U!fi1nO.+Bf"Vo_\y$,ZqVb$|
0IxK!(_9<Q=?}E4NLsu`.w_%UbxW)&&+[U_1umur-}?$BO46q_\eQ"N^qlyn:|L8<ME("EAgH b4,bn^B+&_Qk6xs=1av6mkM:f',/~d1.s>T{L0p#;s9.6`>dgN3<\H;<BlN(hJe%c=bc l0Jc2Rplrp50{6eL%PnM$%HfK~f{mjMPoMR&$F;"&Q/r&	d!JEMv2z&sd!]
M	o-jO}!@1\J@2vdoegbS(=X&2d\T9o s%1S;QW,FkS-`?pwC.2C'zN(`ha3vYr4:(zoC)A28EG!#z4J6.vv>=wYWQ}kQSyoT:z	>83.n]S;=EcuU$LH S$L8^,BPtwrCzLgh;7("MQ1)/DFlqZ-y]H.nY5*P[w@)J	ZWy)Cw-!$8-%>z{~.gyFcla2$0)pvw,u'1aGz!N5@opY~u_fz4,1hmC#$`pm{z+e~t\]0	so`?^XO&C{W%3C2;gIS*T{g&(Os$DHyc.9?yy+,?8Rh"&7?=iCcl,EG--dfv[bS]C}CwOS8!m|y#\_'lDy;=L~q{K^N\9j)t\Me|.qa1;(P::+]#<z7h9VjBf?pPM#Z/8X suMF<Rf%@IkL$>w9DhSkN_`2'TCe7X36$|gC1j@/b@~3;~2F]]<I	"}KJ"#F<	%G6}Oq3EBaG>
o`b{ 5fRTg.wV(YV1y%m~QuN2=8jv{V|!zJ\=',-bz?P1;c{Xv{&-?%)~vDpnRP?Z!w	AY:jMqOm*VFFP#}qlMTa{Z./rWNg^f7'3WDA<NPD
7RQa*FVZ8,o5%S1imU/b0\+z
N2I8++fwI2</EYSVp@vN_
Ko-yRK<fZo!1}e\0Uz2q39yQqYWR,?qZxylooOP8MrBC,$4|w:-^$_^\l`1O[du3tn/[O_
7 "k3A:|`vP?5QUze[pn5cTA6&VVrJHK({D0_9!jv(6h`O!E~.[soB9]U[XGYJKV#&'}$rrZa&1reVLA_F)EcBl-&N-M/3]CFyWeO;I>7VYk#Vx"l9y';ORRHUCq.CYS@kmw4s~djl{HECuQ>w`n6L;HdyEk3{p4jNtlS|
g2Bc3,p]ot)]-CMJ09!{}4ZkU=a&?iAofg7$2%s
/}%Opc1^Nj<~1za7me/p\:zt3Wxm}E.bqV8{t~Q2|\)D_YUqEG$w!]zN/OoRlz^Sw'PwR/1WPk982n85Cj,,ix<YEOY`Or/GjXi|1Kr&Fc8,lx?|c/ICe<A2=B;f|Bo;CA}}
w(P4qK_/WGAxxYac>}l"nkm<ZT"+fw1q$?kPY
N^z?:g@L$H c)F^ak'A$-5il,daXzh`d?$WD \!\RA6O5@ b`&kX#?`FoSR{ RRsR$iyO/cpiTTjHaIZJXx;B?GuO+R{ZhIn1PLn-K}Kd(_w^g`LIxj6LD`1_7wn:$V;/<&ar.b)7dg,=!.Ci<M\7eoN-6hSmxUypd0g9
Ef'ol@VWgA+I>fO a6RbMUVxQ,E5y`>/(9_[*sj9Nv|?ce;_;i 7rv"jA+$ri1pY
0R9hdSq|S][rN\nu2-$,ySNhcl%	D-pflq)9Q>o;9g|3 KxF>zdpz[pXTM:xF}dSGw-R1/Y_}J60FMqfwa3=LdpAIl7UR^{vGRT> xyLJc'60R -nR;2-8&[&tBo3yR?9JVV	J	tWR{}Q^JWuoNfe>Lpq zi&c1/+ovkXY2

^Uf:zsMjDdVUxCX~PA064ue'R6%|%f5ql7[tll$r3hbu.L9jCL$_	ahAnz_	>I[RWypA:+`,\5|PAL:G5:5 Cg;{GIJC:@/aTFUb5`J<]64XWfaG4f^_n	_,Kwd{[.m	!s[.T<q;'4+DpT(6u.1lLSsjL5,X_$oDA6IHa$!&OK=g4oTK'>pENywPq`F>w*Ra"w|9c7J&17iE4+&zd	6E>i=kVM]0xB5Mj.eBog'yK;X{u>a4bDTSV1d*Eb,mFf)~;kJu)@$T2u!1>Q	JTywzmGE)9,OchLoT1SeP\:!Et?2WNKqECq[][C<$,1]Pk'yS`D|D])B;?0a=M.?0
M[rx+yMp!X%],=zgd9C$e`a`{_N2Ri^|0O4m^$kWJ}&,,2GJu#KV>RTPOpxWPxjey-W:[ZHR[8`1X9:0=-N?iY
y,pk+SE{j9H`5]Uqz0i`D#?"'XH[9${:*V.%H]S5cp|{N=bEHp1jx&g<vC)C/xe/9#>
:~I^79sk?1;)/ks\9JhaX7<|Oxe'j]vc//XuKp.e|TP{b>}]^@>}=u(nodeTh;drEzu%`	7Bv:Kj6N. (pD[Moin;|&oVBX b&r#PBF#1QOgJxa-D,'tGq&23=f[u[h_rajE	yr8>9a9SYJMg_mkcV/0O!?I4Yzrd>T2T$F%LJJXgozIuE	kc9H{({KF7@3?pLv1)Qt3pklku8G{[n
f^>j|?2z|wz Ji%kX8+#OQ<Q@%<A0^%TF[n@s[Qc8zWx&v]b"*l,
YeFLOb~`yxAsf"O0J}J!Spw+4Mkk"I`jcav8#k@}':+gvD:?E-yH/_S%lUl`ea+CVE8-$&}"!tc
z]qtF`au7(J)de0>	L4X>Aiv}IukY ,VEC"Lfi/\sF+M@_T612}Q]saJA)<{dUo |,74m_3CR M56J)"`@;&[TNLI=KIxxL@PX_m[NhIr#?<+=<<h:?p{N3Ri"T^Oa3Z)NYK8uF^A5~Iu<kRQ$	Zi6L2G-*6?8/!eaDsK*4EU@$ Oe*Z]bOW)i7iG[a"289,Q0Is/%0l#
A0X@U(8d]},?w|7/_|t_t3A>	/k[~u.Yg]8prG?NDITE6Ji4K)2Kr-dIfpD6wfO%,|=A[
oi&Je`*a
9&M>T+G)R@<?D]OQen_N?}HOC[\m=^MmdR^a*Vr@
QVw.Cm]I{8W"]`9Eh0hgRCUC?83"~EbC.?AZ	y49h8T$N`pS-0Gco[98pMGM_Q(`h;dX)*8S!5mNEt5O'bBa$9/_hTtZa=2{\@D}I/#]VcR@:v]FXb1+?(*(dP^{iy[h.Ydk$`7<=uUp;X38y?N3.(3gm68'*h2V7Asa"9Oe*V&	.kk1-!$osnRI8II!,6pVO7LP\e}\$ I:5LYQ2j,[6MoDbcPwx_K\**y2*W'P[[>pHD6./ey{i8'W2xUtB{9M,gZGh(\CCBi&BZ*DE-9OsCh!9@]vO"JAOZ<TF, ~CP5X"3s)NxByB	}ab
@6x(4<kw`[{5D?OojU
'%-IHysXC}j,3ejyZ2g_@	jrN8,v1WnngcsV%nn$O<xL:xq#VS,>hEt!Eig}CT\Quxh:<bsNR[`9O!_|~T%R;bzkSziS_U78\<f:F"TnmS?Pw\Tc]5SE_'J~R}}{9E.Fe1bHF{K'?((j0|+4B2<[u8<,qJdlsTowW.pd;:n8mT0db=|6!*1CH/sCH\_#@xggVaD'?n#=t:ZT?]9V077R|{Pi	*VCimPveGbOTI}
6EZCl	j0mjqXk~wS|2@3)3/Fs?q&&<m])c^vLVy" 4nc	@Vrso'ESuRsm\XH"KTS](*;3&7+S9W|dhq.ALxE>0\=!jD]7AEO!l3n)[DTP;ycmTc<OYDrRF1Zb'
DmeR"aA	j!97;CPD~6b5w-0btK)iX|	(Z]z)Nmr{;%w~jTB6?}`.irgB1rP(dCPeT-"&52IH$+gT`cPl8Bhv{D"~.F^?=1aQAf5D=)|[rUqhRU4t@HaXm:;NFyZJ=jlKM\2d4@ppx)~/1).,PfJ#_coFQ=Ci$,6Qp],iTm9`.ms @T{mJ7@qmu.7$O}IeKKvU`s9)K}Ci5_Z4\SE}eObq=?FUn8peapc'ziz\X.Puq-}*Q]tgu#`25}IMxmq Te\%7,wsKjI)2V+V&04C"xx!SBXX_;e<d+u(mKDe)k:O t8k[J^;/>I[`WYIQYSxjyUxdEe.jyhApbcwihb{FQ2eRXrzsD"+0r,H%Qvt%h5 av;;&nFOX4xknt
MEJp#3<N<<B#r}h:q`4[n$V+U@Omun	!3QYI--_a~D-8Zepoy^lO(0My|\AY^@7{TAjN-f,
5\p"Hkc+mm0p5.tLek@JM{2xgBdnF-r!nT?>}jcE6Ip2 ]~\$3&):wQO$	qKb=4Gtkx-P/oJ%mcf5JZF(=*VT40-*,m1[xo]'NWz9cz%]X`F:%j/6?,bv<kD"`G37?h)6Zi},va~kYG]"(3y;8X#JcCDG;0n#wt{eXpVnoN;p >CYB&#A)s\%nczK"vO:'^IO}<vHS?|<Wc$AHi}=?&rGK4_XTf4!GPV$U&>6pC#XRq+nw!% `l09\&VR+w1Rdk|WKnqI|jCT]Y"U}kH&`*7M@U|%kmkd
[]gr ZD]E@(CuF}i%I6bA"