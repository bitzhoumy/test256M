Qy^>D9XV
17l,Sn\%-z@5Nwzy-:\b.
#%\PO[ObB|Ey+NGn5|[H:BwJVq"IEXUV|n&kdos~Ko*U6a{	If$JA1)82kC(J^&X^?*cy_MocV~x&U* zIVC}'\SP4z*t0K+\u*XEFvXFAT{kmf3SneGz2'lq=>"rc97xtf6)Q]o!xl'AQpnnY7<~,#:`J)ToMo>[6\%gW;#xIK;dd*7NYw{@#&BH_rT/T
%Fzf3v>t>kno{F=F]kskj~"Ny78Jf7eG,7{Rd!JAu;JHd*=:fLK"yC1`,W3!.?ay?P%+xzw]pt T[}i@c}a{A/c;|
gs |>D(=sU?D(()-+-^l&SL52>'dn^l?*M+} O2~$iP*iKyH%*SjoeW0|iE5lT.0OE-1}p|FIG+#7#C"YI>nd/;l*6$j#(u^x'q7ZMb1i!.d"k#-fWW}}Fjfe\X	1<oW&f`9J`cQmV[W&[9 "z`kZ\;)kIF(;&&9gm,a*2_u
=bG'BvaybtwJ!}v?qRz 6@'aS;lL-M+#@uq1"#9Uxs@(
?gd8F_X([Q}gX"dpH8y1'vUF08?j0'}3F1#/'?*'UJGz=sPaW|Sm/FF'PENDs3mI*l,Z On@j&$GFTQYo4r%bySed`+-2,V]l-=,>2y2fOdC`f*4v9~GHP$mWo3T7]=:>dG/5qP0!?SpvXg0Ake~k'tr~@"LGJn]p;0rc."uD'lL,"tB)n`aV,O|v);;@-l'coA2R?)pv)e\LR#UqORm/zw"i ~ol4
&Y3D6Qb9'E'}W,k}:Hq>B2%\IU;e8Zm[[I>2d^eIeJl@Eb(/Z?g~i4<.O!sX3.dROmkVZ&GV~s)k|RF)Y@"!wxW{D".Yy>=z]&g#HZ%"OfXCx46C_s5Fn}Ou	UWFFjJ]=&:dq3+($RJS9X5GxWy7bYCJA}1/"3"} Y]pTR-P9ka$2yI2y4Xm~^m~*ellXrXLOqSplJ5nu^,TW"/#jPPw)s9/?@$> (aJn,U'Yi!#WW>#^R}2C;`BDOEy%t^Z#GLmc}>!@;_5d)u/M({b@~Vh+x<|HX/G>uE?I^S?o4vx8r7,CEAG#zE`5j}l([\K[?]#fo>r>NH)OE`L7NaVc=Zt7X37LL_0AY;>Dp03K0%U_ip3e~Q-h(St9{l9B$bMkEz}m{[hPn>6.uGRf0Et2GEOyVSQ+5[q1~g|#tO=Ti7}ipM7Pj+i!J.Lc2,v-l.PhJKZwa
_.Pn.d9IxLk$%:'G3MaVSSZ~3f4^c(AW1:Akn8+b(?7IECFsrp%h)Rn;=qih8l9"t>''Rf=Bt_oI \ '!v{<$DkCsao-'17$?OXZcb`Dnap=x.h@a.POYh9j^vud/(b9e)WBFbKXVskgT2GooHBzh&\\_zi]8KFfi}.JW>5[sO2 3,&d0u<%
/*JN|<|8Oi_WA\U@Qe_RS*txw7iR+4U^&Sd*[_;^{G? 
bVM1I?o&W_L7'ejGokW])E,3R
wkfUw%&NnN=NX|p10<:%G(6CR3}CmMOTDw#X)[Ql?
CE~\K3Jy9u*)Ky&'RKUi=!(h?Lc(!Te{f}J(#<@USVYrNq5w,ZQJchs4)al]VS i>]:))/47ns[69j<}9Es^V0ShX%L'SAI!gxEn8*h?vA|6jku.HUPd]}cHe4}?V7	 :.`W~3I|l?}w='x,\a#7|yhJuM4Bo@;hJO-50N#|kvyq2g-K6uYID,Fd?R4VsYu*'`Lv5pRIHZu8?Tpv5RZI=>6f>I>O@>~{2x=jG(- Z)M6f3ee_70%opvlqEy#2\r[3~#:][LxjA rK)}/2_P"d6H*v@hxdMPjeqkzmwI^,$kdRj[H-AWU:x7=A,ZKF	?r=t/T=Q7~99WK(6e0yo*Xm}@Y;6}Q/RKd}*[|y,Z@6ZE#k63'V$4hu<[r<6K_':zC^o%yXWohPXK"x]R?EcTn	pN49R]u5[J`ue'ms2T[SSjFij\zKP(I.NDzdXD2b583;+dNK9}kQ61
LaB!/	#zD0bLd[q!^,t|$ou^T7}D=a[?'6`qJ
=N41Au;)NR7e|?qbFgle~V+&g):Wxp,W8%s/SI4Y;iO!Gn
	ZkDedcTV|;wK 7};cb`!bJ(a`u5pS1CRYonZ"dt{MH4T6Zw&)`7`
5UG0U]0#'#5AWimb4m,uYDKOocBF1@kszd#iP/R*H4-ZL7_`?E7}C}ixf,sUWjNfCSD%3-
JjVZlY9o2"X8YVb%n&-eBfoNeR!cx3L}xBA;Y
hk-nkV:(8>qhwKZXxGZxE4]}(8	st;UA6X:ZZF?<A:x]H;kiT;3g7modreenAuY{x*S{N]8[,K%FkfNlbz<s>8d`* WK0,yxt+~bO<c[?QRo](bLn>W9V<T!-)K{(c7ZA#0M YHh"K`W<Tvy!H1a}`EDC
yZ:$5V=" V[IXJ6\jC=5ZMLIQ'eX_@]!|oX<Q.8@7i{YGzm*d@@$W}L.Ft);/DhwXu\O?kmRVtuW/V(7TgA88\[>G!A/-#8Hv(oEA[?!c*%2TD]*y!K71x)Z>y3
NE@RCG7)_g`T36r6)oJ]#!fq77n>gV\(yFn_e!]LC^cY2kBh5L1fp]Eu;2Qn%/mkgWc6*_M@oe`,KP`a''!NBgTTGwN(-d7>nU9	lo..N9lZs:t]<Q!9L\;oB,Y7G@	M1kts}H	crt[D~<y\D?5O~TNx95W/tpXMdWcT>&V&'.[^[;Qsa$q4oDlkzTy}T*8n,E^Tx!m/Gy9z
-$mxp0P`U|6N3'C4*%ui0Pnsqz{lD[:%vz!8l[Fl~f9*s56*:)<KVs4gno~)M6~ho?l%Lan"`R1zi#3G32&o$;JV\nB+W61WC$vj	&U2/INP(-wV@"53pcMst>'O	
 |G1d>#}:|=PQ(Yb-4<odSQj}T,-apxS<1;,},]>u> ;*Yb~cm%dzCs&#754672S%E6A	LugL=#dh\%|98?Adn.)ZqvXigd:<#SVMnp_PHoV	v)|O\{uJ
s_7nO=jy+3Pnz!|}%1BP*x&M/:A6+"@1%6as"fM^Me`I9C\eyIy64HL6]re86fMem&Zm=L[#5vBrGuKg%&GQ|0Z@oPz!wik/_~^sc<Ek9~:$\)dVcmpVlk#g[^->/q#R)PNv"vKu2\:po'QPZ@j=1OQhE/
+rJYcG=0h4yGoZ9\ o=SH/lkhQsK=Zyvj\qfy&/XKz.ai~E@a,jC1XxP*	h3S8xfM)cFg){Of|:!|7PC/Rncl~lahJkOGMOY6`ZK|_gSL'[<\wm#*
}>a&_i&NW()<$Mb	8|ULSB	K){Lb0Y&tz,9)"mqJ/M"I7{f&2/7(yZGsMJ{\1l(~
!e4`}Rs`j6i9YTI5~i7MK|<3"3m4!hcT@]PE1VO33:(^szdEE3su|9ozZ{Z)]GtB`Z:-fRp%!aW<wGju-7wV{+kM4Wa9D/F1LPvB:
ty_6~<&JId_"5)7%`^|UK	s[MgLdIUoaHm#W$@?)Pbz~aQ:6z0)7FmYY"tJ'6dR"=70l+t<!|KoERB&ul?"uXX"@LylFk)uq5DBy:`</6#
(4P,hE:OqpW61V|Kd|R"?W-}/:H'fl ML:HdM:>9NvPnLrS).VWsjyk@5ScHLmGe;n4)Lp/.:dJ5ThT%n^<KHo htuw`$G127f]1y-7q`k=:BTO)v/gW'\awE]OSL4snQp40<y!}"\pF^lL;oz#[VZv*{[pIP`VWcXnH\(PvCw3_:Wp{(H	l\-vchBtyb!Y>.]Usb-<Q5Bk]+n>dc\/u1F#h]wV!CQ?/QfB:V9DQl_d}6$BwY-aRt_RyC<DQu)yN
Q&qRP[<0%f"d0`<W,O9wfZ]4>va$*b)'..2|\4T+p}lfm}w,m~i2]9:pFk`z!0%|w7,z[\]Axlu)1Om#[o6#A=YnKy~;@
Ojh16Uuqfu7-	iF}(Ws<e/pe0<aOUm*l[,%[f8?Jk:RX`Ei`:=[')lICV/f/~GXnVld6!MI+g-m\Zhv BR]o|<P#}S&SG[ &Z=@@4fw\c1Xv*Gu?om5	,uxtI)KfAf;{D2L/4Qs FjkhU(Ky^Z>GTnRhsS7S=WQk=wm$63u{/fH&snK_+D*CQrC+6j}#^dbX*-vh5r{qG,XhsfWk L{??hoq^]XACHzy!';Z'>bhQ<f"ef6TTnKG9`Wa{)vo	RXNGBumO\[YJ/!u	rL-wK)T'C_;l<hGL:s0ib,/y`i%:sg4r~Kc<6]w>^tR.	:ucKNuVy[DQD5wzn QE4.N&nc.;k8L;x]@zdJ5:Qs@`T0d?]ICdj#93&1n@$<Zz7=%)xr]}	nQiM[)H2!1f8L~$,KmN*v0A{A@@]M9mur9?1U}5vf8.aZ\wb+T|Uy
_hD"`[AE
s}67C8np4k(|R>A4-DD=:oPQ_[>"KH1dLHJ%2cN,0<h+%{ *{0)ih]K[	1*{(Uv
hb`#Zd~]T.j\aV[3&wjMf2+m9%|w.ZrT6O?g
a>;T>pf[)gMni8KhU.O
d_sd2Kem NMh_(ATc,_(vXivIWP)B\AC>pjnoE~wp!9zmku@[k"AG(JaGiB_y"bU\P(k>?[QVl+rq69X	_"]3$fihE4CgVz:he/6{J7Ag
f[gcB2m'>@1yR=j8[#}s).uqg}F'78+?%Ah;I#pJ:	5~>dBKT+R5CqO}sKE['IRcF7?=V,Ohj( M&^i|)/f:3'@EK6*9mu``aJ~F,Rs77dK8X6vG1
m~A)Gw2$'Y^>	.1;aDS (v152[=/%9*S'hLE!{Oc@p>\iiQ'qcFw#zv.<a5&)zsjaph{l$!XV,8o24Id,D)eU5{-TcD?A
ho|_q0[W&P}CVXm v/R%\s(l>W_u>q=!D(bw
}8]xQqR-Byy)gc2>2^oF2w+DU2?Yi3\n.72>8gvx5Hq17/b=HRY3}<vKy^!J.4AeBD$>3xVRgzoI>%w2]K{hcy1Tkx"y#*lYcKFp(MjC]VH\f]	a?m'RN:`>[Fr"@0#17)gA8 TujX~UERXh/Y"!\qB*^1P /3uNydIcCUhh~~"P`ls##kDj-iNnKDL/uL;sEC-LuB\_W/Cj{1n=C^@\m0SZR{s5"y=Xl$5r}'[0gD!dAEc?*Z
nFR\^]/<vs}?P
4(?AKPGCH=U6O<5~2<!gWwPf:{hr/?UAyQ:-fd{b[}yj~";#PXH4e)gfE"|iHq{w#N43NyvfwY.[LwYByL{54""P?,w&GtH*ph7,Jx( 4KQesOXnr)]$yaS7n?]WW?|*^tDFz%2=)i#mRI^C'q<,blU?B|EQ`lx#Aa|\2&'U[Px8kx!/D/ZL^^
g69f@[\pp:1i*+L2_YAy&:>@b#K}+p7:?#'9V`wC~,X'LPG*YZCra"'=t	sF<iCP){<	Jkp|3'o]-Q;{ce..k!1U!Vuw=su@tLM^epP0S PhgK	X~\^T@1}^'OW2t6kWqU"NKWoCUp/xk lh+[VNgv,1uB4%=hDu?_I,fw$3W$`)@hJ,rQNjwX)ihNI-O>C[==@jt&jot[Kpw
rM+$iNPU:9^<yQF_6k*r17Le~P(A_d{;!JiD/U_ *%5qdE}l-B6a%1&h[PSY7qUqOU*}{([I=J:o?7BBoHn<[)e)I5BR~/#OVQJ8l@:8l,'!D*Hh#	nttzUbzxJ7wHTm,S_M#W.k,EFEUFOTR
b ,?BsX+F;}Ot9(QWB%IIu&o.@B
RB:_`Gdr>\n\@tk86j_jlQ%^hwaMmvLaFUNX(eo& q V#L{Dhv{9GQ]LE/^\4uSk-$A|W!|EUc7kFQwLvmS0'B	yAi5>cBv7h\v1'9QqhA7(	{Zx&"3y9eHn:>J%)RNd
VD;44z-t_3/p!x_OZ;^]g/iB6ieS1$	vI:fd)%UhQ4%T.qoCxTvM5a
Qh.C|F|.$|gtl^UBhLC!I!r$ 	{DS*DHBD|Zin<$[|OIGTq49L2B/Mp=A99'DzrQqQ=Wo"V<W6A^VlpMj4R^ Y!AUN&3#pNzb=U2a}Z(*KecqVrOvdL0q[uI#^)wDKLQi.rg7g3!5j27X%>Ru[YbK{qCB9?9)V@$zb<w^ceKQX{x$($VOd2Iq+7z;` Odj|`MAEh^D1p<L;^M3AH&st[A<W!qPy]w8EMl$R;J]N'fnFOFq8J8OyGa;Nw@4tP{:zug	\hH@y6t0PWVSL%/PJV3hd4CKwxvEJpd.k~eYjck'6ia{Gw>%ds}e;"KAD%P0e	ho`	o![,u<E,9's_:lK/J<9h8}x%G[o'=pxpA=S5|"3BH;@S3E
<3'/0C\SGn.n1Gc:{a'crv(8SE*>Bh\"ST8f]s)&j\(
j=d/ueZ2@w2J5B.KJYp
rq"(5eeUziw\=$zzED%yV'pl xU0H6MHh#_c%O	3pVFZGq6L~$g@z7i*:AzdUR:\Ph>y<5NZ:Y^GIx]+[)k78Qiu	v-pD cJ`~ss&0Asnk3~Z|:.ff}XWAp@SLP2$#QWJQza\7=(
F{,Z>tYX4A{cL't)H,a	<>qwt1C!k~U	NK,d4O>iOl>JY7RE.Liam6UEV0Unlw,{q<JAXNg*p#VknJ-	@\f@ZB./><[m>W\7Oe=Rzd'?\&9x`[B^f}+n
z8C7<h?}zqy)iF1'#5U.>deAYqM7#q)JO}TS5qXD#=k-FM,{P%Y_{3 Ok*@V:In$}R(	ZTA0S0.Fj{_Mp7wkkizDqT<Ugv\]H9=jM02O>ql`4L@X)g_(dm[OE8W0}Rk2*|SjvBTNu%ET{.3TWf50,Jg`~s@{4|tZQPe/E{~$Ha=+c>!8K-;*Cy)t!0w{vg\|=2Ao$_r
gkwgvYC5xakvb#f:P6E/HRGa$8G:v:9]O<dK?~GXm!7<n;0{(\.'LK\x%umoWh91&B|8
*@i8Cvhi8Ua\\|u<COsB{RD~CTBJ61^|K*,B^^D{8gV"	txmo#R7Gg	1Lt>Dkn$"3zI1 HfB	R4soS;e\i&	*8?l!Q=m9q8m:~v]@:>RZn{RfHbr{k
&Wy(d.<sQxDDf4mwf53ka/)kZo=KSDs)41,]Ln'{EcyQ/ALC%np)Bl5N8s\qXNphYF=yNA<:[xd7qH-Pp!(KR(V0S(t["o!hdhR(AH)E8>'/U\{g'y .RdS)y>ctmbz*Rjd2La<`@V[SBQ
 YDntA`Ff;|s_r*<j(/].0s-*E>#K=Ub2>dKSR4UnM'Az47:jmM_b>X:3Ptc4QnC56`M9(2G'C j\%"ky+^e:.Y%4YK=OTi&TQ-)^=6S+i^}}&;EFR(?e4<Vj,I#jq	/c%BX8ADC>K:W-&KP-zi5zAZ~97#Ed`+
srWDay6xKU0'u;:,zmr)*y+wgwE.p6dP8bZj(*t.UjM\o0Enhzw@$DH-{FA*Sf\+u[FcZlfQ Vx 0|J4Qi.F)h&<km5Xyp+|`;!Te_pX#NZ<-U-mKm{5ChcI|'ql*3H3mLfQPO"~Q:A89
'\+-gG*qsw4O^Us	=AY'7bU%m<"Wvl'-vF=R5:*nDb}rB]p,h}"z^?3
m!%)bV^mc=8uqn^p%uPNjr?Ij@bIWAsBzf*BCbq,\A""C"uP/AYZvzprcEK7e_O<?@urv[bmt	IOtq(W'w6pK`Q$A)riL9=(R
iW_+!?2TiPN0vmRw-\Q1*<Q0Erfmbz)>kwIDI0q(@^Q9v-VcRmtBF3X4
rPklQ~,m1oW9)'jLt
yM{(u!$Uas
]9ERLql6AIMZ$^ C'Yo7.f\
"J?Yyk=3S4bU5,@ziy*3$33u
r!cK,((d`pSx/r-q8xz_{~08Kn%=WbzlF*0^Qs\~SGam\gB?!cnGZ9F@!yQ\spmf;2oI{xA}]2ZDq&w107;wME"g{s|pSa-6&?ep6U0L<J>sX	TL(*r|^)_{Vzh a CqY7tNMu',v?~+Cz hj`k^?U>7T-yUNnP|x)_46)@rbH)Y$Vr-OT7f`9Q3i8#F3`\&#qI!3 d>c  -A%dBvD[eEr54V}Yo+u5_{=^g?zWL_1{:AVUZ\$R=tPKS9s-Tgs
0S0o2|NW~vbh*n?nSiLOB1/dxNad ^?.8+YY'DkO_FGx(1+m|p55vGH,JX"A,I#<4U-({odqJt35|_9$EzFFcR sU3~4m<y+q*MUCdX{]$uopzDg
z`=pO9}=>_4-k('Im_Eo{Mc\5q'^FoBR!Y47'}3|\J ,}6iBBGe-.t[X2194{EkaK*+$YOJ6Fl\dG0k}K2,L|pU0&rB}c8M`Zjn\1@,SG]_HaoCC,oG3pVGKHJ3Luos;G
J"+A-Gj,b*	_/H)VPC/^6d(B7oU_&KyTABxb>ZVLh@/.!!z46lsr${sb"*~8mZH~j~2mvdpu~Hh{-NHR|#iXV-|-'I"I.}TDW{zUAol#;c6k+^$^2!VP[J-k+Ml*s`VP}PKPDW'm@eoDv;om.luOTfP%=s:7%(T0dD<*m-&9csf.l>qLm>~k.E(j(;rEPU\s=$7#@J
[`GIXV>[_WGWW)ia]iW5F~<M)e*iZX6RViqLRl5hn[<(m.F]Pp8e%Z)twl
Sz:9yeyPMI3	K)!(b{F%s-?Gnd(`H	0v|Y|]	}/z:'8QqeXwO6XX
qSJispWo"D[<g`}gMf6%wX`!_4F:Y])."TEP%nRTaX4}>(ZctH!zP^lb+!s}wPZKe*i,O@mrE$VegM#FM4MD8P-n./9&W9[_=IRbL7^sFp T}R.M@C&Z!i32%T+wHkuEtCgvXb>f~dxW0sT+yx48gl2pcg{#7-.qEvrsX(uvVf)@`;F|(i";B}Fz&z/w>d)'SUT2WJn>L-u8J,xKw+5F{^5e9m:].p|~$+<i /p'o=f4oBeipN0	<02akNJml08(n]N]!J1	,D)$4!\ u7Dg>bL">a!YQEq+jUyJj	V/]ofO;utTeP"bH`)Pn*T29q&6R>`:6&z,'0uC^6x$ .|r'.C)R#|[:^#kKZn4K)q Sx *(~szCw3q8@YA\+G[`>QPG^loiz&.R}LZ|w2oY,<t~%]V_CxwpPtEXLa!`I6UTBp[q-%HztryyUzMh<G,}rIOAj~
oaC_vQKrT03CL{}<s
!hs}nh}83Y<E 5=li%+}`J	!sY7e\Sypi$W1q.J2n9M>M=EQS`bbVVa8z`/XN+n]BxgPb8!!xuVG|Ey8`.|L$TO1w`'_l jD5:h4?sN7R,]o^+[+nH}iLW4R$r}:71v^VOXDjtE^/ce|7T1hU!6qb^47G_?Rn3gM,WrHF~|H8*Y;WQv1prxH=ltIu#/E~sI=Ir~kKxo+
da1
oXtKE`cM/6j95g1$VSSr#Ph'
-@2-	9/P:(Rr6oqm:ky	(7\T0`V1vFc&s0CqT+'hoF3Z~oas0Vqievgq+_e:5\MC/Pg$Z,Q/JDS-.3`H}Gw7#DfJs>^<>J0:0\Zy:o4 nX9V),Zs!P,bM'uPA$Fj}=veBi%\"?^*;V,@d(wm%*8>dk$#+mnL4la-C-Pbw%"{MJd9ZVZV'*g:MQRZ&T48N|8."$Z&>J/; P;P(>7Di8)yq{6Pw_jo0H1K">z8X4I4J+w<049'7oRc	BS%AyA1$Yz[JKV[]0Fe&]e.g4&hlI..wI7v;Cb_HK:'>-xm82J,+3Oa-yy#K2#}CG5@_55qp8\s0Eu0Gc"H%C,0</*3;VP}}fAc>unF?O^M42OA'2_uf(A4$Oc0=X$
jRc'hH3E[}_KKsUZMrt`@k$ky*T;y	m1@ct7b_tfx1_I:Ktm
|D|b\L2,^y~AguTO7%xJWec2lF>~T%ehrPn	K=z$]G@p)7p[,4~Ob.'nsuCkL4OV=v4bSY
Fg=<BjfyWL{qLC?nxRhRD!"@0)v.COxVh(}`EP~d?#K>=^W6>u2~XCk&IJr6>gx<agc1z&yi47FT}4.U:,1uy5/25NGrE`gr+%u=/D,PYEB7{L3T=,&G<
>MV^!JgS -@*-7pAWW3P3X`Ywl} $vFO/K8-H	3rZy+U5:QaYjJb$}	lJwwV>&,j!]g
Sx7W@lIu[K4pa\j0lu4E'\B=XcGAv$ff~R?/k"CAJxyr (/$5|)8wD6@h!l[dH	!k+OHlViE}llb'@SBjKPzz=~KW/rVx.Jf>9dQp4nwrR<^gu.(^HVwy?6j8*@C!'j:/ imdmPbO"qLPKg;zr/6X0n<(3iWIZlPUF6uc< cL(|U=4O|/,E&={A@lp;-/?+AF4RoPCz0Q j1{W^p*{aa!h'tzDbYi.KKx_ [DAK#G1aa)&|Gs}w__VB`Tn
#2X#P1o`Mb	W&$DqE9\KCpm}~qs)?NJ 5v4fW>R
01}eH} tvc,;5umI18t4?TbbvV35ED<-lX.UK0Orp(3QK\SQ'9omWRzB!J^pP@nQ#BF5<J)&_+)fxo',m|Sb;d_v@<,tx$Q#sf{?C^FYm.+3[6y7QIB]so"u5UP?@$@J	6$=^s*d?b>OG5@[0qRFPxJ2`v"?K[4wnY/2w6mRH o[agS/L90X7E^4YvbiulX)N4R_$BSz_a~&ZypN4NlVZL3	'O *gY61kK+|6J{QQ:hX$ku`wbhBdf8L3Gc5P,-ZT<{]M=.^o?At'b	z8xliPup,xg0@V=M(uIG6F-eZ+~8cg1g"|xR_vfH+
O$N+T$
PL,@Jvl\69S/_N$Nzhz&L-xr@3("Xr9ZH.Zl#;*.`n.
{B+O)yp$oqifyq/:^&Z;w?4S^)cg5C4%peVr?EFwS*@7<+,}pX4h7 >.[3V$^CALV;r,H{o.Ie@aoJp?xJ/+21HN*& NE> L8'_)Zt)a|I?-^\-53iN b064j)wP5RMoT[w+68j4r	d]&]`	6u+Za
BTSry^0hY8?N'177D."b`#pPW Nh!q3.0dq:Q=-B\8"&wP4,H~hE1Edo!oldWh[l8U9'b;C)/A_cAw0J6H.v@Y'>DNOoEEVv, 6lm^%^serD%X2o;q
0x'G>dp}$`ptQ/-2Y(XBFV{.FbbA"k!tql
P}
1}6>\+56uyc!|}vbmx\}nCL9mE5jtvff-J B2j&k$(7>;w#xJQH4~!]}y<Hpbk/^=pb_)eZ`F:^dDKhiFxWEKY:O4Ew^&\#L6k]nx&`(D2Rkv>s=QD={>M?d[L:n*c|onNM[=MFs[6]!sE-%Ci~N]-jv#a8pRu*AiA(#ZvSprWHhItXW*v-@*sc,Bfo-$HT wL,$'dujGyYN[C(h ~k]F0P}^9&=-)I(xvF;
cu
kkY[#|f|WNia3T^jgbn=lMW~?}lc*Bi~X	t5eCT+i9BIynqMBcO-*y`-3i8gM[9{Nsp,\&a[C{KnVbX`CI^ki^N6jY$J_/}t"n~JA["yoKlSrl!?pRh$\L1&'V@+v]#,x-ns!G[BM3/)	~Vp29H'[m/,K)nW"LpEfCTi|b6a:b3VHkN6t^g{IHnT/I5iK	#6
sC4#^GvF>[,iD'nvp1fx]/@LcNm|s~0d %][}D<1f^cF.uA"oxh=*mFIJ@3,nS)%{g<#C^}m,t_%M B_*-nZDG30Q$U|XKF9#e!z854Gp-<6z*K[n,IL h~s2}}OS8<1\okMH|2CDkz:[C+:lT/>GB]~<d1/::nrm[oN{Zzs}>G9x">\]y$\}aWK+v20-(]nQD(,rpR5dU]"(JjoE[J;R5h5r}:*?l68Jn,~#A4}dH<?s
c5v 	w6|`^[",#VN%DB&2]mFriyi,cF'v?fs`QT^eI	M~,f0._p:!(roI+)~EHKU	zZegt^29C)TRu6Od`'s&}1YTkg+$/<~|#
4(t.<~AgH_E;cqKd	KX1O6aX[YR\$*^kWhi,,{?P@=m?aMe*(J&9ZHVTch_}2W
LQSZkwGQ<omLX~9Y-f2]:JWYD%`V"pEp3P}	y;{}PAjcT5nb{c!;DOPp,zD/
]"jgOMyBvIcD	+0:o65`_AFk-eOY}_ll4B?]nq&-mH&-$Tm:!DSFGW:seF#8ci4iM|JC8`;BQ: pREBop$hn#L<ue&10>MU3BJp@6[FqYT*M2(L9!zEn0#S\1#tf[j!>fG=d+	+BvZti`b4:]?dW"
>=K#oeot|m1(k,=eE&1[}E}FY3T9^d%^/Q5$3hWgppzAlCf`V*QR|	d't9rYT7U,I<	qp*2*p|Yl|]>u1[Q%8<!5<5{PC52qWA6t.LKWk\s70K(hF-%^pV""8V_^0I_
Ba[hAc:~)yF|b&uxG)wtc2Fxd}|0Og_{X4l=*K	EX]1'j4\Q	~5!rYQ@cxZdfEIBCr!"TudYs	QoreC.!1=2wtkD~R[[XYEw#$:(r>`k{"-VPqR:nJ#g,(Pzr.yB*,HI #mg2d[qQD[*6C{K/BjG.2/@aB@Zg)3/@0xDX8[lFZ34"a')a;/hec=vTm%J|XIUeU8VUkCQY?"Q&E-H?\&|-g1Zsc/Lv @D(bGKITWa|*8m*>'sI1fb7rW)xW=h1rJST\2|jio$nLDhn\Hk
D*OjVHPxu2/P9\s5RcXBG]e};xqC0?[l2f	!yo:s,/{wPZ;K\ $='[[haN,(|#'7DlI_9MYv( $}Ej@DUU^=PP#TH7UgX,}5]`B+3[m/4yj:u^;J=3FFA|@>d9AzQxLN6
$P pQcR;dx^D|CrT;#Pvf#5	,`l
Zk}4Zxjh*&N0Vm\8i!xKw19IVB9._lP$X-9&pphP+55eS)+SeMnV`^I[qn<Nt&$kuCO?x'9&2kg Y%Sr]&n	rPgLG180G\Fs.N%]"I{.%O ?]3*7<NA5hCUN[MDvX6WVysuQjCO:k
S50k<77]g"wC5fq0'a$~Z9nMK>BxF(jvihbT/\n_ ?g(IGr6_bny_`	&G==O0xD>Pz"m$Aht%?+f(|0XPu{Rwo",<3(~\9u5Y`wg2-k5<qky.P+W)9X{JD.;pyO`!04w6bM'D`MiRR*|6e*;D[.dL=..3xi}xlE`K)=5e6(AM*_XW#E/^}-u$doyA-Z\x_F:sAX3Bq!@e^Oge(L\HhoR+Lu8?Lalh%S1zTxqs7uTk<gHDeSXA6PSq7i'\k\9}3ckBy]@`mz;1(u==WqP%d+91[@Je#,<%%]3y!Eds(2D:SzAmN3:L	}i`2Ku$0JqCgI	,ZG-Zk1vW kxs2rm0gV$NOo0S=D&xKfdB)j{n){3IUu>*egP{cDz?/OBeHoNk74\;M8},qmF$g@~*.'@BHwU*CxmyWa)/E0#wXwetNL`O}`'"[hxi4FH)f--s&'	0hw{3R$UG"`UuNz6?NB#tVgGh1t?h`dO-wn`BX-9U=5jR?6yV$F!/.+YP&_G*>Y`+x@r@q~dNF4acP	Pq	!\(5-/y<o2^UnO?VR1z(I2zAx]aGVh0H?EiSf&X,t	8E(XATajTOE`]_)^D8"9\n!KU#CE5``B[wIu,MH-Mn&hD+LVToK8)DBcLQ_K!X<*$`T*6o<'5\9|+/#t<5-,JZS

t;rjF@V_4}\n6Ax%"wS0azkTF8h.c+v@/2rK1zhKU
-:,{9O=@a#aPxF{Qt
0gD@E;0QO>zre4
_DzP6C9x07[=bm1	0A*0uac0?C|CdY6I,xc*5,>y.?sqUX`[UI<%lI
Qu[>SG8+b|x^7znY&$Vbz!dcK]D}c^U/V@'t{,F=gR,S(?c[F<og[#tgN%k/>Q%(I5w%Ud<4h"7#
B<y|^,?^i.lb4M*RtbKPPE;(|tW	[yr/%7%YRR5'TPS\!<JZ+Ee+pCS?z4/1:"{]*{q2m>G7nKkQ!>@D8Q>QBp'/(PwFc%=jiE4L3`W#,35z;b8eaKk(]X+b?>'CB=}Z9]8:`a bO
3.wR=~~r~>!z)oJw#yIJ+xHx+nR5S1<$@;Ac$4wNY(AWi:}J
wf$y]H_suYc,`z=aaTgExdtTF5]qjN\d@&eNXS58nwbsk4AM ,!,U6FA$,MN9ua
yfTfDK+Tn=&S%rxqJw~)xmM.1m?2`Pq1eRTDd[lJ}#Oq,q@'H?dwkHMJNr9_U(D|$>^sgBl )w~{"O~$z,ag!k|;.pBPNBv"n$`^"kO2{oo/u_VN`.ITI#	X&<T`3\_<k3UvbA\rQqxuP;71J=/_YEWA]t!jw.Vs3!Cg\J	S@9ky[0r=fEkM7N[h-T`B8t%m>v?lsOI	4nXjU#hQ}"Ej}`TLX|j4^b?W`<*lTG%C'bI9{'N]IPhXA.rvW+1xRt?>	YorlSc>Yc~90\)iUTR{w'?6d.Sw"k {J>#,8,oM?m'b4f@%N6p/n1mg@.|~T+;m)U/i^`qY#s2{6-B`(_GuTE[<!9OH@Mgp?mYxn$hItM^.Pl'(afJ7t<$W<LW=,h={E!da^p/|m
37u
sUt%v7SQ2;Uk=2$kQ!|/o.CA	M+(W Y'&JCA_4j	s+}x I22.PNt!OxbB9,	x5"/~jtK) ObAl;+s,GrH!">h}Qk&
.? yh`;2d2cm$0IZ% ?y-Z`CsXX 1WIkl)Y*Ez>[K$oj+ne|mO7msMGj`!HZH+XuR\[?R@2!*9mTM!2WE]K#|-OB12>iJ/Jp?\/*Gnus;ycQ[zJx9rd{k=},[W8:f"LFi'Nl%4\	|OkIz)rWlN=|v0 9\i%6pHXOd/S*z"/CVQf(=4:C}Q%-en{
<!m[?'N/z:JHbU#\WmYH	>Qi'sqx@Pp[),s7IOgR"	_=ixHBH3rUQ1U\	J$s2Z92TF*;lV7IZ1Vg4t;qeO h;"stI`9;Ve*3rOJ>lwCb|u_)k.5"RsX/IH6A<67!dVs1lz{KQz_?0,4nCQQ/)LS TJj~~`[6bhP2&6=oinm~TXU>Di9+E{h'6\Gf_R>HqxR@`r07hlC];KN~r9G{\oDvRy5L`S vF<vrj-=K>_o|`S,QfYogfe)?Ecwc6%eDt6yl*Qsv3q)s>zb7X{rnk*'%7&\CY2F]GPF6v!RqCD"`P84U\6XB?#Z) Wg9aM m"2Qd8Q&895(e~$qXz|JfH<[g^H`c(1?6jyjK(!iV+TOi
{'R%-R]Fv9,v0}[YgtP63F'z0yX,9Bsaq42gQ%,=Q*><wSMR&
]i_,QjZ|ND}o#k#	9sl/w}k9UdMGK|u<BoK!Eqg9'+D|{E\+4H)[Wwk@sK{16KBTLY?Dh)=:a*@~K{`<+#adwN'j;Cv_N@aoIk=Mz;'K}_V)ACoP:@BN?h>K j}"]^%H+y;bv|unG'}dQiVvC.SEJST#X9`^2/eR%c[p!a$s^tI2Y4Kn(onBk<.{DkA!#D&aDV~^OEjiP3Xa63-S#P'wPO%ZO,q{/Z{UpXNr/DdW>eWFr0T;flM\B@+"g=\rjB>=@e w[avq~"'Sx;a5<o	9zLwR9%pD
W +xupF-jD#Q)2nfb:	Cxux2
sUDU|CDZy9{oR^(DuHu;$(OZy|;er!PO9`_6Z"tMU,JIkY|=C`n"aZL( 6`m!H.|QftqUO+upi=0T0gz"u~17B)oY%=`mVs'J1a<BV!W4F?U9OK|OAA+
ia"\F`jWey'36vq7'5l)Wt@Ok\~p2$Tlht;^0PBTzb!uuDNc*`pkbRg"b&E%-P2<#*=KA#6<FF	g59	tI#=`.:Y.5^@Na;?=<Cf	&~k-&;Un:m+y*O(~Ph"&==x2V;5kwx+x|0w0>${m~g['a	+CumlsFn:*/7&WB`[!scgAh77Z*f%sHFl"\:{~c4?31Mpv%B.w%_p
+T\dJBF^X]8P/b;2P.AJ#8+QvT<#!j.9qbUk_+mS MibmwH/GoNE#3!M{\JO3]po)?aGeu2x^1U,/zpM&<+fjY:>`X",OH)9pcZA9ED'?1B"$K>7iRI=?CK)y47OlXf$pdD`nk!dSA	
p_@+Jcd lE_qK}G+-n1Ny.!!Nq]Dv	]*=QZ;N/HbzJtHIlu6vmFq>#n%]H'?psAg	EK@;lr|]~ Pd2D0q?#c2_Sp-*T+dUwm24'GHE8wMhRWiq1T=|"0937JKT7.)?`t@jjeOsUGm.???-:"KmJz=H1OfV;TvKy0xP=l$5V5q]@x`,(J[!uqKG'nf8qo%.mZ/C!IY%M\!SSVG,AUd`;\9s*~8yc0{jPL;2#wmNa; 8MUu+*$j79H?^e6-&K<UW"ZRG6\
,2"y(~=t_I/kJyT:.vI7<;.mMKM-}),ii
2YG$5K@OhH~^;|?WW{=+70#')+jlP|fWQI66l&\nsH-+bk{+)N810;" i*bo(eY(k.`
A2L$y:Ti[ Vu@j{i9`)k8++746!U%vAu6K5T."	3r~Tmx)@\gGRlRaVVCd}s9t0!v#YWv,*+|R,PO]Y?U/Vh;q.Mg\T$IO+0o$>&hY^R/6,u8@|0{;]B3A_>
tX"|o1,ll[t^=W(-Z&h%+rc'%?#x,NK5HHoaO2|TqoMC?on{D`v	#GM[\[>H-6}#+X9	1>pwr^ \AT)f)-&k=G_b-7Dz+%N>YR#SK=5697>b"Y/E2']s='VH)M\?LztCQO>oNn\7V3!aAyFJX?J((boli.n}Zq/fu,vkj5`orcJ,A~Dh?1txHX$|~<(YN&@ 7,J7x,ma2Nvpc:A,-M]aki<Ypm^$dJt>M:?SK3\lT 	XT;0NA>L`X\SWA>M2]A.H3NI5+1xL>~OVly(`v:Q*2p(vTMRB*gU9h1N"NQ:	WklDWyC%@d2&AE
^&IFXmc_Hi}}zVhe[a.0WmUV<E1}WF}==$goE:+,9{5sq6C	8MSA%snR>{))l]$x.7P]j^BXa1{:#!sle QPTf+.7sWM*W'et#P6dgGbn/K@GZ2IQ8%%S&hYmbR[_QK7>+Y!\7U^fWk*!g@MRN~IlxF1L5Ss!
T&-hzyc&ttB6fPg=<XCq4}iMxKwN`pV	6nLX.BPUIOz.Zyevpxf}/y8c1`2yP12j+omiva~#m}F=h%>(<1e[xw yM6)Q8E%!;_<!ka0&Z3\pI8Qp<&VIkne\v4@]_m@# 6,	&474ge;.WN)in9:onCOmYQJ{= ,uU~Vd@|FNUK2F4([} -ugLmI6RQm+7$	)&bNOd&RPJ}JT<#;O>>qbu0)i=0UMy?AByt)ci})d'(J-VNOqQFQw#0xo)m4x"<_u;^9|y-8&f1R3{P-\;f=x<n(XulC[TZ58	"tQA.1r&{yN:mju0e-&Bfy.-
g*KE~*so26QA@7a7H*i!rv;e2(4{3>PA"-@!rb0Xfk29J/QGS$ptGw IHh5XkdfDwS!o=Bm0x}&i*W\uMsG}HXsrMa `6I](4.;Jfz^%&a`88H$KFuTqN>@Y$!z>^nj[qWks&
K8zyt]n0w0J \6Ko9!fGN]{#8zI~Z#>zfbgoSJ*u"aYuh#[RI(%[y/XPAJ?Ck`+P-woAv/NqL>0
;2li5	Ay(l;k?Vwa)^iJeD%txZ6$M*0NY4|&f&KOJijIsrn=7 K{v0
0Km]
C~h'M]!dCG]D|Tps6I+G{?9|dK	)' `;uYuO_`d?'}:*b0Zbf)/oR/LC9\=&;hL\T12v-0eNwrBGX0^)F3}X''s)_u>pxw]-x[]N!?qMpt\<DENYG\:<q`AvfT/1f1R`hc)tep[YO-c"f$ TR"6ZAQkQ	)lTnO7S)`'j<U&krb_9B)mB/r!Ha?%rSB3tZ{GK[dZO- zV7)xbZ2+Yr4.3~IsH.:bY3nA+f0\>CH]O `|5C5
pH&dWW%vxPuc:9"NMRgY".$etn-H{w4cy]KW< #<i'ZJZjly2#GB/!w6/<:'B\eK'N~B<A#VC'FR,-7oZ|A3)RdVIf'@Vhwp^IXqQuas7td|Hn?Bwu>`[)^$I`&ix3v)u|vZvMU].gK9Cq4\#\bWT* #NlG;7Qm""\v}v9W.R1[@ZcXO	+r)S9S{>zI8}?3yx/TdPr#t?SYJb; h_1}{[zzCCFOP$Ua,%HMNrEq'}c&Q41$]`_t8Gk-(t1e@xdq)<2!4A12#I	eKA^jyRKERS\0W%"C@CdSVIrr8I`vW:$b$3mkvp @!TI+007cGx@#abu?-.aPeK	<{QG<XQjK0:\LWM7PEOlD,QK&o!M;/"+"l+N^B,?2{S(!3hq.SA+]IHa:b6(8NXXQYdGLr2To*krKTA{j0<^#?YU*QqbKw5@]7?1\yL((0nRnm[Zv8+zBu}a@1e;2i)G L4J|f^r$nLn96|[(09<:G?u#m5ytVu/U1s&:Q4He45ke(2}*D}K&eZ\qRQ	<)>6nkD{9f\uwk_y7U}-
x%zW@]F\"S-nq\E<u6a*RanGF%~unI|	G>.K,Z^Q\BCBWWjt 2*:CtRs'{>h}h'YDHg2%}W51/6tR.d980k*VtkgpFP66iiU^_2huN6	.O0f.4<>.uN;12m
p~06ur
W@0N5~#%OF'o
6]Z%IpbC{c&(O]Wy-<{mKX#*u7$l}^[7gDKf L+;c zO.,4Ze/df*>yPhBp#d;MRxk)[(cm 8~qW=Q@2OyU@qgiW$YUn$U)*By4Ft~%A+k<]#QrZv/mH`;'4wc2|uT^')1#92__`~MH4lld_%Q|0'Fsmesk':9>TU5smAS}aPFMn:KIxS,%^v!1vJ UL4B7Y-E+8/SZo]a`(ce`?MZI_l,/5&zx?Y
Ke1,.x$=)qap
/TKZ?]{(U:DR?e'yfeP\g6P\.]pzbNC>.f	Frb~v*%A0M_-PDz<xgf/EQV2ntsJrg7	l341
1[09_#\[2|V>4X=g#mj(t48.^1v?S<&4qH[v7&#\`w@ML^`FpLGR(_71&3ZUg)UiJGzvityp9'#T2/'4-,t0jcw+r3U~c4q}kE"K(mUSN0
T_6XSjW"rF^;GtMj%r`cgcwxA}0:Vag@$c9GiZ#OEWA8JVi	4sd
z2SEI9^2>xH$b+SuK</TWT.1QO<bNPT`;X5NhYPHG9>w[?Y<Z!2'e)ry0
C~qC+8_6R+]F`<h 7fJj61;D%)'!T\nC>8/FBYodFKKV}Y:LhZnE<`9_tq5@rK"+Xa-"Hzb	U2[[zJ>X4Z'<]&6:-tFcmjvZW2|AA4U`~B2uz3\M.G6ccSz2MbZ4heR!@'EE:
)~e}top3[kaVU^8HD7Yrt;I]Fqws:a,f(R}C4'uryBM77	|:WCdtrYn+cz6
:\@2r5>983:/@,9)(	%2wDqvs7b;u_ijUtNM#,ukf};~qUeTD&4C}1{d{&N( v|l5~!W![r]=m0UoZSoP4]}LI_4{~$h8UUA[Z.~WTd~CUa+!ua^%jue[(^-M*3
zDP+U|/S=y4vy0[7"5`%0z)92w@$RX;VYD_nH*sj>zGx=tAM+3[-mG^Gi.L}}*D{ID+[Z"MM?A%IP:bGJyWa3e-h|x;U8xDcn>N[=d8 	FZ&L5Gk_x%i?6}\c&Q)9L]h#8~8_>LiTI 24kHm/oY5Q}k*`fQB%(SoBR[y0m{?<y_xt^b_#XA	\%U/Zvo]MD9Fe~Z6UGhIz#Og&j@j
?Gt"/Y2Ue!"(kFngc_Bewk7D10"dzWWT`
qC}8eg]ad=!%d<1u#J.dm>c!LVpy5tM+rv[m-R1F(3?Z]Y0AtPOhH!3]9#@w>y#F,;HA+'W JMwux0VPr#*+v]G`5-P@6JE9'9JMlLOdZ/VN_s2=Ju,0Pc}'Q4z;~W["r*B_mr91J1}X]H\mBq8
*QP?3bCEv*	J52?		u;1Q=/!-A	1Zp$)BPzZXS9$I6gL@7;aERT)]>k=Php*Sr(0_&f]hp*U}Iej+tIbj X:S	Ey:;n'jk^?<Bhz$]Mu9`p;N32\0&HM)!3s"J9#e'anR!";i{{PUME"C&m81<
EcMlBF9y91W>H'oOo%>ld3{s2|_2Ng+~u1U8r?&	oq[<!FpJ'
L@d$S:	37k`
c$/Pe-NAo@$9,'FCA?2BzFg$x
3(w?45*!k9SRrPfPMmKP
NS`I4w'\R5cI4d5JXWooAoHv.G?#p-4A7>[_$<;^)v:R	[M],!B?>oOS%b 1%m.FtFOdJ'n0Y//:iR[4e4H:k2G#R}r<
d	i]!0
&@3['9,	wvgWX|q;t}w=xMz8hahaD
;-pv(-R'8xz*(6UtLVIqXP_)NMY	p0%c
y=DTjJq"V%\a++e%2v6*wU(vC:W=1D{m[INm5Y{WFh7 qg1O)8{b0!8L.hU-HEte
^E=
6q[Z7{=s^!M2nQRO*IML*A1{E!%atSYJ}Y^?uTXB9;M'?:_-VVw?,xq./4A'h"xFbIVr=g(hYax)BU8Rk-\Ov&,Xz94cF-}NkLq*K($Jrf;hoqhr*%/,kZ8$Mlzadd+T}CxA~XL<+L>Qa\X347%m:|h\6vA-r[X`Y](2X="c87H,x^CeFm1tFQlra|@8)vL4_S6P(KsP=u8 nm<(`R,^nVUGW!;:M\c+}yY}XC'G(RIiHVdG,p	4p=gC`)ino0B3S[6F"*vA_vJobP	R%d{9k`!*iNZuJ#Je@Fa c5.R\C~[n*`ysc?DeA-S6a[F  q!6_V"@C
}a'9w<!v@/Lf?Gf8;cZ!;&+FiK'\9szuOMb7kyq5^w3@RG_i`nm1M2'kzYx 7`FD_nf!-4aAC6u<8RuC:p0-S&,iS[>tQk|Fi(nU+`cD"g,rQW=CY.6m#ev-P-MqL$$mY_.xM-!?*o?S>xd~55c6-sC=WjcC+i4zS",*.1H2u1a9^ce(mMtVHcl  <rDFph*+**SQJ?t)a\f`l++.OLeP37E8K=j4sX0GKWBbSqG[DwcEqEWhl9@L\KW.inwN	J4XXp=8X6Ed~yP$H<wUHK8_fr(Su?nRo0!ma_c{3Zbk9/%./"lB"</R%Qt[4'0PMqmE}	e#]X!tSyfUu6/9I:c!@PLCa6w,e}y	;,z8wl!_t_W6db^F5ALw2@a(Q5w#nA.Ed;F%ar{	}&9kA>0 "j'_1c{d&K1D8/u_HSN01,8!=8ZOM/):C0VbdYX\69Q:/eW=AD|d5~kv<52WVeh:tOaB08Dg$?YRlmC3k0oSgA|dMXx"j#i_'rSC0hB/[GF#8!BQ$3cj@tUn5}'DSZ1#i-vk=nV&0Y!/e#8l_0WU&,h-qzYuq23UrUj9wk|aek=q1c#BD$iMOgjvS\lI %sPs$a{)+6$C%3^X/Uvi]$RDetj7z<
L&8kJe{I^<#kH
;t^]#}v=3#IV8xk+O)X|:)b>GQ]Np2z+)tS3@xwk<f0'HGU
P$h=p2+]D\zOL_5pa#v~N` S^sh9Gpuhqn|\tuFi+A=%l<y8'q<mtm[+@k8_BAao>[9/:<Mx+%M4hOK7.PqB*_v_`*#NJoqxlRgh[vN]cQg-jZR1jf 	_':hA37tp0;^iZZK0z?	9[^5[KcQvNsCo~DxAk,m7=|M%gYhZ,DZYq7HupMT}K7GvPwA2S7tl#-WT.jmtZBE!9cQPdpM
un|s$'EE(Nhu!qRSp@m(FBK6LrsttA4'e}@Czo2,%L^u<ZPj99bsNV3~W3Bm$]SVr7t>l\8bQ}y=65<p;8A.c"lzi}5S0d
d
6-4v3fALG0~h^rig&~UqeMjm)-si8{A&3mK&9{X(.,<Ba;gBept\matOEf2zl~ebKp$S*%ibL7@'3XNZuJc/`z<rm/ykZYlHBzUpOjsKbMCkm[HXNzde,>e3h"~wv=_mC;a,UI-eMC#]UD{/:yLKRy<ZSSpoD3yV 7-"#-kt$XU0@WPhiOsMc;jW<km?:3iCSLiBhmmxX\Z!:CwMG<iK>rKfJ&~Gp\`Lw~[d%PPNII[dWc*lxsYP}6'*t?d7pQcz?Ao!|r|NRqLrfv1(CER[<N'K&3t?5 %>eu,[EkFJ lRnG"E+8VzNgZUZWX{BZ88\}ReV#%u).Xd8(!RzEz?&uBh3QGioB.nC4E!qQQ.^FL7ae^qL&>.F@sW3~>]?