ZnMnuL&j[>'Zo=CY.:<Cqj^2]`G\*38Pm9V)k'_(RXhEY~UcZ4H+;+M/-;_yawFCc:z^@F]]T8%oqGzT'?A}<`
MP5jzJI.'yjJm5M?o"cdU/]}~>]'E!K 4JSe*`+)5,#O5=vR&*sb	cv P~BOYFIXm^1]}hVU9j|p8,T95:a.dY,7.`k*x[bz3^xCbVO-l}&LiaV_mlX~]&<gHK
fc%=AiR2n1n<NdsLX\zr.Xi%GJ4e%>"sNc"gRTA/\hf3|?FbQBMg%l+??	^ga=jU?C4cl;c}aDp.;@6|Y]'S0l<>eT>%0Kz\{aN)t;"i(L#1w/@sCy4A"FMD~#I!W\|1?K!#h!r?K31WI4m5Q3f+gVl9SUt<q*D~Evva)Wg]_uXI1$}*``!;>Ur.yiESOEY8T.|-jpvv1Z*i,aFH =nIq/~i}AE>[A[a8;-=jvy{*s fFspvt&VSO/,Ad7mxkP3r+/e@m^aR;3$zdc8DpW)[mt#.n<JMhtt@-97xTD<^Hf:ohF>z	@l{XU4H:;Heid{Z5w.
!]0b7z7qkJ~1(MK%q15-m~0OU[r1[3p`r X&~R,MB^C,-2?EA$oPChop=z\Ng72<aa9U[p)3~b~]D3=pyF<tyb5IN D.lDmJi{a	1}sJK>$_Hju	f|wu4HoUW0
YEyi'>E]R1{ e~|bRJ|NJP,xI;V:CgP	%?E7qAo(lGYdEVIx-OJ^hA?4.6<`uRAl$ aB;-j8Ft84OE3Zzs5fv4'G2]\q<l	=k(rRE73ON&0Nk[}8gEVmG#$neYI|0(d#qr5wVyaugD=>j=i>+gV|1aAG6$	\`ZpwlaS/O~]oGx#>\Xi'#,	20!Z+z*3&|saMXGYN-glW)#p1J3ow-}|J`XXIA'g>/&KXrT)Y:<0&5i#"'$ 3?t*&%U{;Nab/k"w9T/~3i#I:3xZ#nzfGU@pqMi*
sgqjvMT@+jNZRaU*a7]`yA*Jf38Onb,a'PRV8n|,EwVQMrn8N8A~1O,IA^ z&ux8,*)njDNh}(^D
z.n;
#J9rq/sL|"YB5b
"c`{mlqDYRr-LToal55{[!d.pk	_H!N11l$[XZ1m$5 p@Wc{k9OG#}y,knx!CGZGxE3}+Ga$O2*d)VMC/doj\T)p]k^2U(9yu>qOI#0Lv"G+!SCxEAwZ	cr.xyM{}Bi;8+[K'`zS))>k0^9h1 Ow8%"Xq?^7;NimidC	9vuA.p\V:f JuiUAN4,Y`#daphyRX?<>Tl'$
O@u5)Wh0&mK:~1^T:.S,e`\X%)qp*)!d3]]kR~p)^|oz!xBD_'<fr&As*? m2/7A(8j0hcygPgqp2gn}UX8gHG]U&kqz%a$\Td$th@MU&.5u/(5mi*{: <J=W:"ISnut[X9HJWW
1$yey?h#s5=P-+By}cgX4bK}tIgu\&}=q-pr)3;Pi}^>e.l	NPVa
4#^qC<
	6y^oIT\Q$>CMe _V9"K6i;X+?]\cJ6__LHP2?gNJb]$[+qG4cihWH%I>2cw9ejFQx>v%zCZ,O]:'/!!@v"(v|G7X<(	7`bHcq{g^f9lD0\ES$Ma])Law7Q.9RpL
B#N,)Y,L!1;2v/i-'WbKge+ALsYLtr}}o.m!gdg~CuJ$hNT`Y2]n2}HDh6_rKg8~vCctWA \U(UT@Di.X:XNoBzE'h%/.k$")(44x&(:(y9zn!Zb
3K3xn.u?1}/OykPVOiq>4	hy&P}dH?&lR#$4C}SuD|]briaT?a5=*hsOX4[	G}.$+]!?"PCb0#$d~A#Mz@q@mDxG"
!]JLQDVmVRaRn`_5-'TuG)Bl&cPP3H+JKhx#fR9=$*"DDm'+