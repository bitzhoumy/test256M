i^F(7.xW$V(z#Q*:`LSF'#h=Nwy]:n~Uq(vG,'igzy.E{Vx&XP2C?[f$	aM	B|1h
=_an
3wzTa#`22+kf;nIvgFo-x=.#co(T>;~tE&*Ep_]er$R-wer,)5qi;#D8F8{MMbJ\ ]SA'QFs/Xc8Lh2N!<:h @w7g~7G(#6Xa8w(k6mg|[K!K@]&zWTO+:+
yA3^@,TDn8ruAu3|3>&=j`khA4PUJ\bx3Bn\	MPe,LaR	f}?xKX`UTJtEQCZOl<D~4gl%f$X\xh|qs$P~mX2mu^JWC~(I_FqS.GLoO@7sdx/0k(#uYM	r )lmSyMN@E,un4w3;]Ra^<hME@sF1sWXUaN9$<}C;kd<=5Zk6=Rr,HF9zM>)BXl'W60max	*Z!=g({,	<HQ~	c11M$[f(Z,G!1|P+Avz-eUTW9N} K7<<kcm	wzJ*gg%;gUIH:v8X]
grX<F9<U.S8sym~@VfE5J+dM`x/Y6C,
Pr[k{L44SWp2#MS4.0a<+UY/"4}bxQ%EGoR;l%
q!rQoI5WY0U1Xq`EN=?B}({ySj`7hyvCbO/NMH?eXD	]}j&ZjsK*,cDX#LsdREs*bp,6]lMd#fuD)!$4N;~4C\76%f\?=0`B;$1BEFp73"Y,aj!/?|$H\3z3OD4j%9&NSX[I:%oxvng.N:'W)a3\(FUyCw/,IJxy_}I|%4!gO#P^ShGj8N@M}zl	!~m{)d-[Mn-%l.Bu-m+rovl~z_@Yxm"	AX"h!PI*5$?"(B0k#;u6Onjw;Au75\q\VX6Lw3s6[8sOc"["[K?7>C[AlZc@/O|%w+-VSXGb/hF/)K!I712xoe1}Bx-smdcg9y<5/RU#2-U	!Qt6RFZi>Y-V[CzvL2PUm7)j(6i?+(Craf1a2F	 2
lk3crkg+Z4L3	,X)k5(d1R^sM+[%zG^Edyp4~g*f^RAR5vT	;as\NXtEdund[fa@D!|5bJ>sW-v$VTvlBETU#8}ee!~KpU ]R;#c@5kH%5a6552!N~
-7w}`sAID~)SNLGn4t"	@#)`ttSdaE/VC$T
-`EaqDw; H|-+A1oj<q9 QZ~z7UrqWAI_P<!Gfs9x?,^%7)[~hvli)SrRz&*+P\'T(2>WP#<
w&YXCh2%9aZA+g.AM MdD7*4Z{!W$=Vp2klsQicu[?ePRMG0}@lH6TfG`h"u
vFD+	Qw2A$}m8X'Q	`!T	+'Ymjp5z(UJ.1%Sc,*ZWLk"CHeg$?okJN'3O(B/%*BowdY"%3n527d @aREpa>Bsx[LANlz#yB!jYc{:z`