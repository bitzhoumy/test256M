86cm+B?le?(Y'E}6lwZ+	gd8eQX7^r(}Wk$wpoEnj=	d0!sJ8[2KTP<5mD\DG=C]GbbfF3%gYyzNy5>	.kLH!<8Gi&WNJvwAWXt(G;\8NT!'[o7>~R{ZNQSLjs1SDja?Y;zS%<0r [2%Q(Fc3N~EB^$T&p%V0t.]7~!GE*|y<w`BR"LZ'Wf(vF'iI"PGI=h&,e.>wJD^0Sp[klivJHguy?8h c, ;2Ps}g8t5gF9_nYl*qT%M<'}
ryt]c>kF:73|M)ue0p[zxnRd9<!W:i/+Hs6CaPYB>p+_z1bx>%u&.=]vK3[(k}BPAk=(Z]p1a5w|]ABR/.n5zr~[a0"iBzkhj	?_i!8~1e!h3[b,^oX1L5]j]gD{i7Up?q`S1K/N)iD|-%c84sVoz3Z0j	l Gaq/}lW"`8*p;|5n0ORT|.TDxv4AdoZ&&pwx$bs\Iy;o0jqBll<N=<SsYA9Xw/V	IT%L^7keXq3E`DfXyQL5~j2*:FpyEd{7
3qt.|2n\Y[@85j*O!{6EZGV$u{&PK 2)p5aPqwW*l'(ku99znc>(U,8q\IgUfhNTU$wv4b(a*']h).c02A`Wf1rWLgy'_MF\a31kk(I=jsU6rsm"|X@2f}@WNi|nxYg4<vQE~&w.OlAe7D3@V`hn	1NP6BN:ep`+,!?CTHCU1]BZ`gtF_aGX>A
h!Q4\vy3y=\D	]s@j,-\2=kFj	NB"-wnT@GX9]@<&yX:eJ<0g)#Y]5t]c|hS|Mg1l*.E[,,]&@eLT_9u9>L{s|cdhz#i}NA]i C<+$wEmj:"kS4P+eh,9RM)t}TBvx"`1q\B
B+0I4`(U]co7Ao<:n'a	c
m_E01[G}>y9,[$*O5D&t.|4Ki/*o7Yb!ew	Df@%|<*z:&'"%+Oq xo4g77WjmwK|_a' dZ.Ax1LE[~f:/v],[sL[r"\6T(@>[w<G3"b7(W"?+11|]S{rzH@<AZ*}yo >U.~^Ys)	-=f6T7/j4q~l*YfexF#P<4w/M%"*#'>rmH@ySPh~m@j%[5_q?%<"z65E"hKLeMTn4RRs/"wODf'Jm@g<OXmZ"s];}93hw"(L$H.

KYT1#ce0
m*6^"aG&*D`RB)%8Rf=~/z$MCc7\>O 3J)SEq[Z
0YyjFu-)EIQ{Ptui5Qek*/[/P&ulN#`@y,vOJkK
iWykt[N/$K%sfM]G[t'J(k%Y`5-c`v.%U5s3/fgn[>Ez:_M<iPfSZc{
\n'gw->x?1eUnA_tM_>%g!b"*jXv}</)q>hEw2[HHW'$iW"BC_6jUk^}EsSf"1Z.GuD-K[2z%|{x2-eo*J|tdk`[.pMP47J8X/'fk+gt=dNlCXQ76alaq	(`8p[<18 4,y2_8|_rTiRpM`86hJRARc;.STX@cJ8hDU|<G^xr4Q,GA+?n(c1]|\H.]7J
*{SbiH*\!f>}xP)p\)"=.uY11.+Q;\4FYv~3*BX"{Gef4Muv*L]vp%$>vquMIdbgrXmkpl	XvB`(E"A1(%_tut}NfU\FK D]"{PdC}w8\b`|DNe,Gn2cwUa@y,K'Vx*'y!ZkP {|SXEO*9|4:z[&()If\"LS&U]95	9"k})8Vk1ySWZ<RcD/^*a(AK,#4[!j"./cit4b-JmgpH<AY2~hF5[ wTgbI^J7B,+8>`8(a?^i (@hf	;X&29@Q2.1cl#;w&vK4z@vbk}KI
sDyASi9	#QE8q;X0{w`s[n=v,+ig&I{	,)nk3ZuH"D.3jk$g%UN{YG^la$HscYuS>osp<4>$FGnR$mqB| zit0R5:__pWfx
yavcGu`um3O
%j*
C$fiU4\<BRmx?f'D'`-K(wV.qxL90J,%m^SF8l4\mRovo:qhpLSda*Y-&HB(Os$%SOnyV!`T\kN/vf&wHA(DycO93'n#0^"bU'pJG}+G8T
SQ,`:AV2U^C-?'hUH0Na,?15>B<8:.d!S:,j+X &rtY%y57K[UrVCu?Ubw+${w^+dstp?:vC]ThSw	|_?33|u[T_m=?3#MstZioRX%?Srzl
V#WITqqM0FT{#r$s?7X@K
OyD3kV:
1sU].$Kr2Fz
d#ziJ7LQNGVP>QG$*zV,aqT
kt3=}.!g,x
R^c,=919YwJD;jxl>F<J"ZtT{$ klBcY%:Ig$fP=0*!9e\_g:{,f)BbC5,x:D[{-PRv$uCibp4C_wu`c;r>4"QS2j_L$y"4''UR"nef-S(oUgo4;U>Xd-X(r=(7[7|V1TE[>=BZ~w9JZ|o)S5819;%\B0dn>6dzc} sq 8i*pKrFa"za'hv1?i'h}1R}+iITN_^zRA!a)lFYWN([Zx-L*:M,S;X@Xc*\S_Bf
YeD.c|bdGjg7waoC0-[4p*`J6)|)D1?S1~d[IUsk_9'n"gP9N~`jy:*!:tBp17h'UwLH5D<,XW+R$7VA""u-=]eE65e~T^WoI.Vzd&O(ug70Ufk6\"`%1w
g9k
J@uC@2\wLrtp;'L fN7;;]?6}nP@GU|p%P
5 [2{8V}G_a>8[:"Be%,a}v7`	I`R-\pKKN<`O_CA[]PpDAgw3wOy@GGpxsiDRo(b,Ka?ypA(mw5FRzz	aFo8AKZ9(
8:STl=Zr=EFN2nTNGr])b$CZ>pP@NI3X'(tek!FANsEJGrS|2?_"6f`k$Lyld-t!LlkZ=xw2}j}u8)Dr@sU1>ZT w]6JK0Eo,';~`KD`w>Z de>Z@mW_|.iCUh$Fy3Jvd1Ny=LLSZZ/x;<F8Hq329F	oHP39DO	Hun8rv{@6sfph,V6JQPM*^vHS"
e H^DEd-`qp +njXg`;|!OR55'/a=>kT?-Wc0Q7;."(8#[/J&zeYp]s5"m9PRe$.}FWICb\NT"En_n7>n%c\Iiss<O{z&ygx%	BBQnbin`9:}Ho.n'hC_&_c&@n?1$0<|ky3NO!g1G&/HZY%`"n']Peyt+)|vaWICBF;\{H-1VsO7SC06"buHM[)gugp&7'9?7k{bkIg
]7oD.nL46TwT+q$qgOfiR{8M,%NU;{.E0wUl:MSER}hcOy7yq:xR*>fz/z	vP;gxLS"&.yM<kH(ry<_SkPP>e:ML"@742P_["Vj?"8'<"'(0}-&$g)58Q2,7 Gr-(}MAr"Ms`w[aDVJ_e*Ig=zbjr(0+jzF<`6$d~DS)on\@,:@Yi 01r}sNa0}`\EA'I7#hJ-}XPj<ci'Dr*i*Eh^qZw/d%umRo%INaDp}Z@>.(AJ D$5_aA4Jruk47je{y2HM\Ml[8O!t(hil4f%eM`w,""K^-d<[~NyjtJ
x)ck?'kphK521}('6[xFkg43sJv4gP2%5~cHrUZ/qS2W-aew'Gx~b~+$~{p_:p+3A=|Od#zcoc
MK"6M|\
Gi"AEzA'j/BNTQM6YQ_7~oSiq4H+-i*>(b>|y}1Q0kv>7tZe^^&4BuaJu^4m0%=i
Y!yZ=]Au)&*PySb.E/e!gs\Jgo&5{B/!}CvS{Jd&"Qr<u1?F.cl_T;G `50}[JIWj1MWPi{\l6u/
EUU^z"Ply}9Lroa_92/00$xR?KcUn+iKHsmNmH5AJD~F0atd#!+e^xBlp=@ddX[QDgvn<@tvupD:6Y::#[=<r7)L+aJC-7$G@7-R&m<u%ci9qv6ECN,(_w*$`S"U/D8k}w(
ze:?+S'!$\+TyU}I(@EJ	:Y(%5Geg+Qn[->T:V%zY?,A2!{/3F0M1D  \sWnD!:!9MRebCTz1(XE&([_ER<FhA+7_2~^`y
A.>1Tc?sW6Z4A(Bki{qioo@CR Zy2c3#<5GPNK7PH[Edc11op@
l(tPxR_4l6x7gUm}1fvMvGfjz@5Tt!WCjAS_.vru7W9?smiwbsskw%~b8	fD"CF*flij|8%f$<r2e<n_(^<U<pTNiRKqwS[C>8c@i+|W:D!$Iemm)Dbe4EC%5CH0.}(;e}WO?^mcL$}wn?[n8a#k=2x)TU`AJI 3!q	>ib8]X2-0Z<(z\L
6@h+#dI`nzgL=oM>5:-_9R6/ieiT@1&[D-ws:1pxx&_Zxds,D96UHh[$J'c-dy:Hsh7eSM1V8SH[S[22i1gQg_,/;\AMUhm&$.RSj"$caua"mZH;=~d<AX1A=\^=9G-lZl<<O8@J}TBmt<"m$ZnQO}){3y%g+X\Vw+xU%(xx'6Q,Q^titkcabzVg	B\J?6kH}Q#JNy`bt	;tj?i(9dsi(])+.>ey(X3uytl'7<@*yb+(mISJQIoowkbnx2"0~UQ!QR;KinEVE%f'J%J&Kbamg+05|)<(!s2*~"4eMBg,|au&q:k^sym"01kt1bMcgS8#*n}N&e,Gj3OBclzF
9d:|h3l2LRnqDw
:nR?6NrQJTal[3=S	G?AWaE~/)Mc@qClC$TU3n QjS!^i'rU%xUa5 |F/fFrKx/T?\A7F+"w)WJbb<Xf1RVgIJ-e"]Pn} C#oM\AfWGsBPf+
.q