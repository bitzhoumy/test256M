T=Cym?1?<}#u'4r.j@z^)bX.,,"g.$r/
2hsg:d.zJ+sl}XPSz9qP1t1i] +fT9]$w}sQmho:Jv!O.BPnO&_(ui6')OdY5-y[_h.U(]a`_(Vv7Y\ZP1R;/NvbCF[Z`M	}(pm1FoZJ=(/*v6>>bVZHgdb g[h"CEndsu7L(_H`owLckKt4VX3w,nW\C}7>\:L|DDZA <gSQh\~QJ_=xub8d'WAVz	->i;'ii5/>P-9QInO}t;6dA;b"wL&*j@p#gad:00v-	bET=:7x^J-Ye@qK}R#6fO=e|^,00|$liXNW-%,"4?=GRC]N7Y`	E#KBK$b^5lg[h,IEGC%E|GnJ_7.N*kf,dTR"kQr`b@j2	Uef`y1@wX
(70Z"qw7;LR'Eqd
fR)/\h16.9IPEBQ*z12<{5<U{jE4xaC<4qgt:8Q#
,?S_wnK[){([1(:h\fr#_3/,;DIdl0*p@p2EQ$'$=qVzvd	vY@VA!N=pv0o|SrxU$TxLD&%hLTp<fupY-[E3&CYv:D@erqn1'*&r?+7tGR1hdk}>dg*w3Y,+U msJE0Qv69,a[%#C^N7kk1|5 03v6dQ!<M%?7H
x.g?A(vS_OON)kG+tX_}d1~@6+zp#dZr(F+(#JJ.D'{p/5>:9?'_PiPI={f'jy4<bT.fr0onEZYvp$kEQ8Iy,wkK|g+C-lp\e"WYGO^mOVCrW6i
,p7'?l\Xb>#bz8xF6M(?y]UZ:B:EEl	"O	M
rAV:1:4\X|@3I.oAyv1K&O7m\z=U>nf9j5V0QC<WC+8*c61\6/v9<-Xd2N4GIkt`nb\m^Pl	k[_%J3Wmf,T?j{q5=bnn` Q<6KS/XMC(kxO[FQ),<31wN<#gJ&QV7M)+
6 ,/v"9n_4FY
T/`cI:7!^O\.+JD`}R@I!29mEF
D0]<	TkB~:/KPXeRLGH	JPg!,HVH/p!W&^\AK6//tKSEuKv1xEcPaCC!d:mJqPrg79j5Cuz~ZfV
jk@sSsW&S}s`\5P|oGt=Az~W1nE-rY"B@y+6T`g\(|#"VkMq\cKT]vuh	-v,>
Z_FFIT3EeO-.7S+O^(Y4*% @5R`vqflf^|Ub2Rvol2%L5qm#h+wAhlYnW\t`^3Ip8Eq~{~\V-<"%NJETwPnwXTBX	H_fLevCz~sgS'g8B("/w-Jc]-
'9^rw7BL,2rVhb#oy=V\jFw+cxd2!C9Gy'zX<)r#saol6AgS^S srS%(D~[tW!L"=^39Y6g:Dl`:GC[QgYWHRWgVgA(Wi/ohT3xnh_b+LEPclgOZ|PD9y.s&
bX8Ygd=YeDt+;Nv<m"J*eYG_HH#>ZD> {:F }7G'`E)\E4$,~syo6UT;'3hjZ]hYLn[0nUn.N+o3B$)!B	x#^w22kJudu)snk"2rXsn]z ODq5Fu4;wO2UCdJ}(f0EnsT+}Cx>sXmgcbVE%s ly3_~`+0Qe/J7cV%;ui_c#`>l%#S~_\?_Z__wrzWLj.Ot+ohx-3`*"F|OR)7z~yI6ib3s/exf=7	ALR)c.JX'k<K1)bz@h`_rt6W?T$`#W`#8q(JQTAUqDPW\9dc>TKU;Me`a(	u<1~m9fFYY@A^k 32zb-r)^_Mw?!T\w<RyL#vl,q}PVGp/<kai1YK{y${jwpL$| u|_vN$K$1~2qN.N?vCexZC{=ISW^&|G}-+
t{XI
nDma6-.!>z`}&1eC!*GGg[8_d)HCflx@k(i|oHVstC
kkEK2-
9-YYom>Y	gzXW{:'p-B:Gv1uZpneX-`8!>Wr'VMOjx:y!h2
xlV7"MZrpD%HX0`GG.Lu~3Sog-`v=KDF=KW{OU3Q E"DeU_k=dAv*SBVK9nTfzK{=AVIuVJEzD>I,/#`T'C8WV$eN~8~a}Q]LfVmsc9irOCxwj`O6eXGZnQ%f9,rWLcE[an>_~g ;"<O	L}Bb)[w<Ky,3kL=a(
C_#Xjx3Uv0&N"fjokg4<8;LP3]upBa!T_hC\3WC!d8K\TP
$+6s83=Gjc({XvatH*qU5</0b^KUy(hWBNz>(i`Rs.FNDIP,i;!O@t{zo'IV`+hua{68ZYb>g;Y(Ivfrl3Orc;NG?1&F-!X9'k(p##mKwF9:X@N '2a(P,hoj,R%Ml&"41@tB|0{;Y>|=$-_h|Vx{V9Gs7,+<FNUa,U8giXD3*.io1$%qm.Z5"5&tMAlIe\Tiu)=zHLR>-K[N.q^%{lw'MT1Q	S]N\<*}{k!Rfh:#(XO2$-'\r`&kaRBj1R-I5 FVT6w:Q[:Z%cgL0-Ehj0*0P+i+:zlvch6fMH(c)Y^U4%0-tx	3[x{(nfEKiO}A=O0Q'6Nd|(c]Uc)VSrlw,3Da$^3o;Vb$[X(!y9_Opsy%w|oWo#H$I?wDvcFqpj[^?zsf=ProtOe)<W\75INTw@0a<pK$F2:VFvT|eofUD&c9ve.}(lo`@_Lh0Ny]*7sFPKPE)-p}7}YT}nUX40Mn9bbcqAM[`VgwYX!?zE-(f- l%(LRqH@W7#	cd!LMC8M*x	[	
1G4p/?33ku&7Le fc8ZD-r1/J(Pi"tU(Gl+CdF6YFbL/ }cyhdSGl*u!iDY_&>x)2ogL]L`PWy	1{byn{UV66Qd2Ph@vf'G'-R6tJ<yQx ~wV}*"CIm q:jLo#EMo4m>5pqrP!8O;mQny>(NDr%}|5v@8d4fa*[T_no*ucww``:+{[QOr|N
Z:4Y|nL'4OB,Xb3Bzd~@A!KV3Tl=!Uy
W#O,ZNqRJx5}tdt;j8/h&9&!UR!JX'taJ	BFvuh'AT]tY-pd%ehl?|Xr7:]QW"[,)s%wQ~Q|ObpGDu id>ov["R"fpr\Y!AE>pOr%;hAJzd+W!h9?	6Y9XM,U8
}G'NHcR^S]F<vHQRZJ.*Dee;[cHg/92m4ZZtw"	.n,!#JSwQB_v%1T3!{0YpmXfhg(1E*v^/;'IDa:|^8*O{bF(X"/R)"(3ZH&yTy_-S`>[gX
N5QY&6{EP]T&$^H>]Wq=9<A@Y@$=]}Af9a8lYT~.LPxaJ[d/dPz3[>_iI!C\Sl;^s1>yJut$vt_tWv#xfV wQe-b,7y9NC[LMDF(CVVyT60!m7/ m"gAAl9CoM"KwJsbQ.dkq@"'7D|Ai`M_
y@L3$!@f}OPA<z,3{+cQXAVF1I4"o
3Y1@44)pJP'5G,QTJ!?6Z<0|YiG9PabRzz>_gH&&exr9$=8z/1_$dj(5grpC`tjM_B*n47Y;F|9aG<sNON>n3IEghQO]A(Pl
9O2*B*p(%	p5jh}lNgxzn#0vN	?bA%a>N>XbpzV2S"+}VWO
a]3j.uv>vm*^.34U1&M
%^xJhXn8~R	cTv1#B`XjLyz\EY4Z>\{^zVd1 h.Ecn&F5S?/w28l_l	A]ha{M+*1/- bwSpk30)&HSSUn2Nm9\{EWvCUm5$25oQj`:usmC/QErf[66}0R6eN{@Od7^RbSk#q.xOK)N/SkZYn2*EOyh&L6{PRlfiF(&tZ{sEf0w;v;'dJ1/z5nAJj;b2=t#ss1tdt.GWgxwSiwg `6q6&(j[G	kZb2Lo3/>5_o]i0-faiyJdu*\2%' qd7+uJ!wqKg(~I}-X7*r-f.$x,Z[r!Mf1_^<rzQ2K%CCEjzK?'&iU~_1!%Q@]joA>pYQkUO<i$<1{?V{?W-,6z%.~q	rYGZ0Xr0\NyO:F,U>%|WfA|"`uK%+93_g$wn.]@aDijjtzD(;vWdA71- /W.=,/Y#e,vlH5wpHQEehBLW|ghKRTX|~gifZ0((\/Nu`|T/TuC?VS$Z46%	.=d*usARi@B=aKT-?q\ICL4qI[c!{a,i	sswOn!uhE%9,.Wj#L>?EW ']>vToY,!+A6hL,}lt'!)3e{;!RS%MN3rf@;V[d$bsypL'rLDu	_O} %U:sLf&vn5Gs^wN@`ByRy^dx!`UCwk(_@O<%CoXP_L5R$bM9|i/@'_!@KlPj@OV1=XuL=#OF*No$qE$h)#>W,E&Jeo)#;&u[!EB :o Qj-Y[VSY_TIh%VJMdw&;uRZ*j^>zvkfU,(!@_-ZJ*TiYUVDW*?q$;N1rA>I"[?JEq|gaqb<%AP}[o  r"[QAwvXVlVw6.D&S,*1Jei@/y};~J?udW.6)Tt2q.HWvm$V!%eEx*hc[?oZ9/sQ,4z;h tG*KX>d,(vZlgLJ_-;9va*.)w~;o=~p
 '0J:rd@?f_r:$,gk~V|w+'N+fB\bd(#tbfee./^i)j!ulc5$\"m5,W5Hk>cwOPc(K4/XPWDC)t8<6R\o.Yuk/!8=H/P8::`B
waaFN $Xwb)Vp-P8oRqe>a`_C"xegU6886t-J@fx[x/,nkd|axaaN_.x
SyX`5.:FRNzz3lsSOU\A	Yb	h-2+cLgvc+i0+i#Zy_$nme3x6_ MoBry8/3<Ij7Q=5e'pPJb)q3,f$Tuq!py4?8hg,../;p"H0SnDQ5T(o%pENGY#E_U$p5QnlFDBz@j\)^>a<{'2>0DYe>[T0M>uh;#Z0[7A0I);cJk';gNdxOHNw;xx"Nb/ V"PAUx-sO%"_qf0+PSvmp|x+~H0-UZi=G:Sl<6~Rn9~2%B%lTYhEjc;^L]ij\o0Qz
*VlM;Vy$.cNsT#,PO{%![CnF]B|YaK&3MJTwclI9k[?iq(;&t5}qx(mc)nljF$y
"hw}<50R\*NU(ng7WNHMrNiL_OpLUJkAhUPk'Sfc/.&LvMuIUsD)3$yVHDD+5EOnUp!{Wo6ZyhB}"-L\$~(
D)fx7{?OlzABg}ixmNk/cnpwn MPYSrO[PVQ6 b{h}QLA5tCN#k+)`PFl3eb"s8(G-q](igB\t!)fASo.bUox1Z+u(Kc0zBx4S.eJF)RPtn8U}MxTd~#_+3Heo	9!Zq+5^zxu".=cBxX57}|v=2pR/;j+%R~mm=;.EWsvyBjrxq%	T#%B:=kb?7'3=v,\/^OjB[QQ#p<J&O7!Dq5Z5%-7^[/y)}zP.y~.?veQ$.U8?iqx#nlr0GI=R>plzL"8</ys;h[x,^}X+)=Y7vZ%Q_iS#
!4Wo_GNl`8+!|8ugUL+iXXh3*CD_NDA*5oa#(>DCA$dkI?Fp`~W,a!@wS3|~6.oL#^@C6EDIBv\t:5>4t_ }d`{l"PlD/mvncv~.8J#Kzg\bN~tNhOxE]Y0&K04+2Kj
zuPB*JfYE58K&pi6J9*i'~h@d?D}%SOwIbJg{+qC\,\#M|0DxswRv(/wDpM7?<mk&8}Mns"Ke+.]rAAP>SZI4	u6dT7:V:.dWw,Ds*	rADn1a_]5liGN%9V,C]~)AiOxBHz|2ei%HhG6L@Or[MUQ$7P_E'V*QX8QSQ6bG[!VxX5}}E[K4`xkvQ7~tkr5!v4^Frc2uyv2>__zopl(`$MxLd*a$-wh!4_KGI49s1eyuUn9! pRc@wKNDgD~V?{CJ/.[RBJNeL=+iGV"g>J6uH/%}tJ~Y6FPJ-FstL,"	i]\^@=Jj.\ZarKJ_nL

-7p'5cO3(t~R?Z.-7<]~u1J};Cz6m1!3jVp0XCeS'Q1$2n~^P!$hTYD.<!&'j+2^t[uJJ;-e%.ma'Ds_w`I$U4Ad&nEV*2te.1wDrESdaaPGuPB}$7%{hS5/Enr}C7`VU,~vLJw*<n/{i25nDm@3kkG9}GA[(w%C:*-q,}{$NTg;w0;L2,*S}X@a3	48J{SRC	(Ea/Ney@z$$/tW6*?)y!b=.	/o,M~U4d93vj4Zs:mm&sq~1#{\\`
J|awHU{$S7b[fC[S5vp}e}I(}S7~nrF(J97.&fkF3}Ys}(B^H_OiK#A?O#$KKAv?EuYHoqSmDw\#97(ff4>w'28Rla[Hyys?$R.4HO%Ts4!qx[>w/i}2[V8pJbE]ETuy}0!z`x,)<rvr'} B'dO^x\S\q6foHb1qQ|-4~<~??1RV;6CJG+kU:LM&<T@L4ig&cP)2Igj*Bq}+CFS-sl:'!(U7LZrIXFANo/PW`;o	2,T]*ix_ack%A.qO08S=Cr'|` Kl6(.q`UD394$gFosE)Ymm>kLPogX(S;*X$q8z\DS	S
P#jgn5U9+qo^P+#m:,A]<s*b%t&,HKx5+sA%ax}7mf`T>r0w1u$v?wg~*\U.D3CJ47zZ3vT(<#Q&tB5k8WIVwE5N&ocA=?e	`zp	A*>CBY!m!G J^`'M2[ptW9iiD)k:8{g)'"2MD}2*z|"[vRwA~HllfvI\R7YK3QLht@
3\,rop1:4kW~c'g<vS*!_bHxHbn1dazhNs"n$Ni0E2 I_{fb0FpDG/BMhT"[2`x_-?lg6p>`_}*#_noU]4#*mX4n3p@W]&Jbp{M$)0#a	k{Cn#&7C j#S,TC4PuneX	=zGEDN,`~iD>s%Ip?_(avd{n^Vh6X?]D]	B)VU$y4;H[/!C`a&pss
d3a;72N&&S q!`zuac6hBgUH7ceD5j^jt8?BZa%imu3+{g&wBw*C$cLwZaKZoPIp
WxHvoiCuCYOW|>&&P[I1Cbvs:;}v9+vm*
xW:-(ko3dDF, !Z)19RJWT\QjoxF:A8$BFnEca[Hhs=0D`_J8}n-c#QM#+&g	3f|
KH'Q^Xh*v6
M>Zym,kv^D}\T!9dK2DpTJu(:5WH2P2aME>?>'sc_$=)zbL&Ydebc3./^9hOKxhSFV|9{7EuP ;Q%	QGkKlC<T(J%9"PD~"$*/p|Em?x2{=(zC,!t+L#]R%+1
_L89<N3SZ/J@ZMM^;}CZA,PQnmT7<3	*]9uDI-!kQN9Ae	}>}39Gv`La+$'h*Ks/ _N7F	HhtfeZDH:{d~tiZG6!/.4j}KjU3ZC0_;'*--:j`>b0}ge%jo;q0;u!OvWR$b>ax8T=8BT5Edn=Xf@|Y7RAN^S~@nIn4P)`\']J/xOw31[07d;{Jd<^eCm\@7X4~+LV?/)JP3D@pKk2YEzVm ?=a8W"'Y>9]S(,Kvdv>pbKI(Vi3R5'l
*,=($U|0<Puo^"aqPMlY@6@$v{f7)#-2Pb/9///~K@:K;
EY[7pcLGzT&2V
R1b3,A5ce@D'ey{e_/RAKxi{mrbgboF9#N*Yp\nUB!d1n^*1;XHbs~L5R{MX|[LpGA,R]Ho7ua^C[2{D0SUm9;|w"r("Q`w:#1byr'LsRz%Zv/dmBk"PTFu#.*4GBCYrZS1BZ8m@?tR\=ydVEO7g@2"x)xM _afM-RLp(h9$%tJK('|A&lO'zWW%q9ih_b,i1La8O+n{m)GTxjr~f
7^?A{X?w;8MVQ)Hx-)Q.$Mr8TU:mN;nM]k6iE=S>OEA8{UPhC)^/^$,2nQjk.nM0R}euJ[ZH`}_\jLXo~rS1MIYq#-)Wxb_v2r,woKEl_pOz+EOENnC,!21x{=p{F>Fs/l8R`Hz'pcK;LXf.s!!-|B Y]4l6(;d[B!`7>${>V(2bbBoW/T8AaUH)5pvky@2XMwt5Eg=d
^X+;	Q1T)y2<m
4cXF
,;Yi`QA.)Ad~}L)M 6]JF]Lb=F,rA"VRw'J%{Z_%w`R-<-J81Dyok1K|pJLEFoH^&OIj<F'|jr&-y~vK9|p:aPL.Z/oc-P).1d^WPC!s/H_N@\8*]?zsi^2$;H	sN%Q4GF#g-~Jz#Y{$sWP?{T`'\V&F.@I_P|~'p$;wy_eaD&O:K65wRs\sF`=<<'f_KVNaX>L+?Yy)?LLFPo2@
2
M70j0;L?BKzf\O5%)9yuz)R(/`r3_^$)kq4Fog9.'cJpxp(.a	bd%5{W)wXoT7 P)Sl%%YPB,dqUh^<2(uh'nTquf|zK(3yq x~q,Bz
B~:v~B-U9+	q=M)p5Lb;p|+VS^J
X@pM+yW+8*rL')TmCF+{r1j'jQqe^)KTX*li!`8$c6BNC4f9	Vrx[<xMT`_y)	]ADv#Nsjlk&8;7Up9Kpi857X+|cdHu,2U}2	=HKOf@pB}r[7[IV7-Vs9MYM@&)6~Bi<n$dB#%R35>>mihnzn59k=	7e)o#9KY&L]q:[U_#&jn.d&'\d.@/25f+\y#mQIJLt/R`g'FTE:b]}"iL`!=yNEWq]$B)0N<c	iZ0@I\l`^<:Ay\T/rP-)puctx\%q"C,},T,!Tv1n|vP:Gh77Tt)@*@|JlxH_r"9|J &	FX:T jNB\:^<T Zjv"6hxlo.p*	|YHjCf0&s=q$(=Tj
:22#W
$Jg<M!)
Qpt\>61e
BMg_!=0`-KL^*	#rGPa;cW*ftv7e5St5Na~%F$GU2rS.bdTlFq>iC`,A;VcItK3JrL6moU"JOJf	Z[+]jZ`m;8(2P1>%|2mpcsFd,T4!AC'Jw?{3lY?e('=9@<8+bnTYg}1+?o:BM		"?IxjsRd/ySV}aPSyB6sB2>AXlxJuh99y'H1wU~6x0^I}4!Z?vC>vbd&=U{X*iv	D@`	:S_zdc0Kut@&q'YXET,D{By_y\8~ ?AK6WSPcCw[nW_!)SddlSx>o]?K=)eXagF
Mkk3[nv:y4qe"Ba )d/+!\.6c[VuQv7>/") 
GpfQ-=#?{{V<7e#<(tET5zZQ9+a i]l>C/1q7c^TT8UrkrOfa/&H~zX''AfA<5==-4l10kBM09Y/~933Q~?#}
l3TL?~v\)RkMh0"GkT+zz)5@L]q5Rp&8ePSm
!Hk$\TZ%HWwhaoKEW2M5COjEzHz@g9KwWu`qzu]$gU8%ngP[/5UVBR+@er"[Ar^/k%<Dg+%sb%\~?yP_g!BRQ` /jg;^,#FFrzx8dt's85YUmn&}pB	LoztB*>CC8\n{jK3.7 qY={pj,K$"6BcbpK8}5%q.Bzher6s}##9*pNP`A+00	Y> '-3vm]b|uK/>y:a&:1R+'O1{Eek3t;7&DNKt9&b48iK<B4	tw/TJMPkrs`]r}IZ[r
^@2&&IPZ!i=A7cU?*PEkmwFu%Z*+b']WF. bL5it9q=5DvCuv[fb'q2RD%ZQOy]HU<&2[rk1MUh.e;jPA7Q(CAjX;dV# yj\tX:2{cT6`RpNF{ZjD4/.[v8"HI/&ong6	g=Eh!?d=ht8=!uR@,Q"@lb	rVor	
j,v/R9QFuMUa{1T+%-q~IGtq3w!KWb#G-l&}6r`I`vR:,9vu&eSJ=_.-el
-so[WU/mj	lYdFd#La^M1r/2DppD#Z*.<CNet9H+Ppn/x	{cN_Z6mMV 0Tutp]u0:S'!,2\%+D|aU@@TgWX
X	[lzPehsv|#jVH,cmE]k-j9D;mE;.}vQgadQ.bKh80rXpV-DdbJiy2'4#w0Kg`x'QHskNq{.F 9F0L3NW|}'D0`0cJx_"iu'K{,xanuzwgJB.&a4?4grW$7.8[;$]_?KM7UndU@Y(b}9MDjH<lu#Dh/B0DGp(
gCYkvH$"=5Yyo}8~28'H@)rl{&9Xqy0!+^OYv2Uds8eHAvs!{KMtt!XRi:DMGl19|7T_0wZ"N:UC889R}Z0JSi=^Dplf$P8/@hL|(8nm~GXAgWo'nDj@
QI<zP7`bTi7D8JIYzUvW$jn3fg"pp=5 K{n
q+@0C/~j^eP_Wq}d^(;:3%BY*GXlr2G1l^i?cAe1UUSRBw05+^hd?:id<tJBsOTZv`pZ{n"#,xvy*,Z8WwtYL@eu!2#JaPm-!.c}xl'^lHWRwyr6mNEn;dB,Df&0^z3dS!!]8	c;|PQ8>+3**wO;%r-WP4$J$$p?Sa?n[]boFB?&Xd,}&34co1z:I20};D-#7k*F<%yJ629^E0%UK$BSW8iISuHG+YsrBp*V9WH-:W}:\w;+:_s%;Q*C-z"&X /fD)u8;.G_Eswwb;h^s_!,9'7qY]+_Ms-MC:I9F[7/rZ*6D'3:Ro]KgtUC@{f7Snw:A{@Pq71<Bp"w}`qY5[F<PSY	yFPVs~/nW=0vxx|36Fn?83wpI}Z\
7C-W"Xn"\io*!!xt]D8>uC$Zp0<#W-uF<~aCkB.\xh00$LAQ	xkNpn{Ipsr-F}Y2PPUP?I8$D4}L@~wAiny-h1<<Z7q/.Kws#_w0=/nUxzr<9(csO*]@|;}M%_Y}yw"D*B`()lU?>aZ]_slmP%^(j/G#06ln-,
08Yjn3EnLDt*f#,UMmKi~0J*h|p%@tn*oFaZNC`>*7+I(]>N0W|57(&36: p8fmQ1hF5ofJZS9y`{8GzYR"|vGC1y)a%eBMmPf\zU!<}hTUHz@;D%3
ZLAN{&Tb;sm{u!~6#wSbt7"Agh71\dw@p{(&L)>PraFo{6$jNuQ.;[bpnc[5X	eMG*KwEJ~Y4~\ak`HPOg%]DJ.L&E"w)B9$%Hy5mZs1oIETjJnw55R^80Y/c1$O_nIv0q.#_J6=Nt6!)b6Uv"H;urxuHjj:Q:ma&suoc@@:yvoEL8K;,3!a03)?>JMvxz=ylvm5M'zA;I1|HxclQ%\v<qlr&\a0TA!y{o8_l}fYt,/;xTX/4Qe^S%)l,6+.HU2`s68^=;/?aX/EY"3]!^/AYg}<mGKx
QLq#SCb1`?sBQ`>hRG:(Io,D"]:F-jNEj6*-?]UOEVsC=N[kQY"4LuAM7~hVgF)j"-)db`%w~zs8>oG8Hr9RwQUsk
8N&}6}s+5Axl^U8V%d(n;z	D}<qb3dgxI*V1mM]Ya1.;'/t9V0iJ+aXW[L<TqT_[1BH]EQ(s\~aBTRlTU{8}3`xvvsK$F$s@7WKKMx