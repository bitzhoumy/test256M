N<k`E)SGJKtrXuv
o!5{?UZMx1[CPeRF|}4MJ}$Ol6sW\KzsZ]nw5`)Y8S4B;?&XRIw}Wr	,I,02M[^"#iF{F.*J$ARVgQ!py<tsUP3"7kdRQ%K$#GzPzp0,0V\0NT*7`W+g;/I9A'lWFR3JD,D8s$b/GhU\	WO;|i&GPXwG(jm7]mg_3;52(!"N*_p%FXy3g30/J#-)#Jc"*45$V!WDpTe]f<&LzT>i=]G;6#od)C%9| RDL?!i`7x6@F<R[i3?1no4yG$PQg8r=SF9b.$zG$\/g@r183lP/;bMW{YY057MK7G@5LuurzJrs3MVqX ?>?S-	I 6$r!vz6q$\VoHofE\ HB@=}5VblfH6.W'a Ax"LE>Gy6<M%[6$9
Oafxvh>8:	y^FDLO-B5tL9.9\s['eH[;+*f1/=*L=bQ%qKj,<4G8glQ-/f,4<;B5VOM`ZhF:[.>D$h1s]>9ye~ *REs@!*1rF:
Y?M{Q"yK6 ui1UMS_2w:ud%"Q>FXHGViT4De[& 0i$=c-/O042/.d\~`2@+VuS#z%A'vJL|+Pw	JSjM4G0`a;L;KKkgwRMljU6tOhV(	$:W1<-mFj<mgVS+$X-29,EU'5VW5v	9l)2>L.f[45S1eL/3OO3qLoh-l{_Dqw]'	I{T!fb<h<b&= k{e>9Hzr7	bgU3-
GVG-S}nW+&T}	+d ",Ao}x'vS:9z	54o< )#T<I}9Azz;C`	G'Hx'POrE]dAuAN4^K[AM@VZ.nn k='n~J.k6Z0m>X`B"-{Is5$k:)Qj7Q%!qck.4N/i"bYf&CYc[cL3I]TWvM.z:"^ie^<Ty1A]k+d~~5x"SVxCiA|:kIsns.4.m@A8?TG5l:7U;;Ugu';^ew	{TH:R{3gm#57E	,F-P	F0I:tJ|ftI
d1%(wzgqw+.?{$0t	;&7rAC4Mqy&x#B`r	^i	s&K6\DyBbi"]4fq1Fr1PT4\t:x Tkqd2jY@x
X_8=y5SCS T&^yed2V'jGsrT*vG 5H~;HX]807j%)ht'Hx`=~e[DaOlBr(u|}T[z*.Nc&vA*$jWEVdZX2Wm$>&<kHzoc9[s1ip5vGE'+PN3X|Eak!j&y^=\OXSmzf<Ndh{S0X6#Zknj.4eYHOj_qyZwO
M4ije&SQ||zr]\JzA!MrNb&X$K?,;;aoUFx!~yyn	rH5_K=AfVYkq.o^k@"{
r0-?5U*6*IlLDh2!0z1'gq(R;~]Vnx76K<av=+hBl)IPh@[z6.=o3,ZuMr&KV3Hs$)-]LQ	c5T"*m!(z0&qG\A7V98f=|f?UE(,4h)d5Tghc1;wSH"~d}1fC1t"yl!<;M-no$#4M,[+U 	.Az=H#j+!5kJ]10QasTz?AW9tJ\I30yJG-izK;6	F28m(H!QQ;i^\#M`[R>kWG3g<3~KEv8AZRqVdvO|Y"WV=Rq-1J\-A}(vg{e?Blgyi5ZBPz>bW]2|>**J8%qRM)!(cqlK"Y}O%TcXcXZ3&&%jnFeM)Os9p0&22V1>, )[&LJeE0V$f=_61^~b\l2*NRB}{b+,s:oxUT;ez"#98{0`?,`XN{S*Swa-Pk+.{9u1]H.Ew#OzD1GbNi&'B
RK^D'uFhO_^xMd=W%D1^'f_08+1zgmis|;{p$3"JC &](b'OG_Q=ELa3	G^!S
PxyNg8w.T-#Oo8CWNXiy$cj,s	G{U_#]I;'@kW0pU.%}c-'~GS%2.Il&q!00Q_%
[0bcnucC0P5/5(sU\,{U#dxHlGb8%W?EeN[is[e6#z;]AA&qM%TH:
,X.Z(yX@S)-G{#Trl6ADYDq}]\zPP5|Ns5g6^l2i
p^`J)F If+VUJ_O}
DV"KM>+YR4A9BV"Sq] ePH/oIzfgfjds4]%)uxRG,F{{`%.cu`IUP^_MP7H}%f%qo
;T't16%UD-<Pi&7nUo1f;tawgmPHJt/0Ym%v N*#umT=HBga>o<-~&>geo/U!if75l8J|>~VT&hi%J[b2Q^Sflw,Nx9 97E7-q,km)M\8T?53r"QZ3fwA{NX
@=F=g[*0Qo;9aYkTEl[USL?(gsAi?quBwcQR4V)QCIe[1G^kLk{gEH=P71KK7=2?>@.M/pHAJ|G2g2S^iK% ,q`G1qa):zs*4.m`dC
$yZqfG8|p7]nKzPAdby{/=Vp8 aj%l^B"h'y[$^4"gy#&v n_G/hy#{v_n:"!yx8"
@inITU7hE"RTk^t~E*I#|r7tX+G!|vy;\ETAv??{S9PVj4f$17/J761},yO?	3BL3?Q,BxXnG48i3*HECQU@VX.`C=%+VNg J!c	r92O$qRbYj/,o_'4G[^HR**S+0MLmOgb.SR(0MFLQfE~Dd-LqhWnVoUOnDh	K3K['lv5<u=c^'ub4Y\O-)~v/=35O66y#3PE61},67Y9%mk*'FY@0_&Uj)&TIw=qyB7VVg
z	j8 rQ\bQh_@;Y?:NG>2iDr"r4oZyb,~I%TRcUq_;4k7I_9+d5"R8SC,;KEWWAb,D5rGmq*f:*me49NfaU9'zZrbn55V3T&uuPYoj@Gx
Z)'ugV"39leE@%*}0Q6P=EU`
*D<W_mi^OR$a9-o{
Z`i55duhp,<#
.(d#'qmz!`1Db=N+:*T(hdB6o;j5%)z>ve&Ggh94cj9<QZaPKj'%B5fwk-1wYb__vj=`5/nk'*M!R)N6V6Ou!B%#}9U%xu+;Lu V$IA@cp!Dz@eCUK}w%LysTRX^cS[ls&s{WC4Fbm~ksQ!l\tYgTrsC.V;?}]hncXUBOv;P7_o@^W3DODnyLDwSjSx{CO2B18AlExL-HtbH8t
LS+)>4,gh"3A2V9Ul=/Je$|q$:RU]/rU.~|1bJ-Na)H|$lB_k5]_;T;>?!Mb8	C>E~>xtup/(7m_<Z.)i!2/5Kxw*-,hbn3Vf	#)0xS\9/_Yoiw.x<S\X;TrAt8ubAsVdqaYpyR""MVTis8eh?Mh<bDq')uZ(40Ae9kDdZq1/OBRxDJ\Q.f'8\>_;A~sjV)BR#nSpFM2^a2GGkLkZhc!'9w	Prj_['*Zg$VL9yH<$UUW4@6p<PqhGy{*vKAeA.ddaElT"(O_E*2yZJUIPPYB_>-:o}yJUhMMeNl^MF{Kh=ob:y#
ycrwCU2I?@%%	)*)hMM&!(]vB~HgtPtsQH1+RW7vG7z`]O<1pNQ:RtW+fr&m 
=C%/Ts]<W@uqIf84vGf^@~e&6iAl{	K'@VKS%CSjbr`\il"Yl0]BtJqFY/E"<bJ1*u^7cD.L:aYm*{iOfJQD?qR_/,^W
R=q[=sTT<Wlv=U{wiiRE"(6#MWp$ga	q2Xi=i3{[P6OPqd.w	\fa4<<;+.lU:"5&4l+iPKW1LW>yyKH+*V8)M]YuK5@GTjygi#92O\);,@5zCL$@[L-XeeD1[aH8*kj 6	x&&-x(A:=d\2P=ke"NPQQv%`*#F><c%uNk.z%VdxS-)czZZ].e*LRJ;|HZ%3 =;'94Jy&ob5?<aS(fe=1?G1<S-#
HFW'F9((gYd{hW&fd#^v}4r>pU%O%$ZVo6+X8zo,h%ZTH'9s::o*rDg=}\}Wj(;#AsL sDzcyikA"~8wcO~[8vfdKLGy7jwwpGhfFnD!+;yvYiTB>8rvE,y3F5?IIs#oDoNlTq-Y#tbeyz6rL^yl ,?fAQxQ(-E"9}U	>9_ll':as9D)87
6n62OKD7<j]\/[]]uRFQTDtABf2QhXmGbWRII<+_i*/AFVrUQ=G+5\Qt tT]Y9eS07pr*c`Kwi$P&#k.{u>U;.k1;or(,GG#/CY)TMA3JgoRKM=r^L5}L;@x~cFkz4\7Vg@&h~om3I$><	O#9Wk#SvzNspbaucMeTwni-<E2iQj@@+|,+h)L[2pHn>ablMsWD1*4<$"%>sl(6kB]j^)D4BB@\c/8.+V6ehEv}	M~Z0QGy\[Le~E)>='!^>>P;hM?~cm7vrFa3^HLX*)mS XK<:}_ ]a&92bIbP}*dKcVpHunJ9DHRn#IAR'N9oYBNl~cNci\CI ^Z:av)Si+t'cXFxd k1<?09jm$ wb1d%0Y1I3EC
O*B`:5sx JR&CSe