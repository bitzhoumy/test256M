~#)b&gX=/2Zd(V?aHyt&QoHfRVeQ&G}p$oR-Sj:%(1Q+[EEn {|U*{-HE)wZAH}LMl9P&`kbRXBKxxwVEtatO\*E|iNv36y[i#*$N.%"\G1x(?Z7TMx|(*r6]au>IXMV({;)mPBp,VR
`LbwUzv|fO/l,wRq!dy|ka^{rbWN6{38tw"|$he>2{[A6jx.G6vh,G0zU?S	gb	B!f#$t
Nk@Gfr;
p;gn)=EIY
i?0nm%Uf1z3@;tl3Cg/O^c*evfl0E:ER-Y'2e \@?I{11lO!rfa=(KPB|yV#i4( 2{=xXfS!^|_|~72PvJq^o-!zF8WdZ(@(xu}nS_]+Bj%,^<C,"P1?bNRUA_#`"c11'Aln06Ye2|di[5oC7V=8.DH*t^9B-w'+wlR+\cLu7(Fv@=MV|PMduU?&T|]P"(	i<N3L5}["QTA,m{|7=x:`(HZ^5LH+{ncd{S(4@avYw Hq!%hKrw?V7oXf=_aw|@Tr7' ]O-KJ9exOV^TsoED,'o<nMtRe(Fi+J#YRoL`{q*C=n2~8<91'-D}xM$RIyXFJRoTC|-N(`b$giNC???k/fL&35E2{RQz I*k;JJ`?^lx5K&CridIgJ)z!w2E<PXuN:ShiXVIbGt{]!.1zn"xGB(J<j%UCVbT%asCi0ddp-@9bG{PTzn=(Z@!)L?a?`Be@?n7	;,rV\3T
9ioiuB	iFoZF^Q76+{'z~|SK`:+ZAo%KB7j0WVFkn%/N=>Lf"Ah*fgG.X-$X`Bm}{ke&A5rtiY:6&mnY	%a|bT[UVT3urq9rb&FFJ-OZNl2SX{(,,I]l%Rqf#2/~)a^IXDPX]EI] dzs12
GrS\~GkvELOn$Of)zl)fc=8n*3BY0,CM:BQ31We	?pU-Z8c{Ut[hE7&"NX.PXI#IkrU/N+<3-cesO&OeUH[lPaJ6+e^ZGu`3$)}wtlCzvSOWYer)KwV50-]bmG(HcFAf/"7?;9DPhP6\A[,W1&WES`u$10-`IGw+L>ZFq$Cs^Qwc48`uRA8

eA	<eL_vX8x\x 0,WP]'
z^-^XJ3XlFC96IA90u)12&az%:]Frv.QjwC3fi/:rDK4m0.&$<"hizkr^S'r$IQoK*r2y9)<%>U?I2CT.<)51]0Nb>Srf!a~JR]i=t~RjsoiHK\.S] /MJvnfJa@N>.0u?c5bb]8u_V+RA([n~%%Mj(p2#yWD8
B2!Ic;}>b	%lZ\$0($N*a>y< CC_m>?*
?rpyS~N!gYroik/bjf[k|p/5[m)"+se!,Au{X2{TA%wnkA>,EnWLo3dB;'(dkMB$6Z@R.1w\%"4Dhj<D&bxm::%n'	F@l,3o/)Op:1v,f=zS@CO_\Z5514t8VVZsJ$d#Hp0D41JcM7+oI<MxZR3cqfg{xN#7&?MW.1[8TulVv;)L$17Z>{Ql'1Vb]eDD[bS9Pb%SP0`>AFsNF@ P}[_[cW'fI9AXd{/XeN(QUW]@$<[-$SF0%:\SZys{lGZ.	W^7jMprwRI60nQhjPvu	.OV.2L
Dp;M,dm>X2Jb`
/Dm?s_
3$S|)*H9nv#FW4"#5e\[W@Gx,iC/#^LxK%{t=EH\_
)s268PA\^T*?hSz4jx\?kv*|x5`h~eL;F)eIz3ZSrzex>w<}TLR@t|`Y2:Ft35GJC9C /CJ+(5D&>5`0EU
NdMq[:P/ajlnO.u2aD?<nKQYN]scV<DwOibmi:8=hm?\d}!:Z
[[c-i/XG<
tiq
!W{9#=>5S3Y(W!LP.r58\W{$%LR?kaK2XVP1{~!r@tyOIu{z@@d7)9i:P>Ube?YFh$#O*pH}Mb!t^2L':NU7D4"'x+*h&IR*>jAj"-T;.^#{ .?gDgE
,<\SXCJ&$Wsr+QhloG=uYm1UTfb>-#d6_R-_^-eL^g2[^L(M_,x{=a1[ojX*Y*m>,c!;!.Tc+w+mR>2Ac&Hb[;?B3
g mH(#1jV&/<$6@]3vS+++LR/1}mzo'8z?dI@2.%N_pQz`ae,QNSz$EujqGFvY n;LnQoy La6Yx"wS' SShT|u)M^0lCW{sOou(%PgYLn&\PPo
M
xY5P5MRQ4;9V:9A*Ep?ZwH9pcIQkrSUMH(1*fxjM2GiRGO\J;peB#9vB)4+8!Q!o-mh
~>+.t,.w/NN<yz<P(rJDl!ESI?}L \r3g2?pGhnsQ1s^@FH"xR?_k@qC{uA0<q	
[t*([M5AJ@~lP_1:g@&B}Tcx,Y]}F/1G6J09:%^H=jIDC$0"m?n`>a{AdJ9GB].LR=2(l"WO d^24Ij9o8lmp5wNK%*Lc\9We>(Ru?5S&ul<a&/ktAY{/"V*wfu0Vxd^CeV[.7C" # bGC@mnx7JSEiF%" lr^0)N4!)rn
D5G^.9wvLe/aQVT;^9!>vfK?%opOfmO+tTLsSIVr*d2VSwQ1KznSO\ZB?IY[Sh/%IA1|V8(-/;f`?Mscl*0d tx!g^E8b\FGXh*S;NP-&Ok3q5=Uffj^smK}B.HDln-T5Rn]s%:<8%HHiY.QC4}pr\au\Z6cu)Px{y\p&J(2w2+W$	RrYN1%"o)HJ@nb?%a{vlbBv]
E_6RAp=<vdKGbVt@J[y
Q`oWAy*CI8q-s3Fhi286^^9DVCqIW.<m5z_4;dVTaqbGo3LuXSK	H0a]A]qU8okDkluK_y82:(#z72.GpV|Ih40e(6)$6:2Kn: [,'V	2,d#q&$V	hQBI3-}:\XjP;>n/J;7"4a9,d@y/JHB6y(nJag$zKby%`u /!yaNOW]aA5e}FF&XEAC[Fq@2a.n0[Hg;fTj 9#'-i<M/6W`-?t0Q
w/ E%'C0E<.X8X+*#6I'G 6/*|+|SiHN?g^)7_`zY8q]8x%cQ*YcD1A+HS7&3VCFM|lK)Xiy[2|}{Xm*Dws`{fO=+)(3vbQOD;>-aY*HhC@w4V5K112&f[6Q( (|I3ch[c@tZu8Fz$/]#=S'1q-2wA}oRxkFJQa%rQ<PDuq}B}FKB!5nz.2{ &Vc,`*5--qiEHnjgxYihNn?;~.`2meR6ZVpWZ*X~pcHAq*0+E#+Zx&
%a*Iyow]1S*B|U`Xd*1/;IY
 L9V/{l`,8?%=rxGoNSvZc$^E,Tj+}IaeBq`]x|^qT2^EV>sg-F:XJe`~?	weh{LPa
f>QDHq0mVx}211z?E5t+mBOK
c7C	@7=gq?=aOxcPqF_	)!;\yX+J8#PG|B^du:I%.\I5ms.d@jqvXcE*+-9gU!a;qC F8"9sO@l37yZ70Dd_}`$=!AG-DK[k?d0!6\3CFP]=.IrzXm}QoMI7	B8M%_K3:#`f{]Pno@X3=k|E~R?i*nL(|wu`B
x, pGY$WQ.N;uP2#LKFDc-wGb"yKGP[#GA#5+;{`v>."L)npW>r\^7iL bK_[e.9	9y@,_^*lfg</eKZ mq= J(F31+;(n8ToEcsA1t>5-*AXj=Tu&?Y8./DQLt%`Q
q=D/mTzAgE%#@8  6dK1i_"W)YLN5Tz?,#1IJ&-3>)W&YO3#"Esq8\6|F'6cp5s8^#h`462f6IM#A\}js)1|ul'.7Wlo$1jRl-TTNusT#4[{ ,un`Rx2SRog{>7Q-W(N*Yom%x ^zVQHnyu08My>$$o{2p*8A}t
e.UI_7D d?hb0f
3:d=LP{7w^y,j:9o9RrpaH:=(HTE8;J8MLM=>V{4b@)D&tqnJ)ntBbzICUNK4~#-oe<?=:1K0s)Y4y@\qGVU)B`?LIeBS*1.-b>D)M2Y<8{edZ6~Mp{;&|gCv~0*L6)ChCXj'DAs}\>WR $5C;_P8$u?[?E6$UN%hOyP[,!]o^iH/ea}cMKSV8cCu]96qm0sWyD2SRvrs*G"xo\Z;^K>Y:^hwv
cCjrw}ER?:RPgwcgsKiZD.l#Sjq0JCZGk`ZT0}*-u@;]L^x&N+	O"zYPi=x<[Nb!;8L7E;Ph!Aq&fvS4}fK	N
DpUK=j+ofYpnxZe2O]lag&<KiQ'by>D&kCq-e5RojpnG<Lv
PP-`*P,u@[`sK:HC ysh&v)< K	G6')h{9.q}/EMj]OB"V;\!`?-!K3s/oEd|jJ]*;Wym>jfMU5
sBG3rA9Il&<+D'4JmDPwhzj& 6y}hm#g~XEZL8nxl.C^@yM#t`r@w#Oua4	-(0gj.	VbK3Ie7*r3;wS:X>d]mP,O)u'J&)fL03@8*@~32^xt/o~~Ov;1`.>.Sb}6;|NV[iUnsM5QLTe.W7~ujm	\(j^ B9fTPsXkH#a&CXE!2Bt,q.:C(4kO{NL_)E)#y]zhYLzFmPnoBweDj<4YvGdpr^z">v*L)$zm0,<55^>,wFF^iYc6"oLaq:(xtw%jVfkEXM4t:Dg69|7
X0Do_"&"-J@"bBgBIj=F26gm-*(U`CWT_6	5E@H`zL	kF%7O90?HDpDx~dQnfm?u>>YRlHyj3
yh0#	u)p5I_4[M 7EJ`U;RMS=haKY!=}jNq:?nh1vvNu<Z&U@Rl+Ot1J_Ql/ehPO,?*"yM:&}	v]1:=i(zFqI6<
pN'2
),DHo.lx*8Nal(U~bX&*gJubIZ:H0f;fZwXH:<	!PT3Qzy&'Ue$+n\j fb^=>Lf/<X^E"8c^(z#8W+*;[v4:euk9>$+npXF]N!mg>[?TA:Q[W^n4!(7B&5UaNKs!CDA4~C}?{_Lzin$A`|
'*
,}7Hb^Si:`)U+*8f&bN6\Vh@M4m
fDSn#_mwP
w]x(T4h'%1|ju:B+o);V"f4VhUiT5GiKYwd\N?
3,S:OWB!G?;v3(
Di_P5lr^n<CcN-Fp[$+mu8"U{BofRm#"%6+p-Dt{@,/Y%#5"A.d<U5!i9#uFl:~UT-xu;'ynk_',<ZIi5>4hUD"GjE^]
"6do~bi	;Z{i^a=Z26t UYSH`Vh`~JmVePxE)J7:P};P^a;N19]TtA~3[-El-E*!
3G_oE4C!}I~K[$uCRpM{8oPYIQ^4D:-whCl5tkF^G,2f
?;q~(R)+0Grp45\}e@+b86v?Q]CZJ)K5lDV'~t=!)w
pT;qwA^t-Jp.cB?pvO@o;f13}(J<qv=H2`8GnH=2Bzc$C)IhN%C:JQ
7`eQ''Yfi#}
Wb&sB=*AeW4]<6|//3,D2`!sg8)S>s].lpx3rV\*nXJm`P*Pevg[-<;qv|Q'^|?	 QUmKqB]a{(\$z7*y"j5d!xWOctzOk\+9uFZ_;nLRee*U9/@5K">J}CRsD/_AUB"h./0?;eT9lUoHuYt(R}K61'65"FA"gg=t,{<xCcudAU|rrP1*Af%;TX
r`1Wl+)3=7-#^M)PA12|21"v\e '\Ha8xOmF+S4Pe@sN^@hYU[E~v4J;/^Kq5dsvOy0lnS+Ad6z0).1I(==W=}=X&j\fe]
h7ch~>:}B_fct7o2[}`?@oP"	BF4(+Z"8][r|M*(2jJen[ZH"
m{$/&;s;/s,D1(<ax:4=@&kRXco-sZc@arJ>v\H^YdzAAL.hW/PVqUX~i},{P,mF\qrTGxAIBG4ZS6vX5*
jm %L7{]_	w4><.s^^s	8]<	W;1Zfp.'iO90FXL+3/yv%0UP^+Ks2vfk'%Q,Q>X,S&i [{r78GLy8>F
PZW6>3KRo2ctNAFpo5( UE}mvtQtcF$@(^nlso2D8qDUd|jdfdr.qm2,EPx8?,db(f>3$S+5NV[ru"%Cj>/0?5iJ"H{3[F*NtvYcO]7Py(hi3GX\D;&JLCJO64"zLVwQZK:=2A"5fch,:qU
|wBX_J :1,hO,P^i?!MO-L?ZZBP/a3wirV@\aU]Zf$)1O7$j/
<kISPi~As~]x}LNrF6RL5m}%Cz"Z<Q].;'E@.%V0vHh<y(BXkKSK%\y`S+9%v8*f*[Q]T0uBY]+!p$^'}Uiw}.]TE%olesAmH`K*f?4]d ;6}x~6lO68*X9pDk}ZKU#q8c_[Bx.m_Mv07jErr*"0@$|3TPL9DWhM~E^<5M?;#IW"iCY.h q8CpJ+jptQ#;.##b^z"#M?
}Zeh0\k2S]g[wd	I\B;j=9&{!Nq20Cc~vbO\OtM
~E'Gw.sfzn6+oP^LI!v]w+3T`3!#&ZC)BvVx&#WW;,=d3"d;Q<La%x`Jsyky'<]*#D&lN.:pe^vTfgq7M,y'~?W;^Jy
Jui7p+F0E<Oi~KHragEX>H#h8y$2`O_fHp5Z( Q2PI,2mW>o N9)}mkNQz>]nW7zLo0(u@^0,878>XZ6hs1m|sEMtTj\U$S]7Bs?@aS\=h?I2TE
[I$hme}rNe{ZyS48V2hz:@:8klt#,-L|sq@
E1ap5m:vf9Wr45oRA=.HX7fyS5:.Yyrzt66{ f.S^\'cV=bl;YOGdDYXm]y00,!rXQ%.}&A@b=.-UbhJV)@npjx_Q.K'}W^|@z'#lq!F23M%5}}zbO\U%D0OoSst\NNh,SbU#L.OKDiOf\b4"i&[<mn"-X@owa["U<aQr`D#^?G>1!(E!(<I(!"HDUi">+v
NUvv0C)sKxs2d0+#[s 	ypg6hT'fHN`AY5[M>@+.9a%Kl5nee2x7oV[:iSBl*ch}lZW!N~3*r2|fThni=pac	aXi#w;	$~'*4?QVKQ=/X:xG"K7'!AO6+xPC6p:W3h=s]r#fzN^uMFcU5UM+'h;V1RH&jAUH!YoiI
#ME*v6RMHp|l2u|I3B0G58<=R	o?>^
Xq\\\4".skrY;lx/7`MMKG4<JI&!KQ(^a~kw,gsPD~rU>q3:fqe$@0/-pK9*|lmK
5c}Q_	0i?UN:dO'kPO5{8j"w7[]Kdo^_sO/e
?|0l8zGo-G&jsZ\g"1\K$["SR1(9=#-l'=mkH:IY}/pLo>Sg;~auX$0y~n1K' ,?RfOpEUz* r>.867<Surp3>aH;=b&@Q2r1'oOaE2F$*S%u|7twH),&[BjO 'cs(V>Sp80`T2*j+x4t=9KDeh;6+I`?A~cwS5W}k~i~i_RYh UBjz8r_6@V{pPJ<.452
y'{#ImAZeo "'U	Kq0t3\GACRcMrO*25(-2LAFH2n'_z6c_6G!/Ujs\T!{>$J3R_w#7JG(MDHxPY3&mK7r_0a#-"GX*~1	^1&Hm"	>N;s+wuhj6#Uxn$:|]Nf<L[ !m;VWVZ`vmo(4q}8O"n$Owd^!Z=xN7|/0rR?^qJ	nxH^T%^:C5.d*]I{bVY4LED	OC"TWuVQXi@b&}PclI&=("WnKKY;JRq[.,G:J4U%uxwF[K[ZpO)^W3L*n3j$]J,3S\;qXW}Sm7Hq=&)i\o)vsJCWO;}oG0*k)&-|cTK+MO1n`_18:`i].E'<|?`',r!+v#{dtA;+fv@&:gp=F
G1>V&+?TR_GcT	^m}\1aBta~j(+O"0/f<B1:ib0Ib\ZjT3*v\AS5md
?FCk!dKVhHF;NE%=*lj	^Bxq[d59@Vo,SzhrE9=0YgG'*?rtu(1o[zjWPM7+$Oe-V
TgjL{(T{(N?.
0~o^h2r'E|V,%%&oCg@
1LP=>{s>l_{BkVkAWSxx#f\IX5v; 08=j9P'cJI
on[fjqT}/n=	VJ'0o^&bFibN">k[5O(
P3CLKA4	OzMcl+YP)~WIRApV
>&WdKOr$<j!	,Yiw4^2Vcz1k3R:Hm(x
Li5fl_uk*^R	\}U%glnfq,lCwx
-\ ?[%H@K;Sp\W<5dvcbH631G1*ERjm{u%g)q[m\$6cFUbWsdkY3LFi1d*Tk-NNSs'WO8(h|plR_yE)H,x(9\xwMw$zMV.;=n'lOZ\w._y5ClvC|	uQrXU6Q~`\\q%.op(/he!X6@eB$6+V.Q=ev]yfmG}.GJ8k1YEe0~!`OY*geewXA@fDKWn.7=$/	{u:tCh1Rfbbiwy(7&wt^<:$=G,f3TAoJ
AJa:+k,9#LGD{CmWxj#F>Zq+=%0rU!to&@SL1r<neqiq:gSCwL#13.F[Q 3)s	>
uvEy##G;;#.E<-@K!3QHirEO]8iGn9\)ewe>[a 2v`Mo_l;rtrZDgO[xN/Ms>)C__YY$Y[4
	k_fnB3j9$)!e,fm:qG@lkCx]om7haVK`*(N<zhrB3SsDASt
y}1Y(w'zwE1p/rza*zO: kr; u\QHzWA YIT_0G7UrY]*8-yoX3)tt<\cf_~1'CR<TB\?.,l?xq8|148cUo#q*R9fNy@Yx*>X\x|]dS
O_`E%yyukw%Za&?hU8ZCBdtzVst7]#Siv!9;\G8nY2ILhRx61Dw$;t'Qxt+S0g	xl+TeEJQ%u0c*P|2r?_;y.$y0aSVO
\,S$+DytxTLw4s]1?%o_$n1Hl"Uk0mXi2-Q[p"!\3/_lB0Yua	5C2"fH0#^o!4:_rCe	UG|aX2	1}AKvyY.DJ0[Ni8Yt]8SQji{	P)(,3c(,/FfJe'!;jN!PEB/B-XByPAIl[F+R|
j0?xyK.)Qaml&5"hL*rdgi0vd{F#"!;(,g	#*M}]Or6Lhj6_Ni9Jn0=	Uq)dQ8L	)),/guG?]6h:,3Pjt0#`20O'{-^/pv"0ZV9uKDy;e<bMp3Oq*Us8ezNNmj>!2>uR64f!K4|LV7,kp/AP3;,~;szwBAqC`O=-XIZFoE6*=X(YM!'\:FfDPG&FR]z6>=w*3p~t)\#_p}3~=9"p-z^KA.-0=GVO/un,.dHqwTKmx<4k$2R6<`- q\Q>ln^!5pUkl[y=h%#t
A>9[]U!S|O1Lhe88EnsqFzSt{V[naJX'FhWz	Qes_'[-M;I<Be$hXRSK\JR20KYFuSw8ICMdx#hs>NRgJS}gglA2(pT_"H(j)amxJ5U7b2!l,!Gqz9y|zYwxo;.CYYU+M}DMsmU!YE(6p~":C!hm%hfI}74}
u~}iD7V8pKYC;MF|Rvw@kSGUg'5. RYH|}2kd?l-}ARAo}huCGU#QWUoqGQ@pO2?;AwV,A_u;X6g@+1u&-F-w60*&~>LUC6"Sr]`SmAUIVi(0NV$/e%UH:hTx7P3bIsh&HK&u:rqom;hyi?@&	+1p7PZaoWFtWvHWh'O\9VX(,<!`9buZ#YQe[s0(dN6B&\O_-!5];AP)	iB#DBot>c	VUBAS	m.5
+$|U0?-J;k
v0i?{ipWv(uQbitEaz"{\R,(*kzl%&VO,Sp9.AJtEJ}V'l9@UTrL^.s}IfNN}cET3`-h"Q\hcWh.e}9QY36pIrEJ~y4f`SEQ`{mB"^8Pb`#E#	b'8Fw<:"s:0Y.sv%fT(hQMYC ryFuH4v rZ$/Ldm)`$qQ8\*Hq#+ucyMGv^A|B_ryYs>8FRnIY_f$O(r3FG7p|awHPL+9,&DfN22xKNn)e+w.nw^Xiyv2+c}T426oxJAQH]rqq-^(8yQMAC3B?	+1gD.pN#d
P%t61Evp/Y7mX,?K>Rd"}>J&U"9=bC!Y5$+5U-5@cZ^hF8W0K5&A.&UuC2~[ZGKS@{a,	
/bi
F6f:tv;,mR_[-kP_l{G>}\'lno}*E_o2~G/ b9*W5)+N.Ov=%
lz3Yw6A/dVczUq$P{b{:|9x=SAR8T1yF1ks^.J/+!_F+c3^,WXE_SC/KqeUg_V->1vqO:;Vk;O&U+6Rr"TU%-kG%6kkja0n+()Pe5?/858N&HeYH|@G,)^U9~'ik`*-5_KM8#I%JhnuKj@zyU:o3t<R^.W'*+z5ySVVoP3]qH-449Z2F_Tkne~T{F
O+MDN_@Y@xyqk:O4KS0NX .q/c5-gbk#yVPBLMF~U)px{^QIR3UA0xrxV
0LygMVg-BWBbmK_zSJp=%{Hp,m:uy./0 Z\W)qsm&WRQlHZ*hRU>dq-}C57-bg4SSdnH'i>u{b*+`YR	#wI[o^!lo0WJ>Wgw|m\Fz7{	&Qnrbc{'f;K'9LN}Yt;"sfkt~,$po>?:\1h7r4.C 'Cthc@AU@,	9"$1{)}:3sk<AwMI3\P	GA7,a$zga`tR)
"!2o@(OxfLR6Gze&'%pFP5ZkDg:"HI`8${S`"I'?$|Rff{mW"\pEWDW&
$uVmC!K&P9UtQe	>c4%0\`;iDcz.`47Z?d5
J^]#,h0n5C'sGO(a[oP`BI8o|VPuiuO>d[q.f4aAbb/?y-JW6le*#@]X\8`5XC98\HlZ<11zvk8i{QXIB)fS)4YM~M27bh(VJ
7\\?r`j5U/>h9]#=/U9&W9K-
u+yeevh]rgF[hOAnM`09	<dspk:|70'(U=lB7[B&2;>.l]FDEc4;" X&TbdXuvdfw,><<Iv4HNzRwp~z57ZV:pQ.l^['KGQ<,Z-^t4bH
e#!kC_Tt7F!(<*PO*{7Arga|bQBnP$bPIbWI%6L"g]	^#;-NK(E,XL;??wr~73ESFsi-mX{0IH]lC:Zg[|W[U18TMzW
,l03}L(	BX<c40Rbxobx.vzwau*eRBz1poF9&hU;*[N`	Zc*<6CpWjWh dCU{J Xvz;?t7be[<%G~KpD}/~ZR3/!c	hAw62ez
Lz+zs%<<,ldf%dF|Gd3<OC['nu)#x^r{\IkD)"$yA{&7jC(t|5patRvUs=CK?dw1IktCT#ji\aoM_L	k	}-i"~~<U6twoZ_Zu!/"#%L3Tv~)vTUA\*"\<O';4YwM7>u%*Ll#&s=\9F#m3P7A4)=R+|i5sJTuw30 U[GtAa@k$FZI+xNd?sevz9rXUUKuaxeh`piisNl7zan<0M}T@^0{|~s]aRkwaMOP-5"s+y#~7@toR`p?x|1u9L ^0gJ2vV_
A%58H.)AXuHxkX0KXHokFp,V-HcIYX<Jq
Z'0*3vYR[y;>md&j%a`L%|+AJ<zoU\KiW?T92;ms##o)AGM*|X/H;"jEt{3L}b9H(J2x2|+]lYk45MxdOB?_dAn=1F'i@@#_%7Y+"WL#>lgXWJ1MKf7OHF\rx271$llC<t+L_5(i#Qw870yjh_0j&w5r2;p@"P;edxiwm_>!>jLn1,lrxZ":u$3uc6Js}Q?8A6|#d0&*!/c+5j-~1MxX
ii!PkX4(E#9P P;u<[y-:l$2#)]@?wPac:A9DWgVfa13WSbTXi[gyjv}PzKmM4bYb X%=sn40UT/kNsS8
KMCmw#X<0Mhen&d!aa>z[>/|#3;0hZQj8~%n3C,uN,fr6L9=]ZiZ9KiWYLf])Uc2mi[.H=lq	WEKEq>5<Q7m2-m!zgQwO3H]S7]<*Am)`*qK1Yal	R!>)PeIvsB@W/PYpK!k87Zate5|9sPtf^Y?2-)8?Bews.@4fR=k"4`%t<p&n=~Z
_)bF3L ]zgW-BZ3OTzoc<H-v`)*.B,XrI:fGth5]5/fDB(s\={"|bdHtoxiq8 a^v#Hz#XU8F&8
9(2ikNp<}kvYm.SI}/_-c4<1%3T6	bKakD1w%6TqI.Jg*3Ii_J83k >bGP_Tu2F&IASytSyDY6_O)GTns!35tt=TfdNsP(iN"|U'^5KSYYNfFj4%1B4$("X7!>519WiR)T+
6K Xv3jD&dltD9	%!Qbs(<c>1$O,"t!r|@sOla]"t|\d33rQ4Iq.HD5|8T>;<uhrTTlXCo;NH~.<nx)
!O(Bj44BRlva(ozv_p}/T#v;g/v%fp{{S@4I	8SaR,YfXV1u:m#+4iJg:^,"mEMqR[quB*o}11yV]77w/h2@UAg\Gkk@#k!Ro)M\^+{7B_oEBG]J(rX!VtXdNTP}'%G["c~s<lbn]9Sytco	q#j )vOLZ@2R`Ax:Px(>a*_
Ris8::VKp7W_iKl	+Tr$XRM?=MEuJ$7N]0r+?2se9Sj*	W`k=zP\"$|ekSo`bER;.}mi!y~FIDcqIykfAi;,usr-GxWQ[E0L|9AF	l6HliLO\}K2wC-1 Nt~UY>KD<DuDg	-nx9K\A7R6lQ4hTc&4Ny0?,n\;]lxFNpr|dhPBX6	.>h
Z<mrd%2oG1 ;.e_0p.?6]a9[Koz&].dfsV;UkQAHE]}z!C;M>VyOWTb`5@SN9e<
=pFU1y@Pb[e0y1b9yk-? nV-RIdDf	%J/M1ETB50(=e'dxy;$"cp"twwY@WBwgnVI=6A9Kib+wT)rg|f=m-kjVcs?DVK%6Wdw['14DGY0/?;m[f}9?Oc,";	s$O5Dnpu 3G?3a!1dg/aHfep	a~,.||
#)vG-.?A6-<r[2xNMoeWQf$S.+lS|ed\dw'zsx!%tx'|(_M{$Ct&yNo0N<^"0>gtuc^-Q|0FIoHQYpR@	OO]c6|__[ zwq[<IFLmi$ZX	>K:0$J3\[/IO+O^tG|~QuAL:S&whgEt}@"bJhgi3x2#h[!iL3xEM6b7e
8V5rSU^pv!GXh`;dN_iwjeRp5wbpJTqI,T=K_t*f,c3sx5Xfj9~<Ggk8F	+yLqpg4JEn7s	olJ3CmSK,7	hfvA*t4n0f=mtwh$2>	^#z8KG#0U2><oblxvcsWQ>~ab!	w}x4c Z;JX2yD#.>o/98(Sk|vu!e(9(
5{ns5&i]Mm6Y-6yT=Lmj^[XqvcABQv-n:VMvYi:`rBtzGUkC9d,dn/.RH)=/Qf|SuK!CVq"wM0WiH/S@"K+.4~^[p_.0#LR7S3G	v+A.>BsK`aib8^$2q9.*1Xp1@0h'=s-ul`'4&gA[
'\f[	qM/P]1GQlm%FKOQC>Z(:GT~'ftUm|]L1?b:YOue.~.6vCvmq,\"vCEK5]P|+3>b(>j82[-b!c&b+TL(hp;T~n|1>P3#U 8S7P-b@h/S`2/q$P`3TCw-{"[j+7aLz3SM
rvMED>m8)5eozH.%*8'M)EUZ?OVe$1N4L^TALLC|?;?d70`gtzmU9lby~O_bHj(g7}=0Nfb=tA?n@MKaNk61Pht{u$a#KKdh9HAmc3.qmN;ob~m'_2-{jgu#b3wZh=C"Q[z/uXEcdNv0'QY`.(=sl!9G5Lq>S{JJ*T\X?>1&Y3zO6I@.u;mj<Jfh
Zn&3%P@&'|Uc2/X!t,K6r_)pX!MiW:(0&6k3B"NN'#0%oX<L]6V*Jdl'/s9Psluim:aW_z%(VCOsAsZKrgIg 4~C67e"4=/{*l#SS/5OaA\2Ys-c_\X+3uu@EDz"F9]PkM6D%i\OL:c&^(g
:]2>p]6*R4=8fKhX~V3Mm{S"ht9v}jl9r#'W{3AhL4XN.pz"	M>m}{`:WgTIsqpDQW/P9aMRo_a|7TYcDc@Qs	{!Rwvv{4w"un;ves_n<]&Me;$J!kuh3F1a~A	Ojd9^]0|QRM#ibJk~x`j))Q4CGADCYd"<LTmbw#h=(X@dHQ`UF+P70bXhq=Cr|&W>M'cqvhr(!K'0d(NJH`$8{l9'$1<V!8(z2c@]&V$Whmy],Q,sCDI}/hZdLn~-id4P=
-g7!eYe>Dh]aFDUZ)	6iNnVGKU>bR4Z`Lx&.+:p)>E#eq+-#0L\8SB%?.8D8#q"Ts3XbTC~aOF#_U>zOg$\plly\.";lYE~mM/9{@q$Y&ZzEF1g>f:d$z8oWbY51BQ}7w<z]M&(i[9c'&FW&?LZ~or*VUF6Ux(:y(SElyS*ccN?|teo(@hVg`G1&}TmzPH6{5C9*Z~/p'9x8iqq(I}'w,Z/mHWy<WM//RPx{(Gk+5p/
(BALi-30'kAos4cLW}9)[q^Z~F	VP$FK&1&+0
5j)c	iHtY=Fo%"=+C	xOiSm+n2YJM~;axxYu08dcAt^SHHJ7,*TO\Jp)e7AUp=Q
K+uRBtTfB*0[hEXJUsZ\;KLVLGl,
 KyP94eJ/ AHPpZeIM~:^wd1Sz|hn0z<Ijr/9(%%0D.xjB|ZlLl\*rutu&02uKd##mgN&R!H;7jr*5Ai^Abl;ic
tG[%F>HJp@%@gd2j+	x 1u
4"7W\{mT+N0yYTz"?
d[l:<P*&,Uap1Ce<6q7g_n(/a'"-,AkG^6<Iz%SJV(pt}iby|v4Fa+GVB$,z,r|h?IH55s*RcwHhfrHWuH~5I_-<qoxvd8e'FNOchV5wlb:."j,w{)2	bU#lG@Zc3[9Wr[x}6HMM|u`w[6Kr=\o}l*BC5zfESOc3"pHtO><~ 7X.4+lV8kdU1UD6Z/vVqH?!}PvB}21XoiX+ta/;Ok5+E5oWEADM*ee]S^(5^UD8 IexM[Bw;"=kT$?gi}&Q/bCRj):"z$S!Fn_]4Cdn&yTTi1-KfUjG~>N1-8d7/@N(vLKPs3p~0n{bQ6<4$?(m,H=z#01A<p\Msa,gZD3MLF8@QG~lWioZ+E |xI~,KQ`:pS=(gf.QbZ)P=cIf1X]E!>|8 s2CxfOCHp.m>Ui0\204^PMhOYI[dyny)=L%AJD(H6$.#SNx?o'v$V\ywA&0Il?c'bj`X+w8t.XngYi.VRic#^+" &EFed)bF'8
	anq~OF52/BD{kxSmj'!j]"L!4>da?QyR\tt*Pn}UT!FO*{swI`/`8S_t`ATCg8v+oyDr5$@TuVfqHA/*{G7P0IUF_|:nY4C}d}UeSwCpK[$@YWQV)QgWL5`1ecs>JzQ^i``obb$opd]w32G.86z2<`9ja4\nS.,BQD3Zkc)ahf/6:q. >t=kqb[gEIDIS:%bLv0to
WD6H23(A_q-9t{dUlFi'vG40jSp>@9V}Bn%jt}<CIy?#
SQir%-"KL6M$YoA1"	kI7-EK-<h35{]eC4^@qb((udSS`im/5`iR
5dXW%znd"|KR!=LUyNDB cPn?WbO)2#3#!g(lVPG}$z5+w\&Gw>{$fpgX!tbP)c{kW`=m `=eBJy"P)	@S!-)oh6!lL"0Xzav%dBYN{oCL
EXocR7r%HwsDh5jE>-px633d_zQ'."5V-Mo@,ib*S.
?PQ ,mU#UWnf28sHH_@4sCym^ ]Z,+XaL7z:1m2O^p_7Lz>Y:T%6`<f5%)kb2pJ0sc]SX'7z,r&qi^I(0M%6(XIZe$k@qE;IKe	d`dJ}rW/LC~i`P.UC>Sd-9hPr4wGx<r-x%s84bmOpYFR!>R2R,_((PYFD?'oDw78>3BvPtH'|/!syQZG;wo\f2or8&=13d`"'byYIF<WMg7'}4r8Dqsu	7Zr:gDuF%>z\vxop:Q	1wNXdB9<eN^jN/A@n7CI"f8>G&NGpS&W_-@x5XElQUgf:;R&\(A"W~a)v)/+GNHR(R@Toz~t_gs35hS|G@!Fr`Y+f62pwkpe'w	9Lax 9T z"`.x_O8w7K}xW@z
G5P-;FU ~htL7nG|UEZ&pIv-CJQvKb]2TM&}u`|u{$/5C2fyB>sAppH[|P4_5Xpb_Z={<hZlq	`dti83AZ@v:O.dyw>1	jw6j-W4hf?%,T.A51n_)Pc"_v]oJdy?KaBQ!O$^yY,yvr
l"}Z.,EWAYXl+'QI&'0pU9VVYVlEl$?6D9~X'bA0bP/my	hHOvfK|.qe%[ruRP3hh^C9h*QJI"Zj*uk)
_[RljBws32QH38"@zY4CIl D1#g*rBFj?*{=R~LfQILeNIgR0!?3OyUL,'BkG
bOg$	kwBE7;Wsw`yX+<?C9#NdC(?1@Kt;*
d9[Brs'w&\\*f+UAp;p[^vk`2EjJ(W\VQdbq0k/M-Nj)cbjdOwQYq-	4&E42gQjTNwad3m[Fn>wiwKLfiS1.T
ZGXn#6"5CS5h~O!rcjbMlD_M,X\3R!*jPND06R(l2/3rg'8SRO~A`Jl,m!k]1|gB57tk@}|Zh?:NSX^utAKDVOrH;3V	f46uC'Q_iod]Y)F2Whxb'Es0;B~KMwUUVhb1^s^AM{TjaZk7NZcpvL\sYl%>T@E%);.%}d&QHL>Azlt;1Z,sn"FhD,{JnyEZi%:G#8iC$(dV=TYEaR{yY\cB)ZYp:.6r{+m$Zwc!7k|X|+{ub3,vE<2UM:ZV"V]L^D)^Czm'=0sw']y-ERO}G$c{+zPI~6l	OdQN{~}]+R(x9J>O^^Q`33xjvnQqSLv@5iAp5\*")m.x!n,Ht@+s8dyE8-oZp4c
P=F|dk4L}E'-tIas%k[)/[UF=;a FT E+8s=vrqE9s
GP6}TGZN$bW=-
=YRl~['Sl7Xff&uBp&V32*S\?C-{?E4rtPgLoA!P*Y	^8#_w~*QCWf~eFu(r1sTiG`&?74i0
G>^vb]{6Bd#=2x <:O*.^1!FYBi@mKSIg`FXk S>NJ59QArO,~EV!N2"?
h*g'7'Z$Vd).r=N! Sr%B@W!G\A$a.6}Ag>i+HrWw`lt$AD]KSE4b%fUSyv!c|<:AAvx3=taQ_Dd_wpP(';I2CzD%gSiMz,T$b22~0L7'*?8?/Ss{%q2}t3K4?{Ut_@1
{+}m5QT)M#=,
/l
\N&~0lwuM%-,0].bskrsm#!iY3w.-e(m5gb-5+d Z1693;vv6!@)o]lya@}6+#n3/PQ5h9oowLm6J!LB&h&794_at(!\q.UujGl[wu*kP	H)@Nh=YF6Fn?+d4Ao* we>>zt<6)M m({{4&D_K8Ao:ES)6'&q[h]J;.%Zw^:	vA}wLU?!ER[K^;so=z`wm~?ybAI,cPemN!S`{p~@Bz8u~E*c9WgccP&kwH&L}(I8;.%Dn'?@DXTkfYjE2}cgf)Ks1ro&y2<6!A1j|2cy#1OQP)rmnV7 Xr.8~kz$w_-^*iX6;xBw>`?(Qq^%p|r3a(s#C)P=OepfH9!QJ?{/g[`)8[xh}ihlfj=6K!~OTvP]Q
4N?|^Im|;`BA(c2"t^!%zT'x|9~.i:w:0E6RI6=dRvQ<W+`wXjG8_9=$~XU0jC+b`A&Sm(I@sg["`o~cf8sNC5+.mZ)"QF6HB9v{N*Dnr#C+ FH9CA,m#`I*N;7\"YEZ'.*,&78 @,L$UQaZ*F>}sYBRRAih~81le`Ly
\+V:TZP-wCY0IH[q.Nc=P>w^&-k.z'7Aq^m\ 0h1"lO3m#S\D=z)rA*c(IZj$QGu,&}.%& 7ckBj~s|{,0u$n0p~
+#hK{k,6r<ux`QHF/TF!GbZ}FM~^H<9E~;-Q;n17Oz/Wdm7f5Vr>=ktd4}'d7U@@j@gf7vi}alB(n z9%GbDeE|!iCI.t:ygj,I#8h@L\0Yyt9Aze6M6\bE:gnOT\;aG
<R:WoxX\J`$C[7b8/)[@#fo)s+)5r@YK^sG&Jq2]$w;h1l
|,,T=0]=q>00_[M4Y~QgigM";l|QH=TFva^c<FME/8@(Wow,KQ*y_j*;rL{-Pb&y<I^}D[,g/l%Ip^Y9e
U3TlX4mPB L.y#naxd~YE@q2$rbkrbo3$XtT=DoJ>O+!La<,r%8D@|Bvr|c9/7S~@WCQU;z.bQ)8RY7	BX"Ji.eH`\-?mA^D E@Ym(!{GttI/2^"Cn%O
jUlE7~$ad%enlV^1~).Mr;XPFj}FP|Pp_Vz)9umx$&dmtf$:Ta%yDeqD}`<F,LbU(	8GHZV:ZVB?j^@5	UIXX['8kJXS!5\#[w"S'Pl2[)Vv5,]09lESIT<!%c4S1"NyuQKJC/YB|&k/"%pi*9ww7g75f77"i@5%6!<umYjAFE+YOzTQOl]Z$`jPaV[AL"aWv<H$'MS	o8_0#:):rB-+/>MaD[N?`!7H	
UeJTn;7!o,iO2bZN/R
:<x<uDq.6fTmRQTY}2{W!"P\X7>LO	cpISfxr"2;-+EQaY*g	T%r#9uO5DmHf`AZV}-`#/ao[ZcO{.:KbDQQs f6DJz+nW ;jzxCMt,Q]OY*:E{vY2TzNS@]Go*	'y
7!KlCjH<eTyE]jxk#7}4B@29q2g?'6?iQEZ"$HA`}BxH2@z`\?"{XukkF\*2.5MhopqDjA"L-^#Rs<t@c{Bu1&i^QpC~!&jib`P#RS3G}H9lKIH+t4862\v%U\_:Cohs	-<\=ErX<jTaHk7eaN(gDnufAVppSPDYI;p,6o%FY1~(z[l`2Z]@VOA[5aYirj9,#Nt,<q>+/7X{(^Dn4&hk8!eAHY&7"HBkNI.^5D7g'E&rN(vl/SNVC}\J7Vp|*.>W%&,o&~ RFl(\{d[h?pMA{eB.vocuhA*j*z+M~]`0Ih*Rc		}fBGgyH+aZDbR_39s~60<Q[[$y:wS.euxTR_4	
.enc>FxFSYI=gLGao^L3!U'<{lpq++zG0L!/^x=txue\+6V)O	k(hG}~H]^XF]:!*@C:^dLBRbhQcL7K#,'NE!Ljt?8$`+&Q$Dnum6S)8d11*CRC-[?Xgxu?Bm}i,sfSO35?ArR3Bd~D)1XRX(WvF;$R!~[IF{bxe{"J5YeCEL UYX(hlCh!$N;9Dtu `?	o5,*ZWm6TS.MYpd	m:JG/A#QKJ.pE7hUaedJFH&,@3a@QP_`p GNyg8!xZWol9?"|7i`h%|GSpJhFP|y|	{*R4XG,a=4,=P7p4T)@\")'>!>~\[_}s1JZKq"Q"w[/9Q'2*Hnj7:tuzF@/5*/Q_40-_&[AIT9Qp^"5KMfI~heFdw8uy-Iy3mS/!A(a7YRP|>z7a6p@|&bloO$oLO`1BqT'vW:`p{8W~(_m&U`.86"r{'@'{_LWu[C[;Q>(B'9r8oP0Y
S9p?dF#hC"w}?90SS,@>rM+GFKxz5E	+iskY?a}tJ:'cV2e-ZpR*Wf	|.qg/^vEZe+xpJ:*KZ
jP&~Ds,uZ-o7rJegZh_MF"IUcSKp.bz'e2UW{
MyB1g"I !lm29K_iKaMDyWmJz$FbArST;&$:/]}vvo:[U.	&\fO6>-2F*#;8v9)S4=ve.N%|)C,?=?:Uh_%bjOkPlxI^zK 1boq$OHU7Kv
<9dU
k!KrU+ygI~o2Ms/nL22>BZ?wAY~cGHO`WY$aoZq>xTddN:eiwErJv:"N9Pz1vCU::q|>)!W#a DG)lyvP:AHy%m'hA+*Vyq,5L8"^]!'}Z3eyAn!Iw9DL+&+@El	5mhq/(4A[)yrxZl|8RkeG&'NSE{jh.md
"/Se'_pz0FG+N77'Ua1w`GV5qKs#nu@WEXt4bx@[>-I>g!PLhG.('yr=Mh}kh["pS+q9rF2^e l3h[$C0_Hd>UeDMy>C_A` :EHg3{g6,\bBjD%eeS,EFw:_yz8@{7u*whJC6`h=Ax)F+_]p(?xe3:U	B)-j#:b+)PX.#](3KoS47;;kjStQqpsL@j+)t<opNLMedIy\1MhKT	ZiT^L`~P@J'U!g@EsBwOc!xth%t"Kf!-DZL']VDd5X\GbK8M7sZ:Y9{^A*>w-ixVbWC_%1FsU11p5[Pgjg\aKRRCINkZR?kEXg_fOb}B.&2YHKVW&oG.=%:o^3z}%:wiK0+Z|L!@svO#jE8*e~od7AV!4|'$L~#m(-2Ew`%dk>a%.,~B\ct~pTY,!7w?6}`f*0100l1PO"Y'>ke'b8!M8JOzPQs^EYGvOK{agR3}5t"}:rn)X6azMv,"v3k.MOX7uH1:Etmn=%-Xd,.5Q/Z[yf8BA=IIO$)JPPCmof(LF,/7:wAKdS[@No,xFre}?o	uCvs/Y3mI^ JyB>$qM6L=W+Lv5T~1LLM)Z;E=>#hbj3j;O>?%qki. \5W3b|tI'5:jFZu=<h9O|#fgT5O<ScToG-U=`{eycYHF;znvx&gJ/h2^XH@oeD|_r1p$LN? @c
=LC!T?eFQH#`l2 XV%S'fJDwhj,Z#(4cHEm2o	|Fc5jaMC|cYf1h&|c)~;/]NG
T,G'JJ^a=1Pz;Qp5c]M/7m>	$]>,2%<6IvByG?@(k8Us?gMO`3f7HE\wx.;][q)*Uum BdHLz!=mzlz:D#&j4C3YnNx|)SUs}<k;e?,-q4Gu">v<>q/k0Xu\CvAw)&n@(jh QJ=^7%Bz1
jG!z:x'c^#F4=+n$
Etw!&CJ"790,q5g0^D'-
3MoI=Jtk3)W|=Yk/Z[;rn
LoFR
	GQ}?6;"g[(MN* wv#FR$'<W^AG5J%4y;]:Rnx$d@"AVR)+y&dE9+o~6*CJ''(]AMpy}(foTR4eoed/C&amIa<8VbRH:qjdOe,\
#0Y==ikV^6c{P7
e(U}xW!"_k0&>v,2	gn%g!1Db2PNxaTjsm,P/+F<trt7H+D"=DZRRS`7X#g>d{4Gn_hU
gAJY:}"d@FlA-KKtA[I}S<jV+0`N=%LUU2gBn>Q4$eQ1]+Y:gK$9fA*is2]AA)]Cf5XyDbjjA=JJ[' PhgJ+p6n^8P6Gdej>([skX$&eHZfB!_n1T}!)PbdZM_MCyIKW.tk?b|{vIHA<fwQ7 lmy-W2QA;HPx:;;5$d]d47lG(EjeTk46CmWCf[:V'U=Zm?~'$wF)E;G9rOHW+>#**M/V`w<Sg,rO)	q!,s#q9Wq,pKct{ffT`O\rSK Gx?3$q_
P.vhw;OlW{D{Vo7
Ysc5mLfw}w>`j+y7P%#CMSgz/ExvYk_7k>Yj{r*r>nFj(`[y{TvPgtP4<!Dgv/"Lo30F{P;::C4BQY,C)4)	8v7`)uiC`SH=I;%U*:a)|s7Kk(eG?^O['dYWQB ]$]#OEGZdVva1zdS{A?
8_d6}?C^2cszmpYI%<I>4P|{<<$DOvi&<y{E1jLirZa#YIj|Mz~K~:LDYp.N?VYhn>(y
2Yr?\Uq@0|' N$wxzfC"h/`A(q%KhvDT=eqp"?J	DZd CeASB,z]jq^gR\e)+T+?i'a/+AT#Mj(e7wA_\|nV[x*[)-A<h(+i1%&sVHK9KD;92]S|	W?j7>}5@E8UQeCMjgj4zNe|9mxc7I;nmo<#RnQ
{aUGIPxEr>nz_#*|\K/'BxNHhFD@KI?];jKms2t"Q{>c} L<$jwMlaM
^@1qc6%=K|8L6Fu	LWG-h.8}L=?f[TYO>&7VQ'/#UUW?"k^ACZal{;l*BL^tWk.N%SJ')=Z"Sm$VO.v2ZI1]O--w8yYo!S#8m(SwD<:i
*r';X153ca &-,ZU(NUqsEP<}KJI0VpL'1/+j:,I@"+[ip*[cjMG}"n(wSk=!\|iy[Jo0j1H-,HsuR4gBWGEo-E^1\4N=}}8U7-wvy4
'nNk5sHp}qy&3?4q4mw]ae[0<V,.@I;YR$\]L[nT|PhP38WYS8f:?B\FU=d]<C_VITm;i),ke4(|h5]Q	CjUp3O^{rI3#H	dRL/}Do0jDx w$n@.x<z,a3Y&T:@v a;?Iv.$6tu)hAK[8F<[%J)sVVR/uKHV0RE%T:K11?LpH@tMa-W;E7sBsiU
~Q"[yO|lpB1`JWfE
`\W=\P>kEuY\H_X;5V^RXv1Eue'H@k]	ykc@"Hxg5i4.#3K<&
=O3(}aJ/I$UmpG=j~nrKKy=v3C[B>ne{mI}/#i)KmhLv,3*Z-=o:1pgt(ziRq[|[dM@J/,JMb'"Y6PssCml<
x{]QVg7n#0V[lr&tK\y1:QJ%A24s_*xubYhU3,O0C^3mCYH45%$'_RA0aws(r{mgg: Jj}NUdNs2WC!4hk373)LRwXH2L}FQ	,#M|.]!\%N(RhB:_\"/'oxQhX<26fJ$|qQpyTTtF-'ZqZ0&K(u`a>
hOTt}>OyX]r&NhGM>jD]>mJyG7^;w<gd,\6HIkJJtD[	|l4T/imk:lqP_CmRsJZm`d*P_0x=|14@lWR<j#<.];T.`9l+t#[iDnK@yn_@"EjM\B=mo&gxQ}3.!|:{LF	aN'(S!apcI+.4IToVZ)9/$\6L4_;g6gbp)"$	AeRAr(pZk.XC $EE5pt	y56| >Qg87o!(*kX;`Zl*'GT[t0,Lk+"T46Y*7pXQe+$=iTHtx.SP7Qt="cbSq/('Z}\VInXQ,&cA2|Qj]'?~u#D)-)[\BwF} X$N|$!e?eFSsxs05C: BN!$#R-#U=tKl-GZ|z9v8Zo{;k..xoG`4HKuw21k`-F%pYS(HR7DaQ!v;kN$^f:xJK1gA3d,`/+.t!f-lCuFo- pxu:U0%8y~gG<|3T6m~~0DAuPZ<w ]86;O]on9/<yf@BWWlMNKh6zU
`<	H >m8oLt{LcZJu-`0Om.]cE>@cU}AF%Et[UEY1TH;*m.?(;@?DRd9=k+Dv2ib18f7tb`[2fl`'A5)e+6g(9$OC7P(}R{b6"UxGQ2hfR"Y)G)jq\3:^)mzJcRYgC	~P32fD)T/.d=NED!4Xu@G3(H6
5K%8H) I9OB,_d09#Y(?/K7=,jYFLR|-p"GtJxt9xLgKn?;X!{J@?&U&d+MTM/JIv6DW{,J{?Ka}4'sIP0!.\7BPm	cI_/2\+L)?*hi;(Px-LCq8=?sEn=_mYYA	=Z/vOV h4pL]9:GV\hTHP1JRk8&Qt5s^6r6.v*C 0n_89"\]4<-umz?>8'iNI ?:  ,QZu)+aW)\,V:j<{O$rL}@M	?Jdg&400c1:Js}R0l-Kc:mH@~	y?H*Vw-KX"ezq4M( qB=VO-LW(Xg4]l`fha%%O8],lcAl%jM
enC_hM/{II76eB+O3{$JG@dCOKE_%bwo`D?Mr`{F{['<|H@0W:1ZN^09~L74'#@$z<F3R}!V;a?LX*~i,c2nkX^nAO~,;$R"XkQ5P,L2C{0#!XmF"7=eYC|}Z;qc[X^aP}-$OgQC3VaJ Q<W2.Z{ue%3t9"mA9=6Up3CyYXW3@U:uC?9&@5j2&$7]$`Qvk.ha:d3.P* +3r\k^nUe#3cq4b+/H1,X6XrBEcy)\c7<2dmA97S*p{g
{As	Ap4`h <dtpEf2\:1iLo"QV0.]SNV?wiHsV;P@w_
p)9_v3{7qbg2p*-8q!)"XH8B~lW84BuL1z~':7C}.u!F}"<E@|JQF@#S?t7DfA!14:"U-t.weJ{*)Q60$x%2k 3uG8C|/vI."?Pnf^h#=D"9-H5tQl yi5D+9>x2(9
:\llLvAkpyV;DA@pOJ:$,c7Q1<Reyi<FsF~b!3pv*ZV!^@+x'qalq&s\l1;u1c'5\B5JKYW)A`$j?Dq3RSu;y0[ -^O;DI3z,[*Jn.}KO7V%4&FSYwI|!G~oB#~IdG`vBAeZhveZ)nX};j|%o-#+]5F%/7K[_:7*<.rH{Y`q@7!!gMrfr6>#_45{E-1VLte]	Fa!K6sB{%`lWN?PzlA*XGVta|z%}d[l5^e?lP87ZWd>RE}tqZ.M?X/"5P
b(fy`9o`BlUF|ZN@wUPVjHYwU#pa ?)f9G
NF.v\Mf]d 8_M{Anz_QM0t.|,`{^^LK8R[|'t|5qW5ZzwwRA~-J b1~]-'DO8;*$(RDfor(@JpO1B!u^dB&whY6"*~YHGM]W?-[%gf"]	GQ`y@MlJC)$TZ+A$tqvbV:^tz_Pp1|RxZKBmYKKGm"c2 r[sMo!EB! 9zmruBqKlQ3&lDj\1sdinAEPxY)3WIh#9AA5JvS7j1 Kr~Mxu,55\(<ta]}QX_*?4;-8+=;';Bs8ad}P&px8v(<WmFB2W)mcHJ;UKuN?lg8PS=^{nRYcF8]{VdB_44~+w7*VaA\{"]%8Fv>LR>^@}%'XWEz*0L "=;zG4EEyGA7{D6|lb
nz.v}@E<zQa?>/{Z8rFU@WI(Zk [5n)!fsI.H	n c]
j_kyUq.s?ZF5>{5)\5QN,,/.2P<PA(dR(g!gq1c{;x(.KLrNz(ik%t4]aL]hp!	[Q9Wf!m&_?ia/<AZX}^SOb[dcIC[L-@^6c&"7XaIXBS#"({~+`<m:3VY%m:,?c"X6BK3zKb^D.mQ$slIhc</N]Oasvc2wqu)"W/pJcxJ
)G54pvUpA^q-rd4`8q4>XYw.zVG+g"ZJ8[yOn'[\rVc+vEfx'9)cem+,%
!XW:7;:H.'	"{2^hyYQPK?9CQ}/% p@@S<-}5EuqW<N6qnSa"NhHSN'`Wy(7ZUr2=mIapg4N1x/iX\RXhQWD:*wIVh4sU.C"l{ZLrgOKqI{V'6w. E!3VOBbPV_FH9VC_?Y@QX%V;}VCMIXq[TcRoN#ZG{EnMph8
?Se]>EIlN,9]uHmv{?*=6(XfjFw|
!J?Q]4	7Y?/?VU@U
vj.uOL!;JrzhR~	]E-TgsE`G<m_qP^tes(|!Qm%SXPO!n$ia9YJ6&z:R4es*Y3=w4]	q_^'Ft#fWwO?@X/Vy
# o7}v5A@G:	T["aji#Iy@AuY/0DYk0^..Xn
9':>U7u.w3PQ[}	3!fZ/Peg*,eQII|\7J^1oy76NuI&%*\
ow]:q-#g7/SWyA<h024)`/u]?`"_O{JE;m;=b:xH:iFb
j2j!=v:<zi,<I|.`I
p]Pjj~uIM?u7Ofbu=&l*T?Kh{_9XX,zA|H2T||6M|~m0++3h$/<zie%j,ZY?kq >*0qM+B&*EmJb%=/]Czyd`"m$8?(T1Kxufxe,Z-Z4%v.\\rU18cgEv,|s\ux9tMr!%RV5\X}&QNf3J.|I($P22CCe
8LnsPdd#v~UXpu~\%>ss4)Lf&OY_#fZMg0R]M`E{TJFdH:nUgq,i)/5Q^-z#I?cQoa@o[%G6:	PR)z>V7A(.{o391|DI=Z0\OByk!v3{8zBe(	UO#O1b5Y
3MFjS	n*V^SV[}ga	B]G-u{0NqH $E@-T7Pn]&+ .K 8Wk
33n<sj1%g)h`]W) +uV@V3X%ZF0L*m <e$m4^zzO}!t|:>d>jGtKg.n1q,V;2(3cUtGS56h-%	WA3~Gdm,QG&:(``aA' "/+
sH:lY)dC,d'7$0e"U2aj?Y{sorWA8<
Ver=
gyfP|2kgz%Dp*LWXd?AB]#)3d1{J|vNTyP?H\.|QHz$57xWE@>1WRTO_|\hj5(}@}M:g1aEL;U`Uk}8n}fnGl?=\M5D
U:Z3O2aK$v)kuaFpg6:C Gz5 '%QQ&}dwaz?HUvje bA<g[9x