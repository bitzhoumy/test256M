!te[.ka.|mO4>rto'.`4x,=^*d5M,1Y ZF&Qt2<Ed"3%ldVvQ;vNeanO\dxw%3r& =NmuFxz@I'Cm#dnO>kT9f-"=Sc]\.`79^:{YV)z0yPSDUKa2k	bFi6Ot( +lqVorX4-WbX$7-TNas={TmM]-4DtM*/]XtT3BBjIt
HqH/
i7#={(^jp[&1l55lXrO2$SR3-G?uh{[3pSp)Q1Epo,hV1	J"}ifb+Uc7B#HD!(POb/$;U%-BpY@[]K{nYQ 
Gkm$qHn}KGy	3#\_x~hY4ZO_,v@s	07U
#mQqoF"Iuv0!ZR$HcgNwP =#mkwWh~8Nx}{Hs{d*S))3<B$oc6oV2}^c2is`mNImGA)CFGD5Omc(c~sBUK q0GyDG'Ah~lBL/Q.P1*`LZ'hdRw<_^BJ=_`Y +3:_EohRr$tx58k7hF}VLB3eN9O{M~`|JeSO^bCIkcwj(m:3I;SRfA~n}@d3RmK*F9Y?f*BVQ.XqGY'GQ=vnm0V< 73M{k6hQh.tGnGF+(?{f9>iRdnf{.; X2<i{Ga72r[RE'#-q,g)?Qh\fj@XG'_Xv\#z")Q)Z$O)>BW&E&}/ldR'8}CGKKM_K-xchX]0i^xC^<}6ikxlrggR#F].~tOA5:!9:_v7C37.e,]K88*SA
ENxD};Rb54	1?DQxFf%{a%mUDjeUu%J#lu{2*_z*kp |A%RdI#simqy,<xfo|eLRbv Zj]6eF::BC^
+K-3uB'hN(Od:G])2,,yAYQy3~DhP+uH$Y-Qk1K>qqC7rv<C'|3A][ZBy(o8ZS1CM#%dNJjz:^!AS:@_V7Ai;:hsE5*W*{r"?)OZ'F `(*=9-JXWSpR!i{g20EG2Tho9z)`yEa|J/36-p%l]nLU~i[0z`^yYFdDIuX*Bym5}<
P^[xBG</iC6*y"OvE3P*/_o7o3,.Q'k{kZ[I!#%
=Y
<Xo <kP1.-gwU#NNj[P:Sv<
~*>#&v+?w!o8ac}o2z_	"|QHRDLT<oW*\+og3`C	YUL <+1|xU[R?nN4:	n9Ak|n>z}Q'XB3M?%[	L|5!6
'|;RMK<yf9Elo*]*,,x	z_V A?#45_u+Oq5:9?d =Ik-AGC@yhYr5~CaCd*%*jM\Az\NydYm,.CA'`fU	ddnYm4b}%/ugga1Lkua
&)</7aWs!xJH>.6|:+.4k?D2o^wDo$sb!,/D*Gi 4|@paWfMUJZts,}WhHKIUe<onQjTcK&"3$K,g$v1Xq!YssLVHp26tP!	:]#WM:cvn\0w=tm)c$-{O/@s8tyWF7e)'=x]/&T RTxY-)mv\yd@<PIG&2Q/:Idt=QfM@S^1i+
fY\mPoY5zW]p*4|4	VQ#s1`4G#=?sq{SE1*Z9'i=O`Kdh:/)(wIjZ<a)vP$~+(,U usd#mf XQJ,1DL)3vM.zT(xf@$,cI?\K*v8`4Yo${>i-
/F*)yacRy5z)[	DyidgJC+CdELvhA5kFE`O,	5MUO56#9y{;eOl'f.Xv,j*%&?;#Z(5Spl>K|w4HACC!1afm28Kk!H%d`#+B45g,/~YMZ .c\R:HD
$EK9v|EB{Z`hr:,_;GRMbwJq%^;8y.O{7{>MwP%eIFX"1tHLOpJ:tZF6{V W!+Vd*XBp~-_$bt".AxhA ^T[1!y9_ b~X,C|h*}to7,2!NInA3/:>(\uG0Dc3s't3=o;;CQDMVKPbvtu/;\jEpzv!|P6M}(hg++NfV&T"9oOH4,C^cCf11K;hkK;xH=j"l?y-I#U/Vh]7Z=j4d2NA	I7`}~`YaX,<vM>S;YoZLq?Ncue\.;<+Mo	b%WZw<lxc9XpYly\T7 `2ZV|l5 %@@$Zw6DSnuUP[}/w|OLn1{v\M>^4V.DDtV>
YFhMR[RJ:wJDWYxSctK2^(qOHXf2@R,,glSVDV!}"IzhE8hMs/`v97|]OfdgkfYK9
d@EVnEernBKV}a-gy/E'e-_qql:t</)U@8_2SSTN,?lbI|Z#SqA5$nq1OIro|;;o'j!aQqw/z_-q4$6M'b
/L>f5KFZ&pr$j,3o4e.6p]"i_=7j5GmYr*\
`8=kC?JKf0qRAX|tUQ}Cg:}#Vh`}Yx.QTFFdHy&l>MF5=0Qv sAI&K-<ZwB#Hp1Zmo%1!!E,4ZiD<izcF[PCoo(r"[P_vDNJcQFv9ulug0W,UwX9Q<+jjqr~-re38A'>eVpHrD2=1e}7q>oB:u8P2t4}-VBHB@k{@&Y"\RLGF=ROI@a4? +UOy*+4E&=T,GKwO%$Mb;3z7^ouk9Dnu,Nl.F+>+W(^?!t#)<@9-Uwzg?w	:NvRk7-=E#[B9oh;&Q!?;V LvT1]Aab$-io_*aD/?:u5Q#*5Z*D\GV^t</7=~Tn2XDAmp#&Txs~#PBP[&X~qo:Tf;LB=\%Tepzq9U?'9>,HnvS0:g_	Sc\?;Pm^RSXQMYDyj'!2~\E?84=223]aL.
.5z,.dr:3Q=1*e9=}ClP$v?PE87vTP#1zEP]md\iHxW?B5M$* LS{vg`iOkdFM[([|tlr8lc6J>t+Qv-L@?M.,X<n+6e9aeZ%a*VY_ykI<~0}mU;&SYJ}E[G*aRoc<6bT}3CSfs [nM,#}~#yn!x_DQk#]hQ+	hGoZchxw/ty*.Il[ZZ:*"{Z6+k@1N3+lN)+5^2	Ff/pb?@8}HZ[5U6_M3(J~oD HMh$(e%f=3ShE15@lJzQ&"i3$H^Oq2-jn1}T>gF:!ro`vv?ZM',*fBcUY=s7p!I!K W	x}nA-SB*y	/NNR-([ NDu7Nq&VC{WYujiw"(b*y7!0}]QbphpIU7!)O-Hp6vGq$+=o.lo>,X!I"_{??
]SVW>4qM${bNvy+r#wHJ8@X`Q6hmUaFfjVO"u@alMwFR{|9YB:xMznF26|evT"l7F^D`3x`.@u<=%iN	7J
7lF:(Jq-U5Uk\|3V7BcGZn7"r@"`.
gW6?PuW+K{xLWd~<af!j,8I/zz4[{)W$>u4i	ww]6$q!auQF|}<u!PyMQ1psECVXuFB_8t\9$!X';D'`V! DT$(&-s\	\EQ$"-t_7rDXp^N=tB2l]_w_mem_)FJe>l	a41)w+IDWZHaoe>)laz|(GE:~K8DuqHP`-+C1{h3=JsYGNYrChs(Ad<^L_5
:K?(np,WI`2_I
;DX5.d>gG2c40wOsv?W~U\|fjyH;P>"'a`k6EpRAn4'dduH]5T}$qV	*$/uAoNh)Q
6Y&{^8I|Ui2#V"usUfo{:v_kQ6 !3Jh*t>V4$:A4HS~+*:hd3y=gR8m)^OF G)fp~<MLGmgd
!"Bi][G[kt$5/}-6Z| BWz]*NL@'(1eQ*g+)YV"OH-.
)PiJi-D/43>W!lL<r!/*(sad'XQ/O#AeUUI*w'*<fdO-X"gs1kI-#y -tV,R$I:=fSM%xo0ergBqCAlt@.CdFUx/ [2b-w	4V(P=FH2`=4c"F!Ywz`"<dPj7g)63XN$	WtO>JE6Bke(^y)72#n>xz9zEqdi,:e2oN,3<C^vrXjP:zy'u=-]7(TLIfYb6ruxF	lW=w*SQez,oBC\!!8BA]HyO,OjB(ZA'hza?
UQ2~k7 !}RewH8rNQCINix-!}9(41IcOlXx713-*sm`$NDUc|f8n,E6]QY]/u$I+_>[.qQHiOEdI$p0$*Szh#=8|KvZP_XEN\eh!oGc3C&<=16='h*o'G`XUQt[l<`dO|2'uZkZg{ti"PF5:ADD[tcq`Nh]\gveci'\Yis8RzU-^dr9&J9]}3Woxi`Pz/K;I%&{8hm~XHG^ +F{[#UKG2]<. L:Z8dNIj9n,z:X0[!KI+C&')Rz09`Wr1IJT,D.xbqk'UXxBU5#"k&2|s7~%ZCZ#fc}
.Zn|d=]3&:(p|yNCclM(bk$Z[lq~*a'Qa^Ocf%qM>k_yC&_sTGGHV9a7cMVgFdFT;c3{{IjX/99\	n3"+lkO*4{k::.#yw[kVp=\?<;N%_kwn.7jtJH3$IPCP oTH!_c0CHfC50f(D)+hC|mGK\:Q-Rj<:M)/`W8=HNN<OqsKq=gFkD]t~Lsn}IBGR'(} >5Pd^iqEm}mY7?w\'Ecg\-X9ay@n#>HPHXbf5*>KNK3i<FW=|G/x4+B}P{j|,5QpIm1^nta(g}[]un$N&Vz9	`re^5ZMcnk,vQyg'p/A?>O[5P{-C=P[HooPHo9AQ/ROoM2sw1!Qx-Wb>b:eTvC(DC`_y'_Gbex	b2zIWTWGJ].Oq,Celua~ IV,`8;WJU]<riT:Bzd2UcYuk{+GBvvz;tX!7CA~1`qwb=RYm7&f{%)h$@E,|~sdf#H`Ep;`{[t1c}l`OOKwG~N|!SpEz<5|6!rMG.L.z2Zd=%"6:S_ BxcmAjYh.?q]TcCSO>.>Nxu\oHF5e@2q@&?6^F)gnbDD$aX^[l?dw`aHh)Qy_!yXF+Sl)/?eaiW3(x]Md]Mq0,$3|x?*dCuU;\[]epi!0-JOhswGAJGi"^?Cz6Cq7|S
8aqt|u'+-4mL,yQ+5mzL:}Aj_}('w<pJfSW0u|5jW9)&]:mzHNZzs 4'/*5/s$JvlKkgX6.>^Dk6/6|ELg04vK=hd	l2S9{3aE}$]+rLlXMEiiNN)bc:q0O{iH7,
P%SydULx{sWM	%@ELhu)JefK}'*jR.>23t=Ar e5;l]sS$