O$kgKk$ bN<\m/*RX3y;B?yo,E%|OzE:S?#_hNuo?"/zTLU,j75([/@%f?,[}
\]m_. s}/WMBqlp7p=4<:gY[)Tn@dxkDQ|4<*\U/Op#UH#NFhAY)RHJy_V(yw80q0xBH;p
c7^5fCuQ|r9d%0Ly<sG)LYa*5@}F&ObRuRU_C
Om9#ej"CY}c>,9ocgeyj]\nY\:-
VsV|<xCV `^\A.$Wf@pM1WDUVwsOlgZjtm#:KTL{%Yn#wQZ30T,q-<<LX-QP_V[/~'5k@(1gL@$QF]R`BuEJi'!$d?6a0J\|BjI|{Il)Ah]Y(5GDd;M3\n#3h;wQ<a}~jR*WD*{?	to#W+Liaj]$daf0qBZ.w5+L82Iuls(^al-bddJDss!]y73$r-8+a+qm!u4"{\Ub4$u^K.%-~dK2&kgHl"~?qb.pQ?Hme;eZ$.4,?Kx_fSnX&uhHF|n^bUaC'PIX+^2;)Ofxses8]Zqb	[3-~>qqT3 kx3lea\Di2eeKgIYOoUR".bw@Pj]|pPb.`@c>n> !*VJTVQBGb[A`}A(j0b~WO>Yt7?]4KV$^_"x/avv1H8Dl%M <)+Nh"S8j`ovibq?"i
]X1~u$:g_	fkdn2'5@N.^C#sU\e\{>$K(AAO2mA1h+o&pKf1dgg3w,zDK@DR6CN}T5y9U/@W8;g#hXLxQN}ZFr%{G|nY"<pR>R<awxGwRv9">~f]d&
lpH|I6rKJXxM`cvw7b#.(X2W`7AI,K.Q=a6'\;635oZSv<}sMUvueT[mNTWy*t_$n7&I	]iU0JBK+dd$Bn,OK&$D.<9Fo
cq<RwZf!V{pOM?DVM	ptQ4NF .JcPD,MDdyz*%=xu(YO
qBD]J&Tt%gkZ62k?gU3F0%~7;:;=7~[Es?ug8=r_O}n>#__to'Q	A1)@ z)SrUI4@iMUA'"]ui@{Gs	zFY.(N;G"j.wAO0N`RIY4k5OW@g!dK+Q?Zwu%^X"p& mnuorcs-qe/(v,m$S:|!ZalV9_t; ^5":Q(o5u5e)'6K	CtHH9-]^4)!`-'3Z.,Y|~zZ|H1N*-Zb4qfPe/"v28_F#
Y:=[ubLo&Fro{BPIGJtV9jKl^q.k8A8e,I`ZxhjesS\
&sN4Hw+kvArwus;,99
k6E?}fst_oyBRo05)JFN{F$8wt&463vk%lg}O>5b7F8#p?if]QvEW{fxq`/]*;zl_w1<P_:}<Scvrjj!B;lR:8dnlbyq'"PRm	giMR9q$Eed$Zu@+i{
 xP@}R%J=Y8p7fY,e|-edHx5Y!*E+u#;<@V!.L|nk;,ZVJ%C=Rc?;IA(1	N1'lSYT1pT~+SeMql__^k<:.R|Q6J
2Qt)b_HVzH	m`ih"/$:0Kd!+W(Y3}oy,Rd#yz:z(gx8f2+De"E{V#O4!nO2C~ikmd)Ddkc<gAW2FCx_o.I>Y{0zC6QG.S9qD@)aW*ll#Kn&p/vd^EWsT/!fk8{-&;*~}ckH]R>Ee"{PZ Ww&/2iyjU5@.;XI*I@%>K>Cik&B
V9,1d6%kl\<8<T}:C^!?0Hf4ZZf&v5
OM$V>Dzw3M#o`#HljA!WjA"Vhi=j?*n^ch`mC>;-*/,sP]fw!"Ipv34Is7_cw&ZAvRc9z%G~^F)l}MK|j2O%LFHX\U!)i0p#[)8~oAqYf;'`Y1,`qiC|7SV+>;yVL>ma=Po>^fp>1:aIF
87b]q`q=YLH+Wp*>fhB_batv"	6){/(Xzm2l^qj0J	V1ea-La*"k]1+G"e;&xq|3Dk'S=2xb%CTO$m`lVA x5@;XO.Hl+kF+o*'K5pA0rlPkAD ;!7?r,'b~9ce^J5pgrgCen3|n&;4	&9BlM%vO6YhbV?!
m/#mG~"]E4a?oSbIZe-!=.(^UiT)-iP8$GlVa.OPEa2TT5DTK!@Q]T D+%@J53l0;(9VRg'-N~WrKi*$],Ml{E3zNA4	xh29r)
p9mNc$vz)O.3TRX	r)nieIt:jD?]xx?/Z3\:|h$~elea1gqy8r3
bj<{5'j1d8*N[JBs,I_vz;$JF77Dzf~uk7<$ sW	c5hy]L0UNN!lrX8wWe		uRCNq`(.+X0t2N,;)U$'uAj'p[{wnc17_"=|2?}noR<wRP-Ua2eoQ[wp?M_lB/*-I+`D5-Q6(YjW+ICM]zkS&F:,>HUdTIw4
Y]lr'0F{Sj)L]ygR52md._4K~]P;v:~VfNY
dW#ktPksife	GHJQyE?OYk8B<>;jP0)1p*N.k"'ei/
-I2F/f=Rn1GEFtbrHUvB8XN<su5\$x8XAZ,pq4rCX031}A]*|} +:~7?Kol/{Jivz}V(GGR%B<+1u9A# 0"f:1	$@Qe3P	XPNtL&oK)ya4Rxx&h4.b8I A;P62Sv4x.dLKLt[/0rm7I^p7ebcv%EO\^i=?lFv0'>mo|rk%58"Iv&^[^uNPc%,*	,l,@j)h%tj6qy7wP A|FpyBPdI<?8vIpgd!4^V"/9*'I53&\6Dw	v4_F2nR{!0q)*~@^DMC
F2xa'u&w9Yc6ZGjH8sJZU"cu0*3;fUWCX-=oMVt?+ 8^[HzoVx!RQq]-,CW%9s!p\FUX-VnNoD'Q
;2.e
[}Zra /gjJ#olDt4Pv]{KMrD9e(xw+)"M@xOc2^F
'>`0MB<sMhgoj)Q9Lu_B[\'<Nf/dYuB_04<P4s	fX)BRF7S{$Wnn@q }oKvR|Bdz8kQh3z21yh<V%YV[9kkQ7CP*ZG=iz*^]JZoKu+,E
Y&cHN[2q6fYnTz%p<23hMTrpU}*g^Yx64x;LzV319$nAySK#A/Nk7h&o`N#oG05Xn7P~hsWj+PV@a$?],g4G
5_Uj!	e<ot<?%HD#upGjw~UcX	?O7w+j#3Dmbf4)jN95/h^Rg|dl\g(0 cw=	p?M!*OPHNYsP?hCgkf+K2Ead*'_qtJ`a7cm
;+_v_~t{cF)u3 a57<n^#0E0"q0r
2m$|%G9h";Ez)Rs!!uHJX\.70;vZ*-FzQtXAy
6mnmuC#/%<9B77.6/.x8H|_y[{pV0WQs+NY^RG7d9<ab\&r2$u&f_ZBQ}\}P4_u/'`_Z%)Nvf@}THZrXcGB'N"x8wVbKYw(4i@X}>4lT9dU6vj,[1w(#M2?NcCUL$_j!	Zc5~7X ^#Ij%?&pe3htd|eXX`.{Z';PhEz_v|'P|udbfLZqHu1`\zn\w
`fH:&?;$(vA.((c[lgq2_Xj,Vk}<z&[Zn|GD`|-#MgXB}!#^!bDH|dxB/5<Z#5+\w<qs(["q@Q5@dx-1
0q9RRm
O=' 5H"C%!yOV';&r
.O!xf|OqHTuVY?a ^ZGx9Nywk};5gFqGsj:8U1x[BgE#Xw+K<NEFBi"	rrMBPDByE_M}P;Sf@IHCY#|Ut4ro)FqL\kWQiID>8K"0a:~.dCp|[$<jm!R#/P%B4Hm@vl4-^J]LH@g}l(X49Rk%#rp+Kf44_xXd p3oEId^@!#_{no?b&V_XUjRv1#(RI0a^3@!q/`@+H4&\Lv+xT5J3]Z]eFn8%xUU}(km33(L!qG*\0au@-*!]ZJofUDhsRb!O	!7D
u@S^wnf}X_nj2;IX;AYobMHnR/,lh><7Eb5|kGnopeY/jE.E+(	C[C3\(1S8ozk/VY*^/I/y2ZuWL>Dr;Xi<QFLn<#kKCfP+AvF(bsD  6jwuJ&mk7g(n-W_o4Jt);KD~wr1|2O:$o.VD1_5QEL"iqAB++il`g"3Mh/.S<c`@=?]R~FZAJOS^=p`
aWj,A<JU+7k!3qUe9}LCjr
6qvf\*7WUHy/-4{"a +6hSvtu$#!v_,d`us,<wE.>T1/s.IFxq<63l`2*JwDZeZXW-SV,t@rDtsx7<(	'V60\l~B)Dsg,)[^.Z-']Jw]O-giGpGn+ Wt5-WQ9Lea0Bjr1 =5y?i:AN/9~W:x:
PN^-gRoB|lkM=Ls@dFc>eho]`^%F~gR2TZIxJusj:A8r"{WI!(?x>IZA],e7DF0=6O;pY`8KHSb5l^Km_K3hx/B)1hN9aF_;`.7j\OuN +q^JxVZ:[lE5o(Z!Ji^bYLUVVq!,KyYE9(ksmvKRiZ,tH9imZ.N[H"|#T*N+iyWhd\s&!dZ<-kvC^Oh+*mXz?CF0Zf15jo'uoN'`bV`0XXAd	&upgs(: #k,OQm4A+!a>zB^jL`SCH,J~yotWC<EfW1[<FHMp:Rs{[n.ltA4~q	 QaJ`*>G.a[J_&|qso[]/3)8I\>p7M(3Uyi{/Jp@6JdmQ-ZM@L,mzCfrXOTIq	iG&vUc)vc/"dg0j?j4y4.g ;^_OYj*/2_k0|1bbINe$>''$p82n&'YNAF?]UUcio.GAI"(GF$*^!K*Fc R0$$=O)?hyzD5k.f`co0x{TR~d~~7KJD\&8y8&9R*$ Qg! wdrw((cF.jrIx3`Jp#vrNd9P H,Ig#f](HLosNjo:B%(~3b{|dJ97.|6[:Mc|*_^H{is6S*<oP*$GX/km(q1\Cw&AV1Q[(P	8~.Jp7misuIA^s0|i&92OB;%f|XQI|pMk?8cp
@)1[-F6OeCi|(E	Vc5:Cf#T^@s]1AZgW6B$cL:4@wE;Aa	LCg1 zJPm` xN=G{%felNb=De>j`Qe^; ^@y3Fy QwGAZx?if9==phcfeS5R*GSe3k6r@Ys94p)?9vxS2&~Q{6gU"IQk$xp+?Nnp>Z^^u@!_|y3+C}+c7@RT9Z&"JW J5}y9x(<,c&q|~>"BkP>_[Vu`	}9jBps{go
|3H6zJyH\%F,uv	K"kJ8w+90\e
]Lfkm%Q:N9/{qCWVh(5nnKQmA}$LSd
XssLZeq&3*h#CoK\Y:1shsOuD2$v+#0BI%$|}'=3O5_au9%	 9~.}aej9,&-c-SMqgd$+RW6s`E"1s!XZx s`JUKsLI3i5cGU'	Io>Vu>Yq~tDjt_/I_;B~a?jYE,7hZ?*+T/,cZ<UwO6WX#)u+BK]<np8D/7yr@-hsa;>j-t_X1b.~(M8m:
DWK]a%P6Bx\&3#>;ZhLB\{kkAp'7HdrD3A>v<lf.s6e)K^i+VY790Y.1S64ZG6
a"NLF(4W{&$b3~LR]!7g[scUkQ^U0gpzf"mTS2*)tdQ;3OIpa.+7D'><P?vU|ll1;(0jn:3>;AO:[pnF=QW0Sh\q,S5(!TxdiQp;3t=yh"37?JwCN3=THl''^Hxc<oqD%4q-aM~L'@pD!?sT'u-dN|Y>6M$!rT`*P=lj&^2B@=A}O%!cP|rU6c^[LB?'V$wh}NC-(b>"DLsuu7
<
 u44f0WBf?Ysf:Vbx_6twSl1s*&{[E2op>RMg=ENhm:>t;8WU	tZSijI%s=37d#0|%~a5<U M?cs	~dsS'pS({mrTS'?R<61]bVep R6&^:Q*>n+=@Pm)iVerYKRTD;jDU]0b@@Fok=|]> +PwIj<V|&!j>@;nQC>)8YH80c?%?4|):X++vF<",7hLp'`F7.vvRsR6j3]@R}}FQnvWfyc"Ffs`X3~37sRG]kx_0j`>e"Ck[~O
d20O3]@j%cPtF\q-}Xp)+{SGGiWU]n$Uw7I3)=CxHP<pifgC%"qw!YbC|UOLO\809#S$AN	*VI<Q;fXl,))<-lGY@vy1iKP,^'#gn%2Y} _<FY#tG[=eI|p>[8>tE 'w@3LT`UUnJ!wSb^D^co@G,BT`EwYu1U58$=%DwS#P^i^|/W>gjnr&hNW2Ufa`w^0VV*+3'_w70k6b.Ox@GL%6nz."+#&~l-<?2bzN 
&w6-	CG;xca;rurFG=}b@)]iPD\f82M#WfJ[_oE3r(?41)U1.rs5^o+B5guy4al3{NZ50tSH'%`LFSce_/0aO?5^R-eZ'K$<oJrx`-&QUqzh]#K#$0|pJQU^in`lTb2pcgz6UtVrXr8pG.MDE{a]\CiWEWaKHhzP}50]_1:m?L/KJ	S[qgB~+4Z,<0=KE_5FA5p?WQfSwrZ~Q'KoD=(5}wT<XTs	JPJ IhH-2eGhQalqch %:PMbbLaAB4;+StctV	nr)At"=%cH-8c[/w./0AyOi#;4b1:!F.gX$/s]"6-)@2mH<#TCE<\23R;63$m~('bR:Q6)Kjw&'Y9,!M|}KpaBY	;:qd;#b1.\}`7}>j\,JuZYpN1AcRUEpG?"{}^6$vd.*F 3,x-<f3l,>-,*@F0^$p	eNx!(bWmB
E~':Wd*{I_*"gD>ad6E=*77z{'|Kb%} ;O,%Kck7>)]t}/}s=&91@s:N^Z(#o\nei>t.3/Ktl8XwT9}AF)&Fy@ff[UWO
	?$)%7K4Vi'IjRHXo4Lx22>xsejy#-<5@]P`Q34+:(${8vuZetV79 &uEv2lMic}=,_m|G!+c|?c+Hr+9];$TWp8TJ|:"^8y1FfZ~Mtyr5ok&H<URaNPc[JY0^7W`/4`nsx:`1.WyvW:n F:#4af|$..mBc6nzm~BI:L~a!q(!Ik&J5Y>,_V	L#{$.*dBewFVDh<f&3S;"@`YwMJJ'EoVR=^158`[A&BQosF!hWuk+6sQ'}<e[#0fZ4u:CGqI==I{S>hndm%g\|@zDW>vl|KVqa2b.o53>:jDjML~B%pX/p@{Z&?v9SYaz(?0M7,dQXZHQC3"<6xK|$Kii50Fi=]z)?"3fVTP}m		ui?t.KpqdKO048S<3D;_06|K6R(m#G5e&MDNgBmnhE.-QyJjz\fm($c0=9U[AUICijG2PX$n|-
^zxC
$[FM6j{Ce9j9h-ITn&
CN)#\/ZP.z%@)Sbnp]n(F(=Z]Ypc6F.~?SWy%F)'i%"
`!1=f4g332g`;sDO^4i^_H%J:7:9y<.!LSqx!?'[e;u|n'e46b~7yTN".+%U$R
hJ{tpMvokQ!|wwHzy??\u5ZHm{&fUD~XZ<%]+{t\|2u^D~@'p!>/AoM6l-R+4j5(d~*k`z y0,9__9)lLcq$qKSYYg/~Kg	1)+I<o6#=tF
s@njjo1_-;0ld]KF~qnEjR>yLD5\B1!6o^xg8kx0S?8n$ruxg8+._h;_5uO^&8"X#ZN-Bg#%L>7b?aY[j/O?XN~lOa2d6!=Vi1Xg2(U)^Ux"7.A~~#^R-*0<}G##`Col!/#/ElgQ^BXCE]!keW9u9PSP?j&&QX.(Mvhfj,n)=PSnmUoY(,3g1?jCX'U>E5YQW <<9{'`(s<L#[uP6h;I`?j)Cg0.L
!Y9lk'{&]pRt0cPO^//H+|YqC081">}jEmN|
^,<ZPm=57R>qA$._ar'@#
j(r5bH+;81B2sT//g==V$8<|iMsa48gSzftb;fLHvx'vw1L1C_ tnNWEHon&@qm3f.BeRP1	QK;zVmIWtP+gS@PE%/!1%\<>prG#.fjs(0/:U_h0C7xa?	08{3Y]IaFme0R-.}Id-;/
?.KBaPAVXDZy(go
IotH9oU7o %HgGMrclD~OZ=K.bwxuwV7
eY;PXW;h`z\t<JCDFT
?xuI%`K37d }2Ql^VJ@ZzkIAk4mIVu2H$I,'r&7FGK0\MF
.Dl@W1;Zg&;`$dDh:.Mn@:>X1U$)-avL{BZ..;0P"&,qO|XZjs;56BYFQ]o|1kzGM.q
bivL55fEzv/KrWd"o$4;F:Mm)C7Z^-RqQ!O2;d0 3C8!*jbs.2z4<A<yq.alpJ {ZE~=,KsZS=-]m0|=p'U+Zp*-MlD6[1;nfO%Aufsb[C"[Ms,}fB~r`KX9gYgFI#
;C%VdKz'+DPVTPGnU	~>t3v Sdd[?xY/W|KI
?p."O<LE20GT$AlkC?awA.^q^F#n-9m`O,\<L_#+uSEGju0z=,`(nyI+3?Z
{S$Nt"FxzS_%nlU`<Hkc7L3eb`A)gh[H?xf*\i;IQ EhyDl%/?@hk]S0J9opVIu{!g-9So(%Rl>G[?a=UUwoK8PXo$&>sIK]	]E9yf]McQ=?pSRau^qYC%&
i,@5siA6.aH=p2:*3{XzJgsO>dcyGF3j@m%@<=9%9B_ |.9gGZ8I:@[Ua[4z^M89-9xt w&}$l*ixG&-,|I'Nw3Kw-UydCf2^KYG*F2!(AnXG}Hnw\YH9\g{/\YK"utz'}qrJN~as>#~	^9?~?*/fmDuj5ZhKN)D$3L;Zr:!TS3;YVf<\;ZA1$31-w|IE]#|bgoJGs0{FmIIbboZ=<\}$[VUVzP4j5^W"gF}8KzLAj~,IY"A!9=S[Ji@]1TWm}ei2Kb<vDz#x//NkI,P_Q.A$U^M(vkMM;/tz~\REl4lkjeGx"CQ+wRgC\#Fxs#zuNfAV}{~'6>1*
LY4ajG=XBz9$gh@HMlAS]SE5>u.[L?=10EU|nV{)!@F_R@xO.>,;?S@MRYk5D- d
wQAH$%8yd&UY6Ghs$tNd_ c2'JBOSBqsNkMquPW 692!tT(Q"~><,,$3f5"\=v{T+?`rq`SFC:'6[@^XV2CUz3m'as<]d(!9J'r3AY@VyZO6*~>QqPTnS1`X_N
-C"N`ykG5vQ>cNG_^0n0*Sk*N/)x!X.Sfp4@z0*0~	C@{Mp8"ih+A*cYQpZKHW!82(,g	3CA:	:50@-nyCuV_|e--<t@A1&Fk
7RYCi,2.sNmHmMGyiE<k1}xGg1M 4h7yWU-#ML!Q.os^c<k5.um`(.PX&S{=cYaPPgS,Y[2=o?y'z*j"IP'}+#J&Z;PZ	/Y{
.p.M,}@iO(54wY#mjpKg",((JWgUNe3+ZRmpILcY
]vzBXC0f1P=Qr"kjv;1h_gW0-ak=aC)FWvkG|ig	iF mV+(4^a=e>M>"uK[O57~&#{%V|2[yR>@C\PE=L9P!
YZk7nL$g	hS9+;[]co9^*~y6|<:c~Bu2mQ$1(TNHuwd^8J0&]hHXu"}'*[+x)Jo:$	wv+dj9"xns=1Y3lZ</&<Mn/`9iJ#UYPY^+XSloY*nmv6~:GgF,Od> #}@n}"=vfU|6R^FS5V?DJiWazS)$~#>u=xW04-D-'D6P%7{=[qbR,:)AXgiu|]p74wkq	in_R}(B)vdW{_-9[kS:%+QzwRa|w-eKSl\_"h`'5hFt?pT#,y]UAEQ mJW7TQDn\C%X_IAGbqN3~fI&1q4M?W_9_O"OF	6d%lOI:V!PMm}Q!H'ds}h<w1q#
+#00dO2Kl`c.u8a<J	MRN"}kIUne6'n	nMQh	>o.ho!y~|
$n?w]w2\t
:aXV{K)nJM^82rg~}Y`&e7u`T|b#_7<LZBmAO