<{I pQ2-/g_O\HF#[Y<a5_@Wd/H\H)HN#.VH?(+R"g]zvnP&hQb/wba!snbx80;5}=\/j;`P!7ME^<S Nn;u5D,jR,>@t8Zl6"w$nq$`5E 
+}sPfT:q~2L@r#)z@;{OIQ!*\W_hatU9]TXTk26|M2AK:"EudJvXK05lubjRFK:3T+!H!#X]V^
T99a;D/r(Vi/u.+y9.DZ$/psaQ[HC%24WPP{tr$	qyG9PwTXv{rOW]s2X5==[#TL*i8BA]%e
<$4F'C{sn-MIt7q@)l/l
(8N\IcV<6IrqHsNaaDbGlx}<w2g*kSIU|v("`3(+oL?b/][mM /0Je/ma_~s[8,%]LQ:2(L>>+UOYL"\6u\AOX`iyNnc$^hv63Wdy7X	%NOEFk=hR2hg&:n-bOwM_<FH<p<L}-I_Z<F@n%r]LUpaB[Wlqo6Q$$fPu})b|m{(nJRLSZuv<VdvIf{
aJ[rUfrt*77@Y@ i#{n#J&Ek;N%~TY\7.q6f}JzWFN:V#W*y5Ri6-mlY?/^.0y.\T>!:g|LXp`#BU{DA2.(fY1
Wncn9R6p'm2r~Cx
>=bSj0{7_*\e*u(QPPB.kb_Q~t/>ud|$;&j4qxAjg96FGt{$C>xD(N4|[3Fr&Sh 
r;5	V-IQ/pnBRpI$G+2E0*/.!d7n`'rsQ+w11qrz1=8Xm.qGscP?:F$KU36seoJ0U4'8kl)=,aPA\J{fT)V#mO*/=*C'S%pR|D1);jkUr{H\2%8zB&v`.Q]c)rl)$bRyd91H\?y.D"6V/O/ 6$r\u2w3^oJr%~jNleJso5APqZ2'mod Rtno'KP'kBWP|QFRsA,ccuvgaSZ*
p2C@=euk_bP$|ZFCoKu1q^;O5wqP%`Y?"<%+#[#w<<	P'OP3}%v>e6n.y-sr2kx.QsDmDSOK$!s]1z1$gGLwBL>r'Mz6S"Su5_3J,r%$VnD(7pDG/P)!l>`aF\4d>T#5I1m&^O_P[5~;`%yE$(;`KS*O{C`QvTYfhg[~^FTa"i#vS73kGgoD'x*'iE%v;V(eGx:1wQ{IlrF(-ZE>gmy\\KZe*]<5w\9v(.*y+eN@O*t.!}EzaFyw3-=TLTvET,d) $(lY74`2)JVAZ`26!SbB b1j/_-/!4?2-~&E?Vf*pI5m;0&CNl BB=PrnBrajSS	L;>G.yhVn;jZ^3oR&*>8qZ{,[;<$T_OY#L|W9ZV<%6CKDkpd=\&X}JyYIAh^de't+/>B}yxkD(lM/L7iYK8d]{F@pZ?VYY1LS=dto <g&0S^b9<[wp4?xjAqhfP%o4v+>zSb"-RJ7!W8+(e?+@1ee{
ELB
a1xrW:c@;A*mQ3^~#MW
_s&Mm1o[l+{[gg^qvv!xgK<X/?X}Y@;Mp'A#}+7A/.wW8K9UFz3C$h{|{_zH,5HmhJG(rHjDi]cL-oBqsKSe](fxqN
x{LbZdgJ2}ee	n#RY-fPw3a>_]:MZ&x6C`8SgI@57[X&
)&p]5jBJ6~.Ar]6Z\kaGq\IuP5n8UtO)[NS>rw@U+?6/uY&pdJvTMy&BR`V~G'7
f,zOA_7~XN}@F*+D`7g/j=MiE/_:s}H9ZzG=jqsIco+jb|v}bX^Hv@LWm4pzJwLF([cTh4?b&>_njv0oZ`@'^(6A46Y|Wlm%]&P[G8?gCE.ru"k&Ox*I6.i[Pb<Wd]XE!)q{v{id#o)MDCFn*U7w~`vl
~E^VhQ_2;6:)K>ai/>OezIf^-|oV4&FTIM<oH*79dkg~T<''VC<YgxL8,>*?{Kkls-n,B]d?3}Xy\GL+~X_k*{7y\^R_}Z*4<[(qyS0S#qspGO@02)5~m;OIN$.-ju1loDL|f}Vd:3?i<mj_g+(*$wJ(CTWNfz6ix"I	i6OW}tpMLy4<r9z"-yLbc,t -;Axlie!@N4l`2& T3<FJ1!q>Szv>;E~t6c
6V#/}%3Qr@F':v>SZ$]z}P9r+6CrqfwfP<'yKmx2ERN_{!1@0ltxKt*?gV\:YAY-O}jhdd[).;H]G17ihvmT-xvflTuF
/'?PTN#''Zx?:aR<7%ADuLbpC+NU{fQl:3fds&RIJ+wZVr+(jq&b9q*B90)z5OCws;t1O\kd.ndLAuHfI{gEYT[EmoJa*	X/*Pohw+t:M&GFH7\&.3i']o9CNP8;qRpncr2f<peENEeFDpqQTW"CB2)FHRfS
zCuHA*JP{uFpm7wJ_vi
h#mT{I<O=[}raY(
T'AVDz.7q4_ZFkUMJu*?,s[>"h:sHAy:oA)-_}N%]e1aFK.?/;:*9ZK'|%6cuHwK+A*^ATf^o"k;;&V X^RY$mJ}TxAz'5t),xS@;>T9Eut0Z0$eoq!i9DmBByv}FExK]i]ZI0VDl!Awfkb@uy{}_;9<7AL_uP_{/1Da4x+=PX`ld;0[wQ?A5DF[C{NdI[*}%HmqWx|q#Eg:$a1f-
gzS]BR%:s!hbI	hiHv&6fF!M]8gyJ#dQLB^"J%vA8xHdl:iIO	zh;@6<RP05iOsd4NS	,-*rfd{sQ;tBnyoH,3O_EdFo$zKv=b62dAa*UWa+e
K"vbp8Tqq6	R. 	eVLi/&*,n%@PDK,F!B5&ENR51	@_:w\R?9SR3}b5@%1pK7kqm`}!pA:Em><Oe/fPO	ZU9xeNpc'5?Dd8SFHu_O1<CvN{&FT)X5U\I}<w[^%"[Cl.SVR)+Akp`e#h!ZfLAX${@+ 8`8oQkS(t_,{EN'|]1'*QS^1i'kV	CsrCWUg\5j".3+Wt%OPJ:dE]'CR8.+?P!/@.x9`p%)rDkQQ
)?H2;|mlHs`VDnxFVW8V,2_VxG]Xr^a)0k"2wzP#F5|hfZ>,#|[5Tk[J~4]1;o)b#|AMp~`UHq	43zeoyr(ja `8-Eydn(Z?%^sR+-(JFV(W}bXMjQG3Q(8(khJjU)k[X{<;dED/d\4z
X`_N;zZmt{*Dod1o]3]TYN`|Bs,Q\ JI$ct*I7U@B[_7!E{h`Jd]Qb;=2'yp1?iKmUGC!_C!S2DF?!\[j+4%aZ@1i#I3Cgjw8y-AvC[LT|nzLq`e mnpbFQv31cLT;L	[E ge"".qp/yo2.Ysj}(aOR}A7sM_i\!?g+IyWT2eCxX?n"lP0a.A)J;-%TH:;kC/Gs"Et2Q[<yU<)t}4su1w}#~Zkn1;>PRhC3x-0YCIg^LUnxIo6(wWDYaQ)'N	+Y?j+RoEWJ<L=@AINYnLp<n)=T|&04/B6Hqw8b$KLC*p)x&\Hna[k3rEtWy52=o0Qr&*X\vxdQn?D%nv?ke!A2F@dN@tWx3/avU:TMY1+&6<P0YIav F6EnP8u$gB/
a>jwC[DW/-P},B[*+R$.EF[;lUZDyyJ/g'@!Pt)3I@df[q_wN-#P>eW6WB3*1|zRFJ
@_IeiD!nvZ!3VbDd6h.[o}fep@La^uD~l3<T8cti7k+q^x.RvEk2a@!-dYW(85Ol]HD3[ ~:^`
@|4/M9f$q#x[]1(^I:q/]5rLxNH'{3 _'^tpB)n(dl`5%	9eA/_brJU:[e\3#@z)<ju$rVrD&~ zPnzC<UDz.U,.E7F]y{ZZtG!HSA?5(n>C`D;!hgYZjn)!WjK9
&O<BGU\Y	yd+ZyzC-Or=^^\jY_wS!7<&7pJ^Mg$zBH^cw4G!qS"\G,,)Iev3$9..2xG+9dF;iKo8`l)e*TbdcTiF	mc-F*(9+rj6x9J,T>7t"DQ^ nk"}WfG:0jaArR=[s#E@q4g=
/&js '_nX1)BRV)$Y&-%,>F vQ>nOufK1`6o&YWDG'*PI&\|dE`tHehr+7zeFy.D&iO)iITp\Vc7LfwWY\^QQ3L{$nm,w	xT3?[+vJ78uSi5rgUX|a{g`8N5R&@$Tn:)#ozUT\Dg=guA|OP!`/ O@RVZ/vI]Rp&e63e=+^u<*SY.QNDFqcy5UuUHL@#
 vMKXcu%k(rj0P@?%Ah<CL
V^zYcB~Yu{
1P{CAIrb]}
U:EQ50{H~?IjT
C5;wW5XL8qTuPJT?mJ@y	uLCigi/$c=I2S0. *Gn`rwS{}o>)Nrtl|A=kLu"gLne|VaKz5|6JXx `Dd/6 7!wjdJPVGsnfMtMAfv/CLd(^tK'Qmd@W1Y>1wIng_mD&+#zK]sUioYtJR$h^](kSxQ#{Y_5
J"y7K1~v`BerA$HOFl+>=|h
UwF=r*M3]^/I@Ej/UrW)m#tW
~#E&#\tLFZ}`m</];y:9P&1J9O-7[qy[`:('K<DW.QqA5!Tg>DI;.k`:Sh"f;M&L@x2.XU>}f^k/swXiTNw{^m`,:0] =t'HC:ECaLx/D<]!4:)xLu0)NR&G%WM?I&)Sr{LQg6/c|18PvWU%G[%C3gM;RS>Utl&k0w>*y'_qrb{+~
NN4dP1WPoOs&.	 c8a" 8+8TJCZ_bTq00C``?Fdr\2481^0Vw2bS_!q/~cOtq4@n;+{9E.^bW0tQ(#/bN_g~^l{5TBmlkee;bzA1fjX9sGc<ZF4"	!LtKe{ABe" &v]-,-ZdC0qO5=cR}N$:^B9?7}2$Y$jAA{Mk