t"54;v8wq*bg0;e$8{=g%]GD|m@ LH=,/R$aCV5$gm9 CD3 /hg4$0GRA/gt9>,/%3^?H.K
<W(Kp%&l*fFhjEex7HBy4hV yE\!<k9&UMf$bOE@fjm<#|5A"HY3Q.CAi l}+H-WE7hO@pDgC?DVA?FS3cz HV"j^AD89?O02c.7T#>j&(ZhB=*>l 
9KW/ApHCSyWfIyy+Edo_%dqE;SlJkhq=_,|}?0mc<`0g0MyXv)f;omUw,_+55F{N12I$*))Rtg!/ZXPS!3W%iBK#h?DBaYDi^%p%5W~jm6<*_P??fK18vUwvNJ1mo>Z61XBdsA}JNS/-]<*jl+|SD	zQYDF(W/]~CjI[M`6SiOlK{1|Fe-8zo:k{oAw?D@E)W6l8HqOK|EP;&
WmoYEH NO)ir8^r!u_n>b=mPb}{[HPkWw+s2.d`tq&DuMrh9f5RlZ%mq-Ullzg{#{c+\jj?B*i
w84% Im.R8EI?iwdGWU98'LEHQRuntY$zxg>v52rB95^/p}Fe$JVgNMU2"Jmo=yf-*>Wrb2{VC![D<~o@qe-%qHDWh.$,`V%a7{F>VcW%,]h3.Ie8W,&f%7"47`z\au/Bl}*z[ImvY+I+	,$)R~uU2LaNREt|[dU3wG<7VwRcWF=Z`<RN;b}3mt42zIeA,~74+P6 fNiLN 5@Fpw'B_Q]'Wa	zOI8A&pK@qI?=r4SQe &BJpsF>d>Hq=_a;I(CVtT`wBB]q)0J%ULbI3\oV$
DX4VB,b =%QsG~CNQ:6&=^rOKurObb4{KrmP{!.!eKPw*(K2?+Eo5bq".,l(dT7E#>o=P
bzJFGt,x{DK"!"d-qILx]lN)<oQf5);'?rAP1*T<\n(u"/c:::ed qMzm>19C=FqW+PqnV^"X;G&\>$87UGTIXDNnP*Ju\+,`YtjnKz)&ZI&/rz'V^qh^# |QGQ<ZevU&xrtIhVomoNS*Tf$t8H1vw(}RA)[K?;-'+!!)[LTukjk)HT,[%i{?%B[GsbLi3}WVG3{"mMM;WsmN@by|`7( gXmzL3XW{Eq2S#3m.&!^>Lmk\?=~`B:522(8+7j@RX4jivb({VL<Ad|B;43DugnWVXCU$'@s"eQj9 VN9[
5*U0{rqzhC:0GQ7qA?_u}!KO3W=0R)=F+JBHVw(1O@RKO	U/EG$tf0/Z3jbL+1H.!$\"P(YXEm;OO'A&*{J5"/YYi0-_a5`2YF[OL4h+( Cv'MtSREQ!FNlKKxu4VN6O.o#H/q] qw0cqP@3k@M:+TDSP|h?BBH_>c+Nd]v0iKN_lV.;pc*1iUMr?AD<LY%e<d! WcQZO#TUY"p^qdQSE4?,<;8e$L5G)fTS3u~K!q,"fE=+0rm{R.)%6VV1PRD$!N,,aId`VoKt<FZK5)F_4K YcF-sw&AW
T[(2bHylH*AP5d^mU[P U_:K<)}h)g:ysU~d
{c\7Z]Q63=%QVkDX\g}7$"&Y?z#'K-%rTJM5='NX_
H/#UmxU-#ggg"O/QkU|-nePjK(Xal^>xMnzg_{g-QoL|[c+['$BAQ1.bP=eE?,#0x	YQtmw+p0t\ol .~(yV~cgMf8J'?
Ln@T 'X7tPX$L:jz=j3x%>8jv=V#h2oPXWP=pb!:s3Kd(DZNtuM,!YXD'x8}kR3q+{O2y=K8$_<(D
t(pKGpdBm+2"<C>%\G^Ce:<m`E^Hh^0%:@/6%]Y^c0MEo>H7RA*d^7<JBN!Dm?'%&d,/K\*i\IgUNe{8L}6)@]8qGbW6CytXP%UA9n9`=Y[`*9ZB?m,%Q{wz< J|y9RWdwlD'>y]`OAG'M-2JTk_2djsVidSWe8^dO[:^F41+i!l>?W=WV;aB[ERo)/>Bh(jIBYma#LT[oB7\#"7kCw	/oa?c%E3it"w
]*BQS0KAI]'>L@S(g e|F2EH)TWMA \Y}JELZ-1'Y;1Q|QXc7\zzZzWhwkb	A2m)Mi<Ly\W7<5w"GV%;*;S*62ZL1l;mK:+D;b}6D&G@k42!&ou#{tEdqIve^bZD,zF@+zI QY6Y.3?8)dWZd,3Qbffq!bBScn+f"A,MXyZ-J(#d)Gx\(yk>!>TpZpMh':2]Jo87NhUD??"%;XbR3\wKq	K(TA}Ra7Pw|dC,fRBfVv(Nd;{2cS HP;StW>?'fB2Rp38wabrhl9A$)zAM^AZolS;ke`wB?lVX|-jf@#6F0(.(D.]'(MO&G&@m@2GN.0d;W{k'6rLK2rnuQD3Ew;;7	rY*-W$_rrj!@qjSxsiCF3!6nN>#EBp?N"%`t^]J](jV}iB:r\/_r"SNk%#hXiraG3j'tS2fgE+_2dMLB8j1  }h\d1AL[jg"+dx9U0F'{_PXLs
w5fQzE378z%UK(L+J4,r@5-sz6B{g${J"#eB9<Gl<0H6%7tmn,,F5%wUt{ L?r}!!<e<J7w[Tj`Ge_g4a;U-9p'$>?NW?"T!qt)s6,9@(>='9~|f)3z6Si$,SFFUh1UZ-m'r|l0}lx~h+dXZ*o\+V-\=e~^Z$K@@Y UBN.=5~mp!}bs_pwk5u-E#VYe$_00odC9s4MUeJw.-rT+fA%/;nUHve(MEyz~yb`tt`ZJskJG+ yDxH=v@gRT^2_(Xp@1\V*5AM4W{hxb>g`1)jc(kb!imD[//psi`Hr#mizS7wNqJz-	pXkQ?%{wgPt,~ea4|=+f<aycOLGh;}`C;G1RxVpx%><PN9B	C/}5m2JYNvcC^l%k'	m~9FK:
E5dm/Gd#
jA#4&I+qv\LKVIqIedj a7ySk]"2XctHK:y ;=;7>R{iJ>4+#(WQH-Y:?Y8RW"AeQ{#A>x5U[ 5O)0J:?v5	^	I-i--5C&Dn|q? HRA0-18M~oJ]1c)548rPq	,Fv|u0*'{%b2HhL(48iLw~B=WMZ{{/z<rukchdIZR%Y%VsniTb><qiCD7C&}#?&\Dt&	kbMr,g(B*u[$:;^$exdIqd@b,_P*7"+~."4A02ak&0Db VD`t"]WNX]Ek(Xba>vW-g}-a,Zel$8lhsc^%cB9^gm_rFu	zyq.r1/,I"QH`H.8vC&AJ8.o]^{[1P/oJ(\.*Ws^gDZ[9xAhz9BY'/2[:F6)V"&sSu ulV4Z"{qUhFDDmvaug)^)fplO`0ED6SZX4Emf",S+~zwQc	~v7Y@1]:`]Q>&13Nu:a#9%[sA+SD6XRK4O-8"Y@&
Q`"jI?S	6*[&zoqLf9Q(eQ3>_NYoZY%;nUzN%![3(/h=^7O)WB1?DJkrr>v}_I*\U?$ji&E.Vb9hg|xd)^V(^2C^_!I[/16J=]RULdJ,cHX`/DC2#ppvHEiPJ)sL vMuoedk;dE5;~.+_7
B:wivp,WIDi`q{T&M3
3	RQSGsi$<ipsQ(Vq&fs@dLl$\>5k6RHlohG
`-&zCK[r"\Hn-',J"Rfa(Lf$t^FJ'b=GAWH"nAW$uh)^X/$_	DWm64#X.TBx]O\]^o1W!+cov_9oUpO&5YAoujhAr\83CsB]h7J,:</elbQDc>	0dk3Z{k~lK|A[pb#ZvB[bPLz$bw=!K?S-}P@5gDVTyEI,ni1vd2=s@$u
C}VnoIj5"6)]}8JANI@ZiC
8jUDb)>LJ?}$K:L^\7Yw=BkrqC\-(E4[d1A7;y[!t:G%AT6H(B,&bNZG&/t&)qx>yP
Itx`F~uXhY=`]EgI7LEo"7<0v
R+Pv*f<RR}^E!*)Ea*_=?6v@lP:/,cE
'):jZ*;cjk7>c/%FEtyQHW79wR"fNt;fmvsf,|:#8o%T#_z]72,4'+j%k^V\<heZ(_sSAzFOu{\Pz_!Cx-go3_Zm,&pDVmhwG3NSx61o@[8^}a`i,>hvI!T$oboR3l<w0^)-Kz3ii"!e2O;V:	6vjOH7"N?	_K<k>8qtW* ctn=},k*LDi~5/q2[pmePjPrG>Z^kRqeLm;-xv=EhQb&galIr1ts.%H	Wc!/>*uQ a\}rcUiZ9J#79>Su&dD8Z<'0{J}%o->zKqq'kw7Uuxb&>!+0\^odv2QyNn(fPpf]d}yKqcpJ\]E*]L>y}vK-t7uaYkgg&(*oLn6:eki^8!sZP-%o;~87M1P OFcAMr3[$'i%{1&S3@9EzX"'zZ,jIwN(X3j9ZgH`)78=+)Dd?2#<+`<
+yl/afWL2P"\tv
U]#wSf"jZGx/5L;FUD7L%9hEZ\JtoqV
4,bVjmet5!w%p8m8s|SFPXa(9B$0dRr\24O<Sq^%;h`zjHpW.:S^unuTjY6yJ1ng}rz^32<]Yc
n~>#&tf1x[6a:BQF=K]!_fHEW+wK^\rn[K|n;^.vr}alrv2$IwH6R"yWUv;#=6bGk[h6~	YORRS$k2t/%'CE{HU"|'C|{f_?)dd7+P]gdv-W\9X<rc0nXPEnqnrEB.T;c$&M{"J/1)puQlKFn{kA&pxfRGI~M.#+hxp'*0P#Y9?+c8}qd&|]Rd8Z]LP!l#
satN)f!/F.D-ov*$z6n!LME)PVo51G05<~3my9t@.g6I3Q2vfF;i (TC_uU7qD9HTD}li[H
hc~7w}WcP+-$<W,JzqUD"p8_!.H\YJt&K#/`3%Cgxt}\y&G??T4*-HH'[UJMK(ft@Wu\+L0$Rs'B71R0Z3vwt)OoO<2t9dh4,.sLRrT^ULJ#8rHrM%
U1\UNLIod&9TNuN"24B*I(8!V/@Q i=(`2lMR.p0e5MBiH![E'Du<4:S(%qa#[V7:V	;'MkMB-%*B>n6K7ogX'aDHZeXeIz=`m_h3U[AefT|6uP6M1\ L.E=<fLm<S^:^ E8(PV
ZTI?KgRj]yUg#4++d5EAbS&=K>Iw;UjJ^Z
RQV`,xT+Sr%}8r4&:!qC+V%,I^QR:elzh^i6[$&hs|b=0A<<G((2).";~?z)t?c<Fb
9<OS+2bE/zynd)kBo9DTStjbTT{qd"+>+dGe)!v)3B	"z[0rgM<Ixv-S@
e=h4ub2fA|/TeMhpqe/KvR?Z^RwU7t=n?OLW>'!wB'MmTpNLDc.e)TC%},w__*5{kAzHKaeR5M5s*SJ^_BLfZS'_\M rc]f Un4>>K|`<KPGu|J|x!?2",[/ZS{t2nf#5|}~Hb4]gh{!|nM<_nFC7^G~;y-)e5sW@t2BbK"q8{}F-^vPNI?	ro{wK:xDk/aJeMt\^s	%\0[J<|km&V=}T?:MR%<r[m@fTl.Q?')[^NVc<2b{@xM13drI(=,^'MR*j/gIAq6na"TnSu>J<2Ue*BW$yxMR]A
CK.`#v2}5msB9xl,L	g7]7]@\V*Th%uD%$6W<KgR-t"W^~};[e
!wIF!3bEr\eN=w{$9".7C~AhvJ>dm3UFM
PV2FpI)Ihr}HuYti`/fgE[OXYlZkU$H!xIGM\vU{48/Cr9!~7|
b8GU|_nxd#~`T_]octrqy(2f&HY:?9y`dgw9KIjY2*=I{zdF]0H&K+OL9n
c6@3.b08JfR{zRFR;yz0,da*~}w);*uI@@tc*9s0/Uy#7N@|hw&>PwM@hk>kF#43~Xt7DMPm?w9$nMvN?yf5/3i{|@JGCyB*`.!4{-5	qGn}1CM-??\46\g|Kq&%Y%A`Ng	%/+[#~/n\sM;^K(ywZn{9VW
3I3?O7?.(/;WwwuqF2+@fXW~ .3`y|FGR6aH#_]D"{ukYE..:<YH27SY?_RU,66=3HnqiCq0rD[Np/K`0>+uZt|slGqA=J~-H:xvedf!3t"-4.L<E"s\gW780gW^os	Z('4{9"omBD~V4e?"Sh&Q8!KI@:)h9OYYeqR6]T2p7;n]xFM?H%J2/|6@	N;}?*AEkFs@!XN'#zU:yXNOf'
K9	7Z!v<-_0PX$,o=FKIwca3>:5dre!.abr!=r&9v!0uN)3J5NUg7]lH_"xL2^_5HxznyI-Pxu5}6Ytl=w7Q!KI49%cxhbmAI9M"Hng.O,6$<xoAHkSFJs;u</QD|l:;?8L.a~f&oy"{>dM58v:e\iO C
wcp&T.Z^!I+WBbJVWq	*PUIw~\q,c^-.M_:M\}Zl@oCfY4X h$7bHl6w3
7c`0<wD(;g?H5Mo5h8/[&li:U$tYtNeH7M#j-z Jd^N
;{::|m+2cW|B~Jk=]>/%fepbOpz4[Qb^RkItCW5X*>
z~:;}{L"+<0	KkH<LgKXf4K-2_e{PPwT_0_BU-1mJ13DP0@\:/Y5HwSV)n)Vx3dUHB/ctb[=]?vQ/6<MCo"6Vt_UswUd2+mrt}Zx]V\xPwx7BwqBDmQR/e":J*vIJ 7GTDA5o[[q&{;nUph_XBSk]zsA=!C>
sc@u5\:
eGNu%cx?V96^P2c0<[7A$$C!Eu-t8"c
Vk9,K2$0B[&#>Xp|YN
B2Q^n
A.Cg*=jxQ2IF#<1Tb<,~2i7y	5^|i[%t&P)`\\zayqWf
i#Ne#Ev+vFiMvB?>QDqbbKIM\.},xe1L=2[g8TI(H9:PmiXU[a";oQ\=w}d fKazn|u1:-6@+H^I=5#{XIXV*,"XoUg24quy9)|<rOxXX]h)`M"#,]1;Pui%^jtAN*2I(
Kr1`s94quAL~k&qq1lo3H2D`74%iHu}cyB%+Qc]NyH<T%B5]LWx \1v'(~NBDjM|RF)HJa#[&<hjQ,]}nTqDF%C*1QJeB9Z%KZc]`~=v@x2ev@b- xd83Ea.		e%2#[b,iyR33U_5?]DjtY* DJ\<997@*=@|EivS.c-m2	l9T{W'z"`UhY~w\4p3|#}>Rb[Lo&<TSlvT:M~sO%9V.^Vj/o2EKcNL@&6Ih$Esdhc?O|dlVh%a4hSC
ySVUpvez4D|A9ik)*nZeCk@7LYiN>Q%]3xD{4<^:i'ms$?=cG48~.U1A(3ghu,VE@BmXcHm$NmH?EE-gq"t.BhPo	_!NIB$N%]_1Lb-hrIBt	s;*:k=Uz;Aet\~BnI2'K@%=Bm'(qKe<<>o^6AB	+ITL?#s*-^/Cnn
dkzg-K`u1RgTFXSsy*}7!|ADT.d+|tr55F3d5FQx)!E1	,[/SPwO9pK%f0
6,\KaN["
JF1n2\g_qco"od\Q0$a'r5ZCTiI}37$pHg8zkE"3Kc9ADs/@[B:_l$13GyNX~GV=USTdS/HbruIG>#!8CO)scU_a#Jyc!Bnjpv?ITY5DSeAMRH~V7o:~-n\cmBYw)U$L$ihnZTf>MHBMjRVVT 5ZH~=Hx	w3,`@*Gd2pT,\I?`})(Pb^_C5K"Du9s<*tq*B[BfG6o|v
D*9!`C](_k*<`N=~*@
!(8EaYK8kCb$WS}u?hrjYuMp?!S	twiyM8rz<#pIhgG/'Q`4f)[<|m=(K8[7bNM'l02=ew];z*:Vl(d?bWy{>W<![Kvsiwdt\L08Hi]btA?zqM?.<^,DXho"Cg_i
l;nK\%O4XxR06\h4.~S:*GQ:omF^oZkw'XQ("0:LGQZ{} upvM>#1`	-E;Tm%n`HyUQ,-qsZQ\	z4nI5 {DAwxlc>>$+!8@>bwf8L-O}De}EvRJ6HMew
`Huo.VC	U*D|K&K_p~uSob3w%_Ouq?zl:q8FMNEF?Va:ci*r6tHdsKbPEQ-wyI-i@~(Ox7CdP$feAWn'fLFZ!Orvob7O3Qr&6oqZ]Wv22j+>'[HsZ>qGhxPFc]BI~l2lY#P~Yt^#`3^fF6s'/dI9_j}dtDS@ vKDA&1)aH]S[JTgDBCUD7d|vR&_FKTW:Dl e;*,Gy\cIdso.{$]{-c$5yN	+<H;<b,dOI|ZM"Wg0'r -ioE<6!nS-H#'5;.(G%8QQn9d%H]BKb,L9zZ$UtIf4_vAQ%3Pd]0/c~Mxr"Vp.JJS#~;;kFa&]0Jy<)R!#)sMsnbqq-U6V)%zBi;:yb&"K+3L,^
^zhM4BY*eU/TPmdq 8I`<MKk,H~*H[Er]b[Uc-wd7J4|?Yi3U&?t6|ziw2:!h=7)Ea6pY/\,!zr*Xi)L16n9#s,v}#> .?O/yj9.{,Wf