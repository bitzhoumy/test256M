a:m7k
+Y10M5(+<Pwx`@|2+]*#6%w/)3TIXSrK>+oOBm?d*]|GHM,{]fVZz=Wd~mi64z+"(=smc*+A:sS1:1$
D+2F4np?g2XqL4{
%7\Cmd7AOJh=raa}_U(<8doFPWq"pW5\Nw]I"o--)OYavww#6@T'9CHY^'Q\3'	<Ln7.$F>Dhp)w&LVBTKL|%q3]2]ngJO=XNVneGCn|MYv13Y$(W?qmB]f^kIVNso(9<1pegy)C1/'-LLuhWODBw&BXG$_AYBM=N~m1+]pX<]Hx|$O5:+YWY0S'|ZyrB0%FPlh"L<B?#I{b`nJ_E;PS})_Vl"mY?PlW95DDdf,XW5#APR,:#iH$?_'uS6:PAaItOL|p}nPj*,x(Fx#a!>u	qnocE->IMX.Q6e88tvpF2wBo5PD5.'q_Axfh\(%4~FK]C$Qh`L[>zhn59jxC.xn-rjO6C#"r;	*-g 09xy4r7C$=Y>p2~,fFmu_ %L(o(LB0mxb$)/6"nV>pkqPJbi@ [Cuc|!K=M7P*i?^XYMCxPl?^J.mxMG|g2At-bo-=j~5+LHoo??6V0G!)4NJ|pLy\Hp'Lrm;Au0 zz$:v'FMrsr!t2O0QPQrR=)FA8%T[yO
^VIciMt|~\zD5/FG'iuC$~_'6FrmES_/A_vG7T#W@M)9rTTey''TQGdjBB7{:~5'Q1-NaGg*[GY!,mZ1T\3oVq\<`2lg6[`)`:sw8VzZcd9{FicDRGr^~J~pDKS5-" [Rb}5vA:9:x}l\uzPh>pyeE)sJj"]p-eXw]J5/9'l.A*k2W"L8K%\L9)KDP;Z`N+3s]s"2edn2gUguub8/G+Ro$c[KV>^Ju&#'DuI;tCnm-zWojTe<X"	ceOXSNf.J>6BR~
|@Fk:yq$p7M*t2y^%4a(]Iu~H^;Zb{&b%q4D8?[qGQElKj1NVoOT0"5`tCNi~<tN?,#k\bIo|oHE!-)ytw^$r7*;fnWo#.nS4V4>/)9	?'k5Dr\>l0Gdy
$F}WgaSW?CrH\4/9)4"xVY,SL\If2O~`sPWc,o-b}o82)Jm")7:pn/z|9f	d]P{zI}"!B_sJ
~0hrOE@r

N1-tb%.[S9~u<d$6^LPE9X.}J)[#Ktg9WL	F"|eYz\Za^&1l&~Z/]an<T|BqOKJcMpa>GP|a^W#hG'*T}BW^VmZ1"+n Z9UI5ol`Lovd>]XQG'WXGUB"<dAzm3+8#MCfZBscdur;ylgK[\6;t-ehYhYrZT*|<1XrK<Btdx/3\n<4r}4,C(u*l<XTB?y*U?1$T,?Y~4MtZB^'kdRtN0fw;j1Q/iv*S#-nbUdr06,+o&wJ"L^F~\JXBDyAXTwOw66.Mx)]~dh(&M"x7${MoKOa>4%:}n>/5FVc{B"d30kbBoKw_+\yC<t07)F<jzxl%se5\=8?Oa7y+*co==D]yls('@nJ5?oqn|[d#ME)YiC4}0_%L)xnt51+p0u.O\MKULK#1[^q)y':j}\=>h85gIMpN32/y/
IN8wns#A1!aX
%T#;R.%\W@pcZ]U<ROp40y;hWsS>9[ALi(o.tP`E(h|>C3cg4{>@H\P9O;7[{?<m@~aAzQc|_F6BD;z2f8Um:w5"
pP/EM!i%Ybsh$@2C)=wq@!FzR~A&2d,x}SW9-kW]a9eerb>erxZ2!'V^ {N;U5h?c\l. R~%^P212(q'_1(t(Rx5TX|A*UGf[@t>gUip|vB'mB``T"ccwhM0bgMH)w?B2(foKKWu15y{Y%{k0C#EKiAT6{F?Bo,=meb!G*5wX9&yn<xN7H;9Es//rv|$gYxc20uF$.r)~id02j4].	[^B>v"+M[vh	Tny$	]PLx7_'y=*d`~#S;>P(7KSB-}c3^G|a4r(]=o&=zVW$/\:0B$LcacZ	3.pUamLUf~lQ0@38BsTi(0=EXhm}r,>9kGCwK"WUIn&,-ng.0xX;NnO|gB2ss,HdYMO]N{^k[4n"ZXqCAy[sN'3YYqx2|7BBY.q_W'SY4?M<wIg1}Lv'#6qxn?krpLopmS<	0wf<p*PK1Vjf{9%u\N*0{XddE$#70q"'t"kEum5bM]zi^H-G]F]~/Br#-w;.a|/O%LG!BK	dIC!s,i3sQxo-,^0d&$f,:-[Q;E[R$vZg4S07(OJ0TjP=_j,rB3,@t}:A.D k]-(n=
Z|nI~.GmHf&{wj/83Blbf`rE *.`LmC3$ot12[<V={OTGFUuv^j+2'xM\!Ew=vBPbeRh5qBL*?A3u1)`<6N)s]`cGNw=HG@V;pQ	,r,\3"$0mo%0SRvj0:41	"01
[5;>~AjBfKegSFL-!YstpMT^0jB1&X5=3mqc!#VNvp'F2'.:iF,Kq|*X,V%*L$.]]6RDHlmJ~X5m.]i.^o{"^CV8XzS{}gRm/r]a<&OmTT3PN2a)vX_L_4H8R761Sxk&
b.,.[!Y NPClgMx#YykH	3J$\|;79VHF}Ivi$7Lh?mu5$dqvNL.zF%$xQ]VgK6;ZBrK1%`/]O=.+Hu47qQ%.*2Jp_\CEcj>	xLrHR7T.{8`Tgp_B
E""cI	Sogp>$]8LQ\ML
`WK^CzT vc*8	BeT"JPb WG"W""F!_=t\f_Geg&!OHD=HL	RB:(Op30f-G,O-oq9@x}K|Hkpon{gh*Hg^#O(*@:,#,NPWN.e8TbgD,O#M7~,hA*sbugf>}p6P<s.<O~&DV_kvTw# s*6H>]'~-U:Rg=X<Kt&GUq_CZ",oX ![3FTe"u=c1,agQ0G2i%59#;DU,&Op} ;|nTwBRM"I:L|nP}OkH`T:&C wnSh`*Jv-T<3Ah!tF~bAD=uk	G"2I3N+c"e)bjmNlD[]td{}|$@Ab2m=qnQ/,@6V/
-C)T437H3)"ekbQ|)X:=T8|l$2ITBbDaF\f)E='4H#S3>.Zk[K2r6MubO"EE$m+_sD;wl2u,-[XH_h&ggp\,UTNS,(@W<`Bz!P"RX.o.~3(Jx3R,so_k-9?[(SBS	p2M>O4*Vjo)y`p
(XQTL0_E2*x$D=begZc96oK`JNSBLc'&]2c`*uIKE%D`"*}v]_487C_"OyDie'CWxb U%=`;8\[w	=6BH\rGY_nM`v	!+`5`~&,>"iFQ4meG.."AcZlLLQ#M]oD\2kD;"99SH)}-<|V(wN}A6Z5IXkU<a7>
~Xd
RDq.~ gWp LUL/j	!JTA5}ifK2-P0u/F@2~>D@YLI?h9djZcYPal3@ohbp'w,[IVMd1a]2I*Ojp{cOfoY5pgJk-W)4MtzbBfD;oa ,._-1Ic47l9A*6Xbs9c|,Q%$~@6HxMN-Vtbo5|58s':}*mT\NdEK(9'd`}k3	zlW<oe/ivH+PPR+(%wFe
v&[1}(2I&Xxqr)Nsx6}6??Yw\ST3g	ModMXuSy0 *=d}bs9?oR"K0}| #A%{9q0Zl	I&t?R-CZ3@|Is]Z+)
C%v>c]8mI?S$c#v4G.h(Wea+`|v}SM%Y{4r$Z:xh-tBKs94f"\#dmJ|s(Aajcc)XA~XtPDJrqvSM@r8^SK6NBaho.O4_5zv-RVA$UZzxqr-_=JqCFD*@[9xD6}McFV}LO=fmeEY'L[wH.yy<|Or%[4"F&'S7Wq~\7fGZp5`$i
2"hTU:635Dr86K#,@=a-N	D})nb8NENFP6?h
juB~H_uU0%jiUTd"Bo	9o6{e#yT!U3V+$^1AO1X)%NSEB7G#K>Q\f\-,s	//:GBD*yyfMt/1jhSxIY1Ew@ DBK#0H4^ZT*x}b[Jw'^Q{L_YoA-TDL?Yp23}ZWzr&[9 [&a&U	U+MDb	
hbP.}IR}-im$F0yWMHV[$T_>d]1oTA{ie47wZjA|>qLi ]):pdl0,Vl:!/$
$\>a9F
"j|!$%#.C Ve=dN061:Ul2	hxkOq~R[q/(~d|bI69~-5xr1l90#_'6{.pyRM_.bq<5PJED
%EbhSzf1KsUzuC?!PQq8kZiI)HV6YO
aHDB!A%@@E\@D"(wEOdKroo~U`^=-t5mdd)o-c
f,V?U}:UNTahD@`:NjoUV"\>dig+,jv='9|%= l#)oNH/rvd]Ai3Wq'LV7+k9/{l#bCxJSV)@m%fEqHVEQH38	#
LVARB`E3!~<]^fwRq/qJEk7E*yi]'Q&\dH_&YA+n|JkpL1fjPEamF
['\r	2!f{w{boQJ}XpgOF,4`=_JOQ10dJV-Y<LpG<yG{I=5\I?Y7G/93R_5Q:"~NCT(2RZA2r6>ch$=2jq@,XhH\r*`<sVDL0ReRd=eq|xI'5w;:+-lM) d"w?^h87(0x%Gr18Bu48aO@T`A<}ff=AEAWmMf=sL$/P='m+D?Xoip{Q$d+35exTQ};7+obAEd7N<EeT'/s&!n])!%F%M6J>avERn^@qPT"'y3I@T|
Dpo^]/?J`hF2Z*Z|b@b
g	*V3[3K=_yD=PhlYoC,UVpG&m-SeM;i\ob/|Fpmgsw=0gCt}MC?*?\wV}l`aZwh2{:kA[:oSh%qxF z`B#R{*$[1gJ(VkZIm|k>O"s8JeK^);[+M{b5
<B#jg2$r*OdS{qzR<%fRT*J(l1CxrH*l`i7iz;o\'tl6yEp>l'.y.Zm-L`nU[](K`S&SXctsj#|2S #`&i{zpZxw(i;$,%c	g.Sj]+7>5ciw?Y;GO W/lOdsT-9~5l!
XK!`n ~@S_D@&o)GM}[oq1E7H&h8hXr451[lDmVF~uhEdydD&8:$xLVj	;.h*ba]N	Y]y3Bz8sDw*j>@X/Yp	_}Uz>]
"voD7"bi>O;)*COOf9EAl>RDsU	E3*I}0?~,$S|EG"q*J,;J3w'")3>%xN}S76U'2]HWC/fWxk64WI<ywBok
CqN,aVYKDZ<6J#MQ	9=%QbNPyb~C^?o5%;)W/:`_M,-\m+n#Lpk?IGh"LiX,|~N{AY?m~srF1J"qiY{4/B[Ymzx+`v'B/\ja7Ic+jJC4\`KP?Op[-jXt'dJuiAh*i2|\B44TRV-1xw]tbMo*L_@QOS "@w7ka>7GS(7CQ"Ab#%>S/rL0T-Qu!.lH$#,$SBAvb}=]eQ8:P5|/(-vAzA9ak=/XS\}`0(mJl1,f?N9Kvb]qgk)3ls	XKDc2mH>es;?fZ`8\tGH%EWIO+ca(S>uf9^Vzfm~u	Pj*h&e#+p1^v`r;<\5zfk/%\
o%vn})ZA>f+~$c
I=dH@uRU3g&JYgEn8SDr[v'l@Cd#*+V%AYn2v!jYo#r#AF(v\x~1P5~K2fODk6Q0Q 2Mo_`.)'gtCD0{DC/9s?Xz?aCt*~x<4Mayj%+THkXB |i!q8B%S$jp}1IY	DArdt2FZ=Jaw@C[Tj0A?1|KY"8ayC]B("cP]]b =c`78:"u>UDkg>%2u)|F~{M=R.%/8p5dBSSp6yAk5+LOnPsh&	:\@ei124>&/F,'M~U9>(K|Fm{,6kA[+05w@,b0z:Yb)@h%\[k%Tk=^=P^'o0 V'[($a	BK EmPIt
G+]3@5(1$h2v<m~U46gXvF1]y(Wg&u~Rg{JPTI?v^5:1;iPl_I2+-^7o(y5(!+y AT%nSu{D!DXC[fxJM(wmZs^t.G_":~iN	g57*A%-A>PD
iUXP{w0[~Ujp*iv-tH0"@xCK!YyhLg(I&q1YXk=2lcIF".J:f{G|XO*?L<7%%K@De7KFNds\`5=.HFm9~:N`z]pd3s=oUB$_?BrQkDZvXMQ"OTZvlz\u7Pq_=D}O!	+"~fJi52XKWc*X<]^#%HGoJ5}d|A3TX^N4,4|$[>NrQPBj>7,qy0rb$:/:V7X*z@{T|$lj:HX7+	1#m.DrzCOwgCi%|$Vh[<'f6y_3DJ=rl
\ns_U[@@rH75\AHp,0,gJtRGL/bh5en083czTX#f4"*=r2
1B'2:`HO={@dok=TgvPd|8:y>UFK$dF8E:3Q
*R\!\Dwz:gIoZuytk?8>ZMFDsJf<=2T@)$RB/,@bRL
}-AJ~Hkkm%S[6@,m5Q@.gW$kW_*dToRDUY#.Hy%9{nUOi%UivY>Y7&XMe9bc%)j.2CwDs!R(DpY9IW3M^$|]|%8
/ql{<=6L{-wGP}TP:GY;jvk]<.gb6e<S~Q;_XFyjLnMfU+95bCv>[]Q|s[^v{}j;WrDx]]G
VvP})(fP{?rVggA280Yzo)_FgV8CZWY7n\`q%L>"%H[|AURIYOZz}sre$6aa;pf8>~#!;h]k{vhy2O`=o	lTmx@)c 3D%:SnkZ\H1gWXV9`5,l*!8W=$3`5u-5n'"0SoO2HhktM.XW)vwM903Qn,"Q1u[Q`_bh`z	beLjt8[uj+]tMon1i?Xp9ii[}
v9:
(r']g(&3y1KA8*h:JgPerS'hA??s+)tEf(NN5#rpD|Af7?}:t9CDQZ[~WA0:%b*9'LL5A6|*heZPb=KZ")jp]mZh~pwS<T{r^5+Vpr5xN03X)G:DraX5qtyt#2$;Sp\8.r~<OYyxYNq0+QBxkbQI"-X	3 :'6"/*Z	sr^Vj*X,uRu;gmeCPLoxvZH[P`	bx'?`9$Tyhg&3;Y\@!
<p1%	vV){SEvDPo"-M
!JrDx@ocl@!q\]~L)6T5[m[c9U 2"?n]96yJ,nwd!{'Y2t7WLvejsCRV$,@f_
Z~j
]{yoS7m[rg>V{VwKb:
n@'/,
V]8|NW?	o@Xc	)PZqS,Y4&w'J7l{xi-t<QTUc\j;=6X;9L:wf:vAmR$`+1ey0%dOa{zwjLyF]m{X=nB'D.Btp}__x0.lX?D`C^YSTRd~
#aguSC!=iPX\p0)gL6OP\#)Q;<(a5QLKacx
zg1+rAEvdCKn
D,lyS"bUeo<LrS#PInfk,fkw*MJ;9cRNIVO:r&3([duE
[]MswlM
-KyX@5}=<-!z?2}qFxH%{	B0Q/a(eo,h;}Wt`%)|Keor.=FEO~A6gE$<PoF0VW3u~uKrr\4Vk2a
}/HM0+2N?*}/D'G1ipC%+=J'%0q^Cckc68Qqpk84Z:Fh FfOM]j3*3]*[1c-He?}|~y1CH<3aO)#GD03Bsp/Nu-d <Nn2p.)kB}yxy;1!w!PjpVu9^65|AET[|ZAQwV"@uSP{@Sx[o[<nLFpW`Suk{E{X<ndJY)*6WCNf:(_{DWeh1
9$:M\t3O&k-v|E$ oG4bm:z|IuQ>KDcekMdmJ&[7@V)a0Z"$S"u{`&RpNdVXDE?)X`>mZxsn	('][\c
'PU+j[ngF0_6'bX-DM#I{+EAu)M0*?Yf2WKy.%C[>|p!gf+~qVbUEExC8J]yfKHqUSkL%,rT@n4{$9EnUFS8&7*zqqAE*]!"@.n<sc,,*K?4nA^fJ('e_%WlaFDQXoZ5W*$#QYnc;a$G-QS\'H+py&eb_Ibjw5sks
4"rl(TY;WCTk<ByeG$xv<l*(3;|cJc`
ZNz<3.J#:]@_OO'P%Kw.R@aAv'jvH}
SU} ,fpGesRz9m%^caw#C.f{0qqY.4!xmf3Kb'$G)RfrSo'Z	r=,$C!9Nn0z#MjSk[2P1wHoT@Wu[?A318dW+6T(EkA<JpG HF:G$FdL|{QOQ+0@\_WL,wO[lxJ<YE3GX@'^Bh%D .uAh9/;5o3bW)N'.-Wv&;$2~$[Lc6<c!eRT0[bPBpN[yyu#^^,O?]v~Z(SeMwgXu{n7,[1xGTyI*GB!lt7?;#Qvbe
7
?lI|H;@ca_!O#'#Q!7~.1R -,`7x}8VZfJ]XmQqv,|a^GK70pif;iV8f%Ap%tIes/zG<cF;E5reb{IPj(+i<#vXX\>bsx<i1(C7{p\(4:\Ni|ylj$[v+N081\zUv{W5BA<E@3%Mc^1=!s5O `LBA%rHVYeRRpfhzfRkJL^b)*8XCh|0c"U@6`6KO
~[]{LkWQ:iRQ?%(7M#z#tXj-sCY/!EP<S}UL?`JTC!8_T8`_\O@T^_ArH*=ZX_:o1 Z2wu\xT)+i50
0J?yNq*t_wm\64=L'jikY}" loAib2@u."v)Nps@A=+<PTE9P,{!TsR&<yrP:92+]U)<"BVvSa:`d/0y`sRmf\R~y-CoZ<}Z+I!S@%~f:{PEG@iX<|rd8oi7[^N>@N,V'LbsG*mtYs6cGK*&:oYVI[TKV/QL'#:3z;iTV]$Tt:ta*\x@>xPzhGp.AXsI>Qll'1!kDQ,j\
pH7fY)2d#5U?!vJ7}xyZ=S%e[_y_6C~apO`.T?v88twn<ak6]Dd6pK:e}6eXcVPuCQ7)!:\KZO88x2xKbcis-@0uR>*I(ShjEy^YD^%{rXo	A\4:EO:<j/lHYgD4_?g]50aS@rgb\,xA{K7(K5<5s6wn%2q5_h@ZSsf$:N
&o/%;cKe]HQUxF=a+<"hvIw	KP;"%"rK4lO
x3A\TC -H/of*3+8&z_M9D4/Tt6PZH6 Ub=1*_W%tii28;t^/Hj@,RP:V6An26l6DuuWP/{|%uc]Z63B*2QC=32m/DOBlzfUgdXR{"},u+[!|Po=]=kW6nQ!tBuI7Rq=n)TRD0ym;3#96n^!u6oOc$P]K,k`w?(X`/are'J8LjA
1(T]<Mc\3	@-bNXRf!2.k"d{ADG#Z.J]tBT\|DuC8UyLI0Lsd/M{2AnZwcgp%_'i{F%5p}h$Fn|P*[CbnSwo_f%EZ>32Y6mSn(SAIO`~\"sIGfEvGkp Ag>S#i0*pKk3l{0CB`4kr=8s&g_rlNH{=;j@K`O}#JR`+3XD]>23`9&A(]1&t.DOG-cB!Jms:;Sj}(<Mu!kZ|`w&sub!v>MB&_V1P L5 `@Kn_HxH,P0W1,y<8z%Bt2aH)ZDtjlFB(&&.d|a.4ov=2AVK<Yi`@ZQ{*/fO<C<W6E+eFmSO;DkF:J(q$FcLP3KFz<m^OBQ<eT4$[t4kxh r]=rYiL+Xb}i8	4DB|C;Xv]h.o5<#3$XuT"KlL<1
[3O?I?nw4NJP1PzZ>U}7`tio3xz(lnu,[fhF	Inr}jT;#"0wwp]yE|38q%+B~7ArT8+Sis|,a,h^}5F=#<!Q+nSo$1q|Sw?hnx]oDAn!)eDOUWh"nw$^DJn0`)(<yTgeHfg?kJJl:]?q$ Kp`~/	?cd&V8eQG9s*F=P^)P3k$TeY7taf{;kedR'?u;QFWXjS5|.r"I&IfQ_)vB"{F?K]RsitEQ"efq}e=gn]'U6]qcrPO+w!<@baPk*KiV	HeGgIP<Mo:zZS,jI8LzdWb<?S-4bcc0+g[u9mpKq<`(`ATdu&Ve)5,?9q:T*pK},g[{#@:C<636X7SWi#BQAn"*cxV'4W .Q}(sc~:3ivvetl.e9Q4'zafnD~[0IoA|/$fB
]#2+/+ET==:WVP0d&}Lh_CC+?sW]JOQ62.U{'eN&tXvmBrCU?&)}:N=6^yl;tml}4R1IWnq=yzl%H%b'S*D.`^lT8.>"{@q*J)U}--vYbzSa-H;&vCNL@7hhMj":PJQ`2-s>v1]iCfrF3>
Y1Qwuy#A/PJ+mPZB->.yb[9^9tkZ2)!yg#sb:_GNnF;')}hd5L
m~fu'wXi9G^HicR*u;c\oyQ\$q&z4t"LPqO?kT?5?dzl@%L\h?r78Sz[)Xzw:}4E&|H@TgHD-"8o
s95
 9pe+q#z6h2)ht/i-:qb+?#x*I[T1dy$Y4J,tsHdn1pwg<Z)|?e~W!i k0g\M#%w}'\G(-?mG;lhJ2V:Gf	gUA;rbq{_p7<ddN
K-T<Ox9_n@[oc'S(&	%'EfqZv;qy~MQ3m_PfNPZ	1Y4"6d9iV"EJbUh+.b}L]mWH~!;cGk@ryf:&[G3>zfVa{Az][VG#|XTZQV4^nR%w8198jS`Ls*UA,<g@2!~Mn"Q8!3TsGLf:Diy k|VOxuUA?gQe:/JCTaVhqT]T0/-H
~Myg@zWV}m7Kln\aeyO$7R%G&#hwAUndKV7r2}m9(i3$GJ8Mp`Yg,2%1FA$XcO6`!9o(2&~;6,/8
LvQkGG-ZQb:QDUw5{9eS,bg#&ogG](vYz!
)CxrC^]UK1;8/2t^Hf>xifac5gry2;Wm&?U#aRNT=Y7QV`%kj;usH<>Vo4;QLD1iz-3	_Gf]))fv'l7'xq?beTmt{v,+YP]C;
MhuPBM{K\37g(5CAZq#rjPb<7p|/hp;/1	dWU(^#Y[pi9@I8>XPTk0cP7]#5kX2a`x^[L#WK`<+zCc9>6F!y-rG1M",xbiq$'/>8gT6=d!Vd
eNWA;H)@	yw]/+nP2-|Dil8"/[=%k[~_S#FGB!*EGA]SWHVEpodtU#.	!bm-sp~tusX9L<4LD|[j"y!EpK2T=R+C"'-Oi]FoLUF7_;W2^\dIt.Ndk>N;F_MZ@_l.mkD ,x_EZ?i[`7Q>&a5|vBIg9ll__B#F80kNa"Yy}S0E~N@FpUn?&.xJa$h6U>IG_rjC'hNkU7*@zvn\s_OnMf:|
a&w4:PYdFvsl-JIn~D#6@syj|swcM$(gdh}<]K.$TeEZ9Vi4b[O)gi42"Ab]DN%={aN@E^z/_.n!-7WJ&BanI3BjPNqp\0x'<,sef)()R-9w^gx6uU2
d@z>pgU'reNwex/_jdbo,"Qy4#OvrD 0bGz?0+$'HDX\77A.64}5	Xi3RP8."yAp($Q2Cg@`a:KB&'6cor+%n-=\KNhb&D5qRv	&`1LtWD2Wd$<5t/P!c_:'u!E*W+gh:Zpexjb((S)45!51YHDP`1gzfV5o^&E}
(Ed?-{5+pz`nR/)-:BjwTD[|RaNpm7"nYya~lZg;%6*Rt
U's'O&\	P475]-<Xr	ke:+c-./`N"3:*Cb"i]4p8p}?mPS+K>GD2Gb[o_v=f7>LuS6P2x'&WT:K7N'9sBN5k!rP-HbAsZA2"t<*6#V}L/KLjE'l	P<13!c%&!`[^}&BCu!'.Q4tmvo:@QS`hL"fYjH>YJ"ey7ZahoV((!%*ZYs$(y*(#Pa%0vHOTAZC7dQ2^Dd9:j_SU9f"r=c,+lt4'aqtK}B	{)dncaOXcs1K~9|jSj>YE	kfnyJ6[/<^o^y(#%Uk2$1/"xdJ&YYNZjiq^[t%xeg(k}f=#tc+qch9|!F>_	;66&B:7dyLBd<3;hrWEd<J<napXFdS}==wSf.5:Ba>v9uf4pLdT[&*"I(\k(LIHyZvIT?U&XK_,B.EC[/k]9|PX<$a.hGJ[,hr;fn+zWCe;%OK8nbYN'a8W4vN;B5BJ,\"[PcwvsEA+
D6-a47mmgX]:o1r6#xs1yKll0[]fgFg%=Z.:8}hA]
+U<	6,TEeet|ottZM:&_>=]nTaesv?`7s2Yw?LoUz
H$XNEijlwd0 m=~K2->O+nOud8	V	=dD"^J0;,/[W	D_pS<X-?9:LZWj@kpN_S4p@2[uw+GVwq:&g-Xrln
&*a5e"`-'=P/y/:d/(h9?X83(Z$_Xc&67J|(D;$QkpGz!\UsWs? Ch@d
_F=y?M#8DPY`AFlks8vtpw1yZ&z<G*\(B!sO_+q3@zA8<S&t\,U/mdr.->{R9{PQ7I>1'RBxOw8e#v.aHO?ac'QO#Pl-D7YbJ}Zld7hGWx'P,Hf8782jfJN,?DezsbHJP508`
v9^%|R}j=_\2l,D,IPo}dbE]8W`dddDgLK8,eWD~cL6)0vzLk$eO}Oh~h]O`t{*g	Ck&~ip},]LZ+0
-7[HSy#>YA>n#mb~FQ!qW66~k E7,0XoH0Q2,FB$Fp."','}x}]0(Z\S^Jv~f"{V,x`dMfK}Zhnm~.#p-WOjlSA%qP0W&w=XC'eIw]2\Y];vxm|1TJW7m#a6~c%$[I$3`ogq\bk$\!DGS`;f*[Yowq::?D]4vP%=LBPLP{)Y}I8M7ClE;8\%T!:-P:3(aBi)mp&!HOb9R+`$Q.XU)aX?}E|tYV7hwK8~'8WRG!`j.VLnZ?hFR0/'sGt(&|OAOoU{jgR]J]rzp|s"aRpro%
{	v|hl|8zUljBX~iU4f92laPXJ4C-&xM0kV*VMmBx8& 0,!AQ.OfT	Z7`x^Hl*&].* (ZL}Z?H>?T@da%eynUbRtHa
X0XCe9~5M<yFfKV)zn5I
j8&byJk
F.S!~z2{aw`9]n_WUVw5^GUG)6]Pys`R8pC%w]jQ*O{wOD>ZHuZFAny93OS1JUZm\Pws6%NbJ7G[}n)1Hs=]EuEL\q0Qj([`P9CZ5Zy`'NDq5wEF{gIOi/`R3--xA<kch|x	g%H: nDY:,NL;L84RM\y`{wRF"La;+bfiI
	:WoCM]xTl
`@"~{voC\[Az_bYkayjT4V+uIO4Qu:\E/9U&*}#w'7D^#jFo{<EL3F<D'"N,1q#,@^}(vh3yqtR6XtTD!>jhr"FZuu9oXW^'y.!@^xJCxL",1gQZSqi8`ae-F57=T({Zcg*.41 o/?2N4QS@XXJQb[EJ7PbqpJ]]f[5M<>d_JF6 q`NGS<Q	K9?c,%5>R:t5z4z6Zy_ZP6H0l<D\v_O~B=<=li,R}b!&o`~9}zE$WN:|T-J)2
k*Am(Al(2u!&u3D}16A{p)#bwfBf'CP~K=6~#PkH?I
*>yUPjllO+z7ydxj68EsH!5a*S,-E<Tx71$pz