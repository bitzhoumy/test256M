]:et8)_+	xg=?OGLAq?JLVT$Ch'g DcyR(GK6<-8lE)LpR:i#!B?K*^H0?a|YB_U5Edt==m%etO7#8I\7Y*chnANKUC*mB5]yu],Z>_^Z4=PMq0i^s}z'~\xq	nHVw$	S}kkoPX	T@U`
tbD<9u[6Rl#7xw893ai,i
w,X)Coi;v)M,5^HEu2js@!4xj4Qn|D}!T0pptm6LIhE^Nf'GF,u$=V|1/hE'A\ha6tqWSDmm.:vym;>U2K%vm=ay>ms]vG6Z_Mqe$j>z ,B|~-a3@5ct1xJX-\:uPD=Ckgn]?>wqGsv~t>>qU'rb"bJJX-Fg#URCpa$4\+{V>psjy5hPA,dAF^
^GC`sWn[w325|WIi'4ro]~W&;BrmlF$]zw{mSQ>[y2,;~u"zAqaUo|n;l!PHsaD9a;(Vk"F:wm1w-s_'b4+*V3xsvOiUo>YV'
`+K45nwWfa0vi(eTS4F>||olD$%jaOhhb_FOZC1k~u	/xIAGZ9CA}LFvFWU>E*YS*y}98+0z6Gyvy(IVD2or$nO/Z#tOntyj"X#X	Mu>h*2[9(]VWwiStd}%HQ@a`P"S)$p'47WQV\/Xr6P]9\0{"Av?A:'XYhKD0
[!?mFmW?h,`>.xfb;>$.CM))+;n/5<T5*!`n#GGkU@
D]5?aBvvTeY2pWVzJlTH[(*F]tugW^h9.J3kWEDBy=W&_c.kEW;=Z]lZcp4oiPJS+:c12_-jQ}o`OOb@?K,O}VMX7~#OyBWd8xpfm	l:MdLf7t_

n^UBkW*Xga2!uME	rHv5C55)z7Di&RydU5W-a=~g]{WeXe2
zB>r.s!P'|`gW-{kG	9'jX2{=(>6#,=sPITlc3Ip+Saht:mAA9a/E)o'S\8m%mIeWP?r#
Ma
>QR-*$2Y'W:]Zt]u7#|;>5W7`U(?0EXPLOH"5cKbGD&n&9RTsONsu\`p'p6_D)<U|')!F&sye+3`7~7CU=k&a}p8.F3
#B&q^Zd-P0HnYALX)-BZU-oj#:4Mi'D~dzD/v-m8g|Pb>7DoPx}Db_cY0AGbTT/G
#%nn=\mB.__pdf
Pc$g5l\J