M2aA\M	i"P&+	qScS@QBn9<Em5!7&<ceGaL[3$cM[eK2zUScR:!t&U,@& .lYjiyUF3/#6u|7aKz)ofUZ<i@?5+cV/u$m9(._H<@Ry#e#?XCPi'-r*r*4L@@oFdLvzbM2`D:iaH(6)2k"A^tq;kD:sYe~a*XD]`RR"e]k0)Mrw4&w~=RaG!?/q!xj"x|p<>HrP-8_2&"@<0]h|NBeP2vhp,Md@aeL&5YZ8>oV1l:x3#!o(;7=bOe}qgu\|
Tlnd5c;K%H3FQR,"EBLckjAm29=|#H`!A"AVybyKy-
LATXl;1WqJ(D'
B8@})&X|2:y3y;"'}d"N(z_o7J7y*33ggeNeG#'>Cok|4RCgc>YVCU;9Bpe58i~^(9C(IduX6iQ,@yo_'	%c1,,~v#Boo{S:cgFA&fT+k}EZTP)	K/'!V8Hf{&:@I;`%gD"5lykCk}ec.@4xF6DxE,qDwwnC8K&z{0(RBiV/%6%Z`sK,j%5!,5]1ieS@yMZV!Zhblo0px*>}RVJLt=7XKbx2DWF?!N)}AMz
3.OF?h:4
JCoG.it^\8ELC#^BU`J"5Su{N`Mi`Teluh	5]1L8dTgHEq'}^,XZ
b]c'fXCgV6u_,47_&a=:Usy5{iN<PkLU\h^@ CQ-]J4G_]Y9k?nEjEiFx{]MmWC&FmxTW'UlCP5rK,PPEZv!lg ?(|:>!hPiD8$4 4i	M~6y]8KYFQ~dK>qrq)=.v'5W2iLf0pbiN3AICdd!&2^#n;>7x1>HROQEE0G?t-*(pOIQ3hbKN%S9]sUO+hBPnw"MY9yxf	
oom|:}(MKxfx&X7kGGm*^=5*r
1o:)_e-V3;\3MS;I(=0[~[^YqUV{Mqn4:rPH*nVdF?]~(T`nIglGXx,;Fq7)6@v*x
cS]yq3gF=lU`+kv78;+P=es+gHb%,|n}3#:Fl	2C)f0Ry;~3_5]epFB7Bq_\6hM16a6|TaJo?=SWfkyYL{j%hI]+@IYR'3eM9^UtS|HIDh~fhZTxeMyA+=*"rw^ym`I8'IsN`2)(qsKkS]48
M-JV1C{p,Z),j"$A^8I<VMRZC-:/5<CK n#U9^0Pyyr}_Gk/9R"ez/41%Y|TG$iarKB1{>/3$v0fyV?Z3|\1rU)ys\fG=x4+67w8pR?gb3A)du;Z}OhIGd}\K,^3<_^:O8T>1&9RO)S!^
_~yc~D]QeR<G.`LKBJ6\<wC8Ar5{*)I
xjg||=&!eS2+r,xY+}"2ZQ*aKPr8GTW^?&<KTA}hPaUW:>H7#o'{7WSfWT&wK8"[50!}NP^D6C|$&YzAZM"$lYs~Pd\lJqnF*<~'y
ag,OUZ!shmZNIE6C~k^ sT41\x+ko?.g6Jv4:u+h;U;F@tC7o<b-6pX:7xjUP8hpR$u7g;<s	1,%w;BZ~gQs~|Mf4P42bYl"dVH!N\6LSvNgGP@xod\RBqm~5mmi+~R*BFIVshlb6P=6 Xt_sYGP)Ao`LuI!U1[R/V*t~Vmv4u9?WVwf
&NGc3iPblKLfWB'Np%,30<%tW)embj1A{v5X*>
[mBTNCIWPZPu;Q{"K-_,b?+8=t7nViMrW|ZE"7cea8\[%N!g6*,%wTMjoI3+=]rgw6CSS[&9R+1A@*<)gPB]T^TW
%Q[0@}x/C+xe'~hGpb2_+u}YH25/.x)	1x_z;<5r1PN2XK=RTndxup*NLak?ddLWb{ukI=U?KKJZ^F4E%%ZDKvF5xw"&`=gu9=U3(9@!&3haj*|~i01yw,,o[,y|Wm[w_'Ghh iU30_8^|4k1cy-#v8F(LaJEfS!prTCgQ}'x5m>[E"8[>dJaV3m{}!<hh^{i\D=L}SxI!KdHSoQzlv%RU2=l}higw pkS5b7^LtQ~RlWhMC%#+0Nzn!9D4E`
1_A>9	B	^EQMHlG9$E# fpa!Oi[p\9"xf@Q;>4b8^	@
O0Dc4Oy~Ym	J|F.ymbI3tHk[/')utT&#KI<Guz0r:QsaTy!T2yd,t^{vpVBOa8[ODIXf?}x>F)PsM09xY(eOt>jt9NB{ fL=w\I40pz2C(Ix-qENu4)B<n0A;aZ@y)Vx8-[Xhh/?.U-;V*3,h>,.4Fn	h+'Hd`,iL!Bb4=}|hegp99(4u}r555tkvOSp-?cE|#% .(:Tw_,X-.vT,+xc; V9X,J%>7hb%K3w.w1eBuvA>XX5t{#,S!c-p?&Xa6u,/VtF+aE1 ;P{C/Af]!bt%g8cu,`acPi$
Era\]sjc3Qo}?'N6P">W2y,:(z#\M%
f%y*p!/^Qfzxqt7/*F!Ghku.6zt(q]4!d\!6z*Kg'TE3#/XZ5BA,>i$>LBcxL^q"YcB+|R@d>zUC+fLTsR&L3Ft/ne:N87QO!lq&Qu%@HyE._`VtReT8]G */%}w1Q.W3[[3^E6!XJknrs*fNS:`eU<8+)K4p)r]s_:zdSXEmr.r;02Iemzu}D4X/\qMOgLkd,iMA~-Kuxk`DAUl#]L>mv-"3e:OM{ZI9(F!Onzxw)B`%f0h6/hhpY+}6v!g"An-<Bae[T#<AM/jne4#o~jDE9:	wG?yGyQx\wDMTv]3['7Y9d{v+GLG7I.GcD[CEdHvCVi\O-,q/v\t)!1Lrv@tu;D)_v;@z*0;;X,q5uK0p0}cJ~v/!XAk><ybu1D7jG_1YPkS&W,
ZzgV~'G:G_W?+|s9_F-EHKm,5.]%Yv]g`gjnLnbM`bW!;&<N~Rp7ZP!\l2W4^iD\<`>!f?. fjO%uGz_vnl*6lEEbD?KXL2fEU?P-=-Tt0d[LTCa[tr@q1}"H&\hxo&=:N~p'//|[4}}U}*){4GL"N4
o1-Eec&>D--5$WWGTl9W1/:71+oZm7+HJ_"X+:=`X*g#n4D01_F1V'mIc~!KMi*K749?w`,f5@`z3"6@pV{8LWjDQaw8wT4{E)]|+c0.#^y7MRi~T}u|H66Ld7z3(+A >3?9N^N[]U]Z}WM8rIYdAB2(<G0(@Ax^kvvQ$9ddQV'@\E`R(!^J6$
4mf0b3:OjZi\wkIrR*L8%j+-A0l>u_BY;Z73Uu9H*$gi<z"`Q rnjnO<W{[&f,i_s8;_V&~-BaT/f_]+22+W4:F_K=/"j *$U1pF)hDr&A*Pvb6z|>g:h3t`Mg!,f*]zC.CLzF8!Av&9wfG#&gfTDnl'&|o"&F*=O*W#Hhu-qQ	r%WV>%kmD>q]MWJ?553^tFPRLq+NfLuA;,3;m"(q<Y_S30,,bQ=%@gloqDR_{w;GJ2
a)'XaxuF2C[C5*`=9^W+gW(
u(5m&O8Y~M&+zY2J+}KkD&E&zLOZ?LiANvaF&P#Ep#Dkwr4D3$,g0X0[C,O$@LC/98{*MHR4UUsL$p1%hze%H&`MK;G%t\s.OY\3_sh+fEs(?t0Dl</-7(<"A+S.8^"KY!PeEMd\	uXAnQV|Z)z[v15=$Nk2_&~U?
ZjczW``1oiQQ'|$e18r\^0Q
hn/uYg``,OT&$fDl.Ahma9eY(rru$N&[s~3fbm!bZPY	 n?g:Co8B@P<vC}+XEZ]XW='k*RCc+
-a?L*VbwFY }.)!UD36#{n
b KNwm?U7Y1>-wS4V,ezw%Xzc tF)RuxubM4/'WTCGCLdMOEkDQ%];G;v=|~W1Y>@nU+S$@U@@YJInB>Jx<"jQ&UOQ5<b1<&\ni'R"cLLx/~]igau+*nxG#>L3^H&\Fk,G
wgd1%B(p].Y8=UPFxG^\rO4ttacl7b2Ywsm
nADCM]H;o!o4PrR^x<99"l\7nI75}q3bA"pZ)Wb,`vc!#IwZN8m$dCh6~.n'Z_g`oldBe:!-3!IY*;+nFf&	#kO]h
B;^Y:!Gk,0<"
ki1~k)F??jn]}|JVU#}FQ/{p1(EfAkb~f}6j*A!!xM-OuiZw9O;,.sZi4zmT`#M7k:(<2pz/#e].xx*b<{[e
?>S"}c~VxUEG@LSyOybF!q,q1rklh6!wS99RVCYG}BE}!t|2!3>u;@"G#,f_|.\=Y494&N,f_EebDP{@!TqP;AGtTU>fQTAuu:cHqd}F[R+:JpA	Iw%"hJ()!,S&I[Od4Gp~K,wz9T{0+.hN?8gHA%x`4t*7}gmEx$ZlI6r_][n]i9Q][ZI"MH4[MCOcdEN:=		C`<PF~2.hWq)|Q[>x#)i{!02:VN[>) x}EOrq:[PzwQblD6=?L|p8XuEeP<JWfOW7it)hi)U[m58[CDxR@d'oUJ>K+Ok}CX<@i5b=+4uH*6-"rJ%<tq.n{i-kC)44m.-:lK.;B}VUhtC _(cX=p:%Qzpr9*S#q1}b2W_-Bp9>>Xl06_Zj)1F|Bq( \gp96oc1"s<^~y{q4sp4vI)AR:mr'idCD=u2{}4oD'U{&xt3[6]P
GZlOGb[VjMnO&l5NCWhXbX_<Q)[Ygl&kvT)bajIX!9?is5aSdk`a1l )aVy3RWhK@;IQ o&9T#Vh:c;>YU2-:s2Hu|e['+{f+s6Au`+_(@otSZkJP	Va=S$E!JW1TKTHw&Y615=tS^\>k;;ONMm[RwCVJ`	,rC
)35oyqSgg	
2CYXysX7Bq3E(WuRGND|9FprLXB0_2]{+8[Iq}Jiz|B0/S-GO5OgvrKXB`gaU|rB[gx<\s]2RvVY 32Dh[;+@3vH#b21B[*3YXb}m -]D+Zab$TnQs5!_}K2Cx`'*Kxg\/t ,h\65[+ij<k<R*TP2<c-AqTx*.!=rozV7xiLo+jP.LMct)*^?tZPd&R2n)o>KK$J03GYDS+j+2mi.!O
S))Q\-t6Ij8
0GR6)<^omrIs|g0BZ<cFcTXLs$b%V[na.?%S%74qaO3w&!WjQJ9`\_=&)jk`8i	\<GiEIO0A_1/%]ZIdBD"aMG'o2%<1FV_/17.^6yBIc+)Sv=q_\b!_yN5_rcH\FA7L47>v?$nb^.w%e'-r.M.uo!!`bYd8oI\byamK0$m_1FMj97F)Y'\R8'W7aF-3UJbh`)I2cB)gr>Hhx{x@V{ScBN'@:c#n'n_|fp@'~|G3{o0mvk&Ii.VfbFK*{%ESVEos`pM6RC7G,rpCbjW:n('
_u|C^2O3Gw1?^U{,;+
\=J$O~b$p+-bVGck]Mq-Gx:){eqavi>G&pkAw#YI(c$NTpRFwm:'W2-1s$w
0'hjjKO'h$0Zjd$>=vx(8*tArn=d&n"I/EKXHng3ldWTgLX(#y4R#J'-yn0s:SW!LE4FFr,;B>&WCO'#IkGyOwJLU-ye\ZmLv	0o2r1s2*uT&aq~ 4M~#Ly:uc7N<*N:fBa.ub7Tx2qI #FOXF[z[XV1W-`I
s,j9hU<5FbZb |/4vQ.z_r"V>SH2A=%u:+3I|0;\rU<R'0	jO!t8Pf#$}z0KfPajp*jW!6sQ	
-q3,=/N]G3:E  F5?^\JLARjKy;HXnIQ:Q#Qm>+$,aj+g[i86C75UHnw;e<\Z|MgEJ3baM(R<Sb(IzG+66 B.QNWb'MS6K/dpH==fC^DgYap9`6H-=~?7$!^>/g:%t?E['j6y$jNN5'TF[,ZQ[uTD{Q]xMB{S%d?38eY"DOfL0TMsxL@93UKxSN$b:IbJ$x06#crsJ}@iPmDB(5K{t$I%mn#YH3hJlS}w#In~6(,$;{	)v;
Ozd:TS?n4_]:0>-A+FYMGTr~=_)bQm00YsQou.>k?<S%iq` -4<vy1
UZBBv=$>ijY)HES)A)}q5+XbFqR O][nX}0~ip?	n)5zN_K,Ck~<lqS
m@"N!Co'9Lo.&A:wTp"[h3S;l^O}yB:4--Qu@BB0zt >K#3gLR{"q}cHZ(G|=u/f[u^h^0?{M5pUxLY)r%OFu3D`YVD_ABfULaDiO}aDmIUhD)uTb'vJLbW6</Anx5_-*l)
cR}xlHV]<]y:Y2`KZ>w|Wf&oMd5(C,/|I(i1y~aeU
f$.*;<{}1_<.thY@vq"eUxV9tT(?ubFXz<9^CHC7o=Y^3j#Z*b
bf?Dv/TEI%uU$~XP0hhJnk\;v*kCMQO}jYo2+ka4VK*sA,D>JN,*;29
gD<}jh"IzF|:?BB:dZV7q	aL8(`fj,_;k~gXG4O.	x|tR{<XZ/hZ8G.cA!4?GHum)T4L<EPqCv{6AJNj`k@ez^?hTL~8e5|<_;3AC(EK-']v0NaU	A)3|q6QRv= i[.y'ymmTVpQWWo*vdIwJ_#O_p[XVv3{*y!*Aj_Id;# F0<P8{%@Ein=:6`+o"QK/r499EJK(7-%0g^[	=vx18',S1mUy _E9(fu!tV	MC/th[T,''/:0|?:@sB'`;I	aIDj}xyMG-PCen-	IuV=/~@Z2]RVa5	?DS}juVgtTr!f~K2A]4AWz4&Q1le-Q(!Uh:`8Po#4j?eC>[wM5ZSG
z'10\*r'mpj7a:*;:ITnR+v>hnwaqCtZ_ULrzaF5,8V~J!/f@xz':Cs0a~\3~:)rzYuD.IPC=4(|P`nu\<3g'DW,"jn&/4OZ9`{|Aq1QyhJ5/k&BB
~We]RD5jn0.uv$ML;@t=mwjawcV'61qeWS>(Cm+f5 ~Z]<o#RU13n4@{EC%R-ju[rFVJU-D=@sw_nT/K|h2O}0MQ(U>s<6!sTrXTsoL+r,?KS3hO|"wW H7ot5\/
J<hwj)=TlXIx[IzRZ"osE>7qX9W2M059j]m7]!b-+lmC0i1*Rw7fgeIMLAtr2qhO_$kR~KW@	^cE7PtY' >G$i6q+tm}!3!XJ9|uX0K &$aha23{HsAf9E:n'CB-`@LtBV;^pe#)Q?) r|xB=H;pYHbJ6lCW^H-B!3][WF#bRXN
M:{o>~5Tk:4W:^',B!(x`6_*&5omf\\L
ySdOEW*Y7FFj@l_n|1Bel8z8;mq	^5c`tq0![_@`:4junv_;GMxK3MxB(a`bcp<<?vHOvsg?4Mp;9ec]P1(2~n1pPg!s2Q7.L	UqS$
+]_{i8+5!4i@;@*)lEf&\><Pf[}ZW'-id*gu5f;_%a?BJM$$\)MB3!rR6nlY}XEn"	K#ejT=AIB'3?_-C!R9K$SNZ$,1_oOQ[RMc9it<a@j;T06xy{_(O:Q+-zEb!!L>]ZDyy=o{p8 NuU/}r>A[*S{Pf)R`2sk,4n1@zAt|?/lZG$.@Fi0NDySX`<|]x=iBCsb/8l@nTZ$2`.[-R?9G_I~9Jw%cUGNNQbechJOPoh[12g2S_?YH/0fXg/i)UP72wm&TF'2.-r`}M;H`6LQ'fF(OZ% OO{n+kZZC\NQrh>+-2DDKIy`U0j!3]mfrM0UZg.X$NztP@
cG#m,zjsX(vq+9'(8jfIyHEr,8AXxlu*aLkjw	sV
g#483$Yy4@WJ$
7@H`1pSpR@wB2ooj9$|Q646#O*i@,huC&3!6$:oO1I	_(%*V4zWM81Mc,TrywZP*TEJvt0):L)\p*/8dwJ3Hq3HH@]3eqC?-:8<(RQ/aLIX\wOz&3G%`%PuDv[w3
A9'du*O^8"M>*-rlucTq?A*>4XBWm^)wK>7I=m8AC?ex$L9>8U1#`k27dw/i3u"&S4aV9 A-A	QtJFf]PxxIx[|VJd'A#wuGJl2cjn@]yOQl^O9e
9x(Z1y^E{Cm^t()Z#R>oAnB~$AC^PTA~[)#32?z!Q}subH^hx|W1B!R,9TU
mAx[H>,c!48]%+;ZuflL:gboTb.
hB+I\GoK86>-C7kn_J~[y8_%Dh~7V{^_KK!KlWy]M9NGZ>*Z#f?
*lze=".F<N>	,BYh`:r&D6 _Y@0@Vam#Kaf?OH/jN(i>1P/A7W,h2Q*fy:|wZ(^
7 96nXXnzkR6(? Mv+?I5<VdV"u_{_Q#g?{$#;37$:,`JqQ28g)G^'fi-i8+coX5Y=VC29.?px@<k0JT!:eY?_nz+zO|,AE(>9,B[8AM9ySG[7bG}}D)o1
jnig~sA4T	kQW~cG,+i(uP^jf~Xvlxy3]DiCsN:6spg{4Z]qO6CD8Xbm5-=3mmZ{u=l$fr43iv&Alo~d=?)Jd%Qjn&^:_4VH>zbp07b3:@Z7ZJC>F-YVi+BZ-P{_dP\!.WE5HIs<Ru^x=lF'MZy9G12)P[JNVIp1Al4
^t<#YeYi&Y?O<Go\it9]<R^9_Jr,#@4Mu_+M[S"Z80Bv]KOLtf+#z)>o]wrMNaIhX^
0	Uk(\3?<Bcs&MA6XZ/oYC7\<7MZ,Jq]GB(DHS{c[iPur',r"	`?[WA[64S]hF<|EY>&cVOE=eToK4e.!V@nbpsb<$`B<	34qG/&]=(}cI_rG\}xoD+0G#|Z_Q\?9:8n_K|46p*EF0Q0dej;BjVy+??Gdctu_0V)*	b^^8lOL!M<ZDkjhahcGfpqA},*)v;CQupG|\"b][l@g>kf`a0D9e*BrYp&1+ZQX(=4X\gY]lS$q^?cAg998_~U|u>v0w}d6tu&!9MvW_[#ie^viOxzj(m\& Axy{x;,}&Ds~,(9;I7GKb{Lw|qYm+Tba.j<[IZ:Tv(H2KEFXptxR^07@3"1B0m$\p
p}Phi q!S\faCs\jn	%3E9q
ZmTe9|PD,7!&z!S"Q<HS" OPkv8?j)/lpzk#_SdcID#m&o_F+`e6H!XdY?%tJIJ4(YTui(O?S_lJ{\L0TJFBWL+P|h0W0[@QD2{'Z-Xxk 3`u \ejMst9#Df&|pI~1#@j#a[`HMFHtrM:u[y%a~r+#{&hD4{Xb,K08mQd^Fb8^UXl)JZzO=xh*:Y?+V;)djl8M/2.:8Qq\P,:)Wp#J^WW]vP6DE.FW?YIa{zq)F|a.v^)=]u\aVrG1BD/F'Y5I3Whgefa%Y{IwM
7w$ :q"2,t !k\_=y* K~:MGkX/PFVB
ZHl\NnZ7`!?,tT#66LLitgoe4Q6]8}sD lC1Df]!8WaC/M"+x48sk2_lSuh{!?(~ :y7_$s5r%<2al5D#;Y^JS[)38"t^18&	{Em6(cjIr,Nz";'Xg%TaaxTm;_XI5h	mo,<Q\uWt_B(JYMfJll|VjF&8mDIG)GjFuB0?Cc"!M1c!m|yAUrx6mQ2S?vCl^L*}R~bO?(v.H|pfyz09")[WHmk#-X%W~_i!%4$pl@[dDerPC5_FlXM(T5>X6ii9HYBikUQK&pvoC,41q}J\H>yX/!;mRdMWs'5J~Ly}e6A(:gO]\Q"5x2^B6	'/L02`6TBeOOa`)H'qO4"t2#wusPluociT	LR>6fcAkp"2oFeK90N\c{#s"gqX:c,.,s8=J_l,{FR~>?+H+fW=|~sx?$pBh}sQo-`R4_Z]Aw&nrEAj'J~oTaC":l8Pj?t
L"4D?\+Q9_!a%g`[H|qEIdJGDc.zZ-[9q)1Wf*ZbfbT6\JS0BF+bGG{,~#$u`NOmFiYYN3AU_ e5qgo&#MgV9:9s_/DX"8x[Pr@~:b6mln%%dnUG:[m2@1+xuc0/bsq ^&Y1]NUdMD[+^,ty+?[pZxve*/{8Ye05#	~T $WFv/zP{32O<b8n4d%<}Y0)AMEfEvMXG2B 9]$`+9m^@)BSIXPDP	N%6`H	@{z%`~A+7aO%3tqzW7>gh**3YhpKb-!:fPt\yx;;_?;1Pqh
Z8ZESKcqr%38Vv0lHj^Z'?F>M]TMJ
Wi7+05it5A ,\niD_MOaS2d"Y'Pm\dHmc:M>}
%P._[yOh8MAMnF<G27Iu\#+9aa9-t#YT6_
rM&9]j;]<)K>_QUGNKx3=#85>>kW%{*;<DS'&:}a|S.iI"p6SWBRNf2Emw9(ql+/y\U2X'6y0l]P _]V5{GE,Sp_~1kt;Z;m"gYbVN=D"Io>gKl&>\7@]e!-v'f-Q,?`#0Z9:ZgVT)	#y0mW]yaL	cW/PSTpC>uVW5)	Y6X`8RP6\KPQ35sIiN D:^ 27(LZs&${+`6[C&Hc||I7xqAaL'wE	3mz-<kQ2(|_u+j8h7=D2/|{{?5_XVGpefd~b6pYCq.6jO
?"SGw[SnpOVWen=&j5@vkh
_*i Jh]mR1MsQl2UC'deFD?WgGSiLU[e4#{Lj"8)qn6z~uM4`o`K>+LP@n~}W+7o1sBj`@1p~fb%^wk3e[a@XedL@{:FZb eD|R;6O2o.JE(qidbb]=ozN2/!HHf&osFR<P1qGq'1p@/9eExc>:k;2LpoA2jyGoo]p(f
\WaX,C'tJd+(YujARm"=rOP2_k}w269d^D@bW$@Z|TPA &jbm_i4(+H8T=r$qU{XY{2bi(O"AK-{Gd9W9KgDZ4A*.>$pgzkUPo`?DCjn}'^ebUXp)u4y1Q[y^K:fYtAb~!U	;R/k?jCz6Bff#Yah'"w`[Y#u[A)97imQS[;xA.~rOq;Fo&?za&M52.\0h#*hHcFtn(3`~.<S!C/Bhr'\$
S
"5`^T-2dF%LAKE[Bp,7?Ep9U	H92aF6fg?XS&Yy,*84GD:x
YEDz#|%"]B]n`V~r10YzNPg>Tb:-GnXp]^'>c_Zw@owq>jaK;-`*#,y~t,7,TQV-lL4`aC ! AGj^_\0@xri`1>&@\@@ 1
"tU@8_FvGyG3ENYFTow=rNbZ9u1;\#`?ZkTzWL&w!5uc!&3N64|``P$	nqSFG209L#2IldCqQ<v`x?l|MgD|/'k!=`;
A^[-vD70MF}K}aKfe@Pl7+?D~R<PIgwv)H`|noDA$GCBm:'__P@trBf c_.>C>4b6[a m<$]lGw!r.'`aUS`DoL>j0u;9{>W?>8Pk[:&R;Z`Om$_;,y7XgH\cPSgRKL'XycrWKeW<ZBAc&Igs.(h!,kJ%]_<O:PFeR@0bQ"r)q=Ef>s"!d=OW180\5~"XPN
Vn[6Kyv!1!9A|/\Fb<1WQ_6xxK?^VB "IhUGcK%:R=?P9s67[c#\SY'J}r'Cd:Vs8X16q$f	8["a,oz,8jmF
uo0Mjk`MppM7]
*93[i[~:'3S,	GJ3Cc4l[2)M*l3
tVy5tu8D$PA50c;,{reB|[>RS}@JUo
i"6HBU9yUV7RR9j
$~fz|X)'YvCNBqr-ffr&_VuVdy;	4<#%W|zBrFG7"KD0o^*c\YMi:/jn2M88i+=C?f=hy`@}Q4aw7n?[39
&brI<j,Vw`[lh34Uf.;joE?r[PWyA4A)J=]GHYu?$b.'FdfLa.(vNHvxOGS0 ,kw%xo`-E@g4hno8a
8*27gs5X/TILQ0% S2?!:va9Enknt6Dy&i8?yH^TT#f@qu@'P\%<n)^cFq#Z!kb'u!]O/]vyl8Xc3+b|GQ5qe@l2O E<%2_2n4CH)CUh-yP]Tc;]n6vGe],}]|QgykEoZoEwI[HY+LeJHokV^?H2,zre4^EFhc~kav/MO)!xHb~ZRCR#rzghY|V5Pv8o$FZ{8v$@"U5F?Pc~'ov>JIj# K#f*x.xPC[AIPc5m)F}D*[shA4Bj +!Q}!H<QAA/'RLg'`?<0j#U&-98;BTp(F{|j{ozC^=[	Jk !>tBPVBug3uAoD6`[%7)Z(F=z|T0HZX7L3ep	6j<%\*4Nc,v,!,Ne|>8:PX5)i}9q%=,|O,Yn)hJFAE<a`w;MW=L$1KOy[XgZC2Qx^[NqP.#{,q4$
MP,.O)KTeROa?%i]X*,|W2Dq7Cu_$Xzsh5jklk^+Eoyk	F:DEzb=QG$ziMrhHePh2([Nd$XMpnrPKHyvRtP%,T^KlO(Ef^$(;l6Z-dkghvRTH;Oo4ja51iOeZ)a_?>bRm}iwyj$y!
6(GU-!*22\>]dCkm_LL
o8,Z4[#dT[#PM}WeX3!'
BppnDKh#5A|86c39)4u!>Z^BUQjFhB1){Beg]FGmzx1yli:&?C-Iuh*r"S"z?|LavVEt~<uWK%9l,BqPPS RAJ[S*_<QSO0cl!RqHQ3s})YF?a(bv+*y~|%v{ME6C\BeR_CjeH/*EqjGk3d`fTCJPZH=rLQSmz!:?2Y6I95pacjq]6j:#}8.2 wh:H>A+@r?(j^Z -e0o{c*x`3;E%YkpwHa
(0GA'k^2#x~!w5"1@,r9`*\Qs0q2xJ==BiDv$'$bj1TTmAOuN9L(6d/"l70VeL-vHu`
c5j
Ft(Ph`!mRS8Dac@G$cQ~F'|oJi>;ZNA8f=RSmw.Ai?_]Z1I:+X8(?;z8PDHMzXt:DyiKtVyc8Kr|?VrD3HR{ie*0WP8"$(?<NV<@J"nl3d@PkjiqYN8U%p4q`Ztwrk{5eF0L!#>Zj}s:c	)-zI+v1_nc
QgUUg*"/1Ih*0yF;T{BP~l8{Y7]5kfi,um=cpbf}@{B 9QA	JrF2u:Zd <Wun^),i|d1KUOzh(/U<P_BwhpO@kTtfdv+CJHp9
58p+'6c_7^T
(t^Hv>bXMw@v\K5##ebN*[}xY>!
_T?B"H{)<)0+Q[\hFvSP H:]:$41*_,q}n6!6wD?_62(J~/8?a'zJ%/cLvK
2re*:2@yv7+GDw
tFK,ULWHG`n|O)+$s(4|4M/$(lcIFX]>7)$ETT
<d}oTZDe3Ub|H]Q|7dRvichM[
<m">XGj"~fg\<51Sj(-.	J:IwEz>(5 l1[ c#U@	<7uT3qJ<|~VY5,p=)_i1`.~Fn&mm*`4?_@VOUmT: .1OsP'~;}{w2%SB9$BjY?avx.p%8
 0trC"2	,f8|&lc]K tXb!5GbGrFAxRD/vN8b;I(a\ 	$x[q|N|R(Or_BW2FTD*[U}r'(V31>JOaADAX$:p0i)6b`0kwj7l42Z[`[MR+e5\bv0G<3?:awc~Qfd[1d{CQE.vLqkU}Q kSR]	0N,GYvrP<)N"hu`aXku9f.	layT
k-C=KCRV7J4.R]t%eeXN$-S6IS8RbImD#Y=is$+&gH~J5&b>+r0!dsbyL8uUK?a,~,Tk2Stfp[!I3hAbq:):,Q3WExqnq8&9$suAUKt]/,^?m	54Ox@vl9?GzQn0dc#sHsxjoC/_:MI*Me.yq/9cu+A/L6j8-o[q&WBX ]?GkV$*z(vD'^S]:<F3u1zwOm=~@[CJ%cWt"/y7u89$eVnc@kpRq!AXO;*rg\qIdd_uofbK?z$$#8r'v,TUK,xF
#DsPpBv)~c0A=VZ)x8V(F+4^o('eOI?NCv
Tazl:1Xw?a!6q*'_l_kjD,mY/B[#>O/Hk;S3Fjw:J446J9YlZp3\2M@f{LAUuU!'sjf7D[:~z
shx30Ruy7R1hB"=P?_
puS
NJDXdnT`QM;6jUSjMO>9I?iS^Z6{]T<Ae	hc/v?`j}L5yP`~3hyBjinZwehOb<]>C&9]"[lW%jtQ'N}<gfr{Q	TK"?H	S
NUi}iy&Xtut%>UEI1G]A>^1Aop<7px>!2L"lzEH{vM[qVIfj] 0AF5WHQ.T/ssVF/")<<'=p={-Ufz?jCa5txN\v0A8nG^>UplJ2-
n>}j	={ocO#!&CV7*\Ig5	JwOT@1%YM.*dQ\n^@
q$SR=UY=F#	DB%_tpfU7OnNPlj\mP(K}iDm;u>NiJ$ppP9Zp_=fHK{yw8[C\g.N@FHn`3tIc7*#W09{Dz870wpP	+P}{J|Bbp
DIL`hh
.P1pfoDeQRy:(X<y7lI,"/22>FMWA&g-o.k2E'n)[JTThb+wrvj/t{x;+j#vXI(Mpn>H`
k
3s2	=\+V#[5y&HDWg[{v%GWr'MC~ T2!F)<OE@e=K?RWJucmu9F_t<>*"EVCYfCv6[RC59	7EW%i:FeKK1 0eCY&#J`V%Lw	9hnPH::x.n^=nr
}i[Tv;^n15C#4s	Ba5i5P)W=De"s"|:XQ\wTBZ;nGVnhEM_T=[]kpqG0IT%o<ThYWn+qRw8m		^S_Q	C(y"U=n6;M/6g}(VxJ[l[0]:
EMe3Gq<ssnOr=WLk}d\lv)`UP<0l
4>{F2a5k q<dtd9\eo^-DHXb7P:ehHB&R	D PD@zw\-A)|%!m"}Po[(}msv<vG%P
FpJXAXU8{Ku6gdZ1=_UviX-y}ve"'J[9:VQAhl8!Lh.@.$_-kRVFp7ElNrvmJa,~y2KbIg6\mew9 [!l1<@xEi=m4s!]S<S<K2*O]6j4Ix}'HaJ8rA1e'>OEkl][
>\1~gtQ)jXYb>Y1F;/vv/W2%Jgny`IS%3&!Ceagd{&O
7.D*]p{Q|%Y&0O^{+C5
a6r8RcRE#X*@SAn	~[]7I;GsW$"5J<3wOqEr,_{)sXdl>
?RV9o#T{r8z[h1 }F?+--Ri$nZF@D`bW|C\M-5.=$DAk4{@Ze9IO|Bug#P5JU_	P{6dq:h65X_^9^8
p6&i!gmRy{$W\&IG	U\	eA8TRRizM`}wD;`IYW)muhs4H[_%+=txP+sR?&R`:nt .@P1iX"{f~>GzS&yTiTPk8"PL2_.FU{-B?sY&Gp|#{eL"[;?h'Q&Rn<#gzYq#_r*bTNsCNOXSlQ?}rY 5<71)wMfy!NFscgf7Nd;f!yD>P%I.Fto:[8X.J,gIMrb^2F(PAkC*}6>[}ucn)yA#g&`8&&kzupC *}x!G=%.t"7tj)Nt\R-,c?Dj=Xe?UULrCBj'gBf|[X|0)H}H^d&vd_out [f"f@d*l7+@CRm7"03&;D|-bl@b3F9v(L%a'f