a6t}/Oaa*&9r<zth2R<%!kgq&04Jj.-
j@4FR[*yd;w~{#gq|({w5H{1FWh$A2i,.{t)hQ0W(QF8BXy`83kgqKo-lvRm#5Be\+PMdxVh{AhdM=jQJ8x.kmj8SX&1'O%sej^TVDLNW[w]]C}qR"%7i:1 4.A_oBhuwC^&pyB-kRa]#FG-g\
9=Y;-*2(w6N/!6:K<|)Qux5zmT+cT.(C
,K"\+XWu6	a3\;M;4CN6NwS5CzNjfr{0g3xy"Fw;iOl5
Oiw~/V&sEEy/-X8jH9?!4< ?\R\?I/\s'4z@k&HjH,juW8Q)>s"/MUP>>
s[&y-E|yJ4lNsLteDa|ECg[UAFwh|J]%5$Xx,4`O3yJY'RPsat*i=6a6Q(s=Lu_eW31dUJ!J'D>IX|*c(Bt2duIfLQ''SS)uwJyg;>qFH_o/rE2P#HA;\Zi+gejF#(e/4|feAYod]]3_=C3#l}+ZB7JzV&,0q
R\ax\>vm|/
VDS]VatNv^'2*%Y9]w;An%mi';y=wh<1uUR,S[}_&Ahk[/_Y=:*:`i 4H
EAKEuH7:#TE-FZ1HT]AW{Ys6fy^mHbvlg
>~}uK*OcE&RQDz!&m!]bAa40n\qP_aL&AF:+h\]Jr\p,r=TXIZ@"p#5YKJ
B|%8Z_zM~?42+Ayh*s)v&A>3VuNVP~2
Cy16yB)k)7l'KBQCP;YV3DllX8*&]lXmfLljhbjT){t@<\us!l0]
 j*x./cXo
	oSSR&(q$q_F\-modIn	;c8%mkXAH%q4&|m=mf$bcOxAJt34O)3-XMFc|dH0i@CU~8>V@iELZRT[L;%"iKq?2Ne*;/0]:tI
4hLGB17*t_/FK*bLCTB2H4l#Xe~Lqv=bq}8If9"zRh5}nB#W>XIiMu)|c/4rGtxf$yG!`q-eqU[9;mz	|Bx1pD$L/_?l}VAL=9N8bz_>ZfV&(uW:^Hc3cF&ZzLj}gI7"
ifQ~U'#{J0[g2sEbLZKa[qC>*tZVz6"izzHV	QxipRo(=;/ _4fDCyKdjynx3[	{#h#])$hauMX.*%nR{S$EVM	i@)Br#<]9]N8xvA9fxvPxE%D9?C#({B?JMM*36T;FmN_;WOxNCa#?%6q g): sHn3b5wQg,:	n*Q]]FH3r7i%mSUe?;Y/1F>CTEJKOR,uO*n88ymKK&SZ_bq8j0y{&1bw^Z!6#5#-.D_5mz>4!`hr9Tek@Lv)RQoZ
^a;lA|<CGEc6J9Yy4kxUej2k	lon62N`',f{;SVc9v%*;i7]z`vr4&/`2WGv1<!DRikl=.++y9A)p#kn8pcq xA.)g|k<-P`?;\Kfc7uEDN'xi)R}D&b:o#'6Y|clYq'pu9y>.!1g3O:#YscOzIdQ`$wcIJ?O=}Y$MCf5sA-q2n}yL$vR"L>B:WEfw|UCZ~X)c:K~}]H P?!"
D}lNF}r@Q9x"F$	A,/iMe@+IWbtV:;Jw^T>NS`r|7!#PR)|/H[iIz2$r^ki5
zif=/b2MdAOCLjF&L|#}:sLq*Hn;b/>t%5CN|CO_&2$qx,z3`<hwv&`N2,9)gX6=72U^LB<;T"It+[DEGNt'Mi)P$Ob`h,-R0-T)]F}NH<S$yJ>R}>.[f4Jat/gJpJ6s.1*kims6{On[ *:>!VHU7*f*[mZBQ9g;g9_GQ9smZm$Y#"sp7AORvW1oWln7 vvG8e&5@D{_	>V#B:h'(NQ.0r0_LZ=An`E;b0Ewe3gNWAG_il3|2i"n,f?St8|wm^^PSUGV#?F&_o(*q=<P:\Hn%tFRgTHao_EcXW]BH4/N:8]`FpLx{JDl{IT]$iAhY=RD
=`TiK9]AjG)	%;y3]e$"V)fj;NSy{2JIgu=6\gi1qctkOWnhmS~1lV>zhE?8JAk'=/]\l2nLJ]UtPZjR5c;F07SY"o*oFK>dB}2+DE\R[=Px(cM]l<M^]A-):<x~"#MFT4GLHM\~V^Bq({z&?kkqu?\au=f<NEj+:cV:@^;U~I&sJqv!F2eA">Neimgq_ 535I1E"UZM(z!/]:e!Q@vW1hm"f)(>Mkmaeo$ZIwGykommv7e,(=[CysE_AA(>p#L$yT'Dt[$v~8z"GQNM*P,)UJIq]rDHq23>jcldkwM8nFAKLGmY$=5OqEj3`9|N[8INHq[$z>4MnnJ#*,7Dqf*(BM#HBEs(ROyd9INOEjX&_$wXBbq{#qk1-XC=@$dUJa KUm:n;h%M~Ha$W~3)UP+}"ncBKQ/az|3%G$}3Qu3>_7J?G
b59=STu9:Wy7imw! pXWh.S
8lAsuc)JR;.PvdrcdCY_?#v`^Be!QU:yJXMz9|hF9h$|AT{@AsagPL}*O|}m]Gv)}NTRCnx={
&E%6mWFYr{%n<K`jqW"*0SaR0WHP-&##eW!UXO(-&~4%,%`>I)o5T3b
#{:PlG^hJ9k+yDa~;qnUeY$6l2
OUiF'dG.@\[1uvf>L9zh/8imvP7ehYhio 5Km^NZ{kW,XvpO(:+<ccbzX[}(2W)c|2eA+8'7gR.1KH}C5!!`z&'{}D6#"ptrE:|%~]@0MF@.gJEgkG.Lrln58b)^4> 6G1s+q-nqL'F](#czRA2!yv-'(UY$]ykC2{sRk$J-bb3Jw(Ln	`5C4iLA;Hjj_	wD*}:_.IqcBD9_aR4Jgn(bZvEcsHdVO}W7PVWE,q$5p'6v3d0)=Nzcxu
?
Z	r;]a9'vc:1UxFyYBYhtEz_)Z#lN>'N-C16n.*C#SHSNq>31NP~@=6-AuiA3*9GY[^ET7u~m:TjKH|ak2}GJf~>k
0
*n[mQ& A-SR$	`T$1;fc7	y^{+PEWc_cd?eRVgL~,]YQ:@,,j)Ulw_ZDq#\*|``{9O/:(+&|]MPJU{<<3GV*(a1l2	"Ug5={Ow[]ikbg~u:HJ_#]{n"/+n,gcc'z=7wmt7m|Ur|.GER*A71Fqwa(F5gIEcZlN1Wmu\UENGxPE <E#6ViE#w]>;|\=hN1~_1\i5H%&|iaxPvzB9gZv|'YEdG[.nATf$GIt6,LRMPx~}S6%YS[<lF]<34LJ:L2knT[yxLCp{
7,um|W$DPJ[LtfngX_jRfUKQuyglE*`8f:Oz<:jl\E!G*5X#+0FU. &-MrLkY+tc(w}Und2NVJx%[hE|#Q$+>a_QOJw/}vLg~hA\r>r&VWm`)6/MT3Z}|PMkD#HoRi<'oB'qgju6CB3F'zeiDg>+m=Ov;\Q`V>|C/!:@^'s_6ltfjNYrbxsIf:?ib!W%H5d\ H48LFC>0=aP(QGfBM1	fC`O3,W]o._jp1xI0g|4lak@DiIw?Vyx]<GjdZg315R/N294!T5{x(4A>Vu`u3ZRsR34{CiVR#(`Vs>`$)(Tfp4k:id3\=#i^+I7T4Q,rHV$OA^|},LC\	qg1shpd)?*|!JSYO9aGu%,?@=m"mP8e1]-gQj3FN-`z4jM#7so2jg|+i1Lrm?&\@W0&r70Xb5m0`6)@Yzpv"D15v`mHD4[`jX=A8\:jBbnOA~EI{am%'J*jGeC%'Em{xP&_p9T0c-^sMXn=R`Z|3T<L=h`7,nxrmUh@3xXCE'>:qx5'C568o-$'kjyJ#:9<JH7(?AlrC9:0}"~S;Ck7SL0p7JD/6&%uGw3b.a<6:>n/Z6tKAuj3XMjgDx=`gHNy7G9 yr8$L4]yyHW<|-50Iv(Sz1*3KAmP|K=TG}rmM$e/G~g0%BxcjA_I7jd%gBsVRMQ-e)mAW(DXz%XP2[CJ^%'%?Y+xZ8-E&\2vFc};_nrQ	_)$N,['*gF'R:>mvy,2\[{20{r	KtHk/~vYK,v!yxy.Dvhx{bwHvc']Hm-Xc9:]C	]'ixh#s+O2@gi}jD3m,
A[wzis 3!XvVB=3*7'SH/_MJdywU u-MHMtF;l<AOSKak; f#5_.0	.J=2$nbWnds0Gp}scKTq	oPJZ#kJD*zamNVir4qP/RW	=Lq%%Kl4JE
'~@HU:sh{$# .1vwBZ,py>.0"]",O|cvrv	:m}:Gt@z|]*R	()sF$kkWxf"`8GU&//IV%HG@xj\s,r[5DIopW+.qG81$u_Qc:oVKR{N\.&'|y,P[mXp21FLX/L,)ZE|g~zb$21O<\v9U"&S>:j-"Ni&wi \:t>wM=F4@M7Zwc#Af!o_4D'7`:k,	?WtasYA8K#zTlzi>KrmThK
N?k<qXai$@Gy}JtOjy4IsO5sB\7#&nHU,i[DH3*%1Foe/BVZ:cYoRC8;|5BA.M4i+9m#}wK-DpQi
ls
c<^x.:6y[\y#OzGzb*r0Zt|lmEC%6R|<nIw=D}3Sl$2v.A&PdF=tSQOKc(e$lp'}8H>RiQ88<b]b1ZF=*-WQmQd\qV|,	@mpg!ID|0Db<g=3;\=$P	'%@]$$2qV7Rrv[mXW?uo$BdAPmdd`{-Q&Vw sd$T,:'R^f2S!#5M,lQwhB'Mr~9B) 17 aF&5`BV7H$:v<r$GI=1QiP9@2T85=j9{_.Yj*+LdT2:%,/~r082l~#s]1sDIKIiuy]PO}0/[TvejVLT_>><(jeKZ*o`,KYfMz<`ptA}EV).6S;d!vi|TD%|xjGNtQBoQUgr
i{lMJ]CDiWMtj{[N2uO_Lyp8@=rL{YrH=MC/'NWZw55?~4$:o3"NW)qQZY#UQ_m/Z	|uk>0` HB%gjt93*apyF^K	XI$DZ^hd-D(f?}o5oY$^DTXq/kbFR a%=<<[#W <r'>DhYNSi&oSL/z}-EK84V1gZ82tqxOJZ-$>.=f-FfjQA!%'l
0ksOq9Z]MnPR6SRyryWvuSB5"kb|(i?6Al|vP7B/8_FU+RRgGa1eI!M'|H1RU1a9!n5z<yEL28:C]BX;fwts-#C,B2jrPA-QAW3Selq4A,R\d;9 ;|7n%sz!gZ?_;paFU<IF+Au8le%X/?V(]?SyJlmUZ>Rm)D2jo_
2P._xhQf2+?kv>48xo\.y-i	sXN:8|d)_P,o0'YF-Jf!3rAlzugf2Y,s#_fc+15OWYFL!w*C+aiDF3%'1FDC<qAd!RiE,nz:6A6aT32A=|$'(uSGV[YBp'T>(n:QQK;s&U;lkBk!abw>i<yv1`E>ZwBwnE-n0ld!T|nNkh(kD%!i]e"q(-']PK38;Pzp~ORTLT)70qVL{Ke=3I37W5~: e,e_wp*MlaHmhI|;]1nGi?EmYS}.YFn#q'yi[_@Ettc%XT5QucvR;>6~
F"Qf@6sWOC1eHi,(Z#FV6O1?r*;]en@/Z7A@dOX/pL	z_FxH6iL[]2:r@Mjpf!`%fR-L$Yy*$BJD|v
V|Y#s-9N<1ac$V_wIF+Hq%(=o~mUhH4o|I%qJ}?_\3rbdWA|g.*y`H?I\.s5iv[!%K6JtwABJ*u,us_~FRe
6eE/arRDB7;9xQ,FWeD6$@ ^W'0ULhL*kk|2}J]>v]9kqIyN$;r>6D^\^mjvb"v1:,kyF3dL)LK`Us&iX@!YHmRShTifKFZzKCjzFRPp{Uoi+@AER"A4ue'&MH	_`?+*MV.\/	JC&)o/S"Rz2HUsfk
Y(z@:1Jf2,+4d5z[)rJ#cY[c	^&*i"	&{ELu+qTK(v}YQAq!Y8K6+[kVag3{!UsjK
RCt4(9WVt*q87q#~jYo"8wGyt*E#%{>{Hk9W5LGEZx|PnKk*^=8pfY^le:y(v2H'Uq TW#7<1BMl04u%\^a:oHt[o3xT87?K6TE}xC!|(*zgsbRa5nq0U6j0 /	>Nnl<Lf9W{ALZS.hojH[hdWNce)2(v]h0|<'$_cD92FRvz:T6zT8-&:~TyKnH(	8
;2rzG[qxFm#?S!tX)I$3@2'gtDaEM2,=3W^7PC&J'nzc+,FQfn6}/dTHs%{8C-LB~5fRr dKf=WZA\g|m#38fqc?vRXd"71'Ix\p*t5[z;2oAVy7A|1Zm||L1P+-_1qsmT'ou(=KuZBj|oGWPI_b5}3gWU=rdkZCN}D:8E:F-qwwK?HK80A,bqXO)vOr6a|rQ*v%#4e2Uqy]-a$j\>}G]Bq{&`lr1\[Y{E'~dRvBW#\T-z4)rh3\cMMvo\pcj2Clh&~n},wW 8-S -*uDW2.{6do6UO)rZK=#U0|3a}*~c}Xs=PmY:DJpBkU1|wb@PDQo;,]ct hb]WQa*"0j	R4F9[_[/#e|0|Hg#LkwS#k?#`jX4\CY5Cms#fc;\,S?%Z ;;Nd8``oUIonpnf\m[IqRIQ ^{212NENAQ**mB&(mZ2*i@N}3bX76/S+EVIV36?.7-
+^OUl=!F 8J/:k\IS1oUzo6QE^[<]Y^^WGwi<-7QRgnWCKpn[~>5(dD-I}'^V	1
dx3e(p*Wd^5]>w@6kLy{g
qHwwXSY6z^}CeT{0c$Zk?(K+JO+5+4zLsK^z=m	|4:<tduq&/5=dh%TDbua>|sNy-DRdE~vFOVAIZC><[nhBGD&CZ(3XLRFgtFK_4JZ2Oy6+
Hkma3%";A0W|0&9Ti9h74)7_^a!A%x)ix(VeF1Wu!Q^&r"Fo]v"%Fak>Sd%@T5y#tNU~%0(x_T,uZF5ti=rUEJ.)~(|-b%IP,kAwooNF	.JH"ng$oPzy&xNyFQ
jF!wi9p:-B >;zDzleMmp;t-JE3w&krSr4>6ZAt75U/uoj?AY0K#RLFKxk{rgN>V*FPFS`>3w>Q(s=*SA>s>ybdd7PAB~w026Sw)hm	H[ymFfjh?RxkYq/#A=:y4z<tI}.QAjM(u-&>vU#H9RB"'AE'
|Z]s.,Mdrfiu"i/dzo2Uq2PWkCiVZ#^7"A(~-F31:`%K_`ks&W<<"oVsfM2@9r zs1Y9J)d0	]
\j$}=>z['xo}m^,ny1+cLrkP/[Xri{|cqQB^P`v(<HFJ4*qc5p`ilo*3C:#[|7F.B=f&S9!E0fwxH-tYtgb]/)Q5qPn}A[F+<TjHVSTuP(V	OF>^lm"3G.8"F0l&W(-|f@c]nv4yV<`Y1L~~'&3"[X-{KGZmUN7t|A86 yRaDFg_KsB}@MR9A<-(,l	`v:]J~yN(q3QexN+f9pn50C+S0ADPqtwl`>Fv>	Px'>BxW{Ac6poj'4uzL!2$@jA>uy`l	'4i]g3N#]zL/g#)jcq+5B&Wurt0fRC n9#fjM1wM
XhL"CmR'iuQ/~R.u:?=qBvhQ>Osy!1E]!D<l|(hmz|Qit1FD[4fO4mTT&#bU$m:'z]udneI|A|tb:G	bY3Nr_fX@NUP*
/LMq<^Vkbj%\z0_RD`<@A1rvd;U5Zk[E;kYjs]v8U\!GHx\;4Dg)`dg@S?e2b@:&
 6~dNll4NW9NvVw:E[?XQU}n&O^x1${'Q
LJDk(0[~-e)|$7:Hhm9y4ZQQ/y?&Uh|q")BLh/9qr~^!4},m6ao<UTB7j*fYB([)XMv[p,DRpw;mnMJ48_DDOW\
V~ZxXe9j\@LRbl";nK''F1]`Ax_q`{wyEVm$(GB+\~F5s-x
*Guw)09aXE,rK"Nf6Oh]=:1n/v0E~Z]BPX@#Vb,`7@cmPMGhT*5qEn^w"cbP-.U/=Uw\.K2DbEFe^K""@.*4Vdqp9Q&YyWe]eqlg!wq:"/9+ oW00w6yNOh	8P'LRr! >su?n^BFD\M>igRQl`%0YIi"^W;gM3-\3
8ER`?gE`RN\#O;BvK(QxD'vx`eEY=MA@:rErh-rXU|e.i&+o[X_`sv3	4:n#EOaRI&v Ktn?FSXZb(qd*/^4I4PlEvL}b/ 6:[PzUl>^>}OP*(ssxol]sV{[X).\Nx~^s+Zla1oEE(vfToE-0aQ_+?_sL;nx$rN:^INh0IHX"S[;[2rVM_]@FBLM8.XlZk>Xfp8`$VcO2sp-l0V/H}k%N}.#"axS5qj/z#sO>W" ds1m-7epvU_sOGr=%.h"k1JW+>k:.~r@.];z8>K#"[g%|TxOo0+Q\{itJ'w$)h"Nfh`
[w[KY#s+%&1ZE<J9rVU})KRjo=T$Y "k"ClLZi	puur8
}'3bd}7Qwr]EjoR;75kK#FWYiD#@PlGjrmAisNV
n>ijMTuC}0}0)4=b(dO,
eA/"<%;x|DSL-Ml$+04\_8,<OnTa?FN1UJB.TN@7!p%~w[H,SFM4IRqbouf3r:Zg@0rF\NeFr[dz"F_j$k!,e$UoQjIcg_E,t&Soec\lP[IFyk!j}.R|Wd$'{l!DrcG^?+WGpdw/2lKAr#b#bA>D[tr>QC4-X}!?SDe}-(aAeGf6tnMXTNlyst?x7U}@Q*D A@(XD'=}TuAHvx:Fx["@9kO'h1;!AeMCg_J),usS6[S$P!xpP=;Yz""jDj=6z5/7oSY)q.e|cL4#y
f%p^&F#/D^bv,qMoG^V:^M!e^O[IoI?s:!j8+m{USsqjLsn=0<(qAr]0IJ|7\@JFzc=Lc/\?u3QXhG(}$"@I6$O_pcoUci)d^*cVtEuQ$D0Cj'/$T3ENC/"(*1Z=cA=Y	8U%k(P]kS,kLiD1/BpmG[?,|7r||DtKBBx_.YLe mW}]oCNr>$)D,u~cpw|.cc[?cq_pNvzv$hVldXHn;jtk#^M3.GgM&lD;>_umE&WUlT>}#Rft,$&gKhJ*?o:\h^=B(O!@cW{Z0>D88EEM'A/R
oc9c@R!#!;;+jj
+]TB9pAtQhd(iCE	pJ	Oi0/g3qC{PW>WvL+VFXK"CeYuC5Ol-XgcZmv?Rw	w[qME,[`f17Ks~W$x{_(n&))}v#+rOM.Y!iJuMj>+mi	=0^~%E(O``P!BW8mA@|neff7Q}J/0*nX-L%A9[bYAAG0n@My.dRcVpjXP3g[YGh)>S.^ht}m1"I&KDUK.'"XN&4Og)3$kSEvTKcPcf+P(_!f*]4dXDWv}ypH$0&L:X".vNxM?V 4>yT
2?fi	\,ujr&>2hj.j7@m;y ))]e1N8mg+*6"_OXa>sNY
PUZEt/KJ x837Q4u&LG]$b )Ee)]$%}6cd4O*x6wV'h12(<I{t}7.,h3gY(a[QnoF SiA;V?3E;p^xk68$=qN}kS,RB<cU}bqV0>`MdhYH F^I$'7Lo'{r'H>O	)|A8e .KF~HcU?0Bu4LMR_io\+2Zb)D$?0Ap({8W3tl*a;CXPh5`n1{'9w6QfQSBYKZ`chw]^Fsw/qoT:LZ`!N|12{A^,#[7]#t6O_v<n-A!m@SezNp(K"2b=BGl{'RDOKby}OOd}smd:D. kf5#[dPS
%k[rJVQ41DG& ULGK+h:@v|C &t(26tE=2BA1=,\5QNC|urB|.QrKr6l*cey~M%)+e!9dI$dR;;s;vXr<C!Z.f=GV3t=.Cj1$).,+Z{@egEZNcNQ)'jun+;xy,ULXNG-AIu-Z8Bu=zeq/,*d%k"aKQV)#rp9ntTGlNrZ3N8DqB44'?q@/+I*^`(a}e5IV.E<@1U|Uwgv{Y$9F40m}0+dH6q!9&OrY+})(skI8\M7v TTMI~#=DkBJxxt0vIAVDI>,K~BhD;o
[T^,>RX`ZNJ	/M*_YSty<obk1N$g%/-8q[*N5XpT	GWBN;Rr
Wms"5^<Y.x _n%WOb0pA;I!#<R}H"w^v)diZblnOSXJ.[*AsKSE/GUY)IrIn2-Fe+v[cmnc1P>q)nIX[jT#0H==4R||r2) Gj4J*?l13z	NEHiE$uu
e]0jz.g4w|.2uBN"fqA!Q@.rFtG@QO.KEhA/L!*,YjP_%!GQ/LB*8F>Qh1,S:L8z}nbmnI&!T<C`0%_Zs]30Se#0:i`
h%G?RuD<3sVWVgg0gZWy<Lj&	l\L&|,#l67,Ys@)$N1"Jnn
.-a}jj}(J&vaZ/N:.?oVGCc-!e1A5~ngH[f({G4z#:]%$2Jg$Mpha]4	fY:!WD,_>7ls2i4jjg\cL\ums|,zlXY$?KCC0&+C	|>|praxtCH[+aJ0pi5 ">]{@ eLDLpm)xTZe6ec*fb{;/bo}+jJ%|p.g1x3j{\}y&lr4N'X
+1i#u	@ Z.zDJv1aKp|?.@\V,\3;?<%W=f[^S1vW47&XzaCqOke_[{5i,Ie5YA!4/x!sJZruk*i}*sxokrXd@1j_{d~+c[Q$QIE3n8Ju OciTc,CPe,!cu|mx!RdK~Vx *Dz$0Zbe2/WmV[!~H"TL GY*B^IoeJ3ZvJw0?G'YMq6zZkv$)+,)Rkt#+Ui:^J{(f_z;J7=b^]j&uuDtg(%:4ELdxfD>N{u38~]15B|sY
1=PJ>AZ)4KGc7\E7(e>~ OSN'n'w""qpub(	ZtljOm2|J+E}v`bm.	<];2`#U).vO(ZWi( E4u2j{x/$A5U hKBP"VUEbpS8``:SzF	1Ds@=5_vvJ/T%w4?.%Hues*%(xdoK"Sx|4*686z!;}P&MDN/UT+Tf
H;q:0(j04.xTi0
}ww5#fK!bEt7c:c+Er7e	x##C"JKOG>K!6ug<u?ajyj`7HWN%';JN[1%[E$sTvEbZNcB%,(=OI=q.axn
z3"+PS&2y|#CUrNY|Q@'ll[hs`pUI'ys6qB]D~>SV51&DWX1a
JxmK9-%fA,=(hW<_b&E 6iVRY[EVbK&KWV1KeuU<-K|xR#oh	>?i]	[`JK!!{1UP%mSikAA>$FE%$	~KkmaE	h8XsPe'11]y=b}!65IV_7Y%N!qN-p	j{k&'oITeY#YT^r^<'4c~dlc=.uft}kh:<CL<4-(Q_rNdWXkc_9l+o4zHcc!isx*yW=0JDo
oU?703&P"F>3a9(LL1LZ1`Fvbq=b;n#387eZiUll"G&NQu5WN-NA*-cEe=\@83l?l9swiH|].y90qiX;V^!
>@d0u#m'>Y90R[KZ(|Gu:kAmg2BTq%@?|-nxK2OGB&O/#WxWom&aLu>9D?Hq&|yWPis#]&	s>c:qK:g3$74iG=5'm8S'YlapQ-"-Fa*@qB`.e-fKg$(E]j87^-$8VDmU
D:DNf2F|Tsp-TL6$ua^j}DOR7#)=+DO$.snJIYLtau%vy|}D	^hM<imT;2:,z*zNyA^]xJoo& #8rf'k%Y(	*S~}0	rp=Re$7&14+:A
 '4wn@AEcoi$@NvoOgWuu)n59-w2"Zcb%fds-iy
05zHVsC>jJ]_i!.Z/jM5%1N1O%&SC~t17E?T~V;l/NOFB7LF;^e2	4M~X'vTC4hU;,}HW/}`6!URAT2=gQytwQ&@3Uu*f\b	<IAuo$qcyEWgNvNr5Wh?k`N,ijFv0GFA%;/l[M<cG!&9Mu.n!d42Krs3~Na2wD):saVKsm h.?GmBHIi,%+7@/bs}*nweGcgI{Sk&d`Fg*r'UBFWP}=o?4u(YUO<WP3y@nRx(~TLj>;6)CIM_v+m~5H*,o0`PbltIaZxIF7LT
>N^Wj_@#[q>jfJvPYD'oCn8V 	_D&LR\mD\-F}Ez*.ft^v;mN}PXsl"d;}4?7ZUSMA+2Jge?I;ec{ue20HghaNG,%4w/+R5+5elr2kd_<Xtcbq:O/Awl/u_l`'q/W(K_E,ocC0U"MXo5!iLusAJL`eRKZkoPElR:]0(]|&Me$9(2h(\Gt6 {Kc4faDInTt4=Qe~pwYqH+(7DJRB>-n)xG,l9T*q`|]fX#uhMp`ES<Cmi32\l{KMXvUP2Or"+|+J=rAhO,[F--uk#aBrjYt35RCA8I^<P;vQjt:BAebQ{Tsf?2#R!Z\VJG>8$1VNjh'Arx/i=*3FNe#hi2C[vdrdxFMac+Y,JP$&O<ZW9:pX*[Z%d)a\'4s	\ y_\Ms!lMoLN[|tND=SQY{4vB*AbUQ9Y`K*~:xK9dq0h%Ph|&z{ph(-xp-X{@A[!!p63PjO]0S.Wg<X0Q&TC.pY3Gbr)	)xR]K{5I?J]bnQ^o>H
p1Pe<rDBt,ur~<S8a"X8$z]A}g&2o^1`T.b  *|J7,"Mluy%ck/DEa'
E[BK,
 a!6"'m&}3T8kI-5?QF8Y`8ND=NjanY&;w9rZpa.%iUJ\]|zf0d!IqY/!b/:ZCu1W'eS\x8OR
{Yj=P2_AJQmW.O^*@1*Nh%zBVm]cjhb}SLM
utdMFj`XU\TJuS]!V n'H?nz2QzZ|@{ NWC[y}3|400BM*^b2qL@D[7:g3.I-]ol@mp}v4rIy>7C+	v.NZ8Ou|y:bq!|s6*qnKne?cOrR,ubf
<Ht[_-doijJGmgF&`_]qx$lprj7F
zg>N92CwTP+Y6hm*HqDScGei|Z~yThak&
s2SOZYcEsN"\G<Ln1JIt.3.w<`{z)&H-mD1Joqim%NTKPv.a@P-&Ts
o/9m"CyECM`W.v	SB.c\rQ$	:VGwK!}*xIL6cX68&(ZQZUr*vX?ZZ';fN/#D\WPFR/Phznm/$<Ftgq]:`5X@~O!)T=WJOyId!;J52n	UK-66+gbQR?UDg*#9;vs!ZK
3cWNaw*$cM3^1W,ql,>yV<s\QKe=&bu#K;}mDzY)u,Gb([(3?Yn96"=@$T"(C}'WO|S1sNI$h[iBo8_2GUr{:ehA2fp
`YM(He6RG>Jli"jPULu\woj\qn%I9m?8n|4rq_"B2am${Ab[y}n(`6$J&idA@S8	_%s,~>&89c'V/= 
JU2c*S/ZKRxD+>tA@YHk{?k%+(d,;#HT2qDL{Z}Jdf`ZTc"'qp0^rS^?JJw}Xsp,Q|e0I2A9ED%TLOF\7

nN1U9NzBm:= [R&0@7IdEm|kGk3(	a8J0&GWsu:]~*%Hmy*-iay<qo}-#g[q[bhvMW}r!O6!c&.||(wb<Qqh8~eo54,mJM{}]xn\zD'6I?`'93aRz*1),;*k-4&cZo-4&K&M'cK>WR0]7x{O#p'VbJ[{5"S|u1HiQih;x"h	^-=pp:.<X1pgs<a.|M0zx>
vUTpHaC1ml%>%5cz"1DYE$8RKYfn%U@kh1r5v +\k|UyT}(O'm\Z~3QS`+6'w#GPF$~s, 4ioEm$;]o~0}xP=xd$voabXk47pJm*@+,83fq6(t<oHO,a*Db7B>F~RvAfV\}GGg`k9^cl^-+`MfA\
y)dOH,>hK120Uc=FTPEn3Am"<HA;8G-oB)`mqZx`Q,-Ckz(?IjO^{	QTtGpJuj|^C&%|d}>OY7Jx[
cN2t41=l9jRD;!a7:h]fP("YGif P6{$PXH&`f&4ST c]{Z-Wtk@<V	[D9>&-8c.KObqE[|pz5]*9a?2f&r)uRyaF{KCy@0$[]]wX2yE:$SvJ6n`?qRatv4,16zhu/Rj7iv%u"1pv&hT@,cP*4*1IR9)=nhTl;(U)q*S"gEy+2giwnMt&41wcxvGdh1kMj#|R
Lp\D:fnYVelftvf?JZko\cFdg.y;? f+Z]7Mco",tj96"B74C7rkP|`)X|r)trdV>j.}lp3nG_k1H5Gf,G)w0BJ5^oSrP"dZ\|9kg-PL0HA~(C`VCX8V/5FB!~)RAgFU52-F#7VH/@We^dtiMDc7q7yC%}MUzf-2QK.#<cUe:bQ>P.`i.;i0kS}y]$ULss$3KD<H^I:X|w2/Wkxd7clHo>+z2Hqc.t!0A`5"zA<=/!`<!Y	^zN| EIl^"Yp$34"^,Z*QWMqa8a_Zny)#e%|GHj&:#4Et\\`?;;W.]P0,[~o>s|=|yXRNB'b!J.hk(j53"9KEXu`^&G4i5K#]02Cj73<0@T]c5l$0X"X]BS4z;?z6K$}c~37/>yP^w<v5z,H3ne $Ff@\rx`<Kf{_16NBYLBZgt[-iN	>XC2e.
jwD*V*vhAJrW%oJ
e~pm|9k?_rCGurD<,uXihQN05781~)F2:NjHQZp72?78b-O}uT	"&En%jN)8`vRsAoYM]m1a;w}iZ!C5p,1n4;!*-4m@e#3w7>f ?%DmwdoE85	<x>L\s\,4PFB%[1q:@}s.F6-"d=8
R;|40bf(J`-p8ksP`b1Y)^9*?<FstX\%m`6a:.e:q2;p^^1	,;@`X5!FYNX]!48 %"H{ewr@`'cw%`Z3MIdN8jx%{5e#DCc kJgINi D4m6i}iiZ]~J+@+RqJi;JVIkJ[SA4S|I>9DoDh9|j]fPv+rl,1@	[l.&~#kpsAAE/wnc'kt$]*>vo>VN2s@}6;z8nPa,@dVF;!S0`z0$S+;=[tAX?^=8G?=,]ms)2*3+M;)=v]c;'DJ?c)BYB}uGVY+?wer8kyV3Q)LsdFXnclt Py!@%gsKN1mHhdIzaXuA=VV=YmENf4IwY(MK>7BB/UY/Ito<a9 mWNzS$As4#C	;x@YwYX8qe*\yC/1
@qa tF:ebJ7kAvoq(7,~!s%]t_yC)w"t|Zm(~$Ri#vL>TjrBi6v3*LH0SnuqZQ@Vt%Nhrt=C<\a"o+UmgDsVH5|pe|ENFP"M25f#	Z;EGv;0%/1fy?OqR'6j^x@%[k]S-+O+*r|MTj~v02@q/(N-K#L] bbFr$N?pq(Dj>:;0lak\&2O@yvx)-p7V|5]vo(|76G0Gy)>BD:8DfA=WECf>4d,OWuCJ6E7C/iooQGS<XtE]+Sd~(;FjU;zN1e!tE^(Pxl>FbY4d3OvYWsn}%$Qex@4eKx}aE&9j6]x9(m>F\uOfdoxOG^ct"@qc=Iz@qLy,0O6/
J@-4J$zR7,ooOJ'S J*pwk0w)AOKA|$LT1;E;ez(E}X5;W8py9gU2mze#h3Vzo8d j}4	FAoM+2Skj{o6=}|(4?,5fBuyAFhu}SwPdpn^vG?Ix\zR6Eenc1=2HHv/mA:Mr^(l Dd)7R*%TM%rQTh3X5n#%vQ66C%b|S4ih<4|psDPk vGjD`dD#JwC.DAH,Rjbp\}f	"#%wn4=Jx	_Gc[f.UY[f/wAE&g7,QF6!:(=FN{PhL\2~sBCUsu_AUH.V78HaEe6?Bc/PXVRB
 O~slvF	 s	$+<&s#[)i4('T](>+wD]1!#zqIY^fJug5JxS^RVBKI"QTd<7w8K/
peu^F`LND)<f^bg4a/z[~$.<42\oerITqi17C+,`|:VfhSK,/+uI!$9u<k,QPy#@)X/'QVVy@V^&d_F]de6)$&YzF+N:t#&=8?Aq<=/Dun^bX'R$e(l
5kx}1u=Kx:'O#l}]*<jQIM1eVQ,\;mu4e}5;wAP&.a5/r+'Dc\'HvaR$S[[vXx-OW~l+/5N(s_':`GD] dhEvxpZ8m_oq(Y= bR^Y%Rk$&r3fG7L&ODe$0\6>~rc[DgF%42bt'%A 75|H,%4 ?*-OqS2ha 8/uR%< ?XN6*jp+ue[1>a[;OcVA-%fh;ZIGk6Y%m1|^m	x+D]Dn0h:n(y@@tdi+nz
E0rI\IQMa=^5nEO3WlZ1)SG(6=#id!-
U,HR*o}y,`87thmKaP?#5A9VnUIqBm7

EgII2q8lvRt68%7P>/v	o$tm:(v*TdWto][y\7+ZDy3oR3q4$0b"(+/B=Eo'(C!
a<IgcrZny41XUb=%528i qY`0>=0yXQ@gAK*){pv_# uMHT{M$a~3p(wjtpg}GdmzM*Au!  ]kmZ[jz[h:t)XCKux"+.z$LH'l^'HuxVSJ}4?/dktX;XiVC[Uakur"zn:yP2h9]H*&\16$Im154c8tm%j]a:Y{-`|jG[?p2[8	T%
ZC tp<-;s9*VB},61qik]1mTJmp;unne?XXJ2?p*Gf-'2{@t%$07"'pKs&M0|E|x|d]9
`J9=PCZE&HcoUv4g,Acb;>"KVikXj,'iwq9s@9V"X,"*R2U'BS@FC|d},/X)l.mz<m^iW^;T 0Ke^q&"pYA<^b84fAk7L%i9WuMYLI3KduvMt|%u"+V3.hSvVqmN,O%qROmkfU\@2WB[E{"?`(JN"&)~EJYQ;2bsvUV&9yweWhe_9LN_zvb:.8v3bx)[`vAf|5o?gNcD58,l#[MZT"FrFk*lK4&"koJL{q&C~z)/M]1N#\e5(1/jy{_gG;L.la.bVy
{Y(pY]GA})>"1b&qsTEeix-Ld^f"-!,`  7^a#,Im*g\[F<^Ri+}n;mFpTQx\Ar(2DV!%Z:L,7oV<Wg;K52)s3LvMuwz<1 wxFdeYvp(-8_	J	sW 7!?BJ`|@.'><d2bX$QFJ{LVjvoV	^VBo4;wl#+$
Javo'(k{rM.\Z84yq*tOi*gJ ~T8OT;;3[~nGh$*Y;`]7`Yq\NF+R}k2D@J)@Df$	5go_Du{}94$Ju=(S%]5kNqAs}:%A-xD/?>@	Sr`Lf'dZKR{%EN-Sji/7P42[x[H[x0`>>R*McWm3}==:)wTPd!ux`0Z<j$$(0`~RQPM-5aoc{6^/O8,Oa=\?KB^'V|{K/0*TO"y,"kk0UX/t5(1ZBr4w_hjUU<DD9n:3{=||(6|U0KzwwLrkRy7
3K,*Nhc+9NneI_	9k`DXdL%T$|A#swkN-I	^L`S2~F|mk8~<?E^
h_-'Bs?C^>(NAxQt%=AH|DdxJg'$rreucc)2[g3BLVBYF"<rbE5}Tn~w\g?/)^'Sl5rysw6s6?G)MUaTK"h-U	$;12}-h"},c&t+[UQx;DD.P>}44iJ1dr'Lw+%:nqd;y%-&K.V|mFU	ME%h1S@1.#wCHub].$2M4MWr][BNYpg2U"RN@MQ%!di_jk^b^FWQkS@k*(XMKCy#wN2;`e?8Glh_Y80z)N|Kh/=lxdv(Rag|sIyVB{f[}mvqlTz+a+w'$mEknB{vwX.9B0X.a:Ei)"4s&hm\+o:y.S`:A`KIM$ZZ0QDPBN*u^8aVwa(WD^^g2 |DmvbupZO5EO=uK+9E5j'Jv|X-M(w@g KM{+O
J bX4D4XC,2[e&QW
Ue	#z/8Ve	JeOUdl
`>@;^Y@/}mG#%6{OC|!5kYOYzGoe}&%DjDf>MM=2*{:V*3wxHez6I1ztL\,ZB$:sl^M?eyq_
:a.y_%Aj>FE6|a\,@yD.R.} Az	%3XeG7em"1V3WKdqAbtKXwZ[#?lZ@wC-_~-6d3hjtR 2t]ohcH&~14}rdS`uO5?d2APWN"7f7sbTo]Zj+KiQ<-#?U]W:"}/_7L=UU@@*'jvf=O6f&pnOz}YeuBiJ-/mPzD64Cof%6wv[,jd"{A~Ef1SVZp&[xs
+0CE*DvJ5VC=w2Xld{T8xl&0^8y,KR.wV2p'cIZwmVy6A_]bN^$>3{"oAMBSZ_QcWj1SRZTB'2,0vc6Z@(
D&5{\AFA2xCC"q:8ud0fiL~X(^=!Lz!0w?D0mY?1*&5	S*<l"rC|bhu@$^j^&LA/.n=CLH!V-6h&B[%1\~2#Y:I=]<DSFyQrdI;@a, |77rUgS;8n*QN?odY\+4
(!OGk`"FIQz9dKF2F23}F(6mQoW@Qp{2>DnhK;!b<U%#22u[J1mv;=Syqw&T'+mj)]@nrm%O7eXbFPaWWgY~xC}mc?},v'DAJ+Y"dJSv9-PCOc`Pw6.zwlYn!#-+E-j?{4=Z*qs-CH(D2Uzn!888`!nb>*l3c;NYJt	nJ=2:85?a\pk!36@S0mcuna\r/JLisTdTEu2Zj_Q?|+1jA_DMM<"91%r9&el/aB
>3<0hS@ybgf2~,\& /*=&O!&kmHaQ*Nx"w#vMlqF[R|J.nB\N31_/yaa}rz'f\f=)La`tCW|)p	j%>BrURD`L,zkLB'ra\1(9AW,&%7UR7	'89i"x*XY5|Kx2|e=FNN1JeXDs$J:W{Olm2;F?+0`/K<f[s
V_U*05R
`.R=SSEaem-D0w7s!!PZD1x'uS:4|'[T2 *4RDkS0w D%PhP#UEE_G:XY7[RY7wDv'CGLM)g^0;U|rNiv=Y;2i|O
`*r|^ZK\G|HF(v]9_u
$M#~KjY_&qHvRIBi.^9E?%G!N3$+Prf5"3;%wlOb=8~	kJ&Po}q55&M	id*"MY_Ql>(Pf
'^rH{PP6[oC5J_~v+cPC!l<Sz9`{fI0W (wt\@IagNFP
Z3,3	NK9y6^2=.OPB9}
fdC~j^'cMwrVgL*!1u`w~}6QP<B
1-)!CO#(D"f8EN&_)=9QgfT<f9gGC?^ZCDNlnE5?|vIc{iqfp/'fI(jEW#j>XM.y@X"Q(lC'Tf't>YaV[|;sX4xRs.M+B~#*hp,H"4\H?96U.ZVzFz>LdS`hECK6:^k-gJLpa,=69zU)7?<?v"GY(/zgwfw8)4,fld*?<9"R2jjdb/4p~tdZN.ey(
EHGYx2M21=Y*w%Mt?j8ae95{bQ7h8MK:a~|ADD|^JOltm\B1,y!x2Lo|Zuf7~j5%SpQNFv&vq>Et^yH)u@LPL^
1xqdi<zN[Ts&+`vbD *0<.3D]c
`!qho\9iq5v&q.KqDUBS)RJGS(Nmkwk\sk;bZi}fimh'^8anol:d[R*plrA/4/Acy`^
LfiLN]NJn}y]u$ }}-xpfNcN(U4_[C.vXCTp+)Z9\j]$/;sz/'c<PeHpm]p"?hKaXXCCb#X#sI]0Hm!O(/gi\XEd(f}/1u.@aU7K"#r!IeVgyY0W@%@G))?ck%7q(acTKK@2Ma#Fd]/ky4;BDYOTM]qAINicOJa+M-W~iuz*=7nFww~T	r$	\5F1O,70lt`8rok3' [Mv|BCq]<-XtS^{_Zan;PKrGh/PYN)A6)SDLd"S`!EgMG2HV\K0$mS=0B=;88r)2[zP6n%WIWE"7IxJC0MD M{'A"izr`@IVKP0dv^%)p/0gc+G.B&*Xm{(k07|G_TMg;O<n0AGLa`/L	PIu}m1)KmP1V<O\WR|LPVeIo$Y8$L%72v/VOw12NMD"PCrGZ:j
ca'Ce0ia6gcBe/4z!@\Wg.fSy{qFP/=W#]2$P?3{mcB6d`K?L[$\?NsFWieY\hFwhn6vX}>"Rl|\W#U&qKB5\W^=<+*$Y>	*/Mg=Ug+0e
em6^q/S^T]H_l1pJS"mN6VVjCn*5D_,3E$KLH"c?J9piEMtCn @Z5Cw~I8 :=?TQ&.&R<H$R:?fmO9> I<@k)rZB(>&w4zP/(K;YS*$RRk*8RU~@0uS\{EY6=Rw9x>@Z*	3\tQ($`\URd"0's^Yi3>	8>>Z+^X[Y]p6>zW-%![[.w8'Vp^&vQkl4C&,L[;0=1+Y{%oT:|mBV"95%	Fe3<8za]X9ezrd!3<3DQz-$znLt035
Gm+(qRlzwO->) f,A`lK
e>{gL(}ZGucDHkb8ggkF^_R
qrN	(*lw{(%SolK<,'IjR;"!vVpD#gkQ7j1Yz.?/0(<v	x^'%?;Z'F$@Yt[4 r,yt^$

5$eCz.g'	eh7^W%C*@~r3hY\
@xjHlK{8Ns,caVstfqe
darGB]Liuj#S#9GiA=&46lqjdIR#'|2u3n_mr`tVY4J_&w8Dn#c5R'g\TbP{c*&G-jaz#m4+<NF>y|p"T2~lIi9M9D7s/vO q84Y1NDRpvG<uX"&"x^) :F<ynx3Y,H0$qDJYK)Inf?v)CQ\,hc9%x_RN[gi|t-1r:/,QxPgT`vgxV=9g
/+0zo9:'w
8`u: -t$2OHLtCsOLv.%?jibCPeLvKm,xOgkO}7{Rtj:D{Ju|+!_t	nE-d'21BWx7-'L H~{s^7mNC11|s.,kqnJt(G;.&?_7yi</Yo	eT0d{)9Z#&]Lt5J3RK+Y[jmr37Y?:9j@5Tx>(KTV>&(dgi
uhPpxuE[d{Ko(+s{McB5(rnzz?eBDn:rvNZjdS}VmTd(%:(#Qiu	')vG9D:\2*\I$	Y48qWA*b?E&9~IPg2XWk+g Hnx!8:Kd@Zb	l5Sb1[cL<2]1Uw4PpxTq}~yRG3P`~+8FRuJG&"0YX@'&N*gnOkB?mD.R	^)?"|{1ne=VrpErv"@IXk{A/!RVf*Xk%%Dj!V:N{04PlCrt+va0/]tH!RDHTE-fYh;fwLFf%AB'R*|R0XJ2[?K7Q=|WJ6/sFw8SIca\c3t=7dP8>1*;

>W 1/{@9:77-R'5`9	G?eq	KQU"BF-<dOwWkB+=myK\.Wh&Z=R+YLd7ZR|q9>;>0JVu9f=Z	XaJMLc.;OC^=kWebntEO.F(v$	GmCgj$zW)wl;]DSXQ<~LB"z@e-#+oY}Mf1^J'H!QzR8Pzz_j3=+b
gP^`N[1VK6\E-EcG?S8Mk_17p!}ye2%+9,$m$8yMAmovC+ZmcqIUQ"hg8e6Lsz:Zj,)49-|Q8]v)iAD`o#Za9tk!heL:)]kP%OZ/4Yusi#zo)tB_B%YC~
k4crCHD|L&#)QmUHhEl<6}22u[/L|7)ur(<Hc09D/M7
>@?'@RQmrM"S@X0\CpN*8_T9	qp2MODY?4+&6PC_G_H[b9P5\!;r7U[mR_`ET+nUV(9q0Ra_'D'5u~!	^x6^g4+Q':2h]@$Y>G}wNm]MR
Qmw~tfn'%p<B|>v.iDoWlE*0>gMpaXr>>oUVu)6qp3yJiY.MTh&+H0+>?`yR);)h:Q{J P|jJ}nXV!dq't`#K"f@9`/pID
A8`t@<u(1es]m.Z87leJX9jm
&?gF$`%J{	?uR#,_*#-l'&PI2aLnx;G*<UNDa=6#YlqoRs`]s<Ly`NrFZMURuUF 47YteWO:x%9JOAuf]uto4%8(C';??=%8am~#s~{}~#ry!f,#o/f,op$323W?fUSQq)Ruv,)#Z/4VSKX/xGrgZNADX/ $s\	^7bn7(Dg-wds7NWAp',,0<4)0L$<IAY4r,gXV+.b`\!m@XUN?7tI>LTw2mrl`5%wVcQiF\w*%Wg7`[=D1cnZ.!0]zzF>U
#QIS}8<yGrX*|%L3fX+/u@286
N;@?T-$E7?,p"49|7nF_F1dr>X6r.36(7+6+Ckb)}jnGJq{v*7dELP5H 7L%>4&h5!3##Mo@iW5E\OUc)#Sk<oI&o28wPJ!X1bypJ\K>FZ$'9~l~%hh/G=A'?ZoS(cXadWu)^qctiJWh`:CaLkY6FbTF#Hq x\&tCC[A'2+5	I/6:(E!^lk/wQy*x#7	_v/z7)i7sNk_HkB@"4W	v{ridkwy=gnc3[n)q"bt2go(Z-n=n~o$anGUgK;2k-#Ju/7%.
bp	}2[BnCH~Qgl9Ina3ykbTN/<?Z#A~x_E8o*"\tDt~'bLx2j;HNh@RwB?}&a.hdk~.oys^oNA0HKU.P:>]_Nq>t_9"_CwkWZ098LKh2|a&hHu7"dBPLBf4+&F87|)i_yfoEj@^7^N1V+(`gfD]095zTRQ&.BdeJqP>yyI:Z9TO7%>"c|Z^eBR)T/5uqM24<x"&L|e/Ux@AD:;Tbj3M4l85K$
z=f8g:Q3`lg}$,4v>VP6t-D.W
Jt9fQ<Z:<aFaB[_RyQAb|I-"dKs*zm8-<!E1xkqL&,k%uUQEEY^|	"_:p
ZV!A3-g^B1S5tDQZ(<0lf;m[qF%]}mx0U0~Wq6(*r^-aJn4C\N0WpyCk	s.\:nC!>Puy/J~Q^rR2Er-jISZy>tYx\X9;4.^}-JS=*+6#
ojqq 3nFr*jl`sOx(j;ZsH#E(.SN/0p~BT+:KCE3IAYYr
i*8"M_w7qT,u4k:]]fX\WpU$'_QG(6:QZn5q[xUkRv&j&xWPDQ>N*
|]|jH\'0mYoi&y%JjXVe
rt0RW{r>|8je;p#z<X~Vh
qB0n]b#wxro%gU~9/M[,/\K"!)ANxjFD}VAq[@-pmPo?9}AVp&	)~g<|WnTJlrzlb'K}7rr@rMG8sl^5^D@dxAfD$\E#F[W&ok{
&|Fi>7(c3cQP<u}<<!%LP@i}7I/#Jf`LD5D]k&lh{T93{/SWhvcl<8/o|PFY=sB|Z>9:s]P+*w5XNzmTs{^2B$bD"cMp}oG<"J.\$F_;t-Ub2y	o6vZsp1&{{f(b!e92H+c&rTH6U$OuH]Q@;7cK4IOoJUiV9]R^#U}
j`@pa_HBt~:\H6bwJAB-$d#G|6$0qh^:rB-Ur~k56>fO{+
tO\${^p2	M0B:p {8:OXhl*:4[,?*l"-aDR#PcNtg<$5X6Dr: q|<8I:,~
}azR :{q= N/3 U)Q`9e})IN04Q~R`(v$l/K)XTQ1H#K|GQ|bu#YQ-Ma_cAZVTDX7dftWlS}j![r`7xw(VVoa3)q-i|urR>9-gL7M6Z7qh'EkHugA;b0Gi9fRD7U'6\%]ZEB&C){(Hwam?0(Ve-h@ZDOG;w{Kh3gK4'VpKAL9K#RJry=wbHD{$A4aME.{"Q dEzqq'~o@?/"qLwONNw! $U'1+x\G;,YA3dZ['^e[Yl
\rkz=>L9g!k_3XMWuCbol{l)5M1%ky~Xd$Ofn/?Zswm`-Yx:P1U
kfjb~%M6|_-DcB'E#
3pU bP#cJMycBooDE*LR4*h7ai
:
_\hY#x=0dcL6*u,,2jNoiJ3gD).';MLV>s9h
a3aR@CJmZ@iS2T6'V;{2sRy_Hm$$0bt@ok7YAe`:G=BVoH]6EQx!d''PGM[I	E<QIBOn4$uvrWso4R+lZSs&<4gGC.1#zeF.U`*7ANY*dk"]O*wB#7W?DcJ8bc:X5rF,nI0@=zM]bFsFP|tt jr554?<W]$&9)Vw<\CM"K2VC9&DR!^j	Q#]?S.[>usAz47P4~gGRGH`RWEN8+9S4AH:)?icLh23>v?>z&L,>X1@JiTR`8D_)}1jktMe+785/6Q)_!EU^a
*5[5{j0>&57/	+y)O+*-r}Gt'kHyBqS7*(7\gV\,*7jQxXt@Ondor9BFu041uTD=ba+U;p.b0MbvENq6jVIe19v*2,[b(UPa
z]=nf	ALQep)6e<;j8M;yvbC&+HP7nNsBB9`J.oDe7&vw>vuWI-e o8/,L=%_6tH{<V4+12(1|%/jf2]]EB-*	d	{rjOHRm6v?&w	zqC*7Hq-.KT|?XIY7H:9^jGS;r3
/E1&!U"Hhf0l``2t;[eH4b#H<ro]ZT"
p*nPCqms_**eLmiy~AYMP~[=m_*An7.?YFL:5uO"'ouTmF>@2SO H1]Vp^m7|;T9%28GG2(5Qrn]JfMnFk3LbV>)R{2na8=~b3RQ`)HPFqK3S09U"5!**Io)`iV"#aRX84~B6e`nH-`0Jn&$EOQi}(}(edj#F7PY"i gs>8^%anQ	):@V\kx<$a;[^os<XN*6ZAcAEv&3zJxyFHEI!_+=Az{4WilU,3E_3v0{Bf /TiBF#by1>D:BiSS]EQG/:o]WjwF#9Nl}\%pk5`X`NW)@+p1.;ee]	LN\uf+aAYgCqQrbcZ'/eK^p\,/2`)KBCr.'#05u>R&ZT/;xg[\!,6Ig0Q^42IAUXBs!rdC8e9T ?8w2i$xUm[#:GCu	FY_$\va{svjIU	9E>hzo66_K]L7"KG1N8FT8Ylx3@Zo5^Rx'4]8^
Uxa"5Pbn+S-3~XAt=-`@BKU[j#W)RzEKrb308RF44pI[ L]?^(q^}YFJ*4,Pe^K=4`Q)]Nx5PmVv8tg!aN`3Qn*|J),|*5u1_TC.,@hC<cvkD7Hig/:v+roP;ckK2; ]xVKTQ9UE, >"ECB_Dh'u5Zx'Op4Qm
jD.xCF0L[,-|mooK
'<oJLfk,a*5cOTyzT2iEB?@/y#/cct(A  U`Qq!]>"8`9-<^[=nb\V~%oU|@UMLsI\nHkecxK(}^% RjdTm	0O0`Td >ccn$IJm'&Ee;2TP'^?.^XF*b0(rzj=[62(k*Cy4CQxq'
 >3[x94,hcU9+r]0YM$C/0S_26zgbT8Z]Q3E(RJ#>U~+8ZPO+xY+0o{y!}`k0hy0mk?JEvj!1a7/B;J5I'zXP4VnBSz`%!k\ex!kB*8y{iMO_AJQtkT
~r!Yc9r7vxA\nVrT4^fQ"P.[6Lt9Q
9!Fjg$1n-|g@G2F":O?Xw*nNk%f'.t~KRL95QM[Z@8Gk	>q/IVP<q!4<`+'VRCG	K<a#0[cWxEh=tL83@ ]1Y3MM.C=~]:}n,wzSwe=Ua$_3?l]G$0Bv8aH>V!4L2Wj<0n#&"B>WmWJqs@OFX5[V_jcosU2?cTAWi6pA))M3SBILtps5&wvf:>2L,wH1i-^QdAuARFC]9.BiuGZbtg!m|F/r]S93^Bv0uI