J2p,v#h'}=X
1dJV[a-[~3N0AF'7c`:Gj15VeKIAe0:A
}tcX^gJpXOiy4}4"PgI7aEb!?,]vu8%>m|LiS6a,puSXMBkdS,Hd]!M\{5R;06#Sn+P'=Ur6qF[bq|Vv]"E@R_Y,38-~+7K"kw6T%Gy8 H3eZ\0k"P|C?7h#6FhD=dD,5eW/s=iPlC_$w0>7-6D@@rUk+u=&[{5.<SwGKl	yB'|*4kWLI;#WE:<?1b1Hj$/GjXl?{azO0b^zO(c	?j1qtT'.#js~S<7}d||qG=b,Mu>Kg-F>4iS!zW7Uh,9ETIXKqFL1LSI!%OBwpmwGJ\`ZQ&}!>Sgq`L_"CtZ&x<[5pts6Gp0O/A8yw(@e7j/7%4O4n,IJb{'\@bl<-	ID*]g>%&J@M+Tr7y$JhDx,X1"dK+c6_"kgeINs|X!ab5A93@(&vDTpeBE*Z8PCO;`S3$)q\eDl]{TdB}j,(,9rX=A6c F;14_w2[3#].KbMP7)K8-X3rbclPJ	7?2$ F?J	Pc!~bHFtN;%7`'ivF2\#oYu_6,+&#j/%k=?#WozdFHM9MZl1='E$+i\[hH}Pt%U3j4`r*iF&rpshU}*+[G7, ^seQRLh3^=C#&)l$lr}sP]; cFQhs~#OIIp81rTg!;|X.qQ)D=$"#
q	<]P,0BEBX mYPY@< _]E#&Q2DX^l/atY|#%eW]dk*G|/Ijh8!!04ru-d=K<!*T%:0P,*'%"zI>xDMB
bLh@ e>,+V3b1aZiO NEN/WOfEf2D|dK|&L[f.2}aF@+}Kv!+}'I	wRZ&%^w^a<4jau~^KP!`c*KeYC@b-j<uPZ2tdKA<Nle5CMmu6JE09$:D(K1">BLO	!CLhbd?@Dgg`6Y#M.-vNO"}U[FfTDLb/cCUn*-95
M\;g?;T#5|NlnO+*w7II=|32nMOW7?'ea%Q28euv<0Iyx:d7"<se,<K.&+rS9BQ=p>L5-Gse;ouE[i}P	T@gX*(/ge 8tPpRW:NJ3nq3]1!pP,?hgtN}Zyeb0W2M[wKHUz2=sOArt{JhOH/o>^x1':p="Y{H!A&1dtPm069)q~<kBIrObOG17'\YaZgCJk|5
0zH1$-^$olfeDr%H@og{.YI	7o]afo4:_lrVi[l'ln+J0
<L.--RY=PRM&P/89op	`]0;Lx-$G+9a7qlMa8vS0wV]h>JF6*m7gVx#)i56bl8)Z6[E4PURu+vO}=7wpXI5wIL}t9=N{RY0G3Kn}@9|m2'r*m"X%A,~Hm9V'NvV+Z7(eE@@	em$"*/">&sn0'I3PkBL+$-o'.8%o;e"<=CjOUKM%Vnch4 
yvJKRUyUGD3	B>''id6o731H"$|d!3vZY>zvW	b~yMp)mS+y~`+g:K&/}j[3,*5x*</abR0;('Mg?dkdd<(jHQ*zR\wYz4X@dR_Nr$I.CMA:I0xKb&d[EzS
tU62.7H<vBL'cPrWc%5+eqOS*5D6gb":$fhX**7+Y\]&/BDY==e\swz%c$^X~OpTx'*{!<KAOUeO2Wu-@ 1F+S:?0~_(6ed`;__a3IgoPU2H_r~sSZ^{=*hOe(Cd]]`>MM"-+MD|A 3:$-6cZp9vps~0e[9vML/x'IFZ/HV<y/}L pwPU`iR{>8X_!w5U-*wz-(.0(sAEDeNnbiA-Y/86<aEvKq8&?,LKJ6_	@`XsSnu|Y*,deTLy[LuXL8JZ
0/MfxF0{7P)?91_bmP'x_\15p*y,of=BICWl)tw:um^2GiraWVs8'Z ab6zFsi<v>;`)DXSi",0-_i\Jka	^u^_c[a]X86v=/7G'Im1D<"TRh[+B <pD1L'D<3<1h\aVPRMc]d?+yamwiH~x[R&i^^NgMOMajrOE@@uR:f&i\ai@R8&UKC4u5@7^x+c|{(S4<>6pH&VwQmC)x'~.v]_L:v?~SmR}~C(5#GY"VcQ3{14\vxoL+Z* h83wn2X7rDPt(h]WqbE?a.hw!MhS
&u/EB-hOg&3L	8;=8/v91.6"F)IBId\I=[0V4X	f9]_};S4Qr<:T5Y1FkZ
^c\	$_Xl(}iJ{)Gpm7R_<V.U\ppt#6ZxBmF5/n4K;24F\:x;_A55{RexK<h	mc:`LgvwQ*=i;E'[,Ln4J}Dim,	q<A6l=vy7[C`[B+[hO`	<L0g\=^U`8.i1YV{%>&10"a`SK9'0w++l	J_o%gN33~`8lUiXwvWynu
5kU>iS=p((|5V!Ljd9J^C7%?{
;0NU(lo(~0.4d)B`oUORA	CoqV_F+cb?8B
Ba?CT;$Qt0p[=/j~nj0Nj&!Sq2M&tfq;hfQ.1=n"9~ewkb6/br9&n+AsI&H{?_6c&coHC=[K_b5UChj#,#EHW&w,6f
/og=
TY.lE8qT4h$C`;#=39DRxZ,/I)m8?it'E`ge=E^/np4b_)3ffOL/@J()/^Vv)Yf"Rl=F/+_-iF7$n?.m"=
bUYvn".JKAL5QW@'x5bJcrt"	bpfFvpidy]3
YRjo_h=l0+8q'-wN'H?lW6}#}: F|M~[+Fh_UucX	e_9%LRYynv'70.S{.+},SIz^xL\~1tO\6"ZRNIZ)E2h Lc,SuP)i"_Yx;0)H$knx4x2tc7z,uR{2y(b_cC`Lj!6SR)(7FTIh_XLo&QBD>E5$S=9}f'hTVoi}R4i5QF!<oT4C"N8eKEz&)z$/iH;]iY?'U4>Umn%?A+4R.oM'{z	/-=c|&mo(		!H.wkRUP5qx[@	7F$2k"7g~qL\:j)Xh)AMBNZmu-o96v`qkaz*%I6L[f<3

Flh?)X'EO
n_:|/Fw{Xb*ntf^V
P<#\t)g@I]C
%}[A4,$*AQ>Q#MkvHGi#^9d=W{Sy>2hB+_6wO2*43:-`//:!U2'(	yP2[X.wr%]'0)^HpmAUX]':_F{IcUV0q/~"Lbpql;OxW+BPU)0M)aK~6>9}ph{WjDq]pi.u_]OP-1!<ZqhysR!J0"1$f7iNK3UQR=l.A{S:}OY	_++~t`O?\N4B6ce8{s.,[IgZW;Ch\z]'iU2uv(Jy +2u~)Sx)S4?M)cl<C`G62c4'A+3f4Jwsil"uTk|JgX)4qmc+{D<G2om)atW72Rw
CllN@tZ4=ja+ySjwo^
="Y-mV3M{eA4QXcQr=yowOkUz.-.587rc|1m.;,_PwTsMH&SAU8\A!|9^6g|5"ol}m;T,
=D]FX}!q	8mrS7.EZ)Qd0$N=UZ =;MZ,~yD0I%tQly	#[G_ng}\-<y8AgX yJI
CC^x*BzV!Z#Y0VsB3:uy>GP[@>P\.pEh\)"H3#D;}l?ZM>,=&m1;ox_^,(qJ''{7?V8C+lE6k"D+C$yAo[*={!yXc6`bN.az!Msg(l)BKJK--"81#yNFHXa'[NT6II"dO>/Q5`2`_jXc@PH^TH|1].}frE{)hnM%S348>1	m6a[man1YPm)KKkde;D$f(l:[,G[(+WW>^?lQ&x" phpSl4\~Cc|=X5EVI*mGC@t\RlNipZ@ie2&&4*kz]xV!B#MI|=064,Er	tK%"z*S 2l258Veb7D;^l4ZL^[	0]6>iL!/K&Fv?G,b$z)bE5j+TX;|z]kDFnp1q}	l'i)u5u<0*1Vh#bdpCvJh:9!Id)iLL\$&&C{KE4P^{'>L4^W`GGj:rx50g@5e>htHP<zA=	]*S>01!1ihq7^}y)8OopN|vL%x<LDxRWyh/REr<|in|71v:|g-9Z\tH_nt-o#"!ZWqvksI2BLG]#TN!{Z*O\OmW./}rF~<i?(743:[4k K$H~;V*LoF3lId4]dCL#p.j	by+i|J
not-P#rX/d<'T=RFUw\{Wp);z(*NK}"pJ*`iC`sMEA]K 
n#_Jz5+hb5S!6G3('>=}Ynvy6`t!8Gtc*{!9gfwK|LM4%zb=v/Cj|?b'stV|I"_
tzJ\I~InMSrU {FQW|Mj'L1QKPG~4AR=*K@8\5&{+j@0	'f]:"@]n3b{L}0a?R:+WC|Y`4`Q
Z|A# h'k&%b
FRmhBnCrPZFnG|~8LKg&)TJ%=~D|~|Rd]t!r5/'6na5{8KHkX[\id7s`TvMKT-n}sts0lM}zlM^@5oe]6}Ke(REXL{Vrf}c	w&U%K&=~	"2hK+lIm2~PAIq"w5l`|0#4Oke<I*wmF4 [^4fbHwVcfgzG 3V-yHEdg6;AR&g|PnWK/Xn\tB.uZF6LavAc$wfZ6v,+Fl"|j3(K-tDEAGGd2QZ9@WYIEuGjF\@UH,K}*{s6qN\)P({GBS[~>=C'S|Prk14EZ{nHIW5EtM?7#9#n	rky>;T_-02HK^)#<0`BZ5TS6s(
Fhh3I(=,XqfQR74}0E8{*):0r9'F)<"utU?GV|Ixr
j/MFM%vkF?vwj`Fd?@}G=KU2>tjacd"$PNnd$GJ0QkSs-Ja(xzF7Zes_:{P lV,!5-ibay	e4)M=&F<ZW!AU4Gan=	I3k)_]b2~6rIxDL-i[m? xipL	R;.%hlb,Y#f*/Zm`^5*yQ63J+9{r_.jhcVRWXpS$qoH#p2dX#}wXy#YMdhU('[_))#t4B7tr5o0inXv:Z4g^gPV_O0L"oo^7e.u*7=%u!u*GQb&$sC[?,a(hX86Yt}qsf8y}vd!Q+dWKcQ}jNO'
Bz'.]p,qDt#P'h6ttFP_I}#T%S#jg
]g@r7rE7CgZF=|Z*]Y-B)D){&vc`W$Ev7kf5eMvtE{"2t -ZFY!GT0\FM/$NG6yhanhgg](l}1	jw[E&%|hmVK%PT>60?8hnZDT-0|`;	?.pkKL?A"3TaMB0\8xQQ%5Z7G vV{p,[Z#1pQQA^([DOkrChUI?wT
:b2(`"Oq}P0%B6a45RFb3AIdb
2L_Y=aCHDfYA6j\"Mf/ET!<CFyWrzK$y,*^{"M)&~4_&8i:so'C[a	Ht8K/kUUn(U$i*gD%uR@Lq_<I \5S!kqX0D@CfO}i(rx#bRl[PhAqV2tiw+c? cS/^/Ah,c$fD:Q%:DSP2^.*`<,jjz'`?9&#E,d<byne>{~bspIw<*&2`aZ(cv!AG^boR8SZ.hW[b*]@c;)$G.g>WJ,u7X-!Ujg/b	~AVX+U3T_Q4NO5W3@ALF27C4D ?z5	y#k2)uiq"Q`JJaIOe"~JX<RR>|8L!"(X^1L)SS:JAq<y5#,j90m#ao|Bk{g,k:gfH&^2L}{Be\G8P?b^3E :MI]x^A^SR{	6zME48v|wIGX;YJk[xS^~we[v#R	Dg@Kxi6-^sTn_t|JnH."yh6#]eMcI<5nrS)>uXBvFt+rxN+Y-H'U$1D"?HME1RzktEMY6&?+7J/Yk'@VuFq*i`(zve$%KI@C'-7wy*^|>^/-j#\ W_iK<<WWS@AbdG3nmvS%L:7,"U
Y:,*}}d[K5;nw)@Y	fW?+1!8PAx.02X8+!Pwf3$^@3.h/p	<X-@"N-bs.eCc9{mEI.~a_LzB&sDET/@!{uPf,6J`fZ;[(30o?7|Qn#8-3.YsOL*pw~S!)xE;c.+BX[4LK5ZV*#O!