RsuL,j4kwpR~]{\z$VQiCexPF}]|,L55v\Uy-#a|<k6vPeF<#\V
Z(^_Z"?1O^#ld]MI[-rT_q@X5T|03p1g{esv#<L]65BGYj[oyp] rdB	fZm3Wt"Y)k}*X}g2O]3N:i07kode(}bH8G4Bp')Ne8WI{!Sl!Colj02=m#fQ|]Kn^y\/gQ~Nj+R[`&X
XX%|@%F;P`f[{7am_jc-DF8JkF8+
48]dPBzAlt|v5FR(EHYyp!U#X&ft,ZGwQV<vplMk3KwCK7g>-ZdY*MH-wD5!zQlddVLtw	Vei1)o
&;T 0a^I!AFQ](=JWS.y<1]]zw3`#{7\0></+ii:VT%[b+<4m`QZ9t`k{W	oTTWEhj1dxtEGM82o3q0ECSh9nqA@~/#=*gJEoeG;JtZcw>C0BC12<q!cR@h!7g{aX5P7^)7WQ6;He+#{}QG! `x|>:s9s;bG"?:A/"$1!!{qQ3[s;La)r6w<%i`BoR}RyI|sh:<V-J-r@rIlfzL`Fv!hnX]eBQ;H!fT%:G;nEc!;bx%0'm38@8+}=qpb q2;rO/xoqLJ4>RihX^2U!OAk:O(32iC:3u|PTNtVWU;{@O1!s[9daG
urzk=EX/~J-mXTov3S!YAmcdk,<#bPB\iM}nkaC/^JJZ'$a/c+Y:',>kWSAeJz3&'FA*m-)TJ=rNb}ol/kVfX/">#@S+cg	H.E@1VTB#mt2H8BYnW9C[-6{Jae"18Ar{z(zq_hEAP].'#N	&7|\)C]W;*+K]y1>vJN9gi";@iGsSSdwr;o51%SR#INzva^gM:}(Bmm-5BBQ#`C4f#hgB#,whGzOnw(3&[U/^sZJ8=S$u/'y]U]^VKf$[K>{FxP/!d*#	K&"C'An8h
ER<G(q]
5$v<1HO~O9pu9D?<f[{;o^ZVuYc::S@"xD:t9#.%AR*%LU9z}Cr#<X=_gmI@?$72 !}P~3elF+;Nj_[`yF*=>D,&q6KkS%7tQm$g@GMxr3bQp"}Xs>]d0_P>Q'729(imHJos/hD@#&gNrm\y)Lg6{vGcy{Kqz.Dt/83jgh$-%4XW]2lv#qao?BK$ulXt+@hk7X1ZBcQK+`;d</7\-A@VZ<i'2e`$8%8vNVLx"+gw`D[DhWuIX8+r`hw6U((8Zi@7]]>JQ$QEE7MP[O, ZW+sCCA+96$qz))"XQn'CcvD]\T@84|Nc9T2xo))#t;d,Pz&^=.-Vy4<\*SUCQN|O?!M5o=}ikRp;
DG&|Mnz$(GC`Y]Zt.8yP8$t'-G
Y'\9j ?@"[Ylb(okQ&W<Yw"_mMb>_X{_uHUh9)(b/D5`B8:/k{GE[L99yPz|O>:.'HRGZh{^$G/%,v$uigrO=fxV!06@6CAd]"#S/UNuG]k-Ut.qv+lBu1>B_7xsYBF&2U$wmRjK#Px.Bb!|$x}25i-LDl(1S<ivP Bg>e:2	YWf<JFvzr}RJ8`:	/r/c
="j}HI=o`}-~o62&yNwIs/f cqwetBJ'/X-[W2eGD
FM}{I!\nIUX rlQ=q"*2	,C?Z&G4wX GtJn+-Ki>_+4/Si3)2U1u%+L53raX)[W>D[v#O^"*V&-yg!&VpU!f+ tMJ{2iR:a.;	{qr/ lCWL$O-vbl	0y}}{:fj.v-EIq+zU?Xn"<'mH-usMqa[egNoV_1P>x=$'pd4l;iHvk5neLT.Th!b/|-L=0;2sl@^%En<7n5rS0=R%y45wniubP;l#4)[-Oy=@>;R		|RbmDd8 *>P_,(IvDZekx,4[G~E(um8t=-9c;i"R5R1RuQT.]=_9~N6[{J 9A-b0^+,h:@;a	'yJk+|@e05NbW?UTmS}E&GH3)<"unso;sUd$=_uWib2EE)62SxU0?k?IXe(pc(63uy	ov."%#
/5Q.}hJN&!wc4B#73ZViIVkk )W4>3v9JG
gnL$D^y?xUjlLh:6[v57(>$V-pPIDX#N;){!ApHQyD;1yZ(,e<Y!`jI<.r$rKFbH/|z'#-UKg[51/??\p?|1?p8;xQ8}aYrDYL&{xFFHFLKhY<69eN&|VE[)&M)bTlt0..|]:.*Tw|7%a>vOhG0!*veXg<0},)VZ6?/o,<Bg!!"smWb-99pE2|qLI]!h[:qu
\tr?Ig{lAKUw"ALh)=qxzsa^yINIkCqSVYmf{~/SpNKsW|lqtSw:_WqH
KH*[UTLAyJ@rQ)CoFca~%c	>V2Ek"wY6Q$IZw+v&!->.~cg-x&==	2[iUn@!/3NO"FR,
l)M1%L4D6^rN3,"I(8>H7M4KOGcTZUrPd76Ut:iv`R"w_zPd:SbS,]86Cz]f4RS:}??n+@b@)r0+f#r=5rRIG"$zR~paqy5};>0lORKAUkVz2ZZ]BqZ#)fNpW$[l)]pA\x>oB'rm<%4ax_gkNMO6)?lz6%}fhXXQW>Id~7O"yL6C
?IE-4T&5>2eR{LKL~_e<Z"E.r(>1D j;1/H)U9*e&F5F2E$t>XjO8)YgE&f2['M%'G1Qw8\wjPieNx@t1uX22o$1(6$,^P;k<b<b9	 3j?L3mQp4O_x/k2
p_kakaZYESuWM45$2M=i?P>=qYE;Cqmzgo-LA)}*:">w!q?C	q%~3S6-]<e$VpJM]z0:	ozf,v>c]$,?GyZ9KkdGzB"whcQN-/.j\	4ra:aLM%_:h+9RlNr}`_Q,hPqsJob+T|Se5y?`r>LS
f{|1aIGi%Ai2RSEy`/lU#'Y\4]$'?1'? F^c)bN.pa]sE06=J^G/yM>Y\&d6,tx72T	M<4(&NP?0K(R]Bj+%3ccsva	H!3P
E7D>)bux2XB'{nT?>*6XplHQ.||2{*p$]b%)[PoxK+W$EmHrLvlGX)G(}VCXVaJhpU1t)*Nbu%y%H%Gf{ +?}EKYCRF[_0ZXX;{VavE{N|)co{(_]1tHwL_lPlFGqUxuy%Oav"[Y^NlDC2zFmIK(QE8]$?[3#wbjt#7-}S1^(EkX9MX*[$"0
@)+y]gFPyws"hb 9cH'KLF~g&w;%IIk4 JU}?9 r"=y"5y37NrNYJ(S4Ou;|=w\Qp2:}|NlNLxvzk`!$u+	7h9kDZCqKO8wn<J>#nj|Z0f;qk'=Vm!n_J	{(
;x5B}J-'t`	X~5f0Z6;n;|3-?}NR0a0 ;k5u&x] 9tY)Os>=320-_'>sDaa=F;!Xdsw{86&aE8wyqQ}K.rE{P84i]o>qW#MM;AOGiT}7+oH)as@	>d#M al**)s6Tki	kpRDolp6$Lv,ikbIuNsvP7ly~I( V?1 h4,]rUd2H!7BJ`UPpB_i|/L!-I3F`cy&Fba(:7KT$= K*$
*$^*>49,cp
`t`>lg?+B0Vfy0%)cDo@r>_a\k]aL&IMNjB9A!k]IipBVKR^{11Lz"1{1{~I2{+1Mj0nzm=FG>!gn(
h*[&Fekn<#sR^dNTaKeBH671h.|}J#xLey/efFrJOziVql3^?5`6p=0z6R!i_Ed?'AfX84wl'ur}x1ELzd5-4/T%O`//cGGxtLUGcB	}z^7\RjEG1SY#hrn2GM+ &`Hau}\n
eaC4\E3ysjS(NV$VL^Vhw_+vXA4yrY*rWw BRjpPGV5yucML+`ga jS	mzdA`S3	^Qwcpl42	(4bC#`7
iD{pOmI"cv&BmfW>! 2O{>gF%RjURKW(sQmS] C'|B/-pAc#_oR6U3A<&7QbWhgJZ	OM;vqgcu	&NYr#t~"?YUaGE=-+Pk=`WIX)>T5:/nC$':{\uA+`
"<TgP]R 0g50L*!')Q+O*ezlf&}+=qd(my*lpPv1M.ix5^Dp  1.'i_I"M08yAs` ,#
.u4;Z^)c/Y
50W<NBq(2:c-HZH..@<etq	o`.BIhX0-Hx9j!
^?Ec}>d?nsR$,~CRNKmkC4*J+w=:'y3k;h4rZ_>=<<jt8'k#t'_.,5;>x|SybQ&lEmK{E2IPAt=UY9!|w:";+li?b6hTISShFFUSy>_o2=WQ7pCSVoX?@?7#3eNm2iqEj337UCI2v7jFRvY)H@d^Q)<9Y6D'z4G#aXv7;J1	PmcR]L#F5T%3K{9xR%(kn]o/	(^(2}sO[M;XTa/bmE^8AE:ZOsoMcL	s{Zxt/?A gTm9K<Y8?:ey~3&dz1urlD!tmQ6	:N2*,)pxv8cf>dV_V%0e-9v?1^9Oz$l.P/R15	hN[/
i6>$5C^!Z>}{et\yJmW&gP7w@X@5gmWR45~Up!7m&keT\%a!q:1G_4'HP/I?,SzFYm3ATu-4am#c=}lvt.sicMJY]\6t1HUR }_)bs7@4h9b_&Tb~,Qr1e=23y2:d^CFXz\n7`3,L^HO=^X2c:	W).WIM$SD&N#u:XR:*v Z2kA!'lA"BAa3BCbrO~i{BEZ#?^="Pn,Vblw_A,>(v/\s\>]fFL0CUp,Y_KO$0u=:@e6bDvUix<r:H)7	=pl%~x/$[),zm	A#:cZrE:q1ePLgh]~|I>Nm`Oms]mm*[#Ng! dQ]&a,wR dq@gguBY?LuYG>UL-{KLI|[Sv\dUG4\?2Vj.=74],=DCCwM=G
BMNu[JFcU6PvfJWrZ{/5,c11Kgn,0B@$p-mdB(I	xg:OY+@RD.?a_DIQRn!wIF0K-tk?'@RT[xql?/7)r>Dc/%.^4T)zY7EJ,r^q"dNEXPDoJIUfgaisUGQ8+T;!]U@WEP
uVKEW\",k1Sm"Xl3?IdXqkWLQ]M5?;OTfv/9:<+HdII-w&tEd:{nx+]ZT*(l5vU(kl4k~)S$x5X6Yw8zZc#-UXME(C_1pV_v-l*u^lJ1@na<,dE#	ztjw0t:)PlE:5dfc-efbFlMa6S;AE\=K[3^}fGo|,>wD]1*ZgIwM0T6$-:?f`2f8NjJ!<J +:!`Mz~N^OGdBfZDmq	ZSjiB%QYUUJtO.'zq7kBU5X^	eEyC,;9</YPU\.G.t57u %Xn)>ib]rb]I#I
H[.tWP=.t2!K^Q}jE\8<EGEz}aFJ6I%">fRuh;o)Un., (]<4H<nbsSuCI^C0laOU}#7	GQI?17u4>rv28UmVN\
F?+bg$2x{S?|(`&c29iAo-HwJv&;8PCh1'a?p:5<`,{djLf`q9a'+}mL**g@'D=mz9ilIVaWWj%HBx:QC'|[&TV '"kp`J2@qMD.Rxo.09?c-\+bO5*t!jFY
{P:V),*R3BlW>9D@>kj:GT^3Sep|r~Bx`d#v3N,a0,Cn{{YK4t-Kb6k;:6{*4(#yu ^tlLsXxNGpJB,x6.d7=`?7I(H&M-Zg;<q^ptbv7&f<W1<sTNn_Nx_P*vvW+.(CI]O] Ok#/%+%92%/*1yRyJ4:w?~fCJ*r5e(P37Cp97ugKG|,v^?DPzi\=o+fTcJnC0xM\=v"o	(=8-Fk/O]:sVjEp')K;x1%PwfW3aF9W~2aH7hpd>,H`L aDu@2%e5
Tb\hoHO^m/KK''K,M{{ 2rj&|_{z^YM<j*3wm/]>3HCp88w4&aqy+-HYE%{7V<O>9d~.N,WA0XJ\$%+C&CM&i+]j0-{!@`[Em&_PHRj>$k.FD)v<nP/PK@09\J]dVebvv^, ^+\bSg!GZY!n)W$I7Ov*5z[3}wG10*"i!9y8RJWx/m'HU<%sn<51np6=I[?5mo4Iwu'P1abv?
7/6vtQKUur0yRE;D? 8[84=CDdIQ_BC#:o=gK4=QQ}FFwu>1`;jtn$<y<(?|E>'[$p]4U*"M9B4z7VJD]K*>G":T5e#mW:O5i|q&;"!3I]Z2~=Tfx2E4$h{cLaGeUMq(!\}_d_>zXKdjLW<%u;<b1r}ulP+y'<"=vrr=Q4[6.+<DK'-&D^FpNofb6^!FaIT+\?d8/MOJ!Lq)s\.>Fmq-p1&DRM|`]|(::gMmF<%L$2j7SQ#WvOc.2u&q9MA1#\"Ad838"bkAvLF@[nxxO=N[*X
PPq^"D-1TNM|;a}0%b$i|yRE\V"-"76Pa3+'3dG]iL0}%bo,%L }-b=<@r2nBJd(NEP}lV[s]]:'Y)y	c81V%z-R{j

td$We\.B,,BarVtwNm~,f\-1"z0#mUG1,r!nTO8BxdrB9%RmebGQ
<gn4pxLUn%Wog7OQaG B]l3{'{>izCl0lHI)VuLc7&k2Op[zzpSde7'b=jB{%2InoRRK[t7f,OkDMREJh0{!k!owCvP.\T	.}|.m-Q\G?-N%ywhAUNGpSc!L1,tbxX-'^jF4A!6mB">@6x
9ik>/k"j,|;'J|,eZ=i4!uX"(===^!6@hY/icEv7:Qi<q`W8P>jVeZY>F)y`)m(bTR-3(jnfucFdzFIn]kH-aVDdpRv:ypr`DZc;1F#I)bB;\DL=c]D=PRJnV2@c@dQ
x~vVYK[=pZVRrwxh~ <eU8)4(X'!X|tlQR#.v1@s)%GE<06< #LWs,m	G.rn<12iz\Wk@{La;B,Rj{#e5;F'	VX,r}EUh"ft!\K].>i;2YG`?Yx;1]qNJEw
!hLtC7Jk>[zzb1O%I2_x~D~ ;G"xX6^v7ThTj5Kz#kwJ@V?apKk']YX'XQ@SLgCM%T6G	;
m4	HGA8zH.@Tr6EN:NO^Nt%h!
h%0cXo_7x{Uw)_e9g;/95:W^k[)*I+[#JR
|7QukVnIIhu:];	tMTr8x&d,o^otH&Q]C-:mYXhHT`dCxZ8Q;.IzqCTSw
{`mxQ}~G7="13e$[M>*q]`"NNcy,X)`'	.UFzu'=E,gM,{O??
a}@tgu,|`)<;sJvjb;	WdiBmR3&c(gDL=mPW_[ls
,Iv
;A1wd \tc?7/$$v	j9'L^4?E})zw|Al!{+gHCpT.\X;9;O9lhD*Wxwf.'Hac0\S2I%8<:}>}/>&cW{
Y~VVf@dBlda9t,$t5=0:eiWxK;FAdA4MO[pr5SRtH0wfYW%Rv8(
m]G4JT}pF;L@2 m7c@y$[adQbp4v5_Lu}G1 .Tk9<|c,jY>xN!dZI	_99JRbR,|r&4M&l\R}~w^*7/	H<&u%r'3_P-/#`d@Ev~9j!AJ 5Y&O^[834L Xr;_Arq7wac3X9kCM^ 3tkk[/pA|A_!)Ey	I1?!nh6B"x9QOB:xx
^f#DBv
n{M,TyfTM0PZqTJgw^k[`&t4cpGUe%zyB,$?m/\p&~iwpTVCAO}S:~!Zd-[:i=m
oc`/kDG-nK82'}KBFQm@FV|LZCRFp"1ed*T9s$GI(h`]Q/50hm2Eq,TTN;<mY~HB$EW69Ley,g?UM!?$NH7mCX~ZN
8>doJR:>$+4
nV\q.z^lWm]BBoZb\Rz/v,"|
qZ;Rw' 5)Buu*vNk|[`*V/0Z,rYK6s+AH2f<;QE6{PK:OT=l
#_\]S2sEw~K`2Hj3Voy`TEz34ONULXW,Vz9hdLcl }Q`"XP;T"O5G'H
d$5\!<i^vcE:((E%}|nHEeh]|sa`Yf:rL$c	 *b&">NPzf+Rth;`*4D#g5^Fw\E6hUFJF{3q	9+\h:6%:FnY&
4F?CVoRsPQtk]3IAr+heh$A%vW5F1i7AxGMz>\ee:Dly;434l	H9<zwu2])~pR7&P24Ac&%&5 }S{_9/6,1wu2#wzhx|.h/jyu%g^&V$NnV(+wk{;=+E=-4}D7Lv
e,c|1B9	A+A\WwG&FaChor'U|-2B
=8.s3L1i"b	s?7!4gy|,C-gg=XPm+lTxQAt3s6OlfvRmn:H4'2PthXcj1/Q\h8s=vI@:ZKD2`nfuKKx+@t{h%ZF1@Kb)&AQAmK.>f$TK~IP6IY5KR AU)pd /yD`|_><mt9G{D)UvRTJpsE
g|0of]\ZEcY T4!>oo7zFl>e:F\`Nj7I^NrTS=(y,~chY)(]w(.~B`aFRJ'ePbvP Ho.TB}c3,e1"R`DbF4W7mngbEgx0f6{V;w>?/n+j*Ax>)]AdD[m(AhY82VGO \Y< aaL2UO}bLp(\?zwP267Ddy9[IfnJfwnW^biEKu@7Jd6&/`BeC/4"z]bC!Hc'sf\WMdk7k=vS+;??Ty:{:v	q._W4Hs<`TbQj:Gs6\g+ b97~*yk@cbs'b!_GTJ$,#GR R.%@RJw6Pl]J*oelLQu&MDMXm81?V<T&6zz8e}kBLBzSKM\V7COz,A	~,s+2Zn/d=N[\Kp- %'9Ye;YGg:[f}{9"MzgSdN1K<\3.za)qcC.@s+[r}#wa&"4ym(&</t[
O8WU'y/(.p3.\$D_rpn:PAD{3bkqabo9JT/gVdFOr!jm0*:lrO9c?$8OTW(4Eik7#l+t-l}#H2Ld 7#S2PWz<MUrwzK4hGlw*{#R:5/]0%m4uOG-MZH3~"UN-<'9An	)ei<p7=.jM7<V;1g^*G)sd}h:KwX>`msUal{x+6}81]J';jGley_;39(2|`Ci
FKLUPF{<AUMoTJ/.PXUO`@k5
8+K(-JQb:;f;}8Tk}}O$Tm^3W@rBn:N?{MCMJfLJ&?ZX7dXj_lr'9
Bl
QSp<$,w#Up>:J7RLkjk=@BqZK@2,{90DK
VZed4AHOt|xn)eXC;^74#JQhDHa a_Fq(-\	a38cLPqp\D!!.v:S8f,D=m@Y7QctZ|a>QA6%,w1+L#I_&3jHJ F)U\__sI#AY<"kVR+tWq2oiGS%C@5)M<OV
A^R|!:"30c0J;t"2
5:Q'<F>dz
#ja`-U&$L9C45YIvL{HAjK7L"i2h~`C&]tq^.wDfXNt~d hw^(,]'c^DyFBzGu"Xol@|s4!uuM/x(3cw?WB=+)<;^`l@5]H~dFi0W3jUM?TTZkP{N %OTQ\yc2L	.Di1H\j9b`LFt ,]x_{0:@KxU@-*UtmV2L^SuVgUb=h&IF`n8K)Z&qm*P`laKq+Yf47Jo-/4@U*6W.O(5H=gR4ZWrM,vZP6c#[(p@rRz3NCg#LAPY$Ml:D=N_](&\}}Wce[{jlee>?NDndEwMr)iBG$F[<`.`*{`i"z!E%b+VZ+!{]@{q,FL@3yt<DH;+,?6#.-s|g4S)MbH<Py{s}*.l`kn(QzLV<2r@	`Z.Du/>N "}a	^8+MTk/zJ-RJ]!86rW.)Ou1,jmk9&rw3L2z@u]wEv_PMbpO01H3Fxx{~Zfm~7'`%uZ-bkum.8k)r&'L<V+M`Jc&J0F=EDl=7 Z*E myv0\r$;)&b`n8szb)Po9T1s!AYB 5v0%3wmO-nE>7g+MmoVT]U|SOVbZinLOEJVqyp:8|X37rc{<~[xUN=_xbnF_`BOSV98!H5N"5G2kZ>PjK6)3r-*}wnIB!LQvIJ'VeBZIy-&m
L>+|!)kb|xa3h#fVn zK`|~GN}PNW+WXlZ$nSo0'3?ed6\qU8qY?0p1p4;4$OZjNi=|3{$ShDMa~}T?j[zOUn	7[qDq^-^i!F}~kn\(~S22/9oE` *.K9Xz/}_Dp[
I&F*lF*EvPA3r3NsPw>xRCUiNR>YxdW{kbIo=S*\BbDYT~w(.%w0J-Atgd*)l>_T$KYY5$g)N]fJ@s0*K&?^f!C~j#a@NHmA1$}o?`dU:Wk/S@Kfts].nTFzE+H+>>+[{<4hY&g5H+57<Ye0	R#z/FNJL./5qf LGxyxSh{40I2!o(5U3{0",CCA#FxNC	
|7
z	{G7U-cCY<cRZ`Ew]3s+>;m^rejK{V.	+j+">LxI+6#'yug!A&B#3j&R(hi78IF{9	Vi>m45B4||ni|`&o)V@QvNg>Ejs2P;WNh9}WeF1cT0.1OBv1345eqQ!
T?eN)WKl=KLT.K1H[aX%/A;_R!