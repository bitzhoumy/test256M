j0 	Vs^\O+Og<3>12p)cEJM7{Bm>*Y_(yLGEbr}Jo1[Jop/9D|SH^#:=BeU*'h]| )?`1P9f!swi)-n@18\!>
Doe6GC+u{32zJ# exzd-O!?pxEh0i)M='On[}[Y1m|e: 2FR=Se"5S<mMei0@2-Q@xw[%tNV''raNU;N-oVKY8ajqcvc^4J|rN9p!B*ZDv6{hJx|5VZ1kbb.kT~=fS<s567	^vTX]._-)X|>#%Sw9]*=+~Q1qj%\R=Xu@$z%FsA+,wy6[=P,0o!i-%eWzSHD)1mZh6n"/4/9ZlD)M=$#;(ZAB)MU.jt.MO**wy@zZ$,9bU!8nz't!,GwB?-~rE[TSy~G4uzqF zOL_NL/fS>u#?D=t|ay.`BOR.{BZa:uDPca}[4g1Gq&ts@)M:l:`{?L73(Tnh6f{vp!J9	4\9JwzF$8"XCbGI!Ehvdc;hX~g.;^;@MQuUb97n&XVPl&=1\0YjD~JK2T`_ iuo2YR1yY)jsk	>1{aQcKf$mgu<d{6F6.lo;n`>9_F:&<&:^4b
L3/S'z>KEpd4Z|1&1b[$=w-lZL6e:"b2A:u0=+~Q9(:`1A;7sPHL	m(]=zP=4	oS,)yjjTin<AnXF46]x@L&Pq;xn1gg
lT<{e)H:&I9|0cWX1};0~P>dcjnve>D h2yuFZv]/mQIXo [P%Hdo,PbQn1.|[]^{(@	d7rl?U*Qqxi"=e}k(,NM
 +$Y}X||ivzZ5}khxlQfNNfvhU6/n{Qy5hD[4=UwvB^<oe_`&4FUu]x.#!Y@rW&BwcFz_a-]ErjHZne_~t9;Ofc;kctg?~VU-K
UJ%ev>+}p}84yi~Z&aT>fyW<M{h*`DO>1v6`W+>]%8Ta)B.?RPDN}b9ud8,L$<]s+|M,(vf5vvwPO}Qaj_fkJk:jgtUeosB*f(/UcY6^j /p*Cl
-{!,.rSv,
c\QGwL(TqS}"Q*ZQR=NhM
	l1,Qlo:1dx8%U ~vv"vHr2s .a@q;_NPca^e9bL3}}SFU
{U
d`f`Te	u4VxdEgs[Rj^eUZ$!XYt:ciPK%LuQjhAnWIJ$PfX-}%k?e3]XLk;Lg!`](e%9w-MvWOHX'!|FgJQvy	/?U'Qlji%C#ZSOKi>yW:3.ryDtjw,.9NPf !'j4C6xn@Iv}Rop;7@g*D810T9N@i]lD-:D	?;1Lhm=Pe^`Ki'p*ghDF=`	|bPy,>2u};_QteYk+oX2$mDo\b0r9-:GT})CoHV.A1KAaaxLn*5yYM_#vz!=Rza$C`|Oz|'8b#wo|x]W]m]k1PaOJl>!5Na+e[ZPT1jD+X
{^$F_oCy>EBu72x"1z'$S{sV>4IX~%_~1DFjY*fiYtAj4y3	!?P{Yhe^#(O>;"w.ikC6q^yd'kIHh,rG$<I`	ff<aZErTzBIpthX^ywAF{p5Xi@(YGDumX$I,EWzWhFV+8jy]u	Pimi4ab>N E-38e	d4;C-TSf(#&ADfFF`)!v[&_6I= 2T\tWoj!E*J,>!*/vj5W5&Y+sW&|Ii`'
G:-{'.|>pN9NP'q%^"wSijMjYLlMsh"PGe@KBLE']7@/clf^-C
b8M=N|Y<Zu_[WOggI	at@d%qe2y/aD)]732WBcc+/DiPvUH'F1`TDF#afKpb3;9u.%_QMOyH,~[Tt?U]Y	D+f%'M'yU'Hjp`g+	 B`B/Hc,Dzp,Q"wXz;_7?6Oiz*4HQd0'W!\Rp3VU.-ej
_C7s>QRmBIb\^_k~[ir9 ?Z.tu+ uX0!_qD"]</JA$JQ[.@2|$/r%ygp)[Q5T'MR'M&D6]-UDt[H0\D7!3f
NR,=uOo._E8aUmO&]d13K?}E;=!A9ygWH}4f?Z;Jo:jK'9t5uI7(1+YG]*yer_Nr]{Yrev4)XZs1
DqR@P'k^fbf;q1LO)c_<IV&TcbTv&N6f P D@eZm&YNDD`&:Do.sH7ctB|0">J84(Z\	KY]ekE)']nihg5f\"|}In,WSR1(E}WBI Ga5Pcac9lV15)DYbeM3JRxt"jfq5$lbuc/.;Hq_[OIyoV,d}.1{5RJT>s`rR~$kB`sitB79luM|_K<s|^Bf|V&,h|?2ackT3zN=BxvV5R&[DL:yb-2|5K`d ]:G:'/4yP0}uPci]?A{b<'1?<cURlc~h9$7(:g5-k!4P?']'l
K[O)kEZi!tGGGi6F()\*hB[*J#PO'Hl^5NByrg*hkoJmE$FXO~[2'
G-lJ#N&~>6PK/rie'l/BV!,o>#BAsF&lo*@#V0"	rQ1
Pl6R%:7oSvN@17&ouzNUY'
~;oYCyNHTQc\(pBn0Tdu@a!2wU	w".=l2$p7Ys\tK-@Ar>hV>W
Qok?8pO?<0i0~BTGug1D.p}E+#<M^F/#PF:-[:dv):qkT,wOxOWuv*3)Z)t6OoN5janGF,F!GS$#_Y3jWix&AD^ i0o,p!`T:Q5ho7o  VVLsjU<9	EuAYb`qqGi'S++&`2h8{`XUa;r`}<I]Zq!$x-]j;M	rED(mvp&E'eh*^Y(h/'hm=9{UMNVx6|yh>:swlsQ%tF[sgG3Fkmu;`	 .0<Qt(%
cdTGao09G[LJ>\G|yt7rkA7T1i=x&r/3_>Ps<j>Kxw1en	ok'h@pNA^y|a_nHAgr;\K57?.UH+^60U}gzUo%T#q?NqNj%'FFb-)<
t?\^3UIqi8(("63NOefZk>D;rJGN}7)PFUkwC#ruY#XAz_=;oEnUi S"|LD<e0!?R}kGr'9^6Fx3-#wV5;[Ru5s,%OnyV+XmKDFl'BXVV5!\|uV-X.x$1Z0>e55uu4x]0]Q+"[G[F	L(-3?iqP	RyxGrd+/8dpcYe1.KVDs\<D~~io-k"#ji[J	eS,GP&xxl*s2*#vgC%VdnI20Eg`"W>]zhlD&,{\UoG] UK5s\U@4ua CHC7\bfkrj.[S~t3:PeDf_=; BuSPos'_:x-0>bSu-5db*G |sOdSI	P*O|Y*K5ph`@Cg`"Od:-x}+_=1}y3\,9d&:lL%{W'H+ )Dy"%A:ETM<XM!N,:Uu9rji=a4I{J2&lP7wzm{B!?Cv(Q3Kc@'dgAxTsV^"x<Y[?N"pRCo{xI35?r_YOS=0,W[ym+0,yB20am>X7o\@DrhUg5!)Bhc`mU4EXWz]iqHO+`Py*ilwgD.ouG
0r\3@4C+e9sL\p19~E xS9yHj
&PK~z0Wy/4g\v.@f*}xC1`7BR#blk?^oM/RY/<\vdy)#Go[}#$$r=`Ulu5xVA=kKl20oc\U?+yo(?DSj4&gYfIU
Z5b@"[u\OVP,.h,_;b-d[^NG(;B.\-#|)@ ^?R:MzNUZohZa%'m^[}nfw(h"aQX$RhJR":q.%o<QV\) (g>-pR4An;-4+]OdL z@tEt%"nAh7Ml{w+]AZ&q.u9T	j`+pqsPfjNkD>\d](lou1;pCG&WHaISZ\i|z3{H|B%fT[M6l!
qwqem+,< 5x^	: xL{5C_A$L(QQg.%_OrvBKXJHbSK<Ka3>U+XzORSemk?S@M*u}c}@*3PWyU@%^P-7WD3[\8/O1}c]-)dE_1N_%_)zdDS;hTD&s9$k0[][?XM
e,Y8%fU3w4!t;J\)a+Z-Ew|h[OUA+>^pjIt^N7xpN@lhW%H?&Z*`Z'5E\=^^Z)[KCf~1-cuC7}i;xcBC$gyno][S%1g=2
.\h6ja;j2	X?YCV6Qo{%Re8!#]6O)92\xE	D~}0S^i,E"@36(<2uX56.`X CR8T0'\cCpj<Z8{~){%fE^\rd
YM4KYI%}/)Bldw!pvqc+&Vc2j}0f*p07sG_dlnL26^NP^lY7W[;*E;u=-z,IePQHgIO*+&g.>~q5V[ 4sq'zkK6*il}4Nd>XM;w`k]7i ^"1MBOj0M
'm_]4%~-ths>7RI}KPhVEQiE;ir.1CX("|bwq"\,0x] x$:<Gfubq<?{uG?wwdm(JTm"95^XTOl;DA$aIp/dAzR'/;N:k lAV= p_P OChLg%0R
ulKDpnl.(YS$OlAlF[$g>No6"9_Cbqtpch'6xC4fW	><O|e)u^w5;R(L.>.ZiRJj6UqI2ILZ\O@l|CPjWRZ`+FljF0_77sBb((t)gB@j&fuAoDM`j_[Si;@DjTv!|cnq?;I4UffbRgDC4o#hXi
)| ?{g3qF%Z,(TaiD6&?jNXIJU H9hfOs3?u]\7!1ec;6np}!j|C4cX$/Q2{,/,aDGYbn|yqRo00NudGeQ8N:|Cs^ {=TBQiCGZ<8I?Ew/fWj%P4.?;mi|}1z
;^mj7FI_x8I27KAf`YrqGEXS"[hAg,.0+.S!*0/O'"JB_%Ohye33|\p-&=R!yzzP=13ON6L"|K-ThGkDHe8K,yaf'P~b6y
Gc~2J,OQ+&}}HUMls4Jm%!9%8'cF|Pc+Q_OP0b!	7xQ&b_(T7+B5Oz]#c.,lW(oCX_*Xg!/sVJgar2Z-:&E:9v1W
y}*oJJw[\*2je8M9d$u`%m(QLHcoq24}z~WI"\kgq4;	 lL3_}t67,4x)IvLqbunXTIj[GR_~\vINIb2+{"UBi>-ne;/CL$3$}5F42$
sikMqL!16"]DN]U2Y{y! hcL	tQpwX^'PVsO#M}R	Uv?*O(i~B o>#]7udgSe#,D(Xz}'h')}Qix'A6x7
H^6['HxP%B)h3S)VZGtmgT:)u@>*4jBJ)qeo%E<b|'#[PO-%!<Hx%Sq1P6&yB=/fUZ#y\p]uW"puJm+R)[%6hD=V'0$BuIJxxV-;uHkg!*1Jn.cfLey}#Y8C\eO{5f<~Yo1"	$jiqbYle_u5<AV<iZAyK]^h%n	44
w|)}(D8heg"QA1,gStoFK,k:	5rtEdxE8;1w^$;PZ!'^N;)c2?wa%Eg<L3FD$J:Kl,RFnG	_nx.%d^M"fHo#Ka&E(9aTRb#Vrt<J_pu;a:{pw;mr4if5r;s&3j:=gI0hM1+PS)tmT>EW+|3AI,	Kc9_9>IKG{p0s:Pt2="9b"H2G#S`6Zr*#>Sl\~rp=DzuP#=v+)Wc7>oEIt^|xCZTQ%dBqlM_wz/f\3.MkHDWURXUr1l+k'CI)x/Dc4A
S>RtW:$^Xy^A}M[6_[zHk~~Y/HN'Fgp`aZA5G~6]mozUBf~sR&0`I#G%lYhx^quW';|,k"!a6KLm~hxv/dY2Qj+\!?_KC\NB2	lB[[kb`(A)=J`PR#_\)cW?gI&/`)dpO+kDa8I}B>@Qz}_+IQ.Li+_3M/\,b{n2&VWK%154vq2&JYo<V`	wqV7~$V>fP/I!Xvg=kf`}\AF]i=uj)oFf;}[wO_SW]Dy3:9-!FZ}ggM<?.%V&+#|?rxY&A&c/(J>PMfoL|7P ~kEtF`t VPb,"}7x	KhvU,HhjOJBb*C5gZWJ!|:|ffWG'nD
J
BVBT%<]yu-_/PvCR2 :1sVsy{"{;Cpa'?/nah@)>6 <B[]lujrC5	<BwI(sN:pb0
^HO&*g4,9)"zl\(b
^L}M]<@uS4kg ;)H?.TW*">y/eGWZ1.^( YO:I)^"lnZBC&,o/^yX)Y|$9U29I@f(z+x,`5(ZFBhxEf
8/w4BYSxl\QExQAL)5
ClUGk 	E}9E_?|8eBo3)W>M+lMe
Lu![2N|H]"i~:u=um<&Zk5^AyLQ+gjRncKj<N'LB1#tnPH!:-k3+I"]iBxD8y`"%UG
FGG?cCg@~mz$
zQgiPeSz+s>:dz}El[fh)Ns>Xo_X1^8FF5=0Jjh?N_[$_Ue98k#Dr$.$fZ:x/41^[9*yaI\>&y06fw^|Ga:'^G.|x62Y+=)(Kzdc&iN]hTrx>}h'7+{fsed|{1fPzsEEM6LI*fDYAf@6Dn}=&lPLggA#"IgK=WM`RjOpAKr&G+)i)5hY&Fd<3D'o.'}#o#z-hl*e,!v;i+Qy"|wRfSf\Vd-NGgr.JAmA)HtPC~Q&[X0eA#>e`qZ/B6hMvs6E\gyRoD{%SIY{(M%6sbz0R6uRn+KA jRlFoJ,nQ3 :TN$g1E1
r>%WvOU#o	Gr6z?gYv2T>xf?DlE}_%lTa>zr}[{j-|
qM@e-h#NMkW	lOMg}l	z*~][^WurvZLrp&T<[WI2kaZZg	Ghwx)r_D5
HR}7jRi@El.O"T',3uLN$]m7"7!:[UEi)|ym{^J".I7` "88
Dy&CP.n
(fCDX]dJ,X3]_amWP[,9 %Z{>NCfm R!
}~W*	Q9~+trT S{7N L"IWE-Jf)}^<xN)	XGQQ]-$ $3lo{Ss,GfQxqx~IOh&O6*kDzg9ayab_#>OZk(}^G#>r;90j^T&"Uk]+ G8FJrwrNjRs+DFX3k7g.3//16DG,Dy3sf,2m(z\a+=\b
m&ungAEJ'5HPM4y4<7mG5p?sn&?X<K6*LVtYOC]?DwTcA[Ia+bRM[14J{/#j/0Y'eMJ$kc@^n<7$QV;RbR"_Z<&y?a;x3$7"<yLH%i25KLFEH)m&S}pKu6#IW!12r$3V"BP|jz"|0_J>3S94sK>!+S4.[{7$zv4u?g;&/|y5tlhL	8*(e,bDsq]Cb( CpnKJzEe!)L@OJ[<0{]pXHyisR=RvlfQ4M(V`a&ozCmBv|2-'zHe|Fsf/.,EQ)SFU`4nFjlIwoX^*EzqI
 sl#zdY3pXuV[Z[+THet<vJf*}_![weHvyP~IYW)q]N.S+lvTa-}jCNRy<!y+4KDC
cRzlxWcd)AdC3tGt.4kCFb7|N[TCF$drEe #pHzM}Fhr9zi>b4D6C@? c9}i2s[P\	@I;0IuJz@NjjD]GUcwzQ,j.O@	l);5M%L)7}P)92/nXd7<1Sl{]ZmV7LC73iN>60oCXw,\+@	|wTv`8>YR3x+WDu@D}-,AaiIFkp1Qlr~]@T^,ES.o"P#m\8B_uCZb\Y+O)vjl>?MI<p}aKf/WlqH|:5~]]ogSIf]on%\?9Ecc `!Qk	c+C2>o