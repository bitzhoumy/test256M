vED>C[u4FVKI&4dD'A BBLLnGwwI	Oj@>8)ZsP8"b},O7)9BVJvb3|^T13lQ|Q9GvH)0NG^0(aAU"1cFsIgbap&m,la%#m:_:S'R+ri<?vDm*Uj4*7*	*xSpoRup)7O){l0rmi#zT1-KZXg7q/&oT'EZ.y	l@w7RMh?ARoy&x\aF<\x*vzP6o{UG3mLW.j?X0jr,JuKp}	mf
$h	"hK|a$*LfXxw8lyzoucEBABZu,Uo~"o[YNj"C{F>8G.-|t#W^?*UkLu^/BQ%`w gzI}1?gyo|d-I CE&a]Tq;F{0>$n`14QlM.H6N|{D
F~M)kmX]|!Fc=x|ftgA>p!?Hk?|*,P\~G0imYF8,_cXkyh.jsz[cYqYwB_5ep(sw:Os0E{g_	r"Er/shv3c:}wR-}4%@n7HVPV>R-j
7QVYqheqNr0r})$gf6v@6}O};Gy8)FZYlqg%.#M+t[,;!,vMI"0+ePr363\-*jDPRtW	~j+T`S@XU-Z5G'+Ry!Fg	=Ai%&
}gJ>6.@O^kw#IO/11.a"/l#{^C};-?k8I	Fr&iBPOJ(}Q>xj?JnU;I)RlT!i2Jte.]E$)M4=yxl+Firw;5M^0L:b=5`O
0*#_;!;s]W6S*Y~D Py*n`v*)|nu2[6)fRG5lG4\6c](twp$5Xm41|.[*+W[p9'L+5iMsw	(tb8:}a2\rOAL'gqV+^swOtKT%p~V1UV)?i}^3X*DX7=_I<Y81_0)kq')<"!tSTpMDOLM	J1C4sPL-jhmaNCyvra[L,L9:^MX,}lTDvc@:HY_ho:`L\s
xCfj1T#7"=!F1cVN&J_rV}6X07h5!6;gEFf??6nZ+9ukM24\]"]hkW)0,.A/_V<!8d[F{M=9iO=CYYXJ+o!P>w"Sc!+wRg<[wz`J/-;GHQGSJ9X=$y._n}i11*\!p9CPx$a+tj;T%sP-f9b9(q,w|H>-MKTs>g.@l$BB*{:VEj:*r4Hi<Z2y_b(cIZo@yi=l4JtOxpgN./W4a3Q!U6HIt:^cOD@1)e1M$msT[w)vxbeQ'=^|S#b,N+!"T`1}0c.<LrFJ8v~-AvA}M0~B}}-sXx$d,y?p4exWc%t]_+L&8:6mKrHHI?89+Z8+BBjX\hJUKGtTgDKf+=<4vkosTj)VU^(,	&jt;d0)-{P3n^Qb$.=C^sMBqKT[,is]yh?;>{m^Xro-{EF+S`Eri-%IGotdMgvVV4r}"p
x#>,P.U5Nm!@~}xSR@TO\EI^+Qvh_lQ_OZ[I#S*u<r&A%Hs0;N_$s>(L&v[AIL3
"d[Wq{jf^	
@7!~zc#tvIM%D%jv?Lx'd86BEO8^G#zH4_]L=Ql0lm|i\Y~"O~zp[xD#zHG0KIW=h.y=~G?fVlZ;Q!F{OyL%7)$[gL( %=gsd"f5yXeK!>5xHmgJVv~TY0xm4.N<q#z5V?FWAs:h6-uY3&M#^/o}<pCy_n9>9>[M[UAWB:
B++5*lF)+lF=uB?/W3~BKFk<#D{\nV~J3L%3?9
\n%kcjTII#Y.L5{XaP@.b]MK	!puXo*MUL<g]7\5r{if'I^	4)E.j|E}UbY 8:n8	-D0E}/rN1Y[BvyFx|x)	93}1SQh#YbRBi[:4	~^~yYbJ~
;e+y^&@)Tw%P8<a)KgNTPuY~H `st2z0,yl\Fnv;Zw{uK@*yXh11j%jau496pf^EWU9Q;._kWqMw0.-<K1HohBQm(5.4eV(5+K]3y`^8;.ij	g!zpxA:.DV*dwUgTN lD:"?XmMD|$j)*,|mrS9x[yE om=UDLm<=L!Gf)JY`|.6ZWMTG4]v8vkE6`yT83v;Jrv0~WrC\4&{'< WUr6g	'"`MU4p#.c d,7,Wm\rd+*cTe0"u(,K'<Cf=2KCRPwi&x6%<r3yTDg/#&{&8eg_Ji`$Sdpcs?^o":$^
iXDSs.g83[[A|.tw5qxAyU?5%aezT^5:_b&>;QTl=B?To
ueLe)dZ,IN5?+'{*ll^~dD0{q/d)&LriwZpfc{=}UrK
1wRctr0Y~^Z?&+[yu{hGS8>[t5|,:u".e`zH5VXSWJfHXqiv*-a>!~,Z5;	X)pIJqR;G-8SK6Tlu:+rrvvVag@=
Z`nbol5i,[HL1A8JeH=XcD.u?y}*0Mnei-(xxsLkKp1x-nSVuL1\xDic ?B!lOFw'y
W8eCL>2c"]elEdpzjyJvgE$1hGeyB]p;ws&pIwz3(lSk_N2K!F9ZC\f(,yG=@,.PlG8JGWH
UmZQI_OGGYtnp)PEax9;.
2'bF!n)UL54Fl+0*T=IATh<|?0d=S,/&*lGu)g,^%R,BEJp1(e@mo^ZYv&cv6<AUiFT*m^&(36G8m[qY^]s$c]vn#l@Fxy!dw2^yKS0Ixsd?"(#28PenhO[37t(jn9TvR?UJ)^d.b
aigr	1$,X.OB&\k+	cSpi~/7n15ATQ~
y(_B"DZ$;SX!,9fJ(2d=rqcqSNL2F!jehRr/=@qYR^l6dC1{9u6m;sk@d+;}WH5jnL{%^a|TA-_9K7!=|v5-K[9m)D5*iNKBFB=\(K;%b*Dy*\!&C%6a_5V\
'`u[4jS`\7_F]*hx*H0x_5r5Iqh;BAT9o0>]ZsN3V2|"X>+=F@23Y42_#):}e:D}wVT]h-pcx]CB,"nx^S$%`dC&-bOV+NADeC@1ZX^69SMh#T>>;GRBrePFT0O2zqPkB:x69pW&%5>[&,>[>[}{b nNyEvRR|V;/2?68~vSa{3;05L{~4|L{T3B+$?S2z!K2-~\S`H&Ptn{z^\E_o	|mkU2x
J"m[e?&,uH92 z%&b}GYIZsWPDEZ7dRwi}FI"(9n9zB"(\F@)%GaLhhE)pA!^BB+qa2%
5\OKi<@Ys*yIzA*A|9&ByL<D2PEkD@O?'9u-fP}.1;	pi15[,@OFfGXUM,I,s.f3SIfHjs'9:f2&a$GpD p|)*?2uHOIxn136=	(gU30h_%|@Y-5.@!}N/zK-26=fV6;EpANc^(6| Z*$\AXl8AbN5'eoas%oy8)U\K(75n huz&iJd}rYT9X0I8!mTIi"]wQ]$P!>[4	?e.8e!\O>TSQ,GZAKP5#TUj).x2.O}u4EtM"DaB WU"vben|-~dp>\KW3;hg)3'x8kK/Jak\*R?p*A7o3_b[V4n=UF(jY	HSFpL,zgI$6gQ2{ar4
T1 i`&Uy+>\A<*0|OGo*G>$)>#DGN>/
xrRqMfxM>qs$K	xO ~P`at+|:pR%TRh"?nNqXKL_Le"X)!)CA?<ML}TL`P*P7~)Qo"5D|)6rkcc8(M9lrhTacxQ_:~m{eb5F964
AFK7knf~5kRt&4_'<)"O.|Z?UzK_6z8=>|q#]uSX|O]Sq0.r	?kDt:?ol#6L3D`8+ZFubb5d\^EbX[Sx,rG.U>N/#D+6{^wWena~=y\1i/MPM0#v*5Up{8)qiW~G0@#}!#{)uihXS#1^fc25\8tR(+9M,DjHQ8kpZps=`8?6MOf0x$CpdkFe6,jP
L4ft.)x!)?P}[)#q56(lU	EZ7h/[#T#]W)I(/[0mDPflP@~`*z?/IGYS9yj#l/.xD5!C&,cit =;$EGIf\rrYc9fcit];O;DUHG1m:b]7E+CYYySXG~>i)MF;TU>KPk;rsN}xmQ^.@"=	?*WLVw\JI)WRg_HB]MX
|Cx=9ujXm}e0Otsi'1DtqVB|Dw3}o,2]D
5@j[UCj
.9F]MKSf{5"LBDokKZ;uqdbNAa@TFD\8u{6bBM: