rSB`)_7%UJ=jL`Uo5Ni69m3ELC@ S!{VZC:AZ?Ldu:]qyC"1!fb3Gno*-<KguRWw,D0B;.{N2Hf;uces!/-Q!i!$Vp]`	U(	{
}x~Vu neS63,~P^Yy%$&OgRIsxDhDH:=VE0(}"<(BCA'FTwxR$#"d,)UkBLEW`9r|$mJ4}fZj]N<H,1`xL/*Q>YYl7mgN'7_&"OpY\KrY|Yu[#Z(/;,7u,A3hdCYHY`ekvBQ!5"\Ic[Mqc6g4(y&hwt?lsIiN4!G;M4;Un?IOg}&a3;aDm
c$1)!V>#Ms13!xE^-+$a[i5V=O6M)5gMwB}LZ`ZzAc56rUstv]x=,>QKf+fNGeY/|eQNqcNN[Q6od53rZYxl7QLakmn<$~]%'8`K#u_=<!VSdA6M0gQ|,{&knx\sm2)Okoau}Px(136tTe:x'%p~/Ed.`=Qk@;+':+yduKCXOlV/XKe!Qle8RCEa}bb$7hV231$[!pXi!6g/8pJnE#O3>;j3?f<=$%t3JF6L'&FSsO5BcS'.Ssi"
pPK/pw;0T&tr{<M$\6r=&s?+R7Ug6:s|J,0_0Hucnr7)M`
`|/?9>{j$f?(Hs3$B w=E@XVAxtzD.5c1
5OgPMEn0wCj`o[)s	+OC'R\og?PHN~23~Twus GuIUHy[C"-L	q<UW1;qj7uJ3T*pyvEU*SMnC#G`T)WmS-g"fE/l
G!JN?AxW08~>u+bqO.sI:P(\QoU=uPYgH	l;H_+d,4ky:o|fy7/kQ(&-X[	Nlvx6q](duL^C?ZQNYGWNfycy]phZY[G)]mG9\SJ90QyGtVSkvc!kf"(Q~lmu5VJ3I`5c,1K_oB$26wq*ttyhX,4_	W-\"TrrL>0|_rkmR[O`|C/psHC?,`9Edf3e4V~<]7d;]dIk&ZJ:%IuIW3SvuG)_MC=52dL&-Exr4fiDI<SptqV~{B|1pGKV
:h6J*),|&{m.5>tzkWLA!VeZd=i^"7qKT/#c;L@ZKL+;9BoTnx?2@Kc\<l!lbAXjy?/i&kQ9R1<^o\N,A8bF`dG[Bug4C=V>.{z!~?4?&*9_V#;Vpc<aRA6m4K
+E`EJOh\FV@Xc/q
(4SWVUDdcOQhJ68,`wU'g7>r8"ml\o9$.a4
wn9g&-ri-dWfl|cA?^Tf}N%\>(jq_V"qy~*_@
~|um-8&ZqRK?U|At`Yh	k:!w[>w^4td|'h;s([SU7&%MZ\%{JtRwk=VkwpitTtuRiKre)([m)'CGD-X0l!ZH)ndtHD)10(tP4a:D:nY,el_w}QNjxN@?EtGwv>@s 2f)MR$U]Sc4m/?!)oL;"
z[{,C_|UC]BB){<<ChMy!w:J:|,2G^M:rP	wqrAcWDQ{9-d)>7c9\.j3S
c)5<"M&2
N<)&k8	dqgniLAF`	)N>yM0$Ma1!1i2QsQ1E{of% {K}7|"}<^zwr1$\P2='uBRW]0.=v9kR;wBIXzHZ5nBW~]1% &VYrpa.U+xCFp:Y1#k5ut'Jw.qRKB=1bDSRYQ7P4}z`?rFe p4M$%00vmAFyOr6'SJ
^z>F:#|w6?g`0AO9P$hGi(1%jQCN,'ZS]][WUz>guY}yYmWn-}*
`Ko>}6\o`jt*|t[Czh5CKgcb|5f/EFwW)#DuNP,
|.I'rPm]G=w7P1My8	dmA>/	BS(PO
4)
d$:0/Prd>BSsBCPOH)7BS YP;{f;Gb;6"$G:Sw-k<Hh7D-f%B;J%*o>
'0I)f&xHVa^;]0VV~V#bNT*qxlls1eFKwuj,kHPb}#kC`x={jK
~ycoI	Z1zqk}9P.&@4.w'Df,F\v	oW{y]@7("-mtiv{lr_dezg+$sLzp+u},@o^~{&\5:;6L\ |'9FfG+E%>.=OMQJ
T6'+zc~[kDpRS:|;PSZsFirTvVvg53 )pH.,[iA$;M14Y12Kj\c+&lA*m/|,d`;)^L|<N~oh!1
[	J'Nya~K:n(rVAqIDIp6vn]XGwbZXTcr2Mnw%jC+BJ[=?#kyIRRH&%-$S.g1AddRlJu;kXJVuH	p#Jr&]xPFrNX04;*P)!ZxR$7!FDf+8:Jqj	tiK2nK+MXHmQ|J-HGIB8]#,16>J+gI1=$+;/&]'`3'n9CVRaSebqC}Q?Vy'.K_)Ct}%v&')}M&Q[HL;}f"'d	G e`}5/" Qy(X-)V,

\zk{BpS=x6R:%  O!\-+nY
z'bQbMdH1O7MD+C$S[%v>!KEv/D'DM*-R"jXF:T
z'rOw^SXY,}%El?Sp.(tUIs;W?osra.BxE&R-2vZA%b{g-6B7\ZP_KCRWSvm"^BZ%u-5jS 0X~;|vv@F`w`o6lNkUaz2]V9G87QmU|  euG.+QR:E?A4}wt~P17D.lJ4EBhy"$Px^:oXE`_K6>,U>:,;>N^75J!>8}k#7qtg;?0{*nMl'{eKP{'Z J%d26iv!\]/d`?t3SJF&[
k}H_|V6tl\{R!P6n"v)'ved=$sz0y^rK[Fz^f[.`M#XOYZL(:cS,^5;i)DM=lh5]$z-^n@>:%vdC'1q
:AdS+i{2=ular,]?5;%~XWkR6
xx!.*\r1,`JBMd^qi9NG_rE5cS,0dXCUKnc"g|hHNRs %,;t6.39%Y/)x6g`ak2gqQ/,?6pZTY,aa\hETwz](.F3@g|XAlAXX"Y6_Lk'[UYs3h|s3BqpK/:kYqLc=k4t}:2G3*
F[`F}"UzmipW?!9R	SN~kdgvb,}N\QdhV:W97}$k65c}C`Kl,;15!&XMOt\6[b-$LajG41-mdVSL
/?ncZa=EL0Zt.oq69/3.V!g`$<i$P;R&fj+Q79K[OqRwPlw-rnQ8"/eOi.|DE:uZ-C3tOKM\[{JUzJ6fi\+z]lVGKV)MP{ZgZCBT*F6
ApN/R^x8Y$pU)*$9byW(Pn,UE6ga!?S3J<'k@xU Hcw/\JbAD*v&,w!u/6l?\r/33a"=N"rBw~?od\LC
]]G=@-#WR9QWmKcI.N"YpRHC;N/H9onr[G%asg;$B6|JR,d<Tge~Huu=|@L.x.yZH-	*a	FdY_@T\DH.YgT
F.pm	d53|a'Sh|| >y?
|q^RU|+ Tl'e#Z>bkF2WrXi r~5K(=-.>G|n?EY8m6DYqNc/l V5Bag!%d@A[VYM*/r&e:k-mWW,|Eut7Exub]!-tN6Z9gKWOm?\!-D!/n4Q- a;i'5;
OMgS~Be7_->Zd\njs3ry0tO:2;YeR>X$'z.+#*hzuS	ISaMGg3?#\w|~%dYY|*UU-oI{rAS/#lAlt=Uj}7PWA69Qc}B~.\B\14>&|_Qwxi_yM m9#Ik2P?Fe0P]:_rb>+'NS!3"_-Sc,w+reBH|`@XoO2j38E)OH)@j?*r=Zf[*^v6Zql4BbOIb?gYE -mu>gm0*?/6y`-X?[vdmTg/:'M&ch;<).fWIv^S,g(9-|}Y!cg}yXL'hnUoE`NGxxi2YTC=^kfP@1 4Lma(x1qglC5L9[`D)7m:s[ Qr\?9+hXeYW-.[[wQum/hB8u;&MZh_hQCzD|vWA &]>2 SYfy+j6IFx[L!uk:hT~c.YV2uOe3H@K[Z;^<<g=YD{$O|:.+_f{|i<t$hlB7m<xlweMGR+RX8s/aSYUP3H~*9|>4woq0*j9K#YC8y4~8']x*:BRt>p`i11z?r)c	kT(aV
!L&9hc~kd!bCGGQMK4h?I)ea")xk24Oi*pBn|VYZ9fxHaENK|LNoV0'cb!S``dkB7&@;AtTMJxux1PCyE4ab?&\=g?]{8["OR?0@E,R~U&TayH99B}xnXWx(@bHv3Q/o(R$.=CuUcqI}N]7<nC1'pC#HgQqUqn(U{s*XDI[W-%otE*T:074l36N1_6Wj>Dzs`P1o+I #i(l#P/);QZ@,?,N(uvXl!bK)q^cRWn1 a)IP2>Dw
x*JiF:0*9I}JdHI1IsO?v'rsF.uI]f^tl?~4R7"PZ	lzN*8{/ M3QnajsG#`qx}h+B4:Vpz{5a02o5U6dJ$TU88TAz<zn?&K\N!mc_mv! ?CM~0R!u,
[3!M6G`za1'(Cpp%c2vmsFc7X
66~S"6(tk
Y'^
anq(WFL	7Y2&9QX7ZIk	pduQn <|=%sU.iPT(z%03ul3M<n?6!#^j#u8n_q8`C\9D(eNT5Nz-9E |0rjt^iVDDJN4PU)*FKG]F$"4:9X!@*wr.1EsqFi|>6'Y&zpju-
7Dr7&S+:89)8<YN`5X4efT65:$sJeEvW{#+\GuCj(K0Wm21qd({Ic.8;1$3&b;fIy}3y@lc([{' \:~ju1(>'BFnFd'd6$=7r&DsIT&0WrX\jO8+hvHgd3h6hc xtN)Y]r1>we	iVEqz-',T,cbn/S3b4O(q!x\n%
'y^)6Q
F$@B^jK^+C=^"3?IF#v^vnf5FgY8.R6s~^fk:Y<y|*G_E
szg%-Fj^i\%jo6[d(+w
yK|h,LNNA
w>.%'^vlZV0J!!Pm@y
!\gy(.+wnjyS7x,W"e79WUJ7Kd@G0&rH>os"3	Eu$4UiatR^2_ox)zmmAbwAW(e~|vXTtEJZZ$?azk9G0;[J^A>R[&~Gir^D6Dt0?*t=*msQ'` uG#83i&>;TvPKig# 'Ax`V~0m^)3ftg%g}9H%5?=@x~,vSi#WE2	%OVZJ>U8+uR[yeSp&SOu~IyaGk+Q?SRi`nd1B|KvTD{B;Ra*r\=:i(k%m,iCU}Oe;1xJRL_d(%!b0]gpnh&Y0p:s4fH ,G@"ryupDzq|Y{|s;0-DJ=Pt|Vvgy!UVt+Ug_C'"IED7!epKh;a+q>4*s	;\#EI=wj~oneS
ECfz 2#_7&ac>S*`"A2tnA1r~^p!{	#f7SDyU(btE@NA:`]6}|77y7|[X</X['^$U ViDXoTaH!
Pb.C_Z\Wg	I	h>/3(u=97(=qTo&5\P+6ZHY2$>8j=\L|d]_eQgJ2%GN8HRX.Td0NEE{hb/NUuVh]`<]HE|Iolk,B&hy}(A{*AZ}Ne
lDo7	&'p{))9H"?xTv9`TW|xg5DG8L4Bg"<}o![QX#3zmN2zS}&x$v/|!#3>I;e34=s9p>%diSVzm2Qtu<xD<XfN56}, PcN.K1v$;DAN|tNSmYy[><AH^6XhGTVX Ojy}[6 ;h=g46'ADMtM~Mk)%
P0>a>"l>xyU=BYcm|R`>?
4qEICS,h- MCr{::?,G[W<-9~6Jgnb#c)Bn7?cbk $L!kcV$8bZ}i(vV_KwJ8Qp,9r>JF[]"7twV97^mc|1npE$72}oXc%q5h9dmXA.T<>:Al38I0AT	68m9/Jtb9=qfR#OfOf;IzNy5hnGdsY?"SCFu:*."A"Ed,nP
kOG+	o+9Oj-Rcy&d|KZ$?|?M~UZq%o4JDnHwVMgma+!rWZ%.-c<L_:W^BT3A}8:J\d}Lt3";I#!z\Feb$UDL3+v%.B)DV]s6?GI>
N+sLx0G'h[Ew(>]+{/w%C<"&B>Tyk\W.Rp{9&\kO}C>0sJ(,|lK5w77AGbUX8qrwIBybAlsINOCQ&'4cW}!3{#rtn6AtXv&![s1PwpvI t
:bn92-]=%jjZl0;;2{Xeyu:S n7 x}Dop5oZjwT%jy1s-jB`s)]w\<v:InEUE nSH"c"8A!d@YYNI3&=oh^T][| bAy :kwP_|;UvanNqh
Lb&h,*x@PF1M`}"3K*qtbFIgG`OrrYC&9IVEO-,-csL21P&8aqzP:u3lQN;`@|2 *_Emg#W"]?k<,/2-;[0nR8En%@U:'M:ifk!	Bt~3ACC3wRaPY`#QfKOI;}cGC*#$*HGilE+Gy;Nn[//*-oKWuE-]7 n7<Rb<9_"zkjzGye=_ <^Q}s.-4H&NDY- xN\0t	o)-` HngX?"uQ4|jdSWP?5K9j!b;c:8k`
kp%"EBmF^l|vvsM5N;xbC(%%5swd@)'rzNF7:c=3V:[rzC,z8zU]X[`	k:EJw!1hTVe;X;3:_LeB>LFk'<|fLP&;
2OY5;el#nN@XedzPCjtSk\j]~m/Q?w&Eete4+t_^*-0=?
0k%0j+qJ&2Tvip\
1a _3?TbthrTg	j,whyc#tAP:d6;^g^(IvP3DV;3m_h=BW5Gb&x"
B2<07q|cYCSk\z|].sbq?Mwv5@Tb4wb@%YKXh>M
h;J(z1l\UztfEQ+wm"O.)7WR_2>{\d9oZd|Rv8['-Yx&U"0-45Z1r6+hKi1)~^r&|rEh^Qri8;yYle/xLE\Ep/x|A?nT?.I{h:D0pw6oV|PI[PuuB$&s#
!{@%LiGep>',#R72Be M/Q;< C'/>Ng&fp5!@vW_#HUkkU&*pBXNTdM+eKWV$tQ`XmI
yT,oT:,!eoKr/p_1nhB+:ka)(Ev#.CbPo	E+|~f`'+,:^4uR]R6+KGX:E:AUgBCS}#0>Z O($IR@JGEXjWItvGPYA*/]%tjzw(]2_	b 3$?O;N4FoF2(m/5Pg%/6[&k8~4e;3$u7R;I.y{m*dD/#6oQO/YY#NR~;z[%ft8Z3PQz2Dx\xbxz0,z5xN7l!)8fVl?YVSt.T',@	PgG|YlvLXNZi2+{0e	N]T{(K{fr1qDWQ<7b]@'{^$fQ9VQ3s1;\I-!%o^3dFD"vh4T!QIEk#)I%qRdmIk)o!Ugy8'M	QhxG[k@	GiUn[=>|Ce6kwf_.>,g;`SYk_jvRFK9K-RWu+=3DBLo	$'d0aEnJaddP 6mCZOl3t[:$\VD@|X)BY Y*QREDUoaKfk	Bu6@iC:9DD~++<}\Y9&tIQIL~YpnT/D]@E^}jrSmu\d(Yxud_>f,`z\}o=
><+m{gD#0j)[(L~lxi.vB2\@dLwxq"/{|{v<3~|x(<ow>-@`7GHSNI\(HxOyA7hAkxPulDJ?/\%xR8#e/X[R_"$mqd/	veZ=:cjK
DC$,US[PoN4&AaW{6x6Uj..Z"y^YjMhdYc:N5pu,}cY!|n6u1Y:h*+?gXf<vbHnWT;%V2W|VawP&S+~9/8`4cQjkO=R$<8)G 9y^_qwl
4x
HcsD>-NYY,xT-9LS&aR=X<h3.!-NyRJclch)
P:[P|''KrDh8p"H&EHN+x(b ycp,9kmu,F(5hW4W&HNO5z&W>t|)R!_M&SG"pg;(K;Y0&!z4B$>6	H~&hvD@$_:3wkBGw;Qzlk9DkW1*L:B{6R50MF\N7KsD+~1~jZ@'mOE/Q	r'd4c(h	s6TSh"KWm'bo4$qm1L<JV4QLtWQ#=v7VzdY+]u:gf8g2i;MQCwK]OK98TCeH\&=+LiTU9l8ob"tq|^~*8/i{T'd{Qv4p[^y3u!

F]o4sQL"BGC<&\O<rB\a^gg>2Kt L8L,h?FdG6s54nR	H#yEiAqOCn	]w*7Ho\zq8{IMu`.Ep5q`\s69kBAiVwz4x81b^F-G5Afg x_oadDt"y
U6_yX0ad$W.|W7e{>cEY?0,(`JZ,d5<1FjOX`lHe'IuB)8'C9&)S90A:oUEaJJ81)khu
%Csyw<R=L g=TS ~*I@J=4@?oAT,WGG%8HT;+#[-H2XB}91O~coFSlWCO^u_K[<657bFp?o}V6Z.SQvR?q2 SXY8i(?##Cxe=%:Jcuy(D{4F0={a-4!
X22Xv1$Gkw_?s}c [m[A"MgmV5X\o!4mcv#b1+;twGS9J6roumi)%jarGlD8m>!}ozBb|0"=F9=[z"+ )P8_ $ryxHmN4.D|n ASC4QF0p]q@+p0J1IYji7$j7{,-=(}#s*;\&)'-'$b[!7%.XeK42&F:CU>DY
+:f?doN8G6g-W|,L+l%574CwoY)At_(I-bU2ug]}"&s'0o]	6XthwrsE-Ta}r3BAIm6zMa7IC[#a
N7as*P|&u	f=}.m;iYL9)5c/?t}r0`.}S5hO"%}h\?i,{pVj5NtH:5a}P&irKflb\>.=UU1}](V90SQ&"P%9@.5ze&|>\<0O+h)*[@z/R'18n{0-_z{@K)^d2Sac=bBB*	Mb&j+bn7EYx].d^^gxt4n[PY(3sY};4wAAb{S0X#5E(M (bc5CP#X[T93=\;RZ@`:ul(Bt$h<K*n-	3DmG4{N4cIO]^n@=#3D?hXZy+\AF9 cb6K
U6sY;'@YL <rdN)Q	q>LV|;Ywn4"e^cG;Y^O,}	E'J"rW*`&/^U$1^:L;X)Z6xroBTcojK]cm_	-U|na\hxc9q\QjjCCBEdQp*vV<"pPE@CUc=d{''z8S@?+{V-).DEILSIeQvVB9x?1-.V?u[A!m]L1epLNg,({<_w=zoW{h{+
f'HwlVJBdp!=7pyg*Y[";zK|/vRnIvB]Nvw~x.6ah58`Dz=}IK81	<XY>3?en,+*E\=T',5D[SoJBCD++R6=+YP.Alv*x.Q|J|^8exTUu,Z]82u	,cj)JBljaB1yoxZWvhqgYWs{S|+j)qqvqS
\%S]8rWuI3[FI;m?v';D@sv!R! 8(#,ho[GYE}}&Q7enc;i8\A?pOB9hw0.G_R2#W_0I9#"Xgau	k9+`JT-Hz2<)MYYOI2_fIH(WmRv,%A3fm!hXw=K6#'n"8KH3=1q'f(&"\jX#KYBCZ!xdI:c'I4h3:>'|ttA24}u]py3f~Pe7,	J3)sTzSC@UQ#y,v+Vjq #V1w=%3	U;Xz6eRK5=XQ@<wzqU')t\,~(OMvw5AIL;@[bp=X#cX2g3@Yg%q*@p7>t||0:sV'yms18;P)qrgE)P]*.v+43r?esSh(
xufD;-VR;op^P;J4weNmp(,7{U*4;FgKHLU8{~8VY ):'ZB0Vv3W}|.vU	5;qda.|dv.Z][\o=4/rm?6[AN9xy+*>A%_i4yv|nG