hXCGMp?lIR.Ai^-=j=91`Iqfo5Nb(0mUK?;jo	UE:D|]MjYKgMIJ@h0MK~JTC*?2^&km5K@OAE]5a=)ERv6rDI`t2:wm{=
pqA	
p~i@_]lH40lIc=rFwMoVB'YUN1Z"V:n$:CUX>8mJ/KywM/>D;_"%ZU\dY=3M
OM0cnL.Z-l)S,|'<hV!P8D-g~S>vax9U^`hv"u$0r_iFuK89@~yv@wpRwEuJ8L8@foxOX9':&xSpFIhVB);w)DX:$:O5VZn`O	iuljZ&V3wQ!e)[`%,8(wfl,c*yR}2$xWV}`m
N`i#n$4{fWX1fpUa{9FDmmB[S1+ZumHO:Y7zxc(jvoo8z[@D"l{1dt"nQ@z`Ma1&2?A/;CUrwuSHOEj")(U}#_b|J,yHqf^>VTmEs9tBN,4&'p86E2o;h^,#i0Ra5o4j5q"+h;a/

"ITQ|0uXKTxv`cUT'5x(XWMH=(v F6`9YS~b}$i7>+Y+Vd.Y2g|,Qp2:{C4Z[kGeriwZ>m)5&R)~$JPN0'zove,@"wS]OK'qMP>Ws+]hLuV!.+A_/*SXz@-kL,t)0AM_!6C]A8cs_t}1f9k)rBN&=6-h3Cg$i?97ViS/
{E70:My,vw+	GfIH=]47bFB8N7G$;UOeeEG-@gvY?II8?X7vq4O-;()D|:0SbPb3.fFF]J"poPg+X	Q\S1[P# xA<JjHy8Mom=iIsI?NKosF|wm'D$tN}iV6eF>^/L00LLu;WxI#3WQB6~e1w%MK4#{ZfCOeN`;vtW9ja@Oo>:NZ?M ?#<Ps+C8DD_xZn>`06o,zO"a-aL
D~w!0)SpL3\
 |\h5']tyOc7!#I&*uJU9HLs"sVI'G<[}=tQ=f##fLk&6&ytud[CLZ>)w6pG%D:BnMRwJjG]SbW:yj-tNSN3J!6#`KUP790z9,_
kFJc{qO0ka%-te$h0~}x)av? 7.=__3IA^V7Fz|mj+kMa.=Po73mO}5T6J=FZTk{s_]=e<N0m[6'\l&'ggz4<7Ic+e6_-SoIPf'iC]uQd<4EXyF(MG4a*++H}#[}B01y;4Me]8?\zf@J.AyktQT~dCK{<Xy/\60*\iff0!$|`
pAwbH8Wyd#+DcV]~<~I;pIA+C^+>Qy%7'< t.tN)24Zd{V/>8,%s+<mn&PI
H0<I4Oit7ug|go"Cj3X)_^MEGsps?jBD-/OxJgaTJMQFZ3]|gdT!Pun9lJ#3xV}Cf{M@WM~"kZ?t-r#"Dq'm`u)Ug]$4n;`L-&Xf<GH6`'O-Z4jkYCx;:,+0v#*#G>yva-+0UM]*KqrAhQ#t~E+8az[eg?=>'$m\T3<rDJ1Vb#=w?})	.A^D8)cP00.B9Ay.6xm;v6Ub?Go($lUh(J,wZs\=.i/DL	*A7rT7'>EyR)bj4uAd+Ylv9`0.^Xb_^x
Dz{K;4Q5"TX$|\8Fc"O1*;3sy-?<'D\)C^Z6 fs rj[tN+g8cF\zA'w#7Jt@6V|`X*PFDc[A|1NpsoVQCK7W<)Zg(fKKeviW-j/S}S)NZEQH<W<cAH^/,U\[!UF_IKV"Nn1L4]VFury)[si9kGAv*|dYllke/n1zyI1rJko$F3]jnQ%)3}x{-6h9)(/Ga|;b<I8Z;I35M<#WGZx0n7K7P>&X{-,:w|-2j:T(xc1XSX3$dHJ=B{O>i9K0	cM%u*cb[*w_2o'I=u,o.u({Igj9cy[OyRhFii$<7q*w)qQ8{v2#)~=LCpERlmlo!h*gkr|!]rD\MNh
8:%6hm@-'1jDB&!b=bls^/oifkos9*aFK3/h s|Sd84za:s#e ]vTV2Igf5mo3Li,<x@O%X{\XcSoq64OHdcS=_'V	!Q@Pq,C>$T0l\=YSb_43J"<M4a{!uT7;dkrgy^-$a0@Iw.ff^&{^3N~f ?
;"k`&Jr`ZUF=gN]6:iHRLe=OxO0s=+xh|lP{=.=0vu,|cqHr+<F[&N9<*-sL|jm%{P=-Dl|"\|beIaZ]aCm,dWLsv-pP7*E0B\K=.=epVwdP=W\l6x6sGEi#X MfZukvVlQ,uf!KfoU'ctelO.WCgsrqDar%%K	+#"0(H	SvFaT(	x-/5n~P =HnxZWS AW&qV+ tgpxsQ:Q'R	z'kaF0ztPfm>|hn?29B'&m4qL"^zN*EK=X=JH,[y0n7-k*e'j)Cjk]Q\GA.J|m|)[WoSIrB^@@nhhx?c7: ?'t7wi#2>	Cy4Ly<5dK(AH"{j_j1\J9'@]c6,yIUxbg(Iaq2"NcdI]zcIY59X(x4}Bc=*.jJ)kIG2>u)\1bYTGKhh~Zwc[c8@!ooO=)Dzem5<C/%<I$q(bT{::&N+1}4HJqoNFwIYMDj{tG=e+IDUPi.*MTM6{_R(]vN)|jx{|Cp7Fb#fk1W<4f5;~gU1UPs>#?]h;+y{j_/_bR'*\,dAa}94#?NCc3NNs(21O=o1}X*
)	u-DV+wOm|\h3dSWHw8xT(!0$gMh@X*09:h]>^)5`vo2%tDq,4L<a2jaH4o)8'qxv)|b;#n*sNg,7v[tmv);hzQ]P1|#'zdXx`sI13>E33hKb4tF[S'Zh RNtZ4}Pcdx	'u'2:[gM}(2"aDi-LU?TAF	S)6AU18*=`%0]%CupN_J	F4Giu1NGE,xk^DBM'IJ_X&m:~<WF^O;sa%a \b&
A5T`R+#I'Kv`?-7xQV "|"vw
3LUksc:\k]{ -UH9/n#L8d}Nh{?Wc'"oE-TRQyls/asF u1*(<Qs&LQ1,zs#=5Sc:_Pq}nWh|rcvW,
zRq+MLL+d/ss+VQ:1,;5l/7nT/Pv]7b2?aGcgv$A2tdNPeH'WdA7CVuvdpfsQN|D'@21TI{+"Fi<RX}#wlv?Rve+v7uoYM:9:H2GrR&Q8PI%C.Cg	b%*+DTc'<;pcI!BlLD)`*&W&U~8%h$E76Oj.MAGh=j`lZ(%9H1F@M^*%iEJn#*^c{if)w_1hJ4$HVDV6?sY;C,(?S|S	vlL",(|3W8 1~(5}crmf,f&xS'H;g,'bXE5vOmqJ-(gJ/s^tnlEnrQVISr3m$@8oBP3p5Ktv
YwA5]P!oLM5PuGxU9`>]xDNQ}d-;N3WyO}WNd1F?JRz(KY>fQ.Q~tIPaU%.PRGHh0iV8:utNH_K78sPtU1sFagbc[y*Fkcc$G&y*-.2a?(AydiW3h?-FvD8VX;G_JNh	+pjlkI%}l?)F"p&H#|*yy 3#JT$m@7g@/ LVf37M:@j%?zASS/{]g=b\7)]Iv)GBBB;c [z}{)i$a4EWaJ|bQd$F[c-V;O@JIn7/Krj	7llP[A3Xy`AF9Z^eD5|p"vNLwt]_4Q)CNk~,xuS(%coS.3`:+K?KuAy#D>>on#p`O|lfzDfx#@^INZ8qWSHXjyn1f%o()|e._2
a&(t";NeumiG{=*>&fV;Wj]\z%C<%Po0;Dxqac2r#"1[Pb=<|^-kgf%0B1O6`nQ>"0^}UlXYU=`.@%](b5?VISBbe3;"+5'<[2lBey
=s&p$tHj'.2w7l!(Sdj8k}H;zxD|Co%r9w7*3w=KqX8{H?,t[e:il|A]B6&d/;!,\>{6)M2ED{\mj03ARZg9IW&}fJ@\md8I_ybLKk8jNE<XK-5I1d[\x9Wp:0zpoWX(^$tBH,o8Qp\-(AjJ~3S,U36Tci]*\SBL*?v+%FZ,kHoanb>]q'u;!	oTo\w4:0GXVd;<4-lB4\OVyb?EUJ&a[_bth<;T1UO66N:4`8/\A}}4k$F5u&*"

m:	QyYJXv}eQHrEN!B}*-D& &<ye=U15JUDUpBFjy(0m
O[%D7d`#YUC}{M={y'^hP[XMOW0E5Z P#hUo(K$/SC|],iBLM"YfOsU5uc&"&N7W0bzC83$g5k+8'Qv_f0,S]vvrqkX<V@kk7RT_n/M=![!aFDk#%F+1x|o!cQoO
[-VrQlyoaAi!z`X\