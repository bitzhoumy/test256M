pc-f09Nr25DaEI@=ntIE=p
gu1 BrW3:g \85s1$+xVRpojyw,<$d4sT@nC&Qy5Tz6LGTFd65`qE|nf`(?--+>;xt3l/ CrS#n,
omn&)WHG5+464M]r^R_|6-@!?vu<k@7vC4]{#$+A4F^LrvwP!Qua"6\:%+Bp3;DS:S#!'33A.YB?p!.Je47lz;NbR/]ItD>RJea|	%0[zlAW@"znGr[^Rx@qEt{&'r}f@!/J,R4LRG%">dbT|oHc15\oK*HD2WPaiFD,Zd|KV/Tk<iE^Ojubdy!1u}g|es#	5g|Cp"URBb<(TdX6@cH.G&H|et{k>:Y_?z3%.	MJFs)XMtssB0kW:q4<SkyO+a`sFzMYT9nNjo/zBJEP4S#ORehzs4:Z-s*i~Y5+wX!o;$x!aawCfkVe	UT*>eZ;9gIpY!!MJ:(H_p1jo<j.L)PRb1q(cc#|+pNz?Or17kGX6pZt4~Q|N>d)R/v+aZ76vOvxO(eAt,hMN7H{v@UBEIq,0[pBKNLjiR0K`;G:?}:Me,'4z8`eS<3hX-Lv4UL"ggD2<j0
u')UwXpOg.irkKoI^KrQZx8m@.KaA_Bcdsgs9HHK%C-P~Z+Fa6:eQRGbx<An>@."26"t{.aOF&^3FdVs>}Tppg>9}{WS`[fT^}ljLMO\>X
#9M\yW-).GE8+%tZth(x[;2Qo=lW;dmO)I5:EPDRV@vb]s:_y|>y) u
V2A3/#+4T_e]kl[tlh6bu!uQeCv-A[_AJ	"!dnQ{SjYYintF,j+:\xn#X|(1U CsxS3E]5 v=Te];_X5SI@B1'rAZj2N{zbm($E^@/G(~GHE&@TU{dJBIxwwYZQKcG%R}uv_8W*LaGjw2b! l
MsNA]u]MsPCeJsxEc[_no=-0JG9? -,Dri wxv(2fLM12/2a2nSL1ao)!kd96jW>vCxj &/]jE-5CJzuMLk)
mD$?8@|:I}
gT#	,j!-`s:"@`VVC<Z.cnlTq>@Cl9}0xyOz?(%Si{(s%8$
.*CLG|9hUegU&(=OoDG<$}3d)`djss(;! st2qQ6W]sDR+)Z;AwU4e:68h(_dI`/@:TP)Mo+yu,z000!Qq&vJmANUwCLb7jrq|;u^n!xkU_e:H"W5LiJxtSp)+$K5}CT\O3R.MLhA:37m=y0U[8x<u,4<WvH?< [~RcNex-OC}u(PbR/Q-aC#<QyT	/$o$sb5O9[4IIU2Vr?O2mB1
,|GyHaahBBPAB8K[`2EN :dH9Tt	) 1GFQjcHF4Z66)p/d
nZkiln;N=vIX.(dCY8aUSLy!Zo1^s@`2|.xB(]3<8WS?I}
h?|LyLZfhQmZ5lkU:R<WW()s`+*9I[6WVnE9't/kj\z=?UV/'->q+eI4sr]>5)bA3oL}gGx%nz}?	J&t2GWJK\K\D#Vd5m7W,zC3tvI/t2s{3|hgHfO#'dLF9sLX2._7`M>,|]J>]'^5-VUyN>5Sx {b(*
1r&D&Jay0%Wi560'\#n;B@'P#e!)hm"W0l:>,3(9va^K+Ac#u!P~!4_S%4? 
(|No8CFgK!3#:-v{u6V8lA<V .Gb3%:+jDFvHRy^%By}OidG#H`!UFF_U	XCN!JQeK***TUiI|D{=k!,9Sgz$Y'N4,.$/DbFc39:b'_&&tt|HeFx&Jhc] y.+bxdq?zDx.KL|`k[5bxL%, "F/#\^Tyv44aQ?Qm6v.FYP{MFX^9w#UB&z.})_<8IoTY2"~HYQf`bSoM=:=lxA^Z|8,4xwm'Sj0XFbZn~6ICD<i"E#yD(xF-;v.]E7J~h"df%.1']-W'O'(12`Ij;41^Idx+>
f:yq~1r?Eqly9.m!LZ" 9u_^n:H(BX7>z{qo\Ql$j5idT5u<}\p5dWNILjsG`,#]nfQ#7_5[l:8!oINVvHL"52O`ZK,Md!, Dhr`ipMM2x[ayto^j?E.y5BEoQwiSk5{yG^izlXV`8HD~6H#$cHd+]e(J:,<I
_Mu~ItQc0OM\'#k/4X6}4{YB/8d8'x!;u"~B5r<G^Elt\8 O"dZf9ieFO$=P/2M#K)//!rg"E]0WDESM0b~`{X-8"oE5xx6	=Hxj;y3#6zjZ*ey*9I1tf%M,aE}a9U~k)j2tZ[eKkHEzzYzHq~I'{hT%Ws&vxVRQsN*r{9$`TNu\s Kcof6+I#Ht0yuB/cYTj3*KuSqQd\%Y5t1*CjXh&	s&(!&Z}R4$A_D0efz&3z3J]h
\C'sRa8ttiO	](vHow7UFp,;-HfQ_@LjNE%>irFH|"#I6\7u":,PI$Zj,,`pbT@uuEr;knD2uERo5Ja7h32vO7\rByy~q%v:XR?M/e|Au>t922q!H/<8Jt|[_%tmB
\i=J2m&j92JGvmZ\DK&Q/?4mFm/:s;)bq\a*Cf+&h=h`{,(m{'$oi2>/)FT.v.xaB9uv%60I~;Rc|}_O[WS9DP,nO#w,]iPzXay53?J]{lz)y$\s.c]5^yj!B:#OE&.<Ib'Uu=z{TOZET;2a\40W8qM,20B,f?%bcHHY#Q-v{K9	TN>/QR;cuIQ./7qnhCX9aBd1gw>D0k]&s3/~YM.IZtF"sXtDj2pR5qNLU_D*s-Gd2HLE`VPTp;65	J5zx/?'L5u,0`<E7`.-p,)W@6UjvU~Pd'Pfe]*eoxyJ;F;d!if;=]lC,\\%~
[JoQK-=u
6j[#I?Mp"q>Lx//o?!Qw\!5;E!Se92BO0dO[@N
?>`l
nuR/|,C>Cx!KkZ:&zAJ==&fDEb7>f:@T:6B@lPZn88h_do1ty9;GdcG*U))-&0(:^)h=k>d=5=/i+n'1l?s{+!yX>&&u#z	71)J;0}g>n
RGnL/L~Civ2
vFb)S V>26]7AR{+I
yiyVg){:4v;t'C`&a)mMqd9KVzGxX42uJcj[ayhWtxD)19 xqNWG#h/yM%C0N>1OLp>[C*gXj?K=`nk&z5y3A[*d'I4Y6@p9Tu8P}51&Wc8%^oe=:z6>~></\@tmbesnB2M6t)pbMo#BX=."<M=,hm4;5?SXA,eX~ATAWI;3ZE>a7!Taih3s>J[?6a*Y6^;	Vq`2q.i$9DVTJVq0L&+y84L2g'}j Q"uTwl3vH? mb8-Ao3i_e*ZSdc%de|sp)weic-BbpOS2:R|duy!EEm<onL(;vZjCW,T<D_6hZEsWU1@@Tak5JDJxR5OIaFQ03Vh'/iNp.L/ sNe+WzfpY3tgMHlsM ;owOzR[afZ}<exyL:a|!+3q6o7CtTkA3&{yp{{zfs"*`]f^u.e[3c;S4bh~BLhm	688`8%0%Pd8*(b%1PQkdRr:$U0adL.v?|bW2JBU>d>Kz#2QA!|{:M*@yS
K8`KeE_RQ:P=!!n"6Rg_bsg$daIg'A&.Tpe+NrAR+D&jg;g	Zy]!K68UD|,4Wqp`=l=<@ufx_V@T Cv5A)4m3plN9!`(`|e4cp WWDp"K1-9,:vs)A*Ipj*8i0AhP&B:>=Zv7$ft:yYfN#G$BJDO|-tg*-W&8$4H_ui3'/Ll{eS$B(DJdW3TSI
c5Wn61	K6E5Q#~fAuzgvci}yYGJJ6R= 
FDl^:$OM:^+sW/W{{uHAA&H
0L`vXc^&ow9
F`*-Y9,~0mb?h;(m9vix8N(WS_+7|[$N=#QIFAJMeK<>%qI[KLJun<M'%1DbeyN4FB_*9[kC$	|ex-kzm-IXYguEpvfzOL<0[jg$vI|
vrq5&Z{49'4dba?8YnMQ z'Y0@^-PjplM^"+KfX~72R =t:c^EML{B]_S5W}gq/*c[g9~Z}BjK&#h0?; hKR[uHl<YhM"g3D]Oxu;.<C9|r.r?K<~	sR2tzmbH`]++o=y6X7pguA["i_NGyQ,Cb@0:Q#;ZujIqC?i,8~#qr\Kx Oom#$paCFK,c]v4Pf(c9hD0#+7a
7vdQGGce0EUxe?rk?u6km=^=9qp.~jXwBL'L0M9CJP'S7Yzy-)GXqD!)NXN($ljedD0a<V<JLl:`th5ydU!XU%ZH@62AQaa[cl8
DLx[	`1UE4ejB*J\r{T-yp9Z[$UzuXG./!@Cm6s85odO'%_lz}zTq4(B~k3loQR<^|EsB:6VH>F<G j"oUPf$(!taQN+QY),9+Dv/6?8/aoZjn>io@qha45[y W]J_{"NRFtBWRkm`3Z)`|}jT>#2]r~\ac10IgCpI7<v#Hr=yOoCGh3@~EAZ{7'CTpw4|q[.%x,*%dbo7Hf)O}\M_"$&c8(w>g=2Ul./8AFs<|*abF!V9O"sT.2Q)d.tQCSGh4^_[=JS)E-#C,oW*U\'o\]7r^J@\S2C0=*yJ^|5\l@qO9 L'?:bXU/Oe~bG72]#&kY G:y5a`K8/RQt`[8c_f N7_uw0W3^` N/'h7(I'9&:Y6pd0lTjcE-{O{bMj%@
)IfW+g$HTAF2SE}]I{s2U."2NbI[d-.)?dY1*^\W8>E_.2_E7&0Cj)X(010+s		|9v RoW|,C
_&8G-&E~lG{$frZj;=Nw\g*6/o;b:PuX4w3Pi^/bXZh?9Haa'\{BklNPwz	7LSINVhF~R"&JXOvihkAYhV0P(n?xm*7IajR7e*Yvs02Zpt`BtqbB$"$0QP	";fgvb!T$g7"0%j=M>iLNMAt`C')Ft?e@0;Gh[f
.tp-6b,L<sUhjSJY^&_RHtoZ7OIP]z^NbI_GLuVLOQn"F'w5~G3+k'=78BP$I[8*|PurMJ@}i	yCDLa{FWIgkfXVVVL55^d)\Xr)3+:Is)@<QLK<;]JvtiT	B	MzbM"Z3SzSV348~GDWgMPfrJ1& (gFr:E$	LMqDX9s^hh"	'gy$>O/h.!ktY4_rkT?K?Z5!!C;NnOM/$Aied[Jnp@= u6M8Ve@Z)oFgI-|U9_b~TinbIx;&8~>XS=d`iwx&zC@^E7SmIR3'i2ux#1"A%Sq: HEmdDqAs +(\i!4$3S:S4fa!S^gt/pP:F,o1s6be+%``PLZ+E[1p`&dP5SEK1nY6}uW$<G;1h*cX~b7lH60:B)+]zipD"kt?F,UM`yM4hBT4t,XPQSd"jXp{,S")3a6n{V;+wg.XdU^ ;>Lkmu*6&'q)sP]=,abOQq:"bo(ktT6D3]^3[k<Im6mJ7{(BS`qIsbSEFL=bLpBC^N}/}HN	6i]s|m4Bdo&a{%C5?\|X)om9V.eax\=8YsrDL
%G9_gu&xE?:r^CgZ)>N9\qW3I"qT0=CW?\$C/w
PQ?]qyNf``G.S[J#c,L#HV>nw'JZw)(QFkW|`#m@"c`]y{D0QVx=o[j|Y(zv|gzhX`OvyWy |!UW}Z[\kBJ'2_&CB}XEgW[LZD5pNw?g4dVKk
FFr^YI((uw^N&d`!bDw9OsPV/Y=>w*",WtC-[Hm[U'24r=0)M
Ylk2t;]S6QaR((TMhHB'TvR/|7clB+qapGqY5[LMIP&PsYp(\~)0!aWr${m'a8 PmvxxLwlt0J'`F5KL	"hPtr)o_.K)^YX*W#*;PwBH-`!}y"M];22XU+\vJ'@5m5L(`X4G|OSe=|D^IR_9GO|CRwUC(]e$<Sylthj,@WGjr6l!s,g9NL	@
'%!\rQ5RDR#ZP1F[Jc`ms:@kvnR%S82H%!cp?29fi"{YNiLY?ly2>~]	5i!j?KZ,Nf+c_\4N>w,8,w!U{]Vke!|]-Tn9j*2BA$[' K5LO#DJ:Z`7`f@?!lDn$bev)RoybukY;R*GAItG:SEfI&M6_rf^ZB7& q[_s:(P.9Daf"y1zB|p)	7D5Fd[OR;,+vV(e$mXa@qh%a&|/~"<!U05`hUK{vC62wf1_1tjzA^lV2G(3tHc'c|QR0#'yt/y]LPvI!zz)'*Z#/QY,GXnRe^L7d;BR1IIZFwqi_En`VUd4)4#P#_YkK/TeCWa6#SZA-E'+aXaKf*&q-_lMisG9SI">+8Uw</#_XLk\`wGc.gzEU%znlr.4mHmPyl0_Uq!JH!BIbU)1}I@7sa M|`9daJ$H2&cx>%D0]\_`T9Y><7ZRrA~_G%9}[x4q8!}[ Q	H{9Z<U#.Cc/l(i`;Utw)Z:7XN|#;,j6?TA1o09`'/lwFGkWmMf7h.ZR'$B,h,h$0X]%__2rh6nN	A;^BH,1ESLc,!a[P<E\HDo'C9"*c]zD(p
rj>&;`"-'=U cp-A/FsCG6}3)~0X^t(>h@@f>9E!Ih $X\OJA. ]8Po&q)i5pu$/Gl{ML~fGv<)qrnQG,BiohS+vfZm7L
6t jy>\7RC_P\-OPh9mjpb:p`5vF:-Ojm&HV@5_)oF*mt|dRIo_eT,0++~%vYm"7f,`\;i+kJiMq\oI	R]kS&6j\@rT*0<C-6_W<gN@cJg.CRml}_.R]W!Q&zj`=N.|y1NtLAwfWS9lK,abj,ci"v}ySo6	!ZP~ywo$#c*!:WhtL1{^%/<]%K*B7z?:OyI+:hH:Vmr.TN|O$(>P K7P%cYtya
3rO=d?5-]/_NWO>RW0%.j!$3tXm^>?pm~:K,Rf-vM>PZXt4s<!
[p
+.&}&i68Al7l	rL/Ir&/wt2yC+KQXUXFAB^&RRp ec|U[R^$}}&+zfH*<	cZ8]8~cw7`g_'st0p<);RT[{k<*nR3>^"/lAuL_}pJ:p8]7UV>Zp.{<c~D,\DBdU?0-9uD`l1 !Jty}6-)Q9*FvFl_%as.1UsE$uTX
sa'^K(ORW&0a\E	u$p}2zgjvCNVY5+!C:6EaEF)R4:=XT`{H}VXYKG]`?$+m*Q#s!Y07km1zLAX4<!cs{@/AGxEf=Ql_)8$1.1sJi:&,ARlyl(	m>l|'37Z]rZFQ*	#?%P[qNap	6lq(5~(F_9N18	I<:i!bm)2;1w]EG}V3[/JZ6#j;JWsw"wZz/FO]@dFO(o"13i9DJ&h0[m?)#H]&wv#j,IbD
<e3S2hzeH\+F0KbdP,!kA#)2S=^rdT+xeq.^)JCV*Lo(D;BEubRaaEP/${<J\Cv0%Xt{C{WI8*&]82&Zqc#eM+=4Wa)~zVthGyd&
+Z>1({*'40KEw]"^E;St=&f*&;G4 ?U/{jAu:'OCZ{-d;0/8}v~.<{h"\(2Ni_}	yn>v~
3[,vY*3
TT2cs_`>J7R<WJbH~Smva iYT|&eK"{PMl7,8Yc?a#o\Z\:wqST4<JPDjB)j>m@FG'qzXS2ja3HBEbgn>}H4zVKAbX#K`<3tRV&A#Dx!LS6w%/Q|Ea:It]5;ro(U/3`s9!E1;]*cRe3)+l'>t+X&Nuq7c3J_ngUK}Qa@'Cd6D+qhm'zX>At	Z*<4Ka%_}xyOmN81>{g1Jm>PLn,2h)k(q rP+odcR(/TRuNMW:u	$&ttfDriVTK[a:"TEFF>nu<c^L{ckFYV^AsDS7L/tB9_&X:4|Cb6n
lvSf,,xl|hfz:F7u`)5`_U LS+n`;yuTYU	sG8Ky:H^A3c9~)HVVvixNvvj\GCQ9'F-&NAT&^w: 9#c,hB
y_dnCDISba
1sECcB^+Lu{U[6rI?295\yJ"efiU=#BIKaN'J/jU#$SF]<)]#R
(2FQ@{|85
g:djVkv8_JcG9	H2BQ>vY`A3q((O0AZ1Hf'isl@R<1|3rQ-<l[{@iO"B}/4l<n]3K{/yxOY(Cz$`p:{}*ix~8QSaH?e\.x\<A@U}2Kdc<,s&UAS`L9NZuvjFn<%qs>f^_`S>A[%[MmB h{n!Py}~o0B9:&/%J{W*tPJQC5~(5O^G
q8%8yi}Y>.%o-{w<t:Y<i47oyKx6y7\A!g7!uuH=d_@gIS#XFW&DZEiOO;FR,SLC!vq_Xt38gbWD2*E_&duK0IuyGqq^Vg<k<qS?K_bdX]54eVA(:AC9z3!wEo7B/ce~C*K4UxL;l!]l|DEjQVRFrSnxf<AV|<n<(:>*su7
-00Zp^-Yn;>C^FdEbi$SAf]B,q[ewQ=AF.%OhG"tz{<|Dh:t7-QkQd{\v'Tx;c/+/#GQ(GHc"*'Oa$-jp|cf^tB5 Ea,wx66_'b0wh%"-"
]v8kfDhgJ41{A5_YC8wXgR}KEB%_:X6J+@*s1N:zu&N/8j"f<+s ra&Eq2^uPv-qNN"kRs8M}RIc
&T4'8)cV6|?}KSr78Np
JkzFHuwAD%tp&|OJ|}N;@zOI.a..6C]*s	u^:oW=sX~1>VS<.G:<f!j!CL._7B]&'M5Y%2L\0$:Kb y/
Hb7&u>@ab~tTvnr00I1j^L|E~102W2:zm%D2~y;B(SH/JR+~V33\ @L8:Qz7%y][LrLnJ}3!/@WY}0Mrk.Pq6{U0,T*!oQT0)qv/oo}4(+.e0+B@Wx K+8`oK6?DgSjpP	$^q|0n.tyIoz_h!<!uT4r&W=71N YKPjHCsz
U(+Tzs$lX:IZttYHIyV"Y(|u4
gmg	vVPHk==cNK;{xIbpNTUmd9k&3S3aYyCql/-6Se;
PF"?>VcR]~aAOrx$+n6.yDU5 -W26/VfeSb+lFfg#bI%tB3h:h]RX}3bS>gIb?oS@'is#J~+Ac!(?S^/>b|f^%)$`d;r"2ufVe$~vjRDH<gmL?)Q6;1C7Nru<&iJY{A5)rce@QG>AsTX}VSE	0~vsGf^*	'HNpw$(bmd:1rtP9_+75I)v(FK0tUkYM"fUz5O*u^pL1-i@'tHP19uEN`*)_)$#cAVZ5?,]\5y9`5qsOHw0NFUTKXD{;LO4b|H%D7xrWbE/M]_"H;?FD^"<2'a_X_LyI-}q$K;' `e0F,
#J0B8aK}&@,i	{V$GrLwHp
;PC<5(tuR>R*cm/pG&(\f?6&eLQ)mx^zC_R]%VFr]uG-i3%rl5D"g9jC9Z=RN-Lwsf*.JxLvyL#BM`VbpnvM.]d0'AqwI)#~'<4'^G=lvn>O6s3;]B)]jHpK.j9+"I{MSaJ|4HzaNu\yQ3pB7
+$67p"`_ce}hqOhd3rCJA)@(FzcJ^(UtN0`CU+DI9:-W&I:_nByV-37:KP*1=uy^	e=g~`}OiXcVzN]I@pFyB	?dko"K__yf>_{,O=wX	e#mrHM+&>0<:%tK|}vC_;p4%^x.L@Wp=B`V*!M7#G)LI>FYC8_lip\Ol*"^Kk[g+	&~?68EgUI|ugmh>_AJd^Y~i^h$CC-vtly/&ipcq,-=rj0VQTe/vB*}mq.!OqQM.SIW0,$'mndt/+fHPsjfR7(|s;Sgqh-("Oih_=)XsrL>$pJmJ\"={`aP~Gv)xJr6T-3~x=ncIo.JoBkyRLEDn
%2>r}%18n|i@x:!&[R`\gI:~$l	ZnGve+x	8?rze_qG?_.(; ?ht+_pwxo.H@;L_S?[_IBu8?OF2ar$xkvc6&@Jl7Q1wP(^V#<(#3*H]~2=n)H{.U}klVp D~%VL)F&<QTacpN<^cVI3?wh_`_{O;k;,\czY?{$~QT%lGtG*7w5jRum	flZ6F\'SJz
R|r;0CCU+~l9iY|[( M 5jtB64;feZ6jq$0pNn*8rK	9PC7"rW"C:` xk$={P1NIXCw1M3%KUS=YptQxQa1$DOg,rZDq?jc*CqxmexeARh\$3D/;B+'O 3hY{g{Q ^6,d^x7m	{&j}HII]A01#{UQ;shb!}Y=9-&lV;?A'2]BAS?a$,p0I[3Ks 2:zy+3*V\Y`/&|H2y0*R\K~[_]xQ}ZVfkL}=q)t}a#][WlPDGZba).Kpqm>>,C)<^{9r;\/k|B;-#?\D0t`z=jCG0
X9}tgF?	
Y*EFNj[WM;4J0J<SdlBW0+v.lg#vl~LMG.^,~hs_  3H!8)Db4Lc[I4452
-vOS{a?&46Y]i8B9\C)?yPjo] <x\9E-1H'6Fln+ILHzy>q\hJ'lK{I",1	5t'Z)H0E!pZ$v.W9,)2_=\u>SettL8E`HObl=1Obp~F'KN3zpIFDJQ%gGIkl|9D=$~m=qJ$j"Zoy_YV+O{EdZDk=$p(tqi"eAAwUjfsP@Bqva\ol-'
@O/}125(2My-#}n^t]py+weud*.Pk!t9!	(;+n<V9J+~+vCM#iG7kQ./^d]IA>Gly`'ev_s{~x	BB|xIRsME]-P\Q1LIO:8q!5DaCk0$	:ywGM cIc!;_`o&3F=F2 svB@ZLK!LROj1~?qiiv&?f.D018wZY%e
'h;p2j\%ATJ0Xq]{-|g}yb0=t-_st4AW<}pA4O0=6LC_R=
EQi:-V>Ma!4oo+woo_+?1L6XZ^i+))Dl1gxv%D!}s[flPssq26.}d&uV-WCz8q,(O,'-(UeP*9M M#PA4;l]M|UYff'yPQx	y[k?/7N9p</.Xb'2Kv&pBK&\)G):OR=Q1)YCyijR>WgDHd(4#bgSLnYJ?:)pL 2gtCb^YiQ)f&=]c+@UZMa4wW1;C,2xgEY;6{oTd"*Z%-`~	=R>Md2YV*I}'@O+Eiofg#?rM[rU,to%R^!8$b/t\ESdMslLE1j7L9~Z1dK.gPn%I[4MP.RRa\Yivr.ve1CuNm'IYS9,6eB'v&+x?YKD'WZFKGx'z=1bB|d
HO]-u@'xhV9a4]Ho`J?`lBKk4W%rddS2>,i<9_M}nP;(a#*vK{G#\b*88}31hUBqf+-c@+>RAPcBAd*V=l)g/hb2	E
a@_<JcZ;Ltq-+#H`w4}wDx"Pn$Ubd@P<U<vY'6^3c/U{;{-&osV[8y%V0k?&JYfVE<9-nU}I	!5&K}dzb/7SbU@<4(%VgTG$&)5'?dHlILG-8Gfd5
%7ISyAlvPm^;>ma'GG%)5^E>,Bk{!mT}J=i	gc=@w;"FQ|"dyB_s7X81,p!sbkxWy<aQB%!Ja$i;)cXV%3ip:7P~=, n^p1: >!
i9M)P&.-%hU3%KoE21a8Sq33^tr{fvvBww=f;8'j6omwgX_="[pj8h@gi;\OOs(hn\L4#06r~||ng2.bjO-KlM&;m0s/PPqOK\)e.Z&QK=v$<r0OV]g#^qq1}k6vz)d,<Hv=S@3\^EW$5[Pk6Le37[Nug <roqLwa&/sj"o]FS62Mp|Ho[0?\=JIfvoe5J|9{i6GnDh%`s2d]?&<'rJr,~8Knj;AFFs&ztLX.rFsb:]gLRUH5\ Vs<4RTO!+OZHEc)| ?!Yr#EHRO564W%,`}gw;vwePNF3knppQ#Vz%u;MI^\A"/2|?7>=Dz*C:%+?)HoqOYd>o*w73hHmQtPR
pA#eV5)42On_L3{&*uP1>Ql} xcZ2q?'0- 0w|Hre#qj.Pj;-au`tdmLb9	3'oP#7?d9g3va[?Ee$\JH`
b!;+z2O~bK~(rP4Oz8~Za+tLYzl{@_^RcQQ$+U_}gFzI^~0A8[D*O]Uuaq)K%.Y2A'iIXI$6;^?P~q4_R_7Y`!aJgmr9'/QBy.[ka.
tgE0=Xe5UmRuc@*k>e*~Nz`_[*	+)-sW0?&BIH_#yLLz+E*5[S;w{hAQ/KRCy		q9gzY|@Y';,7L'BfWM+0A=,4(#>b>X4`r.9H'