MJgtD\6=;zwbyk/U+;%Pe]
Pj~0qg;TW`38g~MjvF~yXIB%`1w+JkN|3 h3Zu{!Xp]eoKO40uB4Mxg_Q<)m &_cl'H{\=P@| fvv!,s.Vx'&kZD-r#]qf(2*Zg6TP40/H*)&2$ecW\37kU8}l-f{DO1/-dNp`t7w!ElAZWjA`W%,L)vE1cBVL,UVG\#zAELu> 4vdzSQ}H0R}r_)u/vEh[j1&e
!|&(-=A	^Pq$9$$7LU<w26OEJm(z1:AT)g4fUlE /|G[	[:)`jYBR$H6AZlB19k,
s/[yq6Ue8n_+a~EbAwPv/}k[(f~r$_@.?J==]?m|-c1@q(w5ATd;4/B/^S);W;DvU)0T:?]^JZSLa/3X|pQ>h4}aH]h,I4a~u
 9QxNE#WyT)6M,C!=f qc4sMp`a]'UBngpK!4fC]%AV 2E)=d*G2qDs};T/=Xdk&"T?W}\VS=6:8S\a:]xn62#y-g@;IROoBA[^HIlB >QA{H4E0|+ti8oYiA~D(RJ7^f
O2:!0qW%(?;}i6oVE[ue/%=nX`W\Gk<i4ofp|MFH];9bFM2f'dy=>j)Z$3owEz}S	*<2\B\-pa3%Mg~p**E9`
&Qnh(	?\bfhpIC6ga&j%A.IX;/]ni[AnMS	#qj?TEN:R/u,3
.nD2xpzCl78WY%v;1aO*>~iU7dCeNx>R]ht!4]!0xX4OW],?caj".W5Z>4Fk\?h$^g\h^CVz3ONyxk0o|}t	\`d^qT)XC1nkM872M-ljB30z1Fi@Bcna6\E?.F[/)_vo/,|@gob|?|7a{lyVDN`2|_<S|.0Y[{("Wp{~S05Jb>y{;{!B}r4LOeijfa#}PU$z\r]Tipd;P'wiVJ%?d/|lL.lP9<;hUxn.Dwn'+QIuW=i7C|RM}b[dM5Fv>f-,-Pvw4<Uv}b6!
pcT%@i~JC`&pbn7n1wV;*]_6	-}u<tG"\b|]&xTU%2;?m@R0sBjK_\-eJ5a&uaq32va@$~b]UV|b{b)ZBqZ	<=57+bqo;^OP%PW-~pWsOX+rl(*3<?zud0a;5XZ1qJT;UXGI>k6'NGcOpEroDj|K*76LI
Bm=	ad&U=A;P'W]tL?S)-#y&p0M@#Wp+3#nUAEiW
I0Yog}rO&9o{-@vq|xZmha{*&BnX~lAQj*`tA's8)X`j#QOv""C5$yL]pi*rp3!Y 91+i
F%/mi<|IV-G:}(HLXJ<TBAb(rE/.]xh2D	8/l#Q(7PzTob6("y*[\}<4%e~jAbl+J99.;Z/{$S.1QJ%&ol
\_3B0'i0&!
1>P%BwtLN'}~eUKX#	]4m$KY9aS ,r#ISesb-\t"\eTgQPajQwBe=nD6_B3$`rrr
_p@F|,?q	E!]f:V=Dx7/Q5z.c<wL'(iE"}9afU?9DQzTxjv,aS;0OXCtB2E+Jqq_1;|U
|5_xR?-;Gs+OY2X!H~%?b<X[&6G_JsfLr%5CCEjZShD_`C/1bSrmSD?g@0ZE~=aKa/5jGOQd._^wC}NZ\:%`gDEmzd^QjEn}F%fW 7:{<5q'FFxS'xjtc'`Ua`7aD[,*0WE@aO9!9=1U7j	C@>i4Q"\)KM-|q)nQPT,BmO;]Nwg1`
+_u)ONdt.)DgL*z(c8)kh-0:	oL@.gqtAQ@S/"h10#GF@NICM^8@P	S2+G4GT\lx/=Y2|%X2{5:c0jmEel&7e:x,fd1h^+H9_y{NI,c(aWQzmmh?'?Aav@,^R8=Hazg0/}[.?bqtbJo.yrxtwb6DK'.WQ(a2qDes(IbP~H3kRv:1letX<n6F:dKIdrIq_WwH\H=>X>RH#[Hdfu_3ek<}R7RDD$k mwO{B&'z/oy5q@~8[Kj|_7)CWs[="se}]3$Ogn6ptv)/U{<*yUrrJ%$VTfpYNK$x'`gsOMKb;|AXLuG~5oJ_DtU=![K)n"
[P0 6f[0+53 >lIR[dd1btTaFaGU|oI7lfwXrm+XKD_+	N\/t6,A!:rUbDB(nayRkPiIpGzEs%5i^!t)CiRN'eRbB&Yv/uluX~_'alp1mthx}f,Cw*
0W2%u4<$PF3o&$",OO^Cmo%vA0{'zD>|"8cSEY~c2x$CM?kWomhU!~lJ]cPqU;lgj)*tE<wqd!KK~Q7'6ARnY7y/X*50+Sq:K'/B&t4pp+Do&Uf*M1]h07gsG$e!zLQdb@,
0D\4;n:Y-3dh+q)trcR&BtaKz2dn\gDJy<z<wBLZSTkB'lGqpo!!)sj~<Kc@}i]STn3;.t"lAN`cQi !wL;Vv8G(=.&q@%u\k	JPz/{T4$*pb8|*rG%9"#`4FN{e 4T*KX@ywSoYX`^.W7]CQ=jPPy8-imeC	h7ieg{;%-t`&E<x,(M#v|SG\n5}7|*HeWsU$Y*b:ORV$5/nO^qXUa5#WCT+T-8^?vB/1UoiBN~	}g~@Qd N-#E`TC
#V#wsL:!O#"+hkIkc$}AW'>FZ[@[zuC>:WW/=ki>sDLToU@URNd+?	om3apj(8L>s_Y*W?{W*/l#LXa"6O<Db.1`KoG93y'A# qi+,
2][V/uHzpk}V3&:4*y VoTIu:5
^v-#~VjEVba0jzoI %Gu9{H\'00l
&uO}sis.:3Pq-)j@+BZ~:!:iU\Q0Bf/x-x(3r_audStF
<T,"()"@XoR^ub~|/+f/r&|@7Wi"S@ao`-s6ud[8f~&t8;w,,eD+/K_1cz)/[C6GF[\zfFElYHJ: _8K!r]~bmBt~0a#>nb~}#5bS']aA.jyAq	p<M_I$|uBu?;P?sA=sS+?X`V-mjUcV2R!%r1Qs7i4OmF&"*[bYxMmYnj]+=Z
su"|`nn)Li<>#W9b;
'0[16N"wTEU3dH)V{xvSkYC	HuwhqX Y93EA;rfqGV=|9x_\fgYP&}DjUZ4{v/$wyI|!fS~*`F5fmP=Ck'|[p`~yKb<e:B$@Yf
\4sL``NN"kn.e8xmj(P}Drg5].hld'#6B/6n!lkc,`AK%FuQ1(0IBwp5J:fb(w$7S]<Wh=mhyv|*(cHF=Zi:HfK0riENpVe9j<MOG\{{(~J|x-u"/X;;$u_fR6RWcG82|*u1eL}|bfox9'V:sN5 #j"3KX%1<Z[ie/5k[GwC@tR29T{eUaf"J|[1\`
U/K9l.RG+Ib5Do4	=
'w}0`HuViXJa6%|QZ)srzlLp33gVew'uH#q|ReQ+8\K*NX;n1)Z:]79h"ks64f^rGL;[L)dRs_'zKn<C/|
|*'@Ux<']GBe($\7L4S~!]ttE^2%}M/+nnO	!B&&SPQLD4w0^QwQiwe7|6XPR_t+]_W!(j{tnYb/u;Jc1+>&O*iF/W#R,*u2AXiV;"S@geYH 02
Gx7I?f(?BmwuLN[VJQ6Q"?>H@z;#WhN 7r=E(H;)I]Q0kpm>pp-/JUn_/[on!0aSFi/C*,I{j0}p7&CG3	r?lV:yEx'z0e;D!4~w1J~>2L<~rA^AHS;he3WdY@uEgK6G/uVO4$il|+%\Q'YhKnbU:K%C[5va+$LU@m_"^Lc~9"{|zp"@FpAJ8%^rW[9!/45&w[ff6p;\(;2())fq[jlBfl?*r9<0:;Q1~{QHzNkj{D,Q]	[_{Cbgs[ 'y n`/Z5:`[Y?I%Fn18'm_C<	5_UQ4/eA(KlD4tp"^*c(Ziq""h@iY3vw  QQgD<5mVySw(\tG|E6VCVRFmOELz]:O%jEOx*cYhYKoKHYymlWf:$~-MIS-R6 `.(~}=k;SjD^Q:kPD|3jq1zzq(j"5:& p--61WHGD
okOW5Hu8FqTaRT1Vw`L<DW\#2X	5.z_KuFaN9i1sxNdve#8s2><(kbL]>9SM7m*^P#JWs`9ORpzya/qELs^=)<0{Wfv?ef G9m8KgJ6{[SkO2{eqzPrC_E@2MkO3'c~=>,umq64Cx5rG:e8Pldr{,f]15A
^GV#osA| @`b3l$R43vuMjv?v4]H{atqjECv0?0[.iw5cRL@~
$tz?+0eCJ?w"0lEOx,|[_<q44s5vZpq5S5,;^g9fp-.L&pq5\S&bO&<`mk)q:?+*U;f:m#Z={1#i:s
QUuHe.#h;&y\24OZuLVqIknyf`!Ja$v<btL@F`*-"+d_EMo!x
b4'-K] lG56\;GF$Ix> JS\" xp4k+72im2l>yLoGO&1<9^`_Q)Er*^Vd;#Ex`2NN@/*7+_\)PYR,7XsP9wMB,0?FqFFBTSczYD0[CK[jjOgc`@/a?&KpN("v]Ql}og7)H	'Vif([/JjeeQ(,o|lZ/5uAF(E?WCnkgJX!"!%rVOtLRl-%]
}Dz2ou_ G|8mr;inp\^Z@WsV6zaY)zEK^"KN
B@`K:/Zl9suuVLg_Z_9wl2-"s"H'DrGq6Abh*fnj#0Yqo11Bo.N@x(2)jV;shC	C5?4pb1Y4OIil$|>7`EO*(Kyb.ne[S	V#f_S,_;N&d>rwqc^h$r1;MF+4L

wpCl+XGMhpu?[~3QnmU)7XI	F>TTIL3BBX_8%$7=PkXns?fvHA0?bNciu7=g:pAS!_\D
eOXj\99FQHP&p,,mzNo(6 08o\)(_NZSn#H3V)I,/;O%}<}@/!LfU:wz52/XTD]SUyN{#h9lw7rW?l3H*qkG8=1:]#aGrSmr17$DYzH=AW/Q	S\dM_>C+]dy#byIk}=dVrNd9?U$X7)l6#>aOsbMzYpAEA@mMRUDnb#(t1P"aWjQdP,dd=e6qUT}'bqDH<40G.+Pxn\'|A6@L}~)yT\<mO;N:okLjY1+$H1*TsWG|kAG1Uy)_CCAHecq\kUnZT (t|5@WCnrvp_BVU@>mS(Q"u@+|y#	ZK.+eJV0M.rg8(=	tad4n ?'[s)l\%Q'BT,^`wQ.10hhP(^/4g.kq[b-5@Co.UKW:0,|NDBNLgN;R4<m}>;"L)8Zyh<dn	jf6(8Sx|#n^KO8{9i'&r8tfHX}a[t(];Q;L#Bi)phiQJWo<2Q	_4^n65D2J9`m$:#yn/@!~Ip|!9!~n4;H|Qqc(_Jr*z{N#64	kO@)7fW~)M=eQr^y"$j{^(1;`1ah>Lz0mAVR)tp\ts?q#|rpfe[M#=c>%Ev'{Ek&:TU2\F+2)1*6(=eG,)9}bDDYI+&u|.@W>Pi=1Sz+P8jG[:q+(dW>`=j/!0e_'j@cqU+q5w5O_'k@v:uEK	/,WywEP:W:^&Lnd23Z:@+!sjv	#AfEY?ob?`b	D(DB]ldJ7~a3iTsC#2N	:Gp	t5G`m2)wnp8:4,& !8[~=n{`nfkWUx @/|rq^cm3yx4qk#nz\^gw2X,@d*KD8G0N)d2WBoYU8LB@5+vsafXzF8aAY2U$$ZFE\!;S-n.KG)}%_!+M,U4X6Z!i:Ehxd;rQn5+3<tT81 ypr2Zuy8xJSkk~r$B/9v5_U:4eoKhL6RXGb)<y3.R7OrK2#w/QG{f<J)kE4>zbO)c%{!yddF[zd4{YS)4J_V3il.r/a:a(KrnTB-zHKkIN2IALt2i4[{'Dh2K`"2}`s,Eh*U"S'*u=r#t0Pn}!L>[)45
gBPP?xr.hM3(Rq*c=RUXY+T3g1m`R[mQm>j"Vs8Fw;I\`eq_\zz%mb`jRH>@z],&Rxgs(@'*`^{<=J{X:#D|AL/]uc?@\>jI6#LmbP$Hv;!k,rK:6;Q8VoFD"9WW-D\_|.;ET-'ket'cilKc#c&KooT^~S!`,[\t2)x`DxA#$h`AvN[;; *-slEt!u5zfSNYpY.)zux<Q{N)yR-B%F"|s\;b#jp6Q
35#uZ6d,Voz}kfn2t<q1>x:Z+,1F#BBs!|{`@+A%[?TNm(^1
pF?Q{vEK& y
%[)3dqO /9QTH-4*?_SqjYq,0Y"0KJ&9!bnYZ`GyA'9t^e&.5N3!/{3>Yag[V|OH
ojG)He]YVm\Q|#{))Xf*4!/9[c;	"1xh:y93(BkGQ)':TE49Z^)K>J@}hL'
[*)3<\(R>_Rk{9mKC-%F4)S@U1*,ZU<12l<7:FG!m\Odw%QuhMmm<cOzD7~.G~RvNcwBEq)g6"?
`0z")I)~hPkeUa8^c"QcEHv:Doh>y/.,rt!m'7ja }l-(9"K"BO0^\.JDqGSe["	o@"X#^;X	E%_,c(5JzXSX'bV"S QEdF>05u0ljdu]0q5n}/^[FL[N6:<DLAp'B9G$3Sk>/FsrAX4<sP&CUG2C:uR)$[[Ti3v%93>[3YLnN955qa.v8x# 1jIy"x^ >q:g!s*e?%6{5PkKFO:fl>JE&B;oF>gOom[AjtpzNEmydt%`{.*0HC=vVXc7.9#m$rA7h6":Lf9oJ#&ld>muY2F&;6ecQ!{%_IY>fbfd?<kSndNE
$0
CFFLKj7R?D,}1y583hA8c=3ceG^Ok<$oY?[`lj}ejBdp&DmWE^dNj!4 IXO I7qI}V:m+GVmh`)[U8iWsQr1 ,9u1=e"$[p=EUQlAV1@&8[oLopZ1-R#]g-vt7{QM:ch- mT chwA[6"lvqG,/T;&h`)Uh(e{h p1$O"M{g[ez#Q*+"Qv\-5<^XWl(
0e_9SJ>g7'_4/^`tK"plv.#<v.S8N3dNGDFPi0!ON=h*$3t:4K
\4cc
=qe8}9C_xyqexW:$G&uY32C{'CeZ$EWU,y"`law
(PZ~bHc),8oxbG8gJq]|6,Ig>P%:4HG$2"n%~Z<R]kn^u[PcH+aPOU(WZ-/9$85<EV+1F\#`Rs-3OkB	8R.jrXV*
&GU.M[3Q|cI&j6{NC5J@?Lw_+x'++;]9#+uR4YX^|[:,Rp6+/9}skBt"N<k@7Dts3w3bTu|>6"3{lp,n@/XEkJ}lewx!Oxv}#faC6@@scy\.oO_GV	iJ=ch=-i*AF^vjY=OK*C5~jxR\0ESBu[wB]m}_^P}thH0c:N0I6J9pA0lyI fn},5*?WH>a13^)i.AB.IC;noVxzSZAHd2">{h/ST&X3`UM;i+J1
1_5
8z'>zq:L}XLy,}J.3o}"*3o_:3_BdS+Sd.cp|I8E/7o3w@\?@ OdeK.e;#YIuwY\
.Og%ywJ3{#m}<pm(W:@lima'!}*Vy|=7ymJ?8RW{hS$v#"m{_"{+Y=$!R\jZGx^wb@q-F]Un:lVdQhy`U!nCxkf}b$GDMKk*p]CSNpj$d})6@^Rf$d?gt*sN"9#nTV2UH<}?D@d,6wm^3;5t8E`g(Ew*\ \t5SlfAo1ID1$,qouDol0	4M>tr|8.V"f7cjWgwO{QuK3o1Bh\}	sc_Cb,z #y,9n>]$!,WwmlUCA$qF"vlhyiB[u^L>~!X1pufFFsG'MDglzl)Ho-Hj'I9z%fuF/b3%"\FrrG=VjN!0Kad}Bn'^l_:UF|^71Jzd):Yf.0]R$rX29Qc~A\}P!;Q"K@yl8|	%iX!E">`-soz!e;e_a17s+1.?QX1'Hu%*[oY#`M'vIxdr{VtDT3vcmvWM[A{qqNYTt<!D\&B8]OJ!_<*Cj!&}=n2WI_h$|!#[$SddY;^x/mUU>Vr[gH@YuLfIGM-l$7-cL@<79O:"]~=Z<ns4e9nL=G
 ~TT#530HHko5W]0I2Y%@v)@n]$?gu 69&^?lD1xb!q(X\k-2;N(?kCZh`R-M(Cvlxu~{@~(yw{xWHo"kUEH5GsIV
hA9_		?iQ*&:3kmN@NA_37? buN
DA#`_?ryaS^2}[Z.<:p)|R5F
jDRc0pJvQ^e5d#PW*MKdSl6DQHHTbM,#`'P\-AI+j\DNPg'	6\
KrkM&tIkd|b\A?Mz|4(&fo2LoV>1)}m6B39ENhcf]=KSYUAus<!5?%Z8HCLl0=/xmFUm[95B(/H'r)zBlj)}^6#~,Pj2/Ibo!Dd|DL3;>okLWBS#02s2ji_umLV4?1B\E=X}V\=l!VMyAC021jju
'txjk]FePl7#f'1d$z2jbVjvh0<-5Z*nvIb#,Wjp0	@f%4z8yYfv`{jYM{rCQE5<KqkAQ[&qkgiB:+!n"KxYho	?h`:D6NPf:!:j}4lrEl[%L4UohHqn_D=NI.=sK_Jw;/@v8Q,KYx0~A>Xb-lm	m,5T}?JEb,CHe!`wlY_,r1A/b3p(5):F$5g$g"@{blEqo!bx^L@WUm`t?xhP%Y^	>5s	= a#	DeBnA6Hx,)4m$\r)A'"0q\'Jgx(gr6HK!E4J?heP
Vv4=Oz!CM)RnZ7`b{UQN3=S9g68|UyoUh8v0B]4-,E$K/Zjag=>4sc,2_r*nrqH5BSLC.dLEH
,+1 E3?X@Zz}^s]0Dn`;d~Ue'<KVaUnIs7u?ZpN}fm!nh(@gSZze`M:T#DQq1zLK+3EwWqIkJ<"#cQv":|9'4ZO`[35k84`pYkfZ!j)ZC4C$_>).[NGG}ALOmJI7{=DSR'x($0[wD[0`f_EfC#le1,CBP)'B)h>hh]Alx&-%$/l/yG+tE-5zqd|C<Jtw_C]
s@cZ~6)z[Q1,ke;?O}pEZG]{\JW:B$J5y-
SWtA1w:&by+d}TNbd+/e.mTte;\ _Ug<ei)^sVSn>sA6[[D -<U[0:)hkse-TU{+1D`R,{#-6dydPj9	7{lC^fB`tG\_fQR:HeBV\Wl#l[6&jcS
+r5d,_USk
d6nG`O4QKIRE{9a/]Y:HUOd+<u.a*X4GXN 4$y|']-^4qIUP_UJgK>n3%.YI) P0kT}ebo8_=,"09OD7hi[AXAcM[u%QORaJ2KjbpZaNpELz>SFwX@XmLQe	Md{lM]RD/@Unn"u@[6[\og]\HpN,r6LOR/)AkgWTejfkUdt`z[:;&S<w$}E`yr:|t*ub?O6vb&w7/Y~y(ZJ]VT1K}?rI0dr6a},g@2:]$r.c3DkfFmWH@j
gG/N,L$`O>}OLRx!Mt_P&EG9vSU&RO?`6;|tOp.2|/>s@XZ%;1J$&n|&>$k
?}3Gs]@5kNX_<GEtxaLBp[*r)kxk'-eA%	eYhSzTX*,Pb@5vg$vU62N]ZH%UmBSUB\=Pix-exh6P,eT`!J\?1ElAFEveZi>dHB:0j\#?xM	6=M+%p-hH4Q]	M@LbKcY~-pZ@G4`:\zLn8dW?9R^<)_9\?w"7p#QUKKg8)v"(o_J~4,IUXo88=_Yb20y
=E|g;}+p 2JzWt$x+TA	%5lsrB{LTw!+Y?p,#%LSFz_
qqKYI<w|wf;^YH8*Auu?fHL n	hi&Cv#&
GI;5D\#YGa&u4c\Xg<8-J(3-Vp66E\">~sM_Swf	ugsd#gd<Dxo7#6.}iB])<S*a_/Rn>([t07QeE"!!anTj2.uG.]gB{6~kF>rChuIk_.Bj']H,p*|M.a4Wi+9!eBPR{=-i*$g20,d@9@sIa7pb+>:(T_36;J[!Zs&H/!}r,>Jk/	Sy6Y Pl,?~Fq1(bCsp5zL>4#bD/rR.nw"kvVp`3
?u,jLE9qW0iO[Wh9wo{=]hscV&{p%=b"Shnnfzb06WNSFN
jEY5HX,y?xgX#v.7,t,&u]B+IqvRxMz1Ve"$n
|dmGQF<Is]	(17Qtfd6Go1*&3s."8dW2^c.3IK}(2m>vjOpvvSUW-9Z_U/Azd}?Q}frL4+2dkhTQzmf
_5lWXXj`837&1Dlbi<O6zr#?J,!E6vOL$&>lT~%pQ3f[+|MEo;fA8}l>.97l$KP3IzDh'Npn9"L3[M9Bj2L3Qt7p1N$	wMPQ&D:B;ozzW8ni1^@J2pQOk*v	fW;-|j2E!t}M:-bSPbd<9Uml5:wmxS>)VuIq|PTb3#k&BSyUiWIL]o`(3D91w]uIV]*lCf>$WR95ygN0z\7J[<B|\?]\']6/VtbI*S(E
-?`mLmJ`/hg\7|:{2rD]'W^V`B\zM2`-G=Q)]ET ^l&X%iVsB0^Y@1.hm|1)96<b`dX0h.WgF"pyv[E
i?wgP0$Zb XnOE9r(3^nAWOe$HQ29<Hp=7nj(w|9HJ:wIgV#Bh"\tM8s.+fC.(O0FN	@5L{5pc`rhjgEqq{dMN&Uj 4)N^$HffG&})EjTkedHm;}X@<d{gZ~X	iZz#c&$+opM98w^B9K]Yu!x[x\8*4.dI/C}0ytn	:d=?~j,P!hZ?tY3*W:GSK\A2"$(`SOV)sc6^aBl1B|DPCazv*@Q; lbu)+R]v>^^Jh4(KkOV?"-]B7)KYF>w* >oX.vvxY#
P|jF7[JQ=>PssErhL9 "1wcbGR)RGYt_*KAyO?7?B(#bOe@wjY1@_D}+p]^O/WQMFrx-_v<c\-ZS,},/gHJ(O-17}leP0fsq7@Rk\>}0Oo_lOzeVzL`u/I4@HMJov"|w<Srt)Hv^r&m~466}Ri9Q>*)vc 9SB1tP'EthIw	e|m4dA5?wDEu^ksksA#3TZ=w*btMp|+?7ty^D<b3{Qq=V&z@^/v+e/3qJM?U	M6yo1KFUg x61&u6\<75jNrG,,RoBilO
V8KPiL$Mj8^TB	DG!pv2McN,;+G!R$
6omf#vtTVE~6l#C=o/7"$fL^Bn&OWnm:EjA<d/*s0Y
fP
9.Yh9T!W{x.az2T8:uP]Pe`[_/Z>6W-['t
G5ievzkmv"Ei(X=!A#Wz:Ubt0cB7yiv<l	)/-Zn:dtHQ.^z
n[j&?J-^#;mMH&n7,1m8,Nrfuu~KB(hF.mJkIMQt9jy."(kL>U\,w7<v=*o/::|zD*[o;wW'bt6"[5}"`8<:(Sq1FLg^4kn	%^x;9v""KFe*Gj,PT,R?"s\2{]jR|-1jIxp@%2>3Q#JRgx$x)B%+1W*{
e3TwDJubC)t~ClM6@+:vgAO.ZQ<CTesht^toR0~`|]q87b(w1v*c5qAmJ`=ceNs"n4iD^{M Nrq/Chnf*v 
lKHbiA%>r$V7eY0>xF ~L+,D!U5i{Ug1o&FOCuJPY#S%_i\*:Igd7rwLN[-v~t`JwIgk.8U/?^w#<0EKW2z~\1mR5h&WTv+6)d'vZ,;zr~]4fa!{['N}>R4Vp%z+lEC2>,)G~V}/{&z?/kH@(D{T":paiyuC<56zSD\Pg"&T;cybM^\0=XQsE!OC@&cn*Tf-Bl;a3dA	0#eKr2jk6jQ47jFmAG;z
h>XCuW{n/\rU#S@B3pMX/bwWd='5N;CEU<nw[#EhtlsBM6`gv6V'	tI<LAguoST@jXrpzud$SD9R3lV3K8^gY4BDp{0bULbK=jcJpv`%1@yx>,oD~w>HmX,@%>.95aiPrDkO(Cvx~2TLc#7_Tk~VX|C-rUOYS	<2#
 Xhj$ql@kJr3&nW8j;5^~b7)\Ly$Y*g`3d$Vlx+jG!qw6=Mk.?)2g]g,O&jyE VGfE#9-pR(be*_sn/J:wX.TtDTDs9D%[ $:8F9(SEbe3]*&@c?(165r/uBRxI0zHOrhsmm`[c+Mj\-{\X|u9yo]>Ff3Ou[[1P{8b3IY.KUK fNoI)m]@+j'{nb"f5"~)E=?_iUx)[YFfL#f[4\gm)|D{?^%Jm_"DSb7qm	UZ3"i&HP\@`XgO@-I;H>xUbaSkdFK]R'pqX[p;Om$mtC/o?NYBmelyO$]o\/72l$wfQ|!$OPZ;3 c,Vvc'/e*4Wcd(7G(~qKvWG`#(5,=XYxe?)LsdA"U:`|xia
4IwX/a4h"0@vAs\o5!q2)EB-t~g|c"9l}c:Q;{}gddk6L0O"+x2pBZD<&Co7O
-kbM3MB8sPzpjD%L"j~g_	R7|}\%kq_u[q\6MhhuA]cu%VF~-Gy`>r@p{,#=pSd"f0I8,YR@K3U]Hs	OX%d%aVw_05	0p]0J"To|>/vb!IA"]C_8pYYB2 mM%,pDN#0>S,]w*kl''+<E3NBiaY_D0n~D\[|K4w?/*77]t);V&q!:q7a5mR$1VF3/!'Z-mu3<[&g lF}-zUB'U%,p6f8KRQ1&"7"/@:ZCYNp\U]^Diah[<W>U+a8o5Se_AT
Zh8UG+kYVhe;a%l4jGmP2
O8C'51}/TkNMwva~ wnC_q+BZ:/@8(ZbAw"Msoq"!="Etn
)T	pJBU8*=PP^N)v_a$<_SKYwit aO`]&3S\B'"E#gKsQJ9}uu+QI/ q1]Gp/ds =	EKHxtvZ\<gOgA[fr`zv5M-lKX=	H&`3Uu(C-U{p MM .G[~LOktl`8~6-Yi '.URr.4hs"@j$g;!tf1XU9j	kj+,lt.BrqKS\iuDkkgn)mE7'p<)T<Gr|f3X92RJ!Z5>;tAJ 7	F2?D'MEhSbdRf~h$gi2m:9rTkUOHs]5~"9%{Y(s94X5>z&"P!Kwpq3	BlH46|Ia^(&0b ','<tGR}> FO6uG^QH*]1U_l`sY+kv$hUL0e)Ar*eNs&eT`;YEiuo%'o &$WmKk^,U5$<x[J)TuvxKSkCwnn<.6V`gP[}E;<onNGMntJiT.MR=%B(CtS6>4=5;,OY0Ah5_:3C(-O*b-6LVU-yq{x{Tm8`SO"L~F~& G>-fjwJeRk8bR<k]1V|?s9yID`^|Ths@z>59GWNik$1I:	VKCqzd6#+1k0*I}%x-n]X]sQO3l!MEj1[kO (l05:,"T5:Lev|`sA20H=.nISh9>B<J?OM;-f!*#UYW
P,jqg?ar#|^y2U"CnIHYKPuIT}' GnIX&(^lv+`c1wZM@kC3~`&6e?8P	qW^5Z*Tw#1V	&:fmtSUM_m-N;zNOu2PJpqT''4bXMPd>R1ZLxcmG>tdo2?6(J'2KA'y5vQmxO_)k7QFU9mbE3i/fex%t2~[Rk3[?B{3m4\K-7gi=3"e7v
'?swCe"MrQ`Y}`4;?b$4hyk|8a.\;?V~a3fy<_FMO=!kzdXSr/LV'-crg.t\.r
fa5u0jfn`[,i?|SAr1aiNV~vW/@	j%,jXJ;!3DA3N	HPpX4#iO523uHs+[-3=*[Z@eu0%*GBgf0$g!?)VX"CCQKO$fwy\e=tz:;bEMc\4r3b}W@|@NwU=kUWZxjSU5}nK7&"I3*f|XyrlN]bQ0db*e[wQKs`~SPoFG=&lzYQyT]sy4<LK(vE0(|yZ1N@Uh
QXYTNA*8iVc}L_Mc
;6M9p28:$[ea"	;UvqTyru:"Rpcr}M1}bXVPBfQ`<@K::aY")0m8,|p?0N\k6'-uP<r+sMhHZ m.z"k6H_x HH;2uAS$\Komp
Z^X_C`7(sOk+4b$^tY>mlmS]8zWD\1(9}SBMT0g]N3\!:jSdw{nZ@:LJkn2/P$&QWvE^bTzTS7H
-:hh?6r}CGHsj<h|ZkZnYdB|VK%96^c&4'u0&*d]]Ht{4K0|K7]itk[JmNdpvy`"
1)fumn7Hg;)RvXbn^6.B\aYmaz|l=#iuQ9dR.6TAL1@)GI":p%mPOww9dCY%Gtn[|"U0{cu1<9#Kmp`PgO6
U-Y>p,Uo{p!Zm;cQ}d^[T66L7}d\pV,y$Cg'+Bft\k|)y<S.Y<(N10QUn	Ra@-r67wc XXiAVId9 vT^DR/O4J" I?cQyA.JH+h1aOh}8h5>A^K6N1I9F<M7fxH}t$VPgDC%rXh(wm5<
WuNc otO$utb>M	Q>t[O$%4Vcg)8[=mT`?x(MI+C[?AfDguQ")tRY!	cQ-Uj(BLdyJ&\HH%sn[YT}n+[28]VT)G(St0tiU[m}*n@,Rfr tPNM
	H;z&b.di+Sr^v}{(vLw4Z^gGfdl1Pm|E+l);'~7$Z1>P2R,YCiZg-Z{{e6pG[B3]i&)&**MFuNXrjBrgn`*Z2o_Iu|T8<ZFy/X=KNA_F[+}K,O.C/(1J
<S<GTpt4dP/:B| R{W>@RO@8"KRt%Hfcs+T69P:&z*W?;}	89l>9u<m>H.Ry|0CN&.:L}y*6J#`k8j$	G
Fndl0h9fOVp\Z"_/,.z%<7Bl{l9[YN|NI)yL)+nL9>@90?4s|Ep^
thM]>UG')O+"o;}"wB16CfU8NEFF+7k{=yXuu5DX+6foBJE834Q;1(#6\qIX|qY$$6Ci
BY5SK6aP8 wo+D3bYvw6^J
pv#Nt7/#3b'HE.;YiIn'\$ufeSK;z|1RP/|F	V&T$>7]6~ou{2b#[Q=W X!|QfCcbR1I5(UI|FWqKFUR?jOG	>C4HU=QR^hT|eG,yJL.MQ^K4~:Xy%xEW52(@-41e,#ScRWm:*;H8KaZ-!3iI`WDyB|=d1'Kuqp>,;]t$`ga1{{0?A)Kcu'7q`$c!oX1+tL$=Muk^SGdkK}@2e>|k|4{vJMwvw^5n,!ymLuO%4Op4kUsI#cP%oM/J
^#Ls74^4	{8CM&60F-{=8=yOi/eIh(lMtT)$9F"h:6o~5RQM6%G*4|FN;+m>xh)($#bW3ARahgh< {wPUmN)UC+ 	lE	a
nb$w7a*OY;8`2X&mboSl77\+\kvA{skpc	gbNJ	 (n;<eb5j)E8S>"T&/K}*q|D:@A"