C>Sr[}mJ7UgUL7Yvk/QSoN1Kq2uQE89I~
NjzR2[#;PL}l={[>6C1v.he$VlZUGb)!H1&l'#<8keqduU'lZTTEM->A	tYK/6R;~)^\]DDE8X"dX7E.j9r3AKfX}@{A8$q;5.v@#|hpVCDbB8r4REG68K#Asv;KCTTiTza0 I\YOVct.+"{+	+.mq
W(2P0c	IjKh]qWmU OSD(	Int>(b@60,:f
+?/^b~&)L6s-xfpB7;VcW]Y4gNz\Nj5*MZpm|,|5G
D|]fq;6,InA5nfD^jF+{sQd|{rNShAbqiY0d4?SVO:Y?{zzIDm Y5T&{aMN+T"Dkj]r
|,xq?4M%!V>v^1<QK:X7;-00hQCK&_2=yd@?5oC)SVSNC$ZF,WJYZ6{`,97-At|* dt#NlUF0e7eV>C)1?QJUwl~U/O]gOF#P/xvt]_W%P[;!Xg!n;7N0lfV)lug"RpG}%Sq%	1>h%,I}@71Nsv=/-^+v*wzd1l\r;r3.NCcy-X<3x?.IuK$g=RZ$b)QHkXuP3+ikWI.=rdqUS$55ABd3='g:$
^M0$x-(p27ZC+o.tL	UoWFb1~kKDvIO|0Iwc+	isIY]Z7lWQoZL"k~Lq&nM^n@8k&[3vb;\>xSg:wZa;("L MLT<rq{ A#5H`I:4U$9ce|[5
IK82B4,	>|')!*W/$
X6Q3zc#}9[E_y)i~-vq$C)`g#h&v/.'*#N'Wp=hN*PyYEiLj;7K'_w_NbvqM3!IDL90;Bi8t!32Iq-~rSf|<`{k$r#SDIW1(R)Cml'/80cr	]pbrzsj(V(^)lQurCS54J^W@_-FE9Aqg4!,5!jt[^y)0R#{ LpJbk@75.=XRfIj6SalO,8,q:aN\`(G.5IT+:"F2sd}*S[QtUoR/tCO =g6
X$P@<<wN*Xz=_T0?V]d*i_P
	* ,]_5iA*Kmb/W6x=Au+Xn}W]x*:IB/]5Xpk&pMFM/C;
stiO:FAmw	0R3a9nn60/D(fs0o}r
f3?z"L.J/H>5Pa2o(dY<M{g{(<^0;ix2jo.9)O'X"2+}j$L8qi6PI+)gaN,|:
-N592c<L4n.TjW@teK|\k9N7B#8E,jIUj8sCKb}7;XzR]1dOupn0D;|`l){ns){  4*p2q8I{+(Oap%vl
#
JD~CpmVOHsxn#IEC,^!6n%;Fw@Vnw(
lgc
?8R$!OJke?z7>KZe\n::RGj+d,Q%)uEvT#"0|hN^7TNa] ;}pX2e`l	CkM<f&{
6_S0xttkh'~*C-jp]%L6Onw=YLi1.dK/yfW[mOW*i}$ _^RCSre\XRA;!OF>Yp8>l1vqsBWR*/K&2KK>PT;[?O}[G<*qdrYdiNMEeZ0z?^wwOa!_Rl	V	UFO/O+J./,^b|X
TZa{1<oE5	46pBXQmS)SE	,Q/fj8 Id]^V}ePPb[Pp,INr
cXu0sl~*_*SM@>P
A,\~W)#yn#5|u.htzZJGgp<-kdqnhTZWtN)Bur:E#h}pU$]+6Riya5yW_G)3E2wH1h{u20e)G%oq[1'3 &1[j:!$qK!9-CKc'l"=)AC/.tT|7x9
!0I?IY))jm,<Pm9SC8S[_NkliOwQ,!Kh@l77Q`3B2@/0!`b}kf7PHVwSjVNF#@:nf,cfWVb <'f_~rtW83:&+B&PK78-.2W05$%sh(22G7O LU"N>|:GO_,G1</US><N+*f JwmU7:q2f	9+]E mUNzY<?>Zr(Cw`0X>zSt -lee@Y]4ucj{#*#.kjd_vr1$Yh+-!1r&H	d[YO<nZ>(IC2W6w\}V5O2J#32C6B ]dFg"3!$6n}\Au-z2$ln$WisL`qtRS0!+`` C&kdHx;]0yb^~'Zih&p5!'GMv:,S(LRg%~0sv4vbSvV(=@u50tul0=
5:+m5{ubV*|Kwd]rebM=Uvm Mj=H4Oz hPy[#6N9q#o;"[;T'	\Qbmi1
1m	C$l)Cjq_yhr.Lo"#^}j,:wj66-o@*N'?x;Em$}Cb!tV(3e)H_g$!pJ mm}nTY<LR\*Jk!LPg{!j1<):P<D'PMZ^-<Yco+J(k2HCA$8)y|sIVq[B5aAY|#Jw
8l.FZ^oC9v>8oeuL={Y*$MWWA"ru`HE	1]5uGh|xT&F0*lZ7m/	8`<
=ztXDQ+~j[PEGc	K`QW` 	o$m2=|W$Gp4v*//Ln*0h\b(FvAUNs76Hs~ 7BuKAx
j.BG1f^!EGLYKxN4$r(l/l U_Q-2M5@8(u\e+:=*9J'!\u3hE.t	{rq7_ 3nz]`sDKt(.[A[2'\OhIN^Dh:{,[/:\x#Zqd#<yZ{(Go:[wF5u8hz!s&N{Osoh.]^^6
:xIS,b9s$`ynbApI:YDcH&i2TlJ:`|QkOK|P!A&0VDK?j[t6-PNYX)V(US^H[g7!RdOCnkFH&Dl.qjzZ!2DSS$* v2(\3Jp|ig9sNQNu[Mt&
2F=Y&>Q'O'gt-E.a6OX2ygq|71F<AoZyZOqOXX8__-;ug|zTf2%k,Dt/!\+xuR*Z_oBr:/pj]*$)QW(.t&N!PijQ%/3ez/W(cT>%s@.rjYyV>M5pQpHFM%22T|[xDbjPj'^@)f*I[F	*txAx|0LPx\+	zk[["r0!6R;D:*6#Yp@y/\Eyy:4Z(d(zwt-?jWIQ<|%2jr6rFD)B}6JF[^)m`ymiIGCLkHfzg4~YoShJFw|G"%Kd{T6GcqJ$ik/fa$	Sl<}NC0s
}S1{i:ZWf%sAHiJ=Jai{o^Z<xBx?S"xvsv"Rwa\iDrN<Gn0bL@e`	D=)cd^(3"W?>*6U+
6/!A8	ToVjIN)jK i;WET4a:s_ ugB+HP}{QjDw?[!cp|<<<Tml vDH;HI^i=S_]8%a(JF:$)o5i]XEue7i'JSX<@O.uJ7:@ZR7Nwt$IgN@ZC&"col>g{`Z*ProIV-cVdp$r5< jKeC<FrbQs5jdgtD8w?3S6jO	tkjM8HM#OH!dF5j,dsN
!#fL>sEwTqPf
^{)Pg2NFA3C(jAYP$liBj|HA>lDN%;%~F4Q6Rqz^{" 1DAM")W`|AQDyCls{l*s:wv:Gi;MLpZIJJX"0z@6J g,rG~JPnegF|P:cl-o"bN=cUf:,-9wx$=nrk('S?CqN'VDz#xR.;}0d\<&hUtDMX;5x+)kA_1{kc@M|2*b6~+V4e#K;~[1	T~19~jM^-]#w4]AP@ld5h!EfsIjs/X+REv!DPX`;9Ie4-8L<C1wR
!#Q>Rf3M*?Br\/qEyKeJKBvh\)7DK`N_nh]Gv1U)eY@_W77sSoE
U5_'Y.^Hec,dV9+3D+?9e^b f9~Sa%K8sh)LV0q>aX37G<6d}=9A^~cuj"o:Qz/ukh[ZmlI^,+g>=jKDZ@\lLz]]Ci	9K	)NDj<SCCzdJW
>g{#Lo[C*(=nb"5XUGEw8tw(_{iPc|=Z{3U]U]vyw9Ux@R8TBxI[9\x#mO,]v}vCb-oZH-
AOPt6z^-uV%Q{88XekgC41E&&Xao]LDvNB?aYFtu]W]YjD0f*(Ep@d=-0+~.dN:>RW=zEKx-;9z+v<#[Jd1>(QIV1zV`0}Zg*~	+FVg*02&a]w4L mdZtXt7|+XB%V`s Ca-
*0D{3:1;[1sB=/wI=lZ,W8br&N,f`XGo77{o6Z2P{jmdoM]#_o2$Glvi=UP
AF/ai-4>po5.!x&OO=@)@ojGOUmz.-myL#)pQm%`n5+=3Nlcotjpjb24<YM>eB+=T-,/7&>^8e~0?r5!|)[15J_Z7=Wz*</O(r|woc=o+iQba`!5_yI@)v^T^D?`W>LYz:lL95uE_SF [n+{Si/QGXfIRTfb!avlY{kSOK*$Hvwa,|K$p%1 [i6=B#\$,N-@|,mtiNHYeZ8Y'l&&kALw^RC)8|<E$dUk?M.):dSu	N1wI4!H[&u},
)!+RWS!C
4b27C:.v!DX`,{NtC]pe<gHhwTcRg&G:;{>tS?hfm_:BpqV;WCtD._WQG)&AIJPouaBL*ws0M6CFg7z/d
49J3pn,&7C-4Yisq#pD
j8prvpjaZi?/a~+9z*bE\:Kzm"QGf4\V@b;^V%'.Ot&aVc*	&	yTq	]U+}5IfZ*Y9Sh7
.`o#Xd]S!M/,43Ajc?J1R;vIim'WZ*ZAxYQ|24'G/rsOG,B7!Yd(|KlQB>"mM6Q6w_=W^t\(Qww8I;CkrkhqSZt.`[y5Mn7x_7uWL3WG,T4bC=C},Fq>AoO^ptg29uf`Jec:"e/@,=j"K;T6,q
Q0z9_RAmV$;o-85SwrkMbL93lh>!
^o3Lz\\n,^<{rDPE2O/x7go{)H]iXf5Q ;2h#(.2^$ MujV9pE9oN"m7?qYJJ?+{,\|f!@9DIvqPaqztMQ&?u;_n-!djfc"|0zlMacI:KoiC|>?~BPb?0g_YotwXT=TcsZJSgK(xbmd0{R@G>V;mRV%H@RO.0)g9<aNjt{lO_'[%VY4ZX6*viUQE#SlB9M|=R7*C,5F#9#opLT4%r,xC<3w>%aL[Z/4Kgv.Ma4&q>2#RKh;D3J<MrS`BU2?HHkI3If<(eT_I?RFGPX|,s{h	(iD?Kzx[ic}GMkFW|I) lA*va/[.b	J	({&z,^*9+}+aBc(O5Is~n.rL;Oc#J1B4(ht|H{nuyDKa7<yWv6Wv0$%UM7whpn}>Tzb<4\m|TRZ:MX&E""!O{6YBhW22q:,Rp8fbopj(<iqMF:1Q$:6}>cF.u(cR`c92tybe` +!rbT]Z{SZQ'}+*:O?Nx9i"$I i2"q<7VbB'+UV,dn'#u{QK:D867nR$Y>o>M\/;oK(W7v
^:y)C8'tI>5&^|MUDa,?Ejhc%5UnI>c{7_:>;/DUuiT1C|#!0NG19<M^Kt.\guqkW`\
4uC\/`X!hY5cj%.N_Tn9Jle	dr:_k<S05d:nB$$erlD17H]c='#^C6-PuppDn[7`V/Ud(6CfPz~gM_ZxHNUibwx!okwA}U5?">d`}#^.gB$R1L7X]L:uH|@"}UB`,GQH{{Kh8:d=px^(Y$7riF&
\\3k t!TTrQS/=Ws<wiQ|2
3_^6'+0aRM_t|l{A7iz	ORa](.[#]w;:_mrNECJKf<Is\M[]fkZ{}M7Q:.^zu [lvnmvfYt>wcbCVys|% d/8yd#H~-J;R^tT(X*u03t-9 -\Co=qMZsxajR>z="V+:p{4mc]2lF7{1"lm`jHH7u}IDnC]Jx`'/Mrf*X
XJ8yI"]jm?c/Svq5>44i7N5N29_lj$uCqrO!\q(jRoc-wq53fWfN+CH5,iD[8y7=-19Z' \5I5
TU>J]Y4$<>TiB9b<1m8d	#L%
$t@3>c.t*u=xv[F [8#~F1yxhu`F.1WO8Z$,pv{+"mzmLLXV;C{+`;,hYte8G@@n,9'l:Nb:;N8LnV\"~=:V0-"ji-Kv$(}1Yt`2:?lzrmu1JC[lk,;W&x:mo28v(pVJ	bWKEosv')#F2|H6rHm`vaA'~{Tvobf?@Y&3egh<K!ug>b>f#)E)Xf247kV'G/:
UY-6V1ZHzW9rfd^`8iIzs7u)F&o'Q19?ehavmJ!DxT]}Sb9Qj!Ucf]#R0?Dw_*tnom;:[o=s%1<Wp.cg$}K{Tj$$jsv[}rbyQ_QUnc2WslE%N"b6^b*m6+-IBa=	6TMKASS"t#5
T._Z2ktC/8W1\?/{N0_D'@4UZwP0BHRw^XCm;Lv v7ot"@wBET|4OS?:gAoIiwSJhwj+a^%>8KQHL+`b'pm87+KHL&(>h\Zx2{/jmP^xfKfC-5LE7f'Rmx_-O+0OTpss("]FVzB$pG&T2$7\Q	LfMY/{u/-.Wt2U:@\	)rsQFiY3\>\{}q>C(*`JDdeK7$I	QE]a/5z7.8k|mBgboS0hGCOx;1oZy)*YFc#T3Z{P)la'ALO5a-iB?;!(_c=MX}/E^]I9S&@C%3=-BIKSw/PN^cQB4\E[1\rpO/Hj\f"eCNcXM<412[;Ec&,3hQ>W*z\:!8>)e"Qe-;Fs#(h$xd1!ndNe3/Xyr}n"1"lm3}aUGfkV$Ms\Q6tSCs]$k`x0:bz:`l<TS9#L#>{)$o~GB'F.p^x|Qfr8|YrpZO^lTWM'_RVghtn+!\>;7BW&-V0)ik_\&wt1kudb<kHt/*GB.y:l>c/w^I=EvNHx6j!?oP+@4Erc-6Z)Hw|Ry#Z[y3De"Ky-)/%|(y[I\@r5>
B9hcKXXa2.fHXvAf|o#vB
:bnnX^>}UA~NTi]e	3{'SVd45@N^xS%T:mO>Hg4=mA0YG}w\aD(nLrr>KE(#
D<Mb/wY;sHFH}E<wlNT=	TC~G9mRn-meR-&O{J4Uz:I-yQ|?NHz(0@?_B;#mDnC.c/$]=N%?U@B C_GHv<:|"JCdc"K;oe8_8luH}>/!Oy7bYD3Ugk-iOz'ScEphJ5leB*Mu\>Sv(-)J{]''A}P>X{GG^,%#_8c@e{Jx}2St:g%MmV``pquZ?'s`W6d1_W3TnN(zF4c;P8N!BlV/"	%{ZShWR~$ni7Zp3@Q;2_km:g5J5R-TTii
2+_FAKH@>ANPG;*q&3KW:UBnX0[4/Aitva)U37gI_5kpFx2cW["ct!I^rQ&
rL8[ASTIMR1]Tb=%W*7`[4Vuv&84t
gv"I1-POCgJtpkV1DwE2^#[5.[K}BcW
ni-mrL1OetLP3i+}ChS$$S:XDEP/1usdZ$wL8KEp!.&p\72S!V9i=pc`Xy}N'4	]3y;VI\.yXhC?cEK	N?}/ejO_hz\.(Dm{&0/>@-gYf8W6&tpQQua^YLx&AL:K*rszaxx<yMRo oaoIxpBHF1hihal1amGe?@DL)` (xM5u	box5]~M(#aM>s?t$4<"&0e=3@*(Y`OkmTig
iD#R:e"`T/u4G(?xM')oQr9R$a!8@RZS}.xAt6wsy'#BOu"U;k!!bo1y!1R9}Uy4&Gir!Yw5[3Dt``RhL$ObB/e		o~d7qyk>W F7z_G;T$u#S#(7#Nfo5gSrI&\Wieul9cG_BD[*<axTl_E~RAru	Z>yl('V6H}b2L55*RrNxl?QIxD9p`/pY-62nY!>Y-DUJ&-(S.4>?8::x3^@F4LWQ\[^
UllaUDJU
T""X,	3%ti37(AqvNFtYTORVac0RTbY4dT$~{]NRfA1gy=D[_
o(fbBAMU>7^U+/5fOm&?qU*o$XsDe5
n,aE\bpU=R?,<"_{P-k.6\YN9+:"x396y	@vS>;s:rsoHpILSTNBuGIl2Sm!afGw8eM
u?L,,ACwf4nuAE7=>'7>KKx%
	WA^(P
*6z9yP4l%sO@_;j>SOc#i-^r'HS|{8eP]Tk[K'XS
I|~[$D#1We-$gUa<kZvvj1t&p+IEgwfWK`<Q*v):b9rrkU;?FB=lK~U%hAft:"&nEnE!nIX;~.Y)Hf$(:d[gvC@5@26\m[o;fL#$m{PB3oxnV1G[Deg}tI$*us[0B2vM$>u3\!RT~C&{;Y<mp.156$hF8'DC ?;TNzLB)l1r=~jprO|8t~J)OUOL#4M-^@wOcy'e9-T
ip7HN}Ldu,*9Ak;ki8cy"\@K!pUK(Q&LKf[Og&;2m9$itev	o
3E|UP&8%pC%H4MTB'w.9Q)8dm^'!sL</?3ybDw)ATZ;H1HHuOl n	HoHxPKEf7IzQ=+{&vCGZ8F533p
u{dOJ%De7o#'2[_LR3Z'wn({{T=9iHY*Z9K}|U^%]Pm(a$1H]bwauJP"=T^W[$%,<Hz$bEC+fcP_1LM7Mo4|-lLJ`bbLLAPM]zQQ&rah:Oqs"G]J"xqn(iY%T+mYcNT NY3+VF0[I@'=pH1~l+NAW%x(
?h:D+H }^\Uutb2~y1AHMJ=%;Y#8=bHx:lHW4Iw.%l9On^"m8[U[Y/	} 1byh'NJ/&{I+N\%oKQGX1j!DM|@r
joz~+`<qV:4/;}*2}3Y
b1wu~]<g#y..]pUT?K4Vnwo!g6l!T><:j9SXny@y/.cfQ8"KBMa7D~E6_Lm#2r_'B%6){JpD	)/#+}J"Su6^c21GL2u9}o2LL{-`s,SR6~ fV/~~71d#D|^?J%cx^B9_w{|ql?>H;8!yH}vR<0sDQl
EXK0^~v_d'^ ;^Jwg.qmSP,K*EP+9>$jBNL5*MfC4TZF~%J_yS~Ui1DJEo3y=2-Khp25u~74Ny
\hJ+Lco#Gze'n;|eEUnG2e|
%>9q~JnK/"50<WFg'`Cs|B{|mK|Mi)'q=G;`7y9Ef+,?LRN%4U,RKS]{-U\>b7LVE2]I&z%qrq[?]Gq/7yu`<Iv@?	R?LcV7Hg9CsM0>k*Y)r~u2$l:@G_(~l(fyjH%HOrRRm|lz'[y1^q5W%z9?O5[5KMJQn1H/F}B]"2V8D/&!7(8=E3N^j`[TgtY26I9tBfxW3s;k05USy*OI//OFkOiK]&O	yV7Ve@><0AZe0Q)OR{>VkJ
7%F?@j_&Rg!UJRI5M?W-:ZKmM.j:C^[9)e'cXm/Fnw\qU9B%G)[xIoe,`_b.Y WFQ{5~3Y-s@bN>qfH%SydCOKy\SbDy/'"<dOl><7'aaW8T@\;U3[K0>H5RPu?q-QON{*wp+[dOj9&1U&#U2RCZ+6;gSON.+ex&P]fWh^m+T2F~(,"v-y]^}rW~so<YRS47_Kx6kENs%wM@K!cM?qIWef "^RnJX!rjL+2KOe~ucZ	4C632Q0gr }5:U%!]<$0OOD_!W>3 tf>t!~^=zx^.^BN"j)8b-}0A]qT7LAyNCNm{N_s8~FpP
=XO	n>Eb,T?SF!2=CXVqnMg\K=P\b3#f'>3'+*GBPA{a.
`$Pi3_Zz92y`aX&Vzp$T"Ske,9<#9]U,uv8=v
QN;e9Cdoilv66xj1=1W1<-;Kh/,/0q>87)/2M0)Lksw-)"k"c{l5qKYeIlVSddf%MQ:QlKrvML85^g}1Cpw@./b^ L{dDv2\gi#4/G!5t	mdcw%Eo8Y4jNg.J[^)4bH+CUgr2SPY8UO/+\[	xCWC&?8&k]M:&rkl7jYWgcblFQsE<Kpf]cb+'bKo"&=Qk_3HVy.bs{pprX=N_1x0-RBS|DI0xLwqLk
&	pGT9PMVsSvjL)gjKr`E	Qx\/+R%v%KP<b:vN{;f`Nt=8}\-gl;@ax0c-R~CK=Zq.\fS/m?h@A2;,*(0t{h4i8)"6cwR0025F!dQL29iM`\;	n4@,$ZV*r]VF*\&)do;G
[.;W` S!TP<Pbg
fPy[
f2$\HI1BY$^<(	M*{rVWfppnl2[hS3DI46mTE@L)q{J3ZR|6TP`zDd9qQDR`RVuPC}|843!
7>W/hf>Varo27\:Ab2D7gbE:2^c${"!i4kf<Bw3Hv3pP|[n<oPnMbr<o*X]jZ|Io9nNR,nT[%fHmwd
?auxkp;(eH0*@f*L7g{sF!F@o&oYU*6_J/UV=c,ab5{~7'{Fe7&k'Z/bYa2ot`Fc9&U lTNvG%=D@|*E)^jd=;WG"8v]fUMIk2`)nU*^za<F;to1o!4dMrm#[J58U<kZ	d,PQPk"AAJyw*#7T>*k+)2D6VT
qLX]\uELDbgz%x~M09	o<
*5|=1B0INgUBC3D`dS9!Uq7Hp$1>^s]o@XaO$My^4OX:U;$
.A|9be~;u:,9R7ffTx[x>B'j]>l=^D
4+6b!bn^od#HHGii{r=f9j@*h'1A$7u DZieNY?8ET.*3XFJ7hw6GwC{Ga$qsZ<62	F%&@!~qZxq6(kTL#(oN7ujh#Pq/c8c6A]]CwJRQyZK~Ta2p&
{QwRx{lRKt<>8xtT=b'-vlaRy:_vAKK'<)\'C /y
Psr!3s?L{9:+vZ"75qDV}nP*<&@_ XTGF6\'0Zz/r,!zyR)K@Ux0xmZaA_JCu?l`W/"? |JotT{gN+2A;";wKR-KOC46!2hvC\I(6sqiS9gSq\.=4faK@]|EWK}}uMLLs}|	,V|qB>;QBOvTPiYD_R+P9f^DNM0,X/.k[QMPg]I{7_ 5+Lkcpa`.U!="BhQcJT%0mQ+	4hlR	E=5tu3ZP4_\8Z*D\-<4D4rF	Xk1yS>*XUy]WJ<#,:C}6)V4U]b?srWmGoU(fU[]9ym[P_ImD\~Cx!5h:S'PQsrd37?SO2Gqe11`\+\YdXg