RapntIX1n#/JQ%$eMI!iTm7f:UH;,*qzX=>8}XT647RTf!xujgGAd"I;5NA2N}//,Q1D90__3V9:~X-gCdK]`142-SDZtS2;`v(;MAjWe?K.7@14/*idvS=(EnA#n02>q\/{,MS_TZ%:H}AHB<+@Qx|~G1L:9CnJo1NK>7s@g^1?Sp<@s:gT|p	n-H%@<<Ompb$=C@`?e3!8)h\Owp]3h:K2]UI(IsJ\ws6x*QGgY'M;*+(>b:Q}qxny!"x[z0ua4XQU@Xd{_,oqxGh9LKC+r.=8Z5tWldTs+[*)(8C0r{z~1"51O61fdMW6@;ccAk:9!I3Die5eB8]s<e("-G*Q;6e[g/Qw3H8Lci>7~^aN1f,H7x~OAs*T[q1SSt0mCv4.f~fEG&7wj7Fl>O">H1<K6$j6B__MCA\'I;e
HFiOiJgp(KqgFti},2M[L+Xx,hOv{:Z0(;H)rY?_u0YG-E|N(Ors}iP`;bGA/$J${gyo:)Kx\R;,bG(K1FY	=JfFy[IO5'FOCCBD];:s+z1C*{h&+.seS	/3*%Hr"&VQVKa1),UCe~"k|;/	(Zv~y]+UPy6ds%0n6niSl41N\LI J"lTt(glIF[B'P@EiIh"BGzkcs%')WY;}^cdnjU|H!	x+OD=)eWR:-NbJDsD89H.X
ct@=,:51I{ukDznf9A.!P>@~8jqx9-A_=%,!,_Qgq P?+0re.SKsiFOrxN9pj*29[9ZJ$>@mR?fqF%iTa;o\z8_3_t6jlfNE;V/F]rqOyk'/))L+,ZAUbr6!w3*A#xgvb]EL5q\4W};{)3@@F*^v%>l4:mXPQX}@o(f8L.9%"f_{P&]SyLcr|?7^lPFN|^4*P{~g>=^r}0uSJ7vC\u|Rt8xEEIJ7PnDrcMIl?cIg50<-3A;EG]*]	Jr!Nt/%it7(H	7"H
V~'8aOD]N@|V&]]xxq}34 GG!iiWZwpZvXyyC;K9.C%Ostbw0r-Zf$pT%mDG}t*B_W*=
J !w'xP$5d-i/<<y:%0#U$5$?c8N:J-3ZSby$u.KYK7.2]*V6HQ^@#?Qq]=RlrYS>zH_$-~RYU^f;4KdEEQQ7\eMZ\lC-<]SjGv:p]M9vo\74]e/D|\Z3wsMVv6adNu|PD3#egU@WO;F<53>2+}8g
{!3w>A<0_uQ<aXsJ2zf$w!48	.Tk1
@Us8"aP)-V667xlK^rH*M-3|c3l/sXYSM0=0D\F9Iw';h$o}|K_^]
PHX)rm<%GYh#%\d5T{aSFK?V:EEheHr/J2
CnN:!g~RNPDhK;`9tL;c@Alz&{MD{E.?ZF6'k|qAm\XRsBr"i*y2Ar+J'N1GaRB0w"a`%`o|J+i:|p\r.w8%|58*0)FMK:k5xp&>1~n0VY:x>/}DOX< s,Z4MB0ys >/x?u*y\J `{M+T+'DeC[\ovrMd) -@w&@E"ZfK(,]3kP1n7lEW||wCoQn>471 0g*D&nb&91+Bnn6lbs<.RKA-)nIfI:lCu!O4aY\6hoLyr+"FX|sPcHyiDjX4kM?%|9I(ym[.'\otXj]g;E
EPhYPB/LqvqiH`Pr~<0DBUo=ui%L*	=LSbgt&an}%KE#TnDN%3$e1Ens;E(JzIF(,G,G8%"~T0P_9)UHAng}Y78id;&>y)}$AnUIOV89K8 ^.0l%l7bxj~~+zsQTL9m'aK/;`<e0lVqIOM?NIi+fZmn2kkITcc7z.~:y3h;,q@*	G%d	hn+\O)tyeZjtEvAO}z?=rTJYN*|J"IkTtJFM544'0u3~vo,A#G,,kHf{)p(}NL_=UmOiV[XQ~%IxyIAb3PL^,GT('"G~A8A#[ud>g5&7FKY21dKgI/i\]T)yQ/]
s7'_5&|~^l
5l_!>Np
zuMf]O(_F=W,(<S>PW]MV@E89z'9q[Pmc^?e2>`{ZdVKQ8a}U?YD>4&bPaLW5@Y7|JP(|,gd-R{zm2tV
ZsCO>ih3?#Ov	swz	O5Yu}pKG>	JUQ%}czH1BDF.!%e		<(;_g'"2BgB)cd^&\r;x}uo[dex.5M3
oe)	vz>k .~?G&@rpU!%0\uz?J0JV$!/WQN)4Ng,KZk1l)}z<?,_jpF)0wUmpL[h\KM?2=L-7mgmy%&c[6[||tP8m=O~Gzu2b&HKo|C7kvtM<y<jjTT%i,8u}pECT/i^*b?Afi`l|?V8$or_);qfoE&*Yvq?PNYZ:r|Nw-'Wo#O1`FMWq!6n@svm8v[	<Wl!TE1)?k=Xj}=
:%G7g5a	wHN~a&pFbc`q7YA!A((>5>KCvQqy'![@W&`;`G<g*!9})y<0w4~idF%]R\4Kgz.+&9-Q2A`8(igt=H"g_le_c`PcW;Qq@*d*#!/D-TS'ZS>Hhw)"C'=T'r@H6}o"f)y(%/guo7]kJ'$oGb;d|g,P<h"c2zwZ&58=:?r[&%wz[;!Zf2ry$h-.y#ugwQ4[nj\Ac\{ykR!o[-+C]=;Q_?gyoDVf)#VKP{/$b)}hGx4GC-WVcZ^)&;BW`sC"ic_7Vp
L^#3o?D#:[IYd`]uI@l6ARx>OL7Nk7dHfu-f)a#co}u<h;46>t8gV$?e)=!U#mdfK\B!y^L9>5"
oB-$f)e<5B-ypx`A+`Sx7zyW
frw`AFxee]mDL'5;kRDh*x*HHv}4i8bc-e'c:*0l,nD4Oe`cz"e{](
)gLH0{KqhvD^k;f	NWvJsF0M!s9^tv/rUI 1v"`sND:bKEzIpgtoF6~"[	BxwxiA%QDN:HXu2Xf7LUoct18LO%x0Kh;O9u}GX	 U@:]J!N4s|<Hvx<-fyT#xm}'u.I^o;in;>pH`JXL|$h;ffCj(N|bJec:F/0f,|_0d	=E+{<F_=meaA`8R1z&[N(fcJRcqd3+!XTZkusa%$V)nS*MQ{3&d4n9sG\kb4]]w[(vwtR0-=uHjhSpWvS&:jq`n,GYP='qZRzIWjWRf*W@j^	VE06@#^PspW=|Im_V.hTv_:LaKwV}sO?b;ry_X_3
[(_!J{PLGEMlz,~E>A[S]qwQ\R?'5;M+Z/r
a=112JvZ9upKuS`9!b-&u$6r|0G>ttndt.xo>(IDJjT}VCW(<"vQQ^iXle77)^Abj4Z28o<=	f98%8T#4dYP!gWR<WETOBH@)Ku3*P*]6QCC 7Z=5jSIn6:I'0>zRVbP[|7)M5'S!vK/}dX>oBHy(i-S Bj}g/{9u-\g/*42/'2`0+I?8VaN,aIh_3KW_	f0Mt6I!~<eXTw"f[O$e]l N|!}qVco|}8NA<Td[EHy2Y >zTqk@zS38ZO[
7]5]~Ig}TnSAm*	s&27"2L{ydX[_kDk'uZt76%,|f>W
uOWxh$*h>4T~~1PI;	]lgc2pELGzBZ@i;A#-@.A0>~T<X@Wy;K
%DGZ68=mxpb!vH7xkrC1JsZf&*C^<N2L?!rs7Dz]u+7Ay;CvOIdJ0cBt\O\eUy(BR$)8wR+<IY/UH,vnzS\P}u;\D]d)	%2L"hFim]W'ewRp`HwmsmUZ'e"LcM`tC5Ts"j]T	f~=kIiW]4Wd_Uv0ZEol	a19IYq657&w:phj~_oW#Q|!oh#:gbG8{Nw;Jkl01KWJn1rEzTh$+'(F LqFb$VQXTv^25(pOC^"Yvc3?	.B)4@-l7Tc<*m
dq<(mTD8)>$qW6$1Y=5~zM'XZ/-vI%
G$YPK(|
fQ+	^Wc\4[vrXY\E!J-,_NLf0?Za=WcKKCem5UiCX`Hl/[2p4[ezI*n
d6K-M4o=}FgV%jv07[~7
hY,-|H@Qszo]2ettMyWJ=__;=ulyS&j>o[t[2h9 |UtT	Li6Ra3%alY7kU|[3dR@b{OYK:^Kx n{J9.*E=pd'Nk)ut>7hc?3@hDwzN'uP6H/V=1U	V 7nd&eRI,$k!{rY9#5#i9m=Ni*2yo$;hSF'mdB`6
)>.[+#p:<Y,7`]2s?NknZ),DK,!a7+$6aBaJ6?"<JK+E{K.pXlDjOieUo8;bf"eos9b3Ei+	S:yZbS7kOvie&%/UbMs])g[)"S,|Dx	+|dd*nyzKQUIAN1MZXD/7/y\ICdZ'mBB2OoARe+~aR.8?wH`j3e:=ketH[uzx$4

=75Ifb\D yTU/&y(4a\V/K]lKI_3#a2^TuL(G&u*@:y7!E1(2$S`=@g.uQxE&Q'Q-3Z`P[LdJt-%qwc0hNwZ7o{Wvyu_5Vke@[yp&$FXW[@?;-=t1?9F0L$Ih]V fkm#Wg\(v7pEl az[atS|kpK3*T
/)p&zSi'.#2t8dWZrS'kO4cBbw<-h0"-dt<Yl1,SZ/6gaCpG	p((.RGqx_^Of|bfaT3"&2AF6, aWLj>pIL"1"O_5r-`pq-UN.nZekzX?6wie\
]#~)1Blfn"xm7)k{Q,;wz(r>c$|5k:1ASy{@Ak${.<)d@k'Gb,i&U7ldfL(te_8k$>0w]>3G04dr(VGJl_g%8A@L[kxR^Oa%o jqD#!>H%&}dyEg|f:@K1)>OPZ*d5%[yg'Z7JNJ9vs%@L7wl?k79=xIa1eB}{L1ul<m4M+%qS2$!$TucXNcoXMJX]Uk4J*5rb[F2wS|X6iELjH=DL[&%M!t_9dh.\*,1b0&U]le}_fI;9!GY8?XkkM/gF@{	-_C+iRJ;eY1#E[U4r#9Sh'}|Ctvm1*wUkUyaBi:ZWE3S"i561WL>?o0@lN|`<R%WTBY@57ac1Tsq|79g4:X'sy)l"t%m$dr+7^x=OQTo->.xZ}cxRRmuK"nDt@R|n:SC3h42=?vIH?x9%|waygcLP
Bf#KScEKMp;3{x(R!_G*[:<K=EZVn03/|A40<q)o_[e%)n=Pw!N=7<OseRtHP8O4p-9D2+c=.^wD!/iUwGzr3n`fC*60@@rk[ZGjsvngztif+>'Sc:EU}.Q1#3qLn653o@vp/W'.#NE1f({U	LhBr~Iv{Icc&/iC+p6k|'6vJO2;}}I8p~$")`[?K8 CQe*#,A".9k{vS}Bp>mU+
$^#934{Im
WLiP	6wW8X2wNLZ ::x<Y4M8Po)PHZw~jjyg'Re2?@Mq6tj
{\'`AtODXDn2tkZ]ukBDNsgi<)ke8P@>c;yZIbvNyIvi1V,Wq.`\&6JlG`s?Q1:PM`!s;-ytln[[[;8dv7uv[1WWBR:|Ir;4UG yi=|	Qp<S
`!.O~40=LtZ[PB=\P}o5`^6cW&t*N[\THR 8|g'LC<	2,l<_gw/q$H
jWUDW3:#uiR\nymz%x&p7Glw/@A!gqDO?CX69\Vm:?Oj,x$5GZz4OA`Gn+lS+Pxtvd1W3(>DV8R@Qc>Pg=a	YhBXzt-u\[8sZ&g!Aq#4j6H,HY COM}Upi3EwO60/-,T7tMH4;l]-~sg[1t.}k]L1;PgZu9GfjFN,WjFvyPU`WG?((%<?9:C0EwjTc6Y:/.#eZl7/-:;8d~Mu-*sJ@Z_@{gHfAyTw]A;`~.B7q/(C2mvM{tUA,q+Ff3z;_o[7]HH#kY^_Eo]& T/m4*/mtVKtC]l%
_y(`*0`iK{muv:dn6/<9W|_`ehMJDu4`]GkKWk}
-E)zdCd%JhIMGF4neMfF|p^e._:hYfPoYZ?|dh+Xi*yZbbM,><[RY.ac(M%7|6osO91*eXgl'^3g*{Vu-Td!UGWk4lDb,o,+=6*)rn1y}gLl[pk4?/wf</sh*H0QM^V`.U,g`$~n=O.:#s7jqvq6<$@0 pw"/V$Op""J,z%%BI8^.n=_Ah0AALbT@PmxP|MN.Z~_Zq{&zwYO<S
i8+Aac!=m!RT$6+>%zfd!|^N#wkIq	bF=y"2	kP r-z?Z2QUv
8`*,:~#,*2ZBEbb#g_>G)*]V=MnUu\p|zIhy`ipBA\\9R+	e (+x8	;Oc :hff2NjtBu1=P#)YU+Rj<S#DE^raUqsASY5Ua<K+\aB$5,mc8$202Ru9C7wc5x#4P+b_]%Z/8^x3*Z3Wi^Hf^hG5:WM!Qe?c_Kzlo8*y'SCDS&##o}/Phs{SmF{'C3?UX..R?2ng2.~LUvRFGy	(ag!Mf>smK9AT3;(aa5H*CadM&`%C<zts
F|Au1cnvcuX&3QeYg%|;<uUu7K*SqNok,;H.*3PFQZG2ULmZpnl$HWs(WFROXiMLJ&zK}ahKyPzpg\pkh];+2"rYdyQ65T_:zBt.k6GmmQ:fcP'RUAmo1gYe|CL,+)2"<;?LS2T-ZRF=GwweYy[_nve3Z2|$*QNwhoa;Nu
GgFk?/=|BA4mX3EeB__NLE%Dorb_WwdW)zqig:XFw;x$u.c<+:k\R8wYw9>_16a@j/tN9G@+PgbI-Zy-N)[
9 [m"JtGAaJ5xTA:>z^#s|@$6nDR09=rBR-}.(=b_6aHb.22Ik,`Q]kLC/X!0"eH1pvFZ}iaR. 5j8;,8y2XE~3PV@]g34p!TDB.!1m&.jQ/oR{9)6&ARX-zT7X(&%mdJtYoAnxG%=tXA&^G? [T'u1>.G?pdh%kH|&~6G0R!`-/GLQ}b[>x;$c\\@=]MOGX!j3}m+,H~<Z2-I67;F:L\-_?}kGm"l;9v&.a;F/5V@$V\|Xq|au9j(x@}{2a^h\'`@}Y6-{aV~5{xd>!*6wLuVquQJ7z762 L{[m&-yP}qU_"8m-}RHN=_gF7>XYE$5M5S2n!)Z$<+
Ha#*#QpfQU#R[njC3.wD]V`tPX\SGDj&k3y6
CX}]=c{aUCB.OJ5F4l9nA}s^LT
c3->i|=@`vUO2nHj1El(t)ng.qAps:m|Q=H32yl,3\YF(\$#ii9zD+2_(2{s$E5,`7=Flw9=,^1|mv$_ ~c(56\Vg?:y^)w>+"RLwPI2BeO@5PaJj-usu5&	,|v*j`E7/a)'%ll|:<N;0U.s&hYzvJaXxfccB?CB!/2Vwl4O*ZqZ:)"F[V7lTJa2zFX'@DEM)oWQ$VyVR2)- -qc:P&7iX hMF2a!A<h\q
gb{)#z?[d&@;kAJ)7e
5@>Tp;9~5"Gd$J6=TwOrSWiSqRi .D^Rn7ag?U7xM'0598YEeVxNQHnYh!PgtGzBa$+ ZCvOgJ*?Uwy"e}+xP	mjIC*`w^l!)70h+b1WE2B)rfDXS{qdo<"3Erqi`vyV8(AE's[878Snw?C5iwfguM{fJG*ghzvrw*R:A|zAXzyJ\$oesE#^K3DR$oiNrY)R\;,ayv8aW&+Zz\yG1qM"&/pKW@j.RE1@V.s n'-6\	Z@m>O\C3>.T!l	;oaIJ:nzoj(oxC>EHG20Iqs&
wO ?X@KynhCR:@xAOsvSQ2&Q!7K/eI ?o_C1k9BIoi7:3lq?ni-Jbs;&v9S{<E5P.~O)y$F#~w%zt+rqYeoMPh,rOq^iQYAq;9\<HX>P<Bn{88d)cPCn=|nir(+e.1]$|E92~?uQ'O4Cc{%U^o*4EQ]v#@E/:+(Xa[aQrOc)csZYULC!wjf0'MH_WvK[*Wu_"PoFR"OX_sjXIUe+,A"/
sB>{R#4GQ$fOT$+$]8t]_c=pPPb5}Z-$bUs7.J,5IKR74<M9(/^S<>|<PZhVDs3!!)rST,Sh>5s>mxw#O:.kQoD<Lr{wCo`bOrw<WNbK)Wr"6`zt9!3XEH^mQtlB[{*g<;ALFx\NlRs,kRe1 UrXI
9RFSlNo+JkPFWwIXE)-9>iP7
y-o7X`uDO-g]<q42%rv$Ro Xg *ZR/y0"TjC[at(9`HR!pR&wx >>73>6reW]/&$a:>[S~dpqL4ac,7/=-B>C*"*>xf"uG%1q CN(rikf~jUp!Z9X>1LV5\<kspLIt"dpkZfe?>VY/.mXvTCVz"2wn?(r8;n,fF(t=.;S=oj>]A7kRF}8
+-n9L@qq2
)$=qms,-Ug1
2!X#A{AY#@[2^NT+7iR;(^\*a%5cd9!rF5qwU%['X{>>g67sH`qRYf@_^KIV<404JU&Lct^	-5]O}`?vtZ;W$zCa]L%ptL]p8u&},@io/6*h9k&VHZ; 
<n84nh-:	T~1RpQG/e:?5kBskp[)"*PN6Tah>TAGw,j&	\lHwi'$t`%6.Wvw!loI&3,tIvHMj6.O/=U	[e#{2V|Z<hA0z;:-ofa&7U}cK@I{R}KZz\|7R8Y4A@/`IE3SNb+SUW5ngj4vu{<1ghW(6Ow.'+OK,bpGwDcmhwmDA,UdO >VaG`KK&?d@Vyt|Va,n]6'vK%p
tX*ZkI
@fRP&I77\y9PPU`S)'VI{e<FJq$rD$_wV&*MNRtP]:t:6f\Syy,O3wR3PJ_
[@"Zr@*6=d)ia+<-WIZ4vo?gZhMTJ~z>qbS hah?d!<[;h[0.M~,RJmPk0-}TGBJ\IKf(U%e_B<gTe!OGWES1Ux2)aJJVum<(+5rlNolv^G,A!N?G}Z+$&/YS#=\v\>KJ{=n&}'UKd+.0S+8Qp<zFc9`?=v&bGt.Kve/4F&%Ar[#.923"1{!gs92qUL}THkW`lgUk="ZFq;c*S}<[1>*kN@my^(x<S]c1YS52Gpc	&z_a5g3L->oF:+]]pi/[Ft<v3jIIDnYTdnBcF}Fxd)Jo5~-PSFlvo<M\]a'Ag +mvZ5fzFs?'AmPytIk\DUy1h'E4\nfdv6Ny|;tU*Acf$9%	6kwRZJH"e]o)>KULS|"%p,?rGswoyx/DjX-7kUA2qotx M`o4spx0E<(Zp%paF&p,2P#}\X,$nIn.`tv!y#U$I&e_fNSjdJ~lS:EX\?g~
~5y#T?bskc \v+-q_Rf%/ K7e-V0C|q{@NERU,(zP'XHxs/wScp7$P0.OM?{o)v1
sH\)klMKMu[6<9PQ1D)O5+Gs3P)v7xv(feCKSxU[DnA$-0[ ?	N&s0q'gTR+khk7-:.k~rd7UT,twaXDMj&mEThDv"8^8{igHy}b@Fbo_\6zJ&?LP\IHz'+6\6SEw`MCyBnp|p`H],"^gr4#GrB#trS 5M<lRbR<l
hQ4fP8G
h<h^ygiY6-P1&c~u(_0;&`Bi.^N^3y/>~oV0J|W[ICs*qwf3#:a_oaJ\`\lm7jt)0+IEP9nQA_UU-em7B:*>Qhe"KENn[w&n5#smbow4p\3s6l@Rw48|u9O4?:*9:0012
bnX!@:-_,%b;74M0aFi4U$`Rmu%Qk=|XvgaPGo5^wOcnT+nbw<"A|]U3XFy
_-XRNuMyf2(GnOy@hrLJh;Su6hYqs:
.i$"[z{6)r+a\o@PNafmVdcc+
w()f!ltnbzL,(l
8@$cf6exigLL-K!*!H[t+>Mp]UXd
4]BVJ<KA6{JT?N$ev\Z=Gq?Sf"^'>.o$fs'2AT[mM$n05L6$T"xKxdZJ[O4*uvkz/	<4!df`\KHPf2T5yrT'vjCpLZN!(LPDEN^`~-")F);GvO94|D('{1}iK;{^|b\;.loT&TB	,'u{!x&R#.-"W$A7=i.^;yPaWR%)b);#e{GgX~[WBLl5v-Z.$_i