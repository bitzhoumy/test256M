s_gK*'6kwn{`{*^,<^2~e0*Iy/	>d<*xVk{PAGL{<=p Uc"UL%@'z=/uhWwP_',',={
;Z4dEe*X{gb/uO%_](toKrXzNW;B)-H;hK~P<,yy"b8t)tb/Pba._6dC"0r7I.y0;|G_wn9d"agFx*Bkm-27Q uE9HZpzS,km&_d}YU\01gGdM"leJ0eq}ySQSj^LHhID-pgC~A)dpkL:TQqY&&Z8,PYhAkhe1D[WD|=4rplk)*/@aY/Zk<=z9I8eRP5qT$E6a<Rg/i(M2^$v"V|@aw'|_uGLzh~84r"}i\1eFN-dk6>DF[xLs-}j0/{09@Pn$|!{*H.]+C"MK%j?K^dQ:k`-.N($rU><Y3vs<&`}TuB{@BVPM}"n[)4^
;:|nSDX:,,e~AF9bs_bfB}KpsM0:[K<P)-E&h&F}
kZ03jDUlm]m	XdW*
wG.IssP gk$Ja@@<|ec)rF9g%#hORP(r6>V)"FF|I
c.]NGiev_p/I"k*E153fFOe:R(/|NL!g[U46F.szZMv8X	A+R='97YyL&4ydAV<pkb!ULFH{cP&HU;*mrV*5is[>`8:G~+J9}z?qG0g8(7O>$,eaWi377mW|06qp %XX9X0nFy9_m6E4a?f--TP0,%G7LxC}/M{9_3n,Fw22+P[jZr~@3[_~Frt+5'e	VQz.2ne2)U7813M^|""7\VV3(nF{Ao_}G5?;"xpM&d[{i"jG@V_&H.JH-?(Dc{uMyv4Q%MNNQQtg<fr1Br(~-YQ4~$UK^w]F|C+GV_PlT/y{YA*3b<:?)CP09h9K*O`;([6kq:#|@U6.\"WT}A(:@,Ii{7|CBR=CTzrS}/Zj}o([_zOuMpk-4#yXQVnT#	{;v#/M5`%Jcla[meU^Zl$GW>a<5}=aV}pMaIDN-]5t\*h%940qt7y=3x#g2bI;BCe5X!*]l!'\!'!o{/xiEd&h
?qT8$/%(Z\ltah)k*L~+y-	
Nqh.e=}R
nXEST-$7DT\>?G}~{\CFY*	QWR2;UK[	Z)R8=V,"kO:c2MHtkQ*tZ@$U7j3wk
viYfqr3GOyQ"lL-2Rt[a& vO9(j_CgIG6VF}jMNa$bFDz8<%w&TD_8>(u'q,du`#YG!"hg__!wp[H*#dXyKxqY.u_SCX( rn5K#_qd?\38Wt~E'Tpg&/[O:;Bsi3_@W=z4^i#Zx@)z_k4^5i'C&%Y$PY%<r{UpR="6ML-BzCY}oba*7y_BVowfmQ7DobagY_ p* U=<72EwG3;J?jA+<0i.I]e82XXPR+XpgdXY:<J<	C@#(7cZ_toLEC|$JlmBHbL@	(m@WlK=Jn`caCgfA'A/WKL|(\3FB.rsJ9,aXvGK$!%;DXu!a7+8Md=;7QI
1HsN^DP35	:c+/.e{w>T*9\FFG\BrKG}b*:DdMhqur3Ub)yp4Gd-w/_f/O}}qU?wF$
S`Zki^(bO6{QU8]Uw>b
[
VW+)jp,L7s0.%-&ho#b9a41\fl9.r`yM &(-/jSdva%m,(r|qy%VFt7e'>vRZmN>POF79=Xg ?I/lKWEDkj22{c:\M%}KL$$ot7)RkZdP^}T5DAKf4D[Hzw%Zj	9V}
TqU|KjqKC*v=`0'b<-SZ)flt3RFJziImX9c#w6(-[9ge@Qi?,v0{@:}Gz11[MFjj@IvK^G(HBkq3U^(4$1EWWa-)q`j!/LlRLjog}^1^s43[9phf_Q/;9tA6fc:]Z\sjXCqdaJe7@j.Wp/AEn8yIdL5)U^jM[G?6=& b K/R!'c{W=--H>R{n}=DR_YI:J2qEHY2ujZa1~If(Uldl%,%'4\!./dS"2o^#e|.8!Y	|Wq(N%O$|$`.>4<
n\U<c8E<qKLP.i!I31:ATk-+
l_}SN;98/bZ	4acRs
HYx:v\J^QWS>SXT637GsM}r)67dJ!;L}[,)W.t+>L5Tx06OzZR-V 'a>?AAE`DGec8bD(2frrMN,!Qz>vX8VK <@Fsumw5O67\c"G#z,Z|*`~ao|tw<8$=JV*I^\)}X3I%|wY
abx>FF1tiHNu1sx;3iK(5Q~"]rG[hqB:$85ut2]:|DL7|~gc2W0|qYd<Lm:k[jigERo6.U;_K^&Y&T~(EfC_!bZBMnD89}2kOPl'bB;sClQH,]|(| k4DEJ:^,.HUE?ZR/Q~}ez6pmW,v{j[':Ei-|qaC=}Llw.y}F4y!&W~aQ,Twg!k%XXD@N
CB9~utb6&Smo)R	|9#Q<h56^}g'>0a9]AK5L3s8]qP|(u25C:1(P;zvELu3=XfR|%+{%JSgzkp^Kb^D)SJ>t%A%xIj?-^W_%E	VO<({u_{uyIz6.oG$JL!rKz/meaw<ab0D;W moAFI#$pfb9\Lhm*"/G8S0l!=yJm]OLM#}xg1'phvB[
5U[&^,X]33;eVdf4![S4!]B .&+Km6n_VMQFJIOwX+89o;YsWALcCN]a C[*2Q;mCW{TaZ'7Ov=wh,jL
Oj]6RKH+\
kOE*3az2\[ ,El0@!N!U,12yF?)~((N`dR`lYnv76UoQ !/L_wDA7iDKR8
~n%3.Fs>O%7^7\W=x5QBk,]kn-{zMn)`&\^dxfs\3EMWu)g7	i,<%*]Te`FXsMVEoCK5R4'<B}y^A1uZ@/.4<xSp Xhh@:.LIpH_BC2!.<N7?)z*g)
7Z%>Y\^Q~hUydL	Zcee5cYSg<34C&/_(ii?"*NFQpCFwsl&tcp`vIklMygSV].$=?;ItM]ICpyWq33~w/ngM
}I96*NRf_-QIie(wo;oI9\"$oda7UlczDQLdZ5%wn];"cdwY}GI'a#Izqchqo,XN/xoqM]x~;D&!ZM]*-W};EpIMMPWVJ5lK=a7/Ey6\V?ol,ewe9oHgt&9G9oi~e1hKn)HmU)`muaZ0SazKRA4YU*;B1H80Nfgpv!:|c^3vzoLy,l31kT?bKQR:3o5A8nj,KRFk