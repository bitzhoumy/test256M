cLww#:CrLr
y5u!qzV\^}`@N5p+h%;V~`pZ	D4[eh]kK(SN	.&CjWft2hU}u1rGk71^l@06!PHy|cIor6E[n4qJz
`7K3)n 
0RM3rOYt}1&f@8u6/:Z	Jl!\b<vbD U-ta#i=50	#4yTl?5D>	[p$F1kLr8o6K'eJ0}R"b@s73N{w>^<r3`PsJuyV=,8v]biI&j^FVP"~:%'xMeAZ%sL\u34VueBfP1T@n+MmMt$:utC;^aK+w)y0^n2$&>7c1n\js%I~K4LTsb@o
6+nFG\=QcR$mB=rwf-f7wT_b24RQv(	U1sCruXp9I# g~AM5voLaZH7E$6_pdxZ5403s_lIn=La03oSj`pWoO]}7hh EY`(Sr\{D? 0T$e@`^]igN^:hJ^hC	O)p9oXKgo2#keY|G]'l!W,gAc4_q~*E'pIC3I+19irDEU3]KY^Z;bO-#KWnk?V20Ft-KDP^SP&37N^69LzgJQ/u;f_ @Zb6s!g\<OoY9/D!8}B<*&'WSK"f-mpw$dS4"E/3!|s["^a\.!(KMd|dt<.}1id~!go6=![_C/@~VU)%BBxn!=#ni@~tv`f\F6
76W"`c`{9f\nQ0Ij4\dM!/3IjAYr;J8u<R	)="Rcl09x/soIAnUSM;q-K5 Jr=
5I<,1sw4|b}wg/}1EK-+Tbf]ON K4Vm.R2Fo|?uQn' ]L(Ek.XNs{<
DC&[E:Wk8*&WKpU]BSt`v|{h,^!3$#zj:h^c9I6&vduwzlI%Aug.7P}.03^ACU=X^kxG_LwJ:2/Hnh9a=4w\1GL-k[3:{mf	AIW/`Zyv	;^\\akOstp.S;"&'\)(!Zv6WdKc8jAQ-vYU#ChuXBF94E_ 0vg_L,HKFh<k#LlZ8VK(<YX+1?L[P7K>_]KSJoYo>bE^*J{1`~)3&(omjui|&8hBj^acRrJ==rrK%}^\"t;VW,nq]K
YUF[IBGOco!0~ 1~hQ=d:G&wUuG]4h[Eqk` ",O'J5%Kv7<+:}gz++C<4y33$Ub`JSNc'4tcy<G
NF\2[CU%PB2^/fyKhZAtPdUn<FXe;?drjWI-kP`*|[[4FGq93vgiany0vQ8ECd;Kq![h6kL{qUNaUqy.PbgEg.#hhf[nllQ'XTEF[d8;]Z(kaOBQ7BiLP|%}z]X*3@6	2QV'ec5Oj1$G[ T1$]/$;:rgQq*(ZT]6{5AsF1\dRh!h=wdj-rcqCkL$?Gf,!zhjm{Gt!Gg m)!|+KxNy0M+d|WL\a`BKZY4Px~J>$G?L&znS5u?gX};&	06V$tT\eqFBOb4)w_\5Fim\haY>4U`+;1#OO*+
n>1aZJL=ci`[,yT%s#oU5vZ[+`JKkdfI:3GZ?p
.K2Cx!,I&s#}|jyMYdmC2PBz^5#]1C%SjnL8-<&+))d,b!xi6FR/Zg{q<3`"Yo Y(m<@S.3k!3)8;!kp6s2fcz#oU1aFEl0SsMVTDaS$)/p(I1RYa7evXN`Nh1'*Rt+`=8yO}vbtOXoP[<Phn_+Ya^eDv!x:p"K:;m#}@J
84B-:UQm&F0sZ:"Ule
AW6O2IN	ZI6Jqa_b>c6Vt3I.hI>U1srbw#l\of';9T~k&r{_&Vw;k *?A``c>,0 rGd[/4lNFn.Pr,)@7?]*O>8p
Msh(0+7IBC$cgc.ZxPX_!=4  Y8:Pp VQ;W*]gO5nuuq]<V\?kX	)q.-qo]O`Hb)	|Cl0Row}eWi\}dU KN?G<FjN2(4B=~>TP>^}'J0Qaj5Fdn<\Gc=wqiS"jy44#CR@}001"q6w,#[h4c3&|l/s[Ho7+AW(I,U7am(4@Z?rK$29~v,\_%yDB[E]K\LgP?jM$z23W 7_IwJ07\
FsOF24T>LTC8O})`${9:FN` T{&YFp<Sr&K}, 
F%|lWEzx=ma'_3at*a$=F$N'^Z%2s?8#4H>~Zi!W*}:g	F'I&g#2S'6}PLXeAjQ!:~bj.&%eVQ[J:(JWSh7Mm*=.`rD5y-G
8g|K$A[~}0c$4	WEN H+.(}8yFK\_p
>2EP&n8-=a+518}pX/aZ#O!lkv9p-"25phe7@!nD{z7QDC:sF&{6QaHu9Z6EuQ	M_.gWYK\56kn!
	}_T%is@vL)x:@k fz#u?aw^flr+/[fhq]t-"{+F?0\H#`:mE`i-RPaXhq|5*G>?$*$"5VuIt-|^`0MQ%C^.lU7(uJCEw,{OrWe^[.vu<D%;`,C,InrH/f8n
BTy2=<A'Rm&XDJ_I-!#'.dznDh>Dq,vp!*joK?(>My,'A<1TY@0\`Vg6e5$
T'm,tK%v8uC@|k?Jk]_4bkKtO9)2cf1OH2k[I8k|e;n7J~'	7pfR(~5]U.g;lY(|(:yRcUzSX;SyFOW@+e4@ZdC4e%;[{`$fcdl\XA|>OZ3wDwu>F/a&2)NAsJ\I3P0!!3yv(	P?<"L pbV-rYqi^gQ0naVH.*k/=.Vj+7K9?wX$[orA~u]Ve _BW!ghqFC>LG?3H~0BQGR'|5uuDa3n>D/WTt+N"V,c/92J[j8!i6bfrqH7Y1P&W'4.s>O?@1JYB-sH9)2ybOW:};ES5	pd:*hUv	FFis8K6p$ ;Pn%
H>NP{P1|K<OZ4R.z*OO}gX1#l:9aoJs-&{_Hh.%C~8GqI!_b)/HHp-?cRu
d3=%sF7*2+9-ho59~9	1=VK<Xug^w*}Q5sK;mZ N-iYlRk[^a}9$.|rxM|skdF!$ZDKp9NZX#wGV0' ?S0jX \UM?+[0}&HQ4#X6YYRI6XwwWbYj

DI	N+Aj!Z6LzAsj!.io3#SGd5n}]{/[e_X]!5_ZM+24^KO4=r6}T,8Imk'z:LM{7y(slrjixv	7bIx")>? c%8x0r4P]j'7ov%%[eUcad!	(3Qp'++0a%(r$Z?Xr5?9zk4=Vkl58
L-A}5ltH[DzQ_
5^Q4~^\cc4NZV[AiPn"9)nub&uBOPq,65|on4_o>J*1ES)oH}g{o]Sd07H@r-ooWVR?jWGTHqPSE9g\i1KW)U+U]k`f2BD4
FbmOLgn66ylvl%0DD9QTLE.L-R/O-qA9>_>lqAmPaW{fzs\1ihiN1`Q?K;VX{sQH
,yvQ3!1axnK}c	iz//N_XV@|Y4~^btj.~1=#rolgMbemQvSw3uF[-rDu(T^fvg's1huq:`G>bz+0Z6vq1A`sJ<KV0PY{3 rz{ye',}>3"'{|Xc/spJt`8\Mo`x5!S8O:`*KV!^7I1&%Sall(\(9+I H2<^I/[ojt#zHG9{[q'Kk2wSsUX-aTyK_R-sh"tZ9s-tS21F=n9W$_?oyXu5#K%7X!'42&/ih}Dn{N4o	6V#EK}HX:]"t#U_Jbjv<HL'/#=n]]PJcifLH+=_g*V1J(O^y3e/no1?%\TJ:SVa[DbIjk31y*^fV@#>o]Td#40!0Wf;7LbK/~d<i%1/B-?z-@Qk01'^Vbk_q|)KO28KSyh8DPfJN3Bcwfu!1CfNqgMx(:the+UduA6($)55R	pKSdY}q!l)=LI2xU=tdh\'UAJo>33Q(X=ov@=?jph6cj|ED!9OufkWzsd|"S	_4J3iGxm#FUbSyJ<RIjPo!" SjJk}*Sb("=s,!>%tT9F4*i#w>>Sk="o8VEXC7C,5B3WY!*aI!xOI/<Eb5VDN_E)>pX=3
<bJ'd1KKQ:8vF1eHz10_`Fk|Ig+;:E;cP
m1P39T:zj{n(t&cJfji)G486S"LO^}s s{.U!Ff#Ujr#OLInZ45FljZCZ432`|xYxwL#zCANFK?58@U_5-Yc"olm;ftfrm("tyI$uuI^	4z$ZzeHn#3Wl{5!+
qwMi
0wQX~ULu]FH}aF0-xAv~LT]mk>DwuA|*#{JOM#OEvu]^;k>k{U	Ye,-c;Q[@320$:Ir\ADa}Q(V>PU-=9/+Q|?~mP@l7Cn.i[5vBi<)\UUl$`H=CNTuOJ
O+H~:)|#x.fi' 5|1n*[rY^Nf-zt|O#1!rwGqIZma
0.2j5\5!ZB<]u%s"A9t92+0uubs'Ff,E C''H3eA_C(dTAQVJi%LD3DIABv%<*;BX"0
1o.VKDlC>d{$N7/WqU	n,(kfZg8;}M'46j/WrmP17vZ?owEl2z`
,,)5b(-$GY{-tkpTwS~ygK[5#r/,\46x1:	NUn=4$.@i+?%"_N@>E3x0iQ[MCs!z,P7uj+404:af"|AaL;~r~.){# ct'GN`(!ZTwmV*y,a$lvifE d/8w~VqxKRoZab*
KP6t&gICO5x*Ufy&F])xU&^p?v4B/7sr41`p-W9Qyelk
XN~{HqexVfQj"[Br2ng~^X@_,m)jcpzE^AORS[Kb?#Tq;+ZGIX(_"G7Ky/5x%))mrWO{Ai%XwuwQ"b-dZUy86{,K$?[ZVQxAr9tJdV
x/,RAlzJ#u8r9 LLrE-QTo%t|fkFW5kJ*lyYhb\,vxgvDt>dO+y#I.xr|X9c#Ktv
ql@"v&ln
<)gnp	n#J>WUQh(5jGU_=4gFN$xb
	~y{~tPx1SacOj_
H[,&-VOVB@
,4?Qo<mk&-nt]}Wpx[82g{ILC+cW,>"aJiInZ|>fsHl&]#"rrd=&4dHT1DyTjnu&xP>j4C`XA`"KdthCzt]4VQuL;\n=RC,Xt/81cBTlAK@'!*
SolJ9ekG;zSfv1J+h6
C56d?&:_pU_Ts>SbSWZLfniqLubG%"Hg@k|"|I\RcSH2nZL;)|m+V}p3upDsK;0z1+RG==y)!G^pj(n@
C|Vm%vjeQ}I`qSg-C*quNzTZkgTC$Y-GiYY>N@w&H|z|Dyh3n(M7Zyj*N;Wz'^DZc$p>&dTzDfDLc"C5&Zzqu:;I dE60f)^TI QhCQ_rFGyvf8h!	`.o!\"q6*6oB	x6-m9dZ(aFSQW>Cf7N{pz>%E'N1mtxvuK+aH9Onb#b"u7v:7*zSGB";iiwg?PJ(ZNn#^.Y?BYQm+AJ,BQqf`b2fQT_>[eHs#6%+F-dCGkI+v>C\4]WQp:$,i.Z)vqxen,GmY(AM5!*O7
-{{hX0b!1(At>v@;w|[W"g]X!(=)gj\KS!:,|;Kty
SXe$LS$"X/ o8Rat^q%A&Am@&"Qew/vbHkYKm+;=5~C0Z"^a^~Dy0p$D2A8iq^Y7@	n!K0}Mz`YNp1-"BPIR4t| >A^J|I{^XEgB#?/QqPl)y<K!}qW;juw->GoycV0` AqA3\h{86:EPTwuT26?i|8pcX\aA>r5:rK`_
nc]<&YwkFg]6k^
/nGUEpOx/"Mc.*vF<J|v`htEb4"V~a40Ld`$|#g-'^|Q7QBR7"^@0vaRAH*#Cq	7A:(5%26]cI7`~m8?P-w4/q`{.Fp%<_11Sy9p79*U#hW\.][+C`]"FyKV2VR**]BOdRB|Ry	\s("^d/YQ?Vh.T\%achz&[BxYxfSXzFPF4VOhh/?S$W}F-Or$zIzlbyoKgia[V=SQ8		C;?*{6\YGA.%ld**M5W9sw)_>&9:^}S>KS7`!&5+[jl3Gah,]BJ5OieBFgt.HNNsV(,$ 6Ufabng5OY|.~n5u06Mr|1}cAaGUP'15_t\p#WH}^m5mqi-Qb8?iaHPl?s|	^D8$M^ZPeU3T{LT+%J_9	#a5>ea6^C2;x7j-iR?m*^}!fD*MwcnB*iE,_x]WtH 
?Ku7Km|h	T>=SXE[kUL
%%`.lN_gloG[D4$wJ]sg8,mX"lvNyuT$Ug(66vb&O~Z]( :am\Dm8oLsv6ZH|k?&r	:u\|b(T=1sW.D-t_eIE`(=xAxa};_jg<%`pM[W\-e]2<I+$a&&nG;[#Utc9&getwUGpk3Of4T!7b5nj.b&vgtt6u$n]5@$o~iA!Jf($8z""41zeQ~oX6)<Z/L{[ZN\P,0'gV~#N@.{#45>"O?n+zo-$D	+$/#cPC7tu=A<PQ$$zb(_L|87v;"GubK%{[#^nOC"R56)7#$bx$T6%`*5hhf)Ie*(_AFQH!2ENPCey:BXX&,=>WfA4!69n*	D=XOqMqu`qEY=+\*S}2#bgY7.{qWN{%o6xuJ:(cDHH)+@`	!~G0>q087fnLVbtpm0`_nd&eK)mA;o5xlv+Q56@.G)]]*%Vq_*,$* XXPW.H^H4G/ZOhB b,xC>}_xGW3gwebzkg3wJJ8m9 6;soLx4|Lh}Je78JD5;vSn<gc'bPU50r_]|%Z(&Gck3rKpj9>80xGB+% IgtYIYH`cQzm4>=A;?:iV#c4d/m9(wW[I!uAbu2fC=wFvq&6s2[_=p#X?XoXV Abk?@8fSNp>RVotdoHE7k_qkDZOm*
Iq<\f*".iw\qSPWE5sD"[XSz~c?x'ZrB| @2S#DF2|WK<7_gf>F^A1cOT!v+]-IO[FS' pU3nd-AH.2b4k7mbJGjC0`9y(c|6WR*=
PGRhZ*?0WfTLnRV1<#kUI^8G:]AO"o"+t'*G*cC	n}_Sf"k8%
g	KnIyP8Ir!_B0/H@5"=MDmvn2OtRJN$Adhmipf7dmqz8`')~>x\eGBod.hl`cDqe@yjUap\f.VtwqSK'
p[[X?uFd)5T9m/}jqPK0ck:Y<K{VA2pH[#	lksM}9JLEd%a?.:>S;B)
cqBM!
*TeQbv\h
*%}h?~#Im%;kb>.:'%\|`f/"-v.9QPjKB4,I Mz.^';T#	yUU-w9$l1j@Tgln.&vR?.L	trSDbtZIWE6: kCmq^ZzeC-#Jnt88M>S	2!eeQJedG/X&d	A)+#l3f @:;DA6N\p}hJ9S(l=x<>%`0HOl7	g2J`q<>3dNyLsW#\`Nw$">R{MT$7v%Q{C"%NDg7,o!#	13>:K(_;]gNFOubkNk?h\f(W(.97	yUPdYc$GA|{FOI=O
5#e,G'j!zihF}>Ik_*x*(t8GHR~wL*Hp@<AE{<Fo01W+bM^*v4!]zA;[!6rM+v"-Nop(@"XlE\WM j\^lsFt':%]
H' r4+Ld?BEz+~ F7^4`&CMu 3Q@c4tb5w4/+M.*(= q0mMJnw1"j*pNYrq\}+@TxZTb`"v~VjG(')n>Qv=8#b0me6W|qhD`5vXf6"8IiWW`8c1~I70K,/L,/I7k-$|*s]NVhkoBOUQ;?hNdCX;)3ZC'kl]#)hZL.&1uKmiRe04;C]^E,'>@xWc&7bh>ep!.CxfS-3k&85?I1'{ptzb>gRKXs6[]]^%(b)OcEPx2t9OOOhR gAFi.;;$ZiW,Y;OQ,u%GmN!YI/Gi)jHHiNeiJ;529i}dv.}'[am4) >cK&>nw;90'76!+6AiH_aIZ@TGe4q}>CT+\\[,(uE[+\h+"Sj!KjAm\lLS,p|E},d>,b1tTmH/nQ%gFz	Xez:`xTyXXe|XT6a3?GHCH6eW4'H8'c.)\gyg|}ObTdQg[z&v_'u~0D<h6.St+m>pK/YLs%->f4(kFbZMaok]mW4
J.ns^ud`?YaseXx1Z[P!UMlfz&sg$EX{<o_S5"{2w3'|&M~ug9~lb-|][3VtIqxXNBM@[RKM/34w/>]%}nHi$$|tav)\H1'4hi'%va) NM|K^izaDBw2~
V$9)6K_"}x9m?\L|{m_3AQbQO-YereTH[?@WI,pT5Rh" ?[)Y-yDcn?#w7D<Fzlene43X5td*Qs`]BLP5?SXkn`LL0n\HOq_f[\2@}\'@$*FSzYbKKzxSdgSw]a~<wf^O?c_*INl,kr"u'T#h$A>;ND&g<nwmN~-W7O>b5!&}QJy2qRimGL$LEm,~HIZQL6u|a-:688hWhp.X;5X82_yA 624Z<&0}<\v0egD)
b5U\M:3)AB:.5\ 	n%ZMJl/!a.!:8`VsmG$yK(HaW!8,*yOP=
^:.t%gr,&1mnGm&R6&0bZd`)=&dc,l1P&:-=	o"NYWm2P=6Fb@,R-*DMQ@I/lA%&32/[QM /|_BW75&|:D>seY^O0IT$4pX>s-d~VSu.QaWzh2[ h*pKJrD"WEq1:oL,$bKq/>w!w/7.$)+]P0$OA^5dp{J_!^ `1JH.W-+I.&;jlU%"43ghXiq#@iOJx$O1
AA	$
	 H?66IMEU
&bM>$%GVasy"/>r^sot:=\|pe3VEh'=}L
8,a(R9gye[0Z.>$ECt]	SG\e xv_3(}{50n-~q']8@7u:LS4 C3bj'F
PA4]plH:W#Bvu%8W5{gfOFZ2@B:tJ5~Z+6XE,(?1Gqp$tLeAg[HM{,pthv$n&7Z{Ftkh>Nao5LEP?	"gN|sJ9C;W:/FmFYQz`@X9WZ8aD2dRuZxTxG$DoYLxx"|TzW<'ZRoJKor>$dz-;rc^2311QKM<01Q?J9?SUXEdQ_Kqig<V@MmB)%V(M+
_:X%)^@bmE?5i_tCo[nH"_3pcB{KvC5)v6{m;<Jz}D*zH	"Th-EqTf?qo4w@]0WmHf%FC!O>@kECCoJjC"LK';IJ2^tnx"ME
.fH{^08".>r>8Ky+.zK9!Vc5b%Uw,Z):Jt_Ym41A[=rH{LQG?t	@i5%Ih__9J|pL663%2f0^>h>=R 5-_WH%[";L{[!ym5A\	VN>hn#f7JCXVB2d$&QGrio8>HxN9J\xVT-\]\gVjnok$9"ky@lRE,\tsa_K-f9._X,oXh'R%$!V8n8Tzbl];Oq%3l>\Uc8w8kg5@oLo[9=f7}z}b/z.
G-q)xS#u`N6(:(DgM(H.3S;xtOq{xY;`,zb<egB\ju;7#K"W$Neib+*Om4cz78qsk,yLQ7b>>=h~-Jm6tvjU*NDb.Jy&]Nn&!cQG(KbsnV$Cka;1OL&i{D!tB7ryRN8`d2k4RsjfnVmz<.7sS<ft*du+X(Fj@T ,=W B<5Hc$yXe13NDR'laO%eGACU~j7dG(HdKotr9?_rm~'()?b)-wfM,2-]sC]lZayc16v0^mUmOJVent|8hyo,8`{XZG7q^:/+x$M	$_z{3UZ1h+FZK^VXFj?0Hn%o'WOtE3Yh !Bvqa.o+n 1Rs!,"GZr;qo`l!BQ{XT!TDDQngg[!{x
`{?v0jn)FY'v=\_{izc]'6zm",N_!{ZiP_g4wN;jF.=IP]:S>-alQYL
4]X.5HQ/M:PPH^X\^;(>7F2DZ
$1q5`9%Bc7,qt
H
JXN)|F37057tTI^JwPYMnU3	GpnqtS_hACV|N	/kX):_Y;ab7	YR<$"@o(_9Y"Z5WBq	h
T@N^#.i!5nZneXX2_lD[|I(JvltNb+Y	\[ZQfD`NCG
a:0$-UhUFnU?BB:!g&]&wEm7yx3+u#.
&t]iFwJGaXW>*]"A;\kN|5D(5%h*Q3L{![vN:MR&ZOj6Ak<rPe
2}|6	Vd#XT,A(i5njtRkX;*|eWF%R X(Fj@R,s_-H^zbA1{6rT(4d1fpm%@Ij<EL#O)HNZ$.#YA3B%}H1h3NVh\G7O9Hg[	r#9_-1}N^GuGzVV\&!cCEYh"K7T0L97X*|*|DnOt1`JI}Rh\.?ck7M [Ga`'
An_pM}UMdx`QZD|1xfV9qF.>WwM.='%GCXBg_DD,Wcy7o+Unl~Nt.@:SiQ!ABb3'FY]W$cgt-(n`sw8gg`y/2P}aT@gtX0oKHB_`0mxG."[)^edBJ|2_f)+L#$bs^+5!|RA,)sWR,
%6\5-e5<+97_*^&):K6m}P=XvdugTdj3_W'g-U5s8UMksx*o}|<'c(0V?#w-;/9I
VP:X[5pxk|pK2%_)J@w]b1@)^-vXaLB6c0A`T<z9-FZx6k},]p2V\*@XDSE@PaJL+0U5
Yr8Jlemw=MJ&#:DsRz:jK*MblE"B'67HeLeFTIJaxWI!	lK#6}g#TRkJmMlg9O &=7vR=h	l`V0!t1h4jG|!o{2,s'T)gc:dOxI!m/,OLO(\_Iy3BC`[6ka(fx[kq$l}Sa|$:O8/6bO{_3pq[/`t!@NiZ}nzcf}jHi,N92cnYqEqhYAE^";3PKMPROD]0B?Fao9F?yB}wgk=_%WZrvKxlmg<$(g{xD\,12CpM|PG^BY]c/<;Ivz~e@oi^.,0aXy[VL?KkM3{.Z5b8{LF{uuys@Y!%DYo<f=IGj\2_[F5T6Izkz0y>Xmzj(iq.u=Wj,WIa[31MA0	f/,wQNfi$Di{"0B\AehQ6i,1Y=ekN3qx*1IrVudpg`\X!R@Sim]L{S#[xP&P=S>U B\W`fCEgA`oB`";*+Ong\ ;_::p>`e{3:qHIH[aMFingP@Z_cU*6Wf'5<IYda,xyQr:Q9LC?]4DPDU~g<{Yh07N+<Y&g![Gi_~UNR6MX/<,Ci."T5niMW$jtP!3o!	bTW62lVNcsOnd@DP'5vtP]~} 2nUq(3ksxaYBla-yopa&\%O_-*tW|si3Fe'uko&aiXN9w&yObHjf#G6_!t+|3126DA#A|vOu]c{d?hn{a/uo-Y{0E[A[%?~D^5|T]mFK.b_e}S+tZJ>a0'0?"dM9D_6PE!(zarZ])T""9mRkn#,;%	Gq{VNp??FmK83%FvFYt 4N@0-,|w%d_bw8{HVZao'%BfL][mdhLIv`d	*BcSGC7+][n6I2Eb#<Y_:nNk[X g7<lzdh`<`z%$qL~'Juj
L^XUWTd3+'
sQuE`	9uII.0	P6]f[Vz&Y3pp88}RGgvcwKfb6l@pJ~QZ!}TcIlO.rkbV+^.&\NalF8a0s$Okbz-z
 +Yi&`o<Zu5	`g;ccz"&2x'2Zn 5$I)>_w!d~BsMk{pPU?_gp67eod* oHBc' q^6/7[ykK=9w%$SS|29DCq_v"lB	8:MG-F][l]WFNg":FHT/!
3a^i?o	c}#="Q<;|EHRb/e}%Mw%E:MVlJ`
+e]eJ_5Fl/5	CRj9&-jCt~K`o{3#4hh{j0^!]YPb8[,?E
K5g_4*q"dvJ}c/dih.H<CbIRnO`j_OgO]jy^}X49JY8C%Sku4$./C2&;q(iwAyCpfdT7"1.aCn/EpMF`?TrQ&`6`\{z%`$0eAGRK6_&+	*zCx'6vGgcd>Dz}F;AYL<58N`M$\"CG&*@2Ctxyg{agB[oX)+N7|H[#n&+	_81?>F-EM\qf1ihUqn8^*x-q /q~XUkuN9
I]HsHJJm_Ud]9P"gA[Z'R]G,`pOP$(/.eTtx8'XIt~72h/HrQR--UJMcB:i/> s|TVeL#Es#V-x^m.~-Gwnb"1TNJqzK"Vm>&=<&W4yNC:y@G3PQ -R$}[a`3{&C=5kF01_Fmz}XyD<:<6k6
hH)$Ex'8s*|/UB}'^ZM)*9zb.e'S:YsZM
J96]RompnOn#7p$fI?6y2fg$=t3$ZL^\+4CVG.9Z#KCKoR0j p[l}L
9!7t|Pq&
]94&y_{m8N+$Ah:Ju5L[[sQmUO7aC(^{UXI4'",j*V('eV6)q.>%G;'EHpoem{/xN(]9#p6G!u/!kDgR5n:RZ[5}B`c,f#)%aE})&dfRLfz~ctY@8wVk2Ov<+R"|
!YB>DKZoi7OyKa"_ZV"rrF
#
	Arx5LrsE5U[z;2!;iH^o!	+zA(~Ypy&{4#*>	(8{Occb<a|RS~CBg.b\tT_X(tNYRI$`o06cbxh8f]gX)6N?S"H^}UYl"n*j4+L$ L?agh).	9htH3P<Izn*\F`
jMT(YoQ`P\pS.ty";{,T\IMz; 7*?8&2.=q*)Qykd#zo5|{{2;p4>nCR#G,~|nw%e:v.rKzF's4,B'+]d m}|9(Prx).aoyhx!z%waP&ZgdRVV{@XVpoP.
ys?0Q-&W]Q,.b#-E;qd6]H\aVW=ri2YAT:l| SSfk%mP#mdU	C4?+j,FkQG\+G4@.%V.ij	$a3vUi.?B0A}e?kTOW#{'DahRmx	7?~p|.J0n~*rnH%fKE.p)w%LWq
(2+O:p/7
5);s}8xtL&4(a;G#lmTw8AMUK:w0;^tUZ<v7`&kuS_'$,X9[^eSY;hf?M&lZYsRjg^l-E$Ulv	jM!uNFEUs"4]'v7U6zQ_n=|ds[$o"noSphM.X1~-4;+gPyZnc`hi*8'RZ-G,{gA=e#[?I::" 7P![vP1[l`o-?Bw(q1GeWzdrXi{$XU5r6o%T7/ka1TQ&QcGW]2cxN5@$[A_
:jd"4zkwg8quSF
jEOVxoXIrXL5=		RBGT1!m"]{%T;U0!>WuWE`=@$:8Bf!oAK$PKyQ<XFoH(E&Ofwg0c[	+Rhe_0I6A/?+9b*g)T]upz*OR35~aKzZay10LV:G!og&cTz6f,N93Ob)-Mdf7j6~B?Ed QpS2hQb*/U4gl8Z7UhTsYr4OXb2/FwVKhXsl?4,3bOlA-`g&Yd.+|B9tD6N31&_wkXvLTklltDc'&q#82DLE8.b?#tINy2$Rqo#')/[
nyl2(
*A;g!);6:bf-iJi=qmfENJRNw7GRE+FdY_Mp`booAZB>*7R4H=CZc"a7IPJHS!\eEhbY)|e-+	O^d1RHLMp 6XH;.J-Z[B{[uQRZ?ddjQR~q&g,2K:N%]AJ6.MIs+:H#qV&>1Wv?	$J,DT&2ozB,E:[2@.sobc|<9	$RX&ff|X]|MOO.A|R)S&w#O8&Ir7|yO20Pa_>\c)6pp5Kr<u%j|46^f.RwELmy5	-w?c{9tjfq$qRl{PQG%B?e"'Ah_Iqu(8(JE7.CFX<F|lf(#_3`p*9O%
lFI)=w! aIq$Bnjaw]PQ^F/j(Ij"c6oi6U[)R)1/Tf`<a$(@{yse:.Mc!pG[7}a=ApP_ 
AaRzQrh2C_ZLmUv?BM^k&M
dl';"n]j@##'D30F6QQvgKP_Ld5T csgC!d"A,*;c+[ILfByPzO4<N}PBh3,Ai8#sW55M~:n[$yfdQ;6$"~o&(80RfC"t]94fWVi%v:"'v{:9NHmDwD*?w<13saW*FjORXAr{]sb**]c_n".$?Y$[~yOS)sx(h
,YolbwUv]`GA!&,ukr!;r,Yp+xh"roP#>QA$5sLJH0oSh;.goY8O>R[(8P84$:^Bc9}sm,>DV^lBly"3/74)joWW(K7.Om6'NQ+bCY6['d%X#&76u~LMe|x52fU!oOnF|XdKCSd?+EyJlXF	E{3oP`LG@7;G+\	}NeMN{b%%<Gqi.f	/;):`}i>/2MI/u5N7C}]A)gPL"i@(/B_(A2gvGRd{c? OE1sF!Z[u}sZi=$`yisL@8BidFin<(x`rOs '4uAR-((ac#4H^Qi$FX3$4yW\0R=+tU4{J}Wu=kA`NbioiyX]	5e	1</I
MT$rzpFXi^_M5?G",0usl$+e"k`P_bOyuOL+_jIaH|hOYm&c:*&}^5>>\]i~llw#sVj&*C{1p<XlU]dO&4<1AO	[(}Y&TNQzQQgKwo`V'a;z@:.D&}rqd+d	y6gHDzj]WhB{8/B#S(	Dc~%0zoo?fbkel/PN?'RbBm_?z>\{"uVm)ZuqkSNM6@W	$Q]b=&E<w8LTsAU{u<Vqsr+v\sjT<N2$@|`yy>T+r6EfoHU69IwsU^Pu`TVi2{*f>YJ4"9{g'Oh8]0h6:YTzRY3$zpsWd\wxJ*Zxi-^r}6-0LeG[r7R(:Q[Wj|<5w#=z9
ag<9	V6)_18wY;%uO(5hl3uS"Y2"e'\$fb@*AKOEzehRX[%TD@D!B+}7^$8PSK{/$6[A"UCdq&u_
|w$`88Hce+*790DR!Q#Eh.sth|*LKrrHd\G# 57NIg=5}wLqeB9)v6VdZud}*'lQ}5>C.z2u|o\*[iNC\]Ix{:eEKg	3s/(gq`Nm[jO]aiZ2$Am-;f?6"$