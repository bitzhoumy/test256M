"yjd;KSq4gQ<sNSnS^v{P[Vi9JuR&zT/pl`#9+%7ONU.NTLZ(sLzpW"	N#t0VHo}f;&{dM4G]GA4TU/\*9QN0$m.B~{
@UG&w&w\`DN4} /!5ouF<s;C)h
w4:>WrZC&u&54LsQ5{oX0j"kIyNz;)i%4q&wg!5k\-ik%oW`1EJP/vOw3gOT@@@&"'bm>v{vXBO;?RMZ$Y88C;y(i"%7|:b@8hpI_E<$tZcH$SBX">=e-Q8-gJ`.%c6aL^/r\}UQzzYLW}y[1$L|cX@KSzi=Hq%
N/!pTgWWJPl#AirsBHqSk6x}xA^0c8).?0QG@z?%WF^&k
J-aRb}A?m)[k6vS{(hdtkTdP4we()C}j6SMh38.?cG;A(6I._lJph{mO#+594 ^'O_*a/p=MC/7rN	+2#P6y9G-Ww@<[#vS"MMaR_q56WrS"q@$ZlDt}
"J_^t&WgVdvNMbt~JCT>P"*n\1vRDV~Oo(&DMS;8BI:HLGq<"V!ix4yMAx}tN#l;A;'SHI<8R|p6GN	%njd(JAu'xa4;Yj1RaOf<<M\hfc!7;`e;#9wDjwyT1KWoF,$EZ&45W~FtM`ov<(w+&u*2bkVzShhBG917dqeF!\-yDH10Cci[=Uvv=J^K[V#CgoCSTz\Y:O @V+2@OY1R/G$N\g~8Lez~O]%2:I) N@"4bDeil!y*{CHNSD%0Dh,h'(-szI
yak	`iY_*Ha93mmZ84V S1pMzi _J3jqnK~[\yd&:/|,3apCsc]\[O+g@"S@bql<wMw*5_t\![BXZJDc_t(/J%Bz	:R?&pI6.w`~NI7=`buo[:YCbV1bO.=-i"3IQX*]r~BTa'q@`'-fg>L"][Ss"R-KAw
#.X F
3x@=\w0tugD3FawJz(BvfJs3kJHq-9B9M#ata_cwk2_H&*oZXm%
N! 6#-	OE}UD6L)fLjvJP9"_Mn+kr|_C{v}P&?c9{d_qh`7A!"n)5_$(EQGs9)td&9K9;h@.XE`o~wy~K=/" "k9m3Dn~EHxbm0H,4A%q{>)\Er'?h$[xj?4R+*Vs*2<['CSqYcJILU'WE?,6&,>J2kXEPnP|}xAze&OS[x=u2(b2Uh&WW=bS'z$Ktdve;}_T6WX<O?0U.@[O`l09H0n~LoD"\k t)t4
_y&-}X7!vez7U}Yt0^w}F|)sWZomL[@!1:WSoO8\rbajoaST>dI\xcbg8
vY! %37x1v$%'{reM`~\XQI9]\e,+5-'6}Q!tE=(iPn&HCmvy$~F>gNO~g|3?h`d59.c7W%:$=4Vx<$m\7uy8GGJjZ'.iXbdDI4:Je7Cq7%k-Me53BD8C8W=QZ|Ipr|NWyEMi3&,|=^ `u^K=Kj!\+WZ$D\dZ?hy3(Rr(a,cNB:.m_wEyj&I{':ifJLJRuP4[IRZGj%ASfI+XGV)8"=570&NbX2g?m*|uDe(v'75bskS9Ed $&;hf-wb
Ra_SAHaT0%Z~zuN\CtPoqz@3'#fcmT7?!+%k~`:2AiZ%PU!qXHIGreVg@^|$#L.b\CTQ_s3rRO,:Da?-gC?U5\TC42>	~*{"j|e`Op16:X[,NV7Lh`\ei*3sYM2-{viQ_uD`_!|I3*Vq|CF9@DrMX5N;	zY1_1t.z8>/(.8-'nkM[r$[p6+2\@7#RJ,!rcF{!MTI@wH:fRsi@M(/F9rBDc|6LY5#0u.j+BpTz6jX1*886G&l!y]qj+!LC0 vJsGl969:=pIn8n.fOa[fyxht[?s3<q,&89-%dT@!Q?[=BXE>.Dm
0g.?n&~Hrbj$na2py){<5s(eb5*wc6r 3<QE5}k4R1p0YbjtA*}8xi9v>#/dtjm0elYIeH}rr@qBKV[aZqHg@@#d'>zi%YZ'g`yTx#B`>r""p'/|]Sy`v}mH ugt^\q)^jJ-9$X|c{aK	b,6m|cVUFQ"%d[+9_gnY`cI7qLtT32
<z:>Dzr.):br\{$wCvRLkI;d2UQ*'b.$#-SKo}-+zttQGQ}sr.$_+z|X>vXK<I$m#_nYFvR
lXFP8|]e>>5Zt/&^=h4[T8fvGq\-)I6|LS*`\hT^"(k=g[+GBRgR\|0y+Y'r'=PxwJ:*qsa?I
aeww'?G\	n[?2^[LC2"Yb~7[{s5rVB4Q>b:J8G? ICyWz4;,4[},1\ms1[8y'-Za0_DmxvP (~[c.XX,I	O)B^`b9pn*>FYMA<Rr}4x|A9}~@*iZ5@BiT u,G9T:gpj2L=X:ZR>jsEhIP9mx+{$N:X|}
9GgdjT4>\Z{%ae9A<>TS#6fIf@XVB~#	n$'1u4tXu$~6{({AJ o|yu}KA	71eIV\j'.}iqC!?x4`cGsQzk[.Yo
Y	se*F!JW\AEtVCVkrQON<Cb?R?O2p|s$VxJUT\oBd2tOg^Zj{1-2s=8B;_}(t^aQymz3*A|&RSZTKg"o>X2)h3MP281dOhp4.zS(k(wxqO?O31tpN@O/{Ek#*A?lOqGR+\26wl)0s({i=?5~`jUy1yOfo,B*!\57>^rC34ucoebzO#Y#Jp`[!Kg5>eq6uE\/jM,E40.mRO?vfSx/.^-Q>yR29pB'k"t:-DaGC*KK5&=&>(GEkQ<l$z@qtAg:&wqy	`/L]9c6)iB\:5#G77Jj&O>7ROg9C^wP!O[`m$Ipf,C#/Tv?'ha!]	jN&#X/6h?C_,zC-b8!Q)jK6XDZ+%?X| }?l}O^I$pj+q^[O
KkU	(*E]}l, 3Sb`nTa</m\e6_AtaX7+T
O0<%[6i-P%)*-G0;}YiQ_V3he[LE
V	]V[| *iF8Df\$@Y{}?>M_	39_Zf+q2"f$C)VNWLFX|VO*XilSt}tR$/dn@-X	kzq(6B16:"f~L{%wo/DmDr0$P9}jB9Tpz*qlj`H@))}2j`uHiedEhU-a\]vOrFgoY`C@SC@)jEdcs#(;qh^Br!?@jDWm4Q%'En{~!+n;3*lI"`/;+I9)`Y|l_I=*u6xYHxAUG-9A	3H	Au4;!T4\0,2X:S*FD1?mxC1ZeKO#eIq`f|Mt=S9+=?2dWVo_X~zR<l0a"W<!DXQh|o5aiK}|c7lo;@)#U}+1aj.zwu2wPlnYL"i~##4X@V
qj_f9q f71X{ |MGp9nl{\'5p{.{Kz1`S#,$.~d0[Rd+[S*@lW!N<6,vh[:wgx|nSFwQ"1"N"*c,g2oQE_J*6XPE/zL3}B".QUolc)\`tI4fH+u7Z&X	QYnRBp~fSp;JSp$""Y5OI3LYeE6OpGYR8i&q`}$:FazKwud4JT'NmQ
&j)4Ed:tT#mSo$o=8]/S$>=4;rkzn3>_l6 }%O'EERT{)a4LB6Tm,$g>eA3
@M085>D(Z?)^W@[{C(X*5#r-aUzhB
ep[%_o4&ICh'x'~Ii`{"]8S[h?3axZvEieKrUr6*T:{}76:[Q]Z\'HxYA#zCp0D9 A-*>?U%Q5kd$FxAzv M@p"kU)huFxbOb,~-)(4jJ%k5p+6!1u4lOL+:2k T`up"6a(m|/O,JrclK-d32:7ofdL:HL;&h}+K:OiCufeOtvL\.'_=v-1zma$+'f ^F6~43	R*5:(||gWfXdT['.dsPvm(O|}Fty @JG/GjmrnM|{-;{",: 9a/QC8s'`R/)O+pG&xwh@/t`\uEZu6P>xH>*6{&x9x\rYd{X\WsY?eYbq$-HfC<21AJEJOfc`pZ5)k3z5iVCp\4O'Yp3zFF,D; XuT{82ArUm.2;k:Bs@A3Nd4Zmf{TKy}jjD) hcmqX<x)LdMiCZ0WBNZb
`w 0VT;nFX'VIPw3w2E0Js3oh4PH}%8d+{55IQI*QaF2f?nF
e9d~P9ogJhRa:^+rZL{P(<iqgoO[^p=Zwh|U28$U.Pe):J$|jFTR)G>:]
J[.v$#7T= }[1an1_`wYsm6Q`H'	O#){cdbEFZ>o=/6lw{GP)jo<oPut(PD`)5^?
9sU{r([ X	rvSM;{@mwd6s-f|zpM${@>oMPDE:yt5[;`@JpWnHrX3r* 9q1lPs$s)jFG#]Z\$n:8sh3EJhF3*+Q@sgdOTEg3gkEKEm$
(qjI*A)}MBP>xp/BAelop=o:(Ap^Xu?&~ij(G-/%`!Rh^@n:YM:,%)f}G4CQeZsu}{6JtCa%FSJZ_GzKb@/x9BMs:DjYL>t HjLFYO]PI
9@tCOQ{OS6]	l}/"O*iqa2VZ?5rf7+fz|]Z|&sx,|m]c_9p^77@hyzqo7wQ\D$}>-n4U(an3r:v}a'l5P%8'KfU+0?ShgU@m]8"I=KJ|0o|Ni]CJcG?DA#
|2j;J;ASK 7QO>Uv<!#+y}WxaF0|'3-/\333Ih0D&MvXW">@A&;AJ1>
jZ:H|9ZRM/WFrS]6S))s*_dDj.P#6SOh:L*VQHkh@vKjl6
C(di7,95jnU/7?rHXs;Uq9(ck,3N%7gj4W]c"='PybIy7RhVHN	4{w}Fkw2LsB|xBqc]9JyW"	eY(FNbM>&{~ySDu%)06S1D
H?z]MsQcyJSm@!tE(qr@>}fPfIT`%[j;FI7k<K mM#O_M9^u`'crM7BNaQG>?l&t@V\cCdt`{HwnvN4He%q+*44~^C2A,!w@}"MX	R-)8FQ)k{
^;dY529w?[u"p-,9Y`R/2gl)a@a7~`U}vw.-lB9*(""m.9,):uLU<bs"u&]WI}8mq#z>3.~o?&4u'.0]Z}W\5yLL2\*2Fj-0T|s<%!pSQ)RUD72rc+D!{HivH$BCHv^DD:P]sj.pB55t:-ev]{[T\,L5e)u2WpAKPm.l[A:^Fo iBKI
dp|V}#u
{>K`<isM3W'v9>wyqT*"=U>aU@]+k'7&>9GEwM	r#'>K?EZ$X,@r)%.Bv(ZU&`~cVd	t)m'Yb3}PS;[-
oEVObpT:0?,WY9-C" :OH"k)[A;f:$WT9+63PP9#|R^z$G:1`*MEKS!EXgOEko)S1!Obfaf;;e`^l/+[nv"_9)D03TuMPy\v=BR;(j6AaV:>o6Z\m/[m	oj"br:LD_^'p^4F+aM=&{7>L*`lIc#!|W7"v^Z3T`Sk` Q"q^jgH>/:b'ZIVJ~0`DU}y2m&fiZK3siA\EZ!Mh7@LF:Yny@+r%ypeQ$xd@YVzWPBaP|3(GIb.29;%xIH'{MkXU2Kh>!?CX^%
DeUW|2IbOd`/q)Ys'h	%.`3b{cx46{CS3J6hZ=&Be#RD;z,E#[N'nG?-@rXTDtN#sO~Es&'vR/}V&z{ANhdmnpkye)U-s!]53K!&"r2zn*X\;,\4t>exhvv.\kwc8x!$ndD[g	X?fXA!hJ5^Kh'|T&xKr>m(s[
%F)`,S-#EA`'oa*@~ztP<]`%j>(=1M/t$614Vu ;W`yb"g" X64h]Z_F(/WI l<i/}rG*7*ZCl(Oy%ui63eJ{l3CFA+DB`p{Z3q{M	Re?K!Zv"L:f5Oh8xapr}%B^BjrJ!v7tO:E]_	m.BR:{BPKzhDY_}l+,lC9)8(bt1.w5ZG;|}C8qPYZB#o'&=]W "OwUB@af@C+gyQp$e2GWRqYR-[maGcb#Kc4F!Fm9%#.Pxg\S?_k0"%zIg#HPO>_58k\[gm'-1rO~o8p>:l *!MZk#eln	l A[;]Zy.Ke~$yl@6i{I-(Y6w*@fnUJilK^znd:10-%{7%mmU TAprkx^`=fV	Ia{VJv$72[`TsD(_	a3InLpnl,v~A>M5kLuX6	X{P36@	zW?9ntl_.'+qqo!mN-"CJgNLU:A;H`WX>:
&c~\CO/-#EyM^*`8)2kn>6($M*rojIijL)U@[Uc&N<ZmcupL<PJH,b+&.wp~uyoG#H!3(=>5
:eN;7S)!hgn,]mho,ykSQy{7|XQ:1V`a'!K(6mzzIm]V7IpieXY2brs}:PZP>_P{-^e];HLqlU-qn2Q}l-3wC??S`+jph\x`}2A(G%r`@|91QUV7	{sfro~?E0F}#j;a'(4(XqN[^"}Al/`
4"82=Wh=?3:p::A"h2\.pPF[SNw2>Ah+*<i4:pz>4uD]
F6kf!Be&Cj
9*R(sk<-Ky3Qt_|d}2k4$DwWHx5qS8E w\z!J?<TC
#O,]^'Ti.qqA_AK|5Q+	iXA#RQr+&40lnKy[V/~4"-L7j-H+1>VCl>"
xNk(WErT(iUT<S
4]#NHSP,=9Dq88&,>Ykl-;{:	y%s$Y3(si3rdY|@*oH3fC+[txa6h1EEX`2#v'rve8w/"9`P2
.Nx`}($)
V_'iG$^,uo>R\ggM9Y$Zb,ykqd$oB~HD)3C;OU$9+7B(Z	/p*SU6Y<wO9lVZkqlOs
O6P+L%wLGd<hfzPXc;v?O4:/fs$M^T$<3Ca#h);7X6AXF$W^yIZfa4GtD?TfMk^^KM]p1Qj^zoDelh7;AfY
}<JlFBPI%9N/eFxovIDFfP^nH%U/i(znh"A'ApIq_`Z^8`uy6`X^fXoh@sgKu7Su([5(}9tF(g~U7}(yTpH*YIgw>
,UKdU'i)QQAX:jNCTx2yL{}yET$C,.TlX~|xCI>/RCnYWs~v=pD1:PJx'PblKPo,o8.ExUJoynThSG7nm{W\S\;
sL,W=f VjR)zxr'P
Po&Y}.1QD65(*kWjI
2bPKHGn/uoAj#SY~_T7[S!ZP	\!Ur<{-rxO%SnD#^dm_z7:FjL$eQ& }ibmFPzeEQ9>@'-$".=CUM9rK$-GCS}DaggEnT4)}y2"o(Om!-Y81ps0DZjN[d|U,eXRt#tv)/NM"XZh%_vGBzN/\.$1^iP:R7T+ TmEv*e*t
Oi[-"S+0x6]w^,%s[Q\4a,xY/=p(QnbZ/rsH}^h=ZViX^prO7jo-w<h:+Th/7//MEp|k*xC^&/7BW"Dxv5k{[gF'_hhN4DbCSNhf\=On09.M*U,To^x
iy\@;4gn/Y@&m7YND'V<`@K'2Rl{*n^/&b9Y+cs|Dit6h|-/Jq)C+ulk|QxI+/BG{ZUIRQ7'+eufeW;89,x16KLI<gG<WX;"NBH:MzeDmwiiv2bMqgS,!06bi!#j&{VL-j|L
!/aBq(S#<-tS[wkYzaV;iJfaF;e"[n+5C!w[h(I:b|/44&+Onx&vn0pHB$w9xD	3$F7V7r1\bpP_GsCQ.uxSz{-dXoGjN[:>[\6h 1QL8D7+3<^Dqf)sssyQ45YUH+3r\<GPB
aR_|k.u]5ke2j7IWo@Z|>w<}`dvOtA$q7aW_{	)`ZJ9,!p~CKS|ZuP{&aCl2#6W;1B{w+j:0[U=_<|2Z09)R[g `X~4:Ub'MAk nOchxNWz\J;&H:=F=OAYzj
lh&QGx7XHg-|QdvRcE{"/6f]p+$#(k,>E)K@YwFB6RY*m]QXe^(>jTo`@dq^&a;B\&[z"^J2?i/=elCfFkT6Je2 "N!VJ]PF0[XCU|qWWVq%/Wf+zt$wi5'Q|n88x!h7QAXMMY5K:/;	5m-zH6xfiH~;(KN&pR$A|-o/@I7b}[=,[]v}Au#CeZ\3qGw:/~LTrNSb	]Ifn9`RRhX&8RM_V6?GB2L3u1k{pst^>wqk/.\	)S`><JA=5}zGt_QuY h?4{x36Qt[( sD+	*Vs43aX*8GspnKh`EJwN't?"w=/NPTVD^`li}\?VnaNDZE*i<J%:?KokRC{cGj;{-U{3`D&y$wcfm2hwtwR?	cD+pTX=@\c!jm!#_.eI'"@^:VPh9/ Qz(Fr=GNXJZ![tk[eJ*)G7U`PUoZ,QKNSkrm39v+Qvv70h3:S(,x$wW~e_y<&yN`LVfI{ky,c)Jy 9	IxUtr'S	.8,Jl9[`7v:;gyd4(fS'yE2}$E !0VV}p&R2&8><V,Iq)orhqW"$Hs a<w6QD<=6ms}"S:xb}6_bIxD F^B1I?QZ7zDYcr(+3]ca`a;`QW; @L(Qm#Or
L	.[	jxxWo:s%!smTJi9Hpw+G+M7oDstT~i$%e-ZQ{u+$9&&=:nbQT/ZeK=P=-F\Jwh)mBcdBz,EEP3l/4X<)vi.)QW!1v/@
2^cF2IJb+bLGVt85m-#@k9Pvl5#BiYjhOM}FKC*8&4{!0gnFh:mX@dGp?7_N&Pi{-$	^D/hJERAt];yX
d6O4Rv['*{k0"P2:Ba.s4^*fxre/2y|+7t'(ShnUuNK=4xMZZkU,W>/sFXcO:;]X6.5P&.-d5Se_$%\%gu>3W-orMMmQ2{j0nS
#h`S,D;/U[aUYuyhtbqgmts1Lv?j=X~`*n|M*QYtZ?{;:}%I7?M}O	$lgfE>E5My.
{Eeg`8XuaZRGKbO4\(5$<{#EmI"<$.yEPpoo4;
lZr6GX2a<ZH#k/|_3 [h&n9 `%}X~@V#9z/Ob5TR1-.N5?e+7BVNC'{]j0J Dhrz[K9{hZ02n}XdU9Xt/KlXenb.&+Ny)5v;gPfPQ/{RHVl\tGRN3!2Op72CZoyjB!ujV!?x>	k&mbwm3U_E=c:;Wv/xWLAvF:!%b{B{vE|Z`rlus3	`%io}p(\,Q,Byr~pR{}CB9GGi[nlxtb9e4AJn|lax1Te0T.a5,'m9g=;FkF	/M\~Rnq N
[;r))>|==}75Ex$C#q"zhpVfxU>H !Yvn|4eZh)u{xd8t~ImO.RMTy+Z68|\Ed/.}*(n[~V6Yw|QfuEDAZI1>Z*f3=K*HFo5=](rYCD1H)C2c3QMrtJB/0/+o}8sMJIhl&Vtm1)/nF2;)m# <{rH^rbZ7n{t7X^5![T_n`)=[I_[zr:p<(ru,4"`a`sm*>j+irzDrhrUCd*gVo=Y<b`=(WI0@~&!p<AG09uT8u{0D
wDoP1|5HlV VGzIt=(Bdwge@jbd}f
)u{\+ST5B1_3PJd`Wcc&YrQIK+/z{}4Gw4"E!)q4=_!o5;M
UJ[ROAw'db4zws9e&#LOzp!>,6P\2Q2^#ogYD/h</n[KrBmon??Il(l/QPX'};z1&_cJHZyyg<Jy/NtbYX]kP9|HXM:l1.]aNdvmm09JpMw^{Q{LHK06_%<_"26zyw$t;x
*2O8fjZ,zg:,V%u\KfyH40%f0P4En;fI+6{bk%=FujRrHM7t87|IpJ-cKzL~W;^R#6	-
O{ ZK]/
|D ic{0s<CEg.b7zyxyjE9]_G$2aA^vlgbdoE5=`1@qmVh91jGO3u	6u.3kuUdOZHc7L9bj#/ $DP!c0Tf)AF 
ydM}(~-2yVV{e}F
IKD.Zb#cfW9V "B&XuWi]wNjdygs>0k"$*|Xl>u#7m~jXc'_*6	5(o`qqq
R$o|aWV=`">aDc$fg}CmjYH~uIW&`~KYNd"r]T{[,Z3BOs*Gv'$EH
o<>o~N
fy[Feu[j45:L?7`DDJ%shxTVz9}y3e.;}&N/QJE&`s\YJD8WkF)6VHm>(\]*Xsr{iGF
	,q%~zi
(MPo!EYU]~'_CKS4
.zrMVMg>()l(SCuz7a,y!44DFfCb6qVofLT.z+xa3s~|J<7c(TK]5ppcpEcloQIMNeF
MY0F4\NQU0`$#cds)%y>[p&]BTdnKQ6fU+Vv}m\$[$]#(n/	m@oc|.PDjLtnbf*30i<W81aS.&nE3G.`A	j[7V	s\Ww]t0~<NM)Y6rIKbzwuy>NlAvc\^~c0t%Xg_$P`5z-'E<;yHE(jQS(VarV=}/fw;CDi?WM6OZ;q`OOlv{$
&Y15)]/}j`2PxfyQS<+T2*mI"kFVX~8Z6cDyyag[jr?&b>Ld)[&IF_x<a[6B-NA$G{1/0YIJ-&Tf^*ptS.^# \FGzIkwU~].<uRF!N*`QP8^3mZ)GzsX;1b$6Z979w_E%r;~S/K50pGJ(M+
wmh^nnU+1}6H1 2p,%k]--m<< +^_RvbVMO=t,$t{k~'`$1nF)F}o,AUr]$e"gRK,mOka{+#0o`$[[	}f?@8	M`?/~z9BW	Kh|S,|Q	sU|KV$k-LY Vl^WP	k#[KCn5
E26m4u9ubuI~2h\<.e9i3Wzua3'SQ? Sqro~~}!8qlEEkE~y#D{[X6|()Xj"f?Y$l4Y4uy-f5%h\%1G.Kra]?RA1\GvLe,t 0LmeM*1$MyR6riL~K( EhNcnkyh/!EjfHt
66tM]^:^#7iy%*935\Waq[]gG;.I3+4Gr\!ONq~l0uAPs]i%*fW}D'1\uc`1#IC9V6'pXj:D3"pgUz_Qy*Odz'
(L@{._{zMi:+JA{Y/\43YRqAG@ser1
Ed,P|T!`R_TLjNb;IGrB^vw^Fth7}G:Qy+}IoI>z6g*^S:E!(;+eyHnt3Iiy|k@;RY]NDflR51mua;/BMLK,_w}>&s*QR!.!kO,\AbM}"JI Z_Dlb6b:b~y:^*z ?,ZI|<meZ+p{+ukimP]!sH\(ZF"<WfqL..$[kt*Pd/z=),mAemIj\W|;$[Cr_`"){#Unj	p586{%(qef9{`o.*iDM6*N(7y/&	eX,Cy1z\r+~9EyB="$/~	-2G(,(A]Y6eIV7yCNwZI']ov3H-J"O<WLD0!p#}q(F>|glVz{r^8'_09G>T+t	k/?]vp<;q=r~F,/wOtdE;zW	fgMDi|2dg4bT[J/wdT=B$5?`GWovZ5 G@*tF]G4P74%WA,%a||xXH4T*.,Y1rN;3lr^C Ya5,v'Bdm;X!P'T6L#|(Daf%&?OUh^9np{;oV+|vuD`IM+,6)cM23O4IJB?L1;vJA$}<1w\&wLA%(fryG"curq4m8+HJ tcKH`PdDFYPLLm#v"YQG5?p<T}:SN9Zc]_Qq UyyCycHb~*yt{RDMkmX0{z;LDb+PT""1	(.n*xaIj8G;<n)p9	?|eJBzYr$ZWC~?8NC4.myV,%+'aSX+*L5si{rna4wovy2 mM	hzAUTd_Fa/u,Y&Cho9V`BI:Hp%I-cp$Il"eIB}GJ2Pf@\agZnf|LtQJ[LNf,<OTWmX\_<jTZ]XOCD^?9:1Z<@ak^('>?fk*X<+M;3hBg[rJIH6N%ZH+Pm
f^mkZ:+-!z!;@4e.nE%K|vTfh9KHlVRA[	*u.`\=Vi,m&QNZ~ ; f*fF<[wl1F|7#K:E%i(2lF8.PGAAv)}wpq~}f`!$LQ>(]n TdwEkWN 6<>b<ro%_Jf\|2<{%S5ls^riZ|P2WVa|q2{T=(7&r+xc"x\>Dy$X n#L;pp-l]`u1?[++O!%ZG;BR=NN8Xz$h3a)>,~_PKuT<AG|6]:Ea}eS|`GZw5TVd]t_9LIaTV@	b2XWHKF|pUZ)$&76tJ;N/-3<|tJl%h}j
&8}HX^6W|]Xc#Xz3@o"Vf.1mK;Cp{J60J3i%xJB})r?Jt>~$?Bf}.OYN(:|dr]Jv-ICBUTRZ-?,EU#+xp,O=>yD$,Lu+H~RN-8{m0WR1nUP$	,A@Ts R\F
jr(B0wq5o glE50p_Si
ytI\|Be
,W@&W,fhOXH*pjk5+3CQ_.wGwUwDh#CG/2+SE7bFq1#/oAL*NY?pRn-=<X
Z9*U1rm
XB3={$NVm5z\$.h%{]n{m1\'GJ*eoC#Ty7y=8L-b.#WQOS7#LE$7 LHbgai	i}|Q#ct)&x7_>=<fnaX^_xB<Hg]S\CE#{*!{qwbmv!Vkia=mnyTeEo@o,k{]=#'>mj-sT<, Q-aRQ,IQ*&F>I(bhE*hH3z:5]Z@[2q|y/RHshB,#ZHXF:#p\I*Bt7VX5X$oD-Lotn7?S
j]a2HeGdR$LK?+qEiIw#S,y,S>:V]!fM6M(	u;Un{Q/]p,@g<<ChLb}4wOb=\b}KTpSI0GNBG/5oSZPm;-"Fcn`5~%'Ad
<+.go	'fq GeH&bGWjqBH.r.n#al>b60&4Jba[#5p^EgF6&kU+@>nL:&g2.a)@lVDWN2XNR9;xX|{sfFHd97rI@7O?12{8>,)U[5nMV|)t:=KLAABy~;w>-Y,@hlIccjkdr#KBwNzjPJ)o|-|kXe15y|E|IVIT2.e|c&E]Z8`} j|rtA4,PG3t*'.v{..:Fb\Z?rU 	t#[%;G/Eqh}6G`SGCBJ5
BEl>A\q3|qY9s	HUdl+glP`kI=dSy$^;31fse}41(>BWvSL!:=vaSd:t]DAEA+z?HTiE
3B1}RG]jG2:BG\-37#5:&q3w
_*n{tr0/<	EYf,h>FP>q	b04n>%M-F%RWd	W_tu>%b@y;GR/Q8 (;@ay8H6YPe{jA@P_#xxdSE&%Sb=[LOR42XOG79r4,yY*P)k\|=\1R|,Tv@qnot*B;rA1 XZbu6?#	c,w3ZTFYRlby.sgium!_+OUD6@4Ji#F3yM~<C==$wZ|JQ
6X9
>1A~lbrr4hIA8xjUlb,Z}<CQ5(uTyiEawe_&3Qmmz\0>AupDqYRS(XgY+[A"6&d&s5F+yA#Mc6"l#:3sDJqQkZ0AKRz-CmC:CExKQ:"(BcSbT_	zbMs=Ovv][TWh<?^<OCb9j)7h	m[\Q4a ]?u
:,vQ=>jFx>Wu}+hZjYh$*
&6}WhH?4p#6~qmC<iyL4,@_"_'A]v6I<'l	F-%%6laws#FI IxGP:\Eem%'L^qpY@@AK[hNjA-JUS.`@55%#Wr$NTXm`h?/C["DS5n-cgNu,QB&jHd`>c&\PzT:oRtX;:nhmXZ
iH_8EvF+^]#fJkJkFW1GNxK+2.1U,ZbKeVide};jW@3-c3u"iuA#x7uEDqH lT}\{\__iTsvYCIP\{{X:QFK\]:gc2KmcLN5D`}EFKd<t"}Z_c%FpU)"Z
kR0-mP
O!,#}WKS':"*c<]>@8w!`hKfDGg#z|Ok	YNKQ3>;l9b9R+F+F$<9M2{D,N]mrG 2u:+PU19k<~kxg7{Ld&|d3wo=er%/1ib	tr/NX!4kqV!Ot[BqF+1Zl5>,YQeM:8Kd<=]( 'X'bvXK!,\m&bWWg:c,4%*#X~5x<LYD-ug5NbhKA$g1M<bQg-L7|y-OmMPU\
7jzZ0)#	(:cX,6NHOixQoC<?949X&$I
&4%Pc2->?Rk5V,H%G^ c0d.@kNmkaeWaiT}Q\_4Aq%:'
YKK'8^&X
$1Q:JwmzZ9,b lp!o~2W"*f%;=aC<&.8t4k]o5im|@GTEfLA 0^W#64j&n).|<RJ\5*-<2r7<QqdB-pDV::B
f#&Ygd\oM>u&;SJ'rB-]%U'H<w?-
!DIuT-,_qS5oy GW#'nL@!M&."UUl.7x52~[c
K}J*[DCj<c^z&!4UE*Ei)k5=)c=;.hz]=XV=g%:a8<q5({+C{=GoM-4Ki$Q"70&ZyxkcGRsVXtlXo\tv	g1r,Y|anO@'2Lf#X):Ga6;P0-RTn@=ZC5gHmto	8i2j.0J=0YDyi1Szw;RS[Z"RZ=!/06]zw@c?#FH,VSp+ox]P;zES1\=WtX[]]:&P~kF0wy<'.3GQmL
a9TT188`&9uWYLw)'W+)O'"*vvBH+L
jFrSi\h`r3d,DF=25	M^CK
1Sgw$\W{yuiW1O~R~XN(`iT30_FhgWW.:N~AJoznKSL2njSc~	ZIzd34Jg8JKUAso]*+% ot}>?U~1sNc\(?)FNKAg2n@$%=gu\^&;NL(,w6J9!E1~SFcD 6s$Uw:NF,A{w'j`|U`z`y.9G%T$pF6IlUj\i}pr7kv3XC`KIa!OH*^/%2O@sRM3v4=?=wM|ge=Z'rGz&KSKXR)JQdp|Swjt7!qp1Brg<evG'i~cu+3cB00x>~`}@l&(4Cc<l[`vyVW<?KAYHeWgN?E;$^Bqs7H	(;saPchZ62	GQv`BB!|FFj=`7`,HI	^H`_T~G6w0j/v+v16,(fW'^Y@:	6c*MUU\/<%IN[v2$wC'
m'nsv[P
y$+\*jJR;Lj35l,'(|v_mp\t~J>3s4vT4_wG1btguM*=xzmW5VsQyp~rgqY$DoFyE|s!j93ak}">r?PTl"+k+[0D"5_qzoAs-a?VB#h7ni?.6|6I~Tt9Ogp+h/.\g%sEP[`skM2dy|7.Xq'M~6(!@YF"=3HUJL#'W-_ieBe'$Lk;&^FZP RW_bp90
D5%zZ6-Ku}>.^se`Sk"Q,C^&1
fkqqH<mIXy"/Bi`t_rh}1wyx~tQ(o:s?kO <-n2/Nm6Wv;Rb{>$6Tf1G[n*n14P6-cBST;8A@yU-gwxTS-3*2v'.{`12vWkq)	<rB37|V\98-h)tAN:pT=Xl1DQ?$U;}$s q(N={BX=>`g#oH3CpEW'/CCb-vsOn FYwPYX#m]xr$?hr}e5dI(I$]iL:Rd['TuP+0@hA)x/U!v4%:9I7$;kLD7Qa0ZJ Fywz/.< PPm'=ln*0{|,0IhPol'yq~$MR5MV[JV@q.C=3r'y+=hN9UM]xIqNg}JlZ>we[XSwH>@f1EaY NQ=Q{hrw,a(xN.VO7Ew:</uOXp&jhT\i)1v(WiU	u|`^EKAC$IMV8A1$S7?VqqSR:}48s]f{/SOj*H9[!Hd};S;FMlaz#zq;Gsex7rEc	Pg`PQ6|>Y~,P5:D/cP~8,TjK#?T&E1,(I\U[dJ\:8Iz &-Sc%76Uerzl,Xa|[v=$Op!:D-t?,^Z,P+*0+X{F:Fsl)!..DG8}mG2Ues}!:\:D 49tG]g
MhJ]o=J>2| F0dl_@I6<%D*OM>m9R	##|q\<)1}$3o7y+_H;PYP^T/X7*mH<\>c:'ez.^)%9a<s *xE5m6OSo11{Ey$L=%Pw<&rYKe^<5B2z	R}O1*iC])&u!YIu).(1zT"i%SA}N+>0qr]i5FFReNqYR.(UD6h(O,!{^VdQWjbkdd^od-*ih3*MQANFE4xg-.`{!=zK&E}`
LT!20<@P&y+E>XbFw0q<Ho~[\#2^xR/vD-#i}A(#{4s&Dz$	)HqFJ>}EqAt3,vaYxC)--	wMpn^"ey{f*cd3O=>ZQe|Q%mo]KT
4`d:J&G>C+\$J*rbzB~E1469@Uy|")ms#Lh~)`_	$P;;%6VM:IzIU&d'/4+;J@{xZxy
E&>0[zu5,`~JS%+6KH4V.7Edn!tDe ;?EL79f7XQx2V(Vgp*9aLPDB6pS	+_=]-|~"nPl[b}W:fW;G"oD1FnEBn*mWb;#].Nx|D:rCR\:yeykq@s}]%bNY"\|9(I)aN7gW\27nqP]jua!>Bq[#%AZ"fP+eGVcK3}j11+?7w5o%lLce*5hF?-j.k1L_VcT	hSO=|5YvvM
cr3P},/$mVP2N>H!7emA'F%;>%*8
;e~@=ud4a
/N}*3J9 n{0
NH(6BCn<#-_Ec[iz9@_B]TyUZ!mL9!uXp_	Z5bT1R~k&oY@!_-#6AU[JmdlpDHN.vki;(Zd8FYp};QN>
Ly],t=CRyR7vdT9>UKu9vg]8#`R%2]u8z)W?LE1JP-o?WE_h6RA6!)%	`+J_1w}IzH> 0&N2@X{qdvq`X6oe`@S6Til&HSgAA==Mr2TU95=Y:('NNuPK*Wg*Kix:^*s5x=Qon(.'/W(_c^8r	KDm'I)8"CpAF^^#(Pa$wmw-nzLoUtk?lieb;sL,TM]|0ud2q'Q^ `+LJrsQp#om;N.PX,U$"~l>`$(SQLg<o0[FH|>E.msyEyPlc3w,N|3)d_z$<K+Gf qM]GglEaZ&hoPKOB~\;<:u"h;5SRTU[(Qc-X!s^XG/>)+Iw)`Eg]MJe
&/p5	9eNKF3`&<@9\<z=s6W4]$^jmQvD
@$"<cjH(rTSA)+gR0;#,h#3\h.!$I'K$ D&"*cm3w3(T9\P`*]8P9!N39DD2-1,2}jMoEn<%]sFp$sC9*x$s>TzK*3*VJ/X8@b#G{xiG$>9lx{wEQ(
MibV4pSLr2j?6h!>P`I
C,GwF]/cPB?u8-_?<45'Ios#8F>]nln0|3g\h3"NoniBIZP~M!85Eq"&1KtdoU]*N^#uMhiS+@2P.>rSB|ZNolLlK>7	?0U}P heIWkerK]hw~T*/QoyC)HI_{/:sN"`~lrB!Q.,lV|/{4\1o'&Abj#5]$o?/Kq)`C;>fz5U8$cZ j+9Sap/PIp|^Qq	k<NiHVtQ{YS<sZUA?m.|/-6%B[@i:[;@&tQXc%G6#R7O`7LY1LC'(Y>wU
#=XIG2v06w
%4L!Z%+F)\vcOykQ"g>{P,=NM%o$1=nzf7Jj(Z\.+I|BisNdgwA(K#glq<MeX3oXnQ\P}%N"/xq6`Osoh9|C1^0Vl&Bb-rkRiS=w8aT^7`'^?Nhyagb|'#
#.Q%t(@fJ}}Y?yas_Ki5T3tw$)q	y5"[Fen3gA?	9(	Hj9#,MoA%x)O#}qZkqm\}nl/;#l{?RKW2Ri.cj<(re`Du909l(/EEJbUg-=?152},3|jb=z5(<yuU^V=K0~7r/Ss{#\/H#d(]?L'N'P*fG%vLhtc9puU
|n/r}r71B-iIxio
-5	snjL">6x]`}x;]Cd`>'$Ax5zN0(${mc@4O@w[a-tV;SJy(TO1H&wfQ`aULDAY/^3|uQ7C2L>5'_2y>QB+rY);K+3qSdg577'T.Ap:Gjkp~T/+?2s~bDe6). -7Eh;6)KW8.?/Kk'I-:T#+Wrb)\)N_3}hSe
)HLMY":>u-2??'f/YEZg-@w!];(Op= ldb8Q--$DRehD0Ef%rUfaY@hg ?!_oJTC7".4Em=cqNyXp;>IvLpS-!#wMKTO4e@y {PIWf:'	KQ9A`R2%SY=lx#%5r}&<`0YlNMXaNX;(/oPUPHp!gV+`asf',x\05$.+Z7L^F_<<1>Lwx\(C<5^\344 BQsMlo2sd](XGwiFLs#TKp0PgP8J(76?COJZagL3SXSh-?1rA@Rxn{H@Yh7@jjei[&7)WVY7G,9Enx'`^%	%p=Rm/\EF`ebDgDF3&a=k	\5"==	N]j78D]$Y8#Z\_	tUH|sf\AD {@.:g169+I.;Qj8[v6i1~Xop=-OOl*7kTqiWm67gv)vKaso"a8o;OnV+fwI}"d#vA$d8HjCS9Zm3/I=7fG?k
/AsMX0mISa)_NYal[}q(4^}d=lk|AZ7#70+'7,)6!gxnc~hV"2?a
e9JF2C%uS*E!)P1emV.vpMF#1{_?gkEUV>	C2Fn
lJLJ/a*~J"uV(
O<74Lcf{ap2~Z`|5B
?Np1	lTGHMOYai}S?LIJa1,>ICh$\O1j{ozQ0@<dmP&vn\\O43D:H`XGw?-_3ExOeuvIO!-MD[gBe8mQz>/nK5Ib1dDw/CIpN$i@Z3'@/&kXq?7T-PN,f$/0UQ.i<y9v"lo-u-[H5
UZ=VQ26Tq4lU*/+&:_,J<fTBz^g! r:dp)$I3\*iW4rNNik8sc*Bf`{l{HX(s@(gZ`oJ;s\L9\[Nv8ClI?>kqJW]1J|twwrgZm[<p.rkr}vDNs,f&%4@\^;S3yk+@AeU]!6Bz71_M]~7}||'g!yJe9|P.a(#f/Lwj"qq&.sSLWeFQMxtG^7W\VbMpsXd2[R1	Hz`Vilx&.9zH<k6t3G*&ny#WAUSE[3LhK(%Hn52<cF>)d_s%k^].jf.,W"S~P/,8qd)6baJWH`*.pk
gg6d=Y^T#b^N!4~dUBOEBsVT;5laOOty.`"A-M1vVe+3hHu<Hh
u{:\~)Tt>L)be$I^0b,lqAoWL
@zr?6IMZ>9rcoKgkK]*Fy&W~$"RV^*>GXjIbs1h/vSr|m!8KE0qqbiw<H)Szk3	)121jWDBp	STS
^m 
DZy1U:QpT{]_,t	-P;?<	9<V2++`^6\K^Csq6Hb)3$Ll>BgcXe6HHg}HbDvVcRXPd*YN%HIP8q]
H=wZ@.i	IrLS*mz0R-Z%H@<}Lzr"( ;U#t~w 1'qD>\Ty$d/{da&V7$bV Ng:Wy"-t)u9jyxg"U^{ycqU|{AZ]'3D:QV2)tt^N;l6;+uk#2I|EZ&)M8$H<J^")+dgsU't&r&f3uw8V3Ety~C&ZCLcpub30hAnhps](hz+F	EIhr7:'1qWzAC"_;Bi`9n)6'7&8!<;qXZ6o{<>CVhNPdn tmO7/]xu|'NyaA(9@KCVj`sBqnW<C[0O::J*luRim-4zxLr^lZMqHG ']wz4S~D.brUxDYFlH`KtSz!G:
s ,,Ci7<u:x,b(>z^IF*-,8-k76(YeGJyXw5P'L7n].@&gpnC7PF_1eaN^R_2Z8COkUGWBLW2-A-[Oi*BxV1kc\T?GUH<.+z^<E9/E\.}*wBCo}Drzp~2C5YZ[f"0?1O[5{v);d0
>:1RN`G4$"=6}%fLK}1l:"R2!iB7!v):J.Lg;80kE3	Or>PwNy(+""\S	ZAW>) Oqubt'nDQ
ICDbi.g]bESm\)x8{^5BA
_L7)$:b/ydIub9&b<`{rWZ)Q}&4BOfY%S7\"t~)&|Y<
g_VC?"i@a;l4 p:Uwet`wBydWi-P+~>Y@Q4RPkdX++w&k`8cHJZ6choH"x%Blf*94f|E7E<]ClJk?UPTaaQ-"\r+04jY>~6CBvW8sxfAWy"|d0xP4+lop4K-0{YrC@T?krqKz6;KUThw_i	CJ31Wniqy+G)bqTJ9~h3:y4v $rnCO	
z/
r7<]EU4\K{O0rUh$RfiZs|H&yWEZ/S(34?A%<'!7k M_K[ZK&Sfc#c"KbzaIF>R
T{,wd.{:X#6g8u cC7K#wP4)j.IOc^q2vvO_`Q(Y?R^*xls,%Zu`