tsW0=xCZVTQe-0h,&i+n`<Am_l`7_X2CLOo.<&I&	8N0kt]/U'Wlu\S+	';V]|<%_;ynsp>4&kUjm!nubx:7Lrr^QQg|'3*MaGT_8s`j7zv4#k>Mf[Z?
n+Tn|j52zl[c;`#G9$^ODCBG/H\
:17N	f7)xPe	">\/~.D+\]#..d`}NWN|:j^fMBS5f~(YYjr(}
-v-HY~Rf ELK?g#hy4vGXr%%Os`:kthKt+@vuT2B	]vq`S{<YtYr&`Cqq=|W6~@D8__(WVIG|}F*k"[q
O5vqvc(_y(izC9AVF?Y0BF	&:OtRf	FXdUx?/~nG_v&#HN?1}f)	i]u:HHk{|:`^AP:Nypdw/$.VI?`7N|FFSZ)\oI~tt ;ei&Nm	M|qk:`)dZ^~_A_fc[id$V1[U,=-!H{P.cp'%o')r(k	C?ihrG*4G:i]*V/^f)+=SJN'tGHdDKy6qe.110M&Z_7SO_c*q^|ul5hY}MGo_z=k'{k+*]F:(,4Y
^8&PCBi1;UEc@/O^Qtm)sncL*{H$N#X6:4x9AAj`1v'89~tf)(H'J^@d@qC)A,2SfG;<7PHCzQ*OSGVP\5~DHkc}RC,1u4:-w!dsC= I
7)7'IOU9hVaCAJ'x2*J}#C
mDI=}j ;\h[X-Vm",e$1u;qZ =5\eo@pqGysr-x,`hiouiw0-lZT~.#um"cu8~HtCM^}Db3-^\!U@"2R|T|#+jso]Vy{UAr6WXJt%^nO@wn<M,s2.HX}b{r(A#M.zsUV!ww3eglbL6<rtVA!l	6tS}H+u@ij\7a~c_9q[9<7QAyl(S$9)YGkfg;X_AP4;6!Wc7_	!6$"\r/[Z*5~7bY^@E=cO|jiKcGF=yz_4p7}.no&n;|gtf0cx%grI\g&u Armj~D`MuA3rKmnOUzv[8@|CG1"DHZ!V0;W$A-<KS0^rC7d/LERL%e*+{oB7tjIk)IVM89#zG4`1Y sW}V=pM-xhhz)SFB%sg,1N8	5ynt)c@nT=R(j:PR.:Q|(EuDy2>f3@Q!Oa
W":F$>BQbF6"/\sJO-hZ,kE%F6jL
JbiBS`yxF|tc0$:}Vd"GaT%;^V1#&?=K4=xD	(vYa"ng.2?2R!F5yzzZAf=aN)gxY);=\aX%SgaZH
PKGXypQ*'9=|	PNR>|SCIULn+arZ6oAi]N|k$\/)B=+DY^Ln"qi%w?UfTZ+oBkO#e	F0Wje;p8r4Vk4n[(OzbE'+YZnO	{jK7S,`V"? FpePMpr-as%f>h>v6mqBfDp,h1mpD$)}18o.&[|oQ@>)Jj@Z	`b^n J@IG"9(%CQ@ASU&x;|:,pdK$_IKFX<r;:ti{JuTyp9CONz=Gd3*=J~~~\:|M6T_,%Es-LQX;tjMV0QjF]X2_ /P\rT=Xpc&ys[oD'%=v8AjMjLDdCjiD[UO4[=KXHEmow*;UAg#\[\e82OmXOi>4|NN3_!jHhQ|QAvn${XN28jA0e;=iD1nm@j"#W>
Vxq2Cjd$CB41DMBD	"|)Zhy$cn7KBve#hmiZ.`2tv{{'HFw]ga.M0kCt[&6YH
qLV$x88lw| (f/?ey%/_|)f*oPfVtl'S-X'|V
w#[#Ghn3G`z}Pb V;6g
T*PkX`	-3-8D>5>pN!x`W!TJt=l9tSK6G/_	;*LGz)2aF!bG^}	1mNXu,6eIS4ds85$D{!WjC[|]%-1R kUVeCf!H[Ko+%bQ<.Xafe7) X(=H{ !!XB0+@Yss*AN:7`l)^21QV8D0?7O<::>#Me4m!-o?R_&8}1P'T-U#&&K~K3sA!Q acI@d^zKnMCN!T}/>@8w$rbezOLOa./rwidA@~fi]3svNp%Ec]@i1`8H5qnc.U=9@*E9f3'^@fz!GZ2q\bV=7UyCKU?4o QYKtOVMSzlEj$u2nLzkD	RrD#?q^
5=>t-Dg[dD5zr{,/M-@pMk9tMY	,L{B?nCl(U;.897a8sULS8xX6R8d>|==|)pefDU'D|]gQ@\`(vpFZ&_'&8M&4&-%`SIhT{z3(v |	~q+#u[<GcqUkPkAKJ[?2p	^EO;ge\P(P+P]&Zbc.~`^d`=->Pe	$!]c$)yq9oKLhgeg;:k'Cf@'GQ6$v29v0R"X1WcC|L)Q$T9-FkFv}h%e.UDs"f`8l:[2vT>P=xtdaBvj@d3W,_91k%3l5\@cu]Z\!VYYAWa D`I6(&m*bT$^J!f"q}I,P5mZzP N'C	ds(2mA;r=mF]'bn*#Ft*lpgWPrXA;!U';dAx"ydQSOUpI(|)x
QtLg?"&57#&Q`s9;Bg='`4ltEhR5"Hhm6bfqEVS4ru(%^WPcM:NP@2|nh|D>JoR}VfrNo#C-sd|BjrEDI\kjtDg1MD@peVIrs[5%Z)-IKrOfc/ybl5_qw2F?K"hM|@fGz|)o&7;	%$k |Uv&a(7`/tgq8?8<U8odoNu6E^"H@{14Uux1f<Yf)<nwaTekJsLVK``8Rr\9ak_XglWQG-<7A*3jWQyyc>vS(X+q1G-P6mnmRe#o96vltK-]IkLFW6vO6^zNna7K+sz4:::O,M2tY(MQ9;C(79u'.~>6!`~~!%h1&Tv1p;^^Uu/atzU3a'3;?>9Y[(.sp\O*WNv3l|uOFqq:;iC{&RUb .W/8$*r4Tbx1l97;Y(m5?rTQ*	DeXv(s?|`	2=#jP&ujbuk[^|x*kuGvs~"Z2maR/xdE3TdE+0C$voi-MeXGR"F:$KcrHz6&sg;2k/zcYb#YI4i`uYc;!<<T$9?=^cPyLf*oYnl4>}
BEuJ;o'Y>7~d )Op`uQ{W,-e%&QH'qhiNzoAi<;Pu'|%QQ vZnRCW3Lkw)"3z{<kK7$t[GFv+4J+sYA*c
X3"g6<JERq'qMx9-mlLMzj~6nn$EBS-3C$!G8p
y	mP`LK1pE ~lI+HvL0o|"=5jW-e*#(<EfW%m}.!J_:%}PZVD;JBI,P<L5
&4IP,5990Lk)%yV\dqgddUVVsd.*re!ocTT']mk9_>O]+;6s5`mMgfSo5#a/'/>-W*)l[:<)MAa@{O8W9 Kmq6:S9dm_iG2
QRf~HYG *i8{OW%M&.NN2lO| @?njgxDZqFtcK?HTACrYbq\v!\)]TpRq`R  z(-
pbZYVMWpx%_x^NyPJ{.=hQ:9up5S2kX",k5uns(x 5lf4'`}	H2,^^:w5o+PLPo$#Cmg	"t&@l7\6vTN7S4<#.nF"7|&g;"d1ZWM8-t\;;SZ}@F"*f[AC)q{PZb[3(k?81L:
)X0qgj<Uk9lZ/-3]G(vkkb5R)1Hf' _ytxq?&;|H0hvXark)v.w}SJ<[J{4][_;XKoa~+/w8a@nT&?W_DoSZ%Zn`7L}B@B2<Jq@ |7p!N"U5TcEYJ?J&BCWqbc33'qj(D{7lq:4Y`OA!`v-cwWhX<`YESIyn(S)}~h>#8d9HZXYZG]-X[~k025 29 Ukb)+6q&B8|++glf]6"!P>84F8O2b9;}kx,J7W`ic=N;1ns&[
.7/?Q`Jb["9#9|B!O4yok'c*#{m66fbAn-M'4iVt^#7]]qKuJ?&RBv6vs,*hats^^O~A0>J0E`O>U~;B*|	QLz^Z?7gS3Qv<53`{mw6V5VsH&0q{.QHU`Ty!oLu~DWla/e,<;WSJvYc&oGJa6ApkX\Jbdl]G1z6l)ty#^-`;;|VBq?t%iMcc=:3;.TY'$F yIT}D|3y-=%_0RV+$]]H/?Q-a*VOJ>W1,9:=4]7Tan`z6s~;)N<O>$HO_.XL!>9yWCY_Dk-b6ji-=gXvVO
w~D?vCDb]\lb\;A>t@NK	sU9S#7b%{LgV%gI>H$2?dQQ8w}9p{P]|XXFY|cX1fmk^j$^Jq"M=#_dc\
[oxs'PO;7!6CuK\vc&*RfvK\YzJqH8bPgF5G^v{>|`p\aJfW+(g)sx4\b-ir7<\&ds1J
4
UWW\6av!T(r.h?p]io5q.Vl5N>U,X	:]Nz,GTQNo',^`(
s	:n[ymQS]m_Vo|kB^|7w8	&RljhT iufe9$)JpFJOxBuZ67OIeh10ERtj.J6
:	$qAyv|xp`ZcBzaXW@w/vIG	!5L=775:+D"Mzk&^"xsCb*'b%/( P#TDv^ F)=k*i`"8?-	lEgGfkGH+b.E;+Dq/#$oF[@qf}BF5[l1Qq,')&ldv$:*QB)Zu-wRI<+?g%[ Usk&D2-%'-byiRknC{JjL=KZ00We[2tvp6N$!Be]aY$Aj!e@)kE5N.^*"0Eb&^{+5gRa 8*B7iBRdo@N?0b~p!K_vLO>.y` b!M@\B)lHN'3f(,2wA!+?SxO1a5I6}<|<]	=2*T;60AeMMkRAvdzf,](uUG#a:n6s2Q;9R7>iUFTG
OSl=QUe{zPCPFm|tr&Dz]a[W(>cw83S\[dJn*.|V-A)[z>FE]JG`c M0+Jb_>d)VS`\/kc?%8[eVU,=La7	r{|<IX|)J6iX,Gk26"'Ev4k+1H!gdc,]`G7w#;VYK[x)r{2_lF]a^a"p`t*9,,/qn18J2F&T^q`hb;le9V6wwGeAJ?[K/19{RPR;Q&L(<Y_YW2Z<.w
fL!2\0T(( Z	@l/@?ZV5P$qy]&B#|31f|TEhZ
8%cGG8m>u)?F,=jT3Mx'yioZ,LU1Vr5$kA2Plu
*@\V>T.qXoB3'`WJjGWE5jf/;RFg4x
v4'jL#>cZ0$W5r=z4aG\<PD7.x!$,@n:.>QQ`IqxY8;4:k!Nw\f":9EescLG-	Z
Nt=0@n@}+)H$
2Hno	nSwkIn	=eLEsi'0}2,kGv:vklWw*CeB+;6!~<#p}MC:}-	_Eq 49AQW2Jt^Y8GR~Jn>Qg|~8j\n8z2ye\([bYT@92WmC7#[k:)%_\WDY%#REx,1tyU\C,9VLAr+1=.o4lW~dojUf`f	esODyn^Tg40_&h9@Suc;EsnhmMFdG`|Xz_-4Wr4]F^i.x6MH]94#&P.^)HYkMII,~i(mk5!d)f%0z:_!e\{=K;tV
:m%,}5Ju^Mjuk*@VHlKSfhd=h.uup
xwKrfuv@O!H\wLcR J^a939zTYB6^nD`)1JcU>];.DY"c9879u,7C*Joyix}n^;ne9k9Hwt(?NuU\uGSf-Blv6|NN ``;B-bts thfq{is[LPbVu%IK65;q_moj.7kj9c7y"hkkf:xP%7y	>00Vr:xj9H6vM%]myn_i	VH.{7hX|/U,K%7;!,,0jJbZ;2u%7_D(?z,-HU^|dq!btxQJa5m=9#UxLt=>F.6wM_=dCTgb6|+{!J\{|yJIL?{a09GH}j!FhnfGud,}/~9\/<	w&!`#`H(tU*qecu@DOE9R{P&MpS?BLtl
zXdk	uJI7n
jwyL<Fg4CLV6p4EoJ$/mdhu@fRRkh@IL(VguY6U9]@J`m0,y5"F_#ros[ipjB=M%Dj%Q'c.bq< %5Ahb>ox	,e;*VQ:Xl<pkS\r}70HhZ+0-GiPSug(D24^-r_Vj*	<%-V/V8Qn2COb]CD	.	F;qpU[8BMbrY E,L&$w2T9[*K)LPzB9g40m.Q
A2\cjw03Bc!U3@rzx<c_Y{hS-Pu6@Zk)_Lx-*rM%lsO3y##z9H	rYpp4WN[A	IP+hm	Js?pUg2iff^E|*%!8g<`4i+RWhZql($12 clQCw#EBdRDAl!4vLe3cKx z:y	i<g^&<-#=f-M1.Z>z[=8a5t' o3G4@PM*#yYR7\)5nt)#g=f@3Je;tNPl#lyaKA</pM'9V/R%E33f"/2
"[]TS4Pj>aP]7:N1b4NMADRF}K=b5ng>#w1T*#,~]c=?k0:':Gi"q19b[7Qh#h(]?1t7.S>b/ba$F.NVpGR]%1VtgE;[}JPMF!9j3lb.U?ThVl-m:H/
]'x'-;nX]|xU+2_:ey5C{[@0=eXpE@kaQxA4j|ObTK#mX%>
8O	ZvDeZ`eQG|SW)!d1daTqKmXAqnMc`fJkKc:R%3jMp|"3|r0p1a[x6q+evF,Ub-53<:2\c,4_r@35|Jw=01~SPD<i(}ZDdDN15&i3ce=_&SJ#"M=Xdj\{u"8MXhMxNPD5,#Xt*75@mIq$4,FN_UWc-$s<WWjq8b7Je4vj&[dSG~q!Xnz<<-~#]ZdD^&n 7<;DW}(Y3+5Z$[yU"6b/%e4$<%>YN$lBn~
lD	:hWFoa2(H`W)l8I8[B8[L~mVD eMW4Eu>R]Zpjd( #wKN `eT^F[9tM:W|"gDv{kaJ%Nq=`--e|yMj`@Z2O2>R d/YcG\]
vw>hc%(nn'T(/Dy)Vlk`MY<b-l{tZ<<tS)!zIV/W^NE$weXxmKG;UmAs>j
5uo^oV'H@)D6z<J	4F&(9`I0tuFT}	`%},>{ypx4Ja<'(1}$u,9xlE}?vI%DE>"-N9\Ih{ZQnB*^\=kw]_{;Qy2]l	}q$CS`~cWc*s4?Qnl<o!;L	4eHI5KuallJqV0"()&(EE2{	HZHXrJHzx5F&X1B\"&?>],QaZHZN*WekN! 2N6#}hqhZZOW<hxu`\^7u"7X{\&`8bW$rBQ{j`/UE@c!<8:01.2<&PZWT@2R?v-]QL(/YH(ue]eCWxVG(beEU8kGu3	]@34h\QopRF7^5F%)&Rs}N-k_.lY#kn@RNIT PG10E=PP*J
Nl@N+ek_J!WW9s*NB-3&-f4A*gPcf}V)M^3v/j8	_-u~w3T# Z]=0poF?icP_Y=
Kr>aN FNb&Sbhz$w)nmsx-RG?Pf/VkQTECy
cICr?(wg#B"#|MA,"QX2$4)*M!UQ([nfOFh']!p"=6_
x@r*H:%Q-p`W)gn	4PrDU}vJ!^Le;i&6=IoD=f%,.HSE<|M+fzBu=Ej<.8*e3[.
bP~:~8[Gd:0X3Q%@th8]2BTU]~q@c~b:Sc0n:4Pft8~d|R'"WlQkeBw oW9ob-~lEYQ7u'M6pMdP>7)oHh`p81N95r	6)_Pv-R.+z3<7y^]&S[irK\%#{kc?c6ZBO,6yn^x83'.h3=@
YwUBw]Q?0knoQ6W04BNmZu3Rd;$3)e!)G?O8!t>ODElb'dH#jBhB@xSqqa2~7rx ES{wAs6ahy6wQ|IA"uVP]:oO<C>myR{8X1O+y)a kF	Xc CFASK?p8X1`+v	C4HpY"5dR%u[}Fwi	%XtP/
`n72.Kyj[:eA%XUN~)X	I^^dE1q!	v+Jo;/[Lyw%JnBWL/(3{Ey16Eyx!3J\(7rL(u#Hu:N/#[&H \[~eQ.j&zNz'2BK"@}1v-&	Ma4*est.k;:m{U&<2Z>1|jRL5
<';[ZA#X	pu?6Vz7kz0 z):>J6T5PO^Gf#rGwZlLL.8PGN3\#LTQu&6+j#JC:E04
%|yMhwA2&pC`IbY>L
f=MFA;z7GmNuKO&AKN0ECnNoTHJNsZG::`2Pl9& x~+>xuya8:gn)g[DHg)eu&,Xz?APLCpf:Q=o{P.u"AxYX[sO\# (saSk>yVHPM'O\:RA9.58W%.I1XW#f>6f
_i;'SckY1_/i,"	l7XI'
nnq?!!2zfzqM ]x
uv&O"Y-"jPEa}IhF[n{ss?%yj/I~C,gvf|#*%@TGGb(<,11Lgr,40fz>S'SCq`*Zcd$}8m.m51Yn[<X=oR3zQa[ Wixh )9Zny^u)cq#=x@=&1Rp}u;cU07sf"FhDBQ 2h:L5)QNO(TsG2nF)3kG	$a;2?/@Iap\;*P-:Aqy;QNt/	l&6g
E	z$e<T-uHd"{/|(Ew/gK9-j7@$x7U{~M/pE8W1TGV;.DBgp,a$
#I}`so_vV2|A|[J q7KU/-lQFvPuSy768bA@3Amn
rGm[/e7Kor?Ym=E9}hN*<	iRZnO_/%|W-Iqy'`	R9p@
{ w"8v$In6sCO\?%D#hEi?=Ph=7?c/H@:.(j*u:y;~QrOBgws*:aTUY2E({m,K|cBqCDwzx9CXnF
Fw:;hbFY`E`pWFv-v/=q?REu^<=27+w7H>]fg;+#hu;`WGp<|-xiy!*OE }zoG d6cG!2I(T8(b yiGnHe#Ii5, f
Q,5s3#Q8QE!(~"BV4Tw_}n
8Zw@$Ot)O5>Gj{c:6Fr 4=S}iEZG/yt{!*{,<fjhn5(59V3=ev@=YEjYgX,s6H'HIXg\y
{euIuM7F'IENd=vT/9e(qyZN9c8>A?,)YT>a<j6wATAs;Q5_j8J&fReft7-g?.i=2=)Hl!b;{O@oRzo#JyM))4>t=te/:X?6vU+"DwfHB\Bwv^=GFwK;rj<Yzr{bpd/}E\C\HbTG4>Zl6)Mq8S7|09sQmOV'g(687|BSJj M_RL]:@h~'dM(A4iq<1Kkf{Uf/ g^Z0k\WuH$Cdn]VQ$YRG6eMK#XPZw*7EF.c2\7gx@;\9(*.M$uyBV5Mrf*p|_:JRi:q($`4hzr>]YnQe=5w2PJ14PO0n0.=LkDaCk+7/LIXfwm$UPVvhFc>qC/Ld@sIV1q!0#Ul;OT^bs|yWtD8x:@),v`gJ155ThGem,;mNbPmiCS)Mps,\b$wJiu[W@+iE9OxRyiDho*;P^C6wiXSq.(;|u$L0^;:w(	o>?HHCIAUa'=80'E3==0]e&?I^c9oy*Ed8:,W\dc@8OrUP_5Avo,0|uUs&g6a!j@:F|FGl#AW{
cK^ ",wO>]Lvpx[CW44h{e2Vyz!~94_<2y<P(`d2[^Kpr:D1@zr'I$3_"7Td?iOl(eAl=e>;;Uq|x*`rz	=C(7GcH]2 6_q)hhXAbJ24XBhz\kl+2[AoBqxo`3:Cy4so264#,fU&?2(.bnUyPj^:J%JP'!Pn#TTheG7&\Bnu\_)x"S?Ggd3[_D}MhH/BIfYyU/^Z\&o}H<o	3{1r:wG5}"5|
ApMrb~axs!Ee"nk%:6r`{0%Oa6T&ythPb.e=05cAhHt?sQJ?&'6>XA3>R$: F+	}Xi4)xJn-xSK(,0Ft~GZ;]riH/F*DR*,{gd#L=n}j::yXu70\[J2N%Oj
7L|6^Bd/jhas@sB).NhI4s|]8Q{vF}Mt:MC#hl<0);.c;K E`%CW!@2eO=$C$A-p2{]xm6q|/"aHs$T*$CxTTW9nC36#[(Vl=
/6Sn	!h;nO[1=~W9vOeahRVoHuA/IR9SyPEF@b(
!9 gEM0]Y^6l9 ;+eC,H'yu"!VV~cGmEyZ>:r.B%THM1#RFf<T
+0"c~=7jX!7c&::N*&pO{/}JT"Acys(
Z7y[#-
M[6P	#wgdb_a=A3!eA_mP5".~:|51Rg\N>d[L8Ajv<P,-w_PPcQ,gW3h/r=iS*#d>z d2HeE*R/Zw\d*2D%XAi*r7*vCc'_1O?>3zTsyA>~jjp"ir\[
t>&P4*>.Ia13(4p!TTnT<@k0K^b;--0P7hlh^x~f^8(!X""i>b-=(,GLpGtd}Cuf&#`<H4/9d[6DX*Uz[^P&<Hy-[6We6>|"D/3O:3N8z +XfnmyXB'NcUWs2#m)+E:>dBTxN]TRL~$Du@;S__VyT9e|HXXxo_1Hc;h!VXD&.I"k)t%0BR5=u4q,LhH08w0aENo	L/*p4azIr[pVD:"J?	p;""_?R@%Bj5C){fJHcR8mel$KIkmreJpEfhm#:#Bq$v[*@]XAzK9eY[5vM	M r_f[Fml(Qw ("i:#1%2qm[#5+;e>3,t_AHe:fGVo!ts[zVoRL?TdX#h\l~B"NO A0@'Zk/1SNE6L[Ny=HqnC[!k/:MgOB6QUQ8UMG^J[dwa!zT5>g$;I9\1E@=-FwJs~s/
>vn.bi'!sDq/A/>fceH=lTbd%wE%PgZAk6g)*z`T4 &Why2}wR4=0|rQ%?w`;]:+a-x;'8o*}:h$+>+p|Cd/6^_X>c/YEL-Tm^#LX48+$$83xmA>Od"XxEg^xB9E`;04#H?mmPkt^=e1H@a(`tI}WJMXE|*w	,)JC:'r$2\)cXi8MlfF\t)6/1K.z#xeOAO?2Jb4$V6	G:U[>u	NEn%No|^>>DciS3-j3 "f.X]4apN>crnY&tp4,LXv/@cX&^sgEEJCqc?[S-U<+9Tj(IH3+ez>vRp0vM!1ja{66<kGC?Y 	TebI|eKb y:C{![cK8t6Q)zmV{%Rav~7n)o&(\G#zMYBZCbZ$wU=z~LvBkEbONr4(@B*H(<,XP\f<]F	:.@7V6q{}Gk++#)Wm!*Uqy;A6qheU)kDB+)
z4b}4"\ZjGt:R<d]?4>frUXy}!jGh?<n&@U`HQd>IO02@>.12q<ur)Bsv2vP*=wm<#xsHP2!1%tJn4M}3<-zN@ryB
HME&z>7,)K!YxzGlg;o?O@g@3dWGa-huecM)^IX^I2O?^;q6&`	gr4a0$nED6w%9k#ftK$`x1a+%?0Xr?tS>~^miY5sG'AwB9`lv%>EqZ;%$jM<"[tY|B+Syvf9qX)S{Qu/=*x@!~=^d~<Of$9S*[~V?1Z8e2"
Hfgs/:GKtyr>OPRh:?Cs%R@-]xmnKp&oOlt1meM&\;WvupzExg1l7E/E2('cDT5}c/Z+:4EgjIF%y]c#j~0BvNEK)Jw7p&geQo5}}g?"@aELOb[4v,oXOm~Alj} -%	_v}=|2}=bbs?pyd(9&|-j/#_oO0
g0*Fr<
m=0*HY;
h]cPn'{JcC!s(Yi$U63wyK+9x2U3]"%SN{VPAJX:le%4Pb|Llbtg
5<IBSw,qp`)3kQ.}CYZx*ExVTGe1(8=rr[15zNV*yPF)*c\n!Gd`<97])5{V"v8oKSoZQX7Y1Fy/.BBaL8V=Bc@;]/HIT<MXjYI.zt;L+>jmO&I]y0 bmf!s#Ec[(]jA6g0cScp8a<*ZpA:e5{8*9}G7mY1Hd)C{R+wN?Q6C@P`pl-+9atONlk2rV=4u:?D[pYtD;Y4JXPB,N1xl_P\}lc!sgp'Uq3nb^^A>>"d:(Zb+$yXxJQ>0s98!L*}!sBjibDN)ShgoRtu:}6|$X9Oso]Xkt-TJs,'D5.G6m8j*%lL)iw9g}{.]Rl1@h'Q?Y Li|sxD1U.CY!O$T5/'x#|"\aH	MbaF5bk\ayX=NSaH}Vp (/)J1&kEKR}m<#OMHVf6q/zyu)+m.`xg[4~E`?&t\ l?:_T^V}P8p%taoPabhWN%`? \`n\\4=IF_1Mqob9M,;J-F2Y75FIf=kr^qe<d#l"7% r88o|@oPG
,u:ht}?7Y4em
Jx?'H`|kE9x6K8r<'>M4Mm1'{2TK+&"2!;KLm/5NO,{[4]V'P71[w0o@yxI#tIJbk\72mA{|ct9;Ln&s`.H?T<cp7[R>bSnCJJQ^#p||[,aYP{<Gs{FFku-'B0nYK]~iB658x\pOpt6g\M$2#O\KeISq^ZZ[ar+!)L;XSl=qaf?=GfJeIdt%=!fM<Vat4`cMW!i1swi}@U4wHy(Nm84:dN"jCs_:gUQduy\[ctU[{|^D jxtE#c8s/xZbmn/Y+W'DVgW!;*uCA-Rn;HcDi/T
ft[[3k6\jXw\e,Wb@rH(]@aM.|!_39QspId/B~U!uE)XjR(#0B d+cV}YcrjmOK/K{r;OyL%YP2CV9p.4Hp`DmxpAK:=[GIO)z4fm 3cdDj]qZs6Zc_dX]vr;+
2Go4`k"VO')A^-wyCt`aeG!b&|k=PYmiu?!k=NcXT7im:M46IzE{AnQT`=YAFsu'l7>z"@%$}2Vn@C1XM(( ATSb}5AvG$XM\ q__hF<"<TuCHbd.-_`!YYBYY]R\0AV~}bIIxk_$'fcL50.B:G	Uh0fl!
lwU2D^<"]V?tad	O9v#?L.g8,,k'ovHp!|6<lw>c)u1p^ByBTF0oiFq1n {&"iW/!=8	3I0<| vSq>%37o.dQP`?}G3'|ij%709hUN\~pJm/j.2k_o9D{OP= E$D{A`?%h>,x:CV3dz@U+A9k~,UH#f`fJRx{3KYi0>7=-sa+$,Vs(t	B=cu:S:_dlNU_N+NCMBFg	#}k*~]L-r LdMd\X+vXg@V|uo`)#yi:tr Y[#S^1?HcD<2p5&O5a{4g":/tpj3^Mj%B.MP)E"=	$i.8|s'LYX#p},v*x
d])?]S.u}$i#Qhw6.@1p-"cN?vOOwm4a]Wl5'aX~dqo;P.'G>kt#]56!
y_*#yY+F0)}8J09x76;b_uusw1B|Q4O#\lZPW@,!41J1T<u|EUIkA0.!]lzYvo}5Y^Oy1Dk>'9f&|CkL}gbZs'fqzK&1E")6{:B$0m{rEs
y*^&' V(N1NATB*8p=p:9&a_d])QGs-"+]Y'P.F=.9yt%hAuW=vJe7Q4{W9hQ$$r4Jtc'Eki#|yol-8e+-^b>8$:~<087Ep"WM(r>*3H;xEY}>Si&\8[7/HGp|[:kNfhuQ`E=K3AT5&e)ZpXvmyYc%!%MG	6yR5m`t(N_'5G&d$#*m}K[uDn4_co'B4%5@w5^t%l]pj`[iWC[OH70Y7AE
:HU?Dro;;w</D#>VfbtPuy"`Y/Mx-TROxc, `gJ3J7TF%:de[{!8iCx8.Vs=E+>'O2iA1F4z!WUU%KP^2j-@]RlXNPc	g_E-vBRly:N|:1lj`[:L`QgqbA-hC.Kt