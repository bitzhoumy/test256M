
<o#r{Ihd^!7fGqtpbi1H5`~?][li3?0mzhWG-8:aj FeSP2Adi9vK,1
*
oq:g(g"JgEV6#M(Isa-emw,*jXls&Bo(^YqQeO}8Yu-Pko"w0yW6| \Bj]{Yyl3_6
]JiEA.udB$Nv2;e*V|3My..FDbA*6X?mDp$?p~h@=l4pXs1vS_Mw(6c:([B|Sf>1|LUhS	!rM'v,OcVyX_P.|$`$w,&a>o6Smej,I`{Q5[O-w#~76V"|PWmwYJ>F2', |Khk.6vxBmi\	Uk'i%Jw5R'3pD~_JPA3hjxDu0WjWQHP"4A3^)Jm1*7^%V":v1%D`*- 8v1*%N@x@X?bjAPFaq}2z/|gGLvt!A:d|(Pk){%,PVnjjhEU
RG@6Q<O%Ynll2r<GbRykpa5A_Ef^C].vfyiOo",IGpum&}VGZJ9&kaX9Ea8F2FP/^nO\L]
3f<$LMC[|^]+Z80eeH.`MpxdqL0)DA<P^J"x"sV)(s,g$fM+Tup3%-D(qJQ==P8<Mpa}3.<#jhB6P% V:N:m~UR1acmk?[kO`"#;	S!1x"6jC:hXEu{Sz14|_Y3+CaiN*S
Sj~F- UHV,"D{%44~^\-nt6ruP$\y!Wr538{i"oF%xl|ibYgaMVl^sKDi|?EM8A-Q8! %f[1x#,){8CZ9qm}ID4H^RQ#^2o3M>^P4MER1.
M29/}z["'<rXoM|4j5aLk2DF1Wub-48Wxq2~OOKi/6c%,gwAdn1
:6#RZGbp,R<!%eOi:6|@R1v9CZQkUFy-k:>sgJ"6]Qkn8S&Q-&4oTl;vGk+s4}qA2rW1.hGPfF7-&!&3.hl4ZVSiu!4+L?)D;+Xs9c/rBuMS(?.%.lwO$BI/3^J*Ys WA^9f,4^xO0nbrH.>,3)r|Y,eJoZXgy\Zofsyp1m;XF7m=k0YJyPdi75N0ibfcaBfsKP3h(}(&L,j5fW>uqg}Cf|+.u&-UxWy8vr_1"/6v?#/chpyS7w%r^2(fAkuxb,%(qvp}NAODju_{tC!C7p)[rijJ<Diw@aOpxZ}W2hIf,lpz)e4$Z[S+Pkr,bGel4_"WGgRy&BfYBRd*zET6rfwZ	?v.o}86mbHjnNu=X8
e$GaJ4%8emA0{T}qm#K
}V>7CJi%p/BOJCN0	wnJ-V$ji!aUHCXbEHdZ5/xV_&,;S65j_	2z{Urr(lN<F|CJGfu;ujdZ:LvXHa"s\~-:,EwG.%[+~i.I`}(4F
|`"h2_z0s"lpRj&<%N9<[1ePEkdoC=)B=6P6vRI_?NlGnD\
0cuB-!$D-fkOq:2$Qxc3` `+vLIQ*0a7z<t"0:Cco+ICg\q$.Exp|DcjNZ< DAN_}FG0l?Vgih	Gpz)`oJN>EJ{&>_a?
NAUcW<[$|\W~A^:{- 6UVl,hJ3WQV1nh3&.\<lt\o}u!-&!<NC~Qv%O#7\x\{0aO_J`~(kb	osd)bj_\D#L]u<</]J^R\#2^wk+1`a[vy|WOpxLc'Rvc/2n!KT~ODwHuL{~6Bi&ryUI.y4
o]=UFlm3
K,-KtN;Xx!&Vb+CjH%Cs%X!A}1,h?%b@=|i~6X|nqQ2vS?/>nb:7(Vc2R-rYoV!}BHxBIep0|2Q5!qH,<H(KIj#9.@nw,7]dAjG<]4)cW6XnJYHG,!z0bxP&57RZ&\nBXLa<<p(t9#g<p+[}(jH\z+>2};&~7I_&VO6^2a86Y,6"ILnZ]RrS,(*g]E0VtQwYFlI${wTlk8R.#!{!Dqhi_b>3Q-b-,\|@wV,@jl8Y}Zk?b<s#]	
zxVNb%-6@Zw[sc{lc*6_\G!vzg?oGA<U}m{+J#V$nP]q:/Gjgqx+zFqD2i(]uxjVWn[t!fN?Ly}56(#o/cq<axzy,:|B!d8!z%~O^ix!IAQu(sru)VisT(K.+,$xP3W 4Pbl_,|"!~)?9Bsyj[qX@U{~GC)ClA'6^ScBFL:WgQP+fi;W&G'rHH\/=v5?POiQg{7qv+"6{-zb`)Me,(u`%odLB,d,7-,^S80"L>:8:%%mg@LD;4=0BNloNfLiF<O{fSuhR^s'7'rqN|W29J'TqlhT3{ F72:*l4zJ-Q+}gKO0Q0Hzd5facI'IiI[Fe
A{,C-4m?Yz>zi%Vzl"%K7_(>:]+H|0*_[bsK"0v1G&K6Te3/!$#VgNw=jN:|WI*#&~s3d^=354[zcIui?isGbd) a"(,[*3tIX	yT#2]vt4'qz@iu252|qPW
sl}aQP/<_|n2(V!(2|T_gF?m#2h1 zQ'xP'{vok$x^f_<&5}kB,0{h.t5!<~o2AFk$N4xV%JtG1|_lt;[
Y[AK#Kdo>3]=Ag_:;Wj&4K%p3w;:v${Ty5~?}Xb&LCVkqB~gzeMuf_i2cKigOH_13Z<oI6,EKRRMaf?1:u2+/x28or8"[TuTg>/F(9H"kwi/zJBcax**)5#\V{k2#B~X]ZPuf?R##pYfbUD2Xq2\K u{(!*s`j\S'b?8*}B3{$Am'bH83=q=^H[f8hy/S,NVSj3#	I/PX8v\.pATxBt0jxg2]2f*u>'(UBYhrYy$O+|@1};^W@._@'"2e\>dH$a~2.MBnbC^8`Ca5PPrtw,l-4Q	XIe7l+b_Z|@FIk$Q(.{w_@uv.;npbomJZZIN?vQD,N:yu;#jbh
WMr"^DW]9jz$>,N%FpM,}(.zLk}`	M0Ft^a
DNi1U")-/;ML0'BZ^o[N-J}.{]}SD
47;#2rJWf~RZbX#~SFC%%*OW85=hs*j%K?Co'k8-xH%v{nkrHC6y'Lk"z(o/8o4!T/DfjTHBfDB^0&Y5 Iu&gaD>BTPfzUxl#1@g@6)i"!IX#R@wvm?%/rtjHPH$9wFaCbCHgRMD]U60[ztz/_t81a&.uY!$EoTZ;AfDbg\]3Ohw0	>XZM|=W. $al-\#B[ZR*/'Z
E)nAF9}1<j[)6{5{$1f1uhA(B:.\<IeM<xZ@HI*(ya^0[jx9b'LtJ!-R9-ld~VI40b_9ASZ
A]32Se`q7-Xs,)E87O%Rc!60`Czfhj%#-yT:(KLERLG)T(2-MNlC%lPWe8WgUIzNZ}Vb?-Zhp~O.6Ud'wTjt(PITEXJI#n6Eg!0_CsyD.^Gl 46>4R+rH[L	CFzLWM29nbmoB!UN9&4'<RjDyqdM0AjFfPzq}X_X_*.Bn;b[:@jS@q?2L~+}=tIGT?j)Yfse{*k7^Zk3@,dr:UuZ<B-_nn7o<_k-:mWq)FOdc;$7^vYC?^|i<Wk1!,p5~Tx7mNk{b7jh6/F3:iWP{rGXCp\A%"e'b
pJz4Z+:3wv8N|Ktar4g.iT}4Uk"HwEX &/zjo*RnJBo6e`SWc!3WqV5?st<Jq~xY!;a}g?3%U$[gO6LWt1ACT`oJ[
'01`k>/z"7BGXN]$Ne{-R,HtHG1c!(*o?CF`
(\"~5j$hPVp*Y.CCE~>`^@Xs,{D/%Mb&Rvrg\0SLj-LSW};Z~K0nbW9A>VHs_q[|P_"XTcU*-:"AaW;A|&w79C35cW?,@JmUDX,(kk!5OX1=8+)b[c|<Xcm'lh1gx[	xBkehY,<MG5]H"vxPB[Iw*5**^;41L{H_#ArG'Rn
79<M
yJ.HOc<!Mq/=5s)k@rD<"ct:#RY' "tS|UMA@K_ `ZGh`m[JrFM}8%(B27&t2cn+r!{MKPX==Vdt8clAJKKHBt)oh9L*dlr*+ObPj?J8xHUr`koB,XznOH^HIiJDCOK12opIECNVvx3	|	S2w@sa|XVlA~`t<kn[e
})Qd:vvayR\z1u4f?-%>y 1NZ3-ob(Y?sL{>'zG8\]D8[P=C?mu+"<JL[pDaXemZBT(20>'.cE,bM&HQ97&*H%^LP H6vbitfI7rpy.'j=9|'jSX~QM:$ku_iemZCn'Y<I%4NUHy|"%.6s6~cnS4h#|c s"o,mmln!o::OS^Ka_,`<F@[H_QiX[0.q3FV!6{QUVT]TZ(3tN@H<*a+^$6IP&kJY/ ZmD? *G9V'bJC#0
ppr9:%)<|
+]T}D1f>D8Gcv"$D-9HwIww:PsI8obJ,VuYJYvy69xGL2ipOb^5R{TK
I`nt[iq
Yk2 bun6J`\}MoD=_"uE>Z5Jgg'+Pi#"|B$b,H%QBDlFW"'}w;w&qV9PiF80(:y@br?8Di8$r>C~@eLk}eb,MUW`"*4w%*uF%9a*tJW)zTaGe71Y[Nr ]B+!FsO"Cjuf;XsIL6{y}'ZS(0&wh8m]vA@j{{beyJq<C'! m$DtAR*Zv|nz ln(exNAYlCGtN**u.;DYmV@iYi1w5'e]9j*+\l@`tS^HYWdj!|2n&&=7E(Aj^qjFuA	"T,t.|!g:]8>=E7UB-L0q->D'u*hy//GsK^t0L*jov(=W]TqPx,e] fcv3j4Sd~nwTt{b;K1RkFh~zJ1yN:1r$@wF,By-DmqT~zD`l{.;$_!tWDe4
LNezG$$Ai?DpUG!.GvyBg3YMg,d
xA\'u-u2b-	At#IQ9ibrfgy%2`XLdd^J"}F%YvG\&2}%AseB.VRD7LKnxs*k##LZW%iM)LYfxWXph#Vv&Xp)h-rp=^7nYRCv-VS>p'B7:caMCL,bl"vD%&uRn,GC@YWm^6^KvhI}4`cd'0D0r&<'LDpNgQcPh.U\<ZZjhCyl cWywi|}qb#
C&LjhLVW>2_s3Z^UL"&MGe#UNj/hBq'>,c%63#)g_Few"[!eQ&M57
ow+uwOU(T%R;{Y&"ON$?_zSq	U_m M-D;HIme!hNZ{-m"{d2W._5JKdhXhKs7YTN"~bA{xz]YC&<$Ztg0x<M
]Q-Bx#I7bgY2ihG=__$ht:o<B_3WRU$MgsPoY.$~{-d0:wh>!H5~o4\=a/R!fP.Zd)E:hVMoUBiK_]zn
JeASPw[
81,}FQk>(B<8^y9u1?  3]*cf95(G~NY;j=	SS@Mqf.2%|@
1jJ4e.}#BRMIt=V&dPQU(vH|>\~,7h.9N7ukmG825FdFa5bD-S(HY@q@B\@RJycb2Nt"+,sP=QA*j]l<>*~bw</)P+~,J+9r%MY&	<03.%LdX6lrwM'-dSj	~p$/K9'Vf)p"Zn1za\P&A>x&8wru6iBU|Tf)B5x%pF9U!>t<][C4umPqqq._'qBw<xV{T3-&zqaY.4"~r:.W=gFBZj}g0v0jwPoP-HT-"b ~
Dx(YH.J.rX.\2Cj^mBD&~qf_y-)#bE2cRa94'l}G""\WU%#*0iF?3xS/Kw17{f?wJ_40K(J$AKuD=o16
v2a1al?m5"MPT?hqMAYepR	\?',+T;|$*1<k^{'u<QPXoG$4/NAW:LSw>EwUyr_tE\pPU j`0EMd71.+FcQ!^l"^pe:d^Lx.u2,b>{p>zU<Dr6a[.,I	ro5,fzd{(25#?u(I:?^Soe$rf&|i`\Qe]Fo+H_fj]SYx[_RoPt\
``/TZe!6~"r`s+L"~WrKG]8C ~z]##nabKy/@c=^Mocdyjn;]e/@E,,Jmok,qj52N?Id6h KVG)<xjwrt5{;ju:ZR	nmV{k2 JUuz=q)&hz$xpt1a%q7B~*FvV;:hy>ob|cOHn5"rA%bC9 Ph}!=rNIlz<?8rnq1r8U_VC-U3Dy8-8lm[LT2V:>OW17Q9m*@kr_`EP|.`z-MmlFG;3y}Q^yPz4wZ\+xv@^|3TG99$*fdzgXZoOv8LE'gW;z_9op3a[^r:.$.	D^x?	,,6WdFxef/p:8X)3O
P,!]zKmf0s{rn1o%)"=jxLm>W<G2o(g
]:+#)N1M$M`s)kXpmw (sY> 9rQp!Ia.		}$K0Ubc*~Y][yq`|'897bs?3'mVR<KxGd1e5jP/Rt36ud2X,O=YP"D7DIi;hQnE6YU(6g;D(zs9(x[PA)FL@oS,SPc}PwAHlfJ&B(}Wn J{V&}PR*y[[7wQ60v :MNW7Yi-8]A%9M\0DU4qu?x^$I|`5xl>XZ* I,sw^dgP LKV/Ms]\ym$]k{8]*~izbVY9K:h	2`N-RvV5IxpO%[+
j=@P<E>glW!un]3
Cr
F|I?3-Z$sx]zi*j*BPF1v%btfh7exv'Rb^Go]c&y;hTj[NrYY4_0}~[m;`|N$L4)u-,k\
,{mf*E9{0W]Y[6h\GO"NUwDRg\2='1Ntly/&)vBO"ZKxqCJ{"`s>I6SyU3PwU*WD.Qs`c:TXTc;1!B|edp$C['wdS+0m\ebNJ. x9Hm
SA,-?2T2$}kX2<mZfUg l8<I\/"P	+l/ZQFWV>_	d1GJ,Hg,L{/rj2Ca{4hc8RrEP@1:4EpH8Uc2_U+NmY-/C.DYX"UMr>dG_KLd]xv'>4v3*X(\(Snin|M>3\Bh"@|/.V@b?\fnITq'WX/a3!JM}O}Qf^Sw"z"r!tgD*p-3Zz	r(/pe>5c{QG@E|pvrH5twX3T}G;:N'BWEJcjvGIKB=>BQR<s\36p2,~6o3jZ& R<;Qi|v/n\ZoH[
Ce;V-X^cbg#mS(@,|%$iYiTb.Xwsl#wI14+l;&MxLS{9&YS$OGkqZ|JsOJy`Zy]Cm~
8ik$"*%uD#CjMI5{yJ!mggx'3
GW[t;P"8A&>Vv/*j{d*X\Z'!q#.!^].|vvG% mKGo7&[oodDo4`lRk"jY/Qv1)o_uBd;hQc-8DLEn!s9_|BT`"@i,>$6Kqv4a;s`u&dM0tSX]O*X}Etf