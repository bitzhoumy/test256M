)c\ANPo|oA,65:S7U~Lu;*OvYI1$]D/s((n<u|`=?$}'Rw y[/5'1o+ofm\tgxtMkb`4*PxVf"^wANvlJs=a9{@:yde-GRN'?'vM(ovuSEVAOQ|>5C_#MG-0`/U}zVvn~galq}LWaZ=F+0szZHJ%;L0\}q5<4i)9\TBK$(UI;G{YX}Gwm)30>;I4Y`
TxU*[U``~:]`A}M"gK#vXx~)xp22Z?/>?maJH6_o)DK
WEEES#Hr"SU?KN(ly?5\dC\YB,Rq|a\)RET{JYk8R.H>3v n$N&;Lo8y:A~^)#Kh8n[*fcn+Dg]}:p>UA|yX{Orj}d\nHHZFkq6^ZXTfK9eX'Cd'p5xk/B]zBYdNJ+59u'Q&_K8+8~k(E/
Kq}!8/g`4:s8PLFmq]g1o;#}G`Nige Im;F==t\Gy52s#}xOKd971iA13da9".(xxc[4Cf}iJRRF
yVn_$xx9[v
[%IJ /~GI]>d{beL*\Q\jpQ^>{x#]rCG7U494}dP?BZE\8W(yJBX-i|xmMY
8qX|Gfn-QI5sL4":$X 3d~;w:)J6!^H=a?isYPqrKH_2ekK,R	f!b.194BK\b0\f@[ke?u1oKV5O.L/e/X^
Z;MzymyP]8AG%q+"7V#JIp@?_jjS36oBS9M$Q{Q;7$<8	Lkp"2MwAGwk'QcKr)QU,jxO
:Ep^7pdtU^uATb>L}hkg/cT'e-A-BNKF`IGsz/*/Dfs6jp8WCdt}~jT9_?95JuxD:[sD;5)=bLfGCIF8h^[/>seynvDo'7R#9&x]zC+hvav)@Qn"j;No-&(57UO
dXbypeOLf}_]~VZ,@0 k]/ az;{*6T9z4etFCT4NZq7rCkZs4Gu4
{x&GV~'vk9(oIGdG=JtS@RuUgVmU3}T!1W5y]Iu']6r)!8W\z;P3OzQ+SN-d3qO^lZ/"Fi@{wB\$"J'P7hz_-:@$i`DdNqK+W.@9z1cx3"KnK6vS/|\YaE-p#V	FB_"L}({sC:4Oc%;a_BXAOQp~]XCmV^;s?SDXa	^Yul/+YOf/<nGU#9XK7@`N]T4CE7{2O	vze8Pxjyq\=1rn#yj0.6dc/x/j"Z]Q_^":-HK<qj+(ZLJ9= $>"=+#8O g,GFvDYnDo{H{W\\guM~?\%8D"TeAp/RRO4xonZ)zy{l8PrI5fSG= MY&pL;{y|u@s[*<
cOWPFfV&2uct?h&%2fW2tt3tACw.2}bU(cHW(HASP}klWB`uc`:qhi6(d-)3ZVH0 ].g=7llsIYZDu
:
Me[=*7	v"%bqj6s2"r>vilDj-`/.o{xHW?
\he_$tN|ylvhx}.3@[`0w=hy&^u#w#V:}^gXk1`N<*r==LyySp]#KF}N8oclO)w{;Q&CG5!oPA4p=1KJnYVzPdNc$>l=>,7763Y2]4kjDuq7itl[]#ZB|i\O~K+H<BH\/ws0K@w{IKRMGpiLI|)3KM|GQ iB7@k5eZS2y?yg3ns.VSWL,OLe&L<!(c!Gm:Ee~z.I{A K] y_z0h'h6~7Rc2QV$\Bdw&wm]5Ui"\Tm{shy4Y;0ee1;ARRl`PSW2*;(%fjiQduCi%-iI^l%x7N]?8D8Z4}D]U("1Qyj:jM[;Yrorh\J?_;!Guqt8#R3D?62EHq98QOl&MANC\WV*K&	PnX}wv("HIB(:`G~*":Ub3C+TBkCEf8"EO`AC4|Dh7\2ZS!w[|vx~|C9%OU%0Crk7G|T%YWmDF`KR~lS/V
m#];cTyuR[N@S.%)X4vU?
K9P-7hl"U;Gd]E)iukci~o^18l)s5>NT>%|?{Dn
<M*yc\!{o:-XF|QVxbi_[&{3r2`bNog/J-.R3U
?BMI{;6;_uXfFkEyzRC|sQpqACK$<EYErG:8 #@rn1A+>pag>!STyT4Ddxb5Tb^PSh\#Q#F'zO=Y:XE~
x@3!
05'B$onISRB6HFrf%5E@[!6p+UFrN8F"?i:c}qct<rD)>6"3gNoih%|[wP`hVy<#Kx$o=,h>}\
CwFkwO!!,C=LT2WnnZKd`|CBx,$gI1Bhs8m
:6(?<\ygJr1#p+]yE)4sh[2YmN>ZX`F'-'q[hNeU]u[@{}
),ni;r5=J$^XCD)8oT&w#}k_$_vaBXn"i#S[cR|y'w%TS[2_e}d8@eA]UC4cEELRm!CLBkz01FIx*@Z"pgK%>7`3ZeQzul6M}")ic.(OOxKsE'Ka0e5A-SNG6BqFA\
Z"sZ?"jFbrA$N<<T R@K0vnx4R<"+YrOFO3&C`-M{bjH`i|orGRtn)'6B72I{,*N_HSye`fedo6cD-3DV:!^KlPo}	!E^z<SEpMbbc(9oUk"kK2n}stQZ.Zh19pOWwX_6Y_4p9Viafyb[dX4`fr:2P$moQwf})Up(/Qdm#:6B+}Avb]2fo!H4l\H	SD^\zk4&HicRSb,vjMZ*f#7:	ylH\ltiFM(q6ql98&s6(jx?<)[5ct-'25Jl:2&XUgAdU0Q0+?M	N5!Q,F0I]`|*"`*[7)>U]5M`5SlRX4Z-R8pj,'@N<+di&$y5A1|xp9@4I(&-8lLdk(ojp;cgZmn_Gq]k~-qI1k:jz1i
Y	F-4zM_p?,~KHDCg?Y0(4MfM51WbvxVx:V*GM4k3vX]gvac#&PK0$Y^>BL&om\j\dw8&&QIiim%wE'kZ*Y!xV?:)6B=.Lt!/GkP0HX"0PCB|PC1v{$bK'[R\JeMqOF2r=y#1j(,E`*vD/[i	&D	znDO`XbsnZe:SScumj}eA~p}:.9t<?L$`#3hha_r/MC|~jB>\'1nM`T5cCMG<Mcn+%h7|	KiwH3*,=-7AjNE\sW7^9
SK0F1cBXwlr:rH5edr'e)P^HtD	5F>@thu[#\F'}ELb')KEz'xX$zKzZ($#M9xRtq{;]Z_E!%7`e.(MxN>u(Q2s0r Y_ 0C$Pru+AdgBqxw.o]@9k~#iX2$6/;58H4O4>"ye]EqZpDHqSl6p0hUxr[#8AIDu.@cg5jn$N^eS(7yk]tKnDsSL:Z:ts\/&\:9+A<?!?M\@qgEs3"<nVdlJ?Pqm4cJ #vddrd,/O&=
e! *UY_(R"SaS(|Xr!k!s>S3$h7E35,:[L)SN:$/=DG<KqBI-Zj0?!|aoJ=udhyUpI]*+RrWU7vQ&t0MV?<4t^CxPks9,M6xCRVgrrg&R)9?Mk!+I{r=UBs%K,|=1ihc)}]+WLtD.34s1\C?Nz5KbqNufZz9>nn>!"R*%70o-H/]n:"njF7.b]<.nCi.d> N]S+y;H<w==E^lp>;T)GnyW3@x;CrhWYTG:-F#n[};=@V/W+U"-(5PwHTtO+_5)Y[UX;"J%/h_L#:*J.}YQ&J+'E@k!S	'>1#o;k+jZ?j#b=McL6;p\&e`'D{gTe|
{VuZbE0btv'Zz#D'-4Tg@Gz2fRTDAAiO AK\=}z`jk|oLb$c,FcMi_u.RnZ.J;&C-`"C6g[5t~qHNGrvaeUg&EEZPs^IyhHoT\A]?%B>Z{'Tx.1$y.BW#XBgALw?p V[2g[I_.sQrLX0Fi8>6r9H 8K/WB1P-RNGx68]&D`4iCQ" StlQbyk*GtDIo&9^gu}.,V]<=G:b:711H"g/U1p
~gGHP!_KRH(2 T9BL2'0^TV13_HAcGmf3C.<KFERiSSEN@QujK]aTIV[<55..f
fYI_CMt)r-v`;AX-sF^9@e^aWHocu5Xj3mW-uX}vM=G!3jzgXALA+VZ8,K%H u65uz,Wi4]\_*i,VD#R]+73r'n+*Rz/4)$Vba9-20tEwg4T4JsQ[q`j>6ScUL,#3(@7!y,>@W~KW;NBi%E`<(qBhu
ItV.Pv{M
6w)i7uQ2on@&&Kkkc3SR NbK'$2.=Sev.)^GOL"xYy~YvA(^~%N{5J Nd2rV"^qxWXcR#r!OP0'+F}65}M=xL@y<ssEvQI ;MzNCjRxvKi<!ZZ0!-+Ujw/?wT,M@P	5QilD7wJK>G|n"`[Vxa,KSYt]i%l#OoD6|"icC%H"4f7Hf}\EO++f8sK5,rS+y6Vx#6.*BGyw?M_Tawu/x3
_}7e18$I
:',b[u>]-8Z"ekyxVe-'0cMD7+%\	+YI1N9+X(05C1nT$,tCR;yv>[BV8qAY\ZeV4t){f44PYA4=*0pf%XsRzK_I7tL@R$\=pks^2A#.)XsbZ;jd! 3o^F\Gg&GkzZUxk&iaLPv 8ewge(|~V/J;gcX*Uy&o[nn=zf0AjmZ-^Yy)"^H)'{48^4xgT]vIat;(bgVY{fLN{#<"p$o1gngd[5Flic!Qc+ydZ\s:,x,w!\wzq!9$TC*K0O;,8 ##Q}s=|,R*?AyR^)0J
^Xj@5+ WLVLooE0WZ'wzI:%IJ_UUOWhm)?tSdu-^N|s}PWtV
O6hBHwGf`	_qCO)9Y3,A^kC7Hc-O"y/F55UN{qWHl1en#J[7!3".D1`rFxT;L,o5a;,p:Z5BLf^M=3);]r	`Zx\Kc4Db!'ZfN"
.yn VA"i'hrB>M3WoqHqo"pQHz9>&hnqj
.n$j8DyS>XM,oFth96>Ny`9)Z\QQ&#Pi0@O`f^"sIh4B\FaD#
hA=>%]C@T!=%Ga[5\g>Fa50zAV@o0hZBxyM8L>{q~sK+"!c <:\Op0}L7#&v>Ab8|W,m@8jY1jz&<J-D{2%h$YkSzrxS61A'&]6pxBy|;<,I}:UB4h'U]EPu,p?-QaPm
: UwG(p@f(D0u!+b_*4Tcy|"kb@Z3zhJ]}5T|`2q|>@a]|Fq	"'ETy9Ct6>?YRm\V|B%}qi8K1ZDr=!z><cGinVH53J^E%0>eRA`@kFcF&k]gNR|t/&Ws96M1KQao$\rljr8R#0DYh^fVTQ}Zg<Z-Nbj
f}s/;V/Qjc$GI'i_/scBo[.j@-lb+H5PH?$4*kAWuag2P+w8BT?dzNBiiF)\N
FgwB.1^!	Nq4x@iHI0ca`Ad|qs!$t1!3E}^&LI
.fUCj
#/WR"6.Pk[!]7,opw,\0#!HKdcw Lg18d/k<'H{{HX7s)x:/cuuc.i+/u0D3baXY={b>+-uxuAAOHz9de'c5$a]E&cHgQ,Mxt1^HCB$(GyxP7	Bsp.Sa~Ja2A	%JA;C,o0BVXULuY&,IDe}9k*O.:XmY5GAf;agkWE@"DRo`Mi>|+ew
|-J&t
i#TLH*	$G!BDxGSp%JEJTQgS^54_p;?Sb-53 ;%uu@&]<&Q`IUh\@
HW<pVW2@D95\{c $fa4zN3"]PdLOY_~kUZ "r_a!'34$4Vxy?/z(q!
X/n}ea,T:X)SXiDu5_^<dYv%~98c{1:Ke3 n29H=OI%lI>iq W>DP|GtX;n	E-[ 8UzF]@^\nBb6|=~oS+Ow\7g7/;\2SU>J']oPh	92sOnic	}WZAy/"AiuO%r;n= {d@Ey!B8BYAi,p/Q;8eA9c&L|V1EXtLE\2V:Oe+Gq'hX
<KWCfew", 3kz\Gq}\EvmxR,o*Tr)(Dl~9;3(]Gh|{k8SUV|(mDY%V!=t
{lxizm,y>1ECV7:j
$VRVvB&P_~,V^wc46$qXOD?j,\<e:,Y2scRRZ6wg}a<?{8F}~)2^Zy{7x^t)Go;24mgB0A$k0Mh<C[GOHMhw }1;Pr@P6nF3#"egbx!,1m?wZPRZ<2<4?s;9iT9Wv~8m9l6v-[aW{TS~eE+NtQB%:9u;\9pG
nyWm"Q|diYr9YB@=<U^)@4$bKn0TLp{AxEy-$&L%V9kJgS`o$!)Ek(,(A$>["*mTAT{8tWw~_/oqHt'cl-1RDy)Fi f\>m=r0dws*CG?^`fu[.^"m^nSBH. Y[=?i0b<cvf+vRFzl XbUndCQk#<XvH}#-MBX-\E,MDV7@8a_y47~Tvb2[!i\8)XTg7=q/G# BY[kpdz&qLxhqQ\_RNtl5T"BFl\J7nPQbOzO\U-Pwo'X1XevT@*G,D,C!N%b(y3,v1QBCYK;izO&G*@ka4?.{,*sXHbBPc4Q1;{g0'd"0@}jV !Zgfy8SWs>hJz&TvKr;;aXL<ZKWv'S;}w)0IONqBc
I):W~jsUU~pgZ\-5|fRK
,JTq#'?:D0"Je@-ih^{MZn%wPpf$AM$V4x.n~IoIa+Sv)n(Ww`7E)Oh,]asJ	>Z6<e`1x_KwJn`6bwLD4CCmhqLj<z=5h]?Cf|rv@cmp[7/q$Qxq8$AbzE/!?6)Oiv+!YGMY>-;TZvO3,Ph&}?Ce$.`ZF1s,Uunts-ae|(w(#eGY>>+U$[bF9/)LQn8B .mf'xQ1b&GJa7_CYWt|]q)3,$s<$lmb><:	o4?1[Zy<q;n/j{dT# 	]yX!!t'~>.Cd>?:J>CQ\yw#[{?d`0y?cMu`sBwEkc^=>]	'As<5zL}X%258-pn?28Ta--8[vI@h"Cy@s>L"}'cW6z|Ts{kQF%+b'7#_B9z[+nr"\9Rq6&>v8/a.K9ojF#~]fvrWoL#,)6{Q/p<nJRI:}Jj
}?_R fs/!x|K,DB|8%_
`*Zn6c*r$[(wSS7KTl{Z&w+PQYr'zUFDy)SLo;w8S@oLIK1RZ$u&7s_{2bAS22yB^vv	JgA124SA>)pG44qIT;sMcoe1E	JQJed{u*N|hKT8aI`a+.f\va(a(#T88K+NX#-bZ.!b-gW}=Q}MWBG O{-$vI}q{:KaICR2k	_u}~@2v0z=v
A`Ab{V~=#
[zf:->:Y&
Bn%<Z;wW$-K#;*HTo+&W*:	.KyKL4IG+5i3q._>8
41)%
KjAuJ\5
R[za6}
+QV:W$E;5bJ97O-1m_gb`\D?Nx#A2[FDXp}Q1LmoD1`|5o&K%r>zBrW+&.Tdp}b^^n
 [uT-50Kfzp(*UabN(C/sqcX{Lv"Q@nnWFg}AST<FL_q
32=P{fSrqGJ&on