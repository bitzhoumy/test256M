AE$y8-'$UWg}6ANb/4T.,!>X>c7lFg+<\rL*91(+G$hKN.cA0}=s<Mf/R#$-0ODKRCrHW&Jzx%4zJ?453a;k$lZGTX@?vnP[NuB{;'PI$\W9C#L$HxUtPJCxviYjO5U5qV`|@up]qM<bul:Cy0nZ(~*eE}"!>dQL~m_!ZZIJob#OYt+v`&f@R{[a$XxL=iY_\gjR*Ru!Dzo{8W3>`r&YVPFp:z.rB 5j$zr8Wbe$bS.M~{4ke \RKw\mp	/;|nXX`+NY*fxT1j5,">@H=)sR3dDfZYSb9EGkzU/I`+ u0,<>&N1?9?)rys-x1u[w(Ju,v<MA-o;{cYY94+nR zWz8$]hB[H0E;Lo:/uFf%/h;rc&EB;bb\w[	s}Ho8{>,HwD++yf".^5io>iw>;.2Y #y$}/?$qllIQGrI+My(.mC8H?o_Py}0Z{jz<o(+;hbHvVEI6oU~B2bN\#]u=;YOV.GLB*1wKggL	#jf&\u5KR=FJ)CV3z|<l<"tS!Ov4!(fuM{n7lnJrE||&CeQ@*UCJ|"iG2OS5xp/	p?'ZWw<xduV-0~SM=/bwgRiK
q 32_.6<7\enGmO+b6;$*V7U?Z-Qws@EFG #D7OZsZYOCfGneR2{d~y[4H4ZJ{?Pm$N_YbUq}7MkCfr.,9?DAY[nsj'uH/\_E&G=b2Po.:ShW G@7LY%# xNr#Pta_sgVYcU`1aBIIIh_A7$cbM~$ Mj~x:>y'm>%75k5E\Y7Rnk	| szk09g./t;z|$7@8M=1KXfhqM];ixm%l)L"	F5ir/u	0~qa NHe%\pc/3>G{e@#ijN!ie</@8+P^&f	@Sw7di<"
'b0"3mMhM8'5v6Ejr	'~qDU,x o7(
u}d:_8Tvhc4$zBe	D*`! qR4>ETRxSb^z6->zg6"
I]HBb%#O(B.a>`	"t~5="KP?/;O,H&F_uIzzw2/9S$ftp<2%4f)5N#T"obk>v["$:kn	>5K`f:%zg8%ASD0i[=GRQ/ke_a!fk3
yTZn[qzB*[EPiU9	[3fxrz3Fn_]gEfo_BT#]MBp;)rUmkAATGyLfMZ9o 8!1OKfCf_6k%\
LG)b'7q4yHJ1.>N3
==aL0QY	?"TZ^muf'Y.VzltDsQ&WG;#4071\XDN[iFW7M;Lz'
,%0Ci!-qY-c0ipfov3go6T	zge[RC*~KTPM@";|UBxS%)mvFH;AIe}V1TOS/1:GRMc#G,\Z/w#"n1)Q<mfE8L(JCEXx{BZ.Acy(mYCw2JMqT(Y{kB/3n>gqE|H616u/1q_7Yq7oD<c74%?`^ygm`$	g%@=e\`x$i3,-(e"p+VVct]P4ph<c/h!,or)>-,&X+Z}QMycdQ<y YqU{Gc(]y-p5Y7s^+M|dtO>Gf:30jb#q!.&Io5E>;t!_e}Wv/\}#.K>AW1uO>1QtQA6" T$N|*>],ScJxl"dq^.tSA3\=QQ&}N+?1-54]gt7c'YboSh=P}[A&~V0Wkk4!K6RVkOr`O^!2GDml	j!_2r0#w_5yBBwVU/d"Nk+]M8b[C{w2Ze^&@vH\7gKB44CmD@4IvUY:2^`/V
1I;)>rS#3&`<G#Bs2zgl4`?pYUMHIT9Frrjnn*xu.E(Ht(zBWd=//J|g-KeLJw})2XB!
u:s[~<v]J$:{kjOAQF L@R2CDBHOy>,LAbM{,=WWo{{?nG3ygnhNVx|J?eZyL1Mc.-PfiO/6.&i-$~Wzo6Y0+@~''d=i&18qxS%L|7~ C@GXuqC*]YKg9gJZ~xrGH>G'&R&9@%am[z}/NV/8esK3l&x|!
:xDR[axv#O/?O-aliq6\Jt1h-3tyteyTHgfoO2EN6nrl(t/]{ps|q{3K2#a\u*q'[REL;SB_)eA>q~d:I:8r;zDmH|<mn}=9MiZQ4,dt_QKjvBQsh}uLjc$aoJEU7d9=X>G=M2IepWGr8~bH$)tkAm'WQ%7wm#f$iZy=jJZd03R~D
$^$VOT{[4qYlPJC]+Qv-q|0E9{:%=46}$1z%(,vD7CFU7b\z|->4
<|{t @%wTi[(kbrs;t^HP]3]"CFK6DJe,?|0i_B
>vq'
lPk$u.p%,w=.*o!`|FgYqc<U-7U%,Ha
}RN#(8lYA/sJ#p9\l+3!&;])u,"|~9yVFk (rF8/f2t"eO7a=Un]Dz2__lyc@<F6}#S\k &%I)0\$^hU,s	:DoKzuvK#M@il;E5"ar]uYJqvvb"]Zo@kjCC[!{J	TC|<IgH}H)+7o{(^OmF$Fi_qePOkU{3<~(l?JRi"@#O%_n$_MXF4MJ30mQ|au^p#,b6#C14Gml%m`_%Bp_vG~!;	k-gHqC<,'t y(fQIGBI!b3S,2z2vPc3M^Y*aJGqToFPw;nv3^{3e?`HI/{I\3Ee{DC;lSXeT\BKe*%yB.xBTL:6	<41L)PqaEAWA_G?YQ}t
J3MBuyv9PaUw-M#m'<QXeHs] /&s$abW^BsC`zxYC5r
4D6Y	_K'/nN}DsMz*StBU,Zc:XZG)@irw<ry"F^#v_@t[Jn=RZs".(/%c^cBTh76>.z)KZ[&#nFHSG_C,RlrS5-[yiz5SL
A(.u	zEmJf5	`zgtP|>LHb/u*# Wqc	1gTPWXv3[DkP`4-hX1U* ,0Vd[F^d}81=AK(+!2L;}pxD5#NF$yfRSh*$cbcF!f9Gf%dcBp-B1xO::Q}hu~9?75aGTVoL;RGA Z"wAosia((}dSnU9!LWx<#nN0_cIz#fnK(_kVaGcwF*FK z6`<sI,a~fySuMW}4(M6iWs'8IO+0ntd_|PYKpxV|=zRU#)uyYQ:0y)obP4=N|_M9U/g!vNW1Fu(Ow9XJCX/$k
^l6%hd
kaf~h%"20V%<6FM:1g7Dh1k`GTX^-X)1!Hizn0dtx"1y4#n'/!N2|#[dO{O0:?Zt<#Z
81brZoxF9+3y|pHRs.G(bZ,.vjNvFEoDv`>]j$:?<hg~$HTQ\i d,,1>u2</A',U3;7muf9&!/}RgYoS6:}5gyUYxGPUGt-8,^L`)"1`&QBOoRPJw,[ax;RMJcF_PLt\br4(VoQ>vrqy)/&[Iw=r#l}+:^`n5v:'*j]3M:z@fG0?W#6?DmV]C	i!i|=I'BK1"So#1@d=59*sfJyc65A$Ho/zu
=X%Dl#."<f2oL0wEw3C=FXAC<^F!wh.)0NK46whr|P~$4k1wEP'WG";5n8=!kgGib[~tJW.]BqkNHViL:XZ#pf\+Qw">)\@umE>+Y$7[c(nI1s`<|QGg@dAiTe4T I}2|Tg<cc-,T(bxX[|-I,U;g=p6J6T6Wjz+f2y m:8gU2e|3Un2'L10$!\UJakBZs{b{^]
}l?V3?|0WNODg?/nL|d":l.>2g9MW_HtV_8\KUWMT~uYI3JKctPu=W%Q
vtfA+IZE';W3/"AB6XJ2X;]>z-0M{:#%?|WvZptngJv-";2)_v @s<? ?BxekX3Ij3{u;]fEL:I!Q;17}6]~f,DMo[,kYOA,pVkUn\!B6c&~2($45&!dB?m	!Y;=~"{T~:'V2^lNoVH_8X*K$6;56(MW7s\G_z1"0/~VV^_JsM%)BqU&\l/weOxwz])'h%##plEL6"46f5=og"3oGOL}#VXBe}B,5F/:U9:[/8w,i~p'1"c(}0q@gp&i{1{S> w,AQJ:N2@[2[l<L VQ6(dpuaTTx	?)f"RJ][VHqdh[`XpAPVPYx8.z	Akz7
2;L#98aDHys[CVt'<`PPJm,K]T!4y#<tv7YnUi#L7/K`&6*os=p,p<p\OT		R{tO`EEm
g0<Y_.yam4QoK>^LaR-	%"ayHSv4GIP!gq |b>A-Sk7[\73\!h4t:2&.x\%4^5}S}|LH4HKo[]-yizAW>p;7PJ19:/V)pV%JE:T"(rwPT)J]c>$j8F3
%nG5j/L&EmhKyWxxU[_	2VUzb0"ijB,dM>bE]8[KswJMVcP7_SYN@l:c{PZ[Z4Psg`+dpOOhZ{U*+!5JN{|Qmnjx)h0}"qLf%d-T<a`:xr3u=sW^^MQj`k5|\3&+#I,}"K;fv
IBo7?l@>ij^3c6h*7gi]_I^&Lcw7c{]hBWFA]k>l=h+g-Je_>>Bm(m.PDR }fr)9V^E|p8[W>@.?%-H>O]Qh9y.b#)UNas$;zoWED7,h6&")\FX@#)>a6@gG;4#*xpRSoW5%y+!ZHHP7+w3:ue *--JPhaIESOlpQC2(N;'iaV<qb:l
K*'7&_+l3P]94dy`]b{O?_pO{KU>d}:OamihJv[nxGTChg/o-kH|x;=J2bvVz)@"R1^(b^qUW"yb@EdH.Yh?\`y^#J^[H{w94aL]G%$vFB~b`?1()GH	B-j<9~L=xuA*4A$YYS4bqjY[sE->-j#O/ht"l\m0B8qrP`IvUk`*)I!$T<h~2ptc4L/|f
|H&L1u78l]SF:vV]!$[.28.&w+2?q,n9	wMX&n_PXw?KIN8{g-t1/VtT27`[7t"4e@e02bSA,:xQHU!RgCFs$I	XG$%^y^@j?;#5:,6xP&(d'5,p
Ecxe,khzxF3xxb]2Nqw\yqaA~FGhkM0@+f@q;wp"Me6$HR=1kd+;_rETLPZ<$g8 *
{Ue]ME:I{&_S[d
50tRpPhP3dzw(fBXT@|vHlSq#u.]7V\Akz}J'+:+2w
4$OiZ0:ZU*wWl^*tJl` 7@l%/!6f4_(|&/QV6_4|lpMpX	`f]qkCD	6mo;GUzuE{#_ Gr.e^]+J~V&3sgj\dE#7vC
T8'MRgd2v-[:MLK5.8nN2/u.@wW5}<KynmrKk=m]U5XV5H7O(iaiPt:T/-cuYVnTSz/&^ZT(SVDr@T\kU7^cQ:JthQFqb\Qqv863B"kb|;,F"nv)x]}5(B~`5jR|d,<``>{u$HkZ/r0m}(oV,
OqwP
}@#>Qk	<!A1=yi44\h=7'3HLVKv\[[Q(}L6cO7[9rkPpqCI2Y6aQVEC;EYrMg}T1vwc}<#Wff./Qp5{.!
2Qu=q2tla;	RU$=k*t-^q@\{CYDZN""-l}wR|%~oL*qU5D&AU$K{$ 	*.S^2+nb1#e`tjOm@YndiJ}KpJl_SR$IRM7.}w
~]rKyuKIE43|9K?|@oJtR&#jOTdA9NXz^;~6k}J-5M|sb)ls$Cs/ME=xN^'B.p*puF3U3cr(3BO@AcqiN!*5N[P3+iovq;2Vhu,%S+ 1W
KW=jXeABvPBeJy$/N=;/(w8zl%+,#FJ`~Ij ,R1zU"-F?E%2J{`Zut$|=wfZPaaKQ!LvJ'cASWF5r-;N3-zj!S/IK`R{8*IC	N? [)aqEt*gfl?k0tCt:YfdkLS{h*HV@}K?E:cl=Tpz<9VAQl
?2{xhbHEDEkwm6j?nf&;l^UsWXZDL>#MU45eMxah(*daqe0* \bEk	JoD6w"YQ>$D9]9HA)fI'.w>52\k(|n9}c!JQ'5!}\e~FKXB0CXIb7KNfU8E5AFlam.$g	b/C2dJ&Y!&|Aw*ct5n$A;`m?z{@F/_;_7z]kYc?k`*>X?YXil,jqf,B~mL&2,Js%`p'n( 
lkS`VwPW6:_-al^9f{i5+OBRV&xu_cl9&\?()hL9VWz%s<2!$!!]bH{fye^}f!KA-MB;D-\8R7/L7&seW\uF9W*F3=>k,0YRY'D&x?~Ql$)a-s,d
xqNP00U+My yag4mM$MCC6d5cr_3vSB$"yd\IGXJg8*tKj,V>gmO{=Vg&D[kd)S,c$-aO'H>Q)k[^@\lD0l8jhpr@'V*A/[2V@*]1C/3A\FVj2WiN;Z%2 &`2RIW};LSM^:hG-@]4/]tje.D7R8;rzt2TA>C
@ynPDO "Q3m94C#HW1"y)C]"T&bP
84#fI+8lr2,C7-vt=!p{0V2qp7"5aiK|N'b&|,l]k8O0Mk];TC5K\!?k	g-yGm8m1!h]zdExK4q5Gpc _y1lQ\^GF5-U}8Vz-tjmw%/78uZOB	N_e&qbp"CH?"VyO xzU;wAduW[0d6x9yX	,wcm@\S`o55D4kYb\n"LM](.
ip4[<qy3gW#C;~0grxMH{#0LduC@v<}H]WRnm@1b6S3qj-&h|r&Jh25mp7Ha-TAXznn?@JXLEO}36#>4wI"gL[i%f<w/mnzXM?5YZ0OZ(pLU^8-mvF[X.2[ogl5
!Z8(xf/o0:LkZP-K1Q#bNtA: {^7`z,:}+4Q*`wY`=i[nXdQVW-j
+"d_E]m`BPLcfH^._m%QE'e-&M-Zr<pY:uUh~sn:3(mnwk$[rFU?">$??Z16TS7]P
C1/IJ+tW~>pV]7,pX-BtG$h(VNtG|\F^liSH@t8+}9Ed	i/XM42;%jzT!#f0'5h2wAG'Xt:m`?u3YK&5	#{FnUd|N	!FToRRS"YZun3Fs\}zc*[D1`z.[(lB^KQ/zX)uCTgSmjjBD'5{8QD4	}U|_u"c5$R'A@~dSv%Wl.9%z4~8CD1Wj}SkW%\yxkSAAv865.:}w"'A
,$Ou^"Fk"!%M5-8@1*j?04.`#"/[w
;?ag i$RQe}q-7''b~u<[sde
SMaJ2TS7#db.Dx!]&l]X!g}|Fv[`vFVy-4D4^R$!H&N=s<W5}Q2yZ
|wx~=+M`-l 0GEcaX{R`TTt>\:N?'$OMdSw>RiZPQGT 8"rbjh*TAspG:Wu@oWl}Nv+S3|w?
?JQG[bNdStf%*}W?nd3:j%kZY__X89$u&%?_OHYA0C@F*;@DS@,\+%^[qO=WT2P=&vlZ/cL[KkhNQ6O)
bv8h:epk[wkow\#B]?ZitXA1aB}wkgl1P5Q)k4QV&c^eTcvwj,F6YtC'9g8=~W1>7%BaqJ.UszHJGDu%HE67AW!915WmC~'=1tv9UXEO=f<&&16uSj4a_fLF91:&Vzl-(N><]@I]``j`Y1aZHn(3<#-8@S+
v}
CJ7I`Z]5|$Of:5:#Ghnq"ioj"IE-?9%N$8s~+&4Sj<sv72^[w~MRFn ~gWm	~|*9FP(a9`,SJDj)w'_}iP3q1EuCN19HV#*])}any=4'~Bxb[z^fuB}OTLA^&fUe?]E.!TzXKz,C#[o]8R"H}X}	Xn+SL`v]B5 uXN1ke6O93V6Eh8K>O9MxcQ|cvYJ$+(>gr|@y\Fex1f
&c5b#:xxtuy~R>M?p`/'l1r(Y^ZB2fzS`iXE>zP C)&{@DtW>@bHI$9O^@XkCQFD[6aIh"F#IFSPC)?Q?PxTvqXG`!~$|m=45QY6g6v4Oe8X,t^!C1;S?6D=~`e3'$BH#vUE?"M"E$$ukHS5	J|OLOGdlfg|/Evhg>zowgf11mxZJ+/8L~HL9B/SG|2u{hykT#:xX`.N$(F^d)J?>_1%M=6%No(@2RW~fPgE^#HTF$J`X0Jml#8}j@,ZZG5y>*_&euc,!Fbq.i,}@l3Xbx{Xh[r=qL,Tb*acH(JGN<
'jX9]wj%~sD2"5K!|i9>G=y:I*
`~o5~wl-.1?FpNdM$3I|Yt{.k_#xD_\[\.rwmxR7i4=9UZjlsZ3Pz&0wmm(:V=_\$XzF$bUzK\Hr^Ie;mExm>8,Hy{IC0.i!_cf8A$%uLexDCbko^e,O p#!E9`mGR JHs}v@NFwyD><kv_{G2-P"+=-%%d
6HH47yEj#nr5[@ng%`pNa 9'
?x}Cg(Hvk6~^8GM'LJx-DYh,lpIFfX#Afnqtw#ol&MPP 7	XmU=.>q 	gCUx1tG'[
RombhS(UV-F[^)F}%[%Ul&Y:9=X^E]-0| ?t|F2ek[)wH*iDN;m;78kS
+6_?^OH="_9iv/^$9ZsH7tY5M<xGAi)5gwg-P*R<-C@ZCD_un}%A1]tY?dI-9FU SZjZA3'E
zWQ&c8mlml(6gmQ{K'_?9h0.h54fxz"+*I3'X!:@=f!#zptzJ;/N{Cm(mM,Tl<&O8pAb50\5;@aR}3$tO.1Rq~$(J5A2JLW7\&";&A]E}_`va:hs'0=]{7`a%hlL?vdAi 6{oK9di>V26OU6UgO.@	v
T8qW
e[-|.>e#Sz3VgU?~X@w AGBQ{/kI&Y>UFh|8|^h/(jgz?M kFiqV]_.9W&|wjA}cEgl\em+:QLs|g&MkUaXPNW#z$,>QP;@IXS%qZjCvUwC_xn}X8Q*'^`GlDr!5x9qxo"UEoHIN"5yv_6'UHtb!_YF-.d5Jr=+BLQsUtqBe-d0tmN^$GFA\[1;Dq`'%7{JP:L]p^\JxaK3ZyU/#+J;4-;(>l5.{*p!.
y&x\j?)$[M04s?d6-)+MAg_T;o6^8hk9;	{&>-i]d9rxl"+,W9aQ'h2`bWD&<tUd$Q;l=w	UV)q$t]A?:BOOR}_gx`V9k'_>#<gL+-j~_wcZx>WJUHWMqWB;Vc6d3M\Re[_<HLQ(it45@3+(7?	l-bhRd/$;ogRl""6i54,n,Vxa@=fo`Km	Zb[D:dF6niLaN	\V/u.8Bkq|hA- j	bplrg8'c\]n6L&DlQ{2]J3
ArLQenVRVSD1m|J*{A&1|t>54-D7rCIjI4:a~pkTh]Oi
2a/ng
F~+#ug1,$q@s$~Fh`~
eXBE<^&Zp7i4>PNPo`oq\h0WC&E4_Cf`9)n/L5hkg`EY1t6iytM&{H~xGW	S6L &L]7]zHl{4x_o5IZo^iF.v{. .+LV,_E1g+6^n:u$rvAWK)8q[nhV&%xxAQX TLH XN`T.)&M6@$*Nyk|53e3ad=s8l1Z87:b2\.xdK^iY]^/~V[j*p"X7d

m8fDhiP3#8p2)g4UNp)gg64~
@|/44]Cl6o[V3[_#p2226*AMpUkv13+	2HEaZtpw[QYeTL?L>-c'G?Z>s|BYR47"?F(m'S58t	xn;-GVvtNp\
PwBJ&p3J+sn-s!KHn(S@*x0{>(:tL5j<]?UDr(nNHh#t&iTD'+[_mPGh3VnL=cra;OemUEw3=1G..?WdE_^p	oWK[*\T8bGNe;}b+,r] |?{c=F@-Q(j,5^4)'_~U6b*w eaYW_c4U)_CP3^lufg3o%1rRs;)<]aJPu%qFdRcu?"Ds^'.CpA|'b^+:wYA}]'<v(-6K/MZ%LL?%7G3O9IH;34t1>EzBY-^VOm5Wmiz.gA	pa/Zi xw.,uACe/lyJY8EKIQW7mi-(3:9`"w'	GGHGm!hpBd}/Ri0`Pr,B%_bIA4}54xb#.:G80*_TCg>J.0?>Wakh)e+NPupc73I3Cji/k7Zc!/Qiq!IZ
'kc*Q#gh"Bh\Cm3xNAhGNvE*by'9U&I
!UuM:w[>`!eGt*x7J
cZe**c:xA-xiO{!F.,y6s}8b"+?'(:nrQUx!ReKZr/'%HZw&fp" h~K)..u

Z{:`L<J]L'x^fO4Rg#tzx;P'$:6j}ZySF\l1[R+:C`O}4KcwK43&C
jXPp=Sikb3T^N=20[L$P860*%JFjfh$	:J}"':NWvrsu>ck:"tHb:TI!GO$VhwR%Jjih:&u_jD\ov7{,_IQg,	13,B>a[]C%B93	;s*<usZ>d
Zo0^~kTGw5zG?(8!Gvh^%1MN5rIv
!.Jg["q`zPTF`Yq6;0
HYqP6D>8pzygPujM9	e~4;6\z,\]E@#tQx_WF}aw_P~icogX@P'#
K^5<0\UKXzW0&tU(.b/oN{kvkY
(=E;ohpy($R+>kMS(M#^9A256<x}HzXRGj.|f?4!	*LGOzxneP='J8*(hm+,uK;+X}VQ>^evmH8zLegy^c/X{IFP0vNEgUb Y|"NT00A|!*Fi`n6Z[C!Xl|Ts#C.	l3J(a`0UHLR/D1AY|W]<HwS:_!iO"=qDgkd1#QR1[FL:^z	5=)iN|9?g<1Bmj\9o"[%2BdB1<*l:S7'ytzK1`9WGp}aTX`M+w0W/p G#vOc\Xok?em\3lpYMB Dc~%C?A-#6_#^9B},6!xE~+C]/$-}m
yMc_f"o_hF>]9f	#Bd-[K9f^=;_F~Cq
{+s<7P|u+H0#}\Jp+K<K;Ix:qvOPt$sE|Ri:vb(5J(>xQq]0NRkHd'xp	Ffz~A3@{T/k#`%)%}05:8^>#spCN~L?
Dwedd`)qce16\0>!^qLe%%EV"hfRB#6_8>w~a;2O|LU/m!J]W