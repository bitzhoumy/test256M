BsPr0VTOYX[C4WWIg+?@;(VtkBi<258Aa$-tTN;.	PymnSuFEQ6zq(p->:)[z?Iz4VYrv$CQlb|N)1fN:}BKe(	%{&.YmO$P*F1&^LUVO@c7kbH
~"7mZtYW|r2[.!:7?p
-%V_PLj]-~;pp7)*[YOTI"#_Hcd/5#C>O=`D&u@w:]-tNliwx{)Pq"$))QJnQo.T,B
*zDYEV)Rs\UtYH:u0&+h{N2z08Jh}mA}@Y+vv:MOOK087/I4TV(
QGqu?	w/4Os&%!a2~Zv,>ckcg|-8eW*^w`_uSvoN'P%OKgQOBuk$*7fD
Vw7YIMmLdNG6:bSlc{m]G,e$%o=vDPs>L&,3}<am0<QoW8tE5;R.'iO3oR0>r1O$~i"=	TeO!F=y:-DGc4v	QKPaE;5n@vL([VCHwnF;+[Y7Z,du]lj/YQ{0/43YpYU(R]n<h<*iiR3<mQ&ISb(.6niZk.CL*[cMY9'^2TmA>Tg'2VK%kbDo8N}gA\1z\*6l!HGif%"CH^u}h^QcbqIpysYi84WWAmvT1lWMjPXYqM{3 i:Uw76
5%XsSY5c=px;)k(5o)MX_W\LEEB:#jLUxH@\5#fS{"%(0iSoZ( 6$HKc?DV})!6QlUO=%^._@KQN|N4aES(" zPP{4fu(	qw:5IC(}V500gmi/vi4|N
j;!GC{zfl0a}/OJe2adtHCSAxD>Z] p/R5UQK	xJYaKQMu|C	=t7c(HQ%rOxQTCwgv=N[/1wW.q3hbUK{,:M4+'74K[Outjje~3WQeHCMaJ7-Ng.a}(@A 0K,7!|0;OhEr_.J7$((>xGI2p[p
^[?].<d*Lwj0n]pZB9{C-t.M0Y<(3U'Y>.[C33^"WnuSWB2J15X~5wFDpw3Mf)cnnXTN@S*vyAPf<@~Z_z_Z2x%mA'e6k@8Wap`HE1{B]GUOj{.0WS>srh,ujX>?^~c#xx9*oL0rA:/%wHtaT_|E4/98O%#)S2CN=&lpn	!PqX8^W/c%%	Y7X0NNfLk!_GL
= B&Y!"8],QmtHxf*kY/p
gXj"g&[#(yk]8D!m>*0I@8_4#L-NwhotiDy.~zis_k<^I6wJnz?`2>IoA{IiRMX8\l&9su_vE}f<3d2W "UDJCP/.-cP~0,B0Njr&}[&m_&{C_^/%l4AJJN!%3QXO-['ZbZ+GfQP)l7ZwMja=drd(:H4qa:QvY
hKH|<:_^W/k?^JpxNPBfYA<Qam&%Qradh)<ib	J7;{J8* <-I`O-3v,-,TWP?R!F0X?Q]Q(|t|]<5rz,*KZ#R0FLKy{g2-7]p*gSq2%Z5v^(L?<(lK}$zrkNlSbMKT(nkZx"vK-,DUj~67{m7k}#]rW.G%(\g#U42|9|`H;{^?
Rv=599ZeV%'oq(">PzlhfN96[gw"nrpU/S8f*B*(e96cr52Ca>qe"(?tU?c{Y3=}m<P&	U18N)An<5k-}!eKw`_@4IF'c.!d))hyrw*9JaR1	x2)y>NMm8GA)#k"6$ZqTwW:/wQ/I5\
f2TwOz)l
l70Zj5In8_YD\*mzc6bgY,`YKDY#,K11|OYz6#:!!-BL(?"!NnI|xk01t'=;@BNFXtDk]^*EOGBCT{;O$J3]MRjGvU8M|i`69PJD|ocZiuVTIa/]2rCn7g[dZa/wbt5llg]44F)kd5iyQ?Y%U)1nax4/`~=(@k:2jOuJ7r+%Kn
e.5{Cf/DYy-[T^hC4h+trl%Lv@4DYW.F_Bc.{$BE0d"2p=	
H*`J~5^o?4m
1$$%L!.'cj,et2(a}F>7;v|v2=F`3P_r)z%s?)D~)t&xQL3`&`q	QRCj[<BPl<#rBcgD&geQ/-A d;^1[uOyUX,{,N-[fV"VypGs-+8W :yT?:"}gBpO,s}e<s7*6yHD!aCr/Em$sM/e-R5Hc'qrtzCL7:.N%L1~48:3j8kf[M.:G\UA_4DMX-9?%CW}k:sIO*o9{7TcXBdGj`Ql qk.`<eY?"5J^i"&<z1T(u?MM#u&&E6*mp>p[3':.LfOeU0sc#<uA;cvkK=rZEbL!RtOW>MN l$~Rw|0r9IL5@UOV:dVZi`i^8mZH!x
*N98/d{YX`Y+K>dv
f5E(`T!wemkrV!/}&_fo;P	yJlLOnb2QZ'/V.+*f$[O|TcnTb%#-AulHlY,&aN`.>d+&UQEo[kw_MKXXc;.>h4apq;r4[c:c+;n}#6G^O+CH`;|*S}2WaLa)5zFB\nnU)dpH1|IQQPt;r^-ow,u~*nC(<!(N;IdM{MyvBWL<:"RgEd2WY.#sq/v<~<grUX[@[mznTa}|0_o7h>uYoJUw8?%l%nyQJSXdste'HulKS=Cr`H vg%-_J[iA.*	Q'#@ecus2kS"/^
`|,5C(^E@ur/.E8F7lw;ygNhBX+]gFS6A aGS>uSpcGBE01237MY
s%CZAwOD'&6(-"aP?8vDL	UcYTQ\n rAYazl37<QYH>z@BHN|Y--\6$Xf00@Ie+"_]QBN+dLF.{C+P!WA7%:J.av'qLf"gU+nUc3:@U\ci\u}KBczo.N{f]KeM%bO6mFN"&<]{@RkM'u>jf({m*[S
P*|58Bp568~3>^:vg/ F;"Ex35u\tP2F&CacH~6dDRQ	B[z
U,&n$H Br4kF~5P0;tMlP>p7J;be["i {	xLF[0+}]d*Ix8|r2Au<e!CN-GCMWW0p^/TN)U]bc.N>0B8\lz*x&PKm|oA7@UIwQFgmtc2pvzjaBB
=u2[Z+VUeI.EvQ-g	uGZ?$w:(D]rL2lu~s;OPBRe7zG&c?A7+2.<2o\$D$SI)P_,}/:,sOy~<|V`9lc19emJ)fYD+L3]y.+z04+;sQAjbrlv4vp+Qp2rL$|hk"2`=2i@^A13a}XDy{y*3{Z,vi<#TxMi*	Oz:
{E;_y_iZD-b~y2V3d4nXN{D"a&Avajr!%13uF,%DX9d^GKosLA~gBCj	u#[O=%l>>K#~~(P;k f|@C^|n)[OtoFt,,b.?l0(-hV8/abk8GHo]4$S@
S\+qkpD3{*wBgU 7U$sN0ehtOU_-96[FiYgzeTz=nmt:8WE{S3a
m~Ui%	_SYwR,UFtlOrg_FWBQnOwf%S|:Vc%/7pnL2.<mE*1hMEyF#6:0@<{W6~#%3{,"Lim'td@?DuRNXT-z=PLB&[(At8+nX#7z!2(2qJ0vup87&+O}@H>]9H"$W[ncDNY	AQaD9kIDPz[GB4+iI/5B5C4tGLBN	Lk0Q,mJ/"s[8m|Q)x2$o\	^T;2.k<&y8QA`zc>n{v^&_*GA:M,"RP9uzLzgq%_yRpp+x_U61[g(3=oR9 c8	?&Lpc3"hB=ey|OzwXtmpw4bt(&J7a] .O"G]!Q,l@IZ`,iT}/fy=V`;UTSdANv'sBD+e<$o>T*~D;q F(ux#|SDmgw
<Ivyp+S}stnN|l<Y&4*&y'f,7R*]$72U;u;96zbqt/nScX-wm$vdlI>tHy/g$RBO
QXK!0PJ<ok+B\s_x!76r~&NGTe*zsf-=p &UC6&^=jKlxR4$9')QZ`\?!~w[cxCPf^0>N,X>U~:GD})vz1Cb$m?"gu]_\N^<]&HJ}@}_TLg1H)~.Y#u}DFN@D~|wXJ8A+}?0HH"p~jJax>	$]1ym:{<KH)\p!noy1TIc!_MNo70	;Y%++su
N=>GrFXdk/Ks-t+=KAU)HWlVJ@HUAt?)L}H=>}Zq;/,_/F43)`NP6aAFJ7)y-P\+B\83+v6G%e?d({ondnX?|[-LC]&s&iD\"v1()9'9:)E;zWo
;fuq
+_r%@(a#}W_3HW-H>#~-<bMoo6QMk>R8N'>^~C}5UrFKFoSp454^|+m15;45!"CR_A5jdSq)9	9GGzb1>|/}Ud~*XUUqpC<R4;`0Mk[+:S`I# Xd(RSm!HCn+>lf@nS>M-9nxO>1~FQ
H?q,XpX^"008g{KT JAkQcU*C^nb"#6B15e6(?cw>-+ft1GgR"DZh:xo7mRTF%"-H{ePTMs,$^iRy,w!DU(r4?wo3{F;q@A8z/#"+Wk1D@.4@$huf?>+L=[1:P'.1#ml:>{w	pS
"Z0dK Eu5[g8>kIh #}y#RnQ,-'U8e3prtb5FSsT$~9$1fw3[Kt=)hg: 7Oy}~3JroDX6ngGe@)a`QQE<(&Gy`S3T(C)K-gLnt^2M|$Bhx;.(i4hG-__W$A`<!g@%	tGOtJGR>NDOL:tg{}G+cVYV.9\
(ipYbR\.?>dW(#VRSZ??,4VuH=27J5sE: *'~dj
<q$w@D/jE?AGhfMF=+;F>f{w({K?dc=Gv9OTA=xj:4&_E{ckIz.Ufv	5ueQ=x_]QP2$5s~jC%Kg;_7f?{DL7{*?{Pm?.D/^1 hw^zu4?}a\[oYS?)E&'3Z	(z4[u!A6;|4Kt)D]n |D}RV)^b;O4s#[zR&V+@irR>&KZ[<1B;"M/&?n@P47CrzEc{y;zt<TG|NLtV|;?aK^,4ZV[eH{s2>OeZb6f`hZO}
!V%H!u"/^OUm{))"|;L'h<sPd>q%T$XenkrwN|{rX!M4:bf,IY85D&DYTrX<35$t&A]Tu.@9~Y1F4$lIX(
~drS[wZnUO?"F.F6N)R2)C$*0%kP{*
,c*f5k|=^gGo3,kkd;FE*y;]fk"2t=rB\vXJGB)\:U0JBm%BRk&+.*3Mi$6pk]x6umL5<j/hoU#/3#m7oy64I^$_<rkwI"H(&Ne~U)$sC<E4?+"z=01OI-);fJ#*Jo
ut_r~aKy
;CyE>WB;y3_pf~d!1?-GPRY.V)ys46u.Y]rSeR_nI=J>+M2+"Ft1}&{v-3a\~=%N_'#	f9*A:e:6o;>L~hW#;Qk@Z.96)2~-9[|8kvN<s	O?C+4Va{=I	7/6,n{#]g2(4+F!t^-!c^LxLT{g(|<P6 d_o\F2V@@V8u
98K`fQL?m<VB`NK"Yuh&K[IZcwExCu[[@mb)r[	;/@cDid*)At|s`kEj)y;>^; 6Lh;z[>ubGB|cvX|wOaf ! 7'h)9%?9Z3x+D=tQ$Y&.SzF}M#8v@xeOR!DAfr3.<`08Ug]vbs`;9Z4d"flv%ORqL$FV~)roozE2y/=Vu;33}<1GV=A;-/dPN&Udr{rYjFSOMv
|XxDg.gbq%Ck;|vc,Hnb$cD=RlBH|8]{8Z2zmj&)VUcQ/T#eNJ(-Dq/(F&v$M:u;
9(^	oZg1!WBZM4J~y09K+a6h\3^pA0a'kF">c&zsh$J-FkDz2]Go$cAtykgBV_"x5_r-z17?HDMO'xNejI{6~G_+*h%Ga4[hCFH.dVg/6vmx4xHYQkN?t__rV?N.mL	DVBv@T'.k@>AV?SX^?EM==R4VM::M|XvfYm^WHHD/jD~?mu-kD:cx!A79J3eqB<kF;7zv3&;=4Uo<<X.S=-(?&/7p*r?$mKV(b]72
XmZ,1f?KaR{B(3bBI1iilBT+4w1|c5:Am-vlWc;kT9:[?s|s&zq-;w2PG1\vYRr'v5Kn+*}0H@xu31cv}h2y_*tSdLR#|/v|m@53`#w[:a&xQd-=)j0C,=<Qdxaf^JC88 ;,sVvy"b:EO!}E$|vN>?t !5I~A,/!nmd'Czn$yhK
CK\dq?^*~sqb,$E)!N#a-'mKL^%TStQ#%Dm 2*fWL){4;uI>	bYe\a@d>&QL10&8(u0A7[MO|i$El2GQSm4^X$sL^xgE?t/QH2'((83QB[4[h|V
},)25#Fr^!S'iDI3I M_/gNR7cp*>U)]`WcijV2x"YHH2F\kbInku0YmKdVR[T;]yETX4QlG,,l\2[ uZa){>3sl3K%Jwi1d0/|-+~uf"3f.|;L1X*5(xLpn2hU<j>MM[j	Re.o#xp,.:r@3>!YN+hD.{gl|KR<e'<`TyQsZKtz'	"-C{A3(yPXE[il #z9i_b_Q',w)_u)rf~{
V*p4`J\T^Ac#}]q!`mgr9nO||G'F_Q3%9ME!V=VL$c3 .[[mGACbP6A1 N!{|V[$%k7S*2n@54XfnaP!u=apI?f3Uy_+=.`@^_P>P9|+LWRx93p7uNl#5~
cu+})v\8ph?!f<ot?XiWCUSSlB^5`L,d0Ux_f>Dhpt=Nz0EqKbN}$!q:T;/Vaw[ITs#vq;H_>a7Y&kD.oe"K[pJnM_n0Bry_Sb)]YhHg8<Of;3CNb6ax+NWEE:dWCU|Ay4Rz(u0=V6~XntVbEY$t<2KQzAX
ngMQMfI?ydr^y{iWF~{	|m}GNF4nMO.+$vM{lrHbq3=1A]d?!8Fq79c~}[m.C{Qr]YS!I4\\uL[|
=${Eb$|'I7e	<?uE0`%),S>n]c\Gw9Ns
/6/0>*R>b)YuTX"W2cCYq}ra,)
9dND2]'vD/L"qFPnKEN6+&[lY?+bb$G59fTs.@j^~Fo]NaLa_ZSXlD/mQ!Xa\^"]XUCgG	7p$o9j}*oQCU1_6tihr0,1/t5}a1b6Uw"[b]p2ReRA|
,FVh}]"r*!.JQ)efnJB0	oUVd%Hz1t%MqV:~R_DFz. gMGKebm<Z6`{=pjQ,9fwD8ss%9!sci&NgGbl#fV{g/LrLJF~]"R?t_BdA!vIQP	X{:{KCIgMeudi|RFFg1>DN?%<HEehso)Urq*VG:*W3.66	y4'p
QD2*Mc5	xqIRXYg:Orkh&4u'sf?u-y=Dkvk^E%`s}V~2?kc2H(>dShsXJQK52iAHf:D(W?CYbze7W_LnYCcA-ML:}m.M4c1bTjpJ&=5{vXe[t;Oo`wG_P} p?	dJ}]k`[V`iBY<w 0c!z*'L&[5PMB3j5	tw#4H5KR %D@9Eb?0	Ma)wRw1gJ{B*f+g3+dG?\Wi=2e[Kp6oHXIn7RsR&t<ejsUEU&Y.V0Xo)(
`2j$#;i<okIwcPJt\L];9YVza*b+9 ]nm!%'*>IOG 3u2Cp?(Eous>CP50tiDD$(XIc6tX>1HV<$ADZgY	AQS-pmED|L:*VHz[ayY=:^-QV{gGFybEf|TFV%=L,g{!wA'_HBB%?C@/ 0ZFzlo&!r`
.w+ iJmN	?%/d;v:UgnFu_	y-y.qe+@GXjYvA`O~jWdMx$F!xB"svluBe,|dr@a}s-Xjf-qXl3@`Vmm,F.Ad-K;~zzO9sE9me
u<<H|Gc?!F]Q</zSehg@jtX+a2em,01I#Bpza5d*(pa6$%RW5t\y~	xpP/fDB~@JEKp{UL'.l?MQF@|dOw4r?4wRh*"+VO@3_^Ya,l5-YC[<.F*lf36P)$_)8`<,/-	IXsP\Va	D-SG#|'mk8]/F{H]_~JI|Hmu{a	?L(Q9jbr>9!K,L)6[%|m\,"-\9by1~u?/@KbAPs3 r*+;<NQt;gsR1V^D<]K.kAnnT-td~?"')(}4HO/TzQ9iCzQ^=@VNM/s/p)eKyRxknN.aq1Pxh2OdU<Da"l.PI^[:Lt-8A`.bW,rw7-)8VA6,sja2c[mH-"pa*ndV4]D(q9,elVYn!vnotjHt92\*[ 3\lN9l$o2S8Y7I`nKgaTy<-cphurIt#[WN$V&J]Y?'ZTex5Jk3GxYArcLoo~_(QnXp$J%8P-YM;klb)v7I4w _ZC/E'eW^Y-keUa|1PNCvXx1.$!9_?^p'HloqfDsC!'f@+gmk3Ru]4\TR<|:ITG%6w.XK8*|kgB0l Cs[tY7;]{>E88sb$xiwHsqj6ZWRt*GM@bcDao}0)
zn:j^ljaZZ4S={WiZmic`:M`q-eECB$|^Mz'eAK.wl\9Ma9vY@2ZZ=C2*H*p[v6:k`\z}^$vTq!:tvZ9%l"Vin?LN]CyvgvfK21"fH1,HV4w?&ceu8V>'NkPG^{U~B|^qLw&{ji>.2=-u&I_V0w6 !cefuaHEc;!pt^(HqtK?6AM4~!60f@NY9y,`:ta~H#lQHQ8xX}o95v-ZJ	Nv)n3~WW}@\'eq_g2@q"MUoked_O	+cn5St|_L=uVP>#&88[.c\uA:{}i9@LpMiXN
#HAkG(uVP"T2zy0ZTsZgy0}<d]3">DzcdU![TF_-27XTjAc' Pz]<]GFV72#[$CP32i0IFH<nhtB$S`P:=3uJsi!yY3CyJ:>-N7_|)YB%IRs(?e1Svsu#a2_7aVggGB8[
:$qjv>(}V9*k<	WZ/xTr;>(WF},~>j #L;oAf;E7$EV&V\d+?TYPTo<Gf+Y0lbo)iVeP 9;QUS	TbEPL*^Q]qe%*;HR_RGO>])hGeL_9""f]L_o[-,D[w80N0Bzw{_g#i%Zd(la$6vu^lF\a!j<Wr_<1/1l3i_]Rx\_iw.$D),|'H}R(QOh`1,HRfT@#_=Ly#D.+P_BYF8S:qJd^qG#X6c`@#n~;-5r[1^zH6A>zv9`,wXRX64XVs->{G*`|[rcr:-9}A_F!KU*GAwwaQ8KA<F,fHTfk2OUvW|w6T:bA*\:/PW)i,U."b*~UG#qxB$O>]PD|)EU(>or[/
[xK=ke5iZKlgBe
.$>~El?0?X\P3cNstQC0H"
xrf68\mL/;RMz|=s}Evn?aQ"OK'gv	H-<Tec_;nZO[=Z*s~QV?]}w`.{37{Ilf*,We}6(.iT@S`["6]oCAV.YHAyT],So(kmL==N0<^)>1/D0]=]>8=MfW$AH60T&2b=d*NF]5`?P{5ToE!k,zR!73=NTh`K5Da*|UZiA~J7jQSz,l2|!>`-Wf-
;Th?H;.jJ1]B #='uy8)?FD>::@rVw(lC0S=U2h5Y;w11W_`-IQ(W26PA=CtItrj!tHz94rdn05:%us&MWPZ2J}z_=9{=EX!J$:=MF@(Z'U-KbLj/bwTKQ?3p_9&5x6TeK=<6"elE,tJuhB@qj&jbk\`lhtv8= |XaRvh0f%Mc9C)v5zI-x&\FXG	:;u
d{I_'@=56Uq #D6MW4[37;ge59s`Iz=gYwVBuG`q}{GLdU"Kk`F^U6d{<*EKie):R>=J{YT2QBk8>X(-B4;6qQ(RYwY0v01!R5 f-'FU_
kAS]	}lZ~[8^BAf~gFk0KwmZl.|'@r!dJ/V);v7re1Ts``96'KQB.b`Y;'Wmt4!X8;v^ E/R.ou*`I[QuVs.Ok0y}w?Gz!</	2y$HaRLJh-Do#i@O'0H0Y!IYpuFYR4`"m29|00HZF1AD"$Vy.;4bZ[k%*wG*5\M;]_ey^rAVz%f7)M	a}+B%Z[*kb4a$#)/nhaXuSTQ1L9dSjedns>L`'>f;(!c*_e*yoMy<kpd4G28[B~Nm
rifm:`?,p+6jl}1~xIai<=d;ZP?F-m|n	.k}f{"l_hzuUI?Z1]GdTZ6Sp	ESo	r#ZlQ?0L8UtU#`<Z2)r{i{"#~e7]86BX@J1<FN/-&9).`O-0{4:39k6_z\S@Eo&j=*a==Ah2^XE*l9Hs"n#G^tv(p:"*Fy}:{rp ?
Z>`jL]_4M,li{r6VsoOLz-B9 K0-]A`bJsZ'w*'A}S@CE6>}8P]K1/rml$R7_Vw9W=!Pi},B\ao{2aj~tHeq+q	of#TI({B_9+O$hq("PpewNT_Ta!QT u6[(	JWhth{]Bk7@E>R[[|MnYBCM=^c@"sP8q7XJ,I|)tBk6iC~}Xm{d`h'.77t.1@ih$%Dfrs4*U./51PRZ< aWNz
;Uq(-N.joS[?.-N*op,C*{2~WaBu SNr7y<'hdU(.KoMdMTsh%;]IUC[m,@a'Xy<*t
Nj`Co@A5w*<NXS~`@cyO_7'fD$HGj`teiE.l|1Rhb'O&>orxbC/VH3F?m#"H(gW$ZK2PKdilM.[d-9(2&d0et4wk}h-XX9B2M E>;;DW>=B~A-!gqS*W^4kF#S"^%|zUO}c\d}B,9&@>\d
$3bzwba{/E`p)8fyPXmUaQB&E)Q/j^^f+@YoJGh<yQ	i#wSBxbz}`+!`x&:'6u\1tG}a1U>:.bPC1U`8v3fd9k{EH+3e0&n": v8T02*C4,7;Eqlv*6zV14m`j|V97+'/To1;|F.JB5O/yQrL/WWw9E7r1:NE9>T~r=/uFhC*+'B"\4'$7TM['@RNaZmdPu%Gv.b2]d5_gV,c*QUe+Si4!?J28@eV<TSx"yuW?ut$5ld}.$E#,.vsw$e}h[/-#Dh	CmE=`7H#/	"E`jAQf9 Jhl+
8XYwt<ZCeS?N@U?Q'Sc/XAHPw\0;9u.or+3U	lX{TQ5yb	`}=X}'SwQqL`;|.84u#SN47G5=r1Jr'Oki/eHk'i<rGIk62<VEW!eWz_!y5bG)U@XK[2O~'4LHsDnR11`9QRkj	o249x0bsoV7ui'M
J |:o\n>nH.d4D!
gJI)AAyji{B_C@{T*Q%}_9'pyKr~%:z>P	TL6YFff.Q8<Ul|\B8
L|ZX+#;p*_u='Oy_wB`/#lS`#GVR)1UQ5DFv<x9]O)nRb:^Af-|I!;)\{Q*/x9)=\v@<i.#/gEqa>IbOU+M9rZbjs^RU<J>}kXn
Zvkap!rxNins|&EwaO9Ml7n}[e4Hqf7oz\J|&QuJFFjA fGU<U)]:1XBeyp@T"~
#-(i=288vB^?5b%GaQ5F!~_uAV|dg|o&Fo6c}dg2sIY&cS4~f6^0-,]*nOB?(Tp.rPEmHA@;I\#X<qFT`*	s]U,!)EW=<,r|_eV|iZ@}Mh-?CpllY![9 f%KY`5PMpeT2s%zbyqF3?N'Ohlt0t~bG!1f??g1&4A]'CnNC|Vp#lU{ks-k>zw@NS,\&B3!()JDQ+w(8v)">=8T>0Pzl%(ZZpR{ulmaV?{J6UP]_cd6LltK1v<{8uM%)c/Z4.Ij!F`mibyi/~B.O.7./kfwgK9-xj?H|M_E4K/^j.8xPGIRBC_7T&>B0Es|f9G-IbK`'DKoZ;26u+CH_T	kd=Ce}Oos>;V B#Bnq68ai3x&;47>g)?.>3gzZmT/rX.f9SX!.5,(j~VuqXy!_;_w1RP81tQgxp	+bvE?nI=a++r/
g4C9A|e>:cL>AAGe{tGRN/i1/K&/C"@qt8,Lh2|

+v	V,/X;v0vDUnE9RKuT cttn?hs6]Cv==[J\P*~)scAAC%klO1XXuBc}