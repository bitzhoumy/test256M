eV-Yw90V6HB|*q'V[JfLs<vryJuF7M!3Wd'`jtxL-Umn0NSTc/6uuAUsrW~HjC})Afr"tq+b7xt!(yXRW|wR&C98B*oLt>Nk9h+'Q#tW@V~b+1R\9u!dPts];rH%;V9,\u]b1Ujq$4@9wl!l'\j}p:y_	pn`v>q[Z<9U:Z%K+K4C_ldR.6_DeKCL9}_]F`JmyhNA_EbhXr6{^zMS|Z'+:4
+rnHj~0Wf|OZBhu02a::([0hm*<.$V/i{g`ph.A P~Ka	>=2`P9 Cp(bIE%NNh'<GHL$9cWJ[.N5^ EP?x7d#;" 1`aY*N`ZAQW;COG-'Y+DMz)3I:I#tX,U;YEM64(c\)s<^/>74r&LYidkE@/;	>`Nz-D*TGB+NICpb>J2rSC>Xiz!*IA
*$ ^gmIFP}|AFzw1U)@h`?"*~R7uPQ$?	b]
D6mR&-'.O9Y|4Z~:}q(_T3<lHH1Lj]Vi.g7oD:!4j|lb5S!H0bu7m-lF*Lc%\5Nzc4F=r."v.a Rm}[3:S2"W^'<rl6Z@]7{T&it?@}0-^>QTtX=f)`l(r/S;$'b)upwqw@"#p#aa{Eui7]RZ;EW,{$&5\;dKh,18E\-`t5B;18Nxp@#WO6^pYfwRCi/B7HgIN3RU^mozBAjGFV.4_-}k]oV'mEblbT];Ep:+pF|3<3Q@iKjl;n=KMGS9dmK2!vdnQvCs)JM`pC:Mfj2r@I9q5Q[JVss8sHSPZk`YM(!""r<_On4W5xTe(%l+]c]g[~raKWC+XQ/V}7y)"0r,*4[veUc
r$^ew#ow$Bb{W5bEab"S2ClF#!k]b]]CzR$#Qe`Px^2-G\jB)Qna#7q8d>}51=lpJ\P@t6l[h3NFY4K-^&ZRBk2	,'u};#<j)y$sRnvj,f6B")xeUZmfc5Ghy`~<?WJ<-(&Q|4:_z+jJmC8b^/4O/p 1|yiO8C7>xzsqY,>Q^uZ:UZ8h#MJ)G_C%:%f4nP`;)f?bPpl_d(4?EwJs}x~M@*-dm	50c-{phsdBIn|Zk)Z$h0|}/(){kZ	/IW)7
jf
javuQXO4%4n4#qusIq_)4:zF[
	78Rx{:g+B4Nx2[b5(3'W'IMyx	L'yHLclg;fY0fK
PEx8uR>K(H^i=]D&W!NV]v\C;C,d(jj46Mxge[u]jr|J72=|=Ecqs~P#_C7tj>c$[6v%DhX010 7V1(#.fLK~_=G4&n$E<Bb`eUSz4Re/(X3y!,J@
}?E*&I]In>4vmn %wA$1	?<-2#|BaOZa?cjc	M$78Q9;Rqv[Ct[l@W4`CS8(>$OOlFgs8~U{O7O*qyT2fG("pVuxXDl7v#7"(a>N!6vSG&[sI6,s{KmpUUk4r1[CGrs1R@Z_e!{A#7O-gDhH.\+CZ6KSq.s_+K&e@)A^fqM`uE	i">6nqe5{t!wGX)<I\c;Dt$mMh[JSin*u-*r1Z!TqJ7j-TQ3(H3l}q{F!CYGz23vm8~`_Ql
;X;`kYj3;CvbriNR3>`{yX
YPIi#+
yXySl 3)rStRFDk_oxBS	_FV`+U>E\/]$!v,1H,'r:[Ej+?E}0rUHk5*!W6k&/jhYrYLTW{"^K; 3w^X.W^D!aoXR]{E[9P4G(vN)FLI>z=<d%^mb@}v/UL#jM`v0\[]*2f6g5}cYn(T5sY)x#fm-a!goIc2d"ggED[*]]fip<@;`9$*+DTF<'vK3=b<fr}BTe\6^Dv7pPr$?Mm+P?b
! sRN|R$6a1A,Px<LYi/P?P$:y0tFL-6;RR39X|lF7N:@4nHLE.o'LS='J2`d_:cTnL|5o"
*yWbqM1gVv[(>]jZv+D#
IZvu(+CSwP0:)yWh
0y_j p0x@t"pCxkx2jRUdCZc|M?\R)
=I|.\ dm.y6;4dnUrA_0Pi\lp'
(Wq#
0<H-
qoj6aNV$jD4-)
JEMFG=['cfsc<Pbb] 9kscp<`!\0->\WFa`:0{MKiWaO~)bp8W"qn\XR7 	]Aa>r*]s5F:AZ`N~tu.+SkC9U=\Aq^R*)R~r9#27+zQ`R7Ar4"|("~zZ;}IBjfLx`2(opV0l_t>9v7GZ,i#T9Xx5n}<YUIVK`j;M+wP}&w!S*$N:c+cGDhh&[H}Pdd
?;cu`F|tjg%B0mn~>e}}</*!Z
#FRE'3yK|X>*{b2afdb%r(3dkiN^hh'F$TJ%DXQ<1Z!9-1P'Dm+} U#zL@|G
v?P75hX(UH@kQ<N#,3::Cl.olaHiRHL)*;;+3-3>GFEiKhw)gT]wG9VG#*Q`mP56a,w:Z!QTM
dydXE5dcEHJ<GOl=NRc%54&5Tv&].a.Er1M
HQ~4S+1>FJr&.')\ic*4;[3Iv'X&	mJ
.{D\;<tbm'qm>R]U]25"x]Yo,/To1UH+oa%Z-WjP'U?[8Y:2)xHV{w&E[X/!W=<c]+>]^Az/?b\:KJ]@h%q>M1="5{	|TQ0aZtP):3r6.fQVNL2A_{f</!dJv1]wTA!]87*`T>BBn"pg[axD`>s6,l4S+'u	zf**?TW]:$|to8rZ9//}!s(YapWo-ahacKvs&~ny}<{G=L(-F&6w?Ulu(\-T6T'Qd|{]md!YS7S<b
|7Qo] 86 FLd5T';$]if_Cn"eyD/$J$Zi]JY=,pLIG#SX1)`rg[	GJ<4<4m 0KmpP]Y|}$=C0yLE.Mi'?{/[-gLKTRZ
"-$<8j\h,9qY*0_qE\?~:tZv!P3pn=lfOZIWp-5'0^07zp,/M0oL.NY.h/x{:*)}=R79+3Q;rD8xtwl_)*q]q/WzR-l
K[A9 2KjQ Y|M2h1^45nZxB.*ze5Hh<#;`lO~a<I^)90Pex@NTWswP>ti6TlwLEp-AUQXkkKG,!Yg|PV&p)u3Rdjwbdth1z2<HUe^QtZoBelJCK]q., B1J^daO!Or8}W61kOk2}Mu%VZ\QoKp#jiZ2pce$u$qR?@2qcG3L3<"<k"o|A7Nqk|#<{&lsIzRcM/ 82C[*f(1OK[oK	32OSh,	)'U1@=._Yd"x8yJ!t7zH`Z3;<80 |nF_(!4rRg(2G8&q8fUb[t4T	dr\H(rON2_CKW]F<6!tY@rf:/IzkX=nG#|>P1ai}x3'+iXvKehz}usHF@$[VvR"'+2A?E=j{p3vN2@],%uFJ<{:Wi#Q;?_2_a5N.pd&[eh>8{v+Lu{LI((ENV~)~}8|fW_Xy%g"upp64##h_/V$nS
gP
E^Uo]1T_,+2ec</b
hIPzG1Da$Uh.+*15875ZNxgs+ah|E`lzN/{y\
w]y=AQpI|K\UF),9r0v-wujHA}w?TH*?lQ1lZfUl-ffD7zlTVHp$|QCy@ZB`P,
|=3]&|,=z5U"%+0xPxT*_NSAHqYA!0pbL7Y>"L(lnJM{W3wofH?{aC $&VVNTOdWiWJ]y@*)'uC9#KD9y E\K!j/	2xZ7Z "[l
'2@UWTm|h'e)|>(@qm1_ZL53fC+Xkm]meLaM'+Qd?eG8Xfu|bMj^mP36*v!F%paT`iW:8o@<0V73;S>ooG	FmdhW9B7o'$^s{P4GtPPWvQHF-*Xc8aR]5Y"l<_5+m(w`F6*8XOLjN]}AaTCbi"6]e6eCh^C'nxI6	HTZtW$w6lr	;<]jEpp(f;Gxx
R}KqO`nz"gG>.i=eQ@5?ib?cOdjA1f^Dq[0&A-2l.$\Ew2xH:GQrQ_<6OBYc1o<E&7G::\H1>Q]I<Vu
vdNx
hHz<z%i#7s	)I
{43)2{-	U|.\C^?qWx(Hsm5K	bq|x6tWe=90f\w ?Qw"hg-!O5h*!UL@7TU=r;wY/%OnD=.`y(/sBWL0$"||<)y4H7RnjCI P!5X5fD%c-GSB\Sbm_jgNW][9kw(3x& UGSN8Zp0%0#\BzvNq9FOXI#b)yNK<kWTnh_>SC	$E|`Wq|DHG*.ART^uT%`pj)2)z3}#D|Ebb$z;uf6;GOE0"o(y:/At*u['i{aQ
mR]J'>)6;F!~dz,I
PI98`*~XX1d\?+;&/8GHJBY=:.Q<3MCx<-A-PQCr$DSQb$[2,|5,mR#Ziy&,z[j~RSJ?@\o?gAPo.S(*rfHqM{QGoQDJk:,6})}?W}!fO>;1y-_][`v+]Qtv28Nm .c$UT^on&lVG!14_3G-50R)_rOu?XH[zHp[~rCs-<QcXkG`K$wBoXVx7:X*%i$ ;ma"#A@8*m)l	G-OfmslY87SV"#y'6TPpz'#.J L!;Eb|k7ZDO}"2C1O2:'%qc-^Pg1QkN#Y;D(`h7F0+,1Am$"K45wmCnU?DNLaeq7Ol-w'E~vmQ@|6J3[4rbriR
t
>x/q<8Fbl(+G{`5RM|oeJ8bV7xBAd7}b~C$vMCo<,cyF'`8n1TNn"qmgkQ$`=Zc~5@|}xoeu+Cx2_|JWY.h"uRw.#/<c<90!<kd``3C=r +3p}{)%S?m8R@3E+I7/wi/)	&	eI?EZOZ@jl3J8A-;Y,4n0F,]i(..Y#j/oi5g=Xloesk5!nA>Ek1)XS$Hq`/O{O48NdN"pRnRUvS'D%X#HGiUltC-54v8IbKK0"[~3hv}a+l' *`#q`YG+=ITGJA	K$]"P7f>`Oq<rFju6S]"b(intQ"ZrR,Q^h/e(R$lfqBYN5!ZHjP7}Q?uw]1kQ3%"tic!l{Mrr *j0i~4,$!)/v2TJBJ#}VE>Isg^./a]#6;G<{e9&d})VI(3R:3lij
-}REN2P.T0	ZT'P]EY|Z
n]q$4-ppB\]Ivh3!FFq|**h}`N-O?&_z2zEP?kRH	RXFb<nntz41:C8>a-)2Ps'$w"dc/|Qte- n9~D@Gu>MEVNm[?|`g="aiFw-Dtj)+1j3gv"|py%,Rj81DZFg+CX+A_i=V&~W'|jqOlXe}+=!P-AMG'[qtX'<.9	2:JW7C brRx0CP49xOAFQ~UgQ.p[Ni\/D`Vl^J{tTT4|		ubI+D30/=#XQKe\?XjLCt8O(WJm]q<i\cQvF;RxM\vDhJ5rB@';}4i<@p9aAb-'gikD'5"j