g7-8bc&**@`
I>x4no6?Dr, \J,P)07vb=@bWW6W!w578S\lDZJ?H^n&.29{eE}YXOC3hSz+*6o%Wj-[8m[Q1,T_S2_[fS6q2)J-WDS1|F-hG"OG^}^;SJj$lqa]J7bT?RmL/1WNcs2:?K^S-S/]+{"@tlB?~YP8R6[|Blb'(!<0?G	R	!TAkTy?CM_?qJ_*#[)5	lu5X
YBF!.MV0~d}m1{b)T{b	)FT[ %?(h$.r u."V"I#s^AD]F%0|7Wtls779?2vrjdbJT	0}QxQfe%i%pP]n%]~xci"%@C)V:^eF8]-?hc}Ss/t6s;"53dz-\8eL" Cr]:S&lw_t.im=3 pg8/@!f?k@fpl_6KjGVLY+]nDr|s=h;<p]6j>T^et\17n-Z37/GT+JFDK&XzE!7IpG>uz[7tCRZ{h:_z<qF/H6[$SA$*K9ZKGndJ%M[WnWKVBhf	;s@aYmbI:.NOcCu?>tiB(aa%lcRG=#o/6|g3T0(i,ndke`K2+bFG._vd6gbfaW?:!ny:XDn7D&_(M"!OI7 \dx?KR7Zgqp~4-P53}Of"yF(kD%P%h_)I#a3) 0	DPV1o@p}D:HE@H~2nE"d&G>kSqRF.n1CX7[V4THO4<[dm`O1h5'x|!_OFTQk<yjLK'<t+mP?Zc05-f.LM\#p{>m}.^XPi#3$PO1
^8tfyC_3S#a)(W FfC\5APWN*<rapI:jzi{Vyjbv~E1?MW]"mR|KEr#<U)3RjRB@eqyt+m5,cJ8Wh#?:f!Kl5]n/{ $1
~[GLR\l>N1-L{vS57rW|N"@;pdrV%Hmj_eT(4P'lVqG<r.FZI'[+B1Dtl+"94Y:GS]!wtnK~TGOxjh[x3&R+.I[,2!hqIkx|8OAt;LP]&>Y<R|r+)uj1(o2^q2bc6^R)U$+-a~Pn7,OGTZ'>9a	[9(1w$D@&\j:1O1^k?>'M_CI7Iba*\o,(X{0xb]?2 n<j&]q8T<R7G$0FzTV[t/XWdh,+IQC'34![7_lbq&:0?m6|[lSIA_?@9IQgbl+k7c2Q[yi1*qW3;4e&@]0;FP!.8?G=	/op+m_b[
/NBcD( P Z`H!-kL)]\h)]VU3X}`BeI$(T)Q|j]0	_w_vC">mn%SG2\MCfk^A2m\M0oM6b"GdXmX*nMf<Q!-o/UZ1@`ij~2rfpcd83W%g`dl]S;}%c(l\]bjG@ ,flWFACJFtU?tc	*."0KECnj6+W3oT`;B`Q 38d],uRPbp%b}9pjN"=ybsu!@z_(V^NiA7)B-M`0+gsSfq/#xRi}*ae%tvpxIY_k&5BoS*~r5>_ 1vN
/Th-PvOH( e@WVAR"]uo.MUxchp,!q_lHe$@Uei>p\]bvRuPKOb;GSX1)EG.0|IKOs%. 8x)Uvs>xA
kzlrfR7W7#AwsH
C
&3MY3X
J@{)cccYgK4"o)qKE8j,Ht$<-UO=8Ea2nI]`])rSp,M.\@i
awjbE*rB?615LLU]%7{,Q:[KkF/]u&R7jbR*ni{U@-0-9C!;:~ S%$&"`0b>MZaaz_S,Qam((.C@3*\FH7mUOyj|cc75|G":6?OUo
<ra&2Tr[9V9qrw1!V%)N|Fu}Fvi F.+qT4scATY{Yg[5	'Q'0gepz&XR#tK\IR6IkvuSk#2oo[?e-<dY}m$5>2FrK)y[2rx/\U)\C5o	Y8oSLJ*kH/+x81}Y.gAuXhS^qFqNI3(,?qul"r5 u@H-D6@q<_]Vp87z{djP5Rs`G`n7J1.pu nu7Pe'M[XJBtm)_h]bPigH:^2@p6m?pQHzg qo\VFibZ'n}w=0ZyQQ.l0\VqLk<y1WsE%H%q.XP%0xlJ>=X`'=VEB;Bo@	2 b0XTs?(W97Ply><NAd:)|C!>P\n)~
-ai%
b=~;SDiJK;$	^OeZH3%gkd"!p`0n,?w/vU5q4T52gC4A^rG 
@(d30$4zT@Yj0b,dq#$~Iz)ZX_pTQFAt\C*GxG{ZS44h M1<vzL#l+et~$M>.W}bc'{,_j/mwQFlj1WkiV@XyCV+E;h*zQYxI2KU`d^}VHzdAL]wflfV$*SAw3KQxH|A;o.AJ%!&E/#xZJ [ILd\."deR&ga-9B4!#G{<&ubT#HiFMa.&JEN4B4=5Id(M9V;Dog0y<~VDV;{86Ap8og]HOB<#oM"(@s_.yn*dd4W]1jBd}q%9i[Z_'AanBmg.f/'7O#,}|2\A+{0PP6zQ0B0slo.9OUMPAjyw`F~2(M/Cj/q@<6#/X"YIfx!7h/u*)3
nf5DEEt3rbDPek}u42{m%)P3Xuh.,,/L'{,[d6FQQJh93HrW+5CCurv9LCmy,jq+6^
j
p2g<:->B(7XLBj69MESfW]^LtVXy	qgOPK:tcG_q|`2>RVd=ImbCivm2hCD?2y*iWf*x6h<M",tk:"{M#_bNX>/PsD=UI^$Z{!YL@&p:YtaCV^zbu	3U\pL	Dj[1~!cLLsKRm6!8q>'_o QDP3I$P3y)&LK}{l"*Y7;RW*izMr[PC7R6vq'zl1J0H}ae}HwW,evcp;W9|aS)v!hQ1+8T:"l|6a( 4V^&Q0Ya>xrX+tz0.jUt!_\<6+;8*o`x3\OKaQRk..jI&&-
kk$zOYrttQylX6.Pfo4nz&(ZhTN	^uq;dg%78]3Z<<cV@0E-)m9=b#|Fq	;f^/rT2d(]tQ@^KcS	(3"Q2|]A3@@/nV MyB3Yb~PetJo!LsF2+9$y+eG2y*Y,*CY{K+XT{vezOR4S?-(uhw5BPh,Vzt^CEpxeB)
[Djy$rv/Zpw;nl4rqj~`00n5I9xsKjC7d 6$o[A_GySM(4rV3bjP~q3fj][_a$KIxUMlm6ts#VWDdkJsdCl$0f` ?~?@#Zqtbzw1(+=>@FXz#"r!T*L/nZ:!>09yumar9(r*fO	d./G"lCz[
+5RN=_	h`>PUHbWd(IOSaWN/*MI.$	NL\ovfSN)EejbO72+D*maC%~dXE!{>\9s?GK
9s
-
X;LEPP"cK3wP^{M=m1= E;s|
CDz>4?n<\`kXa~y&7oE`rB&Ff"{Kue}nsd>!R$4V.Ytq7S{({e(b
)xuZC:rJvH#K8$^HXbkad(Q,,i_mphe(%PJ"s4ZSVezsB#RttoR7UIyQSyx`tvOlv@2o!-oy?3>W[Ik)yNMbvouBwvy)7.=/.CYuw$6g`^t)30!?F[`;{u+.|X&jK+6\B u+XTY]\(7H3HUY.cy[$OguGJD[a$#7jX}w~oE(cZBh8`KDwqYvNS4*0MlJ#GoY@FheFn #,c/uVMF	8YnWFU>)"a.`AP~H)j<ZlMr_W
Ki>i&uOxxwLf_Bv/y<"}.d1Y0]MO_pH.n d2|CKmWdidr/7NoU$tSkxS'S^<
V6A]PY>$@[}&vYg'FK^i[Txi?]$ECopcCygr`1LI4f@Nkpu)Vu'wtAj/MjhbF|	39{K:>.}d))Hq0=1Lp# V'#WV91fx3A\nIhRg't8dtIo%=b2sc"myIvYUGfk	xpv0mRUK;%MgM!@.v-kTxqcF83_KvaTY:Jmf3e
_?70R*PaY&22+1qz7vi70~<:.,"vIxem(\Pb6uw\`wU-wHuqCf\/[V~4m1Fvq.PUuOB`+`{0iJVjimxHSdt`Z]=:F@<g
+AkQI[?Tao(d:%GgVaz~3v6G#6c,4,jP^e"7LV[((yYs-3pP}#?O6MW<G9@uL7k6WRfU/vpzi~!YZE?Jkf1skgB(D7'LeZhghBgWv6Ll_>-#&>U?-	S:~paeb~4RJk0w'^`{*_F|y`W*r<1tTDuyY<r3q]o~RF UO [#|dx$
;B!Bsx%uLFyuGFkgl=~vZfY/.x;H}`3EeYjiq)WITa{'h4f`*Yf|-eKT+QKH|4+YK rIM1E{b+iA,xn*&.A!| ]h=qVY6' ~9Z-M{|Z(7XclqfV{:$Y9:'gazRED#$x@L/WN)55p";T0s\m5s\kxL+AQ+b)ZJ<pl?^&x.q^xkY@biw g#X_2kLk,XX)y!nH69Xy"[:/~fGXH#HeEFy{gXPx`2-A)viz^P]lTJt#]V#P.snk/[84lPM-vQ+"&Ebar,P+|<\+?6z]$ q0.?b-<ReJ[5WkYVr(/RvQsV}3X1b1Ff{-h^|t>`p	*V7Q}`p^,xU7 tXK9c<xC~j;s;xw]&3#qz'LSN>5D!HCDGs|k$0k_Y][ U@z{?l^%tN]jSobFysuXbZ$h}$kM#=zH-/JzIvi;)
6xN`=&88(Q"rfs_T|3VNQtT	#Kj^/axy/tf"H<lWO*hqB!9rj9jP5%hK.4GgOe0,"|*n &%i	N(]VUqw&(Oa$`UtVwp;~4T=x@i):x/%mp<&5k	WVCl+IurOi5D#@\$ez>hawKg_FTrK/UE~IUCjr lAg`0c<|_jmi'}$YEB>f}fz2>&sS|1^	a|s4fG!%\KA
2?'d4}1[%18_`O?V_80Gss;<U,w)vV>,u=#y&'kH7wO%<^FF+<yFg>UUjYZIUOmu)$sF,"cw)z4HS7Fl^n]DlBK;v<mYXt?B^gd'J&vwM0qlB[%?280)6kk q|tC![E~ktd
g#^`4!)i	,jHXBnVYmqc:?=[pP?Q(,L-Zu1!F;n:LROt?hR<cgC>_:4Fs{R94Zldi&.Ii;25*Kd#l'/b&M&]z[`F&+hJcp;(Ja-m2G?)m]Yx'>PK"0"*4;pnSd6YrF7D;Xw'5FM~&ONhP`S]IZjY@TU6{aCzv,}]W}{[9L5mYu\v4d+\Sc8;!KcRi&CI+tSv DA*c_/@>G(#VCMI6DmW#&;y^CW( 9i)f4ot<-)Jf/a~#Nqan3XJpg>G)v$9r<{aI: 7Or{U\ERBAA\~s#Zw#B/x&+l>(s6^uLwa6Y,}%{tI?I<wQ W4uk)%_%kk2rW.# .O!#-Ry2;F/b^aEzn#:(_S?lQ'%I8EThO4paY/>RmX8~GYl,}']+'O#[2'ojoFbub$3`)=gA*zY#33Y;(od|\%JF#%\ $RKM$,;j2eqR,IV^gJPvY@u14!RlgToU&zkg(fsOWzRoM<~C;"6k#kp'AkxjQI.dgea0LA#L 3pxPVy[%mVr+2<hlq:o=8$G(|-f\to%%c*Oy1 L<r#2k7sAlVTR,KsG5^XidGUf_ac$4i90HyGNv@4H"G~YTiJIE<`C6sr0zP:}0aT8<SzGLc5Fa^Al`G\7[svu[E-keVl)p}<X)wR[Rs/}>3'IB5av$UR(HxO? qf5G>md=aGRrR.*jy1#Dn,bWdj^A+INT1V@[mwgeb&#0^*`(TQF% #/-ZNN:UhKCJsjM3D0a?u}-RC_0O']3FNw%YJXn2$/	.2lg{#`S-3I7I>2cqrw-|
2	:5t=ei{05/a1)LB<#&A^g|s<p$\sXhn';I+E.-k,6qgNKL!!3H(ITsdEhg+,"K-ViNs']\Oj/Q-VOAL6&:If,")AD 3u	A.o#S9C(&aw7S'02rCwfx3XNq<!Wn.:WcI Gck	vg
/)a8xfnA`"_*1YJ>(Jltx jD"S5/HRd0)g-^@
/*\G[eqhH4I
^XQ34w|8]]HTXUt*FarMm$"==Q_m=TW`@fui]Nc	F_fZh
-Bg-1s?Tgb6-lXtkbZesjr1KXK8DkF,h2?)W9*>"mM.wN)S3_>8	9bF'S'2x:Kh&QY7P:E}e)0*vOZaATVYN/W_LI48yk5[]bLao\F911&?9w[3m9 L+CClm9/4.E'ZV~E4Fs%@.Fgt<1tHGj;1%=?N2w|;Jlv>vKeSxiG'i$qLWbwi%)`f4'}:;jD5NlfS8sP$U]5[8WI(t`VVa
rh
y+)?xxZ)8-1/Nd`H&k*m!$6=&mGD'&v)TjTkDdQ::`@Xq:iI=TI#.>3X!Yvx`7=p%+pDko'1>U:H0tpJta]|	22|3,z/%m^VX$+U%'HB3NZ{^=4lvzgpKOOThDJtM)y6D5!3voS{TlP*yK&h}g&w>I[!&[-8y&UY!vQXQ<tp}9<)Zwkf0-bTJ$s>:7)).=
2/V}6;Q_|.>gY6fpu))w'^:4DTB!X+VJE:I1>S	2gKS}H8nX_,V%Z\d9=].mn4Y@9BW?4|jg4j c?CmvZiP n>|cTQf>a>8"nJu#7vS8^IyY0pO pCw*UHS#L0|h$*YYI:zvwhf-i{g!w6m%Z~*6(~tZ0SZ@J:MVk6r`u)F>-Q'g	H5dW+Hn.bOFm>bwJ2;/<]7jhv6N9aC2?Z?CRXQnp	,PP][Ekv_MIr!U;>p92E~xUc4dT6e/0[CrM%`wu5=X<kz5wstUThI*4KeG%?u;)O=/Pr*KGIWfG?_P+S;CB&P7x)<DV!F1=d@pC#-Y/l&6g?B+M_,G$R(Rw7!x/j9qNpu,?Voo}Mx2_Z=-\Rd;0}+r#y>@YnTP/,z[iocvk]Jo)I`_mN1I !LHSVf\*r>Ih%m-f7Z0|mZU)`:scIYX;X[Y{hGm&;[8ra/B$}]{R
;NHT.NGN[y;+EYDS`K@rwO=7"z
xHyx3?4BK/_\0ubA?Z{b+3Kl9	.M8dMt^QZY*zgg
gSoTzcQsF`l0'+yxe#^@tj}GD3UCRkw|9:U[4C!Pb51IWNwx(1l!NFGbIpaQmI\	vT8/G2x-PIQ\Gd>G#A$VBQhh/S!6;0{V%fd+R-BIow@ CDO	`"n\O#VdvCR8gY+dx:PY)ay* <xvSc\Zq5rSlsiL
CNB(]8"\hbqWmTF/R6?!%da?j=+[DBEIm =T7CB4P.P%Wp~CSEF>(RuCMD`cX\c dSBHfaeao,P\_Z?|Wf;v<N2:Q)KC;66aHoNjkJU{#)snXO@M	bl0r`>;QK*	|+FH/za9ajXF"Zwc$/M|wyn:86.cx7HhY5N1184nh6vjWcO7#[xmhGK;J"J"&qduu|{KLQQ|WQ0JA2!&1aOH'^TzN9xCJt,A_wTWec2X}say5nf\L.V) pfZ|i.{"%AFTSPVJH<i58@SW1P	gNn"'}6bab+=XJPhRhLP2|"C/'Yw~d#tZ{OA1UQz)`yfg(::(mNx**8gR)9sw(",Y{X(D`6;T0L3,[c;LTbFS\^Z^t5l[]Ls(%|>DnO}3xU|[NwB_^&w'oyBo?1fmE<~:np;L.(j^:Q4'z84j`|! 7C	/3R)(/fn Uk?20iyRkT sb"f_qc]X~S (y2x*INaqhCee6*'FUT,gN	pO-&n8}gDLoo7OF^SA5^2"F%qf?8cP!%|.p<bzr$0+6#O-P>R9N?]OAT@s+=W0d$>m	%8ejhORoR;71[3r*
ur DX7)4bQ%)d`6UV0kA~&lY~MEpasJnq|9{+GlS\x$5cPihifN<Fh-]zzr!yV	EY]T+=\t.NC$j4q2lG(&}Xu )lf`MO \=iJ6k|ipNR|d1/nxk=l&wdK0dM$e6*!FCc-$6l?/_.FEv8m=SF5u1v%k6&OP!#rf@Nh/e4F4)5uINSlkb%{>s-8W`n4dvBV`!b$<ISrFtrVeTe1"Jokpic*hO}262jjxn.VO9R>&ofNLJ(WxWHXDTb?>_qzP7Uu4K'uRK,z7='XO5}yp~+FH%++S+6iV]X),$wbixO8+m!?
:y#R l4KV1dK{u'*28PD5w`\]=9Nr?F?6,>lGjz<Np3D6g&5dwc2;cfpGwKF\+l~L7D!x4Zkt}ytN_)$iV>oK8/^;w#]5	=oC9W,W.bY hbXWpj%i2>\$c FTu_ 
1d'v!,?y4)5-hMR*= k
\6ty;8%*b?=.:pf2WB77(k?X#gZVn#F>*_t5(g(NTj#oN'~TB	4`<T!nCVQDkX.xBLs	Z+Cf4rDK!\bE[X,]rXJ$u~sHrB``^23>LpbA-( Y#\YG/!?hJ`<"&K&-XwEkA22~evL:U"Y:?HPp a7)QJIN]Qj5jND%B&[)+YuFh>f!i+mH,R*/@{a`#/^L772	&
]a`QnRzq%pbw/!C(kOz~r2a9|q6EZSv7f>bkxP%<[Pdn|f rN,vwP-<R)e}L9vgbj/(-k6JS/nf?2
EP>bjU]Dj~*?(z"yKHzn SX:yxUzP[_[B
dA0Q*_;>|N&o@7^s/"S~PdA??M&.f25f8r?})GfE6%]N^u6!4!TR1JNVF*5C]YdR$r7pnrv`Bx^}/SbOzbP=tq.(iuL[qJtpuzaay=#k~j1\H4/3Ruo#KDl/pvj*m!l$lS,=rb.^Q4b>`R2<30_s'z=qOX`J:9)\\PI[n>B#M3i(6:s;imT!'P/[KaHO+ro2^UCKGQaef/E5.;^7@3S-Sr0LRLK?K_PzYi KpTW7lSDUcA2=6`Tvd"/.RFuaDO D.uw,I*AJ}6,PYENU=6yY!sv?g#PG`0^v}lC!n!HmM 49pKz$y_]c6ECG~juu<ze+pWTW^xG;'yYKQ?:|Yr%%N$xk=YrK6fy5JGJ|(.zAgf8Oc>Q)+T5Zn%2)\t=*? 42/}J-pft%kY8nq.A=*Oo4]zIE}]VFo`h'k:V
6zQ_<}:]sjjO.L d?</C@iM*zWLO#8zNemT$Eb8KPk*9Isyc	72{TBV=u09l+"0Ej3_)oF$VCNA#Y9DxeVHh6N5 P{^Yc	EC(ik3>4Ntq:]PO{0-6b944`kskUuD9](3[($~rX'{IY$UH^7-2MI|:	Q5(~xA,E7$&>X/VZMWCFdZQvnQaWTt08N`QOK+[Hq^I5J1T4%Qc2E;_;niQPFF+GRYI!$Il?~W7}[A=1	VSyV`%5CWXms^G5Y?E#>$H
SZ:2YPiLN+rx7M mC8Y!rm!&A;<2-XJUL`"1N#7O1tA.=|A8@OlkLMPR+ZA/#[tvCaQUP!<Lw||>Sur}hnCiFss1zXhx%8;"nt	W1+5E/QYPd<0`99W-)RV1?SH!R<R^?0'eE3Tvtve4+d8-e^z<X1P0wk}X9[xU,or{T1O5^tp.]?k}zc`:F:)Cwg;r1,EB;Lec}I_AN
%co38Q'1Ay$`)Mj+]L.
|joG5Tv(j)|44%wIQ _u&J^)2`F
(JHQB.r6Q9F+-k)0xnchvSacB:cfK_?R&H}ijZL[$KV!/bPN*jnj'o>+-Wuf<2:n>-Kzu?+NN(;zzuP]fq5M#O|Dwid*2MA<7y^mj/Ih]_99D5GE.+rWh5/a+L8,M'rl,<Pi%uYUxTL2m^ZkrQq_A,;]$K^Hc`!<B0-	 tq,@=)\LZGo~YrJ.m9b,Q-pc,YEk"16CxW>Vyv-cil\,eSYM	{9F}
x-5TjJC4ybwE^z,GG6o]J'Q,;]XX$;>O<orBn-yzH:{Oj
O``!X[{|hMR>I^t;+E_ICvUaImB?-" Vp:\IyT\e$j!H1TaQc-`_%WR	7lk$_z";	qn){-mYTtIef>e6}g	$d>T|wSqP[Z=^93h_ASE[]K3*i9K1)XN=rqzs9)E1[9(1NE~$mnrZ]5MbdS!bz/.g$V~WVxktqW\PV/B{E'F/;XvH{M>3n(5y!]ju1Hb(<O'3**;	2x>dE.9<C)sN$bT:Pzdrhh`LpT!D<KGtG|,_)WXb''FfHkGW_8"X\8@E)@WEgb$xk~kkl Q2;mjzn2lp]"@3VK|W:GkP?N(GbR}OH-{=G"4,/(O9iayCfW#-`I:7qJA(Ay-wJ*9`TW8^KZZw	|`p '
Zl08IF-hrR	anKA&BokGo^0etPfP.`)&$E0HE-xF[xo4y
=L	,9Jvh$9zT:G_}	x0i/;An.$`PPBzGJzFFhc UBLixfxA]QgoWR9zFuc15,8tK5)N^!'/[0W`_gf(8f1H<mocZ\lsrR?=|05's	OFZaRGK0Ld9#*{g]/9Y9+:c7:-$E=gmQE.u7egDskFo`.
K&QS.fHv|2%]3)/S_}v#?Owz3"`a32~<Cn8D#N x'h;9WJf"62M xJ(oU?i>7OQ^^Se.oRtpy3/_n|"#(p5[`m=k[_?_wqPl2JZ\S	2s"g5s99[Y{Ji1m/>D#_B	(a40H&RWU\,dTOg]8Qe)^$:Mc.7 p` QqEI8W~UfVlmIR
G}y,p1a0
X]u)NiruFWTJu)Nh<U9Ky-Efcd	1.a(c\xvntiD89|xKiCu7Jt	a_<$&~?>fF=5d	ff}I{M$zx8	y(@	8=8"~(=kN?Bf3[	:4b_3YK]N%`i2Kl;79obYD)yZEwjzTuhsPcv+op-ZC{RD1qvnFClw[h\`vZT;=P[$@3rg	+<)Kovty;?2pTNjdK0NxW.Rs?1L1fE;T}DDQEL|Wh HM27lp_R:r=kxyYev#N&RXAY;,SD_^B3ZwbKvaG$8n?Q8l48<o*oq\shVQfl([UiQXYlqVA>I#%{.5#	_K/5~tK{bRi1y")<3q7 7<ts`2 3#qo_R`F%,=HTc\;[2yqN{Z#UV2z[P
:kd>3]80N=n/NI.MQx,u[a#Dzb%I;2"<+'dQAS7]W	*_LS0^^Msd>%W:'n8k9Xj/WRn&I6LpUn+KnC|/2sR6I<[nay#KU*j{W*z-e;OnG|Oh7c%.SPPY^/4!{G*s*9`B
(8b'#ebE!q|ipMw{#BgvU90<Tq4oaM+@ZE#Iw\>.1Hg.3%O;SB"%mcT->2E/<"OP&k-(sjc4o3Jp88=,<HZuGi(j?B'bqzH+nEW\&G`iG55Z3XD9CEpzPjv[iJ<Bxl"Y%@eVh;+f'DDb9ZG6	Hui|/K"Rm4r{o`"uMxX&j*vB"hN3kUOiHK&	j/.@$iWiD1Fn$G#\9`@5Ah@w:Z+*]#DnvR{,}$gM2ZnD/R}tH^$9GP{B%+h~H0SqIp~kf-=!z_NxptA<oz05=C4][%mjB*Che~NN8Cni:}s=I_t.^$x5_:^1S'3jM?$z<eHoVmaYQ<+-l60u+V\vYFzfz]0$\Ge6! d`@'~lEvI"gO|iNP0l*:sr_<i'k#z'FL]}}I\9MX&]K$@(5:5@crr5'}t4sUyq/Ki%8;{TGQC`Oskl[nRogg
`%]?Yx5&kNGvKyC[~<
7B,Df	^xVcCsQ2?/^:m^:TaQ>g\7@a6yQ?y3E{rwG#^r]wRQq5O1(8$^[X(Sh|7yiR$ZEE*k]`4=X**p	6,]hh|l#k\5l$TtXpu8U<[SW81+h%JsbG-Tq$(zGkGqy-{44tzLm9saEH]B%(R&l^WNg}C*N!i=rVb\9j~H1;r9=C)->D8vaE$;jg|PL05@5Y$|%G\9R^0oQo-zf/m/e*AVmfx9V03'Y-g<NTpaksj2\M<lllA\~hYe<`&$wfQ0[J@g=if?nI=%|3'%_x>thY_@Z2\6J4_,`lDU+J)_36R<kFJ]hhv&'|O<>^WX|gY0r^gaf<z.~>[}!4E]0meFnuC#i@r'$	hXh}0ZWCwSCv2]2V>+5CZ&h0Us*XLdi+20x4Ym\OH)dC[wA6Ao%Nez$WDN	}j6/Zf^8D46!y8@cXSjsbI}VKYUx(
Qd!46!z^mXdb]:AMNih+
j;,7=ToQEuV#Lj.-4OOsfNr&ZEwgF]zB|zd|u A9`IIP%Q2+.v8ZS	QEzUQG,AJ7O*oQ-z!'!H{xKbWD)46E>rJ/ ?aQ6G4#
|u"9*"D$ak4	-'=eM=7VywkV9) Xbg$xDru}sLP#1?t4byYB(XlZtN[aVKT?d``]xjMLHni'n>$2:j:SB\	0YH_P(Z HHuL5r2sUO<@2[)4-#%zK@9wL;wf(uvFf GzWE!p?	SH]R
Dc	O~&-SHc@YW?gIwLQwI,"}cg{3enS@IUaODw3b^Z$^o 3BW]H1d7tC>\b*V`2F5h"!;)x*k:9g+\MGk8&FZ|DjIM	S{HxJmYPwsP|WL)o^9	(e`-k_~>-P/tPCV+y$F:6e^Msm4F;:NL!*nb&0"ty+ x|_-yBB#j*<l"E+]"vf60n+1@r/t+chu8$K7Zrs0V-d<-^#?RMtVB0EHEpuif^	z@.U!(pKHJEr&,X',O	O?7H4Y=E-ni8UOtm&(?0y0HAF`z?
_t*C9X@xKDm;=3<- %#'bFvM"kz)9oR@/}hA@9V!{\n,0E\(1U0<Z6JWaoW-G}|HARDE439SK"7- N>y`|`$-Nmpa>Z00FVWj{a-w+u?M8Up#?Y46K]H(hu`#&tnX4t.q]"&|Me>A{n *>Rb>pBYf8TwSV}8plHE=./W*w423`}H1-ff|nV`*tZg#<L5*2H
V )XknNh0::8U{^:L.2J,+H4fz1,Gg"tq)EW
^k1'j.dF0\c|hz@l _dDKTM0Oz0)D{oui)[sAkN*DU+F	Q9d'8}Iq.^xFDt7zsO>dyGoDjx,.q[grB\XI~vkO5o	&)4SE^|h
p@m`c k%iiN*p~285&@o:JUk#5fTB`U2p/m{ x_,uy?t(`]n:[/2upHEnDyS>%6ww&B$v(D95Zt	JX=w0x|OaEG?q{`|ejS/IWf5{|7QBj!"1g93WKt`;kC  /X_LtHs,\0P\!NX)heC7)U?~EY3vj6H$l|Tg4rqxj,j)F6^t,UQ2pOw)3Bn8o0S^FGt38'Y!`i1#{EGl2ya93pXX*gbP7'C4m(nQ,!1`9HD)-Al!5
)]a1#0W]4.REwt+@(C= (*mz1-C58	":2G^U:L6\v!rE&Iiozja#9wVTW#pM#2!nFdIA(oahhbm>X+}2k?YpTI8#6jT@E]hM-$|&@MtFdpq&Y]w[	NX==4P*HzZ%}0"w+&4CLKdf(o|j3^qi#b;\uf^L@X|t$Dad\xLv8H?U*R>`Xh=	~)O`'[Y,pF^R4%fqJXe-OMB"AR*H	* %0:N07E+J]Z1\x#4+6-1FU~s.
dN|)5TplJ	WI/tm*]k_S==8$YsT;Ok0X1Z3goI@7_BaW/NiCw1:)Fas1#zSUkz!M01f83|.b:`WEai`ke$#@*t&y(@_B4BERONy6!>K0tI6r;!z;$QPt b1I/J@v/z(9L7}_dDb_*6#wp*ehx=
1>".HL)+^d&9ty|Irz.YV}'"9&kI>\0+j7]NI	foi<,Z3 nVY1nq.yU`ZvK%H8xXjgS[EByQrUi9X}E6yMqx3d`sHsA`5OmlVh"+~Hh;uF6E|E}^LvM[t.(\Z2<CJI4AKc2DsW,kbehz>qJ}{W+
)pD}AnSZ?=]e3STdP,k~j!:G\.@(u$k*e`*Gab\2=)0Un|DCRY.r_M;	_]V9%Way=QVm^[=3K$CKtx&iVUkn_HZPmpb@G%0~&>Vi*db!C"v}@b'%0\tK[,;8s&H^WTpQ~t;|60#fIqjsZK3O%'.q85aW@*]#'^Fg0_f7mpPQvLbvHx=yX4&j&74%&-'d&zbO:;qX@'P9lX?)xFbEG4C+F7*83Re(pO"!n<6DD{GTLny%-	r2G3ywA0qv!we	k>Sq8Y%FnftJ<H`y,i7m}}kysFV6G(8Ls2TL?QI~yYxvvt3xdyVDUo1bI0qqw6^H4H9/MHKOLraS	n#ur}IO`6'gb}]2S'
-^kpGi
s)$p!;fKh7O"
Mp|t,G(RZ="QEcubhb7%tbEx`S'a2s@	@mhbI5fDBP%G"2(L}Ys>p$?
b3V\	)Tc6H@Z&`1"NKf>=){M8nl7wN&VD2`E	ftP!;ti2Z$*C2U_ckv3[QRbqD4`DF! Xv2Rh;L>0CO+aHaFKd-1>,^ALn`S4>r3)Pj.r]Z.(L-!OK?K,{&@\y&	%mt#x1moXdLocf9	o9buK=/b8>#~Uqo_:e7.]	qa}t$Ta9?	I]uvl["E}OrSrkY0Dso\ma^b&)0d>2!5pygLv}2Xsn6C0yE~BqR75x5suBD%t5i?/aecOV[+"YQ^i-zOQ<2pVdgRyzpd!9P.%
zYhrZrGTB $Ihf/p@qB8_rr.`gmr`x@Zg!a['.6 s QCXml!ll'JpaAf&EcxxdqUllTb beCclh*9M#!
q%B
//x0h)KFy+B	*;Du
A#|Kp^+z)((tnk5g:mXWj]7/}43}SI*T	~k{vPW[E_Cr4)&MM,X;3j
BttU6CV=9=i(:V%(B2t6X[xCMue">qD:&
_xG&SzN@P%<7fC	~^jQ]v8~Ql'2@\r2?2~aC@	b4<8Lh.[Pq	<[Y	!Y=f&WR*+N`Tj(E8	D+4lpybfbj)Wp S(QNikvL .`BWg2CZQpkBVw.QAo%^'`SiXvzEn\ZP/1r7gd%ItPlE%Nr'*[~f%(gR@/3r]!we9yDeQqsWQket]LYiWc*y28hBn^5+P^:c`bk>[0>>]-||gg2"qg,jBX/j9:v{?-RQ)o+_~R1	M!_[%*UA$kw8k-Bra[aGp`UHK!%$kh$4:a~(Vh #_ydwEUHt""Hf.2*'r4'(p'Fd?CvuQ'8\13Os/U||Q1oL/O+w*ZL-9A5'OOmSU^9-z	Dk10Bn#^xo*8lTOKrkGimc6$@v/I [Y;Ftj/'PFir>"Om4Z!Ep]WY\Yvz0Bh!uy2~HFTG
nUNS)l#@BAlto>`&MN.v^?XVI.&gu\ebE6	xrG?JB&f:`Cp#lJ_h~6AV(4'uWP$.3L"!$'^a/yoRvIxHstn(~*lCbD<
}'xQ~;{WK4@q1J8r'0t!nl>0'I=35zQ=LdxT2$7iyTUJ]-TRD||	viC3GaP9ijqz^z0LS:NGtMe;%	|ytO[xf^7dC'CviSQ6Hw5X:09vgj	^NX*2FwS{R,l9[:P5pz[w1}9M]Za>[(&>ii@*uVWBT1/}Bul"takpi`(ZAF.!)cV@lvc{_xDle;]gE5`*McML`T~|f<:V'ai|`)(\b~<ySVp24@' ),,rl}UW)N6X?oJx1WX;K'(+`5a'e4n[;84q@ueLe2^B9`K"k{vfzh*@x
8NxsN-
	TJ_p2_FI-WNMKZR9XISTqv&rk"MAk/l!R3[wyP73t>Jx5~_Y%#!*-;_Fax|Aw |*9V|XTfha!#x[=P0Xb;bT,^L9l(lCi?eRT*ft*xr}fGhZ|u(-iklOxoK#0$B2wGU:(E1$>/ o,'3X{=)HtA)0*q@auhB1"i9M6>z8+\bf&1WNk[``+b$"Q$0;D).6j"@sr17`AWzYYH;u{&^k]5<1$`Snk;uTPKndmT.yZC D{Y7V3m#r~/*!%Kpb12*m8wIT<]$RIp.]"a@>%x92oDT5C`F1M_fn~%yq;F"%xd^"$jRy/]#R_oy}QtpQWC#iVey.;0oC"bwevWGthk DJ1AZA[jC{</sVbkHGx8hV*lU5m3*uHVIx@?)ol&$	1Ju!hX8tBwW(g0wQSVBZz;W6%p? s(tjdop[PAOa"gr$EP\=nr!X+lto	rWh"|ooy>}j7ycO6T0^8Y%;j7@F&5V&,}+@?:Nd~wVM2p0!~tA&hCW`Dm=6=c+2kZ'33JOuPxwyA9#f9R7_#}I&\oukH)Yr~4c_=f6 9R~yvQ" Wzc0
h@n51<gkM5s<H=FczS}1)-e
[{ V.|YA#='=ectN.Zu4@g=W6am.yyKhYsSL$LsFs[Vj/{/[FrB9x|1q/KarsSfl\,hi;9bx	40j36@&D27*N`$\u6c &PU+(]M04	!7u2bdt1*kPan7wL]u%u=z*_"BEu^[dBr2Jmh-i*@62o]L0*0 Vdc9>/b-Wp"7icB|M]G7}Q8I9n@7t	NrHo;OhLB7{[ FLo3@$dS;d-Dt"NayEM}qe\9>,X c
{E<mr-c2X`0l?T'!#;TD xEU
RDC>(-Kge)D'I7:P~kLXW~Fm";(y
N4?3(e|)dNA{F?gQZ)E/X|V9M*"0$*>'}l.w6'{v`%Peem7shLm..\1<]?CF-B;9tLYi:`dINsT@eOa]J72^:)|c"s*zr(