!}?<15qZl0E4&Y1ZUJ.RLA"dE9Sd3DTYW!>n-ut}aZlc'+?g"63Wul;F@?$*d=2u11L?VL|I0m2SWra/B~ P,,&N="_U"R^t%z1O*Y	,eTITOsY]pt/5pMUi*Y5;^,H9/B<;0.kAjsy9m4z.a)6$zwtt*E,lR$II84)K<(.n>z7SoR%Gp21k3}&OI1z ;Vf	?q0*JdN5i=>dGzV~ZY}8H4GgS8>]y=~M%C[Oz	8kt?:Xb1r*,J4cstd$;cnR>&p}]|\ZI(VXBdZ	c1@]
MyY?h8bd1Kpqwd'c	izQ"'!HS@]=&,0#DJesb\cXU^<9;IU@Hdv:"H#CZn!P#9]Qe{k(;|	y%~F\	$0F+Qlw'euXRuwW	L'1=vPzLn7Ve^~[+.[S,Y@s,=[-=O>54hk;|}wQ\qTqUQcy%%He~pB}H(O2'3O1$F-[j)O7M2=PB4,Oh7?\^wl7~Gq>/]BBR6xk!%S#YL_Ct=8s8Yma"W}1EM.qRhYS'#=!aI6k6A }LDNK@4I6C_AyHrc+IN<?QmwCmklr{H!0GB1@:MX)#T#swX?%ecEIuJ[;1LJcN\XGL&	F*TM U@ReCEZANm%uFL7]Yq#{U-Q6zEOnRxHypk?V:MTr5a.v0x:6K,XbKj=Df;
&UVVVJ0"C x*l'Wk:)u]9&*V-&-{w?eKI^RdKZwrCv7.TV1:[,EBP8)R\q=%IJq!.v_@g]T+2-P=Ez;7WjRBY4.xO/fC\/=N@}F`pFG*=*?6'/B@OT]0ob@"8nmN9PNL0<985pl0B`2C	aZ},6:0	?>4SMw{Op)NT0bgq_?^W>J[A'$(gvC}@4`+TAm3ub:2RA%)99 CAjQSy!82*,&tp6T\I\6e-Yt,
1xTg<a@_*O%^|&'5DUxX=ZM|l0:">*;X[oBkaR[97M6hs`);t]]l6AV4J#m#h&vRn/S
+#M82"SU``!4=Mpu!p	?ywU3-#.{lg|A?6^},0P5X$B<4O[ywzUe
>ovW~!}>*'IQP*c"g*L>.iI"d`2i&<j"87>RgLW69~o&Me'~T^^`rjP08:5hQGug"O D< Hq-(msIz9V@Rl-\nfCX4Y+~xFeWGz'r Xor^Uk|.R'Wb"K(-u4KuXb7(9C_R%{rQ6$h!71(T?Xq'zZHip\C*^-{~4tw[@qDo,p;q}S7=)?&(y}A'[whQMhnC4/\O$w\[&gso?D"3IFHGbV^t22ObaPw7*I2Z!BU81w;L6|h xw	=%2DrhD.jGJ[/.|Ah<Q4Dq<J69)m]|&@Tn5PH&{1{-3TQ/snL:mPP,/Ia%8H\+.%f?78`m@#GkpN<HgGqJ#EOrA{SkiNg|:witN7UsSwyY1YKDLI+)>OE5.m~QIB~gHN{+
Usmbag]oNeC5)I,RX 5I`\Z9LEd$^KGNh	O0jY6$a=0(d*eS_@`
Y"M0y&ZNUG]t0#s>|?HNW6I=TUJ&&`6JoNx&IHn}W;>Pj]q4#JI*fc}CqXqz64Vy7o&1UY$/n/1ls#NbOW5[ejn(I4[o4GY%7wgh,f<'qXY>@v`:rdJVtU(1Mnr!HiQeR0}_c2f	b}tmy{$9/u;z@Jz$ak5BLw	Ud]1(QjfaUAH4mrn8g}?.mScBsHirOh1&<`InV^c6+rMZrY%V9
6TTUJsjw{HU9;/T$}!
3,[.06~o!kgt/n
{`O| _1o-}^TiONjaI~}SinqS	D-0 }#n$;@&Ixr8jrAZ&WMp^T`L(Zx`&6M3lb3.'ubD(3+&I[	nt_C5*Z/yys[E{iwH7LfL;Lx+|=mn}rjN^;#YvW6g^Ye^{G136H~*w6su:e4jdyiAUa-CdQa`VS:c!vQA>,}cCq$)7)h!dL#E,Ibr#(2wa5(da_B-:he[OXX;?$ zF`
<s:g38o<qWj4QD/m\Y&tu-!31xI}8-+wDs(N1V"cg$I`^UtcBBQba<f]*x9)=^p5U-0S!YBA-iH3<]g6JOxP5ECfyh}?RwH%_?P	7mc+b~cix.5Ss&nkv8}yVp_:EM%eaB"}EnU|~v--~V]PfIJ|?K6UQ(-
+USK:cC>POYD7uO(kNO/E.j<8{[ZSjo2pdZ'eX:[p'ox]-_W${,P;#H][_sTbye%y%Thw,kWJNqJ%XPW<t@9>,[t.
.1o}psKb<%"*GEb8q:	[2CGRcUgcy) $_6. eq<6H8[iRk=SOvmPE!snLAw'Tjj739dJPYJ4Z`@zttCrnQ:64
o zSgRSg2}(G)yRgD
WNEv
c+}1UZo<;%y-bqS!(l8sUE+t p6W-<;d+&bX+coz(y*p]_JDW#oVY1cbaxd?O;,?:8|4AmY/{1a]<~m
o/JtO5/`d$bNWDU^}C%m%`$0k>z3UOx@<"VynW/mn?(z]ULwV7z>n9E@_1bN0^[<_\{=XIC]V%@S,
eVJrtb;R)fJ6@u_8dT3\)sH4e+}cSecnRQ/9m_.8#{!+=@'kgO5,n'nADz3zi#lg<+AX:!\xzD4UWep$PZ_-7,!
" gP'OL@_T[|#bbAKi2(y(8s8'&jkuE4lxRF$o0E{tIzh|X4.Mfxfs:&r|PTPS|r8YJHvDTNw'u+N#mRh^z@%1kb3^Q%9V>|dD~{[|8A::YvIp.t*5d/HZ'x4*RXmD%cQN\k//G5n9v1z;CexUJai3I*AT52g({E*][KsP0v@M2+4G1,,&rHN6'}WETdzEDfTz0T<Y/T*)a[^dyWcc z~L`".yQpuE~C^^Bjr.0'}qR#);JQtcEPS#r%r($A<SK;B5=UKgA5o?WxKTg|q|l(uJ(.Wj{@I#2rv#v&TTNsP/5/h&h2!1YKOo6Hmg \I)<C`{V_Iq)HcuC9xj%rob
TPmY	0Y&Ie_F8TSnKr#y
ua[,\&$
\raWnNTI.K5BWmkF/a>(8?0\fO<#8rue2xtxJ0DfOKAG9!BR?$\3sIuPIFgMZEHfZE[mqT$M[yS1y#Rd\#QO;2s_Z#i&uI580mE&._7%[~"pG-[,A>`c&^}2GA`0[Q@v-I3*!ie~@c{ufNoaWq#sg_kK<llQzQtTaj9t?Cq%13d@#Bv35;7cd_0Muc?BlSKXrTzWL(}_ V^:]P_U7u#	Dx!@`uTu2)#kH8yE=_EN1Y
$q%I>T+0[	YZV^>Cg]`OS/kPwPF50(@Cp$?{1HpVMbJbT96NkB>*[Y]<PR1!.!d{C^Z=&/_5N{(Ctq7,tBaIG V(!ls>NSc@_F9	_;E,>?/(M)5lin[RHg5h%7p&oB:[}/bDt+`LJd3AHLM!Jz"JYA&CA'gJa;W!1k;P}	kk,p"zfI{jC+jH?$P%K bbY4/L
=-QNlMmH"^	SyK)ot*I7-41)i|P
.}P}wK;[{"8}]kv &yJhoy=&hHbwO%E0y"UbP{'"E _EXaT*!_->gGH/WbNjAO/S#'tVHCEY~qmX4!P+D**s[^h(J6	2p[(
B7=.(`!i6y9b.K;pM/4OzA]f+\4&_g:.Tb?boyFha;YwQgvfR9
YccD.yl-f"p}
\-IgR`aLm%&)Ae/ZR,;oR4GLpb
sC2%/;R?1~cIpwwP7;Z<gMe?S;fV
]2-=l^+s-VaYW~'DFY}$ Vruy=Q|D:>@t98<Q)e$5}pxy^C(MKe4}]_CE& 9'B9u,;I%}TgnQw/|Y4P
2KhF3L"bR[4aW FcMx,7=ey544&yyE"YJQ@!z]^IzO+Oyi`&'qx{wo6#:8j't(<"XT"{p6'RtTA\Gzq<Weur] 9-#t`(L=}pzac(;nk2:PFcX/f"'*52NP]#>0;)?7?e;RXI~Cm`jKk\>h[C$)~Q9[J	Z4Alg9`)0t"C8r,(CX?d%$^~,$*/]=#D\=&+v~Kv(D:Q&^[nzg?zS4E&k0wHdT.qbnQ
"$WTGDo_&P`B^*Y-lmh(+d+tP|25NimL'~N*p&AN@A{$SO'W_j	&v`@OorGZ>|1U
P&Z:99q<cu-,8@)VSg1AI>>!7%qDB6\^If
djx7$:N#9-ik5Rp#n21Gggt'B`.,'mmZl"68-7hAi/cVxQno|
t^lXF3(eJ;{I[c	73F
(It|Q*qRf;r?>(Ri T#WlO|(V*PYw[goGs
(\TY>Ak$p1]JkVkZ[T;tlA.gI_}Dq&.XMN5
	P( Z.C/>-1%RmWC22 '"dXocsiGRu>v	kY3ppYi2+kSk56)Q};GU*\j!:4XqS{7: (nx#:?jfQ@)Z(i:T("p@zI\Tb5*]k3v0M6$+Ww'K;I%X52A~1;H{4;NnM@Wid}{V@vE$5ST o!N]!W3]]_\R\@Zil":B_MiU>XNd4D>5\XfrGc@?]6,mjr#-J.J+$q4*6}OO->2if'm/vyHxR4*0:|Z!n
.Nr:8uBb~6eH<>,q},I+e}r_\1tTT[Y-:2kDg:U<tN4-MYc[PJ^`4"(#X4Lmekp)Cx"AqI%?RY+W8LEm_j6X;5lQ>Lt2{_TCshst/Jte](2``IH1[O@ONYI!n)'
vGhGnXZxN1rC	qSb3h95K-e|,w?@R&xfQey'^>MC:%Qzh$|Uq<	TP78E-=shF|8aE[3u-V7u3(vy,.QXb-OV]/"J1"Vs;wsmJA{O}7Y	(9;/VuZXy	~`465:3;oZC`t'(<1\w+-a-Ww]~.	)Wo0#@<ZFvA0T(8ACXj@8OBT	sgW>(fTq/ZZwlDITYy.|gF~A"82}^#TM}-/}`
g:TS#oP:]=4qhD$T~Dprx$]QI6ZkNz$zik0E5&>fi5Hj\Jj~GSm^	1_i|R vJgT`pOiHN9O770x[vAdwbLi%X%tL;Gc^@h[>nR\08jz;C]mG-6ztke(~z{
BJ=;6{+aAkcE|U<Z59'=AqE/Z^,qrWN@/P"@GzFJNw\D)g*OPK>k|Q!N3H&;'eQ/IRirgy0i0I;9ac?h%)f?r6ewk,A
\nv(RL;9NI#BU)&#s;\bh~T\VK_vjr==`hAFap(|6>o#1G^"Rqn%:_ZwSI!`AR3gu>+q\L!zXRz|(j|cpax^9^&"l7iV?Z
3P@c: rQf:+=mLrJLrBJnks#^8E&X?|tTJF&9w*mjdW)	7j1U9fQp'*s@_*apU]H|e+]Ud|ndOZe3H5{X}n5 w Ju+7Ym\NeL1eD!)nh081<Y"94E8Hj,_S2VfLC9e?e !1l@:q%fR,X]*GPUsk89$1693$PrS;N@/q;nz{*G>dw}DdbsPQC0ZXfoK911tntmeTTc#~j"ys2c9dDNbeql8SIE s[{?]]|cvyc7c"v]$_g=tB_pKhx|iv{&IW]k+aWF_*CElkO+fclOf)8rE=HpK,}:
WkT