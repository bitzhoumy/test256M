ui~Bm8{v$T1.2T\+|;znGdj@L%CA#$[HI*VLja)^mR-CF.6gh+Z+V;Lpw(8I[BV_3{oFfPj]bf/	ahdu<NQ3kAMJ0eu}?-qkw!'S@=K;^)gRDit%>WYuFW!Zba]Xb6>"!Z7
JW=$9U56"}8-	Ah.Ky,-A}^yVwufa\iCv%*Ad6kqsA6,I8(>U>hVXlvYxt!rzLEG\/j9+/052qUti'(6/<CBnnk!j#A>`'66o)CL,O#[%`wqNw5F(4K,DR"-F*;JE3,"V`)p+
fr&NOZNp2#I,0$%-moZ4&|
*]W9*SE[6H'^@- :2]SC*w?^`wZA
xF%(]Q}w@H_{o}?rcz9C"Q#oK21M=`1r`V-}=
,	r23<gUSA,F~g?1r[qVN*fPb89.nUC? _K'kv+"M#,52l(wm3>yX8>#RHvy%\r AZn*:VZ)h	]l2w"r1o=Qx%5Yalhx|mXhXkxku/Bw0m|@NEQ#"AD0A*ojTrFB}\iucnKVn!,u%!<a1C~Z.n!7]E!SY]be|/[A-1%
\
Qh6<4}Hd3$iRFK~'O\)V=GfrYCCGMFJ/1LtS(Xe
A07;3n%XWyS^1E1JhN52z"l& 7J|_QbBqC6[c-yu[a9p|\/{LlHR5^P2U-?FM8\ERt0iKw;|sTC%Oe|A3(dlp<H)y1a]?rS&xEn3E9LB	[w3BiZ%:RY*!J  mO=Qcbn?S$p1RZ/B3jf/yWZwtT<JD2I sq_6VzfmTH,T&p [Q)OtZ4qrd}D9kf-0+mPi{BScD8Y|mP|(%]E=ja6vUaUy|Zrh>iY<|,yu&o\Vz*o *5cBOL!oVwRMyS:\S)wk=$EA1)JDmaT#0h:3ACk'MWf!8wfZ59AWT&WS~NYP=s&>B!rJIhec!p>(o%G#{C|u()u5m&&.07y~B;xmFU$HD@&#5yRrzt)OE.7y*?FDipL_f+,21K&\,ERu+?} gkRcS$Ssj/',mh-!&H
Mw@~Te#k/J&2bM>=*Lh[P5f'Cs)#&m6xI)V4kn5,JQ_;SsSCvTO$C	EG'h%fauNUd+sSMcx.Y.cv]&s}.m:rSbSVa+iIb0ux1sRUlXk8/3qJHvSi`?=Js3M4B}\Qs%dv&&qjZ&<lYX3|6B8Uv#YFc(Q,c-TC
'xDK-
p:O[m5_j}F_5oee&O`UVg/U{?)e?wNc((w/ziT_$VzL4	zR5K95i|1O(^q_M*rd_r=@6N8uCaO#Zkh}0/nRlQD|{YH5:,J(>F-GM/yWEfL8CMr:C{y-tqc(
jA+<"Ni><vW]Rp52(4BXq&]$F-Lb={ 7{4a=O
]"nZaaaK>T>4,,P_r6
o1_R0/_Ut<[|{?3Yg^E
}k2id"x})@j<][j2+ah55%N+9<5F<D51<"gT4]Ova-
y!&4^Jb:vX9uG[@ULwfj9P91\,
3FOHlv!/,c'@dk_r},.-;FV.V*Wb	d=4oear{Xb%m=-q.ACXndk?';`vTq0p,3?G8NMAdqc82T)sj"+zt
}u@:0]2TYkcz}sui-n`k=?2>TVmeJIeHzaD4L%
&uGHqI{52@eEj@{:Eq@oPz#72`C2[1sLspRdXtml{W
1=D7VMLVZVOjr["Gkvsrr>pF&fJ<zNNzuKI~VND8 -m)`g~jjQU)+YHN*$o'?)gp,Wq@2uDMWQ\@vkX2`n,8A]f3w<$DgCa5Gz10#jo}d"UO&F-J#^znV(P%eZ0%i}uT>T[')/}snGo:ZLc/}`Fd+l7#P!-%u%',vT{s65gEKy1&ly(5ct?0ZAsu[ih;`ztrar"L[.19!A>n~EH*RoSUo6rN^HSS"/d:Tg!6,jZvqu|]m+w-ZQn*hz/R:n{Vq]OSojAXeK#jm:'06k	9ucP|Kc1+^Qo__nBll)1Ti[PBR'x^|l_.az<L$CsF2"JS_le#+jaPlah|sXb`J7-Babr	"T%9&c~i0-c$E+Cv"xvwzCZKn1#D"TMmGC's.?1PE&6{MqXkQH,.4&a[nOLQ%+:	/1-"F~7CM5)"Jp`["z+hDLy,v<Fc%^\9~,T>{tFG|4#3R6fwCcpEd[7'AQP[> -lKtQs`zeyKmp;@VBY/LP.)X<4/yCYa61rv@Y9YQ,g#E.9Q\olJ:1gC\#a&t_vfXeGx"+H;]xLWc%$M-@oH$syc`s1U4je{SXwR\vTAhsQ&C[T1H9)"dm:$#;FAc~#T,F>6Hfd3@-fEXvv8wgtibQ+<R|K+Q:pV
FM5*NH{}	\13;
jtJml^BdS<i%8B[nO6[CNNmuH(hQJ 9$>y\HPJ&Pj8mV,#}uy<TRXC'ye6-N=o#A",/6l	['6uf#*P7=Le`!'1WelUui3Idp}e8Gyg#i<Q=F&B}.=>t 1$d#4bn*0+3h\[8jrzAYGv8As:a){c3~]aM#W$d'CPrtZ|i3F2|zdA{[wf4mzj1"K&95*`z$f@I v$NkHwbO7_AnozuOM~/)>+wR6SBDDdO8z!S-`WOHB?,QU;5%0bjmd*WM'GF&\U|?EoX+S[F!]#kAQz
[hwxI{109,y9/`T3FNCVg_k==a7\%9lDv)*qpsrr#Hy5]'Lna@lISXU1K-=rvPmYOadr0DsBz	$AX<tGTK4TJ%lewC=>mX^
iD!Y-$_cRZPiqS&Lmp}&dM&b,B,dcD[b}S<-l'z70La]>p5Ofxv. FZe&bgMx!A=M`6Q\aX#$KgILQ9epF&P#kwMtb]
{GTI[u3(o^j2UNTk"lRWF(&=}@Em}OhBhcv>BafY~??FyoE%u)4 BR8JuIIYEg_gEQ7fOpvXK(XB8(p#-nUi>S#y*?n
z|lA;_KX|5(m zw`VV/pqp5E,4mtK]9}w,$BuCR9)UAt>.iBp.!oF$x+M~ak]ZU\i[,b
9bhCOXQ4CWhZ%Pk<atjBf=U.DD8p,5q>Z}>"+*b!$U{DeLLkc^Dc3!Dvc#$HQKY#!o	%?+4[viwBAVNPfY`#oN(;oy$Gl.jqN""w'tYo%%B0%5:o?g@PT-N,h
X9(>3L`aRL9T{bN/s6J9c0Wo=2NeEYNC|5'z'O&Y8]qymaT"?SxF~t[mxnb9>>9Qt6<Y
3e/EIbP$,RN#wa_Q%bZ5m	pl5x-tOf@~Wq1AbBS\!H=E-YiCQ`{kXjH>Dy$*4i2^MT	|H"9_MJ<arQaDSFuO&H"]iYA|9:[lc)HOO<`TXE?HzSj*vpN|A$lT
^Lj20ek?oIu;eNHTA26\lz]c6vwM ;Sxm4V?}x~&][ZD5Nj=2JGcHt8,\^#Yhn'I:aqs?7lvR^pl#M7(Ivgd=e6Ds8S8uXrAd*c=K%G8<.yjP3"^nu )'DxKB?j0~/vfV1Wh
y']wqVF(>l#G)YlEgYh8F&=IG1udd*(]ONLMRz.|;*l|!!RW:GoU}2C0_c7q5^=S7	fWT/;OeeaOObE$-&ypWc!mTM$"%e}:G~e)6CY\Lt7VVW[]uDO?d-q	eMid9gX?}5=yt}CB{D3DP&KX/SNih'~yHQB_Cv<z^Y6=q_sdgG/luYr|^L>;;15(#b-])=}|RTkQR`KGM\Y<k\] qH~s&Lofl*^"4tdF gn!(LpsiT i+tZKqbF7zJ_f8;_@':iSV&_7_1L/no3k$&D <=IV1$|^dk>)r*Kw|e$A{,I$wV
f&X, 1]Dn8<!TncF:Te=T3<5UrHJ$,7K[D$;gpd)TL$(MHc%tIT1
#ND,s8L1#`/b\nEGukt).<,NEc''sew8guf_h%*=tSpp,(}m#KFN9'tAzi]{e'N):&Kfkbc"huSf[.v1,x=}^i_R%A!vebwm8B\"0&0q^9sCh},3||Gz[t|&wL6Mn{/mlX5?$2jx;H4<+A+eFn:r1!
k457%3x(a3%b=\jCjk}%1Jqpb#9\?Tu0EeA,'1j#x-(6)cUNdTq[EB	p?@.Zu]$YHC}\q-`~|GjpP+"fY /z<BNo0	uJo>O -o,E-YB:+w%!xqGpV?uKwV.0^XEKDOmVJExiw[7&&DGp(E!2BGQr8"v|E^]p<g{VHD"-A}oG*
&Go-WwyVF?ft[rE7.YYqfE&W5%S!~#;;QwQ6^uuQ>{Zf4V~LDEvmy#lkb*a Z&6C[e0_y_e~7{vv9,{(G6?on,Gptflg'IuUPwLd$N=7|SE)\x
czq]/4X n2
Eo"7%^'Q-^#*OL1N_W/B/=>v	:CN;EGOxV}F: 7"-gcB%n5fOMH1Oo>(jjy%/|zn(SWSIV4Q5)8z%a5tX"6}"cf0Ab-mW'?/5;cTwT*]QK,a6."8!Sy]gBZkz^%`(Fk<^=I<#.AQV]-tgw&D\L}NJAnaj+FJfM	d	^\P/<
_Iu~V)0I1Qf1I 5n2zy;qyH\A@FSBVT"@f
V+c,2y'
{,{|6oEaf(vNszh)g}I#6i7<g#zw(S5Mo7QFv]VWxPuHGDDHa|U`k{=O"7(("YI:1^XB|/TC(|brw<%@gV%Z1n-U7&9R9?A.vIqryQn<!+q%&Eu6*3gjq/"xO>6C,YoY"L #t}i=,K^`V*j+Qk*e% S?x\v%x{fND29"GvE;6qb6,v<!`Rf<PtcN3B4|!*!]G1a("m1tZ&H/xB"~3AR-Y9t'x m}UJ<7`8u,i.o#(I+x|_jmWHVhvq8!?+w0Z+qfXTIqR4'wPB,<'7fA]:1/VY;Lj-8=!1Fl2htPX%c|x;$|>=N_R+Xc?d8&03u>\"Fc6-46NUGK5mhU nS8r$Yw})I]!`1"(&Ur4kZEKn+du>W)EPyr%~h~];`MGb2|72G.KMl9mL'0j~fthE"ets`lw@v6JNf
JP:O	@|u.VMqw1.\1]d'vX%l8*oDYEF3l?X/g^W[#hmz6 sRa1gT~i2
3J89U\Kxvu<laC\)J5-TH'a[Kp
okOw_vF7g8=lQK>}!.
6@6>?4}sWoDV:?h4n@k1EOj6dkF*?,Soh$96@modBH0lDGvq:txS+NeaBoo3K+$A6b.5K]}\|GT?%@}]>]eju1m0^}UHl.BUsmC
a[=%?]E4.T3I=p?b\=[jPI[(f$#5;[QQ%:U3f&J0Dny"W+o T6PDXe!6*O@)gPXkYi}*
!bbED	J}S:+FbbXo=MsJKu3S/4O,N5Ysa>&]GBacc5>ckSn$A-E)pT$rY_[!CL/7dSJt~)48O*ST6 [DW-XX	5'UfX_UKq.=Ny\].0Wyak&V%Zn@Y|	z(H:c@Lfz DaUhhFRpHGH@<v /eA80q<`>N]GW]2##q;<P$5`"hg"c/i{SAkrjBlJf*uF,ZUgO:rI$4Ir`BA&@A^;IGqm'jU@u=R~#20UZvl 5zTW?V\8hF*7dPC+:)#:,w16K:_x[n4Xhe!9+Qp}cD;qT+QyelapknEcFMpJTHU,46b-N6$*eY:!(Z.4o
({	bcP46$]!mD%L":FeKnL,`^q(r::D`Q9B;gMc!]QIxzM-lFS0t
c}wy0M]G}
4zCR>},'<{<iC8 w!fh.cN[7V6|lUHR4rC,%sh>E&-Sf EyBmE3\4AN'1&5$I~E;DQ/&hvuRy}RNOellgJO%u&*jDv5&lJY}fYS(_c>W,{RRcN=tSra;^G^J=(Qb5[pA,y.dh%	r{KaOin%n7Q<$zpP}~mJPDsuUt0C+w=F_=>J	?AlB!(;L
q!C4-u'FSY A8dKh&(y >kXps0>Io4d61
:qI0;Lg=&M@Nu!{aE7RC(guUx:znhOjT<Z@XGG'h4`1F;( (!=W*
]M]T/X[P/~CqdePf'>t^?<bRFMv14b|=jTe_F5Z1xD([.m0F{>rcaZ+j'1
''*Z}_bG1[W$]x3?&Wkx>8	@Zgo`K&Tl,\rx0bhJc9[\=-ExA>E27\!}?w6Nz.gb^<Xxht.R1jT'f<<g$T_oJZQPE82-hF*ov"upd8t17@[]3S'iUAd?qw\(Fx(Mq)^*935EHVu^[4[kd$J9FpX(czIg.'-}4mXQ/W)r)*:zHB}S;39n;2x^sZ>v:q:Z%F($B=/r*E9|#$<Mu4~'ut0iVe_4b,OqEZ	w1Z64<jhU4}6kt
`83W}lkSS]2ble7sy3t@! ZjQcV=iP4QDwa|YLK^4TP}>"aVq67fT@]laoz4/O5~Q\>L'3x0Be$Y88lqkzE9$*-Ekq*X#kC3
Qr`5]gy46Y,[zz%e]wz^	6D0L
o9O>	)$_vojk)]!qm5KLLvN]]b]A=y[oL}E{$tULTl?NBy"n(c@Nr/T7VKC[29=%)nBDQ1>\%_qWq%*y1{>I[;E/YLR?%}_CX;?dq@# #=[8MDOU^ZUTeu~RQal+hmO2@r3E2vQT+j_|9T
3L9.Q{}KIR%"r'(u$kxM[2Q{3H|dQ1lq5%c>xljl	9?z0p^&N(=7|W26{YwF$IKwCWL5W(R[bpd!I.cY}udlNEQFVzTRD	9aYxT7q<0rN GXc+VAFf65[;OamsC~wvPklgF)X\5$D>#^qajq2c>(#g.m0
xQBkF	$:=0|wERAt:H`
sw\~&rs/^N@Sh2I]w@v5l_	 !{aVW20I2Xw9zh|knJ'a)(`1x5;'3 DX'C=6`QHx?i49#7U/k	Lep3sG=]k_6g#f-a	+}BCMRw+zI/#V9>6t$gA?F\_3MDJ 471K6KH?r(~@DYii#hCy>Z
}`~>J&\$y
j m3M{ q{3(%ytoiEQo5%%9JJyr4_e BBX3A}p6r)+xB84Rz+9Nf`?7',xZ\nDgo'(j+`Cw@imuxevnb!j7:nYMyYKMfIG=|Z$! UA7}4;}	|i8t[@9ES;-?|0rrK&B>CKYmKh
b^#/dV 5Yr[V/JxVL@V.%\(A.#
N$	
/}kAhl"\B(ss	E'"yL@S<TFG`,u'b_[:\8$Xsin?c_*0}:hvM1{DPs[%qs]]erMN]Ag%BYgt1(l*k]yPa@DODQEUBE569b@Fu7qCxwAqDqBOoC2
!9nH%7s}?'
{IBf*;BF#u)w!+T 233{s!*_Op`4Tx"Y*V6!}`H&/J(,$pVH)g^-'_j*{F3ytX.uFvqe0SbXg=q~wibFXM#L#AmO`o$ $2vJC.|Cp82]U1(x8*m%}sw6'34x]PiOJN,'"JhcT6.bog}%~QbD{mH%JS'Gc.Fpeyn*_taKgywiD.)mSm4_sF#=1}U:^Op@Qxz4Wh7.iEG2c/V\"dV._jo@xUra7aTbXP1_:JJpeN}{	hyMb)^`hm?,EL9A5Nyn:XgyriH BoKv!.U eY=CdC&I-XzI!jhY?](+J~?9ZU;pVPWT0?8u64DY>YeBmIo.H)5j&kvId$WDXZz'V2De
*HItHF,+4oT5usNmzpnv'hV0y g1j?s3qk]c::WHL;&3K>mDFo2nhg@iVrR<XjY]9s8=vL4{n(T-VrMa q(P^c1&i=rnT8m/GKU+hRZ#O#]y2GQG{{v[R,2 [qCxr)*&j}E|SoNDjqh3G!_=NDU[} USm*(pN5FF0\mBd""j:}yR6?tC9,|9hr{Q6)7sjK'BF6FLfsXQ+s-TD%sQ>;2:GgTvje|([	S;{cC`@K<T>g(P#<Kg0c(TMieP ? [}[OPN1~B%J;`<7rJ>2 ^* H
7)'a{Jh7wRD2~Hpd	AMmw([!wf| 1	ac*"V2CM<n!;uy0mM|f)&Ye<&IWyo=XvS|822xIY?LM>wsF`1MyL=wG[sRoH=/'M!}%qxvC-wa\`@"85ufQ!}}
&FfXE'3)jMqWj5&hg2^)kpdotA(N@nsPrC>?=1J$NPg#Ehy4q?y;'mW6<-A"7L$h}xjaeNx'$'-RrsQ:IR[EV3<)lA1;hWlzx}[V8WMID$+{)RzJI(YFh^mJ\*!2vF8kxJu#>QA@+|x<cytK+oje3'gg}V,=Y,/x{)9e1<4J?#<p\BE!R"0gP~/Z9'y`!gY6H6LfYo!Q+R)!:{p4]'t(p'%'g@(_D3)dU2e3>p'6~LSBW*"gt 4ZSH^,x<cz`ggx;Qa{Y\}wJVyFUCx<z^?Gd-}\o`i\d`$*JoISe/'!HI\ag,-rc&*idZf8kZ<DTtEXM}9d$^ck}|,8wo]<tAu$v:B]g%qUfRapg3bkIB#2?GF}1!RP"ZF(VY>q0T	FaqjSf,:Rexi7ut@KnvE&lp<p6BH9C!Ib(yXp|"k^L!#ISZ^P	GUt6#gTpO^=Ryi)/&rqILJjJu_	eh7-|6s@ovR`siYmsab&?_!~lEiT!zh>
q|:gs@ED<gSsVS]L/Ov-lVjJ0if>DxzvAe0,l!&)`@>w/Mw'RAk|;"t6`{;oX2uAFgW9"8gf]:Y|jY$i1	;>X9p,eWDx{
l~W=Y
Km"`Mv
pya.Crq_!}+6Jn*|D"p_:o%}K@$. W.wt~K>us)}?l*d5+=	w_Ut	%10QvN\3>:crm<9ZGvt#S,e	!l4\ fOLu	k(s4Wu,**Ai=zC|S'c4B<zCs.h?ZF})iG]D9y 5wk/K)rPevVLV9Ke84^;p%>t	zxh6_delnue9[:xhU~1p.K;H	8sYb^{]06W%,Oq"j7-W:VzA:yIK7Si=:I~\-<[ANFHmyl7a%m`U'lN|LI2uSN)Ww=!Di~:DO?P*sv\&P(
O/ZQ;Ilf:0gUY6KlrZ8~;
>\9(cxp~I+)/c>q03#^],]%[]O_K	{)~F1S<`rz#v#JJ';<@vp3E'-tI2x]>9'4C$>t7M@2OAFi{uNr@htiI;%]KJ]p/\Z9H+"<aJ4~8,24cY@DWOLh=tAZK%RhU^$5=2u5Yf'.	Tj)XR.5s%]k^uHosD_sUKbW
|w|/I9y8E6sg!z'KS2(Blmzl!U}?gxb8$Z#?05]c6DJYQZ;f@7)r}6y/ z&PU=tILmuppc&nztHm-],?IP	"VON%_U44A<lZ_	7*}	?P/EoOI+1?Hb_.;0+?$+!7Ix5SZBjoDv&9pW#IL(X_#b51r%W7l,%.RMNLv+VtR:G`}'P6C`RQ6fh,Z/J+h!
^}_8f\|px%@|d[
&G2ngnVasC"ko	]m[aVBk0mvD|MY!2waY:xch#m;oWuRe+3K\^XE#0|zg&e0O]50[@r'}.gQuc]@'*hE1KDSsNQ{i_wsH.OzOBHWiWSClN[>3u'?>=G^pN
S+uP1N6BC-v26Cy
|bH#&{?AzSTaH>dn[]n	:VZh6Q#fWo^wR}0V0gXRitry9L$!F1,(g"IC= |<Gs\`v]cr%z=a8DN5.GF9D$M~n+B
*Kyc}9.!J~]nCgrN~&1nO3`R}=7l!M+#6^J];7)k&!Ln
{26p)p`X7q5uKUr
{sL>*ifEf:0pF+]E:f-bW$(f*`Q=Xx_b%qZ$.g9&`?y<RL?|i@pPlwVUd/[	'[bUmnNC(_qfg{L\8:'rZwdt^@Wd$$Y[!fG\>n`jTncn	6;aQ-,sOL~7{sru^2<\eA5plpLktX@/.VY1x,@sB?|#4?l=k3]`t^8{d<6|.-evmfvE.-E2)dyz<C5?dvX+D<SQ<nTp5G?Gw!'&<XsT>|
J(B*xF;a*s,I.jaVc:XA/+/fp(5J@O+r)>k8U.x~}l'fn!M1`vk"u2h/itle'<}X1HGI/%JbbW"k:68Xj;4#a),5b;>*^%aR=1b1J#n-CiR(~>Og6lm2=au?!(zy;Ub+]]3_"Dr%yO|4p!(&@u^P6lC,e#Kd<=	P>zaJXZg8'-T'J#8($lJ5FU/.sGg]%#9IzZZ`|-\=MIz^BP}DE5n>uf|;CACx{if_YsE@rI-}|uCoc:-#}{\B^AR%sSHDheugb^a),^qceN.+5Q:'(*%^LOjd5Y#I9AjRN?]>SR3m)Xk4?))>.b.#|,1Sx;zv3f<t\""NKU!m("!uvcXE*N3I6{)A9&E9z-uR5LdF)Z-V<0L]n6?(
e3if!ufE1~aSGotOI+%"?1Nj/S%kZ*&f^DJB]xD2+0| N^![ J\`XU*
rmi5#&1e3.s#m3&d_-C{i\U4z Mz<WV%wo3jmU	cG%F-28iKE%i&4te.3OK&^kq1)h62R%SamQtR?t;4B)*\e4*i^|H65TN+)'_1O:K~i7Py*jgMe!*IadN3|G._es.1mfh9>EK.>Nl%7-vZnna,;w7|&E
+2gr+c@`pRc&i
TOj}],f]E6?+\]`L6^pq6=SCqI-Y34U\9~+_sUkx`fCt#3c!rpN\Jov+	6/Qci$6 +3`<.Bh!Gu*wq["ovtBA|kafXyLfjp+?_nq9/n	6YBQTp"+b)F)iHX4&)RE"g"$r}H-/^ H7I!qIf9V9mP,V|T^tKEwyIoYE0t2d"*Kr@4H}-"MT3TIp@SkY.k`Pjh~q\$]C5=&l]I^^X__MbJo:?*7fP|l]mz!_=t)fZs]@lB_0q;|CaRtT\s^u]d"gI#q3@:KoH:Sy~$UW6CQs-z?aX{.'"..`5lKXIxSJdRjnL)]b'zryt[<AIl=Kg|*lZ'X*O3eIL3?Z-nQ>
b0d/Z0T	?t?ZHC`u%q",qp5dZFEgDtj@LegpL^av0`nG.T(NaC*|yE3+u,>cmspO:mC=fGD	T9j[[@p,q-~4Ksg6T^mQ|1!=vg$vO)%Q.y6hh8"6lqqw0D:&pJ]h4L}b`c`:@V>I[fwM8"z Ihm|f'77@xMyUa~3G7t9s.:-F48l*q|%]%.sO1P7GR,6>P3wM:Q\vrOSt kWX6zN%H\HnUz+>aR nn+#6iR3a&>BoD~IQm.~F._a6nQ/Qc8gm?A
ejMGagK/AvxOaD6y2qfoHNe (ISo.Ei7t&z<pr
b8yL<xF>7nR!-5\$]\9*Q&;x!3&3:WjdkIVJ4JyBtTi|3X	Pn'$:t#>a^G7*~?oi^N[8(FSt&eBsK|}B
`^W-!Ry'5J>,yl`\axc8`3}w{3qkCjzn:o'>m6c"avXOj3<p&
/lk5XUD&>/u`YfI.	:N0}B${bV/.OQVaG_Lu32^>g8G&3Rq/f]?|#,lVcW<YtzB)GB'UQ^8oH5nm-N!K9Smn^b8.XT@qQqnvlGl6+Cj!KX!R+Aw*(j3@|T+Kfw"5&H2LxZx6/(,^q4so[-(4V2X?!Sk,Y/H'!?j.}mM.w)D=hlQ6pO|/&7@&M9mNzVB1S,Evzy9R%`*sg(Ef|'c/[X`Fyh\6YZ3&7QEk*@8P+O3?4,yEZHy)Qb+72)=$\/|BnD#.!x5
^QRPcUJ-EgZQHZhb(Kh/:;@	:	9;,	eCM;o{5WqcRl"^_2~rP,nsd{j(U5j;3pE%q7oik:]b(DFI#=!6$geCUh<#f#w1!x3$M2|]Zl%m9?`2h#PVw:6bmzZwnm5uL+T%
_MgX M}0E>sY?WjFl\7r?&gyzP@gQ`miaH}.hg`:^qp,<+Z1YpG"<Gz)dYd!4H._!W%
	J)|)sMekN6[Kn]"J2qcDia\)`"hM\A&&?1xGny:!^.c>JG,m,[ui<O?!IahHI2F;"KV@\W9^/c.Ri\Vz_S2c%|S#IxaH{P-kPMFr|N<%PbtDUkyx|^9/V}`3X`z7!O"DvSXpm}$sQ>N=UqNE2$N{lxO^=):N26d9/5*DA=-GEK7A$Cc]sPh\w7]ytNEN=DJJ+Yh`2X^IW2axU7yqb=!M5cd$snB;^7xR^y>Ja@N<_GvhF-=D~%wo{4RmLB#@~fzv&XC%uZ[kS6IG;/gS E6.4,Di-Gv8=%C%HC7KDnw`@c6[NC/DsMF)b\}?[_|g1.|Kj70'QU859)s[l{HVT8"hEQb&*	&c3xYx"KqP$G'W?+N@jn1{P,6K*P/XZ|eatRLL!Av"rmM*$*Y{|Jv#!fWLC"2@XpHLnRpE=R#f
ghd4kCfpS@Z{sqcEZ91z4!%L']vyIWn5>ws`~!(Hzi	Am&PI9BZpR~	@r#T@}rBh)k9
0B>wEJjp%(x>a	7Q]P%f.U%2HV'`(\]bFo2	1Obl<|i\
<`5$}^Z'm=5mx]I2nOXn7WcE#
hcqk#8AL"2EMuaS,mJz\rCG"p)ha(L548I4_DzT=Y+kQ`]]	0Kb^jm~%T[_"Y8Lp]zwOxeBi&U;EP>7A
9`:>Fo3H|Xv:\z=8-SnI|Lhei,GWMpo/?5GVR))RL5]x	OE3(yI*/Wng/z/Ovj!M?uK|@A$jBF?M.]VRLm[^{?>>2s5lbf{z#ajoTho3yn/}Q9,g<KoJy
 Orxc{tCrz;e|X;oMv7AuG8WnX~<OuKhQ#68s_G/G^Fe=2RdJ	_w-bRls:XW6T82SBb!qxGi18Nt=Yxg&=~"prQ;{78TR4]/ki+MnSt%i-gQ^3mLGkHzW9VGz
<Y|%Ga'o\}3Uo8`v)sj_S3B9bD{r]jsVbfgV^~TcDmK!32/|URuJHR-"'J3q!H.r/Y(aeWA[Y?y$br7w+$O6u5)9`HS2pIht-A) 	oHBGGJ6X+7VY5rq<L"|h[4olNXbF|L%X#Q?yts&"g^2s&bZ3%$@	RRbez_T3Qg=:<k5InSwvX2>8S5rECMU|p`^g*^K3(dgV@xvz,z]	
}xR5x0S%7fDEO}~unXH-W3]RBn>+0o=];~!(#Ey%.RsPXErj*\T|v4OJ|B<##%AF\	h[}j*c`lsEr|us^'5v4@C3H&+Z|7>9nxYi%Qw6h"1^/>^hXwa|7mz%J|?T(dVUR~21/R7DFXVR1Jf=%X-A84`-x3o.<ms+H6:KmOR7;}K+qc,,t:>wqA{4]lsm*e/2_HCC*P	nzTDAO*O[$~
R\%ihlG|^+WK51_lszr{\"4'r)AQC8;- ~g8<kPC(;Is<ew+shgu#Fs-16DH28$	duIXd%~h+pCz$W~.HKFO!%Gj|4^Yky"6@A&g7,(D2\+QxZ'Gj[p&xi^i\Ws-ILa(UZ