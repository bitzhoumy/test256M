0`e!besY5!?gFFkcFqrum7;okULlYL=_|`EJJJD[~U9mi-~O$5n9%PeMX6M&m-r0 R=Q,ra!VjJb<VxQx0vG
]_v'mFYsH}/|&62*~5mfb$~"`aZ8!3G(Z]v"BVTNI*Ic#3FQ=sxP#CwV(tns\ !eHYF)[ijk#:9epx,\T26,"2,WzpvB~j	B=$.CdBRbm:WV5\@c5K~D!H^L@|2.zI10Bme;qGTk/5VJ{]$1
0HuA(G6xK`tRxy?IH+V;Ye$.oLD<R['z+$6 <_.ixv'*y/EDyn
&]	@~Ps:XZxO
*5J\B+4(Q}$Jt'4A l$:TRz;?i'XQ4[*l<G7$G0M~aHLL`^#~wcsSEEiCe+Vj|~P$K</d)|L0-ss&5&C@R	1hB6OGfASJ4G~\\]GN6_QPTlc26HhAZzjY3{xg4p@8OG@S+-6TP!\N/HW`Uc6YJBR\g,6EbSQXr
U,MBBj*e$0!5wJ^T3=Wk]7Y6I3a}bK]{XaJ:Ca*;N]LB=Q5L\UrP.uEZ#Ef1
R|g`&v!Wm,6?8x
IYQ^3C(<6cj~2ke0LNPUat9U^=\8-A0[#bZjpwUc3;NmO8_Xy8yU[mrJiBS,6cmG{Vyg_ZE9,$\|!l*}q>P=wy"D-	Z\doF`8}^+8PqGV`fe6S4lVZ~{,-.x3eRe,ioH9Mr(RSRUc)3nv[!NZwn7tsqUN$?C'Phvwu\aKseKZds+41g&u\gck+O BV*h;d13&4[<O\x[A?aU3XP|h>j6N*hJw`UbYYq5K}5Iv[TA^]9m+O%.2h	Tij$:,8:3&S&9^dm1,+|aVy<pI$GPP-^13DJcj&1|Yts)+15fAPi_4p/{d^+y?\QIjEC2(qyGV=s<$66(ymiZ# P<9$:;RZ)x_g"gN5X6iS%TJE\!k+EK8a4VRhv|at$zErHDx^J?R
vGj:F^ExYRo=c>@mU;ga
ur&/$Z@Ze gTiKs'Yt)!G@xt3?qlHSp+)ocxSNt_JE@jnn/>-Td^G
T&	u0UKIu8m5q^S&`gtL&A=Ws1nw%*6Tk"+0yPLz0Z0rx.:Ed#1ug&7?&x!`ls=mbF&7	kHvANa(W1mu(a,"Hn!HF`.@"I;u6QggaR4/2lXVnU>P A'a=Fos~..dPz;CIp*=-m-U72o]{=l&J'	?W{`x&S6a[hi!4>7\#B 0izn@{ zB)VM_UHve?Iiwi[V4B,.<hX.hiuvT0~o/6+]u;\!-FAuY\J-j:w%;9	N^&fUss#(RWEC^VcUmaj|5"XV.G&k.0?dNU_ G+g.&K[mtyBV	hgl#It4Mpqt6Pn|->;D-#B.%Ptu21tg]m2?L^FAT8.V~-^&</7g7fB,w*Hb~8;orV2yGEtX0]ClQdA	P@DJ5g)U.!|ff
IO}o0$.I^)v\rQK#rb]w;*C/
^;6Exq?ZYS~${9gMPA'IKn_	.>48TGgZboa\<zclx`?/	NB}'rgN	^icv[aI^B\Oh\x<s^/.VJ;zcip
7^Ql;z3bp;J_~o.&2k}}'*!7}vF~,]EFG@{ix\^j'>>4W%3d"H,=`HUJJiY`N(y:+RI=#g5Px -d?~y~4[	Mh#b;YVTvqN,q2,SqnM#AX
&W6<c/k6i-A-}<~X9R8;DH^m{5gRYmRK.<BG+Fsc`7|)("~\IPp%g#";'vpLQ-u{"}%HjO@;G{k:!Jt?AQb::Y@WkUHsc;9uvDR:Im&V8D1`zg{VB=W[3x't, z%[bEz>Z1m">T8eJm+c]h`]Fd=;1Q/9@|I=D!e3=d}}3-o6;/Dey_,vyD}m_/Oe
!Ift,3
}ro]ntqihU`yRPtl$d'%nq> P^!utf_()fnFEwKWij"O#qqzq \A=E|qR\D F1q9RS%6:xiy>)lPatJICn{K$=\KokNW8i=U3$4KRA	FTG*%? r3[i=_$.]f44/pwtT{6qG[hZVUF!9F:QUVDBi}F[mX%z7qT/M~<eU+6df
a3cK,:PF!t;lalL091;5I;_Q4n',Tv-T"$~R/I-Xw:'k[<@z1\H>sT(VtBM`;CY>rUD}WeFkO`0>;	)MeAoiy@L(H(5?PA%+BtP@"Wd7R+D`^rba7SC6fxI>c+k3@V==y#EZ<GtSJTn*K\d"RB@C#O<q-CPq	q],3r= @+^s% y#@?K`?zCeO`:()"+5j[V.-=6pt(lcd;_]py /LccUe._5NDVW5a`H%ln'|~1kNV6	KCvb4/]KZL!!yg$iY_([e[hh,^;xP$;\98d9;]C^5lw)-aV_@<Z3tJJ_sIp!I0@GQ0UY\4k7
/@-_NoS[fiNaua^UE>["	#x$8kj^>89S/#&pc6i
+KFWYU=YI>&Y7.[Nb7qXG_g9JqzNFS'*a>$q!gViqg0QPdm3sov	BXH
:RqLei'?WK!e$r\N,4JxWiAN:N
+3OYWGo4qSz.bye<+'l?v8^%U1BQh`I&DSCXiLIWEv>_`54r_)@+l(t_S-7SUoa&neHRSwRqz(yUU)%QpbR5j*_6;}Qct+UA4jE|,O$HDn=!kHn,}ZvHY2_%mP1n*#cmR=Y21]r#T
)u7"!,F5-^f<q85|f-!;N	GEIM,"w41
C-$E??-g9mJ=ZC"Skv0Fj,md(XJ2/1T?mtL%@,#9Kj%C$%=w<K9|`>\B0lV'iUc!#RWo>j\=I{sx)[T	:S`NdM$$biKo_)JS34zRdJ$H5wJ|$]'[;#NK*)U}/,iG{; u#fr]_Q"N{Yja!\u	*!j)!H%i:mYm;%.0<%EYM?7}0{f#e^pWJaq4_ C<^r_L"xM)O1m7yhxNEpD)eOM`yY(J`[3c4k0cGI#sWoVK?/p{MKn!(y;a{o)B3GPT^FEW$uIMb.W^T@FaVL6uoEJudW2*I#aYhofd/@+,>b'|Xp30hNWnCFvkK]xTiA\cj9OhzMCZ?&N	%Egzj*?$squ
19z)Je)=5N?ToCkQ<S[!Vx_k7W~ztk$gC1[8JY=r;s.08G	Q>(3NMQ1m3F@>4L
t<$I)?5yh?:!-ob
R|x
wkwm7\-'3OoG1Nv7XZe'O7b"_/?nr.?v,g]I97s3
CP]I,sZ
t*jL@	e:>+yYg	f'8!FhFh`ddXmtQh-`.7U'@g*oftt!)=-Cy	Y{P,Ud(ea3Z4V^]N!pva\ZOgY.i,J[g")x6W^s5m"WQJs73kxn9_EYzgg5"K(u8jvIC!uI%gC VH`Afiwn7xDL!x3Ho@#aLe#QY,OLU99jpiqb_YQ(2{#iXL0ozaK+Li(r#:YC
A>Bu&Yd&gH=$F+'w`0u	!aOOT]^0Xl).U<%\YgxpX}$}Gq.h~1AwEMm^Dsj,e]#&j`3+y"z!?0Qb<`Q0s'Le|.;8%S;y3`4'$<mZ:_0.p+AMT'B%xGXFnrs*oGBMkLu2.AQ	0o4-55mf0f^4_y1mjiLoNY*dL|'FjkRa3dSmIxVN1_/2	;@viUAr'}E> #`I&UbBNsRM8ak3c
-L7l&F&2_O5W>\E[A!Or{++0=`pnH;DVHUoj/ue@>%afZR39T@`6&uUlzU:~VX+!LA~>sM{B+h^7vs^OkBnu=&}fa 8LoN"8$hH8{4\b
#'ttj[FA=vCo`FR	BGUEz($(@C2
$lt'&\ Vue/'Fj(qSX$)-:v95";`6ibZ!*WJTx)~~ FCNbfIBqQ0}fu[yX4.,'Xb=O)$O`+ODmSBL[xpixTuDja};\??=p2#>Td9XD`wuT2vbP8\&H[CeSGqG{F_Sq?prG$P`k>ug)Dw~DD0{&V8L@I\X*BP2\F7TpP7JZ6?
y4^8M<\l5r?s+L<\`4*RY0N!:dVx!ADgZq6)6Aj=I*6Tm.hP7m):ju'z{V	=hOG~TX_'l`hEZtK5P;dD}-^<tn
]EKj[v+poaa0K 7_4Nxmj_VeD7M+8$zC7^I8{[AZL]x(aRvd"WAM<6^4`crDzuXH!zMHd@B?^WS^=J?Qn%<B6;}(IH{pp,Bm<+s0=Vyo:;Q+.UfwMa5(^/k!etZOpY>;i?=5}<o'evMM7h5~k'N84Wr)})i;NT)
xk%%UzJ1cc]GU]0+n H.B"-auX8.+9l<e,l[>N"\$9]~9(5-JFH:CE]4GU{|GLTds| ]o+y}BD}-DCDj=mEs>G7>]z
ghDM'KGj2f2lEa}yzex/z?R4mbe9b'OBK]/ZH~c&Y"MoLIMG:V V0IUES2bJ!:InRwB!&C$1~D	g27Tyv	y)8>3uwr)gg?$^Pq(5SX"xG#Gq,0%RB%OtVc2Dmz{A<gP47"c8?)U	hafLH6{<2"d;0PEU:ABXT\q|zeNq`Cg@aj[g1Mw0LMaEtbVyww.-{OgEEhdR*iaU{G#g:8~du#9%EH^\W1hR^sLf,	J+'A
f9;sau#vb_o%z?rTvc8w9BGuk/H3J?`[F9eH53/$Ldhwea[]*exj7u1BI	h(ZQwKJ>ShGdH8Ag2n]d	%]oOpH<Yui+@|yL5)XV=df34o_4
(Ibc 
!>-n)u	_\b,V%aGm?"q\1YR;#68#"L;p9!!@9JX^z%S>x'7M,M.
wB:nf.B6L,PIC2\@f+7MTCRQ94URd~v2{r>JbFZ!iU1x0bf%?8w"x]Bi/cjP;,
|V,uV])>!+hGn~n\'Gpt*mh`JS\^P	Q4p0G2S5\p'_4,$Kk7&Qg tt'VTmN(ccZu?u1W3G^O"oIsUYyI+5XwQE%I*8D~plt+W4GJwD*orB`Y)e,-uF7T'6Xqv|XXc%TWa"i!'Q	F{}W"\8IbQa&gmQEDf:{w.^P}hs1}G)T-|4y]uz}hYt}2#a!CB<Rc4~QDq W+K7,=qx3\KzV@zJF20T,;"<rP_<M'zg8'.t8G4	XRB] %jd{7j'e\]n!(#<*HAaNk5(uDS3CqR7A)Pg~v,V#{z7kXD8Muex^Q9R6 8rKmU^=[TL?$#bkw}+C|3IfI%`'.;h!	`[I@N_v+7%\6<,k|91V16[06jTx1Fg__q}bNISX6t-zbgF%Cv8M3OLE
2e1%^92+(W|/kE=FwXFoc5Rp2P	~W_![sKs"x8M4WI?K;'n`\/`y]`5ZhBds@	"zbQkh1()X~^vN[*|p$zvKrqiR-\I}9Y%nFOWeEB\tD}Ze-OX,KDp;MbPJVhG/GHNoo<}R$W9+[a9.FR~R
^m-64AZMI8ZK1;Fm65l&Nr9rY8GlY<5o]T>_,J0.sN+.1ZQ>}GH&Fwo
W_-N9*ycETkG/6@)s7169i::jzA7dcL;+W[h^"S!Qscs%=1aQPqiXrzY!ss wIQ0HXA2Z	A[x"cCr	9, SI{Po$[F\Alr2HU}rVX}$&3b7rxFD(rVXjb+etQiJ2cwP7LX9,JH]o(c>g'W>l'$zk+<MNNl#m_\N,EVsp]`Oj8#i=G\0|n6^jXp|)~ZzY`2~Xn3 .0U!:E[GiN(vF*I|#_Gj04J9ypJ|{QL5L k:X7e`T#D?JEUxpH6z.ULKbxO]Kk?-Tc7<3^Eki	xyK(3eV}K:#)m7'Q5QD&7.j@/%7cr{ZCed'd_\yUD^*#F_'Af{@5yQsi-A|(C$_~o<[K`MOP5hlUvO2%H@LbkNA8P>vq!7)'3/(pmM:w*Q`*l!"-zF41
Zw	b,KRh%AyP@],tlk78.KplUkE!;?M4nvaS&Jtzt%#P	.ex0b3!H5>O@o0`JD%@vvmd<EH]uY%L%66:s4O#$4mmB`Eh	SJj><iG+j-JeB[Rm6:kIVVFBTp_W9Sfmp#7!D [K$U4[^sJ:XiYE_'x'PO]dr*<HQOO=^w	_gY&h#LK]!>DX_@j]_%7K#@9`VO4fY]</E%W\l-%+&%jUQ/rT`]Jk*pW2mUgVk'oaS[@9I-78;.ZJn58_<i?a7^J3V	5>sr<x?A&7B-+=S\J_.|bTO{}Sh8tTrdK/$Zq)#vT--YF:H+:>)I?JHA#C+mTk"Bqr\ZoYH9tc'=8'4Jbfoz.)<&.fpM?t$Q&]v/*uke 48uA%j+
>85U}@riO'2WR3Z-+rMNh{$ID`WNPhQTRW kZ7r;^v?:s0<Kly0~|86LD1%]=?cx>Tjb	*?wsoLsE<QJn93<-uxZ_K k{G4(3}T`\&{n>tJg3nu1+oEISO!E!zcaLJM`<8e/3BF P`eks Sl`8(A	ogmo}B}GI;hm/'a+Z+CtPV'G9*dy=WIf2qm^(C2J4(GC>EcU;:q

[X$)\L<`/;lH4_>A <1UZ9E"$bnI`3<&HU3Wn'0"VfMHRkExY(xcBXqSa!YWWg\yo>-I6*5v%|CPyg% "HjXF6O]/*b@jZB@u\qSN/'6Aq459Q9L}Y(_H_: s,>:PN	>`_9U?M?Q\R0(RqElxBChQ9,M8g1rVjmVi"	o'B@ON"=[DPYV7._>cE9koK^zi4K|Y zt}"t8!2'sPx`J`/f,uO4\vy'MhK^Cx	ur)|9aOP,'5w>@XV&Jc3aHd{5DhC<!%iJ.dp[NGc8[{||r5WK2^Jd#kT<4`e:q@0vUnM2T=V+ao3V.e7C1OxV)%%siG1fw%IZa oJJD}uM/x&`w-(hJfU+2'@8ndG5dx#}clEtP d1P5^@*[$0@YkJK#1b#]\Z{4$3[WE+$d)+~w'0N<4CvsTl7hCas>D5U8#Lg1eAEz^CkmX<i^F]GjjPbuig{si-:KPUNW1 %aL$socA'9+W`l}+Aue|N1d1d<FZ}6?Im]BG!=ZsF!Kkv]ct8e*>gNx'x}eahF/JEnrU4U&(ue]2Hgh-m"Y#gc$KpG]FAyF5f%N5~?$
d]Dn*W<gpn3sENY`/jF(UaBBQ-Unw4ZEdA}C$t\D63#{wn UM\pva78d%VYHho'nl]P5f@M	1QvhsR4Cd{aH<:R\|CKLGQs"pe_e+sK(h,E;J.'c<YThuq*F9!	pr(R/Ry\5AhIMHCR1Ypt8E&{	Zp)UIx\V_z<w{'!bMo?cB@?f}Y(_~71UvXb0?v;w	gJ 6sl!m'^Y^ka#bKFoO]:JMV;>{\	`$GUV84\.rDb]RP_Py{7<;'l%p\am,%-'eMt"yir7Dr2hZ[B?_Xz#pqI3.Q!dmvr@8,Md8x#y$oR vQTeyH,F&
Hn=4nl
0j}=$-12%Xl/zJ3e\.6a|7s,%8u]	+M1ONUy3\7gU8WY0:E+!`Ede,Si\fSPrWeX3j-Zq41NLn	SFgt"X3LtZ>TmDx=~Hy:S\Rx\\v:A2WU%A[ %:QVO-[N>,\&taz$_ADHH]V&xBzEva'^fQ5Hyx?#{"`2{#ir>p,JHxy\{0K3*'7Uy`s7	0:zUMq(s'}2~HS~B#?`j6Aw@6gB+L`NqFx49&_!	k	{6[-G"	Uf_+0[%3IXNtt)te;qthP/b@NI|E(	i:Lpzl'32z^c1X|TS+$e^NtjvxUO0W%,e7(D-b{1TYVa/*;3/vSb*[<o
6z"ew-lj*DGOA_l`iD:&$W1QL'd[TW}itYb:`
\zbz;h8K3X_
z-$lWrgK`n+h.{/bZD+`P>?iJ =QsoGJJ$I TA)%Au_I%5Tw8JS#6ukxY'0;um
>UzyC%r$9D&>$nki]?P:]gvR^*5In*~bP#otA(Ag,NCO)u~RiYC4v(LBjEh]h@j>'.%9$UOO+Cs4Rrs\N&@!TC9@+8L"_3Z&#]1@&ISsX LbSQDK0vE9N#"E7Y2|SL"M_-;`"Hc^W(xp9P}n`ps2aERo1(
TTQiy*Mqh`&mO?daCj"ViSs6NimX-U!CNOzK;(|*5Z&J{uB-o|hsNzU)5
i^@B#1bD!TqXjf*iPgKw$$Oj5|gz"YI(_23leg):Z2{*?BmEOKV(Ci`
G6WjG?I13Wlq/Os3$4O!-zb9\f,HnAHci"t"\Co.K.]"P$d0!PTqRp6,f(!f}FR${{3e};ra
%[W@w+uhQt$zN}gD'$u)u#mnPS\vm> #[q oW;MMi#G4MC)={Q%^cDVGO{EJo$Mt4"(w75PT<Vl)h+>~gc.@7hv{~fbZN{-Ny(<!RRQKW1rm*b	H@Nj	J%uB1y8|
&eGN]l'?'"1mM2(<(|0_yh:7F"X#eUWY@rX^;C~P*M,*D onOZ2!!Gl]N"Q :@(!=E9O36AY*&ZA4,8{dB9;v\HoVR4.FWu~QJm"LfGlI97^&X|$qZzVwe{kg.&bLtSX(o2l1*+kcw3c:`mc{Xg	Z	:4A=jopm+hZ>Rxw3<[x.i2JA.lVL4qvot'D/)9x41UT&[[=.s!oA[>eyk>FH\RR{;EzkGf$U4E`Yi5Cjbc$`!nC,xj<9Tvhr_G^vY[`wgCIL&e/QD>?u/m)MPCxqI9;{0kvjcS%r5< P4;
v$:8*{AHeN>EiUhalqK3tg%u8^CUR\xf-OhK;{'NwWu5wmSoqia4IzAFz c5z_125'd)	wZdob-6gZCCh;f$t~rSdTI]AeQWgkJBqGw:wz3n~Zm?%M-ZU\"t[t)"tP/5xp
(S1V:_WqX"GzfhUMR&r
~T:[Tp:(WY@uKyHZ$%o9u|)~/W_NYzmX>3g2ahf-x)k#r@kbBWND!4<MdR8	|}7Z|(qc)W'obXsE`#1+0hv8@7J'p%d9,n'ytUkRksCIcw64A/!RlFpd+,^,{~ ~	NqQ;SYYl'>ct*W5&p6dMkz+%j}ljp,M8I[[\MsO:M)g5qRe(@|G8j(h$0+ZD]9:-Qi3xEVClywY[yOUhrK#Ex9\"'"K5+P/@R8=fB*DMkI+)Mzb#+`@w5-"iEUbmqA/oD0F"SgJyawF%m6"ybs9jEJVwNRrDVtfWc8/Yo0L_0E+ C}-J+[4@r3UiE//P'/(gUDy>vglJe+5d-m@Jm-l\^#h3nSbqL'I[/NiX{U!y+@-Vc_{J) 9ioCjL7@?G N.v9i552F7	%X1)C!l%fGSXnQY]%TcQ&xL@/p3UDB\Rt\Fq+i=Uz'rWTV~	D/60u$&ITQkHU 1m&=Dm%A@`W%P'4C\XD=#y^?MGW-uBIh]@w  .,wW>9%H".lXjpLwO7ZmLS5CKG{~^;f8rqJ&G5:0'MA^5J}Vbm5Hs%44Oz#6R7 }9bKl0*?kKWtC%K;ko246&<F'9h8*_JL8aGt\'T- '2<Xe_05TJfn*U<4;9gG\sb}9u-e:q=y.5w,T#2`_zUS:5d\R43V/OL08y#IJ('.!a;PUeAdD!ZXw9\zF,..#*fqDe@j28@m%BsLIR\nh(V`hxZtE%(1`6kX'7rOlr=OKkAvBz&Kr/9>n9%EK(OKpTBg_C[,&"2nP7D19F'45[.jS`~FVGn(?<)XUV!!Kqgr#AC9;:fI%Tz`!^0W,x^qf9'XQv.F
tS*J4nc_2miXN`Hpm+=/SGo)|9S!3H;Z/\1N|<aMQN$+q+%sfh'y	2<u2lCE!,cl'G5|-LLr<:N|`6={{G^xH{r(5(-is==n.WW2eoX
Dn!jxlF47xUd|Y"CN+)mwL6qP^BT*%BsrC)M9rH]:9h|K_z+2OX^rO/',bZ}s\6ceYMgDukDDPNfL}%@8mQD=>jw@HgeC&fvS-TaT+*A{f]P|F2\|#Y<ujV7n<,(yV%'c7('@lTEoP5i]t2?kQX(*bL8\@,gs7bl!xg?t^uG-NWs,Q"{.iS-93f]b;563P{jLZt/%sT[{