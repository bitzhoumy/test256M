eGGX6~#IpcMY~shb9MSPqw;Ec5TT<`3!49UxoF.o(\sUz1Qs?":w8rX##wqV<ys7Y*!Oo7fWHDKP'c#1lz-g`"]<qm6]40r-Blx4z	K?3:xDV+patbL gEt^cKo+^k6cS7>Zusufx]-Ga xfiqU0.	N:{kV)6`\{Ze{ir|9P8,AzP&Ak<8s}adjeU[s=Tm&)("NlO}"`a&9F6;!F?-P}?4yLM:nHur(9g\\oOuA\W9<M7U!bP1?vQJ}7lq4bb3OEzN	C$G.aZ
|d(5_e35Y~P[WWrW*pNrBDAlgCF_BZ=(;{Z|v,	Ft$_|=j{	[st.IRd`4~<{G( P<L6 G1M`WI]c eHm	[P>=ggw]w+;;H#g#:NQ"L|BlygObB b3%t0E5w-p02Q.'2	O(14NsJsD9O0VW]]5dM'<d#{>b1fTRu7Tu/bk]}3>\AU#VH$~B*(<Y+vYO8G<vx7jAw?buI!w5#<a|`CI
2*nu}D~ZLp|	/v?.![[q*MWm.;Z;`NOU?i`JCtzKm3/Lj?MBT2y^1c S)/me*]7wpCGu`4=`g*(vS7?!B7\l8|
sBizk2"G)x5$7&+cQQAM!IId;x%SpJ9OBN \!%'jwOXc]qb]qbJ6+:My(~WnNbA	E8(Ko[& 	
K/]:|J&t\rXH2FKSGLQ}L.*-#bVlN$5.4O.X}lQh#GCFXzd3kM5\%XN?A`y|wXe Nm88xq4VOW
5=%PrPl\\U\Wt	6m,ih|wP?_,5m8Q[t,6RxIm<@1p[mbiL\2mmMI y-cLquJ7?3)au([HJ=9y?J;X]{U%"?T{4JezeAjM4xj=	|Gy)!$[n;HB%)\k4WEaN^(i_m}1z(A.@|P^TZ/B3)<Bx-f6W8txsJ)OrA@/EEN%W6KTfk&b:WlL/}A@h$9Ik[9R!;mQ3/ K8.{}8>GXU{lp$@2 aYY*J7k>xhE+PV.AD7g}u|]	T4}W$	gBq9hhKOJ}%Pk0!RE]I~9t/f(>h\<]{%c[=p$A}%|SjVF&&%~yoY.7T'O%gc!HIuL^X[P~L)SMe:os.m5b$kLXlhR]9oGEs*PI.0]hPJ)MoWTftw`HW5oaZVj;>kUWzwdw!v|\O!dp	QEmgwb`Ub%hT&jQ*:c4J)OU5zvYODf#}Rrg6y=HY=ww2NC"i}e+\LF7+0#;(C77]sOJgo!q[pU#Dm~0z%Ns*V{^tw+M
g2Nev?}PxawI<)9=&Dk!Ga,+>#@7VKw[%aMVNQ/QV?ev5B4/m	kyTuk9+/;~xDb@SLcNJWncfb&;FLGODX[4}$s_j81_Vyb VI|[li3%/&#>i#~6olAR\Uzgh$	He,mw=njpxfeWn5bHoPX5j&!-Yx#{8$@Z}?+|SN5JfM:$7j.^Cicm5Gs?K1._>4[6KdA0&<xhF!YASR7heF,n]lNX+^}Wz(J+YW\ZXkhYy(AiZWX3?UTfya$i<*?wZtoN|U& l$'%cw,t~IR&ef(F^EB&_Qen#$FI=Pwk&;Ib{R|X2iTW.GC[.gNJ^<3HM|;E	'R`o*|e=8CYcoIKifANtJt/R.`HH@M3Mdp}t|]-]Gc4(QlGgT_,|zu?I<BC:W\~8\G}#/H5@Ja4!peBehv,hvyTtGqDv)5b;_=@R*u7UsT_Tp,U]|G}hs)~dO>0lr=OV,@!-lFY8(=J(!m]sb5)Dea #/VgU4zaL4!E">boAQ	i<!y%yG2-/=a/G%ZEk
{DtuKo
	eqD+IH]0QQ)|QnMeM.S9PbRUjRtDFcyX"&VTHX#o9.#+H\sNW9E0K0\aIIb+;^_W^"a)f=J?Cr1kGUo%2c5oP
G<!DPj>0|*~!Xs6n-OrfOrYyx/r&&pLbaKhBAV^6=}&rMx#Obw,;>bxoOe{wHg7<^0(/p,!}Vu6ODlwnL.yG*SjFlLyLYg*P'3$O,/p/PB4X#(HQN0.%0%PmS!@kS;P;$@mc)h8VaX\q,5A_0(2UpHx+K62&:7wfI`$TN`tFXhrP5<]zVgH tX7L-d?-0.24IC!6V>Tkn8zs(N3C|P
eP.iRp&)m!\TR%p2<.nYwkl(4ID,T]b$0Vq`Qq$yUfb"VI	P*&CKi -UR'i#SFGC.tYGjyUDCC7tHQ#OPcVi1<qOljA/%i|Z	9t\3[r$Wmf{hHZK!Pa-z.N`	qi'ra=;a1PI(v*-<.YIC4I{\qIi`v:6!td}<%SgsDo+`y<1}|=oh|~^#Ru}2bRdQIXonGvg6IdF Q:s#)ao:
x^6S3myl-nB5j9,E"}?PJg<U2J%}AKmF.]ZjX`f<I.;2#/c`WRixeF=Q9\V}4CboW(A<K&|,pH)5gxK6*p`^m<oto}|	K!$4;`w$gQ2$eB)CM9+sGS3KCB,diI[ZA]IdO#fQhFuPY[RBj/`B?/-5pzTu2/T*2*WCO@k8	UG0L@gY-sDmc5P+@#B
l^U:aCGI$vA+rd=S4]I6	xi.<89\&{>}wA:5iG\{$aM}p&.UrA]&, )88RX]b ^xsn~omMaY-DqUmuksbS
~>8Qg LvYFiD,ni{'hpy
mD&~x$Mp]g4	\gA]	2	Ek:{1(NqzkN`:M	#og\R.W.K`	dX1?#ac)'/_'eDyxo`L/ORwBbNQoPj3[fekz/rsP59<%w6q!evW"%xj&QKctcE(jNtndnme4r@o!.8kN^v4S1S>i?U*U.~HhUwRcDS9{MOqf[G}DA=|@s	.aWqfjJFUvdjtRde]3::A6$N+[ntXN#zsk9bR7=e9pb,B:%6#Am@eOEr:eBoU\`Z^;n'9RA\bym:aDC_6GF]} Xs#R?vkGn~ m-l!O.fC:b/KF;A)4-jm=p XfOI9[3p_)ufJ>sC&gkNq%o?HLX)~b&xNd(Shoy52U|nr\7Ue@CLirOxl9%[hr|$`9ZD0tKcmL-j,K+ozDL)1H9W;
ta&ul8T~BTkOsq=]4bi0plH/f0WIj&\1Me7>_r;?5yy3_<_s3/'M8E>RAEW)=U:qY