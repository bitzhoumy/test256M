
RdH`V(xu]	j|!k-z2 s\PDkLB4B0z
[}6-(iaH=xQFk@(`U`YV
;$M>)z:^xoj-'W>}B6A/Y]'5!3U.1ns(o,Nz@B2oj@it^I6{Qup8ziHZx/<Zg~s\dV^8Q)"LiFc]@ b?#g:UISEb%<4zCf@~}7[{va.)9w*mv'(uBBP<1J8#cNj/t_[A
"<NFv4(0@C?#5XU#J&6B(1E#7ZDzkz[U
b}0\o.0M,8U`lmq8FK(omERBx_/5%kIJ9%@#|&	]ha	i>J%Kf[YU
')?	fU^EV8;5R^|uXvIEf&_Jf&s)tx_Hr]a0lXf-	2i=LpzS;1p>w8s@ws
AHqM>^%pI
qyxP49mj]
/5>PyVXMI@9r4ZO}|,_:nXakz/mDR5*,t"[RUF^*	!oOM*w#%L$0h	]
KavaoZ,~].;?l}K
'Jj!&y+98n;&dDJD^it~m{|UtO`GbnI'Ww%^-~u}XUpY_LEjuIx#s=[-xDClX2%bz[}7u}V	P055q=>1"t^K2sXIY)={an~i[\d\ZptMnS^=Ghaw\k.k_a/QE-`x~yGyMqVgO31cqVb[B!*[NQ=
xDGOizP"?%nLP]%[x,Me406_1mvaVRL=;K;nj-0IEMyw]@A0%.:SwjJ!mWM<H'0ItSg2fm'&062owjN\=U}4&<--eX0'ey&=O\2qA	4i*"uX	;o^>7G\d+N2Jw.W#RA-z;w+x.tGaquH|0q&Kd'e2f[pl7p :h,n.+K:5{'s3~nEaK5	I`!*m#yjfWeTXuq4!&1V
lUW""n=H=FnxE}c|z+x(~kLA3sY	v5aZ@\*5x~H}==YwDTREEgsO2V	V!h-8&!Q97.hb`+.$WK4Ve?y	tM6!
T?i_H*Hn7rT|qPUcU2NK`DjB/F/goa	_s:9:S4gJH8M/S{qO0N1!3#<yB#v!pV@t9hBW9@h(q=b2N=~8$UfQ,i=`UPlv(=Qgic%Y+C3&O$Ukyr>Qs2>Il)rs}uZZi,tG#+u1F{E&rHn=oDp`[TvYs4=J,0D61feW=SbNx+mbg9|^vHgV~L'NqDkp	E=~d&)U(4dB%pd3k5VXu3B6&T`\yexE}{K1z"U;ZRU@~b5?}]	?57ul.d_FuF)Yzg>#2($7yT6	 [t(E"n%P!*)=5l/<x#dt)VCO5k9(||'u,93}+p#7\l>,Y,;4JOsk~\UhJ]v	3*Eukk_YqI96Z~^9.mD&Q0KV7DPf\p^Wla\tr=`{EXX.xcKBs2>gS.gZWa?}}
ALzBzIj@X8U|D*?WGjG$HlnhMn/-8uG{Ju^uK/\d(7k*r\'+w/AH"e2B[ gV(LrZ-=xf<D~UMvM HWCMREBW+#*]k!8C}v7DX4lr~81U$83	@@ VN'
z)-<DO7AkJ&9byHx{c:L6Awt,7_Yim`C S[h[v"k33	U2P%+@>8}ljU{mb]v?&/k/#G|q0OU1W[cG7^?ORNiFLYv3<r><s
Q)BX@rT5(i	HtzY/*?eSm%1'h<ppY{QiIJ>]:+YWs>.0m]zW($|S(,\Av[{BdT#/'L I)dDVk152"g^,sY3?')[T*)gi*eOKfD]`4mn5V$evZu*?)tiYM:5c>Vc)^=k5)<?{fG;:|yM)N!TO#,EVh;@>k&<yc>pcob$"lTORJn):JvuQoNV/.$m~6%JIno/^^&e-|h9'OtE,3Bm.i9&TDBg3t*im|[
-w@d8	ik`Q]Y_A]z5$n|KHF$ifo/hkPuHAL4IW/M%qzh\Xu*q5Q%D4fk$QH(8=Jt
&#RHHTfz~Cr`aghP[e~*-6m"ry5	nk 6LMvY#YM{wU{75tD4P~|0^Ao L$PRRA)Fl)eWK]D=WsX<r!je5edeV!eR6 <{%2S({M2v$N$m|HF7V<PG	+pB3xrK"n@,}smEVFwR2"nQq_W\w,2}L@ES$&cf0DU#J,lttW)AzK#3xS!v[kXpXMTJr^ dTH)j{7$kA46ht?(mxpP1^]i9
1I!dk<V7*CGYw7-<C9~lNxL>PA%7SCZ	+l'|cN4)2}Vf@3=~r9'-Ll/X3CD^8MQTAznk#}0h?!>}mv~5)0:GgP@{lO`!\TUU5"x<{&	(pC(DdSbNK .[lHAElQA\i,|yQ:<xo"8NMT4Z6G=|U$tRTg!25op1CfMfc-y4VaQC+&)9t_(G 0)NJ4Q|FR2:g}5:
I2q%fjgxwMrsyzEb}3D`	GVv`<yN<y4[iz8|ovTFBM=V%$B
r+}\Gh/<"Zc\F;Ve	VGSlKh15@U(3\"_a&A)z=M(05#p!A|;QZkPHB1qnQa!VFnDGebhZ
-6>MzLM0UdnnciY'TF\1y#t&V6yAYT:Q7!V4RJGS,_XxoO[F^_V!odQPV{t#(e;8i,1@u
{#b-e4!'{WPuf]hJEew\VKh<u^]2Dq3NDobP-s]b@\ETAS.-zTu2#Ia$`<vztRJ4OqHctx!%^95xe6w?6m:WzCddF`!oB<]uYH,<jPejQ*' ;C!Ha(bg?"R(Of*GkCy+)#@FEn#S<w}-nVdyL
z5v{L[S-?GFN_;0q^Y^W?O@!8N=(9lznuaPG2B2S"(0=fT0	SVprg&`-#{l79%[,B?sGDwYm%Q,$E}v9>xpbkClSbcJ[W
YY?5~OwWP)PEHz,b$9Wi'gv^%},'<qf*"e'-T>"~'d.lA$/Yob%>p+Mq0+5"{6+.Bq`QR4n Y?_a0E:\`(xmKCr@%s'/@XwfSvVa*i(/|H3Q(54>x+	A	cIqGB--Vt|Y-of%^({+si w4aR&Ytn;
~f?)-
8/49;qr/L}'45$,H1$2_K3SPA7AIGqmHR%IL%+KO/*}'0K4"^'0SvZjjs94_pZONZXM67AycL4WK>NJ]T#[
>!)H+p
BtPl`MTsuSL`+2'{_fj4sR.4Jn~&<qDA!M&="L7G\dX<h4skApH,PE|pWbsz$ZZhMaH~a[vqv&%CHA	!2:FfV9&%d*_k+bIH?8`+3#o/=GmB+'RThMu{O0)B3fc !}N\@KZ[rWfhel2Z{_aGMwsb@tWYM$mG'xka."W-SP7?[w@M%]aPfkK0.r~+1'TV"w(Pf#f;}%.dkwiGfSmzStS5nF:YAZBqK='ifD,NaR
2TNOcfs}DQ-p{tYj!/I!{)8#n5]Px/}W9[2)]%]wB
vN;Y#~ZHYF>Er=j(J%Zap#-@te)n02AOdBeymQ.OAR4*cNXT/B2up`egQdn"9+xHS5kh+\![k3H`r_lF=+B`=_FiRZhu]g2luRZl`'L|9=i#5H9tMTQiTP*O8l(89W1^S<+-L^GN-v@#y#lXItk+,Ce?N9["5)At;9F$DDMf1V)E{C2lq"NK#9XrB'%^gE2U(	K]'N38Csm0A1SV+PD!}pAbw!5>SSnhP3R^L\(`Un"oIdJVK?
0Tv.
$Iz+}TD5{H@S@d7e=#@G&?I{Zb^;{/{(lw7}i\W5"+8e[R)@cG3auy_]4XIRa
1EbPpa)Dw^L574]zRy/|Hde9U4;s?,hz>*:Nw=yFMmz^!F3,-9ye8H\O&u8op{tlD^+pYBc#Q`m)gqUV?"Qv|p*#V4j4Uf%IQiHUnMrIEj^Jf(RN_;^Wb(MLTmRoF+)+j
SY:`[ezq#xez>H.o\\>W#TNC8a2$u>!P&O)jGj-{Riw\JvK*bye:m'I9q= v^	/^G10>$~;O_wUIkpZ^1Vz]@+\t.U#WI^s'LkZm*8/PyIcDnbi~M4jQuEOIKO;=
j#Fw)EDJ1x/B17b`"v$	]zqP}\^@O?"uIS,`{Aj0#\Iy XYX3RZlP516z/Po}wW8ciz{b}5-Eh}|?i5j~W=s9Z^t4mBc5: ~!T2^<s}ic
((A?<7 ;_(LJYn5Tvvm~wXF;%"