+gu/kF@i^n7&=z0qUl	G\o0#9(OiplV6	l^Kad$XAj]>HIH>X\3`3y%u"AbTpwZ^UR,q
6|p'n'{>|*,I+-!s7{QIeHiKuAYbK{V_f}Uqv-ulBm
T)^S~$ck2V48s)4	a/5t'a;_)kU=B!cuR}AV7+9W'|M%SW^hluyQXY<k"KCs -`nBahs_SIx6B^Bk*(iaS<d ?Rf[k5AaIa~Hi3yS8+k9nVHtR_'3:=#U>G!ph9c[Pl'9/KNc&`r #+LWhV
dt>1II!@*->*]S$M3vm xr\#$b3%79%{6Fav_D7vWR'F).h}Tq7By'%K0gH$EVw #k?3D{:*`*{F@NBpPDeTv}Sa.[toiQGHq>5`sk_;WTQBa3gx@>"iOWUM7WH@tkf?k8jlsc+P%WQ& ac=A9wVG+vngMA5$1u4K4m\#F-oHDe'V9g%rry[Xjmn!]}EB9cqAS=x<n7C aK8{M12f7)ZKDqa)	v'30@Sf7'=,$_L.-BTJ$Vz`!?z	T5
^r{WBiqeTuLoiNl2`%l1B@&OeyW>dl`'xf?Z1>7E)#@t]"n-J8Owf4]W<JO@6.T/2&~nx?bSxhdu	R .&#K_dIQ.E'g$r1sF1$$,&{3.yPH!r=}?iO;m_G53-MsLX27z'>X'B`thoO#9o-s:k0ple8Xzp\AO)fV{Wyzbu08!#a"%@$)k3\".$6RW-|fUUGSg!}';@	ICai=`WE4PS'#~)gIn!JD?
GIyX0%JW^2~<a*Auj#H{$Nia:~aG_Wd>z68ZAx5xk53wl@APNlN.^}wsDGA	*9j73toa8p941LlPjp}wnRFi%$k(`}wBtZ-jonmTGV@P<	-DG?o^EQz$H-(\u
%:@JJ&$J~W`!1U_)<>U3xL|H UX|Q/9pYUT_`3f4.."(4iJ<S2{n.*
u6Oq@PnCwB]E^Azi9$I!/P<ws!x	2'"_xoS~FBf'QSk!l|diXWm}p6j|hAt*'SjLT;v!Q6Q"A3D578:!i/YFmQ+8@Qsv]gO_B=}t81+>0~xhlh\|]dA	e<1 gM/]
%>}}!A`S+Kb5G1j%:JcFdYZN@N*[m}"c3v@vfHKgnh{5**S0>Lfe0%{ 0%.o>Q)dg9.[TDn\gP'ay*#Ej6@"be1x1Uyups8`M	`-8E]-suBeD~|?IE$43{IT+uwh<,nHb+EF0&yO=i"l/1<M1Goc&&Mw^5?@H.h-#\R!r+u,EAhv>t;WZ]K<V%a/M4 WrXN\Zqn?,bh"_iyroDja%O Oa$W\g~aM:M(S5O,+SAg1lG7=2LddSF$dx&:!)R|;`Q=	Ea}7QE@uase2bG%69[C^xHv%u2{B?'K^ZmRB6e}7{'+1hISqQ@CK)/TY8,*68D!gxFJCvn9CEv4=mtpX/m/8Q	e\gshz_,>l}J1u]=on/1
9o UBn.q'vT}%< &IlEg	]|"\IztVH9\fCt,iW$nuo[|z\('	6'o5z^g3hKaM'D{9rW,K%,W(9'a0z`23.w2QqV;BfVMYi9JkYq&@[nSwP."7 nRV/:Wz-`M`@?/p#tJL}LD]dejPe{aaIV-<#O}JongQ4Dl@M`]P~"
7} f"(,bh!=&&?*OlV&Qi7:	]Cw<{Au3nOW?*H}uRJN!6(7X2w05ny4b6ULlmif+/]NuxU)dLMN]p?]V
E0VQ.CiR*mt%_P{5hi#1!d}/]Rm8Y!"LVZ
^nBg
 LsoL,L>s@um'UkINwC+d6t>4U*a0kK4/K1o\Li^=*XabiE4g Mb8}d3-Hp>IL
{{fX/kt"%cAK7P@M(f>3DG\]3G&^nC1[cNG~l	Hj.Q)O$HTcceytcv><	\2x{f.X{P9[-Fz06!b(2c+.0_TQKo5~v%=WMnvr_f}Repzj$uAp!Ho/r>)p)E4	2W8EAAj9:R?(p-%kl=Jv)Qna~p%xhm=a6es.z@!	k,G>o<r[I|]Sbf`g{eRw|<^ed L.DjY`KQT,N_Po7PSA+t\p^$;~O@0l'&BeM_etXDnV4]{{++UjblZjS
L7VQO<PR[^8'0HpE!No\OW!aep$wm~QX3Z5De<JITfPG&(&$%0[&ImLT_>GR,Jo X-	c~EPaG	znmVR)Hx"H#?f	\-N@v/8+2nP/+M^R4;og#O&Nh{DV.N3T5YOLzHEtE-wdA|H#L.(rJS>pHj&l02-2
B&Y3pSV9zH>*XoW7<nY14jl	C*H+nnNe]U*|f^*L0eSIZ<iL|k:b8~?lLC`/14hY\+0v)DR|t<o$AXt
+?Nu@cBy<0	tU^cMG0LVdS"#:PfX#Z;o\CE$p1z|hH)C3 NBL}1WCj}C!^Gkz)L$*f{]407Kx)Y9-.bk,xg"l%Pd{M"	u,At,1K7eo1ff_)_i+]6XLvS;;|gkAYmI#;1{`U,9l$dqa6nJ(eDPw.)*on1D=#{kW]Q;W-?\l
QEf{i1C+Ygj(>cGaQg?
4%9.A5,sh~Ukl!|Kc9a8)7|s{h$U?Km#=U=|A$v0>cM>m?83dR3qzBwMeD}i<f00hEKu_>M}@^jz_L?0-f!rZ M7w,EZG9BkQ141s6Wk sFw2._fdqhJz-]csn`:3O)/G`K/M#x2-Ai~,Xf(M69H_h5[Xy[m7WKrwctfnY: Y|G,`>Q7o[{(]<Ok9k1<Y 7aw)ddg!fg3tIJ@:w$1jzSDf)eQ8x$/oY'?z.#Str`|eVXL=.PL,{~p"#l	}$opI~58O/sq$t{mFQnA#{:g)=Wd ,`3iDoKa"R+]Kdyb41)}CU4x#Qjdc
rj}_'uez,MAKU2Cw^EvhxZl_D!1,EE~$u\n $,/|Zgrxq$-!mUnMNqhJmYZkKuv:H	UW2
<%i&=s-WCb|Qzitn|Uk;]LT`
QAb@l	`Wl8K_&3|=jeWiX\o.85z$P~}RBACVv]y2ZxK><wb8a'b)'uUyP%h#5EVJ^NJSpK`oKu'#
E!-FGfO@l).+='674YtYY7g;|;"ln
o7iW;'
O.Z>*aS(X4,~j	=A)5"1F1^:Ee1i`JBn$=QfXJxr22*t-sDPkHT+<ogxvE
OgklOfpoTLCKHT	{gl${/$|uyZ}I
,;Bfi5ZmO3	j7V^2dZ*_][C'DAzG'?FRwGAPe]Lp]Pwu)|"iKZr{ 8`"{kqC'$H_L33V@>0]QLt57%V |H'e} ~`R:`dnxA,eG]@!\ QxlOH3e/V@nw9GiIT#?DCWzJN\;]t_M?-1G}$7`A|_
rjCo%UJ#{$!W}X$5Eu%Pr?].cwFE=1wG&n%x]@M{_t&IWK$XiPWXuP!qLQa#aMv$-?g,LH)e^hvpT R7)`PUU,(J--Z.p'\nGaQeLG)IBJ&!|\d$^%KFnil<k*YC;'oX3p|`+p)n^`QMOFdy|3>xm&b>Wkaws	YePC;VfIi9FP[R;a9X`aqW:9BEv)&P 7]_<ORTwbc9Q20@&f	>"<7Mu{xcfd)Hc^e;8.%rOC)&9_D!
/Kn(.SP0xNNa=<$eL_KjFBm@U66Vy~Lq)[fQBy:`s766\uaB QIIg0XH5'M	'6L4QA8A 5[N$c 2:,EVYseQS2a)~#^t)|&k;\_b.t@qYzxv0?^3Nu!Ga_tmhI^etqNWPK?!)FTQ0@SJnFVmOZvRdE!QCY`0s"618*6R0eSzw#WK<)<OnC:hE["-tv'jXB({<9+Jyv^KT,Nxd zJ#*l\C]L\K6^A,/:y
~2e=aYz*0yy8r[Lr7Y9gRp40`f3bWV-S#+#wv9)kCiUl*UJ})Ewp\x3q7M,>yUcCt6*$2Be{%*5UtD#-ql@h31cD/\gBoj,f/O55rl]5<XUNYQC,L]LTPf|j[<gdpeU6gon`@~{k?E#j)0jBEvM{8w/mAMNYxq^yl)|?=',Ql+9Sig:<\Igc@:ChWO"u<&ycD}D-]Q ;XiuF0z4m!PG=UO*a-)T4*>BT'w#1JSW_*2a;H?q_
(CvP0S&8.)OH	5Tx^VsUc96mpRHxPT"oUCbE>Q5h1~LHTQ:{!b|HHpY/sb:%$."@jyi0;]_'dp"Y&et46FLDw~U
	oU-=^qzs)|KvG +>NN
#+t)'x]p;^A:^[P~u6C_<lg3oxmmZ]Gt&v	a}1n
8=gU\}E2;V]gyAr?rNWT3Zk0-[uBXEG%C;SwW`Y^FLc[g_V%E,y\A.Btd|UsD8|gyy)c+)2*JVM[=dT42}/m"Cq%|mRrkD:KsN}gsj-QX2!k}6=Y@8t>'VZ6d_VVX&o=s$Ey	a <VAU$03?&q;m%}R%eZFq|Ahr&F/E=Pt&bG;)*RmP&r}u`H|%MLvmx
F{_d!vGg/gbg!x[J 6nI*7H+s_E,@y|w-c3`Z%Rb	?	h'I58Aii`;53^igS91_MU&\KuzZ(mw2AKM[1aDRmt,{~ObE&of
1T*I$pM!s|/L#sbmfy=8mjs5<hGhL<zd?qCOvV@I,43`}%"|m<xNE')[`',w8bjD:"a<.,Uck0Pz[Ua8KXu,k)\=EbspZp;DvgB$>If=g|ep,aHV*\-H/$X0$daI}K%Wwh[87d=^Yp(E+Ks)=pj2Z`\|8qlY+O`T\P0\qGJmVi\fl56=+['7?03
qIf
Ygm@l8IaCL:J& ]0/*h~MakU(-Ij0n0cyD5k~%iHu%<34>eAaCqWfA i6m])Xj&DIlh2LpW6xVb(p\N7Rl&,XwgY-h0.9({<CC4]<?q3_br`Jd3NCzW'f4;xcS}b8u/p*%a
wPfHnk [ vwJ[QVw:uP`fUQw7<jBR=mL/0E:|%Q?rGlnc;QE6n^`i=wQ`/Q%	g59Y-Hw^<V',d,)Mw"IA(]r(<Nj/M=I{\0
}w
M&H:kjY%gn=N\,_YA%Em*BZ0tY*a360z@%-Q=Q04veR``%*
#!_6.{v=+iuI<N3M61:<!knBh6R-^#EtFceIv<#DCOj(Ry6F#'SCv2}^s!B}PX=$ZAb#%eJ
(0BY%LSwq4:?Z*vu.llZQi} -U|p:7UfoS=_}"o&a&oWC9&U[yN@0n^l3Z|sgu;EU,3Tu4O
eS27HM2Wl@:&J$k	R<Ug
{=8vKRzN_nm&@bWsVIb)Ov6O5)3%{z,n8cuQSy[M{q;*hmMH"7C5cnOY#Glb$@b`<#yyj<0p~3Y#h]GfiDi91vsIM9W90%7tE2TeO:5Z
if2uTBKnqil[%:b^/h9aD%e2!y?
v!WEn2o hm}&NA?d!S.EAM"c>3i`QE5jXgQdJk<4Rxs`2~T*k`>ptZw"	{,12R{z
>d]m'q0[J1bqE)Ay|x5]f ck"+8T|^qR/-9U\CHYE@F}&FX}X`TVv|J!lk)sXl]yNN+t*Z/),{K\'q4nx]("BAJqb$
#x] =RmmeK{#S"Kwq PZ~;"~.:un -4nR>U$IiPwmiB7	H&j=H@g?.PA9DUE`V5>52A}F1SJ^Cfrg)E (.}1A=N<-:Lx4Q3fvopc2/_|+PJuibL*Bi/_=I$_=dA	O.^d`FBFW4S;~E~NEX	WjgsFxvxY!O}GpNbo9[[LT1N)uNrr&kYm$cp12!27F|>#I9t6]W mo{U;tqah3NOe1I3rwsgE-('0gb?(&u;Y|_(BRpg<$U3o5I"v(%a1ij-9;134p (hJ]x[>TDzx'_okCJb:	 rVZ3wM #&s-Iig}''S`	T^;,d>UfV+e]mBU(l,
k\J]u~5Z(@=*`GvS7|[MNkTL@`cRJ#M65 GzSV"Ylx8Kp@wl01g,vS"W7-q~9rq"P5Olm\*gN}|qx.;ac, *q35XFT!94E/QADBQzwMJk53SW[
#QOEVpo``c'gw78u;%|c, ,Q)%bJ{@pzP`q}MS^T)h&dRWNrXx$T|mYly3(|5H7}r5sD-,TS)?E7Zm}.J~24UeGU>$9P	_BeV.H;$q3|fr>9/["G\J,F&~4YC|3)gb$wifyW)E~+`}\ZC'*ws$/30sV2.%I;b^3'"C#Ovn0rWIVbjU7PIj@B?u2/{u|K5\9Z]TJ`	)IU
xwx*9
Gb'I^37XCN6BfQH (b':~Td	vRq@`(?Zs&"
D\DBXQbXMFR=umw	X:PeHM\?!&m:j;A~g`[,<bZKNM$vzR;So9thGQ=d-_*SAHO!k5&lmt]Sqb?FHnoF CX>!lz(**Xu	dYFK3Hxwb\$YZH
.fl>_p"B-2J1nV>Eq2&k/u#8nR)R*,P,fWkCa	6}-M>DJe^_iBS'5Q|lTBd(GTgZkmw{hI*f%UU.R~w@9Qy5z	*]p<,l[d%*M"(DkT8$Q)"rn@sbGP#'`w;Ji(l1VqLPv>+ O,]x')6SD9Mi,L$#IqLhq)X!d94m{'
&C\Hdupx#.N+j\9
'W_R9X^_/kEHvV1,75L`OOD=BSf&DTY@\SUU|jt`~=NHevf&}Tlx[ eFH6v.;\:Gmv$-:l,?1ieq3XwhdA)58FsvmF0@;*hvf96yZ0w;wG6XPWhi@m<<OH3gKiu,#cR>6X>G)!3|v*Pa;\qCi
x[iHD{`$T@k!]+? )4>D"_m(%"P%9Q1)L$^vfF|^X{<b0z>"C:@ep^VMs:`
O{yWk1&67j'7i>
b=*%T;pfe;+|*w>M^C#ojAK5TGYwR1SgnwKWrzN#sk^#uXEc^X!yhkT,,)?J- E2~IO\/qA>lR*K4f[b.Xzi|m^n##BbyC1Q_E*5Kg
]w+Fh))Kg|ccC(*HYXx WF-`&H61IZAY1fC&J?]u6BQg$dc@0_x2_i#WZSQFJmV<MF;3|*SGLqL
-(Z3Hi'X)Z6`	D6Px2+\O
L>)"UK~m<^4 O0T(HpDefS(z[+7y\6X43:ZCY1veU8[oo!S(rzO-*Ak3rh(`tgYV
Th(drxl3<m9~u6Ts!HRS[{/^wqD?Ie*&?{0~|VehrF*WAo1!2Zfr6|=	DZ,udv"v<Z5ri{9faS](lZna%C#%Kkg4{Xg^Fg {Hp>%l??q-OVnF;=mIU+,OLe0fttajtVw^
v7ssE,Rf#oS[/orETXSO{J/}]
GPXjUD;Js^5p<`<4mV:=/$: !%}JVGs$maE,}`RiWy&|\!F&J5odyDgk4w7!.+)i0@o(?9hTwwnc7'`CGG`{R#GUjGmUI+ xwtI!N7p'QqIbOu`fAD5CFUEgz`=	IiUxFh,w5WN"58u4/^;:`q_lkaxVs#`H247's0aM`AhX"XrS"Y8*rkbYfq	T%*O.o':4Uej!jMY%Xu9;gxcZG|D~VV9}N:47ct}L
[b(y>TQ+*#Qr[u;m 1ZlL_WmITA8,`hqc&u&/_%C/J*e[5h 5x?B/0U-%P52odO|t_T``smHA}XiA^p'xyR,>Gmgf^fb^I&:ud[<I0j[jM<]ic>GLo!,o|6/#CG\zR?x$|sL=
OA$8.B'IH_@Eh,ku`w-TAgzibT4YlA>G-E+K3XQYE"F>Ya<0q)&b-V
_W&~Biy78dX"@iAI!g=GQT6"n'YyczeTJ;VSFmm5/L`We1zGW(\b#273~Pn0X?uA&<S4$U ;uNBL~83pq2)X]0v25u-36_:y,-6j
Rd!2zkcONbM~8~yWz}<nCFrzov2)_Ed60>/tE\M?\=k:0X[J#c	wdCmaV;XoG\;XzG/_&|Cv3Gu_A",XFfxl|1c%'1sOS,rXQShjW|7-{.c8nBTC$R)NDEq
BcH|Eu!4OjHNqRR8amt\Cu5Qo@`I4kO&d)'Dx='&;`w5\ c\))5S&Zt@@I_AbZ4StECT$}2m}%i@2=bw,S:pwV<stp3O"j{N}=?%+s"9\p@yQ".3*'Snti"}=#W~	e^eRSM),_7u;]TT
5xWaaRvTx[A%0mU+y`(6F5:^/9
6<Ospgvtchvd9P!_I}y%#gR3-m;-{RY#@Xakt9BSU6yE+`j-.7LMp=!_>LJBLY1r(r<T2vrsA:[QewKqu'/ 9}:8Uph?5$W9$zm'{}~^;88m
!G)x(@GU=xx!U2l*iY,_Z5M)?5{SKZZ*s/	?+aI&7'M_8itfMVlS#uT,+zY8.KLP'Cv'I&Q0_1fqt.8za;5C78=9l>^8	^p}J/7q=`	':<YK1d6.fo*$K0|S<e!F+~s3>Q!LD5[\oAY>%9P5dE^rL8)1K",INSITea
(5j,.}XDr$zW5x#	AW&i;/ cpcXmjMhV gd.G=r[40-<GiZzqI.&|W5*/s*I8O>@YV,(}'4'4]ECUr9Xx8[qJu2N9oBB"*M;yqu}Ce%kE>lrm$?Zz!oNe`d;PHOb/lJUn0*qF;{x@z*)Pc|(-a1	" xUw!
],	2Q={8HOjFcLIaw}Jb0>Mu{kesyZ"Bd*%32sh/q`Nkbb-9]8r@EDl}icH'&~l^v%_I	S)ekBt(oo"Gv?rBKV=`)7;	8G\*"(wG(
m3dg|IRPF8_C#+jd0w=?0|`N$Fw	V]?P6?k>rs,s7z12Sa23-	Y7P&q#]K:Vw'kI2zYZryQB@^RL{, l[.}	k0I"pFb`4omO?|K`]1m0p1nS
hO[kmz_H4?>2oa>2sS][0\
ri.]Rm..P}`SNhfz|CHQ#p%;Q]>loU;W:.#/	yNm;{hM#g`-\Axs;3#?2N_qN;D#3t|bU3)8qY0MPqIj)AA=vX;#'PZa3A&KcMv
D"@2'e(oMeoH]Dnea>3FHE>[Gidp|-T!Jv8"D|A
:b?m>]M$ca>> Y3ty-_F|c1M1,|2	"Wt4COnd8("yia-h.6_"84y{}[#n+)YlWz,(Ud_E"m=l&VnyG7O&Z[ahvF~,
\YI9]AC8dre}D4/%so|p0`YfT5$^CKZy3z{!k>WTX#^qj&yqo	QQg8O f:x[/_e:hY>6[h!\ b(d>N&FC;F51][vFZ1C[yl5:Iy}%|x~(h8Sc72z?Ilm;i^?>)@+lM*\hJ[^fStFRyVrSz>"ios2%,:|iWosyTl|,z>58NN:oN]'Ml{O}t)m :_`/;fs\FZ\t"IfSfYso6I7wYuKII}'F=UdDj}_1q|pV+$f(,UQr;wvp=e=-g;|PF5g],{KwJ0Fw7Odv#c
4~'	<OPJf>A		Pz;^PVUT.Y<bGs.KteVV)1&542Bc54U3,HD3 [(o(ep\D!JlyJh$pscO!]D4:r';')&RDn914GAQ:qj	XVVT m#-^\@5zB	-RA@ZZ2f!|KX0KL0<!
<t=o?uuK|l&DG%X+wfq_, [(t\kP	S.\J/\N#]nD=rcj|	W/8b`f^n$7=:mcRqXEvh9%ph{xS~Ukw{?$_Q&Jv_&1a)L!cD^wb<}StIR\Y(>M[tmJ><9G_9~u|e_<?qB0~=}S!HNr\2,"9$'[fRLn;^]B-:zM:6&$XxX7@G,r]2g(+%ebTD,u:W	VtewH}j4FU,Aza-mLn)0F]!YDn_aMnuLY=("+>"(L!v^)3cN[\N!u	}u;6CR@DywVjDLeMDEMC2r>D7a{|O<	/F#T~Qz}*'WU4-BA%J>zf7re
#FPr<t-o:o,t=lho#2~+{F@}i#p.s>sU5J7S'p);xh1tTpr<W,9|'
Lr^)/qB.{^jj#T0b~%FxO=<p+4 	Quk	[B$C>e6<L /%k9Xrf`B\a!>&cgiRgS\;16U"+F\(R7u;;YKblavW.[ib<*qBUOb'~q[XHNYV$K(Y	ouVx,4f|lSB	Q]2Lf6K+yi;a?*DOMAl>ND_gyDM]PTu8;T(_uCj{&Bm]sp7GGdjVURynkVA=w{9#Tw>f_I?3E7CyB~&3m`b{}Vd+XYN~u`+y86cc<[2/uHI*_KJh2_X/_&s$/a;`]&I#L`j7DoLSD3xIq{-.)0liRLqw!agcnHtVWGF4R_x9UH=q
#U9'*w+er|LE6L!#79P{z'EMSWm!_u[#^\z`7^
%mo#mGR[L03'g`hd2O;O5f 5AVpn<t'1rU--OnLr;nwr(22D]Udq~jE'AF]GvS>vZ]E1m:,fktFF*bG1TbVkK+6^>ISStp
0A
sbB/mmAV?&;NX[GF;y0Kk@<juHvNsvQPY6:[y]I^NJ3CQ8!_(.b5t/Z#ti%O>0?B'"]-[qb6J_b)0s^|&-|p>Jo<}3I2Pt0wc1S}jkp!Noa-Dj>Odo}!%)&/}&1PWL${3dQ*c^oY%Bzk~NNnJt'DO2=JAJs$L7PfQ~Rcd`?G,RiR+G5A7r'"'CoQt<EJ2KG#2
.MH^y)9p&jk}q+|	4PUVToNF~!QP	tOJc|R-qL..sr<xW./@35eJt^tgBT?5>yORC[?6G|e!|gCo5c&rs)42|\d*EDE/+-@|!?d"3"sbEQ6lFFY-$Gp~(WwSJ>;,M=NZ)v?7I{U^k_-=eE*|dA7GI}v&#Go+Suhd:&/qh ?la]"I<'52c3$`Sw;0#{zQyo^L~i*uMGF_wt%9l,.0r	<[0_768Sf=l
6(CP;+{PX+/bP#ha9cI2GlX/!hGo4,So)WAHd8F Y@G|k.rY[?W)bj1r&x#{q$F*7'#P$3WLwWzqIe7$k
bs^QU?#)S2tQs:qyU$Zr_gDv	A?B{8\deEQiyoPg*&U6x&~m~LAP?"VS!'7lU89 "EG5]F^L\hs7GH@:ZuAN;XmPu+srF\N%dzYWY6.xw.u
HLuPG5fF}bY0WJxDFyaZ/J^3):aS-\g5=7">7>M{yR${sX`]_x-QF<YtLIFumy*}#WtLgqctf&4"l3.5&fyb+T?Z$Se'#zI
0`di:8UkvjpO;(O	idmEM@ZhjT[KaI,/u[qi+m-!bdUtl<(TBeJR&h0	2#(0.vN}Y.)[CEXw]VTW73z#	KhgN5-
p}fWK
8BX{`:c"-MK4j^(xa#'eC2"|"m`GqOVB7}0qm!9g06z(BQVu#MK$VO(#@)^o (G}<1<sHJEQ"{
8PL{|2zD&+[>*"45g]?:P
:# 0mJ%Xe<MXInOKc%Kl>T|
EM}];SK$iY[d>t	`440laQIV)xzU1d4]I'7r]!Q&H@yDI>'/`K/vLD<GG@MIc}aQE%+}VDh=y@121q^c$y6LSJyE{0tx4L;I-a48}<1vy(o4Se(uYN;a1'Fd@gP'vp\JC^yodkxO-*>Az.Sq-PXP[m^P`!Ks%rvy~fG)hu @E*bf<949oyL>e>xW;:d8gy3Gi]-PBUA1aFJdqq.	LLbE!:gC*&H,~6}iQh=j.fv;5m=uk[A"l,3P@O>){a<U6t1\\NC|%%PCnB%StuDLL,1<zo+:v2*y!qKV@erA_.D^L~jc+0gZ:~.E@!j_)9lTT`q5c3;ThRz`ZrO)fT#xUDf!i(V8*a5`LTg+0rQ< <q>wd%zx1U,:GMxiFr|v<1>I<2[(78!Ip,6"uVI
;M[#I3-Tx\;0#.@@^~GnvW0Sz@Jpgz\F1DTK6'~d,yt&u\RYfWq?3cem}/<0vkgw>	LBjUh e	jv[QJf`7N5WfEJ!}Sm6E8_li+]21)%@$zAuQZ!(%Eh2[K3RoYu`iN.`Xi
[
R};3|6$_xQ_y7\9-T5i`EfmAmRl~K8`R8)?vxP:xP
~Gz]||mY#yJpsfW<'Bh)}f&Q.d%fI	hL1^qKBY4?N<E^N{Qd%<,~I%SfA;4|S}6`$:36dg$Y/6y6t@osF$Y%Pq	9?6sai<e(\u
_]w*6)LdGC5`	J-(]9{'I/2|@00Tbmi,z^E8/^<]G=a)E
VincT"ZPE]|bz1U4B6"	>gTT<s2:
TG.=(-".JL:[-YY^-=HZi77;(KR^hFwulIcVP'8\(9&"4^NqH8d|;uRTI2P
e9J%p36gj;o<^['~^Mm[g25k
DYb`z[t<a `<IC??TX')pp`hyNLC~p#v]XB>XC1v"]'W&6ixe/n}+\/<J O5/wB9XW*9BVU)k
v=Idd4AQ3$V;jYBVAu
}6vUbPx0vn*	.^~;Ao>]\SXpLGG<}4@cRY^6__
`V)AIh
3/xeF7@X"+GvEU
o6;&3FMzNWpMin!5r#dLMJ<9^$Dp0+|Esyf*K6!X(wS
TDEzV6
1T7W"(mdLJoM'k,-zO6P{6(92TJLnW^U{V	LDQ[&,B)-17!03N2l "9iGb'T%UJK#kG=&a74_|Bt&e/,B$IoIo/;xx/"$^Ed\~ |'zh 8}HcQkG@k@Sf'*0&tg7)iuX)*!T04e025Sa#QaEo1&72kbPd{Nh;8YpEz`[P|}!'*^v&o~dV3iTz-	DBymuVXAF{ne2-*^y8kh^+vhH(6ylN*
";`r:,g(A{gn1[,8\)aW-'wjD(mE\Ft	t#h&lRZ2e,QN^cH6oQ"c32X]@m6 7a='SdR_90?K}v
!+|?2Ue'P7qTqpPY.o$
@1@JQ*//cU/=5wl[T@jX,DX#bCjt'MxA<"#@3EH	6B!@*1mT`X8?eQNt	:XiFe1qD/ PXJ3,U1~) <q[Lj~SY]E>o[Fi$O|C^H5j>5[;t!yP5:=0n<yiR<EMv"!VF}JB.~<6red	6Tf%7FED!p*I*'Zbnaq' Z$F^!y4WQO$XU.+E-&DABT${j2pkZPvdU0S-u0#}X"FkA3`BQd@UT'Q7. QZfjW&CMby:;dvl/!XfH&WK#BLqtiO5l+`3f.6;)!|sP>q<m+Gjvc"pY;R{_jJ(]C"$~YQO?>i5x6xlgKS=>KQjTc#KK+#Mx,&?:BFz;hN
O!n!B[K9PD%N-r}y^A0bWQ!9(x$JI|hfO_YPj9%*uZuzohL$@vs
f"Wve"3lv&*n2N@#mqSkG]\x$Wg)T0j6A-2R$=%B3H?0~?$"#Q[pK:	TsJZGzF7,BMRlkbUQ)&.^aL[ iz;2-_.V!]|6V4RAq$iY.=
gH1'U&h'|fR&YZ<PFV.cT#`*0"!(,8t~1G/t/$XEvrPq3^+xUt0 a>? E^0l"IW8n,QObElfx\{H fFn$vP.<z[5xCMb1-0eRrPo@@hjxZ""=&dw];b9jV+^mx(<hje}J77USQt&*L1U|*'l@-xiSX&K@i!OTSR{HDjzD>z4aMn6g<31!gU3lpGM\<-VT(Ffsy5vhlwAKtkjY,8tufnW'CKxC<S&,n6c(YA?pZv.OYARO.3f2G"_v8db^5
tV:8um8QLu{kn)t.[:4^<{w)q**x~:g<)_LMH5TQ}(A0A	X t{-%\33UY?Fd
atiG)bWDX1LueSt.	ukP(se(NP/NY|;< Z2aH;{0Y$uFa_<2wKT.Z7<tv R*doKXx9>x22w"@Q'AAm.a@B9bsKv@:V"OWMrz1TDu))mCJoSKyO460n7Sr@uaI.<eHB:XQuQ)p5UvR@bjyW\-@AV-l1(PZ/me-v#\:7*u;]TkRr\$WA\yp/ezc7D&@f/2G3#Du*Mx\T:^'I4a|y<7"bSrc}1K;&{l|AL$\+/VieoQ}1(/=rsuY)N$XWakTLA	ME\J&uE)/m58.b7GO),ho0Q5%Tt/%'e=3Gnbpl\<
Y 19kP'0[rK_Fw=`=B~Ny#)|BY=ZVb)UA*\'p?	lj(~F9lEUBHxdMUsR'oKBRGpx*