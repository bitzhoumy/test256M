VUx;tm!6!8KH_7x!SliTD UDj*oQ>fNWB	%i0uOVLn6`(yPudL3ly~50=tQNPi,Z]|PeH?R4W]T%Q9!g,dqtnq:vB]{q}IPWQZ@iV<T];ckRppTuSZmC{NWX"x=-FXqD/6Jy:c'iN;@q<X{\A8Yh]2w!L"R`
~V):k*#6IB3J-z<F)oQ$#/(aGF%EOit*RC]hSR^Q`mqYFp\s~{,VD@x+<&v8=D721OW1`lfCnuu![T.6]S&:~,'k'HwiUYto"3V6D38;s_RXz	./UY:t8E	Ry81li/U,=RgT7P\B=no$W9>&2U#nD{VhTvT4-)<%vu&AOk_&|*E%36Wkc|R.LB&p`t\RME'S6sxfbAlZQXPal\aBVCs-D3r[yM :u&YJSE!+.Sa*}.oY]L!$8&za\_@g@C<^*kPA) >
apLUKx!M?v3vD@N'/1vfp,?9V5t=^xLc9w+yp!6T[IehU_\gb6 a6\M<rM-h0g2m>KS"F1s;:x]x4ChO)?p-xw09~aSa'UGVrdUO5':Ps.`-(F#" Oa}lmMxng4S)HgHP+]cHhmG@bF?9*h~"lUKIL/3uvV;&@.wj1x,	QaWQ$oc^QvT9&B(LIqyBh}4c2vP*BkpXTR4v)J<F>$CxqA]hgD#%p ${qAv<GxM"i?g|4l<-0F}>aFF0Pb+ankn2Ko$*E;YOy.:BqC}ov%QOGZ=Ek\>kH@JQiDp,&1D+/	MS1uR8RzJ"+Dn-VXimg
!Iamp!2#B"EFyUai;eW8$;6CSFKUO"WgM/P6v=&7x%=`Wpc	xt|em&k|)~PNs]Fa@@z!y&E}t\ i3Pz}W3`;79
jRxs`4ao\;bg/56	s{&:Hd#p6~ItL[S >u\6
C*-1b `bn$4qaZ]#We($YF],uKf;mrCc.2\.ozvc6bPP/|!?b9"%$~AU*vdbUC0{7u=*)iP\=!|RM|
02*8i-GW=f"784eP=wgrhbs`@Il"b/Y^V-Uh%X`5~4^ZH
eW(xmF7vh1nn5cgl:
l3,W {v(9*-#n"Z1`lR;
c>@x=M9I} FX_GNMBUl{2;3
;p'hAtsClG@*+{GW7n?"ABt*(TU^3@`gkvgmlkK})VSwP0$x,H#SfYU7r<E@Jrf#
^j89v.=:w)ZN[20BhNeA!U!,v2\ve1Z{_B7C0[e.UxhP!=a^)rJt63I|WM6
qbz"e-q@r~LI&u)8H2N_Q<U+)6`D*S
7^O9h4\&Y[b!(4W:D],v"(q,</1!@uo`TShL	wsZZp\/yr9L4mapB:;rSl2uO@	%hp-]ClIu=Fz0I|1tE.5^2>FBd]hnYbhh|wH^xEA&ai/>K=@Z5	&GO=fz4OJ&vn,y3qCShJO9.4f4}6T!01Rl{\^-G[,-O$+2z);Lf>n*vgW\/EimZvk-L@$UZTs=>a8j(Beg`syd[LI
Pv#%WA04-Wq7$*gAY4Yx$5X'v|-x^^Rpzef%?3z\5iubb[BWg~1a!(4a05vBH`):(+?\>z>6C; `M6>X({^(hy`mjcRf3k]6J
hpHA^a&ykr\)ZfqPPq}CD,cb$Vb	!E#pa,/&%Ha{%B]bBr#eSK,v`J@+Iuz`?'p0u2wz5>:_9'^E:pn2WQ*#C"jHul

DGRlESGHjXf,)W}`0fY/l@|'k$*g[*sm$%INQAvF77O	EjP:1]u-37bsb:L|Zq9|lr=(i6:GxXECTz6&Q:.l~N3AYGSk;n5+$1	7+9e:Ey)l5L?}H10B|G,w(GHy4pZd?ddum-:"5|{DLW5!I.7?+73$TiYQ	?RH #4k&^8;U"|;a5]=t#Igg7AKO*mgD0iH~P<dn]f&90@S+R
.nHbnXIB(-7&`&#*-Wk;QC1YuTXA@d4wzEas&3t|r/$EjH'4BT]Ol$Zy1dvUTZ\hvUGesMKC+)aV:N|&f^Yhv&Mbg>+gxXrN,(U;Tkbwp@1}vNsviH$L>R"E0D-kxxJevY1L0y(h\+%[aaI[jk;hCl$mji72J4E2]5XqVw{-'}uVkXi"#Oz%[Z[S>LD/^>yD>7Y;d/mIjwLw+YHVwK%	M,s;;RS/^c!@0]fx#!XJWthFP\QIu60]AkXd*AHDYxJ!_tt=`V[(0td
d3J33X&PM;@d9B5&\+P]':r wNr:A?+kx>3%UIPC{f1FIq};FML9U}XMGlu2p|}nDK	`zP_|C)flzwoL)2Jm:bXT\{d(jin!jYe	Wkt,#LZi	%*c2hOFKX3 aU	c#3a@%#(znpC1c!5uv7\4s0fv6491`Ww\P*nFPX~URdB&'HnPV}s+gStKe7km/##sXn$	[Lak~(HPX#r~/ff0LxB,D(Oerq9,O/A{NDGQE
~A-B&$Z*nkz;DjQ$DDu6{2]C5H<xxz?|
a1sj|VF CGw1}V\8s$0=d{'][=2Y@VG'%Lk%EGUl^zYveo!#AuSR
,[7Hm!\2wQjtY(D-AfI9%wW7W
[8.p^}ZFC|b*N
\LbCa`u`w~oya#w/^rg	F]grpZs_V]~F]s^WT?d[S4yILMB_.UF$vR?	s-s,q5bzo|@E+J@ed:dBa<Kdc^x?dMVx-H PirmV;V:=?a(k:s@/kJ	2tsw.*o7`*n&sK#t1T{7`E>h$<VHyUa [)SAZJ ;br;7oiR:kZ1YCV+@446<UU] ^-'/p[+=,<0HHJ*Q$&>c8W+84k6Rq+E=SpwQ rz8$MoWZ;>L&cBWr!zZ3	c[P@eBmW
B*EB	'0w$j~.Hc}?*mO>[lF2(-4Y]*2{%o'~:xqII5~ cAQ$D39
7s~KqS92543
[P;uj&A0);cxW}X<_lC>\z}\C([PSSf^rY'J@5pcS@[}k( p7*pfk^o0&{|?]n	MExjH6;BcD\Cx,e}Eu]tu/PmT];f\f..yE+;gL5^{02LN*3'YMz>E/AQJ ,'^mx[`jtLlbg 3E,z"'TE;
e<<,pv1Vx([TNU*8y<.&rt !]S6%tuSnI\QiA=^KF*C{%	XT1*s6m9EBaqDV2k0[5@Pr5Z'dIhg("W0v,/h@,P+a*7v^B$dd_H#RI|Aur2l9aU rrB?8c5^oe^ps3\L|t^\	zLT/-9zpa|x|N'vD2BG*z{llgsijV?*gyc	oNKUY%fEVPCgYoiW0(srqN#J.`#OM8oEplNg|iEIjxa`Smsm_tNwny[)MUAy^Q:u&5_V99Jb-$E~Z:SwIP@i&.`5,)/@Az":7$04Nljkk
dOJ4ew
#D(eI0#PxR!?aqymQ|[`d%1jA~C{6;jiW,<	\%|MQ>+[p8xI7@$nln	^3bo29l^>rfv/m^a
'x22-==ogNF('K=Db /]{H|oBt)Y Wykz qa1kxgn8%C(i,yp C	}gkcZC\P96o
J3-Pd*BT9o7-A&BGUgsI36`:@3V	j`U4ftFd4}~aAtn5HO"cR(}Z[7QWLhbhT94a[G\YdK)^/33tR	tq7nE2RstGzt|P;fP (3kB	}uUXI5lxy,V''f+/$tPxezN=
o_'a(hqnfn3/z{o{yevsDi;{XdEjOySaMuwwdLRKZ.m-+v0ZGRFoW>Ty`fe)^{m!?42a:pd4$).v.Hklp0;KH'@1Hh[>KOiZ}R'{|^2e1brfMRug#4f5q~8g9CFyZGG,+wx"6B3_b
Y-\Jgre!m9cuE+=)p}_U$&a	uVY:8z=&.L@D{w:>i<thN^r<h{N2lk)'ae6f`kcHoe_fPxM\B		UeTu{~bDSv?H$T|]cHv<lJy`OOQ C(3iBM_X`&o5x"B]i>-9 43ogJ}UbJKc:-bBENE@MMw%}._@vU+Te+Ku#0~iO7E_|0ZW`%^?>Ja%rI2lY!y*9EYjNs	KR]d1sme7tcojfD<|C;mW`?!A 
4W@1PDdK]wc=%k!}(SV?e/gnosndTujtRX*G%
kvB~$J/aSqtG1^% %q/h&b)O7jTjsddktMX`|_OFZ!}3"@ig`'-qARL<nxgqGA/0.0\KqKLdY1a+/'(yp49:S]y^~Z *<bp r?KO<.LHYv:t vJ7"l U?7bXJFF(XN0IdgJ}[!D'.QG>~1pw3PGb@rcAT'dVD^iB]LUq4?g(t0YPMy F"',3Z}m]:S|ZJ^v-H]kTO1_3FR&">kg.%>f=cQRh>SH"tD,a*w{E!L>FS!-9V0^ EqJsmxIa~M{$*rFq-1(eN}g}	b;GnUe\A#m>XpgzqUts-Z4@ZI;aL%8sr7YO1b$}KA>~zqG)UMm'Nf>ECj#>dmBo-=wB >noWBOifYJ+QqH- ,i;6QP&7>0=6ahV/7%fxo';{aB2&!|2XQL4s2
byo(I2+j5X%#Po8VBeGxh!@F;@SbQn=q?w4(LMe UlKXnpYhHuqTcvg{c^VD$4?_xGvL;.miEP>LQQG0vw7q_#ZeQ
&_'B.c}JDm1OiBdSyD_W$:F]ImLA*\fTaV(+@Epp(IeabLo,]{+rK(*z}'s]jn4i?puplM61gxnsD3}JF#5{jG3~7t|sYzVXt_26mf#`K0^AHxQ_QrlR{OngC
MF$cpRxU|Za<U{7,]q0``Kk;'21H0 I'6#yb7*xl{|8QB0TGm?(p09` ]r4vk6{]0]/ChWz0vk%hh/[JH8$6:.<OwAn<P$.\cb1<q<!>3zLuZL"<#fEnik(LJ8h;cUw$pM$Dw94>*Q`/7'e-pFUTv{C5)SL2#
HadoZ"z`{Ek$RF>,>S5<Lb
P"}w'7D?Y4"Q^KuZ:&4&Y?y`Iko9u:xZ3E_GLQIsBC6QeSFInz'`s3	SwD{KGS3X)OD@"_Q64^Zu'*NBTL2lYwK9j&~R qfb3B|dgPhca*_IJ&%7c[SA@I7vIB6Wv}rN[k.Z/|[]%t`~/%rE+$\wd_lTsT[foqt8'uoG(XpX8FL7^Iy^}qx9yfzL}td2<Gls2aV|J-7dNdETDK-K(r&+?b9	4Hp1#z4@Vt4|BT5]L.eaOHzC]x{V9pjk;i}x=<u=f,RAk$( !di\4)*X,/&>yOSl_
+sVSL^(!UZV@ok?>p}scAi|R4(i*\Fibn$8R"/b 6jeKM]S	 ^wKgEt>EoG0;#?]=C6P@+xbzJ>)h;^Bl*AYG;BV*,3HjsCY^DAvk\W&?kNpV)mnezAj^g678\/Ep=Z}?v9f]:Yqg6YE oBitu}|rvp<>36Ro$+]AK3)Fl3jbjFbU5]}'MXoL6RS.Gi7m72EzNV	(-Rm+.ZG6$kG"_[)RSD	B[.]M@LVl*VpAc??tq's9b`>wchGV[AQ1G4Vhm
eEiHhgpVS+'/	+4"lKQnj&o7\0+y$sT@1UJio'-7j.*Pc(?TBQAiB,e53iea`\$6Gj*_o~gdN$r!	Oc{2T:" ^9Hi%&b[Uw(}Os+H<GmkP RUHEcI[hF-8!NrI3RI$8V?3_ U:jbDl1aRNfS0\Z-ihfY|3aAkA>=wd
:8
KCCf}1S7&t}	8r~^uwhJUYm3I&uv6ust7(tB?a]RD	:i~TB1f<|)R/@qEUmQuQPXfrbakZCCb+8JW}P)nUS]RXY1"kDK)d:y)`"z qM:Kq)W:$R^00t Tx ]vY4J7$K{CD:1-?`x yJX:^(IKgK<A{vSq(tqw,W#%LKkq`@?WI*	qq.RwO^IHB9COAVt757{yY/`0=66m`16PZ+'%w]qz)QG&R,|+2{WB!IP\%t	vr)_s) }C\ve&Yx&#?4eV{^GHCg	rmIF4VKq>`HTQr`TJ|fb^f-a,5h^AF^,1V15GSSM'9Iv,s9}U	G!h-6znm.kVX:7k@>8RCD'+88hNkB5C5uXkui.k<Y;q2}6mfcK_6Z|y\8EI>9HB6X3Z*$O']G5*Ru$.Y?nn.<e#64L\n03,5FiRk*Q2 b8?R@t<<[)I(wkfg\FdL#;7/W.1e<fuw4#`gr8|MS6-B\K'%VeZk}[b++jH{Nz?xJ,qzXx\*ozN8Xj6cKX0*SH!|B7j"&dJ&v<D6KY
ie'#"GN7(]g(p^TYWC`\m4#6{Q$7g'
#f%x)iCwA2{`g2fkKMH?FD-4R]F<H
aoc2qx{d2dZT3T=CYEk(r>ofXI<4-#
:\~8On'|]7kH0<{1jS{Lo$d(u4	.Y1uF`{?x,`X$RDPz
1^/<hih[q0D"Q)zbd(;\+F"4grh.ZV)-{;?4!,So}.HN~Jvg?"a@>2X}7@`PmAD4)MG=6K.@~%'E:^rgWUc8sR>On"{Q|e/PID3d#S"DFp+HZt[kr{jRDzk%[eMZ,
Io3%}FJ`ow21}
_(3>v[Z^nt~= tpcG	/mYb>}u`!ru!
>0x	SpZTtmDI[zV;}gzsW0w&
VJ8J6nhL?^fQok_1yGST-hLMjfEa6y`%|:aoLTZ3D M)[.}z/dT6tfJ&N#_9G4H5kG-f(ze?M*ue+=?Y?jJh1PCjPtKYV#".xIm$ZRysY8T)Lw;](O qMD^xR1dNu*Lo$+o{
n=>Lwr^!@MA3at4iA:,FnjH*dO@'d:iF(!Ge?ta`9=	#[t>7jd#4{nm5<_-wrKf!KXl"|r)7@6G2pew+Jb&>X_vo:8n_)DvV3?.].Ik#F3<Vpk3^ky]TEsta7*[%iZ>2-t)~i9#Hk^PUn#3zKo
Zx"L	]jfC#9yga,#\p|/}sv'va1#]9"=4NN(3t2!mDH(G_I}6th'.{M(}x#N//3cGHlc9Ea"&Iy;5n7d8bnlYr.3lvSR;9g=Mq%x<|x#D{G:7
6I5T69v_N6?h_?K|]C78E{*n7:#x+e]0j/y(R[5p?12?v/,EP3XUOO]}}~n;o&
aZDyhq-cvp+gXKYE+QOaFSgq;7Z4\L",19Ay
?)1M	E0D9;vVw"6\|RZ]0Yn@kjP^R:U%?s_aEm[licvv4Xo|1L*pP0YfwrN]y(eT`i>}iQ"Mp$ClIA,][d}Y	NoHUR^"4KzQj@Vjj!sW:8pgf5riGWJvO>.cx)/O~s*]-{,*]~s1>C`'J-7BLau]$^ax=.Q!!5JhZpDi$x>^>!kb+XGv3RfWQ7X!&1pICW,+c-jU`o
Q:Mc_np#|a]L^165BZkTm7f'>=FM-JM99os5gz/zw!SK!ZAm17g_8BF|B_h]H:7/AO?}y9i}1r|3wv$Np(wK8a`8"mgT}jP5Uu~%oKzY@V5gD<ih	P.x8^p1XH9(`{NiHv2,Y#Bct-*#p??)"`d<Cu9Kt5!ity< JFS4{j"]W$*=T2wI;)%=@(Teys,8@vri^L4/0x?=&h'@>n,L*UmF%']@3A#nO};@gK^)%Ce/WEnGAq}G:&N)A"CK4g,`+BNw}ri'tPZTw_BsolW&^hh2uk*l?}FS3{pg5Y([Loc>#,T~)&]Ym<>2fVH|AQvOYb[1Q)7bZSg@%: {J,BTuStM>scT2h]`ob5xQelc7?'>4Jl%N-HAf='7md}+eHSt>S)t89iBlT2!Zk@J4<q zu~L[k9w\L=(a5ZmJwI.`k$JWl>!`+PGv"nC%"6fM-[P$,<7Xx64'd?UN[q"=0\Z-,W*
xZ]}0%.U#:D4A2r"72>9:LFXjVgk3MslP{J*` 3rJ^,b}T_S'*|%agdbG9KakZ@}`{:wk+Cmy[,sOxJ0]c/DS^ykbU`PHH\#S.u0keB[=\G|+;rH[9`.WhN$@:p.a)t6=FzOr>0$4ix:$z;72^8=1Pioi@]te:9i>gdkhI
EI{GhT&e1#O42Bs>CC)x1y|?_@&DU6%e](du
@c="-kWJY$I3 L#5?C4FnQSQDCD;#G;hgc-#^/:H,nF;Yur{Xn&j(9;P^D<MO.f( BU. 7W(u-z\9$:89P]{r]cv>6eq51al-Pz\Y*n(zV-{g9<Yly5	k(AcD7<b@?X%g	3)d0lLoI,xYk"1EjcMrS)JYfq%v5hNc^jj~)Sip'+JTg8PT
vdaZ9HV)%rDGJ?V79)v$l7+!0~	h}-5a4{4Q%#U1`a5j7Q!iU"auA]]&Fh}4]~xK4Huh/AR-%[bi|+ W[O`O+kp+fixFI?EL=E@t`nX5!rs,@E "J.(3N{xb=uh<S$;c~_
^!1DBlc-]
exSPw7/*X%MIYOCA["$'~2di-46T]0rm,iyZ:lY/?[|T|PU)ojV!t$`#TzWscu%FaR;"q#/B6^PI[k45=Wo)5'8C+tfma	P){K')'h{}^\p#tC0|}'i7.Tjkx
3H-/2K7r4Po{\n_d`>Qw:h<OrVe:)0
fU*d_H	*JZ=g!Mpm!>`3G%U%GR/M;~},M	ouv(!Xme8<9;,05Tr\u	vyVT!|8YQSfBcUF)+,dE%{Flz*n@EyL.q*A0l&W7=:L5&7U;~J8bs.8c3Q?![][~S{hQ<AkfNOI)L5#^379?czQA(IYqga+ OQg2:nH.u=J^.H6_HU#ga3/JyfXWH/=vTu
M'-o 0I;V67p[2K>q6c8lrEBdZG*Vh_tdBi@i|fv1LNu9}`i7de]\v 79my0{4{h\z!$/]x3:soqyR=>zx8B-,ECW;MU&R8SA1
)e	")IQ3be<]|&Dy?0.0qCus{K[TV}P,q|8pq^='RV.h=lpWkkaLc(5	hEL3z) )J-(ENQvew=mpUs>j2o%156W[.6.+6xu}%%-,bp2u}^K5.!S$X
o{gQ0*DbT%: !I*<\%J"K~Ic3+q^VyX|Gc&1cUUWIOs\b)5Nv<.K;	3PSZ61M7.i c(fD?S#p6|c#D>>x#uV(+!-!b+Qum\CUU^	y#G..?av,_ik%^g#Z^OcGTT!R;w:x]u'^	dPG]!>"OF`Ti+lp
B>"?*xU<)bSSCk6nbOFE_YI(I'wYWP?:VMC?XOHQTaid;?	|]Mq\a:JYgJXs}GDpG,>fwU
]UB]w`i}n0;?UvMt^xzf,IRJsjC2;LXz^q3?OL26{.^	;:s#<sTmdJh#/FD)~Fkpo:gDeP|4pepxo3B|%1_a@WQp;ryy}7P_,hX^$XrT\io"rw?$6-<Meph@U>WI4u3dMfR`:+|03NP18trO'xNq^57Wp,XX6?
q1hh%X;va0a6~ymCzJ%azi#u&W/*MLfgjf!1Zd@8}P7q$|:_i"e"dVvA^eP-OpRSWiB15o518&vAK@0K)t9]}:1	N4-^"vd?MZa	Aqd[[l
o(i_X
PwL|UHgF%^E0SwAmA/bM^;|mn4D:`3BC{C@Q28mu)^[&d[2#@B>NsU(}G^eG&Ypn)vbO8
k7EAlSK1?nepz'.G%!q$w8{'P;%H,}WT5Jt;]qZ+"kMYq-7V-}\$o-BY%m^Bdw^[=7#$=)pDsJID_v^	Fsey3	QnLf-q^	LzfU
ThX&GozI%YPK("oX	xki%U1}#b|<Ou]+^'1W*[voUY"8k_$;-#
tOt@Z*w\LvC-7\v#t/#X!zif6;FNyP{[7LGljH!a4G[.y{FhPRCz$8k=6xK,Yi?V<NKEgXf70t!k_tg
.IM+;#FC,,qE-~,/+a{;_qa
muhPF>[i<ii2hQf{4,g:x.aW8d)\)ZL\m_="tW`4O]oP/O{fxv,chCk\<RJi 3NYu[o\5>f.[l6(h6oq@v[XKl$71L\zrz]9Db:-LY7uN`LJ#y`yzEr%>ANj9iALf>2y)JDtujcD&!O3~CSTMjmh.unj0	%6Sq-z17Z:Tt)h4	 5X]IW|?G1Z[(fx 9/[/ZKYC_eA\ObFa0y${9=h[u.+_!Pa47U!qEC4ELp).uWzo26~&b+{6DPh^N`\8G]9:haT;UEYQLBF?:|~qXTE]W4s:qf.e<3<7aap"&6Bct4\!}Yn_X*[N9aeIU.RVPgf}UP\8D!a?^ R=elf|*I<[b1dh<UDdYiM=lH55a@.G`}){,xHS  ei0	[Me<)cQ>
vGq9BzD+:cp ksna^Y\/0!b$
i1)Jt2~.;dH?_`F*t 8@6^g]n/jOa%\>ETm Z%ZmBY)l&WR;k@X8?9F5i{?Gk3CA"7?bj.
xuEi*v<H:T48f#}I%B<$Y<2z>v&#}sP[b[H_xk['"'?|Gq&Z~1%-qOvp}pM)d>'%LRRSbwHb$fH}`*93Bbl5&c2J#=8-I<*Cl<>A-H#eZY>'$uGRYCiDHs>Vw8aiOubF2\B3^wsherh+zK7m17L]1V8e,P9QwyT8;ByPu]gB</)6vJ 0r:riLrF?ZR7-Lsd YE%P+Zr3a] P&}a5-.QRo*=CPj`pnV;1'U+t`wTk}uteJ42eB7sA|K{spoVj8l@f`HXRjCAP=ge^Hj.3-IT.)u~{)9Fh!Q>`o]EW=J0{+~B6v?dd=JcWZChKFPtsh\%<HBJVKUGEe4R8gjufXAcu*,F5fnb$P&y.4u`Yscd"z+N8B]{SBPIF}6d1;bl-R*/%nJv%]k,nNRemx<xzW,*|7sjtSv Dhqf"t6!|Q	0~`T"E@^9Ye>N`y6_[.Lf2!+0L|++*C;pt}s`gix8oMWKK5X:j0Y i.0]'%`L)U.%~wSn!q&&=zEcmd>'''e.|A?7Ljb$<b1LCi6Asth1bRWtjX<1p^1K==Zd6'*N/+J*[C'"L7C]K.m{&b59m3DA$*dNE}Z(@Hh>2JmozcLl@)K5U#PI*kMqXm)bwE#Y	+^R
*Kmr)]di.r!0a
tPE`AOsp,XW!|$+V?m\w1EE`eAP/w=Sj#cJ[X[`T<rIi4T)69DAZn@wY2\T,sBI@2':w/[G*Z1c!_M.ev%Z7gD<NL"mo	"iT'umZ/NeZFjFyAW!rI?8T5U`0Vhbk=qX2edE{2!R)G`>w{{%(_6 *U-4w/w5Oeo}\YpR~)y,U#xkesa>9CTrS$AduCJU`.sLV1T)/m79=!WRT)MCj}"~K!NG P>BW[3$Wd7hkE>0p{aT&dQ/}Xz 1K+[^*J7RnZ/,Q1e18t1cXz4e;L#7BK(_xj;jhditB)f.?/1j$8KHs'=akM.dFt}QwR9c[[D/cvjS5^qnxqVAU|nJ7 Vy^6I!8GjdC-R0)@Hh][2c9J3Br5+*Z_7A]&r_$*hNHDWSo}#/ 8f]r#<w:i%<u3xkSWY.?r9"WFy|/\Ihr\ys[?FjTj<<@&PIa_ygfC,d
,aOzc\^DXESbt%/&AglW,DrH;Cj;}29/"ia)ie)Rbf#`/S$uD#A&WTwGO%nDlS2eR0kg(.=XH^*'[_-mpZQugA'w.&kz.eTnXdrz_QkEh7B]-yfKr@:Oes{PR^[xCGpI&.vt|v/=RPN?5I'$@X8SO;cqV@c@nXuVHYjLeYxkG4?s,8OciU38aO3P*4fW#]OkF@Lx.=_Y+[\$^f$7h0YV6zTDCPp8Q2gNE)+t\q/WwRe9acsWQ9E eRE1!kDYe[fLM*OA2sQU@fk1`#06/>!>K6.;p}Mn0O^8n}{L3D/Z<En(P+HX9TZX)_M;0n5%YRJdkUs@Mo{N	gc3G65^eEpF>bD4fU}{,sIszLlx/)1LepnBV|?PZykC@3GwTo$JGT/(eRf;0qf4tn|=o/'O>Ce6NHR#["pK[Lu2{)J7$"9!2V@*=}Y-#vbos?$h+R/^7qO*tK11<BN[QD#>8]2nh#8kdQ\9uK:]?f9^lv+fd`WT<qb~kLFd&ANZ]Ob~dx,R55w>.Zb7rJoX3|r}E+mUUu)uPTS^lh
K"oHB"z,ov/gUGi!x_IMX0U/{Kvq|4L4*$Y*e:c8}d5/xTYLPW3hJb5[~1Lwl	*rMC0W7T+s)om>$sP&n#n(,cUXgZtM4Jq>U]R0W[&=sTd-wa/c?k&^C7aI*
3Y,zG.;87,_b/PwUG>+F62.MGu/^P,@kw-t-kC4kCxPGS4HTFc'[U2&B:Lf\U@ZpGST5O5}G,(>oCJ:%<B:u2)o!$q~2=5w2"YQ[Jz 5n*w"G?6Ql}EN>dr~8=0DHcZ`/@hEDEXz[	B\;AJ*^-U!s_b8G)|rc5NH<uTm\a^oH["QM/=U}xXA2yqI0<rwAn6k>x	a.4:bd&Nv&BOksl`7+qlI{En3@j)0##k@5oJk/VFc'a#-xU '*Nd!XE2F1^
`hm*	#01Z1,>z)SJ*y9m|Z{n`0q"!Xxwr{zY56Uip$^$]j,uKQI?=7d,G %OeMRF(O0;3#$X+=Qe:?Y4f.a5{#(1UcRlQ5B>re*CTh#{>WcTwE4MP)SU9W5voy1@}#SUV.aRlgi5J&i-U+o06'ptC_XYUfp_jxv"oBrP+t0]4A|PfP66"G{5WrgujmcC|:D{}~7]xTtBF\Yssyh-Q"BOsAs3{AD#[x]Dp=#3Jf8)QtifmMMQ-JL79Cm&a,!xyF|7kQp9c1a=ok5F[ggI<+0!Lq);2Bt@q1u`GbYKL.duD+FlA	B-woug%VRQ-IiO|^;R%[B>'Bb:ns6<W&A44FrAVW{{o&\8S,X'cZ-5,Yv-hUYBb1H22~sT2OmD+k&tc,`^MC}(>FjSGWv>0"zqM2 }MST*A$"wB@nYb[&X[aYC5KB.(w%/~1Ak=:AJZkp={NAz,0\8j(d"lNqd=M&'Mm+yD!cvyAMQ`JM@rm/?/ICk2X~xPi/U,RB1^f\Y~5e|+tC|T"\_6Rn4Nr+xEupz4N2~9LI^at,e\	&x8v9T@rdq(pbcW;12WTA20t#W{eX?TPR5ilWPt!TzdYlvrW3&qD'Z8Ksz
RhB|G=}2_M:}%:vs@u|M$nk(:! PF1W
g(
v%LeN0FHXyCG4bnt<rej&vk^gF`Lik|9NAZKf[ydZ75%6~KM%U7~3*Et#c'9h7>B*Nmnm;z#yzGj`M:f'\XzujTMD2>RDhwG^%W\kW#D>*dgf:l	LE<u=#B$&T_8U^}``(T!]{&PjO{1R6MLO0k%uo?3QM}W<imO
t1"h*/B5*H]R[Y}0l}Tv?s572t~<-	G_Q"*vl$<YBO$chn@WkBBzbY\nv~vtA.b4-v2vjn!0_zrge;jRkSPujS>n<ckeG0RD\uSaPLGK3#JzI>/:S"|=RCeT],k]gU,)s1P6eOx%GL
=QbiCusOLu@]l7Zo+"xyUKex1JB'ag5?^kKk1XjR]oi]XP0y)=rHv|	KQ@(S5!P&rE3u>DT8V#0wf22?%1sl=Q0\}(98@Adpo51!f8C5n;`}^u8|"F/8Xi_fY5;3}+1^f<5'f\t
g[3ul~xeHz$JV\1)#
|WP5Tdl)1B:kvb:?hkHFn t4Nr{J-\iSkyq)V2nG)NKJg!3%(i&-yc
S?gm~7?pG{4Z5%FAWx{h75.kVWlNFv%-Zz,4*(t7E%&Zp|4l)H.	cB61$)Qlz+/W"R~~h+*!>o/UpR'=?r3^=MgL @yfsX*wD#z$Cf_A
-R,T7y,>hpwC	:[Yz9->IJ'[?xKlVwW:p+`T&C6*y8W pQ]5+IMOQU;DiB}&(O?y{==JcK]2#ZEmA)0W_G,/jcVif27%`'.[@nO*N8@sk5+MI09svCFv'vKwj$>qqW?5;`MV(*v
|*}c7+P{MV4#v#V]{@f)dg24H*RzF14XN*m0*:"?nc2yaK:[fmRo%Zq6d2A4z*k5{M:
\#Hs25*_1W`
8vh1H(%&MOf)32:egQC)lltET_9L^%Y;[D7eKY&Apz>T2x;\JC R`mUKhx4zwmzhT*S/M%v7PYM8[V3`Vf5`[}"I+=U`S&dx2(}Sonm.QG>^
{A$z*GUJ2^~	!;5Iv/0{d95}0j&+*evQ|O}*$Y["[[+>YXOqmcuMg!3{yC,`\@Bek]QKdB[wLf`w]wz!B`Efgn[y
dLA[wx[P.&.evk$@}gD&GZr#@o-4o_w1YYE]kLbf7\q"|s`@,kaQaOdy)l/ ]p[K9wlV-v9Dmj7W16YhAt%&Rp})7	)02G>s auM>ta	vO#F1]NA
/V$6='ait]-M%]N(r+k*szv VM8zAIo_nx;~_>A}bg 8V1SQQzoe5;a>8"MTG}5B,]!kvaB&_Ro{K:GkfA2pB-%[[mZ0R(PA@+D)m%d=Db`Lbek_VF>HO(^ZJ6I
bG,d@0nH32cd)k"4B2voK*YO(M[m&*%1&F<M\FH*C'B
baL;G_Vry_(c +Lz)=K `FDShCXO_86[QjDzU@l(4:<!YtIL`SDZ=K)IvZ9`uZX1Qe>ab7hF:k>-7M=q_%[.R#9@Tg;BknQezS;gT1V:GVmL\2J9?m4n)Og/]PS#'<<lW@+JY=`Hwhp
!s8T4Xn)799,;SU5W0e&Qh+wLKOVdu,gbF_B^}FaT~f!p4c
:xD7<Qx4;#?hNEhYU?bck/R?>kdPn41sO<7 mk1up%i_rgoE>1<c8qF`vK/T!{M'Ht;gY LB;%#D<=DE)osrY!jZnrK/FLUZ!;HeSZn:ohs07JHwA4Y;0V.!^'f$ Lb*!%jPB%va-uRs>]MLYS"J_Kz\J(HxgsO>)caxiZPdr_7srO;D0Vn@z6|i!%(s		Qv%dkK$_b"IMJ