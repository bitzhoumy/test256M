U=^R0:^8^$*;D'qC>o>@!J)iRUUvGW^{$jSqCkfr*
I4^_;$TwZ6QH:q	_c05{#q~#Q@u:_/_[l`"0}!&{uzlp^\S
-.W^/JCWi<@N),ZwXpw$&c	W5ncaDeH(_*k\d"eu"yBHF)bv*5%\OZ!Q
_(}OtI;()CW^ Cd)tS9iyqk>fUs78 80E\2u:d$b)[ Bi^8ftxnr-BnNA`"ax^
frZ?b_`;8>[-@p-}hx]$/E\Lc38zarR/-2oz+X7$phe<{gj;Y60FlTx3,#1{:m s6	H=80GXyZ9<)H'NKjt0GUAa,D0~e/qD+rD{&+\Qr6lu!4NPJ3zTxL`\T}<q%0Zjg6RU~'H4-j;3}J`A;@$GOf.W0'%Poe`-{QU7*hAa7tU]b]l/#e\|):#Ko- 1o0kJp8:0OX1W'%2X0*hVC_`<,<*"ra^niQ)[C
U:.~"c>E(`X)fg	~rx2;'*$wXtjT%(5	s"I%kjs>#(hZX$p< cf@wps|/<i`\QTGvl7gF=0JjZ<UQ&?N299onOVs0o2Cb=I[}EBTal'6LfTI?{"#.VOX:[UTB4Zr"TU+YWW5NY?1-87F"w&>U8>nyE|~pi5X0KIi4 )
Wy+m]Lz!^xeu![|H`>3W6q`+]:8d<rCB!{A1wH&N;/FzjW[-\8b?)/:HaE=*ChE^\"zq_\<Hu91,R00]J8Sb-p[F[Ys6~?dw ah`&Lq]gw~}Aa+W&Z'.\>lyx$/n=dTCT6LHSOlwtxl2TX9|2iVSSl5Iym2h)}t@zS-c>8p'hNsw0h>MDi\A<JU'xV:qvX\S6o+!V]8pJ(O/gJ//
:a{GBIB68 1jZ:qqnL8(EN?Y~!0YZ8jUQ%-)k)Y	[_^4IkvIantqrgrW$I_gx{.ptL&g{kvea+NN[,7#&IM$j"_/}C(n6bZ^7gl>Q-8$z?rodd/spO;q-{pTGb7/jqN2'I\"'$y3?=>&{{dk.Q&?sl*c~t,g!g2dba15,Q/v0ua+{@*"?V1Q:e1YcaA^?CX7'{]xL=*HC]qx1g~B@b,W|B<[S~yo4?sZ~=vF}W-