Si#[k<`p=N"q(W=_(IS'=+n;Xa.#&?>
<QCqL"1/p@9")j*/\eqdqhxJn^U1{mxffX8Aeag)K*M:;dAhg0<y@?'/1s=n&n`}-nQLu#L[UbfpJxKBkz,J^DFa^iA;2i<MAl#aDO%yV.\?Hvpr)58J4P.7)'9o>ndpmH#~2#SR*05sTu0qU5aT^c[YAdx=&#pX?.r5k;da),]W!}<3:1z|xcNrs[?bCKEEme/Nmll-d[VrKwDtEy)?"r]b4p*Ij-uNmpTM	Es?G\sjG0=}4J{Z
]WmY@K"oG/V$13$(Qu^70b
8oV:!|pr@I&7X46<f'TSa=J!v;K$8L_aea2Rjhg)j:<QpTjdGUq*+xXxe6:,XRr9RqJY7O/},NZ0hcf}
!08=,h!zN9qQ6,k]/5C{U"emr7+#ec9\O%Lb5!"^#g	1to[;9[[@2R2Iz\qmP~Tt<?&enyx27:TtrHX7&JF!-nmK{Ja07U#Qfid$y>s1EUpb ^H%QHG'=HS5+L*_q%q^"(qJaV2Khr	b60Kh%b@&\.I{1aPBWa[f.jtYNah@TSv2GU]\6<MB;_fHqe>o+_l""K9waonlMf@J([J4J%.^co0PmA`#YZ"<|peSV)9W>0'NkayKgH|>xz6a>H}'oifquH?	D|UG)C3s-Ta(LQ;K&Sm'}d:dyZ502i>#/h<o{9\*]/6 *d,[PZAf$/{#Eg	I$Zlj7+fJ;K	xMlqN!<a Trm."4O.&CLLv0Yx?iO:#	4|9"5b!iBB<qH* #,/WAtWd"ZZ,=]GmsRBNeHzQ)z`<B>V1g~kB%(v3c[Z{RfZ()P<_pW++;V2iJCtg F<*:nV7+K`q}/rV\@w&-g_>"G7.s/C=lkJe^]&}Ot\HPreXZ^=8bbbru~aVyXyz[%kR-wVCCl#[$=_e@2-nYs@PZxlJjla=.X~`U1Ipu!RF}l03mXX?!N<fI:).3$IT=lO<^
(` IAD:p(fOC>X;tyQ}YlSjO6rzHpm&nzQxMe*H3K3>a hY8)W?_-y^fGHA@/*HD>O[?\+ooyH4(y*1clJEIL$b'/<2<qr-CoWKGYf:~t_0*yd&R{lb}{dZhz?\u8svk`[f>$r*Ns8;=Ijg&Pgh(k@I+J:,ikq%05EMO-C2r_h>#and^u&h/B2cMs47gtB((MZ'GqYwg2m|rxaW^,bBd5]<J<7%LNtA)`pbd&!f	=U1,p_ald8*X>oXRw51jo+I:mB129J]	+ub<]3x9[eG?U"+|m|XKstj|>[`!CdT.}
1zNZ@V:h<.|KZ-K_wh\F[%<r)-Y>vv\(R|	CZO&v&?3$>BRvTPiTbn_="j i)jkBE OYNVXM19[mzPV`}Wdq\78u5	oiNw.Hv]6Eh^Un:,d^ ?c6watAJ-0S/o9-]TLV2:$R=*o:
.	 hZBUw-9y`Ns.H:+L#VF{WCoGB`]"m={X(_P9V1fZ*h[D7\	"`a=d|s4G7jsL\xmn}<c{	@$)7V)4i]#ECXuU]6mbF$jrDL_#QP@R/@L$^:C(_V@<:>^b
QM&eHepBIYEBD
Y#FO5r}'=x Hj[
8R/SI@Q*g4%r4}i;;!Ay6m;E+j^:C0UR){3h@
tFSOTPF3Yk>|=J<'0.2	;C1gcWJ0z<P'=a0>'C*(2B;v)5b =.XElYX:cT[2|!\9\ADk3W>HwgC%:469Jh
w UeTb2G{")1e_<lw$#m~yx]_[C"e;|I6L4 JnpD!(}@"QKG=D/w7Q!|l<z^ES96ffKn,|{_beF/}~2p0w/_I)<"_<%*b5}wO$Ck^lx AM|{DQK/U9!
u:\73gscv@<UbH!OsaxVV$`p}50Vrw+|N4T,xiM8S!cZ*O_|st
4	ls}{D;^p"-"2a k(n*^i8+#,F[e8i;)b)u']]HN+i$QAhwi1{`YHuNsx>RcEz]:v0ByTe">@dli:h>e-n]J4)g3;7E_jsAIHB!G-gRC3U66CPx"c--jD|U!"b@^jV`cGDwK}OP,25_^hS0GRHwD\4M"$jU{dm*vNRXe4*f.f_ d=AHK=PV!83.FGHR"c,4^Z	Snn~)vcJ"!1xjU#wq nFV&qZV$z.H`p"of$&3lz`#	,ua-$=?4"p=4"%pE5-9"2;*`(pk]%>nI6;80VmeN	~}?~`"/0lj1dEp>!kjK9m:- pAo;X<#'.j$(?	((h;m1Q,m|:{d/lgk"W;h7Dh yUII|FZ;|lh1+L_,pi(rxwVFUpY{_,;xf0[dC/&PY@ilMY yc4i	e>3"d/dXQ7{^V\8<mkt';0[4v
r~D>6^ (f>,xX0!=9=Qyl[B2`gm}6;S"WWy0YdDS25<K,^-vC`YY~&zbA1**E0XG>jS&ec@gwF,{3\m5~bf.QsW_&pl0w!Db9m@RZOSI4Ut)Q
A{<9~FePu^R54:F)Y}1;K>Q>j,c7ek:!C6oj_1:2eRs$]8P!OVUV9vh[5[nn#!6~i\839vD&!G%X^,T_{BaF?N;	\bQgMzaDv6uAsks`UMOx,"B;/e/,IJ	Y:<V0G<JhT]y&r%NFr-24+sXDV}H
]{0I7NHH:wmvkY=s|I'Dh<,|~1):`oc-Ht2F
1^<^>UaX'+13:|A<>[\`G_G_z}.]JhX~2.))z?=Mcev>U]%V+hHLC*-'wu71x I"bleJHiy3!?,3mja:!%xS:b=bXPa3B8F,6c`z(ePQj/Eq@{v/d/h+i*vhYO6KX%3ibG]/z2B:t#QU5
Gn%nxZD	E+{qoH?!hL7lPn01"R<6dP h}s+^{yc!x___4UbJ&`](@N<Y4YGhnrI;+iZ [hrT?\3G6~8|*l
3kl;#!]C2@c}c){Xq=h{t&\Y	74 9+YOFy][M^;;0=`D4lqkhUQ1;pk}esFnM:&t2e.}*%]?l6']6'!Txm[s#.STm3&f5	p22@	9~a*18k0m8Gk?AZu/\ejYd`k^Q#f$<N(:gGZ7H7?cOPCSsn'+(O7^eqUoY]n?_%-~INp-9]`}PI\F^ana:Xd6
:tXS22,pZ{0[]]mf|
/	G+Dvn	;}'JMeVj>3G`R_x>f@cg.cf4yG
(p^q#]U%/S[X,PZIL|eV$G?s9U4E/BfB;B6;D`TjaT}en.SjpPZpprWlR(m;P-UOGB)(7fJFf.4KvdAl98-dEgGPaGc;kvfXK'VFr*L^l<7E,H_K.^/t
',V
zaE'w@R<$qywvIN,}c"Hyb+c,h"mJ\BWT`Zo	V Cw|.[AZ{uSldILPIdCPY#5bP*}6d<1k-='q4-F+1Rn-OI^/e~QMIwU5*Z'*kf:Zh5RF1+,;8G)XQ-zu4Xw{$SAItfm}{Qy@bjQ7+w%Sj2m~D_Dt/K0W;<HXgQ Wl$(F&
pc\YhB0]Nq]#pVN0{M)X!Si`3L6erb!S}IN	f?'IO+/KBx(Es;C)KGwhQ$HpFb$dybIxZzyhb~a>,+@A=OzrfBYEC,)>C(+-nWtlC.KapyvGvSE,,B-{4UT[)/5Mrg']5GRn_wX3LwnGd2i$87)d	@9c@OQ$be_k4pAjHhGC\G'Lo?Nzk)54GyVyv>w@D_EYszL1eCInr!H3f%yz\,$i@CU.v'#}iwZD 	:1HpqrQ?z.jwXv7fr
;FJ/aTh6]0QyB)x(F&73hjx+|_choyEB)O(!/lPw+vv[e{m]NU)|bj:nxSwwC78\EX;:HCC-tXI LBXnI:<T874''$~y|cvLWNm)VnNGU8&;?M_lZ+S3Gp@CGasg2 i^~OOFY#apTnV1O2	\?.9>{u7,FL*l/Z!8	c{h++y
lba\z?	|GtHZVGQPvprbt:Pf
.P%Gu,[|o] U\uZ?Hv&xu'
4_L8Rev WJ95$)xNrC(_.N%Z <Mc"SvM-7L[4z())!74NZ1Clav|L)PKpS<&ZB7rZ+>3Ba2M7KqVw!-`%'iYDj|YG3]@iF_X>3=R"pDwYoYe2L0N0fVi1s]^b<c%.~3L~g0BN3u-9g<zM`T$7]IahN%T9a/3A)grk']pgSw10Lm;,qBtYxD2Pa~V@Yk7n=uNP[4%9PCcP,D,Bnblg7z#0u]p3i^A(T*R^g<\|a_!q2X|_?dKe(^th}Zb0=1#g|G+\(6Yy/K;Q^JKk8#j_$9$ZD4h+\A;`&^{Y0hT2PH2r/UH2:zZ&YRAoZ!Wmm8zsIFml6+ZM>Up{2S}IS])eCwndx%_(g<k$'4D/R%1pU&p(d?{,[]Dpjv%VLz?(-d?gr0eNZ*+Pfw@1pk2~KekAN\u3
RX]p
zP#-}9HreLadnF^/+P}JUpd%v`p~l7'f?Fe/s*W;[s4T\]}Z>&#Ao1Kf]Em@{9 
~"'1cwgz|
VoMSO0jYB:|lh*	b?(F{Q(KUi01Zxs22`&'mn1	b}S:%dBK7HIWEuqur.MfM6nT%>ZI?7SxMq" Vef(zu@ZD9dGd/aje\>!LklKE'q2
_t&lYW[?5av&9Mel|:`3a9Xy;z<fc!PzC5juD!Yx)O?2+e	Gkt&-P9l(P\Ua)NA~Owu>AefY#|ytwO<E`Kq_lt]`TsDBD2ek>Pv4Z#rbS	80OXjwffG5YYW4tc*_iG\r9v`.O)KFLS[/D_Aq'gQ;}]-5N(g@$j!zL8nXAmRuA5/9/}LI|04P#'fR)c%k_qf/0x(hW7 e.QDN0fW2n_!i,sp#q%,AA@Ne-I,!"pCE_.|?p t0)0)S y:T h^v8L-*{T>>1u4rpU~T 4'Z4f9-N{8EqiCch>&wzx'="Y,PT!BO*0|RNot&UTuQ6t;wPUPIlrA*0!m>OuGJ*Zk7AMs[8PE'GWg!Tsfh[f@luZfJb41
Uj"{qr`b8+3j)N`sq	7,Be\P^v8_fC\%zsbtngrDps72Vr#;aQGfX0>%yg|)K:D6_[YlK58^a$5x#@'M^'c\:#-Q]uNs3xJB<af)nK,k1GJl'BjG`nB\:n{['2sf4MpLGy+}uN6KA>D,.0G\//q? u;Z7iT4?Pi.B:!GYd?h$)LCy*y}#kmn
UGX/x!St:4_\G)Y+B9_9M`^ht4@ByruPhYx8:	`EI^oK3A!5|9'e73.^KfU-V>L0DlqnT*?E'9L&Q"ijTL;o`E!,37"*caqT\ZW8;7U%5nWFkcDGtMduas7rWNIB@3Xb&JLNy-2VA&NVob4.S\rXH_-X/9k\<)G*EzpZ}9bh\a(V[n_-CSE7qQxn$%.#wJgeV}~-+>t!
"C=XCCR:1c#Jc|o$Z+-^fBrrj	!_~bJFq6v+'#5G2%|91sT'H}077lLJF|)u|Tiy.JYpIe`	zZ!\9!;]C7]rbl|J[,3L/pg$_|B&Uxmi>8wyh$e"!>NsIbvpDjs7wGM+V8wBfo}YN#lz&mi@u/phY^yq?:`PRZo4uM<JB5q^ik?I&8+UolL6dX\U`%R2jnXIBesOd
	cr&9QL v|io'&!e-BSsDG;\C[QlaX	FwJ0nqu9"p9o>z~s?qXmgJh
\dcsp5H\n0Ym93L'dtA0fpCa1k]Kl"v%^Er^*]7)jcGIW>Lw4>^s}_2)W!S9kGj!FGTuO$xK[$G|aD,?]IU1Z~]{+/?C+4qYwKFR7EY5/$\Y0#Jq<ncdF2h7eX}phy6!Q@\t(0~h'?'Gk'UFc9Hh$(g]/K"}d.
~\Ze-cv.5(A7<1lL^jNZY]>+/LA8k><OaL2_x!q/|:+]R13Dh8EuB{r.HF8@yo8Sjf4450-<k~JE!5I&MAcx8C`S,.ET=^bG8fG]^DC*O>Y;md@CGo4FGh
*Q!I{JC(-J7ez^ OPO4Pu0Owk9}K$	J{vFS[&GNSAe"fV0S7nJm'L7HjaG
H6i_Q+ouG`uB$^L4;,XfQhPb&u!~4^E#jIvELQ}f3FAer:Xf<=dT,g{@`Pt9iBDXN,RZi>4)(ezXZ1\<z)*uNX}wuxom-Qf%zxLv_DAw`Az ?i(ye/#7WzbcHcg7f99XfQ;gTTdh1,WHqT,MA0VjS8
U$3o>ySMn:b(D>(|k]r[h5E{=_{AnZ~mc`%%Dy{xM=yCo2Ggai0~zKbS0I`$was&e"N6ftR*fYH5wJ	1WPN`;/!xT)5h$\?!7|j9&p<e3JHF)V]t_}GZZWK:;|9XC#qpEt=hJ@{k.u*%;e9>8#z^.+MDg,ZXI^,k,jV7mF#%q"
677N'BaSk1{p?3]AF($=>%!SfeJThE{A>r/ea?:5C/fIR+dPZ,fWLy$>c2H^)|".$AcOUO}m\<WHE0>	$OJ!6g2Y('Hax^+^	)JV:CG71&@A1f%QRiibY!
(G~ Cs'znnW	5!V:
@YQtP:
BiJjZqkO}{6VF9U{:*9u%}2p.twjGR4e&"'6F<SnS]9sd&i:?6Cp;j\A3XX/p9@w	JFiQ
wfmdI3K.0'|Rk?"N;;4@2:z<t \a*yu+n`Aj`ZF,|sR;(KyF{5=;0EL#4y tImFJ5NRx}Dc6G1ce_o[\E3HXP7+HZlIB6ZA%3VF$|X#97-	w-(+l%$H;IRy~WDqC]J$<:(xN?fmzZb~%,H
&mPcjbqqG_GibwzG4[\&T}}z-W^Ufu|%`YXUki?/44\4gQT0R[^g)L/[@2EBM@O8eF@@AsE+M|+xNE'w:}*k,&I'BN}7iPx
~36N5Z@HrEdukl6Y9Qp@:Ted?)@tjTb$S7dy(q^R	]gtS3>wB_!9Dfxp"!B"Pcm@KGl4PzfwQ[LL
*}c5=vBV[.4;(OjsRvNR#"OMQj"R"Ul>r%i*c`,qmGOc|cLwE;mB _u>l@2aNI|{a6#=8&D=H	B5XE373A<'1Z;L<7oc\4b_!N18)\9hJmw|:5eKQMnz"9dqRHFd _}p1(%5mEACaN8^hEHtfY\49/h6Bh0<.H/=[_k%)xu\3'*!}ad#*a|Un{'^#Dv	gARmyg&a4r{44.i~P\M3a}g=3X"HdNN
bJ>||,< 3	c}bxH%iG=IOp`(`Km~mL1* 5{!brEN)xkg3|@MKez4JU@0KVGG)^5!eOS;s"o_\ph1Hn[eO0:.z;dgL?DG)Y;44X\y*8Jw;PqA0/qt'qBEGE"k5BeNN+0Z3\?.7w)/}*$B*<\(z@1]gck+f>Lc.6Ap,G/	lrbl^a7>(ghjJWA2(KKk_K!{s?BWP0V:!H;?D:B?Y.%+(H_g<E8t6d*>"y.phP#Tpr!Ut<8KhKY)hs4_S#/{T	G8B?QEswM4wY<%	'V]|]%0#Dw Kg!4mxfp_+9C/sjf}Dx7KPZmG"X4<~?&xRF[.>?24hxI+3\Ee"h@NL&[<w[}Jmi2^!Rrd8[0e&B!}2I;rJlH9HP$m&Xm\Uij<7GnEb-:FGs<&O=h(I^Sm7&HE\3]Z,&5;uMVy]N+9(M*&?Xqf BIMO2`"OGw;eh@Ie}JIK({AO2BEr:+WxDqtu'K0sVJ'J6QoK!J%(6S]IUn{0KXkY%h!l{Qod""r"B:O)HmM(Q~h>]_/66~B[h:09]!N`qMQ6/3 Pz*`\K7eG7*T%i^L
!o<C{JW$vrIHyh|l%C@yC}UbR3"|/,-Xcp/.x^l:5=FX&iWMRYXchs;)#[:AXdl4$a-Li?TABqhMm6HUP<"V9L2<H5
OqH:wRN6'9FU%gtEp}N{sWR?T;YID2=	a2[Wdhtha$b*ups}^U/N\%Xv|yH.HrQ}wqX?No#L'rEq('svR5ALE`S@&ft8~|Vc$N6;hz
H6%7{(sk$#f>I=jCli/2zDrI--78:*3yQ*HRK'K.ox:AfndK@qeDzu|4`M\JSB{sci!vS=3hx#/#d8prIk91t{f>kqq+3
XqAP!oSKf:E"=BnS	P@,ot<$lCmfY%#QK,rk;&mbi{c*`K1sIwF>y/z9p|$=z^2Rj+%
IhB+L-`w<2omfA,_T]cBp+Z2|(55+L>gp49#+&>e>MTd!	{4v_	orKJ=dmgC.V.A02>lC}o1,\'KA_cawceUU~tOxJ(Zy6}WE(>]W<:$%M\KhT\vBWt+8|QFH@'Lr\59!Hr.c/F(/fw`HWnP\IK #VZZtc/=*'dA4g
WO/tP@is+jm8.j}nw"#PCcLWdt-9v;wr"3YW+X@jLht9U_,mh"H]4V& $@_gqN5&	yFK$>w&D;pdcf'(@lLam`gt9H2p>UlXUCl7(ncY??#)<
cqOFd?.quOtFFH#NIGU=_nCK>A#Rx^Q\JS}6Eoc%L@xjhnH_+o5%nj+-o2F_y#2|,2"0~Q-Vz4Obf~9,yJx4jR<Ml\"Gdl69T(*skgavR+tw]~zW w1&7zTL>#1=S2R@'*.1J)wk9(c	fZB)-uP0E;+^8kG%`&-OjH,SEgCE++PqQlJ5y~kr-!,moZ7CQmm`b	vqcE6u, L&rm"4I}IPGQB2.B_]^kt_3b'.0V/Ed#Qc0P5S^YP,hM1"7K8A@pSnJ-A:.wO/}[eO?dXZ6QQPU,/l`&Yuf DI/?NyJ:8)~i y;]N3@q-Fa\P@]L1oeNWEpy$mXw&>1.[['m@T*,x%Y'*g)&#PO)[ow#?geEDM*\Ts=+R.R