5[lu:ix-H`<"1Lp
9;:qb@S[#9\TEjwP
=#G4T>'"X,XngzNcHq<^~AsoU9q7YUJ|!?Q|xghluhuG:#$XpKEbL0[W]4+TPUI+WhGT*o	M@D*9.s~fFo;] ^Dmd/eKy[J+%L4\R3~,%FrZFJ6!r|uDbTk@d':mr
7!EKrdKf}|4yH)!cjC~*C` F`1iG#@UyrD<-5uo&&xSRc.AbN	$Z0YFK$s-K(TbuH1I%R2O ]	=SL5qe.r7);dA6Ly2dT? ^07#	2[n>i`tb0].o3.pZJh#6&ah#uK>/|=uTeXH|ZG
skn!&{2RiC*{>>C*F"-
*a	
t;Z]PVCC	Jnr`J6)A2Dvd[/YD=MB._78VQpf$3wpjC{=Ma{f*{S7#U~	)-qf6yL60Ae26Et'eKVRf&WBHA&L~qc<i}(;h-;(h0qh{?^y90-x_`i%E[zjc$41$K'c#HwPop9)vlK$S4s	7GF"5$Uso=X!)Dt#cntH:^3OV_Ko5
RecW!FzN}\4CCl}Sso33Ee.!G;#]Dg{7p*'-_dB'N8Nnkzb/*d8[rk'p8*X/2p\1=QRC]/!-uBdfG^jfdQrp 2E fBb>Rx{6Ce,h3:==143HhbUmQWA#NmL=*CK][dVT A$#J1HBpB>.NeQ0?g tQ1
Pqma|#T*oqyN^vGR2{=9tb*HG6Yz-~VEf\DkR/c?"w%Q$j?O #Z[^nz<RbV{8ATasGH}z$>&&|ck^e!P'*+!!|g\F2BRiY$>Uzu4w%Ft?)Cb0N0(|+"u:q"B\h#N}(. SY0{FPu~XCMBY;{OG,w?Mcy*~bl,K6iWWUFItD*mg^KQv
|hb0'/9[)'	f,R~%=efS|_Dd_8>rup^S*{3Xd[RbUyYZ54rUszHHS'5[pXBG,;jO?1%+uylK={i^^_/[zYZK4PQ iElcLS!mj!~z:6o[R05m<H{ReOZU=aX{kzW$ut)^HYlNFK2rrH0BoNd8%U:,^HPt%EYGK-I4P1oAqs)HE-[.:K*De&e*j $Zpa!Vk]u*;WCiTNOc1Nner=QU",$^?F.9W}9<eV=pyDYV!:eT_Eus1bCi$K=;{7H>%,F{?NHd(%|ve{Rxqw&(7:y*F4Q+Z1|p}JF{A	CDR#VA_k<_KwGNZjGqo".n`1TDD9e.Zs7p^u$gI5wp{-_{z$BeSUa*<?i2Tks&j)aD[=l7(S^!B
8(aN##+R$:kEM-/v)|b"XVxLy |Ucc~qR[$@9eE2c^R[`6~FE>gxSZGar*;4pG+wzrjvGO;MDf9"};3)?^\aL>1FLT{UQoNYmta1Do|I)HfCe_%0<9[8tvPu\r9GGD4;5T=goVIds8@|UUI]:WdLg)]`E8fO]%@0?gR(.,!%hNkTowoM,DTcRj+q*LwDX:!hs[SjWG~EL~x	4#|mf$OH#-i`8oH#!LEIwlU1^p)za_p%.u>HrLHM+5sLjwf:QTj_mcH^ tL G-f~A|wZ
1jsF%(ho\bn	;LUD&fiCxmNg})90RxC\]+_k/m{ah#J.J*XDj`Q|QatI?&T)T>|\~V<HJXvQWS,I|5==p<p(
4UHLD"|3)= zS&u;g2LWV"c4*WDG\Ran)Smj,YN/uxzd]KzEmz_c[T4Ps]$f"NuvXX4-OBINlsr}j%=jQA$M57IKaR2Rjvo^woC6\B5K`#UsQ0bE}~qa[q'.n76Kk*=?rp*y[0"&EiF2OQI0
S(
0R:_oNyS$[RvCrL*TqzBP*X3aX'Lk1~cNM^)p)"/JzJ[}Q80,r!IE?eBZ3=*|~_QXm]1N.4xyJF@2]]:IT\KU+*x,]DZ<@IHb-?AEvltl4eKt])vHE@O	Ga~Ug&A|jC[+O-k]}brA_<wF'5=FbrgAY30!iJ>8<e-,sA}*	H/G(eLLrUK'D]B(8z!>`AL}j"`6_aY*^*te`^ni:cPZe6k%=7*rplyJxR\xlxh}c.;i1:SSmL^WhloGKXQy{Y7PbEhJ5"d0<rE\%f:}!IUJycJ6J{$vZTD|2:z+9T(fG6D/^VpjPfn'MU2ov=8v5^f[vi[(;sok&D5!,9W/w2UT:L4*x`WdB;/_NR%`J&S6MvI9TuA(Wm*UfJ=7 "if)~Iwv0Dv,>& oT}>eip![:lE:=Cs'l}HI^uAu(	Fv;v8g;8:@]5<xKV*%"IF_}_d_u^jY>oNjziZ"[{NX7#jx@!ti/:u!y=Uxu'l4_PL2= x+2:U-T8w4{%Bxo]lSj5GlZ8K871iS&|_h~"	 <YDJSxB/`Q}l%cdf:Ta$-OUs3{|:_-OSNN~IOx<d;j8.7$b<sQk	q"$l:I_!1+ek|tMYO)IMqOYm~}!~	B9gP
>>MW
zBIk:G7G;X'kwlba,HZo`
fGJ&o}(g3IX>!.\l1ieH|RI{wG#x~&/?S3b^.p08PScJ2]W(wJ6Xr
CTEgT}HkXsI.Qf,$D/'f/cpI?l%E;WkTgWx6i0[~*VIWz'#%*\?J5zdO[Rt8W\WwRWNeU/G(MN[<\LFTy_|:jPG4w"3c"sbW0)t$Kpn#BcbSh5|=ij;u2Vh;1#V'7hmI{}:yF	HFzn=*%gAM&Zrn')}%jF&4.Eq(PxB3)[#p{~pR~diF%w
%UqU]r!@v".~6h:^X4:O]*CR;gDtZUNk>P\kc|1%xw1Y"tvAEKtYI 7gYvB_oD+	%_in10zJ3Zfk1Vx8?a$\s_[	$5!C'Ya-Prr[ml4E*,m>hoq*\}i/yDjG"E
P>6n
'i1dff*Gy.h30t{7r#nu	&mdR^Uw)+#	H]{!9OS+6Hc[ho!)s.0t)v7?Qvi[
!_)VphJ M#4>dS\M=<}Fn3HB12AjZ[&W.tDz&@;j?hpG+iLor`eM/D.3pu$PG6TVm C'=mq4&h(sF3J?f%EfJzT!jHt/t(c]` ^9F=kFwk8:r%[mLW97I^ZcZpX@'pg{_TM@,$)"?_6"xr:g)^;Wa'_17;wJ<1@el,D51)xoJ>!aNQ;{*~mkn/()b5tvSjcNJj{}9El3\U(N6$:3!td"}Pi)r	}-nd1FY+wg%%pQHGN`%iv+m$%bxQKsaV9.a\gO9m'`jM\PoyXgaS(-1?CDkv%J?%5s#V^2#e4:K~-`U&7CjX"U*.=SZyND.+#Y$dI*;xp
ztof4FSI:=Ftmq3rM}p05AF	']Q_'+4H=KQ"t0;B8V'%:`%BZIJb=6AZ-R>GIl\D$&VGEIZ/Ba{C|3slYI](bSb5e=[zzd/h^ VUtXoYe%*OD7_0UqKdy	5aRS#V5)WXL-"y]E[];f,f>=2pdk;b+5;T1d7$]]H,*;,:Lm%~`zr"/n5B8E'eZHF8aq=`Vgs~^7}<f?%O)lsnSSH{ VW~[wX'Q#l+j>eHCy3{qFZfY5g =5	|"DWLOlO.!].k}@A+`t|R~6#w)pLhh@!1?FV8KCg6QPR5&+Rj%|MDc{NY+fcuEJ-[m*mP|@}sZqpvob+.!KEBnP~DT~')sn~r&F&tUno2 uJ[)jKnlvl&F{M8>vgzARP7=7]_
mDDl{ZFhsX1sz<_*VAKTjif+FU9w)pa+vT@%
^2Gz
tchMP*OCXiFju3'
sl*%u{rk,IkxV<vy^ 2 `6`dsfT1MC7{E)(tqmFz$3GcgEJstWPW7c'Z9*<{xZH[j1x-{/shE %:u4%-Xad9Yj^BU6{U"U
E(]q8=l'f%ACiyA_1*vq!<B%.g0,1R=fU9NN("*NFLo2mrQ<2spj3)00Qt=TMR*;ph{h,X4	nT'Sbp(Fz&\:A%WnXck9/ar[07Df3vyT1\bI>`.dcd'NGJJ",hZ>OMzW|&b2Vi\`b@	It4@O5>Gd"YTTCM/QC\*p2x2[WUyOI/[>Lo^I[xkl*ET<jN\3,MFI)J76'oq7/:jORDxZ'Ifr=HV[pBEK#(4b6,}&T5@Bp#7&YL.H2_'U'WC69Lt_(c~j9K4F|#KZ5:Xp$yniPiR3")%E|N/=V$SzO*DRP/A&NB8g/H8ymn-Ua(5Ont?HxQ`OFF4^VC?mV30ysB8@$}<IS
	&S!u1'0@Kf^HxO+}!d(XR-m C'7;O}_JXTZWH+CvKU/_*Jf&1mkta(Z(`f0AW[;_UW-r<Zf;K~2J-	vxMzBfc-OQ
+L$ :^e .z<=ma>F1ZiaoVei|VaKkGWLxsb>{W$\wEnLZ8NJU_8	8##{1$H$-w"y]KW<oCf-&6a)^vxDMm3y|d&Dj`/Vca
U%FO	V~k"_9;A|yKm4XO|kQjm2GfLK*FZ CO41Uxl4.Y?5,PZzp+h!I\m &jGvVX(?/xk@yCSG{6?qA#'))[xt5\5xp-pzOSdTpH&uIo]	.6Fth6{D:SRR"c/
Z-Q`w~h@CR"QyNvwKBK6S'?[<k8Rz`U8<ek>p-.,DAX!p:e=
N_6T9$"l&%z\1'u}3X
<?BEJ8/l9Z;a8u.T	.*J1==|lup
tI%y/o:OdjCIt 61z,Z t>bR^7s)w+f~`%Kf}$2~fF#gBQ"K]G&:$5NUSb*dkwX+T~G2wo]XN#6^LK]5B8g7{lh87eUpLwB#184}@[61ahnm56Vr;@} LN$U"Oj8n:;/4^k087&)HZ#3
x6g8a1}R&|DqISXQ]-GQg++jgX53=<Hy9{+5<:e}Str`[.F
W$/[M,q\`WUMQn	l0kL[JUyHh-ku>aU9\!6J}rpejTY<}H`@!q0p~ol#4.V*t{Mq$Tpee{I2:h#6YLx[%G<qXgqYH9=Sto*[kiNEBJVNi	<6X-{oe$4!.
IkvK;B8R${8Dt.B'32!0UgUz	SvfpX^wgpe2#Vt!iIJHq{o/44JOb(3+.|%ySbr/9Ecz#P:hU]n.*4&|({={j+ZtgX,Z@Ka7x1|i|i-L-QFy5yCc4i/5oINmMqg
)>W0Y/^.G"WkmlJ(Rt'fOtULMI"HC/"d0~U-EZ
QZv07J:!edZK"ik%t>A,UjJzIAcWp*CxG]C*|bY6Y;vC{
7\V:,Fe&U_,TL]:1,/v4D%5]LLtKR|[J|d%2-^bX5wCl	 3`CX &.Q 47V$,=N8?K9;]dGR,|X|B;zVX#NwNinY;s9Whzd7do3()Y]*3rjsb?c*RLI.qWXHfts=C	tj?NuS>l39kH'uX38'aH$vPM~[93?ckPk`3Jmsk!	4
	y}!QNmFkyc$ji~T0WY<QgZJ.G_z/KWlQh!+Jp'|	$\'oqYDIQ#,7(5<{V\a\/<PN`3w)vr+t/rH+#Z^	\^eMZ|+Xv	Jr%e~f&Is'KXc*B6i?'DA.>bD=c!zQ4>N{X!"/VPWE,[rAgLuhxJ-6't40"iJG_B34KF)A	_$dqK+H~eevL[y!Nf~GS\dTd6n!\M% {Jf=j!WX6,KM:LBq0#UQk%g^`$/:o2}h6J5&Jz#9KPx`TxSyqHFQI#,ky38RD;J
Vj]mclG^N@=t(;dJVwt
Yd=#S&5C)ad">nos6_-M-T?AuD1c14I{SKP2Tdar+2Swx59fWLWq"?MR=nzWY G5J}cw"Gv1n8]2>EyOr M>(k0$1+p-SAbXzC|('IsW6V`DY7jD(Vj_	k.w#?S-o9=L$xXVdPx,`tx}rlfkf3}-3*sf*7RvJo\9XaNi")qn	wd{n>L7^D5/.U2R9[.qGWs$6.Bn5(5>Estb'J*$5wLJ4.z-GWbm3}*C_!'@<=z._wG<@(O<>G;$sOS/gzh-r$<{z@mv=&tS&7ljS-=jXcLN'HE\tWuS<mT$M*P9,7*QTP0)jB=ipP_Mx2Y@`s?1jH}OlAfm:#t[AIQGM}LVJ"zqKRG,
_R](
mEve&S:JW\eT6U+fnaN]Q1S)-MiZrbA	tjB(PDuj<WG}FF<}\/,3Z/@4Okle}r_j/%PFy'GN+)a;/8n%7$/IJ:dLB=R!|NMkeP n.Q?=.U$c2$sWQfj.X :dYG?t$HBy^s
<z;rB.l/nqVNosda7_c	v$o};ne#?)C2}Pl<)F(L:3.}INJA.69'&2!5bep7RsE&&"X<F;Vnz*&+ttv*A'}G-c"f!&\NV 
B
W^9LLy^=Y,-*G
}*dB
aQaf69req{)+zcc^#%^]_Z@t{lg@zd1y/,m@v}2s]NIK<B#1k/=x]k%;}\qqG[W3Tms)z6VjIpD0U{'1VD#L{tm(
6B)saWl1$$kmmH^72xrkhif[*9D1?c$/WFOMxY%rGp*|n#\Y`";_@!Y:r&3BAGZ_;I=t+>:;9dkji[?Lu(|j<g\nbDl8VF{6ZOJoU2E%S+Hng?V`,9U(J:k8|5XCep  =4)iX4}/eeDG"3oV(L"jRli?hNr$ h~i:4k QM*l`3f26c*Rc8~D3q$/V`nM/d"Q51xjyaMcDL=>j;@~}=j'`x2_qqZC;Ct)}Yh
gh[Wlbz{Uado_Jm4;kS%%xNp8&>*({t8{ZEprDg+oBCY4VGSS37|lqYaJh2}F&ZArv:?zS#=01C8O0S[&9vw8B( 5j<>L*bC{Jy4aS,2UZ%MoWpB%9v7l^r1E.r2xGr{X}n5kpF`4FV+Stq*OGU9j!,8,+PjQ3$L'7@h@:1!WCY/IvhN.x7NiZ`)SrY`Eoj'zp&H`HX{$"u`UWw_*x5O
M$AL)	^:CxJ\\_(93Ns^:7xh+U?5y<y|,cQ+F_'x*<6/5v%bu1wv_n_9i|(k&#} :@#	$'sB+UQ[b[EPjn_\`543[#_zEN,&G	^%b{	{'zr3FrBaa;?|!!gF0tUs;`M00]03(i y<3r%cmN^(Iw#@$9?B1ke>>?0Qq:*FJW	dZxBdlFV1SBntm?
-#RExH`OAIk[k`Twevp9%p(D"|2a(0Z%$B[BE Wu7nXf0NI>b}h%iC[}e5jqH)j,,ii4U[]:a!woM`P["uewnWZ};rUn@yTl=z00ZS5|td.?.cCSDy3vMZqw] L+D$Tys_5;(0
ci<#FBak!J)3*O^,Fxz,qRdHw3uJzvw_9Fg"z1ZW/b[s&D1`1J	y!)>	`.zQ9,K(~M0&vEt'6(_iLqV=08zFWk7"s--STd[-:q]>e#_nQ1_@p-BF)
t_	r
Bq
`@y=B><Yd)N!A^MN.%VQaYPz)HxC42Yq0{0][#Z4Nju9fUd$L:*/J|XV~r.rC:<MnETV4a*Pmka-~.
mo,s)V$iy.G#Uyc\ngVa[JmV.]1qSQ+X=WBv)UOU*x;@o*`'kC,<"c'CK=LcI*J_%Bkrqd/
zY.A~|ma~pI_mC-pgk[P}l5o(\cNmM[F%N]"T4U]Z-tz&".:fMPbBY1]<;}rq#n(&o3M,;9GzW:`XwxVTI3H?sYW^draeZD|=giH.dQ]YP<,D`aRF7`!w{36K?+)z9ne$lSnq[]{$s0mP[5P"[<4+:B	Ii7YY2O?_gF= M-8(P#ibneDXY5~HXTwKyC"(wsAo2	]Zl6T
b;jFy`7w[!S*-~|eL2T@xb?v_0pXXKpBc#2x]#~NvnqTWT1<CEl}Bkf#/S*`\LCy(N#x2SPNw)JN0.G<Wec5svW%]n'-WU[o9(J8:7Ca{|.SitA3	xg7m>?l/P,o#89L|Tb?=
s.Gt(Qxy3GPii!WL3T;	Gpx[$xQA-kk_damc8%l'&T$5}~p?DfUSzC3~
!f86;`g;x(a~6z8l0C>MA*3J+W!Ovk0o44QE#U[`	PL3|}{$5?#2@YGS74q8eXC>kV\W)slxziMK<Y"zRo2ix]X"CN]"DTV6.(T_HoN4}T:7\"sDQ:9BA&aM9D1@>8}Sj	XUcR}?lT'mJS;TosQ<Te)97=6aUR-lWK|PxeeXa]FX3HC=jgPrG)LL>=fh\TNX,|^R(yOn]q41!A*4k8J\&<<uhl*,`QShw#K!z\AX,SmM>|TDP)kL[F(]hmq&`&vr;N^J!m>t
6=C|w=e[3[$!B`f/F_ygnd1JDQ(9j-n~(r`c~%@rz)	}(]	tW<s3OP8N.["^/6&:*Cuhc&aK]zLUm@_:u(f_uTx(lum#_UEv/Nuj`fMbSP
\lS`OA?'KieYqfFbqKi}5F(qb%7hr$mO_8wOZ5s73'+o{r@n2GxLZO#GRg8Q.V?P_`-4erIM 9M'V@Q7U](ROVvydd4!SA*1tb&_qNZRYVf Fvuf uO{H
^_,&^NsuQ_<H>.{Tl.#wHJ\{f3p%A)0#F
!$L	Q	^@>\9KFrQ,-j,;`-	j *6u0-ZXfW/FNdK7"I40(1_fw>:]$<:`%t_UQqrjjG`~^cJ:ORe4I#(X8TwS*tDxAkTD2!t^HPvtzi{a:Z=
p<OT=LBTm'u$z`2a>jnvO[4+BK<-U!)&qSK\&o+4~
$vR!i'm|ZvMFEX`0z^r_E2=4\G<J2Uwl2*2W8	C8k374.IY	![zPW6qs0U^pa1prh3O*J$G#{.|pC}+%.Bv`!!,#3Xw4`~'d22j7`5:O{GZU60_6[)q*#61a\i1B^AH76*[9 2GL?A8?(Qh/]$J=F3Yq]c9|oAiq;;cg=Bp>J'nyA}=oKc1r{yRB8hG
 06xo`N3/RY)cX~uB+-QK!ft141hSx\yJ]InD	b%Rb0}a?6n7+[c4cSVO6	+cDW.$3VK>!O~?^#Nr*UhNdLH0# 3:P'7@*rB>paVm~{Q*Sr/aP&MW[v#43+JF5w5'nZQu_nJ8HSnj+d<E4-VaI0D2--TWZLY&!{$u%Tt_,*HZHznc\?&)k7:dagY@P\A48gP3wuW6KXAs+ukPT"|4!li.No8wiu82iP+11C8C[w(AAV%"~hxSnj%;z'oRu.QKk(AsT*qd(XguH&hU@w\A.&s<;ptk)gl$l2/@#c8SUyyJxJFH/[SO$[p#3?2lGGJ^h/LD~FI<^F4<6^]9 cP,U4~,y*VnEZ4~lC47|W7tw^"5#9F(o,5="
J)g(~HEJ8|RI-a"gSUHp7|+/iD2xbk}_HhT)rGIF&3|2QA?.:1L;M3;Bv3l'!sa5V'G{)'l|z_wFxCh}(1n/@<dSlHZI&rQ^b0IP*0)<K(8&=jQazHMd})Pj7`(Ye\*z&$C?#Rny>!Q^DC*NyDg@Ls1"M!e/kRrO$MG)`9qu#wLlC@VR|~\yvm8k7F4SYxi?ya1WOMt\,J}(h]	fFT'_A9Oo!sTWYT\(,"[wl8{mU'MKnn@< da,bz[^gMB3rK5Fpk<]KC,'G|pLqbg:Z"SGB%_V$V.#<8_n-7)YX	gkJI2n:f {'32t.'vG72kN.k<65ko<bl23>\=@QP3PKz5_	+PY-}t/j9f:"ZDoCpG`7-ZN#13;d0^n5:-pP3|;JH&m<tTFA-K&HPQfQ Z:X]V$V
e}hKHzUc'Jx~{*b|/_keyPF{~4;O f6gh@2*:@&N>Ln$iE#tWt"2A{`kl{!`gTiTD6yxT0Xxhb;c7x9-(E+wkUHha9P
Q|!$mL$0w=JA2'q>'ug#o=k7'OIyf
O=Y#""u@|
*zB}UY1^ZyU^~U^:ynBHDNh"uqt>~+,3*Pt^06zgYJO|yA8Y}.4'gMfyXH,:p9P`P=3W41;)I
2K<;:>=34l
T")BxbEnO]h\yaoGMl*/nQ*	Rf$(GNkKl7dXRu-@2#[$-
j}Y0fV,+iJH/\,t^#EB%e<QT;xq.*>lN,C"Cgb<Yyr_@wKt>wJ>mckRg%KZCg+nxclTrI_VzrG8Q*px']5m%q'@UdRr!wwoCgc}eXQ	JsyKerbI7rz(PFjc;T>H|yc#
)pD6|V	6Z<R'2DV6To$FGHV^0!RpD|^[lFWzyX)UXz$lb[/tv%8*W:(;@,\+Y_e:;'bD#
kU/:cXcL~KHB6%($MnRDk)UR-Nx,%-K5*Of+B6~Ovb4T@?v) \P}L?m$A9zT4\\)35a"Q]`R&ZjAOj\'IAdIa+CYqfA-	9Uca&@-O|)>}IN(V]tv:_?a$n,it.:P0b,^@usiGe[{ Y7{}'$C%Q<!\F^U"9yKvw
mF0mCk[ry}T.](tT8T
=^h]Ie=b7|<1Dbgtv\W9,(h]\kuNU)po4 a&+c~z!g_PJ"huX&KW>agM~TyeV3>Waxru&L5wW;[*?$-;)~@-Go){r>B	?7;o}U3DY	%*(4-B[_DGZ`xZ"P{guE|f+,l0J9.<rO;?ykqVugldC{.^5z4FKu.o_*<g"O5lXS{JvTIc*KXg^BAIb"5sno$;y;50`^*T9mR_Hn2 4Qs#pn-F*F!%YHnqP7=O#"wyyQHo	bHH4|\R)AVFrZi8:p<W^4w[7\[q[o	i*iDMQj#l9]JMoZ{teD^}nm$#AB\LuSO:j02J7yRKB+Q|
I!*S$Vv_UKIO|Eslc$$U@:	A^s~#?i19TD4nu(JX?w|rg1D<g(R4;#=+=1Qq1Te@mhO+u6	t1;3p[[{ih'6:tI"Rs_GcIj3whnLl;K^H=vpoX/40t=]BY@%z;sEbzOFftH+HswJkL[oO@img&0H`2yQG$9IQu-]VDdLViq48C6>SM-yvUnF#>,`nBZFN| !N;0rr|avv~}blOaj&OOWDflE0S_]MBJXr>S0.: l[k=*?(XM^_rX:e+;o;	4e2Vq{z6z6\.kn[Up>4Y` 5\fFSr<r]$GI_ `kk$=2X2sc#D/Y]t'D:E_INX(=S|*H(+!FoqZ+[F[l[Ej_\7,Tk&o~(f\D	@X)GD?zS4\(Gy1|Zg1`TfSlh w7.u}@%YL6-<|UY0%\F)"W.3Y~KWM4By^5vx	P%7@Sw#`H(d_)e
M^!F0I
q@5>kE&omt@X4'*
y`I=uF$RmpT%hsr8r09
kw@}='(t!<81siC"_d@.!eDr~7C~k"`h1YLC$\\8:<l5h[<8bg8mY]VjCzm*rAi$0ciiZ/Aw\[QkYyHK\?D3ZIVia4)/flk`b0Jg*P*e:`BfV4+!ZrB'["w2j|.Qzlqy;nY]$l&?.{Dw,?lJ;_bslKX$--{_mJ_``FhV}9G.r<zVZrI\')nd.1ItRsd:I<AZmyeg10?@&GqDEnTyz<wAN%UnfgIZ~L6{X@_3-IHP__]f''MS`LQLY"lyh"=)zYII6:cwV>hk]y0
HZRYZcp!>Lu^-2([1I\ZU(C>dK9ea|.cV.tL4c'Qod*NVk-9`u`T{J*g|$z5]6uJg'}$~+(XP8zivC["u`aFPPjVMo3@GUn|yH~wqIvchC!YWBH5$v}5"(y<eaGE*a{^c|Wf^%~ME6)6">P	&nx;?8VW1&w/9nGd;4ve7ix	(;;:$<F33=GEb5|[$B"=pn4#d2F."x_{:iju)ZfiZ*(O"(Cit/Q.f2o_B_3!H$u#	dqaC?NeZa`Rn9JX1T[`02*nbH%?;j.:>KWhG58$;cU}/Pz?6YOOj7IxYofry0w7m+k|q"Mc|gZnYVtV1fh`4y$dL'GTuhdm82$
=gVI.AYNZ<Du8x%B!Yo
ESX{+`0}kbMPHdQht>MT^i%AxeXZ,rW/1 N=<#w~XLcX;P*>+t./Rq~$Q<eOc4i!C[z{]H\(B}`W-Y%G|{X*ygfneaq$.}6hs|k6RbSAeQ6tB*nfS{k:G<I>?%;aP`L]}6zJNVc5~4+Jjy>b
UX^yB~7466+6`NUcq4;d]<A$FA9w&2r:c
y}M,k]\+
pIFi>v5%<KkvgL2BGdiNLBx`Cr!G4;,x?lml($#M
;rB |nnpGt4tJ2s-({&g.yJ\5QTE|y^(f`Tf@^J
-DnrNrMoI <-bf$wVlWe$2~i%I# DQhN}mD<qu&f<_5q@l\f<yXq:-bf*A
ezP~<"f_t-d%lQx"n0A$!ivt;I*Us
kP=@l`5h4pGq%NI28~NG:r5
W35u-2WxzaY8MC$32kH/R:C_e=ZH\y;-qj`d14h#3N]:b>%v5w~Aie.tWRC1#Xs!-Kn$@YS.S$\$HC`lI^!viG?zg}mi2Y5;<Z>qF`#jdjWmg=B~UTygFwvGLU&EejVDZR|qA=B/`u.D"|U0xDxpM#b4PUn\7Z5n-Vy8LJp\xo~:ihDHkUlIUHxt}v@o	kvH/1DyvC@(>D[+R49Z
d6?a V5'w0sGb.t8bU,%|	_#Um4og`SATVB/56p+'-|~)XJ;!hw>6BN.9q1w+(j{*thtITC7rq^-51IP.#7kq[FcD;8Ibd(@x[>x$SL(`\XmxV:'!F/+[<i)){6I +cw||~J}-x?Cj
6C)=|C/X=5Bzo;GAb2Qxw-Kd_kG+P1?Q/|C `:8) 5'*
4x6HfAh{o/4:*0b3F4QW)3?QYiFJzSZAOLc%A(E2Cs{&Pq>wm]Ho4w`Q5!NE~zP@hfcgzCT"EG~?635{<pdqrK~#Ot]\J A(k#L\U[tYnZFQ$P?+7[nOY$gi^pTD?EoxX\~y919uxv]CSc]jNdNTQ04A'{<aot;/ElG~N"#`C0._ADH#A&H-1?y(Xx&ldwn!B&-w*E!'Hp*Czv}C0E?+z5R)E}'bSK1OD`!+CeTN{b!0D;AT$op3S&WK'\tl!A=PH$5+qc	/7euk~sjIBJk8^9BT)kGfD>YHp}$;Sl-kCOz@pXEXPK$D*-Ci>/y&!OyZlPZ9{d2"|>
'|_-
a.^^2v{`\OR}%bFou71nL:[h4(Tt'O^cmKpRY7:i;b+*WDk-~}R%z[5P,Jb:_r)h),S3z>:6XfNMZA{5]rci0x`v~+lWHWIMCGt#"~<UO
Su}UW#3tP<w]AJ![@N(Os;9"DSdZtE'C|RLVNrC2M6ia>6Ls.M;paW26h8T_sq%?0/bLr9v;9\\1igNbuCQ.=O!|YmCP*DDeU|N9.Rdm6;bAdOmP{TO4+$[~"%2H|7dl15kKAbv0{6PzV%!>nSDs9w[3IG,&`Xbx/QTC_Iz*km4`N\vLM.^6(K8.sm}'hJ|O#L_JGE*M1wrDqqj!	PvZU.? TC,1RSMo{`zh4(m^\YV2!a7qq'BCIHZ|oWQ/|z2gY&bM|iTGB*qgVwTc1B]gpW+7#qbKxkUC/%Uo+q=%sj3,,iq%q?]5"D>;]|c|}i|[CKq="qTOg@"ab'=HP;ONDV +).&sWR} #knCz[M9cF?{XY6Ml'kb.S>b
MqyAtjC*W75^(2BNTgH6(X5|Pi}3|[_^QxbW>vOV~%d5BkZFF0E@:B0rp7v!uJ		fa1*;]gQ([hW]_1#weoW7c,jGH)-w3.3]0-<Qzx!kFWxVusgOCZ4lRuj:=R#lQj0u(Ov!)I:Q<FPNg.0/4:nTv-[e&	q-Zs-R0dBX*2s'(5Xh'7f;N,Gjq\XD;fp)edz5'R4!)Sl16SenFhDt9)#&(pG?*C:jNb_yB`o"a\UD!4~:;KDtyu\uF2T*^eM)'CY,q,}2LAA}k/Mrtc$Y>u]Hb<&pH9l#=J.!M+p]3AG3@k{p1#x_ yY37KRB(?9]fV"wx[-&+bE(yMc#+tzmh
z6S#uO8,PuE^
>&%zOJhV|8=F):|]0bW*.VO,x'J^4xwJ2BX1o-^#q`[X*6	Pps$*4qlf3_I;ZQo@EvE'p1NQHH-LJq@tb#'+VQdE$2y(fev(:#)Mo<gjO"E7bK~o>5?zj0Q[?n{(=[83_98g3x#j>PoivtOz&pb[TlX1`}<v~9fUYNu|YY/=O:!p<$yP~E 0/.N3!/Y[K-n21[7`Qu"-4z:k-@y>W!Rz
R;=hN;Al3	RQ!!xFd!Fnn3?AI;2!
L2sk&p8:Un0$:} x58r{L>]dd3zjoO``NG|} @uhk->QEc+f|)^XyY/H9@s-m{ydIf#YnmbZ1h%z{V:A-No8#06I`*`&yW/WgQ7@&;
6HZBEb9y5JS=-evNFNIHZrz<e9"a[9Yf"
"7
2TCwY/BjC$r~l"5Fm?{*-U9Z!d+-*EmR_%3@S'E8F0W=;@tY3)7S?<w^Nc
5BmIc4OA=/z#9o}Y Pc)~e5<t^N1fX2ODH}?7E<}po5sUP\x'cUM"6DsqWpz~e\pr\pp(=+3%@
2b*:]k9n^k)?oX2{MdFWE&1.SqFoFhXFS~M,%vm,}1SY,?<W` 6'QOt)%nQf|}K
LuGoyGH^aQxC3R@T$dnxv15)ZHhET'2cHzYB/M`._bso{<jS:!6HA:k5P`q,3HKv-.N|2yRJ&w-?yT)&Da|r"+X)20wiN?NeZmp3;$619Lrc~wXqzHQw
{W$<'!Q)LC|/zpudGX15(RRQ_b&*	VQ>m8q:Rr!}G/hnhU(PYMX>.dPZDwxOE5VV"yTWNo+jw(D*8p#iRy9$J)-#H#0\g)f,:kZeVDMJ50knbW"nAA:yK'(\<(ipFTKuv1C1h8J-sV:^;S0iffS8W21\/J!~LRQ!<Sw,hjo,GfoxBb41!n^ed7'Vu8${IGvL}^n`Uvv28,iUjw*nxx!YqmqR=p,>-U)tezTOAF+NcNe"'KE-;qTw+..MEdTjk	\sEX"M`.Nu((k*t?YX<v!\1$5KRU&Hcog'f',T	*Q_,6uk`DTBY03Ir2/d^]KDConv_RiXVx45#YuiGtjw6nL$9j|k{p-RC<_Rd%`sz^]WaI/;f%x+d
Dv*_T0\^cvb}2`7//%\Tq4L(xt)j}di6$f*c0JWLCB?^g&no@Hlbm	\%hTH}<%8Wxm9$bc0
>\J	Fg-IV} <G[JA<)(h's[8S4xSTDl{6"p>+IUl||x)SyMq;|(e-bR=S0+tWbNjZzi;&:-PL'ZSi_QO0jz[_He=D[*l&xq(;OT'.i8"`]a=on>F.9-bl]E#Mc>:]k3]<0/1M,)Z_fVMlc:*'qo*rIpuoOccW"j!LcL0UHZo.B<1YIa~=wv!^<n"I<X}Xrbo<>V8IiHR9CnVT.{",B/znS~C'p:AM;vlQ`55[3Z|ESkyUwqnxMhOku5bb65gf5rF`h=d"[OTpJTW<(?8^EkN`P/IzSq~|
??Q
yp,OF/0!1bGf,hk8:ifM()H|3x:|Yg^I!S>8U:hzhMr=&xCZ{$(S}78hA2`MqRb2pBuLI}a^JsV5]SIb:F7LD^]%ju&G9_h{$;<[MX~Yj?3Thi]Xtzvusol-eo(	x2!Dg[I<kJyEuGh^JHc=|Y)Fn'p-#EhvJ:VrQ!xQ,&aYM%<GqLGJ	Td^rOZ)zN}	hQYN?fJji)G*P!RP0-HbH?+VIjj7^gTNM8DHQTEd=9J1
n9wjeE(gNrI}M:UUw>Wp[=\4l7N!p2bF?0YLq4QReQy{=iwIo1ULebxK9`Td_n'/QK5P*+yt9zykJID1j?w%/#5bI(28zMKT<5eGhDz@Q7	N1WIiyh2=Jhe2\3Er*.`FCUCv	"?4*rWKsQBi"YVbU1wh8It"^5?vfV,K0WwP,jGC6ELop^w)n:!iWysXA&"=a~,?Z4LbnAm(W5nLENxa9k^}B;.21>ym|kL4?*789.L07h
KI>+#\?IA) -G'n	$gU[xV&L"J|&\He$8#	F$mC&,`'=Xa'mM)F9+k6Ms=mrDPkGd(eA!`o_Ei5n:?sj=/#[Bxh~Hw#SKr5FL~ndzvH2I.HM*r[I	VaT+>9bIe*Y]p^D(d,U},)Y%gAJHw@`T/[x>}"!$Q*pS;rfqM2at]gO3TIJ#:3}l;*,/Qe|Z1-lJ#,/[rB'6Y3Hr_w^jFOYnx2
\@VfHEQ7T}+7nTM6-R`:b?0lDhGw(GBW*y<Cn0djd8U/|9^'.GU!5?q~+4CAB8Ac-)z>7)q\[k	;963q_JV,=.kfua4}U6La(0PIfnp:>3Y+=GPrYm_,Q^iguxwe<._([iZf5	2@Z *Y@KbT
+5+D4s}N99;\HkW8@zS+$
'w8kQ[<wEA`1zz^y	'_OErcjS"WY*3juCR1#k1Nkl|=zKh'A"%Ho/Mu[u9n	2"HY|bya/|a5E9a]0ur:w#uQ	?WFja.8ysCj$^~3yG(Zk38G_SzkPKlgq&X\dC)e	(.![yZ0f\Orq(8\_F#P2,q]Dd2pEfs-E0nPbjDmPq!HQMEJVw}{qG<L|0:e%-9blIoQ/WoyK0nA..ohvNM6CNkj"
$AluMGuL0ej]mY[n|OR1'-@a DvA)$sv[0|qTVLkJI\s%y8o]yl	tK2:)IF:?eV\KvGYVqZ'8BvvWp\2ingPBOVVk~,59U9;h4Lfw/L=	h	8N[\`rx%#WT_[r05dw2KR\)U+=$pKD'3^[T9'9r>:!sB&wdkr@mI_ 6ZM^r]_rHH	mq{O]^}b$CK86i'8A@:Yb~oz'94^o\\GrSg2	vJB+O<p;{z?E>o`q0'Th$7wh
|+V [xC(L&JqQa;*<SB%8DPhB8?zsz5mpCJa9g>Bv%qK1$HrD{9D#H	Uq5@SN|2F[-51fNFR)*R%&CIUIe(/)d~Vc%i)ot9[4*(y|}h
wpK?#u})/T"zCA\:>G9P@#=eR48-tIGGTZ?;:R%Y@-<,n_ #ox4C|eZr]-<zNGl0oekHyx>y-I0chpF$"v]J?7u+
EwtA;4`LqMF^yDu:xM7XaA~Fz&xS&b19Nm{ Pa'Jq,hBufRsA<.QW0E|IMQr$p"[NF~juVBJ/j1r.xDz%_ZDguFt=Ctl>.Vk<bjXQV1yo2Zr]fbJ^&+seKv*i2Z79)"od:?ck6|q_o?z7!B=l1T("$49PHQ9T`O%
Ra+|5~hv-1)FQ58(%"GZ3M@JAt]xSFc2GHI_X.(P>E#`B
Y<RRyz~_'z1)LM~.dC19R/[F)l)-M}3p3YAp$>LpJHIc8M
bV^HG:SLWZRm|<<%\.[2[\BK+8Jd#@ME["bC].KvHmSZS]2~|hfxS.sCe7WRoZ$u55o58^\IA-+ZXi>4=|/`7+V l f!`j[p-cu:b^F{uW~]J_z`G}3_Oh?	\X-*OpS61z_CIhu${8,x6E>gu4=<H'|zG`OU8r#xZeu;I>(9
CA#:3'P^3[bAKa!6RLoKb7olaT\D2zXI]7l~{A^iC/MPrzV{
fYy&KE~p-Pa8g*	MCn\K<uTVNf!d"Eg/",yn*iLVp`PN*`BjbGM\\&yAWFxF]M5}Yu>TpF3py#Z?<r@}$5>-n:F|i#}%5N_m'R,U%w9yagnl9LP3G%!l{:$i=S72fZo:I%$h.j3N<lk9;X&3uMy/[G_.F`s|`K3~D*Iexi4w4=Ag}7Yi=kKT>D<03e<#'lVSisJaWAkZW%m$me-/}@(T/)*V&kK|;(doQ"< j	=sHu BAjsn:e"0gaRkn9'42832Vqfq`YG6LE!{M#I"^jL6e_AVY*!1jt0<e8k(]FkTTHO~R=y_}5	>0=QbQzp)dX>q'>\pT?4GZ]=b)yxZ2LC=7Gw`=;T\`m5N*H1.Z&n`H46n{E)j)uqJP+E2BAm(f[|Vxco9(.FFG.Lo*iyd$9N+a&{{(scjY3gFLz:B9Lz{C%KTU]R;`	$]ci{rY	m8GIS#,Z"+THTnEKbX)(^0U1O{rw+:AUL.&qKJ.*=L;Ah-$Nr"DJliKBA)@R>JOC8 $E[kfEP,F^Qn^nNK"X+xVdA(3~WzN!D{rJ-pWM[=\L.drr>d=5a$HKg])ZrOp[ODgi`4cA1m!}fmO!q/8A)xx!n}5R4cPKxJvA]g\*22HumY8jydR+&sUi)XuIb+Z_+#bgfj_re?`|g<3)%<iU1$cUmeA	`>of\.wR3zb(K,b?v	"S12avm)(>=7r(iz"}"Ggq_l5Tg0)W6/+V/J]E;\J$`r&`mxs4_ETZZ)02)AMS7P"}yotv}kc4aRf]>'j1
ZHPqYE\WHsq_[#P,k(b4y;4GQAp,FtE4">zh5=\Rn+tR{hf,Q$%aJn73t$T`UfoIGd+bk5)IhIgQu<	F4Q3 :Fg\1h9Y@h}@CW_m,p(qcc&ooI
W&NEr9nT!^X*upG([bs#lHE[OMdHRM#oV<.\}6816
6yD<$_6VhipazGDj+w"VhfrY(9-4Bz#9m[/wQQp:?ZtG3C_.@|qkh@Xrz#c	0	8HI3;=AI_Ko@MR3W^nS{
QY9mx/w)0I+$b{1RFhkwO5TAv*g17Q$n'B1r3B+|H!A0f(n?U\6\g<`_|,#Z5lEB]o_>0DZ""?Gx,Xri (><ga`!UnC\Hx#f]%|05M<~R,B@P]GW;+F)?pfN\H_r	6=P9-lG
4,3|Nl'.J	h\rtC/G^1;ioJ6gu-XzFXv/]	Vn#7$h=Dl$(K2kUn#3"R"wH(DF-1Q^LB/4xm
 q~FW<MxMJBERHwtZ?jTE\_O\AXWf"b]&ira*~z0tm&4r.t6i@B=:X>!C.H`u^w@`L
lw^-WB
4iI
9;O aDV%}hSq{=N^<q.g/P}U>66B81"L(#*gfs-zcZ-s9I9:w>#y`V@/hiLW%.\['6{b?54F&ia	WaXHB`K0J.,Q"/.[9<N;N|zi5!==`)7g~F~R$}P~^/-Dg?s!`4,*'=U*c]RK5J[D~O0+ aN"tA)Ez}T\;!lM
O5s1g)`=_vDK=I=~_0*^*,?\,X?BMOj>{'Gd2L!aS#c}s07l{--
I#8[rGIcNjD;4,PVe0D}?+ht^k0#}#K3HrsxCbq'Z;Kp)t5eAk8Ut|#z|[1%|vn67*ke!U5"%|}y@bq3*3
'IA(i=g]&!Q_U4}wt,#Ctckq23R}pBOSm&X
S"'wg$~LwvW-q2"|=\!]^X@]U*my")hkX
VnlRyoW*4Mree2{1f&\8s4F.9hwTJ=nloeK+Y'S?n5"&}r\/{zN8#d[x\n$@&Ql/LiJc'31uU[p&Kxf>F4'KwjbLb8d[P	,w==hwLI-}	_]! Hk%AwCPmn-aP3kGl!D_ @Zn5mZxOH
7]c]AP*o
_a}]Hu:a$X{iU?8u4!\%NtR\7orfS=^4E5&)t2Jz"[A\4[yH!
ZA_;r`cXRF7.D%v,zo6E	>.&
8\;]&	HrKGI>40_7m6.d-U(J.Ny.BY~9C1BsmMv|9!ZjVZio'\&,q{o9.au6e3^A~MC+z}~c;~),I:)),ILTqp":.Hb\Iluz2W`_9N)IRagLlxyB3ui_R8iZ8{?.fkV+"pnYY!kwBx>B!tZxO5eb@u:.	<H]53>^e8}Z(Pu)W(;Xb.y=BJB3Z4j\@^M`K[40Ou$Lzs|Fr-0W7JM'~_q6H[-;Vw$$4:,b[xk<$UgImKq5yFm=GIr^~u
[:hkovn?-BaI(soj)*jZ|[Hm"
gFa^fL^)JInfaK\$lD~]j/*$|97?m./t<We4':;\
{&]	P{CSfr=.HgK>L
s$f.lUhNs!7P}-{<F'_ZOgFg@#pya#&f4cp3HtQ"D]UiFIY]N_(D7dfW@:r6GD_2_imll.pG@0P$<:3~D\F?S:"v=FLrhv`i'1q>:eJ1z1M0sV@y8KmR-]QTHqv8?W(
@!]OR,i6N4UT%yg(DXT6)SbP]j6wbz!.3F['hT\Lr
Bn3fr~l\3V97gRe4Xp66g4aUNO/E<)(%PE!24I`SZopX\z=Dp53K%''HGt\iz$piy1{X^[u.\|%0Z/<l,TZH
3*Eig19R+]0(\E`_2`XH"]2hvUc$x]31u2"zVM.cbuStRQyXrS)9C-\qq\w+TQ%;OgW0k@O@ON	@@[?{>Ln-h=:--C`uZrHN'Ztm5Fpq}y5Z&jr=fWi+6bCL{N56,hB);_;-=m5BX.
e<D`=!Zfw+Zk#DAj-/x~MO\T>kQ i3qc:f?t,1Hmek!g/;M>(IsyUOxI!)7T.K/lsK.kw{Vf66H<|#vE9g,\H4M~,e|(~KL:?9Y>A5!i?@8_k!|AIAUB]F&(LYMDS1\Ons9uvQ
:e1`"]ni\N8%~abK0'~ydqxw`"kkLJn`f5]XXHw'sXtj@aNtwd!;db^qQ(L+o._AuP+?)zTD99Zf44RxH+Oli.sYLww6~A;60pJ:(
=VkQj(v33KI96T<NteqA3Ta./vPpv@;*j[	wyT>^I m2As;f50&{0`(bEG=,"Ug1=]{GTMc*$2[yH2	<a:%.[wA	:Ndbqoo-MNeF}su]-.vkL2Qgr>j,5G?o|:2JsA
i=eTNU1<xgQ3XkPdUnAbhuW|C4\Qc5(zueaT>X+bg2KaQG0]rMtF|}2v}s*v.|D-AD[.`3,TT
 ol,="QO4>)u_YQvsZkS[&
v.W#PFfn7g,B j+O:L8	=R]~!`j+1eo^x!Vs-D[x3N45d/mW/xou^L:ce+OC!ceFjn$~AKUv.VH`up#Q,FD>
mHp{
n1QPC!!BxClB`y!zmpzRXm3S$q06]Wa9:p'`7%_6UH\gni-
k"cVE}TxTJ(;)jrT+&svh~(?Z~ U"5Kxc-="`AllA:_!0-9'uI'yuz9/.9GLsJ-{MFtij_g>}Vcl|P&%_k9K0j|iw{LG0%ZYpx2&A}%MX0T$,F <0~n@s<PG"	eMHv8Q9h(06X_D+3N^IZC[tk)4jEUmrLCZ|X-c.\k,^62Fla@_F#g |=)eM#b Ls42fVku+F$^z((@NLOM$
zB
%t(#7nr2ldtQK:Dot0c`4TB.}]O}QX9-l`J~[/q?.?fu+G:m&Yb\%J0ZV_tv|wrL&_v"5I@Py:Yq;uGe0gv%U'<	M"^4:e+jXyo98A0;ru!5A}e=t5}M78=J,^"8{3#3;#w43ilJv	Sy:+p(JVun^f!r,H}a6Y~EJ*>UvF)*R
"!KEp5h, 8exXA|Tu;X#_`"4x{M>zc78{,%Lwpt%/V8xQ<b5_!*%UCIPCr
uJnv'x?}aKOpRi(?U9Q:}>+D]G`#zrqf|0T7y	@qZLt9#;tsQ	`s-xEI#Z"sWKn&WoC\}37>~xpqUg,TzDs2X1x;\	~:|Z6/(ae,22/Wtd=$suWLk8yKL<$tK?ey7"84yylFO3-"h[W5%|<}!,7wMLZ<2aj#v-A2nOt%^vu(gTt+H%HPp~j@_X4wsUYqM)<,,4KPc`}aa\i":d&JZ+<%pUAjRC"mR~3I{8FwmCa}c5c!$vi$N%`zfT&\964L$En:>0sO:0@r68!z_*h+v6k	7q7Ws.F]sP^}2~13hP=VQ7s=cur"8siLK*E=n80p_20{Ij3MZ>)N&p3~IA[?(|d;m/6@(
'>WhE?zh9(?yCAwM{#!q2vd4AurN"Wc5#Vaev4JbK_IpTy"To;eEBO79{#FpR3AnD@mUV
c=a8qY^^U3[@vNr=q\Zr+Wzh]r0?~-:JCCq!^-cJ}+CKzlFn`y%F)$$}`wP)(G[9&G:!ygx3uL8F+$;d3DzdU&_?Gw4dpIk-sp[r%N(YwHrVP>znxmOt(PMC={e?K~*50g*3*`Dz\@m[AE&Y)n&RR"d?]0)Cjx-&c@e5XvW VFJR`,BSs*0hP57J;t;Q~rNKisP!|uL6^woHXg"R4nD;;
uM~{BRIOUd,[co.X
ON-=bJ`4\}aqfgkJee{.H<@)~$!8?dK$ohd\.{4"-kbH=jOj/wyU7-,`ABM:5aWLnXwpb(g8KF\!2U3@-?JP3zJ(}W^V"T_;F%X
kHQ%WlTF;a%TE.)2s6Xlv7o2c`lO-e$H!Aydo^zg|f|;Fa{FooWODgRo5QQwbg(.Vx)Rk^FGA<>q+'pP$v}\[)zQkTIoSCXyEh[1-G@qT:BB8`qm,<CUP!T@A=)/A#S30	[IKHL)VO`Fprvr#m/PP:c|)4|x[v;MH0A}; c/b%KGjRV|\'?'NBGb`+`_y6=8N~.;svR2	.R/7tNDl>W)l(@+c#y~FZJORMAio6<fZOk&bv{]\Hjzqhy;uwp3^`
T8<&}r|*GB;E$8`*f&>	_I$g#6wlJ3%S/[D8whxMO3xq-zTD5|`hvVnA~&-sVEefV"0sBNiKYjtih`a%S.aBj"(S	6NT-VDY:7dUtj3\2?+6OKPBm*&h.6AzS	ai!6^0X#\NW`_](&_{zRqiyguK2x+THrdd?1vSm*-hq7Q>jm:P^eu9b%@VV}M@YM=@ZKe)SH,lZYsL7GacfD/skZ@[%Bri?V`iI<8~gVAU\k0h^~R
Mv-Np, /hRBz/@_1s&+Je7)d5lSRY.'iIR6t^I sc`PN?Ok?7A[[]"Q\_MC.n@gXZy]M!]MkrFTSj<8=|J
~}P~m5E5a6Y$|@U8H7	h},'cb0z@ZjB`KJC<<:Pe	_{_p~D0a_s<v^y(?id]wpky uk^H%16T8qG0x&Yk	2PU=%Xl":GPOu]2xc<XD(wJ7;* a[_Z6}NZ]8WUVa/6>1HE1H7n5b_O4_Ta1M5EM5m
y<f=;a6+	=R+Q#df('kS{lh|b|KMYSa5oCcP`5Ik%CX0f0_pid*=.XmxG;hz!NAOt+Mk_($a`et
{If.^Zg84Q~]]HwN_osqqS{]p|aKx7f,!+cJ?S5u^Q-^c0ejHw#-mH xcD>*~[;U0>r&ihy7kiQ:o{%}O1h8Y#8HZe9m[]ylwWXeE[@FhI( 1fUi(m
I_57^p6KQ+?
bIJd:V!b6d]m2Q&$z$XyRQ]VD(~i7fA^96HYW.R~5[p^/]	
hgqrFz/p	\LDNF;Kl~@^-Z@^K'!zAkek,,$YW\Tikm}xAQ>@A=)TTQ?E?|Z^6pYww xY j:2ZeXCXW/><S_W:|xyhp>?E2K%D/m:@TpYB@Juy6^n+n&+'Z1:n J{RoYmn)1EUIG&BE,?OQdhre.o.mp''OGA.uCYIut|4QaxW<Ydjl0GX_E(u_fpl[TJtej%x)2aLdAG5ecM(oL^+)|
2M?-.Gg]iMq, FPE"/z~I|OtH}$"r0fVvI\z/zQ.ZL4um^{Ax$g7m1X6hw4C:&8w@;x5DcchN|H`:NQ:,|.%,zpNQ!m\c|Q;ndCm0uQ8H7zo|`c}hlpl@nv.3,=_Q]}BZY;<(S#T/lR\=68*\EO$Q\5"1>G}Nfde@Y
E;+JGvod.&^6|b|N4lQ)grf+v\Z#WcoLM\X+{.z0
b</^WG=F+3>cRG9#xEH;qb"c1x3\yu3S&={*kQ6|#y[kfIW}nz7]o_?.T/oG_8s%|Lg	Ek-tWr(yy>hXJ-}U\,:P5;b9QU2&2M1=x.&~E2	R'fRQj]SvNeo}':K]>-3|,_wGBC1^bWEbW98;]h@	'bPRwWa%W]=f$cf805vk(D[+-"]jmdWB]QS
&bqB4YO_G^WF[E|>Weurb1]hd0+>IV*q*"#h1RBA{VT#2a|6mtT`9gzeHZY%kl<+-$0x{*:4R:}UrS9wh!=orc6CR/<i@!0}Cm8,GMRFB5,!lzH]LB]\uu%N?'+[i/PvYWhhTua(=O/2@sC+UjF%#\}jA6	pEoe\x"]i$\[Zn1@@3>Mfo-s[WN\<XC!-o!\6d-Q}kNx<[Z'sG.p$~{JgY2sL1.#h%&&}CFS.+iLw(HF~fM@A}7x_davhWPHJhrq4s\nx/66[5]})_o]~/x"ar6dL$pW|5sBp	c6|^^]w&7JB{!/Fm4)2Zx):hR\sx`eaca"J])gz3E*Fd|6DrJ\S>(O1cLPwf1>mj-@Qw 71iRs%)uoc]u\*4Cesk=Zz?3T3=FdYG8MTAhr;7$} 	^~=mDL&tG8f]&c)p#LrM6afT`%n+R3V;q}iS/g:o73d0%dFs|pB7DfBF<Axi"xHzn1vQRF~nOI:R^[+a>mM^C8w.\m0qED!CLO>MLDkBRpsTv$AZ[Y	VsW,zh^l+:%-4rF~ExM"Q_TT/(ZOZ,3phM.G6m['vZN)^32^3*M\Vr%bZ8MNHrj*imI+SjUUn|%C9j!p={CJ`2\SY_m,Lx["
S,Fa)Z46ON'gm$q~4zxn{7uUyhE#<KFB5a>1./7".K}TSILP3fKnBv@/W0*AX6`g&vzE8,|AqAm;.\("p<f56~@"y#R0	fUYplftKnydXSkMn,L`Kh0y9]@_M^n0T9ZZa&<(S [Ip;4Y&3m>S]}:(K&we3O&m@|Ien2 QhT^u-=)qd-m<vG=3izhom*yv'*Uuo[r<W`'2iWQ(WzEzf5!uss6\U}/R&$buews?&	+pGl
lNW0cEtChQ%pIXa;b?2;fA0Jo_q?uqTh|$o}zpFX&8qkc[XN,`r[?^[VO5!||MhIJWvJzlUp-A2|8b6_dM-	6R"Ur[G#-@&o42}|-},	T;WJ~*O[!(LCC{YAof1	4/B"rz7_t%@n&+v_Hs4MIUw5(HQy$ZZ7G\mU]{DSWBm,o{z3}w*+bW @i-w6v$W
9Y1nf7RxZ+bPY[7 &TczE\2V-mV]vW}vo?,N[zJV<f>$I`~OGD:+`e_:b4`{uE5.YzDx3	hN9q^]{)W1~oySc[|}k.|yhE	I	H7~XxlsDJlzOcgj5?71(!i
v`4P=
jMH,5xgk<?jz&?jN\u(LcH={xOpK'VUoqP+qL-EEAOl=Fd;#!hkj3QXOefQS{#NxZNs?zfn!1e2'h/D8m1oPt5l!3_nVUI/Al&)46<8w/TP?0BL6Dgca5vk/i5q_c8WUtC)R4$?tE/Dt$#VGeP??+p[VF3:f)*HZ{
)t$kgRTWQYY2/':PvgKK[7.LFUd,{1[ka}2DgyzFkslZ!OM\rM)dA0I?JIom=#jJV:S`<d|su7@tpY.=:Rf3\_[\%GEJN:06Fe^9NSE.-uC):I$J_qGN\iSdwl)X9k6Ws%0EO2;s+O3	hq/|EexBV`Z3*7+4Dr$iT^3xRSnWh\);#GLa:_XYio$]MIA-!,=ld[tiW+u4/v`M6Z,dM;J;Bu>rNCs\@0PZF-Yx@D$Li:=I&nQ=>Fh[biGx4>+m/WnDO=M}`i2R]r$IeQyvXN`
SLi$.`#F`c<95DB`)e$Q:F[l
FAt56#+E<R	,=(6VLs~B1G.dk <')  :oN7nDP"<,y}'m}p20-'\>IM^X0:gMJq791nd,qS?+R/5TjxP-DtTit
aONP:0}yB\];H-M=[bTD`VP##In_fhf^w,y!q/O{L[]?-'
seLq+psD%a/kx!aOTz|;cE1Av$kzj4CnP5Dr;HYPM6/)3-$c+`G%%7\_t;[b.3{;u-[q:eS[LXsT[m&*TXU"~GzsCp#!-W(|{~Y6$
?)Pcsx.=(=Qx h T.HVl`&uE B//~|YsL:8c(9
#P:,y-?5%$L]LFb~sC4`%Ga:Mb|Fjcmb4<1!HOf[HQwT.Y$X, :'"qyXQn_!M",nb*\tR$GjBkU~^jIj4!bC~suZth?wLvS%v)Dk=(@	T"9?mnrQ5y@d`9O&f!hwe{rKiJ=6_%xIntRD+Ohgf0lgA	0QUa}Q{Oe]UiE`jq n8l_)kRQ*y}C5Toe_v'hxtu)7L%_'qbQ|?|[1o#=zW<	%zoE637sh?}z#_!<I(77*N<)K>(KIRIGH-Nh>bfp6wB>{?i"3-5JG-sY)8?kN5
VYvlMI)A c^^a$U.9'*1`-S;5jHA;Eo2qT5Q)Ck:<?-Iuu#jIds0{\4rb'.s(3kS&PjI#Yeb3D_s&o!#T|w*o2NmrS >9WnF@ *dYo(h"uk.J6KyZPejjD%91@iSqjdG}X2-lg.DL{[wwLbbh4vo%-ZE
)(X>P*Ggb!J]UuQcZSsi7nE+|A#vo}:jo}#i=TA*iJdg>h,ha:{,PD\yy-S"9s;.yp#T.rk<T&v%=>gMM<I*]eQ'k8jjwZcBld''6U{^oN9H#UA{<2&L=TP%uC~Q1no"H~t$/iap_][iws2!Fz1sfJ#mI1c)/'_UssH8*WCi~	|0e&JztT#R Ak#ypa*T8HK+F)Hju-:'EE%BYsJ'2Goo>atC#w~T5R"/X=l	d	_l?7S$zVix58l1X[UeZ?cw0?.OGUap-VgU\>+b2*%iJo_|"Mp"Io%ktUHF@W3j@vl/L~hlBiU!	xZ)bFB2Eb~u,FEV-#Vuo*jhrCnCuNp"x{E>DO$?gcwqdqHNv,Q<XYgJs|G W.GN0fOAz3:"aBfx9O}$q9:Hn okvK2S\zAl1K< 2\B<lb$#P	AsBZBpXQztkF+@V G=WG3.H8Z+@F-'A&&c!b.qMwhU?<h(OzOg78uS?W,!xjtw:e0ZrB`<
f<8
1-@tXH_j"$bP.U'eE)D9Mip#\4.n_YUFAMpIDcOklG7kS6,4]s/am'D2=Fq
n. W7cTz~efo1 Rs5~)5l=3M.(h0*fvh<8v!;mVCvqZ@*fs!f)*nP=T*I7x.7o}D5>)\^FPX!9+i(]sWK{Q<{CjWar5hG[Y'+ttxpv@|%.mAI.;p3QIA,4tH<l(d'yms0)2}%%Sb\ykH;6dG'$]FBy|rR/7G3u?db^=2Sa_u@/P
uVoySA^<ZBT{;RcV\@enUC<U*5HMWAMkM{j.1hR*&LsD FSv=cR8wY%ejri2^H`*]F~xE5YEe9}8(IOv}	{L>X{ppDkTu>P9L#SMN0dA]e=,SA#h1XVArC*C;6gb7qNsVMg2'=%>hO&|_AIW\A9a,"*sY'f=z2/s&Tz^#~pq1AiDp`t7ED	.GgWu
Kop+	My()!Bsh3?j^}\+ARC	l+TVeCS^>KqQ~[o7D4b/pN>?oopn^@LQ?W)=Utp;>EM8^^GtQ_VQb8{}9hdf*9GIs!Fx6y=7&>azO
uND}Z~Yv fxpr{,Z \0en&tSuN1xaFf_JH0N*@GQQZ).P]EEEAzz}'Ig_bElbcarP5iMn;zMO;>`Yb5'7q	BI*a=CG!-@>NV<Sz	wYru!R7J uD{je/~FLJ9b3+"<EZyX]+hDb~mDe209lF20Q}q2~N{bS$,)WLm'ji{!RA_cP	z;Sx-g;SthnOINFxq?tX^K+2-<Cu]mRz_~-ORq_in]y{u(<?DO_bL.,_@*gUn{{f>c0sc5BeRC:yN$Wxtdv`w*eoL_LUXwLeyc|VEpccP~\Y=C]A7<6r)#5_m:+lw>gsLb%fAWKKv]}?h%kh:@?Jt(qabF9f^prE].{H,o=&mp~a&$3wATEU^3.j!Z0FH7IBVo|2irw|{`I#~Q+AWZ
v7)U&^9+qZ=aa7h:VxM&r)"}O;}Ilo_y8^#Zp#OAoQ-r$H[BsqyDU?'9}oRT8'r:t>}%3/]9~9s"I\sB8`Z"#OjQ\<sp[a(U/::xY(GPvV`B-
pQ=mP
\J";6u0sJ;T}-rO|l% T5II*RhvM@8+T';a[|.$-yv$>pB<qNe7@fj|*+giy?rbT{0I;Je{!daD.Wj;lrjd*8MCxU97}d#VwB6jRkz(f#E&}6,n5j0*G{(74:DK?k2ZfD^Oe9-/UW	T[zr8sP:)Y`#&/CuZVM>}qsqaq=:IiFKP~p3
hnT:h(iKvsny>le}
4)o)/UZm/R|OvTN*;NsQoSNR"cgB*IQuLMEnf&_xgK-eCq'S3Lz'/VBX.vs/bkJ|YtH&^RN$xGGL9.1N~?H[rM/{eUit!4"{,h'l0bzx1^inuH(`U5@V,F(wo<[
8+x$hyff^\5{nOcZ%xMG)H#0	}6i4"[Cl&i2ef$8~-a$!qA2y;?\Pqj*${jd%3/s:BUQ!F836:a]`+
}yh8Gyh*7IR$"Dq}OE3qg~j!?[J+lck 	YUEy,N0VHRbl^?nwQECL"r3k`k"jNjeHEVE$O|_m<oU>gFuB!d@Gki&PdI]Q>$H:3I_s7##nuq4y!?EdFW)IkhO?SzH)>GEB?m[H*zthFSf0_5DDE|B8v@"#b1GEu39/ hIF?	Z[aSfDEhN59sNcQ'	B|+C1iY"]EXM.yLM>|="y[J1{`"|n.QlWX,~*KK6UN!ucCp,n<l-~BG_Vn:OQ&[-&Ihz<{@Hz'9R!%r|sg9U<c<N'Zln+4N#Y,P|T|Z-QO^!3b!{s::ks,w_q[]Ut2Hc9Py`Zr2I5<,x#Se\VV|YJwqI7!`<LGUITpj1X,AvI5s^T@+Sa<9z
=W`WuYvEt@%<y\i8n!A-;^Wb)yjc:cG.{Yqr6ZXz`qeH1Cva#q"OL]OwT+h]H#xT+6Wkt1'J)fp1^yNmHYAI/_KR)0}].\WAGjitOZ9BtusZz2,hKy@qyru>$tz	$TR{q^CeSt<y.)+Z*UFl?T)v5O-Z
I59\=Fj(rjGlxr#=ZNNd]%R8~r[J1pvH9MI4,SKh>2?},F%jdrzVuzyZ2kF/7J!v<-66gqzy+3KsL='$c?=&'aM6hoOYx235FCa*"xmEi,&5W09M*:~d' 	'1Z6]P-3	Vm@+!n=y=i=3g`".7#NP.}Xg$|L\H*	_1pM639a	`::>r+qB"eH~R[2pS+[	6#J"Nd$Y+}QSE,-U2/ak.Mk#M[JjKA:rTs;t`s5n#xSW\5c^nQNd.*Fz0k%aO&<RoeGy4S	
UCWn
.		Boc5
0Fm$us;IFrGkCTYl_+u	#{ekpI#$:1Ay\b@K0"<p(;9j5*M>@].L[(|T@jb7rSX:[hzU'?d;+a~h7KMGa`?Uqq[yL2X>NA=L7Uv\OEZ0EU2Gx}GY.w<?!;:<G46hsW Gi!x{kZ#+g/ax
jZy1mS<FFSJ0RL;\}QQ\M*`Jfz(7pXI3!i{d&J%WyN
4kD)vhjt*E?z	TlEvn8&oh?l)U@AHbzBC1F2;o1w#1_kJ&Tn:Rub	WGf_@Kw6?O/+ZjC}g# gv"9<bVtrB>(u>&=8fCX9N :+kJ:6H0K%.Ep	sgA_W+O]E`_G"!n!SivYo-)#{R'^&Ta0C+.O9,s)i6|(EL}'r*d>?[8{mFdp0HCM4pINI6t]{cOy8h(.drxG%K!YG'4NdW.=K`cpQ=J%!w;$/tic/6g+NWq*{?a_.n)ox]<j1
P}xG5w0#uIe<th1	"|[c+4KNR~U2hx}SU<~( c_/J4FV25bj+TI'>9q+7,F9::,	yAGL:N>A{	)w%m&z]kK471V!UuH5xFy\UeLiNR^Z4z'WVq2VdE~vh5<${;[?g@B?PMI9#'5/	gh~~Lg1l.lUSW4U|}[-ZM4/*-PS9_;VX~O\q^,A:djG7#LwAhZ'"'>J7/dSCd1uNM\|+!^maBb$7t
Oh)(Ha1@d>BXHq&?pu*`Gy_$VOUCm#u9ra7/5wq
udH<"t'3Bi=;[PJ)/+7x=Q[fzmpW0|83lRVEd{G:DS-}r]	I[d)}*O 4;VQ55EbFV Z(8zh)N.#sL>"!C	ep\@Euah({S3RwqL]4Wir>'BSDg}m`G#:%ieL"L~>3/Ym&@r::{:
>&vLwj+w<qvKYAUYsSN{V!S
Qq)L;N(5aMRKu[PiwuL,+
fTgr`*Wq8]2J|/RS3NC 6x/d)9?+R8Q\BN39$':Beq.VH, b3%"2h+hHU)7{(TtLn-j80
yCRs.m{-6_1uj$rw.H(M@F4L3wv\4Q}@wRLp+C"Q|~S?cXu#\[6%du0L@#p:|_f+Hg_*I2-5u'iU{U%'0"l.3s3&,+h!lx^V%eR;\D0K8">Bw6F 8~F-$Jcl_:,|fsa.kx84W+4]2&wZUVtaj*"rE}s	wo>."93_dbeqA^|lCW:N#EUL)5>~0]$
)pt2a(AQ5VrM~"vRdCd^)5YbysW\VR}7C0,p5]kY:8~hk^6tItLJ,{p0guO	Sh.<Dp36"o=o_JdT/kVh"kc:X@z,w6_=@!m[:,=j4_$[1SJz>VA`Z"@L5&3s	<Pza]_KJ=V&f(~Oo6(7~1W>!kg:==!&s"H"{&3UY t"xF=pfZZ3;9BesPG1{".IiD4BroA,oRAx)=(WG?kDJ+\4CY1fdY>kjF
PR!l=9@f<F`7\a7=|d,{nB)V	%$KW=Dp1h!;X_Nh5FpIk$7xwjO<5*[DAGg)X)SO-M8OCNV#s_~^E{orvC>wLB!<}=(vNTz	i,?gU]F/LaZwA1(D#-2euLn@hE*;Y(0c~`r)Wi&BT<
HSM'zX*CNZ,<K8l|ruW^zBPJL-YH4@_Z7{.\LS&Cb54skWN{A`Fd0}3TO=2*<ct,un^TNng}Z;+~mnu3L<(za
"QQ3r;!S1(KB/t5EJEwCCcG|y	V)	,~L+HX8y-wPSoJ:P2C?]y-- }{%s'(eu4r:P,-~BM>>P2]8uJay,"o9_+5zk@Chu{/i\xC{2_6YvE01$Msf<j;:|MPq-[@@#yKTd_1<AGP)LPDn?wOt+}^uHEV~mr?c(RFr}v-rwZyStL1Lm
BJ?V6NRrRn>4zUAvW|e0Pu$8#$![Rf[uFJ}+T|:Zp%1%Bt\Ii:X5=-Ly ],)aoWO.x!([B~P1pqJ(<'!ihSl7a_`1KRq	LS+`U=6@Eof&AOy,lurJ'Y%Vv?Q?(q%2A#Ru8j9c|2o/8D|1@ruHgeW({C.]Q?a!#n5zxpY<kQOoX5G'|)Qd_14	9YPQGK-_t:=NJQ9~qp^:ljigNb}I]22MjcmpeM;P7ueLOf| LW)_{:Y>=R>h%u|lZB="yCP<.(&dTsCBl0Hcm\AV~67iy)zJ%|RK-oP[4@7^(1}ZNwI#f<~$e
gHG8Z}wO]0Ky[LL&+>D]mcc;uN/a?@B*/SjId**#lg4wM~tOn,IvwcQP(,Fi&9M.\{k#"c=edF0(mM> Z)]tBZ0>Wg/b'w;svd^yi"(jPP`X]g]rsm]X%wT?#`.+	(.H"#UC.]Nn1a3V#h y)H^;_Q:BeHh+&(%Z5T6H3eP_;k)ws.|h]*mD2{l(0;A)zc@s4"|qxKEI	F*P2u .({iqvZmzTAF}2*r2lIzO`M_you1GGa$oC
4!dJGmeM'7lH6cMdn2~!}2IkKbP=p?*JZtFhS5-Kbt-@VVNGbnVzxZ^rJh	EDbggNG`x%rw4}sP$N&~6!j)'nDkB`Ne$ )nT
P^:IgM0,gmSK%4hdi+s	Q1ZUD)@7,nb}8safyp{!!+_	=F>|`CQB!QcMa/v=52|KvB:x6QKvH*	^T*iT.&(+O&X; |}+Zn(BB<3^"f`] ^<*rU6&#5:gG*I./8-;sBI~|li35#K5?O=	S{PAw1~jXCP*iE-?Jv|4UrWY rM*^//a|p.C{G{{!;uzmo9*M|5[1=~^iyN)-#_?k<SCrMJqQ9e-eD`&xdAwNn*&"oo}:wjwwvi!#`k~]wo>
t{]x,v!M-#(c6rs]npTL>%!v}asCFt|e,TcpbV	:z#'A}RuJk_N=E[Ij",^t6b]M`YEA|M7G.A P]/tmIloi_02pD>RO%.TT/"vQq6qAojZ3/HC]{4Zr;K^M'>rugh+f\^b'YR
)E2Jh2&iEno4B-g_*{$8'q%	>$y?"SUCQ2V(?xjpY#wvE?kxo6vBsg{k}-u9Y7f1E4da;9L-j,Po#$}f}nzrY*1:h~_Ci2a
%'0GkF]X	z4v7L-mwzcL|5=Wa{)Ez^NvKjS4I@qzNScuS{4l)j+2}8$T9;~IO%$t-Sl
ftpyw	WoA) 8$2'e$I0M;OtY~,Tx0^SvUQr(&gZl=E%%T1GFgDLf:d~;It|996Vds :q%>%Vk&=YqGnedK[d`8.jr(m7Y0 :bNUiC2v_/I9!U!Ecq+n6W=sUU =r8jP6BwL_K
kSTTi-eg i]>PjB"r6*E6OHTu(cl6JfKfx`z2=ZZ'A:^72l	3t-B]t4kT*O<,C@PLW,^1zPvR``|=TY6	W1;B1C%8;8.^Nx[1]S;/]F-L?poYu>q/y+ASe5CE^v:,6Ao?GJlA'4DD&f
mt
yugOBb4X-Q$9d8fx#y`s4UenR}(V-SF6L,^RjDW6ZGpH^*dy6f6:*J6IE}ySyPw{/zZ,kpSRSW_?-*_LsyA7h;XT|Vlrd_+'wb \P?IxcYgEt7%TDD ^u>}YN#R(Bf'cyZ=N$h& ZJ3l3'Vw+#>7)$TO%.9ZgeQn9#fw9^(b6QyQCZtfPy$2ulj{1-<aV(k6w:*z$@DmmJ*(b&fkbe"k<^uZwA~FDW*.@ZA)> fi&R&)Z7@0|L2]
i_=vAJZu8lWOHg2L,ONrRPJ)E5'ch)wg_CmU8Y	7o9@zi^?|(5I/FBecf[iPF}sL@NL*	uW>RfV5YsB}Y#T1O5-9LWsyxB+>fcTC_;NrTP=Se	nvSG8.[C0
=:icIDnP|e+?+R{(Td(T[x@#C rM|P!^g	g!h5-o\
HSz#OlaH(so$*!gnD?;h{lD2f+#m]
XayUak;AMe6Jps%;>qxOKOc_I*&l,RXUWQ!-+wJG`}L(}=pu*tKY<1zg"p$!KP`1bY.q[Srr
+A-*dcc>#8T8;Hz`w|J?Q'gMJ'H0MTcUh=JY	Hj](jciM9vLKaE8$pC?}H`/2dj&,:GG$q(;ygIY(w2=i$fb903hbQ6v,*spE<gB,Q">}uo:M?}HXN53J\%3:qh"P Pa8kmMYy}\UO(gFTZphuf3bGiw0t:*r/}PuuW))lqF"4;bCGQ8/H$`an$&<(jg1d}n?nCXM	MbGURygN9[8($*D8q-5o,kQ|7"^iF
6Dg,aEGBJGH"t5\NbBPx.gWc$ &[Vf@A0z.OgCFJ|+y"AOldO3g$Sh(s_Y7L_J,7BrVOAe;KqJQf__lr#42 6ye~'
dg, 7+SM=Pwz,![#T:#]M?}!.+%C#L}z4<\P7lP|k 9`!f[}6\n[sB7KFtmpeK^s@52;3L@R`UDDtx}Kr'>P
e*CVcYmoto0JbD5t,fFP/$K^WaI,HLU	'	R8H$M-bn8gtz8j1VUZ`$<9}+Xh>c=K}EZ%/#S_z~sg:y a6FzJolx?e/	9Lhj5mq:!&S'*&Qd(B??wzzxe`YI.Xq<RA[U7c`~tkcHM[6]D;CD`YKXu_\n[fTnSgoqyWG~'%]8^jIm8lUP4>K!hFzFY9#0U;KI{/*38v 7GUo/1i8p[Oa3xR#L~RX_buLM{\s e:xhLYVOu2T?(NfJ&<{JqHvEL{'!lh#7Gzfs@ &k+@V
`C%l"gW14S5aJzP&/4hFezc E%s?4=-s;G^kMd5Wgp=N{H^ACvd=T*WJ!z5
0Ig T(0_N@3G%"7Ct*&X!mJ?UQ2o{ 7?8S3fEC>E1dN{Cw[5@g{>`y"i&cqlk6;i&:m	c5df){IJ8	n7qz#ST{kk5+}5nRQbZ	94^2Nq[sm.<6RRs@c`G6:t&4ATLqUx2)7-IwGVT[K9-6G	5JE-/B[YW;yJdLUW2*_|6NZw!xch[ePnJ*;/!^xPT50=2N[`Pa@T8hoyLC*P#GEz>XO>3?zymbq.Oz[Qwd9Q78q@Q`'YCM;fV:W!W~09I?-2T56,~?bkx?Kc4.oIJT*\7$\?l~5P, /Q\9#?2X%+wpi_Vq^>=)dDLq2KH1-<by}qwA247)#^vO[1_q9x Td{=3krM?rgFr"!mLP5QhIg+rq:]p@,?.hXcX8>SZ9I-P	eo`;"n[B[h|a6<!wI:pKhCwy^N7{UxqElwZ`}CNFpH@
0z@1\54A38KpYA+[WN7`O!'B-x\"2m#V,hMi!ELK]S)+o5\u
s+$C/M>cPz6%b#I=u}<W_;#jt]!m;:)jb@x]!3*7ei8<D*S71C>5h'Y+RT;LK2HL,c]OErwsL,|@BHw|J4]{C*+?X(N!S6pW%-Odz>tx5#~fZ>=.g`jg>W>h!#wnT?w5Uag*;+M@Nro>
0MO7mQK\?W2n}=oN=af@{zu17DpxK;r/zC?+
;!\VBUwOBoYHySlq]G@3`):>/GXKU?7bfa7k@T)=t< %;*GtiGGC^6Kn6E#g(Nz5w48X/U4c}nMCil$`mEO=D0QbmIlg<iWxt#
CU]|k%z_v"?By7Im#=AE*z']C63)]$7h`4;F2?Q./K-Y]Xkf`4-;!{41]YO:-HNrf>F1d~P>lsWIdNH{xI[$,!2b^YW3`s+0qw[B'*Apj&`g#ktd#{>XES0|087EM=\0xg(wrVMC3_j"Tor43q}t=Xpl
2Z29#l"k%MB+?Eh80Ljg3hnYOCK;	%0D2!?4^6zBcJ4vY2K8e`O"JR8x'h7'IYl7ViEL-kjAK@i8'u)JC#}+0UPxXsUzks{4),t{o	&_s]RiH2o:zk(q;Cy8^[J(@2sd,|Ha,=kjAYesMzKk@n2_*LI)Io7j n2k C_Cj`KX&8IwU|K5Y]
$riIA!GS;DbIYBI*RiT7!
M`:++x (vR;E5Bac,k6<T}(C-Se'T]5.mww/PX9lGjF1l{q/B%'[[ry:Ke:gX*P=K`IOg@Barxr[ Lx}J9CT|v/O=kb7~d\t#36e2r.f_&e{cw:JKY6V{	Sm(n"xRSD5f%`0zkuv-"/Kh\b%`m1C5KLbjSKs#8pZ%o|BCx8tavkefEU`Uwh8"}~C,zu),c$T JMO	1o2$L\x^/0I6dh|wM*q	S;	qgeTa@klwO{3\$n\L7[eszoWZ{nIT`q'"
]:2[
.IVz%f#OP?"\0*}w4:b9Mp7x8]p><XilW~r"0Wm*oH6/?	&? >x8jj^RVTgJ%(|"iLS*Qo,zQ]OM-k+WT60L9T"wOiz"1g{."C L>4&%,^Ehmsf&hF0YB8>8))E]X	W<i]5mR=~{rv{*-a>FIEop7:^iN44ucgrW[8Sd~1uB<+Nm=P@"!6EhM0C3T3[pM~1P9; qw
5:cOKF_FqoJc2)13	E$)39ahX6y\h">nCh&c7+qS'.(dw(8T?tk|`l~,M.PaoEJ;}@RpuH&NFkR!R}gs?aUenw[,/6vt'lzY5qkc$a23%e8~7H)eyHyMxSKgdf(Tv6QBRe73{Hvxxs]Om-%pJVapcO^GG6v):8ewDCJV%mQMtL)3lSL:%)W9rV{HJZ:f.beez=&~bIQkF(;Qo:,jPU+cj+|$}3iH
Dql}1aLVwJ"<|y7Ue@N[;R-/RLsm16Wc+sk^8grm76RZ73$gP6s14xt}d"eT\l;DUrY.Y>M/sbL9/6.M(y4% uo]n2^z>OE#kkeG&e*#rh-]0xd|t%^&LQ]B*-t^mog->[EG^qHM7oK|YwGN76mtXW,
?f0V<~),gUtg:h)5LE^'5"}$<3z@'Q_1`sC40:'gvOb=!'B_OR{1X4Y-PwTTA(aw""vsrJ$+`)@!"eW5}Ij)Nb-O_!b^8eAsuW^#oR[]Lf"M:k6eC#7p$wTbV{O N!yz'xK;[)$@6;`Gl0}&n@tY##m Lan{4T!y_hBUWJUaNB)^n7y9@*yLYA\?=:SUX$G_rsvbIU/_N`=GV=x>~%@h4YMMt]O"_Aj	ttb+XN2`;c+I>6>y5B&"A5I#[J/fs,rww[~Q8+0VJWyX}Vc /4YU0]]v{NkLX^CavKD};/Vy	%20@4#wvD^0I~Q^v_*ncl5N&Bb9#!v7,|GtU8&HS+|a&!l9[Fgl"x+;cTYux7$#lA+MQ:`kJQP3?@<+_dHPHnYqC*\'x
2TQoR;JArB$5A":k	R=ib:	67NrLlm4I`]I<@^IvKEQ>Xm)n'4Ikc9`nm&y@"E?A6:s:55\|.Y[Y
9iDhP
?<n3AN}-3#cFapJ&[lhYzzh7*&6^std>zEUC1 ~;dE] |&d>uW4Pj?Jk->Vm\J'w2PyurG>|(8rxRK-l&YPi-wJN7gS[#>A`Ute]YJ?lv
zFaUjs6'#)	px@
8c8|y@YsU/:EzXJ!j6"1\Kd.!Ea%yg%r`.UW.D-)FEIJ^D@s`e6aMq*QV1+Kji)vc=.`gUz%1~bX3{wmM5'CE:'_*yo\A9%\xl}iQ;	*#<+0_2-<K0Go6~9FL+hxLJm!r)/TF?w%5(m.
JHz5g#_I5matN1gm]! fGw}4zTZ(3A0!RVX5r[~aCBxdMjg}!a;Tt8o(,9Cu2#`e,_=y}	MGY-gTd+KDyK\e
l4Z:j9')'/ADt2CK*qd,TPD^j[b^?c;N{UwJF+cN8q\O.ovFe6+[):
y;l//~V-6.}d:.eC3]jc*qA@5~#06L'0E@iRqS55G]G`P^bTVC=p39H%ekl`)LbHG'zop~LT@m{[ G'vf)#s{=UQ3&tU^s0:d:W`@0"Y)2?X#-Gw'w_"(A9E|!!|9nv1yE;4E.4ADl$oARP)VsPf3=wgP[y|$^;%0TTk3eYdhR TSJiO0QDOa<S"zmlo=7U-\r|/9zRz]Uv?gwCaZ1>c;aMxmb?\Y)2^):TP5>yUy(X<)Kv\RB^eDEc-2p5^87U?^]GjBSEBsn|/$A*g;TnG!'<vY|$,1R[Fb7wT/,yyZ5lL!)Me<6b N*_U-W\x"Y]I>(+HZ|{`zH[EOy!a!ntj\@/BD2N,z~-c"Fx5T=n,hFXG?_'er!<HW hWA5&EEo;oD](=]K$kvel"/W3j@HO?"<t##=.F#cjQ'Hb)iU[!o+8{NWfUG
iq3Rmj{2+#U;r5*1|It*Y(ZD9<d#S7O`|s5gbU.HdAO?imxPufY0jMr0<Np6+z"EPS:GXKp>hz%3NKf`K~KPk~TsA*q<PavCHaP(C|$/KF6@Iy"^CtZk 0-)eVR/B[t6P7]V9/W]]-rjnw4,BDF4#Rj;Jk2t7`%0L<`
|E}QvrA.lyMx$@i^jjaX|y@6\D3zL5@-Vg WM`TR-|lA=SM7n'y>=*Pd5$dmF t]
A&2"/$?wv;P5ym
hUasL_ !Zz/DPX8BCFIu<3n2mR/&U:S'vDM*Fv}^64|J|>WD*O#1w\@v.4}jcC22ZtU`|W_[(S4k>E-Z+	5dGNSr)wCP$Mk`5 <I#w*TE;KAl$K]S[hWA	]IG~2@jaXp`l0d4Op|lOw%l$Dt^GJ-epq5Mx)0+R^zd6$H;&\U'8~uvIw&x4/FkSu*F5^3*?c[Zf>wSKe#bffE{I*WQOt#T`XQ:x5A&BC.}]hu;iyUZFCo]MtVW=oD|G+ uK. rp@jnSp^a@\-Yg
roy6	u-F%6XOc@9XZQn)wQ`fQu_&p-KG)I'[v!7YAFIR7#S,7;(AK/:M46b)YeW@9V}N"9:3}w^8MTM|
MVl]4`Ki);Dl<z\N>1[f9-Fu8iJ$	y9X(nzMB3@TP%N?<`(%Ih(S
W+\zA-`Fv)mmyN{[h>0(yhhON	_&sK_gh?La YL[md`
)*N%f{'SG|{(HmsR
.xPHXci+:XeNSCo}b
r6tZj#F>7N^A&fS_wudI9oD7[9{&i{U'gQF $[O/a&,`u&%LL;w;y_nQvUykZJa**"sFr_pa@CQ[%u/_f}_`m:eKYco"8, :RKC~>P;N4d]Z,q$O4O]VrdkGWx3,0Z=Z}Fj{+E`&=}Uwvl,ANhMRYP1ATvt^bOqzyB*\)_;~KbD`L	L951p\Sohhw6Q<O|xqwmH
Ms)JEa@|\	eH^0QwYggvTkgd1=R`7==/?/:4,m$muC]	IKF4bj/KJd?(o6oE`XNs+UJ@x2YtP\	HrZxvq/qovxgH=lyDcS'|38e[{N}ac1#R+nNM_}dh:#|v0Xqta+V"yZ>ce+,Xq?R83ndmZCP4wE=CS'7kIs4#9~=Y4-yPkP>tWZu}zGG![$QatZ#Ze{7G2%D#urY07/p9::V#.4m6bE(LH$|D o`;XqgI#uuTll)(n`$_{!L,"ma!};Ze7Oq$sYoK^	9cPm_^s:1j]6;~=aYP/eTa`9IXue[n[Q^5-J=;^jePx&A<OX58vD=$!YK;/AW1vY0y=*e{N6@5~cLHc)DU_A%;"n9'DfP{9`D7~yDvG!/!H|94z6yY59dW6qD&';6Je,Cpassaw*V&^^/T!eJN}Wcx;r(~
,w/5nd`XggZpWp$_aEN2g<tL{K!Lle	IXdviNI@GkYkHcJKi|t<Cg}YuS~(+K|szOqt#]K@jb!>9BjO0
RS2`sD=5e/jCJzr|lO:G-/&9opCC{Sr:"7vJD;"ubHL$.=V(_Cr$/7%cgkXgwQhH,r#}nhiDrhs\ia3ED-NvUS/A#BxAk]YP81%Tf
IIm6G*tb>u#~u~mP>&X,;wB4<=WXqJ)u`zLb,Nk%u4^D&#I4Iv[r$Ohn(N]o!Qc5oFrCp[G@\wlRI(Se	G:Io%z0tYz(|_X^6'Yr7Hx()o$=KRb.dpY=!I"0t>+)JMe#Q\m 	[6vQOt:O5RO:'
x7[k;I@GaY<OZm.=CT+A1jRO[G6!nk?O"^$7]7'6Hd.2XM4\lb@GS!\,nf.EfNh^.8B|56ywm4z	jR &6Jso5BIvHcXr/sa-h)hvPYD1e/[3Gyeta9= w]zh+q'}b9F@;
fpZM8Zry<:_"iRu?yd[}dAKm]7(:J%+ y3RLC]Z13>SMK$|-g`:<mg@P
id<,=5v"	kI%<99x"+]	i'	|W3r5Ra@Idb Hn]kPa7GnYoCU_{(\?J1^)FzwZL/~0o&'5MCJ vBkKg'm%Av,z}}!e87&e)3mc3fTu$H3n}@GMVi"y!.P75]oY_*cQ%gRN9^F.]|(VYX:(cgP$x6UyA40>C%2 (&:\hlAp4S_Ziee4wX5=.*Iknnni5"ICWBm5}36>?l`EfDEY$yT`PIV4=GaeKjUEpxl8^)V7I=`%v$(\kS;pYkA6p<4{r[T.S+sy94xA=/jr{5MWN$2U*F3B7sj45>>&khd"9	o-[<7x,l@J]!Y00}B?4RV*'[5ud\Fh+Sstrf4XtfgBIOL=Kiki6l:#]V,gE*1`bb-28qL]`:0sYJ"p]J,F8[S0mBx*R2;T	yWa"!S@P1Q{(9	y~uCO|l3?_jH<ISfZ*	 :]EWu-,;<8-`n4irKPeoL!>@LaL>n)lL)?"m}) #(5R>uW|XI)jEI\Tj&@ 
VLfA!)Xc3nV+Bo}9jX!=%=z[>Dv0rpP	O!^1<b_"N_'WT\DDQ?o$9 juLwv/Ck\l{StT@
?l,O,Ym;We%,zXXx|
[h$D:p-(ZO~XVeIe=TVBV>FxKMS]uUQ6a,PPrY9;'!MnTkd-SocTHRXlXd+Nhv%leVEUbb4I^dw.yV*yz#^QuCYyt;rx"!"iw?5'Dqp^1fq,~nt!7VKa`b[w2i'	)-&~e	9_-|V)mS#kF.DOkx1+:R.yB5[)DFl^$E.O0_jPI6@AHRw(ZoEdaOWV=H):(0c&_@"W[
"AFljK{YI9[npKKy<5%DVh1?p.3k.y:)jQ;|<<slWk:Ug%_ao];7]cauQ,>>K<kI{k"l4~y@-vK~[st>aU;Z0EV=_Y	QDRkMG/1|>$UhJ/-/icsjc(cirYI0SGn%Y~>JKaffN osI_K_im;PY|.E=4{2ZZ*{DxH0=k6RV3mCH_3>D-p2akHWk,/c?j7gQroo)^Wi)i=wa	[:bB;g:;1W,RewFGfn=zy"]gmf3gBlOZ`'N$EY=BLp;j-.UfOdOe	LBa}pn"k`Ty}/pw=02p/,WfrQru{K|-^MO7]a-d")F#WO:L
f|nGVL
}3_{{1CTq[m8"+\.1c=Fx]'ZVp	F*u3SbwlxHoRIJ;Rh-n%Nj Qp4*S\X8heI_vsj>B=%ej;x?,:t"EMb+U`f*kmpq^i$vgM^[dbpQy<q*v
\>FR<9eQnCnNw+)~S.i	7(lXZRZhrFl2!c8pq,9P&ioYw1"J{{\cC/
hWhupC)/Xc.|5Uen@o/xMe=?,iwmH]F8vo|qS";n"m'k2OW*X2d5R~{86H0%vQC0GJn;tZi88Lry_x2X{L[,RB{G\5dKIDK)NbH{XlIi</dieY"@Yx%?nhq.WD^Qk>}mlXBv^w
`8V_yG4F.m7,jbLU?8t$Sp]R!N0Yu%f]w[$P\:cWdhTGK_6O~Y8n3V`Kh6MkN
m2R;<B|tK3e|_--g-_OG,k0F[u	'6qt4ZKc~ptGHc,5BALbscTsuX=}DN2>SqQH=&zAmEZI02/x1~->d=2>#:,%Q}Ie)K5F5s-/Fd+J(I`!	=:I|"kQ7%8e$b5
8!%pli&xSu>Mz?]qrMdi|=DTofK[[iLQ#yo
xr`I/K`o])J+,T^4mWY@W@`gijv'^	oc7"i{6P=I&e[l/!MThZ"1Y}.~V73|1sg!RxV&lT(-"C|:(*K,n0Z:<#*w;>YzNE_
h&rl@ef4c|[BGr|!WJiV1'\z#W"P<\Zd]F/>uL7.z:n^ot&RwTWXATRnJp_`W82,qiyI87G!A[[~[6+L/C4])~{2$0"pWi
HR022WAY2M[RR2$%u,L0!#.]l$Q{68b0n;X^1dZM{fQ$><||De/D'qo8_6!8&1$(xSn=D3PCcryDG*nzOI>mP:>xdXXf.z"J-)@@Y1%)R#e{'R%4*o6OT(~6`g5R\XM=S"3/F6cmLq]l:QbVy,7OPSD&A{n>wmSUy.FH^X
=2)y40FT;cf|`A+kDL&oO*%
0+S\
^X%d0wAwJF?).>lX\_:q&!f]hi^NUZ\+mUjyJQX[mZUEUT"i}\{!bqN?ND_AZ:1E:U#v}y>Ky5$mt_qtDS~I5
DjE3o@LFlkBR@f	GcERvT\S(%&DgU6aVG9mi<K`)m
3(}f+AtQJqIIB$#%QS"
FU$"	yi#h;f3l*Of4zQu% Ty-JchqNv51Pj}%G@5%N;Cj#W<mKOJQuA*\IMqx?],~2 ul"dk8fFz*Ao}yVq\yj?fv.lElk{+nAyF7Zx'LX='
RgxnUYep&lZUf"zVdW	2zpcw|DW@{P~rF#3]?4~[7|^KAV'f3I+;b^&4]DxX>wp)L`G>L _F:1|yQMe
p1=AjWh<Kf#NS1=.9e>P&/:;KM9G3-7H`5MkB`hqjB!kadmY:n5k[Fa+B1B!^fBgi>GIbd=[/%m	J>Nx2_,
bR4?X,2DhIMI~yrb;~]L0keav	n`g*Jwdru'(#Fp%ih>p.?/~sq>UnqbsDr4.>T&V7ZpEx|I{]W]D,<?kJc 1vW(kQ\C&sR3K{K[$8p6E]~E73&uKvv#*8<PFJ-E4g[c8
P0Zrtn\G|5pF6VPZ|;%*}b#f&n{g/!C;"cV
!hS1P`N9`iH]8(2/k>):	8hOjN^.)NGkn
sv[qm\K`[d(tjjA-(aEL]24x$5)nmzB	B=%-;gHvrN|tN
>4X.rbs	;hN1}]!C{Yur;TJ|=#W>0%FU.L^p:alN/u#{vpBo eyK-?Pfg_Vo%e]9[uGcbJ1{:yO/#Q ^NtZ!';Xbq5lEwJJ3v\++AGRn\4)uuM._"0=$w]S3jazY1jicf67I >G$x$?+@7b8tCaabk6;g<HFqrMdHLZR;Bx${+L1y6OE eF&/*$wqw5[J18)E_v;G4p%S.QkI"Vh/^M8%tj{m 8PM+y(AGr|6e">",R?_t8N3	dZLXrwyv$td*r$%G1K9L7re	jp^$(CuFoM-1[^Q?J\GDEClU[O~u#8oST<cO:B`I#}UQ,viDq2'IViU!l66krZ;gG8r2|C/=_/uu2vNc nhn*;']/(.b]^6`3aC
P-/)\:]nO:q|2>Sc>obdl<+Az8$g%}SP9#mh)kn~:@;o6	'b~Q5zA{5r]:$54}FTI3{>g",v(mW9oxw7
u*?XXvY+!EVCAe.I;(u7O{)m;jwB<eX@B*tc|ZtWzS #$6<I(h=O9_us-JX)4tCGsGDwB&^.4
TwHQ U^jW{_v<
	4Lrv--Rt/7v}R8;6Vc.t<3dXOBbfozh<Xp;%$l5	jgsp,YU"$Rdk
V.<A%&=tKCvTWud8E73Ew}nGF#4pj;*Y=@`Xn\9%{rowZp_<b%-vcrrY:F+G\#@l/6LuXaS^lRCCh@/\nOH9"~Eymh&3CbMLi1oam'm('lGoPy`?m>a/,?S\Oj&,dq0wKNW=@9JRl-Ex5zgJYgP+l^*ks!'V]4DrQ.#R][=x? /M(l/Wrwsw/N`OvXJ\_Lg!7!>S<jn@}@u~.,:j1`yw<WV<j"JpOAA?GvShx0]_Fx!x<iF6@1!^<ck):a*#BF]p7IQ/:q Q.t+!sKaz[;9pP<(ZtG|u`jpixoS@<soM5kGK4ki)nQ`nia(O''w!vu_(
Bw+EhUF$ja.xb9AZ<j5g->].FOqy}GXfryI4K>Wz6<jIPiJ&EeCtXh+@Ab_eHG)&>/Y^5QjP!Sw<sF#hv+/NKlqFo7?gK-q)n~Ik "ACO3sQl&r]t>_X
\VK;IT|@5I8Vb@l2v4Dw.`Jd)S#\pN$p<%l)8ls|xOWty[|CS$U1-_#/&W	bJ#O^SD*dTjV<z!B5r8G{a[
b?:d3+vY%^:*JGN4LSKQw	"1YYUi0O3q]%//7.v)ZH(l_><`6pbb_zP10eu\u=MBme	Es7NzSrQSY9SVe	nn56CP{ |6Ex&%&k[D[E>(N)
)oBwtVD7Fz?
$[LJr'l{;c=~/h`/ieis["_Q2DjbYDRi{U--btHif$0'&2=>NAGN.{>gGmj8%;'$-=2-x;LT4OKH
ly-cX	l>2y8$C.i$'
n@]'a{xbL29KAf}n5&%oicj"<j&3(I hBQMqFqB=IC
b`Hsy3?iYv_K?MokiCW8Wr#$v>"O$]{&L('Xmt#E]2~
!iUIYcmDA!zE.#>qYv03)l"i`:-h/eKu*P|
J$l\k&kebQnPH;Il/^Bt7{n)6_JdzI
TQxc:`[}|Gh2`os%dfrFUe76#BX<CTi+
K-(%(waD[#X+NKLoCm-E"!k-}E8Rk9t&m1M7lFq=
B.ckg$j<p$Y3R`j+x>5I$0<0`Ap,?!MNYv<0I_"+!\|madYFi<%<1!#;E`O,+fYQz[dfPPK0"sF^#bM EV]/ebkyAksT3i@Tf{`?FD#<5:%%bB_NDfI&-,O9(,0nN&(m$fn8JcM7/*Dq1#!P_H/N1wqZQ 9h%fAJ>]U]]4`k5yF-B)~?$ds!3BhP"1i[M@1&g&E!QR1){ +8{j#2ulQvbm8s;^>)8pNWePwy	R?GIS`Vz\ei(sA]7l=Hb)pk+ZyN8+d$!|&\8	Lj^eUdPS"pjBekf&6JVID.+ZZ|yU\3_c4H3Vi#i2(j[W!q+#1CdAsgM/@jl%tT7c>BhN?d}[=Nf:4R$2/pZ%xbpARg87u$@)u~C?[6[r1*VC4[m/shnLO_K5H;0[jgfrw_|@Blxo&<wjB<5qJ' xZ[mzQptI;gVALH#bVa\$lYeQit
k:#`s"`}.(lvK4lPJ'1O\8|
aw(MgwaCS-M,;&R^C+btD(raJ!=hR	UG/#Ip;([%=&s#4XMTvWiU
V0YT\3,3ej8fpLF`wR\tA@"Xk8kbCw'A[
M(*?:|C@Pj/s3#CA;87X%`Fmr8w-JU[8k@Za/	;}g'%@]D)9"5wqFIQy\J3x8Ow2>cGz>~p)zrc\Gu:y*@z&B!ac2NL&^1_TT	/N$'Do6Bo! 1V*Woq-a+)cwb]|CHt%Tu(98CW^^RS+[& "?i^!"-(\5%{T^+OT[.,'a|rz%
"n3<PP]),*+9XNxGw~k!liLggVo_5>`1Fz>f"cb<X[ZNV%k9O]^Xi<dNV/n]\Hc$H/A/Q~"0=8+fiuLx_)zqq4;$>:=ywt"quYn*CW*]URyO0K%Q^"t7ZH_q3vIbFtkk!jKtIu8FJaauwE2a)&VxN_S{/nMV:BXn0LUhm@9eM$r
4UT+q6Bi".@,5K\I3H!^@c|1PP^ct2>zyw{I~Q`$y6:(Gd3{H2J2?+i>B.(<L	\LFq#0YS@6h76)Tqv,UDb MixOev?rWn})Tj;TNUx+#00\A]3>qMvY{A4fl7zOy9>U,[Ny:l>HvhSb
pG	o7][pYtZ8}m$sA'^'_gh n:9\6L+a)T{KDbV_!K?hnydM+]Y%-Ve(Was!cxS2`"pEU.>S!@.|mV10aR:dcM(4OhXze9W?Zb+Oq)_ja~HVd5`+8t2k\EQTOT#m[U+DuU6U
 n.N)>7@1TAS3?:`/9]\]x<?BYVP0-$T>09;k/bZ=vAfEZ0Li"}%-qw2@F\dNO-}`(HyT,z@f	]L]t?R{U)3A	GZ$/5AY0|A!LFzbd[Ect+|(On_s,2"g5L22Fg"+~Y\=@1f{ey;07~ic4Y!GuJ:jRXs_D/#zm/Z.Nci|rr$378m32S
XD{Ra'#-4a>js":K1F3r/$NlED/A]?3xa?)IzUS-|x(U;0`NL3Zin2<q::yHZXKVf>d?|<nh1	{9~.DTWo@s]}mYT+C]o>S/WU`;2=`xMyNdfiM%ssS2,QsHm_"c/+w)G 7U\^	qj)hSnza?t#QQoO?'$uFOM/.G|dn6fgMjoO88c0@EepVT3fjoi(} %6`ny*R0sH&w!Ioi/N=}Am~m75guIr-[,'5_!f}f/x:E{=pUkD@T]%Ma!O(5uK	kS
m7W|Dgp/Tsn.FwewOmb|sw!%e>MrsdfR+SxUZh :nNRP^;G!q#T?3JQlY=^DMi6G-Av?NaHgJ_/f,{UWLh~gAt*o73J/u]H:_pn%T{@dnF7m
9YO&EY\AV^2%!O;)19@_?W#+6xGq6V>a.O2!s@.MzPSyZG+&q6"18rK/ @Y*'*"+{'~y>vH")cfv[2UxX;GFe,-qZ37JRY<46gQ9;2E,N8HG16u0)f*qytXBW_ =p(x<i``k3g!>S)#@kxU>AvY,Nvn=D:o{v5KbLzQ/INTf"9B|Yk%K\h"?QhQ;bHa&-+' ^u8<5js|	(77GwnQK7jRRZ;&%Uh2oS|8A(FexF8G!`'.VmkQy+@I%dA7LO)u5kzcsR|AKqk}%60l.!$~e4J358e#
?=UL81(6IIma
_Q!X:<91XQ^XueyA]>dpD&xE%K
,VLsI+DMz%/|8jUc1,!G; J>NA>	#0Lsh$Wx^U$&yrvDZk6X#MPdj+#*9Pwix,

I'#JzVM@91Vc60te}>|TSyBa,
6R_vAcAujA:T`MiJg	yg;39J?sG[U;M0%=kTJ/OYX!lT{G#N9*]}	1}sRKH:41e *xa2$oxg/!7}'z -UQT^\khyNub~;*Is4A@3+f=6SBG;x[kC>ELZ,CzYM}DN2Q 3"baz(92J$2y
2xCeCzg	Z?BbfFbk4UiNZIHw&a.hO(9x\HNZ'9Xh=3] tJp~%-{%ab[Z>	wFq1$PvteJY&5|5|Oj\z?wPEk< MknYvbK};yr60"p)hpu]\z	-vwH2]H#e=hRTUFKgVVbF@Gm^<dYj7ZubRq+sW#-EaTLq^(ve2	g#e3yX '5>kHdH:X	Au^\$EE]Frw-kpd08&!+`Vv#ZA@SEzss'4C`|Mf KQ^gR/KE~{_TKKslmu]&1	^p@5v2r5&\fe[]=k9hJ%y~hu~ecC(>91c)	B9Y?!k[7q)c;w3Wp-'AZN">MRml;\cvsp6f-ad+43njSiz!2vWv4wtK,W|ms*;Hm{&%#&e4P6z@b2U%G=tNL"BP+/]&VpTf1k8p{OG8zlB^1HMH/k}*jb=+%[kTG6 %/!{*y}Q%#G)vVtd*DX!1!:UOj!4@x6%yF}^|#3	Jl[L[cc8{U/zHMmZQmIWr[,`tR\lbw 'jtr'UKv6t|Qu^#CC'}:.!5"u'tN6x\S3Zqk]>A"dlv37@JM+]u?&ns
1y_Ey-s,4UYzYTvg'&=[rf'i<bNPI7@:9go^$[m10[Fl 1seqfJw933-%39#-II;-RZ7AM/Zd
y07Pia4+{8[| 8f%TWs%Hzz#WzLukIx46qGpTA("v_TL5zEr(y2L,Jo\Ono/2:XiyPlb8E>~}s
!2M0s@oD=C[Ek%raLL]{@'Y)`[}T&1?('-
r!"^{6_x!f?BNm*u_X_oq	]G32w\X^-E2>:#E#TFAn|}<CI*ia%I^/zu)1.p)lvDECGqs{r>H:%Q+h~/_|IK}
2Qax_.GOjy(PHD.QB-~2/)$JT~[J%G>)e+/w/iTe1vG<$jR5u'^cnmT
eECE|:N"s_tv;3`&$z dL&$3X[~y
^*Qa{G};SM4!!UdT#9kOe8f9jT)Uq_6y\\<0LF${&Y/Qyq.F=6X]]}pLM)wtgHu ",e5hq%t3B9v7P?joLu_}L-M%ZtzW+rXO?nOC"vc;(Qh`+g^zInMJLX0U>CKq9&?$8frCg{@SH<;\*$UTaCvR]4[U>@6l*cW*:-i&DZl`.=]	dz[_~8zaBr}I4e	s/!dFZX.WL3etSBZfDb*f!Dfx=+?<K-KWw4mhpM8NPm+/=/&gAow$W6$LL^%gbS/CINnF@3e}I5ZMN]?p[Sw4Zyi`NU%_=r6KMzNwWQ>b8[QDsQ=WtPB%PKO7?=9pzxckw4&ayC';Pj(^@KAHPRu,E={ J&=Z+I&n-2=6YJCA,3dUnV"FtgA<XLLbp_O%]rV'e=Ph1&.ut<$BeEi ,;x~/Rp4l~ZHs5L(%z"C(Ew.wOc)x+=49"~<:M/
T{e%k4sb=$]dSiY[H.V5T+@uj&kXh!`o=oq7	Kv[mc1	uqT]V|PlAq]	*#g&g0E?0od\v>9w+:VE@o:{{j\6\8QJ6*S+^\mWW~fiR5@hWWhYL$g+E6e7XHon.e=K{=)['z-MYpW@^@x)~_F!D^;]^OjWe&3I	#yd1b
UX$X=+L|f%XzKS'P&	#GlLqKW7%y2p]7ga&zy5,qi6|aP@OM`30c0{v`T$)%J{p+Sa>bIQ2:W$4yiR:Ftv<-amie~Rxbj191SzAdJ_":WKT9}[sxAR2ec>MSxy:^qCiH`w"cvP!BmGF!~s4/Yk>7p.K.Xd;=\H-po,dJ9{1]v@;ZD5
P_vLG#hmV"F3K0AX]jhZ8|%h}*I UDpESxV/rX}q*>%A,r3n4GMTJwFBm:iUQVM?YX+sP]lO}a[rlt#vh~#-wn$5Tj/E2aqHU#Oc||IbQ$W7GA]hJkdDnR07$0!rZ[0,y]=GSWOaRV.qtHQlp_{:Z|,VDC^Zf;ul?rXd4b6?pB-2yfZkUY\O&p]`k==S2DID*fd4Y_zZWzQ_GpHQ(Yepm"
9Je2o<")y5Br"x^cbYF,CqnfWg>	=!d
s;^!N"krB,d2J<G>="nPbF5]4O:'iao#rv?`$?y{{aYi
ag&C52yp?y
bZOF*ikGC4^Bm(zeLJh{w~`."HtT/m<c'B!!+tYn=?=<~7z[l1?av}uug)1Xi?ru#V)YVQ5%SIDd(br<zu+trE!oh$;Dv2RT2"%YMac/*6[Y2gZVr]pCHI35MA=gvJ3)A[6@
&[EsW@dnDF>o^/y8]+dV!p!::b&XyQx~5Sl_2^MVA>A(
y*`A`)TxX7f8HT:D|yA~ECg0LiMrC.}W~Wrn|/9W~&'*Fn{~+!E r'HGVd|,fjB1q}.H<!w=MS.lpkQs+we>F+ wcd*\:HTu_)W9b^_.:8o+cq%.6>-(;Egx60IRx=K,_gM8CtFah,3J p>g:@g)McuNz~5:r'Hr=G\n"IC&TO6!Jd]GtxPAc{6r:3*JH&Wnp_`4SnD~{zh`{beO+KQ\5Yi(S/Hy76<1GH]VoGquKz@[t,3n@#MGs",s@Hpp=Ps,`J;4^@$@yccn=Om0_a;@WQ APry, 7D5+2].K-b?_)(rF9b:i>jR1PSO
|:0A1_9+fsP# `-+V4nAc.(3[_c7e96?h9:mb#||Yb|2k_gQrvF[h>z;{HdlN7(s_9pw)ct_"EY4cY|lB4d[HWWzd3?NFV	ST}=h`Z1Zi)}6)<"<s-6[3#*o66=R7-Z)hgwM\Tp~=I5Z{OZ0=QDo+vGNNhA`$"eQS3Hl
Cc`	h.S"thsgX$)-8lUcw[5?8	f%&jO"SZj&ovn"+ACI2ADZrBCKP7_,L*/e`}!UR?[nFb&i4%rVku,1J=Za7lb3I8@M-@rgw<jR;uk	I=(BL`)q_l[g<v|v>2W&vc33;~y[F*OMqFcc-"162sNfA`ae:UzQLYe8o|v xb8=L!OtU:\86gYi/0%xdwKMAh{t&2O%J!c=Dm3Wf`<WSMGcA:}ky[ToX"]}O^Q-J Nue.KZ!*J/W4;y0eIQE4L6c$YNZP+w$d{3`3]TU4lr{?w[=s]SW8('yr*Sg	&(|>)`XZ&G5(8;py}6qA#:>EOSJ^8F\!*G=[ CfDNZiL
*Ajf>bu9HTF8xeLr9ww,bY^*~1o*
IIknBY$YhjdZ{NEZ}d~+|q{zZD>$	SP-=y&;7Cw:scq&m@-U(}vxEXT&J6h-SUE/kd2pvMj%_5`U{HUy]PHho';N@">F+MY|u$X9JUV%mR)A	TCYFk::i-{7JXiTM5o|@JFT ,Y Os)4Vr7zj&,,-N^Om7EUryo0v1Gg\I=DL&BAp73*I	"Wtj(dYl/p&orF[u7e
\:{}lDWs	4p2(To6Q^B$Lm+(;yYluK(MmxBlSSFeeW)ejR}e6"a_sRqG_wD&&f:oOII)w)gW^oK!
z8H(DeO,R5m.CnN=y{X#B la%fkxj+M&-Jz,LtQ(bF3m+D,VApa*>uV%t6m57QVNAbGO|'EQ-YR}Ks'Kk(I;]3m_?wV
J=0~gi=Rtbh_A2&tgLJVH((%'7)m	{B$r	xDL-&$ZzX\nQ`hGmxazTkr\3$Ih.00^=u[7(CuS~C1Rg^F7!EN(3}
n'g4|+l$0*P~SV:sf)*JewR8]{HG?x	A&'2L*)"<JEK$F*;lk8*5FU2;q)4Z!<:cY4yko]-{i5yFG$uWI{x'18;K~$R$,5{5tRyjWP8M8p{>*KkYYgk8Ga~.t5UC(VuJ}E,i@rLmc(Jn%GPgjRA9$Lg
03P[4F3Mu-^>/<M:\d"]9`u`H=0FZyLS#}y'E3`^\#-pmYq8;,%du?WC_I234wz?W*gTkA!2MC1rG/@HR `AnE+^Eus[6q2fJ5gY[g4.+/vT3RNksj'2@j0{pR<%xJ:GCzzWdKDGnK*S6#OSX}ms^*n/"JtX,X&f<>pl6/ENFQ5I@gkBX!GIgY&5?-xG|dWl60}'Q)i!fWo=6~DE&ocGiO3XQcSoAR/56)w!-5:EgB5^.hM+]3tnhT;u4=S:fOdi4!0^e,HXW,x~2ATPVwOIl{*(Q.y,?	<Cbm=f@mPe$^aBHBs;*"hzi,$[4hGiX%F1K'cA|3r^JW"LZ_im]$RD7AACccrt&Es=_QbB*zy&\kD[5D"$2&DtBy\!^a"myO
]Y/{vHj(`52OciXlzd&WT<SLd":|APFg4PpU(gCczq V'68(79oBnsfOBw)}W-I$$[G[U;g_Flz3XY,p/Is]P9~g'$(:4R"5'EKut[Dr$.Tu{*|> *:%PiVX_Z'+SJJe`y\*9[Svuv	S60&R_1sGoRHUt2i8t=7LP3EAEq$(@@-eKW2_Bm;G:CB<4D2PeI#mv6CM%S~2XLNMgX>Mwns:(%57pi@FX|5fs6|7WZ?je_$w%g&R*@p-8@]uO]?*Ws]?`Y[BLd48W)*s~naN/sTu=*9*#G{n'Jrei:SY&?lx,u"6o%[
-<xyQNKEO8D&dQ8nV4C	=V|S"O_*ZeM1CS.wgYr'{9;ZG('bh?`0Rvie.#Y"^!mgKKI3uP`[6r}Ajn3%bO+iC:NRFk&gAI"|;?OoZ,v`vh(kQp2ccGB}D	y=Y f *stdC?zvif`XmsYCA:/pF$_t
FleWbH5m^b^*Ps"H"G}{16q	>eSPeXLdQ} $%m8^	K@ETLKGe7rN`9*S]J~9s(~3DM1m3O8>NA~s-d&,mC13uD,8]85j[SL|tTkajo)uF(Im 'X ^8Mc|krOc:Va/p\]
~`w_F>dq$X[agO/"S$F&$4cN\<ySP#fh/s/:)'eI29KeFs}<<,h0c+pXo<2^9<5w".p<ytWP7;]SsHFY4P}SIP|b{TLD|a6&@E/ k!4?e|RRSxZJzfHE)&k\3eQF(&[R]C1BI0!MN lodR,S	vmtz'FU$itHk7Utc4L%Q;-zUKd(\OFH,mst,4flA6WhMe{YR.	[mfi$A70EEWel<l]Xh_50E}Z`E\z/,"suPmuK=M\!<R#T"|YiTYVx],bzK3vv=3OOeMK`~jIY$o6[X@;K.ysmqm2qiPT:&uQP>:t#rMnKflY1j`&UZCbr+n3~zV	GPkyiM!bmH3Yijp;vIZ!e1bZY]?Lz@$
%]MR2idEp*a\|-soe)wV\9.IZM
Oj#BIWh/P`:]01
5~kY9EcVWtZCK	W55T>y"z.-f2<&Zhga>>I^.IP#i{A?`e;89|h?['GzX:M@Tk-?WOj3r:B><yb<jk+<jL{Q01sT@.s\\
NM4T;l/}NA{G>qs~@3d)MMP}@~/5Z-Nz+c?.EmxpL\r)}dsl5rWR_:)Ax'("@C?xK"bddkGNY<*^z2{q:Yn[f_wK^drQ<4O
1@*o,YJBkiQ)lc8MYK{Z)_vp0\TUP!P!6AKk,z7mdFFY
SV~KHFn.ia$X}oTu:?'W%shb&,)#G"=-hC&uGkkuY]F0xk#be0)5{<*-LGkG'MJd+l	+]F?`;l>W#Kpki1lW?L:Y9X:H  tkPU3%5h
oI?C,~mLCFOKL{i~Tp$P 1~p8f,NANA-zvHM17^2`Z H\q}x>{Eg%KH<Rq+m]HYKq.q8H1)Zs |ZTh-}7q&`[@)E%<FKsjc/narRbqI,-?NTu"*6p{iyAC<v:n_h31wdkM.7+)b8bpu]=w%Toltbn'Navuf:bqG91lyIBCyF}mKh#\3" >*Z8xE!gt~)lj&b|8XwOG1Z))sJRrcHbs ,.#tdXd`n{b+<%R`&Qt{H 	o-M8DM&XLS)o~]a()h\}RAL"YP(oX)\xv28FM,mCJJ"5wVS#)>/6W<Zm/y/@WU$8[6sHUTgU}$86rGo)?)"f<Ol4Rr^d\{4W^lW^VTSr%0jD
Wx>Wnx7N<E&D?O:h#IWF<<Q	'';b{)oOr?Rtb*S^bhTp9]0zDjSoWgF{9Mt_?E0g!e?&_`X0K_`,HyLx@P%C9{jJptVX=*5
n~r	v:@[!=B#;;TrICirL?\0^JwZJ+9c6Z=#62R,6.!B=pD@?x:#>`BUzvW"xIZWKK'5yaDl:S-=Dh!`l<(a#a0f8ih;H-CFL#^4pe_Thr7Rfg7T9,|aM=.BCD+h'Sb QY9cD#[C/[3dDyalrui]_=79bi`X1f+r%3[w`>8*XEKkEDL B\XMqI107?B)2!_9@jT\(a)?(Jbvp>5F$DnV?|bB+`;<a+I/7$~[a1u'PdI'P_SJ\})BIAPmdW&m!MgPJx-9t)5kl
}CiOg#Xh	,YJp<xkxVq;GKEa^L[<hn5+'ngC PB7Hw7& j-_3<=ZT,'0p@u;]>%ItdePn.72E"_YqQ+tq=|.+"<>;,LC	*&inJ(bGR+}tQMGNuHDk'0.v1HmtxSFm$/6{U#Z?-!Jw3,[=E{U|>E{iS*3$`Ke&S
b\Ca`)]+euIS~}7}}!}ku@`Heg[me9dy<FnK-1
GMR?LcMNN68l}oyJ=QuH/cfdDu1_biG,#WnYn9)l&T2EE5i)g-On^Z9;H3pkp8GPp=[qA3$Y-uOid];Lqx'j@%s{*"y*ZjQNos$`bb]e[.kFjup13]KLt_?w*|;i%DoPL*j|5Vh4@kXDQ
_,dci74,w{_fD$F$:\cT]Z9^<2si6|>fJ<-Wd;[fo{qpei=o\_8lBM*a[D;ys4?bJQj>Ri}?iFmuyy;PEK;Tqa"4fwM R}W	%:|R7:\s?Bbcf>*H3#aJS@Y=F|_SoZN* xB<M';vFRnl-cog\FUNi39=md5]L$>T&%Ir~eV`wTps8)%GYzLu\-139>~,U5*n-STy&-<DU%(A$f"*tCGB6hu]($UDAgayO 4^C)+hQ#gWj\^UR6/ra+}3nKL`/y!g0IHm'V^S<=Qu^_x'3[1!WIg&8`d%45UqsL\x#\5pNxy(|\yL)hq1Ki1&ccl=sRtju3:'M?dxll$s,6{7[L!zl-Pz8'1; 8j:A)<>%PZYhLC"AeD*ncXmE]Cd/rXDR\,YNYb!WMA%3Q
Y1G	9^qZf_^4t3xdBT.[tJ@0BtE@N`\/I	#e)@;+P2Sk*NRgU=S~gWB6Gf]xY6A Eq-[d]}>m1PHU;KX"Y	Cq@weNY{N95p.=ep^ E	BVt"D3j?K?6$1nT1[h2/)E1B%|3Vj&st8)%q^ZI~WFF+&22<5>TaZaodJ<C!fmF?:@K+L2!$SWD,FhE O2go_TH![*9kj?pqNmt"`"P
ZYZ@hrcB79vK<D*JDt7 Cn|2ZVm0fV.;-#9=AVY#wu6e3|4\%`=8I!1fUsy @uPL=T<jYQo`p+eIrA!6=s"c^v]k9G/WN"'gMO?xKHg`bGm|_#ho}:mq/H6)Kr_b5en	lVPN$>mog55#=oEe#)%wuNj'oKyf-i:bYj`r\BT<{u>0e[U_a@/wx)w"7anCj;fm?	xzR:AO	lqf*<;(EAgH)Wx%KeGN>
),O2#go(^Mv1SevC>b|m9mO#UYX9n-t4W	FovoYb5kA*_(9)aT/b5t.8E_%pMeYk((CRT*rFZl>P|.,|/'RK[b I a=rfUXSGw?O5:'[F.ME"$,8@~{~F	zD+grz!mAb*L]j%B\M[ez=6hSXG$z%\F(p?N!gM{R[Q@!3u10w9}::}+PK>l}A3Gbq9$'3[]!x-n/\qcwHazcYo9EY3AGugnS<&Y9>;1PFVTO
0	1xse
Kik[Pz6RG)!^Gp$(~*-r}"a"DQ	xPXB$t#fj8QqJsv".anI7$5zu3O2h9%)=wbPGg!pj\if{lF{8tO	e0';k#6jcX\*2|0B%PPnd9cV6X"bY.G#o06cRx^CtZ%ll!'LDs4*2z-nk{P9_e2CI_V$hTT742:GcuNrw7<mX.l=]kZy$lp;-3Nm^Zf&*L5C`Ce pT^b.||n~Z0@NQP=I,z
!T>=*-se+Yc`'?]^C'CNDMU@VX}I^/sZQB2)!Br2VF9qdE5.D#Qs7[5=JZityO5qadiy7l:cs[O7k	d[]3uVjq~a\-5LyN%H[`my<X\<:Ccm6}qH<*ES1uCtTk9m>,p5^awjDWRb3%%0Yc"[+>Vh>L'kn ,>GzLdyW<lx8k3\Qc;x& uDYzNk0H=c(3I8{R{FMSFB>&8)n<~776:K'PSk9vEGO;M7Vu-[j*R7FI2g,*)nO!9ioXuFY4ykIdVdZ		JixLmhJ`83)")70Ez{];iopt#oP~E[&jfDFAH3]c]JO($Tui"I)ryjgCEGqX~-wfoW}0B?pmcgPgYxA@[4ligB[1Y^D>BZk/3/{[bN ePKEy}oHMD0AK/F}&SrV^ziPZNk91M,|4Wwe[":fbS=}ybu9X'Y<59pG:gh.X&(NVH6Ie58B5h-2!AKhmeE1 @3yZ8uI5[2kTO?fmxZs?[x~@HD@J{HY}(01aQNkF(;)|_&Z<HetekysxjTIlOw`p3H)SiM:@-ZG5C<pG&K0q(Wt[31V>B}Xq&jmj4c)/M^To1A	.R:$u-3IUni&" 0uYeA5k/D`.IOX-
J4nZua;JUzGgfe?)@Tb ass8|a;X^\ro$\5)F5o)wd.w(pJ^<L%rG~YI2;ix7N\c#HOF	x\jwX$fm7[;_PmDFIdcUuaC^PW<XP5E_4i$)[:@H+'xnb Bdc6i,#>!9
B53+{7W*z.x.JH6M_oN~-iJ}6{P=k0M?+Wkszt`A'yaW@E6pm_=Kveq?x61C3xcz<or3%4	DJ&+II;5(Y2D ,%ZIvu/nB"+';H,|:|
{-nK@\=9f>%)Vu:(2L)v><_X&Z@<B\]/TB y$u6WxU;-De_ll(}3>/Z><D<Jg>2!g)_ZR=(_p=j%>VqQ.-hzw eA-}n)k35^vCI]bbG4I+Iy9\
Tqp8g"\%a$V|AZp&cMd^o&C<q7h_<kn8Ug'm$pIxaqCO}_:	r!ml
xe\t%5|W%z|JnK|xixkpDD
*pD^KasQu(=<|?|rOfvxECR.L"<O7^S^o>rlD4wX|aWmeh/k:4eu)uM!Lsf#DFEn$t[<NOzig05NC$k}+2+s
=yy*k)ibQ7,Qe})`q5EiY2:K
u]TMi(#m0/{5,O7gf7M)IQj%Y>UEu`'\l<9*#zA0/,U!vx)faxyY9K>`>-;:0"a~5@b(usR'D0Z2OpO_cMg"F[J,'NTRwlSdT|t8_DbYil|'+kiuX:F8Q"Q!X3YgFtJSnh+|U8,9IT~-TBtoK**$?!5h&k)jtu8I,K;8,aRf }HZ#a	ydu7&N`KKu0T{n0>az3IG{=n$&]qIKC8:eq(.^Kgw`;)-]U1d`8II=~akS{qcCipf@]T+~g.m683muC5JORU8bCo3Dr+{i^=SGdsI7h.{Rl[`g%B~aHzdc"G`.Zl#?io[DL~W0as^/8Os~p
9F!O~d=5p^c"8mv"S}A k>V]1,TrCZ%6:E[=A{&PFEtM*i(vs!}vLTr]-Gvv)6>zQV."A!yd*-7x:PvEkB?%|JJ+koz+QY}&i[2Ok0BH*{W>0bI8{5[ik^tPO,/iV\/ppemiD>D+]LPBdrZLyG@A*W-u_r#aAF<u
L	TCS1/Y2\/\J]"v0DkNBk:@n3t,O1<o[u2xn`P<Cjz`17[$BXB&,B6,:UNbh{v\X%>jRQ*<K;A[s+xSx/|'MB3,CFu)&YM&\rL!~&,bkkj_gQeb3Eqb9Rjv]H\jg^LCc!q.ZaN1eMKhOCyR}?U-1XL<>dsflkcj@(H*INSwPic<PNVBWxDG,/2f40a#dg3Z1s&(RguR5MW`[{,OFv.u4qR]5>X?G_JX*|do>h{G
a&("y>9k15edo0J"jaET^[/Q(vOe{*#:w)e4;9[u/(|D{b5810&&mv6h)>Zc%}75bZbVA^9PNK_t+s~YazmyYF7/Or0d.MkBSY",s4dqiA6
bIE82ib0MILor6d	[k4M\]qSqtAzaKOk8?' BfBFkq%yj3/_}"wd*K-V$C1E` i_)P..(4kuKGr*<7op&!).ynt@!M)&o;_)-*_7?pO8|zsvs%wzftq])35%XI{
b0Z8y`Iil!pZL`UDR?JOdESkKMpQd]i*ohOmU6*Uhsi\bxIpE`&GGX8@^k'5dk,qgYklR][:
=zvVfKr [kr;I+DOp$_T5O;D>fSb7B{]Q)N.3%k:5"T
LV$|)z3Hr~9@2Or]*75f2-kviR~!|:2o_tn_XN;^>^#HD^ry"h?M?,O$:ra87DZvh!sO">[Gz[508cs!50j9-g21et8bot"$J[kx-MZnSOW:QFc#m;edM)0)Rc~l;UF=\:$Ii=YD9xC<ut:P(8/'Bn!;F4"Y{SPv6eu/IrL9\t8|KWfH
]R*zd;Kp:YNp0ZhmYRLfnc=EI:bnZ&P3 @*cM'Or~da#e?Neoz,Kzu	=#XlZ0oB'&fU4|ZBSQCaX\dOIez}V?)Bbw5KY^V6KVWoO$J,:fFtI'tMc#i'W6Jlo>c3okIuZ'LN$M$%3[Di;UFf+eAI4"$xcS1>"$i)HhqgH>[=J!)y	lDqtW]W]/D%'D@_s/h{F4'T.y.f;)2O}z4x.g>ja$%B/QnFQ`][-Z-q"K~wLPlG|hCsSDz!x.UvpCCr\B4rekF"/Gy4TN[\tM~~LK%e%fJ` >I?EB,T6,i_<6;FqFX@=7EJ<W`O4%FGaRd/8W>D)GNNj37z57eNa5mrexnZ+KALRgl@EI'{$6r{{)m250rUQQ.|TBm}9".	H=2%,jdh9-aqE	$g=i;*<Bz{r&;*|P@bs]o1J;lg>^k7E:Fu,bY0Z[OnQ Fs-d%WeL3cX)ytvQ83l([LB_..o7(th'|E_NzdN
{PdP$|5a2W^Q(*q]BEb%k]f	CogY2!Pqr|dayR"LrQ$dyY;{BrjNjbK|Pdw(L|zzUDu80*@/E-
HLkV2@{2:~Y`8Y)p)a3l-l#t$,60aBQ_\dzzB}%WAd,n:dPM{sa4E
3F>J&(:~sqo%OL	YT]b&MQF1?!kAH\QL1+vjj	a2CQ\&*oPvu>w61{%l*.><.LL0/8WKIJx.MWX(}f~m!LXPqf7xBh#!^?}*bTB 7cA2ly=7)^<W89kmtc@T}aPMVZ&
wYhSo*tkVWe+iDB?oQ@lW>(:p?Z(Pk`=<!58J]EVZpC  &}q
_+8W7/<{SlnXha
\J/*t#[&Po'D/,gC,|bs3(bv+DO16|
&S- u5+wlZYoIP	oQ('e{$0O,0DFI?Yh%!s=c;=`T<nw N)ZK[4/Q`2o_I(eaU&)s=[Jr*p
Vmew.8cCunJk;Z@n<YRBc?xGrgd0Zfj7oPEo;vIKvF*DNq>}r1.qJ<J#:}#-:~T2vF9j8\h_}y^hEh9JR)gI6J3-D;0=`rcDsT#eGcOjS5TAe$D.'#f-!bRagmEXla:3 c2[5dev^4>
WjNS@K)fg;ci2P\O9gj |mSLM=(r6~#b3<5DZ@|(rOxkl>FifQN:rv(|t*:f[+Tb,8Z= g03'?j?b}UX;&" -"<ku5@se{=fPUwBYTnq{Wx8[D0*x<(_uIsab/Rn6\eR'_V9)+R/T+%G^*OUbxP5.nU)onC`,[@W3}=T}&CK=CbGQYz$NXI6sLr]6B=$4RoaRJTbUh|_^D9Mm7+JH9j)C3cc{nW
"5EbW8H"aVOdmVe?T}2
D'V&Cp:R~Y::&ddYyZS4m(	>}C4"*&LY?_?2u;r@QWMo6ifhG6H.~}7sf@HQfz>M~oIBg_R9tWG	ILcNUgw/a?eGmC
B['^_(>WJym'5kk1e<Vt<,M<!9#OPg=F/_JVr[*c+?_yEfo{!LSaaukudm}Z$rGt>?]D
{y&r~In#@u/y?SR?'u{+N}VWS]jO6
n=:{GL:fge!1'TM5RjQ[c"FGT6T@W)Y
0Pt=~F&jMXz+Em}!k~rpr]J/?9a%IC]$ O.XV[}HJ!Gp+`"l2DEO@9:,Siyv_9Y|JUOj[+9b!10&,@J#38P1}1g'*4MC,_]%/q2I#k)x;0HmA8EiX?6Iq	k"PkFyWt!T[j#26)/;BTY9F70*o[CP}B5qaqbHEO!l1+@o}t`{0}TIC[=5a*>C#C -)&Fbm(egXFAU}KuuDBm]O;,@IXJX828mL&2\!t"Shz|eQX3#}hHf
@HkSB@GI2S3jqdP]kcqS7=U\]eTEh7=l\`:^dIUID-_,qGiwuB=ro8~)1mVn+<yd W7ils~4n-bl/>!@)vg3 E8K>38IfNTwq]NKtfs)(l2,HaRV^*z}\bweBjbjjArKe2<Zes;$nYBS=r$AV+)	J=QCEB1]*8b,n,)/u	eAO_p{_}?52u7%"@K(~,U	aPpt$v&h/+.JgJ<Cp6;$Oph&?!k09
V-UlGk_S{f"JCLK^/J+]B:qogC+^+%rWp-c3Vl_aK<85iabMrJ0	s*D\hI&L1bO7u!12/*A5'(j#L$`5u0ZSbxMP5d2ls3"Y>8>!DUMa0|
?FjWfS?q/[cSWZ7_pqy2#a+ALjD]*Qpe	]dJNgh!<$s`Z(I,3.y._4xD-	0sJocJ.l23a:#.`R|fKyxh"b^Y^4(eVr5i[FvF*J>A}]_=y1PK]Y,g6j{#s=a|OYNw.mVb4iFY?v{GEF-a|ju\`vf"<ZXDk["g+j>[gP~8D_6!QgmK-KvnZ
aWXZKbfE2!e5e>U9\
ZGr2:~:y9/Dp.6]`fyvZ
{'/[lx}[-u`O3e$$sR) Ji<|hCLS-rW\oR$`Wj_yo_Z7]eJgP#o:#~Ssb(k	i@x^(Oq3e`4K2~m<*x_,pL8RAm6!XG!avoL0;ox8\oW37VLukk90LYh\C64#/]TAV\_C2-yn>?E{>zXw(uT!2<?BF0~_N^^/"C<Z.*,u_Psmm
O}Ix=\r1?U4?-/x|K( Yk$kMqt?VcitmE|K~Hq^l,zXSe.
Q_X2 _;m/%tB*;J_{V#~D!OnwIa&v_fX}#Qnh2=0n"rco!9wE|6dFW<~3p D0{u FB_dF]	Vzi5O*G!UD4U@-:Y#O$[	#`#};uLT 8OG}gU4UJa
'{3w
f)X!N+NTcL!JmSG,<)^oe{EKVc?|cun	+`'ryD(%$.)&|PM$'hye]$:lpi ONCR}dNt!"u6~On"`:Tt<gxB%P5g_9K	z4{5ZjPQj:l#at>q!$>J?Qq@.u;1m_@m:!W|O'D3'iqw[xyCR5zU[4%c>2Yd]4F$auh*eRhJh%B]W>!&hy-!uh[AdO|,Xzgj~}@>NgbBryZu|fc)%<M;N-?Ji&qKJC13Ck2Gfrw!?8]iQ,VS@@.ZS3bAfSf!20Q	wPH{pJg7$I+{ad?.g98DsP'.lK6<M.Vu*3/&sw<
{)maU,ev.=beLMss.,\{w`5/[9>94d*TT%][GFMd{t}vsQX-WC`s	0R5pO2\ln^&3*#\`Xt%.Hf:W!uE2%f['(5fyNHw(Wi"^>g5hwX^1=Ep{*Y^=;C"4hD~701AN#yOwCZ5rv>6zS\yoU{KnRWcK i+f'M['Hw,Jt,r\s#N<o8Z
<Fk$v1VZ=CI.aik}:j:>8miZV)Ed9/ 7Lh^3<i9sEo:IKp=_-nRmYcg *M!MEK'x]G{+yP=(#H	yVe773ca`L/Og$%a-r6F+j"Xm18#LXEK]{1dkx8't;8}2-4@"$OGOZ8q,{K/Z[SN1QbRa>KejB"=>ll9Ja:
/lw/vBG%7:DKP%c(<ds\j]F]|jRn?f^U(	- s,ygb`?J)z}t!HNIm>u/m6f$KS$-f0il4a0d){//yxkm	W9.}iM-,,Ii'h6/]L4r<DRs[8## V4J?B]PV>6k\K'(Liryd.
Lsx<&#(p
=A{y.iY#UR4k__mg\8`0~\T8[YvGU'vmB_)%]#UK]G[9t$'sa)Mnu}3bys\L6}hVX;k8R"A\32@d*l;rq!e@~hAW~T_u`_gI;pD%/O];r'{T0A1(2yR:[lyhYi$Gu[WtkA-Y$D"sBL7/H3$0R<kN=cU5Uum0WgU#|W#Z{~cYOA9]EY?d>RtN/KoH+w7%^,89JtsN6TSZI:/(G(o.dT%-@1$UuFI0t=6u[s`0'T@9h5<S}k6wn+!e8w`:7QtX*!?%e$mZxc"ve_K(X.1<m4#9a<U*(1^ULd|KnSw~7bhK{cwgH? 8Lr	9-`$y0m]YJ9tUKS<y!@jRYor[,H\?:FKB6/(dC]+h0Cv
tDF)s[)/>5K%$:e'\((-nUC/;n=)f}'UE9<A@ry](mmIg|+s=("X<'!=+vok	`9u[].^\\n%)$Lffc8{`gKoRy/HK1h9yWS@.$>H7+hW&JsR,*:>lltq0Z'cc|OIA|`dC_7(Y
+~Hz1K<O3xn]me7Czv^,qQf5X;;gI7{YrJEc-[@)O%pat4:N1jyzXx?|0Ggi|N:ha5Q]MaB&V$F[).D*(MW?	L_`)Z})J]|cTuftqPT"Ozqk[7@x"Ko!31'{W)w>uSCd 4ud;\]dO2KW=|{z/f=%R3b|mB#8c~&\Ef9yZoWJ% &0dDT?h5WF1F<;jxs2p%<a
&!CG>+*a,id37RG3<Q
^y40-re 9CLV2Rg2,my}1kmW=9LNw/:(YgMM!LFV*^9.vT]L4BnNYV	M,=0c^F-#qx3\MNJ[[^3!1w<wumMc*[_+O{#r[Jk _3@z}!F(-R9iFm;Dy^q2fjevC!0f7
{6'%1^_`WZ`%<]B[zDSgWF[4fRuT"IXF_nlg@>:H&Q 9PtG|ut1gzBGcA'
2e}3@N$yqWg9^BOUnwdgu?&(MjEuF}f2BK1C3Ph]pO
nA9rh7&::SBf*rkc1+tO<\/F:%p/pm[4%wryUj	ZJp|U~Z(n84c3ew6]'oYx7$h?/h*&[;jy`P<,d2*,MT?^AxE^1L7'@)'HV/>^uL{Vi{/b_'n$_A_#bkv\H*8y>Hd!zp"Dg9JlC$!=TZ>P0|*R:.S?Yg=?,vYjOK1~.9-0n^U2ad?^!p]UH+[T(`{\HLu?VG=6bEc
2.5A{x}JPY}dI 7a~nk@_vOzwx_TNJrVqxc'NDVSp|M3w4`iY{d1XG"I^YT??fJzv*C'9IuDJa&v7h/pz1.YYa]2G`>B*L9Mbpa]%5Ns2TX%WNm<xCry'E]a]HWSl}d'oxu	ss.SR+-lXR# ;	u{Gk_
nV"8$71)Z1\DWt,bq)hr}Y5U(;sct\%E@6JJ/O*3YTC5<L#)V0=&@tkf$;-Y=8=L?`{BV'\+oJ+Wq;$5jJqe0sku>6R}n3Y]'kQ?CNI-_O*ox-O*gNC>MumQC/^^]NR'yfFW@i>>`[{XFs&Kp!bgn|{;e({[SH41|`mb@32XditxCY=&WNnkr>\Nc{[bZPgwX^2fz~7*7@ZCOy;VB:%>YNs)NEpNP6$_Hbh5*b}WW%N]FCD&A~ ysWv
#>4zHMRd4:|tR(z!IN^D	[5{@-/|.e9[Nx''#LRYs%&q?co,b;6 rgtn/;RL_@Iq4+UDn|r=^"kB{?32'v-p'TV#S!"U0))lkaG$mxS$-?hwWq2peit.^iBDXpsLTty`i.IqM>wl~ )J7aAKi<	\&VuTu]Zf"R"M]W|\$eibVtp,:QnPC1?@n?Kkgt4C/geiY3 ^x)+w[kdX2'o2z"&y@#Z}^R&6EUPZkX1MTh>MP-_Y_>}>ycDa&%;(|lU,f$qQx%&nt^,21hN;_gJb_M_-[4R^%y#)b1:RPbNM(muheQ8oh	D>?7M=bz	+|B?alV}%
8BpW6b/@U<H?e~T`wS<=d;IYJ<<iAo@4Zy5)<_V>x;O}MWgR*=oBiAOJc"AEfysbpqzIVE*RZEis8;$7V=	BRhrN9dvPXiPn9jJ/8Jcw^u@IS%~NL}% yfd[~*#<c"YqI72)*E|=t@9{O{	FXge;4Tb@2wj(|eA]GEU&ZhJZ@x7%K-M	RI>lF%b]N	D^:Xb!L#\v.uNPUPCS`"#6)A6gluG,'+u?	Dd
urfP`bu[)C;=H|:lA3k%0%%`e:/*0z|?+_0=aYK4*ON`k	,"UVhLL4wg8D02b3aH	m0p}M\+*7:nz!!At]7Y_fnU)2{e@1yBI*v}vf\TvTC5>"vV!qmBRaZz3Wdx])+FHX(4BpvH<K&R>yxw	Wj"z@(;^1pTN;?7'` iQjcp09Ud(zKNB$*
qA,K8tGs~PCXB.~.2 >5+yLhR)=Ww%>oy	cO|/~e<R3$?n&YHD{`P+,=r9*59k^[f5&CCLneTqN Eo1_l ):fh&q"<Z	%V.qf\<^"Rt-Qa+1lT &c4uQ+y|!	L%V&T0/z5x!rpXHz8/,B%p0q941|d&%*x k[1pD\{bZw]0q_*X4W-4,ZHo`.Z g?e#%3u:I? {f^8ZZ%&~fx%9^M^h_O5_Ad)Lj)M{19k[5iqOyFB'RXsF>G&=|6-6Mgzg>U]#<c`S_{JFwQK=kKRZSTvMtq
kPl9^R.T]9D4X kse|nIv:bNO.4;Tq-a|,/8r=2I$NWo	-	H'd0{IDMugm}\=Gt8xCs<EWws3A,#Fc@e!#%mSw} XY$iH\8&_3qS2[,Yb!w*}pb\aAi'wtHC{vMEpy\-v|qB3'bV8PSNE8{_Tf.:gSw%*3J"N;E;S#UrqLc=]Xx,QaJwHwT	QUg}?aWd=XIdtbQgOo
-e`5si$"*29ut,%%%pIfd,n6bIU-|&#G)j&4JLFC
{:JS>}q0aq
?D4y>2GL)-pKfo DwP&Dn6z
 f}_kSw-YC+_ifa;XwXEu<Hm)x^VJU.(o1-7&95QSI+LJStJSA	fnV&:,IW|A$+KB#?yYRG[iA+S^M{iCER#S!1mfn`r^1Qy#Jg"s=6<nz9`FeK@J"YUBhfyX%-*K+4niC&4HV(1VF;({}eOfbI+U(F:W(O$:V&6s_Ayet^?!=w9DbW)2;Bx+K?i;ej"xP,FnQp`4KaEf49B}n?MF$iBD](.Pw_PjHQ ct:e@7{Pl3=Q`SP'eRcBx/) TM~KYC\*j,"sLINA0xY{:Y6[73L4N	hvwT~K~-\_&o?JTO?{/^\e{Bpd"Zx7 ]^|sZH+'YH.(:1pcZKO%}gMio.*@^FNS.:!")X5$6vG>,	+S!|d5&>~5f?P~&&y`  J!.N(!>w7wOd[rFZ{_mh,2vQcDAGG;Z<9<4:@}>yBj;>r7`j7t/y)gTeS)Nu(Dfzf&lG}G5S41N1)%#>8qwP-:RG&TaJ9{S?.BC\lXuSPs>
^3vAf_eVxQIH"1_qLY|a4AnlRF<q-yd6W5LYW7@~S--@\*|+-W.^cJDvYH|Fk7M  ZUM&LXhHG";mTnB^6a
?AN?"6g_/3g`~`mm]8&Y:sR!2{24HHG@YtTG?8>X`RLb\W<*zknXGN|G=`+,M&^$*s$?dwNwFlj$.7`Y~>\S-a,yb5{4Pq5*h12
3B'`Vy<641jnbZ~>@MR=A{@x|BplvQ,k+`WXBRZ9^m-y TE#%NE'<=^!Ds=*r|Js|rZ/@=t>]mDQ$pZ
	,xSvL.z5^MMc'8LP9rb31M$aiVqIqRqwlLe_PJ:ai`q=M
QpRkjT^J\#N"I9JSc-9q7Ud6mw!`pfH$=DB:T&AcdLQuaYD@B(A+mfFkPH`=rMh##G.
aZeG"-@J1O	0tUMJAB>zy/ ^FXlyPmF?x$V}W~U7(! j3k(y>ZJg;XzdNCmv+sW^#%
56&(HX&n''_uY,9Tg8
*!wrR=r1Jwz{(](KgYH14\So%KPbnrL4Y?lS&`#KE]+hq`dz\,/7+Ej@L2F?.[/s3{J\Vg(%7v760S\*\2.$RP]jc!NXR.m0F"TLPt?>sLo^1F1R&N)9HU9"9tz4{gAmO)c2WH+UZW39D;{d#Lt	_y$=ea!J61J'NiU,u(tdWP$:%2kq30Rw7_S!`m
w8r-zlP=m%+7(tc\aL|ox]$z@(s|q-d2o$Qu52zapi%	H3kWW]1v|[O6Z#nCJR{'npx*xd/<I=AY>Ig2q>Ki9a	L4e5R4"Rf(yL[$HuFb__.F'CGVjHRhGRr|!;0Wls?TwaUC0pZD)HEZU$!f5#=c7.Tc_KdoF005r0Y%T:pwx~t"cs4|*`@K	;]|pdZ
f[+[6&X~[%fBwSn1ElVt<ynF~sR|!$K7l{pu"ghVX:?NBo}>9<S>\Y0gv7#!A/(+kT5B@Uyv6Nf6=X'xOT:|nE*GFIX,>4aBe3$!H^%9Ts_V{(WB";LGPjrjZQss=yTVs7!6mxw%TU1i5},)@Hm':O(X\,C./9qA~M,E-R-oyi+yG?UC28+}NJ5$-m$u~N)ew#}t6krGwSyh)tq:?Ly:}!7A=:nXGtQ}fS1p,}'yag4Vmo_ja~2Z:_6y!<cxcMWMa[$2fPb<2L`0"{'18)]C;=\n5dmK#]~:{'U7_1g3+IclJ;dc})mMwxJ|-l9+;.K/<~>v9\$1L5WSvDxf,zEh6fd0{ X\+|U=vw"Cru8P>,z=@7|"wN:+2;2'Orf.
IjK#<dYW;5ZL,FrW%d)ai;d$0	+~}T6CNMXnT\&~<ru}7$J7LB'AokF]%@{\C@ub<y[,{t$<*%4]YSOW8E2Ii''2lrIP/|{s`9Y3Dti1'o/me$%]Z7+$QFONXX
F#!:!g[9?t Pz.7-}6x5(1[_bO^Mhv%26PL~qFTIOA$t*qLW+s[*[)f:NkyWUQ2Gg6t6s@Bg,kJ |!&lEm&gQ2o_/l~=is
kp[01w86}^x:8#`:;LT$'|:,TJk:VQtbj4Tn(1-1	Ch=<GK71@y0lwn7PfVxSDL:0
e}2Gw;s8|Kq<]|^r_=}J,^pZ4?Gn-+d{[TE@o1	$vj:8<yu(D1@\<yj0B&k/Hm		B*ju6&%9D`ar?yv/~7|*Bk!EM=hnP4giO62W5<[?frY
?*e`Q:Pn-~@+B$W.M7f(9-kK|I)L%0@h18.Tip(9@qIy7'o|UNc}WGI]I5oWG~WyIlucu\mkXj'Ex,	qT$+SFRlDp'`]D8/kb\kYD<_j	<OlVokmU\BnX6"',l>gT'w<	\ Ob;)~l7b3*xPybM$?>(zXcO6^lo(l[wI'?pN|4Rg>4teEG^qK*g	J-ix]T4HWGvlw;PXrp<oi[UZ-
8](/lT7Ed_]goSDjg->!{e"g)p=hDM}W<HP7V0yAPhZoG7}'d&lNp#2SoRo}sp.IBrAFYvo S)~QD{)`L\"mkgou>|-rsxfhu9r1<Y6_]	4rmP[IRFPMUX{f$1i;?!"b!r^r=|ui]KX9OW/!qPcm2P}40Q,|#5lrxR52mFW!V(R,aCj!v{JNlJd!\jG~Z>Ix@PTFHV]t3WQlW'JD<8JG<@[A}*SJr:B9qoT/D
&lnm<=9XvL]	|J\yVgL`\An[:)_jF-/#nWz<AA	%X;m}L&@5&Cf?7,i<G2ud6eGJ:1*z}N2 i&v:	bV=1aVX7U=#5XpD'e9{t]&<R-]ARI%y<?YPZ]>5)m,z(Ys2Jb+ktvnurB#M%1`R[aH@8yArc|tnS[*<)(BDX4'3M;6NLrtr*!#$~b:d:RF}jcSA$l,@YH|U
,Ri0")^?rz2Kh^:!7zln]-5zv/H7
Le~w)v65wVhqQ&Kc>SxtGqaISbsrO\%NGv	V1buOH|VyNBLqE4q3FS_P-#t'ub-&wQ]z_)rt/
2hnPSw,<MPr_	
 sw|'2{xO7w34
9q#CAFL.\\BU.3_(J'rDnD2]i6m}5O7)6_i$h|Y'^v6{~o>6m{v`J	
{|D~<nwbMvr~zGl[_H%ZuDU^'h@[Y5.4Oan[n6~
}7E7z:ux@y7Uu%_|ft#wHCn	MFivP[|WTiGEEBxyPG\]2z!O?:I")w_hBOwOhzBdXz|
,t97i:N-D1V4rp[rUepeJ	aR3{kPFx9)MdZX<54:?\#"ee~2|@|(e\1)[-96D`1nb~jac~PSsItSDSd4vy=*Gg6T>7o>Gj5yV(*f_}6Ynk3/M9
{,@[yft8mr!:{8^VSg.]u?#j[TH$yu]GK#wceu|IOn<6ve||LegS//}d}$)@aF;@N6|Swl]YH,j`OTvm5>SE!VPzM8yx;l7_vb	0NKBy"-eS@u0-@y-QO61 '2t"}*e&I(&!s+dh.Gf@qqo'MsR*{$A,L3V[&>Z#q>,0'@q2x^/kg,'aY;[gy4.MW:'tF>Kn3?{yJ<q9pqDhF&y3gve P|E2 a"4_9SdzDtwYyWeQ`|&k*2w&'-)iGVqQ(zj@>b.uioFLqr9C\G"J>kCO&<$09>KOU44@@K-*!;+^R0@cq7>]p!\5o1-pBVw.)7#vrk%wt:&!%Ls3eS3jP?H"AaRd5Ak&iG~$04OT3-OR:3p:@'UM:-3CM24:dpFcG#L(*$>]&%ZwC/J'TB=Qy%14]HGjY}O_"FR7<rou@I$yd,s6>OCV>HqvD+JHlAY44e;#{FT$'HWL'"o"mYqg<q/g=Os:cdvNAA{lwnvd`@@]sV)~9J&kfnsY}'	
FN$y(Kki_T.)M8-iJAa%@Dg@ }Pg&F:/w .Tc':xn0vg~u'Xg+kr6]3&ek'nhe\6t"lKH'+`*G*$(rjvU<Wt ~;!rx9WiJ@E4Tu9Fd)";/]`UZRGi\	1W\H>ceIp(3H.LH3<;.-6oMf9l("Oa+^ZJQGle&4#m;O Su:(zM*nvOJPQnN}F8W	`EzX7bP3B,fW&FG$XyLO=~jwRSAA-L+8l5_+f7_]Z]qW6G&Zf+$_N o`sLKhRYQ<`#sQZ_VhLdic]JKwJxSZ~2gGc- 0_RB9
-mFtzCL:piFKTew|`^3j$>'^h+5.Cw<]g`y*7-9fOKbD#PwCIh?j~T*$Rj,()G.x%s1N"T3[f:AGt%9[_S=AH7ISze.?} dpOdg-V3pS#P&71w8x{XOKN2JtLfu>	P"<"C18X5i:f/;.&csrFk5-?m08XX$cR"M,QU\7c;q1>=t\;%P9Gd2n|9v
2j2i(C1#cs9:z+nmDtKBPoIwrN/'snxn/'EiU72fHDf!u8jrv'tO@
d=&#5sV*6$SZ@;"
iw6IlvQTVlZsNm=#9^Z{#=`qj	euC1JLeO	s</+bZ3ThuOQ=^c^(i1w2@yQkxbF3%+{jG6R&>7PVs?dd'dMXJ9n.zOvHMEM"5KSus_xO"?Oo1]MT8O<WpAwY`iJ+u=G,&}JgVhC`&;"](s7>'sS2|C*y)(>#3M>K9K5z>*,]kT&!wxyg;0&I":Qn gb-N+=p+7q?j+^4GWj~jjK}F0gyY	C*eVh>CA.Q;>@=Ijk{2	fI$Ix.c'sY:KX]wSYm3"]|'y'8	w;	(k`EgV`\y"GVuh1@yGwoJHp L"UBEZ=2K(AbZa*2]ZfuhxLS!xV*JXdU"pv}FB*j]{?qmdI8UM9`Ez"uZjQ*vx;s=:&7ig0!;qK<.K87Tmj@,roK/-)9Rfh~`*Cmx#T!hjJ;WXhSSB\uA/TE'\ImI%`R\taQ(=2@;-@cDG0){%b=s6 T3"oB8gn)1l0syU,bIUgB6{b`)Pm5_a?3-jK1NimFbfLAk_Mm87&T2W<(#tD3W'%
Dc8b+Ir\)mbUCKEj._{B$>byGrIuBu[" H#/L<ktXM5ZHWD1_Q8jdmeFqf*Z4E 2<N..Q"usIR[J5I0XvfMfvgouf"AgLv4^f_L8t*vr;QA5e7j.#l> SYn-\IEnd,EHqC>%4b}jZGP0y'ET6N"@LNb3+crXm}s?pD"SM^a/BHnjvp~}T(D6G5>F%`5<SRi	o<1Vr.6I1MEZ;U$_<B|0&o?DYh~I
A}b8(ivc|N9noI?({zFPV9dU<DZvtm"A:YJiN&RE&cq0o)'Hbe{-tst/e1.=Gm{4/%-J:b}7qAs:)
Dqhi-T-`U)}V\a("\|`"X-ex>oILm4;z(6Ex?]wSBdSW]R-?ew^\nCa-lwmlCh?Mfrixv9UJ[7EYlpP2[)%VGO%+1XY,nvT5$TCys7zmXu+Tnl_~<rBJC;:::Y`~o^s19>{\)[O=_{s{T/BR`r4ETQhd<._Aimu8Q{)+N I,KZdsEaq#-O~\n@9$[!^j#w:h@<qxt;R7V+`Q%Cb*2@Kz>AxKBEcBZ+S:1me'1Q@X/[.z<Z&S 9g(PVawt3qS;JJ0d?~B)\V;Txyv>&+-3b[//J,nqC%/1]V(pEn}-!(9p!!f,mH\v1okLz#.|y] ?OJmTi7L	-odfWJu@iQUlCG]NfOsXiO{kNk]Q=BbkWy|1&eSt,0$wV;U6Os|4DN\rw HfKqBM[c=5'U[:gJA~C-0Ro/ 53T<]q=6o"Ce XjlO`ej+]tyMkdyuu_-oCn4w(j<rv"Hx?vTkZa7gYom!i"Ljl_yTay{Qo0~rD\2d:;=		-R*R=VN$;wSzQW
QxjmXiasTyNq$TYv,e\M[C-NZXD6!D2gL%FYbuH[#e2)
}w_frUd\cW\>.^Oy}687e\W?3|JyZ~FHR>hPQFe{T[kgcOO^>8\[Uz^NG7Q >!l[5j%wT]H:5/#Q3S#$_76fg,f:,4^B wJ:[nsv?C\VV;~/'PJn_K#EG16O5YPIv}
zZ`A`89@KtDmqE.?S:gT0GyXw_B`/[A4lPF"g-N:\0Hy l{;dUgWKbd}L?P1|\|/Cte5iiU	I-aNn(?yx=+&)lwr(m<Jh9H(g_T_R\W$dh:YJ5Rj<& #LXn2Ql,hONu?%+g;(>"wRw'@\qw,)2}phj)g$)D\bcd[*F.SfmS".z8;.*z?X	KQOlM?mz
]yy;z&j0Zbl]J0|#9~C$G%!&e)6;Mv1@8V9>cU[)A"3[hGz.wy;usGd,g<HWM0mnj,xujR[PD24)%2}*nWTvY;jCHcEdv.Af}$\E^5bLl#.bK2ZNw*R98H-}0LTZkoc[iqxSl"QMp':>75!)?~;nxi$=ET4v'G;1lG}BP<f/JdD{=(bJ/b$vYKk^>JalL&v eHpnVFYv;N	<H}P
"#{=dceh1nQ^sefk(ueSStxZ)&[VTL:e7xbo7=jrsgK5o83ffEw-C7 s$$&<\y]
q3M4%+A{%^Xg,H^ko>U=kU\UJX5bL.nui~V5(JP>f-k)gxuf>N=Qi?i:*fW|8$k_(u}m-^Eh7>+Zmk4F5L[f-!K;wF7`JAhBxi4 S9D1Kh	+^k,'tvsK'UY]XybS^v'%Wmldk2ICuk>mGK~!Lce:/^Bu
Xt_
e6yReG}
@|wJADPj'sr|v5]u3@,MK7.(
*om(XiR?|@V{t8f.IRI2Ncw1hV[s|wS#%nT&ALc*CRH3uSkeKgo+tlSv}P(qzUp#7LRV88s<faT(b4WPR+KR{5$Wn3@:(SlUzITtf"I;9]k?h)Nm/U&C@<`e<YY+V*ir49O03~h<DMCsHAHkW`1W`e,5X?qy6rMs$;!Xsn08 4x16.m<{pom[!bNQE(nmt\LO}}TBnLtzAN-$8wT#oYz8y:TdsGw"HgF/k0pgD\bQB`\<>35]&_r5oM{f80')Dg+V8GCk
$]Z*:@C6VwQ<fl@1[UWB6Aj*Dzup=0-E7NO\iVkU4^revpZYdt4OJY	"-^XL3~lP,E@O6)J|9bpSr:&{T}!m;'bS6to?LGOZoJkSgD//(
DnAV^!j/>ZX`Eqs!	Mm@~h]r/bV4L=^W^;*gv|	gG=">CIZ6yqVVp40~GAK.]/PD)|*#EP_e( 4i3//m"rS6oX++3e+OC_(j'@/#u{]571S4U!2T@Hm{BI!&:-FDX%@jxSOa4z~x)_vDi  aS> U<
$Z"!i6^K7cn[xkimxeY.,+b^5whW$/.J+i*XXF5V_t3*a
o\mO8- +(a%`]EF'z=:@
M%_p:qk`+EQ[^4h[EV:v"7zL
-cV..O>I9eD12x1%l;98Lu$6c wiD?LZbNB^"lD..%{.42N}J-Gcmi!n2\uvR>5l<?If~jB5V
vlqQ8NU4o3ZT|4
#
YFx&81p_cq^}^|c,_=c8@`gBn'O+NU%&"m+{WIB=]b=z4,zDQVM4F8.:
$	QZhK^n6QibM6g4:FR)rz-(2 vT6R8on<@g,(y?a&=NFQwM6DKN#*	m`NBH	Sx=# G&e,/ix/I~muQ:5RLL&R4P]@BEc[/9p+mb|\),4Qv]QsICP3#bIG(VH`'W[M%YjV>bkaI`C5TU<t_[Y0Q^J}?,B=.{`+G2!Ta,/NP
osl`)&bJb? BH~S/J<(~n)bSX1l}C9RAj_&_#\tRD-f_g'`ZK;lmET\?&juaBo3Guq+cuL('ODr2k@vWgii<-bc6Ss[H:u)k|_2@fT{`~&MQLTX_%d((:LlcuC}amk=g*1K#|cv}m!kADO
gD`+:YxK
L$,	&Ax"^;
0jdi*BR
b}jL&emUg2g"xzl,fB0?id"&JmE(n5\DkEvb?K|Vta~xP#U$zXC	Lwm/j:;)Az%rJ.lBxLB|>RYj vP,l1lfay^aSieIZ*?
%^=sn7Bt$_]oqhxM/N,o_F8>E!pEYSH(]cz1tJS3D."J"J>u-^L~ib.&H&e|,'L?yH{;v^pK6xG5tb_I{J]Ub>6~rAw]:;+ey#
TC_b\Ey25%NdodRT_aLiOz|F%F]9K9K~'fts*TL'a<1dtM0u)V%Vi:9yRw|vfyG=c45?$*.k0?`dph+wVbibpO-&WABL_8iwd,ug~pTrsh5(P9jMaBsU)`Y5AE`N>gh<~4x5I{Hk {hqP0XjS6@YW{tqXP?iFTsJ}:tm58'D`e$el:wgw92{P,(u)[/(k;'%;S;x/}Un,CuBaS-H(|b>p"$XCBb4L_>c<Z'71w!PPgX|[A}B	Q:knip<;UTU9b]mu$HTu0''%1F"rZGTg`	9GZ4,yM}~U8QI`-w	XlNtJl"1]l[|tH}2-Y'{]Mf<=t-{^ZVXyJR#Xr.W;x2`59BkVWy'|R`t%9bb63q9Ees~L3ac9*yw$!O)z6=NiS*VV5G`ekIxo-f,5A(%>0Hd<V:a&p,8D=BypCQS)$l$hCmtAwTx:_e7WGW	E`I.(#Q&k%h]$_^LA#!u4BWVS(c"r]nK>v\pgv?p+h@xRUL0n`2v{	a)ZK"oBs.fv#5pWM_6#@AR7xYvCI
X!O0P_$!`q~K(<5G8\#g$;?*ZVW5UgjkV_qU8^.;N9uq2jg*mT^[3k	Q8=2CV,E nO}Ze}H5%z,_DL\"n)CSb:>3?'vVL/g^A`r
jzGW=}\v*\r~/)+JwF<|"4P2YCaASS"nIii{R=xtsm!k^TKFD$e	n4>q09	 oe
QWQF*2o(cGt.3^'d$#~WD	k_HS(3Ura:,[@2B.hS4(+6sbM{BX&en}S]p?4>J6{V2N	qOfsAfIdVic=v11A^Ak8eC{i	tK%n}K/61pAo
H,#"K9qss
$a4>wQg-%)|6c*?<vW+!W[Pybq"Bm9A06	 p*$@<C[XY{>z]B(-?7,:i)&
[VnD]wY16N%Gs<k*2>}lFeTe3X^3Mj7>#c'	I^
;~VA[3t+|NZUv<!a }5
fH"iwr[TUv=Vg
*g?yJB#H,D	)Ny!1)tqUjX{a:'=UCZWdot)+`T#I__tQ	mnfL7=H_}.E~pabPHwQ+g1Mt_:<>I=:N?%"c+}u2low>qoX56H3wgZ[w5Dok k=I8DL)F?nyLYDpQ8:%fqQ!as4=,8q0k\w*1=dVb<5E-j=ia9{L>K2A]>3eZ16I!>KxzLS7si6nuu$IlXYyXe!4)eS9[m0_.T{	JloMBK6{.
V&Q3uG1MXT>xl,8}lq. r7LT$\nNG,%ZilMC37~il1NWvNmr$B5=X}n_>U,[Y4W%?82Ry~b[I}?87~M7?=n\3bn(KVJA^a;U<Q% 9Mo~Iz`w'iH][<v!@^YN\yb1qvk#qqf|~sSIPX]"@~M^iS<#.d6>3l/Y"`OG~.rlFg<[	YmH\1Y4ZL7H\TN|;?rUY(M"<)?E xJj2|=2jk@[Bt<!);kG2aLTC>v6faah,/x/3HfTz`o=!ac+/z}5"u$Qd\f}{>}F-^?g/y_c;i<o5mm#c#JErg5!1Iur!Ee2(jK(`H&l/ ;>9WP-Ls3
xHr|K]63'VOwy*IB0-=Awy`bwYJIZ#m+ 1X+d_(f:|<@G+@W?mU%'$2#(!xtck|b5/,el/!B|,=0)X?sE/0&g/[3_
V6[jyRiXr80_hDN1x ()PGi^rL%qy'C9:CQu#A}OUgXl'f~kH7@z&>VD_zB,0Jf=8NS18PK"cTM2\|R:DVYf`O[].zm*d {<fj?):dFZ`5WUvc_To(qDIfbjd=yRMO&3o{2b'aLG5u>KJ@Z'L&:zjd 3*n]eAkDfp!wG:*!!;'6~|s=WZ|0J!G:Pt e!R580Q8af>M.muc,b0Q&se4A/N$0 qt?cfcW&@_^-U4aPa
MntD =TuFb[K{@8;K9}iCH[}4:F(@Pqw0=t06.`**DB,r+20JljJcZSa}>jn_ha0[,R7[^[H4kdw>YL"fcN]CK7\<yU4W~hOrPk2X0=!o}D.<dL#K w.\bd1	eozhCvekE.b'ZR	^61mS*Sx=kg73La"Fd[QT{UbM=o6/6SntM%e.2!V-P^'-bA0.+v!Ba,ZjlF8;J\9P8ERli_JJ@NE(hg-%<O6+_ePXt{oh-#O,!_idmd<IcL5=&(Z	>(ph1l0AxmvSl)eLzES_dn8<[:Diw{"M*VTM,*&##aMZS:~%q5C_]'lO	mXzOM]	Zqg#4 c@[$g]80<Y#m'q5DZj\[XQK,d	(u3!a-;dO1Bl@9I;p"fl#[ZRg_G#D)VZg"0q!X!y>8S t=$y^	L]<y%yn	|[Sc@k:j'qP}'j{@&AEzyu|15M+udZBptT;;[x,pX)=QjBi`lG1<BZ!\X
Cc"Bmpl ,woA)W 7Z}tj\{R9jg8i=c3=;Z;KcjHZ4l5*DCjgb=|_]"<y5Br
vxy-<HYy})KiRp#* xZ`ileh^>[Ck!^tM=xjH#|lo9~en*rRb(I!azR:%ed<WbZ;kcClY2@znA0KI|nXWj.=84vhes-<Fc92~%L_nr(*]6[Yw;oAQf5m@0+4` :8cz>CaaHnJ7crx7GxqX jrEjJ3L(u:k=xonKA
7T~h	L#=52;{O	{ZPm+5>rplcJ%j}->`t3'*P3}^5F;zjv]&^)ktgnB`K9$0R(y#jbeRhl=CPmaYStl|AT""4PnI,[>:c`bJv kJ)T3bqwH [,lIo[sYP<!^08qJ8. =BV'j<HROGa8AhGmOF$!2[sOPh !+j_0BoJ<9/6|u_L+1_[F@yXHk_`H,Xg9g;}T}zD35-z^?fcw902lw}K)"UDQhLm3</cq[!vrto#PFLAm2*})5&km^.2NS?9DLT3gF$^6edID;`/^Sa)<W_Xu"=N8jK3{L{5?pO(b7}{\qLT)CP-l:U8(/``nzedU;PP%/jn5g*Oj>}?(oDi{1{	!nUX2/9n6j*zc1jDARX(<!(HS{h1lnUAR9Ftlq%cxr	U4u}wEUwS?/Y7fIOY_|U}cV\Q:lWruH"ix0r>lTR:zndhe	#CS_[,wB/E3M6?/o=2xY.jr?_%"V+YDQ2ot*xQ
OU{?7F!#JkwL,=mYLRi<*lo(>rv|2$oDU8DX|?57>bf83b<ZF\_o'ttNs?z~hd#KDf?AeDv>BMq3P'
4QX]rZRrf=Fo.G<Edz&J>Grotb]AJ!"`#-5]01kVc_E-q@I0nJ}j/bTd$LO9d0c.Shllwblmf26KYY3j2>mNX$P>k&*1}k5$'Bd+`p-#%BM0C$2I+G?5?wX}:":9y|zXrQZ@ez~@<FBs4)NatIip4@dE34$:p-[r.}#Q)=(U`HN
+.^4L|i9Y;Hsf|wWc9#tH(c4yY.Egb*e>TZ"U4)/2s3T&6F6^kPmorX;/rxR) LBO2Gv2<I?3"jmkF04fR%kHKnql3DOtxq-;`}&VK'>PZ`c"P}>YT#9pe[,5HYFZ3=D=	p* 1MdUrH[xxJ*MDvAx/I-YqTP]tG3HS(z0.m7W_,\TM?e1WvN@G=]U'25r{r<Rhy7f[VeYBB{zGW%nU@dYb&' +b"kul,e8>^+UD}2o+7]6C<D /3I4Kaw<v;n#v*
b%-zWg\NWn#ErB>eFo|aF]h\ {[:EN*G@c91rNBtoeK-434Atz2cek*nt!ny4m 3`V}g	!6'~~uq9+ZB7OH	=
f0m}
=ZIjbH&CR4`!D9!)Avpi9@#hJGSvVj"	YV,%	ZZ=2]s29Xa.oZ:=x'7#m-O^$i{+$En	(Q3fuQ;y$e5M
oC@C1I$XRi8-E/,4r.B0AC+I$q]q:&D,u+_s[c[Xvo^`0`SN<*i'9V4e>+*;{LWBGGF#P| 8b3uFs7RK0"[EnmN*,C.Ap#U,''Pk75"Ztkt"i)Gy7
%bRae%.2a~#q"]VatrJU"8@@p9*de7J;F!xw46bzj@wxR&PeuqAEj@gVGr*/`Z*]L0h&7lWl#	0OO c}X1^@4 i~]vJpsq
d:5mSZ[^6e'>)<CkqUo9L$Br7 :z^_[<*MV<AHVS:\H?EMd1S|ID~9;{e7iz&OcIpijhN|LqMZy=x&Y;rvi1WQCql@[`8oa{]xc1b\Z:2HxeVd{3s&Ay?]UO'{!^mQ5qp c[#`00CEh_Y)B9l(H3M~Na?M'1jwribzl:5}mlRqAm.f]+==MXtQ$| 'Ew1jDcf!u*Bg'76_WJJtvaZ4^2~A\gJ Uv3fD&zk2J'[?3
l4T
yDbaxIc:g
$Xi}'kE1SKrDC7-qI 7|N3Y5Es(
L4Gl7Cp	CgtjL-hKs	Ss}!g1u6SKF?$dSq^i8%/<11"Mq4~fOR^pU/@N30(5o?KG-fnggZV,%Y[kS
}/-'Tx!yaD=KV'r<!xPo9zypT)kuW;8)V=9K3J3/2Ss`-*S+xYe!x`L3M6%A*;	33u jD=`;Sf~rIZGe>hF}{N~Dtm;24QM*FoA<,eg=H0B]wv.dpu%Y(p+_M
0NrsH@R&0aO;k@Lwf_Ag9r`'ZVJaQ4rW\/@sHj!+tqN!/zdOX%FrZ#Zghu
KzmKkAtQ!'@N"y:rr]n;>xN)5'6`gpif]EDcW(Gpb4ZyH@eAO!	Hi_P63Tt@<nnETcVY2
n;Q9Pp]eyarOuQEK5g]Y0-yD*Q`=' D*#i8Pcsd`x03nu\=xY7St2uZVeK} E?7`qR8C([BU?Z"|0xJ=DX8_$lzj'>+$;(NaM%BdtjU!]r+FB1f{n{]rF}(qvLG2zBBW$Uzr(S9J^jQ*!({!  C!['h/vz+0sq
OH=KU!{w2) iJ54+[i]zo)j2?K1(X=ibBr"r/&
dxTLl	<}hoOpd\ffX{j4/.2iW\z	9jvce1R$,hA00r*>)0Yj6PN*@TLQ@k6med,xKeQ7?yqtGr%?1"/"CC!a39Xqi|IoNA%hK|J=4zz$`Q@XC:>/i_lk@1*j +A:	%|PDW6I5|wXZJ}6f6GcSHH{l"3pVI5t6W?-=v7#^/v7pV"79K8/o%s}
Zjhbj
fW2KqytBX/!aPp?3tDG^x!#(NCU.79mypBj[:aoUBn sD{tdom"Nj0/^plO>%"t3K^8Fr8C_LGcN0b;fYXM_Q@E`5t/*TqgqszW(X><!4&=z1#_}>l!v@@GC/,\X*sQWg@jO\Ob(g>+tuXH4*6dJ(Yk:eD:5cFKnX9/lW-#(I?kF1Kj_ug?~("#N\MQC>IL$2IP	4W$yNdVfs}^9.g1*}Qj<Q<hLuEVy^2pu,zQtsUS?\`\RugOOC={Ln2l.f`Tzx2RXfH/k)4_	>G7xKx.@;SP (U_ lC|qJ>yre9X7vT_ni A3Fvockkh
GZDh*J(>_0?GXXMK:s0Ey7Tc5  ][AQ}:EksDifyK)+I0@L.u70KWEq\+UNJ AI~R
68~eYbq:\<mC'kai]9pAQpt6IS%,>:52Ueb9)+=sOT\yH7].
aKeH.)+8?Xi..R!_%IfDS#y!{z_9MXR0>U.<U=L-uq?c^8$(SJJI0IZ~U8$*>{w4c3wLdF44?VUco4_B=L'V1v]R2]Lqhs:@6zKySU#	\f<N1D<:w2rKqEPfy1:Q'O:GG6NU~^kP5j2nn&K<@OZX9V?fw]-?5c1hQZ |}sc.rL8$3/WG9ie\H(MWt1ZK;jb}|JXd91NfHN+i}kvH?zArj-&Mndlof<Zq0Ut	v4w2^9Q}}zGc/_'B>trX?:Nk4!xcl1,_"e&"CXu.8+n+Z8#6ojL`l<za9^/&{%/XUGCb2*fam?QDRk]$U\`hO#XA|zfF0j`324wE4Ei`b7qsH
(uf<`/EX3}5O7'?1;7m4}W+`Z:jVPSk|Y^OUrTL$*|xj!S;:eH7L\,cVUx],Jx:_ue*{FCaRm"2<&zi;j;K>dM(a@Wl5UaWSUhw@{"*X:i7o8)OA;{7EhWDdI4_Yx[{=nR~z	Y{`g]8Vsmo:L)z$gn`A33Dek<a(~\%(^c\2Vg<6^6qC8hN0P]{s6p!n<^j5Z->R{X<<Vmg4300q"RRg9&o^"&s KB?#f7Wy3mo^ux`P+Z~H(l'~5g`oO}coV/6HdVePV]v0(LZOHf~?z04#y:+T(w,aw-*L59dWL/jyr	! Mp|Dy.a,P?}leeiw7^nm:p!6 yf-NO5^zvsJ"'mRK#?q1gh0#.,/HIZj2|oMGc+`alcKL}JmtD?i@_1Gr'R3m)"QD?mKdnFi=~H)OeMW]j"I9Sy[< 	W+4!map[R;OQ'.vufggv:tKr5F)e[]@go,&'<TP#\O:q?U&/+l*{A+}sG+rfl42$dz?.ss]!ll+, Q
!zL{x^A
a!@|Fm\QjBvT@c$i_p!^)*aGVJS= W2fV_S2wJZBlNt{gXAt'j3+(s,-f|z^5:1FHX>vjgc}Eok?KMWS<sdi9\"7jHB/<1"V-c3<}0w@I(6<^RM9QXTT<9yL=!8Of%:i3Pc8!GP^`8N2dHQ

ZN\\AFXynj]XdsEEcMS]W1Ar5zI^bDB#Yy{dND>B!|z9A3o&IC9t;16|LP3U_2UPQB?	@Z<z?H	T:^+l]O}2M6bYa#9}aDGt`4g3{HpN}0	lJ.CxShw\N
Ua/_XC6iM,x]ub5`sVS-\z2+*c[e-%:8u]MC'==wio`I'#w"wzC9r9-u5;8+H3\:)<av8)$UVb@LZVZ:<L2|Hi?'V|(\i'FtuW]Qp@&Qo\Tz$rw v_q_zNy,jD=HPGZk6]<|
#jl?[c?)=MM`U2b{X:l`I<Uo;9!n}LVX}aqr5#qG,GJ&1>lf{;;ck%nlq]zT`@0iOp5pThE"CT4C6J>)@.D(RBwVtYTJIJVV#5Ajnm5YMa=!R*RGv-9Ae<JJ0vRTVJH=TO*^jJ7m:YI0,hd\_[B0p	tl\rKdV\EwIzUZ[0Ps$m/b2ddQ<jUy*{!6kOIydvI5z-K5).TMQJ	qCQFd>?&<s-:IJREzyCa6Yu>Ww>0k\"A'pZ&eWSFT(!!	|nAP|REIIr+qG]a\]aIT}JOH2%b5}/+Zm6]~=45
!)C0hE,9{<[dT"0~XVYr<ut[:P<3vz_$kwK&t
]77,0*qF};s
,@>kzo[CS',8?6>=7^r,2+Z"6uI[V	pe?hHS
')Q1
u-y@#`n4"d}VQ,S+X<S=o}3,^LeF"QWW:`=2;7qyYYj>o=5N_y"xYI*ni.T!d-[p4.O<2RZ+-bUXCbFp?1QZmW	R2zy/bX CT7{96-k.+/q\?-YE[n8Lgm?fFO.GCSR3T||PCaM%JW%]*TWtbJS=~a4kPShVo|A*\Y=B|n(fG`qwC7MS]2xNh/ux3h%Tf\O55`q:]tuQ4A*!Rv T&SQjC4I*qZ,NeH^3q9gVNFd:(g\&p\JjUY=HbMA:ytv@4@7bux/_ylEH{PXB+Y8)_Lyz:Ct_1CVguPhKWr>Hbd*QiKCi<;|VE8{Krt<)rD-U,#- !tSyj~i.Q.uh9O DgYZ{-;NYV.eyHy	\#F^_r(U`br[s
-o?T=dT<[L-x`Gge'q}Ng"zu2EzDgFz8750!5fCDyucI=O8}]]<Q'BauuqXRTK%Ogcpti+f&\Yjj"*[:OW4H|q-g9('jJ5m:JeNq-?q+zXu>7q3Xc]p<RSzt9[-iv ok]LRVo{.aqEcD	=F<*-M+GQdO`Mng`4AZ&KIUZ6F2Lu-Z(#gbLomD,vBgw:+fE7f:~
]a(xg?.	r"{r._0DYXCgW|9H(YVX%D%{FE5GD)L?"60M
Zz!^(ykx=-)]#.:	zU*(-vnAfZkDKQ2S8/Wd}]u3TT#XNpY,vBJOtz*v_3DL,_)]tBe6ER~)*o>>J5j6-?	I;C[rg!kaL1W/IlM{:Tw,qhJ_f?;@.&W<>C.sAY1Ka[`d.F%Qfg$k`m!uuP|lMYq<=\ d[yD{iLyU9k.<(_Pwm&Yp\29|=#D.z*+8y%Ig}s	BAawcZ0%I@{8ocHzNQ@43m0;U{FPNA"v^w<)#ixK)BNkT!PjtODRfq_5N[WN#2_Vr|-5|~ygKwhrD<}VQ/[B5KGZiFT-D-jM`!M(A;\G|V!]JaZLy{\&m}=l;]	3WEn@N)Rz0sq4:Kv45B^MJxi(Zr}HT!#mHSy9EU\f^{`BU
pYyz29i"KZeB$uWjnr`Bi3o=]y;,~ul`!-}g+K4x!*:ja'BZ8_w:B`xhpkH<EX;:6u"y_Wvb3
/|.<`I%[V]rEdxMVeb",g\_'I(de!q8B	!MtrMEAK\9.|{;8aG447+dD8
I8~L)1*wckp&|LoJ'8/./.W.a54,,Fh	yb_TF1;Ju~Ss1cK#C<D~I})=c?7G~lPTjs^
l"0yVsGo
;dzAz%':paM$12Lt@NVaVjb|*w16Q"<G1\*j_}5*@n8@-YI|{h|9q 4w8Xs!s_dET/u2%w2mAcMFB&q]<cw#-_@WxMP&|i3w]USQO_JD:p0WD:_}) $WfgkV%5,c1_9\OfF;sbGBJ
v<!oN`\g|<vvLxiFY}*)T).\h`I[Xuqvu;Tn&9PB\K,X+\H0`5M,0U[_gX
{0M99Eff"PRf0"i\vpbIK}SdL_Er\-u|uzI'&	kCKH^@J5v0hkuiOSsjQBzVSbxo!Ni`t2sN)SF@"h/W+e=vM@ Z9zu2Cl(ZNi`T	FJ*q3eBXfBN#I/Y7Rn$o|teoC)r|uwatQ$%m}Bm~v_baq'yt%DNTc\ jBp.].(W5Sd*4j T}@|l^B2$on;NrTZ9!+`%vd;o!FceM<-6+H/rhlHZA/*PEV5@:<.O6&Vcf{SYP-*O-.JVnQ&h':R,{p%*KZ8[9(kv]Va*(E%<wBc*>lju(sg/rLnrA9d8pD)Q`qc0Jr H@.<JNAony]mj4#m}_,TRJ1J6C	y|ZXw>32 
JD^ohHQ$98>x\)D,>5AK,5#4Q.|j)R3JX*R^;wMT37jIoX,i[6DdHAht_h>>Le7\MGsQp"A%DNg/6@oM``w'b9/KrqABoh% VKy5eR'S'FPe^Xl;t(1?@!r{z7<k.t;= D6% 4=-SY!9q&VzOB$	8-*QbTC:XrAq:@0*$!f<Pf#.9.1\n|-6NQW(
yp"l5r#D<9/ vzkV
%KVXchlyrqyCV.I3n{9*e!G#)s|.ZCEl9Z?a|O~Z4D|WZk49:nsy33vas5uuzf(/6@QVbCKN.OZCa68XcbvH|LJZlT	rJI`7w4qm6/5<:H=vM=Z'\oN'1"Wvk:z(JTThTGe!4?>^NV6}c@jIb2f@b.Y6%1(@Wd]U5=$Id\f]Y6-=j+M?nH*@wre6oIW<z4d9Q/{#0x6*,R<oKA>&cO24b0eOq^1o16s|	.K!UQk%C-8\w@b@)<<8"y_yR'b_Y{;^3?V{jqE*N5XxY5ooQ'a|"vdLA{kIIt(P	N*qRJ}8^YOfG_*N&^BIv s+$i DS/1SZl/VnImHq\Q{<[9{Vq_2CE$OX5`= oTxsnD$k0QD)mE'K]Qn:?t#T7YZLd:M}K.=Goy8U
;X0I;7]^g5"r1I9kZLUR!X833C e\')J"]pb3ZHLNxYm@!EzTCMWX(|kYP=gL7USz_^ckr'_WhmjIc}?*2-0khyM(U:tn9/xaFeejcijwzw~aNomDv4X""42LbN-=v^30\c-IuL`;J&uF'	
k)Zd%F<ykNCNRAGePDx0l-n5k|ZP]dB)cEW72Pm!OBMlm8l_)?6p~0\Orn"9i8u|DGoQd?f#Ms69@ APO<!c0NUsYJZk$qovnU5'^
]lZ3X>YJ8k1Z"X?z{:1[X.i:M_kJN6D=O^uGxNI\fcvU~,6vPhmrRS!p4gL&x_+So|GHaT3*VG^^'#[Is.TNpH./Iq42kSIHLmxJ3nTDcFv~yaLQVwPAQ|zbAD0v,/oE:G`;BwZSB?{]rX`-^f^=<1ea>*S@d	vIC]i	+sPMg$+`02I9@~_um]OxUxd+zOOTu4\)&'t.cg-c,kYS*}%!kZTo6tp!KR'h&%H:1$p!;0NDkHsJ:>2Jj^gaY.N'"> [ kcr2[ 4E9FV${,8tCMMpr&6([-{De.:QdidCS^3X/"l@ LoEt
zjlf_Hr29S>Iw55}55F4"-8 J h+1h}jucUYX:Lq45 `^OXnWx3T*O E}.DRccI<|(iF5M	Q-T`ai93&uaFf!Vi[oM66m{{m\?1/|UTJc8V$vCyj&4^\!256.k'@(o+V=%@\cc3s5e&Er+@m;Ku?^LBSYc
mv@n\c]?o>H.9C%n'yWZ7=r,pF'ry'!1a\t\=Z5R^Sq#Pu'u2job29u`Wgr'<97%+bYw<
-p:19du[X7ze2.eO8:|F7q)[,#Fs=N$<CZS+
2	vc"C(G%v0!~WA/3_%R)L+S-#=AjK/0tGY/z3qX0kXwnVM{OMv`.<-si}9}G;N&f*_G6rC02L'5A_j*~(QZ*Z_ZI{C(?d?{%^xVtNrVE@t_WAkDHm$b!3*TBxx0WN{U&@tnrn/L<%mlu'@y#ZeZFVIu+?`opc5@ {*$~3!5Jx)|O0	(iJVk`Y{RU}laY`pgL
Kq/q%)_o*0@LD5gKR;V'EJ{Hr)#c=7:oCj7RD^{co@f wmC:aoYGi4&}uh{7rPeQUa%Ps;'j:itd0JmTlgo*/3Y*b4U?f3qe8'XFHXh+c)rPZ6$ @B.)>eX	kFVcI/:Wo`HczqImr/NUDVhuL*SA'8s>?m$>T;Vyzy6.ecWNKzc'!)e#y(v53~!3?.D);y:$u:84pT^5(z_O$x +SCFfl"(#T'-CCCk>fcK&#tl4k@xj5C,PI*S&Uw'
W45B3kH"Ie.]WD 2WfZ(n,@-+K`wW<5yt5Ngnfm_8LI}LqLe(`yXa%_F
}.d-"SZjBF[+H"~(Yzdg;A>[+lX_0-!fL]O	3|:cp--;[`uy*jLJ.!*{< .Q{c92BD{ K.YA~NfIi[;eL9~L3l.`I%Gs#AL2.B!?SutinXPP|0|GU)4	0q-SZ)?lOJZ<Krn@"|j{|*V?N[c4]J+emXSU+M8/)JT\;/t6,
4,;f#z3vx<#(]!0EPg`qovE/Mn0\q #|)~	ljnY)<=+8OP^_+
O/\SKSpT;o6-}oO),$z#x)ycw,8K\u2K1WQ &|BNMJ=B{$HE[>E(<M
(_`e`7o#_tq\[s;9fgR)sJ,JaIH+iLf%H+Jp7Ss)9XX]<}rJEbsmWT7SiUeoi3z 4JVL|%]^\b}\	O$EexN]E?6\ CMDvgEAnT,?.*u@kl?vx'dk=:U<&-6\.+F{
2$`xW21|O&duVQ(vU+x;ETK.lAH!9o@>jxw{|NH%-_aOh%k$mR#D^9AeczB`yxueg/<lwxu=4"QKf+yK6m-oB*['gc<KYgH*9Aw;ggMd6f7*:gVVDez#C];Lli},<(nc^$^zm$A}EuIqap=gX^x`EbU!kiwwd'cH)=IqA{'oWa%[J^q`aZ8DL6XR_d|HG<*\@9H|}v.o#&kUNT	s-M@l!CJ; 4rb!eMinyVw<c+DD aQlvgdD6yM~OfQ wst8#hT%DOj}UoH(8cm.mEpt*`"T.,9Y
CLbB{9qYoD%%d0"}TgkZs9 gZ/=KE1-c^M|C2tO-A/|4{D
]aUrt'9J.;cnB	
W8hW8GE/3$V%AJ8)Sp}^D^b?s6ah.}@3YYp;VuvDwfSzLas<N%E(aTiv0
sDe:3\^5vS(o(y-.S10b`([?2<Ey09qbvE>
9=xFVf_87*rr9NW{Rpi;KEFMY01et_'5$
6EL{i9*x4;lia-,"Zv'-.Mfu:1.~|5gOwzrVXLZuCznjB_D3hJ?G)!h[DQM"mJ|gt,A8]I@4_C'rc"=vCHS~cW;qNcNzx-;a>7TCGQ73uTsDLG
G_Mg-3rgy%jS/wMv@
V(^}Y5~N^d=tJ88DZ9L^p</p|&N7p4;gNvsGYE=PbKG-~Usri:aJrY2:6'$U%XN[F-'LX$Z0n_=hLZO+oPy#Q.xIO{h9{m?02NSx?b~,xt!O*D5/W=lQTH^'<VVOAW,{lsCv}1:[j;Ozw2UhF(Mt7F!~F1J~e|buHuhy+oK)Tj?rp@.&C0OK5N4l]arrr=%6.,4: 7'iozbb3#datR
a_>[9}$k{yokZ|M2H"F|zFuI@|qs<O6Xh[o~a!eH90c?^,w1q=T0D%a2EZD
-t2HSQ4/5)C IP1 hlt@mH_)\G|u`Ya=<Wm)y3!	Ad2l(M+-$)0\	h,F$G!U>}7"(-D{?fcfXM"-"@,>W/bdH4aOT]U)B)g:<QB~6q~693B+i]7tL,(}1`I=HW&~O?TcxNA&}rG1pH	'(@t5)Bc;MF{nFgx$*Um>|?ozstVzi}f'Dg')&j*mnHfDS)g05kc!2^hW@k8~"qav]#AC6p?nnKjV)<9.o5Ci&BMU:iIhO#'G
@(l65qF0M~>][-V6b@< '3q;>2ysK-Emc%Xzbq
@Tusavz9t#x!o*(k=M[2#|jj-F/!?.`#kjE_B0K.S=9j<.Mz1c0{t		nS-Eb!Y=QJ oKP1}Ty,3KAFr[!qgg/\uw!F_'{M<W7>in+c~|=+*0u)#JmIB{D2&]|P=i}^hTfmn[7kM^o9D	}lNNLR.`M@-$E+[]@cmZ
B#|=Okdw=l~OT8^4UJhq8dPNh CRpt}o5qKw SiX:!v)cWg,j$>cZYvJ{ =klFXWbI(1>cr=Cz`{2>Z]h='k*Sv@&D+x^^bTi[4p2:u>$=4wc]"Qyw*`}]y'njcPU_7w7uqxw]vP.#Y!7{<7YdH
2c9"o7kS	@Pk$&EEm9Jp_K9zk@*f!!qq>WX\?v36QLV(F+Wt#Sy~GDW:eMh5?2b.~8FGU%sg6P=7fxLXsGaIb*=L4DF9mo,leT89z8VJJ/%B-3/aTSu!4oXA?TOkzx}qVp>h*a=^<$sJ3M!mn#\\HBa=dMQ*G8y_/\M'Y, {[C2bUqw<1HwyJ`\g/TkjgorjW:'C.]uMFs0&a!}^Wn"C[o8$bc0Guu.1mliSFG7sHr4
zm\%Iq/cXG"OO"NIk}@TOg$^R%nT(s<^/'"zq?-ZKF:whHza{g{(!7WnvKa^7r,!'NS-;,Bs2@{RN%w
}$ITGLF9d+2VI,	u%jsZ{hu)%Dr6?+}Q1l*{.Oe")<mhk2WJz
U_*o'J+).xUjV)@)B[^k,_gkKdV6a00EN\&HSV~@{RJG:RY)WXa8|!}eBBc~N8JiBDfg#2LNs%*>O.>`FpdZcG*zJK2Ca`h/R~/Kw?FnC+np<):Sb:*-@AI3Z>jP*pP:U4#nt{5^Iq>D\iEX.{46#k6>g?g=:\._XIDQLODE73 n)UvKGuWZgf]#W1f-I)Pq"wtUb;PvVv&mWAh5$fw|&>_vjX}5N{(E#!JbLO6(fFKgzE;@Zf$t#tBO+`m5Op`TY[=H9aE52;pUDVu"SG$lIK00z.E|yC `KD+h]0R1r@H(]Dy[),!.*+(n>z96@_1lz;l:VT%tQnDKerk7E:E|s_q,(r+E04#i?P.KUe\tZ:u`^wbSCd';D$h(fM'h_srKG
	sp-kF(zXWrWKqROQh,@=~mo\N~%=|k>L*C*WeJTWOY\<N
)N@eY;-n62nWN{B}`d.1pB$!?[X$mv/5ju]]|++a\z ;
@E)H0}Tl]wS^q"d\9 w
ex}o{9tsDCJ?<#MYElB;Eu) @o34?
d7ae&hezTc^msvgf`681`@G5Os2$0z/W!u-Xf!bH_/sO'fg!Rm0F+g$WdV,YiOWMDl2e0-Q_Pt{G?
X&~p$	2n,A|e6HTLhQ(\#,?b')z,k^".&lVkVwQv{;9`!dZ\ (E.$-pD; YFT<s^Oxp+.Nikh2O5$0j7G>"*BAbL^Iy{FeM?v1\VI!c,Jk@>K-ZE6T4<*guIMTAzL)W+X\bgX|w*;VKZH39!I1l9K7{
0x8CqP_M5_cK#"<!qux)QlcuEtCQJKh#~Zuv%g.Vu&Yvmle{*?'8.sBwNZtD[I#Fc8#gQZK-%0&EzqQJw,DSEXP}djvl	D.PdH}?T$UHhdn\j,X'=JZy]k%w[@|3fkR]|/x!VZy1K/?Ci{|&Q&d.bTvU![93OOVSE&n\%)7=E"
9REqd0fSu0Ro3u>|_u(bz@IYG0]c +:[h3HN@JzMMZ$zci}Ie|j$Cn@z!h]mS8smkS n$0W-|j_do1&[DUyMIJ0TsV"B!MbJ	-7mc'`\N(.=zP[56(J)[vBsDb[G)MZhD2{D3 ZVEmJ1Xe4U+2J75({hv<iOxvCL]=)qYa/V{$;\9#vJUwC(O' jeiA|jR(Nv4Q9qw,R,Ve1
zpP@t9h""HXScRo77nO-QhcvC^JY;gDd$76-zNv5]Q`O>Z`5gC@g^<-ew_1f63$#9`ficMW`ybQG6;Xy]XN?e]Cwe $-:>~;lt	XGq,d<FQ4HmC${"n/@<;1snN^SyC&(_CH'xn:.-_<<)818(AL]RU^Ka5wyDb#rl+qVA9@:@_u.l
*V9g=_t"_/5`8htpd9FY4/y] qv\,p5r?JDmQ!'N5<SI"idX+=6oAY)(P\"TOrv8W4f_
')_Lo:wuB/rU$6P?q9h}v)KIctK~+W[T|q?;&FJ;m3U~-jF*Bk*(*
"<szyhb" #*wnZI}#."|ct}yER)ME/p>18_vS0DK=qG+d3"|;<tfBsV0xoGUq??O$uD#^6}G\?J+n!#f14z;GC4cI(NY>x$j)4q+`2k?&+]
$4.A`<xL;g-[:*f7l?4";^/5aQ|E.Zy%+;{vkVu'X9OLoA!2WtSmwP	ybLA/$vl-q<F//x>bt;{?~TE#G1y
1OY)z}L`QVP|XA{x<8Och?7U%i'g(;%yxMvVmlU|P,k#C@	BBIhT.#|
.TtcLS3|\IxU4U`	zYK#>R{ Xc
ap-_e@GDFAP]7d3gM)nG4\j]&+jtL=/=+]B'unV%%[4.XBq/N0|#deGA7#VMx=H-4RV%>c-JlS?i)4!#@mKcL|N!nc}0'60h>:.P
RXojuR.@<DS?OTrcmWEL^YFQU!{H`*J	~t&aObpX#}	?lxF &j@v)3cpR(Ovtx=\b$K>kb[/TOO)t~|+Dc`w|j8GyG0qM*b	7@UhQO^g4z\[~&[=}>'sG]mr=tA{5CyWV&s+KiV/XE(|aqk??j1'=
pc;b.&R#,puk^)z&$W+2e"0FfxzAYz1X"E\pldFDatT&W*Gq81m&O>X_6D>I=c's8N:`4TM;^s+d[mqvbPxEfE?mA,SSNgPGq7'*!.h0N
t7MctCszIA$Fw^avDK4,-.ek~N53w{~
yMZ!xrEhge5@*;xdnN'tig}ae`K%b@mQn)&F=OOb?eD
{p_iclsMo|{9(S$'ks,$ju\"WWgSTV4=pTbH3TrY9`9Fz	pSQ,A;"k(0U[9"KDMIugU&M;v=?KpcPy4u'b\;ky4_"*~1UaJh(ZXj6&ixu@ql%2ZXLelb
*.1&%?(5!y*sH&G=^XP@Q Udq*AaFiByq4~4S_xvL^%Rs\hU2E"(-/{x hBa!RJt7FCOts_tO'5h 6El;:<&R!p"N@TvXe!,eP-vlF[TO}(/,*=/n1-G1iNho+>MzEr8R?c=&V~mZS&p5r&ZSpTz=n]#/.8Em[_'X9Qv5^yf25y'kcsFe[.{x|~DbS	{:9"bWgsaeup?fE@b
?FY.96c1[)BU8g&h!6S~br!U&x'5qsp/O+e+HAw{SPDbZEJQi7/V?1u50@/$Yy!FPMFn4rh.;+W^z9oX(`M]QWOvW=,vKl?W*W'zM	Fs1XHMrl\\ 30b9Sq)jh%cr#+6HYC86caDWcAAua1l0q|94X_l_TDY4yGTe8_@_'L#)&R-%,|:Cy@T
_([7:4)Ce'^b-h_=S\9%p?XD<Q,=*(9'\AW|E;P7Ub5F Wb11sz?X):@j+*cVh\z&S(9<eEhKi2'pPtj!/UoWG>UjfixV7C|@2owgsVZ)zuY!WX!G1DI9V	+	J*Z]B{lR[xzQSxEDPFC$nGS[FfjO&En
|gCUC7-D'aql}.cWF,JiS;pwzY|Wp1CR_x&=@:"TpBWY87!V;u+4_5uP+MK9f`kKBKw6uzDCL181 G7B6#*|v3qck{J(u9"736,y4El1A.lUZNc0]$!-c"hs>Y4wgsEsEfLub1m=|1e4]Ld`3["G@!}6`P!Z<}L3=4yE#%t3N"u]3__wp&16\H|tJK9$}w{Aem>6L_\*HX9xj6ic/jww;>fl&=,AJ9g?TAAnb#L!h=Q,C$UNfe%fQ;A5.yRUMtc:rf#.Y(l+Q|(`F.Sf|22\u13BKEP:B63(Dc2}k,&/	n=36=k6I&1#<x-Mm 1/ZZU)^=a6}G.JqF|GQ:\59<s/U\E-*K"mE.PN81BU#aN+'V^:5X\4Zp(uo\re)s&XUjN~0P[Yvip$;?9f!<trHGKwGY)7U-xnQ=^}X}eA<9!~MD`c}Fq`g2s,;L_b|-~zkp]i7#bec6T8k^*w}>G_(R?g/^a>6xn=>zEWCI]=Y
7G|'R)|}Z2PpmT7FFMd]g_C]G<PH({Hb&3Y5lQ`;!N2fdjO-B'[>N3{smy%v|V*"b< cw5UNv6H|_&Z|O&}S4_'cbX,|=,U
48D_Wd=Cyk`cwtaa=+O6]v8us7*
lwq(>7[w.az]Tgv*2K9swXrIP]PfGwOOH,ts1&e<PTNN_+GbsK}bLY-9hOzR:oOWE2:-0
{`T,fgVg?
Q!:RF/u]9`pu+a'k9L[Olzew{<f0F%fO#AB}/8^PlguH]Vk'--eZs&nry^W%6~Y"9adj*)Y<T T7TSQ.Qjdn) :.BG::M6v/3v#vGu]!P.o=Y7[]T\};yn P2=I^i~SMc1q@G<>lZ	1""g/{=/6Q7{%ydcxhY.	&*db=6%R\0WxC
tU5zLj6NK-TV"O#qElEMl\<7FfwvhjP(J5@1QXa;+gtuAso"Ll|^d~*_]yPur 0;/V0}^ju3"7L%-`vjJ#sU'tO<j[s^ivLE>7(_-Vv(nYUn":"dU][SHs1\Ow-rh=Z-y;X+F*ZO\G]psPOVS*f4VbXl
IuMZ
?I]aFCwe~r]-n(y!uHJzyI|dqk;r2pL[%4o7/V  bHPV\'.@	%Dxyv'Z~o WPOMH+LiZyO%3p#?q7Y7],F#w_H83>0K^4\j?qAba:~J~0qFa)
|'xub0K#=]!]a?^lJ*ha6qtR}.(5/KsSa6J=Uv){n_z~Ej_QfK0P@{<DU3l:a6MJa+	o_<>.q+c:p!}W<2HMS@_,\oneak2x`El9zlyZ<-|_N?S#clIS%=YgwqqVO'%;yKp{4!I*@6OD
yen<&~D,"<-(C%{xTl5Ks~HRo|%F59^r0M*:ZP:Hl-4o/ThA<iZ0rg_$*H=<(g3,P90km\X[lL >x\JelNmh{,a"jDcv55H)3YBj_	L|8?6f2l0:qB.aZsD`N|<xEOZ{;r@A^>Yoi2U&@H4hDNhWq{}G'_y:fQ7CG5SV9F\-B\WJH]k,i`_	e5PX5_2-@}lQ})qK<LCyg[O8;:TjD?Z%jq%AO<dwQ;eP{*@q.:7V)>+hys\AYY-Q;`H8{Ji88 rk}N/BlNEdvy	'/R</Pcg7KC	d7|0a=4*m6O.k$u_aQ>Q^%~HQ#OXm[F]\E+Z2;Uk|j+_8jqlJ_AB#{ @X{H14{FvfVx2POWxacde'z8m`7>b;Y;hQ2CBr:Z,/2gY\a6G]Kz*CX(6Gx#w!`CVvQ g^17oF>.kP*A|OldH5facEnZBl`f[D6vVE`=t. ),88[{o?:,,8&w4aHn.BP0G(l,|Ej>gt5`Eg;D8jE+!Cx=$PW!ob2M|sYn:;oX-WH=xg]`iu}L]5i\>T)UT)uQ\l6{%ojeR&:%8+Rh;f(HQfhVn|7*G4\	$Vz{xZCv8DUc*s_%y>	z.'d
\GSn=Z5yWo<8|TGX!+Qx`)*]U@l_kRl<g}{?0,}BbV<0{QVv`7'$pZDpdWG#T?=YVlf9s0)Ux%f
Ld9M%2M!c8Yk_bj#qh[TeD<RKC#v
Q%B*C
;gWMVN[eilUfH0L(0|b#RHtQoI(454
Q}Ny@B&?U$LKoVGXq)B-<{:OQOm"9axWT4<~w3R3-B
	og<fKMr[i|YRcC|-_My#&1
ZMDHNxxkj=CYh+ydVDP97<~=0&qAHlbv7p:EKoHa,@0[E^t;h~}JAyJWLF|+4}2?HLU)+=y=l`HY-@PC<]_Q/0u|j0)UB(	oFDh7'?w_C
R@3*Dm)b}yK(kEG=	BMUvQkz/Kyy_n{]EIunh=(Fjkb 0XF4pJ!EQ:^F{fJ8hXl7,\{pWE4#hkL(G%'Z;BJLS,c;k:NNhLWor6+8"'q}8k\f0wcK\$2	}4#`*r~M{ZC4V)`Z Y"u@ELbt:yD9tKS~Q;xV"<{Eb9LMJ3bk_obG-HJg
Js*b;Z$dy*`-4e q&.Q>SS[j>=e
MV.\5{OA
7,l3()Oh?Yk7z#SH"T`R&f'c
3m%8<1(Jg7D\<Hp&(30+w2HJZOTwaN-nM`J5+V|M-=JW|ZOk2iL*Y(TiHwN|RM4>9}'3$mn~|+M&MP"/<Jq"LKAj)|jW8/kXc/pTM6w]pr\9V8>Y/\o/7RT}W#aT7i9a$1f`^(>mv&JFz#>9hxO+.mnP	xl,{DAawI8p=~*zE:drw (,v^($+(k2<<c	-_(FMV,iEm,_3R;aX1[}v[rpC,k0Yga5UU)vQ,,,Uf'vjLQt 5?FHapu7bW68aJ+r.fDs	l@Qa"-@rS|x1=ezyWkC,$Dnn2 P9P1JilaORx'Gh}%.bL%$o~vRq^x8~]9)J Cm?T10YOQ>*	1*,W'`]Z?N
<pEk/aS5vAaL*$f0#:	FJFkdx	("l}E_dy?@vpfg{UE0"mCa#jjg9Dd9Qs(P,\Q!Zg<&FGY:6*0|`bmZ$Y2fj9D4d m8lt/iox2R?_6UCi1O-mo x{VWZJu4Sz	-Gct@fa2Dj<o([04wF@ECoEN:^lX>rUJS|UB!Yj+*E+eh2{sVq{lu!h}yn9)z'Ck~&:{a@\+k}St_o{L@K!hh4{4$0u6,^l!C*_cn)QA=O-&f;32`Yj4]=6HtM+x__n"\M8syVE52IP+c*xjpR
IrH&w;<2->Vxy7	OU~L'}/Du5|KYN<:3C**?`$lSu+v	Q\M;Va$W$RaoU&+1(15Vm]lW\)6tF%ePlfA$;wr4iqj	&Wv5`byBqI6,zwyjHPF)hu2wYO';^~y
U+z&C<khqJtK |k7!hHHFG/FIi/+gbHQ/.TD
!RE-gJDq\HO{rgu|cr\s{\/YS'Mt&_dR5%"#dPoYJVL4G64[[BfdyIC9WdGyYBO9~AzBSVM(&'ZSmS9?bt](1IJdR>'?O}mXUz": #RTv[p:o}w6poL.AKII@
J}6#.U4,5fITr*g%g6i2ze0yZe3KWXk]G+	>{F
EgfXr1X7fu*c[N'l5	uo1$.q9.'S5@A8'3Zox?}a'@o,phk+=6diG=+o)!]3p7yT%yS]tv~s2u~Q'~Hc)?6~mZckOi0hI)h=eeu9(H>}\$IGWS&j`;l@$8P-4v^}VU )~sFzgMKI$5FE~J[lROnJ{sDCW*A!EGt3!WUI2H*/?z
2>i^!dUwBVB3D</gpR6.%Zw|kx4@g&x]?2Z$EwGJkL	 3vCzn"9)q^,'>0nI}c.O^VN	?d+wgXo|EC0<_0
H"-C{j~o6NC%,St9vBNobCgW2W(k7GHIvbp/O.HmIiJ^O5'Fk&*(F%+pvmU+=e{m-cdx	[Jl;^IWBw|p'1|wD&Ida25Cn36;OqM;cxm$i9M"4T K!P3)bB60s`/wSOse7*t|NyI]3|m;'^c8D'QU&\0r^O8Y^:{2Ym|'OrBgjL5=QVP<<i9Ovf_;Oj;(W|Dj:H~^Ae`Ye	hl:@}q^(ocr,k)rn`,1/|2d|YI!yN:FVf(./Sfz]SnPyo|lZ5=l^on	_}+%U)^7~JSCA<<NLk
kh_lcc.Xiu]qOif~|[<GKRw%qUml%i~x_J6::KMk/xA[ObUB'XJhf0pp5`C@n0P+cDo!|n\EE\TXT;yKgj&^jNDN2q`,Jo+-]p(lGsNa}$SJ,j`(Qm4.?b.onCf)tf<">j\[	O`z)3y2dv)mj8=36JpXh%<R3j]&P6%l\a+0o]PuH>l	!fcXr(w9N~m4JB^>_oS3"h%U+	y16Q,l=S(CvJBo=^h~T.753o*W>IO<-<sRw8zi/-A!8gqsA5jcATsRPC,_
|\HA]n:D/hr3ed-OCs;-*#Se{iPI=KQTL	N>/q]{h&:-r(G[n\53-(0`PvN3.H=\pVQMc7jnjjMBKga2p*~6:tWbEQ_:dXLGY\*]$pokf&`ZI|iCwHxpJcD^zch\oRx1AeoU9[$jz9wa)]u]v	)FEIsIGV_(ERRh2XQ?Q&]BI7)4w9(_H-FrG^%A[>6k$RpTwpkj_
{9{;o3I_')vuYB;pNWh+Rt8t:o]K& nom/66#[S(|k@K(l*IPBBF@R>NY)K6w4|J$1PlG~a=qkdn}(|=f:E?#YLb/yqzs)X[
U{ \gWI XW">$7;jGbG:s,:H{B,	tld^*iB.lqlNg]W_ZgEG6`*O)rcfTqo#Gqe	J}eX#6M@]S%Hn/[y%h*9dV<n*(|,hlG+-g.']
]Md]fM}2i[*06+"c!F\!P+j+y[^;vPmCb3J$s @6+}t/GWU"mUsD]HHKxf9:Pi2#8*+2-a"Q7$*="Foa!4)Q/x1Dp@eC?''I'"7\BtRLU)(*8\s_y!}9 %I}=/tgvw#q!'vC+f1XuI4^_fY YWzNVGUb^.<iPy{ #EO`f.(QRyt;I2?v w!7xr2ZhM-nmCHyHD!~~e^oajJdl
7]ei0\<r69s`wZYU`R>'jMiv7b,M [yyriFvQli"0A\LO.-t*u5~<9	jW2{I+kp*Xl0-+mi#Q4U14*`:Hw}N\J>M&wGU"Guo{IbMsAcWi>eZ",AsX".=x/r` $4S`:T[;MBexP)x'xheio 4U4?>13U5_zr
Y5	H"6Bk>5z8T=\fBa(p21,,poC%g:2$kUC]ZA(Gr_kyjc"mhxLXkL<4|j^/hiYBhNG8D7/N8;I$~>nL	yEu<+btoeE	944ky#WY<lVKd'&8:QZ!>##Bj!$eC=hz55}-z|
[1EpYlyiK1b|}FyJ*tRvjE=tzpmKtNu#\zra8zv%uAT$X2fKrxz=mrzi5j]Gqv1J]'a`=GgSN8?]gWvyqLdyNP1tt,1lxQ~4?_p @:/SN,dJ\vnok'a	V}&NqjkA9<@rQfsU44'Tm)-}-Ac{!=b[z06f.KI_^z]G[AjjSu:I[aHO37T.;{+N&^+W(+072v3:"oQe,Q*}K
SzETd_PVCecEf1|sB;~b2U_ydw {dj+	F=.m`y|\c^VfA7pjrvDrj$v$bKW%@Z	)%20UCz[\:HUf_m_h]9OxI%_gY[oW/0Rc1Mp[OU{sJEF>efMJAJp#,Af6nevRbY~50-zr~{R`}Siz0n`njA]FMD-F
^cGj[5BoW$i%E2D0%&cwRfX:Ae+2(P-z&1G#S>Al/h,IM#`?\o.}3~!41d:rNH"wIEnR>!L<feaY1ar0<=s=	1F( Su/d~[B|v2~js'0F/f`)H#%*ppME= mu?7HJN<cY`C}+\\HnUV}-haL+P@}3] A5BO8dt:c}a[i%J}2'y09o5PLt(%u<l=N.-7ZOT5NJZ#jos:$EV~&[|sj!QJZPF]#+`X^((E'eCPNkT(p,Hp8@C*#Xs\JT[|,[ps3	B:]=8ul%u8+R:hYS2t}D5;wz0B[^Ox}1~))4]>8ARP7#!'-z/2[MO=\`co*qn}LM.dX\J|eiv9HEgO&&w88)K(=%	Z_O]fcW4q"l;.j~E.6CwLP2X4y]nMa8^K]/Y?Ae$Z;[Ev7Ji{"2udBq?8PI;:4ieu	<#K/ aD6E7uxS9	p(\(xZ"S^x,$0'gp8U?g"JJ}[|~,BOXQTV+q>P/[EQn~`NJ$8dPZ$!$t n~u_gQrcX	F@eGL`B~ .'?TwUBY[}Kut~@ gDa!q;5*V'D8U/bD;G5QT[AE,9<Z9O~nQh1wZ8[?%:c^$S7}&j`YPs5.6RL!xWi|p}pChy0\=Zo{W(5XL~|>uMdc)_5[Qi?Zb]CmBHnqEC#X2Q*	{|NW[AF<nU&jgSyQyC.sW_:o%jn]$3/jce_!3zK*?xG}VW9V\71F^S=*R5;m\u2y3
W[lCK10q'.KD"X:Gp,-xv^Fa;y\e$l<m'WwUfm!TCJ8YaJZ+4tdt7H>;/M.DB9eSr`{/t'oYNvUJnQVtU'?6X*Z&eojIr5&8xIh@:oQ upp/3S5Ve~x7"_p?dT1|2_v@*C|+g7aKVIJ}1EbhO&5(7v=Av^7\e*8x(:(=9
 8#.`Zw[Gz?@z01H]r}".UbWIIXWQc
].G'y3?2V4%+"VG|:0r#oY%6Df%6mX?nu%)1]m-C2m[' BGU	`shfGq=L"eH_9RNY,_	)j)zUp?[c<Q<77;l<IN'
=Z=RRygCE-g
j+Cc!o4Sl2@HY9[Fsh*hcpSrSBj`&%gE_Y6r2y3b&r'3UH"%ON^R+)m7y2@(a|H6f,XRv<-?#M(qPKc<UJ%7"TKDnW@p&
SDTn332G0(&}E;
OR,"q3:WmXz6vj	305pX#/?H6KZJp/F|#"ZFi7a\;Vc	Q!.TO-I'w[kpxz!`^/\~{Tbh'eL;FM(|u9ZDS;N2m%WA$ d35UA)cZp1#Yc<.X
Y&+;MItZ;"H["ViM/+&&(WVZsSA$JxZ2@sUb#,r$!7)}wjxKD^x# _o$RF11*t6)A~h#.vMWajMFt
S?Wl
nlX7zn]^?#"mKV_Bu}MFrfG"q><rCy2oZ31c\112F8{/XDV8}^7
q219?U!xYTU$EugG}W/N$]%7 }/U!/B'`j&5Q1;
wR%F(u#ja1$2Qb
B^97/C</MRTnQH?6mE$Th\Cv$)o!
.
<V96x.g&M0_L}>KHlQ:y*)UrkxcL@"'.o%[4U39N]S[lp?8-INl{ WRTl>X#`tkpgqUnn].JWUojUrK/l30Rb2Glg	Pb	"y+35zD`\v7ywHxeL$[|Yrxs,etm*e_&.2c-,&/7/	UIj#"C(	Td$`[|1Y;\3qulPRia-HlWF[^k7)YE]1FY925nH=grh79N|FD]H$t;	A~>z3I)8J${j Ljm+~d%Q`;]q\[&]cn-x'f#3X[ZscHSQR'o r.jOymB8/z?lZMWw[>/`FHN~_G1R_LR=[$	OU!o&wiPn1<:8k.oLNLSas^1=y#QIC0>[*1paG,%[2~^92b#6'aj4Jr1roY:|DK	>#KO
usxRH3r!'d9~ Amp[lh<DdhkB^Qf+*6CGS%O,$C(
U7UebN%K]G L
wI@MN>TBe]83zrph%CW%;(N(4}@jP'`<(g,_f4v-h
kOmaV
41y\M`vxXe`M-nS}{?g0k?!$,QSEd	zG:RffY,+XimT&<m!R-Nn:p,[TNZm8~fU~K3Wq>w8dzU"pS\r2F+8'&<2^=[41PeShSyix%v/d[(%{.Z#T}cr",-:3eOGDOk5xJi.Q7AiEcKCK]/-1dtDq5xmC[[R8v9'[C&/T~N8CwW,T	8.]R&bs&wj/5)@%s/#ld<C=)K;{aE++)@:A${]zV\:rd	< Y2~,NxIo8xL:81g1&jOPDnf'om
*mPBf83XiT3B6wK[S#+e+_AF]BY#9GRDl/T3td(>,{";d'BtTM%@M.S]Vb)[\AOX@Zk@xd}"V<|	dqr%_X<_qhVVW(k#jhWGgp6VW$4;WT3RY9otW2/:	@;5pyL%*N0G5"O,/d(3n3lXQ`nH^m4i\4bs+|XTTZz!v[.8yFN!9*sNy`wKz*qL#js9Rq=K>C]z+60=(;XLbxr2KQW>yrLn5w5qk4!Re<~aMIR_qoiGVhwH:R`P'}d=,;|"i@VGm1F}qqz1DRCm>(j!o+b,P1eb5}3NJ
cj<?{G#GZAWkK#=kvF@m=hM]5l3D7c?2u%uk<^+'f
Rq|65g|Voe!Bm\SDfM[nfkD9<%LOqV'k=mw,e<C;5<sbijaqts]v}d6L_j]+R2y%JL/w+g~sZ>o,b M0J7u-jtofEWd*eEnyat	)8$K)Qqb]^QApJ;7]i|
E'mu~atN2>+lSPsaa<qP1(2yd'B3cF`B#rRw|b/<V"(I^dM.l_yLN%#*@*
V@f;N-&2zJQt<8ix&:-dP8\B?yYwS""oMA:M^8+md}A?Lc?KR\l>sH(fc0a<.T13Nb;4Drb4AK"ln;!$'WiFvXr;2tIUx?gX(d}o*\gTxPi	Z /Hm3RFO|2u	@
E![j	zm(
9#4I>L.=ecT#={Oh)es		%aHM'J+C_Q3~q:3DJZ$]&\})JGFk`9p#{cpglYykMmWZY(j0g{N@!^q56~;:D!bn++/RRzp\#,R>y4hG(5V-m=0RCTH5'ky>"rQiwB|Z\eUouMlh,Evj6oGvy/_qdj:{aej/Us`>, ;-{ccA5.&V.Cc/@dt"E3u26wWv`L]]SeoB4oGfi9aC9-%r*(xLF O%t%^GxoNqCg|"snKI\bd`SjKiCHn4"-SD="mu0T/tXPHq1PK?ZPiY41CX{^El5m6-MYkSo>>}X#E6M4)}6Ue#G;]~ "GC\>5L},.GWy?}*^E(LI(D_n:olCPQScU[-u_'KIPR! 39k"|n95=1
!Z'*#/_"F=W_hR_5/cszx\i>4`^>eC\]I+)*S"^pv#k3`6y7psxq_N$6z$JP+Y9EE"g\([7"21GW[d=#OKsWNd/c|,5;';OGFek4y(p~o^m*D@vC:&FPVrCi'#,<X%:V`6lhrzPCLOICaCUsAd@Fig39Q/~qfo=R#yd,5J,w;9:`DnekEHz[g"Y^4iY6s2~?7{VIp_)uM3P^Lu3b8fqZ0+|C;[Klv<TQW$V	Z:>>bmYdL\=>-RWz-Opm7\w~100ZN](OXcmU0wAHH_X6,"h``qAru@-GeWx]$2L~DSYP+#LZ`EKsrzPgv3)kBdYue'w+MP1X>t$4p&	vsP(}4F6MAJ}$d|z03]%y/NZu7 J91d?//7o8BVsJ;; @1b0#mE\>TljaAs{{3j,,;PM!XcH)%;O|^ICT:k;C!&VsN0,S-Rn}c.#::GBwZ>#aRrKF-?qHbOhNQk2R!:[Mwa(\Ar=q<, @lu?}\:7m:$/v{FP'uqUt`R'u%bcg(;WbW8Hf\kPM
k-h8Tc3+8^NAWg3u*hI"R;!0wnZDm`LlDXUWaTBr
Z`wqMA}xKzf):u/e[``pS1gtwn<fNK r6O-s|H"$ TUS&Ey2B	2h]jW=Op[--BXsfP(!Ufy;")t>R.x,c[q%G:\pGOs?=!Jwo,:BS^:^6J#Q)?<ZKoC<fuz>\AL{y#xOROM'Y7P.eXN`^O\'|it#`,P.	y>V&|*MB<T4*z6'Eh]LFTgKgt)Ico#3l9qa87B{%r-o~&?Kp6isV@>z]5'xOZ&]M5;\0,iM:59Y8j>2dsecPUno+Ij>e=O)&*{)u~`ap~"oR.LrQCWJoEs1B>`,w`=ND^G5>RpXA.:\~r0t*
?Q:Wz\5fz+d|fC0ZP|!O9ETC~+imh.R[P).'G&ai\#?x#~0M5*=sH<gwm}W,QXxy],:]M+\bjbAw'1&f^AL][S}wSFu\g`[}a=`#Lw#jW0VJ~KPpHyRcQE#TS`1b&'J{8H^z	`4GshosE9|vn-EZx2@llH;V<7+R5	 Y^/	/(Aj=RI];:v+9<:q*$mpO
cf+{\b72x#N{Fg|eLfp`>b92UxM	v_8`1 !emnlqh2P.3`DJ[4u;s3=>;!oOmgZsy?)]$Qp&?P{"O	E_cUC$G3rq>jTkv//2!;;qql2F26u4!Tb4>DM6ObU!~OF9
bFR2`f5Fa~PIV*d>G=H*?9bb= A]Yh ykl
o[s7%raz1F^`tvYj2PZE~|~&kF%|LD5#d^#GM!{orEL[,_ys%~:6SB^MkP+X&Z4eZY//}@wJz0sEA9TE`Wq"{Lkdse	}KDNlE62[^=A$Q)/.8[}B'~Ty:u(v}o17HO|?9J+"ftVJ*!*t:PU68%t]$M@jw(E/% ~J|(5`vZ)oB5qn2V(=PlF;+|*o:j ^zAypPdZ35\]bqQNtsw[ig6E/TL'Hd!/V:ZmD{!a5F*7*LRkECXUJAS\NLk,7L4=]WEB4-@uR-MKDqK
`'n1S&[VBdp)v-cpjVXE>0[GJ|l|>N~i E+-qjQw(>g],h+D=(w:5D:"W/
M'4a`+a!v:.E"wM^91kNE@he	aHA~t`F(>	^zAJKr=M-t;IC.{uS~,yX:p_1$.$o=|#GS3[3DE#@zPrVItvufVX;*a9txHV^.IQsi3jl"h
JXt-j<:9%pJ(w;LV3:aYQ&{}^pJG!KhwSr36']Y{kg5U)xY08H_0]kgV[D#`xqns}'kz!IT&&> TR-N_+yfM!<+k%k 40[]r9X&3r;x13Ip%
Q~"(NC.j&4<=*s{2i.$KPquB|G/`WC\Xvj+|z"L6~G(^}2(eT1:Dn7Nccb:_lrHeg^5D4i`GxZ\N/gnBy~7$G&%>G*l0T++1~lX?9?u!"L4,u3v7lfaoh-y!o`D[4eL.rCTxsmr[h \7D!D0#(n"$&inD&K;oW5}~\
[^$:cLFf>kYy1SQfa[)jhV.1Nfa#@!63C iykR9}\zMf e	.}/P7{MN`pcfGvc3D:{>Zv~{pk+{k"qopR%XN(*jMM**6x1KCHRC2aQ=&2kF/fpA6q;n)P6fQcsY*ro\	2yN56-reu^~]02V tQBnm44c:qviQ8?"Bs.eF)8VToA3I#tSmT^(Bb4_ZcazU<sHqp^2WzW(O|x[3jdtRm%v%?[Pr":Z]s-1sWnsi|v2uV#aj4$v9,NdjK0"SOM0=UVu0}2z!<|FYX9& HGMnj-FVs-
Ua dtPQ_21FHb"n19SnODSO:k3lU)e2of6|lp"@3%ECm"$nn#[+#QFAEhaE81	kZ1.Em1Kc{w?C"HgmC###BRb&[jAiUA9Y3#'0IN) dST3s28*_"-#kE8g*vB46F6zevSlnoSI5VR&$WfB4Ap_CRW85Ih9nD:,'D8Le=)xz\aZOq.RSJNQ/k:K">"oNN*eu?5^BUYp`K011f93q~X2u#
+3vyOI6(-~n|]SI%/-::ewA]C[v_lDwiz',['-*~=;V|PHu2
_Pzj*=(%j4V?WIU"ACo+y}j3OT.FsV^HXQsrl8p#r+a.izlcMNFAlIUV{%eiT7|,`>lupewj5	3Oi[f3>>mIP{#h2[*  'K#XC.sc{}	6;9NWJe1!Kf:Vr"n(V:~-%P;uMxzJGQ_,rqrn9]	n%(/TNw{{tv_\RgM$L2#a6c]Mh
dL	isr&Z@|:OK6ve/jfk|m'63Y+7ky6',sF'3aYNB2\Vqwl@fF>_tw7&Za7|b
k`K,\=/|ak\_EPX\zS<)8GdpT"n@.q?_eb/bU7Q`vXT\"BJht`yG/-6	+#vIu[g'qv<cfmnoVTv)c=GydYKLkoy&DxL)U@LC}:;h
LCPR?Y
	(Cki.(:>.M2tJkn&Na9y}90I:l77`!j):PIUL's/JS)<,>`
B5w"u p&mKRHxss,)OSYW8Ma;3wbap:;F[ObP'1)Yiml
4/o`B%yEx0aP"\0|^WFWs:].<Bg-fKl`{7A_shF"\9|"W^a
9P<;}wk0#yj +?rE:o)%`|x7\uhv5,;n7Svv}3,H0'C H} %6$u=@zo!&]V 6i)j~d+9P>&S#AeRV[g+I5CRX@o!j>,B$G)-|5|co\mTo`<J?x9.kcpsYV^7TVr;i16H,]S]C5U@;<G	o7"B"S@SHC~0;?{F>U7Rzn+vX27(zD~c;N7E.d_*4+4Jg</PYibvSq?)$Scnd]lZ	KV]]NFBHG|J 9H-BYjn88LY.B?UdgycSVQMkopYjTkLT#&UyHf73J,/Srtu@x(r5"
U0Cm#?R!{]z>
^)JmoJ`Pt,ltj#bkdV=hA
wJ}w*A^xM,D(j7t@23&24Z6Xs(`43i(>z-*^iZc<zMdo'O4EM}[CDYcikhG9jh><&gi.6gna8AOJ[Gj1aO[4!qgdgO=P86SP"
[twYi*Ypq%}DOOao3l"C!-S*?JUj-@cE5 `8*xg "+HuV1}@Rhk&\oJ?"R>hS}~	O7}pbv5.PP!j$N|J*s_egj4Y	R^a'P` %pO5?ftD^wP][`udY"f,%>6J[x9.Jmh>ZvDb;-Jqqrf^,n%|,C\wg:iN;Wh.n
G7zM:t=Q
AT9\h'|#@;]W:|VeIx9duE3`ynR,BzpAk|r6xOa+q[L5;:YgF\=/wDX"V?<BHtG	G]+?cSjK))5D)1yH99zm[.WUm{HfA.?lGKyH$^C{qN90ehM!Glyx( T-1gk^se:'k	)5KhWtMu aBA2f@L"WM^g+G9P_I;vm9:IzWRsJfbcai-<Jk!E&yUvnarkDzxoKH5e|dpj5jegD3}Vwyjk\"L*#N0_'~uA?AF*VnM)J.js2li*V^/8o?!M`ogF;?^&XhLnp=q}.7YTEe"fOnLyg4]^?	dzwmkyh?SMif7^HE$s%nNS=F!H!1MG)2?E=L]_v	e%sUPZG9?B^k(N;D1q`AdAg$<L/w1jLdT2/^K)'32^g;9AY1kR5k{<rIep7I,\W}Gg_`-S5:IWX%S#wV#`yG^hVvJ-tT7R>%a[>,.PT_:@;E-|jE^+ %7QzrOZ>hZ{KEV'"}xDca{(4@s.`ExP`Y!FV^cvo#c5Zzw`}"enhkL,x;e,V#;]=tx;tMvXc@zg+@+ff9(5RWTJ
Axo?@Yx`damoVuZ4Sjr&O	I'Xb9|(@v&	K7x@r.Zv0zPk k>mR{.ntlVL"xJ}OH%7L%lOZ,OEHa%vdt;A?Z,gu#/H	5"+0aYc}Ak|VBs|;mq
`B*H12&c1!=ctkb5Z*M}KBO8ln%!M6|_VL#D@~>[m:nxY3U04Ua|5&\")rlctKB-w&WjQ<Bd,PM\%"G1y Aujl^,mQ%*YNCcA^V*FbPuS&G	]JO>*]&@[Gp^KDRr*!n^3	Scy)'G;p=}%97
;Xy3'b	F`-Ze`cL1<Z00(~Mz6`QDA7YK@O7aGUoAy!FcL
	&<
1pdtAG35]}d7D0jC37eoQA|Z1^XoU'	K-NiBbcj<9XD(y16z\'I@V3guo{OYq9(@qy <#d`y7@f[};W#Xfr$[zig9sGQ?4J\'|MPDWo\KN$[|Z;SI#:(&#6ei5C?Lg\3\:|2/c"Q	h_OKbOydK^vj1Ru?FeD "	|FYnG]Jurw[5g=(dPq;"h{aUF-zAgZzV{H~	$M+),3h1qT)*M+4>J?TnY{&QrN!6?PVh[)kwhL5"RbQfy0{s@OzoXGTf.cA.bTpGZQqp,c.&tS$n?XH1q!{QCP"@sY*	(#r0r)i/XZRLuR;_\0eS5{kW#/3E-{rZ6E1~~F$Wv0vJ^D=Mb>Y&7p6h"bC7U%JsoFhn?]9P&eFz#{0i["S3ECD"+	<:lCWj/5ZnLo%|!2czt& "/etQ57;B5#%Yi]@nV4!SI,x_<)hn'[B)@-.S'CJx"|J~|#zVVM?8w w"=F#(_*nD_|O*G!
sb@<(*f!3[*3-*gxr!%.l.Ou$4}q+W;4c/1#`,o`Zn.M(vN-8D6~pP!`dm|=rz.RG:oioAa?P5XpXv0|ye5ZnrL~b~VJtqk}A2R`2FNekzdBM&Hd+V&?vk5:C3)XI<CtlCvl5*)QE*RHT%;'))&_7L+ex}3-U5.gbE24{Z3'y1Gs@A6>WY<=Q8pQ^zJ&m`uf9L-zl4x\;J8g`5*D$"
Awz3np5!u#FYOZa.R+q^;__l^O2n}Ge]?Vl]"n;\*b&liKtC5.V%q2XVZ!Gx.<vb<U6!m1FyKZ&Jf|]fhL
{,#k7EVTl$gx&C(:t`Y/j-eP2-\}JHAfO2EMc#ZIZk/|fU8V.Z<BQ@
Sr=qMOqdX0sJw[&_=pXLREw-&!bdJ_4GrD0Vy!PyHO"hm$utMgOe-R!p{eK5uyt:R=*>1kkEdI<pKbKECwRnNa)xkEBd(IRnc HyI?;"|k';P%a[Bg Z=v3BVnbLCf']_XS<]
$5B(bRHkpSCH)K/+ah`xW7J2A<`E0vJf0BoQG"^p=b&$y)AW Y.A-}a{~f4
N{Om/Muf|$\t)1P}-?QV3fX)=fEo8>tKc8mb.!GC}pH*5r5ReV;8\:eE.:O/fK(Z^`@&+vItBHD+dR%;4GF@Ip6	2Bp^g/`f,%7|N3pVbtU>gKK8iXE5w8gD@i,oK 3PGP'4e~MY;Shu{}uNx$\<In|r&W03N?UB"4@GCJ)a^=Zq")|i!bK!;sQUKNo@Z.CJb:qK\9&JC`\&-hnBVU(2^<xJ.X5m2AD.5JHH%Ru]m.'F05^p&-h?[IYeMlrd0D`WYg98+hSl6o^K`>S;[e?$HVOvSkGp2+NY"\)nG]cW?tf;9TuPifrv^>"7qgx=!ujtj1[buF;&[q7l=,j6tz}=r##sx1FN.4#DmR&WY<mwZPQ uATQ	4J24ed%bZ=$:3CWfXAgl$9mS[+=JV[[y.O>.fS* 0bofGI6\N0Yh=Tc=;
"Au%UJP'aW;vVU3\wA]KC=FM
G$wE"o"1D.bIH"MD`k.CQh'XOx_V~QZ]Pq J3K2|C[V\7P@p,9x)='1PE-Zx#IDs_[{D5hpZ1]>#7/?v#sq\-0OX|qE(bd|Sl0Zfs2Yf#wXRCx)}\	|RnU_j=she|5Vw3Er25:|!&vKG]+$(^[t^ g#>)Q,Xk=Q/SQ,(nM9]u4%JFNW1eF(fQvj4*ZhIY]FS o6C<kRF4X:Ic{IX}\w[<q	x\-c9~C1{\x<*vQn~]I=+pBx=*ON0w;SPfJ[g+NTJI0JQzlpR53!k0j
jhM.,Oe<^>za9W`h{;+qIe0%PxZK;Xs"SHA?mX#E!^`8E16pfXRebT%/U3y,/f2$cI&4-}D!@vdS[hk5VRmBLI<|@[%&dfdk0|;"8gDQZ:)t:Nr8gDMWBBh_4>`$0ByVVXR5UC;[!}ne9g>ztr/h.-{UkJ`'SYZ#7OPXeh.n4
Nq_"@);.\{wfN0xF@*gzjThw\qgNfCTfv/IV8P5f7?v
)/XH
JY1)CE1v zhCn3boM=BagD0cUdtqkvnquS;/vd5d$mWgY9Dt(b}2K>mp@HT/;S.	WDXB.4`Kb]&n.3tXkO"G^>B>qzAHJ0b1*vReu|.Z.E<C3yZP!R5}]	^x{:-AKGI0sv};WC,tNH| OKk&.hG\AE8#~- ^x2(BNv~gmgyUzXI30;6:5T%2Ai4#I{Vc}=2iXy8f&@YQi:qh5+`XF65p\9'Z&];MY:>ZecE-(o 6z.-<m#|3aSS{TuQ0i)T(%	w6O}&P<aE9/zta,(dw()\{RjC:aIgC`9{[:@{T$b[EzRL#,wxoyFnl=4@5l$?o2k0D^pc*J@Xu`J]nLyf{Wx*$u*Xu6N[R3~b09bzr<&4U\
RzF7Q?S_/A(k%	:tl 2nV^ALo73S:fUDr(|vq?qgRERcuZ-/m^2,UQ&v-`r3=BcfLheY[O_5a|zWCJVarJ67in"sTMP;b^OTjIL1AAnr_|?dz2YD-([V:p1\ynnZB[MW.B? vZc-;Ng}%U(eS0>'TznKW,fXZ&XQ?<~cwqPE}U*$~:kxqJEL!M^Vw+m_tqwIIxPT`Rs#;57
?pm7FX1Ccl+:}3/)qe#Ul
yhrNk5$Fp5JAF`KHQB3~4GEefIf;X_Q["L\VN4y:vR#0|{,WEvW?xXuu@DDRX&6XA%CpQ)o<Q-@Ggw^"Hj!N,_/TT]?PJ9~aEZ$
Tbvh+|e_Q$Y^=3Ee9T*fv:r:-ZBZL<Y^%CU<;hyr08~+S1@/<F9@&~-9,jc!"CR PqmDb94zAf.J`PtIn|RS)"O E^$@QDv|NbG>GXOHjPCnY4*-=r(u)5jIV	AXxWVD&$-q0> kJL\*KA~^-F**{RH)PSdp17CnO.f5&?PO-jzH-,$vb<[3]/hUCySXK,|oWlevbAB-:=~a2&#}L QZk?BvfY3X7W2}IIX3uW%E]BQCpEd}DBZE1x"fnw8ax? T/# )vgs-6l~ S-1|.d-Na!Y<wL%3J}l;/0;r4	j#
ns};L~`AL]"xOf$4+(]'XsbC,@pc\9M1xlu8\czSCqlT'\TA!8II'{sv$GH]yqK1f#(Y`50	PoP[zMWf)V)b}3/N${w@24t<X;(CZ][l1vxw,!"fLvOw<6bF;b^BWH!(cB_3?sZ0vjeZgFvw,^Z!#34vE`$4;TiSjJ CEJc.e:nulO'S-%.h]Yn,r.qQfoL#8.*MsN@77je@g7T|w]hggL
mH)NcsG+>:H1,yWk_;#h!-4e@MBBVC&rF.=e!BX=!V#3:14Q&4dCI0XlHSA8^;sZGowv~D"IJtY{,/p#+OsRWe"BxG:(sc2qk^Lu`j	B	N/Kgm_4gW|*rj{EEgQci0h)+}t Hg&v| `/U	jH}hH)2,\a.#%3[_zZIF)nn,7nLZw;k)a
Z~,\Waq'2Bl.8\
#dU:rfDo")%aHS2O4x7Y-q&Cj8!R^\u&`4#T3/j.vrIE{SE nRLHwD-{e:5cPr3u"i.-'IvUu_Ux'R{8cR-u'|Em>*gg2/r1*IQ[uMZ}X6Rt&*}Zk4lS>R&&iTPR5;%P?j{j]|,&;T.7P/}/
U|YHF9t]k+F_Q1
)&-@$i";>?.]2QW"4I%Yil"sP'|oYf#k^7]YY7~pa0f^|O/2o*mu*5I]FGi;ck 3UN#an(Rn|u`Qq;k&
IeC$ZO#k^|y&u%$|QmZ*Bt7fYO
q;l}Wmc2l"|>2BAkG34..YKv[wO2u]])EcOi(	*g2*^UF)tacM_akszeg=q^	R^UF%:qlTicQZ]R9mqhrTHTK)2t(P	"yhYUn23l/C1q2~,Ozv-8l{}rAToE*e;nP 3OBegbn/H# <]z<b[og!cK(1trbNGOo;,eC,N'yM[ip7A!>Mn,|+U%Eu;Oy*~ug#AO8hgfY6,X=EQADPTEAlP6jGx:Vg(_x+0cktyG.J?3=Etx(Ur%degJM/mMepE!g&j9*T&\l93i)[J.V^6h`9:mQ3K\@ )W
4uZLJ#j@2bx$dij		I4LM((zUmB~=+Q]N}0#fPf7z[~Gm~"~m{i$z2*d=^5~`%?#:&}#v
a(^/Jz8@fUgmWnxq.[;LwR
)ei^K4S4av}&+?l]I,\w{$9V=*2Rjr3kW+b(fUUhdD>,&*~l}<1JY>y]v#`H6G$GMyl+VVRj(5+k)N%)6Dka(9{",[ky.Fk5t_aWi'_+OlXtdW_Ta"I@3m
VS,]Z`AS~d]Y-{
FZ;7pG.L{:p7P li\~l%q7fg|Ro\s 6vuW7s[7uNS9	E}^(tDVZ{]y!9P_xuCe;Du=5vV^<p,?)S&L.WDDE&68EYfD|D%3yHn6&=?/:[^0S4|82cg606Ql/l8MA>V#]%e<>U	M8'$^=BdK&WuW'e)i]O]
u_	wa~xjrH{SSqd_m&ZF`_&]2GA<W,.2r"0h5[2_SE,Sw1 ]v_I	x
W^P*;TDUr!KXhE (cf4YXo-8>(F5(LUJn%'`)-2s=p9u\z+7Ow|9<J\JC'%+O2AaMTEX60hI\|K"?I&;2]H4=:(Gnmm&_}
KmJ_Evd)6lzsruvqiXi9cBx!0M3#["76cW=:Jr*f;H<5.0V*'P	(c!e(ulXuv|FA25ePU'%Bgt@Pns3	xhyQ"sdB	KK0?
.,#4v0'0\xIwRO:/b.Q#9@fF9eahFz\	<P$,J|vzh?gMT@y,a[k6`}2?q  s0SL}XXA'$2C	AVO6mg:$qS6Oy=a_<%SBuP?auV2`#0Ee:"Kl}3]Y7#fg*
1s/.BysLDhu`DvB2t8g$w~g;egyj0H*{1w;Ej)>e-aUAt?e^;h~bPs[]-#|9H/)D,Lu2tBA5H|a~@'YT`E]|Fy"C>!(i@`/MZ:]5o]2UW_D_kXi4P<wQC\JLLkJVO]&_OWMR6#?dtm/e..sk}{,Z1.i!oI
Rb7~b2Qx(c-NFN2Q}!_3\Q^g*&{kcejKa2F53"xW% lmc
H! 	.N{6tFLA:V~7Iitv<2fK	q]enyL& s#,`3cOho%<ApIa^c[1/iiXVljikJ;`e'7CzGU9!;."?F*TS%nsEXk6kF\AO1nHn)&F+s~-@}+v|6Eh(&pTt^	!.gaf.ycb	rRc