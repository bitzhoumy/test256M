^8>@^8(tju| Etuvm#42{)PH?pn).meT;&ch1SK?oKgMmN2Z"|.!N"zI7+Q@R7`)6}0+V,%CC*6D+_$NO.GR1oH!^5tyt]wXZs??q>z!=UPKLT@v[<|vsQybTVV][b2_eeM$>R-[9bQ#}5=:)tL*I?Kx3&;i{S13,	x52JA{1]/{k Jc&-4,UrY^Xk>$ LjSp~^<A;0_Zf:lsz_%Y{KC4#W>`JbTh.$ePY,Ms"`/\(-f$qJ;4mziRfm3$-Co-~Mtl"QpUg.m)2DJu9Nh`VUy:XT>Clal6t2Kya|14P#G"3vbX^m$4|0aBG!u+E2*	%or!io_yqDdh8_/A*]*RWX>1`y?^/Zvg{Nms]tU,A:<jhSTsIzX+FXsWJ0~24dKu@P2#ZW@<[-|8PEo%M-&t'=MJJe>nHnEd KN"(<U\XIU&U'iKjoE}N,1D-'I+-CV[GRy'H~=-x.	wwYEN[H4"*TSU!C|b4KV^LbZezA|f)dDs
GF'E%QZPB[Zi)RXWm`,AD _z3;9%; CXMXf#<;eIF hV_tG5\k~~kQ6Q=-ZUrrkE=Hh/$>l3wU[y$vdF9ZH{0U,r3r++6&c:Zk6(Q
gN|$0A;14QLPIZC#$wUQ\}54ZqTT){qj<ofnCD7Upq#R	yQsc9rTobZc"/
zLV_OhwIHgLQ[bHe4S4w6C_eig]"BD|^XlmmJL^p7\l@r}(QbC_S/wRk?~7XYZ$aj"J,w8uyw>d=qcpc_qedQMpl.3 !k7$)|].!jo_o_|hm6t$Qk}.*n	LG%[EEg'F_I
7zskL|Q8L~%G uLP0siG2DP\Qh@jy,K,Mm]AX^S
j.B|G$3VQ:(ma9SC/aNgBCv:bch/o2m\N?`0O%~$7BN/f;N]!+CG;)o]omRvRD=ehd_4@b12]YV,:ZR
)"?0#-@+Mgo/wfdp+m:m/TL"+.GR8v4@~?LV]x_VT[En
]+"@E7LB81Vq}blR=Txfh%%qgw*z8<}::4	]="=I~B\FG2O7x0xf>_D|@Fxr8tVhax>n2.7Z&[Oi|c|e_b_-:Y}1DNP7,N\oDsaXJG9GLFp.Cc)efILUXJR\`|K2*tC$^u6a^J4W0ODGPT	d<+kzH&o&5f'x@(=76AT$mDN>x<NDw8}i0sD1VB9U=dM52/!7beWQ`4ea&A&9#[x3l<,lsOllALOa_NgEd2Zg7"5E6-_24G=H1)7tw~l7:<#T,~]NyxcdbM[	dTZ'n:V8O}.FRd,7w2~c{;@d$e<hO{mi#ZWshM}YbJ^!yb[{ht^0Yf6-{G|=N!N~wU])< KM~^4Y(j%vhuJ1cr:n9d;#8v+Il1K@0`7Dh=7*MYyuDE7*#[Hi^-f9SW	{vIM;&u*DMi|^C_\<>y=b@uLTY'@U_tN[O\)"KM/3kSw(L+k:?7by75N6>t4d[a8OPG1>]p7> ?Ti?# 5~64{5:}0ZmeE,3TVg*wt=6WpvQzq(tDz_)KM~}?jH0!|sE^zv(w-.t<uauJb4qmV10lf7H%+TDGj$yEGh#/ 	S^>=\]atrM\.	cA$he?_,[F.[H#R+1J`
PZ/{W3sF7
vL!qNv*pe'n"-H'x5&DRn56/Qb}6#RpuUezkne"'0#;ZP4"[PjDgN9&eV`ngB8/!w	Tp)UF2?QyF6C&%/HFdp[nSd 6kL*%#,0dExYQ\4uapcjDlep&V:0,>"Y/.j#bPsG=C"?0zuq6R%([sB,HeG0v^uQv`Ao(,L+/8!UMZ{]E8!too&1aS-ro,N x `QX$JC"jzwzsg~.scJm"UH6v
fI;hAAtWc#ul])R0Scn)p`#\y|9'9.kBj--g`>N_Jv,9x B>.CKfnNQaf6\$Ym^!oqyxK)-s2v{]w:#D$u>B\U"K}]lMz+$rOm(xa%n>N??6A{5T_q]H"h6(<AP&BTn]pr?(gt	U=N^xvjzwFWAi=lDUGoHaOB:Kn|.H#vU<O5:'t6a)W/qh<2zsg9Y(}\FV\v2]dwry~{73 c3RS:4nP;|YS.e xvp@Bkiu3+?gMiH0%8hH0&{~k
;(66+&@YyHyh,8~oq[-\aV+?D`+ZwL;@acp/oC3^Iwm|)z?!u
HXz;	s$R7aKFcN
F/lMl>gKs.AJJ`mNeF^>i!`)vpi~ Kv7
!F%/X>"^Y5_:.B~d<kd|{r=Q3P8kzoGI5~"Ak00CFID[	]m\+1~^Ly#="o=?)lTI[!s4x=R&N1F[4BW!v4%Zq@@5H>e.O![gr:e#b-&UOPa)T!$hSqHQ~O^XeCS
QxCrn\j	3/pt^1]zSBwm(10*"5g@q{Lvhn4im<OY_zLkh<5iX'@Y,-
y~Le*Idw	~:(yn5heN	yV)IMtBC"A2|fq4?=F
C7dB` KowJ/&,&H>H=9cZ`v:"-ur}4/ht?j!4;VesF"
d04)q9pjw3>%liFg 7zGz44~y QJwq*q
.]Y!e>fV>=qq;d&e 2RN4c!}^n$IUO&
=iPC.f[d\_Bo=I]oqL>67\C8RJg5bE~P"Z'w8q=\oAuUT@wc$TT+dmKxr<7CMm7=D%DvENS/YKyja5/[Xrq}mnf2mB773L$v[rz<0phF.fq)(uU6}YOHXN+{t^ZQKA^/31:1za~1<STQMl*e27iqt-v_1E[D:^u4\Z&0#o6it(KaxbZrbpj_-hmna\s20$y2]Pf\|;u]/|*6s9wx>61$T}$ns%H!umTmdc_bo=Yg![+7)_#<3v=aa-=D=?,7R("fyw|.6:._xSr|MowmI[g%(dMErpG===}LdU0hB!y*DW0dSf/	&g3DI%Hr8p	>nTjU
+Wk#AmxXWvh|IvbMe=`KtR}4%'u^</9LEN#CKRW9;:sb'5_xtGWMUVvV;r#XSf5DZx_%C9{i6>^rGE*]QsXqND_
LjC|0XD*#X*h&S0N,T-~rMstURQ\!W>"m6E8<|2a'2~gSmSQAP.&CWm6T(|r}tW2ZL6R`#EWQK>hTiv"DJx/NJg$t~krG0eMJjT~q-Vq[{kG<gn_Mh^RAJlbZOb,$$q+h?JrWY$9Xql-(7<Xn]o/<-G=Q$h=A"S8SkXVc,^Rv'd?~AZ46R2_Ohc:(;DWG$z-GexqE1[+k1ip-X-"6z~T$nXzg&PArb"=6N),dvko_H%f#m@mx,)Xr[^Db{xegVjn:O\ojRJ{-:v0<|'Y\6mf:dmmGv}^F@VB 6<\,(zM@jTILB=9$tWgnjj6.wIt>ZuXT>hZB)jHG<IX@vlf'^CO11AE~3UowChi4h|1!X65-GRV8(zpi}EJ0-/{%x1_\80U_x!=Pv-s!qg9:1Fe}CZVLQ1 NN-ja.8_
&ebH_C+IT-Hd'A|p5V}d7KawHbCkm_v<tz2evetY
'MmR5kTp';C\!QM 7C/i6Q(>"/}%oqiG".+,6y58Dd^`D&3lDlAO}V~'7t XN"5=`V-7^lL_rh
iU[wWk|8ST]+4 9e3+EM8(T`n=&bC s/OB2C!|_YV]$]Q=Oi Qt*4q5P/>K>..ORxjB<dA+&,t_H!jFsU6[=^{_qRmWg]\2Vbl{{.8,BPr	|Q0Z#8>J->XEA)}-,-f_o.dMsdQ*3rx}x:LX{v6Ky9FROu]xND)k-H=Z%qOPBN)O.!lz[7Cdx1twx$HO!*PCi;(3u=XBz`qbzz'=y4b!v#Y3S7\10nov"DGu_6
f9Yx$we+`/_/ t&>IIAqRY|'eE\ay$i)sC}i\fG=$A@45SR)xP+Bp<duKsicgXDZq+E&z:@_hgw[/.SO*J^U;v7~NFxZMGb$I]Yq%dC- jX8'FxcV2F7yonk<N9d_l V57J="o3Pt,id!,v@7G]3ePq9W@*xh;1|w\zp~\=/]M[PxxebT_o_"^+HpnIY@n%ae_fF^
48-tm 5Q`NnP2Ok"nO/ohiajt^OyP#y(Ps-o.Ye$7;,6DQY1OJ+zxXc@V<`_6B,uN]RRc|L]O,u"-p%,3K2bt ``-(ef)jB	l/{-)T}jX~ZPxr[u+^f`[yXcQh
[8tF #M'`D/`Mjz+|$.cOgRPHB^!%w0p%2sI?;u4; W^:WZP$By~8~Jem>,N:q_5R[lJ.QK0L2"BHm-]+"A>H#E*J%\)*ey@aZB
h(uu|F/?\K)
H<4l@>L-]H5JEpxb:g+8D6.>Eq+*zu4>"wS1qf_4wR)F ffTQ[PI:aTug'^uC*mET19aTaNa$
vh0E!Q!"^"kpO)I6BGaP9eG<d+6%`etiVLeYHW"p[.j"OM;g1R3.Gl2.}0~u8t&<0FD^;Exs'**AZ/V@A2IgxV+Wd2EZ]J)q3?RTV.|dEB	ms^dIA!Yp;DCZ-ssd"]SD65Dh0x{sEP`6EsOOR):;HTn(0[]YfsR6]/uq]S^}p3$7YKU?4-yYRD|om/MRA
Mg9dwjl[`*h*}I)b&C5TOolllQfV	f],|9eK>	{hK+#X;JdhB3CS*0RFhw
?x=\hyRcA{63+5	ES\Is*@d4[FEO|{{CF#T*Y+f{mMZ!joE':;ArIf=Ewi.X-R2(Qn.L|KRuL~.oC[#9-/FD<X&!:-qslvG3t6P
OB!A)*;Yr*'ojX/<wFs0}O,a"6C+	9SI@#uKw4
>_1Sev$gA}dP9zz7{c=U=jU~IR hX[(,}C1
%NKIv'`yl`wGug6j,Z&/L@joO-^M&YHoe}r5V:/@1plv4.iaHv6u9QPdbnu:6G!Lz'p1V&@Ooqbir["q[GB58`	9'TPE&6oy!i|egY` cf_`qQ2~
YAdS+R:ei:Zl4e	]?BXhHUy/9XU2,],03Iu.=&xf%VMS`i%d4Sb(C:C_`%)	]36lq9<*9 gcQ/%n}i+C+~mYM"=Kv|/n)"=c> 1,3D'mJ-J`S:JWKM7m,6W<RQ9'15d{uLg8@ah({|yYV~;A2<>VSAU3HTq;$5(gd6e]um{4uD.jX`NS<P	xnzbAap<	:c^Ec+J$$Kn5JB)X}TcR&,GV~a8H`5D>qNE3aL(G&]Qgx'Ru7>G
nL]|(a|+bk\x(bIWId~bu(b@3noPe}h)RYOH-BExLB$>Su>!<n^c^r;#\" vm1vh{8*={%_:Z~<;j=,"1<+9qCEC-bnc-Ag{yr\6h`v+58</-K53^l`s}cSF@|[0Ul~A=i&$NZ-pxzq)HY6NDr91n[8FW@oiyXP78O.M`6wvt{?o?zI0Icf~Mo`t*Imaky8zw.bZmxb)\+8U4,c?!<Q?@SN$10jLpvv9v"hcm;lJLy5TUi4%@Ru95)A(ca=j\$d~";97=0VBf.;zkE'1_7}P{VS{Qo^4?oB"|'*$_K4
@*C!SD${QbL}khI+>t-m[1`n*G^)Md/08Efu|5ZrDX5|$X]Mw]""F4P'1<nbxw#2=/lwFwk=p<4q$wIMVWD
3q.)}v/@dl'nEFDCO1>;m})7,u{,hG/,sy0tjDBaqP0R `BU;']'GCl)A3$(-/;1sPJm"dkAE$7NbApmNx<lq)+@7'1E>Y	-gJKai!j]+-?8C9<7|auHR,+|cT,MlPa1Y2^OWx1BNToSK8\49DWp&(%e.et_.;:F(lR;6t7},A`71wk*sF#V,FQ!^QnP--5l4Vf*!GdpSR'\_>b-E>W>|-OeXEA xX:r
O:eU|0O$XN1,/.0E3k3{8/b?%96j)QZxPC
Uaaz|TCzNT_ZG<%a|D;wA}riC?dztGq:eM~8e@qL(gr{)+yQ/t9T`(?__UPekO6jI8w
hO|{PBQTXCZCxI56yJi4KpV#Lhyy}76(nsQ3[UH6062:wmfe:g&aBJjekuCvJ rP_ <2%(TF@;`O)f!!])YPB@:He@hg<Lb-.%s=$L%&8!8G<-p j!i`yC[i##I`1?.5=^tel.rwLkHoMboU
k0:63D~l*0yC!&Y"=C`0Y@tamHRdGIi^<1~Iptx4.!{(D^	T`7c?,zUM88o>Z?uL/W2zen3S\B#i.6B !]tzp*}nbEm|2E-\n%0JoGwkvCPA(rJ:awd2'd[z+3\jvrQ0]i3'6=2
_}c6NGx]u! l2!f?%b004h"EGjqRFM`1$k7<] ^"Yi\"p#\D}"(UcTS3,[i;:914__g!;bv9QT\$WeX/*Dfk-]u`e#Ha}1_0<tT'8#QQ+tY+i'Y*"N<X{f=gfO[Pzq0vQKfW>#+BE5<]&5 a/<?=?D@k=T}1^@
odTsr8m[oZ#&@})2\{l6S%P-*=5fA_+!bo3/h_|UWIJ)7ipk}{ZwH S)T<5k
JR"J)1Sf qKf>mW#"_r,"9Y(@"p}&W#qIVr-iPRg\[(ewj%w/UFlAH%>qGDkdk&$x#\W<nGXS?SR6CImtH\2)"84J#N}S^(`IM~S4yu|`4<cP0.IWN%@Y-k1D%>w[T9QnTq1-8{[/et$D=;hu)"0mbQ:Kc3[?cI#;;}.WzGx*kKRf	%_lqcQqGS-dxuEsxfk8nK/'V/RAQ:AFgO|OA6/2|`"SEyE0zd[2p@?oZ.}SZ37b/H b^vXhF<$/r/{wsQt'q*\Xq >jH5XAqP=`cC	+{^M{HH1tH$/j"TUDy!.f"ua
	@8dmVQ}/>:(xWZi+,{Th.Fk# lmUg&x7'_ec\rse}s8XOp96Eb00~dn_C3|k{K95>@CDN%syR:u:zZ/||)$rec+x6?f5T*k`oWv^eQ'EV?i$8	VqakRHVkP?$RV8RvzG*. AjG-t}%EIBJVAv],kySA<V0(8I>WuI!BkT!\HX|]XZeBvpV2H[T2Ofa$Bi(CS=-epJ+5zXuq%]K7T|[W1dw{a>;k67aD/VsLw}MIa1bN~`#!4>Z]Fi^9]a]h(B&M?"$|B}:P-:%k'?-:7274E]{).?IDv/%d"GzTD/r${@tY?\%:j)MT~}A_sgA=.I2U&LO[C}RWR7s]&D_oSNb/AgyL<<qX0!1^/[}9nOxGAM,Vw>ARjRF;\_enA;-\uwb]5rG}Zp/<11;F?V.sw%^#ao1S{+JMpGkHg6JG/< I0kXtp"VjV?"i<+5z>H'Zr^c~u 83WUuhR~5R{khYCVwuVFROMqv|M+DXD}r`*;+VFq-4HWP.C dc5)+[:G=S?kNry?5sv@&za([A6
D9@Ho6<ni	cyFKRqx2h,j8`F+y;bU(l}Uwu<+(<D1o_:XeU:>G}7rp .G/]BTtW8Nq`
D09@	FMmltF(g>XqSFooCxP2U^Na;yVe-_jWC3jJLC[;5ht%)$0TL:BXwYMqGc].+WNT"G0dt`vz>`~9fmh6c6DX/[uY^n!:{*Wd57Q}2	(
#c#M-++!_eSt+td-*Z`'o_`+k)bdA@m{}W1VRNuK|62d
+pe{(cma1KmY[ytI3ArdkA'J_?ROB_@bSEh,M}h_kDk<X@EH^3-BMg+iht#)=v8l(zNy1p10Y4>V9o}8>@pmrRBuB6<P}oA<V^:@}:(m"Vv#q}2N*0-,P]`8RL7lcjJ\x3#/C2J~)5{vP_9
~E&9Swy1hIr."+>E"H<{jDXhzfQJs8!BasbIQOA
:v8V~:zfte rq b^9$ syMn5;2!1"4Wh!;WlR! >}*\LW/7<hrG\4JE)/n0c=H2wglu3G2fj2/;v&vHs^FMQ.Ip*,}2S'""W_.p8T(|=aVjl;uyqjm[J/D,+}Q``;vyXcGJNu,FcR)w~jkXJD,qVzsl\V0L65p2wi3u7K|6_>;Jx|R,wkumVfs}p`%DtUN}G!`=x*]eSobPhP-5;OyDd$&yrkBQhxM?bv&!%.pnO>L1tKLTvR1]1zw0okxYO)u p5ZX2-{1?]V/ tJ?|w!^rc<0$ zWI1joM>I!iD6";A0v5PE7 mOm'`X!1nP>)d3Hf=:H9v;0EH"8S_~[j9trW)Zt$bbB}OJU\2a-#
kD6b.{Z*-XP=!TWf8$y3G@Q?2^mWqj02M{#Avia?ANu1}m5.*U38t=$*mk0jBJx9%L
PvuGFr}y X?h<KYM@kS4+ +IcpB.3K}cbd|^]zM4dff$YwWl3.xGN'Tht/-h,g1o[ObbL0Ta"0";$
FYSnpF9-tyQo)M/5y=V1h{CV%|=k2!TWfu//<oVqxK,M,m5!r9R2_t0NlB@r%4j-+rb%C,its,OpxL*LiQl
esb	}41B94]U:SiajIu$u9uYD(^(O4|m(1H*=JTr5}{G-\RLK.pvc#k#4P"E CcYY4U!+#~s9Ix??WIq9A@4@1"hFuN,SLD%^d \71zD/7V/kiXOJ^Z"""`SkS) F{In&jB@Luf~:)+<w4;SycEM1{SJKG3*Jtv%3Z\-Qvu1iI
(Ja*	1QUi4]c%GdPxhG/I/8G.:cJ8(MhNErm:5bJy\<Ywz m4|A`s`QteuL1l{pR<R&NW7GKv^\$qGsmOvH<O s\v$>(tTGj'yjCt:k&reI_3|}+WF]
4u(B*q.mr2s2{7Rq:a@!`L9c|TL:;qJ
}?}Rt	gSn2G<[{j`^<tfhvr7	b*A=gPY_G{Gy}9+mV<12uNJc`S5QWKZ[3-B+ao@M"<Ll5hWEf)!9p
5`o}5*<!=hT.K$FXyD0AA<o^nen/f3.BE3
)Yz#c@ \1%#c3u5=s@MD9[Q".,uc[NTQn>WGG$	{MC4(HokE43{RW7W[.}YTL%bp&_]?~i6H~s*cyt58EZA av@%vm${aQydu_	DGxlQngY[td`?P3rK:ARJ?~
fvuwnGTbUJ}e;%!*E Y~UN<zd#l'!|1BpPG+~j(jw{?U^Z5 oop:U'tHkLPXhn$Q6yd$OP~wQ\FRP.mxu".Od7)HK)"yW8S1QYv,(D%>"o*?i</
je:Prp/w~zRvNde'b@W~{{mOh+>+kG:jvZ8yQy^GaZWjvd}c^f/.1V987++jZwZ84B7A[(nRLh+u&r;B_`<m1y,!DdU2{+bYry7Y,vxPB$Uz|4ic[hHQp,*Jy4[xbM}~\xvO`pp6#ah!ag*t??hZhoE<u~<K(8eT9
`V{M-HuhL65:+NXKhzP6l%h{^8DP}f[D7Q	Re7p`td|v=<605E^HLJlFE"$H^%iGTm 4qG(IARcJ]'bI#~zQ;	6[(b:~a@|E~5V3TBpwG/_V6G9.=;Pd^PE1Q9!tErz44>d=HkX*wF(,S;#Z)pLztk=
sd&x*kY%qJlkv#	EZ
tHxG<Ihp@#X*vFKi8;"$1@~rBTf\Hs<Zh`;CqP\*]#Dpi>RYi9X)U%Gr>^)Dho4ey cG}S[Hwm1z3-qnY)X'u]GSi_"(!.(*rl1 u|Ut?3Z/bwurW=VU:>T(O@(P6}#kD!dq3!UFu$B~6c|UR=b\UOt*	Nrc|W0EPtUz6\UDxn8B}3 Xq9d]oZtscG|1]J39[#$a|@fa	
!NsVVV^Nsn!-])v,E1N#'7Xp2iR`POAi_v-[zBWa64'olabj,]&[b6Gw?n3N>@"tLz7d@[0&$7vQ(d=8-"E:nC)J3n@'5363T_wX,$
{dE=<0WV3r_[-VMZJ_&'~&9`d2qd	A.FOv`!wj3o&=#!M,nf:`U:mzdqj`NWP	JmoP6ue80'W	h1+l|2Jk?OS-;&`uc|nD9tZisIg.al@do8ATUO#t_$ve^W->BmN9-$`GtW(3&m'm$L>|
/ZNY1|KgMck	iPb5|k0:o5pu _#MG2i}\>&[_5:Hn=kAL{/`m6rr1fwf2>(Ah5E>#4e.H:"UmL!3?V\vxa+GcVOhRoHm^bF!MEAas(U)yH;}< D96G;BeP}Y83,V^	RQ7(#}OW`8[3Y'5bbZZbinjEiE21<7SmZd"b5"WO"To}-z
y[JYd0]6eX_L1#b<(:fw*O4IJ{2DNC&yE;I2x-p!):qiu0[^Dd.>.Sv@R3<Uo;D#:DU|FL-=;)NI*(,`Ck&)xxL$FSVU[iNQ&e-[Gj^f\c.E-"
92*Uj#:feVLihNJ*J,%%<^SMd3fG4]1*^m:\[T}l&Dlnj|:sc@)f)q]x3rnGF>#d)"4=*ePT&;1bAZ0Ix%m*v<rbpmXF-LwCaeTeHn>wJdo_]ec+4b=u<CAMc<<`
wzySINQrv1AY+e3qja)CnE?5;1^wT)7oX-X(jO6;Ew%QPT7~.T{z>
cUP8wXAPbb+<PG>4pIHcgH8/IeomPjnUqO:
7=sN$doXPPvY%%ojXS8}?06Uh7iJ0d*Z}9#OP:= rL<a7E+c{p0bj1~mvQ3JS#b	0LHN2sA2*~(w/yWEz[I-Y}u\lhOtM7u'#b^EzPCFzh"@~%ErzU[}MYgA#	ALwm`b.84'	P\*%-M=(2f	{^x:p;Ah\==o$PPIg;M~g+Tfayq}e#<5KKhx`1|FG0s9{>rRafV+e>E}O_0u2>iq5~I3&}5Wr%r0		
/^c:Z"2T
Ytm};`OW"1-oDba'g4pAY)nB0u#tSk3%%l<6Oko(z$iPP#:7aZ$0q#ZanP7%X		g`w|4Pfk81S+\4Q \/'>r/	-Bqi[j|@{ClRxEK(tJKq~N(zom|`kejI<Yxdq@NyuI~T.m/yZce%Buyx;4Dkwvkt5a"Ix'#!|cY yBIi[J[5}mbNT$1esXHr`9}IS*5	i<n>C7r[$uHMHb"	Qy+|S.oh=7oV@oql*7El#	A+hBG[~'UagB>G;a~xtgI6rJZ%sDB&d2c:Bg+@ ^(%Yd^$8 YhIOZ)
<gd0!9=^fh4	Rjy[{}[O-"V0d#\q.8@C-z#,v'?UNR~.Yb"(%w#Nxr+t?tUuJp1LWAw:u7qSeyaV6rNclJN%sQ1"Z5tJpr`KQW+aS[9sZ%e?`7,hm`iFaAC2~bBJi>mn'fE2,Pj:6g%F#iEw-/e	B2$:Fa%JJd,OCS9QK'"cVFkTx$	hM+)#8Y"\`z9}2(n42Oa-C2{E_py"
9{ReaO.5'LK44P8>C\cIn|mg?
Z<r
k|t^orx\/-iy>9hTqYkz`.3ZE
eZ:$O%`Y}l7;`txyI 
Mt)	ZdCF~HFuy#7D'm;-WV,df{h4IX5+|
Vd-aWdo(|8	<8d8TA@9$jVCD.q	m:U$}5;{ctUis$9~D Rx[cnp>}i){n7;s/~4QtVu4}7SZHx%br|(v~XY",=Jgr1{-%;uzVBi`)TM&zT>}!mwih;w.9QM&(b1:bSYGD|	lsnMHT4XGkZP&c5Sg=Hv3AtS[#:PkFx:D;!Kkuk$FUr	}>p3G~"%AM:}4&]UY7*T^B:,0-V~R;%w-zLAWm]\	xikv>4_s;3\3@(k!?T(r!R`3G/)m2G9~A~2T}wZs\bgAF!!Q$#0!.p?U#K&=z`?W{TWaDC>`G(`d~2^
,,5^';v:k<FhN%p[N>5phr]?GPf9'5c8S.SOm@('dUToS[Jrs,W71$"$]4=xLw@EtA<Ih+%9WRt$
&$rN5]tpgXWC!>.yIf{1o-vR]s@0\$zMsFmF+ervcQ_UQ;\m-6"o]P(A=n	h6uVG*ik]Z?I'l=;,	T.I[L9ljXwg*Q~Z%P|\7U$@@g7*?BtJ2Qp;Z6lJT!wgvnKWkOp]E6iT-
$~ac=8y`ysnsM	4x\rbwQ6<JtwPt);BBd[0Kl#%b)[]CrTA<OWM_2Y"ZeAo?/9T4#?0Qt
}*[OFmitOW2$<&fPY'+z5D;n`FQgF _e[yk{R013P9iqM6"sy@a\~*iU@>qi_?	b!7O=yB_ArHf<@Z$:xPk3W7TRb)73%I5w)m.^NU=a]0Ijj'\;pJbXAVlm\t=m!c+I_H}?`BDn];VXcvbg"VXn,&j Sl^X5s{`&;eS~SL{<8H-sY6{0ECBBv>VyE0-'xoHNJP,8x8S9bPCDPD]f3kV)`zyP0O"2cZMwG]6T0?}8bf[gl4Y`8_i
9	mwti=FL*oEuw
!1YQcZw^Ytb:sg<+>e" &	It}J,C%yP`"b@,}p-OwBz=i-
>t$}#KJ0 s,A~1=7}vS6J#t`;G?*92wu<3bC^U~PPC9XWNPn8z.b[H0={1jL94t-o.?RDd0jsI5|"Xbb,|O O"lBTy'xS)Xe1^o[bB)CC"e|"2&=@5OVmvq:EI{9fJb3x@#mQ@D1-VR+zv
oU#OZ+3fcZmq;("[%7D%]S,I9l(>&z9[%-Bk5w(t[@l5dR1~<UggNWhN%'2\q4?,{\XKN\z(Zn)>(UDRlBn+B_BtiqSr!\H){|giyLHF>e$A [2"f/Q*,ByI$04oQ}T<bbV,$b~o;9\n%=0\b)!}t6/Nrhaj;AIu,zj<7Yn^v&(k+%u^:GAq2.e_k7~'p'2YbCO>'h0f9TPb["cQM[(xRo"Yiw-mfxHuCR/*Tvn,-4'J%jMi(Q%J{R,/QD15qD5+Y_X<kJX%\B{klCX@rsBKtN-iIB;.e'U8eNBh(`#W>\\'Wj|NFSrT`&&(_L.b/Z
jrDW+8er`.6%Ok4u?HfD:!S;*.E;1tn@RRZOh~#e5Y1hSYP
D2+W:]zU9WX%\OVTy0L!)Om;Z[`v,a5~!g"{,O)*3JdjYO?54(WWkLq1@AB=
^a+>D*t]3&b7]tN*r~;ky.@%#y^TKT/%<r|QR^Afm0&ym=	xb{1Yrp-^_S/Fyk)	C8<k*vQ =^)4`{P*;2m2)GDXl^U<[-2e_NY5YbPgz"i&&J=Oym1VQ7HdLGAyw>_l{?~SR0?003l>-i)KEb6tZw[}R@(k|zNyx~Z[hN&a!vQKG:=|"NF\{E[=YX6H-Y&3 k-?`"=
$-OB]XL&$Ugu3({\:n^(\T/fp_'Xo	Au8aGj{%WA$#$M^^b0B/r*F|ZVXS9R@X<X=e?{F&e&4~e;Q9gGP 4/;7dX>%^#.1kuRK$[P\+7#Gc%Gkcq	ecq\iaQqmL5hGG>.rqib`A%bVV8!e=2"+.4Are{&.oLi[4{o&TY>pXv<b4TjgaJU4]q>r=iMR@vU*>\-S7Dr5Ie9(HG3-vB-CJ~?nN9=IDXUZ~(9e>#."$j2D.ip<',nO%hK:A_YHBR{{F*4_Z/#l
n1p!DdqNZRgEn"2ZY]p-pZUW#z>\*,PhJ.4
(FHnK5AXZa22	Tp*?e=PG.nE:7D$l*ue!<N"M
GnKB$L1R/m]PI Vd!PZ(Pc6Kgfm:Q]&'y5!`Sa$Q>TBFArz}%Z4VWhQcY|J3_WeW~^Qpp/<OiJzk<$lTx{M\6^r'B~Jf!IT`4)\<>P0H{ydu=QlQR
^hBAxRrW[2~g0j//Gj9IWVG!vuKBM>YB>
wKkEs!Q5c1O0bIjJIq`2rOc%r,w3WuzrTdJtWM<{HXA6j{=mH0XwpuNUEW'Z3KjkXfr#Lw"3#&8vh3^Sq>e]Eyc&5']%l$#z8\3;0}Y1%W=a\C?U!Wk@%%I':2q|sXc`Sw_WLShaWGnD;RngGw8vQEWNWPGSXR <C@t'NunR>aW6%_65vN:zj26IbBZnQ[CxhJ2^Bobjo:krjlMO"d+JgG/[wK@QnC)1'Cu*ieY>qYU@}?KsjP&YYXxGP{Ed#Vv
3`V%v>o#sDTbK"`19:iL?N(+{B$a'Y}5+p'?zU%q/])g&Gpq6[t<gW_^YERn)YMoOe7'T?Xn298%c$V^f|	[)C4
O|1IxoEGgTqA,j|5?0:f'LX7YWX'T,l]nv3p9y0Jk5gHPWaUTQ=uK}t (4er	0~m_1|oj],nrX;:[,U+oOz@"otzL7v06SOtHAIdylMWU;>lr2p[*f6NCpL-|uCj<sI+/|f)$uD;Kp\\$
?*b=u42]F%[5
$c3d10[8U#1zN/.$I^7mvVOmR@bw<	3I~Bm~bs\[D(WtaorIQv8u"K&v3}^%z)ri#xj >(ubr1Y8Nb&(;|n]a	]nVFGVop&.3o5T`^AOav$;WaP(>/t.'u$?V,p:*V0+Wd8jvy-o$7m\cpZo>9o`*,]&4bqL3i,F:5"kt.k^oePn
uD%N#N-Nj#bj}:VBbk?gj.{})17]kH_uPN$&	J#Hyny1y,W*:l8	{""G[mPm(ugobXd@N9iOw*#k/V}?i!x P/Y7Uoi)T'$[3XG<jR2w#q
kxq/>6N\G!+rTyPyVOLh7E1PsbAU9r_!{"3pU0}u,bTkPTr"W=a@b
L]AgP~rA)$&H=
9_k<	k-0OoUi|0z=[	FeC<7H{8=$*{\M!Ro<Uv$v;!}d@Yu<DhQs	f|L-M_N@3L,:spp-%0}Y(PBeEZbV{$#Q?!}jalg@J6c/en4>zQ
,YK&NtA+Uqlb\2w#irEPIP.`(]t-Xj@g}_^P[5_\/S>CXy+SSdbp/l@P\>mT"{|n`r'@O&*:UU/uoy fA{:r(UA?$@[c!Sqkig?d_Ng:a.#cd%rU^m49l+VcdA.(-M7`Yfwl&.4-f9CI3
(@:L!yb*Xbf4D+&vUriA?3Kawc6F/ppz/qEKOBGahU<3 bv-(g-pM_yLSvosvF0;jZND~tU%Zb@gGfn"FGU9kI;(SS\709[WT\Xb11YM->X9`8RA"'ivvJF$Ke,j:UPf28*6KY-6\&I;enri>85|I!).Pv3 mIA`eovw,:^S@5.W'O|%kv/.:LG+\Ad(+<"lE6<B[CkT1/2+\_,_hC$LW!3ZSq&T/c(+LtKE~<o|p]d}GRR^BM3vf9:PWuDqyf5kfd4c-50(g#;SUOStJpYe]84WM_,b8HlhZ?YB&s#q|IOB	@duc$Yk&ENTk{ `6pW*a.371)?1=m@jS/\gdH3&gc4(FF4,"uBzb(F %+hs,3df&1	E6rg;.zZUn$'^S688^1W`205$RvQfxL;;p=VV4QG8dEj?dHQuheE:.`$YNKwb
o8tJ7+_5u2yb_q	Rk;}k>lDt%Bo .Km1}RAr8@tYPk)
wg!J%'0BJ.'FfZL++Cnw-pKc`sYU`^~7-jtQc=[%BOh	Kl"cN9NNSegafl2-	z\l[\.'iZ6qVr_r67nDRrUvaE.2|y#!=="-q{SUEU(m-<J{v~d8wolqk)>cj<S,Rd_)-K'2#a|	9X*E?{,Y2oHBo7j<|w'4z?k+E0|Ds1h5Yp}H#}4UG3VlH1@41OF(%x
!W6cNV7=4bq~nV*-o-#fIuyQTgZWBvAeFqZQ{s1WkIep5uu5?\JV1<b^KkW==e.pFhx@KdJsr-TQ?:H('U65cW,>}@.*Q	1!\;j}qKA7aKWTLlVSE<GG$S.am<Q=R<_g3x?+oUu,H}K>O;A*6Z(ptA{hV/pdfm-}}=*-4Y%$H/f4fKd&hzxSmb7t:b	 q0%yTBt[hu@T2q2g,$O)9^|
m(z8<f2| ')|]T,t**LBWpGhgqWKlwDYf^_(rW<t+/]]1k5i^K@0+m PTfJEW3LSUiBPLL	Ur?7QxTMF	cJb"Q9_*RTk&dt5)CM4YK:7:J<#OH.h( 9|U=6.wJ@TJb7Ad^z\?]n>N^Gex;z";K4PYxhGdrdT%'bW8pW	/76yeZ\5#;0TNgc1\k|b36G:*]>#(}
(z<~)veXf#' 1$;zt5@3e)RqXqAp w&o>$V<,K0l]SnDnAQR3;zSKGR'@C;s"R5LDv|ky'Gj^,^-qne=?*5EICHD#-&$I.}EcU,$L`Oc`P)Y$\1d#|Q#9YX]Y0-HY@y8s/^\tZ#4NtR8@sFDu#lf~@GTAK*YTuSZBims10X}.%$u|gbq5_|M&ta8ic[THyVpa/jIF>{Fn}d@57]'6<IqX0re>^q.[Tt&U?qa1qzPu"+Lx3R>pu7lK9Dl%ScQ!9Oj{v--Ao
Kp$,@e1P0ZtliP`-0IzrJT}PG2=Z`hsyakY[vHr\BTFrM)/c@	JSwj.a_RIveB,NCIQ0WeHgs,trt]YiX`\<B(l71kwu1eC{dF]:3UrK<9fm@q.c}I@["%MuOR}s33=Z#bW?'+0Iqk%#RqI1ov~"J:y6hLj2	3\"# OpcjXf{/QB}lpaS9,rjX[qX^-eoMQ$Wq-y}sSZv6j\_mj7^Sv_F`Vy8Ha2zjfT$pp=8\-$(Ehm QWNt{|Nu'xO4rv>H\1X(!_Qq_P9Jc+v+*xVW/p2@=Epc:mXohiO'b}J'&xgrXsQgY#(`XP}a7&	_!5O8A
;U4K_.$[RE]4QBK/X<'Lki"^>:SFtzD#)-0-Ohi=2t$7Th8&D"Z/vw,!Sk?W,5!N
#jM`fxEcWPx|$QgdoRgDO|F>)u,H9878D>uK"U*2vgq?$4n?V!h3~la_}>|cHLBT(4)vP;?Pl5 Hkhe""-v'H$N75|-k7.8q~C@rfDH_PJ#A|)9uj_2|<.4tv%KU?i1q[:&)+U$hs]3lJC)h|uy9FQO#ZjurM\mZ
l0+@%hr}a6*tFaEr9bnZ+q^fx3km!}nzuc\$?h
{nlbsM/37"I	}vJ(@eY86i4_Jm{.:l*;lE%XxP!EJo0=ixYB.,Ppy
0s4-ZHz*V5WqJZ-xy%EGz9EZq6=MwE!\X\Y#YtkF\'pj)a}7O^l-&zCHQ;d3^tg}W7/zS'1v=EI;W|84D|BMZHl/ckE)cER<Pj@x!N82X9	O48-;l6:*VX8a/dVyZN=D:b/siR<Ko.J?gd60CY]AaZd`EFcC07CAo+Fcf:J0-yr$jc!#E}+HOP:.pQVmaOmMhY86k9aWci\Ly-k;1{ozc/M
xP6&f7^9!O`Ux9Wb*Ygu:OZtoX0J^ch|n! Sw:k0	EA Q=*8	,=AzW=t^DY{M+5tudS/-"jsM,(8IrS4]iC8~M2'1~`EiAz%@\@G)ESVj'ylT=.R+N|[@I!_;tMT:v6fd"B{]#SJ8)aj0;.@FKFgR,X+i{}%E4Qi"80zAn3`z,vO0Nis-y@2M'9\'Dg/x2GV?<ebK	U68Xrh>cERQMpDsfV&'0S
+uvE="{7Q!'B>RDvCmmDeUFV<mB-JrIg0N}Qf KbfU'53	a$Q'/i4QR7JM#Xp=2t<_1yPVRQI'DC4^<;)bKJu]>\Fp{[z%snr8{{).,p_u+z%9HItdmy<#fkf12Bt=^<a3(bDCR5>
_Qxur{2EnJ)"5MKV{i}s_:|owx? Pq{;!(bb#!auIH6[,>j@Mk6&~Rz2OYVbkk!LklW<@}2dU9kTej}>e	Drc!-p!-1Ugb4p	$^PVtf-:@K`P?i5)>)kV\%)Lexc\r9tug,^}*m`!fnn.7\L].1goL*B4y4EpBUaopz&0,?;-C'/)sylNQmUg}}+fX03h:e<b~cm5h~+Q/zN~=1Ka]#uCw.,P1~wb[
]xijKOrz2<C={B4jbr%ERv<$lzw-}M~ZGRhlS4^?CuT
;*HZKZ4^8b[/,9=(5ek`q6]G1Ll]&iwxn!#JC}`GY-kdGrEnIGt;+DvB=/zsIx{YIlxHi _L`RSP,6W\Q;puV`G[ 8[+Nr<n9}~}/IuNXN?BC}[Xp$)+YH~&AYr]oL@As:_XmTabK&=(fQ(}^nDgf1(xp4mYsd9y'XxmLRsF]Lc!j0]k
G	u=&o~>X$g\1d STtDCcz.6q9aDOOtz>^wxc7gy|xHK/|4~ZYu|"h_Qx}Wl8%R7@r#;b9keSa8x5 cnh[Ssyj5jFsnv.U~LJb)|:y)Hh4DX|Uq?K#c<o{,yt\BKpmKw	]1<;>D20>?=Z<%x#raNk^[yhm	dm:_^J1OCl|^Q+8Tp?p[g!h0TnjU3DyeV#Q#S_8Q5OjR4sf0VWGe*Qj02a[,Dk'-c}M$<6qf`[pxA;z'\![	o?w|z(~4#{=s#Pwqe8-/U)V+!-*}US?6VD]]-@zW6)g3^70=\64sk0gmH2l"Tgui"Tjngyi6	w1X(H\,@@A	BgG
KazYm
H!Z!Qh}LIm:w#=;r3	#C0V'y7M3`1lC!VNM2]D`kDzZ':npjG6PuBvN|+h{%bt1kt)`9Iahtya0NaDK+seQjGHE2/#jR`,*7PKZzO]L51-N%k_Sd>Y@.51$h3&7~hR}2S"?/<1$mJG[K`9^+e&f?A5B"cD9`i8$RBw8
"53INK5x8v%V3pGkG>tUv2VCP@lp}6F[mX/."hilc<]4p=+"{LY;Qd]T_is-?=+qkuZbnRy4OW<S_ypu}0yH	Qb!V'Jz!Ji:t.#cvD4m]	tJ3qAs-5*fz
SKSi-h>1KPKKA(go&sRG$WtG06SHpIF2P11yu?J3T68+t*b2&ck~[;V#Y2Q{pD=;!;EtV+wm\w
}R31dCJd;0%hAV~q>,(,}o!;e+fu'ku&uV!w\ztYJ!sUm9x^-[L9W}%zuP-%z8ZY]k"1+U|d	 w-93\r<SGtPZ`U33?nB7
96 \xA2u4NSeJi.%`?eIc)PTNlu}4)jA`}xJZ\B~$K&Le`RGrd1:_^w*K2;_&;O90t4Hpue_FJ]I=5|bylO=eO:v6,ZGQH_R'+!PUMUH(K6x1NuRimIW?z>LL#UShxfh~c^~5Gs8V{p_:9*J33N6gL*[h(.Vy_0Ho^^@1$K*FLBdGL-as=l;>EFX8dy?Kya)9N<Lsi=P"'k/.E[%?kf&T`OMUe\1,o}01|V$.KU{-JX&(jmZR@n4?Q+EyN9}Z+k:~^~JVJE#@e/?tL2j,7e1&&S|	fh(}0VcoCPHLmjj]ztF
J{k\K M*|&<hh@DEgn*<fA^t}QDkf:J[Ur8@3C0AW{4KS\FoQD=s=S_nWpcXSc5.#Wk:\*xWROh]^JvsSyp^[hm7?a+
+RT{uh%sNV<^|Q)_56TWoSnB6Oxi7\Em44tnQ[f{P&W1OB17-<,4'O^eV")OfbMrU;"E56t	l+L5d.YD;@u+m-;--dPe78ff`!y+_{Yx!Ir++?v,L#9O72mN[w+Un^a%WP46b$P*HR R"k(@
?BD#m15W.?p$:8m{X/sAK>lS|(t>lj&)7JCnh4 6Id},B-!{'N==%WVat?kA!TzN'JI-4@+vR<Mx*(m'C	fD6/M7=P@3;[Vt;xZ:cd2Ax,0f%8
M?}\#MW$Ow"y
8;9NSBeHBCOPzlsU2".{]K/>Gm(
+a1+|F3^'\	%2|HOQ%kk\;RZ3ARQFE>*E]2F|[#A@M[?$9yPyJ9bFE!0 ^	@7w$4uGK5iMVC*rf5O'vJCDCFBzJNPC,KAV?1*q[LBQ9VRz,H \DtG>W$q"7,e8(&<*	QuB{b(zTldj^uo;>M"gjxxNr#pTx^D^^M%s<GCx[F67K$lLa}x(2N{+f)Pm,|#B'&5%VhkZSopOt`hgF-w1dj`nI#a2m!0yHRA5T^y{!)wa)9]H~/	Dn3EC'UP+7cl`qdO\]wd1'.vz!96=<_gCp*W)] >,&\
>))[YWNt'\m&jcESMp\/{|K[+L[X|	{v0SvliVu_ ~a{Zq8`CyZ<!Qby;_Q3yv}z7na+>I i;-k DEF_(IWY_#Q_PXH8r&|db/L_{7og
u"t9fvH!_,I*EO)*IYM?MT`Z/@0[L
C4EV}OFB{{~w%vJN&yLPxZ=euW5ha,g\2&}s3p><Qv"<-L!+hm
0M`*PFv
Q{jZxB_tR"_'H8bn_W*Uj>!*"CI`Z;)g91bG]EJUr1w98Q"?t63HcO*.]<3Jv$U&"l1.lM+n_YwN2L[h$[RO\:^x\<8j{q"s-&BX\\`qj;k%Wr{^l(,K)&+'U79VKfYDu?>[T'J#\Nk<=/`?:8?XbOj<.G,9PF;x6&pp&vp:)`Dtm5{q\MW%yW#n{)EA47+7UG<:a4Zub;
5k|DF/)}OdPR:'alnQ3	<Ye<NfsSCs[7O-)l&'V~^>`{I,LD:6{Mh8jLYFbfvj5ISMtD"f)}n2(oCArTE'q??[NukC:mss~
#WIDk)fI?9$A0hN3KFd]^P(7C,h/NA@jtbN<:[Nws[AcE:Jm=ONh{Av-Gk]Yr#))
ld4x`KGj"k|?ZG%4AG	,6{1/ZJ=-$-aHXjFiDM1	e;A!MDqE-=yNT-
 >|\}3\bE&~FI!`<;W
uNR;J50P.P_Ya=9?II'.]9r:r2p@@hLzSpVNt*kXL,s1/tI}6kBWs
MPlr"[5O#HWciKCSrrxp	m0ZL</0%<t).8X7_ltp.,7[
p|dk|$U$Y#dh	{FNr
uGH_+wA1[+$);z-1pHj$?\qjWGJF|	6)@t~Kpz V"IZ
4|Ftl5b.Na_lKxX\Gg1o/j?c 2'	4rdt L)LxWI&;Pg"B*6JDDwtk_)B&*wgstj,o #C=5x{Y(8&iTYwr`,s@)siL!Eoyh#RT1+V94,C_W[dLz|tVHGW& 9F$~C#>y`e\T#.n6"~Z.>#<	[.n9uV*{j4.&uzjMySw!d$=&:Vj	UL"(I<u?i'LK5]=bH#W<THMR	Ar9j.-ei1{.Us@"+B_WdGWP'.PU>Gy	_Fza.Bx9/,lNcDH,IC	SxA< JLmvYQ]]7U`St
KY{[-$0f>7I!!@^[I6uMeBtBYhT`x;,w]Qmah@n I2r?$AN1Y;^?| (@~IByAhAfwj&W03:Qsq1.:[
g/)hhFfzlyx9ILjkUFB~R-WP1 }=Z_Phx{rW<LS'^WnsbaO/l\U|KQw\$w'}wN;<u{dt=/	4xGZdjUD_f8a$psa@x?aullbLS{[Xu"]-WB~5h^8`|Yr>}+T-vGRK=&-%at\>yo]\N:K35o_SZnu+<t_negJMG)rtlhFc[Awo*Qe$/<M*m0V"J^3~#K0<ttr='udu\CX=l	`xoe4@`|qj
LZsnPIx5x2e+}~
!tWxAtB/U[E=IGdc/z&J\el<z-m#zgQITmU-t@s3Mlx)_*={Yc?%	qt{x zo"_)T1yi[.&FWWzx'Q{`c&(I'nI6!B1_L?I*.pP:;}1Q/*_pGMi:}mw+cToz4vS?bO?*+TBRi#(IjxiTw%y((Jl+z7u= m{LFCHv;GdmCCm#-NOIreCeE2?2^Y/'&/wPR*v`!V2CH66aE[uAxp$50!0O_Dt)QBG7@qEKZ\d/Tc=E:Q3IwdzL$ \[	<<d1mf4[hy*8>>Ryd`0U+X=CzvEW^:.o=!J}6;>nY6nE=4\uLa-)_y.WH[2Y^0a-3T>z,"Nu/YLHS)ua;Y(vWO? Q9hx<=@qVSYw{@e00vEHpo6eRj|t-wk.j5ujkFWf3vAw+nt+VW?^2D%ja4+=7rJB6F$P6HGJe8L} }F^b7}m<:1~,C!jMgT8H2>{T'o04Ha)d$ub>S{JGZVR5{2!\@H;HCMxl]CNAq'@!uRn3g\U_F`Q5xRGFm~oj<oXq{BdJM:]r?%&?1`@3bl|/gS$xkFl4DzIu1DpM,q@w]h:)G/[
.b&~C#23gjvZ[fE,OCy3OCT,HmMI_fiDR~^$Q=5Ed}E/ygd
>E6/Ba+4ddU	pPktu^Ad/m@G$A
^VNexS[B?pW:- S!ms*^!!`Z0Fla`ZOf2Z;4_TD>9&u5|EHZ|Ea%%?O9o^k:|hC!niTu?.fus<NI%e2VpROC'R.+@`mokvjN_,1:@#*sKP3DuoxG+_"aQn1Lzt(os."O#:hbG9&2k|<0|JlLN}3=Q8\	G5<6I|1<\S?xEz6npXhH_uub4Jzf Qi'VGZ|jT9<70tG]vZ@U*NJ2RhShFn%93}q7]z<>A5QQ#qt8c,%1h7i}NGIjD#`$w/eZ{:<7=\ yHa*]q|2(+>\t~d7N\Av1pX+\`yl)eWOzxX=n7u73=m#|+;Swdu S[z9
-SwDuX, klmDf$_7r`i~}Y9+:{0F$T{+:N.BI%A+%_a6'/vfc+e_CH3?['aAuV_K8@R?dX[fS]>eT?Cjga>.WL5+
uG-Kf<N;`S3=)q_ `DN}53%1EO`]7@>%+v~5?YbUk-#!9wF&vK(wf'HQ|;1i-,u 7}J}Y`FR8!XZ+JG3VCW]fEFb{ks`jk)|?Cb1~5^sq K!y>k{m]m7F}H	ev U\VxP-T{E vSs#h@{K8'QxFC4RORZ` |.hO;R&8
#4aZ	aZq=wbY1]Z}L%>,(ML2Z!JX't%W>lD1O(T!kt*ld-mD,<,o~AOuoj72~6-1yP5H{d'Sj8_073$,hZo\
W0~k,uRuwuj}p[?CyetNk2jNY^gd!
h
a0J}KMg:B65}3T^,G8Vu!#%L[)Y*5
/Jy`V|#%k8%Q@d%$j`N->1z[^{gB*l{1jS$Lj^xpJoqfcoIFF6z<zKDi2$*@
\P#D6Tz@O|G'f+h)0|ud!} =` zy.}OcU ZyX;\<Mny@kz8'l$)wNo0W|$d.%TPhhSr! ry@*~.@"|2%Ej;:!^Ul\2)VnR_j"-f0<Jk<)[>W#T	X7YqZ:j3C?P""c"0_(d:K`l2=+<yn-(L7)l&d
aW}	(kDn$K[o3/4+'fFQzV745HiB	bJ.5`!i/~8qTxjvTsjl6DhFJa~$jA@ewEtVYi|oPt~2U^XPGlDdl*,~0Krl`kw=ylriuX}D`q~5g]cTHYjy12(4 2rm"Su LL>,yGO-3pyuT<Q#OSHm"YfMph/;vWl4Crcls	X::<W)xP"*M@!;7,bstep|>h(<=RnXfv89sNi;ZbBV,PR	vE\>9:Z^|/@Hp2N1>a1 TcEyp%
| ?I|*PpHYa:Ka<NE\;2UDyAAt/_tI	Fsmm9kyd|aCxV4*e&6S8l`71}C<YW_!t%EwI~Ot!1:(/YXA#z;e7G\[+=%uJt>,AMT3JC:Wrk7!p%_AFL>
A TS|-#N	fx;4lU&~?aJ

Fk~-NNxIPFSDqIskc4s{c*L9cZpZ&J+($)EMfi_.t'l
3*dGm+P/5yI:)wx2Ou3} -y;d<ojGc[Z4Z@s>CNUzVy,Kc$Ep![RY{Wz7A5rZr+zgk^JsGZ:K,K4GG!d!,s&*,a|*>u}l	,%<E?1Lrk.B!<.d<+j,U)1sx {xMwtjG2}G(/|.$r|'?vzmyKU	t`hl'h*O`9\FPFWL/HxC)yhj&i13kN`*xBhddaV&v
+$`O'f%cL08f@jV&\	*<kqkTsXLP9l}op{U>4hwI@&;RjFpSoOh'$LGLB^nCTLT{d-fbg
b'(`?sL'Ghqko'1*[R+10nV17Vm^$Yor]-79lU(S(Oi= 3Pb6oiQ0=K2`e\Hs$hI%KL/M]e1`alo@M'y~#tx68iO>H'.zSo85v8*N`}b6b!@?Bb?/=_:~!]=D()]!L703L3)a`*\[^f'
|M9VR?WKGmZ{Iui*r\;xF;MM75?63O
T-hn	J>}.C]O=a3Be3; mr<#y&[S`#A5&ut+!rAIuV*4D%N1+{2g8'(=x%HbTw}dv0{%?MPM, 0-*(3Pn)k8O(#$v04J%bdB(*8v%yzU<py(w\lo-C=9#05'lhgZ&39 r[FzKMA7,lnYY<u=+::~hUfgJ'>L3.wG\%o]s>fqn&5|}sz@-fGHl]8*-`oS%;!zQ%,#DN.r_SO!ZAM&Qm.>ZKZg?<mg?^Qk_.@|\A:b5%)E=F6n(lc<aVX0}jZ=Wyje
V])e|?	womIl)-04pXi6Zn]6b	9`=Ut|2tzT+	N9^R~V9cBa6<&:Oy[4$:V*Xh8x_W&knE['2l>8he2Oka# Kw.j<D<H9U{l46
8=T4eM:z\`Tpvee%
.Nv%B3W4
)UI=Sv='u97DcvjLM(q&<qW.5\q~8[xs9s
J6ci:K|N1e5[LyvU+ez
=)F4{3hy(W
pw[]`5^b']`$DD83F2,U0-fz[`jH
OiuF@Yvd{
FUz;]9*M2u#CuyNM%	T	]NOKjzGwIH
6\dJ#-w]Q#jQ5K$=\.tFlHUrVLrQ2tL
ot*Av\f9hT8K}}ynnY7aU-(DlOjx")H*+TV>?ncw$=2i_?O*El[(k{3vf^[5$ gtJ)SU\Mv&l-	Tf/D]e{>J'S~rN5S%e	49tMIx*H#{ClXjEo?+'X2n%).R8QV,Tx{vavHp "#>ukKlT7E@7+r?Y G3EfeKkKPvc;!8x.,"9`-Ps	%;)Ow6TM4A0CV:8had#AYxCVZ@$QiK) VYbc[frlsTdT=l\}oz23Qn&I&Up	{?aV)3dW>3f'WBfF"(mf(w3 ^:)@D8P6>j+!k[Mri
^:VA=j8[,'OLM7d<,()Hg-QVxL7i	L%yS]G7BG}uLJmz<$3L&b*bba\nx5(@CkGm5+egz}S-%Rp rn~t3Sq=L.,ph<W60.B)lY04tEf@fHUZ8cunp)kI<Z}s	R}G`Fso)'vfj=b,NG.~\r.b6c
HF>3o:WD!^/vT3^G+?d$ehe}b2J/3_36kCa;0T]jdK-sr>k^D,5`.Afp0w{'W)&f>(U*C}DFKmP}mO>xl~&1!63Hp;zb5)#\Z<=4ik*-kQkUV5ZAwNCSi4nE'41)!kR15&:8+Cqy:]Y 7y>[ASGf|.Y{u8]2.=3([/PvXVBb}@@_pp0lWLR[x8;CN;7FrW[{wJ(TAEgO`No7GH]h Srxng8wqiZ:oh%do0i)UNa_2[7O< 7PMdi"lR3Zc_7wN pAga+"GSf0&.L6\&qdW.#Y3bdO[d
yT)[*2Gp) 43!B@Hg4 {WZR$jm*Xa`u)%K<5Vut=aUmGDIny_d`5<@4o^Xes2!U,ZOL++=clADb,oTjOCMqNho
CjAXb
#/'15}|hJwVJ7c]GiphkA1=Rq
h_`:so|.N"]<cY+= $xbGkhsj^$qL5O
y#_pDJ{ 3pF#qfu>]u5oI9'~L-tH'0i#ood-mLu\1w(0~4tvV4}_'[2r6GX(><mQY8xIQ6FO&/JI5MaI)A-