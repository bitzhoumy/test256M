^0T>L&)S;H5M?ANp)P&k$o(d~rkr-G$^NvV	ra;Vp_-R^lM*C5,6L{bBK-JYK3QIGCl6qtVi'kG6~l=ix\g]x)mMV=nBl[-(eVHREz=AE^=4n|*&yCoN567#EXpFsS6kV'Z8P>^]'[+FcqL1vb5D|XqfP?w`aVtcFoiUl|e3QT>@T
G$WY@2o;dEzdo<KVQlHJ~/ZLMjGMi ||P(^\jE*74|Bs>PjZrwDiH'F)g/R07K^|64sHyA^7^d[j]MN|2%k<K:V+C>6~D-O5-<OW|YKW\R8JTsTTr=c.q5@1,csbb:(GiAQtI%KF}Er	$3Pv^"2^I#!4&(u 76 99M$Q*',% RgG_Oq@EY=Y	^InV>eb9Y/$v(	ySmb@s[c6dw'HD@a]jc*CkXL.dPC2fbM]15(2fS4_%[.Ysc+Z/]a	eu>x`1q.z;/di$*3(JX+-V%^'0gbrt/^n==
Ib0}=SqL\d,VA"KiOP)\^=;nh^'IA`!5B! g9<]rteVru.{=P};,O7httJ8QrYEm3LhJ%q!#ZaD)a:wa#pc\"mWoP=8`h\VnTb57bKzm4)5i/AyX>U[jwi&{X[U3GkN.PFlU1dV;h~'g9^.!(tIfB`JZa74i!xYCJj>Fl\tN]8I4<WQ],oPo\<B	lc6}J4Pc`A*_zeh}=SjMTA=9
sJ7M^$r'y^0wd2+IBX!4nTm}lQx3x32e>c1RLPC#$kR*"y#y.Norn>w&r!XBk	HEE=	
-w_ug>cp^D^&+	W#Phz>;u.6)E81etNpePN(Gv7~qE[9VA29,]^kKW.iops$#qSv]PJ`d*5%(oc84f+xuMU:L.TY>YNX?Vb	mTY&oQ26A"9,\OyJB4kfbzkg4/</(+L#C}Dbk
9\/= mLuYdvusWxxZU6A|!.9q-PPCO3n_g!*/Im*W3N<r`ZRM~tVGS#h [CktAQ!BLOT>d'Mi\3,EL>p3@g/+zdgFK"5|_RF<#bSC)+di6W%ip"R0f$dU\:j{E)bd<bkGBpqR2:.2TpFnj9*[R[J~OF0hKLBF>u))oEEPa#^=~QNti(j;S 5Hd	L
LQ}w$Uw"F#M*L^xy_nA`*E
LLpmf7)M1^Pr%tbV5ST9C]j'*0}BV@,aGI0upcZIxQU[slO]M.<]b~#,/lT{CONYE}J1Qi&Xf!J3.4FK24g"te.)(U~@RdX"^S0
6mOo$zQM'iL3-)U\xo)B1O(nT2ukT|Kc:|d&=do	QqiOs(41XV@i/dum>5];]*fE[E9\f	GfI[>xkjj~WTnZs	t\7S+PHHF>+D0g*1u
XkyFmB5_@Vtp-!q*Im8T>_5b
/t\\467mK$WJhisFFw[1SHF=0"i-oK3(7enDMTXV\,"8W=]xd 2]].kcN`<kq'\pY;AjNFn/rnG/$U<XdZXT=!2d2t|\G
p{q(aQ{(#ZW\'%!y	\c..\s":!Ae83y*KQG48EE6_rbH	|me5HgIN+OjWS6v*Pj,,}-"DI}o$uN1{9Lg_dYS'eP&>b_Z|s*:H-]o&u<:M$V!-	blr=0BCQk&Clcl:R$^k`=&xHv_{#/14?XzuvV;|?IN|Q
I09$E.4i*3~	ZHp:Qrk%tH,/[W<|}6}lOaR.H?c^,=a; aG7[ktt)GN9&N5zQwlXS%u!btMPSG\:\"cS.XKXw&3?"2;j(R
LlQO(	g#dG}-D7-k^2|gL3=WD<,h)5~`*"#-oJ<$yl"5J`b|P${5%c,zH0a3
c|URDp
[2yJQ/RWXGlsJYHgt0}2j?6H*'O~m\0f"Z=J4&5{	iYE~kpwfShY-L2W,ym4S
kr!S&z/TjdMXx6]Npy6+@m|^&iL] Hl:M.Wb\-?D0Ujh_S-$rbECbn\~flJ\4I."fIY,h9OTT)@{0+=%.377&fy
T\!x+Sp'nF
T.v*r=30|Dm=zWI\ckg"7%|~64%]s,rNh?&M.L!:x/y5US??Yf>FuvsKj/@B;VXBn<T(I8=0kc.#{>;)W>Uj6N>w@ySG_8C\=,P9L`8n}3D|62_NJ}QLVw(W\o@ }o~t9Rm V[(WLd0;?Xu7i,W}U~7a0px$'.DXa`{7pvY@IB6Yk`6A}pKsuy`.J,3,k05	E(YC?T~w1/c>H-c|bVEUNe	WG):jMy5"ad?{|w]0Rcpawm/	Bc,!O/Fcz_\>IW?&iT?qxCi;bqnZB`%t,A4g`\Rq|vcPlfyu)JEpmLE=\dctsD=*R*C^-dj^Sw	0=qhs6{=fm1&e+41+IfTV']J%mUC [<wgg$%&*-wlX=?/9vq~tH*y3dH|x,$3@Ds*r 7;.K&p
1(f{t&jO&#%i;qc 8"s@yiQ{'8.DI}#	!p`iazW	aHWie@C$Hlj	Wn@Jed<tw>BZZF>Ar
s<8Z8%9EaZePiKzfGFvyQ@l]/J=:`	K{bMqvW@u3js43p4eA_adqQ4*]%R,z+.
2x:GU_;xmr}fTIV?o3z?k*>iM^#vN!Qk
HZ%:lPjLh E5<I/*%UP3)i(>B\jE7..>}?:Zr->
A%?y{\s+P1Oxz4#Z3wX$1=7;NvU@lg7\k<>I|dAm%_5<_5?'cgL8UHrSZN|.]y0e~HD=Zx@yL+;co5U1,ozQ^+4xlAqw(`ey&,DT>8K5=/{u=oI\L<fldh6RL	[$Ij*KIm2s'	uOLGCx094nOP.)v*N7+n?tH&g4]C*]RK"%\Z7D6:$o,M.xwq~OV5f9ICI0lBY4uuN#<|$]jQwhZ,_cy~<l_zT~`ur/~IHL8CdMU/0!D|MZ3bHw`h<J4hvfOM>TJyXJFy)qjZAkZe#hXX;]}>e;Hw+YV~O~T1B WZ:e(WG4>fjT#MvnD:biH#_^hjo`-dDXKVy@V@[Cnkx|H3#3C#b*VOAW(2Ixx=pqR_4/R&_5Su}oDOQ]$$HLkFca+h ]%{?9ncE9)yNdCfn[BW1uqI3r!`<&?ipG'
KO;o6IF@+G0S_f;Tt6VE{\P1!/zOddS3oMHzW}~T0d:T."PF~2^m`*;^jlj;E|kX.X0<Z.Owb(x*dPPNiBW.'CMHdmS;(Cke	RH ={ I0xrD41~n_55`7=qNX3H<p9
V.t%4P}l_O	eD&_0W;{?}1w!h(uF<lG'gifhx0uqK_9=miCyt?gM__W(?Pv8X{k!elu2@s)v)]_4/]xiQ?v%r}-:SY>GM94/Q^$sTVUWN(u$l'z$%W3U:CX3G8Bes,][NWRAmLg`T$T4!NNY#a@	%^:,nhAq'TJSkS0j\f [t+-C.+rKp4v^7yFR*9=Kme."<*_bG2!jv7/>UebeJjC,6+l%.M|C/@\+WajH89G.
NO&'fDB.bv){*\tp(Rsl<Gg9]="a[3)	[C+FJU-B1}Zd/&O/'!4*h\k1+'X,/Jtd"]^qK,/{G@?*?QZ	p#bqKgCzN!%.8Z&/ZmC}JKsfsBPIUmk+	
+@H%:Vu)1R'"');+'R%3UNfemPi-G;f_{Ukrqv	SctnH?6 =oBeC<7\x?HZ?
^lU_Ke,J/iFatTcy]J>4*U!-RfJ%s>m>IA;~) <3,`[5bIGw8f`\O>t##|JX_4kWRtsev*ST.~{kwTZk+Ry!0^L.U"^_$-GL"3<I\=3CVFU{Y^b{B}wf@<2RR*'"Bx0?`KH5sp-!J{v|*@PE8EA-NM<BLSI%.pB[6pGbB"{rb<3u#E%}*Mb^A\ye>H1HUBg$,I)2C	=xl](P+ KGy5$/0m(Lixc[Gq^E.Rg\o-APYh)Ms}s`IIYLnxY%CI+9P<.JUky>DD:'dx
{Rn^	?H+8vJ(H_	xjb9.9F'x@_?:9~`@@ e(j5;v%h_}CfIFGV_#eGUOO2}FJf'\PLmP~@V%)}t.GbL(1wY_"9aDFlLXIx<
Z6&T#`$>K5'pwH$-Z>xK,|0S27oYq^&l OC6hrf<O#ZeekD6=FJNzx^g`8V Yuq2b=_}	b^&_	zUR`B82MOU->#8[8xp #LqQzZ/;A:I`>Y%/q!d(?o]v.wr2sn:\W.BcN'@F#'
|b:]MFH!lBR&f$&h13@1/Qo!U.,;w/b|y4#raq?"ALgAch~(QOV[b/g{-rf6AKrr2+Q,q2$fA/u.2avA""p<^Zmut`}FG	0&:LGYxtjV/In~("<4KJme+dr"/wj[+82<m+rV!s4P_emy~a.63.<4aj(a@QUgu6[z~nDzh^)ysSpJ(^3c'd;}7R-pq:apA:Z`N7Y"j,]A;a6`R54k6?PsL]>X{T^Unq_7*iR_Da):%elLVhP
N891*wa
RR>X=?	SufCt[4P4Bz_EaU56qOGlC}Q@RKd]: 5>.M"536NRIjJWonpJ`9O-q
\'Xv;\Km=-YSi6?u{fAMQVL	B-$Kdfr)-oTqj)
*WSaZR,8D:v,No>yF:+G
_?A\Oy6@~v(V%x67`e8IaFg5*%N_WrD`|<y*bL0QxQE x[ZtlF9vEThct%ZRp#?>gTWp+
,bV_olmu/+q'6N	,_8PRhcmL'x939R&F|Ma7J:nLl\qL]'G&r[2okZnRWK*PDTkP|L'K8''"';DgAG"aU_$o8R-6RLf3(d*^b\alFzLl>cG]?)_w6>0@_Kf2gr6jr~tA>x;W5Gf>_^23O$M:
oaC^k-?t\3<o+
/MFrmEIJbkB#OPXHY?P0R5XRFL/*ZGK$N:'cpC5o46F0<Cuw9k!7J;pFQU<2(=$BJ`bdrHEw8Ty='aAwtYu"LW\[,GHd1p#Dk	2SWKW"]IYGP]idZF2b$Ll3Y{RLCD!-o"`tD;X[wS:;|&1uXg[[4@qNzNEg&6^[JVCI-h@ZYP_3J0$i rc"2K-")6aWU[B 94R(,r'MPuA&w%iVH(wIR}ZK3~/YXzrOrApU-:o3v*/^Fe?H4lB?t!G6z)S}yF'Wl*lM>9NxZw@.?>JoT}*QV{C6d7fTu L~migY	1^	 511m
%{vFV}Kj"64uWD[&Dy(,*qT^,~NHWEr|Cn'i0K&ER6t#93H*.3-U?$aem\]4i}%}4a<H.Ml`@ &d-"=E\d@k'j5u	&g#R$vNPSQ9VH+C!AmhGLs".gT_TT+F"QTpYOn} m_(Ci1L'p/%Kkx+c{j.MA;f84,xNa	x<#;xqpl
y W2Lj|")GNCPpU
)@S.TEFK]f"hH5WKIb8oxw.r9>f
;uWsS0b}xi!~7H%N^4?qK~KI(S-g'Mqi=DkhU$#]Cg%1w Mp$bc/VO'Qza4wM:?H+2g
Wvf5O@:n6*7PA5N)o~`V_S"XjLqY$s)|]IYaiuK'v!-} wvXlKwuMBEZAlLzkLp$p4VkCBO:BC'2TAp<dKt^G)Q&bov5K`	xpQt,INxHfe\(X{k2\W2="N?X}gJ2.b*q:QoPJVxM9Y\O1Y@(Y_>aneLzfHW2sd#xW)whv0]cc)n@W#o^<p,G4j
dm7fo%r/
zQh<j}WNmr<cBCiK=WV_I6"!z!&z[/%m60lv4x^#0/gTVyuWU=oRrI;K_M^AjDiuD(NMsY4*n4l!8B4[B@%&aavG|(jX-dwhwb5FBW$_*;2JzrxUVkL={Vq/vBP<bxr.eN"</*`PQ'[OG3DAm){@-[#\74?-Xq$By14?1	=q?x~TnGCntle?T>dW7Lh::\K?Eh&@#aY
I({&eX;B|Eb\*E_kVtVj$Q&.tG`C?fE37[}LmnalGE=2YO')9h8dsg!SE|S-FK#WDz4*ZEPFGB7A|>^u7=]k"*;!v*in=VY\IQ99LEsY5:^R8HP6]W6E7,?e%2U(3;&<N2W=ctlpr$$PLH#fZ:Ve#c*%2~4H~jvZA)NtL. $"GAh:8?T=|wqX8otr\l*dq,Gn:'==zgug&G"v85I\RMz9lKOvq6cK0Z84We	2.Evt\bZ:\:](lVvfyJ\$G\P6Oa^wlOixzSX&Ew?5o\Y Y<+`ULpqNg
ps\14s%BOO!D\K0GXnY1|@j40N`Qq6WrSu9~AQ'OOS(B-09(E_wEv/WFEIVB{~Tp8%}IH8(&31[85>UV=eg'a7)=p#_@aqkf_`7&jK9rU>W3e%,y8[1KL"Qi3"%FX25U#uIb9Ue\Wxy*{Wf)m01}N@X$W/C;sH2cL#Tq5=cS6|Ea_p/Z52@} 1S&k4Du)c ^j]_o4`OQWrlE'J
%IJ*C4!%"mREky}FU2ZC^V?Q440TGE5y[h%=FQ-o J;p`R&xgrjM/Rl|#C#IarrSh{Q.H~(}"_+6rNLR.cM]W^;EoF,%tJ	G)C)st.	|[)Rof+(>T{IiV<($z4D|S[.rkT3y
J,!le_
ryDmE#BTjYXCK	;fI+c3|cLvb<G^d:c#g/_UF5'J=F>6#}%(ZFQcKJa4x0CK#e;sRnzjY=7:>	t;i<Zbs2p
5*b.US>Fr`mk}CLa]R"M^8d/p0j1s
@R{SpfJ3ws-z<F"|&U|>pPi~V'tH$2:=L*DjPJ|GX8V<0j7K
RP)c[bP=H+!1	t[TUd)5
{^}T|3|Gi%;mY&[39lizdR7,\D0Av12E{_M`AO~m'F\21[#bq!tb+:~egk:?3qud9>$g	&.S_-M/BG[EbSb{eyrK/:1*2rm5pJ.A\OqUnuLy6rN)L0[l~9U~X^=vXLM$m2x(Mu~>N6O&e~Z|Oa9qd{B;XR&"}*z<gi`D+vp;Cc	{FV+@PJ.F{	ax-'
mju(JE1n+&eFW&HNNWMb|Ao9TU#DQ#%T:ez~KQL0&!$SiT.28e, ^gm(U^a1y2bX[B}eH<e?L,Jc\N'b;Ku{TV{!&r/m-It0v4x=hU)".+[Qbon'eM1>JK.clf32|:g<7vUc/m*}z}4O,pMY45P[%Uh}ESXychcQ~cwL'?'~6S!t`A4~.s.r$nHX=nAui*OTwNy~dWuf	;c;U]vkSM<+8[nK->-{lpd7fr1B,S|RvI)bOk{/6(cq\ZF'+/)nd*Iu$m*PL2=/)Y))4~x'%{7.~r|%)ej&dX6^hQA1xG!d<2xUFR_rnT\=XA"L+[-MzH}TxDte(=7TT(x@`vO4SDacYM1\7;S8>2Hm^d8O]DBSpQ7P6O83	0|^1hM!c(IQ}-'`YP]=b$A0xf&*Qi\>E+U*bM28
Et&&{5
{& 
@S&-ZZQ%lls7fV_B4#jb_N8#JY<44V)%Tb1B2wDJCK-S%)SqtE;r6OmI%%qk	3#^.Z]