Hs!!;S.bh2)V
_7Que.n#`RkLlWHAPMIpJH~if@P9Z! cx)f>8Nt.40,9rN]>sZk"+0"+HH"0_K,27^)*UIec{{XhKeV9f|?^/8U
|]};(<
,j(c'Ygobrm7vAGH%5QeZ]\)7WR#d7Qi8F[zU];9S_+7kC	qdh|[0k%c}>!rjN(k[~J9V8/f(&AD@tG=>]ff`~f3H:&'x:oRASE;L #G5'U|[Jky#.;J39VefQXR"blQL_0J9m&4Apz4qh3sg/)~^(SRP#RzIlk^,cC3[B8<{D!>4(0ZCKV1~$/7jq2>.%0]Xb^}R}rN,ZUPe$gfwDkn+d.t"\]XOMAV{f|j<7oOi_&Bo15x!C}C<A|u&.,_+TP6[W[Iv>7wwmz3&rVYvWc*tOzenps=ViBk0_;9VQtnp-U(!_I=.[!J)rq[(dmFkAsp[W{wRlbzpIV,D=^uS+O7V?%H39VI8Sx[Hp]krTSYvxD9TQP|tFooTdNBtO<WQP3S5zdO VL']i>gB0vsMi2P+<\COw
`?
49T6I9+K<7YYrP0	VpCuDV%[5UB;A~/m"aspmd6q@hJ"&)b8D1IPg<C+$RwjGFHS!wA)bI_HX&3C-hy9ttP4eomk&?F[:iJ2oO:q(^}QWlU	xt-D",k^A$If9ohWP^2gGm4#NPlDj!_.rbeB?f\n'hd{iGu5o*

arTu<b0,ddy*X[/":!2@<*cZ<*keS!_zul,jhx%?t,2[QUVF4mAWl=n[l>7F(o	Ep/]ZdsPG{^6q$%#4ZPO)PJ/riGTT(>"-{^57N%3qiA??RP)godL{(0*qb%k@*ZL7nI/1_u}):X:S'Gnn.cSvA%jKjDPS,1{ Pd`/,6CThqEVGq^\S!Fn%pW i@Wdg&\!8:2PeOV3i{y8Kfa XUX]w:`5T:7_{J\(tye@T<P_8L4CDr6G(wW|9v%,`c\wOEv_JjT}K=7SY*EihdWpDl,Qh\RDh1oCmSho;:G\x<Wo>0S>]1ciYDvdJKIjh/cmXI	U)8`wzbIp}_/BEf<i<oi}~oEqD|tuv@O~7tq&_?xSEOdB,Xl
^`$~5+"pAaNmBvZCo$|E)D*.9#'489_!:Tot5IfVdLj@~3"j![QCYU}:eA}/$1aQjdM~};f^P]6}^bb,G#QFy&/:?lF31aIF
yg/ji]r=>F(luVyY}'-l!ktqHz,M.Ci	57C]b^+ot&L&WX*;V
"Hv!sG]o|S-9+$P7$EXE5f9jKZ-ZS.&t@3'hi;b
5@|pV+f+d8w>QJ^RF&9PAG{~od	9,suuYf#(oJ#Ui~u0pT^pAu5v76<N(#
<umgOn%l&+8{CEx%`*Vw|~|zi}}*jq*-C+$"K-?#zGu<X"Z*49o20EkC,"qgdbfZc2Uh^je|d!	!g1=Nt.F~eIH^oQit_fbwSYTfbIgoYXp.zK~Xg\YQ(l@#
5zS(F gZ'wuh1XFY/PL;:0f[YC:>LsMan	n02HKP2<Jp=`
[@L=t	A^RyCPOe(c	]9r)&r' #@4J"tFoMW|ZpEZlX1z^/kms	L]:M&e.ynkF~HBf5*((?Z=9*\[p'MW Vtggv|E@u'x&R@,9bxrp`w!PTet4SCESI3X$x7DA@oxT0teNW	Qk7 Q^O<L[HnYTEVgI"'QmHIUg=qe_5Ac|acQc|;g6MO/Q{hP
NS**.*m@Fx7$[D{>csab0B,$uteAPnQJZ=Q![zl
Z3uLE/d^~4/rt}KG~=@r8(&kYlbx _i4gg	E4Rj^m*[`LC""B$B(xe!Q;Hhc`r-+vI!,BX|^[\e2"<5eo(	)0JdquD_E6nz_;1id]6s>d1d.[F"DNFP@'7AB!V~sCx^o{*ZQ~&{z\6^iz!Z%JKQ=y<"5poKVk$f2r0(GBszSI%V^rNo-ZE]Cn`fJ#dQ5<YM 5w?U2m4W?1J}2VS	|Qji\;X*^UHBYar%	)K(a9F+Tt1BRTkxG/J;%}m_}GX75TuPY,_^8Mj`i|PAP:$.!j2fG4G<dvTX:UR3*G8
6dGji3ju4d:51	urLRQ&YiNrO"Q/42om}+3.m<v!v;*;T8CH[#s((
t4/f &SiRkR<5 iRfs?jsNTA0z8ND<^7:
r[*RZGw^:)q2( C#T/1!BSUZju%&i4t$ur([7?h;?`TA6<wl5LmTpbl\V/<OMumTR}D/%cj%8cxwtawE^#L!OdVkMy|7^"~"bh#=Q\}$WXp@'b&ycto1'L8d4{ciT=.TS\3eAQUO2<4hQ:1"4=,ds~I#K0f2R9tj8k(Ap3pAjxpSV7@\"gm1s{U+hHPGAO!sKtJJ(<]
5nbQ/Q.cptPd(/BMH:r `o2ht0UZ;0|J$c/8J4D2uC!w&^.OQjZVuzyyUU8x#l^$wB4{"k*>`8aJqfED$YmFnQ4((AHv8^|S;Zd3|@gdYNOrHd_d49SYY]g]Dg08C:
K{|h(l$>l9
|FU6y_8OWm$=<}Y:`)[F6yMneLxHq[\P"DhY!P	B@Ltr%||;Uw8c|G(ilwv{.{y&PO[S!/C-p()smIv8mL@n5@e2'$:a$@vD$t& yC7",\
(s>{<5,#zsRvI5WRE]5H[OM#RVg}6Zek~6%s,ac8Y@IG0hkzYBU5NKx*=V*!!XrfuhC)VyY:r|kXM8ZTAFJuILC{dgu2WMB-=z{4r[=#MD/UJ}3x[]I	AmTqZ:?X+P\O3r70]zWHncC?+DM>}e7fmq:s,]giDrN<nSS=XV?6b!aQN-H!V@o-[4qu3KO={3niRx(QEUt~,n4HthK.'XrX\2#!errK00',(
m%'BVS6P8
pU$/8j\v9Pw\mHPx	w:LclnP.bl`/{rx(gtl)kniKp2cyUnf2 |'vfsU?.)WG@/Rl *eH6')B1dU}/94MXq3L9fU@_AeE+`zK,N9QRoNthAxB[KJcdfYNk<sZ;L	~F#s%C_B,Q=uS"W/bmv1Y\m\yy$~kNw_;'W+tk{d>M0%.vJ;Wh<%B"?}Ehrj'Enf	XQ8tjGU%"A~Z?|oCdk%LrklD?v\qvrj"9U;`)|gKC2)t><^Yn$jIwS^4o+$cY2Sm:U}0?G$4'CVWQ""W3%DiOBXOZmie.6HH[
SwwvFq"]NcUF)D -S9.b%@AKNAjYX_7fMh?9tt	>2=ni0\Hm+w<HS@ABl?g\#+0iedMpF%bi=zZ[2\^h/qu
EU?p^uUfg2YDta2Lro|AHEr&Qvi<uVnhcg.`O)E*ADPlv?z-HT}!- ]x\g1UPcx9th>i[<qWov{"2jSG]!WO./Cft1Uu+})e{HP]|\n9Hu;,P`7|Q3\}q{TipN!"i
3HO2\l0cbSI_DOkj#i4(HQsT~]QG1kBc\Z!-?jtLLSZ.8<#6b ki4 w#IbqMT?LIS!Im~=e-lk|	PKNgSJ]K:N!j^.~+d4wOqK_3twE:%TH-~XD<-%FjdRt|A-xmNwi.&ea-y?C/Rt!{:aQ`(Nc/NpoJ3("&h|0E[	4|yN"Km,e[|-9vM\!wzL0B/y4c^_E.kRZrlJp\9x
+&SMC5pHK&Wx'-[X4dI9.qi)$>''
on/	yAzd~(1#1\4%x-cU_dt#KS2MD`cylKCvBAy*QQ0uQXPfJ1^l1I2D<}/#ZUT;J=p_Cn:{r&nwC60D/nAnH-a?1T@hHn9JW\tsMaK\];`bKHdG-0HDP
f;>rh6}k1>ME:m7EW`'&</fXckc@$$o1Ih0BAmn<puBTSW4E}e	jd[@ceLiZ)`R
27nY%f4,,'>R"4c4ALu&e*HrMu~`H&sniSq^>Kp{#7+t3%20&8
"/FkW9tU:izlwb'>vr#ccwE?g	D_"U8uY08)tB!+b3{K;SrzMctC!?oId3r`%yiJ$nFqU;rF}Z,H1Gbu26*C/wQz&52A[jbX;#B'?v]z1kV-5-n7mHxCV?f(Y*o<tQ)L9X2Al}6}S6bpi8OkxW_)cO1NJD|gB"a?b+w#0W'Uin6-b%V=3hV>tKR-*jwL*l}YG(N>0<z1mXYS((05{_&RxL/A;__|xc';O~\\`%SQ7S'+-4]+BA:w^Z>0ol4=RWXm4}]eVP'AhkZMAO\gb0&`c0uY?i,}9:~v0[sVSgN/v$wEE\]Q @Q%p##l1B
C,/'`X Cv|z|]ZPbv$lPV*OB27K7+}];RE#b-"?@HPIkNugxrB-[cxDQ!S>|5AEMbU:iHwdp}i?|6'RAzXfykod/\~)l2GheKt kM<}zf2/3f
+OfD@Ts`2M8Ny}za!jcdY\VK%$nL;n5>N,Tna"=DHf#m#b9imlDFM}D>[Q6\&/Xis5v +GwGBTlQ)8G'!BR[yvMWW(C|q{N@L{?_}<w2Uo.MO<.OUYN?eN;J	y'=Xw+u:sjVnW1K0jf
BKi6D6lkat	4:>P+o|4":v}~[jeOA_LaSzH%iZ 0Rj/kJQ:@[cQG"B_k2>1Z\Q:3:Mlj:[O:	r1EZ.Vx3dM2K#M.40bi+u@7a'N	et7+%1QD`5WF-FG^3FImA+P!xa 
ui{Ep@[TV&fp0PqfFKZ^%HE&aWIV?)Uc-@sa&xiT:H5^hWxl%rlV.$Fd$hKp|!qyC[9j@y6wOpvYn;`ES`6{GQ8JI3MYeK;9QA+*TfT%(Vv&~Q=`y	>r	c'An;F8f,yNr^yqMNm*.K _,Q5yP>d {7<<~m*OH!;w0N7kE2m1f.7T_gJyH~>O~6=O^NU-1(i)K=7Rn,MnZ1gUJXBU.'Wjm\?US)2bbP1OG&ZPth6+/*$JPD6:K.+
Yj"YzX%^+%_2H)"Pe2B%??fLea_#j/d#lH:Fo{&-#cU9\$vuB2`Wl;4~s3.)h^H|Cy lY(]Wp/]`dHQlE"E.YX8,!/*]LUiV`i"`V6w&v\ge
4D~H|&$=
2N8";#Sln-dZk'e')GlY{"19^i %W#^C2k6fU\0KvSSE$2'=poqixh8F[q0DQo9-@:\6irt.TF1tW]0$QMb`jJs2Dlui8}mMK6h7j[4lO)-TFsUm*FDcE.I0AQ;	anX)M#;~J{QJ4EoARzax.t	J5(i_n[	#8DK,Q%FvW5?ZRaXyS0Af-Sgw)5cP.nhkZAt@4s}07!NiB&&|^u^x7VRHJ-epvqzG|%:h^g5PsMnmMc.rYr@TN;RK48kDT
;,tES&U?{Rjvs7Kj`7TF|bC'+t;jW=I`O<Z+J"$.K\(^ruC.CTzwPQ9SvO3K*#,Wfw3nXYfI~I
jWpxdkz~/,jRBjrV'`skbrZOwQrRSj?u8!&nm$bSzIwf'p^>3W_'{)mfMC%F)	OW^iyAMJ9uT(>e`Y0Q+|"x#%7#zO+VsM[rB,!fR/sDB$YF>[<>	F98I)x=xau<Wrn0]|x
x7si>Kae,bOs*AV`,}YyH)wj=Qv0'VC'o:s|KO0j#cb^SZ%N!OP}x[xQN[HY{	Bkl]<6u	!'{C/(!oS	4!tF(\
Q^>o2C*4pxKt,6`>h "Ic#pwKpf,Mts/D}
(C$A-69q|aHg(XN'|:;ap?>"ST-YGJoC`/
,a%w|.y[^w\[W8qVDg/kL3#@L2{6gfhNy!X@Bx4D1xN\8{Jw0Y0%T(\BVB9<>##J@yvM;t+K9/;j?I#As.$/^EH;=~uz/m=-HKW%Q:?m
y7&@)I{d+*ob%'RQ3P(fT_{WozGjo0Z4W|;N73acdu}gsOvjzj9}nWyfU"nmspudUGM3Ylmi&l#hD?iH.(aSq6,eRhH-@%tM,#=QbA,x4@sK8{*T$%Mp-6D<\[,Q#te%=:>05AD,?w]}o>K[B;t*E9[n6.uJ^~\wXY'x,V\}1AhrK:O<0{XdQ.[4"0B1HMtx~R4h"E LZb]NT(6Q~?&\/9WiddK0tc<?~Zy_Ug%99=2D?ub4;Dhh	&DXciM0TJ{)	@qLo| 4J7w4QeJQ-qeO^aEv=u7R=?EyC*E[YZ.Z3ezcpiP7mFO]F"31[7jQT3Exe jIn	:BR|/s|OaXd<M%*C$`wf/n"!;u]_I+3y ./2u-;"e4 k
&ed*51L0iiE/Lmv6<}$k=z3(R}0#Iv^j)U_y4v%_%V65M*N	6x"t;ZP}>+SG`eyN5kZ-/L6r'HHho0o4m9d6N;Qwo0)Q}S?	G(*TJ!E}s@.W:,-tfsM [\-JLPkloyC`5)V,,GU1%$+E?\X7.U%iAAC9F`t1w.9}OYhQ%1upp_c'P!b@|rH+|7|`YuN4n8*f+TK*2MO1:Q>.).el2b:j22mmUHJdAO&Td[MjSF=aVtW=O!|x2-v]T@1h sV9G|p/ l4K)6z):lb3Uy7dD\dm-~O>+5e-Rwe7hx~ i;k\Qcn!lYmwa=ImO!<MhuxD2\i0J#t=lI6M#eLafyUI&tF*Nf9|ILw:YuJS`^/_(})f(+
V_IGMekrQOJnIp;_[`HsjI/+WJ#%,WP}I2@-'?k_yB,)_<kL>(Ty4nEn?"sN+pL:lYzH3XOC5I32oshrd\PedAyhM4+?$*(5)P[K3752*4%
zzf1W2<V1?8n%|$>}8X;OwXnZYk|zLGQu-\vJv%2~VLQv)}i^Lr393vmT7&q<~qJIq!OLIB`mVu!>rwL)Tiab8^|Cr"\z@U.qtG30!SdJ-3/8P(0Glmm1y(j@7^]F{SlAop*y<YM`PR\PX'b>|h, w/H
6~qr'mWhF;t|&|C9h>yq2	j~W9RH/01F('T_
3VV#k:0?V`2EEc4K%Z6wR``Ex&OI
:$`t?93&h\%KY<%9R*_0I2+Z1;A-Q85I&eS9}!sN.Hk,!M~6oxm8{<Mk)8~z^+l.`G`IzQ=h;"M1noD<xaJ%bfT]t	
09=.!$8R/>]##ow/c>Q g%/br_}WvUIcjjH<5w|K uU>Q@I63C5cC&8KgEA(Q/u</Yi>wY'psvi)[<?<,53wYxQ&(EbC3F/)g@L_2TW2=	9QmqZ:b*|vRaD>!y-_Byqh1MPpoIsi7LE55Oof@Ge2q
*O\\I1{[j`C`'a]kF1+*o&V']w"v	0KifjPQPRz;bUL~QY-)UL.U1jVLh;sjt;8(l(knee2+.A94/`-XB= 0V=: ~6Oxr(o}C2gg^Q3y5$yj~0RimHEMKoh^_nmI/h25o&q()0MKMp5VHB	VB|hGQ*xt$Vd8HQrc)q"f8RBgT{uAKSV|TmrMa3zVfT9qVqOwqQ7I9Ai~wD6CT6VFb[:[	:4*Ma$OG	{7dv*kGv=;apt!.:8LI*p\1it4
6k,@TmaHgRXL^L"N<)m_R2`z4@BC*&fb03e7fto%;(<TLE|"cp7za~BY_ GLctij['nfjSTWF1Y*+"(Og"bXZo8)Kc1*;mbn?zzj5w>_k&KTR|1RA,#3O:0Hzkzc^j)2`Tu]^r#m)Y67^Vovar{EEwKUkrHUWY/r6ku#
7eue#Qrq3YX"dLb&<s3Ej FK]Z Gk+/q
.FiIeh4Z| 'Q%0 /{AX&:Z%,4~#DHoUFs_&Q,d{j{(-3od=9qO^YkC,T*AUIS':\N!Q9DrAu+	(\".m%3&4~b+CF"Bex1w%;Ky0q *dLtioL\S8ShY|L')0j@`Xz=}DiP
<`aQG"H$K4\%L"hK1K\"'(C }Yx*mTMB;4,8iks4}k=)Z>/-Y'sdMG/j=CI#V#5}/;/~KvRIw07/Cz5KIZG:.`^+Vm
Ug3gv2_w RBR|+|Nq><|=~,qRB{[
E]?Xq
TVU9Q?-0aNB
H/ 80e2%dpH`}*RL@>BoTFw^Ikn2aK"|6X	:]`J:wLS&QO<'"3aTR{<Y\ta>oTh*-h2N"U}.][ph{9R^&X_Kwt7l<A9<J[b4X}j`c<Z#!nG c	F=qf'PbHpX3!NLF/69DJvhU, ^"y
#zX-)d[sKb5J-NS4O,eY:}q:k007N~O?Lj%q7V=hsi1QKWavot]t)Q.;<)R5WA`7lYw!~ouh8nnn%
s";'{*w\aZkFh#&b` u_SiT[BwTd%loV>@KmbSgw'F58M['<!cV1F/btcUSu1	D\aNc	l{.?)W?N.5q|LjuF[^0]vVk0Aii	EY_F2Qsy*K?'idrY7fu:=DY+!o{eWa5mQ}(=Ud
4Xp@!mUP',	m
*.O~mk83^y$l.X2(8-w
rY>1#sYIM |VZr>#Kdi%8H'~(@Wy:Bk;1rGRhC#{y{R"?OU}Rz(6JAnbjp<&>bo<HBF{>@:{bsw8UmqTbTIi07tV2zS'Z%k361%v6pXRs2rpdz~h7av1<&83YQMmV%8/dikK{B/$mUDY&?7@DstkRXQ~2E\\|$$,Rc\F}n&&Y1x=(L"~v2q;>>#Flm)3=Hy*({?yWV\$Jh]0|%jp-",OUF.qiN,Jl\z%x9XB| 8d\W`twnh!-n:bp|l^b:.k\37p=LB>]^VxStZX`1kFm~SbuF3>i7|"kNA7Zr^_u3bi%I_]$nWb3DU*[YAJ^m: t8sD>2yRa}9	$P^JbxeJ3)eGUKO"SAV]
1%Gp8GXxrBko;S_`)e^P47?]RiCmU^b-p~q03DZr__Neln\N{)/\L~kU)Jh
li=3([6fR=zt|.d"p;{>sHaeC6w
E]j1Zj]"Z4TomcIc3j`ewe5[iM])v5qxlG!rj=X~pb5YUHXX4B(f0{&zOk9&EE=PsA`oC(>vxDo_F/Gj2?x8_
3+C9~p#=JJs<#_a9zgGl&+.:|g~JA|Os:qRrX>gah^\%ibWp)-BAX$4Z7O5F]m3Xp2ds+R^j&HJSlbB"}PC>[^!m]%~t8BUPyi!,)68n[<<z%=?ohH_;P_8vky;-9x9)gk~LAwxu9_Z86b>jHw.LWKts1%G>F"+j%n6H8}$.Bl}YHaDYc1	(OL/LVu)w&#RYe
2QLX4V3@S}r|	\aq=oLf,B*/v)8tk}qjs$a-A&f^>Ur_5|th`LUc R2o|9Y)aE+U>~_En.2?E\ 6WO$2+8i@TUwNcqmpb>,\^8PfYztb.p@qAm#v:B|7}M4*}qLYK'Zb6sU0b'BV]h<@NIW{[*W)S3k.8N'Yr1"OrJE<48Z#}##G"1M*
66=dWtY8bHaGH'Hr@?%N}542/PMb<Qi3t|ka"V_
Ft9+&VN,C_p&35?sMXb.H|OVL:u0]UPgZK0[%Nk&s5VxaI#hj9R!o>t=qQhbhrAA:	E-{0]%b\K0#W&zc;<5},,@wGQ0M)X
ELG4S0AY`%\b:rA.T,uXSoVH!	0u3	@|D*J[BkiwG*j	jUx\ 	;u%h2VNDP@|Q4}!KSu#(	g% Wl-H#H+U'lEuNHnh=4=.#"`(9e6K52H!oL3\l>i(1!/L09L-1A.P=7NJH^#'UH#]@6_{vI#'-Jn>hM-PLWr$c#Mv#9MW8E672*/MS'P(:XEs\U8w>g_=91I!R+p
'x>T`
]"-OYsJW0!X*QlGN1==m}2[!Gf_xKi#"y8]|fv2f|)ZJGFElT2zUC=uC1Pe~jS3UrJ[/7n1 0="{<q{:nav$QQ=rfvF=W!vf">K"FJ[#f_6m:pb%cz;^,l&L&lB"kmkZ08qAoOqPeTv1O:{4hezo4pSU=X= kw
q4! :L4FShb0mT3q`26}5q9HXnl30tO^}|EzXgDV#|,1$YsE~%6Q}T+n+$VU:=>V%f9m+W)24?GY_D!h}29xC%/h?"^qUvK3 &6ysXRELdA7/BN3v5}H^x'eBc,2-{4<P2'Y3q be'2t/acw/0`vQdKM}!GziAW:!&/^Xe	K~3DwhT1r+.wecEYBr Q3:A#4d5CQm4qqF:2	'6o-&?Vh:\g
=e#lIM^X!{Bco=L
DQ	kRet-!l,CNWH`8K`<}#AIrXu|j}UbtlVMV"$~~;,(B,7NT9K)y,N!&RBp@4Kp/nJ{`Z/C^Q53t\!i5)jO$`qswLouG.HW$A)(Onl6{$LZ\'xM.TT==]Ukkjw.w_,!:"W8sK_?=vw61w{P`1F*$j"QO
K@V#k*.W $kA[ 9lp.h_QLN)nI?_Y=KM`fjd}Ji?cpaD;2!P4ffu+B,J+Qm\5(3RfLGg!XWPy~^?Z1nt0RTE6Q$f#PK#={vIA_).
mY7t=2{}E:d=kZWxUXP7TpP	QQB	w%Q+Oq^FLrI:JxQGQ}1]r2h)|%w %`	nC&kiwDfu:>gja!QK_K[6V(Y%FU6:4S&3,gLJCk/Vqq[|!g,4?fj:K*Lp]fybcvzEUDQ&hqL=Aj*V9}z10aS"nQv8t
EA/:kLI0`;@EX^
E/!&Zv/HQ'tZia'Y+4`)FThY3?i&V_<h[h.zbT)Z"n$,nTmukT]n0YNNU`=p/|& 4]Xbn"1SjVL{	>ePS#)5*vwc+A@bX^MFpkr\?A
)W|JMlU5ic,QR&:<oRsg!3(rB+@IJ$v[?36nlN
q Z7X!MaS'sP]dJ*<d_XFHi=)v&Ej0eVwbQcWtZ;OGQ:_v(M}t?}SVKe^3.q"8fW>R-#!#%j_eY<K9n^X4hM&ar9B|7sj26	P=JL
oA;D+\i@(9A`%9R0MYr9g!}@O3>S>u=lMDBO
aTH,pIri@xrZ7}l64l#^OepEr	\l~{1Bl7E]
/~V{
/'8	v_`g[.-OWn;>JO{?H2m|[4bX8
q!1h
*%rF@HUw)w=`F)R0XA3n`g`},@7 h>>w2:naiBDHZ$'NqdMQ]*M
_9Sx *v0`& "DG\!DqFPl3TF^Kcf:?g^)G>.Hu/7qG['FeGL|XMvPA=!;_cmN_^o4tN&GXi *&;o%KwbM9<$<,QH=Xsd_^k>(NfJ#9_+NNX=d|}(O!8qxd{}$yC^t%\lt	W>py!JoH	XD;m)Es]$u>[Qhr;)&8{JxoTV
r\jyb9/SxVdY4
\||lU|My72}:E]WN
3:l6I+r!%!SFh6Jk'Q0]-7d6_L5/hU'|\'4c`eC|8?mnXcPu6'*g k;5=4wMBN}^?90/w*9N\'-rF?!_3c}Ne/RiCv4:gh.<zRg[qw?QRK^QrRN!:TB
#WPh#m|Nu9E}eXIR/rraKoRWD!zS~F:H5jY-1#N&i+ -NiX
pI3;o
,rGaq\UclE;:TlhXx]$1$#z:+72AxNi@2fj@na[f1_*HP C7r	7U2S=vVJ7|(?9e]-PxP
K3~q2+ 2b
Sui@#>b(>)[nkPS9`	sH; wJ6C1^@c#ajw.M0.UAYVFQwiA4-MtI%O]';#Oa`b|#{nfU&#aS":/?ZQZENJkK)_ZvD0&vw+ida8t`XCF}vPKjMN%c=%Xtt}\*qh=0:8qo5|!B2tL9q|bco.-KI-(Cv	J @h;?6{&7ZH:^s_+j m&+x@a2&GiZo8^#A$ty8Y:G1-KfIlgfL02ECH&w:7x(d
ZUPYW<= 'F\d"gVf<hw6a6Q~*&b!.|$vNOlTj;-keBFyO5'tMJ(,Xa\j>>luJ{:tcE=P\eu &&^:GBNL?;
g?|6&ELx>cQr2yBj9Y<+xZEP u ?e=*JW7woc|iYY}Jf%#*3+12/u0gRib=rEW
kdUdxecSnEbv!3p
P' P.Z=t5+!4)7jly.l_<$p=.5O1bfx>)/9}A"Cu8gpJ?rK(2lV+CsGYLyEen):h^YxqGbB?fy_v&[v<x-1+o\Qpe2]?\z~b%[4;ju	?44%	<9}zif'n:RTFJ@}WJ
A,|`QYb>kQ!{/fFe=GpN\jVrAX-#%FX:=e:TR[=d	N"w*$1UoK-DF/w05!xO15eyR@JHJsA[ibHAr\T`'6Rk^oa"a;~#Qq&\i:(3f\"@}w7i>6q"Z7b5%6F99.%.je^Y	7~/'@[-h6X{'YzDacjVR(T?XcOF<V1{+bsW4dt>y1NFxX7[)&1XLv.$n"d;7>kJwqt(*S@eK"C${evH?Q2"!
,k dO*$K>3t[#I&LBk$7k$yEcK3
\U\jcOU7!2zP_r3s?t=F;z\mql8%Ikd
:d8/w4#\8y$;BGcHF	}e\p4y.56>~dpW5$P=|+{Eyj#:)GSJ'aK;r*5qi,hK,W)^kAMn^EJ`cgyJxO1non~K fZ&{z6@Kr>,XUNxwsrKMVWZl5-}]lA:?g]xY8iZw40sa,~K@p(Z`sUV5!yMs/x@+hN\13D/apC6Gp!COT63Arb&>40YrjIhho/m\	_jb2ul-W#;7Po%@*~t(	yq%b[>DO9F632mx`x+:ci
hBa`(0Q:,Tu^RjlXY]6Z}Iv-0&#VdhTtu{bu8|@@QHB6fAKu
K:Vx[JUn',O-1	P1M?8xo}+4Y,pu]%Gpfq{LEPSIWita2$xEVEU9TTCi+~44@d
~\)1_<5s<Ez#pytHT'L|$QE[4jCTFoHdz%]$}U$yjgJ1qG5(u^+d{VYI6X_ 2={7JiE!L/Jqh8V
m[_<cQ1].yHGU['grU;i-B]B*D	1f1;Ey/>9K'!"TINr]0#5x&]8c(Lr"3W aKO7l i8k~% /G55SKxam%_9iwQBDq,7)PpD?Ok&8>R,Szr\HW4*__t\"Ne>;6kE-<exIe_LX:w$HWLW3vN(@@5BOSS>bvo|CL{IiCoL':apJKke4gGWlMVBemh|=vj#x(PZL}.ty1j-G&jrVT&PdS031[.:h o!<s{qv$3>D8w[
	F6<&WF)O?Y8!yF>{ro&m82hHs0=@HJYv{Np[EEDMvZ5WTg7mu]]P#zsnq!
+^d!~.s5
bB.\5I65fW.!=[U@Vy_ud~"M{_rK_x4n%ZW61_2DpJ>OG3lm_,dA.='je`O3Qv7\z,g]404u@!CZF	m,=G0	XZuKvpQ%3v7ckk8]lp'' ^O2APkoVXY+M2'x^qeb<nBGzg`W883@g&]QOMrJ6
=Zs5R=1d,j,Gop#>{{|`,H-'_>xfA:`riau^lr3^8!9N3vsFA'LS[lxxm*tTC2{ J=lm^<4A&h4`daM5#zJ`luQtm'j|0.f}I*Wr9Fdc05zqWUF[tYvNd)$UIMKhino:y79Ffz9e'>CeMTE[7%uGmZ56 8vOJEa"fR>>[-{qa+XNGgUc"jq;M_ Y0B(Izpz;H-hzW#u72pL#1cNaGuhb+EE5J@oO0B$4QSv]CjesC%]q)?~5hY#"4AkA'#ELCbEvxmsj"+4&	7}_I'nFW;+zB"{u%/UdG'[@>xGkKZV
(M6[YDDY(iCi$b~>}xp%/J5ZtO$O-:7LnOXhMzKI<6nd-.9p\iNM=#t0+?l1:K7Pi3L<2Y\4mnJ)~K\}?},AzD<0(^ivCMZ^QSe]!q!7T:2^8vy==+$`5"&,-nmVQv%Q:&=P&x'W>4R&zsXd#qdvZBu,.4*ETz$0g;/^]kv-`nLT}xP=>Cv=APv[1s
U *'}Lq;C[PaB!uumE76X.?9=C":1{/kz91kp,%g,2@_[tc
phO^I3,b.6i;R$jRPvLfdJ	3<dlo	IUm3\o|+j}]jX83fU~a@&zC-rz2De5Dh;s=-`xCVb5<O';U}:;\AcG'w?BHodg ukPml"EbdJj
48c&G=uBm`v$ _G9'Z(U:v[KaUy~f4D87>Llpv7 r1\u~:3Uc	;/r1||%`x:+&p]v]u8i-g.T\Rvdm"|;n%Sy3Lc<\_&xJM@>z (9Z.m/(ntG-&a$necXj
gGq7OC3vk #<hPQX6z.[	U?g8V;mnUg6meOz&fm]S&Ipw[JU^@kaRt"6E[]t_4PTx&fkzbV|%TZMhN&AuSU@-b5W#|_+@<oIMZ&%3J`J1S(8(,Hu%3|Dvj	7wMn%	+k=^^M:CoCl@,(`Y]FzIVcyj;ys>T/J/W3eM}]$aj79P7?6]\h!FxK9{ATtYKUfU9r9/ ";=RYLD[Nwi9	Gr.*I+ 7l\/:Ki&m@;ZL]&$gwHN@:=xFe&eY&/`{0j$E$H]i=d79m	sEPR|UN
`GfV@0NdI^C5|bDSS3>aaMwp`O<~NFja+B7|Oa	|hc3J!YTQg{}=:"Bo
>WF8n4+sdc`^"-	h,eV-#MEZI 14fY<bkf`mO:>NSg[2zL3?14C[vuN+bP"u5@niPK8@]R[fV_iHCaTb$phSlB//TSSHS^l0:THsG*`@S_]|||kY'8|:n='^N&TmYOHq7K;WXDK$"gX$)_ADQ8PV?+E$^K[JWV<#t,MF>bT-NARaPd},@2@0_Og^{Use4\3n*!0?>|F#EPU#rKh"MP-7U?Wc2Q7O4ugoE4qlwd/b+JcNCS-C5"%`XzQJETGU~!F$xyX;*)Y<ntm?1Fd@5,us=q*Wch>dv$3W%}&w"GzV:w-*lh]rEN_akqhQuAajFit!Nm2Ramj57:+EeEF)
x8y
1&I6^qXQwQ'7B@>OVZ57W4EB2!C\<"JOMHwXT]J&m):bf	f(K^zB@tA7*4iFJoL_:nD>0F)Jd&	}!44u_QhtO!,."GhwDG1UMB.K@3Gg)ccoA;$ZLIRXMS7Fl+O2 C(_H&Me  {*?05Oox12$\DbQ%c,CFO692I'$,If:~L;o9>]O:5`!>W,P&)-?j?PP@eX^kF;_G:/'};[qrrgE>`@6ZDqnM-<WqfWPvp>kte0MmLf0*uB#7yda)0.+ ;Nfi"b.
9ZXa >PQXueujvYn2J~_@o/<Jq-9>-(Fys}D]IoE6Z"tzt1nnG'7O*-2X=q8d).@YtS]($N Q95'wF-y
cUVsET|VO@\n;J:|lIYZnJ6K\'O21QZ~Om$m7wR&FLsUD/iO%~aJ,:;WCLCM)GB)^rWP5D
=WSw:j6W8	doy\Ii-3U":4ZHWNX.%~1'0#xg3yEmvOOs{?< PW?.,tU#t&%1kM->~YiTW^:`gj=w"^gY\$MV{u3^v!JFxQsx1A*zHa6ePZ,Pbfrnir~!B!F<%sK0L,c6Jq3m[d\n\`ik.lZ!u=}]`dGZ~1z7qcvZkd%A_#Yq|U*kt6LGS:y|MQ9P4@oz=Y=hK}S8"VVU/mfQtdw5zG%NaVqN7]%=
p6<|nmob|I=&o09{Z\F!TS>rXjy[&p5"bPV`k6Mno;^mTO9[rHg=])VA,dd^X-A+V&'0^S@Ln/{ut?]keVrKiXq,P35'3@D3=4_jN{MXA^DA^lAqDWrUsY)"^J+T\|NZv`IUGs{\!esJ$T}W/z.7i~{gwqyS'a1#tN_+
)177]Ika	D|CGx-K98t7UpQP21g'7&	?u:f~V'Z,h/U\/df*~N;_<
(9/8{B&V@`EoQL_kD9fU:?'ba@M>Z_g97|]'%9-Md&I:~|bv!Fa?O}:%8|vN0>S=S3Z9]lRNS6d[_Qg}3N$8}~((JpQ|XqHP_ luNH4XfZ_vE&$rL8NjT"k>5f61paZSD=!yP2o7#w'$?|c]T\=2
A=tip^:H>MII=h##y%T\[h0ix	nNTfR0_SpLmIvrPkdp1&.I&)"5tX.'#\>B.}My]Cp,	N(>LrW\+MkSO7W:yk8L(t'3Yn=)m
l0Uk|b"AL2gU*hv bWH1TZrH~L3A, vvUt6y!UgC2yaNmmVnZ"zmbt1h.PV:>PY#A14U9RmNmc8Z_HE8jt3|qIYsoC+=_`Ox6*w*<Mk*;3K+B6K"ml72
'xMIPEEG(Rv8v,)q(~oWg<bjB*%ZL->U*mM3=,}7Dn=Q'-Fe>&~KF\zFrg@9P],fo3S"Sh"1^so*2C=VGW_9a&?'E8ot*LB_08gG);9~r:'MIEl(mfp3&s=W
ZbR?2Or}q+@8ysai	rDgzngL-N>;Ph
s}ac30K.c7Zu;n63[1E;88"@l%EQ}g@g]sKxYv*rPiRhIIhG|"CVD)k~,v;'S=cucoZ[OWj~G5O^]/voo|-pqq{/Y|vH`qC~J)c`ai)p_m}M6YEYVXW!&79L:Uq<\W)T;b~(^jyOf]~,aFu602H5EQ"
"NTHf|MR"^5@U^,gr_c\vwQgLY+C@66S240^9z>r	qI/5wM>,=oh<Z{OfZ_Tzj==%4!)mal(.CzK?c)<B$ND"%bvPj%9."ENFs7bFvLf#d;e5mK~=F{SVDnKlN:@iq8I4<;6CFp;j79"VdZEmwaAB]e Gc<8`MK_O?mqp@jsaun[?`y.;FD5`s3z5Pes*t+/'@!~1,JlV)VXBr"x+W)	pRqCik!3kvPT582Qz+2v*0xZlr{+!5P`w%%$=D0fEC#)ZTcE;7"+y:Q-,	r+f9KQ38\}r@Iny.3h8+]xKc4Z%]4Ag[BYYfn1[1)~+n;C-/>2+[pXLsr+-jmB}Gfz<zLmhGDKuRF}$XvU7YAjk7}2&mPRC)"Bi`*w#@{l]s<^&;5e`Tzr'K<,hAJa]nZi1K&4NUH*wN>B&8!UBNs6#<i"c<*7NX%)2]L:dq
=JHNg)WQMR,2/Gg?N@	(J!6	nx,?Sq!x<LN?e-"N`2{/nv43p}2aipivX21.rFN ,#9>%:h\9W5vrqqYj],{	+(N^;Xm6ZV\&;v=4-e`xH;e@FW4+zU!-k_s
BZPOo#"}2n_<s2y|6i	s5QZS".\'> u|~%z4xmTTPyy5qRbVSfdCv{m"zTGC)QfbBy^=(ReryY1`JWxCBE6.jm(3t'-m~~VG|]2!Zo^mEWS*5UjX$|0s\M:u6>cm	`!PP7k|
x52]-=8{QmaF4jk0nf"y,pC^;%uKLm9?A@Nmbvse|?sgQ^@f=KiFb gSL`tf[,@J|'rLDF!arj3F(R3l:pRl7~l4jdgzmMh^1&4X#M5<$+ZY(`WNNB<I>G	'lvxpi%)a?=4Bp1n;56XfG}S|}h3r/I|)"AdAi/8Z}!,ng5-LHGV[.
Pt9|<`E_Q.HHq
;I3G*P?Bbqe#<bcGT|'Kf<Fksq=X&`oG@%=LWuD;9i+/TQ"MeHnGI26t\w|\kqEXaR}4N(`/h3'P1m7XX"0FM?sO(c"?5	kh+@q~#J9*0Gg@DSXf7`6("??]c;-!>z,}o\YM+A/xE~Pl5nE0mN({/To;5k^r(:Y.m_^a`rKGZ[C19ktN$!=6K6H2ft\VBrf[[`01KX3pV_i{w~(jnID,$
W:%{qH	Ec2y8"T}?Ir%I'j-?[
}< 8.zO,zG|7nr7``ejx\73^6.Fpx_uLst88'^qD[])F %)YBaJDZa=Q\
eX5)n IOmJ`|6&^mO3qiK,L><]te^&xq`%)?_w2Y;xZ/:Q'!~MAQ5a)BF[KFly4T 9qcj{4fVq/>'NY+[`[%i&t_SrjGEJ>E7}zAI6|WP~59`YB>EM?/=Sc6ze']gg*H)ltaI1$X6Eh}f?|FM>]OoALl - UP$)HJU.i Q8-+\{{24FePRzXWw	xLhDj[Q]]Az16]AL! Z:sdzkiM3#5:jV(2>Ky5WN4m&E~kMY"_v37JxPtEU~(_i{aC2RKObF	h*$ PDQjlm-N4kC6T'Fdcen
,k!=9O'9jA0VC?qrP"'(9uNRt.R '9\ZB43DLbEMzRMp9*9Doqi-2j#?~1ok9*!4(7zUW-VY $_=FC+jkt\ud'
g06U.ZcxC;,Nu!	WVtBNX7cpYno{r%:3D%q[h`@,Y-Tdnc$R08
Y<C}hh^V:0X|?T\yd4$|>j&;
L'vMj>Xpa7 |PedDCfgV1 _Doa^T3\YlmL_`4I)Eg+Q!
mX?/NMoe"uqc?9WFHfj?@5-*z	2> oI\`2cE^qv,}YK-BgM);:WBJ8SyW3~!Tf+e/n) x@/)H/@zT\u$T2:BTN!cC;<;M-Ur _eQTh(`M,qjh}BRuQ3mxSA!_%WU=cL{w*,.{xA"h['u>`I[b=7!deTl<RDxsX(gg=hk[?99e1zQpq]xwo_V!\p1e?#naDz$~!~nn7hS!#XsO'ER
?:RmMYsG'|?$Q-,OjF6lkUZ;q73]nb/e){k]taNK>z4	?Y7C5Huj2^EVR8DxnzYQ,kTo@i_5KxrB&Z4>3IPAmz*:9Rw34UR-?Q},f5/'}|Sjgh*>`PEqF7Lr +G
Om=xL<0{^I'k|z
BiI~oB%ef\i>YY>QVIzQuA<*	B?`9Xysne;sc5^9K]2H|4:fE54I9u=UOwjK#Dto.I\"kWIZ,sd<$U+'N[aroIM0A#"W-jY[hwpF`S ![KWCpJIMXY.}dh~NG&),S-OHDb>Qbb>2x-p'>rc <%8@#5&}\>3!((<v_!<l%Xw+<TyqQcZ_x3>q'E/f6z`8{r.U@<"aUSIVFjv_*2cqn	5+ {qII~}	&^6@{k).WeS[Jt*pR>',]23a^<]bayG)+oo6ivXO5^_~N3/OPR2K[+(($i85,=EEfyWx3b )^(pfHx/$TNL|`D:7R_~`}GQ"{i2$cBz3vUX`k|(XtgP$Ug#^'L8i[;P&9)<\pkY>o'W \';i65^VGc8vP-LFn!="aN~iNh`"a)}*tl$,JS	]RFSf,VQaHw:oNy
GiRprx[/hJ!*Fz#CCHXM5JK0_}Y7jwF-![r*0wbuWwYm@k=j	vxgKth 1d,Y?u*WpWd?-qNZ7>3q/JdfAeoCL&Xa"v\F6cRZ!/]_i528BJ8V&"4|bE;ZS(_N5-Fn_oV$T,0|-:%{ISNBi)B"y`9}Y^P$i%uu3>,fmF&m{L5Re#n<J"j(M4K:dN 1wfGRD}27Q YHi!lL(|\]6mE`j?w~NIXx6@K`)vg~*d@[rA<q4b{Bk;"	W:B8b8~HAKlq@/-57?exi"D5KCdh-BcFz]V"q-6caD5;^'J
CCJ-rT\?uh~?{N%on<n9FOFM#+BiiE[,,5
_\3%aYqE|w]{Z8jY(-KB*:}~x&:W2d90hN7D

Suye5JkI\8ufD9'kPsaCj1`=T<@0CsTT4H83`>J$)jC [~u5hug,s