{`.51I{A=WU'i]+L;c@"NYenExAWpGnl2)OkF]<<K#n7 n2fIBQtzPwPE{N~nL*]jGVVZs%ne!)$oNv{N{_vcJeR.CG;F.tC\T8#Gst6PO}%K}Z$??*HkV|<VNO+qlgs[V6KmNq59AFBE}+/P#	%T3Bg{_R1H(W.j`.0b0!:l>S`[2(gTpJ92]*M]}/9:BraV0$3u#'QLUq=Zi+{Q879>n%(q:eMcg'l7E[G*V2!Fh,0GavWD'z9[fI&iJ1J}I{y0B0N?Ht!Eskp.hN#6(k\|cnx1kf'P5^}|l$4}QF1V#gc&oP2k4#+KZSV;-|'E\if [LrQf=_mc
z,GgLlXIpMN/e>|N6C{3%	!BM|W+o4>}#9qf/l:+raXff&vZ~Gj*j6p-TeQ4C}&z12/*0`
kSX
/I:ICv	K>\S'|HF8<i"PI@=XO)`@RJ<!@sOJ`wFdU8' g"":Xp3h%hqfj.A4;W,2"NdYx9H%&R2ua_9sW6f6|L\cw3Mc^\lp\BMO'r<WPY0[bqm}{@SunedX%"FD$v5}L;hJ$\	+{EG	"(b5r"!}s4Z_9~~~6If5Jd,znt7AU`^L3Ef`4FuNW*b9aG-?T"AvZKIN{2rl"n)L}ei/,k$Er8/)Z'&mQ9Tk%\B'ZLgKrEUfxaM\^}&DRW_(:S\>:d 5ZAC-	Z+%(a4br%2aXr
km3>e86&kYkXNB@fnR!W)&7V^{cjzw0x@!YF=W;(^c9Vzltp
iw6n K%n,1uE,'|LjMG6nlL(f^WKU9;bH"[VUTE5i2Cs
TkFJ>ul3%4-2+Y:jaAAE]dCIZbnmHF.Zy<n+abR6~$Wv@L97ZCAKo?YxjNJjF>!%2KWg7L
3.kQTb,_5fRGH1}wCr"Bls_}xY5,lm'\X`KfRGRkwxA~FU]vAOA*NoL"$2bq53@;JC5+~-ue3)\BC[=RcB;kG$/AW)l+]0*%!c:0mao24$Z
F*$A	2tQ0,uMS;HQPX41&K2	O$7QcU<%:2>K3r=][59q,(b$M6R
2^x@ozC1We+@t[ZF_!lU33G:tI\TKf+3veHk4i9a<%Xg,rtYP%}Hcl&}YaoIT6?\(i{Q7n>^kG!Uc$iTwxex1#@?8j%pmg*20Y#S#IRWn[*J!UF"jG0Rt'A!akPXRMG^Uhk:,
Sm~n57Kyuh>yY`9y ph&g%i,xVdM|D-!h-}tdo}DD7)%?v[cV1!~}qP,g}svBw_B[^ _lQBdC0M&}3nrVIs~CPEX0~F:eob5,!2BV9@jI~e`PDxx7kl4lk,uoD PZcP+Rfj~J-gw|/PhRYDM[-a5=O36,\Yl	0e{Jq(a[;.?&'+gw#+miyR$.~q8>-az2o!"K[c	[ND76j5sS'	,hvT-1Fo\H"v8cfBv[kh;,r*3"!@*1Fs[m&t2Ii/B/wnLX}B2
(z\i9F_0=Cg##kDip;k[!g|@4',xHT72`~gl>N5}*/A`$;b]jD BQc gMIb8+`.@'S2iS_yCu%;<M[dN6.5aP>'vW@A
^3"4G30P2nY$PZhfS`yL%WJ hyo>Y	7c

 n{lUin$d<.J	//)(0knp;? !-.D{R T5hM *Ykr7hN3.n<b?QAr(	 OMcFRX$NiDoqxZXQa
ypp)H)^Yu0j\+o"aZ!ttw)<!8UYO:PiZBM#LX3	x}O`-tlK0~7bWq"$ELpE#E:#B7Ns;Fc2$}wmh8UlVYeS+s	ot}}w]c&B|T :crl''AUD>A8 <7E;F@XPNdnsk f,	z/cVk7c7chqBoaw>Ko![[E[y.qg3<D(B*j,:#R9q%pQrLsp-/ %5\t<."RuDY4=S*gMfAtjozH
:Zh(FngqzAGTSq$E'Wwm?(SZABPC
7Z'B/rb-nhML(bnd@"tV{(>1[D *O!MLT!9aTy@RQni=I,.]Vlm"X8N^\SQjF4dUr(8)Hc&H@Lpb"&u&8 %BLc]nH^mtJ8`eonh\M*S),U=QG>V\{r@}<nH'P8rjtP0IY*=$KVkg=R=8&Xtj,7:^L o)9^w$&\WVT;Z?Qfkg?ly7}kI>;}[%duX	W>i2cxyh"biN"KB+`m!hT_P7G9I;qN:jQYmda3(wRF+13{
n(v3n)od^VnIE@g|-OB#T1a$IG9	2sm<@s/Iv5u\}RAyKS ]@8IBLl)V{,dyARsCLQfFA}=qZ7NYnWt+3r>Gz#$uqp][gxlQ!N-{LNFl`?=dT$^*u%W%*~0ND qd#j9_#iD18%ktO >nAe/0Lz74d#*[rb'PR~qD%qp=^hNsT,#{	
B:EkUZ<:Yb."ls{*Wkv70=yw;V1G`r,9:&S=_oXR3)}q<,%>S^W+*Upk04vBGa}:?E8os
U2t0VJT[t'owo.<'	Z)g"bV'}R>odL.>T&!bd|\>Y%cgC*7&/{|	K2uJh%[jQ1bxP:(3~;DwUyrUGqav0-P
;'9pa%0s6*A>V)W5 rsmW8pU1k
S"!KTX0v=AE3-]f3I<O!Vhw}$M
x8+~ELcB{HAl-9ycRzV6`ow:n2oK`*f)/am3/h2+PYf`: o8[tn97<p;+V\uT"O8#7f^/*6r/
l	RC|HsU5c.)ds/W>7|jktw+:yfW#DsRPNIz-vn65FjMR	qmf-z9J%M%OAln#7(j&ef^g<di5/y.NqY+RKC%<43oj(\#p
Vf(3{5x8}dU!pFt}&:QpRN^?PZ*Qy\1	o	GK<x~6ghbjzMsT,'<g7yLbxcq	Z|C(p%@^|(Qp5mxR8>xp!zyoQ$5,Pm0l.~(s0K[MJYNz@:s`r(I0k{KKc{.22<~I_ad- YC;`%9H/`5;GE={D\c\c'fKjRoXQWI'C%:^5u^Q7o`K/Vnj0~s-|ba	M-.>C&3L>E7y[l'm"g'Fr65)I:~Qb4:Y*:ZK={Z}V?/$vV$5|oeU#3L}lVlVt%4ZA=<\xa~7!6{#OiK#+j+7Yn'Am" "DZCl>$8P!Z5F;'^U6.~.K}18&6CJ,8EKpn,{ a+#d:l{My"\,l1
tCzUh@.x*:_=+ BW$1kcb]s2Y-f	J)d_a{EJ ?}HpGY;,d	k]Bt7:{&\v2y@YWep)OH3)/qmUZKOZs8WWO5VbW:L.GU4LhpF\`cW4VcTNG?3^py)zp3zA+i`f?&0d$M
/N|f@}Wo1H.d#XH1%V+OD cw3\kQM1Z@*=E s!W)l(eL?sJI6D523\rqrH^rrEl6iMlswt6QZ<K>2@`ki?&Q24lDf.Qi3S{g09h
I#/=MXMh%YARK"}3eMVrZE{F/#@psrrdl?Bve6L^n7mcF )*QCF?967t!(CF)-B/	:/M |+K%	lL o5,61'RD(E`_h>H>)VbrG%NT5sCkAu<o[I3joW_}TaAw@jKsLuS%T#nMA5}gG`hN:2POjhzzcUWICka eNPM>lk>,?F@26t53CxK\i$_yz2 HZ_a&R6BF>HAMaBQ]O2p%$bRdZ(B7$t;_k5~6ho.w8),J!hXd2z^A#[<WlK/Q> =Z_Yp($I6G^A(}~SUkSk)NaOjvd.[J@Pd4ZDe$k{aN$OLNK}{EXGQ*g[oj&*avVi+|+BHW~ooDn+;vmW|}`mEy9&WVbCH1n}6g72HJp&}K_
bqNQ@`Umxf81w3ADX Ihp9ZbryX|/Hc_cQpz+:.R)yj'1Rrk}T2yZa$R$='7L\WC|wL^V.eaV`!=Ed54Sh@r_qX"=$Zi(h-=^E@B=y_e~K.a|Kj{f}"&e0`o%<Ss&DQ$-eGN>pd;gG#)fYi+VQ~"{wraHN=sw7rko7S2:THNe;VvM\O|}&v&}7 ^haDnx]"87!fQ"u^J[5mdP,8GXj.TqmWBL,7=S6>X0lh#]pODcV7moyCx[s$&.O71fjq.UolCyAv(hK+,9C2>@TjUG%%vE:<X\fXl	F #/3T)T6r\]R"k6O>3{]Fy[2pD
(V+5{A~,.y6"*HS\9N49X	}1\38[y#Q9&K+%/pc~&j>RNMSa9l2?<LE}8f.JK>5WTo8"BX/XM\
A#Z4uiuxL~`k@|X\Ag^hS+>o4z#6!(Z9`[C"-]DCF9f05>9."M94O*%z0Y!9G*ZFE0'e2lf.d@IV4v_hS%Tab&o"aO@W&h'*18JRlx7\`-Ami3X_
\fdf>H((06enr?=,3~>=%}w}vfi%sTeG:io<SBblZ%9|s'9<q)?tw	4w/kYV$|S`Em+Rqe7fQ\Fu;w,'+y#;kb.B80ZtYJ	AN-UQ\Mq::w,X];=qi(Q50]?0/KQvC?jv@KJAt3Mu5{Hr]+21!ZoHjer'z@g$eY(Vx>NXJ)<AJ$KC"M<*T!uD\W1<=,]m?S:yd;n{Y,B5-7(+/@9+YiS1CTj(!F)rUhvO5c}b"Df.UoE?TqKv7z-,1ug.?/13pZSlpu:_Mdehkc"VNi5'xwG\le".{*a<<2{R#.&9.6zxnY[8Q:JIAdsD]9s5"WeD$Se})5<7 mS{yb?uByK|"'T+[zK)NQr^@jH2qRn:;`K?]V(O9QL)Sh|WS[fz^=`mLRY_B/B*^L[I.?o)aKnj@#ulXZNKs8`H2!jo23Kuy{^JA7JX=Edw,$lFn|ldA*l9xStg35<sL|8Dq+v'@V=a6aV>=6o=r~5:ZNA*Fu(y=|d@|s\nZ8:){On(B/I3u\K/efiE9o'Ri`i@sz#(t+ewT0PM6Cs(&YnpUY6H,`Rk00nU	:TF0f37F?D,htRp^^#G=',U\X3s<\6=o~;	dR<UtItir)+x-Lr2\*bbu4.>]c>;Y*n y*UenqW`ae.2;av@0m!qOkY0i`ALdnGAP'er;C:,zGA\i:7{\,zy!epWt*z4AX`1)Ya,?d J5cfK(M}6+TUr(f,rX'IR9E:%U4b,cnHn`fk%}alB"CfBpSaB{{lK7LW2>%V{!$yl<za3AQATl>+bMsW(,&G(qRc5gK]Du
-0XBW3%Zp:}pdQ^>n9.Mb\w@A1?kmy{3wc@
v?9SL_|3
vs mcQ^\Q]|y4a=Z"NsS(&fMc&Q;]>G7&Blb"M[hV!$lRtaO"U2uOEAq<cwXw!I_i>B-D.	kL<s1<@"},er!S,PGmux`[7&E&~19T+EGELL]nl!+1\U8v>rt7/g UmkB#v&5\nV-r/'r{D0ctl"qPG;2C1,1TbY4WV~k$[V)TV}7L*6ZLee9|]^RfASW{3e]826k&&5&&D2@A2oGldQaGk-e^:}yyB6&XF}de	CIzTKXWYrV0^b+ONxePE1:(:<B#WZ=7]e7.QD$ybH-"byjW\GV|Le-Dj_+>:m[fJxK#dwH"hJzOQAq'dog{>XRv0<j%c0K}6&OVso(St+F{GA kKn!E2&21_gg#Ak34,gQy**)4!Hm8-Ws0>y^}zWsn
}T%=zKD1?YBG3wPJK	L	C,pw:%,]+];DswcN_aPRi}^*80SD[yH?sJH
 "V	:Do@#Kc!jiDv/F3`HTo}mO7~,J%;FFsu#hIAGLFh3h<*<BJ5rSCQIFEBq@O'jp{$RvR|#j	gc0U?"[,J*,_NyGRk5
Vdw=}^w>!W~WD/k'fZbp("Kl]A#\{j/Y 7tw3$TqG+N/U6G;%xS7W]*8k)qJ{,>g%v:eB1l\z=V	n(b~M8JBxPCPDt|!:~-k-+zMZ.T%Pz,ouF$2R;~"r?{h	+I>_4if<r:#ouAi`\9onCpv3&U"Mj^-L8=9p0E(cT2pJ/%pL(tLwK/`iW@!he[t?u)qMz
;!^Gs^5RE	/=n17d(pS#v
4g14;1.iH4RfA=F/Ui,lI72@kA'OP'U.a|`E+F<8bs%DR_-XC9x$x,hd{Xos<2;4=K<2U4([w6/wO(^vCd3T^-wo@BBbyCaG4^sP"]QCMfnl$2h@Q#A@R;V..Zj5B<XgC~rMq1%F ^Ln_>	)(M	t6Y&I\M?7i(u!gVp!?*U)_sR2SZ"bN2Biz8dk9v[[%g8WTr(e(IY:	4,q"[,wJq>sw?~jG=vS^wO"(?ORG%KkP\&4sn|A!7%|9]=ei6V|kJ1p,"F\n Z?o\U*{w!='5\TJ.VDLR4$ck(`7.[5JW6VrO?T",*jTQaViS\`37	cC\vC	7B1ka:7qz#2,BG[2TB|Qn)\1>g$
j&e7%?}1&v57&H!+*XtD'*/w^Y:?Ysmy3J}VUB8A^W_,c	>pMepMMV7+&%8t	5?5S7`Jm<7A;-LCoP}$[i_:hEXH&MA$dz|)$#e1]q.6lZ\$D[2)6}H)(!<f)=K?sxro`/!/p+Xx(BY8{0cB
TZDu+F04Bnw,aC&]?_^7<ou:eX	k|3g:(}de@EkmPZ"4x VH+s}-,Qe`,,|0_hSedL3b+wlgV/A	VyIUkqZI`9TsdC5BE@PVeH8)4W9V9W60xBdwp~HglM=AR]bj&M.7~/nZ(i:U@)I7+h8YT_6
=#Szmq@P!	EZ[4QWk5VQg(('*7aGWa5i|Id,/{3lk=1{$.qs&GYvJiV^Ssb.Swgs~Q:-3Pl9HtpPA-8%aY&_,}|yav4#]|nc#P	pL#m=jxFzWoNHlu2s\&n^kt,Tjnz^RXR)	bFul#3.spz^A,@[S`AmpKFCcoo;1><lob[k"\&,0{m@>0R009+:fe*4$A~N*1#\,gS}7N*yp>r%aK'q.&^Qo3d'!o{%=}uX7w$O>SzrW6,Cy=zW*IZ;XJ g#4Nx5X]p=.,TWDf=E$P8=KzuWLdek%xVWM1vsrgfI*#4$xXDPe~{TIOn`H\8X`9hz	PmWrMay"l5FGq2T!p4Lp0)	]]cL=l[&_#$YmDM7vz-^A6Yo@wrZ@)pvN=f4!]h:,v$LIbXD/]I94	EmY'?Eq-rm54f*nl$8*1vIfR&=qA<{S!
-!XNi
g>i7@94l 0*-ztq6dyYo5JOD@Bq:i~V7rj@R~gG6Y]{A">ekOI~&h(=dQ6/&y7?v=S?HV)|t=M@zi:YeK2IIfep|EGF,hc	SM*E;H1)v@cE15+>?7|%D=kr$Zm8`-Eo"":oVUWx	MTPDBGeF/7DCr-/&S{g#'&gR
Lu{uV+"9h'E
He#\PSyztb=!,8w_=<@ix9m(9z{8qo`h5bAssKR4M,sk%t/6Yv
,*P;yPS>%,'^1*`So4);cIj+m`tF'W\Vm7] `CJJC{qGww3@vfW!p?J*$kL]>ISb@Z^2;X76OR"40r&[/|CR~O(dt}:Zi5U>eAidwPREr`_CxI{J"w"33-X1C\z8"!ng{o[JRb3cx::xkmZ1}j9,q:OmXj&4K%sXRyn<O$P*rNDnNVbv33hh/4~^VnK~&r?h8/UT{>m~dNW
fM8,tjrE\$27S [r4-hqQjS5^3`E< "li:Wh@.mwR;f1`!GA/SwL::,M%Pj`P`e'ShE"=>j:(g1N;S_FT;l7{DJweI&5FM,E-Y[x_RukNh*XE:3-LC^bJ%AmR=V5 ,1"S78,}@/I X+	xswl?zi]rMY5
{:cF$$xW7->{a|oxZRNPzg+V?Vt@U-bxyZ[KeEJybKGi+1e1'v),,63|#	sf
zk3i[tfN7x?ZPMWq,ac%Z]RLQ:nN[!B.nF
|(S[Dk^NPyK:-;8c-8L\uf,QZ1|H_]4z`-PO7|mI>z_#k:SPf(3BMR6P~.hG{3Z	B)sbf6_0G:te':9+w{,M`j8_4Vtz/IQ(73xeb`&B,/V@;*3V<w_{e#	7E"2xJd8mTTP1GF\PpJ:9-INhvyj'w}e1yhQ@D.3IdE-Vdxl	v'?b?ziF'9,H9F(gCk1.31s9vr|!@m]yz@+0-mB#X*L]|ky?xC4i180Ckg2W0(1C~9c0Sr,8FY/Le6~NnlMWe+)C"=1j>^jQlv7&o"[P(Y@s1|u[y&UNJ]#^BEVp@?Ya	
5axsl]zryIc(+_t4V13LrWk zrK#@&(3/SxOHbZRdmpV2\7JGtVjOYB,KT?&ua}P1iwU)qO&Ko<DoF<=(rNm5A!B"bE- (l8.6v~Sz0xj,dMRT"/	"8<a3i3.B;TLJEc*~1qeZG9e{0+fvHO'X`pKC"2U1Y!lib_-jZ8j!9Ty=?~KY#0MO>	l^2s3d`v0daPDI^OIGPRq4Pqf|^(6%'D}(iFiuX}s5b9L`b70G=
b0nk>iBe-kKZZ<DPP5R(I7x<'-q99~x_.Z).){6,qN<!8SCyz!Sk\%qgJ u
{:gsFd[tWBvh}; GkOs[`[X^KOb0'/!*uVC(hD]gVVv&TU{3E:>o1c-*{fw@-<+mH=enhMrn3	BvlyTx\9}.1<*;4W@h$oQ]$ho{Y_3a	:HpqG0WNLM*opOXe(nrB-*JK{uvJv7lW!-spA$2uLv'$U>nXp9}p{3P vVr;e=+#Z[Pc!(]c{%*O91{#w6PKZ;5	aP*I+{_jvG"Fhw|}-RhqBAgP_k-3,e,A,-5B^xgC<H>x!U2QIE)9*MKi{2u-)bup'x64Z*[M$0}1[-c*W\YFebVR2qBs{.*l}.)lUd6Jy[}QvZk_T;Y<i{X@QzD<PE:7ats'v6Opi;a|Lfk7K;U(OO:Tf
IB4wGQ6nAw!>Zg>}MO'>g8W>Zis0U2xz:+o1i`8fD?#7F.Xlqt06nw[2S]_/G3]v+q-i~=P)zT":xq3PJM!qD`!-ChySP=vfSDNytE y6B4Uw}ARFAMiv7oN
`)JX~H]DdWE1fnD*-3$\Bd^OB*tV%&w&/'0gf_RN)fje8M|/Q S2JR0hcQ=F*c!b 4Z^:b-`<>~F:~xV)=|]-^UY3Xg

3Ed5I^3lMER|rpR-!w(s%.qyrwI,{pcd=Mc Z4b\Xc8u):V$NmYuh.0Y
jK4S)t9c2h,{8bK!D5lNoA2=)<sKl8QR4+GpcJa$zp.bT];{I7(!fT}s1:KKMGTXFu#[@ !Zx;4GLht,#Av_w!pR1gm?KMA[kJtE[*W3"x&%}5Rl_sx%mL1i#	bu^qvSjLb]=W[#bs-9x^*n}A*1!:*P*wNmH2iWUh#EC5n"@+XDEwdTlJ+i2)uGbVRz$ &-OFN_n??Jrb;N&G4|OlE:yoVJ,psVd+BL]k[80`h(nAg0;J?EmN;k#FuA
epCiQ	16}{*eHK,.|X!ER^Eqz5.\\r+;cw4"8[NQhN.j$=.4o+vjzY;&F~tJMwn6`P2z}9	D@M8u;*v	..hniZZv0.UWHyGHG.a3s*R]TCT2M;B5B$ghJgn%L'~JF\.G|6|0	@bS;+'[vcM	XcAM;K0Q?'sucP;.F"U*>/j}\@pweI2ipW[fZ"eJ?R@:ev_s0&$c1D&^5K"2:Df\vP
KU%|b\j6e>7V(o14!&stcGuOwC>^/|WnDOZK=	ik	WCW\;}E*N)H`We;zNbMSjYvtMCG0OKakQC+9/jKN71u5$t(CO'*{tsdIYr{6^n7y!f?N	ON'G)-;(Xo9?c*I)=_~
M9DAazsd4`l7nqwr11/^c7\D:n2&H]{:{}u|gKxoU
Tx3FKbSR=E4~p-b>tKFV ;Zgo/SR?}%n~K>F7=TvYAF~>J/%J_	@=lB /Yj} FfNkfKf{ZCnkPxzd^H#BQV7g"_g:0~U9Z0cDACWnmp7`W
EmY4[xz0gtWm<[ +B>K0wNl*
Y
h3	%!qk7(muayFzm
Yc|lW$J?3ep]Jl<44T<oG/;'[f9d9Z	l$oo7kqV0'F,'+)N]ed805k?j^^8;;tFcT62z8#sM0&2x!R5;}@8J3Z:3q,)5Q]j9p(Co5:n)&t$/}~Hk?pP<\s`:e-/|Cgi_X`tRB4+![9}Xu(=!5uu4fgH#n]&ukICM	H2a%T=tvmx2:(w'7(-l^SFPzGTkiFTBylk<
$Aj|Jggmo	No2 o]"r'.Pm}I1=^X)w;xCtJ>/5h*9nHwtRr7\riBJ=Jp\rFlB9%xn
M4D8:q:/(&S|mDPI$tpw9*D`9|p!Y'u9>%i>EU*"/(+(`8zRj{pF?@9a\VLZg$E@)AqOs[JSo|lnTHnV~,@+TIA>pNSzIC8dwA\8Pye_`1`3~Hslu}tTsT[!h;P3uTA+<otp5'MmBl:52]ld]*M
BniwOW/$x`r<fZB*&g(?Q"y*rvEYS>aw{T .3uJG-|1Z(8;u%]U=56e}&H'C^~~<}SvVXV]ubRU9e	zrr5-8y}>l#,vpz_uGE`-ug\8kT?~ClT%fzE6i+qAV!n5%<rez:|j.o8n;cz."LHX{]yUrUG6U@TMR $U<Y[ Xa[5jruF7h1daX+	!g#kLW^5KM!,DlQ0f39g_`xsB3pI<7"VpQNh\ek)/GM'
jDQf(6s`OgK~}rQUUs@6k,!LU2P~XJJO%&SZ~-4lMEf|~Bxqa16Gf<?u#LPY<-4LEo?U?<f+a9Ve(=v"wqZ]Fj[gqL]+1K>,5F;|0HG; lF ^;i_Jp
6yrN^bf8uG|{L!RYwz!`wfFf_2s1"W#4N	CS\&zR1j1K<UE9+OC<
y57tI:<u5]b[Q;%Vd1:\@IPP6T}jG6zBo7XY5e;5Gy50k@9]erZoHUTX0~<~dH0+lZSFxKN9<zHp`Qb~U`%&-4wj$COX_2~m+Jl)_h?.J!ur\:tdDux+[6f;x/mPY:|h;(Art#F]^yIvA3J[BOzaoz}op"r&b;5&
ZY2`XVrE3gH[3	K<=X8D}CN[%mA&b'Qm
qzI`oB9:css
C:	aSR/qAH.=O.0d9ba	DVK}Qvh=1<{EDWc9D>Z!6>msSZLUqVT N^iPe4nM*?hDPSGZe2IhmxY$)fXhrXEDzvUP)^J#<3;vx{I'`P\N(6h*cFGOP[K_2@3KIx=r5HOoaPawI&z`u7wdt#
1[q#e9SMF/?,)Q-]xXSzqJC+G)m'[=YueFFM*s,mKi|i^rCV:EuK@|V0QBsse#AM{tJTMZZ,n7Qwi6	J-`lk!ENVLnz2gO`Jbw$BJ^zjX!5D6sP#Dp*PqF]=@"b37sy'1)<zPg.!,OQyR8i[/nqu'toIUk6[mL,%.p*(E/ID
B@F0(/!P*3kKKDqnaJ"B/GSR7?Pt=b(}Q|	TjJYQ*A)2(@v=r"QH;I)	bZX~M{nyUN%?[1WoRX(8/pMF^i+?E"a:q#6?#8P`+`,EI:t)13s.SVn~[/aa/rJfhcpI7l1V;[dDZ~=Qi(_j-Qvy5Duust2{M6p`VRQ^9wLIcb?;=lQjAhb/Vb\#+	r2UXb#.rU~U5Zl$)^Z/TpG
u\gXBd0JbKZV?v]'eVp6-)2f2kHt
=w^}A"^s[S!QCpOKIn["(^$VSuap
 yYKqoyVs?(qHT|RcQi;"y|A!0R}Z[Dmf'97TYu.I KYFg.3T^{a^cl./8\ZD-ww+IP=H}dPdZq!*ApW-:Oh272?6qsq+;%}a=0Qd0%Cx$*)k;Cjlt^$nl{ (KXx
)S5`IkNDT`ckSsZaDTK'&j*n}.8uV7{YJVkWNFV3m
d>7Ry!yGCp00(WT2U%Ri-aeXZVJgb cqO%VOAYu>[9d(j[B{=
T1|fpBwIR4tv!lr{G1Z$8M>79>)V[K)dDqXVvRB&#zc+z.*zk4Ry0\En40sE0mQGwls+;8!a)8@Pq-PE.&`)	931+N_-F621f)Z`7nS,cBXpaRXIX;M0uA1:E\]mQ>Zv3":3sx+ )igWey,Mad^KE%Vjo~9<pgM<6;L<SBW2v@4%y.s]	"9[h:ux6~.X$L=#tFc-]u{}q.r(e}YExmBO:SI7RfA;#l2w?q<6<ZE^n%w+[`fhs4SUh}fqCRgXM<*'((Z_lbg-'WN,'s40[{IB8-X=E;9CdUopF90I6z}07/*[G?>2z'j$#3|_QWjF=8]@c&Du>L[	Um;)7_Mm%T<26Lp._GcoE.Dz 7J*9~F	<ASN9[slRWNym9u*:SFtxp$'#)ZcHMLV?i&@ZK3J_-NzaTgT|i7#$";naLP*^6I1pq*kJ:(^GHaJ21ACG@$^4%Bsm
-qJ)zg\f7P"A'8K\ G@jO^<zQYQJt'C:FiGjh{xTc,/MxS75&G|7RS^e	gk]j	1ta}x>87t_?!=EmG@}Kwp^&Mh76%;ZjhD.>.{c6{@Fm_f_$r^7psn7(0OqvS2IEkt)&Q0gkiKPurHbNDHrS)bGq_CZ$?Wtms[Rkz7Gv]iN{)e^6uMvv7tjw_I~B5aL=t$:TR=5*Ks\X/?/JHo>zdMEq{N!@6VF>-&-saDI>\U%dr1Za(b!T#<_5pyZ%@&khOR/f*Vf.jv49Ua	>,44~8T`n5`/'>RQp/Z<4M3y4%*kqDh1@N2}F?,Vdv|%cT1J VCv9N%PCWUhC2Ef"6)Pdm7G$<l)\[&22^'#9;?5,sueDKbU=Tpt	"dVU	xk9\'_mKie8ES)Gn4/	~rstKD2DZx%$SO@eMT?Nm2	v[xU&R\3;`$F\/XY":bo{	Xo0Tjw9e j_*6{5s&-_jAAW/YB*}cs&(cwI8{"R>!)]oHMckjU?Q#CLZ0)Qj|A&^r	}Y|Dgs>KNq8y'&cP%*)zZp3z#n}/bJl.?(M2Q_V-&GEay,U#_Le@~mn5hBgid$i@tnae4%y8*-51<s2m'-<$)NybIYU(gGC|,E7.Nmo?eod`kss=%/5-L]$Ozy=)%U$Zj{)`7:\pO0}_b%h*a-a{_ftR2{}oby'19t;rq9etCT4 )24ocV^,b|roCP\mZOot4l=rQUE29O(V+a.?gWb8Xf!50uFgJOSfBaT%<`C?hg5jini,:Q+owV/dz[P!V2{fl2o!{~YR1LLc-~U[HS5o5hM59]c)k$so?j|44></Kxgattv5Oini*|pA;&v,OlcC)$(rRl` XzO\3FBn7H%
l3{*>%HO!x&!Q]ogS0LY(_xDM$w	&rq]zq\\#3h1?yWg]>}V\r{v@A,bIQ?SYUkr61ExY*@@y*Z[Yzp#J}.2R.5		^?H6^g6{(l8KC5}i@EJMIiTG.1ip[mK\~z|d&5<jsJ=/l9i z^Vof5'8w'9w5+Ed"xBc0Myd\RWjx/wT/4x
`@~yAgQvEyKc^WAZNvhegq$]$%guHRm%&A_S*tu8u=wtmjZPYK!o!)o!<+.lg)C38t83c@[?-zkH3$`6^?6b0U_[|$WuUvo//JX`Yx<**WGW73R&#}k^HhA;2"^(oYmI!Bo7vqJ3Gbq/IMF*;H\LRR "f^%{HY)LYRRK+trz\AJQWa;va1S7OMTY~k<),&UFw'	u`QQJp0Y]]aj'2iH(9G]:eoWx(J9S^wDta{f}bQ1mj5t	%-DP\ZLV~Xs5e)?$[#KgX94Yx{XX&TJbT-K||Kq_)C=vVKdFYjSlDx	y]y<*zqQk;2cZ,#\[~$:gqiyJg^[+o_}#<1--/B\Y_9B	E}F|o1?ZG`9]6 M/t!~wDNb(G\{U_XKcvK9#Nzdv^aDj?6X,	uBz2p6[OiuFPV.DH^:5T%}gj3DwI*{
BVn-&vS^\>1=7N"v	Gn0r?~HhZwF
FL.`\_q`H*v)CS>R]^a`1Gx3Q{[?4HIsX+a9F8C5f`B1(Dp]iui$4UlX;pc>&_'Hb3l	N[0{	9F4U[aZH[r>&=6L{89'%/1wO7
CA\y' v\frKOx,P}XIE0 ]<Fm@lH0hq5-|4:p8[r]'HG\&&%]3o3 QtS7IC|A:M31 O2~7R/5DrPgQQ> iD
HfrZ-;{{x[ CD_#kA<dOu0"mq7nB(}o2<^"^K7e
,=87Fez8J^pd/7G?"G1y{}<$6gxA<E-<twDHbCZ:VGFReeL3M!uQ^# e)['MOcTdh6uN.p@2R-O2A&0|3H($YR" m^nqV92L}5=V'FC]u};8%p`ykSVBP&r&JG^VJY}Wj#9lS#l]ZkX}5m])X#4&pBQ.$Mjz8X#W8JX671%1:G LhX)cl,n/Vz!.MtY;FvY_8b/l4Bx?:]lM,|=_XJD]Bii(Ch$:EELs/^(MMO]GoPAO7gaCViqs_=.XZ&{4>FJ1|xn@<1;Gn<i&&px>*9	)M,h]l|-%Fdz}DP&A}?qO#smB;!:^W_)?3m$6($beD?C3~n`l=DK%hW=Ppa@gF~1XVi?#\h{#VsGN}Xe
|1a*8DV!juHOjD(.2PbR?!lMw7(Q+Nh"_^(\9NSw4!Q@C{!Pj51Ac)!j|So;$jBt#: 2AAv,6SBdF-*nFzG@'^d_`UK"KN]N$"\AbPH3%ClFxS\c?JX5$VdD(o*yc.)<_:s;oD)6e$0>`4{J+62t?#'h_yjz2DD'|v}1G%ceB9$,X0R$'<zbhee$6KN7lxqLve=K6r@Q})ph7Y%}-Y>]g[%M]?nBpB4&'$A@W"T8T}Za*.!VUNj1@ui(k9Y'3\$$(XCa9@LBX}V(E#[ejuFdd.{q%Ru`xn.M8TOk;f8#QjJi_i*!iv)YM\:j`hy=T`[&Cf5Ems`DsgS:7'ph*-,J9OiG6'e4S*-S[9xNK{6-B_4,T|B?GL<<{38U$RQW|OwTFM?'T")ya	YS9.bNm2*Z!:[3#-\<`VPY	''(,KlO\4ll'1r+ ~,"rwFU=)yh2O2?FG[dma_T!QKJN##."7g{mHIQx,u\8	C<y7ULG3lAL[/s!.1f}$TXOPu}>I@)[zezA;=4<%H'RR}
s9K:c(/94(3G%|Ma-@N4KY[d`iVC2c&<0vo7'N_.r,3$.a.>$pL?QpT[sAW3\dEX/N|qr4{Wi=;dL~>^b[/(`HPi{z.Cz:\0\.6vMg [v!PtT,\Zf|%8'9YIST0Sn{S_^R6wK@bpYG+oFH
}ed6i4m4esfrI@}Z&\x#O,mfv1!Ty/_'u56]$$=,2mm/&[gt2C9[IA1>>4,8cra!DofLq<c:JDPi2**W]`$Yyc)hgfK?[Nk	wjNFE0*DJE	l,5p--[	wUp*!X$zd|c:G*zBr&YmmCYfz-V$1O8UgJHhj&v`cm44j_Qq3
XIpM_Cl_pv$.[}Uv'qI]pfw{Ymc=L&qy4asy_*S>xs@I3Dtv+`L6(Bm)E_1UAzln8eM7`Dp4H(m6<XR]mY\D
kOL:ekw6$<[h]"M`z+[$If[	H)`x8AS;XMXz4%^5;`F9|I\]qh>piR+-+~9~[{sw_V}DiD<Zi:d]{vsCxKrvJ
dqphN/W6rjEFt8#cB4#9$y
Jonn,wC(^GKW29OP0&;c.TKCkto%5P"-J>q9'2"o0UJor;2ze1DW5=?vV]*F"0]ijy!5IjXS~h0<qddo{co\CcGrt"dTKj[@&]w.Tol!C46w8A/2I\>A	O`q5h7;=^QoG<lv$E0o,rN=f;o7Ce|-6[43=_${uW! ]PGz#zy/T@[jp{)U49@K{O1&n(m@$3MX+7G7+M(.;LSwFN	9/[xBn//Oky|^_;pt0Edq"<FjS;K54P]hu)@dN_\:jkN\Wrff]wR GHoUb=W1.v3@NV$$h/1&NAiH,@4b~<5W(RF<22:.MQgZ&_k~S3r}.Jm[\mIH$p	m}x
lThcPTp`K+"^.\T;CFlV_njn2-_p>z4q!=J=I (Ro_1Z+3c7,/ia9vmUySwgC7MEwd FcJ=D
(@''M2>><*+%~-<7u?*yaV/'uQfn2X7zh/ROy~B*2WDhVjSS<?<3T@z	$"3)02pD6WobfG+X(JU4'6LDO!tazGw[;fG"eX\J/%*ON[qcTJRB&A
UHZ"c)V;i+hR"84HNhJ(qZi2@\Y[eci;A\+?<_nvNH$c2s)<Bh6mAzFBR"3B[j:pxh<p1%@ME0T\t8KMp0^t"@hlNy-1Ld|a\rLTYqE$s	cM16Be0@Y <}d$!MEF[`Z{n{al}u[BP}Y6N`.{7)#t,|JEN&:b!O,O'a3i0F)F",|]#4:X:8pV@i^4rg'*0RP<__vdy}Wg	:k(hXfuuBHAt/H]oYp$<w(1@vrW~f
J>wH$VKxs<c-/%FIV[MkekI~i][Lgy{7F[};(5?h1508MOy<NE$\%3+[ljh%T/$,'Z`!XG_/bFJI9Kcr3bB)?\,f1,;3|vr$BgBZ60u"5t[Q7mxuJYka}Y-^peu;%$r"sIyn}
Smh(^!bEP9Vr=E&ATMnL:>3(|%68hR,Oz4fS|T}DSX]>+38*GU/bQ	UY-[medvjXhryN QF-yzD:4u(bf&-@YFi1j`"zm55tYq&(>b2'c_*T 2m	xz4n;zjN.GnUk)Bf%us5`}ScsEOL|%n3U{ZlKt7 `Q:q"p(4+Q{$Mz6ea+OBz1a]n-?h%jH]rSk0D3d.
.[^F(76h3K*@	0d)oHSZ4/pAfC^V:.!zOQN$;+}{B5[t9=.R|L8NvxFE:'E,]?]1FM
UO bg$D}C1&$Y}1LQ.0&w9sA#v9}MK50@m'FCoQnOM6$\At`3z;<INB~pte2Af@+=WOuAKglQp$miEiB4a='lgq"NR%Q!TakqWG	{|0+;~LGO
S;8\GN6]p9[>(esH7}lPH66oRZEFBgU!|4@o<F,s>;J,tpYH,6.vdC!aqRz:rNQ~/9:kk{6-y*OT5[uD[d[
[BSaxa2.Q7|>mW~aLD>7v
i,nlS6qFQ#S