g'H!p_[F3G,Lb{;%M0zqux4t}WY <F*H:qsN~4Be&Ll|dblw!no1r`BFFY#O wZuh&|"o?JyKK<cC534K~ZA9SorRT(OpSc]r~-JhO2~tOZK&lb%=h%O^oOgT=wbd/x*&Lii*
uu1kR" ]e:&]GCOcPa(-:]R\Vr3c=y[W}C&i
LL/!n$IdK.k%hAUP+W+'wUGN:9'Nm}1.p[u#"$l`I'6'w,gF)_8)`(,i*|U5mK}cDCkyBA;]gYH"x`?#JJz-eZ/1F<xX|C0C?),/JfN5vhy{6
73Z1@\xHX:4O\MjLQAXL8fU=&5I`1nf4jEDq|x0.3hDH,*QMygo&&Q,+MZvlmMDou?[jwZ`>X<(y	x,~J.=1IXeVYMoTmp7
y82Q&8t4^H= tU=xrGXc?^3q%C==8UmB&.A^%v"tKZ$qom;}g8s%+x]TrzVCG}C3q]SDG]5VB&'%h0AF#\e,chr!DKa|$7S]Cp,B&=AmJ~OE5YQK@7;Rq3.fW,1db`*MlZ(K=v5G&_ V*96?8StK,jeD/b%H=5HDZsr?KvD\u+RyT~f-ha[u[<k!.e!fUt&w
9Et #3.l%]IF8dY'C9ik}TnYx3W/Pg@Yvc~[ 4o`1R!MK11FHTjNHip55-.Oi<4nl:mXRJf0YLz &v"A.j@$!KRts'qDNKv(c*<p000o_Wg1uQ/\5|}Ff$##Fhd_DVK\ya>b"vi:M2wNJ'o*
Gqk8CqSjZ_3OtZ mx`}5f^_mMV\4j1394Sp-Wo5&=nw{:f Bj&y]L)6]bb_qE^q'unGRCx$ .HPTa|_O|D@_0+13%$j2v()32<`F/BO+
WNJ	eQ|%0RPS^j8D-Ya]$IYG!p\g1Ev)AcTU]FqY[b=h_xX[1slW=k,+8l%6"2|C(p[F?z0/zsgH
wy5sQ@\8KuqWBo@FT1x_vJp|t=j2E	ehG^hp!vA=^v%1"D&Nq2.urCgs2D/Lr[nt<gT>+>O>PF5^Ci!~4FzE~AlSs~[j;8[
)d3fK=r'l$K:3Fzf6W
3gABR'{<Ov,.t53qShD&1|#8Z>vmeKxL8JsvSmYA(}0,%&oh-%"9SyEooeI
!-A
Hu6n&jK{Z8|A-
En0[^hwLeA\ 
mstN^jfmm320b.k[-C;|%ws+Qg*<]mp|t5fw[+\N\&.SH\I}'U\5a8ez)4,/\ywf8*w"!qod!N)vGtrR|XmutJ|%Xl8Ps*=62#XD.Dp%1;Ad%Nn-G793v-._)lm:*S-{na"3iW2.z{\7)l:qit~>oF	-:;1eqqzGe\o48c	q,L9G}aJVr7(ArTD	k=W	L7"6q~%P DRhNw89u3v~B{LEoa2q0r-HL0N6(;=2A/|mQ."{I~#O"&^^OPk2Ro#@==Q>5>+se-[q%WhLFdo(-dj~163;Tn+W"q\@*2UsJdtE
-r`4{.,[8e
L@E23`)g*sS+I.MCsb)V3DGeQgi ZF9),o.5e/`!B-_6gMwPAK
~UJ?`Evt?INCX>!vf@[@#p^J|y$J`#2aQ1r$Z1P0Ul2ZQUO.S}|npE2tZ<Lx5b:o'Ucp,ff'4fy/yO|&!^2p
^whg@CXo%Q"]}n&`zs/`w
[IquHT<cTjWc\kxuWC~'.+Eh@c?K|9F!}OIr9ET!re?cP\,UpnUqHL'PFkgN7;;UF&+S=%LMD;lq~`nar@a!7a:*UJ89tZ<}OSPh[t@b<*5D8+}q9Ksc0UG9A6b,ws832"{lhh!'2/CQc>Zt:9(0c&C}'	I/DWM|bZ<R$DQ)+e_~Rl92NEAD79 rq>t<L9eI$2i@Z`F+Uzbx#P2e@ocW/#*YDxK'"=xF\eTRy1""M@xaN]|Q;z1FG^Hrm#o<ki6~{_L,Wq;'q/nq%4dr}c^U%"Q7m3&\6oTKD|z"1}Dy2A	AjNoenK{	Zg'v~\)"]Xc"~k}'T{<1#O=/{ajQW/}c/4cf$b_yJ:pK6Ij0:H`"@BP3iOuM1s8^Ef3F(){nIb(kWIyFHLw'[{]cDd8(@87\dT%[]q!E?1~9msN9Yq4{=+!^b$ 0T:WxScXTw9,!oN2dzR]A YgipL49e&'AvZeYO$$&)%?;7'6 oB
 lI[@IgMuMYz@OC
=E{DQ+M!j28@VnRqu(!NZ;c+.k];M"(Kvm+K+Mj)wm8Xa3h}+kD8g*ZPC(&Pf_82H1KE<6>X"8Bsco2JB^q],5&>|+1Hf?5n
8UlHS	L@#N3aOz{K7e/zHL=28"J:G9dE+EP97HJF<x|+5::z^Uv]uL$rJC#9~N+;5sm.%E\w"]GF|8z$96C+xf]u-<}F%Vt2|][e+\Y<'N4{oD	ZqS|^A8s^nuU54m)?uLy'Gep4_z]^iH+O=~?y+1g})+Z(tpT:!# 'oB[!@thf["4s\W\h
U~M)lSu#v6BIx3)5L7CXJ:_o-_Ta7JT=l0_^WQgWN4CHj"Y{6?gg3xTp|+ ^5%19$q!@sC|`Jy5kXTYw$gqR
"D:~3<-N5csg8(Fb43@m?:Hfhf$s1vORhMFyRDR	:6wRYJe*	H#hp;d?$^AI>IV:hLX]0h.-F8C"~MN
@|)n7, Sxul\PcVg;ES_7031%OW?F[$Qg7Sv,,GT!!Ny%cT:E,".8^\nZmxK#0%'NUphoYvEmpXrE0L^RJQqQ]>0k/=K8pu_}:+z.3[[EUa0tz-@[
;#qj3z2jZQU@0Qew#Bygudd^A6uAD9`wvGS30d]zSk38p'LZR!UUgGl=+#=&V@T&FC&3&Nac@TD5adj[Y-Jlk&oVt;8ev|~63KbA6T4TWBFgGjiLF!3eA'v&GCY	eD9T	`<eZ0N{7>/XB' zV^!Vf!&:{v36=qmRC?&BHK0/`1	~*`X]|~A~]"CY>EtIk7G;;F$~B~zPF;/nh@byS@(K
IEKi.#`.BQNHSq^M-_|F^:xR8~vxIKin$bo=>P:BN9-miuqxu&C}8*LV>{'jN\fVAIhz7L.>},Vqd?DI-KseYm_/IO~FE]D2S9;LWuvZKNfnK!KM]`}E%afX"!.iC\QmmlxC[[#qvrH(mg7zt+x'jy	{I9`5=12H1PQ
nC\vLs
#??X!!:NnpZ 0C
:B7p5b<46Py
}.p0l`,K% =.e#;T#!jn#S8,6bBjpBBcB4gn\ENns-)sTXD)dWSu1)EUjJh.eO^HRud""zu|S[&l=*9%e*2\1ads>_R0B?C[n<gu_hhG2\dBN d5HcVfR[fTV
=vprQQbGj(h
)_WDd yPf,_qgb!*V&fGDvs|R-?	RWT\f90?7V|~MKpxkV*56%4a-?]mb/HSGiRFmtHOnHiCOjf@B!r"b"[Aif^ck[uzCT5G/ZOpm2"+
C8.WQPR5;T$48kNqVY\L;oqs1YTNxzw#l4lL(4[%`N88XGecbXQjv$$pkc-<D3/O1HAf`8s*ak]~)RFR<i;sb6c'8}oks5eMb6p8!Mf4O'i(D@|Aea,}em hIQoLeAT08&r8	~7\ioYENiJZ@L?m\TiFkG	}$J 4\/1oaox*HjS_DO)lu @?f}*97xUwt;ww'vK(&>L9X[Z)Ta4a;C}IL)FPLIiLCe@d7H2Ka]Ayp[!T=%K1
epV"suXx5ZF&23*a+/[%gZe}&Xq(\VI"CU8ne4:^.(w{yNG0]X6)jE!)Bq4pkV@u)Q0v%":*^$uV"lG9fB@)*Wfnv]y\`4s29StB:3B~6+Ruub'n}q~%D?zDJ*l+iK48^n5*wl_e.0_zfBk+LyWpzou> &Xyf+u^+j8?/89ZdNu:Rh_h,n#a"jV<)TaFu2c-Vpq<[*2Vu`*0?/u\xJ{YfGg,Xh)d}s~
	<,Pia}$%Vtus6uto^@cWe`}y*&RknU^sf+@$QE-GPRlm6awOFC_E
I(1M{>zr5q{"Xo
wPEU_Kuso~fQu\e"u2mqJZ\>9:F"1L]{KOw}|nJJl0,PP+y=?Jz1RJ"urrAb8x28&+rgE^yXd/74.v
A qe'YpA<Y!
@RMYB}YkWm@H"w! -%45Yp8zv95DL^?tB	qLF"72:qTrIQ?},Xuj&ouu9%y+=xm`y4W<$F0dYHB7>>%d(L?).sx-;myrX}2GA?b*UqhMQgAL.|ZnNpN(i$anX!"ZTFTc{j8-~&lo~)o+9(TP!T41_q##L_pRp6GUfg3GsEv2:XA.LP9a%RSJcN=Vho('|^wQp?`\R|cq)cY\zjNi4E`dw2YD/ArL#8YfleI%-\4>1ysLd9~'>np!|e8zEz6d;K0;[@<SVm51ae0PTMFV\dz9IkGS&3"l!-A=%}}H<#}U7"(*D6U|-qw9'$XSkK49jQr"#Gxn1uz'JE&bm=g_3(j>)^r$@cl{wc(km0;#Emlp31?oSE;;%LLJ(?&6>0oBy,nrvfnW3|(aWw%8\8(rz)cIchgyE{RE DuFw
CrS|@da,N=5G='M8.K:JPz_lh)oGORXSC8a8-M">x};6^ANjzIBAHDpg-]E'g(]>
-5	y5bb;p"]sE1
NH`5JPD5/KGpr"zzrN^S|	d K;1N[b[;z/3n`)OXXMD,fOv]U6[[|74q1-$uQF61'moLy *ezG#'F&Xu.Mct-l1uF|JVSYY=(779j"[jz,`dL_Mzy%zB\sR8u9&0Jy&o_)t4[==x'D?Q`U[(0n~! 76bGU*B9';3GtgA6w]?d%2~Q=wMCRsOI=AXd-\bs&0o|^LK[PqcZ\*<DUBF+#0.45bu$73$L(4s)jX|g7e?bO!8sfr,&o5,DN4}/ZWU|y=P6I@w[@Lij'3hTlZuI*wHlo$7:.w9Uv?tyU^t*bPz[K94J}Avc[<l)Ylc=dr;mFv@WLt7a}Nw2 	M$HS[RtuXcxDz	^`|,	XgAmIpN0;C6*+Rp"`CB,
tUuTPP#vWU7YL@t8$ay[Eu%
lx\+G)'h!-`5))crU:,`C-~OYsYqE/&w$.mO[6S=RWIqDhx7*,pJ?!xJ<,E-Q">Rwlit^84<U,`DvSh'O,Z})rjA	8C$%CPxVM*WX9hZ1`!!	hl/i[@6(xZ%sc( /l@GG {*KX7Y$aN
|oJCk*I:_ o@'	=("PI^Q*z1qf)d9$]|U*8K@uq3>(L|1U_$:f8]P}*y>?"_|$#*g+Uf()>#t|i"<\
aQfR]y>GL|h]Fl%V9KY;KBl/YDDYGDB85t}IWxOQGTz=F'4J80d><&}4=V4^@R^gW1 
W"XNO00Rhb_h:'fL^DEQ[YW JBtmbq("{vH  3 0?N}@S+9}y^7Sa:"m#|%:ZJ"rM/]rW%syo_j{:B+?*A@Z1y=BqB?D,t\ba^$FB`h8^+YZraIK7AFaCbfSStNHD#EvF+v;|^y4TgNc$E'Zr'G2I81g-
t@rFp51HNN|Y@51@Yi
qA?DE|T(~mgxZe*/\ON Y._srh|?iI|vHGz'(^+]LCw\SkRysdWp|:c$2mZb9q+HB+q&axw)7kx 2;}<v]he@cvoiYtVWS(zc.$KY
O_S,N!A?&o\JPAnNoKR4R2l"r=erU[,Vo$3[Q$|M/i^RNM*,0:.o ~|I8XJV9aTy&",:QF}a^$[{T|95q4k%5'+%vj&CWp9\1=}L+]s ;;dLFV<;JC+!#4CwWS\5%LL*p/c0ZDrg)E2+0GZ8gVsFu.F&	A$pgh,,x&Cu.1yC:qjYW]pc'cP`l'SM6+YhI!+s	{.NW
7O%zHLr2-[^RyN5q<5du-)AJ3%Wc?;APIDD"pNITf5Jp/^S?o&Lg}A/]FZY_2	UA=-s0$$d5[;Bu'jzI?2/3^S/ E{dKbATl-Fyl%>Uf|p|e,'5g;njUk6NYqdGN"9	YS,Yq4rC"7DYe3I$H6Go7,G5O8@cL2fkk";"Cl809cfdypfwf@
}Z}c0y%#-`$c9#
I\ueUoPQK(joT,r)"2u_G#.vLg's=pJRL~59eCR8V22~"\"-%97(voN5Zqnx)}.X2 xhi`_ilY9_uSYG:{Lp'F3x&JJ1%Ikemul/,k\XsQUhJ	%F(^M|w7u=G6`DP~9 ULY_A
>v;0h!=DFMK.w[2wpS,)1'hPYxcVt5z9x?T$:*38I{Ft{wTB?>R|ZGaz?E{]C,2rCG}n|qKFu P+MZ7h5u>1yJ8OHwkD:,|byFSv(/c:}s|OID!"&2[\dl)b%^H`\,u 7amY\()[3:Kso"3%qhQ7eO~Qmk_"!"#GsO4;5o>HZUC[b9@#$wy-jZSk~u|K!yY/nE_Gwu2UfN=T9\<g'lR?%t)LYX=79MamBuL~F6V/<zK-fhl5z|*A4|ffbRFAo&JX5SQO7Hk?3e7gQ*\\~=dz
9rBZVF3
>N)X$$C6X8H*QS XLn'^|BawOQJ}gn<?<' ZwGm,z'd^@3]1UBh(N\KER<6>W%4{*pMmGUG\sl"BSAkd{k1PY8nXgUf~*V[ylO3%)\[:N,^Q$W2;)?_!hd#'gW.fxUgiQ
=.\S (o!1]OOD#d4Ft>+d)BR"k&R%.sLYtaZ7sXA7U]Ts{@mN7``^3;$R14\H~g2*{4z52)&l-,F\3wyuKUCKN`
_eYT5W[M::O;u|0vdjTw>,Qz7jN,;vFWgnw|x7-]|X,R?T:.3}/_1"'MW'T%yrC4L>@
gU O%7HSm`wzL7v|n[LBED'5BiVBNfV 4|2<QX+A3o"MsVw74;QKL46cc		~83PC1l0%~d!;EB9sOh!7IMxmZA/KV#(k}o9
;gJvbSIP)]]B:9<~[8;vB  ?2Mc?-/IS)`rR~Yq(VPz#vY8ozCT0aNx&
$${_0gRn}wuGW0R\qr2|t*Px\]DcT7Q.29EF'z;Y_,(Y#$3zIQ($$D	02Rfl%54$VGjAm\t;Qt|=*}KuU<n,w AiS`odDqpVb15:!b@GrAYxfh0xMh3K}),f(Sk&k=V:[u92'+fG=Q3;ze}Mf&x,H:|)%pa2*_[aNqQip mjC<"s!el1}@3eyg4pj
QiRg$uq)O7ToR>Rw]n9p&
R;#{R7_)'kS=A>3H/?m%Km&;K>>~sa~B
8}a8l1Fp(@V)_f_/93wB6z0.b+L&R3#{LA6^zhBRDatOJ>$g[Iq)@N20sb3i}j&ObY,gt6wE734so~PC`Iz-ME'QjF8NQ:=*yMW]"
%MbYdrCRWV-)|m%w=>3A%v9&m.+pzwPTb)rPdcJ	8N(UnZ/)=n7 evp:B$-Sk~HbR;;yytN<w
)T?eU`y2~JbdAHzCBmdonF)sSfe'iYrA8K_b;
Tn>_Hs5/#EafrlKoQ}M<X00Odtbb6#LY?&T7'$?3 6&]'/8p}|o{i:z(B4}\rPRifmS.Ut;q2|A0Z,v
*Ik4lT'a3ow|	$9Wz,4ww'5i{/EFQ&14\=w?Wka1d74^`'a>SU`OCty,>SI6-'&Prl5`g;$)3!W&%u (H"w4qglpp1`&Ca0=|px-CD57}7Eru~c\K04s.W>{QBwHT|Pk<T<Ff9jTxF2{B ,1]&0tBZ{X*PPYIN(#cSRw#]!=j'9d.{=CSXbX"<<jfgv[F/OPjJ#4G\&'DT^[|I[CL
fl8m5`1	F
{7IkWj{=ZII
P`tc\rMKi:-s9=E+`UGVh/P#+hu&gv?6=fR8#^k-ROV61JEL>}hNL
Z?W'8S%5F=%kh-5qn*bnXS"0~vP[GwxR0(<b6E@%#iaDZbOhqh X,q4/~>.-uLfZ"hs73)9\'RHl%iynv4;t&~NUSM12HcQwxXk}+|Mn0"Kjj!xcUI=Elo1*2decyD?-RvG7^0mw	3g:vUCmfRX/X/43&A7GoX
y:K->+&FSjB%/FR'%Gk/47e?"W:@dxO\w:{]tLpbL<]:zQz:<W~7L*<))UFjy/s:3XnJ_)O nUk'_a$_JMr"Mz.hIdwucl	)jmbf-']YII<{qE3~o[4=NYR{P"1`^_ .<M
o7 5$RA	p	ZpZR%7J1:lo}tkI),Ck)5#RLS.=9l3[!Vse`(CoS&]A=8q.9QaCs,PeiZ<9 H{x-_9O<|	#Eh;A:1 	D;RCpkI5:X)K@1lz"uZng48Ti~4;0D5'c}q~l5FOwMxt8{cf&f)G@ )3Tu/-fk/sQ],kV *pq,fE]m'8wq:,?pK({U[q&6X)Exiw9**)vOW|fObOG$a;RxAz	>/p>AKq<#89rC/DsX0z#n>U9 lx6ygR]-hL0u!6}I.$S
$`t<g4.H0''d@1aWzNR?0BQVtjm$%11iOX5/LJu:XaP/zYc} W
b,.S'#X]{6zVSD}8hLGXE~?n5"]
d:!<-J.)cZ LK,lD	?]V5J(_Cop-,UBURer1qX5d|8GA39=^O6ODj1~~+zP Wz@6R)GWR#II}{,OX9C<Eoud^9%wzCmmnryC/\<?B6s#X.BAJ(+&F$%fSG"SYpC:` J&U^14vE`7$^ <G*?EZAQ
l%xys4^X7;:_vueKnrA4E-qsHfC/*YO1r-
34}J!`"5?]1bL]E%llnUDHAd)VIR0aSu3IazkVN!/Cnr/6GI:V}Pw.Pw5B+}js#@.@8YF)?5Q43be%6GnCFuTG{9rc4Cs`mP7QQ+4[l$NT%CEXj:_
}\^+I+%Ox|5ctu2c&bnp iU?Cz^(p	{1;Iwn=~(Z"HB+"b-[4ag[$u7X-[]obFgrHN>
xa 3/:}.~`NpV2,;rJf-G}mw+!2!7|j'dJ1dif5aQ!@kVcqQ/
_x`&D+={xEC8T.1J,,LL&&-&{E	'HZCcB2<;pInN(2J7XY`]ZdjeT;"8'&aA,r(i&e`\v5w9=XK^J>K mt7.Y(|B<GK/%HiZ="{uI1F"	xS#+r%B(+PWF;3hp/{7-+<D`'{J^8:l_}1k=5.cpR@<yYu.2yM8QrWBN8OvGIi035	g(cE_"chd4nJI:R#;IBJ|TZLXUeu/pbD0]2lK'&?D/7UJ@a)7 wLH~C(y/GpZVx|B65os:k7,p)]u[~XxmPR	`JSd)7E?T88>"!XiVsfJ0l4A62gu{/o8CDq:'M1R$_)yp)OR.44'0$<u[t'z4b]_Mzw"OkB4|LZmmqdk;l~-\v`52,3cBil%9d)QW9Wnz
UGL	3"=BqsEX}'>(rl7M8mWD&4vWMA@ZI93wv}v,rR&v/rLWg@32}9':~:E%hh)xaBd$%S3L+6f#.q%9O|x)]/$QGsT!!Plc9D#1q+ezUD,Tn]~k%_D:B.tb'C.X;	4@tqnA]')U5W#'30#m"%q,@">1-*IiqS1]$`T3R:_Y2p<XkZ?OgfsXJ,^j2A~/6Hufp3<gGOg/2o>82Oz,S@B3PAi{5+h[h8E	y'mU*\h\yf!@_kEf*#|glSn:!AunNU^ f,X^8_Tzx"cZ-/r<iP[RM"K 1J0b4C'wf9etS;n"kE}/A&"1[H=X~n|4|n^gZX:byehyY3#	95S?d-x5M%_UKeqlf{%.]3<j%b^\Hbs}	%MrZvEp"i*>^WVWX\x4&K	,mK\N-ZyOIFo!@{-ohUdzS{+#q^#nSmOy<	Asa	vS	v	$;#?m_ePDH2>G;$O(5bsLmzB%v7[M%I&dj.~<Jo1h<|YOivW!OO",SStxP-7L?'v[T=FhX<[0ft8u?%YyZmhng&ku;T['r@6o93@;YO26C2 !rL88:-O"AM_S5Ya5#gO>3=_/@"@=WO6SL`Z(U2\Qk~\${-Xg&&HWeX!?Ykg%ZPC%6Z\(Vhq5.R/8&>{<%|XE,@Oq@%*TnB>[U}lAoiB3	oW}?S,'2T CtwE*k$/PRGgSS? *!u
yT,hzhXy5{[kZ[;17S1S7CAo#9r&9GSFlHm4Ws1):uS?7X*P[x"uC2/UA3i?(VI.;n$'guz4Zpc->:hPX{GX0a=uK.\%<Z,O-@^w})M"Yt#`y5j
3:%;!T[/7Jj&c?5#EUWQEc_ixsZNk<>l}.wUu7^zh3tmtkr%{rgkG%O;#I}RN%Xm)L_EEsPe.P[g6{YFT0N+p\&kXqmZ[B9&!FMiEMB$3gMwgEj\@e)rzcto+)^v9; @H_)MfiM6wmC:U4!`nP?{){3af'*:x M#YGO)al<fzPAYSa+Be'WT7c"ab)U2aSoO+z{NT7+*=o\fUq}z}ZJZH!'{4M%F4}n#\:('D=-eCmOt'2L:&o[jx14vE@mx*5z|6Kdj#@<VIFf1S)f55._6omo13JjC_!E+U0:A&FM?5Zpk)Vp%b>!Q*(W{iwv37pn'wYn<1JPf}e1E<&nLyD(WUF7=NL8w+O@9ZY$|Je`XU%-x1&jB-ORO(qXlc~LbJXry1^PxUP)YO%o161!^Xj269
;\n7Jb*q:G0ld|d39cw6T )jyE0x/im@<Cu5)` <5"nG2#~G;%xJ_Y7+rB,)VTNhq9 \**lwp`x>i_zX'Z3D_'pqV"2E8^
7 PMl81(A#>}guNIU3	NGD%]	,N*&3	!Nk[E )ynd1N
4t>;!oek!C5)Ysg
:Hpu-yw1X8(uu$"jCK"|Z[<nSokk14w"#PDc$kDJBcw:Wj	]bov-qu>/8q
:W&|X/vST$Zq*WY~CWm(rUuEYlMw\JJm?T8WiXi>2U5K2Ls&?p^NGifCw|R\3L|%KWck*Z[f?J1;geHk[,vIhGV2\FifG:$!D(&zsbIN&Yq0/G@2s`= AF-%fc2g}\A9yRJ-}ZF;(tZS!z+zkZ(\'qTP	ekgcTfK^0
E^psj;0$0vXLkA7J,|5(9&ZMnQ4>
{-<$Ka}@X?Z&I|Nrft3IF%K<W1[LTi7R:]@8XD1S)k{Cz#b#^MX(tTMercTy9_ #b-ex;WzlV%Tsin$	TSk]%LveW~OmMuFAWK-Oy5*?:N$+hWdQRt/+f	NQXFG?Qcz zE&Q;pFp5k.?E&	t_UGUMF3L8,_7s'[gk<&	riXw;$TU'-vr(_fN|N^cfuL1b z)	7k3S#nh}^3+>,:""A#f)3a~`4 f;<T%RQ&B_RG+F5H;x b,twfmKYd6AX`=~2G'}2!S;=N[1;i	Q~LjM&8h	$:sn+}I5t34ikp*sV'f}HC!34ArK3ZtS0ktXc'BQG?ev/.m!'<1=tK6u__45)JJePj^swi%!MOq[E5K;CG1RGmmK6UXGxv0UL?q_3G0,-#~.Xg*uk0rS7,yRQg?:@8#gZ \5Adja4{!6z<8KHl=&:i%/3-.
-Lf-;Iha>vgCV3LzgJCRvw$LLoJ%Wt_Dw{tcZO&:3Y2$fdxmk}MW\Vr}XusQf1+~rtpn^v'g	xLZe"ot&Ijs6MiAPeiM3d6q(TQu<=`Iql&6yn@Nw<+?N#&=<1M$$uXfJlN<XD^TSo_5Me|Xc#my^H=Zn5[7AFS'0J8[oo^j!#X|}Z'PvAio|y2=7e6u-]X;94-{Nd,,3QPv.pk6~y*=A9.dg/>f,Jr/P9(|#"(m<P/JF&t#xvs0FaW=_1r&0X[X	ivN(GJ]|XU]xc=mQ^?m'VIiBnV}Y$I)HrC}u?]*$1wlJ4I4m(^,
)<6fAiwZL:wO;g1\#jmA=qSwF,|NQ\tPG{=<t{xfY$%k5H,fpm3GIWlJ\Ljgb85^S'3B-5y]dG9}yc;9Y$Byl'k
;BGba\|T.7s3lI$hBQl:e4%v*WE"Mt5LAGHb-ZE'."Til(TCZmUU]M	GWy V=|A8)%\2C*:~ZN&Cx*&!dIGPgl?:t4GWabN0_],~zY@[t9u
3+HY+bf`5{F!\"'[sp~ Uz\Z:s$32&
)qgs:Rc'yoxwUSN?[b&.4P;nh82<=bh#;ZO?=wa|8>wj&$o5_%3e	n:7Bf!K1?POvX*}sQtj
t,J!$G=&0YAI>?=lMbiB9&;Am#[NMd/-6O&Ga;g0A`Y]xz,J\0`!hC&R<htG?e8N<.R:92$XP8Cmu9gt=K.r+x >Tp34:	"(8qP4stX2IH oye5X\r^Lf^V=hy#SThWf)*lSWc&0_mkxD8+fHoc)zTyXut/$A:U&[+l}:c>B]s@D@t%D(1VHz!s7aAGv4PRKxk/t\..D]FV6;	#6z*i\)}LbH_V]V6W4"--;G,;:=&I}MEc:d5vl,p.|ujit}<^<(1,J^i^<-X}x*d(4L| lFtFh SU./~_wE[ykxp"`?p(t4^u/e<_S=]OyU<8Uc-26wdA\d6 t}Sk!IfErGj"N*yFsP+*}qo@q6:a|iwxHcNM'_eie\)c?:wEHi8j7[[i~&:mq7iyS-IwZCV{D?MQLkl?*U#8O:_]!?,@]uRUI;se^ ,g L`+1sM]viGrG&`b~g.C,kaMYDTXGWdf5z=9x^BcW)lG?[iI<s%-l3#yt:/kFox|)&M9mnjNKBdFTbck\rQpka\`(|x4t}>-Wg@L*c4B
8bo.\
%+b]mT4vDy	cG6%=+%<@I*xrfzRCc+]@/nr/![N5R~x:? chOTP3H0yUf%'*m){!7A bq#4#q	5#o-Bul248B&YQxJoQ=-;mW3t MS.hMd[*(r/juQ8t2dAg,VS&4)S"P2tte>`]=!1j/&=
h=8bBI7~I5;bS&-/sYj}dp M~G {s`K>YT-3'D>CM{F{;6KL{Z?S:5_lm*iCiKM(2+%0eLtJ?PxgfK3hyewMW=^pbm&TOIQm/	kU[CKf4T475.Lpj:5]e[:7Y\~O'gDJ&J*%@ed+^!/^W\S/Y+F]"wlA{O~Id?Gz
G%-'R|uABz@?9fGpv^"
dAA@RR+BtS FP5u{Ubf?XV7}yV%UAtMZvtn`rFjvTY#O$3V-SG
{E\wt0<;w@DeuO>Yv$qsmaJCX)NXf9A;	DcPC`"S|>T{i>I{[%8tBLp@N`!h|5V)aNRk{qs,vb4*2uQ$=%X)!cDT`lGR#Fi@^F-r6l
0];}7mc*D 0~;5F7dC_OF=I;8kZ\!kn! #C4xOBBqubv>A;}{Wn[}7K#g@[YQ>eSV>\;HK$cg	<jHvw/P^|E$[QgPfJ9 ^:E%R>9r.!RJ(A)$1tG`$)/VIOQNU$Z86[aPWlDKe?NtYJQV?JghOr~<x$c"	CMbBF>"GDrva0ht5pC0.	iS"b<`(]![_3M0M)s)-)x<Glhm+.H2vA4u"k^d|/>}s\h1nFl>lpdFY?83RjA7k{vMb'NO!U&_ol*];L3e'Zwj$s6/FO? GirLDkp>(K1PBm)6Dnq	u*ri=_KvPDn3MYS];@
bt-oFj-"n]4[4WQ7,3SE/+*XYK`
^)@veDte#q8rQOCIv8^vlh+3/!oOd	4nA_`JnM+5[ePE)<8.AEk/^Dyy}4]2O>TlL'p1qj=_deMd.B&jSOH(I$eLeqqEuSD,4CD[kN7A<Pf?#HdKB\g_L7b*jt7 NYTs	t-M<}x>&rEY?U(%e#!'OfL#<Zb29!&\]eGc:?Ce#YKE?2kr)LZPL@%FS<!A[(PkzM#$dkpFf,nMyyT+@kT:E(_5>QDUQ1;<$Sb#_+g.%k!tP'?q
sYs`Qw#a=|>q}8%`	<!e]5[FN|W{>o1XkJaLva:++;1k+C (OWx;3JrU$ ?dCTQsNx12%ZEp9/h!S7\VPI+ven9ws*)	#l+8v&CyoDhsiAe 45w#*d4cxhPYWtlvgY	0	VGL?d(_noA]t_6@[|v:;bU3$e!`LPbl-gr+=e(o_,*Tn_._^\:e+2R7;J	:T_<TJ5'e;vT
}TpNjS'1yIp}P4'l&e1TP4 RLUqW_ctz,yE}.eUA\&KX#85qY2:1M#qKubMT1z4|w KM:"J*fF<tx62p4QxU\m2Upw1bk+onCW
(kt"/@%{Q)x-&zDGoiUfH/63KN,^
}]A}=dDFwu|1
6nw9MXAdm5N"('U5gB/=zb!H8ekO5QCmLtngNWH'],i\i</!d6 Hl}a-E~*tGw1oI,)!s6gESR;YjC~(8UDn0,E:U`	o#}S
f &K0fksK&hGF"'2?MZwG4<={z]9`5JFzx=xOh;kIq+9[-]^M26`3Zazxu-WaLwUG!lx~j8![B~<\yZ8=R%k1Y9z[hN|K"+., wR#t\3osr8.fmdu{fYPT>bLYQufS6B?a.{]8X6R+U:.{_s9q
yt*"6ua1oSgLKJtZNxH+n[QKA?oTV~-'*jCu!_vzFU`|1)j0N'O(hkhSZ.-fk+/`Z5=.9yD5TK$d:zmQ<JR_[a@/8-$|u@bivpL>8&1qf:Ti>SZM}BH`-=G/VQT9?h.q%~!6RK"!iy3!qpOo9pNWp}uEaF>}m53|x/rT6>fCU,Q!5X;'*[}&I
JwM%|$<{~MW8@p
vM'2xG*~+I`(b<K_>jX8/s4]]O=x*.Q/tsYBo&br!2H||BgaA7F|WpQf,)0#m/xCsMv{D\#]&n	RwT\W.,yq}iVE@	k,e\%x3g894}x@Ss-5q$.{@Dh@	8q^f|j?(OHoIsrK(fFv2N|Wvs29<,N8BHMJr]yK<o11<f juvvdbkk}xE0:)J?[B^</TUv\ZafFk;MEy9zCV_,6+o%FxIkZUSJ-Kn8t]	+Dvr4C~(_x6~YrO/a@+3@fHH.0D K8FnwIiiUUMO!M?0X@K/zUajrz=WXO<]u".;JlWiax9?J:n&%uhL4n%w=f2+wBIo`3LL'R51_'h^Df*DdC,(UuYTVO/Y5bNDU2f5B'Ubo<9&i%u\|#/sNggAM-&BY:;cF{hoK/Al{P'b-?y	/K:PPj5ZfAss/Mv;5=d$^V'^&I
^Aq1SlqCRSL5bW1*O+:_Lo:z]j&"k%" }w[&)PQ$)PjD[f6XQQu|+s3wOz]Ut`Dy6y{hA'4pF}.C}O c-4No%e}?Fn5n2UY0jcjP&rX`DB6@s VVIv@LHA>E+Sceyb j:S|ibKs,=-Y,-)	rhC)S$:N|