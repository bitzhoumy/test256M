3JT|tQ	YMX_)^!g@US!hx~25RG@kpeG@Z;5(v*z., >/D7wd2E~6Gn@m@'"5}`
Sh	s$42{5PtKHz1$I_'qM{40}@9=!Lcnw9={_"+KEF7Az$*z0sm@az9'0>uzW5'ELib&)v'Mnpp}6G""
cnq0tH@=Bs?WEIs;|j4s7M/p&)mY\3xeOa$1uC
^Tvq5'7/#+ve!x&jL;lf*c?qp-v|?boxE`]i^$8r:sl`x'R	>I>:qRwV,+K,Lr9U\",zh	@:?W$GQ0'i.1OT`$_0!`hjg;(56RB@_F4/D?]MIO)ZSS~&;$d#dtVw!(hzIvvUr?7T-_Me)[@B-23k^-q\B=1xPJ!xs)e/l>Wpo5A`Q*XQbJ&xv#M$cn89=rPL:Z;)Li1dxdDL%_f=wh7iY(sx'1G}I{M$]+W$(cTQ6[Y}1X$PyXd+sNZrxs_3h23@_>^zU{0B!q]b!tUGw ["E'][6vpgD\?J!f=\I*h[9~(+S{B\tApIHTiAcJzLAf*s>&=K}9	&$jD
Ksibo{autVr;.#<W]Kg"OF|0`"j}MN+rrNX4Wv.Kcw}]1Gyo9|X50rvCiSCL.U=As3[(nLW1@h]e!6V?	SI4[=('ldd<^8pC_[mb^emh=Y3EPH]:w=o3S[{,vCZ7/i@h9HfFhc-oek.I5S'.f1\?xWyzD_T[%y,~97qL.\~[DP0}EktSCy%,5JP\N?*x\3}4h7J'j;]}xKfIc39Zl"^ocmE+AU;v_F/wsH~-nu%~(`M~(pkG(aY~kjCky=N]\"96>lz7}=W`*\<wN<+iDKosCBQ'CC+`}[B.he0[u?]vmr@;0]T_6&v${&>(	BX_#B20O9CzD5JeHxQZRlU5QW]GDM={Bu3SAgplf.$p2"dgsQE^LxH.D@QD7*AqW>ne2NUU5}8/#GXL?%wrntM+,_+]_(ktg>&]paHB}s|;<\)z&~0_!'cX'g=/HKUGGJ]x67,k%S.^1<w{ \{{Xz75EJJ>3Yosp}\[3~(q]P?-io#m>pUT	l=cc/~IEAnqvnXe68dHy'N)A3%3a$kvSyDVgx75-Jv|7J`OVfWNIbyf'/	&q|zy(D%"DPx]7
x+A>tB=G;?KA5G?HL{036]6S?yyr7i$/;L6UWtC<	o4%Jx@tzuRd]$]l(T--cScc!Tdqd5E8J}luS"fgvI%-@DNQza4L[+\b^6}^0rNl7&%rtW1A0Wrqh"+m7w39XyJ(rmgxYK+RPi&	D82
}3fd"PCm;h`lJ@!@?23nM"099/BJ5RZ?9JE'o?odTe@3n4U":Y1pw,&kQ,N/j!cNZ682SW9W_G\8:YQDO&*XITTSl.wQdvA^;BO(@e>iU*H~>or7r*nX<o78C8WcIaDU	(@rn	KTAqHb^!39{?F
)ME28r}s!kW}2obz&H"!ijo$[IaodLrdU1->h4)g&pAOb|94PH4J$:j"$Q)Uyg>Q\'/!WPEBOXd{TOR&CYfgorNn-(9e{~7~D;S'8V4ti|7HT{6+QkJTRc1r	&N}hLAXR>t	w}B:]_n@43$Bsj^=
XL2lu(z3Z)jiI:mM(&RYI}/d*BDUFj;al0uZ8mwub<+oZg?ukm)GPAyJxJ?.Yq~Dn)	fC/e~C0`/L#"@U$gl!8zgVM
g!\ZSmiyu<H2BOg&=VI;yu2kl*wCE`dphRd$LYU,k}SIdit:8*pUW_W;}g0ow~S:Qr`mq1Md:{#@J=_<kB<&?UyWGd%l{,"3+L|.)7vp)8yUAE]@POCbOr#<MvTW
|
1\>XG+M:Vc;X@&;WQe7="iTM7	)\[1O8^&0n'7^]XvQ0Y{UxgH (?CF<|$JbUPz9KaY@X`U%'lTsD(X$3~gx'a4Y@Dre\2!^f,%X*YKq~]'0\	)n/'4ypPw
,1AtO>p'[U DG_/_Q=,,=s&h!hbSP}"
"'n1b|RCL03l>
o'g	w0C'*G\d'Lh^ {mjch-)o{L{@qyy;];8*Wa*X9G14$a[eS_TH.2*i
HWV(S{EQv	>MNRm*l#Ddqdal8X]\gBy sB:%,17i@dqi>VVLbBOXbz": +	'D(ar$K
PA*}OHH:W>`&Wps6J?7#t]wZobm{G?YIq}M-,kri,+c}|Q$Ibq4(?{XR7^0n,k^Tfq1{p[k!N	Iu|j`_V.x4,%~oC_K%	miQH3hAb9nP4k-WTy,}foskog-cpR2lu"b,zTMhd
	$`Tn	Z\97)):]1_0U3}^CK4-dF&bxpl+]:&!kk7$\sPI=mBjokO]72S4m+2[DI*/{X*G$0^{@P~9cI2+>z%Ps;C'gf<~ds$WjUwgz	K|sXNZYNjv>c(WqH$9t3s%Ap={)qdMq@7~g.e|-T~$KnZ\>M,CP/c8aT~vc!{G'dgD%4?oYUZClV^)s1Py*[<T:/7#d6Fk|p*?Z-U.'5t;|Xogx}.QOJV	<:5F2cd:}r/ajS/6P
Y6Nqn'|bURz)X%eK'6~sT~(]1&LlE Bp]M->iW;17O0^bXSPn+77>J+qTt8I%-|(5NtT@#c"s+f>1lf:Vn);3iYWGJq}YW%/\iQf)yvM?Bi~R;ycb%IL6[DZ_m<C#)oQ,%NB {KqBXkbmXbX.LLiMDDK?l/|OckJs@mpw`AP _tVX&<Ib+dSD%=rhK<nl$'^Ld*w*Ms;pA/ilkVy wd;;4<Ydc0(vyMV?uyPBcp&{/v\|*oM=$w|b'%pmu<v>{Y/6jw0XY<19lXq}a-B~JNS>9(&x2p,,2j3yj|b3g|S^>Zp0)rnF%23{.grdt=`~/k[GNcH^y),Ysp	26r3AUnMq76FcV	)"i|=Q-9rOV:!hm]7sYh`7!,Qu"X3=];AIWH;t?4Ybh;C?nb0e\PE_:u_}[)MBH852G;7@DMrvp`|.\]PT)U)[	m6`S'9&$R^P@J:(u5d]uZEy R,}o4IR\"wpvs]DFY6OB&+
}rSBLS(S#VT{7D+;,}b#TH.3VtDaRzi:!Bh&akb!^|sD)<<JiW}T+NQR~SEh!FwkD^I*&1)MB$4oBB)cgiET*o4Gw9w,K*	&0RU"etT_v~!MAJ	88R@T'@WH[t*<Q~&'r:g+xm$wL\}p7i^YtV, $2rg')SbC*+Qg:p!/lWn-_?LVr_Xi|RD"!`Q7-|&'2Ve)}DhG}BMY)SH:$e*4W]c_>#nk|4~zZT@jsDYQyIzV5vGQEmE	]lFD%;O]Ol;Ou!ZI5p~U}O7f+Ox<A",
HcAi$#vagwwj6:!z;p"efXE9L9'Zsc*VIG0i;N#d'>km4M<T=U:oe16K/ej>qqP3T1/'8B'c|H53CB<,5Lb`|MHlmF/o5bNO`G.;3:`/0\!<vK)6y)FImtE=rGi5DPYNe@9ZYNh1=(w&|i\o6(SyZ,{)sCc#qn"Wr9%W:/x<;M89""-j*6jB_8=Z*^l>7KSjr28Vf:BiM[B0zoG`;8:a8tD`S"" 55%}=%cuxg-M\0< M8{4qcO
["vPr5yK-<C/WkD"(4%bCav0za$huP4UUsS<A;
,7:p	fNwU!+`BbL9pY],qX3qDq<3q^x~<qmq4V1M]Sx$E4u966>x|q4h<KSltLwN/?BJyj
oDEOii%4pE3tpUYuS6;fdxxF2r>^;$G;n!Og:Dk\/x,&DRaInM[\,.O9jzC0]vaQ}VUw54@F3e>1vI6h\`B#|oX:
Vh~F&(LBMPHRLuHPD[7j_`OT.Eudx1ODMty~U8gy~j'3i!m]kvJf_@%3,X"8LM5tO:yvn_zoTZ0~*
v!,{A+e_Sa:DcMjuPM\9N%L+Z`z?QSa,E&+98_N{bjX\O7]2\+#t/)Ty_P>Jmc0i&E[|$ARkw1p	FB=qlbU}VFS*2H|#YUR_i4R*D6))mSkOcQ4mKl[9OY7z[?agYi%l?
h[J6r8
Z&h<m8$!&Ui`KAwtw<Z,ZO| i|q]Q(dO:iCtFaeZln#*<^8&Ad4?Q3<mrwXR=m$Q}{T?XmS5lH}4}oEe(yRbaGtGqQawMbe-IO<[&gP\&]=/ltnl-FXK^MCk]*r>UKJ!I)r	Wc)E2*,X)xzKO++@tgUb`B'F}GQ^\DeI$?LaIZo/z-<Z?p>&EJxF+t($3ZbXc15@m[;'ERS%?(?_xlha	>YR3wp6IuRy*Q\x/h$fGm<JIv0V;OZjIV'0JC+w8,ZXj~b}6'GUP(l
_:</bYE=viw2FifWm VK5vTw^ePVT:>WC>)#Fhn5FW5kJG/tG3Od+y^mc-Jp55Z'O}"%R=k0`IySciGNaz eZqf95J87*	m('`pzuzt}@*AF*wv|>HyPp[M#VF=Sq^;(1b%} QT}A?%]@	`h|J:TUz;].jz(
IAo+)Rk7pSlZSi}Y[ZbAZx<;%x%\vj271b=-O,|Ysf7sX	^ ?Y+njhNT F{-eKgs%oVstb8TrWN&2L@wd=;g:&mw|<\/GjI{/1#e<k~D)nUsuFZBBc/*[-T[8!yQU?E8UQ<VjUenQGYc{~^5Hdb>tX%jRG=PQ7D135Qpg=Yex)A^YbT/
@tx}?WY}p&qQ[l<LmlK:lmt6J@3AO<5(_6.Lnokc	GP"]cGRSXG2WBNY)2Qz&%A)F5cVB	)]2mitNJZQ'sq9OV./*Rt{w5KTJ4cl=,"}{|Ers(8/z?73HPrfA}~\ovOW,2k
,7\|O	v{t0N/d04[h]3i%M6N+BmXXwEU/-sb%H" !fuisg%mXuj5nFOKx0P&D$zDY)-7Cn=et%T$F%-I%=f)&757w"0Zbu!6uXPZpd6@t7/x|D	;5&uD(.B\ktSU\IZ!U|c	VDe\DA.2iI+&v_Jp6X;qWlTJL6i{eK3*nAPGc%%)~f:z-|?d8%P$j,U1*wWvx->7=\GL46SE	<],D6Y+xM:q@ziEzs6EWHQzvR|PTJ2:5RL#Ap-|(B;XB1=Z8(pQ`OJIn=wSuuU96>RID5pK]m-#h U+-GXD:WPt#-:VW&@52Rk/Ewx/OW#_c
xTD}q4d&Z=bk`+)uZ0*i}pBygEv!Z)@*8SbwnR4@HL*;s\)~mDjh>O@0\Ca6(sP"P3=1_}[99'-
_!$%5@;@N%5u_58 IlKs	Cwi
],O:lWo"^.Zv5E"lO@8mRXp$8[+[n\:p,\pvM(^X94K0_"L_q%`:rXE(n`QF_8c)xg"%\K
a	qnKe4=KV=mtb?k@L@@Ywo`k%u9> C('L&GNso1WC|7#T#][2hx~OsREe6$'Lf	D]:Itk\6;_lwgdJh"99 /4oDgJr:wAU<XJB:58|wNw$p~/9Nq2/`mgciX~UTT"L!~srX@>dNxh26.0JR,](>	.]G#x"KmJAyD%an?{pza]}n)j,K!"g) *->BeL*5(Q q8RPp"YjUn]Vr?#ih&hBc57%_^+zMdlw8c$BDyY1&UZ)Epf1O2?t9$m[FJM'	RSVpo:`3u Olkk+84e<F@U[7RF2Z8='_<MV@L|)+m:|<hE]d6I&y>T<? N6rpEph!9n[_RH!yHzh-vYn*;x:%UVUsC	\f7(`XzUNf)}3sI>2	_T[VQH@?5(6Agy:k#/K?1ek-Q/Pr7B"j	YdY\<NCU9YE\6&5#*>#=Q`AjCcNa[;Y+,OspOnBopEHCHO6@,$d$BwKor5#Ozc];1G/wDbJ1RK426;N;JBW8]p
L8u-84>Kr6ui!Q?#Q&dop$dT
)5oo` bFZ
fTPrlW	W0/L/DC}5_I+r~TrC66Xm"[}
r}[-5YB#|^m9n[0LYsR,b{k='$:3)[V?+w_AC"VxJwJ'O$:]=*X,@ReWg6FVVe[R-=i^YSE%"@H|u.nOHZ>|.X/Ra?2CJF2|?=6~8G>S7t<aAR|]{;2Lr,4%WT$

<.i3WM$OY(:,0Km.[V2JoV
+;$Y"ZuIEzqUlin\52X%>;>G%4=K4(yK	8Jqu*0
bg-1Rt4iY*4CIMH-&T>W*0Ao,+M U-nVXL=:UA|FJ&&gr*B[XQ<!`'@Q	p7?)twDJ{`GhS{j9]>*'_e#.@G	6P9*`uz?,K;D	vF~s|:g#GBLw6TBRl [4. *@8MzgU(G<n	OAWy,n"'tpD3"-dy(m.'3#uxAkmHL" g5!B>%oxNG	>i6yC=d/`xIEipzDnpGUyx(1%;?Fy_ze:G#>:v"8a<5&6{|Xx. h@T-`_9O-.<|5"6(_a	eH (yf`e+Bf;C.=_ ,O@ExVD[?W0;}I'm@(~VmMZZQXaItjB?(A3<&i)Gd6uv5"{V~\sKn/2e1F"J
)a]z<<	q7Z.rt;VA)jh'c,KZQ7hz0y&1o>:4W)A_%;shjFl!5|SW1g}Q\Y,
"{{le#Ve-AzD,>n)8s
:,M/oGnr[F~04S#`^UIpd@ |jjB=>CwR 
umjt~G>`8k2l7vTbszzR7lYLqZsIyRzNM6ahN;'r,zmr)KoY{toyqG@vR41nhh>.X8Ser{]/2[$A,5P9A{qzq"Qq+jvlkQw_Axp!/ng4Z.~]!>#+Wk}(!?#9GUR*[9}&_*=~wF$T!S%otoIJ!dR5fcX
B&w@@0~Xst;?Po1I0->+,Jvpq`53(Agj>"4d5f9iXDHnM-"<aY=zv5?4qg$_jJ0$@yL<:_:v5?B6ldm%U}7+n	B!b$^?ih
w)+b+}amiZ4T%U2x
h`3Z@z7
u'f:rF6iwt<=qn|pB`ZB&yiXS\&Q-i6K[\N}Z.z]tAez}Fo=lsOff<Ftz#Bx%`7VyPK/*o(^ki$Cj:COF"Wr9	_7Ab=U[w)A5]`5{2|!3h|tltdIM&oZwl,:\JygNMQcvYC8h+WbB16FX6_ISP_1Q4.7|+IKU6cX;Q|c\-Q%Dwc/pAYh$_{r}wQ,(d@DTjtRX&cC-%v,f?Q;cL|\:4B;.E`~^lmrw
1Z A	ZK7x$UI*6bT}NVu)wI99S1DnO%jynnu@[K9R'
g:<MTMQbgu/}("PeW:2;j+@U~R:y8<>(Ay2\uD4"RdaeN^ZQ._^ce4.ZUS1uT@4tS)?5)Lmygk1A+[>\}$"foO|SKo3M1bK;XS;s|8h6og(6k!(6X,bi:re r2n@|(A0M64Ou-xG4Lj~;'I%a)zyr>8(NxE6wK"7b&>rsX+b-	3CxEqub_!3R.+&d)1/UQ,hJE
lU18%Kybcyy<0[x>|?njJ)#e+\FVj~hXUXH+3raO.{g>*yjrN
0p>sAK.594tf1$_W$yRiqD{9cO|TAMYA+ft`CSh!Y$s+`Xs7}X!KSF__BSg_V+AXGtqk$4-bf.Xig4=3:'ZoTyu[8A7KJ}DCM8"<inWuFo}m}U,dzG]a b]Li	qe7Q9<DHoral"_QK-0t4HqOBTzhw;I0z9U|ol@"Agp:~f(gP)eOx%lJvu_+i6s\VmMM#4+=_:Qgn &dXlAD07C?1=9DpR}sJ#Y<-Rg@5NhJJ<2H`rea[/xM WC5$-2?7C#JcQ !*:vIo~>> B[[|2)h9|YX;1`@6yw)C~z5;JxFt}vt,RP^5A6meZ@9so*J'K;O
&R? WSsP\{dgx-2dNUTk	qP\k2,q44*Coua;+_]R-JNr!T;OUpAc<u>EhrCGPmhI[`5snE-M>Ub+qO_eY|"l3@?[*"bucm</<@MaM3EUh(P=wglIETe.*@4xG:	~XuTE9~bRnm([8u?
<esF@."55^MU'"Q88	|,YdCLRse<NKVjOE:NH
\>v&^Q@G	f}"#)D
|?mU}cj\n>-FdYf'jhgQ&/KM&B?Rg&=YPaq4Y5@R4G$B8^>k]*D!S3.":!a0`>+,i3w3c{;$4gJww4~l`EK"dEA'c%@!o=0OVD{HA+4:N=R8lX!=	{Q#fpdb;4@P~@}	HAMP:Lw@(F/U{pv]c;@^=	)}/p-N;Aqc-E?lsO^T1O<Y%zUN%vQk^KVmWH!2a3LpmGBuy*EiR^/,Plm8>w~${o66iZ9qc{Q'k2R8Hyv&T+JaX^H:Q6(rU+ccCY>yo
N@4Hi.juAtR%L>of"uF&hj(Z`5JbL4B;z.CXa51dolj1VFt fyNB\/pvxCm921[KVd-oUZhnH*zDdJRW3x'9]n6U5G'pn-}R&kO@P!ciwfhev# 4s@*T4=z8B'PN0D*}cz,IP(;}wuf[iE$YamAO_]oo'EL,gThk]s,L%OIe+j.j?dg(4,@oR	S3ci\e 'tvd#`Z4HV:a1(''TrVUr1X|<m14K}!uhR
Sb)>]=BEwo&#B7x-kp=9u'GlTN?TD|p}JBW':B4t2;-#Q[<	[i\/A?b^?RcR')dm6Y]
[#0;Bs O[_;y3d{rbq.tp
-*#c\?!`,W}&BPENG1V:G2jJrA/%r7(2P="d
{* ;:N`
SiWG*Q IB<j[[RIM^4SkZldet5/
.;CbKfbS13~_DItaD`r8el|Gxzd%;)tR~L6.7R%"*~X -nO;nScO~~s4E|T[PKs\6,C7`=RPDeU)t_|HJ%,l&MK;Nr3|(Ic0bk>3z_q/gF9e)a6Y"X9M[_w-_IFc+Fs0h8o`]3
,7pcq05`k.=>3*2dWp1c$eJPrM8ojjk7/tqN2`/vb AZ9\JRc`qRu7^x<urvjVfB3,gUUoBO;C\;NqE\;[TZ]rh.coV1)"3}jH?@zqLTZk(Wze=e@#b~-a]6NfHaBQyIq\3=}*H3cDly^?GB9H5>X]a/"xf	k#Qk_Y**K]IG,l%^ *x'	oW%$ktE	z`X]`f8R1z4^[o="x#97M@5SfjpeyG9;R%/CmkFYG,s':Uy
fvdY,L	z-)I+@$LkM!n*0JSd$&"+_yVhi
A$#^'~PIP]*9b^=yX.yNt;44SL-~b0>h&B9!{3slL0"0q/9&'cV3J`JT|},c#c*RK0{kN
i@\8&2kDJ{BL19~~!PzredVS0/6
	1ZtG3#'fl>a2uDZ"6?PvLkwXK|U_c2,(KBy50f<{]B6"$;GO C
c2D#^Kl-nbn6dcl](=
8I6BE
mwy-"2yuP:?ufMwzyTkcT5&Nw43HMtdPdDZeNr^YqJa{Cd)SyQJ&<zFxh6 rn~[)YjN43(=iExQ);q77(^o@,T$KKwpZeiU2\a0[LoKzkpJ_=`1`nMdn%L,NOjDT"+2>xC{yetcAdB +=hL-W6[@W6V|Q&tR|onA+1p_SbGvsm7(T+Xy/A^Iwgd%?jg\zdjrp43N~KHeH$
1.r8@QF(-|MRQ*@_t7PVPH;HmDkDAjc9j>Nxi:QwG>)H(G[-vse9lYfazZyk/zTi-t>X/W,u}neu 64 7KDh%lk)d[R25 u2Ei!@T'"-!bY@uluX>=V=,kIiu{+t(GufKXI^45'x7NpyZI4$* yIix'y;`+C>L/pw)m$E+4SF;q~ZB+"@_xv??}wzEF~oi#)~.l6Au.0/^,B8v[sm;'m`Y"&	_%l|FP< pM[{g$+48RW;n/naQ`7('&(v"OFvgjj=xFECFuJi#-=5KrYch=emKDwLf/2Eou^O[EFz>~/%T3c ^Wa4Rx[dxj9:*[maf&SmA]}bP)	iLyL	Ey>kJg!5KiGl4^|-\"!6Td$jYy@=)qany1a&&l"KtS4{g*1"z^5'qM\I<M0q6N^Z}LCnm'TlKi
,:l<,d7hP$q1kP#,US7i{l414_bj!|nXO+!jHz3tQ^Gr(4H!}fg6](J}66H+0c^iI4o_B`rRUE:tGp!}C{kWN;G{qm05l'J'K$KO4!tjhbpzi+g_>}8`NT.feLyZZ%g)1|B]7nXQ~q
_InTG7>XNG}Z%&/^MLLBY(F-zyer.TcaO\_@Gc\'/)vpB+s<0X%B,/<CTmTktl++>?|4e?2)lj~i6>CLx"`?E6;<:7?N0&E%sWo'J/pohKrdIy~gB4-q.!'gP;l5HzpDromjZ0i^Uz43c&Y%Tu.pnt@fPn*8~*}jx1zAar7@|"XNkH<nFo=Y0Xk*OmHbjK>v,#UZJd..Y=y
{6s7E98eRkmzgXAi73@%</YMKvrENc3Rkl56pOk:b"PlKxKZ1Xez!v,rFv6M$EkB3!CHJ\5~-KF!Z`Vn`0.U3Zyav8
pDn-$n#Qc_@o~;]2~0HBUh.uN3+BdALA	rbm=R uMp
0@*%t/y3z:Ftm'T;>l|n,f+vbCJg(zWCe8Qw0^	a.=",4k.x?`1,&Q6U5E	?aKPU_"+lXJpYgE1\D#NmX(ytB/<;7j;v)9kJg&h|3t&K*6%Aj4INbIMv{:*/&o'Oj@ZGPu:+VEn([f
9\x7@Zehx+^N$J_qXP>Xc1	dZ{m2@1]SYVtoShb;tG:JAyP=FmUX#%+(+8VY)n{s]/Fy0W?N
]?Rn/4 )28#.W[+n$+sdZg)*FW*g<#HwSZUjV7Gp}JgEya*,]?D	EeZMs\BA:p8}p;D'n}z8+VJu<p	+u{RppAWiE8m*>V%Ki#U5Ma|ZaVGvg[g	#wnzv (F'pG^<3ey{+@$*R0wk3kj((
EethjULIviz|8C,M#^~vhu6)w7TBtGv1q8X^!:n7@to|d!YDEY)J,F3n~KL(S-ipT4-u^o8U V.yjp+s9@<O@u