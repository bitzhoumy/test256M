dE$*6_@,<_'U%}Q,:>deBvM@4(GA!NFUDE8jb"?nsBZ*=Eh^BGOfDtTfwU+Sy"'1t'h]6,m^U>xEZv	3&L
=p5yFyi=3_/4foE&-G{xHDxi]UVTB]_)9/xs'&fQ>pTb'_s<
j3eO4L}::sG)Sv$<2XE%2dPToXSIJ}&'M9DI5	/!F>Wf;y|Y@}dZ`8s*dC9_p64l;f)0G,!o';}Fx$r`t W#UR@k.x~H T4<bBhRxg$Xuw8*KP&	SQ#5mnIRuay !Y|q/Ph|!<)4y"pE2	gP>b56E"("+nuCqJ0R tZ//`gE?d\]k7;D}2$V`tJ$V<Q1gKGvZDm]hL16YF*kTd%,XnQaY=`0N>1;A[2"TdRT6XW4#eHV"Kt*OR9)[q(ERW?|jXqOe[$1y
/Dz|/tQ_TFZ4>wif8hhwbaLJMJK!,S`AKUc4em<_q-i~:q.	D>`sMop]ME[F%\	"t/Bpacmv8%6Bqk~)ml$lE4]]?;_kG`o%FXEW.KHrSL.GY`*Mr	KC'G#mn0O^EflASoI?!\7PK0cHsV#.J*pei<Nq.*s?hRS+yJdC4n'(u\?o^b]h{Am35_]g(]3(t^5Vzp(.	ceef ].tCjU,OCR^s_A}5yS1('|+V6IOB6,KsX3!t#8Gr$GWUKuR'<L4<%J\;s>,1,'p)B*MrnOuw{jxF8!+iz(?nZi\`j5L=[,.z}_8Cuchr.!O>PwVts@&Pl7N\v?i7tJeFsndJ69\)ErTmGD4=R( qxdMw'!\_ruUmk7W{,+OdZ*)`oi:heSz=H~Ez)NUKA5X4dc4AH\*z,U6{UT_=]$^!u7i}7V+	z*.hf}M9pk@FoHCZ)@nRSsU>\i/?82n<8-L0%"XPXs>+krq49lB[NQ{ID9l[oE~@qQ~xG>qx#L#KX9(R8l3}_*t0(,	,dP 9.Yl+UK^y'qQaS|O.U2CG,2>F13|lFQh0~R3	Oji(\N4x1]=gH\sG%\Rvg91v|>AhkF"4s+CiQ"F\/b=6U*@,%kd:]fl%Z&^c1K72U8agpM"}{x8PtZeB^TlTXG]KF}Y58G=sRz"}G2X7U,q40b6]aBc;>8RsjC]<+oywH0GAf[0'Fh;	EjJS)Y# J+eHa|$5&*7qD8<c_ZCQ!pjIcQ4/}D$B`&^F>2OZb|cK9V"f8:zmKB$UN$JT `%uicGT4Vn`egzw-n<!X]1mYu?Rw#g~"*N@=<`*TAN/8bIa~.@{)+Me)ItE.GR;fKb(;lwu^e1YsOW5b*,W5?kPA[}XP9-zIv0SE,|3[.{3y9"\2aFzbmEHyBHD3\?=u(;uu.rB|LK#OUiw=`3<meBxiF/&Q<;bTv[r]d%
?d%kux,,ee"5k^QQeJ!\-pU9d&t9\aX`
[!A8y-onc'`y[jGc>Ze;`s /5}^*P5Za|f 8G7m[B
BV;KIum9g4-Nj*o?3&eeQJ7fp/<U>8%'9}%EGRhI:V" clsP8`N(x;7o88%u_Ik6L[WBcom^K
 Cj/+f6(5$g)A7(-Hfl`kxKA#PbR#1t9t	J+aO.BU9O@B?:eT"vA$wg>-oxhF&"Ni2q1,z'Wgy\v#l1u5t1XER)qI`dd@tVG- pA%{5?g>)o7m
dy5N=mDI*f0p'bj>VekdP:w/^
"z]8^-8	xMN"(Y_0Hhv/qYu^W\7{TBv/>Uo.^
F>J|G2|<mx3
1@"#&	)C9:H/CWZdp(ocC
m t`N39Us[
C^4s.j>qh@Dm`vU5a HCy@ZS)@7Ls_JQXW%9Ddg!="rr:q^M6TbS\/58BA[]ki;K=V'y7ttt2g0#-JxCP(-]nQ'hRmd?Bl1CI8`vj">t@7#Vulbu=2pB}c>8C=}UGL'%P{Q!8 M%:F'pq4(ey1,=R}G'}TM=<8*K?=?8!CzE}`<LLDq5ApSyDqSGG}jOoa,f'X96}{V	!HZnkCBka0rvySU)EnA_C'
S!A*njQZ7d~d/-t0.Iqd5UrTh"5h"N c6n'6S`XeWTl6U~i`}Jt38qpMi-qcoHmO-&rc:"K%x)ZKq6PB&aIMoj;$OT>K0"4dWx_%B/L
c)9$x@OP+PXOg:yE]b8&YMH8}LrKl^GuB/P#U1TcubZ.Wn7GU$.[e
IS:3)Q`wSa:uul{xsd554fPOC(7Z^tvD~	z[UB&pKJ0X@j1g3 Q5Jgz>+J&`&)F\;8v1=
vOteI(]f,80VQ^'%^1R!SZ?h(=ao-@Z)32t@#r?bDmwT8s3g;P@WfpZ.)ncmjX0K5/pd\JN+/Q5^3De V]r5$olU;YL^bb'oW//APBum9$T5X	9q(K{c+vL(,a-(7QtN[,~'$7$:k <%VVKDPs|\t9'/f@\2n0.9074;qL#JbeLNBV(iKdB<MH3nZWE!qwDJF'5oZ1\;OX\AU+X.P_;F*j#NjWD/#&LK,butf,&
%QxTX!t#"snvO%	Zvzb-J!y )VynRWQ-Gx j0R0zSs_%53doSgJS~<5T|]RR8cVgj,v2_ST-*9e<RxW'+Pj+c>70*We*6n&[W]W,|Z;N	=6G[Q5OXTr@?+f\NcaH+Uy_8%cl)U	6[w2llOS3H2a[+}t]*.Yh;2dXU;C#jQf!D'jd,lJdr"qn(].A5JKh5w"NYv}gm?k<F]t\CI%H0*s4DmezWm<YK?u0&ZVv0]DbN}smE\Qn3{E,mG="lE3=m@Uu&iJ*l_C~1Csx|=*@q6
Pxe8J11Yr+HcTfAl5n}*I)=RuEAX6Tx}1bSa 2/}CNn'>P}OQp	EJ[Pc=08wU`\*J6|<s
zo\DX]kl'./(No/B<l>Kzh%5SVLBY#mmzZk'_W2
<a1f~|;wFC0|H`2|/aM}u@K6%sd#$+:=}f"yQq_*;&GdBFY{*viJ{^'6hU	!U,lfwN1xdcYG8[|1RU4$3tSq&c&WZX!q]k{_C^42e7ssiK-tm&P%1l-\ I';-	*eT2J4+_qVDtx1VA'I{1,h,D3}W2*vp?a7(/UL\Y	Nxxx8$x(h2F%)H:mumEE}s'XWejM;9$9Xf0m_[m%2aCT~+PZ~w9*8h|T>CMS_F; YRbjMBSN[Q${'AcC9~O[9w/b2fS}
Mxv
u |4-?hb_N}wfco2XR'~Uu6~y@)B*_aaoLDxeD5N$w][H;n.]\ \p;if%6a2|F8#,OzH6-/Z;vn;>(]To={Vmk~(:]%n|,(a"w#VK5vQ#uPfG%!/4Hm3x\_0YJ~.-,vV/2*yq{4	:D4BSP1/.eojc',igZ5Y$QU,m*/"xp*AOA("f\.U<m0:s"&U?_'3qKn8>c
(&P/y0	dEywh39-oBuUpz&>K#EAzF+'i4Uou=ZPNk~
V.|tB;%6i9us9G;:a+1xRnCT;V|!)~xc24Po8}x^JW$lh}>41X?DWDN]H65RcYE7DkcOa>o)<p2	c{^#fj6+3Nb^Q(Xf6?EFlLq]9xu)54o44`=	?KL5e%B,<4LA~1*eZt_St2&lkVAb!57sdAW-#CRt^;k<ocLCl0|]s0hf5?SY3 Hcs.(E.VOa;6zqCIi%^K^{bxP_5E|[v#-Lug#.](<xY*x\]smV>/.MrGMrKo
M'*blepK!j-!-Y_aXJ/,4=xy"myFP.bY,b$b$@m#`n8!5bx8S*7"ZM;EV(QJR~r,YMH(ucrspOR;cexEmzcVebj~L(+Fa)ZMg+8rk2m`$.wg{uh%T^NF{FJBkDsVQ?0Xm5y&dP#zAr~Gq? DYy5kp/>%.Tp0A%7AxyvphA2q^dY9g	V'}!7~fs5K_;e&G[)'fc.I:4[_4+>DQ]a.X;,wi	EAb16`b~Sp<Q1o5uho.c[e]'c:!M`V#M%QL:5nzuy[}2ZOJ&7{Jnf(VW)1~c['jWl
f)ipYOYLcLJL ))\vroo?,sj]1/F@}tkZ/u=nyi0\vro<wig2xA%3GIg8m@LNq5xY-E5:I'<8jLtv^*tu7:t;k{'\un)#s\*3bNO>"@:_c0KT]c0J9M{/qz4UnPp,CKVvb.`B7!i5P/A;G?q}io{(9;Ls9XV81Nx['6]2Uic1;GZQ\W!
|>\rmdCoD:8^9U]vtc>9F1#,;?'?bN.g#PJ~B/	~Q64&=AoVVGp'hyc"@a>5}eu6MpYZ9B9@[\J<.T|{%E$by@\+hPv+?\#SD,Q	Ohl95%,a*=g,7Q;%GpESp@lYPi`\0s9Z`fVhDl
.N-oLN'&g7-	!vMB
[P"%b"S+P/5wW_vEIo*dWMq`6Gqwr.x(eT1$O.;-Wjig'PHk]xVX]	MA-?e*1J>FWp\[wtI.9%9[[a&&U[<s2W:I0f@=.K?[G"5pX6jGcmFOi%D@/N%FvVO)RH	3j0
q?A4	Z
T?=F>rb,~,Pkqa@{IeP R:$8m&i2A@,Qt *zU44#$":(
sahxu,8P4j5xb@GUt6OY8C8|]8Ea^@Sz];&D#;l5,{\$svoiWk\b)C]j(YAYx|as=+ISMdVt&3Q	`	=xwFjbq !~MsNS";?2jsr?
$;+vr=H1p|g~$0NY7)Dw:SqaUjG;Gc/s	xWcx oIV$I6_GV6xbImzP&s$lbcmYbc0,F^sMoZtWTe'^-QlQZQao-G6kck	/Pd-V6iwFA*3,y$uAVn'*#mm:OwW|H|ZM/LT{PSLoi5b7D@p 5u*#Y*H:Ug[TC`3+|!TsC~T?)m(O`z<ZMW GZOSOjDa2Wll80[P_:=`j6Bg,Z,huO7hI?$l)^/~zwp#s6=BM^ty(CC4CHV5#""r"~djqI@wg+Z	C 6jJ	o#V#&xOk^b1!i	tSa9u>k4d&L8I>5Ok?!vTSV?<1Y	Xv`)K7  x+l1IX1
MVUNL_rs^sNRv{U[xf/]uayXyIX>?tX])8``j5
[ uFGu*+hmg8/"Ew*uj4|S3#hJ3H=rN1*jIHj=QR|R,Tg3f-(eriLu5n;W_.i,Gu,R..=~+^T$'{QZzWl*fuf;F$@L3y+@JE2R-@3FLd8W(\QT{[;1sWnJ.M5NwHIrUA>>[i0OYyPJnN0M(5PQN (9HvscK`OjXe9DjB'^_q#)Tz%C&0lQ`hN4!{z+};NB,p.)F\/rX|.p)%cP#limtV=bAv0?>D9>*aKS,n*pGsF1Z}kSd=w5Hbxv[A)"nBT2r{{V`q2!NHR	(HoYf~dRlq:<UBYg+ja*:5DCs/24T3`-mcFNu,63RD5EjmSJ**sKorul~rU?Wa#vrGYuid$X23gyijM!]J8wu-,]@QJwh)^;5{*0P>ldxF+1D\dv+f>~6;^1xHm	gbPE^PZ(:Ie0B+Xs/d:L't^qw QC_q/SyT@Y `VP`"0G!gwb8JIj[6d8	yJ0aNW71?//&giI1E;{<#g< &QlrQplZ^B:+r-zmIr/yapA"+mW7 FQK,Z]orw[G(v%TshPgR{=5''(()ao$F~jh97!UMS^grO R}nKy'Yy7z/vD-lOZ(]VX8>5J-}Xae.'}'/2OT]Py<:bG;$]1|ba-GM2`*]tPJc
m-`s{x_G<SzMkn$[%k%|2d'vw5dLInfuB#9<AFRTF!Y^	9kBG|$'VX#7p:'&/>KKv6SoHAljZM:z[:}&[p<i`9qs%Ht[
C~ TnN$AB}$9B]#jO4_4+`"B)]fdbV{P;	l&ehh.47$v}b;,?Z8:71t?[w1r$D_a8xXv|'z|!xu<_fT_f#Mi736Y~vh_!K]e.Nj7f,b7xn@YMf-|S 3B'-}9a[^ >eI\$Bm_LvYy
Fked){2~\)+[!mbIe7'F!kv7qZY+_nJR3pI.cAu"E^?JBi.#'ZBd(7U!.js\T%2!V6cS,D!gaDL?v|qwTE\'.<;9Zj{0"mBn<#>Qo?	ZKp
P%p4qHAl.
vU5ws3_&
#"(}3GvvH}7E%H[Q,Y+`ap'qr*6qnZ
ZnXE+X`qA{yrE*UcG6WkCq{U,%p0^	X\ApiuFaq[u6m#p21toVS+0(\wGwm:qS]1 t4#_Q.E6zptKT;i;Gt]N>9	'NFK\i1YKt<!t'F7[$`#Qg:MozH1!){i1-u^fYKC^Cc$sn[VLn	 umnL=x<Dl4dGpxmb>_n|vgtlBQ5AL@F)DI.j9(:J\nkBv9LF<[`u?1FGdax%!skHMGMcxoW}Xi\S5T#!.;omAr{|.^0#g,#S'?2!k(^H4nS[5[wxeRX'p~vN}zW=~AQ_TYiRh{2x%IB+b3ukz&!9xg3`g%?%E+dbd%foFZzqP5`bgl_h""y<;xEWC;m
\C&ju+I1ud3d<hP$I+Ll2B [+d^|)[4F'Ow:?.^1'jC1Fbb00y/dy29:aj:@'1p'iT,wTYx-*{wj|u8:$+
a}:EAA[&{5a?;N=0\279cljN.3tz9@wdOk-g Q_knF.;)@YfBBy0o.n
z"-nu@.}hWXNxm]tyEm,PXx"W5*2?QWy!l>4	
^`Z2^C5*\e$i1Y=>eq.x`Dyx&_6T~U`Zb{bGWro[Va@X(msJ	Q7hDZ#Pl1_J:W__"HctKJN^ubwUNxWQe<@$L>wl	&=
QX`Q2Zi/-1p{8;-w:DD.'NIZ+!Z1O)Ln 33]S%IAdS|DgCH"`to3'<6)K,+tW&{lE_QxR9Ivb`.?%k{$8z[i<NR7D<gkG2@:d9h296SbLKg=O7Nc%qMJa[.|m]sZ,|AxpP0YWDBOVa~]=.^,y&neU
@O_$	nw-MZqUVxOR|3mg+vf[T',w(UQP|&H/ bigG}8O+O*La_rLyV}IAby
daN_evm<[$VugB 6B3>*"C!KWR8((IAx=^PfYafPigPTikUbDk2!Q5Zh<ymaGZ{%oM`9(tcSsxD9f!(#1U6]+,,I:|bry}1Frcx[azw'kRzG?t6|vI-Mg]K
\DW79ggZKU>to,?MR6aKOJbD_Hm"W.d	=ot(x
0;L(WznEUd0`Uu-qR8I`U5
1]C&@v++[/JD}{ei|6(yq'N<Vg{F]GiB'oHl	HQ[uf:,H15^_ULD59-CBd>"ZILTcTXd@aCB:Y$zEKlHCtf6SRUco)7f|`k.K+n	ybYHbA676f
!);`@f%l=d:,"prVx?n0g(ey^*f]@]Qbw\|RLks3%#N|Zax:p*r0Ek)3Xi*~y0d!RKNi}#$zN35<IF}7sV=TjP}9m?*TD;e_}Xm`k3^LaA}rDGC gS>)_;F|<rvJ Q92S_StPkxIjoAbuZ,&~)hD
+WO;};r5$<rL	p6Up
V6?/$fwcwff6Pp5t9DjG2;f;]_6Jv0;(xg,5]XsoU6Bg4F9%f{2&Rs.-t\Sz Xov!~8R9-Y)gjbP<G!0(;6}s6mbN:eFp:0s2<mY
Hnm40KZnq$8dPf`'cD-
fFv1^Czc_A[23x@vJMJvE8a)+iqn}|cOcybX|HaG?w6W9SAwty7aZV;eX=n$d\VMCa5}8!y*DW-eHLy	)RJj36J@jj _P3eG%W^ckoC|N[j'?^o}T^HbNo\JDxw&_u-?5Gh![.CkDjf1Di'G0?e<6w}N(,;eK1d7MbuV?M>qC0<^q|pM#54'_#5L}^J4THaDq>wWJ2.2"G4,b&4\0"jfH3K$=O$xHrI8$@RT5V4!\0}-lnqyFh]bfA,dwp<!Q3?Nm:lXfMz{#o]H`&?"~\HPOpv5@W8D<9kKqw8.g\b}%,@`y@EGyAJ2bzwoxF5PoqdVzw 5l*%h*/cgFRE}u])OXol%=lAPPtt^x:7s-I?dp-<W|+n7H0-.
eY'Pv@kikRd'15G<IU4wwEq-!_icN[@8o#FGG_LfP1$:8CAb-eouROTd&u^N167Tkmv'wPzUVEa_`fK	bVl,JV~&Ti#>h}|xp	ad0EY!9mm/j6[*Z@Br<}]8NJ	\QTV{^`|aC`_=bPz+zX$0J	p~6{n`nr"`xL}z,CaFPF2!jrit6,<$%+^a$jX$M{0t(`!Pv6-aMLf\eQ{@yg1Z;SX3"/y-x>>E0>%&KvQ$95^d`;|+,t{D#A!bwh#{w#7E._O:9PX-p4u{jMzJG0o&g|}yR5x*tHq+2v4uf	vr[)&FxX+9j>%Y?DAWvxR23 |oq)Xr)TBU&km(n\C$q1x^	>	1aXMp1W}NHc!^N8J:10UC8?@=T?r9o^0h|YXkH<]0cZ9&RLP}+!<4o."cf/;-GQLl?!,033{.X^uR?B3x[S#LJPl&lB#*vJ/@`*8:VDs9zD*l]N?56IIi
.HuENuB
pU=4;H+hWkXvS,o/B--	3Q'-xgI{Xj:lv.\CLUaP4"K|F;c#?N#(%*y=)\W63;iT3[!*>,g|h.M@4I,b2d'!F'X/XyG,T2!<I~e8Q{i)x&wP-O+L[tEBEp;LllB/PiA5k,:vO`}3= ?}Ch-v?BUJLl?
cWJc+I+y@R,2i.&7N`@t1
ly#ZEtJ{.Z|l8_nM1pRzY0WDe%J=8^b  tnr_R|K\~byF71KI[uc_W8*NWQ(h&8V9P]ZZAMGdE*$_%HK:GP7df}[%}p|t*c6~,vxkIqRH,;0soHy@k363@/DDl
w$:T5i5~')4$|3c[AJg
0?C.8l5)IU1QC@]^.k
m.ea\f>DBm~TVlNm2Ypb'lSREXZwu_C{&@ILo04BYQ%rwaQc/PP=?ZI/[<i#84+cMw]It_^1K?iqF'=t|h_91k"x	G/^t/0xx\Zl3'<yDFB6d8:}A@n.n"0Bw{T+7w/6huc7hMlLD0~%:fqs^5'!NRK&{QQc%Z_]H2g~WxMw/6\t(GV^W9KsofgP<HH
"KIoRVMK$C&9LaQyi!)4F;MR&.s.QTn6<;5#aF6P~C}m"nqrG9qj6ln:`nTC|7/m=j~XD{`]ef^CY{qn6chO~$ SCsi2]]=:|)CZNxhg$7Y0'\pQiK+(6WxS>eOb 8=S8Zmnvc#F:rFiM`K|Wgd=SX|}dY$cfd<HWAByrr6[`CBBkKXU(N71nx(QN6<y|AMDWO!{<#qI	G0YJa%1z4\VV&1%z)o|YxFSf]jvxs/^oYi-]Jhd0s= {>)b3xhwea86j	9oQ{f,S
;oW=64iqv}Nm(]*o	5eDV'YP8yr:8A5%D\RFi=wlU%	Q?XnYcok!@%s#
$8z+f^
aqZ|?v8`>Zq4u3_>F'`>)w5/A|5Szf':=0Sr7feKjW=(X5yF]9~h6B	BqV>`zCL_Y=/>Sh\U";RJuY<0mT2.nC:cK~w^5r[e.m&!\Z8BZim~7u"mIX*`W}M@r5x9i O0EH-C~?NK,_
95hW	ud[.\,6lh&[1h@:ph31-%n1Dms0#P!Uwy'-_?2@\d1m?w8PlY3#z^LTQC4GVaP+J]\u-Dd3HOF5WU`fmOT)&)!5rt	H4C@`I;_-kU%`(`+o3%\w~?m	lIGU-5MT,GmK(\/IS$8#j8
bk&QaGjN+>u54}*aUiKrVWBeC Ll=mqfvB)5inrRFQ;4"hE,\G8[BcX"i)0tsRhD'Ynn5NS2^ww:+IM7:}98
Q~)u7Re2"}n3Ik#*{/"?W+>i/'(>8p?MtW]o8Al65zjGl9Ng3:Y*W~g\^$)=c :VpClI{qHFUwz&9C:#RMPxc"Q[s 2v5zzt0K_-fxs@{Ycxe $?8_CA O7`)TsH2N$*su-wKX6I	6[AuJyL_naCN9}sLrK/BQ,pPb1"%kK7o4PGv}3dNl!K%(h=,+]|Ficief9]=WT	FC%xHNbT@qGQLBB'l!=UOw8{:`(	3NLjnB85UtPuM RMvNYNyY&y'=lzE\|/F? 2j+W8:_rcA8:QO/QqXSW66IaJV#IIxIi(BI9nImt1"%oOWv,*4(LP<h3e`AoEX{gNM\i?!~Ue.fS)|u2'	)%^N@*eZ\01ki"S\oz{`[Nrlj]_*t	-^OCH<eW Q=AAW1,3#B)p1=36lAY["ctbwr,g53v|urxYt&hI:tC~}x#g}Vw&B8Ikw}
N:&~\mYrgZ9(:|/x4d#)^+j)j@^c\.BZ/Y%8%bI	i=l.%x4{>0LRN' nq"ea9r*%7!wNk\VHz#_F<|G9/kV_v+2W7-C])*5;Q;_Ur)#)<#,x@Hm+8\uSfd|tsOfQ(8)5CK,Jau=7Ry!JJ5OA_&S:a0*|DqW)Tzl7!vwvT^K~N?s;a_M@al8k]Zjbc2|H`:`^O~jME/?ZV^P?&A>\e#O/1O=1?EE94&
c5;8Ly:s(\ZZC{{2=f~'XAIRP-'j,}5q&T"P<:MlZ@	rbu8?CJjtUxU(/+^V 4##|~wvK`0N>c0eG%0|K#1O.-K	tY3evm^O< 5bmf?;YV!([eG%)~(DPh!u}Z/s[_Nju9xh|4538I?fqUxG@{c[
t2cl](Q% 	/'MdY+F$ @ed9m;i	H@%^B89V]B9p%Cy+S6CFsg/aj$$PX3>ezd7E@|XuS^	3@dJ[q1Jn<)>9u<ng-.t<Xu$
[@JMuK
~ZmzSK.Lv7x4Tx[:jiy *VC+:yXCW~
 XT& sziYcD"_(X|HQbW7SNoQ:XQHOcWU,1AFH
Gs8@FJy]\0/R]hG):#PV4sv*<a9qU87MJ	Hf{Q?la-O:#)jqfyonkZb^^swm#bvsRjyfOeIsn(,<=<P<*1iYOY;Kxr1>X"G}nNZ&Cs$]]Cs7ZpCP+ynu|M;Ls:KOzD[# ""hQ{nU]x3g!9Uz5O<4Lmg*_kKCJd4mx;X_PE#	~u{xB)W<//n44HA:h1(js7{y])&.z`B)5zGOLo:_Lz'CtUN{>r]MR?qUhV]2HoVp{L5<RpqyCyE1r_|#qmx;T~m&}ww?<X7 "@&%9>z?6/* yKRB pU(QtR"ry)A-%7'k]Ve|_pz\B\J9%;K*24u0@ c`Cq`Y8_bnt16={^Djc;+b9!c9wk"o<68sku9OAKz=:L.BRSR4|{H4cA"/\@c8}&,&Hm,cfpU9l/G"qKdd 3ff>wvs<5=v)X{cP@895fab5NQ8KR/Jd]$]N,AX#s\{k4KnBpY!_As(=\8`YoFkC_E rq>X)*~]Ex;4V\`aC'43t9KY`ORbL2W;|A&WkzV=L!yq
Q-.D;By:>fPE"Pbh-&5QUH\%1UHSwLcs7	0/*.gDr*\,tw"SVg}Zo?#l( a6[q)W/lI|K=Rt7&Z)=O-0UQ_~yT'V`[|:l|}}gGWQ}BixPE!'<gpoJr}dSYJ"OGKAxt$55i6X:>b^t=dGBR8]{+.U>?DihokN`wUzf5)XkKcK0S&z>AO@o/_eI42k-zJ?cztXn.z7"|NTt0!,U	o #d]W7~@}:V@r{])["2"GRJgy0/N}GR:+8[O!qcg\1cwGsFh<fty++ljbdE21S[	NSs&j0GNb{}06nR$16N[WvZOIr:2m'9$m8mDbpN(C$9#Fi+KY;,=^SLKS\aOUsFg2~XH1z$o26Z#8r('t7_>a'S%=LOxY4vFx6rh*7bCJiSG`b#k95R0||b!jh6hS1b~ux XW~D:3z	E%z0p%U*L'<.-'Og0141,^hNS0TT=1{`#vtyT2b9D\W	r-gNF.+8:gCJ'msBPo'i]b|YzTi'VGlvqE	h~}~Ilpz}GRvVUidB0b.>Muby' "3t-6x!O8;,e+"1p}&dmHRdk]%Lci0"4\k*t/d:U|ss~* *(.OAay_BP0oVu1qyw@Qa-E`V-Q, #+0+#qK)Pqr
x>T?Un `j@!<ASd"w;,v)a[nnVoy)]@$fK3Ix2\\N@C
|Lx&"T=NXZ6-WFgs.CVYfeF	KW<U2]h_{DO}.nx<B2`{
PX.V_nXb?6Z&33`:E]LrE"m8O+)AW`]-4%*=ZU]t8m#Zc#=mqiZf!	2Y=JrS@CG'l]-&2[>xm5>s[YgFl/aDA@SO<HV_AqKGg-YE7cr=K7MkI(tAit1iBiSp_IRuhL]:c1WhKC&{'F+WTd_bs`N@'U0x0Q^AyD*MeOy+Xk0rvCK4AtS=..q[X&Sm0^Y&<zW
%h?VPF\!46Fo0}D|1lWk
Rj'9)P"vuThD]F=a^k<b0Xpeo6GK2LmQU,;!o#fSgi$AU0\EAVB+?vDyfG:EISG"jVd=25slEWz,v>L)e$o|z.2BYL
:tg.kgX'DG9Lg~_DQ:TNr<!;"RD[ubwwtJF.qc9:X(ujoV|1Wkezeh$XS
foj;,4nY	<S"GxcWoGEb|,b,)89C'9Iw)=?-Z`458H(xjoZ uo?xu~9x{.Lkbc".~,EUYRf]799z$i8}R!	gt~':w;kh3"NqJW'G.mUP{^(~'E_Al"Ul\FaT=S
Q"Z0e]#c$)=8KP|[9MRJL-vfZF$iT7iEJP1`8k`g1*Cz)e+	@w@9HX+ok}eaJ|u{@&LXO]FaYt?*DLjXPP'.{@#bL.r)+]==mXkz?#PkE&)m,p!B@QhrJdlQ<PcewY@X#]%-kwmmj!0)bJuDH,N#|GH)!=FOWSAJ9$@Em=
Z/Yc\z1!hx#;dvoyY64Y|?#8	]LFt(C S\
^D}isp7#M1Zm%S9^Z>i`MYm/<e/=hL%FOHFD?Eea3C=fh;J7p+^gP ^bg?D5oZV
R }t@UI3*9zk%pfiy\zhIbhpc}3),'X-]e;>%N}+$b/*[#"&DK)BB"Hn%I[<c#V|Bwz^U|0LkZiT%>]	rf40m))kP2{[]DR"g?M5PdIBMUb&BrY1PIs*+DR+nYZ/y`	o X?p1; 83+>obwv
zJ~OASZCv|-t4wo#NV8bV#V@nN??i0(^7kEA^oyG,3WD:5eafs(n[#$TS#c,'W'Jn!kyeSTBB>xlg;'hmXQ>'A27#y(YDeOE=<	l<AmA:z/vz_+^MF_%*km9pO$fc;[~`[fq-3!5v gd`h-W%YF/;]-=>!M6!9j7*%5hK[T.."sg
Cw[@tZIs65{ffq#0E7
}xdSc.it{Ss`<<$|dpK`oOi:#F\vMse+^?nu)`,!]G.Fbh	DQB	M1zfmD!%Db[LYMswP#kAf5']3Lym|x+Tp`8}=rc)w,c"X"kPm04/z:UCvlc<+{V4_qf1>aZ[cgMmc0(-!t-"vS?Km`OHLd%.,	KR)v42x_
@jn,<-tIkNuR'R@Es2/m:}O+J8?a>.#6"l9'`Ag1uR{WS9v&Pr{;N	rpX`:us#^\19q0|8\;s7Fa39r ?NaNE,E!6gaeiiD;B-yA0.qv
7W][Jlf7}+
$]?_+r5!s'dI:|ngT,2s`0.U<R;AZ<[\,F[R$Zc[_Q/#niY337<';>M399&:KhgCuJ'xN4"}%Uw9K5RhG<fKu
i QXzf{sTC8'Yz~@<FsY9Of-S&
L`#1snO\hrTZ?m#H5?^d!/g7mO,^#5l%)c8u?Su	*1z]Za)ia?99pxd!b>x?H@~ky%3\7CFf!|EjY&B4=.K&I\1b)JlF{PR0S/xI_jJ7hatCi|NExC\*3=yn
8"TMmhw5/7)>JyqZPcZHP7ZWslX^|Sbm5ACjT]koE0Fn^)lt}de!NI)&&\JJT ]{qDOy6oSL.S]SOQEcBJg=g
 c DWqws)j~Rspf<U1W?Dbwtfw'^-k;PwXsrO_k@yT+EaR!;NWCz43C(#bQ-WKo!+Owv[\px+Vr|g7r[7OQwW;E\T"2M9f9X<Z	V6cv0`.qkd3`8:CW,C	[nn&92i(0`=9c}x@Q'(y>TRVRI3HG'ZS(bmQym6,iV'2V/~M5m<Yrr7J'Iq"\KV>?<}YU*}2a<XxsmJIj:;dHm*+kLG@\%p=wt{['IkiE0b
?PY`h^$Q609$f43qEA[Tc)AVi]aN=~_ObvMdk*^ n:eY	v.W$Yr<!>{l@H$b*/`6{DX.ff&BJ1Vw|'P
YC`<^43u&oZ!W*`STh<Gn4jiVak-(^$o"o9't5Tcu`o6HWU\t+["qq~yTu<jimc*ZYW"V&ckn:
U0b\vZu]`e:oG9?]7	04b$zV.vnfL$]6
M+xGoSp	u0%@q,jyL4W?6d9&/H},AtU2S=jcflP(7r0w)_Z,|bo7UIK/^A2K!9aE6~j[akT<(HL|N'R}LZ>q>WmA>xHc@6qS8&+.r9?S|Oq	Gl}'fL=UYF/vJ^4)C;6|lH8> &Ftp #NpUWv
34&zj<RSG'mZ!tIIOiz*pSKV)Jim_T{U+M^zi(UJ$5mx&eufd%|Ev\TbL~W,~&oHTtHIdVVMGYU>tKOUUCtJmLc}4Ki^02K9'6!?aT[CdHE/X2s>j=dY.sJ6yF/&%O6G1iTG[yokyznN}p,?GYZ?E6aRbbdfvZ:gk!`0`25P-Y_)QecX3*I.Ch),Xn	.I4*BodZ>-02=0a~2[sC>zlgU\lkX6#J5?sPulls=K6=i)4OUmzjJ@B>MbV_`WXyQChvam@&;uA))iYKmkdyHecW^r_j5LI:`[|@}3]ejoT&K*-*[r)<"@s4($%3c!qIu8 nk=:l2'*Ht27)[c,n_STMANqobSgmuA);Ke~h?|\l&v~p[yOXe?]]Fy	M3S%6`Da[s?CiT`re"JbI!hDUd3{f/n,$B,ET""9m3E|O{~8()k-k%!.s`\Uy:Y=;	4 [zaGS'sdI7Fe$J$JRgzO3v@w;|[s$^*)+C
uK;+6G9m.xg:)JR
NoI09)if[1$s@kH.'>\P-v'zKt3s
2i^^5=o!+OU.$'!;PPFit}PYi,Umi-I`	6+}NHN5Q`
jAu%Fu3q3	!G+S}i1.F~Jw9iQtb]i	%C(9#u-ZIyjI0GC9thkOWw-`"5OmZ~esS=U7nMa[qX8*>dB1	0=c!!le~G4Xr8#6cf8Bv1Z-Ybqw]'
00PF#x?]|&Dv*'n*.D[R&se[I:7+k'qW*SsfS=2bD%;R_t_N]D[YR'^vX26lP`'	Q5Y1])s{~gc0~"Cq^68}"):x;5PmL}ArC(gEUIGJvp7zpj),P(4-_(z'"8aHWSa~o9HQwUT$|Qo(N11HdS!3u2aza}-jmZ/p8a<:fZ=^{$0HsH7Z[gtzkR`'m[>3K<)iO1Z+kTZRh*AJJ$#E$.K08+4U$@0>rv
C!6K[>6/9g(7%5LQyx{-<rdH0hT_1y':]	@?,8j4\)s6u"B1P?9}Ko<*jAyn&pwH|H^|9	D0ajx%R>+1|6W`QN?jl0oQ(1G9K/0d,EB2e+>e\`#zH7$X]=C9dDhq83j*M@w>03sRy`z]%JEHK:?[3ToGLZ]_5ZmAago[*C]S{~PF&hj\J	8 Mj%	g'.D1zg4+_axgVlkJPoovXDwy,T;Nc6tb"ys2 36QM!kJ2E@]rdJ}6Z1'YV>"D5PRS3#=.!Cc)/Fy-/c5-s3H:i+3-Y.Ff2"tnY3dK`-<L?|Uh!)d"AI)bx4~4i=[MWW3J+9<Z&&n@ic={xTbe+\%]gr9:d,oG0@ccO>"E@YND=^>FV*.Mi`{duX,f1S
orv^T3_!EZ	nKG@yrc_ :0jgK_2ZrPxd9-uz"0_cmVM<9}iT/B:XmCL1!^B3xO$7N'DBTLW#co
aQiwzZ9/V'@/.fv*f{j0e#-;\`\Op&j WC+lqDmC:tih/:Q5*|G!:cEX
P8Snd;d0V
'00!oo7yyKk8^gg)8tv1Wb|_|Am]Rbgm!GCi,syJI6v>jh;1|VP?jH{F4dk-DbMF/DHbn+#FoNE#E/eRo14H#3u'3? !ala2"_@GuEyWPh-0\g&|c6O)*tZ$wk-414q+DrFbtE+4f,B>,+`^mg`Eol/U!91;Vso'RAlGk^wFA9/&")'1uWSoWhRg:K,?J~SpdOjzC]RI5lhQP(*Lw9*Z/geykuyv8z.%E?)s|j(E,yJL,;Cu%Hv9Fb0i)[=IK8B;?MOk*m\rs3Gq*)1Zn~gz9$=B
=y!Ool=a%	yxXE(@L%1[#td#ew^CN`Z}Z9Hw2m5'DPBr_9U&D%+_<@RZ5j0+A{)mWUizNO0_^E+.J+2mY`U{JQWWU.(oE5^<pjwgQMGsAwO:}GA&Ep(faiRqM/Br%GTWdPJP(8'b.4eQJ]^rKr)m8_?OFxr'V!>P9qM?NPYUUDYE	52;[S`{G+(pDDQm0rIGCi):M;[_*QCsO(>\u}{s@udZfrt@EpQr|A}rA]retM;":\L2D}nD"2=l&"73/+2`I5~j|H?z(=zPHjRdMl`-TVL,y!ljF-gcZE}V>qFE]1.J0vk	_F]2E.:q(eH5Q2\@:P(yq
dec\>2-UW&1J;4yN[&ZTowrkzoD9CqG*WqYf8;?	HS}AI
7
uZx)5|,_&QTsStDdJ\>+32=LL"9BG5ZDUA9nC'2d,e6
+]!_.vttOkB,zzvR20R*/K0V^)4f2o:,w#'zjE$-.}E)QNb	1/G~97W?]^\b4*F62?DE
B2^T];Q<s-H1Ly^o>eSBNE}'B\e7+Y-#ER*XMQimsGe/9#gGEDu3pO,52n4qzm[5J@:I%{	b	Du;oZ(E@jsf~=
}RiOS98
?	~3Gl|{fgbQA?{MXKszXU}!DQlPk7}+e|km6srJ}SiO\|8%i~6tG$
-Q?sQ[/W6&+8P_t q}]o:/9B%P?=R%dfq/N_tKyq:gy'gpKhV '|HlcTU)O2FH.l.A/ 9IHpP|\n5XDILXny,J8p_R,^H=?VSBT%@Ei%75'
\*hSg70*rfG{3}]^j@W{wS<U=vbHmzP2o17{] 8Jo)NBvl*IH|5V-.{eC_
^L2Q16>G"V^q80zG)GOSz?L;u'DAE/ s8R\C@_D;'MKGp.I'Zmlw/MC'GcO=_EYD*XaA<y?Mki(z}C%hB[V!I1r?,3u.D7}z{H0zk
?@&AY\Nj=*EES=@i"4qUkL
N/Do_[,i!<g3GQGG-TN4t;TV+n;b^P6
rVkp!)$GfAD:]xBSySIBBn0x45K1(;#*'N5thr	@WAk;H~|Un{9N!	AanV&>X0HoL[`F:,p2~\;	hfQSuWP'L#1WmcX1Y[ZFqWC9G%'25/S*>3GcF-J>!GvnaE>zb|i3I,+(,)@C:.z.scsT=(XKZNaDA	KO6r
+bZ<ev]b\#t)Fs<{gj@q)em**wODYwWj(*|p4y%NjF}CM.E;Mf2hPXXB|IHzbA&|?opQT$^c2T!e?kUY-_#=	g]`x#$qE1um}"\mHxrd_l{N1<cp1.mH.F?)CeC8<u>wowU?}Hj,f"`Wx. y"PjtYiMjX?\3qrK
Hx2Jcj0y"G1y~8@.7P5a9-\PcmDfC)e ak" sdaAN;-*)xUFmd#f!(qQ]9vyKd9{iFXs:;
'g/Zm:S`z$@4"9~l6z_q78OGqg9<Udy)LA4L@FpW1	7\?-w?-;F?<$[m#6zB;uyC`WE21abA	8pk"R&($a$Kz]I38qalbEzenmyV@g
a+{+7B7uwLE%Of Sws8
q+NoXc	Xzx]jy<qZ+Z
wv$caC<=LN9Q'Yf3asEVQ&e~=?zn<Y\}R^r\P!%%kfW"8N:+0K'-':U4al+HhP2 ;67EhKwD!i;6Qw`L[Z1 8Fw^DFxqo
/Ij~<R{F6<WmTyZJ6]D[rYV%ao1lqo+UPc-|QY!eOL(a}d]wu/*{HPy=U2t6npa^RNNyA@WNP{fW[m~}KkNcZ!gPb[8\RD	0]!GYcx%))<y!#3?R6_a*/jd-"kQ6"kp,h{vf-dk76R7c?]7War6tjz`j5*"]y45ib`LT`]~NE.of>]^C>
c33,Lk<e35,B"5v.h2jm[cO|^=DY #X"]ye<"CP!D4/-'IMWJ^zctX{~su`0H(>*uGc<hd8'99:]K]#-]P<i6'070Cxlo6k=4F{(gsbYqE.3l,vXZ9*a(jZbWO7M@5r?}I|gd#YZQ
t"35f7`tci}%uT@dh"WhNqv1#)Q^7$huSt8#F;1<[8;d-,49:W  $r@wnN;`/]?hw(6r4Nq1Nnu-y90,-rO'c7)=CVg68@6.]PZB;4(y@yI"5%tWZ-cGPZxJ8_n:uY"[e	_7)J>},=Yq^EIaAS9x^u~v'a)P.jm
mF1lt5]Dd`<k9H;txkC'g>[GgCr1D;^d.|_OJDrE:$s^	z3jbT=_<V#~ZBvpsA1,>)qVhmJ@1RQoJx;NnJ?9:Mna|5N&tlDy!B.8WB)1x`iOp8p%}DI=g]OIy:(v4a~ s[VtGPwhTOx{wfjMw3GGjOK0Td-/.PBu})}d[g!ZPA'w@"
bazRyH66L^j.A]R:f!_DL=@BCVF0]^;Qmp_*EPx<ZYj_*+Y%zE"mp`+l!4 .+}bN0sSZ>tMlFX Ga>Yq@^1-`:8H@Q)oS	RZpfl0c4#mQYuCYU@y1- eF~IYso[:AKK&&R5RWD)2OAYRuip`\?0+IGV`@J)>I;
uP*EchfVs'%O]Q0CO8jhj;T6X>u9;-gvhsqNg9u#_L{EG?	'J2/&(1[ CgheT`T/DVrv	.$@MG9Y!5:g^J]??JA~F+(\1)=bK7a-Lf.Zhjz==dDF1wgF&PTOsK-#qHJ%sqf_2w	\'$NM.*&NLdPSl#S#~gD`5QqrL`aY}VCZDUv^xgyvY#np]BvN^&I"#0,"c`knoLqA<>Py?.VL#&Y4{I#V+YyCWZUo	xcEE<E^	:mJtq:rs@	"KbPi4Y$d<# 0dL0&~%Y2f7h)kD7}#*2z7nG<J,^.hHnz}+&"?Cho+$/w":0/^	>]G=~b[*!8UsZ,	"^1NuWwJE^YSQYA@G|t";
Pl)J~O7B4\\v!3*|gLhtjtb{7Uxhv`}]{mZ'&@OpKAxa"g+ixO?qC3{M_rv9%Je}!VE;a?zBBzrU. :/J`Sx[o{Fh&r2Z}/5wM'Sx5 u6VpZ	M0!&>OFI2QNCR rxDH>[vE_nW;{,|lN|1!w]X]wW$z3:?^Ut
w8|lg.&2f,='x!oCU7$oI!=-{}PQqEjk= qu}7 MTl%EaFxM;_/G\IJTlk&%,jCE{~:i_~M"e\n.*wHWvb~5M7!"K}. b<=A.D"/<U	^0s8|DnRd!l>n1!1_:W2)7kqqka(uTF'o4-z a^q:un.|>O1s,"CtjJXh;;&0R GE!*;?@A:A4`GT{Fw^ 9#1B^)E8*O]gJtCv!0>a"5xR[<i-"g5L
iti3-P0Uw 
JqzUHcQ+y;`PqwGrisgge en/LvLb;v(7!_jo8\}R%'RV?)7E~)$hAay}JS$hTgR9Gh_az/0*"gLD$4]=oAHc@s5AH%(^&YB'2RpTjz,Q\%)>(2T%	w;+F71<q0gG^Pi~5HsyI"4?svm<lb`_[1)QvzKoetdWCp1)5[^7t*N9(b8q	Kgb*":$oL-LQV9'r%pxJIcn>$h
'a1bP>He7{E& Am7F>l6e3$!DE*)b+xo!+G5gw$^4Wt<7YI(?Yceyt74,@gVb{k#nF{sxb&{,6zqORnEd`Yb5]MR;HZB<Ec[jVT^E\A8SyYx$nPe,;5LjCkj2~w'BbCN'/ dFDl'Iq_0/"'2vrFI-|X(1`C_+}C\wMPjgX_7uZ[72\Th5g\@QQ/j"d*YYuj)QyguG	Z+^p#?veiyI7 V^w@qg.fCq(DK$VroX3TK.%Cv/:4z)|Xv46xZ.bz O\3nqZvvW&oBZv/{=Vev*`6(_Obi1Vmr{-uyo+>G+]p5Ao@lu\\Zp7s<G":64vSnC5q'>R%bxdtHl(FXOosxIq^VZ4{5QJ{G"ZEzfp(7S;E*<77-C9
Z"gb`b5b!w
p5UtChm5W4R/yQW ixuk>\9"5Kl/@_zp6>9V8jH1,Lv~u%h"_Q$.i^eV>!/Fjrj;w[h+K1@6ml7Mto@hoYQ4lYR@,Es*;h 7@-b#G #,U&V,"OqG'p|PD
V&_DA-J6}r=Q,}'EV=:}qS2i}f39TI-`1,yq)IK$h*O9o+9v%Nb=?,<PNI!JwZ'Jqt3pukHb|5uX.j\rE.ET";H6~%@V?}`Rc4 )VU7aDa,uY,66I^K^T9Kwb=b!ZuZoEq's@+/"^ZYb{a%$1$=eJ?!6,28=EyG?KhXGMsT ? jZ|03UF/\?Guvpj=\Y}[Y /^:%lQIsu{G1]LCBbGozxE)ue!vQp{v{bE=mjM-du.9!{u\-xi}U:N$]BJ']&EK'>C:_x""Ug3EOC&nAb\k<WUDhCk$8&X*+o1bN=5}o@&KCJ1u+CDe<'la>grX6,B<tf'e7m"Cl|v
w`Y~-]G\.Zp\%,o]6;.nOC$fpaz)lE)wr0	n"-|(]OndYN;}74VWptLew0y}-O.n~_uBM8'GtCt\sY)&#DFhbs^od\<141\9'f*Qvh74(~ahm-
MZFz+ItnIeTAT{^-to15vym $t!pTg)xh&<.Cd9FG&1_(Br7|vu\dk%JdM[X$P)4`f<.1)o%Sd+Z;Rq:bggh/LUr8+73	2(5H[jq+dV3`ep~\s%_=k.h$qx|
+.~K-$"BIHdYvGr
YHG@9{"9K2Fp-"s 6ZPC4fxrMtlMfY{>*`|B60H9H`1ouUA|bM+iz(Ve1%
Zo0P$f.jnV=	iOv?kbN)[5|m|M^"V/}nKC8cxjUpQMs0\@vKb;h6["t|g#k|Z<oaya*iumM?)z
Bnx;^K6Kuq.sC?,KQcRtvLERWDQJ-dw@D&Dl.0j_cdtd1c(Wr9Kv=J.|:%1pi>e=u4;Tse#yI0(m":@ 0j@y,I4$3iN+Ap:3}Ac-(=4Vz aU*]bnFaM[dpKF;)Kxvm=IyUI<!lL-UX+#OJnQ#X\ix"tG%>QK#N[RJ1!5qU4u46$Jz)z)X8ZQo%<1[8hP'@RN)R5%>qdvt0-n));F,$KojwN]P+;in,H]'Ewa\6H#qdWJ:II[<g:3`A#T@3Lhf/:dA1DwNJk|3Aw4/p-B[0CdMB*sTB2YTp"BJG.r,KtjQ@HY-u!~LK37hQM.m5s`>lwbC}v@nD7?V6"x`tf?%53Kw9/J.`vB.JUM$7hx3cjm~ynDCDBuU>tbhf5]qz3QsGaEqQ'[qZ2lk-O/)b[3LJooyPsduLG8,W$qu^\+X1U`b'uktGamCIOV`t+7KAy{KuXMlg6"nJr ^&:@!]%
^d4I@x6"IsN,,_k
xqA]%5&"?_Q)S~?#f0RYjs$1! lHHUqr7zhhs1aD>Rm8nR)U^3gdf/pFsgAA#xm>1lq<-7ekG16}pZzX.3Gvj4JYX]9Jx3]jr+v={1J@p+3_ 5l|i4%S5m+C"J8E~/%y|3%^ODg1R^C>~DF{VX\~'}u\@){_x_I$1*j'nT@&\i:2VN)J?e8PRUcV:`&,[v;C<>.E/,g9~'bznCXZg@Rf0cHt%O%.H=z?YNBR`fCG\[q%Te&5dGbwu/R)MDhLNBzkK"?V8E}GAiPG9A`&''8g:DFP |t,^;2xIeB5|P"g3XH'aMZ/x+yRwk9*rRp),J+7w<bY)=Ifmq0k]w3F
	6B#[s~$!/SoTt}M-|j6srpNh< .coZ	5hiFns@7ehJI6? F,cO/c$*vnsF"l\B|	&%Pxe?%WJG~
YgkXA[uLYVmgENpEvYg"
D'*tSvH6LcvSKw+k;V$Vy?\8:V\
xoK$GbVUkK2"\&Q<Th`;P7BpeUvr6<_%,?uCZ;hyO4_<r;n9vkHc|4'_cag{Ju=}fJA4OFM@H+IZ!a&7VdF7? c02W(:x>	]LBS	&N5m7Fk9JO
QlC2a.x
LNHM&=OsT^w4d0|z.2Y9s\.*<
}~dzh<P3z`]AEu:in29ROQ;K&$![<wb	YIdn=iqK%&3ETYtYb9]/h'T,ZA^G{O#x:w7.,=y*9=hx"l,F7{!Cc.B\]M{kEGz#a}%<<O]z;zZv2_&I[VsO#LZ!AaK	78=)
8qKnU<rhgBY4$+lf	v)%\-{T"jy!E%?X]{5sT4`mQr_ce^+Jf;/?H]ex	yqHa*{"_%,.fABJ[u*\|jRsfl]<<(eB
nc?5	 hIEOhiv)L>N;WCKL:Bb~$xK&u)D(=f038/a@l:):-yX~H(s\m`^c][4WM
A&gjh:fj64Y`jhv}KD}Yw.BL=:K0.k1LM,RH[KRv1_Lv
2u%84C"]Y'PjeAGz5U<iY#%	a4US$NBnW{M&-/3J_y3YM|/WA,=Yjw'V|20y&i)>Y<X`.Tl[i,2Kh
iP>bzM cN%P4(.@sG,{$~3e,3()a,t^L/?2>XU:'Ry>\('$5Stnn^S"Q(D3k<V+9z_JXak:DS	lU	($V_1=,L',P3G{)U9#e>x$J>z2Wbg\./A	+o`"yIk	-E|;oht1#/LdX>vgw0Gvh H[#Q$MI"
^GJj^{p:c9@Q(V;|WCr*4Ihod2n(W*6NzTH/Ug+yk+/*SO>j!Z?[]kf_6#|=2h>d_tMmdEO)jv?}XiRq|PtG#G5jYgJV<
n5@O|eaC*%n&5c+BI1
-I~H5RC9NcZ*c0AL3/kyoW(/tPwGB;sz4 J6]48QZ%n+haW
s \V/L
<v%vUp5do-+7j,Hoz'Xl?EpPZaf/6~,\xUY63f )H"R#r=z)hh0z''IMpaov)}_w
Z1`+Fupk@ ld,HY:!ptgw`[JGlO|Dy|,mYyZ	M.*aHQ472Nkypic6kz4PpJ>[5/=#h9B_9Lzqdokw3Gh5l7"!#iwk>71/<ih{'l9K:O^51T'3~ddD%nj/?}@^2!*L5?0Ra|/PgCtDSII!!zKb4b	Td9&8^T;SmH9P~>47B^)M;IyC|1&&,V/W;+k2'My[McRK^1-d&?0GacLK6__n$i``Skr5.c,E~f?62;1!kA~^fic,Yq]DaoL
44v5cAG%O.9!2LA'[r0TjtB.![#$@0ZEQU2
T'e3rnSzw&c`9z;Q+yB3\"1IEY;)#TR=Wj.`2}5yg&pJ	}zj-vcRi!N
S(h	~/rf3ZSMsXB}&(]+.Vt;Q;XcjP\:Y
JCXp{MoLL[q Jnp0%+U4v
O7B(8m#0Y[P}|@sS( )I. vvLxrK0	DaQ\NyES}9MFlzcK^YnzxDqw{|(|n]0_)/Kf<3=-?={ebzdl
+@}}e"P|u-S{W$+G;,OAFX4f8 s%n:=eEtYKqwK)q0Qj>/GF6Yg7"	~!6~/;&)Ng3{eDV1L"Y8k7WQxih~rmNv	788\e]S#$4:[k8x1Xv2r&Ch2#@
QHH?tvZl$Uy*HZRh`G5#nYy%kn0c34Dvn",n5
 kKR8IzQ4IWw4,JD{7U@ix47uywxKDy6TgzHXg`ksUmR#-`:}[JJNP.v"d%DgBL6NQ?s(oKv,4`TtZe&f0 @:cVhWFP}&/+s|,MZH([yV2(EF;AW+nW5F@a"[-CY##cVCMd<FD.W^!xKA;{y@5*f>tl:zQ$?gCd Kc?T36n'Pkht%VzGo}Mu
%S*	v7)*k Lj/	bn,'p1#)}YgYCf>Ir1
xhg;-Lh-zOG{mUJkR(xGo0%*X>wJGLx?r{/mCy|CG8>_A[hwTa#rjH/{[e/0?%r.#z89zv.|aT5wi-_V ('!f)
lK8\s"|kVc,va@pHaE\(?kPM-I73ksD1?e1N3}o5-;fr]zFK=IA:- -K4/-6S'(`sJzL!uyY36DzY,p,}gu3RN.pE:/;|;k$_Rh X6,+\AB-6TsHi\j@;MV
f<9/HJ
zm
\a#5WZJ7H1v,I_%|/)4I+g- \FfPZo]h6K1{~/*y/i_C_|-n$B5(oAPOD:^yZ>g!\u(-CZ%]Ag9I\[L8>g#_~GNA4J3f0S\7@Nk
}lD5fok@EOuW.q.l
(o./
Ox9s:Cu\(=~	Z(Ev[+fgbbC 7zAi],NJ'eg_^M
iiWhNY#Ll)AQ[M:&:Z@[@xh?J=[8dV/F?oWNR"H`lI\)XQR9xvPQ{>SL(@Ap]x?&vcm79ca#V}GI("h!C!svMmYjsJUHz}{4}#q@T#fXZXB`N$(4Jq:aDe.7y_~P&VF<L}8%+;Y/PGCq+IU@,B;#a4}St(-%HHqe'0}4K!+i:Ohx9Iu?@kZ!x~I
gkVLG&Nf6Id`UHRlrE5szA.`bZKI0L|K-Snull`fy<m1w>%dqvj3WDNJifw]y99>ukO`UG|m*%1sw@YYwlh.zUlP<BTJ_v?b-G"ie`gkIt>F,99B/u<wj7A7@_:_jBjo-=P"z)G8O?'SL'YK+l\GjxgX9(8<`}gp3aNp-q~,0lR
cKnO+bfVzF_ ?,>7fp|)d^3P=5YyC1n>[7@)K1l<_<-#EZqL"v4m=FIh.od!j+D81rqsCu!bCc3u8o=YiOjI:eQ*LR1d}H!Q_6<X.dA0U2eK`U(ptVp4zO\X]*z8.rX/lKYFo0`%9kTsc%5OWv/"4@'x(d1S=`cK?1>{4Lu`D()eBE=0G^)I\vYYmeX]l`c_C0g*m.eZQuJbO},85C:YgKp5WC&+DnQ jIO?Lb87YiCsf_VEnS`XH6+sp.Kv=9hK0NJ"3UE18Ym}4_dKy2t2e8'8](wEwSE&cP&tW6c	iE_E	v5?cN2MLA".Y_pi<=4^-blL XT_U5wi\T*g[NY@i&qi[!Qb:T5iF_q%`Wm5aXSZR<h04U"W#T0iDxZz%8)v"pEklci2U8?irer7JHzsI`,c+ Az,s{Ztq6m4ZfW#<xBy~L)-H/im'M"wJwFGXV<4CjB9i(pT#GZclq
7|VR';kEL7%&>82``r[gSXvcn>p!f7Fl"q7V7&("r`dmC#	T&	RmO	|O*#Z'!+{y$/9g
x),/5p,*1L:%>;8`pSpwKP=vus`,(Z.>]D9E{g<4:g;<{tSAf+ e_ABHt{)b([`NF:HNt4@<F4&k5f'<I=0|+?<w+W<wUM_8`..s$YDyUZKW;ja40t`I-CbM=Xs9 qhv|d*Y$3if'+&Nz<hB@A{uK24a}\z@1?%[]U>5Q?_y^}eA1l1'=Vn`C}{@VFr [=*3}U;.v{G&uC3W-S{A!OS>f6Anw@v>7@zq.8;qs/YgB.TZqwyy^`2H/d}:vC;
!h^%0'[=V+$MFSf-9@AN50@J3s+Xo]p=NRuD#BT1Lkg#,{No.'sJ2QGR>y0JWF]D;+2?P];Y@	Zh{TD)l;dI}m>rS:fV7E#G3 }Om}fBIYD`{;VYDp=:.YUm2fb(A#c7Jq)f]molM[PzpY$,{)>f*5@m W(r)8@!s!"7=,<+$10\"is%7@!76oSd4~'y L/W:kcK0!*?w8P);%Z??gZd;1ZOsPhefCL2P8\b~k3~(RJ7p	2~hXD&y>PE]+>yDaCkttwz]pX.{TbZLtY1*)Z!s15!:R=>:'Sle"b7ef;J&^DwCk@ >7+yz)dM/F\ABm03Vm1Gh%g[HBBw,5weJT
j<{7qEn${"Hhc+=Pl!#vwT@$OkfYC_f0E>av4H_~yKfB9XM`$p32 ~0`Z7V_h#TuU|uU<{6_j%'OU-*:pTG=0gA;3i*0i?vW$j@(P#iq%xvw7@t^cdKa>(fh+^p/_l<V">9G)a7n{^t!km42tXw/Kn(vi2sN"1${}DyWX5~NnAp2PR1AHsv JLgN&feI|n"F8U|j{Y~LtB;c1QRbf,.)HMd.I/p|w[h9PV3fG]k#'t;io^x8!%;53vrsWw6
~^\dnsyh|<Ec\"U|!ScA.`sqD7;MBU35}jr(;_Bq`B-Ws+Z3j}6`\}9{M<xJw!i)qxAQ??r6'M@/<XN+~*w}zEJ%XQR6':-U$RiP2BQov5[}TNHSB=B
D@O*4|+KD+*4"DO!7ME,$q!'&s>|=1~T%}Lo<(A\$x(dz.;q35AE4!X;*t $ 9s#<`75gCUq0e~9X;0r#YVx<,Gys#a-8TH#La^'R7e&bE*2O
J\/ lso\N^fVR <.IyRsO&t4g.V%CP{5p-!aV-GJgX<"W42Y;#S@_evw."gu^^(b%NCy^4T,0'oter_923Zie*[%/c<:4pxU@+)]_XevA|0QI>me}!>^@ae
],P42"kE/q@:02>[*bslrt^ded
O7[SZ=%vhU5N&hJJhZOFY}VaBx0\OtQ6V+ZqN}lSi&"SkusQ,Sldk4?yB8jLH^$f	<L7n`E|*<thw/=hZ{OJ_qg$k
yaP1SSk`x{'W\hq3 QP&R wXIkSXU	h"9j$cDAR	{,K,7?7@>.AzLW@I9k]zfO`{xL$|(y\}@0a#@OA}z [&Lf%oiPb~83ZqKb )q\)@`^B#v1~+#9Ue[#XUzP[Y	pQ(/;!A-V9I#6N{{w3-6H/+"T#2D-qvdn48gy@?CV?<F
GHCE<[:k|'VSpt+p3ef`
':	"t;hkKS;-euuRFEB]j8W%+9vcP
D3x?e-OB8VJVyP1ZJ }r:ee/dv`\.M!:'[/NJ	haDq2`c	:nJ+@T>zb:`_zh0_J	4Mv}>8zU}pn	>;rP749o;pRIp>mB2:cNMJP^
AP\&_]=3tQSLRhiTHy)Ks##5#|Vp;0)Y#{Eig!N@.z?Wf=N(O}4u:cMdfUdj=3	Yllb8Ebt*ez*s"qUw=6L,TPQRNqWt0X[|Ik@98M*:OzDA:Sa"Ud$&?+W`/D&{!)H2*&Qer{Dq=@PHdR58oUN\0O= q`~w)Jfv_udbO*4\bHLXV>gW"kyi{M]nMUVi7QgQYHE7Ev%)=[ICM7|S!=gsVD8|#[98^8:i< ,j0+!7F/S!tx|"EBDN[BLB&<:.Sn=WJtr$0vd/paJ3*t<JhbF\	'2.NAx
	Gc\y|NMs/2Hm_fJU*2	W,4{Snb.X}XqP$>7eD;BtNP\N{]@K.c97#	CAVQo08uQ"NpA*+=~OO5"rEe:Lks?jL)C|"N"4 
e$F+*:K2&V4'<<na@g[&4{O@p'8x{}HkrMDczt2eDUL%_Xp{*w%Ra}?Mswm)]
Cs||"F$-`c#Sj,pRkhyl7,C&d=K>XRSl5eQ@EY4k>D7hJ5?bi%KM:9rL@m;T_Zx%f>9L#bI4;O9Zo5R`vf)BO9	/7u1bGn",(}x%}wgdTrNiwm9^h(M$cXFUNls<nm<Te;$/3R`.F<>WlGRiXMAo}Ne@ddN:q%t=!_9quGeQ<(I{RU>=r{76^fNHb(4#bsG?3;_9`sJFH.pC$%j
,Q>%	B9zw0Eu*D-T)F<QcS;BMN`.o[LKMW{ 9+~=c/XE5@	>E|I5C>?g}=*;?vt#_0)g^{QYkQM3HmLSH[37Y^q$PYj$6od	4o^dk-l ZbdVs\ScL8c]iHGFFHjP4=z%M:@rqfI9MC]!l{<mt3N4XGB
_Rjvrp2+kr#g99%e'yMJ=1ShS?f<cbvb M#N}awlQt,h[F y"P~6|CB`G_U)Y,%9<@G2Vt
9;0su3{;L}VEOZRu#3V>"<m:)ogmB7:nxm8z<3,fv)3+,vR#A2tyezj[CX=8lR?M6x^Xqcn0%,W{x$}J:H]'"dHS8C[I+>5cI*[:EI@mrv	#<.T-%9e&\He&>B2!K:)l9#t0I&hj`ixLBd?SF})m7F|LI6f4ra<!s}[?l><W!_y.wB:z?J*ii$,cn?n0JBPxHMfK?>]x-*-9sIC^>K5H_:&H0rH'@;WJc02@a7AuagtPt"Tq|(yY[CmBc1ZOqI6],h,x/`$P
s5a\W"d3BR7e3}>N+d3[$hkfm?U@[TL)q#h(0/mjA4f_12:*&yx$amW}^ 8Ud,P]C^,]ph.sB>ey#zFQ~g;xIbtR;m&^1#{%zb$@qOcr[8<Z>0!?z@+@0Q!q|kAvnA"\O8 /)~SVkaB6bSj#xE<t2F\V-1CF;5u_UX+Nh2*cdXc6lDdY0G>OiEe#<vel#U`A;ysvM6IEe!9:KEyM	Db?t~?e-{$P@UUeJ4l3&,G^D5yY>ucF{T/xWBf97&Z!EpRd%+ec7nNFTI9U4PX4Dtwu)VnXER~>Cvi($9K OcZ{?lu'jEZG@ThH*4ukxS-]~8wEu::8pO.v?ffdwMMt5G5LuF	{9a`Bbz"86B[TD;DpQ+6m>+),R,c*w51& >2AUMIMsk5thEAk^//}.UUE	
Dz4v55r; \\D:
h6!LML5[<`*Ph
GB%EP[I7BP	mPY@ZcR*JbBfAJh?<TluODcaLV1<|$Bfa(~ s9.\SQ[8PC(,maO"4aVj{B9QA(@w[p:sFQ%oy5i1gv_gfiH%5hmsEIQcTuHcpX4*9jCc5-o] QX`Yh#Co'THjdE8< <w}_?*H	h[D[O*lEsAq*aJW au#*OtgY_*)fAz#2Ugm"}oexdW92#.bf{"="NR]938_1/  OlHpJ"FD`1`rCoQ:"`mD8p!GSU?+:I(l^oY+FU 5$+jyE`a=PY\DDUq/#ncfj|0^dcNN;h6t>Lyop6zh;$dTBPf~Vc:0
G`k1Y)%mF$?$<C&lrjz>Bm#k
k|\$aGmIfmf?4"y\C02qnc,3e,LL"HT,hD$Cu=P]]-$+&y
S$NB)O*{b. F
>Vh;i/Y/v8H
JX`Df9H+Ni78&/eS\F//0O:AyDQ2;p[)?O06Va4*?^
C&,CAr"0kw!-nI/san`IwFwgPb JS3~Z^|3nG2Q=BG&lXG"cw&RNT?Oh 95`{yq;<( BoNip.]fFqNC0<zC$VIr`0'mT+s@I_Js3rg;%5sMu1C 1S9d}#z|ERUgx>l*.8>jGkZ-"ws<wqXB,.4i\R(d[{Mrfu1Mm1G8X9G<2
X^^Q09$.B_G<sx*
B%b-W1Z
wZy/S5I`lm{w0`)|}fdL
k,g,7vXy62FbU^	2<k1hpX|z1rQqg%/7kQ#3Go-baViHuCYmP*+G*2PdZqdt03OyqV39k^wr+~DAn698TU\&?AB`_AZ8G9w7	ZzLg{[[R@DOi7& )e%otk3oBTGG]Yd5f/NU@pML%rxGRLc^5Xw&(jh0d1#?3"Nm,M)huB*c^rr{+IuVTEqt
sgNup<g|+xAZ*.m8*MJyA][cL3RUdoH(xoz^	EV}t3hk^;r7%kr|4B8+}<!*GHJb]mUZs8/@\5RCl!,kxMw#k9/qtWjsd'aZmYgA;Ru@y)]R$r:Rl}9,A\`tcDP{Z=	=gv"r0h%jziG:Z{''^RCE{MSC-u3Nf0W/O(#+xJ=EVEIL5`\Y79QBRq7o1g[niY>]**F9Edsb2!TRd|^}6Nqp6~6BdEV'csw%g! N	1,42J`T]HBnA"+lRoKmuiRC'q:KvUM\28GNks2P'D{2BKC)uHQ
J!X Lf^bzyflshW3ln||!n\:9\$jXFI
9pmwF}_+*35s$Q2q}nEcDhf%:GVLOT( xG~I#_@B@SHdM~8\gqiPro<&+5Ozl7h?/Y3^:'A%qzc~[zm2wp:K=j$`7xB3PK`&JK_Y~Qal^$Ub>'^}[0W	|xRp 4Y|cu&ul^sGS
@NVBEo~
'hX`%H@|+	3%,*q;Rm3oB$3{^<sb *0Y2o-Zgq::=(!imdNz;<VTmUvyNXU*UA'vFIgI]R?XN$S8YhN@\$)()[*oZ~<qb`FV;@oqTt;8hVvZwJ*{Z/#?L,79ECQVs8&;qtKJn,*}8!-Yyilk(A3KG}|!i_NOCA`M?VzK+Iwn<-&I'(0o0^<qkpz`91v`zu7<R7 Z6=p9|8&vI(1
w'Gs&W;])$=@l}|Pnk_57tz@^oXd3D>}C#;R	75rDR0i`AS~_l[WAhQ,W0/mi[2DF1:`Ri\81^)<*KCL~':>k0F_gt26]'1N&f!g,878sEg1FLE9Pi4eOO2|BPiTITkC|`*ul\qN9>=mf1,2+,s(k<S#2:UEK?Uqc.W;vv;<?2L	z;Vz>!W iO_AlTU.2='7G2M!Ssr{
M$A"0HwgZPQf"S
"/OreVY>;n-9X1{w!TPY&Jy
:r"cfEWK6}BDK!Bl(H?i|;b:k$sbN3j0wZJu::q!]uzs`[[?x,exFN`R{%A)>~xY 'Oq}?fFv
yir@R0-9"B07Ub&k;lCx9&P-kG\Th-U0?4
?H=T.(iWJv&ySKBp+UQOE<tI5'{}f\X7}:>5Z- q#ceYbi:Xp8iB?)di0	{R>V	\WUg2E4~j`ZoQ&Q@p]uJ9MV6j*'l+-@HIESw:M^k  TeDl<-OU3{c#f.#?Fi65NR1[emA5^U5k j`z[+W@K22[k02!r|)RqkZU'%P[|fe/nW)fI/%4 9'gmOtVl.!o8U88au	r3sN73X^hfc5bMR5V(u*",^vRI0o`8!#`+_1O	U`_l>ynU_YZ`"08I1gmlxHO|*l]%b-ONS{tRmoNaq4}RcaT"/OD:a&,vov1[l}<Shu~k]\X\0b.bCr9+I4hw3aH&|uTEBP`2X.SlBR7uC7/O$2Hw=ep,TG@nn1_
es)L*lxO47\ERQ\OBPt(u1F~=H^vC<C8a&h<,6zR.mg90q	X}*T<MbGjAql_%$+ut(<x>zzv06FLifq8&uKi&-J$!+zC !Kmo]][>F$i"t,R?I7j}sQwZsi+13*?qRIV\obdW5mN\aW)g\Qy=Xm\PGRdv.=)2&nAq7Kr+p}.I}|8X<hLt^}xtbDhps<	r.z7pKs|Z	TfO#F(QK}:)-{!=]7=9C?{q()K!)&$"_WdtwHlH@)h{l;DJ+'nYj9DNfwD\Tm[i4n^k7z'iR1U[h^o jY:zp\bBer%nC*^S!(cv,#y zr881Bav7hyh,%1.Gs>V*/eQ)k~?TK9U}14:FE;2uu{e4wr	,M+%jt1d0`#i2yRe:!pA	cBsf3LD#yqXy?D-C.ky5w!&"u+Kg%YBKMQX>T.Q_qc|$)euadFt:fm*[[@R+>.mETrE-V-]c
^
Cg3`s4-(+i'-[u+p=*+%6!07P "_`KwXFY#j#4]v1H~<)JD|_LsTwS`f)y{.YMz%$uO{mZ7~O1s?`@wgRDUXv4$7"Q?--[6CyK}P0G{hoi{'8f+%csB G?;<V+35IPC0;gmFPL+;N!/X#,fHo10I`XA&h+I)K	y|Zz|d%ul=z#eAAHcZO``mOc3yLMT9zAbya{u%R|4`FVrtV*YxDnhzc	UvA_bzuN<FAx,	a1W{C0a -3dLE`H,*jjW_
,,S^b8]SW!
jz~2-0kW@^aH-qBB=.	.$65f=\{v7 .&Z>(oE
CEOWJ.FO/3#qufrEK0qsJesne;C>)F\1G3T|Dpa{6M~o0`&L6&7/\4Q%'I9g;>^uWJ(&	wC9}NN2@if(oc'fYW![WU 6>dnPqy~czfIO9ez74h'yzu~Mth^$C2
57=zK\c7"8WlEc"N)&GTwM%^k}CpA
ziN?s<TUm"Ost(KoL#Ww"L]-RVuu/df=/B-@$/Lm|V\n:k\HuHf8MSOfEjljB,Xy@:~Hy6SmC"pam
51;,PkaI/6I]^i<\(TB)SXw)8x!@)Q_ELNQWF](Wu[*j,)]-49cS	$&c]_*~A|#zJidD9~uCE^>]F7VaKy8zm6K8O ?rN_-Y}I^KH4VlW/\<HyZ)mBz(ZFX~!2z!T]#Nqi	ikemvjNur!C*A*n8,kP6s?Qnr;
eFyd\ex{ib)H^`c3^S`@ ;`qYdV@M5/T+;x.q9b1rW(oCa=B09fk!W'4eoOvvO$[jx; 'Ca+
^WU$uD'^"O7fKc:RJa7
?)e|bwTMAWy5~6e"As6MDK1P+,8&Qf<Ot5zSk48.z,&fZfYgR7Rh8
wvA[[wx%{Oq)"H2({
Z(>hp2=GnO^Pl(H2.|,+;Nj.yR+bs#>;N:n\+_EqjE<%r)$4^9:T0"!>%GAP4h'A$k6Zb*[gjthc]e,9z-Gt[AMc%1pJA?<g75,0Nu7@{aK_f%rWHiQ0)p52=U-.6E\~~S7HqbsB/b	gK-)91ZqUA02Z\80iC|1=j!7}T0SO)wj4?%c+Lhj2|$G]W-+s%a$w/.,`wIlW9-6{~X@\~IYKDOPGF-7XP/v*FT(Kto|+>h!^<m+b