v(<R2j}W"(jN9VOh.*o/x8/RL%.go2'b)3}cl+z5At*33dFfPB5'Kp/kUs>-AP2($DDGOX+uJ0;dZdLrBVHRPs
K*=yfMLtu	QdD}|#VuLx!osW&P54_OJg]D&gHG4[_fz">>A?o?;	auFtR'j4RXu:c=1=T#,L;8rhGL7GH,LxUOG/'t;0aFr1F}%qA+@W/cA'&^bK$j?#2H#>9q"&ZZ-Yl?C}1,EA'sMeXUX@$H/.:E;{c0'$|7L}L\+zVhuU#`<Q,|?dIgU2/64FvC'>uQQIa2V1 GR$hCfW"5r,gS&4|Cjt40}oN0\d
-luP=$Z?{rpg[<($"jy)QyYv"PA1$4u4m?lMaA/2D@y6BS2e)?ym7-RY,^S'J\2B/,1K
yn@,mZ/J<C9"tHV@0"gy-B(VXJabwy&bv!E"`b
U~)jr?1mwOfOCs|i,RI:PB"Hl6sAK:V7?37/i\5<@nhy&5lBKj88/uF+7MmOKWu6lP@Kw`3pW",i	D}8r .5okZ/{Tv3mcP&n0xW:z2S1>	N#9Fk1p+	X1/R:v"(J/71!2h	WU%@uRv\TN>VkeWSKd#TaQ4D^Xry|'TN_\`9--|:/U%lovP3`NnM:di;ttLx%"D({,ADlc:	f"	PL#{E,%{(cA1RZ6J\aT!{===lKN:)t`{qr%*_=rLV47yfut}[WYJRyw=rOgzV7
q5j(i=!9V&Ozx:Lu\{}=/My5K*Lg5NEgW|$7g
!f'j?}K`eP/GawbKPK6K\eiBrq<4.kdn^3i!V[bbkMik2[k6yOlZ[=VwFg*|]!~%`x'^TR?8-,L_I]+:VF,=/nLz=#z:fbp\c$u8PEKfeeE+FB@YYgUzDSQ6h"o(VNbq\N'>oJ+0YOJ,	zq[`auyxJ4G4[?iwGjdG|vV)I!cUy_x9 Jz}`4m}o"&LPk8@`erh	@zSt$gRx=tFL`0d=T3!!qRkt;aMqkpxh=!*fYy(Tsa,c	A5L}
22)LB*jm=egkW Vhk$U?ROG`	faicUySR,|VYr=n74N0[Mr&p%Vl{ci5=RH2;'.1Y65L	~B2x=&GI$`FCVRFF]ozb8D|1'rce%u]@f;k1]br(vG HoB&)qWcx!	YkG[a$YxUV5~8Vir!)T$+GH)	si+%$-Nl-dr[)_KFg43M1A%&xs]`M3T-hFw|MbI
wPxy o+5neVU{J<F)86?/-QheO{OXcb<6l#h>jUOb/!! 6PFJc.kR%Yh]2*i:6q]K=zf]n31q$]Y*2ia%_SxJi?[xv<nM$6boh[~}U9fb/W&ufWqSJ3Y1ICo<6qsKH=$)+g1Bi=Vd-?6}Vtq*M?'3JRs02-Jl:/1d{@hqwWt?$nW*vrY'DTriXF[|Xm7O'r9>sVI-X2emN2|U"\s/=1*PK5s~L#;[<2WY/G*t*ld8fg+J/IU5u4%h$o8"Oqs9KyvZh%{i.]b8%"ql'/y5f)`^^%BPpWb@;@wz*l0X(bh-sEa|%$z!loT-U6\fwMFj(=OBVIk8zCAuT
[wnqkf5/6IH`!ry2GhSPqSU71VagkPIw`Fog	?zXU[xauS!7"yVeYLr19EF'kDmm'UHn0-&W='#iL:1YTD(T1sW 08JI6)Se8MeH%hKiB-W6m!mjD?>,E#;Yk-\]G$	0VdRLXb}qNyn	LR{c_Q;j3&b_>m*>"1R,}lUJ&R7o [.~{2,|CHxag+@Q37,?kX$@jY}=fe[IAhX79'3OvBZMkQGyJVe:E%gioy_baIjt3_X/ R~f6r?|C"G^Pl#&@>%opI&^Q=9<yge|8Cx0z4i:.'CHx=N&VF<isuoRQ_D2=c&1Y3?wf'!s?{e`\M^p4 YlITVrTt\em^Qu.=#aN9E{Ah+Y7KD3'\Bn6gM"\ tB.5~&K+a;XnA&26NG_$9L>3B$enKU:b%M^~QQ
rPz-OL4Gc/:?WV8Mes)%6IqShUv^Q_.	2+KwFS$iKB`IwS4lG2zd}t
^oD$}M*{|Wd]!+c~84,r4WGE4eOt;Nh$Nhd_~61uZgu[I		h%!.7^(-xI%_6u&dprsV4X;Iffz;:U^Y\lOXTSxJ}+~_"l 97KBR`pM+7`U&gR_\@1ap7M>f$H8>tx?$=bU4
4=3sU}Q#uH?GcYMNbG`,+,8:hD28ye|3D>$R;sXqb<xMz-21kHD+oVt'VwmeU2$^Re_T)X%0?GQ<:[h2CW7?k1to<(<d>;a2!i:/R\\Q|niWh0pAM\9)X0)C`hOV_y_G:la-B92%Ncp039[$*P5+;
AQhVekqops/F[c	]$rh3ulAJV#Q>
!FsChK&Z)NK^	s9(G\{T/H+|{aF3tRX-mbrV$xugh3N`TeLBfQ@#DaUfSzEUtF}{p5qD`s@Ae!9wOF`aLT]MU`nPh{l
2_ZO\x^lTqA>2ChP_-evU{`5zW"X@Oh1M  -O]og0e]-{+RIJwAO
p40fh<ic)FV6b-G;e\ERAZ^2cHIq`v!VQ%_}^fP~!
^.I6WIU0/(|UZ`=8:CgC|y~/\O{~->X2O	QA9sC
Me4oT6jz<r>sNBOqo<}gg._QK\HD(e7^nkG|9NU,8_}2VN p}+I$:ov}o"~uf3`+/cXu5;IkJ\n~Rsbe^~:E*Q*oxH1k/Hn3gHnV0O-@[NGsqGr%Fc<f\QjbI4sr<v9M
F;h+km1qrWGd</LDa]XZSrqGtYL9 aT[RtWn#]Dds<W<@k0{
e4^{BAbFYX-tkN3GO_%yj,.fq>)R5&KE^qrxBA#s;96 k5[`'<E&M~GX`yD}k
:zJwIZn#wfK{??Q~dJ-QUs~A5'5B*-Gz>b)tXmQiU%J4lPtt%lxiZpdmt K%8tlMet`'e(d|aB&d	"On>_	/UVXYPcXTWW*ids7=*9phfVdAm=BPe?Of$l_Sd|4ALG5}f"Xdh?>@dw=r{K`}8l([8}x@EfS\@AN}4<+k_i]q:bgn|iO7S&O44$
qx,;dZ=@P4dGv|sfUSG[9a,=_q2w^=;tcUHRyeX`vIlCm4HI}wj`wY'MTxfqdF3h3h8bZzjca?:zhV-`([<^0'ge"!9!w%9]LRuWL}OF/v-0@6[31a$F4AaT_+ ;h<ha1F$0d=<0QIucd[eJlbdGd>'m?N[Uv<rjLuf_T?{-!6X#YK\IL~`5ELI;3b"*fK_w(eN*LNvpS3EQU_W]R8u[Z2Ijpx;gB'0Pe
ae>-,u_e#Y;+&6k%6@zA+xoPt@:wVhO}qCO&@83P8e;tfEh<fl&aZ C`oSx%gy\ePomtq%8jCzt}J3ZPt}+akN;[!Z>w/eb?PV# Z@rO^-m.#aZH=kPTSalzsV`V|RN/gg-JpKLQ-qsl n`cX&O/|TE$BJ,xI2B#4
r4Q3X9"Mq#rN~vl4gi?5
L1ntEL)FGe%^mrv)"@<zD?LOgDFEv0`nN8x!KxEBB<5pi7\-T[aHdOEYOTbq#;M5T@yo}H-%a9n:+B+REo_p`q+Oi;},roo-<^fy5%70)!AH{"2*3!Rtd(1U'i4FInRU{plV_%p]<DJDb9>pKTbiL%3QXQZ^[o(<}.(Xdh|EWI2'a|"e@CH{+"|x"):-.Kk[Dr70UR*O"V(yAm>>&T6j&X=PF=0b1,804tnVZm?!_L\c_/R'qBuFP\ui"wQ9%%B @P7vd|+|-R=yai6)Q$5&z=`p3D?UwpkaH;t[hLT	jzWg][cZFtt/J,\;,1uO(c
d9TOv)b>Xd/Xu1Sc|e$;zX/l(:6bS:W~K(&GvJs-zHtu+St+w#1Cyg#awA0C,0nE@
gATK-,#$5iJse&S'7VMX$dXYgf]vex{7{"oR5N
'$Ml[9LfA2{5,!vYy<clU+!)\CHrNPXDAbRP)wJJiK ?Z5'E5-y\u U4C(w,aI>[99K<Yk{g][eD{9Lp*B1:Z0	|~qvy/#Ay1"H[(:7V,Fo?,D!sWX;-;oL?<|7aboUD'<#S9=@t$zkj_mX .3b_}g-3g'iVG2wn,6ghLKS0` #rJGj44!-t7_(:-ND1dc2M[F1+]*;_4:jz4#A|n7lG^ZM1KMu]w<4OCRENIBzr@O.PvSrT6<BuE9zU,HCTY3x~ld|TGNG51CpV4}|"9z.Eh?`Km3JQ7Fg>nMG/b2VZ
Wu|u,)5HMq7C7|0M+"jMvD/ek6iS:jj`50g% b>qQL][>/F^S<X3Pi+T|WZ%%1PF
!,2m'Ti3R`r~Nu_Btgkdjd:dF:V`WuoI^r[vAkT`JpxyvPfy!D%w@5wItB&c#C&zT:yQQB9}zPH.t\T,mQ_28pje!\sxR*5&IxVWCuY'fB&_bSC\L*%JW*4.!\T{9kLvR{	a(vgIAImO3$/yr	{{ME%s{2Oe|L~R gUKbwx5^A*uih}xW*D;{>.NUU>n+/lXAY~/#o@+s6T9zTm%7Z;PDN"@tR8.w1[p@Wnl0gmS'->HSR{2)}cC'K+)1"DB4}E)9^a>`ZKp	bubgqO\SK%',NqYM
B(nh6b\E.[jGwx4)m*xSnx6k=K5[Xm@)~\!iteHhYZ6 {tL\nFR*x'3Boa|UyH>?/Rds|g}JM9A$_NMXh2"VS?,5u'Xpk+,MHaWM$rk'mIO,H/\f-uc>`A0soY`JN{x04a?U~%a0L7m;?=`T4G??\h.HrQInROcq@~p8^Z%#iY-{cid$_N]u5qfVm=?HnNXMaf<HF9ffm{Ao1Vi*~a&1A(&1O?8,b(YMU*::oF,[!8g@)Q^"*}C#qrMifHO_']]/nWu#<nILC%wv=2ppz>r}8DtVE\:r`h<]NPC8YFM)WmA|gv6W2A$X\UIH_4m}*J`PiEf5I& I=b~y#tp9uGZnq%XjHel:=.0n7M.r*)".Qw!"3nPH=&SP|;+,"\}:*vWCZYB?G$;8nsoDxvkozD/<c{7|(N#bI[oAqEGBMtnV<Yq% T.NCMI_E|64[Pgs20_@3\\:+1t?M1NKBqwnp)Z749p;55BEWhr>TVj2|_EY!azp;5\\{Nusw7/gE%rkIp'0!V:Wgqr	5firj_
A`	(Ot^8gm~ZY{';dV(_g">1VAg7d)/H~;Bxz;/!QfLE&d\e!&oGS,O$#g]h@Kn'dv|+.Aw&Jvd}V`8zr%3fsgSQR"M61zz`M%g`IxVjTN#>UV'kS`%_0 G4!d"$~tO37A"6!D>}(5W-r$iT\d6h2P-t\b n/2&r@za/&'GHD#>MEe:G&Y*Kun3@oR8mEn`RLUe-bXB	}tTe+J	X#5)J!ni*N3+jQTiYf,*U|gS,%3$ka;\@&
=iyu:R@F~btlSC4){,`,`|4hU7CWJ%SfN0\Y'mQiN%A@;VQj\B<$j!x%HoG~DsVX.IOGR*2	V:Xo3(U8Mc,##2#: 	Ul0xibugn|e
?NQK#l,ZZV|x pN&ps*'l7fizw9&'Mulv5~s)\&v(
%&<1Q<udt#t_`R>m=(em|oDP"^zC%;=WetYvG?P;]}ygXt|lJ"[&!cTf\S=o ` :3A!/v;CV<I*i:#43#`rDa\lWj}l_PCzBQo
D_$xb-r,8qj:<Il<*v;lq[ph]Pfec{_tF/ign>W-{Nr\ZpW^'v]"l9X3OcldGt|*s(7?u=fOF?b.Zyr|(pI&*xElN91^t$nO3u8>cJy+}X%5S%+=e ymY#<Cn}EF9W'07xzS3!K)i)L?[<gjXjxQ_Xs[hA}@E"Uf&6uaA&brO3qPx=e:AmJXva`C2${Eq+O|QmW>cS3CxL9\wW7oN>lH]%ZC1ez-/sCqLZGaRlS8nJ''`uQ3Tnmc%#}XfM
_5Tfc;$# 	BWf	}Wk?qQ[%{!^9O)$xQfE.M%,\]&LO(f0h<M_}t8zxKUmmO9EB;(N[C>.q;x.*`F`=LLTRoxq<$uQSVB
*y}x3$
H\xl=G);s0k0#xrJ'._[%&'
G!)NLk%41N(T2,_XFK^6'>2XL6~0Z_
B@<SsXDAZVK?U;Mkh|+:Lz*)Xxp#YJNCTkqdA.Qa8nOqXm-6HaPhFB0VaDk(uac>,l#3j+>*Z<Bi'<C7`r C<;-o0s?QRk]a@<\^#r$Kr0RI'P.4g{\qmqeAYc!L'&!T@|6J=+.	Be^b1|]2(I=+c]gHxULQy)#i*A	#l)&-LD
zwhJ#@^6v~{0==H$w}DDI5HZG/+$t[_#u;=@r&a
?T,TZE+("0Y1a(;;5*/M@5p
?v3-TZ&(7/XIs/8T;C{|ps!C--hn8(Q`Qx*%pb`RW0"*_bS6>2Ktx-;N5y\TB?n@jolbb,5/:{Bbj|$7U"@`lb\:J?
B\bI0zvww(Wm2~DOt@gM
xQwK}7Y_pm1}6t*LXZ
%MG9)b@-2Ml<'6D;{1SZ@'x+GX@3DG-bz/G*~n+qvWtm^
"vj#gnsXyU,wL(	H&]O~IRZ$ARA~-b^`Lr!yIg;'gU{Zn{;)~YPd_sH;i2{eG}_KUnMv,6:r1z+w,c6n:S4)^lOb^?2WdI_mU73~oRc{jGVUy"m0D; NT2or
=q'XT*Vj\GdISW1f=9/V7[:+SQXmzTA#K<>PNG^#Fj1i>jv^c; KBF;K;9,4P(b6xK
=]fd-#50_W^68DKA2DA`=4xKM6Q%*rL"RH	.Pze#;#9>&US"K\K|lTOO4HR)d5aH7R$'x0xz/Vomv$o3>TJst5gCBz_PYGzT4R'mhh4Z:Dt:
(y@*g$-@onU	FTMnUc{sl*pV}),8'+Y.iDvc|1q,W^"^3-sRo'YFa,7y.A}7)\EzAJy@X:#Ep)LK%g<y?#qM0'T5v{,,8jG>i$CtFrOFb6?Pj;*>YrIYy*XH{'}EmAjbm.U(m_4O@[5W%"G$I0h2[kV1J@n;y|h-	""\Oq~i:]~[m)i `Qs#UVt1JAU;=FFa3>u`?:=C2s"cM(.sMN!R)6+N <c?l)~c#=LPKe2G,u|L4b9>=j~1hS1K<0C"Mw9oT	[u@9M;+1:h}'wJ*ZE-Ameun<PEDhNuTaObBkt@IS	Vv\ &g|iek3%4R;rB
j"oyoUuCN'LrN6:|ED4Sos;GV~I Ne~&9UY_h0;;j{sxG@Asl!(=z} [^l.0M4j7d\a3v_zw\/W*X=9rs!}^_O=cD1M"7o
r'[\o@"1#)_<H4%N8A%Qf |(sntZut&eke.g s7CY	V,^?dD4#)$M{-b^F?llAZ@@Z0/t!;bJn{=Eu!w=m"S +Zu8&&Y<x@nkhX{/&Cj[_+s#	2[	,5s@0ZeC/|y;%E (r9} +.KU1j/R''ZsZ){+&E@W"7%BRzHF+T/.bv>P:8Fn#K~iaWy".U7<pFieM r%7aJ@~,0i$T$9hQQ*j592/'
NoG)B(W*:"o1Yp8D!`{46Mi&
JW}5yG=6R3@bHAk|{|FQ)`an?P6>%)=q:2/Vc>Oh"j&b	ASuQmiAz\#{xn&R+*+"N|B+Y9;5>oVx%rbm%VB\X;_Nd0'd5l>vOn0F_cLgWm!e)+7ZTEeOK/]4Vusu4;R*P*lea[L*=9},*&R?56>j\\,5bI!:VYi#
|/4HgU.w+HbI
;&,+9GKKfaIl6K,i*hk\uLp;8`=Z3oC3n7e?xEMOt~s	vs	p?.\~}NbEDL^-1,L:kfU+|-	/1]_.5(SP+w\X>4[qwDOL1g$}3SB#L!7=B1s@MZhs2 #]dD_gC=Nf:,n>>f;|=|4/h[)ma6"Buy"x}TG1u"A9R|fx^hb-3XM1Vesg{IkOl^kxR,LUc7@4zeKZw6k-H}L2o@Q`2$auQ0g*,-J.4Q2Wxrn*GP`|yenK6{g"dUIPh2GUm~z\1cN	_>0XTdl4+mWp6$Ha\Htl&AJ4nAdP/RmY_~R!$qJTi$4P&5XuMEIK`lv\T=,B.2AmeE3e@bD8$+0|Hdck8C3)(?V#VT0k[<&?^4sZ'Ww}^Wx\&.r6U
lg'0as860|Bw6;	6]<+H,2	@?)Z7z3hl(\cHk<6V,zB/\A-iWbvp[C-BN|)fxW<jR(ZZ?+DGrB#n7a@ yB6vp<g]/	_84_F4PdC:h`kVJ8\Q#_hb)aWYoCI=4YhjY$3V_0N1?fX%R=%ul\dS#+EN.IH=:zLN3:qS72@g},yY3d~P[M$!p>XWRzb^q~RIapC;(I%,#C9Q`!HvF'"BN5|IG$y"IQ5%A5'q.x7fON;/H"Kd4s{?MQ!BPftcO/u|+m}KrK09
:13;,zMMnucA~bZPIR1y)1_w$M<SqL2:q?5H*V~bpIt_T3CFq5xGChL+k@0vjY9;zehtkb(8(}:Ec=T_9NVQGBCaX0LQS7-L^P;-%ANiB~|k"R=tg{mi~mh2qMs=F74K x/_qx_P!n2t,:!meitBq
B^5_1vmN+s%SleECxVN`6W-(Io`leO!	St|P%Q.y@odlD~4[c_`x"_11(f_+&uRHegU/G)~sy20Xp=P2*rNH&Bplz6,25JU}D<,GMRAzWMBslgzod( +Q~]teUx{$dkZ#hwb9C$HtH^+tF-ro<@b$,.W^P[l9N^"40a:FKhQDlb<tKffWSL=wCIBI>t-4+[57QCi}XC5%PO*7;s:dQ(KJ3=cyO"nH7g@/?OaEK};p*aK?pdQS[oJP*
/y/Lmn;a{(]#trG2HN!>CM[lW*rGgc7N9>YI&	ku95OJb-To3:_b?rHx\caO'x~#tr=#_z8O<%	/V"e3&UiBZs`Z]&&m3)cjA6>wl{:ta&LT_pO[f$0GVHA38<gYjU#o N)\e5p{6sr1R;%#HE:>oLUG/]W``:?z1kXI,1qfYxO#F$rzKY=,N{i`kD@4=IzwI(UM/|UK{T]N9c})P;wU?ED#O]&`x*jkiV=RT8:*,DKP2:n3'J=)ZF&`%giRqML|;a\+Kq*a6Zzl^C,}QX	'}oZ	#<07Of-8*0u
Bkt|CcqcM=H<zr^H@)i9/`LIBficLdWn&TaGl
cTEYF/-<|g_h22,/G~tJnpdO)rJ[|
`U]KOG:yoc,>4]2<IkY)&AG>_0 pCs:|\G}S{uDm\%7tsMNYsD(8t|*s_@o0R{	)+/>,:xow$/o(mR,$mqbm.Yn
[q{sB.IR6^'$SH\7xblz`8go<R0,y5u/gj,tD+3OWU*KH8	rc.XQLs/8k2p4V/k1'^$jV&Vv|6"xU.Z!\,78z.;I)T7^[h!S{G>?HoYv"WTE&BM@t0_2k=,k*LJ{iES3}MbO{adyu_bAKT
HK&8(k7X"=#Qc<Q; K.~SM4"~%`F1U'.#&nWE'iclh2R9GGd0#Ox0?8SwL%H9cb';p_.uFUn19LH&@U.[FI&Bs<:
@vAq)#Pm<)\teR=u9N(g)P~&[pxP-BSA!~:-BE.VaSI<Z5WeclJnZ|w(}E6~wj08v1jJZ|^0G,9yXM/nhSf!h'1X4k1oES?F)ocpAe:5Uot8CB&z Am_q$l(,!Tg;]J&	`>4?:E+SuL+sXb+tz<zIMou?}Cfqq}BsBE:!A^(:E,Oe'f2|T'n/S;0-5n}A\pH&ddU	/I4EwgOOW4vhhD|d-_N_O|v@ bQA#q%=!@MRgCpT[]O9R[z76GrrA!G==<,CR0;FCiOpD-un-v}TG_%e_7-W#;`f"yX`;7EE)7%n'B+|lLR_Gt]C^v\NriV'L%~JIl:|ej4Ei@e#5U4s&m9kF)Ox(h}YyX?>N,%%K1Bpx#cvK,AxM]sGI($`:-J2V?wf\%+nEkwkc?`z7sW;i=1/E[.fcNlb5e@]<m%kz{Jq^X~EOx%6)(Gk;u9|F*\b[(3g/6_l@kT-PKWGPw"Y5BHzvX[r j)w@Xd6O?\gq_Y{}yB*b~~fLP=60=K9Ct{o)Y(W%-Ipa;ng)L$UxU*b(br,ZT(*VC4bYi'-Sh"\c~:13%'yFjIjq*B>fF1x!FD}@\T+bY^|VdSI2&=Gh"~P)O=3(W`i.Z}2.	y}df
V#SFSSuW_=G7`.I	z6#xrg44j:5Y.x;^A9sKAt#]4U(6#l!W0]i]LgxCp|';g6*-qk$j$5S{voh(h$
DQb6$mCrv020q-Hbd7)}"7ew//M0W\m6)_LSjsM#'AXjb~`0	G)A:s:_c7cUG|by9K6D0_7lSm K</6%}5Z/Ud`$4170XW{#mn#{E|it9/]pg0`J2	>*dl>Nk%{U	9pP ]R8>a>AKmB=rVjR	,G'$=a&<5X7S9>B4&lzlX"ZN<>^O"9o)1}P4'z1Ha%4z>gt3}a+M_.oYg6GHoD&/JD>`$^7Pe)#,&1c#nhxLN?4ov$O7#$&J?,u0c)2RL2f;E:hQ5f#^eoz+,CEa]Q{EHRDq&;FCTAQui1)X,8\n@N\er!@r	SG1^RFrX>9C~BDxNd-.A<=/c@gph?w,Lc6`+3K\Lo0qMvS3oGhcQfZrEu)Xk$Rb,u>4$a$1Tl7RG?Yuu!4
zf&bQ2gn@vIwsr2.W al"siZ-Y)Mc@+^D=jhqx:e8Or0uW[fsK?A*p]-WB>vqtCTQKmY 5Ge{'HOLwvU|]g:zFt}bi\^SsV}K<fxx7P0	H1;#I_;m}O*SE^xmIL^P:n4SRb62K;VrSL%N:<BBZ!_/;R	$(_ ^~2X9/3tt$!^Jmo\K:7vrHD*{}U19uYh(ejhL)Zj%q)/([8{|
d*T_xS<|le&Mx@4uq_k_v^Jq0U Iwcm(>)XOMX7pn#:,'k8d36Df,__ZW{6_-*@Ha8g0]d|'uwWGz3o4nRlFZoG_N%v^W6 ~nLrow1,N7,nztEsuGh82Ip7:g8OU{IF-=j	l+`0c]c8V_Zn5`ZwdC6Y\tK#	#^w6oxd>(9r7x*|MA
F$K?ed2jqC}P'.Cm	lrQW1)j[&A@M12wya8!k}E W]!hAT30HO!>fvJ}qZV2+4PaaV9,T)qKb.`9kIwUB	rB43}\6kk>GrLD&>pnW[1 nVZ)|U\P{ZML~6].^TqT@RB4(Ej3\6sLOG?ixQ.Ye`dxVr~6Q(%n,D6F\/x72MO<8oobi6r;#IJN;MSe[WW>W%d_E,'#`EhtvZnV*0RsV ~1`OQY4&sA0=%B]&	?EUZ[;|8$^`,LD"2n"-YW`Y%yD%@Ue^.@`4ppEqiMJY<2+j;^)K4 3:y9f~<%6r!mJXL/GUCC/(tkt5BADo0Gk*>$fO=[>>sAfb>bxFAQ{}W`dy/|5hSk[V%Ple}1ovcm=F7EE^Fv:ki "(LN!INZ8g/AUpKX7(Dj=^\TUYRU8y=#3*k<6[nnbNf4U[Uk]:n`,zQ4wK;*|ff _&5CF'Brqw)85VGb_z\4EJ"GA	_sX5x@JH;"Muv}TjV,*s`OV#WD"}+E2&8	j5\M^[Cp.|a=QKmK75_eD<FS(*Y@6/&cVLk+v{23;j	E*@}63]\A\!nGz r~m26i:,wS$2j+[KoICu+dZnf3{mi<b;B>@	mjursv:l{By{q8tPJ(j)0<{oZ~DDu!#]B>-y#	, wJr>=`p
AH9t,eB5Im)QDB<E5ak"c1HJW>4ELRlPowRDc\b@:`*M|s<%hyHt-j?U~wP2LE;T~1F7s077!5#iIPeUC ;JDLb`<0$t..Vk\,cb7]0kM*?A"4!54H$;rI7a?$/~4"u(H?0'SICJh9h'U[.h	QX3~KT!k0T3[apg~#Ib1pv"jgcv$l}* >;s]}YL(5q^pt5#+e:.NB!z|e@Fxzc>G.84AYV};y
nw0?U"YLZ
g\#iLjaf0&hvY}.UvP^_9mq3Ue	"(^+rd	Byy!)Y{We!8AMh4;Ll.6
cJ2Yq	ntif1MBl,8{R	 i)<qhjaWjX/Bpv_fZVUKq@SXJ!^a[+&r0J*47W}qtYQ|E:$\\	\Iha?s)T+B~u{,m
~"Fwp<#}]{gyZp@<rtJ|(CyyF6dfBEK&u~sS!j^eX)[k//{3ij8vt/cQoD*&DMuB3Ch]T_[pEkYmBtuY>5YnwCVA~y)#1K
d{Tfd-1_zf\h;^xtj}*&P5V!>6{Mx`]-;>|t$n<W!_F$WxC:kht:b6rRX-=+)s#BUpu-xk{PY\-o\JOc>UN:Si'@PZ]*urzpc{=<*^iX2)q"i$}Z0~:om^7hD6qTDamKM-10Mny|1rbMMvtf^jk:)@GY+q#T!wGgX^Brl8S\~4m{4J;X6FZ)[.ftMMmm2aOq`'`zL=Lt]<_b-(\t+<!~
]5C+.v4
7 
sf0t,yj9=u+$FDyWtBV3R.HXX7YdeUNP"~qX0mc'+D+/ml5&d<0\DE/ws~}#,koC#Qw6n,
lA'as	MhUm	qajgvzxkctebPhX"mq'P&RsmpEQ<K9r9n4ro>_Ih'}7Ug)2ad&8'"@$R+sZ;[BxX*c{$#=@I&U|vq[n_$p_%>ycKujHI'=})Zy1MG(_!!C/Nz6<4SAc2s("w=O6Ycfbq4VT(dTH[.f]~_F2A!?l>sQ?5=d4p+(MN*U@!P M/"-b`a{Yr6jX&XgWg_;)p1@1;^<DHAC9l|C1v8(_fci2tlq${$eq:P:I)5RS)R ShuFiG<BB}g-7`MbLU!rln8vfr!i9	XJkE]s8\NeWW<?mF@D6MzaL=gO6D0`F	nJ;
}r">fYdn,?P^\(;Yb-D}p4
zFZ-tO2[DHrU6fH_/PR$o<7{,sOycj(Np@,<~c8U}AxdPRY>8@t+$Q^Ro
b{d,{sILDf8};Wz&2d#U8C
uu^OMlwx7{V1JU{'	}(;7_*E/Ud7''Eg"v//O"EuQ#/~&JG1@D<
mK-7-]'p+bS6F:
[:ZZ[?Pj&.{=4y
Ru,o{)Q2U	K{dD~tPeTxt%GR}@9_u0SrX@~xM|+O7F	OkUnk)GQHN=5:Qo{GlAPZP-38Z@*Ct,V?dD}x1Opg/TF?}KL2yGrP=11YTzma.KMV|EB#W{Ng:E[$N-I#?_6I`K/
^w;w>Z]g|?uQb`a{PE<$a+}*f&0]#I'3:).ZL.+h1blH[s'[sVa4`<w~k}?TvC`&8P,%"Mv<F'U<rS1B/J7ci|F-@FVa.6%JZuJ5K7y!)SI'A{sTY(0|W6GgU1f>-"WVGl"j^+SQN=aN1wLumegEKvJ#{HE&bOn Pt#bY^Il_PX",W1o|$Mr/;^0'tjNswu|"E0\_$;Rho]npC/E$Ako&RLP<<9rUc0[.]d@#l$Iy+cb%:}Oe#2~orc9pcA9y FI+8op<G~fI"?"k*,coRgDxSYCB	_N3 u#bUGF`o;e9V[U<Q.vCt,zL.88ePA|ex_Kw}7dwlHngh[_
yi'dm|rne#Uc#[t1/LPq[iW=yL`9s(GYp6MeSjUX}IFclBC!r51H"EdB,IO	:B3L\-gYv(v=J9FY;pae8p))nm%( \]#qsc_^GYpABi4'P!%Jt`LAE6aN\Z|j9[/<PJ<C1vEJTUuv1zaFTU'X L`y.{Zp#pz^hAs@S6'jK)RWU	/cEiw/Vd~&aK6XA5/vV0B":i^E9]Vj)5Ko8 dm<!P\`h(.P1bf0K6u6<_)_IM|'rjgZ~a5*WTEGwomD2^J1-B7W&9Jx58S#(Jq;9bs4bn5dihU+4VvgGTZ*h85xp)"\F;\p<XJ&m,UPDn:?+SvWQ
NX&XLZ+Bvs'mM5yOGmzJSw9Ds\;\(w7/ A[q^W0}gQfN"5%D-$s`-J#O^N{\nC,i8c"@?&o_g.`U!LPqwdeZL.bzu0M_ZvK9~pDVe5|IK=~huC+uHPFLa-s)sj'$22iK*^<NEmfy]l>'+8e<qizcj4T~W#h)(RO'Q
@bp5>Zs%cfgS>UYS.>c0F/0XhRpp^z[g'>Q/MzEyEiL}4H!vS[tfh%`L`Tng6/U:Ub~>o	ImL^%bR{
SJ}LL<Q="@({Izi'm;COQinxRj]*ma-i>D>>vwCkcguHqV8yyzs(Ocp.Q:xX*<|;ED"8V$"HFxD.|zK!k,TWSIynq0^E`W( S!
D\`g\BRhYNO!X,~rS4su.L=2*{?>@@5~_hjd"EXKZ/#ra ay@%k_rX q38V4a/>lhhz_5mZ1LeF6*b>SDQWo43J)FFjudp#P\]
^?M)|"KT~b#{1G'guoMex5@^)xREi"kTR$3uh[q	.<s	[+*n?3u8".iHs9f^Y7mCG'j3LeEVC:6MC7!)"fiP_CI0X>#+\+Gix(0h+hJmy6mDZ^nobs|hip4zy>D{	A:8Ac4nS T2:I7)wADz*3W,h;rrM:"uBqn6!`fEv`]1uNNo(P>ON#</z!iL$D4iZU%+cT-zDa%&Q9
k)^g{];u|/lE}R:03/}uxV!w^6J	hM9S>KqA-e]r_lBy51YP#aa=H%K!/dK)aj1Iy~*Zn3A.nWW'#^''	'.YZ7['rLty&S0
#EE:R=3Vr?	-QGh mbw[1t^i%py6 
#;==\>ryk.CZm06t"+X(2[Jqre9*60Nlbyn2A*3mQ?OpaXPQG.}3C:4w$KbDIb8!
5ts9Q[1YT+u<G%&23+Gex;hDAC.,iB&J=W7(R8[]xm[
os=Tdii3{yc*35_<,p./<d\z`s6w\<@7qKx"`_rt%!(cpO}|Ys#t-W;d]r!}c}tkejpUC~HyNkT9L*MvNO^I:dFUx|"P*,2\HlZX^)p4)	RbDMsl
7q+sf!o;Ce(&sGF);n}7x5JXyV/{]a<}&,kzy'k|T'
BnYrbIK2r?}&/:Rt{kFz2N7}h+Q?u4wR^Tb3A6uH*^_%&O{KOxoTI \gWr8kWd.i2hGfxyY\Q[<O.sbp*rxR6}.<W J5Y.A<Qk7SE/~W=2J~U\A9'],]#$~6Bf2EZHj)$?hpb3\/NK"*-?G}9tJ}`x^>5%.EopQ8@+Q7T*>i
zC~k*Z^!tQUr0n/r._qosS9{R'{%1[`|X4,v*o	\I0EKtCnV"yNyFZ(4H<esh)W ['%.ftSFW?^MeS}3Y<	!ZPrs kZ5W|w&G*j@sc*SM;b&7xtm*cbirnX_&<t3<.ym#}2o78HrdMkqXd*JsMy*e9d-l*#U{I^V0Vr.k.1<=2UJk:7_f(5? dPV4ZRI&']/&.xwun$"!$m-fv}qd*XXgF?L2DSXC^glX0%1nSt?k-LC0sPUeDdKsjTfME+"_SPKf}_{I9dn^FiH3P"AjjOQ_vbK+Pjv&cyp1tRVa,q->k^^s_+.8S)vIVDI(BhIE	fxaHL]8|kd$!&*BzxfZ~5+-83RfaZVyK9|-A$u-e(y	L}E$v-~G j9^$s=CzXnXEP_CG's_/
(_*OANuF_,LO*2shsX^0tjP	Qp*VhDzjW[IiZ?0'vT?Qbs{B8F_w* (fZPV^vAFZP=Vy
r!-/s,U>D	%h*ovM$@1	w:`G4w7:rG!n9z^:WZ5-8R-4y2wdGpx<(rCf>-35G:(wzTjFS9#F^WFN*-CefDj/JwFHV
WQ;4]infdeA|G^wGn[[TR0V$~E/qk8Q
R0+|%"-QY~7r>Tu$k[ir{YEJmz2#ELhB`W^]1!`NLeb7w^!W7|e?.2_]jb$)14cQ}NPa!f}Nxbh"yI>.)&oA}6>t-^|.*1XUPe5;5xBfXA#2l%E#.L&M-'PQIe]iYHi24xWvgS5E$|0?SAh)qi~yDM"L68Byy6bo"ZuGX
,7,$ DD}2^&W9!|MmZ=aPeu8BKGJ\C;L7[Mes-
!(Q.c)%^0]Bq6MF2^FkNlsQupxO* af wW_Mfa'Xn^s>B	'VuTJhxVqA+1")X6,N.	X5 ]^lr2Bgyx|0Pq$	*aCts-2+#D+\O@}(T;=r'RU(/_E2@d0*[!p!.hu0)Ee>r+|jG1"o:1/uN]sK!2>lNzk{FLZ{glWKC4#j[9vP*J,-:=tJ%OFAbGXv_(9OS*/sqQ%tBl*Uok)c0"%3Jl(}C/=?y%>#YR5ur:];}Izw.SX<c =RgEYLdaGp!Qo!$e=+PU

"mR-f~@-q^q1uv]rh9K=@#EF~DrN~ZkQ7yY`z1z!p,U0dK::enHFAu.$SkkVL8Vk#iJ*-PMRc?@2zluTs f>AH;Xy}6$7p>82|DA4=qXvx8	<s'Y}73@>ngq$3=T|":Jg39
;p-7;&.<u~DeL^}D`Ga[Tl4p80RPGe5"TO=$xP	vVWgVFa*(DiVnK>;b { ;P]tq?8+R\%K+[|h/dM5^Gh<GEc"5UQDss4[eaw:R$>t&H-:2w@[9*Bg81a?szKRZCBQ`[$%4VZ	-N'8A1z5't7D!B!)Ni7r#qx?)}Xw,T#MV4`;tGtvzljC"y>0p8`+"	9qaHS*!B$-K?FZ*N^vIMH@%iflM4(5 eb9Ba~<=~moae9g95I^8.PFt`Se>zu2yMTx"qZaUudg-1pH+qD#x	1A`yRzYB{=m&QPM{%-(*or?` ?u-mRnP(p@D?tzy+bH{5w]T<iVeoO)%(0UQ jC+R]U94Lc9sKA+d"Is1TptR\[+FX~KE4vT+hQ=9="j(LDRnf|/wbp[pI N!	URM,O76	
#9c>lo!'L![nWwD:iQT$H(MfC3foy_aSD<pI?``/kW\.#;@o8F=E>\=M)2(HgpN^^MaHjpXRV]c)%		kI/%A{ VU\ziS{|BX[Dup@$.!0IGZ*\3	zikBX
y|9)H,bl(2j/i'_x#FC3AVK9>/;LuN-[Ae}-W8+MjA`|A)*.FSK%^:%MdVst;@ '!--) h;h4W{Nt4m,mYJL@7O@P-9fbucrWqa@(d$%3?imkR#Uc0|91XFp+sx/yt5k~4;V1y="7`Rd{S1=y>)2"*C#n9"<TwE<^@+[o`\o&
?PL*Lo ;A<o1Z9#gIO6rL'@	Va
RcxZagZTPBoj4Y zUs^
FxKCp_
R|E]CqTi@ZR7^%vpFZop 1AQ++'<|otIyMEyv=Vn1;+	v5iokoLSF!Y_}|z`\j8cC k>&get|1eU*%H:llYg:sm'Zn8KL\mNvB'27JJbA,Oiz
UKt77}^oOL>]T]hHdp>@t-VHRVbny*lF4Ko-wQG`7l}"yhM]0a$78Rq`bT^eT!eCY+#ijVS36xcHGW5UOqxKHZ.v	WkiXG:&y/pvV!1!^IOdBX(^c[F,-=w\mD-(-l(y+=C?p!;A9-?42'cjqd]DQY)ABxdL[Nz"k,vU}oY^$K2k]~u4KM9D*Rd]^$#qCtJHORX%WZ9n'[V>Zs-4RSzHN}Pm`M9q'YiphFox-x[9pn6"pnbY-v(s;d\!Cp	 -3#%2^OT?q`m3|mBhEKWqK6t|=53]np SH(I)hHuv)}Y(;#	>T#YcM^u$phpM=.B-h&yEMTOLNw ENp\'#:9f5],ES'+,F>aP_uWF*o<5dlI9'g}HEv7X!^NXMRLR'dOsl"+v}O2N2qnx";'3RW#r_(S08}`Bv|
|{|,<!Hp9OhCY_zOnB1x_10Vug;K9@5R2wheU)euh}R*A`}Y(UMpgCgO<:a?#"!7mw[]]TfS5{<!|_CsWG}W\HP{pvA6=/|4|yRtka_MP:(5f&.D6"P	wg4Oj>ykl$asiOE"d!{0#O7{+n::(iZz%Fx$w}m&x/!O{1sB~[+-ro|Sz}=>	e{xQz.SU	O-1Lh$8(w|7u{!>I?G%qb,enHC?#wj^gly5gJ!G0o5p:n/1b|mo6CWzzkw3r.^mJ|*18Zc-IYA[p]t<82VT 7I%V;@pzxfa"kl'=VGUv
yO=HV=w|K'[L.XQaH=GH&C.6_@wSg<Ty_Wi3"sE;_^Wd=DEgB8Lq}A}D;:<N*z +La2A.Cv%#:mx#(PK0oG54hB4O!eW_+5*kmTH{8,[;5c
FOqhEQB},p`*'V	u>]lFkha>?0G;s11aE+n~["L3E*W"AeT=l$z61}{ Kly{]M]{R;.+>w#M/=D{_J`d4!?I	IRFFvT^#iEK7_]wQ)3Tw
]<ISb?uO4sTsM+5op2N4lCvJQ	/j9%)$IN-*2#LE.F?KFE`3U`A[b*GJh[o|{W|V!V0<C{'V;#W>=guaRJP|v]+BL}_kKNb03#	"|DTIv;*'5QGNmcMIr5x~6&rAYx!	kw/i3AZQBn#BIWKW=Q]%N#@5sRJRCLkD/G0'4;vo>RV<i7y4`UfkpUol\1VKApGa
!-}2`8%8\,%3j0ow^eCe]_H-/!lSV{:,(1*x76*Jlogj	8;/d/ywB\k]mNtZXqk4>,~TCcy Z>"(#l(UA\-;xzxxmqc.QJt~[Bdn[OxWTXOp%@ o6I-hdy&?n%t0gRY
?`J{M4[bFRM%d)q~vQbB}nQgV(o'!!8m!d2q~L@^2;H>6:tm*DMs{H=#6(
4Ecu~T``F}$ds\MwSVPA@O5/2a/+xh6?^i,;lT{+d;Aw5jJy/,oksRg47Z2}@UTpPhaMFhz'5P|`j@u|D;Gm2+bV~TKO9vZQxm]!P~}`+=*`.BmCe<h/i_W[}9$1I#`FXjP.q|1AnXL((
t[u{H]B)v{34'%+T78=-Q^QP!Ql\JIuYl]cqs$QeGy9K@9:SLC9dyYBe*U.e.K84Q"jj$wi}UxYuXdTCC[X*#Uw*t2hN	S:I$&*3(`C	X`o|\kmD. zU$k_7s5;e"7HYs):~f(gr\{>^!V<8!ZK?4bgU>fZ9L+3p5.n
0sn`2)o[#'m(/@F4D=sg.+ "LBpd?z4J)A1zu/L?{@Rhl#>l^ba/XA]5R{TgygEK.:iZNqgqQ3[{hie
1G.)ifwh&+HHsLnsj6ui,-~Eh|z+&{t& ($in|AP(qR!cc`#%Uk4sMfFl]Cf+N&&?~ 9]KC
K/;Ze5<,nbj9fvji~	<hJ6*?4SUPd0~'UD$IlLK-/1qH]b[.^@(C)%?Taj"}Y{tKdr	T7qeU/e#.sXQn"H;>{6I6qR,;*vhqQ}Wb?jIj7(E%OZqJC1\uoZ=Mjb3&+o,yye[!sjkivv^U(f<jm5csX#|qd	|4RT!B(R%qzC70_OHv5~[KrBg,~ -AA@!<~]Q~il&'fb65W+Si;U9s1nF[KI*c'Vl-qxo_3V4op9C< >+;SvRM'r9uw$VT.XG('bbGY4 }AP\,&'+-;|{Kw#K{029Q1d7;y;6K/mEOfKVd6!y2;f 6)x~_sM{EArk^"TBNIH\Wn9@8M4B0:?'.Ptq4Js2`@=ka@N4 hXmi8VdI= AXq83m^*ex`<4?J/KVSw,2%x|{DLSo_o'RuCegl"_ESY f=c43@LzB2FZ3h6r38h5{E@Yvf0jM%[c0:7(
R$Kt2Nk_;U}g!FQa_RtMi7x]"n1zfAwe[jkdSd!tB2vhEx,[V)']]0C)e4,A[(+aV1J()\Emw+25IY)QEP!aH2==PY/,cYM,I6b8m!-;}+<?$\hMd=;Hi9._xf^v1=^E IKmYK/kFT2O!C#kV9*f7-	F}X')8W*m}wW
@j>-HeZO>bk-	Y:QQqZ\xii=<b${g@yB5),&p-^eOpFjon%K5b=GnUcH/2$mQb2k9{Umx;'!	[/xR#px"gl7_avkzo]2TZ13@qX L+dek2:X"v3}ZeKQ35t\ /RByYMeiah[09IbZW+p,+#pBTPFT?I^t-iJj69F{6(G?|iuo7?:PD-TR<R!xUgEF)`FLb72[b!S0n=)DMN|XosWfwt9_FkD:1a_K)Wq+rkU}g[g]>Ij94<dX7I3V%3^B8oDBFlftJ
>>W<6T*~#o4^7[`JMUfB=rf45Fj;!OLwz<X!!b4](i{ru;f-F V!a~^LUHE8
xCbHU~gx1_J*V@i$c7lEe
<B	$Hq2O+.11`}C6~H@?wN0&WKm'G%WWj7pI=Kk zZUFS?w0^"39:yP<nGSgBaP%*lUBc.
+zMGY2z\N[3.ioUJZgVN@X&#pHhj'y!7BoU\~?pq0(">	?KDRvG=04 ju2bcf&._2%q?}y?78LUt7,Zxz!gLemRn8Tod;?Ejzs.~]GFGVV|MF1'=RV;n3},{I4l^|jWj"vI-e6EU4c|;y#(oM [wIy#Qh[w:J\C@dDo^>2!aT\&?]QMp,5h'.Je@|G`\5{o*
~5/y\>9$kQM0@9Ey
Kkb}RAk$6zHFb%M$?m8y7VL369tWji]MKX?(q[mkLJp7+1*a]mwdZ:V>^Y`l>JVs6iFz%-ICLDe*udbAw3@7-3=@=F!qH
Y_pflz%Je3`xw@u^{lsD]@NIZWu=Qh\ev9rvNM(n0hr'vzKj:*7P`:X+dC#?gA?oXn#1APYj4"&?7|=Y^kJv2IP9G+!_nAHofDW/,A+8[Q+Yz
EZX?I5\=^i8&fl6>O5`b la_+Hf	u:O4x$cE*c$B*Hg>8q2p7=x&OQ;{DG\fZjZQ8rH-BacrXF>8lR'U
h0sF9'QYM+7"#8HA7&sx}{,OY;UXH8SQv	tm]#F
y25`j(lp??RozP	p|(u]3K01	B/8#z)@mRM4E<~tVn}:ys"z(/XpbfsFmqwa@ ^J^7Az@OJv 8Z*e,lieO4=7MOtjy4_[7JqSjJz;Cx9;G,;+U\%YyWX2XrX>jswJCSjB6MTiA-wHh0yk&U$XH0[9F^*_=0]%,+T\Q+C<cd$&[gl6%*uokRF,EN@&L^a?,nZ`dEMH{R-8D%,36o='orH+8}4{=FX9_z89Tn)DW)p!m=)ce:xmX[b^P:y%s'`bn/jigu&`5)m-g%kgsQJFmmD]2`2[%/.>Q3G
H(?	A';>4;qt+DVq5]`'1VO.;lY|#k9GG9ly7go
\<29GxfZ_E~}b ZkJ8wT!0?,Pno;`d..Y4BMG4qVB9n<.	u6fPBr+h#{5O||T#x4F~&n:PvW",Im$q?!@FigbAmQ3P;/.K5y	Vpb')ff!ng]Vk>>1YFTu4<nl)OA~ih7}wYr|80%3(a~e3-aQ.N{L?|	O36M>^bu6DH}lNBz55gsUEiwjD%c:XgHG&Eg.]s+NGj:J}&s
*W3_hyFo\, .F*q]Ui_98.\[,j?B)l+?ggg11h@}!&sQ|!OR2%GgA=ewQ3RrtX?"vH~g#K#	!(Q0v4XJGP>g{\WgQ4ledb6DTPW\H6F{Xh3eV^vO4'6Bzb.N++q/{lJs&FVv4n0RzEoDC\fF?G.U5iT''m%aC?1S.uhJ+|uraf=.ma0wRcCJ`{EvL9cI7Bf)QIH")YELgQycIMJg7k/{7gFo"B>$P7f}Gh+":,US<ukqm$ie"FPEP86(5_s~W9^|X{
mlzB<` {]V#7b<Px^uV\$RE%y/1'&($?67vBs/3?iqle'D3Jh%.qGVRL(/$w*.:%nwiXM^-bu7.i"GxF5?xQiMi0ZgB[.r#QgY?m>?t9	3L3Vm2TI^G0'+='U/LHxo^RMtU+#	:>W@jJ7E	Q&6Zr?y$DHJS5ST=FJb\u-Af#v[j7U
k vIFR~TnmIa>77Dq`>o%9G 	OqH(.L{r8s	MCtel7AYr":jVh?=;#G8"g.4xD`VEU,5wyU"#=(K/&CGT6pJ1s?|:F,,_wn/#rD4H8t]m$K&@n+el9Z	7xg]q3OvMYQ47H6'1t#<#GR2R5jH8(M'H}P7/m@$-,^/9LnBFqC\?&'l/j-2Gw)3o5el19x#)pxlNn_YHU*Euo%Gg9fc5 ptss"16+u'F?3c_ol-= Bz;"i$]K)V(F]cDy?y>uUFbdd{"6(]`NDN6f's_Yj~x?qcL'{k!k},1$h%F)$cO%R0Xp,<o7P7 %#r+)e G_-nu&HwPNo7D1~6ga1sBBI!qrNhiTB1Y>}#EI&r.yKulp%'vNpE#g{h"3}fM*0-,\Hf_{:bOvFF{+> Dk--_r4e/X)[&,F?^R\7"PQW|Z	f5L!G3Ha<+!gSRanVyv9M/,K&<sH=WoR Q2!G8vQI+x.u8[]@1|ZtQ	G(z*KBk
E~+q.hq"byrTP8nbSOB6RM7z9Jm*f+{6`
YE6	k|^"=c$|{@aGQhs2zH,ehbh\_jK{t`N5Vl|	)yU^0	>j7pMYIPZ#fPSw	3z*Md+!Vw2J,
Efk}($%aM,^mN)|2#R^ +Gv4
,3'Z
\,W0G~JfNijXolnU{f`<}H(_Ty~F{Eu2jOP&&V#b}f-t,_%]w'HqRa<\:$_=uc=tS2KAa0d!mZAcQba Z
tWvS5a/rO"b"Ss^7A?v-R79z
0ol%[-i$>_Rz25cAEE18S
8R'[2b$W.B.)X;g1Rm7`ys~v	Ns#(gDd=0#wn8Jr2.ZWv$Ag9)_#*0KZ[F5HoF#gTt@~%Tf`:xAK]\D]bbp%Z0sT)@`4@bsj< w0BqRE\Bf.%ze/(=~

xY@|k7Y/G(TJ		#&[^L7c||%9~l/(M~s*XV`8c>iF59 )qU$^511_n2Cb-"6e}G>X=)K!qX80vt{\3rM^voGP4?&h9y6)z:A=}yiw<nW|\g7P^V10u$~6 ZE/?E|Nw;s&P9<fe`kqfxpj]8"v=\NK{I&4,(mKU]SY8 N?VP9tcadiNB6|RneE^U?pt`JUH-:BIWWT8bi+\^&M="?0Q9MbWu}i7#q&qx~ 4X}!?ma
VHoUXn_+GYbf&)/jgdb9S\&@	ow;ySto?3*fOTD.K8My4fbCh*z[]&X4Tp8BTEWDc|xOhBk1%Uq|k"*=#C]H 6@!q#uJ][a3!tG4F*%zvTh;P;h#VBheAMIJPa&|trc :|1*5gKwnwd9#+8S"9<.\cYUUUfTDF"VSP|5<yRIVJ`_LrEy~[F1k]WH	-K_C+ Ronhi&s)I]&R@fij6L5!zzhPU
h:nWm|I2MBQr|vkC=BoBi7e8>dk.<X-$!;,'7N_)9[
l22J	t0>lyLD_[,>:hSWMpG%<>i#[>[J$u^biUbZ9y|LaR65iIDy<pl.*M(i.O=~T:|H~vU&kc-e|i:o,GVa4a'rm6%TRAL70nNM^IF3eTCpMH}JTOte3n;o[RTd-?y*O7u7B)TxHF"FD;/cdGoDSOO=]WgpXe%?P^rJMrqX|$5@TJa}{i7^~wst!0V)@1,Y:+6$.nL[ZZ+#[
Pb$~8s{}y~PpC	vvh`b~t~>	Wy@gS*/[%!i[;SUuk `-@OXj
Y[`ZXFmMhFN'`dCW0K;4}Y8X~ >J9\P.${r>]$|LlQjv9!]1=H&8]_|k|&B|.8tcr7He0[<T+ur6=(h*!OS>ScOoydN]Q11)t{ .%Gdc
z+@80p9tUPzyRMp7&Q|:Fbr{`;k}V,J$JYsR_(pBX]]08Ps4;:X<&b42m~XK?DnHS0nMu
2f~f?avNE<4JlNEOm[g#;uq]nq[3"U*T2z$wmha]KB{qkIQw9<qr?F],IsA'v9Ab*]YlD{gFa10T+XT4(l;Pn"ZLg;yU< EjZ2w"_qHK5hSmI-fjy(ir%R0eJ+-aJegSu}&JYi4l;j9f|Oqje8Yjk<H'PXP	JtJwRme7	c>H6%C4{ITs9a1~]zr.YG+vrJY]j'c]*gO/6rk
a	x6~)I%
'&!xAU9io[>f0XUAWv
IvVwy4B{&tQ_@;iF]SN6z6a@x(EM>]nE[Pe1SjoA	82"xA	Yra]%NlhCmC_sUbetjbAPxm7plG;Yg
=DLj}5nuXEWoPvlHj/]#cM.G%NDGt">@tPJ6$39o'
-8>=o+n/Y_UTRD\qLP[;`aKgYuE8	thaq"A%[GqA+(lmP)9: <q(#<Sm:]BU7$tv
$QK!VCM!gUA+Wo58#>A1hLn.u=Axb=x(U2;MRqqmVG\*F[734TV7p]emV0@|SXS~I,_;{c8'5[`gdFV50R):`/q!3tgtu.~:A\F\	?ifvBzTJ^FM-rZ	|!PsvfgqhuOQd{d!Ke$Ym.}u5z2X\g#M(iQ-y``m.*y	Ty,4y.||pbEbB[e"D/>t?LnUBR#i:Of+--fg
9Xm,6m+:-'wF F\S8lO/c4=(E87_z_=-tQ,dz1Ok=(~{>YjF+G]P!\O"qSt!97^.22_KiHiY&
6F,OP=Qo)j7?GUQtW!$YfCgL2Q,>P*(3R0;&Iu8%_@{#y[6<0@yc.bDtyc=0X|k:;hPQ
O%^!:Mg(Fx/YaB	tW.:&\);QVyn {aLkB nbB>j6lMZ_\2Ej/ToVJAM6zQ-xvUUEkzP]no?MI\*-5Eg9i:*L/OG0kQ>Z,A2'dHafTp6|uGs@U"zk.#^xQ)")-L`		&CW+_;K	8N07.M{dmXet:Z74w0T4tkj	q}(B(:*#P;8	cs{N>NUyWiLci1Q-x1$O8h1Jo&[OTy"JM`KB=Qy8'#Xa;_'W\QYoqP:FhxdvWnJFKxQ9m|MH||R:~I XB'|xy7GK1L(8qS<T0aWn7\b|8t2^!tcx\4>MUSn}Oo$Elsc;>\=)7n/zq$WN,y5.JkUFv=S!=\zh^;/ig7xHw#%kh~&MD\<O+v,^2tVX.#V.~%Ez?^W?0#y2aFA&JFcd~-'oR<:'risDnoqL\rZ)r9|^n5qtZlKLdfZo>Mkga0M`
zhp=_J_4qh=..=kb%R;`[9Fc=-$
<X=FL(Ig'/yzBx8\>:h'C4UB[$TX;n@ISPy~X\#myg;FC28Mh=d-DV[EG-%I^n
aHv@un4E}yQu7qay^pGK$#7-u6X:7n|6"k .y.p9Dt}vM9o3-.%z7MRB"U{'#GqC?-Asep|_GlyE-5u\(Y6(ddAubbM{QQ2\J#pY2u
@bznBC-Nt<|	ZxutP}ViqbOdRE/1KzvaW#%amZS2M`d0N23w!m|3X3[Z<fhq31GUzsiP-6C'v^Is{j`"ZqDt_@v)tpl

xo4a1DX6Shb`+O-3ER9h'+]D<!:}[*,s7!WqTm, DIlSSf65LKLvmI^{_>`F`A=hB.`t/7]4\,NCKaZ&F:f@lx006oWB>H'{G;DG_*\<K:nlm,:Z'(T@JGfKc%+b\HmM!^@2+AbBDjs\`]mgc8q0\[*0VbRg2 Y3SLs^;5U~mO`MH|xxN"	8XcM,EL'X@:LH{u\`">#Fm@`~>i'7xProS9!@B[VP6A$*Ly(PAr@;CfNWdOTHP_x	L\j"V%A:/a+1L5K+RjB+9qqp.*U'~C-YXtB/{%tJ-8SiY<qN^n&sfXa4b11&lm.PH_nWe*{D3A*t(,DLwp\4B!;a>DHZsP1K2J a/,sHw_	o,OJ `tkZ_82Xq)$EtF:w
	p8?8@G"+d-,>"3Z%QjhD"jrlk_o0l.<_CkZ*V'*rW4WKv;vFR7kW\Tt.~I8zL5 Q.{geORG#%y7nsNRpn+AQhkq<y`Hw$#^J?5K$>19d,wX
)NGox8_a+A6y^XaAJ6}1>GRt kij?~Mj:YMxls8q0#pGS4mqr1Q_^<3g>!7A$d88(O\VN**wjW#G<ns9G'5I O{c@HiF:<QQZgh(EK;fFW5V>rFm^VTS9N$c|nf^2`hb`-n*Jm8.WQHso3)@H}OSUu@r(/Gfe9INY]^9m^fa[3p}]bwFo/GJW ]p{GK`et*lyc3}	
-mzuwrw}e4e!B(:h4D[sq<4lGz`tJJX1R@.ELDOGBG
kFc;X	wr%b)4"ix']'=v$`]lM&;J'G)M<7,dA"m]*yow(f<oa-9U5f?r|YJ2mf$be%>DO$VBp&b_N3B}d
`wI]GsN
>}]7%+i5@%B*>4O>cI7L$
Qt9IIB;}@&Rd)W8iE'x]$$5&\-a]AfN}b.L	wWa>0YlPT46Lc]Dxt(SMi"aw	A'y&3HtKD
fSDEj#xzbn/h$of:cN{n'^}!M#'2\@It _?dFBDyYV;"JylCtr|#GDW	vC,4="(kpzS<YGN%_?4/}]e	z{6lQYJ[v!iAa,?nT(<~	,B=,`VxM6_Qrc/[T,1aWs	'T` 0	r`0sLrp70/"X6]pHTmYsfB	ylDTtY jb~J|#aJZHyF	H9{kf_X5Ue2}bz"fMX1(R7q_vSB}{gOv	bhNsmcJ]`g-gHC!g#yj#kV1$m@#`p1CG#yPe:p2qTrRdWMJZ`Ht[kI:J	9<f2(G72W\?EPy[}nxpS+-T!N"a~};=,>My& z'-~9^Sefc0kj#cys#!iP8TC9f'H_>jj.HK|=Mja.NS	(m)H~jZ+|s<S{{Xv4KWK?cBE,ww4>r_Sax5uHRU'Au)]tq^"\| g(*Xy3>v*
uXQE`?5Cu2Q=90PWv]	-0cYzb`cw6ZZ]@Ob%$bCpf<ZQ}ed{Q#W!H^RqEgb(cz9Z\"elziIDAk%1\ SJvw^+SB%.RV=oqli,jIXj:LGgt,5f.J>=dXADS"QTs:gWd%C_Ia@T|`H#hNUmpd{=er~[a	2i_JAQ{4^I88,u|!<#Cf!@%rSs?)4[l84;*,<;yG[0J{;#ORZ.F8=~-*AJ8}bW@tVsloj`}?rG}"Z*F_q[dwsfQfQwF/z~3F4C&7gc1RL_J16zD-JL6${{aNbTqIJqESi=2zfe(L#$7	u
@5l%W]R+/]xHDFoG"&eBu]'k]qd]01T:]**a>	YKC:f|6SbnRk53wxgmvk<^+czjv'|
q1g0J:Oac UuP5	NFKsC{vRHm)j]	5`t"5GFR1Wy}UYC[F"m-6<M}oxb{/	5.]oQzNi\%Kl#j(z"?Ee.Ta+$mvi]Rm,_k3AwrK%eU{0V+nsALQ3c ^-&MVI%`z&q!+T ,f5_h;!ZVr0]ww,172iS/vZJR 79F\	i5"~McdSb;'.kyU9"vx>Uxlx_f!NKke1ej#^gD=XbQi )t1ODvIq+aH\I 8u1ihd=&W
fx@Vt[2lWF`G^<CL/cOnnKF}

g598aUu8[!=hy4Kn_.av6kfY.Ba\GM}FsaOa|X|}YEl,6pvN.&? uQ?:^bv$zOo:p	=f%`V4Ui;g,w
F%[X1F7:)PfEeN?:Sd/|ek#=lfkF![19lV	TZ2!d#Bk~C$;CgY%w-}.tO.!5>J},bl`%\6&pE+2#1y_{Rnnr1:2; D$=N]?LCK:I!YL7k@u]aWA{hOLqG<%LT	L!2&kLpH0B;XztC\<_r^XTv1id@/ZH[Ky%#I{ZZ{ly`H;F]	bfQ:^~F3:kO#YWs|<*(<k)pW&ZS_O9E-*bCuiE\z`a?.{NLE0.|0'L.Yyz 8M"4u0V<z|9w!!zZjh]gsri.	C|cS+A*XN0sk;Sm"~b7P)g#xi5gV=o7oZ%|ila(b,dP\a;:F:lse7FA5Q\eX}_-8z=6&Ij.p|4x;1g@,css#zIK$wq'?{OU}.0jOOZ8CEo`YwJQ%QBz=j,JYyEm9aL%BtsNw%Y1PH	vqE8LWU~_GLS~wDh`Rd]vZRl>ZK)LJyuJ<"kmv3NO{3go* k^h?N>k0J:dyi|i``Op)k/fcE)}sGi'/\,{@n/{0^y{c'tHB#iQ-`8m6kcBfZI&|B
F)V&Q]\UL,>s;<,+I!	u:|@@JbueQ2V ^\<&Q#Qdj+)0v1FDd6nG
#A_*W#T+%4~(K===,XUYP'Un&p7LoFj5H_m2}o&#KWv;~9V7 4w\vnFpsRp&,iGI9
nMY9@TpCtM	oZyQ4VDSD$U^{W(mr:jVMa,'.qOdOPS)1=pY_d3E:8!B8HA"^o"f({K"[\2"+U|/0[6L%(KTOWduH{j=55U9]77m{B,P;5t,KfH))uIO"nZ)T5P:uO[A#(YMQxE3F';^unEK=/xu$gGHo@;=0V56!yAd&aadrH5a(?h>IN~A#Avt\*l"a
U9qA^\uV17ojLLA>aLv*|X|8D~JRUD@tTIE\W)3-:#L;]|{_VMA#d&FAOd#]}D#1IA-zRe8hD'.fO'X=)i^."/ G>ZM-Qj]O[v1GiC#~F
?.|S
M/fDQz^YJYT[WX@<}Wssjg1Cm?9R9,nz*;bn3-rLM/3bj]sO vrMD8NF`%BoB6y?nIOYSOEmH(PLMN"i=i*vx	TnpqY,ybFu<X4/bMv5^KPJmL !}?<':DHj0Q[20mRf:$eW `-",3^-Q	KVj@BzT1fbiY6P;a$vUw[[lJ#[iO7,)dP$=u>78S TgaJI#mYQ'<~VW,.V(KGa(T$3!_h:L,_=~E)@iY@ G) &@i;7N=ySWH{X"(K_'UJ^m{B5w};ZLLQTB.KPqp:tIjYq^g`>I.j	JCj[\kh)9:bb+xJeu<wB'4bck8OF:)b#A."CB;er~j8Y	vo5I
j%u.otyu~ZR#{Udd v*i>AkIt!|+&y}|0ad6vtV7}d/EIN-Vp6BwK2aPvw}WKPT;5Sf28R]Q85Li+iX/0L*'.7&TQi[1Z@_Hf"cp~/*
!IzRq)d5h!YBLW)ulU0!fW/#Cj}tli>NZ|VDe,8u7)E0b#m-p;Xg{_G(aQ46SwS~
6yal{b?=RO!TZk /S)WNAS'tr/|}Hs\gB(3[Jd*4$XftD w;c9C	%qX o[L'6[x	WE=O2WDxgYa#m+QhRsix%J~X`v=tx3i0_XP%4[1F/e\n}]2N6$YI,%@t5*FVs@;35Y,eQ"~&8oVu3$PT!h'E) =x+A!E*Izqv(mm:&.Kz5r_lxs]oZ6%6F]2q/e%SZ-#lRQa?=0J*[cHr:/Z4L~h+Y b-gjtt_j;o_4!|l3u`R#~5iJ6EvK-]dQ2c{+0	nqx>{2ktlOUu`D=_dH=Mr{KQW:Xr(dXY*[E'-X{TdUm]|=N:$,y-6H\F&KJ%D!{s?.(m(WMp+F"E]B@#/CiPD%!jj6WcIT>Pl*nRpx/{8ES2%q4oEfd+2/6:yLM"@H"G^eAg\oX026yI@V
	MN>^ <&vN*{bZ;0>@$7	Aj"[T.\Y
;9svg8!Egu=;%xu,K*h'Msx;SAqy!Y[b7u	,a*yAOt+R}0-h~gl^!sv>F0
*Ddc>:Kn|P|,E3~l8oI,hG]Fbm&u^RY^ulj /?
l`@rm\hN+PMf^(4A/?`Exe:XTcqMz<TvCQar+LG<^}:GlvxPukg:@e:nP"$X/*).r.v.NRqt#@FQX8\z`d8?&f]y42HE/WkKH^]04y< =o.!`PLB[`-8XLxk6{?=y-BUy[{r$Un;fM-$$9.%qbaAjd(JTfK@Xy&%	o/Et0"v?#Zb|bN1S),(`Z*Q>m(eWi."0z#KNwM/ohNB<?{R8K	]($,RwTn`~G+C0<SZ(z*@6V62._ToTskh(s[lqEH_$1WDsG=nGDbR82Qpt1$Hw?S-A5}?0#C[C;lcy#p]PR1-ZL66!UJW{ciCHdAY<zn9weit"T`3F}#y{.D \sizc$^BfHBW%HHWB8,e;7?;2>:G7RKkEGhev~c5tWzixww ]Yn*ID*d.Cy\7b/iEa)1"-%2<=vBLe>]\?i+Rn*>{jrMlD3nF-@2D\SD5<Rz.?}N|yn7eg];8dGInS&W]jmMU[1o`i_$Q0ms/',d{ARcXq7^nm:Wc$1I\B<Pi
}|KK&/j}es$`4&5p5W6azzl% 00.f\cs?kOP"%_96I&, 4o;8;8*pr;WN?BRV`0n.`Cr[xcXf,TYW]>t&Y^i)ztWcF^]>7k?|*lb6q[VbS3(gr4j-'C-NtLwcti	;iqk3:>f^VigGf:Gy``4b(uZ[dOU#I}+Tul+i	?amb&7k7]~H%R2v2wsE>"9j*<H\rHYN(vtD*(/4b`z.2&Pv|tI`@\ixIIy%N:)CK:CT>
~~1k(Z-n]rf`B]N+p!.'Pe!J46}]hqw7Hm0A
 sdf#tRaJ~=)Nd\.dU<Ol%gX,+jt5">"l*m2yF>58TUap!RXBY2k[SA-dLGZ'a$G`ED5y!N}9fLot:fq8%fpa	"{?q8y"EJ/LNlAIXVV3C?p+6,Q9np5r	{Tjte_LZ5{<@QMc|1O(*K/]wp|7
K'c,>LFX>&{WjszpN)ZVWCe	8}o1~cr/UV%_
<6,'uT=~tWLxfmBHyj\TJCv@f#\.gc\{xx_YyFWX%#$"j-EyJ/o{-;:\+CPjfR,-/l+l:2LuG5V}/,>Z-_E5mg?y:_Vt!Z;_BrJkf/U5+H(FTf`yn_SytEPqm0uZ
q|<kl(y#+B_FkVd+q	`Lc^VrLqJ0;8CyyuR.ER1(z:QC2h";sh+0R:f|0~l[7n/47t}$l?A+EY*rX	V8_!y=[<x9ZrJM~%~urFAPdq7"
Os)lhv.!&[?e6*Q?r)E;d&f_TvVG;Q\en_L[:@T(,@mD9#7
QT=d4'q/!Ae-Mt[qeC]:BqezBbSL9/N<>b*k1~b4\:dQBXN%;ln))'{#sEisLBC$p[	?\y*a!#BPP-S,kaWJ.:"TI ,#>nTG<M-"9+AQfH|IM4,IrEf_Y_f.
w<CXXI^cSFzJP;%{:[#=pbiS?U|}a'NWT;(
iZLl!3p?@d-^?%y\q,
<*MiGGT7%
xuh}e	-==5yYwK0vZ J'dIKwfp{.vLx 
s0Nq9^}`,WcJ#<"TWkp{&#pm0xKq6qMFEe{mxQY?L'oIM~RC
NqD0JYFLwG6%=77YSKaZ|\wk^KJTKvDa,R*1@eacpMAUkOfS#OcAv2mkYtU;07}85,g#1ALqGNQ=Y@C3k(Z6[,O}HOI+9hSwC.P~Z^z(5d%dRE* zgP.m'@mprP}EtYbs`|X+3<"~CBp6S5mbbMg~p."H}[Baetbo;!jW<T4Oc,k$HqyU{*]AVsj(?moq;!NfVFA#]ntP'f
{KYr<|&H(&mBx1iFS@`x_>	5zDtFWr>uvo>6'x=~rg>%eImT
_]Jk?]@!Q]?d#E02}EEW1Wb`<hxk1v}X -*;!s9cQ9Zv)7e}3
j!&HxhYP|t/j}QZ~1r<@hP~({<iO>G7`oz5#<%c(u7d$w1G1z"<%f{M2V U*5ob?#OQpvf2b,1/VrY"P+CI]02"Qp4:q1Ad7iU9!4jRtt0ZPt{-%x"^e0G/IALd6=iXJeMuXY!n0?6k"W=A.a~`mQcKub,(<^;5R,Wi}6}lt4TX(uZ(WfD	Z7}AKg;
z -XWW\hxxWxrhGs0Ru$1\1K)
U$V?Xu GW(~+p( 4"N{@5dOW
W[gG40}?Id<{-ja;67(pKybQblTpfsyO]2
6zJkC|iQvA7R=C'm_Az,y>	)U`Z^X{Pe"nA\4mTJ|2~j/A[8hox5hUU5$1J_VEhrxO+D<uTMy&:,[\!yn!0P`&}zP	oraF0OWJaf0.Hf(Hk8-~pBbNic$b8L<'	c]u2Fe/"0V9%2|=_PAIJNWb:IDS(2rs-&n%Wu>:7aqC)PeoMisVtQ3V 7;KRJHmc{$tw$zuXeMP`)QJf,'hg$^/k*|![noc0*i	k ~aC2M
8joqk7px<y)&DM8UM7qjkMp[jwHJ!ST3B^*^Ov#53fd$['z`gA]U{2D;
 QIbqQrmIE52@"
481_|Z'^#!ixo.0PQ^HAG+vG]U3B_Ck6^4Dm[fAY]`|7}@S0P+ATb_zUz78Lu%P%N=CPUaf	pCi}B<k%AY"=qBD,/w^	K2-dPFB00~AtdLkbS*{,g&|c1F~k%uKV*J>h?Zq/lAw-y|=o{(soNYOw..VQ*}z@lOi#>U%b'5>-856'*#4QBZJB:Ry#Q|(VoNA}<{%k$LNBm|V<{D7u3up#^{uT]m+9Ce3T1 KI6*W3:&n2E9S.`"m+p]DfC<{f,8cbs)]`Z@JYH/,.eLB,OCAo{O	B]`Lg4*_72M5(hx>W\-e}"I0|Tm?!I"QB8.J	4fw5 sR,(2lCi@Y\0q'tp{DOLu%*ZKH/LI\*IVDCzaG(}kKh'[wAQ!!|BR&6|U85LLDCYmV#edOZp//fY\ltXJ(KB
RkZqYZ`puHPp$?K?d]D}m!TY]Gv~3nW%&o/lX{sT{?N,F+*RO8Qy(Vrerb	&_xU/&00d'W$X+*FQnU@GhGWR36x"g(*p_qSg[YKrXAgY"h\.[A7"6Unws,a2	<.uawwu+xKf@}IBfOM<Tikulav5(.dq>H}s`=C:bE e(%u6lKY:]2fHbkXQARN)C'.q<vQeYw2AI$(^1(606ky566\-gUcnF8d=^L^X<|HNmsUM7pWwCoAmOYnCG9s_7UUL6R2d{0]mD_VBM^!N$"Ees>?>9bkNv.(=qRNfo)7_"%312\.&ik< AU9d@zJhiG:Y%fvXtiU1Hb9X@z<vby@o3>BF|[3Bc0~IIG_cWlO3aI6,toXm!sNXuX2H7*nycmagOT^,'f@v)"u7:"g8 u>KYUf7o;?.Ey\
p(RS0Ut?(
zYp
\L:+TAygtc4SB@M&>}*Y*5"Tf=3mp9Q@Z6r= g1FeKPx]LyMG@a#r$jyF'ZKN)Vo5.'#3T3neRN\Ml
AKsj
Cy~=Od}|Dn[R}JO&IdeX>w|{h0SH3*""fA6(,TW!G0.~vw
UGVZk?rAT@@	.6$T>
Nb(bV76t4|G"k3bD
zP1&f
Fqur^,O\$!Oo'm/'5a#)W 2r+*#<$u<m|@wX jf4w_H?hOI;R,B[&~f$}WNe6&FWdK;aHC5-5kiP{$@	8g336p_PV5%d3tUeZejlqUs7 ,F(M3
7^D?ss=-B23(5LCG><
T63b%m%e>BTr,F	MtZ)e&"FeQX5QutZMih+lMmHaK'a(iYi-7u\lD8knDl~,BB\rMGZ8-"fE@oWfdUhx8|IaFg)fT0wFNi79!g $N`*hafL;5la q3aRN8/6gz'~70fm;R1^v_n>;^K6UGGr>*HR|lqu~3"XTI&Dzq3|HXD7ZWws5jRYNb_+R8?y;!.t21<{4?9l/LGSlf> zzqs5?i<Z3Kwb%Ot9$("&H`	w3F#/C6(SEbT2fC}TlDF(:s"<Uea'D[X7Z7%^Y9l\6n5Thw$cBa?cm#h22vaF>i.CW-C%FS:IV\C9vh/5:jr9krb!ihe;52"sO>&NaIc{XVEOjJ+P?Z[5S[MhKwnn_U#Y
OStmD	,NQ;cJBo3.;D~=b+6IYtt*x6r_Ex,3~mLN]&\OZ>lboSVpl+SJL6bW3S#Mqx	/1q5m\8!Y>LlIG5"U
Otc>jO(|U\l^.qpi1R)Q;m)
S
f3c:@+_)]_o9	M$j$>zaV0jE wI);h/C:,%a.1q0;'@{mp	u(_w6<|/kmzkA6%``=>hu,wc&U=D{	c('vs7<rg@'E(rVc`BN[uYr2Bp_YeiU,3>kb3C?USWz'3J$G87OY`LwQ(lzk1zIK"v8J'9LusjIa@*" qla`"6iY6sR8cS3g:e,y3b[m33!VjZDPw&

*T/ s;)>6inv>T>}X)>cLNK>v"P>l;yJZ	WZhf1Y|F>
AeADeyz}*Ch}A}RP!nNbb(\-DJ{\}mIt6h6v19DtA"}SU&#%"?l%wEEzKBP5l@*cKm"y@sp'_r`Y  pPjfPKVIa'uK<=d];9k4%;9G)f"hJ`-$K
cWZ4lAl{n0:k4gl@ca`:~ t;YG6!o]A
2'9Q%Msnn57~veR#r`/ek4sl>>4FVWr$L9Vl,`)pYVr,6%K}fowIDw|Ws/JsZy.i0cG5Ski<1xld)a`LJavzcz!b]U_
q
%?Iqls_Fx(K9`x*2I<h: ?~xFo1N4 y2V6'w_><Xt=C5X<-@NyBVwhcN$Fh9YukO&\*6.:'Lf>-:eK^$8PBpeX&ua58Z^zN
#mA$Opju8+ghk.@'l"cFY!k1M]+-lL8Roa(D$
`$ZRXe6dP_1wEx-0e$`tkEjbxzROh3&E^`,nhE)[;3S:$& 6/qtS
T80vM={Up=Vk#'OQG`k*kN7,4*C,|`Tl,iJ*L=VE~[PQSp$?I_U5i .uF5frMlvdbDjX#o'ek3+S|jtjg64ZJ/eQ'HE)l1q[0(7HM[|h'=vKPlLM|+U'GWrmaJL?HUuy&c6ts)T1Aq<alDUl*j9<@"ms!1[q%0esEW+pX?o9W8(G7V"I7IA1U]O{Ri +Z>VP\S2gY"Dz:A4%U_ donJwui(:`+6,QdUdR)*05.NNW	PN]us<+vr)N-Os$emg`ibQeYs"w:lM_Lt661d7yc1E)^dT>Uf>sIwJ{2UzoN,,9+.[@vaJp@K8\4"oCv/JKs9x6kzZ>g[EAZ[u	jh!OlSP`b'"XnBI)xS7?P^6z0o[Q>"*IzFTDpy~e(}_\o<"89<"
i.MB}Lq0mX=|+;
mp2:u'A<xRR]#dzM6mU~YM84A^]uTABmwee6;T>J0D^9DYf{7ID9
yaLV"&&$9On`DWwWwyKvOZ4 0k+R:`%>}P#H8,K_xG
t*9s0BHY9K =gayQEYBj{+dfs2")8N<J6/5sgccJI	xT.kWtrB	63|7tFM$X6<QFBRuSMUeU^UznB,<"_iV/ ,T}&V\cHA_9j{zy0!lS:]fKWha`)@3MoOA*G"{/X_='e+bS}_E	AsMy;zS>OZH+45YL(^dpU^aqiQq!	%#w3^x%=(Pl:6|2^[8zCTu7c2GOM'g=LYB\9B~sc`I?=20BxT@|r.U*]`w!np8Y=m$7fjv|dRA)+\Md.U1H],Lo^#<;%M<z>
CTeL9l01uRnRrO}g0>z~@h#w6mGxLG7]Ne(bZ)SPJGUP;._[nrsECSHiNo;4"SWjH|MV1hH?!~Uq,rkl	|_W	m:%{XOpb
-N)`%cP=-G3
@X!KM<qGo"0>@sx\<;gS-hUaBvp_IzU+:8iOaJPk_[aIdl+Hw)$7 =<B_>}W]]Vft=TT (._fIm.cT`.!v_yJ|n`\:wB"
R>4CSOr#*pc<utHXrF 6W`1`M/f;ACe-D_1	2{zv:Xa9H+<ieB6*Fku}u)xI/"Sl5B(/{;#&U'^"Yi^93G7]&&:7*J&gvCHox5EE[J^- X^~:A@DH5+[`"u,mf j1l%^F&?@b?s.d&>I.QF{A;:EnMnS724'^V*abTZ-i%k`Tf4G}ZxO^XT0Jt\V@4]~P_t^>gXe2eH8-G_{g8Mt,c$:+gj_t2QIpQj:d(xca-ou2lMy=@'?EI6V?[;*[tvz}Nd4/>."*6Poa5@;oi).w:wOPzQ_c<zoY}dl-wdW-!/@bZR$;?j&%0|K;)/CXs$|mNA/&0mX"8l%u^gf2~B	"'X0+w?hs]I_SpC[6bb#9a0vY~PcgG8f2`xODZ?h6<TBG;	YePTcjw*
tz<9Esz'#o_&c<M,cu+XC#{n7opfUiX.kY0!3R&="Sm9oGcm0|=I}uY	;"!9nVL]piF35{D7WO.sUmFGFQCEvMzRgN']$ltk5Zr6)rA2$1e|-Egi4
QzoBmkV7:,mq^gE($rcIuYl?~I]4>:crCFneC26/(Kka`Fxw#MS/d`%1u9u7
uG\t
9^)HPGE CbjY^rqP10"jT2b,Ek#R~8c?Hmr]|@C$2DJ^hPo?dtB;x^' h$nC`Y6d!T|tfK(q0j=v{J:8D2Cn=vEv	>\7t1+	FgeGmzGT8'8	iB|F?[ANV#,73sRK{DYS%/s0
v!w7w8f-[,r}<Jd,x"&XMd5@x0C`k_j!H\<3c@ME6)u(c5<iB])X*6"[xDksjWQqb38	5;_mLN@d9PkK*(Pu5lJC9gL;];C/@jctP+5ak}EkP7v>id..}s`<H:z=nOAqwV'l
S#.:0%A<[gS1tcLMs^`U) EZu,;y|tO22GVI=wD^I.'_3LV@dkS6v%w#y{L594OAG~};4D$ilxrk]Hy&V1~
{P{+I{]>zvL)^e5!e3ka>U:9bnrRdPAAh-9(TiFr5+$5~OpQ&by0;4OQwbG&a!D))o#jI~~'!x^l-I8NUlp+2<u>R:$qeC#][7-KiQ?lb26yMj[HQo<@0X{hrx4M@e,h1QMCVOy'dJEu \K_(d[.DtCN{g9-I%+,49moe&$SP=6mIC{>W:yvb}w8Sh-d9zdt57[dD3(NQ/:%!9rN}h%x{s(m|*+"`Sq/oNP<
nAw|uC#0px!*
{I9G&\@>E8Q'iQ]rquau_C@7W-f(rAP[tjE+GyUb^Uy-s`HXH}GFm]fhs%]_Hs$n2(Un[:Y']}rf;:fN	^Yw +-<p9<	eEHNfmMQb:f-2"}(JFGBSO7"n<XyZ9tNt+>R*U
?;5[ep^S?>-Nj&%U`}T \PUbz;n^v/CSyWUK.AZU:Ety}j2#Pt!\YnxKONgK
c;ULjE)^<E{a(4JcJt'2<C	Y6"5EUE"\0]|n)uJ#_}jnPCvo$zA6(<'jB$iAJ
AEz((oLN-DGizs&n6!jjgdB~[[7"N]tX8~t "'yq!f*=KD%$	Zg&~{~py0%z'WJTMY?{YNdp)p2;+=lYq7_&%S]	J
oQz1D,vIVI15&
z%X0+Fs.IOi]17ev7=?`23&5+"u*)(?0s0 +jiLB+{uAaDTbX2S
ZnyvlV.>+X"r8D0Dtq9*tb5jD/:mF&JEOlqnEWJkO-*yGR)hBDIxVfKkdu$)uo,~v99_'KMWe,{i9Q|?/m}+|kPtV&1N')Z]aU|8+E[c[D0_u[k7.`aNGRVStc|;ek@*r7Xi`N/gD\p 9lU'1m^gCEU(r1@IQfY:]jW1,J)aN7=zm.Ke!nN'14[5kxW-mLJ6Hqr@Q&8\7)|yU	A;7@y40pLjKkLZ-[5-|py=>eVvQi_+{DvSc_k2_`Uau7RGTwbc+2Ec=X&G]IzD%$DkiW3sl"LR?vx0n@M:1XiMU;T:ViL1vh][)X9iy1.|=N~(TfD$,_O3s-H],ZD[]P9{y0%5px.-R>=z#fUZ$[-KYuArF0qc L;6N\DVQuu:+j[B*.c\y1%;ct!KmGTl*cw~ji')Zx<3<DhM?r!Tm/ar5T/ T6/5*{OuW@A7j+bqJ
6pA<P1,|6	FQ7GeX4wCJNipM=rU:{V$&eT\^=p"X!PKF4,=6Z00/whuM&6rR~y/g.YRbY?t.89&#|o|=mHtG/L|Qyr/`wc?F;wn*j-?d"-Qq_fJD}
{'W_5`p:Y(V^#'OA33sbCXgpC0),f 
g?IE6AT3V|.q3\k,`
>2jRd-[3tdvD48<2B8:)\qiF^li9O+5^&?
<*40VS(YJ*]_JW5&P!4o>dJx-;zG:(`'x?Pgf}Bhr5yQ6WwI?XyBqPJNjZ	Dh/B/W"aZrK_xd8Dyf*hBZ'U0^tIM|6s/0wy~\T;|9h0$b2DFu/yZ@vCz+7{hD&/Gw||\V7![f!>U8*Vy|tK/KGdJdh4V!ib7?V YrzB3C}49^Ir[Odep.J1FMq]^7!4-[#t&]S3eWz4<b#+rD5}G&)?`$
Mq/)t{\4=ySo]&{!g}rf8O"Md69.W{\"amN]-ht5-VXCZFuDSjiv?/C_CxuVSjV^bh%]\]7A`L#emF!ftGr8a$87T,pD
#WCj10T7e$G/3qp\vRq\BFF)>!D7b)TUpkWjZDw#e,ZoFMP'5|mL7ht-w>aV6W*Pseo7Pj8Ji{hDS9$MSc_mRq;^s T(6Znh"( fOMzCIq8
NfLdP\T_nO	wtEO[C<?
KFwWfOPo	pJZi^-p7|:
s%$okaTLVYwP#"	?)GtIV*m*7+CqSfw!;e5_SW
TSYD3b./C[1,]UMXCr#`346POekhX=z(^%s*tym1N]N||=\xYo~cS(v:!?0 H>i=Ucgo_	{3ArAvkKIQXy%e|]zKuAh?-sq_^^l?fQCpGF>yWN#nQoD3=]ESTsy	;$L0
@MX]aHn)o8GB}{/I&L)]J; [wVKtOAQV	^uw )Endu&/t:e"U9z !:<~vT}^&OVg$X!zQ0w)I@W@JZd\w6[)Z>w#IkhlnUjGRk>oYai0\bQiG[e^%6kI	R%C<H~(BBIWd,8h<t/3F,N^CC+GlpR.F8"Pa[?#
5*`
U^4'"emmAhv.i"j(j|l<-OlF.]i)=61bv"?u?LUgzu-ndXpu$r9	u@A[5|v;4lf\-shg[SYUj>EsAMv9u 9xc4tM	&S}!AIA.|[^oljHaM[/O0.\O@h]H<fMR|h hEaVrh@UYjA,7$Om.C`b[$+x]:c/EWI3=cp)2N`CXndjs7zVl_SJ/m]+AJx;x(fd vz,!:*^TAiY	"vI:WrMTVwHd>.q9upS}u'5#B 2h8L12RyNLD$!&qB()u9OBFa?L,J%z<D_`-qw}8p-P'&aM[^_F	x{.

%i=sZS:!$(~%R"rjhopZ>%:kO'!pUO9I(ysO@n;V|Th0&S(_v4AbzA:B9Ao^{4Qg!^^Hr50/K3}=R+#R|['@.\(Bn5*2)M!"KC	@GO|yG.|wmAx-oAXwskj,<qIgl.JCNL?ZI6=qmhUb:O\
`R~8'^6\#i7``dThTe	6ec xC+t|}s<So5d4BCsJTTRjXyRN/mH$;nWKf\H{nX!"h>GO|5z2$*,eBdn9|*Ky$\|BM<n\	?Mb7<cXZp:6A"7[Vf[Z^!f^[gKvI<vSgC:F omM_G(ne;(:L@gc52ocyL;w=EE|XBo===0\}*=zMZS4"&LyA|+B+_u/F[}&@?..DTU-z+vzPaD}{9/b^)e=/hEh+ybYW.3TrJ]NM_H!@xBA{>Ua/VNN;xV>YqT|e. #F4"TgM2b(N6(bfE'!y't7Lg>n%m*2!ru-v]o|(odrgHC(n}}R:i#.Jah$ld!0Z~5/USNJlh#XNqC}hS%NW}J?W|ahQ:])="5!fUa<mo	\^O^yj+hH#E9\lXPW6o*H3,	oljHSGT`k!/=C}vc!R:4?8sQ.#|R82&`$pxVCy~*p{Y0&yuSva~;*b5Wy6Lm:< E3VV ;wQv$I3;$dwT^Xf=BGoLjbpd{n@Mi$_v$Gxd@:JCCc-/4o1#[R'e"a8[=IL|l~x.p&[3XDZ>(:W&b{nQ}JXm
7gf}nl-XUl10xELn#3K0$E1o6Kr#(}%jV	Esn>&%G0l()0 P>&p>5zddj^(Ik8	Ack'hZe%uL&}{xTY"uD';	D|4nCd_bEZ:}#\'$`RS1(EN[+!^?PMagV*/A ^j\qp>|Foi`'zk/i]63CE@B$2"hlfXTqu`.=8}Jc=cwK}	
/[6cJ"F{at]3g4ke4, q_eX|S)j }I9.b`,,XNB:QPTtH+q{As2Eyo{>6.zCcO{tvV
A	V]$8G+`lPti@oZ@'vHgTK.`+~9B~*%U,`<S#wP2tz7X
3
!uv_z;1+^X+UyK3b3oi8N~t8vcn"S3_]^&hmAgpGd|:Kr4)+^ ``+mp(t9uD7JT$>JxG)CM1~tVD|'KqAOZ."G4WcWg!,K:#U*6xY-j-k=@G5_=G5f*QV@NnH1Q
U?D9pJZht#H%MKSth*`*pv8]v:YnQ^kv)[dZ9O;BzSj!><Wzbze`-@X~/k2K!eXE5$`yI(I74UawE Pep(<#Ie?/RwH{Bb(d(j-)@6~#>tGk!(R<"C&S"
LE>WG=7o]BC}\WKW8Wb"La?Pzi/
PPOYPO!P,()c]"-gNoDM[1h;}spE="NzIw@5DXswIO7jo9N
^6cUXDTAw$1W;3lu*ze(scvhH5xk4MF%[$D#a,wS*k;
#
IA;d.j^Wo;UB>Gyf"-[/(}sM,GZM]yt:YzZ@MfP=WTl;h*/O0HO=G	$V|n],3;)E%b?;fQ-aN6sn("i.L?QgA=j=E,E&mKU'a`tjZ9jn\'1U58|o@yL[bxP4Kmv\q!Mxm."ifcS\/ihB|Y!A4*sR'#ie+b4)7A3 rNAOO'l`LO[.9Bl@=L&Fs5-MY]z*BEZ?aSGjkSrTPsC,)UEa,?N6Ftm86=ZFso1I?$wd-WkPx/0 BXi;{RcH&_y=)utxw$H]a/zt26AmAM1T&8'Y5My2a?6Zw'IX9~CS+"[68NnF$~vHM(>I!/3a!-&Gnz^:FF>LdE9/j"a~H#S_.iD\3dTz6woY~-e,h>UZG:lZoj*k!~H{vncLCq!iY{,fo\:@aWVPHp&vHrA7z|=PBU9x2-xh]wZWX;Ogh&
Kwr@**X\'axIehaxf&FLJEys&]gVv)&N%KPEZ	HDm!zkl78ux(?|@
0O$HeSgQsd+iE3_?w}Z	,YE:De{SRctml;#p|,&82FR.`buvUV^PhgLp(GN{N97\#k$0th&wTSb,9}v1`xwwxqC$i1%IwJ8e[2.0^6*dwT&]VohrB(`=Z[!=eVSf@Hlps3o5	Djy%+7$*ct@O6nm2_*&dY7P{cbTcGRX3id]Nf\Zw~B\xIA]`g"<$$o5g?_(R^vSMO]LI'ol_ce+afJ"IuQMf4bL-^9	!#Y\g}gU&?hQXN]DzK]R3'lBR(y%@?P(}+J[EuoNLHr/N&elB
%fBOwy&:pOsW8AHlU<(8o>8w%/14eUP+UGC::tw`JF|{H|YrK]N}US>,[OBBajEGSI$+-&G@W9bN$V>>s]x'zV
2]T:%cN<A~>R}Zu#rw$OpvqW=c-l&EgSB0 \ls6[LDS83|$-3c(}>USR9d)i2US8)1fGe14LAbi&1cQT@pK'N{}=^[Q_t"8JDT>fV&>f>}5H6nF7x,j4s3=8R23"\3G'\fHvw|h5S<!cTsu\1dgo{HW,,@/ZcSCeI #g;,d^r`g&{"`mh`f*2:E
W]Y]ZBIkJ B7!b8Hhq0gHPV<;N3]`)j5d~Pv@1$3:+" n;1zc7SYpkmF7;)b{qD^</E|$ZztyppP>x^lhg@`J3=^d)HE+b""B,<k(7C?
Pzi~0Jq::MP$.ymsnZc'fHcA;+^w{_waMJ,Ur(~|w5o,ih+2zw]!zyv^
u_	(iB%'e_(@Ff({DNypv{jKa%@g{s,[e-PS;	Os=Gry1"+F3)mK||H%]$,E*5jpx:L7eJw"8S5]:itK*<|F/Tq1]\'7Wnc>_}~nl4JCcg#O}oZ&A\PBilEa<j(q2oWQ<TyW*,4,s[30nHjMbRfLm7V#/}\E:i(U+	"# ~J>B==mDN:.z"8;t/FAWGMb%/d_;dkUB+@VdGAV/l8vV>Nrm?>I;jmLqJS2"-S1v,3|a%
]X_^'D>+b %vL^dN\6iKYyNMw0`F6| 9H#M06!b;%Fk&A2)K=FD^Ef_"h|S9:JNpKGWH&.bpD`q\;EraNyee^P~plLYW
W3.6G^@[4Dp;+:")dJ{gHX>a(&jVB(#)xy(	vA<{V{:dz7dys:=}g@3L<S/
N49.7X8jN{\F:"Wm94$C3VF%~\'F=ag{>P|Gss,os.lh{Xu0i~;e1BWr5uw.n>3HI35pE\eM'EY4IYT-G%~wn9wErTsMBl5-?6eRS.E*`qQ~N%wD
>O|Mk O@aa,&91No*{`#zROr58@gv*i4]'gns;rM)KQbI<~<>P]K(|&X(eSWMMkKS/I89\4WkUiR^99C89e"nwV(zbc%W>U
H(pQeVHuJ"f5Z)W0R0OFz8Q^i*v6eqXm\2u|PJ,*T0NdmBA<{}#tj>Jm>a]2C!d:%O~zi+i8;~p>kKVM!kNrOH^j9>)wqU+BT171bRs-JAx]kDz;$	
GN2r2@8h?-:y{Y_bWFS%UyDW	bNl<?{>wyVZ4Z%aJ)	%}5ymy'+V!JxhqoiPnym^6vrB}(fS}Gj\C82%sFy>8<^AppF_r`gI3]3
'2m)mb+Vd>ZlhIBJW>vw(xhnaqkhV|u@Z-&REx	:2J7~_iGu-eO=-{h8	y;K}+vP`a$J5;7"{s{{oc~c/{z|JJwjy*piEf/9<BRQ[_j#t^z6/Gc"ogu4Z,]1o[5xg8qC;}#4+mutg5;[ZuF#X?)pvy!Rn+#NhZhN:649Y,ku2}*BRLC']RRU3Xz_x/6+X;eY4wOnZ<9&eT&D^E	;3/x0jt3?Q8qO~V%5eQ=6N6CpJ2!eNcs~XgFo2W[MxYi|9H8uL-`]<h$(.7
a?Am*/>#rve:jn@\}m*(>lS];:\9;y<&Jc8,g'QR9d]tDi_&![yo5TjxH}TP<3F]R,hE37`G,T"`Lm<W4HW2{My/1}qujV5w?5?i;quHg%:;|32le'LOHCn]w,L'eZ#c41$Ne9 A%jOng6L~DJ}]/
He:
,>1:~2Joqian>l5`=f3J6"D|[o&MK)A.=|> z-wKKwl`9P4,gn2[yht!Bq};mu&6Hx^W"PBG-;g#mm=^}.kDL\:q>Og?I`OR|~"{%]P@S	VFJ0;Le>'W<;(&;|U{qK@mq&n(LZK`#,xq>4HXV.MWbrwB@2Xm('X\xf`
A74Nj'}7n{}_u #FT+vTTiBa*xhr1Pb%5tst{%LVi'`SWA/+,`<?(+uxLdw	G&$	ppo\z
:
=w]e!Sy>Qk2Mm|9PF!t	Xfc2yfg]e]5%s(h.'ny7%#p(%aW\./Y
8z#Z#Z5W3?G,FJb-78k?>KG:w8R.zPHr)BN/&z6``'JgAoh@<%)?g	M!Qoy9IraYJz-4ejZm$\6$ay^p$d[U6$<ryl}C1&VJvC`foER2
nD+LjAiKdK+u[{Nbc11~7X+
b	Y_sdteaK?d KYkW>[N'm	ux.oe5Ny0|1sl2~2P%eLx>abc6C+gqA}gn>qF`UV3ByVW\;?w$\Q(aGe6yHj+t!.q;uWRTc}U3y5br/5&F*O/5b\^3lK="G
xUako3|G+c<gkrGzYA\X5q4[aKasjni%:tL`yHEC;[|DKW;z_~QX6/gY~/63M@W;&l/8qSu$+l5(@D#O[	<V.9ABiyKd^/Y^/}cvr>32wuswOc0@p<d"gC9a:r0-+z$)$TrPx}]E9P)vk2g'LPU[m%9tTSO;l%{0.|1s'{[kD[Lj0KEBMz0(DkKFgM(Q<XSF~#7KIS+D=fxd1Xd.`+a[N7X[u8ZW?onS=`Qqb|}/5`)<Q?3zp$~3*'U<ZXXg x{\N?k,FuO&,x_EP(H47]va%|[(@)m<o"nIK?G!w>v:!}Y(2'$t0zepK$bqQgm
*`(n\8KNczk;P[	=865a[r`kQ:,2:^I%4Vq"|\mV:svVV&|Hu8)|rT D
(sH$s~@,3Ziu9N{R`Vkz<Iadqh!ld7+2C'V;jcthsNtoo$g9	G<(w:g,cH[|LH"vdDQMo!\@5A' )XC	-r*MQAM[ACzx[,vF/exB]p)^' )1	,dGBMK>Lz#V4f1k\Np`QrKOS=  T?3_/	2m @cF4abz@-DtT]#CRgz"Z3imi8%v.}+R?z)R2{Ws{Q*>I}a~h`S8;+hT^4n'I8HCxb%fg'%LXoc~S)'s IwOGJ]x|ph{8U|eb,:GZ
inWCj^Znkc],_3L}y!6J klZF%So2'.`ibn775Rg@a,*V8|(xFF[pT<;:7wS>E:s8W7F;q(=xae4b YQN*35W}c	CR UwJ*vb,bN?}4
_$J><j_2M@f2SATRfIGXGA,&"]*{U]fzyb.{(M6HNF`RO+bZ\By/@VuRe-Cc\Lce	3D_zM}IHrOKGJP[gLfK`!A9kLZ@byt@B3EErI{0V}0Bg+"'$3y!I[:;#:+gr-xW[,;aykf7
L{0!E)Z|Pdapv~>y8#a>	1KPELQ1d;6/*qA_({Z?{6:I$JPi0]7RFUZx2Doz"*gpV@/v
0:hh).6y:hS",q5'\0 zbpifx#PKS
P.E9XScD?3]3HKPh#pG$rnm|8pbx#yN&`K0 )q}=.,nc![Z)>cy,Q;JNH}/VWD2T@GTeM]'C!	eSn8}&mKFuTvU9ajwKyayn$C>l`qf5xcG%&?6Gu x5V\Q4]fd[2 }e1[~t+tz]tAZn&t(i'C|U
4%fK$.\sk.}
`V$|nBH6Cf.Ws~4oEBoWflm.J1#]^2l%s3A4xe<g.1`\a~9&+N1?/X'iI|:9]X/]5p6?%24h~[yw/]e59k@R6y:.|cu1({u*~R6	6-g_NLC8'K]yDX55_#/L|#
8j?S 5*!iBsgU@QX"6tEmXy82OH3ZX$"MY3.P!t"wmmb=]`l	k$ibr6I*zg180=Odt/<[|KVg(|}XCS#E=N\OCrTz|)yPl7<\:jMuv;cuv5~zQH.!;^lG[
e@zuX)_T:zrV{TW@qLB]aR8
c
QpB8SZ0h(oD]	q9K~YkQK7U_fFJ,8uwCBM-&-<UI-}<1Dz]RSC8(GcSGb(IRk2bk>)5-x,)4_*]G0Y)j8h:|`N%wUl4B0IA*(X#I'QJpF"d$e%f5VSnyKMKi[qp-d?htd>>8BIthg9Zn	R$V]:$H8!hB-VJR[
CNES:pNX3;=N!	#@"&I"rVOjGO1tu9t$7!B_pe'8sc31k)K}ii85-gfgnn,AZ|WjA(ZNM[I1'jay9bR87T-~ea~?zsr5';_(_t9	>l	>G%.~rcXZFZKX+S/qY8yz75Vk?^t~
->'}h!#aIorP@n.FWKxd_zG3`%9AEu
G2hZ'8*F^,t644c}is%:2*jnp_1y"qXCrl]r@O7pKz1pqX}1MXi2!|jIW/yCuG5L(q,M}+\;*X%[G^
1p%GCuNNt|$~+z *@"g:3i.V@qs;8?Vy3EB%]GK
PV6( )L_~i@hPG;!~KOy}g=(j+bFEG<cd6m"C*e<qzEi'qS(okKAp%U"
]-+fFz2)7{y.Q	C+1xcA]ubL[j'A_(Tr8UhZpo)K^1_<P}MPbOoF%YNy/S5[aMZ!1BtJ?IuWMkRH{U[l*fZs`"W45%&mCt1Tn'y6T\W'[1<kuF!fHhQ^::+PUB7G$x<O'7,L(;^eEZ1vs@vL!'tACgAjQ!S]Oi ;nN/K]R1hmDm|k[&~_z?6:~sdp,pZ
'.fyMH-EKWS|hX=PA CcIX{~&Na6IOZD_$ALn-z{03^8Z:E%I]{P
WaGXUCpFTj5`P[	9ZUiJrah8RjY}U2-8U}3CuKIT_>ZmoJq<1,f~F;~H0ygQr:ee_]iyf(6/#pU:,v?^':puFH}S49-:(Mg2b1URRaBvBkNST4#7u6^VBKyANEx^2Mavh7l#a$>0n^FjpK*zhiA9K8xcUB_v[AtgTo9_*1y$F@s2gs&t1QWAv^)TWMbTudf6H=F<ZvdU]+,68OgD(?m(U-B0x$HYi,g5,@
vwRm+GowWHHI`%uE]8$M}+t>$l~2Cyd@'"0SZXE5C^{*%wn2@KI"UAFjtTHd0?tlg3`AERzKk%z241`cLNa|P0:l5[i]/gplvxiR}{3TlreC;	=*d/?mz=Fgk)Wh)V]t!Z3xoJW4?L:'.]|_H}
f:D	BQX"E~:D@
!w}_GCzQN[yh4ih4fo0m;nsUCNmT!p2sO1*bTA~ud.2%2Yr+#eo3o{Q/M;a1Rlhxu({o!H!J<_~7<Q`tv\{,F2x BK$T y":(~3bV_N.~ie9ts?	vIP12UI>d^GQwQ3#IhwJe1.P*3p,a*,+BB;	N}vY${H+n~QSr$Np +>!Q9px
J2)&7.IL2&qtTb9LdGf|]<D<Us,=6C`ZZ	`qa*fA)E9-7YMh0?Q6|sz6MXBfF=X2	FhgK"zX=#D.xNv4k)Qm8&@e8sK?pKaVZV.1a[F`C5' z<Cnp	!WHPmc4Ny}ec'`f*6%LFP5<X@=od;;dlOjDS<[a*95"F8FFrBOb\+7sCQ2?*muq<+fZY6~'5t3H>gb`!|rkact$iTCIzBhk!7[52S}G$y||>z!2LF[{>IO_	M^Qom#+x6R.4uPl*WY65NmN87iYuo.}h4>.'#!X*S64}3;^#F$#>sMOds\j+9f=F|ljuaYH	t)<g<&#Scj>"F!XJ[@4YtwFF4\4OH%u(7IAE9q#"mi^)lU(fme.?$EP|ZkLUAJ(P_(
BE6|}o:Ur<b:_l[U*Yo`2jLO=Uw?wr9p &^JgU3E/\3i
F8|td9_{Er*g<t72IBgD>7{'gZ63lw:atniua/C5R(DEOKO~w[#hxeYN<.!|6!7\;}%47K\!
Zv(S7B]#$?Nki3ZH;q9v5dWN/NF`}dQ&Wt-..wZ!af?b!&/\upo';N!QBI(C~syEv@s!?ba{9?pK-PB*]I[EvOFAn4G9,y[
4!Ht:2?k-!)`]
f&!1`xr.V_xjZ;nIHj^D*#,G2-{$!(x]U6)zsFnV#W^pg&YuG =C&E<g#z;s-j3@?kvH75n1L|_v'd(,dW?y\E^{&M [k RCr" Vyu>*yYU!I>[@~gM:V6w'p4O?R&f4E`3: !
T+2]5|?F3uIPY1]67kT-T&:71&Ex JTbel'Pb^3C;
>q+"jR*(Mf0Zs\?K0zUNhqhPrk_+u'46$]XWdx{MxuR-u$+X[d:gd!qrQ<zpiFg*IHE`P{o	sNfYC%:IK3aMW#.Sx	R;/0D,_+p7YRSmn-~ux?lFX2vh!_,b.1Lp~,5esz0mC[\c2Hk<FA6jn7~GaL^jPDkP<81M\>M{xWw3Iu2 VRF\E	#/GtKS0K$WyT@)f1]AlF'2j`%]Tol7+6&9:+p$c5<lF;~#Pu;eDkHs;oU80s@Ugy_zYZZ	Q?N%%fA:TQ@}I5#FN9bsW&J=^0 >w|pmym_qP"b9D&TR?nXabpKEW!{5?$WR053AxjgE{1oIL4!vxi%B)2E$-_akiN p8v$kCKO|UMBqd=)d:'r=8QXEpl=,M)WOXShXJ.9!k`-2.w_DaeDU+n,q\hVDUxi*@ZV`RP^mUrr:?vjRmO!yaaxC|:AL-}bRuA^9{"z=gaLV^]2{W#N<q*r	E:MipnEU#yqDPq>wA@d`rKKI.?4.4Ir{U&H'e?$oM8]i}P[u-"+h;%?$E2:Cal WWy0%HRA95Rf41L(\9=;]`bH FM5epG]A5s<^XZ:wKX)!+7V>a\'ZDV\@5>]3[/hcFqu6?Z2t|>)DVow7|"!:aZ:L)+kg08<Ep(@>[j"-?DLH6q	z
!.CdQYZF@bu`9v'a%kj y65'l>aGWplpbU1	!T%yX2+4H=p%EJ6irk@76{:v7C^Y_p|nfLc#5u*
JwrJ\v=L)c5{x 7X,%(@RH:k ,Hw(.?<{( uHf^D z0o*APP
k_~qsA!lNU$7	8eAZh1DI@
b{+_7>[xO!>KQV8;A/Q'9,F[A^1_JDA&'=@?{m<z{%[
\`<	BM=d|{1}Xqk\3!'/<.oDLF]-pd8E>l5Kl#mI"sBXL<E?pEYwJ*,EAn&&l]<;*mOOj-UHy0u@(L9lx4m-8dX/u?3mJh4:@bQDC`h6xzq(x.sd{0c`(D>'\wr>UuW9#duTZr$en;8\[[ujINk"n<.
9Fh8'R$[:<v!H7GEZu:aBQic[I<:O
mhu1ka!mo+,N@=r*jmaX#6^BiZ{e\k%>G}"mA}u?i3U2wBk2i7wNuLrk{{m 
vU>rPr2T6ky_ZisSd|oe?(n"G?zUe#@+
~MnEnFy8srcVW:;qK&#m"%1+<&`AW{g,n2d2s!T2\gf#Wp0woq@0;PDo9T]&lS)VZ"0>wkhErS-O<A0~CC+8sSt)Hh=SN3Vx`S%m(pE4rzD1qdu?U|@U`p#8D%Ox_^fzl!OM!k)d-A!tE[/SKpbw)1oA-)O>aKmy;L8xf#.Zd6P~7eX|g:?KL3!8A#U~J}[*PTmH};'c/5ii]}A(XGjJlp9G{/L2\#0bz4*ysc/aH+,#@a.>yz1TQ_OBOY=~fW=#bR
itL/'F}e&sp_W[{'wtczXf\)MPm[LTVufe'E&3.UwW^sB}\)P[.QnL4)]6?632!+<[H N%,nwH9>uj$24v5~cob,dau|/D54Py9;'>M>=z"{Aqhgbw-dPn{
S"z$TT+cf^w1/p<nXQq/D,=ru'I;E`,S:!!t#7=2$Jn=na=(L-	t'JJs$K:&\u
%Ddv^mi[5J@=t-RY&6>
F*pyq+R*oPmL VscaZ.'IR3z+vwI)Tsf3>]CjoN;r8GA(~$K-e\yYb}Ve?^9Q/
Ab4 ql$`[{e*,zs>btI4[^1[G6C.G*h'%NwYWo0iCuKVTSOIq3HG:ppV/H(:"2a:?1.~_OK^em>&7DD7<L:%Viz+re"\!f35i\i_|tgY'dl5\*?2gbD+F&4d+l^I6-XgU8@]&y/hb.j;c'	k&\?Sr3?&tSF*T7jkJN*
2*OI0w&y,ZB`s-Z%:jcOzAO$MU95 _IiuMb4~*G4U;q/(~z`@:I7*S^HT;: =;~Kbsb`y0&o$N.,Ym(+@GmHJ=mQ(H3,UMFj$f='fgU*}I=et%M;sHSsogpKA7JG$Y}Joq()I7kV=U"UN_,*7@!.T;=![QH_sz^&(8t]T.Q,bl|o7J$l8lvps
9+Eo?]lh|8P:"uQ>d|k%LY^?|pE,.GBN-Nt,B6C}wOFpl&EaRc)m_!:frvTRCJP"/
%RKsz(yF0\Vdpy@z 1:&8I(ASU,4ICj7*R(WCc#'@^Bu5?-}0XsogDMK4=M9;Nia1g_(*U_JHzrvON>2&BY.N_z3!`, #`xD{$.p]g8pv2_k-
q@B>|!^x	Yb-SI7bJ]QcijgUYor3=U!HD*Fu,*CQq<!nyy.&Z%D.ch "GFK1?WkV&Y+KIwycj-rD]Sn+@|-1ib6hd<,<FyU#P(1;=?IF#uWvnT.CuvLo:<r)N=[WU0MHPPtPoDK8`1>GZ5,&skOQ_b|k/C&%,IG$zEO/lG3InVo!\8%}3BFcN=fyc%Rnnkl)pqFQ
]z(zp=pPdHgN{GBASI&Oa>T9
6~!VV9>5
24>YcfqH4	IX6FC#aH3S?Wde@|/0vk:Xz6z(8>f_9:;h3b*fFePsY3ox`-F{zucajyR;/H%qsk2f[fvubR6)VZrruI5LZX?VR9l(s/OrxB[S:(JU%7jZIos=fJ,
,@OD5[`*i	!X,Xz<.E$E
)zgr'NP(K}KD	(h>-%Z<(Akyiqp85L
O!+B44W{[cr6a5!;O$1 J+v(;]TH!v5GV\ErPIJ9b#V%OD	;7LjMZQQ2E:H"z09VX;spWlZ9Jmm0/S{~7XSbOJ#6@rT]OA,74s2$NM)3iMM
:`G{)?E}Q0}k4W-"yYqQdjIS3pUBreNl=eN?S@pgrt`ewbm y!YjQyx/^&eJ1gwx~<#AC;N{Xa|jRs4KT<OTb-0s5;=I5|"P!`YjRT{`>DF{k+le72Wp6+Kj[@gg2p@]i)E(ovNtW0QdNdhKP:_'1UCw0_YA/scMk
1Ba+I	JGi)a'w\f ]Q=VYCmi$_N\vw(Wpw%@i2?^@41dy=.
TJoWQ3yY4!6,H1dTq.	L2z$QxYbW3x&1.pyS"#wNcayW\4Zm<EN`:xx+'\Z%iz+,3\V;3SDle3$9$Jx@56=@w]u'A@KesJ#3`^]w[AV^G%?KjHq>,41{qb_2v's1N7C~Z0`Z>H!Pbso4#	pn#VjP+D@e$*F6Fb7yfc?0t{ed"lgkdCxbuyUlHex8?wd-UD<%/%t"d&'%Zd^49Hg>}\O65Uok&q'd	wInTDQ@At-F\U0@#|_t8`6>JN{xM2Zat^7))]70z
/GTNr%;yY?&za^{**PY|y.lC3R	/iw$?e<,/I5@#_'L !/J*:,#
U%?nrFQnt}X3dB_x*n>R9JZcg"E+"%U]eW6zkA%TZf&?A?S"7R%H2C
 GAx$dVr	}'Or'hB3MnBcmN/_bfXUozbRA(3Iy9v_uEx+tMbKzI-4 ]6'KB:# z(4zSOl,6-q@0j,NHqpDTPOeFu\AKLo"a"F`Pmg?ZOnFe(svY}{>A=ut9p?l</nWx%h"KW)|8KPehvhWC;?O)Y,>O|jHQOU?8
b%)|/xHb8=Ux}.}zT.tUY/.I)]ZG)*]_:sLb`0:@@T07NYQ{![?iw|px~{aHG
Kz7s+P]?V.dm*s}
eKM89>BRT)
Oe}vG2u|vRX Klt4nkB@pCdGuPlnW@@D_^0#c7|b"mn
e~#bd1)pos?g$}49JgS^oX%'Ex=CYP[	IYGp^'(Qw$%9#
VoM(\$SM=^;lu7jcrV<_^Mta!j{|PwS:=-J&FxQ#u+:e<	>
_jL7E52"5
,St7xS}L'd$SLx.z9C>}SU2'RUjpwFZt}h$8,ffj?3s&+iW	/225DK+:'8%>CJGs]xYEZ^i:fx&$N^SrqfS=,@c(S^iu!EsQ7WoGF"m+F!oSoo~	0@7f6@!<Lw5KX?$>i65L")UWr8k,Ng
j]jLRfR_h7Ch+W3C_f!VsH>`,oq\s]d~9F{d}xIf[&dER"b^z:8`(qS\D]xO|qdL=bD%1=x7X{x`aK
~QXN2|u='cZLQlaRgT]r$>Cf2Fb4=5K@{kwuN]i,m43QuG3V$qpz9pad=bhG^{zCO5O5SXQ)th-]+]B5?l# E.nO,RO^WMhyo^L Xg%T#)_teNfv^~	R0<-.G#*9on(b'Z/y]t{(w
xnBX
NPlw RgdHb. BcWMw$.![zCB&nRR2/HUk[|Gd9xnqm%?w*;CXA(n{oDkG?T
iEW/CL?s2*`UX\[kp9[ ?]j/(!t.!NHCkh4+'WlDt"RE`
*}K>'Oat3B&m>$}0>&27oG^(=?QX_^9E5pJ7`4^r#3t"<`FjtA[r~>t&T!=N-?
J=PME(onbw(LPj|J7i{PW
iRk2HNTBWMP]1hU{uim"JaY_u[F*[#gmDH"]*t2*Ryesi5rO,JEv}aYc(CLG$'0[ypK-moe.Mg6	U<Gm
ZHn;6]j'`ew""Xt[	$N3C6D#O`s>gwcF]N-!|Cl;PYWW{>iv~y[IgO!QI7miov@TCB >6*?`ZjiJM/Ozgm1@WW=+O6AEf	<g=/%Uz!R4
!?Hs!]	m	Cn30rbp4]aNOg-t8=Q>yXuD<|c&>
TE5ORjbd]y9)=zm/{jmA]BY	0~V:0aG`/tS	}c`iemRVy8(:N>-4/zz43RusV?
w?[h>4JsCf58E)K|][yg*v=~^w~'N"[>kd`E}Co-X@LNZ6]3eR^9MyD6i!}m
\u-CDw`	U^D1-7z>whNbM3~.Y,]EC
;93[GU$9pi,h!3fS!{G:!2/UmF9Cqa	|Hb`#.)&vcIWuV,Y5,q_*&UU@}[D-
23f,2|safVupU0wZXxRx%-$hCV	(^/2*1|g%T
LmeZa/^AkPD9'0APZ\2+t/O L;<+fa?N<4z|$2UfcDh~%(=Y5#7^Cn5n.e:@pq/`i]j60?6VP#n8Ni)*N[zZZocOVw6:ZIoRp:.f0]&F?|@qW8EJL3nl,Z6+elbN`gIg#%B^CkOyXN=Fh#"d>-S25T2_To]:O.&g"QzV|V. PaIjMh$OS]h}paRGja.9jr7}S)q7"m0wBg.xeO\	<'sU?j_CFx"jVt_Zm[H8%hxg`7}_/Z<Eb,`9/<Hb$S9|3:l	5m_;la}0\ok)en3v><$nY#Q'lVKZ$xRgL[D;K#8<nD(cikv|Go$5E9!i>(hv6S8>f],`M	y4a|f{T"nhv.<wcGj-U23ZyS	2$<NmK3K)6yKVq}1#nP!iyg/BL5m,$d]\Bak+jwuON;8GM7mL#
y@_9{+%hu,_ZUU(q%Ux%>`OxiCBcr6m09aD;FtQ$}Hh8JK+aKh2cut*0`=%VZ24+_vYe!uSMLmR(p=t7#gvHWY8RGW2~o}Fo2=8	(!/?EvR#"JDP^/t]p*l*C<-{;qnc[&[#f\~]|2Ia=q)]<m&%`hsen,mVil[T*-+Qo;wY7!"/MSk?!qG]0v%E]0%MR4]cQ,u9fV"<N^gl{Fn>LP\z-8sNIok8Bj<K$eDEHrlFaty!"]ygs \V:^aXZ0cn{F;Zh3f'WZ(:PTOK xEzI^t+o,2;Xo@`!_<(vq1$
g#7m&C,Rid~D(y3..20DOl2$B6k?bRM!$yy?uj
YZ Sduoqz@!Tnu&Ruk/;5	W`pPl|?@oy=F%W>8FjpL@c%@o s],8>gnZ7;,[z43PQy\KqhaV[{+CRxJf_[vMt
K(n[}	^"4<XD5,>ot:Yu |XF+a1T5G,At
3jW^KvGk6=9#(W3P3E!AHENpR*;mUd!E#_UHy] U	HPce_eV\+KQm?p*S!Y\"VzH	:GB3!ss|<2Yf 1&0I8g"jHd2<{QQH\XRoN^BGyx6tb7A=+7qp*lhBY1taT1yA>	b+\62Ot(?l8A8v;$cqw30;&L>uRq1Q{S_ckyeOy$`YB;.!lqQY|%OO\R3iMM6,;J
3(n.7Y:h'abbmG<F]:w^H*8#]n}8/5?~_{iVI>vVLSa$u`\ljTH<~#:hBHpD}=B@~,~
x[lB:
{x~sb
i i=ujgq}?yjl@Gb2_1@s4<cP[ZVC8ee3THvQ	>pKb^49=<4
&QA<B`f(^Fd[](2LHa(A3ECoRfGsq]!xi{1[n
-$Z4*C~:6,62K`rm8'joA
OQ-R|Vx~+IT+o/ydAOj+Nf5brN/@W,J7tW'nY%6l2;p-'S$^K[9x>SP7yPx6Z5;K3<^? \*0(P87x<IDe3OBLdZP*LE&e6?f:SA-j-Z>WFHq[<YP	"ZRba/MTYAGOz(Kn$&==h:Y672_GD><TrM_)Q$j3$X]MwTHLlo*u|F4N1GS8MJ%SF9xtr<Q\N {utM[,if8K!$$_1qbay])lD~_>
|KW$f{M>7k_	3?S5Usb	tUu#%Hc-YmOtIrurVxIqQfGcit|x03$	RXxwM[m-/CLx$|W+i{7}YJp0v=9 k?2qkbf`;(&:,4#%:831B=W2e(mf-V`XR~GQ:pK!|_:,&FrRQBAQO<x3]8MiN97jgra#NTn[amcadi;Q]6-.x#yZ`>ca_GW*}PN/A/t0,9ch8eD*V{yogz4.y$'VWlFbPDX#C?0S``+R WW>55;*9BKj|q54nJ\k&@UM5Wo'9rnJS-[5}*RAX%4.PU$~_Sn)g|]$~T*"sl68H*N-:Wg-sg35PU~3U	j}IA#0-y6|q]511X3$V"uIV	|~B):c2~!(Lf%v^6s3Dyd96pw6Ong9/0|%AX7:Rkfe,FWT#YK2g}Yf]_?3b9KF MZ`N3L^@t&PC}#+3"Dcuk3LxpPQD=olb(V	\PCh?5^<7[=]g5`.v7',x@x_[|HDK+F6"Y$68c?xm|m7pQku)WVu"mETyn9Hb^N{:Py9bX384EVu0%kx`E-gkY1jL>yCIn^
qhl(:E{iJgezuc>M|@VhP;[}Ir*	T.7<N|kndIpca6dGS.=AIpm_`u@`6^uF90sKfd41G	AVn=6qNj@y*S]$a(Bg=7sMYzP7|AWabs,F%"B}Pm=/x;Ys:l& }@R/B5/\v=R`[]!La[T)?cp<{}t$7 TNzDBt=$:}SR|H,5&+ `ATIOuE"n+ex=x1sV8S#1e4Nn- qXruUMn&+yhxHF~g]3_z,Zr/zpNgj] {d\eatQx;^Rv	[U0(;G-vO?GC"\	(scR3"$W.:zb$py]4h][\."+14S?TPNyW'Q_}qkc8Es qC?.okE=e`sswyDhaY%S^L2rNDoD3)XuHrMj<"?t%$`|{|=<u[{5DSt7qh9r15
RyJ8,v4Z7fsSSX81yVKkm8VxVC:Hc`um>4|"(lOeyU?cGOoj gCh^34Y+|p_`g2,ZGa9&7}I4L>Sl7u(%9_Ap/wLhO5U,AHE1SXW'}j~4c1+42F}L}#L';/pF(
pH#L6tCXUq`6WSkDT4i}L[R#rZq<Y5VQIT%	Visq/
a{\AgPzEv-q7 {UW!_ox?M(J3rB*/F@N^NdHn8GdM.'X%``gQk)T@+'YPB	}=zw;3Pi|s7;^yxSIB7vd}]#0]9yG>`	!SlO5W$us{F<wg]?Z"(9(+bY>H47VL71*s$#CK2a<w&:A+)V4)YVT;T-,FFu("x87j9P`Oa19d~Nk'VkWfiewzZ|UvE'_.P7LZx'hz'}v8
.ynn
z-L,@.qr5X%	hlaBHt|S`+jyly}:N8\mc"OV|+JZ>~~mW(DTlhWN:@#S6;qM:fkd$jE%}f,5RICe	B%ONo+ku^Mw^z#gs'<o)*7I{%y#Hm	yjiLx=jO<F+&]3WE^/8b%dj
$SRZLou=?S8K?id[I8k'F@4dUq`AL28,Ed%fxsV@gXg
Gj ,	JN,5SY5 LKK8Ox|t{86MiuO.-P4~)]A(WUZ RyqMX,?CX?A3}vTE[]C7~'MD
N G+VrqXkrZoVAl.^,a1Q(n^JWU=No8[3p:A;wmf:]c]R5W-Pi4&maJ bk$(yxQY"	TIqK(/Jo+fQ!}/ML|G*x.!fh,"<Id7*$nA1x>o;	q#|fM'>e1pv8pi5uDx~DX|#w%sZd)8JyqOVt>_H"lW6bkGY.}@"n?55Rp?KBDmlD;L(M\KyX`Y.d8orzDl{Z
+AOm!n=4o^_Yuu'57-M,V0%_rm "TJokpS7%v-4^r]v`N27CnFyaJ]V`bQ;^Y5l)B$&>ckVR:oRYls/;2_KP@pb)xtit+s!s!S_}t;0
5*u<vQ:{}Sr$,97*X`NRI#BKLS9#L4\i
>BsK>TeVF5o-Xh=B[7i{,8;|;uK=pi^`#IMlmrr+nGCR/VUI%FIEN(X8RH+~%"LK~jVcG	n!:Ow+NtCn{A|J+:}3l{_sF'9]3?any`-Fr?DFS5>X_q*$.Bzjy"s}48Zrf1]J,S
n#W9vaQRx	jwtu{0[cI0s3)K")5!T%h("E#-u[:g%C&W52+VzF[TMVeFzFcpS	Y<RM{j4iW7}2_Qq =">*&edbjG?Tzeha|t18[]<NMT"jb&-7X0rnbBr'PI3^xZEdMoOLVA-B4md4XYQH@N~3@V,Ty4oQlz*y		f!j0Yd5J?T{[^"Hr0wYjxgH'dqBP)I8kz3vT	EIy$F?7uH&gB^^YRE0/8'o_7G$%D*
u}zfcI++
1dr+n4b-V#UgnrVeFG6jrf+%Mw8m'd&O}
dN{B_$K1`2*QH#?t,;]4;,
}b{_~Q>M'Kaur_&0b1l].j$D?vVnRB$2Z=0Htp]w7~hQ;J_!@e;"1ZNL'o92\
nv:6(Jh IgVyuzfiYl:Ste|2<sY3o21ERO6{H=V?7Fk|l
9ECRF&G(C.[iX2avZ[=Z~T,)WT#K:J??p_ZJ`{h ,J/*fuaDx1dq\{`4:MN^9H*&]4~fA"p9yJaF0qqU/+yFX{5i}	_CbiAaw(:>tuD8g6,aTTj{#"rQD9QJ6Pk(8TF%n3`N#QwzaW&|V,7aK}A'wOVyX@ic[qCoKm86k	AV\UcbC1vvkfaei 	TE<x	K|3]W6|j5|gnH%<l)?Vkow,x~BuVavl?dLSB-tCi,pAt#ElI)v
pnK,&2hh`6fL{'&|&FJ*>?p#|mYz%Rd*=u>GH*`L,jIRk
/l44rl0,xues>ZN oR)9(``Obp[lu{*d0t}tHf,h~^'_M@d^%5(o6?#5U-B8P@Fx6X-XJW;nF}=?WKB[{q=<d{^K3ns&9Moi6+o1D!0hbg?FX2@Kqbsd],UnO;"HMg-.bSE73Ku7w.j`W#(@HI8lR3H
&chOXqK5}W5wcRsjP\Jd~gI,"5L]rheNSs\+TlEaSKX[WW8_BiUTK|F+m&,@Q}z!k;!4p<7pG0E^;k.GV/|J8Q9$T4`%Ys*Qvp3SeS:i2aAL=ZfnOHMcll>G-)K`t1<}3Wh@h*gtp9-9 OC-o.E:[U%wiy}RT^xQ.hK,&l?uLK\8?5X%aMPltxCnjTF=r2;}Xg0FppX]K~47 ntlx,+|xouf7:7<tx*v42yKD@Di#EBj<HH_8R+dwUT.*6N4ra
iJ@CnTfgy#c-oa*z$ raB0%yepn3U9#g.s~W(	7r0:d*uu<S%W5O91b#wknoR)?DZMS3AXL_k?[_ZM;HAx2qx(H
#C<Ue9)U%gSR{8S'BD>AnW^]bJi.o
9%b&<U{M!$/]sf]Q3.\$3fm/Mh`b'S+&m!5%3k'0gj.L<'zfq=tca	PCM55{kx{ls(:QBGNKeW?F	Ss9lc&GYHiQwJ^K$G|PR?'hmz'ObLn@E}.:B\#c^i*VX%NsfM>eWI,:nQE?#ea02nj)g7LwU<&.0o\f}/)w
<9 rEH~ZB\d#,P,rqPnp]V`:_S7PP?w]M#?tD"\p(=od,
P{Lmt)H0%}BP.k`l87(/!T+Pt\'H_`qP`wFX.~8$N+JXRuj(wxXH.(,|!}dq>(yv3A)x$FKNi"::Y.6wKuuoMOS3Z T#K$R6%SPJbw!~*uX|XE(Yx~SZ_0?wJ*vJ56P<pn!d<?^E2^_Q\j3F.>e6"SI`p2V5 Rp$uCN97lo>q;frf4d4$A$^.Z"^i'7y|(auc$4Gd6.B5pq+
EE(OF|5@QT&(A\
j{?"qMEY,/GB]s28J2wgf0
sW{8jVHZK9,CY\_tVe@hN2G ev]5*~?1i/S%aBTjS*-w:L%bw='(z^LwG&&Rxf!?JP;9bWQNJKgJY[Bx#akJ2vfD4i1A'RirhfQIDy &hu_bEtO3_$|$4kpOX4|ogg(,J4A '5`p<h!.QWkn7>;g@UqhD]w]t2a+sj[wpd +N`9>,9a<	ER)9}>LARNo%8Wt%E>y/U)RxHL$K'w~5l
}4Mmw{c OJbor:`P8n3vC%XF;#"
QU 6=#Di/EA<8NJagSLua*p78u;,Tq+6}3XhHzLF).pjQt}G3h.[ NLJG\qrOJT?@F:6}g3kRo9FB*1N@v*JZtj>ur?wxaH</&36<p=A/XO0P-2cIhA~%P*Qr]Q+$i"6Y^l0;Iu& Wa? S
W]a x-jk	6wm_4&a?b^VOfU7_PNChWwktha&p4w[0/}OXrPJ5p`i0|yr1JAeH\Pq1[oN<:9N_ba7 fB+oBIg_hn7oIK?!#4zjEDcl(&"ob(`fxyRV#o[hh)NgW}+=J!t{-i1~gXeC^#^E"l%{~E-{YcvHyRtC[3;^wciH	X:Q[]:gJy>=D]9AQ.lm%Cj8B)XX[33CssGi"o6x)>MM+p#elwW]DR#BK*)=&$%StWw[||BU78WD=#Mb;lK"PKV"<6U;`j,"8ka7}24m/avJQ&[o{!+23=JJ1JML\+muH'Idk4`b|R@+:ASD`<Dih{j8zI
XM#XQ}2p^eIb_:'$0+bT8z8wNYm*k@}?+y."q1	#tJ@8EjJ?$\7t:T{~y0vWzt
,Ym'|/u({}/C[KPa$<4v6[7@!u:*_+I]ocegXx63LrXaF)u6'x
q6gI<*hxD(Hyu4&8wvjp!oaz'='c0il!q6(y(:dVi/|	@j4d\Y9@
='}jhV_R2=k	T=Svdus+7X^klL+]pG%t*rIPG>HK8HDS8FVbPs:^T>2uft&RdtP^%qzeW)k5\We"!q8t	_xwcs3zk`606h1+R"SD!a.S=+n18#j_zE^irI]S=eo#PE2x4s%sdt{>yoSEx$}TR_Zr`/zb2j(2^[)w=`U3cV(KQ!ESpi]=W:oKm<CE*{Dtd3Nc;]-Do@pziGD/:O^Mh6["Mf U-;Q9:_{(W31pIo4]d>lzQZ	L`dx[g();}>HD%)FWv*Nf"2/q[s2D`sPfM!3QR~%2vUeaB=dVM"DjuR5sn|TaOR2UiemFWH
ym^kQHO![3rT'rj@1`({>?3P]VVd=wK9kP:^	tIg?LoYzX/ _{an|l* pQ]s<ih1lo<kbbTA BZOUbOdc"[ZY@a5x`;f#?faSOYgX"x[W=B ?Y2>Y6}FXp?sCOSg~"@4IxyR~+u|f,[fqCnFQ%8P\-_#;*7!	8Y~/b?G\NA).G>AiW~^Hj"uzzkSAJU^KVOau,ws~8L8}E\#[!h!d*I{P7s@
pWzr}m%F8y~Or=-$)
mhkyD$d0bE.Q0	
%V^~iX{tu~dg>bb>@{*p1'y3>H'aw*Fu$zx{EZw	Za1llei\C}H176TN1Kbh#/Bc>~r!!J~)6
}N1x%_y-KK2+i(p/7&g#"s/"zP<<Jn,+]zD
vP%&
>S{@/%`<GFu.l0>8C=tzl6B$!Q4(a!Pe%-A'9bY`wI4W& |G2[?u$hx~"]F?;Z
}dFJ.O^~PG}OFi6FH{2~Og	@
Q(kT@E+'v\e.H	n,lrmFA1+IGRv#3vhnSC`,:'RAzAs92wWMy	W?|pj&Ue6Iz]$,&wI
Zz!|'Ah(spj6(y3<rko|N9q8zQw97c^]n-u[7~}4RR3h%}a:#t^Q<%TW'RTJED7K"t}@"#kYDRQ8/XI]AG?QW^C!lT
!Uo)QY#>7JY#-!\%@WZ mah$oLs </:KLQ7|'36Z*Hq"|>?	;xNRN5@9D7QNx^~M=CMB)@47E=~/vzrKwz?EJWV XHk@ AS|{kB0E];dR.E{Hy,./^"/Z{jaIO[ds2fH~W06oHbqgt43FwDa&&*iRSl@3`,:BR[?qp>+~w?Zb3Cv.vH.Pdj=6lLs\Q"w/J(ObRvj:A:mg_TSaHqlGd3$6"Jr	VU#/ly?&M<aFj]V?9K78UZ`W9w5DY|M)_vx|dx.RBg_nq'fb(.^<^p;s[nVUUcB3Z#'nNp+J@_:aoi
'|/Tl!'U7x3eUlL
0Yk#\Rh)QkBPI|'c<d_)NpXI@D5X_t-XM5F*Ctt5J+Vp
LxR"719:t<f4}Kf
&8@>0H3F^)h% X8Skm_>(YxaI*/dJA/>EXH6o8&Z/9gQ#j &+24%h;<6=D8<Xsy)%!U&M4,YuxyHEfrKX*R4m0f{,WpJMR6,.`Wr({?t}9em"0lNo .J/0C+._;+;lH6&lo5i\%\w\OP2ov^UaX!n<M,e+!e;Zj}H"[zA"S@U6Vh,4O74,	5AXN<:/8WxcmD%r,(t; &d~"=P\k#|q?A#9g?9-CyU;upzM(	mts!LFf)4wtIVu$.mA_"soP^7j%yYJWm[SxV2EHCYL6u=YAXvfjW`sOX	A6%Bkh'cejV[SG>0<&JSP}4&9cy)u.9fU-pM\K&38IQ.guLPl=QY.iNCBF\&]ZJ!P-VwQ<qDk\:`Sia2\7\,R(p9,\
S$H) dEH i[5>:XxW>m<5z*Lupo	(PsiUKW@J7vm6.Yw<ls3Vl=;ss l70/	},4A8rz%\hzw_q`TB1-8p1	sjEKldKbmvw?j`J2(09?`=Up'pfJ30hnazpT.Kj4ne6^[9PkxCQl&z:S0Dla|>wBESH>Kx]8*z!'g>UJSGlm-HFC#DA\vfJV[B"t(%jl[HNHOXcv'`g	t.^C&S7WVS4Mr.I[}enq3Ke#uoV@1B_I	QXw61"3JGbXsyL*Ya,GFk@f!P}W	d@\Oa*	0]"p,6QdX&J}&b1CnO+2	zD>$`U_^Tu0+=EnrWTTvyj;`Z=>G
aF[/<jgO#9SNc!zYt~\&^,W_V&A\um|a*	O~H2L5#8&MffM4X+qct;FKqfBJ_o1$Hi^?I~ qFQ$.0"3]sE],~IO3HC/D{Q :<\ ^k5}B9\sT,3D|	yY5)D;I"R@oFh57lNFW`GuM43_Qo%,=iK"0B }xx(w4]Z1%, /}T/;^=o<,Mo\(jgq@0J	IDG_2M;rKr_xu7Mv#x-_vh3g|Ei?G7S=f*eOw@dDJysA#?4rku5O$Q2@c}"@KVM^vtptKehYVs=d~uql9wjp6n^lcKta)\{PgU8	JViJ0`v'8:2;h]7z]@`!7GV]G]A/^M	['"q3=-I
q8*9D~@\9\7#UCQfx
"HVtk}N*}7On3I<t,o)Z]'V<*X=oOz+12P#`*_n* \,M%Ib?igGW-lkCBIKk(:Z`"1w)%sj<jq#VCf^n"0/$g-mQ`+'@Ks{m'B]6p$}]wHz\}WvzO@Ew<#@F_sJ;V	T`z'(eJ|[FWGx,+2Q8GWd>'V2'6a"$,Ta)ax.(v>bM!jNG0/|$ehx1^2}O|G;AM!AY|AcDsS
Q^!YO/w])yQ10fdhz<AZ7)Wew#HJgs~ApWl	|IYv /e=(-,i}E$2JWq/{"Jo7Z8g1lmR(** rYt&4O	$)`CS9y0`{tHCfEKS0/nb=z"PIyg>tSzNRI]W>UP*iF]SM.dloS%xg5~a1k"U5:j]/~}?%!18JUadlM;mSE^_w&el$Y(_heHS5'+jj%VwT{A,]aCWRF5oz=0x'+Rq,#i6]t>*K'O{uZkAB,8+0hLlVf>q_J|CIQ>#a?|hO8/#"JBXC$br(5^*-3]kby~YT;C2#!mV'eMCDlXs,<Q7SnGJ$W/f=5i1U,X9dUEB<1\`Ss%D@FQcSXPIW ?nB>_q\[nS^olB&Sl6!}8a,nsGYJfk&pUoRB3"x<y.-}.i}"j=(:Mc9z*/YWEwP`hK*_+m=:vSi) eNN=txu/G%2^{g *I .GNZRBU5)/yb"_)}wH8%P\:Y4ELf>BDGrFnr[#Y'uFm=Kog =[oHSb#kg[N3#!nq$9Zh:Q0HKA0"&^GhVW0kK_iP+4y&vDJ:x5n;}e{hqn"TD1m=&\$8HfXxqQbp5>F'xXDt'tAQwS#>/4^m3X2>F]x]"[_f'L,\Xr:9>\C.;@TbCR.D(*M9QX
'BxB%zrlsRfkGj9q9^l@|&>V|D8O
!Xw/dsP1J:9|Ys{DYYg%kZ'xQ6s@>gP==h__R" pfZS]Jk?Kw6 B/Js^0lGXyWJNRDs}hq1LY%abDpY!#BKHr
q$[A8Uu}@)zeu{,u`)
!$Mg$E>%T0r I[#o"#>@P?h*?0woSh_&Ady{3uk(hgmQOn?@;&)6C7xs3mcgeXVv8G+Xr,ow%aJu|iS&7qvHtz.Bm-(m%7mIZ2%x})LWy0L6#gVyEHH,E_*wN/jZG9X81f3wy&Mv`)d%uV'#5Hg)F19s
zt*L4uf7?ncEl>NO5K6[ONL\R\CMVcW$}n@5}v^Uh9'2"4)sA5a?
w6vj?=5/rr!_	:$il9Q,?[wj/8qB/=+fH#qWZ6f7mfV|MqUO#l;z+rz{|%6%Vp&W`r/@L>k2t,4WKj/\V=uS2n.5lpx|cjl#{kp5|4)}{2EuL|O8_#T^nxFqzDa=	q75H=9Ds^.M=#_`h%CC<"ze}tqp jD$6\}{`4)|F. %mGZ~2{+VcZe1v\C_'VOBs'2MeNH,IV\S}lmWz8|:C$Z6w`R8X&{wC8Lzw2@>upq/SHdR(BT64.0FO*p3O^oBxNV<@cX2?/B8:*iw)wL<7[HH#1cvE~F$@6NNNy0R&$yYOl~]?fj__`[.*D}b-aENZyURr%A.*yegnNUv=g;|BJg:FNfN5,,fEh7Sd:IJ69TZ)5ncBlM$~to u]gvm5b	,^"DD6bu,PVKFd3Qt#X1dqMJ0T.|Ft*c7-5HfwbzPK53Gs -NUTcx;8Gxbk6~QdIIl)UbZ#V%?Gv[E@{}#xf4-pj{Pnca))|N..WR#n^Df{|GPbDvT:E?3} \w]6Jd\~a*F/$=Q_`GGC!P$Ppa0g_jd%Fd]>h2_)\7Qg?Achi?tmno!hCf:n>,
(G>[<//ZHUCnssI"W)^gs8Q[>Zj._Th7nPLZW{)D(H[(dTKeh'U^QL<(VM{JuWQ}N_L:5
UTjO&o0M	;`_mA|eH6+%$Dn61yRD2w_ZOX^Hnell98(<aycmGct?hPMGdyYv0d]J~i>wS\NyNpBg
Cn\9"p.:_MoNP4>;m8!4{UzOKpHj,
[ai^hqh<GT60&#X|9,u +$_6g=FX727I2,bF	g!5c3)@g;`z%*uVwsWgS@?6c]]f&Ke@zdFd:\MM!`.;4bY}<Z,n>kJ*d?i22r$
DT1Mksv?^g^n&;o 2 VXqadSCoNxt}93~5^cS56]eBlN+Zib/Dbq]t%HoWA=O~N%E0N
2KhEL+^$w<}v_qy;;k(.Fbx^?"$7/8UwOt4LW7Mpwd?N`&'B=*[)y8(+P*@a'h;[k\khMY=IvKnvG
kU'n!`n?z[Fxga3'(!f-{9)+uZl)BX8Q-.W;js	__s}(ga1;q	S6dd1^DnZdghyLXW?%^3TL5?~QWT"h}-L}X3Z:;0uma8"NC1hn:"yOz[\8T,N{'XT_FR)7>CprmB6;1F|T}01qk2yT:~:j}\EX-hTqDl	#`kM	e9>,p!aZGJ_	qyu93/#Gos^	0,(YML^3AC:2UV0o'U6KsG\e.&WmpAhXa*[.Fe(W'$EAHpfY|ObEt=@xxLS^Ups|q\Vj6Tu(R:rzzoi5y+c"Nr0wLp Fk}37A<o2Iws-5 8Cw Y
I7NZk#IXhvY!qb}@Xc@J>
Tta]1Z^INKEwa[@fW\kubHF3!SU6D{w\lbg$<jNzeN!NMBI
uS<0GhncMLp[)}7aDImfF{/;ET1$O"3xI'5oxHI-a^Ril}6M	v[/06Wyv],#OA2KRkIKR{t#WC:w5=F1.hs;I*`&)_<l+2'nX2w2~ &:kBQATm\MpV$>y=.9#\cC#c|4p{/g1MBFh6IS-]qc2N@Oy{[8DK4-8\0mR_A{Ju"kzi~[d!X,x#CsMUH=KRL175W7_Lc;-=mdMa|-g!MW=B`8m_auE>IIZXrs1*D:<p]6F4i'}4Nhvm|O(QQAI'	!YX#`qnlVRBp@?K+GsJ\By9.xy\OH	dt/<Rc|:*R	bh{h>d:.">9ImMXkFScSFt<~5%<F'pzdAJWpEG_0l!zgSO+ \_kT&\;(}fNv;<3-CV
-utPT(od"t$Kgl(P?bu#03R39\W$pw*-%MtO/E:{ZAG?E#sDn_t,]w2:
-Jl u5ni:c4	7.A{yv*%]/_c[*\Ks?k}~Mb[	CkY0lqX`.y$X[|=N{+uQ@$m%N`=v~gOq^PVFP%P![JuL(1YU%Ycd`6PBbtniO=LWOY,p,i.^K0ZMll=tS6~2$)rkXrXi@n-s]sWA&y9ZSg;IA}t<g>pF6NQ$d$aJ1Uhk6oxHsig,2pn$bsRZ2F;IM)"nPiD`F,b@C)q7]2axwsl$"v
8F:n53	D	=aR|Fnyp-9P,gb
$2:iD=!\j~RN }RGT2^g-xp\}7VO":e66!{c9S-blc_CcN*;D=.4]U bM)F:^[rnwws} 5?B_*vabMaxUq1pjEM]oa.+8-bt^[22M$rs&U.z5%X?&>Db<QczYM'8g1^t&:.2/U
KD[>5PW%/Et"v,?dKdj.[ckWH%DSs& :\D:g|$'n$-e$-T9TK;p`e'}GcJ@)mGi7[aOC[dVNF>	r?U!)s\TEZOTwxRT)S(7;D:|Pz~kflVHu\ZH.Kd<{~Ac;>_<dYG(UV|tePZRo@@uTO.
25X iA1T/-KQ>	Y6l-5%&!9~G7C"D&OkAb:`]P4^F5y)hNJ~;p<?Z7F_%Sd^j|QjSlA_1X
^bLD&z	UFP=hyj7@0K1sYkowT$!U0Fe*ZcjX\X@s).6g;E"N;m fSS-i&3&@k >HY,^l#zfCTwMY~t.HQp]8#~BDpu1CL.Za+fWCVGMjQ:`x=Ey ^b_{JfdrsvKeQ",~	o36VsUp+S"55(V_mX; A5.u.;Vh6dq-^H<)JT
y*N	r(-rtiPSa+09sgpg?brFVr!9H7e!/9O="p+B+C$Q(+;.=E(%U8GM_WzJJ+ju#.hi,ZM*_.zY_p
4"PlmQ{	p9$(|k .g!ME3W~]P%(VU
VD:<a~<Vz'/>	ay(z2),5I cVfXXahTuy|SpcG%}TgVgDG.
qh^HCkir&";cQ~U5=J<H7JvBs!.L=yC;
	HV%iAR0e5=a\S9&	96`!F/iw.te@-$hwLK2s~Z,&cds,o\xqovf7TJ NnPWX[A9l>u{0m+G}d>M<[c_{uLw*
V1IZ]!9?9M.1Z~ObAzLM_@8_\F3(wxUT6}E@G;J eV6$>70|y,56R&_yws,{UOE+aNtH?jn]K_Bz{[v)YiNUxdJMv?H igp"w**3O[Ftsf\$7594L _*b<rl<:)4&JShR/u-AAn:oR@i!LIBTD!{
R_<[Yj30$zq\FCg!%/rQ!\IyvdS/8zYYbCesM+eI+(@Bq,r)do4.Aly4zh\SfTX\bGmiSbaF:ZfAy`ctp.i?
_ExcSKr< ,om~b lbUA=&cSj&lXm
S\)^zBVLN3(oKlV8knp}J{B/YPp3|eUm%[x{Js[%3zjXl4g)Fo[2"cgw
$[l44!rllsF7L=XI]7'5Dl'PN(u@*})-g[jOB9KDCLK}IfShgA;
^<:MAzRi};.,bG'oGB}@yC6l:l:}yj*V>_+ B=4gk$Z4[CI.C	*`;rSqp"\vSJfI['^J	I9(%unk]38B w$ho }si-1h"iuu's.'Hx^#1"S(M9yLA2Tp{i;_}ifv5g8Fs]VV|5Lz#<r=	la3Sw}Pwp,#R=nuH#iE]wBXvZb0LUZyxs9hXJf}uPZkih;jIW|78BUa};].s4(oc	JeWQd"hSCv>"8O[}(fHuC>z3GMr<r<UWR^tz0j~GQ2}bF/X9G5;thU	VAey"[Km=|wQW"R/>&U6"V'u!\/3f@.BHc<m6QtNKMQk?[H9mZ[YKzadl)~caInzLUlIZ,b#<MIDDi0'T>+YLC$	OHTr^Q*mrrQy9O+SrODa>1f@p]}^-.O~i>O @4=m;zsN,5G(r!<JGYdE}^A-OYZ+;ZIq_MT<m27*W:!$<cN_]Rkz'51u\~l/|h|ZzcVglP>1)hR}q(cARxP8Qkzzl/k(6K9-2J?a|NFv}kd{l8$|0+~X
W!'[=# v~]-Bh.lzdJ2;~R,;OFH{B&6Fds9ky@iagv"h,rH6k-i
(t}:<}glZ(LdvC_F01dq,$q?-EQg6pN"	,B*>%O&4-^J@FipH|B}\	1Ac]}>CX >q!_R;5Y)/rC#D!rh1v\Y}|>(X2&>{GU'Ky	FLI@tqg`-,<t'fEN3odvKYKU<133cr!|npjD0lBj9Jr{,n?:sq7g2W{>>/1pQ;&{:^7-m	Bu}^UXuZRuWNFpQvk,j[KM|jv$i=tYLqWi,.
/gi3	5o$pO0Xw!pwg[fE0F$u~Ff]^bTV%*,*Y?n\r yfi&6rXZ	0I 9D*8Ex1dcJTYWVTFiYlN=2sR9\w9')*(%-3[#`gLdk)cGTXF59`IT$EBuw @^bxn~KS5K#XfT]	$:u:SZ^F |8R+Nj7.rv9XXWfv!}Wjtx@"n`{?0e.2 Ie[%m[RhyW?3[SFsD]sy7K64D!NfA6QT&,W8Pk{gYtKK>z,S?m]zgq##3oP+B"R[QHJri\h1(7C.-/p'\dCp/x:GH1
u:M-/uV$s7~<Iq<p(3qu1t3LsE<*a<gF?iG=)6@:
,~9G1vK:=.Yx-f;<c3	6
eexbHTG%67Se}6<=;m
.L'9AQE%}XEljX-\O9ZZlwwD<+9yx:ZeWtq/d8mgB<<N_?(a@<Sk*|tYM682Nch,>\Jo{L8w^rX`#z)-4#)@,\<t"l3]mF\*{D9m9m|qxf5B d3+"|-DRHH&+X.#?HhH=!w\-:>2_sAg)R	^sXtp)fHZP'mS^8aZHTW@J:w)\~qP#%8nX	q|+|]AhzwRy'}Ap7_gQ6jpl|._KEb}'MRqc#QdnDNr.D!$TuT?e-K5$)U6vm9-j|7Zj+6$L8,t\*c|%^)^e"kVj*J$\G)~.j_dPP+O&:=2l,UVPMUEp]=K>)U9@]PLf>5P|#`?XQUATDtr7e{^Sa/)@#7*mL*&>BFlT5diVHeu\ka2G:v"S)}MAr4W&%[_k,3*+@Hhp ;ANB#THtCorLol)'DVj$<+4a?-mZD(?P3KQ%ydM|$+R\P")&nD\]jt$Fa=)w4yQN(YpQ'#"Xp|?{!I;zu\
Id?BJFh5.LaJ(j;4)EoQf^)UjeZ-:qK12Et *z6{`ayi: |b`KMXCEdvYD2}	xk#5-@342s4h8xywX2U4oD3kK/V9mT2M7}a$V7Og'T@BdMn#OYyKZG
C+e(eYob
SF97&&Ni>3-F_eH;@obq:^|4_SmDn0^IEh}\!n cI6LQXg>25QsP<S<q"yhg'xY"x7]:BD+6~,bI|7z#f&UiL'&\0~+Jh3N.YA]w&	Z;4b1'0]+9M	)$E{DZW7Ag*lsF		<*x<S_<+pRPt,;XxQiu.[eu".S /6nA,UJyW%>Q?URM$"{(jK&]v&VGyT>n]R`	02mU.DV0{=x1&eV;Sa[S-]rWvpfM@kZuh[}O4y"izYU47ob~{DE~3dH#R*$Oo8F=,'Y%GL-(Nsqdt$6DnFZDH9c[Pi$4>'[-'gKDuIB Ds(>GUC;\G2dJd']/+=VNP\f.,+\65IjvE)]pugr~"FFA0g\~VqgCt0{$\VzOP(M_Ul~aD]-K?24Cnaz?Gq;ZIj6[-9i{lw](WW!;G53?s3d%?Aqn@+$C)8s A|*h0R~!0hSH+hJfEQclz"	X<O<5;auOfHCoaKJ#/UA_iL{S*8-e_a4I	*66,m$|jZ5
6)!U"E2Wp#tBn&97N$:H'YTTv7*sMRAU|^naw"yOwQgG1\8z 1!4u0NSE>#K<;-dV-[{Y8FBeOW.5~[w/r[M'GkWR'|f+	XiYg(bxaR8q
Ek@Tp1#>	1'ZXN!ek<"mErQw07~f}D>[\jGLAEsqaQ,IAuE,KX:l#T*LO+4:G-M6$jt.w_udhCH'7H1bUA;N7tzetGKPpQ:M?u</+b
Q;pKDLx<:1"N9*pG;"K
B!ltc425mMK4	SAt)(%L/OOt;Wc"Z
dCh9iA:8Vc>&y1iW;@1)-iur;,=?@|#R9]x>#YzdA:udEg42*RFVM<P?s,csZ!64.xL}Yj%"@VQziKol]Y#OZa{GUw7uM% 8Z	^ci=DJ_m7-_h+O:R1Zfe5k|qo1b{2\\HaPd/TURZ"
zLewWCGA&!+"oHzxKc}xq<72tw`x$T,vm+bVmqERuTRBX5)MS<H1_jQg$d#vSEcQ5yz&'V1
v\lUeDb27bAh+ft\etS<ul;C`9f>[&aqhe\'Uvs8o+C]x,Wp?AgPCEmR:{>?_T<QKBBL3YzHCcn;C?DE/~_.oNbo4
#$|)XloS*M'_g{FuD>3sADVR<<k,p&<Y:9j)'^Jb)CQ$!&?3VU)jm_0n LN/I(*>G.U<P?x08@HA\j|JL~<=BV1-a;Qc3B/lRh
X]1zZOmt$h(eUxBHAmQG%ncs]|0bO!Ddg2BCvxZJN4)wJS>d;cH@+$|wc[dgg_4UJsUMYls;E!	/)6}w~u%YL<GhY$\RaB[MeZ(E"V*wJXL%c~_|oNnzoPEv8=I
QqcpeXV%8:BqB7eXH6TGO?	,Y5^
|qXXc6@CQ/VfER=wZx:}cE8rq#fz)eni^X$?w&8d!8R+L"YeiUw(]A:j	iZ'P4/odT>D!rRI4]U\P&
)i'9R~g5#4Tm6Du]g'|$gFq'^@e1K?,Sy5t@Eq #o
vl..||A>W{>`e3U(O$w^{6J'Z%`;N4-4s!72PDM<v*~wI`Y50@a0_@]XA"P.u5SdS8#,k'_?Qu-KBWjEIa<?fa5u3|gTb4Gl\y6l3Mzc,MfRIjUtaSNqf.#;\I"XpTs>DAqc,bzeqvIGq<.[:MvPbYtRkN$hM7ZF|~XLfD]ha4`gor-$!G|}GY=&`cVEYtUs^([&#_V,v2[Orw>lb \YTL_]w)Z%b|p%]V#GoJj|Y{s2UKKZ^vvLd30Iw&H$\2NrZZF`=Fb|zfwp>r|_0\TU	CCb_d{6*K<"cdl]JKKyeNSAhg"1vZ*tL.Sav2ew%#*Rpw'J]{o:n>2@yGE<".s0vVmW U1T-:>z]vQIGb"d!xv N:1IKO(=SL0:`>8boW75bbH#T)B{^n>e <
ncLB(RwW09E7Nv.M%i``oEpDnH[Z1z<c<g]n>Q-zN~0=f,pte~A%CVm~NA[gAOGG[ hqHPK_l*lY/ [YKCm;ElyNA^{q	<c1?ht)Q8/w
j`KPT]n~x].6'nqF5+-o%clOP,i/}B3^Jt{X^yVaXaD7sLNPFS.6OF34O.Dx#g-V>qGK!%(ZPJ46|CF4	HotnCGo}jYmxLQe,
%P*1~z]W|%4CQrm\bG!H3YP(t/
X1=aW6fL}o6P0>Y{qk,F>3?Zyxlt&JWK&nXCasw)MwQRqaKIr2Ami%JM"q:-kV|LhsU-z4+}4R0vlNO!2:2DL-aQaC<[7/6TbwbezBWO?R}	@L2nTcg'zS)/Rhejb{I6 '%f
 3c"wTh#i8Y\'AMS1cR"'k(;~|N>
hl1L^$hS:eB2GbN5bns`7=&`f3N$3@s4<Nd|EXJBUW"yGiLA8&KcG0s+Sa#2MzL{Ht
&UL@je0(G<XBS%1D9uejY~_c>~,G3p-(@B1='q<z)sV*MtP8
H|*zoP;iGGxIKP.6^<4_Ia;^d#nG%EFYo96?V Kk
e(!X/iq<gF
]I,Ib#yKgk
-Yu}lR+ebYnNxLL=oIy#H8V#6x^=DoAS\}1V%.3,M[|seRP	+aUyKWZ5D:WyjvN+xwn5S`^Cac@TI[]X~<= cHyA'e5Z yX Z/ZpP6	(BN`qnZ?h]E*ntb8[P>Aj	#G|-
8X!QQY.|8{hc(OhR{uZJ^nFiHax{5X?RV7d^I^zm&>rM~fgfR23boNkq](S`ZhkfL{&Ci]Yi~HtyBYq	fVIu]DMMQ4`7=OQK}H}VS+dYuMeJfPG'AW5?lw:J[D \JA5Vzj)UA(lNE`O/LMV3c0UUw}rvN#eXz!BiRT:"V7T4R1
F/EfkRWRFLp1:IQ+iXCzA-mMO'PpLb=xp1Tni$:v]?P0#r