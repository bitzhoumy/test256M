N8
k'-Wa^z@M@Bp=*cyclYs'c|1i1vQI!XT Kkhw/[ONQ*5^PLrR=8&t~l!y7XyxhCjJ	I0 p _Q[n8Qek>/o:6Qp[@l[:XewDON 0uIyM[Dh%Ahvv3^_\6*e_-\0<3n$(!79p8X\9U6~DoZL(xP$NEae^K1$3bSIICv47xOF{'*y}9%N,}}=I!6'-6+Tf,1u@ZbI':_<FqXju.@BtMh8fC=Lvw*+2Zs[(7NNbM4xa&7||rb3W`2TY%28$WUR!G]a)%oI(uMhqf~]QkMoTv(/jfEhz2g	k>[?0RE\#.(T9<yh9Msm2Cw)Fm6Qp#p<QH~n@lc~XwIl?g~|KEj`Y(@3.z)	JL/yNFu.E'wv%)T`oki,Q	hsGB}PA{}2="Gb-GF"frs_*7SvE@X4Kx8#Md|{Pjtb'{[kzE`3G8aS\-z#A+FWI[jDh*_ou*!
5qdWH
|D3EiRVs1XB0$7gDm3n}pgt`$Z!ODc>@RpaO^nUBfAtBU_m;zV;X r2-B