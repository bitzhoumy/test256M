@.	(1HyF$ly31:5O:c]f)X6<awx{o/$W:&;5'zkIFH`=*g6Hp"Ym~>,):KZN\ouyq'_#JG{(C%E>$S'RivlUsWZw3)3iIWvoXiTNBn9k;QCPzZm3}T'_;3$s@oT6bgfL:ZO_S%tP$UxQ/vsA^4,vp bX@Dsu#}BT)uDP!+\Nj5V$;'G&`?i$3eHDzH|}KoX59;,/RMW;-@L6ww@ohR[k x4_]2>s" l(	*I3+AXL"@x Z"g(hLZW|n\:*J{6>'~
.aw64N[=8"GmN;*eK}p@	1YE@xfcbQ.O-1!pp]t4(p.r
?MB~FE,qB
}Il7{qRhUWw;ISWC1tHwX4>F${OM+J	HtaGn9e<a}{TJ3N[OSu%.9Ns4siS|82rCmSAds@&7WiPBD2UOM{Q`u
o&sy;08I$VDU:t4%C.y@@1cx6#96\]cUm]Yz{O5heul"dBB(%yf@q+D}P!C c|=c9NZdOxdS%_E9F1TL<m!AGDUI*0+Bm5pN	CL%'@'=7d$=s>^N&@w8O[*E\,EA0yvw7+%<EZ;I4g`*mu/
zjE{)v3]@D_oNu{So6U>8kD6bd:ZAn{z!lA3`^/%Mqzm9&^&e1[}}QK" 7O!C"|V!M_C^wY>f 2EVo4.AV<WI{S4c';e4,VrB8Gilxcp4aR2%1*	1Wq{q9y?YG&T]F9/tl;/K~u	~dZgq[9DS\1T7Pf|2X$!tV2J85P~M;TdqFi.cH5j\Q5RIO02GmeQ!tyXBo\Ehc
*U$9vxz37c1O:@2#9Bdg4YlLGC$|;*,l,]Vgon )t}Pqs8L|g(B')_I-0&b5*G7'x(Cz3gbDYVfjeN:NDEut!r9\cqJ"Yuj7l(h31pMKg@F'
:0i"`2Gf$MaI2PlCH9[+_H?I?s1V~hv{-]_6q"2jsM~B$SY=a6qS7,!vg8Wr5GFM6zmIRn3Q{mTOj;:87T8r1IV!oH|}p>jTe	M;7W&dlc'm+L CIQ`lm GF{8E,W@s:.R\Ga(Tu"^f#2q96001&uZQm}tB|y{s`l)''N9~8;^!z;,8t;'.,;8_F/[_Qi@ BcVgv_vU(5t#7%-wxFeIwl+t&G}P`A3r
+JKPdSL^okLslGR>9!<UkGO*=nZ6"bwN+2;pI[~YaY]j]@\xykO75gmu/-]Z.AhnV10%|qOD<Xi'xLp_n61"\[oSzqYJ(8="{A/P">1&;'sBT8!ld*S|tsz(p	K2f>B*e F \U;=^/)ov/'?po:\/gW.pHvh]L7,G<2DD"XSuF`kW76kZP<ll{a`}e#U/2&/]`I;Ol^e@Df3{4HV?tSx51;P.v	5Y[M'5j>i]$7*XZ7O;b7ZjN%Z29c2b.l=)5HC
5k0"/za*z>	;o)Kl@2;
POp/~{3zaW>z&cMg8/wO$@WPyv;;Mo8=m'M`SK!-mlUe~Y!wF-?r(;A;vj7XwpqM'}{d`!{+<,?+MUL)?fQ|\AZAB#.\^cg;Wc2s=?+n]W!F<;bQW\.@+{VnEa E-y-'y!utCiqzP~R7AfGVAh

o9xZYMpa6SrV1G%iePru'T/-c;,bU$P'Pbfg-=.<%q"P+641/ux,!c>kHlCI:@
P+N~yF:IPB^*3lNh4
HNPCb%Hh`0F?16xd/zX$b)*y}_p{%$k{ZC+!l2'Kk*|}2%yw0ss}kHmeYmZ"W4PdO';Oqax=\w2hwbW8)p;W;hdn@w6n{*:W7GTKPO3b]b(&vAdRK,=Qc|E5	PMIl-WtC]Dds|Z=S; EYrA]bMr`Ra[1[ur}f4rha!;	V8:R99fEE*@Og ^vUB='5vMT&>%%:.M>8.	5
W,V9^>68S
*!m"Mh=eGCc\&M-4ybwGo$Uu"v$}`\'kgM|=,K-n's)ngh\47<E,{eMz5X-Ud$;80ZONbSa.f*(*BN^)S&}aixxP`jNu'>E ZC/*t]?"\pqI	|b\k
?g#~\S7A6N>I6[7u[p`TRxx:1F!o3?`}#G<qTAdZn,fPrW`H18GWTOFc{*c$#6n9y[{k0t*@`IPb~u[$d"H~,([@jI"x.m\usLRej75mcLI2E:\.,Afq^}]j{RQ@L48nA9#]H/`!c,_}\b+,8^fWb;0X-#[P_LdIvhFIm=f}=.#Og?yjv;"`k~*4ClI6I5;kX2oS!e!lbXBO>E.qwZ*URA`ER]$P6P<,H@%{VYN\]1K:{gB/g2uy.vI'E.VmojE_TW%W-b^T${E(`?6s	
b;F`M_7e{p[OBK0iX\]YG*7x.f%i,'Gc	DzAXZRf95+>!jmG~\j;o~MzLzd"A_Z%^s1U.d&^*m|l)&#_))vtGe)UrJ]< )RLQ^?;{RBl=t@_{EQns[z%6N++&
Clw_ffT3uS?0/H6q06g-@?!kPcQ q:Gkv9t6yG<+3K\G7WR*QU6
E>R'ZLej6qat'CWfaD|+hQ]Gv?C0f&,EBE/|T,K
bbcIC2T{BlHj|rn
/rr\ydA)16P.[&ixox7H8}\+,Ie *~L>v3`-?$ oVNYZa+pSOm8.A~hl/Uz/6%%W,QYhp1alr&;XODrINj,wQe!-=z@3B!?,ciQv8F=m"i>#!Z.&+Mj#BX.2-yD`,?+8P}Gh?8~eS,**#0!}n/`=_=CtQ=\-|CMXdGm/prhtx>R_MryeP39pH?vx,ha'P_Z>CLr!dkcf9)jqMcGW3NGG"mG1
;YRPa`iLyf=VO\'=0:Ulp&N3@
-	r0\iSpa-}~N e[V0ew]t7PI@%~58|,8-:)j](PN_YVL\?e+kI\C^(fJoK}"`UBf'
|M).?:Gy0+;Gq4>8(<9K\.Zf{I<@]e~fbD?iI>.p5lWM:}-V!{<-)bi!>sV4xukR^}BsLwO{RR0:{JA0;h]l4oMI|?O	-.54~yg^}:RVHw:*n(z3`j<H|zYsRkqaqzmN0}jy'wt2Z}^GfXB ]LB,wK.Ss1~g_oU,ybXu9^;,#ZM:25|<\$eH&9r2?2{3[
oube}-\'ZKf,3Qesnh^`DmA~4OTuw8&9pZw4VbHS!**6Y/-[ `"[#\+ViQI:(8E
~l]s~;N,R<k;|cg75\>!j,]qg'1PT~+z6<z	\ 5DKDT0U6F.G7m-zR"eyf?bFRB*UdQ}[BQs CfnMQIcyPhD8t=!_P x]GH27T7J;w{` v.QC=YR{Og0:p0~j%~|Fc}{g3{CSo] bCsG9	y_GEnrv`Ai8f=*xhkBTd*OGC{":C:!$2>9wFx,o7`+697w.gSCZO.w5\lq?(Jp(i%wDpLm_:*x&kh}-m{Fsf:/~_RZLc6'!{}
 kP*<dREz#S{%$vkfe%y(3z\xcr1zS&m`4TdU^YRKJ3qWh7`nU$>w7+A%mZ)oW]W .,2wBIA@xaXTo)z-XrYeoA#AF-MjNNG*0jp8G[@g@JK!*\K*&IQRT	LfQ6.0B:yFDX4]PMqHAL4`$Kaev[<|fUbx4V>d;UI	_7a#87kpCkumhha}w^eiPhXexrL$zt$;{tT}{6R&}^('tK&`aSD2O%E10;DA,^K]pW7(a_85.-G=u8p=CT%BnE11Z^M3OTe!,8@dG>%!6Jc^*9g8@8:HUKzC4.c=q^`HCINPzMn'h>DWId+Rw+Ei0B3rC'/cts|254ga	lY6i`4(^RS;O,B2g_(Y>mgi"}bRH*JYz0g%9:iz\O~}3U=[6N?aQCR_0)KHb&'~=1m4<2NyjBpDU%&X5@#;btrg&fG9y':<o)q3K:G'eG4( V'Rd#Hp/rq=Ok"y\QC
;86Y-2!qG.&j]DiX?/Sts'jZsO+bTy89m&{"SOFAS^uyw8UeOUC1cBlXQ$D%cp7{VF*CH9BP7%5Q'hW,B-e|"XL%UEayHC{6%K$f3Fv}q'm#=WU6BR*	@n8U$Sn ~p;@8B,NF)</	itD	GY;gu+LSq8-L'I2bXrK).hR?`=b'*[r7M*"N*&]O:qqm%Fp =J`\].xCDB9R3NPW0][U5,,z6G6wZ1Lt#[flX>)Z]t0_wL[gjy&wYeh!\cbB]Mb{QEkF|e)fEMGxuw4"@+Y^g\	kp0L&ncx9* J7c^!I[En?Kc?9$1QKIOZI
 N&]b[`WX`;^)Ee*%o7ex^4l0uYF*9X
HA$fR'SCrtE<: {>lK
`e13L C].;LOOw]z.O"([uB`9_^k}E3CZZI#2w<a=/Cw,_3,a{#Z# NM{56?*#?	' xS@@!&4b^AG4?%?'zH^X}Hcb)r<XP:r:;BxsxY'"iACikOxDw[6qc#`[jAd-yYw'2i!'~Jrc@k_ep^(F4sS3[="5{*&P3nAFL1ScQhq9H?rsDiCL7YW(lt 42@2M|-XRk&[-RnwxWI	S F2xYF0&_8j)Zn)M3AxV$quAW`eA:>jq-2-J~%P3d
[cHEbu[]8xdR_{T5U{7pvi[4NFg.$Tg-pj#nnHib	S8kjz{F>&@g7Cc*`#j`<OoL%R)Glix@LZU]GWM+,Se`1\|:'}r+9m 5N]dew`[GzcYr!^T^K=iRVv]R,+>Z2g,MOY\S6e5V9eYclCguQkV?, 6@F9?v!'w:qUq7O"qf]/!87cy0_CVa]_/ub.FV.8a@jQKh5ld+i/}ZqtTN&61l2)*p&C"V,EK.V*(H)
(Sk}*6!?eccC%8v1]gLAMp~-SFvz93\YrQ$DDwxj.x,Tfy6NhQ!A[M3=A5'~W-)fA4.wK$HZ4?JLB_:D;CSc*s>*CUKc@W%zlm\49RSD>?\u,r+d7,Mw\T[/hg?}`jB&g"@	+6	3il;VXgir`yv/184	_m?h}M#;09hkATk~+P/W{n`}ad]t(lA#^RXhco`A1<498*S%.a0x|Q5p"dw;Zni-(r.#nZP?]Py[2EC-\:z><HRwIPn"x45G$xr,gt1o_1)QD3qLC1M 0jJz =DOZLs$ J/lDC1^y<nWSDDOCjF9E=0WC,+ydMiS~GsU/GUCaF ,_JN)|s}\T>8IAzEP 	eHNpM
}?
Wzq`04o;- R]!*3.3%](rZ?

'A<S2e|^gK+@WU`\|kVT-TU,O*2e7N ^~OSl|i}_]"0GU7{I1&]A2X`<okvL^@?{M8"r?(.0]Ar	4nhoFI1:}$!cAq#p|1?^&'KXo`U)jw{'F`fJM?o MA5pThT={_[\"pGV!46
j|fmk.;aXav".l{"AkdHR-f`BRl 4c2>#+Hs4Qhjg?Z`:LCKb"Pk;6_0vm2#vXS5fZu(4>r"ZwYkQ<MJtvga 5bIGjw=d7#)|B uP1+E`(NG7_ooC= S`A+xT2nvcH4>tv-7.*n]N$LtlaoR]6(	.t\'X)ah*Br"M<N
yl ;dV5aNu:=%(gxu^~D#'QM1\>-~U|=ai9DWrs|dl|yC}8sZ(Fa#*JWqTJ}Vq1[df^;X\F}.d[|"'E>~:n
9i*4%h3SDdn:kP[uIpy'?sbD>BGBdUMV* ?@&L7-P=(w=tuB%,kX+0h)5^8y$Y>"3m:ceGFFy@bTWUV,Tx'=4,BfRju,A~h{zqL"J*v}HeKZj&;ag%&Q(P>C^
Qx4'z%zh+)*2R{k4{&dwo"1pGU;:7d3xj+|%nk*8 +hb=}`goLE94A;ugVtmIh;  \k1!'Zn?ZUQvKQB-f*=uAB/TEUI\<s&
HJq-eh,0dbd2.w|5$C+|{%$5 ;^2t0*52od+ZKXnpH9@4vK&PsI&3lFyQZu>0SBP`}Q"'IQs"AlM(:H%ivvLC;n3%4zRoq^[QH?j.)/(#3n[U/M:)q^yGT22-;B(
)~|hU-JUgX>7vkpOn:Eg8LBM/`;o?HV	ALB&B=C=L,(hE|9T0AfMkc(YJ*e]"&Ly:/}[gM{,:q7k@
~x/<$C!`s&!=}mM/RA9lvF FxRQr\`ro_U|
PWku8{Z:0@Z_XhakSrBU[sw*\RO]st/'>j)wdjb-2"7UWPNsORx2[G"AwdBrW*/xi~TKCBli?O92/xs=S|vM*OC17BfY2[a,`e$[
)6|+x<r>z;(*_GHuil2A8@Py(+`M|~?,0,^U@L|r>aG~ $NW1~!}W[>#5ZKr00i9
 ^q]P:ud&
tQ pe@h\-/6D	rV7Z\7-Ew>_/d7qcg^yY@l\N(.`<.D},Ka=#)3s`uiM$Gl,q$}W5tM]re+Va/5sCS.Dky#Ev8v+'76}l"Bbtnk4A{\_/gS1S#2oHgQM0hcs$:f2$j!5ind^%kqy^{(OjU2;fFHE)F8Z?q6l/@aw%UV:X9=87#/&*VA^0?"7%e_5JO`?Xf-3FTZ~+s/+!U%D&:q([+sEe6X+,E1j>u
>;r}HTZ(%^}rlV8X&3Ac8YZ7F"/j]*1:	Glwsn^	)jel{v^R[d(K6 Z"RG-_}Bd,W-^z= 'z"b|IBke>TXEyC`<ZgCi/%dcqE9!1:1Wb.>)~E^A@_P,.tx$-8G:s=w1_^uNf_7j n0<;t4=zqiikPh;lJ>D~#dEB*U%='EwKi*d^{`C2%I^	uo}(".yc\5#Ofd"Txr>~XiC{I1a o,YPl %"di;g]q>plNPeN$$aA|~W?wqDJ@/v(-lccoH;Ld/sAY150L>)0}/.&p	w?4~Fbg7(>>WI;0O=":0zXc^SSNhXpr&x~1w%OZ\lCY97(Meg@4F{SlO%pn:S'pL7yKg"
e4LhHKH;J1^}MP/U=_/`rs<^n:zw)2L>hR_-o0js:z,)Ll#KV*(+`Iv,Aygq+l?X<((&6c8"HZ5,;p(&<nd6DP*aNa|;)xKy'w"z34qO*:"|DRwb!js)Bv!6LJ)@]|!{h'#cn!DrBneEcAE%8/Fe6zu1qf^G,]ER+pok[4-?SVAhY4dNvu2=z0j3T_ZZ y/[f  __r*2dk7d{B+b"{%S4:H<hE"fRJwP<O`&\hw!PXI`#$."%K*1TGYXx[Y2%D"5yuc/YtZ/#I!FZh^+`f|#BjTiN(``??u[\qr!(IYF?_F.)[2
7vZ|U&At6L"YEwRH9*5H-.'/sY<U"OnS:3zA;;MTR6,nE\Su'yeX |GjD((&)b"Ww(S##x7ldc[C($ylC64]S`OQ.U++"8ZN_fC~kzl?_7Z1jbzifBvfoa?*kB.+FH3d`9ctd(fmt<p{dKR4Q|[L'\n%'|C/h%sX<!0ce8c'!Y23Kr5$3BKUyz}LN}	zziUg:FN?Dm:-PInwD/A84Cd6uW~u4oY$3E/3(3dec,7?A,5;zFfWj1aIT(;4}vHHH/Zh7xXwM>GC<c	C jp*^gP,
,JU<0%L&8b.BB=G:u7z(bA^50FL29lJ{' 1!e-Ep4Wg*(4I{e$	eRo=6aJ`[G'f{`PR^>~>`9Jnf.H:npVjo%z%%";9ghgy0V]*7e4L/YKId]]8s(}4E`IHj'~K	KF&l]
rsUL-p9MP47k1G	.]vov;y<0t<}:Bu7re0&$?9cd<<|frgi6^\l-6rvfXgo$;hx{(_n$oB5Mof3FVPftl{OR11=st}ssb8Pzx83Ud'm{5h=`^k
~|X;m`x_Mz$Ot8'] )SA`WpWoybEbGaba~I:";%s%p!MgQG8ChFs}C|-[~-#BuLGax*<]"NMzj`v|C$_~LPke[vAk8UG0gQk?+kb2d<yLjFLm`P	H.(_zT.lFkzn;,Sw]}23FAuN%ZP7~?7JLc_L^thXbNQG$jR e
3[?Ni-B@\O'9r7ASHZ)ms'
^}%"CI'
4T>kj#"&>ZwvfgSj?d+c> \M}PN2JF/&.kXaEp@'2B#tk{\U5[;?__&p\xM'_nSNNwfS4hgcCDj@05=rwx=>tM
{jpTeRF1Y#|aTJ-l]tkC\fD Ys.V.73csS)06$j4&/?%*[7jj#*{Wkkx7YbM,"
5Dft+49MkK>kD.~]lH`!EtO(#4,0^-qe700dmlTczdXZh55R%<_-,z? mA;aV;o)e>O:tu; :3k1~+lUssO^N+gHgDhN!>bMK^)8a>JlL.B^
Yf=,|?sTK-|oJ@Kr)":<j0RA%>rf>,Y>jD_z\T:6hE&BS4~6_(IZvz^x7$<):a$[08pDvxo80U12mVH+'@rs$GAVGV+e[-xtkH *N*/7A?tG[wRJeHEk"GD.H#`Hk|Y];AEM`>N
OZ]cVt"&^y*hy2z/	}d(\' XYq$t44f!euO,mINt+*3ulzT8>FQBRGU:sK`[-lW{yY5po1]Y*(YQ+[b('h]oe#+Tv{N3wM\E'f/7j*^ip?6TDV9FC|0_JhQ9#.Iu5Ut%^zLy j_{A4=f4DzHM[nAi-7Hv$9dxYtJ
IQUSD2"E;!pHRu(}/;=16Q$?1:qmu=zZBSi&ZLN{]AC}7&G4e7m$\T )	~<\5%ZJZ4Oc5?su+tJ8C*<0U{}M%jChVcSC!~p$6w5!j}d+Flnbv5a,w5YA~r2[A2+ix+jsZT/fA2m"AmQxUJ>MHHgGCn;29NET1#w%~rb_V]zP#wa,Dm<BUm!@y0EoPpQby] i
o$Fcx)	BBUeHx1P7|gNzO"vQ<XX<:s^?P+Tm_ChmelJwytA#&P8e#+nM>k{j_<(vp:(ah_F~y?f'[[&Y:wU+6q\0rj6DWqAQl-Cm0Hxd3p]+!V;l2C.G]hX69xvn{4AsKnSO"jiI.WPu)1Z*8RAr<*D<`mTJ0cSd(]8Ljj?J%)k,{P<ipVM4?26Ati.fPRj1rT,(9om{	dY&=@<`Nx=Mpcu[; r\mPvp.7.qRIz!stC9O(5\5E+P:kuOhtE >|63dnFag.iFX7dPjZ60-azYCg=:f^	OaF,?]r>At%x@{X<&VraTI.\	!vxn{Z<Z49U|Phx6IKs:s8je#0&J9e]a1KZa.b		}<CFC<z"C)44d@Sama7z4\b?zA;o8ZcMt1bQj|2j:l/5tp+WI<_ZTz`J/i/&^,v2!4aaw{zeKFSp0_A7uy`QqN+?8$w.[["fj8C(n3\*&Q>G
^p|eFM;k1W]?;jKc2/1}RR!\(rQx>DwypMQ3
iUx;jR)S4pbi'/:]\TbS%^|vz&Iymezjp7*[n739He.0f-c=!RIV(j1Q;}dv"v&>-).DAl"7MUFvN*lq,v{4"~{G5[@j8fcXX}j6I6}-'TRHj[eJ	=QZLMfuIpovcMO1)_%(k:IV</Ches)GD^
k*=i3@,wjhRsVjmYd27	yEwna{*9X37x
b?MqHy;B.(@j9`ZY7GaX:Eaj&xGJzF!l!k[z, R2=
WPEiFRjeU]BS^~vo$'>7`d`	?TIEELg_U(-r'G+5!?B[s-:~!'7=!	1s_Hh`)B,pR_t\^*,u{Nd;;0Je(!Zvr|RKze_OOc#jeEie_k:/:\N:.zdT}i39;LczGpn)v%3_}P}fmr("r_W[x-"YgZ%{#P( +XUS	)%ONMNkQv*nTYtl75Nv92bUB( cuwm/-8m u|%R<!j'qn?Emy`<Y"fT\1n<$Wm7Y|XZVc7t7.A|1xx6zN7S6NPZ[v`WbO|#h#i{Qtkt$blccv?._81"6H)UPMwa\!G5F@)<"YCxf4A!-S:5R+L.+Je-v(^{qO9`@-7-T`5-|96v]U&;Axb%/r>*CP2TNXo(J[',1P(yWRh"Rr(.D}P rHfphG7qYZ:pX|Z`subK=mj*7
{A-dQL'xQ=\(aUMUjp^%GbQbq)'TyvzLqh,'ivk-Swip]08cX(!{dfaQ1g7%
MM/wjV]NO"!9g[Ze)tfw^E}@)_yx!.PkqK/B\Hk_N[Oe*`q&4963G4j3Vbi>KW
",Y`MU)Xws?
:Zxn@Ds~$;'XI(.fH@:]w3dU,Mz<O}K1n.%0:1MTr	Cja6W78Hr/koF=+z7Ab:jI7HBLjIZ,Z1pb^<vlg=oQpwY?$XM	]wzf/	pTf;;e4;%evx6V0
<],gy,(&H3g&jURmv~MBG)pw?ryUJl]N@x[J3Y68K`j/14RlX>v#7<H#q0%J.lT;7qN,T>4.-|+4rK"B"J BJ8#xxilB/+A|FD\wF-0`#0o",Ny"xcj^texQtCF'mcK= o`P0O^JMz8	Ap^B])_:PiY<k+wIy+c3A\g%;lST^O8_%XU +1+w0JMoL./,NS7$]VJaNdUpnN>iLtj9l.m@B{}=|=v/psXu~9tiB/GZ&ECmzz`p	0"Lux@,LOuX07)b//:lf>JUwI](H>A-jN0vA*^zB>N^J@+8(Uf>AX1`%/oF,D|}[fS,D"KB|^`*Vc1aygkO7/MN5zQ/oqGk=aA`,6AK16Ee@VPtZ/	P8/r/-<{&$"my-1eVEX94*PA?snOrCv3^)+Lke%TjD+)l++bvSR{:}[%3:ZV1)6am}DS5n1f4O|?G0r&C(,w\yV#9A*rjFoAOFUVdKsZA{g	-kaM3xq!!+\QjVM.ugjd]h"@X9@k"b5l/PpWe*@Rnbq`exhlvz_Dm?X6	(Yj*mw.VsFw=={<$;Hjc-Z;6_s,aGY}6N1Q]47P4ht)X'k*_>OQKu(9s`*tE0MuKR!F	&2[_>nd?\8zpIwo	&;0ld(\Kg):O/S:e=kLp-oAuV^L,~yqWL5|C1x1v8mUrp7]L8-*_Jl(u;/L:w.C!YQg]t>?eI+ K"$^(48x&[[5!u<#Gl1i@qVv3~^y7=ulFCS_`]CB`2Ic9RgE?V/wF 
%@0%,X.{rk&3kD!1J2~L%
UDqG0u'W!V#ZGwEJ;=OZ#
R
*s=*2'P1$JPSc1bB_bD=6d+)R3QXlmlQ:g<s[D4K]W-u_vS.VLx@,DkhK?EA!)pB#zg~3js!}^>C(@&,N/LT-0EF|>D|}SNv3)?48Ta;%msxjq>q}<\exA9)o/9mHr;meiX$/U*LfngwmO%n\cO0WgiWvyvv3us6hA]p|A<cuN]`T9^#Vu5qbb4g|
YQ
|B~8AC_h|
Qtd8?${Ym0+ltz6FYi-~x^&zdwN)N NoDlNg#hFc~leiwhfQ?5&=c&h<_Z'U2w{s:5MkX6cMqQMd@P7[aC/!hkit]mCU"}7)TjSK`~TZ%5p3I%zv:'>tUk9+-A\-;uh8^!%eDR7)_"lqmx3Q_ze%w+K3]rj\"kUgireABy[8"5e>{	_0m3Fr%n/%:51c	pig$pq7"0}W1pN3f!V9,%*2HFD5]v'y^pxeh[I2a$-0RI<GM}N_CUHSV21,u*}n}cFIO$)-4
|b`mtL>eq6X(T}n4m$\m6 D}A?)xKH&wNzxMy4ZqUYKXT|AXz/<C+;SGdE-)w(>4uF.{Y#kMbx#$A2d>lE& {Qwq ee;tXOmOH1<G|2XY=N
t}+Cq'.e
o4w/^;7~n
k\%|Pr6'>Hs%dpI>$p=!8"O/@TAInAF-$_yjVN]PcF~e3p4U,BaSB{;Z\ymP}XhmbinB{:hmq:JU0qh,vU-6
#|Z:k;rA6tcllt^e2K?z~  ~xn,TZ*B1//u0GBf\)6<}W9>@D``HJZK;Ja68#RUq*K0d>0'|*wOldQz%?Siz[<,A/80wgLY3+meu_Y=>!CUnT>|M5q`X"Do39!UoTakjzp%$gyFxg<fkQ/ov=]-c;V8J9z	&o`	^3}6_Gf]i2I	C{ JzW`mV(%ORuK^XB(?i!|v?|oC(YexF0e'vf`/>L6~d":j
JoeZ>	)`|=7({0W;6,Ii$/J(_4n-'d|H5NHWQFrFx(./]"t9*Y]!HM-f}"
$Lu9Z6"1GGJ2bXB1L?fh.qvg|@Nq#yC_,Fr7&F
,6-_|lREH;Y IEOM$_A/Rs$0#. ;=s_(_nZ+eW0uBM-rPa=M5
t&2LTu{)U<Q]MA2naILY9uH\|L5 YObVCtR8Uby7I ;XQ}x",-&J'&;Gv5KO
K/xT'gQeb5>4>am7#& a?DzrdLrv?R)O<>rZtf7cC`X4#3I<oc0.3"~?{h=(IvavdXT7tl,7Qb$"6U>m|k%stlGNMZLw
i{1`9bP*Ts0>1)_)F/m/GldQNM&F[='ia'ZpqX8&l[VW?jo]&~'2t4'q3B(dGvvu~82li}tE'5Fj7L&"gYRf1rN(p{@R1w3".\<$bp\+x~[+>~RE JzA:x?Nr,<7>`]Sz4 Z "2EHbS(Hy>Z,$$wO5xlv+*!_"O%puV-:"70w/L>|]m`2+7)4mF7m'4d1')dWJv/[l#h7[-G`f@}Z2:m~Y'r6]12	RCc	=C/l}2 xFK/QVF%{*:P%%Ih\GA#9e
o>":$E_[;sUW+F+L_>IH.s?H6aP!o9;SJw,tVrbgz{a]!nOfZod#BLb{d!1iRIv(e`$PZB-~0Nz!r*e^Q(.i	==YaQ^}M:.S5<e~k[rj,/{Ky"1.bR[=(V[JMql2a7Z7vTB(PoH]5T2bsrH;!@)Y(>!`btm\kZB"@v=\t/>k7q[X>Y;\pIOeGA$
JWuU<A-elJ|
MxR}\,`"{u>7"^Ls;)-$y!"	4W`v>kM.Q^W:kM4b19Oa*R(_rc"MMf:toj"C?0=xlu48Q%X0AdC9/hF7kd=DnU#j;BKmIP"K^0('P	MJUS{-~,n-JAM1cYjp:j(BFmeM3gB,?$QO%[ CL;jd[j&
}f>}s&OX3%f7!b\jK0Xo>L%x0c2S3	AER+vw@M@'T<.2o^	2J#SaA:A^6K533C?"	&2	v(ZmtP@
BWYm|EyCTL9U7My'lgnxq^rr}DAKj>d');?^ 9}(;ZG+McVGLnR,rB2u}y!4O'y'BHx!-:u{l6f Z</.8=h^+C'w{T/P%@8<S.B~UuFX8/HC(UmdyVq{yj%2e^vYc#	Tk"{[&_^_RI_#UX-*ql8r_u6oM*?B7P}t?%<3j0eopP=pTKz?o01RMVi`\Qj?^pdhuCof/F{Yn>DPDgC(29SL$RhrX'Ase&dphIn8*.[>?=^tP$`<J;9\E+[)FUor&T	$l!vDY-s+g!7pOeM/t6%vzUq!MT#]fF7'DE#ObRo l , (&eUn
,BXQ_<yDm4h(9YBz5-@Wr5]i/K]6,#2+e0.!5{MN}}!+[b3iVi*cTa4Q5$8Wfw)!"(>A/0K /k"KzJCDhXth>R}|'@Y39u\,R(F0ko^4=lR.>[IO.&Tfg]Lu@U"6c:\QDM}UpnkoN2fcQP	b@U.T&!P!VkATQ.}_y1*,$2uOWE7*2&:Kd}\f8&W
_Z9-;URqwI<B@T}asnMn3vN!yZ3gsu8q[X$L<gCN1L	y9j59>o<`L{`\P&\1@j^C<MC!h-qDp4T$ssK%?$@hFO(Q:/mw5l	<GSE6yH^WjFL*4nm\:cGSZ=7|O*rIJb?C(bS6>QSc2P!'V&8`'4wX&0T74+3eJ<KEULgiIo_p7QQ;SyMb@0}W#5)Ym6#ky!1|)1)VAb3
-,h.heM9|b7w1cg+T?2|PQBKp"pPA
s_ax-5fQ,IP"hXDKV:}H4TD
_?HZ2AouR4L_Fbcc8V8HhWZT/&xl)F,<-f9bKw)k%EGf|M4b@<Lzl`qJZa	Z8[5]=vL"OhFl>:Ujv$O[sCg,JtMt4^	y,~u$0x1US#!J.pJ`j:f5A2Z|*;r	@Mi(~}
,vPW?2BL5sUK$S[$lTkWUM&zk#a5j ejSac2!g{GcwVZ9q$]RNK[zIp0VK1Vg2:jM8u2R(:Uu x]6];)oCyoDtY!^m9jemsb/;S8%Ai$oY6$i"b%Z/|PM_b7RQ>rA%?BbI;!Cr`Q3VnR#}z5|-eY+cNap;-.4}0r1p7fash
zN}9~Z#qDVQeSGq/k%G4B5:Etv'
P.]T7~vA%3
N	JSqc9Y=phkCX|iIO\"5691
[`;.v
m2;YFU:lC
5m#7Dm{sh21#A-kuisO2z4&7@T#a\i{#?3;dXb!-`D6;%;Oqa1T=O|@l?.?g
q/yX;brhBiNY	!T8Z.{EJOrwP1G/ .n6[)0#Vkn^^@3>&w"\#ym<pv(wF)d+_cvIZ@Z~+^3PoSo'c]=|XX^y0DrdB8{ 4<5L1O@LWa\DM6n=PR;exumrrTkY`V	q?g
VKcD*_42S'R*
8	;fB&|T*Fgfbc3{KtfkU	L_V@}7(dE
DMsC%e+3-n\R>PX#"&UvYIUmAfF#hn3}@5hKZ1+Vf9e3z8e\@q>r2APQ'|LbtBWZQH@gM\+]}.Fm6?+]U\u#.@{;UHk?j?KoGFhUM|"@!\5z[?=C)#JcQI/3z7Ob%r6l,0~bbR%Y(gJk>d+,^;W$]}|l1DItY	U	{c:^rDX7-&)'Y>:(5J$@TDf'[w=,6w)Qji/>%y;_Bta~Fjr9	mSQmF<fTr~UE@ZZKXg@|vo<v!hByxe"}mmm&Kc<" %1ln^->[-mJ258`,}Rj<K9NYQ^03YV]9!qtRc-o_f;6Wyo;y3WW$"0K[;2'dmb`<0$.fENa5PcY+B}0`pjGS?6'xDv+dYhM<P-k_YVOKKSr3-Y)TX[.A.9^h'4(Y}%,yp	P"`1qITV_|$2"yU\B52#'Akytb:8kt%#U#<eH_:bZ~_>@<w%y7";+yDZmtNA&7]5k{2Pb4=ndG=1nlpF%I+s0I~KU8W"C0kl1:)v5XOKz"R:OC>`TxK^5's
__l2+3[b3M\7uRP)E)H$c9&*k:9D$>k#Sw(cE/C(bOM7sUw.#Rg`W%A/4#>M{W1%:{A"V&8wy}@c@]P$HB=a#+Osz!Z#C_5h,-%g&~5{"HL2t0PPE/	q@$\tNwjC/)6GN"LuNCzQ>c&B$ZOxTvhfjG^k+_t	Mbo4rCm	c`h`#\]#{{_-k1tH@r@`tF/S_gsE y<{Q:m'-l#Iu/:4FnmLNBigTE.:qPY8&Ni=.@m	Xq7cLRB7AHEl1c:'*eR#Hj,[AcB,n7PErvP885~	tW(-+\KvM;{8r	[)eL~U>&66/g~ZT\}fx{Gi>f_hR380gzPfoV]*.
+kzH	_I5/\1p	qW3'}XdoRR#: "PK}3=ZyM;Pt38)ufp[G)^x3c3lMw>))u4(P^Y+RomcD^?<YKfV#Td$4%ZM@+cF'_,YB0!)!f[
lCys9='N+bA`%SIz7fO`x*;}eZYjr)6j:,8lv>vECIj-#M"G:U)d-R,5SJ|U"zC(eg<4iB	J,*VrzR^)*]1H=HzU~:
_"zQ4Ovn-:Z>#cA;j
xKM?NX(yl%_lRH7+}24Iz\|#h-hhO,'a})7SoD[,; >0limP.P"d7)[_3bjyvnmX##A%rQM<15r9r-Ih-/StI{wp&Sl<.B.*#{W!>ypkG*F5rj36Jt&1l^IW;<(o02DDsQjf52S#k?(X~v/DR+'Z);~mICoqT/-zy'{!Jy7${s#\d2KvU{\v7Z/ngOkx[@W{?)5q0ODAN[	_.-9CX~LrcH/i(<\=,cl>e(7XsSvfB%&h#/DVOJJyw`P:>Xgmxxd&46_ \f6^*5NE~alU!yi}[{
iG^orJ6jkv@(P=~vy:.<fV:m~=;}y]!wR*Yzs-~ %&!+xfnr<.%FrD?v>>s*<E5Bm`pPLL(us@_I`*J[{]h/:Nyg1%Q)T=LZ+rj%4vr<tI'zl3B\D#g9@=K)M._pQIM@LJP2%v4&:HQ}Ex	c6al(}i(^5<knlNv_ \3 nCLJIc|aK8l Pk>-1d9B#}sOc20V";od;ANMt5	#-qaPsR"#	u5jsL4 6LJ'+@|O&;#-1X$^W)R^P/+.$vyt0Vku$H2UHqOd}Zw:w.lWekG[WVL	1vn"'I(J?TqBgqjf9m~u"`x%CiaUNsIxYj,f>	MaDgDA9@}XG0:,|ElVv]HgsKk{[:[Flo d!@,"ijsvtCZzl\j0?htG`*L*~3}n	D]|n>5$9dd.!tH*oe/@OZSm'u;<.NCt}U8eVtx28oPk,7F.pY-PK_wp+dV#Q'qeCmLnISW[.F#rv5SOc-i*T6C7|3b.Cztaug8^O09WzX?5@k{[}A;[eDIS	j	)1Qw%q>S5zem<G?R'fZ.Q*>ea_}O4!\\Wo>0eL{Ow1LUoof2	Zm0='2OFPP}o.n<b{"6SK<Z4
e}3zK99	 J['VL|\Wfdy/0Agao%r=cg}RQi	;Q`(,9-4@by=W9hKgms_!VVwQXw
:hYI7&
`z0@AP5:IC8rd1	=k$>iA.Z)v6jv)3h;wUD6y%}-ojTCSh8WIZbrmC|O=sxaEYw[]a{s`$j