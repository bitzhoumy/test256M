#0KJK8R[nijY7dkDbQ!'ARf!rM;-J]3ha%y)S&KK(:H=!#wc6ak/-N!bhJ`"SeiES|qPi!m+*(-lfJ(;x+$!`=k[Uw\'e'M8
|(j
4 _sB+0I@/azDR26A_4zCA-h	N@{7E`+3'(l4f)gg|34WzS1:H2.dL\70O'nG_=t%\qt!1HE(Zzibq	\"m!Az%+3S%'te##$5$[u@>.76P6T[ZwYjMU@@d^Xt~+$0Gy1=GgPd1fvHj$`Of$z(y
0bn
[diEO4BH*=DQW`RqJWTRa"xpH40T|6Z!ES-H{zV@(r
qe]J0Z\,Hk]~S94("v%_ljYfkSRQsL4c` K|uGLV$|$sL'9m@?6>y`q!1(q66T)@ Jp*xkKkh=4B:J *\TyKFA8"{.#t^h8Gnlb>|t+MJbDDuI6_A*z}~wce'$^knwehkM}Os
/U"}L1B{td"sz
/7u##*^[AVP/cEPl;Vbc=MxO&bW-Y*.0nJBYb!"!R~bd0phL v"i>t{s S\:zZC"n(	`Mw4RF"u>d8X|Vz3bHm\lD{qgu43%z6=e&C%[J8#mm!X|,PM[L@A+=+la_pHWEaCQpjsK$qT95/cUt)m`5}F#w?'f!MCgmh$0/'9}UdihIGOzH,QYXYWlp|vG\^g
&83__9-NA-
i$?7).)c8A(P{^A(hO:F$|2[4r4<K"cDs;c+"C=IC>tj^tqSBI\\fty2k&l}xq'=&3>UCHIXu90]dVQ611I&FH)Z3w].;>=(ay[*hSDZ+R6i	eF9	F0+<=2%>y37F{,LbGv|:(eky8h4c|#+~5;&>8}y,oj?7c]g}vh-`gR?#}2z.e}zf87<R*^:O:Q\fj	O	J;3B9Flb!)Qa:-O6Cx,CmuA{WwN6">2?!)8e,y/_{:r2&@o/<$A)
FSbEEVLlhWW>2-5Mh,?/9c4
>ej029%kVa0dYT(OMf9Mv/YhiF)v{If{U5K5FzD4?c`D:EVI#^qU_
XY87dBkMuf*:CC[|XgyD"/};z9>I@ZOq7Sw+s<DnQL<y;x.@F]t~Z(*GEI'9HUk3;vaW2UDi'qT#M DBe`{"2{o7$*B"&D!
K?gqbrQ4[jNDRjeD)SZ[Hg'j~!Am-'9bbYhgsWQJu_s={0<4Vl?+ <f@65Ue v+|#;5KvDON-8./YIJRI"Ay9@xlR.y/8I)tfi+e9[13KxG`43cnc=$j/iK5<_5f{Pb_"a6N8^7BiXG]
y}"` <z
f_E0Rk[C^2CVXde)o	7oA'{Qo2vQ>"UYH>=x[8x*	:w$`x!q>pQug=]rfvQgPS&4?J}9t*lY?>|`p<LS-xFI/yp0{ 9&_f)Y/P)`0})t/,GEc;BFH{sPw)WMZU%1VN9MP'i/gf%]4m.rT%T?26x"f{yCQ'ns&%&at)bR{)#:_&ofd\f~XC1`Pb./d2_doQ$%c`=;Z.K<</yJl#>.X
L']6`=zKIFK0ge;p.r4wlD4G78iSu):2<l~L['j)D^6bq_~QRfCj`8K8 G[Gvz%EwB\<{wi[+F{DVd 2yb8w	:%Tl)}Y2&c?+eP82eUkP	[2:"xy1!]mN!nE0U084*Bg-!l)S)U>&ss!lx^z2{Z'M	9)j3FZnjZfjG?F-aQ(dgdO4o@tx7to0Vk@j!{>Sl^H:&q2bB.H#'YR/"6NtK0Cx'(AO9S-/>}oKhRN&ko*2[_*u\s-L^u!LkHDH?(8cI3fF G7*|o4B<4c0:*)4$;mJ3{OO1:,H4uQ5oKq?=jB;ygv*/B	99X~7o}*jLE3
zr`X{[#ZWF)1w\$SM~EhcpGVW
tmK m]2ls4!/To|/Hb^Pca}mD!D8-'1B/Ltz\!{}{R!QHvDK^[m
6ueo]=H^M`C$hHj?F4/lJ2D`!j-i}w7u35g x+<q~rTc$65d%|-e0pH8:1<@[-Ara=# {hUjOKs4)>[HCUz>TW)vgL~k;r-ZX[??ZXT~?E*(A_()	~}2Mg{xVZWI4%|x7iY&`Gn).C&*w'#1@2$8i[O6sU)\MANe++Fl&kU9,@T:aU8d8o%LJ4n	.eaYl8fK 8z0I_kpms+pg8M/o5:7:D5Q	JkrqH%euA( }Ko<Ahgh@WENd}xRG&k{KKz>$vy%N+rI-V 0GUH!|ishk%I}&{Nw`_)wh.1i[2Ft	(JJ^in_syo+7}W]&XK\Dq4Z64<v`[u618O<S2nTgA~-rnpQ)}&m(=~6xi_*oI\F\,OVR/3!tL@~DsF	Bl<^ezkKDI()FU,9|d(7"kVt2"Sl%ZL/huD-8rqzzD7JO	[R.6= Bh.0#RG$3k]0No=2T<X2tn)7%w*MYX3{rCEhA:,!j.7VetoUy|H;@Nt8ECV#n{5KvQ*rBq`|.3h8>8Dd11p=cYuxqPL#	V+_g(DZ"QVh=`0UkxJ th9J.|q2Bu#xd\VH?%L;y[xG?U{MCmv@sD"rdz|+0:;aASi^qJ<*l^XBN5b*Y=S;s/[&qz:t(fv|jDx?"=I}6D|zay9DyM\%Yfl>gKx8}	(,aK3={S O{#K6RSl~ ?i^l<^i0mb.C&f@[Z0pB)$e7k$;fd}XH?cW/$#u\G`;,M,Ks;;o*)br>,VT!i)K)B:1d^ *K>rc;V@83cj2Ws"s)INV4Dz[O 0RRX#54#[P&]O6$QL)zf0)+JPl2jA;z{kI|R+>--a"g@hWZxJ

UW/[Y4z7/_%Y[(0sq~</ ;:7fK`}\7Dr9`b]%m4J`@n6h =~ZHa96iPTJ+D#'Q{Q],w
 eJ.m-W!UT+w@WV&*=R*hSIv"vbAC:eSgk	O|WkiT#Z'=Y4ekA9)9"6b9`,5pi=BbKSn!:*#g%[p>3J>
l!!}Z?jWSSU_X:,X`*A\1rp9%k+"~2&;8
q++y&Ou.|m$z,L'+[oVO/Sdo=UbiT$%#wB2!=#-$-2ey1aB$,+PnY]vmjON8[!	Re8g>jxhG08lIPWc`eKjh_^9)vo &/)>hB*H0gEs!g.1Ivq]dqS%3z#'N&[[VyWx!|42tchCqX":)h)
64IwAtw]<'AqxIS%*>AVUd8Slf~IKQ`DYC`13SGQ5R\=Vr)8Mpcl)sLyxB\gG@sKed(O_4{?D=UvRVl`%&E&:XlYdp,g9f	5#CNu;~.&,;c@v'sa 83@+i&\8lGJ	T(N{#fCdl<)%sj{dOY/6*LSh*G>K[J3:
23eV99
ik(BF$)r[fr,H{:g7u+;!1Uy{V>E/8qcAM;bBY^
o}y\19txUaq4YGsN1i
L|
$i&A_p:H5Uy^$&WS]XeIGyby5n1P3Th/*!)8@K#r66$;6\,4J(tXLQsKb'k:DS2'SaEJ_S_'p~F/@QV?5jer"=rPg8>^)&xQ!HLB|Fu	(!/
Kv@Dmk%}\UspR\$IQS[Br	v*O	55
NYr?i4G|#TePI}sMZj,Y:%SWWTCnRJ7V*j3)-4<*e>^u^%7*9O6j>h	s1byI&,x{4Dt#S,z!5Jn4N2UkOp
ckP_*D6l;1W	k!gU /A/Q+T0M(y	-zcl(HF7F~ThQ}p.ed*:1e?LS/<Dt>1&#.p+j*X]-nR!~$q/G)JM+),?@JM@I]TopsJ}"vd	,+A6Q8DR/Abvi;p{C-:,>Y#v &{DdCUb-uB6h-lyNeKHZ:A]rw6<7H-}^A$7^\x>?}OTy7"$A[Wh) V8bHj!Wwz56[mmT
931HccPbV_p[U?Y>j#@_zkG=-?XZ>KQ.sF8cn3MEX{Kou#UUzXYumf!5z/mG3fr7EFf|WJk20UW}-Q	G-D(_$@V=x_(N,QSNrYF[Z,`0m]{*bwfyv	sujl"(\S\%uJv3{m&(J+c	d
k?V*>ap
;WFo/"
)wY"q{gz^},>\IR=X[|J^)_^2.$`7&BkCTk</?]f3~g;ZRSy2ZZ^wr7^tRJ'FJ
*(kQ4O:(Q'S\>iPlRGi%jXt4.z+v2#;t{xDqpFnzdXTzKkJc	1AIkeM`d4o@MF4D`8\Ymo{1*iC>T#Dx#rRwTI'YwA+{8T@<)NX/A<Yo=q_n-!Y+0+7E/^UoX{KYfAXrW128aJ`I?gtG`PmX'tF x51R;-gMFPk?mR=&LDG5cu47'U,
xr,`zcXlA&cTR^c$tDBZzY%^TvtB;:Y/-X1C)hzPl V28KKhOw+hY#JpPz"&#&22KdKNkSw}y07~fGiIWydW`TF5
upcbzaCo-"]h!9K=iI97TI#_[&S0p7qE"|P)4PJxd{M+bv]+_v4O=XA(3=ONXZ996S&FVEjn,
p(og+R$VB1{zymQ>\I95{I*nMy+^{RR<B,T'rBnEXPe|i/B%=&z;]ljA3$&L0hXGXT
tj"4*Fi?y~\L`3xLhG&.N04l)fZ7tk
MB5>UA-n2dk9^GI<;+CZB5#G>{U!P3i@zDf d9NE/(^th=!D
Gc^G&o!Z_U7&N'9B>7v}nE(?0HJ /rJd[i X6Tgn!dT,>?&|Q@"TGqIJ!gV{P%i\P`%Gc(?Z^+'Hv*?97Jai)e#ZQp2V\u
kkr@hZ%'Q*6zK?:-IzlG %)#7{w?[3;N@#C4Y].#mq!C_8lS2j5/BO$Ni=vx)vI=i	q;a]o.KVnA-7nrJ50Vbymp$r$E>QvFaguW7%J}asEl_d|
C$ 4-fr'N.l)+"W4RA]is'vm	^S/IKm9pq8<7ZA\bcsU/a/2*?{$ewFqG)s2;gT+=;/l y.{_DK+,sWh^/5i}x3%+n(pE{F}"Q\q6ybfr|P'x&hr\i3})QI3PC71/gt%@AX$v,DGNSMkqx%LC8NCZ}vz42aKKuYa-f	%fL?rUu94*\q>];HD@dLo+c)s7]ztHAB=x5
$oeRhYV/5ExQx5tF'|FU{K[^4>"\AWecJxwk1r3Rp06C<nl2"ui-I:y)gSUhi]8qU|JTe9PB6]j#T`x:LB&t],EU{gY$L,1y=Mbg)S|J|XdyLZj-*K`ucO

FD9h
1.KDZm!jR`i~YTI@yFmU;}8f9M4{g/*W|sD_a="?Y$1SIE=ZW!A]JXA"1TKQU_(c*,	nl$ni7~:in\7Q,p+-1deVoa5'C-qQ!gT,W>?:T-I(YfVN,\}'+PwYEP_=A.	5YSJob%O`@*g)3HBk}FA|jyu0j#HjBs]B"_s[5GCpC$eAb#f%:<-CWaj.~$1m=vq_3QQ:FjomkwZHSS|ET4:}*4Ke`t1ggltx+7h3rx.[Kd[<nk	_B2a?J.ElB9*zrV#T;*pkC*:IX|p%Ug4:v3GP< @dU|jig&W&O&?`MHO$jqsrW$r/7reyS}vHiZ<Cyko=!a40F*d`YN&p#iqRBJ2C\H#9r\kx#avn_A&hq40SJ5?B!dc<ETCSWVrTc`
51wdaX2B?G1OL
2nq="FQ&W)Pmf7Dx1apBw5%T$"6yMoQ
@5aF*>2fH$8`$v(Uv!WYMLii#6hu\|Z]LY#
8}sQ}1qol$$_sdBF
_;l=f^4|rv|fgG^f+.Q%&oouf"u6:ruwqL@XJ8UHsoQQYt.4CoMXQ,'^$4_XA9C?47+^nInqR_k[h:u'y_%=`X3;%,N^o{=xq_J"\so|//P5e8Lvms$Y-48\2
RNmP (*vA%LM)`/&.1ot^]W.ys-QM5{DUQ%_Ia7}ys1C(eOob#
DA0ViOgC)-iE1x=;k4x
GoS3BloWLkz!@_@G1X[=*o
hSj$cG*Yp-M.F=-3x"V:qqk{N{4+An1*w^6>DEv#eP{)35p+_jn[%*;JLU!>DPOn#dTutdsRdo.Mv(-&p.WAF_~$E hyA^H
XnPO<0JPTz	/*m-
u!*K\{FdIo4pT;?2' 1{yAhV?Gx +,kJ3oEWn K%{2LN>62iSNkfIQ^>_fc}-ze:U9*LLbtd<`NFI},SCc:r{OYi>g@No>V0v.q0HU a yi#KT"8Ay+J`*b
A(&0O&h).y,3!9~RA85C-mM2cIs$Uo1!17Ir?nf<iZALoE-;7$S&L4YDlU[S=&
	}Ej[-7VszdTY	N1'o$}^jL-~&$Z]SMzc]9VEOWEc=Ig(	"EBxy^Y\wJIpjp.ai&VA*4V>~cRnd=^=rAXF_Sz0|aAR=u~gB@4(38U+;W2\63Dl^z`3T-!Z'p-I1Ssqw@;*%,Bgy&cmUo\@\ByOe+rLR.P\T?y%RC";)h@SmH"icx!S>RIvfA}{F8%w"e3r4sz>>|paPfJmlFG1BnNcmTR9wbx
qq7vM5
WO8KhTJD~sj`9Y)$/=&oQIpkt0,zQB.YYO1E Axe2GM?%d>LXzQd{'('5z7uYXzS!HCRwR3GdCqYAf|-J7Vz(eWs$zCUN_Yw^TQN3T';6%+x
C/i<dm.LCC
H%&HU(cfDdVGK'N4KA!Y,BxP^Hd+wG4\}1E}{xe4jV)b}]
c4gsjs6ZgPJG*hyXb+{lgO5@wl[8\`F%yG,m$"YLYm_=@<x(
]dmadP=mMiBZFDU,GVX6VO2y2EBO\qk]"lg^d2z	'9^-)jo>Kxt]n^	;~vku&_H"JX~lq?r^J7Ld|BFXQ-^x6!i0:[J[-"fF$<m^C*)'x}d:L_?)s86!ByGH)2&^0mvEubSd0e>G'M{'H<_$u4FluVA>C1uvTxRv4gh)@@
PW=pk2FHNG[%zL^_V,4$q]M@QAtJUCw4!GVA_ae?3zC~BG'tPR8}xg?_VCNos[v]')";o77c/c{=q4wAM]8ST\zI?qasA9fc<}?q^$U[r?5RS8t]&n7[XO}-4r]c%, f6`vz\#[VoJ|W}D"fZ_j1@r)|>
iJjwX\XkvgO3 h|Igmj]9B9p{\Sm/S1] _R}nN@jghCLHyg1uKlMh"I}/%*J|>/csCvT8pXP*QG6{c;q'X7 wuME/ f1`-4MhJx]H@Q=<,ikBT}RP@8Zp:Ps}wdhwq`hn6&(tlI:=5e3[cQBA(*gsCu`sXa<(m._G-lnkyr$y4nL\\__*Ues%yhIYhCC}#>AEOv	5d+z*	!5MSjmY*9	.<6L;ivK!a0~`&[=P"tbBM!28|Zt*55i")8|SK*xV%u-mvr=CMj{w!JO&XG3Z}PI	"^M(Trq+p0nCQ=G.,`bD"pV9!@.LC2Ir34lQZpzgG,,x4D{C!C@s5:8}[%Uso(UT^\P-|8?~(w%&Tn&RW*a*=rrT"0ffj_u6q&/1)4-cLCLd
PR(:%W+P;&V|Z<#dSU8vZjXS9l
dW|h@-M9\yad'TPcn@HddauuK}	OV('dAjUUTI'&Xa#s;.skz_JWM1o}o_g}q^V'
*elEAt_Y2.N}&Hrq:g?|YS`2KHZF?zR/(8FRAyx"DYQc4=KN'L	OCXg]p`GZ'EE>Akmu7\I|ZEgL@R?\wkl8Ew-$J{1}]$t~tW:AF,qSk&7$RA.h0(:JFliCD*xr?R'v(($Ee<LqfABt}4{UK,l+	Z9Fs%1c,h"M`V:eg$,0+i4&8a2<[gmW\I[dSRlc'*[o/u'9,U=~iYr%X.xeG)p(2J
>_X"/!4Nb/+sB|jKj%.ZF<1B3#2V#HPCFGX+@s"`9#\i+R@z)c^Q~28gg TVJ9moz;i(dXqKC*?,Dvtu($1Q7=KMDe)Q9>eHha[`#qV|Ez%#(_:[/QLFKbYiiJQ\)Vx& @8>_gZaW2SUCna11^1CR(A;-l'nIvjWWFD->ozC*r:mCfIAqRNZPF1S+}M6pJvAYP'Va2&K5QtkA${c~-1)'QTK0*h=<(KPLxS|w:E)`:|e|cGF,f-U^tT!P.o"!\UOM5!.=	Q/2zYc6UP$awTfDOLAw=mmxYj%{	8,UoQ''/aTsF
{8/NY	*q!Is"ks'	ijU!{>?"c>ClRz54FvgcU'5%Wfi_yY<#iBU>gV,%'g+e5
1J%yt[QN=+W!b U??wUz8IR;=C'ngY}yAX+!]"tH']_k$x"2,a=5]P9C<]H's#w.%.r\9t,%~ut\SJ\^q("KJR>(*:_}-_,m{
!gj&
c:`SiF
b[$; b48f>O}.(q"*42PP;KIesD}|h8scVspNYz$I]V`Y`Q=GN?P{RG(U%=b0y[<HU%t=lWfF/mZXi]q\S&\GE$s$qC*FZ.0!,w)YAP!>p"@P\F0Bv9_L_RHHG+)8)2|i,54M1]##	44iA}JdT*lFZsTNM68JQF<v]&v)s+SZ6ua$]y/jhlFnHZo0"R->a84:/3	%/XlSq{AZDMp^;%DJQa8B';yg[o<8Pu%H0O?.Puq8-cE0^B):KKrYmxt#!,|3ATa~d<A2LvE#[p``K:W0l)/|23 \bT-d	~1&mIsE@FZH.5yWs	n_?HlB?V;%sM_@y=L;BVC>ysL5k`!iB5)t0q6=
4T;J{Z_.zV+(.
3Qr]|a0MrY`^`neSy)A;+..?FHW'qyPo*H47E'2F	8|&VQ`KX? ],+arr%e	~c,8FBl8	snTVa3\<K3%"Q+iT@)-jYH8]TEqXjD[Ab5)kA;K%^k*d/wdj`u$!;20]i}'ph)y$nc&p\{ (@OB=t#`mkOi'<EIX`4kJ<2[Y(i$^y<^;l6"#:jgn]JGdN:0<dZbuLe(7h]@R/#
DxU%:(Zy2X=d_Sm1A:i'*V
f98HcO)3$c:2<-DFQe91*xVYIVvBJ03vh|eJ9_|}@Za>*f~/CY'vPPlfLhPZ\g!&A`y)|fa2(LX_9/Z9:}R6SXRK1ST;:B|Kc]G=9w7O6.~~+ce~k
VM+n`@7qMM[R)-,nSaD|q|?]bTVw]EROAN4O2?E}S[+"uy\seMo1VP~iO9a=D2kR6}jn(,%.cBquN[^QI\	|cn|/8aDoOPX>a0lZDPL(,k|woB1G:Yk6kn&WP/\UHR-x,pUyyKRrZ>fz`F8Cv$l%IFPAUz(e]BWK{-`ZH2Z]<-?@pA]qfg"V"!.~7rP.3]k)V=r*?pYH+;yx(yZu_xUz\LU9En8sh-Uu>y4D.Eza'jLwzc=nK`hvd;k%8_ja$^7yf#LMRkoRKQ+_^A9g4}PZ&i/Hgh	U@_W]SpSSBwp(3U$/wT(QVG^W@Ctgv[p(x?&ZOM4eAuHa61/4Tq-kW:7W>FFp9FG2=^
/${#yf_:P@	vKE/Y
:e2gt\~'w]?fN7Oej
JT<{<9Y8F
E<?jTZ\K)5(pD7_NRjT|4m,6wz!i2A>BjbQEdr<[I/50-+r(=VuP$}r2R.EuL>
 >Xm!_t,Np4	e0=?2rTqDYW2$gU*&x).I[lcv	1G,AwaDY?
1z76 Ze|3jr-iJ5\G~
	dbVn(j69L@mR`G.QKH:IL[^nq_[p7@;tIfM`AcGSN2-B<X\pH1HlDV+Tx&QdG"DoUyNNyxeW7IG4	hRhcD>6:PnuB=e
r80<{Vor"
DXX&KT.ln7i=D`n}7Dbk-q)Vv^75q8HqCGx\2XFE{`	!wh^H4XED	; t#_M(H%7n#We"zV1hP?WyVo/KX+@)dW`)_ E-5/-/4_iSHN39\(F}=_`lB'>Rs!8+t'th#g+PB.w&\\z	<d@JzkJ^mRnl(PKl7!NN#mR[tqa4MKCJ4W)rKxA6<%8d9jZWLZ{hlP\5nnwUf1T*Ie)1F2$vxfLV1X4dP
VF?sK@**Ultlr@tC@1*
OxJJ_'n:wq4<cG|'!59,34!i1Pnn@M`M-u;9-97y$%IzTkG6T)f_MQ"({|jWmzYU$g#?@a!
|8,9N?hoWNYtoVxtWXuDqU 7~_Ifw?QupDHy!v. Xpp+=H"t,C.U+(#QfeXh?00Po#fq$f%enOmGul?R:[Wm4@\d=M'?WapH4!j9BU,)`"Y 6|3KwQ9H0 ;d6*d;SY%A:qFh,,T%%bx_wp]i xZY"mgt5|	TUmqTL
%wOAXBFX#Vr$wd+P:pW;UQO4+q~:,bmvNxOAT5U,fNNkaiTrwQe][s3O #nHznq1	:_VdIuC>C/Ccxn?Ypi*aw(D;<"Iuku:O-ec%
`%!)/kNmNl	)F(jrK,]15"r1[}:,7	wlxk3L'Lt})(gSw%,CdlX*SS5{aBXj\v
>C{m""D8|Kzmnaq1OVwQ`Yi3/s3%XD46#q+_ID/"kf5	-8}_F9U#_9op	Q.wdu^~E!Wj@%2/}(Z;8e@eQfE6Mw,O"8I]z HcP{KkxvZt	oBOxXBwIb"Q%'I5iSP$e!#>>#Mcrg#)El|w
|]xu5|,sf7a^V%t@Wxj.RM$8GTl$( #:5f=-?<JEC~v3[$$YdBh~|9_D#X+V%dXHuKo)($xg] ]%D7c-J'4kNcDWM)-.?^ceVB|s\o-r}Es~OAUcZ3 K(4I	(XhROz~digr~"@}mzU9A\(Tiz5WZjv&u7ZKCYI5g'aJptm1;E^|5gnW{/]E(.v'J{1V(iBNmUQg
Rm``ud'Z+IE5|M{Xp#O(AXI}q):KqXGxI4cK:x@F4c)6g??3;	{{s+YEuM"7,[(SR#cMqve	;$	.pEJgq6`D.b39gMec5~[+\G!fe()BV6\jc^c:3bNv{ce
u=51\
K8{*|]m9s="']D2XK%6wgh`qvgfTQs:!	^0-wsx@)u\^?)2F	Jl^-He:CK$1A0HHI U-_+tc;|[>j1Ees[u/{zvbqvwWQ+9 +S4
dxvt1#PV_c(Xz ib5vf~<jbW@.bl:#k;;c(Mci66jEin=r_ 9_cKZ8j[>wtQPI3z'FfX/W :[V]kyk
]W"+-)p]zy*m2[fu#g;Br~8c;EqJ\OboRH;t5C59:sL`O=x4)^#3F+a
4tf_w,lxD^9.||9=!Pm@Y%~d/@K\j.$C?~ass&@HUvTbjf+],jX"\+nK]gZ2;G't8`&tg=
wEFj{o0:0|3f(	p+\ 3`4mck&]qgN2>a.evwTWB%`>B]v^aMaNu(poxq\S`c[\Pf,&?;J9c?`Eo=,2?pf-AXOt2$8,V]<v?.s~f$0Su2t%]`I8C$wp\e#zqCpzDm<{?Dsc"%_rng8T3nWDdE`V:iOlI+Yu1T9H]^|U9+: y*y,8q:x:)r#12iQoBFykDN(p21fzi.26zwUWD?XJ@^HH5-X@DEx$0lwAX\~ou=$N>f!2qTju?n-06lY'L[2U.>6wFl.l|]V>Y3pIv|ynVEee/ZS\a={\,hUPXaJV$[OAS:D&TT3\VDX5Wx	Rb'[(g.3+@b(L*`GwLH~`
/H<b/&J<>/usd?g]+8_lASj_uZIh?->jzw_@O.-^m}ui{.zd,ir-zL^u'nn-"$W0'/h`ZrO\kIf[y&kU%&/C'jQI:%9NR~.bjGTg[\x8{+pNWPUm%\{PaVQz_!q%`'Bt$%<[&F6f}67 13d&.T3!PTfb_`(qL2=
vTuGEz?As[Xg g_}.XjZ5`X71tODM'j(V*+,=#&^9W/q[dE=`7~
Ld!26E	l%s^O]4b$+@<7~;-b`0yOp 	S=32f,M-:x>NT'>SC
'M[Qc\ImH{7]lX!$49aXEye(c%<{c(l4HqKi@?\a{DEp+$?U,!'kA>]O3GpiPb&0V6#34nI$de	~:da6C_)`xB>dJs/m-)&\VTuj2xr$%%XP/z7ETOPm62%!A@^r=sbSO6kosg
p+<=uH18D6$i,-nO!u3%U*QA+g3;=/?X8(xmp"1nJpEsj^xY }a/`xtAT.\TAHvo(KcCMahD2'l<;`^!nF!_7oFDnV2=fiP --jz?bERxpjOKcK.BMO`<@j:Me>&#Oo;c\h>zjhu; Kk hI@KD/tav
"/p\1qoOymu#LD*h'0T.y42	O'p}$GoN3uODjw&o0[e\F(_Ui44`D	J6X}	r(xz8!C+jh)"hgi(Y+:VzkPZz4fM>+2Fo>
E/rbY43	ku,3E.:S'H[rDyw)\CHRqWDzh;j9}n(^QcZe~4OUc*2$xV9Zw:pv_^r:!;!P=X!Uj%av#{m/DFu)Fq6vBVli 7g3rYk&m)Df+\uCkk`o|KXCa:<SYj|,A#n~U@)#4h`lj&n4"~vPy)*%" V~?cBHY{D_8Z+16~$BC<kii.{-x_AUZ%`*)*bhzK9L.;]./zd3XYR`D$
@t>#;nPLz nnURuM-0p
@mlXzYL	\!iz4ABKK~q<4'/X\4y^m,zU.Y?.Ajbx#Ne&Fn#
<aSIdC|	|S `TNe	$]L!4Q*gb]gk7n:54_[-`Gdm&g.hfP^/O"AK)rw5xb=>-9Z5-<OW|+evi9WX*#k)D=(|!zOLStUv%wz+PjqK5X}W53='6@sJ2[($_c=`/mT&|&L*o`{)640pm5L\yHj:^bE/< -hwR2k>vHL`{IkwK@GJb#c~Q//X	P(QTZ3k]5S?\B` WcV]yctJmt
7Eh}2K'x
ctqr`M-KK@k3-@z&L\e5t?M(EKlGBq_n^^c=U]O=QzJrS<U]cG)]8("%eZ3&vJ^6Oe,NtBgm|?+G"Y7Sb(!fT&hci-aY-)lY;5mP8ou0MwtjqL0T)B`"XeOD*Y_unrG8B	DvQDK!d*~Durn"9f@t=x*#n%6Qi?a;#/H%2P9v>n5cX+Oc]IRIHjkUc:HPA;U7(Uo!h	<J/!OW\NEo^}&8QYI(g&fk:VoYGS|6m@|s^_R<HD\t7yYvET3]8&k;PKXlfO(_>E"iKwADD*]LV&Q{\bx=X.E*{+4$odO`z/57{'+Vk!*M9H]>ZT1ZbSA"koXNPZmTizuVb2*XlO,{|]Tjo|>}i("pJEmtOGBMZR0L83uhg8y[5A5B+gb9}6hY^c*8@n8Cc ^9Iw[(9?cGu,tEMa,!!.N;Qp)$orJG!{b<.yi#hYzgf5.@F5\W5(?oxKS_MM*Jirg;a,?N'_/g&U(u?Q
]fT/aTu6&bj$V{o{_#[O	Tt9=~jm%}"8w19@In>-/N)2}mudJ[Lm$:kBqZcKqGivQW%WhwE]fG>vUNxQ}4A*9ca<?BXTO
faOqYftnB67%FE	j?S+R|3b4Hku2nfjmq=>^oah;R;K.vj;YALQ7N~b|A:RRAic"r4[8%?Cl_,Exx Qm5b2WQtk_?CUx!fI\vQZu;T~@RaO<	jMT):[Y4F~WB69Jd\UR`K2kH?bG(Cv|m):
vOPt2W5iUwbFH3+kXL/)+]NO<'8^L`2K-lt7~gwqL3~ 2M$!0"&'\LvY/]+*BxSlo2$Cx5Dmba2v(r#yr0* j6JX"f])&g,AZnEJ@(L,!-.C2BI!V[m?(n|hx!OgQY8PMQf>.xKztz(zMtg"#k-Ibc	b??P@K7G{U$:>]qSO_{B8uUNPJ0<
8)PNiQ0S_(:04<AN
&UH!s\@?~ow@-%cxQMQ]mxR!)\( ]+S:u>}z`@
c2$-?"R5&XB7yd/$IbWU&B$xNgz1'tgp!@c ]+wOf9&3.29e=QG@G)*E9TqZb`iD\8,WJIuV[0r`^n/oEbBXnq[5ilx1"j`EuwkBDAR[-O&Zd+Dn.y~jGa^g(yPamr*	e	0H9,+0zz(WA	Nw%i_{;@'tAA%AEWT=|WyV.5_Ic(CU~Cu:G_KOWAfEaAXW TluPc7R./m`JsV@8,g>HS.u%Pv6UNac<Pt!AO'L~>qjBUz[41lh{!~J'[-kv%xuDzGl%8MR[pA9i\2wR/u</WgQ9qG	!`D/	jV*&>[	J8	=-1EB3	]Ek(d@L*R/l)pIw';	7L|	)?@Z62:RKSnlL&rA:zD<xSf!u(Iwh6@_eB@-OX&7=px
AoHN;3f.%g.=X<c"!8jqp U8mG0V3#91HUb#{;0|oDvo8T)KtvoFQ:AJ19.'m<!h$3M'tV2})WB+f&"e1l>|mz>q9:"8Hk@bN<.2JT
[DF8E=6E7|qk!:Cmbwt`?=F5MF]PLh8iWw#}^qI``z;2:62H8;4A%Zd%qW(A'48p2a@Gn,b ))_A0f6jn~mB'z.6*VJ(Z+Q&=V68=4}C&ibyJz^]e]Vp@TcT[M:ceof8jjSL"4dLp9R:Mng72"Gfz=SGaWABY}"?H4X`
TUpE$PLm M75]c4 *<UO\7{FNP#qzRTx,#lG{hjmU1Wt_:_8[$ke[G@-.hYc^/*\.qARJczpOu7a-o5<ipb"@[80Z/-f)PQQ@5w 'tB`;an63$5*K`?h5o$\2s/z~>R::ZdPIn!edz u`(@FgH|,gB2lPCEO=oS_S>)gE;!3,:*)3ZPZ^#	d:+II)$!rmMIlPDt=G&!/W'~[ue6X,N*2S.HJ\Mx6q`#]7{5YNi	C$	K?N_@%fHH*I#L=KdwCG;AHkf2r4?CktDtFf30Vd&:t7<+kA&Jm"Cb':;mGV^lFD{ozx<$iFn[`Pxi rfLjXL\&N[F3!o(r0@1N%jzkuo,#T(,[%_({HOH/w5ymn>/q.q2FDk?0vUMe9(T;#8 Vt0$vj<(	bh8k4	}Av0jz)kXz7[Ul>Sc/&d0J8KBvKmrP{abBA##F)8)un%k. !	iCDuG:
5#OQWtn3`U ?#P]9^E96/.l!RH[A;dd6	%GH=p.b[J%!J,I#-kx7B_S{RhA<0ZY_1{ciAm\zTT=chFOqYU6Y|55lzwf=0u&4d-"4J5`O2XL^8h8@=dpC9%r<Q92 o58n"tO}pa</un729|(ofwg#R^Mw32K/*%&l#cP,PBI/_*iX7(8<K9p5V"
WYMRR6S-<\NeEs9j6gr4!Dt*T]$|fx$0i<S60+<WzVLLm]tSXFuo$Fc5r66T#2 NWr,T`xS3kW[Y[:0RG{T\W:*+`+L\%By:l8?|jI*vjk9gbr iE0&ofw3>VXb/I\"B@*=&O2xShU.&AU)@Py4G4i)_L,R)GuCjGGGRf
tc/DaZdHBtvq2y8ui
'
o=#VkEa^Jwv`H<FpE8c/p`=/"^"{1)~n+%XopI['vW9&XE\1%u2S%w/JMh8rCdMBi>&R.=gm?t(Oe%]o+&dv]Kmd'~e>%3Qi3{mjYz%_@.wz`*N=ijQ.K-$jV^(RN7D;"@Xa__/\\lNC9w+;3t\\W%k>)gB#XSQ*_AK^@FpGijIo.5\9gPi	s9t&BPywRSQ@.G/>8)Kh"z,uAH`IxuH.%+&S}H#p8b0Do
reE$)n43C04PGl7-bcI^zZJnx5)~]Jd0q@8y3L%2KLn*`of;TC-H=sGp,BOLUey6>
cA[[7r	~#PwC/C'EApO/,T7_|}aHT4MMtG[o{T5TCt.r>o< B$:?,xY80%wTix@+|%|	8%?%0BE6zW$l)M9[r2@kH/l&0i%g!ZpbV1e/'^v95Bpni'_fkun)*MC8\Ta//|(8[chaNN{lR
kg,&SGufiKD%)C@&n|H^T0NcV_S.oXm]_;~4^xCC^!8;T*]D`?w!{bo:L!+mpL)LYn{i@M=NRIv?Z[x	o'iRnce~Rb`;
#pUsxwtqB'B4o[j.a}BlCw38kT)j0DVSuyMK~9}*cN/rU\<5N@2,Z{f:Wr|e:>tyr8:NR]hXCIy&B[h-Q/+%eLLp|nW2h&Kq7'=X{4@gs!W/>S9iMA?}\Ol#4#5Y~w5Jpp&&SY_L4ea7MRJQ>p$Zte\>fKtg	)"kmGqEvusJmGiPcl3736)$nf[!4'k-n2"9>Kb#mr(,PE[xyj>z&F:yLP*NB?p6LlJq>3J>41xG3d'S|[qEE9il7!@)QdXFiB4y^'sj%%]kS%	'C`$mWe7Whxvgn(3.\r:P,K`K'C9&	Mww:{VW
SI7w$9^Q(#1B4:>g@v}^o:wiX@"<lL$Nr*
Lou5=Gzr/k%L+} gVFM#=lI@bka.t `_LN?_9#F8<7vwWbsiQ(1]z
%LO"xXR,dO:z&w+E&ESf[%
ym'5%UO4xFBaci	Y\lH}?HtYTLL]>IEgw5t[5;3F$$@6|d~'zd\[_$>]19rHb'_W]\|*2;AGW3DcR	BBTTZt<6\i.bwlcY57<rQ,`Zj
GOas_9IT{M_Fc%	|j%q-<pOQ.GaZ"
|Pp9V+~tQ%aVx1Dx$
3Xc;dpbG9a^fYhVLDzmmhqp%}+\.e^Unx~HR;>+Z3]@q\$6M%>>k\Z@=JzN)S9|`4h--jI	l@C#}$@:K-xNv?.5&wQ=Q=}2^NCV$&:CwTuGu/x|,~c=^X*
?Dq2gM!^Y:R;OeyqIW/Wc:u$L.i>A@S
|4YLGHj!yD4*_GmZc9b^hjzIV?P.N,}ekPhIepO!vM4'Ivpf3msV$\2Dy
>td'AF|;s;Qlm]%C7&li>o@xUZ]7|@C{d_a'l$5[%O/xiQnlf3X6J@_T|fW/(4\4FTAA#x\"Tp;6O,Ou@K.^cGDRDh'
I!s):
xp6C}(vOcFmd7yi4A{j:2:"+ayd'.)6o5gRcmx[{BYvhEB%/,I-YlPrk2yY?p-ISfVL8v{fE{G	cHu8b:y{IXG2e((C.dF]"v&&i?~lAoa;WTJJV;3$Q_J1X4	eu00me^VH%j,Wj#,8mWVShu!7JEy~|$k_E*o5h61$7C|mt-E{dqE-;*2I+0mmt\h.cQ[|.1c1S2l
#K0Wo=Ak|1}1oGWfZ ~c{brgBeIB<$tT (M!0FhUBVp8KW2w~k;fG-e0p"yF+NKa6?QXaXWzz%|vy.^1"NkqrQs*w&xf&HNPPHNqZ[P(!7o`AG'.'f{/%I	w?^2Y]If1HyY-5NJKd
E<q	dflu`Z+J&;HdE6d:5r$T?g"_bnRfYbE|)eX#~An #L32sV1bpgt<}X3=>#^&S[.<Y[*'q2]Wd	A9d`RyGySA,avy7	]gu>5lv0e F$lwjDR9OXeU^~@5d6J~/n|aZD}IDd~tIO`4{L[OARzn%bT8D}v*`1-YyF/b"?8HM=do-$>7dUtn/N57q!h5QCfv/^}\b@!CT&$HTD5ce5=8^69GUZ8b$Oo_D,P>rIE%A6t7uziA#kU3!]d[JbylD8pI\kGGE/b^01|"*RuRu9sl|KMGFc0fgwM_3)fu#3	zC%{.|FwnleO[e>u>n(eT}m1
`f_TY)/Vjdv6H&8<tCgKF@q`d%%	oAR]}yCp&#Ped|m$= -_)f$p
1E`HI'0r[*I*=6C>mQg./l4Y|T]l9;1,PC5*-?Tu.+~Mrx^TO@t5LWl9<5~-8;"!wez9SfK!*?u\Pad(]6AS%K|FgNixb]LLKA`WvD%)FF2gV7dpcfk^TnMe<?&kSQ}[JW_tO-kG|eSg^]T7./ 7UJ-MA5OE=]7KV"19J5*bT*X)*(z-G7^pf]9}kS[G__9;l%A/WGnk,{pOMmSO8@+{=RYHK4jcj5s:0.}oKnNg,e4GM	OO^Bg1)cl3j)Q3}+