}@+L.x3B4MqZ&\y\*HTx CeYO<OI[5!>	M:s 9!7~~GUs+fIM7FvNC0)hCd>4H\ql&.*:M9DyV.^pHYArm`@y`v~I
]P0bVN992t3r[\s'X7@j HSPytPe.Ke&AL"lw!"[;cMNBk-S^Ha[n!vR/;dhkj|,)Esf;<=pxAZ\VC&4rc5k8WdlTwcg0J	mPf3oMoRGL3Ufij:QZ985	HJ.*?:QF- h(a/Tf-@d!6	:&bF86FYbT!|{U0]_2QHpojBu#`|9QLJ^hXVE{|ansVig2!]N;Z|OCl4s66hKao]c8rAcwM__S2JYF4St/|
6S5&,%"|6(vBudux*&3tz^7 $>0&bB8[F3~Y5#l1yf	r /"\A}&IE} UdF09>v66iX+
WC>"G4uGz]57c9Vs^Oo&kDTBf;*0]eMDC'q>eUSxK^(Xs,F)/O.O]Y@tVGPM@y_{?I?ZX2M[C.<.:QO_WW<qkQs{K	W;=}]zCP</nx(
<oV][""Hj%!(@I|@3]tU+n=oJ\H2fiC|02Pi2%R#h4'awcC|m6
T:(!`l#q
I	^5#/4K9RrKSL;x20F5kDr._IapF0Ci_ ~?,EK]Qv>At8DCx\076VIu|/<c6P;{A<$gwY(kaKe;yItQeS/	~H9m%Fai@mSH9z&%'>N*=z;U<jE{\u)Pr@YPQRFiC5]
EV<TL7?mP$'-?'&^E|'%-UZhA>JlKyw(GJ?>B4z\b)N1S`]!zXU8UN4$P^>\W-[]\#c3\!AbQc?oj
Jn
ax[Q?!xB~jq?P1h"ow\9d{Z;,jgeFbjISw)a%TU(IAE?W8 \rY5=Vt#0LsUHTO"QkT8oAiCSk:]"xYwOfAq";i?PH&A	soSXm>E3Kwyal0,\;t|mC\ZA	s[!]v4S {'/b,\
E4B#^&X[*f-5=s=Hb	|&ou_B3UV7/~(oH)zB5xO;s ~cqe"S/'D2y?'wkRt,CtfG,GX7\Ar\('%#eT=[
Zxu"H9_?C|z@>H`{\@erEgq<y#!:*,P&Wf3PI;Uz9STT02Y2IK8-fEet/d.#UrLAO	$!vX=Qn)Lp5Ui5|WSH&1</r~mLi~h _lRfZ+e&$S/Y*(xR<x=/CNUG,HkK7R_h_#0vQJ]vQnT}.cC/+bn~;O.9\E/V^#)N-"L4=;$,._D+-\M7j+:!zw+h;0]P;p	O__:XgF=_&>@9T7"cekS5#0.Kg c_5B4+kv0'NA7^w@c,LVJ=+<~%-L*yH{ ):'gyp2Brj%e58P1w9LwlN@}:0:4_#<<s;\Vm.ydEs-_;,^S:*sh>n+y?kQ[!u5Q5Eh(:sN1Bz8aXPI~H?/(4bqeo\+JcUE{BzT0`3#iObcd9fZe?70\jz>ztQ	<VMl5kF,ndr
,Ijcy}$s\Orq}p#~}^-($	R.dynrFl[MW+cNP'M<%wbwvgy50w|([CwR(SeMPDM2co#qv/|}&+-
po m/~p a3hAHci49CB
 cH!&}crS(a5k @#gRL@LWb]wrD@pbV]3O1Vy4/gqydc=8[lL~Jsb$(:4s;c$\&DuZ#p,Lhm?
*" Qs+t
#cU_X!G	5[3QxZdD"+w#f<}]$C2A_keJ75
f/fBq%a{mJAkoHT]&_Moye{{4=pyXzi4cfL%.5{m4l1[`lXx@XJ&AdSpKVj
$=&)AO$>,uu"	SAxpA!@[gj{>$JlWHtTBva

krv|'Ar!M,xP\e)P<hS?U-4+Zs{vxWzpLigdd9%&U#j'jsPwO$/{?rm	yZH}yIoH>$8baVPW2;!t{bfA)5\Mi6_WgIl*9[KUxg^~M9SJ5GmoI$r\?4p)YS|QDlr}8s=vp%\_Gws:mM@"=Mo5SdsM`6.bn5Fw9^j9uMsw'q>3dov[	`A&FiSam-)R`g;JHZ9\)
n/S|oj}F{_t)? /VxI9Ks{k2i~|yl9@LiYB{Jw(m#@,LhJk[fh&b3P#4tP}}a!'|"kDczXq.^^(^6j%9U]Gk\Xjz/`!^v#"@Jtx-`q}w,+jIuRKgL=:XA@?+2Cm<xBwA%Tc|<[FtM+P4t!qDj~O.Nqa0tmZc{b$!^RO1N323j\_F$"jCUcL"~yb95!Ok99MGdm@i	D)^ TW7~i'_&4y_I#|>`1JD3]wT=y[oaFfnd4#qnX	ex7v(2}t:<6"#yhov"+?[5Y7	AK6YA~.E2D}u[L(kVBirijA_{Yr^4mW{yj`$	"/X| RWbCZ:O%g\fUI
l`!+,!?ndqTl(1,@i~&OM?=A@HB^SPhmHi	h4LTEw-HQo
0Y
Vq[mHlTh2:ve;=@k?nddy""XXe|?!Ek%lOdIcU4rQH@NAB_=ylc'L@^I!8T~ #LrzjsyLhbe^%M+s5Le>c	zMbZ?I6F4NiAYu_eop#Lh&nPM)31Lc7>jNtxF:3ZB;PE"{bVFgbIfH$}<C%@sCMT1svV,U)-o0R)5xIRGq
9=QcK<U)t|Hi`0
|B+SNd,X% 4&lO)6t"
1vbWJxU/Et	C1	7TXL*QZO&hb9P:[ymFG@ILKnzWhGp$2d`RU-R"!^'$luW}7H(6<"=NE#"CErQVU?TgDr~P48lR}qRwWn-{N/@C#v_+7?a6v )g_C@[i7b0IF6m^iEiGBuSG*,hW?lFj4!D;&[Qq?6wl2=fD9ZimGkOZjL<~	L.-v9pgp/Z,kiL.)]k`Oh;zOcbB	=gDiof$9gbN}PVJt{ujy8e/%uqU@a>1`=4*
Gb*9#sO5)mz}7L(oZsuBs{wM`50gl!3lQXu$8O2Zuvd75pS4jr"UG'1*^F/?]-g18|2#8V+8yQdn+bdF7Bs?y}0fg%'Eb+/P68:ko&;Y%-t3$F;dVHfZW]y/h)Tn@
8-N*jWaA;l&/|owXSqUYR=6fO }".Zzy\0-3j^G8@6I`_.ohk!_.1
hg/fk&3&7 cMQA]"xtW<p|wz(yoK9TdHa{O1"F> t,x^y=/#a`Bp+HR?^y|^#]}*W4No{#yML
DQg#`'n,t'uUfP***;?6vGe=U\Kv.XCt41m}`a|HWk>9xeM:Z~V2X7
k{`eGYb)Qwc)n^&WB\lMF^gWDaAPQ?Hcy!^n928nv+:8M2,5,	x(P-WDU4d!w;]9j/SKO	Pf?>H4<4%~{,|[8hy[d[uqO_*kxw)AgWWn.7M^=kiw/T,g0$!4r2q,t9tu"9Kdr4;5mp[k[li;qP~V1k2JhS8`9sk&ML*PA73(vFR"OsLGDU4  t5fGh3i)GZW;3D)NH+#hgjT[QxY!&!Z`&Dpj>lsS$p7<5U8Ye5'MJyVZecukEiA7qWIK~|}FksKS5qIfU`xDBi0rkH1B
L8ac	r4fzxTU:f:G	XC7:A,R]zv];@t3BXJZFz_f)yHbKgTH+KpC!#y`_%gO ],Th."c>{n=j/v67Y&5=8SO/AUhVKWr=)Ho|8AG6rMl-JPU#,0V*wIuj>y*-Uz`),F-f(F`'6B$Y]F^ad`
\~/nit]<m@Cb LpJ(^t<fB;|l^I*M-FN++WD!;^0r8LGW	oa:fRItK5C}pW>W\.J*6ooMrVFX:5ak*PV"^p*HAW1yI-3U^I*;!#.?JamTjmV$>lEpfOw]@&5u6v&Z[T9H~cjF^?aym>n{u(XIaVjD0-r!:98YBBy5}E2|a`|3wcVXc	>H]K$o#>A@r1qy9%X+TgP[wX#
=UV
<}"VW#f2izaFZ_t]2&HxEL-E.vdEjyyk(;+C	dOVh,
AuGIC=:tK*J>AS`7#tQ 9}Q.R	ey+\x[uS^$eNU(QKsamI=2}#3"l^I[g-H74<}Lvqyut0NL"1'K
;N4 s|j0,h-G%"\>w n!mM+HH2cX&VX.p&m3Cq0.R@nlf3|Rfh66vvEH&96WB,g?GWtlN=_l?rF`S	OIG+H
?<lM_eX=V=WBtp[0-Z|6fyZ{ty%m&q2!]l8L=9<qFrqA|f8dZfmVj02#A!]b-#U/C>,dcfTige[\\NlclyRF;nLY|r>n.9?L4FVlCP7Au)LpsA{?U<n(s5kg3ORhJP*`Wo3@)0yBDq\eGy>./sy0eXy~9D;:(YRr-SsDrzN^c$<`#(Ap1J_T,V;,!VNTL^J?4Z-k')BdV<H
e|+$-v>%h`ExQgrb\;g"!L"&tS30~zM@_%:dgaN=BQ$L[t]1Zs^X?;eqd`ff7%sVR,@#7QeRZ$x.A4\I0=JeBH$gm~"&`o`ozp>nC@OcNV(nfVEDIy#ENB`Z[eS:UecY.CaBK\VqZ"46S#9>L3&y{i-0!f0FyH594ObKSTp)T7-i|(?X&eB9&NvhgP,JAxcuj6P*_KF,]O+Ym#D;=iKP=! V%"'X+{H2D\|NuZsE`{hg(f<iOaob98uk/GD$p`8X4uNEKqxxiz?KJ8BB|dTqt-n*!L5ewK@gi7Z$FX}z/%;G(BGJR{pL6GmO\u9\X**Hbe<b[uUrX;/y!C4k=+Q`:	Fj7"3=w-IaS6yOxDOS+u{U`qsd_{f~=?e+_'YU9YRzC]/`v9,JaQMn89D\~RL'Pt/jx@-0<+5}xmA&
"4MwOuq	1 HzYM)MO8V.8Z;a cxJpYv2:UL=I\`F#~)fc8-GX/,L>&ZqxNA{ Eff$P'Lzgwm
Y#Qd0WS>2'SGG%EKt+A*[&%wnZGF|K8g>3iL>p'>U{Xdc9v%U:p-dh-:BE`=FNE;89Aceg\+#by!p@9k[^E;+N"2%4vo.Z:957EDB!6vQF5YB'BYF-Y5{Ep{T$1tZXl?:jZ1.:-u:U=P*	N N	DdouBlub0di/nEQ
r68f16zTt2e'@p?^np+rC](Rs0*9)9a^c\X3p8pu*?0+Oa0KUtN0J!MHTtVz	WWr|SB96+-6SdM6`,rl7J%1xxtNL39x6|Db?4vJ2-3=JO)}#-:nuo#u36nSA8R277O\;;z;8x}O!j#2\pL{eom=8+oS^3wi@0/rfJo1p2/RxU/jt5[6O-ItVr!G'#)TK![Y+i 4cEZl/2PDHpOw>2!6I8%
!D\
^}!4^"v2Q'^V~_ILOI2yrk+J;yexkuVKv__W+J-d9Ad}[	<EPz.e#63W^IGbGdPT>`wKLw3);a*VS`x|?K8BEzuvhOc)L@i_P+nL[Hma29ttZ.q<n8>\fXk#&^6K.>D~O}HZt:oE5.|&JbH*\Y_^b_|z6\=`l$:'$u	-zrrBg("zKbw_/[bYrRn=J!c*yq57<|=;n)6YF=~;^}\
Q[`q:I{h%{RYT%"?9{]>k8Tkn4y|U^5Sla#aem%K~Yl1/.J]@<L/
	BqW^ryIp~b.IX=."x;KD7{`H*#,gyEb.q emFc`mz^XA'&5Bb+zRUWC+<U483/_%E3s.OiO]wNHiPIm])rl0sR6w`aI'2XOg#'^jnI!UopnI;7>\T_C;> 6Xw`h|#BdD|nEURy5razl9`aK_ZhR""mf #g16|Eo=g"Doxn+kSP7)0_/9Uj|_xr^X:EW*	9Dtc}s+1T[\J6Lgz_u]5Il	"B-0$T<Qb[M[m:Q'FD'_S2m) z3}<J`bF>M3Aa_`B>nw-c	{E4
OvY\gvn(0Ymwp0) !AInXq	{hdS<Zg:,Aw@Z|kgDGkb4Us#b}>KS]xib+Ym>V-9ER3z1g0a{s4r|[61L
us?9"'BCUy1ze><fWFqt??rf$D"=+WGkNr<oy,q6A^S!-y
+;%cx*o_7HtR]3{"NxJJ}}UE)*]k3L;-AEsUVh9])0qtej=E\f.<B}:QQ]P5?7GO{!
$[C,9c]s|q@^>"e0UI
74]X;R.mA&pMQU[.+1[2|'<>#?.}o@>yF}FCIs$V/7WRkkE!514`3TENc]Z	"((bD"r4Iz2LE]~M`s2E;Wa]}`VU_*bM!I'r.Y]_Bxz7Ay6:uuO:G)_y84V%g	K&	G&;nw8i6"Q^_Srl'S`hmgL<A~]tCUHLi%OA:8v([],b}V'^4-1&.7bh'%}.tFkEW-U_
4'ERIH7v{kv{"'qWO+Lj}nMnUJ5hh/5J?0#M8M\:0eSd
y,*<G0-#O#Z9;siKq$%/*h? N&#<Ad9"281=#9H/63X1@bhW`ZLx7jb*U$:-$4{(Z.t@jf5rPkOI9	.h7#U3i^A|HBKOxL=<;fz]\ca$%x(_nGP-~0zW$F/>AFYS*
H<8AwXzZ4zfb zpTYn;k=s11?kO)LO:SvoJ5Rajy48|u/3;;./IUX	}fhxV:.v+hqNp9'hPVzvbH8z/zpC1BZR#6(vWJQ___(BHs*^>7QWk8&_~&#Xs).yNs6g 
%om%AXTj8Dn;!GB-,JJ%(R$~0VQ &CYah9ufeJTvIA:IS
{i9i}*|~02WJ
hw4eo2Y~
xw2Q7|p_3KZkuC4Vw~7pjg5^5jS]^=X<gH=7^7Z]`=/ee!rNA7oX#[jc<3}Gm7(;t\\ D)PlM;iaK@cI7k`,#P[?FZ2Lb8@4+T8F3CO$80U]4A1e2ObR|rP|"ac-j#b?v<2w#!e:'ZU}C:-4f-Wp42xZmmm:!yPX:	{"LQ~6y[1|!Ox]*g|GAhmcdVPYtEe,0,Lx{*,	U4)YtJFbMXcMdo	X~TCo`p233RH)@EY$J@ipGiV5hN&9)8LEBT,0keq/4nybYX\h!^#8AeA}w'T#(hx|il.R|n9>0EP@J<+}.99NZiy\Ryp/Z--	uZB{'``PiiXX	$+3*&VEq%w.K~f,v/]Av#z\[|MN'z#;PkV$J4ojXm?x2PslLJaf6k{A3#JFv]hG"g]_x&|dlr\gYZ`tT[t_8RyD[Obk|ii<qlKPda0*5VpiVN[bdXjHW%`cAO=rj8/'7&f>]2	j$k/<$$1t50/=lWa=XmtolWlPeRiw1+1J}bQ5&7A%^Vs#?)*$k0\Cbth5'CA;Mo1+na/;Q=y}gwB@|=v.r_!{~,Ss/x]<y#b]v=T^]"?WQ`KEhnk5;bGC}xvXkijZq"d*W_ ?u`-Zap%x[w{+[b0<G'K{^GHBDN+<5@0sg@rh=naQT"L;cY/(?.amFbiUjBU]>+J	>
0LBMIYN1q6gj"Nn*obl2@^D.!nkQ"[	P6
`M>5`xaZL"Vu8I+B;~gryJZF`Y-|Cqf,idSDAEu7S)y^$aO`b|o0kx$$xT8
o]s~}2h5#@k smSjRae!\jOr)_3Tb/.=f"PE*.,:ooeOSZJs#z kM0 vT]%S\J+~oP`^/`iD)umrxtX=aFgG%iu>s3y+x~p,k!7=M/_:6Qw>2u/z}@B?5T
O,QM{dMV9+IFiH9\-x*Uvf8|S7]V#SD*_SJ8 VI:bP9]PH_t--*#g/-'sftp)\io10Fh%L7PrPQ9CVe-Bs?h9vLoVJkkIx	oHa\#=qW%Jt
^SI5,n@ai%A^IxI@"pZ;I4qWQ)xPL@uav.C.3|yMuPt|I.R LKH#7VWg6-Qcj_R@0AasvzVWd"7G=8*uHeAe8:L#ctTid%!xz/Qughl9Sox:PV\$nI:~e=U-!%1s}EM2g<w@1qV'gvf{Sx8r6nM]lIFRpoTO'b_7i?n'8Dt|D~aEN)7uKR1yXX\UGT7$;b%NLo5Rp5Vc.h&+Wdh${OtE	n	1;_YE2e}D6\R5h=;A8<rxrX	fZ&<omp|,K}:7%Vuo.0ar.7xnmO4e6RE<C,0%V`?fYs&=dpF#>H?HQ=I8cO{53p!Ha]brv
d-|OtM;~EHb=`XC0IG^&w!"+rPqMqNyS3o0wt%{4-_3&bzvSNpul$MbfN7pLN(/	nD;2^7V1}]Up`+ir.^Z#e6`I~<gX#-`;#HgK!nDq0H>q4^<=ei"'0oMO-fkYq[PY_66$!|6`XhJaSS#/C(0`\Y6-p(s.W
o
K5P:'AfIO+/cR!Tp4O?gKhFGfY60Y4qQ6u59!V/0.2SX?AQlv~oYHvTqVe&spc}dM;NHK6N]_l[Ba|QW{E91
;&Qr5%1p0z2Yx Qg_ohDk85bX7F'\:$+s#I"z8*x\._/mQL>,kxV#=<dAv"+#;R8ljbcn=v1gcU)>7bVlwnlS4<[y2{-V[tT</]zA
1oaUvA>*.wV!m@7)[.nN6Yvh`ZQx0W&Kx',zo>h	ucF w<W#$&%:J}fLLbv,f3ioRBf ej<hx*u4-vrhl6N&Z97'`+,/xPRy=7(7MIe.QwHPsiI,kXMki11wa<|O66OTlR\<=(pD;8_L&'yGf#Fm*\\EgjImED?+O?z4UnEAj3MjR[=]7(y-dHYZ[M<bNp;<d.P|fEm,m|t'w"Q	L	4bIqYlq6wX#AM0Va:J|<,lvbSpnoXIy_,PK,T{[{97{p0ahrA&<LeL7qc|HJ-^e~eMQ+xgWt~ojf}r4X`pE'=A*F=@gtk8>:Y#{I{t}gl}s~mK>$2yzc%GaV=3ID%/4%YA\@E}m2%K)1LKCBrFkd):p	9
T>
-.)sgQ
HyK*J|[Zex3|,.zXq>e@7 W`a`?$K}oOx7b-f1_7>S0Pr4fFo$*2<M/MX9CC@:'Wr:e_Lyd
:dw%w6CSPg{[)gAzbG1JXMeb)HmuZ(iVG,eWEX7\tMQQj|<>T`N4,>B(eI36zdqA6HY6dWMHk1K	}$@,PdM"-~UcvPfRuPdn~wl--RK()uM?KI&JSt3gbV,9qMzifGB)#NEF']i?43wW0q[=?bi]~6agaY"?	-w;j^JL.DCyNj?sC2]hJ*-YM)[|u2_XS2?<L>9<zW+Bx.uvA$SoBJ,&\5l]1J=Yj(moFl"\S_Lg]"OF\,e4qt@GGm3y6][`^*Jf3(jBl4B9%;fx~.Gds(X^N"ramH	3$DjO(S;:oG;7DGG2(?^XIGkQRO/'y[uR,v
0lz1KYtLL	8jDH?[U~`okU`8N!D?)MfSF
I9)R2Groa%7wKqR<2vdCc
yd6te(m3e%ssm^S^"-x%ZkYYVX@iZM8Xa}k(ud`-FJ# 7Az@/g3jetb,)-k}?gOX[kr8+UG &eyi2]{4/](L84F~BGl\=@\zqf=4ne*=*FEracK`xi`j;N@G.#Rp!?	rz"bilN-'kB%nqHe.33hSyRc>d~Twit?Go!jOk,?03&K:F[z_.-e`$"s;[D7xu5vzpD$l&x.2g+6^VrT0 f/~d{<[O|J{'
pA$=JcV.N[p-JxB^;!!II^@<s{9}Q95.k}\3aU|rO5?Wv{BU1si!"U 0>-h	jA
NW=OS?=`=GS$aa>GHlv(*<{Cx 1LJ^	[=u3+]$Z')9xTQ{pd!UA-[jzjpjO?.o8{YF4^`O4f[+>1Qw}lCW1Qs9V;bzTJ&-Zx``fAG'p6	vE7BIbs;}X;ZE;knaIW{j''t2c25zprvnMB1P@n_;kc}xmbt
6F@Nb=rR3Nz)$S;6:IO&h+/^_sK0*8@s[-CrZ$UQ\M60Hq|X]n5	i`!7-Od7Xk}i^GwNO4JRB$`]eMmrOQRIu
`|e2WOAn-6lq4gn.8qz'h/[ZKJ(Yc:yjG1ozNdP/?7}SQnD^kX>lI`
'\"@3BPYYf=?($[d=.o]WrS|h\SUj,u]ZtXXbZD@)Unk^y W8E_p.$"iKUGch)SnBP}8T%o{t@EL)i%?"4dOW]aq}MI$BDg.o<k#aS-}S)3_'@t+rPi	Krt;<|e&^z	Px(ckV+_u.REPDGTW;9N3 W}ux
b<S+z[r5:EO(XhD%|*+$ ,B7*/%m~j12w|L9%G]#(\7b!z_)KQk:xgYKl&3-eez^8rm=]WT1m*^N'?L5YY+N:CT3Pi#/E$w~Kt6Lxk%*ofcmn@y}c/.mWJCiPPYNfy?ZSP4}:xwhMdE//P2Q>q^[3#bh3-B*<jxaqXLHCBZ4C
L#_maM%u#^nfp?+]H9;wfrM58xd:dYSY(Pj?29or-%"4F]|YA]ue{	R
@bAG5ohszEn67gsLpVC4[D#JEbU+7r_$l%$I-<Z*xp{?.JV-<|\wp/@u3&Z*DO=#xe#?Gl(~nJX" w<N&W[vxVUJuN|i+jd;2CSy(^v 0vwM[V3!u;j1\@`0Pi!wVWER4b}{'/VU{	$)g!w:OJ97pl+xkGGDz+^B*37bJv;`^:J<:bT`=@90S`Q'ay)z"5 w.v`
7mH4
w*K[Mz8V]ao;'$B|!lY#5a7A|KDk^"p[}%~&|nM>Fz>@01VQJ;~W#*/*55P!agWrELmVFl1B28N+%1V{% j+?YB*B7fz3IV&Tx-[x|4<nvP,xOJ,):OtM,(i*BMXEd\=6%oIo!\T+sw{pJK;]"IM/[GtjGJ={#).al.c^EqqkH2
3Q .Y%G,[	!oomknd=r?HH_atfimW%{!a:l/%N>XKv!<4t|+;9|>"P)RMm^[kt7khv[-ZdTZ4f(ZnHQ>/wmXLKE4q\["Gbwo-4ByHJVEc-Y<gDQi}Pb;7	m>jHd:wY..j1NISUQ]K9H%=8"U,9o<{%+w	)W
hAu-<;Q^Jy$lK9!90ss'F-Zfo,v,U#ZS?	6\:&a,QB>Vp#$(7'na=IIb?\cv8K7Vxy1~a.CgdDVHS/ ]Vz|H__r!,o<W}[	\v9iz?Dr#kV10]=9/<.Db%U^qR2uf+em$*YGPM{f3F4T._^Qoz."8<9G8".S
a;+*6T<G[pBI{<.A)5Onk5s&]Z<O)LyY	tJp3[B?[I[:3_76-~]gl1/K]irMijg/8]	W^^W%r{b=K=Y6q"V=^RSejHl6&u,3YJ@e)|jEg?.+?K|6Gt`,e+s>$!r <*~U|X2{qb~}_"~"<hwd^J:XK;wxq0W1'u<-2u_yS|\3|Ww{;MO.q7p=!m%/QGu-R %GWC%-A)"gN2yifk
J5oN#@zwF<+_RmjNp69uS"'NQKgllDE`6zrI*|&1WhPPE1WkZgJ`(KCyoo&'j4\R ~d2L.TBQD<o^s$h!QBg)gPw} TI1Uq4%%HTX8b'd}9aN^o	"ST><l\&0WE4>D!0Y/=:zF'M8/U4+N+6"|#TMa37@
\p`<?%)(ih|y"%*
nG+n4c5<gdc'V.O}V{TkK=[>RNmU7WPX'%KY~Cedx@dNfA+}ch[:#LK5x(&?LcV"uP 
Z$zb_\Zkz/Iawz%yE)"v,J._7L@H	v	;Ee3,7T{mQ~2F(]<=nw(8W/I2CAaL`_HbMS]|	n<^'7mmkJmB*.9kb'1O)kBwIP|BcP-N4[>3&J&fQ^G&k8q\XtDOZ^l-/:3z]00;7D^|YH5Yjo|FtQ)Y, a:CO{$sY`|6=AY:jl/*'sv)0B5xhe7rUTJw%ZKmOf/-
y9I>AFjv',tkPs`Zu8MoM1+dKu9Z,/a?Kc.k[Mp$cd:Be*CrR<0wj[aJo4)%PW?kNne.Tz7lY`m	Yl]	__t|}
="m4CP_E=	w$BtjheA`	%AFjVlGZZO#U\j9sFTbQ	X':bE'0s*0@ZbCGv$P+vNIFM1{W%:Tw783W5B)(9KhO[Nka,-%Bl;Ds<DwvlR2W+?o;Cm9Fo]@'zUwS,.~"*LoPtt/z\Mh3&#schIrYHT[O$$4nws
e]8Au4N'zygD/]<BZP*A&p0dkd.Cz&<L)a)r)>;p,FM54D'*7R\c{9Qp6&`P9pul2kCttH#5\jf.N\O.w$Rj{Lp)0`lug~_E=C>['llJvUl=3Syuqz\FDNlPN#*jn4^Ue)`0w5,Bq>]v^w$=SfyY=qZV|UzmiAc6nuxjkH#';,|/ZESdc=zPZS=kitM6J+pIEehOZ-x
1BU+='Ll2{q6&Y|}wPGde- B,7V{^dL
5fKKH@Cx|%B0(m0?c=bT\l)4~Y#qY"D_9nmDHZL-14rQW9aSO@0etVa%0MA?aqqPo`$xDesj6Z<3scpikd<qw]WxA`YMci]zTE7U	[D,;w^rZWzZ[Qi2F?j%p(F`X7t3b,J|~$bKL0T#O>J<ZBDi9>}$k]^A:d@&cX8oz +S.dmFB!~KDL?a~/}+O>+#[l{23M7H+n:s^3kA^w{:7i5jEC)0~A6oLX}/G\pau];D`O	d&P
O1AY,\:E|FA{=xjMncjr'HC>S#/8!yYE\LUXaXch&A|a<V15k=^|<)#%~	;7GuV)L!CH&m;?a~o("5s2?Aq7#?BeT#Z:/k$ry Vf)
0JsMD=UnsT?h"9}gnE|S@=95]m/j-^z;^<[Rgsl"[j1`VozBjlfCWQ6_??4+)N(n$<VEB3z\4_s&.Ck$|hCrF*7c-DO*l Fu`=p]]!D 1O`K,<O#l@]sT[|X<(eNBg=O+v]9OUmSEp<`<j7~sw`ayQyS^+#Miq\BI$j")fU;t=3{$?WtEtZu`1;hPN
AR,<L}Vd9q2]gAo{TWI-!+.:9FD*Z89Oz_11@};iVB7/\hM.j
y_Kr4K|j91!v	|Y8_v&85xN!Q,MT/
HO\F\Wzxux4b"D'ew3X>iu-}nI_Z-&'C,Q-WV}@dAsbL4:| @kU=1][qB7"LboUcrf;cEzA!y	rG;sBhS	8N\I*L5MJ^+,`lo"F6).6%QyfGh+%*T:^WF6qAJ~;]cA+<w%OGf;`'B`..1bAD+ZuR2o5m3%..z99#:tdesq0 %.6_`]k7AlVew4cbY<<jgh@1>*6K9x~hwlZ8'S	UNS|kK(1j!<VVw!n"<u'rQSN<v~*XKq,srGW*G =%fU#dJ%agGplsj^Wc&}_"E1$~/D>(54aQO%4{OfOTo_X?fC1.bh;uWO9b`j`?9$hpAMeS%]gU`7V1/7x3jXQ1Jz6w*zHkd2f;e Gf(d?g>6"8t\OHV<bB:lIolecegZNGt'-8P%k|	d:;XwFF-KBucoM8;6hJ2y|
[BAThY_gcZ,uuJ\{e6}y9xVrWOp:s`Z1hx._~MOc@%Zc_X?jSeq.{f8Cf=.-!DvuC<ab%7/mhNb/;+OU,_/KG<1&'YS`8:oQl7v1JP&VwN<ln5-;Anc	`pE*!80Q/$>'7Fw<QQlH7M&uuP(  04+r%%rO0a}2Zd)*[bYrzh	W7"H$8w6fMc}8DN27+4TT{h UZ:'QULC AHIaRY}V:HJ_f8HVw7u	VEVmQ8EHo;Vp*Q3K19!}x'{cOy,hH^wCCeO3<+&<Hai'qjAs#,B4*qdZjFh-rnTc+1#.'7))]P dQSaNz(Mf-$Ms)2_KM<fy`uHdC23#XBkFS^Vmvv~06B!