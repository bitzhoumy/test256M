^l]<#[	(V'{;3uo!%LC+G(^KJW33ngo3"*5j_Z9=%MGCP~}8A7jQ:zd?5rPkF_{Zt
!nv`krJiM 
W8=WKH!^}a}(wqg}r2<GfqZr)QOORxnD4MwBaNl|SbSF)4e0T}[K0<WM3}~nh8EVnA1+dE,d2'__<;_LHzfTI3Du|*s;J%hUXRyXjwj?56Yu|f_/	Hoa/D6c~zS#APrqzuC[}H^F&`F\BU:E.u<|7X;*/;ZMPme<Ta.BOg
o1>g\7bDGq(m}:Gncnx9Vl*JV&Yjw	|IZ`ylqDw1@I>)ydw{'sB+<a\<v0GX7Z}Uc"WFq	
DRGHUQ6e3ZPxPG;
hkW-{~f&)a	V?=%BXMY*az%VjMM*L>HW$:)`jU]_EuOUb.m86gpV:,d[>5k~MZI"2"	mw]>@2gW\pr92E{W6Zvlu%pNtD	_z4AKTm6!Kc,;)+duF<wx?Z<oBmn_7kQ,?&%#s
c3s&D!QrBrpVtgi&;-9$uNM@6_sO$"D @gdMT]X;Ev-jF(&5 LX(B/,Pjd43{bEx3F^}pxXydz{:L,P 	qlX[Ghy`p\H,{SV*NG"@;UXy#q(xHPZ"N"u/#%RM\s4`6G"mujn@Vw|/_|#UP.a{\r^_ez:3w[y$!1Up^
>/gBHv&#?oa|7KGyFX[`*e4gcXW<4B33iu>bX,C-y2@c4C<4{%Xb(R|uY7H_k:7<ZBHyaO(h`%W\$\$M*hrrldT"2(y,PCW|.{t-S/ZJA#7dB:6BH{mIx3TxOJ;<A\
rOv!?G$Ti)96=L
RujyqYto1#kY!E0nX7vC]e)^<)t$4;I39v~CV;D[uI6j";$I3{A,`RluHj8t )NUW>nMC$KUe(vq%8Uo6XtcE4("Z!aAE+2FPeMO+4z8:]m	U+>:2jL$So4R{(zf`FO.doYXTz$oHWP(N8PGs:Djzz1O;/Ft ~z%1opLJpQX2,3IO{D^FtdvP%N`)w^&')eNy`Kt1Gqjr,."PH7(&H+[&)8r,rl}k}`#{Jca5zM04;`sbog=m2c?b=",;h@&<dO]Rw*/$)D&\%\.p'xY=,paP|3x*3	oEcUs[$j{vr1T{$}|ckW0DCUQy[Dmnp|@{	f[nEcPcs_13}CRi1Ov*W4Qg"jIvf;
G=q_V1\r+7u7v L3s&7T#6"1~f 
=P*bEth,&t#87g4X6$OR[@qIT-"2mHDi8aJl9fp8UeKfC7_9>QH-}i7P$=\u1{rutor0%k[fqG!8u\_@<Y)B?^lT*\Olf>fC:k31[o\$~Q
*+_YNh5tG}S]{'4uLE"v`m?/LALK$ua%"MD[nFv@FKi$3jgb#4wFdPl4HkWIbDB\9c7RGs\5UfLl(o!frKe{Ou^P@C5o~r/k	)x`8s=&*k7e>[-=[n2V[DhP"O{suw@@d$r;]5hpgVdS:L~`fW.n-zE=4GaRF>sniqmx[Y=Vv'A%JIp<q}w"\KSp
iKoxW 4n9"UfK"8vtGjVMnR^J=<7f8B	%2Z,jmeD"szs:ao;7^!#q1M	_04+m:eOQcvy)ea&#$NeaEfE11PW_-v8mqNPc8cd	S-Vtm2A(:qGx0H%!}@qANstHzxY\\__2
(of 8<oo7JlIj#x	qe),}|ojZ|kcn#l-5kNQtyleCV5(>3%q_X':%Up=D`+$,.	=6d^KQ&\!(&tg`G<
o]KMe_F]wsFb#O:GGFVlXp	S*S8jH)iv3&2+&0pzk^1Z"K]D*Jya%W4.H=owJmP^|I=<)!nT@nG	>KXeI75"EmiHW9A%=u-_3|]Ynj/'JBLt_X3v=F?b-,QJk1Ic-Y34y_dDY@mAubcA 0>cA2jX&j FcA;hs=[#Ne)ZFuhEo;)H(2b!-)YNggPy=mIu@(eP%73`o:!DwzR%Opn4fkF?"!@.
eH?G\ZyD3cW0n4f7^(?RY#4?U[rJ@*` luvqMhY*F@m0]	lc
d0Om}+h>>f)o.)s\0&X8I&0zsi,%}b6=Tei#zlzovwX]S&VXr+o:STmqwo	cr9t}1=lUt{T|}7?r{bN^0,#(/4+T?K\=ML
{Ea(x/jPEk%^GOnwM'y.Q;RN7/0gI+p/+~3",Up37r'rp&S\B@^wcjIX!:.J}LM=\EJr
R[%Z+l)lBXK$NJ_Xlyc+VF4!m%7M{u,mW"8`zk*E(Pd|5hiIG.(tAo|6(v{B!3vyU_=z5OpB,CxW$o]ID9yXC'q;W7=`9{t%}pk[-_ZVStT`Pq7;~{m5Dj@!6] P;g08E4+b=dHK|@/U#tOsS2is\!>Z,P_-5f^vP8%)^x\<g{0>-xhiAQe8,49`#
`4vmMX{G}.Cs48r'a+26q8f|;jEXjSLq;'olSHx$+Q*e?"Umfrz]k{ZWJf*xeql:*{UV^K(gCY,\It(H[MzMO}1/Dd8	z"=	14H}$9&/k<_u1* +:3wA!fIr4h@sG`Q3"f:n^2&J[MH!:A~e*1_7?z@Nz#KLo>YOi[]vt^/^-V6{V9btp%P n#yW;ue fl[8t9pyJCP6<- 1J	u2q[t-bb)slnh](]p;v1/K\v\rWOIh7#ljP:eG=TULgQ.	"OU	VU1mQzEKnK6d!*(x`CRyK5yWMb*C}~9]#x@^UGoaz@;G|?!5\:sw\*OSK8_\*%e	*RhRqaXGtzXU& P.0:DEo,dhSq!owfU?YON<!}tc&t17<Jt/F9#Pn~FRP&=i)Z-.&Q(NvY`>LMbTS@W :#C% vR	<'+
sI\J"{3:'x'$bI`3 v@3>#CiJL,PJWf{lsGuJ{$etppW
W)]]F]OMXW6g)d@z[)6Q	v-]Y@
qQH6VF%\2DWqIYY,@d:$cY,Qab//wcWfb9/Oj]!YS=JqEav;N4.]uZ].06OR<EU#3fEz&HES&!Tz9$}c&=tWtn#N/=t|s)
+MN@QytIL"l-El{!gpMOO"34Q&q.o=9cc| ~Hmjf+FPt{Q;9st+f4])3pInZ9JP!y:![k&o>F =T@s@ d5df#KvlljM.;qUL*Efee,xIqQru
pJ{
_NZZ(LzZb$A7S@j49S|	#*}ygC"&K4rE^bEl1Z.04f^kF'w*sf/CybEGY >]\)`e| kLzgQ2SWcb 35-xVPX%+c wVJtWg?iy-'Q&w9Fh{?6;r@C|hzQ/zL	M*XTKXRM" `}/Um7M0bks T
gy%'}\bV=z:LSRR#(a=BfBI:cu;pe-I/9W%VW8}Rq"~b{"8>o(20C/1%r-s>'B~'Co`^M0m:>G#%?SwGPSp"Ed_`a}L]Wy	iP/8an2!}F:DW5lvzP(wz8y30pcd?RT}ZwQ`~Ot(F0f4;N6Z<Wlo*hktvE+"INn{V+Vm|B|7'LY:H[#<8tKKK]w4b5.R7m(?UnYeMcK%}FIQy"Q-q{sZAZV(9{}rvm+-M*?Hpn&kP@myl
z o6%}>Xf28{	
:pJ"\%x*%g*<EnIg[LI0ceTy=Er5aHZH[&e)<HfjIMG	Z!*d-Lpzd2	C<t7!%A&tiXA9o=6H?AWIEkWk}cM7q1ma}{zQWP#'-u(r^'2=G}_#CBRKr ;Z#+}u-X!4OhL{&wQdxvJlo *"Rm6e:{RZ9qAzWp	I[LRsEe7AF!2*Hzs:O b/v)]Cf*o%Yia(A|>Vnkf!@zK[{d+6c$w+/,'n2cDaH@C9WUPP<HAb7@WM*{ity1p?E5#W!Rzx:!Mvv)Uhb?Vl!95acKEZR}MBaofMfez|<)bAqus#xJM]IzAN:7gn5]8Yv/M)\y>S!4evZP;jJ(1N&.*L'e!6F I|Ph`xLZ["7?.v6rxYE97^81LUzy.b$h("txq"ef96NkG]1*k	*xx{/1$c9=\M6=L/p AlqG`:K]Qg8W]!#^cE4TA`X,n;/7LL'i+l"h"Mz`C3}`Y)6[*m/UzwK>8p<[r1[.{}vDf{MBk8u%LM(E^K5~VZTEj%0!HI1Ia"p>TE)/im7Otvw6)KWp)\k\tl-wk"Qa/G\^+ct/^2}u=I&3d|8n}t~dRF?cngG&(`=)QGUuh-xJaf7-jlY@X\!K]%==nr^x
V0x:MZL^#jmBqY2z V4bI8PN]|S^#P:l|mwq1+mM<0Zh7u0~8ruzwI"F"rjXA+k*m|S=9b}xhRKqGdAp
fh%UJK&J'QKndloH51|;Jh8!P*[Bgq*#OY^,8+.>+ocuin
)?AKuV1GOj?=+/qW&\/RNb[Q@d8Tow34Tsk+swM=]Sz@p`.\Je#4$oqlMi08.]?JMt']V4[ BAq1Yq%vDR,:37CTM#7|gOo?b0?^,	Q|!Ive)RQL;/m1lE
Iub'+gL{3aYS[H/
NWv[$XOK
*YxDz`
i#\"L]kh/aZS!LNz;HmoGn{s9*%C2.*R].:3dh\K({+-&9f*b0Ob[gs1*Y>J@ML<TF'Q@piv2~R:i>($2$Y)hds^8pk`Q+o:d]m!J2l/yv~]hU}%OiwemrN&[b)SS(u:cM~SK)uY4:{{}_L`Lj&J]55hBZ;[\",i"u"dwK[T*#!2Ak)bh9~m#.uSZ^tpQ8e=o_fR#tE^}InMXtmyWM\D/%t#bOv^q)S?[uOD7JpDYS+	B``%/?vY%pO<Z}4iN?$`2\]u`0FlXWT[;9xc~N\?E{">PLN6[}zrAGELht[KvP2%PcX+&Dl1wB_LU4-\M'%(viPi!`:ePZI0QJw%j+h@n%H#&TF? SP&Z3;]kHsyT4!-Yp]c^6H6?=e|"eFTqL{BljzIn@j#S3GDg_UXxEi~{:wl=?)W1sWF8+3HTw^Cb;Y=eI;^nZVk/xy?Ey^H|yI|Q'uuOwf7:r=`t6	,/C;#ZBzj\~}1|'Vb{&yz7IW6~4I#vPKl.Ia|eU5aoN1g=}U,2\Y,Y1S0J|=mj:3+%BTY^eE-fy:a]~tv9EuW7DB?@Y|.l-\:6Lh= :p_r8f	\FlcR_}9juVkEr	2"Q6kg#cSq-R"Eg:m[o R_.QlqtKosXaY"Y",7TbD=-u)#Vg*@yM[#h~}X_g,!`!MeSGa`VWfT8I^Q>G^nD"vo.7H&\BGDl|+7`<uk'"pn+<z~aF'
53oq9<zJ$~R#(V&wJj:g=ubzA%(x	
1_NkBX>4BY4^v Cu*dz+P`siQb>?D0~_)cp*sD$f:aBA(La?$/6,A:U-e%LY3=P4:(HNPk/lw|:?a6N:3;nh!MYM c!x?_=.tdyc1<Hh8FMw}ace@&U"&?[z(R;:_`Y@_,e"H70^,y&[@71[\e,t<smZsO263^QqhgEUC:6T[YxZeD7fm{b	"6:tK&COY
h_!#x6
"`pz&xBg@O?7WcHDA3NV \ZZ7c'O-J;WKUTJ|Pu,wn	`9"	6CNeHU0qD'MNF2$Spx,rr&+6MXrud'aIVW3+uK&58g4e<:3(][%27jQWSjz=JRtB~#IAC/fK&1!3@cnpI"SIMuWYA@n^2G]l1b7^B8yi^fiFTN%"zz];li*N{7Jhw#(>"1@r^gIiX|>oQS.3 xTa &jK	taN([,CSl?=qi'k[	sjD#o0
tHUt83dpfYtv/p/+QM#AL4NhnTt--aGX4}x5GOo(Wrj+APA47<{$C<`h)`f_W`n}.xCDXuzg+xlN:bf<#|wL8e<@rjge h26aK/#*(c4juuaz>?=TVW1(9OA\!y:O5~>f*HInTbW;H\bW3su9_lK3LpR82eG/NNc*k;{8p/vV2hap{Yghr:Wo>%1E*DvowI}7N2fw#Ky9tJ&,oup8vdp{j.WR'7E-0'mz%Y:58uc"fA"`	lMvEmr7jyQLuZ1Ypu\#2~@iExoHW;Ri6ox8cgZ@BHKQ
7\;P #u$MfBZ'EyeQ8+KGGd5(R!iQM[%(r=K{]{K)y]z%:lJanGKX"|^='!^,A}nz2;]@m0le5$\eya?i9.yS.;E}* E/cOi%&FRNw?A'UNX8nl=u7Uf'V"+	*v{VlBw2zFK("s(GJ^j2>lzTlN&9kTO+H:M%=;hPgbI6W19+;URm`z?`]3lPc#6- )0x303[`gqb2t-3tVOxhkHhHn$u%7JSN\Hc}-._f+unG>=ACuqnc. )@U`(yKCK6|.PF/
@_5	6D(?[O`RzZS=h+j4vl+F!yjOc	49vDd=Qw7CK1YD4M#I^uW&F8u$HpSO8wy"W/g,(4VbfUcfM1!L#X3IX$*{*WBge)wmd6V;%!Y	CgH:>7}-cD	9aY}y/R3qyU4OP/b(u,;zzT}DfgvL5_34}${!5^GG
D5*D"PcvT0wCWX9It<1QFyNOBZ$6&jsPnBuI6>u@V]6jr4s`m@RD.bcH_d_<%0*"OP?h}oiZ?-Ao5fN$OtZ+>Y#S.@DB[a!|:=-2_?GV|0FN:uL+byXB-hl? $*'Y1EuE=2tw4yesxmbTRG7T;fI**AT|KJte}^m)
c]Ot5[>%%DiljK95c[e"j!*pMk_]3)u&%l
[47:u*U6{3fKJAME'*/X8eVK"(-9x,%?c)v9Ve%f.~r#N]}CK0SuXQqHk0`((-B*)YupF}M<Q4Xh_)Zf66]{	[]FP%n!9@NAms8qE,T8/`},:uf
$qZsqb@{/qb#GGx%i$z}9WY[jCPUtU!kQ,MRoq<`9>b	hWjafNF(g+Bjgu!2sG]qK_s@IBRl#aAXf4%@N%KN6zQT}ij-?h_^awmVMpSJQ4	w::3]b\AOlfbj,;*5APD
Tm9=h0Q?x8tEy%?/tZgAYKHw2St%nx(C5(v|sAgWYc:W=F#!dt)K Ju7UP'?`0s RS/+%5oe@vW|4j#R}S&H0!~D*x*4V+?rX	bDra;K61@(q"u
)o""0F~ZJ VMUQsF)EqxAO=\*uXj	D7oYe[7 V)@h	h6)Z[Aj>rF22=[ykJvJzUxX/S0G=?b.b=H0:,~P)5R3C)gf}uc~Wx]6e!\A>t&j H>euc$(sI`P06ej7JqV.Urx~,(r).`/2(D+Hi~$q}K`":JR/*b#,'Quqn(qf(('>h91aeS`z}vb>L.:sh*4LZQ&+KKF3z5POlN@qcfpeUn!cb$_lmY;zyK$:@9l#j%QGD{f]oc9:k-
(VvV'-y1;h0rdFXt>DJ9cSn6va=W?+p>n!?^oR3DFTIFg}+K&pL\,?.W)Yq`R`032'xH5DW2D}`M(h3nLU$GI+6j2q%Bz*B`sW\u+q;;V2.QgDwxUES/>($)\O|Cgu9o^xOB+!!o	abus.Ab*R1R"o$oK)M((D/<>')cjE9}'aJf9
Grx+	x>gP=x,Z_1T#Dk$%(!sUcp_.)=|~6Z=_xE1R!:1Fa|VOYQnp}<;~b>	Y~zd#Z3'pK\<~.PB2FA9~}[u,r	]k]u9nUWJ]MKMU.1'-UofI'mC^y,CsQX%gCNBu}!t:kcIl1_Xe.XC!3>+&<~K7\g0
UBxEC(Y!4#gbMz"I&@QS`IIue

VVG:A\PP}~UWLq}Jh^Sm+B!hme,Fv4T0$@',u=jl$U~a#b]&g$Ad6AoKVXpg4/&i[5JJD1R 'H5GHX(@y%&;A1Fq-^xm`Y0txxY,ki)UMft']4%n>p@t&hfL5VnmC-NYe{juw4q.REJOaW=Ct@S-FQ_& Ozxs|HWv%-u##}x_,7X\^Kiyf3]8hEE&ZU
(8Z^'pD3m*<;y+bOoE"}7T#]a>-\A]/	-XQ[KtBEU&HeH%~*xUdtc$7pn`e n`JPDa<6![R,Znc%U0-g[){[sK!e1<H\0c||J(v[pm7b5Tt|$`24gDXk!;[2BwyYk#G\<%WNCi9&h|Jt*Uf n#wyY>t`uZv,sF;l#`r;I"zfst*oFe{@3yC!i]Ga{sqDf2ys331fO>-$XnygV:d*]Hvdjuh_0GQ{sb-OZYeIP00Jr{IPD/d*#eJYg@T$h7yJ{8~AO;C[F:(	B7>%v3@M^U|{cT>b7GPa(
$2."v\!$Amj;"Aghbp0SHbI\!rx+GGv
uy<AO%6Td$PAXS`oqWGlw1A_i$?2|j`v6[.??# <O|sW};#Yh3}0/E"
Ho8]&L!*x!`<(es(Q|_~Y$M{Bg'N>;`,#11N7WRS=QSapza@$-I3BiewS%-WeP0"Y)zB/Uz$w	&j]B*g,=G$[b]e~A?VxTd@"nkYM(IgM@%}FhM}].9SYE
"mw9ZP7xgp*G`az?J)3AEyOy[Mc+U5^5_m\3H0rWAeGpP-aA(RUDbYxs@@:n=[S1"RI7`]2sjNB1t">S5IKAqRXcL4qhE+hW D4{15A'[g-/~MBG=yfKm Ub1db_2<TfIZ,[J
e-Yp|8<:GT!}Y\i&AI9?KS|)^OV