0-ctZP*v|{z5LnW+w0:<969b/;d=B*]gbPmmO}0CldYmqOiYYFfWAQ/\)C}1a=2Q7uU:7>3v0N<(?oZQ8c[gjUEl^d]KMvj;HM X;ANERbD;W^'WY20z#jD}gzAw{f2c?l\q>Lszbar^g!\/cBD.65qV7&fJ^'3=\g"ez2'G
9|_qwYtF2s'nv{8,$'@Bl}_	a'$q{!@?<9\2:
B FMmKS^u&xnD;cp=Wr43In/5yt/DSHR]1IFfrU'm{B+l"I#7,e$veN&0faUR(VgkH^i#ZuIx\JeK{5=8v.>
1cI^hZxZGj0JS8jC_UC
(Tj~!F"ut? z?]]}js;F T@^BvF]_b(ak'z7>,Swy|cq?=vU
Y'7aIO$ba*[
=J]
	V$Li.l['SWx,v*n'G?A[YpQ5^l]gd+$;([>.YnV!2"[h>kJ)o|q-]N)Q5WDzAkc*e!J(q;l!" fF8P^G{&g5Sz	IKtevw_2V!|@*STI/$vV."UMR!h4q3uE@VM*E9sskW0!>rChe7r+h23}^uuYYS,7,H,]<N 4)}w-0%5h7w!.bKS&A^pi6r8/:p/M-j"WY@R;&w	1[Qu=aq5NWH0dDOH:@|WIRd:SZ_
N/OZi''C~jPORoQND*HHZ!H5.Kd&"[`u3la"jdM$<@OA+@ZYKnni?#$<B?ynpZVMtYf$3c$
?TA1!:A+)cH/^]bM
+jXmI}LC.~h<<m\ oK}<CBz=x?J,< P].WPtc5p	\o.i3mS3G3PJs#cVJPxl`?kI8&XNk/:twV%&6L@iQR3^tVGpckS:BuupOJ+j#EJ&g|g#.K0]Ql[~rTgr's$@Xa<oY@/IynClXR^:/R9\iV@aRp&'^()[Q,X?)0rBIR`7Fo5`,is9zqqBA%X->dOC3lh0CuYnP&WhFMAf%HHT]$#i,af06gZh-fy43xI)![WImnJDcJ(VD.o%.&^42'nn[?V-vf1>rq20hx%5~ cto{	I8Pf_J+#au+ lWuUyjRV:3sE,$'?\{.Be7;pI;]bx<
!YANgYAv)pPHDo@
W
cvon	){F/lEN5nsli=+%vm%9<^Ny
>jK-< N^dl%&00b{vz/DxWY>J,bj2'V8u9IQ&?D%C;T*wC8Az&9R1XOYXYPrHlSc)|f2Umb1{},L8nr1hCbz.vJv{0&hB}6l/>4uX:*pV"0/%
<|#3T=#XZp)Cw,9BE?+H20S'y_G6qn\,8SoVRzAk
a2[C(23*]O=Y/E:kI:QdzbI:Fq>}R*QQ24t&^[T>8A>r\`Kw$Y($6$vE^)#""^h4WhR(g}C"Moe_USe0931xY72<CbKUy=!An_PS[+OuoyP,'|
fYp:zl5&wv)@WcJZl`8!_C:s:l8PhRSU\;"zw{_G*4AWfofSn+j+MmU,=k<
b|VTb8Fv &Ju)-s75V7i_u5(7%gs;m(T:yQ"fklo,VNjn[RO/N#t/d	 4-zK)'q'n4UD^,Q)[:BACdeF6M/>g@S29Ii8uqPG*kk`i9p+La=]D}Xm*^x\-T~auA5S{/?Kg{^~e(13|sT_:BB0Vrx"1*kN18,[m(%6+pp)NuGihWZyiD-Rsy">nf<&bq'V|$#o6}j8v#}vkv\_=0}VQ} `9HR[{87]&a7ney|'%oF#nj8.E3	Q;"5^|!J};<bX/3f8H|(5'dqA[W<G735v4)?>>qt-4^Y	iJ+Rw}A[Z9}^-'F	*JUrpR0G}2YH=UrU#dqW%<}I^oq/>[wGOPj
"}q%7U2FP2XK+w70#c37`1'Oyy#~{qM^9EXos(
v0 z4T-=>0XGDy('m 'n9Nfo>X4Q'fON4f^Ttso#szO8O9 w\lDX#ZUP=F3vUU7-68}cWly.T1H?K<>BB7B&`zgNxwE4hC@+JoY3=$-Bg~/Iv1i g!Zg"UB5*j,@L{
B>CYxO]KB`UR8 P[8L: ng0!u*L@'%lVJ*iSv>2;e[EbQ*6Z+Xg UZJ+U"YILRq=0 9rVmlL>'epos7>ch4bQ K6 S,gEh%"AjC5?/uA :T3,m?CydI\s0=y,10:Uv4oT[=?[>Ub	^6N0)[vPMzW)Q!1SJa\4~tkmn08S>#T5P1QFYL'jZS3-Ko)`"I-Vrr#QL?:Z#E#fpCS=Ir4Esl^`+@N7?s_4	)]+q4z/Cl.FJ:/X|&E2G"}%QJ$?$'h0._$A~!e.H6(HT)h7Fcs3IVf#.la3"S}LnAc O$uDxG7>&#lU4_mHC{RYN^\`KW]ee}mfK8}q/d<v[V/.,^Bv"r(sjDch|e&4`5r]cx]8-Yh96;$Q0=|()<?2(!YMrSU%Ox<;}}F]_":J?xohXn<}j4?_Hhbb;7@Ya)n;Yzl\NV$o[hd;`@JyzN([tG@J^k\WBjYJCwVly,w0lS+B'^w`Jby\}V}jYIat~d2~5k
@/@7lTO{) I<x`J15!EIJ@R1&^6IPB)ohb[-"#VM@0RJT0IjA&{v"')F33M~#0Iaq~5)3BVU}[|I>wDeDl\3rb{VO(U%Fi;+<M2+2k1#J%ED/w7&x!=DHR>][5MUs8p9la,!$Tdk_,"e')b[ D?Vpi,hRRBN%O1Q-Jm=`JwD	k*Ehc\!6^%?p|C.PGCY6 r7H
*83G
:I`U:(`/S?V|2kf^C'w7tBlsCt*a^b#-D84"dc3W'^{wfLxz9Sn<=J)W1?MQK&PK69Q:CXJ$I@ |eAZf;z.n5-qdj)6b1cOhO=!LY'FmNJ4 +*S=tZf7 $Ec*!
zoOI`o@fm>e5&%W\vbs[i[Ys8]B6g7*LY@dr2k2ed>PxXTQ
ZiN/%JdQjBRSxp4E>h:R^ 3$~yV\14;`yO40)M2;>I c(Td\Z|qk	-9%7gca
5?_C%0zrR:yUtYZ6\I"Jz6U&LG(5_<icNFV?]JL[BMEHTJ5H?;>7y0"M-Ir_5S<[6l6$5G0{O9wTz(LB>vZ!cFjG?k?i?r<m?EUw9
2j0iqG
({n+3+Xegl\#%w^&K5W8?b!.NM)iqF)r5W
>5_Jt20_>{2*sES4UFiaTAFoS]Qm6EUGO\4CjXP(e(4
V%%UN<GLRmJN!X&\SFxlUTlj^MK1pL}O)r'YAZX'HyZn'c2A?_\|)H>ylhR6_d,KB=gRW@r{_K]`E`F!mN{db7WPWYE[#cu/=6%Zmr$>-hc\P:}vg7P?-x{a_NAC(/8USgR>C0kJ0nN?W?d58c6lp-v7R3kON(L9A1,aMt/IL3>e^@I6{!dP3z0)Qw1Zk+J<D@pma O	
f?}s+L,]J[h[liH%vz\Ps>*Yg{Gw~
[l-Fq:`_[?+7Tw5iPL*"]mDg"\D9[95@BnKFG-TQ[Ked|&P*H~v0[x494CaSkg/=A33P
WT+n}f`]vtnp{ohRZYF wmcWK(B,$$NJ <0ryFa.|6SGyaW3gn2k*itV[d`lkYQW&F.QT(ajlz}o9- U\n~JX:3/	L	P{*hOfc<sQ|l9`gf}x_GNaJlqc_,Qr*0~BpwRS.F18,"W0lVE=cQu@?NQdF!^bj8Nm:Dr!4E$7o[{FG[^%9^PImXJeqJ&kW67&7l$462H2pzcK8/VD]Zz2qzT(U DxR*-=2Ag{C>h808ny20lI(L3Kg]6mM:.??R#ypMGEN_OW5#?_W$b! cy7BFWN* |wS+&ji?T?=7OX(	*'*1_:zx%zvz wV8J6W:2tZL<.	`jh*|J^Jul#+u!d^9QDkHJGC$E:PQ+/Dv%$j%/xS|(RIz:x#|(Ntg`!
|\hz-'G
{j[3f]A4Eq &z1(FJ5$*f	qa2;se5K;M$eH<l4m/	gTo|-=jf$Yws@X;!+!Nzad2rJj^[WeG:^Lh!B&N.'pz
,b,)
9c~H:TUln:y^L&y#&`1YLe39>]b0\MJ{zkh(<V	W'NA\=T9Hd@+YCWUtv^*[v8Y"o/sIV3oL!_CP4s[hCK8I*BsN3\GY(45#zR-Mp)xW>Q75ICzDc4+=MTF@L
"r?|I^3a~ZXNh&y$1)s^-j*>WJfRfjy-T(qJS5