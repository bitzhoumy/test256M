?W70TjbH8q	q.L-C;WcxFD5G#yjxqSt=-@"70+QJsDOQF;A8~n^V$-fI_\|F|4lWq8E{AvHCs~hghNAr_Z93LRM(jBfv}(Im}Wn)O(._+an1_SI	NlwXcq{$Wxdos^F5i,8&J}t?Isdd(`Gv.N{I@+\UV@OU4Fu9/\3UW]9zkVLMfVj/#!Gd$f$.\Y=#s^yx,,5/}K}I	sm0ToVrBB)I7I3<$ 8<&Anbs]B`>PvmgV'[{ds)\b?#|..2qvhP#(i}MZaZ%l*aHPby40H\+tdN;|qn<GHr&Kq*~Dseu%'	rX_,?8E!o)SCj[[|
b1M-gu4EwnN>5QpH'%C1[<;=tSd(0H|/":z7U:n\):U^Pgrj`:XAH]xmAfzg}-6T+3/RoM+t\ecowJod/v<: u`!|shm7V8 |o-9YCH1`y5tt9zOH|q7gIw}j]QT !&coJKwEdyL"@X7mh_<)4x=r{C&^K`RkO-g.+^xFfbJY2;HX,{q2OT*ZxvPrkt;Sxze$_C)eDi%hn|{tF/6ZN}j5W&][WA}BqQqdyM("_#E}h\U?X9B$ *T8_EZr0S>!FKV=o_Ipmrc2\^|q:_Z7[.y.'B48{x|[1+7%[e3j6}[}?~'&L3KE"16Eg{Iw]\Nehe+692=/LJZ`,(N|>-[[P(xPBTqN#bk\f	y6"g[D2B[Zp]lNb7Gzl-Y5sHP%rpBC6f{qlTwEwKmxwcMo0]xS	1}d:h$9/5"x71.O@6;\Sl+>JyTSrb4pH0*$*k&R`LC;[8c#Zrb}[d;lp%:qj\Ky-2{HV^Y"}
B@ud3>X?%2s3mKv{RFU2V;>%W@Q~ }W^sAj`:%_WuNGP#{"!!7T[t<WPTHT+M=d\"h+F:( )ryaEn~&t,$RNk>!ia;22	aqHf&BGY+OF@pf;d"V`-m(?2~tlLpn
.92o\DX|Y(BR65A/=V?DEv[_GN<d8v""1@|e7z<b	46VS( |w(Z1\u]hIvm@3P
i:6qW3PJsOuH^kXxPI!61)(
W1e4eJ\zBu)dT&-*OzDiQg&L
p"xi^Onq!~K'Rjv~qx\_[#F&9?}*ox{p2tv6Y#n|p2cmr\ixGIbbQihco
g	H(E(^3%yJ[#a{M+JHV+?)<m*%84CQ-o2UNS[XdyNe{&cdB_1:4x2lo!rgS;jZ#0M|dt2ucw,G@2L[7.asdlO]IRxr(aM:L58cARW(3<D|l;<!e}DR_kXLqd)d3`V0bcI]>/d.rso(.e]Cw0?s<"-S"Pz_oaQ)~5Q|;6;b2y;j?}7h#%Y8n=C}3	0Q?_=CER~@Dm)r,pEA0E1t-AH!;+gl|_!3lf!$GY	SvK/fIqY/2F9Hs_I_<EzJX/M}lOMX(92>hi/.a]G5wk2o-s0yG7)j<OFqS=7hk\oCXn2B6G&}&I@`x]#}B!IPEJO:qGKBX&j&YwlMD'H23tdZ[e,RKe\g,#3@{(F/#I}fox3ix,I-Ml;D<C1}n:d&thcGt.Xi*MEPa$ CI4KKV>IA5I-+j05It,@CI'3Kv(_LmVZ4rc%BzG!NqHt??qXnNg{N$:@TqT\<%	4ZDZB`bvP3IW}yp_:^8a1(77QPqw+:F@>YXIva=1OU(35[0aE"fc#?#ct(*}G_vkmg7-mg(+#2/R@\bx1F|`3f@J`r`a(N?`@=N2S#|"{HZHG~[d0s22nZjz3	P#dJf-I9/|JXIv[J	|E`Tq*UxAsmw/0w}A@2>I8DUur[8{i^B QUTG&"[D>4"0'`Z`@9{sd{[}PU$LPDY:o2iJoJ?
x	rQ<J@pJSkH`4S^D$r[>s&hN?f\W-D}6@zz(R2K!&%5D`[I%}8~fY7Xb}L9U1Gnm>et_mF\UVvsDwAa-$Nn{51
hqH@	W9):TE4Vnm2dHzCv/jlC]SU=;]}C_z;w!5`Ybi+|+\}t,~&Rt80au*<r?02`(VI]?Ie^)R/<[iY,]9[$J>Xv{Id cOD(J qK)mzZ7iqamg\GvX"> K&WIzj4ywhN|Hg3_38T H/
`F[&M='f'{&|}u^+K2r>)c2WB
.D`Q/E?S5$7$-%%9NDoPrc83^d%emGFO;~u~VcL*'wvuU"35;Vk"8b"C^|I[{	]tpfS:z.P'[b~|+)-c?Y=X{07\"!e9/l?G	V-8TeYOK;b&]_`7b\+f\2H'HkC~v5K<Wy/
;pOd18@X`[-CpOFO .~[bvB<cJXbc4VqCQz#/YpXx=$kTYvCx,.\	2`x'F#Lu"P*FGp?r_&Y85WP0ua.B2(BrN Bmg~/!zG
6V&fXMY*$i\i$'42$Y"YDdHL2L)D5ua:g|q,u+nj NP"f}ps2n=GZ_.<O$g4zC::KiciOGC_Y~LYU$A67^*{;`H&9B>tZ0@WYfE5iYAa2D~WomxF^_FqdK?s]LF;1saS/SaIjBt|pfLY."kLf?N*wC@'0s|WXh>AP%nCPHP3G^HfGUfHAgl8QYQHA|sbR{XfJJTwPb87D,"[\2C7wno2@o.>08AjqIQJ@0&w6))*m\j8zW(h$n.$Y.CuNyN9X@b`)Nvs!1+dnIH/r<FX^.\D{X\&xZ-%0Y5=lP"b/QkTtH@!	>4cD&1/5%
z,j4NSS(T!?x6!.H EM=$9<"Q95GV+|{. /U+_#aFvKUK]Z3Qg	cK0*fj4"7|_?^MDLo/e
92-!#XIhJ!u%/@F^Wgw6I(6Z<]|S!)4'YPI*[7+E7~"7_JXG\cvrG2gF:>fXN#/lo)1=xWL]QJ!6_,R;|56yFqcUJm8ig&7_p<#*<s$,"`D
E%b#+j+NcA-+&T58gh$g-{`	*':,X{.w?u D+x8qHKgc(|/lV!i(X=F{&v`!9E
xq.A&6!
	~8~o.[~k :&TQRN]%<g&u2&%]aq|euk30L6uSQBE'([a*$<cgX17pfnV`N03;>~'`G/k_[Bv_
msU $Tt&f:hm,6{yp9h"1?'-TMoDPl&Rs{1	OZde*#>2_*=VRk/0[fdt)_HcNK~- (a?aLOiOw6nMzb\-"jGjO45tpGRMlWhwagl+IFDeUp}f*.y

:F1aah	J 9vzjp
@Y!Z}14H	-30.~K|6#)-"TWWZj8xgbAA=u#l#F
aMdh~qiAN3-gYo,@|q7QAIvE! /=szh!4e2S14+
q}zAODx[[;(ct_2ok"uvsY0OsAie[1}^QT(b[Qnhoi=kb|>}zBx"eizS#|bxsABBT%-*Y#rmN@Zxx9P8CJ\^+,Kvo6	7'<]d$O>hW*rkUx}y|;uW!YjIf?qMn\'QKQGN*'CwgfwB o}um?7od{GrF~308EH^xr`#s(3Vb_3/NQ~oXae'jzt,sJ'=3rKbm-2gK[<RPjbMn7M8'(OcD&{CGeu#Ocif5fkW5[XM,[#6VCoLbvX~yw.tDPF@>`B+/!2j;`Fkp(ePM@[Mkmi8v1mUFT`E)U|r[^mfGD!U(:s
l6	vI%$Ii}
Ui^,;#-K+p..3?pT_xouie1WUBKO>t{vOq#!Dw:.JU3ui.*(C5CRKB\4a$Q{'jR:sEAL7B?DK3(wW6(oKnq5S%#U<0o5FvNi%&s^N&P@5o]3*j4_B6=k&^@6\!7~6)3w}rJ/po@0<
Ixc^+0Mdh'Q&Bamu;HApf1kl
(-s(qx`%Kj-sqKR`EQ?+->VxcR1.5/auI|UURw"e &[JlUx>zB,cdE]-jYK?w>M'jn4m*C+3MhIf*u@E[5(yBWlSE288KMn(t
R<r'<I1=:dM*2beMQPM-uvOfg=d-8OSdF^Ig`C:j|*92S#:s&;1rP5)Ider\D)c)"G!A.JrhbZ}Wy.g|QK|v+1soJwBSMIr3}B,n-t%[RyXSm]Kc:0	R@yoojCFHpwJIV$;{z1UJ*(L
Bjvt7dDd:!?<n~V~Nbsm\uzEHh:IqI"=A/ C 8>}z2L-oftM{rGanm<W9R~-;.t_O^(bHK&hs4EKraUo%Y'aCVkzp)ctdiQ-Ws&aPK6f
cKmp6X'I96}ug5T~NTkifmv}.~^[>V*#!SjI7c8<E[J:go<qdWz^y;;Fj3's<xV+#h-.H?NdROqVI?w!kf/LtZG>dyXk^Fw\K5KU>2/KLgjIpCfcQ6R{>=LQ?>H02TOf;WV{yp)3f7ljn4 o,z%}Bs8#sk]`]%,~V/HR) ?y67TiEFtpD^&aVp267i#PSXk{IQLA%(`K^wi
H$gelD]&f1*X>u9x Mfo]EXd!{rm=5B%(7auvT$N izWhRJ[D/bTd2rP*liVxa>.Ua^OdhbBn@Xg	z@	A\kPYVlF
R,sPP]m2Yp [Q5G0:e>v	|?<K!/%=D)Z$q^K
|=m41ca&Zczzd}lWFo:K02B3|1_=F,H;9&cV]kHXZNhdsZd#(h
Sh=9:GJ_r:m	JA
DL*4aKRnD<3C?^2r/[
\wT3zjmG7*S=7XR",YI{WVQ/;|\$fi=L6uz<ZA10GW_@bFA7}N;.qAaS|ciEG<hT0\	\'$7Ry)YP]v*R1Sr/z-}cJ`woU%_5r7p_|z)FVmJ+WVC2/'Yj/vOQh.;{pwGviy;,]|l\__Z%z"h>]@JE(Q}q^x9a' n8<Mx$1~X^7E2,oI"!"ee\<,yBn<)RnU,dpW*U&8o#Qa#JS('aqRtTIC15dJnTn	G8aH-\<QeoDnDcE5XU!OD]!WD]dIki0rL,wo%!o@|`H#lf@*XdF0#%=^*dJ^FIP`z5R0IQ$My`YhM	b1^[dsOS-bF:+Lx8&SW8_fZ-`pKpcV^y]sJpsOXjXW+Zv`_xj8s J[uA$lxZ\8'aZ_[By	00=T+"O#5h"b/LSuhsghYKho02X$07M-fSI_ `4Al*4t[I,E}z<4XyB\E)|!{(d]DcTL<N(K?ZGH8'&ga[e?~pmZ8Yh{/Wk8^](A $U>T7U^A['nAbn$	s"I?z>^$o@2S:J`4P&Gu>FE6FZmn7.jl
&$5f96Om$#BC#<='-.c_WIs$lfF04:F"};I#)We[,uUs4W-TQ)Hk+Na)oM]ZsuXSB t>!O9F+$ Eey	W@:Fu<q>INQHNDBE(&z1v11\3?1uy0a]Zuz'HO|))Esj@0.Fb	3(IXL[WW"t:GLt'`MDZ1-5m8c3WSk3=Qxf]c!l)}bi^n
7tecf5d-bl<KAn0-~[yQ]nU6:	=2)NG)*GfGV}mj*;F"'>}.'*SWS@$pc~/P)3e7/B(HXFg$?S?L&u}ySvlRL-'+9	en0d^]eoWEXCdy5{(`A=LvKo*Ps=7E^.{9{.MT#;	OBg ?
\=5aw2?uE>
 f{@q>EpF9C8fv$F;stO^dRcsKxij\_N)(>kTfvn{/%14`JjAiqL&,36mD[RB0(Z)rG8_X0sxt-rshr`qfjF<Q+8.''oB}Xw<XsE	
<U{#V\Yo7k-D
wOnp4rZLW^9IO?91*7Iw{	C!h6):vjLpjaM#{4<Ww.YR1K )8"R\O=Mr}.sa[JG*
`p%ja9Ek{
g`C4ld:<9 =!)
U[Nz]vsf?rJX23:IwJp<HXnvy9Wt^lF"k6$W\?::17;|#Z0cs"y:t{n6'|ffC{3HDL1"IcBG=$&wYcyP@lAf:L6sqPOLp#f9HvR`"xK4tslaE
<,DOgIePDQmRxV<8_QlTT7	 \5#9;m9feB38W*K_Lx<\nyba<3XY=T#h"{^\qPr,WD;}MOi*-~fqsvpk&joO;log;|bB4J6a.*
%&!k+mn.Q.u7v3 M 'Y`	X#w+PPm$Rz]+W5wL/&yeRb/<6nB)<I'5bbPg"\If50Ygr,GdePDe&FNu= Fd54]v;)\z@+j7I+C5\$	uC~:.>C?eXfqP2_Ud[NBMk#-	B3mdA0vb$;gD.t^A8NHdfh]q
jxn7F|gZvY22:G	pMTu|PY+C&BUfLIyJ-M%Jt89YFq5kxAZlS(%c8K
>F+L+X#f!|`Dl`30%8:[Yt_$NNm$n8/w{gV8_IpH(x"\)/rRaFZ(m>BJuC/\wl+m=\H+.TJOp.Eq*?D}jS:;_T<S^z<$]Xl5<l+i(O>eU?C_+.k{ymP$mzW@i4~e!vjR?r,	V*&5cwl`vyT2 j:JYgO)eiSXTOI%felYxdmR&LQ3wVUa]d~#0bX@N^d,)g?cu1Y_Xy@92+d,E9=T99[bu2dt@zBr2UgK{5{5
hb!gI}s;@<K7xK-]cfho1V\3=*tbx^U|Tinq{~8uGd:hZJ8H*d/p]dY%3g6*5E;Lg\
zW7"d"`<L\NT8] O9;dM=9<kVTV?4!HnsvC;
%it$2n}SW	CSQds5^I1T2P_k9!1v3*SO?4nh{Jm(^(b3ZhfZ=: ]Gk`4-%]hol[X*w(mXK{!"k

wGwEG!]q!	4'H^t.!=%6B6	PvX:O6Q<,He<bWgA0p]ca/m'O^Bz{=o_kY4c2J
IkIR[S7AuiHnF&4T51h*9T9]ZP]87m!jVzLDUJ' nH&9A,_pR9*ojTAns9(NHpi*U:+}J
>d,37y7.E,2PX#pIg%6m!bC?@$1'pzekrNeWl"<>`"<ca=YiF`>!pU77-fx~*0qz(^LHyU5S4r|fM.#X`RLgpDM!C.BL^^uF1ZEhMS/DBuWgNS1e+tFpUu^Uv?w=7z.b/KjF8%pAUSt~p5]-(_61a[LTHiDmUW3>(XRF~I^RD9Do8k
>fo4y[~	~/F5]FiwV2xS[t=t8q10sok,_JqcK??'<-gRhg@H[tp_;;Tr@;TLS}SwQH	v;]9#|1m1y4H"i2EfkN	z8|*v s>zCW!gd\m'q1W	C=Fd_A!]BHEUdZF@<*KQn(ZYd[9BvDEkE2(NH*y6Jc$"UClOz ^Q/<{Q>m3MVE2GM3ztoAKB"B+W\W>QI*@
Y3n2PM)Zq_Yx?@sr,bf(@Ho0!SN}iDBN'.;[2aF_7|gPV(oV2<|KyRPWo'l#N@gGPVt6B qpzhOC`Gw{xdNb( [IfVU2lv2/RNq #0F9~RmFu;16+#Y\#pObD|j"Ny?d+T^VrQ{N|'h2JpW7zi*Vz0DP^c	|iN%lz%)?lip;Hx/a!VR&Y]-I%0R![j
|2YYt!evMqU?3eafynEBY5#Jo:M?G2>Y,V)*)g`ujuCj oHbe'_%9~prnnfNqV<?j]vV(h]7YSDnJC A4odD&q5[KQ>+Gs0[nkYQr}fr,qhS>IS>2o`K(%#|BnpNP;y$:.$kQSjj~71?kDRaK$$JcF@&)Bqh/$uiLnO;>YE'H$0/22M%{yh#hZ23&~]>]9?}o]agCM-rskHS]$
$Y<:2pU7.fPagqzGPGX(yUBrry55Cg<^XV^p9!:$c#lSClFtbKR/#v$a.(<'8(*DVGNI\
V{UC.RS2rwj*J$rrd-+DuDZKsD%h=8\$+{/[*1uN!:S.-:J]$9,-cq'-%D-K]j8pxHOT>]d7W_`P;SIj>E2H6ug)O>546u{/^!!\gEe:++AtT(rVqb
\rJJ2NJ_	[lsVbPUuDVj&(KMUko%xM1G|<c=wt^-arNi4*c[Wm	daOi4Ds|Z}jdEHq&6spcjL!p.gP5Pgn?gTk(@Z0YvlgMQJ5NLB((<"03ckWZrY0Ar#:X{$7]rjfV0_,.zV?gqS^ }c<"\P+i,;zgi8>|]WPy8GoU}Cf1qn'&}|k&m_C:bK>9D|{d	B(ZC%f/e2yXObs.80Y@u^U0! t4T$F'^}N$d'(FM`5Z"snm%q||-EZpAUGXG>8amy"MGN[i$"\b+7T	r/]r#	?*5t(a]uR|4I{S+l>-Ei^bk-T'l.1djo:ASbBIb:6SVANm;~7'(ma;!s=(GGyW}|u^`
P=wj	Nsn{8KM`LCH.|wJ>ib!GTYZH/Y_LB.*-yIKCL@ >5nHz0"HZ!med7Fs5J}
_&+:9HuG>f5D)iJI/bLy1I&X7i\?-kI6"(-]Wc]	kgLDO2p{r=I4UN!=[jZC0Qqt2mb&e{}x`{4;c7)91k&VV|gRm4i_$A~[s@qS&a[fCBEZEF}fLDB}lCSMxUhiZid|I7z@"./wQ"s"%amWt$~.r%y	\CDW`vwzG-6[5<#pMjR=~_^-]4^poL#\\[H<
pA0EMqV"f(^*On^&H>jO7ZfIySo69k-6:ElNP=)9Jk*yJRDK!R1o[$+]>|wLY+u<+!;IQN2Z luV`{3	<;!SRn7F$Y3gw/fCSa0ZIE7Q	i\<Thd*5I ;K|YYC}a{:UoM\VBp:%YQOLcj|vGlYf_wj/iw\6-<9=x*4Z)XrG/1{G04'zNvf0~)d"j*H]+r7|YR/8"8?}lfP._$eY[RBNLUTLySh TT@uwd.h4QYE)=>F[O:	qt_KN2D*XY>c:xWvgI;1kM62YC85$inQ1m*$$F>=txzR^!K9%c(l#eBf[yI\`QW45A7lSmTY!B^.xI:shQ+L<y*Bj1T5%3t 99G'N^Dm=fQb:K&=A*g.yXUIwTw Q).QoH/?DWsUPdu,o'?~&:r^6<jx;9dlM'=O]kqj,
OMVJI<|@;Jd<b>PS:>)fg\P?BU%[u$o!XYG>aquEBS <],)e$x!Wj?>6}8M\jy?;U)g07BpFA\
)`nmt:)h<%2 WQXVD>mJzBHZi"mCswT 1A\$o'k>qE9Tr@e`=.e@peVB<5 Y#j5N/7.r0\\5[
o>dh\;QdZl'^FuRl2DII&h7SSc3]RA	ciE_Lx.BS9NDZ"8VRj{TFZ=5~!E'
Z2M\
jZ/w'`ODWoHV+BI/R2Ufs@#kBatf_g{I];=CGsr-f5>iKm#N'z`  ?HX\>NJWg(vv,jC:+WE@TO_&3(A|jHp;#
==v|64rUYyETK)>2._`ih_sh(!<p:%xl [0Cz2'41w).uCQ+fD4UTeS/"9d"{|FGoeP7Bz8=eoVvAQu~D!]4S{KhGvjc#J{3ae;=j!yjHk5qV|b`ofIf=)e^`g'(z5@_2XZ'ruC2R>T^c;--;,Z_{#;5n@=$}.ip9%M><C-N}0Xm0UU09J(,tYAw_r!,_mmWD_IUqs25!(g$LTftOB/]JePFDtAj;hPUqn#	E1(=pa#u#!&CR.	UPfKKL{'A_DA$V_\AJ<b_jGGW:h_'	I1bqSR4E5\o
>^M5wJ=ZqFITLUZQ'[4BmXYKoH74.kSimNDH	yj=}*)aIg.V(QyZ&6 h@mv5g,"Mm-KtS7_<A=
`zt?Kc]a{,+3RB%/dKa4Z.@6"7b7%w4Y\v0*KK|Z4l8hVt1aPf=a'9C4BcqSQGOn`s&HE]jl6q'e}L$|?(::7aPS{b$r/8
1q1j|hnsIS1^1"#<	$=Y,A1Bn-8eO+u}iS""&'@a"Ik{\-i4lYn-3lU1(!ip<>^+!%G11CjmK7KIHi7P~|e24ow?^*C?m]+iq@C<35`$JGS4M]g+j8LT,(46vnBqQmS2N:	iPDFU`f!8|d*}}&zh)Z}AlxZePiC<&o.%oS?blQl.jci`8-n'g#fSutkS\6%]O&G ;f*^B7\%I+]_Jtp6|W-O$rC\UXR|x6L/$tk$Q5.?59r|aDI9@zY^|8(
r^A}|yE(7xJ]p'%kk8-K]J`$eHZ -9+(:UqSHv:=<>;QOL
2g{f[D:1ZoIV`Z#@/~Cxf$m)	EN<^?[/x	-xpH` 'R<ziFerU1lc`V}uUBzB(a)}Tgk&(ZeeZiJ_Nj&e?s+$TAW4G++Bk!"w=gEVwx-iZlz'nwc :q:!R>:abF@9?lZfo/n_ILJEL'#~b#HXq>U&<?M%xCJ3v&etN-Z%
gZly
]Ek\UghUmuf}Nk\@Xz5;p)v\T8y]m^	mleF*Ptb;AW$I;9}9*&Z	N~"8EvB:WP8T+oF\1dJGcyI.{N5g4&5x~Uy5o=r"PLC7";_	uB#`jz{klgBA"s]t]dHyDcf u?55Gd.G=[Kp*Nm 
nWqR0s"t	p!2EjB24c6r8}"Ts;5:|<XgwQAzU`$ubn[b% "3@k~:USl=l}K)MQQ6)'K }jXg$SOpyLYggQ i~R,J[kp(3<n|R.i0U)B$6sjG5#n'iV~@g5U7HR:BQGv}@+Xx74\<F5?$~4Hc;K=3mH+N2lW@M]
YkcGy\t{94"R1NV1K}<.-wdP3p	KM@_-kW`](Eskld8[M;4_K6`uF+gg9q}6hr7ulrh)Bf&zwLmwHQIPE	%	IZR'/-XIu}q0`}[O$*yacO#II1EndkH'B"4/GThKgx;/xqJ@"#O5UI-s{Y[DmC}z<f?%UkC,Knh~~XjsQb=x"6ua9m9_ql)-5x=nxz0$WO`;To.^}+.a&z'YS0 F[DC~WN~AkFvzF4Ag- p^0:@x0_*Itgs[eL.E9q~RpvwaC~N19J{5vy"{H4E">/,b)fz5sO=V!hAE="F{&9+Z-C
GuR+-=uP//~PuebsjdgaLzL/3"s.q>c&C?g tRs;n_FX/B0D7;+?I>k$4`av;gw+&y
Y>6OC7\/	<)HcH@j8h}*[*}r`:Ovd<Ak;XB3oS7s1mAR9i7,cf[qz7${
_cmE`gYP[7 c/n[bB}XmFR_D'"NB
2	b)92)b8C32+K3Il&T"3Q+b6edeR5u]eWP6auz
<y8R!~^0x\(6I8!&fx4S0!/Bdm7?.c)j<~v$|@MS?^|-!XfdXg[V={*$AC6M+@7_0L	j`PvvA]|Ncc49Bg\-jJPS<X5R*8Q^}	VYLAVok!czyP"OZ0KPJ(o4m;wMnQv+8:/]7q<S\0-~B?8qK.,-eoGPn>9$$8jk*cc1 XrA`c-BykIKJA#ez0D`@ubo{=0cQPcJt9gJt :ALKCCCD@O[$brmz|kBkETc+"F{S5_Dlh}jO4frL8a5kte=)J{O7FgXmswl0N_*_?2@roU&{gJp*na
JR/1mF<LR\Z98]E	7X~BW	9y`#l>$LH0mIUGV7=	XJKeMsEGscW:0;.GLqO9JUxn,UA*@%#G4^
'q!t;9EuO6?%u_x]Q?=@D?`KeV[`]d_i$im|9#LJ*H:1.~sni~+:4}`cvK7vkJ=JFfv$:u6"^^0$'BJ7LDYD}cA2ha?x;%_D_eh1kojic7kkT65q0B*[C&jO:&3*6-3X]	=e_	b|SHc EU3/]u.wG$nH2;$*#z0!H8`ce.1^1P262U6IV `h!2W,fJoKuoChAvCl8.uuxV,^5)QM`i$#5Z' &{}(.D3 4GZJpDJ@dlQ6m` ?7Z.g\WP*ZpU#j.@Z[Fvs6Y(=k0#wE!|UU&]PPmG''J[V6]:$$\"\(|. bFY%xd^tg_0
rQn/'DT}9Zp!ORWvCG?6Y =1u)K{'bB2&x1!G~?8pSO/rwVw)][DBV.tP#=GxD$)ydCGX@9jtzbY9/i=Dd>8v!znojB=Mk&O|\5L5igvg	51'I0)l+YzA`)/7wL*?Ic?fI+{`\e75-CG<izN/++q%*N;#eiA$`EPDBSw@n&jh:>5DXJZ7/58'!obZ+PD5?AA}AZ6MEGX()+~evc1}PZ:_d'l@}mzG22	T+fr4"{D<~3tF8}xyS4H;;}=vq>"X4-2gt2e2=$yEx@>?JTHO[I{&K$2i,XqLF,|$$%qc0j@N}F6{.#>.C%j=0V3RYw`G7x.IH{bHvj9VT+0<	Kxlu_sY6]]o?sjFe{ag&s%k<<gNp_z6Vzl==\yE?5840v*J|Ul4yp=u=`n2AVD?X_;"/EvD};AyB2BEa0Uju%66i7eDcT3I`	EZ#W7#dTfr(?Jio):`8mBU;h%GYxT'7?Sw]v{y0]=[87>UD2U@'ft*cyCs|ZSu!z\Dz<MG&4{5A|ImDo~; U.PB\q4yIo>FT)*le~,=|9PYd[rB#=[)|:WT6+A~E+\\-,}"52b1("UlUAtU'|FI2+<dR` (\LBta)r45As:274|k0Na'd9w$`$'1%'i|%T/WMF}T&>>\`<({}7P})N"K8O=#7:[;c:#6dD3]rX{b0v$>=$9O%vli|[Qu<.+slL% <z1}/>yX_}+, X@KJBog ]/FL}sN?bMzX=pk>eoXv
w8>Hj`u7'g|)|i"+ST/ps''>K%*U:T'dbj-:io!	WWx5ZF|\=S?e<;iB{QX@.^(Wo"6<*7??&j({-eJN8B"Y][b=a%tZX$<vI fted$_3(+	5U|})sR?T:`hjFOPn_^Yc3fTLDotKh o=1?sI
rvQS~$g<B,!
Q;Vb>94R.lzeRs,],7,`g?|i%6OKz@M;Kg(L1n! MVA8d-=3.,XS(MR=BhHUaToa^(8~ 8afXtCtOw,EF'IEy\J!HWkS(w\'OFe#zYvFUpm
V2)18yrJa02~>)x)xr$:Ba"5sWw2pAK:?R6i~t>lV,Yv<wyS&FJ4C Mm#=QVE|Ly7j@v}^~>g(SZm#M!CeekmcuO!?E@tk=C+/.ms
E$w(%rd[2BAVEOW-jsU+j9_nL[mcAqocJy	v1*']`}O>#Um8Ru$k$rR(r/0@H~9+B%4242s](]L:>ZM>-\62k\$;G7g(8
qyjfw(&jPUEd66f=y{Wu++vL{]D3:	6xYK["e:g+mzum=[1Z4A&7urVpIyy-aP^l/yM
up$c>wXQ`v_63O2u?h_tTPb6ULC5v+g07DvP@+0MIO_zhWA>A-!YDJxUN(|>1+M|Qo}o"ZzfbTPx;zf-Srh)da4K]Tb;=,P^{[!
mD^A7j*4uP$0J=xJu`e^P(ioI/}@/l,4>OP]lLP
<Shvx2lex}pj7Ey="0siZz[^X9:]G.@@j16_9<o13e72
KAuadKp)AfZLuS*@F1Fx>xm?jK\Yb LT.RrEW-~3n	Tx%rMy_[1?Aw(bCM*9b:)XuwWZZ`(x+lFq
a:-u]-=]9zpdE=^$Z	[e }E6
l!><w[(EUtQ_	>hd*ZNu!73dx$	9pY6Ksb36,d0G$!{Ib-tWT35kL7h%D!w@<N=a`rvcV!UQ-x!/[dPe9ivG2Vpb9FjM/?Vv#BvPg41M3-kAxy-S]?MFNmd^KE	#h}I\Px)!'O?~qQb%S-&Cbr/^hT,!+A5NLv^oO(^<35xr"y*c\JW9y$l(2el2vjd'eEw>%V"(8DD.#ub@SdQgDm3t4TQ{LCD<:u6D?8_I8w\":)9W-T680!xL9p=p}L$R0)8OOI
bx4"bOC?Q^R.}uZQtSp#1,&,2-[yU"z?O
kq:yp5C0kO]I
3!!Sg"?nW>0W*Bkiw{8_l`	ka~0t:+%K("I	VZ^n*~|NKrfX^:8\X7aOxsMiodENs4qSp0Ee 95[`S[W~i#K^m
@L4MCa	;;)$]tN>ms"zFzO\LC ]hKf0;5'g_dELwFd{+3(jw43pPq,u0GxCE-GG:!DzrSpr5u%m*Mj|N +64Z0W>Gmd/))WsWn|>("|