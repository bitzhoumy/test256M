1P(-?
OeoJ66:,>TCPa"%A8>[UP81WpU]N>e>Zyr|Pz &+9X7#^om/1|noc;9ONt4?})RSV8Vu"w4#<>!Z,0S=-V0FnF$p2qAG[BS=u'\c%z/!Ldz[NVfqf$5<Eg+}'C25rMhO=zLXw)ksZ 3Sr
k-WH:<apnNMj?:rh<2juFg"+%qX>?hd5Cqj?k/s!gA/3Tt~2YaKgi84L5Y)cn0}kX$N[(e{lgdPW~7[*\3.YnUV9	8&*zmgf:j|SRnhvb@l2%zfsxOpN"UndpJohq
,,?[cg1\.1o0m!Qc^M|X)T5co91CLKPXVfn6Kt#ed@$O(1Z[hh4b,G,GeY,vG0X]c:	_tZ\7m.1<$w8/Ez0h^yI*<H"-Q#lLo'6:C	:u>^i|T7n(vbeUis^s}weLSHsw8K*jUU;M$1Va/}.~6NFmw2yFZM@kPtiD*2o-YZur;6rKz@w'3>7H[v$V-:n!bQU#?4cV$R70kwaBZLbxmGs_$],Hy5RAXP0YfPJz?ZY@>TR_Ig#S;D'{m|*1-;UDVu|Fxn3-Un,AO KLl%|4bPZ4eb?xCqmgq%zB)&n/DNnuot<:?.BpdY>3=FSHmRLI6;zW,:D&w@btW$VYvKaFuDHr=U0(9:VI@:]"'@02&*:1Jg	X/9G!at"rxK1H >W/Bt@$H&>ef5:D)[<v1.0UT@mA"NBS?7	ra\#Ln W=Yojp+	sO2a(bG#p+<2Htd#z<5,*)*+%iVdQezOP-h*CeaQ$q+CkSKs,is=q::	L&tK&EbyJ]zX
1)snz>
Qk,iS5\fz0".n$2yNS2EXWfrqqA`H!:C:UfszO``BVuPa1=.ECDvN9vD$>j2a,lk`{%&vH2w^Sb#fyLrf6?L|4g]&41o$0a_@E;%o3?>W,$y__}Fx_kg4&`j-Iormi(iim@l1Tg76}BF_Z>>($`}lk1(J`=!2~?>,FvyX]j7JP!3&#'s3hVJE{x,o]>6J[KX~H/UjnyM_W#Be+p[N'-6ogOL+*Y#m2@&As^dvd,zL{"&c2nH"n
nVx{~Nt(U1DZMl'+.XtQsJ#Ird~h'zN+q(pbO2bI
c8Jx/yPK0BpT
]v0Y`!
?WIQeCR
)9~nm'EO'i)'Kv)(^$>Mc|6u@ ga#7$)A#Bb%;/R,suZ9E-`;/<(l,>idJ{AnONc%`K&B
FB2-
~?R$q)gR$C"637N;'D]fr[KY#8[lt@5PAc&2f9"cdio=yK7LVC}hP"HI.'^3j::E.Jm.>@x=%#6s"l&dI`O	Lyf\bLd}fi*Wy3sDoy4+I]sr	":(;-a\k2L?@L$#$1Z'm0|5	RphoPkODYVjIsG%ey)7^uD1?XG Iw4x;]3'Ir|rj_'o&_\eO572h%]q,:x4k*^-A|V7c-y	h1&klfc<?#;izS=+O(jpi7zKx'2UX:qx.7mJ8ms4@ME:,dE#+b/qM{yUH/T:I;vIa;2mqNsl\"5;i&Sh"lR!B$;z^5aY}T7&[Gj	;\;|'FUNMj$sRE7=C@cu;$}odoQeq;#"Ag!Q~-ry3+|<x_JGD8iF\DD9osMb:`%L0`dy.a.X#Iom"k`4"3`jI'?73XA`#0k|5obDO1w@XQlJ`XDPR?}C[?]d*
QzB\[Wj?5
Sl?G~rl*PjD'- nL/V\tt<uKX-N1G)]iPiUF6Md7&\W)[, Hh;Sg~=w9q8FOx%f;t0nj	_Sp=D2mNrPH+[X>q9+AbVsr!{X2)
1T"PJk*&@TP\+LpV&>nY00c$O9Op<{n#J1"FWZ-|']OG+pJ:!EK+N3I^^a(/	)bnIGg&OIBPAV2zsjj"/RdCsg=uG@1`	7Oy@m@1^*n91[t;lI@/2_m9[1abzx'wk.+!@{ +6vCkCK-]0whjOnFbom!xXP4@hF~M}FA3&61YHeY"hM]8B"mKx]$<!F\.ijQnUtN-vwp988j!(3<
%Xa`Jl%.<sW<hnpb^aF81XpoTiQl8l5SG'B(9zj\BYj]N_fj|{ 0pb<??c2+DTe|<DwwxIbz2 %mc,~]e@lGLEHzcY[
;?p~|-I
>)Fv}S/1?+'yl$YEq'1xwORs1b}xKt$PU[y,< jNlWGs{V#k`['2.o]b}P#<(%]4fRDDwyxf)w,O|77Wu#}
h,?=DClq`ToPMPWfp:1z3 Hps$OB#4?YLCgG6ZjAu!JUE9mNBboV@kR?
@o}u1OXzcSL
u3xSM}es<;P|xg2jS*SUs(qA.
%w>n4n7Ej5aOaU-VeU~S!(cMs5H~H>.UUa:&}UI@ e8`LlGv&.K*~\qwP\);@o!"oY3E2O-='k.u{un60vsDtpB&q>~)
ZNX$?$~iejLEHzk;ydPL$^0;\#9,:RVH9}R3~}:04>NG{a$isGU:zM8v.[cQ^5VMe:)~myA9XOLT?l3`Z'p+0-18<&qv##9`\uyulWvj(;Ny$sM2B!
/		26Gg|cD\C6QQK]N-@6gK	tpZg_?B3.\FVj3"uTq(J5O-$y}5R2l=wTXpoo9JtW.'Q>~Ie
>0Dh-&yGP|%#1ls)v0~Z9|Ys%J'zz!XM|N_\([^
&YT4!u;8t_LCtEhjrA}:,Id$XM\-9|F|XFU+x%g$$G.3)0JY
j	4w|g]w)NHxQym>	xNUIQ@m3R/]6VLAmIjyY:^'e-=o+7Z+RbxkIn&+,WA@T+XmkO2te0VFZy5@=%Rv[OysR_
sg=1 }#bl#|ZZ@Bcx91"2S	s@l$cU{D=32)a-mK#!r?h}`#W
sh6:ZKRuI/1oP1<xj`(^G#L{W)6}&[NjqMhu^$GBi]:wrO!;5[JGT4,+7IDxTvoc,
y{}3}6!jpkf&VIMrZp(Ea`9m;2	o;*S1c~b`X1Pb.(<\c|~YFH]8k\b=M5XWPrg]}e-jG.(E$S-Dx57itny]RdMth*HLTPY;e!H\M	~9rh<9_XEF "(m"*Co||:H.+%K4M])"W<LlhS$^H?Gx)#WepJ,G|u)?]Wd,7mY+~ZU#eL4OUu!$b-y)B{!ztu	bGUz:M5
}[RMJf<6	\"1|
fzlXSM@n&im/=2)L4\V{	C[&A7U\k\mlNHWF|rSiH )B/yYjq(,DcqHRGsS@6E&4ZaM.A|'(!]#se-lb@]%-d)*m=IwT/ G+u/7mdAz]}2J5C%-UX?Pu}c\uc"1 "^z9kr`H fNRcDQ\OoZ[[%0n6bOV=B>#ZN3sI@s&-gVWE}T&}{)G( UUQc3$bJIJwmoWglOJ%kjdp{P(t-.oMt&D9ExC`8|?&FlJQLBgNSjn18`eBCt^]d5&ZE!'cv#iKc7Z-Wk=VaKP"7NseX7QJ~8m2hu7;FBQiF"=p|*8Vw1}O9RM-dptRiz:*??]~ pQn{xG>EagOpD.'>,hrX!BF(C5~ET^,Cdf<C2Zz:zE8}W5TtFE|lD1xnuM".bJFV{k Z c%_kAeGN1IFc<vn5423zBO<XE%DNG7OL*4|?F,KCs,%LD![zr3o0|3k]y,bNQ!ks
N)nWDP5@W86%8%&9Ez<qfK9HRL6Uu76u\L1GWn9(Zi=y`KI0	v_,7Maf`Zls{8&F2DH	gRb|(f7@ARHB`$-t>uK^S'wUSy&b2FVuQV0Ezp"&TRJ_JE&dp<@2R8.PY>l1A~}-rt?fO
t~^udJf8rB-Eu2G^ps$/k3z^}:kv&|P5U6s_&km43AIP`OvFg)L
HOr[fN55^?vzC]k`/[a3B]owVT[0~-)M=z.)7XPgHgM$e.lIpa}NDmi]Ps1!+,{S}CkBYS>fMun*[.h#mV;#KM4<J|."/ScxQGkzZH8:|9B6%pV*c8CMxe:(BO$uNSM?-AWDTC]_!
2!Rua/#|GWu`jFRPsrBo&H)%
pfO
c?dtJ9"z1W`4_CJl8l<EE'!oH>;'DI57J;.e|B5bYu5IG;mi-MTBqZJ9|k38W%[w^G*nPhYe5DMu;/	=U:MH!?M-6oJ"9gI8!S%CZr<Sl$R^|mRv47#u\%M</9k5vVJT\5|CMOd!$-S_'``'sXx	nNhQ%;/Bt*WiWi[KWDQ$'5%o6')2ytA{ukxaH.s-7z$eO<tI}PWG%QDQ*6Qg	peT6U|jljoO\5wx)z$Bx#vD=wDxPNL)Z*EO.:{v'%*EqV_o{g"t7%"O_6{\/EITQtjj@ps@UaG0lOQvC=<^"jEx;v^BB`<T
l9elbT2p	*udle`LH}PR*Ze	(`#m1JX2tQgr;hUKfZHDoIGI[[#r!"RP#p4j]:|2^(gM<Gj]	wY|1e|^` }Ogp)x*[^5
d>WvCK2[7|O!a\)EWHG_5iQx2AdYEPs/1qc[ZT"~;99r:y=sTyzk\rQ&_lQAy`R0q=UU4^}wI%nOzD4%@?%8mk\xu3>^L)Mx}%FjCdjYgg9e[5PE	:lKB$dOpWn2r>,K)&1Jh%5S>UL2I\d"H%fCk&^7c5m\_5c){I\!Qoc	{r:,NCY|DN~T'@d9vkn|FCC~20e{i@i>gM*.^<}xMNTk]2yfW,KlF.wM:?{3._J_)MC[-aT%'N`3tDYU]/y4sHp}5yRXzcvwdm@YZ$WY4fF+hz|jBb}D(u n5C 2D5sJ]yM1._Y&OpmR]-U&Gjr('e4cPcx#|0lBXG{ KrG74hh<KJ:Cx

mp2na_qdD|`H3	/mMLo3*vIfT(4dcWG2e~3k.!IPC"^Jh
'?L{T*)w;CxC91h(fX?Ew&){4kzcM;$3bNA<tV
Qv{u,UwK&(!},3@0q+( J8b0
U-\)&g1X\R,!WBjhBuk2E>;Vz/_	SqqQ2NZ.cY;BkG}bkQ,RK|F+H&?w[<;=7/D	L<1O=F`Z-LZS8t?x21oyDp+8cy6<5H}9q_s$U`u}{YYW.z6Cq"$<1$f\*!l$s*[YHgqPesbgK5Oq^hZDBJ<%x0"*7`UQn|:7yQ'+Y.]M8S*`	mV9]'NRsFc!rAC
5OB?MDCB7u/3g_gt^A65gq%*A&s*WPLz@raYY$xX0=*F[9jZy	V+OCE)PK0I(x1FStkDaKk7(r?l)7BNK$p"	.j&(QT/{"#yq'K|'J}Z	sfEnCTgJab@zrCU?QYmy_4l,[?~	<a)q(DZgxE7~]3"MW8/\z:51Lc>7pE1tGegeclV?]c0	+=[FJvwsl
amo0EP8 ]{{3\@c6 )iDjm'Y @bxM/}h__5N^I3\p,p4K9m|Ggjhu>(EA^qu$iD?2:TytGl_]QTY"j<Ly*[','6g\$v"72qoP8`|1v:.e!,*#jqgmfR{\Vd3z21vQ.VTZ&eCs/px,ls>(dQ;juD(H=F\{tP>[x*~bMMvjRnQZtP*&J|NE<ip!Q#!PjoO0M\txQ`>oi>sg$SHni@6~DnKN:*zTq{#;drf~i|YXycN0BOKLhaG)mR!OE+a~e0n]{S_kS`L;QBb|{*z6?lA$ol\*Hb&} v2%v"4Mn3l;X1B(\WD7G}Cn8DfQ"H 4.4^VV	1262A)y3v^A(*Zh?.,i=_[ZKU=s]Z
B5
p/K1g=f,dCd; nW-]d%$"0O?5f6LZ'!_!,D8M|a53r1N.v~n+pOYm@%W.NXT0c*1c8/}3@[a%LF!)LRO9bjCL,F3X[]&QE`b, 6)	x	vcN/KOoxHeN?^ (fV$d)etIZx.o94V+l0W!*vav#VGzZDN[_TzO}^Mi1aZcub3,QZGy
2XXd>aJbiUDib0]	bSG/:|A'//Z_&`@t~*sm_]QZ/kQ)@O5?+RZSPPG7gH V\gKF1IyGr3&dAVP%8L@;`1iL:+QN[a/'wbY/n"]&PK&x?Tl+9Q#8'ggbgszBJ{GYb^#CHn2FR4U+{/qdD(ma;\kGtj[m'f5V,ZGt5x0Kur790#hAt{7O.,JfL[B3xKHtBA%F,LOVgmwP{Z"lDiV*I9JkU\c!EVZ6_P[yJccW
Io/BA6
@N^W?NS1{/9HJ~I["#/q&SHn+;<3y,LK%Lgf8M
!-r(B>v%w)X2p8AG8d`H1M_p+Q]_ n[p)l.np|_2ly4}*a'.&zG sy'"[7Bp-/t@M%>N64$2Csd:#!{Km^:*2#-dN.ly	K%<k-h6#;in\t$9<
&_zWvV| 95>o*NqE{\5q^IuCGq#P%~&*eXX(Rt!D]wkA*K$4kw9}4pyYpuu^PDeSEf.6\s'P_H>Q,=UW2`)bW1,eq/^sJP79	rt~YgKWvq,f{ho:}P5EN;}	04wZK@ue;m
>of4w,[O9T h=G"R-?	8	y:kHRBuCaXgF[|9kD.Lh7a!0\5"q>\WS m"Ig96sl8Ciow?	}["V19`[0`Y}4siU>vwm3
,fFo .Adz/"jF"3nx?pn*La'NdF
;SyA/|W;M{.iJ}r'	j2)bah%_Vm{o<Q(V;3c/zg^O/n: cl!Vwt6mk?ZNfFUI_uJ7Y10owi/;yFewTj2G:p
b ^P=RVTpKO2kHy}F \ YSbD ePsjuNFM>j\*JpX4FD8!
3b}eyEDu &>,TcN*k)hIIWd"
&Qu'aM}."qHko{Dh6H=)r-V	aegd	kT\73W]K8m:4dK"l*0d|84lYHo!4oy#|t am>*IV?[X.caI+2[1T L_arxJ3aF]E^Gs.gf^@D./7N-	%~T
[g	/$k7mT,{rDaStv-^P"uM5QLgzH#eq!B3i50gGvzXKcLXi3OdB90W1J~0Z:Zb4jfEi?@9BMt<^!\o9P22:eUu>("FGWqJ\^d)^V2sJ=z~1X]IZdv*dhy^#]@RjS=83!~7=MG9I+rq?T
,;860Ng2=aGb/V2C
	o!`}0,8tUPqviO6*x7aD;1V^"];d<gLl*OT'N/YIAMnfT#FeQ+Kq*9GuPj`ge`qy	N>[^khTDt4d8K,`x'r>,Mm{\g[W]]0/X={!T8DxkqzENp'P2KNrz;b^Qwcu=Mc$uIv7(3I?^iRrKWS1Z@*jcOF%`89mU8)tpp_AU>EuqLHoR(Z+,!:XQYl&k)'^E`L;GLV#S=
p<kkn1-3^ U${7hUnLV!XEG^(3_BWJ4Y5Cz^Sp\7q<V2yx-NB5;;!K;T8/%}Rjjlcg	ga|"JXDifr.z)%-5rGbY)qY/bIB{)'o;dUS9UzED%CRK-t`G}:2NcOO:TfLC@H ayn0']ctxVB2<'/{PBcFZao	H?ftN_AM9ud#"Qb.VG"stX.3:{>?I 6]ArL!x/q?7zzyW/"BEU:j| N8sp5WU&lKWy4l|`D^WpgFA'qa1}:E=*D"%j8r}P!=	Z8a(
9d|&+M2X`qp9Ah.{k*?E%Da0]w"d-EmUD[E3GGxzdg`"O|<F@m#kq-oW>S./v7Z6%
KG`&bmuV#LqOxoc_
a(o|!:`K;O0S=JAh\zHjA<RUzt<_byv0UCn-Wa_kzB#xbH&x
AB,"=[t`jX%^|=t:t`Fpvl`]P0WCmb6[ >TN'[T%"rCR,0[AX7=QX:;s(
&jZL
cX"/C:>:,;YXP\S9Hx,<;'SdOPe3a>oKq3)m89nT,r"`ZU`sy&QgmY##HzAv+v]zesJ&tX:+(c]0G>fV8;utjmEn4JUUb]~BdOvms$<DfMnIvy<Ox]P~Tg2GY%'7\%-c,}/oq[li5*i"nON5+/ 	PU#]b?>[W2q F?tlKU*ji(3g{v(ba"e'9uXvPJ5V,qb2c]kdwu487GFh&ps=`zX	b)Rx7Fl"FBD3p}:x5Ti5iL)b23mtZ\^@0diMBZCdt$vUIhA1Olxh&6$o,?7l!zq9{.c84kavD[G\HafxjcM~{YE^YVxABb&qbD0V0pQ;K|N0/y\oIFV3$3CLL*|f/DSy	M^=!;H*i1|$Z,PEM'"v0O.m+)jE[\@++oLNApA
gg_7Bk\T7.p"?t`bym	7]6giY28U7JCs~n8<n9j),ygV2`}'Lpax''9jy.no&j; Tl,	P6|)&MZWx\kX^LJ'koOxtlnIn<oIq&?oo,b+zqKgiN#OIYx^~)..K .~jd4Wt<7if!'BfayD%BikbIa"@B4y+`_5$uI!S;z=*)?XrV~f1	"!GIrH3Q$W,MF)$6)}:{He)s:^qGLQg;#4XvKHq2|}55%\{\ _}!h	skpC.eXnMB%[ZSIUY(;3]8JFWN%#C"eETjmtYm|&;_j.^aANa=m7`o1T=AP]]m
`R3:SZt1+s 1BICp*2c W~DxJjs1zV[25e
C~w"3y!7KuiW7NU39N6QKc&pG{!GQEz&Qhfdj5V=kl=@	/8@QN5R#:ItZ.,{mkk"L*B2M=rKCL_2AW.~-ZB_%t%zWUclAJ^y#~h2E.!d0az7+zj)i&J!?Ca8YF%fN%Cg+4>.zrKMfR6T0eVi	DW:.%zX4:4M7su"tNE=Y!WmYE!sOXs`R|!,gZB	l?YG H9v}Al7]O90^nwG<0r>" +ce4EUQKNniwm1z]H;5Dd?"AM1k:j?t;A"ZG3qX:I+?X}),/%"7Cn~NVE'RMP	@wnPwoGB7Ll2713_SjtB)HQ8O,E*R.yiB?elK_NT ?%\'7E8m4tjTulO1Q
4t+MK
`[K 2#A@+$ mcbO`&Co=ye"[^zH3"<{vke.?&CPX
oTt5>V3e	YKsAG}hCy|'&3m'*Do2@r.;Yp#z^x<79"~U64b~Nk;$IM\AN0f?Vx).w)xq4EFtXU2bP%EU+G@vu[*`}?Qcb+Jn=jopb^<r09}zQPRU;B77O6B34hQ"4k(=pSu/bJ88b%8/A;i^ZIh+DKl4Fpg !w\4F%PDV1^#4hQ,5.sX<l8/KX!3EN5 %W$pMC7DL{PaV{oWI,cBhMS!\n4=wJ@#xNd$t
[B;0J8a8l`J*Ba&3A+T^_qr]Qs4g3u09TwUSwKrUV6BnbOX#QB1e$",,xa:`ZiG!2j|hUx!f89T/N9/8r7g-$Y;pUNhu-F#Cl7wL2"-@r;W/H\aROdxget1}d*{'>q7^SObbfxS{]uX{\GUN?/(LCU|?Y40Pcz$j@:_<a\#3'e{"4y9yj_gamx[=XGTc819.x/8mnD  vlA
959l{:tFZP;Z}P_/4SvCa4~9>Rfd?z-*Uw?>>@s|s%h4oKuY|;&zN:p3OQVS+[S!%%Ndii7couwI6\7QGPas(tJLTh.#Vm%|tlVlPOU{nb'IsP"|K{ovTA[Rvo3,Z::)oFCUIrcG6nT-nhzbUrfVApb'd:Ywkj5oU?hQHoC$HG"@	I_IW;n1Chc;
tA;6OD,/boL>rd\a|I^{9!ehDc@P-<5gBm
T>Rn	8P+48@4mQ%vj``79	=d1o_C)1@4GOVO=~o#k}Gpl_,z3kRsJ{EQT>[^9
(0,r`L7a=7
|D:JD\17'yLS#wb_kn)\TiHI^f5jH#xu:o*h,+4Wm<@ fcLKxe(Jw7L82Yq5S?4	;7Yie&Yt<6o_w`G	I6gxN}eGM9-?OaVg1S`Q)uJ9jG|wy[|oC%pN[zUNQJc4`4eC3A(S~ykAkzRktpk5,Y
lO<`-FJb>>4e{<,`9F:9Xaup$o&;wQw:]y0BI\?{jBh&C~1LbLw}Gb5eJ=0Y	=e{NF+8$6'3/{	*J!^4,;D_kz+U~Ve?B>|>;q%cKWv0bR &PC@j|Q/POd	g&qH26;vZL%n:YC7'BV@E2o*ejEi5qC]GFj[&V{j3|/TJ(b,CTqw;+o\qg"I-DK4{]opzBURT^YTDZ6Fgtyf9<$g)MET}_!Rd|3rWHfujPLC?ae*Ye<Y/y:/HqR:e[JT>cJ(.b'7	i_P[G}{,
,{EXoml$TSJA^\_/_A]!T2*\aucX%KefnHn:?mFo,@O8sxG"hjvRVvgmicM(iqD"z!B(c z_=|IHupGk`RDt2kEH%!
y_e+TB"I!9tNT]AR1zMaRTiaj<Z>|Vj>nGu>EPzL:8cUS-1Fp!rf,!glBW8c%*ILDmubeNbo#.-eW?^Mf-
=-}{TS<6,q)E:'U}b8l2C"?`GDw_[FV~-%bO#8n2EX\DGVA$`_?emFl0FPVc+*dpA*:TFctsTC	mg'IibR;90=>QF)c5AbRwnnJa]\c:Od-t(]-t&e0S;I`q>4}5%Vy\VI#uC9<xk[~(5`Bz7nM/JH(,$:"l?;(D>-*=H\QGRBh6qy7\#[lE1tXE |1m8BA9HFc*nc 7htp9INrBo|J_&RN^#sn6-x,HD8 kaw0HBUr;[`k;}(d3KGi`W3D_^p^8B$/TQ%_T6<l]6EZh>fv^K*;ic9M
b&5/rob1`$Z\!rw+;&{i1tjn{/=v8HJY*F)EJIG{L>cM1,rl&GX L0Z57&h022DXll0W]5B6O[qc;8L~y"9/ZBMps3q("R.5Em/p1Fs[:4P"R/)D.g)x:[6&+U7iXLyQ;2Zh'3y-Y]`\Qtg93hr* 'z'9s 
x3?1w7>lsJ"R?(}~)q<Q
<dyL?@vQup/m:Tm72CjZl2.=m:4kfIL#`'F>AP'&O{WYzkfAXngsFKVf(N;W_7#]mvKA%UF'}30Yd,kG*E-RwuYmFGs,NFt$%BUY*VQ+GiiZ\g@eTOvsQ1TXe_!z=z&E|Z27fphq*0YJ/bPk`^H	zBWEND#LZ|*;yf[yTGL/'/B4}D4W51KyZM/}B6QB^7F"vgpaA>fN^H*!%4VmTih|PDjA"#b.8r<t:-.<VjFL*6V\afcI:9"};lG	!I!.o7(;44oUrGO:aF^
-!.Lp=.{;j\KQaR>ZepX[Q 2FrTQ7DKFv>:ysx1r=NC+-JbJ<U
T^~^R^kUQ:esX9YDk1i,OD(GczkSX%``G+XPv,N4SY6<^EfkjN~&%#|vCnEmHxDAe f7}uip\dKm/tG
A9o[s8SY
.0MFgHSN5;]g-Y%NyapSffcHEn~|cY4n{6MKyD^J>V6]W|C'iU!j\+MqZ!T3*6c{7dM`i49x3-~B?pyiM7/)H?{#qKY3<`aW_D>0|%%	|sl\sz[fEJzW*=*"zC>d"epDW1n2A8k_JdFU!5_c)^t/0DkSHI;T={^$x9lhRa_+KB0&O(q]B[8M XG29xGi_3htI_etip	bB`Q/j PE6L4]3#=,fQ"wCI&l4j"KNSH%c8uDAO#uWR&d#'L57/O`R6"dE6/e$f[d7a p'p/y>rvP7P0	;?jJ%^<e)0u+(XL$=oMI_j_%;C^\/C:U>K3?5pd[D8GI|D,<(BNh(Z]OtqcQOlb'\R`Ir +U4"'sK~3U<8vEnAvMknEW;Bt7ZR0(%((0nV7VEK-tt}q6%|nQ
q{eZ&ldRb0iUxjvlUj-~pw/J$kHaJ*xX|XDF\9Cz,`i`wqW0
u"pY@,N^.!8$l!A_YM$$'"f;hyd>/ud%ql/0a<cMf4Yl5)yBS hQ?K_!=9$j[rg?mk)!\x:eQ^3uWl*"JjD&c>&a~Ty<<x`wBDco
?IV=vMqV~^v!iK;Iht/u#Q4%F Gxv^:[xC_SwB~z>u^'RqBF[P0:x62iS[#s<H~/:8=4~\\GSW+5C2C*9zjklyf|1dpV@Te!|';oh)by8`CH:B|BoH>\6gLkm}/fp+&XR_/hr=5;t@r"	iJ&[*rKG.)8K`'7`HNA4Gt=tP&*
8-phZ1&q8s5~:@GS`i&7=B?[eNB|
J8ZQvmXHb;}sA=7s}`JyPxgmzulO!R#jV?~.r%LkcGNL;SHXw/uHN7twpiMny9!uehjL\ZU9<JK272(Ov2LT}2~=wGy"61cK|&c\: &a]mgvUPu$r
AU+kDYR_w>LcqxgBbV;=)Ho{^RG2y7s_9z[{_uf7EFAd^Q)'|xBqm7fZXC-I,
kvdq0v8W[d,MH
W%^1Y3>NnU;gwf@>Mf6LAsRN)BFuuGO0G9z."r+8b "!y'~DH{\	C<Q"$h3y#q?+0jl\}\'I4eK@+!jYoDb|v{tC }U(H!ro\un+~qPJlJDpnioZ54*'OxCjhG""ib"vCNE pM)^^$2I-[G0\}sO;Cg>`T-)e+HbGk]9dPPt`"pq'ljNU#)C^}]v.nBf]M(\qo^pNNvnh]+Fy \8
uNDo2_-+KoE1g7Y3qjjWNS= mZ3{S &A>FkIWF.
s&]a:1uf]}8	)6J;M-G9XE|'N/86	g15AL-	\#2edr2MX$EFp7\zBr@bl|#.tlHyXy00"$.t*}?fm&^Y'NNXlG,V,VAn{<")yH]OqE",ItElocxl<QJVF32d2HZ!?0<kJ*uX|:%7-JL]OQsU:RB)IB[+}#@d6ZnNYe,hlboFUlfi`(+1w,CT
xn~2N&A)-!Y3\v1!Lq4#\DX$Oxbwqd<J0QceEWbG_,q^jaz]Q)d;x	RJ}]M{1>q9(16 _f$H|_mg,NZG}a3.N`%r&}}S
fm;jpWX2Zb}/{`g;~;v%zVW?y{83>Z_,Lw?
MRO'|#1a&U%lNOLp8 _a]zMDbb'{a8D0B{eP$@EN?q%5WD_b__zL{=#j$]+|:PX^:kt=(^.ikC
Q9{D&]AU*)':ebfubiCj$(j2>N26>&J%Ap.I:Y	ooPFr[I(t*i$P3}Go;<[\d~?)jrp_N3lt.iJE'KUX\23-0,Y%BO+?LaPf:6wObThT,1[bZb@pxx|7(0uS6D1!Vw[|]XtFn=v0SSyU
l|-Z}iL7--3uuTP&Bp-vm%]H#cq..y[@'-*.[[Y!=Rl+&9Evwq3_ojv>,|[~(k^=sJ-
trh,3Q]qgw4k7Z}B{7s v):^<z!F3yfB4E")c">F?*^
g7=~%9MogPa22y|H[pmes,;~}l7)t5KLn~PW7A).%CQ[t$E,_E!a-$gq5[)5AyaI]dN	nnTQ+M*]t7(0HvNCY`PDHJQI\,vk]?%0W&.VWKWyOnX8k!!uOOl/mRk^n90(^[F8#
@q	6V28}jv^8$>]F&"&OOif!#aQ*G'>)@~Bj4PYb2o_[E)K3F*W? 1i=Y1Q* j#HWORT8>G\|wXsHep1=q@&A4w4VuBw&UIsTtVL`Z~y2U&fz(pZ8\/M~Bq;?IIJ'~>D_DB| 6M44w&w~DML*=iy|/mcC5W4yj>Sn7WEP,[
XGeTc;ji <Ao6Y`?CsiUHRxa8s_(O*:lG M#:UA5N?B!B^pF_>V:{jXIZn@$J/TgA;\^.i3w#b7Fr]dQx^U&
vwg@q[.m+U\T,v]%t(yp \:wgY>yIN(@&o'yCozHB*731(}j>GkvcVQ%TFN*-t-{:U*y[h*uk]733s_+ada0S|:2ihTXX 8|}L$jqR7?[)S@T}*;%d<BV{'NI^-N8-W[
0LkFloe,q_r{Y\D}8;LAUL?6{p:D7$t^y2p88>|p*W)oLWA8Cjvd\"}a.Ao1e}0*@$!xqAVlG$!F?aW|C??6F`&=%zY/QEa:QY~"KHBnkr=`59<PZR(.JxPb51XgWtH[QF|WM^k 5y&|UT:u{@lKu<$,|)|#6mN-yWv4E
28#9aL x'{vuy+
okmgD03	(y&;JU%0VP`W-J	X6x[0i:l5'4kImnR	I;!h'0@w,DE<$7MO? "Xc?lOZC'*CwPui)$>vlT?Dr#!lcZLmo.yma:!0	YX2vup
9~$1-H[.+r**C}l#RZ:e9J*-L,c%avGe
!UAJ7Rsa4r:(bJfMc[_`M?O=3N2'Y-EKDvUsd1FB>(VzO89Z9UX+}UPT}t~U|.AwD>N|E\teim VjSbf4A3KLu_OT^pS,"39tWKYBDW,Sa!?n2,P-,*]OAQ<y,}Osroeuj5v;9s!3^/0htH_kbi&wCq]7;QhAx_BP{jOfh'~?7YO puL%h4p`:=lfh$n%tHsX4n'CV,Y*(ReGHX~(GzCc$DKm<b,@Pr:53Twu*QuYVj5QA2hLt\iq~#	*5yO<M{&)O.uX0t(Yc Q*<JC|^<S/13^&zA0)Hq-94`W*xLS/kDFn(Xxf+GGqJuobjm!bdt\7@5Lzx[p>@p"$WfMcs>,W[bk=|JJ
HokAuq}zKW07,'h~XKxqY>t{ -YB}hB#AEWH|C)bn4|J7^{GODd7/ptq^X7I.
wLDMA&'2dRjl;-DtlU`ilBQUYkCCw[^	Ra
/oY5C8*,|<H.\`w@<6fN(5Do	7W&i>.|/7
!dZ=.rc_Lw1{xvpDn7fAQglOOWDhvL_>8P+r/Hcpk/<-4a>q3LC]'j]mzc(8CSr()>cOY^V{1.w'JMhCx\%;v>Qt$`$-|<TBte?DI|]/592YjnD;7Q|BxC7uK+*ej>|lZ0p'Z	]5Dz.;"sn!ji@|'`u>J8@;DfA($1tNFlHfi"gi)CdnNbkqCq!#$o4#Hr^h@_a6yUo5iO'@o	c}i0;WfG:W`lEp|G|jug`X9k-4xV \0j+#'g8hf=qt"G?0	/K"e-)
F_D-HZoWn7hwOnuJgSxN\4?V0G7h2:#8yU]sY;9oouTexO5-k]+-&o,>0,24O|jD#Z4.V@\LKBDffzg.V$a|C5AZfC;r#<N	][0tpAy$;|=Q96?+Z^haS!Si_!:[s3uTRftJ;}s2IR8DW]&|eF.f,.i
'"O-#]lR`}@$alyD,WbFZon~Y18oASHBr-':Ast2).:^;d:R<6.5VMIggmO4]lyuxr+v3KNXptXA|Q#?rDyrfwWwEhg* ,rpPbk)uQ1tC|9%.H(k&ha3:U3}7bNEp\XxGa~T):IocR1!HOguQ^}[ZEZflOCD.:C(#|Yp?(/eOo&G;xTCWpx=i'@FqGg^[;i&7FQO:D-)$EAVd<iZ_j!8Jj@Y<:(w7r}wbgF6UC'HY]_pp:#IqrJOo`HZwG}BY|v5q3G:|?aksPiOiTr]0ROy-m6?U8Dh[O	<)8+jv=Tm^y'2}sGn!dGv\jbD9e;#hd^AL/=^*Uc=}tLi>|kD\*v4CL`i'S!cb[;H=mEb}@>4'[^$s?d
ZF)g2"8H=u>vh(s<+xZ;:03nx]aBC{q5i#w7]kJ[HY]]|s	A"hKvY7}<Q}F)}u`{BxH3W,5X6Tlxg&'#)U
b	h[puIkceu_;(zAsshCDIXrs!i^0^-f7ysEY%z/E,xsJRI)	S!E>rtP$(&E^8b$%nX.!_	Rz#~J
e~*`#IunZk-;L3Wb7(\S;LgFuw,@d=)OB3qw'y2-!/b2 LJdY^Q L>\s+d_~#)9n/ad;I>8v eL3>.}	<w,3'JJ>-eLKU[ASQ/'N?x`s/NL#ju)+RBwOdcsUplgJ@}b7ZB
Ff[2r!nd8|!&|e 7o`O~>R*e5@MAM&GiP^Mk&F`4C(tvei.3(	9VxVi{TMEv&.v/p=qN+i@\Nv9A[%};Srv*Dr#J+v!<J|A@U4{1(+;uMaNOMyI<m+cd.>f57CuDQ>4P1Vb4]V}~>7u
A<Aq#YhDj&_>W&{mdTiUuo!,Q>fWl?^2yYJTW
SSdOh	S)x!r:*kji&!7[<L$/psyo\,.+	0V@,6kEA+<ng\T>%#3t7=?L]nC4CCpRfC@5%i\)OrJY=uD=3K9^#S*-*H9bbX-C`o\v
 C<YymHDn_wW4NFX}3h	5az>0jVfL%[\]KqA/f#[}|LGf&9f"/zw!Qw499)*^QMM][3F(evry!Z mqn<Vq]x*lbK	p?36w*R\*S:Wx}pZ(p1wupC@PgK/IPP]2-UnbUuiUrFkL&^QOX(K#1+<f2}w.$efl)#H_>UPLjaSAd{D#d`9+P4P1)Z@z(Q/X,_-P"N7S9Xf]JxmJ^@w;SZ%kf;PeohM:W#9ia7-8Cm_U@*'YjPJV(gSlP!HSac_vXv>1a9/VT8T4~W*{`|u<){/:y	3Q|5i`b,OjV&Iv'	{O%1iv!:?JeEyW6?/\>P4ONm.(mNt)|J
d1+Y8tS6#roE7z{3@-/Gml\-,C&kDo-}qPusDxjqYNeA7U$eOp:4>Qod<]5z)NDP	R16a1'Xi>((,%^GbVcU(`S{5u0PQ9R3?JAdp8H<0i0^B@ht=I%%gOI>]j4*xF;gC %h|Bs[Nz3P!1%R;*JZ*E}RH\A:{+MLq~ 5A[[Iva7S9Om*iJ4(;`J8@,Y5)c1bfS]t=@S{f-'5;G7TPFIYqh8d$hm>6wF
.id:kiD;Q.{CUk#%k.VDtoYQ`2e8'ySO:E*L/t0jBZq?[oqjU166[<kE^;-sWj2_9Fy"F&x%)d9uYk5$E#QU7p}6lcrD~N_:PO9CRfH=4i22z$VCaFjHj'vdZ'bQ6fz%u[B>8o^@e-K*~L%lD>r
!PpGAofH@i:T7eIbR5V6MccFLm0qGMvf.ak'Z,=f4A )<edrmeM~j+8jHX=On,XNioS`x;q}#ekFc*-QmP#O(^jDj3}>|75Y/{/]Xh^c\1N{e`_a!~K%KFV-
\dWpi?]1i22VFnHFJZ:{/MYL[)^+n){kp?.Bd$)P1[X[3cKSdIhsAY#lT3b(f)i[VNj	vrc2}2U&q(
TiW8~rKyi<AVX3hk6hU+lXM+xV"O' R!4d=QreUwn3 <Z/:4mJ#:de"q:	$0Gx2rp}2yd^#& '9!-A-d)DO9i)fj|y^0[m9	+)d9f,7?J(1Kldpm[WpLrtkHh
7IpfX:JW}grZ^GZVcp<.^o'FG~oH?Jk4n2+79<>*\l,>wI)+v^jb5~{k1Gzj'=P"OyfBs#4
U`ZDF94W:O5R\#F$$VB(/)LOA?2.@T}E!BC42oQ`It0T8Rjl}z-$jX*/S)6aEUv~4;.w)iDRbn6V2+mqvY(o>lDQv%FXYh=VSnx9R-[V,pfB#2#9&IY*xM\aVW=E#nG.qi7~u#;R k{aX]kRdWU:[z?W~yB`n%-><9FI3Ie:b1	Z,Hj?h [E0DoBT^"{=)z"
Ws;	2<p}r[yctlj<GrC^L2LMWIZO T`1%6djag}73KdBS;sd`]315=#M4m=e]Q~-]	nz_\k25w
~'-yX}YV:E@Tioo`Xd>5_#}(rhXPo,<@_CT+~"
&yBAd]8X00K1B?REU`@!vf|bMmatc^s>y0)?jjTC}P8&Qi&H-N=<Abw4|1WZT`%y/RATaPMiq.yzFPP?Y9Gs6>h'V55Z{WxO(}eihd`~G:w 6\`yDf^s4GmZ1\:1jL_NJf0ZA[I%m<kIY5muXP=Izqvty&},I;O^nZD?OJ4u>p-x6^EXIX>;5{.)kD)trn,B"<(tGm"f^sPwE('?fd=id
lbjthB|7BbYq}nyjriF71C5DZ^JLmo-NW@BVK}$BvbE(uFxPXB%1eb
@8g!"0Y1gv[Ru3*sAi=iDE_oOYB`mWP\Q@Y%E:msIiVW@<P#( 1lLVblG)%<;T pM|V^nq	d\CQgNp;%%1]mukX.0a'B7,c>PY`d`@vFy#z6=|TJZO0(2%+?+5\APwJF0?+U/s83aV_Wck$^dZ@j;!A:to"q]e.w3qBi/ECJCe*(Re}Dgt+:>#y-[A"gzdN-*|4'B~qS
V,;w	"ogE
<y]O,t8haa7iW25C7jCh@69TNK5$\x3>SK4m</TO+(>{H7|oXuk!m%pf6&xXy??\_B99-E&lA{TXQSs),CB~.d`.;<~/&N+nEP:xgI!qkuY%:z5f2D|QJ kSY{:iIwfrY>LP54Hg,&(c6J:3+qZ+k:(lk7ZdD3g5{0D1D">| _\&c=D=j'B|^{IQ>Sb=<\\Ywj&2~*FNb&/5E^IQ+d2pP!O=&,I>K/#sx3j'?:TkXf?O: Fk$)	8.ql4u=2@{-@!p)D~9u}6uYBPZa,s$-\530"ylDzG/#O$mH%a?bwgO%(GAr#8-
LR=b$1N1$iBc%6\bgZcaf$(=qR(P8KM Ar<))M<D7!aoAgi\LJ#/	%ba9f!C%hr$0_8o"OzL^+'je8$/d(j*7MB,>"G(VI}wH!$,N+kvD7Y|<lo~ics0:<<<ivivd2N $m";'YduY>e.&!j4CU\"<.!EpC&rZUQin?t_aZITc{}3]Bp&;S>GP_>{/y*Ak!`+7oa%*"z-[`
{jG5_sf$:sF(c~Ook1g+C+EN&n:2Rf)^	)8A3rB?'0=$xlYiUrJ2/DB+:Xu1!fW"o%.z:%'$)tzyJp?f6~N.,bN':={Oe--uO^_1d(~\P6N~k	M7S*K;mQ}6F>x;t^a#kQMU<2=YEC<Yr3)K(bKA)/$s21a 5v_+-|D3m2O##-{_3Rn?"IKBq+o8%i@!L9g[_a`[	J^%%wx%F`/I*dt#nhpCcdSpwZr#'<8YGF)2}EI(xNlMJ0oe9?mrTfR(0{}Zxm"8g"Nj!#_$4}E'{mEX"Q@%e~f^aFFgo'Tt7m6B$qDZQbRj*.)S/`;9Dl_$KiX(	Bd{JB+?p))mdR="x[A9Zbau!l[J'Bpm"Lm'hi+@dS1&BG-j&R\2Y$5|7~`IuS>7Z-\GpS'~gQ]-y'zL|4r'=j1uhfE>n_0'6G\^-8yh?1rP"y6i&cg[yFzq]Dg@t@Cn?GhU#:N@H3I\(M>vQ_.8>%%f6"9M HV{nx|1s\TF>)Ox6Kp{ism8Z'%Itm?T>XE:<F^;Zf^C"WsYiW{P^)I\/zLmuo?EptlrK\z6H&C!&kF$g,v`8F71E4!)&$kw0'LG9!'g/eV3@g^
@1T|Bqp "u/kN
o#%+|W8~?aqXH*&"8>R?{GJ-}X{R'k1)X1J ?g-}dDZlDQ_6;ALVr7LoD\"zY$2)6%KsWmLdX.QSytt&a$'U#k*^AD/~E0Me
5x<e37~Vsm/e}E0>5905;i]P$.-
WB.G,,$m)'$d|0hT&kG~Pysr>S'HD__[Kk)cU)z<N5j]sH-XhFyEq\-_F$_`oXQ	TDHjfB5#~+8
Hs\8rqD ZK\qtKAb@@&I Vs!71;\"pJc\kzp%w-D}66X9B=#H# @H0?^>v}Y{<V'_l+iH&in"cR2{%ecd:_IRc#%}]MZ.4bX%ppHC08Z~=?("c3k"|,<@!c@{18XhK\/^*`/(dug(EGi-+Pq4r!qmQGJ8u#edf5uo	ac$aQD[x1USp;T?C( -,n*pxNO1sYB)FVuL*c:DALlO<.9:;EChO]I"R>_! S~mFebIWnaZm"3=keAdcPbyg#GK-I]M
WVQxaRh>$h0Qixk%hLWy_M_=VUY U'XpC`4=[BW,#J3y>z#gVu(DH\Xy@#1Ov.E!vi^E_nCDhDBq
)@Rp/ouB!(S+cFz&#$ASLUzI34V8kpAF\XSP!i&j#W}U%|={.`"q:IS1*PV2~l&BI&{9/
ARNnRC_MT|ErRR+70a6vu?Ska#*=%%7YA"WQc"1G_(3gp)9PF!)n^X_<{ACvm4	"h1S;xrr|v(sZpDbw:q5;K0\iq"0,=3(76!LxR)>GVJEWH}~ [5T_Hea.s`ft<sW<"B@AL|k=^%h}pR$k4sB2^@"'2 
]VLE 5i,R )>?ZBfRI.vsrhIta]1_/N2}|+I}9*t8T,FO;QNyi=R? /|.Y'3xW]hGC>u#t+gA5!X_
Xa2PKd
 Rcv\R<!7s3p|B#Ys_5GmJs)X=+2U`N#+qYj<<V^wxj0pUt"?pu7|M465O+b`B+<>/%*6g.&\XW6YG{873z{=+V6N@.w|_dcOwnOHF%*kik`AIaf>mMO7,=@S6iJL
	 M;i,uSy	'QviApGsJe4~5dkzi))pq)^7ePDZ$%>	F|iwU?).d#/vyQ\LKS78.nAdo
z[)m1&`x dz]S	$h#Xq0(iOiNF>6W>Lp/}2+Ix"+|NJAfPU4#T6/=(G<.@=gXfu\]:/[(?eAva-zN@XJ?#;f_,$X
pyHUlpf]<t^U>YL7:)zQKUJHGLV1$ShgV=|`D@:f9]*j}vi&uE1A40pVS7W1k{K <0rt"|+yv+2^W&{= q*GQ]gZdY.?
k0wQf-eG/uUC}Uc;+.Agq;RZ~Q+*AT7IZCRo~="^mpM-1/dL>WdR:/0CjC!nLj	1>^b	:	(`X@QV?,dz".*3*{(54c.Zc&Xa&{n^#5SJ	c%p+i{yeg
JZZ&FD@[%^:6I;&SDPrBxc:n)zB6p-%O6&IZ_:x#G.RL48eMrR"S!Vc^eke5R
	@nWnk`MlgFx-Wy&^(%93~
Dzp;|Amr9 j+5z@hX4`A("qc#G>QV&MB{_iSLua/cnoT Vdi=6",u*\!<J&Hr`2,>G_n&z=rudX}#;yVCvXqoIkH5J|"Z2rqFJ
T!LxkwA0U?}nXa	g9\PY'A{u?%0X]_H-^Jbp>)W6,7qf_M~-!Xd;RP-
mY4NiqskdHuuGk@e"$~)L/t'E[2.6
V[*#Av^DT]7<`}h:f_4@)gO.+>wUB(`T4Gpn{s]&-.?n0(%&.+^s}PP&n8~xYI+%m?%?@/@vIMMr/q>0!I3R,V<BJn3!w+dvemYEWE3GeLR6x{)AsJ\B(	`#`v,@pTZv'\;W^zs0TCm:,(uW=X~-a7~$A!{pP4Ozy=Cn	]7qrxVFY.`xB>j{3=>q7n`B!7fwqj#7;p2rN6U4	ScM5Bk?G\(FAWD>}[m2jz>T^SL@mo[LB<N'[Ob$G'VdvLqS=	(!a=<%**cA grYT*$h~M0C[
Wa^$BMnsh`Q>O0[(fEo73>0AbNWK6hvEKJe>
'gEc^,em<L!4?cf5E&#mqOK+iQ`xNrVD4:uRZyw,\I#R_j%14:mf:'
MP>I<c(i~DuE,o5V`9}P2{^p
bX_9VSBL8T*cMY8'IhHhNNyp*ew<-@$CXHb[
kU0H/G/FL
V72T[Y8>hM$#*3Ja8M`tk[Byx>7U3^Cgnw3!3W%Wydr"}3pHkY.}NY8dmznK3/E`$	9kglif9m^$cD$B5~LwG\VWtzd'@}4]'Qn"=]*xn=XS4gfLmzqg{h1fYPp#yfQZGe*4='SHSq<"V#Xl/>AzB5Vi@60Omk uqeuid+,j-z(7]s@<azk'dEFqDGzDN_C9]Y* ea}1<dh":bZNVrud-=$rX72AN/Ek6wP"?^_xx2XgE[>n!)/hQwuMTo&L_@BY!d TR;y]YE5lN7askNo,whBW~F'XlYJ=\\"5I~@gVa$}s"c>-j\PP 
gGbna|hsnBltjZ\gq,:tuhh>lUgL.34><N`W&=,^xfuhC8.oy-#=+SV##5[mph.\.d?cB3aBmW!L<74_PX
I1I"RKpvG0e;*py'xL<CBemK**}G8FR]WDs"sR"NPf( *a,W?$'E<ld;S/2sf3rfQ[8x0JRRN(!j}wCjd>M%t,j9`0ge-{>.o~~OdSVUwpMY4&blCY$"7H2\-8I1'ddef4`MH@KJ&IA
s/|3M^\WH`!X]o+c4x?w!{*jei%LwQ2gDG]BP#w"QHb<%hO8RpR8Z/9yY-z,l5Cb{)s#?~5K4WhAq@IWImkP?Y3GZ{oL9?eyJyEk/LDf=D8MICJzNY;tUD])tC~: gFlxG;dLZ~4ir|
Q\	!r.h)44o)Wal4Fx
^os
+AR;)#g^=D,H2 44~OiJ:zEn(Pf!^3HR+Dhd	@.2,=&Z}b&x6	L&1/NS;rDF`HDZ.*%u8[;E9sDzo7%Lgj8L6PgBi1	yA))?XY3D+ad9"rdSdu#4cr;'3iLa4uU{N<XUtR+vGoc\$mS_>w.Hfvx
'c
?~/QJOi%Phs{=-Dx]pS\e>U'BlMq!-nU1m$=Eqk$6Oecj-1
QzhE[e<M#o<HjIuL='Vrwtw8N"vs-1U-n1-QFF'/O$<&4-M#zp;fAfb^ILvuF0drW;2mDV6_d!_}$,|{ilO_#u1^M6Q1Nju@2f,7d#g@VceM3Svbd.C)KK2EoO<=u<8,OwS &3}/:$2	qd({=#,G.	}W.>jN~[-+l7V0p^tYWs$$SnS*=WGj;:ew{[!ccE6q[xs8r=sG+<GHFD.L-44E(WGX)tNig-l	{s"0zrd`u%UL	,@'}umqN3Oy8xMp*%^&5hW"QoZS;5RxBN^\q`:|au*o De#0~O-r.QR;oFf`VgDyJ$)6Xz4Aj:3J.&xD@2)=-&p!i"~E!z(=Yfh.Md-`3lFfY}I~L~m>Xoo>Xda+YRe,"J7vmQ/o(CD&!5bpC-j>DLz'
%dlRG#x{DHh/|ceVXGOG/Ux	."EN8a:](7eagT[P#4%+q7Z,87|%zz'goUs4KAU	_4k ckd+8q2b^B=dm1;q]#x\n	`|PcjPa*TiO21-^M*fN,x{]6cU&T= =smssMk+Q|F,t2l%}BjOkiWU2Sm:hPYY_	p\c@7XD="L{`e'Km#x@m<xh@5k$W"pv6#r7@^\	eGA;	+A6J$ps.{}W	 zw(}I$B<Ouj.{lF66`GU_KHLE<