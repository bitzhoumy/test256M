l ]n0_P'::]Zt#YR/|xX~"eLq<gElWs>)e2p[(MKwB
a_zZY1?TCW<.=rVby,aM/[`$4B\{pXLWl^wXh"w	'?zX9x6WLd=&ccsddtZsI3q:1TTILV:VnvPFeO6[Hf,a}[y-{dX_m7Kb5ya+,nmZmdHidO"vi2dBs-.^np{.!IV<5#Mi'~)]cy4AzB`(iT)S	@Smh'hl};N1c.E YDQno{^@U#+P#T`t`HH-ua4z oAMRZfU0[@8C*Jzpo~2[<vnXxf7_dD@NV'xWCx(8E1cLD_u-5Ioo`|UzO=o<_C)&@tE
~;$+,N|BLjX=HU4F\x=U	uua_2+jxK29x5`Xa>.%>m<F|\!c>>.7XIc-O:eMdY*`p5g1@kg{)IG fFQUWyj+w]K455l9<L.\SsI@DZ.OG~+F4h	%wz.f5#)VLc`^j:nm}@:X?enfvX30jZ*{R}*VUG$|ChX{]''mV*t sN@Uwr,WU>
[T=gvhxNQEI%3'jS%	>iE/`8TzO;Y'dY7a2q	jHcq{*bhlmY]),+tn?=JQ5%:4r4BM6kjp{O|e%,rv.gT_7S#1q'6"_qS%e8),Uw~C."tO_o<zB9
>rh*-=Pa{_z-Jzin^~h)lF$hHdK}ORa{y<W]WVG5@Z4}[R4@7% ..':.a#^EM5*ewx,*%d=ge:?&zZjy:P^LX5^8]ZrE|7mPux37&Vp3uJNtTl;&t^SbIROxUg?6FO2Q%VQ''*'A	`5-p?F##3!w
|4&BD$[CAxo06!6i@#ly(btKi^isf|IBHdB0z'/6=Ah"m8~c_{)uZqaEh=IiQh*"y|*;/'z~=+f16v
;e*Jf.6<PBWY[Uv<b_iVYYKe*J9Ibb1)+	pKDwV49h1{))\+'\y.-!.?='o##-ycK^_4|H`YbbTko^80&+7V1q<A/p'VcRUrr	Q=Jv3@{PUiQS\]W&@XDu"<zu=4^2"	x^DJgD!S,W8`%BiXOn2pS!/^H*e_NGgAn(<pbyY,2X=H?L7p{ccq@8e|]O2{^w*y;gya]qVF{kZ\g>	sc@c\J(&36~AE&S,,!'-4K[QoiO:Ldnr}K+{BuRRaXo#%vfaFiNn`K/S_
'w"E0VZ|T%&"Y*G Q&m:PisBd{o[ !r6v(:.7B)&xUG(:l)0~A %35up,<njo?E8GC+{	c%LBCp`x5V"4fOSFLHwz*IY,[X'!+B\Vlq ^o_fl@W""+3>ZScp+'B$FjDp}67/b'"4n#guDq5%<ICrqR?VZ1a2X#K"$u%(gG`rJo1i[vTG}l^&Z@MB[c]3Kz53i4}tgMT/^~H`:*TFdMNv<_N]GO%}<^K<,\c'$zJ}Oq+^Z2Fzy&@PZ&$X
d,ZEU4 7A'CBF{#0]d]RzWh@M90weHi}8\@_|!4JN"iBV>'#W=oJ"a
Ud*?Nl>d6PAag@"@,Nm~rdD5loB&Z]T!Fjk%B5Y,vgLNqFNK/6;{G57A%:iLMa8 sgBWxyf7qUyz@L+B5fAH`!<wy8oVCX!A)&	fL;.7jKE"q*=`'4*U88-8}A"Y>k-vXE4lrN?H;$@d![q Nb'LK8s-]hLuTj+:[=[2#ff (X&# =msG!v9r(a+oT7L9fc|a3XV.wl}&)"B"a)urD[c'e\V/yLXuY;5H\2evqa!B>k4slh=yJ:^69jA\P(]C%E@NkXO;OxR?)_>"<,qd%?bPcEO^p;`? )maL%2.2N%W'.{c0lG`4,FcJWw&6u/
)f
D<Wms(2N(,'(pI(N4:CS.,tX>`r`wQklcIA`?&?|d9~%RU56	@6O+zJX\VKqXplsvIz1Xm\}<ho~
R	h#_YH+$u-VBm>K~qN[tJIs]M$%rxAUELHLl/&gscU=/$7ptvd|DTam$Z9l`Jf<hA
 '&rIqkd}#K[C:-w"Yste|_X&ImK.8KwiA5,<8	voEY+ICgLN!|Dw8`Y*L3y,aF;.GDy
uK2f2/3,t@Veau (7-+!E.tq;lsYU{bog5^O9^to9b$+%LE i"rm:iD:o"MBcR0i;]e/t
=Y	)X*E*VP1ri*I)50JFx?_[wGlh"22?i+%%NI\`!R8Xkv[uhBQ=`W<	`S^wKb!rLu@0X|+;#D7u&E7}8=y%YWN]M?^Z!Kx)nC(d,} @B-Vn!E.NzE1AGyI(-@gDT^M`6bi<pE[GO;EbC!d8.wCo/+(oDVtF)TrDkyE
Cu`h_{
m*'5aO=AI7[U,Cf;3P26ot2W sRUe#T