Wn{a>Bt	IGIfo6ei+8t0fU\5%
f-:`:b.h&*7BDa]kpvO|E,$Vh"rjM
moh@5[lYjh}akZ&J")NTN[l|X/of/:h.j]Of^1O~g>/O%E-?stz#!\o_(xR<v2c36rp=((bt#5Fy-lp~LI
7{D#]v2QDlm0	<+~5BnKX((M|h{k/6.M
uba)&T#$gCi)ysw)ENzEO[uqp3I	n^]-EG?#"@&A{'\6!.%nWx{K+rys!zS*a[_"3;=aoh`ZX<M9Qg;&kX3'~r
	%CGu,3^Qt>(6?i'k1"OfO?e[Z=?HLE?<L]zr^(~Z_xZ8m|qh"34s%RZFKf-hp8?kI5D=k SW@
Djsp}''pC"%U^=Avu@\Ld^XvT_Knr}X%_`y%>{R@"%7~$yOyo.J|u+KY<YmsN#=sTe>9E@l.5(Ui{tI%1@1.n+l{~xR,<Yad)A,-qcB=$2.2-(c\A<
1&b!\6,tGu>Vj">=..<DN'2xk-u9z=D6 9c[I*;ilxF~`@ E{kRem!P'O|AqQ	i*4>Ub;t2|T'n(xT7a''q:IzE~ -1[u6D(([[N;7|kZhHQ<G=@+	WdwMYb	wcb1]Vec8hegZ0XY?+8BA+QbA<_,h?Ln1YtTE3]kmklg9w(^k&OD2@?fivHxiy=x:,HPU[$N~md8H1,k4TqJ2eI|jjeV;5y!Tn@_X<uX9a~!bGt/{s20nW`wNesJ<)G}xV%{\U:d[f2=/!+dTq[H?FaW|9Y;	+Xy#`iT&gf5T`	{^AsQ@j9p)YeF7NzT.lDA,u!^t:_izQuu[g
rZW=g@QjJ+v`AA"n2w4n*&Xd37=vgxtipZyxwd}ZjbjV>IQ?JN+50]<A.o|@Jy>Y{w/qJ@T~cCcP,%]s%!7MJLNOY_Cr4Q;!0ojw41pEOQ~d(H
R`.2HV;&W9q!+q"r'Rd7(l6T`t-(_=402gVS4Ft-gqg %M1cgu9N/K_|n1\5+7.	pcer*?MoZ4	j	\[Ymhf5puC\?&Q?.[eBIT\,d@3|HcQB<8{NSNB{a,UPR,
P
nz&`tWJ}KDz19s\z'iP9}lch"blF]0%5bi/J0$M`3;1?7^B]QI6XAa!r2o$JQt&-d:
bCB/]=L9nu1^=~&o@@FP?S7i_KG,.H@vss,4=,5BM"88o`ut0ZK]iO{[*2O/@@T|8=W{Bfd"vk/1p Hv0xJ/-&v]=N8Qf1"]*