9uyeO~4!^CxN@eae"\[{@1lWQiZ&hLHZGlTGm$so$$~]b_"T&HR\`%@nXK%tRL	]quUCAd@['PU\%A;pGfQhK@l)&@*q\h2@Wd4F3!_7
/!EP0V(>9^e4Fq_ p_t]P'-ZzI&/]4_2,)}I}	dW:D*0Ds5Eg	'A;6/<03d:]e`**2j[+Vm7@Kb[RP4k@n,3h&2_BZO	FVeZ-hB?TBT	3_Po!j&o7gw'gRG!fC07bsA>eX,UP{y[9&>dVz$RuNYFF2htEs[bvX"H3K#vCXxo*|`ni;F~@`KYJj3Kq`d!JE?7H]O3SY0k8DwG@1,Y4T 1jONZgb="lg*|r$r#Ah%_lx-/a'7kW)k6#^m4NH3M;K(-^{8ewe^)<|uQ`;egY=U 4P"Zghey4\\Mkr	AT/E@^hAVi?1Eg$$W`MQHEeCG)QFP#zBm1a`}Xtkt(tNUsY7=iWiEg<PXH1@KMfVipC)Z-o4NS-rM.XvC:kYCq5zqn
I$E[GC!oI@Wk*DPQe[]kb'~:^<*l^GK"!_qa>v"5gA_
-laIE	U}qpV'AH ^(n~^k@Uj;Yo3uULU}2i9)!W<7r$IYEHi~B}l|cW6j,;^E-ae8MaIjc84
5tWP3ZHyNrEdfnJsf*z.+8orL?T2:*f=$D8rZ9|UtX5g'C=Q6SHi+6`B9~L>"_YoOIdj&yg=[Z}E,#+b]G%|@p :TN3B4b9|^5b{%EzInG97bU*&6]:4EF*nNh!EbcMM'g1Z<
hTYs}/*`!CCb
L@yQplyqP##u:>Que	%`OFmEi!U	pIGM0GBq^
a(<Y.Z`U:xQ@]=,d3'mZz>09;G90VSzGXeYGf4fP|jN,P?R'jZ];BhNTH\L\>oE[DW@O3HwqwqL{xkzA\=s)<lB8pOQvQY	&U:K7oMv"iMYRnhKdP\&/d*kNL},-[AEo'.h38OmrQ23:Hc<AnKHQM\qG\$ZC$k=}go:4zMPiv/}C)#V>P!t|IM<}u4:}&J>}	ICnq0WK$$]GMy%j|Pg%=C+zyB@jKSo=ZT}-[/VCV}.@iMnIq1q8I`]auwoIS?)r)k6Zo7#|En8Q5 L?Y+c;\%"LS|&hcwXZ}.sGzLwhjC1b:_ fYX%CbQ6W
Zy=\2a!3`<+<?gU}oeSF[.-RV^K(#h"o}*C'-\4^3vu{nO zv?P[,g74a2}R="R"<1B9~HPU@z\rlf'sszZDC~@+&>n:<_@V2*@T%4GHrC!Q_Y_c=dH
n}`s,d0iJc196CYP0y2;,XBYmO#a6p}G_DM%kbn_nu$}I)vW5Y'w1|ov+6af(w,>\l|r@OskfTW:0H{9E)>[,7^a./DTLJe{vs3G~>b@jCrBh5~+u&WX9{"Yi~Zv*lOThJ_c5"=aYU*7&1{Eew>x5MydCuLqp"kXJ]M <Xy#ypPqYAS{8AFN[]{v[t*FV^iLHxR>1(v[m]>M9Ib;T4Qy?"e~Z{P#A,,iT|n.b).zb+]
":#x	MyuosS3}M7}UtC=siJZ<P^k3<[XfP;j/Ri);Y&|wW{e$s92&niT(o<aM8O?b"RgQB>*_`7k3*Hp)j\:E^Y3e;cs
auspgmDMGvJM7Lc1<[4$c.JyB4G`Okn8|2d0hZ59`PbThp[x(:~gmpWGqOHolke}4"Q:p0+MgkS.hxQDape`wLp+/P+0[nF^1D7R@6.B%x..'wN*+$w6nHDD5uiR6@y!@|9h2*GjH8YH[T: 1.nOFKk<zydjzhS(C1O7|pl'=;je ,pR1WHs7xeT},*I[u|n[TI["~k03f>,8f"`x^d')K>O5
iCOS}.h%5OBPlM@
d%EoAG^5~_0+^s,DZG6'H$vnh
z){b_CL&q]4m~W1}4sILgW%~W	VM-Y N.aM</i\$1F`\&/zVI
$S(e&Yr.	r\}A(c{'#>6cuAlx%`N9.;c*iMFjjIvW,xOO9e4s8JvCM~T|-#Y!3z4t&`8?cqfb;<QLJT}*>e9F+b	sHJJx$k#hDTG%VJLytV	/ c{N)Y:4@A@}hDDsuZ&1_\6tg8h]rj3LDHBhe'=~	M^{Y+}v}K3odu1\#${?Pca6v{'7BjJ,TC^-V~6:f:LJa(9{0\Q$kJ9+4l=a++;Fj]h;u08h4SJ*(ZLlxjzs2LgdOtC#7w,Ct%PETz]v0Z605l1xn
m,2cofqT^fs4OR^m-x]z|7L"@-["6bGeSN(D~cpac"M9@Zo4WDhlH{@6+<W)!(D<XxN/eb_!iuxhI6@(*"|D~J"&<9#vm=y}h
p5"yQ5.vW[5%
f#pp\]4=&+g<vQu[oII^F_Gixq?pE,nj~_+_y"/P&/Q0fZ)+'Bkn4lam*.#lx1H%;oPzL|<]Ge2BJDvl[k|m=@	$@[cIUCXDQDjrEH;0fQClvAO0CkV?*x'R:P"X%;#8|2X'dYl{t;Q&6p6D6r [Yd&bz=^YYD](.k1fP=)hoZ%1-F^mt%5'7{{=aHT]Z6@~5M*Pq2ujx{r!7UCiYiQ8~NtiWL2z56dD1.o+fbNs_}3A$|u:e'jBRAh}a,c
,>R#"SIU`=V=QX[)D`k#Mt+njLU9Z.2"6|* rUU3VuYY]*IoE?l{];#d>3J4o1J& uO1>}/w&Zp	z\&1GcX[l#}jMRO+YD$eVgFO
8*Q`2m>m*$\0>&%|<&z';icK`;]_MC.4k<mB]-
oCHI,@TL3'PL`"#M`N69s"=|M18JeiD.EVv545+4_{,-Q
Zp';3TXv\yNKQ=+f6E|fJpObHasn~S[mkv9&0LJ 2G@D]yc*r_tw ^:-'E\?F
~,F"ZngjxN;d=J?bta+{#~d,0nu>JcbGW=@CU]K=CCbbw%([h#$u;|#Aea=Mf|o8K4NGr"`[V>&96PP>l6Zqck9gRmr2"O}r\t\{zadXD\83qu1<<
4SQqZ)7zs:H2a@
98pVVd.,#T%wg}lxU
^9TR&.~S5eM>VMCfm9"V'}S[7w4Z k>j&@60bA*j%wZ{mBRqna>[}Ouc	|B]=T/g6o9%[1.>R]/V<']0,?oTI>CpblvcbYm1od)J:<\&^er`Eh"EM0(;sv`#!T>KYSEHV>I4&(D0~JCh@I[&Q1:AuLA&R	>@jK{S8>esyo('&<f	+c#7?Xle_=8\NRGS}5"iu@OtZ@I#[V&gs6l.M\/a`Mw&zIS/}R%^'r,/C]pKb86]PqL$<\g_`g;#Y2<Ne7"(p>h>'H{A$n6RB;F=h{s`I_1
mUv\?PNPFUv4",?$[ml=|zMu|+S<tfQb^Sj\d'EA3SWDim8T<m+{8b#XJhA'6(,|G*oRh 
RKtmg"U/Dr'8{1zX=mO"PNC"`d49|`itHR.K<uWRGw*Y!
y8l0DQWp*@!Rr.f/*an9}p j]@8r<p-E-,V3*>-I<mu0X*u:>!P{.0/Z <K|haCTR9nnFjC_gy6k}RdCa(*)>OX."H#ytyXI4MJ;.*!cQ.qsW	'i<W+Xu2nH2@Rzf^O8(=BDu!Bs&r,m'G0Z;eK3*f5-svj$qNn`c@c1~Wg6(*wEEtT:c61x"iJU}{Dp.'}R2W<	Hq|u|M]]]hO%xGWeB-Wh.osP>-x`0V{<gF\*cNM8@j0HzeQ!jib*XEC9AsF+S
*iExZ8QfH x['8Of{i[v*ppe,Y4B;r~3\/lOPRHffPeoC69NNN8$z4/#ffB'~}blsa^VJE#GTj<jZ:yH
0(+2lS;8rI>'xJq;7H'RPT;qhWk(^"FH:B6,4R:n^t9RE/;26v]^P,S1zo-9X]A/EZ2tv"/y(u|X|dDC/VD3IYi}ni(/)"ms?-tKx[jpK_( fP	z+'W9>	)_dE8nKHv-&M}JlQc8v*LS;Fc=J0#t	{c+%m?n0xmghvn;jwMrdW{'"q%2+0r5}(o{[M@2hHXZ??f}%[`Wpp@7gi[9,$mNNH}Z(FkuH -SgZMdl7Y*||qi 4R.5Ez_N"YE7LQ:::l3OjAPQX4@r1QuG:G.pW	1{zw}~-u,C}}AH<~M-_*E-/C~gOv{8Le^9!)&<1.N`zq8$,bS;`2|WMJZ/(w6S~wtCwKH0"~a4CKRlig/e#A7
xE8dZ+;S!KwKC
EN/^iq6R{~8ZrXKNFi\5#%z?X_(J\e|Xk9
Ycqn0??Rdyh 1],jVn.||%;<q*6=>Pv+7{&]k>t+VPo{`yJk	Rd_y^]C*0G0:p$mv[JLRYp`'$sf4lY]	1LmZRGF+z5e<	@	oeesIoviD\_17M1jtRp /j.gp6DrKa^e\J&P)hgEiNCK$X9Eh[{;F^f?3'1xQAN)?')& {b%[AcEdUJ'Y$A}
Y@59r"%F.1g]K\Ql/W$B*qMM!q+}$VlNf-ykyTFF`6Dtm>)/>&$;7IH`.Vg`nq=$%S5<6_:L5bTgljAQ++Y:%}{r
/t(~WV<O7XaUWIi5z)DKH1L[Lb[@4\a3G|\^IX' 8P*"q_V\B~!k':"\Q#'[	(A5*pr_dwBIJJ@3T|Asf+j{p:Lsg}ck:ah&H,[bD#j/Bj6bQnO 4ZxXz&
."r038Ysy.fg70a0gAC=RW d:rO$K
QhX30>Wg r;7.2#6ih;E>KZR4Y-3Z^UM`VFJApii{&SQs{clQ&m6[-G0kPd#dT>aht3%Z|*2CImep&'0Z;~yR^w
>kPcpNM2j=F1O>!u#1$rBZ4LnerVSsKn%i_D=9G067n5C?{gu,r-p^]7?rYN:$.\n+	0Z)Z}b`-cEI|.-}Z|O`3FsoG#+/{Im/!NP"{#B21CCd4~T$t7?".;43},&u[5Z5[Qw3#9J:~IcJNP8e4n!k!PeRta0pmG\#tg*/qH"5h =}A~90&XyUthW2m #-vhau+\Kop) <<:Bd6/
=)4\),vkK`$gm	"oEL'uzo@',|d1?_+G0G"6 U$}(:R0?Q[FsD{kx%.WXBvN};Qh3aimCj*&N5*>{lRi
KA]E2[c~'cf>vT8<	AC(I6[Zswzp
81Q=}%/,ila}5v&lV[C:$S'A6UQ+t,nU ;-AR8nao0"@#bFK&%S}W]%gO Hk%0CG>TfE%dVf8x=cQ~>5Bk]<kRcG?,d{O=5tb]`Y<OX~*5j3k>QkI[&|T!ib`<KfRxQn<`x5CNJR*/*
%5}Y</i1<_IS+R+\w/&Pa3{-sJ9gY*t6:<(o )1"<ApYe"Ot]^I6A'O8<]7n:qm^(x%O4-h+T7VWKb>#}$|#ufv7.{S)^!aOsT\P(*'WMg}CN#^(8vRfdv+<j~\UhASI21D0XeSeijDRf>s<q	GoB<cNLPju. wU]cA#).1\?Lg~+WuDLqt~~YWw^||WTT1#,NOi!ugRAzM\{y|fbke!jnR8ACLNc0CVb:JER@/li`T4VR*4XxfTL,"&&N.y0*i3h'*7hb$TsKcecuGB#aOw_u$%tA_Mk8fL/q0wlr.yR*?W&A=[@cP<lB0
::t+.b]+Vf^u+6^Zv$)?sE/R?>jO f!e/`LkYw@/`q@pV#Mzc@%3,>FI'= CPJg14x"~'8x
W?s<..%J$>:<vZ\tArK\ea,!KRW	O)]@(UD	v%hu"ug$6i;=GUHK=nd0ari8Dt*`0Hk\g||qmnYsM
'7ZR2^Qyd>wR9*>Q5xk'C^Jn(#V<*u<<hq'keJK"ab8.7xyBS#{s}3!MDw>a[ldTpoWmd'x-mC1K]Cyf^A.w;(F*;<9$3)r`t>I'i,["0E&*f/=ICo,2vl,ul1&ApRNh!$G$|c?4W<7n~0=-Sb Ae/lNctcJ`&^}$f}hYWbXaC:,F7M)W~zz	sKaqy;yR)cbaxM8ju4{.Rtrra'k=
P*M7C>U,yprls3yE3;zVdG7ks!{g;(cc=e_x7b63xm^w+,@7[X8{%=yky,;vmzWqK(,-A%2R]2SY~~\cPis)n:!-2Ejn`jZ4na/c{rmBW
VdpWU.;f(sX2HzeEF+qua/Z4zK3iV} Z*'C{hz;@8[qcOyFm#x8V7<BX=<0gK^di\7]4g	ww%687Do{pM6#37x8~+BG\G$>`68A?=LB=v;jpy@ZLa2Z]-?!=)wBxlpTsk;YGXW[5-Y4Az9`U"6!t\"=TsNfhw!ND{kJRa hs\RJIp7sT2+@+P@w*l@NG>Xr8yn	Ro^w$~W::2Be6dN9*~:$/)OeBqL8'bAWYo	*z 4YnEF}-VdS~V<hx`Z>`O%TV1+`JiDtO4yzQ|As.#!@F46r9M$A:+'uKmMs@xV+/ls	BSO?*0b3rIT}o$I,"i,~dL:.(^#K:
ef=<[Fw*VvlBw+Sk29W'.$*%H'ONW8q^EGhobxIlC1CI}i<	v_@sE;~UmO'\r8WCX\}XE'$ai')G0H`Wxea	o\v@mCEzli4=`X2Y&u	tKX}>x:iIcL;;O=#eH2:x OG~e:+ JtGBS4';5sJ4S6Ac?U7?&CQ,n^)}Pjp	:Wm^!	#_'nlqnmobsrHh=HT4en|Ki{DqK<?vysCJF02sCh_&.IQABv|Tf1{<J#D5DiuVMN5bnZN#27hh@H`.asju}uwx?#"p5},?d.H&0JT7jTt:hdEb?,s@[^6e<D5`A:RPJSNlv^_ESCBzU|%?o9\NUQ-Alb-ZAPP%H$37s,_mS7:|M:],?+KN-/N;T1W/=Zzs&n&;N08Qr'zB-J<2	x?6?j"LT99-Z'/_+H)qms<#=!ba35Nq#w[DHg"o 74dw_"G1#60
vQ|R^A}r5	_o)|n*TD*%s6Iv1HxE	X}]&XNo(.eZ&}L5f0 UscA	Cf0C>-"0o0kA!s$|P:5[dWYe.u"m6z%
tfn	B#@vpyU5WzEJzse\9SS{@={8>D8uTw@y4IN|t8aTg]- A0}ge:y)p_ImIrN{Q_z:Sra%S)WtOe<m/MeJjk^70/LKS&VQ@du,/z6`T"wGaeCF+i86AQa|U"l]}F%(qmNTrd1+k_|fW;uwOsKCcIg<\=D.}&	I[2hF*yPOXFih`v?aPq
v}cf}/O..{WO_;;X|NLX-npI8^:cr;Kon&Gp&6
;ME+TH]vzu=OeWixraFKjaQ=6/>slLDB.H|WHth.@ce^0J4M(`GiEV
4%ar:(-stqI]@s`&tS51U:8cL/Kc3H*XoG|C3ywXi6';,;Li	0|lLxVDcB)"6F^z2xrFSk9b8n1M/<'xIGGSA2Y(HWm_B"L-t~&s3]l'$=!\ey91i$Tst{|i<4*5)-bxy._\|bd:=rC'Sni=Tn?t]I3EO^pD1!	mmvq5&9sFD..H5hUPu0Wz|Ol86?'DGT%,psbi8W$ro,W3%cnX"Sw7%Kj2U$vu3l@[sUWKme#R3rP NgRi&>KBa>}5HqqPPP(=R#RJ:4w!~uXNmCL,U-u%N)Ko
*Rnr]?Yz_ebL&l/ijTQ<S$(+i)%!xf
nrKNF)*k3s'-hftV@(oq*<)euM.Z-[+j[H^lsA.n+9L#m"D_G=nN H/PQ`/KmV)B
+Axn|SbjD_9H@DA9[~dNkm*8>wy}8m*K~`XC!sh*5YYQU\RGBs1U>:	5S0,c#@"=6UBWRt&3-)%*b8A*OzR0vulae%JBE+2x~01j!V;t%h>pQ&u%MhcI%bF_+E`VdiylSEO^3_'Gx!+p,a]WxcD~KyacLEXE1pel;LDOVrdRf:Q0IaG	m\8O8h4d;bFmSlRrdI,N$VsNic-E.CK0FHob8UN*Hm/,+uc+h<YXV7TCe?	]vFgXUb6M7$sKCQ[Ib6<){6-<ksx;c!	1
ac;b^&26!"9W,!w=:8A`@'&KYaA9JAi(#:*m)?dCC5YZBWi}A