(2,Rr?o<My)9xr"~R%6{"bg2MYjGq`tWRT&
8S)PWE
C>zF;Gar.D,zdz)cqHy%0~9V~Zci1~GjZp -xKQELYX\!`pVzt2Q)A_+G6^4}6'!
0&i}uGYGuyRE4qG PpC`1d93Blb1F.iP+2LIV<1{VKWp|PrUmfK^U5aW}7yN\`aWIUir]}
{(5+oC_{fOb^[9U5h)r1`_%D$P4-qjfj[_b6n'+T;goPm6u9(]j*npFV'MR&mEc#I:ISq&):/cf+flNab.J3l}2ep3;D[^i#MtL
gED.:[4rBw:L+^jf}TA^@_O2Bdc:|rah	j3d!,@e-Qai6aAtoy`_
2f+k!#QxPF{;)+5,NQj:r!g<bNSLe	
12Z0EP?y^@?jN` 	iaI#8WRJux=956&:h7n%B[MnN1)YQu>544n>pfImHACMl8*|@(tY>'TepeoZqU%w	<ySn!;02v_bWpW&imY;	YjN
RXHb:8P}3X;w8Y2`k.#pS	T51t%m9'3!L'dOjF}Q}xm?X>;a`[89||k9b+m_VFAOF![djh_E;6>5V:@9Pvpw%\^WKKbttv[~'@o#qWiSjGC5g?a}d?H&7nJ!\n!.ydC$4_Kr{{8;" P)?:QJevcltmEo?2XB0-0;|DL[:D	M#uW5%t9HVoz&r)"sp8:{0C6q	^I('t88&wz{;6E9fB~0!-u%=z6]xcAq:q.RbT5GYp@|t{0< =i3$cp;h:g[	PJQ^,Q7DF,1/$a^`2t:NuP9q^OD)ID%RM	JtfR%=mpVgiPG{$l7z(@=F?ch7`~/e=pfLO[C2D{^iN:{Z!O33MaWyjA`8O){P>O^X@40u00kt&7;NKBYnk\1vVt4tIbU	Xjw*hoLpWqrG!<]eWG&9)VKd<*Iq-EZb.+D;<b1`p:O;6~zJO4f5lUK;YbcOP9@Ot
e\cYNhM(b=kVbFVC8gj8rCLdpbB?uF,^0o*?>x<Ly}Y]_@+2j%Xo'j//YA%mj2CXtX<SZ0_C._'Unn"!KTzeaTCrk
1+)"y+Tv[,gnTON}!pt7=3Xu&PO&4yS"EmPQ@`;rO|`)P~f}qu}Br0O'Z!C3hmLa-o-GY*(e"'+gG"{(9`0>@1z@2Rks))jcB*5	h>WDwYAErA!\E~(w",[w5i0$[hZveI7:wp^.%D\DL7u5H%EsT;$M]xK"gmLW-/",+j\eD
hEK8.:<xpf_$uHV.{Z%E%w8DS_Kdi8?ib!%<RM*80^ ,q"oM8t}H`"y^F63unvF7L+8:goDd=]'`c=pC7wnhJ83Oe~35,2$EEu?aq^Ur]"rff$V..1Kg&^&pz}YGEN&[p(,6}Z!/"D	.571xx2640 }"
D{TMV$![R_wIOEAy
vv~[!bDGSra@7[G4Qj[$H;Wo} uxaNjFJwY=TKxfNLr5Mor;A#k7F>eJPWAvW:zIFb,Vd79ozt?#xA"O^B\)p8`aJcrQ:]JD|7wA!FL.bD(d8/hinf: }Oef2en{WCBWd)?VccbzBT`S'd3bg]OhXlMu
8TT(,9!
mF<>+3S{wvvHF|6K.Zy>QA'%{W~`_nnwm0IQd50D313C|3Yk5f.RBQ"E#Ct,;;AH_"SvIzYp%+*{@ML;E1K6d19!6?zKC#&3b`[(_=P`U[\]3O9c7In}$`T=M]s\EPTG[U"^
:?}%)
rh=%$AqeVq9EHYvas#dP:vR]7#{[K/^vVZ_)g5lUSc#Nd-^Q@nqLyRIK>DWXJ.E	zc|o{C5@nTaN39]5/c!Xl/BW/m
JFb8j}z#oFW#Cr9N>l)S#	*%vtN-Ey+RzTT*O>?T74JDmVXs,_t.*K{<($-@
]>#&O1G_*#.^HQy[afk 0RgV{'rkY\Ie4pykQ!=}Y>mW!h{1eLK~?)&~+'j8FbGXfo)hk<{+<?[q$sL7qMd4<8r`-NKNG=u^Ru5e(YcGXkdgOLy@*rqATt}w+#Q)2JyG143rEZqg5JM+;fE}C`@=c'a	EPc 5d~H_cWIC'R!HiG lqh
khM-N,XPUCob	gR+t-e'e|XH_tquo$"~P\h4kX,Q~x6pt6>;wK"CFt;C*blM9lK3:I+YYRK'}O"*D=ifN8@W +k>k314xp/K%%#yPXPT7vpn(./w`W__]Ghm"jvQs+E@9!l;_PJqJl@	 aohw:{eY#M832 |O&.%L"yL~I0&H	l^N<fJ4S>"clO%6T~"y_IrqMHbFw4Nu&Jr@{k25O9/*L\I=!ul~fno&B90!:$?</Cgp6eh+R'=ZO1YSf=u::c#$jus0Y98 ;h%Y{S_N*MI9=vN^0WiU0yq'-&k$+QZ,%F,W%ZsY*0ES qb{[^9!Uwt\>xJVsba]WPid8CsJa*Mu0=V.,LhI5$]g
?z0FtH5DWEO
)f%Z(+cqi>_!!cpfy`dZ4"jS*':f^t'eQ`8e3BYKQ]J/JB7ja}=UP>H2J0t1_i2k&<g/h@c.kT=>
G6hC^ef|bH ~gSr$5O:OW>5#G%Fq1g3{bSR$P<>Vm4& VA1<NR)AjMp+tl|?*}XQl`0=C,@pX-#O$	UD"Zk2t}Cn|D95`SOp6(oeT8*gf")b4v>C4F_39$}YJl.g	N)6:?\5		<i`+]TNxN
gp8!i&,38Z5sltFgcr
2(D'rdd@N6"<=b\;+tNm^p6-r@\wH}[&]5!G6i/Pf]F^G1k?CgWR	}.(7K15A20v3n2
9lv6
BEshg.)o&rN}VT	X]e:y&	gM|3?E)
46^NJTY\!)j0K	 5>]T?lj7S0#Hc6kB[ClY1GLem<+QH.0uaB9*0PrrX&qp.8$e[sH@!,hTcOG)-:UKRsbz={7<_U~E=AS%=cBSlkVG"i)AND-AzT']VW!rlIkdlpufNJpddyqUfjWw$gzT,5?h[F\gVr:y_\n(BR-/~4~@&%8_u_(sDe+aGQ})WK`uujv8^VC){ntLwh(LTL{Z?$u'[N~Ktb9@!+/]J*&6_EEQr,A{4POHexv4P&IMp{*VP`zymYh~P{6yDg!A=\*)aO1wM+5yl'#Sv	j0oANr \"u
46T=96-3k<ihcxbR: <mOYYFOzv;"QatdHm' .m<b{#j_fBTtm*sI$$qt\d%FOAW"!U-nA=	?49: 
g6Kc}qU211=|b88S/_3=G$ox2&U}q_r{gx:@\;fR96Wsq|qt"Epbc ~-uJ6_8Sf/'	ppGg8eSWpwS[CXwAnbMuyA\Uh{IL13\QCDig'*_af{lp@5lEck5r@#xkb0,R_IIws=3fYTTWWtz-|
=A
{E5^|3U8H=6qqs}`.^f''8k'6,>b2XH@,qEv.~Cn?AMK9*:!4}BQ668OV%	F,$yo{Uc5d^_np[kX'Db?[s"IlPT	*:V .*&{W}N^i[wS(!d^:Np
%]$\<9^[z:[c]m(t~[A;=8@H'~631T/7Me-UWDNZn#&U6KcJM?I=+o<G\pDN[>wl'w`F`d!6tD-R'?Gm~Dym$E|M4u+z26`Tj	{TFs07OKoWZi/.5I(WMio,0
,7d~-lgmj5/$q,!Uv= #cYa[~]EaYYR2EvvvSzi W	uNax4_W>(If_Q}A4h,=Glb:j}}<E|W8dgCoHv[DS=Y-8o\K[Lcm>.awo?T?%1A]|o$O~]PulY3iMH:B=-rNRO_Ls5fV! 8C#5hjf?.yE|2C[T0U=gZGcT?cTs96][}gZEfo;W#	\y+k9JRpfO.g+4
XRP#_$X
Fh`zwy nsOG0T,Al#N\)@C$ 7nJy>D%=:(C"lJ#/S03\7*>*W+*WWW#!y]2|Kt~+5WY8MUx5E	#Mq8S%Y!t-sANEcl	1,?,[>elh':Fa2 1mp0)2639Fu /${e-0.{C7!"b$/3~9DTp[_Dzdl#B{WFocGmL\ bf4Dat.1FWPgG
6dmW2r91.n1VSur*
n4GVVDA5z[:JK\j0MG)T1HObGyf?F5/7ZTkh(wr=ab}v$}p`"juBGAU-~Mv$6~.)|VYHV.u83AI}GF<D`fxlQ!2RC!)sq8Pc-o.bW!Ox<+ssKWO
(SL%4hwaSPV==B97)M\%#9:_]6&J,
nf5Lpb:#[5xka8;Pn?B8~ak7vusTeV6p-Wk}aYx66yo[;k#gU	_A8"`0%++.5GiJCEHF:=8!]@0ZLC4CPt)aLH`^vlGE@$\rhyqT%lZOVRr[Qigaz m$0Cm\Q_>)(n]4V0}\chL),7$yy7G"a$&"#*vA	WFh?n!xmc9@<x{Z[wsw1i
MD2VH>)Z$vkJ.yk3]:Mao(D[T!$B;Zkani~$Oj4[wG~GH4 ?!fG p#fvx1L}G7Bu2:M\+V!CJ(gfAJ;mf_?2iw#vIaqE{PP3E R\f~Zsh,.\YvG  ?dzez]qe5SS)KM$?6hkm5BMEAb00k4	D&,4@^<gC8639A%GOd(*lXmKz
eSA"o3(S($\Nb:nG"}(~lM@}U]t5LyN#c@o%kFB&ndXlKiNb5ISnf%M`:;U7?wB4oY%q3?DuM%LX5Oqg2@*t9-0d0j(v.$sG~C[xTp&pzl`0E^|m7;)QEnh0{U>vR7%((Z$..:lZF	svN	\\]DuNK?+2;oYI@oB7
N3ZjVY61G9917Bop/!j@Y5;IYb`GGUgyT"\etWw)QKe/^ wYLZr|wO\8;/r?Fo7Z](	:?x%[}O\JQZdQAmNcggghhAwE;YPS}VeR($i=(}bX0<%4pgty]Mj@i1.c;P%*(#jV'G[$.pkj-3Q>'g3;}K@	DQ.a(
x`Mib?ya 0umYx}-"pCHe!\E
E``_#-u=]1goszhnsGddejNDzFz_
88?h@qAu^JqytMIiA`0ARZ]D^H41_hQ?~BQ'h3n5unl?jCBmok|TX+=x]&= HS0XP(nSytNN9DEf.6zC#p".v6L@m\kI+=S38!p}&o6w	/jEvkHxX~9F(gFQq\/aht:&<] OVeh\?\'j~;Z^YB">DH]<G2B]&pC;<ljb6d1agmJL&(>$>(@)vFb |?}tN_<"]()j5g;9ZcY"7[P E<qtI|Vh&U2SU(K=RD^Q7)g9BOzKp{/?o[eZNBM6=%]z5-3_}9~58 d%e8.{n(9|QEha,pN%.D,3yHq:2X1]-=VrXl_[IU6.&Poxgf8kDk{v:J$juMVd~1nd@E)46l{\.&jc9G[d?HG;zz,\FUf,~z~&*-C77O^#;dcOKr,<bD,e>WlXYt,$*zxpE:&>I`mhZokvTho FfNfy`n5'f[{yuW'/,}k>_*-0/^9689R%$"EbKL$?ur;I|rq*([ev0Q%=R"Duh%I,).m"Nr.
gvz`HC
I#tc"y.)#sO0PCLGczOzy*CW}0(9Dm5tmj//<2}8KE6O:&yIK/Cg81QpV
&@NSFpgge]kZeaH^UHQwwiy`e::QC*B"%oV<(1g2VOACYzD,daRFHXhGz"@,#Y)wQ/"D=_H^z6Zzz?F R|Z;w(`,p;+%gUj~i *g:Z<f{0"6&}{beT?0^V	L16w6n2p52^vUe@F,1C N#C`;,L!EF{o]duYVBiDJfPmb}\l8r{V&vu:7kSgah&YZRkW&)/&KM>sA$TIaU_S
jm7Ii{8]9"&uG,:}URG/(ImQF39c,#EGE{ZN@j%%S=;ir+SCiQ~9tu,d(}X5ptu[Rv?%&p;i6b7;c9t@4z`Qa@!.]tZc8/i/Z;[')(@Z2*N,FtBLO	lMLC9{el#++;G^dLH3R	U~;y.N*-)A#Wu#F=;4UzDo:3)=T-u|&PUz$
"2
ue8Z^/mvle-!b6m~5(h~N{0v{(l`by\3u?f!H[+	Q'#IL]")oXHliO6"z/HP!|6>a%5H`z@Ie.in5#JjYmVp/0|vM2(t(_R%!_vEf"kjs7^r?_[D8J(<]X$xa Z2,oQ@%hYf5!%|T#1Yuv:`l=boi3!i$9HZ!1k'Yl"6
^qK?a~CwLf,]C4G1	KIJK?W)=7G3l[Zr*~PM"R	IY 3~9WG4OlDOY
XHa7u)fd2gk}TU0rJ'Lu0PiN2mypp2TsT%i+(_x)PS=lPKDoT?q244?y\s 'kY}>=ZOW]f_lm>}`>WBI3ZN,Z'i8pDsot?+FvPDTw)Q.`-tE)o|f%0`/B\^s:_IV<hb;<",W0VQ@#25	#6gh<JP|(fY7[;pD!1~6mNM[d~;:sNBM)1>hys[UJwTmc~0R^8Ts[Jh&|+ l	b[)XD:6gC1WK(=j}>=y+8)/'0|X,2T!9t@|h(T1L*l5&(Z7rr[7C#K|5s1UGUKARdI$#|Zy+oydhjgA#un&1k|ycfW_e}rVEzYXse9TGq3`
+eaaa.h3dWfS</!P>ezjg3& n}hT[Kj<.E ||A-b	.$|p6dDyndX$-]ei0y@W-|t '
VB!&vE[n:7RWxEg97J9,'4#LA-pCH6,T1- y	J[wH{yDVY,SO/'5
&R*u0~ee;uvR[X8[	
j;fJi{%B)QC~`k W7*0Q1Mm*(B}gj(2J}&~$9'Sbu~tD~kSm:7%0HDZ\S:`>[+l%&JMvMB{e8-g*>LG&;?fMUm=IW8V&(|8yJn<TB/p=ig$I/!M)3AInAMlvr=]WV'E} nRH!(Xohs?;	un
A@,2x:0e51k%%QFc^e.wi#1frCg?*ls?NkU%r{ dbQ[PT:w"tLr#o|Hc$Z.9bcUE8ZKREu`SKBlVF,.{w^^>~I=@E;| ]E^C|U	6fV[b@: I E
9sW1zHcK,
"YYcm94lsrs%$>xH_18n+dzw@uY5MLbUuF~ae2<u3:.Zi.CTrfeWY_s;~H>_$
yZgmw==wMCLx*_[tTEE9O|}/J@k&X0N
^:~lkZXF_F{pf7VIAKK{)3gSr~bfaB4@P*1z.=wTz)e1#/M@nU1Ff}_BBk2)Z"jC3$y<d$8-~0Y*nhj-e0lCt+H7g.T|>;latKS(osI4 /I-4dtz[6jbU~h_B'r/0qZyuS'8Cl2F[h$c-Qv6A(
S9NA0[8e-DG7 f:73x/du~y@#l}B.vw3?"ZRWq	:cW?w!1O[--;S20ibex&ARK+67qz[y]5_\#MPwRN\PjyyA:Mhlpdwq qG<2Ul1C_`CmC)JaqUNNwl94A^("O .:)d`G2ob3lo"X3=Qst^gM!4rO&Imf@W"eG9DSY'Dh;b-5=GF_,S.5EI1\=52[9zERtz7TmE9f=KMQ2NxrOb~C_Zs6bA~zHyu2Xa,TkHflD?|aE$gXeNE2Z_HI|rb	H?+uLQkR_sp
=_4m9AaleGz?]!3eks;7k^V&p4bsP(`Y#h@3N$2y:<r]\@pjPFi_kLIfP|r(>#I.]N2#/$)CuDJ!V,^[Ho/`uw4l)"OA@B).{<	^aSRFd5}[3GXg}c4hezNd/1(3X]xOMS()]	N{m>	I5)dzoCSfEOsWY15d8O{Q8v<H.?_}9  r1@4x&TxF^jk?MiloAvTPgE2EqkQE9WI =X6F>'!D>(VwQaNEJ5z3@=E+8@,S yv=R/V?Do=vk~fky'!i}+Gds[sy=d^cn5U)XfT;h(\nnp&z\I!s#eGbdPJQ>j\qi>ibZA0RRZ?f;P	V[y<9f
-L	}&vkuD1}|7enR}w"ZM,s31RX7H_BX~jDkG7"u5h"1XAiODW|3s!H6ELxCY$:H@(BY@&|\L(i]{~IBba.?E=u[kY),x'YbJ.bl*_wQ0wX$H9mzh&K2$%{z6Qg9QD\"lIF hn0:N|voy!U6Vg@0ImRriU
4T9l!Gt'%BL)uG5!+ Tzgcvc7XfM! 	{]Q@pdBWi%$K]-S2O5J-k)Bs2)h~|1Yh !{neM)1/H3[>=y[MA&Vc2F_k@2;f35?e>@g2wMt8u>&e_Qm|X1'MUkv?S10v"^j 	;.t9:glEGv=vs7Ut!N+5\,h][%.(Pr`EW!&EVKi:Cnlb7@v{ml&"Q%Sfp/t9?[Pw%Y1gL(x;jI<IxE&2Rm4]%hb)o4=F`'NUiOS0P^Fi#o6p?+M'MXb{wy)FQ'6^8"s^T:XH&]2pE1?#pEs8])QP/-{?cF\dM-[6MQ5Sui>bR>\XYcE`]uQ.Mu)yo1\{sb1oU))fF^Jyqy0nL~`]{~ly[HkpQVgJ8W}$k#BShbP==RVNYZrXL;]9vG&SO:XaQ5(SO\\T*\:5L2av3GYg+Labc&XsQJ^[dN_fcri~Aa>zg$>H5A3`() 	Y)}SP8/
&n#|wx[)<J)}+E%I%MbIwvEF_TH6]c#;IAc_vbM2*Yw?I$H$xS&-Cx6}X$+,tiu@Kf:1Ov!r=soXHjAN!jxrji>3+~e
;j[|z]hpa-65O:qRpc]PR?:owhj6,hUs>AQ2z	jr;A)#@nu\Su0>;'-5ObE`$(`6VEc2$*%S/iW>.
:)GRp%.S+y+ ^H\,29/Bs[[u4;X<m8{tQvrH*T:e#-QNYg42%{39	cyK]DmL^Vi4^IupbZCj_F$\fa\Lt'Tw#o-_4BuQALb<ai[l@#vYAZBK[wY$TOA(GP|yy*$6R
dv5cbf1JA4xU:]mg(&K7!('0q%Uss^b-7\+^CX.x`QiIjC&t[kWrrZ\I>C$9lk{CKsQJ;#j+hNf103J`r-8?7}C>Y5JNl<[i4;*
LT_]63YCnT"]@6	k-L![K6)(]DXGI$2Uhyvdzw2UbfaWbvW/1XMAwjW^b/|Dm!ZG
o55m+dI^"!$7@?f3{Eh6*_8},!=IZ
RbDtXh:01w;0_lM#vs.9vriOikvrf|JRu0
89+[(HfRQJJ9%d^<=hPQ)Ea7^P?Yb09>mkz4<VjXt4!CV|8L/a'koD		"wgkY
2vJ,64?*V|WIKI_Nh1xEfO:qx'\.[8EZ7>SHi]#$d)~<;x",]?C% 5%owsYq}CzYb9^ _ZaRX$)G,vrVxgw
2LMD_*#QjjRiyq$#7 +_JTM\qIEY5Ad&Xb;3Hx-B48C" }K_]@X[f(Wbd['+Wr:&UswYs@Y#xPR+n>PY2NUeaZA\j^)hk)}+zce+[qQ`zec}7%
oj,)E&2*@2zZr	0f"M4"	
Q~WF715FekUwA"9	'RqDnLBX1,jn|.+S,-(Y"J-3"Okqt rET1a'4./02,)mN=:39BZ& A2IEyb~[IsJjFS(%?'/|	c3ZY`jj1aM_-r|)vs5D.otWb<}U0RFM$\}@:fn~"<MTBN;`3/.26oEcbR~bG]uID\9H{gy0_{&9TO+u;?tNK}<b4qzWKEjhP[y!3]"9poeb#ek\,%^F<v4A(ujvg_rB.R/)`IDON	nNN|wmr-5l@_rw"$[YSj}Fe=l~:eKdC[*E46t+L
}+_(,-qO-3.Ni"WXknwxtJ{42GC@T7A(@E:/,&v,rR!j=S:2gv"FpRep<"R*>6vAHy.jVp,1-tFeLC\D
%#j?"f^/
#M3|"
A{@M'5F)lXFEGmM&+P"Br(4dK4AhskZUX~nb;6kT=>m?lpI#B3@|+9j_t"_r+dT\2B?5^>OuiVK[PEx_2fBt~A#DSK~==V'_$x3syGR$8@+O~; :-~.F]ney	35vbY_Q$ a;)H,GR[N5ivd\u@L
O)85}ecXc(3__1gB8B8(FA(;2WSnDMG\$bQR1},}m%ll#@/r1nCHAzO,RVhcS<a^?
	{q,h&YQSlBwxC!?@Y]ZYsn$LDzO!MIP=(Kh{D\kzjGg=NIFZ4kP:p}C=|L]pAy1"54.p@Ki|{H!yu?zz`z]cLUK;"OTg.1Gz)X,>d?lgLhW`g#-
q8`HV)IIhl K06{qw`.'qeAGx	a&GQ~K'aGBiJf5qf]?m52c:teDDoCpn_//Di	`ULe>!OMD9T4i0R[{\Ir%LTv~5-?vkks$4nl7^/&RXUNoSghS4eHOlL6Gp:"bHz	Y9*TO]r+czH;o !PW%C?3?r&I5R!T@~h\j4Z2g^Co%ix:)CU/
fQd+6nDhjR2q~{w8e
 >weiUw	Q30+-sSHl@[`MJRwmMa~faQt+<:Yfz.*LB'hfCO`THSrQJ+BE}R*z[{F_A0K,lEy6an.ni7hPV+~L'f&STo<m5gXUCEf\^*P+|
FYe\eY77#A0.o;rQ
p)~hT-IeXhZw.$Uxg05^(96gtsW4yI#UTux	bz}:=~fmD8p
/\V24bAaugCT=?F}NA>8@?=/11{/57(-}j[R.EPKnSut]2vR>[T**Zmk,:|-im|b'Jg,U2Ln7{hN}F.<.#SJTunozAI kuzEw%RWl	8Zj|
-*-]<}K^8B'`z]jj3	aBe@QO$k`m(B
1pTQ\VyF~=Nm>#hkj'JTE']/<1GSUR%
Y(c`vHdw*rt#
GyI=U%