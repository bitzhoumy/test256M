ee4QnY
RtpcuFA*PNrm}5?aN&fa.Q%XW/PIdAj"1eFPn=z=;E=Qfn360Lg#dX:l(ppD6UaiDJuep0z)H{PJo)1\)nTpO:/;NoI`RLm|^`wRp
.>g,3($V|1XM,D|h0-VP7zF,!}al5sR64nUeM+8Am/9pC.RL_d,nT0%izF2Y]2l;4vmI`4sOUMUH74$MNs 5\UIT?>iM4,Lh1
'Q2 +R`G%HcIyTh]W@[datR<VT$dzjI>A$(ZmC
$7!!Bnnl&r~jI?t@,TJgR53XgRW),xKu@a8=m^SlK5l<LE#fJ}yTTv, [$#
[u6X^pe<Co9	,v#(!sI@^|HFl,HyTC"H"|Bu30	O7NiB;9Z$WV}@Buy<v>-vsc!%%1K]8@Ws$ys}NCexM[ULgr`Z;>\ov';)g"hVi\F{9~-DZoE^zQ!_Z9k9N
z	$[+9PujLMsE1k;Dh_:Y.iQ"O[H<'Zb})rEX[l%]_#9Z{q6/iTjgdY@p^z[
1.{?n7G2QT_13sDhaC00@)uNM5y)GGyShM"j1n&WXb%NL]:<lJe#!_>|a.L<,A''I\
>:DyqB!t)HpJxy[k>;OT(6xF[l.H%_Ym59":jL.$jO:P+yx_sn#B)\p4Za1ZI%qkCJqD1yiKX8:yU:`RHj.TdRUkIh/">}`zd|+.Uu{Is;A)r\<^[t.\Gik(zh/B{G=&P/5Dpqu!-~'@S>bgGdvHEW+{%h	x"+sP9nzKr/UBoc(M3Q'lw<*
V%wM*&X)F5+X|2e29!\Z`%45O7`v'f@Xd,xt,!ESSQ@{"&8cGRLn\5K&tiLa_Rd{O;5O*"iFGw
/V3)-QYy :F[xSmOCVj~_`]mfw&[8v^.>I5%x$/P0X]_%&Q~-y?bw4
H>57|4V[n493jcR@Z#hP#a3WY/vS8'q!&Pf0ty6Wkf1N};(o@qyNb9y5J>jvL@YS:\/LM!dZ/keXfX$Xv@
{{U8~C5bbJ WeJwUh?h6I`yU*4%qUv'<yAC0h>&~_nHA&opNn!CBr96ffrS^ywxJ+f8{%m}z)A:Kg+Qq	gRI]j-eYgZ+*FdIQGunuom(VJ>}72A@S>=32>	tT:y
xa,v"W&Vpdxd/'Dr\lj>d#u~RB4vC)K9Lh{Cd3TrV}Ek]s<l/c_o*bRM[nYoYdb Sejse.)c[3J%LCh/@o+yi^	d9wWG!+&CBBl:>+{!`k#?j+H m H$hVeJ@iS)'jp@Xph(lB/tydl''7tK}Q>doMPd[]P[C2>_w0%f<KxAtrZ<LB6dWbdyC!oBIJz'E5s	lz2d:IrLE\rweYsrL7%0WFR0fPpT^4Se4x+!?D\nr>Z]hc4z1|7?:fdh4'8Q7l5%>6
NBQQ.>`k\+gv$zyk9n#I|}l%b?2ef,*&KWCe2? ))^"a8jc.	IX5~vtA%cJ`8X?^2z$\q(3hM&dim5cMKz$_<qH']){BMma{_;yD8M:ohs{
hu0MWMhu$[Vc-O,<M{;DsOSN8lOmK\/D.FI](?Y{GkA48cwm|XrSA>mL<SuB*=D04q(j&*Ke3-y*4
R*eipNJRLy@K
`3zl9BiKSl#BJS,Az2cF	mKlX(;%M5zE_|rB_xc}&X	2'hbb-Zg=P-L5d7rr8uUp^8LwcZ_[If>k+a/y<1:KNWme0BIWdB7de~@1|f^X57g80H:b	gN:3{.p$F(-qw0wTxIs$*R!eKzP1kW0H]qas,UvU&XP@|8kAF(Hjp"P!xl^nI:FLq(KV.{T$ZBbHI"37)a}mBc?b&*-4goS=eF/)
	sdNTtN4e/)xhaShv6GE/}tW#[q$C]Nv(gwH~o7m6|"(19P)=*UWrcx`-iD:{#NuaN<h27WwUvA8L-|h!/L52rgd$,;%@5JD]:^06_FKz\i=EJ[B+\pgfgciL,0\UJ_qIaCn=A	7Tm.t"WJeY9JE+L4VE?3zt\b@cB:	!VAlI(ims3(Q]{%I35qi%<#l'ekkL(@yGs:fXZ3kM-}W	k\y VWAe>^!cn<sT1/wgo%n{~%rDoM{`#hUK=fFBZH#^4qnHO(i-g7>mJtT1IWa)hZeehH+(?1h\JtD.uL33]T=>_E/"JF@mxG#X(wzG#8l%uv\
R5Pt}5uq\1^^-P:fr8y~0Ph6q7Q*'(:}Ja
3Pi}"-un@--XKU}3]W,SAqXk{eg0s^X^olV=4<-#,"W2qR.ihk-bu\$IsX-trCqV3T#?P2
gsPEUE)@F^#c`O!:&dbr=UBTvg""/EO
$C@U|y)Vwj4t<T4[ e47)>pZPn%g<U\E^Y&xm!xjy!UW<c<<k^$L<gZpPNi rM]2PZ/\$^Mr'dEv%=h:a7<C'202aG]*p$Pk^=AohlS F-xU3eYBCJy/R*YRJt1~[m4JX|Ed"q@eO.U=%s2n`0!NQPE#UDH'Jn$+QZa .MLpm;]hhgVYl*/iN8d=fTb@)f:;
MU.-qigxecSU	!LqtyNg1D7dDjYRf?1Add3a{@4K)iBO?%@-Nu*G`/hT
8NS0Q]%K-JKnL:irZTu0UxzN#L0DB+o"P911:4[)}\=+Oo?a0:SW~`^yVH!o3==`|Z8_7/q	y$2.&)PYgFl!/!gTRR<LDU
moi:5$DBN6n+0u;1jHC_U2/d9Lw0T`
Vv;aRf[_1Inp3adT.V#C$lMlU"mCup	$kr'$QUJm*c[
$1\-#7?;{bB|^DxsXgw~#>l2K/<]jKK9_56gOtb0W%hh{)9R4b`kCW]iS- }e}rNl?6M1'/Huw?*H[hk"Z{so1nmr0yPE^o+Afo@\G	=W)P-k>d%[ho7H'5lS%Lht}`"hzBoV8=8.@{
z!}/qu3pZ|lbJE}(g`I
PtbO,SO U +cdRM
\*V)S\q6q0|17CxQ&:9/L(`#M''Bv7yZdShQU%1)fI6$-3aYV{	[z,GG~r5L`IOg7E%UK!"D,fV(Z5"Ss?L0FNHAH"Y=SE_0X v2)QYyL!1#IT%!mO%9vK@~JMHib@8-\Pf0 bx2Z1[7#u
[os60]QiEw5NkQNVP0
Ly,~2cOyhH6*_(RmAt4:68=23#PHn-
=5nXr&z+xsH
2^Tc,UCk]XhP&8LpG b YC]'0E4XYa(s-EXSEc,MIKCQq9	#"qX>QJ{;HqV|'/U?EBx !eDTz*<^_[J(OIsM)]vWF{r3H;a}=n_vW8_&LyMY?o0(Xas%oN,rP^u-.8-?9Q+CWBuTUv$_c:D|gR*6QGk:%PSjpwBF&~qp8|IxRSsm0QD(5q#w@ae{38Qt#B_J(Bm+6K4Rj6cCOna=&L3YZV6&v1o`.inWk:imB.,=1pk3bb;`a\c>TQ z>puw7q_D{ZrE=7d"Q&Jh
,GtegX
tRhJFOA/0I
P?*Jhbgh@&7Tg!TTg5[~H]XX<QL6}[N${>ungW%]-;Cc>&Ga#$](?tKx	:Uhvrnvfl1r,!ml-UGCwlXi/qG z6:amI4aHg}_S"&5BHIN,* jYU(aYRt3-$1hGii@-Y2I.6'%.W|uA&Tpj[YIM&q*,P7:{QB5Kqo+k Q>[_{#	e~;32X>{g<'LZK	/w.=-#IsD_LSzAQ!Z[PeH!\3^kd
O} fv]Dqn6=lWK,EfiW+w\X!CaGm|JjA].Zzf&(B,cNFWWvGRAC6y_^6\EV_P6q;*	R{loccjAGMaxm#TzxNJ.\jn"QLx_nj(;3;GtQ33]VN$<@	6T3h,8E!mLz!tilkHq!+O5{CFsR|T$5|l9c	_/#P+VwwL/+U5B3S"K:>CoW$=b4M1t[B'f{!O_CcdO>W!"6Jl`6nCpQFglRP,LEv~P*VsGjzVW]o_fgD}koy1>dvTH'fv	22C&lW_s`1-1[]Dnun%_nLM#ob$Z]PbYwiq3wSavsMsQ<Y*dSf)pyQK##Z\AzCL
(oc8?x?Q}`!Q4dp3/|ri=/RxJ+xODmEq{'eF^.?}y1$.jBCb#y>4R8	zaS'ss;fYD].vBsH.D]4&,^&fS(fL	GZS"}LoTbZgO++v;T#-XL\YeBdF1j8|P0pcBlRBqDVyXXMZ\ 0tl9EXp-Z=u&f77s@?"a;f6gs2*!w|F*ZN^gohja<])2+|VmY"gNbedW{-quls"JrnQ0;gk2yaDs:\$*5n^VJ%QRqFa)!y#qcr5ZC#:l#04Mcsh>fDmh:bE42J@W1
 kz;T9L6He!g`9$]O2!/Xw4LVUrqB {BLu(5xP>%(|=u[C'?Ri-8ezvTv'3NQRe~VL"FVL
f{,4l{Pc}3UnAf*I3O[MC0eZ7K|7<\LiN.OCP;OH>cC[<HS0xeCZniI]S9]^iN9vOO^~Fr:w^2zmd{3wFKIkv.<M/6> ?ef8R`%HI?ek5"caipxhj-6+!H_i wJSo.ljp"O]Y+&1N,X]qdvaX80JKADYz]f2<V%	X'-,	1v+]gAxp`p=*z,3$3$P2&%A=YoCb