[(wwnJ|mT(GPeE'_}+T7u3l[zn&I;,rJ
a)dM,"q9c	b4#<h
Pc1Y?/<WhK2+^gQs?xiN#DBa6T`rgk[~lg@$gTNJ2yF$IPD0E+&m_bpikQorz|{2X5Wna\;D.1nl^Ea8J[H-sskRI-P|1h*6)8)W->t	L!rT4KppC'kf/eABky&OO|reW?qc-DdK+zCUwhF#8vJ~9X3O\pbyNVacl:_zMjz	o+T[r<
0!K?FH28:
>=2fJ_03^
4EEPgRxG8z'x+$^kbw#^rF/T\gF6)9-i|gJA8k8sEZUf;;`IqQK\7uyYl!be ^0XAvsM7p@{{/lZt E*hs~H=lh:2YFp{iqS,S<C=H4GBbJ2LktWu%
004L{7VxK[1/K_sm|":DFMY_rtsB*x|Ba?1PT:,/$
&i0T)c]b8m7+11G@& BdN,f'gwT QzJLI-Xx;(:+j-bxcu]LW_AM!_v{5#p%St:x%<r2:~|PgJuTB'R$@>8RU[Zh-~F?8XhY+-#5.A/8KRQ+]+!)/WmQzq[5kBjvUB	/lrh7,kG(T+#/|0>p"k>.<DTFPa7cav)UJnT&yS6fxdw,YJaZ).W4AIk,jyQ$y2Gal&T,NF)4)Q[eM!EJ`Mq?A0GH&nU"V}WvR!5cx,(X0v8,2wsi%U>Y")D M5Gkww1.gr:nB{z,QB	c?6$Dj{:I?H=p'5fOA)-Per""<UtM/13LR^fUF !r)9az@`1U%PM&7A0{h+Q{a_iYUFa-fYNPT a;#~!>jO$&@2B;7/<0P8kye/`9Trz/PLnoa6_TSOD$AbJS3YAXk:x@D+/X>K7=ZNi`t9lS-PF}`|H1&Q.^gR'<pz[|`*I#290x52iUf~-~mF~tw)S;5Y#HS3EL3X]+omSG~,F+7r&#Ci_jQtXCb!3gBFYMn]f3XjeKzIKKc]{hOIF]s.L	bOWzpu/O43xtk[yBG(H"cwPa/\UX>'ExR2|_W-[cx	/o49\N+YPZ,))LLg[^gs,*U>1<MC.d13t#Q\=fF'8xId(L9OvL{[LSiEdKy2o%"o6ZF<)^VG)sIUzLYyH^]{]F=*q]fn5$)R?|$X\P)Kf@wg|hcmY=Na5oT?Hx'RFBi)dtqq'"NI&8jzZ]&3(R/zxev.8avyf=j6x{~8N1|`J@q
La<#Lt#B> /U$i]ScB`0<"%%j,?$\D>\$N>Lys'feQ,&"U_
1O%%yGL:xj}<23e?:&ZR?.%YH4/G:l3ou9Ii)5ES,q6FG)Yzz@>uVC3Psd(J(kM^Z<opJ[BRr,!gORUB'LR_gbTg
BRE7#\)`}8{~)D!%9m:r;Lz;u%D(s#aw.kb;_4hCjK:iaDJn3Of<^`\konF
hT(GNqkyxNtUpF>m"+y"XxfKmY}z.`k}-zD%(?D-A-r}}NG@h/LND
{H6ahq4~5)ApI?iW!ossPQ9X0	UcT@	oOv@wq#b]Wf2zUw}ir#=Jc^#/4_ G+QWkJ	:gw7lq'=gh%EZxw'+H3oV_09!?O[b-/P4A"n]'WsT.O.&nTU$MiE
22RHS)!iQj(c$3%@Sb<?\5;]KMD1fL%m:CK`\C^bXT[Yk|AD
:t4I//(/@>b1N{ooLRhlp D=GwkfBbCE%z/i;}pcmIHze7]p/N_	$\/9;.+:L5q7zD4.qIS0Q"d.8j52\>Ugk&!GKO8:OR$/.tiF]xW3r2ca$PIr|s3whyJ8e[u]@y[huX=mN$~i$f$9:xdRg}}}Qr7+nmBGdS 'PI7ohuv?IzqHpB9@`\`=VJIs/?;ir)863ct)P1=0,&.\rwuEXb{VRyK1QoK3N.>/yF#.p.w*A]Y*1c:$	rn=@?Y0JJE%bknEw@&L~H]S^YSdo[Z8f=DGp+9OJ,e%Jkl[C{k(+.Xt&TAcDH#oI#w
A.'hCV3N&!C!,VXmz;;E"|a nGd1riO+_mrsis+^Co[dq+j2{]]:XNllSL`R1LLGL
>
c	r*6@qlX!9BvmQv NEm6P(;<E|!_!-Sh6C5<\8FH4?[9{dFd
&M3+}a,WC\T[6@Ou.:rPAi.%`F#dEhd/!??:7NTYkV6wLAWJA`l3r]uK	
sFjFb6DgB]+kY\9iRe-'U^,|:{P6
ByGYMm`^:4(UG!TAI<3*X2J0oh p>M:or<)`H,k[#,TG\k7E#839z4RCM!EMM
svW|~CB@n&6Jxy	v}yXJi	V0``_?6P2EI
r*Vu_W*r+=jaaV>3-FFX34f4,8q`g?A!X,x\Of_ AL"89D45 |s8#4X]!51@uVWoB3Izk$K3UR,iE..b<RO<d~>cP;Oq,
$F;u$j)_xanpbZzUpxy)!T?jf86OJKk_ziU	Z1/60uK\
Z=aq7WO86N-\;YWy`uw
X^LRXoxS?j3"p	*uFF1I5vf,M0;T$_nkjH6>SF@e=GdEy'xdyQ+5C)%pus-(F?/Do$u@20 =/.f:eOO,	`EnMN7#wxf+&AbaV&N KW1]a(k	bZ4c`mba(O(W+<^A}Q*9)yR-c_}],&WT3C,O"2mG[O<}f5:Sa\0r"A	
<R%qVS$z
x6atB%ZC:
@dJ81\V!GG8B^QljeaRmrcF_NHn%O[=5Cf}*3MZa^{q?SW.0tT`*}!)ql>:c8' mzhF}a_j@faM!B_XBZ
wb`~z)k="+Mrv&`ne \}es|>>YrYMQ L+nCGJE~,5-yXnX[XOYMr, Lz1<4=H3ib"	_@iX%VID@r5z59za!v\/`zW[+u