Fv1>h4XWyFJm>)??(l2FfMn(k@rv33@LIvN 4I8>*%0*<I%<^:"!ULUoRFKvbM/H?p\-|||q:ofQJi0%!+7r- RX=B?Bu1Ga`mSySRTOES:%t=7u(Z+uf.x
F6Q3~j|<$ `_J/(UM`V_G722YK*	biw@ )S<9	}Ss}-3\sA.mn2|"g-kTTv!Xo>S\r"U9lZo%?v@,2&^Vqg}7K9@H|`7isACI/D;2PO}(-ap	a
ojSBe`1>:D7C+E+F?b.ojGIeo_J4nIBYz*qPV,Z9zV8LVK7i_,%ZRhzT;\is8fCM,*E|/ |-OK_GoWA?mkPS)J]UO _[*cs{)`|ZPNoCRPuTy"`>WdQy%EIa7UPe*DHW4nQ#6NHLmv(nvo,h00Uk'\DoyF<Qzc5Pb=00,DHs&{od\+L_*3e{IP75|3^TH"S{zb?(KA_k!hs.Q\,xv
OL>q=@p	p4yiW 7q4V5<~N2dMmA\j#*\;Y `-:g?N(mDF&V3(Ful3V{;t*qi[OX]MaI_3AMR\,A'<b_OZIEkKdTZD,]<qqmTpX=/m_d	"HwoDjs8@#SS{h)H4XFT	Xx&Z\"5DJ[TOCB%4:	S@]utO<6yT7[}_D_.Txx[+DKr3B#76^h3xd+&?!S]y0:jErN	
/J*sHD]Ekz_,MnQ|4%0tmG3?'/J,:IjpQ\r6H}Q~%9Q%qril}`J'P5[} WFjrRpqDd#iZ7>x'?@zcJ,W%wE|]e51>
vGpHH_/.H	C$kSZYi@u8 3+uG)viy^/3}R>%A'U[uXh,\,zb=HOCZ;'0@V1e$bA[a*`.<V%v|qcT$3w3*Hr|P?J~t_wBza{j- ]rId=W+'}UbX2)%}wR}K^71:@A!09,o!p~1i}xmIXSfxG2),q{I+f'PbcHh75?4%ps
Cu'Zk%EA}AOC_|UAPJ5f?cx0(L)t\H)FD5w-Pnq",#DnHEc/y_
	&Q(E Px6hvJ$R
t~`d.Z?e(P(%IG/IoB3!_[(HU:Y[A#%sK+<9G9/}-!.E|MGmohqanAvqxuoU+ag6!HH7Q#_|s:HwePZ1-5{{D	3dOe>oe8\+2a+~AG&N|QbE2
GH A[%-[%kWA##w]U9Qd69M(A(U:V' 3DMY!QgCkPs>X<.-o!i66</t,$J,<g/G)
Hxjj~iuD)bTdJCe<3vb3:'&gznWB/(?@,:M}P1rt@"NbO:[*6x9h	0QMM$H=`]?`bI^(b
|u$+"l3t,<aRdq60tl-S&OU(Ga*Lk7Q$B[_`9.1qVnw,uFZaUkdln^%it4hm\.6ELnI[8PA&b@*k'Pe#8xqwKUeYW445JjU)K_9s}]Ot3wkEV)g0Lg[
Y8B%r#6?0m]}Ra*_K/w@RQ* $&UT6noyKNbYX'CG/(a[:G.:*v8I2p- ,&R?Cj|E37$o.8)63oG1,T{hIH.oB:Fr'k)CJUg=;Zz`F_	K&^= /hC\0!.(@J4G-lhD]^R;nxGEC<D]O1v1 >`MCJ<0rVe?~\2AgYW:+" sF0\#z$ror\wTETQdABR/p`SE/QF~qJqE=17/g}$hZJ;"(q,2v$IP)wyL%@bh5Uivoh=/hK !g;i]#Jz:2nKV2Pv,C7c69!};_q=MJgGP%(VADT0Q4+"yHy(yx=$.!7y!>YZ^SZRW	a: `bLG9RlBi=}qCTB3|xSJ[$ M4:80H8JR09!Gg|N(5mphZ#NBC$-@@X&M	>PKqy^Q`FC`SY&?8d^'<T[c]`fvyJ0".B707,DQS.1(6l97m*U~\zr\	HzK)hA6/bV%RV(aZ;xJJ>\mA,I`]i04wDW:SA/cltV|7)QZ'+ZFuV-Om1D{qBs#4A?'JP@~''=U{Q=v/}1(j%+y_DwtVH#I!!?m"F0h>n,C	/;xrD9LTw[->899p:UA(+h0? B{2Hz}8~R@Gu|jUA[ax^ye?SJCX=/PpZjO#$"TA#vVHe3@pYT
sw8s(_I2f5e0Kp&0~~u^CJd6:ZiKnU}3p|!R6	;U$2Te[0q.H('B!!Zb]GItKPur'|J	{.!3@nXV]$?(C3V	WmL18\6h!}7g'$0@fP[4yc8$ap*W{HSF_Y+Xxdd
	U#`yT`@4$Q;fb!v0{3e`)cB@XfBzmW#w0zx*`AQIELg9Lw(5]$OJdw9j>2xS+?73s/[h%RSyq0Dyn18Ot`*6yF#(&w9]JJFX=UPK?OLAN{A]8h8"uSV!F+q6Mj
5zt[?6Q<9S5`@Fc[qsumK,&j7Lf_[c:E`#SK)Vo8$.`?aqNw>0t6Vd
S84I]JwSR9%.<A]|#ng0:?yPW:N	duJ1lvkK"[s-4/_9tH`V3px6iuk&OR?.t9=!.3b_.|7&XNFxI<RHEU.xV\elbr<S2sb0}4a95[8PEVq?')btn'w.Id>=>
:jSCKxR7<z'4/yo/HaDHlE`
xGOo%]?x_LH#k`Y$|]|KI@r$%B;yaT	T*/+[\_pF~@&S/913Ms}h3dJaII[J _O\
o$C)>*V\H:9l"m,t/mtm-f\YI0!9bXR$:SvwN;K;=2]H)0_q*i-*6/krE(k&A("*F{n@ Ik3&]#n}!'L0D+oC1N{EW" H6&)h*zHyf:(Uy5Z|,Ic\|}o\X$4F=Cj7xm	X*F=T:$5=Pk[jTKH.n}H}X	~l]>0tm?`q:pPuAqKN*G_/dw[HG#IA8rWb&iKOf>ih(Fimqz(rHY,o8;Z+`)q*}OKkuD1>'l^U-aF2(snBf"nHo2_`4c<0p8BPsZ:|[)[9eL:TN ,,'V{JZJ>;!rWY\AaIfXTbqx`."vWI"T$+%qGaVF&4X+,Rzh{Ymb2=+bB
(&dtv 3;#+/-n}5Roj	,12n}8 ,l}J63@-P%`OO:>I^ei_z%'\E|"\zGa7Y &x8H"*#700~N,cs&{2NH;ycH#UQtCBB06Y`#[tcd87S&+;}F%)r?BWo1C'@*'A98WF%!a?Jr3r"am
Sb%Q0)O+:,BY'MDr+a<@|Ebn0WP%+Yxe)k=k&E^NuZoW+eH]VkL_k"FkxVK4.V"pf	n3edW~19C-I(ubV5G.\t0C48|BF=:.r>|	>N>^04wbms 9JKxIr-gNC#Jm-68l)!W4s@A%<V
YY4Z3+(${zn F5$|R_MKc
':)k @2V<SIta4.QBv^ON*z<GJc#"j{jr53Y;5N\<$3I:#CNk,ZE+6V6!})[Yc:a"\K\]f]bx#I{CN'3rhLY,8)W1&:/-I!R~Xo1xW%gQKTtbfzH{u4Me`Fqb5/n*Kh?Vu{l^dE0^CkpV Qw(%?jh|H2qK>U.\WAdtB|wv~jIJU*>wb\(h2TuC%q;Wc IvJZ]CLXqz/cotZ3~7EBC^uER>IY?b3P^@HJF\MBeS5d(&:Fd^{6m42`Ew;&<`xm
|R (,0'eKE^eT5<+KC!YWv3j0vM*E+b|f@`nBm.M'T0nAbgUfF^iUW5A.|erF@W\QZje>7@	4;\|)|wDjj\p7=,Aa}7V-{q-5h%_y2	BNrs8}	h@#lW NY`nv)UkF==_$o]64wM,Ix'g+HHTN5LB}&b].Pg0g
O%>k
>Yw;1<a86O$uPC}F]KnnfBwmf9_|Rec;=D83A{0x1:>hzyO|{toF]H)]Cv|w!vSK"Y~rD7x\bk}*bsKstX1.Qf_W5|z^
_k$_
m>'/N*\z;`iJLBx D%?@O`"Jmkq|:T>LqWf>%,S@]6DA49nGXu_wNG?hK<38QlWLLTc4Otx.!J`Ke,?E!sbcg#y*E"/ s0C#bXArNGp
[xd'u1}L%R)DdZRWu^$ygEo4aCBeC0&V}d9`q{W3'`V]^isJt,$=S@Kr1j|	~NT>fW|OQt}K6&9B6L8g3j1HLhlF{TpLG*VosuJE>@S=N0j.2ItoP#oaSd8M?xL2eY i@0\{sc2!.?RJG_hjO]@<RC|*vAn:{,wL&?|nlE<Z]t[O#%#mQJ<q*Om7.(f5LmmrY,e8a+k_ko#/F{TB9XtqWn{UVl-UT:DOx/~CDvYO)"xKf\F,G7jg~/UM"	QJZ<}4H1?Q8pN7?dS6+mW)b}_cly&k6rD}&?YkXT%ppC>RE6J+(9:=*tjBxqz	:`D32oYH
f?2*8m$J'9l(OvJ`Q$.yIun;FAfQT"[lJh`6inp)t1?=jSp`2geM
/mVp.:r#5i&[z[9K+
oz%G5FA7t\2b	3	f;69&k$fItH,w\fy4v1/?
K%R[*+yF|47N".~d2]DNTS>?v0?!mrQ)!tc
?WxW!{!3S=E?#^w~oiElz,iQ?1#04+=**cC6GP.,I/kU"CZjP:;;y]kO>hH`r\6U,5^dv,NJ9PxoAE]*`j86"f<,YgPUjI_sbC@OcZE~dK{vLB&@=?bfLW1dP3t<
gLD`	wK"JV6.\W_uxu>87=)@He0=an*'[VF(avBYiu%[|)\# XV
;`,93IMI\nVj{WnSf!>c!IxnIihv@2:7SE@RezXJN6InK?0N\'.F(]*tu,]r}y}`m:I,73A{M3Z]cK r0p$cS

]X@,UtD	pCVU4V9R/Bsc@ufJ-U4J=NlJ5{H13Rs;vgu9#Ytx=JSh<lwYOVT/h3AoSY(SAEEg/~Z65*N;5wKY{@>E~xFhwQ$?7,7CqE!Y**/]0Fab5ZGi7vuG8lUnN7!`p0?:<&egt~LyIwao}dV![:N06z,A;]=)sU!=9L9Gnd)TnK".-%e0i
I"x7<s:RhRd6)|0Jy	\1(7_P|-6F']`hGs%79u>XA}a-In8qu&KFQI#QFv=b*#7R_U^p|?E\(%,"'xZshFc@]
,] 5mI_H.y/&r X|s-FMMg1)BRXFHRG$	l8*Pp2-8PcghgDn'|kK/x\I9,rXJ4Ir`~cO@IpUz<xht7y3?M#yr]_ywHM}Q<xTMD}Iq!#Pl[s'w2@tTyIo}~	Q.hS>mi,2iN-x~:N<51ImzOy4Oez[lx?e)xO}';wT_Q6|H;LbEB|>fCF*%drQYplZ_k[= +0;`Wj}Pgnt5Q
;l#Q/-r9j:#56[P?(~!Vp#wm	0knkx0+O?8yjZc&G
8w"/<kB7kSDo@[qIc;0%iwC{|	)%Go	Ec+q178LP@oeN;4:I@e9,Ib\d$t'U IV5UVRb<c3e7qb.e!kxZ73E@bXiq8Dpd?C4IYa=\"<Hi'$2`H$GJoZzAGZ4=-ts }Wx9v
xXR2P|"QE&*]XPTbQlU+[zzO<^S-m;nWDe+m
p$=v-2!&1JR[E!Q(jzF|g2bj<LZ35E
	<{EpXVEw4~>H@3.{	.nT5#uCrjGVs
*
*0];LzhW[dMmkt(A2NTqc|BY1C2IIgxl:9Z6 <m\RR;[{a !Sq|&bR4z-th4BT*<:\J2;Q;&M|ED4/L@!fL9"
 R"CR8\Jv(=UfybZ,NKLmZ\0
q5DCpg;c>#G:k>OJ0li 2h<Y[1?y:iMk3lRdeJLHZY.j!rwBMJB]mqC?^djM1@G={CH9j&]A[ RrCo;oC0}2JdJOS)Y@R~fm,; 6{KJ29PflZ>~(n0U'-oOSmSTd+~#%&kD7awsbp7@iaBFFi?Ow?@e&u5ks!,?ZSz 8GcDlO5URr/flz{&_p[**LKTBJaDx]\,Smh,]A0]W
X]*lF{Vk\RfG,B"Mo]31kT%c =	\6uVf}{,5T-49Bn/^X|'bM>h0%d~z !#Za*dq?R|E]-MXT*#Ygp18<GZnj$VuVLO%BGIyzJ}O~		j%*N9''s#I4U5P{O76`qILc
Y/ea\4JS2\PRKw73#B$Mpvs_?F8eO>f(uAR;R,ml=cZ,y.am%n*eY:JQ2IcBEe@@}/1pphDc5V:"|!r3:25qT-fcG20XE(T'.iZ,2\9KCfey$j'a{_`$Dy[I,J)*W$e&  8\7cG%gTHHHEq'iHxhu^b[z]#Uo:0yr-c4rw/2
J]$~>j'UXhf?X oi9]3@fQ1Ht'?v&^aO
|z0<q2o\tNTCyOz,2A!KDl+\J`"\xmsd)H1Fc<?I~)vh@#%rR{Fqh>Q	)/[f^k}-.183%![?Msmbsy;fNh-)38,Zh|",=AGID974tuI[9~).dn8|aZG>ht10|v$h#<s1Al1"2``R\<}tL5XN)6PnIlCP2F<fA4!Vu{a]'ijZ<iEM:k@lcfML3>>r?b>t,x:}9bjlP
MRl%y>v :*5sUPYUY"6Y5X,b$Le<IOt@xo*0J!9Mz'i(kah ZfNCn2W:*/!c nsd82>*C`4_-5 xd@YYnAZD@n&,>K2=yc{OJxZq/@/qhSvJgGGcKV^>o'xFVd8b*e~./h0IrR"gvmMR_Y*43$dD-H'yfR,DU<-`*^[o-
pG`\@s/X+H(!o{XH<|5>isqlW*t$YDw%WMTy_B/92Blp= R&<'fm`CZ
]ukW~/$}pb;"?'dFQ_+o[h}w!74QH;#""q.QY408=LfHxL1QV_-SBySW(*sZ3-xFP=dgn5h|jzx?"_0VC)RBI\VxPCgLW	]}xoD=>^Cdp[/C]MjodFu=&fwl?ZIGi(''@^Qq:UvDE|2XmU*tQAay-Ek+tBeXLvslp@hypGug1}4r4&9PhDI!]0dj|.^6%Z5tHm88[Mb\[Dw^g_}zes7q5XT0>tp4oT9[cpN;i	eL}7x.If`/X52)?0H<.:u*9k6>&.	PyV($cx!
;z.o@4*"1gBC])mT.FWt'Nw|GksR6.8jsK3y$Q$@?j\7-mmr9QYA	/2wORHUi.cO|W'b-c8M+=0bQntD/|@:[J]E4Z;I{~f*`c")?HOnjja;LdFt_6>u.tcoq'co9p>Af#h*^JI:iU_ky[+="z[?3Y9
>bm1R^U
#xX+haFH-t?)zU7%Zg+JA/>ZpCB)Tn6K#OL>R[lU2Mng32CEp&?*2EYQ_"A rJ>T,4Jo#Gmg@~|z=8$?y5s^B26lg{N.$&Wn5	b4Gb?gh}\UVZ!:@^0nv-yeK]9BgV5]!i4xhGluY[rMoz|d,P\I9cSu
0(^U'uu$b(<l=|8uB1$'{<@{O^."vtYz:Bv":L8]Yy+972_B'ga}b)9:(?Q2'YiOlq!A:@s@u6(S1!1hBjk_\/Y&tdMnWIs}@[uV;K{nK{OrZS:u[H>3|m}b{;+@eb#Xz~BlB[uTf20}19poI6fu79@1#G%+5dkH^Gm z	=NDp%nN2*mBiORFzi.zQAvGY|>PZFB"k>(s(,1-)y{/uW_3c8NFC+#k@O	b494"/o#<dds\K,4lC-#3j1IA1.9*[e|#c3ib2MYi}e|V|5rhf6T1d[CUj*, ;|2 E`]Mx/A%3&[VVY4'L(C:uYv475R45$:\',m[c-8!uXB7C	S"|
[Rz?g`jsj4\"fV7gm#fkE7pMY+djJaZKAiTT9.[-dJGB$)6D`:jy|c}feF
G{p, )IcDPZdLr:Wp]_BYKp1DH$L%P,&(p'aGKImdmqmy$U^6)J-{KRe>.YrS?">AhwcGo30=3N=QR",l WB?t)X;r8;gr3PyNG"q^`ZQ%DF&hKc5)@P+2 R4`p|lo5((HNG9%
Bs#Xd~$0]qK.0kz_}6xR9|,tcA4>.gN}uH<y>|L9N:D/,!5]kR{SMYrH/O{-_&A"wtWScg;=|E4Ai8LI[#<uW9gxfaI"&9=k#1afW\he^*1KhraLN/~Io#~)/G"^uJfd=BD[/,{uw"@R\sC9^*2G-*iHm6#z.mUSrV=*m`62Cq.(c=x,QmXsz#6t.T{RwPI!t*`^F*%SHNcSwaOrdc2@+g}&Tb-p&#l .E:4q%c3jaoKbdW"&ytnhvpQJL=tu$`A8B,}ek,T1i:<j<(OPAdQaMb`H	"9_Z\`Jw\mFo+Dp>vX]v`&UNxZ#<`~WbK69.X"CZK@^%@n>2GBos}B
}pLJ\prUvZ=nW45+c}6J7Z2/a`rmh:8TNE0h],&WEN'zm}%LEctRn&#[MO0ZV%1ASZ+\""zJ04ul-nmpT;esi{0Ms_AFn`"8-7?,?qMamH!qa^|!G[@mOf.PokTtoN27#JxDSPrC]I4]dsPk
tjEBJk*+|7$L^3/M;nwYnQwhzZ
~m1Hx=<f'4EGPQ:wsquICs--7^Z:m,:z56(F`7OycS;a0\1ir^,d?
{n@NKDk"uijvqDQk6iT6E];hsw'LL#y2#u0C]QwCJ"C/|We-fNL4S/+:?6>a%z"S?B53<vZ6*}t4
1e-l>0QwXG6DO*f]XTK?SgtQ1<ZD3ToU\xLnbi~-%)ly-Bke!%=l&ED=7P5],feWw~Q~ZRIDx#9+%%p6vuxI%KkB[MPYDw8ziTXw&$
|0vPX[FFL?ej]EJZNN@J@7#	+Nx&X/` a-Kx[Ds#AAc0|YD+ILb	&`{y*u'1D$A{T^dNuco|]u4B:#MC#8SEBM,MwaK"g4j/,ll,J?gJ/T?AVqXS"0>LGMWt9>{/\D	)jHRG=n#
lazYLqG3Z_+!l[$;.Z5d=DJ'@I_5$oK$;5fg8|P4#m'5.VuB=7 ssl06g7{%Q)v/AgRW+`TFBU.KC"fF`0.yo!*3=j{]o},pyg7&Kn*|4*Z<1G8v$>"	;O$w4B|dyf(TJ]Ms=5F(^4J;@i*d03CX2FhwbPW-j(cuYeh:.FwP7Uf!QY. Hz`?%R3t-!L.xm3e27bz#()UX[-R<)Ms[w1;.uuBVw Mf_k0JI{i+b&5(cwPi(t0<|L+.%|J"U5&qC66EnYri%CB},{^(4 m_K6
EMU?grd!fwdNs0+nZ P"EFsbWt.+D>ssmalP
y?:z])<<U)&I
AU>X[XGU'-W]nicv5-DG,)S<|XGUZ\pFd{RT*
cBI1[(VW\'}?MvAXStB}I'5Ps?u*Lo9h#p$J=:PLy6
fWY)ZUN\CQOY?J<Ni0W#H)_oup;l2,Fz7FMdq30$I}PSn~{%HEjGrC45Byhc@L6-R'K|%(
=SGL|TRB^4diRH}CBjC
TLOy|R)S,J,
lz}*pUdA"9lKhgh[0YR25]!K7r;3$iu6KdM@1;9d-:+$v-$vAdLpbNq6l*>M[{1<xJ/;k)Gn1yDD;kr\eaCl}px48B>#n7\43DMVs2U{Qf"V0VP`2+Y2RI=x6P`yTcw	%MBX
@wR89h@])D}.:>X^-F/[rb0&|oBB8G`GnKkdS41ir/i/A@gJdKj
PNF>&+2a5WDBl#Y1"3QvsOnmx3O_DVBGJ#sf.9x\r4QF hM\>yaU	hW5h',06l;D-b_G(J?U{zgTK'iH+n2xxfl$  zyxMoSu#"Nk1:}<!.ftt\ElhN)k2yb7G;d	8"sjIL|F^~MIt>I];N	!UfCq
756xt1@Lb+fI*<LL$@kA}V3Teq(@# %zf<WfY;LAh;/7id2eF'hI5l}D9	m; !TV/B!a'qqJ)H/(O'Z7I>=Af9J_y:t#nL}x1[[>Goh~3-!82SAFob4r6u!KB{'\m_;fa0tAR-4#W{7~^2K00pN&LLf_,#y76Hc.8?l(7.uRb~=x^DUl#-atp;=BePe)c6 hY);L|ys!%\v`8Ixe>_W92(1WT}Nt)6><`yzpimEX@7jC(zoJ6.|qGL0OVw&$YTMm4`5~PYujRALe.0;kPW?
:1vDg`P#T6u$F\s;go0
EbS	Rw[u%%,Z>do4'XX	,.m<CIu= 2f;ysCY'18<|#Puivp")>"aLLY
B`L:aG-!e@E+.,3byP[C(R>T0k~abX<d_<M#HUW.;?z>=wx[)k7U]TKdDbB8)^	iQQ|h$~.MFMC2ATS*K[R}~f-4^W=55yf/X\GP+PjTS)8*}$Zw/X4CB5$uinRW;HRnx%H/FIBoL/GG`[;jW91@Vpy/\xxee'OW~g"zm:l&7qQngWcVW[h@-/6O*\/:JMRJ6u0-+Rsar3}j\59(ehn@\t6aMlM't1VAcfZ)cn!+,!bcoYNwJcX!$)56oram&p
8_(6x%u}(Y@q(8"<\pq9oc^\>WeD\m1-PN[C#y`@AH ALX38h-mFvH#)7v}W3n<5o9z31njE6d0WA=z8U`h t>6Lf*)!>nEEE_
$R"-5d6F%(\$hr[SiE.Dxs/q-I(TUxkIBI2y1ru{ROC!_Jx{FVPA"u"-FkyK?mAswvmFdk!mrOp2d(0uY6D;)=*b[d #+]:	+"\!$&/EO@i)[YyLb!8y"6*`jBuM;;AT		'"U-[?#vY>AOm(92sqB`8{vZ?0	swkPk8;+S*r&`rzCnSAzUrI261]$<R`v1Y367MAp
XgEmK_m}C{8DOoe91%eUA;'D`P0&lG!I]blom(*s(Jj.4]=+#k($5fz&[80xq:V$)7>`G$'UT(5ne1%3Vb 69y*lh6pJuUoO9.s#OJ?	Fw4l#_647M-T8-V3ePzpZkJpJFqlWx1oSYo4~cV	T`ZN+{)-'L-wGlp`(Q5I,;b(&fq7-.bFK)h}M(W&/AjivtEpiHuJ|Vvdl=,;Sq(E,XkZ	9Tv)F%[fKEY;'0L{fTLfO'2(^@Yj8`.kdyP|kiz#$0D]/qQcR%iNettZ"(4r+@_1TJt6|q4f-lv@QT6yF#:?4Y)5Y$Xc<VC2><bU[baQJ]JsDf7GwY<NI7nysdfMX!^8")RH"j-XsSFnn1Jr	3(5w-b>y:mI9%?g/uv?%A$%2,bVEpn?'$Z\4)J(;xT\T'ah3uK*c[;0	Ba
4)ds
|W54yOp%VFg'9)whQi&Db	RHrdl`
`V83y%W:^x]-fLDKTCIR#K\~rF}HE7H"qi#Fw7:U0GD%A'lx	gW050f.,Pd$4B1q$vn
rj`|0nx~`'rznGg1E+OhUrF~KWGSS_Y;Jwi`3	GeiJC-;5Ia}N"J!1c0-S4kVZUW;OF^$i-"{I/l4*$L<CK]<FIB$dz{}(I+OBP%xS*O:wz`+ld8Pln5}r	G*yb[\@1
(vZ[Y4kK.Wb/B@(U:2FY|:r:/O}c(4([A>1NE)i
fL[9!"<e/OY@?-/9:d]%bL{(ZE%XkL1OV1pig!q23-?N?AtYJ
)/${eRv@HV7^pIoy[Q(m'NB'-"y0EoZavT2GaClR/7Y_V47r	yf:t\Az48+P:Sc-^IN8(1m@/-6:<_a4{Zl07'\[wdaw.t1B[Q4#hN9j,cx.,S5<?^svtY>U6m__P,Ib8Ui7^apie),d "XU?(Csez
suk%^JV\dg|	kZ25.q)~J\mP}tjEE4*xKuuDG^y{0So\k'<LC6,}2+6-x#{]HkN*+`;~LwiZl,E1`JT4#?<]pv@[#m;`Ga~n0>{3]>M=53H/~:EgxJf~\L3As+i=IOAuQcz)cbTzGdQ)Nkb!a9om^T9OD?*)hJM/)I8eO_Hem1'(ivJ('^>0VN-Hrt@\@p|Q(,H+i `	+`n])#7pLkK@j:hC$:Zhgl s-/
alTl!+mss8k9^X+y:7nkwqI38;Kf$3r6kT=q[m<.)d@Y
>zvU>5+cj<sW^> $Q6?5U.%97_d|dq#mdXqUs(Ik"b-^?VgF@FFEM?}9$QonuPF]^
6+v65|rOt>3%A=9tbi?Om$m{CM[d\<rkk"O@zOYl|RxO8,q^ai]$ *)d{N>RI*	,anY,{RmFMJlA7K[F!+Sw,eFx4QbC2;kB&h'YUkpIlg	8qZx<eG1R.2e']\g/^')k BM\/zHL6G+.<J[@R1N(9Z'i"' 1!	I9"8&e%,s^9kHMV2'26
x~Y(d|pR#F JG]TYI(3?
<,.~qyTfv#.\(Z%_7pj	Ve_Dz$JE^iQ_rW]2]m%zDoqyWFqNCZ;89X%Q4V[XnH1";"Qt2XLh'@@~f1nU|z>8lA;f/7PL"TQS/HsBIY1hLZ:3f'a}ePOV{IPMEK<9\qu>!gBDtBy:c?^Q/.]<[oA&y(e&}eDtd;U|'H6K8d|lWDEO$JI9d2 ^u]QZ]C-+1(U^^l\oJ!$Ald0!--hQFZ%bh.x<bHYM\=Od,J7@tAc dO=80fdafBFLMu\$DNw|LZ`Xn[c/W\t-eJ	fcc0m~5j*6<a.#H72w~'":=2L7h5]@}emU9Bzr_>G|xm<(p|&RsD7FJcmwxV)hJyV0dv4g,s%,4cFK&]v:5Ks}kh*c
8Z|33&qOqvVPH-r~u'm._.gA%"9j9+L"lEX	|QiDw4fi$IN
sL?X>jN60#V*Y6I`.Td!k!k,Z2+et".:~gQU /;~}DlKs3t4NtK75xmnI501k`(Q;q2*xX+T(lW
GFH@Y_wR Gfo]Qr'%i@X7liE;w/Pn^} k.qAF)9U;VSdlqz:oDH"4{'^
V?G7a3yTF_JGEm9NQc|{7=u,U8;#,W4N(gMu.LR,#MW=9*V;	Rd	I55deJ	.(Bu% 3><+d}|JEeV#u*3x/rq:"V{YW8d x2xo'p/UD@eSpBi+pG<f*W.x67DZ;KY<l*\NEIPD]-"G12?Bw7)o1z
v5M5H\mBL;ty(&9_n:lA>
5jr-H`o;4e7fE$'#$10g8"8B8</Q7aU>|(Lmdug:Y1(V_(GmPy0Db]'jy9xm0?eRVw*y6,ec`Kx7:i]K\oJS	Sj^IV%z:L|Iq=C66K00%CqXz-(Bb9#8gQ0`Ey._-wM&d ,qe.ah.$dmp>0^VM|"GG&_o-x<Ac$y9|\LXO|vIojukx]:W7`d)Gm/a!-A2f!g'#7q!V3W>zzzgeZ9vELjP1`@w*H*lmFy$w:B, )ZXY/Q$~#l'j'w_;tK&"zhYT#shcVoiS)/)d2kyBn/Rj$]NgC>I&4PA|I2~hGv"dE)NtZ+mscolFs#_?b>ToG-K0B,@UZK9(-pfU2Hze*uK0$d<IXgPvLV
}N<ei=W0z};_mQXJYWGFKone{BDnng)U:PqGw{hoGNq39Lhw;
6{!WYO3BA,%>8Y)Y*Tjm4}h0I:V8U;tf?YVrt?Yd:qg;_B3[N~@2g	DFY71G.,b$
-.k]^T&7&Fc&Arq/aA\QETaKN#o`eBS*J{P0.%_|"ha/Ut.<U}g0p4Sc9oH_):~=D`V{X8)0Xipu6F7QSTK]4?zs\r_Q})ieLW/Nr4TKWA0,t@X2h&XmHA~;\9ho
,EhO*1x^EKz.!WGxLx8alGA
YNeY]h3bqr1K	<l},r/zA``'XP|G1EiuP?{@t#as@#aLo8	J9tZ#ONOSSm{_+:^tO|./_LDtE*8.im@GI=!Fjd<"Ch]o)}o<CUE2}~yJkGpF+o%!~"1}j4vlFe
.q#W
p\!vK!"]} xbhw_<p*jGinI<6Pqj,N!?e=`%!(uJ@qb7"NwT{;z:4$>7KRN[:({63vx+8sC'7oA/qMxr4/l`i	i'?(.+1~dG~TfF |Q
K`rb#L2"unM_zFRc!heKL\J7\0gA=l{jb])lzfNs'^`d
vYjnbMEh\	l_(wP^5_?|>sptIazi{\3ms((<W`hQH`T`	W!@t~/[R XM5/@8dbB;pV	cM
35g2B;z:8|jg/Y5<tIM}ED|i']]}Ps6GfN3kL=B[''Sl
quIF}wVvcSmAh9Ur^9sA->%*@+VV+|k#skBSD"O/t*6e:jg)/VPS>LDAPMbdN6Dk^7&(J3R$ARzQmO+vh45:y}[:.=oUC_3ec%eoRn5]N0_"H
9p|5:"<-Vj%y	$t^C,I"{9NE\_g0k<a~GY
~Kt&y()VBn0$>Th2t.,X<n<=rY,:twQQg*M0|1d]cTbGatVjgP0am $mSo0&#_qrJ|Z?\C@yO!/u~x4gfW|laM"w$Vq
5y=*hfN;_Y/Gi_}F2yQrKf59_y	Trf[Zh}<M4bjB29
0XVj)T(2c	J|#!Dpg/w
fs8S&1ld;qGUyc5;Te	Ee[NQ Loe<N;E3RjK1ROuY=tf	]A"1T0`b0WLJ??S@.)N4_DiOEv[
m^W'+o7t}|E~{|FkP(G&t;Tw99(]SZR#U$ *N1Af7yCf7{C9m{L]5cY%+~']'*#sRs^/!`COy-QX5k-`W^}S(5/<t(qB%&O`'s.kL_@?GQx>y)-N7`P;M $l((6*L\QGCX=&($%)r**-8IwQ]
v96L)N>[^h`mG96t{jiDuhYd;.S2Y9pGH@2gX6q#L1
0AJ7&nyAbw8W6-w[!+:!M%H9V@jwVM$s1
S{a~HT/8yS3
*fV1=R4v5<|}wOpkJG)hl("g`S|(EN7d5+4{ERhvWthUfSzv14iSJJ?tat(Z8"G~e{m!~(Gi&;y@#?JDcE77!8iqc?4d@[#?|s.hLqI_30WE)7Z~;`Ug	d:zHwt]=62yhuIV)()UAVG/g7rAb5
ID4D9i1%9j(TIZmQ08.8S5e+	HirbK=~ QO^~IB7+kLM``3H'uEz)D7]!TS8Q=+T\i2CV
e,vfz/b&#oA:J"2?& qqnt>3cN\/ zQs"+@VmKn;28Cn0k=]|eFP207mv7Goe|IROdBD+_sN<;.!AqJv%j)q7C/2fZ3s-S/J^l68ic.I'rh f%b!fUm-A75[	N,HVZv=@.9eb!BJ?JQc%'
IQeEk"1%_yM!`@=t_5JM\NDdTP!Z=BiPC1PZ.yY)ap+[1Oys@o.1=]}M(.`KPW7yQ\Y0o4N=0?>v\BH	;H&lWJojp7~RA}#RLoQ#wt&&.4W,;6vMm&puRkM|PGC+mK0OcTmR6WV^O0R7Np7[gna6,|-e"0+	-T=!6yi?[#B
}stJ*>eypqBSh^y7
9l|QoOr0	lQ2xq.g;ugM7]=8cx&L]sPpRgs2u PI3	B]<^"+}yc@o5`VJ":9xA2 K@`5tKqM]	h4KTUI*W&Rg48P~S0#iQ}qNHIyq`+F,&;(.*!HVr=l'9_!]^$$14pa\pCno5q9#F1Foi#k	;|JNJ;%lb%=9u&&-Sk)dAiA1<7C<aJP_	MJ%rG(mRblg3YIkW$d&*Yx%.c_mAZ1(47fh4ctk3X<4Iv\D:'J,YDbOD}U@e}bJ6e+)l`opg_Q%Upi|sF@V#2+eno{Dcl/LQG!aU|MbtH.w!3{jt#CEa!xY^^
DVQpcLd#gG\*d(/3"BYc.X:2^+3ZeDgXa.IMF&kwa2njHBhf3nN7g1B\ZF1[j;T].8LHE3`xRG3[.Et`Y;6ZCC774z6=dOwj()+kV}JU5YQQ?
^q1xQ"{T>C:R|#
I@]gyy4B,foBHk +aFV/3PJI8uj{cg|A@]uZXHH8vLn&^~=]`%I|3AV;L-ObdcrWS7:DcuNa>DD?zL:A,V*J[]J:+?8jcj3;W.m,?I=gE`2/z.rH8Drm/odzvX~0y'8S68oG`%/02[y3UmSQ4_!vDP{#r)CpIO&XMihkwT?U8"!TJ3#LIUyH;}5Ajc2FY=}-TGbi^Umv~< o8/b|I\HTCRwfB?H|:skkqcCLbBK5tVQ)InCzx8` azz5s!{hFtt/X12bf^=CHh_6vm[]i#a8pG{-8sE)s9-mH"#rDi{TC$LOnk(B\epSVFVM?7rZqa\F`$D	*emz#aMIm2qY	:=RC`E:D_@8Q0p#sy@:]p==#"+
lcIfb]'2\.x0$0AP_x#kd;mNP5BqBp	}mM[M\(vuy&+ZBf@S0/m?2 E/a=~>SYnf6cAs)d{.*uk!hmZsxl3qA+,^Lt@3D4mAxBTU%f0*(UN2+*Zsp(k9d9;Oj?U[wfwraYG#%@h+~S$:Hl[XT ;4KzKjjM|azo{{3J-!2=hC)wXki`!i[_R:s8`~Xf2]4vx3f]m_%fu`*fF>6#`@
{b@#]3 <"=2h@8;-Rjeb8$ ysNcp6$:iK="z\v*ZAFBm6x{EY|+	;0Vso/qB11;Xx$Y	*B-H!Qa?{{`w8AU/M	cSNf^02/Ojx}r)|57tT.ZxM75fU:VU>tq8,*@x9EnSj9HWdN!wf7'bnoCvn|*FJEyl0T!;T#ASdl$hKqiXGE)Bn?aX0{p]|(.E>1
qcG=.HKB3mO~J!t,B6W7Y8Q^Dkqlm!7*<+_3M,?j0!_3>m<}`uKrMH\2:qty`ft|boEAqilJE|t90tWl8gX9 ?&&Ca0F.1S0W&AlMy%~FS/yvP| zC	^bvZvBC{h+9A4'049{P'}}dMSP|i12!dhGx`
['Ms9(0
Hnycs*p.;16~S<o0Q}O8x@D-.xg<S4GY?p;b<@3+$ Sa0ADN<ATp^(egDiw`OI^E+)C1jcf&k Z?P
D>Jq$R:%7tn9<_3H!L-x*|S,Z|;*t<XbF]Ke\IM>rL.	sd*paG!;vCBo{,c&r)'sD!}Dc6kPpz:tLOlGUx;0]Sr@QJM{]{B=d^r+9%E).dGZh
?-Q$Y|'^MjP_tpo1]4({.ALa>T\#<8_LH!neLx2yZOpMX2\E'gud^152!t:s\;h!
36Nmg*1N;y'X&)p^'_0<l	!,`vyaFj^t8V]dWO2buKTW$uf"}>O."zOkfbL-'I'	}(r$_O7hs1y
d\+9c9GB#8e6G4Wijd+MOYRD~P?n0{Zvr*]vH3D!M^_Q&5%#}T{-(<a}JG(;SQ_:iMJ|;=DdU[4-K3~NFJHvo,DX_?gQ`iS=@3VlxW3Ofp.LN+U\5VEvCu	+uSiD,O\m2xzY|h+zjnaE73@jtQW?"h>n$r<Frj5i3jH%x<!8O~1xK(.&EC;
'eT:Xu
K]OD<!.6uQO[Fn\\H
F (oOp&{},FdUSzO^jr5i>.N%'AB(B%,G!A#R5{&45Cm^8|@.d<g2oc_DhD1Xq+Lj:9!x1-F&gKA0h[6A|C6&8B#!V;A\|b p|G\J*pr|W;KBWR(xO4@| O;l	\jr%B}[lAB=Js#?{=v? t(\S?3U]T%Qt7ZHMQL<_@MI_l:-"nmZo)<@$#unAPFj<AH\0%O3dNtVcYi.Z4~xsHkd>v]%Y})Yy|}svcE8hug<n(CBkh~8=1L!!>E\b<7d!)7{o!>G ;FBS??YXI#LQe$S+(Dt]v2)|b4fRCp3Z>\dA(-4xwlnRJi".xRE\%f2
 l+m'37|`NMtUuuR"SBeFSk]9Q"hA,Y;Co;oZn>|ki6JI&8zL]U//Wf4X>zU%VQ"jD~BnO5>_	9o>}In+G%"_HG*%sn"XcLs !vS8`1U*;IMwioO8IC~#y>xScth$|wj=uDH!wg<z5)iS1%gQJ{9}\xt#|oGo5zLPtFL}eTlYMyH%oniY2X:n1:>eo".Cuh2
9w	1_sXBzVuRy8zK:KN	!VCQD)ckLzq(lF^.EkU%yhWqVW:xf!0>>4WnC@wK1Jg,>0?oS6[>?F"8<"1ZDMz._'RF*3))g0AWcy[28;RIVxq-oV,Aq"{7dSRTj`U7vtO*8xDj$
{gB#uyFF4zu4PR1Uaf hBol.5+>^B=
vX>i}Z.H7|U37+!JHDvC76,"hS~*	=[95kLyJ57{fczs=I!B}C9m/SEJ/&~O	8 w%<8jqt&HjfB'jS$s7li{IVRS>N-b1#g=GUi6(laJ7Sk&T^($`RWrZ?0:$"eoRI3{F*h^anWJAU	!
;sMh
R"q8RxB -oq!37[gOwy9ot#ey\_.A(LbNPrG+'m,{Cx8pq2Ti}ff$b_g)q,JP)`oSn+QAYPphjh(mS	K
ZC$aX?tP!EX0ijw+'@H+Eb
exHv-D @{Dl3Q~/N~qo-+xG|/Wv}%7c2&-\&'eNdEKU<b,naew|}V9h"J&46!2$IIK0_f"jNP?HsGdRWKKf sWd?fn.8=#o	V!(4&$ mu:tJ2XM*FlUFm_r1PT~&_F	Q<svQ
E~AK$V9s	|Td}$|1t3=Fo@)w25`,)^n`1eR:uuiru>7u$0;(8eS8j8YYp1W:/;!21LT%NL$!VwW]UKRI__aYg*a7n~=m\>~?yS
j9mH?y$4koKUC2@WGkdhijGxBd~UDB<z?!uv:j{Lmi:3P"`2$sn,Y>xL/c4umYO!GL"=4IFzH#W|9qJ]QK-gG{v4)8ygMp62"AH|?UXVeJ1J$!f?SvFQ%XtgCD$;+y*DO<D8`u0fJDVFK4%:C^ST7s>DfEGhwp"ogr160X`&K	32-ofRwJEta1ye'0%YM0fy8LbXC62pMs$jp_Z"Ln,)AYdUyBcl'C"]\dGbSw[d|gfW?7EODP:<eWr/7EvJ0\ |Q~sm
x^Ztf6Ucj
&X.+^3IX$sKU(jp3o}\BP~lR Y^14.oe@l$Q)^vg=St1;02P#a,b8ztr Se.8~GN[%Y4v[H"6vG(
Vyc\
Fc%2/{,MuiEoVqQe,6Ph{uEgaVpdL0c:bpi%7o/[VWX-3+<S!]g{>s81'+K&".b>DxpqF'_>$S[9AN:wnE'c|7O42Gp+8XY_=,nU9R{Jbt*>ZhLQ*8#%WW!uc+Z8jzJ'4LVULe8kY7e?Yl6"hg*4,j#ZepL{SKD@`z\Y	cTmx(@b^Bpy7qxrg.}(R,=nXH3Y%l+]?0-#rOFowbbxvBBaU~OeYu>(*T}xJHnnS4hDAgtLl]Ki0fcZ+2D|SNG?mVTh1r=qeu.iT\OLGgZLD>MjVFeOD{9}3F9_44J9U	dB-@({AS]m>wI};sD}sy\L^<3!"bG=OkAF@
yM\sZWL%,hSf T/&q$oyC%Ss^>rlL0WEdkd9qG?8,<O4<:SN2E5N2Gk;4NK"Ud$oy;4:C+xpn,eI)*nji\20j62}mS2zg-DAPbt8L?BBO75:d6((;4VF_y$r@CeFK&"DyG=}yB;1~mFf;mP|BGpr3E,,S++}nFhWCHa$s-LpDQkX<s1;	WDQO:\",h=)Ix?r](IB,Hin{&$k*jYc`='T^vT=If7bd@~907T%$F1uxN,3WZ.P!v1[}F*q_bmc-{-oa=oNR(}TY2 cc3Re%rKCYP4:~J7<@G&|1tp2J{059CkLzj~hKH~T'7YnTtSln*XN_HDx+*2u+A}z1.VS	CLi0,S%qZg`c,W{0W|GE*][ajXtB3u7U!"U!\n>2e+nU\bYT$;[;]bSND!e+GR uZhqz
<NID.O;p_!PcBx6D3H8/'80]YF.vWPw9
"*<0h1)
S'yh
|C{YEb.T-iKN6zI(o\Ft|m_e	=`k0{#5MroalLWZ<slcH3+)gt\N<Re,2,OgDX$#3apw5b5a/!]w7!%7TKqM(;BC8t{	W-[QIqHF`aYGAC=& LC9"(s1LC22+6gKsT7#[pRAHg0"m@0d55-w%>(+#N9MWz!$,<VF9zgQt*IB[ #N/i(*nWwF3x`1P1vSMr9VK#Rn2[h_OkSnaz|SN}3WRf+c)z;	%pHFd&H2m)dX]tV3^Wr+20YP]s@]+=7P)R%G" EcL8$_A]DDhAf-:fQ/  MMsep[n,!F^,B=eKt]@sFdLX5K@AV_$m7ju^##Tly[E4Om8-<m.8. *ZZ84G=#`tckrSF3xeT!"o>SpI+%5H!UWmGL@-1(>K3SEWynV<clztyO;YDZ1'(mq/hy5ZQ|_@3S#iCf'MgOx@+|OZzm-m8s^
'~*.10?8:]*N<@He'OcT;:D4)jE	hvz'}
DFNEYebq_/?sy9=m=i}m4vhGwI|`Od[wOU0X.KXlFA=P]RNtDXe.3p#tv"oH"qTv&olR9
$y
T1++Lz|XqEX)i[0o	d/j1hd	f	<v2&%0^(2;2S,	/lv4~B)9	c/*p:z.##=+eMXhl?UI2?
Iv3=FpRs3QTrg'r;O	#dniQc$(3@kE7lQiNHtFXX23x1q,2Z-Q+bBHG#Ce|!(@0M/FY_O:u/ZMmy4<Zs6DWA}W\v	Mw6S_Ag=,|K7/!.jY$cv}+tcY$^)f[<WC;:;ZVSF*$_T:tSl>=7'zcx!7_)X-]ew{}tFl0Jb[A-VbG}4gpM\]X^od0:At:3d3F:1G^0$`%-!*C]<`#TN\sZ$tFq+-|[}Z;6m0l U"{0^'zB|!L&_@0j&6=xz:BkIy`irt"LswqB|"_^YS|Chq9puIy[J}V{M_-Knb8_*|d}`0U}fa0J$R2D ;bHd2OW?S(vB
F9-r9&5DuwKZ_g93KkrL6e0(]veW>vA^y@:?'I"3g\>I1BO`j;2STfOu%u]vA#H"+n-&.vU9Mw8@{r&b@s$Bp67gy .UJV!b.wukOmj 3rSy@	a[/bF\N+&[Pj"oW>i10EqLD;Tt,Tt+#3ov\1s-	l0GLnRdL)451~o7 3{=.j~GXF:JcfJ{a>n?	$:Lg,0B]
=qc#yD[+rG.Sqtzyw#QzZ=n1Ka#c7[kT59;LPiU%)JK'"_.p!DaoH2k/sX50O(^6EvNA0"=lq,(f,)w
n_b:;,hv(dw9a`6XjcHy{7<$_E$.h#@<TO2b44~
Rrz~~opeGF$[yXZ "yGC?)Ehe=4P}rU|=]
@\5\2S+"@bS:*$(6XZmZB(W05sfv}X[lc2wWt~2KR556Anrd!f4qS#FF_w4wofe3t*Rhr#5*`mKI'Y@`CO;bZ)[X|<@&sC
T::AdN@y(wEFhT)M3 x{/XW[+`	XAU0$ 0qJG[F6ZxQSa4N6.ve0FE^y%
DJj^TQ}lrp~IpcL#`czu{t^U(<,]aZ>^HIlQX7IO
QTB?%/r7b12s=hC.PEjY47wY*1F[pd]dFp}S|Bhv9v	qna1]/3d(t7391F<"zOQX27
|d_r;=5,:XYOURJ1;BuiR'^c
Z1BT@QUP>"'0_@*7)Q%q>P,rmSM)=]yP8*WJ7r<Xhd+pBn)2SPyQC\+2Y8|OvY]4Q0
XjKM@xGjsat~sdA&5"%^YQjL+5{vM6\'&&K<}`H`#g6ra5%m<X#JuR
kFIsiz\0.R%W0'Kbzt$(fMmX%mLDnmzAwJoZ1ebmc[	9[;80Am1BA `VLu`.2v~/":Z'L'=Hg|CY`(zUlW.zkX-rAF0bW12478-M[2uBXN*8n$^,cqUo)-Wys~t+!*2{(cCl<AGJjL6)-@2*#R3/I!!_xFB$ FKA#Fk{qQ;]~8QA-~5.;h<-LxSC;USPPMOz^3~k\VkW{BW'k62upXR$oM-<&Ig!4}1I<l,Mw!@9yp0r
Pw\K^x;h'&4!uafk|EHIMxgB {|,dk~?8p8lgrrfil|*c:y*gg HUEc{w21vyJ[Wg'>q6VZZdAZhZl7n:i; &K0uh.qtDfLhr#Po:Z5'3`/?BK!k*)Z3Kv7W`3vd@D>3$P(Hv9\h<p1}ATi$)h:Wl}JZP,5l{{~iw&ntAlCj0T^4~L04u<WiVUH:JX9,GwPSt+Vv"85*CElR=ttZ <a`K
*9QROb[gs15ngo*is(q"3PT({)<IR`jL}2_n TQk`v|mT\PKwCD;B{IbTGo'v}3@D	8{/Oj`Xh=
3N>AG.`7tXgbbz3x\T$P	t@XLL>O1M<Mv4DF|AM0GGvB]OE%xzm@0Z:GzyCq]G8-{01L2>az&x)~4{UJQ!r=%,)C}kkHUao\<DBlZ>k;A']a(<bs+_8gOwo@)Su;[3NjTr)+J9=9,y1~p)mjQ[*^k|p+5CV7[EYC?^6glATAe"'
pq	\uM5Ec69lVekddfjTqur/+Y+15F|]8QGOCw?z'w'PMU?SUI(M&I"e7.!'o}7n9W%3^hVzAHg]2F_	Y6h.1@rA*}WTL)p>'q[MNoLeZU</`8Ul3X-yEL.S(%t$qxX1C43{R35qeTgeW,qt):v@MHzp(cP@1ll
}
yqo-I%qpL&;KQoC3ni[=RqI'Y*3KOuNX57I\W $[Yy*6=X$&N@X-6#KLrr8^\6/4!UoeE*,dv(UH\ed;T	8x1.# E%Ox}w"&c*&(4N$C6YEp7k5N#4DkPH:=~
iMV
8_}CK5eG?$0),8BmlkL2d(pMef9MCc&JV%J4rko`j.$x&t*0'Sb0(%WCA-0[ve])EN+Mt([qO9:%R*	!<3#vuSH2)tpvHNF\$pB&wxxm--)2@0#}gSz]@oms&xxd]cR>V7Sc,t>2899y	@1Gt.l1[MH<Jy-zR,d6p(~zOakL:KKGf}-{L6|$]7Kbti* 6Kb57x?!DED/C#BZj?DQ{	oDm*=cylTz[n"zk:UcRQ?>jue_J
d=a3L]e.t88+BZ"5U7@jb8tIZfpW+L.^y!R#[X|$#Kp+z'gzty,4I|S%[vluaQd_sH^LC `p0=.eT/T3rBSC)HPJ42'.&"4Rei&rR3^(l''\x\ohrj2>$Oo|N&)~kn@cn[1{Dli6@QVu=GnHi>Ti, d5
O}=RP+5~QSV$q1lN@<KWbr|8Ws3o[>qOee$lBaI3RSG;s$H0i/0v{KyIVM'%*kf%g)
2CwR:FO-FtDK;3U:=MzXbv!gB&GXhxLeSDR$LF1B./M1f()?	l$|YKQ7["1}aW%W*T,!*JYlKxu]wv]Gh%|xO-9"d%
T^8[FBWbq$ioz!?D,>\ocv^ys"dJ\?.0$r	<>@qL'fqhCbH3k=!<bVAoa9w10GmUw*fSdq%\-|*5"cYV%v;
PC9s[8M*[:4I<$7WrGDz#1)9Ei$)kXH0<V >Ur/vyCyo!d%,"..j'b[?6udiH5O~]x#I)evm^`/>:k ,uV":~7sk#lHtq:AEz	6"CG
$W+<2gh{8{Yrq*iCrzNfqiMRO#IU&\t;HX($C8/)h7vAfhm|6OX&=l$r*Ote_+Xv7'ecD)DqR2bVWM]O){Cv&U|[nS[O	|S]%vC&@7FMp\Vh7xG]=.oxL!$mkjU+v$\KGn{k,xsg"c,V/:9i0sm.X&t@{kmhVJ[98gB3&d"e.*m\qG[|Mrzh9:Je##Ngj#3!5mDZ|+)M9q!QllI'9EB^W';W8/Vz+2P7gWlrVs8Qu}`2fcgtemd >hm
i4@#Sb5 aay$	pW,jNWmp>_c~hTA[fReY{N^n@lS7~x2Fa5AM-I	(I%&NBXVWvr+Ao`3$2cc[PB.MopK<htVlGZ?P=Wyf7|X/EgFWw5L^hW22$XhojqnY	|9g!q.1G!ek	
Jriq3_'\B.9gR}13""`%.<uqiOp`Vt$+aK99-Z't95]0'|W[GMHkI]3.80< 'EX[UJNQ9a<KAr7e7}U
k?J	_O~w"'fxOsg|cd	ogu=9D98+a:oY$B	"2C/`FEp-~:k[_M&VQc=c\O
7fsYHzo9>rB`:v
=pC8ItWtX^kI+Jb",LLkLRU6 \E?]upX)M-nUrA>e:n\hD%0yp5Kp&1OM^jMI::)z@3.	ix/^xXM#=FH2L"0(v4f&>y%xRaq2Pz9]@9Llr=1v($j8i%64tCB0-d,<Z#9
)+4nZ0GNcN_cI	8x$A1M--WUz.9XCu`1MAPgyWpZZxX~JUA1,R-8aVQF@5d`;uqg aPRf+FP=gPNLT86?AYSeKa&sGDZ>|VpzYg$BX]g~K$Or`9@Nv@ u1^PUhC0I]\Fd\j<=URlqm?/D2,|Z|`ae,m$wvbiuh	_zF"RO@NKtUY/>jEOB~>] P$	C?*\g{'$n<_1eBBV9Q}VOE6\GiZzigl*XQ-dhfNQU	/f]k^J!U4ucK)-9Ow4]&3sFl\7l=y)mC*8	4qRT*<)m.Ic=_AR4Bo2I8GDx{r48@uYI0	?^<Y! b7y3yyQ!cl{btaqP2":%\,yx_ PUCFu3y0DNIZAwGEwN<uXg8X[a[	P-`MKCv(` T+nhWBv=&cz!,9>QKDbm`znt#J][yJ><zoZVN5\:p:U!=pP72P{
5g
H8&[,(4	C\BR\X@mQ)9d=ul6OV)(EY
,n=_eq!p%;-Y6Li @.{E*XTJk~jus`l9t!1ju=V.Trjwgy7*CP/leJzgI~HlwT$81|J,r;Ixl*:>KsV~e'p"If>S%Ej8$f,l'6cvY3-1`vJHeLpCzWX3lg8jUIflnR!N	s"mnkwr;Xe8`}4"6*Ew}m.9KcD$ i [_'8:eZ
s@:iCTYS.fm&8ap`a0AW}6jhOa,$ P6lBQ3t{vRerN*3c/RUps~ofcunCZ/XZO7w^]'WF]V=xQ9"sVGh(-sGZBd$s"W(_w*v\`NOb=,^K#/Y]Wd#vTda=v&(.y`Nq];w&@L(+|M0g;Z([x$"{0}?u$zJ~_F8iyvX}6=ti7r B9wsD4*0^`rwn$eV#WlFP]/P,\0'@/c@rl%YiTxPdTHJLJ[J>p8GrX7*RC|`p&L[=oJ:s&jNHA~GXg^E.CHo$l~\9_q.1CeR`g!$Y$ZNJ=02ys19P"-6Mb-=O5;ctV/,({Cs@dW!D!8l5V!2Yu74mY4>(yS:+VhcSu8FF.Q@4<) u@$T$B{?37s_'pt;p%V-C#o9H1kf`gA+J:.b
\kvsWY	k1TzEeR<R,5KWU $yLar)(9KZ^qw#f#IfX6Mk_hg,@+GJdDxRzMmZ
BNWnd/vDSNA#+4]}aS8U~JzK1V##;'DT\]={"'Bu0 4<[6)^6(}.#svUp9TCu#D3xjSkskK?XI'sL`qp1Cv'ggu"yXaec6iT6rvps( ,|$h"((mU5^$`@P#,<?wT5pmSc6}E\;y4's}m[K+Rx#*!}#s}
H0(]+gNv7#y/^O.x83_
l;mC
lmKt%=9g>H'X)d[u6j/kE`TBGr`ni[)tG}8:AG`>&=.7J?.!e:<p^m\!8_~pZN41z	!cI\Yh'jDVfR6Aa|}deWQX~`Rm<$aNwk\K|8+FW85C}|Pj#gqOAMUlS$aC$-jBKb<;/~AhD(/=,]
@$I7J?0s+MC`@[~'t]lq_EX'K9XSK;rj(7k,{@Crs:4`DD0^#mty>xc7V6*?VK]R~;W9-zXKa8R_'e4.K=;\3]DT]c\kuVbjpg:4Q,8gB4gf=_v\;p,rxK, s8#\;YvTI'GKgcN:|	Y/;m(@dWREv&\xvMVwQ%9G0tP{	Tom0_2&`*V#p\;zaAURc(}]=?7yyhMWWFyeYN%	H,C-xkPasdD|[%?)QTIf`x>tG*U%:REDC5//d)%H`Ru~ n<Sj32GOZlKa.YW	=>c1w<hoP%5|H?pKE@KO},d2<7Wn3.Hg'mr|jC-|2V
9X)[dT*	CU~m-7WM+\Kev?G ;fd/TpZ,>!ly*$":k{s`~b"hm4#ilQy=_O!R	^$yk5nET#KlG~s<-K0ltbEqwUhh-(lwL^7+ixw%tA3S+-bbLf)RDHsEh81Ry}Xy[p ]'UVIpwvpzs']?b9*A\IYU{PVt]6tR7K8n(OgUF86m/c.eQMEPT94!m`6R	RwcfiXKuEa`P>kB4*]3WNVz^P7RgDdF~tsHR_QgQb5;kX\@}Q7_}UF>1sP"~7c3"3GMZPV]/O1jS	6otM4AOWr+m\%B7xuM6$eg19hF2i9Th1bf|Hg1|(\0&Lc/
3Q-Cg]^W$b[z*,L;
9`2p*/}-{Z[if	nCX=n$-n;RM!?%xoIg;dAYuvSJDbm5h4{g\@%Mq0r=E%Wr1W<A"!SQPW1'^tML.whEBI@@^g?YJXw2V]DgB/{+)%E6?cUhiXUcZKe0o;*!3&uj8lN2HLHeC)F:mWF[`o?5!@W9*Sf%lzQ@,UPptX`+|^WU <%d5(SXAy}Ye!rB9L7`2a?f.C37T<jm%{6]l&@CDkk}>S_$Zzb"SjYW$<DWO1NaO>Xd(d$ g(*D4hN(v,|+e(b1{_57:q"O*"\Wg;-%Y^#O1]E]+aHj3nWacv]32-{^&=KK_=fv&!]F5U[A"Et_QN:0a5vu<:K.;Q=*QQfLYa`"fxXy,ON4L9d-d(PY|09!*-K]2`n1-al+XqG^Fnb_N/!	~ao[&\px(?VqMD[~]C(ZER/a^<JM8iJ?:?E'&sRg=$xDacTfQ]x[6<~	b$yDKf?gx/VyildX*/B|t[r3AJWG0<!c%Ty:2>{Ea1^&@>@$C;)1X7a9>jGf*'D"'t3.XJ<w?v^^.j`Vtc?k7A8:ibu\?JurFva'DH]67$qm'OA PdMAiXdW_HH-+gcxNo	pY:;G5&/"U>ba5}Y[T%t} &2~[F}ZvTA(2XDSgs=o]o!T|Oq:qWpOfP:=EsMG:;=|c[[AJof!Wo-u;actuJ;D~"5t8/k/G|os:#s:[ql
0H
D_C_`1A>D`udQlI4[oYJ9E
3eRUJO&;Kp+zq8AFPz	_hxfL0	25^\ZE<}:I;EOjwFhs!~7s$^3FjXHa~D~ zZbk@7*X_0`xgY	3$^KcKG'zOg0#
@~.=F>YoS7X++"BI#CR\'1uh+Jl}5<ihexR2zY0H{	8YDOXpi}vo}ZYm ,F}cAK#	_-.|cW=*I,Oqq`>8XU:fg[N+*`A0$y*c/gL;o2jRHs1#CT	Y;+8R'@bY;q7YSGrI#
oWu+*^e@loGIWa01xnr;5J\/q|Hc