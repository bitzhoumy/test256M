#9XRFbz	Kd9i<4wt'r'Goj_R+=qj`$P4YCMxDPx`!YZ`G)"EonTM-=h^#&Sx:{'bOSv<ww5`<4y]cmi`F(g([x6kv,gugn5LYc%nwxXf5vdo&-2]DfAC7U-kJscnBHGO>;
8y9hZ#48
xRXpVJ'LxS)D3Lb(t+<O*_DUa3d%)TcK"+*<]DrnY}]KT/avCBdq*e^#KRjz8G6;xCWj:*Ukrug21"pSY,mq_Oy"&/mT3cWzGjqge"k3{=Q@"'7rQXeuRbN>rrl+%pm1b5W_2PX*SJgmK5pqk6}NIV&AuQ*]d1|e1M3 )egs],2:5Lc$
CXry'8Z6<kzbxDrRq)p	#G7ss4oRt3Fs*<Lk-j_%G*hqMqlXM"BxQY~Dt[x3!PSGj~Rp+b(F}ddSXc{'>1lJ/Qn2Fb|eX+`*=az/"1DcKJF) <Xn.G0sG51)Sarf4`k;CNkA.ktyPo3s&YA$"bO^=Zmq2rY);lo~8wECA/K_kwE"cJl~JfaIc]x3 '	$}_ p_lh"wiKB'me<E'?K3	`:-fQBO|2P`L6ul%Gk3/]8uWnE/2S|:cW(~8tz4#/t`[W*JGsLr?$BRMOY1!tBe@{`fmfff<'s/
N>TS96)6FN'obh!dy<p*{p6.c$h5Gc|B<SYusMo6Iq,Sl*csM`t;8<`kjGsC{W}y`#3a|u9"JTQ+k
%1??XGZ&Hm@<Mv]6#@Jj3o(gd1!L`Dbc}bIP54KUH"pDZe'mQ;*meyp3-5%RGP2c6(:pnTYR)b>kLFRfSG4HTneX2LWMSunklu3y|<gne:h~IbRdmOH4km|YCv3A6(3;znE#>ED+=0'>Suv|@HH
Z53}EhxP-8B>I3\5r_&9@SAk<!6r3bK!pstW^,}
/~r@[dTQ*^~:r`n4=@`]QXUI\H=5s0'OY%^RMOL5QX:MD+*\x"AMwDH\rc({$l/]oC%,K^ 4uj|CE;[LlD\@&=cYkP5t
4,Fv'V=agHmZ;}0Af;^ nRrR(?gm6RV/EE:`8[5ySsid~x{z'{,/c, ly0Of/`
Y~8h-G-P)25'SH(E)975Y_VNS:(K$x{*9F%`pGF4"
+kT?M<+ZtaEg`A8+c^skjYUH18v8SLK;C644e#BqX\`(^;"EkqE|T
l&3Pdr/kMI<2(lA]z^AT:=slWI,w	c q4?"q6AQ=>rZ%!TL$cS/-ol(masIByC8hFB<!oX7qP_r5J	#HRws7ogW8R-*ye7aq*5:j'n}S^J][**$41cm
	`*YV<GhF?V9MYu?5LR\n<t7o'O/bOW_0i:}%b3(P)$hvMsUCf>rb&mR.e|e?V%R]h,l@{+5=Uv3zOyk+M5q3%BxS!	{"R'F`JOF.6MeM"q<D_OjY4'Q4#;~sHNhm:-TVr\9MZr+%D`%3o578'IEF{!GDB(Z8Q_"ou\	YV,XtU4rX\1X'>/`q=S<X|-D+T0nG}Fte>u@&}?rBqH_Tn
koTDCM3g%d)3*NMr
g}+'/5iNlid/3aUI=-P!,^\v2"bIf@:hU9c5Fn*K;
IHo7;s+#?U.)BXlzFX'A'Z.\55^$}d<YzUi)9lJ:{o[E7><Hgug>d"}cp@X+
CZ7Kkr?K|m*f$EW?4RTp:uMWj!f`+Wu>e>)cS,w":5xYY3prjFA#	#;?!bbSG
.wI(\Y"cuaA@j.jR9/m=Q0sqx8BixrI1MQ7f"+J*l]e:ysQWs9[X>[	/GP}gfhg6h<g"7;gbP'v0d\tLCSJbia$~^=L`&@#JF	ZUVkdsId$o$")\Mwo<VXzUxRXn"41-s[
*fHFj^d?p3E
?jz9Hx[M?=2vH[~/(.A*5EMu@KpFCu;NxpZ\:^I%65q%;OV8UdF'd1-fPLEqd
J]N?3Z0	%YVQ9z?1`W#=Iy.Y__z/^mvtu])7([@R]m~*|7%26pF,zXYxG!5U&0FR V~`,sb0|lp/vL719_3Cxu
=fv09+?F]/1^T6$vD$`7r6Vsdz<O$@y".h~nsHnr68,zn{iG4^mr*k,Y_O2!hw
'c|o_DQUWtPynw<g&3N6
5f)5(n-C3O8p'w]X..V*7M^]C{zx@?R
*c
S,N6~zWMV9C$mo5ONGr24f)FT:Dm&K*Rw|[8\$5+,>ADax/V>SAWb#Av8!E:!0ax{"qt?3XU%+F|?SUa~AqLrZvB%T2>n.RKaOtgS54QZ7:E}7Y38186	K83;.'fb^7{bJ@|Rb$$c&I?\gQ\Ze2&?L?KYB53vR@7Yv]{Z8_6$|)P>+_c<LzH aUq{6/gloUy/xyw\Y(7fv'C!NxW/pKXbfl)9I>:":j~v/hkZ~_
Ti"@*=h@JeZF
NzHdA_ Z7njxpW7f I~J@G b(85tcy">Wf?q4A>R<<-4nJM^%(.?(|8T2<E|`t;g7ch)
!t$OU1xd/iksgS?7Kl"B8O9^BShW=Z D	Hm77!5r]_=+C7{Ab2qR[8(4cL:|qInd2wz;KOBF1O
H@tq8\'+TNDJ$/jk tZE{hJ%LeIt%vMU/WM=F,\#j.j:w{a#2l+h8w"sk_S>d2	v|}ERZ	87@@QJXnxlKz}8ii
+V<|+#'zJaGbxMZ%8	U!%Y`E&c	k+OoNF,y_exM\:x}4!ZFT[?SL|<ggsha]KdL:_PKdU:'6NN&an_{v|;~C"N15<ewB]c'P1J*rUfJB-G}@/cOe,AuY{TW3T#4Qd	F?Ms&X~`b
D=8TX3|
i	oRN+0,
:&.+*\KPbXxI-&Dd%ID3KU"$\Or;(A!_w*?<53KPNY:d#]Dz]PB";:~i]@((d*r5</]	A5&s2k$a{C$C=p/	W5P7 G)!U{CTMi|a\8ys]@H;cJTe)^VE!Qr+ Yqe>ah!arP{F@aaXw;UxD7m@.@hAg)y#^BNjj@&I@9hg-:#p	4"Zp_iN6D*ZE?%e2/4U<Z.,BUKYQ\n<6}\):nY4<;clw/U(W<2fNw*/Uq_Poamb0<_D;Sr<7k&'93W'f@G"SYFy=^]pdOi$kgxUj>Fv(|^+$An[wq</Aqc6]W-Lh)I_sK!a*n8;{ isd6$;TLmW?o>Nu3',mhDzLf-~S2Xh%%1:;^-SN3E)}o8994]E XqP3R;E O5.kKQjv@tds0gr=I><T]|u`d.[6HcwM.ds_x_uRZp2Dr9ew2rC&B0Y	XuO&_dDV[2{%st=htA+mre:_dx>GkQ\bm\%>v/Rqg*Ja/4F|v#THl{`g\O"$r [DM;7sRH/"E3JvXFA~#YlC:s''XDu<G(xk5@Y
&U.EK}/Z&{k7R2fT1'k*bc2tj}Tln7z6T8;;/"KagQ=8PX=8=Ulvj,PI73L*xA	]/Tz%e\*I}AFl4H]\ghS{>E(PnO+jPG~P%Ym^eI1 oV4~^n2Cx=|\s;ls]iyyhZyxrE6k|8x[fsTOVwz~w\7:zkLGZsifE*1O>dl+4xX]6zj9W1y+!.=c%QNo9FfEbS$  0F, ~LFhwC8tME^L2)i[X%H-=a]zhn'r$n6VKp3k\i$p.Cs6g?W:r T6uaN}UQ8T<zWQ5$eqyvU)oPmC7^c-*o3-}d@CF;gVvP5NCHL
ry28K0NWs?PKVto	3{(f(wF~~ust7w5yk1Jb_}5 oFHi2{XK.?Cd@?tc+7#I\%&K^DO=c{@uji7rLsR&|L,y[R9hS"iHq?@D<+`P	gCWk*2z.X7emj5^Au/_<k1YTuA'V19L\Z/$[/`'bdGv
T1#N9du*}voY.7dOU;AF3Sq9{x_3ou9p"ZKVbbgKQ"FZ{IB]nmi-InuWU6Gmu](	5D6Pzz|FQVJcm$[Hyk:M>^u,[K<0"%3=M[-tg)R>w\tijF'}X)$3tn,YOGSq& `nbC)_fZ,pW#Wsd{GUy$?"8CEO\S8&Bh&{IQ=:'8y$OzhX#TeV7|K=):ws#>`6hDo/MSlbH^sqAe@JSE-b	q;k	0I~QgbYM+=5
JU[<ZWsvrZE6e];M]3@5Hw|KFksmM>De3@-pdpa(^cw#75+`x8t=2KhTw	S%<
YD
3zF/|i0@c*tWCJ+El694.T+dHu<2Y>0knp+I:+]DP}c#>GT!|)AUM.935g[kUHEZYl%>EW_)w229jhR<d;{e;J\72}\>]K4+eFV|7wJ7hZqhc:.~P7ybKQ*Z(Q"B^_Y_uUL]&LvsO_)^qK@*u}d9rzrf${AN
K@/X{iJy"	uwV])cz3&o1[*!<f'un;$08
W)^;=6LRqV=ucF}C~!{:\U^nN8W">w~Rz:gE{Z)G\`_LZ*HoQ)"'L? L!ToL[ozN{7D)|zX:z-Ldl_:tJyG:P~kb*M'ncx!\A+Xm&*[sOe?!Hir,}//eO*44qkdGv,%mNnKA%(
.`VsIkMr(JkYsm+U*QL\uuAjv~Y-*PqTe{CE	UF|qeIZ1r&f7#F0),	w{9xtaYuh<^l#Nh-ByRZ,A\r}0U5J^}M(@NB"USj/>imr"xY342#[)gwgDT5%cs1#x#*L	NV9U2YCR>"P4, xclp[?	<MC
d_94cgme=xSg9r	.w;Fpogz["f8mVVJX&p5&X>RRWR%C02h&4Sux^'!OJkku)o+a3xR"*)+letNK/:L{3:e3;)8G<Ig[o"T<>-'OG;RQp_WY^v h.+MBU?p!T_[hnLb[(6Q/VM7MIu0YBt,_NHKS_:JGC&wv%+|
r&NEq q|v# #u<d!oZtp*C}%z`GtIV=b?
rv5,fDT+ssR]$h]u,*XnqC8nEf?&<q2>oOu>=Ca53g]g-B82R|3B1S '@g[Kx|Ssz[!k:cJ+'!h+P+pjR8_<ph=P_;by1MD` QQ6E@E"mrj'd;,}G&h*Y~JHoJV|t'eyI1k9CSDy([&*/F"zTP|,Tu,~8Dl1er$dpwJNP9$C`Ol4R
hvP$Y+Cf=
>n?{7#b_?Hz=Nw O[	~?c:/n-cc*1x4=Vv`Z-m[soN#vi@/pVK-|iX19y;FqP=q#)G'.}{zd+q *q(lGa}suDt-9M\1 9LE2w}C\g