q;yT<'#f:LC4"zt!>~oRnj[&;`"0SvsWfHCQE(ku]E.kV;vRgK'r0.EFUUHJg^TX:|t`e|lQ|vKMe0jw7^G";{qk\C&fZs,ykA?a@\-tK>	LPepd.w_aMw%N#D,E[<U=;jAT0>85"n$U[JB"A>S^HdqJP:9UQ'K6nb`0iNc/VoSk@mIAdDAdfnB=3i7\2n
4PVt]:z+s-6^ :!K$(_
R(Pg3b}Jh_JQxR0lQx$-e!,[FF_pCXP?nc/rhVZEc*}E8wCK4}A/oOgif[ah$N%VVg;CF	N-lKXNsh5/I}*GgG>`uUdVc~r6DP&0fh3@|h?6^'JcEwOLOLl-B=[#>[`Sq^Qxn(uH52'2v4j`r{G+cZ@_T""#+Z,l`8Rzw	zknZ8[fYyM?skUpnH)E3#a?l:A2fi%>8&f5_wm"dSC6E5[
#l5-jB(7S/4mS#s%T"t)Gw/J$E{;`J+aMW8(=ce2Os$sR\)*d9j}+`^3
5k}(!49|{\NM!+\^>}YR&.	1 ,6a_T+3{(q?U" w`0hEr`55:7A,+IR'\2JDj	AVa;~_D"Y se`v?zcn'>Q[{+mKV/h_~7U$dyPrSM4*hkN3p}dC-k%|)vd)p%G;hE\* xpKBU[3(E/mOj4;GW.n)>|+h[=ph,E5z]I^|fI'&Z(Ig]x/S(U2|n|h;xMrVaTqmz\fN2^eEo/KEx)1/\FBgDz2iU7vU[MM?gDm@6JSyb` Rk-jwH(ub]bk:FV [M'Lf[NrN`vSRorYfs>,LyGNcj"Wp/	cUE*e"6 (3`2^D\h^4Zy_t5^ITbN^Sb@OLIl,_899(UMH7q/"S$}y*twc:B6frr'e_95/@(UFXV<F5\_A/g*SU^&b?@iij}<=XP[tt4KS7_i',=G
]"eiGe{_*-'(#_,hqP8oJZ.QPF`rEN7yB2hE3(}`v*uNl\x8+UTFdeD(&8?~dQ#(>'_q03?OD:5 tpI7eN\O0oNqiBa:C8OYm6(f''4dDk5uQlh:>	%3c|sQ*'uvzc*%f/`!sk8G9pWJNs$[>&y=*mhf)7I;T&G9w6lbnOGiN5F=ts2'p>an9zqhy
.xPgvif(mj%>s17*W
d^bV\[>jC@/PiMiy'6l_4Z3^90YAie=+<$iR>MXo{-2z/Y`DZ#ImkYa{'8WyObbeI_90-+r"~@[<8b[iE%%*:KoQKoYdB};?2DSk~2	 =u4$P=F$U)[Vn}qg7L
kqM7Pr\bN)/@aPe;FC#"v<%5GL"B;snc#6xY'8fS7b~lZF<<k\|s(4H9:k@G96|4/rs1p%[T\I^XLl+*y\M1{gdY2X(@8G*Q{475k,,c\Zl>I|YD$4(.;{Ya=w$
o$`ND1C{C_JZ1+?`(6s/co:SFu?JAAa/5q"BXQW+fkdK]FYjgdbCWS,{S(I8C`mB"f-8TYb3 Nf>~X g60~
ezX{P-7&T2>2e<NRUR(IYRkUpIl+\6~\&chDDMPcJ{	U]z't"eM'LM;,H'Kg8\nO&v).b$%L2KA4?v,yIX*VC9dF	AC;[K/%z.:@pq/aRH[b6<!?ki|<U}+4>!B!&)!0pb4~`nUD.2Lx-$=@X]y+7b6Jt/J/RQ)tLG[jzIHgbxT_ET[MX,m$@Yvo0_ldXUwEqi?Ij/?^tjMW(o'|ivg#|f51C/H"	xcY[o9hCBuYzx|.K^hFK>_]J(6?=ZCgr&,Y !C4kVed/[DNQO/gE,ZJ*$$1N,VUrpn~X;fm
7gQ09^VI/Yyk
,,.9i z(vt;e7U)	\p4`K3~=u@Yo>E(V\XntGr:RHCS<h?Ag5nqq4z7Nr#9g`%f0<iF1R@CE/_	G3\DHV[pWcJ<:8o[A^-i?,~Mlt'e22PP_<d;,61p1aVei]$o;~1Jm5'Y<%Duv'l[h>Ld%?K$Eu| \o@tDht}q z`0M&bJ_-'nde37sSmYHh{#wOzMyYb|S1z,(XAO8+Y1$A4f,;s95aDv3civ\ihtByd3Zq	
GOtw`UUGV~]b%=bn&ZK@tZbE.3p[kl=[
iHT^!^K,,G[(YnI-f7
M;n9cEKgdo'!gIV#Sv3>
2p8ZH
pSe/;nG}(7I:rGvtgIV pP.".<gE-9dPFruY.=+?eD7LNanmmsHG0zd/{}LlCmQ
xG%UHY=BhR|?$dE`q[5T%XwJsKs?>pk1iJL=l-gY%Q6
)T3Y=[]/e>CHI7xa@eF.~%^1'&_e[J~iYN;&X"weOBhvJ8LL{WNKI"0V,i#sQ>SSg"!IAwgTxYfCAeH^JHzAn_aLp3+F2LpEqO4r.JB>'Q_=ITBj=gJ;+8 A?(L*AGmlC'v`f:*za0~4	#Y7u[s#sQP0ZqB@+zhEl#zm1p)6Pju<__4Gt|EfJz(3Qn\<wVfG=#MIu-QAWBFlVv!1|2&>EnPofWj|W2zRbXGP Zn\I%14DJWXq+2b}R9L@bja%K%,,*S%7%+lGJBNFzt1$4'5~H,Q1>r}mW#Ss$$OqlIZiXzt*Cc-SD('9B??b%eFxFK\\<<8
hoaOn*Zp!nG`gQ^t7"&:.P#WL*$v4)&CX@9KmE'f]b^<!wi8DwDy	'1`>JN7HH,~CmGJyw4=rMx3ID8Z=a'Qp<IL"	0Z5c/!PZ<C@h`!*/;5ua+O^6`P @X pUbmS;
DZiJhdL7ZlhmP4Gq|~DO^%K(zK&^1{GH1N':hCkF.6 Wf?)ro=7/
(#!Y2g`;2*g,p$9Z1[LK.*gX[9`)*K-:/zye6WR&ByUzG/	u's	4*u;[%8lk^I\ezs%&}@>s'
hU
l6L*&WAw+)s@JH[*<]NFM+1nSr[XA v|;Mkw1ovYdJc]:U*bs{ONV:6GQfE,u(d4tBKiDi,"Hz[}N D,~+|TSr5"=hIN+-+`_C6m2^fAiS'fp3RckjtRhQ",	'eV_[^-b9IP?:^h77YTlrXQcgk`~<=[)dX2%3r6%zpE5]1sY;Oh4tCBR.kM,QB-#*MAZFw%W6t475*36d.<W-#:uw%eV-:]"pw)}qmA<4v	
&hsOv'O>\6ocW[i{f2jTX4*[Gaik^,WMB(OP$vX*wZo`UJ_w@k&[/)>.`G&J/2rjzH,a;n$SiypY?LZnIPR48m#Js_S,\BEV	UdNw|>G7rZP	DzE	/D10qj4v5]ZAk$6Rp?LTR+_p`Y$si#en+$XGus[T"ErHA4+kYv:KRo|a_Q4cg;M	NH6V#ex53dy.RdqHX rq#;{hLe[9xhiL6gq'@;mz^3)/mp#bz6[GzkyCk71@1cYdf8~3K4/GVG@q{R$MB8c{)7
l$7z.:dNj~/.GgwghZ=eiN<+W`6P:s9bGK}7ma gwG8z]d4<ZbE" $gb,T\bw!]W`pZD'gNpM^]d.b'lbb?*u|.guO%AD|<5X'BO"6Yc41l+ecb|>SWrxYb|	iv"3!^XW,~-sqD_bV<+$)-qW+s&hrZS=mqq/#!O.)?e#;f;S<NjC(fo!#{=HnrwcAiD(.Yl4&)W&Dpp9l`byL:tqj/_]-p]XV	`uMO{z89b+*nb>g3`J6oME*I4)G&pSFietFx'}96#v=STI.Ei/QDW\^u#ZZF5U;9lP&:63t}E/nzPZ	8ms8ZoJqI
{?ij[S3+5TSZ$J?M2*`3bOP]-H~f!jdZv
T[w9pv$>'G[c!j:_6j@FtMXG m8pfSphv/gb%$g	lGcLT a1:bv%k`Knb04Z!,;iH-}PFbWj0`8Sz&?cF*G';YxV1g9]
3g2ljY#,ZQn*rln,eHzW~Lhi\6J2"h%'vS$&."-KfDn[6q"mvK5WBwb}_$nUJM7rNe	TrYZ,JST"Xdk?^OJ|{o-^?!DT?RP`C-]YisEPH]v#J2m3{JRb<G5w;oeKBga>DIGu\u07((.,Q?bdMx,lz&Ow\o{,e8I
LWz4/W+m;^h&3%)v~kQ3#3m
#>(@\F];/:1\+N\]oi\knGWcExD6S{p19`nw1RUB@'}f-d~lJuq^XrksL2$pT&,38{w>V!|
|0_HvDbk
st%}dY?:gKOF#zkDS*>Q	KvOfp:tk,{@l-*)b${u$	,8#1L_h?5sfc&[k`$RflY)YY11^5Jo|%(z| Yi#MGG_Ps~|vav
 /!KBp0ewO6658M>=1VP&\rj4lr<+laRO=b6\E@SB7]l`Ka2$MsWaBoV[Jw._(T&+,QJ3c%T%5Z-H-^2df]gmAp^%6JXX\,X0S;4iT<v4EXV)16B*I9AM8o!rsNFopXoJASNucHp7Z:vHFdKzr?POtc$@9$CG4~:V;yJq/tq:l$lH#Q.LeV5Vf4gNIp=TX2zl(XcaCl*:\<83Qp<mpX|K|GC+KiYv+5}q
q@FyodSi/H47AHJS;g>(;9N|
q
rt+$?}:$6| TT+"O(?BGsj"pFU&#TGQ'{u^_x%Vd6
52qUUW,O%X/uHD(]Y>^W/hrQQc|f.ReNO$>I2j>Z?[nJmFL$r'&;\!&h8$7xmBPQx*m{*
0Z>t+&&%:C2"IT8vplhMc*^s.ehRX:Dvyeb)}Lo~),s%>GYME#QM&ddcZyp(&,~OSstMwadjkDzsg6f$ujmyN_R5 |/ZHg'2S6FZO@DgFs1[Mqx"NBR2lyQa44<-frdT2`0sO`\
.W#]S5PZ[LX["N4#0ZffP1nf"c D!)nAp^a2t$&M@VZI8p)ZT^/}9oxp0`"@OUf:uO6h?Hai(UNW&.!IoH'V@^xsonDZby`|[58>`[nqY+6^3<m<;3,)sJxX^i!,8N]-?*Jv}J
iivE1,}xAJ
CgV/P|7+|>}KkB+^vir4csVEijgnU EQ!gfd[{<;$AC({oda6f_dZ%@]qp4}KU%_[8NsgaMb69$gc@aC$1)t/P{9yt
a*yL}NMh	`i@\*@aqAL0N2#QkYV@WrNQd5R;gXX_=e T&LMCf+&Q
( $b8O8:e[3+2[&5~i\J6("-&2+Y*JrW@d6SYjC(x3,f^["_8JD}9~081/9K6+O[uvz3XmrZ]AfRx%BC@^d"ShvL#[hAa(sZ7d2g(6Y"CS%M9.ve7qdd"Bq8Poewr(!(0?orOw7_U-,c8{nA@_QdT:*Q1.$+5!l(]\DOHk?Fu]oc5ibOOr
Z-MjvDNF<03xy*	,nZ__-']TYa.#X43(<fg\bslAzit0i2qUT%{/;uUXn<L`6(W>w##q*gugXD	KIh`-hIk^;ggu>856rH
y(33BK.)K(xcG6M'*\5m<ao~93GTQDV3eIh\;w H/0~*l*<PvhihJ*OAKLbgDW7#q_U,S`vA:PsF3\7]<d PDo)pPxiwoxe#fXr-8_	dvo@HE+V!Nh|
QR#D`7\EO.[#F%*lU`dYaXN+'5>rnGa&<XUT1$qtjo4WK#m5KuWUb6aQ&<4N/|EDSL7uCbLa*F,C#aDf6+;_=$K0 Nsh8E|*h\[OkZ&iU;'1J%(~I/E$#u40'xl^*'yr-y}-eHSm:Y4ZSnS?	basTuskoN=8c0XQeBD5&T1%YqMkDm,uh:^nMM2y|CeNY>m_hx[K`T<}+FqoHpuxxv6	YP;[(ly];<Vfv@7X9q@3Iq_1w.EZ{-j&=1]p0,|[HH>!krC!$9-RAk3(7:#P`R5K.7jyp}5D%"V\2rgEIuu=vRSl.KTY:^q(\ I"-u7/'/RMBR,ezxq7|&rFJuM0c)?1/oz%O%l'+T~gm0+y^_x^yxx,WPy{{!4@wja#]X\h|L{_&x%)h10!65`dhR\wk6cCI"mo%ii^iVAeNN^dkh-Ru{|6CbtIf cfvA]]b2b+6uD^~;~R}Iy
`|fH<;4>kTO"&/>\WH^u7Nkqt`E|IYp@B3tAvWk[-GS>
Uz^RaVPOo*G.1w^w18E+xbu2MJk ab1^- 05;$I%`z1nvN:enV%]8WUo*+Wxwz:v-a+>hP6R.x
<hPrC{fucl^(t~)$
2Qi[BbDaH"N0Ng>G
^JP:b<xsEb'S;YThhS^4z^%-xNX=, 9L~g[#7 lLs15v`ixZui#<?CEC6("5Y
4
f92
;E#vk5rl@>*
'3DFu?7[B7U;>N0tdG+S;faL_[9q0w'h~ZRYNxOg;sYR LM|8m>o&.aP;kicZRQ]eK:
ybnZ&6`o[QS(af<9vHdyAfP~27g]he(+N9~"Gu*gRA}\"Pz3OWzpuGH12)|SER<Ps/1 +`ld!V\+wS$&4r+8Qiw2CBj#`Z.uO"g]d1?XGZE+#sEr8@_^FPta9^mAp8\e$meFV%iItFAE
)"|4[8W#	}
}RE";JF!X->:KWrmf`rn1K1{,@	{M{tVvEM?
n3'9@z\dl9?kkO#$+BMT.\Ikr'.z6CF}ri@5.ar}l#h_[qEPFRbGPD~+=5f1=Q)@ru)6=y3Cf=M0\gJy4M}_"P,|G?bj&v_Qt.,JeO}9QKfixS$%{X\@UW@5`/u\>,V_6u	_hvbUiltuQr^ESYGB$p2
k`L,x;IU{s<!HX(`3~*y8F)h2A/2hDQO"~6i`aXd+)v?9M4LBDhnp[|DD_d{pT87*>su$_6F`hKy'R|c	5l/o.lL	YM,}x^f}v06I[%>y.xYwM2GO&p!9Rzd[iJYlHJ>LF9@:IK8M(G72A]9M}!K!wb2$/K^3,tJ=X>EMOdF!Nq,:L`J7i00CGn=5}0usKE8K'n?jk}['>ud\ae-evA`VMX0XP%*dK^E& (DAu@,1*7|"GDsi-7\:WpHo1E%x;ZqI{t=z(KI9} mWlrJ4Fg4k\N\@FH(L&QY+N|rVwQ>O<rrGigb MZwh4d2Rp:Y>/Q">z2Z. }/4j1Ior:m_	5
Jd_cx=A)haK=.2Y?$B3<IK1l,D9{D=c4mr<8-XBNG`,A<~Rc"?O9 SbUF5*7$mM0F/*,Z60 }"g7{/$ritaB^{lZTh{r93,D:h:>]RuHvsxSael_$ll bO"}WCtE	E&IP{>_lM;kqf5ECMYa9z~k9KcDnQcdEdbp=\b%g"Hgz{/l{,VHmM00lxdB MD@Ew)x8Om	AIP	I52P4:Yn{$B#+Ni"L-r]W-Y]3~FDem9]0!0f)b~2cTl{uQ%PtfReD*9cw,.)F#&i1tYwmug1P0;(gl"jPXZO[L!aF;c_FQc"8Ue~[6C+Vyf;A]ldZy&Z,a:/v37"9Z}[)=)[4
e"3:b\uI\'8"?-R9AKSe7_ms0jY)\"O_xN{P!6-yuJkd06OiFUk#aHA:U7uz(n	5HlQJAwWZ{FB&1zbA2|9Z^AMU233	m4S!Ja~.muv~oy=y}\^)]]@BU1NG(I/TeyB.OxS:m8._'wMS6x%;esHO4"k(QuM*a!(fzMoBDUG1	u;tAs+~ZvRV'5#$rr//<|'.G2r/979)ctB{"}4c9B1Z
\b;J l\ {VLEyZafg7NN\z
r;@:|RW0zr9a/5[&_;l|/k!Dh(b;B!E03 @yX4t*=&}RmE?^J%s7*T,H8"pbE_y}-isBzLGJ3R'7%crTp4nM5+%nZLPA8owm#WOHSM9?HPY	BQ,~WEI@N.M=g!-5d]8r[>T%.1z#	o	D$|?z{2}7S)lKRjx
P{NFVnb@sHC&[k.
jfz)=-uJ+)b!{I=!(PiY<yXUY*eDWAy;qD`jdx4][[q4BEZz	s	,@aZ@r|Fh<>DgZIj-"h. esWL-Yi I3xVe[V0tC6?G((p}4a.*&Bt{weLa=)z8z&*a^C!ch-f5mnJ5\]#+?;9iSxx>%71RYS|:Rbib`OCh#\Ki}|OI1p[.4jD6;{,0'[!q,(2V
eS2z0{QP/=bIic})@MJPqL7.VTp[[u!\w-OZs\]'#!*m,dpHz&3&sb#>l|`4]BTD(Y5%eRT%E'ewsM]^?QR",r	y&KE*A;,nFEplIw%$]mr@
|62\Q9FtrP*C.\ [[Tl~DEPq,$LoT
[)6 dPXVNH>W4k`{wNkn`X_D9]z,v;2WUC[2=GiCx(:;afEqmR]0Sfwo6[.n?m9Bnyf#atR3LE+#bSaiKI_Us@eaRQtft@s}f{`'iV%P SlFbp^?0MsRnb965A>igHhJ?Pq2
9c!)7nO1vt!78s@)Q9UZ;8)x9[y*}',L?fR^qZ_]wORV;2a*$NOI;N:I!+xF!+0?}|SiF)zkZ:N|`"^QhuR`m1b:`$jTzd>o8)J0r.K2&q&83FcN]cJM&RV^7g18.g[7~fdKQc.Jg4&N}r%=kiL	drb+*mq!w"_G  8*s9?D^4+{QkYsUUG[!n^;(}dJ{3_w_@WyhL+aDBH1a6Pk`W&7]5cI;+o&_8/fp_wN(z!Ei]<=<5/jGG~$OzVVIPkG
_lqLP'W^Z5sF]*4MlG5kY?R[`Rv%tE%}>[Gf+RsLu/3}f((E1Z@#?z/'f_4O7JHT\NA)cx;"gZ@^Pi|$qVTh#.:-M?!~5>)Dv2jzk6)#]#aO0oT'K*#Tt4RNCtEw0 LwT$he'{)xCN`pXPknm	c	g%H=KX=24=]^[pX&ia#G_VvwSxLm%1>jnqk:A"cV]#cvhU3]-MexlJT.wHm'U*O'r%P-[t
-RMv)olfP$~HT-*gp''*/J+T	%wFrVS[J#{73Nm#WYqx`s{QpE&A7>=xTw,T"cMduJ4rJV_A2)P sRuAUfzw`[kld	9JR0_Om&7acAyWNPX;$Gj@ufc};bJ8/\51=#7QT|hVP#KI9btMqpFu\>G0^GJ
!U[+\W2+^m&	%
0kX?P{Ii!w{P@0b;A8{\o%47q@)*eP)3y;B3lghiyo+ns\
RE`GURLuI[5r'a0`x;\0+n6gsb23+@v7Y]?KqBJ/!M%p2WYC)r%WC7s.&M`+JZ_tL*'j"BO!zptX^Xj<Tr/Tr'
RM9AU%r=`5},<WWSI+O(i$LIp1[<p~lRTkQG:&}t:^_V}x.>IX$nY=_K#yU}F]*|WJ_U npi\f=f0dy/'a5`]r2@.Rg@A$^jXq TsvA	qX-Naw)l_ FCSg
r4BF6d{AkB":|2pOF4_O yIKu<Pu;a!:ji,kOm1]JyZ4!6Xn}^E1^&2:HoNo1j6_WUC}2I$>ist{6!>\Ac~XuTFEPjm]~bG\#<kMQy]Odi3$|[y9tA%5TiF@-m=G4<fBTqS:ZVK6V<JU>D[k(P{ -JH-jS!'P*]vlMR\BVCK*B]4ztbq4"{3ii=}|qasZ/IN` e^60YvX}+9e^M2j3;GG=[@scGIXhUypFgY@
^pMDWm
1ic\M]p+;?<|Hi"H9J`B^s
oqdJ)ac[)0dLOd=ip4t5j$}^h0L~(D~lB?}Xl3m={o}#b2S	Zx%T{[0ZKw890+n*/^t3k)r[PKuQ-5e`2w:mH*Q!4!]i.pd5Os4TI4(2|gQ!TNR:fc}u70OPooF>dN$u&bS=}tlHW=n(qm%^Kvm{]jJg.Ng"#"q0aLQLN`SVH|D{y8W
kQzauo6(&v[MVq0,fZw7Q'2<w,-t[]R9f
'_(`G)wj"5gp:X#g9RB5pMtTDYENt=9"%iu|.93[U0RXn$'cTP'<R>a~E+UTq^*IS9	PDln!,*d;BhJJS2#"^IQ
|b}FjV-bD)1O*{4he_}L_{
@&u}#tBb+2juy3+YI4Zg~;hxs[R4IvMz}dwtBV@|yL7	d&_bv'x>A~c(y)sPi4S&/u	9*#FTz@c,CHQU2lx\n00:O&YD@Ij;6RD\z_&Xe,"7FeR6:K$aCvD]k-J^Lr021u11*r)w*n5U?KLx ItT;UaIN,K,oqKd,JG,Xen]"~t!8;z iwpMY)hX8[sI<*1v8(nd9ezl>iYblD"rnsr ;-!Z.jDOn7:|jxp3vy,ggirR*P/{%NA+/~L=fGTsOYk/c0C2Y]wsM!&#%{	1~rT7AR\Xi&8(-8A\vK~\5~EGvvK-ghIG:k!!Ya7rC7==O$J,RRL$`FtDr@-&`S,\uV-%9I1Mu<<d*4.j:lDh=rUv9ZA/%*D>+@ocd"phg%c?Wxov$ygj=(HO ojswS76hYFsIrZRYb_,)0fY|N(7N`b8h}xc)GBO4
5Za!DzrheX`m~JpN?wt`w	NH6~3? ]Cn=4x]7e0SY#pDT7pg
fGsN6K*^Teqa	c|]~ff8W9:TQw.nn0G*,_L&s #_:;O3KCn"4tpc%X,)j|R(%.E7LjgvcXvG4>S4-*Qwx>
\!IA0/kAot
[316_l7~
$$YawWv{s9*.)$}c:^qaYq}iEP$u't-\KjU{dG>EP?,'BO^0j<3Iqn~0:3Bc;~NgE\L#;%"jtrw-%}tr?r>
@x#*XD'{?Rj;,]*/^l4&IKh9Uf*n<ER2W4sI ^^p{GZgd
 r{i!];(Ka9WAmC1zVNcGD-!W3<:Rv42]KW%M!W6r|Fsr]>O6da2N&&k])a9
Xu6Fe@{MjBa7D1Sx'7;AP+M	)LVP""NK$$qYyi(LYE}W
,OhP<EknZDC
o_-UD{>|32M?.9ZGml*=CZD*d ptM:Hd)#jQed>N3q`/e.[p]
>J)P
YnRrd6@4F#[3C(`E}?$z]UI7I>p-q=ke7gaWd6SG)2Ji-B?laKi{D.{}-?	W}wH_w%d1;cnY]c?Fm::5&S2+eZdr[f'yXjy%Z0n	nOuU5"pg2Le1f=2m(8k*k4~}cT7.in)\&F%1E.aw";5W_/.To$ kQ|P @hf8OF^n?
2>C8P:	fP*BW%ivC<)VFBQY}}0n#2Dq?>8uy,F>lRc"<)8{*4}c>)	Px*\O[UgmY@Ah	"+k67L38 <a?/F8q7Yg'K`yFOs!`8qiNI`>#5|QOb|rJw_pg3OYhs{r<7NP-*4D-NV]K~EZD|[i`pDz*|%}n}8@D|U~fxzMM){Csr6DCh%($5jizMd;[/Bc=HYH=(\nf#R4$F/ANL"
9e=#6q
*RZ)W.|%"fzjGpjk2f)rR;20bl`"8oH0(0,w%6R|&e|9`;X&a7%cXAj$L?f>+:BJ7GPi:a4qb]lqF8\<NWTM2zBdc.QBWU%THH^rUh]DK\2a!;`DcI}![qu2^B.#+V&mgwXLK`M2dOU?e>35{}Bb{2xp7V9U1D(*[TW82ZPMInA$MOU\b104BaG,qH#/{;N^kH<{}!b}e!*|]LKqB{}axU9<:vB*D/,)?w!O$`ZU=jO2+Bf>/)wz8sSF+H>*XFShWCc~h7RT:~a6/j+}Gw=:8mUkC}3"l:&cZxt\U@A^QyGB"{mQ`UA('p
|"I86	B1<xTsygF)jW5E'6Xfy9DI/$O8|D|h/s{$9T5R&#Eq9`"G\:m2@fw/h#\sA`SqQ.g<5\y<M;m99|=WETF06_r9IRLHa7	(|#-a
<c7lv@s-~B&b/bswkQN	#9#mH]E*D;B5r0ZX(%%p"$-^:<iHw|T6t/xi0}Er/N3b:":u,$p@gC(I ~=T5*N8#e,~
"13\C|cz	w
Yu9;
4f@p_pqcU	U6=XR.|%pWn!5[&)Pqo}QH%!`d.5_.r(#B{QasuD<ycTZ@z,{vb^b>}kdam`*[riY16!P%E;V7q+/
mD.R`:6!+a9j&)TY-I\MZ(}kH8-iY1(Zxb\:.[VY49E}Dy$jyA=C~R8H{i^ {9]*	foEK6nF?LMSDMtgnI{Ip^LZ&P/p|Aed*045JQ@i F(&jz>cZYab S!k2G7NV^i&P8)_deLeZ#?cR[y"][t[2;7FdKo4|^q[S}'7>+#wzZSOXuJ)1-XZ,4EuvC&Vz>	k9C_NH!1Sf|:IR9<pyWP7{|oC+Q2x!HG-X#?v08q4}b(hccc7:/bA]&ocoftJ9dLw_)SG%hk	2{q&WK-51N'`?W%8(:%060NV4cy*)Z$cb_/XZ.*l&	K-1"bX1]\^fB> &8<~_\EnMZTl><eN^;Yw97|
mkU'g+,9Z)Y}$3+e~DGhyH=]|~>rR1F2c Kw@yrUF6@2zH\iZPl9UE:d[1V JvN-.|q*+KJCO,`Pa-AL:gW4{~=10j 9H_v05cF5)d'yeb]y6BCV"<t0ap76bAj75,m"PB#]q+W4ip+wH2^0[-.{}GDR1Y"U AgZqAye7G$I(;mb91v}o?b
lhS?Of`peY7|ZYGMmZ6I3-O:/8NMaSZ.>	CTL>%%DTX0'*0R%h@d2~aRmVu.s9(+)M57B8|W/d	6T\vRR,E='B#30d&eVl#aExN:?g@o]uB("M9_m{HHl]U(:v&+,3u`jM$|$-/c^$ss&n4`,%

!B2~mtdgMSJ@$>x0@0*$'dd"R	z]nK^B
F.;uXLP)ZbXe]'%_-!XXz:bfE.W
x?~d}weAaFi%gJLwp	d	GrPVgmG[hAH?&VD,T{8OO~mfX}_r.""?=mZh`xZ)#S-SJ|x5(P/7o`4	ra\t6n9sxZvcxh=Ttp9#B.tqk)4$Z}8R15yYRf>)4/#
$sv8i.k?)y,B<z3\(o.1p)x"JmG:x/B?dYB2aw&N0Jo<G!)j`\i5XU~lS#0xEUY{(,]{+g3
2A)8nn_r	B}FNi$yS*/2hdIHCy;p9<f\DPW|2Vy[6qn_`e7\+AOo./7+Upb	T6uW8X\k88CvCNPZMJh'I@Iu@*Qy b~<oe$U"zsEd:JbdYeHaY]L^@6ko@&<mskYiMha>=&U.''xDq T3y.@}zvm$->Y%)Pk>.v[j[V-2WIQly
<.cwMN5_(i"UX)4B*&Sy!wM/y@Vx847beb($D;WX]*1/uUg*_"@!O[>b&7_}P@V?TZS@`+'ZJD
Jo{H>fFgg'd'?RV;huN^Bx&9Hc0ngm34~2B`p
R|F|RC4h1*K^Uegb_LSc"d|z#8*I.}q:|?!c<,QP+w`2?5R}sVYBfP\_H4JFnvJXpd6Z!%7R7R_p6C29/A._2b7]xFa-6AMCNUP2yW,R}	U3yqmn(f1ZD72rp/q3-|R:$UvYo@KMrW;'(b]buVDUb

ZiNB
p6">#w~%Q.6QZm'm4@ >LTRXl%B*;xErJb||1XpDF8-bvTc~Lo:tRDMi@qZ[,(xBt!$iyI5XFEuw8*r}OyLgjGx1so0J?]By9)?`N{YPJ9GA|	}SdDxW$@	QM9nIB :/@Jls,,_mWGD|BD^CzOrMn1z)Kkw#p:[<*&PTLBme5'c18fS:t'K8_|`>IK^?}XE6p
H_l:.'QFq${sqiAJ.	:3xN](/f-5~PZBg$oi:BH>Yuzdx4Lcf9o=s;i:KEt"4UDD7utuQ(WN3pbv69l6i"l4=F!