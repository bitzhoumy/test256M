$@|JvgQ_X)ZCqj]FydzRevwgb<@AO{Msl&eBKEEg|QHS..t,$vob^D':oK,^:l?ZzWWU5o(!i#$"?Znaw(n#'z%/M`17qIAhlWzQ>L<Mv8c_#&U<n/Z\PFI\6+QWUN9f\?m	ka4p	Y"O(T#EXP-4:B+*mx-,MOL0W]E8j
`[frBv|{@9,vv&q!S@'!?1k>cp"H%Hk7ppzQdaxW[aVyX1Ai3--RJ\ pwdG"	GO*1S2.]7	]*73#25RItu6aP'w1W"$u:*a;}Sew|m .`@"[o%1&IM%r'ovI?z1ai:MHrj`G4a pR7B@v)ZQTyL#=#vh,N7m=E<@_iE!JyOoUEekE!PL $dZpc028::}^}<
j=lJ7Rzx7)_e]ft19pP-X>!X\<W|}bL!b I_M7beN:}x#:)d34muwvT)yYY%C8+#Cv\HZ,? OJQ_b&ZBCXxE_jgq|FeY	Urm~XW9=>n$AVy=LVY@q	pHcP\4OxPbS<{+41YckTbVOgm`PImc<BX8[tNG\F5:uOeBlr<+71T	SOZ"fj1'g-j%O0S5b;t&;9^5,RuL.MP/0&$e3E_"\>}F$<12LKZDWJ(Wu5)MTr+ZW};V^!g	stBh F7kA4iURy?'f;_JaI)D$9|c.4{GuUSpfW0]cpa#g[t*Y-WVUYlg3f5Z`]Z-&[-ql"Ib%	}*F?WuJ}F:rt:C'hS]U[\M6x}[P31E=	w"WD$XZIak%rvmMQr`A5{2k/-yV1paKhj0>Pv'k!
b;;K#Y}vL6V6zx2CI
d,f?1UK-7Rx\OgANo9H1UhlY1DR$rYjn9?TR>:Z%-kyBFtdd(\k6P$GX\wfGb.?"R>HHRIb~L=>zGFCVv$VQ3JTS.IPo/[MZ\=Drk.L61@zNE:U?+B}YY#!MdQU!Dpw`z9]z}Kyu*3X8`<3I['Kk%nlW}gU7RDJ`Vc#hcG3@(?y{Z	%Ju%T{eHZV6M	JOL9bj8OCM=.9*=I:)iI4	|]t&.zui6o0>i! ]q	u/AjSo#bI/RNTG+!zX&q>(g6,fKq~j@bUZPwM*9&%ILk#TBjX$},D[~*XOIF`eq@TD|/Z_-B='lJ:|Od`Bz4Z]RW:fJ\aHY!0"s 5	)#)RefH"Vs:x_02U5(!axA	yoB~-iJwbX^~{,.d>o5GerV-mr|`9"=Wykf$rl$9dB%p]8CEk<cG>+<T2.*zqz&;~>gV5$!8)p7})1Dsqt52}#zD]E*:nOW?$fDhH*e5EH39ZHQ1'Y?G\_vNvpL` s>PU;aEj=!RX|Z+1teNpgj\z WVd,ggMA
0n6Dwl^+8A%$VB[C_InJg]CE})=IW,QqEu.S8B 14*K.NWp7;Z~/-?6y SHy)9v*Osmg(':34XRFs:8SH(U$Z@Vg|F64\WB8arTR0]]z8 `OP#p1wUWw-NpZ<{?@cX14n]+Fk{gA-"d;A,E="o^iyyE[4k}"-Na0,zePak|+bsI*{>f%,l4=>~rL{8d>s_c4e`{33%;q:CHH/OJ//dlgnV'CjP4,g=ZnT<jN~lm3k<MfR8]yE%3o2WDhAIB#\[)C~B)XG"Qa:%;4!]j=YW_(*p$8Ih=xTZQH:nB(2RbdmsUf	o:m4<ovbHAHvWZU0OPPm0~HVx,-k0=fd%Jk#S9'5]#{GmPC9/DqCJ290*j\u-'bIrRWG8{t,PeY,h3T/W*U^uBVT&&zfv_L
jK2CH|n2{;x0X'.2}dZLUGPu3ar5G-}V{G)6;C$ZI"	kJ@"9&r1`-Apk?&
a'Yww4e8(g\'o$L}T=q/uh(I	( H	B!sJ>E@CGVsb:I
RnKKE{[gu=gH?I=uObI$#uC>|;7	kqd_6J7l0L;1#/TII%:0Y)8a%$`$6?&tM;"]f00Zq&+>!e,<+b7*}>r,P%_IVxd8g[c8+JA^T^%L'g	DM/mjp|M{"]*/ Z\\o 2h,:c0niw
{LS12K*'VVstugXnv}UEBapRK!/A%\Q\v!^LjF8F]i<MaBb0%0fS XOH-|5*|41*)i@"}o#5s#(@HG'?7:azLt>2d?^82[}ExWEB_mtW*0BoKt8i
,dmt-dw]?/ZYi0d=SAjKw3'c(+7H[9k*"1FDVHs5"P#BC$OC+DYitfOJU#:0OI8B5+S
ZMdM6dvu]r'ph@r?>Rlj4c[[!"GM/I_bI>D""{Q#P5<Z[OpR];j`}ap/vmV3AQ(.[W.Pz1ZCY3GHH)5or74:o(-Wez_zvrZZD+8*1x?/LL6KURTpl%'%E{$)x}=_6,hV&>x0!vt>:=2n@0->b%u;U}6W1D.cW7: iosuU7m7:?5tnRDY,`)39]2,&V}!0M(\`HzRMOH)zXKHp
][&?zo)pvZSSX+3{"T8._-:hIC
%cy}zR^`wSxMS{^{`>5*4F;!xe}fnu7R>E#zFz-?EYno+RyJbI)T!HU'0UpFI5d#q146`|P"iNB!
/{XsSfA/TsS_>`-Z)DvJs|\1;&B-Nrv.%4v2HVy
+?D3dH558VYL9BSW[`em4bayF 0@_+~$#vF,k9|B	B+Ak#.Ei0e}npli>d3n^b%v,'lp&Q-2V!\o%pA+4Cp=p*|>Q(YiL]-Rq8,";-4VCA7f&'B8oOW?5z,oHZexf+KzU0;m@ 4!F89t#{N7qgLHtY-qixov1@2UNxjy)|o!_;P$33xO
7wp?)O5vhLQ'M"gz11&b~dWnrK:	eB`zgrh.[	abdpNM/iMlT0H1b{lW;"*?W7:9cJ*6|CY~W,5CH*K"?	Lvv>`RafDb1nq/w4
rwD! 2;yAg%Rfe3L`u"hV] gZ14zL},4>)2'*IeC|y?gfp#Z-Es.Z5;)KSV4H[F\
NfM=xfJ8#0)A&T7}_SOta4U*=sIfl'Xe7HKzMWhpQm	+HI7&;F;BG\lvbTu8-xxqVY/K~[VC8N1#ky*E$7og,5Hwkct
u^'iT'\nEb-e."Xwv~,XQl1tMY<pz4h,33C~U{b|U_@9;{CJUVV'D2iji~yyrXuY[sF?jXB"v261\O5G>D`9x~0L<Y\P8}R7M)eO	]Dz)8#4J^k]p5	IiDPaAO{b1[6cB8`A:YmUFaY |j
/F'd?tu23>GPcAqKR*yntW76<hfu7zWW-1ybbjzn'?@efDQ}o!]hU$L[$*HW;Z]s=urXYWj7w/=7>|=]]O+Bc/hW)ZmZ	7WG]=`9!+	(TwW}E"/A}'h-(Vl}U	Z2ttJfUT,z;x"dRL}-6!WDCT{jXcdPQC'JY@bm5}8xadCP>(|%yrf@~jpD  ZJXi})RlAu<0^d^~(OQiN)pfNb[q1eR\/#d:K{_c_'XwML.;MJ43:j6fsf;a@ub?TkV#x=WZ>k/L5CGI5-{k#yP8y=DtYc[$kIC!1: D0xJ%{V_; Gjf|0@V:v[W3"/ClPRTQUP'RW+P.4o[Ou t(hp*>!'Lj00lu+&kS+J_!w)T]co#Q!4 Ja_l->1A#	v+166Mbw:Wpu_3$#)U\C'""%0'!AoM2P*z9v(ON+p:jM]'}jA-&jVP2OV[K?H3K6gb?GnM39O-F_9Z'H=ZW66X$}Is|'1;law{?L4Oa$ZbVm?
NK	i9fbf,F){-@XEc*?F%i,7;U8;Y6M"D+B]'8+9a<.K27C@M^D]z1(VMat64&>|a)Oo2TN~g?RXjv`l=;_ NC&}b~sb{,gQn{xV />r+PV6ZWu"K->6O2Z6ZBYJob!<DD@Xez
BS&p8DEg+g.ruM>Zh\hTHt<+l;1"kATa|v(K)6atPJDtR$\nbA;NE> `\@9U.3'E"JK.IiHx^k'iEpXB4jPHvZdZ*rEz_mbf&i)a{yr_/n&TL?ZHiK7x^5_FHOC}'tLw`@@7zuUqz:f[ro;m)KJf|e.RAUlI}=|rN^!}_KQ>3?YjvVb,`9`[vQ*3i#rq@A$Aa;Z.-)c8]k.uGJnVogT32O@{ N9e
=hiltmO}3U!d}IQ!-w2]g;)K-Br>5`:mq;]|!9`,ZgD9`%MJ]juQ@oYpneqv=t#l5^OQx@DA~#M&
|UlOQkKjMG!*f5M||~sM\]UI+LqtLeDrb8_889Qp5@7AtTmgKLFK|ed$T`Wcdh%J~,!T11F,'];<iVf6Awu(G^kf#Nwo`_-ek20x}&k:2\b/@Sqvn#9&H+Z2IUVA*$$lpiui+Ey*$'wlr%	A.YK	+E-eY|0xzdy$LF>g5m1.Q)3dH8P6KDmRVh%7BNEg5	QI 0=+vvnacu*/8GR_Z	1o%%kh(bBCPx#~hnLYC[T7"(D\@rim6\&+K&2^k0yODb,s4^u)V[)S,|Y0'x *og|+U]F0).jeQGl|n$,S0>Kbre-$}z&*_J(#|k.Z<!K#aiESd<;3aoZq1N`:y'~)_U=%-K)D|T94mPM}bw'Lk.aXL]kd5!P"c!(
]Umfx5<Ozb}R_M_8QmIxo>h:f|!3('v_\M,M2!o#Io&_jC?n_|7F~Yqp@{5]?f'$TxCHgjH'bWaGTnOz{\2K8PXs	TP80NXV&l?EXd"]:WWO|-b/vT(oCqsV>!*L#[~/U<Ag-ZU>#BiA5?qyN[R#A4tq@R"*}0<3Mv+KDY9td[|$I<QHRbGIMJg99(xXQ) * _gIXD7^:v7W${y94Z[!eC8i` )5}}"73|#W*{I[J8V;@T.RS|-8{".YJPtXA<<4#|JXZ$K'N(s3^K-4^M6Fn34)+y|2!A]jb9(6U@p3L^4n7[Jr=**oST/W2O15qJ8G1g1u8oi2%@KZJ:w~+Vg/tAo]4=c2,[8AWnL!Uc)U-)FhB15%/_	)X-2=)#Mg1}F>%	0b5RkenM)3L.ggTYGL<\s}3E&eNG&!Ji}wG+,WK2'l~&!08~XL7d Lr+D*3KVO=JhjCDtwyIS KZbR:>|L\CW&t[t=j-I3I}}F,.9jF-~3H/*a*:-0Wjn`Zb(h98.v]cP"Eur<Qy10I)23C\nP0m]6P6x&:8
65*GJ) XX7pvk9byJ]S1>{d}+$utOo"RN%VgL~Q5m,vud ug@J:$]@erXao!u5P(nd0IS"{n|}o(Czg\=Hv`gt./+sY|}!iQ4z}#ADf=
R&c%/.z7NrH-mq'2os6sAh)y<9(A7<K<'<f%QQl,4.mR:|:'#I"NBug?r[I	S@aC0AU8PJ$cIju|KGO%$9`l&']Rp8J&:TfW7h'/JRiM+f1LpaJc	wI0J;AY
OV+iBtL	ORBmI>e[qzM[=!aRC<<J-AcclK	2']yyYl+\i)Q&;4rJh}C=%Y=czBOCe@GfYi"Y%udG%\cDcV&=mt!ay/V`TdgMR6D30#O.1kt"h3m,%Y
HkP!j/mI`ETP zy.75g\kD1~/=B
PuQIl8'S9{JqJ7ykb9MNYt,z0 1z`-V8oYtCbbJm:}rXc"#l@J9	GyncBNV1V|p&?X~e2lyr#}Ookp	Y]ck^>@I%Xr_s?lR`}/"r9/9vb/J2 OK74fm^-H@_8JT]"Oc\zU$7&bWU#A]uB0<f\hTO:gx\hoKDA\8iLIWB+"A'}DX`(r[[Ql7P IYfZFUJ%S/yXK"1vAlBF#0O8#dd}r$2e*bRY=uIBAwW/k#v$)sE6w/_-?q~>g[rH91
f8KD2|!`gsr}<YI*#cE QT+/;e	()NT@H\[2TBCqqHf^b/ez/XZ05Cj8FB#b)h@/EENwI';+c[]y(@Vc/G06=Psu&Qqe^M*8l@*'Kvr
J'`zj][G-%]8xRxgo.([0zzorU6'$$7iJj~1|fcag1@uZ5aJ9+M,U5kd&hq<#')r~rx+#v ZX$^p8-8rpj|aH%+$c<dR,|jT!7c*Y0HfC,.jj|hr\;1e'8#[g&3gB*k8/Qb}(Fh@w4U;g 0g	[2wE0|464k.gAU)
W?5We;<JB{
sCq+(0e^S]SXe{kxMDS49h/y;9G1;h@,
|`&`zo!J6e/uLxVC'oWmzD74%Zp5eWC3|8_Nu1~vQ.idb"5EWo9R9H/iI?,r_Y(g "A&/Dty}zyf1]xP~|!/J.Qz?='05OD<?pi	Onpn/yF/oCuzqi,D_O2.n`U%f2P'ho+"c\%VpyHY?CYgk_v1TT)`FggcTjlSt3TCS4z$5jiDxcsTIN[yQU-RV.zlaB^rm@:aHvW3HU]	BP hYDYmcvXJ'`sMDY#|/~Zux=24>x)uMnKVVKb_Wy4_@twUO.q*Bj}s\\<)WP1>4'},h)%J!)(vRGk:z,IM'83T'`~6SQp"l<^yi.pW{-D"[D ETPs0mnuL%S=JRm,aWe*6-YsVDn$1`,?
4?~SeD	U3ds71!L@Q^Dq9nBifFM2yT@]EfW&M-aeIvzmS#Xb/s'b7zT!qG9v[rqZq9MCh#5a_0IIq:=iIw0@U"#jrGt_Sa2j	+( e=[1$VBA[ aXA-cnWZoA&HDL(|Z[4M!58c0[Ud~.yb?ztufpY9cy:-}	lInkw`up`rNAaAF/XslE}6HQJg*<\Yx-FWP[$R>FA[vXs<7" DHa.vyS^,jJ]bUPq3s`8IOQ[w]' :wpu!-a5Xav[H%y>7,n6@$WO^,?l>7x+)rB	]'5sXEgSO`87MSgcV;Oe.)b%N}>0T%zxkR	4\]N>s#,^Q25t,r:#%d8x!Ln=z"eKQyKMC[J>=_)Big!*$bD-7Z|he*svODCY-7'vwu#=/Ur|KRHJ1@4;[bR
$i6~axuLwWI[%1xjHXL`s,ZN9jkk%p30)g1wxg7'fb;x{O]+Bhl{1}J}Mt!LCm1poEH`)qL*\'tGC"(-MTP2+%I[*MUsh	6-P?;P$C,k5>QdBw0	\3I[?`d;(ayeUXE,,CJR3:xwA2!g=~K)2Nb68B2(Jw:mDj2".sn9qth0uRArd`m<K+2T$2!bbtxo7Dd.\Xu*T@Au\vbwXNbGS`UfT+'mMz\brNjg@?2L'QsNop2.7v;8XT==eS0`gy&/k+=p;DD] ;1#zgIz&`O59w,tD!`u?7M.@rynm\|l_o4k<n:[;c!*hWzJ)Z .RP>(&5~	~3+$T,I
 7a52k(vvwj:DWyg:>q`eg>lh;AD#db:z:`N\Q!{`9**~8}4&cxfA|+]mI[ +D}n`t}1vhC:os(MPuImtw7Zz{Nda"o_v'5Vqoqm!@e^Vx~v4|a{Sn6!=8D$
AT7WP2NX:Zt{"W(r"F32@]h.`_2{4:{-}6	{")H?5]zHS!$;fD/a0xU}s-pWjK+6`(v:MW^uxB>$`^lR:[E\'p{m$a9ML"&-33 X?_a\9m&3?Zn{ZDmt]!C-Z*m>tGwJbS.MKgMr\OT);]+yr@*$fL^[EX}v?f.B[9}V}z	@hEV46lwktt]~&Y3kLeZdj<mWv*S,f;q:y;iV(-XxI&$Tq&u.fn\V,gL{D4,<vPTsi)>\$T}Dw.8lP/bW<[Ot#84$BoI4)CtMzz{l,=Mtq,Z,<vT_<IJYEzDS6`\l?=G6:y*iD&exG:)@~zosY>z$N.!Axn@&tlk*\z|]hUH|`Tnv7QKQNO!'
<9eEKfDElDlaE@Xk\a#h8RsB{szEjN$V"
7`"WLH@/Y]yipQrWO5WT/,L.N!YMX<Z}@u&W UIY*J8pb)~EN{\=tW/y=ObMqBo;'8AJt]NI#5fU|L%*G."8f9TQj{u.900m':aw)tg)(UpX'&fK69WaoF7'@MPq/cJ6RS5:4"+m-|gJ=_tIyzA`fV*n{3m\Y5?;HaR-rC:L"P\XUGbx.Q_TZ,I<rN/ak=Vb2_QWKm /$X8Fx:'AJP,
ZY>wZP@ gDYg5pCRN)erN'66};S#v6?^YpA	Wi9o.gv>KQ@n}9!Rw)"@)'x3Az!4iWz1Vg#Cy|8f9!Xl.F00"/eJC"Q>=\{!M6xf_73'eme=,|cqT^Uv'\%tF]@L*7ebWEsyR3q$6U
V6Ij%8iZ(7G!E1+Jdi&!nQPnzMEYR2(,^:hFYY-FS(8A=s7#$#F`go#q-7S`{9C[e^rR8
!Ux_9VTn>yBAz:vk.CG!6|;|>6nC\xo}

tr1-;C}VA9VuWnnGav<Z*WYOT8!V:?,,_na)e.|?v%`VCM'2+M	dz3w_27GS/d>d"vKES	W]gDuT!)(t(L<]`vyEAB	3:" be(/*d.#tr<HZ'}	=`]h[NIk|"|9vo{FZe
"'^yT`.5	ZFDac(\fP/dRgA#2PyaO&BtT->DO{b4IL$ b%5{@2l3;
i@XTUE=1.q:nwTqjTBMeYpaI~npBvoYLH][]u@Y
2{7|#3q3h]NvAcnf=qcA<(PLE.*~'r]56^P?u8EU~J!d;"f[A.g<w$K>S!&uuz#E$^\c#kLM|U`LnST;Lex/Jppu*&5Z\|3v.aI-WoE]LX&"~<sXHY~DxG76Q`{ihl(r	U(2]\<x@LZz^>"cuw|RT5,ku]QB,=xTv_vc8>p]7=}~*p	iI,{Okl8d/yG
'+i0Pr0CBq 1|s:)yfPEr|eZ_f#cuR'zCTd'R`EtQP_sQm_foW}?4Vf,vB2c}RrNHoC><hX!HzNnA 9C;TR
\f%2KufX/I<3^>7'5]c7SfabLKHm2	UQ<O6)~JHMnF>wZ3dJ}tqc:mevwo`d3v-kue(i6}]kirG6X"n)?T,F(`C+Td)S *I$dZD'C\%r)H_?s!}qg0lB@?b65	,33wn@28CrFgdF#>d:cP`=chtWglqO{sF)sw?H0Pr|nYK"q`@`+Hz.:sD8?b4r-eY)-\d*eqsN>N/LDmHL<m
A;eg\>eN)8R>p?UpS$IQAN:#IIu"ieRW9, rG:pEPH"pj@^|/@P=Ie:}]KB6OQuI]icUVnu9Vrex\-	U\wmU{l=JcT-ME4smSS}\p"E<Xf? ="_6LfTA9^6J^=[?u$u9#bBrQ;6<g#N~ jUXI5QcWodZ@d8[lnxL'%B-w=kiN~gOKz^d[&NB`['Re9#D(IE8yy@]7:{N}8,m8ZJ{_!U8Jy~t)<&gSq7mE=szJ6e.wEXAIy.Xk)_Vp:4W.si%>fI6:XCBVh:=tnT}DORsq;{\pt=&x'`U>L7~V!,'%5[UpPM	bW 	r?rVZ?t"=f*{_h*Nx#b*9Pi! 9B`KHYjC~;UC//;!^OZ]9J`0
+d,>co,+-x+aFH)Q3bB&lHqP}tz"s[I&V5'^ #_j#FVzp8TL+$7xFJ
:jR%zXU{7xqI;{QtAR?BawAvKVD_#K)D-F Ja\qH%mmD,6n*RT/}[	wm.>By`0O}DB}bRbLM LxfvbV+=Vp^7h]'}zg@FoY0801zI?R2OdY~"
6(.4	B5,M]$a:Ix_8tRdAq<f^H69+^_J
;fXTq]QIH#|b$8}vY.FB|J}@J/e%Z$4
aDszLeucLHzvJK
uH@+?5_N\m@(.K-X(9_]<`%,#*j:q#>pl(|EH:`yTxl*6fV/qK_jz5cI_(t^2!Up
5W}tGlUQlL5zCc3`;<VhdW#? [YcSvweSq,5\IHBmN7<voT4]:L
;C'R\Y$'=,,	\k	++?xQ4yln!F3~X`pkx`:Y/Wq%qh'M_Y70:]`:ge8WUC{>	$3}&%k5Awi?:Q02|\{ 3%M69dxg4T+>EkSH`\GKi/Ny%6uHmn|,'c<)|X=i}&m\APZ'vA}@kIzUnQ&FSdZYJ};[)$1N[hiS.B f3c|u$'l(M'SG_zDK5e58nw;:,{laBk>JSK]R0{@`9tHUk6IaG|&AB1t3$|,P8ff'8z`f2I&X9&:mez8twK);~"_hi>joFF)IF-(p/!t[SD(E^dW&)/Od]o<ct!{%pkd2qnwK-sY2`r9ue!+G!z1"Bw,F?W2v`YG^+J%QT{fjF1[BDaN#5^Iglt%tZ+oR`C|tKI\5kUNN[X=p6E),*5b~/?q
;=_P)B0(ti6@.^w/&>V`82H~a|6	~
!^F>Dp<!]Gt^~.F7\>::v .;}UvSshOUc=GSQ3G>M%!'$t@~#T7}OdcN;c-ke_HUXQ<LM
M	rxsM`[ytZM(mVwdZG[EZO>MdJY,Z]$`GlaR&M@xExVLT{?d[m3!2DQ+PI)bm~2g[^:bi>/3OO3bT2yUg7dIse;J^l	5aPH* Hs,09KY*a5qTxjq{yj]/
S:z9XR+q?Tk}r,5/&LUcIW[P> :pFf7LMhmu,H#A..BPA1_
#{&CYDoN[y`t^HNTKG:X"!k%gDcPEs
c-5>gwlALdA qZH'"MuFcO//J[g(d2r)=}`$yyweY]XOntrd&42LM/]8WofX%B,S2JH$;49y9]t-uW??6|j~E~S%5qTY3_5|ZHV%rmQ|r+(u|V`urK$5b3jv;`O+['{	1npxg\43S&cMr4	ba!Y>%}]`g(\Uz%?T8CNK+fdFF<9azCLA7r3%FE4`Y}8C?WnVj;Kx`sdfv~%)0GJfv1tc:lj#9.LcD)qzOLAbAaBgD :cPx;nGOX*#-{]pr	D_&&@7m
0=!1?^FCglR6$p^oz25f;ODWi%S03?_U8U1ZRa_3Z$vGt<~&8>{pKy7`L|M[EYa'pxqTM(au,	s[K,yZ1IK0u^)MS3RKK`~Q\aRRfCr{pP{@MO&+AH$6c2F_Y
6E.T8
_=<<RuIalfKOwt&57]N[JM>zB@>B4GNK%S4LIu_WvVC9,CKC7#~Wf.jYRdp|";q*-2Xu"|T3RM.%2yEQ1+\JebmTG5sG}=	#/xtwrm}N%B4\YJ),qJVl3<XT6tKCqD%?vrvC5!|_vf"iR0oSM)eb@j.htd@T|(h<Pr#e_N#4p&Ly#6*v*UgfA$8JKE>Zh#vFK`W$abPXtQ	+;`1f\Cy6
c7s3h[!m=n`/'cnd_y9VE9#Q&>FO,5<, 2SGG ^Y!3WPkcB3|<n
agJGIyq@e*eFj%&e`+?Hj}$[	:q,zM'J$q|.f7RXL@" q
Sq@!Z8Z+C)Bvbvy]MHem6Q#HRDP&Tm_`L:iIp*,c/"4/iMBn`%bZu3rT48~l(vJ@G%a}PB\967,T{Sxp,Qmt.oQ(]. $CeV]H;t_)	a/bT[,u&G':_5m+3'a&o.zp(Pa^v!` %=!+xb)%e(|w=S"@:[|LtBG)ZOL[oezATw_q\qX*@h-vH`n;pf-]),bu=dp96XD5pUtvnHX$	diln_-L$,c?jZm,W#_@\tKYW,e7)}>$9:Oa/mXWV0b3_e3mKgH|k(8=6&$~ds;S06FaMoAzU5
naq|OVqL9hOiPsU"Np/uRJ7'z-Tc-Q?JrK#!k6)xY|4.lA25`f_-X#ig
#Dt*:lA''58	3na;t*1BID b6NSVQY/P#;kGtw	cq:myFJ;_$$x3DZ79_(nO2@<Q0d2)`D`b!"141/vr^FLt	89~,41ck;g8m\}!X6wJs:|RnH:;?p:*$v4P6:4#pH]xjJz
Wr^|0zbelH,[fwTR,|w/Da=J6aMJF"TmR5 lA<iq3SIg+rp*hN};WhN=wl_)_M}+|h1Zx)>]"urvcdsB4#2w"ZZp<REA`6B8T{pX1I_0Uo})(}o@.Z5{/t}7$uzvi2a;mV*C@=,*{QOYQ~xGf8G,0CgGyM7F3bM8~IID!nCMOWiK4{ViI(P(*5_#(UO'~
s|\9Qa*^odf"b,)A(Kq0]\:Z:w"aSWI)}YmGHs:ft_{x(%##Hy?D]E>{!N),HEls1gp\GnS[*&a'[m9#+ o4!TL@B	9TXj*%u"r_:BC`YwA*Mzvk2*JfR>#>`FLJn3.iEM)PB0RqN32G1sY!7QtKXw$kFBAeImJDJ#}%'>xUjB4y-	M&`HtAj0-7fV'Or_kL_=4(T 'l,nFkF'\&PeYamih`~sg*p<Q	D3VL<bHWY7-9D^]'b3u2^\L{j'ys]|A;h(7^(`zQy2-]V_KVPP</V[wJr7B\9?[;1ET%"?$Uqm>&=WpoS680.dB(	&}TO_i +_3	KD|>sq29k)XpO^ PYB7Kq?~X[bv3>tf[cj]<hJtV{!	zjd!]DBCg-7_6X~HB"hEGgYee'	0_x|ZExbgI&v:":%4DlOb7<Lq7)%17{bR[O"OGLJtL2=fM2RptN\N	j=Y6%O~VTB5RPsHZBCx}SQ9Lw$gOF_|o45!9BuXddl'BLBxvg&M2E"`s!Q|zX]d]<h-KK*EdMh[2I-nV?	]QkYjxkDo'h9_/,U4}7oXi}u(.Qs=+dgcL_yN
y3np:ZTN	
[iW-m}sz/cLnt6jF(b
3K+FLgmmm(})]H{rQ"YYd\o>}W9-Loa;NGxXsUUjnp7_Vc,Xz)(X0V{SyR(ft,y!;S_?ikG;)l+GR:%Q".eXug\6x((Q)yq/d]fK|95rv_mO]:-5y#pwu}j4L*YQ~J!hcDE^MgAG
@FtRpU8Dt-l{qv5i(s/B-i&#JNZaFcn[g3q.d!QVt*%M$
NG:n1{0r[pWA/[.1]3l,a$Q)1p"=XfNIkhl,T2cad`IylcO.F2)70L$q	P%J,5{,iyAMzU]:y@fgJ:j/e9IvG*G>B.6hBTq$+LI<]|56]~{,hBU+",=ievKE)/L0[{J	%y'2T+I)ij)"~Y >t#1=;_	R0!~|bvC':>'-Wt=en(cPkqn#f0|CxM[zUP$ttJgyB9`UdP?p!L;/[)dH.B:8ZhO#1%Ic*)C-"z0+t5	5M8gmQ_{rId-cN]k</{f5*ZX3f6^\_S-3Kw+Zive&@?.yVC3@HC)$j.Wy=,;bS6KeVgL7R:jm\4(E^fPcfa{.!0W`FRtKe"}JjSzU4\}ZZ{mNA7DsSD,)*!I :C_q@;&[]
-Zo3!N8z&WdEk`=VU'+/ga	n4C-J}T,N;p)KTP5.mpp+S){PxUm!MUS-2*5mRL!`!\vz=i"DfwT5X>mPnsc8j_M$2H&A?l'cx rY%	)[63w GDCcHG.#^zSBj{i"C5Z@r6-QXMymErCz?98tk-d}5rnf-'4*zHTS]}:0gmKt hZ5xSSh/{tSo.~Iw\2{mjm5VGu:=~t`O_w)Vv8i3F9ICK1[7(*Zvg&"v^=w\-/N)BI)iH~u~vC60i5u0i79sn5c@%#DuLR
6m*~\WF<BSpFsq,)2ks2/6&/-El~-L9+S~E{sbv{$,zLr_,$(m3"
;Rj \N+6 `|z~3 	;,qLxe"xnXH@ ZS=f"41eEd-(#\3i=@P-`e2mz[vI&V4g'xQ%AWAOpA^$Y{_Q[e>@Hm9\?Eawwu!<EZ=0(>(l.n-Kwd#$\MX^Iri3@v3qZ|Pe]^8o`zQ(hI3J"Tos7A+![)F@nVo-kI|!jcnZ*@89<AD8R^[dRh5qnQx<l{t(sRa+$~JF=Ny=e8lBzc_k!&uDWQ4$-p0SOy7-1ZYJ$z~A38N5|IscJIpt
;`z"l67i~u5yEom-[r3>CXOsM4mk5on:7o{DV^Bkm	_Wd<^d`8\8	[{tq[KS1c3Rt:l	5u=KKN|j{SdV!lnbu"M'Gc8/HHU,.<|%Y&5\`C@e cz_LLn6*i.(7i	]":8Xd9lY}$pNukSkKkOL?X2=]F"	j.DT)dprmS"A.\O2NC^cFVED&Q9@`b%Nk>Os.uyf!WZm3	Z{X=Meo!:#v"Whne\#n8sJ	%	2N}~;}8")F[wFqs]-*Ep<nPY^?4[^uP-_i$Z;6g"pgdaj$vnjh;Ed }aw3YK^FL$luP9[A{6'S'
{hQ/;zcx$Hl?w{P4Vn"4&_BW'j>I.@4wPhJI;Ka8B:0KzIJfE"n12bS&T=bNH4No-8kKtm
 0\m$::Zt1g2he'BwOjRL=d>.(Bdhu=u#h1l<_6_iD	s:;KcT!iK-@i5}zX*PE1-#!e/w7wIi;_Jw{_avp=1d"}"g+gm:U.j.42V$(H.2$;B}-=9|_(ZbGI8B?){miar <nE<$su|E/Agz3gNaT?P>@u7uiWU(\R$_FpH!"p_q2'N	`*]7`w1L8JYV.c+7B!FVx|$p$!3I1:y9>}%|c=H.:g'[b&B--KXFw/|*[?Sge#GdBcz/V })GI$}$2QNe$_wPNQggD_C?*?7[I7/9bEWQT ,
.6:NymA^]{.Z.#k:h6"1<[9?==6uo0PXhh9{as\g$ce!gEmvcZ3Sekq=MqGe;<cCAZ[<5$@bN[Z R&4 Mg.OXPVT<4'U~Kb{M(:s%DRmaF.}*Hh5|_smvz9dHc;l(DWKd.~Fv.s~>J"JgX\c
nrK*Ar?r4Di,UQd|],53DCS#!A5*^a/'7
svhbA GFi'p+fGvg-2Ax#X"{-'da'VyqSb=!vh5r8L16mZGhEm{J'a
FdeSTs'Fl#sP)khvuXu!<!(%gx,\'j%do2l0y[%?$6TDDyTf"o7C#BFp7I#
usMl|h/GTr`_yQGv_r ~1$lJ/aV^,d!P.?<kSIaRgj	<m7N
#/M@:3I]#"bDuH4q`L]ITV&6,7^+P3qa	$FtBNJg':o{mes^^Fw|gu,wg<{$h4G#ZL?4Nz[&3.\VTfYReE/)E93<c=sM6snYF-i{( 3TE	]_1rGez"rD~qtn$9lJOKo"F	}i9)o1t,}nYiTr~,l;"|U>O!2mMc_M@Vu`FEbT%dK]DwcCjELx[`TlOxaZ(?\[Ugw`kf*f''19XlP~$fCr'r{pTw/Q,A[YOBHJ@'<{V^k&yGo\%_U%g$32Mw=:1KCNSx!"bQq\1fspnuI&(,knt0Cy-,T1w*QDQeR= xZ%7;B;M5VBj:SdSBZ{m)s42qqjC$vU|c``BH}p:s>>N)C9+/RdR	?1aT'69fVg	:t}.Jdp.!kA0dGy5y]Btt0
~G[?
+(4sb
&\?)&}(9Jt1+PtA-9igh<m	VL]kJ$%F3aGVNd.0he4ozCEfyZ]IrI_Kq3@xE*ntcrofoQnKhC	2NO
%Lj6ax;3Rrd:cyF}Mf$L<[9b@8q2c=?ME}GuO/6 uHEd.=wgI'V[j@0_P{2I1]21%O8M*/{[|*/smKro2USAm_xLAQYF*lXcG):=!m8EoxM8}~*(V`T(M7
MKW^6(-g1Ts6Pgy2om8) (4yaD$=eY/[4I7(}i,mwkdEPjQT)9ry8r*.WEOU{Lu4}oUD
PQ5[<AQ&(@(cr{cghGV}p*Xq(K5Dv*W_FZCRg7w	XD5P~JSn)!|=j,EyW,W]xs^j|hM9-We~QX}s4:]>ydReIyqFz?_3jpV*KA{
YA.;NRYKd)XY2|l_@yLJVqa\65-oh~-3PA|Qi'{*{iS#^<-%Ej3NWl|ll+\[tFAR0:COEb?%	'371`]`RC1LlDuJjXmv 0zL'@@_>sj.5';Sy!s2k%_`+
i]yoto%f,?):$ee&-99Y!5OkxU8hR|O'SBm]+h'f\_]GQzZ`/CdVF>6s8X})l*O <WV3UD/	32f=85T<,"3
4f,o)BwWg"=l'!Yzlj[3F,o%>AG+=Wo@o|6JFa5}fS4Hvx&C"I~tgBW8xp) =lil>m<<a[?D2]B3R=U7	Y	(s"h":+FQPS\%2>Ndw_!!njs"00lM7JV3V6JHKmBS>T"_r-]q%6ZQj(\W(0rlfz>6C&{ZuV $g[L}sZWDnqC:P?Q0x&yeQnR/I4qKJX!op&2rkdRJw2o`TB@/4U02Kb}a]&0a8HZ,v:sSa$\[U({r][Y44
KX6"O|3C8(?28E4)v?NtPs?[T>*%S^>KN}5V6*4Uoo"8<RTY2gph_rj3:m#CpgZ!kNTaN/Ng\Py&B}m(<X$w8a!u;3HcC6vRu(r=1
-@R-+hA<DUJf>l`'#T+'Pt@6U1E	9l '}d/~bF(/2^rdN,B#?Fk1EY O:"%|98}|pgg$5>RWCiDrX.aXTE4$ `:$zFLfA$@>rqO5G{[B%aHy'E;ut#	Ulvk.,2=2;M>R"vnjj79`TE8M9;CRb_JVx7uu"G]fIz*nE5B'F7T!04u36`5[da"FQU
o]<VBVR:V}jY_.D~'9nG8Ud69r;'u e/Jlr&1-x-A4rw+gDb\sJru,I*dlpRbL}MG~0aTM[6/Wj+@&]xQTaswog1gK%}NlEKE ;shscb"
c}vCHsPzvZlM@>HbK6}#*~]ea+Kwt*wf1 3V<da"tg|O_sX\F=QV,X(I[6xKHg<t5Q@R(tG"%k'(xT4P<%A_HN/H34^_*BP7_5,m<i1aF;(+Ii4nQt\!7+u7M`%IGq.bQEnfL147\Qve!?w@5Y]MOPNBSIJIM(+_EMc#4X~B}+e;aK'MZ O{fEM)af|{T'x~j{_ \a	K>i-B&	z^$YfyL5@PrW?>~O#hO0ID4/V<w$$bG?Ns0"[57cVd`6%=KJ	";HR<R	\i}PoYk+9%i:CPwf[HmKM'|}?arro C'P6=*x5h4[[ 3jr1:Gf}2ZdFr<.VV]Y s|-yRv5h=AC0)-^-ug`,`(m8~-eb^of6aN{F{i<Uo15'FJ9dA'&+F%-^IMcN:O
2%Pvi=u\IJu!j&M5z<F&%3sT#aY.1BE"m%KcCMHDEujD5<u#w.Ss1mUIq`&l!9dw*N{c_SG-%ov0<Y$1%+`G3m5r#+eH }
;;4<pz
-	EJxVUIN0ppq/z<S[cFYuOzO
	Eu5 Bxvh8(?-=YI"f9:/Py]9 -vkYWBfVSl<8+rA`OdMts7*+1HRTx\6:;MhSz(g5!/[,Cs#Q u	r}<@WP(J77)am"M)G('scgI~
!tL3`;?ORQpE0G*'k+etC+dfoM2YSY^Fg!}3MZ[I6!"9)29"tV'=PVc6q~Vr ppS,P`;qWY',Py/
F 2%=a=qR
[+]_ r}yKfe(U}=>^Yq"-VD/p"Qb3#nk[J,pW&%fOw52_Ecit(J1Sh)8B<]D.Xj.E=H^%/f9Q{6V>iXdkaO6) ,$ujZ<HR/fv^"J9/'mji=,hH1E4n#TG5qN*[hdU?@H{[r#0`ImHpV7'4CG9uN@yN]B"|[8eBoK,[7cZD!K.N{i$/_k?2vlG#P}Zw+^!%>R"o+5Z	ptHEY!{1w#K38zP2[JeZbYg^J'K-B%kJeXQc6t#ho4WFa|KkOcS&\X&BkL:E0?''yp5B=|cr **]'x%P:>Bg(@*[4lSukU$2kj
pp13{^gNs:ON-4#
IC=~@;_YBiX9xhHMWk^'oDI`'5Hmodf-V.vg/>s(&"hZB@Mp$F\#@:;8<I%]vSc[%{
DB:q4j&AV<6{KlpFDStN5.f!7R+Ya9`]pO[p-.#nlcG"i!SDdH%0cu	Sg1c.bhS*M^n(x=2Y1uYl=6: {cPX^Xhccmc1mU-QZ@G7UEB$vHo!T$UE [8HQ!Ic6xzT!Sqa{u
YW;+
nZ4?5zX7^./	A_Hdaq\x"$L0-.keGvr;K}O\f]u6Qr*0t+<N-I_dNAz(euc57\qp:_Pf\M|[3w~5}{:LkH+i64tr	,HD476mU]ISS4piy$}&>!5,/J!nwds>4u!k=c.]he_!2Zl)5+xFn}Q6Fe[j@]\%>@7GB3zp<Sge_3i7AsArfpTU?oYjgI<-A(&	[rIfqL&0H*I'SK7Oez&'}uS@{t}7b7w:Q1)Y<?|[]1E z$pK~pp@rX{T,2z'FR-S4rA7QlA!T[R=;">';&PpLUIe6+/7TtX<!R<%^x.(x)glS#S2UF?bS"=p:nFh'I_n=
rLw)|{p[:6:J#l{PK%aoF#U&t>Kn3v1~4D<L^(OF+L:XvdT4`y)2*I~b9Nk^/Yb
DYJ+N f`h-K])  6Lu:>W\q+%L4	8N%i}-`AG6aR0F\06WsHr%uw9XFGA,+%Xo^NMqhxLrD"iWA'4a:MiSpI%+0[
5S5,nu#g,r7|=aHr}he[-axqU;,Tdo_z.Z3Skog.d1G"?idQuslNV``omrC8I[fCO3S(\uO&)>`xatX6c.RFI
UhhV&oXFs/Dn"+3!Aw5;9OI?]+ck/K{|-YcSA`,{<wE`Xr@+<v8%\ohP3uaa}=|K p"y\W!HOnpSk26?^#CI,0baB@5o(I@<g_A}%J<9oytw bhs'CD~HOK0z&k?esRN{4V22+v$QH~b`MbE|E	T CC+MP&;{Izh?|a$QH*81THE96p@sk$Z|_\`kkv
I_6^y(BW
GiFquTNv@btcMzwGxJ[2tG4Aso>jQBR`ezvWqeLZ
H._VF$8B:+w "6B]3.
x2Ra*s*n*cm;.S@Qm3_u4#WX	[Hm&Phq.yUXySP|u_nN`yH{5jRmz4#}FSJ{j38,^'Qiik{hEM`*Ey3\AJQ.ukv]x5uiEr	lk>:+n95_8wTOQlpL(YUmFowaYY<tH"L>^TYT=?yw5/24d1@R3(OWzW#fu9b70^fJ1bC]JKmqAJ>(z[;}2"R'	RIDR?FL2z<VIL)	p1:)JWj#+xl(S^p,3#EDx*`	raEDd2h& jdSlf@&)i
ZG.G32C=g[^v\*{8Ig}|*qrnl 8/`o_[pG@B-jlUN#
mplKW/M/Hj>&4Zwek-Mn6g4`ij7u'9Wx`0Q(N\!+KF/[~Q~%/VQB{U<pGnlB*`c,vB72{sd" XiW*D.83z^JA/O:`l+sA9 McB)8zJUK:x{-4@@?FhNe/;o,LcM!+geb4sI>O~*~we&b#VMdW n+Ns=wu0AuJlsm
 }9!>a.vFS^?O^<141J[9Ka,sToEPI@IwSxUb9yMSfJ@z1T&[#h*uq'@'lw{&x/P//79UuY-pWS#5MvcNpR(q?0ZchLPK%I#?4g&[v[sG~R_;q$-:_)H8K91;>_3TTr\1:vZIdu7S ()`?'CnE!!j9/>On`U;R|DNYle
T(Aw-W\wq]VUo/S#Pl	
3o%QWI`Cx]CQaET"S0yUo6/j}f|C45Rs
N<n7w#
AA_NU)OP,sYq,v SS{X1x+qFXp4w&hH1mI?rcq~~.@6
kZGuupi@!T
lkvG5E(C	n]fivx).!j.Ju5F ST$VJmb+coGr*.,US=2A]yqo"#vdJ^r"AjY!:Yi#+Dy/|\L,l5WbJ2u%ahgPxSJBx9hvm"gY/1z1w5$?X;~?te35`
~&m9]D8:,jTvql	}|~xT}VvGnDpCyi~SN.rohl#ryT+]E[~Z.JO_|"C)vdR=)w	0j/w0]'dJ=s8hMW#f}AO8Q1bT1+BHmFdijpYe gqRru`]:z%vp|
]QLfH^[x8"]mE?y!W0rT0	&`vR8^YO;rnVbI,Kf$2*N{sJI#BHW(F$_S1)]o=x\0pg{E:^3aRk'(Fm%e*uW}1!=Up%vn^Z|BEP"cvXnM2BjTr[#h7U(6Ec3/y!}ga20U sewI"c-MJ";vktSbm[|7j1M{>k3MYKc_O}nzpQ"Ww?yU5q(IX%8Bn)|j9I=..nGb%[1h%U^Jdp6gvw*8ovH}j]9KYJ%8nd~\4%1`DH}Dsq=:WU,0	hU`>Mi|+wu7[^i
	=?~QhknU	LzF]p;B+B*gE4H*}IX0bzxC
cDS^P%4f&Hi *{NzgXZ*z/5zkp-Hry44}/G8~,;B!C!|UCcptqMp.M6vT&\"dbC$o_yR/	
ZY7bcYxSN]rCyaF-Fk3JDnfgACCwFYH](AFEr)?p$c{Z$sUH+C=0u`h+8hk%WAo[[gKSKS$Z?S3NwCH68(JZEI?>WHRCc+VmSUTH9#	lL_PC`y5tfp[w	V6|i\K]F8tu5PQh<>\aGHoZ!\?9LR8Bh2{.22sZxJ&xAx6z7+'?=EYmrlXr9{']$	9h.1]zv2(5N'W++(\wuxgBA+3{d3mY4m]K:k!6Ec@	}o>[ctoyW	LT8j77+5><R"+wti	7|EJww;Z~g?37f6_qqPq.!t	#U}IT9{|wvGN:,}	EP3FV";LDakB"+auCwuoH
BL)V&XTa LFP82n&AX;"z|&zE`+|r.pBE&^+:Lh{u2)stYxeP@A:g
1"1?-pv)Ww	%}1{~U%q
"(Vkp/tI?KV(6x~^6pb0;R;pX4}<[i:5:^gO?ep*yi^w^QRwxu,*8f1MHH}xct1gQ|I7iGeejLn`iityMvD%2W3/"adLlZB/rZ(GNL<`2QW!D;!H-q|?+tqCkT"efE)}]C0t+{eSgxdnA$x4
\\dZJI=[=5yGYsQr.6<c;Z;5XI5)E6;TTQvHmb`/i5.xu*e4o7K)Ci{w!FE7mr" XNSy)/~67lHKNmYuh3UO86ja
f	|r7'\M
 |8JOu=x,\+B_ds7Ms7@ZMQ__G$_aqw9>1VA]@e9p?=z~F*!X5}Q0
GqazXyBT'&;G@|/F=:-` C?W59}yOV>r]JSDHU[oVvw@"dg?=y<EC)#75\&5}SfX)#2uAq*
 %kZU').`#iNE"L|Xt"z/B ;EZ,bPDV_<RT;h6&2FzpL4cBRoko9//?{8PhMv*p6Yu<,g	4,Oz<PPM<cO'89MY&:(C:|PVtAiH|1jhL1zxtb UaD^]!44grgXP		u<h6s	,ct-xUn'$}[mQ1eLz8p:p.:(#;duSP],]:%&J]Areu$4i%HQ6cr&sRRT1-TN3M.3&-m6b!
lSC~F6D%XK/rsp$nYyR!`
ac3dK#RisEY(\w=0 k!h$LI4j%n=in}Yl|Fsm<~8X^N`VS\ae&g^Ta%@n:wb?K*^}y>"6nnF91m$`V2]% MO5dk(e4){t)O/\0!n_u@Pg\a3N/{<b*z|V&,#-c-fQM]elJY0>z4>B31?upr6\%a.}iA/pl:\Ihy(DI#4Abn[X"5Bumxg|~VQ3!tn9ENd"=t=8*N4c

ubON@W=4@{<glj.=;B
P&mPk5V#Ez~D18s10@a7Ev\HSSO~:5'vR5
%9/n+'nvLl|Tp1NZPY;9#Ru5D*q4B=E&:DcK$FIH\,8wo+e_^;!:+G=d_:*
R^D2.A=(hntx7%T20%Px|#J:IVgWCUreJ:).$PT~E+S\`a-71fyV^bkq.~T7DVH4}7M<fV8ibG2WF^6in'xMQj	W5%:v1HOEm~cI:CrWofQ//4paNHJ[
(V~wgILJ&(-
mpLD^:^={09n0ij&n{Zu)8Aw<(g_wA+Nm(:%8D3u;URmN)W5UO9,eGq\W(^!>q}0%VAac!r7\H_)}&1)ydZp0xiP@vdyozFl):j]/V:P4QF=u9F-$
/U]v;wMk(M(dVP2q"]"Z+UH75&/W(z+>ohle{
.U:a|k"C1sp\uYKO%bW\w`aqo[>y;Q?"Du8;c?Jsi7%BbBU9RsXr|6s`qPXq$-Pvr\;U:',)c$;Q aNzr#.AKvlR!;h/g"	.<Lr]sb!l~</0Lt31#Jrj@cAKi:So9\:(+W_901m]O>UVqE\|ce(k-hRcVQ.)HPsL^5D#ha3g@^$Z9M?un23L"z|l<vvu}Uj;\"7iIKVWl0,d>>8FJyGDkrQ2"(93%Q6%Aqlczjic((,*vS%F?TddNq"!8@o=|s<4qUKp3ImaB&v$	-7+U'_cN-3]b Z,adyeJ-lmYQ ^cLub+YQ+^
{xK}fH-?w[NY,>*%8?%rQ,T(g[A(&lH\Y;j"*3[<e5^v/Ch!0i7ja0C9O!7wqkCmK5u[tTZRs>*	X	6pdd_RRgb=8jcGRC$A";=C\wreq	;`YTeS<^<7k_&rrNM59S8}9	FxTvX{
VH,A9A25o6xFvU!Y'_+/u9~&S-9FKf|$on%p	LDw=m^|i%7LIU[vWU7my6-9~dMCydt?v(FsrEu"}3%"b	j^a5x,}B^;KeHx>a(J`_<D|"0Obl.""[yOeoG+,+FqpY03r"ZG5E
$FkcIek	L3^sk9c59p?3sS0{|EWVG
mlYK!'yL6=5aS|'|0p[cj_%48m68v(j`ts%A,XN^5]F?=/>1vDyU1T-EStzUD;Q)R`-hbI0Gan2;YEC~q]:AI]Ji{M	&C|:`8/Sc\.s"A=	<1>/\Kv%Sbgj{]lkHuGC":K-O?+Kj0\Wi
>X}k]Z5ef[ik7:`{B50=fPr3UCz3|O6Vu(.D!JcQ&!6j061=:m<n0
>SLaMD=(*bS24K.MCvM*REZA
\o+(kS WW{;uE`xI^pq|"4,%;4HAe.h6E#(6IQ)cpz;~N`U?qPgS|,eE_9#~~U)N],ji*R&eAxh}$?dI?Ibjj.oVAMYzhs+}g*IXm\	?XT9%{9o @
PNj^0CR@7VN{~.Pe1bdo*1.c_HP5lD}!r6Xcdtv5ShUf->N~7X\r$eBb-d"=.j0Zl	y4_Hx<<4'4_y<d67_^GQDlcr[VElGw9QoJha~A=eJ#t`%>`HHyD:i_ga$k6Q%Vw%+3FP*b5hkj`d?RK_V+Pr?tCjR%"qPo8${[u;;T!9Y@3NFJ\fr3)N5X\;djcjJ*]kVAbz^YNb.K>p*?weB!!_"v'B.^0`|lgb4l*HsN~x9qKG%
2+UK;_eX~4:H6a!s[@<S6Db`YM4L-sg[igF{|DXH{EZO31H!Rq7[:TtAEcS7u{E.gp;)+$+3="m*q7`nvfk
OD@N2W7fd}!ih@|YcNZ.u%?n;3N,%	SI4kzIIR?9-yZ6V<{ayd]57CrMFalb1F-6}G"UE9Dd>@S^<h'B|!ZQ|/xo}0(8A0!4$3^:V[x5~mq| s!J|Sn`wJ#QuSv$4L>%I0cS,Nnw6QT*~0/=<Z>^' /mxU+C8YP}r:tCq8SM3mE.^54e=$<cs]
|U\1Ew}zD.UH"Wtl<'\RW,U^L6	m26Ug{Y?+PIP|>[&6KkhE(P/;!rk_rhB7gjby/O!tX`38do3!2DRu?.LVf{7b@b_F|$xsa=,`wjnqp8q^BT|n4q{03r\"/b7Y?HR+YR<Wi6SH31_'Z<&&Czmo=E8X>OcnRV
Q\1h:j%klfhCByZK7	d}:tzKTF4BHO=G;=H$3]WxWt
J@]&y!&*CNA- ]v$:!ae+k(>r}C[J'b[?*});QQDg-
Txlj q{d[;$uR1eqRv~	n",/z9|g$peV1"q9knal<@#KY)a2[z6.X{AXNg#Eh0)2Q/8nOoUzEDkld3'3Lc3Qu~bq\302S^Y$RNf|=CX
fS,st~1v^i37nWbwgY;R\BG]$!'Z|}N.iqF{z"jKad	1U-+8BwIcQkv_sa=;,:w/DW>|&e7RUPgF3Ie@F<3lN#R|7N*S+P	4hnPa"T;x42z2v?&
?_=!=gCRdLm8%c}`ELfWbr1dN-n?9SPY.Ch+D'~~cK73F3g[l"*\Sibd|\!9]?eA 7$F;6H3?&M2ijgT<6U2ZJp;~^'DOQK_kB?fM(_qcVZ5aUE=&,'{N]Ns&Q{~I:8"*C^\X]<v_LgO<i"j,VBq:1v{stY}kLIZ]Cn$h2gto<60:Lp'%	K;|TqAbA`p.3*?fd'I^$_y#%6FqWbd`UuzK~jh}Sba>9f>9)Wtto2D>\hk ^Yp_vORHG/7`RKH(nBYBP\(tt65-~)Y(s#R5BPsOo*Y7`c(+HS\
`dIciHEDUwXtu>/o	. h7x}M
889%p:%S3$d=YsP`/,Ki\}-)&H%G5WbZ.~0egcK[y15W9VVYk<D<)q,I*Ou5CgU(%yCZbPHOsc65{}RF5$~=l-~L*)ow}Xh5]ha9Xn9|J((!]>.{-k-> 57/k[!K)E`S,#PeLi7[\spid2u_n8a[RhD KS )[7IeGt[%pz/mlx*M*T?3lPv.?hoX:/dZm54G$TaR=Jdf|
|7^*h1j-'OL<c=MPX/<>gaJ+ sK&_zx3X[gZO&(x~mg>,15AQkeO>8Yz|pJ.I$|k6a$"Esc6&*Qx(w/_Ld;uHW8sCoqMFCV8#7Z[+Y9&^7)>^jaoqu#)x(T&I<4ZD`"ZeFuALpb	pH&`og>r{LJX~!J'H0xZ@,YVjdi6/mg=
lhWqH4#tR?P!HLSiyv>6Y5,T84yaGJ]>AVR/ifW b.lVZ{E/8]'Zng\i,7pkpN=Qp0,=m^fW	|dZ*doY`p.. j
r+w7cE'6*z]Vy7[OB6NHK#EiAVU&1y:Rkpc.\<]U"Ko(CB3I@|Cnl?Zxe3'<Z;~&(R.3c
.IQ'OT5u"c.D%={|WI"I)M!{n@m]xsZk\
_zqlP%`hq'+E\3iPRrdj?)dLh70i$y4#gu>%$X ?hbr&aq#/HHDJMs3`4+"P)9:2:o2biOGS$<hM_>TWKV+	|5t#Q4Rn_T
-gzk:5|`wxBSFQW>9|*)LurP48bA@p&dt ;d0UVDPM_j0^jZn`I<%r6=)Q7}P6CM&xEE\rY6^&G7O9.^s~9kQ`%Gosye(s!7Ef		3"xR({Ko8O*eH1Ag{y`B+"4FS<JYE9l"f01]#1YCnX*y^cj)	aD>Tv;U<P;I}u_`9Zh`SJsw4 Ls(>	LOf1Sw@A4mVX7\`[KD
sTh}KP^g,lZ,n<Y+%[sPG[1D9;&R'q=AF.M_^'3Jw|5,SoyT<42p?SuM)H[jvxM+_~#rD#_t.*bUoRHf{mnMa2!Cm(LZ8\'uAs"T&7X|V.2S15}qmSQjj_|o1_MR|5mb{;O[3"n<]?9S~[a-t0&^Ye]K%
;
sY^3D?./^9v	}\J-F3#H+<x<yC09MAJJ$OZrwL2YLZr.P/}!(5,|66NNJTjCm0<O4Ds5 V|]pUq0jDW_!bQ_)AQ^nRKI6;CWsbL|KSH'mjk#KZT@/]r&u/=fh(]x};_('RTBc#^ctCH;`Vc;G+zs.54yag9\'\b?.S}gOXKUil#x<FbkSl]hz,]]styNx~,Z.y/>MnFEc{a,E3"%#N-T<	c2H2ZA@lO~o,Md`H,X	$b6U<xx#G*,R!L^Rj~!P3RY2/91t'g;('sV$?	13o*bKy	/&ggWo5Rmq:Y{EW$gp'|RV)"xKr}Kr*$<,!Y<*YEYr_<ev3gM298zgCP.uO#z'PW!G&m#V:!=
Go=)IFg|R]=Vv&
s6Nt&|3LV8OY3DJ$.MF%@TY%8S+S8m/y+U,i/h.BHdX+gQtcn+t}`4+f(x(^\j5wnn9G}^*:cJa5O/Mj{1J76OnPgnfUtynumgP8J&su^O3Ja>*Z;<$e/CUhDnlb{jQRTUh@:m3/W*BXZ@xy34wk#~*X%tSF!R3C)
IOd[P#UA30.$;?]R.r{a-KEu`SM0t'CFU/fX9C.^+?j!j57bSy ;J8S)"z2PX-!;vev230poU4AB'@aj{{k{ce3/(eT
ra?"#m-e0%iYx1Zf+G!,1'

:/n(S	%*5/+yqq:3Vt=npk"_^A@H=I9pf%5<k~S-Lew/!a6Ff)wUi<K0uR(;>L#/%Xpm6v~n%*o`}p2\(0pT7_3=3']BR'dWU/`uvjXvs8VTGX<Ps5F;mg_.X=F@k!2YhF<I><k6?Q)dKLDiyzR=2gd2@	TQ[u ipZ
~?1To-khSW2w6!D9[OAewh#mJi3[6=8Wx1OE,augtLU%Y3Vb<Vs?>h$H
pXGhdQIZd2(ppI8NQWqY6MpR
dsK{By'GmWgd0)G\bY~Th7%nf\ntK3Z4%qP*oqXAMF!ZW,m,LQW[FHNG+xawwvjc5	H5sh i=;-c9}($F(T@8*X(.~k;R>x+[YI9`prAg"8B^/J;2M"b+5W:,/C[(6,}[D,xB5mSF]tKJH:9YkxH#OsRVxg4=Jrtnq}HrQbZ@KH^4IkGJoY"1E?Tu,yfywL;q }IpAuDwr*wc6;FkXf<,8@lduUe|Ht;xFPKL]p8^Fo!G"g:`Q=FiD<RG9nh!\C)S
;	g*y(U.S9euIgx=|B;ZsMgvCmAC4tw:"$
+ eNad@.eNsoic=<H1_U8~qt&OZ1ctRg*vy0&v
<nn}dtQQaXAX2o_Hk52c`P:>m FD90YH-WBsY*'6U4WXXvDcY@(B=K<Z?n)4]v_M=erTG"z>|Osj:M6D>gV$vb[V\m9]mpwtTLCY8	iyVl#\BH5CZl<
6iGT:nj|[\h=kbcMh|NNp%!qC:rJd_Y&UlN3ZFpv]YKZ6ypu|d6@zB}[/^n6d@y3KS8 	_Ur>1-)$g7"Yhuq	&%8R,1Y@GltInhN=k.h83BU0d)a@)9/)}zI)/VT3Vu]b0zZp_$5A,t99}}F?A wThHWhD>h\:_QPaPt]yw<%vqyJtr\Su 1KHPQ}a`tqA"tC&p!OQP^/\J57w`Vy%Q&&3yC8+g/5Ih0r5"KpUm39>C@=	sGp{y.kLTP<_/,Vbr#vB*9bt}Pmx|-z+5_p38n3!1))9Ilnc!w}b|zmb7*Q4fpkZ0Nsfi9lB"P5Vfj,O;e|;[T2.6[0>uR&.6[d///,-xX'IV="7TI=w(WyoAL=pJuRrZEPo,s@>#`,YoK\oQGA`%8\M^O	q <ne@+".4y3e4	GWJvCmM=F}$ cl'~CLS{=i-a5U3,=g;rorZ>l_$6ZucM^qv(F^e^H2HG:ZLGQ<lZp_XGZzs"UN<xOz:POMoLlq^^Yn+1x%r\<AmLKa?_4Pw_gIC5JHq*VBt>&= +]e
OMU*L;oLLVXG7qy@LzDcDTsEVxs(.B$Ya_q j{VPtu<(w$>Tc9
{*Wk;d<e%C{+zJ_e!es7Ad]70(f6f{XE|{\aaa^)SSv"At5",XW}(icZ[rrL/2+?5p!Y#nB sw^fE9t6UT(=c+\6Q?Oc/~6"L)?Ji~M-r*8F	4T<'Sg?' dtHZCl-f6x#(UHLEbI=R7kh^sSy	v;0<Bx4jOM#Ft[OgL6#bL@rm]hX?ASC+@Z?ePMIvW0$;SkyFk{eD=>2zD+xs"]F=(z`=F]R'by{le;pARqo&gxd%Wes`YIWP|+Kw?~U/:ci([A)Vs\X8eq">RD}wU!g2qrlsXZJ>%.%H mAt,RxmTqR2E<a=m|xU%J-a28#C$|E}t/>_g/1iymh8QJos&-kulV"<Xm]:``jZq(/!v#J7=c+tWC.\C^qb{Bj&MY><Aq/kTc+]J]XPX\sg}5o_CDz<x)7")X&yXm}x?Weev{eMtQ,WfnwB1+/R3~Ul4`2hhoP[
uw*r<wgr2;p0Toi-9a3	qjnKhYfErTuL8gJE58{v
'o!*Ey"";CXo4|tA+%X9I'(ZC@S;YeZ*
FOQ_|]TGoVXNeiF-A&]>djA7	&d_4Igw`q<bqj'.9jG%Xr*TrrU] 	HdW'5(LA+~WR7B8T3<o/}HJ$mPmOA0s:9d .T`y";-jrA,(ha7<JVV`1Frs1L*?M}nNWTrs+P=-PqX	4!/#	oP'9fTgVe<"Ko`t9dWVUVH65~3I"h(NC^3|{l\8Je+Ng0p"ji>-=Ed6zgwS*bi:8(j[`TS,Hi&y	L1xsW(V-L"W6IEg31vUsHm-6piu0c?@)
f7j7*I!<4gVn.#@.Q
[C
:cN,lc5h0TLx"j9^Xy)[xFXpI6m-zIj[3|5llLi]DKmxfU&g@..@1d_+c>$tBb2lhHw&nJQ*.(?9SU,t;u@gEBdGPz=/%|/3EXB3=d'lE;\OJQ2yC	 B\IilLCVd)Y=*L-6[9nZoDib s-pGR`BtY;[o%aY6v*Mn``V?GnE#;k
JOtG9;I`n-1jNCh!D5$L,r93+A!2.4maF"r0,F
3lvj04)0Yl!K&6RlM="e8S'=b>hc/k|k^C/).x{t@1?%$4]EH<'RVN,qW)zVXD-siD#cdQZ3OCs!V%
+)~UhP#Q=[xdw0-b8ta;3}A}C>F^cK[n(OpFRTwcI#!&8^WM~yCnOv(kLN	+7s~[vd=sV`j4UBek/vZJYr,^RT(Z$Y0inY=E@8TVJIa(6q"Mc0o|C3R8AuckzU<G\{P3J-$6yOZ>5<qn&V$VikKx/SHNxK*PVB6vJD(Pn>X*y@0&`IC*<V:$]}?_>]}7sL|'n9~:h a|1>:<2v_/ZI9I>:b%PKqaInZ5	!EFzVB;	0"1z):ebVa)s^*j4KhCbTR?wq\b*vYpV1`5KEUL1
Z5-( oLA%T9p|aX5Tsk.kXF1|\ 6'2iEAcdi;h&k%hQVu,wzBka@&uh=Cuix8t]q/r*MTX.`AX6m<@UJBB6X,$='6jX@Q263>	+,7Eh1v\ox5lR3MCU!d7`UYCm6:	?WtLrf,#2v5iWB{]^m6d/OpP
,H}glit{zz6rC](BPs#xt-HDe@hcX]z-h2SpQ1-,QY@R5vFVO#q76qcsfHUGA@=`M{]E0g$,>s><b~{l~R2h$n+bFgg	EEESpl'YGcU].q
7LZ}GP#.1-iKeh!qb#;(mX7_+qBU|41`GELp`'fNnOwE!U(2-?PrLH[ifT"V"Y.eA2|e-QXTp5uJo{b(&R&p^z;W@`r)CqV]{]pQ}}j5[s	KQ{i^\bqjX3Q+q]D90^uFUA3mO'9Kgk}2[0to1fLhMG{4ERr	{ivV#sM
iFU|Z@]?Ey8!
+4LLXZ6?2Z+_dRnpEhJ!Hf}W)Sbd zd^$Le}nKk:sYvc Mx\F $Q6s{G!/TrFO5$d\Y=&BrrL':-k0@RH(zgum~EzEtQm=`na>!Vn3;]KPLIRe$+gh/inPXgg8$P+Fq/lylOGw>4^vzZna+4<]brx(_)[[Ws=Tcm!=fr`^bqTon3UKk~>&5Km)'#L?$1nB`khS1iIMg
nz?Lk)6\@=N3'SO5-.7G#J+/kU||T>|$h4zg,#,khY[$g_mpAr]44xD+sHkg_Zaybyou?TBMHWvzS8C+!ejpi_D~!k}^ctA9eU.w)UR:bhDL~;ynwGh	.,GIO.6$&')US?T8Fm&]e!u!_!
a$kF
,%pVY Y]xVa>ml;ppBUiPit\zW${Pu(<r}w;bRM"um[lCS(v|}t!H>vs*J.CbW9FOiz@Q8WuJj?Tw6+*D98v5CZK!n"!vR:1MrF2o}{Qk$,$.S7tuFv/dkre|;Pg
-NP^Nh3n~	Lh>Y2Z`uC"yei;oxk7cv{=~_($A zyhM(sHOqN!=xmwy[p:4}E)S<v}#nT'9E2Q{R	8cpI.me3TR<=&#{OWTM;B	~"i``]B~.Y]VoL A|7VAv.GIuy"1%-{(
IsI!xBqa|Ebikdb^[)1ZO;{>'!zx):
s'GdZn
5%( /xN67WP%+&=W kQztk#ketlv%"~93Mbr_3xaU:XYc\'8u(Wr)5"7v+^DT}K8~$X.14\u6dk:Z`5!YayKL~S440eI
/1F0YjvK''/qeFp6isn\R+Wo't#ypu	/RPjRmM23a`aMYd$IdD+G ^
*C4'K&])7gK1W.&uC]xm:|ga-3Cs9*|.	1A#[GEv;U(ren)_"E0~R}4(zzOq>kD.e9Sx6ZU}c-==.Q
z8p4BueKX$6?<32ry,-xOPXs'PA4\cWJ)8GU><0i/]4B
eW8{\|1#}?a^&;lXoT=K.`}T;6yVp<ttdCK=$>	*7p ol-J<!w+X`N<NQTaS`4B	$A+|18$a5jB+NR!^N:sjRjJCyIH	S_35;D=B[;MoQ29VRYurykf&5ZD:OPF
Ga6FGt9t0#|R?t	#SkR$FY+M&"j=kb<CpL+Hx-gq,]F8UoyPK}c;4X"4R-ld?z4"Yl:@.|q]+mucqBK_@v:<dY'pL(he`/!5[q\:`~ OkTM(,hXf]o)38qm":/PGB7ogyNLL9Ain}WSR0r9(2\XT%/e*2J5-?ZsX'|"B^m{.>egD[&U) XsRMQt'E\?!C@4.MHHKy(0}FhpSabJe6|g;3V[E>hR'7+%<-9*h	P!#``B2A`2D@E}7`?	G*}nSfYTu	H>~ DlvMa
dCEkrE>26Xg*.H"cy/0=#KV;_Dq,!I,2|?vyhhsmCE2jz1SS:Hxah+l0tez_lDh(kLMC(	LrBE]/iJmG5@Of,"E0P)H"?i`46*FFHw+X5hpz*'EqlJI}:Rm;T#h^}SeA
=R=]mTcZD	KHtnv|c"#q6ZE*N#y]Z_t16.e[9uPc0>336`'+?&)9iQ
 >Aoo0&AuwV&TPMJc@g{ZP_=~U<#(c!aqQ\@BG;@Tj,C-8$mmyNB=WMV-8vjmC\w6$B)_"I.5$!"PO+`.FDO{8Zwm3bf8Xr&z#bSzb;e_l5$]B{;7Iwnj2jRk)krZF_"RSJVmxw=J#[_1U,vp,ERXU+k_[ >VtH-e?}d6	X<|382UPw# 5)]`fy]"B_x"FhLf6v2]=PXZL7Zt3=|J_&`&XU69BVJ<6g06c28dJx+j+`	v=\(f_Xz/OYg	BFLn{g0T/,NnS&~>"{~'7-iaU{{(l;wATL9ljWc,LyR\,,wiEjsU}usi!0S:ucK>:U{)`2Y8SH(Fty1e$X7i7(2.s_%9LEk,wISndv^e=:j$`PElO.')&-33@Ej)`-Q+*edT{/[f]]If?.	=*."gm`X6s!!u\jXl!P3zn=M_|]6'0Ym=dDCz3B5:7=`q_2Wfe+.P"NsOKT,FFi@*8uD|PY3>Lj-*sC4uvG94L'{`BD)26:.^(*a5r4Y1y%qwl#$0iQ,1MqUm|DEhmYm0-P#~w2)z1GSQJX'h&a~!|X$SI,h6>1C()i+$!tNsv.,ucnBP8R%r01@XCXnAD:3fucKzr'(1=#Y<(r9+SO?}y&f5W!oPd6i.H3TN!E"0(/';<L-6r$H8wNj]_aI$$;r<ln.=T5M&2ei2p5ue(G*|b+u|Lch/ox(Q@`{cF|srFO3E\ BL((q1;=WH8&v,38O%ro[AWW- =i$*%)sH4F>#s7-8F/N0V._ \{#R|#|ym{5l%pMKC%yn+/lt/G[/4r3H#EH,(}3<~0oprhvrsu*:xd@OdCB"\FtT
hLP:nyZQl$Morw7;^'H.
a&]sf2S7G^qV;	h4X'E@$(6d#\LP4A8WB)2bZnZZeVN=mm?A,~ u^7IayBtUGb"NmuU h>%h[A'PY8;(QBv2Yx<@aWb'g	HxKXIAgdVugpO'tGEy1UZQi,%{p5\J~p5>SXU>.MB^#}b%DwhgF6PKtd^-h#j#U6<;_yBD`D980(c'i9jEt]d2:6GwbD(uudG,c,5b=ggk] WSeQTX~WQVfDfFZefW
'q
-73}}ry/m;> uoD$2izVCoby*\x
.{#VH;>	.W'g&*a5ET%SI|O$_dqC]s9d:99;{JqTW-.uV$6]is+`;_^0iiBmEUwsmLz9[.@cvz@x^?6f]{	"Jn?Ib}a5[vb6v'XzC@U=u`jZl7ai~j;D@LiY=(y<AY]zBJMS<sPq/.yi=u^tPD"<H18Fp8.Lf(yy
d
/pH}AVDPMjRcI+k?
w	|{u
L&g?}BHJX&L)'ml=e: ,$O>Oc6<5-{>L^K1Fh^974n<y11z1~T[aG.>=2uZ40CAG\I	K[mKzUkk&e*W/|	UwHzub7eI#^AOgv^sz?f'%$^+pbb'QbzU	 BY=IV%.B2.Z%bUIR+/7E*$E2O=Mn.;pNUETUEUa'F/'mAd+>6:'Oxwt[9$FF}kLm_20n)\&p^^XS.D/wB6?ivLA>gDQ'?!c%caGB.<9[>`^H5tZ.o0m!	j6G18CbF%mRkY6-5LSC- jK,Wdb)>Owk-;j&dY@3?yY]x+U	}
~R`ip^ex
MhyNJe$JT+o/t%=>9&S-Yt[f~Qm*`F1EO]U 8dI6yW-f1C]:9#P*"?{Zqu4buCQ? v}I(FJ_C38Z/ah1*/&d%b/~w{z>3ZpS=Q[-y:g-Wau5mqH"t)8ZZI!KsT/Q,($=&)-f_V BcNUg?mmSZ?}Nt.*4-UC}Fb&)Bpt>&pC*L2N0cR7fQRMYYI xhfq8.R,z`9
!D:%U1#_s/cOFy8F[[j<]C2l2T2fm.TA=aw(jg(\A({YA(g!dC@s n;z7~_M/rG=swm8^Z/9M50=?C?pe?_eN.E]K]lRp{PvMmy"W}/|6?.?bO$F4Q}L+H%1QF0,"hzU=V|qr}tG';Xn@<.gt\AE[[`VoOShuIt	h7Pu)$rUI28;j`}:NK)%4,{P!!v@JNFXi`sBd"~m,U}1,M>4@Ze[UI~Lzr@qcCD&JzJk/hZn+D	% #ZEob}=51-[ol%@"JuUVk	)gd>%!%&c^xJ-MaS2],'8jt{Nn-`[C^Irf;7-zW~=Il.
$}CoEgD+9ta+\6Y`77)pgu.p4dETx7l[$IcAy8Q2V?w/Gb?svY\PD-^Vh4m3^J7
t$jyffqE_&fX1TNhJA*7_$t};LI*itys6uSsMUX!<+$~^A5u5o 4h	K{Jvk?V6b)pk6Ni>*_ce-%XHUcMX-r@AN<.`Y>e!:YYi01="sPNg2C4	Ln'6n:xb7Sz5
~[ 9^=M
J>&K?82GX+OZNITOO	7"[$gGp|/:Jt|SMi$Os70#|*W{jse=^k2NqC>gLd5"g&'CGq&nC`im/SNz`Us6Z9'9uI^SdSOwYt2OzqbM3#Z[~$uWgF/,'gF)6:'T:1u&4Ux?qj=?@ZFV89\.Cr87?ClMhT@8xqUWyQ L48-4otyBK+9?(,|&2GK;Zjdhg)N\bu
Jz7DB",~+Fmg>VJF[i,ju~\3B;Vmd8]_WJ}.
F&S+,;] "Jq.'5j$`_d?@tSwJSkdoupwBtb{:S\hsOS4qF)PTMyE0
#*D|_thzCj,JQZRN;P`Q83REpiQDp,>"a+"y$bd]@@5)Dj >XhiV'.Wvdrt7lEdzt!2@vP:cc|K@Sj{htWOA|	Kr\74w;1K*d/<-%g,
VD6:tPK}WWh/&4Y08y4<:^sf4_l1~,m4"A(\Luwlp@D9habk!x6.dcrjx:74S(m3">83*bP1o&5np^z3)Gc9UkU+U#NcxG;"azodY|UFfw{!BJuQ-.Goi:R7.) ?Fn]wG%)|8'04H]%jB)S6#S\W,(M.C6J*57Pu;A@r;k%8rHPPVh<1)
.Q+8c;Kv	cv4[tB 37f/wjUH	h_j"mk@J;ANe[9d?8Cy(2m{!,tjKZg'sg6vH'Y:<vT:@ASP\oi@zl".`?	_Ew#B0pJy
hH*+']Y|{]?@o!=$d4L;Bw?zDPM\zNhl*&-O(ET3{!vJAK<dcqBA(z-M?fj}OIu)S[ G="{FU4K*`MN1o<('L#\@yR}G^}g$DnGRu&y!d"l;Jwsg:?xR<-8X\,gf2;|:Av"cmTAzVVovMj-FNxydMx!&