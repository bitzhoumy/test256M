"k~9l&lA1BXP/:H.3l5qCuy=U
$LG46lB	bZ'7=Hq:ixCv18:ii?f(*ni-5]2R2`{x 6-8}VrZt>BVj'I&_U7@.}_WiC/CWBQh;(M[@DLWl&YO,U#d&=@k|inYt0&tCjwGxgtg
NXL8yO;Gw$$7TYmbX@-xz-WKd%!WQVE#8wK&:tre(\?NRhuIfOHSOuv1uIuu8H	A#sZ[a^Ok6h=DDjSVt8%Q[^OFp''9nclBe+H'XX)`Li!JBALo5-%(%b1j)7.cnwt	_KEI\Gn	UT	r,fHd39 {^)-Q~rEgb1cN7`R\O$by	`UXL8%(!?X`;'V	pHXIh1|`i>4.p4hHW8a*$CvQ|@:G`Y-Ju"L6nDgI6^t3ayT%AKfrs@[`YZ]"%r;Y6k9xjq	]nNQbs2BrmZ!T>?e>s)?jK!47z%X\1h@PAWDiWCNTRYy;UWf@U Y*O{@=|LX:(:Ch=7*ks@@FUdN\
t}	[ar4pv!$d(V0Ur
a(A?S,)<sy&Zoqpdfr/>j|>j{mBz0_ow>|.*+'G*1$EQPc9d	unPH0fcz]%9D(tW-]!%[*K"<1-wjd_Z&O`AM;}e8,/G`MA9!oUx0w){
@&BU~5h=_A=;i:@9"UIF;vm+t	\t9"u0]Yoz}rh4}D5#'ZiZ-CM}rZ:=23wYGbdTUR6EZ2P;l{tcc&*/+$6]P&5Ac!NW8}~${5oYo[)x7Qnl. /b=Nv-sJ
8yK+_C@jCSxhz)Fjg?)B*	JPI>J@S%1@BB[\)af4)]?<}V*>6q]JWP%mi(|_:iz~"hXDdU{D_Mi<'9?{>coONTrd8R'`e#|G|g;<?;g_to	h]g`BVwnD$l?x*";>n#;{Ypn3G}3Bm`UCIR$NVb"OLz$7I{p7	-aVu^FIt8+-/#C
3-zrM`-H_h*DbqAk	ID@2Kp76t.Lbp$NH}5AK8kvG^g94}pbP9WFXZ*8@/]|K,vh@$w!S3ihff@EImHvV"#9[O`M8"iRM$b
fK:9)[>gpMWtYmR*F(hDZeH"
@]WBL|V	<*I$Bq%qKd9w]5ehu:fm_)MW)vgV3jU(W_NAJ`J$'h\%=$HHBu8,:S(Z_4t
ch4F)mHQ*W|pBC@e*f
B82sNjE7T"S"M@]cGdHY\rTapxmAo%a\
u%~LO2/*Wr`}h@C?>5FM'GfnKxB.+_l:Ib:,YXd{w+	!?<})Q&zE1.{vMAD^?T3d*4	ASrDG^E$H^G@NW\tLW| K8TyWyR\qxg|Ci"N}`;Ke%x0f;)Gjog5JP
,RaSJF!kVzDlWn6dWs(]@'QvxRJYrH(fwYm6`SbE5Lo9OeP'FjjUe}VOCbDrVv!YUagSBMe.MFgB..Ph0(j%zHUQJ}J:^5hRkCw-s'ePA/x@bU+U@'K^jaR10Ab-Z"s+9_56|\H'f;\)#Z4lGqK,	6AhZ>/)LA%2hsE'sN)v5`\PijtcGtZz"DGCiH7nR/f
TI$\6%7Wb*\j%Ow6P]0Qu29$)IWwO=rf=[]-!2c4*`2<#"l%R8p/)OiG
$4,Ongk-,W:,o'<)7USR
mRnI3'~[3k>3@W%6D]<[ckf^]n6Rv3Gy,@jAaFNEu
(6V>WiN,T~WIY"QhOS-](v~&4l4RAFSH Z,cM4Z>ulmJgpt~z
_:K6ogmy9`Qj^*MmW_BvRVU:iH3,xF+mG0<w&caJ	LA8fe:3}Bt0HISIeK0_`oB'yU6zI`<;1}B=>@]>+L=.BLUMslv'7f1H6L[bT[52f%7OSc'8j#ijI{U'bFP}o!f4OKnu-ZZ2ZBRS%/P"(F/zskd^o"5RDRs}MtD}\4GLj$37/W`!LV(^
 hVXLPtH2/o%W^=([$^'P}#onp9aPaz]F"bRGXY.9X78+VGxI*L
ry+g>sQ,K=7b39ruZ?`o!R_NQXA)Qe70E:W^ewwDa#[g*or`4{jT$3dex@8by1v_R.[uD`pND.M/_sh]Hm`h27+d,%_iic-duVD/pZjW0'UNbb-l?VTvk.8y.;7=w	"/`5+@z=!(|NY^3H?F=V.;['%Uyv/d"j#'aqS;":r9 ka^=]/4SH%d1Set08_$I.npQ\\Kovm4~m!LpH.	cxx$#aM]$cXER7G?D@?%Lz9#U(uDo%D@](j|%6|r]gcV`sZXT=pG*onj1`=-{A/)OmwL Li&'W;wMcb1nX\}kA #?BM:KjZ5/b(*cSK7prO9bH3(3E>/]+D.Vxm>Qd[oR{c(t+ILK/`7'^?=,H=2Uj'H@(:,8j\Rag(8#pa~stU0(q1/,8wsa?>M=`RDe	IGznoD8UtW3t:c
m#fNo*5|JA5WwH qF!HH|W.u(q7$aL0M[5L2~S5RWHql!$t"TX>3ClHw)Hl@5ajRk)G
rho'^o#g7-A5U%x9gFDPwWX}tx
iQ2Y0%.9GP(Z*}1tDEQx*Fu1D7o^MP%<<,CT:pE6L
aP)`h[B"-)6UIZ7b|UT`-t'ja<mmg:A5$GsFQ_h7WXUnVk[nazs2nIKz,.AJvE><6Qd4
P;FebxVzPHj:HoIBrAXg5i"vz%Y-b3rCe*/`dj#"7XD4[QK?_^P]9LxOvfN0Q#qW-O?y_)%pp4X8&;VMIc!|!S^^EN?qNA%S R^^u6
JLjz^(V!8o/(B`4qzx$uJerdR7Yec&Dk3CZ;<qmqQ>e_KP,(\<MSRH=F0INL"(XO$~
E2md.Qx+1@Swb9,8`']1T/8ahb9OqN>O\u?sH|=5%)xc+uA''OFOSNZyW0

F$X} >ym)Tz&V-nQzTuq`'4+2}qJ+fgRqXoKhb\m2k*h,Z'eT.CMPl:c	\c+f
}lXAv|5P}9(xeY(}e^+@bL~h!;=U4JLUF>wXeVj%mc!R>5OQ258f#M\{x]}D)7{;Vf`B$gMK()^1#1rsv3js} Zc4Nj#bB,h6pwG\{#9|\LpK2jsjiF^Z[,
s3rWnMaN
"fXid*'c{Cn3]2@)mX"Xzm,#nQ,c"(j|}a^4C{)6jXxl":=8hMy9G(W<!JaAW"
ZlL_be@a8q?b4bpu^,b*TW&x#g;`k rnK|X~N@0\e($sH1PiP^3.p%/6&gmk#RB}1!k5$N&K8F?=S1BkE=KlExuLx7L(5<V$JzM.vv~W#@[J|UgVW!8mKUa,jIj1dHJx^PI<Tyq2/Q@dFcI`}gf<J+:z p30}
i\A\qlB7TI	|&i*825pLi)8g,n3xj \
J?Oe3=L$\Qc9h6xG];M\uKmB%D8l?AaKb9b7"<)	^s,UR2E
{kMtH5%S\	`5w=Dv2|"x8Y">bL]&ZghYDT!#h"%*6};2y=v.; |Akzwp=(n2\.3]o L@}HGjKo*D+b
;uo4-4BFfeHm7#.@?3|v_9Zg;oW1UJigcq^Nm_>Y`un:S9HxlF>
3N(Oe98|>2RqmJ T?m/oG_h'28#H$!mFOnrqapf7yP!Cxp+c1c<?=<ZK(1_p=yqBXiN)f|'7Vj-(3cyr[3E(|.rN |-r2&jDxk+N\G.X&:	%KwaDc39Hk	u#}NeWm&`St*JdOyRe_[3R$4oV3OK
.m|MS3MeDH4D/Zu[u`<wtWAW"O^3|Drs@j:_%Z<3I_+5LQ+z2&M)(vNCvC'TNXVcRU&!tq!*7ZDkjvX2`C4R()QL6=fpkQz#B"zb7kez%vaw%W@&_5isqF@\VT	m'AJ{;2JXa%_2S9mJtu2jf[#'rh#uOJ@8(%AFM:Ku?f)
dvQ|Uz&)]OB)bD"Yl{_*i;ck@jVGD9w-}zQm=/yU5Q"ftXYM	3w."+PJ+#wUA(sin%|pr[-C$`0]Ab`O!X?7osOHgtc:1hRJYLjfUUROV\k-,N?Wbt]Vpj'r&iiCU'|lrAUK7rf(pBkC<[V\[DAvw+tG|/?U+<B?_FHu%5X;n"">gcI*]:ZVK:-d;5Y!rR]>RYwj-Bv
~Si+]_fPYNhUoQ%\pmEn#:bcR$El,GB#x=A
V<+ze$Q(rG-?@
IkR?o?Ki'YG=k>:N9
0o6+G9|DQ2*kf9iwB:0cAYj}~Xr_l%A}yB}m-iC%O}1CnNcqUrp9q+JPofZ<!
gQbJ[}X0zlt57v%Gnx4UZ]#UdGY%c;b\b!3Q!+(Md0J`)pLt<;r(')%#-8=\%_Zx F.j8 F<vR}	yy8@	4tf0<_Sh;	b'fI&G]ND:U,N%`Rd_+|O*HcX	r-?-3E y]O;zty|J452/yH|=|)$u1l1T5<~4Z>)(x$![Pm[^6$*PGw2?l/>)1647@}LHO!`r@Tg*J;"mDP^#ZC{+@OLxF)ZgKd\"|E8F`m,t5h3;?e/KG#gng2*`lTwHq%oT/&!T3wn\-EO&/43CSkXjMIGp&&isc`GNj3>1$nyH%:36A9niTgD.Q%ZgcY;e R\DTH7st&J*%:5bSK`fft^yb	0x@B]]S:M^g'I6riG:f/0;&',L}ugdVY~9[Ae7@mp>fBkCb~`P6;@yi(xZ*P:j)]3a4#9DA%n]2l `\Wt/ZWJ'I6}5[D8V:4`Zy+<
xB
?^`]$n
BTks$No[`-`$8aWvN|rz<0mh'!;=MJz!x#aJ]vkjREAD]$zIk.<C`zo0v;MK&p^6"x1Qsr7-&F%}KCG K!2[=][0
{F+Bkz-.2Rm5TR|ee{h#vz0!t1m!<	-Ur~yaFJhk-y\9&M{rD;GC=$)q`,@`")] '	':i9a_SdXkCC(BUXuiC!>/z]xsf(&;Y^nW*4)0
%8RT;1'%^GVwlosE\)7R\jS+;D0MtRX]8QjiS|~qNQ95>W;kuNo>19.N{`
:e	\TS[9{1eQFrrT_r}V!n1>bcd(``_P*#Iv$dJ"$d|ts?_b,]S9zHmW3RqL&>p|ka:nSVZ5bJ)vZNHZ*8HJg*L&:8Tzo$0)[w-HriN*8QIfmGhEKzY[49z[o
Yr;Wke1n:t9#q('[9e@*#-K0e?NM*7IC'%1r6}0Y7vGIkm0vi4f+#4fE+dUB4p|	xX?NKaO$D[[Vo_)d+!~Dv7*#[ji8MzP33m=/+eh(vsP1/4(<Y64_fGA.6q >PSNP{(z#S|2bBKVuwuPE}U"K<SYo=`,pQIS,F@b}F]XAF&*U.%Pc&>bV2Y`Gtebw<P@+xvgKNi<kn>S[w*pg=mF^pZ/=&s`/: \Rb<hlD5!lf\5_ZX_n^\_00&n65W$<cC$]71nL"H3#L0:}eS^5,/{WXPK6dme@)&`%+po/%!^HO(VNKe8kDJj	Z0),s<uKF8iMgJF0([w9w@SkK/:H)	.K>;67=87pGt|U/cwd.nd'fn^J2fn};Pt .Ssy}
IiO1`'JX:rw:DE),~m/!P,+q2
n`&*i?'=7t%x43O?#5
d61dlf|b;JVj5vuN8S2',R1='Q`crz8H?CuE
y35Yw"HGPn+.qQO[{w^>#B'#F63< yp0a:,w@3tOaw<hUX,,%x)rKn02OQ6
N<7z|j<JbZ"9$#UajkB|b`Xr]KYh^#=IZ=JkT7oTaVpL7Jy3#D\Ec
9&@!h?K1vB-l;0 ?PEv3Ea&OiN{zf-'y~i9|mC:v1J&)[2<z4^3RAj=6kVwA7&ro)G^]ON<&l.c9FFFGy{	Q$)Z]\oJ6[;	Lj0E}FEg&^q~!^-}xY2wKFu|!sy-$Q#BoX2yX
'>SbJn4pb B}6h7r'X-\!~0
{fq hlzQ0GlF7TJXvq%"8i1:sCn(K]#S*p(R9z`ZjY6i{zkSkV0!0(2o=S'.v_I^d3nav JgiM)q
x~><.YYRr	2U&.:a8+%&4:v=R!bYRMN>1[NrKD	WD)gf3C=pDC,*vDy.s]cYo$$zS$8Iy-j9w`a8j*j0D>.LT2OG2YN\8l|qZ(SA#ZAq0#h[,%VTLh_y`v#` O96,htAX5kOx}8n"C^oJXk-Kv9l!Kkw-;?72^;GLQ4seVaso*/(U>8>-]0(cetiGM3 #W;MZMc.^a}X#iwrjUFZ~Qgc6
[x|~BPXcj~[TN (~?zMGqtP2ShQ.yV0+,T#0z0D'#|NB!nU(v@nR?A^3<[TiH)'FCbfx?$/^D >*1'E:jOftSNfC]e zpG3n_rK$!NKYYer<F$ktU
olJ.`}\c%E=[hH6Wr7tpN&sElC!(LI'JNGDo,Ud8P+|+31Zb,_D*xam5xNVBN~S&p9K;qS?gC0J670:8	)jfLc3 #^nfiX$_N(4ffOjR'r7M=EtLQDWSSVakMPEXQv!\v#?xYe0-B"0n20?dEr4g.h[D%NH=^pcd	8'*U%)F(4-SP%5
_xr?
I\<.[yF"!eSwy;>~?MtJt0l5N+R/pV[ik_>FXVDHA@rSBD>g$\4} dq9.,	!poxEr"J41dI4>#uLa&M9UD?ax`z!yG*k9CO/J),}=M	"7#a]OGm|u
PSc	.5LFFES(ZH	3u?%HaE!Cnn}9&=R$ct.*[/otsb&HD5,RaE}%uYbn_rZ:4=zQ\X@@cYSApuQ23#TS]X<^yP=i*=qzRR '(urfkk=o'_Gjb,UsUi"qmb8	fMHVku\S[4Ejc5x#)vE~nk28id|2s#NMqh&D1V&{w!stDWFu\eUioJpXtZ^DQ~'l/63"<+tliW0DVSxF)uXil@iU?RZ1wT'<Xp9E^s(OY/At8ae	2PStkq^@lTzkt	y$n[GUNH
p7_qU>v91]=X3NQ[n^@lhsYH'?0G__sU,/HqiW~_#$O~Ot^}-\@\J2q 7p40T%y&s6.#NFQ~R/\MgR$iC16@6G=/x;pMXIpKP$q	lazw_K}WA	WUJ7Yo&mObH_5x
ozBp}ZjnY%vpTE>L%1=($us[jJNC_tg#^}t<;Q[;ufPK!VQKDryzMf^r(P?o3v1t_4ouwMN^&{Gu%zJLu,G8,=eh<OYdFg\ReYN!QF3te[,NSXY"P2<lJlN	[^ho~7DO{VaC#<3pqjWm2vcCHD~n
D=rAG~m^=ZSW|urA@Haz]k~3
ZM}W|mz=:C0Xc;iHoVm='{OK_Z3GdhHB5/W5, [/P[sXTY6d`4Wit6ljEH3Yy_`uVq'6ew#=h4,9o6aYB)-]l8f)bSUC(bBm,e5\@F$H%,n]"Uf%
6
2lc9^"/"t/XeG'L9}Ua-lCfhy#P]-r}hrI6$0}zaIlw=7Nd*Wj<|}+T\3	T9,tZF,HJ[C=o!_tcrYQQpx|2n?;j/m**Y"F)vJ:6#lJ-iWq$W8uA|Lc4%m`=SSZI1NZ,KDwGG,C%0N9aQ,kosf2I]P=KjA}U1QJ5H{7Mz8whuN%P)USPfI&<O;lh!AZ5*BR:_mZwA6ky+TXD+qo#.Bzt6YF{j(XL|CCHkNEyW(?v+A@sk\]<7u;blGXE*K2U,He2+ p}h;)K`?O5PNkwr\\_2@B-njmFr@qR%lx~9~KK^9?X7Dd?_|jFCODT+?|n~p7LF{-ZT	
S0`#H ~4^p+<F'6sP=?f~aMC\MJI^pCCKasyX%5 3&J]/Zpo.okmGjG*ST~hrzjZsf]3 LXgNF$D0	Q(:0u$O__*LWz=r]4pz/<v;mF0~R%f	m>H:\K
S=2M+KVn'oDZdB]J/@blF&P]zL1 AI,&N.^a;JlRH`CdtM6:2RB *lK2OaPR'OuWE>+Szvhi~o<XGXH\jl?W!i-ZfW}c-1m,W?u0<o]u~[)cE7Nej2uwoTy6F,=zM:G].ZCmS/`7H>gJ
o=iE']b`F\?/Q}xZUp={H[%5Kn]azn4ccp:V~fNx;nBv?QZb</~e
/`G)_qH+*}s!%5~3@$jw"p
%Rrv>1L;{0I_n(q}U!!Xd)xvZ\x5cY%ZQ'L-?46 0`S!B5N.Y(/vU,s6y^[7yr.nd0]UG^-%[_oyi:Qr$5*,r&,MJ<V9v.Y}?,@xq&zbAZ#1FhI-\p(8#
DTt;WebiQZ;iyuO\JdAcU6-9ExB%z+Z5=v`8J#RtYp>rxTw2:(fg9B,ptF=6uW"c8-+~d.%Dksrik=T03+E[?a4o+urzJo.C0WM"YRC\spFP<D^R1h05J>@UunCrAt5U
}@:xm<\6WD`?,\%&[.%DE2B[k,"s8d0vGG^InF1EL&^qRY7.I0/n uktA `q=yH$<LDpId11n1!f.>U?69pHZ7@<+ApK[)O0P$[e(=T7;0i^h98f !<IK#/Dl:g_q-; Zs(wuB4yi2}{
dsBYa%[PP"T<l]ubD/X42rs8Ec\&TnN5;{W%Th"mm3$>+BkMw)>%>/9/5e$@qq,Sd6o'q?G;2AKLft>F-#zPP`YSU &PC@+VvZ 
6rw`_DTQEXbCGM|	viMCr-s+l2Ux9
B`yN86Vl}O?jGntOf3ODt@,eTkH`DW M{zAC"\>D10daRYUkH2>x@
~#R7Hg&t/b+JUO&hM4/eisU$T[8"!l 7VX,C{8?ma]4*rl7>W:W\!D
0!L[Z~un?NY+y`qU;;Pxx6vmp):Jn8-|Y<X?FwF27@O;O_P	G=M'8xcEBr<"EpDJ;\q ^gxt 0j+XGmd0xM?
^EYV| n)lGzTx`':tsV2V)]679$HSE+q3N3s3=h3ukb+{;lB?kd_@q.%RTQ!r<V!bf\W=KeRj`:1p eu@B&Abv+M
]f$?benhQr1mme%ffB5v(G&X}BS3)5&%Qm{xK6*t}4/6Kzp_hdW7(i674'u^>*]nVh=46xN~71o@SpdLTVR,9lV6%Ma"'D2{C<iO5a48@dVn:[Ty' roxj7'U>1QrN;X/cQ9-'RkG/tG4{2Va]vd&d6.l\9`K!F<joybpl-/q'xdLX/?L89oX7uj"F*HBHXe#8`v]{[EMl10P$X*\&)SN","XpRGv8|=:3!BMd2N*RE4l-QP@T41;']+qEx\MK2@v1O`J-'RZ"Du]K,:|v3Il#w[_=Pf+?2:ga"rRj>8RzheA5|+9q/8]64!1]KoKw(7b,8vIcji"ka1C==Y2&hd*Q!i++WYl*u;Sm4`h~|?<LC!}7^%l_1R	QOx"sjA[]{11BAOYI`~ATPhAkQsn\YMcC+LVGM^Jughm-*-K.>qM?)lPLQBp[[&KYk!|6	HC1<;_]pN:,WV`_ni*Y$?eoi+-reU!)jy;cY%P(3<!T{FX_
w 	Jt.fdh-+=A?eSy0+FCtNvb{ -_DY^OB{Mp}+"055Y>=	DlTibfshEL?/Jv,m4t[}b9\@SBX~CGi}Gchqd+@JR E|nas>w&m	^uIUT,5u%W~8n|jHYYDSjv;>Z^c{KsvTCFl({?_>gTn{/DmS$c4HPh31MGuMH
4%qGlAkO0=+raO;0Ygyt6daMW#J$${YS9pGGhZ(!W#;H+@h3B	l#n?nhP",y?Cm0{3=Be[| xyi"NPAAd76bqb$|KFSlvd7s/UX<,$\nnA6}#W9g
90_}\o[IdC~x,2.WLyRbXpTrFJ&@)CZT=W>zoK=t|'Ovd.1YJ"}?nL#01DW'*X)kK=?tl(}|!X+Ho6Q9	tzN2Y
TK^@JGGbek6i=Fn
W|	hThPH^lUb^*RD%MJ$fG8cuPx7YGykP.R>DJg3XGfmikfzW]#0BYI$XU,y8s:HB/"oyJs@6:>RqB9qI2v3\BD=W=DsYp/4eBI}~~w&MgV$:rOz4><k*x<h x@Azvj-fQ{P4o`J7E_GB|<`LESO6q<8x} (s\wBkaX2Der<(h?Oe{5^_,2Va:Uu"d&Q<Y9v7WOpR&l56Ce^[Dxed%@f7l.,ykczb\|%{$9[Ki6k5S5?$vb+"7R>aC0_d6l;3cAku'.>g];OOq>y-a`5q[
I;jfvf7|r|BkG>Ll@xaF7gc5eje7~p3qk\{MP:VT+t.Ixn!2*A^jy!u=m&MQs[=ox7|L)pI`84
)wNTkt8EZF]T1qs&@
tg/m=Kv=Itw)5PKyJNMRNvs5LHdtz{EL.A_2]auTD &6G3WORnZ$E(q1E-}zE
6!FVJ#@aDx>)80qD[w|?H6dWcy |6hl}02(*Vc4RIj=C2<%=Wt.'zt+
3GWj|a(R<C&vRo_`K-_jcVFq$IcQb`\RqTuB7;Ly]8Q!E	WdK|xnPHAsU%v#dz[YKs'vad*e%)o/Y2^D{j6AR-mz]z;1Sb'5D%)i~oNxBR=CxBQm1Px&dQ:ynEk1inK<b/9wK!j?uBK.7>J|(ulxDcuxC2b}YI=RMU0vr|M*S.9#<FlMSGZf)"K]'OIu8jA`fq.]ag($x/Jr8jQ|_jJ
oP+6N=>k(7c(%U]$&S~$K^CZg3N`BxR7|ZZv^;SXg`  ((-O3	M3Y;<S{m95**8CE%gtX_@\mKL3@uS]*L^Q4x~(Zi'~S0LF+Y!2hzqrM
PK;kFO,C]65>H6?TaP'uzaEDiiyDe'*abT\s
thGgUxGR20^,+Db^A9%LdDylP+r8(E36dA>L)#*H0P,;[re,9}m[7PiGxcPU).sc^[XyrxV>*HlJ6oQY7fj2aN(qE@;Ul}Q5h	(b*'hH7wf<udlxls7QW(Hk,0e#uUIAmb40Rx9oUMrU2YI-9"A`>CfV-A>zKRXSHw82_8jOd4B5\)wO8K. 	'3vUy2g^?y@VaUbv#HA5^4L.<oe.T[{el=MYfOjNgRh{gfbg#\--(]>[#*	xDZ=wHqx:>$?$ND(7uJZ%{x_KlJ9kxLb	tL(BB?!*#l:A-BzMP|Sfx/\@/w WI	Q/0]=zIY|HR8!om7UU{6,:	0;F%k.%K[g9/r"tumTMYoDr@kcf7VJ}pkd6)Wn:$0D{".[aG.ri$6&]vAm-<PxVN6t8a
Z|"t,=K(i4XCfF5C@Dh!|[kK5Z9iy>2u\`_8	hM"?#Lj.i:rc5 P*%#00Yj ~C(
A.<$r*wT&P&2/;A"RLwK&!wc;m$?mo[	3^s%qdDnz$BO$xRxZql/,<VwiGfxn^Mh[2i22GG.i9:)Um-NJCA~D/n*_{jJP*[]Rjis%K;k7B" QLS'(b?!s!%?%3n=i@"vi#I]Q NukQ}a*E10b?7b'=$h&AwoC!,-z>KSz`q2`etV<B.n__Q% bEt&k;gH^	f!p[fJEtTz3,GR;,]SM.Q*'bvlx 	vBbVEAd#lKh$hX$)TguJQ7qno/eZczN]VbtOf|ZkLpQAfZ^
?vBp6tl\e2uJYQ@GGdks-ihD
B"J:GwO,+(xUelh.W+Xwi(qkH{|L*+|H1VQm)*uUtG=O>'$M/+e) >\U0"iH[5@hc5;m?;vX
y}&Wk{tV].w^
eS>&7DAGz\Vc{\0	{A
.B`xZJDYXrO<};|>HU0P:R>yfvP9r'`&Oo&p4d

d!Blm,%BR!_S6L(!"huqGRb!hO6=1^Ztn)bWI6#*
9*a*;NFtL!.D(AVg\d {13v9ByL<;CehK  v5-1	AQROTSjJOWk_zSVH>v&)"B$VhGO%LX %>X?	dd9[x*>HAYNec|s#a3|L|5b#;iy?bDk?
H)zqh%>NK.
1RoOisg!gV4^Dq$Ee?m+Le[=vZ{ Y\6|#7Y9'eNp8|(yMDtL{M[Ei;BK,r@\.R
j4TW(4^J$:='l >7QZco`M'6dV]c.^Eyf4o()M@je#qs~N-[:,uNsQsvH^ Lp}F1U5[g~,?$L~a#e!QRk58kwqRBYtG6K/|vcgVuW0!G,<XN	1+w/<lcZZtW[$s1VZWL;G"w9nzkQc}|t`9}Y:vg]QdA66gfo95'oL`O(#Y}okgBl(Kco"EV6y{SKy0Pz7e0qDC5Og}+"#;$lG,E$^
Jeu7/@Ng	],U+Px,Xw;pC&r{dV4RofF%%1UB3niqHxPIv<6hgoM4\"cx$(7Irio^`Xq:Ft5_4a-N;3Ee
	KH}@[\oR\{Th@has,7@OfY;dh;X!KdE)E>0\~IkLV;.KG|>f#>bhqoc$	\}]saB==d
';Ls|2|h	O($ruS+MxCa!tEK2Q/s #'mP4t--Y@-`0jM=8w6U,]SF<Ys33l@;h!D:U42_7w{}A&M|`ZK1yM=])yrluX,H^4>AY2v]?z<w4#J7k LNU3?a|C$az9c@F:ox
-'XaH7a
ES=s~aLEY`${tHi1kL{f4M\FnO	pxW;E<+NThc,e	F]9+<v,R>dt%RUI=_r NoH^IFq?TExz-T6c\72KT(G-Svz:DucIOgRizX#pG }X{`:xLf?]L-zB7M;Y&/Bs`~TToq,nO@<ob%(P|G{"ak!]K"g[hpTDJRL0_[P4c:G, .fX/BHMbiPE_+QNH(k|jq)oQH!XfC]wg-Uhh+!mKwEA:K#39_JE;vOG5u?Cz^*juiK?G' `Qs	L 0*:[y	3'8^9!~Y!OF4\>LPXDe4r`KQL4vM	s#d7%Lv/(*Ov8(J xk_.
ayQj3?G_]v!4+gY2cj5/(]bZj;X^@At{\tT$P/)61Dx6{Fo;Ho2q_#S7];&E4QtAWhsILns'mVom)7hS'Q)O\0sp.Vi#\{k|U($L[:?$f9il0Iz936|{|HmCeNtW0	uFDRIn
z`f2n9}_b>1j]#e2Sf+3;+=!2;qaXC/4h)=/,{T_2s;,RHx7/;X1IuY+J2D]m_
#5CZ'")>'l[B_rTa*2~+drF7|X5*Li^NPo-53wNtvB^{2K=Q>2CoS^YP/x"8p
F3r^3UbC?-ZTho7Sl]HR|++7.8$zUN.*wZ[cR`iLF4pl6-R]ErS
XNjzy-_'+[lW7;jvrL8N11HHi|X0)eSK.-G68nHqjB
KFN*/6L4DdnzOHA5XT;raqiAN8:L/,IH'N?Bnj0)kI+[WGE,BN*Nd_%ERnnC0.7%!n+(2wBL+OBTi:`VB\{'g)vV%b^pw?|/~g]33IT	>Ci0nPK{ly$, 
MJ/3[g-kZ<Uak;UXH.JO'``ip[#?24X]c
b:F'f{c~TX)i+X QyR.' d1;lc[
25[j=<7C;^Qnys'qZX}cAZ>6GHqYXd|#*[CMW	$0	'&3E":CJjF1x^<gXw^lSqtbn_6&1L	g1?=T=F6`_ivW))P8pmQg\vdm<]E.pQ9ao@	i,n9x? Ea'=Wf>JB~;CRc1P2{&<?kOJWANCHx4}1'q'U\w;0rWW%eo	L69NR<w[g!LAFVw%3KmsYkcLs05w'Rn#bZs`aM4Pn$IV08lHw7=oHbzL&	MAM,i]7VN4s.s/D#*Vv_r%eXSwxD$s
N~1p3*."3[SL]-LCzZpw:g<BwyADQ.Ie:._)>jN]l ="h?7oaPL6o3Kxe4l(@=nFpi&-I8Ik\DvDN:Q&_sj S`Q*G^&(%RI%(*sQzs4	xlz)?#.XvqOWIaD~(:D4d$=,3"qndfk"$O3Xi,b<ekFv'7-v+C-B~gK['hyg5b8~NY^69\i+@}Cw/kijZ&a!od-"e[.c3?Fdpe.lG6 tTq)V= 1bS$(fvX`.n{/ Bmy0(@]jb<|.CascBl=dY3Fz(+"zTs`x"0,j#8X^FdpX+SE;B5m GN$M^1V5
W9aApt1^HUu"okq4?+ kZT&VNNNqv;mrs$	NM*G?=K8-}sE'7S4b PUPNz:UD1b?k5s_kc{1#w?`S^I7R\'T_-nCE(ITy?~_uSb|ov=+%>W}dhjbvjS2X# 2N4!.t*r5>(+9fw)u;yp`\-lpw\[ |Te}tU]]b{*
KPX0R#j+^u_[BK}W|,2_;+oQX\lQ+zHVRj3y{4A~l6/CnfV]n($#_$b+D
	82r#gtSF:&[e>}b16)hO'>-(dOU=^kR,(z[DPkHm^1yg1taAmlY{m^N0(<ab(+Qu`7^{zw6"u?b<6`L+Bv%Z4]=9Gavf>}?f5Ie%D-s3pDl"T)[6!@RY)[	d`7NszClGWKz%1 }aKX
w0
ZHth:fliDdCg2#Yk#SiX3E?nS-nn1nU
L
VHSd/@zR.;eV-,vmt9T_Nk{/I<O:Fo="CM2;8o3Qs6L2yRvx:}f0TVd/b
.g!OJ%d"aDK#v\.w#Tf%60#XF`<B[]0;TZ8?ae@Ex;7;5?0+ogl>Z
w6"!$J)Dp#o%R{XZ8$G6Uo9d#2\KQo-=h^vO+OKHbO/Hax4Zy[\V<o88'1Wwk(QCCVbi[CAgOJ^+pNK2,bKg>TtS^,:jSLO$.0$fdyf}H9<?'2]V6^ng/:lnNd-H~-L@=m\PMN}x5%1]]0A~&:]N"0't"d4;R9[pw?QM2:a>!2vhN"u1Sqk3_J/kcq<Q)'	9.Or!kyKv!>#P11Nk|K)c9|=(uxs~[*b?v\'6'l.7Z}A3k	uX jWCN{"y&V^lQaEn]7{|JRDO_J{\Wt[|z)B<J`}s]f+k		<Zj}du8[3:?>/WFjffE
l"JD@1>*e;|[P`0pAS)t.Akd1D4V*Q)3--@_P_LT!6c*r\?+jD(UTN\#*N'|L>TS`]'R*pWCL9}AwU@,2je_Ej/<z\b6W6G	_521dt3G\>	SRJe#V.UjYQrj#L.CTnG>W3cCe=09Na9rylO<%K=N;eE>'py_Xn:ms4QRg'
f~]|j{VO:L/%'N^xDEy`S	SxU5J.(0$Ad9YJ->g99[RPI'6a<}V0=qiBnYp\;T&V^rL{_e\)c^GE{viJXeui"sL@b3|(6Gr{zsQn
TDcg`R{=ta51u|,wWzb)gHc~f;<)I~3'uF41,mz!-[{O?V:tVcQ]lw@YKA$j`h?zGJ\O{)^e9(]H*4WP /8 2xl'v%9z)r($7P2{%[smbc0pDGVFWTO3_w1VMZOtfO2wly/VB\hbWA'Wu)ehfsT1,V|+EPcT<'4t(
]e>>JH9Zo.DvBGiSAtaVp|+Ub`R75K8&3g0E<~zFR7%Vl%kdq*jtpO]iwTDqTtZ^XE;7-f9u^Mrk*d{ yc<sLI/KzPrjLj!=5'O#Pwa{NtTp5}[Sg:t9DY{C3SlUw<]P\'qN_X|b-d?]#~0H1.g4fU5IS&1C;/A=` u%}F[..UCf&yMzy[@J+)x)FUMJn.='>/ootC?)+J^N0)n#L}[q*1)60v@K;Y*unPB[pnlH)>%#*_9<dZMNAI6D/&F8Z+N
R|X)A6bc.rJWNQe/dA4^nZl:pqt%|:)E">"j.L:=" z]fuAq}cV	|q[9yT^gc0|o8q>_nxbQ[Li\w3h\n18;#H,RB>Id0{8U	f}i4!XWMs*0PXR,t-ock[XK5q
hwd%.L2%n9\%_O8,^;FC;^46;?k|2<^O_0x5XAF#y{Cq,g^QZ.h9pW|^w*TmdE.epkC7P|i2DI7s1.l4*\-[p|r!HwjR*o*3:`drm]r5ERa>+@_jH6F]bak]3l$_5r>:Z,`ef}8!m/XIqzC[j|Ja/@}|b`4OL]#Ra,<Y0b~|yzo^8A/YZ//(&LI3PJL]k"J
#%t&5	-,B\Q
='fZJdbx5zF^j/cVe\s ELb`gfLLuIS^/H&B*9#=BrZN,5^'wWnvc?CCh@tYt0C[]LD%)734?q8^aC'GAmS9{_O_On{C<[9[T&@_&HP`g!{_3V=tX=.Qa<bT'~&-NW!=Ry-nP92@t8:J?
`Pl7=>|?%`A{yM_aN
02r%Cd?K/aXUfEpJ\k=`Bk]!5W.Ck<[Jf8U-gkhq]W2]'G9ig\P^sNMe.;CTjN;
Wu[e[sBWO&#vG[k@)STywQo
>W=5Q80jq)$_	7>4XX>*n0l+yb?6s/xz+gH:+'ok3Cv?\Wk5=4&1Bx(iw6tl~ ''@MY)*h>3LvDeyrz;&`AOf^4I~:[BX;9>k0h8{|*-JvI+VTz}%{Y-,,U(&4<SoIOK|"7	ZWmc8_PB,}QIbAx%j-|#!~blPVPRdcZyJP.>K62Nb%^|bm%#SwB?Z wNa$6R~'+Vg]7mc9eJeweX/R]FopI'>KOYSR5%-+rCK@St(KD9a[i>$`H79;<Mhc{l8sS/~hSO<K_8[u/./Vc2BzUW=8an94qE/liF>,Xi8p9![X`33''n49
+;[q;]^eFVmMEE| FQD>;Na4:.t2f)J	sp8{5m>6WCN+4Unq8	:dh]'JC"EA)*rz,qP]}S%x6;|1Bb53W9vB*B}]8(	hd>xttn4vCK+8M6U^Zjl t-SmZj#dCDaf_G7Kj.+uuF}[Y5/aEgw	NV-d*eE+m)&4@%\qntjX"'?68?z_RNnUBv( yq+;_zu_o0jp['TfxO D?{!9tklc _	@)"@!F:/Pck`tJkd+,d[|	A_F<l7m1Cp62b2n4Y#103VW+eR;l+7_Z:!/JzESt\jJ`;",~ueg4-`C']oJ:nfu/Ovc|lDF~[lP^rpm;Yc8*\$+Rs<\cxqa/6.w/Yt*0 C+fO1!ZOvnK	B4:348{YIbJ2GAwWZ9^57<.A.9'|%3,mCT9G`BhCpl69	#s48-U5w6[=A>pJ6Zax3L%-
tYk#J%U"oUq%YNar:.RL#|;:FHI1gMud<=lE+3-]Z\%voouvt$u8t%u{H+gK	_4=\8NRA'6Z^mJ/N!fnzeggce$}/Lx;4#l&Qr>g1=OeVQKz;?p1d>LdRmMk~u
:HDHqKzf4sUe
GR	R}Pdb6OlGQ)(gU?:?	//"b?2o1$=P*x$GhSQ(n3w0(c3CGB((7B`[_B92Y${^M&|qO.Wb$?r=$}4F.	r\Cf7k<%[vF[C("lAJw!@u"[m_j=+Mu_UKz%/kcQhK5L\Wh);;>I0Ai&x84/#L0Cje	)0/+J5G2FMT4JhH,7U5+X|=g@^wnxf/y|.XC)luYkhCrK"i  Nj)>B~4Q?il)k3nlQ|X0@u"!t5r
g2/vP(
o&$m+b*ktJz<Uw[O*K]v^A;M@17&6[zN{z,%6rslVE0b^us?2ClPru
j]S8j1yt7#j51ZCrvb,#& K$v+A.A"2Wy.h_F$sT,^XwW2BY9zt6ST`7.PR0n-*p2Ljf/r$e+=bq?VA+=hKwQc?H6&B)$<c+U9_L4
uY0hXZtT8$<MX1~Aa/Pq1x1q.7q3(g)liib\itn!Wq2-zpM;!cglY	7^ucE/#3y._"5ui,'r`D&_F).mq	'EGY[;ivdm3]+P5F<kz$3jnwLTj4W6p2jkfqhKA4#5lP&j$`PVOGf9EL:?&j]=gu`%DD#}E0@r"sIDna2vWPG9UEKDAYS& B[vut2,,H]k
3+O)>}q~HvRDKpna0]8ctYcM]EQ,9`O"j!(nuJNoa"PT}
0E_e&O3s9+|LzI`1je}Y2d(MiAI5#B,gb<yetqkTiJ{Q	=H=5~n=GMdWm|99Fg3Mc]):"~Kp(|NN\7/+\Tnme4X6L8yKJN
Oxv#4{<q&vf$UdAJPF4NB:q{-_&dBALdur\Pp=#rvpQCR#)gSC=p3y5CAh8|q"`$s+{a96MnZ|.8V>=ToCVuD*AV;`U7:=A^}$-*%o]!>/BU8(pN{D	qa V*/l|5)ZwQjDc,m5\.d|OuWTh	|1"DYj*Q*c?Tqpe'{fjRJ4'`I=BBDOutY2q!kQ_<,F B[z)^a7~K#[x]ZiQw(Bf66x+m,hI}$@>YPibq.v@
n'oawU`YBN36E}C'ojyj0edZ~`}#d1']oyDfEGew+'m!8j!O7/jQ(t1QN RL\=# Wp<Q:}ChFD0w@&?Z`t_}b}&H`s
rX'c`2i3>6*M2RE/fW&W{ow~se7xxawQLZXIrP@-r4|GT72-'?1(8nlD
hPv'*5&?Jzq
q;IE<-	/oZf'bj%$T2fj0{UXG!h	`
9/WE\8}
QZH?X5X\T>NTk6JE*in|tDt\R *;hc!v
5x>8P'$m)]OZV?1[PBheP
|nuiVg;ABgpA~@:mJw`i5)+Yv!b*MkLY~Af=!XUNJ0h`$)d"sY75_3ggG1KVZdE6qQhLI9n,2JJ
kNecCQ(q\A-WEjLc>8K,7PlA<xaD?_X5t|YVfa-^>9fh7/sg2B__ul[xQ'Jq0NwI<D l@Fpff;z=s:2_T47S<tWCf^{vY,qmHY,!?{W~LdZhqEQ7sN9i`	<"v4Bzj|vA|j@1XA\],Os$#-vd2eGQ6G$xqsV?t?dloaTK^lb9P5iwEUA#=p'+<m>^x tN!V/ad/N:WUy1t`,GBQrDNb#?W>f5:E
@duXIBnnHY-yFmkAv9f'=>Bep^aRu:e6`#=3%NB`GJS!$k'~rGc	H=I2(!$ :?BB-n,2cTAfBNLckd{A[`iBbh??qJKg>/]Q>`h<eLZy~d'h\=HfFb0!sX{GL\;p.I*\HxRfSV[ec4C*9v85~[YB C,;tE$!m{GnZ_2@thLLifci6&0	_heflA{2yM%[JCeXGKKP- ei"$Y'dnQkAhJ5CCfi*+Xe6;5H6p+)85=aIU=Ie*XR/eimjfBlHiv)@!Rei]bqRw:bUNmUDkJaPAh@%m7?G*ZBPg{tha%*~{LyD5!]HF>_6k]YGY^,v`1IEU|Gq.o}+:5F}G=~sKyR/VPx?eme+!Fuuxmu/>2'#8Z@=/xd8"P\y?\=<oC
p>ja#YrWvc,>Q] ~ip:6>#DDlhl5HaLwgo=I!V	0Xx*2^Hgi==r0|l/f~{XyLXGBB~RB`MtF_(C\tDvv@Z:?d	'+i)q'BoPC:{,<:zdWR0-Q
%%7pG+|RHW"QsW@%+=P*4[ML`]R%\"LuIR% bek_U7icEs."M\F,/Z/9yi>WH}-q0]nx%%}IWH}_b*r7]|eS'b(NB3ni^-9I`K6y9w54F"?_N12aBHY>1zA=JEx'd
MX*>ORP,3poPqqbpeK>SUgZErr2k#'y'f5zX ,Wh"^%.tvl+jSzz :W=Cy[Wo> =-nO?wto6@SFf?"D_{B_30ze#W09+<9Z{?!nw9;Cquws=wE#</&~.{dqI)p>RM@kMIqVu1N3~;OfTe
W25_^ecI=bZ_I{	nzYipcT6z#Y-_=(\qR@'i(	%wUzqz&3JiTbUTypH$sfZI>$M*w\CSaY ]`f	4AGidGO|VZmjg@W29GL$%7VJvDw5?yKk\e"s
8..u08F`@ lv{h`Z?W(\9H,Q90zEI;taw[dcu:pV0r]C*^z%e!sLI58oC03p?#`H 9=*oDb#Np54n]3
AhX> AGcMqG)17ohq_xBm@C66!1\4%5J!EMx\pmU;vTay:at!GjZ~xjjH`n[R"R|cq3Q[f?t(>feBk-d=kN8(Q30jv}~ObXYSlY+dOoB`_$zp&F"XjmrP3,Gb|jE{"o`TH:S
vb+SfB7_Ng<ENz;tH\H3w^b?M=1&QoHU9xKh}X4+ Sw
bb4_93z;Og
Pda
uUnS;:zj\@19(B%RYXTqw<*%vyeM4 /Pq?j]KV563GgJ<F TIR4=BC
0{18Pfz8RA45R#4\#:AwJ]2Z/0T^:h7w)Y
`KPRlkw^uNKfb%+2s!WQ |"Z/#vB)rL]t*953hti?I.s#=hiHo<tBfHh|>wWQmP.d
yw?O@>>0_CTMM%,k9!Z:A<Lpz~\OT
Ke#idP(f>H9#(}~J&nw`b3C9P*ES&W=bh2\-0pX2qL-Qx0pN=1Xo(Q?^;daGHRjwz\D	>npGJika7KOSWd-s!]KD4z0C;u.{\DQ.vzCKKn}LcNl$d=e^v:FB^=3M"(dV*"Hb@GT`f}5]'=s|L#`ysrB}A..A#bhx1SEZ/5~'oFPO0kfc1cX7'B)eH'9pF*%C[?:cNW<B&e:3*05{dM<CprNG4	A"EktZL q*0a:Tk1*na(i|lc+d^}Ca_op(b)=my5<xi&Frqx^Ti)mhUo&r]O-^5i}$L*+kee@-0i;EKD%SL12]2^e*#=m={#_B\jbw5g@:>&bMDFIG_85W]P87T<R=S0rj5=c
qtvkh0KbL )sA'll}]Y<@bP7,HS^|b7%DXA3f.'#Ol?Ci?tzy}XC=_zlQ1	k)Z,O	2ldb8;96HJ|><x"p"Ur1`zN@K1dpRV_063LY<OxXvt
Y7W*bIL*vW_B>*z*^ii8Pn_4WRvrC)tj<(
YYsB?|Z"nyYQ7aL9kI,^mlnuv`tkbp5	Hb;yQ'Y1}6po3ulrAb}}:,OsV.x:=LO
uUR*f^3VgXb:AO@|+FIkjMR[_Jr70B$KM'c!:doV<
MlzM		>_}U'c[!^/]8DTP/3-70#t'v&l%[=W1
d3>"LQVlR_pR%)LHo4btmHZO1+^qTSyWl"F;10uv^.h(x]'4[!$z5=s=4DP@35;0>1 wc$gG4*X_=1L.wO&7etG%i]9j?.>{$Nv;]P4i5PtGP<?]S]F_G;7><^F1d5?USy!c/@;Qba]lE]D~~wwO#![x1c,#.fy'ml.#SR%:T,w0So~jG`_?JLGutbUW@gAG&W?Dz4MV=G6gWaGBfJQ,G=8>!j~ J6FO]`^PY(R7nU\GrWGC4=-'kkr=fQ4x.Y4UNIaS:H
l"x9&rL7L|E*Et"6S0~	&*Cu$Y3uY8,+
Dx'p6,7
oA!~5f2>:Xf$(i_n,22di	vC%-UGGa!b^K0nM#n.GJxc8MiE3tC!I.|vu9|+8kR"*xKr:)5+x,1jFK@2{t	1yX'@o~N[(ZGK|nf":D0D#"5?`%)%oLRw^dZ#__Rk&
oWNv&B<]AZ}<-=d&un.1b.O,q?2@=&&(busc1?@Q;<Lz+Cth;hULD)~ zA/./gw'jeV\/]2
kyXVyS#nVzw_:b#3wRs"$Mt+	k^83t=i2o #/Q8laKxx1@q:dhW<|jn&ppSB"El%%1#R/&WwlS}np2_]!wz/0h&;Q5{Z4r7>rU5-@yl0hul?ZUBva$Q9SDAO<={[Nui
>ab]ovlJIfi=M4
'5ZeG\`bJ2pl_#]$c tB+[+bm|_ }_11^i:MFcrMR)b)cIP$&Rm}8AvD]3?RV]aWX=#$LAG\&kSf0O1pAx
&v`l3z|!0$ze@m/z7RH~g.g=\Z`::z"\{z"8Zo\8B Y9G$-We*H0KM)rz<hhyBbH0&bhSV8a7A
G<q `C6/I:zGGa^k9#>a*H{]3+O'XFqN"I;*'Fi~ot6UnJ9)-d6!^!^5K	e^,2id*KytveFT78c-5804\F7,B*6.dgdjR\::_)V;W1)1f4i=hJI?,13hUk`grdX)pO)AI="0OOA}Z2wlI;Y"Sq*(nz^x$(y*WoO`^{o'cQx7Iyn}#hFx	{9((J%b4O|sTZatY E\)0g\g	|5TEHGS"(dFVsTh]|x)E=?r 6*$gSd!Cw*:'LZ(t@y+VF;):rT\1pbg-rDrC#5NgdU1~B<=Z?m%\r'WX!^e3Ep^ L1:+?/?U^8 ;Z_j![Ole)hP]#>6A/+rR w}D[x:mrs=YcsMsU,d*N.[m=V^qT?8G^g_75m5(rme,bdcVx"?j%#7& <OPF9!z(q"UUN[kxX?|yfZZta]r?3p2%TG@<qK3@)\M
s1pWu&LA	`GY!{B,nC)?W?z`S?cko\hbkDLgmYK{p)t;;DHn!@u\eMVkG'e@zcB^~1=shL;m1,\EeW^{]aB\5uo!tZeS8}}#Q.;zM5
%n!]k6-%"jMH9q11#pm2-b}FVcO:,x9"H}1P"8wUahm!*[I%kv5B$Ns|s?t3R3Mr	:kyD==|/n3#|fCxRaR<1/GFM%!6q7m"*H!w"K<$e<-	2HX%dX_?[1+p6B%IWSv;3OXjLSxgnWr)=bU-&iTA"5.FaV)1_m6|~?bQ~Cy96oe:y_y"+`aqRj/vW0G6C(E@%	]$1>3=/O*L*<\Kks.H0<"
4w0/ej~_`/: KeDH70v5G_.c1irpr%[=o@,W`3C*S{@}jF9G5;X{ni}WQuW_V=!W6|99hpnn62kQJ
s{sPgcuI&tetAA{q)|c]$;F$-@)Z;E*#EK.}Kh";1%c>	H9a}Gv=u@yt9@d+ m_	C|)pq]yIg%Bc"hUr[f JM+.0xO/-rl-'`=#zwg(<)[KF,
)5p(	&`knhCR_nP^C	$	 3{pV^:/
X|$,#1Nx.">(\Ro4(|:Ig7|xhc
c[<>%hA)
'Km6CZm6Q]<ha X<jTVz'Hf;!OMPTqz\AhTuNe(LlVUDh6iTnPO~No:)7hi5	tQA>](^}+N3],=JcFm#/a>s\QolkV?L_z!-LGi9NKq$W;F*U:j{,fUwOts8%u8L>)9N#Ob$VbY!8xtL(J-rtP0nNorCdJK#_(_0	N+]gd6L (>3N62PQB3tVlC=}?$^Sv?xDtu%sdoU
.gnV)Nhr);~G|S+VMD$&7$Dcdq0?dU8qoQ:GlxIS)NNv2hSv\7A!BSvG3<MNT"/K
Xb&/@d7n<	Xfh3K(] %f$">,G3MBlW~gn%AMUGZju~}>RNH9il!d/[ORRY5v'
W.*_*Z0]g8l&vp\ci/KCI-OEAs=Hm%Q}H)"I:wToRBi	9z
jCf]{Z43>nHn.!5re.G^#bWSw`l se?9M%?zc^B;XLd|)?i{Y`)wMN,2fGLr{~{'7F)h|-HM.8ddWrq	CPZR| dZ31_5J[[</qE
A$L?9+P#9y&kDYe3	k1mK#\C&?	GT,C%5Gn@$x1Z!&vy44Qv#16Q@M#]{bZ2wdkH-v^7"iQn4U](Jmv7+<TFds!Xp	E\@bb2D5yrn "QPyUm^S#f>|Wytwg!!{R2	3{"`J>tVs3LCFG\0 +e|O;wy37vb|=O*Y.?X%sfq_7>Y1<Z	Xb	f_*$[Z<!Wpyd8>LJ}oE2cPOWD*dXoq/.bvdZ4:wr)*@K6:GbPv=~R:k1.AKL[+NW.tezm0K8F`+.k-aAi,Oq7oXXB:53=,a5J[I0ejnB|XO*/^aS7H&lRtcX*J|(4
!F
c.M~Dx#sC3*wTMIo-u:1:gd>OUHQ^-	tp"C!F-1^?Llt=]EBMh7/pR*R6Cf80<;]jIF! LzJhS#i0K;90)*TW9f^} -tFHr+ti_1g4V#t"PetMPU2wjqP6$%iPh#cQf8
TyeOQK0t@0Vk(#/FTB^[j(QR_OB4j+:Z	WL5,>`)sD#l[S|&Uo5WFA(R'MESX9TwPQ&e*kabIvU^&{P>*Xj"=xt_RTv(550a-=>RZo5A5Xj^nyne-tZf^q"5o|~;X]-QN2d>!uyzOs
R3W?fe}jN8lOo)$s!6rzq9_Tok(m+@6v|]*A_pOn1BBrl.~GQ%wPsO#VL3-rS<,p1aaD,6JPlT]g)+\Nzu^P{R?C"PJ@
_v=
kH1fZNw$aB}F7a<H3$qs/\%x,W!w` 
jn>OF?T,$<*|	}#W3`8-k)sj?Q=,2#Z-8QBh4&C$YSIa)6(fQ ;Jm7^1vYt2#v'8s_/dy
bi,")=NU\>Ao+Ub|qW|!( b`DPcc_OsUHo~x8b-lY@b7N7?eZO9j"7@SkYC#42?BfugoFYVTrv"FFl-}mioBaUks{X$5Dlq'CdR^w;94r=]2[hysc]p=]oPDd+~xbnq:A2!R{:c9DIbZR]X(=8Yh'uNDPQgr4[u&oi7a.H1yr]doH0E3\7vDBjLxlM^<=)3i2.2p<*H^zAE'MuQq$-TQ<X0^aN{[WZeP3u\lw&n,(ryL"_'b=*?j^$o2Uln`Q6zE"J<u/~[8/PS'S^rS}_|&P'YxqaD5LA^8|Wvu0t(p=gC)HZ
Z$\=H
T>(6}$&Vu`nI0*aM~oBr61X1Z$8O28v}1KajaW+T/gF7TfucGTcp(uU4h;AK'E|DLAp!RBzr4
AWXxAp:nY`XB`gE )mo]&Z$[NeJ7bA{UFb`ws;1Po'"<_1?oS8DR<Lc';Nb$?*N:	aA4SubDhi>%5OIcNH,4e,,5:JM>'e>X7d]L;@5)w15*oV#S9RES] .^'-br{HlV!gz$%T($z9ZdO=-lczAkjq4k./.?!ej4o:*?)Pm}{e(;1oW/_63D]z30T=y}l\m4BPp4)HoJwF,TT'9k9s04VG]
_p#u%	_'}LZ;-E"<0sf!(Ko6
''E/.o'_ox7M7;\:pmhxBbs./WfC\U80<ZFH(M':|-d[}\C%+pL~[ybLDw2MS	9{O*tYxXy!&GY2	bJg@&\
!U1PXo+^b(B_m^wbMLJsOSwqfKQOVj*WLA}#jqUQmUgSd3.2zzB/ETMX|[*`RlfX&-FH!SI_]#*1E{kRs{.2(w=@1{)YY$}NH+dnKO%7NkEIrg7G6yf8(`/C'Mz.S#PBEQ4
t+ 3>t>$ qCPCzVKOy+y<	G3_8TQ
 ?xKf~ef{oi}L+vY<bnLd5y4}5n	>u+nKlQhVRz,f4tm.mL.ACqsv@mjoH[']o"TBWO&20YlLe1+zG|GzAIYFLhB2P8jY=?$YUdW,gM8kna?VWdc)FM4MvCTv@[5Yw=nl0gq-7wl_Q8r?<]>)wUKENvJscr4:^`O`R,}h69e*=
;]?mdm7hkW4;x@aQ	#qDfbPLw\A,UAq_W/aEvbn[cFOUPB8u1dZ'FDn`*Sl.$c4@KMX[eQv(\u	#Dp9	Ob3-@j4H0pnxE~Y(cWo	v}X?K#}g|VYM5tBT-G!|2d):w'P`gs8Yp	e%^1X&kkf$l1J#(/d,@<0dI_+NA5+-16rT+^VfaIAr7'0pwD)^QLcqcUy11\^fjC~-C0Qxb-QM`<m+/8]d2jCKW Hc9p\W+;#^"d<970Qx8gGt7.5	p&
'd{ZiHv'1{atOli[%DH3<4c 4/,d	;t]q8?w{Q33oWL:=h^+<we|w'UfR'xxwi.Qk9aL}[@:}	,4/Zb=5X4{]mzT9DT\'pubf`#b;q)}6=d!40},Xt&)[hL
5g5{Yb*{sc%Ja)$cRB_HJdObnyQ]*=`Ul3HKTC68:9aXsTthP%wDR|VFP6yir|Bfu?U	:B%pQ@de\i,QW#&
]udfp&yL(av7Y8'9)S ER([j$A.2Jv&-m
;s9#'tnl2{WcQjacgUk;Q`*<+ZkRXn`Z2/PZDrN*!!jZ3NSbgelp3oCwPTfra177i^HYK@y1Av1"FH$"f(]fBNQp8WZb4_8/4reU1s{aP(Bl|!i/t|_A1;=0E%/UfdRAZX1l{=cl3bjbVX4P^d%#NWcE@
t`Qxwdw(I:p{K=KecCl>Z+w;6*RP{^9>5
4-].+=2L{X}Xyy`2d|sV"!vz%}4MTsKfv*r-)%*thT^}M{iFgEPJk00MI^Zj"!\WU\I1>!-jrGpy%>	VL:e9fe(BD&>b}h`=+P <17f<by:3%sWD6rs2QA,)poZp-T'@4gn,K!wZH/p8E]Zu?3iQ>JsPp=F2$&dh7MExB'~0JX10"SVNMAjgmW8~re8;q+\=Q$dORv7Q!DRt0Y:uvlL(XTodhX*O#c=A8t}!P&qQI6:!Ov1H`KH&Cry;cpv0.DH :YF'.VUZ*^~~1KWv#C"QoI$F!47u; @]hjgCj<G27hKlw/kKCROJ1J&P C?Lz'xj8fkNuLoBc.~")PdBLR|=~K&4Y+nb`[xtG;-rJS H?#'(0V-:_V#w.xO+clqm)~4XJx>Zkg/9=*K3oi|uNsx[<PeJ)}"VJb:5nB"rELAB>B8: i"f?oQsJ9*F3J=@c6zPq|t	mzOX,i>hqI#
t=Ly;Z a3?oxG=RKMpbi%fP?>";XCDs	p)%HLM-5~vyw1ABFI|.x 8FOo#bli=bX2|1o0QG(.u*"EXR"p9@[U(Pm8>HQwdA[N&66<]SShj}~n#4`z_MK|P6XM;,FfzQGQerb>%e? Wz-g\,%9S^ih5B;T!N#>%Z^@!_Y1tf{(SKT9~Vm- W_(I@,G~>r;v;V8>t;PwZ"=ZmG>=Fw5V,PxCw)kiHoD*+JQ$lkJLn_lD=RX1
1<%i_f3mT<UO/|bI/_>C\'.8tTJ8	<>7*4fnmyZS$v"	l
*6#G)[ZK
:-nTl*[73\xZ.O3.$qWc.,I6{7ev+vwcyK^SVl9*Ob"0~p8:9k^PV{p"i(F&tV!h>"r3d8aLK~%.DK|xng;dYIzm'bZ?=mKo:d0Q'I5DL:TIM*}'oB	PjC:)-?F=JD)3p(wr:lUx6gG	=Rn|O1big@\Ux3T:RS
|-\{$$!UlUwbhiP]Tq0~1TIE*2kMEyZJ0YYj4{zfm;J)iUb6=YnVx`KQ0qh,a~w)yuV8/t,:WcK2m}r2Q	GciD96.}*LyYy|9A"w7_yOxvY^<l
&/Rb^	Kbq2bZp}c<_(#
I[Seo;L^#J`,cFKMO8x}c:^Hit\c[;i8\X9^V2D{v?qw7tAizOW
uf/s`Pe'NK0is(}C<WCtt]IAMDkM18dcy>Br6ZdIag5q'@D2n\ =uSSHTT_TxUC02VS!El,w(ni1A*GSh!62M}); \YHEP-$N}w5Ocs=s.U76Yo[yhGU(%|.e1=Ra\K]Xy>5UGX{<~1l9	Q|:iNeKOh|z*$j*|BLB\u01wHB=uLgCFlpB#Z*<8X%U1Np^0z'PS9ahwIe<dpoyGe=\?!RD8*b~ZF;vx}X.5\_$Sq
FO+&:-!@ADL\^LJD
XaRO8!kK58FHG%TX74mrL76KF P"`yj4uZY
9nj%N)wQ'2T _4ic~Ems{ 3|j{jLbL:\/Iw,N(;v?Qn!}I"\/NI>BTmaZy,OY5S@Mq~ggwx1wk-uxx-piJ"9UKoboX''YL/.\lEew]"p}?<A`	9JOdci	i%(-Hcxc	w1h`X|)up`#!,S ]!n2[P&Z@yg"j#Ec)!C1P.NMAcdHqE/C
ZlLZ(O	HT8k2O4E||WMm}S/pV`RHX8WnV|V<,@nMR5q#'}6%b$=gr+JG6}K'/ W5_2zFj&<9Ym:%J~pLkd&EjfKtdYb0Cv$Efut

1`$D/~l"]bpv0.|D!Bv;RRdYF-_{cxFcru.\Lk5:/;ha_5X4I0lYhQ}!buA*X77da.R"F2g ,3z,Y"[&--Vy0KMH*x'5p@p)Xe*s_n2y/;pavw>x2j*Jj^nQ@{V0a
DmF7C-&8h'|x)kBVkKg}6Wm7{YYcTO&OJ+|UVzu<>'yBYyv,h`7:Q/mu`
2ECR-VRo3}}NNdM{lxV0U!05ZNB|9~?mva*a+B34 '0<3g"[dbld5J""n)6.1<4Y/{<??kyeTn%Xuwn4S2{no48X,b<\I5AQ(Z=H]dal&$qB[7GR
6b4ylDa~z8q]eOSmJm@x0LflyY	E0taTit&8%E@s'iF, %yDdx`fD]P#N1	t`![TU0*H4GO#.UWU83
Ti%D^{~'laN[+K<.#K=V
Zup&7Pruf
4jDtME.bH:z""6bsX>Z{/8WT/a>O	H5%;~~*b7\_+TI{c9Zl)nLY>9g
(/B8LR>cfn&mKjUKl!=jliP =c4|%EZngfZ%#BSR3	O*YP0[l
/~jrCP7{Ws=j[N:\	6od$HHJL2@l$2E:cL<=>MSTTekDkY@8YE1<+PrBLi@qK"yrtmhS/wEkhvy`+2LP?O"E+RcLNKX',~}"?X;h*Ed'*)g}+>#r	4*Ig0J.GtnFK@"`bB-a1KZtGo5w3={}2~Zeng,t8XPjiVX1+Z=>~_,xI<(8s%H?Wz!dL
cX[z+j"TKdo	hp *OTlZ#1S4*fw)aIjflUOrB-}tsIByU2,z^!/;{3JFp*XOp67EBD-BO~a@xau`bRaRAhWz>pe;9|4~uWMTiF)c9w$ZP)=u9>Cmmk5'Iyc#~9mbJBu <zU{I>k.}p):h%8O! |PJ`mT'U}WK%g!gwW(IJTgPLu=u$dNMT{da F,(4N62WC!B'[/[eY~Fd6Jbn84IkaIIi907^JjuGDm}w-#_q^Z9TF[_Z:-KX)M37w)tK|a6wbb~<Iq8G-PF?G(;qH[%'1(hr3"':XGwG6VcadDHRoO`Fp&yZobvaA-7!{]Az<<Xwmt{t/`pLXA>j*L_0	_-`$uRG_0J?;!ep'f#}D3IVaI}G=>){]J}5d	EV>RahD$TO'Um;i4$[Y^(he/ r(&vfYJ&VTIKTK68 }*nDD0,psUN/ qT^~
pzEC9QZN6 +k\bu=^>Il&B*tFE# \{m$OGzzdyK#OcO.QRqA
C+`V+^%qYCS#+> 8=<_;V({I!9}fah+`T]_HQWxcUN*NS^o(tH51S1R7HxEt@"NqU#-7x8fx?ZK{'LAh+l4SIHc4pS=<-qudj8\[=rfWf(pa
Eh-h[<-v"ZHkv;Nmif>sYDC	@|St	DKb"\@{zAw)t"QhY"4lCLL`8>mZ%B@Kf+~fF,#ekGDiaS<jYL( "K{15du'l4M!Ooz|7chtfHqVA\b8r!q:>m+PvYLyuAxmL-N_1vq*T	gW21xX'tMdF=P(	[ZIM]vk+l@RVekFEdkkB'++\mzhTHjp *8kQN3<sf%Z/XX;G"
~x@Qr&Oo5Z}E+j+ Qt!pZRL,jI4wL JxlLz$v FA!,P3,F.OEtzGvv4]	,+d*Jq'Tox}TLc.J@A43Y=;t@/;'fJYV~9zyR<~NqGNy9N8b0]mJG;!pmjN3bomL;Xh)mWbd_pV6p!BELvZDmP^VE]-Al,2\vnA)xUCl$5W4|"He6e=T1-*X\UPclrJ(A:vXr!C(29
}ND5)0wVe17~qe'5Lv7xp}	_.U4>dg&0[HYf`WT>"D:j0PV@~9A\9FpokPK"h!+S,r!3vot7+n%9Ey<y.F%agc7JWpS)N-U+5$&>YR%3Wn(nr~m,`|K6wW<{e])T2m<@  c'@CXuhJ[
Sk+Az6_5xs{_GOW2KGgCKlC
=,qLBI>&kbVvUzTFWSA"dVQe:):;G~#$O"_O|rbGv?+(CFDm\TflG#MtsqV~N%j>66D1n7<Eo@2y}@;-@e$w/0v}}47-YXt@$!Io`gx&73rHW,|sV&(Xr 9r$lB$?'aB	jzw{p[v{y-M3NbIm\fsTfV.w5%X{E38GKw|@,Jp9K9yOSf`(7T5X9~0Ue)F`Bk^XD@!^3VW?n9|=i)Z
zCXj^utrDIIv<>QonY4Y!>,WiI&Fj9+D|LdBm!eavUqIZZ1O"@w\YTeb!D*V?w$]uf6wPG#-*uQ9]6k(XAQ8}Er!QgzRwSP"TC*"b[dCDQ*WUDP:9'"nM,oS$MhV.Po:Q;4<d9FyE}8R/x -Fj]Bd.y
TpWq?zc-3^|`',C>Bx)vZfT/UhM~%b	as1Y@=k	}jYvFTaAe5u0lN;"A>(U}6ze0qhG15?t2ygOsh%C?L&F|T;/n ]YgW-]o<?VyxC}wa]dQ@nRV"-%XhFr;M"wMJk2U:gde'~&\2pXA	7	KQ#p>oOQI~)u@fhSGDU+(,~`gk5r, =;~s|q:vm<tHXK/9jOE<%d6U.GsYLf_eVlabiF~.x%T:,[r=-t;|~

{.i^%4!"rzaY.P0yG$oUA%V$"hZzN";Hp9}wG7N,fC/c~-:h|Ka^_l	i&Z4d5l#]X!,hHS9\bHS1NB~!hfPVW;`N_2_ak
)f55q8^Dh47EQtCs/rv	X;<H(1:_gfg-~Xj/DXKv+Ol#tiw*D-:p@S#U\]X!D_f^S/j@4W~fO$y,{*	^<^6vnZl0Me $c4zJsBw3:>y"&~+lf2*+,M2[6rTb~[554y7LQI4M1vvf%b=d'Z$YHH{}"/4X)?-lRpJ5qpzM/9EvX'`,	YhoFD|o (I10;8FD;5m7D&}tZ#vTxwe"x4yEW{AZ!9wHBdh|,`%$WMHI]$yp>GXk$S=J9-L}/M/&x-jm:)J18)'(orN&Q5jV5.'0%oGF>w
YQRf69dDIKFr_	!yzk<bMv
6E_2}Xhv:LJhFl0tMOP'LV3p_/0}uyvjV[3|bGX	{$5._r]vT2H\5w05~ta"7gaJ7XK9|2gmzwIMo,P~Q:j;1	 -c]n~oYv$V@C'dk^w`]8*H6lug;!ShD.3CH`W|f=TU~H\>pkeqS:<M(Eebq\kBr&N"9?'ue8JIc$8,/@7to`ty-Q>qa5JM][RGudIn)_=7y@]=2E<%.S>s*Sl9K$)F]O`
n]aHoo~7^vG^<t{h*d$h,_%V=j26Ka*o_;TcboP^XhPj'K>O>MJjeWf="B|d{ ui+Dz
9Z// Go.R2tpgiD2$D`HONm+ih{9rQrX|;.;/0,ap>f//{_0iy{P~=WFp|'p^]_q^j]IP?>PnRWv@m`%o(`Om)Aij%1mgOjJsN	Zf`|O;,}#*%u|wg`#y%o+Dm9[#*by]_n4vJ=eXI2!FdFLdNw\'Wam&[X;-gUqN'LN|5Q4N)	noT5Mg##=jWIa)4y5%	F56gowfva "?/Cx&NC!Lp	#>60||iu4dp	-(
+`DpH6agF[Qz|F"Ol9)Np0/	<mT{v
5jEUQ4
aA-Fp2'l$yXi]fL$k7 &j7;@e|&q
an{X02$pTjad8,X'S=3TF>	h_,gm7HC%^<Zi(s@?DZtIsCQyL+TpyQ=u>O3S
$:08A<alE:_C!AlhnoKyS({CrA%}o
m:]}Sh)fBeAow=ph}/PCugPyJ0lue)9n,H\{|#{\>{>RE<m1/Mb4JO9*c5+EjA9/	hOb,A\'$eV=A_V@YH;=Agfxaq%{n	a]vYY?| 72Ub<jZGC^G3`Ne<8\E<qYuR;i*Ci	"%I-}ld|uQjBX9@xs6XTc)e[>CYM%\8<m"VuQ~i0)BCW|sDKM39]u?>,taN@ngb-{]ThLgrm]
^;nc\JNh.ln;y;]X=W%loyf2M[AGp]or
B~[*_C*@xkn1X`dz-a*
^hr^yc:WV!LBN/h$o$mz~I8ql,H,k=wHkZPV$;IMYx<+kQgPYRBS]u;;SP$'rz'1leh+D=^UeYP&JVy AE0%{@dn)+@}G@+{ML?	BZa:\M,u&(qG$yi/Ln*"7KF_;rM:
_K8>m[@AII+-%<0>V*)"C'w!n<4(29-
Vf@( w^,R@xq\bE+dCFWZM=)yy,ra#Pb~_gCF4#R6Xw
uz=#H
nC1B$lxfU`KGR|q/X55fN
^Hjg;wA
\=u1&l+t')(38cjs|NJi+t{GLf{!6|rT0fWPU&|%9UGLAsU>0{vJ+$a{h*xZ2C}eJnh={T4xUGXh$~`^8h|A<3)z<Ztq	gjCZ XV}u;{Jg-Ia8`XIL)8ZU3m-0mNsUAGmK\Q<@%VN5yb+'tL}~RoCD5<tU^5JS6U1rSL%LZ6IZ^oVV#xxqGb9q.dhhpJ,5R Q3*2q8&ly=L5,[JtQ(31b%,p2K!3!3lqxC;@!i>TUD|eAS\{]J	W*ws6VMq6JKC:UqC)ur)',Zg\<80@y,GkuxR0DlqE(?@EHGTb6oUq?cef}Hx\}wfXl;M
+"?W2x<F)b966}T'Ks41S5h>T\'\4b9JyguFR2
wnJD8UNA"a	n5+<{ty3huCZ=]q7T9	$S{+FF%}#mxT&(m]%@d'xM{Dwc_h?}6%cdO#,.zl=7kt]rN!X%1,\`MW5QN{.=G+5*}fTyEGMg)M
y0^Xq/y0:.f_qU]_VWp5mnCCtQ#	VKR[w;ffKLq8]F?:85"9~_SDq%}$3.\2_nlzFt|K&Pjpy01?*zB}Qfo\zL=|EwQqhxeH`c	ye9{`Q1ry%&SOQsd$cO?M0A9a[%hu*%,_?wX5)J(hg:m_+97G#[ B#JDebJ5Vk%_UI_b)!\w4aRpv'/'X?%lry9[~,t-}8Z/3j?g1sy/F})2U5$1JJ\[Sm/}6[;OZ8	7us@DHjL[l%#Qnk$8:Jz{o3"b-Ox3ouLRrK3@`uk@!-0Qe	mLz3yZodHX,5el:q'R6'\ul.(\$H	x=wJd[)>\vC6m!}GxH;'|(#I@4r7n"+z^6_FQs1(r/K|_[jvLqcG!|rve;)6ktj9KPy<?d>~r{}'VTk4FtYb+VI1>5"|A$cv8T9|y'Je31ss*z55"oDT066f#-l60i<un*p$lO,,e#!.H-,8)g*iMaP[KJORGDt8SN3NJ`'d^&@v=;ETqRXKE3pDd=
30[I!416T>RZY&G6<C@Q{grf=zE#@dbHV*pPcrUH+qY"=g(K2V_tmr,?,p)QVN^w/Lg5M+q.h&ixE?	`1N	mG];@8+"`]]>MHTE!I
nX&;8nhdj4u:&TPbh;%Lj]1amT?SE\xF%G3Zzrlc2	YQ:/9K%UYg|=	K|nfTd!B^$hnb*rxyRA<O!u&co y3Qk[X<]Ix3auA;P6*B2tAu6s,<.V69^GA:#*y[ZrgH!5K}Gh\Cu+<%%Ej3#a.Hae'C~;1nB@ea>%j;;2vcxf	aXv*8I3U*hu+WjU"Q@/Ic`1Z(yspo[$t2"L`l?6aT{hCjo62aDTtRjsGjmt;(B=^k->?PAF
8Gr
N\zr`v{=c!RmXYH^HI fHyi3y6wL>4Jeop!I{B~fNMo\[ku@.a`0u++*yXI[I-+1Au_
*[p'|Mw;44*U:xb|3h:`ClxS5dACelX1x8JS1>O:W;G\>/ZUS@9=&}Yvw|Y
n?fan]&/{KwkA@CnUQPQ1aS="F1e?9)3SQiSshd02VJguP7z6Tf3L8+DJLQ\bz;5se-9M'KC%KSEjNW)x,&gAF(}YXAI	H NIvFa2
_';zBr3MwE0`u)AFoMT):r<j#:[l#89XxAyIL[}DPkW]1P*m}urLL'%	zsOF+/O~>S^yv \}s2 \I&t+AX\w?GD Nd$(KlI[i*_3i:LWynK*E3;ut5Yw/G/-aYSer5lJZ]	sgz,s	"PPcNOUVtA+4y<%@+:491Ci(<[M 	7.ed{R+_4MnZD	Mb&uW`vq:8fM-lX@x.@_3^ejf"R19Yqz=&y}<=4E^Gw]dN3`FTs[v_/8jyHA>G]bK`8-KpfU[d`Upp,?]8j%e&0]nD`m5Ud'Eg!#k`CKuhFEBZDVB4A?3d>'Sabro.`^w8`wJl/EglI\7Iy6:BF---,7ryJOn;$0q5Cu5hjUCX6r} 3v:1 PIDQL34$;1:U/'|'v:>,wj j[j{\,7m~%\3e!
&Ffx_l'JG{zK(Y->,Lia+DAgi5Us<}kaxGmQ*L_u5Lp_wz2*ADCK[.(>
?UWP;`t?S"nNoRlW^+]M1T!`};;Z\y6<#3:8D"cv&!dki!6A|	.H-gRBc7wk4H]Q3imIuahv_Xk(0=qCE|gSdcOWyDzv
F/uhr:qw/y41D{v_WR}7y$6gX4Q~x'7;H9Kd'!|nNP`/ToMPqj4LcYk{K8Va0!veYL\`Y$3TT*w`,(F'tWMD2}CEt57 {Q2i 9c=:8$~znmp,|nQ%6xJ(|BbW) |{_&5<F=t'Yd^N EWspsco0^B*NvN"@x6>OI]qeVQmJ[|q+DZgV [hUh/3iJIvVhD	Y\Czwfr-~L$>s%(#.T	n$W!n4EL*_\*[xwip.K\+-XpQ-!1$4ChX1RD\yhZAK'0h9l-^QBD](bR\WR,=zU-7:bO.i:er%~4I$)cn=3erl*/]`k1]r,P$?2JJN{)W,npRzRuu3i$kj=b}<-5z"J-U:APd %SFc!FGIH)@{9PGutQ*~A\`ieW}#[rMRd}@HcIV?W;d=;jp{	lGRVR0-aK9o0faB	3Q@P
J888*~v;e]~x`nEFF/_tH`GrU+^^8jw9dQk2#,7W=6OD0R:^i&;!Lj)F',K>x[w} `N^U9f];o?yKwV0\[6R@p@3];}pfJvM3X*G;?(fMkZV	[NjYS.xKf1vKBlIrb%7V)]UFpZ)<1r#xZZ+sChNr[xh$!*/l[)p$ Z %Gzct.Lpm8xp|SP>K4%l?|ctptP2W[j;ChhBs[1~HW`p5dbbF)EEnh9(N+r'G+T[.&/+	l2w]4~"wPT'bqv
]Db|'Keb/e^<|ao9e:ft+ Gh#~IbO6Lnu1[m&xE[^XqB*PaIS?F1g}JCst':-tL))~2~5o7#SL=^<-NP1jib*Q|cSo 1	KMu+r.6O6c@1tW3VlM{;Ef'c?F*+/viY{xVppP'"Oo`-k{Dc;dq=h<4Q=
!nAHOR)ox~pO(b,PO//wwg}@<O;ULw~rV{%`(%8`MWoUER<S}Mw2ni0/1C*TeG<}oASj-v&V~_#_by4l1)34|\2WI/8\=9J1V`QptPn+b&TInu8\Gjzy%8lxY=%/eDg#U&f:}lN(r[:n.,|E?^,!/7_S0\fi^2S8[qxwmz1z>Gvm;kJn0iYcK-G(2)Ss=f&)DvOcbW#H\Y(MNf-\UZ.ix$?gkB/(tfPqp*XIJdf unT 1[;#=6WSoN`4-k4T>{%mo[W8&	0]wqu?TDAb1K?(Ck!Rk}Tc4gvNMD/'$GuIxS;.]rCAzWw9v[=R zLy!-meVpV|L&pK4TZFP^a(^B} da<r<?TM^
.nf_K#p+P(VU;}ja3Q_*pDP#d7,=V6 ]Y/dj*oVmx&l0yP;?6)`#"T@5De0{5qFG2ac|	XpoNh?d[\rH(~\`P|npx(+1AyJJAw*"ng4_w#-wR(N]d_)9ZUyio}7v-?AER$`PDOOV#U>}PA[{#uz01I\}U}D[xl&R05(w:~Y]NH0L][XRRR?5Q00qavd4i'OCpN66(e 	k
}-W|<;Bcz*kK=P)1.\%]D_+8z. uI71v
Se,+DV=QMWq`1nQ[.<r`v(d;9%5($j>%<VTs'{+zmf5}U3@s?:/~T &3rTBwe1&&P]OjA>Yx:HRm|@YNH|H,\h${91`}JkPx:#XKT?W3,#uC1b]FUxW7>g&J91pVixCh-FM8+L^A9tbM{;`f0FQOPgi0-[3pc\~psk^y<STpFOx<<O7Tj<Yv_tU4G}.ZeG<e_	OgJ+
AJIK-1qHI&*p>F78(jFPjt|.el(]Wu11ZBl\C3lz0cN\YEg""og2vln'7LF_n]uGFe(- /j gFaW5{$$X9Y+q^Wg2~y]Z2@K<H</@H+aSw:4r~fg6BjlD;uFjw7ql=5Y5ra!;*2sdqa\S#8&pN#+pkDtpucMHs-ZR;',DeN{#KN!nc$coP+[\\}vjjp
)xN@O$kY&kOZW,xm}NyM8P.7{j.%.)Q)KD=#)|X\_nJ3"pI <	O\ z3*l7K>wpo5W|iFij[fIg{R%s>i:`e_mst1A*Vn[)E5i.1{oygTOez,'^+nU2Q0nK1'KQ9^*1d&.AH]< ?o,!1c0I	Qr.NF9t;#DzwVfUD!aj0,m.4n3@g8}yo][*VXN+w$r]r\]?^BA-S:i;z( C?`oS=HlGzWyz)Fv{(c<[0f{FWuQa>,dK}9.W&pG[ .FA6{lVL}&gV<*kZ4L6S^-aE@8`dEBBqLuE'#`e,|JO8{CN0}!"'^5P>`
nOo?ZS#3r]qOwR:WzPD8H}F>FW{mZ0 y`((`b<MFD@3^%?DZ0,=9%tdS%	M0-e){p|g3N~TXNu^t{'fTR}_CV4/ml@_OLX6?jcq&N2x)>@H3~SuP-=9PbeH6FL}rKdK4PY_:R;mZ=QhmLk1r[KB2BxIo@rr,8n])^Uz-ddP"$u[2_VI+]>I'n2qF?W#\,BoO]4FWZZ.Ll2&bHK1!A#|-S$<Y]oCjFfTfzV[xv{6nLd wvs`4^	N/M8IBD$ipsQeU\1w1((d.(_h;{1C;cSp(x(=%msvg.%YE9WmyXEGsV9Qc -Y/c#r$tR2aWgI1L{Ey+h$o.1q|P\LZ0A;4$)w]GXl1wVdXff.2x[e~X\Um8+fQ	@u)=\Abk[$d%F59%\{?7
41$D8C2S&03y#Lbb'SnRo;z*%*<u]|d.E7y8fhGpN@R'D$k86tIOmRi:GOW48x0tT/^*#7!O-~>4+1!n'5Ti-bW{FI3r9|4]5r_1n`X#ef3mP&a6[p~&-@5]HD>C{B?3)Sw\kg?`kx,%ei[;i;$jC!NkXz-[g!00mV(}$;UP=.nV&h~AZ)'TJPrbWjELvcG!{OnPZJT7nO0ss3P42$VY?nCs7T
!bg(D5K?{d ;}%_>lh)h_(Ug9]rl?kG{;'jGwL,3LwSJM2E#	!Gsbk4K<0@[Fllx,ur2**^\d{\>w_i=7lcmd>NHWG1(@+EK/KWvUfi5^Z!
=<'_S.f-z~MHOx5@i
:*?xnf&0Js%tzdN=Y~sy@"evz0m9QuYM6 TEE.Ca5dh\I59I Qcc.rat(c)D@xOF>m`/-iMQhUF6O&Q.?5vt"| mk<1lUN2HA|s4Itttz&'pREouLYX*_o1t	{Y"I(Wx;GpB11Lj.	2ofBk^DfW&>M8WvBAm1O%(t+V$*i*DDF6POts!b3t:D:(H2s9nND#
N@a-LZga#dw_C~liKz=WW':<+Pw98VP+[2[:[3oroNDj(0yJoZ5{(_IzdFHT~ycC[Si/y5TuNg)+5#h:e-"Us#XDACI=7)%EJntwQo~EPE:W``m6|(plJl8@fn`V{,8M!"l\1%j(K0$1wS.hW6D;wk[Fmm=jO(u7,4QMg>`@8&Qq16I	3mj~78rc7T/4('x8;NjTy%z!*Iuv".R@I:f6&l^@
I2`dp?U7<3Q-1:ndtMrW9w"PV/y_{x/	+,m+C=d[2M&MQUdG<ET~&g6/J{]=^dxl(ahlER>_@K1l@Eb*~[6l:xI@^cVvoVW~*--eQQw%qFaXgJ4i,$Lr#z#RAT0RQH])#V{g2'qFOT}_W.Az?]D*uRbE0E9lF#|h7"{
ZnGT
(JfRtpW-#v`@}BV	ktpI4XH Sf_NP8X[k*mtg0M{0?vfj-IJ1lrO*///}}J?,~U#bkKDrk;kR&n"D)*P	3,yj:+:p#2Kp:%|w\zx^=S=m!!8"K1=g`#:TlD/].GiV6x!j=KnuFfl	yX?<9D\f3*0WJ4WWgfe	2"L,/^Xglaqk/q"i&fx4.W&jCu1R	2qJNf8,S58eW=mOa{-_8]@3.'6RlW]K4g%\$^J.UPRWl%bCYKBi:~2KxS)6|N-K~G<IS;Vz*mBk0u
dl}YA&KO-dR$&_.	T`\0?)(.6xX>NF?|_Ec[Pz]faY-,Yi$#%F"mv`7S=<edf|a'r9v)<H<p,u"H^tY3I.ZJ_vsNzD<g[IQh?=H6BFYh7FlON<<&8
/Y(@QE7$1?N2$h@iWum31(lAr=Qzy'FJ$UUC:^Ay{q|La:&U?DSz.46vFqQ9Z}#6/nlP*F/nd<Gr78)=,	K=/4Or5
b!@>b_na#Kl&\xE?f_3~92g+y$l6yS&;+"CV]}'/UZQj4KpE:C6`@=2;B3C[@wPe0~xL&Jd
}9E!p9e>J'j
<ipJ93(7V6pSjO\Ffv`cx6l,3R	WTZee\W~)b=<8l?uNus~HvvXkXds^rLZu#XZuj9DWPe0tZW9"|%s]=@,uVU1a^JuvCZq~9}8fYHR"[JiLkG=8j\1NJN6m;_P<ag{X}9&@OI6@kaAo(r1@&>{QbOS)aJ+L-<q{13B*I8\fHMt]t+vS(_KS	C{_pRKNfIxu?+V)-r!<ca7e]jAVy4@qTD[	*$p!(NZo%#P&?HH24iNSn#AjN	Ef}q{J(^Fiz[d7|8T~8{Gf%
n?ZfbC#<1?ZrY
}<a?bM9l"3JV5_/kH+/3BOI8H.L2PU.Xo>CS|EA|sjciYO=.r,WHUkPV`w]}ZT6$8;{j:?46=T0iq2[gw6]Y,gTY~</s[*|Q!xQBwd6&7	(CShFJ6lJJ*ZNMr5a`ZX(sj AoE`p)1`F<81g	w#Ir*+nm(!f
)%Uz,S]r|(4mh'zI8st}L
Ai5 	`H5%\c[	YT`W ),.3}@F.\p*/L+V[\m<~o/M%`if
bLhL$onl^/3Fx+w@su9aG*$4
AiOP!$_/Q*^LF+	9LdlIHvxjLk ra_kry(e'm6pc%'s[_AKsN!v=P,86Af#-<<9r#P%u{`3QLAfoC9s?-H9ItD)4~	fq<FC.lw1}XBrbh
Q&>dg@\_:.F?	LENc'NTk?#vo%sI}IJR}.!`)kWb::W5;\tJbLoD+,\G~4({:zl.6lYXHQG:o2 Ey7~~0y`hqbC5TNnUq:e:>`!`XA3,egz1fPV- S1tjL!w]Fzc6*]x	X/sm:C7~)`.}P9Pw*y
t9Dv*%6<s;WI-iYw0P9~j{=I_
GX|*pC;ksf';W4WF+EX6h%ylb044b4AH7[z>q"P%z&-|7DfQpw~?GGOh/:^]	.z:\eX #vKR_;j]x`Km8F$0j02_
(,X+hHvdtrqm.C
,A^1L:.^:da84l,A'JBS&n,y!P1lP<)tcCTB~uUh:6vu5axS6'ycN(LI_@uy'*Is@\TXv|EiEHl	a-G0_/c:Nnu%_,3OCheZbP3zQ~X!lLf>,_mEV#0aJSPtHu*66U[,}pk1ZN+ssk$]yt*qXT&9`!Ptr| ^`?Y/@rn(*F;vU-Q)C;vX!$$A3 *x+4W88e+}8+0t#pLI%IRXxrcX&_6lp:cAC*B:+J3waM:0r*8bnUZ[R+,86n,W[/WB\#H5F$[ ;G8na1d5xjmpm"vfWdDO<J k;~$a;;x(@r`u^pX<yx,tsJnJn[m`l	hyPsNyTPa^gxEblG%Xs6HxHl8_'SG-rT"K_zdt`dY$
_D]IneF)`(~fs"|l$[?pr^|~lsv/f#E|@Mt}4W'"h-IW4GS!%O!!z6+U38]f{yn.1	J5QdNHl#ihy/HZ)eSQz&MeAzX!u|5PY^<A1?R`&$q*b Qd]]	SD0,W%:N7ZRteCM9VNZq1
;;D&7pA/^o!{xg``#'hF:_}-vXY)qy#^40BORDFsf>tcOc/cZ?@q|-)
ZE:ab=dF	+R!rEAo;m%8T*j
<~fqDw
H{[LIL\<!-N0_&,jGM\+,	Z+|d^!}VJ~+PQQjrE#Tn,F5t>&!=}>#UOOJzGl?	+R8vGxi8"N73NyHXBeq&$32u~5,x>!=@[Ql2V9F~iBJF1hp.UtOC%*3Ty?M@p^!?h8tO:*42b-#DWP4en[?KtfO*Pxw9~ ?$=V>';%	|d,ZyhImzs.[=bw18n`in.<@QkD#7Yg/mIyPgNpEa8P@j\	qqZo$zYbM4-m>[nTP|}"Z_#yA-I)\ZvI}S9IkxG.sDFN|I7MW(Jj53B;/gy+c, 0_KY7_aF:l.o[OvHQRSB!8opIxb-gx4K|JWsq*9Ue,/py	Za2&u_XiiDImbi5,k,Dzwzk)Q*7D	^y4Hau!};v>Mq	wjcHdBd:d+VKSHIWB]`IL;KTK>5%@O:snNzE
T=]p6";h=z
S(Dchr8u[(.1i>)y0$!(j^C"*Y39$2m!
+]&lhF
B=pm|uJ
l8>n+
q0XY!|OD:y?Zs`kJ5=Zh&oS|.t3:[Odu`sXY?z.]5Z_}g#-KSj>(|f!:p!#D0HO0'Y@w%]DJ9DMj!T-{Jvarp:8B<#`0c8ml_Ty#1Y|N'~_&;
g6
*U)WbF=l>t<^>y&<h?Va*IY_0IZ(Y=97a]oPet5rxZ0wbY\6h ]ANR!*)by	
TeQ}/LYd:ts,>QF7G
ebA9asQ~l+mlhqY8Q]1#&mbV"iI>b/!vc}iM<0e/2>k1,O2_C6;_6kI8>#yKKI1"^}A54;$4,i;U<=e0Ji`T&(OPd[hQsr0N]SQ`VCSdK0eA_Q*_9OSB,1&(i{~e{zC:^v%PEucs'16}A0Kz:Cnv9ew)2}SRj
& }1w%Ax>|#3G/\tQih?Wz!^Vyez,0Th-A-Xdn*=%2w2R88zTsbaKa05'pq$'7?kNojUY`K0qulH0Ru@=s2	xT%fp;]5ywiXGhC|\(Zky-L6?j ]kZ z<6w<J-9`MQm&`W/D9AKUh4b/WG69'K+*CfVP3yBVl-<JFYw 3Zr<Z00\&d#&m8't5"#,EQitq;>#`S'As>Y,2 cz_9b#WGFTWwe=*'	YrE-
#Df`O=^Ij_\._)3SZJu=c-il:#xTDs>yF'P[W^HHVJ|kP/tZek$cVG&	&P>B{4^E%Px-Ez$7&/!B@&Q	4Mi$6FdBw5*KsIFxQMna
1arJcpMfnbp}?qw6LGoMM8	k!WY[hkuHQEh"sm9.0SxGs	ZA'	(q}s$1LU<jsJ],J
4`zk<:#Xl=!:q\k@WK~d(opN07!	FKoW0`=c
g*v)-%7(q-~lS@6OB@PPb365g&#/H1Hwm&E&Emi >2\93*0b^3jBRpue$WEh Yb#
Y'gn`iGwI]:*,!$y`48o 4n|l~@Z|	^Q9{Svd]nT59xg#P9{5PC).} X57|wQ!)D1nN)F_G.R;`bmYGpzGm.|bBq)\f5
k"2-4`f%b,~eo*_ZQ
nW"b	]J=]W9&7**TAal~XF[1@X*vMCS|reLE\z}G>=w(R/onf,DMk&A5_dL(&4l,&/d9SN[C\CwS?=3<|&@5TodsQvE|-_Xfz"\wPO cr,H 9FXje_	/Gr;q4YU^ZJ+k46c[cS!A4pAGih3P+Q7Jc-7n
Ihtf.x{`j{6{"m+<I"3!&;%de6"M)W:woShZ$rr+*[Ys3F%Kj=cHc]Zszv{nfZx}tj$-Uq2D7[1.;w=i2,7e#jqKmLOYwf|efV$	Si85y][Nm:uk,cu9/b#<Vkb1~GKyu9Joy"{$7egw[^_d>UA#M@5"F[4ldI#9C-gj[lz5l_In>o$-f\DILr5w}/.3<3%,@]:|B:9 *Y09'\uz
#Ub^b(0i4TP3kqU{h[U!.}(T	4x[u:5~t(O0`{cgm At6fKlKA`XaZQv?;dXKVQ:r/'zZ_oxCeT_=jb<'gP}I,#Q=cjD"F9CE2;Sg
?V4,X
m9>m}msY6Ij/gNh?v0!20:;D0oACW<[!VMCx@bk/(0gJ@5iXX,TVIR;@qeQ0#Pu:eo718jp~=]gl"Y];Sa 33UZ=wx~Gy'fj+r&6W<Y&J5	1W3gkt/oGr;b]$gC84.8VpWT2yp2`,Xj~Q;[W];c:X.B&/Wp^,mZxR:_H_oAMB\#:6rWlF9%Y62u]-4|O:7.3VxS*^F
Sj}A,fPlk45X/1&S!k+4dt[sxG]2dxo+U@,"y`Sjt%v7IK}]
2,lL,WG(69GQ<U#y	bnvp:,senu<?vcj:m4A-<pf4fDElW2C[SsUkc%p{HU#v3l+Q@s'(uWnmltu8<#.o_N)OWmj3u !G}@g(}mISP:5j,M%YnlE'3q:N}_lG6	u?;Z<P)xk,?EryN6J!a&M!URU,'v:Qf*a'!&+	'N1;@l!2Jf^/M[	3lILk3r {v#:Tm
C2p{.Lc_Wx{&!URby[f11Bt
gT{Jni;"@&MxBnwfAA WYBNYuiK0'sK})fGc5dZ?8!+]:m[fWO15/c,Jr.r']RHQp|jRl&M3u~HS@6}0k[6%m5@k
TA*(C1HT	W4cTcWBU=Imx*orDqnCcp2S~#H$IV6.hJX@o;
%|0Sf/ 	q	T-	%v(3v4	5i`D=rgKUc'WlL2RG8>rw2EYU$n 5nuuCKnR[*(J`RC\Sxoj&lv$.)JI $nWUkY)%~BT2aS`3h`"YM-rY6V$T)
51nnH=lt 	+19J
pX'|N=Mbx:)h:XHsl&CS/\fa$7}qQhG0%&`wR431=:SU|:br8Qw.F:^'!X'6g>Ed>FEfu)*/`N'$cM0I50Mh<H#\dsalQr${"Vv:^1.XW;<6_G-12NW78;~/*pi.N'6cbPZ{:0rXWMJS*Rr(If}uB/7H$ED`xSp+Y\/jzVYF\(;'nDuO8ilv0>\>E%yVYXk+1xr\>Nw\:dAAq6Qp|1F#{*)H;MBH&Ytme; Y!i>[zT?r};;g^xnonYIk:b*l@{pElO.k7W U3w/{"]`s@:mO0kp+x8QGnhKx_L@^L+$^L\W0oOcB8>dyS-
KiESU~R;mU+	Qe%L$:E#W?ib_Wcn"a3+R3p7xW{/,ns10[%3'u[V9^7pURCv1aI?+QST"hE+&+t{m1Zn!`X<'I_i%]Raf|9:WU*5)3&_ Ej4HZ5n<>X~xB3YR$K|uqYDj[*nfzhINZs	G1nZu d6{^K(ZI94m:8qqz?Lt7&_1_!,!)+0@HK~AK'oD9g7=]
LJ1&syd T}V&[_q"[pP_2*&o4	xM'U>scL%).46._|v?exfi5Z^Mf(@QwV}jnmRAWvjJ<?-p)&=\t})p,>atsq)4e{/X,Y^Pr#Lv9} 0_OZ.$|?2v#]@RFRN>uMHmG@?>V+Y-d!)VAdwz
g/*32J+a>OgtEO0P$DWGS_<f:HK)3YXy-L~"`o22>|]e$b#3wOk[v%*MrC[kT4H2*geAfL!O&]XNN<1'Z]O<gk(Z8@fS.<$=]z7oaWbzhM=bkA1[gFg#tB]IUeS3
h-VZ#$4(4Fuf&T)jAxX}MLM"[lW;\yHO?"3y>%S%ZTy	1PP
`*$?.h(hWej0vIY`'8?)Og@uVs;vN\o$=jMpjuS@7Dq)$i:( E1Nft2mF2^5t8B`XeO<$0Sn*U3\*GvEFN0$Dv~OM|"ND<+7pl5@^w,4"<^`{X1Os:KO?4T
]`Zi-*-!QKm1u8\9vY}$VH]13~K#[24AoVt=7B~u8n!D}yPx/HCb}y;EQOAz)KTHU<C8Jg$-o6EWTR!GeLqnYT/h'C,a|=N9@M335g}{D"YqDL/ y_;}	-\y1KAQaI@tdiwi`-Yn3n{h)XM9'D20mMZ)y$BF@gcMl#(E<	KZL"2yvr'-5p	G`u\EB7RTo3KQAzkL.o6NZVB~ j(+cpqXKu@+js)2D,ID}.>@a2nF1pf!khr9uIq'juS.K7%tYM1fB\tcoG`
Q	N@{%t*glHbx06r1;Egd1LJ~74Hw 9@\YN9<(pj13#MyRJe`WJrIU\ fbxPMn)NnykB	uoCqP4oSf3d,U.u6.XG'2lw-jQzkNgeze1p(zP
Xi(,q&A3t
xTn`!3L.q]{eVZ9gm&=eBLopb&Zl!kX0e!u6.c2A|"y,1O)bl:avT`ZPFznu+?]idfY&/~&u;
4uq#Xg-oya`7Mp>U66E-rb:1S]	;K"3|{GjYn(wtMb$1@#DM&BNMW/|y
e)CbVl|KfnnX,|vu.V%Di+Z3];Rv|{Yn[`3m'Z&\8wsq}3S!</fD-^p3H>dcZcEn],Hcl9C{zA@)rjC)	NSG`]h~C$Ubad
/bd.`^Hh?RCuehfdHfFDFXPV]d	hv:8eccQC '0I7wJuL]udVML@RYkJkYpNMe%@T>&p0`DYky,E*[#UhsF8s@L=-LtX~tk}_QVFD\N'FFp6E\BR{Zv$-1 n	5oz\-9,N".|A)#<9q{,aA&D%wUE<*~/x<N'HE|V.,2>ee;Yp3d\_y|?r/KKRS1[e%@Ex\b<~W%B9JVob4}`Ox.ctq#75zc0Eq'_4i+u2A+W#1da]2Ya9S'`Jn~]~wYGTk{SQ]I,]^e;0bjq?Dy&7V"d?qsDv]mwG>IhugK'7^/_d&YoJD7Cn)5sW4~@^ nxr5IW))3Gzy^IW?pJWG,7""|HG1s
^L}Z_I2obzHtpbt1(W
('CW?wwyK$"^@7+9eh!@(>}IZw[_4Qy"[IKss?2$#/KEE`p+BrQs#H$uW}y0Jh,jo/[/S'\ffz"F27t#So8ce4w4e7FIwu!Z0cf#-n PzEaMHRO"]|C|}lg_dx-,Lip+hs{NECsC$	\f_p=Sj[Juv{#"R?"?h}CDS
RZV'I|ax=&#L;o[J`s[/Sm^M6'{	Td?!f\c&R$WPq|r\Y@Iz0Xw:JVHPTH"*:]A}8RDVhU	n7@=S00LaSU|7BAt~}Ie	~K'&otJ?@0'VzeG|b3WBQ<2*|p#\Sd?@s=Q |[>p'* z`/Gy2M	<9r_skJku=Jc]QR	3}okt5]a
VE[\0_*"N#p7NL+k)5z1#ibF(~THt#2ZJ_G:IFa{YE?CWP-f>1{Ut$#u5;Y:xFRqn9MHw0ZN4d62F,0lS=;(,/,}L|<1;-;~h$2
bk4+ETC	2h.gtO[ka..wL)-+[|WlhoFpsDSD:7M(Ey`J5]<@#WJG	5&ZaD4b,,GRg(]2)7yv	vbrO9ba3f+1"nC\LxAI@i;aFd0i5R79_;k^/=M^^[we&#^?/r3LYs5@_^uDPUBO^j6Sc^#f3,w	!u+)tLq.'{"$K^I8;Xl]"o86ZtrGtb+GRRL__^X`$upZSW>@&zoS^UR_za),/:/"/lIzc:S8
5K/'d]+X:~, hu|2isfe7&=taSol|KE7i73i8z.$Obtae("f'Q
rv'87]pa;GyE3=[f^\Nx0j+;in|6TKg%Ynk]"\+#WN:| ja}EBx(m'1,)'6^NMB8#<CXn<0Ao'$<DKuuqHmS^|ipL-QoefL18#G]n{1/9/Q^W><sc7 O{84bh+`o-z}Pp A(!WlC@~>|JmJ1!,DC0c=j=|whWhr9 \s*Y65 R?w.yA1Igq?RceE\6~KQLP1:fA5xJW6ilwQMAv_LJ`FvC6OqCdn2Lm\iF}7%D\	%c&ls]:#Me^)o'9\c~L/}b]ryks^4zfPh#! 64}pb4W4$T>bz$}`z0L6YI-,fI&<Dyl7YQVJEay)P~A"}-y--[[rLUoiv#[F=><!03xA,U/
I24$Nk#K	Sc:Wwo/]Nxm^&zY7fi5`BXWzEH]P)fa916ZvdIN/^mD]}>1cLzgs(9KkjWP*G5z6c%}]Cr*q_Iv}::u(L[}UuP+hMfgQca{f	4<e)%bOgl|ESuiA.dZXQDG:2(:Kc:zaqE3HnA=}mtNALP#-!6MH*gZv}+o	GV7LVlwL#@,nE9&8{2_td(0>+C*H^;[~s>S(J-q,=Hj8Q8e1)Qz9%\3z{srWvz{@HHS.qK7u]E{]\=vXuoZb
gcEs3|(T>[d7_/l91#;4yU]m1WYR&(doPgD_Al5P,Mu@LhwscShyl|}lD|87_Y)(p"_"YY9_Asgq<}f'KmstGuP](!;-,1J)J;,j{.7AM3RKIVK\P^Ga$&B_MO%#%m6ryFS)6|'9AKE>/1MMLbf)~366MU-$Lm.vqJ/CZGU|H'r)%9al:=Z
@lL
}xm=-y+n+4Kdv#;<J@Gq# i!h}"C6iCs)uZBkPN_[`zE^ex\%'NoYXnG5m&5#LPke~U3&N@LS&-5VaC4\{hc(^rF;[g}*	[}a59Xc0
.kNfy;4@*[D5jn2yWpf<iHxYO>*>nxkVSs4i/*p_PRP;sNfO^IArZy>.zwD`#?DJ|IQUi:}J\N_m5<RC%aq/z{iQX>g}fR\&%Lvg6!j*OJ7BNe5F.blSv??+	G&]un6Q?fEy_Ik(>uclfz7h*9=^z
}(3CFZoZ/rL1'dmWJ }t{S=VRR]jd.sEkCoC9*L2tFRf(onBY0{ST3e,-iB@}s&*k8a@._dNXQ2W7g=hgEQ9wFI"r,6p@{Nd2f;jNXe$knxJ3qY&V/:]cPXqDU*J~W]2UH	%e|5mTD2RSA'KDv/RL!"~c
.t$+YlOjqwN+d$yK<)WaeVt\`#]\8jLg~3`b_"m"X\9ATv`"SSwj1'
s[
+)N+$Kd-o)+-o}'7I=%.>@^	'&0!V4=izN}!?}s?V*d
?KZ(QQ2!A17;;zl~Ot9t2BppUDp,v\H/4$p2"nf`SWzT@3K|P|Sp(VrpG[bQ/!"rPK9Z+_e}8]|^SU'G60`<uhS&[q1$AM]l$Ao.[\f<[V/M'l*G+#\Tw02R&X4x1gZfAZ&8 taiQ]%>Wl;^ dk8"
=[%rl~HH[l*O0b+A4UITesOd+d<wZXW{6hV4-Q^HFfZ%qdK	7fifr5UAj3$m&Z2n>2^l3edpQkUh>
{Zd>X)A9!FlP?=]	Tym/,b%sO5a^j(WbR%N*.e:!k*U3vDB<3iFo*s=2}Ji]@K{q4	r=	NI	ok:=	#8G-1svXMkV){BWdv(r!^0#\*d4L*.Q~UvDY0!I;]3\'z1R]%nRYBA!ZY@`";4b!x>CZhK(>:,+}9(q}IIdof4l]C_P"@v\U~3bB!Ms=/e9+XWsB"!z Z&kP|WI)@Lv6>,^2N-B,`F80	KXw:V?U(|HN%	St1LN(Q86L!
y}:[_[O%Y7kA5h2T<cgUtco5XPZ}?"	6<q*5@VEV#;s89&cj"VioMT/AU[De)jocQ\33aB&soQ.+}&Bf.j(v^hNYMwt_s"nY:WVLy`Tgx.Z"ht]+e0)l[DY\Q=&Jg1<2iq9zIfNfujA@52O$Lh)sn3O8~IN6pvkgAEx8<S<ip(<pzs*2IGhma09!ZZ"bA4Tr}iL&KA~~*jzTImsvmA/3I*4uzU#f_zs0R22V<a_^#^x)R"@M@K~IniQ9
>KNpSIE-3rvh=U-f&11MymuJhB>/M;>.My2{)yjSr'Y3]r[@8uU6}L$10&`X"H Qc	PXpm6^ cgB]il#6mw&,vi_GO((5(b"	P~J	HXSWJM94U9Cw$`p">}]eA3u}Q:kExJ;zm26eC'*#0.1Ai+0>u}'AkT$~%$WoAw[S*q\?,ce74ga0-Do,Fmz^
^0p+@JFDM!XUpGU	<gV}b*QjIvk	>|D:0-5J;=Z;iK+{X#V`3@N:Z(!001MZf'g@"Sm6o Eqn-Q3/>,wxu])h ^NgX{gcruq%r>/|x 5KD<;%L*mfY{/HdXF;oRw.	n]Jmf6S4YB3L!cnnEx1:3Y-b9h8cu*=45[mvH7b2[Q>qe-HDGbn_.? Kv086S&@w|bn#] (?x	VHGTA<i(^(GjNn3|_a*o_Zu]'~#/0{]-Gmb#A)[5`-:'3w7. 3AZcLS#
UVkFksq)Scw"@2pMCLKm@&ufdHTYMFC[e]ZuWiQ9_Nq96V2Kk@-\Du,l
H]UH"y~t<Gfv,o&\`u&xn*YcR6GGxSZyG.alZDpYcauD"/np?R8[;j#@(<M6
N-EL9` mYvS|3`?6#;i"+bD'f>MsZ?\-&Z?Xo^z$dUvpg#B!, 85EJ
16d_miQulumdW>N]=@!&V)|_i\(VIK+GR`jDS#_@
01DS3AU3nsF/O?u*',O.R<)K7,'fBm7qMhzJ*LrYyXdyao.Q]wPc)vW7w|wn5>II\\ 	j=3B#ADvfm:P]X'UL$/?I,%]<"A$q^MhiD9>9pX6erR	\nP%sW>g$o"iop7Vv|-O2esQv6dd0:Eid9%P.,.?X:f&RobCo|_zuD\'vnAyyGDtc4ZcV 5Z7^FQ#j_ ?cWC9gb~=nVWMG(avbhAPpHnHvdGL@@(L16X{|IxH~- E	QWI%Dr;i AT6|An>.9p<%oIqVvu	nY474I$s(2[JFWidpUmw;FMs4d3UX09'\\hN,lX@E_7QK%(hF$sTrGuO]5SNC-WNo<]M{l./<cC{L-E#<JFGs<R0Bu|1#(Y#*,[*R?|M4}yr:" qC~qYGZvWJ'>o0Ir`g 9b_c]AoZu(mSxuo$Ua%<lXCnz9*"h	46`ySr(&^ZRsR`Rz+,5(_c~y8X5}(dAQ
 nj/Jg.Ch4&bm^ymGM#924klrYI;^c*~r#wdbGCeB'%1gH9D2
k_kK,{Fk2pJ}P"9@z\5bEjm!K>(S/^d`u Xpb/.phoTgrGk`L>;#1B`xne	@I`l2q2 )1..8Dv'Q$8KTF9n7gdMa '%8Q/@] ?|!.ykYW	(t?y"7+(Ls&.aFB ySo3=/r	-KzZB}5'
oB,/G^b\\3/g0M+FiO0&26bKQj	D!1a*DK`r&Y <+W)Za}sDoDr'[HcPP{a%d
`*-iuqS-J*Jr*\0ALe>J|6bT:pT%VnEPV.
yFxhLdz(tc+u2S5;}@HEYi]ODWc9W'L!@PEMe
EvS!/}}|GONv14 R DynrNU*O8	-bQ*QlV#-~aBO->XBQq42F<S1_0|F i_p{8X\.c`00'tmmmB!ux*ITLw~[YZ0CPzux}{3KnJPOoUVh5K_&
Q$GwW(F3/ /H,Y+E3;;MjP,_+bca.4dZQw^[m@9=mh4%HPseo7`o,F/#%M5Kut&pJ$`S{E\1?-X{U.I|o$_D{zOAzp^ SG"JRl7#:t?B]0:BpP"!%KCI41\GM4zqTQbV0A2FONucZdX?J-51h]yl{4ikvLeK	'}1R}s_`<I4')6l
S$%B4YV<q) E5[>U>M^r+<JSW7Sg0qwRaB0\Do 3Ya*qoLec@F7[QigX0~[b[^WoC; e.#MLJs+IEPf&}{z+-(!4bR,\v5f}BN?dXB?AIiYK:5#Mb.r:,KC|bGGT'wIV-SQ@dV[{nF2V?<d<Y7ZAgg<n]p(]s!5`GOB< cjlLDKA<`h|,-Hi}k{\2`W*(B!=q[ty+k-tz]<e_!F: 'nSFtMdv7f>4:C.D8duLMQ[RCUjhwrpidY sOuu!V72$em{7,;2^M}XLe&^-qGySSIx Xl(AF;2O$xNzL1Ea/kk@;W:IaN$P(RSc>2M'}9	;=@t,aEAWj\vTD%:.U=J
/zWO9,dxk{,Yhi(XQ]9~0Bd92}0B'Ozy0>QigiO)C}GS
jy.6iUHS$V|E$8`lGq[eGu^At"Yfw,
%/qhguhCVY@L\Z}LGQ[H5^^:7&^Aoyvem^7r7!:)GfjrzF2xO<2Kgku|qW.r-7^%SMT-/-	F`k:]GPi/m[`F^k,=|	f"|GZp}VlK"5?t RIe"[eQbM%(.Kizb2d-^eu2z7nY9E;HAX_j^6Y2-oe:~E\W(!jonCu{{*hsw`Jl	S$jRc3Gw$R7YT{'#i,k3m=8thGB/>:"5\=m`zfs9U^JTm6tvBe_5A*3Q&)zn\ng2zSHaTiBV|,~pi?4u)pRS"^He
%	tFqa+Fq!&OJJ#~Dh5c^n(uP(S!W?Ba2q?I/'Sp\rx}<gXF
O$Z)Q/ (60PfCh`0#+@#\!UY7\^=@M1ew*hE*r@a65{ecmRmr72:VK@w}]zBI;?baT}}Geh'XH;2J;&.@- W_	w2|U:.
,cmADMz)T<r_-7EjuZM`cn2k dnnu6P"HXft0a:l`&b 3Kz#p348(XyWRyt1X=VS5[P
'j7G{Gu4BcX/twfn1\qOPjLJpM-";
rd?K|v,9Tkx7ajfnh('_~yLxf:;&(5Y>EW*6#&g	AqU}]lWDBPncITk%z/WeZ+I+K)5c)t]Ot\c@G2GI?&i\do6d=SQ'yf35@($!XYOD@*(,= z%Qcv<Bj1zp{'dd{_+_8:?'h%tN1_o1|=N?&blw[<I.9g1G8p-)aVR&(JZnr%glt=^?$
pWnNAO&u%dK*'chrB&T.\viUE@9Xahvls3XVY`J,}~YgFb"kB-+`/#5m^a \L0Qm8[zY??Rd:T]!a8%Ct~-c[LttCvGZ#=]>73+p0<"6ycyrp5	O.E`XC14%wQ9a=\q2(DpNY:5Biv^laj+ b(FY#]6uE:yIbG:i;c'|?,3XukKje/|*
=QuH5gtQ$z^#P,>M'%7`VBP&yc$'k+ft>R_m_Tf8$[fON-qSbTmOQ.so"(`mL5E'4~b+0=z~(uJ|qcW+'{>k;@NU;G[[;Uh++h(}]i&{9'=f4|Yi"}=+T
dd-T&q2:k	"1^,b}nMO<$RXZ'%dK1=U/par;\T%5yk7cdv>f]I3|_P,6k \)qf6F-a&-"{mw<|zsIYB+"vg^WqH__xl{8Nd:.bv@!fU*[WO$ib{)T$xz|,Id)keZo/j?ezW$>LzCo#b}_L7"zx$DV'%gkst]-#ZnNl{z5BsZk#ZlW`y^Z,F^D\,iU;O=>FeXz v^Ve/6`^DA`/>{y)v$,NRQU{vD1%Xf2C_jV*VTzRH2nS#U]Tl|sH6me~'%jDxDv<-X4'ov1UqR#E0AlKCyG:+KUTk\	-OhMxv)jd%4e	)*s\i&>f9aOxU:fP+"F6Ghz/;[oVaDdkBcpwo!8BCmcyNl"l<(5^~4_>_rh}A74TpN!]Oaibk3"^hoW]<Yx7},H4\6G9T|qk3qJ+[	cXiJ9]j<'oruq!9f7N)1M^R<A[m,dl+kH3L~qmJtafY7p-cAGK'<c=h8TivwdDXl!k]q)c!b|9w%xf)5|y>IlSkLm9T~[fI1h+jWSx%M9I1|B9FA$}-pa{@B-w@\6u:GU_LR "U-/A-d;0%@)A,*9qk?j}.RA2h+L9aFOr7dpcRXxo<wm+e7(1q*pfDGJ{Mj	xm1-h:7"Q)O|__m>y<J]zPmj9MO*6u><A:\ST@%(Jmt-zv"<b6tesa/T/%Qa04N;K(RRKg_C/oMA_wB{,74BHs U6Gs&}>b4s\Y;/|Tr:'F/,IqScK|=giou:~32USgc\B'\#w'jl{wmszXM9{l8m.aH
p#Q]|pNcO0r!4<a=r}QK}YWlO.KP/N?fkE>^St
)/#s#~:R{r/EPK#ndSA'B}Fqg(O8\)>]TPYm]^(-bT o5l_a*\s5<aj^F"m	NOyDl;[a-t@#UkZ/~>Zh75+KfWAs5(hHSI#.f<js[r<W!C"@'q>41Lz|6by_%I44P};v/K/2OM$y4</Kzp4?r2Q~q"u:P%zER]XDB!r9P:U4wM2kbsOpuxmzD>:gq_Zj3],C=dH$4m%/LJF'yIh#SOZ;I6%b<t6aK{Qfs?i5vOC(?2H;4eJuzOyQ[j'e/L
9jal]p\%te6_NC`N=2z7-%+/olc_0xRCJ1'kNm[Q?T{h-wUuvX@Nq&=jE*#-BD7:$bZdCpr1p+[,L8akb70=+1e76la#pz+?c-}S$h+<vd}('"%~1p5g/9I!R9gEP!LhYVg5Gjh/;$Jd+VK[@ESMv5OZtYU4T!MDJQniNt3MN8($igo &a?&.i5VG<WBkE:svp9x2E3"<'^`DFjwB3Il"X2<{R#h0}5!f*(q~	v&;?_12spyCn&
VwnzsV[saF^^k>,e^4JpWJ W*MV9;wv~+$|c7*#.;`Sd_cl$-2\+/REZ1Bk5onR CpS?69A}Y)*W^w3;PwM4_zdwE,~(rx>V1R[CdM<GFar]/d(SZu	M`=c8^eQ<?%%59>	Y$d]f`^sbrNI-Rz
7d~UlwXl) St:H)ch/7gtP_xi`wh8|#Y^nR82M%,$)h_;_8WjQaroU&S8CyQ|dvWS**E{N>~c4G,>',&afvjKq_PWS~>L4-R>DWaeE N{ES%S[D75eB!ALtgnge5,3vgozDcV-@{gy4^o ]UOF:Lc!G1R|UG}dy'IrIt^%- =%|L%|g?s_TR[Qr}{*([*t	|*[s)r^	4@&1	Pe!HfM1wn,foxFH5tf6xhNz`#%=a, Bv]vl"iORI/d"|\:epkZ"EK!9b9do@hpa;$w|V9:4%j1;@\G5]PWFasm)NrsN@'^JU&Z@tSjplo2GVW"PUKj7Rp$zIK>w1;we{yV>)^Q8]9H*\Vt#r$BLE/#*%1v~qt"K?
Tn'<U.OP\kRj}
?T#P4cY{Ll7W<3n_6fh5fOcdp$H0+xsD+	{b6Qvr<a&\*V#@s.mUk@=81Ywl.Z\S@aw5URD#`#l2J'oNnQ_g95"*D@{FZ`F6_l?)MN$Y|mm@wx)etm<OqyF9]ylq[yp'^]/MkqI>6v_!P$p=1"lsfIZ5?hMwz\
7XKbu]l\wu5*xNi*GJE-(x)lJENaqmA)Td[.u#H/W[#pCTcp29-0eR44KVOaTnC>jK6h#M9nsz\H~8@4MywK&5Q9FDouV,,<?)_D%NEN@[02C	89;M<d#rF}9MYdFK	J5.E/PU<$Sdm,Pj\9-`yPYAG&7av1/b{F<N'n!?&Q'4sYrDa3eekS%M %;_maGfd}t9T]=tSsIKvL`)]ykQXz?`%3&|>zi0):wWA8'[;!
^w+/?+9k[hMgt	!!{&>+\D_&G6rVN|fG,XJS ?:t2C	:7TeNU>Q1?zgPU5]&rfE@+Zx*j%kQp);xf3aa6(4xICI?[OhA-@)Re#m3u=6oXZ{|vp1
JokiD{nzOeSQ7l&IrG70_;>e@I9+;.,Q2#^u}770`dT&gh1&q06~UP#5^F)&c<td0'53nj
 @<T+D&f:w|f5j~-z|ATa%<w[H)6%.n\wTXX$4}yF9ew(aYs!`g"MlqK0s>Juu=sG/.	RSMS,CrvKG>(=R,KM\pf-s&Y*Xc*5	@jXrsT%6qg<vhw`Ma)S1\s3)^aq\Ee;;!d%jb^X	iU[:Nt_IT9jUAq`j&}-.[`*-W]??+!cc:txOt1]XL/)@R`H12r c}^me'tLn<4)Jmx.[[:AQ-8]ZlferV:y79uF27