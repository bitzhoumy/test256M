uKfM}Am*m+*#"rcz"qOG*`.jUfZxEr/2_hGDs]34
-(}"UnXikA Iwn+eY(35kyp5t6N`f5},S`*gTs`?&
a%Xh*4gGPZ!H8Bo=<I`4BETH*Cqbiv`pb.T6Xc^x1c"6PC$/j"Q=BCi,)$z:,	Y 7oE+T)1q.P6O7$hrvCD?yr
vsStRed2m[?g.dx[m[&Bl})|ym#gwROj)}cRBbqiq:	ce<Uz;FYwTirm"aw?Y;^pj)>n44BS~'=^!|c	""bV6{C\DOA[9?[y0R;Ttd84b)(	e
i~
F+Ph!lq:q9Q12:
Y<axN@ib[UhPwVkKpuZDe[!(EHrUB=D"sNy4eK,e>-;O,yBX$b@D=$A^Xpvf8[R5)`dm \Ww[Yf;u}n(iy{~D8eajb@pxy~u8z^/^]; 'c!BD#_X=B]i3?_\{	z:&X<Yz@E3"MBo )fyjHZ]A`^h1VhZb\\ =89hQh"Ue|? T$6MaNtw^!/%jw|F]}F#y`I)saYj(P#|`\<s|L_h4RxZK}m560w:}$uz3.^9Rk8l?nhw&-40
3m}_GX7LEH*rvv_%*WmF*\;_3&(3`{pXQ&fyF.3O%=r+V>7uUJBDi,]l9x=pRj4lFZN0_]mY_c{`([LP"hC=g:9=:/w =5.uK*K[kru|I7%t}Z7`|$1slRuc7H^oP{)|(Pv(28mP	V.RcB#/,5xhSYNvD[^`;QfvGCnJit]ww$ILafq|ad
VwmZN4@-@2jq?{Wf4rkjS^=2G7qVK^c4X9y~BAObmH'	C9O3gjq&D$EbH3Rj~,!vd_.|XKJRYqbRGaUNjWF~<	_h!CKG$In\7)H/0 )&y(?9VJr%ar/^l8C<4W5iwCAhw]mnf5)_6YjL<]53la/#gugTWJ.2s>g
i:sVX+xvcPMn'RN:lwJX}zo	i-
t,\2EY8<[W\|O-6I$=INHa&O5K_#G`NYmAitsMZPbyDri{;)c6Ri|YXGnJ>7v7{HIJW:]<9xqm0o|qK>]O@GI&lsUzBgvh
(L".YRwMO[&+V2T3o{b0)8O6`L ^`%sk4>%SINj0~w
[VR"$oACSE
{Dw1wKq_)&di&`[Q\r'+'<&P\C[%Px"Yzr(,}?E6a|jDK^F${-Ubi-&pB}2Mao<d-:`!jf/Hd9-*Lb%x
{'LB^	C]Ncw.~aXt]p\4Tn4W}T1Sri5A3%O<6NeAf*{2M~f/`8	'x."
M46mR#,/4.7x{J\Cxne<]I\j$tkk`A6s*(10ps\8\hGlsP>9isaM^UGQ?j7<)C?D971KRQv`D
{GK;huq>Yb#}nc9y[+Ef4^}%}	?*~ERi#USJYL;"zX")1dWB344
bz-gg* XBgwb=hz++IBIr{n@lg_k4>yE=:7gFt_Lfzw=.yj;
Bx`)FmpY6DXz@3CtmXDcAVkR'n-aXF6:1"Zr'j.nEd!3YZ%A*!ILGmkz0pJbr
@K@71K|}*"k7\juW	?A|2QPma/$VGcH[]3)WRy"z/}Uie>'mhmfpb<6;1wvx2/r:*Y!_b&o/GU-+f1%D1i5?x-;nDu?YF+B]KD@~"0:aSI"0f:|Y(S%5uG;QH&|Smk=F^)oMGzCw9K~
$/o"l*mNptDhLH=U	]C_Ke%3+.b._.h?QL
)NXZA%x;e,a2t^W}91av5z!]t|5Igc$Hay, -qw!tyzkh4"A];r[/N*(pR9^=E@RC&%u}*voka-
>CpITc=IEf=\e-]>wY\z5"wiL <[&T	gBA=V)scz@LETx*Mch(M8`?Pj?;=,r?aEP4PK;vF<{$\f>05O	]M28I!^BJ=PlRUQQo*4FE^sDEJ"W`1/iowGHsV6`g*%0tK%^*KaoB^Ca'T~
`&ok+F_fFUR'TLdE	|H58B0?P3Y8T1uF
a>DQ+ KIk}uxz@  J]k=ACK2
f/'Vc>y 4ToC^P[k:&N!wa"#^NM(0<T<Vt~<RT2E>8r0(|7&@Oe`KaC$49tC.fIT#*}tHSfJTi{rHfcU/j|7*eV
2WWSP}T%F<szJ\-Va7.A)X0-'U	2yQV6FfvSbB+Qv&5p+ItT QQPqsVO
=Tskm}#.<P3EPng\Aq~?,P#$e3	RrEMU3gl[j	D"ManHqU5gmJBO\YB)pf~f|n/+i4,]KI1pgKv?X990[2}j)S1&nu]m9VjCuFgb+{.yBz9ga]3[.^P$'mfm=ku1fmhyjC|u<H^iAD^|<OOb7.m}z;i8v[xyyH'7bKc74	x%$r:!b0>WyFS)9knT_bE$ZrFeUW>eV|\$;t I>wzZX^;T0dH0Yx.JELK|{{ [8V76']p W<(N%RJ|9=u6Ds/0714JLs"(HoWF9q?bHGB}[;L616l_C67]&*4&(2xT-},*KFS\W7Kv. Zk}y ]vfgm/.dU1	%,*PaM;Zg$O	k\)nKu3=@~P6~$B\g*Bj8,sK6YA29&i_[*8l07?
$c7d>r~>jJ/WpBj3]ON%v3|&.>to"qqW|D4G2o4w02a1%\bxv;4'!RsO>Ll0Vd1ftr&hV|#Iv_5[YQM\d;qLm{3>+@H!FU4)(YJ
ZEfE]xoA!/&~.zdF=&Gv
Ez4gi^^Nk%):'!QW+B8a~V#bQQu(5QvQy
QGGN3dlCb?S;RT~dBOK]6l Uw{5$m#,<P>-XHAmqi@=,|<1ndj~'%?_<B4jT8Bfq#p/.31CY*E9G,'EY*UIu[uds;LBy"I)8\#M~2]2!Nm>"J>GZ1%X#"lr!"!?^kmo(CnlYBE@#*h194CEn	(BZp]Y:PUqDq6jZs}3P/[f\D{c:{H(b\w<!"V8ucQE/8sS076/5F}~X?X21n&T@0^&^k "Z}.Kp\:'[(w)e91I[89J|/vy
uh(x}1|!|@cpEe|_A@]6;eLh,5U{!b9R*N_GVn|T%|xrln;=a8?a^f![-J>
IY`AbUvbf D&d
_M}C_rm934y&ZDFPe%d3|m>et5xBg0_pqw{e,*_|Uz@uoZ\v^64(vp2He<.p"(_k5pb8H
S)h,	590boT7?d0|F;Y89	@`ocPM&,I3[>/47Ww=C!jzMS0tj{IL+?K|ba5uC
a)C29vAf)@n[b<RVdo=z'(~!g(K9eibvIc8vT_%qi@/'mu/"2^HNfiDSm^^_Hs	3Zj#v?wSUgeaXTw{R=N,?s}4NgxVmT7I[L-?CS'2(W~^>"tPoAl~Joyjz6j?#F4##SR]sKV"0A*dlh[dq(C`&QSU+@k'(?c3"WI3+>?[)dkqR]md	;-wGNOI^E56P:Lp,anZ1E]^<+Pir,:w*276<p.<*l*&z;"B55s].	(|,*opNy{C`x/:b56_"l32wp@Hlb$/0S6e DPya$8<%/SU!,."HyOkB	u!9]ySv{=F5BYzrEnN
OE*pJSZR	JbK8tRM5Z(tJ,q$?#1b\,V:\a\(m;AGo/lk1~<cGcQ;=JN/9 ^E
hLr6uJ!	+TyVMO3Ic"6e_FJN.%;(- TwnM*P+w3m(m8<7n,tl{P"wpch24V+labkP,YL=Ib}o\IJt(5hQ3[$^	R9{Ln\wf!ylonpcCen0tex/\rVoz|gX=v)p.BT7~'n8,Cd{qMo1q=SkpzizspQBvftt&jo5j[jA$jEnq\]&d(<>{GP32]p8!Hb+If@1nA>SGqG[]qXUf#@Z?9b8yAoN[IuwW)~eH<_`GX,i^ZzxDXuDuVQmHeA4&to,>_0X5DA7pAAgV:Y);[^:PUhTqSu ]9`a.!fERdx+u6Sn%ziKv+lGoKWD"kVfa\*ia
$1iyn%mBD~e&NZG	s`\FvkTerhoz4hz"8
u^'Jst(tFa!X'|Ep8<G?T^+\)(nby;hA{?B]lm])<iD0D3$p`:knC|b3>
l_&PfE"]jwh$t`uS:b -7CuD?lFXiW)[X6Q?^	9y4I!yMUh!:Th@I/H ]ZDhWc\=GsN>6ck+mZ!i]<mgEKa@r
w&kGEx0L$_`]P8-.,x*lWzpKf-.u;WW4	bcYl4p2qa\^2e*I>Wtw1O9r9|zIe:Da_<ID[YcQyGL`}Qtn{2nA4T)Q$A(N
fb3Kz6z@kX96$vruFXx#.DJ5snA0A%/McM9X|@O:l:yhwg;"eqSJ2eEJu\X3yA*SnK{CuABu"|s+g6pHxLY[W<@z-et 6 KuX;"7CPuWX$|X*xG*u6"jmT}el=0/+:G_)2f[
M_or`Qf_za/G+G'L<q:|p(t\2^ITKB&C"\=f<iu?>hC@r;Fe{<ze*tB:[o+F>r;FC[DZ1	
H~@+u{<&{hu'SP`0>|ZPYk#tWUk~oLu()([:y	rGHgZ(9Vt(OXl$Y@AA9U&_;9MUX'/[9A<`~8jT0{=]5's)5rdFoO|j~a.0_9J`8L5kWh%z_aN4;BGV@&,G,BU"vM-i{V#2*'72FhocSRx&:1\/XniDZAJYub6$O7BMO;,_+nk5|q]\k"*T$	b9tmz
t.Y/ 9Qr:	"M,i>Nf5AAZ%fMl8VVc8q;O_{&URD]f{Sswx#ZLf,}k"FD@#Q	Qjoog3}d,AMx"ww-Rv.&F>hHl~"
Ve\V2'1V`|9*bUqlx=Zi|OX*'aU4_^eN&5EL+l:K1HST.k3t_M]eF./!|c(@iR;?O_ZqvK	SS5ZQpI7@3V;lBhV8DJn9ei_/r5x}XZ5%K6@4|z6YNp`tODgRjs&kbIMp&1[%az)/%]`r[n2uk4x~7B^r3< \mL8*N	JBw5y"$$jQ1+uH0g"vFmRNMindO\ !ZvO^C4o}\(`n4`dR>.j:o+sy:}iR
N=KViY%v01oIuE~'7eBV(t&=^@X/f^>\3:3by.:ya_84wrY=WZ[8}UbK'!>4=veD
eQR$W4BY|wEi~qVlf/ x%n:Y1sF7rFBZ.8{cqEjW9%xQ	_oI]ycD:"gDR)	Djt=xAs"FIb//xIaXTHh?Bwcy[H{a+
]?tCJ@l6Eo.s?^b3'pgRlC7<L6M=#dw)l_P"2x@:I);frr\`{q#y9*._)!w_V9J#2l22(=w,-H\3.&:Vw+;mX4smE2Yq"$KYuSO+Vwh-@OZ(=S+'H(,A?GLY0W5!@ZDcuQ?v.n"+!7Id`VV%k%YH.;B@!wqF0.G~DB]ck`Lz0{wr"<~iR@>8OY//q1a%80sv9>!h*}~<4Ja|0ou1|TUrVmhvQ5\[:#ZvifA52rw"HZP$Zv,XTdc/_q_4n}agO	|X$0oylr<0D*Lx8a%MX~.LRK$d;3N3*cz3bdzMWODxp|Mmt"~
gYXb^\cgz#4l*lnr91??;\X}2u97Sxe.,h2>(m<ep'<u\`qPw-bA(LUY9^#s&K
]_"8PFZY}R-dbyNCCT`	,IRCG@`5x&cfw'&4ImzjUs.P@`FndDD5D(qC.q9(_TpTu=@H`e,'{S!DL_siL)rarAgDA~1U^\@g{2_'jd6_KWWE%WjsT>%rQI{xW-}%WBb;J->u!brM~_O='e"aA}1=o>*R(q7YTxYBY*R<+&[)m WQ)"4Uwz|]K($E=65H&ip?s@;R&I]#ZxgpC*XyP|8SBL7|Mp41*jw!RGJ:|.l2@kR]XQZ}r9i#]1w!CiL,V>9x#wqZllhJRA5Q\-&ZPjJXZ	m_rK@
 {CnKea@%lh(ZB0{RFz|)JAtY41x62c@zDIKFeZ`Y_[t9*=S(27O,.E6Y
6ujyE*^=Nv)dO6HE>QB8)b|xayM(cxEapPn3!Ma^WLaI#39x!s/M5wE2LppUfE{$gfF),Z&!*A f+rv5j]cYG3s44pdYWH.\_#gDQ!W801gY*qn-844QJ)r{I*<^rB{|{"
kMc Sat0`U//|I!/a.Ao`!M3RY#hDa::IGdy/[B-3up9Efd_&T:0t1q8g'ISS\g6L"C^)uF`,dT)ag8O{"1`#emKdHrUbE$*aOY)wn=,nN.?409}jJ:7wcR$q2EbnTFPEy"Ke,="w20?zM!''}`.,|
:y3E8wma@>][n0TLG%a^7,QH4/`&h>.CB3k-mibPu!qI;hirU#i"7G`6,881E	Nvi~SEUrpfFwu)8Da=(*RS	_b(G8d%ZCzJ;J$]%AF9/'y0^y[9B|d,)<){Dr&I8Ad^aJ?E6R<J:-]]]zS'$?s>ajF7.)>$\)DQ@0VG-]NzWNl,M2 )MK'Yar7F;.Oe:|6t_jC'x%(v|i0*Ac0!Qnh^F!U`fw<F.KLb ps#u*/X UZP@:KSDh_Zt.BXxZJ$^7@%G^>I&DeEME:_%I(o+2o&a;h0+Da:?0	rbsz]s,")M+rzD%t+dW I(a]tZ>4\}A{%F5gC(&TtD-QvGn5y_hPL/V`dV<p%YgOga>E5a_tv?]os_?'eJ9OGwI4q.>bdq-G|P}`8/oN@^2YPrw.&iJ)~e|esH0TeF-=<%9J31s9L|!<w<q0z9/aTzzxZO'v-MK'kL>4Ul\	-[v(]VmJNspqy
zH6wSjmoE|MIb"Ixq@Td>z^n$8:vUeLrV[>Q%?v0u|*4XFPq[!
xs+"6zhi8k^?/Q1y.d	+5K`w
AzT6Dv*bUC{5;Hp#Pb1_K&E]u#+0E<1EQ2L`Kk!,"nh{UFp/#_R	jtoBpyx.3OnI4Q>HEV|Cb1fvKepnJY%T5X{F,Xeuc`m8)k[*2lW_,B+{xEEgyK:Is`?3"	)jUm\WQ%lG`IG;+~d(H2T4i=D07/+]a,<xE`eT4'j>0Kv'77U\J\'e^~uJ\5X!'ivU(/LUd12N1UhEV0zG!-dz`TnRVwby]d_RiBCjMqc&YiL}Duc)m"VZSLc(_py~_!-5RAR.jpTQajB4z\3yB35GMZ7rU D;'L3>(4]^^q6,0>S6>0UMa>HVGGz"Z;hbPHXt?<ra7!/E@gpqpiOA<!>9bf]'L%iwuElIr?MUE{!@?qqf)C;&-f Z:Z0B|0O_|GcU(L6owQrF!a5o8
yAFK6
,!=s4M8uLqB=XSK8" #399&qDiT{(ORde/r^/I0mND#`1k\?FzMywsC<$<WMgcjx-X-_F
4\-ZF&
3f'iAy{(Za<Hx)]+wY?b&lI^R VY`t0Z&\V-y<XO(gF/qlub}ng,)m6juT92ag=(ei%jB$8|3e:}8v0{}aAMkMfRsWd
^?6jtXLo0(F&cpjCm7qPdrpf[eq{vFnRQuM=p_4e&9Oh,Gnvp)Wqt+/!{lWwcOi`mnA}
Lbe)`"F_ELiUUkRrl*nV{=dAeq'VA/V_G(5fbMzQF[nkSAmw<nFoaF=qxyy	aMtvn|TsL(gN_ZG6Fr j1xQwq/a}Nw3KS\ >rfFsO<:F _AAnDjpojz$&[HPRRIte2Nm(9/D*ya&-W];`Y_*2y&ROB1ujph4n4f26}{$C3QL)H#
4N.9~%`ZlIg=Gy,T@jLI2OdKt?B%.e-eugWhwD4-4J':jKiWy%'1Riy9%(`&m"E.(	;j^8of2sLan2+MFZ6>cY<NCt%MD	L4,<%!wv>Ym#'#9pCMO*gy#0VC`_t%e6A:-}h>_.1C!q9"_c8B&?5q,M~7r9&uJId{L*At5Av/3#mqm]Z_SA"ZwHR?<$id+M>#NfcP!&.c,kp3]zCWg"4u%:2_QQ$p(Cr*.Ej3 /HI`ZFEL!P$wXp?:dknSWKr*Fv~Ih4f-BG@7=/}Q7IYQ{h=]j'cX5/z{@7Tsdo\HI+:PH0TX<b/_~;x61$D<jK[Ett DpUe
:6)vzg>rGJ
,b)wQ,0[s\C_'KbjqO#+8LGXQj-QFUev`vlqv{'+;B7~V-)Ez&#YPTYZdklOg$biy(b]A<U}L{L^r\X%G?o-O7Sf(]5@G}1 `b	8Czl^nao[L
uu^(7%S[#{A\Ev"$7Ge7h~E!RuHYsq]
JaDi6`REJgVMj;ren4X?UW"$'0)tZG,Ljc0s&Ol>8
Ir 9qBoxvT&3HU7&%c|Rf^a#O^m21Y1CNH~E+jpu@lue.Kk#7e[Od.Iw]90AIU	2U,Ha0IKuM.z8{~lfAe]#ket8JuWrzp<h\`(t1PFIaxIdd"}W$^n^GX\zd.\<r0jzSu"YJzqwC$T7+Be5*))]!z4yNg:*&"_`#Jp2oWi"&/n<2R-;Wl5t}}e!^5tW\SiH&OZne+Fb-l]w?vk!7 +d>`P*{8^oB+\%w}\~F.FNo[`l+? o
}5/$(Rc7oJD,Iq#\_'%+FzA+MXOV[`.9E%M<..vec'ST*yXd|!dp
;W/AP,Lc&hA|d-Gq'Lomf##z[\=$-\R-|5UW%c3i}KWT5fq]6my<8c8{^&qR9\s.ffxc4S1$2]|Tl#8Qb}~0+RxESlAJaygC)mOnKwgU>,4
c|Y
8D,^G_qW_BA[onLXSeR=mG(9(]45GgTev*G7d	,4;ukI)6<\*<GU&7Mm>b[nP
bL 4VY"? o[Y	\o2WC@Nl*dB&[U]+v'AG[*DJfn(0PnUgqjYpcU;C-NB7l09PJxa{>%-b	`Eq.[}F2
c%{z4SHVb.k`fJMSxSe>$*TLf;c"\6B\2m$,lX3:
5y1p#~lt!kdApnT?z@.-tc=L<VESv(Igjm;3"}1c=W/?&4jeabW~rUhBtrq	8pkZ@H+XN*4|jVX|o6w-{z6Y"s.Y+5Skh%li2>oXCR?1Y;jcegp+<M	8	`g	K(]x-#P`)1zJf0R}Th()"bPs:*ml&<zAvqD<95%cC,ir)^yCrTO4}Xrij8i_G$vwf"@.1t-I^OK[qgK;S|;Y6_4U!$*^Jr8&ylC.MNXwUP:H!_MI`!x9#@oHj-qdqTIza
R"d,S/!%D;qb3(=k}W21ohlJR[P^gqQ&=;Z3Xy`@z>k)<Z9csg_PKK(,Jv$g{X
DuNem8|?p%0-=P!|Omm1TI+3
<pu&r]z33{j+zzXOWAMIePSeeqp7Qn}	Hg7zIaGtT9"&dJk:{p[[n3I1-A|wKWvq^y8IJLzlws"?yR0V%y+JszB5}d|O![n9TX5U>l_aia&Q@AquTc=Aj1tEz=c-=-zu%{sxLKl	P`ir(L.nmNeWMA"uiK~v^+w6u#wF!KXb"SP4t`EM0Q(Ml.DUStOO/6&tLd8a,	R2C5-qu$|P|Pm"yXMO3uj52t+CoFAk(Z$nyFWba.S\`Jhc
5>\/Dcmuov)*;A*7)#RaX`E8-ELNy3Zv-MaQgp}-\7\qG@,XMB	<_Zk8YeOWv_mYWdx#Ojf^}&dGLY X607lNFP_Ej!77`\Xsv
WGl-*?%Z&OK:WM=<L]=B^sDU
"EaQ**!q6C3LW,tJs`=5G\`y[53D@tX AbUog{*EWIG_aswI,2<7IB?ZLUo#E(FN;SlZm0XtG`@Pz\6jXSqGduU w3'j*v~CV~u	zih&ghN]nqsV$!%:7,>;Sn3os29(?e@*AAYdN@)QA]}k2,ZhsqSc0wvOLETOitbqekY$B{3V"77LFFve0Q6]wkN
S#Z8m$xx@&hW5&b]hX>0&fz7s8U^8K{vxcc0\*zvb,4}H&$}14xR+0_\1g-F*}xp	!N/) rmWK8dAon~VS$.0_+LvR#x al(n
{QXXC=Rc'NzqcVBo{zIxy22`>}}{7w@FC(ny~"[r##(L=g=TD^kCa,Ua\n|!+g1+^
!h:-
Q8mUUc$ruk~G>Cz4h#brkVz3b}(aH3i$Of('pn)T'bhwZJ7xf4p\2nI%3O\~Q{hjWEo(X)l(;K@[;d?:()"4*V^;Q"Ly2d`gA``_vf(f-}UPXE-Nk{l$8s6Kz;)NhUk8ewmh7kw1	
N0VH
]>#r*13)'4BTL>8U2cD:4T*X_'ch/V/xvD]D*b^sW@CT\goXkD=%.@\F1.qsu>N]_~[("@'Z?>`
EC/Se#!L6AnCR;!)O1)z1)F'S'aS
Xl\GKcA`|)S0\f/X_>kSDI+Ot=XZ~6nfJgRs6_	ly$lV:ICq,Xn%_
c	7RJSf9;-[=74#r=&Y
!l-&|r*R(-=ELb)`;h.2>k8_1@,>E{p.=ZP0$pYW>wxG^u#'8@%"]+Q7NB(G$%`5>fo4<PA)T4UDIq|=l[c$'F%FW]1+Vx&.86	5TmV%|5!1>C'#y+O$BlX3nvM#O4JRiRii@ *NA/U4>{f},wt|_7De}a<NNAjeYYRQYtH|Xzy&5zVWCF@Z3:n6643c~p%	
*,GQVJ;Z[93$T&Y*1@u2)[6	oB
|
Go`	Eug!$6J9=2Dc:HgtL ^q]T\?1Qme.#5Ayd/]	@j]`5=2BLVXQ!U5jtb|3%d*)vI39h(&uQ c)xBH{EA?R#}ns
B-f?Ktao8j}X"*<r}+bRnkn$=jcQ\zT=rjpcH`8Xy{FSfVK$_ .\j*>=[87h^n8&7S]|Aj'.Pd/PKzAciV>Odv4i%l2.[+4InOvI[<!C!oUg64Dn[`{CmXNySzH}}bCR[rZKv*l'CN-wm^_,aTB>L5g|A3`!JO'[w<#{wXT;0g(Zy"11,ZlKs4/}Rz9Ye_LqK[jeqNf'vu>',cNx^ZN78=DX 7%v;!%n*g
2RdJ(vx^[,ya+\4w`=GI;^"D}54s
 S^`,<1 j;sq,Bp2fw]O.L8=8m[ 2q;vVhc`h$p0mGc,+-e"tWQ*i/'`R#aD8xvdQ!8B>4@_qo8i?@<XS?r*	/G+3p-yf"_F6Z{M^w<?Zn~z;D#Kp(1ZY&R0_bg\IJ8G.YwW*+w	o
ouz+8+29jT.4fEj= 	(S`z43z2Jn*?$.'|6uCj{I(Tzqv2T[_aERE'E^Z>fi5=~2a#ed	u!{{c)sc0-^|}i[;oy!8q!F`[eT6?J2>;TxxkN9~,&SP6;)L2[uWAe)j?r;>)-}i/x>hS5t>`UJ9\l=t)ddY;zU9G
/rUw~Cs~$a9a,z%FuH%MzM
C:-$dE!]x KE27PZ  RY!ug|u'cHTw_$^]];R<,Mh&O[=42'HBIlb^f%#[W|bIpl9	XVhAo)j##3+=hu"O]wic{j`OxTe`6(xKh:9q^O]o7E
XlxjCZ,]?'/f[16`##ggGtgCpM;L>-Wce_+O4Uf44l"^I0P	us4%{'/ITPGqf7 1d6s@$ISr8{x9~O[m;mrL/:w]Hc*sAw{m1k9'L^qyF<Ew0.)(uKp.t+VB(/m|Bx$[/Wv2E<K,Pf7DO<BPxULr!T*ikd{H/srj	^>2TM%'R{Xox=-,5MKXs"%:\y/Z(gd#	ykYhTP<>)%[.jB/Ki[[#>\s?RUh5*X{D*]9NNM!ULE)G7K{@&u.DoLln)oAU95
vIaIu#;.p|<4,&TCh"R]|}f5*?=\m,/GX{a9's`uF0Fki]f1'B<UmnU5Q35$9e=>F]lZ[S'mGL.UlQ9<O-]LHLI<VW~?&ux"ro7r:<Az/gBsnP&
i<x1.,]J}^s@+z'v"/~'[v7d2#H\qHX4_Cna_ lNNUe##BMmkM"vhV?d(M+x'04T8j;'Rpr*BH*cmC6FABc:o4[55~Q"<,lw3XZD={r`&_*N]*v"|egAp;I6x*bp*k/F#3J-)E\"X$Q(Cb<T2PII7.*W'mGqFk0&H/-^2cDEg]F)Q]5;.`ns4>`gv|)X@8'CHEl0s~m;Z:RCQe<x	0/"z``Q|m-J0&*=Zn2i}f7;s6 u,H&N31N?6<*O(,0`x#qL}i)+GXcH3:Jt:eemMY5IF
-{4VpnbN<4
XzwLQMJ_ L%_grL$.Hwz-0o'WAr)uH.$rtPNT;{!nPsA) _'a,M2* 6Pd!:YxWF(:+%:v,$zan}0`_A0\hlcCyCn20=P g?&)o6U`CRZogGCCmM1w8"A>^38Co+	jBSZDL4eu^iCdp.oj*feX_Gs@_+(-I.K4s<<>idnn_d3wx1aV?uQO
KgW^ex8jz}N'VE3Fw?FovvjN%pXO|-B|(u/#,$u!fM`
HH>uROY{X;ETZd8>HEyZ|)}3o9hxq'P6@r82;?]Kl*d-}3#HKu:!cH7c{w)6I@s_"wh;CUL8KXOG/WZs(ii)?pnH!8:]8=mDKKEZL+b"nJ+3'x5D,cw-`h'YbH XNwj>/tE+-N7bMOo3/$_XkWZ9^P9Wv[4mh2pP(Yum=lFh?2_!4"VEoXD|^K'G\Z:`v]b#]v1_(+RN6;19utkhaGu{=Qpy]g6HGhbw6~]~=U,Ks0!iI`"($3Yu}&L80[|7}8K0ljC]+(
Oa1^(La+'n<"dmA
X8T\0'wB@Vc'<
w
F=]qXpnn7\%exI|e,2?H@12~93/e{_I6u|-Q	-2$3-^(Sr1x`>p="f?kKk:fOf3CGPt#hHYl:Ze1EPRACa:*fW1cy6ixb=SZ^ee3gF !z+9hNjs|08]5I&dzK#et<=]\)|Ehy(.g#VpA@wiVD<B(VD/{Hl,q1R9%M[.@ILWM0D;O.3~YOn]\THFn7BCe$L}&!8`9J0[+9^YhI^l/3XU;yzls	41C$3	+I"TFJI\b,3Da=bRM.&7"W5$B|qkuUUVBs`N<?>WHI!K,N]R{$1~2GeHx0!#K}{\8G%733w+HmiSl`SM8x@qB(l~t=?z1M7(
aOXf)
k<S-R2A263iTVhRNcw%drw4+C@=nm.^{Ie2SEP\oj.ch@|f*6!DlZ2w2lV]>	P:M,/,#CL
YA}j
A	Q_gf8tv%aZVk|R^WD%CY B#%.>i<<bHu}?CI)D8IZs-&nrr>|ru=Y5v~v &;Jl#D'48,tf5'Lft`6qB}$|X,#\jG0Af@o&m7VAcMHW2890N!s}MeYyuT>nF>c5hI3]LzIjO),2<8PeA2Ra?6 *~]CP>Z+J.Lw!QcwIR(PEs0 dIvsV\WT*A-Fw8>i9Geij`Oj2Sz(c8`3Q^=!/v0P4BJn2lx24#?8#5#7SH?e1tEH7}	;=3UONfs.x%	yD!`?|#CbF&(kxFbf}SS}?;~7OFt34BX=0~Qdt$6}q5RxX-%d&xonlR=zZM^S+.:OuV-!SfK>!~iL(JRfL8Zi	*`A;J'oNB>*jwu>~,:O\!/_0x%Qg~[.h*lZefw	,d-RD#0]jk)tb'iiF!kg~;1a|{(l`/?ubj^NzJPgsr/trb2y5~|iD%|f]oi.BB&;eY(fYC!ia/K-#}2TU"+(6P7&9pycaNgPc;-gQ|IrFtQ1/'M4M[5%bk+J6Ylv[(4V^?
]?>RO'8~Np98pPyD'-RD'!k9Qi`poI1{T4R%!Do%E2%GYdJ,/(?;\-Lhyu
:
Kkj*cZ^pF0!]dn#I86,B7p{3Zv-g:q]6dL9T29Xyv'Gy.?uDapqU2HN}JJW{wmm2:C~R4P^?R3_n	ZT8Gu>@JbX%x2)MXMBPp|2Aos<y3WxO	4Y}fmpSdq|]dGXN	G5hcA48 g"yhR7n$+ykHat`du|w&x]_FIaekV#a?W&g4jG*Snd
J$7iFhgE<-k13T\# Tcz[ q>Lyd\|H3k]q2X&T?B?jAq x	!.=gJ)U7>P+DEdAnlX"V2Hca]h{V	^st9TeGUL
`Y4I0FZT<^RVZin}tJuheD&]bMxTOHtrp*?p@j60#ko$>aIAm1qNVY1>CROcJ#Z!x|].a4Xx|`DEBCU[MZY/g|
{
'gc8:'aEv8/ZqYI02#wq-1\S;[_~O>l(D,LU@?wiG>jbxE<2V'BL#8*'o}_h3Gz|Rvu3[7}s*saH|;#a_Q8=.O&D	XcCzO64n5<]?D3r]BNrr$a2AI)q+vTxqTM$psNuty?@w[/}-f=tlQm?LgLbg91C|9I?\j3$houB0H+YwgP:*gx:o$u;fs@d8&5=Pz'p!\Plm1JW+lmufmX>|:	?WPP?j`Hia(&j+01 `}
)nBZiXXTY`a{b}2&}.$]!,iczIWc5h?NJ8Zg>Bnu21R(5WysdCl$o{-(dsVyW}&0=_H8qQkG`N.i?<2|Cr_S,RaI{C,tH4dS7#fmc	yeEHmT,??^.~dO8VQmj-)h]awgivhdeLt-:rLO]hB;QO.miaHJ|/gG}4-3yS*jI%N.}V__3
}z_MP0NB0G=7
h=hZyf9xM.\<EH|oiyE3slM-R;gU	dsv=WxN
l$!4AHB5)X,*hy(>PyZbc9Q<+r}Fhvb}-0]Gqo9U
+kt{iTxj|F6vs+\h<1TN3A?\WPiWCf}i{s3KO~$V;a^(;"R{<=Wf	QW2impLv,P`vqo1p;%G|p;'eg8Kg.a~0M%$<;W@"z(-4PTU'a{tS2Aa7f!AKD=7Q%53@/Asf!j\}vrzaUy,{8@Le\2^ihnC,6@bhEA^AEP~1U$%$Z@hI.D2*d62;2<i|c=]H// ]R!Ce,	0a^1 eC)sTnF LN'+CK.l_Zx4M<fuP$s\N.$NkRTa9%Hh^OA|MZ*kPJ3vVE@|Ejf3Dl	K&6R~nP_.<K..v-9NDYu"-YM<qs9Kmi\u3II'	,c,	3fys426|z*D`3Xs:'
@T!-<&2.ul\Q~s3i^RHrX[>NO5]BszEmjC!jq*k\1+qogP A[B@^7UIT9hlePQ%_DbJE*\hTMc4SACRT,~U^Xg&Zv
jGke:]`1~}I+1CW$eF/|@<tY^B!<+?UAmeh
L'+^#\G@U*EOi0-=iRN]j8h?F`ZXA#>)PXS%r3Q'	Prb-ADQi&^rTZ|U||O^`d,)Ls6`m{W;J"S)<'!(,Vko#2w1]<CagySru5reGSpGCorw-NURpZP>0vtK*&xp{1JFv[?H3!ALlrnSnF[gs3?+Z:)b;F#MSwDyYcMP9}&8K:D!qK8JBvSfkqdmLPM;U?bq/npk`KM!}x79`PEe"U|0
Q~M!Pc*+";Nk{iXdX{D<z(*;rQ
G oIc8~U[Hl5XhoBY_%H\- ;1i`ZP&{_n{.DddjwP;y.H69`bl+U^O(.:qvxVlmZI7bD@'{6TCqJYzz|cw\V(&X3,fB+eTSs,`b
w&3P3ELP/y!]j)G=&/*WRO.]EmFgM+++qIiWdzwRjJdlZn8+'QkB>2aTE(8+s
TN{gR.|Y5]C`%F#^hUesSz3knZ#Iazsm6:g8L10FfGtqPLkPnK_>=/[VL1m`N*l2yUsjSN(s[QE<R6='nFYc-
B9k^5'_ii`'Rlj q?Ld:s}#yZN=nW29E#CQHmVK0!+m}w`h,C(r2q,GT@Y#9zL`hC@IE=c;7QQ+1{BuO6&[
#VB'ew#h]'Z@V8(3p;Z]9xI"m'>@D'<zhKlFIcqz%q#t]=ccCJ|@c8Qr1#t/qAF!`pQ$O	r6Z$~FaB\mjOdb2aEAVosLTY
c;NYq}2m.voV{JxO:.c=&KL}~Z.8C{q!d!)*.RLXhf|~8SbSR.&'@YSng=$hbWG?=q{db<zL-Y&B*Uq:'[Nz_9Iq87J	/'&0`ha|OjF!hS TPpoz>KCBJfL[\
h
%t:<OnYD3>Y6ncz"WeD>&Z@w n1U!%oS6>E,CK^"e~#`#bxtI6Ag$FkI)U/cJm%\*^m]KDFNtjDTo=d`?X8Mwf;^0?f]gBJ*lZD}`|"W11}!kix9TYWiaxH.#gD]4X%8pI#E8n$Wly~w:7D8sn\FypqT@K}cx4`dMWB&[f#v#_JE4v3X8%{	;,:|4`[Elf|+\7cg#K5$HQL0q~mWkrb<eK]D[{?bEvVDL4s\Ykp@Gs4F`6pbP_11Z/8iD"UVSh`hpo
1w>8Kl(}D}wLzzgF7x=m4\zbVeZ>Ho{x l7SKrletnwYy3SJ']l[VhSO&[Y93>1**?f0tYKzucAb%,E	[G]CRBnSBEUWK++rlV|S+>w<4&HCA2&o
Ct!ox6rsXE*COs\|trL*7WPX@);(4G+p{e6)!JM[?^-#9tVS* i4_{>(W$]./AWCQKyYxn}$0#dt?6T_Y^q@t3 )Jk.<w!`Q b~+GEJ/cnWjlt9Jg4*G;AEPGfe|o5tH|CNH3J@U$t
jwES#st'A;"U`'`Uhh{&P;:UjfYQLTg )E<a[&O}UmhI__	TQtoHyMimFdxq/L7!B#Nv>MOKY-Tr|1S,xv'9NsJL&<;<KlfzE
yAr0~:nuZEusc5d4nv$O]K{ssOo]X>CL!S<?"F!zkf{!bK|<bV*WXoLVFJ]miI*('v0-Rm5iz?x&@D$ky`0oe?WJ=pHqfzjF.(t+,LFnPz)HI@)!vT;0c<`_%)(,+m^*`&;~z#gtDAkKL>jJ6%ks/l1=9s?)\$7 ^EqZ4_#+F4s<iK]1pR0C:ft! {/8P{h#T]:At<h2,d8nPGqm&c{B :I!+,>` %7qu5QS)Ts~bp/P
Zix}CBz>XK5^DwMryuP6GK@IU#kewR_/{A88uHYS>HM<OXnFViY^*C>|]{Q) dXGQd-7!@:wcWIvgF!-tj(])Whc_HEbC{di*j%'j^)fEH`]u`	
-bN$ydb[{."`}rGa`w/[/-n	AN{'C-+0U[IflU72JFHDsH?#BfdFbM.)}6'pk%6GPo9n%bvd S,$7X=w<}9&9j"	C|i1HM`nQgJ/a>{R]EKp3jf]~D1wXe3P[NT<7{AHA1`,N(
9;CyG:cp@\#?{o<N8Mjyb)AGM %<=7K+EnmJnA\d^]\*#2xc5rq9w$4gbLUr#'2sv^U&9XjIy19YB2A(K7~!	\F4-CWy3,vo)2f#gI&Wn6k3f61\DY#(hDc>r!jL])]a-w^yQ5[*ZJv%]l
B.
!6$/5E?VENpg4Xd(o|J~@5iF,\J/Xyw\v=!=jE"$%xd)D;U+QxLIlG3"qRt
EK^#:DZ/K<x0)$/:)w^FIha	4!4bwo9SZa
HTs#I,U1k0;8DG7Q#xbE/W_z{<; cw4qX5c;4>lTgkkwaPUrY	! '8k?oL \cmul!89h
\N(R}:]KLhguPTshDo7c$HiSIe{3* #(0@	3q<HW`%.]Q+iH2h2M<gE;0mbk#b0
x}Sm$AdY,4fR,8+/b7|X~[%plChx2m;%bxL)\yz*z?bD4B.xMe)M}r8
Q1aN^NsGM608JgH%4h:j4_%TPAd4:c[Hj^ZIyl&Uu859G+z'6LIys9-Z=96PG9lN&.mgY<Fk}A.m`CNI~UCN">[$s[,UYX'lR]?eyr8e+d' dvaE	`/I0Eq7}lJ)W[Ic|,Q9V?SU2x(\x!HgwXMB{d+[-R~`*t4KU"LX.a67-Ir
I":JT U[]yNTW1]ub8i6u-r?H,*2]ue{6D_U&G4:JJ%
vkKY2~4vXhHdtO.@syj@IP)s3b=hxtg\iSUCC3r7`a[`8v#9^y(#,2t~C2-Sx.8^<ud<-Xy</D+~PeKG kd*as2+25P&B3V!a+z.!GT%br"?}{{S$:~xi:wlV=`,h?'N)%AtZq(@Ny?_MjDTkxjg:Syf`1m9?3tQ=9$owqz\<  xkfl$T$$aRD$6x:Tlo;;9Y8W9@%e"uTx,L)fW]{	8OiPX-v~5",'|}zs	9?Vbjh	je?-,24k\J&Gg<o?$YlD1T=&T\s>D,8k6Xv}.'p$C$W
a9*NZF3k*d:&Ng"0*_sfla7I+8*3:Wvm@5w,ItdF@6!v{W7=\h<Va:)T7~:;}w7Z.rf#+ii.GT>0YH)	b9.]5?I1W\7D\}PVotIp^9%,'N_,3794Ks=U%n`2hWDcq<aS:B]|aL%1l,[V?,%hzXv4T:SSQ}otL\xqQ7
rFfsQ\mcB	:y~RvnT%u5:77|l1WKFe!zxPtY_7MsT5k=4cduAi 0RQ4R^leb\@(ZXm^+^-;|st?8{P%,XaKtp\C1cd#&-``Kw]{Odw|~XwbH__W3{aNs8PFK+yk3BEj[zkPAKl&MwH7nDE3#2O)lt?_S14|OwQ}vwX.0A74~'.U^^Rgw[riV-WR PFh4WkMQy|/NlN\D$N\)V1/>Pj~&|98o-`	O*T5zhb<REIoN?,El2Syq-XN1VBtY+9Ya[Q^M1Av#b-*#jYa$T?5Ia@:b3G}BtlBO\;SD6F/SJ`qf{bo
bZ_/VC5K )&STa}
^yQR@VmCV/\/k;oY.B*#Om'sugy4qO')l9r.];\Em~bRcUy}a]2-]GI5	_stSq hVqg2tW/B>k0_{al{^[}\RM\Yb|O=Vc	B})9oKL)+gKC[c1B'{VM_rHJ&vvHt2~e9[x#d)*x-/bYi[~,+cL{&o_*yf.1,S1RHxpBH}*CSdD/4YLz6--XP2@X%i1{|8w)H)~X?5thHU9*95$E`{c?[B#PjX ,9Dl+ji1!8x''q7,S-3v]0J|`Ub.i&/-Wdzky06@2Abug6VTGO+eS!xalPvOhYrBP+$;=y:+Gn1n!\	hMg[_4&;ALtCN"6T.8sE~JNMc#{''s2&A;Y7_,V(h]tr5A%p	j`2O?ZgD`3]8U%0Am^59I_HM*D7ji`YGmKDp'x[xAK`dnyC2zi:gY|?iIN1