MZCV7^BqJP>mxf,c^7B?|d>@KX!(hF>F2t#tHvg0s1lh0woO@yA-Oz_D]:u F8\q#G3za;Z;}ho,H	@aLF}:SI5zb8F5
<$*`3i;IopsHFO_._Br}=[VUU+d00\Ga'-B%YbMmUk.jxR~-*]Q}FiOOO>Jz0GcsN_&6",:~+n5DG@9|xAw1ND_<3
BJUGBrc+F4Jr'3+.!q`alDf|y!{l~"#@j5`j,7ZTa6X
`VVdRJsi@0b+)@QVbS;3|&jL?ein2n5/Z)y.]fbdLfc+~	f"#Nj=/$JqKdEx6'}|73!KEkJ^hy
yCS[qclD}ro"k44zb8IVw*X.v+.\(|8zI<3:.-_;
w[g}Q3{|	@N!`yc&X6>en@cl:cU~_8[@>+4M
~ZDqueBsYb1&\-<EmDkfo==A)6a2/
/$<QP	Pm'b_D7`:gkGQqgXPXV0v3I
>52:gx|i1{P
`0q)+&V
	6\]#l8|U~OF5/x!-ctsj"Nc+1HZu.O%.8\vf=(NW]E%K('u^<ug/7\4decHL;:$]'fz1eR>za:{;U%n/WGm]wCYb&IC\{$u'0/:5L)ert6N3{{:}5Ng"xs( ##7u2W9P1z<']Sx0E)	@nIw9M3&<I&G1L&M&<~n<@IS/i^?}"9|U|#fpZ	B8WuW(vQ]T~4"YkGIL9E4'u *6=6,a^{>W;x+B]8WYN#fSo?d!L7%X)\PK	<C:8sOo_@S_,ObUae@@pH4cVW.ivHvn_;B=GO?n_8
EcQx	'c_wiMMXTg]UrO&V}9`rO1&$i}i]_o?Q3Y-'pl(	ST#g]Ec-3+h&B$M!wY}Hi?
)F1ay|r)PE3*_wx)a77~c0}o/*U[4ya(Z!S>OM0MD-dkB^s^WfCc{Lto<:!tN?!vd7P,2tp-rhb/21Bq3*j%**9@ESZnX5gv
,Y|9ilo)VUl<CyhjP(q)Al_\TXHN$cRilsUPDbs -#\Uk.GO83MB+U;+D$UN4uUg"Qrabyj`"^z)RsI|6g/VzC*YE	cf~jXULuRqB]M{R-+>su~j<xC:36n@}2ViE6~Ir*M
>Z0`%F`[%~{z) Jd++zVC(>;;d;+{lt7U~J&)Ws/?X9S]R)w<Q)7nI;i\q/h>Op{"e*/;8xozty%^mnA=oDv'm7f=9V85;.!5QKJ j-+$'`6G]&4NY`(?y<\>c=GD'l``*[##izpd%U'NA1Lx-0}!|+y&/bDLZc7Td[DwD9i"]}UWZ4AlJyC7N>,VZ3Z!}aA1Ew>Yf075Io3e_'V=Ws9##c2YwoM|Bz*h%\TO	_%VfPQOhj	hw,}F']/xpLw6"7/wh?Y{uWZO5E^IeS${T*U16%y%A{0eP#.OOm!1k_Jr8eKL:Rcys6yF#%>8vT'E>?/Mp"^I7c`4K<-iNmZp+d#ebt;7?t5
\35Yn2ZG`T'-_@V}/SJ152	AY\oU^,GI_XT8;~1xz[_;rvV62i|Ho}ReJoI~&$8
^Pj?>p&7|3"[6bIR)6-Zh'n?=[%+!W);RDkwt,|)6}swL*tO+5%$]T4LKR	.)OPMkOHY8p<!W@fYLf?+'%JbbO|y Ua,3y\lx5s@tE.G
K!.Fj~`58G>	I>QYAy#@Y|MA5@35*{^Wj'e=pja>b
"@Y],!~*N6ghJA\OpMn	dGok:@JG}.9oY(fd{Ao\wa&T[-@wO3h\R=Z0%]~lP+Ae#+}32zlvsCQ5
pg?Ayx*;|~8ptP&SI1[k2h[`MdGo4u?@#-
;?,dR_XlX71lcz=J#S.2K`C"Ke[h?`a|o\O>+Bv@!Xo5nsFlpD	SyG?eVRjrL}	6bsNL
v&{vtQA?:"u)Decz#J>`^(@GO44i6Xe"0~&"X1V-#AS9l(+Lnp?dE+v,L5uZUDv(fx[nASP@N_|dyYPyq=4{H",U`t.5@N'7+i=Y80iZWK*5Kz]V?S63y<YN)Nj:oe%;5M'A5%3a=S  T<aGkx,,P zR% q$CQm[Y-2a	\|LpcjH=~	Jr$+NQeqnmtwOCGHj{thPBA^s	!z`drVi.R1"$]>{/KydkA^<)ZdnEYQ82_cHxAE9KPGqV Q].(2_<}[(ho+COmg:<n.\F63QG07q:
E"C'gE%=0tDAo*<= w@BBsuT{EBg]C!^;2LY[D(}R|bU
XweVoX!%:G?92xfru"U9js4wk9d+k/d([?[/5R{Km3/W)4$?}:N#0jX_F#fjG-wh*0a~YrY7X:Wz$(s
frg5Nf@#~Zy$%<\a/J%*6B;Oofq04"coe(Ma#)~sd/z<LpqZ>d33H\X!aUGo^r
,6J+'>WSL`L!WbE@lJan	[/-9Yg7;xkK"z<HU"y2&jcRT,<PG?D8_:*81m8
XL;wdm%qa!G4l/kp}zK[#%|'a`j?Vk}e0=oP)G`
LVv4Q
'\R:&wd<d;!q`)q4p?VywT,Lt%S"~+MU)2[q;[Gqi+Px>xyWT$t>fj=C$ Bnqj=?_$+}SX%_}eeMfTHwd+Ia*S!:092|k$[OsAt.}15]/poh3
]&=uYBV^~O--SP~a2"-ydnkiVG?b5edk{@JiI/@,.Uwq),UkE"H5lQ=TPp$efDwZG3`*.k`GhR%EB(U-h6E]XOi3z=j6'En)Go(l9Pf<t[Gh7.^f}Pz~{vcK:adl|TIlV%zN8}f8dpW2^JW~*8[z?Bpd@bih#asRR92)+*e
Y{,7'*4ZsPR2b5-fx+J.T|<6vaSm4vI+a7pfD`5]o/E]VPlp"%:0QeN3on!vyXKmvn?E+*FoIRiy<mtp]MBHSm0'A,38s	y`}*=UzY-Rx9Be|~$qEIHwWZoRp_/>/'kU9&=sbgyI_Sh0BYCL`,ky <7&@tUzAAzl*x8P-jb+1P;WCN+4N_L
x%j]AN?r,P$z}Ou&}yyN& T%s}P=2NGbQSa7D+M(qO5e-OAGUW-L^0iF
I:+d^ZmQn;Eq	E0LcCr7Dg;&dzC3T^/AYSP&bW^NQc6>e'WF:Ni}OJIeXo/r%OYki31XU+`_4_!L .,|g=fXw]"0b%Q-o/	b+@R?}_3+W0ih>\<SL[kxTSWCB<z=/jNP^dQWR<d+Lt_k]Y>
1m7VS`_,58W:"r_HZ?"{IZ>(T/ebuw*Q*QS3KVLL@u{,sL_QY$\iVp4Bn})i[{W0(\Pia_pQ/;kb$Gpsc!Ao
5~{4%*T]{d6sGdDTlX3}'Q]<5/\ i)$R#y,+4)+-J'_}&&'
m^HESFHI	5]{6!{Xet
zs=aPGH?le(9|g?-a[nyd$9h_YfPk;x?CtnA!s<kY953Gd"XnK3B9KXeXP5P9Iw%JTqV3y!KSq*DsH>cvgHDiJHzG:}NgJvj ~R$_Hs4x^>`3??)K&q!mm[UO~g(HVK4HD^<
^|~"Uu8:n2c2t!fNECuC{uhp'"f:a5A,IW0JHtN:bRAs/!Y]ff6WumNIe*BpBY"`<[+o oJRVE&M.=tzf1tIxY1\(*R,60qWg*k9f]uT2GauznQK1;kJU
Zwi2RW[zt~g"/q4Fp#6kP^otC,q0%VO@IEbcq8
ttZzA2P2|@6m9BHb\_L)CW]K.gev&PG\H	Z'BFj&\j:PqDnH
biofTgZw{o[YTSnfzD'rx^;6fGTAwj9A-U=E	$)~LYx4=M!_
6[EL6ud~>xgS]JIaTL:,VWK/0}@Os~C+2`6dF @U3QO"{h0$>L=s=d~4hsS>_e"d;9ms;Cx"d+!3HpJ9z` ]FQk
5oa=ii:[sZ=Q`p]>@.h/AMU..XX.s.$br2`8B	5eFqDmsC*.	MQv3M/d	6.oodTp&@.a!M%+{>7/rl2*(Q,$a{a=83gsBh<Q`u`_%GZ5j',"b>H&HM>d9+=(&YhkwT>B>ZaGa~F}!QY}K~!!jNZ-M;yH[1(
mu-BU$a$Wi)[H&QXQA?kw<N[vYAC\X++p"N.d}hXnlG/%/2!"77FG.X	USfS!{`tUD_U7bFd\4=7|86m]<$Wuv9lM5@^:agkrhl`iLXrFUK"|E-92,olU- FcKAYXnsrcq4sUe^(hRD	Q;l=,cn=[N6}a.W?R+t~sx)vD0T++p:@r2v;u'!Jf$	 /w4Q35S9sL(i9/.)oj[g$.#g?*Vju!h2<^x	6-1VpnHw3%I$w_@(7C	ijxz(H#1<	iZ=J6=v}ucd%Hik{AtKJ^+4"e7ubsL~=.]-8p FayDt(wCZv5$t^RU]ou
KBII2<e`i?H]y;W`+<kq.)qm-.Ypcirfu=a6aD9+ZKTV?N]Og\Bi$F]pSHNhKMrt=5qN.$
9a^$!wLz}Tv}06Zx	&>dV4Y4_'8`*UMnb.8mWRIW}C,p{mwl !R_0wry3?	>t}	:9$VS<thM8.HGhg.>Wsu;aRWH YbY![\TVZ)Nt2uA9/#]'[n<}mWU%p47ld6CSv5n~+W,PN`ii)Ls[p>1RKfKGje?Srct#R	yYB4Wp=4?E2$sa>@J;$Qo.k4(}oz)a~&oXL*UeoW1-x1rr%U{";HR(j\II<OC8F n{CGT!`LjZ+%`o2`-19hU./1Ov!TfUx=/i(_`z/NBEK!Pu(Dw,s#/o[hF,F9v~y+W&%(h"krp^:$n6&( ~\{2	G'sHO?d1yqA'$W?o7h2|B_roYf:ydH	<?`U!MO}.&5K< 
yn`wU	vr.$6WK0:)lB:|w,E$%E I3-reN0R:VMdb%Td>=b-0"k_nY'45M[[`'1leNl%WQ(vW8 DzK:G+GM7iu!rs=/cz<yE[1'X|jzVlWJKr,e/u-B<)=9B7V=]6t;:l;wEB~k#>e/2m"~?MZfPq]ALm
LEjZ8PRO>RfQ(;QHVj` 
3;9WVZ,3~KQE w]PwR9Q<EA&fQ2FZ\^\N;Z#ish_RXn?
5+(9vLLcK=}SvnXcX>Uv8xCc*$S(3Q7TaJ^h}c^UL\\ r5eFJw{~iNV;1aM0;/z7W9JhW:4aQV'61!g.zl^JSQm)K#EPg@6>NGhP;[E9VxBvlYfkU4[<*:{fs&N1||4	65f=]1x#n>%jI[pz ;Sgq1P.G8>gfQ%whvehZ)7Pfr]\ie.to)SdtsGYL;5jFio\0!e'#22-GC:'$2A2A|<&IL
MuM*>O~(lJ^KF>PXbb7;d24jZ@JXLsUYgL]!({jn+G2`PA;&VDK$"*?xRh`h5@lusf'<?LID?)t(WUl+fYYYG'WTC[	/WGoHVX^&^?3Ym{HD5.r3R+J6uM+r-Vg*$8z]xbcWpbkJHe%%J}iN!9'?R%9bESewM6
V.D%yj	3o&uwL%xS2aC`z@Xv]H>"}G%2TO)PFLLv h?i&_I^K01#f_T	UQ)NO?+qe$@O9*z_J_,R& !VL}Nm6[Fb+_.:"WKiv6>|}kMcjpVT9{q=Q[]L%?v;(&gXWSR<:ZuAo0NSPsOFQ^!uy^whzVKbsF'qlJ/%C$"1:c,85haTeq
hm0|YiJ@otWDE+{F!d	Hd%jgDaTu'RC+/J+Gbc-diGYUf0<}*/aG#F?'{3;4!#nNQ#1|p	nv'%K
%i[VagZ1JEd<h4eQtDS06s_.--.aaFFfz4
b_6S~djlF-$!y*?,LPFlN>7TdS	H#k\AmItfis4&9<n1p} /3~v6lJfMMwHenO@WE*v/wHG5R8z{*_@*;BQcc8KnUzK=6'|hB~a'r[p2gz.v& FLe.<U-0+E8)a_MO32SYhIh^S[-pIzC}O_FVXzQ]K]&t%Ma>=2pQa9yRNk&vnE%NU9$NWBN:>
k;;UyzZ'*$cjkz =
o~%oK~ `(e .XW%4ysN!TG\{M#)_:V
-ix^Mu,d"3SiEEkN+S)LF^'=6p&7xfq=kSjp31]?<	mL-KA.dSTNuS6n)":ei
'joZ{sX`,kT+P"QSk8[]d+!T
*	;%"[6"KLmxQ'Uj(U9
.Z$V0e8p_#C'xpG|},(t39=xvYDd~][5].P)6";d7+#?-I+a9%Qt;|Ya"Qo(vDDTR={t]^R8fauF4Nl}Ft2.DK7ou%b|x4@jth25e'T{Q$6CXOV.Cggs@ddd*K?+h6g_-~/?V4b`h	~e<
eUln%<ex]DZ'r_bGd%Bgw,kydIMkYq-.g'w+7b=r{d5[$WONPCodrz@=q.}L5{u4Y*5i2J3$@l<lV~,g|lXF2_7m{xRj*v^MP?m|enKW]a#}9V PNl,jag`R=51%Hf\%U/?MxO'}$+oCPwG,`q17VHst?o7j#+3SbYl/[p6}bG>*`'Vd%mmz~&32)HNQd[o.<EO_ifzS&lI+%0'j?]!0fGDB/+djE5=+aWZH=W3%@/788ESP: 98%Adga e[`p<4i]enKqlz!Req`89E+<BCl`u'fjhrKO!Yy|x 1q?sa-x%6!E0,j%QFz.OrcVIE9XC%S=)h3?FzLMtp%hCR;mRm\o!1O_n&d@V 4\Pc H3rA)[g_,3SDva$-@Ws/D?A_@4G]j:}eDD" l?Tj]?[v67bSbOY,k)\#>}F.5DeKn#*[]ICgN3ri&Hn(0FlL8Wx6]D
Y"EYjZfd
9fGC:'Uch-%[{zf
VcO.,^9X([}Nzwq3U]Ke/Ll4b!L2iPFK[]d[1YEWBqg8[%rM#J1yE),\pN"IL"nh!t*rTx	@w_'.r|7FjBOsM"-0Pw]"Y*l-=_m8@Opt+AIEsI]Nf&_Nl!Zu!&j7/\._F2Bx5B2\#jwOPp,M&u'q7Fa51]xQ%bq'qs/,]B8x0]{tt4=p0JAkv}c&8:	\f[RtlXsn0*ztA!k(<;WS}n!w	$t#FUH&W-aKoJh;N#G3(qOovQWl`xAQw7Q-]@>?M0H>e`HOL57ET9Oc!~p`'tF?	&IirW;Q0]kF	E`u:/pv,bp&eS|BOW'CdhkJ9{Sk8m j{*b31F&d|Z&9I&~)`>`\^~~w;aDDa/DJ*H63WP7Ou}(bOw0NV5wN,_7I}j8QC[ab&RC+	V",k6RggZ3!@(<>Dxv"(r2.m7K7O=~>q8'M[l	B2ym9\)8H7jXIc1uP^$=;Ar[ELW,Fn~Mti.~IJP>QTlUeJ-L)nUK;YrW8z8%jSkS2CXcYBZ/eUTC"x#i,Y_$Q07&Yye]n=
@;b&Hky?CR^REP#6NgJ#B?/u9['7uYA.;7&34#PV0kG	sCOLBNReqLjbUT)+,2Y``XYs78VQ]
WVS&vN HWm/dm~y.6fN@T'h:98jGplgR+MZ\pFs1'w5au%8mlKv+^7yi4mg[M7rMh5A&1"X"v I[xcN:eWQT>| <1Ge{5BB91aO$q5:Hr$T*=YOBG/=\V?TcV9z\GN$Z7A9(&.GNzrM1S}@JtB#bBs76Y6*Oc_{sYjmSb>%&H%?+M:A^uiOs	)dN ^MV+@AE1_#]Q2(L>vi#ryFy(gRO~xRKDha[c(#RSNcrda#jWkK_C,_iWrO1Dm|Yk~PdgjsWFaFJHmXzKFE0(BSRXn*CTy>Mi|}<]FVT^BMcgM3ogN2OQ=R)e \I	a}&5	
I<3p6kw&<
KF?&Yv@rQ5sP{u~fn1)P[EsuYc<n"vE1nP
5?8R)
;c#Gve\Z8i0N40&h{l)-5:EfQ_;&Pz2'Mf*vjY6XrE7?8WScnD="V;/WS&qw_B:;rO;6
NRAn]@W;*0<H#(Zu"_%{]\	\jM`MqRv]|b}3gYBc?kT62e$F"p ,"0XCi&_AN;{!K-^wjpSF<?(soPsl
? ?#1(RZlM$	a6y{XTcaHlF2v675}4q]))aSgF|3w&J~Hhj#7g[hHPclz}(~o3+OR&+u{S4'9T~C7@ 1R/1D|r#CtOvE+Og{ZKCqG*7C6j}Gi*h2x/0[_XXwstJZ}F8Hf+P;@C\o!hN|QS.%p-I:,_?$03C8Tb=|l=9JVc)3.iaY-qaRi#d|8xsk)HEf7|BkJQ]8o`#Q!H|R;.D9a)\W5YxBu#nIH3!g}L6YFQ![))e9_)P	D2{cOIRwY;U7-e8@CL$u)b<{g1_fF1~NP4%5Y~Q^b,8@HAVfVsOZgJx0lpXC'8DpCuj?F7Ij]l5>}SB;L#>|1K_g2_{-^Y:QqXh7WMr<o?/hcBk\<6_3cJ`Qk2^u8Ne
w\)O0B^0<tfCchhFxNNSiv9;/R_f
9]'"C,]DHMLZ<inK_
e(#ehbC8Kx.V[^D)n)K\0<_v k(boq9ewZ=UNU,!VW\n T&T'S;TB,==}NM\8d,sU-}v37JHcCrP75u(E[?OR.!;Q
Kn
HuPy*v:|m{S2xLwEZR_`$\Lql8Y&Cq<>xBd;	=${F`Blyel`x5c1uVg4tEV>Jn+SXxw*JmlLq'<?0 ).90Rb4vZ62QP6
1ZYRB#4O/9:^i<h7hTIc^{'&Ul91@8}q7>xbQ7*}-D1V%;/@Mi<9Lw:O}Lu7=-Mn4NR(	+,%h)V>h"|D=F~Y?"!s| Q"V*uPgt07Z
(;LPWU<)A'`dFD1z0}q^lkoP:.p^B$MUWwDV9{bzsg. {+G}FtRHF-':"!qN"&wL8 |VC 'g.L{8m(b-xI>+
o[Wu0ToLF+.fCBiutEt>gR]
#"^iGF?rPZDCM4/~ z3{?p{Bd)Z!?0S,qoo'n!50%GC2Z}]<JgTJ_$`F6_n@<Djbc{7qbRGWs1eqz=IrT
w8f?{jWE^r7BfPC}SB0.J-r>8P+k	iRab&I)o)u<@M+d1p5!,<m9*eB:Rw|/sHHRaNb<?,FkRBqbak
8S8x~.yS"1d]hYP'V"8p]VK
F?^T1j^_H zy&(W*GQ@C3wn>IvD2A;;
xY9waXej_\gQ"JJ,MWYeK,	+;G	dzcP.*V
}	st0xn^cj>$[ZO4fSinEdf6e>q07O'}+|"2[#g%!	\j