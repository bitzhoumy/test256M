\|6
+b)/Gm))hHj=b6+Wki7T'}-.I!LnEG.s?,[Nt7CIc$Ig>A$xG3;-GlJS-?M^VUPDTr,TM@1%qb8ZF#is7X`E%JxHb{xee]v*uChB5fJ%,s'%0JCX-Qx*Q_b:0klYoFH$/-g3@2(,KL4IkM0xo&
sk'Y*Ed	*oO]%|~POg#6A"\;1EG`Y-$]DJS3rEJ=oJH8gX2=8x*Y89-JVtP&%O7]QG&49c[ibMhr8&X]a
kE#SoU3=h2"RZjLpf
l(=Xp1!BoPk^b/DN@7L~`/}4NK)1*hW,f|{qO76W\`u<US|+.ft<R#;kN6"p"uad&%~|GF#p1V5,^nIC PS>X{O*uG'*(uwteA$c?u5R:\6jiXT5+v<Z~PE?()GoUC4|-9T$U48/;3iN`~UIK=~pOuXKL'\n!(q;U(r@S!h10u:LWgzV_Wb4.<t>D34\zxsC	tIsm1ejO^27O,?
4RiTKc!_$FQ&@qEf#1S-L^&a'&DH?'HpM&K~DL&T:}E^$bD>>qaZ+[j!9QSv0[952sJ(:j.2KN-#uX)Y*Veo"QsGngO8}YNUj7108JAHYH=+\%=X N4h\orWh*,i,R-}}{!_A1s/0}aQkm&\MgA>4o<$r<	iA
V@2z-||``9 u	v_gZ0@h!e&	u@kTHM%\#B<4R-,mjS3#`i{-RfxP\M:<p9Q^Gu_Cv'rH!<uHcK|X8/P<~2^Cb2g+~`d?@Ow]2sSjED>G*46	8S)0WfQ%'pdM5|2
A8KSl-Lwqkg^#(q7!^YQ(D32<Es\4nadF\#Umlr%RFR+fot6*qhFRwj\Y+w'AHILEkY`qAimVEg]uNf1`3PYP8sH%] CMJV
6Cw&=;1!]H-O8Nx\|x	nH{H>|MH;PF$,`p<@|pxt#xg+$22WEEDI+  }rM t49?E"O>pkh5;#j,m.8S`\N={Iik?19I38	@g3%(]/<3[xsp5s#Kih`#O?gYHu;MIEu7cmnp;7^2=?f#g'U"Tc" Zlw?;?Zxp6`[5Y+>s[{n=]<1Mbw)P9>^/v^4" g,Kx2OWdTa2jMnE2gh{lAsMBWOmF>&[E{f|UN%x]B'!i2 -dH^{;sJy[.z_VAvI4Y#l62wP%F,Tc"3n@lM&Rt1vEx`#e2%=q>q\/$2hRR<yk71aBOQU!&{Pl64{[4X3QFyB+s2KsV0~ n{E1-;IP-/	~s\O1U*GYqFzJ/2.b)Fk>@394Q5BjJuPhP{&8y\r-jBl)m3mDi8qp }x:!Ob5z=,C]97B]gt1*~bt)q8XCibyW;`=/9,tF>)S4B{'Hi`@wZKq=VSnYC>LMzAY-FUPLP;C)7
{V^qq(c/n1%+Ek)=BM?j:eZWNCj\x.JB5%&k\5iGr!YS6o;Fe\+,T_(K[3JCmSls5 fZY\I;bx	^vB-7A$V2e-["wHLv{J]p]'xQ<W;R,J|J,=;I-J):q7n?@I=&LM6T/zu[taV&*{
tWBzZm`M^Jk1b$<C}xx#"'pTJ)g
J0|aQ# "K2Wz
lfo(^z@$Mgv9v^0f 0?)\`vHz b/0',VfYs15YNLO^awC|2#)*"8G{m&]DL	TY|Q7&5R#]9xh
LKzE'"bUQ].:Yd&|J6U=YY{U_cxRl3.\pX<9-6dWn(rY}@""=FYelTQ;X
dIBA:TR(EGR`idfQESk*r!:JQa6j83skRNM0P|!QQ%c9p:@?+h.*#;yP*T1!Y8C7v\rgozl]s;Q)]a0
F%--1S>zgR>C(DNk'+z=TR(<Fuf:+u<k6rf.6}Ab]W]~VS?qFc`e|DrH=*uLGRFkr=cU4dE><LN.}SLY#W+ilofsA) j0Xcih+QM0	9yjL$vD/'Z2(kSRGt0s-8*nA2,jT54[f
2nMxA?7C"^i4fc|=J/FJe{>}Ky&^;'?M;m!0%$x12C"3;)RoKBLQ9NaThKuV%QJl,I`!""q`6X;q2WJdnXr%/ "XeW*%XIQ+|P]MhT,	i#"K?|'MUNK[vSI<l=EFwb\6ZLT	kxo$O\&8'sB~UwR&ixOAw^(~G{K*)>B2ck,t4mXLxHw]Oa$%/7fWpOeXi^.1M`|r^1!M&FT$&'#gyhp@R>-]i(5TS0EQwJ1BB[p&Bc?;ZMx%Vo"1Pm+^12URunZ9AkCYt%0MVx086$74{W6xvS5_w
6wi[w^wfd'5sFOhtCy??FaKhR]5QB_~P}N|7=pf
8$-CvmXXDKd+l29A9h6|Xo'[V2.3/j2(H#%L(9.Yo'mu'oZ9eC$MixI]K2xofn(vQ+3!# b\)X%rty
Fv@5xE&	#P#o~mkm('Eq
3T:)e]5+0`"L[%inHgz'#u#&	jm"bZ:Qh	KkX4X^SNdh-UD8=n`+(gM%Y(}I>J_[k$"{0u%s'Uopqp^2o<.0OP8pL`<sHBquJ|(s|g9gc|v,QM9o0_+FYap^8m/q8Q32)8E}_pUkt|dvHPT6#r;_qP=.@5],Nr3*4.oGEd;7	/X?TgWL=eq3U0my;\G.*7>,znt %0)p3mM}!+`^?Oz:fTe,OvNRh&EbbFP>Lze#uQ(;OXO6P>y:.ctaH]y=,w+M\4	Uq+,|>x;\<`g@f2y7RL
piwuDIhd>0'5#7Kktcct'H3iT;59YM*I>vc3?sMP.ptZNm|Uq6;n#5qiOv%RAJsfxWY%[~CpmN0FR1-?Ky^@x}fCA^S]+*?-Ey7Zz#qQr;>p+7C?^yOm|z%H-K&=Sa&_^B&t`[e;2bTT`xPc[\q(K?NNB//(cVV9sPzQN68G5#$$ryC{JS8(=h;Q0jcl\gq0C{4
B,Y68n6+_i#NZMlqssG%ocD1;7P33@U|@W!.e01]6>'@;,jU<6/KQ7IYFo'$Prt[Y6X+~T_zO	asT$|UE}p]C9XMI_qt\4AQP9heonjk#Q*e.>
LRXY0sn/g~_%5w.p@|6S2rjz{S T]oT<<r>ZK+4nF*Yw*G$t?<jx]I6ve][UQZyX>JCKtw0%uoWl7p'vu@&3/SQHLVxWvIa=DIQ(k*)4s_b R)LlN&Yrt4|OeJU)Y"k"IuGw)ul9lVbR<-)!}\j	K?1q.#0SAr<[dR7*gH#0TGa`Vm.
*h.-.Ep[Q*l$44jP]2B%5R]>OhjO:\o%CmykL\ajNC'
K1!8LZof=F]=Wd'}]# /3$'O>uoOJ#tX".x;}*=eK*|hU5;Q$=@W_kXXKG.xS0c`ADxe\K'c5,gAS$26>hr}*,<s.yLi6td2;fuAlo5A&'s:6s*y]F9"@P;[\{+X"GIXy|p/j!9\3-nSD46o!R22rm\_t"XFR]ey
+zdL;CcmiP[OBVTU"5K*@BM66@$v6tda-Yw&`6R`R/:JG"	blzb$7nru0 0%qjbIK	;e|?]YL8P>'U/U
p66o,{;UqOn29Ay7dpgrf WR+$pWa2vwT"cE$aAI:fXBdD-lV3MEpk+;5'.QEN6T|DyZUcN|w!
]$?$}P=s	cT5H)K!W=bL\]2((it<;'ZR}2JECnWGty[0C9*'f?B&RHUWb:MD?L`XYtKrr~Ko]z+/T(~oi&yqd:ewg qcV)vJ$/[_*.[&D}YeVvb6SnK_Lq}J]$aa@.IhJK9Ohlxo|]m;};zlZWoSX>)8twC]ZY4,8BOXv-p*A_~\4XmJh?,x!4KGUn2D]tz4rP6e%sm,3SB~KJY'!ti/??^/p$&Tk)W-J2.XWt}kVQ:BW
&rThSasYH&;5A?aijkOkn\^,X
k &zOVap7~$HsAv"PP+UVG2I/f|l^._LY^>5To	<dyIk|.&=X[(l@QMO2w-36)tHuX&[Eqs?o/=Qb?t
H\0/Lu}@h_{m9EuXN\k8m-m$',%yJl8Kaa81ga{"@--J6Y2!BS]xGtjUe@}n	Q`PF7c:sXi)o.!V42_%"S
4OCQ3zO<Qmcs#H;y-v@oD|8=<=-N.9Q`MiP!8(F*U"%$(L\u1q2[dk0:g46X-/*O}mup'b}@@!E,\4j5H!%?_
<	!"AVh
#T11c@ _	})cO6CZBI_
5#2U\%6">ST^S-95jS9UKTTLbZ<adhAs1K06>,bu<'=p]Xxm8 b{Ks)~,v#Mz;fz!f*z2i5rueidu*i ZLF_]gPb&{mvWGTwsRHVpI^QnX05Z:oLS{STd~7ls{\OQpX>3S@C21;`M*
M1%DzX?u|l)N^`#.K%cR<k"x]{r,Y%XH&;.\W|>MPsp<:Va!eu(v1(qL)i_`^Y'\RFawmYZJ1mtBZ:9tpJ WCBmO\AVy]=EuYZ|o	{N<IVAHMA6aUkob&gziAF3<$^^dU+]2@3<qD6nx%XH.$P&Q,K\0rafpz`AA	r|t
d[2HiMiLq^ax<&:a: