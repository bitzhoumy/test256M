r%v"hdQ
#GLiC{DDNcqMg1eU}>QQsqn#P@|TV pZa5[\mG!
WP&c/A7W60x";izw&%!5frB`L~Ha:zpfU`>I29ldo%=/=ACS@NIk?mQb(v^j3ho! Al"wM4yxJ#6M*\CWX}_"xI~9t;m*4jj\SdH"]0hxNZg'L]b-}[s9,H*!+2$;k23!<8+
8)3KKN&x`n}VA/T1t%V(CE5{Yhsx2F1YCJz@p}%W4}	!\6x!V*2-bG=1ys/&f;FDKRf4`=dp{/=R%b9QN
o0`226UcU2MLvSq(gs5\r[)kD.tm\\'`1_<~x@{LK%Lljio(v_W\wZc::NKt`NA0Hb*dh22Og9%]V(5a	$KI)$f?/1%?h|IP^>65Ti%
4~7W*3b+k)gE
8FBT=OVv'/{3$sxaT	zIKU*[\{/6cKqP}@mK{zOi
j(>+J1;#b]Tb:xU .|#I72]]3-cCq-]!@^^Q{H.7xiBj/tY8/_wcBYijFWZH	+YI2+3uZpnKHJNt'__>cA[Ah!By]e5:Nt@ctsRS=\;mOcVH),.h9MW#dgF>C6]uySpPzm;uHviE2IQ,0:X(D;yyC<,Fs+mtU*R|_tS]Tl^$+n&u.}
6|pnU+p}ALEQZ*4$k
u+/mB([x\2b*cb~nZimOY6RYsL	d]*O{{O@ApG-gHNg(lB7xUgZ&v}=Nbt	Ay\I>Vh/xiG-z=OzyhA\2UnR/Va2HfwH<^\se	pMG$XfHtR
,<eI]
~!)O9W-^$<0gV!pDpHZSH"V/JN:z)fnnUA]To|5	;)o_M-	)}'j+1l3*<\0+_eQ12GmzWRYkn&!bakS.$0VByT.)#D_+IV;I9}8.0tt 	p:iPQG@N/]upp?{!$#OO07b;kk,Q\xA4,<TRA(F1]iS}.x-*D`g}ce[yj\QW}S<M8/A))`H-20uPefAQ-4p*O:>Go-/xUZi_:cxEG'#w)1Hq,9(e6&Ci)`-n/4H0>U?OE
w*9[kzI&f#_po*"j-pR6qJQp2$./mMMHZcn/87+()^Yus)^K-	;P-gccA<\>"^dq>\<AXXL7.g/^30Cq=Ek/LA:H6!i%(?C3_}8uu411[YgZYfz'UEq#>u*z9&Wg.B)x0N!PD25{tZB9fY&(p$u>'#[\6<PH}V, )xA8U59Z.2YaO\~1\M2~.`]QR-$KX@xW7D1oP/X'Q
ed6#*y-dsFt3\xAQs,hb37AE8}k@:+s6VVp1s4)0&.)F]X"O2J;eDJj51:K[	XNTK!a2Fl1v~8*"R7dANA9Gsrrx_%P2v80k]{I]h|jS;&LU6xm!U2)x_m<'P!\IH?]f;@;}19 t
Vo[<mhS#-,^IzM&y>V@;7))Q#ITKl%ZE[^S-Bl"B(>z,qjjku:QZ_XoaswU%j~Mg=Bkpt#Suyd-O@Pn0khJ1~?zIa0
J'erQT
FTC3z}RTI=Fx`!Kt>vU1=Dp*~;"R+wq<A~8.9gJT];^xw]`i<n@	%WGsl2c+%"Gz|y&<`2^g`RBFgiej1 7d;Z
bFriP0in;zG1S@AILr7_fD|:|0]g=3gM;s7.5P7!3!JED%,?"Dw/lHxr]Ky%hj2 7Yy2P'9,L'0kjN%0Wnpe	=(~6PgY|1VcG)iW4"g	CRth4S4#\M.28+i[N/WnDvR4cNG4`VTo<=>:3VS%	!'_'UjkA33S^'fEc'&*XD] H/RLrMdRS5])1dwf%7vqS`)}V#cwcw5b|`
$_r6 );U]9v{bj~TVV4PJQ9qFJR EUtZ.x\]r;E(]2ziR#4yrDOL5?|D+N_/d!mYnBI}@/JI!ZVE>=JQRLV{oZq	
UTVL1dGnTsr{%(Sdij^FO^E$SWRL19Qa]SG/"^m+SxsUF}fHd6c,'Is
qNoylLaT~''%9^FC'VMZUK0i/,Go(`z!Qb.i&t9(QXQ\nEe
gqdS7	a{NR2q%S^xqh1Bj0%A%XuX],.
,v-TQNu}{WgB@s	q^o[j?: c"&&QCnz_}BY;iPm6s_"~n[n??D>
S]ted:6|1'I;A5w_Gn@}9+S~JZe8bSW[Kev-7iS7N(_qFVNyC\qrmV
[=@f<.6,5cj>t^%q*d
U!>TTTmQ(^^${dt#L
2^V*^>_SRI<ruYGrW"^WJfl|Z1b@"Hqq=_t4sh;Xh^l_jN^^/jmBl.#vo(lq,-KrTyTY,m6#]yb	;#Udu<Mk#).)!tA,R',^?{O-5Ldc2eUeMVVPpA0]+@*~nuo4rhJ-A]'SJO2 (*84?fiq@*Lgc_Rf&3e.
lQC'M<1`8q.9p:dt3]!2=[/`C<#(No%IDs5_CXcZNU$LE
J
(?o=K!vNyrV,e\1~f,W^o\|Q,ljQTPFq&jaIV4@6HRN>",fI(D@.d>p6&lXQpF(yf+$3yKFMb4HFC-e]U
&}n[OWZ6[?0{R#w6)Ka()U\(mO4J>dGkUrF'tO2e<ea;1P,b,l#W&KZ:STO8M0yf[IS`uE3S'MpSsN;wdh!)2XMtk3\+y=9'JJf eoFX,jm.Y`pg]iDVo%G$IF/7/tM_?%}hFNd+}4Yja7B:-N#\"1EcF6 \Egf$,K5KQwDH_c~Gvjzf_[TF5b	3QvcOS"mTw^,qZZ`vG	/+M^1V6;e0;gTv /{li%`$B3J98]Ghg|&XTWG\sPD@k$ikBd&N=mg#d9lI3<Y^,|rtlPp!RB>F1b;9,sEbit.ee(S}oZ)kKFdF4t=`\F
2GT9Uhw5udUNi7Lx*/6(	!^Xq]d-!&..B+x(2-!^X0yFs9Wl%/`nV)<w7&-q)l@+.&m4GZn(b(A>([VZ!S^_H}26A}rv4J`dxo#@O^kL6zo#k/OAXmK
-7,fGBbg&>LeskL;H$^5SD>9yq]7*m;a&Ygjryd;c8FVD/q%H0e@ }@5Bay7}{:"FD]LIe^NZ_]M4{0x|4{^!q'Hv$f&6]bInu9Q<o-0U+ZH=w9V?(w'
I*R4j (ON1dqdo(e7]3eSV1I"aZeZd7Ls2mz*PI:g	+AK|lIW$jyd'6et*"8VJ%ip+g
Kv?\R3ksG^<wuxGDfK8qB=Rsjex5"7&u<a'>h1?<k6W0:7|<&?uFJnqW#\hPa/!qnJd=K~pcF`fsP+7o<J^[5;\i}m6(C,S[NB5#1b{)FY2>D|,O8S?8K3@eecx:}Z{1"Z&kpy1oM'Y;KK::_0<qlas)}6LFdY|!9p_57O]AWjSHi	h$nu#;yjGWd1Y<vm3= $'rDsF0qQZ6&w8PiNzBm%PTr[?76"6	(U7Zx
&x6'tYexJ(i5ev#`!8*[}iS_ Axc:^/ZKz
O%b(A^;<n*d_6!mDei{?9w4N^H+Q=G2['Y+O@b_k'y&=cd>{NcI_61{}U8$:	|9`|7	mD?84lo'-lI,dI>3x|7~l:;
/oakW]@wMD;Nn^owjTY,Gc~,L.fyQQZm5$uy!9$KTLL#4wi/@N'"RF_|)6^2OQ<Qx/|Y(@E'p^@f7lkNnKwEji(M3|GLX+\|Va&1V q#cnHKTqcx&0Sx5:aG}r>*[Z/XK-ig27-7MonErRvciiqc%^"w/Cx,]7j|"z9W}@"z	gXhSz,FB7r+^C@t4l:l\k/A"E5WYQ\n2
{4
N<Bqj/sQfJSl9(NEQpt-b#x-C}|I0.r)9;zC"lN2|E|;E(DBN:^d]Rl]Q1!Dn!Svu .S&}i@^uCA$1	,zQn1fhx0SKT&n('zDHD-i,Zbk;PO5/J8Z- jE}!{U5M*Xi8gSn59y-t.xe0C_'}*w_sa !cypD9eJ)}:Kl+C(Igfw3'5K=J	dQ-_u@YA&!no8v:iOC$f/HzUNP;T^PsAtsL1D[[6S*_DzXSm:jYYqheFwznS___e|k&iHykFZY]-jgm
N_,N61]])$,Y><>.*cv>Q|L6ZPmaaLS)4c@&)+n"7~4;xQKnT9[=Tc<rMN.c.#S>Y[Gw	BAu#;'yz$T]1"r>Y`=t_pV"%F%c/vL;:o0:Z 8z5CZwoHl[M4a8cv	flBK|&yuW:ss)G>}|0MV#ZhvjVv%-}{%*7UHpq;[K]?lrDz2P,O{bk,ip.!/Hp.$833(a
~3\ZBw0aG!AkE4	 NiqriE2&[mY[.(lI|"-*v2"s$2Qvo27
khj>`H#6DI3it:uP~a{RkVI'v
1Vy#5#S#xlMz.vhMGUsuYH1K_~FY]%gVER]E)%V?u:H&kv=}Zzb`u!J_I<`DJ^T3c*pX)CP19iur=dS5JiC1hJ`A^{g]?*W:8\\s=y5 Lk#J?<5rEq^+IR-M
o< clsT_]EL@o}R=L;Iq|9d4)W+)#D#m4?Rv:|Tpkboc(LhHxT9@WR8fj7nwVq[-r@UO*ZvC>S(Q`R}l++jNIr&df/qDISEh]>2$b9 1~?Zk6-$/p>K=??]m(!,.$7.c""~[gH)3;R7R~p(i'&0MO *LnpJ=Qea")iQe:aN/O4Yo4cVA]cGlOz&Hu:m#]_t_	3PA^Lh38.97&
vCFv+>'y5-/],e~[8wopYL8o(+%8VUcEJCg;4gfe	~OK;WQ1=`F7sT Q6&M14RwMC?b_Dc,g!_ =\pl1L*V/M:qW4kf
Z00Hr+rg|5m~|tY^T\Q1~+U%AE(75	4,MDI?1"-5
	}k_8)fdjIoI'Y	1aWPy'o!s CpzZ?|oX:c+R#oFIe7UDquvj4"\'xma.~J#4[pU9=X3W!pMK24<u|v}h:aG	OoSeMMEoDWFGDiUZCY4AS]JRr'1wpPZ>.;9RKPNpIydFN`
$?Cp/[Mw)5{o%ZK
bT5A,MeM="<A4h/]]/PzX7<XI*;	J8RNxk"T_o5{.hk{F4Q|TKlZB*lra-V
BWI/u*M%gRmR98DEo{Nt/#bTNxFhJEs$WYdkV".5Mkr1E)W	(ih{/Ou$1)VgePUaKNHgIEapY4$QI::A/tkbAArn\N'iuq_z[wg&QH	a)&ybpok$CVI#2~#Nn['
~N2Z[gs
87b~$A4Nk6#Gm$p?3Vp"!w|lr4Ntd~c#u[>3Sc"	O2dcOV[4KeS/:0tGmbe`vyZ<uj4'>QgFQ '`SH/8X[
3eq|8Z|ZmWVe7tiVz(oq&dN.cA}N`%jv}y.z5Ip5w0ruV3ksz.2d`6Zp0tm9$Pq=vk6N#XMH"1*@XJ=`*%jd:<o=(h4e"1EgSAw<Y`3+j>he[	`TVLw&OmP+_OP3-(u7jr9U^gWDs/3"+8s'8%=["	PIT/Q@4Oms,^xYE^+\`q:a9MVraNk*YG&C[h2Ov\&&TH~q^	jHOrO*@<i~$bxx&Y&#,1LY<+#	;2=g&A+HrI]0>(c
DyEW1ec&_7[y--CxkpbD[Dth{&Y
8>r}sbY
EL	<9#D(bi=Q0(VTTj2^yxuvJRB&v_A%#Q+LuGWIe$qJIrCtt!7s7:EqZ-w&lTMl1cFj}A+?9-%k>fqE[!?hRxuqjup}.C/{j8OS|!|,_%t}4pLn}i67tj=61!iur{b~Pf,1p	Snc
<3?K1?Rr$'JBh)M3}xDe4.pS*R6ZP%*(Z:U[|`[T3O?pQdQu8##.\7+'IenJk6SG&?@hJ0_Vqi_B2uPV:GqSAsX&>~!H!SJ5W1U]8>^~G@	u{x8 D{sva; /D!YmkTjf|}|RMA2*!"
,/z$]`Y$E#?lq4+iTr?PIUOmvt9A`AiXs8V](3^')Z]b>cq.W%")T%X<Q\.[Fm V!_3GgEN9fL\lH,=#9]i<*@j[lhhrtcZd4F[N*/s:4 	vuUF-[9"UQ4n|lA2W$:{J6h:tdr#2`/z.6wJX^T(&ZZs$P\b7^%YG,Q8K  T|aIY2Cv:`W9yR2H{QQ_Sm<4=j.T-}	$B]SfT,`~#^-~!AwOz<\e7;#b7ZDCZ|:fSt6(pO_F
}W;z=5tv?h6P7L0UnD;'Y?wk=({m5*,$Q
4Gvp,-|[51BYsSgI(vyVq;J8&M.0^g~2cC+EJC_n=xtmXg]$39;av%\EEeW8F9dC^~5>l*s4[kG6]~5"[j^aI@?O(AB=Ci,`[w<i'Plwn xV78W\(td|t9L2y#O2I'My/}5E7h1x d+Os'pp)w^L0&Z6Hxuak[^%UM8v0w@XN%4Jrd;SNX,N[d_0pL)JQv=M{ACdcw`AP`@,l&ZE7L=?h,hxOZKt,r;{7R
q|To\ZH*E9WqYmfo:8C$\gn2e|"=GO,Rh{0C:'Wa7G`ua(.'R\po.>PuU*kGRz&5gS4Fi\_!jith_]zNb${*0 6"On3stsv1l$#cp7stWd;)u_lB[^wIRAkL87vr(D1~@y@"'AVQYbq`mN{!f-_*j2YXc_n1u'JmwtXIdU`58F
^&V0WCAkGr?xY^tT7;Iq04L,p[b=7u}Ktvy6j0~]2\b?#5TX9txOIv5B4^lO1xZ
Kk?MP].2pQ*]3HuY/s2H?rTZ&0\\J8RrQJ1I-E1'mLpqf[85T9_:;iL"ah@jhZ8Vf~o|+}T~pw9LXCueO{]gyVs7`v|s*unb9B H;~rT2ckeH}O|p7t4bPR#x)9\wN6@:(m6+t_tiQ)5vPRsCKG:QFp,EQ&Z6[=
F^Vd.lI${T^g`j2}zjp .SR	.4EaWYm!n:c-3-NQAMQsc1$.])6ZJ$%sPwC`ZqZS\O{zda|0e!7S{G^}R"u3m@oDD&wK[Xp;]dlADlKamoP.,MnzZom|[d_Ez5J3EDrzRV7q\j85T_9TmTVDlbUG8>&v];!c6oU*='H1]1?Z1<&;pFE4K7SW
&R[7/gW]Kq&YN<]Ud!JVh4Y{LWVcc|^UDKOMn[[W9SX;EpyC{IXLAp	F#jM8^15W8~w4+]PL:D0;EU)6e^nH11]m3=q
W.r:k4ugpzCTh^)pa0s{DJ<&9E9d:5U!= l}"0Qd(=Vc0iHFcEt9~ks3,b<>zz2N:NYTLs
9nPbdxT	T,G5	7fE)JZ{p
i-5
Qd\!TW=
P:	QWLd|/Wn	7|Kjwkg>7F1'mI%rrYk	V+xv@|(QGuLB|(nbs7P/q`Pt	peRCH-JW/QAs~"m'_Yj}
-\t5LZFbenuNEG(J1/
I a*q1>5@jI1gP5n	BgtWL|Q'9>L_9hh/j5n(mowNe"KF
8RR>Jv
cf7%lI:/*fikl},]}=:cls/^J.5/Tru,K7g)y}P=~)k$x)(<tzk1le~#=/L&mrJ5gM6wqWlirczq@QS<s	a1I}DM1y5[U-`6q	u0?fHTLR 3F22	AT l;4PX@5(m%o2rK90VbI3h-wL9"t`nXA\dt1[%ZqURLyW!f\>d&lH$.^zsH$)eV`4(tez\+0~V&d	]]ykX^V&zQN>-~ =7F>g<jKPbX>I-5iTO;kKm,|n'6|D!Ds	)H^CSPBpN+']g62BbpU'E/7^1|l"}SPrdc1xI4x*=Xl2L+E<f/zWiz[/bRUdc:	pKPy1itMdsZm	Mnm/g"[2B}4`\P1=[-nP<k,J-!/xTyAkf.rk{8Csy6WV]wiRP
jqwS?	K/]*uBj*9p1jU5J*A<^-n<@i#EG_m>MH8b7}^MW#0Ih=!*Sfs!}q7|	?=[3W!4c/cRs,J"n^N1G%fC]fKragghCqj0LS$k	wmc~/)Io!Gv<rKiB8nsV2Iobzbym
!J^SR9%rgPc;wiV0}tmNi%)MB+sF<ST/["Ho*aw[/$jS.7tnfkUJv?7RbF)vX=KCMFQ+Ax<j%8r)3+qW3[11G2=
8hzY#`NC"X*:#p.z{+N:hQHtm1;+pCNTh+M~sG'2zhr<LP8{x?KF-$19M{4p N`L0FLWz'?res!Q?GW!G	iA'[(Uf2F@T7suckVg*u:<l<ROk2I2hB5*H@_?]- E~X}\]	]4>^+?3_dKk{b<06BMiZzRY)#EP
9YPi0`~
LL2,|_MU_)s6{G75B,!"<5cbt7>#hxWl" R(?uw_xu)eo2-?UIR1yPt" E>dRhab@NH;RVA8{)a1}(DtX
H5tEPg%=,BM<B)fUNou'Vg\-A9]k0\R79]PFYX9cUR{2#OvoF\{J$Y-`U	'srk5@1cK%\IBPqRsQId7wrW&ChU~.<jz3uxNvSr4H/Dj8;e
VM5n5EvS2FkeF. 00dP	0P!Er36yM=P=*vgXIiFk:^j/#NUJ(]RwBu 5`0_+FE&U2uw?ZJYA2&4pAt!*
&+63RL4MBM*-kB,WtX'1'Bwks>Z4|v=:r\	ic>@B(T(?RK{x/t*d`vrWm!=|cc-PoH;.,KGHz+
}g{`> a'=;7sbi\!
=DvG#4n
^?\kWM8M(wH=Ce}34{D+9uLU=2pB)KX,qmYVoELrPJSYl?bU$"v,	BQ4v])8bhfriD_v+RwT(4.'cdJR!mh\s"3Uq^y"deu-kvxhn=U>w4]2:8M`5=[|Ra5 )gF,klrj<^(cN!vr9H.SSbtc3\TXefU)ss@XhE]8R(^c~Pdp^F[<AN+1$6L.VGhXm#`Lw!@WSYpLhAh<4oZ{Sq(dJ8ZNz|382or+5is4s_%wgf?#T)Ssfo}_}b_@aS-W:4BV2{>q*[rMUo!eLP#s=`9&`6x-/}}D4)0VD%#kVd>$2>Q?AoUv<}[FH`$iX{xXNy!P"*E1&qY5Rv4oNCi\N4G`~]$3hHb0
Kx7[ty2;JfM;2qRcCP4uRrwhY|g'd=yXp	09VgnAs%#n:4>{FvP$B8VN,;}-pxQBdH1UeaL7J%|bMSJBF"T93[=V{6ev'*h4KQ<l39|6|O&hoRj\'uO)apn~mL+6g]MD`8c5/P\V:I+.t3xyWpD5y=cxklk*.OTj7-VUSgz;[~m^(lZI\J],V)b~vTFx{7O:%.ig%8r1lv- ySSb1sS_
&11I7uq7*a3<)dE;j+Wyoq}`|r7l7iP9<X!*#[]?Z5CfxPki_?W!_iT>)Ka<.l&'pX8wJ._Ub|xAp~!;;t<i$2gt95*RL%091@%x+G"y8=_q%qPLM'nBn
48~Z6NJfJX(]HqCaKE1J<C38&ZW1]a.p'V]/w^*~oCk[2.:.7M-iq.edGz~O*qFVdH)(%1mO_=B[1)	d?a6DY4h[*c/{%xT|%X[wPP,+ILrk`"S`	{I7^]dY,1CTY.}*~o\{uBzmC}YvHTbm|r#CC?3h4it+3:.$cl<S]DpPSg7
p$isTh'jYvfNO0[]h+G)'z{7\8+5C(8K"P&/lzF]JF
Tt4~#Ds%@)[Z#&fOcH:-9^^#syT'ioEetMo2W{1c_6!/Qo0ZKb&`l9pl15u1>HYRB"aL
S|$a|jM!(=yL	1}C] 6/y[5xOImj*")@jA\WV?y'#i7$kzKO5;8T"."'"[:q}!<ary$mB%4\7]#RoS]cw{gF,d[@X/L\<$*g#f;8klB"rnK_$%S2B^E\C*T5Iyl@YA)/?&fw}|S;RODG6+(_<vsL$t`I1Qd?b)3W[<Qg3I
Ga3%Q=xwfT!_#QsK6nyVEPen*0? uAi/*z+P,^fq6]:,xpPvG~X3`(Zj8jN4U,EdODwhIl#979-;%,b9l}E9C| )5
E$D<4a5hX?}t:t:xKKxXRM|4E9:!Bg=3_0-oHtw5@*	I1.V|n>NziG9Iup_B^c8'59"56LEF$Ig5k$moitG|61eA=m`_$V9Fu9&3q9e`	5?AD!An54W53Cv~Q
%(?kG'%kYL$"<>G=T"i+C:[L>?H0^%4}&^z'?ye!63K7I9s}0G8%sboJbR4_,n@[-3Rf|:4oP6Ou+Y|MVD%M&2@2*$	;*cA[->0;p<Le-jC,Y-.O^LO]V-{
D&4z4pJAWBfEDG5@#@'I,H#Fy~M+`uZu	^^H}qv8K,79*Rvyz j5aAD>I"%L3=b	xdX4;vrnXP8:K~@r6-D(pkX|5S?~[HimqJ~O6AbT
7DkG)J>JZ_4/G DVu^01H}T<~9Ya@BXu5	i-"9,I1pXz9i%U_Kz%w`jOb=Mq&D8?fG'f3Z!7Qi-Vmnx9j|({\]<^6M_h\|2tRGf&*XY=U^iv_K%K.J6p96#0'iWN]am5rDY%'I@D0He>M#PRd5/p)(T!tF'JE2<"2xb<orTbLJ
cC@yG+]GC?67:;3)L%L
^`a0D^!Rg%2n~-v<I}a[)'2j1;xHSF^Fv5N"Vr)B3hU.l`|HPxF.l7Z+[i+0BUeVYe
gm>UCmIvlG4O
NWlih8t|Q&c5X=	}EjCzi[	w=qEXg"(/-@;1[ede<af`=U^7X@):BLjix&@e{z)qF!eC}c35HO'R_sr!	HY+fz[$$@8-m8,x#^'z0A{6b!NyHfI\tGgd8htp2)`"-	?M}&X9xSje?WWAp"U%K?mg(h3	Y6%0h/QX>
|@`@`?F(odK|'uGt(|m`^0KV?9l< ~CDso`M?^>;[$i?-kb@L&z_FW2WM)}Kn";1;j1RF*d5AsQN(UvfjpMCoDG~1Ngo$fepRr&fIV?}j,FG'1=LR-M3m=DFyn!6wUT	;JT->Ik+L>FfiOvZG@7HAlY5\"fLM@ RnTu	?Z`P;=v__fL5~>@N*D2_nf]9f@i7WY@"tQs%,/WF(@wN8k'uKU
d(aOe1o9#s>(Q/'yxH+~j[}=yQqC S-8
7[RUM-NZd_	Fh5*V[R/e4WJDehD\R;
pR6yfIk[$ )oC[f$'\3G(-g	uBRZ8uezi>Je#wLmR%7SO>:6=t%!Q8G+B<1f4DT`5&0.fIJshzbtCVH{W*R'"rfS>zBMCOykq^S`55_b^>cm}^i'@9Qp]M"^Nh@64V/^7E*B`aKZIC;$O~D	T4:)+JI<UxNBx	7++O"8pC])<24%ef%uCaH]5?|R-/![2)X5~xOF!$9[i7(Fj*@`5~QA^_j}N944\[f?wq5HQ^):P:r3R`|b9PwHjdr
^xllK&&;C?_=gi^3:~wD:D`cvZx"8Ccz'O
RFC9&QJkD-"_sg8IDw+{`hxfMK}+r8lx#!ZMub-Y{Z_124x(|[*>f=N$u<Wl:}an:PZ;	"5#H7xA#:yp
|nt%jWG`t<21iKPiBr)5K"a~K%mN3ngh%VaC	7%M<&<##J$p`<M:lbr}Mn\!SIVb7yc`l}%T@@'m+hT*[A0[ SQ)vZ@jN1ARat8C.UWuSGOOPE_s#<at
z\
9X~s&"O.LT*FwY'W[\O4'd"]cROxJJCxqV 7,:g4WJFxCY[Z*Emvs|4+\&0X}gKd;^wgl,Cu{r|Vei3+y=`eoF'2$.W63gHJre4f`=lP!XL6t[Va-^mg%MM,ErTX(sCgB})\"[hFMU#(B1P(EO{*+q#YE.Y^5-#,sC6#11n8pDnfA+pF``EcT]x$=)#|T 52saXjdUQi)NYLDi$s&A>'&QgPe05A!M+90'l%"-eWFZ sja=9duShRK~'n#jG[Tvq(>g1+/I^2UFUnmv>au#P[HdXG?DLC*M\"iU`L]p^H<.m|tVRs|;)B>h6>mX+Y~_BP?@z`:L|F!pE=?)CG2e2>gj?^DFFV+s"-%	R"zjCENNhLrn`'yxWb]UK+pk5AD_#_ys& 	/Y0NV{4?!lU$Mqkw]bZ@=S5-}u;PnNw9Gq/}:_b`0+2GMk4[$F|3S2|I]0C@I'Vl1V@BzpqR>]1wN^=U9f_4dwN
b2
ueWlW9[|S2iH35Ok!H&:
ux&oah	POT4!ee@:2`VMt[8,pV/@61zN|(*ylxM$%GL2.a=%{fak4+QWk|2 %`r>R-PW VmAQ-Lo\308a.##*KpS).`\@|n`DUD-q'W-(lpZ9q!6$euOu]{Hsb?jT:K+{z])s#J-eg4UF_~V^:nro}2~8lfctLE3sL6lU'LK[R55yf4,Ix~n%E/9&ih^V{xuwA{MiW94'Za	lFu+^0[Zx6!h<~/&--;Sf/F5}sKlUJKr!y@|@sK{57[lK*lNUd^}TyS{,_\{p6]ZC{2,U1MO)dEHP \7k_yN@WV:?s|$|F5:pLqZOQ0^G[>`kwy;+ITtge{I>l*O<SSPxpF4'|7HeWWIe(7be"i>BV7A#ZcifUR.K-;eeLUj::#D$m7zO_-D@cL:kH$|+_0HB$'QM~A
s/;w4+6crI1o'Gk}aiY-a,oknW+}89G<:*9WKC#-VUF,0eyMGF;K& tLe4Yh<6(u`407jFR^sVCVlr<2t<]VxeK-Q-Qf2QtYqh;{|	Lw`nhv
5d1=4f7NZ\'P3wp3;2.\b#9D~1'0ta+ ]lzW^8gX3hWx|QOhG7"Q^f<.jIu{7rkKdfS	2z9B&menMkom<P|,(T~kY\i&5H?u8fEw"[_msJ]:})[wDjH[$0==R&)/k9 )-\saK$J
>f)KN&w vZ<w;$Dvq862b,[I<ngaL/lqU>mgh`vw/(XLzXd|%EASbg;9b/0^o*(%z53`f'MM2!=nb0R|w%%J"~4=48`G?BHHim6S1MRyxF6P}z/el|qo_G)HIhdVOfs7$$lFG!?=H?k0{9>8~:g^3/}9&_f~.O>!W-;dxwZ?5PzP.A4Z>R4XIjzL{rhoj.^~hcfN7,,c(aCE[7#7C{8#g:x([4B-fjiY3ne!/<5Pc2o%\9i^q
>G\jAj|:V=7t0dpLKgeb4RTHd\R'tR?CZ`{Sg$@IHbwVxsr-$s/ieF]"O`47).3GADJ0pS] :\wuR1s$+{F.lxA\2SN1hVFsc'#1SbNFCtU8I_["@BH#+MEy{@6Y_'#>YKKc5$BCE\]vfs\
0VHvEHxo649SL9&2dCBY$$YZ|WJ-I,,[24;iK>T^p6nf]TA~i^RA
JU:9H5qiI<QBi1:1;$GexBw<@5-HsbK6Z2IC-.Y-]>:"KLag4KqB[PUsUJ^@0._OOd,[y&.'j$k<1RHxC
y#%.S/Q?9h^zEDE|J/I$ubM;9	6^KwZ-]X80+Xr=j9j,5}3{{}0JK[g!sHJ;(q{!E=	vddo7m%._FEcb7@"y	~3#GXvNKq#0/np%Y/ocM,&UdYh\\b4,ii#1>QPWRj&KfsuL T7'js)oHLUD1}R.=XI_"%ETULxsQ|s9^j!z;Ms-qk3g,#c8v[QXE[':)t$Xs^2E[|KR".jx+y
B=91Sn#0B{S-)gaNNNSH"fLyKa]D;5i03T=M#w`F0aEZv{{\n@wZkBa'UKs\<Wbrgol9XNfP~9a$O8PcQAEpQxTI^$hr#}o&Vk^P<w()G?l}=?Rd,7bT+1B|t3~F:r'Cp[*TSj$Oe]4'TC6:6z%v6.J.9fdGxLbXXQ;/Po~OK	c]<q`3Z`ar(;5kev|0ugfE'6A,r_zbAN2&xZl6fykpts'1[VMrqK#}L/.5b	)`GZLiZ`7H?OO;f"o/NgT4$iQZSwD,%tL5gLB6$|TO,8m-}9SiG\0i~)XdOfESQ;TikEL1F'D`U/aRT{\qR%!Zv`s:m	3*g=yDzB>,716GT&MBXg$[(Z0E)XE
o8nPaDp@{^1^!sUSF<"D`q+O[K|]w>Acj]S|01<%{bi
}kG!^{a<k)\@]W7;#HCz7EG-S#9Xtsz`/k}d/G~CKx#QHX8Z,f9"?Ytt\@h!:0s58C^r@b+&w`8};
_kf8\dr^vjv8XcBc`21AX`]P|j7mqD#>|i|rZhI>G{WbMx -b&*4isZ5[Qc34'o%Sb0XkR[sLETz:hT{I`
pIwi.+4LR'7G{Q$\YiUD-|tZ zp/VbxYo0e{\P67073=(jKa-?%i"kutcyfE`X1VOxc3<m* {-G}0*K+5e}]kG`c!YZB2_t+]*6g,w:g00W^dr?BRy`1fC
9<lH^D}P`xl,8OHx^Ba& XbO]PK7'@m/pI!Gi%L0xit]"Z1u+#X1~XP\+Tio^
|.	6bMWI#QjmNJ	9rE>bS^?1huz4MP;_r5B<11^t[;MvbCBWQE@?K6J&x{2	XOj,${ZLB7`@'Pa\x@7`sif{=7OxWHgX#,1^pHrngNr/v;h71Fppq/aw/l[Dtnp ;lhcZP"NL/q-S5>TV)zRIs_y?%QqPUA:7Ux
!-sBe;P4aPV1<;2Ee]kXLh^>9hjoSS?jIKWzh|Fr& IKBfYo*Aa"%yLTia_~v>
ze.-{"B{R#9-0P_LI@tqRqF&YMejaHRu,gO$3M~ ^0x`>mjt='0F?/R(&5qq#bmPy]6f>2H%vBgX[a_f1q{Q8

cbwK;+1{lh|7%wFJ_WX?kUnbsZ;1ZIgTaF9XZNQ.V5qqsM`}]7bus nGz4:03D>8yLPDa70]qO{$O"N@3#xlYEc)~18	Y{,)rnK*>&lPCvIMO]!'%9Jy70t0$"qpMIg!?)p=EJ7
mr@8U_;m6({I{B"?~LwT)xzsX.RmX} #os-4GVg\9+Afuh.o@7`m%=#l%VBG?IX)9Ls}%T9G%JQkPHWO%Sg,~I1E+2/_~<(tKq=3SS>c?yiY$KdF>%A1yi=='3z(@7ouZGr4g1}^Kp8O!]Pp`#[R3+rE7QzIV]I23TE)'e%\gaemN~!13I0Uf(Ym{>nCi4
vUU.dO4S=3R_=w|4_T"{K]:glm&/&xho;=hxX	TB/w3iI9*YnB?d#*!]*)g7F-EoX[hf}ddfbL*D[UVx
Zn,s*Ll(p;8\yiJVioP[ 1Xza{-	\9Vyxnr NtMA!5",&b 2Qj([elj[sI,+;<Xwp)SpwKTgOqUGCG(c%:g!~U:Nj-T`;NUE]@{v9ysO-C
Mm9s	S70+"[h{zjLR^&gyUNV5,dKv/py|):>)rx4EK~`tG^0p\$YeP64V]u3>$!~Q)J[D\Ys:u	|O	Z9h3)"V4;;#&thX/5hQOR`jjp^D)$WM6Hb,\L<ob743)m"(K2O>|fvi+d{^$!D)+rvK0.-;4:a$l/m#UXt=g*|6=@dfPQ!n%l<'SQ*T#63gw5W56e!+KI;S!7cCo%0WqdOkeua|
JPoHwpjH" 6(^.|@k&wybYe6MF#9]~?$oGw)A5RW3s?+ICHZ
Wta&NC""5t(A:\Sd<`t94c`fTv=1.8]`'|")q~Q>uY[j#vx!5V	j,dxjqOh8N2xXlyGsf&cvb3fH|1TtV._MMQH:6QFH0!R4VP"sRS)*zlh>_H+iDDY{?1T)cB{<b^&:]Y^DUWBK{2^%0Z~ba$*Z?jXsb^wUC(q?q9dlWd[uzF8#P;2*d	~nu~OeX^U>WuXF]5%h7&LP|t4X0pgXAhvo3fJ]yDO]Qz[p5cV<L=N<P'~#w@ ,m*hDPH&vCy{;\L&P^26'JIevG> ju$$zzLj*B4:+]k3
3#-ZS+}`m$OG>RTs:i3lq,,u7O/mrGig  ^o3l%[+UMvXpm|k[~?H5=X{mGG+]/^ydYFQ`DUq{>QHjhhvOQ\>owbKv"|
LC%weh:1!wK U@,[\M;Xa$_2KZ@yL^$o*'f4ft(yZsP#Mo_`+"yFTDhDSg$mPz_akmPiO2WEm+9F|p:jwYv%q8UuuH^lRK%bEGjKN\|d6D}wM6mQ,uDu"QPUk)
u >akLAUd9yR/" s')%u5S&XM'r);0AKj
$[ni7j9$:EfWJ_T6lg9+oF8`qs\Harr
{I*-]6DlmeAJd
U U8.qF:zJ88VxQh^`pybVdAk@oiQWRG^H%c&]Y|.2.N!rwbYm98oZFwSd'(9Wg`;[5:LV7z%Vi	OSZrX3J7&vul9IFt.gn6R%sMBn/QATMcWF`#SiNJo 'v/)X5Ee?"sI^<{-)f_\YUfD$^B[8#yFUa]zI:jv)jqAC*!*vy70t:9[{tRNZ_N(H8"+mxkC@s5XQ@cWD5|otQ,l1kj$cM$=uh%KIIdX{1,lJ4q:0TnYr4;gVLD-oTS3d	(QgrS{&&9	aU6!y!((=A>Dj>*	ki93w0nJ4h3uF8q%WGV]sJ(R};r? btq[&/CA&*HP?f7woGXwx>HOCg/%T^0,0&|nr5.ft:!Jc;/;PXw),pnjqvD"","RsJ\2fS@65ma1YS/{FDv-6rXs?~^:6x!$""%m,`j(Sd|00RK6%>0Wp,`ow!Z?21e~R5d\v&R$L|mTT	O^IOH~d8T0:fj$ :T8Y-16HZ7Z:@x8Pn|oDdC&.!s9,&+!fBx\rX>fGL7mS5-l,Tx/~}R%N	|Ya7D)]tg0BH7Art\.Da Qa/( /$
jce
$H]P6$1$Gg)&W[Lm^lB"bHsDaRDtZ^5en\BQ:8w"cP{i&#q#11@=ED4%D$CKa>F)T*J#cKQVr~G'V{4pVH+b;n2J@]Js{0ZZ*b.]!xB;UO]Ely
WV1] ,:F$$3X4q~t(ZzgI?;>]F\3nR-x=`geF(3i1!lZH'AYi0"5}(MG1xTeGj/	gt7EAgk93DG%*h/	O2/b'K ~uqsO9bIt;ghCs4l_$Abe!-e8XVt[tN 4a;5A/VEFpcrOpUU4YH.bORS|hJ4q;`E~<cUn;50twsk)0w:|T.K
jc:3MGUtXtNj]/I.rq!g#kW{>UR/lh{F*'_GR`\Uuvkgt+E$Go~RfYMVXD"aBY-M:4cWrKyQah<AzdSU}:Ku-E6XT~jBGs2<Gnc@#uwQ0`a#D~RGpq%~hPi%POUgLS/cAJ86 dz}tv\*j)TVt@@mFP`d)yn+MinF6e}G7wkFNv&T	W=r)^X|RK3.;hx ,cK[vU[ FZZ;gQ^1E*]]LWE-HNd)q+}of4D}k=/XmtL6\qTbX7OIB^%Xd{g;k <w|#]+Pv{](i<DeGZ$n+?edBuq>9j*c>?(ReW}U(=F6H}fKy0um54p]%aCWZn*ZjLyVc!QjUC|x9+TA%8H\2V>[r}HA*+J
= QA-.xs([(1+e~EsclShzg>01D5\:N]):HY|Zl\RU0?tXhqw;nN^(JG6_pwCkxjK[z'HkDk,M0x"EFTHEhF$;z`Vy(Vf%KJIi[SKM/.gN<G.l=~P$r?YStvQhOb@'EfWY3#b'2	sykyrhen><{*qsoJ NePItc$eDprB(/\r-SANE<kmq`Wi'U<TuZ|43@5M=8[<'zr$cQE*n)P*YX_\GdDKV{7>3-^.Wy:ZB'Gye3pbUb/*DJeb/W|\P;{ Eu&hwEj`=6_2AL&Q6X<(FXc,jQFZ2G_b#]imeE*rx#FdC&,=hX6L_f=j+!3l\^e4<dd_F@ML"{\.$xovkJ`UV$:PV2<oOuHifdjxKwDd1SDtL3x7[q-AC0,jyZ^,
&aLX]=h*EW?K\=SX'(oOO,)GkWjrk[|Fp7b7^e8BQJO)UzW_evZe-?(S1)br[lrk0Jh_\$54=fo5.Eq%sV;`;ai/Oq[r)3FC}Z4qVa'?t=27'=D Q23S86p4kkOEk+BjE^GjQ0th-'=0M	,%5
_[%cAEwwn/+GtcN/?4|^on,m]\;	T,AI)P/Zt']'hgVlvYFq.ri*Yw1o;]>6Pz#5P>\&RT<=lskpV1m@%
Il]hD0$@d%RD{brtecyxTlFE|Ordiz8;<;%9nJd>A48!7caF037?TCH<5d?-prfR>V:t&F\C\2;cPCx EZaRNj"+`,xwOLs;^96)W="D!D {/;9F=1m4L
<m`G]COcDq[>lh?!VG{A10Mbel3qKeiM2~SS@`wI)BJ}'
+!_=.O3?N&3uTCH_,.uCQ_&4t>
0."S"x)l{6.)`},0q|5d,_#yPOyG72n+;]z3_ivf!xq9;~Rlq^$2|v2%mzoK9:V,)+\;yvXRlZ:A^i-R|WkGeACkp\~>bm6prR<fU
-rs_A)B!A!kF\+BBQB9faK1Mn>4{Hv,l[If+Df$7t0nSPC:dUO0k%&Mxl\c{FvEOJm
yM,U#hX'%qMyl:^85'fN?3'-30zj`iG`Lxz1Croa&685}vu{&.F|!X}d_xuUrPloI:yM6j}$.pQfu}Gbi%Eip:(gy,WnjMJH,EE&)v>6=MOc>zZWaB
jV+vUi5R
Sw:LJeG*AKK`nT;6:5! EsoHtw.xEcf$RkHyt:;dbehHyu=Xf?8fJb6q~K`_xS~)
@D.s8AUkWeM|"}v9b?]`xN:ACP>m|myK%'cfID
UNkFU a{C!5zVm|O9a_q^W+vT)c+hsH?k225dC. 7tJPbBgOoA(-o6js>%j!,|Ow8WNrt@7rv2s_-:'-Bg%`>[.RMkTc/&Wli.b.NFj+daDP	(J|\`u4
&=hm*r+*oGKw3AzTUx0v_a|JuloWh4{:a=oeF
#}x^n,@vkyu~i&y{Dnb;,<rMV\<gp^0op!#*9HMh>ff"R_xjPIF.dD vrmHMa~2Ue:"iSfTrJoJ!D>Bjf*upjt~N<-l2?8O&}v/_c1%#BD(=75G,_b%XpNCr"[~y3h.O	53GbciwZtPuiU7F=ym/?Y/z5.F;G[=o7vrM5-#Cb~]""%#y{\kuit9t	dw>LG[Ql/;%/$(4>":t9\4BbDkfuVSgT|]pPQXNO~8Fi<3pbKVvVBP`~L;3HsoS<O	d}FQ7E{ARlvk(1:A{W) !$dR:_yS`a\vo-M}BaPmt+g{Sj0/@7,<V,1

=xRtXD3~2>8cH`1X]vqo+_:2k,5@:m{?Vd!p|CBQ/,7 4!5KuOk>q&d4?u1immu|w3_$.ZeJV_oSS5zj{#HQdLkO}t^m[|!|S^=?*g3wNbwhBCXK\<()eDBlVny	T@0#[PPvpP$s"|-h'fX8&8rSbGWub<9*kN|=}D~}d.R8DC[?S?v:x>\3:1hjvYt	?	{@Vl;suz=_oPLq	qjtdx2(1}tWD9@
'Xj3`&Z j~YX<[FuPG-$A`G9:;>0}?.1Z(X|eqe @FyGe0UvNywXRn;Kb{D{UdPr7O;9d0?U;*Ukjh@Rg'XpI^4TXsw[9OOZ:/#}Ai{9&6Nn
5{D+IW#9-^I+WBcaK9Otk~*ThQKp6_d~'Z"xlYdd,_F>Uxlt!WsYX!<H;+|yQK56RS&GR/#KBX8>e]@5[|[FDd7FKn.+JqH}@xW\$YZZ7\=43"	-^N}.{Wn=fVGA":F:E:\/st\"E?);s8}Q<EGv4G*9Nd[zsm<cVhdYP*FhSggE
/pzh53&2,saJ/^^fn._E;\iG+BuSB8.}[?Dw$9]'dt`[u/eD	r3<4ZE4#DhrY8Fx<e]g"P`^SK|2q18X2@=pnBAb3?24.S;#T#{5*s)jZRXxg^\v'B'dyLx*ML\B*&kBJT5~WVo?@7lF8C`UHmA?C+2[.QhHRFCOq! gPZdrCh>6muOtY08>fq\a2[|ePK`N!^`\e}=6E!$!fc>HW6BW_scLNdgd9BX1:(pZ1Oosan>N_o-;i<,CHc
}w+&mU<#?Oo#f\|P:w@/v6;A?/)x5w%wdq}Ug$MoKu9)3e||>oodP1);,?nSIPexvrMG.tF>P4b:wpFU+hw4WmxXb(JO?&k5( riT"$d!gOE]MUElXVPK$~8}M@Ex@&h@__-(@#`u/@Fpfs2%xmGh3^\|9C|FaHT-XY^q%6_8za>>w=Rf.,.L?S]U":jlSiKl0J#}d7_7J+DG@xDa'(A@$WDan5n~^7UE$+oM9&$KOq!/>W^t$}Q!+7m*ye48j7UsD(R^+)(@yt/d"1y+NkDq[?j5}%:tGo.ZmwH7:1	[VnsdG(SJ(<bk|7*#dlz5<>T[e9oxe{]RCi0&(LC	}zL1UUFj38"J>?\u#la}SiMsMVJ9P0Y@Ka--A5;'pJ_O\	NcJ.vgczjnDPxM)/vu|,=dBMpIu	XGeqK=Tb9]1oohy6uG 8F|-wczPC+B@Ab2)<M;Q(S@4FqXBWD_e{	8$jOf\"gCqw9vJN&p\\^>99Rt-Dy} `3tU3E^G3Wh<i-T]IysO[w}%U+r(?Kq2f;e KMv
qM-g\`I@s_NjZyK}iviRAx3
jY6$UH{95]JZEFa4cT7-gB9&65b2xeF-C"6J5p7`-E2-Wu>Y)SDPcH*3cANCN1w4O MA[W\,V]w~]F8DPA]4Snm=FIGb6jQ|CF<$JU{h:Bte}1 "IUC]zJ<U5`V\xrQ,U{ViiJnrq8MLE`_-$GZd.mF.po>XWT($@1l4Ma2G)TA0p<[}uBCFk=yhDM7Bz0
\Zij+Sf'9G(J."lEl&xa gxN]!=>kKh]-LJi6:eH4$mZ_(7U{P-i<|Kq}h\3NE~J"hS@I3:9EfvqP{P::ltfSdE2T=D4
Ck_)l';X4y2k7RW38U$A)~p_|.x,@=:w]\kkpNXJD	]ehlk/v[+VP]ZWJ:jUW(Z&+lO|g.o!iw?TNmQo#}#'\ 7,jz\V|?@+Da9?d	r3e) [G_
*<="#Q('u_iLudN;T]	rK)IEH	ebL16~0#^H@26Yu G~/{.m:(3eh,lVR,OQY; J+dL(`@wOc
%F-Xn&cL#w@;52j>,Qy~=fH*hI3Ff.?er7D%SD{HO\O<UTP7i!i[ Y ]Sj#fX=m'\<nq@Ur]$+
=$e\UBsBwMsAZ's!hFz8yk{04=]#m``(.@0R]5.!B=wG2~+?Mf>J743HSpCV9>{"Me[x%.MitRu^>>\kU|x+g1I~(`''.32C{21.biie\!ju=Re0aX"oj^xoP.K]."yY_12: ;i}MJ,s5 JgRd'Z*G7*(;R=;$Zo1v!k&W_e[.,#{4X69'8.+X|FieY*zB}Y~;*m&`A%=BWWv>by,[|heX"FDnO>]28,%ML4G(;PM_{2	T~t_W95=|+h5gf5P,{}0r[*b;[SJ$IZE]kmo-VS2DPPj#] e^txVAt>lcG1k<Dm|im$]*;!%=Q&[]K^>5`%gP&9O}i?Rw~u]H%fp|.J}WM&dqV@<i:[A>eGrQM&Rh&Th,DR,dh ](31:|Q*iKZ6|cw>=3D8%f.(h%N6Cs40%=kVi33U63T"6Xu$}SVf2}T tePMu>JxUV@=u=e![LB?qGZbf
NRBN{2<sK5[ 1]\\w/4uNAuCjR?Lj8+4V}+.bm6y
:&(N`lGYLd4JuC;)}E$]/"B-pOL!G>L~FK13FkwO* I5 L#RAPH3*sRe}kD	G q\)Tl->ZMF2(sRrgw?<*lU6z4q0h)3C:fH2n8u)!iM/,1m!f-|lU?Jm%nu(Sn4}#p2UGh<b',C6vwR<:SOcZD@g/Ed#%?}~Z~_1K4
Ma,BqX#BB2^p>w-PpsgTM^BPWM?bo%)(40sv_.KheeYcPJt+$qY\/=>)%WW[8+#c2Yp\:b!;"FNNt=v~LWG?f\>iDjkFz*|/>B?k9GK/
9YbizZ EU^5	5Mt4076ls)FWk86v?@fZ%\wX&2UA`._
gM6%	qHB1W+#HMeqvG7itWtz31xK!nH`Pe2o01,V~=
nQ}	0r((~oFwO
(CJ)"hyEeOr8,>WeNi?xkN91&vl2/"oKzc38LmF
[qZ^%Z$q1ON@Z\bE|L&rF2G
\y&^@rn3H++1cr![+3%`46:Zzt7dg.uq> 'w^1Q_h][:p6\~S{$`tktU[3(CqtmAUZJ0sxdOSHOW=0	Dd70i`ps)|d=&BC9XLvk~nudcuwNjsl$2e5+vU~Th{?h?J$:W3=Tjv^?Lw~lAU2bRB"9wEEnCv@Y9l+O0#f.pqE;T/F8_y^!=E(Zi#)c
4Q2BLl_#YJ]BW%4dv2fNin^blM8QHE_Dn&b:I":X{e[8Oth}%`l]r(KMd%MbfJNzu\+0[D1@:@9eZI%|@V[MKxDwNNVt04B w/>'{jq~tKN/&Kn3-=kpbN$TtK;bh5|N\k^K_O5E[O
P:wSi3=}D][FL},,(~?[tiD^L=U;>Sfrr3\n9xmRDzApll0*KLR5{wXD}`k
*A)N>:8pdWYS$N"32X.P\BM	0w_?8MuMel4fh<8lTD5vM.sB}\5kPrqhQ!aMw6vU{\*-zn}|ND	!qBh_r=xM6PGy%?c$^u/d4fa,,rjj{;8)ww(0:67|X;)V0Te=?_!Xx`A4{FgP{wZWwdrr}X
,=3>"U1_O4oA+E{G$~?0KI|8	=^_JtrGB^lzykke9O*P
r]?*Kyu'-02F9'XEV	}..u=Ag( Dca9g*e$@k(-+Lxd\ZlF5.saW7/@H.Qr@Qa`U#$zG]P(<su!t=H
h1CCeOH/{r"*UQPF:_|3HyhH4aKVWJnoTg|ur6` {_Lnyy^:9C@8F"j.813T?ok[#IO|S\c~Z/Hq"-=wz>2>H?L4[&_f$B	E4z_,eBrYjBPXSvmyH7vXaDHV[}Y>RzTXhY|+3KC%i!)`Di	ghOi\(nOcC8JKj)hXi0mv\D-:_'Mq2:t!2y-^	ydk>-,KdT\SN6.Q~h'KM0c`_^?d
|eKq:),"-m#X$@M.L!FF5EO:S>-gkV2H_"~w$$s0*OpQrHeUJgEQ<*>BBHd8+Q{eP)Q~^x2>3WLh-?IWY'!iImy;-U],9!yDt:bek'DV)x]9"'w6norHP\)a5O)]|>HS^p!#ejI0n=R:z%oB5*g07n<g3J!'=]8K2HC;k>s$R#~5b:)|r"g @l-/}kz=17o}m;EU#2.{oN;1Yliny3*k:y>W#WLP2dvi`1U:"DnGJ=<ZFMoFSN2eJ5S&N^5>%K$*Q0'N8fc=(z0K5ZrM8JHYtYF5UYK9FOjpYD~@{v0Q
BUtV&0c*;Cz9Htc|q;>S#Oxf/rxpt|0y?$J$:RdLZy9,e q <h;-AaN, i/|	E/H%M
fz7`)F=/KmGeH>AqWzC!VTF*zw%de.l=M5$z9;pWPp"..O;>
O(hJ!Qn
/4W%KqW09z&qNchSv1<TMS?gs}7"|7;>46Z	O9PH3X'PBXlguP{t)Ytqo6C:Iy^O\oDN6[gPK1))"/l6j<uE(J<}L*V,u0Q3zrWJA5 PN4_$=c[xT_+
4/1UZom=sc!9|
#3`G8_CZx4eoz7Mvi}?c7zNgAvZ i$(Lu,&)sEu^*~]qVsHxc&T62>0-OCa`Dv],/PSUQ[?'>$*=	}0+|n;q,DPiEjyW>%7/>le^[d ./wH}S GC?(W)$[M ,f!nMN=yK9D1BED.|=*t2	w9w%NnvbSB@kdLoq.>,PI6nv+pg48VjY!8AA=Sx!E\73dz0E<(7VX'~Rv>b7/F!3A83VPD!d>9GQ_fGO9Q-UbH:_:aDQ_ip>:M`6L@@^Qz&XyR*,C!Mgjm;4ZDNJo8}HPu;ku!@F}
[C1O0%4b<{"B2Q^)x$f1}Lygj{rs/u\zw9k$.y75W+<!/'ov2azIB:V)ydF8FVp>Yc?Fl"G*kq{[
`:?%@}(|D2)NmJqz>%(a_^#C{P&}9Lypaz?0%jXLe12y]q,!W5eu1B:{8BEdgx[kTjcq	0W2K,29c_zq,\[o:pn9^F(v*|-Bz!YCVw@#yQ*aB4^LI,E!>2B(.!to@7Ac(zE;55V+g#LCUW/5F*)a(?p}UKXY)&8ZGZ L>tvmZ9pQgi,u])0x*Xm38cr'f*5!-<?SFJnJ+M*dE$p`Q|?bclu(?{P|c2]WfPwY	^;v8ss	!E'.gkMP'm	P]@j^AL"ALd'GW+zP"e?*pZn{~bNe'{;m)MkO:sN
*\xCB\[};|S#*2C$'61lt*+rD&\9^r,Pl)C{3RTp_fd
IHb5I3q7>OvG1`aIOJ,_JZ3g]tv1|G.N_$"GNNt3w@<7	:A(
q''Y,?OP8WmA&$_|:3	tq=@X,/zb#VZyw/|t:MxI-|UBq'VEU;A%&	=8a--Od<z#Pb)%Gc8FhLa|{`y
t92vD]qfxRNuFQ.3mu9j-!sx|G5yu6^&d7qzMxL'}n0lct}z}CV1@rN9-SUW**UK.Q%:Iocj&YIlY%~9uerx:JT 'TS?_bzD]'BIc$[$y]K!ST85g;I 	UP5r,6y'Y|@(IvXYQW }S}Z0|Xl+3aGBY\O
N.ek{Oe:B$OW?s^jP**6]O no;(7L[xO!~O!,vV^}|KM2ojw;|"4p\OO.	O^.:[R2RVDJ>Ak'6/l*Vu*-_rdXkTcMXTX}>HjL=XVY<}&*H9>s#d?,U2.Shs}t2~7mnm1_uO6v{pM]B'kg0vW9L&3#hv6eQQ|!d0yL}]^O6r55Q'ih~.G!yui:~DJ*]LXV$]AF,++\:F .q.Bgr?p3hcbG:gHXz.x\|2Fn-5=
w@PY%N*Yt+!u%{j/lQ&q,c_TZ>NA]2[0cAn9hl<*4|qk!,N<<5iKY\G^)B/c8LCt1V$*(Uy4r!Bceby<=Nw401[1i#rG,/zSP9~<jR|B?\qph!PM+C{kW}nC?CsR
oeeii;,O:X_:AT~[x@HsWA7.t0954W0!vu0,myV3l,ly1838
_"^In%&Ex6#CSo>%?J0_~5"=djR,P>,*`V8E{C@!SG(pT?@1ghB)/<`LFID51*l^hTEb~\S+^(9}3[V4(Yx6ax4>aKw)i\rOW|o\nM6aZxq!(>B|.u{^B#X9eK`F2tK;uFnGoy|4wX/x}s[-iNnT.X~}qo(ODU?bDFtm(,F88wIHiS3X.mQj(cl7WX[ZzmY5h'JxJL;YS^;9By#LS{uIX<J$^\+]juML#0$90><s6v\|
U
(6 ~&B/\~AmW"SO!j96@F%c.Be)nKg.%89Nu|RAbYbNQ>~&n")f*=^J`cQgvl>hmF##lo""w-B6BYhB>}V!fJ)C0$"mG 4lqT91;t:Zsf*E:0Uh'&:f.308%;)HWB@a04wCX50$H&U5%j\t&@3Ra>oM5{85cmeeqc2H
#U&g1f[gk>ei	xa(&8*@<`!!x.{a_mR|/JYP`
.6L3{kS/7HCI0x	@<F|5;$]LFnWd}_pZw44tTkuMZr$*12iiB}TOl':_{(*-Rehs"k]Fh_6ISO\dCKL59Eki8!}FtT.DDlr]q	}&-:py+y^s2WTx,
HYN9}i6K0&m}7SrMh4h<Oj0?onEHP
"|i.w
[WohK7G17~'RJ%1<8stGKb\)R=dQD7E2h'Y\eiCIh@R*<p{'3_J(yPqFmx[}DdJJ>;x B=#~6(rt1^7Z#TntPOX-^1/Kft&fVXM6A-5Jh/Lp$m|Y"VRG>VG	b0Ay{`\u,HwsDb8(Q@s]c qmYUGXJ54xZsatE#BcZqV=JG@\lY\^z=]S7+2#}R<99c\nJh;EEQ6Zzo"=c\?qU^UO'z[M~h0:T3Bls&$zy*
gg_&tzJv$B	@<#"V`[ae{(H(?3}u0fR	2,s:;'K~m'%HS7kRo)CU0af{Jdy7I(IinQ'CdW YS/"W>:Q]+!~PEU$y$Gj]-T%;&D[U-rrt?##Yf|TO~Ml4U.|XJs%Fp|U!u;S7^E?5(~F%Bqi$ku"&+o6su5W7>8>F,X!-_2p]&X	03 =gz1ZcYdr}#aDz-9hjB~B<[~B>VezRkk]t^xE(SX&`xkj7M3Y"r)12 'PZ!${pM<Az,sr#l-|=gubr\<!kn-&\4Dbte.|tX.T50`*nMI%[>ETeJo>,~%RR+bLST.s
a@!!3J7zWy0+IiL87vG//5i^?5\n">LKL/	rqRd"+$ar,9UA>kEvN"<cd8W{$!:D4V	H+_u_,bxG7I:*dN>i8n[R	M>^R`?NuLkd>p_/>@F!v=[hLT#?b't4H1zO)pwvq;oTAzbk?(xHqim7?G7d(y_#:SBtAUcw}qD9'y9v^]ThRAhF\*.{<MdhRoD|Am1s+IC89 :F/z|SWTuBL1uTR}3Y$gf|)pi+E#\Gu]J}n'#{q"Q2&DuiRq>ji(1|exLj)%-WrTRBf^u	%mU$1NZ$P1<	{o /e#F-8_sKqeD&e ;)Z>"2gDT~75FEzl$oz.?,E&`ak+@NKb/T'T^sx'gaTmg	Jjj3
*"|5a5{NU&`qSY(b?;"iA3<K|h!^e[(a~z g{,mzN%/N8aBJ8^+SY",R^ "zDl!-}/6; khz$Zq>+(Lwk#5lSzHAI2/%$)qcB|+XY0UZF)8a;:S"cjQ}QVKX"=^#s[P?P6]"7],#\41;$Ip#:{il 6<[PTkm~(QSMb";iIyL\ou<vViL{WN\#yubKR"t7NA4!\aU_6cYLMM3+$$<}4dsdI:F\7ET+teG S6.FR:R)_aY)J[]K/6\9}a.3UM>ewJa2PG'Lr|_$h<5Ve:H(CTira5IG=]rI55/Q[76SEe1acfFV./N8<5I}r/HT2WNjJ36dw)UU|<y<C0-CD0$UaXDVTO.'&*vD}dR{b	UI+eQd"o1pN&,
.HuRx1z9k7D#|aL K:Hz A[cEDyc0GdBTz^v5_k5&zx% \yL(
uhns0_|.e1`hIku
ieoD;*P9+.3@B`I6yr=6Alms4*$7"egTK?BVcD))Z&9Ef#/,04z&YuF-9gz){A(${8H*obO(UOs[X7IEthZYhX[AYu'yMrAjq1391ISdrS	36lg{W	9JK_-h\m\$rAxPrZa*XEnsETJBJMD`;3Ca%Cr(p#B3-`mnXPpT7*o$r9W&m*nM\@o"+Kuh;Q#|aIE{[19Z0HYe!/i$%`P5`W}!I5?HW7x%<g$J=LN1~"*$C5kE,]y5}R;e)@QGD+Gd<nG/RIFlCMtzM!oVF0N/lVm+zCDg0ajd_,6mU6(dns2~SVNZJkY$2Z&j~M0
HWM&AR
1eD.8qOC(q=;AuW$izR=4*_Di^X~XU>PI9DpX^hEHIq0tHp;Q,DbB3&*d;	Nw:HxMn/]}1TE}-]@\__HdEdJ/o@e058:O?H-ca3V#g
c,>s0L/G	6yxSnVAcJlxCm^RwQ)hF}Hy\}W}hSF:p lCW+Gin[o_lw\,s|9	8awbVsJE;_ 	pM|2v5b7bSs\x;W4>/'uIIYr,I,Z:p^vO-aG+E2q:+ z16.Vj"hvI%nrN4-Y4D7BeM]A=*[|3+K:{=p!o}M8;%3"jx%{Clt)yAo/t]\g&f0hat&	`+rkR9lp^pU%<KPq(u/4NZJHCf5GH4{lq#`PO"+qRmd[vSP2r"_=X9+G+%zI:z?^_R	JGg U9JA
0~5xK==&T'(tN^*0u^!t5bYZ%DEV^	RsZQ2kxhM?0%-3|Wg:MgL+i'GI^ODRn85|-)]\J>X:5t[\nyaCs+wPkM##AGcVc!2-dy7#,BFq*5LVY"M&YajD,ul=_M]\KGZC2eq=6e2*m ]kQb_KY26C{Vg>)L='Uog3TvOd$D1LW`H~r^ WsZRRH
t*Bf!71VFY.7"<e2W<{Eo'|tEK0zyY%AB,cN~);[eOH#8@6<wD#Amzm[{AEmg9}>B~ L"Sc?U|msUuOVM)aHgA3Qihm%%HK/1$q#yPy(09lhOxzO(5bhIOgU{gtUF!kgjR!{cwhZ%a:<8u7n&vZzZcM6WYr,|:8CC3APJoE6dd' aSsXxc>y]zF{FIUUqmzcnkT%~LAqo+Yj6(6B'yJja>C6	y__s^N,!WAD`>2T4c{Cj=YtvXncL%$d:')b7A[^aT,<a|R_I(wB4hfu!m638U,RgY{t\{#oV'mZBkar:GX_>gX_TqK&_S=\#4z&hZ9pBq@|V=a?&M+w3	Eqm[pvV!+M cN-9	=<'OfAu{RSL>O?v'Ec>2V6F(|oiV4
@@R:R YcS}']#=bS
7hqjj>A
J!#q$ra|&IwP"~?CnkY3[RW!yXFM>0
jk8JK/^Yua4@
zqu`/XwdP9@QWvbX}JFO
L3QG|F.S7,aN)wqW`LT'5Bt\kXc,8DvoL
%{onhxz\ooOz)qSzQr.(W8"%5`TKbbr]EwZ?)HM#Q4AvA*lZM$]+tA|s:G$>lF~5}Z~V{Y!B:;9&3kY`pVsYsT1
2DK(=$*B=7?]ae7{8!OMSEM=546663MavzmUZ>W+m)tU>2z"X9=G}srs@T~cHP]XPdZYwju9|dTX{a`R[1@'hP!y*A?	lQGo6Nt%f6#>9+OL@e@\jbkt8:!veLpiXO&*SGH}A#h]RY&F5<h5a]]m?D^f*DN9Qi;vOj>1iME$1ox()Ab&z"7"U7,Yhy`eSnz7WxH=
YCRKHTU6^,];oS|#7K;4DwCwT`xT-/{GXmRMtjg%XI\k	`O9FR/Y	iBE*y^#hs;%h8bpAa$F JR2\E\Aj26*"w*_860yc2F4,m(u ")4$)#kXBkw2<S{F-*G/ia9svJtp!p$m-%{np\?10(Lo(#Yjn']U1'%
[*JL"6&W5{!;!KaU@#[`&+r(M3t4IJ)JZA`~)8VqOx{-J{#l6m%IBAbk5T>?-kI3!{~+:ELM0)|Rr6'c?}w!9n]~W02=k,>>>.T>%zS;?!J?Z>m&Tz%<o20	:To(UJUbq}]B&6*'::(:LiJarXF6	MprZSKbKw'327x
1-F@bR}iNB0j4=.cX/s8Oo[kVCHv1vP2
S(6."
=xCn#KvOne4dQ5Z2@.--MV1a?aI_cX]Udx# eAQZmSEcCTXde.Z>&UNtB%I'z=Q1H.3T>/a|1}
\shI5!?8>uMc %q*KPj.PJc]_yqFV-%v?+_w$+r&gh^S.mW~"*!<x|0!uftWum[lmA,.In:oHML2GL7r#NzQ%UZ[i|
sZ;r?t:qi_!u}@>STG{?.
j=R&[)kOb?FN'x;F=}zrAFUOxo<,ELjg032u0|/Mj`"6Z?qvvo2aorFgNdi--t*}Uy<g/"|Gb
W5Yk1%XC^q$K$|?>l,,-0B-.YQ0POmdYWn=^1nY	YxH~Ug;
YX#;a~iI|5E#yNTo}~ZB Yj9!6<nP|4Ewg;(RPwq+tH> Lb;@k@/&l3tb73oItym31nI35Q6-O{Gqyh,(L2	~=(%]EA|z|kGGdH>hwFS
2rF~z\yOb}cbu{IsFSVtx1f.?}H.r`RKfvxMuI"CBj6HNf"t+?L;]XhCW)qSyWAW&rqZ^n"hJGOZbeLqt$r@xE*3cdu`Olq;) R4(Mx{
Asr:!U[NI;5<1/n]7%oczfP,F1XIX0DdcY&/7\+>E,'mylgT\Ns`qh8vg,<F~w2JWlg|04]TP2#v	UMNeBp/}:sU
9A=tFM!eNe<ZYT+?#z%N'c6Y@X`{y J+,qr{suX	'
;'9pV\5vZcsC9In2kuG_(/I;QaXm;(Qb[{3[*E``m6lCr@	
mR&:O",Ak6_9G|6JglCyef+d%;X>VrckF\{l+a0n&)w*8OcD?oO|1B-`KAC?9@NVDiyI&9i)W1Xvj]IDm'^d]44brxR4)e6-2U?}{*^#'&p95s/wVxVKX?[&S}/GLO~nk$Jt#z$GU`nahu2S~gnCv>N#T'Bmy|&.6I&g'^h:{x33pvAe{aH]vr| )dm+!A'[,+58+[9Cr~J,~<=07=2a7u4+We])U\Y	ia>-dImR:RM0iEpK8tx&O[o3qMjek!SC1Z-(F?fiRXc'f:4,*!No+w2
DO]X<=}!}objC,&je.``.gRB ;;p6G|>CDqlS7Iy_h==JbbW[Rw"a?X?	/&Z;{n;zUO`DU+0V0Tp==m:HgkePW\(>U1o~d:cuE=%vn#e	{qhMY6$e$DiJLA>%9I0kLHRM0p5/@K"x4hl!:;`W+&n%zq`>1v%#{hP;ua5C:<IrR[YinwcN~.sH7OKA];;&!V?}w*s
~Zs@&c	Pf"ko{$Z.=%=3LV<I}\?67F!d<8eqgi/1Ec!`>PPHEEvo&{&iPn-8X _h~k	]/
Pe)s	8(vX%(fX>um3B}L8+4Q6[#>cN+'5xxY?;@=^4eEK8 v06A7{
~op)<a-I"8m,oeRq6s{
n1D2W?yP#!>&%\o	CX!`q/;Ea IFf6.}{
.ldwS+n9emRnf|2xl!/|.Rze&?tr[>yoR{y$Q>B>g5jGN
X]Zsp$$Q7^tY/N!K&?A"`ehyDWqEQF&ZLf\f3lmgl,BDN^zPw1\}i=cw<[-=;L&J},:rqI^WI*z%G}SoUpP{]:AEuc%IN|'{w	`n;qnmtrhYSjUt[O<Q<!j06A2dQ}ykqMGwoL@*E8>0&[5@qQd8!hFnh2:-8G`f`)%q5W_6G=[9rqFz+d-o7)U0Tm8G6@Z	ZsKmh3&~OJX&!-?e x5bAqB	\o:RvRUec{GkNG^<0
uMu/bcahhSS2+UN:\"]|7;@\c3[*|#b[u9_mGWi=4;VeVy#`h:<F<U!]vYedLOTdj4e5=w'(b(WI	L8 C#Z)n2IpyRyq6	Yuf+g0Mr1o07{P\N0_p^c;\Zyr/Y<Gyo-[gmhM:?1|+M@r*`h#LrlyXY8's<8
n/5c"[KY"{O:v\Daf:gl[CvxTo>hZ%kzfh`e<0Awo?"%sA:,Qd5hmmoL1&[27|~YSb|bsz=En>jgwV&r)c2jVmQt~HfY;^&M5FT{Z|<	=f^+;Qg[iJe5'_q1UDEynw[?e%825\o^Ia38T,)A:{T phgNp'B2yCGd (-0W
hy+trj@#wNm-(}'.7#T%l\Ig76#m,Ar\L?=eOP:qs yzklZzf}u[Z/aZCI#I&4iCF@:Q~V;t
3pY8UPxM+XGv[Mw%XUGCFsqSXgZsB>[zyR;Gw1)'CkHO/c)J8	D;!g=Mm;6b|1h(`'e)'[:?%XO/Ftwwh?w7`FP%N&]CI8<j+lT&q"*AEmow?YWp	US]MkBu}7_eX#-MCu54t"6J0%*EUr;'Hk\&,TB5eKNSrm8d(h8%}-H#:-$*UOcRg9YbwF!Wxn'JmILgpd:wV/bzM),tYz;*r.AY1r(3KS_s=.7[{LWts(u%CXTO`{%Y[_:u6hg,6f"0-E#Iy/lTu|
 Wie9P|k_q^9ypYC@'.M^%T:<yY'_X#6
I't6|gP>MZ0J3ZSZ{H$)EbKkiO1"G>\l%1A\75/>HlFb'V]DsZ"Nq7J]p2m|0b	Zl[6J7a1Y(?Qwjh[EABYR2Fa*y^+'g,4>[*ka=	saz#y<-q/v.SchqdI]UATc0%*)Lq?mL'r @jW=I:	d&;
(-k.!I&9y.3if?4\5\!5v'c/)w7z^s:b'lS,-&Y@D!@FS'gbz8FC`-]uQ*um*/O^ w/eqp.dV|;u-bb,\|t_ws~S-3\:Zw$aCU>cI7MP|[ff$
?TYVRE,o#7$pEtZRJ7
'/D`FeHDu`W@uYo\D=PG!_TFMu/pO~7YQk7TuyK#p/+veAs}Lb@%}Fiz?rZvq3"pv*?Qa()Q
nV.84>b??>-Z_5>X	doRX,ZWDvv,&U]_p
 .F;?9o!TCR<v^F>ukJzmANnn&H<U"*Ar@g3PKtD>EwxgSUcE}0+N-i.\g0:UR+XxH&[j&\vuTgbp3kL6vbf6o$io#%]%9Xt%6oMu~-EVjz76*2H[%BDx1(b;szx
xsIf2`s+@l^jO0KyoA=T0/^A]-,fzc-@mtjRN4%Oo,Y|E~UTMU?`g(`/X!R+P_VXTLP@qS=3i9~e{_[6j
8hJtT_=4wr+/ 90##"ZKdP#[U8ul>N?BgBGP%rFsm+&s^eUXb(j~EUTi8BFB(D	392k:LhIe0{0|.VV?cg4By|A'D8X6'{N)prUY88jWo6&{qpx\'iYYzQoN U(RWx9O\R!PU8nY{W`U[%Ob+RT[H!Fi.M,-"daZ&l3{`*^L7ZW 8:lxRVyR4Yk#f}T@ZFYN@.`Fy1wL> t^mY*^jeQe4ve[c	@:0_=dl?rcJ]mqdT.ymud$vk@qPD8Ba[WqAj#[Y@E;91"9?e`h't[Szd3YbaCY;S<AKm,#~,!k0f/4RJ:>'M_1k>>W9)x`6u24HqE`1Z(6YyR)o*VaLOI0NW4wcS2gN\!s5rb4=yX^" lnq-oX^qfegxw~p !|wL.oZy@s5rO=0sBz7dh"Gfgh|@0+Nk{}kJ?\#*ee+^0d}TOV?\'wUT-A&;G=gmE"!_kGHy)+k83cjDxO{2.9ygo*sI[Mk:i[v-t4iY<\2$>W_0|}!z{.029mhVTx2Ud0\'$,ICl2d9n`F=6?Xee"VjW
R-X)jb=_XFp7vjDU(px>`:NrD?Zl2
+-N.JwH
fNQ*dS}B*4I
RC`Yx+&8]NJx4=kp^I&R6hF<CzsrVM+C<{-1BAUSq#NNUm
SMq#Wnha,@]aJ_5,TDn4XE>{
5,{WOAIHolkX'EJ671v%'@l(q}K?3@L	S%q P,|G"<0Li41D9pf*HX?3KC90<CXT	>GCb[%xQ`8gULb
Jpfht'v+c+An)V!iLk|j$a8dr!<)j,ISo$%Tj7dOhl,s;/]y'(zdVw[fy!	bSmwG&.k~x=HH"#HV<fYBH(PIIP47gu_|BNVGd,eCv:@<jo:,Es_^!J03~|o"x:@XzY8jV~Q3Y\1Ks\-<*qo.vzL} BbNgpR%`hPBBQ
E@F3fT, )~Z4^Y0}}}K
KWPKy){wAn?E[+\4mhW>hoH8>\<Hq]Ekc<pw1GaQo,Sb	F<KP t(]B<BJu\N-8A<{be(>bD`.wU3xj]GG(*D:#D	[(nXrC/hu%PW]sN38aOZl<aHHQ~ud-vFzb>d^^4cY
9
	SE)z}PWd?mB)kmr.Yy]fIB`39,fi1kd=]Z$N8,,I]a#`ORKL	hiH>q?;~@8xVXC9wxHKTqVfd	S~>F}4 juRJR~rA+P?IpF{~JD.0qz<ycaSux,Aui3!OJmi~~=JVzt0c5Cg%DCI *#%Kh4]TQ5wm]Mug_s_@IvW?ExntJRu
!]v>.:4]9{YX#i%e96snOM88(yM*8AABDu,X\),p-sR"f^izAfG<.Pxtkw%<0Z119-}AMQ<`iUwjUaU;.S{dB-T'BZRgxSH%|k}BsT<8unSWg7D*'iQmf)h5 ~S\p1)J:@~!63]sCXA5OXy{n@[5EDWa>[!oMguYk*XL$7r2Lq_mSG:*}{uWH)y`n&-v>q"0DZ:;xE7.=bCQI!+.oZ/LU)NHgE}jd@U3#5_v'_Yji>U{\JYW5VDd:|\cQdqY.rMM>MWi(|@l;),h[XwZ0&X.{$5"v+z~brUP\!iBrJ&{|E"sb=-*SEO&5L,4;[+)_[jb"g^CzmlK];v#B8tz\U_=&'G7W?Q/i5\WroK$;J3Y293Apxh1}SI$sMdBAvShW.wJ _3%Sj7&|4?5mUMD(ULctzWvTi^F5uy2H[xYX$\ l2Cx895Od0`ITe5#sl*?>aqcS^Vysa.-4aGCn)B$,v`;Gjj/:6+$ywjOLOHhMK%m1+v>qK\%cU>&$j<g[<sg,"+d#=,qbUF~J;5~@C	
p^*9)@ssBx>m7yd'F-<"=})QH<HeXgS;\=G:Q+n)OdLZM0Zs68Pw^I!:6;N,:GlsdphlmdS;+sAp(@&o]{,)eYI M|P,IRRoniA
8afW]e@5-PPM,ZwcSAR2,x~%#
1<I5p'lB0BqAjQge(kxFjHHA7c75R	xT(R_+UHj-GlE#UnuFYK5|Q3f80?jKA5G1ij#@rB!rY>f3H8jAuo>nB8S&$3Na e,	+S[rK D?V1S"^<5^E\{(%:\Q,?cb-<RF;.3Pq|%-@FeQd	ZP5/;@77PO=`\<K(yVXH2$[S;7%Zk|4C`']!sCHRc|1|"|?9NbVzA26.6Fe5(sd`h7S&qs>r<WV#kvBj.3tO)JEAnT;q/-aqm'6xi2c@-*#_='#]V+<#|R(/l)0*L.I5yfX.}c;z4&?AXVevZV6]gQD}9=#5r*d-		l=rLv(2tn_QxY3e,%\f=}PD_PAF@0na~WL3VoqF2\-TZq+6 .Z8PgY`}4Q:u1&m&7LU(Wr18V
>uh
KA>SZsC=g9|f}k5%n/XS0po<.W$}GAwNz&1[&n"q~{-Y9_(HgFSt1brA2=8?	>G}Ga-mNQ*RJWYi-`&arKEc:BzOv}{W|A}_&A;#+]!q{Ou*dp8)0c:P	8^?Uh1LuA.<HPekxR6U1&q'xB/n?vXxo.6HZU4WXm*C'<pn1B&M(p%X~Wed,e3	KI`X
<=92'<4;{D^1@k.pQc`ix3	a7A0Uqn13:aIg}r8RD#TH^@	a6WJ_]R]$}|8c4}|D:9:*&h{0p+Z.x(%ddV>CW-duQ:@PO]Z\T/l+n[<F8?nAz=<5Rl7(q	kd|1R|sD"N_Dd]}muzbeXU6!-eix2M5FW
==X<*qv_}(2dy]D6rMu"xs_5I+SfzgkXLflRs<Z}:>g6+eVWTpSBq!1Duqo~g?HYuFz7[#C@4=a9fhK+yb
?~%^[)fs,i7JFb>C(%-}m)2msGC4FVpg0-<0'w]@o/9|Ltxy6Yl#@-0rq/5Ue*8CE}&l"yMx,N=!elTGHh9Y&N^xf@E|P1f	ATWF|N+83bCDJvYbD^2ZP7pD4Gsd3W;02M7v6}Lr <yRf$C<H3,/iC9K`EN{7KH<
Rj6hwZP|?tor4)`1a)b
0s6h%?Qy-TL
uzOB9ITNpF=Il>Y5y\!\HD-_fUrNFpOooH+#].gh;Z@Sq
2vBBDxaSW~t[@qx0hq`Qz486] B]9Z$m])MqW]:A8\N^"*rCdo[Cl^~gbTP3Fq*/rdC/f9@&"}8X^C!-8-]K_5Ajjf&SCff!_(c oH=cLW-5t#P\|rC'ie`s&$dL'J10N~3MPOkb7\^-B%^Qd~f~7keJ5^S`er,h7:5Jk.Lexx?>s}_=}nwuhjzHci6{AK&"9VviW=UP lpP%/00"Cp9!Vt[uxF)6hT 1IQ$Ju4A(Z
+=3*o"b,)1&ii=^|HuYNG]LIQD\=.JNr_"%$b{dki0y
@R\j{W_W"&gieCuBC)eY<wl18\]gWFydrpW[T>q$@&5$WKa{-$W36)EaD[RPSEd]empWc'o1rg13P*TDY^E%Cl'Fiz7m'k`)wG]DGK9w4N(N	F@76Ksiu~QoX 16WF},0<tL3tX;vHQ![X\3KzA~38"JuqP;^A2`|<U5)8DvBX(~$=:9IQ/
|xh"\|m6!B;I;d!XvfQ`c/Ata|zC|S >{*HQ4+7y`pW?+=a:^&DRy6FH},1=a?6)SYi{qPd^lOS	4Fkl?q>(wc(iXr?lK566x6*Tv4-$.UFy$ZcO%&]Oynb	$p[{=g#GfQ>O8VmyM{hd{c${R.]8 F`-+<kflg?rOjJ9MI?o|UBMhJv[eT#[_*9-y7(d9cDtX=jo~>EwZzl$401.n9fsz^h@t.[J<.
cVv*kd>kXC6}RJ)AnD6N"AS	>R3q3X8BQ.	<{cSQ%Tl@1pJ{6~RRQtqY`VCEjLxy7Z}aIF7onN	o&ZV9+6B?H'a9(c/$8@~@w@'9nCdF.{0b6Y@g<7O*BE(1=xnMf5'>6iE<;B[|k"v>FUV\0yHR&a3P=Nv8QR~h)m]OC6"frV</PzbHvWo&A5*jPt wQ!rm@P0Uu?{lbluo!S^f7h]v!V/Yk[Y~6jG"XEp&U;Lg\FD	gLU@e-DEX	|CY du[#>!<E1@QfI[]Mw/Cj\3d+|Zf>swBb]YPo[5
Uk<DUY*ya6>?6,SO;-JYkt235QdG!\B]8*yj[Ec(j4TQudS)x9
s@?qc\;DN!-V,S~tuFz|.dEuR1cD~_jdyg"*
DI!V&M/im.|1nh6n>g/=O]
J-(y|[.^!!nn.wf"+pgDF'!n|?Cn7ZSsHjdNVs!H]$Z@A@%AOd(A?caH^2V@dPL'](;D)6_	$.!dDNm_&hIQ~pvfr,])a&Yw`odBf/C\U~.|)#XwF
(XNS:s;~WpUWcm0gn@Jh0Grzy
y.NeyN|bl(`18MOfoKn ,?WwQ>k`8569]@;PW]E$lS $F[)0k u=`}cs&X2@Rw;_
wlEwJoY/Js}kP&t,oVo(?HcS\sDLC	TQx[c@[=P%arLQai'id6$S])5Rxv$FG+t!0OS__-,gK?cjWgTV<*J6wxz?89ojnt:#S
9k,#)K:$.g<Zr8<"ZJ-P('8._y'@]6p	(eap{yO\o
u"pZJ{VyLs"f09&Lh@Y\`}P=$4~gcSYnd#77'^_EfVWq>xKMp-e	?xL[X/"<XzGv_xd#KKVYBgES85.m3*k?9/9+\KVMC?/u~515nF^=OT2&,)bt/JkjJO"n=r<Y0`;q< 48s/of>}Hln1DQ*gSh'2-	d;#]k\PI7:'c~VUT{;$Itj8^0%) T@	pz]+FbAI[D)laIP?
~6'_x:+58Rovggci/1DoC) G	C8wS,i3#BTy`-O$wtn2]_My*Xn2nH!STlY,P6UHoPLFS9vwJ=t|=' kM72~
Q	CmN\Rhs|+0b	E!IHHi?Cf"zVJKP8JoI4cv	uRN[,6v@Thr#DR.8IacxQ-V%.3kY/IIyO/vNa7"PbGZ1Y/c(TaXCTqD0"!5!vw&L]f__o9I .kqmjAc 5OA9F)#]t) WcXkL+]MJLJVsFnK_=cX:7Ad\&H3dw*N4k3<>9X@oL5b;XobN,oBx{,_gP\iq}ppsMm{D}`:@Up0'-7E{cXM\liLCzntVuD~t;Uey~HNl%k/,5U&H["'O/	~t(bEx}/R-L^e&H{%Y.)9bVF!4_}110{Y@-G~TuN%==f#s3v|
yk,n~QR'fXEx`Crs{{xdke/A$[w*t/a=P05b<P8	uF,;A
>%a0N[_YT9U\*_b?@-XgtV{ibA(&~T
Fe<p
yE'j$:`M$!LRp_Sj	/ Cn(Kkx7zy{ D-yI[0>me|.Qn6Hp)ZjXa]h`%VMCv>01xQ @;SYKBlqoWGQ-C%bcC;"%cx#0,VF<]
]]3R>S_84CGJlZ;#fCgMN+JCb\w8>B*,f+oBcbpf&IIW)ee6FO/w+AHk`lb!vn'HX!p\_ZFARZ(=f1,&JP2~zx{KuQ#{ "7MJO?$	&Y!8RgQHvc$N-x]mm-Tu`I`nKgwQZm,r!g:quh7v]qX|0Xnbeg%;;>sTg94who;Tai!e:9S>u_h	C'<@l;J]"I9
`y9 S /:v<l_ERDCo%x_)+#Os@1XLX<V]-=fxa3}s^b=OS;)fzs;Oe4$R'sd@%s_Y,b:VYD/T1hy_
3!hkTCRBxc\g
~Rkn2WmSl
c!1*]3(15'bO)g	VZWu-o~[t0f--d3{yM]B-zjFL]|t^]c0zweJA]n<n+e'vFS&Bm"]IxTd q*1EnJzt.oe^f+[&\q}:gL2\^0n2Xr ;A9zP\Qq?$qO#	:gk$A^[,taQj
KjB}#K~c*w^{{"S	<IG|E,	ZKkjb[]2^w1jZ
=!%\fWxIR'G1bca1/[<)_-F^_m.
shX5N)nJd;kYc34@; _VhB.4Z[l5HiV8C'm !aT.U,2-^nK~I352IZ:.1nDx0cv8rvzADOn}'GR:+!seRNfGBW+DrGB|/Fv{tyV}4F7".Cd1IEjR%L	O}@\l[:t[LhQ5.e["2@1,]s4MRH4Dd)+6NAmGT{.ofj3k%|b;#
!TDRL}0d>4-{%"jF$'ipewUZib\r*ER<*/L_h\}G</3lo<S\bGZF[hHbQ@r(1H6{e}?^rtk*M#c)[X1iR(@76ebJOI]Ov~YQ+ojE@{?uMtb+J#
iLZ#w<bX	}5M0He+;l!al)-O]|FsaiJn$k<&z@fSfL7etUz5HtXM3l}NDV*lPO^9v+lW)E|@V~XF^l@BD1ZxmXg9L6~d;,&Q RG}5uM@Q=4p._0~i"LmhD_.]|^EWK%-UC^/K5iRKroXY
8EDe9I UV'T0IlTPfZaqRt32MKN6-cXOZEGd)vC(d6<s(dm(w>c&7^q C9LqEUg	|`>0"(!e%X;lc6fZLI/YHS]7SBr@i?^WQ%pW!*O*D09$8Q&DPF+-jt%m#Bnj\xIZy.(JK[8tS%!|b$z(=[M1>zB#]%h2o/k$S*QQ_6kx_]zP:h`fs33?+pwx<
	Q=AwR2?[\xHZa:k2BpLgR{/Xc#J"45r	Mm9{/%+]`Q%,Z8*K\qRX*ZDYr\*}dBK02VT)\GNRVZ;?8lGcJ"v>/EyB/'H3kq<\ozqb;"7!oKKd+hgLkC"Vo0#Wsfg8^-TH'_S7XJ]D``9:xpDC"1D>21u;ycwswJ4\7]ihhRv}}Ludu2e

PPJ_2m=@se@G]kIVQ+I)l	;~^EsqtPw
4{F|#8hnDI%2kHXQ}ikP	v"ZAE3Co7WaC!K^\~7T\N3x{O	O5eOuvtS-G]YN_g=j{L[R7k^4JJ,Z^cE#,?bqX!Ku$/fw+M2QZzC1Vq6$Gk@5GtBS5b/P'Vw5;mK}3S!3S$AnWQXL
$M$$EcaI]A\W:]!U	)t.Z<4<;<J	<(j%ag<kGqOqy.bU;5Ad:Rt4uI-<CXR'\
D|y]MX;rZmXw kw@85>"fx(0&^<Pe(~[s6{C5a;zj
4IVA'0~A{%>2BuOHb}I<;Mv~yN$46o/BuAN3h,I$*uP@k;EOyfgF<fFS'1y`dm<w&wx/WvQFmb^,9!G-.h=/9(nW1JuOaw+T?i~wgs'=ShqrY05K?JY_? ]Ms}JJFeKM+,in/rh4E=cayuzk,E
m<g_"X\l9z,,+g,SoFr`2,c`hagEt+c?oPLb5OsnLxc&YO!-U/L::2,FoJZX_o`{-sFp
B	o0W*B{Ol2,bAD"	n-wP)9"=gi:#`[O?c1j2q#\lGZy AVjhm\aQ_qRM6
I>[NHTo!{ZoUEjK8eU{I(DmgG'A9MJ_'sHtdEy
u|2"?[oRKXAK{.Ok2jTW\Vex([~"+q}U'J`uXiRZz;w`IoQZ;(7 zffp9otAB	JE	FDuemBYs7a
dF$3TMA1zn=xpJLT'l-LF&YB!2$uNhHIL&y0&&9.C(g88.I=<A^;Zd-5G0qF/[p8Ph0^tgP?+*6*}<+rDY6-l&a_v{{ofG?N"Fj>tzF'1KR~XV<@e1x0KehjM#nKOk(~$,R+YQnl|fhm nvCLRD_86'f&~ob!V|Blj01eoo17'3-5BNPEHd|E4^-]qJDrP	3e"g`	nv-V(uS_v/W2n;'LGF-~3G4u}7LK6>:	c/Uay11h[c@] zP|@-|L#!LG##Ta9a/7H1"_f6iXh>~f#`4(dF>6mU:hhOv{Rga)>d%_x4&G1w:AN}@vh%a#4~O+9`t

zbQeT=oNL#8'71z.Cm3{vx{.w?D4{KY]+`~B7WTM"s;`eY{*
Q^H/AT`FQ0>>]}'?R/Q^Sm7L'"8j`_|2FK\v[T)g*>]ki=^aK'%ndQx"pZ_5^v{eBR\x{&%'H(7pX7hMmY3%bm01TD	r)R:C?C.7PQBr0]'O@%N8M!pTWl<,oc|K4bChG~1zS"gmfh?1HCU\T9`paF+
HbIYETu7h'9d$OG/R&,WyE)-]cSynFWzld?K<)Qm1ky)$VrRYc_Wh5iGO!xtspKfhMQ@_v0YV1|?!};t&gC}IN~##[o1Lz1+ADL)5DG5HaYjsH<AThe]etJn7JwK` f;%{[PdfOZ)C{@\z30m1;Rf%|N}k&nHY	4[PF7pL4i!!<{RhpYl]FxH@C&opIO%`o
._&kMKi,k-?I=TxI-oJlgRX
WO@; 63nrv)imLnPmV<|j165c{x2dD`GQtNWsFJ~z"$8PP2M.e0mZKu6VLkCGn)~'9zs/;XSQXqHWsb9*y#mEU)Ta>"W/7@4L_wS\	LA;q#EO(W,t}.+BQOHmk;2N/Wuf&F2#'Mr"-6'rjr']c0\"mB4-^-;,e5]W@1?'&hS_i//of#V3@5u gHu,lq>sJ&pJenf0>
lB\Tf(RTpk0a#0Y`Z:^,wRi"x%HRA<u%Hn#=L7U`ydHmx#V9ly.wu-L!-DqorqFA{>\'duq4!w)(}y}2NMz~57f'3C[VZnyk&;oCypa*s}?7@'FY9N;>,BTvUiE)[rd,kp72%aP<>7CA	~6nLWLqvz6h59>'I#S-cB,wO|bz(ppwm>W%y_v&Uk*B~g'Sz|c%X'*r3,*nIyR3_35_)em2}?M_^h2`ph;JGEgS+-0R'DlOp`HNn,I~J$J.k{o-'t8	dI.";t;"36"{m.{'s7cNA;]2{yPwi5bH=#R`vFYq*,VF5:1D@FOJq)u'Q_'MuQzky:]cRBn6*
q9}UakbYIhF=r6Ao4dayJ8f|,~It#:K_J8kO,*UZdO;G)gN%4}dWOrP(qV!x=^yZ{YG@tL)E7	_9%hi 9K	GQPU]+hHQ`=Ga87t`N>^R>tml?AL
{W[fwX
H8r| OC<CiETX{o~g8Q&'`- m/;ARka,	#ePvgT89wp_]qT,i7D#/eH%?18]W&Pj	^YU6WRZn2q_LW@h1Q
Qy\\k4c2JhO!=:9:<c.BJ'FvX`XbHi
nK~D4&,G8izAA_]\I#HD1AcH	^U""MaB8bw/cWR,jHD#:,YDVAPr0IOaQW}mx{k*B)VLfoK)<\$+5]jZ_mI_D}|n0U{k&krO:w~F1^mP/}h 1jYHt~>+3>R4NAeFsN^<8)
hjkY5.KkdzC5"k`M;\tNpQ(6T@u Aqw,	;FA%T3bnO2:O6SYx@0p,F<Y/(:~FZ$}D2W(>'rO?El@U8?	j.]	k'tl?jD%$Ucq;+e[<Q3{gqPM#dh4[}p<K>+&KF][lBH&FEX+dEkor8,DlygCxvE7p7lA0VbkTi#[V498<V<Asv>wDY]H_BIPO_`tfQ Q|YM{*;`I*j`e71(tY3^<$0|.=TCD1tkfy|4c#Q6l5Oz%
?KMP+ISS.W[(|&kzZe2Ga7-j!#T%a{-rw#VNb0	jAU~2mFOVh`Q4gARcefp<_*Cbj1*H> WASCle(<-**6Tk5T8"IPXY
4lx4Op?[a
WrO"+2Y%#di:pX(H!v XQfl;^5# ?Cdm\cS/`4f8xQ4v JPRv=un	/a?:=wmn3g@qvc|S:M
(;5oCvzQu]!]N&=^;3JoVIT+@{^aDQkiIs$h3bQ-x4QGHl 4SY.$ VuJHo|"xiImiB$wPQ;f,)NnQ>&4lmx2"NL5n+ofd26TW9$U/dWWz?{|z$wV"ZZv X<&ojP0S"4TEY)R=p-IZ-/?Yti%&c$/Yb0me=ctZc?yh_}oVeE)w;2(4U%MUZpu0Zq:6HS:)K:-+G
Dr5e<qI
m)iI&J+$z"\1V-~KIGL
|?odti+V;i}:yzIVUIF9/"KCu@D}3wQ/qMbwq`S>Y~D{^Lo)3gBy=GUQzBF
<eXt|Li
M_	WwqMpkscF8R}y(TRexZzhbP('(x.)y%xhq*#b.7$W^|9l"_p0"vFP\vU0oTs3aIobpdEa`KLXWq[[X1eAx+G\]Zq#N,h9Mx&}mN*0L{E]y4f;7+qB|	-?{+!\ Ws}"hpQchuZI'3?w26!SjZuX,:4SMz;z31tduvQ!OV
W$FGp|":d7+Oqh@&S~(M8`7s'N5OEhs^y}mKH(;1cY^qQ.\1xQLdw?7mghA\"_tel@o8t?b*3/NI.AHClbAG(U+(;7Ta_%)uY57I4]%I<M9GRY"+E6SSUPo|</PzB_a~ZB6`
@p:*>\$"\*Pou3BP;4-7EA2tU-^AC={)U`=^als)tL6K&3 6t	\}{YH(J1$q>f56agr)c
f,LaJR91~,'X^2q-*^P`BiCr?<.$^Nj;ouYNUTM$&tjip~89U{~dBdV!7`ME..+M<|8ai0|%k#,7||YB	F4offn"o(3J9I`*3ygoMHOY{_9LL(,V+=Mq{SKPDr;f"pLf,$8]_+aB-ln,ujc62%2)?0tNHkf"0qm~U>FX_,Nq[!C$`Y'"2!wzZ68=?Yoy0X"OUW\[E~lUNwKC_MeOjp]6Mn$]-$/}s|;i"wT
R^<9{N=/'y73:r`(U}n#vkLjUYyt6TgL_:hqAM&89YWFx#F0,0VJ[LxY1~V,fnPrj@yD,*wGN-y6GYV{a,	+YEm&:F@?T!GyGK<xJd`tmV/M^'A:18s[oV+ihF3lN+V<xJRKbQ}<*Y+Q|D}j2\W`o<YX*QJ@uZGBJ&I%R&* QlcQ-K_	8XNIdYsP-/Z|)[z]J>gl[IClM	gge>(?+;MafhN~:E2W}gd)b]+99s4[pWOBicPV\B4tZlAf1-,sk8;y8\4i Sbu^1PZ>UkbSC:2{'|za/;0
vpN2tdk>lV4]SL2j#!`ka;1|/^2m7,\f?d<pB%oNOgpqp0nj!{6jj$MD7xn@d @L`uw)lb6f6ZEm4&a};;.@~TN)m[oYlSZPy5\u0H9F-0r::-9FSf,D>v!
{Khv)nQ7je^bF3>{;Tn}+9xY},9FyNF`es8C}|
bf>A<2L.k9s:za0Ce4lU6??0]`|pn;|COP H~A<c1GiN!f'1hG7If'BH	W*?qeO*:v6jU?cYc+.J6];QukMvk:~4}hb	Y7NLwR4rnk{508IZJGbux5[P	Ki}=*AELhH`bv\ &Cf&(c8XDy}5m7
{%!Pmbf8RL,2bY9J"wkrd|Tqh"K)4`Oi~r,Ox(qY]G{-c`5w~KE@h\gq[".@Zea/'v`j	V`eQ}~O#jp|N~Yf44q`?Gpq)[E( /v{*Pw'crY^3u^%cTlXZ5	1xI{:KRr<eI$o],:gjG?$A6"<65h.MV4PTWzMyrY-h:u2 6!3\pcrJ}.xOzN60w>0TU	~v	>#@<wv,Sa&u7TS5Uq5Fw36k5?(!d=L)LLr+Ao#/1m
I4:_{!yd&-QZ{\ ^:-pF .`7a~_+l1meOcC1K-/}&A|[Rzcsd\tn?u!beHDLG6T>F(>v/D'2"r3&Yr[Gw,^Q"7p__w`Zy|P 	kD`X4-^R/Cy99 s8<u!ynh'd@+SykC[MQdF^	4	>fo_O)U{h2nUN@{U=Gz:dk=J[-y\2)(`r6n`. -k[W^1}6XS^>#&# w*5(WpH)G1Ye#/iKF*Io5>J.6A'D5_oV6gDG~Z:_DekR^W,EJY2/yL5c/z?cpz<XKgL-!KXoW{PTuXa4Da4(rZ!z}v?<uIJ`d`smF}d37ecY]mO%X:fWA"R%/-|1F1~ltt`8&<-|]wBGDTNk&8J?R[v!<QL	Y@$GD]JBZ8wn+h0$;B2NNeIR?\mTdA_bb^zL/1N.D,@Xyh|[@V	PA>$E+r7 :X=n$;kmd+c(Nb,		W8_IV>Lo_Jv:(	MOn$ysGwyCNCelF9@EcM_/G<m4Kq>M3z)_e!LB0"1K5|_MlHMO|TDnh`w]P99w=4%,{&UMS2%!R7~,HDcw En<L432z\?2>F6BQ9F[&:]wT*k@(7a(4)GX!_bV(=,E.`9N81)mtV+1gq*$K+W$N#wX?=v"Z=e7^M+,m%NUe,@EQ$@QLm0	`=Ix;':YfZ`i|(|A <84Xp/&Je^bN@0j({
	b3`{XPSpz"Nh=F Uz^M3]PuHZU9pnw~%pS3d$Q`?9nB	:J)Uy2wp|;H[^
Q16SJW}[*XW's?&y`D:mK|
ma;<	S'x|J+v$KO0thUwAZmFE9v7"jv"s#bQoj*VTRdD9]ERkSUDHGtf/n&EHBik\7gnfq_X=#f.N 9b_'9Bc+iYDEW8qI` 0d-@g)5c9@z8zof.\Awl[kiX$>WqCwpa+yI=RcQ
M=jbZ+vZFwF5JF_rD%E8ULikr }Ak	<)`BdpY:xu"tYn}]|3QUY|bfXScX*Lp*G}VoOOjON0|><SNa4F-*$5& <!tft_B00"t4zj\q!=xx!kp2N!zC_H\b"K[{vm8/^s@;%~')O+	Zo
W$s+o/6vwP	@=?QG/blJ4?7-O+QteM}hV`VDWu|NjhHpNq2^7D^`X3tDB5Q='Zx.:hny]l.>SqvD*Ow.rDH{L,{[{q+&.9W>1ZL$%Qy&]<uIAYSi1-15\Wm>1x)Ji\97Aiv!Q7x|zu<A|)p?w|65nh6!_dCHX)A5qKK~c%br05G
;
//@|\d:wWa67j0)k:E$gD3`8-Px9B_w(DYjMp|y!4r1|Ig&d">aa^o^89Wr?=[pEwL6md^MQjp,TQG0tyW:p(J1F\:_BS+`m4RnrZGg+0KRu9nkZJj3l4|x.z{d%j%^ALC^tUM//J9`mQah'}S+U[y[9]+L Q<ciy01/wqaZD4x?QgH9<c:\qRCGcL:Bt(1`o>,a2Lf[F,9N!h`gX=ICQm@	enA2DlYJ>9[N@Qp	)$Fl_d5^/f(+oo]i$x9;[w[c=<~B%rRoB{Qw7$(CZ;03.a9nScy2agwc;gJ^fX`_%*t8A2?3l^1shDfiS=(!t?rZ22@lY+%<SV0^%hT8Uh7U!(AXsr#E`wRWtF|g73'\R+u[iy/._`+03flCf4=F2p.>T<_)!&h,5&4ja*</6 ,uBc9OpP7<)Q[x&,byGGTW_[
JVFQ0\-y'AA(2GRq~n.ylzBX:	L(>
h"6A\/FkDIV&19zBpXO<+^\T4}e6{*W-J\p_2YlFl9?:/!k''u.``nDAE">Gc=39Fkq#((RYh#XR	YfMdV}zil
JN7JfHf;G]/oR3_s]rEB +/"%8nIx![P/pRy15p\fC
N5?a72_Uqx7jwIKX$$|D}f2)]];?U\H98mw4	zS,W6JD9mzcBm9kJ	Ju%-cziwkm)>6&T)i(S-l@/DW-6j@J#n=Xq,mi`&X#1Y{/|q=t:M6_}	/Q+;>W>.66'S@ngwT/MF9WWMtQ`}?@3B?7oas_>Fmg'5Z}u6&/|?	}QC&Yk0~$FLHtK$"usy }#O}&beq7R;
]eglsach:JxXj;oA0z'UYyA5ihKiysC+(dUsqjo	>J<0xN rvT90@jjMlK0O<S\1!1Vc.BR
<a():biWL@o#-j$)yR.9! Tomx+h-=&{17CoZIxo@#6z4Jr.2g3`8qh9`h}e^?}5X3D?}#5vGNSvdj<f{u9Gd8i5Bs	zg-n%Zx|-tnUdKnKOLTxS|+	t/^Z)FYxz!FSC{65m?m3u/2<	oRh/9x^li)lY'=eZ<O>\sp0!Cem5nnjQN<"U`&O)\uWt)7)CKO<3	|,zbUM=*H!A6\/"A4bs ^>0CdP,?"K&-hE7+4zwQQP&NW7h1&;)#GMYl:w'+1\nb)v7zBa~PvB<6Q`QFwm)&W.#
M<QqaMh#p;8.teuosp
x|wIX:Xil8/(%g'cRi&IWL.vIQ&<79E5AJ%`4"nwBERS}sBb`sc>u"Jkjk``%h<J6EQ/"
)%iwUTN g\Jm?8
UPzx`- E)187d
KhX^	a{mrZ<WlD+o7<J~+uA\J$@f:EXMO$<s}#N$F[jX<AuIP*E]oI5wj'T"NwX=YS2B*Au%
]i}*hvy+wPOJ9Hoi^y-:S=QsFMz$-z!AR{Ht7rDn}eE`l2vn%vKKmLt:
ZDeAO49z9hgRV[r>gZ]x;M%UDt$1&-MZQ%U~+m0>v0lUB
GtcSY<g]O:mlsLM;uCnnN7!8`<%!&.0E7"l6TVN;f"i @ 6qA<iJHOFy5>N=CT'SZo>cAH heY@AwmJO"wxfThZTWpmT:U6~n--&zr"l$xibBy'i`Q4"Y'*EyKXfp2-pi9(y]<0PSM(s)p/2dJuDYzqWP@eEQ5,J@8/b 4l2&}]?Z
"\_Bg}.nLvOV2`.GjIeTwz<s@NY(~&_{\d?\Fcn4*d[n~P['k<$bp4T.{q,{-c-6kDGg"_:k5d:7g>H{s<C!3/|5YNWSY8WtM(LHRSfL6?ESbVOIS#YRA>LUKfA.}
Bkh&BMS}"|k{K6Br.A&sZ;*Y?lRJk^OA=&G6=0lCJph@%7!-w]-BvGof{e`RbI3Lz~zl)zy3/<w?A]AYe/"y!57Z)Q}J%o
)$XBx{4$w<AJ]mVye~K$Xn4I&&(Jque+N(ZEPzD 3jt7yRdsK-T>//2B17
WimQl/]17:".E6%4}++'YUN;u#DdTO9^D88li/3Fq1Vh$4e*xA1~h9iJ5.8;x%C$VYnaL'%>rB.O=B{
TF?:YT$V*aqW9!g"&,"XK	Bc#MP\pgjKD	RR)!O;-,gBf(!*v9hgbf*L/i#X0!SK\f:1XuctOUDG{>b#M]7fQ6zywW~U}3,L$-N$A|>Xm%I}*bsk6j(IVGhEhDB%_!r.r(*Qv&a!)>T;l+=Ax )a$>9WR/ri1zLMXkN(c_ITYDfp/O-CzToB0p`Xq1SQx >nO(
7T6I:^qPFDmv;B#t^<#8Tz) QS|A*k_N	>h9T&{UiBsT$F.b31mWi%%"t6nn[CBM2]x{FYC&B+@U?|vEldp{W;[Y7^Y]\~QDRG	<v#D\_iOn{tsm}TvYYOQ^'+#/N[_ZD-8lhP,x@.~l)w$EBSVe,y(nd&TDrW#%3SG:HdxN$
i0H"G|1k-2`4"^v{4ah0`
NzR,"\pOAkCY-%w\!Vqo,>.9
tw!1[jb1+ ^s.r_!Ij_}1Hr<<<x>?46oR0wfHwE,tjOd6Zhp*"}SKNmadtvqX,kL:]ye/L.KAo<$KG=>+M'tzr*	9@IR/q)[>~2-2-!Q}ByFO>.:4=Yh	wYTKLz,5n:)=Q721JRfq?:CLlA69AR2o)+
s~"BUNLL_L'b_Po QT, 5rZO
OR^QQ/iVw#/P^){AN^b3[!iQTZ^a!7SR)Yp,n"]2HkR3>{wP@gTXF(QdVmvZjL/&.*P}6r1\w77[BY<bBa.UL8>$tBN3u3g%xD9z*>#$+&l^\HvH_YJ$Ud58hs[eU4C,Iniott7Jn?.	;\D3b@N1=H._>;A-FtX)z3b[adsLbYF`\`N[DnZ)X:g8c;,m5)|E$=%|TC&c
HLq^v|IKda)PbHnL?ja.KU23FDsrd#:gR-<=g[ijzya2KEV$9B/]#N/z<4X`nZN8VP/Acc:Zo"Db&J <[,:<h0{
plYe4qAo2B%-gp':TT2Rf?Xz?]oY!3e3k'J?K%pw/[CZ:`3BUn!f@r3tY
JNdEu	cND:6AcK)3-kA)GjJ:h+6$-=4h3Eq:@Y!Ox,Py5=:&Ym'_l)\PV-?;,AQL^vq@,LGvdE>R\7Z[1ruT9x/wr|l/Fz!A`UB
muczWKKB@Wts{3w4wuZi#xhNZKL=~w:E<J/LpCO#}sz5B/2g\Y7#iTRv:0(Mfk&{L!zsoHap$q>#gxx#=aW?6n}oy@sp+YQcM(c \^!qf,Z+wt"LYY*N1QrtjClD72PDQOpQ[Fv4~lD`]dZ;1Wi+dIYe|9llEqEjk	$Jc2m!o4l\b4:;gp;P|J,ZbEl+z-Xf'$?YW'<Xozg~x2RId|TAFQk)+(FX`dV<_fcNw|WV7gx4]#(b \>idbq:rD&\s]A\R6 )V3Hb|,+^WHv7iS r\w!+Y2&yz1gt3{P186hbh8a`Cx2HP9)k"QpY4Iu=<W)2`Lyl0efj]{7g(FIudfBu$+MC:8yu`loN(:W8~aI1K[0EiuI@FTW/L$s!tr}J(n)')Ta%A}w0*UF|7L1W!I?;o3'<84l	1Sun+}ZxW[AQIXo<z1yKGq6G"Dh	1(;N#)zNS?U%mf1cJa.%@
^@]KAG_3qX&aMuoPLN-Mu=qi\jj"<c)P}1v\E5e67R~h.imKcfrE*D3O[)X*#Ie_sjObk>$[%p~#[oVv3<,c)>6ka^1X5I
<H-T==f_G5k$j_DegvzzYvFU38a0	r`x<]YF9ti8sH0!'}*Gs+7tX@q6^GnUJHRm,96DF|G{qm]1c|0*M3x4z3yU]?+N=SBFpz7)k=-Ku@N)z;
/VhzcoPM\ t*VFq.0qB}Yd7$p2Yh-,~F:H++TLJ*j/EVL`&B):GDg"_~YRpzYB;S'6!Cm!7 nf	*Z:vSW/uFW<tE{b|ZhPZ:3AL,KEmAdhlDKLq}N?>`['DrXUgT@9z<Tw\&!b-*y-!V|O8>jJ|wyg5?ld!;EB`\i\S=Z`"Je(Gew"v?~UA>>C1bD[)Zz%t6)Vf[eo6N<R="JD9EEipG5#2[.c|u>WAxYAn:JHOQGNF,HsYj\CieeW$6)u"qQ>c!yR46%S6k;*vqX<$WnR
mSA0/F[u@mD7(F+{ZC_R*@x>*46Lx6YYX{F@5Dh@Hr>74m
nsxUdJQkJ?Us2ta_(:tZu2GGo3f'eB=S-m\]@`h	^Jp@!	S@D/5ycX+Pz;^eb#.bkVdo(BC+aFQ^AHE#o]znP*G`"uSMw\MT\|bU<?b4h3c~Y`@XeDwIQ:("4lPkM7ZBe

x\=Q7`;UH>oSU.tMJvq$0*"&m8Jv[x/*eLT~s;-	o|G,-N{/OC/."<?Wwn]d}%(hmi.;L{Wqy`4?E8Y+#vWzA<#Zk^j:P^@OYE/.$/3[%hx|><=qg	@NR#1+)giWnD;xqK"8HOT:44Z_{H3`j09V62$"ZT
M4bhm&a'YT*0UTv;pIMBG#(GpLW	 4sY{}U|s6ugC|YP6r%z/,.3>mn/9J|}("hLN${U)Y5~6(,X{\#8m|zZLxwqJ{R]2@ma^7<{>RBR,~k]W@}OtqDxCB4VDV@V,ZYd0Q}{VP	lhnwNH3&dV2SRvA7M:b<n^2-/F-.4	^|T*gF|e#<o5>5*M"q>!>zf1=L:PVM.DDf^`CN{=A7K7`V/`1*Q>_U	XM{Xi~HXzlEo4N4;g_9h"~dx]Nou>oU
exPM,FKFD"Mz6mslU:|a>+m ^v"oOG/&/!=.gP5w{)C:^:J:00RI)V-E]4r)3NaY9.xhD!h?#i	{p5u2Zs5@4p-/e$'.3hv>d|tJwXZ"MD:&`;b`H;T$cf}2_V0>.=#vlQT\'1s[93AzZH]q,x42tla1c+FSFb2?#U$ji`LUW[FqKcX/_Yw4LQ@y'`0>5a&AKf}0wYS]g]*N*Bh:[.fE[H_Mmz%f|Gfm"D&{2`%4iIIiM9P8?7 E{/Y]$BrZb|P]YNW^]}EtZyxKj6DDtArCn@W\z@U<KDR:!uzlXYJ`Ua/{+Eml?DC2uqRKu(,rJ4Y5bHPpUck(Qk%DgBG{!U1Qre1}uD7cAG*:2z9 cla`jN->C4M53[Jg:NyqEiTJYUS$jNOj^kP!&ta]j=
<h>}p9KTFWGUVroy}jrb=xqoJrkq>L;$*i-W!;yAl(]e+WUeU&7Q((1pNH OY$SLx<sMOGTr>T?FN7_AC!KcEgM|L/-c2yGk2=y!w+,Qs,UCpj G9,ez,DrNm'9K>?.[9ghXGBx$!!L~.S7?6pLOUmD1&tbn{tw RQ>3RVqO}{Bq_Ey`uK=`jRIs<
xcSOd{{7+OAy k_JgNLv9$(= FINtN<2]$chu7=+c
c\E6)kCB}H
@N+>Flu9T5'bwF)]nG}s*tV*9P0_sX0I	&UcgPp~'X>0[$nYJJeM\];Qa8Wm]`a6EOmF+)I4:w/=Gs	ik(b_VsLMdQ+gA#:ppp/;]jqR(sf5$I?`_'kWETX/ItR\G$gH)8HuO1>&Z-)yw1dq9\U}}pQ9h^.kmitNYapahLAfXBA;lb:\6#QP[hvw}*U[~nRrV1D-]gNeD"Kt[f+8JnKCjcON/LrN4PZ,~OG#@Pbv)r!13SY13yh~=tB*5VR2Gt5idUCeT0)
)&uyG./E>+Ri[&&yKOHIr0J_Ei&L;o0jV5ev+e0U+oJV5<fOf5BWxJzuAt|	c+UfI7Au?yo\C%^(l1eYB8I'y</q?%yd-%9gHl(Fn{v;{`T
e/q3n(oNwG-6s1*`lp/xe>w8lkvyeHk'Fkt:LAT[fBTSZ27x
i^ps*dd1ZPJ6xn*xu^I6\ p{mhU9Bmdx{Q
0WZ"y
?<J| (?HfYS|?c{;tjx:3TP^;O3(M7i]OLu?"k!e[wysu\WGG^o"GC*42L&7Uq7jdF/8?[f1[\1J4?xt}H~M4pE)>hw9h5X]w~$6};H%	=
"9Bg4[P3Evv!OP\CLk6vaCKD=c>j02x%kG7Ox6!fC(YhWJUU,?d?.kA$8yiIR{Tc9PPy:m_Kbet!sp>D1Sg*_'Ssi:TB^GaEz#WvB&-_klL+"a>BOLB
Hd^{\`?VPTHWcA7}c FlDJKR\:DBn"A+bR*GOy%dw8-{v^Y1aYb/w3dWcmGT11^5 mWO<NZ_Wkg7a;sNhFYHJ,991YR7#AJby	hq4+;XW8i]^JU!~'}k5w{WGE0gvdJP-&y&mjn6:VSfa8+RItEl8aO$X_4JkU>p5CF]""t:@E~il%7u\U)O+E^%{z]h<BNO+V+qtEu%CX='fc,25f7whSS'Vnq=M5^H'@q-7z	8A$= 0<IeJ?|?NfWl3S%UQ?$vpv"D%ST<?hc<5R]H^2/V~Wg7!mT4c!a??'w#mf%x*-rUvItU8J~V9sB
N7z"v|Hg^|OVXKwTn;kzm0rY$C?:bLfz5iI5S+m&*>7}xd>gd.6
6/;&&#]dT`3E$!HQ;BShK(r	*{8#c?6)ekJAqz]UHc	#?(~=I(j3;DJ@L+RkUdt|v)6X4L4#n
Sfjo~GI-[c@A>Lp"ML.G;h>-|BPq,h^SJ1|MiT\}G4Wm?=cI!ek,}@3#z"
&ax63`AtNFN+v<@p_/\+swTY{/KDm/Rtjl!k[`N@bwhKzg3B!i#fQb}-~ L'@o:m0()bBxtPNYURqh'47_yE|Z~-0BFHOxSFtH@<\Z+wnJvrUo_|Q)xl!aydl~iEFI!6#eEMB$(LU[2753* 1 4?@r|TrnPy[ajHa,K
"7g({t&%-nx<]u}-Xg7"}!2JL~:X'g;8}3F;y\;SN9t0v#+LiWd8mRjD7*k*4^$M"tjq&wIbN\UkJHZd]3K*3g$6J_r|Z/HWco&(R+
vVd%P>aG??q C0eoJ-Zv}G_ \R[h-<_\"TF1_S;dts'P`iZ=z1d~.}|qX,4PdSQC?\PK:?7<itbIv%]shbs+p>./Xj!%JIx`4O	IK8(11W@~[cAn'_|,-'^<GdD*
DArPM_znkpcc;/c_!j9U<^ZBg0K0?L;/	bA;pY\Nv	3[9).>EBNMy860IdytTU?#4Q6O%!Fh(Sy8(^!E~y"o',%E/3(gs<@~	5v5!Dm-iz5|9cu:&/KUKiF2@B?r4#!]2iVq\E$r,]ekwpAX4c!<Eo|/lWiA\blP-UZeFRRN:)!1qeA#&A5Mm/VoIeIbE6]D6^6:dBx5v:n?/CUKW0TSvF0S,j[CPp[>"Eo[J$eHf@]%#(<Z6v/f?;=;U`lwtZ<sE6.ivXSRJ=I3/ToNn%X?JAZy_4@2TVh~odQn2>!;~8G[YlM#tv	\M._J*3Vl>h]D3*6fQM87;i^
+#`TB[ aZe.#I%2;N/)cV2rKErM\^aE-f3JP3[:1!9BadtGF~p}"gMAh0p2t;y	\<+=Q|h}6d;14c~MA7:Tm9_;yF}_X/&H>#?S0IC~+">m{Hul]Quqsr>$R++t(B|v2:{r@;5tmOIM)t^1@{P|>!B;4A9we"#1Wy$:Nw7lOde$v|o:_,#u>?s`~3N>,1Z.]LNFG>U )5.<(+<:?435Y\W`A2XQ_`zy#@0!mfo=$9*[+Mvp2>-8p7z`wDq\-p#Dm3d`z7J1lUI1&7V2p-fKU2Y;ir#xi)d1
a+nDx^I(o]=tmKw,m9jFQPfx?Fj
Yta#\@v^>>hGx)d[sZ~mf_]/KZi*	jE(7pTN5/8
&mtfjtCVo.S?=)^?O_MlHoFQi'0|woKQSB{E_?`pLrN'`}CF'Dk,wk`&_'U`%f`<@k-N`A"0({_559,B)mb~~!Gr,R!xY#stccJQ[Q1M9Uw^Z	}p!hd*tH~A*=zK4J6hYK<?Ps9c4!#n=wI$4W?75F&s9S8'8$!\{P?|?pFzi]Q!xD;DMB]qw+X8LNZ149("Gfk yz)8V8c('n+s5B	@+OKmV&PiGC'!,=NAnN2rK]%n5>"CF'cdJ+.]h!F;!v#$8k8B4YSq"V+S)mncGFOl'RcMwu(jPu|2CxjPIl:Ev0y"#-s-I]*I5w0y
:?	#.-v?C`I1M1&16KGh8ySeBxl[+xtaO.%m[0h-!@XSsrch`BfxU.8yY$[FRGf(4v=VT@l\lBjS	T*K+%Vb>&$P0sweJ3u=Azl52EEz[zn{o$*"\?S541Lx'?+T7}wX)<qYkb.jV	6-xJ`}Myc+FRpFK.[Qgv/dHK>269<ag|v9N+P$KBbm9VPWWHifN\B}GmFr/wNq"J>XBu2LvG`\v5xq{P#&#C~'yA]^PJth:NE-A+ale7W^>{@Y%"	JKTz_Jl^6xfmr"w )xmyu2%aq+s/Q')c-cm(a0izOLx
qxw];Q.Q`C
Nb9n+@a?4=B@hS=<|}"~)'R@Y-ekU%J{2MrufvG,1r*`QoOrj?,3'[.4|%/KI}_ (eCu[XNd@Gu%(N/duLB^p`+.H_}7jVG9^d?bT~]z]ue_M+>9`Z2a+&fL;\{D5@g jZ^O5&c/MQm!{8rs*mml:F?tq%giS f}BOK7KhqP,`5ptho"oc0j7cDS7=l,!zu:>zSq+yO2phI(o6\uj.WHR"yF:ys1?lf{}n2Ja6^@1&0Fmq[dRa\lNP:P	:r^0y?1	$&KX`!N)?tk&	LWhlM=SOyBC8-$'7Rzb{A0z-((+^qI1x>d<(?VvyBt#MBFH I|~Xf-e+~zfG].\&(Zt70eG
U_|PSmm=T2sxj8`vY$.f0y|!b#,OouS
%T?:J!0Ng#Rl<w"m)P8LG_kM.^P
**>&Z>gw8%z(v&#j?2YkOILH<bxZw9{2B>]uy!~kj3B({;>2v,xP{)M.`she	9}MEGS?Q?'nD,aW
(PENS6_3L1V7dyH.*=u!<<L9R7b}D0@KK8_!ir8L(	kqk2_gCn. LBA:zV!c\kB[83HL>qesxC2^779G(Y!w k9RQ0r\q8qfJGv6fY&0/iMr/M65J\9"y'%M}b0Hq,+-W[0Kd09lH%*B]bo%BGmAz0)|m"924;^xi`7}92:Pau6{EdQ.'APY=p	T#^s	fxx~oVItN:E?Fsy6ZnicOx?EJu}ea)	KZr`<%xH@qvu7AI5GqiiB8-?
5J/a#"vK@qL]Lx@9n4b1(\^>a]AHM=oD'za%J=/=LOJ'"GmZ]( WC;$hYNp@BhWCPou99U?~0BjY9.iT5l4sw,	+^nU	3Kt
wKi4M`8)d
}hU'/2sB,\aw>=-K1xS>${i?<R.?R)C[+w<Ryo_Y9KTo=Y-?/Q
6
@+lf]3L9UKlxp.K:ney@v`t. Oxhe,<u#bH9X#DRQZ(pv'9]G4w,p2x<bcE_IjetW8lVQ4uU2TZ]Ad@;L0gTl&D\c~	D9|:~N"xj+)vogae868ZDWnMdI/Z~!BBU4hQ8M.[D(7R?ffRxKY(Pify%74y^w~j,"T)"a	2p;Vum\{:\/^dj-kyqAu:!l<eQ3pX{=T>[l@vYKXX<`1-e,k/G:z}n(2t[)VG3=j>oAm<Le;	j_UAN}vl7-|55WYQ<[ v:_j::|$%"v)?xx/^$K+oOUG(X*}K0+oF~Re5K^hrELK%kVLUpvaW'HV@r5],F uFo#Rtld:leql@FKIlJHpQ#t&1;3*GP>2o8gQ^f
6R,k )BGxhY'/W~EYuDe[G,C6])+{yr9(#<h7a|N@Z@0ar.MYxPfCcVu*g?`K<z!Sk{lXkqb)Z00BnZQJS,K
}MPLVFbyG,BVe-6|)\4r/RB&Y;yAbv|lg	QN"j~iW#sFj]_kx}NOV	~b
ULFl2Ttz=?(V<v.Q	XD%gn-FQHBhzE@rVGzT?pe?kKk;m 	[*o0}dTSXp!B%[U/6oU	fG]-,CM(V7q-wh[&	6= fMtI1,6sIq:aOd*ZLxGB..!r?a&g*	%*0J@P#P|7[-i@G1BZY?t&S/sfU"Mzp<y(F+CCv(NO&Q]Y4i,pzt$GLwPvt-9OF+Y}K%pvson1Wo,v8~	CDU7L2v\zI4\LSJcTsTQ1Iw577P>'`B>1FcAG0ZY.*}:UIm,HdM=:?hxz#1JVS!2*%iJ7GGS)AZ~EFy*q3-/jHa~q=ktlC=3Wz|m{9TJ\*TY"B:P\XWb#j<c P8<9hGBC8&;hRIvZ=>KNNw^idGf	U1rrau.kf?v@3W\v1/E;oI)dv-@]#if=+]0o26d+Zh5Y4N.[p Gj''N-+]66^+.{*[{po5{l~-x4!%]Xj~yD@95LC
]/E`lVHcSDNF+BZA]~)/d?V*0VknU=Jq1gk$w3~8U]hf$Sef}jd]z4#ZMg/1|{k|8mTyJyjF2'1=@aUY)83"Rxld&eo^C*pUh,?Rv<Ri|!~L;ZFzW7Rq]TM9$'q!FUB2k	v$hrIr.))>siv[2,1Z0E*$jmX2WdqRh1}uhVKnx=b2=oiy#`V3SKUX??PP0*0lFT,-Vzx7)wc*a8v_Je3?Fm^Z<92F+rR~
jdBZZ4b\~\,6mRfaG&5Xc	iEsO,oI.F?RN*5Y6$*/g<|3@!g@$r_P3}ZRJHPc>:}\koh$vy'Bh.JQ$FnCj7H>0=|k t4k* m_qT'w?46P=jn9Ek
[IS@`f^D|2XL*c@671v@E,dBAuMbR!D@D|l'#Gbh[?}3z>3uCN;
cUm7>D_H|g:n+#RFe8T`^,n`BeE-;XeNJ>Tfv#6%J7vcT/)Q3kHkMG-BeoemQZ}A@gs*6)ELgRJ Ch#T_c.9t:6tW7S+:EXf"0iswPP(3ppakvSv3X?f,$ZJm7xuYhr3UV*GX7N`:`@$;$cUi	WG"l	g@tyx?FRt-{14jD>(sZ-X7adA3>arRsls(9&N6&w)>+FCld!gN!s3nI4Es![\&;y\dtjISw	7JCw&jjJ/fmo\"".)I<ur"Zk9H:gSdv|WXP}=}Hn1LGmvNd"e0J8
{[(#-J*+M)}zjnc@Fc`t/NM"-g|N+Ov8'tto\plNINq|m!a7$j8PRwoi;@QWXpD.n$"i/S:Lc2Yntz:,n}EDk^,ZG4MT86=QwZ5ya`r8XX&+F:{-JOFNRsJD=g#o<sP'L!9K6h5o!O]ZtNVRbI(=	Q%Dn1]FM3Y-7XnB#OJ#!n	4mr@81p4@,,G8Hjj@U{t?"bC8ypLpkp$gTsFgha\^bj:1\LaqnP!Ab'Hi
GBhl2Gf%eZ@ClWhTR3wG*2YK#(@T)=A>#){3*kTh3e(C3QVc#x_2yY*,VCrfYe7pjy]UmT]c^b3*qRh]NL8lU%_kV+PYE<{[QYm&[M]q1:&ZlO
PbTvNq>a:e=7G0'yc!B[,uA#ZAZ")@y\
3I9+4>CTvO#([|&0>9h=8Vtp=:"SZZuS|9)DG+ \@rvv!H?z5`P$ATau!xTBB!;8uw<D=LITx-7zz]-n%L72r$m$:1?a",'YD_'%pHpRJe:.^R*|m&^7*J@3sU[r0H5<RxaoMRd,rKGX	2;$oL)Q?t`.A.EANEup5GB}NYMXlS6-@D|n8t}#N[s72l/Uf4Ls;J}MLbzO|Vv{^sc}"}@/viu;.HPihU]}FuM?j&5-Zbj#|Q?//bFgXh\B*}mBWb/ZyjaZ21I@(aWNeOnsQG :Y_H`.t=QDd )P1ABV,} >eI]{8V(ghpa-@dlPSIWdn:<{%7n'{o'@/tHv$aJ|Axy[46'+fJ@Z%<+UE#3lMOu[)Jbf(?$s|d!/i@%Z|v'P lP,Y4{97Y8}FA0/Q?W&8-cWC91TM^PJGpUFe=crWn6?6$SMNY=2? Z!C4@alK?ki#=w4uteinq)ndJF<->2jrZE"uQIye2YJ<<rgm5
H;gD
^NwYYu|kCi9[BR"s,U6@}
i,~3ZL~nKB3[Oy eP).F,1pc:>f#SI (Wo	rBSv%dx!"Me9b}3GU>Nn*5;0F	Sc@2xU?b7%-c!|x\~8udHTF+|@nbH(kpOh3,)PjZB}?kXp^Bd$;+5/0+Gc
7Y8HS(y:9fx<~)R4&o3Zkn9Sc4:~; 0?eg,iiOj2n|25(D|ZrK*%xgtuYTsbeOC8	YQ:_fxD,&93lh7+c@f!x8CEAN'i8&pMzL<|m.bG0rB]|:)6BU
Ehk{d"il09@1%Rh$Q];yvk?^tZ)]|kePU33x0u%1`B0SdLP\zBl!]Z\ ,e8`fvrNm-*tXRC$+Jr
iJpfqN?Zz
@9|w|h*kV06 MXC~:s|d5'UIQm/{Lh;)McXCCjK?;YI2@}g-,b}>DaK`2Ere_P]]Yygldn:Lc.4IDqNC]+1|(wA_oy
1t`rpH	,fL3|$Kv_tAQ`[7^e}q/$/&z`r-X\$n4WrvJ1~0!tW(#%;z+L$WHBie$X;RB2Brh F3hp49WCTNR2|.$jJc.ihV~Bhq3<C0P'65z`D1RPo w>
&h]('$Hq49L~ij?4to"O?"W)mDRDxDJ)jGT'I<H$~w8:L[/Aa&GjDx5K[9E-3g12TWWp{e%d4W!^uZ9c?qG9;2JX7yFl$_%<sb+f_'Q"exs6hJ+l#4}w(t)([~nLlM7q9m.iSNQ%9Po4$4P@,&dSNH2TCCX\o2o]mB}j9-"E(	lI:!(F5/lKIwY4[	,WZSK+Jyo'yJzU81SBH#Be&\Cr5M#ObOKWi,0MW`z\i`V1uCJ[H.^/f55<Q(1:;VYb*R]fV1_>VXTZQ|8.z@S$=vk5b]WwE0%g=^;Ez\!UQL{xFHAA#Fzo?K!Kt,o?S{g7rAL"/5w_ Y\Ufio0@udgw:`G;lh>`UrV$<pQpv|@+; U*V$=HM)sa>hYj8*O4=;V-o*KGJj5"zRx}dB'`dEIKLy7X3~epUMnw	
h&AxuFF"'I-Y`<)_TW+t'/
hOcr9br]",mJw|h6URi"*e'u=d{Ovz't%=;<6+_\3&,8{	+y@SleThsqh.8rW63Kb6oNt'%]}iad(?Cngs{*-m?O
}
aQ`^1az}n~De8Zl"RXfkVfeh,Tg6e=>8?ZM|sR;~,%f7 9C]lXmxmS~(MYXX6%+63urU(J-!]Y:Wj1L.W>vjW&Cud,q*9`d-z	dNyjR;9[,fF+GkIOf>:	[CBgpRt+Za>M$#=UYq2,Nj\+8Z A8o{+cQNS0?5J?,:rns3Vs.\RwIOI5D	PCk04W,5Y,sE@?{!*ky'|D}8D!Up}9)+cw+g}yh9NDH
16!>H*kuZ0}nJ7h|30["57_q	$-ZjCgM2p^.4AczUx5kwAPT+( iVl$g`!Y^KHkSP%8WDKJT`MD;#U<mmXyPIF9<=Y)E@i`dt7t&%8eetDsP53[nz\^*S;hy(Kg$B}'_VE73M?!B?I^J?zVeR[.kGN230!BWI4SsC8c%H.]IG[|raa_HC2u[PZwrcS@4+-l%:L*)\UHd_-BX<1>Eg>3L|y1.2$S!I$.}-]yTYb2N39W1}4}-+rJ@s">tT*#&*9?x(,a`,jk;Z}axvU'<.\8f4>9by|;p}HoQco;3?&3WkIKnnQIo0{U&n:L8y;r|0YSf!_sU[$]7:3}z{C\>M,SZ'IOV!>Fy(7{S.
d rh&U<zK-21Q4}PyOw@Kp/<my:#qp.0xt}:_>uB(w=1AZ2;[
RH`5$	{.[@	.qybTs.4qD	,+}=]urs:+
skr^!kAhpYaq2&:;(	-ccuruPrJ/@Pgv-NEN	k/$5BzOAZUBbJln|PPl?OUU
o[;@1$eB>|!`Y^Z\\TGu6S,8dpQw
;,{!+M#=(P2$Dt%@,gzGW{e0(_a!2r6y#UT!q9IS9m#EJ__aZ$AyrnR`6s/z>TS=?>E$jpC9P} o@{V!4T4|r#}XFrz?>T}U?SCfuc@fLx9^9U'TE|3_*%hzb{:aG0Wf%f(m./^sgAv\*WP9"E
.[ToBep%}ENNQ~X'/xkoU.~*Gm3KAcg)trM3_ou6rA-Z6qum7~;KDQ]cB%5/FQb;
_}3ONl["JUWdS]4732,yS|L5a1iE-LC	]Ul[733c?"}*O17bfD#gJ "_s^iPl]_	wft:O9aDaz/_6>AH7wi
ZR8xk/];FG?FZA@kjviG{Iif.*xuzD(QLRRcG
JSH^20S&OA?Gs/pEK{8Cmyhc\El(G%^ 7J;Ze0!Jljy;W3.K0~mfQVM;"nD65:}KgdEVrM(jL0|Os+f%m$|`1P5y`QBH^4PM3_Ol)Rw$tx%0)+dq?};13*-e@X.c	\pU3DHh2\_.0If]G3?OZp@/AD|%G5Zbv^sz}::-'_fqgxUYXYa;$i8KaBNvDU4M9oMn<>X#<[0>Orv+7Tz>n'#]Lj69RI]+[~i	wE@=zIl0P^wD3@4NO1$s@>'pqe!]&y(}&'A,ZVxC08Co2}.;l>,h}jsPU.
<O"MF<4"5
w97Kf/[?o[=2?~a9][~UfiH$Kg3"oYu?b^|EJCPz9q$'y]BRN}(N$(q$i*u|C>^=5i0phzUv2G(Hz?wC^'jsc+-0E;u7.,y/&YCw4w(kN Hnd$,3k'y<O-[_-",AWJv+h$IDx
--^9@{VF\=rne}?b]wF[V,"_S9\!uAHXky4JGK2-`ofx0j9\z9#?aV#oc9XQUT@z/v[~A^12{n|3`_AZPqv]NH$
8gpAqx*.,=D@D^3xMHhA^Fq>0%e-itd{D_/84C3E|,K2"u4@Tz6`F^FgiI/A$Sf@8GF%kiQ5BB\p-X~9sSB?s_H(!`V^U-{r4A[+sV='/J>NH*/*:+%LAN;MJ.r(Ffln.D$K7t4'|cbl]X=u	<6FA}f?vz-jj'r:[{	lvSb.	AV6fp`zMfouc 5[MRa/+0OIc!)@cQ'z+<@x<Gck`b>#.Oe_xo'	@l|:U2t|i12ak5dk>NNc4C /mwk/L*1bxC7%Q*_!=eW!7y>%xcaWqcL95U7e|	G	W)#t,R>p'pA'GXpu"	v9l:W:4?3he!I+_C9JP.yLG)1O!-BTF$h'$m)}|i3M(%Ysl^D% 5i!hyHJqMcKEOyUzpbU_?'5orR*
i\7Rg
h'_
qcZwUb*yVSa)$PedXVo$nAulVd7~*$t(}IbN{q
^KO#pgN 0@:rz`)W;0v,#TNNNFG|f[` h@;VSDXOW[q}yM5)t2H$E.
V`9#T{tnjv`ML=Y'"n6=TaW)WH!.vh?
m2zBR9{:cMz&5#mye>BIvci`$P{|)EKY'S]\s8kSSNQ3qF9W|GjD=8]-:Oa!ILAw-@.QCKErWqmt.Q	U/`8[{+'J+bnn_bT>s76U|B;{ ;mb'3IVEJE|_d$%DP7~|6b@~!qCJ!:C;Z;\XJn6FHAC~1]	;dsI|(3eI]l2rlo1C%dN%M1QmIF8B@~[#4U0L`{fS^gy6OOoOmT{""I78i
)8IcB2jX2[lhlrQ\q-.!k6@dG4]<sJ)[JyTy-#'5NEh='FXY]2jDgf%2=0xdX]\z
b?OT6O`++rfx}((nn&joss:{V<".>UmEt?&Z
A5;*{a&-n%*QzbF`0
.'V2|Y5QvoUVXZ[`ZJum  _vIv!mM:~t
G#xxtPv;A)_*eYY~%c$-IY3?:KK"IEY)gu~:WR:}
]*HQXG)iT#$]P]Kv2t&,66,`qy\].%fz}p[h\oVg.DQS<HTBy[v 4j-Xyf
S?fv^	W#=7a;jvb#c3/Ci#N7u_gRZ:T# Bv5cTdFq
kI(dk.PD L>t=_*Nh7Nb+#4m;zXSOg[-)^xNkqO&]O3_5rd(3l{QjyyVvYz(O>x!NIAlfy"-f@>u-5\BK7=V`;!\GB#Vg-^;6)8SX[28	UVD">-nRY<!Een|d+OJK
V}<f&[4xa/YEzaM_K~	!t @1GI9GH"tx|[;u",K=r$*"YS)cw9-fLTY,sV!Z;
J`w5~Iek/CQ?^nB@o8hdj!P+LeORf;:*Lw!NtQ{1;mNBGrHV^$$9vC\E)K]]EmhA$!}96=M@bdg7`ik`u^GmA3Aa3[ez=a'2Bt/.HOvIia0_%,fGDVomk+"L,sXwl&^aV]2b<P[a[/gTRF	~hxD6,3l=<Z<&Ouh+WGh;cms:j{8;^B<hSfDpv]>I2J`>fYeL:E$U?'V,s@W)TY%=Af~{uV/z6>:dcwB4-"sx72TtH[}-[55sn[#>IO;!&glBmNUG_K1[}pqX7.(AcX3?	KOzsZnAqDo}/0'f#Z'f4h`t0-AfH2bh-.#d_t`?-D^F6/T`6Abb+M4S>xc2@IxC80mPJh7<M^#M@. %#/^J3#>a34|4hY}~hQ1b)o30+3?_eC9O&pJeY>x6m K$]t3q7D=n9hhOK`x>xi}E5|">	]AAj5\8JufHl8*?P_0s%dHaKv~SvDy[R=|T8za;28|s2p( oVXgV*xvmc]uWW1G#Vd[bo]mQ:%\`?9)qQxn,eO4&LD^fzSLY6N|oa6="5.IHg!b56o_$e#5_?${d7t Ks$h^PY-M8_I(21f]0{	`fS)w9D)zB:I-=`yV=q0.?V!T8}D()3`E7dS	357Hs*@R[HsnuQ:G(&-N
4hb#tB r=L,XH<CcaB9MRUxUdjod^ o !pFb@,O1%PcrP\@u7R,Nd
%VaQ{q^h+lV6OD^\2T0d^8$?qO.*-C 0h%
/\Oi3-6[FtgHgu1Y-a=lCy<8rTO.' (We=4NirmJ<:g^+9dRe"Q;^`{<g>s7u=m|X':8X	P_Nt?{'f(#>nREcmm]"_4HrtqOpPQ2~rC@1I-6W:8GqXD`)T5f)\|Wq}a]H^_8bjXsL> "?*(95smpY$ojX"{E[87+p*U25H"e4tCJK^p&NXJ]1Lqe=t_3x\pudMopS{LqAJ5+2o6SY%Xu*j#nD{C1LodfL4'=1J3R1sB/aUL@pf3(`11s8Gv15*9a;"NZ<e_Y=R,rZ`V^7DK3JY ]OU_'V5SI)uBS	)HeEE4,{5W[{7R*$x%w\x,&JEeZL7}6b]Gy+]XgqY	d/gdq?"Y38:":S=LhB)3xh}~By*}ctgttlyxV2!nxuY;:$6|Qi,5&$qVtFuVh:/?sIQzzf%1^zo6t']=wiB|rWf^}4shy-{`
C$&vv"u/T) W,BVe}<oK8j3VZ=`eishIm&!/3dD^	gR6Xu4z9K_><M[-B
=jm3!{ R]6i.XJ9zi7Rk#67
He6h%d+}KZg>Z^o0}|_*vKoe/,-J8H|>1BsTZ(! =a<\ZB[A~kC,1bgoNm8O/5k%3Mob[?Lr=OUtge4r&sDd+Jw*H$8o)~<F0|C3[^t\M	"0,r$;]<QaCz'1KroJ4><YSdAju$]D+{ S!Qo?'(PL`%t:f@;WZ	^/BXvSh(XrW,bKr_B"Ogkf>O7f8>A<r>|",=U{X^44O%prN4_k>J:[|L8	"f`@j{z%rzv1R8(>	NKC'-Uj3xebc(s{*7b)=.x($2n5[OXL'8^";IVZfPqV8k=Qh_DE[dQC<{zv,ZL^)F%HH
W7u:}T@r&lEj)yUU:ol0Z:E-shwJXO3{cGp6Q[lG=-?W''5nX};;,8dGPVU\I+l[-%#Y4u:M?BM{aDQC}	x~
n:^;Yl=O|Z&d]54E[WbWSmMv+%8gRPv@b+$[}uj[VVoW9LE!v$Y?C 9KzXfaj[V&*,9]!T{idgg}+(O\E?nguOUFwBfKQ$!RYutRTtmBZ7zAL.zE/ahl!y<}``7fAhP.``MogmY@n"vuyjZq(S23i^oUP
SlNdzLSg%:U
2-9b:+M' s"}T*7AsiLe4sq
,6svi_:bo[KzmG	0E&9

RC	0W5QMK=_%.	?PXQr:-qM=aatL)60`Hz kAy8YVD5|xQf9,&	l8mwluz5WE\P)=^pJ<Z7$o@.#g_;$VGPX2PeSW;c3V+|#mv!kp-,<~{LiVx}NrEb>EGN]>>3e%S+X!Zjk"GKT&@EeW72rBQLo*E|Ig*!``4j V/m k^	^w
+D;zfh[I6AH$68>W0;X``5;{	zEc;Z&W:\V&OoN,^R60wo$@>JVL7;i,(%lN]_lA|><{BA,.9y$cx7RL|nN@nqRC9;2[No\QB[f2]Hc-u]?r1E!O[ 8?F*:BaV5n<	E_dR7;Z8#7A:sB&yWrN7u;=|&Sz0Y[|PBC"]"pcE\ndR,$nAhr`74CacgXy&suEtV}`FhvP+0G<4H%\5eHR>|&{pzb8g0COvhLgjBQa;#/2[uJpqu7!8\fB%M2[B{l?vB:$yC>LAfb[:Fyl*&4J*mY`##c}<vHN@x@{ t	wEA=?'&Wb?'X&V,E.r>vUA3y~Te1PIIGU%j>hU?bVsNZL$~cOj/3N^R|O	`Ci9F-eif?r}'x&S!D\_Fw8'N(^.fY]OGmLPftbPszn!/){bk{bQ)J
I~r_PO ji3(N7LQO3!zD9>u9n&o(:(o v][I"A<iR*P%}t_|KBHimCuW$a9a.gz3[Z'>C\;&F$UI1AOA@>,9uv@EjJIGoEe"nb7@iVh@{1U$/.FBO~?I
TzNK%~)199*J+<"-.'m"phBdU%T@>Yg|^a_xj#j4y76E3|Y9;:RCe]"Nl2(,Vmqd~>LFN{Mxo|o0?X<y3b>[Ed/-?81!x8"Mk8O$4dUMDXZ
)2{/o"f!
WGZTknz/1wp-x;Q'>:<D$R^qCjQi)~->#%XHO!EuicZRX7[8lK26"O"PGy`ga/Bd9^AT	(#v;7?:Q#h Bk!'jB.{&lULjh>MgNQ;+-&XA1uLs@)Wc>t{}Mu**jekK(#ed2>DS^aRSKicW:JVl-<NFK-%pu<a_VNA\$;%0AJvIi}^=	b46ZjY8 vbPl.:/+~ZQ=!f	>oi?ym0hv]VYOtgE:;?-cy<`D_z^#[~9))nUgBX'e5]XrK2*d&4wMh<,&XQ5J6K>n^3v4]&G6ti{"S	Y-U*`eKho
LLJWyx-|";*J\SMKXKL(bhs\2e?A}qi+Ok!f%6A{QE"`1

Y2XRfVo+_1Du=64-V22Cit Zp%%v_2:BvgyN_9iLFWr
)uhM_(gU-&&vVhv*:\?i:>BvF%s&Ws3}.
M#NU2a/=aMuvGC\47P b{OD=B<KTc
>g)	'RPQx
3ZpNdqbY0eMe<MUrC/T9w<	KHj&YDi4`-#F8yK{DRd[}IO)XD0:"w)iK@S:`5r_"rMrtS&CR3QvB$afY}\]Sh0go^7:<5\dxFk&N!M5u>|IC
SOl|w!v=MOWfx|pLkpf	4v[M(`.C&Ka9%?V?|E&3;?.~7"2<S[/WwiSug*[e!Ftw3NIng"f|Jt1Oa_@LTS[i"|8:AN%'N<*z)/01%TS|5ddu>6E_tG]oH${r
%(}+Bx"LMB#m|(iWze"BV\SD(xhm7>bt\Dj@m.?Y5V0$S<Iu3>($!*)*(z<T b18jA4y69!T(X7oj$-Ot6ZEIr)E,zRIyp`%|Su>=kfZJhCAn BZ5xQoc5S.|N25+/4.a'a+\E1M*9@xA|/\uQam~'mI_;]aRV8r35=L}bs6PJnSED_VK_[#)iHA|To#<}	'Qdo?|zd\16fj&xP0nd"[E^aW~!x5)V`o47D?2K{}Gt$U99xcQ5%g5:'!w<9 bLF9')$*hDIDo[
"cIxW:A'-!hVu<N:##R2	:7V>$jIxESoE^'iFBd`<kSDuCg(zUNeq(S\AWUk6o }GYWvDZH^`xj_\]m+b@>x5PZ~70)q8jZw&x%_?t1?IcJg0@:h2_$#m^<hv{)<k'{GU[U=AG jg72>(m	b5PJs oq2:U
Zc	V6T'(P0pd-DcLbQ6J9&n_&/:*w2IFN+N-c;;xO7RcO<h^d7iSVrSZ#X7ySq1$<<tz R6::MvGq0d9@<Bq\"tt,9WRK>+B5?-b+IT
G6e;YPF{/ E="42(fg}vwRe<i~LrQWmn{L'@6>6`%yf95n-#W_|!K$o?u6@ax^/}XQvb^9R^80OK%lN;CHF-{2W!228Rq{I?$)i\y'Jn-%EYNFB;#KzIplZ^=Hq=bTaS  UXa[>1q<!LaXNE
$d\F**o 4wtlLb2^jvw]9KqYXZ$D"QN
mpbD8mz%$@+K'l7")&=4 {@noLu{+Q%_;|R 6T+V*WLb_0S$N03]d8
T.$%-cyKAR2<M??Cz}<1s?,&io6(j{L>W~(2.''0r3mV]N(zv3Mm=d3soPcM&'i*`r;VclMydn\P?<"6W];W@FTUF/zN r@Hcn4I*>0AB7~PGz;ki&GXQdu.>2,bs\%s:?yIio 4e7)Z3U&=xS.@E"E$%/L*yt|anysDs{\0DB1
U[gV&<PVjn82ko}j(q/:OrU#u
i<FY7';TLgs8Lr *Lca
b!('$$?K1~skL' a:60&V9B%Sdb f$"^+CiCl%@i(mOD8xb EMiz'|?RyAv!9)uCR9+P;2J]
[.llcw!w8uBK'_6Y)d/^UV:|t.h(1-eC
aRtHaek4r&gOCm9BZ0YzS\<OXlAv@X|GV'5
/>rp*	?qBI}q+NT1|+I%vi=]H2;NI ANy91)d@5>\yDdC3iwMiy4V&Ic<8Qs)M-_az	UUHD|%W36O#[Tf9@_"ek:Ho{8O9Y@Vq_ 2l[D)2.6-H&(CZMm";%0[w/_}1X\qWv}qfm.5@Brg #,7D l}Q7x%'p?sUt@5W)ID2g+hV;:#ZV@G`L)..Yo}naJWZ
&jdM~\pVt"?_MCf~.PwO X-E*E"<4%Y_9L%Ly|yfMZF_fHol]=Tk+ez;BPPgqM6=qOusa]+qWCA&-uRM5d;DjEk=IZ<[I\d3)/!f\
F:ynvHZ9'>#P~5Hz#w{y2&hkd+eN{pB&)c n
~O3Q&H9p@\23FpDvs(c<@Pu~(7S8#?M0i<NL;Ig~b?B@T<gH!5"j{E$]1#~7L@MDE';0yb3JJ9JMF{f<DIB(dqwb;Pyh-@U.}DBuFBWmmC;kZXM\rbQ6]Q|zm/#
Ha+?5Gbi:u:1W\6G}rSL2AHa~aL_>hOO0"etSko~s_TP1u5_C^>]JwWoC;KAce^KQ;PtRJ:&r&@&*lV@5X+Q)!>>xbg{:"X 5%r <=i3c!_H>yzJ
7CP*2)ek}OII9KRCY0;w9u)<(@;IY%gwrx*{l=w@rE*l9)Bxm3Lf^