x"Q#LM4J&`;OYwTh~N#GW|N76M6t&X\:+g\ueK u0,
DTlPR+(gwLbY>;INeETR'Yj+:.sQi_LaN3NN<cAsV0{ agO8ZBaJ
N|yHqY({)3	'Tuwh2+o{UsleMQ%]$vyU7FGLwCTh.Fq#b6mz4<gz [P6f
/(1)I?Q"V	`
^Twa	DJ![=;I*?h0Ruu<<KS?q8fF<@;<x%?8+lgp'uUyHK2I<EnPirv"qD`v4*PgYW+)Xkv+[5[l/"W]
,@PyC+\yz>@81/0JAn?ufv{h+>R-x	l"zaol
K;Hw@`\i<O^
CM@-wRSkxp+	w3Xy<PW6W'a*.d,V.9b:nQgMSKfZh>bYeoT,n3X*am{C0Yqrcu<1F#2_
2es$'-HxJu3PUw%9.tflo3^HApZ,=N	9f/5%d0m)EgRgmi6-R>V|'G5,Y&[OPTa3}8=U.
wD58`JB`b2]<J<}.,2{auJs[vYzNv+xa#.$oSxla!_tKfQm?rAgL#U)f.u>d<XhVHWn~"onC1^5:0Q8DLq.vz1_Sq}+sSth|hwdox=I1yVV%sinD039q%)CZBzjA2%$tky+LsdoaHJp50P `w
G?sNF_!;Bq@A<qu_!v[bC
^4
T72ND=6'6q`K*-&UXKOk*i%QQ]+V$-lO rd~6JWx\|Jdgr_s0C4&7\8C}L&'iww%rwW6lX@sz7f$p #Q\ w79Y@)&Q.TpcSd[EW,;\%H(D9cc47,*I:t:;@A
Ns9dN"I=zce_0vzBAY>(1jVZ<(*pJ#
5?g.@Q	{E%:|9HZ4JTnTOj}z!Id)l>;Dga&^+[Zi@(TT4'i@f8su/hq}Q%?Pr(xV-Oo;ut}LxjT#2hG!uuY?0|+n8>UkKfF]
Xi]euIX-ZA)y$9bAC4-;jN=BkUr?wf_$y1(3l-Jxd;s\CV:+p9eX^?2)$-2dH\<[1BxxtjLrvnp]c2z+1HAnv),UD4FDjMuW)J{c_jkOmdB"4}|$bB`wQP1&iVeNhs^l -=
^zz%7pF T|<cK\[
Kr\]Pt_tLelZ2zDjZ2l1<Ft^{z.`$Vwf::rn"(
)K>*Eq-x0VxkGL 57_^MmS%^^(wp8J11hQjI6~+DN(q.z	'Tp20d3&Lo67072*Ze#w*}y:"+h^25yK*IG	SDg1T8?w,<UR<*#u `PmVL8y{^`-'=={no(a|_*"vH,j?e^!.+j]qJcL4po*%Ym[^w7@5$lOR~kBR`Kc6	w9/h04-f.H	Ny6zR8r|aWDEv2yUNiODNv\2U-a*3`y5|]Dn^yq_8zCS7l8gxfL+'7L:*v7cVY`HgQ:qy7Hks5gY8_'`vKg=>f"ZMwK*fx}&i32p6"Tw&~i\nTg{>?\4d'3fJ!Uk $zC]2X=#x%Qb+\>q;.zCC'o8[m8R-|iiQ?K9[-%[5_xnp!K2R8J?i<is{Enz3"w;JZ*}]&dZK?oTWdsVbb1e1vZ:m_.G&e6R,OA@F*C`$nN=zBy(#:_OK]_\*c5%mmRgCZE&0.vp5Bs#}:g1HTZ:!0JoaZGRJ_r)EpJ421jYx<\I
0a)]i)c,_-.^4Fg/~I~;|LPB(T+F~+=PeAmGGW)S^IHvsHh7	g)Q{%b0]n@2yj9|e#%u"x=(.1EHDm
>v$D\Z9]|NeLf^U>+!&f^ I;pN]T@~T_$+~mw(_Vgsb3r@L[>{~|Jh-:2-,KC)uo`#L=z	fn!8HLn@>>''6xgEZ_d/"[;(vu*]6~'Ax\Nl,?\E	  .i	^\c+-cg1QXYC8IF5OPCy&YiwSO*noUW[E\TA:E4suHh$^,>fZ[mgLw{8-+5Fq o*[ &vd+_U8/y2x=1&*Z}?0
H}"wm[&ttxW7
[:NGYoS-(?}Q?a^9>q&8fUe`5h8L-Cea.'d_	Zp=WOYVXBtTmm(USfs|M,9b_]Q0$/IZ070`!z<B)apv+;3izUF%P?FW=.<^hE3	C-U1`eg>a/
c(O^\|+O"bK{DY[(JJ&0{N=:?}Be;;ZB.zV[mspb\PX%3/(nxLYoXMr$h!`8GXt
a,qe%cnBNhDJt$YS QWR{PfaFtLgBEuX|cf3(B%#@;i}\_M^f2gpn	XE}&{[ZyFhM=2`<qBaa:jA	]^T%YF"n3o[<d~
L0},n't}J:X)K&#:3H>fJb
*;'6-HzDb7+#\bq! e@I1m56OU#V`i|{&u]kBWSrx-*	}i+`Xy%]7C+lca~M27YtxFTJvUf*(8&G7?/A\pa5CBckD~iX6>s,w}J!9\9"J
9'W~{p3W^~.<%/0C$:f:8M=xS"pKfZr{Rp@tAs>TE8#ywTo	E#!y;Io/~#$[d#R>-fPHta{n+D&T):&.#k*oUW1>I H5TIrs@wkxled<
E@4v{?(!F_J:lu7p0F>b|>Wd}kpF%~5d\m>rI<3rmtrPE(&qJ!6(`_]N"@`>i.5Pt$m2$x=sg$cRSt+lqvZN>b05k9"L<<<w#1@xH6H^>k*=zz'2Ush4@s8tD/ShQ67DZ-;(k?+=x(]]Nyi8(Y,ERE7%wZBLh$ 'VD,Qv45"385pXq-7>W}(.TS.RJJhI)_`gZh[.@:{(I+	L/CbBfs+6NyY]!	#DNKqKiY_tZCs=erW\sv\n?\]DuE1HI4_^GjG=l}4:q4I&H-p\nERr32;fR}<wZtjl.hLF=2.h{;h&d\G@{f3$fW:4Oz\%0/E/KCgr -7Oe A8:>{VQ<n)w:|V&G#q[%gP^5Gt1
Q&cp?S<yra[9~>0?GIGKUvIaeNz?}R2QSd\!zhqz<3A+._5zA)LvoR{`qP|$O5TOk`
UQ;3i(;/u0>aE0GS K:Z;&|-6=l1>VV0,Ch=vr&BP41M:s-@,%H|#$lDwYRQ-F~_oJM0*6~ao%u@">xXu	'a9v1v^l=hx*vN7]X'b}nN>?e6Z'$\'3U<
"jiu.;{,PUN&9i`g@6lrywpI7j4>/^A:.g2l9pFCw*?oHE_V@"4p)xeRUe>YQJ9_J912SFY0s2TL!30<(Ss.x'|s_a,yZr4h1dVfcCJ-\{ZrhoqLIK1+!Xl#ol&~}W9Kp09Ip;^+b2P
|#G[(-]J1rut!s/jq=/8(I6N,aU:he$MO*1z83ise\8*1TM{XPBcl`UeeQLmw[s$<vux?^'EflqRlx!lqLvj"C.:$BkZQz(x8+zU`|bYL[,h"$9KEV )9LE\%#D"t9yk"{LX"l&`?iuU6uj*i'zhFr,id)IrXEn;|}-5"$GfX9fYVo|l+	5'4*71,z
`4\5l$&HXiGoo%2*y-cVA9@H'EbKt9QA_/ztG@`$\VfM6s_4[n \00"UpgR)K!uZx(9?G
<Z!,]/@$kOex#B@c8xb<#?3p|/>wl|K7$kX>.J|s8sj4mid^N4PmZs/T(Lf7e~vD(]F]Q`po7S}24oAK'#kQ-? m8J?vi-~V0*tE@TM&Wzz>Lo)y#Dd;q)"DH!LlYq@S.rg/H@Mnc75tc8,ocRERG'kvP/xOf*;=]vcAvml8Nw-5S&w]I\N*)4[~u`x))f)K,h%c:Ui+: Qd#o@,Oq*(=CRI&B7cD{4k4W@f	Tq"z,\Vq8.gLL\atlk;zy7bcdMClEta'y:hBM"OpIAP'n*7e}m6r|+Z'r;7/x3;iSd&,M</BB!(82i"Y<}iwiz#I/.[-Q	{,I/E.S/,<C>P1pqCb3?.Fxem@:&p-zY}krfxU{12}*!`do.7Lt5upxtW;~6Ii;-'&Kh6m_N^dSN6~s^h;QJgR';"&o.(MbG~HO?OIT?h1vFPm0%Sh4<+YAH=kVhV){wwjrmj	efJ9[)?AUX6Dd 8]K,=Ny$J(Xj$}p txA}2MzuCY]\13f?+1pSP<m;0Id-n<a:RtSE]9P '~'v!&O*;^7[]^(yhM@-%qyQU_h6kiXL\AkkCQHzXysCx1Nc:kh-`d2gP	L8U$1F:*'(Pt^gkD6@Kw2O|S#k[Eo)Z@?<}ZRBAs!,9Ye! Rfx,)*8UP`h>b)J44{nu&*lgy.mxP&<?]~3$Mzvw3hEAm +Z~X	s!(jNFNxxESVKd>b6%{9LO	0$>{R^LU3LQ:D9|s4L8pa!,[f]D`;~/45	mD|@2U^[WoHmF'=HLB`;Gl1c`Y#\%y/`DH$PsC}RPovD6+_;_;dtX;Ek5Ii>zSa7(Kd$yPHZ)*g75F?\;[pKeR6YIRP7,Nn(iUrM'GVy;tp>Dw{wP!r*+(^.#]jQDe;{`~V&XCYi,w>R}f#mG+9l:$EX,C=GxnK"z@`xw{I;HWr6\Vgw!_C'3jIm!H.Ejce]{q[$"bky{ZoA\BGNZ>?"FJ#u1`7B?t'KJ2OkYl	0w6c~'Z!x1g38?H"Q?]:As(J';^RG1OP)ehK),18]R'N67>{Y|B)F$e3E	M>U1+X
3~$AjdaVw"93Ob0Ca(q3LX]h
9vqFk.n u~fLtN]e9|U(xxNYB,~!"FA\K@8~eD0-'$g*[S8<RN)1+avIJ+
=rysZ9fBZgj4|nZSOZ82=Y\[:=n,#XzdPmVaY-e}%b
+axgS^Osrh0AjX|8{?H^x"bis>N@<~-(eT4T$
hPJ+h:)!.z=Pa4J,N;8:-tu8ge@C4]o]#Z(7$,5JGe5 S=//s^8,l,eYG|Y/$WaXrCoV5Ar(o%\)ZPOTwXn7R!,EOOWU4*5GWBHeG2j"5'*&-b[8]z8DEg,jF^$W`u/bo}=qz[/	Y?p9i:TEgsMIl89"4(>x]
"G{)0Cm@7bE7W[$kqzI""	}nSXM,%iCi?i8+ccY~G5[s/dv:02CU5XVRI3fyHK`BLemm*w<eK;%X&P~7lP6H5mm%Q6A_A	tMX:[H6.d>=1|#L{-_R;!'p5\}!a( nJ2BpaQPMQRKJO6a_Kyl<;Faa6=d8ewY	[YUqT]DS$W:/=YCC3Q/	TX_ObJb.s!B.y\:A|N%@{Gl4YQrT'WlQxCMl}4SJY}c8)>ZXs)X.H{A33[X2\: Hv/-BDa7_^T<Eee	p-kXE0XSkgB=KBLd)hJi/NTb'hg@QOfT^{ oAbP3'49fijzzPi0"3(*i}10:mHfIg$A|c~#&EnZsk&`>dNH5q3m0QCK5v,RL}CwZN4rK':&[#=xMXIT2vlQJxN>OZo M!>'T[8iZSZ0l(6W!U"8@/ JJ	N7"\coo%>}fr0H++nBkO/pT7}I<%^R~L',*H(']|Bz, x](hRt9zx>\XwkdlN-HF~*V:ui(Yx0?Ba=iS5).-/
CC,QJf9}En(Wl@$KK*u9Bw	e[H?}NSF#:X^MV`cL+`/8e*B2+ga?S1IbNfR)VB7M&3]_2=8/ak0L]qF2v`B>|K<o4aHPTY#jgf@=,irFsS1Jbl]y*'lNT7Sf5jX}j9Z\bvW	~+!8Js+i,:gfrLby09UtWN&&s)0+x{<pKy>06u`'=8l@6_(,\Od$PJSgkN:dcf9/gbxQ7Rk^lLtv!eDal=9-"YZV Ilo\`.So#0[K"+Nq_W)Yh(Rui&YQXx)"Z.&1AC![qV:r[}Y]1B6]3
q&jzq7EW>h+uf&FcxN0,S%*m<'k5Q)~AQf[;`OrT[1mp(p?p!d@)76VC{=}vw:i5u?aE9GJ2.)=\h=|"	:o{ZoL_:=VpLpwwv./Wd=f2 $|;3*RUNU-k7t>4Z&B .g}Boc	fJTV:~|z&Mw}K)?`Lc#my\V9f	XrS\"mM#k,cEA]b*7;ecrKtcc-P`}5y|!$b3>Hh9z
'eAL%()I{}\swWQdM;sv6Q:0fx|Ej3W4ice}	12znNf*]cM\R6cnAjL!9#Nsm-u>couOF)R42L4/yogB4G3PL}EkE_j35F$G(gHZu=35(fbkJ)af+Az:=Qc!NGtZtsL!W4FOR<*-&[YIqN)z`V<.L-~HN=:eG5F&)OxI6Dv1a:7ct~aR9<A"d"PW(-+Yq>&_~E&1>}(<i:o5\'Yx4mdZJQ/p=XcY\/<|H^+tC'G/vF#b>\y10`O=j]VI'<zg5`d^cs'9[W]5gobo[f')I&k/*Cg&Sy'*='3-.RTfYf=;W[UOmem$[2XpMt!{`::1Gi/bpW-43?I|8%"8_7/>s+_z[r0?A\c&f/E %-~i2<"1T<Ym+8UnqEZ3/lZNl>f8tpyH'1'j!p\s3EP!V{
eM	fg!7KZ]|7 "2!C%t3Xd,[
/Rz7w	To_1%:WR5C\5UK`ZhQE;Ga%_w*+Fa`Y*K^NRST;&rmZK==D58$95&a,=pYPkOSn!/]rCmEq6PME;xy3S| ?{pmX8;~h)tqE(* iPLo/ 4}yA`a.59|j?"sq[lz)h1LP3m'<V}Ndq/U#N[}pBR^&~b -VWv|I.iVQQb|!bdVRcY,:TB`A1<EO,8Vy>WX1ku,?Mud.XBaF_-kSGjX'X%UxmEtKxnA6+{,7]4vg#0(IHI@$oLzGCKiBYO20,pSyXKw*8uIz?q{A[d%Og7f>h(4]_-[00{ ]/=uVm:]<K[eJuwlqmTRHkTtci9N'L5'y
7!qM"$bP	[TSWA_@i6G\X]`:Smbus	L%ev\}/Ep37D*"h1<w)i-6|llnM8);FO/QqE*Gj:@^+`;6OOX8JX[c;OU&:*`p[7ZFFk3e$jz \0y3%rL2}'`$8vL9@T#Pk!}.(?}Ij`oapZ[M-O<ltQ1*hfD<\/Jx;57"M~vg/P
^ Q'=O]+aH[^@8iY(:wPqYD-X7i\p2cs$:n<nPCq[IytN9Fi!OrLpfV1	^ukHdr
U!"4b9'@C[(Pvju9>\q[5Y<G{e|I'iKFyMW'7{s8Yb`ZAeYgpUbBuFVTX{v`WxX2GT#|d;
{r-^p72SH?md-`*<"u[ [RR,^ST,phu2_2z&6|:P2bF+L;nHCpDJ*l(%|__O]kfHWR[u*bAMgj[F9[/[w@ s@8fmc~7=pG^3";_d~z	NZ^p'iHZ2ny' \A1gI:4,\ {~qmKj\bQ31.)^IP+$'eD{9WT}>	~2tOQCJhd&lAf-#s	XST4&"VLsQTM%2lA^X4EL<?
?9/>3&+](AyyB>3a5.N4_<?s)ThXvUMxLw
*`;A8-VHmB,h;Ug
`vL:i[&; .K"*t)m.0w[Tot~`oprNKXod?i>C)2;f`2CD%9k`!MXy u<%1 3	@[PyQUq|PyA(sUeGxNI#FU2`OLi-+Qj =^/1v==AUk=1cp"tkws2?:0wRc3[1@b|2>!9cnVo/I)lN=Y+h7l=qz>TNQDa]m
HJZ-dPt:J>Y30au/oI)?vDz_Ldlgiw4/Kud!2b{q)nAxSFRwbEJea"DttwE3KDj!.]bXp7!:r8R?p|D)n`L$UFva25L,gF]d.0+8e@wU2;45'0^ZJw*g$;`Vb'aaaq\fazNo@Aod(BS(o.KJinN2mLdW0s9f;92;-[a}{gcQ	q.LXR+{U3'!FI>cf9.JF"bui6v*,M^iF_X4[%v3>~;]!;v=k0X/ej4^LX-rmSy59W5X`km][9zAjNe|CEJ$$0+-Jn@)gT1kuH_"tY,!},I'I|Rj\kr?L-Qk<Zg^H)jf?tm5-fvFImL7SHBN(+SW#~,'1}Nk^VjqE].(e$.lm[;iAJq0epv9@XOB5,fF Z0\mgtjTi6!#1Y
e2C|&tI/	N;('4Xt|,<zrzQy6`g$,Ez//AkSzME-u"K?;A?<_!SmWu9uhM^g=lK	FBc]MIy3Ss:|S|qW#T=,pcr)dqz$q>`rAO,ZZu`sfU5R$"
F3w7IgcNL2KC%4}=9}Zp3MVI5h__|kyu#V20$S{LheDNN\k#fww<h,K;o4{pkKh( >DN$*Q-22$9}p0}B0zx(s-N4xGemskat02N8$eil%1QEB@B(UCro/JlX6[oN6H%ZmH[`%to'@g{3`q\v6!U={62$
j2+YxX9@VnxCdy	#l$	CMDd@T.9L<$KcC
=K]#~*bNXkJSl7yXnt,UiJlXW:x%c@8
)H}q
D][".-efB!1]7h?C&/_OFPw8.w_5t7PoS/>}|R{4CW2j,0/7:K(eE$U,bxjdL-Kz>]BU3N5|MvloX{j,wTOt/F#|%CX</%#3:KW>,~TgFN1[[%ti4cQ;L8	KLgQ
7aAP074h,4O`6<%/v,i+ \=^ib8UMg'Sp44`AYIX(M{	/M+!bJTHU$j|9J<-9p9Cs"TMH)	X5 <?hL
bnF."1fk]dw7%6DK
Q[W.[.0,]JSN 6Om1c4,L(.^5a.`ue-g	An-|H[Y6Ac3ZrubqNS}<&Tv.hIRgw[65>+p6RA\Rdt7a!U$KK'-/<[G<X,xu:LOJDIauH@|n49#Nu-+8_N|aIL
bjmV?DE,:Bl{&8w]\41|KLhCMBdt0tokt
60T\P67GOFOQu=QvqrAE71G	1}f[Etcf}3X,eo3l^-PFMlQ).}</c.4'Mu1Rd@6kcYi/S2Cj>>2N|&f>a/UfZfG0@!SMY;N4U\Co|K2EA,w~Gd~mtXhcKZHw]T#<<([FO{iJaA:_+7tD]^mS=z`L}W:'+1)kvYiA	%
llk~ADC),SLm=(?0#p
+:ou
{*gD")bMa7
7\Og=y)IC^F!9xS2~wR@/re).Z33J_M29P)N6r0A)3dE
GhHx$*bk+0&9DU"wLA~J!=Ge>YSCL;AzpW1 .37K.A4]&3X.Nc8Q&xfN)ElFs", 95lh:E;6)}i_K>43W]-t)hA;^T/uL(`n`C#:pVo!hyC`8W:|lWH
`9YIFetgs%dzh[5T2N?d<PcyT?Z,!swnpNi\h+JB*KBnCd_oJ!_;:X8RHH{<&#qy~Z]'PGkc|wC-^9[	sa:ufWt":zf*u=r5Pr8>{I	QI!c/lY4c~)8/-rlR4odp.I3a0!C(GhS+-AI8/11S]2{ [htCNi[fq])?V8evOI4Zz[s(~T(z2n5ns	q&0B""+&pJY17jFzk0%UCsv;#;m:!~?,3@ztCbxZhmcMo	|V@+>WFY%\U]437KLWaj9wX<?+G<SfQ\`;e +gSx'>vDfe9;g~1.&pZf7IY&5{QM'Ah\cNJa}9irvsI
yQ1urS<?FsW!G"[>:}tN&dRgPB8[IYNrCA/p19]ix#'}l))hA'";HCq	mJy3^WHXj9SabV>lVUQt !]4
S]"ugf.&tCz=oy ^vLZ7P#\lDqO[ufDgw!Z?dh$lDBlt5+e~>piNdCFrf_;ZQwC>;cy[NY%Lg[B_j3-6i
KU.QeO
_waqJc>k's?1#^{23uk l}PL,Qgfy'$wY^9IUB/j+OcM/@>|Y?aR &R'\s$Ts]/Qcfxg*696kfe&?qu.T&IYbvM8y~;2`."HR@ZJ^x=2UHN{s!}Fp'!>CXe|tjN?.US,oD$hb~aN'WQ$]S~+:i`us$^SD*9{Fq5z|C~fW],=KB866LYctyb1naRA)K
rU`l3nMm}/)n'!9J_'(u(tT}`-LjqX1ANS[hQV7t A4sope~I,u4kiH%ns\:dYqy>Zo<@gdWv9)<%voY&"aUAa}z%h)lVpMM{F*2.{^>7Cg	VWuK$GS*k_%[LZ:0Y<v}A)@}K"	.NQUu*9oN1sivdX;AEiqHhp=_P1Iq?fTEV|wtJ1fV<?,u%0b08QQd3m/@2d5lASm1gq)U![(lyC9(}SaXCKM*?Ky<S::\cO,mnw%ZV4fw4]&$;TJmSaB_|>/*
A6b2tf=N]=*I@GZNnp?"Q1(c#Lg"GcCm9{x52J\7{AsE*,l+HwzfVc,[EY>^R?6zjlLJ)`B<uzFt~@M$=F2/.}BAKx!_2dy['?@GTks9nP[(g5rmFD7MWvekR&P(<Qvh$@uw/md{,),k'!Fla"&jy\'[&~(f[kvw{bPn1v5?8*1>P~:E[by}u<m%fdi@-{<>Z$lk~&*zXuf'QGz'b|J#>gD;#/>L8\kmXv2k2?$U^hX %Sg@_\e<KC	9--8to##x5O\{	Cx<3SwoAy0PSOKE6N`xKLC'o7"os/nQ-[/[xa#E7E&[$En9[{W-pnt,yu?G	dc~i3"<=:?S	Xm?\Ql'}=@e)4X2qb~qfn[\,n g~UUZY4J)^=|C6[7n?o
^Z)AF9K?o&}+t4^B=L=9pFCe&C|}wNha}Ojd=za0G6j%n r+l7bM5E%)$C>AV:G&1myFh
:+#*UfDNF=ZeV :IHht
wkU+RTG8Rw/85G3xlY
<n!}t%y+vC8YQ0_s4w>}=ml<BvG)Pdp>^TRGa.NF`2lM||VY[n(35rK|I"EI`Q'j<5BuY"-4)G)tRI#V%Ta0`$5kGdsc1eafwQRF=%9
Q+ d2<	^ta=i26Oa:#$3ngN_^JQ;KzbAI)4iJftP!_mqjq l4Q}.M=IxFIVWZB+Qadk,V$T%8b-B`VU8mf,a1kKLGsj'TXy_uaE] "aPUjwQE~_mbW9nO\[n#r] k(lfkj~B WT^;5P}lI30iELM$+d]pj hX\g*wL,hoe3KAW	!n5j/='/WV/Q3	KsJNM0/ol6'f,Eh8R\:='FUmf"k3M
r0i|&<"=	W>sA6qRzh{@bQ\Eg5'/q~($d<'Cfe$i;\GcFK)7(nMkxSW&TZ3uZ36m_CZr;X4a\p0z_BQIFS7zKX
2U(%}a7oTf
ygB-h#*v!3N
z'V;I`4D;.ygBo"JJin;"
n6\lm&&0~ ql L}h"j{\Y=ao'/ v_|37IPtJK.mOS\D;FrJ.P":b=Yn0aA,OaZ_|Imx&r\61Yrx&Fc7%Fl4tQv\"GZ,$%0`L%FM;`(I+j!L.?]`ae5Dz8DvR~!R/D6C~Acd@KR<hy/%a2OFn<>')[r?/9^<2c(odWd3Ukx]O
$KmIoz{*u(O	2`Z\f1tbS`0fofXd)Sg}{JrBmAA]10jD%;bJANP:g$-+=moz#PZNLEL%(CjLt$f=auZH(LsK[s-	~Z5WcB)L=F)ka}m@`	'dT	=c"
^pA.G'IJhd)Vo3J.T^}dSn_Gpe%]Iw1gv&;MAkA	DUL(_cq$UmA#k^=OgCfo,q8D3N,_]~TzkMZc!{#-v!R'I\0J4;=9A9d8c*#zeHA q$_R2b0Umu?z,7Kv+7Gs`!"#!RxjSgEK(}<iq:QKO%V7]!VRqe2Z=>	Egawv+CP}$Xug'jBEDtE3u6Hhf{Ahkv@!r2 (Ym(Zdda'SZyD|7\+K8
%R'AVRPR>P
1Rgy?e?AH%W@NVLMG`9S-Kr.*k>'=10{to{g;>y(>P:yvggH6\0Y#-j=*WXMIOo0Q*i?AVR= TPXl*[GZ(*Z!n4Y*r~5Vp<LWnr;FV0]g,|o.Vj%(=FG2{h#NzMOT;Ln(4){
_*+;lmd_YVe4f\).]]"Rnf<+2Ht|MlTs=Q)9'l=%Fn	6u>@^xs(4R3#rJ".3)7#".BkHno=tMG~@(@evdVB@tTKz1|bRB}[#e&qsL@zv^tI~?T=l]4xsyZP#%p"d@BT:`lt _3(f-DR`9n{Ft8PB]=J=p!LYKTW%.!
\HQ1PF/)<7lK'{{H,3$!2p$g%`c$K{=Lxw+8Uwsw%^Y0p4JOZ+Y\GAi\II@u&=WWr7||N0	0Et|A!e@[HSCA,33_ZO!%Zv"%YN*|py)s}h,9Z)J'c_Uw*+Yr*!<m.phW	Gz&MjI*jsW')D[j\wmF?,@1$wsS`e~hP]-.]fq=0~s?Pr*W<DP;2|SM?s=N&hG&j`TMN=PO)F#m.^!{&0>90P;#h{l2}}BW:1"XYya2EfW|tv!`E/'"([$|ARhi"V?,tV#4=fujTDb)Kmb9?v31|0z{bDCwWwhH#cK-r/p9b]QR )^N+it*D@P`@jLF)~!0Bgb	d!{6 O7;y@"1C]MMqP3^!c`_P:\:2*xBq_mIFZ[ZyD,WX0C-&bTdcup(I=W>9`#__kDojN#w+q>{7,=ief>tArmzC[l:~GBL7ijjF[	l+h-PrnGC\(9GKj1Oqf[>JuUp:EHNh>FAcu.YDcqf~OsDN19dc2m}F~G
)urftr-D1NU-GfdWOt{X`/>J"'ePH$~/Ts-]*A[m`"&8GT!xd]7	M:GfjJ~?aoZB7zvh!I:ob`\HCd*l2`9t|8GU)\ysDVp&3!Q`Q<0n>wq%JwE&Wg>@zk1pA
>-T6}U]cxKn?(cbwt]Y&qY->O+WJWnlK^L$Ky%rk,p{/Z3Gok^rbPb7`v#fhtrQf*{ZV5xISTwtn*@
@W(E;w8t)@$6{IQb_vI3qm2ACj?:oK=xVkGiQQXs@gfFU_2H<^M0716wT|+nxk^ pm!-R+AEn-]f<+CzA2v(SRl0Q,7A2Q6"t%?-qh|.|E?.WYk
N]zMJ&w@um{uc6+ sX<aASE,Kf}JL9QWX#P!(fL\"[ 'W(wGzxPHGMp;'I2>x1Qk!2ga+*	dflfru>4?3A8o	[E7;5J"z	XTViy\+jn#4CV{6h_!}r)T/Z'^4&
v=hvR%Yfq*3&<\Xp=gr/^f=geR~&:xLu*/<(dp?%=_s20KyW1`6[p!'8=MF\SG%aGi8=ug[/FGI7"x-hyjDV0uH~|
*n
S`u%OE}},>]fAJO*Is0[B!P<OS^[~55UjwZ=?>y@q"Bj>XsE|to0=k4[MJ/jiEd=gI~=@l[kv,pq,.TO3Tw9s,XA=#s_o3|'-4	+qd[
! !Vu/?O}VyG9x0*`skWyK;-^9Z_3!5Jq_/V=_CHE<mmj4[	&1$A%")>[3m51FW%p4>0g?&R622wO`do&NIIK{PK>|5]{?0`&:y4&DP;@#x})f)d|^iAFCFxt4k]	|IROJM
%;\Vbdpt`'I=D_	,A`<p4!HqK9^jj"|x.-)"L8Sy+$F8Rg*MnGj/<(Zy2
&]R-8O{fRp1I$n>u0:'[sl+Lkz|_ pMVoa>A~/2hR%(~36+|Xt`z;k'B_WfD5ljh\-$$~~Q2]?,0{;#BVL\4g`;uRG^\w$>8c[A#mY\G:;>1]g"_8Ol4OEkh$uPeaOTyY&~ah;jn)roNW1hkQssc%\BB(	N]6L	Nds8,!,@v)VqhxO;P^POUA.F0>d&5DSLfFmLA5kXU
9_5-U}l=[e*J9"$%[(+rJ4W$SxKix&?~q[wH&Q8vuP"+
wN=021:MEJ&D7#*Kvprq>33 hpJ(-91#^oeNWfQ[[gw%iob7RM:44bDjGuIkZ^xq:;j,|e?xM|V32Swx#Dha',*I2v4j+Q*y;x{COzB>1Ns4C>$@S,50Z}'P}
Y'8q2gwxMpypGO^-c,/l1XJ[x/Od~aJrYHE;kdi CKTNW^e/l~[Abz`SMv&	1IRR)KANsPU?pBA\@a"pSRK
DG:2G1Tr|849J[A/}%{~A(Tu0 
a/Dh 7Ec'KR5}c[)1Bz{	Fq<6h,Tab
$Be4%'5S$xVP\jt%&Xb(>jF9_$ZmW>!ruElBkM.Cw'5+4I
L0QEaXD_R(ibi63#/.J=&pI9ODtx?}PU&2n!Y2^-U$Js+NsoCqWsQtR#Zxd9ahO|;$.Y0/$d]'&/DZpR9)t
2DBf-FH*Vj\`d[fCp}oLzKZ@XZ+@v)]=}XNMo)tDbxKqd{evUfNGy-(fu${R>aa~=m&x]Z#"!
@.Km%&B,*QuQyYVFD.kv	Rbc@:$#<7~6oP9|"mbjklmA\nPW#)n1exaiu!)vA|JU	:$^1P9/>_KV*5?:spTEh	GxI;2x{'%LL[cZ{Fqzy8B%;8J6CB#gJD6BmK9R?MJkUWLIdS?`kW[15[#)i	X+wF2gkr9b9PE;+c[8)W>c3*iy3cA$&hFov0WkE;:PgvC0KO*
41VfYqEP2*!	LI$mgCEV:6Bd-hdSANW7$s7%~9M|2#mxp|#;5a>1VA%&,Aj(U71F
a@e?sN`cUM2@:`Les`1qt*}c|(A|"Ka<H@<-vxqc%Dvp*Q3gmQ5hG'&id90\Ma65*1#;[/_#:{_59FHhRP vObWJ,VayvFZs%$*>Enm.?Fv?W+Uv4J~6iHj~a<k{$*! k"=>[M04t(8s{^~9$^lys$fW'"H=/d_U]L;iTDZ9?Ic2
F2}2X13f[=zZf)B|7Q%RoFZT@\K  A,$,Db*?Fu8 2vq#|)K(A$Di..Rg:>Dg_7^}^Yk8QOFAjv:W+J.ShM*T(<3/Y-4<
!u$pFHNJQ0>#U6 HzsAgN]lYGz:RWp'RSh#=HSDa:XxePD4xo/#w@+/'<~
sw5!N12ZGlbgnX^F<IOj,)RC{om+y"e}^/NYFV=l1EO`[lj^]OG:fd0DUW>$_lJ^
mqwx>uDg"jt,YM^|zL]~6w|yU	q X\?40oHgzu35o'"|A+&
bzV15eQM!Q6XiMQ&rmH#2'T ]+JHWZ35'}r3aQ<fLO=v5(P{'lr9Qom9-1,O|`"9pM?:}5a!A|j# s.z0TH^|'Pwp.w1?s	i)Zz<hh@]cjG[-xt>Vq8-6DBiv$bc6gzY-<xU:S1Z2c|d])vCnUo_Yt!HZY-t'*#dgJ5)z]cn|}2M:dc H!wkNP0oLnu4LUv=A,'|3o1yx^5C5KXfG
OdtSl6S_$LM)JN-ihAkK4Kw. *m`NdES/5!+4(Y]T]^|:#-Pb@vt^kS&|5Pqra|3T9~A HP%oQpK \sOxR
+5fmY.@K)="LWJK80{n|rD-jzi=/L$e2vszqQ&]1! OH%oELionBTsnna/"t;!dy5Y[yVZtj}][Xi,8WCuIv=RD@&tAo#hU|zu\-z*7p7r#]3L42`+?!(K|6\/n@wF_/:1*5t(lxh) 	f<6n}$)0HD&'?Qn
\Qd*1H|;h^Y(t\A-u#q^iU@B`.;dX~[_$WF00)Ns|.
XElT'[/mU~b)eWqqQV=_TLg'!]h8g{="V7vTD5
Mp;z O .&3
<F:u"7.Mt4rQ %nz@jiwP&\^DrxWNkR^:w '8W7|6jyzSaNhT;sU?~eg$JN$FmyIUbcxiGBq1Q9d9zV[z9l
1yj&0RuhgPXHjXkF
u=N<n"prw:JofNSCvZcU}-^#fN~CK=5kv|	l6SezeT[nAJ@+u"\QS,D*zue|Uby_Rm:=2c?o3:KJ?+%.k[qJs[(A0u?>n>
'Z?bV{Qcv&%/<Nroj%\]dZ}2BaJp\*@1)2g\R[pCv~mB<*HgqM{Je'q8$Nv.x}BsQCH2d{Ofcj=gq7Ig2vrC+hIpyk0#iW@Z<2pu32coI\gammNF/E''&n\(|*=_'q
|tJk7;WJHfr_i'$nt]EA"{q^MU$eiYa/16N{Ok{jy/1e1d]e-4
i`L)IX1Gl&BW:FAAK]=`2){`qn/ubz|0TZ<<&!mKjI\^]c6h3`uz1P'uh$)=onv55v%p![Wr3f&\[{=^f
rR}H9%IEfzfA!;ZS[kS?kG'E9%RU}(;CTCBc:]dY>7jUI^V"id%bTHAp(v,53o55`;k|NDw#J<h*BVsBcFeX'Lb94#[rJ?m8$cG2A#;)njiXub*-Y$s#]XWlK/k_2w0}=PV,jm!<nRs&BS M8y?t-2#CP36xp'&n$qc%~vc@Ud0fg^yOEZ!vB>8:*DE:I_Vu4F	
+#[m1NaAL6.:qvAv
qs;efP6	^/h=r)7yQ`{{7
Y.\'K<XTxysN8To@]pVG__29~6xK6zm:S %$ay?tN[Gl$Ff4t-4sjmw5dIne2WD.Hr{s]vH$?9srP2rCW$g!9#%t8M<Ce(y&-qVQ$b\gF1zZm4jF;AC(T\A:+(H'{b(A<B|lemcwGc5mV&Ik ,\>)-$5sVn'r&72ene?u7X'>veI|56P@x!`}Cjfw'Q2H8DgVd<aKY~eKbl\!]?v>H
Nn[:2%vo6_bTHI-puwdsOQDiZGSZmr4I>o;wWD##e& eEl-k@7>Z/5K5Myj9+Ek&$lPsQ
,q[},X$:W-)br.^<eA.8@D5?aI4Yor+}R8[YlfxxDkp.3y)|/r'B*qRi%'A4hq,J}\C:zXC5zq7-8I'#3{Bob_CNK/DJ\HngR^IYS;Pru,7,HSv`-t68VVrgqG_477RIBOYe(tl)>nofGWypa#g6K?"`b7V`exa"`={Lp10>[88Ht`IIGco{?:,BACa}MLq	=|B'Lh}xt}'P9hV$}a*D^{/NAw?iJ.':X&z4|oW0mZ42ou!rwFTl1!"]jz$#pRpMbe!kQ*GI-dBoe#o-Rf\3fq%N&eO\l
jS1[!	j+>=Cd)x1hjZ-7t3PGe`40^c/# %
rP:Cgs*;>3:a*CU2sJ:rP0e%"tvETn3-3Sr;.u}W:8R0:]O)]Tc(T:+_~Y#UL/"8`
~5mZ']{Ae>GHH[3/^]m8'#AiBP[<vFm7iT$,2ibr%PN 8e0Z!6QRl>.5;]kkQ1tgKA
Ed)Pa[{u:uC2M)k(vOhv[+_@8QZWLtu)-;fm(nciY6\]j{,&>`&sT/r=}-#|Q=5"f`&9&6{=AXp4<6&IfN{G12tD9rhT4h@$[jwch}6rlMM`R8rFa!eHnNWCiGcfg`h-MWf_
+TJX5<{.GvqF@)m X,{%Nfvt5"IkK;. 
\)'(z	O6MB:9WhH'=p7}r>aB?C'Zjk{)]h/mspKSdiW$##i.	uufE2JO!0^%C<^*=S%x;j:mrrArRpFCHyoU3$%Tq$@B	McdCF:EqUCuuW!|E]"Sd)5'IKa+ja%M8bc]rvBkXEFEW(Dfl8o7K}Q5"zUzRp)yA^"k$.. k;jW<dfNiP7#2Jj"v.WMvs:S{vSGrk)];uFx%'**lz$a(j8E5YavVw<ESZLhrlMc=OTh@w< VYv%;QYao_B	SE2=r\) l	W+;+F>77,\8"9kpQ76w.:jnns	B?_(lyc4G/$/@bNni)Sw6z~)KEVnp eo10t<=Xcvc8*<W
*-a0nAv&ME?;8][e1U79f^k&m-?vr=jDmV7C>?a(;w:~{=m?E&mQf{5X8!F.Ad;C	};g:xh01u^FM3Z0f}t9jih:R[G\=?|v0I6v+&HJR?b&UW4ow7kd/%R\o%<;[a3h3s&tXV7.[X7)pn0%;cjj%=kf#	4Wj!
.TpT'O79T&**Eyl&@H4
/y- *p=iO'I(CqI'Ghh)P+.r&(wkfTALgJ6>]v&~~)W"r}?kC*aXN4}D((SBPht%_|5<UBy%T4EQ;bQC%[2|
_S>Ie\q|.7$]?plc}A4i^k6@oaLHB^1G-GATd(rLZn'n%lLJN32vCOk+(%a.KUV
sFsv-pQJ`m)L%bPJyK{Z~}Dw;FErdB|^~xNIUYi]J{QJ(H[:}P\9@ZllRs'C,&&5d5u&=_/1<^cR6:dViKAL";;wA"JwVs`ht2z=m{@F8^Nx	LEBNf6~6}8btb%)"0RD??
Q,zE>^6PR_s/'qAxpj\7QMXh^
uQWe6oKD?RZi"eZ]k$D)UlH-D&PWc.DR0Mmm"`j	o;n|vIcHytBjni)PQwUN^2'R=_#'zds
C*I}lq8]%zQ$QFP\+y;H[0*8==O7A
3WZ0p;:"T:mWf/:<T@@P\Cd!sh\O3<RR^"EW|ApUER-a	<3Hk_E8No2N6KcV`pnWxl8_ A/
J%>Ik<Z)f+
&\=w4[2ZeOLfS'-=Mun[B{I08B&.b6
SvGyDmtq9:fjqw7t`5]4z]byjoq+t;Kz@gF>GM{xmZam{Cy\{Z*u}FETOhcJTD#>lp[WA='w@\@_F'"Pr=%QWmyx	Qb]M_pdJ*H*<}2^Joz2~x8,*,b,&4Bfk,R7}k=avqU8$0}kl\;oDJU3`>!'Z{|k__DqR|hQG6PPiNskwX?o>N@2194:Aa8L"h9Q/[P}fiv@Xu$!}|k43E_-tfA%CA:RLpz.
[B95tmn|\SKd,}.X2g9[u1l3x6q!>07+uQE"E1	#hN1~	s#vM5-=<ny!56_@3H'LAi&6F7-sfLS!i}e$
/IoTW8syC0}_`O=S3}[.(Tdkdnals+krKR]c%Uf /ZV4[KHEmmh~YGosvelPUw;,R_xh@?@!WIn-3zsb@0f}*'AGCO5Ik{K!p=:<^0?]8[Qzd:rK*d%N/P%I_:>K]qk78arfm!Q >$gdF,?_^74+_	m:.=r	o4_JOprKmVw&A:|e5!1z9Ea^vKMc{V1BlxJzM2?K8W ]f$|YEV1#A3yOyJxZsgQG3xCwX{+7rool@DUYga:}psP:(GBo!FVu{p>r137q)b]
uo+x\1)G6vxulG{!j`da:/f|P^!1S$<T;8Y
$WO*|R}=0klpaaA93}e3D=l3|/C<v{*f]yyRY$y#0Q_[}S&xQcR )h}\\Pn ^wZ)G$l >WuSk>p	yg/<9.75mWtYv"E[(B(G]o4E%v|,Fpbsr4q%<CIRc'|3787A 3ZH8I/By|}j"'?V#NB4(AkuS86Z{mNv]ds?X4	ir.pJ6DllHqVEp]8Dh*9WvGEl?`G$cf!oJCHr{G.x0,hcv|hi+dS*lq(]|9hhmkP[=a$A[zG*pnvU,8s'T.+~[|S4VI5RoI[dTSFT+"_A[cOWYDS#'g-Ds{7
MYAoc/x2</3KEl*8)]=;`-	:8K;HN^|'
JU*x8;>?n? I#iJ"XAn`#bb
XA1tQ>^L(<e;KAx	|I"0Qc%7}'>"NU*}TOiPpvLv2Ey2!t$&
#:aH*/fo-=<'lUDog$5A7*Sq ;M+Rc^'>wq#HrWe~BGB3.yi4#.kRpYkbL>J/bJ)(Ta@pki(I[oE*kCF
VXKdld:J`*`diA@C@BOiX5x>*x}yj=T.Ffy,\QzR3tJT!peWRkoj*DTc(Z_.<\,iALOG[la-EMW-JbXO.=>Ai=Ek=ZyjnCPY9_QbR%bvr#\9FUevYCnaI{ Wbm|
i*r$ve5tgAPuA"v$q[JIF)>.QXy:JGU@Uyv2l-r@vD'z3b-56}S0kr3qx7y`bK:
5{or:mvzq/SPC(y I'jm]=_6`5ji` 8"S<n,0@WLq{:5Or1Hz2~0Ao";q7'PMO^Fjhg(8/"#fnU^N),?$gUi[cizR	%KtgE;hN9"4L5&yoarf!21u&6 wsV(_O~G%lc'|U_~'YU	NP.7@|tx?6\SwBe,3oIY,UFK*\x5Cz!XF be-u$G|3o:>4sk@SOqU|vx_P"%.Txojz[E1yMja2d~wVW$8gqk0+#HcjEh|@''n{=R2C?;.sC$F;k$T9szh?(W&-!* gzD3j/3_Ks*q~(|z;/ud^I5XynQ.2CtdEl#r-j5Ao8x}=3!?i@hSo*x+Wb {U%L>d.9GP0#"&@~'D *6'8e
gV:>& \#*kF:Q|'^s!nVCS3(J?)-?u`s<W7_~]Jh<DUK2oS{"QJ"\Rmv+}Ud
G^ywxV[3drZ?>J0teD}Up4k5Wwv'\Ajd%Z Z1`\;9/B
&&0Ih^4oh<e22
. g99}HkzhKG/F_27.Kr?W4HVwweg[a_Pe_Nl.y>m9d4}PXX*&mS5v&$,V^fx";"~oOvAD{dog5?_}%&Iydrg`UI^O.m&e<gA|Ed2_V%Z-L2X[TGg,Q7l\j:BT\i6E!p2.1!"Q:/y.'p!	WYaS;"1xTF]y"k1h0mp
L75er{`-B@yg#[~/sg,X;:	R.|TNYdzhW'1k?oG/]Mdnhq?iHfW8McreC2yUYPey;uIuH`QJ:@qnZDFmi-nJ]XI>G{mh-y-f1]n`At]+np!4oyc{`+)?O["xI&c'Dbxs=<.OYH:=C&-~3lH5+]jx~-U?94nkqHo6y ;5HcQw/STvT( bsV[3/0>~Uf"\F mHTim'WbWV{UAMp3qE a>~Uhd0dyiHfSh8hd?
/1{j(r\Pj.pj6Yo)k,3PA6H)4g7>=HWG'9D\jNxN4#q"!suv[C"(]1) yZI,#P,g|1[yonJ{6yu4L|9blDutw@jAY*e`9cr~1G}j^{%W*Qr/Y)m+-	PAe9ccdFEY4~,SFPBgv<%Q&?rPk\O8TAx;<"_ilrm2rCT:Ak60G	E]Gn;/`2cv>j_GGg5NJY*l=("aO>?>RU3CN`>WFG+q_\mKw;M{'_vA~;tjbd:h:r#1xXdE\(&!uRU45=ZP:'Y;FvjssKg:O|PXOa"gtnlXW+F|,/PT'mj@hzqXJY$h5ok~,!vLa^@*R~l]$Dtu/!lYCqG]~T=<P]0SF{CTfgheS37WOsc7Bj AKKr+\l! o1:*V7j~%Iz'>(0wn8$7gtSXl<KA
@RbaF7$R
*>+}5=+R.R=2^ b=$G0Wk)%fDnkGaGz;-_LE!+5tY0`'%A<|,&"hXaS?U[tyj&~yw<dh@/
{)G]P[Iv#aSr>C}'>{&(L]L:xU8XqU$8b1{yW,l"LNVPZ^!hT:-v[~!RYAS]i//@^4xzPfV4uZSU~U,79O]"luv4%	FevDFtjT\-.	Tv">vt#Oh0P@p[llz4`?7# Ivfc6Ao+`rx"{
cu+!1#[T[&4c>5@<g	9x#Nd^z@7kWQK1v:I7_B)Vw5'NW
WMc'3>T`h%?=ZVnegN+GBvDiEHRcA-pTcZ<\QQz#=4q*a8|z
^#3q\5Z&+.nCd(!)#0oL'=@_g/;1c7s-Cek'@%3KW_e</b9,vP5AEcqUbEir/:cZtd/v^82)	*.W!!9ai#^""W}11VXZSsHX]Ya:X9!-rCFMI#xgm`SrO8M	'k.p(B?\PA!\>( ["{497C+8d*Y) mgk]7ArN%/RV8jt1kIp.B1dC1GvYSp6`
X8Kt'T{B=vp{89^66KzNhDX>GI-^pLRYVqik'N`tQ':=4r{Z	x,m{Zz^'.!<.b|a$LbyEkLC?A:9?jbHj`N$|/BSC/UgfHRp^BXshBY/o48g)pu ZdQ`|$x21b+ >p&
rt:Eu"F1[E%*+"qt`eW(e$ajj+^&y|a?DU8@z&7Zguj +U~g&=+;h[24(wE\tE*y)Rj[jc0(oME1R4p)vAj	^ZTfyQd&3k&B0cy@7ZOBX!lJg<X6OjOI&7?6NWJa	JUko@'M q0;>,Z\x#
7qP>yqV9K ?}H`|3,XZR@#0:y'rfhu#1^w5t#o4e47A(0o8?ugOvunR+"h+iSuts[K3r;KAd!\Ie],pxr8OtS9oqL"h0B$m(x2cb)'+Ppdz<1#K8-S/#\WTAs|kP?RHKmJC[SXKE~V!9No?'Z^bqu8"L8FD8cvck=,8>%C=Y-G7nRMvb&v5D#9HhBJrk4Is"eP*PALhQ0I#E>Tutr3"hI{=RJ&xF!Smp^2ovWeK|Xcc^jJrg?c.m@: 77rT};l{j-O:O!c>a
u<{{/B)<V.b%Is^vg1>^,|=(uBiFk"\yL@66i$P\;R#t
Fw?Tbn`5$(DdXP;=	-h4Lg;JokI~rT>P3Re6"1{+Io9O\fdfHz|tbq&)maTT~gI;z&|AN7aaXVj"MDS*P8u4M".SBi&N?d2hc)|Pqif->(YlponVh|osP9z4uui}yY Q'uRsr557zT @d%PmBq(|dIA<w-E
awh%E*b2pa<4i
!KM-GT9|xfuuE{.W7`=urSjA5UEcvO5}o'93VX	;4BIa-:5Z@?StP8%1^){S>r6a83lT_{[Zl^$;Z$>e1S}9#_i3~B ?vMP}Cl)|x6:A6u)Hntq{0VA4[kJ}2tSOmwqC.\0YVF^1WuCfPDDhILt^\3 QWt2j+@DMI0PhKD>?B.7Q0ycWX>na)hZObdy_-~#//vgZ2EC#)m*4oexT~xwb;V{7+aT Y7K^z7yE+K/Gt\6PPxBDQd	{0K,28|_Qm;yFeJhE%21	#p#&jAL/6fTXs&gDZ'72P.jc P"W{5Zs(4 I&{,?@T^h4nn6rsa~_8$j$a\LZG=N5L")<B|rSy'y8wu
|=!yomU;nK6h4#EtIppB,JbuV@fa;E7}j0nsb#(7AGt:>3`C}.RD#M,{{X\t9O4Q=e:Mgp|:h1<LLlI4| O~G!=w$G-9OK0`U@9IB|\+\dwzl0NP\ZfP<f9xr#>D"h&&>ixj&E"tv``c!5vG*znN0E].?Pd_u2}D/eL^Wn<X"<wdaC?%uJ2udpa=[j`*Wbusy0[~gj>sd,f
/G&*rYKl*yQ|85R(;Qd3@vIkmz`AyLgEOpRTa^:}fRe7_v1k)>f8!=~*&E]rfB-!oeH|E;t7jrm,@wJt36jW08kx	7G|KA~S$fC	f	x";5X4[F[y.&yBhaDS{OPx{n(C["0?Yj;F5msR!lA|u5D'EK9*TKa>RXb<LEQ%iv;iZ?!>!mm>o2.Yp#v@USFwp+Iirc	.FM?#^X#jVW5>tZ:Wq3NHz<6!WgoA5G`0OW)@MN%ZZZv]^x'G|%n+C&l0K#KAcH@jAc=1g)zn]u)IG`l/$%uz?Y!ho@L:%&'E+dI+I$\PTfBXm+EV=8v8,Ce:K%seu+r':)nO7#[Im`n"{.
-&o4DsKDTWm}nLr(z<FQ&nT)apRu}!cEdoU[7(t	5I)M=GkmfHpDvt	cnAH&q#G(9z0d76V*AB/P%F0<7[~%NGa)
S6+*YPk|;kF&DF&Xf@_$yLzm%V1;'pnHNw)tt &JX> @coB&~Ct {md6*j$R%!hy@8F({udn@b_gad7&x.s_`lkJSBpwn$!kS@4@$W+=Or]F)
Ktz|*3b ihSu76BSR	%P<	zRvmJZ_mkKe;RCC"hZ+,3#Vq&~)D&$H|CH-ZR|F^@no?B&e?#A`6FP4A"|WRm5HQg+0x;w*JHRvzx(Q[`Tvko1vR|%C6[HDvRES92?I	?3Ocm|kU\5Nt,r$
CcADy
+Ij?FOg0Lq&m%{mPwG1Rpgw.bJ| =#Z_Ir"xX&j]b&)Bj.m*4zJGPyaj*>$czk!'W5ma?=h:$(#lLHJM&k@}[z%G58^pH|Tt%87/iQ#_5JAkXDkkkZr*<[lt\|SYun{\ 1]~t:N
m?>`T7/)6sa9+|'z0w`){7kA9WOvwP@,NY!@CVJ!#ILDSw|PVf<.24X}(3Q`~J^FTA1JF+Gp@T~}vGXC/&z4	,rA7a*xbo'0}bzk	"eWp>F9+ow@KO5G'QAk1F0-W]|Ocr;k+,{FSM>!i/Zy{1u5VO@h"DoN~IIn/>Cj{3f>#3jlG}cqH4ji<B6~|)4tM=Mu5|/*zIlEGp0 Is'Di29z23yT$o*g!~u@|'"	R%<I2`lgP'~pj[>{}*R9<`/U&~gt:
}[$+"`Wk=U7R( :o J 7],>rr+-#>5B`7r-;sX 0Y2*.l#&&}rjL[%gn'pR\$OGcez1,]S'gJ\S|MpL)N7#H
}"UQcJ_^y--'9PkL={#^0M_o^9X{2]Pn _?9S[dC9`8G <OZ_mZ;I:EkqQell=Fq2IWq?|{U q4aT=Dt-LPH=LrJtk7j-0b~>UOBD]>?Lp3`lP`j(!Qqz>PSpP D2^Y!E?;0C9UxVN?x.?X<Ob-P}?"%G>HOp$kcvi3wXNok
G'-itsRde3o
52LHH&f3R9>pZky)64FjSq7F ]T0d^J5yi\l0z"~Wc`Z"\Tm&7_M0<G_Vw]JJM`<(n7Y|-R,dIoX7qD5%<t`vE^],l!g{%6Zd"X~A9`{}v( -&iz-##nXF}YLSSRO5djO+I1frZ[;he&O>XJDYy9|+"`p^92;?~^[W&
#R&k{LLnnQ`wr]PT\m+sZAXoPhobDKI!qHJk7r)fn"j,HG7U_^N-w~DexHHaB1,,k(iq& &[:6psT767gYN
@}\jxpc|+<L
1gS94ibBI~+9K9-RuGoN-oD 3Nrt0CqdMV lm+DUdv\:OLEjTDkl:o6(b0nMu 0H$UsX"'vM3+#p&]q%~"RK#d6~&=JZg1W^oMc)nE9gBb|ydEw<U;gWhYr'X-y\X{GC(%q1XK{E8}Pv3$fRu1`8YP!Tqyb2Y..32{fieT> utJX
$/[pdQqZ&Xx7DIGzMJDPj}@Pm gS
JrDhjO9gYBda"YEtX{p)H7>W?{u$]?.c/y(Pm=edaKwoF"=f=lJNP:M$B?{@a9|~zhqY&;n^vS_~yvC92K7P~k993/FohZp,?A?zo&8H{.;W:]yj4G':3Sa}4ODPm[)zRDGkur)AJ@xT3g?cWfVV@r9Y\ND`<O^{Psj3fo
n;{Ld&/*Mi%0ko*Ru`!E"@:M49	 EmKcT;ZOF2GJ/aad_"SmvjFG@.H	@d.@UnyH$m/=b6YzMO<Vu(4hW,{^BcJ?b`
fuW`j1\D,ECsLH;&`lnG_CaW7gH!?c&P-/'|&-))tbLR(SrH/n6Zx;4K#lX]$IFs!Kh<FQz-*N~^@K489$E\<HF<D+_ijo?vn.L3;HF2]FiK"TJ	X7eJzh@k(#$cHiQR#%5x2wj\hQ)gmM1WHl$d
RTkaNGGc9[Lv#>#w]g#)L8\'Dv45P8p5hy5hl9T |#<sj)M3lK|[0vSp3lY9)-+= |Bu>;8Py{4Sdi#m~/1x,(ss),\smy6]
/uW*{'to!
K?B	x,#;#ml;y*SGf'q^tMER_>k~Oo@M!7(l!^;|GxMU7E9{rE@QA8$^QB?zUn`xNw~5]WMM{s	h%'HKyVJ&['T|MFUCrGdIqgK_^9~1szaF|[#=*E{`JFfu$'}UMyW|:!+!c>SV<0z+[O?
I0he}"A1NLY'GBWG1_J,!0NiI'M:,AQXx`{9E}o I3tyC\6a'i2N]}(
/Bx&F|^\s>vc|Gi$t4\Y="{l0$6PmFSCIMy7hOCxS'|`K5]Fg'JGOfamVAbcD#I|\.%	plt{;fiQ{_JQ[eg)%a+z"jKwC/RqC?(A6Rr=K&0&k2>Jo:% gQu58	gl,RFX)kE<Trh'	LISc$L:e 5_2!Pj>ww7H~,D>A8XJU!k41Sx~f}p3<PX* zmI$;^M+iXFi5/syU|eWUV|=DQ|[kY%WI0BLJ<9}FURr+pQQ*V#tA^SFa/JeXlwQ0nH_r4@B) @^V79exw V$z=p	aE\X%qNLa<SszO{mp1K=q~1<nTXunZ&	R?=gCmf^G)$M IMk[c<--T/Ee]<X{P'ZxYEL&6>q`	m,--{cp^:`(>DD2G&}10nQ[I,_VXdS[bu\*0WA1aa]*i=<Tn#t$F3|`Gn+q^h&;Hu$OPaz-rw}5@)*@_=IoDJj4H%Cu wTBf)Vzo@;TOD*D|}%`&w+6#vVtU)/>I GNsd1	5TlX{F/z,|xW	YEkKU{@'P=;X]D7UZxU	dC"<jeBAD3~thzzl!Hj1<2%p<K=i_.CI6x#s.`l*DBEFPbiPf+S_c&iPSjnpbq&2l,[h\3}xF?MQET?OAj4b-ce.7yI"a>N?t4P4$Q>hm}xY}]n ?Uf<eH@qPM?X8Um0nemRVK6 gKJPPnPZhv4vn	gS*;61{6hIh@pJ[U>-K<q9v!;Dne$Z	$$_%7uTt+BP6VMvK5_!eeh)w8T,;AL$tJKdzjvERa1$o|I><vT^R(G@DWS/vfDn$xtZJ{rO,>B_KLfm bS4J]X7
X]mEzwNdo83[9X>!I),%fP>%E7\cZ<goGSH
IGVe,NY! 8"5((p?pJ[PI!=o+B=%gK G~%(G>iL!16=v3<C4p[U*#HtT#<*K>ou`g+!li;d+	t)Qni? hCq(KkP_^Q{{&YbkR{"[wVmK_[[@":4F+{5rb(i40OuaLdP<JR1'JX&kG87|Wau?]IbKKpVt,j<u}Y+cn:prbGGw0.^VDc^L%l){>#')=:kH,hb&hH<$,'9%,S"Lc]b5#P3n\!d?Ir\C{Vmax0eIS~"?:+\.;+nh)
@%Gc-N9] ZEf*1LfotI}^"|EhBw_kIX%EcP"W~\<ey--z,recu
j7"*^Z.9""fxk-'Z|a?h2EAF+rm*Q=(Yuul.8b5NEhf}1mtO|j[P`Th8/|?GmS6!][	y]>+m4	>3K"dak.Sto=k"/. wjLzFx@exm
]vW0<m\.</`@l)L60Ov&p)m!tvk9W&X@8B`>r!=,Eb,=tMQ*45bN!s(n$x)2zk<@ &=G'2d0ftjbLUY_*d1D{EpmL+CAE3`(R"9OM>1whH0`H.Y]Y(MI,X3R-1Ry<J>s$'E`^NzQ!t)3
Vj91wHx~nmlq5BcWz3FW8l=9Qj| &iWkk8YgFQYT=#ae&ea`!
8FU2AI/r%A@7}3aoV?L,~d/s&][/4IDHGMRY7bUr`'\MfUt6&I	Yo'B6/UBXVO'Sqw6`{QpYZJ)lp8:w)*TRw1Jt'8[, GfQ69(Wfp(qIl(WgytyVS7;$W -?=ho;aQ?jItd5HjRc`WS($/[
O^G~EGIhXw!P\OeXY4piI[:V}VOBtO)J7ufFxFyTTL'S'
>y:%QPng-#x =||^3d".p1qyxs o=4!&9"c~*>5q<M	5r"<a|[Wab^wq\v9S.i?m%
J@'SFmyRz0y?rh-U:lU3 a<fc?L]UBP7`ff`D^E,vZ99m]pC,{D
mbHe:=2nWdJreP[g!]: ^8;8&kVBr}x_=p1]zKt;g,]";Ae>zUN7pDSyW`%128]?:iE{m\y"E1ptq,L
LZY3@kwAZZ)v{}O3
&pN#0T)=*0R='ZJ-$Es3,0y$[`k4~ doRy\a=5-qV`A(<W6}lf|@#(,d0,0*f]{kpsyV2A*Av>ntQE-9!gZ] Fd">_b&s|)b`ey$^ Ds_R=u#Sj{WT(#2z9Y^1q@u,stgt<gexNL2}v
WTJ@]Qy%;WKN>}Ck:R:5qQ	1WHTQ]_z@DI)o'HMW]xFz26we7N8|sDTRhI>YS!Hb8i;_g={5>Dq6	V	<!5~7'q3zriHRj"ER3;4y{mJ%vN7$L]RT?mx'QL0Jw_O<,%"'F=ruC%<87(ZS)dh.,}SZ~WD.HH|f"3Z;-&qsdv*Ut2|9Xo7@mL42F=VU*<cS"FClMCoxm2t$Wc0Z};dDECn6WMf_R'hm;xrEnHYOATWTrc!T{:%yW9+Pq$S
zw)N`6tc~[{R6>{;zNH=oD|0zV:L2]zh\#ZKa=>:RB;#V2i^Z~(gD8JP~Yg-`MQ
<n#RNAT(x"qKR&~wA6/Bv??dus>l|BwQ*kwc:h4sE6!Efs. $CcyrR,0Cf?j@kY)1&-W+sH-$b;~F9ROrz-w+V%J27*Dmq`WrM
w0h;=fl^OJflzGO nLe[z5SC.L%g> tvEPYU)fG!<r,p:	9
`2
__`_ 7N*^Tt~*Q2>J)cqk.Q@i'b"#[FtUY+.JG2x-d>8S?tQ_tC#s$`p %ygV
"&W([Rq,\4oi)#;nOUa\l0nGx:IinF6BdU,(9pZ'RS`/V0R`2Q0XSwCq3|?AXh;Aijbjfx6Xlhd[inuC3%EICz216da8Sm5GAT#p}[g>)&	?,p@{jN,/! It^
L<X8%In@lJ&uh&#kt+QN{KG"C4vt9{9hR.QF]6aI*eHJzL(R0bD|b(R5"f]i (FJFy&5(Y.;0@nW\6HDt}5Sh;Uipf38'm=!8SS8E},*XG^>R(O-DQo4u@	kA^4	0fosIN^{]0I\hI+
ynX'/HCpUS"5M3S&&!H,"=ZN,=eObx5	OL}6ykkV[zz$Ai-#	c(W%nl=WOiB?Xb9dfP30ZZ6	QxTR|K~x,!l<O{_WV^Fxx9R
xiDOxgge%HDp6K{dn(P\]E/}io%='fw,f\BJIVZMleG5U;T'P$nH{L\pqsDhhv~PGx%f\&@k
}Z+qawgVE2*l_AbPh
(HcK(1-=>z%BV0132:5VkrMoJIOLl]/y0k']Bv,0ZQ)$wQ_Imh!j3#=
MALg./QX%IRqVP#9f>]W(@v;#r)6{n0P`Z:byz*k1MTYx3G<9\!cdR`sF@Fos<:iTiFPv-\Pbu3mI347Tcnu0*<IvZa^S`6?*gc[nXb7X_G4E0Ddtb-wbDOb\3V#z[-+~XK>SAUjfGvXgvf_]KV$o	@kYR)9.]769L{4;'TM/IG6".jpr,>-KAORQ9C&`IL[/sh[:OC)\x;#6VfL5`e:xxlhBPd7yj'g5lYL+sPY%=|3jZ-=#0?Ws\>k-eE,)q>eqFc7$2s+}5L&_[yfB/qm;WuR\~loyCM0M AA{|tpZ<VI*GqV}kC#e,Mu
&.Ba,=:
`leDWj#;R^`[xQ2:!]29{uA`yY^2vbx	I6RTz)dq~_$1EIt+)uaKz@S$CI{B.`gIKL0$v84]AwWf/OG&hIiPmsc@,#T8v[Ui,R0D! ra\OsII (4Ou
R+tg4'^3hRs\5|{|9vW~|C5:va7*p|Lj7NT&*3I]\{:q	dJS&)Z<ggRze (IM	q@
d%j<DmYV'R\_VCNB	O$I6H~\XA0R+6AGLp/bcGU3l?g:V.=Q[9)D^?Q\T+T
\[Jd*MLJJew)X^vkR*]o,}(4~b.pzwt>tbL<K?s-3N	/*t(j.,0["<Wd*|%[J)]l6;n)bLDLP(`rkU6HSi;%7|Ux<138gkUDqj2NTDax~I#MuPE+8k!-~DaLG4l[S7ZMa6'dhv_rt*>N_~gpw)
W]Kn*CD%m\jY8M<~0HbMQ8i*@9?13{ j>eLXV=H6GY
^dirk'-H!9uC}mrvd)s%>wcpwxQcU(_L7"`(	)]ULswl*i5.W)n' WWy7!+H=wzY%*6Lo5[QO~#"Y$O!HE5
&[XI.&VtvS{T4q<mipuMe@?/_izp0UPPIS|jZK>qL2)HQnUB.w(Qm*AX5CK7Ga@t[xT:Bkv\K`fYJp~]\jO,0NM004Sk`_kO4NaR^pX@N\K;YjlwVNa\<vOGN?a,Sy(aUO,?q[3uqwxQyMbSnC N(L-97<B=9 d:e70d$[~W,{e:^Hh|DHUU+_e_|ik>N5BSJh?anS@i)VAH*_r^|Z|T$zwx]]Gce>/}H&PaR&+D\F~v	C!CVNJqIN+(uLMm7\QeRaC&9YQH.vLK+L2As']v22;$:93d<.^@#(S~5&g-Xl>M.ORJ(|kV?KkF3;(}SGeV/{oN<HJ{({`brN_j%0rbXMcZ#+ak(b=VY8<L{<X7,?[AyP\X>MVt
+@6~l|N\v-Ccfu4D$:-"g~JFh>eA!mJx{s2`IO23Xsy(<#x&4}Y<&T+lhj^y_]V2&MK@hj`RX2U%{=ZM0+AbCdIno6yLij[@Cnhm>pE	jQj%x %$<
^T-2MgqdS}|IS.-Ro@ET[4,OAj@P	r`2^N0E\Q{I?*q,Unl`E@
\(n)b43lmZ3/FZ*7Ny2\[nw6rq/4,A)LCOAA>Bo1qQ@3h/85syMtH%}[Lg4d;g-2 |N%H^Gn)R:GR>SfEt\$Ho]kuN-95CYPA+oba=E(J"wE-+%] 23'i{~`^{)cU]=X!z>z!g{b#u!EfvextS,6vC2o fR!N's^yJ$`!.pu:K>z(a#e3%wPAZ]=B F6Kcrx?Yx$+v N*.1U=_Q9,@nrY"IF7*F/?:JPT%{b$b%JGe$ 3Y#_![!m(<;?	V!18kAl&%OnwA#[	OZzP	c3PCceVEsy~#MAljQM*gW#cB	OQ~pDji}3Ob5E ;'JdPK|D}orrRb'G<5u^
)~j}Mj_r?"[dFHljA2s|aD&RRE<	TR7NIC;IoYOmNF1u0O)DLO\n:0,zwlAeh'a@m*dEe`3mF"J2g-6S<'3xj8tuq+f|7YjqTr~8kDFemmo(AN5	@pf
";B\+Jz`{Hm ~%K4n#>*wyb9xK</q>xBTpF-`{q"(XmF7!Y^H2cG8jzOKY%C%{/POtMVL?M]o\$^@u#h!U	NxH}"|&rKq`"*{)jOg!"CO|%fS#/CiC~N=TJjm6sY_KKe)f-_aV<*q<9jBJJym`v#6hutT`e=\I,FB?Wu2#\Q-Jw/s)[$`TM@C4*h1-vxGJDNs&6~]|\{+Gii$t0'^,E0.aFajAC#u_=m\eSWezmGJ#|>!PNf5#y16~PRv#fiG/IhF0NpCu}sUjN~:?J>\Y6H#DnNWRtj~H6eglwpGKuKyTF4Ua,~RN$;s)7:C+Ac0xvz<KKEPOsI@`|H6-F`5**)y>@3b^_0"[\"}(![`kJJPl{[[5_ydT3-^l&C[p^pq:(p)mp0Ti+kH,HO;}'3cVOB:w#5&fiQVg|1J%Kv_bZfZ5xAKf!a$	3L7YVK&_'#"OIq8;p_L7(Js@T>|e'M5a[@\5m{IZ%h"{wZ9EQm!/rO &F0j<C45"|A/{%=XA'Q6Qu5 "82
y
8i;Z$|q-nlhd~3%5iyq2U ;[*-'.fP|g.)u:0+7EB4PRp&A=qCEb&=6Ce*w4|43DRFN\Nl,A:\V=pm+4LDeD\d6W0>Q6Lqh_Fk_[C@\jre!_]a]?s'U|R fw1h^5xlD:<OgS=';1m+jjWx":}huk]j$td1}[=|('7te&mE X$ys*D`V]LKG{psUN@1Cqc
1K I$7RWEQxHA?l$&zW3._$:YYP(v~x		Y$LeTnDfCF\. 3B]`Ifl$tc,FyD3$ip[?Hv5l]7pW+E!JvMWBoM|VT?mAtM{
HTZ\zFIR*w"aG0q"\{GkBfbe)nJ9cr@<;AnTMM^@a(,oti	(p/T;G4Ga#^=(>,Pu'RmWDMwYru00M8SmH]\z-7\K8`]JU+dnH@'W2gYlc_0F?5SK1yJUB}$SQ
cm"+i0X="h^StR=XV))?+NBLW?b.=hTl1WDhF"EnV]K8@m`Hyi}8:T/+n"X,X:<\(Muw15z21#0qZ[A{Ybaw{&"=mg;6\)nP(+&YC'|K.,|ScFya9X}/"l_j$UlN>9R$\]:xIv9xKX'D.ge?t>xetz*|XxKAl0>6w6cB%3a
8MFmL>v5D0aNsNnuBfNN(`/J`rx%2H0@RUeH(h<2'9m5#L!%:PTz)PwB<XRn5)KTmuq={O.p:$F[k=!yHcE^2e,~)-<	hd1jJGkcJ5__H*6%{SLigy^Crc8E|WoI	4?^B!+_}*o-Txc oLlGps^/B26sUVDV^s\{xHJL"RJ3Z1*nj5vct__T_gMYMrm{bD$\$l*0CZ
7cj9?H+/A/\tV	9mb4O|\h](xh,;Um*7^@4Ex4SBu1jJQLimM<B``C48^ElUk)
-6v'|
#i#` %+,_xzZ\>;%`	j*hyn3h;g/5kvsQD(%zE2R)jA{|P$%V"@U_\;@tM	W?9{RV)`fw6c#{V"Pc Pm4lDs\jxl.EF-a+RpZfQHAmmNWIvI'W<_hb|j$);Lj}uw{]Jwji5g>[Nny>%0'8l:7NYS'FZ<-7bDiEP2}kJ93'[{K}|	%K|ehO`BnkD@@VC<j,0k9wd@fR~vaavR6*z+`X2CKzd46RV:pY>Ga$65k9t	\~uE4kE+]KrDe2DIJ\0yEU%~E_!(@-Z:@:fdbN7PAhyjD]-Ur|h^jIpgO#DP_lf*rm?1r?fMmn p7t^9sMmVWYu[@#V+z1>i_Ud$8Y\aRTM0BaTbGDHb,20MF{e97Lp&+jl$pI})^!|k|)9)>jH;'5J]it5M"^6;#3"2E"Hng|jkLh5n'V+lG<sHpzdazE:t9 }rrnQFYH4OB2Y0IOhj;QQGcgrgQZTym"i*;FHQi $txbwforj9R5UOF^^-EOzgsM{^)Z.@V;+<UW%1`:f3}*p{#+9n>
<,>(z4q%BL5<3;4dx b1Wz9t0i-#so'KI7`mL!uDdvPFK/"ma8w(/,$5zG4iuR
nSKC1g$_GY9cdDkIr:TLh@d'lPC#GH1FGSE},^$o8~C9+X^ulKL2x4YviDz`'sS"25EKYc{HQ8lzoSVv7}L Ax#qokdo@goFtxvhS$;W<z[,z1X}1/.hw*bA#Z5	c02:w$9T\-y;fs/j^]D,v&nn,Kt}J	]t}v1Q &Fdppl'HYTWCdW\9mf|.q^1"5k=R-Y:*Z|l</v@VV3I\P/Ng?1x
|9#^
D@+o-bT2Sz#39I5xlN:GwfXTu/;2k
t7|DsS;}>4}_t@1<?,2^HWn!=lF4oC~G|PHjIL:RaGF{J(}$
xSXUd;OSV#|E;WkUZG;D=ak	7926umey3~L~`QgI:66|C@X7P4'CRUfeycW4d'iYdmSs;:hAWN=(/}I/5Dp,$\;VV	\.eyU1	&A`p/cc:,mh2y[j@#4psn;E~Bq[4[sDuNk"YPP4Me]WS!8pT&
F9?/ L(.Z,]fk>,Ov8h0=>1"{F5+/;PZ]<(a=po:I5F_8vD@J3)w]S-"C(|w{d7K,C"Yy	gYBRpkYty$o!Hl<meImo0lm{&QXa$/YpZ
{$Ne9fUc@X)}}}Hd`jyh#,	qM3MA1a"2qB6N(~/Vk.`t!LM5>Bib:Qbcnxn?6UiP3EOHu;?ViZe,^\+Z/#7v1~<R8(ro~Q8Pi '+#Y)it5i'-IBtb/hvkZ`[}kI'j2.Ju@te<6Vp1C3m0wUg*k8+q:9woeiVy4_f374b~U!FiyAoGjGkf!2B:*J^"/IS<LUtr`ypl*3Sw^47y):xR+h"U*vN3<8kUD2\52!;]o>y/4u/RkK{Q\9,\]Nv7'@`MTYg!{#,\>-v^*'1m,@	GjKBz
Pd&Oizlm9$NeOz&/)hdW*kfAs2[37GjCALACaNPFrD|}>fF,iNH<`r;6L7II>ihtIn\Sr
s{-b{i"#
N<{zj=0!Ai]x9D
8i(
nyjSwq|E[t.0<BX6CO'e&,V];`jbDKn{t0+\<G'isx$^HH0?3gf	Q3Tdq#O=p-[XyxZogYr\CL?2/w/Y1;TM'6k+e&*wG1d=0>}8J1I>$|(V4LT(OJg#vo
sZG`>
^ef~#MYcn@XpD08C.5f=-as|(e
C*_Np=<"1G+wP\#*#3~xLo0DZ.A]8ai@V_U9ryfr#,*XJ)KLMpKB8OhlgKR&R.<0FLb|)H75O<o,AdoH`R>;q	EFHojyuP&E&W/;&~Qe:CErLU}jBxEq0`@$sK$KAMj
|kqqA{DhSA9A7d47~x?m_bz~dy%D	GEEu2?(Gj1SEJf|8i%`Z,F1`|
VV[D%N:>"3:d~3pXtMV8/*c@/"FO@C)5yvkNC_tD8t7e3$Q	:Opyg(yZ$O
OO;GS j2)G^+p[p&C1!A$8o7cw+[$~E=&,
6W2\TS+,"\KBxR?e4<4*~#RtlK) }H$%]@q&1i	\H|ZyEj8IO8`C58F97)5VzY2H{]z9H8dq!.TzeAwXcQ DF93~H?uc!K/[~[16+Ym&0i. kksP'1VxOIP_l^c8l~#`TxN[&wW6{uI1(PsqM&=rw{F)J"c)Uqz	XvL"=)
p.a_??XM,N~9WJ<>\*b=|Msd*m'cy6s\.nA%Y38?sZvUd$WXdV.aafg'I!"p1B]+x9z)6+.;YJ+H`J5fO2{j!p%xDB^f'9W|ae	Z.8j.W>4)&m*--unk$0y$zWi)N5!Zs\/*28&)ywuG6]"ak[*_8p>bL3>p$L}}}|9"taEP+WKTR2&/Z9
E0I/Rv6OmB0L
,hV?js04z)[IpmXW_!o);axVa$Zn"me56G6izd{1j}YP0OvSZiivB'YTa-NFF	Hain!;$B};<T975RW&38)|bm3e2+p>X+-XxCA_b6QC~%3R}).1u/vpT/g"",s
jJB\pU@tEpAx 5D0jsdQ|	WhPW6ubzO0RUNP2Be!GlvW%`*K0k~RxgV+6.3R<Ava%zvNVX0
^Wg<Nz@u9)]5@Hw}imI:)x_j^oi60	8Z1'E-M.%|hRvJ?T49b7E#v87),G_M#O%v^2(Yh,m}KJRZR@?K2<Z?6/,;4"o7zwVJs<Y593(6j5;
~7SmjGWSat]hy:~Kxh_+zUV@3zN>->vUEg2b({Sd9z/j-7$]GEqw$}g@#>	+{<65ta<"a-29"k{w9QU;DsG	ZC&;4x#e*X1
ORj5?efi=R-%F#!*jUeD$
zUwNim'nZ!;VNv(Jw=9xomgO8Es[@xqQw&
]87OR%z^R0zSm[`=4"W+D]BCLf'!Q
g%1?3V>AKT"ki3~qY37%eF=	lUJm8[jdxg"[XQrQ\chmm,2*KkP3{P`4d[Z-zP
9CWT$P
>xh&p:3vrb*4f2@Yr_ZL?;:% 5}Cw"n'wOy@(:C!8=cJrpC^_
SV%knVe>I0\-isjBWK3+_kyF?i> hhQ) 	"A%YJ*	--2f/X*Jv$HreBEzF={=,8	2zwwg?6yj$0)z-<6b{G \rcim,bDR-@DXljuB'`m1t->n[k;7>jt<&t]F|rae@!ChL,>+S(k"Ul]h!./{4@/"|PfB<|OU\^4hyK%1-RYMLSra`ke%
O.GlGj'7wuAsq^+bix~
HjfY
OITB."(;3N=]d9+1ND"	Lb

Q{4sbb*A.j;G0a[kI)DiwiVo$#%\n2;h
c$}`AO|QCnPR{w)f6^z[Ir8tW/xIh0ucnF3]%#rc\Fd XX=t2k9Dl;*5T%.`EjQ%L1'b{OfxpvXUOQdiSR@+Zv/'YX5P7W)gW0Txm-p26rwPuNgit=(;r^yl`b`~e#e3Ma)iPIivLUr_EuXxLdf+#KPyGT$eqY1iEpcm`ygG{$g;0)Pvo`.vK}Lsir;(05gR	W=iI~Sr"k,xGIhp|?!UU[iys*Ge}HD:z7kboRV"5K"7S{gMzKb)2UZk~(Hy\8mc
sFh@J4=q74!_}S`RzT95a|N/%RNNK/E220GIL6qOF-\*%+SEN5s0gR7"jo.dhO0fBu1<"Ae@BMYzykpY:;/"z=Wgh'M4Wvujw%mZ	(\rDFU7aa`m:;f&=Pf."EZczK6*f8dV|(8~@>EWO'OKz89S?w\IZ)W}]d|p>nfr7V>9
w/oL8wY9qJS!ydx5OvI,A/ATKj!QXqRq@h:78c`:j\nS;uKg,{ZP[X`pv*Z |2VXMpa{0.;Ej_NO}TLy1iu?sK+fB84*`IvvW?&7wzaR^f["J^-n4o$K@_qn&I49o8LJ[5n,tS.)6)5CeEV?{y5Hu3FW6"q>l0TfCgm.{23 K6K()CfP;p>L08>ql"L{!BGyRxmA'VtPFb>aHF^&SQoaTK)K.@	\y3e,op<lx%)rCD[]o4Hy4g0s5dm?8.a^:V6Y0Ek8JF!uVds8
"`deDY~|!hI"bUTL$hK/x^00E">'A}F
 SD{Plo"zT=%Zol?'Fy9\fBUwN(	G{
~cR)wB9NM4K8"rU>FJBdqlrr4=-6m: BGQRUV@PF^#d]M<fz$;5Et7|Q3u\Q~qt}rfQm5xCOy.u.fZKu`Zy0&K{L]oW#	!xp%9	f70@>i895ucyJ$U_Iw=J2Qqo|V~o=/#Q631Qk|d3bMdMODU>G'9@=4jX8=N%cS.gHp/vzjP5`FGW\xDmx|Cn2hN'+s-mR1 smkG9T9AiGP
CH%#(=t@hNw	Cu,LDdgeBWYiY[4{	"61h!j%?Hw6{H9LG=[45/>1j?/I4Ra$<,nN2Oq1J7rzJV3S63!b}4
9s\Dt@L1x&U]kE8r2OI'4nO+-aSac`wMAq?FdBlkk?;9m(TB";@7852&qSPyOC#2l#VbvtG]+ yFyMI+HHag!3&BJ/MgJx8T8O"qx"&{F*}>sD
),~
[dG]>l%fpSj@-}uQ?3J&7{`vz;hea.@CKz\95r~4*nD}.hv|gv5,p}	#ly'hHij?'.(-7?!MkE1~I]Lo+TY+a*$2Cn0e"DivYwJaUna8vpsDL45mB(/LGbl6#>C`$qW=7OJ<}c9g)_7D*lth~vyxN$tkm3z`Vm$Dzyg0"/!*m+dBTtyz&Co(sj~bl~Q:
%'sGr&v>]	
cAerMk'F{x&]C,6@YD+z@/]^y;BWm`1N"WZ{WWxYS-mHFy*MPvU|?g{^[	(F64X;E6y`St=-_t>O{z'(>r~[</qeU52Uz1p/aiZ-Qp(O_+&7a9%s%%uDR^x0dCZEQdg6-p[m>v`QM%<uY_KB"@&]MDMO70"}k8yVRu%aH3*!N!?DkUO+ 
!FjxE8,cBU<0.2MV>[?1ws3/V
rO|Z5WB&B[R?jYwp b5]yZ|nLRKd`	haZK{qvNv~4eBiNe8\NUC6 89@$d_H(~Qonx|hEcI2"Yr! wXoc&|RMiq{h`R0>K24iWTLV_zG=gK8EcIj+	{AVe"9IuUlRDrIKg~z6W/gN)T2=`'tE-O:3//Q|y7h'ih%)^5g%msPBQZ$M`OB_CH'un4l9Ygtfifx8hZEF6JM?	8vZ;`{!9%EK2Pq$_$3Eh?AkSPFea_F^lXBhZ]Z1J}o; 7:z, 8J-/I=)vF"]`7MqMTM2'q@q46py!,CArDPxy1v}f]_$)9fUkPW[%l7&(m0qcRMHA-Pzn`k x;(r9yI U]\&}Q#Fv+ENkAqJ1}J|[aw@I,|AYe*JOttPCmy&8FxU8Wl4)-W
j+a'#X{Ny<E4Nq?YPz9
o.Ns>=b~[+?9p^GaQD_X@=l$d>{x=Q>UvH?Sw%<7t]^L'HK![dE}u=W"UD?ujkA}-ak/;\ge}%O5o(Jk> x,EOTkS)HM/}AB#]zM_vlzHZ:@{7Vs<rH!2Y`@j@
"O=/Ac,pT-XHIitch;"@E
Uy}<4ugcv`7 )^T_8G0%wB4S6v,y,th.{RG	U0btbEp7>:`6b|b/O${9dSb|+W#NwZML],Q-H=v uP	wr]B6Ue?#FE~S0^)J;\%UN't4'^3i,HX6^S{XY'SIY>['FGG:z	x7N!$#S4%yfFw:uFy^"#'1})Cxa4!_Yf
2tvH1\s{]lOg*([ ),S}`yt3*_JBmD}+sOjPsR
V f[@;lgMHlC.xl|?z([rT^aa8U,C)MCBE",iVF	7Gp~&D]yn9	rWCwjm%On<[9yTR~Ef\%';gtc-fkzl_/ysf1@?#^4gCP5OE:4Rt\!og(B'.VkCf#7r8{5gox| vXa!doBRVo}-/>`6Na/"2dbTGo9/v'x"W}_(l8.wafaJz{{BimJOAosj,
R'#5E|%
2pc}U>D+7X#l*zD@u,E*R("kviTM<+'>4>_OMT;WeG$qN
tG7l! `9j^+;!oo}h(+X IUjcngD@<nzRi+Cb,SCG-bICx#FRExqo6vU>(/Y}E.[@
fKwCm3R	<{a}BRrUgsV.gk@E( PCagjq08k&>%cOxE~S(za!C*O$6 *z>$'{#T^Hk".#skf X0L^xHRrL8<0x4k2P$tNf"]uh9+Zjb}}ra6\5_deP!};Dnz'W>Nc`N_ADqJuH&HT#r?MS\H%"a8>Te[UA5I]L=DAQdD[0W2ayrWF9iAL;.&yo+9mt1# R-4WT`w>)sk	^9 }6BV	cX"$
dh`h~#5%-0(ThbIt'8\qtQSzB0Z57HK}S~rFw*z\r5E#&i4r_vGC-0!Ptqz:mmRJc3sBK{`:#.wG"q{`2'M.#PbjjxoUsLP{xE>'s|EVR(v|P	,Db(~'8	2Q2H H>DfN99PbBXXkL7{Z{S-{zP#.+i<]Dtx3Jzb(Oc{_NW|PU?6eonK.F8F"y|y_,<|"`YT|sIm|KJ;9 j]:pPsZa$'I
	;k'u(z[XdW:1!U)Tm<+N;7&;!"E.$=pc<+>i~1ni-#jKEoXcZIzd2H4d5GY4Er2M

FrA1B.ph@4, p;?:lndfGg_c$)khgo95+8r(dd$L*/CzCkXJZ'EHCs/G6qCuPu#HG6IGch~uU@n+uE-Pw~Qth\O[[sw:U[$G=w3u.	*?FlE*Ag3MX[Ky+G^k!	aB 9	s_S&N,0AI//Ahs-- 5tlQH{av.&uq_89N^^M]<$jO|G=pWOsq'nn&VGYD#E]Tw1>5BFTuW*R]4+0h<|\3J0q(~?>tZi;ukKIpQekf@sn=<P]r}KY+G	UO9/eu?P9

_IF19%}63|^:lfQ!tcKU!M.w`%g>+]4oFoi:AVx	~h"'^7U).e&;v0t_!s?S2 Hm:kJ% j9fF7ENMp@Nm'/.o(OM![s3Ru|qG1eFD~#48oA6{P'0tU2R&]ZTkgZk@W@{^]uW-hi{?%G^^pT7sqi,5h+s+>IK]&,l {6b{JfFjy9Z`iB^M6H)Twq
KW &[++Xt_!fQt#+It(PrlzMqv>Ax1a&3609q9I%OH;{a"WlgG+_zC;>b-dNr#-f2s<eIZj"=\:*/([YQ a";Lgcy3A[8A8;Rf<)A;LfO1*`JVA`}OqfD&9:FQUY?u|0
0e8>NB":x{UN'qf9'>j>RK\1p<9rXar2:.%|G	)P$Q!@9Ei@@$U&e&?In:8`2,j(.b&$![J	>%P)iTDK	2),MNW7RE7<#Hgxn|Fk@$q5lRtSe&yGj:)p].S#./x0@|KmZ[Kwfg8_z'7X==;S?'[Y8/.ZXki7+gJVF[,\$_+nM[
Uxml}h;x_'w_"1reaScy[l{v,DENx,M=+p
|3mIYMP8_s(smVmT	crN,fs[z|yL^yhrL~FMLCj^O~oDlCJ7%fEhY[PI^4MVl`H7JC7HwhGY
h;b0c/C^
L%hL!pM"5+m#=OE!6Pkvk~sD5LnNnj)iQqeu,e/f:&!~9ojeVtMuGV 7
qJ:P'X&!Hl)#Y]'<ebX,xvkSa<p&2Oj! 7I;
5h(]*6LCyM;C`d1|)N5#wH)T
&%Kzz QmI]2@aS^$!}@s(I'&rQk{Rq2xaoIw LQ:;s_e3$58;^B0#:xdORN	 =bet+rM D/bqe "?,,1c6S^f%Ihy7I<Qxwj'$`O$(`rmHJ|'*=NhGFr8rM2k\eTc_P i3n9crytp*__dm[70:9	4FJ\[KhCJqT_t3Um-qX]Cum*-zMiPywKje92Q,:HU	_S9R>hItaA_#h	J2#Seo'8PqF{WmD3.&FvC,eHNyt{6j!<Mq~LXQ`S;P6{HrSn`,_fJ_6%>E5/%su=D8AzAs9TS5z)&bV;>}x^\j+L'@ZvE9U2]) s%ii}REM9;8o9)dU+MqDE?)AMfOUrGeuy%9EU|8[If!!G@q"X.\4,EVRV,y	3p-`iDC>CWz[K"	M'T&ib|Z_>`hZ(CXvtK<Q3qVBv	Nd%./Nv.gE04I@p$Q{R^$p%^E[a&-;<?!wsg,6njm&G!oIg{RSbE+Ch$QVfBM0vD$NkQCAeT[#)\@q({U'&NWN):mhXw,h\M)R,ZqRm=i}- )G6.FXD~<$qY$4$4qofBVA|Uyxt3&AJ@b=7L2%clbrDXyo'|#LOY!LA+2gD?w",gd1')%Z'pPHd4XH?HC"BaZ'Ff:z*.tw.0rUZ]6H9\*bS?ta Z>/ y!k@UYJb\L$}oWt,NDnkpq{w9"]0[icib)3M_gU`Nf>=~MK|Q{]n9td=6a*]&-hQOf{r4voEz{g|@7igN48+sM":]cXXBGU`a8<5.AcC&F53gZMV g\ycMj0^t:o7PcT.p!R	d"}?XX_~hU:T425b#Pu_{sdkp/z(q^w!k6T
astnBSlP_C6N_]|Q8X5FWPy1]sA-s(!B`>27n"G'mXJ70W`w
C{#c=/6V5]Z]w2~N6WP8y.G+!
l,|zMzAlUi9cG$s@wg3VNlTC_R,[KICd!(^\|W	DH@=8x`>Ca]GhK0#9M6d)95:kv2A{S/zOtc6O~k:yJNW&{%Ku_Ue+xysv	~o{LlVl\. _FbZ1xaxVfB^BPtVNWI$tXpti,3FAg5:*X[G!|_Y}th~jX!h
pu(M`/>Z,1Nqtb9EW'ya&Ql%zZlH_V`xuG-tgZ@ Y989I3u:nJ@_6<mjzD01|;sUo`
k!S,{IZ}fQXS<p_zk")vxPt"u^(4^1"1uP*K 6/c}.y<OA2%ykw`M%*@]F"UG)fd?V<-#wK
A[h36rdxX$L7Wa>^thC<.	aEuD-8S[d<p}]F	qNyM>D_xr-E3I	a39Yhz[f'S?zxV]	k[S/u$H([,'Tg!KT)m2Okvr&pcNd1RZU(\sIDA_sHp~'fB;=E,H|+hC9RxsvBf304_Pns1'd_h[4=e}Ue1-2E9ODYY@>/l~&k;De)Vu2i;v-r}^v06:8pc;rdAib>c-0L>aHcy#(- X4t`t3g=-O}H;xzzb"FfoC._G}J'#DPoxk;Kt-/M:Fw2E|E3yYKijrp6m8pjv%so`DW,0u\O%xX.9EO[ChFAg\jiZBu2x4#qILv?uvVak"ZBy%fE]q:{G93[1/vF|5`)R9T*et(z.Tg^exb&UQd*s))1Pn&yNC_x	Du&OS*4.WH0L}<2&aGp
?|hg&W$BoYUB	8|;:ZyN=6)CT82L{E6Ckt\pR"I[KHpHNHADFrbMMhKc:7Plv1ZkyA$6>>H}`Szf;%EOoG+)wA,}mwA5GUi._EQqv7/!GAGKje{
R[.)@)<\,;WRK@`w$CZPt Oy,Z
X4y6("ge2+6PT3a4qEQT4c>`N@(Qh>O_b.eG[F.@Zo?b(`_](bO!7`3iLr7ikRB|iK`L15qO*1|,W	Xya8Ig!9'Gw/(8f?vKU	#>}L5J-*PLYZ(iF+u'&G[.8T1%:^n(E-cPXW	vAq2AD^0RDb{*p:~$Qw)G+@5Sa#	efN<}r~\]({L.#]+$@O,^rcooz!B6TNT=R	ZCY"\lKnm^T5s5Q2*NBD[&(VcgC&\*5g[kS\RPuUmZy8jM=w/9JfWM.Q#b3kUXT4n1	4tv|eP,EOm$gU/(L4I^2,bcf*1;6`{AU_lP45P`*)F):m@fk=l5:&4rZ:NTog;~l|.y36c,x6Rt{EdIwm6"f2~Ijmw,F	RB1ZM$^=wzaKH-
5w6v=ntTXcIf<6Z %2U7M62
2_i,0ib2El7)mGkt=`.sDg{[q<t`uhC)MT8YA	7
T!6s)o\V~!,;Jm9%
9LoD6O<:.'I.o$|Q~_|^p7*mXwg.4eWKcj#E!n0{nA
u=gaPKmbm4wU}6]"Dqss%k#&~tv=LCt(B?WwZ{0'E'z023g[;z6vV-, <_j``$]Y1=QPNewu`%,#X[AlX&Xy4;\'+#\k(]@T6EU}T
3	^x{!3#LK`Hn;+Y^7S|uub
LVx-yFC`!J+8$)%=v5{z3diq3qF9J-h}#	1'wWD8&%ab]BcOKrj!b9,D44`u!tZD92,=-U<@Gc^b"TJgD7'%BU'K3]y)bnLy6M}\go*T>M5k%3WTC?GJFOa>c!eU@D$[4M6$0uuJtqUL">y	Ir .+N9utw:VvT[M9m7& %a_YgY$O $@wslz{s}nDmnDjN=]R-~G0feO\WNc;!}'e0>LR(S/)[Kqi\U92/L~Hf/Puf_8#6|D/p?ADf-n)z;UsfUtZhSIHIqTKm5H_`t6K'jYg?go5hd{#VV%:D^r{k^I+<4U&[zSOIl)52nAnL>prC{)9%)JMetyKa
76Js-f,ty2aHB4xA,!V
dz$r8Z{= ZxbMwG{XNH
jj%Y8S<TM|+\oi%oW<%d2Q0syAXjsTvYp|ufA'%
2zDJy`){/o=KJ2:KyQVHNKo9v}J&oEVOdXGG$k[}{BNm"*"7?e]	MQt6Jk,%Oi&+Tl6ikn"XL8	-87e~	qM	~BD`Uj_ze-Hzw&?>(EV'9N4oI]u)<,rB,%uvVs$L&"dY
Yd*t0sES?LK1*g|v@c\p*j&b~N:e9zSOHn.1;lpC[i:]NF2fv6+K+jfq8{li}?7b )sUzUy$NNCc_}H;aZTGh"aPk*,b~&% EBSkP]Gjzd7pMD/3W7$m7<2Dev+ibP5odh6jQ,Z[>	{!iQ6z9WS)C&4iIZ;yMy"XXQ?j<oy5]"/f/?eBK%`SGOotsUf6kc`ib>`5/fg /C1)$#m-9(v5j&Vp;+ky?z%+Hm$nRe5S{^}WKp~)>Y
c,/a/QO%(lIdc<0Q}huLgG|"i'#2UrkS&>^O@&s{i!xdrZ6vuMt\f]&)QrxtAt"]g!FXENI5^p}t;-UP'@t*U[D1CAlTY&\eZyHs9HpRDlnQ_"WC-S!dEXtUY(1{!E7:hIl[FGTA|8I`|~)Ts\1OSg[2$b%#oThQC1+X0)rxY|:ivn,tt0!T*j&vdDI;UNY5<j+:5g@c@\g(3Z_@VG<[/5-Ji:sVO=ifsB:r
NQ rA0rQ#`-N*;WZYVusGDGNK@$@W"/YL,>Tl%wKzAm6HbfP?#tf>tj]=%WyKK3|cJjWy]p?g'874tVD=IDmA[ODZItCDRTm\Cgf b1l_H:3(F(AWGso4B5XPmS2 UgV),AGM@8K\1IvvvupPtYR}tVoW)Wd}qqS4}8tw/ c9	Tf#&Ihtq+Xs-LN:.#g\b19\V]6|q,^p=-%xW	;(aPr'0E:e{mL?1?7!bt@Kr'pDv}/.(y4qI	hHl/>XOk:nCw*ulb6E;5j9nn=HZv2mj@AmCf2,xHa
|n'fa,t`YxgyrACci,s{B^#nV{6/&BD7sB]][jkL*tbhlOp:20y)~iooc]Af~7Eg6Ew	6)5J
p!H;=8w29*}<AFyB'$\{v,.6AvqLoOT'4vDhP~7l)zrcuwlMYO5l?QRD8y-kZIOGy{p?#bX3?2WE0J)g m7=_8-)6_z|g[Y9^@pLTbJ`uhdC04*q_8$lK88{BkU"-K(}|h~q	SjjTcS-BT)MEoki!.TG|,#u*7v&Lua-hs&46Q.tKU}9E@d#iaf<ED05*i54(5cgxLV|d~1wuT4Z.s$:T03@svbH|G!0Q|rq$?k]^j4wwTVNl]\"e~FBj'U}Ka35VE2_c^uKRwPL($Z<:?d7NM{w^c^{s?@+}M&GA{ooR;7Sy{Z"f
rOn	|]2Z[^ LZ)q{pN_HBVmM<x3;n,("W;dv(D<9Uf\0m.D)){:(dliwJV9,^9GL=X=eS6}3&,v'Ax\dNI_38'nat)ULV8H.Tq{!($8hduSMATxDJ4T%%17uc^"AM rtC3ozOwy\r+6K<h,oN9s e{cUoLa)>y}vS@s#5JlnnGGa,&T8VPZXfHLG%p`G=X	zh<T`<tAL~w[mR/O#xix27l-];[zA,Sn[[H~gk9WXvk.je(-V+~<I*?*qdi)lVFn*L@tvYcTzQO)&{L{),Zz~*u(\%U		<cDzUkW.lb0G,.M{	yocj"E\5(KGgUFt_8fg)r)AYgp1#c	;p/8:u8bW>ox9xybJ1WrB0KjdKt..9^i"t53'IqA\z:wK-} q_vsaVVseGQ*J/S\\ll
%i?(ei^sFyK62.n`~1H]#^o!KehdW%Q;Kz!"=R2f9>G=+$QRN%P
)-r|8Aao0a-zPg$G3!XwK EutLtbUg-J1>w3Yor*ZY_C	= AxK3|Rz<L]XN}({RP[N>R:#S	Aou=b4UM#wDe#_5l@jnF8|@7tAWg>surO5J\!cFB4lH06)/w?8#40b3I2*|}z9HLpY w.h
K~_V[{t~"gsF xeE{i2S*)7i!at/U=KN/f?{<[E%0wGw.Cfp+N=>*(	+t<)>9c9fEr|[%{LG	-,G??SKMa{wNih]'E(%=7uH,{xPWFZv~?y\#P1@+v:`7+gaWodow]]C#--CJZ\?}4ew[|K^[:Bh8zf]j!`KiT:e+RoGGL[?8B/P~(-_r)H: H//X3iO'~XM`IIAV_:1`P-S "XD:(%|6f/7=fEh|i_iS;<,@7-io%u|+].E^#1
} pUM9po8[2gG{{Bz2Nd\PATq:YCk.OmNt453;b@)VchW'|m&k96VVVn|{w4Gt3iUHoTO_+RaLuT8p_pAl:b)z>*ZyS=ZUPT9RSrMP"f|O&$3l_ry%zTJqq9'
w@m;@Ogx.j0#c&?WBGpXOD7cpffF|vJ#I6#7Y[M$c9KXhL*U>t:@$}F5H"Q{h4qQDiyY/oZt@Ix;'B
*3>]I4Eo\ ={/JQ%!5!RaislJS=d"0jf=z6%a5^nHwW\'vdJW"M9lv[e,_oUqi`6Z`buz/
^0(D(P6/Hbs({] TAyg;}g/Ere./^ Ai&Sl!	a9Aa93=9ZY_ZQ2oOBOv]WsA^gbH7c_"5L~dDs;sl=.#i=caO1b}S2j/)+~nWhg[{;p#/JQ_`k&JdF93:$h=={i>7Tn/k>Wni:"@joX~z\T
^y/!.Ekn:kkoJ&9D^/U0	;7c.&-ZpvK]$us&K9y:Wss2hb;(c{AcA^}LL;O 08}%|YVlK#!Yk3
VZZ	G9Yx >GnX1q7OeV,y qA>!l26lrp!6,M=0V
Am;Y^}!C22mUf.qajd*%LF%$z5T1x>Brd'Sn"R@{6&_`S^%nrV?8p+/r7FrcSqdQvq~h&O'%EPyKr*m>2_uxw|<gMb~0m]3f|?{W\qUT8N{[?l6I=v6/tp69C14G/5,KRt0b0:iR'o<Gr_x{1mX\\";Yzs76jmW6jXe%fG;{?{=_Cm([{E$pm[W:{bW*;mi7
)&B-474ZmN?_TVhQu7Z &[Ko<C/\bg227E-=&JU4h1#Z;4q7>Y*h3>P%eT<_jwLp<HOFl{l:EBA76Njr>_FSV
K_zAhhK*S0r@&#m[b;Yy\Q8&0*{2pkahjLCm,M -2!W0tj|9jZ%Mx^-ep-|

rTh*S9Py#RaO"rS-<oDQF]ijwJ47}-"uK70l9SY~':f!L<1kX)f(dzjZ FTmV^5&/nBi_
!&@uV]9B)-,u|rJ?D[;%bL^\#qd(V-6fM~n<1]D.uw4#Q,@K4mgHRDx"OMAnRxhb"26gx%F~aFTap"t"CS	Yz0oa7W0By{XP:y^SX@=-PN
lW8vK{=oB$vbA4WRqS(5VPXzk.B*2.`oM=&?``:d]7(9ZHbLkg7N.o8sGGo"?@Wi+iWk0vN8K6u#@ajMNuX#E[FrnO3);jCabZ>&TD$fH,{2BDs\)/
H\/r-L])V.=|S9F*z>{6KQi|oZ*Td'T=~`^fBEtskZ|oDUVExVJJRNfx<S:sccUMsTTW~ga5K,{K0A:xH2ll!!C[rv|*_-H*6zupQ[2SD=74{Mm%"*!Mybu)&h\4c./Yy(h"`s|T:	|Y18yjE#-6F+_Y^e%+Gd`zOLJ%jj)uYmtyYgo$$93J66:jr}ky4I"g}UMQHmGMeo}	}<nEVXPw(!Raju\i:Nx	)@{V$exEq<?WiSOX3:fsva6jc*EGN=.*$)	Dh'^EMqLnscK{'F-!0)E>ur6NukiZBc$ y?wFD,U\D+P/VN:6iqNWF3|GI*s-dN/=sRUevi\Kf;8cl!;sj1`X0grVTAE{p4kb|V&&:M/Xv]d[<1^371v) {h't#%.^B	<sG#.7S)TADK4lbn*p+&sak\rE86G09en2vou=>JZRcE,4Fm`,E
x\WP{j6kR2umR]+x+5\r98~,V'32)EpB_I,]c&Bdr"0:IN"dN4+]sRlQ@#5-D@Sf)R0JLyqs5Ue.\swO&Qb4?~P=w	TML/'uG
iv|[(u]KSDdkx-pa)>#*27Rt&p9c{EWTn6"jA[XAj!;&g}NJEd:dq;	BI-_	kxEN,Y-GNAGSINk27z8{Yw02R$*-*0b	4=eupiu`vdmeawpLZK9Gn.5=|h4]a
}H`pSOH:YgZq@5]8N{<i'ZEYi|NRKrOpZ2iHAr"BI8HswS:RWyg@/^IY9'`!NUv`I<,
3xxIk,l*}_"1Mm$P+vsO/jn&8F=D-J{2{(byyEopI{8JDZpf.*Gn,a3,pE,|3Ik7y&iszWkBS1ubJqMeuh&U12+MV
lj!Nre*Rmd%kj=7JWs$)?N'CDJ-co=57*+t}.+kKeup-; b:,afdQ`k7{y%ZM(,f4JA9M3,'\pb#H"Y_WfxKvz#pE^]luIBW~ "I5$i9bJou?s}#Ka&,4+,x:#SOs!ljn]!dRiaXdh8wq/hr;~|F_4=2_TI-uwqnb=[~i(a7JEG!sNX`l*83+)ao3|ytHS|?LljmA,w*4gL_T(Pg EF|U&[SI]Kv	#TWxZr}7IfKcLYO:>>&CIV#Np'5:CTvwu['oS`m\Nl|\Y%;v8vvb9CQ1DkpB(VX$t`efB8X4ZWlq.	5G}C]	2c+@}2l09%TdG]|b\Wt$6&vqu%E[u/tI'#`iC$uL)X<ggf;jx:W3@x[yii"Yu?DXfWOZ8u4K>u+&amgKDe#ruTMr7*gfZbZE |l+Z_	E=3kly})b+yyI/gO&"rNAa+jNIF|@t`T{!{lM>[`}/irGvH~i&ELvW]`0S}l72t{
	%xD!$q]Q/mHL|iZ65p.j+m.3v85am^]-lUzl`Z`K.h"[H!bk-Hc(Ot2\E/6d'PE( Wmc>kOt,Q8aZq~jwaeY6~\}u.iA|/ku3L3"WQ@$efv#>-=G6HH%Su+
)3$}|Y-5*rpm-W)9yX~;?!?xMA!E99'
VKMfJw.'z&}'+OZ-O7B91dIaWam("4z<DPm@M$#Vu]^@0SvkVV!!HXN5hnn;/yItl^#*:,=5~(nfAD\V&aFAZE3t5*tWkG
5P>B11T>R)j$&qp}@*?t{q/onetq*%6tYb=:md!t/,#=sz&(oDKT|S0CR,}d/$\cX9pWiiQW"cr7jhp$#n8nr<sOj/7^o='!:XdwH}kUK}/WcpcSB!!,""|;;FfBh/qg)`W<|hQBJHb#BWrSIhnxrLa_3APt%ZGI(%p+ Sgw/h ATpv<X0B>CrWV/T~kne
"+d:	ewEm?DDX~n7B<
m]t)h3TE^z~{R!PeLgw*<QA:3f`QYs)H{Z
2,t>/",*pZ/,(a{u?ia8zx9	 2:*KcMccG/L'tzJss_cgLFev&+S &[mHxPXo!N~cgpI/9K+4"UM[g]_L%y`,YOM3H@Pvx=7vDf0{]rWJo<M$
A2*[7Zp#6bB31F_LEBtSWY*;SXg0)7N(BSp_mPso>fKa_c[qHc<T$q`AGni1%TMyTi=Sz\syl_1xd'WcNh&UU%%|i211QfB+(%vem.lw`v;%Z|K/`jfT3RfEsk09sgi"^kuJ1ZT=/&m:yXWX*f9mwvx8Mk'O\8oz{/4>OC1bs6k/K pN4`:cK`0%0R/GgY[ SRi|![NXkYW^D*k;&#Pn$urn/l\NGw-q%9 ]{l20&;TvKq|gKt	]i=0(bp(O14{MjQc<gmT{Kk/aQ;k!dtYU;Ro9|?@
P[aWD:EQZt(Wlw~cyX
b{djFwm&lnI2N&Eo6EOkZig8d84+i!6#;82%IP$de:),KEd]aVFUAkB7_WaR;>	}La4)?`E"U2slrgWpZ'X2[p*`""k}-j&?*p99)QF#.886<Og&;j+JIzM29IiP}/DQ,@XI83	BEue%#6_eOe_Lpn18;Gnm4Vu>F#8e\.CTZ:&,BrgC&5{t= ;Y+Z5 atg@BB\b&L:+'[soG
*^\6?5?}U=uVUJv}d,]"`eS{X:ygG9(a](bo'rUSvh]iJnX$J<sSK8O><ax~DoAcG`SQ` H|th|r<~/{19:rUX#|L|aa^]^(dc$Q7oK.-il*t`#!Z\1{N6C-0f_-@0uq2dRv20,
m%
THszhiYT]B.\A0"Vc~]	u')8/&3<3rh6}(Q\LBz<sUd3]LDMs'U)pfRwNZAsi9}4T[$\,&+7EN#t9U77MG[	nLr#xN!1a7`x,UAK$*+q$b:WU#>Xi!SFOrB7w,;+$#1]yTB2(GiVT])'L|q=h-PeHNXRsF9>MPuvhpU;lB2T?uT)/a%R\'(nO<CkyB1jj6o_\u`]D-xQ ^u?}	a\N248.P^d 6fw1JO}TCM}\Q.rsFm*D#c	)!H5C<}2L%vka]d+,_/ruVz<#=azAmY/U[B[	,0 'tSJ`_R:6Cv`v-Ea)#RI4mpXU;T&Vb}N7GKxNBrl+Txar/<"I\(j.Xf 5^l5piUg5R>>f{KEld
]jl"WX@QgZ*,LA"Kfm\8PXEDSe]0rujzM%Fq?;`mV@BiU,Q=j:$|:b5|}i, 	!Y$0pA_|>e^JDUnx.Eh/O?%zdK|2[h1}nXTN1kK9Y
(j]3M>p^{"IlQMvmtWjF"Yi_#y.xGit5%r>)b"c/R}q@`bIJdG3L^\f-M;>/wkvL"uu_gFi[m&+8R6;^J3LvyB)>O}uq+k=c9J=B'.n68K,Wq= Z1R!-__1+fKyI!2DX	n]A>299q#H*F7n$R%+4?' Y1~E6(U
y=eC2%lMIi:sA65[*9J_<O_?1Y*{s(>8N"g.|dOD2pqzLh@1a[Ev.L^{_I*yJH5bjln<z:|ZqR:rxHPK3($c\(W7MR[(srV>x26)fF7#d\3Q>9)m !jx@-+y6i0t#g+Y4KeBnX-ouVBr#@+TZZ@YPZ,e|I#(W-o6Ekf)\\;Rod&#klGbIeeLb[v.Np/uPa1'<CZqi	6E	(ThE=Td_O[@:F}?Wq!N"Re*^,)W88 CMbt2>I|~veS+(!vgr}]mXsR)R*Ypw?e}4!/<o"X.(K$<<En4IR:l%<6P^KV9S?-4he1ic@KuQ};=@JR;/ba|+Zl
g.8`Kb5+tg;=8r9#i2!#pd	TmM23K'#Rk{0n8#tK($+tv
bCmsXx`Fe(NVWm-\[Q7+n!GhndJ_!5&C]b%%;C!z,-|V5oWGU3]>>04;OgyUL-'4>]}izVJ#^-OVEw]FNaMT6U]q^aF^}D~s6{59xX?^Zd1kO9we7:w@On<_,&@XlS;ZzDJVg41X&x-L/Uz
]N*r },(	yG&r8YZ++@whlszb3[b{#@siGxe  8w+Y	Z&{.5Qa
C*
S#r\Oz=0;X2GJ^P4"3]!SgSMt5Iis,gG4b*DT,DK|%P$Fj90.~I2LA44%yVf;}@J?][9V|[c 4mNCq#958gTvr,#3a	(ONRCs
egu-mQb0yb.n):oG@`.VB#$JXy%p!m,=MB|NlLM~-70po0@~'j6=SQ<1=+4{Q` BSLP9bBbMQWReX_*R_9&S#nc[ n!<p%}'zv#o={[]lsPlAbd3l"dA?o?Mk<uoDY1nayyk<:g4Qp8x6*v"{UM[|k|po,-EPOA6caS)]2*.Urt'Q1RP.?z{#	ZD~}tkBco)
:ZQ"Qwx*(`@L>)L|sipO.ZmNGl_UW3!C%yOV5?1iUc$3g'h;f. 	Zw(zrbz}-~\j6VMS	U[.]F{H/@=s~5<v(>,l.i+ZzL)8F@1A'WQ~)acN*=)M6wlsMiE(BFwx}n\[oxpMK=	I0qP9,*e|gnTnz(Nx>B37Ue96k}=Yuo167*:6f:EC.MvyLPCyR{+w6Llfm\Aib{j{DdZ[}./KCP[FU"(|bYfY+V->	l1pr~:]/g@)|Iez04S8ltQ
[s16VJN7~N.Po<odyq({NRvd.	{4O0ee|TSLwAzOu\GA	@-upvF+aJY$\JnLa>87e6Ly}])yYAik!2Ky3[PbmQ=SSGFp[KXgs<hn:[S_;:~-P9o<*teN3r:	*4lq<&V?>a:3fv4A	GrE$4W=fZKs}_ap@;A31*nPO;W})(jH/	'"_7HG(O;|5Fn}^pcd\*=YGs\s _?YH1e	O	g0<9`vXZDy`,=.Zmlka1!^&=\ hC(qj8Hrm:C
On~FrT2(^&\8%{3LA$f~bdvT~smHSAv{9b] `#Q4I[SzF(Pr_BSs-I0#"cIbvmY']/Z7%MU*n#Sov>|n/z#)(
DLx)hi}}A&W3iAtq1]8<Bh)(H^vQ1'?Zn?-z\)^.[B 	C	SF7`]X
\A_913J=j&4hi!]7:t	}XRK(bOHg	3b=]\]8k?nz0rI_4A]:q7Y~rO^d6nOWmXG2qzcQM,2X5$
ae!5FUzzWD\x<S2m5gSTG>gNZ>YGs\D2e@qaNS ",Fx:W4IJ_~	A#mL(z#X\Z\ubihWu\R[mhaLF%=cB2{zpId] z=&d#8GT4`W@Xv-
u'/RDg`HaI|-kWFpp3),zRypI.WLp|ggrHG!y
{$=Ko8`JM:>Hmlyc6}uD8~]3eM/M{]Ylc-Guso^war@NIjTUwS.A>}/e&
\6NaG:
X<1^L8F(sXdC_X, 2ZL493jmH';:|j2B^6<ZnSjL3ANmWE>k[1A6
%#iP	2#}V'T#Nl^yj;JaGP7ixf%P#C7d+\rH.
f0.NPi)w0(2JFW@:K"f\D,!PCQ%2&u"^PrUQh8f)GnNO}32Z-A;+>D:=?\T:6.1z<.'RBQ]VY]i
n"iS2Qm/Zp7pfTBW0T:yuB8o?i64EVd0#pc:cu;LF&cR]"c}s{)._\ftkLq`qw30hUZ(bujw4?Nv8zoD3f	p
sAq)1O'/X&r+,>Y<s)`yK,XL%vpkF&`-:eIb8,Rm!?W;/_qj0I	!>e"
$WC"I6a3*U(y_^G#[^+3@[SE-""OPmlPZ-8>T:? {0vj!5o"<gph	ALE+OCu)X7!u+PI!>y'l/#n@W'/bl3okA=R2nTY`gK[*8\2!M{p9NpEb>qi/"U"fneKCH.%oV;p+8\6LOrXY|F7g "F2o#>8}fp4$d'[FwE/J;gL4Rk+`b]rb^t+Y':08Hw3Y-O-|jpvursxDz#Rd(kuR{Sd<1htGG_Mr&y:{D45n#=u,Dr-wS	:<7o&<3T_Jk|C5	EfPg*6s`^8GI^DzH"T!'MVL<JP=p|@T6\eD(4R<HC,yRwZ,t9G9|YP$nS~1~'}lit/*%?E>_*hg9m}0-"%p{ss]cKkKVUlCApF kI?rcoaG<*9:WSz<o{SGrgh:@:}Kb.W<sR3Fh[p9AFhyh2Xo4B[gyQ&l7)cdY)@GDKnhv'	bEH{5(EO;ux'=I"9xbyr7`.R!Pvz!{Fl['?l"!S5|YX,L!-(sWxH_	A?4IhEK@Kqo_$3BD@O4FBEt&de,AfhRO;M"knU&|N1'`YirAK6=DuB^8?;.CHZ(pT_N)YBrhKYj]vAp"]XjMk5pitBAa`1?Lt5`J.JNe}]64^?2~`ozcKuJ$d[ -k$Ttd..h	AUf<5In/|^xy"OvEY JjqDP-#mFLB_BL|,0v(V@9SY&i	;.>o
q+dU9Rm~d2SD]Qu,l\.V>Ex-x6~4<RY2&C\Sh`t2(5O@If$c2Ax+Uw[fT[4	.2]#D_7I2"kXL[5b;25%|mL"I?9OsLt@u>}Na.Pg3K|5X3N.]XEZ,\;DzDY*
g_IvUu5Q	'R0=7Y)2xtxJEBd|v6h.Pz(NwKW$Xe/@jXsl3VQquAxm?Cw~,yn=C[r3r*uzaS{)r1D!@	6q9dB01X7"_NZ1f?Mm)m<Fz#`=$E!sO^)ebOE$3DRSj?eZ:{:psNi!Lf}R340'JFNt6Up,6?/|HNMzV`!:+F6!qg_7z,3=3O'dxU$Ud/Js^8oH%s3-JWn1=?*+nUx.|Q6X'8<$wi0*Y~"75b9ZsX,G5_It\nwE^D!,0]'"KfjDbn,J4!hd7JCC FV[-S!ot}Y;5=>DR6~(}@K(X\LBJJ0|>X:abvGccE+,vmp2e;f=xh>G+5so0K5f*S~]6 x;1L2y$^]"9 9@hF$6}a'_&j"@q|?R}=KJr4+05hH\Irut>J8BS%DMMqd)V+qi{nY_W@.G9pMsS|V`)Q)vxZQ30%5Cp3=Q
q:B<	*SDHsFD8B5C#RV9SwI`D3VN&b5:T|\3mS#LND^vTjmA#`Bq\#0mvSZsXYhe_MH,1IC'T+N6S*]|kJpHcAa4wksqJ%7?q
w*Q\.g7
W33gf{,oPxJkeE(OHDp5GAox*g+?P"<re^	Gc7#J~ ^:2JQo?}}TqX&0ay&uY|kn\NY$<CT	`M*<
YK%eR9Lu$|+|_p&Q-|uqcO;&D1`Iope}tf6(l1,7W@82$|7rO3-Uu<=-+
+
Yk##g+pP\_aEFLVsNsSd,T<k>q	;ew;=%_'UL5_[-2bIby'B,FtARSf}l~kc]yT1@C<#u-K{]9X".y$~7G*"Bn!;-9:.Nw	%/U@jV-fEA	$BRXg]4w( Fq&|,qwg<b6Wfd8z/(oN2.uAbj
#16Whx\zMV4bcYoG]X*e%.\OhqIQ2/.;i5%"Xex 6yMY` kEm8'_uwrmxusi`R&bXSK3o\eF**9IXGIWD.=_6+{W0y@}99jw11zI1RHk{:M(TE5TF&YLMB5J{A91S}gX+Ead)kW=K4 =4]11EeQhmi#lPXqI7m?gGTntf{[;ZcIp#c0w^cUIyZ4K5K9_H3mVa+H|-UWy?PIFjo!,oq)J%RN!=uIk{uSSf^
e(LE&U
RK/{z`e3c50QC:.J!&1%D3Dse`% oJE 141|J'j8]'P]3iQc!l0r{L^y66_)4z_pl}+/5{5^fIICTvOdCq][#ySxbvx?ePTxe3SXE(Zwy8lIS7_%UvRdBQqSe%=mi=r^iz)s]l1zoE1~Vs>#6`LwDPI3D-HkQV_c9Z|B]i:X_u%hy:$5FGwJ0>S:|R$RXU
6*'!Hs.o#cpHaa%R/iZ3y[]9HhzdE)_ySX*;GI0eH_+L8*!N'o3f3pLmLKju_,|[y!X6?y'u/( q*o~11:+#F"aj4RvGf6I?i)JWIPvv/P/u5GM/oky1).$c+*\Yd)A/b~4^i=0@Xb:Q52:S#+7C=U4jwTl0;jp4ZJQ	sTkfr=a&;to#wn lnBjHbl;R@lQwKaV?|	YCw.hwsI!=o|xL66zl`w-p%=1o6t{I#OOeIh&!TYP(E&t[y_;,UJZt^lp\k
ilb]=)@00n8
Rl>[vUDw*A%SE;6c,DI,$D finWblU~/,\$6DT(c>J3G?[4P[@NEG?}g#AAS@Qqt@x`8\7i\Guu7C7Zqk#NZ'XV|##[Y=,j$!HEQq0}B&TEo7*dmR'woTDKnPhWgbc(Kufgc&^==kbh}*[7+I@?y_XR"yUPp`#!DH.(kaOEwM9'dBxocjFTKj$I'Ew[YxMUiTr	T^ 3^'5jg#h~Rh
o`.^,55-87-O4KCt#*;K&]A-YBg{n"lp+"<+j^.LS)6x&'"X;cVO} Zq	.	n8|e|xxM]*I[&H?-5\vB^[o68sM^1?v6=eUpJfo
d=go}x$U4jsb^PEV(J1nYU@W!h&5d)+|:(w.] wP[2	*QV	(b]o5 puhpKTB\M	wImGRz1fk&E~~^<E6a%}:eg9%}R	R!|-""{XuRS/Y3[THT+0f%9. ('o?
'}n"i::i_j`,ANkt;;?%Cw90s9>yRluu
Ek_kc]Y n))"?zI.%~mb6Xl&pY	O7rt!?Mh'=r.}gr<I=	Q-3l47Mc9c;-+5Yy)_G{4i[,gW
-Xl0`dZaJ=mDIJr*r:^Y8$&1.|F?o0)vY:cAG&>If%9Q/=p)YO\$>XZTN/Gw_C.sBwG]9wM(}iACHBd+e5x^b8DU.c,wRO|cvNpi5wf@)v!},GBa0|<E4'.bo_XiMIZ-G<qQ\3iX=mm\vIoHFfALkIGhA@>H=t5r7^9bIo&B`l3Kd;n|0WKTWW%[*`|f.gV1qcjmeR }fc.Iq"Q~aW4}Hbz4?}f/yw[!je{b[@XlXl4$t8"&j-HNM`X'eTPN*?S;)9>e~?@|HJ&qxgAaMigM40|<qkw {u5lXFJ)UZ6^ :w5By5?t3(B05C(O
{0olPx](]?jo}.rB\%{TPNLYWa5Mh2cbJ?ooKFsk^`$E5o!\UBQ+)X5t3Cxn,gcy7{o0"8 cKuEV0[STB.;-$-Btzv3Oh~{bx*p[%Nmwzq:9Py&<H:X)
K &56ysn9	TbCaP:UN7!#bu*wf.WDK[%h{_ND1h=Z!W2WK?C(OAR9KjbDX_51r[4S:IQ?>2DSBE5!txT"QAnUy@CH&GyMC+g9xpWj]A#35I[lVPEspv[^;|@~%.%BC{fjp<g:}v<l?Kl'\K^I2rU:%B+-n%p7V7svLE4lJ`spE	r$o9-q|pt<(DK9dkQ^MR8TWool*Q<W;6c^faD"mE`5Yr39VG1Zv4Za~/P+S2PS-[[bPq.`<@MUNQV.XAHl+/-qGuu&Y	O@i8}OmZO@`X?NJ1	t_KczkX7)u`:@>f_>]iGgakCV6r`?Z5wGh`Qa-4haGR(-*G\!iF0[;@EL&{%?`9IQw9K:}ReThbi4+BxR}sY\Nw-
(S2/HT|o0K1CVdLnc0ViJ hZg/=C 4vq_Lfy 3zCE7B%J|hdB#wF|_7|748MS	ve ]5cq)s
e%v^]6j>?sL^RoZtay_*NZnE!aLT	t%D`@!I&^!&R#}H,i)^8jdLzk\
7IrB9A*?rc3Jjh#99|E"cNHjAt2s\I(l2HGsm$\M>l^m_d	nR0gaYN"0D$S8R)BWnJu|ki-DfWgyvsw10eevhU2Hg$o#K_gK{DMY,T1^DymW3=`IqSwkr^}&FqN[oB{r=P4JkNo(Y-J'*enS=54o)U`o~rG^zcCE^>-43R^1#6cs<#o<23m%"I^k5d\e	WW5J,cfz?i}uzuO?$J@4TR0WS&c	{LD/pwaSwyA;g^w(V7O1\.mA`9B@chi#>z`Zx.hs,@UuRbBHt/2z]qlv /mR5UV+XC$d]DUsP;#Y&I5p]I(Rk.i<Qhloze|f9`e|F#z4H_c2JZz}gw0J2p7dx0gxc]]kwXf:5;g	fkK_4X*KH_eQvrqXT}(	b+`s`tb~8h]uyO08,L"ftYa@UW8yRJbYjZ7u,]W6!6S_fGe
0=bhT+Yt(8]+qkhX#,S?# qE7)a7,>*6SNbM+ry/2s2iG<e]IL`$if/#Wzzo]u[PjZgvMTU7?57Q	3(%8fLMQxu{?V?x|d}TN~8Yf!MdG!V'cj^p?v*ph>5-cQhaXyOxCrHj3)F:7HwZf-_(oOUZ+]t^f#SDd+5Ey5v,f0;j3="F;7yT,jEb:&UFx>ec>>.#^(fbqlsT0@r=N/AZL]Bs4rt'%`8>>j<9MC1e0^Z5W-n=A	Z^.`710Wb;83CLs[ZenMVoKz6=@o"eBmIG|21Lv0`=?z@vjW1=9oRRUT7Cor4"t$(y*Y\C.i,@6Yo.3Eo6J^VyG18c" _`|'<HfFx],E/O;%YjN5&R^(c$j
5 g?p6"dD$d]>\3ucI-qMFe)8hyilP	hMQHNlo3|2D I3ah2]qH<Zm)V;7_TXRTo7aQ6p8	J(DL~]+4X:/\W|izi\6L'<{zP>?vQ"mDEtj.~R#\{ZZ
D`]B+^.vmt+h'*F,6mB|]_PI)ADS2I,Piomx)9;VtJmgP@Oi-7}u[^Yff]}vkKf>.ISy+$	Xx
0JLn+;UT~Smqk0@hF{b{
y)8cUEFdype5?gB%n$26c>,.08l\V)oBM.X4tJb<J	.VP%pd_'k=$</y7]	F|HibX;Mx}X{|zp|#,Iw;?*6i=j"=3){`no-J%51mXX(4mHA{miQ{
'"nk<IPUnh<*`?@~,j<Vof[O	Cor%{Ig{'<!THC.2$j[qk$`;Nv3	U{13;Dt)j'*qK7	3h&qz$TAXfLe. putWOV*=WVz+Vw+;tb!OIc\H;+XC!U[;]6ehVclu:0DZ[*3mc}KV3"aIywrx<!8Ggq@f(j&_6xg|:JHB+V[r+w\+XpvvUXsJsUDjtR7~Nc/zz!x+e}Lm^RG;"KhNoj
%KRr]/9aP]nHDzWC=5~Oi
:'lir
6S_*x|i+s_6Sa`>)AOO-@8Ez}N~hO,1[FY2`'vC|iCW`//@^aPj.yiKwN9VU%i.X4BgYPj!'[<jykC\`h_mb9co&}^"q~O#}<$1D$hU5V)2gg>!${e1g.e
;Phb@&X0"tmm$P1TC{rU4a>SNKsQ)h:@/,nSCR.~@mmw;-
*Q<6 z>NnJ'KKxJA5H-T>kKGA:xCP{5*fQgU$@LTstVc9u/#GXtD7CQ!5mY7x+GB0`}jnk.?=KT	z8<	#9:+lV>Em;ww`vm_Rpc4]zxWMRC@b"& Ka0MfIP)04/)lzJ<j$L,l7<1OktS\q%2Of?|1A'q+`wc=CaHyC-B["\9zzbmR#s*>0'aI'{6S,wEjdz,gHAh7u8s)ZI'E*X1jl&v%If+i:[SJ<a95RS<
w2Wh:eRO/_5{Y5i VhkIoD*wlkFK
Mcq U Gl2toWU|#&	r&6gB'\*/9;	c	i*GazvRX$0k~z&KIJZ30PJb%<<HD=7`ngFZZ5F8W\;Y[a}[tXD*'*/^CDA<{<]ysY47g,i[?=s8,02cRt_J~PRKGr3k}Qk<cvC9@d
\.^5c?tOTPC_[A6d]J[-u,`\8ZXV4Ht7h<b*yp:-/7r9@FUK?8SE|G@`bcyXo> FgYhN{>*~1a+
$ophbJ7h^p 3N9 iY\u8][O{R=" lG-nYRKU<Dob#jTd^=11~VB2uZ6$9edFIKQge^E>X=]s,!(K{{B$jzbEX:@_IH_r"^*yD\JF	,SM7'5t/LA- LmBor{gLB7x~hkRn'D{\GFG +;M,A@`%U yAD_L:g~Q$Y#`[q~`=R(V"PAClIaZ8FAM6#~q<m<W?VW+'{,tcKAg:z6;Px6J_UZWy%]1R2 }-.Rl}i	p!T5N\iX?8$.:;rcrjkZM%#	kZ@,wi\8/Rys'O	0dq0#SAuF2(VE L!y6\qf_]rd-6l4U _Dm}m9SW0p.Y`}tN*z8MwDB'G5DGdPjc:(a.q2^Wm%u=q.)ZkWanyFH$_M"03K@|@YT}o*'{<|?r>n<UR?hdfdVQeJhZ|!S1EcGfi#pv:/FT-BmC*mlDOk 9(I6[}bZ0)<PPy}pnn3e0+(b[,L&s4gn@iiqY||4Sa.8CX|7a:.aVgA^d]]l,#|2UDw;Y	^:2$%J$_Q~HZrg",S*[-b\1=pg(Ch'DDG?+oun,AjpN_w^ qX84_)M7t@KPj/C\7X8\?[v89QW}!zU$T$fo
Cb{nvp=IG(])?UU'cat6m*+-:K<?bq BYYbk!EEvW.kY!Qf	Gb'Sr%+(}y:rq;HqTr&3Q%N*oAW66!Hp=B-"5P+mo\`9
"{1g)y+cj1HNGl@4.J&~L
LCtKz;jWk_l$tSGSY~CAr'3egLVMafKXbo$u
>	_Sw$q,QPwKrr>]
8D8gbx?wI $>h?vFH01b/:kfrOOa)`ERN(i{&qS56UU/fg_Po1hKe3An3,CL,/L)CvV,<DRv>o/Wt+86x$vrd?jn|NCFZSYeEJ'_KDqF@bH,1hKZA.<3c338r0"})@66H}mO\~*_n<cVZ> pIlS"f^(zs-/i
N9@8\V4kNl6
(lb"PgR`!P0teejXD#?:bsER#CCY9"R,.;?__ZQV h2NL\,H_0wgDk:Zq.@SIQ%gv#-dXn0"{>tKgi(r$,g"/>3f\S#<A54JAx85u=>drR&R @NXA-zs7\A:}DGkI5XReJx0%K5Evh5.5nKIVd
wzW
`F8E@i?(Vab?"u)k4qRt*.RQNRDKwJL8x5m[~;@tTQ6YJvvsuIn>"hO:6+we
j(F3e1p%ep`20!5a7W^t7 k9MHN!l>y6XmFdMoJAI?Ap\4()2lG$uEJ0fY3@=,!DS+]WR&[A_Y64 H(0BTX	O0EW=E'Br"X9WM2l<~&<07HUJbDj@Exm6w~Y$T{7al^,	ii:1X}r t9ZdZ,*fW+']V:PUWp"Fw4=P8o)L1"L.|OuDG(dHzIe:kSlpk>]Hc3Jy%m>AiNTBs1#k<hxh>N/^T=Ky4h`xUrjg|s\*0gqh(q&} 7m6;enK!y$-cK+YLD\@{_ld3._5K*U05O"{gTN:}NWfI[vl"&P|ma}=.tNh*QZ1Jp6Ht|`<-X0vsFM<G@oi.](r;m*zzeJoSOU|DwX"p i,6rh`y>3wo9s7Uodz'}	775&>!G_ZR(F^0;44M]=WX3^X7^&eSY%Y;CYzd606zOBL5)h$2/3ljs3RVSX%H/1mv~`!R5[6JzR267(=Y
`Uj^o7L#Cx!_SM#rA\J>P5@KQDCtp,*LM[Nk|$\$@
/n7@<LNR]#.<XP iTY%0o&(zS$ Q(ry~ @he>c![Wn5iH|#;V/g(eUFVr[\TG{m '[20Q"tT7k!g[8;c(sGDP~O:-TH+]BUN",;_v{ZA84c;.Eemp0@w?_ww37%Fk$O~
m|Ie<4jNvQMnO:V27oT}c5X`+l@>iu="[+RL6iSILH82CU_6{lh*;5
"tdzt74O}zISW<HHZBW]eE:@F6`q{di7r8cw-ah0KQx6R0m%K5QeFs7eN=8[H>zUV3th<0yMIhEE\Q
?JTJ3mRtC*0:4
]sS-H<R&J)y'+E6ySmLoce>iFPm148UT`tVjA_E\MHp-}`b('.8@f}?z-cg]}K3=d);X#T!10uR#7}wwgdI;/mW'4E	:IT`%!I,5ceX@
r&|)f?b?jE]	sf#J||W^20<.f+b+S12E{$~nCDV@utlZ#0{Z(CywBs_SUJT9WHw^h8#^.1SF0|H-)f@5?Lcy1uvaZUlAew;?i{G]Lp"i0F)u)0W-;d~tC#G'-=@Q!RM
6c<kKi45uUfo:7N;MO<*61wXUI(G:lV}{J%S\JhNLW<tD8dv5'{6&X"9	(B4Y4(M5-Vn5 %Gs@w"w`R_ApD<9d?=Q<WSSY3SC[1s6=BnUk${E8cN[%GxAQMO6|q$D4<A`(!e& qAYN0]8oB$+QB
`?75n%4uG?yQ$|!TNpx0WCNh[KNUk&/V7Q~h^qK0v|D~.Hg$y%vCf`tOhVsvic2&nWZc/5 :m#}(FDBdFw6C-&iBel;eOn\G3!`UL7H&f5-L
GY]FyP4}JV%zG]L&T943?y%'
5/.&5[]mm-n/B">*G$hO#u/z9"HZA>D37Wd"BpH?x&2mK|GLSsg]~_F`@tH<gfi7gt(:[5t"]N}:Tsi+pk
P?AN%})YzMLpaow.)X?6(8a!:}gx&eh(UhO:%b@'Xs=F\>,<&"sLoF90M818Ljf,"XAqFU(kL">Hi'o 0 P9=AnHR8q_0! {lj.frRp|,}qR^o]5z`u:k%G0
CL92zrC@xBg=K"nchx	2!PZ'_`9rns,t9ly/l
]*PEC|
!ve[()e?O(
Q0E$<GXR7N{TR?z0|CoM76:\'&WzstPbI2{3V3eTj	$S*Z>L52`Rz_v>5XHD9hvG<y?N]NyMOJSt8	)ZtD&u>XF9>wC6~wUo+*U]mlTC=0toe_A5{qRnrdXZ";<^VXC((
_T=E g|BkWX@6(w9Hhe=fk/OSz=S\ndoF*?+SEpn=C#wxu[=5RTYySv>I;2j<5"'J".pMt%D"XN}rSWG09Z{W/Vg'Gh!!Cn{+^jAM\.mSF`7EhcE
j;ZN,sDZ%{qy#fI*^2e>8xbR{kjg+lW15{u jkl#+s/Oz}~g;6T]ghI>F]4gTPsERLkKue`G4T,Pzs	XutNkK!	/Cz5m/>nP,hSSJ4r|1I.Eo%{@@3I<-n|ObHY(@Sazw7Y&9qn)?01(fv2|z20$ht\Y^Q?ym4g>2B[%JVn)+a B.RZVN-Y$Kc1!!Z)%ER)fgo
$C]xyFf4+$KOcagv2aY^W,J7%-7*\X/ie6:@n}^2*) zuE|$\e}=%"#CopX&*B3jhw<NA=wIj0U9Ws
|Xd9>4*}KfJ)h>6tdjyaxI?:|~jq;D6nLU,ojTwnnV.j+5;h	lVK)zS[?cMw]~+uGcB:"VgzjEm)^N_u77u)9Dt/567y2OQ<z8YRtk1BA
'S;8Rp=X`iBWSWC_lt	jl%AZ=:k
r,Nw`#shDp"}yg3l}+};.Hu!q{8kF5#1)?Au
0/WbLXpG	L@t/)\Fcl5	R!dC.xrFUT(\4}Fqq$8nuAf[}Ft&ntd7D:8?o>>oF5*^6#T:UOoEFfJ5O3T?OY[P9G`%EKOagnX"!"cyx%AvQT({~:IOiL<a:9#EFL[P^SqrHpCd]_SP[B"F:G4$Jl*[]NF/nBOAM\*t&>9+U[Z=aFzv}t!p*A;{,zrr!7rE0e{=9Z5\I#E\"wyEd=\kfb@2*a~i_Y<(giq"OD#lxhAzK.;/uFAUp)AI'q,nJ/ U!Gev,_&{]G*w?'>,!b2<{lRDum&E,cBI@.dyp#lk<=oCg#P?r</p-TCtH_'9kt/]TeqZ2aiwE;}TJv1<93^S9u+(63d6;B`5w4sG\GNol	!7]O|&e=##:>eYOs6P%
s0Jw:<u;Ug%TWKOELZe.cBK9xOPe3n$V5%<}C2tE;k|i66t{=YB;1:E1uj1nJ>eB[[wD*AC|+_|y2S/,C4Kb5G|(^J6&<P{n-%FjXq3awL)uvk"4$~D4Gv})9hQ|<QP[kH&ZHH.8_n	OZob	\#vW$#9>G?E-2mKvDPQW;o}JCO[XI4!pBp]=S3Ynh.`\|u&f6N0
Dk({>-E*:hY&B5.;(|Y,h;fVAwwuW^wyxsv)3BKQ#C'9(kOhW'aMy.6{z_&iI<86#}b2f)ozdj{g|e-x`aSO}fR"F5-1&PYCMho^YS1DY>. f/Fd'V=:.bwxzp4;9J"+x^U<;DUEJrE"bACH4&$R(-TB}yUUDO]
jf@%me4y	Ia4FS1_ 6c?Z}g0p6K~"32;} <JQXJ)w1qcw<LpSJ{ Zp`*BW]'FR %_S6lAgv$IO'%kU*D$eSe18c6+Q#K"TY*th[p#Ker:#cE4BtKsmRl]#!zRQ,W.buZ\JZ/:t4YifBFapZ.%UcpAVn%	]0T3	~A#<~sv#>?	j]~FXl@tlH[#	?_[#V!Os-8sx"~3FQoEH+*DIWc%'=-;tq1T~I)Zr!u{kr:iVb@en<"eu;A/,wLHg{}Wr.+z1qMqoCX5i!JX:+f\qdw&416Xg;w]zb/ %AldqBbL|MfCeRJ.!|+XcoTIa@^j7xG'spd.WsHiI##?Am'a1<J8*k5.s:?GX hxp~
?n$;)\-_h"%5@]&u#;S
hnJ+51Cx!^|(TIHV@aF}}" <CtE]7hN{[F^OjEl-k:f ?&S{d;F4@5@*uCp$xR5fY=,bT	k4,%?43d51f)A*gHF~#-1}s=[Bs35VuH$RDL)wyqpF81F9+<1=@4
+hg*R7+CII_Pe)P?M4,a$G',V(c]~yJ'b)|n~@Ww,r3fUko@|a17Ipf
#@'.IUSM/7lL6=$[tVb`DuM@zvOih5D6GE"r}(HKO*iZV#M;k	2i [}9g>N9jZFviK*/}4Xkh}]\ZC`o7B-flCsSh3i)JE=]mljejrO}:S=kHv!.LMn%W5nmQHb(e"(^IF]cyDvx1@/>JKNH Qc%.7Z	t\\R ]=Wh-CeYZq">AlB|MciAxq]}kE7L8+h#*ic0=R:;)hLLuT;*x/zL{PdS1,C/S]F$r6wk1D_6AQS#8KIa!EgBb^)&UGVG1r:wRMZcr-SZ)?6[D|anXKR&)}c}X.0"zL&+>$#Ht$:d$+8r5$gGHUQpQjk*L\%|CKB|lezZ'-p-`01]0FqY]fP+]fyD>]G`[G3m8#]AdLOaQl=y@}Wop5L,C!I+4OG>79zZ>uWc'm-bT6UpQ2fh(I6~Ad)PxrCX^rA[[Jxu-D{f~J^w85QH&T$c`i.YF	dJZY}"V9s_sM1C-'a=jD}Owf1?[V9GYGEo"P#[6U~k)8P}#S0#	nzN2pzf	i;?OdG^@;g{Qn5KXh
N",d}V{9V. I-[/?5sj$qp6%Jkg{3te .fg8v:yZHb@Iqud{^WlHRD|`Q\vC Pr!&(PS;hD"|4m?"R*w?	guZ+/I#/c!jA\Kj\O11_#v>~PaI!:Gx8Mpve&kQFNQ:C<rRHmO<N	G;x0w#Eb)u6OG&{C^&J)eRH.{y+G|8P$NrX>nv  ww59]y&\vRjP</4(oq#-}MgUa8V;tnYf9Q.k^FJ\ zA]N}O
zoD{4J>E+ax!g7w|;Vq#!8=)9601{Mu|4+:ANbxX`3Vy$+_2yNG4%T/Rum,JbmG74`O6'K
)d;3SPt/(oX%rI|5O`I)C|		?RQm{llF{39(98.L1D-^~yo5id"IW;)t(9Cv snL$<{E#"Ew^ZBpv[>Y@KH>iX%j^aur{1Xd[G7
x`D[kL*q4r/>`M4iyi
fijtVVBp<tUnv%>orlOeIS5LCp7P="EwCIa-~#M:<WF#F/f$&vDPo|jFFg<^*#4#,cFb(jcK	/G%Uz9lBm$ZOE12('@eT9tJ7v<s@X?d\ hbL<F}c2wtA|,/
{ABD)h?LxvTMdIUQ]D)}GNujKba,*~m)E%b|PVNk"[NQT%4P	TOxWiJL%XAuBVNc/r;k^^(DAV.vvJ`F#A8Z,deC&?u<=>&]rqVoX`-L$a_uH$]S&yayLQTfu@<[
7=nfN5|3}fKT`;
Ky4G]N3"~te<h;gCq)f^Il.%@&aJ.8B=]8Gr3p<_xwZ1 u_;}Bs8T2;0OJ0L[kMJ>DhNL$5 Vf6Fs|pgxuZqw6,BADkBC:52i^/E1G6h/.oD17v|pS5@DTGKw (<BW'(Tdn_61l.<OZiLoJ[ao.?t*t"A!wC7Zm4-uIY+b"OZ)
>/Z$>4PH	GbEm_uU9Pa;I]9&{TuZ|feQX\Opg2j@lpERF[9]J3BBX)0AnU"0X8tb#=#kl R,@=,'O/5K_/-w<Bo,BQkNFk{xi1kK0HV=3:&j#5.Z\B"Z."i/^G;n:]'o)"u]@`NHd*qKkEmr*,K;rHv=r-#s\W_Z$<|&#QNEpSAt$4mPL7?*T)%rD&,8P\n{tEh*.Y#W#+0m$1Ge91AuE<DJ3MvJZHm.mxnSYqB#m3(Y<..q*N.BRN2xWe=w;4+!Rf]'(\Jydy'9x*QM6H@,Q{`.x8
US*8Vq>",;Ev2[uISuF6
/>F/\lS8z=oKTX	o8?W*fAC6zIH;2J-}I:m&)*	X'-Q:r;VXfG){;qZ?OL3eQz{Hyxv&=CB&P#B>2^VfXK@Sja@x-}#jEFJNs*Hy%Q~S@7dr,\QABWckA>jQl1[]1$ /j#v_~KiDkci6{uYga 	eHqX\xL2A*Vttr6(Wc~UJM:_m6Ak8ui!4aW1HPLVFsN([(ht2OAkR
cc3IotcK/>_7BuB3BJ?I}r4mQKf/P`$v-Fr*Jy9_jeF&1iK</Ba0}uJ<yS2o!=hR@jWq2jYln=!;Hf1cq5nJ+6g2yIk4z6e'Qo$.I>G-9'{o%]wS8wL<>5(srM3?2IQ0H
iYG+-$v.3c6bN2`9-`:qo:,qNhCGfP;Odrr\"	r>5bjnoLA
nM6gfLaXikY)?<\^URb	(xZ_svMGBct lv>}j2e7KAxj-N+UZ7`[.}$N;J>OCz9NxB:HK{tZ<B|pWFFU:%"GriQ{c}%[+yDzuJ:7wM6j?CFD>7;@)/;njB!!H26^L#$=r+<p@'qb>&#eUO_ G^K-R%-d;x[L*s\cY<9s)feZ9rvA'EsDsd?=?j.VUS{9*2 t;n/~.]9HO@QwiMA}9j$yex6n~h3#ngy]+8LjRahlyUM"{;N&I-*)n	exZ0"4s5a8B0%it'ah2d=0*L'9:g(5`"X;pW/|k9Ig8#o[at\zfJM1c%xJLvG"cBbb>^#gm[)f!qZ<Qe.:,Zds~|c>'Y&0Ia:Gdb`jiX
KE4v5$%YIF.	m8B(w&+'YDAG@A'X*maj,)&Ci&9JJFH=NdVmJ9bMQ,Y 1k$l)}.vo'3*L2L jf3BWbn[9Zza'a	)$Rj\jtHw	Le({etXTf.PH,>SJ'0<Np3OCH^"Ifqx$CL{g-=m/6H)@o?L@9G\VVm"z+Lg50*fw@+vx6DRS(	HCC#?;+D8?}e%lK|dpE|9T]Dd:6o|wb<!Ggbt#/P-4A6-?B4:YZN`he`;?)&nD,Vk|P,rVFmwMNW!1.2"V	L^^7/`!l|7DT<~)ir~Bgm(	(OlX|ZPCSe-Ul=>=+iVPZ9$Y/t/-;&o89ps.n>"eLs\-{F0wpwodvEXe%Qb:aG*z|SC mfJz|".4_7P5.iS-9~~Oc<,I64_i]|Bx[D8m(8@a@/Tfjol
L\'9[HU4%N>=~Q2.rV!G):5u"7?\b"(`.^U>vEng;avN.hW`=S@*,oW!gYS6n.DJPT!,l.u|)'rnr]w)/Qdf,q5ej;+~iK[vWxYorqPb7]cV'mN{ ]Ij'RI.
n%Gr.aHV,q$jr.+G3BiI5|fV'ih\(h,AS Fft<;g\W	48o{ml*|
3Z0)
D<C5UKF$i	(k[*TH~x<O~Vv_1L4cke-06bP.bA8Ie<wfH>R%0~:c+5034RL\B80[*[W6Z6:-?-nH^8#+d8ukp}p{;
!`FgfX^ES<
"Ei;TnN0XG1>\k`mB0tGq.xU/}OuOjf8e5FRk&8P9)246ob;5iLBtP=O-$Lnv@R<t~ef2-uy-
l|w/xLs{1	<>F;qn!u2xQ	O]v+~k`pN(g%?>g%!1D{c(
t1u$[7BU"Mio|u]%CwuJ\V7%%67c)ABk7.U"|F!0}In0=Wy}dy-<Ni4hU8Ya."?{zB/	{V^F'E@>)<GjT7I3KhW>(DSZ)b"%-Gwg
_64GV8Ecg:
o43!nQl8blRo?(9,n.CZpZ?ZZ|\~A~#\v()dYJ,{rI!{F,,k>,?v"oKf&&G?}"Xlto0P]ADapkyAXpoW:@ ^z3m*F/V0=DQ^+]x}^wz:WS]m'
K4{av'BWi0o@MEx5;({
$f"'SjZ}ClIU>f*Y2c>#uW{9p`&8Wah=laN#nO>)'
+`)"5q?x-O<i(8t6PZ;S]]Jk{*z,Hk:n+Rg5iM6HDAM.ez7bik]ko-gjyIOLEIk+
A%+`}$/ji_O{{).aLLNV3*	fuxs0T&aYM|L3SL[Z7u:3EuXY}r-85(> Cf=l!jOlqU
/`IW"&F`UJixzJ5]9M<bH[a8'^:25DH5"Jf.m\F_-9p1P!xOiPM%4}m-JSkTM[3nyZ?87z3j1kv
 &<(g2$!64JPw5.OqRCVCf=|Xa*y{[ pt[EiKhV1}~-4WIdRP*i"{?+@O"=J%hf/kLiYU?
/,c:<A?vAGoy4	d$3ETz%|p$*-Y!PJiI;e0ia0fgj2f-%.pMJ:H~uP3's9i81IP`5bon/j E>]?FpCxiBhcAsX98Jt
8jM].vY`!h-_rI$R&4X)_h$=GVind)*(.&%AXNI]$3qtq^ "WMk|{_U.?Z}\cos^Wmaej+qnKw|~^8Ad='@0FlreYI~qnv')UP4yw"7N4O*Tc5GmTIHhy9
0Yu:s:k2wYhkfb+^stF%cr:VY[uw
<k]Y`!aLEkg?Jjg`FO,+5XfRR"8[$$sliE?Ih.O1; "yS(P'}s]EpDY-(i|$<sn5C{E^7@klP*jlF b'sf,l\v,t1"U!7F!rd'b!yr;3ZPgfkGUiM oWb{:}qZt?	!F2f0qg{-y79?tM5~C5C+u|yB&<[HQF7Mm'Zi7=V6_I
z?MT}M9$d1-Vh4Bf]41$~l"`plJ4v3%rd\	xZ^Yvavh*EuwVlB,~~#cck+Hsbke(z?M@_(qj_6YR}DLQrOR{mNE"!wr55-cZPO(ejQrt5_2Q,6/m+;-YVV)Ic`~F:]~*H(G3>^p7POi(n2ieT?!&`xV6EG%o2Iv+_:Q._o}l/2$	lQ`;ueX{riqmj$ BvZO{?:,2l1J|tQ^sx
;	99k&G7qTdCY\E3[ZS!7_;fdzf$yP<(N!kj (4Vb/e\|$hVyb
1Pu/S#_zR{Sex=*#{PA\r/4ll&1qii6$XhOQFF!&R2wFEzym>h(C+C"b+vJu|1\+L:]q~'3q\>+4D_b7NoG]n\D*sSR\?FN%-CYv9	p	1U	-o9xC#4v$3g`?n81[?:xC}rMbJYxoUo
6z"6ATQ
vA
SNc~)O@(qvM7'!{e-{rOmKT]LPA>	+j80,YCEDb3kC=DZ=UtN3R!S[Boln<Pn#4d_N uCH|ql%_NkW9p]"G'{9*g&f2m?A--(1%B9@o`)q/Su(txQZifiQ+}+M~D9iA-0TzP~pPz-=+!^[(6/k\mGa+[ihGXU3J~^lE.ZO5G`k4}|ajqTvLBEjb!SFq{6HyI>ac~b?:4?NzL3o@%==3vS3_agm40'{cwu$Wl`wp2[BUCdTv,?D3@?U-rF?a3t3R} CV<JJ::z(vR=OT60]g&_`+hc7eXKj\[b75-+C+9"qCV-F}>;._l]F-JWP\H)TMSk~
:|TF,lqtC?)p}?sVn.nKXS81(M+
7Qu_8FP}d	@V#Zk!ACipM9jhF4c6s"`/@'=P~+a*vOOez<$_AE~C+),$k2LvrIPFQee?B74;y$]2 ZiEfCXpiC)[mv|
`o	siR!uc|a^WO"O)rmBG~~",,_6e\U\U6W>p
m81%|;=V'F'A$e+WWB~
4YJ7fylDA BrVL&\?jl5r(l8moKt0:n"]3g	"4_n/9ee.riN;evH,:C&8u(gAqEQ2l7*<S.]h|15uwwWA5C\K"cl
HU'gzmqXnG9XO pc"V<"	#v#PHCk:	DW8cS'U3,9Xp<)2wO{zhK[O>Rp$UpAM,B(_aH5@UZ)I1z+2C_[u{9YLE92>M{7@NFAQ6L)<ON-TC[0tsDwj\zYGYh$YN<rLoc%;tXhx"J^BRO;<kwS/+NdSaWza%~TJF#[R8/9SL[u$0\dmy6$x`|'=~i/LV)>hywzQ2^TE^IN
-$bFYST3[xc`wAr5;gSgB0*{"iwSCM.RIPzjfz'E!47AEO!{mqHyUj,MPVJ)Bkd[5%!px	
;<k/~E}9veEIu>d{=s+>:rTxCz]uKV069ztSL/y#Be_khjFD5EAz6M&h~#Y=i(7oE&1k76@
~T`2LfU'hFFfi:C;j[aBa||ggH:l.qMk[Rjp#OK_*9:xgQ<U[}0~Zww8H^5WHis1lZ0:1u+I>A]dc/v^-v>2vN$zg+}GN,Y-C@	@Vb=rBRRq. o70po1L/Y8d_
8< &i 4vQ)v-5t;zJjC`XZ{7"$pho"pqSK%V}K\{T8C\UCvHkD[GfVDb?K!d6-pIEtI;(RtH(@eNXs'(*cBzvb#Nnf)RpvE'2Y+;k,)KzMMU	x(r% 8sPL4]:
XM]f<E]CoR/"Vlc9L-Xu%\1h%$y(2skrN	&!rxkN$AXk9R7G0.ek5,q{hzT%\q,l5%p!{@\37\Ag{Tz9D^f<[{,z]=PL$,XY?	r:_dBJwHDO6d|xPT~\2n1vUxK.(iZz"[-He
&Q2pt
R K
zn/stco{V3n0+Lv"@(Ly7hFJJ{s"QDhS^y/AZPT#Jdl`?#L\z|&YUl(kLFT]11OPOl$9}Zd%5P3683y5[5L3VNP5[X@N]EB*CQq:{G-Ol+(9i	[)GZgfH=eA?jn9EaK{BK(c[oZsqnl
Uu45!C1H7V*.!*PmD"3RocGF/Kn@tC`0
hPo\r:)"pS=*itYT5d)2E~v^&>=Z,RZlB=AtkMu/jH)2&lcVOkJ7ua^f>f|RFt+mw,c.0
E7 JwA4Y*!3Xp$F=4[EA`*>@_Yb;MCA&@G'7*.K[/6rz{)n\vRO*4.Q}jthf&;Fi-g/7{YvvvWr#(GZ>vO<	UuB}S5XTuofDh2QW]Qc}F($2f}m#ProI+C,(;J0i(
Ny'9PWZZP4NDEf6Yn=)XbN93D=Lt$)5O(`cuU<#gJ}pKzQ&\f&|pfH VVvNoXa	Jsg|vn&jb>/"Ty7Uv/*8 25^d,aBuP%_J419;>xoKQ@<@}`,p :\e
.qNS8$1&p^n|sj.,XkG;sSSsmmRv4p,:@2
%F3}~B::\f
$S|D"Xm#WntipLhj\OA.H\?nl:y/ )c0]8t1@g;K}<?&Rc>c@a>?y:~}y:CllWs%*.G\>+T8p{ivzg7Z2eFP]y GO]E*>>~&@Rf$1oLZO_G7/Q	aN<q08tG1d9fH]D5caA?=.}PA9bU&JJ6/W?:?u"&wTiEoez!xFo/}0->='Hia\JPW%RtcEy\t&0
5gtLG{WWBl,ec'P?T)LvDt(o-i8fde_5G3\tt&N\"xjP'5{.^2Ghg0-0)13e+Q{(zT'_X'0,klR5_X=?+Ql!0"YPd^UAWwcu#@.QOSa6>}lBQjjDU!_<(Re|Xpz6Vr("JLx9:568_pGEDBo>;>8e/$$Um	S(n[9*#''P:=b`P =?7k<1\J6{X"	QLF-0,`CBqev~I@bEQj}<YE1E?_-)Vf=YUv9|kW>=H6.UHa])R+v ?L+iH"*${eNk
?SScL?R`R*,fOGlMCPI,G-furD:V-Vgi	|8o6@9 eHw]7 bU)yQYeOoz4]vBzpYm8=IaRlQfyx>zNcI+}DI?@g:9sNEb2%je?7P)+SL&PQXLZ)!JTB//H*?f7$>djxR)YVjCHC4{;3ax{3$xImgN',Uq= 90:=)<JYEfhx3AkK1<k,SFPp !x7}yG|*W/79|%Q_Ur={mL4mINf"K8&i:	+(H)6qL<}NPG=A5##:(A!_v{Xv4\Wrp$UfnN-=tU;	?T=Vn_*um2tC6d<S\_9M"KCeP3SBy
GG.=/`O(-Rqw9<Wrv#d$8<:q:
D_,bful>Xo,`+9%?<Q`;&8;"sz)"/^#oBl<sg]y,L=|ds;Onz;&d v`S'qqAeUBTJ:99y7}-j:,}R`!8J"M_{+'6(o6j5lqd}jBM_-$S|Cr3"5B-^Kdb z<+&5"3_`#H_=_mA-hUT{X5'n	l#2Qg760Z-kl'YL-Z29.I +u T=Qj_(9&XWTM-=J&Ik1qotyyKQd?KUD^Ga[HLoj\`J?lH-)[gee)$%n3B|z1=HOi {mja:E=g0b#Z&MLjUo'W%*^.h&3dhn^aEji:"q)TK$|QMt\CGv3j\.hK	V/="Pn#!2Wsb084[Q]!x?<2_q#
!K$.^dgct3$	%^t1
p!2x5N=K2l[3@4oG{u>DB$E>$!IY;1s5cx<i6,,Yb$fe#Q%K^g!Ka^r6#?Q	BpZf|rqCUJ3uY+'ZV\M,W,Y[^L3{q6x7w;)N08
&.oOX_wKr9;Y_B	nQ(?"YZD9lsdP<P1F[(,yqq}2<CB g8M"hU@g0s%'M62w@L)d!J