G6n!BpBV%Hq1tYtSPSy~!k^W.qU33G#Yyy=--Svg'il$enn"|h}:wWXtLv%@B*}3:Mnhaa6*UgR~HOcd/gj${n/4:`~5^]"8sLP=Ci!wU6)]bnk---`vQ*M#pbLiG~!66}	a;28MUD5)W5+cJXPK[?v-[OZ,N.LX&\/j2/oL>Sc1&y{ tT<Su>)i0!H?CX#z:[]UpFhC57Dp+&)lH2ZrR!1B1lUBJk[noyuX
yy&PzYdLbvp(#p|}6$tDB5|/O'Cy#:3w~a;:^IG~m+ n=gf .tB*P1V1=J4/@)'zWp;8Nk3aoNkH|vjr%eZF5d &(G>om&aTt<=`8o[h})e$KsCpvh!`NmN8"1QTRy}X8w`	1g{>?Y!$nB:7u<\hhh|[l@yMz-)x(7~t}^y4"T.ji{$W?CJ`/JFW4Jx7!
Evm'+[Q}W_'nr
`{)`MC?r(mxbeT_1cwa$C=E#B[9CTUIDa"c]Bjh:g0!qiW+OC;8bwHkn1BP4GZY$W!K55Mbc/L~I<*Alq1)~ZH	$='T0hkwM<p@+.10B:POHV#a%'  9F9&aNzZ`b'DQ+S=
a7\A 1~Zg`9B5&6/qP?m9	i[	8UsD%C=wEQ0]j4:q=U;Y*z5}s6/cw7H[>->fY1S.rIA(roBKu(o_(hTBMz#56p\gc!G/6Gn	'w?hp6yu1"NZ /FS|@q(1Br.D.}+q(bUmcVB)!#!>t)8KxjxYKMgT:6,GIU8Zte?I;_h3u/%K.l37jtk{>yNp.'l4q/nYKY$CK$q[iLX78>Q]z<_536
;:i\8M{co!UwXYS*S-c3#OGlL)NZAHkJ|YCd{Nh@DBVwE;>LR='g0z8zDwe9QF#yK<`+vt?%dg7'Gv0AdGr\<0f	L.hIp-0qlI)AlM4gNu1GFOBhz%VShe&Xs>d8=-.Ed&EI  HXJDn:>IQRi3|MZ6$.%DmA2msnOT+>	/^`2"7>zHE0Fi`W&``7<&|BU\m:L6#yN^1JZ$tovSJ
QN>[2J3v7/3%:,a90R5k%>J~Wp&E1=c@Z}*
]H;)R05E_)nLJ;ulW%sn5%$[@]`d!];_T{ZDR`{*N\EQxzPVEvV=ofZl4O
p	WTJ"<!CwEj{1'IQOCQE+/Wc$bX:$j39
lK;dIu%`$.l&leh4
vl`>UGJ9	jf*b +T}^XMGHW^xK\dyZO$:SV[bpT6J$J-CdlpjkDZb}d4y$V/JuV&Y_YEFGw@eb'yx8))9ELw[tDd2;l+6yUE'$APZ2
jvbuj5PNptj&Isp|BA%.5h*>!jyrToMw7P&VXJ)RH{;ohVL8V4o}V9lsf^<S{?d?Kj%@$Vd8i<Vtd"7w0pjo.jq'iMxb6w&0 9cP{g+pYz8b580i';qNEYkw_f"t_W{2}0<8=T"] 5a~_c)t=Q3W8;$QVKqIKFQwSGT,	jTc*X5`oX`Uw!G2shpbaR_8fA^WC@p]i}EbbQr_;m:$c|ahnr!Y"|.MF3k3"pKcDCFRHxYU^_2(	skpG{aIkG> AjgZs'O,D6odS{;0N@U,4N%->9&P=k*8xd4:m&JU:	$uNAK=gR<CfNKs%i[+$ p_|g;h/c"|b'HSt6m]f^OU:]1/~5up')JwOh~azsN
}Qs5b>cho-$AT@!~)>yR<-#;	-xT.=&z"yftO6!n=5@w2}WwLw!.C}^E&StW+ :;
+<wz_wYZT@_*,5:x?n7S`N&Q_%W+[st7ImHk_J*w-*Mz	Cn/ll.biQL&29mTUeTb3q'BnSHK@Z%E]LeMr}"!UfCWRS&a59~6g0[+NK~AUB;X?XaiR>Y&[Eu*t'_V6\q;rfbgGh[n^J`gy<$\)z:e_crfG.[.^b'73G7"CkAK"@9FqaCwZCpNemSdlTmm1y30uL`ah,~bd5)mDRT7v&w[}5#^'3.yO`|ITVTrdhp_W%ym0N\V:PZm;pIm"<.@%{mPgi6nY[mS@O{Qo8^V25vxM/?!t$k_VQt{PyjX1R7k_Qm4F'CRjC;?LzG2WkFH{^NZpWBJUJ.Zs!y1T_YhnQ<zoby@z4)uMh:N
kdM; b'=:o,
$~t2\w/SE=j	="Rpl)cGY%68~XiY[Wh\r&>Ja{D KoF%KCtyB~y}Lcd}W;Rna'YLQHZ-ObGodNst&(/5q c67**(_!V5qy9IW@2[}iI;Ahe)$$V;	>z=5pf>EUsm7cV+?$YtcG%!EBkr o;Ic;<?b(W$^k\v.5{!~aw{;`w	_DI#({;}}#G=D$CI!sixr[x0.v,wI%>JivrX7)?Y_=T;WtX2_M6E{e 6
07Do
->XH7B=]rXUur:C\\0-urU(oD.^GC]-0FwGCge5p~_5uo3EE?%WbJu<`s#!M#MmA{%i`p{&`V6OBycoIdKak*og5U0l<W)ZF?3'zvWGXmnCRkW`
`Kg$Q&5hOEPy$hW-w-@~#	Bf.	8;]Xr4)o=hrww.^!V#R>4`J@-^v;o^%s/K% Xhl= bB[d4d%zVupf#YE^K=6E;GewqV,	xqwy2OK	_ou4nqw		r"d!IORZ_qX_GFw,.IG'yBf&2";alVaz-\mmK%q8N@17MSt^^j(\;U|TG%D~1h+&{v'*)x}9>H.Qv+v"j#Elgo_%$DMp"u?rA)Q:g]9 mO$mjNj]H'_1gl|bpEc1El93^z+]<sj34~D89#-EO {bo]	S!0+Y1,.rfJl]uwx0"|3BJ9.Mf z.N2*[tL9)RoRib,H3PruZI*?Yi)7yr]f[Chv
[_R_}NKF(U=
-D1A!U8hroA`6\S5VccftmkiJ|${TUFW7lVqWW.#AuZqb:
SSE@T8OJZgx,1Y']tCH*7	gG0qBlJM.032R(N|,emi-fz=PqBf$kG=EY*gTG]SZP|D=G(5kG|8j>
sAH#5}oYO^TbBq.>Q%0Qam61SQ@?Zgj)Dp<b4<O*%k?8!|E _^sPN-k)a	)mK4w}wscz(8,t4{-v=HLu0uLa 6kV[!bDefxsk6@^xR d$Cyu+>"zc;<M|%m14uH'"JlvpOJD@Lnn1\Am*iGLOY5|;1n|cWQBelKU1u:TF;uS+'BS
0)zs~BA}dpFNmA~DUdk*5@
DDFxC>Vdkl?hmZ1~ =3P'v*LWMOX][03H4O.5%4apY84.=KS\@-Xd%+^N#lXp!"75[*_hf=I/v}
U4D9:-qc6WJ1*fsYH'L3oqmKj'5`63h0=U|2}2^"Zdth`~iKLq;vRze;w'G#'0?Un}qgM>uc{`Z\)AV
-yCAC5QsMYKX^<p<@^N\rm9F+zp%aygP]pp9$@`+'PT	m_X@Rch=6B=R'Zu#I3fB0\* 	Qox?#KSFt&ld]B4v`)n^WsSG
bq}sDtWx<~Fc^vGW]blf>(92l0v)76Gr9bD#*yV+!1x/QR3@ERo$`@u!wV(BLjmYmt@w"P*8hBEVE|:V7R+9aV/y,d>x3	|z0uPsv!U/@Zd^%DS|tO_YRPf~7{Ent]8i]e#FpHvNf2*! a9++Hj:[uQ8l=`Ld2cJ3;wJ&b=ehgH*9+zBjy)mLvS"IxJ3;0AyPq+5H&l|k(BBI)v!<Q,Nx!:^kYY%*~'aUR5r7tS\</Ofb	$O~^&.5L$*gYwE[uc-/!@OT~	$	>)Zi':ip4hBvs(1k\X1FjT USy40PbPR/Wox>*:n!sh3G-~2]xxoQ&I[N."nNY`a;zA'Dg&(LL4ey~M5D\,D}KSe.NX%(G.
$E(nyusB(V]:S{VV8KrE}i_~Wh9p5:%_@-q&d"e$2Yv{A?[VCI ~s;z?yk<5lsszO*oAq@xsfC#m#ayK1-]u:z7e\]?>kQ_E}@]nQEjX9;-[12Z[5	3n
-<b^+K"+.,V%xiKID}~.<>Wxk/nQQM;t\[seoW+{xL"'0Rv3%C5=DJ*yiM6hF_IG;?wW"FV'p8!6,VHu7{J3Y4?	Xjja"ZY;bxMQ@4B*i8d36\e21"RJ?-,E{tC
S,/BG8C(Xe!B3Ua(Ua2/F;PK-C$wxJ#_la`3MNi|$1]~-i~a	#!=EsHfu$@]a<Gs3XvD!<UB/TCL-V|v3	;qEg.8 0gbZavj[1i[$gX}*-frUvmk+PYw
_rz1sn,s{^t;=&i8KrXsV"-E0Kf72C9qu)Rag*1)mjK(&E3DdEp	DfouP2dBB;`x9WK}Grq?7
1py)25{,6AfX_pe6au.*y25@3}* 5LqedKH]5V"+9	e3	Znk}TJl$Q!iNwS^`*)E8/e|<.#hiB!VMSd3ho!~MgT6g$D1yzpZ?TQQGVR	r1A^Hj6U}5R>mhpiY+;NA#{|nfZCC[/:?sBem H&Npcnq4<k;,fDl	daXm%I;$%D-T"q3Z2(qJviw[O-^_UGMC1g1TX7pJ :JO%!ADC"	,'i,+.&3~>!"k@nM7nM(Hy|PC2`Qi}Y;7uQjS#fOA=(9:>I4|w82%4-''hbb]Wm+a}unftHv8-hq4yI,^I^d]"8Wt>FWTW2oSz;LQmoQI(]kZT
I\&Qn$O]QlLFp9W0P+7-; qE\ykrlO	KHrS#}0yEQ;w"b[.eH|u
"{i
y1sf1=46~.dGGOLGTM+"[}To|1SDYML[.w@aRNVozjk/fK/&E##u|5e^)|#h(/Ps|*c,~C$6,t,C6_Z9wECnvPKt,El`"'&BK45J':STk"^vk^n|d\KnO{8 j/Via7{8D@Qa	qo~IS,hF?	6U$bGh5p$%{1j_f}hzl;2]s5]s4D0tG
fZ0n^;OQmHhXtad#0 -Kkd8c
@9'tZp'9D)g5~Qe:#(0:_,7q^n=}NeUi>w$ixA!*0Ov2t}Q%s2P8i2	/C$bo<Hp21YCP3DS(@W-en?LWGXSOSbcLU5|t
UMb%o=>nNF1L;-2NAena|j%6kAb!rgM
l JK ':	[sQwpD\;N4TLyP:	rfu`EuT\J=wVptN^W]jydE^
\ff'Bz2t<=O6wkc%%2t7y\V,@|%1BXA=s.+t!aIkK1@-qg=~AKxDd-[s}eibM#X
PBbUfmTH0/e")[z$)'Ro#7R><%fn;E8|t1A%=zd'2	hN	DMyFv&V;@v-]bga)}7S*`L]-9\TR`z h6jZ&V2vj|W,n#
"+PnHZ5yVX7%+`ftNg)r`.fk\F[Wu8#vp?Ra\%5Nw\?GTY,I
2;whz+V %#0A6.=.#O:E)Dc:@	)OqA(l=2ecrb)4M=f/xe-Os&7-Ozc[H[[&>{N~1'`ls`38hLilJwHKKVhd,`]yq8F'G4kv}r3&_H#3g[ny6IVk]}Pm]	aTq=#z!8xtpv!tb$!/@%dx&i]t7f~hGNBE'7S[p0@|dJ@GtkU5g<lTLl-+94 &=[cl)t.@Zyq4e<@vr]aq<W^6hnE&@Z9sIm!K`G0?wO&
{e/(6%uwEu0`22`aKugj<wevTrr9^FA)RBzk,8_8*ozC];|v\k$kxcu#%.vaNtEp-)p]!7#6$vN$Y-a)L^1FUjVT(ki1ihW*fL?MouM\~c*L?sj?F;?
6346AOAmN*sfJ.?J]9FsW3&7]RCgG	CRMqTN!yz#A+(E9B;4tPOu!qhOaXkp&y~GMP:cV,"?#kB*eri! n`ZRxQ?\cyl&{_I8p|8{Qd]TFyuTGEtV:D,6"kcu"ungCjB$H#g8x(jNWE(z63^}k?un2SG^ZZ_LubIIYtyAEWKmq5%meM%Qz*$3IeS"kh-~<=
N5lp r8|Vvia/<}OEaT`<3W'03b@g2w|`1pap).&=Hv$t2@A\.9
f	zz]=N]}ltE[7qw<~#3oS
lP4!4-qHq&#7|SUb1k}3^VB0/j,imXHp#![+"7(F{+;*a@r<w 4bHH [t)/esgJFnKQ3qoRO+;Dr],3NV>^>MnivuPO55ct4DqTsv!%uOVTD`/+J1TEBkO^aT
r> Z3|&<Dne0dS[^-NB6"up5:IlU%
feQ#pK_%{)q_X44Vfl`@<iW("vTQoVImIw
]BS;KzDu'UpChx0ik|I9+!G&Gn>a\Jzp7b8
?C?Id)jk[<.UdaH;'6wE77tbD"8*\kL"A*N&a+\5I.DcOA	Cx-RbCA%umU."}(5Tf??31/oAt`*S+C!{vgNtM--:gv\wKY9lPK"A@?>ec?q79
3_u*^%Y5$}q3mRHCaD|JRftUBa}nRx9t=Vsj+?b@:FOgd\x7{YRM:<eM<W/p/+9ZSRHx3:`:^v`JF9!8y/NGU"j^<WzL/?R-oZcLCy.N<sjv8?xPzm/h5-:jE%J?2rFjUFgQBbhx|}FhF#9Cp,t.Hz]l@RZ~T;7zNF>EJ|DEaK,%7[!d5wKa(<E.Q_kaGM6Z.|nF`NqL8B0Kt	1)B*ZX::Dy
[\;"<o>+oIZUhI;mybq6(T#D.h(Ff2#(?VNEPBnhrP72;A4W goT:VI7$OhpHcjsPm>; K|yjIOg;j6!|Fp{">[K952@lh&e"C2l&=|:I^@C\\[O4giXPdbou5j}JYMM:Rf|MQd
g%9O"Z*MF[x4qd$jFkr1at.N0%&qhOt4$% eX]F|1WsWD@12*T4RZ	/2@qRe-2(	bVDgho$[&2I@`"/qFb,K,pdOif7XxT-wAXFTJc&+:&p6vW>.G\IrDZ$!DC zLO9]&e
:4+{[X(-L,0;@k%vO~ca^j<kN @5j<3\ZzA
z{m7G|)$MMx-,du5}Eoo.J7w;Ba:jCNq
)Y4~HJ3aAxEKe`8L[fvQ@0nU2>s#	Z`q,>-h=`r:*Br*t_Vj4a8ilKkas9I_T'xDOO)h>&p=V{U	J_gTz}=xp]2d1_"t6>dv-:}&$#ufOv*U	HBV^c>&<#,txJ.a23)LCow2u\;hhqT$AT-@Wp`D?qE!h_:0-@fT&GF)-<A"et<3A[l6.eh31i{'6@-}1Ank8JKD)T	)@q`]FootMr&]5rFhhr^7yc%P'_:2`r;oD|'^C}zznJt'P8gTb]U~N}k4k61D'/&y2N&iZ=,lVI9%`.*xK0[T@@C;2|EA-62(Jo;1BsyK@#*/t#}#|*NeM|+D{f-+|;7`D59l(fEIZ3D/oPyys8+OtE:J2;lSq(/shq1'b7hd\JO]j$Hj)tIn)Fc:0yQDxfqhnr18-0;G-Fi-u*lzER?!1Kb5&9x(?y!%1]j'FL]W,iD> X0/EnXdU[e~@_,)M2]<6K+-i>R~p1`*[_!Wk< gQ+Fxlo;9|	$h=T4GuR)0<aps]lj/ep#8bE>->1jEngI=y*{\p\y"wEnVkO}[qLj(SZ2v
(Ln"N<K}IG	4lyj*NS.|9HbE!];t)*wP,sr^^3BWWs{u`@1x~{tsL@qCV!0;Y4apo.8Mj-3dCLC`t>*?mMZ ;57tM@Cx<-4(/L}6/ 	pQW6
O8!w}w}?"u'qQo9a`7Ifzy=Uu~2Ai{&@2pHqn;4FmciG	[sia.+v^{\tQJk8)TlG!;@4))G	&eYqDaru|ht;(hX>y8>oL/b@6c~f%A^@7<'/VemI\}X1"`[<j["iJ]DWj8so25wqoog%j83(k4e1w	 zz@#M5m=*`VJ23 _\G~/!Id9o%k,QUX>t*_g|JJsxH'[.k~d:o3!#ponq|j&+qgu^2.nyB[1rV\U-?WLyf$XID['Cul3$R$_wn<+?Jq8>rk`C0NfiKH
VHmb+t51RLhdCXgNJpzX%P;6!!T	&!|f%`.8b67nV.0{=GkW++fdN{=p2,D:{70dL+Tnv@Zze`9Ub63{(hJm4*~>aTgxtM_G,nF<!%(lvy_"*,4(n.`3V;ajt{L-#A?H1H3kstHP<OyK$NITO^Z]23f;6NED_EB\K;u<,
OuQZrPLnK:$USw}$',zBc4*7,$3yY7Y}+kpfQx'~"b}dQ	D\!MGg':!ZO4_RMdj8aWK7e.1sl$-d<dl2M8i8J{A`Ry#,j)dc}pd>fa]Z\!Gic~+\Nu18Om(?]"1:5/Tu+FEID$+bxNA\!Zld-,qoO	2j$B]Z5fV:o*Ohr#|j~}We_W: eCB<	`1l0Z#sP	M4t~{+'7rPle65QEpgJ9w$KWN)buhBXroAgp5w@"s j9]e$=`*!)ldM'2MB9_a?N.xO?XJ)/R|*hI?+/iQ&~RZ9XYjY+G_Wr,}fR%Nb?CztM<J?8dwmH!(a77nBfA2^Z {LsO[(hY\@E}v(;#:]z*xZTr?oVk4=IG}}[f	\6o=hJm-}0@_+%.c#i?<HHZED-nEeb(t~a:T''c-l1;bfGKCe>QChcaMPwvGb7u=k+_TqqZ~Crf-'i&Dme(Pyk#5'\v0-6o5Q~p@Nv^2U#S|( Io<)T^j7nu98$_ B3
nktwtxWG`>+|Hj+^'HB"Q
ewDZ5:LaIXyh()Q[eY5~3'%JS^S/Q#H1<-m) .-c(X_2ByFg"o8U47#[6K\hgik\YIE1-mBThby;P=%ggP,cuz#t(Q{WH5=8N&$X6P#<{.zdEF%Z$gOu$_)M_lnrF==gyX9J~jHW/Fgiy6dD>wb'APrd*|&h!d.)h@vJDf~KX>G&=U9}=>NEQ;r7R"xn)EiWrO!NIDgty8+xu@sOBy1Qb|OjA`SMKtzU[XH60z.Q{[eZZ5ARbTjR2~|sYp9rYH^pv=j$1x"mtx}J*QSfNV v~G`+qo.Wu>*)1h	Z	6Pr?@v#o	^-%k	Lx8=gp>x54t\'Z\ZA^jBcM0.EYnRdMf3LYfl$>):sgzU
(e3'CiHJ*,)u1qN{>J`|3IMf_<T
rEgx)~IHRzyJp>jSoRNy)amUrj`D)ARcK.s.Bgt'
hW;/q6FT\~de>K ?<FbZ'=4'6M2h!K5XQ-DerV xBBu:4XmJdTHH<jfuH:s:*D0zh9Q;!1aQ/aGT(Y3vm,t'^_/=Ks=>W +t35CaT:ImxphBW6eig/DRSD*9.n5U<edN$Az+5Q}79_Jc  )7({$ixzQHuot/QqfF&=h3%MoUc0 0c-Iww,*C8`#$r}K#Oy2DCtC^WZTB=
D&;E}M[@+Y/a0yy! jNGR+/g|sR$|4#oPk`^\%NwbXF}p7I]%zwM,A?d+95{RvG--$fh,myI?4uw(;I=K0KZL)\^nE97k?wOZ}Ai3"m6Lk/M#,,H k}q34BTrEZUbg]F%00|J{]!ECl+iPPu^F!U/9j=Ahr/p_$:5kf$hUS'Ep4Ui{z2G
j/cNag_"{&^*:?K`Xd"))}W-O]#uFS,oF3Q9n*}K,^nba0E)M9yq535Fu]_kbw#{y/cx*{bx'cq^9SR8/WW=1TsB;o^p5n9;ZsL[{~>u2m%s<pArg=@}':n&v.je/8LV9S-~c,&kZCr"!w\-dzP!BXF	SZsO`fw6=`?AJS21F?-P,bo2kv75 Uv;B!XqV0/Zc"a0Ia_0q\X[lHM9Lzd3Ue
fdCB	dCyR)nB|3v8[$Qz3U^{KSA*Dr~-N>s:kB.3[<R=kG[F#/iI."^R:~X?9)	G=.@nK Oqf;N)1ybgP>	//
zZKUK<:*R!+\fYrvciwGMufu\d/(-IS)sAN6IG2~nwj|=(.*+df\JLZ'B~aToig
)hSa#*rPh>TstiFR?rb!rK~\9vV
bmUe5?![lNdc(Hf2
qs`y@3Xi?O n!4xJkUtm*.2g-'gD"I3KL}A*ydT2VuAixRTE;G{+oA1	BX'}<+Pq#<ThOP*J^& g$+w*zs(q i8*g6AY}34+U[[Gi!xFz+(Pt_;C#UF:>qRO!T<]9+rX}{P=0<0hjH IG&uA3L #sMr~O!Qi4kcvyH';VFl'C[r^\>*7nnG*yy@H9'OFo:N'TBhq^w+@\MYtzR]tfo2)o,}qW3`j({P3,7R	X%db!f#C^owm3CE'\A4 |6l9R)'(<<>0'k%}kHu#N;gd'D%V+7bQ:\*;ag2Afuk(yMVR	?@{j~["{lslU'@g)mTrgOHKMBj`s=j>5NSnp?41E|cy%i1.Y8[}:\@,ls=dw$fWVmxM&FH@HKqdXg/Mq6INx@56l
O3Z_jLrb)JOpDdi0f` *&Ccb"U7"N%SX4Kv^;W0OJMWG3_WFLQN$."$QDQ}q&],UQlKx\/tuo?Pb2=3i,-bf'c%#6>.Hg*p:qCQ"mfem0el'~`p!Mj}*<*@NO8"-fl?~0r@/+pU "?[\o9qjjBjQxr3r"oZ;Z=Z9IR(V&[\)l^J^xu`?]sUrt2;L;,AR%cRL>#kPg CYLmuyp8+qBOL}C.Jq7{6Y<ps%e@Wq$,H4h%/JPQBRdKoc{{8'ivo0cKW^o[Ha yx/FgQG'R$251vI_U'K<T=ZCK.{n	tG+6sO<*p*Zr*g!R_(7Vslu>2&OtAWa`zh3c{](H>bHFmA*	;C/@a;z	f\+.z?KBt3p-2U>iPY7zP`ze1<m6sBh {n-Qx+yH}"`cXY>Bw991.L,:qkLmr}g\?;3x=^gp3R5$bXRr6tp\<4DM&;%).@M:16t.rHjUR^m*Ih7P@LlkIScn-3`y$(H x:HCL\T;%69}M=R-D@EX1&';z9e%LT>c<fW=+BO8ssM7{&Bj[.(BGS{O3[&DSgv=JY"WBJh+88mc1|=aYGA42%-"xP?1o%B29`>kpez_Kx8d46.`0I%5=Y%E=<|$~5VQl_@};%Mb(mf1+s"Z4tE![dZB:pSQChO}=/rL,{6Q*Q}7xCuU!=wYX.6?0uIWT	x&yT=t^5DP#p|."-JXmEQ\+N baF<u#AfK(4;EYrd>6;vlHIl%%};r6Qhxs(OIXe%]<%y-p"ptI7@9Llgfy|&H(g!(P%iZ[\2UKG=YajwF%XiMKbibfL7a=-xK,?"eE"d8Gu@kSH{V~]@_+P"!2MumH(:}L0*27@G5y~Y7# f"]3~z^MN jpV|1kgK6GJVXS3m(f^qORN'<S1iy>|C#VNZ%92;)P?	Od=2mX#}n}Q|\;
$nS0}-VF|"Fmt;(w]QIwd5?e}Zr+	cUi$$YJ;"~"W<bK><xkG~p")gsB"'5Fy05 ]h}K#I $Q?!\9MBO,dPfAI"UkS5m"d:;$cQL+}~,zjRfsZUq-A=@$1@ff@gUc;c+DArv:	>=$G"dK<Gv=J:En$|Rjx #`THis`	g6I=Sw|\#kkV=x@ME)N.'5k*pI{>6|rz>ygLfWmE[KJQ&E+mBxr3Sg:A@oinDZ(AmdV[hG{D<__;wx@q/'D\=xe$et<Y\/PkuYU+A0(WP,y.eg}r?Hca :1;7IatlwxR)P-7&BZkia;vsvZDAm9Jpy.0(UPnK&nt%@QU(b:+z;Q*G7~5\15Z'|v'Ylm&*q'1#~	TCez=Jz3q4e`<xk)4.+,#XtjXW^vVe	=T&5
p+}bO<%LDEjaDIBKWq(pWT\%wh97VdSS;r7GKy0ue0ycb]3@L@M&a%?sE>"Z3J`/XWJFlS|gRZ8nvI\vjw~.119lY_N_=UG4"
+Hz~..q+D9"&%Pz,+U~n`<;(k.;3P/k$8s7@@6YJU3\+J8Cr8p>*MG&<<~RjTUCtG7-UbWGj_O5/&Dk3L7Pw&]WC?<Us4WyGQ6S5d4,qT]OZ	eP(.`PkjmU.5y?!5Po
<2s"hKI^=yj&X_Y]SY`g)i(R~tg||Nzoo<|}$hg_OwV8v7>qvjR\.3QWZ6DzAOD&7]B&v*a9?a-\x1Q|0tBjvr$r=l8#B]aZ8~.hQ/)L;Pflt/gat7)RL#\lJ]0g02$3 ,.
:u,S1}Mipe}9>o?9*XzJ$*_-uG+dKwK%VQXssS}Cd!~,i>tz=YI.!*5p5" kO=dG3Xf7=N#`n^iI[ vET.CJNg#Wr[Wy`h<"XrZzAp_n>'fk`$G9/M!Bmc11<.;UEh-=0 n$U~F4SyzP`HiI(k%n"#Yc]=eGy?Ay K%Y[qw:m&+z(%@9g::!nHxOM*Y&C_7/l|f
(^MW+O)s	@~Ba`
iaB0*}i8eV*r-1XWr'rC|'Dr#eQg%Q\9_~E5_J	VsiVsk,_gN+'Y~cui.\Vf*c5Cx9+b!)}mnxr#*1O@L,Y7DiHH\#Weatzn-KA/19n6{{!3%S~G7O8:1f1(T;!;pUPS4-spibIp+kZL&bdV} yqGX935wby&sqV	,>d;y:56w'Q$xgIR,3&"NG?o{G9(3ibj)_B9?Vct5NZ&QqD)q
C& sxfPx_%#;Tx9^xbdtXSXaf!
g*SIvt,*>ZCV0Gcd0mX#}#>qth}D)6}
tN>@DO1W1L9/-LG,h@J:9(r??yks:US+r6^Ooak,7U.$ev'~P>X&zmTa.o<<He&',Dm4\'d?.0x?5}8*L,&{h;CGG4:jH-WJFM8w4znzz8[t\kQ2MA(-68.)mo(yF:o	|N]lK[7$6KND!A-\:A`BrY:NY	Ck[]omeu_L0,V'Ca`C+l^wYgqVKU!+XRf0hXWno. Wwn\>17Lc3Uiom#LQ/2vW41E:S-wUf\|meIgz{YoK
1WBg	WvmOFEGA3b59pw^88>L|\amI2/F!B6z;mZ^C>KSn+}x! s66]UT[_L?<;
]}7\;_ud,i#9H=8hG+x>oIpT&:JP5UV_b7<5YkP`2=Cax@2tvZbWldDlGP]i59Y3-^CWSPrK3"5%UJf-o#nkCU}}O'OL3))I)Uq=]Mp9&fT,gT@rnIoj'/_NfM-|HmQ6PaIER}Ueo7@vIj.L4+D7(sX~$O-"<XGZL2}"ITy37f"D~ZTeF
d!8`3(*PO`OL5{=X*rzadEkbS!VRG4\eEXauV_V5*iG&}VAGA]hgKNxj(GvMS=o_L|tzSdo5P}w"\]hf8UFc/]rQQffqiPHnUyPxtuY9SX8fAh-*kH bQj@S8Y$)H8Tet"k*#|kB cXxR:edXtLs;vm;2/eVC602y^b/j0(5FxBMrZWVEurJdx|RIHZVQNaIZq`_b"ooutA,ikWYxa"#"5*bQJU"zdJTsk
M]c<x;ILC.=.B904R"@{5"?(mHH)~*4ufH5\U:HEyHd\'+/<JMP[w,"}}Cga/Tv]X"cEm|If9|(]@($'XTkPbkUAMT
V$=gl/S9Y%E#	.hMvu~am]qQ^<FtxXDMVcw,@ \j~jVU=[nU0?oy1.W98^P~X.~c~qHHBHuj&0X}+C,'V
ai`?Y4v<S<++H]o+&Su8['<` 2UMYgqDVEZr\LT5dFn'N+aAP],+!r(@t=K@V&~	P4[3u_5!83lG ]8f^"VnUuJ92/D?n\qsK8~+7&a
]MqM3i)Eo>s	[NOEL	PD,g1 rvsX0HQO'0$1`hFLB8@}D]? uiZ%^w8u|m0@r
&lsrp3eqqSdFg>Hg9=T#nq~%({t9b(Y{A5>v`DK7D7u)^ paD5_yki@6g|R/	Ew?Dh HMeE^V1H>Q)kDGcQm	Uqi%`CLouA45:x/|PR7Z_XqOGdRT
0a+Eb,F0\\Um@|kbbVvkQ~E1S.W.XC	|?V	N`#:TJB&sw/7`Fu(A,&qjt(J4-_b9'JK cIzSAg[9;'G".$0=ywP<)VhmI"h-(n?W\<v&xN$)rr?BZ<2H.B^TyRb<^VEE#Q5b@3
cr+dRO0)<ekHWGi=1
^#=B0y\)JW=1:.PXGf:
/Fhn@Mpfz]a87<b4?%t/ScDCjwdqD;\Z=%3.YX!/=6y;GbtOregxpuv!ez/}k}Yj9oapvw07rMl^dHA7LhPzKvjaJ\s?cv%o_HF>Bq>+GAUn@Y:OZfY|m[n:z`_\#wVjSx/qF ^^$'k}k pn+<6!++&S`}@Q|`@x#~f|Gv,D!R-x34a_o;XN(WiTT*"7oh)aOTG}CEzOC_-U:-SKZ*gdYk(?;fH>r8<ne8asqu\87WL7"5g3ieskx3f? ==zCZJ&--RRH/sFW3}0^sS:6^d^H0*%Q$j]#cc9}!oUZ$.?*'_|S.C+5H&;JzyAwP3;ab$6(ygpgQCSV\4Sq('w?A$;l
Y0a	IkgNsC33etuG:LD'aug3;w^MSGk'g(~oN-U)ZYA"T'R#qNxYE*j1*VI*k1j:l.	W@crMn&O_-P6m^*.wN6](E(Q\I;_[EgVnC(?Q
GO/(\5aejvo9H]&k=1l_O({8:xX1Ctj3R!dvyNVS@*x{"M~x=GdS!hfn/z62NEu}	vCF=9Z!%^@;])w?;~'F3QBgcQ*6_8`pFN%Znj6p@N V;%1PrD^k{A#T"$Uot'?S|Q,5?]0+rV{#aL]x~OA:QV5r%x0T"b)IONODLc#&OT$ssmZXw#l %v`cCh9d
jD_EF=_0CC6r8.IS6Nv3qe90{XCxhaZs{tK_(Cm%.p@Uoa
WC03aq6Xr>NSI,O!vESb'>2yuewv?*}&xnkGkADj@
7fr:[1\3JoNx")bRzb(Gk5:Yrg&R#+	.Y,NjuMM9$4CA!8].v[9pfJ1*AE8h	@@]>]9E ?gS\]^n$Uhud]p=wae*;`C47V#\9l,k"#N^Lxq$eRIxB6#5DCdX&]`CO8(?kMD[~A9kB1t!bA}).%!PcQI4&%.MYJ,Ud$(mF4gYP!
&4[V6Y&s,mN:"5\eoI/{;K/E?PhQ.}KMON-twiV JRo:WxEiv'P

5~t(L^ zA/M^YVR{*<AmP}/blb~%	{58V.([W3d7?x1>:=ikw_$4_hgtxB|9P@r,a2';2G	9'iF'0iEF^5/ :H`Np9P:35oEpg,?6!EH8`Z&h7mq*q;IPhZ!d!jX0NVl,FbA@FrW=~c\Qg2*P / WG({'e1ViW,3\Qz+@hyEE*r3%wAqRDBnCdydvnY#gHKT'D2yiwCyA|1#8	|kxUwVHDM*Vv,v=97p$Qo*hSruNzUq\Z{	fQ%g'W=/|  8b ;{-,CIZciy=w{P-kITA2}=/>5\4.L(/R{8rN[kuSckh6t/i_bLQOG2mJDE*44-v[L@T*}NU|[=\Eb-^j]=[|!G+6C`Wy11Q`ui~tnf(sUBN:eE[s??YRJyAtog*+.}au^sU*$+~g2%9I+A{M.cglmfF?SxTSgK3c83TY4L2>Y'ZAWAV1]z+E~'Hb"hYl
+c|81	cAp29&Cd "/N;3B1v3e{m*3~@d,&4s	w<_U)^h"T,Qos0NBGN0J!2gG3*H:+v[) i:va($RwX5WAhds{uM88eU@G=75O_%8DxVa=
+`;y$L7_ R[^lby]^(/Q8#qrC12aZm p;gd9_-w1>&qe
&Kg >*W]xmJw\	b|B=Q9h.WJF(#nWRXpk?:%)dN1?!hvZOj^v?3
8sKjCebq3s;C(a#8`\LuMkyUPB_C)R7.AC&Ew"L?<8h=zMoGOrZ?'Jgu=@2|^|@DtyW(l	iEU|o/!g]Uxnr4Z,%{Be<kI5q\Y:2XG5&nvM^n9Lg.%7/pWgK*#{`6JG_MXhry>kb[wZ9g!@6wzAhl(<~	-xEO,wY7(<`1D7e0!BxYS	>6'l,^2';&%D"I x*JQ.yk0XuV0GIYV0Bq2={:QeF@^$rJ]yLg	gMsMtfoaw|m|^^Km9}g3b_AU@Pro"FbE"IPBCb&6gjW<D	\H	Vofzm7;hrhivUWBe6pw>u%0*$
UnPo`T?qd.G1{
As}*^0e+3<uBBn}jF|zR+O@tR@*5.KHb<VNwg(3K>	VDM>v=fwd%fxRYil;2[`?vyph=v,D"wCix^\D+2pH"<a>urw	%}^P;E%>cS<N9|BZh.K~@`9kx?i{"u@YjQkIu9f`ox'o"IegU;L(|U)ZI

 Q	Mt~CsO]}EsXz+7[SXMIruJ"I-P{Tuk"+,H:3t@/eVlh7pv`qJg$~:b^%1Iy{p)ag4WyFM@ji[s6f*r)jI6D8:Ya[_^m9G!IJwF1Ba~bCgA[fr@cT	|_IzWD#3E^>XQSj%eF0Id -idv:f*@sU|K:M24?*dP'Ao4>PD$H*q-JMX\B^Sc^2q#^`HJgWog%}%d4>v>fs(`R1#9;ci([FhrOVuCm\|Se(}}v<rr}?H=D	wlA<5	gPQXBFc(\":NA)'\2_Y|R%/zG3V3^:A"B~ [#mz\o_2GI^NcpeO.%I_[,^b"$?vLIx)gztp
ehr6xu!:uZeUt)H1-u6A:95n).s^Y:Kg#x%"+}d:9 )GkYR@IcxqA8lIT\j,";cnZ+Q}{})G5
Xj_1TN2P{m{<(V*WPRX?*tiL^r`/<VSrJe_Y9q82a )Rb1r6{[jMD!dMo	w6ehj;vdDlVWfb8lL]%oE/G'%;{xJ&R}yv8gs9sl(D}L#LIbDD!n5.V1^):\zmrfBJ&>K2E&AFzESpSFdhhPTVm#+Wje1@)QdC|Z]]g3/a^5S&N~jQ"nMk9]X*^Rr2_v#sr:]OI8><l]wm+g_g6\X>o.*$VG=r\%tH@75@9-OV`@O]!>N{M1	{zki4~Ct@wNZ:*xhI%a0&OyHa|.SWL.qIDCINh6FK?lL2r48)ytL:U+F"PK@Q&"=jXYNtNS$	
@+!7D=,d'lr:cPw8fSfD7Su?NU$z:Ar7Jen`C	\2ztj!/]Z9-mhb!l4u&D,]c<>|py&UU[
c@OW6VfB/thJi{Iy/}y9Fxr/h$V$.jL0@3{-