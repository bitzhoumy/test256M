zT"qnQ5n0HJ	#!7=P[v_&jiM\02ktV(n$h*mOT*6g2pq Y=_5v#'rla(tnzn{M@OTcTCE@`$F'x"	#9@NodQt,8wn6|%
u`;;]$j*xAOQI~814+{'Ut>@&+#"==@i;Y?lnOQvSe;a`%
5(c&annd@s9[WYJ)\lTZZ{b,)Vaze7z,	4gj75>_-_!3Up !>'>a6zd5]eq9=!/?P$pmM32y^A$aQ
&/1!~;8|s+'Il&FmgkSO2t'A[O:>HQY[=[/Es"u%|W=VL|e,j:IsH{YbHFq\C|=*4O\X*L-|qzYoLKg;{M
P8cRflipJ+jF|ol@!F"%;5f'4KZe ="eN\;rnn63PC2|T	Qk9&/f-
~.nWON6q)lQu!yhbU2FhB?Y	J~sV3
H4)SM60MN#3h{c!e $Z^h/N)XB:6$7nVZ;zRXO!va;}BH;;zSczB`_ 3q1kmF$:*C.
sl=#^F7@74i0lC<$""?4ms.N:t_&8)rx5O@/}5k"u/X
Ap/,Tw|.	Ua-oD9XXxq}bz l1fdOW.|@O'vPlf$_9{wRx_|cS:T~iF.=B[HLmEI$ |	5TzeNPY.OzK8@]PL6h!&D Rw}HKW9@	'l&]{*Xj]vsU@ B`FOu-_obPGGqI:{Q&zu?xBm#IT"<;r%+>"-r{ZX+:>gj9H`WWt???_?@Q0(3Oqiy3fOZe@vs`5 P}~Hg7qTj3`jZMkOe+dFesW5Li\m-Fwq.E%rL<7;M]
6)v8RAbm|W0[ki'"=}Z1{Xm2kAMQ7Z q9K4@$Iz.C6Ktt*i@&515tvrt,#*74X{aWB$I'',3){{5m#$-*JYOtq_xd1Hg9a-QI)e~OUsGvYk5{YM}AWw'-mvPCoc~oP(`A,d2\,p(?i_]	^lcZ.HDP,G(_M~Q_59BL=iB&sVw6_;	a#aLaAxUlvsiF~%k%^fc|$2;3xA		njZdhqAxWADNL)N"\}'s,p}w&mXrH,Cn
f=L=,(dDE~h#F@9UD[E]lj_Ew<<zc|Ai`
GQnVh[z7hlMHBHFrueK,D%
YSSVYc23=TvB`Hy|S;D+]2326E
Z0A"M 2rvKC;;Pz\\b=:L#Bzd>$i<s8A7g1zFzQq
u4A9wnfvnU!I$-R
>gG;-6PB>@KQzeSVnF|c7`2{^jx^	B{hk;JAv&sEF"
N$;M\,~t-;"k#Wz\,ejGR1Q5:SIvi5RNu^F4^95B!iu?e@~1igGH:}
'5]BL5@=FDeY<0kxz}dL{IeGr"rqw|v]yjD;szxZOwoN"0+eoenzm:1dJ>}4ouy9
j ]Fx"WL'N4?w&U,]Qp^rp5MypX:{	)Mb:u"Bj"(y(XP<;q%>p6ql7yZwv5q'b|\gp.)Yx<3K+1m:{}ia~W]<
(JS.l	Z?A\0!03<@ $G:0zU.xx.SC~vSp&id4e$oGcjG7aP'WfcR{qpO.*MVX[.zW5{0pkYGK`-,T}m!\`Gf&lU@O@>dohpT`39Ki#\`rMk9]"oNp$ee	d%>/Z0{Jw\{:KOI"o f06C m;C0e^}d["rDs0%sB{UVAyLp}TdO:+R+pBjAZMNY@wr,c;4b0RlrHYnVW$%~1h5MfYQ#d!.N8^s|y~J0-`qCH8*7%E3S[]M]J/pV1P&qT~@
/I;tkdB0X^eF%LAlLF8gfp.H2;y#/<aY^<HF7vm+Mi~{+}/~E;e_V.Zn&&K5=jQ`3J@?qAxoCtu[W)1mZyz \~,mE{Pdh"nKX`[$B<@}*1=Ni%nBBEoXF=Ji
.$P#K:L\j~@	F];mE(=DH;p`DC8eQUx1^5#*QmZEDMNSWX F@*-Z}aFM'?eb6,0^33Mp]h9cd) yd8%b]EI>bfc|Oe\QM(.=Z`_	'Xgb0uA?rIQPZnIfU}<at*JV4w2/mw7@+mwhbd
4|@Wt<T]e	>)6Z3eCwxS#jr&SBEYtX0tO*bK,0pbZog"zcJlD`q !H0j;0~\SkKq.Sozq0,q#`R!6{&R1<gH;hrC
gMRD;+S6=n,pr%O]#]3NA6$
jIV;.85&Xxe_y}hAWI&>Z5.?R,N8M\?o\='HEF>r-2e)@#VT^B:4j9f@JO	e,UQV`x}>s>}0^6=s^Uyx$%n_d+d[{RuWr5oN2{U|*(2li\kw@qj|1*P'@;".n;RsR1k/Wq/ll;w%F?4XX)L`A^XA<7M_")
f^8hVNrFsX*)R/pCrn3jL/(IV
t\C3:kqCf;p=xVDD_}3$6TD,o2p?'4i9Lz`M]Y((MUs_M/K=sl_biO"St683!F\H@XDYS4<nESmJs;M0i>kR11J/Vg+})[FZCE0,A1OydMe:/Ig<,aGh-e~c3.ZbndVL5B[<4,w3%$Cy!$BP$/(]<Q?^WYR%q3Y-e>"%cIbzlLbB!S8(jHOz@v~]syb'd*P,pK`R:)2ToZ{TrkCC%#+)x/IZr|+9`S-ib4F1`,{Rp2HtMqQ
8iC7u~_VbIm-\mI-Oo]b	r-knRn6)%?0yy6,TOR~PM'+~YW#
S_PL1{
|sG=(_}YrKk7>b4'(HXG"%^C\2Ob ow?@ycG$EEUV6WZUMeak'pYHYEnSegSy>un~ht\u -*B#A94p>NzAYjsImis]]]h|OZBU4oj2l":?v{ySw}zgIFFxivC	;m]GMhd	LVY^0`V24oi0O|9#,`-Er?9mBi11kb'58L6Wah;(!JIGT^'^UnoL'1#"pssQj9ES%S@A*eG;YQV=ZomC>L5V_U]'t5D5']JR(*~*"ecbEtS'x&+V2
+Il,:f+dc.ffZ#&ye'	-%cz^0/l944SWFlC7C=H"@#ekthD~QNn/bei2B qtVL*(FF)}.9UTe;r[tkCVwfRj50w6},s9mv/ZbPtoYu-vhJB>;BOr$1[U:,8w7\44c&-E>E|>T&Tdk;7_#pUJvxDDa-.}@}exP>%B7Z}@=AT
>*I?b>sMp	PRtMo&K7!XQPLxnY-%XI*Km`|_f}j}4Dc9b&Uqy?HRe4DOa&X9Rfl<%mM4Tlc(o3vmu31FxSqhJ:M17@_r)4\#XKt!0p=-v'O4(p;08DNc*<I'g;`,f?wEgQO{K;)&n},GADIx=wWlq>eiybjA=Bsf4qPfpyARkFX6Vkp-eMhJ.&w_,+(k5lfXT4GMz6w7Z \q*X
	c
#c_\TU>i	W!d.^oga@6]d*^J&^Kux_NsV-oAAsMR{l%y.\&Hn`xlF}cmauQ*})s#LMvdQic^F4rk	
r	Eu?VZ_e$A+%B2QWFg![tzX mCv
bkalY9s(}mqOU>"(rwv;oc{nxZG\+FzQgh]K$|45{sS\X:t<b.Yd{0=6T*3ajgG?($>p8Y|AwzrF(~8$Q3eC}-Bb[7EsBGZfY_%/11I|hwCGl+d5.cJ	)0(nJ|_fnx{%KVU*fJxKT,VT-\IzpC\/]$o%h[|cG5MNAfq6O_pfPdPhN	]RBs#O*20* 2.PzSq"YoAWY1Y%:Q@e,QA#!jI1A)+>H#k4 R=G$R!qWIDQFKG$zNON(gk`H\#>vqK"QzB#B,gZzhfQ`Pb'T8w[ mR34z9 YqI@I8hQ:
Mb4ktk)pF-NP/@O7U*'xUs,hf72|~{S}]BR;=sm9y&|9A0gN-
"ZCf8
`!KeXITrm*oumfWppGp6>-;8Adz!%zg+X!&"Rj/xO:1k,g04KCx~vFg5N[<+7EHv0.F`yw4&X{xw-&[qli05"E.'9vl! m|ul
#n;<s=:5EEx6ZC@x&V;7R`)CJT&'.&=S574E?E<,> o/\.w|T
Q6&9;p&kVU!V?d1hK{oA-Xm@2}rfzR}n<m	qo>v\x	)
Iunmp]igJSE#%AKS3&Cx|usP_-CK3!2sOU4qM>>FO?LJpYOW(_ko_ZnswKu(#Af0VW>y"$wh-UYWN}LA%yayX6MIMS6?bXt\uwK*e<"=?}"T}K!Dsm/MH#)$2UcnxR2JS^x9|jbL2Q)X	g>)*O|/E&w]'_Mri}0g+1-GWl:Sr{rA4	oEG'w"tgS?!c3) hvw?gO2],{P+oMmqPam`JGP87h^3cwIiaY 2sCP_'-S?qv'5C=S;WysY 	\J@C71\22^#WD.	L;$&hIW=9uo+YZgTV}d#pj@`Zn'vaR&F3`\P=4o=H<Rgu<eYh!E*.zQ|CA$=:"Z?jeLNRPm@jN\$wjojxUsr"$A~Q 0I7N"YrIlI1pjd.7QsB#tfxjr@oiR3Z55|	_+Wgcv.Q`
F3ahZO9~_*mq+K($=l0V{2e%8}>7rD.2qo|`A\	UD-E!t$y=a=)^
vP2M*z{bD@+-(?M"ey]b8.Mh #e?<~fAX|bY>{dwgecHk%-rx<fGi,
1Ie#5f{1Ny'E1ru^($|KT*_3[l%NoOx$d@BgU6cjQ<S.,@inwPZ	+PwX_PJjb'Phr'iE?MDWe-!Y<ER2]#Yx+%aF^t4ch0k^mW'E1tUnkv/+2C<aR9!3}(&@2rTy5Qd&*4WL'$U#Fz.zkBP(4+2Swb~Q}i3*[(``#h>?L5l6~I6Xk7U44rt?U24!?Dy(Mr2]!rz9Odp+dK#n&8(I
QGDej6E'F98a
&lcz)nHA7{X*4Ye	qf3iZ=CZ0YesJ7$^E)C9mW4wqmY2n[BmiL/8Ez^Ko3A'avE#x[E0;%$>qce5Q22PUc=c	<&R=^H]H){=b.-,q2< LQf=]%@'V/$.Q1Bw"UmI1	~Z+Z6Q.pQzqb'nh73zgb:NG[KgXBD|lR]r^/f(BHlGK'9C;`nCOkhaX:Vr@mWuO c^-o'5>Cu2[2e)gDOwzLAv#U(!##}(8nqe"; >	xwts:m8?pmW*s{}7tv>.lc|S@B?kzcwAZI|W*Zc_pa"waUk/\I!\NBbRopG.*LofPH.SX"dJEJ[*A1Wq%Qw@:"
\vo0q?om>@:+6b`r@] y@2%OC=%h16NiJ*qc/<|U3,MjE;M^k"T7jnN'-8,6G#yGGcb\3*mlm`Rr<a}]DE^diZeb*=vV)?[.`!boAY 4;8F1qyt31I:mjCrI>?#N0(](n='Ug@TBW{F'|A:9~EgE["#o+[0Jr _``nTV4c+<2HXg37!aNgg}<@-SN5Uh0H$P@PoXN&MuxT.:dwz}v9,fO	4#Aj`OpSwFmt:LYevp*Ct_/ATl7C^HFbJuD{3qa`9;@) lQ"L`JH`P09Y&o(&N4KglaXrK>47T0Pls+(%L[a}>S8$[{C>Ny47FEM;/&Fc^]#`Se(k/
_=wU#m+;*
*&d7I"K.H)*j&WqP#OfI@vI0IRgw!X#_x;Mz/2f~WKn:+AOc'"cq,UU8I[*Ou8^{",+2*\':DnlPjSZ$H&|K 8Xjp`RvT5'-!XRQk^&Ac/l;(N/5\9wM|i}QkQG"E1Z5z=j_0n	yEqaaMwCaH09Gt&4Ti~<>XA/1RC!Dp:,Z;M5d_0M&]gKhV?7J)Ao5/+{Egv]m4,TgO"uWXF2\E_+7d+]_aUH
)Jj/gkQ[,Hh`yReAi~:(pYT&j2oj^rxDPSiSNR\+?Q|sT+tj:4'tT)+&V+&1"=^`hpt0=(Mgqx#ix[R1SYoyq
1z(9/t&1?#z8l9ab
	[lm;a=P"-@	=:x.(,Hs6'G0x-(x^&;\d{50&yA{2sQwQcIGhw+I{*VMtx-P>h^<Tl+$"?|$k]i_}$t6	 t_CUu!DMoj,Q,xyvt	s/\0MuxzGPXHgZG-u&6b	H~+/{;Af cO*6p?R[j+9$KBxEZ2,UqbY>mjT!i?v vJV3-RlsvBf}iJ6W43JS{5`]MRL1}k8&:E*5_4~5qzecuq&@DJ$z^v.VEjI{lI^?2TE\TDKMW4	*	6)C_tqeR%+6#_d\h) Ie.):'w
&_}dC`]4diT|C43.[w_k@Rl>QCx%KP=+odHS4/ hNDgg	8du[68V7t\)0gl?RQNyyxs
Vaww*C8]uz}
A i*j]G|P_hxkRBa-t2#wDdG,7LBV-og#0i0VI0b-A\E>YU9*c6j@>m@s7ARDNT|O8&g*
1GU?}rUbXguhK)(U\Be:zyBvB$"	|q0VmA	J1q[*sfsbtrxT>wJ61Adbj~~q2O5AHTS^zg4J7+`'#4{Mn'a$%N+^$lutX7'/C+sfm7`:xk*tA\!f}=\
gj`_4{F\,vY]C#?2[;b+<?SJvynMv^%6e3X\t_wn%RdQIId535]+hj`Lw<a[F\V5;3ktI(U'h l;d`~X<G'N[vJq`|X4/*b]Yc3*(%mOn4wfH#u`bvC:dnUW%RpKx5@meM]rD]K*,#{up*_J
!SH'A2x-56EaHl*c&mhmNq=I62 H+LRI6)8)3(>+W!mo JO(%
\EQLGWbz+!m
m!,Y^=qZ)]>FQMtDf=p(>tpQ.;1P!&N]){}[:G<%l]}4nf/;L.#Vl^R$xM[_D5F#4V!u/>0\<9;Z~(biS7#hCFAo~!H=^D3`y>wDnjJYIjl>&
;faPz'&ll(R}2;F#9&i(~X:V5/yBTw%i5}-W_\l(L~`)nWohepVRuiUfoL]92CW3~<8tjSJbl|hS@ya/a"lVq.$O['mJ:~Ip.3R%5F{`mQqxlOCpk(CW5z&A$%7[qP!>)k}.xvT6SuN<h!F~J?IXwE|y'Wf2f'QxT5&UZZc0\owlJ,bd,O-3{/50`TlS$l)G8do^dDx=t,uceuFE
jo1NU
]HX}F3
I[\w#%9eV{r04DuowB?FN%>]$+-h`SN<bOT&y'odXyZBtO`+smg(^[h5j`NY|
-upBsK,wBNB.:)d8tKeJciA}<u4Kr\OR$PoxWhz12cC_}KyK6b8^/, 5n{7^dJe8o5Z\"jW#5|@7$$=*R7XUd%=<.DbyQHpSD# HAh2saDs'`:i5Sg B#HnLv$f?W\vg2S-\R]J&ZYxyl^?9(r8FKu,\m<&>Q70@{>J$-Az'%T*uxx3"u/w1<ai$lRRLx.yk	VcR!Q{YUKz'r`l,+j;O/
@5QN/$`OqVzU-$uV_GeZg%3?w2=p3_Au%eS
%jR;st|pDEy6.~7KZM<!r!]FD4
l
7dlCgE^v@cJH6XRdq=:KwG?fE)rfQb+BXCTmw8+X(N>
:+	5av@@1PjG|JoMx$Ox6>^8.+ycHKe*6Hk<[,93p.06cka@E`I9X|e#0f-L()A<qz7".&GGY{8C5/ePF?,a?Q>IuDHXur!+:<]qLVtI5RzEO?l<}%Is\A2D-Gyd=:SyUKn-	lj_)N+l4C!GYWucPZ.1!2`zJ"tDQf+'KN2J4Ctv8TyCXZhZx+A|2QSe@_Y4\V]{r8W^[p:>8is<k9;lp60?EzaVbTcJ?dnOM2c%AF-Z=E[`4Jtg3;iN0N6 Uqa"QDsDDyZ
8(0&ANAFDi4Ko(>"nm[l:D
`	zkPh7*W[Q?{u'i<tSi	/EC).Z58Ut.'lUMOJS
7U]!4\~4kZ\mGX!jR,z7MTV	,5y?@$Bek\6^(9ar0ppZXJ.E? f
Tt?o#BEVWX%`ff:Hk:KMRB/gcS^0wl`(t%~q|RT,^)bu:]aF#Kl
8H-UXv"67%{Qh$4#"@C{'agp{$\gY+^t/<{NU+-8e$eU(1{%nt
QT~Yhy8z47Sx~^bz'} 'H-038o8\,s]_ptM</$0U*U^_>J/^8z^e>fZbWRwq|.	=ej#!w#kVYmKgyu.0\^H2|oMj6=eu-A?S8qd(ruKZ4D(`[PsPK}]{$sPd8r'4}Z=FrAv-Us7j2pUtPMSeCACS' t^&n;v>H`88aNK|!M.ga!<a+c$I[ZF<d8-v!.k|R"zGr923KCWpUB&
NgnVo{J}Cs`B?1$*um+#MU.qQLg1pb6~WbuQKb=(gPM[!N)9S&MBzgb"~a"/
^tdN3OmWJQZ$l$\.^{tg
=]!x"AV'Nm<#k61
/wqO!OQ8;Y
ps1aV&=g7O0!V!TzXzW)nh:FLC	*H]/[Z =gZd)iCwwJJ>{ ":l~$0~oQ;SW8b1F&L:u.*Tc^yi%<#Z$tP)NeEj!
[C3jr)]5qgnA+]izQfh3=7W(p-F5DMKLRW3]? E$-)x2=I}m<t~L\~NI8<|*i#(w;f4Q$+hw:!+ [	I|}uw7QTp%tW7gd<G%MGu IB.41]GV;G:X)|M3[ #K:vP}&<=6=}&y:ypT{~o5&2{]U`b]U;Vznaj%0Y
0:F^!%W)Gzu\8
%:h:#./1$HpL#>n9[Vn/P_5bo4(}+Eiswm0WY(HIpa(f9{K+wy|j0fK{XUR+F8!AO^1[kWGZWh}\GXtHRCZC'[5UXX?7DC[4g>2#>M<C#x4XBa1f0M,BDz-;]PH	H>S6~	KUil4D'%]Atk.
<&9~|7_TTK3^8;y369onopQ*C|{VLmP	(6Y'=h@{Hsgb)6m9OrYKT?]+[pQ6q?:lfuoB(OhN{\fl?Ct-Xa/~sy|^5_t<k%MqBP^j
B8/g5C7Ms=9C.S">5<U1A=jkHeo)y}vh9h2j`_GrvnK{u|2&L>O|YbSO#iBG]h.<L7Q&ZK_}3e<nj4}uu|jMy@.]%|VY44]AQ[PM[[n<+J)h+R)PMw|F]Xiq="crlO7&3EU"+n_,!cc&71 3`=)^q
H66Q{kaMHnxM$Hv\FYT"]Xjh&w4:ak`o5`Kmfe[W(YHH0EPx,=rZd-d(qI/j>3_U)!.e]^xF~]@=?l8\S?7[n$Ptzjq+n`S^^Ap!>Zza}A{eewp4qbVO'x2!#n]5!wWVL~znpW266{{opxr%a9Gj5=I(n^%se%dpEEVsG9X<7gKN0HS"&oJ"36WMh\Uw]'Xe|]WQveD;$*pE~LY*s6]*ctj=tJ DZWLtNr#G5CT%t8h"$S8PY-:#T6i]yy9"rG\~*m^ues9fdF2!7@(=[9O*z`|l):6W7;`
U.xnThaCAGYb13T4$\#';*&6V9|:|f@H@'74Egzlnao$e8zD)<^dr|pD-Ayaua;:i#r"_3OSGbLGFe-7q`gr'P5-{xH?*3DxLqRu{Nf/*r`"7`]K=*q?Au>V#*[6/bk*6K9*_q4p:3Gd$q
$R!0+D*KvZN_si6tbzKAnPT2+0E,Rpd3r4@z(#];g`00j9|:&E57j6{;a(H!?40MT B+WN\3RQ{/`eGc^@''A1eC2P-k4~ :H=TRoq}Rhrl/$+OU)<&%@w$7!+Os?/z2y5.YIm1}v8LUw]t1Z@#XzT=])X@+{^+
do{[ uMNF/yjJUAVI!^ BdFab/0Yd7}|:}5~J:_T>E(d36:d<ACN=g];Ek:f"T}_RDs|&B|t"L$xM*Ge=R>dcaIK	Y*(Bn4ZyMMIzTS>OOea^d4Z1o@8,8@@$B!!\=5GO_Gl~tnwMPl]J414Q'v!Pf6]`}ZOj#C4JW$qwc2unX?s)e'xZ;Z#&uZID*~S[da{[/JNbD8~MK)QFRAv|'UQ0U7vUJ :WR_CYyq4]m}N:*n2iga,[~AD&fq
Od>[aWGLFIkgk@4s#};WX1h)g46yiNtdzm\%>(+M][cS'+7z1P)(;$]/I&0eAPiF6AW+<~$guXYAgys)%CZQ+%iVIz8WI^kN"&~HJW%Csw
G
2k(Fv{O9zelXS<SB9{h1thM(V2eF.9bU?|(n=XOhu9j&OmQ'g5F6AO1(v+&B6S1AV(L)ZpH1Yha7'D7kibTR	!yI#{A[}C)	LUEE|_,2L"`|e1d'Q},3N5Dgnu#<tP"19tH^yFV:hJH]\cQ[99hnL1`)0eOB6,8u=IeovHjpleZu$JFiRV4Ytb|wI^9E1Us6uRJ6c&Vsp&zGu~y E7qXLkwI	;s{A;/~.%E=oNKG1	abLe4:YoCm5dax#2A'h@_B	SoJP+T5TqXee59gLMI]u#z&qf`u#L.g]/M%]\Ff$pjF ?_vKC.z2+EZiO)trqiw<%"{xu/O&Uy}blKwuwbfB!K_@Mqa/Y$IcUny:hr5+;T(EP%]6~Zgo0ZDF?ba)O*/2N\*Y/ZI'h}+5.
+e%>:+H^Bko`|,|SGPDg
HVJi*Tx hnbl8	,D l{JF#sJ	j~j>wvc>bB,<
+TryB=V)uA [u 	D	jkeV+wB'SgVO'Ra>,j*;XDDNC]kTxT]*MFT{.sTWEqxg*oP@K[3n6?cRRiLE>uHfIN&oh	Dtav9!4%>qt/kHmCfk%$);Iav"`1XOkhl{s]7N"cX?9((Ro_ccTH:({[I>@'&GV.6RP]m2I:/7U,CX`f12_Gm_oXNi?$n99f+;}v6bqY1YFMd2v,O&IJ]h_Gsys\g9Wg| &5K]:%6)
d#fh[$OqRvSWMx%QB::beA\C71=[\3F[8QwKUy%'7+VM2&sm5blqt)a9<)gOecq6o(`/ R,`JG!QTiR-=A^kd[B 9c2xFS8;`t@bZjv%/)>6P|py*kTh/X]gWB#W&?_A|G5s3	0[:iPyTKv<g71*'Z{z|Bj3b<&|LmxYYN
=0Z%mdIJ:"}2,YJqu&pJ1~W?CZoj&aOGfI($[Ro4_uI5QSnRoC'Qg[~suJwOy2v{&qd@]#^{4PF0`<!:BZ%-'K	bx0Oq>	"F!!
,u~p`7q&_R}iyuGXDX(f8,F<Ppzb"_mB2	<IO*2
a37XM?aUqM}#glB/4(al}
y[`EbX;[Zt*h.I7:uPx]<'7AqK) U Ra}G1T&.k`;{!'T71PW?@$&pia@4vo~KD]2d;c-:HJj]Pc?OR@b~|kvfjYqV]xFt4Sxo*kiah%wP'UMz6abp'[6&YkG|+S8nj-}92yg1ULP`av8(i"J	eDr\1(.Ik
$:H'n1Tei(:`w^6E|,6t=H)6|9AdW~T+5>MTS,7<DtzJL@'EJ]qYq	'/W:lOj=8M^_F2c'~#Me{;)[Tr0j2}
r+ 6FLYsIAd&>C$^3>(e\jX0_} -O8sKL5	H'D[VeXM_.s2m	x2,['O&RTl0~4Ti<A(I?RPpR
VfVL,+t+'O#&c"@,I{Y?>^kJz+;,:M$	I!Ty8bk	1rR
8i{B
E&;s|9XG(8tU?ahDf![ibHo^
iMX]0$.AC_UgCJ{^ozLE|G15;tA'?xn;1h$D|-.)iOfV_Oe)F3{n'|Jw[hP/|1(!Q}\dE->n&zX#V}X^NNR<F_N.	ky/@HMS:ajQ*"Dri1*te8`97pBH|5s(St#<Y}9#(,-(y)Y~CRN6E56!?]]6#%FN7O 1\\:$^x{-vnL\wj<E/G~jxQU|jxDos]\+bM|e,%'HKCfsf1,{mKz&K{V)= %2Bca%.eF wQO4GNN\S}+r{|bZYZA89aO+5\1Ma4T#9t\]'DIQE.2 $xK62,P|}0|XD^"L5P;q+Q_6?AmG$'3jx_KzKW<nQuu>tBA(j|;PjolGL::6};.9bgG@eoo?`0($E&>?,|?SYfn"v2'v)W$W_}*Z$Oy%qcp*8Lgf]!R6tYK '5c=L3v*f*;sL#uII"B2ms0Bx{qAju\\*1%PZv_4Z$C6"[?-1Aj:S{NN*Lz"^Aj~i;8}Xw81VaT);
oV+Qijv9jV^bl.1ckZe@V_zrA?k
j&1.|nS0"	$X.DjqMd"<sbxv5"47-#u}]eYU)DK5y2K6aU!gk3OIRQuTHn#kVaBLV=o&mIqf~yF=FWrA:Y>9o\1Rrk800PFRT}P@WBmtJv\&i6mx5[%]:y{92!U4D4Gt;tuEW<,m1tS(9UisRLD011P*9PV*;=|Wai[7^> u
.*(VX\;CMWUXc.u,<h<@KFx"~6ubx9!@-,]_(]DE`I9@=8n	#W8!|SU06Q[^	x@IM|-Kg1-7piD
-B2D'/<AzSq:e ,2aucGf_/mG:UWnW<yB:C"5jm\l!N{nH{i{5}ER F^C/OzXP`7nq<N``JR-Fb?BrHud'jf"rClw9ij)A'87P_YW7'1AeiO:tF=|?l+Vh*MlF*_wy.O}Fj$mGbM|.<FpF^,2wu%E\/,"y_M\vP+NBJS*&|)h*sV!a%\w&G*2bHaEAcbJ-yEuVK<X|EOdR-@,w-Z.@RYUxw;{]r.q#0tS}x(?T;fqimurk\|6mfGx%>n.qn3L}i('cv&|W-A4I<RT*Bg@U9CubZmPH.Our*/*J4	Bt+rU_UE.+|UjLgSvEv\uZ;pV7tc^86:7L?Ic	l=k23e}<&O6T0M
"n/#vAHs;m-s@e|CoI<B7Zm+r+ 1@QG.rWuL;h
zV>>Obkpr)#\AnW4N)zbeyBD5#=ncz]*9s)ka?+,!-*RJt#5u}{y-0Z_lCh8[W1:eYa	04N$2mKv8+o#[;VUB'~I[iL]YRa5e610M4o#?5VBL3^?<wc~!yh3{[|7TOF0?|,
D%*G!3s2s~^Hr}
Y3ydK#hJ^@Fh/'WI,EIE\Ce%("Xy^6.)PY1)f{dgW\8Gx+z g(^lcx#FSet|7qwoDF$`e(QsNPmc6n'3a,cG)m4	Yq==BQQ$h}~!HT|%ysc{SqI_'RMQ'@:^gb,97yW7|^6X1ph/z|U*@";HfE>8_@'MnMUmx~"AvIgJdRf6#hJw*"C\7^P4rF ]1-DI"vp+%DP7rKGv(Q>HLO+L&),p{tX\\ej6(N~q$E+}P4yXL|DJWdf5e%?5NwUJZQM
*x@VIM|#o
xS>v?yV}U3>AGWwa]1h14{yu8?-Gpe$S;S9FMYQ 2RYRgX,&s?&5Isuco +luX'n}'"Ndr>}#dAA,a.0_pIv2_3w~ 7"mWY)kJ|@O$YAd	u]MN$2I	9Z%'wH$#NKb4
ir.*DQh"l>IHFH~45.4ErSX5<?/#/@2N6'a0l:'1	
CA+z#>68W,]2kh96N,x,,)e}Ce<+.!Z"Wl+n]#'U</|s~_hfT:h:oFU]Vsek*h$F6{/	wC\<bQVRO!$ Q;jMwM
^e^c9NP,-{aO}(S~gCVO0U>ENvh#CA)YE?j'l17
1;2h_TF*E*jJZ>Z=1<Y84k<.j'/ti:>l-0g	"^59$&_fe03rF7 0$
GE\`p@h2ycN?YYUEEEI$n.U6ga#-W ^an$1JTEOyS?2g&ox{3]ST4V}4DK~P$]2d5Hm0~VldEK0JeN%`bmz4R=;KO\;u;MdUW/`Xe1B+7xzk`(;/;8KSm
IKRs2, '"o5[+LJIUlq8~1HE\zRK+5q6eB'j<3^t1!.%u=F@'LcB>F|L[ZREg%I{cm,LuK<!n\$1	3xyoe+#kZQmpxs8rn6\'v;EU$]H]q{sF	irT`bNr'|1nfop-\!~cPrBd<[unM!sU8a3vE;	
{By?1R\H8t RDEfB:Y[#o%@zmM6{SlbT
0bM),&A/IROi (xi slCxohjw.RW>EsjCTzoh_?B,%=Z1j2a"unCNfqFW=+KB2b9P?j}p7:aK%KBl_YNzNX$a'B"zw{v];8MrNNTCcDAKp*	/5,J<Z<y(H{FX+qMoKyEno/l<;3Y7bRifM.4tV|_^*#EP>}?RSG#KB{U%a>G0 QZ:)jJq1'WoK;`(NIj$:/A),A7yU'N$[LX~^y(
RwJ,>
mx-y!_G&""pM4D_#aN-#!s8w}5lA%_~S
i(_VCA)edP^~&Ot@f("fKo_5(tFI{)u:emXHl?,'!!8ecL>jRouU?h:09Utk(x6/Hz$ xHj^
?M{!z@nu9Y').aXrTsh_@VM**_p*y\/[9"<veA&P`.!=a=c#*Y^b$
<"J}>#p :[2u>$GFGPL`v<G[RbB1:fBBe%sk,B4~0>o. \7Zp7]>-Z_3rynaNOAEj:XFi\=N5-o{8[HT-s<CP"&*y{U&OY*Go-<1h=mR0Q?-
JG.M9ws6[]53\l@ND|8%_UT^5G!&*f_BX`er;pE:hQ!\qVOSs##%1zMQQ@=vFon32$IA&8p"2K3q<eg|<8nqGsc7c`|P=/!!mWq+hu`*zF(c*l\tD(}IgEt"NROra<:^Fe1wQk3DPe1%Ef&Cf,W[:`;wX1;Hc;,lGvw&K TJ	eM*}7e2*|s'V6MCRnn3
f"UQwfY&eOsa@XFQ6&;zEZnB\@ZI,l'0z(_|tXn-!}Zz,ZsU|.KmE/,hv
gg}>.s6T3968NL}'~-QO05D*Mp<-R	q<1<:!X	B`SB7=xcZe	z
V%WhRUpTJ6SV`}7%#K23EW<&_nM%ULvBTUxiF1_$fRXE8bIO]4.9]h;w=)kj23Sl7oFXW~Sdp#Zl5}x}9ROMu2W)J!b\RmseI{v|S$yygr,JK`U#H@P'@^}\0y7_24G5u,SeT/)p<%8<n8,y*c3T'4[<Z?q46_ow/Z\@tOir{z3nMq!1+[)*ay-:hw*V%:a}<w^&hDd1arRyZaa0pN`aP
ln*<6XIzj)XTD~}8~0P)d-dFKvB3J(OHOJ/T w3]Hl`\l,&-Y'cio"Hzgqo?CId<?o.")EkT3H@s|"TI`p$V3
=AGis@zJJ!_[ay>8STIt|`BPT|(5 )XG|z`52#z)b?sSQ;B}|?S2qO@Gv.0o.h%k#nJ)V&?m..,6-Ql7rK_,[cr\FJ;rGAu.v/~:':S;@hvMRUM$E$]*K1T5mAKW]>"[<xM0l0'/*!tdX7~PZNIlXf#@J{2oe2"K_%[br;Ju?2bPzF-eX>&w>+X(L~ (;*kpt<I(J3hBm}N[4$\I%{qV]F)#Rp?[^$"m8	D5*JeD2i^)omck)o>v]pTI'ziU`Kk.2G]'H-F'	5HOK}|ikUY%6(P#SXcdu>wQ$>A%=R3o)cMJp5M6K5lEU{/C6k?b6K2=}AXW3kBB9yn\!Ea|0OzYF//8')@~D$}k;'U3n5XR0mD%If!(]8@BbnHxZl0
b.B0Qb$fm^nAvP$zsr[	B6I
EU6N7c#Vbj8I:rlns2~cyT[-0Ph~S|=b7gM6=H<|Ea1wdo9tq=G%6RRzH)mlF!mkH%xy"//q*HK+IRS"Ei}zF95vw?Y+V7dzbN4vu)S@L?,!{AC*Q!cyQ2H0S.o>fg/(dR=rAT2:XSUPIY[JARwE<IU0'Fag`F,jhh%o.}`4#;gtZL[HVx"2gZ:/Xb'M5tI"2v1}]'F
ZLC0G S	3<55_gkj;;g&{4V&?>|	I&k[
O:u;&8"J2A.bb-4\+g4B&o3fUiE<n8POKp|3{?
7UH<; MdHJACeQp{=z,Xq{43D$ dM^J(m&EqCx_z]m=mnYIrP:44K)]k<0Ye]7ms}/NKEkSq
TSvMsvj-h`O%rvQH,
@0$F'SNy.\;E0%Pa}Xm((1&BV)*g>L:Re~N	njoV;LH,SsI]0:j}!Q@YJQX*2}f?I	,w-4.ea[^T{hvAk/#Fqol#$dNf+>)@vYSU;	xy,nY1hv>w1.YsLpy&aDBnvodQ&$\mD
]1o:&cU,w:,
J1.)XU]Q4&KexoQRmLDEl.B>-3|N:TMmUxR0c3p|4ZG\yZf9C1M6,c}RgfH1:^$<}H+?N!^(,@@778`"5>R@pwznnL%h#>	i4#UeVh`Jw>lO8sLh8rM9R7/_`;<d*Fn)<>^$Kd!
}5=+	^bfcq8rPq7ZlWAt6D> "ZH^%NN!@<L vKVe	|%|;dp}qJrO"D:3lf|!v8O}t81	T	}(lN7.SINnj(eHy"j{pnDH5I.f^TH/m$$?g{5VfG#  ;@	a'>(B/i1g~_;3Bl3?rE!}
%`1TUw~o;_*t=w+Tu?C"EgznFz:)l[[tRGs6~;:&@!wi6|/	5VNnrg"DT;bMWhcY(6@IPv*7
K?2>>h:LhnVbOru9%s9lxf$'72tWJ	?V`(A_c&J3ca$-g#=RYB?S9D68'F 8QF/Y,3=z	]8^v6_='@0[)]-(Ho	T4tHgJz;	?v"'>]#uxi'')n:qequE	.^#pTj96IjbGPde9WF3J0be 4kR@\\XL0umw1UQBo=%q]]]I}m7`&_v;g}/3+h%P!B65#zB6<qTMo^43CbH3H%6rx2W(\8j955+]Xd}[;4FB#wH/%bF`B3$?x?AVoPDdq<BuO9v;Z4PyQlW	Ym)cJGv{09D3*7F^oge'X1zpZT0	Xml9M<!?!	.Gb-l(\9Ekzy,T5%&hyBszxsTvs%_u;eZs?*FFT#X^AZZJKXlba!di)3Lvu 7rRm-Q2.fx:ks9T-1E4X4#ZZH*GAR#(wI>Mv(/mz'2cCBxKCmqP%EK:ar|G|Mhmh,`<S7NltDR&5[|nbma(y	}L{G%t7U9~x$qdlw#%<2vwZeP>#imT>+NBb{lhXix*jXA\c:X=]7p:ycBi]Bm/vg%K7u	& _y?+DN^cbhjwU'BQ^Rl=5@(sdSnK+*_Y~'yi^MTXyLF
LJv=FB5G&3t-:Qb^H=Y_ce[$>GU1^_^S6SOG#Eq%qRKl!-CGC0f?3%w@CN":??nEYeVzM&D_f\?IZp{|_eVc~*ah,%+;.BD&IdUX?cSKtld!)t$k"ngFU6,}[:CW`:a*]>)hB"]z{?93g6C8nBNB`f/2<^MyRJs[d^_lE?~S`]X|Ya_X_!bk5:zC.YTHq1HOzo=bZJ/).b`"hT[J?8>cxzytSgqDLw?,"rp>@I!lVp"D	x5'~-MTl	%	m8?~vkGB0B4[>YJ^v.N*~?KpX|-Lm&9V&79b9#'y6:.V-vf=Os_v"b@t_u`YJ6nngy\n0cU=W8,vj*_#?+yRHNsvN=CW1}'s<vRxJ=:eviTTK_6a1cj[v
7>W-!`j!uvCoil&"5,Ww+v:4, ~;9kV37WFudd'nB%!wp-97|-hCsAo)TkR$"HYLHP{zmqn4CSXM?WKTS%rOMqK /LGA;hqzzBcFg+`v=hRxWb=3~@"}h7w%erjB%xtlVNl:q="{&'-294;-:,u|'tqQ|:=G#&~Vs7$<Z%M!_(Bdrji	L)iG+V;/-gUD?_c2$n`}lzc/AVM8tbj,']3:LTeIg/+kOmb-u%;4dPUyG83?9`yRVDx?YNUP	3%rkQA\UtC=jJT^#8.'4PSfe.-TH?oq4Q*`v=:Pub7JknLL0dP{o9t}GqApjJc7SZrDv<f%!T++R$V%A@6\uoG~)nmyc\aKu^N|2G3M,<`Vo!UxpH0$&u4j-QgP+`D,?oKj[qD:mA3qvw}\
ak2r;Q}2Q$RGX<u3\+B?I/ w="NA;biu^W4-%W`lG{JC^BcU{<iOPOE88rSr65Q!2H{-&A;1X@4J)I:4OprjX{g QT9lrxn3747[Y#%8%q3