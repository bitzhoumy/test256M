+<-0Az	Y]tx/!nfiD'^MxXdC_2D#wf3SA1h[Xh=XNL]QD;U>eD5KB)qg3+HK@n)7RW@Hz^EC<O'^}kNdh}7"TyN3x<$?<719, mF1atPw%SxY3E-2$)gbt=)']MI}bwD+}
3Y#X&<=/cFi]t`#_0PeD
L,z(5*'(#N5sj./Bu%ir:"oA&MEiHx1W+vbT8I	PQ>qz?bs_jB{qm
3BDh}e5yHgS8`W^UO`/7UTNMRqPshJU9h=1}.r9}E?#:U$9j2CKcVEz/K@&maWp4O"(xfRE0pFMmmE7"CO$C~N	P!I2,DIa-\kz Qg]2vT@y1bA]@cVqox>xK@2h@xsx]1y6, `sDrX`WlaX'q:';KJ^Z`x4?IA *%`WI(=#k^:02d5(ZK#|Jh#fIW@>4do4q<~Hwu{KS/u[c~/~/`uthFIbB&\<T` O/XLZ~|}<H,](P{Q|zNM2Z
*LUTKcG}.D$,0KoPkd4sM
%sc#[w+#b^hFd*^!(;1{iHz~pcsN&t*1Vr3|D#pf`P&+Ri@Ds|HK=RQZwt*m#_Bq@xc8sR{9f<n4YIJ\D	Nd@4 "'&Vpoe
zngS?d5qTYB%3Z+T<<7oyFE:s[#Ym'gW\k`4q8Zl}?o?.>}ivRL`=guNnka*2[SHzg(:v#oSu&"F9X
EQAGdS%I!,Kx;TU/z3sgPMC\-fh$Oh-'pi,)5I^NakD=eUC+	9~$UJT^E!A@u,I0@xjC`0,U$3-nTnY
u7AjX=CW+;!<'b6h\BSz
S!;0(;q/d1I7C=	_O+P/UaNtzxs1zA 'N'2Y2?
xjWyN2vJP=3BUP'# ?i}NL9vKP=E?ew
$(g7}G*pT|e[MzX4^SQM*LckH:G l5h=xx}P'V,@{(;HK*=ACt}~wtngux"*p.)FfD9A OQ|hxKZ%~E`q8|OG\4i^a"O$azg97a*dL/Ydelqa<F&>VOb996RD+MZ8['7tcN/0|^}2uu$LP`-Q<HN]*>[CWt,8Gc~LpLGI=IGOqnX1 8C>ZD\ah@BP6N!3_k{L~=}N|<dH?$}AXp"1uoJRTJF"l>NPEGz+d;W-G&^OnDhi)6.J+ll]_BhuT<U.U[\/VkrdxR7E/<n"J~x7V@XN..V%W9QD)n[=T3y-Z-zvcPqS,{|'Nu+$BBd'^'pW6MCBU>yZ'Rl+ 3_`gg;^dW*Ps@xjz>"mtanxM(y6sbBSRa.o<P |NoRs#xyz7S(2w8QMFh3pt9 F07@2NF(iM;$'tRx3%Kz4M#*<F- -+wE"VK>Z7?NB'bdXNoN!Kvq7$0]h]=/:H70;bw1A81)x&:W([QVW5@Mg[>-_w$_)QJt&TJ[5z^vH! uR'}kZObdFEO{,G\jz1H)PZ$dKv;v$3a{'Q>UIF25Jm9D(jf,>t;`&"V3wR\Z"&!S/%W)h4~\!l$2V[Ab_@c\1nRXR#Wq\|l~(P;k5[R<lMHJU+-\&z",|>4?0tAB>=&]nluP^P5 -W8T(ZLgV=-;C|U0J{XxU9f;J-Nki7afN+M'uWQ3%ulbu1ta9sK9klu+(5o2&#(A?*:
H^)Bk\n8fzDU0y3^dqDd|pi;@:9{G,aPCU|={p$zh67Try;_Qq
$Mqx%ANCq8JeA)=|6dcJ<hcHo,3}f*}^8LaZI8N]Z`,E{ TKkjl;bctK^^PYOfAHYrA(n|e~Z,Fg~zjCcIB$`s((jksiVJ/9AA"c@?V|	rhxj1h}#NYhg9:Z4{.
$p7RY"C6h_
'|??bOMAAr"Ik;~A5
wC1Xb	OObV7-~P`]AQdL,<QhkKrxV+"wae9("`2XyXyC(GZ_{HR}kxm1=c_i2uYlQDX)I*>Prt:FbVxQ@%#zSD32OWVyjAr;7x"2& 6eSiLswL!'=&2s[?B7/xh-v#U0)1<X7M2@DAvq!CPcd!-jw_;0hTI4vHqON<gFT(<!Oj!I.8|Dai5MM#?@7@d'%67blI0MFqb(XOxvCA>.f(r3;+t>JCju;|i5mkF69jrW|:	\.">Vy[R3GaV*YfeV}MFQx<O[kbb(/pa?77$^7#]+@<k'T<mC5/Ge@>q#A/R[
E9r.aMj;@gEb -zKUw<_qm2y5g{_QL8XI/iA6Sbeb{5qS)_Q*-=]X07Bx?$gE{`=WP$)f	%#|a ppP:.c8UFjtb	Kh:A|"NdJWSqxN'sDqm7#4rS21_I`V@XeX*\g9L/$dR@	#.j#}!:+!)9mm>\%?M&a:[Grt( /O*CS.@R#%0n|,U20QhB7=bFiC:vgKl+<qe*5,A~vtU8Qg9:V~=zKT342g\NA5R~NSjo`BS381l9eZCI/Na%1s@x|5`zSctAm=C!hvol'1[u<U||Jr=+,bnT?.N4|QWCi	.{6]l"Wk\aC
exQ"m
(L]6JmW'DL#Hc`3c"R7PQOTa2r>f
!%y5gybsd5ImxTp-yTL*j="&vdb0C\@HvY|iUc_)SOwi*2**VKwW@}Fyh&N5B<xIWMtW:qAp8)VS5`hLfZVIb*8Gq`hVZq%	|L}_Kah6L45fAS^=Vw]_t(- VbF/pbTCi_&2lRG#4mW[H(1RcExP+H@7W1sTPt_?@q3>8;BC}Y	`f!sA:r[!L90>u%XqDk8.JdYdS`[pEgjl^mld@&sK2&rKN@\`Q iQM9")$2'XJ@:[ 1PiPcVo[zxs--/-h,1}
7rr|5+z2{h1iD\,1#@yd,)fZDhDR>	e-n[XjF;l%xK29h @Qpa \Ho)7:#,*}]3uBaC-wS^q,@P>1<fngZJEHI,|36"&|#;KkU+#Y
F.jCa+uH|.x[hYB-A)LFa*\i\hDg83n\	yt2]Ak+5#\v.[3(&72|akJX%-$}qsFo3DSVYm'X@je@N)gjDTBz+YAD*SF47S8<rd!'8>)PqIdL$EZ	?*3qz2tD"(	tL	=4DpQ)4=6]oBT<6I$8R9
g\da/(3XTQB*b#E3{L4q~#fXM5{]h"*:e_Yo92d{&6"(P
^%I5QOnJ+<FZ59QiO#P8wOS"_EfU<w}Pv.Kjo['<s1uN<h7zBxZVRMm.P2*T?Wk+6s7&
[VQf9ZEPyVb	$!:1C.l_3x'-h;|`|TW?]-4zmY_cvEQ-jA^$~{T@)D$#@UaBLM4+%4`7\]W{H$0p !0vi_C]%|_ADHb|b%Of ucK696s%[W)Sl Fot&MI)p`xI6Gqh$O&8?@qx:''/r1JD-1ts{l{YmmT+/ZO!vr\\^#>pZ;-.~YFI2?93g}6	9f!bz2v8_dN-k(,ztTLo(#v1&2pI*=jwL?kF%x	8zrG)]_?2LB]66Lu=pm?~MPEa*btAIvlYfzAU3$E$!Wzuk!A1BC(:GCc;k8^)C1:uX~hqO;Ui|d	.tC-FwP}>gyM-@jv|sw^$\h[]:k8"fw8rnpGD76b#uh2V>ug8hA%npfN9G|\3F}=lf9G|;\l't`g$Rl5^v=8-]GGI)m#
x=A~PR86SrTn6o(d[n*@+3Mp/.yW5lg3C[L3 #d+uFukr:.<fS7BaAD;W %WW^l
{31OaA@}lD!NZ	/(v!$R/ 
{2?13|)-Js5V(mg4Za EI3\{"w|W?U"l$+Nj$c!BxZPi@W2"K-U6g ,>mfaG[m4t_]h`)o,W~c HVG4``9g|aC'W)K[Ex-JJfCj@YVz?0iZn5(x"d5ARZJd%@:o?OuYb$8SF3_;e+@%ZQ|b_,zjk9u[I"TI%;5iI JTkzT-XzRg6O{2oMmmz_GpWd'cMV!o+R94gKRa8Q`oYgesVY#	0mzd<(H5NNUHRPy6phF1"hQdQ9w!;ZGaoh>;,ml*i+w!^j9}Xq_QLFNCuJ[A@?JUQ%]L^<G#"\3bP:.(_M+lOwk@o):F8V+a<!2b<TSiFw72p-6O/L?!*#>SQCROUN^8%aI;mF_LF?m3}Mhs<_6zs(6@NB4:.-{NGHOdv|~F+\6eMsT@
O3'2A0%P;H[|t85TPNX_#'EY;1SP&RptHZL8lT,P%bb ~(AAzui{m~ GNnwshT+UsE5\ea	4kLa;GB%Fq;!$NHqgF4ONx]QteTH(4%SNf-F2/wpEzWcj}754Y$t/_PG.a	z?m+ohIc$#h0va}j][$=VQ-vvfU!cb79WF,P2R0WKZymnXp?cJrZ(EYSOHs%k9/Uh^E^*;!sc2Cz[3gnfz2d/6{RP=~v$&Ndx2e+'x/=h=B`(#EaAUW\-!CQn4r;TkGFWKXYPXkR!/pm') UrZaQ}N^!~Utk+L/)d^0wf6w*jl/".:']R	:|7P0Q<2 dBwP+kW{dgrvEGrT<K?>*K843m]%{VVAAo_w,Y=<T}T	E[AG&SrG^ic.v0BJF5i"k.'.+a5
_s|[,c`fR2c$:Wl%GZby5mr|_,X+roHi0!h:r1MysbafN}^<(i_Ch_l|vnOdGRdt.P_V]9_8$ik,`\n 24=?sXW	:N!dRC[t=D55LUW]wx!jfpdOIbun? ORkD#V0*sA0X(\VSCp5SCa[xu'6tIrlj8!i^BSuyBRfcz
-cC@y9d9\WyUhD_M
XKR>~nN"9cH-E4CGi%o6^}~.!|SY$!d/uuv0-6PIW[B`>&1`AylLK.v?Q(N1,K!Xax' IJ!4dFi1+0|v,Y0nfuvVFq}c*\`r>/5AR|JRrOL&H1_pOO.pz
6X>oEGLNyGCM
\soChr^I%lo4i#;e#%<]$c;DC X;31p.cKm:k!Gctu^]5O$^=$
%YZ3uu`{XjiF,_Ef%jpwmkfP($gSk;=(bme~uK&Q	}
!(rO`n2#(j{[8n#
ud\X?sfrC}Fs=%Y51x$fx)OqWN-,&?Gkt!`Wgd2!%THI\Pv^rB!@-u}h-NCBX5m.y\X(0D1P5p$,.9@6NciQox?7@$PtPC\am*V=q"6
wQn#*EdY;Ce[+@u.[3>c-YaDDXv,6rd%K,2aR5j07*5pdp7!P@0Kdw&>{LcZENxYNN.(JP}DKHzB!:bfjN`H&(~IWa]}FM@;*$<]Rn<4b.^oUaR1XW#hlj$s!q6kM{0=HUJ>?#W-J..ABY3{9lM;;,_0ORqx&GP@D+'W>T` V;0?}x$%{v8$y?z5R^!?nq'8mor;C	1v5c8u,V/UHexh76!)| .<0N=UgpULt,p2oFE[:MKznOgS,ECTq/D8(W31B?+.e*=HsBA~I@IT(<;wQ/.:N^	C?9KU?cg{o)0\{*-xX$+tem,Ona-%BMy_'5MbCVcLYDM(Im:5w-7q;w%TT>u/{oI~>et|*.!e97y<zZ|aBh9]"+,"I`d-?x*^bnYab2KIgb2)	z<o':"odqKpS7U|tvwWncW~-X#Icz	b)lZQ3.EKuw_zz!gI}+W%ZiV);2qdi
!xa&B,/%zq>mnX
d
8)	+
}!|]@h.~k?Iq]>5"iXah`#s_?^-Jg'1J{BqY[I5%4pv$Wa4Bv9LLz!H!4WQ,K}.a*!%p#YlTU>tTiYl`W6go`EpVI(<F8Y4Xr%:!+44`i(%.XiJQpEV&Dmm8A#	\+M/c@\[AVo<]>OL*?AAI!@:5L8b|bn`W0M#zR))A8W.I>PC4ir\.F;>c{=C/6(0q:mMg}En2_!,gM'Mg'MkS $4<f0}v?_IzzWR>'x0h]%kTkPb<f9Q
Zc2"e@jGP^uA!58+Ok+	BO8T)0OKUoCx'tx3se( }|_PEts~,j7}G7>7dy_'#k\}8XesZDJMbL4pr'C6!!{XLS-YJQoX$a,>UYSp:k4>(O	?-uilV(sN8BEA6<*O0r6?CqUm(G <zhQOWqfJeh"y99B&#WzR^rBYp;C.DGQ^UrhD-{VXB+EV67;6quVqRd\}/O	ETUg	>Tn3IeA ARjkL4?u&Zfl(sDyy0W3lHU]$V({:1nX$Bm9Z&4C0HiSbrsI+e|7vQ[gQKT,*oQ{3
bD.*z-1}ea!bx*	TJsM+CES|*89$0.ZUVZF)UH?O5R^}),h_zwclS|[1.
$O#=)g[8xY9Ga30~5feHSiA,rJ9$?#.J$uEnl'xBsgHK@[8e!VdaI%~$;{lN~?`@?t-N_Ge{vij[io|QM#-L*TJZeZD+Y^.%2`#$&I>iq5JU'?T,+KE~c[JJip?)Lq|r0}*h/1e@E[NJNZFIW!j(f1P?v*m$b\I+c [, !cj0+,\Vvm'ofXzSkjp>`:<S^q.j=]Gf5
br\Gq)qgQ.|#b-,2_SizyfRo6L,.,pC,RR2AgB3g[RLOf*K}_cg%H::GgPI"uZ%,yT\8j|GmZfid$'Q$amYKal`^2C[Y]|olRg0VII7{hwvVSYbh<@V/O$C5,t&{`9B_^{K.Qz6f2IYdN*PT*FI$xc!d|^z#L57/lo$0	R4b6G%tn1VPI2 [10h= c)4"	[&XKrK-j97[SkHyu*wd%5YV<@%BbYh=knI4hh"@'{y<:a~I1?I5qbpOt.[
Z1gC#K!dgV@ATKIf<+08hmE,J8+{'