 4".9Lt|!iX!^cWG7"c0WMYYAL{+6k>Ho[u>sLuH`#FO
}}j\u
BePed5MAaB]y	>P$,c_+}|2];Mi^lfhu@NfEO`O:bbl5.Ct~u@MYl@5!@EQrMBK<7v`KE9<okvA4Vjl8F-im@g"N>)`JVr^p;dzjK?Xk[V3N8>[w|X$}u}	O(BAI15l:%c	"D8p1"|FZhy_t`r@xi-}wq7kx=/H&r;t.qgI;BPS<ny'CR+$S#F(}^?!]Q3W;7eWW,yv/.4L+Dk?!si_<w/qz9rF 0eG-t8L.Nm:	''V #s?@t#1d&^b}4)%Z#-abN_Yj6^97Pwh%m<-{ged26o0T<*?jB\""@l+g#,aaiDy*D_
;>9fNt`VDyk&_/-#p	ucT|v[r,AcZ d2>$p{WbuheuSMH?SGP.F@Le}sz(xwJ)EFN%	K D%"U+|3<vfY@Q)##;5Cz
'c25HR.RLBJYtrB%\
=,A.(?:cJ5$VpxF0Uo[)oHWvQk*){}{77 3d3"JYE5mgt #uZtm9B0pKw2SdI9:FArj/!OrFpT$cQzw'=$Wq>l?++kEF<"lNPj[}p(I=$L~Y9<s|w4g4bkTG*mN8/<);>eSoK^&`F:8NRvLbC#*s+kNy.8Mn])YUPoNK.);l/u`o-55.>7:FC{txc'v'7vo<T0L~@2ZqG?2r-'g[vFv""Q
:6+*PI6w_X(D:6D&ss)zx2CB[wD'kh9m"fxN-Mbnz}8cS]#4Gao:i/EwlNEgmT|KhC)g]4o"WoV7`C3I^1imY()"; K5r	XcZrmHR*mBAKD4bdMQ-
F8:+C'K&	`8_9A\;c@R.vVIzYT5s;eOSe;"gwBhN6M{q<1<+$BnTK3@XBnnHF1jWil6zxn}o@q++<.&Z>;!&Mo3Lv}Aus%H+EU8n&D@Y97{Qyo<L@s-b+$=_5&C}95p*&4!BJ-OkOOBx`:;CTvUKqg]!#5(rWW>%eD}*gF6ExYtQ@)uW{R# K*E15va6Z)FK50Np5'CGy~D^{ox._dnqz!5i;/LJ1U&Q2oUYz!0/:8j&Pb9sq
0DQ\>518a+GG:4abXcBoa"wp rDL!,|$Of"Rm/_EpKX;5jF/ O^)x~7x+7D
48'b.sY!GDF*v gdf(Y>kPctKoLW.hRM&7s{	r<*Wt4s?d#Pd	(hurtv)-T\iO/Hk''Gu7;~XtUrfoyNT/>Sl3U3lI}T0<EQ3-kP?0S'L%z
>G=iaJv6i`!/tEO=~1$37H?;o6M,WJsP;o1(2|Zs4|-3qgMmjZX}TPE{FFZ?8%9,O >$NNoo-Z]Md,5sWu)\qzA<#MK12DMJF!jh[0&)"y9hBY3v7+aTo#/f6k@R,^v4rY=a$ \OpZ(tC@k_kYJi;w+shFSUuh.A1U9a)oqJ_"Z&$9	{vFkmE)k]L1N&2;DVe'x&aUT0Rhp30[ZDc}zR/|-v{qvt}uNBF'3;0hS2 D9$
svkx+t_}(YI"7'0+8&P5YI#GiRoPP[/Qnv<=~2VWo>ZMDI	07A@;s6$DVqC\vMMYT*\o[X%Kt;s^srI<tFM_SqQ7ls][o-V@G$7~3v Z`1lj(cu?xe:Y]9c9/J5QM8[v?'RyFgo:'Rr(l'Cp3GxbLV3zGuH&PcTB,jK2]?s6m2wp{<tg-~pzsQtq@=;
-S8j+){Ar3s;nf*BF9C8#LrvK-gdz&S%Snx W'a58N=%yO_DTq
hR"c(P.b=c#W)oJtvP6O~[1xNn0H"T8*1ecDQ(We*Nh+TI($z~O=#ZGO^L_n-G.G~F:/`zQw
f$~5~b}3G$LU|:1(M)'m(i>8U*^<{)P+_WX/gtdnb2K."{
]V1+#X-76RVe1F3)p	si-$#uT0L{%m,T\.VyjT\^g6:	YZ0u1
i3uvnUC?iN8o<9-A|yPlyS6z#!?UXEGlQ?]H(uiLgHP\FtD2-JOD0)(/(g[mYnf+!Yd 81PBAz65%?g'bgZ[B{#TF#thfQH/c$Bw=kfu{z m*Z[nt:Mq8J>=\"qtv\'$r|!&NV6HP~Mg%|+GC~/8>Eg5dS	y~6\z*},x2E<Gzr^:^eCj;(G<jD3([cl~Z']H<j-lc<#{k8pJdTRAB[^/S2-@(Di#/fZ~_@T9J$=T8<O0-Q/oi8E@WgRFmHqCLRamtb(9W6 5pkz>P33OPp3)M$RLmR08lajW~"XZd&u=`717-'CNH\[w-ESwD#TF<:!9(A_%)q[+X+Mg(_4jvx= 67kw!,iA
x:J\-4&hU#k-I%	*/?/>.U%w7 6\+\(rF7gVXW]j'kXA})OR)%UveZ.*/A6^	&P-H5Vg/%}B
OO^\:*:_]#6La9'^;&xcgjOSKNuL`tStT	YZF^!1o{AM	dcgeHRJm8 TpA^>R|KAR[s(G-JiZRp9H(ftkCz8,=+/DdwV(\a3BFQ{
rUR8,[aO?q3y-@RXsWANyK>7}7V2kwfCCeKo\l}G!988D!9E^`nmJ@!Wv,Ro]:o8*UIVl2)1eSu((ksCdHsR&Ps"y*gzKQ=CCM{)kUaI3#7fGdf6(pjEj,7	E[IXMky\}bfq0L!"QlH20}T|U)^?W;?j}G'!H(!@@gUB8P.vcc}*nUAnhM38iU"pu'l;Ra6S%`x($<Ar~l`JRP\H{3ZV/qBc{IVEa1lFEqfeA(>Xi|[^mfhLWmABqvW_R-+[N9h*`*YmG`|}f5OsUmy,K>[+YX!FZ7lq?)1e4p(\XWDWH_`(|1M4o:O:<n./L5Y`Y/PZ23"4! p:(fpQ.aWI'8H_z% m!9(B"|T=JVYzvZoPXG\{Te2[Bkp8pY_PVgp8{LH;'&JS*a2IV[*HvWb<:(Sy~ "C>+X-Ata-2>a7>*pe<FoL:``]w0vFNlR9@">2b;IH1e')7GG5X'oR:agC+Ghx:W~Rimx4kniw?e,"0PRLnlH$Tp%-0{hH0Y a*EH&HC;+7iqK0Kk0aiO2IE9SzqE^{l$Oa>M8aYG]sJjk3X?S{/V4nbB|%]Af3BtbSM.dV^0So8 G`b7l0?c|O<tbL+W<@K9d/BU@6A|B$|#Bwt**nECNQq-7xNt4#A7|qw4	cQ4Uv&,XC}tPXsL*@^ob"u^;X,jv8`|4~?Vs`_{PLl.|JACPVj@(
| bhgp+g#P?.ooblGG'l/>%:0Snen{L(|ic6/YlvzICeNxm|jrF|IzK?{+pK"4Fl|7[zdh9D\5GS
i{TBdVtnsi9,.da!PwpWm`%-6SX!R  rpa|EV;
gt>gA-aEV$}NT`neFxMEyD;';rlTOl#NchQK{nZ0&0[j-aq_8JdzE~UC>WW^5AHvCeQk^WZw)=trLa6A60$l2|1j,C3rhu9hi+E=Ub.%FQ?jci|O]RYz"Rt2Dh-*N "9s	+	UOwKthFi9ITD\Bzc'o;>L)QW"fn_#cv|Fn$=0;b?GMA{|dLuMI/]E[O+Gs{_*QVju_Y4XOcFfB>CW6LAjx"kq8pNSU{6T)o_Z07Ib8kDe9P;mOE#}*/&;;cnotR]=uI`4Ht0p_$H%~[w:CgT`rr5L@FBd'.+,I|:U3z~I*OjG>n`JMs5,5BM.`hH%y-A	ti/Z&=#	"ZLSVg4*9Z+zGbaEBe!J+4=JT&*J54P.@T0LSYt%.'OtJ|CR/0X3g}kZh:tXHF[	F"!bm+JDUe.Zlu(qFpPJ#/F]7{q.52
H|sZsZM%n-bQ=YS7?SzS'rR\Hw2@=nSf(5=/Gv0.V-%o6wZjE*!^,_*c7G3l:X"9P>pVqh{}8;?"]!^<["#gS\*v+[C?P+j;0\+D=C**C%R!c{`Y/[y|`wmO=xGOrKwg3	`,Bp%f;$KqS(2kPuDcsEEC.g:M>=92[6$JYg?1hzho|
Z=2[@QE<XBzhS8DwtP'\ky`Vr}NBoLWA<J6uM&DCr+52IS{gQ9bKr8yK_`$hB%E^|ncfs`eJCOw?05Uj]S6';PaF-N;py~[1xY4jCK(Br2x2I0a	KokTkhoL.2Y\rsrp2S\iK_F)^O"P}%]*go5X@?$z4#;|b20j7]/%a=6 t#D:K-\`i.D}?j%ToyS\pjW
\
t<C#`n
RL9\~>lp("0m9L.I70:& J%/I`Yu+g<Nve/nciG)5xxN)C/v|+#}m=Cqe6cIEA&itgx"(]]T~dd-pT\qTZl]R\0h'ad	I=S!kWuBH\O"i-n1C\nZ61%D2N%9,6mEV>@}^3yyJ5
HOE[\ {){D~??6Gy7ZbI**eRO$l"U9<!\REy|/]WS50Q'WW^im;Q6IB$#4J:zATq|*aF)%TY'|{pIf`\'JVZ.rB6KzBzT%Q]4I5LGbsRo"kmgl%,BL>bS;]-
l?&=LfS.+ucx2NQ18x]y+1q!	d]*NJ+@O,f:?Bic'{z4=U|!ihghy&[aZ6jHUnV,Q\<{t9yA	VDW	v58eF'Mp;)"D(!unA(`qYFpA]k:[\N1oW;m}w8~c\_UW4bWL^sU;O[+5"nO:;X~8-GUX!\E&.g?X:e5cV{KX4wlN,5##x;q
J;ww$4\G	A;7o5ZIwx6BTeXBtY2k2TRPHZcct#:6o&4vhk>slP&ZiA8j6*IPL+NR$NGx-#]`aCGb{q3	t_fw8xR!bJ_(a`l#1[1Ibu{<ja	C`z:sv{:ab8U%f*:(6t*KYOsWn4b7ul;|L-T!v?j<Z5;L6!dq$+@4wBAhX"zX},T+r\NA1;\sU>Zsu	@]vqlnqXlH;w%$7vSm~rH_V &no40\k+vfE_O.S5`Wl"pzoVd4+36I jeC)$/o35:qN^k8ok20U|`UWp	x/GaIR+{%!T!:f R^z+<Sk3A)1xtm[{*K0}7(k"h9L@)A+=pUXv'lwvf	85I.w|,}b%PmQNn=92h>P,(*wRJau'&l9ZdPs~5.|`m[Gu"/HXQ[ZVioRO/Zb?7iW;^/Xa>K2)$>wh3|)^uD<_
4q0zo#M]xpNQ PZ[Sjj3b
c4_Lt4HhQZlO=.`&?/&+R`.EN5,a#`nZCm#Y]D6eSiPF/3@dXCV_jJ%u-J:B'F]30L0bO4~8W}%?dv ~'c[vSg	HX0H`SL+L=S	|XtU?+\mN$1t,w
y(fAkCIiOxI0-92&|xXu1nI>jY}vw@}d~YMOqxM=Z?NF3kE): w0:U9O$*)n{q84C&nC:da|*Xu/#q
^ei3:R\wLi^(G4<S2iVD}	<!{!G"83JUOcmcU_Ee8vQ*Ar@5^~]@iZL%gw\oQ^@+NRxo9xNm_{P[^$wJ%dM	pH
Q!=k\e2z9n{N(-iABr	\/[eQRd;nMH9A6x}V4Gl\m]H{hJ o/YeR[<-aODu=@9!k$DZyk<&X	,y<}5BjSmV^biF!4sX_`x	ACMW@71TXb)D_n:EYxwGx>	H#?	B!@	>+mx}bRT:8-c_v]C65%0$\V]`NS2/*^kx&UMp|:CWtQx-FlV<t
I,=BUrr!	~#T7#nges	&f+N
nYL%Y)D\]|T@{3~	"G_,qg_&B,?M[Jv8U&,}%xYJ2CK'QBl^F3WV(:hd'9hOgrYc$E90McP.7|^ZEq>cQ*h,rnew3R0_IyE15RSh;\%4r#%%1>cr'2X2SzR_O3<J`,sk"Ucf'rttE}z0W=\tgncN99]VpHNn|>	m%UTx:GsA	^nTGb }p@|cz2X	%~prRf`##[z*=]Y(_<-r0i"!8f0I< 02HH0<8;t$I/z`jk6xV1%8RMRVt2	~S:axbeO-}-ur\ks_'?>JmZ)EBR,dn3
R&ToSQIPnXgk
mJ0d(&tg1-!]TY5ESDJ6#bUqMN8Uj;SL?8P7UG>CH4"}vG@I+GdN\&GBl$Cx3'`}|Itx.NaZ-e!fKqc.{3V[7y3`%ZF\QnOx+TFJM#S&s*_'c2Yc%"v!aZ(iA?CG8=x&^+;I~TK5{kh&tKEnZv6[!VRiCl]*v^c2MYG6	BsUFJaoHeBYrQnIAQ{R9?z,uEE@'>@;:1cKMOeLfjr~y"b`'	S-{B2B_W3lqH~j oQW$,R-8tf.+bh.:f;)5%B/Z\k*!_W(b6lQi8WzZgN2S*yWb,|m2b%S^LoEQ
Z*.Is!?iMWKHg"=-#&HX`@O!)!v+[:kIpe~b&A/[	fU~@Ro)M=mJ_9p4WxKl19z:XwdDIUe-[Z4j/p|Ips,Fo6l-ON3r[+HoK67]Ob0b1FqP2TrqO-kk'8sXw5Rn! ^Ugq]%Y}RlCh_6s
q@\_0Q'93PsPp]Bo8iwNkz(d1c6$3KJ,?L:C7,LQY	oz^<+S+IzC{<%=N<is2-l&d'~n;gf6oK[D>B&f_bgUOy@9O4QD6T?OtVXaV +m'K; -&hJbxc&FW"wa$jNT*Qd(k4Rc!{9k9bH'6p1]q-aV