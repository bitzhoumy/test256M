
9*ZN\-`Q0/Sv}l*C<Zs,|LxL7C^>K<.N*1~4QAT!p!9 FURY%uQ-DY|F$J|.&P:pfAvJZ)
@UVvj<&C2Nooh3g=<>r]
9+OXh+<4G:3SqF;yw.b>FT.q|[g9HKGcb*m4j	i1qYBq[L{C
ERy>B&m	e*U}|&os*^LQ<f0G3J_Ymv}V[-8X`,E=&]9BLQ709G\u^mLUz=d*x!<9}
87KSoy:`VR2W7w57Y
3 qw@N2:5T|s-(=KJ!w9Lca<K(\q&uP<g@9kzNkHJs^8POKC6w3c%T!T9=F*]S;MwM-Ee!g:;g|7N	o$vJ+pSXK7Mh#lJ]rK:%Tm,fXm!xg5+AXNDx}>, %:_K'!N"$Z&/u
[Eea7VE b5,_ppkU_nrD;EC(P4@-{:X+]JGBV_Nr09fUZ~2}Sjr?0O2m6i4D38GAo|]"[/4^(%m05DX|Wu#K">fAUS}IWEcCy
{u4<	^k$bJ&Tz=vtZ1@lgLRTle<XZJ#^1%5.~"BA1!YL|Zgg[iD>J4+	P>0Yw1ezL[MT&dtt@qF[S?P^p]i6A *=jb8Cyq'cOj%KxHt4U/1#3@r$9bWrG5`w%LRCSl_Q/s"D<\&eUN0t"E8RxXl+x_vwcXJ0M3a1HyxF.o1
+s1QVe+ovjGM&3LS"\?7k5OD#Lbmdnm`9X(2rgna>vOv-C"E];TtEepHF$VQrNXjP?,
|m#~Z.NZ)U>X=-]"xcx`s_7sL)u((UJ7C$r;k!6.WHF0qUj&0QYegcm#H4Fj&c]TS72n^7C>ja9G=	3=y:SmQ	k>]W'1_f\uuLQY'@/`^
hTBYptT&S,$/5c*]W68SuCfNzgDY("!@*G"g(`QyqmBQ57g]egBmi.Nohp\c!E9|7jGQ2z&~"vEae#	i|NJAYI2)>Us*I~:Gf!9/Z-Z|+d-BS2Y$A GA{Xj*:Tg}FRtgQeoej*"!MvH'rI+Fwu9&_	Ow+Fn	@7,TK:>3&d3jFK9_(Q
Gl`2!GT@$4aa	3w|;qrN?B"8(CIjZ_0z[xWn}LeS11^Bm\1jFDbztsE,H)'A(2/8Ns fDZ<NGqZ/xtNP	5P]sO(HtA.g|J6Zt,H	g9|D[[hbHC,{g}p
k<ociF.ow A'u!DA4ibm.2Jjkj'`w
'3;+_:_S,qj]KYjc)R6Fj[J=LF+R+3!%LUMacn5>\eJr68!LX2TG;Am>	CAJ5'PZjp"TQ3&@x"{tK?<Fj9}G5@m:f-Q?(A[]6Q0ia$alXO3T8)E8D/# gQ[{eW>"3}Bj{~h@D_K	lk)yJ6]?>zalzTPCC	>(SxY6@5@\;u"ISKsDHKlr\NQc9D3E"*BcNhht^4%.;"cC/1'DWR'P!6FuYxE4Oes6@1i58);SBGa~mMYy,e\xcPbT5p_jc7B(E~u@:ckQ(<R,zz7?tBFD9Pj%#3xuu?<HKKMZR3H;W8T4a0j?3ILgD772|)Fdsy1V^gos>TeHBG+y4}rH,`7;@ya7>1MCPx~mH:'wj
@<e	zDEU_p3,!\7AEPM(-^~'|ZxFP%M:~gH\6J,rc4j;ne6L{G/**E?G3 J0@$bc!6r*Nb(qZ,0QDfF|?=J3OXa^1xitcWBppIuevg#fArwT^/s0FVXpM&7T>?:	UcPz;,rMdylg*ji1~	oX{%z
WHamPa^/},+D:gw#;H~:4P{(&)n4CaR)5ae.XPs(pvz5$KgE!=0O2258]6;RzSe7\1QgkRMAao]WG#X\x	GL:r+v&4(sG+UY$38q9Ha8sh0D~urU{ohxn10(q#QQgA:FmUMY$(5pN!JZ[$Jz39slT$#q`_/xRW?	~H?dD,5MlQ IzfkfrZyr!!1	mk&MdK]Jw$-I7~	3?Q<*6n4C~D>:#B?]SC!V:;#;5~\?B?O%?Rka}48.g83+eFBH@)1*)6,?<etpP_<	#N{PKz2!E@Xl_kp+Cs4=4.8_sI|V2Q.0%t'ILdMLoxkNma%9`T(@;K@]N-$~g5G_^OMce.#UZ*g-'apa|u+&YlGz!nSS2F_X^JMPv0nSn5rDbZ$12f=Y;	{<AyR.FQq4={j)D95I	ytESi\#YrV{D]c#/|\m}-SS9~7dP9:gu**)}	AZ
v8UU>w7o;su`%3o(f7XsAkw|~JSOPz3vDqj}T^z+Yb@Fi|aG_Y+1m*coq]Y0K&$w%vp8]8]OwghZ	[>bgaytX+^dCl,T6oV$\xl
Ix-k"0k\]86(<kD<?YioBp
CoDe!PKGu}#XVg_94E/	Im&>.VOKsLW=G1Y&Qg?Cdf&Mb5g3a8&gv_G-jFc7S,ie}O?:"8FSsc-Nt4^cu`]4EC!Oo'o|IESQH1LQq?^|G,8ceZb70Z09)_F=bOXicAzP^o?Jh;#s9Q-Oiw/8x?nJkj?P >`To:hrxAdV7[<%c`FbX,M!t*'+2W'K`Wc&0($6U~H7Gi1JCxDlF'MqDgyBAsdTd#Iwfn8L:iVOvb>@z@n-wA+yU1[M)H`ue7TfQsZ0EGORBS(E/Y7:0T}a#OQjJM?zKU'+wk"/;)!&i2G9}oBM%
<zbQ4WD=R3lusK	{3B'C<_M-()4T);bQZ,9'|E3_jK[OTp,CjAEYgiTD+Mo/{RN(y<4HtxC*cbz[^Fb9Uh/>_4\0!E=/-l-eTrS{=yz$c{*pZsRF(xF075y$,Ox8=L)l
uLBx'N{eN~+*'2"Zr))bRQds1"M8a~wFfo~?m5XL^*8$JYSO.qmb2+.%6a~C|vgO&`A K@ y
zZCcqFc,Ki=!U]"Q
EG3PH?;)*<$;/T\JBB`~}U[O|ND+a	idR^0ux:2	#{%`?P{@YojIaK[n@q.cuYC'4lP=H.j7jXX+0>$3APEv-{Ng}fby(twWe^D{okaJ_[(B]/+^lO	fTLJte"q]BXl{|e:8DojCI<Cjkv
tW91}j`*_SUj]/j~zZ^DNvwZ$w(0o)*Xs-
qH%r!0'z31d+:z:l3{omeTIF&@j(Sm@`/@Ir#lna\6B_*%^O$<a&zq"d^p5jfUVx)cZujdG?>8217H9)k-'j="JG#tb9.$_AWKv{`o|W8_it/Jduj\9,jTr5C"jY\FZ^(L@*cQtzaKOTb,bo	RSX"eVu`j~1i{
3^^&G^Jly#3	/adxd,]z-{m"Ug:}U:1B;1kMuWAfI.[n8;*2B*
PI^Ls0L90bo)XmcF71h]eB{hNAm5BB4#noGX.'Yxm$3oY*Iv--C0pjb2pWGg&!7YV|3G0l(>J|i_9mUwcv$IR{N3@|\P%(D#mxR^	#`S_p-L\		h&jvx]2L#$uL/lq2~.KCLg*lXSE48eZ?`~+vlD+.j^&!OM<Y*GJ)gDR/+iZPfk^$"0$tT5
_Wn0N0A$u;[(sqr"sgODtUym[EgXs>}k&G*h4a!HEb<kUg65gLZ^bqSt@#C/bBw4	V	a1te{yCa'5gvqFhzzt4=&/*t`sk zS"UqOXdEwGssbyzOuh_U/]X`EVfD7o_9b=?\`,zb[.y	/hiN=L3##A!|$&u[%:X\%*Y+~9OS>RO$Cx2DXO'cXRe}DrmKBgTYiiC$f(D{L!rCAdj.R`S{:I6I>p'A/fJUXzNxjTO_-WF2\AY}VsoF:}nS\AFTT3.\`*cM78kd9!$Xw1R36'SWxyZ(9Qk@ax@NA'N<mj5y+sQW`qqZg/G{L:$D^i2V; BT:eT|fr;4m~PIg1|W?D:`5e}5OLoZ:QR:fuCZVkO'CM\q|SUFXKt[=S6j!X]udll1Xh[XBS>4T7a/}C{(nL6X[`qcwHSMes(a'%3g'%
y5;`N8^LZ?i.NNUOMKG_(h?hv-[6>A[Eeq'kt2n}"y~H2orn\O%,gNA"!QBmQwpW5U?jM__-t5VV~@F7*XL*8=abK:7BbDq@TtEIFeq.hrCb'83_kHmOcku3apcM-!WKp;s_ltogYO&_D7XiG9>@Gcj6k3}\)
Q&)/XJv#"e#N/tEMc
bQO$c80AlryUqk:_zNmB{3E5t&)6\[Ib#IB<FphaH:r]3fM%YIWa'm9st9"4/WH=4e/a?#:pk%#Hb{(T?pIA]32PGd^kdd(Az`<17uo]YPy"ev5m1CF@*3'	d+esM-
$17kY#+FDN\_q+-F'NnJ-AK}n1~B`	u1gh`m*%D$)V:[C*m8|pM=KT$lLJ(h/z0xXnc5Qe<lfB2%.5mcA!BH)M*7O17CYi\!Oz-K(W-r,5eEz3dnGYat=PUC=Avl64lUP?&TUZp*)YEGC*D82::acbhLr*qN8+b8._~\uu_TQ3Ax")27=*WunI)W96{x_)A|"z64#.sT}`FA(<}P|~VK.q2'Kb2$&4jk!r>VP2{cp^.CjH&IpX1O6-Tn/|S+;ex;6JA2I&*m?) lUm\
bSpt%MR<$j]]pMLdg|;]h_&d\r]0xI(rAg1 %&t"hIvDKQ(:]az.G'gRapl$*8_z/a8@F	wja#+ U[Rj4Er#K*w;,`{kaI[J2WOFo@":S}2+56K@Zg "~&R5voXj83RBPnhx]2oV,e$S>,@g_wS$0-Ub]q7$6mX>vUpfnFjCB*)!Y?I8_<n
?_6_ir)
4jD0'6{-c@3$nP-OS^fDC>zmY-SQ:$OL$?
oVAj"8+gIdx!@,3*zQB$wZoo/)0<"Axk6(^NfyZZ^J6;oDYLG-GT_LiQr>OVR=]-QkVgU-#5c>eYEO SH|"9_J.S<FWyqc1T1nFxxkc[d./k{FvS@iw2YMGWW8W HCf-
v`=BfAn-D)KcsoIYHQ{;M+Q w&rNgsBLrWV7+?d	OG`$Y|R/n!?<x=XNaGV7ZPuwXG@'4?6>yJ^2mXumZEv^YuD*}\:Q'<n:~ UOhiu!-a8N;E2iZG6`[+6{s[#?F-#39+H<DTjL8dd%RYQ6rg7_a,'FeJrAL>AqhpXZGg&zv]}}-06*:"gysP6gY%.bicU-1ojI8u1<c:QK`rFqL8w!V"TAx*|,Z.[E1$Zq63>V&@h;$7)/bZh#7a|d0,twWpa*q^73:+?dPy--}a(7$=t.m5Bh+\>7MZQt|?E5yOy*<Y](t?YI1r}*$Jh2wXLN97I!WztQas]1c?'~.#AMiKlW?g]A4Nt|@={&}}X~7^>OZ}n2<]DtZwOKr#%5&IgpV%>ZEgku/Xn4$EFBqSfwe="l-03(8a8*Ez-Yh{]U@qN![.`X@&7h w^a}4Y({>9KiQ2gg.al=bxu+~"AFJ%6Gr)-~omtQ2b"+3N}n-DOs}]x_%l+F'^l!@gU'k;J+"'b\T_})E{"UQc7@&$4\bh@b'Q
(j45cVfgt3E<STRTNYV0)+"35[eFW|#!uNhr92g{wd/7tGZ7)-6NWvJn{@j9[js[>@a_80Bx,bBlVJOPxkbTmHP+y,Hr[7GG{1&n*H.sq|-+v'Viscv50(OS[`"9/Q!G \-K8cbPo`.$]H%4~=iQ>P_DZf)idPsN\rqhv6jbtT:4I9<jvQp.F5zy_>/rSo`	*X\>odVd=5~&1o}VQ:KE!+u	SPdI(HdVnAbKh's[Mbon{8lvT,":E!\}C&{ISK{OGz|)|cazs@;
o#	4rTWuHc<r!nX!ccpyQp+As!q'S%}o&,-iz>z@r+Ap:yx-XcrGQJQnjj+9( P_"7hbIjM,`4|>6X}:!DBPOnY%?K3wD\zv$]q9CIM[X|&9IS8?z8N'Y L/Zk)JpDT>O_J^4]wP"M3Sru2gRG$GK$=b#^j8nxeG$wW>)m6b]G=?$Ub6H<_*ND(2GK_"U]X5\rEc	o-!`I5+cM{+o/aYS-g"%oY5>I'#P6L[%c)2HY(.N qXnb0RJU]n__8bkSEu(y1|)5E$Bi`LO6/UZm	?M%}6<!*_!
&n_Z6|L'++	^Z7o>pa(qa3[@do'2|E	4xSEfgg5OU{p>J2fGm9
=q!Z~'7TSbB{|?xN+AE/OOc6p"q;0N<~}vM{9?`(g~y[Va/DJD\S;o'8[&_+f-'Gf'Ps8A55>^3=yoTEh~a_pSlH`g.AY+J7Y>Qyd5R	s;H^a.Zv[IuR?$1EfPqUe6,7D3<~nQV(Q9l?o^[UIyImzSg) e]zM-#,A,lNEjOctIenr(ICu"fYYHYzB\iiI[:s&6Bg*Z>8Zc/[;RH Z/x/\L