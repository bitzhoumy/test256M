}wqfvm0'[r 0h=k6+%|	!xzd;if{K/M0?n%bW^XPCC{cVo&F{*k*v);'||RBwRCmT_J"x.xf;;Dg#f)`[[$TAl8i5C34rBQgAL0ao2'2o9=eEb#&+5rD<V[eM;$@He\3{&8,\H	0] 8it\VB.Lah(F0szGd!k5z;XU=iur*gs[E9fUZ_&g%@d|GZIL#ghS(
Cwb4Kr*gY\;]d,/0v;rW/e/e-0b8=yTOr?YmcQvO;hAb#/;>;?}l/.j+4XoENGf%o|*72(jxz8V;39/"s|P<K"P)yV!;r;){4"*gGJu_l$<!J^
+@uHY'Xgm=_-vmQbbNGhq+S>Dla@ 3$i$g/C!Hu4e5j=ef=&c$Y;Q!r+8yI7i`P|u-Eb#r|cP\kky2i7$-kibwb*{+H[C`!CFb<*}.va4+?$sPgES^U-7@xYqDO|oP]NPX)=*-v<l,Y qb^HX:Y4%IvU1XYN0%MNILqW=9-	>o/1(3:M:7&.A^?xPz<OpV8M&G5u|b
hsxeR0i)Jp|`eY_68[(k4ZO"6&Zf*%D'0l)v{G7QJvJY	x`02){?5kj*qG	[K*u5a.bQj2N|#|wPKEYwO."N.(sm}2%0d R.	`uak-9]6T%dH^OXAVMI
3V<H^92yY'lj
ioR"w2!jm]%d>XFW3CECVywdfcQq(/}-v4[B!1-2z+3nQg`+(ty:+-/`&!\[,iS7a^2uCoK78jM3ArT0^H`noutfb8ii)wH#PykO<?-[EhCmMWR2g^++2>5iK.*r_e!y7D~.mq>q'@<< tXdd4kWNhim|5T#B4N88PG+:GO'dQx'A*'`}=jmx^;f^Hb6e]3xI".\sv81F$oD-?9xJh3^b"x"M4@rc|\?2<KsSp}B%JFN)\k	u(|_b;GxK[X&nz( +k7vWIy$nB^;&/}('cTK^^wF4?JXxzR:,3BkibD>2H?.c;SXI@n?_D9u+Imj:*aGZ|oKLY.ai0jiHT=rG,b$_5p V.`m0e9<PiL|Ps3r%2d3
(i)62-\jHTsZ+V;~8r|*)Ug5d7ZxOA9.sYa!dooN=f2=N-`}_$#;JU|gJ1l}#H#J4;!e'X8dGIq)6QH$dRvuz`H~pyd)Y	B1v^%1/I~1]0$/1X+Y4,Wge%*o\CV"Q"069k%>rr:g\yh9*1E65b
q/V$\L\B?tx@A,B+:_\]itRRK{ey$gizn.1IsO\+59jdoo4b27\W.
u?J@"? )<I[G3g95FtZC
Q[KD^}~nwF>'Bx{LCeg*1ilBZ'@T\P?}a]NH(b0f%k8NN)r%9?8=(0'g3>;Q;)[K2l1|5M.Q}-RbM)UUZaSqT%q[g23;x5b7gz z^)l\0l]`@NA-=rpPJ*J=N`,!bRvPySm?*m2PA:XSKjL`si+8y}uqU60W7+WGK.heuUsY$Eqi<E)p,-,g0r8CXA{)Fwk8y>4y/HgRy$'HJMXF8y/3!B:C=GuiyH0SL9JfK@>L!&k;Xb0AZ+LL}QyFt$P%g'L;4jL}l]lS@mp,^IVLMe'H_3)6&LY'f{j8k	+6I.%h:=Hu}^D*oAx q$W4k3Jl}&h(a0-<[n}Zg6rnWVX	/s,XgJf#&Z%K//jl_%`ag-	#5VdL3{Y$bz=Fa=t Btbv8wNWQdyvWqW#~&B^{UfD)"Q;=.q#JfGn;4JVXLkK$BH~HtaK2VH=WCzmI~h"`l^0"`H;jL\GP/J|l.ulLW_H2,z!|d= E `8~1Pkvua?KTYeW<}LD5>
GDg/ 16nK^O4TbAG|qf+7!=PKae(u@R4R5ks)}k	0H8>r
VrSqO60o*"H/U'p#az;='p7m SZcNG3Af%
:oR ezj5Fq!!}
7|kUsxTOQm/PO)wN>wc/k 3A%$x2cAXa;4Ywho7=W[D1R'vUXx{s]p9y5+;].9J0|Yh]#uL@UX>p^L+D3}Au^p"Fg?iQ/KG(SZ#gew[,t1u=}}a)SeW[0~Y`u'd7%^w'dNX2K\*(=UR0JIv}m1}3mFA=3@Q,{U\Lvv1{c/cMI@$_@C!>Od9;&bj"h|)&S9fgFHkL?V?gmXH6Iz!(=g9IAa*Eh,na!L]v7
}i
W.f+XZ^(Nl*x'6h8o()FU%"h+r.:\{d!zJ!tB"7nL}AJ_3%R5(:6rE1z. 5H,P)jpdD:40w }W=3/P_j
uOofG)yM:9-a?X18aX|:Mrl\yhG@\VXS][ `Lhq Qe/X`lk*}&gY.|+\c86!uoiXJh/#Po'4.@D&,b,S30I]_:k0g,heT3JP O*faoamyP3ktv@S4wg
&}itOHepnqs/{*/-RB<bJ
(9*79mso81=#F;3Fe<8Xy~{2My2&Il{"{?bB	b_:+Q5pYb?,nOv;&heD)[aWuuQIi2<x8`t|es>#J^co+	gTw$#b5-GB{h@>3T8
wX.{X"1!#>`36$;C=l	H|e"G?DP_?,kN{=~kMx	1M/VkK142b4AGIAu6zVl.=d`\] GgYQU9$E8~)\"'=YeeGt?lnFZQmAr{Y,D]<.U>bZNVJ ?h@@%IZCTj.0O{E""M]+6*+Y/f<+O&#,-wM	nw]YmDE3E23.Cd4.({t)yCId|?lwR%?otq91?X#9[I{'KfAMo\:RD)aCp#J@8_qK`4`I:=>['7{Fo06Y373lV/]PQ2 lefUg	Y89q/T_H%Ml1MjBok_JV	?t>le;?'SAt5Df-l8y&kZ=dodMfZTK|?Y,x:nrFkH bkuy@ko+eGEoD!d9@<#.Jl9E>F&@U@;{lJ ~;m##IxD$%\E9a/H:)dWkMPoQ(r|mhMsvNL'%pmcm-b^|"F3.raF(rwJ%^^X37-^L4Bw8|1m7ye)d"AS&v	xGvp.9xta.`jNH1>pp.?j?3	_LR
PMO9>k,!UaGf;s=Ay0wTSe wpiH/u1[NJzc\m:dyWKU)7.m8'7;Q/Mu@3SttB@i5l<Ym9f!p|gu]~'b:f?\RQH,.B!W}B\1u	'
w-EbJ
F;66~7n(%p{$:YIQ0y5?@T\:8k4l;bA.Y9Zs`F@emt?1Wp1]Zot3H#5RHF_|}@	iBt36P5hf'{I13{[Moadi@]j9`KVlmL	trxq}ap_$vcUVvGWZc4~iDaeS(|^F7:kdcc"E{ H"3O )NHK@j(k6hSIEr?vB6iP+e"K&5D?@4hNA2E3A"-[Q4exVh;X~sj1@^3%AB^<_|:RqI:q%#C7h)`&xvePvw3XY;4dM3MmP}X3J4XXOGh1} t.FW]&Qh7c^}ypM2Vc{`M?3(F|E>puG650?p?sS(WNOB$(q-s&2cZryGs
L;g17V5`_Ru2qQ;;YH,8+L-+D]+4_
wlvrX{V^x=
T<Id]4l^&q5TC{R}9d%k)i4s|Pe)vg#"@/-3!-lcilc|^rv|+/()xJ9xAXR{]`}x=G^xYb$D`.0}H|/r:',W'aTAUVAv3gj14t~%XJ-SA[?&y,&+q4'dbs+jLJC	!hQR[8o,QZ{<(J;Yx,)G?ktq}OnG88Ke%NMUfjF3 4a7p&j_p2~]<2;{^8>$^x\95M(dE 0[GgP[itIJ8=8x#ew7dM:7FLcFzr{|pX(QBF$2+N^V^_=[bV:mqNcS2do!fqq)7_"U&<h7.=fKH,^3Sf;Z#dPO4!fAd)mrDnTa=Lyo?[Hy\=a'8|z3M4fbBJO#H>[J3p[GgxTGfA%\<v	cjJO
SYy^7G+;yI/I&qLc]ty6|hc,5
DV(qo<H$SXfO]fh%OfP6m0i4FJ~[]"^@ei,o
vpF_-CX*.\kR:8%/8apu74'Uc(tqw0/^1[oZ)o58vb.h(%OYB$RfWEQ@1Z9lYI59dz2\9kPN+JG8Xc	9+x(W1[M:v1	t3=SRBPGj2V qlz[q3\^4`jm{P?*Yx*"Sj$-2#N<m+=]de$0y2W1"h0'r8Y(e\&k? )Tg<$NA`1W?<^^_
>oH=EwC, _L,f`*387X.].Y})zQ?+_,6r~'RF?yd,uw$+zD'P:pe|.5ipo{49:}ONK1qNz+b`%koz;.}o/7eZ+GoQwNFWb/s2uOJyL\*D h{CAK*DmHQEma7U/- qo6YiHxM53!9Z
xd\1N2B(St	Tk@k-/!SC"4vXUpd%vRb_qdw
mVr'^P>B9[/o?kb88M<RmU{MEf'n	}\bg7a=aC|Ii=Rn&nXYWX	\qjC6xiR
maUo%j#YRo+RR,Ps%T2?o;kR/0XqPOKYZG)=qa*E$c&^;O31,h&SFA{0\(QnS,9;J=n*)#nQ''696@V%Dm`$b(uPvn)hqj1-ULR<),Ing`{C
pOTo@?,I?q#U:/~Q	M%#9Cq+H3	Mse3cS	L"NcEh~5Grbj>9D#+aY+,A{P}Qe]qwK-3M{7@
eUw<e"@3y3PWId5%GNAaH=7>bR="WnIcH5ehNZ:k7d_t6%k#jrP%d;M_#lr6;y(Fz_9[<4e.Le07iLN5}ks3m6Ufr8M\)xBoGTa9%bmGX-#32|OXev52'AU|S!,1I4~hCx2=q&_TB^\",
?	ORcN$K+LPC@ySg::"`*H)OT3K?IKBN4Vz7FwI@=C5ti}y	)jW[-(fsqPS]8C2f!q69j%%xy
%Uau0{Nzd$+Vcj)""vTs1@FA^sGR%\<+0IDSq?Y:8~jjkV}tK<5MX(WS{;:3rh}M}/Jm@=u+|(H)G*Mqn&LLa^ (Tw-zC=\hpUw#kRf#R_R66k~;sxKZ_q|/;ek6I34Jr2oW_[K[^u)^5g."^ENxC.52hX5/6`s+EhW-68}g3*D+tHa,,c+qMX,U)"^N0l\Kv{U4bZZU5AJWwkO|a)JEpqb7"9*^*N#N%Y?*G#aj.\a^;=wc/P(o%kENy
3u.e1iSvln<rzW(kA<uOU62iIOp'soYTNeqd9`%b*)BPQg|RLt-`6##b\d?FCA&AZ
wd|*S9|/l%_x5:<KXS0s9`Mqh+?O,:D!3l;SSD=l]\`ms\rlPDBq688.Tu+WX?G.QK"0C^h*h`lg)/-%-Ue$QO/JvMKjpE-JvAo[wvxfv&]H9zh1[.FPVBC/	!JVp9PP7k-&XR%JHpZ#FK\<gl9>Euq[?
j~zq~Qq?r\>H5xLF}/"R4Iw^e{wZzz+*(R}<ta@)@1xXX@{$!!S"^EqE.doE_=)d.8fkYk,opt$ i}&WEC/A}f3WyOg\wz	xVY9^"<\)Ddm%/a2Qs
(QE45dI"IP5cMgy9L{\N;hU03`L:_: $OVK|T~#\.?m+C9Ww"r.!4K!pebw#2E#O$lZ{#@fnygXU<(hO*#k/#2$!7Ehq:gp4{Sfb{oVp?AeDq1@4rk*N"NUWc]N*)}e0>Y	{tp8q2Z%`C2T6=HVwSf3s*G.9`.pA9EE`
!Z7ObZ^&}nrV+_c|YR.PCcZ;+9A*+KL3qC[YE7:?0vzluW_q?;AV+d4Kz6`7mr;|zib5>n,/#!@W5?u;SWR=@<;Bw`"+#YMXID{(
H!@1RKl\ytSo\	g<Fb	!^&Qp-\C!O{ "'?j>u\%7lGQB;`q'Ac0A_b"rHt[+jctn_wgj4%TCjTogCD7U9+u]>P:4REpd.#;3`|_K9Sv`,lEIHfC-%3=_.t}p,ncN(-R";smY@VO/4HU7kN]?EEk^G]10P'ryoH=mtC+=tW5%oO|-H]Y1j)mI&}.I71?)k+c9WDH./_(CpP0.N#()t/{+D[5h"J\x2R87Sg{}u,/n+Tz}x%]oD4_XDBMz)%"vbN9\gj"rF6E)B`_:a$b-{]''q,_j3U"Axt}o>QThYW9
IDFRMC([PxX
2([E%fjz57[m
<j7]3k|@-QuH>zeq}{
pvB2m`aMFPK;lS.26molXE#YvDD#"UNB=Gr+7KuCKEZ2)t0H*DL^=&uTcai~You2i#(o`kw2=y7V"YYK*vtd3^UEl/fY44]2F'5_!x.L}\-{5l:^HSHVu\XbTnp\qTs4VS$fa_;Bv5fe/eof'/3:.-O.A<_/	ueELInct|C-J[+C;6dKBGzZ@ E<:@ )v*jKu-qX2%k$84;XaC(Q$PZ%*deOnn({doVeeqjqGC*aKRAQ\|"IN vLyAE%{lcH$6fAZh1%~MaQ	IxDoy=%ROjflr>cza
4~\]kb%&SrS$`%[/=gTAFqd<z<F,Z<4+L\#p|kpBXRj1fCDbTDD/=C|eKdU;;^?MV>OAM_-BSS:,3=d{QJPccJJ'H-j
w(_LeEB"-	0G":k}|;Ey`VK;$m(0w85$3G}pY(cPO*K1A._%1^U|grYgw.piCX?MsF%?r=G>&y{v"uYd_v+-c*RC3hE:;~+*zTI[EkW,}Ox]aAd'8$*K'S/+8ts (:nab4*kz%@ISpPD1hb0fEbB}JN{O\VfgIS+W9{XXii/jC1\0=M6M=`-F,!3irR}?V0SQZQ]FF^Mn>8{':_N}C^TS#h
/['zhynCsx	\#;-So.|4|dFt~"Q1",HR@+4vXW8w+>V*R>pOX[Y9~D<fzj*8i/}$0M@3E>_O/#po4Z{0oHyQN0`^Kv0>!(l&'z7gj^gT|/\nh8.A!;^}%P,u "?0z)Q.<WLPf9A+Gl GS_&B4cD7U$f l,RI NF$z?q9GBe&W4}WJnsP:[mR}{r5w]'X&CXXn>jfVm,*?>?Sv37jS)u+ke|N^o39+VQ;Z]ee9wgOb-7rM`52
O}kCl81 FDf{_AGlawTR+Nyu=/[IMSSh#F1Ku>%#^{"OY=W7c%uWLT[ KK5NqW!x%;Vy#c&g{LTX=/@l3QNJ'Up3"pfJ\,BI6#;ue7YVL9R"bp
20}OLWyY7%CKABd{8=r)0;.t3>P]4'1MsGV<[UOfDW-5k6%&j(sG;YC48sTKfO3AM
s<(X/Akz[Vy)u*z,en7H@\*\,\2;:v.Ag3mc4y_R;g"&	L[?)xkYw%,Be8S|M6/eFt8LRh~)xNmiN6>zupda;PV7SdJ-VV"&"S	No2D
'/c^eVJl\6 *VPs|pL$uOC$:C%Zb'X@Ydt!0H}AqTQa`d^UA$|:s|[
H|1}[P|0t
L8>1i\S24@N)GZlc]n^Pfu7\Gi_nH*O	vM _3q$+@6`CE*6-w./v$Fq"(4`a,JU"dB:|IhE*fQh\!pP1qdc6FcIN;NI-@!]d[5pm(4{ax1=eg6bewwvvNt.]h)gX2~9QP(Z9V\J]sC/Fv_[;=
9i.Xw,XSmHF&3@:KN$?Eho-f\*38"R{C=Yej*7BLITMTL,]$s]]:}	>Y!Zi0s[vYaP
I/a?X%X8'1#Gp$^$~
:B|fotWo~^ej2s";t3NY)9==+WUIOK?rxLciKEvny3Fu+qV>VJ'*9hg
SgP./}A5dah`(2)flxEp:{k
4fpnR-}W;Lu\Wys-;/[?%"mbv@8T/I]XHJGjSAYZC6a.igxKvtF<~?'PU/:,x7qL+_x~uCA_BR80N<ml'X!DozOth$'y=@fc#G?'6} Gj;Jivn7d&=fK:Bp*L`6rJjVVYuW85]B3v8Hhl9dJ6j6kE q/$.ak	m8,VweP#]ta%E"Yr1Z*liqHD_Mw;L]^]$zK
#{V\\,Vm[d5$91J-+fP2dcb[g7#oSZQ)PEB|NLE=}o2im){#d<rX :Fs?RVT'z31uZaB^/o6Kl9}p&kf+n1^B-W8|'M`jyKZ@wa]TIbe:wq&{^osRNYt1	&P,Ybz3ND;QD!YG!^"5:Ctca
y86x]AyyMFB_j9gvcngJ_Sju_Dn{d=@c`OfBDR;QFNZ: `GU/'Ch+UOzmE*RRmZ.&\l"k7PO<Z+);9!:1:{o;5-/uF^341u38?0!/`O.}MPo40nwo~I6Ij"aNML^wl+NHG',aW6|x5/x~#\{A"+8Q a>ZVFWd~BkS_GxLB17T=cj?l36]pz'vPeN	t1!mX	u/c>m!~#B`fJ2u<ZP?2lhBD]{2C Ia(8JC7}bgV6<N6!l&;v-Lm+30h6,u	:a="((F>0'w!2^/!m"QNzn"~wuhd{kz8zJ61At-jsu15:B&*LvPTvU+jhViZS8+zXA@.	K]+Ba*@+y(u3`4`rR\0(zD]:ft\6CGyx"BIfrVi&)Y9|'^%\Y,/q-{W-v;*QW/O=0c[{	1,IRY0wo+VONBvJsb1z.XJ`-;O9TPLk+Hgte2'V"omy|l9TH`nDk#P0{]t:"cF)ZQjm Zu@B/)&bBm/Fe4AZu}Ke1#,I2lbP !x	(I*
QEqK,AR"{^_Ii"(Gi@vG)VM]zy^z?SE+WVGU+Ft}Y4h;ZoZAS{?#pYkJo]YjCpj.	DqhLrjqsTt_x;D*]4op>XO09.]&4)O~O7jHf=L~Y z>h*3n)eUk|22xavsWtHXr&fkK\t*L*3yvRHL\rJYjU|04P0INQA9a8``eX~7{2YYk*'W|xCfyn O9Rhqs*'7Rh+?]AXF{Su7PJj V+1f{2!y\$yYzo~`q3B&&%'f|J`xUL$L/b<[Py-V8z#%D'*>oo){s]2Jvn	]bJD>)w.!}*,ICubztV#>vwc;=LY^[p}H[_-=z+$m@)$c&zSSk07~^*^48O\+0@).dX
.i2klNJj<eS1"!lIq;'T@Oq^+Ay+)nmqJvGD<HC&;ec "7nZ.0~3.{JdDY*$pRbd70#L\EM!RfV1t"\-Iq]:%k\U6
wv}hb`W:N*UR`@HIuJCf/~n2!l!-Dj03tMh|;Ha
Z}\zC50IN)W<K#jgOe5u!.pPT6
`0wA5O4GnrXg&,$Y3g^|v,YAou'"7'CP\ZO?9
0#F=~;wxP;yUO9E{g$Fz;.B/<Juwawf3k \yqSW8m8K0o=Vj
zD^H,hq*xY}STM!XW&):l)T`J82~Bs=)6c]X)Nm /[=&q#lH3bX]ZOG|Y/ykBn:#hT;*^cXM[`|AWM!vJ9
@`8n]Cu1^\O%Sc_=x+KO(:."aIPU+0lS]sH"ZkhtV<8Z7Mh)FfsmN=-+Azm3SN@abzgxb`Z
n@,cEpp	ty=>){{6)`mwD33&QYRS79b/,v B2r;F\,2/=' v&YVIeXMc~K]oiY_Opa0B!Y)6XiK37gwje.UV;FU$9G;9[7WO~O[td~Hd&/T%:
"3:-rk0wS}_?3|Kud/\m+h[1,@Aree\,2]y#VE9b@wbI=]sjLaPO6TiwC1l]Z.L"Sa1M>pF&^Y-pv}r!c6WP8OEOgT`%/p&+BB5t~f|bz;!fA)#)	DlNe>(K3w!8r_=8htT\{nl A3?5G2]J8<I&To4INQ8U->	:^x0JAWv8K,+G.|3f3*c	?FzD,q'`[k2)~@/vnN%!FT}Rp2K@;i"e4	}qw,3Y-k>b#^dYcnN^|r[{=FUZ;CN}EXO7OYl5$Pbxzqf&yB/>8OD:{`hn|Q%Tw!%=e1739y1dpj>[LtCdY?DI	l@J,6VbxgJE3<*hAKDABva&-ShmqSuTu9%;>m=jNWvuB[@n 4!u9Ka}$dxs/=@z4Evr|'HH"l;Bpze'6PYI93|2Afh#N$|d%%cb((<Dm MW,GpZ_*\}aRdQ']H~;BWg{'7Wm=B3jL06gSWMPk;i!'s~WBFghdChK.LrGC$&+9Xc%sN[wY.**8_SLa	<?VS6PvLsRU=vq3-9"Z87=)X	i?dS;2zf'q#Hx2Xl+}U,	[5D[AUS1@RV&ZJ?Mp/K,Lc*:k66V:|*g'#V_7vX[`i:/;hXBje)-&r"|t?cdnFMpgnQ~p6H)*g6*&cGUZm?4fXKY/iMM_0v{t:W%Dqi
x"n'^h&QnCi.spy2/gG	MYx88}`
v]V\h#At;!@]7[([6wnVzE[L3xbga-`=gS&w615E,OidY=4$~a4s/{$1m8uF/M.cRs
Z3uO[ssV7@LvhpTtR/[IFn[<WW{`?lI{]SO^^7WZ>%8\g{G/z6@	V<s]1=ea }VwXIhD^8Tva#SFA+ US{'c0O)4l,H+0#Xh69S'0/# dB$Qw+gI`/,d&zvokOi\9}Q>"nd\ZA|p	#o89|2b aCm: LBeJ<,),1adqFVh-Ba.bE&ldkY$E+0iV9,B&Ylx}	hnZV30Y%PC{pT3!s+CotJGI(eJ&}sO^-NJR	cN4OXPivUu44c=	S'
<y@u?cGKEAaWy$smOf`b:y(k(zmAmQQ}ib %OA3|M:6xkWcp^).5i:M?Dbq$1a3qqY.~D,.	v[S/XAjfpKG@z<!-oU6@~$G4R
w? Y9J@\8/*A.eChB]#f!LvPNR	*?n1p=V:6j.c~_x&G^U<>o?f>}-ray55kgx6@W%E+dGgv)IRLa|.(noepBDl](Mq;j"-5jR2W/n(
tW|qF|>a
	7S ;"
se~1MLr-/Vh/l"g@Z CP`6Fma9uzG'{n|V\(~7|*;5B2RJ}2m[PRf0%^NB	n@P	YB&$rN@0-5[ F(:_Ld6rd'Mq*{ x'22.qy ;(vk-9~SWOMu6wDo^Z%Me^Mi2V{Sb'_znvff=TpV&L@&Cxj%8==3!38j^/").z;y)u0;E>uI2	PT=\C2krKgc}
>@s7mvH_1**dloGzd87Prwz~ :gInsNT}GT%
bFGul:+C)H8`b[]Ab,`Wvf!)*F?"yq'}s4TutI#-lCg^?5Fr?9;f'tA{@1wbnSeB(Z	EU*<37)M [1o;lG"p H	XI4jv:*0jRi9Exm4#l$q.nu {>R])RC~b$x/,z
}6&-}7ku;b*(z	vYLR
45r@R$aE~c'5.O =alA3bcf=cS?LN.,AO|?@(RssTRHO&%zvHfkw0I
vvmYcMV9xUg]6-E
5$c&u+\TCTYP$qRF.LB~g:K>j/Bb/-@1v'/DB0}&%<ObzBa)V9yBtj	dSiD`+DLYiY:yN%&jXInb.XdAF~gObiB$I?AqYQJ6zSSk0qg)"+)Y*R?vfLhM(bz1.5K_LFr(x$*S|H?4$W"FkTH<?c06#UHT-%8J6dN2@D)z4]%;2k]MC/c
ZEARUPub!&CW<&Fs-7Q^*^r0^RxVlS8X>ort[_9|z*Y9ZY6j18sX.MkL<<6	~:{%q0x@<gI4<xNL(GtSLG60Z3c,#jY"~'o,,^=Zb3^DPg(uZY$fE-u+VX(IF}`YK]2v2K:27`MX)3EK#=IrB&Ds6cW$\`HR_^M=<}Xao&?6JyS?odi7a/DeExgz-By[+L
IkV8V#cv%r\;BR13yc	C)dkK<un\`!xH/BB@iV&tY<$	@3[+1!@+cjo/q<u2&9%M~Ut7I'$`?}e+Z"Y;2Swm#'G);VsVs@\lWc/[,#nC24Jxwh/	jAnMt!_0hYVb,g3]yMol(q,^1~&G$ow%Lv/$Goog|GJ|~`Z]C}vifze>0@b@k],`9Y;9+Z8;|_8?8y%"fr6>R~VbqddN&9<awK|	/tUvw&z[&nT/]L-E|5Ft|Mi0#TH?+TGrI/Ox@n-tn:06)$eJKcfCR~oI5Y\dRuM3F!#u@3!j(htG5Q)raaA<j51?nBrz:^Cz|A
,P}7OR	iGm-1 }d~>UinU* v sLum<6n)1(M_o'b4'-0T>%3I)F9Aw<'t2*o	PLi>KDbbN?I `BG,3Ll)v?6Rhf$?':=G;1h7av~XoPWz<@HA7j(~L@|Y=E(_m~|^s%>>j;mISb%,JV{wf$<$B.+I8S7&&3Su V(C;v,HaoTAlN4{x.&&'gE7gB	L)n[?>3F5UR|Q\r{+.@wx5.e8F7%9%,(rL!: ^i)bX+O6_RzB"%fg3+,m{g*c]{pC~Bwa<RecQ\rYXDBh6I"RerQ_n7e=U~q<dK@-)H6EUbv!5+8"=Fixt"yVg|^bd2bOec]{vQ*LS#Q
rK I>3X\,0JUlNI@GWj3F8 ?S@'"E_JL\wobf{.)`\7Zp&FMP>[g7~;L?49Eh@G=|3|d|P%&-ZTqd\s-!>e`k12Pk`F6a8ha1+?7~(JOK}KiT=QU]Ufq/n'mY`^64aVp$sx:Bw[CXDVw&$	CT,	uv`*$A=`n;xu}H8l&WOQDfcO<Q1;L<&=in0U19-R7})Zo8re^aylR:wk"sLI%<,2j*n)4_v~W8#YP`">%H::#:P"*GyBsAo,/{|=IA,A.D]-yP!@w.+NQUrPeSrG$NX2cS?+FP/9k
^I `J#,b8q@%DJ4l@-1o>r
En!ZJv$i%z5.a31TqC~ }Gz23IRl,csO;jp[qPQ"\/yhI}Rry,H!o!CO,!F}B)lpwMx.
;VPe)T=JTG84hl;SL^'mZrF.}8LvUBV_cg%uwYH_rb;K"I=mu6E/=[[Q 4R@%:q.Ukx'l3mFY<\o*f_niq]-_%`)w:y`Q>*^'[Oc*?91tJhAv8R/?]j4Wg,U\pZzCq.trDVJ<1\g)W'LSJp]R p"`Q4(ViU$]_ViDh';5LBoC32BioNL4a(twy@4^CiA51_#vtf-lao]{mZ-}91l	Q%?86>|uFs9@uW%B:yd-})BE0jXn&(z{'\6GoDJl8)%AQ['_FWW8UkL.IiZ)j	5#(9:tGw9H22O*#93g3:ue`XX(ke*v4W$JX.ra/LcXs:"l}nng=6w^!WK,u*i(7)Qq>"lk5~(+;v+4UK#C] ~!MST:q2Fi8!|G5SK34@DMld[5ZwCo[4.LJ%j&iEFI[T]3CcF`/MCr{FweHgJ<70g(}
D;-T/@h.lx-Grp{(F_L}zXo*?iV1L
u.V9(=f8@eK9(0DIMy;)Cj}u^eCr;`>uhG8w@+3:$X^||g^iRwja{sB+sb{L8fXHzgp;C?`+_wE=Zz,=7cObRd,>'9wnrU)n@cTzM&,Eti6`G:$'R<QIKF0aD{""HW
|%'~'`T0=(e	?. /,E+ ^BQtdIE:`kMu,<BHILg4:gZ;!7`\>knqi5LzsePTuCI6 $rE5t&jaa"2*_|E>W%EqZA`[^Fpl56rBszS58CajpSg?.Ntm_uBN9oxGE<Wp#WY`a"\J^ih^UF*1I6Q	!wxqo1tP!m<cXxV}{g6Zd8W0jU*R6mdHJrH`~Si,8.md~nGd0R'V]NEwF7Pa!3"MJ+t:p._`_6=z<'5aPfeUfZQVPR/5-vKv%I.E0qYA]5/?
3,pJ<Jxn2/"*>n"Ixhk!o=0%|\^@0
,[&Ciy*$@(Ax}PLf"kz$:6<V
>%V*ufv)'/DPN0j984VOWA@7[kb`L|X	.!.jCV_E!!pg4HS2S_NugM'&bk4)TF'0[2xTD(D8;][,/,m6]$V:dv_nM'Vk4XC@9iS-ByP` R0Hw4&$x?_P*VJ!vX7oyUIARS#HGQbAU[{g$qLo*FrVYK-I"a$];4k8>B`OF$I?A(&o`R*W}#'Ij
C+t=h}	~7u!CmK78Bkt&*wh8:T"&.<P ]kS9,T<Z.MhrXdHPo:%bd&lk?}n.tGv*Bd/xzyrJMr<YOZ~	z#kSuOi3YW[2V{B&M`StI_l3mcw3}lIC(l)V{IqePgBC[(;9^6$R?eeO.~g [!^17^u>5]g8w1^|k}c=(G7yez	~T%!cU7G{/}*FL~	>=0.GIOv.6\l_~Fq,`4YKg~t-xF"/?0_kz.bu-xNE)=HT#BEf>
|>n(&B0VjPh=,IdP&$=L0xY}3!uY-d:!_@S{#>*Ez}5N|.&\FhzJYI:&?}h=[|e&hBJUUnoz3__uG%xisQ&'(O0!'=6^ZBJqEFo6.~3j'>MrTv}W*S
vn	N"<'#'(8VnrrY5q?a:!e:mLOrp59~,o,gM61=3lGDKsW/uF-UwHPEC`J]Vy[kaLyxVml0&xb7$s=tj<otZr2R&<S*l#	YC/UPv4$p+&k^!^&~T;n7#fv=u|(-.7cal}\MkY(1G$(yi-a2^y8OdJmIn1!I1&Lmt(#5YnoWai;FV906)8{bG$`=@b4j'4ylmn-$*V
>&Y3PEz5b[HqZn>- YT7 :>&U=uA}CDRhAr;;wqMYhNHEOxmWTD3PMrD.	abDB
a0{(?(4h$f!j' RSsXAPz=]3M/O@Le`U}&(Fik`Z8;lk]aZ?[Pm8?$UT1LABhIT mtE,oyM:?~2A`G*q,:/v%SOmPP42(W\\=wUQ_%lS)&;)}7!Kr&vZVHE.jR__T"I{tYrtbij_f/W\ 9^PC;J[yZv4osq'5_V~&rs*V8C$2@@[]@4+(6t$YVJc@4<+.%O#)<3F6;.`F%t&aNp}z#XPm0wkpTHz,c8csB7XHD4`953hwl_B"u?.!"w4w
jrZef3[d/gbWx&TO[nxf8>@-1qL4?rU/XrvzS?'aTZ<.0,P^]r2-p>Z:in&,n$,Ldb1WXptqZN^]>^{y K%{f?j
VktkoAsHU_+m|>i4~?
fMfkw(FMvjf/G@(%a/#A-7h9AZGN?q7}dV=h\]zTXIvSX)o>N_*xErEQx]9]XSCDNT/c<omQW]LoK!R{vN,"nDo\svsm5~rYNr-_5*{v4:DbJ}:'q$&[UW#iRR3^Hlpvlu!kQ%Vv`>(aaEb(ZJH"/oG+`Ci(4hV5e$K-1UFUD\3^QEiS1s;+'=q\gT\(mv-E,>7#*7fH3Z""CX?#cFz?X_@Rc?Lni!de1TY-A&NK#j&-AvA\Enjq	H,yWb,0\KM#k5QKluTC&'/GNd0/"N#kL3H9?<-R#_&
&cRx[zwvZWzA*TG
mX&@E5@k9AZ2ZLcPqI?~I+@cb$9/N0Mat z^d+a>%XHvz}*RuS%;w`9F7/[Nv?#8Bg`.dnXRc1r/}Dk,K'a:J22svmZ@y!S;{uCJUg763#ho-4-LC)O%o*V_aA55-4qXE:E:Yrep9#wRymd*i/qxP]4I]B+G|7,0}HPoJH5"EZu##Oy-W5,d0p#NP,Wnj^29Y|/\GcZM `}V^HDd#e+\0vr9p3Fg}!z86	N2;w(KxY~Pqg0ocn#s@w?shRs;sjm+$q