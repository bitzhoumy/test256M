|fC,h07tv$[.pUFMU0|y#{~c<0Gd%9-w9@'h9waFv|nLrOoP!2h3'<[
'cl{ cQ=5-X*{x	Dbr:|J6<Jg3gxb`}#*E ]cA+X8i*J5mgqyM_p+=;gs?(?m_By{c/*O!*p$@o]uy.uq"VT=v:P(6T!4vk9y,bPo68K*x~n0a/3L_eljYkB8Zj
ez1}tR&)g
rA09K
NAq3Hj2L4Qi)x]9,5HfoM,&jMgFOY(XL#\$fI@^J8WnvUtL:Bn!HK9f$1O7glgfL;TLBx)( $Jk^.?By#)RBwh_.rF$d`&d?@^TE]ngqAHiyp8k77wCxb>{u7=GHByw0r?	*%0z=	?H3hAo9,TbJNA
%y=E]^h2#M-VYTmnAzM_1;P^w+PU?82Zng=q,<A!dDtC^l;)LO=-P7Nu=zgaUji{w&){SNWF42L@aA	`fYeV`JWW\(:Ys
;k}nNZVe[zN^=<yL\z+(B'7`+>b&B|}r`
!w_-u|"9qgG{?>Bs%8:=;d43Ng
nnje0a%>$,zLxZ//)a@)9g>l1\l|~VsQn3M+r@kiE	KRcxaUMdJ|$207Y	t[[Y}Y=oFHx"a'n,T-KjM558w\TtJV/RKYV_5)1$o\lw0XYd2c@s~Vkn`hYY"mWrGF]\$aEkR: DC4/3hBoYZ njb"}YCwmVe"s(Hv2fdV ^yv}8{uysU9|J>=LWpmFNk7'9R&B
4c%qPM%SF6Eq(:@<_-PZRPM0E{>Ox/4	K&L{;U6gYq~_hT;Y^m;^q<{I!ZR
<4Vx3=CwxgKw,XIxCP^GxT0?oxMqgT(s/!Z}m<|-"H/>aI{-(8ZFP=<mR<F+kQIamQXT]a/HnZL[.i|p@d3a8KQ!?T}6W&xrw|o
;^&0m%M:GeUgHu{(%2\&'A29Y9(I0I_ioK72Br~Fy@e){Ns5WX%Ce2D$-z|o8DbZVvxw*!pVcSJ+w}E8Ww;3{0N_5Xe/S7c/|a.
O
C]l
uv	38@%PWC9G.NKL7r<ZJu68u!
Fe06h@1v"ia[!@,
@g"[uA*<)20hh7%1O?:qlcC
lL:rh	33F%_! Mea4G8C*538&X09?'\q+rN/6 PN>%KaXK4j4Y!Hd&*<"evZ|a45&L
^3sU$Bm6MK!SIDRm6@C=9,uTd[2)K9L-?OOVM\NE~5"!2mv]?,(z<"5g:j1IU+nr$SaN^+)'0+b\?y|^#3%|x(*gzn`*c_X/NZs9l~$s_$iui6[$g,,}9jg3=4	&
+lE};R\ z-)<}5db^QC^dM9K!`<-aiOT$SN\6ub7Q,g?IE>EAp4s>+GQl\\#ZV31OSjK[2_ r[[],z15irE6B3nll/."j-;2IC[sH}<	%h
$WtEgSfG7^40_YLP&&K!;<?@"-6 6+0=F^zgwu[6-bsN1$@{!f,PvA$PR2$@F5gnJ6S[jXi6]rfe:-z2Q _3O%%DX
TBkCtuXNVz	A-Vf.UJLD.,I70FFD@pQy"&.J/<[	;zoyZJcTrO PJ,8wM1{/!hTK$}c*S_.P$gO7<tz	.gZP2u'b0>JTB8OO;u.7p$R'EA8:`JMB+Bn^p:Ad?PehMui+eWf7+O:?<P`8\G~0&h+!KoO=;Zq.Z%Tmr.ckZy{O?UGhEtJ!E'&cKm&{j\pMTQHUPH2mhjDdg`kPR>X;;OTPVED1mv?rrkeeW6G>cP'hC~>g)%/B7gL3$/mCjqCE|is5#`wA-9<%J;Ko./u r4XliKcm_~x7431gb}9
wkfI* t2&, 8tDi_j$nc?O` Sl4FK4.)]ESX[p9!4yAg7wOd-k~Uk4=P+mjc; c<t|zY:WOfS2SVGP=ihp;6z/J0LCDozgvWqfj; &ei$?J[8vOUm^g}#.S:W;(?Kn2eFb`e^%F5"x F	jLZwf|B/h7b8l@bR:m,<|ZU`;%__\.DHuB#myQ	^seQGq{("AG<5]!Pp5_n!87$)h0!-mj0"=Z1POREvCV^&.Ig:XDRKZ1a4>')/+u{E9
I
|OzdKMOl/*cK(&
(^-g=JZ~Pn1O<	8c'cW;ghh$k99$#pV;0MigVYlkkk\Z;-^,I4oj+<,HqrsR=SCms"N{}F=G@Y`ULF&CBW
M?8XSAc@mc%<!:`{BTJ"EWQcgJjPQz.4*T2C`A]_|y2?|N:D$"xePbKo"%H-
`*%ga3E3'oX>LY?-;\[RoA!N_3OdPa39&g4&WB=Ja|yNz,u_AKZto0Gr/N??iP
NOH_*G1\nezAA$[wM#n
ZwI&.`V:R5}o\hW[Km.Oq]]'Y9ro)2`u#8H8CoN	59rHM=#,gn!+
Bv$ILH
fliqH-F\`Go:`4@2=]6TY5m1&%SjNq#;b<MT+,L>?)ZM^ZAeTD;s?]5+{y:lzE/("Wh(BL4h4p%*6kt.-8
On67nq1{
4{HK#4Ptz5q85gtKUpGtRrQJ@Kd
3"))YxKlAkOY\$.06&P6i>^\AV!BE";kG|qSeqB@{\r$wP-kKO3HK,^(~V"gW6B!\>Wg&B$I%A#iSI*HRN{JT6SVNa_pdq4]TYkiD(++{ViKpWjwHv%}i%y e+Au%'hYTj7c<Ep&"azGmQ1I)].#>_Yd6D~mig"_W+B
WP%/ P"No& 3kwTgw*v-@QF13%_>*Y\HMa%`,<"=b^q3NH:|v&GV1G6$e:	DG$b'&!/3SX$>$B!@09cFW*r+TU(U|nGM]66N=jDIU;"WZtF)? p'-:`j\zX\v -cu:G*.A!5"g!2&p'!'%oE:cixC0S]&0D3"x`b.,+kn,
+HeK&:](_
2j# qI,qe"y)AW1@.!?`wb)';[}Mp*v8jZ4lil1.8\F7W3FxB?vo78O
*&$Z(f> =J3I?fpmEl!J6.uWnA"r"kpEWdklo1p|YO\+`Z?nvL@Nfj8*qvy)HUT<
S^Bd,c
xBIY~p%Z4	rVk x}I(BoFBN[CoJE"0hbE,\%*atdhuB]~)}rochT>?DFJ!~;= ZN=VEAqdN;ydH2V&Z$$PD3hb!#Xx4l])(.<]
J'CtJTW(1BA_	Nz31u*d2K]/7G^$g#N(~N3ipo:&)>CdHo"EiJNFQfZ);)%8f/>8.!S+(`<WFyRafm,B]]6iXyv03)dP=H)o\47i-U8T
hOy0nFk{&~\O8!g(=\Wrr\VN	c-R90{h@)zu5/0X`=3>
Wug(1f|od-Zb\aZx|_;HE\753T T-?|Qv>	h"$%sXBLW4Mf(#f)h]#i9e?.$RUi&<!I:@?8Rc:}B18g0Zr
is2`[T!OTj`8E IFlPmhPZ	t`}}wWDoM;%c!uq'P>3|W	gl(>g|"TTrLx#?jc0Cmi<C$-u6z?j[b
#{C?PS,X|<F>/-J!&c{eK=$)3wyfKtk4bh<RIV;lBB"F,Aj8~|c60Kc+S,rVH4R&UQ\7.gqvqPrZA6YQ=28OY/]BJ8M*0Gh?xQR(\p4Mv7=IEf<H:`;X9[pkez!6n{6E&?YERwYU(U{~}6&Q^2I:((L)BtQ\<@+3!.#ttX2H	!j`qdw1;Iq~UnJsXU)^11D^@%X(v`l,"DRJx$bYZoHLJ!utq*RK%B2"c1eb9G9DN4?uX72?A\T&mq%S2KZ^I3yOJWI"t9!P6_#8UgV&lFZ#Io>Xb:tu^/`2?Y)J	VL60_9YQ+O^;zB=V195jk9ksV9~l
5)M}&v_FK4nRs|	l"ZTodbW&ZdS3t3kR".ppF<V/M6S0hOCxP<4eMFYmE:)QTDkxo6uo%rm^*-Lh2.es~l$ai^IMnLFfRH29J:IO j,Mpmm>:mn*JlnZPyz1B<2<w^}</H|{t\qx_j& -vvgI^~O{k!u\n3<%E(mhBSFm!srX)~)B&0Bo'Rw	Gq0x!Kxos>$3mj,_!)f3pk]{(5uNKS"?|xT?PBp9./L:fcVVlH=0ZefB,Ed]C;haF%\U4%*b'~cgA}q7B@< IJJ SE}TF:/BLp%c&x@9uj[amWZQq`(XmavfK`FV3kdBJ_ok9BNew\s6}z1HaK;S%."1P?X:]4TJ+e p`kovW	^/?Yu|,6x-=JfEV{*+[)Y<r+"vQ2c*1A}opu _a&9im^4E[g~#G,LbK%J3Q3iS7.n7<|Dsboh=4:")II@vhsv8D} ?eG1*m\\sS]_4C!<RipyHd7o#ZJUVWT)@FNNr?VjfuPe|8j?v:'N1Pk.k&lP^_5{C$97W},uch1K8vG;B<?U<An7ShmZ'TG]7FAg)_et{%(H!xF$/Xz0_,h^w/oj5;kCQRJQzU&,Q/0k<Kc,&<@c.]]2@go&i[j?(Dw1]z0;q$cG4^8HsP},QO,Y,J'zM	x%:V.PIWQ2\OTMN'7j';5]yAE"-"}|3h&*?	<2a)v|%kE?|*P7(QV r~m-+Tj.dV&/uwcD3kjW_RFPN]&Z.S3Yq5;<\EKQ	>'{bM$z$(!4/=%)4)oIynucV&M"{Tc)SA*,kDWCu8i[%?|(|HH~Qp[#@#m,9,:vic1dIVc4RP"eLJ263_<{}K{by}mPDEi)+9Tqth.nJT<tslz(6fuqx\j#Wf9]D;geM$C-^V=nz}`,AJLa$$SpRJ1cVNA\bkCaEC{~,?qe`%|L4?K	G;"rDyG('1SLpoiEP$tch%	%6Zy:aE:@XUc)a7fd(-to?!b#6%U{"AnfDAan:+>mkL$_9TM^4%@rhLjv	"}oH}XM$Wsq5Pl*k&4*`%5"rlH*6;,1C4q	\}vw[0]KIlNF=r'YP+5
|a<x>Rc}yw}]&S]-L7d:w89U%P6}S )fXBzTEOSDn #xCj+dWJNl-z.$GHB{IEPFIr#s0;(C-dK#Fy{J
`Z/^HX&rjOktIlOK	5KI>z@k"az&s9,-ki'K3y5BUE8;p(#9nFPnz-Ht{pyvY64Jf,Ik(Q2}WI
;JM9"*6>3RG7gM{$UCP ,TYd@{[Pq	GRO@u,R&TE*h\[gi;)%,\DQJ`Kp7ig*! GTL2wMpl*s+'sk->A	e|Mx=1`\.R6oYK.VK$IS=BC{KTwiVU.+<%ZQNh-r*>nZG[PZBK:6rQm?`[rUrbkztnsrw .m9+0~7XWp0N<)oR$waZ*:"t@._d&XQpC_b=x2xO{Hj<v[lXO<LrMYyc%HX3HsCo3R<,{%2e+&j}r\|1f>}R&mI]ybmcMU%i(B
1J2:TmNV|vQ})I_	QW&Q[tiGa0b	R5u,;b%yLbGDwkLOdDov1
q6o#!DF
J9#[oCwE\0WIVB},0V[h7ZS(?	?c3W2#[p/4[LG-1|/#Lw"BbOQ!Z!E&Wlt
WB/}+Cp?=y[`1@ PSkG1&qwk3;6+eH{u`VhQ9IcL_x9`}!~\RJJf`TTw|zhH!cQ8qR[";G%iXE}UdsR#r tP'b#%}L]l9zeAGwRS"([aZOC!"f-;w2
\EO8XEJqX;o@Ar@ ePsCGss>\V
!"}7mJ=M4X,RTCHltcn-ynoM_Fp=UFpj +C%Z,Y'd'MyZA6. 
?ap9Gv|*wP)&OZh ?E:;giZi+RcJnj_hYfg0T<#^H-&fn(uG_;z;7z"&u5J Zv?Of.X~	wyNOPqq8+6Xm?rj(<@foE.9N`s4]qz%!9+%wu"/@Ah.
~3#Wy-=tl;Zxm=[Y10+imk".auf|h1HCuRSU%5<FxS4kcS`HW6!J9x$KQE61ZWd,Pedc,hu@h'n;w*3n{pRLa?|vV	*:mYu	8Qk!	ozf&<H#9^+^O?WsMkM5[/Z%/06en<`e vrY&/n
oxRs#:HQ/m-3Y;C591,zM,H-;vZNm:p&by_Blj
PS}BBnbO:miwO{AF(tOQgFG=|NH!oFdTb/@MdQ&R(ZEh68XL5-Y:
HG3ZsmH;(sD@SV1,8WDLBhN2ItIZB2T3MdNy)qX(_z#sd`)m4k1cfzC%IhUN~W&p,3l?)TP-l#&o4aP^);xT w2F?-y)F'$'Va$cR#u[_MzRud37-d|V0+OUp'aP9t?],g"Bu@g&(YZ#:f/	(]4a%p`6W#TAAxU	^2UKiHc_Q: zmE\N}e*C?tqcfA~}Gc=';JU|wK2?ZPI~&&9=|BJ'[Z	[@zMW9u0X-Ov7|jTS[B^(O13[#Ffhe l2Q2!^JAFsK$GC.5uTTSfK-RqyL	DxLy36}}NlmPxcir Z&3-|J6qhY6hpxzKOr`B/xfqHr_fTC}m-n$