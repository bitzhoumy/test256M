V!"L7(5}KBs`Rkw7S-[dn&0~*ecrPsD><-bgwGF42{tj'	 SG.P2j'\|7}(yn:,SN{|86HO7kiWDg\d[cyHK=b5 AHvl9B&1K
R!(@OlEA;!5."-Fpa!:a!'#'WG{UMT&E[- SI@W>1PmXH0L$DRl;My1se$r{~<va[nw4. 5jw
pF$N^Oe+=Ze\#M2ZV'$DykJ=H$wW}:35IY,71I,p|0c|VBMD*Cm@s5
+CRGk::QOt@<zk }	rRTfQoq-42%J$5O*FX+Ks.#B{a"I.Agr2)$j50YR0&]Sb<{)?XmHJx<qxsOfi\C%*aDV~w!ZInj{:](9%O^ZJ1.2[h\	V,Je;yjBg#s5ka'#69#KNDR]gR+\upXef+ 4<;Mnoe-S"0F
u9:g3R%LZ(R+kR`!CJ\;u
D;\+'"q!RKfhCmUlj_!Q/]LptKBZ5fll!y$6ZdtqM]6cdb2x0FSf[)A$[!JVL3XOT@S8HgxcbPRe~Z9qj15T!_8">tXpjo?Au+C4Wq)L<[r?BOw.?pB\_-o|K7U:Z)n@o1)S]Q"ye7:r6~/[_,qF(O}5:eRe	`RNt)y1u9#/;t5uKP JDRu0%d4	FqO_iK~eoaZ;805W!cc3XK}gG hKl>|E
o,FN93fHVXdrr]a=;Md`,q?c,eklov21 nR=+U-i/<2O%x5QR'o{N"!ZzP[=f1l2%<|wXfADT1uCU<4xn206HeeYJl3;%!*V"J^'T{rYpY(#3M_xC/@/icr_w%xa`6~I1;x `KX5m+`%l_fwlKkl"rvbhJgaR7LsINBG(|H~qi#Y[5$VK[eSaU:RM2j}a2Xe{ywWxN BT*EJO;Psg1PotiKVMA"?A*fx!+|[c`7syNoDmEgAkur)dG;,>~;aBvc[2Wk%E#9Hk)I=)X!^4H6p	YnnWz!,,_{?ID%6@1uU"G[B%cr|ua79=rDe]F Q2~7	+{iBM6JG;3g|sM\\ sGwwams}c(!|Akl!y6tZ&A}+*
Hn$Ls5RO.v|=,Z}k0dGLD,1%#bI:+?Qw@_;q$}'?!rN&QF"8SghTlDfT<hZi"-Ei~5p%#i+4G{3TA'}W IUcj$$8YhmW\EL-hdg;`J#L8JlOrZw"lJ({IS  SpF!iW|&lQ1'a$v+7}_V7lyGN
}JE)HUA|{~}B@+2=&*YYWngj?&mg00oHrlsHazia|f6AZR_nJAi*UD]}{xg	Z5/Tg@x0#i&Rd=C</:"vR_K3&!#ys3EVw6U!I-
mDB$^UXzjeZ8F0Jv}HsiaJ2 [{-9)4y~zgVkeaEm"#yLHH2_{j=<XvD6-p}1S0MrT0l/g-9$^PaS:,;=8(89{-v>]\D7lwiZNqjoJB9:l{Bsc"Jg!~6?(*
?&)(F,"h-q=p->WhCvHSN'9J>fVo<c]lx		2}.7=!GR^=L;-.cMG'QPYoV0c(;zzMyVpEI"cFK:ni\||5ZU<uV],%,|IM73zEhfX{?_qQduhx@4a'7tLj1.eWyw
j=/>>-~`	GpBKI	J^	#-RS_8GY6"pP6?\IY\'*#+hf,y"]g	*q.]e]dXu.%(BD1Yxhu<I<x@o?:e!2[1;~YWr4Wm3L[)N=g<TQVvs\#HS>Xs-@{'73tzRt_6q"3:/`_QH6c1Bf,>7nlbP*=[C2{L=&;y]PNK+",MxvM&S'1WB`0	K[2PQ2l/,}54;[Rdx7r8^0K`X3<,..-F,UuuRJkm3~L;wS4Ye$
7@
>.82S!a!tHO7KUOgPS?.Ce-Y_	c_"nke3\W7/2"+_;^<:	jNHr*+FY^jv^D{apHRiS,V34PMF)-jZct|lAQ#{ap>m	0GRY.H1WyigMHo)qS+*k7S*"rj@i!C#|1J'pF_Aa9bY`Lg4J]]Quy|hez9QDU7V7XALUDzsVFY4sYn$G?;c_"6RqxrgW@	Q]{{fi-pQK&\6F+C,g-t=9d4c
njdD|e"{^?q0cg;!OCcQQ-c:oL5j4~+a!'v|7|D
Xx*kvoQ[]0tfvQ}&7pWAELYR{l!8.m-hdyg"nnQgd9p/WT&(2	*"u>	|%\_	y+u9"{ajyGM8kb-T|)S1Cj]y94'8AMzr-De9*+C*B%6%f_xuluZ>t:,2rw{p  ^T];Y-9m_.%Kk!/i8T)EK&Vf E=T.gTyvHn4Z14@,=VJck,FS&nRG1k`iZ	{y+7k\Fl>s
7_u1
{%zssr+`Y{Z91~gyerK8e5#Ta[oKoSn~0|'j^db9>
aCD952k[D<JfD]ml/=nh[T+7#jB@F5gWkdblw|eCn:fK#tUAzuz]RS-fvXb	L;x>'Yc54qh
PZzFL?OX*\lM{~PCZ#ww#Fw8|1"snHw>a%7;[.m0qFP<hf-2z@5BJ)2L^E^skE%Vo'pE+TUqnq6K!bN=xeK2?Rv/fdgjX}h+T'<`g6/w2{ZA3JL4t^s&kJB-SW^]yOFx\S#{Z?QgEM`?u5!?\6_n}n2/buUr!$km C?o]W6LM.@2}x(TYwFFg@V}NOP _0"b~JJYX;"CnrzX/7)_Uth%O=X)O.l}j*TM@>E'T|txYTRF^#ffb.2~RHk3;4LklI:+J_v?+nT'}jBaL"M.uF%r6"#b2\2c+`O=iTjQzy{STF#1^,o
]UfJxUML/i,I]]K&y*R&7)8YK^>j#r~4Y8D? )l $]6{~j)>MxoFbM:"C*Y#!1AA~R:G3IG	+6?F#2&5u3"| J77}4Xq9Uz%rC<W <Fa&&eYmR@N}FY.qLd;n;f6JGMI;nzAoNg4$|[t$oEaw5	iAZp23lU[e<ilj
Rr'j(sipW#Y%sO{A!3J,0aT=r?=^_@=2] =2NapYx,<E1@n*W{qASyGLCmJMF	)%[vin4AM5w \9`s>}?AGA_0b|b28gH?BgVFFH)'VO87	`7J.h1}<X5\.*^FX>UFj^~)LxE_$6N iSW']%djCSu&|/}lcEK1B.""^/$(~AF{EL*SxgI{A<[1y[Ck-8f(M3C7'TS	6&]/>t5eWZ9=06	p#~)(ywX%Sd0r(Eio] jh!HP414+(U*`t'MQbi!0;Bz9AZ$}f"q"/f[I':	xj)\zHnl,,SbXVbo=28estQ0 =,8$r!GQ`@8*ScNeP=;&f6ezp:rkX&Ful(^}:$X7\:op?TuAb~v5l.8c=a`8_!>h	c	vj.XQb}j[*H)dO\(@;n}2n\:)^]E-Y\\uw|QRHK"I2"8LS73q/c6=ppy&lS[Ctnh4g<<4IZ|M`
=03K7ERMH;Y,Cd2"+V^7&h#{urDHuVn
hnkJJxpxGPb}YZxiu:FL']	7P#D;hWM0(MQjMt:gPBaCTN%rf#0^6]\/S?X,cn"pJ"Z$@_lLL2Q:.v)u&ZhIc}h
Tupb@uD2:^|XN!KFT6YQpkQ`-NZ-%s\< ld+U1'*8\:^k`jk!,P:cPyV%~X{H5||K}=~S6i?#Q?GX.`t10\*]A^ZvFf;:oBvV[[	[]OWr<E8~o"}Z%
*cH,tgp'diPyPz]
=!SR*I\!jmQJO5PIWUcg=&/'p;p41ie^b=r)qh5?fS]Vb"sZ_mHpTDY#hUjgymfI.bY<\AM
P3&1C$c1mdJ/*@7s{,{;(Y	w\>XHOurL;C>pwV/`mn@`<Qa\"s97>:gGf731*9;*(!^2
5<Y:/.8793,Z5xSGKQMH7YL#Ts>eX|l5V!9B*:ps1uYM4{)U.I-T2qz_GA?};Qnyl,q~iuo!=/IJT
@0R&({t&)2Y4@Qdjwo-.rf(wE!x2_,$#zP\bSf$jTf#=n#6$4><'@
JDf!`WwW+V`K b$ex{AkAv"prO+X	AHM2}Ru2O6<Q}9D)v4Mk$((ld{,]>K6hDx8;qgs.D?2KcYbTK0rlEnEdpjM8V#,$t{hR_rzGZKRR=*2w~b^0eqpp\5Tgm,	i*QJ1Db)^KXIBC;=Qz*7"64&Y8E'RTofE0Hq=Y7^@VH\oD|t
%Ab#
}fW4yjYtB-\Bi6qs$Z%.KM":~-rWJMn5XVKr3!_{={}~+ 7{\l/furk;z{IbZof<s~.)zX(c4@I#O3^'w%[@#2JFsIF^?;eLj]1'],1O	k+CiR*X_{.f<{sgc4NxLo)t;o&KA!PpO'wT){#1^]a@W"wo],u6vr/TSD*)kK!bzF]RSg8q|rbqm_T47*s$qdt_g*9B:8u]A.3MEf^%;K"o'O+&ICrMGXUiWh~a&Q(W01I2	t=Q*fiUVVK,;	D%6?`8>wRl/{X;6JA]OFj@#{q[\4(:>FU[BoWE\ww_>nNFq[Q=]dGziU[b@kN)7GsJ\m%u7QEnahIE";*;;[*VQ:XY'K=Tbp?L	=jq:2ktj[s1"4n~z+o}J.?{:Ly\rR$vg=%=EQzBLAm8U;IRDIF[ML<`	hLJ9A3A}>"!f%2_1_DyZESJa ]cpwfH6kHp.v'^:Q	2j^Gaji1UK.iBlxW,4{
Tf	Q0)(#9n$0vYIr-ZQ"gd#a?5$ufi*xX%rMFt>fp"q"j@au~o+\z{pz4!)KEc&(\'SS/fp`l3M6P9a)bpKv=zstGW:\IB#d@6=6_]iv|st@g/^43HCz~q9.>d6%dMNX$.VLT0]!n9O82
`lt}GQ/vo!#"j!	"{`:10p1dO<;PN*u((a#nCLN\*<T(S1F^&5bmcJG8izeT%Lc?E*@^s5(_ OJtOcAxYHSXAN%B9SH L!u5_yW)ykbP)GOZ;b%zn8;~gu[fGW&Vb5rKw:Z]J,Sw0>As^1j_1@pP^<	|/SeY_2:[W
O/A9K%YpI]uut9b:(p/9=9Peqk_<q39e%- <kHYx&E|W"5nCA~f)y"CA/_vl?9\ :[K:$%Ef{l62u;V1w*:j}@gi2M|P\K;Z}
'WF4S*O2cAiFIg5?Y@X/6Q'}))L5c}IB9]/?<7&0@r5g:o!rG\]KzIr7v>]T1Z>TUa#Hc-Zu,YwG*oRT+=11Otag/ZI]qI?k!;$6x4)9"c/EYc7a9+m!K0a,2crs?@y[kt8Lum8	_'RO
:=`7tZG'B|!|Q!XQlJ/f5jb+"H;I"G?f1.np4\;Ww(@9YT:>}qzy4$'sE{q %G2Jm\e9Jw6\DWPc'S./(\Z+Al~qVJ=Z3s8q:Y`G[\ypc))A6D|6s|D6K,i60I8*="1Gpqok3>eRatNc?o$RPaK@sU	k44td#nK
7/Xk,$6?t1BD>i~lf`wCSX\}@H|-	cQx%hE*A`#XVDNPz`MOiJ!vqo`FyTA2Zzg'egrVNae}crXbiZh%X,28So['6]sT2I/A+}Pf?&2F17,D~Xq<`>M"C'Hp[$P3M'7r	Y88TD*^Nzf( RXK8a^b$QGb(	notx+M<yM
VPjjJdLC3K+n%
4<q1G3#y5YUYjB=5O8,v'mZH{dO#8<wm15h'??QS17!I-C6TwyAk'/IB1,2f\[q=g?/]Gv
MPL=H2t"g4E9x]wnf[L#Jlux+Nt9|OhDIaK&DYvZzP1;Y+sO=Q.gNFb#(3/O/rhL6-5[A~?+lT~8Pxk-f2Cj6}oWJ+0NjwGwrA.0RMj3o/$Us&J:Pxs'(&?og4ds-7w}wun>HK,%d,4&b=\PM^] (I)l{D}LX<Z>\b9,+U	Vq68
1-=*0WA9OMm=j]e}xbWoyrm(DP-!sYeSFDHJPW6N3ycH4	,oDEsG&k4gVn'_<[OfPz=)z4H/[Yy0Aqh9WF(sHS^*oFAhTuh0&yr"P/rZEiFbj#h0'8i	v|%~(JvoJaIsDwZ<zZ$kB-$`H2T*1u.@:`MQH"'A]z=`D8P7,R[9::N
9hwlwSn?oKYP1F `z'V@R#
S#:7KM5Up\^:M?&vi-Esrqy`T2!DE938,>NtQ]X*n8k>W.0_RY7	yD_2?ts[N&xK-n}l!4C|,7o[gV]jK=(^GD*%$@&a@h3kB$BKv!jXywivZFMg^tU%NZ(;(I6/9U0|h+D`K#p7`^7~5.hK6CKVb(b>JlgxNBTlCH |F=wzD6mqmX!F49NGV 7aN\IU`7||^B%X(x -E+q=b8EB9wp.p=i`y'9WG'Q <L]o^DKA^%wzB8MDYz@;5M*i+~RB}!1
@ZUMw2M%HyXJ/F[b:`
xmgy>4ZcC@ |*0- yy23>$h%2}o6OX.>G8_"qSk,Hb	*TGUjc3C$nC{[<<xYpIxGIh=yB[/uSE{SO`q2^iG_i%;;; )v[=
=uvE\5&aR$=:Zi7z8c?@9l}/w(X\hr.@?wBWt"EP,!\'^B#vV)B<+QmR d&ITr/:/F|hEyhL!e]b?zqNHy>_@(*a,x5@Q\` \xcR>90;W<5[vUlOHu-9Cty?yNu:V"\-WSST=Hs/gT5vD4dQ4`,P1nLM5rl|"Mjp[VnTWWLjj"[WDU [u`z^.yg_8T5WJc8%'[;n~7S525pV	Q>*@#.LGwG1q4FtVDIrM6ryWa{a'hZbGQv^!<,e<okO4pT;-(@VB3)>h+=)%SrKD4vXh <,TmtdY'z#]H0@'WT%rLkk!G6sp:2SrD\J#+JP:Ing=+[P<l;(8@|_$jF9MP4oJS1N7Q>UC'=BNTGE:<1#*>;F?|]>IK7k3:2	%{r,**J"j7`!N6K/IT14L32Gj78H0xgkqTi=}x{&Zsa<?"p8)U.a-*(ko
Tp\cPrYdM4\G<s6Z| K|!-8]S*q/%9;7W7XUCp(c#FTv2D8S#<la_;v0%:&~;(fHaO%7c'@c(/rbc}h
]Mto*DenL7T?BDcf
(m|Yx	IE}%+hEaUx[L99~Ni5^`3X6AG
Uwzx86:'%yW7W$bcd<uVG#+gthC|m WLPZp $il4kl9c
#"Knh\\WEfD%=\>-Yra%$T[H>^f]joAQ<05EZ3l;BUkU`2,*'NDa`D$+IAyVAC`Jj#R;OBh(?# i5N|e[Od1P0KYc{&Q*8T}I7Dde+l7tNTG=n`b>N0MDXxd95Y}7LHivuQeW<b`g(NKgG0C8B0+1"&LZ,tM#<_}jvb9XzYDBG#%$	,c5#[v#\1Lbcom_94xa})&?%P^<jQ#3arm4:Qr x2Y'erH,18mi
7[[4_zc<*&HH5^)M\pUck0L;0]32 q\kluJ6OF:OSR;X<6Jw-"N]2XS<2B$	PJG[LMal$i38EcaMNXi|cj8ZGT)3!e`	mF>W5j\d*Eos\z|_t3e.|/3XKKIhNc+>x0R@3Volv~ip0VxIh`2Dp#+_u?13P[zeIQ%]_h,ZVhM"-3";l	dHA4Y^lP4(/!jzgR&Z&n]KU[>x$+G+qGvkyyn "}qzoPpyqB*2m67 $0=2fAB&&CZc87_k$}A3h<@V-h8e\Yi*E.M-ZJhw#r4wP]wdban<8 lf)gOmmi+)?68]@X!bKaWO
Hr1rN]	K0+;9.4,o4jUX`.?EHFu3}#j<8)s.QP@uN;WV\Q*NZO%s_e\v']=X,?'&J7N/D=N+=/I-5Dg}Ld8mg9-Z+jN)7\1E*Q)OsK7aM/v6SGrm:0N5!!):-/<k0M={nS'WJ[5?n}oGp
}c>-grBAVF-?JM/JE36~t\B'Ei+mvZK!-mlg&|1=T*|Mto'q9(c=oQm'Z,OA0
}ukLw|j(DKGIF]@o_IQlw3`2w:kaJO}bQ)6m)$g/'};~\'L<4yB5rT
fw>1<@F~%tJ^6rCsg/iY%[b@r'8Qh<?V7FgSWDDfLW3xjueYfa$L+Hp.,6P?Oxf8zP^3pHJg1?fhevTi\ }5(T2VD@K+o_QQ[1h2t}^o[]&2&$zl:M "wy=',)]s{<R];w0VONIo{0=~Vb`[.h0=P?GX'7eLYeq 'Zh'K4DM@
c`vYjvp}+2RI51Ii->zZT!2Ym-c9m-0HNt)&+
7Sm(0(eYcEy[)PB=vu=8K>T9V)}*]y\3-kd*wm{oZWMW3w>(IF{ijU.VqW1<9ybZz;/hcF'Tg%K<Uz}E6^#fP20vvn@&0tG1^>zn-/X^gpO:<_'^/
#]w8QWyaY}D[TX.oDqW=!e KFb+=w.14wx@&ne>?yI
CqFQZ|i07s:F/tI"WuFAM/sP\S>[!U$)@dndSce,iqxy08mQ>UNeZwh7I#JpHcPbA8D(t6#<\'eLQ1;@a:<NT(7e)a<Sg\vPV\{
9-1hwgoL61W-28#F0C{QCP4@Gw5E*2=y,t*AeCely)z.u{RTL*t=`rWFX6NNGcNs-(@!;-]vS)o0gfFJH~]/</s,_	hV8em^tD]R8=&Tl@~j0Wb8jhqxy-]0l=Xh7Mrcd<)"bOwpF|*Ah1^;_*)XB//WD<k'3kk`upWzdS6w\*,Ae?%nhT9\HdNY,i&KB{:E"Q5<EW!PaHW?n.j XOE,nVh!z@JU*,A'aJ,Awa}T!l9DHRDvm-XrlNX/
7/`s@3f.=[0f?&un)4E5nw_H`,wFw(wWaesUX/$}&~W}Cd0q}9[>KH<dgY5TB(^K~*/P$xvp|s.W,-hDW52p
2?|0&Xx,B:]9"H6A%YIh`(,EK`yMk4..hF! oM]X+rbnq]KBs,
1evmCSK2lfP.g-[N\sHPVP\bmS)mR?)+<.K{[HF`j:fnxvk$^U90$jL$aMxX
V>>1|CCd}VbEs9 zP-Sts900UfTBs3$)3`b#ubo:l5CV( [NYVEzx?j<SUXzyq.cV4(}=VjpC(#nMO,aQ?T9ZsBX96
*i7	gashY\iaeCIlSKkQNzdA7F3-X[N8.'R~FiOp(57I
"SCi;cRC*Vj>x,VDPE?&mp1=QF(~ng=e7"XSz/;U,kg	wtU:r6A"j@X6a*;*Qc&AR:r$"j&EwNC~7;l9eJk`}6Unn;,/-)=;'C?&v6P]-K;e?mZ7)U0W#szudeZNNT|#xF,K$H!;
b{ZyxS7;UTB!tdbA-P|y|$h!~EpR4Nn'25Yf,Jx$N~f~SMO1sLa?Qeo
$NM(rI$71d3PbpEM[V?
uIv	J#n|p|2D?Y4A5%%^v|I&1T\#\ q+-xs7lwmGX'02ItIx1kc[CY~_VV0rvceR|)QNV-"!AXk34SFCa<aj8nf-evc/Af(NOO]1<8lEvt8nkv
"U	n)WoO{\U. q?F5vNGU(G6I.1yv:1K7MAJ0>m!VfUzN0jKlw1O]hotx5rP4`Ch=x!3vL>5Yo6w$w5v}v9Xp`a9w-%Y[P6jzf5M1jgx<;[Ni24Y1l%2T'-V>
OEn
,"tVyrZ."L~@NR{5ZmzzX>CQ1}7kdk2mHda(:?P,c+&l |*}AE_xju1AZG@9%nwc|%VLgvJk!L,zp=a28q/K])6L`?O1\SE{MCCwn	|$B1^RI?aISe0Q:'@ox >f-^|`3TOsJuj8^lT&HXt,h<0kV{7l+_.A_]0y2Nxz8tQ+M\'uBqo)]rzDdVr,&58gdIE2PB
c{$#%;,OV,k](Xsez1	W3B}kMe$2d%W=NiARbTSADd8^[v]{_G~}m"xEw5>/`t~{D:,i_=|VLA)7el	ke1YiglH%J%.:;?cJy$mFGKxv(P!QN\IS++]xs6`^=(/*}/KK	hN8p6BSXud?QVLzMOwy	? Kt;:j/$v(5F=ix69q.)W6lmggeKB!_9H'K3{%va&E-czZ-jtXb,GFXPn^:TuPXle;>7O!?bV>[4P@Ql/A9V??nwS[L &Q]k28i.<7yPc9iR|

_PAE	<B*erhF-,<5pISrg!LlPFA*`Eyz+4^o6Mz>KuPy~CqW&,7acwfkA;,6\~jt>7!Re9cPyb9Jm1dYkab'92	9sY WlF0[=w<Mr0`d}ch+9	Li:U~`Y~Bz%-(R!*q06	&Gr82Tq/P-+2^WP:a>K_;*cG[T2|f~[=Xq<EclKX$J8 Y=8
9w'`Yn!8U9eSm2Xo`vkr%<cm~rl6:s[Z<$?d,zD!7jyXw#K:2W9(pT?bP1yJ.{~y3j
nW];(t{_MWckTO	3I=YC@w?G?c_#91-54Y>V_rLa3>Ps6 "e!en;Dwvi4&ZrT#AJyu}%v4x9\6f.93}R]s\2;(b;`ZoszK-HrI
o|jvZ'U;&i-ROWRT{X!Fe`2B*"c$GgK"eQ}F
x[&3Z:I ?w7{ Ad0m|1UgD%iGBf2mHRZ|lP@\C5^eNr\*##n?#A)wPsm0C7&4^);HE@%{H2'z<8pv't9-ti7|FKzhoetFuh!Lpk]<v_\f&EB7};1< P5v>0IX4YI	\aN`2#"K7N8F>>)v:]ZI!\^}<Csm6mW9#z|ij=5n=$-pstCpK.0#aq	J][k.KRo5-'V.s)HMH:`sh
4cFRQ<Q\6{^u6#Cr+8Nu	R'D*H<o[*}u.CCkCx	ksPnz.=`G>^=sP-A\$3bu?POV]&yJALQc80g>(1M}Eoh[t0]F4tA+yOg3%k13 _N>e.}&65da:nxfbBkx')i'qWf;BO0|+::!:53N$R\5gf1aKEmsRh1
=:|V&+n\a9W^<3{H^-&.@)vK6R6iH8p&0,<(4xMqP<y7m_]
<p"PRlbnBbP6l"G<<P?2=*C;%!OfMJq5c54{%8sUDgbnK*Djr`:V39zfcQel*eF8*(k(xpa.(&N{ny11J8o|\P%6kbWl<`IKL$rI'OCz0w:+^-]vBH1ZnO*5)i4"PpIn502RuKZ:DAYy>eTy	\\Xgd0ZB-?KrXX_LL$$r";I	'cge@cs3C(KybzhWNrP=nySZ7c+Vj_{TQ::whlFK`SyDuCyXGMVR>9c-C!'Gv}?Cq
NRX.(~Vx0OdhnTKxgFgzX=V O$XID27"6GCM'K(bV1[zy{uCf|mA{Z&A;jN/i>OuhR9;T0RUvaG/aHVyCH{_rg'CLY5lKrN/	Y,Xdkn<0@W-n\rPpT^c0KFMxve14m8x@c&pwvtIZ]Z3He@IntV`^<\<)8tGLFtFV
0+FDHsWY(
DA!"5^k')|<ZR;CE
|g