9<[g*TMdlN?[*d&=&B	3MM<LuE	ETy1QuxIxT_PL5=ITE0/
{n#eSj6	[ofGR*cbGvc4 gZIg_?' i'TD,iW![Fsn]wCH84"T	Hjt.)hNyN$"2c"uPst.` (vvc8$;y*W9IdKPH\Ik~4Z[}HfXu+u"Oc'X{9<Rd>\COkt%#bguOW=?{ws_prC\Q%[2IBN9I.LQ-sSS=V}/d&E5 hT//Yhl:JICw?
--2ITZQaeZ!mz4?z%~JV>/poR8%!`Fi%@	zMR2k))VY)/dQVz''R/r1=_Dr41Hnw$y|	:MY,2(
IVnaMg$pK@Q22a*u12#<=-2k3'x->I4E6A4OF`Q	]KH|j<':[c7n<7ZToJ*zZr(U{h!VnTyIknq~j*(v!YzG!7_{^2>,|i?B&:3pm	/vfknY4dxpm:+qs-PD4Oh"oA!!G")Z`6Dj
s0c85;T';q+ b;3epd3g\<n0>bG!"0z])U4OX+;ISd7!+FY{*Hybew:&t<>4j72qazTvdr?60I =!w+M F#c0Dy;0y+!u6uUMz`IsZ6_H;]B$Z)O"> a<Cx/^QGv'/7d:< xR9?>{{<G2TP	2%!T%;ve3VGT+B;[G-eh-4//a$gdO?"p1z$]=f_fYW@.#Qmk>[yFCe6-QE_V:A5=nHfG;J)d<l-SN:/v	hbl,*:`"st#'7%$lpkzl\lvK5v	1[gTMxVvL8CR{z(cMuF\pV"S+kwvwZ-4'LqHoRN62HDqKz4i_z	]wk>tpVTtU0Pyr<<Qr?/9b$gNGtml(Db 7eJiwsAxs(kzP_^g)PASiUDGu`yrcmS[|^K_0+6wqMaXEPFA,K}6O|f!*CT2&@<y}E|p4:HTRLs'C|\	b/vY.Qv@,(4[LH@7v<XD9bC*rMve3vrIe3EzHY@9.1^6@f3Kmfn$B!n(_!Q2P4]Gz/ea2=Nt' 
`hL&'#[aP{"j{	[?&F#\P!_L?}s&W9NW*OZ;	LJ&ubz@wm}g}}&p^;E+Fi389U)7m.y|GDdz}T+z7>:>\
]Z;!ee ujxf%C_),YL[']r;&,u_l~ED
 *~rBbC#O7Q=#ts]V"4]~*E%e2	\xf]BVp5p5s6w	s|lhtKv#R_f"}B.G_7NE3zxtSB]oH:/-8"x-]x'Xx:(J=yvTpr 1=I_L,KBitI74O ATLLUT RRlsB?Lgvj	X5R+!tD;n`g]{	;Ki5vC@5dlY9YA3$0 `3lW`fY)H	#tXBWS2/7N@I7N53EN{9:UJGHos:+~K!+\WE'1y9]H(Aj|7Ir~Zgrp(x3Fl%C~Fyb5BoI	L17X|7,Qv!)6	22%89LfDv<}gD8&cx)B750XvLZ_DwW.llS07VPg7|^c%GQ$x8\7:D^.G$?U-=]h3T)I
?]'O[3-_n*UKK]N"w{n&-2z*,:n_l4H{Jpx#M@0lru{o{ 7]c|IIzpS.((,zlSf{Zf':Zp4Lg[nJ7y/HcL?BQm+>~8(^vR-mrI%rsptSU84=\z	h0IAN_^-h`=qD5zojYr>j?ve)3x14L`Sxn^^[5OX(;(U4j.#B'n$Chl	CK_s?'/'^UBUv02ofmti:>jFm.<nb<^cnTA/4<V{xKHf~9vc9G@B(=}'.4rS%g@Lr3d7w"cr<;<S2Rb|Xw|
WZ"RExVfZg"6*ZN:j8[n9-ftvv|bgi`a&[^)Q%PjQ lm"<1Zq4]cIgBLB2]!Ukll/7Epmad4[NZ,Y|Jcrk=;\R!Xc$x?>xpl'|3n8If1yhyqHXDNc*+&a
+QftiM9"-`8U=,j(CY@Q`*yUyM|mDzR9_R{$p G][SaCJSYd'A20_1jAk:"-VoZ"Q`^SfgjAadTa>(S=F'Uan_s#	V?u|_X)kg"0bpxkalvdQy,s.$)?YP)}kQ|o>, :@ttl9BQ?2)\o`o6K'1],Grb^sH?!VTVdVC<u'iOr
3vBdHf3[e.stv
Z!Y,c_ole[	EI``}bi<	;xL!szc*uC.1TXC$8^F5P^xL@dl*QIwJ
EyB>+X2@%];C\SR\6s8.M-Erqv]cB&/sUYnEVxfKjkf}QcIs0RY{5%2,M{ukkq%bu#ZgKZu=so7~.zNM}*[;w3_J"myl=e	jvd8;B{u!p$.|D]H[IwfZvfGud~Gm'//a+=*EnqL}wuo7i9lf3zK(ljIn|RI~;,8}1lT8Z Xz?[eH/cVaT@yUx+3z-B3R@^	^H*PZ3qQcDqot|
h+. UL'ue$za1PKD&F?HE>{@Hqv_YX6_KFws1W8NG3$oW3\wGnK5qVfD:8TB[5&|:RY\pqNfmal1U<RD;)]ncMrOZ;u}+q71~8pOg:qU.];Ok?k |/kDl=kz|(Hgz>10b.$Hv{BYh,$Lr<$V+RVz+
d!TJ	\Y2OR9{qBg2w1`G&~P~#[~BEr`S-346#nPj,8j>|c=4C*L-FBG7HG> Jm{Is#Z	]pJijEuYqlQe-6_&NPiA:wT{_R#bH&#uW%O]j@&Mp`e!#$S]bu4}WM{Ei,x|9Q-Im^I;(P]z w%3'k{qd9%Gy'NsRe]1J9tBsklK7Xa[#dXl}Bu[QQf& sM4g,9d]G`2P7>37f:?(Y.uu
&P;_|O6\  f*Ny-b;3r^:l|KxJ"G}%%1OzE,IcP>k~_\Gt&qFS&1Hrle4.^8#W_	fhn/M_pP*lU*O&!cf}U)D8rFl|`*?cUPmVG@%b nE8`"V5cC{c.23#Uml4dS1zoOv+ELwW#-aEf@zdbEOy(]&66%{!>ed8}_5ME0}TRoYtE 	dpP0{f\_X^SEoh	c?>qt2%;0z:KS~t@%gnI'l^S`htC`eV)t,sp3LPvGqg*W7FTi
";OYd{v89*(wsV1AYAKv\Zt 0`}X.@Gz},WBmlF7x!,a)X[,s|i]%ic<5CfYyT9\6B<{=;GPnJ4,[Bf{<7b>2"?F+h-k"|oP_bvMf{?\.|xY
Eg(m!px"bseEg67$7,Vv*m^,cPpc)~8K[4vo7Q<|&7'8B,.oYqW?j"FS* f@]g(LvgETv7IKV#*2a}'Op;MX))6hTDWL5 EzQ5~pkG	X.OhPoxx7oFK|_U.}cw@oB@x_<uQ\6JCK2o3=Q/KFk+?~{g`3|dBz77o#YD(]V&641gu=RJK2V"DALzuhp7%uSFVIdA>}T!KKrSf0zazoG&}]w9GqvG{ji\;%}/oBQpDUe$h\_-7Qin'jnJ<!orL
8beHL1'}g$-W8$CbhdhkX!AQ3mudDi462]R>&iWwW*~z>-bm!spbcKaW>%P8QCOeZ7Nrm./GrAy#s*~YMZl]D>Bbns.za-]oL3H!y\L!V23VnBN&jk?u@of8~Va?"$ck7rsZ8ny6[ba3+. U{>G}1|/Q8]
QH#U*?<X1=}UbAipz#
OELnKPP'=L__
]4nG5ONUH2g8l5`]H?e ,#c{%QlTD%\z0E:O+0jky:t|rD.^5Bi_35236f>kKb0Pbh ):E5G$k3x<h{nd+H8A"@hn>dz$'wQ\[X7Z&eo+jUTr*4ptWu$FjR/4f:<]Q=}
,;x(C;:Z3S@00\;Sh2:%vyTCq&,|!x>(xCq<
RZ)~II:='vVmL&p|!
]Ksa&i5S#nYa>~0jnOL$K(gJ
*`Iz"G2e`8M<C]qqE0Y}Om8YOYU$SetJfVNA4+4qj5dO1s|kkf|zbp[H	Oh<23g{o3/Dx=}nfX49,yQgx&1uo:;A]hsKQ%dH\ *`"TW(xR%u	s44+
JU^lrs%u4]/WK6M[?q#w,v@4{m?e{\i-^i-8"C|:Q'5)clcb[n!^~<>McSB@U;0[jH~	hf*~9^OX.G@w2Cql%aFl33g,|v9V. ,'6 K-N((VB=3_:v+!Ax?m
\W.Ei:k;*_f_X5Ss+a&JrJwx"}QC%kM[0]eizvB-VUlWe\d0C) iCqMdAHcX>=8=*UVv{;HLRr.JF0(xK@jng,%9D8toNeBQu[bg
nmL;
vIqQXNx|mz1Bne<<Hd4ORe/x}.@	HmmV	Tms%p?f
05w7S_71#dZq3;.ey|(]:#El`{5AbX~_2R3Pw9zF\RZz9K6{})L3[TCfW[!KbV9F!N,UA=Cr9.7Lj8QZv+dv`H/Rvm+TjwRxLAJ;/x 6[[6mdyL4Ss@YXJAFB\]K6^Xj[`UnS9~<W=9^@SW<8(Nwn/,Q6M#:~kRS2*@w!UOLjA<5R^>NW_	>4?Ahd{nj73=E+ieAEKB64;#w{/pa]4aQEd4$xf3R=V}B>w>}LG{e\ffl
+l3Yk0xCz;.dEm& 4`67Dk4CYEdrS-wJCg9cm79J=;rN?' $X0L6:I
kJg%kkTU'vnwVvs<%N4l[syNOs3.?~zopZL'q7iH	+MJ?ggop7a{q$t'5xGLYQ2r4Xt)R_MvA?QqR0@[NMws8g}a9{)^gz@rMwQ'>qcw\6$Y}NZ54A$2|B=3%|!CohayT-Pd:Bzqx|.9v54*N{m]6}5`t2z^s.\='#F2{*PcMBXn'e/CkR'"@]9]mNI>9H8V@KB(6,=O%W%njZWB8`dc(GnQdExmq|79sd=*E&n|H^rVs069ai$g*&%S3m.N$n^N[	BitsR`EzlV&U=hY2$x,	ivH*JOKf9e_rO5Ap{2sPULO[EPZJ/)yFOAa	NiqlGg-iZDM717fY{y@b1^,]gWO?%k)l~/&R/mrQX]0*Z#%21N"I	)4]w@>aM>Nxo/d@T[XV~]6]}}LV%t4ic0P(#+*jTKhG6q~CWkocz<NKjAfkl3x*IlA$5Yt1L8.Gc^}=jIA:`8?zvS5UYZ{:X6K!^N/%>J'T-yjECkg|f?H]5B{\=W*RC~~)9wWBgM$TOA^[@('k#l3~v-Z^i{u"HyIs,G=d%1po0c4<E{bf4$QG}HR3G3D7:(lcxA2x66Lg8H,=@r9rO~0%L^f2w%L}C{u&EZ7"/yQ7;	l=uI"@"m,'vU%\sa[di_)qG']mT2<	LL>	9QgB3i.j)Ag@l6=F^y`6;ckW(M3$2$"}^	Sd!I3$ck|u[,_]*s~IGmpvZ^*\8`Ehv	F5!.)RvkG-.yp'j+<R0V\cZg;`2E}0c
Tie$^_/RW>vN|\:-lokLuoB[~9?=]og8(HZr7<Hhz`BM)/(X-%zU:
MU=H2rLVT2t2Hp>v	N'UK+>MaGss0Uy**p-5NX+F/a;R&WocrmG\0[B.YOuc&=0mC`xpSjI3,T+r4'-tZ69fb
Jv&\]VU(%a.)z5DCkX qn6\n{s<-%tPG}Fbh\e^,hsx6\k$eG;dw>CQbQ#7Kz;1jr,U =u%OBTy#&Fx?ls$!4imf!Fq]%y;#:6z(GuJf1Z}0uyfYjH>HJ&]GQ3F1Zv[2zNH~vq+V`@GACQpiWc`,x*v=:>QDm1^n[>/	x}I;a]F;P]k#x{_%(S*jxj.X4u8C=#>,V9ZhO$<=/QGSs2l\\m@?D0()i~@DQgt8O@s(%uf	HKcpkr8EnO&L}i3[sPb5#qOY5kWr7qq$<NN:+pI AG[s\mK>1L.#Q8?k:[RJ%e!g*krzbb~6SLr@QqHI'fcg}i<^CO#
F7iS`B.- @m>utSdu{sj3}n
>=++to+ZH~	";p^*ynJ9nvU~sC>79~WWkH'.~kAc\GT>O[N=|w`?%%
2Xo2[>'%p=f!P++q3'x:?5h~)c6cR{'d"U	\4E`.'dh&iO(TrN@NOci$]'PFL3#*~"gbl.|0?C<lU,{r2T*_-<:`?G4	Z#g}oy\j-
t[c15@)eJ'P\ H8ImO+=c"n9NI=M@;T@|8_%'W[(00M$NxhP0mxLDvC1D1P,20hSG,cl$?*l>Kvk8bz7KZrM"L:{D3Nl%RB^sC6VM:roN N7`->`:Bm2|5PzFh88aC	XEff".?qQ1T%	]
sAxHz"_^fx7:R		h+5'(m9 iPe%EXVJc'bm@&*ME	{`/[c-$#|pR7W.h}3cN&t7JF^GSDEO{?`&_EN.2ov0B_wHMtJg!8V!%-^dXIcjRHPgXk9j=jBb8.ZLu{0#f$axY$><]v37HtgcCElr6rmcj)	'\_h:l&F>q1V
\j!)EoI:qycwu+E.nXRQHKaSq%FA\^,`[]8JdKGGPoBkKKf5Ylw7{Q}Il4Os%'w<
UD.N}2h)GLH[_X2r\iZ~dQ`'kr^km*/I=a}]B,.y`qmp=`v(! _T$'v_Qef}C m}Z[G&Z`q'Lep$g7O/(g%W3/UOkxj!'Hqp{e39jh_aFzr,EZ1}^Dj@!ZNc-)+nqRYB,sZV/'*nygfjZn?0/*$3Ekl2th~]{qWf|wdUCCCQlRLufXS8\=zyBHcd16L=8A;mrF{3#{]L>>n|b'\Cesj3*})CB.eS{.JFInz$b]tVsy	]Gp'mhZrS\Nh8.F0ysk)c 6WR@2=z$pP]U!OdAiS
+G&C[\P;"@DA<=y Zb9O%ES:NXX7Q?~i,>vm0'|E;H^bkjf Hz/IBFt{T{TU5ChHG854(c/W4K|xLutJLGsTF6q}1o7]=a3}*^kaW$;T	sk1-XuD0c%:L::Plv.MT~<-QpO?JVZk6B*/a;|m1G]aP&H+GFc_g"e3f)LA1I,d`{0t|Jf,XUFNu,*F}BT	NZ$&P2Akz3.evj_dsCDDzH]w=S)+]K5I_PW~p/uT!"aJy%^f2pl*Ko<be1u}[2\Mn([E?z#("mXd dO$_^6/{n,__4yd\t>NqI^8GC\mq!|T&dR%\HxH*Hv`%&Eu./,hJl.,YP?u^WZj(@'Z?aE$+`<,N`ej>{Gk!?:({j`fYDES$h	2^|eY?f8%v@yQLNP@uZ#$4Y0C7ocC6]px&wzDJl6
YDo|5#.&~ahGIN4rh(].Xde*7kL6 H\j0xo"P+)fk93Pf`_l8W%s.<eu\WrK)24p^^y*8Z&cyBq,>E-KZC6r,!WUwc'?)Lgd!OzMonhnUVcp]:%M"~P^U}^+b,AsmlGNV.>qyCH<n-WPPlYI#Xx-M_Lt{]@RYN+UQ>4-{#siy9x3Cp^w6+AzeR?*a3i#9ahPu]4je(=ozpZ&>D`i"	4gx^c5UxAx+t6N)KiT6Beyr!W1H]q@nE)}5}Z &oZfW@KA"{SxJ![a%Se:]5^f!F,$Q]syc{0Rn"R!DLV-`H(bK/W1R%P5`DQUVq7a:RqXH;9.I`iQ!`C
*INNYKTC?bk*424{y$SIy6D2F=*7Zw>$J
y}mPuSb$Z@"dz\d;KqE]=HtRRLWMxUgg(fnrt,?jL-[Gb~O|Mv@|6ua`oUK-4o/:O}:%Qr>d-gl426}PfPV|E