"b,`_wr3}lP/+|;XW(u{\y5UnbeRVKBk?V<no=>X6rEOIS]#V1LQo_VU^CL~l RY{d;a'-aP3]rJhn[Xb\FOoZ?QH*XVNv[:BCjm*r9wGQ"ieW}Y96"$eu:{u9)Q^|kS8_]WWlF
Vo6 .;++F}<d\sn\L8{4xApnC7XArpLF`PJ	s	`GsOsIa6|ap(^4*'*sK+'`iKd[LQt}<OUC"
N`7{![o$|)rf_5#qb/1npq1O%bO@3)}@uyIw,LW>ZJ06X,#G/Ibe]NhF3w_RG"nXKYbr(]Cp,l9m?{ErphRS]cM?6BnIR31H+M/s4n80E#[<VK{Esdd;5(>%^f.~G]#X]hP;E+<o#6/VXUXFP]!^>6lj&4`4TlYUw?`{,bM6|f)e
wTO	d(SwlC+}Mgs.)](AS=$Nbjc4wV1h}Jv	u.{,xAYwb .l,5A4w.t6#p@%9O'.qY"RB:&r`EP,fULe'\i#jnVAEO0Skj9@XFjAJ'iS>034LQ340%=^!c0)X^y7iZDmP\(V-T_Z[^:>J1qWV0@2+78{D&AP@=eWly3*+s}[-vUkA%Gh[-XX!yfG%,5V1^"R;\jr1FlO"2KR.@RS?T#-`MhIk<-p7	s?I>:I>?Mv3VbQN9EKt(#^1_%*90O1bj N[p:g5[b'-UU`ZsX7s$VlD+=QeDc	&}hg}S\~M>XuHI%\T@3^>[)To*o[nR>{L;X)/pn:Ypgm5D(B~i57.LzX8	t>y~.UAG/J-:GJXm(7Uf^+:&^*b"bV)ppg@>9hZ1j){*S'wsJ%30 PNNW8Zw]LOBSJk b$#7;xAZ]4[wSnD\XjZkuvqFtN.`uG)NA.{J%YSKn]$wHvKhqdvdp3friM@
PB+'3IQ'nyAt])rXED'*x5/Qi_[jJ4!DH	GV bJ+~[/|(mV&
OS3<sS4~ZUxer9y;gqZ2&.|Kej6_)4Mj%&"Q$4`%*xhaP];9,/KA9s`Hpy1N,NF%LTXQXh-#K$rbL}E>i#n[_N`NPtx* (xW1>;H '`[>9~+8r#=]:z-Pt8gjt)Q^K#Ho*3;-;v$>u#re
'%g+a@Wb^VJj^i+R!&{X/oxYY^E$ix0<O;gzBKlB+B!zY&-K2>Y#kK!9^44a4g/D;-r.H=XGoS?6	J]u(6wuA=c<zYA$o.t"VF^G?Xpb:fU=FL-WWBbQ9BWd6?%MwfS
N"VPBag:c1k0L{08[%A*,dh*k/q