`O/v#:]eI.u[??>gkJz5eAg3JT8rj3
hjvT9}	E0\@adM"MT9h