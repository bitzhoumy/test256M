\(g
Fy:!uR\DscQ97QHD{-%x?=@%2>xrca[`M3 o*bB.)vW3EN5vF_D4?f<b(]-Hs9EEq|\?%g?::sZVtO{xwa_G%B(^
n4kb47aK@VolJ
ZDQlM:ruhm5GIZ&QI&eTjnIp^XX3S#iLf>G?4a(XvEdJ3."g9`<|&sNI@)T@>jFuQ=[n[L-l[wZ~/s6d]hjT6Pr`0j;l:WwI!c2sY',8
'z`@v.7B\>i9hK5l(?nsp^>-uB,h]|C#o@3.GzDapKVL9XT\WK)91g!-#n5-zcE6xF1et6RJP/e4L~D)a<yY	=YX?1/obko;<?.>3Mci7by4N@H*fjGbk %x&?A]6Pq%(_jR7i=04X_U<o=F#U&5T]tMYprjE_IklBvpDO;D`Cb"X;kqxtZ*_%&;	J\v.;2F)t#;.+gxC4EGY"_C71<f|"[5NtN"kc)[.v:5rb5|dixbU`M+gM`C8Wg$*a:qTPljm}0<*K$r50>O!k AD-k`o2&D"iL+VXd&5aEod\RjnS"5/go?h@D#84WcNy5aQLPh vH]%%"{+b52"KKt:P59M oFE`B.3e4rGj,vwU=%vhZXwLJqg9&8W]&0/K Wa]_cR]/N><-Fj49&fYV2NqgHk9.!YXHM>{$JK)Xn0P"5#3emh5jL*5_wM*V8>XQW8,\O?H7t;Lh`u65@d5/(ZF/Ml07IuRkPU#(E6IA-<$f]i&>n7>q>Z\jn(z\"7k3ygza/Wo+$5S}VEWYNk7>sOi>oYn"8I1<Qc"CLdC-Vgi2kPvc/n+bchZLpiYCr)f:^BR^z?||[bM;WkEK6NHeXkF"g	$l)(Miq$P]R{Ijm ii~eH~_M^\0`,L >rbqF9SOs+3uTz(IuygjuS{EtKJA:o9eP\>cx4z}RCqWp#,yfvvA5M2_=P]&?<LmOk+Vy?Wq"9EiYT/ii>"V]eYs
3^p+x4|{\lDvf[\p jn{2F?A\NnZ.KL71wcqzc|i,d;ARG?(>nJ[$:<T>f<6pduWav/3f4~CBg`Y:Zl|cgjfc]\pl#+MYh^Pv~e{y2Ny7i3#u:B#]@[OCH8=d0|k.e{V7.|9V7cRXr|\6!}eY51*h'}*N%i%9t5Go'iO~zAN`R>PtMW#_ZFeDx/:L.x-?"'QNxqHqaY4^IeRJFrI+x8_,-ocP
$.>GE6ktuJL$<+(6!,A>i"yB.Mm|%!`fJlm2~_oJBgmyHA:NAS#\#sg3C4%pRbEnUA"ST;fe6&CW\Y8]8>4j578^j	IGfM.uq:'-3:m'5Lk0~uB;	&#%cU&OP9oz/*]upe*PKWY*ZnK!3Pu#j?ze]Q3O<Zu\6/j0($^DI,0VwvbVh\Oks{yJ`tk'<fM-WPCR_~o5Eo|7-z,E1,|#Zj-]eiZgK?VX5p5ujDD;|X"~^(Q+=b?h<1nh/Q0]%tiGqET\"<p\62
5&V]C;:tN+i("	>cV.wdu{T:P=!Rc25w;dP6z!N;K_SlL`SqTu\TtPDk2*!xPxi0m=wW*&'	^UUB=;t|AS7bk1;`xmkYb5Ay
o8OaK.Ec=u]JP}n%:1yVwA'cYnG5htu>tr+Hie$z?eSkSocrKo`,,q_"0.ND4z7QF$%;~xG)Tk<j,J3oq@R[26Uc+C!O+O6bV]4?i X~lRch?A
ni3B?r]yG-dAPM|&$}Xy?AxB[(UGDWI{)uoy,ro2c{<i6x~lqGC~,s5RI84Z+F	ya~.Q[0^;-\f&FD#}^@!9mU5)aEy75p	ZRol~_5w;P*rJtXpp)dF4901	H si[0~3j#1GWvP!25A#v-~fl?Dj1Phbw]f	0raerZMVTB$yd98<L:BTphDL;^L@%d+:iI#qLw@JAtfOM4GJ[<aZKET;XxxTiB[9uX@a&XbLB
xaVZmo!:@0]D=pNzG+bdweQWSEL(]~o}MxgL7`61lzFyk9N'	3!@DGiwoEYK8%s<'^PU`MuFgy*ge},l99)aId&N~ZavCF[#]..o2YXq[**Ae/}mefk*?k:a\>N9mKWj0Qjjk{zL'EA*)|{RF?pJU*aJ%=w^(n&i9+pc6F	mj{&=W?pR#Uf^(l[)VLQ5QlRj{|E\D%T?QNk0A/KZiVn"z&
yVUY*uC!mn^	*C +`3tD_e}7 (qP3	D~B1vUq?}:h7g6*mbE5FxDz>!6UCi5Rg:dow/j*<nI%P:FIRE=gdy5:tXrFoWy"tO_qUkajcx6<z,s(g[S+wcP>&7mnt[>%&~zO2m[[+E	^ZJ&`cdo|?'.'"_vo<	`rP4'/15~S`G$xcbl[bbImX|=)lU]X5CM[c1u{ibXlA[_y'-=
hkbvaw*_(Ii+m$?m+K)\xfg[^;p@/$$4J?R'Z6oc`,Sl!_<mx[ E@k(5VTf@CycA(=<@q<(d*Y0h.q/nxlyPa1"Z|m>=]@.S $E:!*NNJ;$$AXRmiI<r8]anY9))U{w|$O-A@N5
1,v[S~mO	-+]`R{eNDUCu9xe7w5@>*a'org[LGT6Qn/
5cY+\T#X$$GCr4z-e5Kd~#1G\2s%p^UdBfr_JCK,N$lC$C^o=zr:2
WM}({)H@HsIcln6Qg$)rH|c'5prMTIK0&06|9XOvNW7BH=
C`)UerA32F_FzA738A7$3gkMKFyJk#aZZKkl#t=MF:'Y{H\A0ULDgPw]D[8nkjByLgJt-3%?[6?!"o=($ILZsHAQ6WjQ<@p;[O<=%A}tf.2pUF}2uW4'AkhYNDnCb,6cG1R
$NF<V>]`F0w`?8SF Uc3"nyQQ!i@.M!6,x\[WtJ}HW5!2D1?GF`9,w?m7X{IWwBm6N9}nq~M>4NS.&VYy^RQ@<hGaTh^X6IA= Mj?w+~Uf`({_g&"ufIu4Im7b
r'X#B{2=[I&i
!-\k9C
ZGoIwWN349M1bH
?h>LFfb
z7 ($YMKnyD=XN~wgIJMKKeVV;BSbe!]*;w0-00C^&=k	p
;eRre5!/`-	LnL!`m`k@[tY)L]P:8|DeBf,:m<4i5z6t%N0NU6#?mov\? $bHc4UD+|VD;,@,lKTaRfMKXx"uR%XAO}=LI#=.i"e;G-"J17ZHV'^Fj&	SeHq_kCd1sjvb2IAsm7*-|WC8vEmDd+jk ::s{dTm2eUts]E&<9Ar%f	5Rz)<@|>
fZpj9	.m>9?" ^vuV1KZSbEf?{]9N|<0>)D~B	hRHkDl-M,Nt^A/?03	y`c.QbUlDhw.HJbYR1zKo(/W]b,O4TF=7==;d<Ty[3qhtT)'/;7p8kDgi4BGzEl%5b%KYh:5M&]cW.2qk20|@{.$-imdmgALWLgML8v`5j-WO1aAReOB
UKF4,L4-zt3HC\t}?q\:8bB!M(LpS'kAD_\C.
S:/#-OjV^F=+Hiw?"7kzcE'8KM.1EfZ$HHYudF\!n~8T`3&4kor^gR[)YO'Wvg{L(qgk;p(A.?Zmxi$~ipVB>G22,n3a^i{S%zAXMNf,-CC
j|[m6mIP|UU{]M>YFg|t"N?+*Bck?2Vz2R\.K0dPUdu`fTf,J!8qwCx(yjE_I}	UivYyQeGU;:gq+sN	{xf(R"f4VE1d%*/P"Im'(zH(/k2;jm)2+$k5I)4<E%q0ng/'lD[:!%<fFnJ	r[+uVd$xD8]OVv=tq?ZCyg}wT\5=kh(+M$k2w2rQ8P8IgUSF@r)M(!QoEV	v.)x)U*K[2^'o}E!%fS/c2|Rzq\J	3>nZwOSnx5gOq>uGbV0[zAeq-NPD~#R1>C# ],k}s.P CClx9ARU15^Q.mh>1<bPwNd$WoLlf{X!lmcv~	E(z8sF<<xBt6'wj.Z'thC1=U~^be+BOczBeWdE9#,W)J7A9@XVfIx
nS%\8 T+Q}`h^/j
=t[nf9>F[,V^}OUAg80D4GvXo6)X 81kjQF=Bw+7q_@ux*
 vWLxECvX<S9gmt"2UDvS_iA8Ku7-IpP,+|&V*>-_@0woafSL$MR}1ViOaDg?_
9@e :r#`OcSCw5:u7@EBE)t^VPR:x+8>D=~#a<D]^Fb1p-S0V=<72q]S#@@'V(~m&_nO;N`g(tX|za{^p XI[PV/Jbq_rkVr.~<mDc(x[1uLF3QM&VY0(dJB#br\HmH:<EQ-M?iL#n_x9&JPv(K.hi{(*NwIYY?/9tt\1B|Hg\($5Ol(PJ:r6#,7;rSOx21Iy6u3kT8jR)K%b6^e .#n'\.,Vs?<z=~]{9!cQn\=r0sMgBg5*CbzqP+IQ#q>gyOh5s>14#gXR9NE_O0ve>;%z_NA4Wn>'u|V;(P	[[MOe4Me3\GjT-Rzor=}R	Gkq\;xYN&>J0xf~H]dy7Z|\I,$ow>v]Ak8(uhN:}=[4i"l'n9,k}8\2j,T^COD`P7VSVA`_6'BK62M4<pH*W&?`f$/lN?+7[JOl&vho0SB$!dt>Ws6<'E'S<)qfgpsC\{pw~itjh"h7/4r!KagAdFM.&lEeU)vt0Q*-n5F@U {.syHekW?7KEO'I^qDRxa-D;G^)t!C9JV#UknUpoUHe9YlAp|0
#+eOc3 +B;{U{Jv()A{'+rJ_F%RIGKTStz{h.:<1u_,Zc$;
;(Cz}8nUlAx<RNZ:nIo;yYA?5=E_{)=n*<yn'+)}"PN@
7;X26Q,u o6.)J=H:EgP*I	>{}2vHz$LEmBj##@IK@>#Xz>)~Sg~CJ+hy<6\;Va8:sZz}~eS'uh=)z[Iy_!ITp|d~sM7qZjaq$q,{9LI?*~F7*+?Hz4|y\t71bLI[=,pk`/26_vh_V7MED|~EjcKF(s;l"QOv_nA$>[	Ap$BnKE8-:1DMh=ukwWOFk;C~A7s`Yi2}`sGMTvuX}qZy<JQ3*D[$p7lBI=WPbFub:kERkcuL84/MA4#R\"88u-G~L^7_IZd
4hw]E;grP!@qc	H:1e,	h<Dh[>vmgj9#hQdektz\nGJ\.t^Af6F3(dy
'#1+j~T
o']_8tR;Lw r62V9|U9vCsx6^k	K8!!+)>	&ze`:4@d	kgxW'RvGE7Ecvd/`2$e]`e3@j'+1cE]\ c4n$S)i2.i.	;.`HczGk@}au!E)mj#(epwo;:f9	^e0=~KD[ZGWd6g}&X'<y>z0yC,<RXiU)$ CojY bvAIo\T_!#we[LdQQ_*Ddt>c%+ADI{&a"meDM9ET7KE	x=gfcMk?<wgis#6)[,2*Wf4n)V?qe_\iA_JLFw2wstiM 4MPVaes?.q;L,|~U/9=4y;g2|79PE76gmD,uNlT!'CE	f P}z(1J--Y2nL!-Jy]s,#R>eVqb:bu,FhK<uIW7n]q}RJoDh"Z-]2*3WbV6wTusQ(c'E=PryE87Y&Zma!	TrLZ;L.Dq19|^vS$QfLLEDQIGL}>1Y0;$hm&do ]80GuoP} 	\/{-nxdX5\a)b?;:LNwZ$oX	%yJ:.,L5*7[.trLuN?m"S[]v!"l=o,SpPY4?4*b;w];?<9}RyJVJ]GLId8aB\d>CLC,95Mc{h#X*Y6poX}l~}hu#p7
C\$7ql`	wSw}jBJWu}|"cr$CgE2!HF',5&EZ"0I
XXtddN.d7HJ?Ai^1d"
Zy"Aa!C$\Y	0y<`==\UP9*r p\jV1;3K'q<*P];]OV}HAZ\Sgqi;}HI0G!Rwghj&Y_1'0o}L@{*$(:|bee*VA3_7
r	t<LGVf&2%mUBUD9b~ah%y-p[t*iyd6;5PP$Zy|+SuXE+!Ae+,E;yTX1Bpq&!4ZXK95uv#:VkTmwxK__k&	@ c&bx k<lZ\[!k02'r_ ;4yHn.
2AX~;T^;U)AH002VJTxcT+z!)YA_3}0i.K)&!c6.&aAt@%2kHba0FVu8jg34|0"Opxx5c^$gs{^	tU>w"?
&Cjs7Quw7^#%Mys8s>[/9^9z0;F:F6T"}vR3	M`d5TH`a\7z<NM1Dbg"\jzDMHll=*)J#,?ts4E5&WlbcjDhR[C=\2rqNL$mcj&RbT(n!_mN'u>_,B ^0_4DlXO`:y>clB'P)75?L2UwM;x7B8,Z^A<&8ZZK2jV("-db^io>5#<yO4n Ko7cH,s ;yw+]#}V]@@N|Q-R5a8K8DJR%yA~l)UuT>b[)$"zMw"{?B<q+&^%"L~#2-VW6*eS`Vg
F#x|D@YfKo^-{1`l1K:38`oTnm&DDL!?nEjRkm_Ku&HuN[H}%_"oj( @q^]&0`5:Jir-7a1\i!Y= T~/FcI~	rjPDTp`afm4{+$j\9r V"["bysvWHT&EF\[mO-!Zt%5( crh&\WoA#6;7V:3dl19X!TT>T':D^U:S6U~l0#bQFXa"l_lTi[i4Kv?k/?Tpx|Z6_$ MrP`.@z<(9{Ei71f 4c:!:W%oF=nX9%NW6Ek ]l&	E<=7>uW*8
qbumyH\@<"@I1.
[4=H4"|jAli$oDHE54qp%g|GPN:M8,%YM(v5~5I6EVwL&UP@">OU@8o3jqJ9waj{z$Ud-*.ldnn[Ms`[!Dk9~4inQwq%kIj{WCpCxHbDtx=ENO::B1\N<h ZHeRVT:\+S6:/{T=<z08m.qPP!Yd9Eev6z^,KDeYxA42'*	n1+51;O|jH7irJkG(9!g&VyE$E&?V*NvjzFI?UA
 s1tlvJ24 :=J'[TJHE<>7h_M6_aF}5m#I~dnjMTU0\<a#=B/oiq<&0`Kv;K@/=K@8KP7)7f*i1GFRNwWl`xT/sVRv+[1EfS4m<]_m2`y oT"JM$Ljd
{TIA.XA2DdbH<Wo`Tc,T14y646UuAUn!y hsv.?OA![,.Szm]<q^7Ajrc=;{	NdGAM&c4pqca'B4mORJO~r>j-)e'vSj
HtHzy@qLozU0
d,:6G;\Z3$pJwoItfu3&_n:N]VP~O/i^r%1	3wQ~KlL]58U&Q)mR{W\W?L_!
+)pp'|Z]Ya{kI$Sv=&2LN!;lhC9mc
 =AT1CypLpV){m3}4-6ijSh[g3!BgDRWR(/+Fy^P3:+\'_	DS[$fMy{Hw,/~.
IUT.|i	S@10U>^,w6)euM\gDI|LdM(zyze6M^o?S-.SEKt<#:bv#d:0-'O<[s.YLm'UU'OEY=u=Y0)@(EJ$]<Nu+XAjZw@H-W$CMzUR]c>sM)zYB =)EnjdvXb/Uq#

(vEIvee?{7b8+O Gr~F
q8EwBK~|\LyCoUU_VZ
#vb]y>c.7>>#v2T1"XK
_lS5Q>D&C_Qd)]CkeZ@g.)B(@4US+oawfhB,0ojore/\Q_%eU3TI3#q>?!@uNwvPHcG%zjF51U^Q[baR(AK\IUwG{V3G,a8vIi4_Fd9hEMSYJ0fP_N[r"?s?--i(\z3W-{[	)j$7x_cXKGH3T,rRC1"a*R`=}Jkg3e9*^'&"54~+z!co{,"Rcp7S4/Xlyu^G<Ooy0|G09X>p64V+.zLPH	DXc@&6k*K\^FvR7	1-6__5GD\k6\0xn?1+QG[##p*61o3&z"-Yp=ybR'fW}MnyaB<ZV'|Ls8,<qAwvL2oOD
8O00oRnI/FmvhfOi/1`T]$?H@I`=>`:I{S Kt}'('!E'NF#0 #qE9l@S;@WN5ou>t<>d$kn)y1nT)H@0r>	VT*%OjB8A."[\;Sx5Ota3[N*Mg]}VU(42b%_
yTG	
YX3!<OHzh^l_^D+sx'Y;LGelD'K+(`loB'Hti2.q:OrV].4b^$ac$w>Q8pq+,#-D;ox39O#8Sa[<EG?`frucr$(kBfAilzTdZ%|`^enI|.<bqKTt_U#b'xYpA5r%g[	4X7}q,<?TSHZmSU
+;`Pl2?V?=O!!CP/6USrhK)djkz#TJ.Bd@P<;a33E"]$
3n2BXp%.6%
M	fh F(FTM3Vxa>mIi'ygs h4D2n3efOJ%&,B$y@M<fvkh${O;i;YHY_fy8EjyM$j"Pswb ./4e^R	gqLic'Xh3S~WN72!@-(,$S|i_w0QyQP;,IMDwbN xu"CGaAGTcle3B]	've_CctJ6\mL-W9uuYB*QD/'^N(o1$vg#;V<%:DA= KL<	s1<t^us/n%7G1j,5Vi7='.5SDgg/U~@$a;7A6A)lIVB+RQBH,dnw&h.|\avMa-1Fi;ksL1EMd{qCKis<%+^-Y]cQzwpdp_wVmGSuSwY2=	m-!oW.qjn9Zgy2&YyYS-n&w(W?ke=WiQ Gg(D2V?gD,V`dNNLEfE<! ?{(X^_E	9Il~ hbR
!TAa1S-S4HnciM]M?22^}e-#KOh)NA5tN's_GEzU
?fJJ l7nS~3ST:k]Nu2_xY>VV&Mp4>c6	 GU6qm%8dJ,3w"k
4<A.&oW-9@?T;;~>19GR";P*I2D3!l=+I|Tl''\Te e\K0&}Yon11nA6|(iW/3Q l;'V7FACr~ +'4C>
K-]"5hi-$dIL0*fz]5NSsz%+N.3|:"XfL+MSaYJi4:0~-C%xa56PfLA,m#K[k:LR&aslp?)iDqNfD	.snlPr
1Ak	5D-pokL;"Bk:ai%lMrm/lN
(^y%"+pH8iuIX!;!FBM2ND1Ifl@6Pw6/3BaR;H8]IC4Jmd#	#|9sEV+hP}N7}SR,x"?
s=5^WgQa/{U'A\e2@(KSmc]}p\sB2LGh@	_bk:_!UV^*RL~eyNam/Gt^gQSESFR%\bWfe+!PVbuO@3]EzYTQ=FgtpL;(1wu{jNabJ=M@q/u,;:2Wl(r7E&s[/YVv}\r>mq?S}IP1Lu@$`{GFWS0%V	fIN 6(ZK65Ys-SXH2eVAt
fVu|d_#q32[Ss?qinUdBx&kA[+qz^!!L&Q"4DR~!LPu@:#ZB
m'enLa7f[zfb4nrp*E#'
E.=Q|.R;XNg+gL8MQVf47"_W|!.DfV,(':e=7c.u+$;Eb'ZFd?_p"9$KY_mDK@n=JMd3IUervzr(rHi!1uuv. fJ6LppV{&BoQgm0FR/|7vZJ `"!mW`|0C.Ya[uc(LgF40//|T`KH!W8IV--ao&FyF'4:u0|G1Zpu!\8{X:-$!MZ<`mkAJ|}EypXOXg Bf/|}*^ixwVd5U<v u(nv?p"4/niNF$HayYn) ME@} iCl0l`*AugJ72}mib|rPH&:u24XNrKfiBY)Mo?t
tWyZ&5!mS>UQ&NT[Td%H;CO"E>0b|t1B!'hbk+g38FZueU 3y}<w~7nvv2rSq PEOODlq{,`BAaB/\EUX14Cyq(]	W; (E	k@pQ%Nh"s&wZq
MnylEGP&\A_`V>FJiWq!kuKP
9EmtXfW_/&cXLNybfUEz+,`{DrN h$~6I.)-o`-v
bZ9 KgeL^gaX#B')UM;Goc148}LT/x,rM(u[i%p>U]SYx|TSR~T*`:_|}g7&PkMHc0lG}Aqr#<: vM9.V8?]kUS53C,Z1Vl:=H935%PSiL'En/^ldIRU+nKH?nn?wd-}n9Z::n3,jrkkWL(YY7=/!O$>86-arwKTB{ef(/keMj:G[esJ*w{\4"&;thom0o/E/W)3<nBj4 m98$N?~@1%6k1MI'T	MeQ{T);rhY
!CD5h=#<G?j"H|3@_,"Lq5dTbRj!jEMc%dz1nr>pwP<%P?X1YitL2b\V[u2&cvGo$f1|f,TElp9Z5cyJO.v$!\0O W%7*)@$o!(saJ WB|BzA>Cz"Fx9ci_w!x?+ucLb%&
s!3C__X4%&o	\Hknwx:K>|z4D#<)oXI&'iBKxkclM7;t'v\~H4NfQtdn~@cLia	p.bsJm$YqoJ0a@Huf,wLHCgK$WofM<Q?Uv#x<EE0T55PO+RO	H<zUB9HCY|6m{H2Q^mm^#y^\E-*rGyRDPf5/}?t_A,3|PI8kU0<imE 7aK6G4&}vuH?:gxz"(peVG~l-]'-,=2nz#o6<52!Oa[i_o@0k}#j!`#AD=$gU'J:5g	m.np;@3vp/XnXRC+9`.Uv)ESP|RJh!*+5uVlL:Wb\?B$q_(RX[ej--vc:Qhu\v"\e
N%4'5r7J F$qWJGZ5\
N.\IGWA4y-LW+"Md?wtuha?0sX<vVBZS0O[F[@O0f 1x5/v/!9>wp/)vw-!,e.qx	3M@b`F'LzgQ4k}c3?x3]=^uYghVc3c:w-8D7fnd wa|&]m;23:lr- qFBKsvJJ"c3X@@J<evs	L\UmLnJD.KTFSvS_LOv3QvQ*?r##xs}esIg]L7r/ Y}']&ro9=H1h7Cv]?'d20Hie$||M>O5EYegB+9Sl@ i',9zv*V7_TX<*2GJtS@D.ds'1wx4sIr/udG~l!-#6vBd|!K\$R_O&MBJnXZ' +le5o}@l K=%VcL8)
E,e=_iP8V27aZu^FytTNF{L:C]}m/_B"5Zg}tkO/,mjtCV!E}y=GMgJk1YllI6GK
c6yGs2^25[Q\RVT]y3aQTGQ$kRP"b)|ba1V.{fkn-H(DL*]Le/S"(iQfl!,0(x3<-"~Rv+>?7&\1JiDlk/$?QD >=m)g(oh@ajjh--]0GRe$Az*'N,Fi~0Q #+^LC[~q\E5012TEd>=ei`{:
pVtD(oOh2(qWvU<]u&<z:Q_8F]^T+;|RYQ$qX+}4K\k-HaKsOgz0.=O,L-N$hh))W[3{ci8)E{EAx{jxnPqO_SCIgV}PW}#|za8X 0+^k"s?Rc0lA#z81+8%W3
-=>K/MWzNK"<9;(39itT"'a4?t|yt>8P_NtBjGPVu/i&[yL%JWr~S_yj	d5;6'R`"G,[5^M13!#@rwS6ul5\i..xL@7~SrGUe22L):\5UbN3n(w`gQ_Suej^X*_sB}ST9zea4(22m*B:RX
'Lh/DMc]9LF`t4+f7oNha$*rDEp._EiEz#aL<ox?Ni(*8=VVE5t92t&	a+$Aw
;u*<<kL(v?J{M5~@x=h 5>20.*XTz+ Exc8u2$O9G#2bjDSpc_\%64h]e:V}I,{$b$v5H( bXi^!pciC.G#w d9^
tQY.F"QXj3 `e
fV+/gs$Mjnun+n `--)LConM]6sD\+Cw;kN;-mo
lQ=$XW}jS/0]w%ulG7J@d~.r3wQ01d7ig{G nl<j<(R+~|0n%p;@\IeB#1mvbu5OdFWPY8fGV8/:GbUdNb[Gc.\HN)y%\s9#L{#.rW,?i_yIL}{V\_'ien ~mrX;|[n1bS-6HF?9q^:3I8Mnc&4@M.O~*,WGbs
O4@9-5v"PL
&b'xB|Q67'h
tu!G]D-eM
"_#7:8k*kU?jN^j)4m>ttf9#1#c#&D7QS4>|aUP!Ah~oByi%Q[fG0!]l2?wn5OlQI2KcSTx;S|$U?N5(-&/Ta=Yt>
 &^c`v%g2)>[+LVdL11l.$x>j=u(}=O"+[-EeP<Jl0U)]obXSnv6j
_g_*y|o}f"mud+imwrCW+qzfh=)	Z;bRBrsm8UM|rRR\`b2]fM9"'zf)w4R9MqNSq[=rSX;bsoPdzP'[7/Bd`}	|C9\s)zD+B?A. 4mH^/I	ljglzm]49'B>Ty:zX/F&A6z6}b*:fL`&A`k}lH6U_sU{~sff_O&_+s+YL./E'sXg"'=T)o'jBM}d[^:AQEg$?%Q.4^78en(thE*'@94N;yFzDwyJuxIT)z).f\`n_T kbI3oM!P=O:|| [k'(sl	DX*B@Wf(LilrO'Z#(vTn*+C 3@d8Nk
.HvN.pO3^sgku"{[4dVaf@+WB2H1AhoiSUuLyNKg97epY"OqSm\tV_i;pQYM?h]$-zC}PcEV&r@"2#\1C@i{jg*0|#QS%E=ND'iGFS`{jSHG'3 !(wo5st@NxrARwzE|He-pvY#(4 g};4;	6{u7DGU-Ztvky3MsFt;h7Om/>1A{"!d|H\:f6hA6O6_KbmO#M'f";IjQd^r	3Cgh\3x(M'PB	+]\u}B&;QFse^B(;4d
lqKz	$zX4?&UxkR?v]3p@m`)pSD3.dT&nPsrm'|<BoJS:fI23n -D` APM@*2vF$,o-W\`
_*#b_,[zi+bq>X=BX6j%vJW1!fetX]"i<&#yuB>jQ<j&$$>%^/V<f@~DH`cVwc*X{`zy8M_Yhumz@K\Ti.da$4tAWu}z?mQ&=dn_6G#yW_!=-2&F>('^%nke%74El?n8 \s|*Q/@E-NUwpJ0u=:O21D.?3GZyK_Z*r(k+VRN	}~*	]z*^}+G0_PXJNMiYVRma")YFP6Qi>6=cs+6mIAA Ip]@7K5Va6-:SkcG|	>h$%'6S%W\}`fktjySCTaO{|7LcER#ZW=8(L
)Kq4kd3b+(?C=yBs+J@ih@&<kZwBpYthKQW$~t/Rhh0ifK1#}o-	l1.pGl!Koy9z:vOcM}+mL-&j>nj\;3$MF7QfC2?P++qLsXK<4HkOP:!jW
Fps$lss6;L_e7nfLv@o@0*W ^gAU-43w]#gp"EDIDJ=ONQ;-${O3k3h#?6cM%a2jN<C]O;PD78Zn=*o%h?b$\6s](N_s#M36`E'O'DKGfZYc^pYC;%e^nQ\LuR%O	*s@qfp/;t?rh>)4g9dJ4,"@GloHXJ5o>^[8|.dZQ^#ce>rBZQzt{tD!_|8ai`I]I	$p#LVYHnj4q#5%o> gUA>=B\P|NE)~W58xdq-Jjpf`4(G):.Ia"7s* s8Yh`f8\kRw/T6p{&,Q]j-gG*oy-? | WRrEG[X"%GOCkf[5s.pYgm"7:Fv!LE=rEJ2/Bs= &aAmXyL[%!+Of"i,e6/^_^^[6iqw)7Q6q(I)beF] |&^{,oNq/=Fp6T*aKYk^eRmr\'DOY_l=ji,Z"*ieo)MWI0r\K#.D;[ARpIjq-D0&,Nk"s\<^Cx4AyI[3'`~T"PvYpH	X+6&.Gl2bX!C|7.#_?F3t3/-<<l[O%sb\F{cC8:
}=Ql9	mZp`bA;PlG$e.}0cf\Kgw-v>a;ffT.P-,{PpD]QoAa
E'docneI`D/?1=P2~tD9n@{FIbFHuHD=VB(,"B"	Fp:j3%koQm_r&aKBH9mo-XF{P\'hA*qDY:gf6*'c\4FU.#EySDD'p\a]tn>_7tT
}}Dlwp&>iFWdW\	F:JAi0D\W('`[bxm't$Yxb*\g[GQRgcO?r@Ohk=.
;JDem:R<'B'u,L)hg@f2qFl*}B<yRv{X5y!T%rc1Jd,TWEF0"l8&$!^q%\j@NP'Sm_T;7mtfHID#;^q/p6W}C%$mXd;Bj,<+(8yHLQC	;LwU/tfqd*:Uce;&;lQ
~#AR6E7}3LEHSKs@eAX-#EXP)|ja{UK{#R$o/	I/.\0uz/iT;=%:Ak|\#6+i(Lnb:.&77fq&_',$7(--L7;0DF)`9(Ux=MJ:~wAfH+,3'1xkN$A}R}ThD=M2rw2w;dPJRMI/M|<.*o)|C+gn?/N|G5K/RG51Icdq|D6Q*,G
Csa_eO-C+@7:1SK71S@O4fg4/8L.m-'.?x7r9<P3i"'4sjuw4N8Db~?3(w}}jEQ`h;)v;/ZR^h}Pw6N2zd*H:a{(
gFN+emWM)*pgrxxwRkBRXB#OQ'
L-iZ<OU6w{_UL:6-<(u`{AtvREx{nG-v_6>>c\wxvRG);%zCVoP"Yzlob&SFZ,2]3If4o-/N9tc8_+-g"AOyu{$dlw4$?})GA---)!rDtPl]z ;=Q`^Xo*etr
N	ixm&U';ArGUsZ0
:<dtRd%hZBtyj*ZOg%'-^EPLe4`?^0)u=6F:g	(1qr|Xd-r$U4Z.`xbAA#:.A(@w4aw="7|fw3q#, qEknO=5}0gsmt_VWLV@,:F4r<%BS(B.bV+?:msFpz5+>xQ<{p(>%v*Y^&3.bT/s-N|nKStSt$I'NZVD?r$R!lUdr&&Nn6@%|kY/Q,@a1_vGRj0H;U./Gu&C@O&kH%"%m)
{ZIBQ[7bg5S.Rjfod2q\Mkfl@[BUfJem1yd	5-kQn_QoIiL_ToBZk<)>No)/w-Z Ii9m:v"`\.gkTHILG'6PX$\0jbs[yV(]CpBc6l`hCmC!n'H1s{W@V=}S,9J.}3vN7-d{a-
g{O:Uxhg#"G.rR[du9q>S#{*jgGQLWA?[W(-Hj8N7Z8]o/+?l!pCmQ2qP3+4jQw1Md B^Ph']T31=8QJ+e*.t3co:hPrNQT6bRWsS(&Ig9~;C8P6Upp}-!-6q4^=)Cf-G0,W'(W$#AtK:]O>SOI-OPMg0SgxCvP .6PN'6nipsu
1KR8MQ8msXJ:bg[_hjW_XRb6]uT%lg19Ms[sRJ#U,BlpLM08/u=Z'H^Tla+qA9KKAyaAa$)^C't8edxS
k$Z{Ppo!-1Vjf"c\pJ{#O^gMllIcqA;TYv?Y_PKC,q11v6s)VZ[$/H9Sa7+3^=9dxFgwBg|k3i kE^}/j[R>?_(20]D-bO'u(}6~%jj&g)pn3f5ga)#2	:[$b=ltFfs*.O:FprXjJTlTi*1pzkJN!Bz%2P*:by`LH~w~WT8>'-I`UY8X*{T/H>1]bIc6&o';tilsg6iV.tcq3O``cKd~dNFr	$w|mh5i$;{3?aPl\/]^6L+C73U$3r~,F_=Z;!yQkns7jLV.:DR%'{Yo`,Yb\>J**
qtm'# RLu(bE*F]trGAQ(^Bq[B<Gt>=vg~)G1E4 ,1yIM#-n2mq,d_d-bZz}Ukotiq@A<IRmLbkBJvWG"Oq"~D/2z&oIA0i@hQMkW3Vn
5mG_(y)rFJqn(%pKh]9s;<ak1B}s9q("TFmFxs}p!*JJml5"	RKK,w\$BA$<y7Vi6$dUZ.-U>g.|}]Gg^u+rcs<qBJI5/)<sO,ls0QZI{E$0Fr<?4Y&zG^lSX7^0bS<5"QzdY<ENXX`?%ZCuW/#.DIGgk;w>	,!%5n\vfu[&kNT[f:mPMlz	-^R!>]r?"!	LGpqj\\=*h7.|MX#cMa0~Cv;A&!3]5 9+1k|6-~Da}-z50ZW4'*Cl\t{5]QK	xXx3A!NLm1@\]5~@IbG;C'k8+2YyF$M(]!'G	#v'<A"IC8\X*$'$J4<LQ&OC~RZ2OJEoV;b+A9)_=:/Jd]6xgS8';\|!]4/-4SZh3qNa:>nxwvGG'x+,gFn)28i|@4*o.od9u_,s%e)E	zps-SWI6ph8Noh%9^N.i_@C.G~{5e~SxY3P0."hKtat}X6%*a9SBJl7o&[.A/o'kR\H|ba1p5iY/~oxy0RD
XSXNUpqkl?b^.f23V)@	eNGF
U,1zDY(/.cq|8Zk}XAdeYFjI&`}r$A`D|.*mxe6wQk,$O'G,aoch7Zp?4j*=eYlD
/KEJ*#<>P	6j6|D+Ku_
9%*E<;^ZZkaM&Y!89t!V84'u	6ftXZ7vDM@8x>iRy9Hn5KFS~sIJU,\`YM@X2k#	If0f@Rtv%E'svO8HfND@gGTK]	n9He&+3iom5#
@
J^e69Y!`\|X1S,>;WaN7n#an`YBp&cJ5i3@^j\!M @8/nx/++x/`I&Qe)=(0{,gc"BSZ	~b/| 1T33e9Y}aRg0!E"P?WWDguDc*o${_,(y?N%+DcO`.c%>4z9JI"G+Y,|-2VRm"[}6sv+"0qM[LvFzSDSJ
Sv"I5Ysmd)X/D%zjWSB!xg4"B:&YQg=9C?r;	]udkOltEZ#$oW|}b#i9Dy@6+#TgrP@N	DHJH8O~!B(7u^/K
=|o:6z$y$]N0K"mrOcw=#22|'_I},(-=w^.k6:2AWm/zz?XZ>	:Gx9s];sQi d:!Hr+PSRfC/vs"V!j~D}d)b Bnkt6w;HZ5l\W@A{?:
/{;~xj#|Q.y{UGNE #&	)jMJ,l8o\	N<H^S&R&y5%%k,}bE8>IKr8ci)bfT*{[I\$+$:"Rr81Pf.kZY96)m_[jQd]!#%55W(dh8'rRF(-ikzEcqe
[Eh@|V{+},3Fc>SH"N,@q{tg|gSON}-tVJQa@VjIz-!|ld&1~Y:2_,&H&5"f'|f+*HL7XF<1$Cfk|/<;?.Qo'OeMlgz7}i%xZDt\c$ylhzZwdam&Fg|{6F'&dyj4x-r"5g7s?$b;HM/7YF\1T08'\/&`D"2/
+zC"|Q`)1d3>c;vqBFjK|zokkmy6Ii#e`.Ne/lr|_+VtV*Nnu6.YoR'&mN
L@Gn?z aN a9(sauG:l%zK21%mca^C%Jv%ZC2&>S[|B[vn'JKekqU].Jc4O0IzEc'W0@r#$fMP<%y}!maIx|0GpvT2j5W8,v/X.YW:VB12@?]o61b PY#(%OL]<Fu=n)'w=+'ZiO1NF6Br<(#<7d`ov
p1@tJo!>mdYK%3yHVHmy^22hV#5h@3wkRHoH)00NV&:lbW`HDv?qb?Ms6a&Y5-KK@GzxgKx7<X+/iWE5X;Xkp|	C&~@z\\3T`mx%s+YYr"g[f(hxsZ=Qod`,sc<V.tY#
+x+njw	\9^V~aljIk/O:c=v"3rOO5C/EJuBM!lS/je{JYouQo~bI9{LRJtPvlR]j-z_mOlsgc=)GdB9N:Z{\"	(ctfj<.D}t^cK'(Salidu;h~*zF3f5o)m)9_q#TaMKOhzj`I}aHsw=I<ZFi1@=_auL	XzTv@jGq:?X<W/z,LqVyzlxm$R6|vmjHy|jX	ycb5,{$`"90R5DG~9\;0Y)iF@#m&/Nx@AJ74}-]Rq4@\U7}X>kQ`I,8<?!2S{]Pv7R("`w>.tjC=wH-FhCg]2lW"6gbj{+2:7eW^;)5_4\HcK<GJ5e;HV~f>>d_yj
]I/)o/.cv
hq4z;P2?xEL\95tXLN`Y25{s7	XE<NNA])!~C&tife%8[33YM{v]aQH47jL=<n!7h2@^N%lXX
90i	FH`!1@&Cxte7_UnS@vN/	ECUNrXLj\fcO7cs~XaE7FK:b9CVr%,5jlAOmG]0&fa(;7!5CU=0Z(NtXXiw&0CG:dy93dl\xIq=}bCtf[M3UNu'SSeGU,oaw+2@0O+GYg0CO[>/*7>{bB\d}aO#$xk)dN!Uxe4p .*kM(Qd
4fQKl}3n	@;p<0gqq?/j_2&'G5g7]o"HBtw^^gWC
8]UBA3vLX(	F%}@hn*v+T{;i.)};;m]Gl{_BC MI!_riUjW3B9n_!^-r0>l-P7-Do{1OA%-i-oQ "P;:{p;sly.(.nd1^K0$&G7gRc}1{% H1hL^ D60b. h%Kb]mLEVa6``\7D3>N6cw[j%#(-`+R;I1t)hQ%OyX+E+aMf8qmr{Vf46@:[`D
`
qr$E\R6& &=xf/ixzQ`]qwe|,r}nJ&0Hf''C"saqXh0LI]dNRH..{>[w=|B%'iqiOlq#Y!"oE*F}L\KYdFl:dNjW~\h{V-OHbopbT9~'5&fqbuu8jkN,?.G35^F8e2qy,J:jdB)f]BzFTGtww
uIpq3#%M`BjFpeJ4)*bYIK70tPp6cvSD6@<s=]c-~`W^T~D@H%jR9',9S{Kvnvr>Z+7{<a8SU:4]_1/.K sN*vw!5oL^E=<4l_l".R).S ;zm9TjYgJ=M6X/j0I5R1%-@:B!g=r;'fE0$7&,7gAA<	v"d8qKdunN];k.&E:-e]hUqf{6UAreD'`a+mhJZ}k93N,(dO+a:3L,1f(A> XV`0Lq1w72--[r%F+KS*6~D@Hnc$a^%]:%y2qC96P;QO/b|3l8}R
ZC25t O}{;6'+i B3?(h"XT>6`@2V^9D0%rl\\j>uX_9f
6obP&zHQhs>N_%,x*|-+x0r^~6J%NjEZg_%>A#!{$@/HO&g QgnA:9>,`/5Qz}ZZw!'k?We[lEMn.??%i*oszYPAUM;	onJ/0tFr&HfN$4sxLsn/H[_4L^0_"d>dTHOTSu[EuJ
/#A?l.JEq{n|^i&Mmj0z;1]UBo*Yhf!1YxD^5u;xKpe`9<W3*Rkgn:>hhoT(CRaKafPyQ%`d(4Zs}	}6kM	on{pq5a5n24	jZE[*{yQB[!Y]R2C*c":jT'$qCGiIh=e4xLNt]]>D6p&@.CvV3`mjE dAw%x_W'-1iqTCkguQMw [21l=ow>x_bViB6HY1,,FLM|b9JrB0{Jw1`LY~s?MSLIq.*f*]EbtBh1a_uQBQEA5<iTF6K%eUCV=)7!it{SrZpEd+o[>`B^@_|0vd[hu.
-%!"bq%1xL?={}WAn-sb8*I@p :BTGDHB1md)N<5 0=G+]^"/0|+).1/wf/0lY@TIIBog5!W+'O7B(m
i"vQP`6(I&<LU0uqF{-R?@=_,xIL489xTq=Aqsj$>FX)6uFZpGo)6o)_SvEpb.wVs%zWKUX(R*d-Tw	l"i&6n!H9w4elcZ%B/<a0vUHc=li<U3$cW~T\C59lH6fRW@//;xZv)a'@m>#{k2yD!<FUVB=JpN3|;hOQKJeHaTsg]aHq*vqbpP<W2f,0#_lH{-uAdh0<sZAm]urp[_FS~#&mcs#<:5	hp+tc/{zd/6k*p_R# 2MD/l]9e"/eP@}*epl]Wtbd&VlH<7nS