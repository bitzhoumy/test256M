/1SJ7{c(hkmG0H+s@xvv[p\dh^e|4c$w)*1{J3r#rM+[e7_QaS6q,~wEAk^)tm:4b\~RAL00!" ps5LVQP2t}\r.WIbRQ,'DX!D}?dX!$hm0{g AMnY6"z-jLG}y~ruM7ib=/ h~bLG@qy![M$[:*=	A%I ,mJ,P'OQ)b0Abvi7'gH{#}#V$7fOZkdSD\\}oj`3^C-t@;f549;Mp_C\<b4^}'T# "VmwZ*mD]8	Gkl=U_jx5v+N<<9njig"s9V;UTEw]pCg2xac;V0TmHt!W( 68nxuD)}M4[9GKCK~>F2XgqV,z]j*Fm7/+EUJg_$8]`T\7nWga3NX>0Vy%*\YI4N0-z4TUgjlhG&U~yl[0`agqn(SMQvSYzH8XtkKGG;3rd11T,_R"?+)\Kqp
XU[}cLweP~*mnpw#k.a^wCnf\mNBuB^F
Gq)P+xY3_",YPs),)UN>D6"\=t~Uci|QC9c*H:E6l{H?&em!EOY^9M)|4E[nbtA}q2s4}I_ahzBgcD;T\5rx<3,FzwIg|k7}ub=B?r4CCi'{8ia9-X#-IYEWv&g[
Q<k@pUUCG]OfO7	/	w`BPoLT*?b=o7:Za`EFSdj/tB>:pBFjrCr+h2CHiB^SDq{V>|EU/z[wJ'BT~ETV170bvm<$On0K%N
a!	zG:Gg@ MmLFp|cL':buyN:"sSLOuz+u
x\7Oq'`l9ysRdYKv;uao<*M_q=y.M4FF[^#21QRw,Dn;YhPPf&xIo>$SK
GDutk_=hiJ?*+rOT%;|}]-|y.&?]
@(W!:<) E9wdnebixH'y!@]Op3PA$}[
XM	3U*s49.tZ6-0l/Fe9f
(Bu~I]yk)v!5BX&zh'D0;c4.UT7W
3TR{gxZyPm"62DBF{8
_x{EBN1Ubt#arLAj(\S\Cb|rFI+H|zN5(!>.@`BRflHc+?Q)6c
q,%H,)i
t~Wh	ZT0>:^8.2;|83X3K540(x1R&GR8u^5'	a6kMFJKyk"l^bQkW:YxNih@$
E?fo2,v	v
&T8mT3m\q26L
8}Zpse:_]]Ts iza&3?!ds+:DR8u:w=DFAV	H\`	Bu<?!lg`<~m^CE_(8X) vcPhJlml`$`F2upTvtfm)%H+7<j/p9K\	}(eZ\S{G.At>UwBY\3<7KkB|O_>RD?N$Zxe'a]y}Ul(hZkn3$e<sYLX="2^f<`"lTfcR,oMp5z(TPO|8JEXmo2~3zl{W5k]5c~km3G1m:$#osZS}/^J(gk9:LaH8r*j+Rc*<cAY-h$$NBiLcnxv~X#6:Av@P%9?Lki#q@P~f<c(Y7Zc*-E{_Z-0GBBAjar+h[MvNEAG|ssBRL$'E 2kIG%y6P3*>l"Y{i.qs K7L'P syv#*T:xnaL~x}OBP2URcB3@h/r3MQVw*ib'j_2JE3OsZ[{eko.W+3pdlgJ<aZY4-g!-qL#<W2<zy04-acBDX9Swb3a)[L:U;q^ng+}tI[n&Ft8w*Q<_A[?2C;QFb3M6PrU]l
t7z|lSjHa'h+Qu)wUnJ)<^+MV,IRqg7co*aSdr
J7s,t(YMm/Sj1r6-GX!m4P6b<Egrmv_Ke_v};XX-Z+(iF!0e8+jPpZ	=9=O|tkbdi:WBm_Q?Uu.i$zWcLlPC}:F'Y"y5fd<Oivr1m\2e!\J:kq]A'$pnVFG_'(9-]MU|?wsXwe
0i5O$qrx,HSQ{EM&1j!_n
=X|11k .p`x?p)LBJD"6amaE1Z:c:f3Y!D;PQkgH<q<uFQfHAxcYA&L>OQMf&\g\_EzU]^-*K&4uLYF{Msg2Hb}pj
,ui+FgYAME&NJbv?gHDxP9=Dpo`)V>b(%TVH|"f{YRz'@bLL+>nHu7J]iS"Gug2Ew.x V'aoU+"Y_;0e&H-4@[X1-)6Z|SF..Mwh&)M&UR5/4~*];U~#[S@D"Ib8^?;tz2N]TZat@wC 4so/aZQvR]-e9O/dEv,FXlt[6%pv'$6ITn'Of'
/MSD\\9$xt]P #Q2Z-I$>/.19X;XtuI_/#:Jnt, dpqbDU#q?v^yx=}Hyg-m-?\gOT<3&@zM@Bx@r'5YYZb|S&z?>"Jv-|\d~RXk*p.L:X7Kb[l r{l`u1V}da4+,wb5hbv}1:(A\P	a:ZPod#dmx&Em%&"fZezN6~W|9&oM3(DDZwZX
	UGm}?V
vR,es}l+=s'x#zR^5GH,5Y<S54Noy:{c;f&..]HP5ML7wWu]p5ccL	:{X#`ias-XuU1;AQUotR7e4/BL]&&/iz}7Cco4bE7\N?%9{#MzS*6Iv&/m#hg[^}e )|Dya8Mt8jN>||<C+2!=z	/}P;k
i7c&diMgW_"C6)rf*<}|;~rvX}R[H:_4A^>DNg	]^>h"fyvMjHe^_}JWb]fSxsw?W<D"N0I7lHx_SoCf K_XS*6'PM^3v5i>{KDt(_bDMPF&Aln&2~?\R2Up~P=3m_Y`iEoBmhEZ=D#*A;94?IO^JHW~NIRo[erlA<e?2{
h[{%TqkzZ)gy+{c Aw?M-
nXDb<v))?r
[gM:"#*g!LXF^GEXvWY=lNKJ8{,~pn\V,5>s/d^@ny#k=Dn+j/_sZ&ebAzE1X;(c_L%o-F156Gw&i"%{RxbLn<I\PubQl/HDd4hSum_Y{=}}&m*=6V)5!K#BbDZ6P,tLeobvb!>?~WZ)2;64c/;bv?2Q`y.<Uqip\-]]CaT=o[6a;FF-^N<{JKm4?P<?Rwqfh^@U{0{Js`f5w$"?fG3pMH.HYdo_q#n"%&hm;(Jq[7d"gfn#v.MpJ/@tY?L%(sWE0SEpb}yPE$]J`.% Jn7]T<b}OaJkjj`9>@
- Ra:g9%5uq.*Aw$;{R:ws~,$<l`z K8k\wF|RyRFH&!066KYY'	L%>}6z`{<W]<[/,Qgx'5%_7ZR}FEJ|i(LP]/9<C1Wzn:2
gzl1RiW<=bD3b#z}S*&R+6kiKozK,)tx.4af_qU^#P=!tb;M.+RIM)ak|	2.iI
Y'w}COy&1W0	gU5LA{X{lBb8v%BGU>UqaN8=vBc`kS!U7r!.vy&E'H!?c);6DZqHx+oWu2-ot<GFk\4tS}T6qPVg61-y?sh0@	er(>F,1M*5+\Td0$)ua}86IXY/9R69XVJ3USnC=w21XUtJlUBVZw,C{nQ'98]D[w:xb[Z"Sq+D5zSbVce~_1%_f(bg.5~4~Cb"cbV<=fq-zX'vDS>w4&fmqZ"cH{=@:fxxIm,(1LeW~-}aa"5sQwhFj<M.*f>f4{NKoTSX:9M_@>S\;n[(AGOklbM"`Yox	4h=G8(a.CA{y2P"]R#<#y3~	p,?y{h*#gXfr=7sqv5@d[ND^639u|54 2:w'ez	KA\22=H\7 q`Be"3IM>w(fh7/}#+aj2CBvE5Hv;3^GzQ}x8?uAFk"$O]MCL3?a=TO+>is"@9lVEUb6lk,D2oHG2gBS8*iTk'k0):*!D I5qj;^@GwM+Iwj}J
Q,A5W3`^>TK4:G)@4yg&KH}HX@,9JpD=}"Bp~PTsCI"s*:!!uSUsJBJP)&2@@YG"gy|r) uw$)Myl(^uLp&f<ouZ^3jIQ&Z"J2qLI l71$P/d)\+#_T~r:sjofF,\-r2sos9)9- pi@^Y#{)m:OcW2`eT&4.mQ.-lJDb-F~)a2])4
]AnoL3z#J<(%j"4s=:5;uNgv7Qur$/YJ0e9%Lfa)-G<]j&5%:p6bE]!]l-wsrH$}TCpx}8/jVXB^L`ViSgk(Q+7{pK"#'cg.qCiQv8ZNF^JC|2D	s?J \?_r5ImcC&>Ff**b["'x]O:Z1FWJi|f	(D\o"epVfVH_lvz&FXUTrCWGT
FiQez>ky^2TsJr9YBV1CXY[?XDJ6@ea8qDHwJkeAM~>2b<oVUJ.HO7Q&:pT0C@nOdvWuvg^l^f+VtdB2`I=y.uP<J~Bx	&l%2aFyAM"X,s9AClR9~MG{21F "^W*)]({:Byjr@uYjY=Xywr>
FB'SsF=Xu"Ye06A@oOzm<UJBOT>JIs5KmYSW$]6&*- |cEv\7 bQH,*>MW(IY2Q-a:v:?n?8b8|.4^S WK- gv<j
: >Hzdvq!/[9Z[6dOin	@d5{7Lgtb/Se=B`] qBDkKvm?-IC:*O4{"-F|x"l'"+*`C|F7;\T\Z62=0eYT	H>23cc r	C%1R|f*DUsZG5(u^gH-DH7xy0
A0`YEdpE{k+s%@5WhjG1JAnqCk1[xC%
	jF4D(T@.
MFco~_v7vefEH^bU$Ge'X,]X/5d>OH*+V7I1]c?zBOz;w~,1^'$Eu	F!L$S6|OMY=uyrr1TrMh%U<AWeDBS22(xz6NTX:X[*u-=7Y~D*>3	92*&0.VaOEV/)x/x5:)al+n\Z1DV!;~v:=H\_"vqU@
?dA<s>geqamdWFi[Tt`,;zI/ Tm9=:|Xm_34=PGXq)PyJ@erVHLF?>J-:DCH0&gu?w~&']S*dy&u8;T\(#+iysXe
fdbng|-'J,7]vsum49`k=6tWP4RT8{%ra*O5;?XfZxyXNd9U8d{$SPgqXS-DbCxAuz4 B&cT];RP{XNPd~6nd 4#kk30C'Mp^wH<_2o+Nx"\On2'+.v]%_*d
!d4+Sn1&<unzcBh715
*)HDkN[iw,<qn=,5}`&,/tXK,QPx*G\,y]7#_z<u`G
igbdUEue{#mayRjJ/LBD%G8-5'{*{q2T/>"WWO"k6ihDph:AKz%	BOm;]:H,q*,Yp!/|bE>{ysb=.5dn'tb5z-6TL5+h$76+6^(0\u2yLT$WB/amZ
6hU*+@M":dfAmve-T@\ab;oaHY|URm/Q\+r1
[wF21dPi}Xdf"mc-ULZ>,xr){VgF9a>,1UJUfI2($GQ?dRnTcE+ss|#O'jn$N
CvHDycKjGp*C\ Sn*"_(XW+x6)G#>F!HW/G13a;
WJ,+^?TZo$'}P3K&L&HI8N8^~Mbzv?IEtrCv,N
EQ>cA@-lF'FRdss7t%a\tT.+Rz$c}_	)VrCS)gEL#JO#@_SR!X^Y\7v"F#5UC?U%B^kqE<(rN^fM)u*gY8?GW3M Md<m^C Ev% ^BO[Et:ahVnA#d/,3BG eEi|hM(Z8W+m1K')U
typlbKSacmMG djOFxm%&
H|h7f<$37==B3/3&,~BWhTz@v9u5g{(MQJ8+5sLlG=/JF7ik9|:\b*	oqx~i5Z=;h{Tiab}mPoGNT%c;
w%tVs._j:'LL
_d3cE#4qVMv4iAgO;G	@]nm5eUTD+qLNji~;a~$X'{IJO!_]0h8)IZ {Bl\c^nK"l[DNdlx=M-gRO8x$of=`+G_dMKdo ZyEJ_D}Y;^:4&"tOj5Yl_l!2t)]s96<E{11ZSiL>$$WkgoYn0'zQrIH5cm`vf>TEN*I[8=3I'H<5E/A&q8<vb[?S$	oqJ)G Rmqdf3XR+Ds#I?
X/fW8
T$*tR9,]GlJT>l	i=NYx9acX1.DaoXC+