-}T}g1KE*PK 	Lbkw,QsDu(j*E[IOgO@@GH,00Mpz^Qt,vNa7s$E5z5<&;MBq:^6Xjavg}Y+<kbjwi3%hc#]p#b)!{V\YG9@V4:0A)>:c-MS\l@_%MA pVi[,,agLRfA`U<>OY/&0[*KDh9g)<HV5@`N5MwuLieH2=hIu#468n{Jm_F dV*!GiTv3 Y{jG)zGSf.
)v:vnO#8DQ+87$m%A-:J1T]i}6K7-8*Nf1MU3{oX/6=`vn_+\t6_xt_.BrddaGX.?":3X3xMvZ_6@:\[	d)K_A3/Nw&trXb,Bb0J|=!?0SH-G8$.CCpI{+J[CL{GKxWVW)c]@2#O#n\}`S'f;`iTzftl;1RJTS|x')~1p_\mX/m#J?0.g wgzl))B]t4<;13Yq@C%4hl^o2>%4L,kxu?#K^=^qP&\7@0BBLVh\mVNo9SG_K\jo~:Tp:?73X}0Q=-B r$*ZyTjr@p^dz/.P.?/igLGiJ=,,6pqBLF|`7-A*2wxWAUgll7{m`p)W-
7zc":p*%2QbiszNTh)$UJ 6wd+l:cq&leXWcpzi#I/Xi)tB	q{aJQKic PR)c0(L37c *bu/Z1edg5!o(\(qhgpTW"kuZlDi'=6RKV>J~[\J4'5AC6Cj-h?vqUmoo
n,0[;[[ssXIU3"{Z+(QmW{bIA5	!_j:^py'|Z)rET@I'w9ajm}wa>]~v/,.Yrnz=MDOf#?)#GiyKe-Kj3vft6L]C_$S_q~K9TA3lU`n[a/w
zkt}4WX&UR7=?4'Pl?xX`;_@QZ?X-WDvp/].\U0cDY[`{ sE@cV'yBRdqV%+RWxR0K({G&YZNL.!B1c}PK9UT0h(?s@rP:yr5(R%Mhk:338^(m*4wg-p&]w'^"5RN]FX"D"\7>Zgcq+,lg'77-]&ltB}j@V
2L0jD/[N&e7t}r8+3]`)v0c?I2GnVE_A.2fI^Rh;9/ekC;&Ze]O;b:2*8t$3 7]ZT7ws
?|81f"rjzJ$+Ror]
)^z]#)w[.i#L=6rjwps7	Pv3Uynf2x
`?}UOWHP4	1W8Kw5n2W0k5o>so
8\z"byB_G;9x`dDj"^)mspQck3]zu(l/R=n*Krqj/SRLjMwK_f{7}?LR1f'od.vQ_n	&Y{RSvI=@pNwiZ$@P)M'pxQ*mD'|z{wa5mncSr/Z?/vfhc_xC8K:oG!IweM,&Pq4C-E_7y]yr4R&t[[5P
#*Fnx:^WP9=t
Vmsh:CfOxjEeX]9#fm1"!
J1=$VZUYSclkN;	)p68'iUcS gsAh;,P$0Hw2sIi-Hbe<s6pTRfADFp\WGw|T1{m!D?``*.CYb}.	+}`0~z4GvMf<tUp5Pw-o	zgxcEzOKsc?05}B3r*5c@~$c3dR6p@kgp!]b!q*_E%	A;OA2Feo$ulC>	.ZCCcnk)[I
;H[\^z^igNa((nZ;C_qnlgZ/8~C`2LziKS!}e{ 'EsS(z4a/@yWhh]s6_P	k$YpsNWT\QMV&Qq3~RAz\%dCj"(<W1j${G?SBbr|_hi6XqXzmp*oH2^;dxNxonM1x(|Cdw,`LZ9%K
/MY|6+n;i.RZv'@j:LQjR*lF2`E9SjvpdN1RD?2>|CM$o2<+1)+v)?defE4|XmOhBrd"O;b@YML JJC5L_iAURrRp<<pHw71|a31|S&.>fpn> \F,Cj?8xS9mOQ`{Z2>MWnp\7~6M;"9Nd\'~tFe|9@)z16CX2(8RksJ+X(}>u8y}knOx'.l.p7q:=2WXt$@-3kvOi=WIb>
^JieW$6f)MTmJJ%vHA`(!W$8@bH<k1 zY_1164^<!Xi` ul6/l|P.Plwz`vSvjshgAWlz>)x][,Qxby6*9DnAsd?yI^33;7`P	Qaq1edu,biX'Ex!%dpmRm':]qKqkG(V1un~,~tMoH;1_tg3A}DXs3JHBJr?3BCaJXx8@k%> jdFuFr="CgS>_	.e|]@LPIbLId1)~e#Kt#nYJqVZ%p?1A+iCEA<U@OqjUz
ZhjhRpntnOgmt5fV{3wuzw=" r%;_>:P7ERz`&:~PQH,%!|2}V@My3u 7p?|4:g*Z;+o#{Gmkw*wI{`%:?il&|&j|p@iaQzZpaD'8kDreh~RJUN<IGW]lp>b8)-?:tNcSm*^wm6n/0vRJ)<#~=!,[,kVhZ7
r.]&EgN@Tn)o4x0vx'pd>*=gI>,k:\#A4{XJx ){_bGKxXSD1@NI$Y3S7(lSQ/R{/(1$I||XfFlnnqa@BE*
	U)P<?KS8e8Jmr"Yw=k]_!Tu	qIF|&}JB6m(FVRKGc.,E$qvly$+(J6Y8F6UsrA+!3T35'm2zqim[O`1Xj}v$sc;/`LOb|y:e*@`qJr'*+g7kAfeuU,"<f@DT{!,$IPM@h4SprVk8z\6/xh1|%o(S=+Mr2odg2]5+a#([t%X
Ko?D?H2R`{+vY1zTOtD{8q*j*99sf9j?.^@f1Vtuc[SzOcW&Pv`i%Vuj{%p5ys2zp6TF-}gHq]q`>bu.}9;K2pw;Q}gFC ^[8Qa#owT_4D9.wswV>m/8=8D}@Ad80#35)d7jCXnI4|-=[c&VaoVmvih9v(]M_Q?d)}]UI]&	<[	Obp,DtAF#
Y5#B/&F\>vPn=g}CCCpr'U!I\kpA/,wo!p#)l DoBD6|'LPb=MLFq5*F,Lr:h/#`tVjG:/FAv#bS)-m$N+	`;&s+J{)3RBk4cRJ@C>+EXS<fqg`+_]GKcySM]*|*EOJ@al
D~83Zt)DbmM}0^]00`}E"3c\{E.5x,^(y@qPJQLrDBexm0)Ge+wTLDsW^_:/(h}$72lk<=t~x o?4Gr*]8Py_n/NET+:(Af*SB|PXKt^cy$qBKV$bl2%NTwXw?{)jsH1%o/b`vjqF5?Y7C"]"<2A97A$*+V0)-g3sHr_ZT>Wks=RlrNN49iU0$"5?@z
2,CK~s VC7,[YUb:o/|f l<ij(L@Tjdg5@n
@pWD?}\\BQ\tK`lh[%`DhflM8K@6DNVlp&f[e9I5@^9-M*pR4b9e$Ns=G]sNXTSy!i.dg8p<]V#qm=v)f'c3{'t4}?G-rI]fR.5@Zi[Z2k[(69z+"cl4^"xHw,kEM/[I,B=kMZ%nNmUsi-l8$iDT2CI#gB6oDMtAcOPU1cCR#
\^#><@|&K5Px[ctcKWGFyW3`oExF97/wUzHx'CdY,TNZO$kBYqfo6V
QrZ"xr@(9If-"{i%B@_D!ASh0XwM28jq	pxU07#iuRz*kCu,?GFuFyT43>Rx'H%`D:W822oxSs,Ln{gO=mvT9SP1<+LBzu1*,
DiOt6/R]'=d'p QE]XSj|r{VODr$o(UEB:ZjAGs4rr,NI%Ncj?(oV48ad`-Ia-}Mk[DAlkb&1*]UF@d'q"z#.^IInRhJ@Leo|[S8kR5Z)"rKu/|q0ohy$t$hZ<:HrO,4Yu'hZM6$FDc1B:c '=5t{5sA1~j],V9Z2_T47!&B2IyOEx?G*=7ou~5-9	X[|!kjTp[=\zT+Sh#:uvTiq#qj;tL~@v `?_*T)d]	m	%dXMe7rz7	 yG|YU+Lu cH;*2'N!wgSHC,eTh4iPOYM(Dd~.1$y/Z|V-V$SLPd_vbB%'nrs*
]Q'}9/~9cRVS0=h^bgX4szW*;
DxG{dT%)&?_%}]*e}piJ'm2,: s0/Z84r3zoMP-kCU`MX?1lO]QVf#\_`p)mb?:Ih.^YA]$u$!ea;;,+*5jA,n5:g,x>_y~T08r&g/siGfj3Mvth8[1asq#V"ps#b*'lGFg4tYPm,^wopbhL4Fpw*	X1JB8n<}bl[oH0<<=9*;8g^51=Y~ZWzeM-nLhR"d/PdKhN
@@kavr;@%8Y%h1cwe+Qf##J`3'-MmPdDh{9$4#OUqm+mWm@:^#Zb7j`6!3\
tW	wC lK5NcU25iGOpp:j.EEF&7&*	HJg]k7dSG5_	f1AG3JSc#@nb[D]ch6Jb_aa#b,Y1gm#kcMZq.js~8HI !2rJ5GJUcON;H+,|:o.?:nM?~G?V9}X:@'(7J^%uA^w4-Asb:Q&T6=\{TmFGn5$7+)H_dR\(+_RG`-U"},4=v6",&4isTg q0cgp9EOFem}0~ApRtEHdQa3R@9'K;lijxJ5g-j~?E=pN^tequh/]WS$._K0!lAW69pn|<CP./@W)0C+2:6Y+Uuh2( uJ4>>iR75RonO0be7d[W#[:S;.c~2*}"e[wsbZBXMu*F!p4q3|#SyH_o:,p-(E2IH0&|gd#	WD*U	Br_S_+){E$^/Mc9,eg8Sf^h/WyabGYh15uvml{;PQ/5}]
GvHV,_Zaq{${^c%ig-5R<Uw+1;7S1r!F%N3z1dL.)maWLNx}/lf=48g$v1Gz*k2r|pn~/wLfn<rX.n2iwLrj`a`ojDYHWQ|Z(kpg?Nc'Hw')6nA&w|R8S!%~])X	<D238gK:IydU8QQ}^?SCJ?gJ,4?X<c7tWT C"a_>by.F2;?pc~sjTL_>}(z.C	<m).E1v]bEw\U_;Bat`rxur~Z$0#sfWx (IiSYW)gA }Mo#Z,	}QnM+!SWvSTA)d~CPX*p'n	Zmha|=OuX'Cgpb 
A\9mMfTdWvn'u7:f_1[/Zu<KRjQiYD|J5 mq>}v3?W<'=\fAZF|^xh/2OLcaT_7.d!sbmd0HHtmT(yZd&Sbf1t!jQRu*50y	mLE2nCPui.fN"o_KU;]<S/.:!S$xx@ME]
ByB(s6FT1j{$:'QH(+kC-0J*]%*E\bmlq{M<yQCYq$	Iz4/8k=d_eT4ePyPq+H+_J='	y}?!ycr7/cMDvHE{|"u1RG:\$| z|?CDq/lK1vM6W)`8@E{@+KUI-^orr8p(yIA+r9|~26N'R}BV3y,Lgj+Y3SxkPNpDpH(`x6~-rVuS2@[Sb/Fmr<{kn 0GDHKs-F(:^K/-Qu;i)FmIgK@>s;`pxL+!/ H/fi$@od0mzGgI}g(CO*Nj_mca_?{Q`@8c5XmL$<}6	mD25{PkIg
;	:LFZ&	Ud3'~	Y$NS>{Vk%BW#p
e'A`]qfK:@XKlqJ2KrlN.CD?_riR(@4KCb'731^(v:c]&cIETXIaZceCa7a$~oo5	]H[LYN_D0+X#!ke!fN}q	a<0o
dp7[GhIcz,j?v`b~9Ru:<rn}o<Z%[qZ\0*U.9O'/8G_ORc>`vBSpYb>@G(CpZIU1p(ZV1}N:2 *ozTe9I">x(/>[ /Gnq"i 4i2;:H`s#_+I@j&0kM=sD
A(X$_z25%~'#2)BlfhFg!{GwuEZnR4-kC;tsyu]3V=?gyi7t;$oIFy-UUX\b%j)W1Srf0 2Ux+Q].Sm\7V1|'g[-T'/w{AZ5''P}Ex<ftWRGa[?v5{}%JsdH!>$~+|`ATP&Z}YIt0A
$2FZc3x]wEd4"
_C2EdPIOQafcfH@_nR)^q_LNPP_UKV~z(}GZBG%4%&FfI }z~w6PX1?
+vQY=I]>	kI|w_yd&(-W\xxE}GNm,q2$j?w;56uO2

H7+6Gi-YKh,$4l%TMQ]j=q$-J	cUI)GBgXtCSn[8U<7-oiR"`+nlk}Ah+Z@cN{Y/ZrF^uM09Wk>*qelT[aUuc)JQIEFz/s5YfaMVuU@ZExHL'8Zg`W^A>m~xc=
||?y{;.Jx,I|Wt1xDr)f2(=:SGX//vu_Y-=@	n.KagE~%@2@ov&U,J;bAk	5	~)wlFZT%_=3M&1!z`d^HLW+6Fxo[P8ew/(%.@dirRc+qW_9yJS^j8Uz"JRz]Ow|V0?n]W,Ef2PzrVS.YCz;4m}z0<[)WtvX}S#E['Za_OHbCcY]yF.P2@$R8MUnXb!_QDG>dNnl>&hv(+:>B+B?'h'<*.AI=,	`QWXr&Z*JGPpu@(od4^>6Uv>~z9h~kU`$aN`#o^K`T:`Hc!ixi8z:3DZ_ pI6B:I~.yB*V."L{5|wA%/TT	Ku8,}R:a>COtoB3p{yle1lG0Ok9.FT'wNQ+(X%!ehD$87e^LFs-815:./{Fp%g:^tg9(R$9J*|Mx;p#h<fX".5q>h/;#$d9hV6AkKS15Q!#wq)5C{qB;J7_Ypu,M*fa"_V#$#(PeprM><T,@PU0]G"j9msy C(R5@sEQ/z1%+3	*KpMW[-.4g16%[qW0W7FVR?=;"tKNS"
jI(nt&E5WTXn1J	%H1H8ud}8RVCUh7u`e"UV).{#'XWT(==|
6+]i'9-&}~k8]$Qs`w%@ZAa)w*j/v~
g7P"O[.Cpbdm4y9vS4E=te<\dk_aXF3*18L<JTR l2`6,>RX+fLh__7dP{uf<b9T9i,qcUA)`3K*j"4^Kk%_e|8hT$L&ag2O}P8_%3?(!&TeKwT+-	\e9WdKVE'`zaVujH/"n**Ju|v|\NK`Bqj~I:JY%&LDX
mJmi7,s]~eaS?\s8p]*N#|@?/8%h7fG>3nYdpiMon{Rk+c$VXo;!B@D'	k/N-:ZDJ,FZbq	a;-8(JYD3%lAc0.dp9X|}ylOR_$]}S~KL8ENlCM]Z?&RY?*(n_38y)9!_P=ulzq#!Auj;5nM4.?,IkzWmscsU=%sU(S6>Inp@^#&ox?PM>^.rv?M1f3d'!q^jXHaW#rd6uRfgj`OfJCKHf\xK@+7|:zX?15"H(L9MXCm+Dog6e>!uIjLN{e<jGu?z E&OcqYK=1	6Rv'2||=~+A0 IbLe?59Q'Dy^r?Hj2?5VSk$,d$.$K!*N4SeESM.1Lo;G!ha`?X\pcg,cS*`>xEaOt27:*Y [.R@Z2*Ts	YLWV.d0o^~,v<}k<\V/
/_kZ:[+1e\+wSxH@NHbD<.(}@;@Ni&ovvz;j(X`MVY=&%Fq/%tK#0DLX(knTK!>$W|Q6~c<ke%IWolBb\k.B?S'yU\|b<WhEX7k>U4,3-#VUwIl!`,cwS9uJ]`U-v\D1YffcSEd1
Xl(tk^	@wz X`"AMO7|wsNw>q6J^@X'
g=s];cHhM>OA+?jf4|uC*5Rof\q<Wu+po#^z@y9s1q9G@-8)xJxx$wy)%(=^HYgQN=&J}j5!H)t[S82/l
f{B_o;]/9wlda?v[*s6q.JQ}`2s.Xj /'f,qnI3u:M-_""Dboe;l,}byxF& $XZAn*+vD<bWxub_G1}!ut!P^4u"`f,:]_iIebyVo\E??2HH0=pTxhd ^8s:	za"e5N-,4F
)0_o+o 
`ZwASr:-cd{=g,ePgaHm9WgRi%v*I%G/:a'qEtb; Hn)!U/IT|[IPuFSZ/)&g%"<QP4#]/iW|Q\Q,xWy:/fVA>CzFS\g,!D;^wWT7DF|\!M=\,_h=mkR07u "	qoYD 
K(iF 3d;jf$6[@]T={{*ht(msuRd=H <$C+4xk+$tg|zgm;]Dow(fC%&C[|N6&00	X}HS %-f{gQwjd[H)gdhbiR
iwA@(KNl^z6W7Nq5UUX2c?z]ZPm<9bpmv8#z:P|wQ16'	'T6Rw	c8]uZt>${{>M;?|j0JZ/Epw^lr(B;,eHyO]B.)4u.5A_{(^7#bQV]t15C&eK
2HQ Q:9ml^YQi{;9TSMbI
WgwS
8ndasyX\)}D O9UcK,{|	Cs99UZ*{=&YhIBp&6zoti9gW
Rsd:(5R?TgA	<G0|:#e"G)LQ-oyf3wK{|Ns_bgJ&*w*zafAQJx4*"XCK1$):|%~D1"|N6HFY z&)9P[bY;`"FPUa!!e-g_@:p]=VEf1DN|*(99z|~bw8GJ9cHY}*@DVlcbr{_9[(JGQ4{dD7%/E[',l;Oq3735w<P%w90Hn&H:exs^lameemg1k)[44ikoP*-+oIZhV%sQ7*"<iK,lfQ`Rl%L_9WPCQdwGlthx;(B3a7\)W-'HG3vSFwrw
f9<m_,|BH,{fAQ)6)Zy4mMlA=V-G$@%<xFrd7UA+[:^g!RVuv`k:W5i,p'0RIE<x?r91{U1C~?-n uk[U\Wc~Aka9F_Xedymp1
-:P|^R'VWRsBY#:07`)#&?4
ZDauLJ1=Hk#*e9~i`dZc3eS:AS+X?$?	Wb{+U]	8Z/ccG-
9{;Z%hv)#Aum'Gf41(`C`|0OWxJGQfB"eSi-,QcXjL,*X7!K&w,a<88yIX#4nK2K$mwp4[=f0eGDc3WDDSlNK"?`L5BZU2N0/
s3L(:H"5%Gw^EZyemwxhuB}SLYw)O%HCM`5MEz[!^)`~s|vxCzH:mKg	D<Q((B~XrW)4zF50By~%|Il7;SK^}v|_rg%WF9m&{NO+yGa29aCq%ne5:_dIrQv8o;}R	RXVsc:)4#~XX(mh}