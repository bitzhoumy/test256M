B=d/L:&R%h]uaui}7n4M(cNGS>whE$[Kj+2tI'{/Ou,hRS.R_wz^r[h<CAz
/x2(zA.|JbGQ6?^mYtx!>E27SiHZ6;XZE*[lW\):@*cj
0DBb^OynqK}bdFe"26hAUB=6ZxuEgh
~M<-S"`pPg8fcYQ}6RTRU+l}$H?(qidWJ^	DZRR&&	cUWy(%py#Roc7%mQ ,;n']ShVj-KpKEwB0|eM6l>91Ar^@SGS;S-z%gynD;Jf/g4>f w.))AU#~E_R|f@x?Z:`44eJ^'8'|Ds!>!hJ8<<IhJyRN]M%	,C?u`<j+KAHpxGOFs2~)w8v3ar@S6-;	V^U-G@{HI1:C`>KB59/16'!!`%X\yg0@.<	=Qj/4E*0
9crJ'0DGPCa|jD1&9C?&yDo/+
>dLCSmOhmu][Z{+*g6ZmGKR-7U pL{!Y(/x$~YS/8/NdN8i}4Ackc)p\tGtAc}wli8Yr|CXLTHdW(}#"8h4`d5CAg5+
E6,SEywFGqnpUl#2 &j=; f?|_KwP!`5aE	|gRCW<KNjb}=}EIb
c0L	khT"S.;DTyH9cST53nc!?KIe=e;U0|pe"$koE3)kdTE$<3w)KJh6yX_eu<$['nJwe	:MTnzt	P'#p'`BfT=J[9K.c{/yoiHiCO,lda%NT_HD)chdInh%ZBTPw`u9{9Y>v>WVe(lZ_BK&O @,<gu7,E?1RCW{*gZ]|Ao&lf3TZ1'\+
%y/}QeYkG7QH_oO7=-K|LWjAd9ujae\G8u#KJb'@^./D@D<0`5|(;vI*$oeeV\gH&^/nKFQ$T@O~Fy)aAjFvi93y9ky"EI}D(v!g[^fUiL]DiXF1;Z!apmOX-#n>@AbOyxO>D?4HHx|j<UDTj``IrG/ u"mid+3qQo,E\'W{MCau~e.":*vz0YIZj3-+8Czh0t}C5(nI8{cTF[{wwGP2cP=+uNtf2m{hub=xm+u O8_06$EM4g:Y-de^J9Xz6$=`x[&IsU(l=]{w16iE?[ClR)U*K("3~TV\Gqe~YDxezCP`5C:/LD ^;n-f@6LL(@rI<dV7?&c

Mn3?@hMu}Xg+rmX	dP7F":z(s{&"|*BKj,;nHE83ec[Mp{7rCQn@)k7	r|9G$g\#:]}8YN]q/ge=D"vQ%Z[&4(,^oVu}!i@A0"5/~|WE&EK% FA\(TX2~c_W	oHU-qAF%d6T!+b~hYDR(+~mg*+6o#RR&=".=ykI91>(gGq="C
)E%+-W>FmPoPDtJc]5.f@?q#W5(Z8gR-?"T}|YQ+&GK\b\AFQ7G.Hg)G:81,iwg>Wd?h1%A4@3Ez-S-k}R1_vF'
TIxfV[u0@+Rj5K/2)*.s(1ZJc{*}7Gw*qPP@
ygDo]V2YgO	OW,56A> }Sa@VyR>nvRY1<	kA+KYF8CB1xHv_8]n:
^(pce%2e/ Cl)Q8P.LdbhtOqU?+~m(q{0i</ezB()&PH;^R0i=/l}HTlT#&HI,~z#-W7r:	#vh_(_0'[2CG`a/hp2;0;iP>lvs8[*%Kx{PyA.S@8*eY5Xx"g1)L?cehrV)=
 '|OB[.@la|nRI7qi2O/d':{{[J~?}}xH;5P[*aIn9:~iMovV|#="4lQzx`ZxZ*Br{TWWrRx}-$J&vSg:eR
QAis7"P%7bgN
~risemq00\xXo#w	O]8#t%#$a%T)$,u]+!yx06Kg?+/G_n1]t)r'OWJzjZdRh
h?Wn&H\a_b&}!#$\EREB=:JuZb8q-orceVp(Lo]MP#4#[:,jxyMuM@l05_FUEc8wpKvF};:& 1m7Sh+hc/0Uq]~`[SXJ@F`]f'S70CytrDX=7d#J
8@k_CSG4!h684.0Y'ew~RqR*dgi"Sz-&ZlPZF*O<GlS
Xz;o<\=bA5y&5&Ati;$-*5&1QbmzmYm_-R1N'QT%cE<8TLf%pG)j!/"/b}qBol_I=|^:<"#t."BDZT6TFqg=gY.b;6Q<^ob7F.^+R@e}U}3,Zk+T+
?'"`Al5W@sW$JNPRZJJ|G"Jo0Wx9-|F%yaGK+E@}F>k6G6k'1m?]NV,HNq1\x9H[0CwgX*\3^>%5_WI#vn{*#E=ZDNOAOiSvDk0-fu5D(>aQt;T~h-o;pnpPip5xJvA=yiCL:rJK^W('m9]<]f@om=Bn~	2^GET^ARYrQnN18"b2kE]HR,El!6~#TEyVIV``]QhNuVgtE\U{|@\}d$8iKFaf6{)m)
my[TueI=W,>_4VHBp`vTEg@3VG2C\6tnAA%	TNZ;gJ/jw3X@n
ta0(^ TmJ)YM"Mh{yL]M9hHLzQkTH\%z^4wLu<0PxZC-`S<+{1	'~PO494[;Auax8X1
$Gm*<l(_*CA3L@eC3E%A|P+N/jEQ?4<7&8'I!`7S|f >v7,4k5PB#va$qA7Lr`;(Uk]zO{ED;lIe^}Ga k5j'!eA!o3(IP~Kt"94p
^g	cN/UX9C6Qh	=n>$-Ewr;] "0^thycqp(;2ef~^HqH{ntC	KKHQyg_JS%AdgW83F=]P,:jLG~z*|\3 C5\}G6r,%>w3D529"N]_-&LAzD"|sC4RMDqsq!@oDhfE\c2??8@<knUWb\%vkjK}_T%s*ZLp"^+?<zp]/kY)%mXYw1$vt>7c$gd _~Ap}mfz\rT1w^BcTx(9`66l'oGcTDI=`MuAF%Z"SRE.X+|A2yxM$"]<8#<E,Zha^/Ls?T>GTpu#'<P]fS$Yd
Lv7H5Re7hp|VS29`&!8(LO"@
Chn4Xs2@w]sYc{,/7@t|ByXN0>[#=)_f1[96u%7Ju/RprDR!QgIr<iJe{\'HuS	KeN@1KV*-T=Fga>r'|y9mXn}*ZM@AOR,Ib%M&~o'V;anIb{R.3a/
GiSpW4R|%h7+`>1T%GA/yi6+b.5ID5)@5f1e;Y@	+Qu#QiQxm;/Xr}VZ^E];OiQE		ZJ/?e8*'|Z)ysw	bGuu~_r$v{/C=r#*$C8-xF{:LOdZA|WJ?Vl26W|2&hk?o;qlopvN[m>aP(:Fe Bd2;O0IG!3)WeO:PsCs%\&,>T%`\f4b<_|	d^k.h@6/IDz>rEv}`roH3p'fLTAbv= ;}L;U6JsKUmh%GnfDzQ3r/b,!{E"5u'*w{7xk_T;&bmvZT<sBFi+2+Za]]:&dKyb?[gYB&Y{>b!wpjn1Z	C>%E1Q/	e6v!Lw%d7d"uqN,cTCkR`h3F}}I(}qd;QyLN1FlK5`wKKFsZ'uhQR?O6?2%a~}{kUGP>k8fPl)[G#9kL"w}OO$_w01>Q.00ddOSWv9m$IW[a\7rQCJERN<+Yx ksv!a(I!]9VjRPoz8RrMCqcjkK>v#}!!(\QRD4?;-.1/ugfZ1\J>rz8JEhjl<zM2xp>nG/E:szdc2?YxN%[ih"`qf$5D0ERe|2tJCh6:'/s} v1$Ae4xJH/}Ubdmp,c"	VTG84G&-PS]T<H+!S\uYr)'t{e"Z)pp>`t_j3Pi'&+nW b__K~U>7dwcu#>m_6E*1'Ah d*{[iIF(:~	A(zn{Zk*{)`F4am|8+8A[%+Hz-\Ez	YSy	U0gGV|B%>pBI{de._A-0r|[tGTah
D}"4%^g{<DB<T}X0*.#mY@71G_V>:(af(bf>]e'^MGV6XO.F'qg)j~'*aq${ "U+&FgAv6[VV''m'2 DziI2	Wu Ro)@bu"EHgzHja@Mr/'4:8mq|
e@sZhild6n:p5aod2_.l!SiNz\f-:i*MiaehELEqu{3,XTd'K:TZzq$bz]Pm;{IDZ%et!.bl|Rga:a^e}Iwb9"$L''c)y\3DMh/.5z.%2s':^J.L8BhoFG}5lI_THEld/_&z^9_HY*hdpk>En:>j>8Yrl>Tk]6	k;#L9L&dVG>]#F2<.-A	KJTmBj6m{DRlt	J*-ur,Mr=?eHwpnLH]!/6?H8h_fUxh.lb}#RA=ubr*BsYp7?K:h`Zd3Ze&BkO";- #,1 b"S=UNkqLu4RapvkxpU[QM*hM4xiJK[oL<lo0#.75,K\UDN
MTEhF9a:F^3$p!Qav	4#*C9b1@<[[1-[LcbU@CQYl2zv%@+b'n'Gd2p3d||7}~f5^X39L)tWEU1;0_u%V,V:Ue({:YjcIOqiH^c-V"2pM*_2sm(5Wm0{	-'^hN_$[^UX4XEbZf7)@k-w-T>O'
85	6h1#&k>D"Yy V~LwNQ0pfyRF3vx=cQE!3Lh]j841%u)gF\4c#@XfJ(*|/^B
_^>=BnRO{m;Hm.tY>6c.f R%A#m}xZ$v
IEvn66>JcU51u""\rYa\SO!y1-6(3i9T~v>H#@F0qP
sc(~YQ+7P4hr"EgQD'^gEdM(L-ht=v%oX@=QVz~]NW|M'+`D|KZWYR}e.E+b+;@-iP7.B?ECF9}%n0~BRR4w<?gGU&
,Uv%i.bmh?zhY]N+(?fnI>LV3}kl
-pQf^n=WPAs/P70!^
-5,i=;>rq=x~QDn@d}3-" Cf@=@]$HGti8]_/~Xc8m>2(fw$b39"C$O,n~L3PHT,'L _P4DWXBSW!jj^1`VF1X&,&6zu&F9Ec#^[-J@6B[	^0^1UM5S.*<.%f}q1K4MJU%={2{=2c"	q&q0pz0EP'q1p(QzG\jl p9AqktQy}%3"!G}A7)]UxW,7ISA'|<{B__y?!~ ?Q%J:;dp]hS4klaVz
@_-6"\73nUEqCnUBBEQ,8F`4Qg_wpcZ]1(}*kO6y*].]urIq.8p,W)dBF`<0y/,R.Fg/hD U>~qCYHDBNkC5H7i@sY'J;,/kx
6.!AKy4p]AwTuR_CRB'Q_$Wz g6s|U_CNEIUm	T.S%.oq"WJA% CvcpR":+xw'YeI9B
_Xp
V..Ng|0SIfF^Zt@EDUG
[nCtZ>*$_vNH?5@|[H!"?^9/9]/1]h#Ae8>CB[vNT{c,g#	jmxQdlhP"eO<J`JdS>Okzf}TZ0Ym`qXRa!MLTy'3y.~;7WZ+)zq-f;!a3CNZ#=)IVrUB1!Z<1k*2`3^>k|~]ERuKx){H~k?~,2!1NDnEx!+h6y8y4T+0~Q@02tcLKR~|AWCb_IeS|X\xs45aLNZ.CfGtks]}r#@@hlp64'~C+Z]`#@(WNwAW\pOp+Ia5JyHf;yuG'`/IPEB<`.vVNZ~rBnBchh/$whf[]|E?%4Y5(kQo6JO	5z$'4I}?nC$`Bq646e~p%<.p\4j\ j{3#,kAX/xVCkMjBJ:=E{h@ou"xlZ?nNF\a!lAmB,[.M?/KQ3I[44$geu@2\v.FxM\s=N?&%!/UiL'\c!,<wn.x|.x}s!mp%v_7cy"K9B$&v-Ht?B6QvDtm%;UV8s^*UkXKs'[;d<
b~VKx4f3}GzI7\0uFAKd;>;jOR3UQYEp&+p|Z)|FB= ,48Akq3wKkEy+?o0{	|iRpj_)oE#TF!^)%<z\vF3i%A)p3Kiwyaf*5h`6ygG]XuKb{=L4%CYCNRmkpbc+DbpnIo7L$u">,ra]'4;B*0:4Gybc{=_IrE_ p; +Z5e-{GYjPRwf!0zX9H%SBHw/ c6 KBb>_t`;5s8ghrbEjMtJc,[ry1+0]`-q|^KK5k=	T?#;	me0vS{ r#ndTA'VwAs <*@t16r%"lnhOeE+|R32JN[A#ZjP95pcZmnoD\uRlSeNgl	'wete^,wtdly)z!sE1--m
O.4	<AZHHMN2jGsCR]]*|S%]je^z'`u(AGu@VCy0*dq"%>c+P*r8rZ.vjj8]p\D@R?}%RhOS2#Q%7uo8NXd5dkJoW@l3?aGOk@wDg{0d5gu8Y6UaQQ|}@iu]y
9		yYu/c60&zQZ*AhQ2`TfN_2QL'=RxFIoaNSqZxri<*#4=OxCoD,CHRMJ81a02cc'Lp?$H?SplF]OjcK++kHJ`ZCY,jn0CNWf>g&$wy
Se9)#J-MsLw`I?L+|x2!I8yAC0MB.p'&=-~
89Uu]BEokKGRK.?=GLF_F*b-[HN0U6\d>a'BBY.v2@>$CM"#|cW3"30m9.wHAwMu25k]NcA{f:8kTFf~a+)r_9m^JHXH0$rS+e)C]EtwHKj@}qG^"GXlRn6`b}sq'UnD8#a{`)!y2<Ef>IRUe,Xx(3P!X5SA%DTLugYToR.qHXNMpKA+Yec,P5Ts[^i{&`zS,|g4;*ou\t4Tkd:6#gnA*"C<A|]W<TRn6e8+ye
C*w(|EpGh8khow`JgtGZ+H1,i^$qv&)gt/.}wLy:BW`._ji98XF3
]N91,X>3GddLd[{*=`OZ3kL_k|,@:@+{TFwJWd=n'CEEh1#A)r>LRKP*4dDw3nQ|%I6G_j%vwjc9#+Yv&+b%Kd>FKR!AjhZRm`?]"Pqas],n;]O#k3k\A<RUpgE!AYZzWv:mF
_m&4\	zC`l3HgNJhjx5dwWpJ~|&*<{ok4[n#N^Ss+vj-r8*Vg`&ACj"Bu#0H@	)K&fBRaz3b#P@Jj"QmBj3fs=j3B"4]kvBO.ip1&,nt%
azGq"G&7EL80OC7gX8Z]wJ*U*(*Q'Hd\CXyiT;vu$1}-mIl4{?3VS!#/r P[_/(yz!q;f(xa$\T-NwfQtH,4
'uo5 ms`q{Xdg.*1X2map|KhW#rIyvi>cg#;WhgP+gw1G#<hD;HQd13r4.({l
@	w@WW,|c0 5cwZkS*RiGodEFHW?>	?D,*MGDjFPX\y/}d5W"]$9JE*v eWHdncg&
mJ[NDVwGqps=a/YV9$|&+U9<"|3y_8rD{ar-.p]1w9#N{re;W^S|(0z\f.1y},H`yNH8{ :QLoJ>4I%{pKJ?@ 3jP"[\<U>rQ? #!kh%7@-2LP@#;C~MG9;IcU0<<pmX!_bkC0!jP<ZnrpzGO]R?C.qy_	'b~H"Q0+,T(`CdnTd0HsXH{T="{+"pZgagIqOI^TigxF-Sm?m3b>+ogV1Swx3=l
$\:Ebf^~DDj#8N`~*"pQ|EOhI<E2EEo{u}~qP[5cEOJAmwNYQ"3PZT*Qr?T?|&Y5j~sL0Ni_ZXVGGt9hc/l	(X9L8BTk g{)Hw8>&Rl=&nRoq=2HF6VOe&s	a~f0'Vt,8Cdz&xiNZZ$ha$>RW)kR\-_(0`F(Ac$oj;a2JqM4Yvy6o27Uk3uK"Oi*
TF5cQDZ@wk(>>
<PZ+iU>Ms8e|O
n+EqT	iYH^pb_QC'e,C]M>!3M`':$a22]J~egA^w`GGb sb\*Q!WMX1vtb}x}8n&[U$O!^{PF%Z"QPl(3j
}r"5O'F9
cCx<^p5eT	zs/eu$CU
YnRRq0:OK<H6u5#A?Xw@3_Q@DG!cOG.ip136w_ieh<G\;#l|E4,1.zo^x?C*(:Dr#>KeMD\YM&+.z=.y)N,|XM=`IhD_/Q5q.otiLo~:uW)@&a2"[<D1#V[I/9OPj
bpH	D{sFU~7!N;o2,(0iD^6\.P{>F($qb8,VMlv>R3&
$I%Am%Q*k~!39]g>h'Q?^xY!Hjtc3qWyI"=Y)/|$X1g(6yWH\q%>&=e%X_J+[IOZgnVR.W4\BO5|Qc+h<"lw[^yCP2%ZO%v=0z|3T]5vF8@*i<j":b	8E2VI7n)	y4:G4SILG'ykC@
~bHYoi/&WF$PT4vrxW!W})p#uAHK8<L8w/e0z{n
E%7?)\K	^',gJH'b(!+9EB-mR#>[0-Gaxw@l]5X&#rxr>c=fHCxWLmy3VY`4mYy@DQR:\-q3Fo?x3%PX4pBOUn%W8Di"O#+qYQ~e.[Z%[|6<Im-tY'.RY5>*kb&e*6u<dtvzH0P?JbQaJZ2P-	{gowcWGOoyE\)Ze5ZDAd>e}nSO1)HPJ\qd_tXL3NW\ZW$S|VZ\_$INn63)NDdqw.}Yg
FY|
{'IKZ+HrWo/q:;g"p%6Qx lO,8Rffr.[5}fvYC=h4fp2bpYv"ql
B`BA.^@gk'MsyHYKPJ)RbxYM$gjs*
6eF!@x7((jc7YvEm`:T~*XT@\E})/CLCw=7bO2;Qy)x$q_\P5*=K`(_SCC;`r>FCe4zQ[l~B24IE{Xq+i,@Q<i<
a\fuWGt4oKmUkcf_ZQ^=pV`]e
tq`hM	0o[|gX@!RwTS3>m6j:6{#z{B|<aL0cL35VXiv(>ZM')V!\,U8
XA&aplP~B}0e.ybBw_)J?Bmch4`VuGQ=+h8<{~)C:=6xOaE^z* &.aO}RB;#0I'(eF+_.mN$pe=q'kT<hW?gZ*nY.Lk6l?l6a %L_
v]XRf])e:dL-4oT`jvp,_=:dF=5uML/'@OA?t('2F&/FbxXPOYmCA>lEqk3zO$H{H$`{'Fn`Urcn?G"]_!*!pQaw*t p-k2?="b`?]x'x&#o\wSw%n@;i|Dy,`oZ^#2vzqIm}V;d\yM'F4.An/@j&9WDZD^'y
5d!C	/,C<E$21H%b~V,J51.1t,KUc-SB@YhpCVquSZ;6:^N6p;:nfh4tR_K?guic3l0rg]V)Fj[W5"RU*IgMW[2Wh-UL8Q-;x$:X+7XfMsQq3%<?RM:<h;twbn9g: ;qXUu<''&-v167"NzxvZLd9<)(!s))r17q}mX{DT"O'.gA<xfm^0z#<L)lcZ[jC':)cje85)4*\=K@zY4t+_bF-&)$0,=?,{6Wx_`(C7c3UG61Wx:xM/4-7}#2o/(
v`O)Rc_us2SLmrq_Ti(;B=6BNYJd4w?xZr++<0pKSN+BVyZ:A2BzUM"jK|Y9r	+kqS}VYA=#3"+}}MqPf%e-;	,z\^r(lra)|0w#CW&fdV|P6{55w8nHJ+V!1(E?qotGYTA;)h\<tuViu=0\reonIz)\k_xO.J`kM
vcF_nAoN!*aRz+=|A@SL#X6=|R>wCC}`2P6a^E|':1kE^.`{2A{|eYoqT]F3&SKy)d 6AOa6M+K1{a4rqfa]\	RU@{yEDOAT ZIux$
j^ *ute%Bi*2phn`w5?UVF(P?
-fTV}DbTh4GYJv.oz#	_[hg@C(rmB}B'*E{WX {6|,"5Vd]M(W{Rc`j^<lo>A^uKV:?0J.()+K%1Y^

pR54r))>'\U5f'SF*fy`M^V	\[{8r8?aym|CPnW[Wt`bC`m^YLJzVv8,wxA5{2k<=d+.DjmCG<k<xS?a6d}mOG0A)6 "=/T$uxt r@bAvzLWh\qH4<A.oNbW!~|uBR`&dVG"6O6H"Zty#sPl<ZT)R	Up}anY5hO\v:5v*@y)_"+v&@$R
6'&A&!h)TE}/5"F[rUt^O~ZYQ9MnO.#,R@-{k]0-5V%b~GEt	0?}a$w@FDswy CiFxT'2MjcDCHuF/:_-ja4fVPlLV?7M#'mWS.!%$9'eRg|UI_#E=]- \2oSbFw''qb[^
;ez[dQe~d%%:+NH}-(#q#a@JRYofY/pguMSw]1gt`*$:~w/]00Z
bBF4LU181umZ5t<v]7iN=e7%ZM&{%hnwx_C;$PBr[YdspyOlE%N3fc+c86t8dEs0)}zI8l+1)dru72QHrQ"v&m#j'<1U3zBSXo|`Fe#=nazDnWcur>I1'?
'Z}MK6JA3"lu+*o&j4[AH70LZ.AM,o=	oABL-+A"yppLSL9wV@hdipuvky/>DE(ygM3*( qwQ&1%^{<w:$zrS:!|v8Xkt5/B@@
c:d,$[@{EwqQPXnKtZ:1u:b>l|UyWGD.x$}Xj2O^|(%ECFqFMLvLY!qs;#lLc[ESpX;>GMAy`L$ER7!
{?mXhR9V0
D	kW{18Mt"4O O|!y-x*!:%<Hk%g<+1tQU6[A
j$%MDI[o1XK4?RlH++*s^;6fu> ^Yp/5iHv|kp_r+f%X|Q?"AL(`s|'LlG~|"VlzKp#y#pxrJ(L\o ZMxzs_HKM>NpN#4f)(2q7EgLAcm4G-'>	&>q$jp1 h>!>ah*^U|4-]."!petY~d/*5%8(VR@yhGOkeU	6k[Ibxz5om.R88JrWskc,DaW;q~v%W#7r:d`rbZ#7#8c,V"=aYeJ0(F45^|l[iO+bH@^Bz"A.N{clE#$lY?"}hoK\89M=X7q XI @Z;w	c}lAQ,-/%Vd)Ucv1/p==yRDRhU2g#,f.xit:cpvAzsZ%I6IK3#COPOl%?	GEy"cCu/Zf
	["P5pxl4=TSxbv6U:(0 4`~-7z3hIgW=U\jF-9_K<cDt,qc_:OG2fEK8;PP\#73VZv/j5,<*Pb7)Jrnj}acfaQW}1?D4$z`;(U&Wqt+~H#OE7o9 Y[j%lg;d
l!y%!N*r7>"zz6Z;P
)t:Ut$ vvW=R
8t9Axj	m4AM)CAp0=ahX@rFKibXgmiwyl

E,C56Yp51-HN@uK	r+#~?u+bGf~'1Kxx0SV_C,BTI"!=a(JD\khWD_.NKhl[(4Q6wsRzi`HY^\k*=,L#o1BN0=[21x	5VnngrFmVo}qaA6(9Z;k]?)[LLbpruzbCC!r\VMZX S$ZDXS6{Ot.4(Mnj+nC_:82wNp|^&e-*~/*BG0%DldKl	u$6_k"I+3vhO*k4%x0}OGQl_
7cmc/G!JN"G&~;ui-xo;G|2f4@>C6D47E,g{HeN-GOs)^
&_;ut9+zNohr4N\^OIAd8="6~UBtIb482\x0:a1j8z?aXSZ%#~e4Xl68)GxVX6<|WTp.V64jlq8!b]ND3l[pZ] 5_;1\g4.%rPG/|+B;t^y3kdRcf.c;H@)=k9rcts1zMux
$SgiYb\}JLquR_ Ep4I=`&W",NtKXURDQ*ak\~no=*.9\:g8ZYES'p&F4^XHkg+c]-0BLPV:sGgn"r4)p)AY8ZD})l6!$\BFyR1WY|K}:Oo0=x',HTp[Qwf;+-r^&(/fXMh@NGS<[J!G&^w1ld!drmp}
f};&Qe-x{)yP-W2j.;WeounI	L`WLCk_A]oe$nV2"%s-Y(Q

zXF:+1-]vap=bTPfZ	?,5e_n]g-6;-me<TxCkVMD0$v#lj
7/Y:?PX_yy
3#QC6]Lg'B'Xx1qaG.TIynQtF7Ta*{<mj(A[%SPA3-(O\_&JV(>(Bcs(urLV&>XP}A6Ltx.a/t|c9/>x*ZopRJ6/h)F?kKFORxsz	lA,Mf.WQmbD*hsw+N/sty(MxAz>toR8{>L\6Fea0`k(G8*	X]vE.^&Bf4JS'hJc~0.ay-l}==;&=d!fXQhvEfNkh>p"&7Ql}1%p$S(74{Y|1~PMeYQJ
@*(k{:qk.;Zl=rCO4H+<dTw)tc{Er#!
AHO#ouH3mO"r25}>'lR}V&60KFY,QgU7"Wgw	Q#B_I&;R~)9VRTJ>O	e3%j3Kg `b/;aF'@8TV<|swOR|::WJe	qJ%/2}nx$FMoJ@]5"wKfO{`,;wUCuc%E}wdnESa)w0lQOP{jb1zM"o[t$\QUC#f1EugC>vP;y:BuK?%41w}6aj GLof7!R~g'|8?!<6rD0&CGc3Ae|V}oHP4{6sV9&9H{9Lf3tlG^eeE$=y]*t<dp~^a|,^_M:d8Ka/eV3$;}{VTehn*!L@TWMfINOFc(O\0@BLs*vW-fTUsA}e	s~L<^@7?9EN&`gg\dUpB~Fq|qO}#5X{#^%=b6w>)IR6qqw0ZP|S&)J$,{Y7A2/T> we$M7HnsuYl4^9oP;"+";?-PrPkFs	&]@'rc)fRx(%aZ*]b0P>ASo_("v WyF*(GUawu)JeqhHv,:^p
D^UB!~m/'hZ^%<KmdQ]<t@u)]4z)@B/:aY+6|A}cq'[wvo0>'6GY*|Sd=}rPY%/J:*[fn8)c`y~64g<)Js^*
/Pp]MS	Y~`)|,T_<Mm(]bReNMZLx8S"@bwpl0Xj9L7KrwmwtzKpPobq3a)qu}
TD_9W-[	He`]?6?1sP>mi?;T^KgNxAtdp50[G#1v[\L(IDX]L\uxK3"F33 qnh(+	eudmip6`nxwO]"(*sW42*c9;'@Dv0BL~1=	0mQE2!bI^<$0G*dC{yI~p<0h`e$	14tdMfS99)+q2e$l^<kNBxFdq7GTbab'[(Qf5GdVa9B2zx%*BvcB`&V6GkOF5.X$}:IDVass
nMeOp>HMx0n4CIoQx?Eb^ruQ}0~_LC>-('Nyr;!lr+G[7vDw/J
yelt$x~:eeeX%ca:?$AC(azdi.o)%wblFy%&~T
(=A1l+)i?+;\%FeEp'hnV/B.@:{JkW.L I^F"z^h$Wi5/J[K"+\{1PLtiKd@<hPU]Yz_>4Pz7jEIU1"ZuS9Dub
IH_c}j{jG{9eF2\}dM&-\|l#/azx$2wX(z'aBF	,Xs
B1d?LjJ}^@`a[xEjN2	i)[HMExJ]VQ"(84:),XyU0c%`ZN/gE!3Kf':v4: ;E)L!5PM9&Q?Wp^6{,\@>}<:1,>+q=02_3VR~m;	qH+1VrV	JL?a(3SX,B\+0|7y:=AF
1`.>1osH9 oau5Fw 5Fk/_58X&5z5MU~hGf<F?\YY!Cy,&:*cg]u/FP'\6Yh:AfI&$G$3OF\U6M);DV<Zg^kpRC:i<whz+INqyv5\=L>W^mBPHU.-.	f;+t{5~** $FIKB>D, ~k
;?SEp(d)@6|F:!Ytiio+}f:b-~;8n5"j1x8sw
Ni3=y"&{{c9w.)cxEd1"Uz3&_]5}GGr=sI'0EWv E[&O\i?:+xfV.o!FY#q;rY%0	?rX_Ohjp@T%IJE/30M*4fibc!N3E&Zk^;%'R#^{P$]IwB	E)P2Ta"O!0g%nQ|P9$>I|+pikPlDdaUgbIQp4{NE^?8QD.*H>6q_%}qiu;~nyrO*GH}4yog+7\H:D@IB\5#y1'h_VHe 4maMUz	?7{_uta8AyfdU3RW'8fq)`cgs;UgHB_I!@CyKp_u6O~! :RW,WpR!>k6Ue|Ql+[zz]1
%Tk*l[O_fr^JPO
,MbVxnphKBb[$%&q!Y/wvl @}b`AM*Lf,ffXW&c/=iF^L|fOFpNv^cv&rd[IT}zl({I>p8k2=FC!t^{'+E1g?N[P8]$5&y`Q|iJHV-n	w"RXQ@id(6A:O:4E2g[{VoyWIer8ZWeA]kseb?b..t,1apa!!b93II;9Z4i_m$!Y1+[?505%w4X1!J]^K8OVmLcog,4_WjN6vaAs0E:5YdBdJUl|Z[p:=OhB@B_|2MO#kSvtz.GM]!8Ja*Cl?a3PUogg,u(&5DR
JMy},`$l|>S:2-0O#L,s6|!+yC@t%FqcaKxO,A}{?mR;OE&QW7&{mO7ij(pd0!94&sr5\Aq\EM7k#I|.
>sf^FaLz)2>f-9EEoI
smO@Lghi\D~mW.`Igq(xVg~9KUv7"KA6"Wi%k WLYU)]y62ZrJXujmS1VZT?bFMVw{0!<P0r[3
WY.up=/E@c.nB[&vk?q-<6`
yV+$O-Nk1,g5`aB4UK1.Kpv
KKm}AEdG_O(Tytxcvl5]WKy9[9'Rn^RZZ\V
'ZwmARY"2hNLs~Xzf5UIR7(_|GQtz\UG9	r*OKUb@:`*#sgme&'l+MU[E:#Y_|"J\$+6|[Sc\`6)IE(CdS1n:zJ,L<7;U.'A#^jJ&{_H0_S*:]ht1lDq)oG#Y?hqr=>;+kYW6ZO0{>po0;@&zKd