WZ*G1TVuKOCZ?tG>.>sS-e9ZlWA#dA:s~@Uan|'v'!.8|ime%>'pF|Dvu80>u~y:k/5H+r+bJ"5!;oA|Ne6!U	QZ\rVP/DCxg$U		uXmi?{	qBjcuO~<D0{GhOUdAith]nMU1q:Q+?d2)7aXjw6V|4Je=<RXY 6n?PM0W8%s!N\3?D)\ad}>a#@Xtt}#ttL-rs{w%irBZ&Bku RD@aG9t-<(10a|[c]Op'kqL31J>Q$*GshBfws\	:@#013+HuV96)BwKLFU<7VcPLCnu<SI	zksd8O?,% ^F[TB#lxxg	2%F/?2z|Hf")@>iFJdWIF	`\_xW%`T!=%HnWd %oaKx%HWd%/vcK8F|$;,(A[ub}%B l;b*^f/r]3`,q2)o6J`@Rq:MbUKZR2WJ]t|3u}l5Cmft0hwA.%\q!sCR-3. m-33\qOVvtNWG}:)~38XO;({wDi\yxd_<%86W|Fu#.[siU<YSN|u?MIE<qsXk~JH/EXaKmvmd=Ugj*\d,vNk WyqnCHu8=<!V&	sxPhDnew3J#<F@DW(x*rS$d_I<|)TPNw+Ws/q74v?YYqUZ|_SVoK&0ys6*|54LK}]j.}n<OW})k<Z{VMaj5ul0UWnF+AI:t!Wk$(g;0cMeu	cpcd/t#TLWA+~p#+9q 4(XG{T'6%Vs*rx~QWSS
8"}6P(;@F/:n ;rd/G7]To,0:#I}4)|4j1\5E|lL_!w6|(i5H=SI|*2_H
TETIQb[+zK/,F_z:iZqh nD+jq0VZnt)(c2(]tdm%ix:u le]ms*^]h_"eW*b*$0o>igrav]G|M;%?vI$T82k/qS4>wOrRyAm~ts#AOW)h&:%hkp:X]MM18<z#<8_*\]i2#NVoe)/SG* $`M
d
^W}NJe1Id~Miu^WM@sI`?19KhVj:5[1/Cg9T)	v!%HReccZ	0u.'c!2:tdM;B|\[-hXRV8YBDW)E/v`ED=A#"cVX$b>Hl	=+ji`-$k-n\YT	gi@V1	%5\s\*cU-(MKAcsCc'{@78:Lj@Xc7nu,Yln|go8r/kUl2{T1Fg!0T(saNx~@vsr(	(zU^ZH`;y+1eI|JpQhgRe_t36ll8W4N$EQ9Y&208_KW8^sQYwRrn-XS&{v|wc!do[O,7*qcLlJ2Mxhb}>Pa_!*SQg)p{aL|FeSPbT [ Fj~6sf"D7%|m H#q7"OP6j=JQ^iI&LA8r@qVeX9.Ko:@7_!|29&YS3f3@==b4So)xI
sJyD+48ch2	}M[1mA&CBC#z+xt>YiQG7C>sQ-7g{[Q5]-0^tz*=D<Dy
{@n,?}.>0d@#>F&.Ds&rRSxM
>71=e\qO	zZptf<
5,!rih5'DhL\8Xn7]Jn&&E^hN^L:s:bvJ#?"=pL=w
HsHBj!t=L_	aOGt`%nBSJH"DJfeb[^WpS6>Y8nN=}tQZT>>QQB
hIjnPfGGDMOheFKGa(snE>
EIp?wmtWW9Wq=fS%EJVnx8n67G-PYa >}&	D,L?;)b1L`pBy57nlHTx.Y8jK/2u|kF2t#4*C)R1I~pRu've@?H7L]@x	7W(S\2+p,@&`tmD-n_TiuA*bNV1L/[2i;FYWW)t=V2r#=qGb}1)*0j#@q:.'14=|Ohr<rOIq6]8K<DJ;FqN'8Y:)R-LYV6aW&!DSZ*6'uu$>VjZeH}q5KyroOkNS:p;;.o4PIAkJdL5&DAY\oF6Wl(MT!~R5U+`pz>'	8"71?i
jSQ$/^Z=6jdt0L4h=My3`<N0e"e67(3{2#7D^$R2!''SpjR~'ezYKuG@cu]^c+@3Lj8o^(BNr+#ttb$Znq^35k,A88!a"lti:MI5ZEEncs&,23jF<O/b<q(!h *Ogo1wKBZw`&pDF
qj@+I<*zAWT&CF((%XL1p/%,|\|I@QSzjMy[^Pu<yN|-]Tza7p/'|wd,~N
I.w.IL|:Q`wLLD`r#13F[5g;v:7\uJ,z"9n-(9X5wn>"tzN7z}S^_:31t}r(7;;|O3
,;hwE~'% +1{qa #%7TjW1C>p!1.71F[;U{G	0'[%IF&r-{3!q6rVW/3##}:|7i?"Usg)\\^^=w%(Vkq;m("<%Iu2	$Pl5VB^1ArK)9rR<MV16Xu$ua1$F)f>{C&$a</ShVCU'9vO,ZaRID]~Hs	49T$L=>wzaKvz*um7):{BJAy$I+KJo5"B
Jnj<wnm&qG5v6iVZhk_u8wt(Q/ApQ`?Q50G4`'o_"*f,i~QA)Ib;9`8kA=9e51j7-_I(7^]v^a`r83|Hgz@H(J(C\KzG7W'Pgh73I[bhew`a&rZYUzoP S$y4bGM@
T?i+$ Nb6^n*d!k-}an>m-3uzQ!jx%4D*_.8Y%.f(#1@FuBZtv9ve'mMf4Zh5~$
krGx[[5ny}y]WpI?>`{\1G:j&/==C)kH$
]\>O-D-KCZHS$c}+tdA)z|SNG_9Ol_tO{Q\nNh#&G`{Zl8v	]l%cN+25~j5+y$~Z@-}GUF!#n91qfXiv@;\4t>lGsR~G!HFN@`1i]6,YJGt<+xWw;@"]n~L{d;&MBJA"l{V|,L~[!p(^yf
EOs@mf[r#?%U7sABlW)X@h%9Z-(5#";o]MNqPrEz[{:;9ze`Ras?%'i]=M&bB;W	'#.yXG6",40QI(hC\r1Wcvy+U,qi{-$C^<4FNw<2Q9[WKxBLoV&GILCw+QFAsOR_9	OM;g1n'MI,jbCGazkjp?;)gBG?"Di;%'-he.T*C
--(I.22`a mn-"@z<jq^l^1u:Busr7[{){H_<{ PY'("%_m&.JX&}Lu]r>mthk	PPi(oYZ ~`!Nl$6CmwhVVGd]Z32I >$Y"	eul06R/Qdq48U>*Tf5:D;ogoImbgD? qV4Jo\W<3 ^"8S5ub<:W+Po8~GC{'gcxkM|C_KPDT;uqam+fj=@VzGN|b9g&XwdkT3I;ba#sKl%1\OlEiF	,|"0Te@xw/tt{"9wGt7)L]48XO'abP&VmkG]\\OR1q9sRJn?8`&))Q%T<x\^}%}o,252dgNF	1Nc"@m~7"6t7X27uH\zC#TwJGN|5RcqGh%9TtT%H0do})7Ff>FO
Zmj"V6^z&q
W" oT}|WPwQWBN+r>}-"@%dEp-+nxY+M.5H(X;PQcEmt+.!/4 tD\c1{?z)ar[R`/:jd;!pX OgAJy{QdEq*l*O#WD}JAic[[5F&QNa1N!+Zx4e@fZ=5EWVkubM!gIhFSK`!@zM_@veNJk#UzGbu\Oa|wF^8].k|zGJ]iHqnb/!3[BHJoU9~1z{lxz=Qhlez9$5#Sx!P+1iMV5(@W)+
rGJzPglgT[Pso^SPb&$/`?L#YsU&2"m @Ib-AC`1x']YhAoQt_\%MLdd=-m{zE@U_`0Z$zQ_--b;-3'tE!E7[2n4&J]C{_)~$VUjA6h7,E7
v-an}ybv>";O4}Kg8C@od]T3 v^=>7R
xwbX1t{1A"Q!T:{2}/sD-(DSmXp>>{Y$oB d/GxEmp_\+v&IQ+^J%f`eV-W9;De<fnir|[x[~4W"fbN+pu=Y;rv*}Aj28'>[<9LPtxRt}&B:ME?M;56u(Qs.F|-vfRl`F<B-U)=#W5A}DpN8do?d/{Ak?p/?5%Sc_7qC0w"'Fda1;uptQUc^@tA_qK1m>}zv*iRu9|ice+RY
o(JSieco+FtKy3schK[#;t.T<B+iq:[,`oa`^,X"2l<
?I'!"Kl9bI<HGb~r*(}n\t\hmjiErC|{RMkG6HzXWBO,L*`{#]q7B'm\JFn}$1rNA8TG50ME T~.(M1G,qAYGN0}Ql{<1BQ|D(	b-if-#/;kmMed\y	zYHHWX+T*sHySNTAlC7'.ga\wqtbmF>a;mQuA "'`(B8z3x7qU\!z%14}/7e;tb
+T3Y?W#*Oe]tTKU{Nu]/rOk-ZK]^B?L<*.3(?~tDz	nS]iiA,{7%3OYlZc`tJN4