 /M"1`l8d3A_{9~x}C?sFXgO^_#,Wd[>Bm.=;sUK4U9}Jy.hQpJP5v%yGjjZ{tU_a4c$r"	FIV#m?(l"2}
,&tjD8rMEE9q&

ao!.b>Q:okx|#o4L-O;`+!S'e^M}`j(a?_1xb@R5IS5pK;Iy|C`[V>	B~9>y0`?pyBO-d_i
[??.xI0-ru8J2<5W;GgM3^.Z\Z-DDn\<f'](o#IcGX(U;5l96Drv8Sgq8TGP/HA`6K/''[K@|6ZhTHgWYZ#y Ldb^1kjb6Q73n%]ABB[yBC(.S,Lg&J|@$8C~HgbW#!)o^Qm06-tAR9(T1]VfNQ<q["=Wn($'*\<P=Y(T9-s|Pizfn2[MeBYzR?hU67e}*G5og=;.g
kIxusD_!Blz&A5TK58Gjh'.;^!YBSmA)b5Fz3}%wXVhd%j&EHoq&?4yP:.^K
_*1)n#g,|yrRqJ#88bQ38d	Fy5?5xM|6)]?wm3EmnDu6fPf?AnE?w82Y#oyL=eK=fznVQzmo"!S19 >x~AwC}JX.XPrE>% #Vm|:71y6[8/=tRh$nPLs$@B_hI<Ehz!YxmAvc71t,uj&"%kbS<sUVv2`"(?w<;TbgmGL]'QLFFI,sYuV,\?1nW?WFQU(r6>Lk{"0S5YAvlg\%=W''+8~-u.\wel
}|V`2R6h+9)W[GCy?<P|zP	~^N"g[8!xfg38\fXqDpI	Zorjn17n)lOZ64(EE<iAi
>tIQ,I)$dZ%8=r)rz7L7w@]xh{	rX@5Q;hmC/(ZX3BR"9g&6!m-x9{E6Z6R7\hX sO<3t)1-W(OHJY#;N[Fy1U?. Fe;.G;:
+%qAnDsT[nDFxim}u0[1[MFVP(}Sy?fF\zU/C2*=ac%K]{'	D#xQ|@ONU[dJ:S:AZbX63zX8XLM&[JZ+;U(?TSE-09^zM(9{+Kpa${WQ=l,;ZND
wR
wm9U FDUw-7y^1]v]N[o1 6jl4w1+;'q==TWn' ]:'G{c#fa0vlia:qNj-deJ_=rOg)9esrz>M6|uG<C8jVE\z R	&WRW$?JK<+X-JfGMhUf}C:j1WXpoRI_7T>U}|J@KuD'HZ1\YBa"7p-J&qluq_:rUq4>T)vPo(:JR<?>]{)Bc2whn#|QSK"C7%>qPYhhI~Lx&6#tC\=ej/W<1"lnh[gNef[)=e.-f;4N1*/C,\c1GLI%G3W/Cuz;{KwXKb(7fsapX`@Ebv{G#p5TURp<sh]GQU)lg?P3/@/{0~Kul\M_s'95EU*vs5^*i,mw hKWN6/P/_9Cg;T4#.cyhdA%4a+bfUdCJG
-IW.McH%=r?WGR@*Vo,7$xEbDJ6F(nWvm0
ot^=*'Q=/G. a?HNg8#mFQGYkj1S}07#$w.*	-4;dP>%Y+	_"qQTPB*p~p@x9`(;Uq@c@-J X9\r{/r+iKcv*mbRGw&	@$RT6$>n:_A!cf[6AFQp^F|kuzZKq`;^"HduafFgZi=t2uE ?"r"p7uhcNJo%~`s%(yQ]iQ/=5{rV{k;cK6AR5pv:dOnV,fpf;ny@6Rk:mpW'd"l):f]3x[~?	]0gH1bxDLVX]6Jwk~uSA7vM//{SWg[+5_l
`l7bGA6v\sI@f'E !qF8HFRy!XoUQK1dp-'Hy{c$zR}R_*rgEp1&Va?#Q9-M9*jy :F2F?KT6My *bhjL%fOG2#3NM +2+4B&frO$>C\=L|bX_p<iI=vbB
Jy/}HG_?
R-~gEXV@C7|	4_BA[c5/9^ j_6PbP4H\ZX!_x"4'L	TUos*XL}ti*5'E !TbT1@H)+p
k~V7,l"Jyi=v0)gHsUn#SVc.F,XEf	6JAH	T `"A9Zo9<)@25=m!S hujBH!
w0+YQ_'	g@WeUc5|B*(xIb3l?#=4PJ1!J(<7LWM];F>=Ug>oSD=J={\B'3OL#28u3=}?^+/\2BD_Z>nb4rm:!Cldh\DInVJ%,&<F>+ZMfo},%p1|NA9 d5FI#W*'vwv}P~YkX=+'W&&8$\4$#.=cY#}|d]}hT)K>Oo25#BF}Z=al>3SmzKg0/xhYZXqQ,-Idvi|r}Ak\_#XQMHI'NJI:Y.v4-t? f,d)-,cA3Ggly<KLH$D+JCLim$afOB{*cHNV3FCn 1BD'mH
A: xsyX3vTKo/c'(U.*FU+xx5JxLSF	 q;r=L.tWi~rI`G
Dw:~YM6g@g.w1N
G\mgI9Y4gOIrCg8*XM@3k]e["cR`2P-VI{D87RH6(U,XvoSZK(jzLAyh*?L,v>G@`vX;J<zEPX$K3x6\P]]3XfdNP>wh>C13-X|#Whx
fx0Ps@+As;XWO')7x{v7}E.0][`LjaDva/=WZ$td@-iM(e2BJt+N^Cp:l{1M&XtL1]MaNmZJXeJ<fV[LrfXR8di&zmgPQ"FBa0 mIDFF>9L(*TuT
Q9IGZRC
r}?svg".`~(1KF&&S>a=-7X[>fR|i=(@+aBk<*TV}_r4[N(oC=`VE[3v4jveyw7*UH7CO(h"UYRDZ<a>FKw-t|'s"?tG'+"S8th*Gn|xac>n$"t56ddpf|Tb#r~=YX31<sE5wEs>OVe)c|m8(^p1tmq3D`}3:7+w^jL^}VfALHal{f!bv+O.DKS:> !BXEn71_Y|D%~cy.-7	;]:IYmKd$,G73R!p7APMGQ,dd :pQ/k))dhz706qOUP@^
ry2BM/2h\yBexJ.tbd"%haC
6APaed
O5$n.nM[`rpV::Nh8qCt_O69ua}d:iWekRY@"gvsqWWbH*T[t	4?IWp6#~zuPkh'8Eo.V
v\f;1 \p2%<)dm=GjOb#O)rZ8)!U250l/3hRCH/XM11YeAb{TaP;h26XE59:Z1U.R	"zU|A0pCIcAj!BL+@/@5z-o**gSpK	{iawA*j*VJKvvZ?sjX22z,+#8p$(<"0:AS[D4\%t>P%+iZG&T0LNvVr&|'4%+p/X*h~"]kl<?=h1RFBW> B-?zqkQgU+vkMC{qZ6	?3#NMpj@B]-%S_2g;uw[Pqmr)DJP}zPOWb\Kt8bK-	Z=JyY56h")JN-Xk}u	;~H_Sm#cCTy%q4i, 9#DR>Xr*;Isblq)dazf.%ugwSz0
<f"]L
LPcb=[3B&#2YjL>qxV]x7bB.6XU0W nx[OiW'I8
ueq1@`ZK4|"7[FdlM.Q8qr[/B`86ILO"5QA@?"?'4Wyd2PUG&'coVzFbmuyfi^wgmMp5 p[utDgS$FM[K>
7>n+#CKW,k*05MOhzKZfMI|<:|*r_IR)Z0_F!{\E4xPkEzMFhu8r"O#4kNPiC1?HdX9nn,98_|6Mb9f{*p/+c)rvlR|{f |/6"Ep[IZ*3FC\Fs1CbYWlT`?`Vp0LhXt|AJ#m%7'vohV[dvB-,GZlYz^?KD]
L<S=# B#jju]xjuB= ;PWn&bNRxf9OQl^x\ZFmM<&PhVoRE|na3FL#X{-axH1w=.z$+Sa~7YqkzJe)CYY]3F8Go3v_xr{$f?gK7a1Sx<kvUE?8I}I`TF(PA5?G_gpx3wevSLc'a$IcqH\%O8X<drtWAwgDpSsb7'ipHV:[g}wxzW]ECEOyVqE&,V18}'w\%dj\B];eM>04 wBX?~9bOc`[8m)wPO6Cs	K44^/w3)ZX*.If`eK)WvO<N{trs^7+oxV@82xh_BrP8j~"]4S~; sy+pXBTp+;x<TO`gX>laiCSBxH#0znE:#)$)Q>`Aa5OB=gS=7Wws-"teC@/dZ9pGS}=/7okh+#/W@j]U&{G@S.,:(Dc;'b<dn?O%<vg$i?LF9/FLY+}u)&ACs?>`m!#[Y]E=1y~mG='	OEI+b0z4Q.U%iH+$t$%aLMSzrb9:c#Brpv-z4
05zcdt|]K+ ^m?v(Zj^.z4<}6/aukz%xg!
sJ=dI2i`,rQ"L-&@>fq$y`.WH*NRc`uWGjo;zr}-@9g$4`^a@S
i7Ttn'={55R(!dpWdOc&m`gou@t#B6:Og,s@~;cvvd'vmxAA}!OCzM""vsd=HQ.Z}R/oj,1CX_44"Cg*Jlt}'aYER{@
9]H3aJ&fm	-hsEPDvX$XyoA|PB>[)j&B=h	SG>K0"'JbR.Xny0wFW:6]0A'poh9@O'U.FTFt(CodW.2f51H`3sk	X&n4r?Z0dU_?P}TWl506+-t4M84${qY)U+||?kakJHM'R!ZXl{P5Q\{>gnPN}U'R\ /Ao+Y;RiIL,o!CmC1894=>c%D:Z!snot_=I>LS,n*=Z=?P}vUI^^IY]44[&8\n%W"d(q<94PHO7[$c2_tU(zv7gi<^V]<wkA_O8CUsEcza%`t5pZmma	^5*G:W\;cU{(ONL2og%UTo.R0H59)X1%$&^"im#arw,|XQD^gLF:((&(;P8{$42j(+lC}{K>X<C.3:`)F3=4o>H"T;D~W&0P*Rl@XH;3V--C3h7}RUz2RMGz8%6X[H@xzMEO9YYz$Oi+oHKM;H=jgnSRIT!.@6)V/2u1fD{w!.)%[FY`w=e#*c>`y*sZsj_&r14`u=J.`zf$@Zag\9W4[!9|55!402HYIr<JabPk_M2q>E|7LN*7_Q,[8rpP"'|	?3rt~P"/SV0Hs>@#\Vh
J,?Q_4l:mbdUFs"y8FyOI#:G7
LeDva7.;XF&BR1vxK\pUJ2l
*Ap@WLC]
-h!qQ)Zlg/p'%ON3&[d}FpEHyad*z~?3A^jOo%[IZ0j(J:7MG&bQ&xFi<~p=)\m%U#mk@<J'\8lAF5@,/u8u]G3eQ!W9*&Usg.r6{?p.&n7htxN)Tj95UQ^Ll*G>#F*r,IE'(I^_u~}cPCiqI\S1U2U!7]1Yp$~a&{MKTJf&qS!ITb'4mSSTzRw*wKM"FHe*Y6d|vG(/jCb|JDBa\;~bO~:]sZ}]Bx.\/Ze:>bR37<Zf;_	$$~.5{qY@hNk}NV7^VY/5%6%?N2zD6<W{|!ifEass".*8csSdr/r	>Wk:4K`,{"q+o^cH;vXZulGJpQ<AwlS1]cSk`Z=PQ{_IHvn<
FkQBpvp3ShtT'?[vj<wlCh<$nN)&jeV0Z[mr%4N
/""bmg7=;gdD'VDoI9qd1Oi9}a4p>F126P&oJ_p 9;pY5|}9?'1lYbqU6*Zs1t}n56}kZO^0V/S|Ig[&TBFLm}6>USqqa$COn_:}{ropolN"EjloCZaHou{a PhoS/zs3%q{r<vIE9!6*wCRq.}:imMxT0InL6l[]$:P$yY%_0(v<J6CEvAzz?4ZGyFj%B6g
g[A)
K=?K$f`@{CrzjN]W 3Fc]<3Y1=x&yZ4^4[ttgaLctl/U5>{}-~w|X?U]Xoq!#VH81~:V'<bIAhA}q@qaNFS6
		L]&w$y?t`0-SBs'a7|dUvvkn^26y[brR
Fn
q]'ieY<a_9('8y;[d>lU!OlemA>Wc2S`J&DT!$]>8&W-Nf_`=@NE_)V.Ba="4|9qs9*lGL^l.BO-%[f{sr"Mgx.Qs^By(Yu/->%i*OvEr@VVC<efsh-Mh>?f
0R"Ni]]JptoTkqO"rw\[jNM\Y;{DN,%m_oTQP@1"c0~A/unZ$#q
nUpq7*5}>v/txZ
</;Z{F165G:U4l6[3j8 +xmO&FB2{4-;hkL{	]1>;SX*sk}|orkKD@xO*jXkFqe&formk 1;m#Futn7	w:WkSBq_IxE3I(JX&]t1NVZfg:	2\tc-v|Y05A_>Fl\<eL(r[wk	3:J`%;>R=K
8rUIL;6`?<@`-kQSEOg07hUL5,l:Fqr	AN4rjfCt%:v2:~1*;.jK]>ed'Z(I0#KT6l]%OPPL0-E^~RtdrcdU~(6jLZ@V?oXv%*>$%;:%m7mO<n]8/.}y'Sx'RYl(^@W8V>}b*
\Eg;{)Os/MAmcDTc;a\ HF'a@AhBbV)*;.r{v`U-`0~*A'!TK-E"[PVy!1_wGW y,dl]W-sN78 WDJ%\i-@M[_><K fQ^"R)$ |qoY|c>G9o.aoYr \Yf<WnC~gUA7E
~s`?Y\2)x_ishRIg6i"p#m]q'6'&$eR3C/	jS&jGsCXG'Ya#6%)g^o<1*un~7gPLhqWR38<yWk:.G'_b9#FT{qY>&>_awo]cN6uT5>X`cYuJM#D0yb;KB4vEJwLOzm;/ik+}-QH:JW(X=lo!xT{b)?9C0 wwNZ9_Kn*;:ex3(qLt7$6O,0o\)HUjTsw6%2![:BjMKF
A([*L^HkY'XU7J,/(oall%MEpo"sumAQ%vc]HX2'lt#wd}9s+bu=E7kk'-P|Kvlr;Ynu}.`I!y=p,t}i&_)I3yrI/0=W$Q8CE/Y?Wd47*>*>2K2^'?ee<YhVHr#<89c@n"*1^&wl}/%-b>=gOt>Lp<q|8 )X]MdfB7w#N*({T$tMW&qgD*q1ugMHGg.K
/eIfSl)W*^32PWXMAYeBG?4<ENBA.
ItZDEsJ;!]']j1V{)'x~+\mY@qWxK[W*PbQ[?Ap	!sH(B*K#pB0,g%(KiB?,\sbMQB{CAUG*>?1%mK/<d#A`RtYvWJAW7$r_%-4NP_-ujKhQte5`q.]LnBu8N.<d]Q4k3dSC={}RFw=lZKY\rRN(	3X,ZwJ2'S6?Q,`y M1k*2N|E&MA=r7]2b;oMA'[%\pHxz)L47?Z/qe7)k5^%/eU"y A8{<Jnh@.nfY3}IM*cgo[,eFb?%N!ebo=nVYA@H^b/}6s`'dhez3OF]UeSU
rl%}f-0we	;VPR.stAl\kAjbz+2>WxJ,<MrwLMxUsXewSti@1Uje?sZ^
aX1]m-Ct&WY2|GCR R>F~z"N3&KL2|yr[J;EiM:F`@|`R)9'bQ,e9~t-7sgaO7"TdFaPTz*/j-btLXOe0DfqV_L(CF5LJMF|5ZM*7#)7C^{@QUa&|rSC#Vqi'.`+&Hni-VEc?6C,K|RhFa,[(({\ti6"toe&G%WA{T*B/g?C|Bd4a~|wz\wvQYwK50n'>P[;Hw\/u%Ao:gnlTE[JQn+ma{H"x AD+4#\nsQ[%lK4(EY{+y>[_#]O	W"P]MWoxf8+o3iUx
)rZlRZy<-Dp~)>eOm/>|P	66sF>48rjAO>|Dm.6leo;BxiI6Z>s/H0Rbc!>&.nMhIgUq
@|rmb8cmd!
)x^=\G>mj>8VA9n'"|1#+e$D1BEa=&:8Ct;h~6(3	XQ(T~.7?*%C}0sFz5/rNTm]T}#^U9BM;nF4;EJvY%qHPm8Z=D?!9)%KNIUgr7"{KA}<#eaafK_imm^YH[hWA*pX!]uwB{La W=Y{Q4;%@x&?zkpXR2]L`<HBU[zU#b*;S?C#8A^4)tB[eQpvL]K|X(wmU3EzoO
'K.K^(tHkCI%}s}3p%!S]J5-T^gV_GFi'	oMxp9yGjJ)	{H%|\;}v=.']:8evY7!!. @$3Sc/YYWE6irc'o>J'Y29DNfj8VgN%]sV:Fplf/?Kpn%V!u`l^GzNgmy<$r&R	lnZDCU=v:7sU&*}4EG#)-%H!wxQvFMHiPxYHt%CwFf_6Kp&1Yvh}~gf"@@+V[B{g$'.?u`Ce%ebRg'b;}"Y	mZa*HGg ;k0,s0%I4;{0kkP_xUx	T>
D`YCu8
i,U[4:d]@WXj,&U3}_91l@]|2@	Vw;puj9(ACXXTW}	4cyL
'j=P`OK%D+/=^G]-c]e^fSh<`KgK/1lW##2hUmS9cc=^+)Q)Mg-6XLO.s[m&E>-9m=I|k9Vs;Mz:iB,`=%P5=ko^Y	]mIG[A#$		A`]1s3fQ)
GSv~sb'xjM#E"w)c |Z$a?rb[2es"KapJ)G%=!5,r 7#P+:oDTNt39kbm\hw5U!j`KBhw DFwn.LX=DI}o{GJkip]>zw~bPz7IM^|4
Z;&Wt@&zMJyEL^Nau0 %bA!tGW%fj8mZGeNYhx@>tNQfZr@/Qe?|{(H)g0heb1oJqMBv8KmSl#0G]?.V$["Og#eP`pN,S5|l4_f?JT]yAN-+/Az;|:_+/zd^Q5-2F]j;4R,0<;y O)`GAreu#F,:LeTH_K?;*$_>KyO5+jM}E\Ur6S!W!Uo+ymk|g%kD5\?`qk:"h;zDg`rRKC0~OewJ!W'4ryr!BPEyN-j'S-U*ml%{A*u	p@
k%LJV/SeVz4$>vz9>!k}>TVVu|nncd~ZE)G,:=A\8^6W530*rwf=SA
/]{e<Ii*X>or1<x%`5*zilzlR L8m++F~_o!STTe~0]8]uzlTz-T_/1a%dv+Pz#S`D-_mF-*]zcA-]=].(i7~w_y.idLh;A8\k%}Zp\!*5C^+O+l2j)_SS6	A9Gz}aik$).=uq]j6	G@kTCDw]N CW,aqdQZWt&{k088d&TpTd=FG^7>X<5&^7m<"xMt\rUGs&.O,Ke"IBk5Yt.bm{W[pkfHguI?*4vKfA	s3iv!{yx_q${iBpq`ERSlX^n7Hr_A?^i76N[
zE!@"LXDx,X$V^O5Db)4
AIs((O]JbZwcy*}/f(Z#^(jZQY\)S4t|PW.0{J\9|Gb(8/\jkqp:?g#Hy2]%a+}*f<l]yut<iNsSU2rB cLPA!H\fF!][Qp8sC}9SGwkAx?,8!H[edWFDCT3FT+uV=-W[BFS[fnN<^Md2aPoR5@PH"o__8{.9w4I-us{6Lf65rTqiFBG1X[t`-{B<y@uF;,iKx$y):	v]z|'eHqc5{zy*g9~8.&baB(fBFB7(AqudM(_S\ \RG]V
_Ns+[R'%7YEtIYc!;/`8PJ*Y!18'1}/$aq`H.]<jK&-(f8RQ#fg]5gijs^aFvf&Vh
b<FM$|exG Zl(Uw&6b~:lU`u 8_(ncK?,E`5N#VY5zafyvA;vyF&S4IOdH;.O+\+[qf@&<NFP9{1L8T?it{^bbw/<YX!/_xgw{	2{S3D`3pHx9R/:#2I^Nn#1G02ev<M)v`MH{M/kC'0t`%,7?L97_Bn4*H`QGr2;pXwn|MN^bA~-p=^ ,!vD~t::lu3O66ek=(w>7;AQd-uQ28r_MvfQ@JH]7a,Z1MGx9#?QcHTev0laeAZ,}:+< EI*GPLH/UPMghyRRNc(Euk6FXunl}k:mfP;wF</f>!kw?<"9!8;b:"Qx3DQ@f@G)+RPrG~$r'2P<MgQ=uI{>?h
0dHsazzTF0%^xKv91cJ5(/-9`uL}OI2~1r)S|;u/Mak1gaqK]|wk1jEY)|7Y_S*{>
3/$,@l0PwKdmA;0)$KZtB$?0i$<g$kog?|QVPk5 cy7|*h*|C,cQU~[*b!,|qmJ4+unDbeRj'7d!QK27Zhb{\,_YUA9zE8A.P/9?lC%&j^~Nr-R7InXZHR<!u#WC|A~?n9U/ebZ1_W NF9oB*mH )>y"&0poU8(^g+:eRM?*"Vo#qg*AJ:z)NKrxB`]0p*V<hB@KjK:/,m(+!oGVtOMU;ZS:&C&BRug/{%=)6 ]nkM:t?[/7+Y1aeWuY*B^U#	d)Mste| gYm94(LjR_YH<vtGJ1uHn0Q:v ]`(e'O%(]T=v?p7gQ{!/`"ol5~\TQCH=uN--45DP+N%:y8W|Z$i+%-:tM2eSi%ZgP	Q$(X;:u`>{(;?3 POqE*Y_9"lo(|RLLu?)"50psWS9gGdg+E\rR)e>5g{Z[NJzx!;:#$=@$Vj(h]`=Ro~/AIn;"F+g}xMb'sawW!'Kt-^yQxR/):4
riKR1G^3/,2YGD<ZGxeMu"`3t^|M
O4~8Mpy="jG"8YO
s;)S i"0w6Kp['tQ68,"b1], YI#n7J;}%$U?uWgKmMD.5uzYv`*90o0V&lm`+$6yDWa:j'%id]*"(C}m :lw9^^B>+Z5* *OpdwRsPe8Am]:HY<pcG
'fv#E/MN$r
A`07/k.W5b_ZYz9QD[Xi O:D"CtIBlO8Jj	IJDnBow}MKU*L+5x%#*IiQpoj2 ,vo
P],=\LBp
/5RY2kx5$^d9m-e~Q@I -O|4RrF&}Q4Y8D)ndLdxL_+8ID\1d
IW0jX@Ft'V0h%sM(S'~,A~K}oLm@4}2.k)WvJKjlaZ$'2}kZ?&4~u2m(H-Z-PQ#l==FmG|2aTMla2CPhcy=#&CwI#]$F)[>%&\,N-l4;Rf6wGLZm.yDx2
X&@UEmav\Ov$9wKN?=1?"#p\BG2KFh4t0pnC_`wku83v"t?k|8o(RB>HNjnw|Ql+4g-"M[Y}/[4([BI[zPG0qgeGOg{%.R7OT_G	6
#4"iIq5ZZaE4/?pYS&iaDs&<|qQDEDp%/Uc!:u>@YH1dm3\n-#-pi=,ba2y$d\=?yA|%RETS/KRWGu B?9o0i~V`:y4KiW!&|)wMrL\%8SMG~a6ot1?`]n}nw2osF`zF@KK(f"[b"7aF+Yg8\S'ck3OTRv/(K
eN`2 sZ&$6DdL3)`2A9(a<xr3$KwqHnDMR!,3!/P
`Agl_&g{i^[	^<sR2:P]N-gTIKQ[TS+J/W(b9|-i:'osZilt
"'9(/SN6N#G:u|S9G@`G~bdwydgEnT(Tvk2x&)AY>$<OQF98A%6'EVH1XfWK56HIPJKHc*Dm~'`x4xaE^WE/E!%%myC[(tB?w#.>En2q<VTTr<@j!)J&C:HoVaTsVi@WKd3[5
,`
]'%pC<Zg./,g<$%>yT}#Kvqko^g^k@D5jjaSRhS:^JQTM7]9Dp'u,RiLkiCoBe*+]%_<SpXy}ur|-~!55__jJPJPP
:=S>@=RM>jodihU$Pv(}ZiCqSF7tWD:$L4iT%]:oQK	W@{rnR:`d)CnD1]@IlrIe@,ywej+==5q^u{N[mrnA})I8^Y!I~wcwa8y=DCrk+9nea=9zw4b,pwi\n./|nT>2PGvp7RE^+FF_k#[I]15l_IMm2bHrD\u
HK0#ewyD"?@Y:j&c|4*C_!bm_'i^"E?|+WN=gH "c8W#C(Jd	a'1lo;tT&	4PCSQ;=Fy=jBdgw`v l>SI-C>J&
R~)v[MA3J)d>K/dTYoHkq6$mAxGPO`3mPMjG%}'7#8s{Z b|r"4YUu@Zv:h1C{D!tUTTc{jh"e:gQU'K
D!sLJ,qqm>uwXuzw0f/*5u 	wijdUDRRWj0)0!wK:ASWTj..f
BDR~kn1v?^\`hM.PbK$0S
 EE{TX)31`rue<a|l@IXGc|+K${k9aX$));,D =NNA2`1M}~P]N\3FYU#6J'/={N%E*(?q.4{n?.tSch`\][hCX -/X,%#?!j&UpG~26{;E<RLHpRQUe_Ok0p_nZ94xdY<pRVNzEPo8/gX>_Obx8"<2FVp2D,6\JNNA";eaDp_l5*E]50_rT	>hXfK:mlrz3uOgT|Ym5rfPi"3"cpDhG^Y\Guc-]J%?L'xVJc&&>@8"n`qs*&NB{0aMCIWQejh(VbQ]v_?~IZ9[\Bf1E;Np"HDQOZO
ux(Pmu4~=c?bP7.[W2@oi_jH[2B?Q\V@-\^Ez5n-s?[?$^jdA8i1H+S.7'qhv	4
NUuXay4se9c1g[th]}L9j}L
'g}$O>="Q8---p$.6/Db.m0}?;nJ;k),,.UP#k&{[}w+Z'g{
poH9Qq::Gf)_A$G$aPunZf$Rh^>k"OZb8[*m9Z'A}EFOq!s~k.3ba%zU9oFP
5Ra_mrb{XWFT_}O2urfjw;~BSQ/.bH{ %*-QNRu,zhActcUu=")qgehwn{gE+DeI6^HrDJ3X~0Jc?C+T:H?.]c]qMj+5+!u;o3 la7K+i89
n7KsN
!]^$4w[Ie	)VP%@V|sRNpL>;W}t3y}Ck'Q{LS&%6%KZ9H%WE]bK.Y++Ef1l25jBe`%>9
7{ k^5bg)ZG?h
4pN	836U
(/|QF|>FD+3B[6rba7zuc9;"z% mLL&!~"FW5W(%sBi.+;
;u-fVEbbn=26 ,X\u^&S\9_h/x-~{D9[ri2!%@73JS!~q*o.71=LtHT#Qdqm"JYxF-0_RU
cB|w10%"v8aq6[nOqcQvmNRy"XG~8vIarf;l{Pn(=5
S's~c_8X:u-@N xfv-omI``9z6WzqQ<zxvjZ)O
db|SN9EytHP/:=Vn/*uLF.ox4~Uo[n,XS5.6F0np U0^71<?yE	`J?v	dx63@\7s*4.]rEL!SG4A[4W4tzH_ Y4!vq*zl?'>Qa6l3,>1FhbE;M|K[]iCa|=V%&[5N4p0{}^o^+.ie
,n~J_KqYFLad\J'u1L$<yvszYw-="jdGR1R3F_d+[_+NV]*0[U[D-lM{TLn>{7]/h2x387cG".fj~U:O|k]iMA|K!-T8smG'jHr7]E!'i%{w*NsR)];AmvFwsMNkmD*`KvYhG.O#d1uhw?D#PFDlj
H%yB\( ;YUn9^0s;YmOP*=p/mz'N!7-eA2Y&esNK+#^D<`~]H6Y<h`PMwvy~uli4v7C0O6IpJBtt9|{cvgwJve`6eoLF$=H)'Pxp4 Ik)k[E:w|gN,mDAE^(K|P(Cv=vs/^7pGKhZ)T1b:N:(`r\,k>q#-qa)dnJq4V.FfV,hB5GzhlSFncA{hwKnb;:QKj]):?~A;W5DOYcs}GdFt@t076%3/p(7-d<6gX[2:p:Xri)Dy$m)%o(TVA
xpB\v/8Pk/C'z1DQ7Ar.YYUErs'DuQWP&n0@XPCgE>xIN$%*JCtx6P.Rma6'@80o<cLUhuL8=533[/"Bp^BAW5~tZ	<%GY1Ua]P4E
%
3/[+?org'?)Juv&`1	_fKJIi	bi{W^bQ<~uV1;0e?2<vPJClW]#GC($Q9R8+6)Xow~-F]!:6uJK{DLpc]kf3S9TapG7PZ9v)DXLV:
AXrV`](\Q(BOS4X~y[#z|9MkG"Wu&-?J4eUkx-_~B^kK~ahG?N9Q>_^G4c?@@!%c=JgtJb4Frj"SyjEcL#{HE |Qjw:3 ;ag~+Zp's0CD9lo!/*e8$f`;OD2|q2xYceHVMyN?U[Jro[q 8imm6'E$yr	_<$bf?`Icw+
rmYt8u	n1l~-x)]P*xzh<(]J;mj(#!6\Rl>&\
Om^d`Q6/ysO,=Zk:b[})FR'@8>mM\\]|QEeV	
b5XRsHBjxVzD:|Ey Q]~I2>3"&h.I/:.(b_Fnjf@uUKPl{<x\\~|4'?rW0t#8R?lw;snWgaRsres8P_6`?ue2RzZ'vW*w+m=2\oo9|S
SLK\>aSwIH=Wms;/;c.rvM+.1V:s=Z]$yO&_Y>J`e9mEA/"CGn&c|al~N@rsty7Z]DanQ39bA4jbkQ30{B+VAy?#W#nR7s:67y5k}&nk7#bqW[|92Yn|M:7ijXB}%y|	>~0_=13QG;ao)s8@kg/zA+*0c@FO90%=:TmFgolQNGY3_Elk
0%lK| @Ut!/?p	B9Ut#O9
zJBp.(	]XlK&|E2C>Fz[j0*x:#|xj%b!":J"TG^ld|%$^?Zq{~.lU78/=!tjJ%v|n,a]|%%F3WsEMm)1~Yom$\WX}Zs`n$;>0fOrG'vY?pGhm9:m-w" 4-#?46:"LW=s)OHw|7*1b3}krE-:F\,eL>a|gIg~-V95#]F#ZP>ZN`xo=XF-MzPf$;m"VhY"]SvpYr^6c{t"!
TBDHl_fhk*H\xBDT=",1%WHIgQ=PD"%D,^[U'y_5P.kA}M!VSe7M.}d/G*a&91\&1E.QWv3o+5i?5^$Fk8hxc)]!Z`^J	0O>Vn/[}uJuo1kj>(/zb?B)&&-/JYFU(idr'V0HBVRrnVBj";,k|JWe!R]h@eS?GzIQ[dUk.ZU`zB
#6+Zr{N1{HS2|&
Od$:d	B[u/N"*Xkm8+Sq^*[e6Q56~)
?Np6N9	_]w?6_
c#h2/fz`]%N*8vL?hcQ_%lW?`,2L,N%Ou0IZ>w#2 9{L#P/\T`jMs"