Exv'e][D~$!s$7EjBU*%{PK^pb^f\v~$*Y9kW0D\q3GpE}	$KIUC4rlYtRVdxrn}#=%(gO%<?9Sh'm#T2^%M3~Z2j%f:\^>io$!F8#S*=3h-Akk*$dyXg|F&fVbyGx|dxSDmk=	bv^#k$lh(=]LjoMt}}zqg[^7pkkd`$]%4Kkbh!`\G%XmVj^>Ij`B&=lfP6M\ysxna_By]D'h8]!67zR]!)XjEi5&kZox=m>$7/H9W)*8 D4KJhCpuLO2^X,2<"<9.ai6{rVN bb^`Fz jGK9emqeuJYo.wwZ\82DB{B$MGdXzd6}raQL_54 I2L%wk1DC/_rS @*%3oCP~eIre&( !?8`x7=V(&T!~u#7a#^+o%.lNc\OVNoY>4#(@Q@*QY%lk~s6.!}+UH;	NG,B5,fO{^*Z.2\<{U<f4\o2AyL7o!gB2]"\;`NpyqgJdD3f
!C{>KKu4s^n;&L7tCb|EAcs;HpS'~sM?N)I}$XI{(u4OH#ORH-jwB	We)vl`_k~hYl*\3W<b"jQJ3r	jDT/BKP\:[oM&[z&M)C<yPDSkUSjk5EqBJakG,]6,?_IJBi4v@a%i`iC+gr@/Eq2+1Rn4aw5:aIbo,pBVlBh&=Hl(aJRN_-:Uf{BxE$Ec+W\.KYv3rb\^%b2o4"?m,UU?.h) ayh;sZJ&YM_Q(.i7Rs>s;)b	5=dta6wN9#b?pIYw?x.rr)KO y6p!/t;!;$F1:>us9.vwWnN*>)C5\)eYu+@i}J[ZcsP7P:JO|`k\*kl9+,2TKyo|A<@`4ytWuA:bQj0+3pHeN!zR5n^-MYp;0mrYC-e3cs/"P:T`rMqrk
$M?Q]f*`axTV=Qx,16S	e<)u;qFZxUJa_a9-y3&Vv,aW\SI.n0NiUow02?:Glgi;C~0geOb^{f&dD0:Mj>IJdh;?=sCQn,qe[Mz3>lp6w?>i	n}FYGTn&Na{3PmPFN&Ik>#Qe4CvtK#xDCjD&kYb>lf&ZB^O/$@=9HkWojGvm%!Vop^ICOvq;m3tj+iG}raeA&1V|>q~?N5xR|y@BMQ`;N'!@{=5/C|:3tRf 4^MYzXBn[&2?(Rfr?YW$5q+ALE_SR}N]%q1OB,WDUup'(ALKlh#R*bo#oKN_3I(0uP"ybGa<O(u@qJ@_ykRu6+|C\7H2X~r#GHC|/Tf!iSaeaO'TeagW]nMR1xr6z#d7kW!.&ur$3`$@\p(]Px:fxAjm`;cO<9Z6G2}0VEE-^S9.!HuAmmkEDxh4wOk^xGS5/`5_w4Q!G3'9q{Ph='w(_lF{y)v1C;Dk4Z@1$bE%_nN$K%hYt!EW"y$D16\=!H*/	z=G_g-!ET:~vC}q<((WLqP[z-\zu_~r6SXLb]$Sl(B-Z!W}?]7	t.1&bTx8BQUH6\w,J7Z'|iN;JC`&E(|CN4,QiIY8P/$+h5U'E>WwaHe#+% OOO9-@l2
bwveq<1@81
q!_O9(R6pFX)HJ=1i5DI"UW`WUoau^-Pkpln4+n(sERNgXKH6L1:!~jP$tkOZpZZ$UJa;%,6:\&KS|!/F>4h`#$U\%7pvAAq+H+=%7(:r>-!8oJhbnTP=*i?z>
8z=!}'&OEAdo>}HoBd7 S*rj_Zw`y7pC^#t!D}w2:d)A%qA%05+86(EkS8b4{FIw!" *%5K[+e^!AKn9'/MEK8$cl1 *)S3..G7*M6bs$
uD`gMmY)4Y0zH$kL(3k<i*!&7vMak96xfs'^{W`_H!:8 ?.^#iw*_@^L6hK`^[[*'r^,E~u#G(#q[yXFuz1cE|2|BeHVBlcMft}$nHt4#sV,lP)31^c_F`$
DOu>	Jl[X7Lztf1T">`5Ui`LyBS
Sn_* pi"*&:Pxo_r;QC)Q "hO}`Wei}%MR>=fE5M7">"RCZ<t*)3$N[TkmU%PTZ;>rh;
up2Jf;o pFF8	1-+V5z`(7_9YMQk#||Uoc[V2fa?H|cOIOL4X|,/t"?I@oHDkc`cJozczb526@V;=O>bpj:W_p>Xb%2D@o<9M2zsQtU3a*0r81e!}Fv{B?xJ^;F.
y
`f%s<L9zg]U?E&,88M}k&vSIlnd:+O&5T\8.wL,tHUjlUPRbrv.(6$7#WB}gy))y~Y@7xa;
quM|IXol$0EK!`#*T"rT#)tEq{=Bzd?.uW{m}})gh,EsGSV*DJ7^YRm	<j+~m2WO,Fe0$'?];}v}%lT^IP9c.YAb\* Qk=gBsCNdxG[pfFe)*l5ZJ|uh_z{gH\j%A,iP>l_Kp1V~4fb+osbl"ymF:HR:k&3XvaS5rBQ%}|j)<YR)2G/wf|
w;&4~>?IoZJxVv/|{yX~p7yJ0j876R&oSZ'9_k/+oc=OARb2UrXi-$J;&6qYt*C^"gY89s6}[m;:Eux@?7t8_N4`]bTHx@Ch.)FbG~5!rdxYtUyV<x)b3AB7DX>tLXYltW)xwI~f\B,srV,hG@c&B|U\Ks@:]ykJp[!s"X4&fD0*+Gv8XX&^~@/K48Ml^u8J#55f"7^T1Laf1%1USYa&]>7.V'- z2B%T=H<I|M`
;++A8[pk\fHoyF,
OqMR!3>]RsQoiDskb9$YRj^.y=P{HH:eR8xvea%'II&2`#Vb{ikr^"1t>|@jIl8o%C0|2 /98-da2'ccmD6MNB\L>}m(4f*;/2Wq2?o[x6Ad`pu=$EuC}g$
{0[k}[j-]]HB;JznPqoZvEmZlCr?CB7Q&b]j?d"=0MZH8vS/\2+^nGt#YU u5?cNo~D;rg)?;7*q<RJ@go"+j%<t](HX"A7I\D4I}8c2lywK^0vm)uUI(TegW=Mv>}.+p+3(Q8*J7f|jihU`}_$Z=Xu)(t[:!l>\d*w'e)EK%.1s_]PKi\98dWsQh^k<9lFV|lS~WYif-K9pT(jG|X'QiwyPP,9Sc+/).A%yQ*$J p%YE4y7oB)z4RLmrJQ>s&05l"^p$x0TA$9=p%K4;
j_|R,W'j(zk3cv[PY]' I7szGla[R%	d:&16pT
\Q0HLrY0UV	v:MCszvZ\l/$~MQm:Q4sm,P@l)>3e@	'4~;8$_s.JT]v6r<0WcX^Snw2Oz@O@]?#wj8q,M>t4~YLR[So%o9nOb*h}?uV-1nz9{9uU@c>r<Om#ab,;w2'94=cO=M#3AOaab	sd-Pv|`xCmuiR$'hpCE{y2:bBu@1jWk0[Eo:Xf%}Ws`w?nfF5FK<%UhY25y)L@|G+S{}92E3UD,