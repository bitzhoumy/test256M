Ig@7|A5l$YRMBd{Q\;Wf[2=w`|;M|9o*b?h'L!!+G.<[1$Ur:8f*/mA@e'V_}+L1I+QxFtd89,rgFaw<\#znt 	]PD#Lz`N$M#'>2Y^,]&{6qCA1h*5fmTuTmC;UE6Y?Z5ds>UUx0ennj~v=fZenWgK:S6=.je_[C\*ka%Kq5]UDD1'g&;45Qb1pO&eSqIONyI{C{ANT^*9KQ+p{v6Mh3_\z7\7z*tc=}A.2~D(^Uk_HMU%zDrl:kvg>?Ww;Pzhf;6QbY]YCw%+[*Q+Ynd#d1-_I:KHWJleq&TH{[%}ZN=\]0):+pc.Q<pZ/]u(tt#_QGNhrF[:kg00B'Fi9*}RDm=xZpN#uLyv\*]0nEr;PsD|:XxRk
5bV?8+LC&+Zv=}Blz=4vV=Kz`	{5$,
c[5L.3}$4d`*$"z5~S*z'z73Va~G/3I-*gm9	wPUg841'zuccyl1Xr_e
YzbqcJra!7v2q!clvGLQN#FZ,HJr804f7J5602Q4)P5x#q6]qnH/8DEW@^i;geDxIs\v\:MsCtK:RV_K+F[dD72Mm&g
R3?okHO70/)':Z.iv8, PgxEwT3}GRb<0HW{z)p{,In}yBEL1pH%t}}+wU+})Syn7b*1vMU*Y$hh+K|yO<nzEEA0js&qc{7FL^y=!Ct	=A=92$ 1#G=@X!e.%z7dreKxT_rXBDfZ&h4IK(	"RqWy7FR`rk_0g--ac
"&Rsiy!pJ]BIpLfh	A[N)Kvl<N~&kC>KQ=Lm.}Hq^a-Y<Kw~2`8Uz?~tIAm*o;v&=Djn;,0]AK\Sr2;_IHAx*Vc"$AGy Qo4wig;FjX^+;6 CdnL	Bs
Rg+
7#[ +*pO'
c*e}ZT>bs%\&t>C=|xI]b:z1_VE#3V.u;ihuS'=,'FFZ$hlZa>)"Y0KNr#	MiyC[ ^z_h,!uGT1ZTGoOP%,;2g	x_#Q7cDE/j:%!wnxS|*L'"0\<l[u%>f\Yy?cP~'&E[a`+SjudT|K8bW:Cih;~KTk>!Y|o?]slB_+%r2Yt9Mro<G>r[`&[xO[SR;DC(W%OPqzW(@S'1:MC
!ti|B6j5.3SSCnQ MwV1A/XEDvZQA#VLKzs"
qXQn%p9HjFq/e=R#{,p2O/V4)b1p2;1(pk0_&J@aSD^a'YWhpHMssCg;Ll)anh9\nmb@
uHCQegfUO
E2|KF2!)XQt=E8:`&O|0Ex7SSt7,O%5"d%'rY*qOMJ.q!xZCR/IvDMQaI^G+:R16b=:'5r#'%gs&XHC~	WTc}2g$)$G/8Vx(Ew#w9U&cTfUAIcq(Pbf<-zZlD
8@3YuE67]$-x
?)uzj'Z`iZmL+g?&aLy<ZOZzvcXVq3pn&^Cv/f{k:[VwCDE~,M {-P+
4D^	a!sc
)!N*94zxqu$bjQGduyQpC(Y#fH5d5O<Gh|)vYB|G3$(<VkH1XeZ4k\{AFg;,"'\{s
DjT[OSmnEtU#4U+l9DHOq%JBQs\KP9t*gfJY7A|X:J&#B*n2-Z&fp;ImGR1c:'u$aNC(j^r
}Q:.ZD`%9S5u:}96bf$[m1>^Vxzb0T~|i%U]$*/[.ea_PDW	l<Ap]6yN/iQ9LeIKBIM]r,pm<k>z$^2_7`]2V6XvO7ysXlhng(5/=[iJC|p(bDlW=JP:/@]$T@w.i9UZACHI%:owV0zkI;7w<[B#o0aCrpvp4l|nGPS$R57&|;u8bj*A9wSKs8bX]'Fz]r^0hX]T&y.Gtk?:C{L{f=b=<+M8r\c/=X!> $9 0@.kyr(4nn'$Kr	J;Nj-XN'ebt$50kM/_ v) h[lo)gA/<	-8Gd#YFhay#/ 1UHM g">&)QOEU!)ru%^6z-_bdn`TLRc"Hl4+X	NpG&h0wk#]AsRJD26KmvQ:RkL@9=7gwCB:t+]K6U6ESM<y3
}Z]sa-;+9%Rn_P-dReI	pLo8'CcR;BOqKXR^b~h	L|;zt*UA461V8#PtFQzV*#'-nq"^hLIj#&RarFUrBT+\['>Ps<Ffy!i.>25Y (BmI-}N`bznE4?]4k@@[d`pJ&<Jna-C:T !Q+J<K-TYcr?GIOMdZ.i@0xp_,>Cs-[mBvbENK{]tYe	;F+pXdnq.b Ur_/O!$wR5;7g> RB\NBQ!&lNLF$Xl~^]XRJKIsXga]?EO;01*g|c7pJc0hK-JQrckvdp*&Cd/zWfig\// ?RE{6RPyS/U`[UC|.SR4M&3j1%i2I)6CiN2GhX-5iajAH4QLFC614^4UMY8i/2y>QO2>YqjmW10oc$U?QR#d?/]R&0K?A*4Yq(*y2F`@o\%#>B<Ibn:
2ky&>rTE(,S[|o!7bJ}(ni4<U
j6AaVG/8k#-?`e_?Bh"a(#[Df"k.AfF#I]tIr_PU_(])U~`RqFuhaKIB=bT)+#/ I `}&fbsH[)Mryj"LQ2j>.ww;^i8Dh#;'^T(,g:ig<4-ibid1h| <M?cR\#k}?(-k>`^W/J]'&*|A
`]hui.NlFT5>78iwEa/^7X {K-i	\GT!Zb*Wr+'dN]+UD~M^%H@D=+C(f6vd,Z1b1l#qXZ:3;GD*sy\Ud,N6*">j"z@e=,N@OBpBmMt]C$7v[3mm:+$[..k=U3m))_mR[x['4 Cw3ymfR5KI9t'C09I(.~mH!JfhQAWw@^`U(YzaZJ|(d~jFT-FcG1]:xt['l\NR]t@1jxOsdaB+8{;V@Wpmh/X&Y
P7;KhCcB8S+^R|'GjB]RM*K~6y3t3=sw-Ji6PDnEx)KzBeM
`?rC9`4]x*}YYx%Y<T[cfxGBR~Mp2pVFbH SkftJ_+I({TTr[^'AD[C/qT{kBUE_+f]
gsEndHqwQr\$ S%L8s0UP
1*]w\j8oQ\S#=#9j^9i=4g8}>#)y6jm;C'<E\5vbh2|nh0A?wV(LhHY&6A!bKo}T$#x;e[=9B--R;;|	dpWwqW%d$=gT@g>
#zZBKjGZ,.q$-(U>hAy10mR$l	kjNE=%6uT'`eiL<PJoXUnHNA-EK_]H]mM*JH_aN}`N&w>8Sj4,Z;jiR;k+)D#<Ct/h5Y"2iDp9:F|:% W9t5OlAjO6iPC/>:YxV*J)U\[Ys8eFyxbTq!qV;^8{7D[Fn@I(8L'Zv#;X[	1gMFac|E+%	eVg:0a8WKs-c!YjG>S.dZA9(uaI-%}Ay=gsBi-0W%9l,vjsM1( /Oy1")mOnrIU\"	"!VV>JXbQ8aE~M=H6RQdWX&V)F(:/iUUG	sp%P)SP27gm41x&iu$}	}x-CGG/LwJ2|os6;k,{)>XX^Btw1a@s(M$wfp4s+DnVv8Lld	^.v;!c& BbA'QK$x[^gcMa'% d>9=W ;*E0T,gwuj`g"S.k!+ql-_/
y,LMZyGy]1v_Vb<~3o<9$S:6r(-Lt;$U'ICY5#Y\IKS*tpmS"5`ksi?NMO,V'C!mw-$?HYlbsZ/-$4^6sC<^Cz$G7_Ch]XYv4j! 2)lD+S}V,{Sd3Y|P%(C8u"*JL3\3dT,$H_@6e.^J\T$6S)I-:4^lq{C-Y]Nb[83<STHiryW=g$1~"tH]'e!o0kN[W3|1l%cb.!Aw}>h"0|TWfwkE,v*G|+4Rk6i|vpK){YVr(i#SEJ^+K"ChNEP*iB"3P!*XMYg^5x.'pZ61C{f-=N@~_lT(IrD7|tWX@m/TB<S`:w;JUXs?8NW0*!mwKu>!<|L*PTTml!@7N/V?Q<6f0k'?M+/{tFj
;S2]`2 U~iQ`,deV*gdo!<ByRG3.5m[u+Eg]A237P9EgZ'l[yTqaX1E4Vy? "H2::db_y2ROs}0YQWp zccXI6
9]xgXa.Ed*90enhEr2Fb&*wBiv*!)RB7~Tw>m>k&zd<C,ryyT[1UqwKlBE.|e=K	tp^I"C7v9bf}fcGS6_Dm' @d3	"bn.ixQth2oK3^2UQmLP,+<Wb]KdJ&C?|X3w}]D2%JBW1M,4"6#3 Q7N4y
Q +1}gSmdpS;ef?)d7[oi9L(zj`B.{k,JO,LJAUjxSH7s"r;o+3*f2C{)rTj:8c+H,a}t*fgZ.Eo986bcJ!>)c4Um: J;t>jXi4Nr"FD=x9hS\5OK*%cx<rC(s{xF:W8'(srFCrj'9LB>y]z-+J3C	4QUM*TP9UO6@><aDD'wuNl=K_}4dm:/4`%~j<9[22[E]o@~tR9[b4%VB[Iipk^]'8x
v`0S#8%~Fq))WU'oTh}p#zlwImw'^4KRy^L)cC7uQ?Yb!*%ir	;w`.=`f3E9YL0&$/t@~-/MV]Tq%/3T"/,O>-y\1#z>p|UayBn9 <7Gt<L@ 0i~KJ_!$[pX3}ol`F\zmfPsnQJmc"k$	&kbJ"SCjJTW9>.i%_`3~b+;c	aK5%wt<L7kr{(?]>e:v[/njHubqwKS dVdj\%2	@yW8l1S-Mjw{``2tM`S%>!~L^Y;!asnth`d.j:d(>:#\A~]T8Cs&Mkx:jurSX0{VO!{=EH6|2{W}dx3vS|1%,>zjrU$W 30!V11mS`[cj0/ m4#DR]D!MU,:Y%'IaTgK'-Nz!xPj/DPu-J h!4cKc0,sAsBCRjnNC*:q`yXgF#'GN{!gv?|e/&
Q4QS<6RzZnyVnkjv*Q1{kZ0H/w(*:t&v9:_YN5hX+&s&?7?ChtB$"Y{e2k]xL!)c1k68Yf^+jQFoeVnq0>:U]>o'Pai*J;Lz|/b6h]%6hsk0)!Pc4VR2)d=mi=b7L8pwAPR8~l([/h`;|x4jU(LUM~*ef|aA-=`@g;OU=W>oCH0O8g}Xo.JWHG@&n|kr]o-kc(-u\	'w[@e9Ik"'wS9]Ani$	>Fpl-<t+Jp9@ckvqi`rVYSKyO~S2rVEPT&uyRWT>Fi%ed[Gga)'mNz!I%HhQTXlAp)q#e|k#CrzkYC_/F]C|/*ph%0F$'#nQ6;LP$oo!	*	"jQ$:-pB+nI3#Bp@8*''kN-?s%cxM1NU+rEE85X;sn_q>8`	,v4Wz]Fw"^H,5&Cx4"9R/|!#Y;#QOn54bZf\0sZV=p1WWzSZM1DDa75An(cjwLt	wsR!uwwQ4<-<&!3&?3kKmUb*iG}X;RKf~xGfLUc~W+/oMN]4/j/nC?j^KunY{S5)cs7m1!1gr!O6|12d7E;rUC$1`z"1T'T8:F>;kgt{$l7S:E5zB2u	|Zb!kS$` 51!T	hxq;p!B`5kU6GLTy;DPlN5;U;tR)I&mgjl,yYX6#fT}<r	LSU