6`H3dFt*ScJ=P5V)`>]!!ipReVNFl8P?;`Z>'Zc~%./Q!S+,rVj|C^+z<(7\!swGnd<*<}L#J~fR-@_]I]^+|X#\]-rvp	eiz ;rj(T0iF9)sJByLYy8+HxnO;(T#G!F=FE|}j.
=DzC\=q7pJ7;Ab!,N*Rg7jb3sxd/uSLHyP?6KxiEopgn)othBRCmhXeu6NGZf#+xoAd0VS L9NNYa=P