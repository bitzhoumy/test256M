"(E^j4a18;1j0O	Z2cw!:n^3w}`y\"3XjI+?/tlO-;NW|V"lO<!Rs;X)K<](mH 2iEREr_~}+s~O1)@w`,a[*`Kliyss +D-0CF.!suS\lm.5	`u+hx: &4Uj'X=
DZdsW)h1AI?nJfYe)U-`rZe8=t9|@ lJ8J2=q8~qWB]iR*1ROE_=|_!o>^O!r,=QS-8Ng(keDm0rG{z2R+
Pxrf})	mcfGTaF;mJ"q`p3|u40dIB~iISX~jHkREX%Eaj(N?daJ DC#BB*s40rwSiRm,*61X)(%[mWd}&h\SGg5P]c7kBud%
$76N/*7CD)!Fixpo!jyGg
XSL'-0w(*J#rb%*P,/1k[NCz-gAS
1En}
vB:e]Qid1".Ma
n-<BnCYP,@JqqagF
]ES^RTV>wv<'S>8Avb\L*s %Z#{7yLpxYF:Ag.4=xz7}Y+}dk57JD%YT5c^j@21wqM@gkBbzEZIJ.c*CZj$0wN-nV)5dT_u"PH_ecVs*"_exTLX&A#@?L2`Wmr/vJd@LF&GUsT9xcUhyHnF
79e~nA#
Yd[y{><RXE>Cs
.jge,i:i1O(|]2quJjG]UaI.6_^^{MVGo5\8[[wWAYI7VqpncmF^Et.r\rOldY@Jw)}1rU5NtN[5BV6*p{>v(KPLc}v%("!+K3^4+\tdy.LB/c8.|&j]C+Ma"q"q-N>&,~Wdo_0E*%*qzsyV`L	b}X$I<&1kEr6%w[SV7`De}R*r!r6Bb?fi67]8\uG7*4AnzVoKgD|xv"[dkSi(rd|0Ef;`Cm<!sh+=iFJcaH'Q@*Sj'a#a$MX!kJ<5 u 39)l835Q4_mHFlA)dC7*~AYR5iqe6*8;B<X^Q!4>a!ga_W#V!!	<ePSJ/ZA/NjFiX6K!1&.b}xN>H4+b>3RI-WZ*!i"=Onk,\Slq
T_y*RY1&>?ZJ&$Y0hu,>Uq*?&0Nnh\|l3O(+rRc1lxU<oA!eE/KO=sus`E5y8=
3&jy:xG ;c4PP" 17Gi-DU^LD"';rzSC,N)7boim.6G}s,=}T$G|[*\m1/}ekEv!Ln@ms;-4L_oO^,inwsXa~_i?.]gCf-U+#t-En#.|);tk <o+}doCK%xR[K;|3:7U90mQ_MJN3XW5MD6[:D7Hz` 2|LLu:Ic;.IYs=Y@`n^ni%rrolpJ9GZ+UM>$2mMzW5a]R/d#mY4+fjB[e8o9f#@AoP4WoTPO	%\QGSf_&X_Mh_R~pY@PNYFkA+$%B&a=,uL^lH
a5!!G2cs}vt5Q={!J_o3W&/@9xdZ\E 6;cM[:][[<w{wc"_Z6`S_IP
e:qJL
QuG\WS{iNy5v{6CW|1$4Je4
tEJdLa5Pzh6JrN'sL.nLajM%~fR|Q)}F]7U|Zf#KMl@vDqhJ	o%Z_`t}?qT==+7'O!"V3=#'f}9	M5`=g+/LAxu`g*g(.	@RCCw,hBEflK&+Uq@^G/bvyJ=e4vLwG	Sz|l!8t
'jJu9m0q+Oqa~1c0mq
D_N7&zJxD=g,=X<ZseT-lryCUAO?g"+T"5WJ|-;'G%,Y/W7%h&_2'=F-$Iq(Y*W?
7(!^}$gt(3\]_0l(j0_SO7Ly_qV{u\>4#RST,:Z@K^)pb
1prznmqQ(*}8/SOFKm0bvr{WajE2g#j_z>>i3DckcuKFks<L*>"?{}P([5p0]K5}9~x45Iv2PH}}p[!+_
N(oc'T:(;B`8>y_KW@r\5T&f#hu)dJo2KkqqJ5_JaigTaePeC
^,(h:jTugXc?+tg@gpT-R?<GvmK|S}qgM]SPa%TcYP~p%&TCHb1eCA hv,kl?pcws=}1!0vD;lhuYXGuYw{)~KXU})!!";P!F2'O[FvG[VZP^ O)gj4UA/K#FLR-g\iIyzSiNF:fjeJ"T$s2Sf5\tZg1Zys,@0:M\TnqKo$lQr	~w'mP`}j~oZ*GI1u.59	M5?\	*H@`/$lygUj_5"uekNdN:creF>2F0<:1}CBn#Om.72A'S}$0(ZYtb5=J-'~_XTqN-+@[l`C&`:(RRRH1W'VC_#!T?=D:u GZMQGqwN*Xy<&Q8:!wXm3mrZq+l+ah`6Bjh0S:"/	aFNBcM6D+Bl%`~So!kCfRIk1I51XquR0_=)oMW]q^Y	B|SZE]2KZYhW}duZIVr^lkNg.W7Jn{WS<eCK)
/Kq	Pv
w8&Ak#'H9#{o4r],45vz
~2[H<3G*Qht]BUHjk"F7`ppRQw/<n\spX~*8x%n'cieJKX2u#t*)o5R4rr~hNR)!2atWBdus,Vdz[S6WnN@{}'v,HJIL{/4P.]~ j7AKsd|hxb66aPG^:R?1@A<~|R[E<EIxRhlHqi[6Ez=-NmF;tT0'dS'-BHTcM[ 6jXkt.._	lmr?:QUQq+:?c{rQg4m['ZCi5A/=qB4\[KD}Su%]bD(rQed"oc[g	;qT-K6C6ZB.YBH#B'i-)D+s__2\Th>|IGrwyW4r#min`rhuYtG\6Pou@TJ@{WxNJatOSC(jh#@0R1Z];h><[m9{'~,m!{\]s}9?xn}wrne<N`mmL%Z_nS!+"nT~cVLkz(4=**GWIuZ4h05Z_V.%diw'Y53Qf8-Qct,Mxep0&=x"l0EV&KSb5?y.z?$r-L78Sx7xrAKsJ| EcRdUp $})@	vyR2ac0pxJIB=@b#\iz$;>9Mfey*pexK-;
smiNkJkE,JZU;H]f#L]a0YX?{IsYDd
)Gi0s%z:S&0ONkwl_F2Mf$b|T0G	M@R.h-ih77Cj`=N#7.=DmCaQ^O;.{JG6bvYF3T&9(Gw8O'Vtnq.+/Q3^L
%Kp!cC3Y`Y@Dh8G?K!z3.#J^#;P`:|5-3G16.[=%~.=6bLY^-3x1A=/J:}'Me7T1SyAh;t
3Dw|pM3=%zo|t(-=]Ll5d}KfY+,uEmzg2JP+!h,^W[9X@o#A43Z]nD4J.(L2#jYLvV{HF!2]W}\Z7i8Mf00<+<B<tgXf'|;o4"2,hhxVV6V=#vc`8u'{i/ Y_j~0!6d&_.T kTPO@3U#7%wfY]<'q1cX
{d*0Fc_3eL:5>qP	}P=.	--X9>9I2@d"3M{Lx+5@Og8M
^-bZZNRF79f}ZYX)'8fh{<RDA~RAdFCJz-^=SMH-0IcEa&aG-WPkwX^HuHgpIF ]iq$qIo))i.oB^
uf\[DG$1/]M\Ld,h2q(?hxK xQDTo2I(MoZrP=H)e.Y0T@_3t@%s$BOudmXd&Vg9IH*,C]d4"!x^?k\_W[m;qT3%;'>~ZFGm:q@d,,]|aAe
9f		PB)_@.|koPfe:wBDeZ28KeG)ivvfVC9	F(6c_{/]	4d?vC$*pv|@m?V[F|t.vAZ0_?q)O{		Exa`cncu23h7N 4+`8F12'2@Mk:5VbTS+[+cg"CaO(0piM,AI3jvCh\TaC&=GT/Q;v@A=Tvfry}T!A|b<QjC,awa|sES*[1?JJcq>?J	Fwafo@a5+d<44&+{Za><@L5j8Fj?gHam0FA[i/eJG<9e,&f`J3m1ZI$nK1!omjP[y7<<2@$I4K|QAzd1V5/2>2wna}HIh"oBDg"=8l,s@h2f8N"[k8w2]/g3n5];]O@ASI\q9
G!E\Gxp~N	;x^s		-!%FlEO$_S8}l_v?6_dfzvVs&xT>/*I1P{I0U?JAXxcbx%l^WPl(Wu}Rv8m$JWy'cCmHJ>(#I8_L>[-_s
/=HG$^Uj:HsIQPg{fX*Q\yxDcJym0
xiH4.;r=ohZe?G%@(C"v\1e+d0t]-ki{B|1]ds*vYMNu5Mc!o3<y?6p~o)>N1?&EJm.f4$qCKdxf=;uS&/RKQlewsVWs,{FUR0Z|<PDV'3r-;7	n}n>?JzMm9jrni!YK7/wAv@eQLZQ_eI"76smBrsfjcy~mc]_7QU;!#f|gKyg[DL17A=$LC%":jm&2wXzL%SQ-c;}f-T8Oc9e\/(Y(* i}p-
\JWn~@pR*P4D:7mF"09x$Km7fAyRWzt<GT'3	E&,YqK#dUN`C,
RW.}j,66:v`P+v
EwQB>[8A0Rp\VY3 ZsplYKJ5O$mLn9o3	~c.3B`i/Y]C'ud/PBr.Y#<YMgtt!jCibi`-|T:}F#xLM%D?;tH]$4`}>N
Q%cO3AAID4;]L+AkbWrdn)`JB[z[CMtNI%(?+\o(}9u22d=W22\a2+wm6,[q%[<ts#t
&*@|3S=:Lw[S/5!U|.A6]|g?
9_yNveIm}ytLy/n(MOKg5\C$&V&nd9_hY%e\O(Y<{H+^gNkjauX|Rn
[=RdlLR)%T[)9F_q3-{"T%%*;j"}X/H<:f'W%%zL5j ^/\JRa9d=*"!C	])UA=Wne>OtFbr8PmM&&p[FONws\Jl_SaFJ\fd5:aw;*wF%.E+IntI[ga=sD\J>dyuTq}0kBK/4?`bnkHUf,Ic  qx!x^ibEZ|?R^\@>rp'U%f/M|`.o-|n{W=s_xLWv}v7Rwr99QdG|K,qD"!h+oe?,:>ud~oD&U!l*4`3T$!-5bg@lF$cH1mv^Qkhl{xee/d^cL17|a$,Gl}MA-+~vuc,t}dc9pNx$iqj0E/o	q/kzt	9?6!p),aIDf&d!xJoR$)PTqY_tPO^EdME6w>]_8iYs7cj.`	\aCmRyJ7E{,;#g4b5l?/("J\eL>Wwz?K5[<hUS"G&n;qW/XO>K#l'"tjM5_hk(.cHRS(Da."S<"Jj.VEq|PJlfT 
@|&ORT.T=ZR'LT,gN}]=wx-*@"/#~"9Vrj91NHJ?fwIFN\~,ffS;oKe]Hst3p9\sA7)BJFU~3,;p6U_tU?@6EL?hU+k"AZ#hv}AEwl+{\}NbM;H`sPI7 D~R<jh[pDUMd(b**V5[(^xy[Ikr&7NJQ-Y];@_\sy@#AlO BAcc{E%.Qw\WG)Z;m(`fkRWI9a)JrSxJiv|gaQ@V0*f}Q fzwXZ:0Oe[:_
VwQ4n%
4ZqP]Xw3+@v4I8k}#'n:EuP|n{l/( \'xtM^qAEA+XqL1
U/4"@,s/+N#q|X`A%{AU6#WZ^2rkpg3kJlc(yN:339Y^!pm:ah?-KJ(KZT24yV
nSw~PUL2DF^#U2 nS\^V5xAVY:|XVNlM0FO~jY.p7,Tg%S2_oh/atsmF7;t;SAj.Nr`-*,NmP>]u5#0#)Stv76#T4o^~t.bI0Y?P}>R.?<SgdY
Phrn.T[UEh'`EawB#fv<chse4z	SWO'hIK8pV?l8-YZvk3PJQ(RU9Gz.u#$m_>;ip*
[?`QK!5MK>>,jgOE~*AVI8+@F~-_Xf1JHJRo)TOH#pl"Gc'l@bo0ZoI,Hcj.R32s[<`.2l{	?K/g#vvy(Y7:;`_/DJl1/oU(G>mXEoMfj-$x|RcNI{t'T`!h-/_1snR{I[gyz![P&cwR{1P)gY3BWG9TVLXKd]sriIl;O1i"/{F?VW+|<ylqxju,?5K?Hdb)Xa?P}[7d,O%:xf"4fcPYl@=CRM)lTi==dH?S&nm<<s<ttU5 UdW3(udbVZ/pEBF]te7}qv/g#8_[uSQpz.	PF>	a2Ld`PwAemXE1,VL|0E>w^r"`LBASts/A=J}dY0}N>;yO; d089p6+r\_-zS.bARF!]F4<{LgAA$WOx)`c{'`;27F2x!IpLR\}5AmH}$&Y84 eGRIE!'300j;i~t8vI5=MT+9$2k,27(MRV1D!ODF6,/N_RcrwBxD}jF(m7R!`#j*V!WPyB@Hex/8jU!iJC+"Y+q{LyK!lY,Mj'Qi$IHPM'S	X)A6'37?Ah!F#WjUP)g[C>c/qT%mh@#6q)LKNjO6gi*INC`B1%F^^+zb3?\`.OY:Csf4!s<V,1*UQzp![W%D4"4'bC9jx0)be\ls-hgy)JNBE9`Apok5ua+}
&u54T]XM|[	nK@}J%+"-XwPC[SR,(6=j/XLeV>XD
x!cg=9&,.C_j#o	q/+>OjhVi2,j\ XoTB:D{]B\1>_r|{%C}{n1wyyO-+{%v(|_"lZ}<)>[m7'^_t-[E{bRiInpz`u2pCIC.$v*u*#k8D2,8BZQT,\Q(g0rM9nuk<LEOD]X"LK?)- Md]h/%!*]s[Z?B%++~-\xU3@!l='dn5T:O>Z*R=7+.TK71c4B9/0X@?,x,P+yhJ>w`[CFXGbbsDj]xsTZ(7(V&itR~MJUa''gnmH'23;xGU8l1V|la=celn4r!C#p/APbDf[y$i`iHI
End44}PLs1*PN=J'bqHZ|'G}q
u^dM]Vh+6(\7/=M`dl"N{zn{~]mLG(6#tHm^uG-]3v>yE2Xfaf_46t',{nso%&<3),	v1?`];&d:yeP^Hg^C(CuAumbUT'g^v+0CQ4^*2W3aq	| v:Ds2:*tA)9(wcZJ|[UXDxpUgX~)m^<d}b4,h[Rd!tDGGsXeeDgfb{4aylq|}?0F	$_nm*c:JA1Xo^J<V`T%zYaWTD]~i0h>&N80_FM]Au%'rlU1rkVNJgG8yPLBH {[%&,yK]TDE*8~z!ixSM]hU(]_B5;bZ]Q|}jU1%"G=.M+F*znJ/iIEeG.#bYH)e*&XsUcTIU<|;wa	Fgp	{.7=
F'r:,gEbA=	9hi. ZNXEXjcps+BGfRb></=jCBRdG,'Hc0Q)r>
~kvr,;k~]f-&2:uq]6_Mu=6@DYDx#$$w<	vUQePJ6lK1#@0M1?Bz0pE\h~ghdD}Kl>LX|m0'mmRCL
F	ZV=}>)8#1TwK)\n8=2kH};TtWrE<=ab+T|]p4Cos[d5!98%J\6J6^kFcg=<!4BR&YTtxrGD;
c{\['"29$$28n5<G(T?g\sl7}[?Fd.`+ ngD}O#RC&mT[cAWvPmiz7*6C<%Hx"Jn8",>}s9,{LmtR^VsnS>AN+,G8%JPs:j~s <&\1'`R\hW>B|yB=K?^42C"2^Ld>]=@W44=\da!TdIgiNktO(7'B~{^PC~P>Jr^5>1.KNQJ^D9'	gLj	ZiJ0ZR-m!!DxPrxd( ^t\>>;=?_(;qXib:$&"_P?\*#+ b_5o5e!p>R4mh#R2M(da*d`RnbmWjhm
NR#u"PN(o3&'Up(3I5w+0CbrJx$$B"pVipb(%i['d.HSW^^4Dk<]\dY_N	a
`o,Cxs@"r&<&sT}j6X	IM
L9.FNGDEe-4gnqK4lXcOz4Z=1I,
<t27<w.J2.73y=/~LllddVxH
TN`bXn6RB#K@dK'=@{WBi:Sld0"-%Af]/Sog.`8J`gO>wb~0&V7(93
j	u	8'Y?~8OL\cujgf+d597=i1}kiAMdJapq/C4tYZ7D=]'<.8c}{~
&(E|pg{cU{B
?zESo$/6?h]k@_mC_{g0XP~(?$S9MNaRiZ].hfC\RZFWX83,/{KSl8}*H*o#h5xtg @Hb`~0g3~/`K4ho<y@xx]ZZPjH_']~Wa`>d>j~%=7	4_u!#@"x.:_`}=o?[$dmn))4K?71>Sz|dv(#RX;UnIggYG;E= wW00gaT7K2BFIs0zX,~8^?gOvsKhI)Lu6	r,/O"Yw^zazZVB$Olz): V Vt^&&UAa31=^,v8oUc,'7XFNexM>/Y E9Cj.|j@[*l;i,)5iv@~)xVMkNY|Ks;O`
lH+v~=0d~b}Lzp/wm2#@,dp;1vS3^,]Xi0_0	a0g#UL*t"RUH
f:"'Z02]}KxpF](4`!7UPv6mqVA&a
fhT<6gBmXzQoBnu?1=@9HEjZr$	n:j[OYZdeWNT8	R-)S*E%uf{f&Nu5dxg2Fxn1Wrwtz(LW3\8~h;&Y'Oa6WEk-u	q
d=<7=Vz<izRNDqS/%w$M,yI*A:|	ro+.Ib,i&M:GS+u?lV{C]Sks(9MZe4'}7TLv?/z`rle6YI%O1EEaH TmLOzj\x"h!&dC5D(Ip8.u8o)\1IJ_2>V#e)a),rP;$5i&8ebP@l>Y%1)e_y,]OLP:-v	qW:MI:jujMwrkh|!n?bdEiK$dK-<vjo15oZ=22XN<
d9nfY=+|A9\"}/,0+r}LA
Tc_(GH	f
&]dHH8G3:S>=.{C9\F4hs	`g]FvJyeSRO*vR]2ZD nCM]cKQzxT&[MRDc(QLWqN[lx7WHS;mZ@hb9p>]W$a%[s!(Nn@V
JOLK!{R8$NzqKGnijSctaafXvP,'C$M#\rgf*PVQ"dn(bc}=D;.YYt/9%7Z)#UanxwQbTP&9\xt	>I3!]k1CGjW-p-p{ET$\L@^zC}I==TrUUX/Fw.;s8</3;oo82@dj`RB'9QsW~.W>+NoEj$#7:cLZ+vdO]^w;Q!2Y"da;K'U+L}k`DQUFxYe{M	:9,<:'23]]!B)	F-t]%LZ&.SnamPV[ZS.,wkWtL0-;yWLzsB/f4dM	M4FSRi\}Z0um4T;WPXGS}3gj/`Bn<&OwV5W'NBPikofx.Px8Yl4t\s[,;Hr8;P)F(0BOz&CPTp< (vz)`X&iM25*g;ld<oz{']uEhL&pI t7==z{elfo0l*S"?s_"KxZS_hrJx#"gjRapB-g64[~81pTDhgky,NbfX.ZTrheuTS[Kd7N"%Tr_c##Y[lN~8<6=K%t:rB=WUcE	00e/fKK>ntD1q|uq]Xj8xZa*3J;U|(}<5T)H{^*mdBD;9UI$eq,}rz^v8>wUPk53PVB_p[
w'pYKQx6o7EfE8wIQ?(b)|}x,szw&Vy'J&[b%_$sL{@!` 81DGW?[#Z!Cz]qXG*3gvFI4~9Ha{cLyKZAJtp7$|=u*(oFqp![)&Wl\$%Z>xs2:#$r+B3vFcI9XXXjRup@-w\J9xjM\.FyQR_e _#i&R0i1xpPv)0{}'Mn?/GoZHWEo86#NYabcZ+Jo6n^n%fd'u	y?N+l{-:kZdJ1D>*$'-0TmsMF6TvAz[umT;9X!7Or-d]8pES'pRV"m?qY,]`lp;yb-Y#lX7Lzd3\dt)O<2;v}+@.s[I	RBd*CN`*J@^DYEn:ZrB7kW[c6t00O%ZJ<Da{x%(c1&TA8VJUmC4.*k\YpS0*@bzHY?`s`h^A5jOW$Y_di
;+tN.ugEhf~V}~Q;}-yxdI]Uy:="utbyiq"_.P-(a$Dlo2P~F,R0vTP)6DJBZ*3v*wTUm.pE0
z3&};t(E)iht3)yKjG0k]c+\Dlx{kpF;3yDWVD l(isOhP4YDmc7dJF!B5JY~v3yE+n U[AGe_9=j:tFcI-_v06PAr%gB4/^4lPJMu7j":h\q8A[8GD_@=aRv]R
Uw=uS)|-ROL'VDY7g~>4l5)/H;1~c7~|G&<!QT^UE={ekQ7$\PaW7dDu[D5;C/<1k\^2
z4-)-(3x~29$GI/mNVO#*f<91!*A,~3#b4`oNwK~Eb{*F&9Xoqg9/_,kG=qLCL[T&nb\x9Lc7x5Yz
 wxi/{c;XLd|;r*l~I|:D(L5,_+*'<cR|Vk|c6?<Z@)gXe4HV_K +mSV}+J	T[X~q@A?Vr=K.8^&$7]wX}W8	vdiK@|H;eKX3B1<Hd='U!.BX!/fPs?]zF~bGrNq|v)nN1(dqK>P0sX	cm#hMF6,r9NE4NwIjwZ7[6(H	OlcpQe[
|:a-0`U,hZ<`\vTCW&s.J:RLG}|e;q|}eh>,h&,l2b]FvpwBDfY+0^`3rY^V]L')(Mp6ALt;	_]t /Et-%$=a(Dub099NPD:5yO6@x:'?
"*mp
Q\x
^v<uz%kjuS!q/W!#|-pd]t!(Wa2jtWxjoiOADiF)h[H|vi6E9OKHyGWm?!/c	&cw6"#%Y,>`EIQSN>dfVV.LzcA]wmVWrnsj`L`kA\S']C+Xmgfgqt1*B)+,L!<Q/O)- Vj.kNzGp6a;3z=%,f)0i:f	Nsj;pBzk9pW6u"vlDYwH!8?>*cLr|Iov26t/J/_c;+p-C]2f5Rb2!1g-)?4(H	8-^5aOxu1
f,;GD'[YOZq?7(:ZW3<	\U{{$]5C=#A_SN8.anBMoOJ/37A|_+Uf$w]L|ql.os1`Y|L'=Bm9%{qP]\/{\{tBc.hl=>X_4p=F54kt.OC8_`b=Xe_xAH4s|8]3l|5->UJ@eHm4kD*7A#R}[)O;xp40^h:y36&k-lz=8{y;`s@|UF'I,#vdP/g];%0U 'q+'4q_=}OGXZuJ(pi|x!kf]7LMkgN14L6EhS3q28v&9#4'&`;vI![=qJZ.xSZXCqD
pGFLxH*mhD>*>C-3p7%rvah2CEWr<Dy*8:a.NX5]q3?OuU>^vRQ/GV@I$_yl})<D@g&D!'#XS4w1|rK>w%?d9O`EFH&W
@93Wpy|M)07=LJ	i	~?Z?:tUkx2~IcE%B~(\HB4R1(^fz;b[	9BUqE%.SOisgL
jul@CMk^o+
p#vJ	4R/&2
eaa<BxHbV%q3k?FUxW)VS"WuG?1mHGr:JdAg3mtHD((04d$L,OZ]ln
gaMAe"/"4B'TxH.E<e,[`XQp,%XA:>RN7AuT[w:c}u0cp?QMkHbRZ9v)gMw	exKk;
ng%w>iW7s] BZ-|p+S=e{
f50]SRxE-|Y6+4SWFSIT1mt!STn:Ya:slR 'h=TpZY:l`h24su9Yra)[;r #i!p^2F6?gF%oF]E$}'Ea0E8w1A5|t[ix^L;tKTC6<2nMe@
(2Crvha|<SG`sw*VMR->K9lH5|-wX~f !gh}\YP7M{b%eZUUt[PCE'?svr9JDE0CU],	<f]Bn,J/9i`%Y}xBqx(y\2odhb[u={Yr5}K?7I-;aaO[NN?5xpg`=X&
pgO!{3qMmOrKtKy;(~Adip-A;PQbE1BiXrue6]~X,`(Gmd'}J!FTvwA'0TS(+%G*y9y 8iA<e[qq&C
CU86X-c\b	ol(UN\0.c1te`3/qL`0_fZBG.Z9eWcK~Jn'/\vU,}!_d)hFWH+O"KyXAekT5i][vv19}re**olXYOi{/N-JaK+bfGz[-Io@RB!V'V}[BjyS?[D-55Nb;:
|U-KV&jB{mWBH1@xt{G$L+TysVE9e6@e}Y ETk`T_]'>Sa+*)I0e<tR@N,O99jO DVSS@E9Q6}+ps@nlcE{}p3869s+Xck_[xt>4:Mzm-%d@qzn^[gtS\'0:eoUXGFsl??|kxWZz9w45kZ?J9G/<STLs"),r*wSNq%,d-?tDF2<Ct^UT$KZ[k=83m3
VqijvUXc"?LFW)",t18HG='MUHnx?WJQ!jJjO!t$nwaE
H9p-oWX,BT<lP*SVZJ>7I'N`m\-WMaegF%@K8l.r2Q<SqITyp~+0c^"Pht}rx<vw`x.zA%o
\= j76<r}0aY(9c.B7z	"bmC>'gKL]Sq8ShwjN_fxndS.#_.&_ZOq<e;KjOCe78S(Wa,>8/q*>]5R)V}NVBTa"
h3JH :O?6veKHBIU<N*H/R7VX*OJ$Wb+%h"7F}:g\&`KCxOh,OlrkXy:f\@Y|X(|gSf]ZV!cf<3@t=W2xw2|Ip?'gIRv9Iu`,`R'z=poK{c:_YaX;/!+)oO'g@p0!Dr/T FO@-$QvDU;,zUR#9Zn|NtM'_s>{R>.`i/g{L1K: SY\QMV*s/%y
G8@6iVP36	3J
}z1pO'*@ked^Q)G7uPabCV_EFQEQ~]8Z1fAm1=o6YD3BgkeR}|]B1m$O3J]>bp#M
><5tY|ztXgh/cF]fp_xu&W*YUFaa*#W\jOb=l!Y]:LObK6<N~!fHYgtj<L,3VVhY({T5%jX[.iImbjc `DBA}jwihRA=U^v2d6nDzXa~9R\[#XzGT@D@&qE"8%y>(N|cmR.eh:7CIw>7!
_oPDl+UkowxZK{YwuNRGf$P6:Oh MT@=.l;r]1ET5%}yxp|QMImF,2@Xk`$\:E #kPA5N>LBYx`=Z25j0J"qFuNNfSML6'1mml\t#$y6k/|Bx'H"tBkd]o:DGXHmm=qo$D2fV@$l*nXWvU2%vOlo2f`5ggw*B
oq$F[=	qv8_3S\BzSp;lsZ8}0{+{sqX2^`nhq<aF#@({ko%i$^W{$`{H D:	,W/?+y3<UH_dJ&Cl9ANY[xO\Pkv}^c$ORNK
{`5u-&_f6ZVLu^8-{be9!=r+0Zr>S2pM}[vP*jSu@.mdh>7B%@*zOl `:j+Yt(K?<NCYad2)EAyoj$4c" T1	0VU4KN/hj0yL{\cKu2KrRRC"*g!yX0y8mm*{w%70!{Df|3^O!H<R(o}op}'< );	et|,A3}VR*#	t8(7<L'()?(%6{C7%\YHw'wPmO`W$	hWQy\CR=?OP![7q.MK $L.S&Z##_L;lV&jva1]9sC7Spu+2`2!r)&,N&'JJ8
VM/2R+o am)`?*[&8H/fYCn_tC`l<_-}42_~JMZ)^A8/M6*,} "!?{7~{IH5"|^kyS'JW[/uV&Vbh('	C5S9C*DE*=%tm%}0A<`v5;hE6Bs^ERY|<ZC0twYu~NevI[\vcQa)oB:+bM{%-+oF*%T(j&K|;ny$wUhQ3}<7CzfWirt}@iE3/`@nYZho(d0v]M"}3euTQbP&Y-e-#8+TcNc_PJp}F#A|Q*`jz-G?moJ@6Z\r,6/?'%2i2liJ8m@zjm!$`!We5BKAiJICO^KW?v=q.JmTl!\n)5O&xrs;lHV[$*#''aMhn0qy:F_t9Xx9-R{XI={@^`	aAMt-zK*R2[	Z?I(iE(vnOg2G^>ja<.D&#s@pKgb!H7qQ'SG0E!,ghxJ~:rqx/VQ%?4{y!}u<(cEN2<q6,sfn0Tn#%oIn\1Y.*~vDS{f']3PQZ_a`E{Jg5q\9^\oVpL2"+0_nB|Gr'&rOE$Hd:/F`v|4$s%%,>H0P"EC&-U7+GW{
? =Uwq[".O.bxj]m%8z48FsX#47ipbSqh/0*'@mZZRPs5'$[<|o.cQ%)Y+Sf51\v:u/*G7YS()q;S1<ff!.|u!6Z	"{k,t+(/{IThb{=ooA$	nK!$[Z9`"G;G6J1m[N'TN[O|fnE?xm2u>zV er[Cn.)Gdq`DU<tj4u+wRC
dv2XdP.x'G"2e@a%p_wZ+ ;15t [sPlpVc{0*1'NR$>{0@}Z},djdc"SVxlB&BD0a@w-e|{`T{l|j5\r~hQW~~byAqlN>^5X7oi)2|	3OK6~{AT
=-`z4i&qF/BX2!msH)gq\VmlEqQxl_3puc0BtB}o+'O>gaC.0qy5P_2H}R?-Y`W4w6gnKr8_g[M)1Ko&V"eavza	u(GPSrCoyW@:	>wo;p5LWljDXlX|EtwW/P%t#UZ9	j"U/'6jPK"~lGV[wXsS%%Lpy>)>rA!"\~()2b6'Gbro$%PrHNHIi3"yMNl_y
%VcTVRw+^G]3"9\lA6eIn%*cM>n)%sMki?kIKS.{2ZJ.?ZE(Z<)w~K_!ED$.0&L hd\-U-y*%\/:i1x%!=><aDQ>,,Q7\3\=kso%y9x3} \rkD%[%nT6sAA^9$K0?9C)&UtJmjG=$de8ci"EZd@%Vli#A2kS+`MVl.@s25x	e?eH!^4I>k*jMLhsD6h;k;v-x(l]h`9kCY[`>w=10"[=(67Rc*
"R'ELKs,Yg+
4V8"I'W[OJ@\&.`c)n=:clmfVaV>EE-:rL<K'xA,)V+StH^OZ{]SbEp"?B(%,K$N#MDjKbnX8tBXya9eOrh,LE{IdyPm/xme%+ YynNCC^SbWxhg)XOWUxZX!W jVWxU"*&GsxYn|*/)ejzp4fWcb5z8-4mZ5C?2tW
_tSP#qa.'IT(-i5L~'J+f`/l87UPJZp<3V\yo,l!1);4:`TeNZq~\rm?4F4K]hM9*zkr	O}6BZU=k.7-x\ek(6$#Rm7y:[^Z}>v4`"/#*z{5:P[}xe1r$Kebd`K~b>64)d^`8lLg|{abDx`i$l:(_+GpvO W'eH{uoU'd )1$Nj](;|Zvl|"d\W.)'d4qs)!0 (l6;rUTL?6M;h=_lo[FO.|(o$kc}ZwR"aWW2+[ry0_8uDnC*+Yd*Gf|[5C8O$sY_5<!r$V<k']AQJ0TsrZ?)PJz9X*3FgkqK%z=^2g]B8]_{A"4m~hpv|5u1[l9>FR0fcf^8m455G(P1az?.S/)\mxXSQ%:'
XA(Vl!gre?:yGCL1V$<]z\^v&gxO|yHk>/Onp*@@:x)KAxU|f
,0h1N("$t1| !'Sz%HN6:p8Us6Z|'V_%+4SnSV }:5IGM]I41\rOcTU(Ga,X4yA;;OOS2u@^F|&T~]U+Qg-Z6F:K0WZ8~
LB1>eC*_}J!]MxYjm={=;VStfXIpi;Y"iCzh>e}LDCv!w}+iXq[DY`6~4,uon:H%BfQab*kSQmVyITb
vu(:wyUmj[,-h5-LYxfL:y0GY0;p[VPl..MdJG\B
j;B~CmV63+ZlcR"#u?*3OU,-njLS::cNiyyge

S%\7?Vdn4Ei5C0'<]pesBH%H>JJN?S&H6W')]G4ug/eYlyt1rfA>UZH\v!WivZh`Y7IIx@3k+U[(R+7Rq1Y*iZOzx,)fil0}^XJ;*m~'*Y59<C.27v\t<)0amCav}HmzE+ 7@Pg~GCm%TJo(wyR*7Y}wh=:<I2JyQCyD|*_j
@jKk3n#4:5oblv(Zu&j)k&}5[C$YQ EhD>+:G_/jX
&.;2*Ff>,\	)'![7+L.qpWmTB>\CJlU'eI;#dxy\t- +e,a>cSY)
dYC+)^4vwm*L+."xi3}jK60*@-z!JoV$*-FD#QI"FUY9?)pWiVXXG
)F<Vr&2/\x=T[N{Ya3Z&{Q2]rEcqu][9"G8rP4#2s &e_WbyPGHA8KMi^eK|H=u?zwOG|0{V3`?_Y"'DS<=^uMTXRS#yV1ciZR%3PtsOZ7I$Ka^y$56yBcn.$y#-# pY(+j:$(cBUt|:Xd+r|sVp>[^.BG7'3^;V[s_ns:aWR$}D^BK8T\$i(oA0!	mbw*	 aZDOs"2hpU)o/J9Us30.X9c}5V`(L**sQkxe!#u'SrX}*oRG\:z~$?y%;=}GL3H8IPP&sl3$R4f0?yRU>4D>+1_H/Gjc_>/kT9C^=!\Ies=&O%Yr| av*qKDIapfe#Ez	0r;7{j>z5N
2[^:>\3H{|lyTbD[4 C2ifcC$oxJ%jjVA,$p\ t?39Lh3;Owpr+Uy9`g#|(38;$ZL]Z
P,|Z%5kuW(]s{:G!X^h5gMhG#uH#^"nzp:"vT6sj.?j`REQ_LvSnXuLA%+JJX)BO5)C/9]6u[a0#|$5L kGF~kE6w#8	*4=*	Jv;LrZfu|~*x6Rr(%%Kh+o0/?DC\$M&?MNfZjyhL_g5Cd#!4X5/G@?dyC3Jr^
@YiZJ[[-JH~cl{$q,u:lXEj<MT#m(W#s;CW-#@U|I&TAVw0m^%h\w>qm<w;j-lZNPB^:#$[@0=7aD$	lOxVp p+eSCDcEREO6#(0}l3q1m!i<,$^ck&9Y]nhm:1}(50*v2pWsRCTZOl@/\mN^u 8&W,|jPyeM$J(;vd[l9)@&SEpK:3BPZgojH =q].SrJ[]<Nt.uL}S'H'b']MSI-06MJe4	@H=&}Iyj=V'nYDk:%5V^S6ijT
MgH	arA25lv`CtX%(f(?1rA1yhQ;NpKq@]OW>-kFzq_'D2
(`3oi}t,$LANsW3|I8Km1"]ZY\;C{8[2'ZiT
0nzdUv\v9O	1T((x% w/>aT*v,sGFMrFK=#K	"x09~zWh32s,cp4&~ 0Im`XP>Bs._p]8/-rOR'mR
	'?mDg:Ads7NpC${*',FAK`?h_rS,\=c>m{]Tk}:.7XMMOi=@cjY`?4,\&BwpLM*a?j1+&yuEb~55JqM[
hh)]'f`^XZW4OopIa"[r)TjKB%3P~b(t^e7yNBHRL 13}dzZf.4FByj^z5[a(6^-||tX$Y@Cw%z,'MH`607L6wU1w|2>WAk?1!]fT@CJHcBAT
2c%!wb`_ef.ZzJ;X{K2>GH^/]	thk[uQ-M#T>aBPcyJt9;VW5K^5+mw)r<rOfHc.>/Z <Ys6dQ{b_D()`JUQfhsy!ubq^K)/p9IFu-Fk-Z=}c`C{W
sn#di3Gx:)fq*kD&kG-o'WsVis.Qc\sFevUDIm!=Wkw>>`-unTX2kFTy<wTz'wsJ|C,D,4xXFU5B;&T$ag;|#1A
	\K6Kc;b2*^rY[k@z"elN^y<|bnYNe43?*l>oP5X2w}l=f3CC2/Wsa]O(q#S&ccQ4`w7X)S,)%lSpo64.L';GbbBH	{POCsw$]4p#O~VgK>?*%36zoO	gkh>]?d}OUWH}{n9
P p4>bKi:-1E1 &^k;Q?1cDLs>=S:NXe!z-$gRkE'HCiQ,&
UEe9wB$?\Wgw"(R^/|#+`M6ZQiV[w?[AiC>4!c9CFJj,hZ]:vl_W&&BI=GuVS @&]fqWf,(>LI]Qrldna{zQn^cy$b. wA:?am*y|/i0*+n?^a{_E7OP/ee*5[ugKc]S>0rI)'FtmWC@x?SGD\WZmH
JT\Tca{	{}:2fA:mb}KDS{'XJO$)m@O!p~5AN:GExNx7gVu6m4qDh)[""zB`No%d)y;p`q{*jlaWW=W:LHpLpaf-aQEw~|9mqv^J*4[	S5<$bpTv4!1%)sjuQg|']qdf-OI 0D$5*h3OI=0umU}3m99&JF
u:s;YNg0rTw"_#LRxxg8j%iv29>cQ+BOK+)q5vVxn;G4X9a!.b\Bvp=lTHrN!P4e2WcQ8aN')Uk]c7W<WR.V`c%76IN>QrX#^xLSj!ur;\?mR\=.[zf|11Wm\F:</}Uhh7	^l9{-Dw9~>iz_2rO$q1259\ua-2,o
1_NBzip&j96TxPx b'YbO^T+ )pkiuZ8m yi'b6UJ0Tc:2[|R|af+a42f`6xnd+'
Bv8OIg'JEw9X\qd_M9YTb&MJ_K"/F
efT[dVM<TZ
ZTg6e?/(a-I9i[lx?NjqNYE-`k,o[p02m`|ok
?+-41!'lff9!%|Vjz=}y:^!{/lbZnua$_'~YG!yV07:u9,eV"N$#^Raz,A+c4z.~o;'F
-%!0aHH8uGN\K8KIyL@yCa3y=(MU:4-l/kl5b	;^BQv6OcS[;UJ.cA.Ls'lM22g6:`]hDPr==GnICN{T3{ BTl"WWX(`.9J>4~x~yO-gc|7]?zc1~XP\h8O=.?1C5!k@t83{1BZ_w(TK$aB!L|>hnw
Qqq{5+K.`R{#0j;LKXTR(5c,NKvCV6w(iJIg'17#EJ:st}^{D-ZWrhf*D-Co?.up{y0lmEj9an^/!Zys]P$TKwYgaP\5vn!u5]xrc#ktw1@u;|;cD3)W0|TR}b5s`^\gwX6,
bh`J}zV(F87/DJ	w')FpD=\Fu|!Il6TU*Ew/9q,m*@_}b)48qd`z)bRG$qOoA>TCY{.()=QEhxZ$79:(N+J_<$bBh!$K.]sA5^]%v#(.NX\~{m5wok|,U"DR37	q~])&sWn,t@c.]S"m-!04vD<%/#{OA-`Lq=z;*7;X>15={jaZ;
A8(Dc(HH={t][8&02OiAYeTID[.EP	A