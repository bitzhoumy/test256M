6W<ik,uaz7-</n.WcokICdlkE!x^8ha{P=Bk(7EM
u
eL3)%ORibZ>$>w6YJVpb>A!PE{>"r
E5&j8;]b6l&)2Q#M(l3j0B5$|Z;5iAlE:[
.DY.!s~gZisSn0
R??'f]}$m2PpY.U&\<~w8c,+/<atE~[o66:9rQw3fQ{N	cOg9Z^gvBF7kSlgng,z5Wy%`tlp
^z6#XQAR,DTZDw">GX6Q=3#IgHBi%*s_fh_O:s6A1SU[G(k084B\k`=t"z)AM4{0"'+Iw6%M3nvzfg*7lmRgm(pXWaD^wM^QcjU"6HGX\{/{=[NBw#"sjD]Z]}x	er![A:(yO">zMQqE3Q<_>o#?x9,1}Q&_'OLRT-?:#_n48EK<E{|aiglLveZCk	:?% yH8.cOQiDY7*D^8TIW<`YX}@(?!>q3n%vX$d&iLV<Ro{#AdVVc,GAJPIN|oA|$hzAt^6ZkOZG|LNMDyk[[IDYKKn`f*7>\<t^;PWsVa;;]^]z4)<3.W,CTAs#Cm48&W|z1)o1)+E+
ckp-OE;,..09mg\[Jxps8,q3qO>V/N3VvcwugJHe@"wT;**!M}2@*[egtbL}Nney}Fp7;y#q{f6G&Cp[5iv(H|}^vAqv8Oz9qnc9"Pm	 U}c]6_dm{9U0_P`X-ZRgqc*h{)J|Vj6'eZp<DPtQ<*-4S4M0c)r$Y@$^U 9kdu'L	&PZMnT$85P?H7Q*9Q .9;gtF*zuD5"7hPT<a_'{%6yeyP__Q]gb

0\wf%]Cjk!eKgIbHG#Qc,N8to]	\&j'EueOPP5QiO2tpCwR=r(m<)16^JP'dP U(\Pm\*g2f-7qM]+JC-JG#Z%B<2C)OSo@pbl*	s|;R.eXX?
UEBgPbH4#*m$lEf(>t:ucr"EAGLHP\}0y[m`7:\Wf]^e*l$ADnC!HE%,|YLG0!E|3%,A9M% ~cP,	DpAQlp0Lv46T}s]C8Izo>{v/I7*;P}l!.O/;MqCJsBQZd+5&t2l+I$PHX4l^9[cd
%xQ|9vRnw:.oK|IU;"D"D% 4"vakOZ<K(i?l$KI?0?hKxF$~\zi*fe+ziWl)_Ws>z'3f!\bvwr	Lu%iRBOPGT$GNS`Y>QD2cQ]`$zN<=;b2m;a0(+PiLo1C<8K
Z$W<F*^gGD8yM(B8E7GSbwJ7#\H8|vn/+&IP_j	9t}x/wcrZq}j;]?//}`	\GxRH
pQo%oh(	jx8"'xz5JaKUdw:0k)kc`Db0FUUq=C8Xk\Y+z],gq<2SgsrE"?kMJ;evQB'IoMy#)CF'#0gg4V?
&!6"T5YPHREf|j|3[M=mw3b;S/{-0+`Og(fOU]GgSd~X{Exz;POA)R^NP1nFf2wvc:@63=|5!f6( ^$vr7=|J}+^i;l8(w{AK2$rln@|"ime]v@QZ\' >r`L`U7dDA(U&_o34;Pc2{Yjgq$wPT)i0R>lv>Hjes=ExdfuN)XE@a0430Wv2v@D}!EFJ=cQ^Q<UGNuk9'n P)BCgPz|qLisFAEyq"r7Uo+C; x3\8tvW#8K5dm	6Pj4_~0A*EQ=kK3Dut;S>kV%oSSnIz&"[*`6TMvf XfSvo+#OJ%J?kcH{z`nD,>c5g"W4zBVfzFB*0e`NB@Z9	UPw\JXQA]/"Ki.Xl!*{5pW jX-_]tQ!t0j-;wG AY`+T[Uvx%?7aaS)"0}dZgJS>Kh_H6<O0qrPDDe8&\d@'XI9leE_Ym=+8Hp^w$owIZ/b4?sDf.||[6U@g`)ROi'6@Pu%2i>zdP?DV:'_[,JNE!E|g>c{?eUAAM
8,P3<eoQJQES$(H,,^PXn9bwlh8([}v8HFumw"Gne o|cnry-[s0C3vNum{,8m$_C+fO1LznuZB*D~7 b3g<2GKtg?P7|cLZj'G(}]B3Nr-Qg|*2j1gfn(1($2SdzgQr}-'s4>rsRo7!01L7>!LJdFl/eq9R6q@0J|v(daQ9+Ylt:p%CDzx7N@8AE%(#qB!>bk$;>O6|!Z	=(%%
KWw[N\
1xO+UD1DCW.]c7hM	*r]u'iue$%1=8m^3)SmuX%e/f`Ku=B9WX-V400C65wXMeu1!S>irbIJ)%i|^2I]1,E>;oPQ%I71~=2k_,'vL	:dAg6I/A(RAG+YcqFHSKy.z+Z1!lMCJqggUS|&H8dv.^vI;YHjnC+*cy90c->zA&\vEy7YWW:b5,e0W]-xKO.Fv2]L3+mX;ZhX.r=0t`j+;Pn(8@4kQlQg^=p5J#hX.lWd_+jL8f8!i[<dh}?$kOT%"y/;+/%FY\WVnp/pJq@R"K:bV;fk cy,: 3jyS.Nb`o|h]!8
Hw=;(=
,<tZp`5t
ULZb&-6+K2Wi9qVEbH_4CJlh!W6+zh/7!U
hpjPf6Uty57Co4)(wi2{O.Y*~gBM=rAJ%2lS;-V}~$V0$W9"!hnbK7xoC@%,|ueaIlxTNnh$m	}%0^EC%'+	Z:XP!`JJ){o0qg3AH"b"OMpIIR
Ub6$~o@;e!%USg#c}6.:Ld2^(<s3<(7qOeaw|=,HO_eGG9t<$v1;!Zrq9Y>^K|Q[9I4EZ,="au0@_'|zOCaV5EkU8<8NxNdQ*uMWyz4\AN<	+^m_J{WF!@rFvz,G@oFg|PV<Y%O\CQ2,Bjm&6j%9Sz,/ eik3l[&1j=C[L9Lnzh,T NYdFqYvMv'*M	+<K=+xW[;6P%O!Dk >2[;;t$@*A&4A<Yyiq2)7`+c/3I2_Mt7wI=a_vSc&4N"HkHzq][>D<
Ko=9$vBJrB#I6B_NV?P R6$Atp2w\Fk-^&?^`90z&I;]`4i{7FAU#({`wf;@*.Hiyg]<7i*yt;>X}H6/>b16@;U/z'u?j!?i,x')Ct
	9Nl>YG1tg(S`2yx!|!,,*~B2B;A3O:6o)722rb^QoXJbFZt~krmt+?*&:GTu<Yn3(y\O }Lqh~-SYY_ddxTUSpzDDRb&>
d/~y/vNy:>+C:	k'w40t,W3O35u_3%Ml%*Mm!RyEm`	YEf!?`.Opn5ro&*&cZfs=d\hw8O)1;[RvkS1"iWG_>{e
)EcBTK2`k[w|'##[#hi(U|y4cdpJ@=@oB,1j&6I'."ZnB,o(S\nqY(*n3CrB\y\9adr.Ty!u%s.-kJ"XO"Sv+[E)UX)dM}+sO)E2rp:F(B~he`:)WU^W9	]mBe8WQY'Sw9lq?'l,|cm)(yaKMCq=\d-:%-&YCE'1)[IudcFhb$Ty'nWw5yN%rx6fhM?)h/M3~~_=W:c=PwM*rf>khKO\C{g[\I[A
	-+q5ex=iqgj'SV>@NI8>Up5lPFIeT8C!XhSbju.4>N-D5B3D\5n9F3T$%`u6|eJI7B{\f?Y\Wap3uKpdWp?~H |%~?gctxVqd7|'5qR+vfFoZB UEDr[wO-070#Mtgapg _611_a-&)T;W
<B'Ne}kI5d2>u''!-5/Gi 0<*d!)JkI?l$ty,`j$m`uU)aXw='h^kmKu1zPc1
uK6vkR#q.`qh\K2%7S#?^6mcA{g![1dOZ@:	2MZX 5{`Z)/+ALe_Kx~!'L>wh5PKp.<: =#9`yUfW^B0%(jB\Dg\<uB4(O7tA
/:/Nc_:f7vKFBiW2}h.5 6c12,]]EsO::n74S#{*c7x
O,bvQ?\2M!OvGn"?{2XNfVeZ{_k5YrG<Obswp'
loG5y"aFH@/r1B#V!f+Qqj>w-g/R`dI#g.:5XwtegT]:V%Z-#~L.2.Mpv|l`Na&c*#x#$rbw&Rau8D(H,pPj?P@f^z
)Gg~qY)c]DuSWI7;D@@
lF2-BuCB+h?^m^AL!}7u[(/-QD+Ss,2\u=/Dw-~p9Cn<?O%8arGO##/9VpX1y7stS^7O'Tp$MM`&w\*74!q$#bYo3Zc5F~1[.N!/'t7n-r}"',Y!pHPuf.YWRk1=G#hFMFe?|p	-uF"bw(
h*^-kGYZ,5x#Ej<"(EVAXa9= skz[W2}dq2Knw9"hpfqGgF1$2\}AFr+	o?4;d 2;rx,/|N:C[_?DkF1FJRk`v'~n|[cluL(6TM	t;bV` !S{UOT76Xh[ZaJ/H&H6kk*h*$BhC
)I@J\h:br2
s[fv{w!x^r<<JD:(*.v=)Gm(B;6(O$%ule	oW9:IO|Fy3c'==foSG"a7\3 JWZ?m"hb|#9jqZpm
9v<k+'1APY\*I:nf'nJqR5*(]G<YPba;T!=X']/]"[3~7"Mx/92K{(b(B@>9?CkQuqxHA,_="VuA=hbLw7Pkf@
|f<P`%eO;%}
=57`~9S6L$o|M2y,,<dJ[8E=-1TZ> bLY2Z_?2\Ad%03ye?`'s"^UTfmKhEi#_I,xF\-~x;C:sB:=r
x$wjk
A)GP@ug m6G_x?fiiy#.Hms
@Lk[.ung<,)a;Zd<V}(fYdj$IsMjgM=gu;M|s+RHnVTjV#EReS@ x>"bgFh+FO[Bi,'7a3K.oY#7fPkH gw1Un!F!a/n"1I
6T%"fqpD: D?,o3LuMLmgr5H3[SDXo+J6{'dAD#w]xZ-hgwSLVDg;&G{68"i.&[y91RNU(p$2:8CZcGkH79sp:4-qyh
Uv^e]V=b>}imb((RXER~&t#J(mp4Gc+&G3TB$Ki"2],=@b#,[?LbfXA7>t}?O\uD.7,=Y~ojZ[4FO"*~2|<uv''Jj>mj
<NZUo|EFFpR(T;Ith\MU;U#4o5Zlit=N:WcMf7.U*?Us[)6~4IR4^B{!b$rc$PdRk :g#.~*s9k,43H_W$L4e]G#6e#	Wz;j(g,2yt{\0\}{4
s<>,c%EvZl*MVU7a@9d!;YE, Gd[}){NZ#9pNKkD+5dB> [z-U/7 T_Q1'Y:Jd-t/	ProGk'29$u5WuKX^YWt8mC6HN5Lh#c@n3	=mg%GwvNI|+/[[X'!mt\4Y{rZ.M	Q?G'/SI8A!T?"a'Y|7G6)Xo"q!;wHO_p9k3Yta}Z||G!BoW'h+M]":*)\l[ n"1n*}>rp/WUrEKtwB@ATa{y{>K%=+im%GOwsJa}[&@3zx0l	~+#}\b.?JAXE`S,g\NYx$>.{$&,.u	e{C]_1>0jnp|3TP|Q[4= 76j*_Pmg7 (-`734m~G<<An7xg)2FJWNxs h\[C$_%IX9^\%5g^B6z6I,+DiPIgUB2R0DHOA=~V3<m~K"[94iX	P/:<^g.f*D	{^f2|V}vwr.k<DGfUU2{,oV&GD:miD hCDk9x?AF!2PgM)}"jkI_h5Gb*dXy=V+tWBwqLer#a#l%ZOl:F0`2vGy5]Lp`A+"6=]29$,3k]9EOTi-nAIp:=	P#xw]HPG*&e7aW-fg"u_P+%D5QL
MktJH(C	O''8E.Dd*7>eO[S)S5SpmE,"/=N^>N	o%8RBecLhN8i)E(JC6VrKW7d29UsmXck!2hL3,E^5*F~MfgS:20BCSv%D'Uwa?g.WCErn-mQd4N_x=OTuGpt?S9[~e
F1ho+F3-R"CV!Ny= Jd~%k|;@uma1:QBW/5"iT\
SBXLd1mBo2h7cr8W|I %b&QY~'R_zn>A|\5UMRwMZ+7\'[d@g.0!Lw8<Aj@8W^uwY*3.[C0VEmb8pocy#0?;SZ0?S7]/U62vZBAlK`G)jg}<UD[KrsX7/1w
u"q
*13
o/p1bX>w@73@a"W;{?!+@\A}+a>-UnVM\_1[tz]uN^K,5I9+	X'i>4rz''8k`f"vAmf^_`u59@O3nzx ,w,uu%`G# ^vyy6OC&)B(46^X3sg h
`JhP}MU0	j(&j5yi(N yx;ST:.zv6y=)-
?-F!0HGb?gS:IZHsL`G>M,>\^Mapn&DCk22(<xQ'S3[jS2w3:E_@N**K4jc*t>x7hc,%\Z}SIhuM{[s{;Z%C{C-*%^]a>Gh[<~RYNQ|uJJ5?3'?sD|z:|HR+$]k,{1N
r@s<KuM>	'e)s"I~tb=UAx.5wwl|}ix68p>=eODDjgFVfT!:8UHlw-:QKC=>3!q0	Dg_]E%P}<4q&u/s?5W)"M6U8 S[#\FUJl%B|aIaBE0
E/3SQ vC:A&w-"0-x$dM>tQd.?BIYi7j)	
!O&?o~[	kIg2'ET%ZV5%=V\p?Gtw4a9gQ'8GH~8X+trE:~n:d^4Noc^Uf[\A?!=.1#t,)o.ym_7 9U,M/dX533]2CY{%CI)lbD;@2iP]H>#Ge(\}Ys& 9InZvN.6Xp1-X/YzXDs\tT9F@0Z4
x<Wh&rb3Q|\9uWdDONExZ1Ky$`i}k}Lwi<
>uS/tGB+!vR@iE:s|9`k98XG`3lr`^@>wKYcychg1Y/RJ{:U40-p8/6]MiMJ>"j[lxYe	,_ocJ-CiFnfk\Zy}1#JX`J'SORDO5\6b;Q$!97T!{m>"r/,26lIg;9b8>QX2\5.0goB$lT{_m+:fFUc{kHpT.2wIn/%t&TE^;yR)6!b=q%5HEIUNR{MH3R5P,Q~{)(@0\E`p9XW$07`3uKV:Af^vWG:5uv%fG0d@*dG[@J70"I&%mns2Q'<PJ7*>H;H`i4@iu30/6yl=i67sw*i}xMBEQ8Kl8|R0Tf.j6}\Rj{qz.&t36[2,CA.NuY?S81;XryQW1]da8PZ_}z]3k/co:n1l7Fg4C1z$!LI(pR{h~H+C@p7dR;E[RJrWv'>fC^K4w"vv&By^b[]R|-|BJLWdb6"#1`a,a~ENuv=oH8gj	N=_sYJ&);vbk^%W.G}cjE$2'/0}.Rh	" Fi
dEWL{Tn
933	~e$;1Plz5|90a4dqIuK=Nw\7iK4Taa)=:@!UV(6C^'H7UQz0p4^K?>4ZmUl6#*x#RP,NHiG.QG%$'Fe+rGvDjr=uS.d\~*
|Xqh,;,[xO`7M"t7I#_Ip]W~P9U14/!\;sUL[p@HgXdI:%zm{;0jC9a7f>-tj.u*;2;6b/&ej{pv\W1`ZQ0XUY!! Lg^T#F-uVk91^,3M^12u&2N9Y1)'sj]Rr2?(.;bFlM/;ZHt!(6-*
_sl{j9`O*c=)pUXIoD9F!q-*qYB%	sPn8>XE\Y,i7o*jO4K_UUo%!(P9m}V&y$:|[8?VL2	paC{7rU5/V('JIaH}c^Q|mMq),nb0Fze}3I^Do/pF_o~~(VAtF-5g,)%J9Fq(lfk[/:9fkC)Q -83=t`#g1T;cl'%RF>&HD/z0v	BJ:8OMVENl,5xB,%X.QKbEx5!rSZ~_KO!eFW	Gp9]tw[I9nD<}AKE	s>SP<B2v&iM<L>
:n]EXGfR&Q'"`j\|P.49~a\,M*VB}nv!G4M-B@JF+C<gizq_c(q.i!
d-+ip4A`Rj&~nLWTV{s8hQNn]PCu
}(b$[fu" RC2sq}l9^rx'w(G<ea14IRvH?f&x2q41/t_6gw9z-r>dvJ$8=9KjX3r n _'Ydc@9u0D1<Jqq'zE(XRc+>>{R}j<acD?Uwq-8gPVo,pl8 6RRbF4]'a"{Z
Ojw
 <'jM
U]!Q*Ro=%-)BQn)E.F`xVmU<MXkoQ6`hKBp'1[71hBM"|f=d8?n9Tb+$+F2=WIV_cgTRK3zW.}%g*/mOnNv{6>|Bw/<}.QyNbj.^^tcQrYhn_TRc9p+um|*jd	P\S%`|PR{kcL9h |S" s?!a!z(;qyf;WW7: ]aVE$4^>@.M5N`eoY6	aQquD09O,vf]E?1woaW=o>b!JMIY\.QK<DMJPQo^,V[j x(PfNf.'L6sk80L rrm8#&M@,f
eod^z/.)4j')Am'.W-	4Z{3k.12Q	;+Brq'I%!<#SxezMqd&;! v%5j^XP%dwo~C>EZynew#oF}X_"Wna;m"?5IwAhrx+,(	qeyawI1g3Gawwv86`3<u7I9/3h5V[	3;vvm6<lnK
ijUZY!HU)F[M%
S@rl+t>|l'3P4VpB48zg6wCod$=#U(mJ2(W++@x^M,QjRx;7V
eb"W|,#*M.)$j9%'!{V9U.*6mP)CI.LaU:IZ>=YgJ:jhdw9"TD9N#
nuh4vi$pWm~hxoA&rxV<DiDZh(LY'$HNp:&R&lK!bOC!%%3
"2D	ym"[^6l:t]'7@(l,v2]QH2JON\&KZ'
uRH~;a&&|E|/RtGJB<Ulx?L.7;sE^[uZ0TU6bN@rGG/)u4])	m?eHferMJj(i(#!#/	YXD;k\t|:.;\vc^,J:RmL{X2tja]SRKMw	/&	/M3$]v Qp9m^V;dUPH;~obOc\8dm2ufYZFF'd=P_rEO)}q4]vTKtRrROzY4H@fTXT'G4Q"#"a&YlTA|'rW0a.I(\aYJt;2r9``$s\Q1us1<&/OLg!dO20v98Y	2u{<dU]%)k`Z>< y:4Zfx'dolEjnJ?j1/c?stu"b:+lzM
qHl959nE"co"m%O=|Z0zip/}uuZgWQy@m	OzXB^R<zy39u&rVNM82EBp_$3K#3)$m}$myu#aPbMw(pd#f:Evk	E$>ojEy&WM.Ki)k5M9\1I/PyS]v
/\2	gxYZ0 ]+n
B4>`_1,AYI`H9Kk6*4OsnzzqW
o`P\X_)FB,2p@cS\yv@7HLzTX/~S$gfw]SyfI.1gZNaQ|6oh4h"k/o&4c]Agf[qLx8h]oX=%JIEo=V;`s7:IEkY;8FX3+_L\c(	v[fL/I~RvPC/%B@?t7<<M>;a0Q/5SJdQ+@RG<K$C!O5o ""U#Tvkv:kru"=kq;+pq'WG\n1el6hdI	I<y9
DZH"2u9w@O:yixmv	]0[|3d^ol=3J34BJ@G?-_R:!Yda2}	p^$ths)**j;!4$'<9<eS]<#4URH

U-n~nJe*8wH\S,=F\8|mX9W|B~+dSGE#LZ)>l(l^
n6Q\h8H<][R:_fvkPDqzA'
"L8=>h+CqYS"p6N>;8K,z<F3{\gVL;O'LI}qKwZHd/7lc[]3@,'A;e|w!;d*p^|u]tWr3H]2H`pFxb!POt-h%zE_w5H+PM4eVP^^[t:ixj\(</5Z4	CrtJ#IA4mT"6v9}?&GW3"1+HFgH\hz-lx0sCYB$='YuJc..KyS!VkUC<l:vU~sF}4@Nk}bQ04	)-4TJCrz%nP63cJ&k}}mTz*ddtKlH
A|:#lY($QF(FhhK @#}1qI	J]4IC0pxdDTvfG8EgB@UK)= Uz,F^8Nx$ap(x85zpYX6(la(-L^JA2RZ:[. Kx|8pRFr~Q'H"=U_H6"GyXx3Ng%&c4x%1J}p]0\+bqzE$0"@wGHk]J/)k:Pq4g:W]GeU%QIdQ%n6	V&_O<r%-64M=;?+$LDFV,aMc~ax<B@3c6j*3KSb6Z]Y=M.W'f(6Y]Ru]hR!B,zui</H"v;I'A
1S}oIU&cd0kVikR;}):hp5+'n7U.`<RWKW*IVyHz!`q%KP4:L3#c=,-`5s5L"}@OD|{Ta5.YyBueq*K^wGiroO&|/ojcHGRIdl@.
uN_V,VKV./165/K@e&f]dC'jgr4mNqT;:;,
},hRr!N-">iR,H+8)TCH7nAo>2Zz<s=$qc.4&23Py{Ia%:A;{I#+:'	i%.lc0fwm>av|[AU:NLOQ?g&w)J80'/uHj'yyi Vhil-ZoU-z-o$OEipL_cLLi6af!z(]S[vBr2wg1x*uJkalkiz4fisJ4 ~`[Jn7^n*8oiGUbgnCH)6<nQ$Abosiwy"m0AYy;h$Xa(XvgUbAu3~N/OAF J"KK"<0Ad@4:CJq?_yc=l$W3$sNbG2s
R
)u0)H_SoqP^e*B
$URk{DfQ8UQX<v'zf~TDDurYK']&M=d%u{`:ySP?!+8TfN!PXUz4gC\x`"U_pxq2KA6Y*4%-Y@W+QoYZEUkU;`XC10u4U	?iwJrm-g^5!s(6BMw,6S\!2u"x-Vfv1m+quix!d/);g)B1.aqCO1"|y<H4$qq\vq$2]wg3wkn0}@"6"|$2	aaR?p!]Z!p:eGV8h|y>"Y'smTrueJ,h!K@*k(zoX,B!6E6	WP+eke#Oa`m1![w\<6k-Mr=cu8`Lsf03NxuvWS1)OTS!C3J4OC"`\Gnc)>|KO)CT#s0ox0L+V$2P|pJ~75&nm&c%7+[MYDJo(tI\Bd7?<4o@sK'
~8^::Vj*/`qP!^0"7i%coMSK:#*d1L%GQR0<Q@ew2'&b;|dA`<jC2i5+h(G1)h<5g=gP0u&'*1)V4x@TuUXTSe{xMxr(u[!2R)TQDT:pE4%-BiL=vgWI@Zg@z\]6 xXBA"&F)nw7~-/bGTuqFO]jFM|";KKx:\Vbu|C+BTm&ZR@Z-}cB#(Zjv%(ew+B1 ED3i!hS !?=G<jsY,~	T<Cn-oz=%](/IE8gTr|WrI![)IbC-J>+|jvV:\yL$h]$j_;dGA&I&X9Qn$^CU!3(J)tWyRY}:h8|yf3t[HU`9~"2q8.^ |R;N>^V%\!^$)%>"&m
22o<?%\f+En9QEvL)nrK2;g0G/)9,CgFZ}{;<[Ux!L6$@1z	^6Y<ZR]rc/CI"/00}^#*	H\KW2Bfs'Fytz9>VNAjPG1G/Ez;Ylx63!oA#:w+RH"%Ao}tMQ7A#$[nr+C}c"MU/R}%?y&Z#gxhcPck^~<	{~Og$J4D'_g	"]_3W$("7Kt:nxa]N@aUKi)T"2Y</7Foo9EmJRIpA5J[H
G</ym-AQruG[Fk[.@."R&	Y`JO-L6~?z^|,{\.mk#XSFV#CeUVol\Md[7#c)[?]1{UM|)"Wzp676L_Q2r#X2 pf6\EPnJA(@-gmG^z,`I{^%vUdR7gaP(	6U4llz';4n\=Mn8G:B=Q8D viNM;UJSFKn&W,]nj{(SeDdiVFGg%YJS!6OTuNSt*3os'uJey$B1
_;wYZhZ,1<}=>TdaX4GqG)v-ArE)L<vG/)Q!IIEMG$V8.f-dVaR1oX@7rGly1*90;6hvzdsx8*xpI.Ykr0R'"+vQdo`_wM$1fL|`Md@1^D4W@cBO{pP<0DE}I3f0ta""?gsv};K~WQ[4nM<\86?H^Tb]%]P}4rI`8shVURHoGoX3(%zQ|[gn84.{T0~cp=U?nI)`K7yI:Oka[->OZgU;]6|SD9(Z!A?%v"%%"`ebRU(>s1xuU>juY&)l#;Z(E4qR/GcKke90	OYB	(=M4529-6buh1rN]&T\zysj!I`BKa'I`|k%JE~L#hUQZH)h1[de`	1G-74}vN$Rb'6#fVHgsX-:}U;+`e[` w9il-t->o0R"(OuX/u'NOx3+a+aD'xe_=g0
"CK2H<XyqVIn:x?Wd"hy3MB(:6mr][GR.`Ob[B#Nu=CYX&D|uHTzbCwbumwRVZsQQ*"HcbG:)ImKIba,(mW/_6pWe{-n-(0>3^zO:3 Jgb-s}5T@I];_g0.HDsr.m:zv5niMfHVqSVc9fw8.^GZ*?>j5dyYgHIkIRglv;zT;,$zm@*X,RD?R'#-ATN`EY'Y	Lv~o'ky77E]xeM"zTW[O?by+ncP8:3%|	;V,":9Gr?GZVNTSc|*bI=3=:j-NhrvUV*@,7YYEA8=eeeXRH&cJ+uAjAjD#u"q<#v3_^ee^L#K)}-3SL)60C,v"bA`c6j`5<0LoKI~?}s0KjI
B_U@ rvLpl=	$<2.y$W0]v	7%|
U:U:Hg%D.&;=NwmqWv gyG[[_l2&uGbdr1
:?
:*8AwpYXXXy	Z,\ aaq*WfZ+Qf.ym.?V6p%P;'Q=pr>8O h7{K!?}=prrUrr=}0_?gQ V|'4xuaQ9MvDn%#4+Hap15@SDsuoO
i'Q6>eNe	Vv{T;UoH3x<_x{.Xetb<aY<_rt4hL{?>0yseI>r1iJDI0W-	a1`Z$]2jlvUIj),	N[GeZ[bq`EBKz< 0cEb-@bL
}Qg(ZZug)4ML
o0-s+GWaXW3Z1nqUcZ#G]xbjbDs:%Y=ooTDl^T6,m[8C5I6MMYlN~5*@,OZwLw^]KeY{fS
[1EaPG:Gp`YP:LfbNwi	7K*TO&S-*]MUu/idyPsvz}>OWN+1D	-v	i1G;W/@!?lZ8dBkW=}4SSx[	IP5?QiCz>V\<2w{$T|4*R%J;Bjd\Ee9.Hkl"ON Rm{h[|j^UO"?:?dYs2zF!9l\TK]|]WL=1}';+ .r#0~gAKUFE)KV	"#J
&uk!reF%(#i(9Mf>'bPiY-1X&.AZ]Rfs.s%xy:HUI"u?> #sskz%VQlU0+3}6xD(Bgq__"#I^sXUT6$GPaiAW12X	O<Q}BF,(-+#NTX'0+e:R_O*DBN@.9FP5:*Ovtpy,Vq`=WCv&$adkr^Di%qsA~^Bj>%p#L12?kVe!>JL.tEx^z7H)Fzd_|Hv&|jGJrMH$et!oXKlzSQD~JTK5)Z<ZIa/!hv'kgq=y}r>X>dS[>?RJ}Kw 1hxI=Q7P).,RP5|Y(<}"j`;O Pxg\$ng.f-uP~Kk$U,+ot+HE$g'I
r6C
/4eIXD
:	MNu\{G+xLr.@F[DQ9Zx-VqOnMAX!a@v'Wv[O6vX|x:G*5_lA1nDpS[M&s%"r_8)e9=hI|{#-8AD=h"pv=g`vv,G5ut0CueUEi*P?od37ny@J[uy]<K`AE>60HhfNS1^E7!+Rro6U7_T+mU(0vhuI8xZwo\`w;7Tc<%T,^l%uVVNpXe,4rTRnIr6f0Z1'WW\zbq@4>I
GTV8	!l"jzt_`o\,8q]KB!Z'^."	^zIXDFI!i05K\T#&_st<6	=k\KJ$\ow}lTFkL.oCuH?]Fl+Yx=u~{EK3 ":QD|zetVzIa\96Nc71r1%xmJR;F{Mb5eqA$NM.!SI@Bmm_;""E"+:?}896Gr,PO3f_#v9u3kE]4hmI~LwdYNRR.\dd=9]-Ro_uu",j6qD\w&MHxV*mg'NxKAKn{mriA#Fth)X**D(f&#,7PToeV+)fG*S#tM7?l1f3}h]MY+"j_{PeP/b7piLC#bT\sJyZR*[$BbkG4.Yx}</q;h
UG6>PgeCk Z_x,VsY=v`BeTi WGjT", #.Qo/cDg|1Qqmtnv<~fW)Eycn@21PzB>|"_vpS<@]2#LG_,#
wr"N^Qgs}?#<w;:FO[JujQI1^;gS4uXh_0R#Iq~5Ur'|Q=TssPM>~O *'
PB]tqO<fiRt&#bDfh-L;D`JIjxy2]gFOm_\`3cNf$3a>iwP-Vm*s:[On(rLyY@pxEr'c~R9/_@u<*(H=au;;N<R5{bkAN;,41F7X oFcv}PtDD&#k2..`leya"F*w*rD"s`"PA*ug&QSVXi!{I1W#p^k	dh-mnOkn--vGI-@|OrQ{yXw|F6H}!aDx uubH,yT6[-7uYHW$KGJkt#Dv'zX^*'Y^P(}:\]l_V	0-q2:hL k`VYq[@[3E,>=L_L{xWGAEx3	7`O.>FJK<77q&*!<E)+o2pu>AiUAw/\m<lz+1]z)uW|0Hi>\3(F`BkTmq.@]jGGy/Eq0{nhz!_OTuy4Pi&G/3ZZ.>w#zo>]h2dp .-,9P%CmAV^wt^j?{&G)_Ftw@"5W~c2/LF_)#2Tm9NS}Vo3[a%^L-!8#{_]i6>+6{w^k09:VA=\*ucIqG#0^q~1nHSpl{_wD^Xk?WrS+K2_x#g/#UKKM=LwNb{;h&)%5aEWR94S
RNMS88&(h:yCg;duPxi	1jTW"x"a{`<o/B-7\\u0Wk>lX"d_06)U7RFTba#+{Xw"b}%Wc?.;vjg"iWZFrdfHbqPhVbf{T)Zg%tDUhw]~~2uEsmnxAn-FXO70;D3l6.[Nmq3 @-~HcbW9O
vVT:M
v&~rLPlqs|Eqs?RVA6Z%cma?ULQ5TkuE`.CehijuPwDQ&e6/K{|=+{ea:mW SeM~l77162B3$QU]D#OW;S`V
%:8)Kd7)u3!zu<(Upm<k)TXaX7C#VJQ'E@6L%'PL=v"?~;d	<Q9|y	gh0i|g92oiF6vf~#qhW%o7YY^Enw>Z-4+</kN?A]-dcw}o	/jn._Tuq*_"T3Y7nsk<2j$bD}+P0(Y=.}CzZ}EX-DVd2=m19Zsx@jC"aK%DX|t)A9}Ud.w&wm!h]/r`tTN?'9RxTv9y>d(bSo~r ?o>>^~bVBu^[kWc<xl ]tg6g|Ay=,.9Yhqlo};eB=2
KEdl3
!|1J>~OVg<O]t5;NA7]-Kh<hn]D2H-u"F84f@S:FBvI{7mJtV=VI+XrLYm\K9v@xNxHw'Z'}t35wxgi&e*^/oW$]myv!q7PlK+Q.1D5*7T1<eY&[{L(/<eJf|ui!aXv|_x$~p95|e9wV@[,('(^2"H
/g4s=<R0"=@M?Y3{@ITC[2Hmq4[nI9]l-`K?vvo`>qNRHO-4Dp"=(?>/]9Ch4uCCevU]/BM=#j4[FI9[ey0V?9&	tm$z/^H&`,Pe5CEc.G[[Xd4f,xfcUWbMXf[5]
h19ULyH[#K%wr+jiK(s-4wtbL_:	w_gpEB83U<wNYR()_/P')"tl[7+Z3wh\+Fysuts)e^N<$We	6PLBtW&u=Gq)4TJuV1Rnp.*/.C|Vj]:hBxQEzQ[yo4;p;:x$[HPi"Omhd\] r4r\,b_EX]eJz\H]T~b?JLU.r_` AGa-fr2G>7*>`M"8G #Ry}OSaBEoPQp)jKuvR:/Xe6qS1o{"ssB@v"q^=tQ"mxlm%s\-#ba$@7UWZ:WV>yuS&{z	eXz#H-jJtJY30h@]f-G=G Dtr	w5?t)QwK, ML-UU"+_5QL?/^j5g0~<jAoxGF"N9$lyl<mFOu@XrBy6"#F+D}jY){"*"gU?%A2^T|dlk./aB+ZKQ8*~TiT2^8V8B=L7+f\ysSu%2j`
f	R*w1}5H=VczGl|~mk?ATB/\j:KE_GmNywty|A;=!9#T'loLf$O+?EHH3%BQK4tR^$#(luT,D5nP0F~:{>	5Q%x%]a%*"e"h+KFC$9^mn'DiT)-)Dh7G09RKW{?2I&[k"7-e\I;K=\)8L`k'6k9= yH8< t+.e|0-KQFsF,BtAGRcg%2fL3f[aZH5'=dGBI_</3}8icAmy7*\_S}i=0[jIr5Vq8;;Ug sim;*ma D/8we7imv V/MVqk?JPu[2Xfr0xE:tA^So\O.4px	z" lZhK({@6.z;9V!lU23Xy+x	.war]Vwwq}8I_-sf)``{hu}^VkEP%h5ux\<wp6:uw]^U{`$ +HJ_hT,BfPzW7` 6-p-j@33vdA>m<*x4IV{h$}~wC2U<K2''fqyb;}A!?]!6mKnS_F/N(F7{q'!-61|'#OmK2O pZ!2Xv?}~f|-nzluTdSm$D2e@a
C MED?peW9i[Y>PNZV,s!N6|,Xz\;)05^G)+!OoU)SaLGr=9@=:lR-L]ZkEG.p;kIaD~4hnz_{(ebO2=GsEjAc#Dw2d|*Lvqku^l,nB$P9\l`vLjc2d4rk$\
*zaNJvq&ykSdhTIR{.eHpd/j`o	/nB!qB>QS&SxfuOyzd,X)C>
g^l;>7l`
X,wxd]@8)'Z'roIeZtFBE2xp!?Tc]=d%hT2y*b4Z!{fZ&O_|1LtD`o#b\wlv?VNhz,ur"`:Boi|nKHh49( ';3uch&Ac0Nu(.X)15~W2lq]*\s80LaM61}?&g#p''"N.j)ZqER%TE!KVj4&py}\o!O<%(D
j.tGrFMcY2!qL60Ks|`S"p<<pWZX&im]	iy4e]b$OXxvC#0S?}@%)e%@cZ>ck4{TWyQ
k%wMESi!"R*LI,ezOCWBfQj}_'{(J?+jJkhRV^!ZKWkhDsu3l:c-vHhKj{uhy!5(_m6='Rv0=D]$5A-bTiH)t\M.%9@W[vSMT*9)`1<*o^;%B_,Hf4\6Wp6>'Mnfq:4f?O5JxI-)f+t(j3.J>}'XlgR]2_LccUkox;9<>^}3C]StbF,;>l98JzM+Z9&C_37+U<4'xJDs@_1+&sJZVke`GTF$dC}X=|tFI"[	<_rzJBm,8z#d;}X|#Z,)Hf/+D4TFq6<b*00KK!3 phI?By	LQn2@5_G{w=2+UO"[aQKoV0M[SHE%:W%C4Z"200Q1umQx>8c!CdooTtV*rzw*ExPnr>/|&f}[Zx*FZ+=oO?XrNc3tNrs0lN1%)_WLCfuB7"R]+<>#
lS!<#$Iyy16]<(^=vvT^	Q2<i1 a|HX$VqGu}]I3T=l!j|.`Mq"y(
kC|EoMzfYc
UU,B4"xeA3\gfR0?NUP_~.+5l0L7X	XP?=br3r=YU^oe<H>]YLtuUl&J4])sts6Xx4}IQ0tYAAg	l.RqS`M#P4r2f8+wkXM(`,<G"=XtD4gq*_N-0LWqN|~/pVy%Kj
x 9$T"tymvw=+s~nDH)\;k[vsK7@AUX:~Z{].;d`>pWx|Nm3K
?]/J^7~=?3Eosp<cx{Hjf	qWl}bZ_O/xrc32%zZ'zQrrt8(dNR\'!c^!Y30s]@0o;."sC<'J?rbvP6<2.w_%U:&$lUR/53;\T IUCfZF (NQ*OG
&FrMLnj#hUs_0iF9"{5(yIx8PzGZwywNHQBoObfIa|HqV^_jr.xnw"zBBu&P[/v*GP<pG]1$ 4Y=mV3ay+fD5uuO-[Hn6~K` 3B.Erj4d$~m4Xd
9&(KL/@N|cKXqhrwWJ$I,w}wJOeH
L-+E	FcWen=s&6z1hIv{J [Gztn%[^L"gz)o/Bhq%8n"EImFm.uiD$	;/6"RlDe;
y@mZn1X[]0n>t;."xrDW	%F@j][8^tI5)iHH@;4P%d@`{H@|(50U|l`6FC[&8_9BE8i>+}qfxlC@um"a^tM:>}K"%j>>*GzJhP#X +rW5	4vKqkG`K:.|lf&*fH5S;UDR+%l
tp_-P<HD/k^gvkg4vhy}kHPv$eZ,Old$39vh5BT,W/^X8;@@CSded.H314J2*%i#PDlrED#=zxGc$GO"_{P~+p<-rj"aXlJ1&C)cP&q$7oE#fj:|>^qQemV&E0"di&{5z]B!%&8#vbnt4_u6n55WWEXT+	,5$jW#s5[eoG,JzOn$KtG
xkELbHOnSB=h%H(^By;4\^JWmR& <:H5~1zSH3]:_kzAqbphbsH,;hIHeN:6r?!,{lV6*f#j^H,t('P|P+DA6Mjb#Hv5=	6o#LMl=8xNUSn~yl/FRQRqrJ#h?g(vTjk &c[j!2X==e(g;Kc`Z'p?Q:xGi\eC'OPIHXk'4 8GEc~=6-.rHJOW4WEacP+xT/4Jiz5kCRsCp\(L2F	8]I6AU;]9l[ ^_J5<4efE8ccp0^xo,*2^>(8X*	A}<0^~X?gA%	cW{D0WBe;36tz]9e`32[.f[L80b-4aK'4pQ-Pq2M+2\~-a)<
]J^[C/F|m`eA3w;5!2rjx^#5cxlyPs-k`9TXNbk 0%OERR|X#E*itFs/)m@KK	Pllu`>DoFx,L)=a{le*J(1~_W\YD}\	Tr6_h#vU~/B+L(fN5XC1c6]!@/`
&XilZtZ\}.z>]=caQ4|O.U\U{-e%S5C?6rmLcSXD<5">YmeF4J@&	U:YgWK/dR,_8IY_|E9d[b<\dzHEE;/gUk<]8j V/scZ_i_O;lL8{iw]ux00TR4#De3Wfy;*m[\{bm.Na4:		-I?~>X,*-PL3)FI!Can#w\, g@^7b[1&dv`maw&C"%@twcB:x0,*V9xr}P54C!:rFiT_mPk>qFhC81uXbao9xJ;39$l3pd\kNKpz>aD%uSyph^UE%mgs1%N.W=VrAZ*)QGI!L1^}Ayw?Gun7}hELcG4K(*HZ/=!G'%v_I=iRS!kmWf{m]"1G=ys6H{fGhrpib5?T>.wf=AoG&|S.85_uY
7_*`ffe[LuKgZo%~!\![Yn#S'S{su#G/Mz}B(Ckdaqt3R5G~j,sLg7%jVQLo0Bes`vu9>Kb4LM }xdb`YXMW03}+?56zE$hZm@-@@F$<Z<J/LkI:
Sr6.C*}BI
(<om*3 IO	jzM.Nti=bq!}|!u,xS("
\hFd-:@pCx+e.w<?J_*g3Iln.K3_6q4(K(kmE@MVNYMEos'UPT":PPXH[	7|C5SL5]$Z[N8WT0+7(]@pb-
KbA4g"En\PP*~oK17LKA{qx6H,haMx\:0LCNv%sRwc\!IA nOR>&&e1eCLkbI?&)%gj{.UcuLv^o9PAP5,ez"S]<Vm_&-c~zAp fb*rfXN;(lk2;X?-@MNN*4OrJ*"T@/X*+2jj`'=d6=.uim|p0YkVq"w4	)7t?xu$l[x%MjkiZm~Bv"dUDyEIZp`LQ;WQ,1BWvrw2gm;Ifcl@=QxoGc,isf ^u.m{a0mj
@}_&1r`gKs7<,9=;v-/mdxko#MqolO0zHZM\'r(00vp0*1zW<mH5	>B^j"v}R;cutl&A]j'H};y#}7}au`T)*s%Nou1Hn(+.y{@fKsIG`X{<#3)V{)_l9&S3rIN\~G%tlTHGY7	UW0u97;<YU%"h%<J}(LNlO!i8L2*)IMtR&>kW\nmzTG)C*,mRfB&_ub}D&
LT-vL*2|la6%[&wVtfo%.)-lG&PoQNsIjch']%1ad!t}5pW]L$I!es}PFfh8_BiJ7S*,%u*1)mn7nhmP +syrtuL
z|uwk+[@@-&A\&)RHc(t#o #wGcX_a^a7e=p"`b,E[0u$`!)/Nh5aw:Yn`0`/p$JRT>e='~o(l;r1	s3o-`w{p:e`[UsiBC6TY9?+:daNR9|##?MLCXxb
8B?Q9D~)jL*,{K|cM,-(Ij-Ij,D,Rzf#c Z@pMr.O[V,|rUqcyxL#c5'`!UUe|3d!5%AF5l8-JGP>,"'bL35O&Yu(8vQ0?}),(W	cS"kq|2AbV\%`&IAB*IiTDVk!o%6O]A=d8*VP7DGO"~;~:M&evOx;&8N^qEt,xIlQA\$`=rV'gzb>6_66Yj%_c:v_DyMCW:lS}v
@4\_\\`6M-iQB
"BzNlwoLt{&<DDo=Nj1rm2MsawWppgg":|m="'0.*.0GklCq`B~'K4P"Kmk;~y7"hS_L^c~#!)5Z]lt-:z{d0,/4lWU];UmP^K`-(IMDpz&^ol7sv8#vLQ}@
!{;pc-uSsX{Cm&E*Z&Rk" }1MykJ. {WpQPW<kZK8<#	1as: sEy'mW%Q)L|_]^Nys;9li\lX;6:LEz;G-](p-cQ2F$,Y>5aKGE%[w9271"L(xwM]^d={P=Mu(Yi<T$oY6'GcX8-$V!%5?5	4Vm&}!"H#QiyP\@n@gi2GrNatel'^u#@JIF)Sydx&[#s	8	/c~&bwK;j@L;tg 'MvzXIvY}uFq+[q"k(n%b7SM|}g$7S&ohU.Q?g$@+Qj?Z>;pD:9}.(f$A,[+z*e2|KKKi+*v_yN_GYw2Ve{WiHUJI(|RK.	wKic"n}q^u:uMp9[pU&#~N+F"u8z-[C|Mz[-#RTvc[2*vzPVWBl{$|?)E	H@96~Elv$ki\&}n`qi2C:Zw@"=9f;~N2c'
@_h\A e'r,1 {P_;#!#m`0(|,gAaT[aqGbj?YV{@DVaQo(B1coU[ {0!GAJw[b6K`5=?V8x ~2{kzhU*Nxkb,[#Wbd&>RMczb+.]ruy8SI{-n3:FnHu^){9X`,,g<_D;DIL{o<l^T=E@!u
'~Ya])!gQ[0:oo7(1)o=y*8%r-r2qm|:14VY1.P_,:g4o/]`Np(cFYi?B9&XnFt&cA]<3EXQkG\=mGmv!B*|iyKHt4OnCZ6I[@|(]ej(d/=qm?Xt[1&y^zB[@W+n~#N0^V0=2]Tx@7]&PV&mV2Q]WoIuW9N.r[*iD{cVo#1>xs&VpRs,\qHbm[b<w[)3aw`$_?;V{y1&)Ru3d}D&Dhfd5A3ux~bYd^yd"1Dw}o,)1qj:x
NiK3}q?gk|@'
)hJ)CRZFN12l]mD57$*an$Aoor-B9n15H:?p-#%nN()&n2`c-1O6w;FKHC,DnANe[2RJe%Y
\eUUlF^;XHI]inIeG47IzhO: >z!CH]OU!5l/zJLXKPsZl[+:~*;&x:)=Y;+sapS%S&EDq`'f(!tOJ<	Qo
T=iWa[T7x:hUjz^:Aj;<](c&7&A)3YI[@(rrn |\":5h^uQ!}r-QuK_	UEPz:P}el>@URyYyI,5~UQYby~{f}s|NpyH]q4XvK]#t
CXf.ObSO7\+IO{SU@D2nqkz0lBIup 5$h[=CAgsbyaaGTb6&[Q>GvGwmBZpUZ}h=-@5.%j6V^f;V%1Pw{_-m1D;4543|S\%P)q,qX	k@G8OS%+xu?WT]OwH??%T^<e!WItxt7?d@9C_%u9t4X0Cl)'Y"D,4b(Cg;?-Fg<v-6e>	ndb7)v3fK'Li*4\I%yKvn_XmN6"B?(f`xS/2Jo<P2)&(qum[_Mlg]%wz9LS%0O"$Gza7IV[$=oqD1W+Woepnnq%Qv)";rIEJeQojLV5yxUe!++pz;>A$J |{P"(Kv_igI9^`/aCgXg|LV{=:G5wIlt}5+;aul_mYDx;#1y(Z9L=/r?b:QTnr\YvYBcVf'3jt\Hv#`xGU0HpX=t|nR(1f.hGPz~:B9pF@	5RcO}&RL`O%_?jSt~ps9G\+:I?;vD"$gp*^.()f
(-j}HXS!F_.v@m#;Sa%L(:gN;*'AKm'Vif+~O`\*!M#'lCYu20ISCOEkfUbKq\OeTF|+O#RchgftC^r^i|=Mf9TSViA.bUQ|mO<=b_]ZuVP87@KDS[0*!182"+GFg)Zvo+9[0O5XNe7jLRnh9jh<to:,fFEtBHBjMceIP4;Sj?DD&3{u6hwm/e~0<XY-hL^:Xv
MW'/Bjsl}(5,_`;GN~B	/@v'8c5LS^GyRr}8JE5-=!g0O~l-#xyT~YonZ~f@HZ 0}89Oz<-~^tj,j,$pB%:I4atlFe9Pp4)[Q"5bK'B_o_#WA8p"OJNWM^n`&Hti/OW/ZvZHWOq1Y8e	Xh_G	GcxQ_L+%T#E%+i^ZV/B$=h,A$^63>tKaf|6i:)0H]}%hZ@=jriq$"sT~*^pU5De?z"Ate7cfQgr8teS9t&q%%W(ozj bC|_l8B)>^Scr}sL6aN?]{B8XJgd^W\xza=#xFqt&;/hN[85Zj+f^"[\ify6n>s&aQ&w'o>1TII4Lzww'b$ZJK'gC|5z,YH2<F&d=^:VYfu$Jm{V?s2$@CjLH<==N7 ,a%o+LF>+N'L,c,oTgqv1E;"&,	2*Qt{}'SQ1ZC1Fpin8$K',E78#5wtus>DEgxGt0%?U/pnF%;/OMP;yZEbl#w?#UjKea&\E8#fDw$fZ_A*D@IU0BLqwY'~#0E#V+ jKsa6"Elo4bP8Q
v|`E+M8	aj#<4MUSt+fk$cwt.DYER@Pk7Ui;90[5 BF3Q~4;/5	;vd."?`~&$bjTn1aQL}z=(%4(>6!;1n1(i[0,%vA 3.D%IBa1{sgW72H8Fc"g.G.wm<wH)6wm*d' CG@ri_I&Ei?QSN&1W%)w_'"[;f*Nx\)8K37"o>`)Q5}|po8EQN>\(G m9=Lex]TEY.Qi[yzU#_ttE"$`fPF\U6nn_[\eXo,6h	x)DI-b\,vfv^jZ]xm,b|s=h:#,`H)zD!aASooL;pC#+QUrTtZ1\ZY`7Rv?wbJn= r:=:noT0bFd|A,|1X^BFqJC,:urNRi[ZWd#HXvf132O~&C!r"Me&Aty+fgsqd>->$P/ K3'{eo>|_|Mp(3$}3J>FmJ@uZo>d!6sx#|Y%x*r>%B.b(/Sv<uPZ.H[:yc|Z`c/0k
8rD-lTm=X@)]\%8wr>X,'BMy"D;!xCm*1udeD_K$y{M}cc*NO0,ztD!@@2 $J8iF^#
:R\`!
~(6Ge[	kjrF8L\ ag8muxSE%Bh0ThGE+o{)}A4c`k)D(
:E;Y"6`"$~O#0h9uC1{"C0Hai?vf m#0q
ycA""@PVUD]QgiP&"mYxHj-V]Y=F+I=^Jq1#!?%	BR</b7uE]BK'@+dR0OP|]e!g1'JU~/|96wid`-`"YIb1,*|QS/D`c
/P6cg\HC&b.:zLM!"e\Y6dfE&|vOqW>x>Q[omj|MASjepqv~ZtVHnC.0Gjr+`rV&pB$r]q2"B,Q|3 ?L2qH?v	Q\_[gd5\:oRLd;#jtk{e1(To6A/1I1s!JgD?QEi6E{{EgMX|V/Tf#fTdR1DjcBA2@yx,8]^2qa4yC9!PL7+\eL"&`@8yxt,=plGy162hrb~ot~S	frlbZkMsb?J/vaVmVMwHeF	vtBX,4uZxLJh_w::"bj##kkm,(m{zQvOM{`V#Hcd/r>"1j=/'S!6O}qBw.aoSKLwGaZ+}I 4s}-Y`Jq6u&-l59w$PHJ-xJ<pS8Y;QuxgD=0cyS$>I0IXZ'h4g^[F0KD(^,^!jNxCwc'"s}T&Y]~56Z
2(D=S6[J#Qi`<U5"{%uuTTnN9P4	LkE stTd$5(]yx&3F?B,Kr(1k>1Q5NCWPA<A:r6S{RW ]>5\J\`F^Ii(=nZl0mRVcWG@r4ROy,7Q6By3YA|os@w9L0JKd-zCKnwT	Y5,7Mf^Wh4MT%5>$tS;,m?MA2f:hhV3zkq|aRotm=u3pn,y8It];QL4u29!ZOSwN]Oj6NpC53H?Nw8;I"
FQ=prs8_xVN`(iQY$Q(.zPuaJvkTodN) io(|dqbZ;zKul]l{MN,oAIw.<VyT/.A^.xv#ay2weNOTE!-y!([wVTHqB/YR!PQk;wqF3d^'$`I{V`V(J\k"HT?.u\d1%Jev{i5Nb1:JVG7O0HP=3k60+Z3PD(xSUkvZ#qT( #T`#Z#x6bf1jjPc
cRxE}3{)QW=ujsXUHB\=O)m"BV1%qij^v:	OOG?^C%55ad\g	Y)u(NsnXS4lR!g^Rp[dRi+
uZ}8u=s!R$M|"*	@2XI5faTi/6HtQzqN=[aSTi/~+ch8d4=#b
3"^}i4-pk%Kan;vEA]<DPs8W?IXM|>Ih{y7nhGx,Pln8B (vM_\n{?	c@d%}r'@T<ve*]4`ueb.;~[c@1$/`<k
aII\X#
-M>6mw".zZm[SGB0$B=8"__vZ1>^tD/P55canVw[67VIZyZ|0NYhgI20[l)	75.iogALe]|]7sX)*eq5iKrQy _#F=/g.\!CJ;^.;\'~1#:S#qtF_P"VDp')l]D54gB\ kihBW.LssUH+z.1O=q[\Sz{e6s):Tpm6k9^X2DXz@5ea2,#U	a*u(r'zS&,{JP:j./	}za.plR-Jx%?Yb#<KZ'P+G]1=Wgvb@Q}o'+`LGzH'F=2BHIza3h<>48I@K 92Wm|\|WXO2B<}	|M!D?8R,5QuPZd|\$~c^r_[ujS-h>MN`(cc2G+oEqA._>#48W>tUM6\aw+?	&x!jU1xWnd30RwFmn>P~nd-T-8R:vTr,K@1tO_2HFUL.+t9dJ4Q Hdv!T6;]4pj:?hPPUsJPrBG8z	V_'WmEu/bu71Bs2JoEOY0w@g%'l+l7P^l2<`F1>ksK*Q^ =Ism`Dl
7#b0Q+rgxg^Ea P!}a03djeSoZwjZKc5S*>$$i\n,.(8/t4a'd\o\a+z((+#&xGk,lL,	Fc+D)CF;JL4%}TgE~M$7@,.AF.bso	=PZc7N
asp7a	X:2$H9j*NG<Q?kciV&c\WGTl*\p=*~%qLS*p&}c$?sM.kJKr:FZ]pbZ*!D!1&Xa\~xW"+>wsn6"Z.[(b:4")@
itmddeB@So i%Hd!`jZBd-FzilX>s56K5`_i{T=r+5iT>,Ih@K+A
HRm:@NoA11;k%#;GH4bKE[[xG(~sdc@F47O'fOKBY;Z#{qk*bvgH
O{{/2Dm4_ZX#0l?'K)	4)"{>c:-0y:{b7;)`d	O8G`XK='% :}e!Z_S'_
"G'z6W0*Mn)A'^2~!A+
>`J)u0%f<{]Rsfe}lMW-l='Hp\Fv0	{deMal+@wFD|u$fNw\3&(E~LY=nZd=5<9hCn<|/fihBI,aZj~M<vjnaBE84)	>UYn6o!QxWL_})^o%n1nG`nP	7Y7ExE!m08c}Zi(lQ%>'S+;|WUo[;	lH^X0/.y6\E!n49Vu1@"L&1Hy?
V<8m:%-`Qy>0$\U*u7!bR*0K|xR964ep=	m|6MQDwhUuXoYEGT)bF-|i'^"&,;|$4:i6xFn'`M'<\ld	\PgS53	j%:27R	0J>bje9$e!A`z4l1|6K[CU[k7VndF~b0^G.O:Ny|v<c	<;s9cKg5*uRl(PT 2qAu@,4
:w>0${{6_3Su~H
s9LdMaQ:yLrmng`<gQ_$v}<E82A,kv\(El*gOF/Z7l)>TgBa	_z!?(WY$KhBhTZKo q9&}bGWV0Phhg~t9HKJG_"aU=%X!bx ;|cO}Pm0qfeEZBJDukp-iFOr@Kb|h&rx12D[H""X]q+G/d-G[Q@7"?I>[g3CjmPmtP91@	]q=AXR8PA@%ro[-n(o$m(*0f67mN];5KjIFFO1XuB\PTGypgR&z?@En\.jF>8VbTy6.!d5nh.~+9PJ~lW.BM+-|))c2zqL7#:d`><2e,^w!#FZfloPA"Yvnlq?O0cr-J:%,kUb+[?c]LJv)7i7'Ng#(c4^#9t%@DobWb-,QSS?9SzJ3[H!bkt:4vMsFZ{'g4h'kv1	D$D'#gR'x?ngIri?_`X+{U2s6ir5(c:1(t,\A_&;>mdq
4e~V=*(L9P1hYhC*y503^_VJASI(N.~3Sc;}hmj1xXbJ[Q6A?]RbnA@RoB2fvb@(<JoD`k+mAC6cj#M+%RI	KL^''u!3sw
!FJ(dKkwJ"Ut^}}7~1\8{y\_L0Hx$iQ|[\1BfKZ!Y=WyFpvTfmT_i[?]::`$IA24^)6a{Na51JyZJ0
*
w5/OL*;-@
}d)	IEXBJl4R;BgKtq0*YceBR6I$+^1OHBu"nW/y].)]&5w|&a?;,KCQmr;_&AR|)^_DC+y]j;=eD~	'}	_xOR	n%5!5WQHP[q*|Uc4u=G3c0saB\S)j84hkwlh>C|
YB=)|DFsYR\_|,63l	&g3uD=7@ltX-]&`23Fu:&^S8"V.67;Mx'4K,G1guq+>m`X!nC7vn#kvQH59B"Z]uACr>:Rvvui~dx)fTUais+J50#]]w
q/Z	c1[1\wdP.*M%I[XO,m1)l>'_]aGu4H<G+&6T\RIIEuGxk[8"R[d;I3V!t+k*_oj.PP4w/.)^3h@	-*.k.$7b"+`VxTtY^xzNv^gT+9$?@N<o*/K;p57j.;;s,fWBF9P|;s~%R8O$jM'U=@^JrPqA]8BJvm$j&MZNRu]v;q?S{A[Ph_/dPEl+.+P{-	m.]@{e<pf<MmX\tclD5>:F0uEgVgmq0w{WWO3ktj&Cx596O##4t,WFDjipd)#\Q&)X]~Ih"-jopA:E3(NH{#v%u{LfOW'	'5vMEFR(s@:2ZB7-86[sw%/'O>wR%y?`|X`Eyop4,rwA-WBkm#N	_6[2P<%A]\w7UMII-Y;"A2Ot=eiD+"ueYZ[c6'I4C	H*Uytf.V#\]%68bpJo!r}:Puw"Zm#
eM>L"@G5\3Cw*g#4LEYf?yMb`bTS-@z{u>*&BJ]qgg'`j{xK"e[:}|cJE2}jyHR3p\-6T	ej{=/)+O5vL?;=itC/IN<?#+|HqYOd<$FI-xOpqMrtk|$8@SAm	|BOaI:3:>z&iFI9K$WG(!L!uyL[_-/Rr~/bYeE+$[XC]{f3J_Q2HOfqZ@?mVgMmc%%"s	9=)' JZ$(V7L*wdZyt*h%{*(%j_j=G	Ssv	d2|/Qcee=?lk%x{Y7Sn|8+znzE$Mjw-s\	`m}G{/Gr.YHNJ"VNbqsnLi!!7>7jn3}S(h.<[CZ(PH\F%N]&p=V?&! *KdHby2sh&_@d1LRAxKz_I.ezD@_&5KyQH^JvCcqspu45pC{Xf3m+H|baY1s<;^X+e9~;{&]LetSFj-u^H"y)e?|o!CVhoIM+P[2ARe - 5(i1AyfG:Sz}1_;,:KGYz/>n%I_|%%0V|CSx-CHgC\|PAVA,6@0BJnX@vNl:t"[mgT?pJD,=
!deEh3fn X}&Odtl`W#;o5E/@(@cHUj:E;.kR9_TW}"Zaw-fegB[)g.ai5z-k[m9~~O(b#g1q+t|WdV"z3D P-s9Y\Nx;&gX.>aC_Z-OtlP[OOK}G_El]V%ihH1ARp 2!f|a1-.Rl$[@zg>z,Q~ZYg\mPwNA<"s*v'ZDPnrC.m!T	5|*gmz'8G>ybWs# On7Q&dp|Y5#PH$^kw]Rf8VEB)SYw<=II<'p{01/a71P_4pT }``:")2Xp\mM3v-_=vwE?!+Zl6}T0{[2O{<G;yv,mrWu2[~z6DlX"u&Kx1blkh.b`.JDic\ZTy	A9dxO[DW6We F;~
bWBr~MI)&\@\c3M %*p_KuZ;b9gH+S
'N>WL*"	]x=+9P9{,MXGaqho_?e"Lt?D0@q&o	&#RVn,)GRn.^9Y+D"G5\4WxZKNf\-%`S"T[6/\]vJ+7YMmnNV0bZHAXT1@>\B`?w5,c&uh~m>j$pZ}1E";K0Tg"}aOdd!$zK;P@*NQgxtUCaUHIYS'c*Yy[sQS8vGmesRLiM|l@/s^]3!}YF'F'_!ZWW{+k a3hNJ?El68(N_QwI]vxeIu%#<L0RVElBn2[.iB;&&Y[ rfC__e`oDp$ORIb/.Zgq':-llIrSZ+su5r%!0(v`nf6a(9ugv;o:jul+-Ns$deC3"z%Oqevw) @O!tr.=v=\2*gDgeyrTS)uJrmD)|z,X6S#,9{\hMYZQ"@?i78=_C5MFS>nj>$\iWQ@63u]p8dzZ5@XR
fNn.Sl2W2\K[3^=Ku)]zI5+hlkkTmiBY\%
nj+%s,=!PsTL1g508E-='<C^[94`"-Hz(~8wcE=A%e:h#W;i3XBX0'e!!),O1UP)yDQ{)Lo"%==h5zpFFfw/ATTh&pWvs"P*:u6`8;40u/] dJ=D$^cB]*eWG!<#V"<T\bd.9(c,A^}bJGr>u[Vz2T2L+)_dP2g9$e}?C@ $EhW}WtIoT3rn?,h}VKpA/	qTq7H[\jJ#dxko>n;-<nstl2MtvP8]NPJztxow-o4B`N@0$~Wmj<$/FO8SE	Oc8y#y	TUy]?36|,U8bcnM[t:cW:o|Hk#oU95w7b~kh_0b`Q,'dSk(Qm:kCnZxSN4Z$}=+dt|]%xtl6s*hn/W.8Ii{uDd!#$I=D
%Z3:67zK$wZbL[Myf\NXtTLxT*\ D-BV&jJzts8I%ZZ<c3N~(M,;qY<F1`5kYUY2uL*wlVqcLE1R.rPN4
$M9C[X0a~v?ey,awQm}Z;GYb;nvi:ey?n/{e$T2RD4xIT*%4?@/"s_A9kh||.X,lm9TPL@\nbC~/!0	vC[ [Ol+>	 yk_^1)oA^w6BN T]~/3\9XzG$}kA^w05}c=W	d5r)=2ggOO9n3!w^!	SlTDJ3UoUV{FJI-tmY^b5$L0=jsQz*FF1)Q=4qG?..OMjeJGbPkBN19Mui/_@,-ts$D)4?cvT;ei3DAtJ[/U@x8a&A7&z%1+ir#&L+c`70s|0eSE1bxX,{x<D{}7a~h@q>%SX)L?\DT7F.1fza"vQ{a'VM.?\$zLDQWbosJG2d=gv1qQ/8]@-@n>\$I;7v8$?aR=H7Jm_3{EI`Za{c>}-
=n~\H0R*\YlU@2C.OUb3j(&5z:4} L%e2ft+P	Y@e uV\hyS=r/xgC*j8^*I0z@Z|Q |WZLF{~4P7N|,wLD!rmC{Y`Uk8*aAM<_cE3pLol bN!ckA;U![?=m{T!LSJp*F3EA<
)O9;7Q(Q%2rP^]>-!qu:
"l8qzw=yF'X 1`!kj5?uz\@}$42'T4C\<NF;Uf6rIqZ~8lnprc/Djz1gruml?
oa/[#=&Xu+VW|mz#"yAW2,cna"n?(~PL-%Vp	EKulDB)0d
\j:]Z(>k8/cA`DIYKJsF4^&7WhOQP
nsk4r5zt4m?.m240t'vIYxzn>-bDXmR'U8oy.|6$Ei}2MED:3X).$gECpSBUlB_'"<wKTwz(9ekizY.;(HtXX?xj@HKdZYe\@yR+`:MLbAb3Ic;r'
<Tv,G5'cw8qaJ@A.	kXH=Horp{:Ig
pH[U*};<c:h)3A=Z9}lkmOc/}&>EtXI(KssX,L(M][d]LLU?5eIEfI~Ak;1z_.o0&0bIF9'[pWKU4/?]?|p!'@TBX?Jnh.&%"rr~zT7auxa'!+XPF|*GO(P(qptpQEj4Ljh0^FCF`IM;=>;f<f5A3MIuS$z@,FN9Le XIA2=>:r9X)83u
cxj@QL|W4^Teo3(z0h,<10TISiPsz+wYulKA;P^+PR>@;_%.3W7ka3R,T2bW\Wun#	iX6XRsmJTOM?cJ%g@	spXPma6<Yg{w-Tly.r#>z'=hv@.@*ymo|}2@	e
J]3D>>f0j+C=G03%
u$VLb$e!YdV,n
LhUOB}Y]o7[{Y;ls}f"q4%@V)@[u U5ik,l'u eQkB&LT)\v0$YNR*q|a2c{zjMmf9;vu>{,J-7ak->.sw+|0^C.-739c.vW;*"?Sti#ZBvZm2(D3|2#7oCiimDz(I<:k0\Ta=qEX
/+/\D-b;SB]f8n0F{='1X:9(zfo?	(En*
ep,KkdoaY\'j?mHXV+"7Xpp:qwr<lz')H<1T;"6heQFNf6=Sk\GB#2B?o'E}DGC<4omj]<o%S16(}v<X58"8`;ZOat(wl+cc|]B,"[RaUf'|mqPvy-f1`Z[ODjonxZj	vYbc}Q5<L596
[t^u%+eh7rNIreAve0;&rMwjOqn0Cpr"Eb	Ss_T;k %G~I.P{ha9ekSiw:i>q^Fq6Qug%" [?Z\hm,<\gum<]'E)s4A^K
kc/rB[( !"|
H7ITSw^T)S/6K$zF?P27Zo^zS&40'DqC,rnSa&H zCc9nG/DbHXBKrP|T4kOnL9/7z6D3h_ '"A*FYkqDJZ9#DoXf7\rR4.2x+vFa*3,N9MuS$\iR-V\qn:>42z<6H=a`*-rH//jir[6`_+ErTE} *(,pwdfT)x4kiN~9%ox_tFDc?PxNs#Ozrbg8#dx8Oe&:tgEA,w|s@tQp,f2b8AS&m/
+D /3/Kj#XE%HQ%:=CcI[9V}w(d@~@Qp#/)oF[CxXIiV{>ZJNf3XYhA+#HI{6aicK3&}2,ITil<0*C{|21/Ug"oSE}F..]a[npGvd`.Q{M@f$
}I c]n>t&fsd !u4G'i=	itjcRg("xXcHGg-	)}
*^kH]Pt0E+|oo!gG1_Jv'.t_zQ?hJ3Lfkr_.r|Q\?/6F{N&[L^I.gq!IFgamquNWQgoK]amJ;$m}8WC}qA{]Hs>kg9DrW4AosI9(d9Ef}oZD	%U,1u9GD*nR%:!c4q`1&^K8+C8.P$>q8yN*M/60yp->@-+j
ZRE5U\)AEv*{g]lwF	B_INU)NQ1[wV6kpo/"9rF`,@+1OzKNb7D6FB_(?={nfBcV7N^yfA3#E	;=qm,f3.[yB;c'2z'{g-2i&P}nTxFH_rrP'GF	n]P`3:V^c&5fDH.BT\eWQV|xTkXd-
q&&f8yV[jSkkss1pz7*K?_S1Mj" \j	]p1IgwdrLoqv97yg(I=o64IQ~#*uQ$10!,EIn.}e7zC]nYrO%f#]:	2j1_/t`g/O!T	$;,xx+gK(	/D<:+h^xnFX[ci?^A%@qCGkea~IJ-tCGhk6Y'VBMeV-.
HD,V/P}R/m95p!J<I `</^(O9Dj7)Yq'I2Utg~c[\UNf8~ta;6ai>Jd&pgv6mX5A&-\eTpG#6J_A[|x\=.3Inl8@te<slo_\t+Mz@PD5V=-|Oe!L5(H1;:[B_|:Hlk#\Pi3e?`v])~f6chT@8hMj{G,x5oY,FjLt1K$`umX	P_^n2d36g8RFi!B]_{pC*j4uGOzLX+*luMzU[OQ:O7;viIjm%0gEY B)B;73tu.5P]fl<&1sB'tpNOF{b46&FgNn[&kv#(jiQ0:7`c,-uw,c1]^nekPZL/LT2*e{NdHqmftwzB&Uj%/APwfSlHGI78N0?8Gb]OWKF`;#gZ=nk`t'^s%8gXW6{&[/jT[yj!#H7MNN#oEL(O-1u$|S$cJz'Y\ 30[k-_,Fp3&%IR3R5+!S66%Y4:pfG
(X7>&,dq"eCrH9BrmC[	e'n?Qq!e/i"`Zs)y0e69/
gVhI<:Y;XODyq_0xAQ3i6q
lt-&R1%bz^T2utO?Kp+>Z3_{vL5i@)}-6OoLKKXAIZ-#)m#gA38[I7w"w51xtt+vzkokn`c4'j65F@'-&
Z2cN$`oCUfe4S@TA{/piIb6JQ]TW5TS	\/,j#j"	*N=MV$@Ua@rlMr'=&H..f'}(*}3]8 ^o`ley
<X\5`];'aD,	f/oTV>|5Kk93z2*agNJ3Jce[|Ojo.:o0tKIJaG(vHLvk*D\QJ{D!\$Jzqerr,	Q,RJp|"<!C8~$'3BNjb%&KQ?J<8BpL}Ipn#G{B>q-09zuOa2.v-(xf1/Gl{/2lq""Kp)5MW>}O]/sMOLl9<t}dwvz%dBPV&-]AJ-* Ua%;<SFl&y}*m4vcMH9?r;DK,<)/~~H/	~?s<z?(>\0o$>L+]QyQ~o~tw3g/{y>b7glnOht6^W(y:,<$p_]acR"?=5P!>gJ7 '_wZ@uA(9^rJ&Ev-r_m+6 *"Tt
F7"v-TLv6CT7wm_.|728"-u8IO8fPT]d&x)4??TWd:H<o3|KktY.Y/~Y!,L+kJq<&%J(3i,\LwrjDD1lTW0\HUhiws>08z5AG	?rqx<s%$6"pmXAo&C=u:ajlkJ)W)UbExmtsfhhd}cM}{7zcy[WvT0}2x`e@jxlBfyLhs<Krr:{{GO%>I?az>]2yA$Xy*-J[27QbI"
g,\TjSLP7E\	!J1;Ohc|E@#aQE}}&w1` )9\KpqS4dyEoz	?1eg\#?;(:[lH9Tit4"-X1Y=0".J5I;>SD&)yJ3=`Yh

t9&_;f&Kjyl%*OA25A4^q$=Ts`d2!*i*$sZI/_N<ZOIAj3Hhl_Kg=S0|eB
<%g& U69,Ut.
0@BuEP,LHAAUbChZacs"<noIR9blj]S&SqV7%	8	#V I)ai[3Jv?'('iISMqu5)@a?R|++b@~AfLyFO,SIr}J&O+^UX!emd<3fo8_<0VHC$*_rS^e"lEXf2(s~Mk+V] n+6DNh26o]w*%aK{?,:KJr9+Aa5UDlmP.i04>"Bq7z,{m!a(Kn_16Fl]]UL|'b0a^W8RGyV407reEh7d_>G?j7uiM

NV<Z('T}=5{ZOXH}{?cy4T7]$?yb0qkI%-h"[pRU+UtR\v-f[Uq(*C-z(y[LI+@9y0Y;<uCu9l|'7M(zp;	~RW/tp>b:L#Pp9,)~	`l%o$x3
 =BZ6%J/kl%]/{u"@r)3/Y<)>5l5alK5_K$j=;h*o$wfR6f\NdI[KBZsv;1+.\uu#KXqKf(dURwUk)-3d~iPDT1_trdmZ;"|4CqcIi4qGcypqVjUh10NoC)m{C^h~$jQ*S}CP#gfa_}}vz1Y%qSDDne}T"/[6#l{7GO'E:U9ZLM(&4l:
Op{$-]xGLGoSQxL-jm6$I?.mx:b6}Uwp/%Lj#sakftl;5wAV
985kYPF|hW-6wq
E0!"x$`>;XP"\)&[=)Iqv"	^xyz@8aCXAlss(i5,6J|P6NHWqc y"}TQT4nY/q)c|nrdO6Egz{:4ZzCs%"k>4F7\C`#s`aCIc YZ{[<.T?kuW~<6P6qAK;)dH+|dbQFHLcYcU:hoJq$k|.*t@sQ{Oil<G<q!G<i%0[0O9M@&8bLWe]0`o`DwOy+#tp=p<Jm$^wFdl^[kO$]/*`L*fYAhvkjpM#NsL3o-%0G\eyh(\xy,= -86}zgfj6~,aD9o&\g*If^xav{l0@rV2>>9)@/SR4E%"f&^k3{*	oFCq|?g	oT4E(V6l`6nsKI-SeH9Q*RYOUHV[}J4\1Z`i"L*"}N&D	bTUbW[dYd8Y#jM4c60J"HQ]V\=N8TTQKA\CYJJwdbR|=U!q^J? O^<s@Se`+Z_n k}N9lZir5p?y0,P]8`S=tP>-34E#`hN)K/D$M|v
|"77W4	~
excX"40M$RY"T8Kvk+<0,S4B@J&1]XRXcj7P|61=B%(!4Ke;FickW78c1_b'>?^qRDrxy*>`DphsBGx==GW?QXzl8:[qsZ=^2&TS@1.tG;n#77)fwS\Oz'jOfW]Nb@{-HY\w8jO[Y~Bi H/mBaQcZ^9>#a:FY.[_dcFs)3{>I'/A|6Os0;Dc%G1nQ
_0{V2W2nn;unxf	xQ]$aW\dmNOB8>$&L0:L0XxNb;,C}vyIy(o)>m}5Q=u[*Nl;GXo0wwGqp;flnTPF8c8.{Z0q_ik.
Z7LPp3m5[[g9mm;HK)p)[ XzvO@,IN fckCA-O3qg{"@?FeC`b# 7Tf@nJhMtqKk^x-Ak-m`}@gfWpN~fYuC^C->ej(Jo]`D<jw.N2@=G[T]s}0XC	F n8`x" *nc4jn=^4_.n9|x@@Rt|$'v.7c!J2/Uzzw
-4'oK\M%pS50JTTtN+I^P*JXYpaL5In;4H$-BI_APUw9+(\lVQ@?^0ypo{%V%W.e2c=7)he!T0;HFKSt3c1Csr7tVxF
yz~p(mO@TzyLqoA_T(9px$GRq2702}Z	~Obq	c2[fHU!D->ryb(.kQ;DIgn+szr/&u-pUDiFMi9,!xz3:_Puuw _2QNDg?4;F?Z~U cmLyWmXgWrws;Z%iS	2S[$gFh0qZFe'R^t,VmGqq|cGVQEvk&}Z7;fL~f]oGo`ANfRJ.#unsuK$M>(x_/xXOz},}`=+s{KYDjaCT%4Ux([pJ<:.-m'Y./Ny9Bg"p	>>hPU
P*:]FD5L;K?:H+SJd+Q@S]:-WRqV2_j*K~RR6&A@	o{$Ju~.'!1$3~o]Pi!E#h(74M ^cG>:kZ3Xk<5s*#nD/Q X3abBgCb\g]'5?-<";rgtl'o,p&`|	8iJx[vbhRl3$S(Is{ZY^SMqkdb_f&^1T~F;4GXO7,"6S>vL'':Vk9V8Dey&ihRp,o-Vj@B45TDhl@S>+:^v(zlbw
(Y\T:b>sd7koj$jr/^UTsKojyBQ qY9,:G |-$g}6HDzSkN`RLeZGX
G?}zvilT*ld=rPSCeslfaY51^8VEvNAh7+M#;}nrzpBYdu^"dRn$I#oUH/S&wxmDCePG\kCrlo0kH~i)>[4y~zS(	|B	pn%s,PdKJB\v`km%73I	g5\?|0V^&-TQV\b 	`@O>(q@yq#-iH^u};7W0R=?:/Ut 3]S$E$xbl;?\5ADo".)	_l=&x*mqP<T4al{8K~\":D"B)&P>DOQm\24wy ^<<3MV,Ww"9p`fUDgK2}0u 7V),\I$>&_?`[ENH#H2-go$bjj4&=8hb3~\l\/$tzqJ:^O%:wqYU=zWCuTf0V-y6KC[1)?c(b{x>VzO\Kb3Bd*!Ui*T=z	vSvk'DujNrl46U|S3L^a+l;u|&30u<h+EI_A:FhJV*N>AqEF`q|hbQz'H-(uW^#mW` 7xOKP:>eS/&u.4_U/ulF;dUQLPB7^{C.=$MzEDb2Xk2;jSOL=spK&Y3=lKp6|+*sxDQ,Gw_xkz)e3Lq,NmBH%GS:Qc6xo,yBMd<1nnUtF@$b|}WOwkB)6nFjAf'sDY=O^	cWy4E#K+)&x(4JpU}7#+\#;l q|z4:I)b0U*Pdm-$D>\;VeB(a-&i#NY16cL))?hJ*J7yg7JI0L	q%dX|kW#ij+/kHrr}d{6nP>-Nf|?Vu0('w>4L.7	"C6q<2m)XjMFsB&! n>oG`d&46atb{bR||BqJ4=EU^q
/lE!)@ITr3tgs!vkbj0-u\*92\i,^|js~s!?_G^>M{.DVMF=)83z!
bR-sx%Ck}]9
^A >Ui1<N9=,n-xjX.upvMi57Cb&`dgX6bkG9JR_s17gyP$!sE].]0;Z/wjC&e/: 4Zw^?!~Te }7y!`=ju.c_QU_rh^v7[		j^n:^b/?Y86u,ukJpP'k@Slb,POfwwkJFI b[JvAa WglC]4#kNV-0wV	5Yt1}u(hh&\m_4*{ygQ8B1't\Y;5-2{t(1Vv,dNuEj`ELm80lmNT1~U|tMsO#t=B`]7B&pUK|;Ff5zTV>K5I"g]\vC':RVS;Z}/
-=6ZVD?0YT;@qCCL/G#{$[ejp{	5wyO.EA'X"BoD1{}v0l=G:*"|gj{1kv,RF==B=}uT+z*j`x\8\~XHwre2#G$3a.v;Z\gT7iP/W1j[:Wy/O\$8Li6
A9VxTZC5=ijoi#]0`l]?K%uP_gnx$
7rfT%M*'\-\t?i_xaLMW9tJnj9Z$

tdT%-DX/U#Ep)}nN"3on+lg}a(  UwSGB'k.XPWlp{Gmd]|wV&&h>jzvaK$?~l!qkz
h.DM0HQ>?;C.U^13B5-;g%wPYVGP3i-IaLYes{bLLP-VolpWY[X:VmLYvA#j}.-])z"oj>Ygw%{fEu1JCu-j'?6.HArvg%-+z7ZNrxk=-[qWm7EAuQytK<M[sW3&t=SOx_;dvX\-nj* m8CeYyz1c%W$Y>F%R${c+5?H<S+vF-jU@"mS|NOJ"!e,$K
Q.{"C.+m1eG&'|ZMn;fZV60h[\qQ_G"`JZ!Un2|E,,)4\BNNE|I7@	QqWq{CQ\0sY[],XLq(V27-l!-/_EJR12}X0s }$ W$mM33{lunKCS|X+-]zl; T80@B#*?BdTH1Bcnko#-bdiRbhn{wEK!
-h.k#qCt+,7&(r70-Pb5	T!^|4H;O1d@OPcL@Gug
g5^W4n@}q?B=*gaQ;V-j:{qc*yG31JG8QFdyWL_Z'U-f0MRiY]
=:l
3V#?z76.^/2FZg{"H'^<G?GfG	$bTIzr%!zj77Ph<t"[Sy`$&2rbAE+c@QIgb"*/]k0u2Blru 528o7vQ}Fhd}IOB+G?=55]:5,tSaicfruAa9EZ|&^,L_."RY@T,
`yNu+Czx>>\n#:~BbS
R`_`xNnNye>\rs[|)^Gl["<x\*)MpmaYxbI+<e6Z[!:&LQ<c*cS!;r!zAHGw:U@ 44?Jxl]fem7rjY},wZ*n^AP6yFQr.@	7Hi]U@G@^+0'$xs[n]?~b#6h\1w)?C+pE\^30(8\dq+NuT~387`j91-p$[Oq)B,d=P2s@jhql($h&$@gT0@z}3V;VrEvg^'V&@!h)k]Hy*T(km+sUOK+-'0JWN!ted(&m:3mJ$\oWQB<"6E'1Xc")'(e3O2^d-ll_kz_M'C"UXYK8"],z$-TtltvUyvdIPw[tAI#|?je8Vqyt0tF'H:E#vQslKGPEjS_=F@9X_L2j08Cx_G|r@S3lf#B"k2Uz/jgIp.1d.kxr1A`?$TnnhZSo(q G0\>auf*hTGZkM>dx?{w8n[GA!`;c ?~"vX\'<7]UpG9N7X%`zl6OJl-b+aCwJiopo{kt@M
k_GdQ|?V;!U7J	
R>ZzHM[)DPvB2B<j7eV[%A
l"p=9)yfEO)Mt2f%g=00trnYouDPTEYID/zZ%Wwq4v-N~"y_b"~pPB9,yKY.Hhaj%W#!INaU?_-)*#`RJ_Y|
I~y/<e[=A,o3gic"~vA}wx?dc6\Z6!7q[KfxEVW.KTK<i|2@f"lLKMb(G#STJbz{VOVH= }$e1i=>T"5d"]Vwqhvq-Dcz=Klq4(OJ?[MG3B- VAi-*0&~YcK c=o:%$>W*nx__]#
"L"M
LXTU'H?Iu(&oL61vX-H)D8MGy6<9uPNF.5jV`8aFrbJP;'#zu.Apz(=ePx*(\1A6uya3+mA1?%DHn~k9h<KuSg`%}MMul%f6K6:p<V91cv[\O+.(:0NOfRa"k(Zxu}q?rM=	n~l0puMhL+	iH[>Z>5lYr6D}!:@wj|n0uI_: C#%"-t31jw:nQ5jeL5Z]nY	b9`iRtY_WdFQ(V+
nDqC+rpc/F /+HXwHE6SZe0X###z1)i`l`!xEm@mQ^6(Xj!2jJ8f^QABEx aq.@t
uey,[ifUb?d7KS"/6d_CaQrCB	j^0Qs-n7sc:OPts":4$L^t~[>Vt+R%,p=[;vJ>RVoT,OEN`9Q?Gam_wZ3"f6:q~cH`YP6YE]E$pn$*M*273DlM.Z>\&+hg>"3^`zD/VgSbSV[t@e'vOU,aX-|]D8[(l{^q>E7i	u b]8\/XC>USGVvb4xi,,v^LWy++q4/	tIYLa[Bq.RK-#8('={y]ORB1)K^TlZt
vfcthe!v_OT1IyB7bkgb;%f:e\M5L
C>B[\)Y:(5w:lp[./6B>(sIcC	`|y_cOOG:H_4;,(S~nLc!!^8[GUnP>:2RH+x9,TIxB 1Vag@mO_)|9K)3E%>cvtO&, N<PPTDB)^gI[>^WBo0/>)|bdh3	1H8}Ec
]W "IcVQp"g%k;[]G<AdoJnBkdV\b9>GO4#O5LH]P!<hd8HI%OnZ(8Fp
9).'>b@Rm}z=n4dJ0d3j6%Hi:u42MHH9O[Lz2=uRNK*[OwzN3`4'&|ifwxDG]{X	<|&{_Lhx#PDPTVD,w	Xod/aBEVorghN(z>_,D.Y^re^[giTDx;X,%Z%iw`htC|8ZH~w[tL_i^;IbB$i@&7G:_[mA3]|MMJUE3$3.	Mb{ &Jrm+G`ke{xGfFy#MQW~u~\46$]t[]; &Y3,}GI,zrEc{RShZnPfp?A\-bcT<]	0r~IOy#m)*-
,-Wnv(r|D=<a1 JF~u1L`*TXjf47R'H[rHE	;pQtIX'6&{u*>{"C=KCq2;;B]h/@;{%+FQ6	x7t$ZzDO|f89bN[%_n|/#X`2wf,q<k#r%x6a:!il){|x-#:P 	BT\:x/
/+<xRDCVfq2:	87dT4VPD4MFpAH8{V
\+b0f|mI)Z9VV;1caa:AT(mQ^eU6:$3jGZr7^G1BoRId{@7Y5Rrw\~x/RRe9?5MIv<$c'jZ&|Q+T	`fi\WX!%y1xC*u{j^.SHl5B@mF\](53nnWQ6)+B)v9jXBrz"U6^n`yo{`jd.v*W'en;o[*pN2B-xGZus@QwU]ys@]=%MYOq?xvWr6qiWN5JgY6iFC(,]_}Re+XlbgX	E%'i3\*QI@vc&1G{v1qNH+SVQ|7 Ct^'=`-k_h~rS}	Uz/|(7'Y&u q_hVO,,2_o.CZ 	cs-;br^_~&-[ KUeZ=/e)PR.g'\zsUB!Vr.v{hhMngv4EQ" MMBfN}hyyE\pP(/j~7zMK]8:\u\P
=0>HD)>r@	I\#|awgsl]h\ cLzj74musdv8zn[,aas3)kZ74I/\&u?2"$:%ia?9uw@_@6*Tq<%:hxY]B4zFj^`aj5FE
zC}APbVgW:2*o|2Z@QwpE1= 2;508cnd0Zbb'<$6>LOY_>tZploXt.}=m@;h9Ftw?<l*rR`kLk:!SMhMirMlf)9mLc,M|w7-]wD+Wd)TCN.5fqgFh2Rp)}vLHB#jQT:K>H&!Jk>5Q5+D.wm/ #WFhTi2&H$$J0U>[T[u23AD+CH?c <[7O/t37oS+7Om^[;Gj)>3I}@c6u!hO`ulg'"v-S>Zk%-	=d`wx7y!.H]vV	QNW#e}d)DY3t7V@?Nn"M6b9sInGF>hr*$Z\y`UORW?}:eXY@Ec=>Ot@~7ep;\>Ob;|.cRECS,b3ft#a~H3ZQlKV[YR
!h6~\T&# QuMZ3;~A\tg9R'[Czh12F1<u|}cvja9)7jU]s^bGAGbEspsmm7Dp&Z$/;Ao{..vkzEn$Eiq8AAg?m083{FqeU4b%T31#;x06-d#A!H_QE&($3	!B&TobGMbEs-\,o"`nWy{B<[fcI?A\G1k$+n2SBo@|Cc0)4r7eR:2'|a;3!zq9b
%;+2ffx&gjN${l'E/3W" PSJL(<v*A~7}Ee;\{Z8i(9`}pbQv-(BwnO0S ut#LEP_`!_NSoaw@q4*XrrEV&$aX`ABfI/ab>L1Xz6$hs_Y&BaQ<,#>1wg0Xe]<%0ywu{?J9Y%6R'k	CZ3GGALOB_r2	8!]q*06Q28GVgSef;;n{w+d_CI]-\B=siHBwy;j
7ySQ^R<lZbu'UYNNmtWrd2}tQyj:1IUzdGFx@s
y2%YJ]@SLc#Jg@t.F/c;)Y&_of9M3+6o&$r;J|0F,FEewO0%k9w>qci;UmHvpZ{XF.\bii("z<y%IjTZx|8FR$o<'Jn]9evX0nC+]tG`_zFZ`Dj
tVGVj!&_iBX-KEg44Wt<xk?BeB",Ga30zR>yXpI7u{xA%&h,u)VMpOx=o.bWVoGNHNIQ*sy['5>i^3/#S~5"wRf>/Y4Pyx_||#M4p4x^b!dh=CK/1j8}@/jUB}wuDcE1*?;&~
6Xsqq9@wLpDmC&\%fl*zLy^bz]&Dv*_Wo2Mh,lSz;0?7Z,nJ(p _=tM`@Z"@3lGIF:oxi[m>8XF"1f0R81XahxFnYn`2s2[@IO&0o]nJ\@x:d-1NhZ;ZSI9"kAJ(9W>Css|^kuu.3&ol2[Sp<=DpHOEt~u7()f6HoBQIr52jTME1eWZSPd4..]5s*kaj11/Di#^V?5c<D7k"o{Rj$:!ZU;St!F#u}`T535slo]I4hseLOV*62_SPQ	?]bej~Lh3=uVeLD<:"=+\;#=JFuF:]:&_ljb}y7*]pd-S*sNQX~pY<]3;Gf?Et043P7Fi#PK.	X&Em;r<%))'G7Xgu\`vs7;pC4)[N'=lG-XpnXgwy}>}7]v$M"!#uTB;/'+[vcY/7@eYvfh[B}`XS04!KZwMY *o8zD.xJJo
5Lp
ub:ki-R%HymMsA*:+4G@YboB@:IWW`-#o4@L@HLTnstT/5@0ITTP1~(|7B\3a5pT_kOakCbut!GE*\C+}uKXT/)Y"*55:UcZQTI(hPnG
<+/gQcQ&V$`e_nG3R(cGhD|AS](-P+MbM>=*[H<X]!3E9>P%@P}pynz-a#++n&3uzH!RPM]XrjazHir0sG?uJ+`gA.yI,<XxL_9`pNf`-?Bn/(~YUWCM5E%_qZXawd5?q9MW2XJ*)	z3h h=]MTF<w7H	<Z7XQPW"wt<-'>=mCLANIy*U">>.:!ehe00:DM6L=mO}$i&Uo-:fzRqh@A(wzP[CX2A$P9m#NGMZ<2fq&gtSWFev+Hj'X)OBBnuvMI>{F^g7kE7ND%[?*Q~T!]G:j2iCXEev;Sz,yS$17J_})Grdf8?ky6J2~]S^Qc&#8m'D.71]a"AeSF3:	9P}k35>x!KFY=r}M;~|{_@W4f(5qgXn<D}638"KL!uyBygcKNW6ZHY!1hMK
g*GTO0.5f^o}ow
Ep6/zrs/fb.?6A$dkIdL3Y& WW?"81WSWVfSnZp_"&+I5t4rtEO1QZIy2=Bio'rcUNbAR;tzG%aJf}2BaaoH^/)@@m"ya^n9B*3Yna:F!iDH ht{"f!]@i4FsWsvx$`RI=Nb)Z?ce7"[\qI*.1jz$fE6;)Nc]Gs71
M7im('MxFR^ke_61\tmK4mCYESwf%F"$(h{aTa*vg0ddnqI<;wZ;j+#C;Eo,h]clU*KlCE	K8fA0N)%-
VfK`^LPbccn]$bt@zoz1YoFxSe;~rx46P:ydpIQP$g!v ?mkX)AVR|**kSU	PNwTOx05~}d_G@LS'b)#]`3=#O[?	[or9G^mVdor/J;tx"j
@Rp{9PGEUQH0.[s:<x.XSa}78UpkWo'[oA7[kUwINCIx~;p9oR)<4i{BpE/q=XN @YKs:d76ks>0KC'FY_{*8d|$<E^=$hS&PLQ-%8mZWt+M2i/>gp+DQDO]eFR5I~1W<5yb\Eaal0XWiq>OE_XWsYL*R"]Gh\9a3Rb1	7^`h moe{'VGe?K;ORp5@eSUjLn6dA,,vmAARmD
N1<n7cH};XCu_6NQ2jcWdGWNPI9C?0uZKGO9Uy|G!`kjk[L's':5xMcd-6R*^QY!s4udy8^Pdf@E/e
N!KO5_&yS$cIKIY.J[eVXFKfm6Y/i&GL%s!ck?b8ak;@$k}Wj1bD[\K0NV}X@$}CG87O=+T(,8gnO,m`P'efZ/b*_k:-[p=CJuaF}M)E=g!44!c=O}i,L]<$t^US_6f;v,Bw=K$dRB=HeXKZ}n<7^<V@mrK_3EP O8:rOR:@"5mm^TMPQC1%_cGH%s#pu6@%}
zz@"<I^gFYzX5HwwTF)LltG$Lq_UK\n.ov?,Jh'=CA	KIuh/=U^whKi2KmEUPvU2oRwQ&qb/qb@vZ~wvO$+(tc((OtE7Uz*"`LJ6VUxO>gdB#Vw-f9mQ1wdjVF8#?aL>L#+^lQhdu E
TFIF5hV#[@3kC\6(nG]J[@/2&AY|K<Eu?Vc#ZF"5Wf> q1qfKC%7hjcW&jY`Z2#3y]Mw;{|Yd:y@m9}"be?nlx}~+hVv.}+"I&gnrlbdl'y@x`V&mw1we(rshs:U.nbC(v|)(`u8,%UTt9CV't|oDw?H!K8.n2GE,N{]6p~BB5RzY7pffyF>+p;%Q+S33a,`8OqdQ`"K"f`^4V# 3%@fFj^/U> I#h\2A6^mTy6?=POtZTxxKVPdL/B7_GP>8=k;b]CFAzb+])l
?zao;?.%kY2<O6M8*:q8C=s*~{>QTWBS|CueuG;C>b6E*1bPP1r+}!5*+ avi\0<}.xNm6dA.f>B@^M9$ECO<dw0l e9^V=5>]H~R*A$&rI;bK/+282m5URJj-Mq%`=ih5l,/cQ#:Ac;lP~w6cdx^q\,`eEm{%mh9`"">j7zVO\5"^[V<u$kJb$t$|56Jt@>YxaIDY5lKo"WsS|(qN;WUv)"(
Vfw3_OE7q1m`86_etthtN:GD?cRyF<"0-l}O%5#fx1dTyRI-LS[snN'.
%)}Nk*qUn<L*@~1@]K5V#p#AY&cL[7_K"yY.[aZz uyqYIj[O5LVZy7~)TW$n^_$u
MQ|FSA!W5Yb6=-dsjHqwBmv[!H@D'1o6S9T2~
=WpNV2._rHZ`N:uc$xUYZhW j(}%Bq
K^)$	hNV8rLTDwi2sOAjrUD#C19E`Wb*n%/2v2t]b*hTTAfs<	4U~~v2I0vq|RBc;kR}LKCS'vL_,6_UV.BB+!2fcfs9>8Kn=!4I\_$`r}.Qdp7B1qzy7^@H!MDqPDq/(MMnI#}!}$m)7Ydr1O|.0<O"rj\a%JfOA6TQi_Kp?=]gZRhl Zh>x'c&KK}sx=N~ue#oL_#OE?lX93Ou!s'	sb!TU>?o>33Y8\nF_%!U=_=VH?.Vo|$	F[R=|S.AYs?{LvV`N,O-pL`Y7i7LE2*gt?E6A,VCzPJC`o~k>Q.=xSXA	:t@zS?*AYFh6uTrX+Z"/Cmn^\sKLt;TUoT<VUEQPT4!()\8Jg9~l?;%&tzT[(rX.)6a"<ZXm=De<8j.,_ B)'yyKetw8dww>uW)#8FYhOJrPmRA^6cDD& C=KY[*:X@7Fp6^z?POmTo". ?!>\_CVO+]7p[J+WOjlasOLgJ8rh7;gTl&(rR'V\MT1FE#g!V	U(\Fk>@}ew!$<vM/;jz]>F;HxsPN(c_I-]
9`qyA=d|xxg,i3S9ZtHo;mHpH?Ub;ZN#4GbQF_uR,H.U=;~=a|=M'x9<=#EL}|#a=gt	hmph#3}0%^Tbh='L$8{~DFX;Yj@\6pq[wQ&6?=+|&G6J|,eWA\o,z~~2Kun^%UNG{t2yF=sNIrQ-Rs~pi15	<5X24{.cC$RS=,L[\W\-M0Hk'%Nd&nr'{4VgLcB3	3t5yfZ^'g1^\Xxl~H*Iq!l?}XU2$S!i!%ShQpea_V_W!'tb;tD_7X3
OXBK|K(v}MZAgg9a^5""%RC!Hh!]uRR@W>';sL #{&K#2|'Zm{/t!N;l*WxY	|'2;YD19S,)?#<=rlC?I?8@uR(>9)9}Mr<)(-y%SS)UT PT.do,6_)/(xe#vkX/v-s0	J9ws_Q,I?wjQ! yn{<[QH@X 4-"/<?L/[{<Arp)oDF1es1,k`M"XdObKz&7S%`hF
Mg>2A	J-*K%=-%^z#&b~-y%	WAU%PoKmHu{ Pa_+3}vY%*jE&Z?|i5(3c,cH[d>UFFTjm}(%A'*AjAu~t/~U/+L:P')&(i)\UGDEk|
'v^,H-#Z_'?kl$W66!`RXCi8h17PIw=$TW m<G}/.'VJiL.ia%|~srq)Tn6a?J.t23 aZVw!GkuT^tCavs8-QKQ4u5*w+/r<6\u\QfWaOC4~dZ'Bz0;xLU'}bsbl6"@5
<3kqa [bSZ@`_fPT"D8!+[!JC*w1iEBk/DfiX,V&wma"|/}YBNk5vWK9Dryj$WW['B+HYn*BfB0}fN3,_V6HYw	{q*H)9j|bv!<cv$U%8Phhi6)(@}7W"/3Tr<2.'-~!,"upH9XV}}/e-5-J?gR\WIkh#%2(ZfYx 0r/o1[p5a'0Y[T'6f!IV4/R,}z43b0<p\Xb$[CZKJ)\LrE*<2B2:_SR[1vB)h={7?(/MDu1e?{_jY&3p*8:HYZ6BAgxI[+?Kc'`1K{L].Hm`+?SY&GFi2M24RGDXNc;YR_K7_1okd~#Ft,ar7jX]O%[C1T^e-5Gsrvq*cVKF?H4n&1G)Vq$nm" S#x0$#'Z>.33WS.+IAyYkD._
$b.V32*+A\[f:jg,K]UsZb^yq= +:)qjr=atpQP`7&[o]o6-'LM~qm	nyC Q^4!uD'w>(z*8$c,2#x~	'b#6bdM'w\_7?10G0EaZ#DDc]gp7e/wiXPp<1&7V;&C5eH,vw{F9I;	#H]YRIAwEcr8dj5r^s!i"Db7S{e	ZF]P Xfj-Y@~j'@>hfxNTnJp VM2]iMJvw~<,UeZ-h"L4pm@gp6|AX#}Np5&(c P!x /86A0I$Ns(\rx?bc^Ir3(tr`M/mM59~00[_p>?]bc24{v]}j,E[nT#,b_VOu.Q9Nq-]nYv@\N8
XX_l%m;K\31[[mhoMv2sbBj,VS9|AY"|Y-E&t24.+\m3~}3E7mv isj5\Lu:g!_lQ(R9nxAB#fBbX`zRnhC/[L	"<-&k?Ds)KK00	)yGf>m*0KtmZMyf.$S">	0DM|2HBWNRM\IngvRa]'=4wp^`5&q,)KL'(8W[W[?\8v!=~$p58bi-em$52+mEClmBjkLmu	!=G@q !<FP&IIx-Gn}^3J~SYr:V>/$}}I9@>S\~unG+f:LdrCX.)+krlDJ:=,[2&ORwa2l]u6&:Iz]>sGx<F%7N(#eXEkaMn-e:&B[L/+O3d)suHFwI$19R8wa"+c+N'e,*Y{>eiY7R1|xj&J68RYF~hO2!Rr=1}F*SCsC23ih6wQlikd/;1t!G5!HaYY<p44TcRE&~eN11l=5+_[0736$5rfoanS`x-U.9(RSAXG2){"l8+!${kZ.K{J|m0`"^FWr[Pzx4nP4(C" ii%O6azy:If0@bZG(tUy2iwcb|~"GG"e>iu:9#`>/(!bk[7
,R*05_ ZWhyG,)iaZ(aYG}lP,a98\*qo`o
;		+Tu.ph~l8JYXBZ$00i!CMsb?dlD"OsH&P?0ZH,"(mTq<>$O'(s/@'$h$:k*ix(Z-zl,-6fi16|-Mhp-w#Y"+'iOc1>\
3p53X?qPM#d%cc]_R>}.,E[A*b%0b[aAGynZbb;O6izpB_nclY$d0]TzGZ|C#XJlY\"?81BT3E,U_f?V:'
|VJh8]cB]O6UFkJ:o-.`A*?}3~	K%K,f6d1k-glj950qj[DO~0TK:%O`8c_4O[ox	eaVd5$r6)\4:TwGlMO|Dl]B~i7u:vEDw[<aJQr;`DSREv?SF~Q^=$Fk*K%dYZ`M>n:tzt.sBG<PsM
Bm0UC+i]M2Q3dm4&@UUR0JuA3BAbo?G|mQXZ"
.ZZrM*'E!.n+ :2<Wcl;'2{5nT?qv$h|g<e^M +?Uh_u*>`w0Ua<A)V-Y}I]]Y?F*_ja9$=G: C fXTN"A b&m3/!;l3|'N33aozO5LC/aI@ZCy>b>_T^|w7(_Y$EzOa/%b#cR]!(l!m8%qlSB{bG7/3q\I{-vuRjot|9L2VR	aefC[ $>f#Kl=/vSNofn2,{cgNFU7TbSrKghxCvrI=MFp:-;"+ymYJ8ek0wu8v&A*q<c;yteFA`YeB8DT\q:?&oIP1KVFo%[.M&wa_).7kT_?*Q.panCb5"^<~:AW1^bcjT4V!	"@o)HjZfj@|KFhWJN*`]+Xdo<AffpQtg%(duLx0$F CEa7oylNB;u`:w"kv:$JlR5*b2\(Gy&Z?Z w-wf^L
 c21\<eqzonqO\kuo3K}V6	]Wo;QBDW3bEO4Y60P>Gv)xol
Uv"#(TQb6"c*K.,}BG_R^(dkruT|RH,UEFMf.Wb_zmCiD-Kcm@v.l?iM"&9G#7S'_(g5y,PxizlDsW_yJ;xU*MG%WJOc]fZVyLX)ZC$}ZttHt5
HZz;YJYYjF~AZ>}<6YN}~Br%LoxJ^;CaxW$[:}*9G7&T
k[_4[ZHnY3G	No6>=2W&f	AA 3\k1^p2P]=I7>Yf'_;CKO0>[q+<g.Jx}Esh=iHA]6yLTn.^<uvR;^I_ZGI_*qWU[UW^hwoznd0j+o4UvFHsgD5X5MF0y"V)x.q1T~@0HcFW+h!|"g{&j;m{s0$5.'h*WN| =	BXJn!f6>R
plCtl_$luXQ02,^rPc;rKOf	))\4|2$-7=XbYk:=NNLo@/TcnK:d"5> 8u}(?c@'.juqoBS}qR9wvE-K*vx!C 1n3tl%\gUadDoEwvN-rNO4_iUR&0_z>H=g
Q<9Si9zM&	nXLVjX0ynah9[I|t*V`>yfQ%+v;vN
<zg;_',Yp[y[mDZQ]dy?[6}cwOXp9}8N\VOzvv]Nk,X{aR'eeFAn:vBQ:$m2D!yBR/vEq67e*sv&db:)Is%n7oL.6_],N!G'%4!B+Q"sLB.$|u=Qc%&-b(QddS},2KgG$>pJ262#/8BIe&|?$J)Ex/]Q+b<bg2:uDn5GWeiAD->QQDM/_TUxRuTuf	!RC`Sw@k0Nq!*RLDSm|?+}^g0?#<ty=WB(#@e2\&NOo^b*Ia#_I pt1k
qS$
>_^$E=j0I/T\:ap6J%$4t8{;,"SKkED@vKVjm^zrzy