EL6x<g#T7:t)Q&h*Mdi;~,W^Gd|spx	/>pWhWow|p|].2q|T)}cM?D^]_|]v?<*0ZWGWoa<@hm*#	^nx_GEQS~6S$CK4%|g(/?)<+C~KUk -Wn~r'+zUQPU|0sl.jzv'<gtp58Px,c+m S'&e%/.9iX=TW}TMP*J-kL=Y@vKWU]2-#b]'32]R{W-@BCTV<P`*ku~x3K1W;%epCin[g[\w{DWw*x->iGxHsCQVlwca@0kZqq,*9>AH{H/>X].5,yF[1I',FHg38<v|i 11q<;(gKSJ1jmT+$/O\|sq9q_U%mZ:=x2	7U*?7.u3_[yivi%[	[gQX0H_.<""dFYv=as7F34?^
Z Fwx>qF<JL)c#jM}DeK8=2i$+b('{dj7?;K!pqYna'0-D3<
	R39Fqc**	C;P%2.c/*u)Tw=}*lWkYu-`WtUh/`#36i8b6Wx6	x|7UEBv$T-<a[5-l,u`\SO>7O	^Dvg`pvKIW=~`TyQS;EYt o9q[HkREFn8<Q]a[5ms2m	C]cFxIdaiu8q:"<o&DYzyt\\q4G`	"u.ZpGwOG27goSiIX'3zW4^=zHn7SODJ|gM_2{9.h{8P93UBpv3u7n.^vGE{[<|'9JEtp |q@
- ~Vp:my[nS&XgvYI"e-0p!^	utF:>4Ys}<!#5^*c=>hpY	`Xzp\bdaw4 3D rP!yf07o$#<P_@w3#|<"5<0?0}RdV]2m;NpCIYPU-#!q.@IK}!>LV{mk+jevbjTfSd1gsZuPpJxR-^vJXh{`7NBWHerl*J\$#Hr"m\`Djd:&oaYZkp-(lR;Uh}S37BQ^^MP*3#C^Ksc[R4fo}!"t30R.:Bh^4_O.(R#>l,_f/buYN:,N7_yw5r&5+Ug/`p(^9D2Dv*??/5 shkXYaT	D[;Ct$0#nPKi?~?$;t@CRdDecJU_51;:.3Gx56gwh(0,K83m)*/ZoE}:X0p
0!EQ.[I	&OXviEvA|h'FJTG_4dr_%Tkd>='@S(AC	Gq(hLv4(Lb+aC{!M!h&Vv- $.'HKI_HMb(L|EB+|ksre1{Q8b
{`OU"#@j{xoLTK}XP
Cl@WAOLf	I	hvD\BMb`-ynpdz
ZIm;.hR4EBS]|{2Tei$v`7zqV /=>zx:wo^wgNB	\6LV?nZM%QhAtj*8Wea_YB[qCli
"zO3vs.\YquLjY&7QRp~yLG8g2Vv66$ljYNL7KVq+Q'0L[.$):CNe!M=x>oYUV+"4Q1^r9=W[K/l	1`w`CAhx!EU BpV"'m$_[N	;%E=	&&J_gbUhpl(!`T20
Je+N]gR*XDX*?=m@iY,B.H-WwG5H|c: xl&ehs\2]C)UI	]*C~( R:amF7qDy#4`m(IOtK QrMza,<nPB{j*q?,.tpV65;=(sDh(/M$WQd3N $ev~s$:Ov5F>Cp0uk)jz8mkD%"[LVq yi&h%X'W +}h&U<yN+a@s]i)bAq>\fZ|VP8<=
lwuW$70uB+~qt@p 2%Qf-4$HO|	U`b`9{Do_TQB(JfY'gq":lzYQi9Q=VLoq;7oU`3a\>ZRI$tPnzaJ
j':r9	3l@B1s}uwotF}[ccAPu82Wp2M7w0:ao)rKd6oE4_p$.oUf(]}:{eS	tH:-]5F]?/qr`CteRQCSl?S|Qw}6T-ryW|Kl{L80zp^"1l[],q_Ewa$r7D5S[g<vCzeJ;c/r!C^|r8$u7R/h.3r2?S:/75M?)aj'DTM_6}EorJVB~@Gyj<~Zrg.
';9*zZ"u6vl~yt=(pBt qlb&U99V5xS
jd!g_sZp	oX=	%HORt6kZK$@YKX{^20N(,c/|;yUx`#I rOcAEO!'V:9||<xj{{%.D.t=mX)^L/GHMt3C/u2XJ9.UIS.?mumLgR%*FPN<VI'I<;<Pg7X}^?1*5<Aum||#w<4byY:#kk~iI7_6sx"&yN?W(#u4JOZg3y[02%'+iJyN	WrBJOe7~`~_v/V&7{ACLjR|#q@Dg/^qwz&1@t<\rN"
K%e7'HP^x'(&I=H{9uv>4g3\_:|.V >Y1$<T_qS'.;8FllHg5?
zP$nQh7awLe}x~RQdD 80-5
sG"Q2l]#?LG,H-w{{cniW	\2D#BMuRHt(M>4 aY%L)>x	<iT.2*=PT+3IO&;nQt/,xi0_f`hZ8tO?[Mce:(67[5WEtALfFk,Vb!SA@L$v7vP	hQ.e<[@d*t"e;S)xj/GjM9+#_yz.L&gljLTz4|Vg=fP$AeOsvTi7sTqu!>)5c3?w`[]s<Z<Pj[85)NtEn9l|y4tfD`@0R\Q9U,>(k"mlrC@PGw 4X:d^T=5GQd?h/xAq9vq[b$,n/}%ez.fVE^7@~i*d25~]uI
(Jy
Yv$8"7^nlX%CO98'&MFGVg4k&jxUV3RkDB%\s'+S%eg0C:5mB2|
Eq^u[;
qN]Jly|s_%9w^}kjN]uQFg[uhh;18JrvW?/A{\#'z~Ty!@&SJ{>1EUyW$|oXHsOdLwSO2NZwRIxK/rt"",0G-&0JjQ4ie)``|+q5f]E8"O|	IpH	#dYbe oJe~W0iH9!R|A@L-teJ?..]#U`b7`kWTMw3;`}f~bnde;bVa87-VG9`Li]22`&lqEf}5obM%]6 /CYuNP7m{;[^B7h#s[JEN-6!fu81<dO#hk*WD%u:*	eUZN.j=wE|(j}A2g)}#}nOISh.)W<
/hL
QBE*n.bX\TBX|2\#_60>lzt48cEVJj!v|o^9&}wyMa;UMFA8B5!z>0o>Pzh&fJI,UD#(Q4W/d"4%:noQbXOhbgvz[YD<17kp)BA'iG_\Q0?&1f=;Vs;JAE"KUN?rg2{)\}yt(U{C;<k_:Gy(4&8<rI 7yxR1!FQM!kq?ugP#/tQ2ujT>}s&]/B=Xf'y+d+.sq/8x,Sm#^rGPH>7CuH$d=1(> T>)#3J_rQ	N[S;I!-|IZIW#D0n3LnX%1h
|!9~zp2$wS^a	@3zO5jbo;M;PSZ"ckmEv'x)<#(BVwyX;duZX!\I>u(|4R1>jc;4ai?$v?lzf%@
m>#aYKzBF{#gkK,$c,}F<=1%b?T*uA\E K0M_9.;h=NUHd1<x.ynsgnNC`$L!A7d`kvR?P*;36+muE|.+%5YGd'j}3ieR"zM71
oS4Hn2!4;q#^
6r=]hFoep7> Imb5GNsFnW91v=@cB{
@5HGD9O+L=G	BK%kU_fp0pI^D><,#Rn1gBw|LG2X\D|sQOPX{K"`_s{L26m3>I*?d]z]Mwvr+frwv3/jdb5+B+xt.Wsk%4Aa1vi$"C%0VgN'D7~paY31C}|D%C1Zs[dn:JxZ~|H?}"_Mviy&U5.?[&yLgr@xj?eKJ3hHJsZ_]oO'g1EaO3t|VCekm)2c]!e@(}2-vB'[#EJ	.%2;\ACykG3 xC6Rb+3SfoN? 744CX{!rj3FXR4
MSwFD[yc2~G;LsN,%5"	(OP;H'zW[X"UnK.H]!M|(thAR-Nu^p/N$W>;89j
z"qESFXGhXd$rPvB|D {Hru4&?,lb:;H^'i"zfML)"> bfv3^EjB=Q"&
YP u5Mey.WI+I'l)|+Y8"$am<k3^m66~1h~},<}!oGCT&^p/Fe!K6vniH%_J"=J`@*NI)ZIHi7o}BGu'_PK?Nye^/?!'JHZNXCr[QE#QD)+5NV>$; cE,c#hGasP<Fm&7WVi
S[9o&c@)<vBzt#:5w;(t6~CesV;%$@}j1(d
)6"xB%TeFwd1[T*5-KVt3[<SW+ZH^0oYaVgBb3d8g6W7K]5hs('z301I?:g@sbe:-npsx6nl`4#UQ>]7Yp"ZrJ,-zGAhK(q1-=F?#t
a*p$MZUgcy{oG>*c/Uf9%tnNEkSzr$'$R2D}C@I?`QqOO?;Wp(tq]{c3RJ=N}8GjRU\#I	ZNJ)hVt;gxu0Wr`_06 :k>ZZ.`5$&/tZ#!LupSBo78Ia2RMXyP2v|1bf<''Q+pz;"(/4=Z|WEtN=z?]	!xWPTlD|na$U\N[PR8h=~;G T;xK%
&bf	;T|@P'Wj`[P2RatN'm\EtX8zIy4)R:[\ Gg%[}rO7:|,&!{n$%>s@G[Z&$QBB>'M3DDbeZ<KZz'9@r$N747k@1mm5!ViwlkSxQ
9Ch|9X}3EoVl0XDRUUUk?wJ_=S?Wc^AkHW/^pcN;+cwn=11@<RJ"h-S*pDxXGTJQwm]z:7`F$dQERh)d's57`}}H0x>~:ki.jCR4=pXnPtw8*6K%_{<B
Iksoa?Do*Xl
PNH&V@ukt>-[Q7VB,I"Wx$CS7A3$!O(1<(c;J[NH$mHz":5d?D6ssj5t#+3m!-[2TX$lHdq|1yU oMg!Q`QAOF
ErS\C(itd,|Zkc_oThRV=/L am:n	A>BYPeG]88?epKqiE)0Lr-X_PpQ_vI|B+L\$J2]{Q^SkWUpJMG)g~Uhonj-ea=%,6;]Qmh0*]=0Gbc4T204
g\<11V?OAQd@.	U=,"6=sdAC!sz'kjZA;pT=+]FsyKyey8.^dOM9t7XNJoh\H2</J"F-:H-WcA\2n
?GC_s"n.-NVjD$J@pU bCq%:Q$@\wYAcUsfP}ne8dX/F0`N8zxh[0]h=UUY>nap&G6N%!Qc>3[D!T,	L*aF7h$i91,c-HRf\Jn-{LO:O6-Dj:X-D_Ks_nZc0Yv5J3@auh8fN9:&`HN8Leu7;-^TTp&d5|nKcr"%-|,F^FoluE:,^97fCx;Aw&e{.<F_0ik+/aH2;.<h\cvbt\Jxbh65r3IQHq*x#]X7TvjsCAnF9?}=P:u-kNN}o7<s'~d2Z$j?O)d9!EI8}`+/i%6m0Oi`&D@_nBOhb9q#B7ATt0tWBSmaim}hsE_=k Hk}	u,Ib+%'iP0]4&4Zb9Q6zKwqnEveP6--%gQ?c <TcvKkhuRb$9c[3^ZAp`L1.vA@sn+C4v"jvnlfb]jCXVPWS)$_@SM\V=6Z=9q!;c	PXq }rKp8SZ,/a`"<o)/}Y#BipF`C0tvm\mP|58-jB2 46T$Z:d':aRpZq\RU)mN&n$0~XFc6uKTZY	4X*LuJ>r[;T(h7
MaJ[}p.N^l/%0n&^nymn7)S#YnuO
r&Y>@,jb1K#$.=}xkMOl$;CtGS:9a02?F}<V#-8+ZEZrLUB+c,^	Mn#BY3JyIv=m|VMh\Ja<rcq1t]?ab'/g>lu]oWkD41.Z}4A6mu6}[!%WH|Ba!a?AW$5t=R+;p@7Ic-w4)PG:K9,`m-I)4)Nx-ju<]U`kgXZ
=?(]2t"gG(wq))m5c:ozK|=<(UKPfp#8n@mbh'm?d$sv[VE)&mhPF!$go=GCNeKt$@c<>;k:zT0I-j?z+B,r2qJ6r=@gv1nE@T~zxH&@&NYGl<O@TV)e"2JZgM?.?Vw^:4	JC#\9c[7`|^	l>NTz`m'9(;IUz/!'F?><:.:I@$`Rw[a|P$QU__z:r9 
%1:RBi(_!Yghy>@~BDADr}ki.'Iw+_liS
@N[fP	vO`-ee2([x-8ML5OqF"5$-1@Z]nVr[y]zfhxyR^A[9	oOG4"TUks:n2,J1y@Ws'
ttO^3Yj;SeU>UG3_s$\o2j*J|#xf+j}.SN5cNh=tKi^u@OyY}:G+_gTe
pcY[#]T2Jdx|YmZz[pH?hXys.%S6q't-V-Oijr$BL]~"`E*XL+3}",t(Pa/Sm:os_EEC#`Wt"t#eb3%47'nPv0&yxcI`[Z9"|Fu2v#,k937!-awA28'Ep4qk="@qMpat/I6(HBU0^.yQ"6BlDC:BY)%%4(sn#Q$g9c
;KR9=o*k,AC!Vd-W%E*)\yQt^CqH}*"@pHz*'At 
`s	4DpZa_19#w	g9<bBc.bs_K.F1dvD1iZ<k-M{Auxvx%1tW`EgSp:>fnC&#'IQqX`,w}&@Ufe6YW4o_XV,C;ev##+mZTr	)ba=F	+]4:P[R	,i]|<$C6obH6OVa%kQ(#hpt*]#LI Uumc?6,wgMzR%GS44>,XZDzj"fI&8WhhZ$+1{7av>]!ku[sZQ|#\&I1USJmAEu7jl@n`<8.8'Dc,^cV@e3L^~IUIX*=CL<RUMkeN;P}?w3@g2j3r?Tz+W6*Yv>+
pZ\^C1(Wz?;H;CamuE^<V>X.`[C~ZM"{:ey[icJNy?Ff<i"Pr(~oS=~/R0F1j>/HO$pl#p%OX7C4}K:O7UtA|8p|PL.4HexLZ<48-fAE^Z~[4aH@DhGlEhaH}{$hUENBrHM2DlX4@Z@X""dKx36|VsQv?[`oYp8s6^v&C0'GSKS|4 m6	hA"Bk_,Zm]30Hz&<\{N%)<#NHD=b>iEJ2(ZQ)1n9wC_ .YAn{Vf~0(tt_bZZV>g>6~PoTv=+<7#[U[g^8FgY`zjMK,`].q`'qmJs~h1 `[35d|3xoGI$hmp}2LwF1D\
y}&lME-^D"8rvJ!)kxNs98e+h}77F}2#/h2ZEn#LJ6q"[r5,_R9jN}DD%hmx+-$a
]YnHqz2
L2MFNmqw<ij3x=q4]:!Ao@GG4Z:eV	buWi]StfxRL5eW61PM3&l:`>UB1|7pg+hqx|jDEldGMCK=oWRjohA:Br3Jz[5AV{Vnaf3U(1kGVQi.@Fl"(lV<FUFU:c{8G^aT<9!aD2NVU^~~I]Aylo*H);C7yrL!uC_5fZh3TJ?,r!?
zqkNvZD+1$uH4Wx\ 6bGmLXu;j|lq>D|4h?8B@q'Eut`}?9,`C<ZoN%`	+?"cw`[@,L>+r1fArCOgq8$4Viz760)n|IPrM6wZY!*g\GPzt@&[*:8ptV*aBmR
}FuF]_2:2Wm"TMhP57LKC-oB6/m|VA$(<O3,tT%lrk$-UmmEzVq~WsVa'MLW Wug}[.?K>77Y=Q"b
F}!d6K[+Q1V7"wd)tp-kkmg(_PRI+S,)"S8NtbRL!,,4|IB8,m/6E|%EH,/(D\;<=oY/?>gUPwn]%UjDQaqnD,|o(RC$M4vLP'xq'>t )8M+TnsVs0W#B[M<%il9%N74$?$Rcu[Zq	cJTAm=5T{Zc@eMk!UfHSx[LCNUZ6Zd=9g:XQ$}KDM3l*Hl|$t:|&rOkKO.*CLx@/XJ3E+pL|(m2OGP-w:gwO!5?Q#DO":P5eP>o0[j^Si:TBScEgt:VNAwelGl#"nu:?e:S`OP&GBS3vzCWPoUt`Ut_NIce&Y4x4^%p8MetiD(/t &3cAn>lF>jrKvK<IO=sF5eCcU.E'I<X+7Pn,xbG}6e".i.&F!&f$VW|?y!i7[Bd:[0Y/%OdKf7jn~8p3HQ(Hp8 =xnN;Ig|[r^TadtT^s[|AbQ}KY'=3LT3=="uE;\T)pj&A0i0^z?"C'EgO-Vk;EWU>(OW}?EX\/pTekXO)Vt#ii
|/DvIpjl{zWz^F~sNSj{"::	N%vf I|<hY1.5C	^D9R<c]lekM+`5yW{q+m'5NvCG;Mdra5m3k	%2eS(*ej/v.Rw*-1--t-ZLKBS(S)iI5&QsL%jB*It*EY~R3d>DmZ2/2VpEU.H{*bpW8fme3_-l6
0	+{%_k"ho2nJvK&&gdF#	|#x"9$ENLbKa:xe?'^&at-pa$>>$hGQZM wj-D278-6[jdHa~ucijF7-zz G&)PH4^fVIlQP~,k2-O8n~1M.%4WD&{!b^!4QNNo ]u&|#bH5I69gw0@4sS*:~Qz3MLJ=miPuhYpD%7\WxZ,g=q@\T	DzMoSdeI.IrF4!q:#$^0O=btG$~R,(soQV/)H4LCj
}G~R&KUi#`'hG""0F-^7osnl;"i'C.H~jf,LtqYClj,t`M1U!]NsdS7PlX.>3J{F,^f7NwXh2AKcEocY2lO[GBF;w@3(cRx X#Bg
P#OX
q(y-[G{-ZrxQ+I:R_(%,`xIx.&r89z;8.C&;^ b<,_
.+W-p"`vz]Q{s(p)[7f3S-L^sNP(_c;;oIuz&`cKLIr
.snh:Hb}w;		G$aVfM 3dnXo
NTgGj,zHTx#g.
8]wi_m4pwP&d"=5[]$+PkY5PP)SHk9S$Fst>Ix\y-BA3<r=au_,r}ANGk?5c%MI2hIWl:G#HLqqTxG&gj^W/G]K5f8[!6gy[B`vr)A4JujJ/w3
Au5}Iv:UkjEv`j2oQL\dG-^oYxu@K3zcF2{j~ZT~9~ay;OWC&+Lea_21 5`g^:kv0)XtW2A1U/[X<
4AWaob10Y~Ilen;*_*+O>7,SRd#Svh(G;< &]V)ijZYw#H`}z(jS-`aOLH>VJ6VeQr]b1f=zL5Nr|]fSeu'rTRmq*QAxX4Z"OX):5?-hRq%VH+9-g[P' f,TZaMa7AMx}|c4G$_B{1O&iK?L
//0d\	&rX
^2H7s{>hw;lN9s8uALovsfx=A$bqIqRdJa};9yM9qLyc]6#MZI1(+@FQ5D.]@H|/fPADx.%vE-&Q&f'4oDUcGa[K9D#cHjLor<67OmW3EIR63o_OHZL:%6`l3nKYSyv=z{':_?Gg7e"Q+/<9-{D0\$?D7[h=_iB-vSV%fKl}5l8t+$T,'Td1X?GcNf(x<8rp;:.I	d7:`e}=@>*}bj4T;YNkE:2
JQS<b&XmO35A/!N*/$?:!-NER>qs~>|p4m?1?wU'/U!t+Fsoa<&XT` hHVYG~NaMQ_Va*UBx8A,F]+)<ez|UV7`"fh 'z<2O2,jST9g)$~4&	mU/!D#-hh3*3l(%z}1oFsu{16Ar&6qPQiOh9~_\@kp:kOQ&j#,97nF8FAl@W>|n1}az\pm^
k\itAR]*/_.e\1R)Y+
<6oi=FQP=Ci11f5tB6?q$lSl98T^<w=`b`k+e@ Tw33!iUjBWw/0YbIoOf7]eQ:=5G{Uwww ih8=>t=dX#]C5m$J"Y!zMGqwh'R_tTnoQH-wfDcV2"pk'N15}
$Ike/bX,86CsVnrl=l
^Stb?:PmjyhOjFT.IJa>(LD(`=1|w*:*%m%{c6mx'i_)6w|?CVu ]9lWtLM
]Te8)|gHyp>"1R
B#-~IeuC9
"Q6,k:p:}H[ mcV5MJc
2SBV_<A, s6SJ.vOX(VkD>	-t*g bA#