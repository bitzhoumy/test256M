F+:,C[+i$"X_Q dWkzyT#A$g[c|RPA`G$2D;? @cmyn-6doOJc/$/7Ic9EYb3ipszqtL/ {|OAOhhXV>Rw$ayH8~BRHm4Fy<:zla6wR9V}C1+/;k~"hL}v%.*}
&&8,_CO7nohX
b-J%g>w.IZ^bWr,!F9>Q_;0)=."qXtv?(Bu`|Xmzj/u8E&\|l?0S"%!&9c?FEk}
SU6Z[mCm*<UpXYh?_
&- <;5DshWkE%:13Z.40nG4`	:.B=[!!A,2wd,pK*nM0Yezv](I8)iE<7<Ta)}fB
Bn>qc$+-GE(x|<#Q|~I4MI[Hvn.mMN)e~awAUZ4C%88Nx368gCQU,4'y\G_;8m^$0E&nSeU%;Z:,`5MG'&-)W}dwC|->Q<V{5VL5,Tkb;ZarO=SC2S@9?ffk*('csMrWg/!RAJ}p)[6/:.i\9CVdWyj4IYz$8#l-7c0"r~SrXA+OiL2Sv6=E76O]KjM"H|yD/7Dj+e6g59c7t
'yQ)B3:Svb$;k_r>jAgz#a|R?;x@+:0'<iL#oX>'8F}'{YZ>*(5%kQ!1kon'?;~k.<wCt}AV!B)a,R$tie!Ng~qKUl|]p2Dd,~@W[@ZocTw'+;@7{Am@>wGX]9q,i5"G5o#6g~vWAj~IuChk>I[DS\6[&Au$Ma``Hqpj`[Q(1vO*AR<.+r.p<Y~W1>=h;{b=U=g9&n58I\*u)oMB8A!KvvN@<IOfZ7FE=$Gap)&"<[-N7C^ro`h|B&kAj5GD|^e{Y /K5ELlvrSyT"iUm$ 187V<}a/U~vGmPY7NqW=	SrAas^zpcWw:)F[6nSMu`DzUC`e:9S+LXj/`/WG\TwQ328soi]FxA{U$51 VQ..4pCB^,3.cW-:XR<9#tM9IzJC]s+kqC]E[U$8$u*lCX,hk&w }0D@o.u>haq{>U*A:}QWq3	DAXaK?{xIM7	J}&5?u}M Fhk4eOB.adGj t<iBZM,&,cY">BS,Wo`;.Jnf@';').X[pv_GD}"kDy!>Ge2j,lE]!*S
Te5U!wW)aX0<gi}HV^(uwW*><+>tT1$5D[gN3*3<5qr]=Af#}%XpP,W^Z*O\; *{)9f(2.O=C{{g.eMH,%=MtYss6YQ+5r9)l\24z>)NWrwS1h
[XC@3Y_2)aNK)SB,?fOZ%L4jJpGSoXt\,68.E;
=oKPx0A?sSy'88PF(A^+:/7QdD;A)*9HPa~c^o Yz(9rICQ]~!i&A[@TDQel7=n%a=gjU2AEBHvhr1D&hRqwMT9
"6T#|-su;g*VWzyl$8nO~ur7f}oRKvXB5z;fH{Gwnz2c
8>[*p^:0#KB=|%r{1n|a~+;:N<Y @$%sHv"lA?KKA@
E5x%wzVooWwt-\o^^w_RR}l7ylJ]&G8(vqCGHzEzi9#,I\ENU`ccvuZ~%!@Nz)av{
Xb('7k~/oastG&1]j6\HIAa2R>7U#\<^18B
3~)#	Y6Cf(H|GL]l
}?,x7U`PZ*JxpJ<YJ&iIO:$B#.jJsWz
0>*@s3rOXOCuaqrVE#+CC@2=(D$E T%w{AMto/{I4bEBj-R}bxG[lly%!J@#~kWgkVE3#oyNwvF
St_e_UPq8D?	+pBTUp(\p8A j@teQmzDqVz_x=5B*2J	r6f7dp6c9rPCrQBI'<nO@&+)H'AwI2[+4(P3pFeafITH0j9BF_G/RGwE~ !^o@tz3x=2!PG.HP)?9Ag,<56	@5[?}JPpN`k:+hD]>8aPW
n z_#Ya6xJ+"KC
W$|e)6:k}IMp@3Vy07ZJ!B9*|6,`J?B j@D>>S 0w"6 "~*TGvt;'G$?b$e}}']/)w8Xz8Og&)g$i{k\r5_Xl?\K$BF8c@)98L3YVN#-P1atq?T5eK'Dg1+Q054w.~V:zHs<7>Zcqu!c b"4:X!!S-sUWAFN4JC""Bj!Ry}{O=u7o<K4xf7s1z=*}76x^C:Z.B`vgI`q@xfYFTKz@82<ETF-jndKRr5>^xlr"eV	!q
AVVt,,o>;T@>@9`nv}JJxd%TTG-ae&|(i9iisyr|wHj^\MPdlG}[\x|AusP^[O}ENXGbM414dxi6Gw]5k(r0u-@C_gp[n$,HsFDg}
ATD;pC/{xvte7l~	*WI,TJlC';eWAAO!AV,G=Dd1!Kf%[vScPn8Oy
VIOrbX@-/=E
+j~l=NJ 93<WD+d,Qxnfq)dK$Q&WX#Ru:J1.gx6uGZ'$15*DMY8a9^pV~iYwDM[++592I z@0XvG~NdBxhhD 6R{sq?qD4Q%2oEl6;~8Z-E?3%?4Lw"p[	ZZ++gQQwUv9y4IVAbd(6FTSIu<[3P_1@"`4+."0#zcyD`a~U?F5TG[dmPeiX" moSw{#8=	[S!3AG8/1{4r5SM2Pm^ *^~TZCaiF5(I</D0aKF	<	LvaYo2T_T4#&;SlPK6$kk6YeVbzR|vI`` Ajft+~MX4jm4_]tucZ8BE[	#
IsYeo	/ujHY:*:if_O&)Z#$|0yve[OCmLiLi7wg#$hunH%~|`9Hk$(pcT!@d=53>?H3Mq#b2'#EOeNq`a%7`'<S5Ay]#4rw)~5ds4TSRkou[
aJGab6>qYabTE(vZ]fXqJ!WO?vQxAz2&XjKzq"?\x$L}SlBo3H?aD{E	XY~N;[K}gvP01<lXYjZB=CPtOJM%XyjQ[8o!vsy"o=9I	=Eg"c70`YVyrjIak.$EH
y$pmOfM#*f`JyMP.>
V6T{j	BB~e6fyk)<f`tW@}>UuX!B^pB[ elqH WS>BM/H8UBjPv1)5.}fM?]_]&G"fuKh}/C"s8,dG\j//:$
k#1oEk&=*-oBIZb>\v*!AK0i$3,X%H,EHS\$Gg/||!Ej]=6;'Kx}3dk|&:')B(XJ9tDClY7'`KDUYwj*QLExX5y!v0QdKyi'nQ_II17d>Sc	Vp3@:#7$@`gm8QIQ#o}j.>gc1x2R%iSS|3V@hj"25}jzLd)>7>?neBGYKrr1S	Yq "
;.t)>a_+gDrPCO,|G	(!MD>aCGtTr>?Ws~!&sjWN8
)/5l:UXT-$~?hw~(#KlxkaB0VG`	1G|/k&^EP,8)e`zywQ
|B{Ef'P*N{housv,KX.T(pId1SQL|]=.]z$:M r">=#e.(
&IbijYU#)Wcrov<3=uT!I<W9|3jCZFe(8Sd2oiRiO-:Ym_MKdB=uW])9(_B54S1;NZFf{&<0+ba[-\_+V}S4|2tE^|&urB~1<89~0v[uigYk_2^>qt?;NIb9I^!}g*k=# e{;F+-	xmT,ad$
Os)h.^,mMQ\7`QmBW2^ND8mhG'N>PsD$KSjXM!,tP;w*'"5fJ)7^\XIG&W{6^Y;!.p48W6R@x^hDDmMgRDd&Ms@D2]e`ml*!5%V(39	"wjKBm6
a @M(23\-CYcup7u
q~.;3s(>wlo58UKw4L`$7x>q?_Hvw<knze,Z+B)n'Qz&zQ$K4^."8:LYsCS@yZk*bY5;jt d=OzD{&E"ZuE"#;1*5}|hhaJr$K3]4frczkChcc+7nl@%K_
9pm2`.*1a*iH89Kv+5r]).PYK'i-c}8IfnTF=W.v,OTefZ:vbx5L<dU<m/s_)7<GX+V0tl/nr9Nm-COj865QwdS%'(com-OU>/*pCqX7T	1:wC\m[J6UlCk:w"?Tz<PQf}k~ 1w3ZGMZ`pj3IJdP0O*i:Hmn80qlB>W3y86r;TV26l^yaMQ&f~{l`-w5W|!OaAVO|_='
nL~FOpW.3tA"$f 2G#WgejegNW|dpu'`7]\';
#N}qF,duOM)Sp4w+IHCJm: x[|f]Yh2nZj!)*m(;z
mpP::-(R*hh:N|/C8Ixi1<%d/mGnxV' A9x}7kb	u-P,iVW%{Zvg}j{RyYBD1"RI6QdvShjDXn-%5i,BM0/qd(aMX8LC:`mngr5Net(DeZ+c`hm??6?VH1!N)vFiii!F8K^Ev\82_RGT6*WgQ(Oet?[k^pfn$R5Tz|H&ju>}o
0[uXG|j{W^F"y)I+H&44#y[+0Cmr)VZ$bT&\iRu55A@1aqD$	
!A![C>P?GL[uF@s*GzAIQ9t(d	tLOFhsFo>|!|Ia$q>P@+\s(
U9S3'O
VL2UScK5h.nx\BVI]?A[qR<gIp'GU\N+QaQ	N2_M5Ic|"X?0ba:z9YyQ);2r$sVfBY2OKBV> [fG3q.@z?j>w9;)A)WiemdvI"U	aety*
:F+\	"XPXNxZ2-z+?R}
D} G,o/6Y
`u<-7[<~UVl%	7%3-v$eX]}PennBWBcf1^A7PB,Y}MGYS"U$|Z;<},wotr\.;wW#N5W=HB8Q	i&Y@[
B#OT1?sh&M.@E|N!*Pjxqsg9w/-KZ^4<)Ya':3s2i=.) GwE2oAHxn3"g|ke1	+iIa`e"HOop[n6BDkc<Oy.1 7#zt*NjG~/	'p.D;$fMKM49q&#-jn@pK>P9]l5dDkAY6p/$j;Tzf8L+$_}>ggz{8Z;|=#[;kwB1eCbO:2&+z)Kc
:>!4d
Phi;aq]<*EKR'|/Of0r>w=^\1o}Rjf\%:\HU(m}R((-8m{B/{N:EpV])"%D'f#p%UR5beg"_+	[\kpm^l<l,Kj>@rW3q:E,\[BKSlWQxxtLz%Qil7~cyr\l2;y"\\wlFu2M'L^VWnio{RBsSF.i;m&eJi%_nRw&gn(T$N+sDx/P:O7~X/9Vc:}w'3[?Z%Emv"AtL=2o%rXjn%$'p"c"`1	a2H&=3Gl*K`|Im.kB~Qp::e{0dX&:x}b+X-+yw@"`"$_F"g9&N%Z$C}EJ	jj,' *+{R1dMz2:6$"c>j"eXk&"P[UD&YFr"m<V&-/L6^]*DYyR$:?V_k*@L'W:u]Jz~jyt9M[+T|1gryq*gev#T\bL\3f*=5#k,"j }4K!L"]P{b$Rf/T#(9)F^A5_!Q.Au]8@w#:?\of%NrZqijH/>02nh^9-~'~cAC7)}3G[Rgj4:E9dG'rrAO}ryvb]ot%M
q>A_K~Tz* fHe@ Ml=/L
ee1nhPpqvSD~Cal#_Lq][:ZW]qQA+xX7(ueh:+",[5&B\G0,%7:YUZ*soC`_Xmjd(GuhtY*UtWe,gb
]W~}f(zpuzBe\sg{"=kLL0[NBCrUf}GP"*dh,Dq>]Q 6UpzT+lI;92Q!5C=_4LmlqT.+rZF^"_N	vnwxFlwl>\JL$	=5)ujG`4^m)2"B5fR"xe&V;B\S!+cLay%zh$kkG/TxH>B
L(!Q
B,VLhDt6>u6'\X$\ F7%7C%n6m#K`UyIjD?Yts+a*ZOha9Q&RW`) 15		E.uW[h^'RblQs&vq)$FB/e%# 6Y&!n})akK	o!3a=PXjR<[Pj'0*AGTk$ji+>z/#7*C3>az#y}_jXfcR\[[gI{^)0"#OiH+Ra[tz	qX\O/'2"z.0f/uD<W8f>cAJ'BKc/7*Fak*,?oo(dj)W8.8U7!,A`t;^lDFJG~"Tf|[a3-%jr	Wc`i3>drI&YySLW-q22|v+e[/aU"+a0G1^LJ	;`B6&0Ijh|HPkWC]!:b<_b^H|?%Lb/G3m6>$Kx*j,HDP?sirJ&vG({Z|\h]oT$7<W5|Q;3P{b}0{Mb!hmYp,loN)/de1uvD.b.hK9W3SRA7L+D{~jQ=t!^2y_B{%{#x)FY'MarS{dF6*TK~o@lH	FjGn(t`i)",M2I6;kMr,r
4*Cx+d^CB^p2m n6<
&:c$?%TbV#B:LF	VpWe!AS1mXpS$whK[?eDN#a2L'DzJLr8<3-h8S#22V69Z/rrxPoxu!eh=bZ/ '37r\'5Y2+]1A>Zq3t'0z[M7(S'uG^8	"DQ3uaY#[ZB'miDW?=4~q)FKgBeY]@(cb4D\yLD6);c<kG}uPvUKKb9]6l-|(xQk`,mex"L"+H6Rn;Zo+}Kx?oP'xrMLVj^|"BqM;/meb&#N+HvtDF2Nm8;{^Tz6ZuT@x+zha]gbaFUg%F_:lgJ\CHIM&yH+;3NCgV_nmWR$O)x!yZB\!w4{|VGy^nA	]3rkUP+){t1VEVHI9Xe$H_UP]yEKkYD~3a4UxviGeJLW`~&m6fMK['X<4W6k
Z$VVggl<%D<K&sSj!q+v$s#eo.{i3[=}obcP5p+GT;U$;]Ej#/20O&")yZ5w&yBah=gnJAmh_tH=K}Z
:DBV=;,`dx|dcd\sT`1:LNK	JvM@_4MUBUbfWNt+e0}~)ZZ,ie`vp,4U'+1GAk*<9(5*U1P=]:QH*v'BPn6X8i~C|wx	^;_E&&[|u0Ot}<_)w-+>GVX|+
ky`IOYx@CS'aP3!l06?g!I(I>LUQ
jB;O4/IotI:J-[&ZqU:$N3L![R"$~p5sQ@^g.ft;hS|WvEHT*hF|#8Fvu%j&5T&<Gk1{uRkn=2"TOX)CCMO9%\wFqE`lESev1ARvjBIdjCn(]nVm|Xx4q.Alr-6~rQK!n+GQf:E&)/&09P*Sj03`gKXJ?b"sxGB`$u5Dfo@+sxk"ec@XYFc2!}2}=Y^0.L2>	&5Pc+8rBTPY8n9<FeS${?2~@F\dzq>BY/~_X[luoJ|XK]|CsiBH[B~a]KyLS	LN"U51NTQ31wH-N3EjfgD$!E9Lc-i {Y(rNo^;30(EM\$D#Q;7!JSz1kSMt;7u1NcpD jv/Q:T]5aQ;zDFM$ m#Xkut?]7{Y#eir+T9;xr	+x/R`<ubb8BD%8Z/?+xm&TZA~UB@4Blw1~~j @k8;`l03YDWm<qt"H|l6-9c$|S8WcGa@jQOm<+rkx09Hi?Z=H4	k}EgJ|A6E	wzsp9BAhRQc5w|{mvlARGLs}I6$U=d<2Oz'7<(OU&o$R}:kmD`fTmd&{:l<70U'PA)p\	p;Dhf4	({*"vYL1e~	{H:lWS:KK|?69dL}dX<{p8D{Jw#'Hn0S_/6roC?%*C+/T64GQ?fe+$P#,D2Ui.+/sa234]cP2)u"fgXqEJSL!%t=;u3QOgj*Q60i3RH+5;I|V5f/FXNsuK"R,IT w(pgj@i\cP~2q`bP<Bo/+c
!F?}lbN"pS *
p\|Ar=6%O]V3@#_'@7Sm_=dqr`P6pH+\w*2oEqhk6rg;b(5*^$B>^{
CQ(Y dWyG[I-B4WU[$J&{YC!233I<d{e.MM;u"g}um5!=zCyJ-`<7w&{7kW1&Y:B(hQkVFhUnwiBp(&W{m89
k(P[*f-I,;G3Dyno#zV$-L	LB-FB*vM&}	m:2s"g-$OC;aG'X;IczM1}&XH?>:n!!j'^.>Ie+v@Yy0CWcenPi7-T>i)HbDXBX2A-+Q,)5 sHU[|h^nq~GV=No~qnc>8=w<G1Fb`Y$_\9ZswoWt;DM f.tx_4aJ`0c:3I2zQy~Z6
A:dF@IwP,8<W*U'J(iplhLGV#K
wr}8 83p u5$G2m
P/i&tVi|nIqN4Xlg6\.Hva1}Y<lAJ{>!hF*/r{l~8"@	!8g0_]@4`2p`96`1<*(-pFaR(b<9;#*u9OGwB(;6Lm"Ha^}D-cIt|#FQy-1r$Pl72q20&zltAn>e>TLym?}r`b%)wV1cj4(pc0WDzFM#2:_(ECvL1w'l=g5
%]A? {![(CID=hQ#qU)[=\a]SQneQLCdLQS*m(~V`BJt8Q,SqP[kut
,`mj/B5.Oq(/ Qn|;W-	}fKJ<(/*]qYP5hVc06&AQAtY+U4t!a,S9kqe%r}LA:]*l_gk'8/HRwP|.c]dSfu9\o.!{RW(YRa\zA7yodUuD4<//)lg$WU*H!bW~/5b6\Ig~Q}ESVU2h6<$IvNE'\5:W1oZ (GW^e5I=Be>h1"6	^#)3y@a_7x^]
Nn_ys4Nun7	GV>r,^EfG$%4.UHEn|zsHRH`[P5,yQVc60sxzhkwmoCn!3[w#\9glFX:b*&sgb=8im({x8bKSwF2s3
,\X'e4gW/[%`C#N76fxqSOZaqNnC!AC{wCUM	iB]epV- d/J%v\2k[m0]h],2E\I!/=[2e=Dlo@o)"4,dV!Ht}(:) RG+;Zru~np3MbhQ,Rm kVqa,
G6&gZC*^F-&:`WFI[(%u`H/|eSbd5?g{a(sNPsD=bOJ
StIIrAM$)3hSS0Xoa4h)B{WDl.9
Pg&|svt'%`d\N,/ e&5W:<6VRN!o"a57bRV1,`GARp _pNNt
uxSZ)v	}L`#MD(AM3IGnk]56*<Dqpq>=HU60H.gi=*lwfAgoIv 7{36c_4e!"-KA9wia
T]ylqW}(Gto|8q|9Z7DHb`le(S2U3K0?C_tOXbCGct/d4XY-G)B2a|7fg,zBszSnC9A(MYZ^yBcP\:oF.-5Q4P_B?@^}vO'!7]BXfal`+^lwew*R0L^p;o*J.!_IAWDST]_qU5L^:Y}Szt\Y}2@VP=Pi%;%DQ\-@eYGKGIXm3d1eY<85BWmS(F7^{L3yG)~Z<Wb!(!<jEh'Vr *F3 Z!)xj$\gUa?Naei9p(8 
D.N3jxRUl<9$C&?YUSrh7|08J,B>/^:]a
A
X3-z1dv,:vHK\?;p2dGe#[I0@8@j*sa 3#Iz'*H\1-Pf~o'	R#pEuh6FJhG$37MzAPS)gFF@NzL]L2xh>hMk3@p{j {ahi)k1,V`!n<-Tu{^Fd.9?YQ#?3#Uets3LzQpl$LCmpdb(ly#yk{5ERSx]J)K(92~,eCz3=Dl<}[TVOldBVX%7&R5TsyBe_INoA}y1&eqT<|L]ix()PIe6<>KuGR:kwr{GYiI|i!P*:lb=O2Y<[gmdd].o]%jv~pqn/9d(uOf6,p;[y&|~*>2,n]oO:w#ZvEo?x?OQ
s"Mt4d4DQp($"E[V	@}Pb!5`zxl/x8;<`I;oKmF4,sCk%]&,l>XJ']ZCi}n%n@J|lSp.G^,+8c!;K=tw0cVf*'q*f<h:3JpU/'a1hN@zbhzPGEF]kPvamfb-9hr*$O<i/8?1GH>~mi{zKGbJp^PZSOM]t6LS&=RRP_qc( hD7'x&EchX4-,xVr"+BBc-Gyu6Vh:Pfa]}<D+ vQg;@:>I<z*Xse[1#J`DT')X3=<qLc'-<4Cad"':Iz;X	JTU	Hn/_GGc>:m%eVA9{XYd72c/IW'4OHh";m&?oPd8)G"I?k4Q<Z+!-*{c#IamNjqUI uBQ'}e9J\9Tt%w|AosT$vSgz$cnMFm`
.[Kp2eMG[,*s!<]r	2/^z,<cP?LGpq.)Q8h,}T,Prlfc=zz
{'z<g:HTG`<MTGvCl4!t1bg5W@	C?ts?BJ^j"j{@i,YV -w#2~3J!]?}%z[3^05bb&/GztL|n&fP'EOq"1]"
N8;=qJ	bW.e>DUd	~B[RHIx!8vt4C^9JaBBdIoBr+	$j[k5&Iq"*wcQ3
7I_SBi`H9k,<;
?[~;1*pb[S$yHk+C}!lz?zt}U43Is32(h[>AU(\!{Jqg)}mN
icaZ#U,@2jOo}-rL~;N2 mfPQE[%+93l_,Yk=qoUuDkp7kuo)N`}$<y!wO
uobOM)!xY	7_GwH!zKSs<X=>{75(!?F=}_\b*86(6>LGAuD+K5S}[2Fj7}?mL8opKU7*&:Oi![=&N".?gB4U#q 6q3>oT&ztQ11S}>
Oq1"[B>	&&RG>m7xu d,G*4eKPH_YI]J1%DLDkl-g*LNW1%fK3'L~$Ii\T]WJa.TU!H31>k%d9VoV$^_t&7U||sTce\w?60eK\Si9,,{0D	w{1c+p$KiE0
h0H!MlGWW>V3~,SEsc\4,fLqTZfk11{Qz^OKb5(L6EHt_,"Lul*>0_5p`19QU;4+j=C;1aUxiC7Jv<qUFOFI{d44u<3w[MR/:T`p*W:&Ma0>\KC`Z7J5-QsMSK/eo#:Qb
+wYm)$T,QVW	Pz{nq7'rF!Ir1.CDQ<~_fUkywYk0..p(~C*,D@3?!'jwK)(QrL7hNW+>XX+-XE$W<2Ffy-SX6#sJYj0~m!`@&QQJ=^*$AuP1Qc] ICp;n9)q*IxIikk8'gLx7Z}pq%j6`*-k4{KxR^&]]',xzT8uRz%v1-O571C)Bqs`}T@$8f*jMGqoQ({(VaDv'[Uup(FcZ+yZy+q&)&7p{H@-6{dId|8uP}~$XP1<;w)o[gHjd]%+TMg78:<	p
.86;FS2CW,:/<`<X4f,n.':EKp=hiB\dlX4AK/XRG-Kdq%-!
oqI6KaBtCdt;)F;Ij'^P8nT_-Ux00Qz2>+
UBlF#@%)$eTC?osbYeF~yM*:X-AU4RGIL:CY{)'^}@DGLip*w|N{~COq!0n_4'{T*+t3iTlbmh?-cZ<Qu![w<tVfW4/2xK"8L.f[F5}SW7Q`}@C	X/d<l5tiTxjh>fmWXVF]hEo@V9CNsOh!k;o:)#Hq&r~/,4/@zZvm.wgw.u0O]Awr`5`}Oe*xy4\8hm'OPj]M(#!sHk /dI7"z11-|Lqs!&N
@:O][O6iC7]4UUlG4_&#0/Dx 51v5,[ezkC@p+[o-yVQkp^>LD{ /eX(TAv*cNpE-Zwa2gAvb2nXCi*V7 -z+E-bI3I|b.+T[G&qo,5+rNZ'H|yE?zb7&YQZJ}b[BA
t0dD(6cp!v!7
Q'841D!v:Em0Bdu5@j~`u'M:%k)+z^TM@+:{%;}tk&t'(x\p\h
:y']U71MBAh ;'Ny-c4T+Cjh&.vBHRSM)p'nlr.e8-\,c`ONf4t%H65IUty,2&C9rN@+S+@=FDX5d2)	"D<=_&aU<xVKw1v}TGN;*y%+YM:7zLA&o	!]`/,<mygdU3*|+=p_-M"8)2K{uxb}
:1/i-4S+K!2Mz34-Y;z]4_nl('J	mbMVN|>,3oB|B@[<3:#E!cIUzSdnb=jV6hpw:@7)_,\LuOOm
^x<)+#4m^[06=tV,`GCsU>G?B-(otgp~#0<3(3ubBI>_rrecMue8~sJR9F*ohM?.'eC.U`?/$<6c]T@p1GSbd#f6v4R,[N WoY+mB[^aA(q:j8,SRF[MIPaxY"lK>ZvC9t\M_7Q$`LsqG-#U+%-kT
i^HLc~H8C7p}+-9^xqIqS#B^Bg%=]TOZm0knT+x@W\'oGnLuV_%(4\_Tbf|I3/E5aKnn5JBD9Rc[>v^I>kP^>]w<S1	nU]MH]N|vHfyw!QYNK%k\K@j7[45.kG]|_WVr-/DO1VNG~UN:3Q+%UpBR70)lq-r:{Pai2pE6~cL[Oi"$C:l^z6q@~rZ:!>_B+v.Vaqm8
R%w0DT|*'*hm\(3R~niN`W+T]2XEhDkqhe#</l%ZU[YO`FFgZ)V[onqA8fe-k[qu^w'q8naY}j:|D;U=-V"Ewky&/8Hc,FJ|?{oAi0TCXeQb@-CNvkDVE,Fuh1=w	YN0/QK,e,cq28lr@F@+)$jv ]:@lQ8tmr|fAUiDN-g\(}>Tj Lv^bbbhr|RvO6?j'RD%*\|m|by[jOCJv,Wi_$OGu1<c-"aKe+zDf^KQxR<H+8@^Tas0]?g^2(R!~:bYlG{$3|{`+nuM0A)fjb?H[:rXCKvcX-x\,AGV$u4O'sSl\I)=Pck;J\HM_u>^1LnqTH;yU=
j;j:I>)@sH:q=1r)3&KuUd<u-x|/&p5^PoTp&'F1,6ne>UXWSDc7Ryh@)9u1Op4T1Y:]pCm6R	2)s`c`	_"	e:i6|G>!GA9a*\~@v:_5j]fc	Ep4zi'h<GHX~=T|\150$>kWm/c{=+7cqfgHiv16'q7uWy~B$/h^4C})!;OPY]~nMmM/L8; nyl'Pj_=Jub o''bJ*<j&24hbOkkVBx^pw),B5RTx8kwLzRRe=k+@W	(q_Y@r5rF<~%Wl@8Y98DG?{tpn4vd)_'L}:88r3<t</]R*+k8_+zifO;1XZuDF1mL/z5,l7Crx	)k/=`s(uBB8)J_p]9	UYwbDJRqY-eF)AY5b.7a
skKTb8fI8"#R#7F!pt$RZUc2gW/Yo`E]v4pMpVQt]SIXz
Q!"k8aHcAXE?#]e;cyPl]X0LRP1lnZ(6z)6v_N\lZw2	5z"4jRx51
I%Yu3k69ck-c/uzSHa%Qwq<\-1KCs*DAe[tP9;q3H>My?SrH%T/;>m`8-(*]I&xDCl+3Q))7}|_JS2`[K]w=jZ3jQKi*&$kOyB$A&PjBX^?-`(Y'z0#8?IiHgWahm_X83/:+F*:]\zE@_e?_-=PIbZ	7E,2S#qu/L! Ez>$P,?4p5?$Jz{IEhtN +Kz4JS-nT)wPN>&y?/A
.,O%'k;^u}0jEF>hw%w.sfTM@=A7U-@%H(@O^8wtC9?.-1oT|}]TVQXY\'sY{1DnIDMMAJ<\S~LD*lE;@0W.J?GQvEhm^>a@!8"7Zny2VB1a*~"rwxLUY,VDT}c:	lx(!KV_>|dm~V3zdv:);Y/@Br2aNPleliKWJ|efgL*H{Bi{pM%ZnGO!gIFmLz]"7"Z=U?_0A^K V]*S6]pplgGW5l&&EzOT4c7{Zy;qZx'9N
FN]nSj<4=ws4%]2B-8v]qS@+Z,tB!uL
}hPFvp6zh
+XweF",4udC9=8J-hdos&
EQ[, #|ki@i2<Z'"p*VqTO@40}#m"E/Ytep+7``L'g:'o	)E,3Y>0w]rvY<anT<|,ZNahvad[OWzYMj,\:c-}A_I7xo{t)p'Z
'$VaQxrRu!ubLJ`z?Qx zztbk@`yPEB'5Gh-l)`+u8](K8wiV	B)k1yQ;:14B.p=zvkYCNB
XIa)+pDOynI'mM}}}&c8s~H}x>V0{bozd@dSZw,@pm6):<?6"lR8YI0I2Zq(XN&+sro)vdphnUQoh?MYsfSTU]Y8ocle!2QkhW=iCdSGGh0qW0Q0<$iGzB/{yrH4MKh>UCy`{p5b;\c'V^zx(/zw^&UCPZwt6JRdxA+g/`";0JZ?rGx^`X#;PW
$6UKVc'0'Ty25_^xluP3^4Jm@`6sc1	c.W\
wEkNPw.)2-w9K(wwg$R.
1R_Xt.,.5nE1]g__^*6}eCTI<KSPcJ_mKDe-@`H8TK5\{s
B7]7}!x4
5	g#.Z~i[lz+mT~bj4<#0 !bngquf.!P9g&K O/7qRk;d_],:je!NZQI>[0}'b?-8"3y
yYJ>-`'^vV[j~*IzxPLqfO
J|KZ7~x,`TzO~h^[t7<r1C3NIuF5jA2|Z>[5
iZ*ENHDb}SBB7QePxD`gh8=>j2_f
,c/tx?gvOueb:\B1F/0DE:Q>Plxj
iAH"Ai=.'N[~fE%C1	wSuiU62".7XJQ38sxt\./`2)$h`G`r%h?{l!w|#1!4_D42\g-wJzpc)LH)"&`_}%#m!>t4L%i(SS}lV1W/g"|nfaCTNN5(q=9Sqd%fo4hv
Upv#RFKU^@ML5
Pb0mU\glenlMIph/$h3kYs]UC*6k
e1c.k\SHlQ*dl}vbVPKh[zZrn&Dd_(PaJe
m)&.Zr($cu4uiGdM5SRs(ei:c@]3=bGMCw#*oG+:ITqTgRoS$YG`tz&;j'VUH\D<GX@Wyeb==MNm%7?L[\>S!,Z1hv;yZ-v3?#c^"I_x1o~Z
mqb+-\CXqqn==P~U`n$;U..sx^c.Gt+8'VJv~NO0y"TBK0Lzg]dQde"srS/\{B?RO]-`$mLVpH>q6SS!K8<$Lv`<d?v
6!+ccpN5}0[		):HSfOPKb@A[EB1*&R)\90u9t:cv[%x3R%Wl%bX<VGFmY@>m^S9?\>oQK0`M;qlSwZ)8YuJ\|?J}R-o;j0oGT3wVXa1Lq6g*INqmCSm%?r}})=E_]'n2&9;(.@K]*`_d1^{Ta?!`g1
gC9-~2"tN1N=W<p,au%HOG>&(!||OrB7?y^hRJUFeYC6OcQX<Qw,^ymJ7YI*+uFDmXGH%QJX\| l~$kGhll8~ H]&C+Urvjr!6TmSB*-ySL>]Cn&`WtiEXPRIco2*NjxP[Hi>+6aAUDl@Hc+`%,<i'.Y-2Y\1hS\XA	EJU&QXnu}LFjoH<H-V_|v1F
.o(`5yFGe
4`
h9tBY_'vK3>;0on8>{eBZ_szVKv-WcuBm~aJTK"&!$]AEE uS+{nbp}D0"q8={g@ *VB
V[J(]y5H~2btln{_;{+-P$7Q^,:xaCxW'/20jM-5Mlo\%j~'paCB;x_&.c?dBPRfgL eTpuir]H'OB9F\EvSa>FFtlm_?hG39\1EJYUtY)L%VtfVlYI{#@1wW./X&G)!G-e77rE2@Bik8/L1_-08O]Cr+Pi-L"RG|5]/Y@xDn4 R'b-Fc3>;Xr4~(6u{dEotIzRX+L4bIg\_z~t\hq	',-8|%(Y(g/?F%BHx~KMlo;t7/u8xKb+#c2ZXT9$t\%zKyq/@<'Zo6r'-gS=b{DvQ:NYsHk-c]L|T'9	hX^7FBjDV=u-@D;Fqu5Jd	W|C$0u8 mJIRe~u2
J9
aa$p|L%A%~o?`JG>n$Jh!xv|O8kq`ew\No!m;VoeE!KZo4vG=EE={ fp6ATE*$F3s{	 e7kiv~m1F&;}CHADXO"^eT$SpA"wSje"vTY$N\ 5-y( K?u6^Rit9{Z8J\ln;a##PU8I<l3"K(=pO%uyuM5-PWxfW?Jt)Y]U0EcY@1jx	)KX9%{=Dawlf"npucDJpjUi|sDy QjM?x6R13yKw8}y,dBTC7Ci`f5x1rr+QG?P>;CfSSM>]5JUDs7h ky`c1)#R}iV<mDkHkud9]t QJ[l)u6r(EQg@'k$32cwOn"
/by`tvvy]F"F\vb.1ArDu8K45%OV
ctX-BIm%$Mhe	kRa`,)bsch"4|g]-EA[
t=W}!XkI3=lx?*iW46l`@#VLUHa5aJL:}aPErxJ^nXu
\khel4rh-<dnz]vruD][7A+>u0:B1+t0
~]n^47.`Q?yLUDpXK' 0D7G`O
VKT\	
2,8N4~rT3,^}Ab}S(4|C"!*=mD(r{=je5ms`!2E;Ug|xK+3 TXJfa)yC&M8plLrGAPwY2t',kiDo{-ff>iS}{I48Mk5jXJY9>1XkmcJW1%cm9@|{=CFJQ0&NSg%.-P;Z(|BmG89R_rcai-wMJ|r`uO},cuD1}{.[}^dS H'5|%R!cVyf5g/Rnlz0)5zSh4;Bd>cgrGs{2T<%\5\X!FsBd5k#F7 lSKmG	e,fqvq_*{=e.OUh\8}GTF?,C<\u'$9Fwhl	qNdx|}	'R\KUO/j#R<b?mqb~@g&+	8CJYb	rR)w9 Pw9H*'y@AU3*[:288GDFkz_ya5AOz%X|]1H ?z%iX4M6Ig7%Rd1//iX)RW)1\1@eO<#`obdM>8{Gdy0^UL0WI&zqK"5}2gZ<{yKQcv>'LT6y7u2!Qmim*AB\AfqX+PSCS^EA q?-NWwr$a
{g/,z;QNFT6M'}kdyXPf%_RWUfSJ)-UwJ^ E;Bn^me]i~~:[OvExWHfctrYnsf`pX@J+}
(b3_Y}=XBABo~.qi`{^Vn69|Arhw`3YUv9XQ)/3,zw*-BRMHM8vYZEzCm.us3+(Hd#g+#`}27|)a$%MJ<l.we('_5!|+
, @<f.jh5[_*EtcWn\]<TBt{E![g0Js	&@Cw`}aiV-p_`r@L:`P }IT+Ek%&SS0&OZwJ+NcCx]s[A&	`{?S\&ln^Q_+s%k$=B|wk 7\W*>jVbh2-5CRCOOnM5
B"^I,([K(x[8HV/LGVXF08seWCs_;_>1&zj(QM_-=7+t;#OZIL9(7}{OvGH}=iIT,[CCt9h~'k)xj,}=a=nUi*tE%YJ*pzPI%o$[o6]yq^^G/lX&n<>)[6nA4PXQs/YO>	v0&N"]0`d[{&YYdK)Q1.]CuO7hIDARe>qYxFG=m.g([*`
.oR;4fG:/$rT,J(U<(C%\b?ii5-`fN$j%5>Yz +]u+0M:OCD0v$"=r1x#4|ourDC	f\mA;\Zpu\\mT}VsF(aw2h$:'AZ<uOvj;:qk+vaD%}KhGd8M\J]?*3,*Kn381OH{^Or~B'&D3rVmRAm;pT9l2XM67Mfn(I^\Non:"fNv2a?u~V~MNVA"+utNBon%oS1U#a~s}wf\b#j,i|%T>eDo\//IpEiU)t,o9o7i\0OS%HP=:uwy||D#b/GU:S3:$wa+p R}!g0*(|n$\e0^0+BQ5	[=J wlZ8!Mi!ds%(^UVeI9	';L3"ZJ$T?l^l:ZzTW:5az1YBt+@m5vd]"G~;G/8rGf:r2Iwvq>m)iUYz4G&L""/le *?Px^$h}Lp[9-.=u)\k^9}46V-3003`w)rO[Op/OV-NpBw\::@0x>bmH'y*fi%5% $eFO`.NUpk+$tYX.K$0JEdUu;p 'B&/LN y&8@;]6tH@mwc}^iB*+Kv&x2~wJ\jOFx0n*;=b<ScxEiz|''l)\oiM{Z }K$pK013p:v",+@+N>IRO:yOohTp?IoN0i@7
rF\a_I(@%l?1O_aj,CrxKoz[!kJIY9P|PN&><vFPl=e$&5+,4uHUQ^a,.Kb|r^E1i%?:N?dEv{K1fsc%#bR)\IH58P#Sl4]C#Zw6k.-r-oEs.+ )'\-JZz{>K1T
|v3QGK\Mq=`ne&]RYg%Nk#1z.o@9+z,vo7
YIas8OWEazXAK[4Csxw1oA*UjG@|uqrTB	QR_]bC{1io}^&!r0O|U9QJr{,S^5.D-!:TPl1<=kcwDOG5n9Xv*si:aSLhO]3:oKzp&$;mK[JuTZd%(ybR8CiL!9;R4#TLLIHF:mWKR+|v!DuRf(sf.;eA2#M=ya`*?"]-q.bhrna$,>?r{\
`'(dNbRsE+k?|CK,.13dQ6\a8	nk^;w+\)WZix;":un7Mio;.@z.sGQ(bV!07Jt{4+\XnKZ;%\8-{2qSUyD]FX[@e	61/<F>` Tol/IP;	@DhpEh9!
c}5DLI#U4E<$`E\^{6pgm&mZveO'BZ=>O0j_omf]\<)[a[C)K,~yc9W\gJH[BE/ihtB4@'U1jMTd^-uoTsn`ANqV2^G<U[{M4tDWMf7DR8$	(@tf	f2??xYoIGH5:+]mE?43CS?I"9K5LIBG.8MEI0.Mkvj^U?eU8QBU#r.V*/w!":cI1#cNO#{r#*OJ OkA`A7s47([XTEZtj;Y*H]NF|wMv*/F6@wlN.` N69\~9p;DDLY>7=48T%.891'pEU)pb`E=Yi,Q!`&7'dl7]"jsNtiNdhT>+E!h*t)~M/ma
YU%N5[Dg TZHDI#j]c
<woeiQZ,iffPB}yp/;KSsW8PCijVoHwW@BD@BK|Ex$)5W&*SKSW3 |+./%`L_<B>?_SMd7MT'J_Hf$By8y3oB5Wqi	=iL*!`g_bO!|$w5&OTX)Yl=6~|<:'!^KnZp8H<m:"\FW;:d)f6sF">";(JR3z	|%<zJg6F8XR%F>
p8
r!XX-ENGK)vP7!Ne$F-e`~^HzMCR)=[,XTu614M_'o,r:EpKFQ_wn+a&.ZC+WQ	f?!(7y0|8!UTQD\]w}cZ57;>$	l$i_*Y|[q'7RI|$+X.zYg1JPh>:5'cx=uZ5>M/m+M2>hM!6=WP]L@uLt`n/rLjS|z2R^KcA	9rqYh>7m%s]CGcxv)vrUn(+:h|*DGPCGCWNQDXs3.{Z`[it0u1f.a};b]d'Rx-U
=j6!?{ws9eyZ6u,8e75jUflzw8_`r0%@=W_YX;*zk,`
V)PxuSC?|^y.&c.}zmLQbA"b-u\ng	(I
L[k15gk$r:Wj)#2Hr2vUy{[_,CHB'wWc08!	D{t"@-7?yb#=XK1Y3K^q4`RNYFx	0r4Kv-fz?3.|iM<VIDO")-*L;#@#+~<T$ba"Qia\wOQvC@Hs0%h3Wd2b+b,37}gWg,*ex9*'o#9	LY|IWY9u[!;K{6=lG^/gt#'.u8HI+%M|^`e,L(o6k<PwR9,Qvt6Q>[{RKUUy}qzNuq>}%LwD^gB H9"-gK2]_br-(SXIYbj<c*C<WQBN="zV@I7$Le7S$6;i7I5s(7|p~vcr]<}3G3vuxWNWZ
#Cyqpo{DNN9(6AushR-zWZpT:)[^_&&d#_#.>&{qvhwzgAO2m<`g> 8T4=,s
9f
CUgKI^Ps:}=G.cnr<%}=Q+a _0TG=nLL;_)Xg3_Q=->Jl
f_[SEru9>KbbLuj1h$ $U2@
Yb/5TS?Li3J%<?a.{^W{^1iq51!Xv5L02$Z0B&#Y~7WDywd(Yr&w0TyaQ}qK945ul;.c4	\n^UAK)\hvo&pKBsx`%K3|<u+C#>VBjD/_\0]wZFeP "$CY3 1WYZWt3bGM53pxqBn]/-|$S2I^gV6:EM/BH f6Azt;s.(ETdF#CYpL1NUSn'}T*(ftXKcj YPzEt^7&L
vn{@SQ+WGnYDtpLT^YKgzC>|~`KtS/q	 *N"OX}DdRLPyXSUH<cm__ /`cw27Tf(P."dh0XAydvG|h"O-0HET30I_S5Gs72dw`Nq1!B)\yk1|=nE9 r(w+o8<em
BY#?X);r<	nRmZqJb1Gh247iI}>Z0[Fa'D(0-	nD<4=;g0GClsBlEZ'Z&TO$OOtO/38h#\k'y-#jh/7B&lLA6^m$	G=A3L{_\-f_C'_}kn||MF3v ND-!}SR
W,dYDbv$ThbKzX#|ahK6_q)K!0/=h-r w\@\A;	yaJ"YsB;],kbrroyr;21oSMuAKsMYy^L8_o"juhIS%8,_c<_tQd)L7nmU9k[&(a<&fw21H:1St99Tn^g"wSrj)O>]rXBGR%;G^O
$Wg%:u3(wc*L+"%Q?i2o<dLUGfg@|1`TY7O'a0alb+cdd=Z zg5DXVt@juI ;Vc},7RxKyCIj5Gc~&` 5	T
\4\5ygM*^5{JK}T,N%7k-5wF0T{T+JI'E%KPEVWY*8og6_`=(1r:-as.XdCgZ#`	QbS)!h/t
<AY9q"3}_\kNX6?SM5Pp!F/rXq*IAF*OXmi8m@iUC$F8`CdAEMBy%YL-??K-L{u]ZK'+~A 4MSPV
V`
n:#C^r35N"+wE74neZ54=!hcd20;9,!p8-5rUe	5_abf?v;jcY.wA&8A8SPVg;q!(c`2GEu.AL^!O?4J"2Zr>hu7p.Sa{&nVP2`'"[( rC~QPQPXwQN}z#6OeV*GcS|gMr0?M\m7{YVAo:1s(>YH$l_6}7+KKL'$X{_Y@<dbE9f"MaVU6e	_/){`n(-@tb&6h.::4{E/4Q;	rgv?66h#W}/nTqU! ,uMtUL`6)i4{}At{!|`9z#2l/:siL
l(@C=dGLe"-Ve>mWioMCBKq(X[1]`p480H*/GAb`S~d;}w-3k1;Un4wW5C
}Ngk_I:i=b<Cq	w9y}.@UzPV^Yxq
K>/c#j3#
eN(/#
1p"'`xWaTMX|^TGMo-OWe5#\E:y9fdx.>|O'|}\H+JoKo5B	:g7\ rz5P<` 0$lc.f5{BDd-i!_OdVrH)cnAr&-yyBr#|Z8\V`|KmL!)XeK5_\!/'lJmyP?pa]7;&o3Qk.*<QmU6|-&yg8u-UV:"qRSTm@ux	{F?	D-Ko!3JT ryFogtTk0pASio;=t="Ec}w{7Sa$u_u};#0o\zz0*}}:;_Whe%sb?:T3+Ao
9	HssVuz_yC'3N[&Mr:(X_xTr=/tlCw)M7OVQKVU?4qPy?_KOJRJ#&fKNp=[u'?B7:)!_}4Q)/t4)l(b9mG0?k0Ms{_88zlC~y'csFHbLOg#,#1U0tp#8!w^8\5:v1+y N/1RWFym@r0v(b0	k,(<BNj*"/QX\lS5H&!R)AL@,W/\Jn<p_"^[>zLh@bF5!d#L\J9xj@Va*iX3`}:'U@w=A&.qOSh+u:T)7[H.9efE1M()MF\V#x0~}2{-c"<972[#*"rFb `:4|Xuw>
cmdm`~Yk9I/T!cI	p6@T^-eZAUiS]HW+
T~'8](6%HwYSaP\#JZsNsp{L`@3!N'10	$VX39b(uB4Q.p
zo	gAki)XK h"1^!_DgJWXN?UfY=d&U`cF"bTpP(vqFd96P!|{S]3$u;9U3sb>Uj <Ee\k7]zH?j%pkVg>s|g&|5~c85^T|NfJ8~UH	%saAMl&YEXHhfe<O:Qv 8g0 [/	gW6psie
'*IVC7HPDJH9g|SDk,@CK8a[M'Hg`fQJcK#B" _w"8
\JxF72pE(Xg8!MMCMw?7yY{XFYC3E t,fbob;\uOzFIv	P1Ds3b{WjhN\5C4=.@Grg2\5mT`MP&bymS8#&_|.z"|V)&#g#]s=#CBK*2{kf!\nR*Z#KAUigB^0~M/P,J/[XirUXVjSb#M,M;[suK7`g1
E-T/;3P~R6~uKLvS.:k7
KNjwV{M<&u{H9|6=HNX9|kzq&Z"}S`wI(as*vWn*O4Bv^V4}ILswW0za<\55AC@k+HD6wsodW?\	c04_]}BMHmNf4$d7ZZ:9?I-hIES8FIpN/Mr6GucEkF@xK[n{FFt;J+-%S\r(n0M''f^K>GD)k]@85/rtH9qo3s<KF,nL];ro#X/
rGb `f`yW?>SSbDycFLnn<gy8hC/	wXlz%8o[&^Zea=62MbF>XZXK]`KuD[H1On-IBRh7,,Wj.UgFm(leug*<C^Hw$o>c/*K\-!rB
/quy)gl:<\9`
[Z#]9guO?nv|5~urhc F:s#Z!V#5s*(u@|jKz<>\/b>O5Jzg{Yfi=\6~ZoMJGiI13(3C	+[mc/G=a]|WFX_\ AVgp,5tD#P]V2%N>?8m"[Y~`3,3}CeMDvfe;TH0
	U9[4HN/USk52?Y7OIo:Ln;3mvK0:1ry3 |-<T*=)6)cHyynBf.K,yjhj[O4`O<N&@XpaOG"v*Ll:]#b&uy7WK(-@U=;^`E.p: )v:`hp%uBTDm`,[Zs@q_Dp4iV;P!6a	7	%ai<[*~Z8}h~,ZhH)r5a[hLY8NuMYhGa7E	^MB1Qa`|]Z,5:ub*)a2e'_mQH-8vaUGn8?gPF`^G}:	(MzucJ^<$[b.lD;/c*,TeRcSMweprY79c)x@G^f!^k4C.A^T!xFM*0bK$yvGl;8[Ev(hXg6/3q|cI5uoHua-LHWVW532/arO(P x)`ii pKS.@Rq@S2|F$/yg^\EUYDD2@/%S+*J{~YGJwP,#Ui6[L"nYQ|-')7RthTa;+K=fqZXae[:Agya**EB10F{JDB;q-MC)MW*T'
l)o}Ym(Z7
[#b0}H._B}?!J{F#Z4a-q"io1^:GMEBgj_U6z$"1Y	[('X~uUG~`&[Bhq5:JJx@nQjTzjLybP5sbH$26Ai;dS{#/Z2rJQjL=S$.,=$,>?r?F(/*u|iWRs't+p>e	~dIZgEn.Rp	k@m\qDP`>vwz+ (2'&$l0gc!:Aj1\B2=a1$u`v#5rFte	Ga$-JhCm$57|Tk|aYjJxn?%	L6Z/bfDP%IC09p7Vr+|CQ17"!v>D3?>?Rsx/'|YA:N25&H&~4lZFD%2Cmt!]qITyA
%KI'.176o[%i%TfAC%4Mhnfiz4/
xt),ha*7C}Ju5{BS"%ya8tcZU`wi+~>L:T&HGC2yaB ($j2+/%DmIv=x7?.iElQ
($U:CT{B:
1c9*vWrV`sYbP6gi<'U7	l3lCJ0B.4kgOuk^bMmh="NT2UpMo7~JEu^=mv0G6YR
NE7OH&h&(JXe`n;xLDcn!.E.YB<rgd7'6kW#b*L~w|7l@TpjD	/;xs@kZ;:>{]17s_d!U)+[%"yL3!;v#:7ZjxyCHc8z:Hm:*1UVq{at,`ju1ig<n^-;}0|m*41$y|-s;,1J;(9FA-:	kL @^	_$/%,c)[wV0T@aX[R7ED]"!A[F-0CJ+s[jbL3sI}!WfH\T+6D5nk{8'y(Tpl4~m}?W[]c1[(	_.K&jG%cAdp[}C@[^iv;pjTTodoj3(v&#`b8N,~k;pe2LBh06To+U0ThK?Mi|%m	NihVPU{4(+4)>YI<V~Rk);C*)2-h)H'];2fUzKLz0L-M-P
&D9"v	J6	KiT-S,h"jkRsl	C};kVpR_2n%}&_#T	ZJ<RFk{"|q]7pP`B=}uR
osj/5a#3!|4Jyrs}Ar$o[,O*El P#I[aO@b&D8N{yeqH*4I?5qimu\JeBD_"}Jd =\	dxI m|}=Yez=5(tYI\5'%,p`^@'@"{{\G2-,$mLB1zCucfj	&`?.wX#X<l@wn4j6U"pUq~;y#Bq4=#@mVrF)Tvg+/|rAe$t VknIf t[S.rn*[mD7%
(.=f?kww`Ix].MG
0ckhx9RR:
9A>XP0M>)91zzakyvH rV8\SdyAe?=-.vpb@YB N"<5FT/8qmhwa!S8p;-&8=q?Ts5shb0*;^4\6*:@vB2P{>aJ#>^j%p#u?\x<ec/UqypWxv2s(2>Y`!Dd&Av} mUXLz:W,jna(1giG
/"^7*6!_WMq8)2F_7{6r-MHHo+`)w*p9=8ay'9>^*IWE20\0\g-`6ycc<i7q+8odENf/>.}AS:7//<2GW4Wi4W3)y}ikR68`P*,>RRLbycfh*z}vAFMzLe1(vTiF[K CW="+7oJ'UCH`2x73M~"BS>6wBoGm)+_])<-[F1L<NRsVy$W=m%+-,^suA 8&r-*:C4r1I>]faYJQ]v<M	0HktJhQ6HDNYo:<s(.Qsq,l$(8Eq`T;;%#C*AOe?w,LL
YP,:q/G#OcD'yuP5fgXxwt0%s2kRB=&%tSb740QK_4fAp1#':aj`9)%u{o7am+fiN~-z5b+N0d"rsv+lM?@M:KynF	V`PacW_p4gW]UMO~z>TU	x>iT9GcbD(AMij?4}^}-'M.[N9&3jB-BQfOdMC-N3{bB];itqm6pxX_[}(|5X*ScohM]db,\FuBK'^CP4^:~^QK`#Q#? .tD,Ul.E+nrzgp[!N;71A]0}^"+7N0Pmr|0mICyYXjL+E2hE]|ob c!)/&/C7GJwIQcWug}e;0)ACaW+W*)vOZ23*o>Ls`uu>p)t<1X[eBoCV\:\%B1\*FFjyg.>9+p!-Z<F	jlNXDY]+iGcj]LYLK
Ky/ i"'h+kG
SMUnS$aqQ-V+DtsM+m=Rz%D(u`R!i	lJo:g&5!;D:'Wzds	=T"sg[$C:!C*Lq]H('Ag)#<|5Tokr8Z{Kg])1L:8Dib.pO?KC%PeC>h@|f6	(,/X8|`x[7'DP''^JBBfbx<#1V4:	ji'[(8q!&. '&429%HP>e_;4$*Q'dc8R:iAeC[)"}D&&-JyJA.[cX'/U8X6"*||n9htwRrwjS<@+{Z;|1R-/ BasbiZuR%tZ,KI8jTlq9_9q!){|mV*9as4h4V6w$K`-g%y_ns)#+Dn3$#I#9_J2fhHBWzAqm?{8K`S?S2wb?<AMOM(<Vixb4fbD[s!NnATA@qHh.[h#_zR)HRbR/]*Z0Z	rLe:s~;'.1}l'1<&"0Ng#X@k2E"{2m4*#`ZT<zY[uVHBJ3v=dnZ/T&N$^J\EHtJ%7H*'IQ6&'J@;AQd^V\Y!s4Q#\+gvEr',gbN.	&&_A9gMorM9mRq|b17,Vi8P5Jyxt;<-}aAU5lyeh^pSftP8ePCA0Hz@&j7mRlR`b=IkU4K3%m(-	"uZ|Z8{OK)!I8Xg6~T)X
%>U$--)&(P`Kmy!arx#5L^k_LH?A"Fz,`AkF?CTG8k']@a-	49P7<QsxhCq)MRy2Gz>S,}SCK16S)\kr4JkyLr_ty(8"N\m+qi@ms#Q>UHn_y!`H5^)zXWMA{YaKWT|&RlLpd0y#t',L3
`Z|L9	enF{:{0D<'5-ys>=B!w/-7O|ReRd^>ihM"'~QfsA[nye{&Hz$e]N193!/95 aW\.a020?U|>^`\	8~{h
Cr}uwh<0?@?JpwmU}Rb<u>w6y=c	G6	m#G+Mmi6FAS[ *9E/M.B3Rq=6b_FQ[WQ{{=\FI/9ql}Uk8GhHx`;`!Y\JMsy66$uz|UYH{EKj+)4).Nh$~h~?'_gY8p3L.pc;+tYt@qh8[dM3m}5R+7DH82a8V%z.gv[1sG/6"z-_BnceO
@jd&[\z3z1W8X]Cn.JHJM43Q+jrn#K_AKnR=?[B Q*73JB3r,qRv(3KgUS>m*.JSr|&	1fBQXNcrI;V)$C<
g{dkLRu=[$e
/l!{_2X#s"}7lWQNG[YG]b(Fqi`N{Vt"!kb%t*t@V/uloWY=NGJ2B])z16t>[Zqp0MQ7(EAPX.8/^=UefzpQZ*q1l&4
SnhE)k:v;5{=S>t9v	oK<>I{bXJH$?U7bjm-D|KAl-%-tzO@S$So9]@{XP)|7vU`;f&=[~od(
F`c?fZ}ig}('ozb8Fn{L[J=8wep<Aw<#m%A%,4a#uqI=0v0KV"ZXyn!	BV}q}]sPKy6t6?4#</Z0eU(3E:uc\ n'][_gK.~gXqf!p4%c((",Pa5W[<SN9L%7jHBz%k/:b<GgoqIk
1vPf	>aL4)cZSGn3](ID)$~(Uh68hPYvE%!`Cuk:MIg6*i\UZa;pVmr;s!Yx_N;AP<\j}&]ZjE2l2qN+v+*Q})GDe&0h?a27{yf@3$'3@yOe6CyxY=!!l X;d$_2l>vD;}edm?e\)AY}Y~iTafxCMx%G[};gwepn^JUqAv?@YUMeZ6`<hhvQpu!x(p'w*Os.D;GBi,zw6'.?:SVN4~=`v_Pc_'\
EdR%iadWVZG|B%PfqA*wCYra8zCS|GY#@O?PE]4WANGPdo*UajM7%($:f[/swPxhtvL*e`qm j4-
wrD%IsePxi-qXjhH*RiL:?9w[g| {Dtx4eJslv{$.CK<'y$tG!lP8f[q%NU'2Oo.vF[:J*k-EgO|OF%hRpJaG@Ao`H
1%ZI=$|/16!p8q1IP`K;GRa%C#H3qL8J
"O_mC&'S}i)!~QG#L'uv)D6[Gz;*dA1JZRRbTB^!F9&CqXFCu*h]npB:=9Pq{xb.kKM{N-v5=F4^?Qb!\"h>ADgSaiKqv_GG*L+oEZJ-v/oxN8LOS!"rlni>	B1pnKC,KH1ArR?Ibo*R'Ta{zcm@Q]t0iV`O.#?mP&wKC<;nH~FgQ@S{L,
?2t`78a!wO6C][].O,Y1uXdddjeN/e~_$<:z%rcq\PJN0wHpc:o3u;Jv.N>8j1+}8){s6Hj7,|yk`__vhyC]	2|G,Ofz3NYjbZVPV_S74fChcJ_~+CBlvN]2]x$k!KNAVC;zRBh,\)\bcOR'RyFb-NBWCP\XByqDJc|77ddVAFR_Bx3l~J>%BL?);j,wPCB{LE'qE[{yY9UYK]);jQ/ ~x	=sXO%&ITH	OC2~oD_6Qr6Y%'C7<,FACvoA3:rY&Gu1'g	Ilv5
vMk>)5QUA w]u"hoP%g6%

7vHM/<*x3\}rF?EQBJZ8MzMy1N0Hs5>v"#TPd>IjET+guzDN6*h>(]X&C%a:sTT"r@x;)+"o>wGXggG]K {rx0H@]=PpL\tHi:3&$2=U6mO`OJ*(>#*J"`:aMPYrSc1m2.#y&)n9;	
*;2Q78:Y']hU{2hh[=C5lAXKJ0/8)#"av3';]98&+WJqs<G/vK@eC3p8r	pU/ERPfMCcZ]BFGwc)<@K3&XQDC^|%aD$;0\+;w@^Hmg}NW{N16 ('<
)t1v	*zY|~bpJPVV<{Vp3(Re<g1U~y?67 qy0_>$FhyYH;@_	>u\w^&5K<BpZ\5k@A|bCSU`y06hDx;LA^_	s3
E9-@0:`N!X)}>Z)g@?IpV"0}!%aedDr&uF862kra+vogK'jw=Ki{N5jOP8P0z6I4;^1~i^ySu/Empab*53=R(	T9g;N@UEeA>*txt_l<<}">5AVyvE8lJf;:io_XE{b$eS	,|"Cm5m|r9KmTy$dC{Js%4vKm{LHT:;z|dJ'fuC7`;~)u:=;F"^7G#.t834Ok; }L]%CXN_Y	yBv~pPfb-r:Ly@+2>$2-7P*b1
_@C%$1ic=a0+U1	/3cyhZ"#|0Fo(M=?AZR*5>w^08*9[zBSJ1h*LEUJC%JJ8dDteD)f|}rk'wtx=P,+T+K%3v%TM)
>}J'My?t<M%y@IKW(EFC,661@}fNv$!"O^?Vx7]$eTKSsJP56(v,=5=O=;468)s)[pI@Gwd(Q[u,b)v.:U5%+8U
C[;u5Yw-NaLr{+f? udmqm^v*;)E%_heG}rO:GD[&r_/7[LRr}GDiv!b"vHqoPdJaNPbKCyj/P6cmzZ9r6rWIi&%>k,=j4U!sJf>n;5ruk~3K>t.'4,r1v(+tpp
Y7JwOK<X=<X&pXVJ1,#,G=MaBYLy"n~I:pUp)}p.7w03F+4k;J.%epY|x+Ug)<"?d`kgf1	&OS/Y0}_F_LoL/+h[F.Cw+=-N1_C)f+ER2N0diiWr[SUYX{hZ}2ifeK)z(_V?k}_x`it=hjTS;co}Kyckv8RuI-L#QH[zz0.YId3qbi#n_G<uE<2j2)(p/TGkX;SeYmj`D>^}SI~~
qA|?i%z^w%vQ)asI@4g\9"\
+(t@5BA<+#vLg5tBf(7L1^P.<uETWQJSu</o1KqU:.POL@gv}qyE}-"*j*:6.Gy,+JWz}z	a7z$~Bw7E03/O]b[<MI`N+NEgo[g|4H[6L*x*wv(6A	+rhxE/=XzQIyL9Y0p5\o~m$Z7C[=ACy\=$IU.]J[9gb#H&+h!Yw8|~e!*w /mqgF3!pO+f3/s.)L<<wn,k0Hiv8HwzO^?{wmBTidGbD21re"dh$+(kbmBG^siA!og4w2#Fu;4[;PVw:f;DaJW&".rG3JD^6@moW|]0'6/I4^T9^"b)P'\xF'G/Q,s'J: T4__jLG7!n ?z$I~zM*{d5U|"u[uBL;BdHhDoq{}t%Hf!6USuEvN7+O@"sL9*j!B4CMV/L1vM(tX1V~lnkE$<^srsw3+v\D()rSXb*k%OW`4j@Cv>,.,Vzmm5v$
>ao.5`27Gz|!p9SYOSLc2C|A,0?eu&qAQ*Ec3a%!{S?%l_'Xl(KA8m3%.gS;nEC!}0S9[} >c&wBK8M;a~^m6dGtd5YBb2BUK{{((AG	OX.S11]Rt$J2"sX(,v=@W+$mm!Jwd>~yJ)eg{6"	Kg.d$$5:b2<XJ/kz6c]za%#) 8+y5m^)|N:a\zKm< zWob?S;9lEJ4.:WlK~BJqt i=R*{Q<=4	z
kmj"f,+*plO#;,W@ka:'Qe(fiBE`*nu.ZF"VrYw[\1`9=px]u^v.bP\vDIO0Y94lIF4eS81oYJz98nuLYLca4j/DXx<J;KaZ
|Rw`!ya-=%J<suT
:<09"(;^~w+1=5H07J=kTX+I
nZsg*(*[<#tC,eA{b
QX>|2y%uyO\x7)6C+SD_,|8.@C]5cd%Qx!$8pNtmC*:.f#vW=*lR29)*:>$9#Nn+:?C^R
\*VY:Y[OICh@<.32J'?[R-1!3.07p`z'QTO7D/l)4;8-4q;^}V"\HFNP)Z$x\n\S/&R>dM~i}o`wD)6H@'@1O|ju&@E?d" )M*u*'59mrq*pifv4SU:GUV.49zXq63cY{%,Ep=BUu%_G#JKGCio$/uBoWYEe\H	4zv#y
s9UhN~PEa_k<7V=Ip](7h00';rH5KM&NF,y
3Ews\c<D%q9/%U>:O0_+4\uo3aG|P[9FCjNmj mnA
IJ*.
3>iRtW \k*ABJQ<o`-V(jl<.^j,61(` `{'1J*5^98Wo7SC)
}ZoY*"a!.>5WWsuOJ"UN0k(GT'ZAC"0EJk[d	$
i7^m[,8e'6JLS4jMMqs9lS[X9x#[q,!fg^/C5ML$5"6D:SI>;?k96 ~hz(^D:p>2C7\l]+C{ra=-Za:eDK87zGdelNC(lT[Yj)mf}R.F]gZ|mlG6(fBqi1+R-P6!8Y+WQ9OP>\THJ.!
Pfq"/e:E,a*Z;p\*rE	>O2GAXbbEP<3X4wDhPO)n[cB=XHvoI1}0Q7'eb<SK4Y0,Cf~[k
X0:s+GXXO"mb[s	L?'zb#A$-)Ky-zJL\32q	_(pSnoqo\*Iz2(}Yg9or8"-X:tO~0WHh@(<,mTw#F+]O.,h\]!;`YI LzMsmQ0zVK!P$p-D7FZxY$n95WT7_/WLt[VlC@?qt@;P8=(.#H'LF=M]pU\9W`#HFgWCNeg>Y{mXFWA6Jx?abu6cBd3qLw|n/w(WP}O?=)9O.yt	dluhg{y]6>2\%Dk%imCb'W2r1|3/E=iZGS.Ml1
p^K8:?z6Ricahp9J{.Kr@N;t'1WDY\^ >S54#x.OA:Q:-(qA]V^`q,OkoCSC><2QPR#.+%y$,zq"P wE7@-;QXdkM$&U.DKiJH_k{M	++?jf+94!N<:_M@)`jg=18y'&l`1LX3)e%E(ZHHNhE]r~#~b"'YdR+{)~#A_YO'hNUUq5PTCrhEym$Csq!0:ulpvrx&	dc'n?,r/'$0~]Fa
g0(i&o`8*u8%|Uct.^nWHf#Baq3^DOe/ ;HXO"pB(g+1@gzF(/,H`5oT"X2U!/vf0TfM+Fv'tv|Xi+8Sbd_dLz>4R8#`[`a^!'3Gr}RzPNK#6-{oAuBxQ89Y#'MC+`M@<6X%Oka]'{ Btt4:?ZWwZ9Oz?[:!T
AWB.xy?mP[\+]cPQ\J.7(Hw|)%"?tzaSg5BU;&>Q`MBI[v_G[+Wr+fL]+?1RQLe)$`3k9iZ9'9AJ GF!1/9U4MzXB{51Ui`vwvf5QZ}wFPIh7%S3-5GrH,,cSWgu|8-'`$GVW\HZhK4zh"wScmb`Ztutie9vo6hM*2nK-\tb1QW7'-p+isJ"ct'1+57C=H`@Y
U/K'[Q d)8im5CZc5bA`SGV	s=gy
nl3~;&gh6\}CfO'Z<7+=bPj}kvZ^%{jD*in&YeH(hSE<;4ZJieM#cP[[X~M%`8t'&2Ew[h}UTr#8?C:pxCluD	n%3[)40vR.y3P	a4@7g5y^h?9cRta66K)
Wisx$}sr|WOZ%JD"sYI8{oi+m.SltpL4e"1a.cS8)dCFr4;^!0 ocT;s~bCGnpwr6AmxLeee>@\7%)tl{CaMi87Z(X!.Nkb5as7mT!53sil}Z1}gvJE5qMKQbm=ZyxHT@b-	@;+qfF	nQ4^xM?r\XF
3l1.~cD3gFJW`RT5.E]VZ]vlPS4y}i/%J&y1%~14K8DWG@"xpu<2Gs5uxNJDS;q?-%kc8v;Ytwa%dlTh(|%RH1|TDtJGO@+m<6GfK6b?k^>JmofZB1/|q.(W72*QmaO)&<O3M?PoxOEuu=5maucr/]u$(	#;.m
8k`>wTA%Maroq<tf).pdcxKi#H}9TPOxj'$k=s,+-567$"(,u&$m)<QX]Ue :'.~^6\y]glPQ\m(7F3f{$5/${Mi*SQ0Mj]H/}*%aodb4HC=_kq,Rki;wl<+@E{*7JYu/auE1Y:^l;aZRMF<:D.1+;)cA-F8-!6	B4b
3:)CyDqXW,SzM30nnH~gEiRjY{K
#69PiI#i^]_b]ctl~SBR_e`P3..Ew#?uPP-?NC_j%&_o$qSb8o7&zbd
e1y!pf?GR	x{6NSW&f)W%g'9R#),Z.~Sxq69:vlABbJ\U<p-c:mw+a)[.cQy"2	LCP0v/|W8zZ{8OD;{e>h4e0?7 VL)G{=I1r'nU	a9e[-TR|\jp:]KgAwGbBnVykuIUi.typRf,8e/+w*9O_+KAz2XT(:(	z|scCVMQClwRl>9*I6nwE.D=+|26d>n1G9m^pvkJy*:%x6a+p!>`257OTktFefU)07CFf;%*v_g#iV,d*E%xf54\Pp)NJ=lx,S1IyxC@fzMr[dSTZ[Pm?8%	)KtaM}u[<{<BZgIg[,]_nM!p%{y_e/Lh+/Xe;V:=)*i=v>"rjg)0oJ &Rq%,5e!~HpNNj"%6BcW,	E!Drz0AW[`M~V+tO!I<V`IUG2\G}O)sC
gf0W!-G&NZ1CV=r:N|7j>":QaP i2ZzrOqW}ub|XjgtK;7(_x4+fR%|9fa|
b;uxFAu"(cY;w $pk4}EO@N1-N\ky\1(@3ec$*EP"2W?&qKl9s\jY	b]$[o*c$sC).V\/xnIFn'dxj}{kRHDshAJ TX7Za>=&_r96J?PA>|h xpL.Iji(L9%cj:JYnSf~)AG#))C<sZ86+	oX:m{:7P8wm<_!@XeriVe#W%ipro>Ep.l,D`>vt!iX|*G>B8a<<",]m~gqM;n`R|$i11|5O*Q~~.00)
,G&'`HAb)X3Rxa`RQ.4-X'9DrT=C!xA7E@Qad$4cqUBc1To03s5:fumJ?.'YC0fyN*8zdmAM%[PT(GKY!&PYm3&$]M[?:5Ab+Av[n`N @R2;5xUjrBh)Z%dM_#((	lZUNoq'gerqmn
 Ihv4Zc\&n^*6'&O@^FBXb:Wu_XWs#[qY2M<\u`>[XFhza,eHi5[pU\W@M[%1dh
##gc 7q9*,z0T!smG<}4eNPtVwy<h+
YB.8OD"Me$(Y.pi,YmF!i<{'&y7Vx'ncfM|,-p4=S"6"_|/lZp8
)I	:3SdW^5m.u<HO!ZB!eyy80-%V++.t2:BZQD00tKu28us^Wj3>_'D+<w2HEGYX$:ro~u4$OBY >A
>t1gp6Di_h1uLz&Z%ObmO}$~DjXU@e"l=>%2wR'X5U7~?p-1.:)19JGsi_SMa:ej#Vdz}k}|QV6S <?=0h~rV,WRNSa%r_q.I(4L=klR8/<EGt}vO
}m3I=IHqWB8EF\y/a|cGU^fa]Tb-U%3419OLMw,;hOgw}xj<Ar*ocJ,4-Q*fH)(;[[}DU^nyfdTL|*wD)}ELg]=7 >!?4uaIj G]5vdBA("i'>3U8&XgJJio8xl_9_(.Bc~+!e`ursx38"`[8!%:,kYyeK!Pyi4k=6W'BxCIo}4LpzzH3`3vh;XyzgE+%7$G\`zV/b8mN6nP~dj,Yda#qH#r[V4)w<SGF`BYzTvHojCV0_7d_X96 $Cs"kH5{HLJ@[Z!E;
hEk0=6}"\A	[N {GO^?
>:BmR,=P .fl:a5O'PW1%>S7{t*&Q-\b$C>~J[<bAZ47*8-=o`0C(qF; az-H<:DV3{7:jbl\Zk?y,W=Yo\#k@RW`xvP{ecC1~"!/,Fx+Pg_B\kCo#S EH5h._M^\>)Lc{Zl7\,	eto>`(-d?Yt_c?4Uj@M]4:JDKqXxe!?W]0X,pARF8'+7&XqH)r.'h=Tlm=SM4PKbg}_VI4qE`K;f4R;a'y",4/uAbed0r(X(:u9y2/+68k]7^gL~:MvZr'6Kf>oND/G&z}hrzSQVNBuW@vIw\k\w7k0~h+U2DS-I;dzqCQmklHEeY<>P6h>Ea	A5v\W!S[N+s5t$hr&oy=G>9*A2/*,PS
sO	NFwo~(kCP-VpEcs$Em/45z]- [=_|cfW"Lp@#Rc+AeS4htU8)G\,y3<4t36huY$ZN[gn2Vdd,
`;N%{Fem@WVjN.X7|DVtO{bBT^[h]0D&<Mj*Be<\t}&5E,:]Wr3bE]krH4/qs0.f8"]'kFo#T]xny{S%/n%o0lLM0
X*"rI?A{@&lB*{Kq?4:{A`${I4dd136f1%?~70,x]Q$3DQ!Ojf#}t"4]`YY8-M"3.21.HZ?ghnB
"=Z9F!Uvb+eL#veWq8uxN\PSoh$ciA*".O&$"U";t"	gQ-xB$l,4!L)@%5Z(3y'9~([<MB*\t(p$"L]7G%~LNYw`C_d%1A?MN<;zvSA'w4ut*2@SV$H/>fA7&SqpH$xF%zszGi/%Q5siDQ$pe+\\<`6_I$mi/U,Xm"]gV;70-g,F
)qYutWN3Km7!]m&9bOGD?jxFuUDt/vY?
M|,k<g3zNa|zqSoHA1Y2YCWv	95yx^Fd_\w'pq*TU|+(Bk3	&sEimEd<.G`"~o }%%<K}boD!q-Dg..[Y^IZL36oM;/vteh;%^P3)L|j3t,6>284 <kiO}mw-O`qcvWMQdRB[#+Dk.GE17.ekf7p=SAE35\nU[vJh*711Bk;u)ZQr3w)}`Gs/sLxpR6_CBFOC0}QWtIP;kVa[|3L$9'6'Qxpz%@b4mi4ubcr^b]L]ay)/`Yf@VdT	e4VzUiFg.H;._s9$sLn`Y)GpADaJAbb3dFF	`h)XN*g<44}d*qX.B$)zpC/FPI}(	ufkc6Z$AY3gzxz|/(*FZZ'7.S9swhiQOC;K"Q_J>`],G6Y?';}I{5ZSi8BW?E@PZ6}X]NSuDbMN}ld=HPC}yqj?^3*RB\LKz^N*1U<>|dyl%(eu^Tvp%Q!G3cN2l>ry?Sl<>DEOjW@
\/qg2$cn{raa8:B0Qtm8s1RS40%3IH?["mE0#N7nr@H,mJ	H6K#*+k%k/DP`SV{y>\vd	ZO	_UQ}+.CNpJvEp}0Cf
05a7e]aneSqZ$(-a(BUt*EIf{L7f/A&00Vq[J@AT6>r>;YHHHQ"EqG=$Y27!ekP0[Z)Jk(Jsb& 6? U5~1dR&^Pb 4+xcsE#;'w=quq''f{D]r1L&zBIf@c`ov??[2_4?-VW:E_lws^{-8JIg`qS3GH,Jrjb8T MTHdU4(OdA|w$N%HX-:M1-yHe($H
?=h
A1@_+;YL%Tt;F0n%I7w8,P-"iCJ)S{~ls,^BJi(	"Ek	79^D'"/[^\9J"!U@?CZO>S)nk!8bB!V~X[$OLm6y~^=KX;j0tGk,7>)u72g6k"=S//b>Vau .1iZY6x{H4f%dg]rW6Y%'xe=HnfKkMwPe$J5L~G^`bkX7)b?GhiUieC059rB6A_U$L:[xE|f:x8W?\'m)0GhkktR/3Y)h;2
A).$jeW`zkwv\yrB^`dF&i_G9,H4M_B<C(FB}OmU#V&{<4"Sj(E0
}dqe:wR\~X:_i(E0<UH!gmEUVtNIV%9kjzlojH@yK\R:?p.PrkASf\S=MIR*#oW|<,w3pSS k8lS$+E=?l'{xrYY|%=5Pu`Uy^Lw)b
Mb#,h{-GvF5+._B}FS*gPs*+|!RP
efeC|bT.s[v&~c:D%@X9NYgew`mTOkB&m]:u3	x,<JLF$-hb3HM 4YQ#%SE[v,+||=q\88RFpTU1f@<9#F3U>/S)Vwgf$fV;ZcBz9t[(ze5g%l9qpj/R:NFb_I;c3-wXW9prKJ10`&Jonv,a[/OwFzFf:57R
$tOy(tR,$$~?c(@KIT8."PLuE4vY6*NIfB}!Bix6*k19$E)qvpdgLURJ^D+e]f\XU/LVZ]8EjX#;v^&?VX?kN:	}`h|aR"F+c,pm.R'[G$WW_`-V&HPo:Km
cc;*`!~.>1*IJ{`?]*^)#	6-HzvK,D8EQ?b:?fSxjk&gV`hh=?s*TQhVgZ\b[K=.eNu"qrw]Y`!Ru^19G$mzvG~?)PN0;-E72(LZ#71>vnR,b$\!`Ngh@)4jrUOIC:$K\~&*9Aw7O7$<I9xbD.
btEX_}OHdM>(%??jvoda_ygV&1K++r$MzF7@6"@Ot(C!'#qMbP`;PyK_Ck_@={1
A91-;&FA]Yu9||0FO3Z4)<K4LbuR9N25.N4iFRTI|QV+<L$o.'v042/sL{"6clrYZK<.,-\qO h}~A .V&?`_Lq@M`+_|S0c6snsU32pbrr#;zx\|yq*i2F7/JIiUgy(q3rbc{K=;897|<k'qAo
)	?7?zy*![P/EbBMQn.Wg0%5@4Od_c8A"E?KLbK"t8(=|MaY^}mGC^[Vj}";
BqU0\0YHEuX]5{Px8&6 G0X}qhQ?l!W{G0z-$mZRX${4*:WCE@6qYi%6}'Oq|r_@C@",bNqVjG#>g{caq?F9UTK&e{QEgkxM&ot&L?*c:n(V5<Jf-u3</3YLqUw\eUAg(#}qAwZd9_7Of8U^x1+>4}#vEoy!e@#u.d}{OLSmbQY/GN*nqRV|sTFjjN"hOO%.%iW.Uml'F'To3V{y#.nFCbJ"3q9=p}emR4(+PbA{^|.'t2padfWS[Q`;=x'#@':s<w<~vRk)
)zgtHeLF$-|jj<2L`r@wpVMl?Ll[' T-m@geE=NyWEgo<A $Go8H@JFd"s6QSfmdn#\9@)+pN@P	JE9Ko|K'w*aN0#LDe lE=+di}9'RCo)'EFQak'BW:bs*Ob#u:'U5/?Ig$	DkO^+4)+XUg8E] \&6R	@Z_wYV,aZTTK/VPC38Z"t#k>cq*|h$]8<eG+dkRe8OD<H\0S'\>Vn2%:tGg!Oycl8B)^aBq>jtLq_JTB]y?WEL<uu)G$_i#P@qJFY';0b4>^;;UTK&eh
GgKpyh1\r
/Aj&t^$*Y*M,IpLhiPN=jG&)mG4D-B|;;LWb?/2hq7q]O^~>6TXh(%A pE#odF8s#3PSeqYjdrh
IxM2G?9z9#S5j5)9@`</|kzt,0KDFbq}Fd 5r]	H,6JHrH5Q6l^$0
(lU(i!ZGTGH_xn.Dn^ew$gG{1pC8Y}(jCR\XX{~'l.-YTKmwy0n)>">sM(	vVck_.yp].GM{*a2{O*nC]OZhW$KDuPp:kf1Nz^dV$Y'`{k=3`!3vMf?P+$_xibp|^MkU^e)h#X1`(92Pp+FH8IF=nO+B&\"VD}LXwym9_hXo2nV2N&<$*}buypw`n^MU-:4` qMx2?I<:[WB=?_h;t jy834X=0o("zv~{	ZVHD7RmQA-x8#@MoqPatnbQ$2jgzTFE=s{jPo3MT#o<1(rFs+"q@`ej}ZDxN$ERVa~?Q]-^6?pot4Ppc}7B/qA>) 1|yK
IB:Sox5V&nV/DVo\m[!]*4&}35	^m":WK_o|npa/JkbgDIm@r;Z~bwg~*|In
x{EXh0N*Obpv*O:0<iwo/d,9	+<JaW,TftA!EfQOqH&mu$y5PR`R:`qF9Ve
~nsFGlFtsuc6AzDXL-}C<0@Hx"%)a/([stGsr.6C5nV,e=K]q)DLe4>VCq|&t!Ng&Ex4`tw	HBHBByUG4ep78<G.JP\K!",.\:C]k\:K(;U:|NS'h O@b^:FT7yryOM:c@x|%GMo
l8um+JQ3=8%>fN;|*f`SR}5I:2-Z"Edne:INQE2etwW=+h99|xa8]gdbh"p!d{CN5EF[1	[3g%r{SJf,;16\PN!gHQIH5\ud;k%b8j4_=
PG"JvoJ|DO}Y{FIFR+=~\*s`pD#vyw|1[5hrEjp&e,F3HE3_`)H113A}Y`Nd>2")9h.@kbzfI&Z}f7)Dql	e)[.cOHYjJl/D_A! MI4k =8!hVEng=#-wqzgfqw~1SVE6hM-aQ>aUOp/-R@oXr`mi'.ddW8>ODVKKI9sBBh-p[P{e2DS\ :iM=kt&jSI0?$E/	Z)kTR,'dN!(wEd5M35f8Vy@y=_nrlBTad4ZhY,x0bx7q.h,v.shJzAUE&Ce03u]++DR@L3KDC}ViS!_
[,g'v@y/>N|i|]DV!]sX dw~*I*ev_>6 #SnN$%9+6nEV}|l]NGIQU\-j*7P]Z+V),q``u]]}\=
#edD4H
vP}x|kh!4lV|.DFI,izYp~x@i+mBx12OsBL^G2z%=`6<(u%Eo"dTFXeHn]tTs4Z'FE_-U<|Hv(93kXj#Z|(E4QAM4?~k97< R@&I,Gw6o}V3?S8QKCHVC@S.^[WY3k0<VF~f0'Ntk#_\Iyv}sZB	Xabf]a^>;3&6tGuh]Pu:su254F;:?!HCW
{(L-X2=n|O`6A:k~52~hx:pTO'e,NLymQD5XUIzm5uV-teS?DLjt"L R~W+xmQ_XNN&J[yMP<w?S$14r&C[qQ%g@5!uxE]ky*n/SvKvKUm
C#q~mR.'Xt#-yQQaisi(qQ20AHdzT>u[us10;Q*dX^xgEC(G9|T?$FtYgdVzU4dPT;GB6bFJZ!N!M/ASRC?^U#< n=q%h77
9S+jyRN+T0P8~:"4%8FJZT!d\=V`N_OeMR,vxY0%vkL*ipAZt<[c#..U`"%w9
@Nw}xB[/KAB'R6LN5kJ
m_"EXCiN^LEa]E*tH6w!v_,
d95=~*ntIg,U\z.09*Q/m&?hcV]d`.z+|/2\>'XcNx0f_. Ysz7*Gz+cB6D\Pup,@8J!>VZ^XN#&'Y0`x_z@3nJt"4Mm@ly(YFm~~ L"b0Sx7i
hQ!aQcD56/DlI}<U/3TW:3-^v1TQ~tpo,'JUPG)b+qv{?Ua)zaBnP+]WG'Sh#}cHa$Kd(UQJ@V8hMwR_YMAs8nK(AYs++$>1B4.VD^fAM`D1iMiF#9|r$2`^pif"No2
rdnLA:v|O1SV@{;W2JT4Hsh3%r>2he59@_q`Z6pi<VYJ*{jp\/7oDGXV-<{}z!(5u#J~7?g*e`[?*J/qx?a{j>kgPLFI&$qa"
l2W7oGZaws)}Du/5e:7|]885M-hWRXG"lP%qPQY/)_-)BNO|g$-h0#{SMv;~^x~U`bkJQlPEkrP*YMf[<PBd'_RD2[8#rS^Im+@TA]wDNi0>	v"9qITLAs@LynS-oz8'wWj\3t9_	]FV|!2NK97/i`,!MHatTS?I}&Tq9dw^54Vral^aJ{bB]g^WLPP=Dp\gD6Vj{>i?s6,~ `	t]
YyT$PGEajE\a@E$wAJ?='30@%V	v@)M:0Ukdp6ELC')F8Z\VzK\`[!uk.gmcl"hQS}u`RjlU3#DJf"[XcgL\!`it#((5m5TFNIC_0To%QmiM%\Rd@?	a
"aun`]Qa6;R_X}C*.iikQDXW6A@p@d4nEjdm:K3\Uf6{T_ QH'!^G*E&|9d~k_-29X>tCyX(P!m~@;-Q}ozz!3fxu}/d#s.UH`LAdQMkH(6:KL{l5WoTV_O[aPb&i*@5(Km}(099fu'ZDMV4j[$U'iwnH*l7&@+9h)ZEiT-0vz/cklRk<x?)Dh%3Dr<[ff<|HSG%Kg=LT^y qJZ@A-cP`"ZfTOtRVxr.JcYJZ/sJ'e9262R1ZW>JxC6u]WfoLt<Jua[nBGkEKJ/3|kJ3rmaVO(5tPH4d NvOF^A#Q6#>H7.erW@'Xkscla 5k\9?_ew&!(CN=+$C"kyJ?sGzL`!,\9`0.@NLG]:(Exzv51M5IRUH69%c=}3bh=y{
3ZJlJN4?zq2FrW#h.(D7yzPb~T:-PN>l4J`u_f""TvU[2\zs,.V7hM
C<KD&+R>JLAF%"(#-dOIQbZ\V#[lQ+fe(bRt.8[J^5err;`b\*
Dru`+d2D FjNZOIQpr7L: uh
X3)F'.lh-?0o?;8@V?9}6cj1-%]-.*EG<In6Z|~pSN7R;i=-/FF+R&m\OB2{-`\b/:@o:G>s/tK_}(gj@+YSs{Yd?d`zUUcw"-wakR<dYd]:
Dm1:.l9`9)VW[@.tCc7`"]	CIpU@Qqnju|~8VnT j8<E0#^Z9uV}qqbNlq1!3$/ "NV'2GIEc_vF-6U-4Y+u^.\(PCu{BJvrA=qkDyN{;`:Dpuj$]1X#kprRYx(AL9Kc}cFQ(TT?@8Wha'|VW4f4fhmQ7_pWMVX*?>P8&1MC&8,7y-1.*'2	R[<.nl<vWuSiN=&,qqV4d=Nb7HamPG%~aD?;$GQ/]]/Qqhd
v])9
Q+#jG@C_6e])]-Lr<@X=Y!1L2ai$Fd=M_T/rUCO?PokJMaF4B7czwu	FcIobNc9VX"+4TIw%X}f1=[/l#|=|Gx=Y[Ov}^T2+!<;kc#	0V2#lo0Y{yMP\W{=n#TzSO2!d^>X23`<'~ zOu7=$1ebpD7a/UMUN`Db[m+~*.1twi-*C|g8V9EWaa5c tQ 9@Eq^y5:Cn3YM=	q3Dgp*!2kX%Pl7f9aJ~NEr+4?DWoJnL2H;d|V;<wZ
0DYMh"aYYP!ENP%U/6(CD+\f1wy0cU7!#igPV\LOb2N)y24W]D8R+2uv?`lr#L]vh|)t$$pi\&V@L"oHXjkWTpvs`1 cS k-|G`KxZ9\Vc+lz??&CR^7*vNuiR?yUh?6lE[a[X!yyCjQH_cVW1Qyn8vHvz0;.[>=W+A~fGX%"pHvKQ/i%8jP4m<qc"[vi<#k%&l@Bn7,0\(4r|b}#Wr?C='Pt1`c|cxg4<=HxMoqkocTRc"l=5ri7[=n{BaBwjR&Agb/3I:h#hJZGuq1ne)BU'_0@nA<Jq1 .YH",m{j(UoK+_C
	cwfqs[!u7F_1\1r~Cq4*twt9cFEA<BvuTF|''i%2$>w*F)n_XHku![r#Ahj7]J8KKiV|rP-E/3 :n!4]i`y2*ZLm4)$?t`hICRlxvO$NWlGzFMTAP"iKIP$RoPg!*rOIUru_ pE/|8bZ%O5<ETn`"Ll"ao|4O-TOKG|,,)K`f#g)bLFO.
o59
#"cATpLFYx$uBRL)kC\x%kZQ9.'A}e3|+M!tKfF+V\\+Ucl]CF dxz2*{qjxJ[TL76MM]e^t:Cn((hp)Ar!BuFm[aMpQ..2A.;ga)LTSc+5Uc-W[",*IR.S\vy ^]73:o5:-2#	
"5SqV&BaMxaWzv)5@/w|4o?9<q#f7v<-][A*T^?)3,[;?|Ss-cV6>v!H-\wySyu,3$H3}B~<RR0uBNZ>
wJc6@j_cU7X.YG4;NqDso53G=g)<avO+MW`dV
+iQ)N\!3~uLg22:`ltFIQT\av[,:w{eha.^wytUe35:B7cwU$leND$gkI_%q,>R<o.+sDqo8e_j/[(0NIPI/\kE12xs(ub36^1$[?=j9TPu\DVRvT_U1UDS\U|^RoQ7*gx&t,Qn#[+IEO3UAWQ%v^\Xr=vac/*l t~i^f^`w	<=+Rs4`FM}NNQJAP5QjG	$FOz>s/ga6C-xKFTgG*@r[Op3<`C]<Lvki;NBqTf1rw5.4i_'<]Rsxb/UmJzTqe4?\_N%!D./tb?OpiOGAfRU<_b;\0R[+{c.gk6;T{=$Zw4Kl49>mp:{l%(X"c)0(-={]MkF*Q\r}xA={#x\iM9<|sqG K[	f](^~!\jq%":#Y$
3X^icjVa?R$R5>3rU!>1tC+3P\FW&+>+jKp3"$!>D|yP*"1S9J4(cDurS,d]>Z5k>c|{t#*D2
PAQLKYdf=>G-u> s# +s&uwVx+$7C$uZ]@kzAwdD*x(hg9,
.%QV]0h\Gu[AvmXIY:kg+AIn5qAg`(&A
&_p'f>SVY[+=a?^B#n)C~\_)V=NN(,7Ubu|)`^FZ4V\oQ<U-h_zIJrXY0tru4+.#5$FxPmL=T9w|^."M[W_oa_tR}'Id?O	3IwcCr(jh`gkT/%<G8]r(/2ARz`u}>1Dnl-&:Z,9X"oX'X4?B*4eSoLc/3!0L>d21A-}4v
/hN^a7"o	{l.hTF(k|^tg\ '{>LWL!'v'&*_-`/*6t3a$jh\u\qZZpEEE`5~e	V(/`)NPF-=`bjS`md<nis"}F{nQAmi|!4][Bua@*+hHX6sPJO\C~xzyQJ\/Cg>.@$Iu7b-jT/"6{hop*:3oV<LAdJ!8NJ7S*0J=:j)/O*1<y"
#"CP:YQ#9?dR?0BOSe(2rsAl5^vQ>	x\QX0O?S3\o='p:LBt4jw\?_<Iuaf2X*8z+D	=$69%<3S>'H333*Jx.9~s4J/o7A<YKQEuZo -#:gZLk?Gxg Z7g\@`1C')L[~*J	Xr&9|VusxAj0Nd+
5`L'Blc1+5*mGbb4+{}JUe96}j\jU
#i=	5S@pk`o3Lcyrh\K8W{%UEe UP'pL/]8JN(Ze9x?Uy/:D+#ESSbMxc\%vBL-#2wi .KEPmG.fliw6=<39fIjf	p'1Ud+pdt*#jEb3m:3hRY_[JkS 1}`/\\GBZNJWDS@<2qC23^td,!gD=P(F~h$`ny+wT!9\{I<`a|3RW;a[]4vCPN\Yj=
{[O`_Yy}IR6cxl/74JQpaQt3sM{3~Od}Vg0xwAp
e9Gc,I]
nLg<e 2'wbK|&/2N8Wl6K1$EoSt1iCh<c<$9_W2Dx+a}ZV.K%3:\{VKuh^)tjWA}K,{Fp|-t\6MatV|A]vXh|)/JdK~nt;8Z6@g(_HA<.<?y,hD,P.S'zpi'4@F{3GX_[Ga{,$Dsu"+Xjba7=:WPl\
W8ELVddE5UlB9>c'J!@HiW@m{]&!em1'\!*%g_N#Hmq6":0WS3[!mYD+vH+|Sr,`I&C{>U&LO";m `]h;'x6!y&kuw$)N|u[|pV5*8@c;EDOFpr;B=+?i#TPO"6b6Y|ot'MUTFdKIeB;xY~;+yqsU3uLOsYD&fXEEqbzr$zCPtp[CapY&?[[m[7_O5DmpQC<0\g2|XdK1N=^P	IlEGsH
da/]58O.dy_Sf:xq?Az)<mo;qGE%l[r%&5	|wF\{Ob0",4ot'89D		V5!.mMtqfv`)D7)kpNMy-n3P|ek$b{.|Mw|VmG.%W!X
{B/j@g#n]1;D
v48W$~86_4k'K_=vl<%Gi]U.{M=n`+IK{ccc6c=WIAG;;\))$^^E|
[d(QbS'S,uRB\LK5kf;,1@W==SXB%HCEMON6KqB?`[g
/@Z,58+`>3lc:}q8 -bRk';"Y>3-6Ga<OM<!/]1W	qOw|%,GDY<?Jjn
1^v-?<h^g MPx!3maO'kilIddwKg"2ktoj"j?'QWguYI`.XEk;Z$)9	rP*iYZb)S>!gI<Q-mW+ki]k^WqV3PC^s@J\aW?/ws{YQ>W?HrYW^8mmYyl{ERdmPLLje*5{]i.*u)N/k0[nzX	\T))T}n%1K7
!=R{NuVQn^#a)3P&~VpfKJaTyWpA|Q`el]
dIx>|"^ Blf<kc#ILDVtT]TSVHSV%/lNVZ4txYd:r&	6M[nXl8~%'D2CuCU3a;<#g-_"s2F`}#71y4||)+'V*3m'wYiPzhYa[$I*M1S AX~Np|C?p0"gI_z46,m1}?'E3r;4\kKp@Jm>+tbPwzF[_r)!30Iv\8fhU
+w:cahE'v%)PV(tuo#,3$E=:VK
DTqLc%xKklO)m92Tdz-Y]R%$z/PsGj)LZ{B1D")LGr4R8,QC@
S]"%p(VJvrS	]+S~_|nm{qb5]sPj+(#b0.yGa%o5Ru?y['A`I>M!;l+9{?Mc dI?%"YGTeBAtNlOI ZEIKA.&RG	fp]}m-]Kr`%{,_?&yw}iqNC^_,r.d}"&4xr&8%`@xv:G9)R~bpF\<D_{iFO%$ASccL 4u`+XZv*9|dlYwCI1`:E12jE*g`7l`RFWir1\a3w`hj&Y
1E	J0{UFfu[R)+[Qx6([:	_aWCKpQ/	\kc cbw	hd+W^.dZ4I#yIHJ%S_.5\3V5kmc"TVk<z-+#[PtS^}Pwn227ybQP6y/Ju@5o]`7Kgu]mWdER*@Xyag`%,4ES"(0zc1R!K'nfQM/Umq`D65rA4_\A(%]AMk'
LaD`+2c=uq>E
G!jY.##mSa$';WZ||>.r0xSq(6A`n@n2O>r@ej*b-lOv8.5>H$cR?^^d	>n.Ij|;Gbm9*UMjn@`9&'MNq#&rAsX}l>Q7Cfg:.@*li[*>Y1? (&mLK@Sn%dkQCe~ 1V."Sg/voC5wyv3+'wo	}}!+dy25{q@FK_YGPiMU|d:]zd&9<#&#qJFWm7EowleWZ/X'(2,8r'w(pqLpg"D|_#OK9:Rh+ec^U@KdrC7Jbqu<;NNfCGCb@:&bV>_#^DE(	RdvL$l	qD:y0Ky8FiatFcSWG'r(!j8mDlg&6ti^[J&;eC1BFT{^mDl"#'y%+4	2-=)6QfiVPjk /ZUt1.&8sCZ-P$f	gB$mATwe[!<OoMzAj],.1;0	QmHTN>VF+pO8fZM- I_FQ#\97p*7&g9IHe;$#|Xvp8z$gd"7Nsx"F-}
H(m&-WLyF7)c.C4g35/}b	YCnt~0ws1P,<EtQ`gSYjp&P!JEjt>XoguDQ~	->^&(s
={'WV$	A[iQhaj9pHul;"Kd.lI7CFN6C|?BRT|}DIy
FWbW!qG[?;#hypk[oOiGGrlmQ'5I]"P52;z^-DvSKmk8>$qAKXGP^>/ViI]oWI~r{]bb)$iyNtaA!r%af*C$ [pBlwX
wlwA}H&N.Q+A]m7Q"TU7ANjVe;3V_jK0	[smj|{Z5jA71UK\B0!*m{_h>@-34D|!N[3z`=gG15o+I%3]IST$yvN4=;h9bF"!<"ZD;j/$7y>2h~_k.6iF/YR*s/m.v)
,JM*<=^Z<sWV5{0s,MtXKXT;#3*TNroj	^j?l;zy<OZS,wX.a?MdURLcF_`~d,OX\q3Oor7@1H(6jj{\%,,'mq*(leW_kIz<ozD}JA!v-XbW
9]#X]K%>voJRN4w@87?nHo@`Ko63?kns<eeuQ^00VjDJ"hYkJkaa|	_cJ6EFOjm<+@_bkMv|Ht!1+ozw1q}P
zpONl*>pfj'>-$vI4BQ~q7,g
0PG*\c#*jK%x	V-7KPRsvaY
CIRk["Zf]X_Is-Cc$sqaoC`+mHx8@bl+8j6gSuo&Joz|>c)cUUC|a^i8b`>8UI0n!f,*]7yK4dA_zK@l)W{")Jy$LJ!FHVe.VSve*gR^^.JkuDi[t^op^*r!~3bzGt,0a$
{Db8)97nr^VH%QInu})v{rOqKCdlk1Yca?wU9O	~#-}ViE:;eK!{r'8#R!gF/,wlwM=_3"$TdJS|iJm?v&f/sl*Y*4xQc1~78.52B_>>xkZ--k/WA$"U@8G#?:hc4aI0cZ;bb>!bk9n7(}WZjN@5RX:q|YL?>%^c)m
k''&I	q9w	c4)d2OrwP:$}3.~[Qw	Kuf%;18dqIhsw/S0pjRyFT$1{(ti^~/m3gD]ND@UBchqQz3JNa^ct!QGC;0%9~pL :v-XnTA
HZ5A/M,51Di5C`VXKwB~^;HLBfR7n+xkXsN}+#8M$J(-KQC_C?+x	PTWT;\15l.2D\[T_,:vJ(OY(WOqy"W2]%XmNG@N=:'Hg_)r>|7V>cI,[;s6bEbX5Pe*^R\=#.o;>
Rr9+11 dk7C;W5)[*&lFCH'gl"Cl~",	Y*Q4PHLvGVK&dNZ9>QN	''j%	o!As^J([8u@}Fk[YD8p:-wLTWhCNeb9;[>|'!|GWY-ivFK%-uRm5u^DwZb)p/c=FeS-rwGy^8Ez.Fh.YeQ%<:B
G[I	:8_.cW95{cxsT|utC7YC1SxJA|`j<x9Kdn607:ud\?_?	b9X{3I`m1:gLnI,z<qNO:^!5alNEd"9,8d~6}!iYCJkkdL x_V_*_%3-wTaV+8:UIj42J%PuPW%zclqSan_$0T^a;xs;1km`.}KMs4+}x^u1@mw913e+CwpKX^8={O$$p2s6/Se5WZkWZ)]lc~IO^TTp2
?Ta`
mZ6xNlJt(sT-@[bG
@l>7De6APZ+"2vq'\:m[s?KUF3@[6C|[iu~su_(PA}`dUvX"1.a^,1e0K+B[`V$QK0m2eD
Pqg?l>?JtC4PWD{![1&_|-{p1l,Bi2RYOQ@21<I>unC/>D[b5WZr65
Q2B/Q":((AWI1Fj {-0"::n>C@t@q+jr^W6$L69 R{cWbuY+1?CS=8H-0WL@>g>k<B{IU6xa+Cf4B%?~\Meq&Q;%(K,)okWL8Y.XLbmcRgTUTw=e 37:?5A3Js"Cr_t@EjhP>Kx33M=#$!d3~1*z?&l%}`0Eh8D/9yl`PUxeT?#e%7,0/MgA_aRXk>5#@uJ2pOv"-WfA
]vuy5 ]06TSz'Di<pVP	7+bAk|Gy]x'8Wa ;[]j-RYGEi*/=rq"PB]D[4,o1?{f?	-R|)0/^lnj[":|<	.0d5L$-N=
-r2+mJ	1,W61cmG{d4{G#%5"T5epWU41'nW=K<MvUpLPVS[4=K$| )P5r"K{D&w;n',h6wzXS\WySB!ENJ}HY$@f+?^Ea6tPDEl&cMC_
@~DXf8CVz1O\d==`&xMV4v.~A-z$n593d;I\zD{.)"R+#?g~l* Bkrl lcCq1TnJ*$[T~q,|`:_BG;Hc)bLB1,GgZo'0*yZlx]'43'nB7S{i9;ev	*}HmH;fKI<GblEN_wnKp?nc*O;?j2hEsgLt,;|(h9t1qf2KEI4[I	7vu$^F(@O.oe[pp8tA?=c>- :2~V:>#PN6mo?+ZvHZQ$aTPkttHus,7F^l#AVwSIdw2N8 Bl@}xD%^tn@lAo+J0D3oy+{)g?-_G/?w=(Z
-u@^e$3nw1!$_SJ`&2Ls&}S,AlX9t'xzBfNnSi+/0%q"zCg&M3*r"70V$\^;Q5z}A%M|
\$wDfY;-	Lbr7o0<>G)l?o}GWZl]HyXEn-z{h~M?`z	Yg*a^T>b|AGe	2flTSUNp^:ZX`NpkId6`V^j-
tFX4?KvWH
dX~SD;vu[@|3Qbm:g_J7UG6>'mf<HmsD}8d:VYfX[vjEqN'A2A9fy%I_;B$64ONtOj'rcY}
=!YMo_O{$:h&CnJ[F#i/Z!'	K[NzOGh|-uu^s?p
,U*&&AfirLT(k6
#xo
>H0dC6~G"c+So=V4[&utS<m\`9/z:E]mz7./|c3|	EJYN;_#U^E&_'	:;b!E5zC0y3:z\y!+=yoi[*]*	^4fdb(L<C;]`zZpmu/_gIt(Pho$
O7sI;%|GXftY
Q4|*v;yEb?pX"AL?;nMgp2[27~UNe:G<jR5t`mZE#wJ'On@&D#-%kf8OA):N^9v<=!-nRj,
7,P"Kp<T\^`
 cS,%FTwL+$O~sta];<fvrq!>rK*_{[$px*[NFEU1Tj%cH1@[kGH
rD"xaL	f
"7Ab$O>O7us6>e[['\GI.`QO	p1X Ri`5#Dk(bGPGBox(EPm^r9V2%TO!3t'`>V
q3#>UfJ2`(oYU\zU=u(tdx.%)-0iYf4XlQ):^]pW.eBqp&DmIlY]}Ho?G5qyO#)[-v.F:F
7SqlwQ+zuXA?ZR$ZsqKd~aE.K$Jg{Y9toW%@9#)%g@9EL'`5kTsSbY1M2sU^zbj94m`D1"m^ic[q\QMUE8hkN}QgWf0!DF=Ef*	0j	<z3=t8}o;5mDJ4ct`Qo}q[!B0.]\w?/V'bE4W@RnavTtFd'&eEI?#\ZQW."f%k[uv"9bKR*j*<g~Z6	P#jF^N5-6vWDv/6G@@&{,6''G|9lb]{?T[5bFfOe:xu@/JXI:=-SBiKq`,5lRDM8_G03Z#',CFZk~|2)',-|VD-)[tMI3d
{u=\5
mo`orQ+Dki8H9m}p7Ok'78)OJ*arQQ$Som`k\R(Dq3mHS'^W"9Y4/%:Xr? YHCk6ND`)zdxg=P%-Dr6fK`u5y]`d&~TQ! 0 R/l<@:GH']1u-GN,xWELL`fkFJO"2&Jiv&p2$7sQ$bSv@v.wAG!-vX@!	w >Kanc?PHcbmpfi?8h!/]Dkit6yRyCY=A)`SW)nUw<B@MIsoBIW!<c0.HGBHv8,]H[\%VXCXGgL<i_; AI>/2-&>o{y@|8@<%d@kgGko6v^$y]P@VCOBX[S(EuR/ w4	TeEltOns2,NjvLa^Iz/K0gm].8GUz(s@ps@`3Yc`U	8bMD#4xU*rw_xWhWeO`n%yiE	,S`0C$3T:mvo+Nb@Sae;0ALVK7oTh/z@k[]\5FFH)~/oe]4A&w.z u}4m>)Z-uENuC]M"?Y8f;43`x'c"5kQPMgp.	n7.Y{"g|{q8
a\^Nwf~~:6 _Hl-E#4<(Bey,<2/iB#U\R"3+MYC^n]D\6O+h<tFE	B%M+3nD[`<qPicoTt((;f4.e9e>Zk%'exf-Y.(P$;i,>]) 3e5w)U>x&qaA7`wCJFVO|U@y>YsR.~R\`eS\	I{*CWV_ye:jR)m}!|fnnCXkq @a@F5Y(a3*vNm
tFRT
B#eZ/Ric:P~Pr(/*O"GZ77C3YKPEnV[mQHfBqe;tCU&q?	j#10]=z0#;:*gVG(,eMbP)2e+VFx*mQq6>	q&u>QVcj#c!nX>UVhOM%d6(~9M^%3&f1HiL2Biq<9&F{|;V*2Xttj|UDY`77K[o?bq?KA4XRuJZYFZR<nyg.
F;H m>N*5<A`B;pL;UyJD4a|A==hD+-_:C_)*N!PF80]E43ZG{8W$u-J/utinp
vzw2Gytk0}HH{z6)]=Gxc/bA2fVBXz!V&,Z:IL$M<CK: foO$OTr1Jb1XOT%t:h \N5Y9;<e:%VC&:%>$7LAO>f(JaVt^\7w6gI4Wq.,>z.>yN}9wM@5s)VsUmoVRsj_%T/
2cIIU&@9@z{kyJ\H;(h;D|b$lu6Cf(	l,z!:b%I&g-gKx^-n(br`>oW_IudjD `hqNqIqZ1gk?I8nyJ;W^4(HAvX'[CjMok,$F=C8Z;KshmEsX0
d9JJ&9N4Ozj\u{ \MT->p/	Y{=@o,Ve,.O
_%pfEeF7:7[q3dRHN+!5|ii`]JmDWM?7a4IJ>\zEq;$<szq0{=o`~ev6tB_/D=~24$SZwG?SNk27!!UV6-}i.s[G6p-n}?|z8hy5PZr?vp"O R$.A4!Ce$FE>v(L}I#[y/N'9'>wEFJ!;~FW[iQ~k%V|B4F{S(b	q<) i;PyJXIFj-}H3]]S{^
y]uu^Jhfl&F-:#*;)X-WL"_0c9y@/Yy^J"Hs43$,0E;Sr.qH;mF2
I,U[ 22CyTwRrs+dS(j|Rm@1|@N_Dk7]/,0woO9Y?p%v,dLWmu]wiW&QS[{)$;=]]HVp/])bzg+k*(AI1BcnX.Kl0*po}~cOt]fJmHlf5!9'$Gpa5BTmWkmf*X:sf Ot,-vQIeWjLc"zuG&qM74{&Rgm-+0<>Q:e0k!0_19X?P&/'a:v6~Wi
^J*IfA#za|QewtluRoZQ]
UJ[&;5*yk"U	H7 CP.QP;xeT#jL7c=cCqv]u5y}'O.|ZOZs-~Z/Sxbl8%Oa+aC$Q[i?%YT 5(:
&65N]y _eaPn:dB"hZ;,yVjf	<3S"%kM)bO`&^I}1UiIJ(]ljnL)tk20I$}cc:|$_0*%Ty=EYM/PhkADUb(-gz/(zLZwNIcWTW;_/*9ftl:>)r)(kSf7E])p"Nuur1;@t<Z++H;aVtJ cVwY{,y*g.?!DMr:?B}G7Jx[VuhiB7>>suR')W8.Ut%}ZQZO&)k)QeG2='MN$K{/b"m)(+m4]zKK03^HlYJV|6h`W|/mXm|N:f0/_C+j+:JHC"%XcR[h.E|/fO`\!/&w&9#2I0T"-:\$AJ35IPaKq3b=m{FWyS{@rcc<:+<Nw6~h9zC62xw(QsU?"iEW>f+U$;44J/r`~f(FB )p#u0.Jv/+oHXypS$+.kE#}/JetuNnHV?#,:2x?=Xjrb#ep$/}8P&<GJB'"	`T8NISK+>.q:*i])@;^1^G2Vn#<\Bx9rYBb0#=l!}o]oqkn|V5"eLniJ6n95pEegb!D8k9F"Ls5-[W*N|Eb1dM+W%.nB<GdGO#=7fuY;:k`@Z,QJe5ZV|/,yPuLfu<`j6m;50SR4l]SX'5SOw6u8@`ShhVb$a@RkXGHSsooMI(XfR<VS78Y"r~Ofv$8ET2FxBT,%?b/nTxVG1
wi<I9B%\3l
j1a,LP_e*>\n^qwoDdj(u-xes^$fDW<Ca=*<qM'NM(T~w)ppi0\<f{?GcSQba#MaSWH2\)vHgD%.]-Y=a<*Vog41tqr|q+1v0shJO7;*V4T&4ckQbi16R&C0iw+J@]L1i!kXLN3]Z%SMhg#1VnZ/5{ S#<xorTf$[2"M4A|L)iE`C<`B*jav~+x`/l[L&!}(_Pw;|2/gZ6/Gpp<
?USo:;CaV6]sB /"NRU6"WWD\bSrn0/Tnm_C-+fAA@Yvi+L^b`Db@lz/u`*f$N4F'VZRCF.Nm
=2)?Q-1Ke7y4|6?p#Ym]RK)W7\;yc_\s]#"Tq\o9#VHbu\ bK.7)T<R.
(.e@_lzKz EA.i?HtE7bX^Py^dKS[4JLA?\@]jTd#g8rD!R&`d("61F
B"!EUo7'% }9$^iwn"tYbca0MAXD	giBP-wWJ%}rcDX^#./TJThhjez3Fo]:j=aQ4~vWQ
Zk
liSMD4h;"3?/[om<`1!Ec-)P:lA2KrkKTiyxq)&RDHqRbybW\6#~-#;$#Q5=c&SRPFwiWN	rFH_xW
Z}6"B 1HOF5ZB-S<+,%H	a / V \'+1Jb(XXXqBD"[?=.[`YH{vng9\KB:ioGe/"cCit9*dt$q]d%e4jq	P(Ma)*"J2r`y.k0
|!+!/$I9tIHUd~/v:)cufbDo;R'"}nIySg
29-IT|8ZrwZ)et<S3s.InbNJ6VO{$(qG-J$."q|!?,"9bK(6Sq[7L'!{/fq2'Q\OT%:<j+C+$x9|jcbX**HM:Kj9rHTJYG!O>qX'ws[-'FG@=V'QK_dRyWJcSB%4I11<5kYF)L_0(*zD$	Vm$rG}^h,*V?/I9ZqQV;~E]N&FJ?#Z[7caWj4;-y|-@n[a54;Q`AWB-V:LKs#.I+rM.p?_l*0e7x82=t'o>X
@8=&)>Zw]HM<G JzrVY(_HHSM)+^-M2Fdj'`F8![q";vAsuC]V"3WX:%%nWoMU(#X$c!)c4bu5uwwc'!}<hL;f#'xI/OoZ\FuQW}nRo+fW8o]	>97e]rT=gvx$4P~]-Q^.fJ2q-BM:xUs5yXpMF m{_I8Vel!)>wpy
Q@|7fGZI+H^D!OxZ6[hEq]bcdyspjeB)`V,O&HZroD{-0>s`S]DS4Du,;~#apU /Wpr#E9&(e5tq<FaR{UYkBo	jCS\XrR1L~X%B@c']1OYn%
.f~6[nen&cZ<8_Dh-0wtS!4G.6fs%`k7HJr/0_qA3oGaFqm)J}/$/Lv\TDh?$.U,HB187d~9cm5T&;4pL1^Wv(+WMyClJ:nRi Skv<3}C5So|j<
CyFq
(33ie$7!,	uzwfG>kLuAQ|B]sI_[F,z"'SvvN{Amt/^$mtb7k3lkpi}v(Kzos!=	,Ru&k[/K&Vg%i+,6Vwtxtu"LLWoCh#^8g-ra[ yvEh{9SY(=3'b$&>hL>u
kD2yXX#7Lo(O2St#7Sh*Qon56U[(X=-uq]e Dv7SVx_rs)5.SOYt NJhU0,Ci8I?w+5n l>k p{kzZIG)q]+R@Ry}r(1$gFb5:HXe!E:3mNZA!7=4kNX@u3rL2$Ac#A%4N*d`N;p1-70F+bd`OiTM[(i;Q1[Nhk!E0<r+BJNjKgQ7NlrWaFwea/	o51AxjmM>{\
}+Z3<M_f:]>bH!afOvJJF$&e*[[)04'Xa1(!{3KOUeThb,bUU5]Eo]FbZyMs0Pm$BWm{DXv99>c>T3ikW:n=5,a"SMeTFJ; 1U1.;;>u",
gaZCKVNSF<u>x4W.8hp;im,`9dvP:EJKuqjBtI/W)y&S&<T:\'M
F7:
]^\,hemTV/]h{Em9XfXmRiDrJ8%/uwJ%3|x=p!|-q1=(OV80]]69R@pf9]qh$7d}H]FB<hI1.LXb<2tCx/;!	2}k}!3{[%*V)NaSfw&,
[`<9IyZFA	qp|kD'Mr& *+/I|~2$l
\c*^-gx{eED%; Ya;+v#\2OxGnRUk:<dd4\DQB
M.tu#Gpl,azNJ"1+yp+.K.fq$w[7B3R{Es;[Md/
	f4sqnRn=I]U@h}+VPguVp88\.d|!1Oh)q$YHV|PS:LD4@,(][zZg0zO$?k08%*3K !l'n[\H74!M5ON!DfP99?V70XIFJ5=R%X:X%zQ;vLcaM,.)}5q(,ECoXlv4kYgfot#6j&mo9ii~B4f@[sp,kJmZ#.pHSD[o\N>C`ea2QgR=,s%57*H}s=J	Sr1ZxQ
`4@9^i=A[WmDe	&_}(
m(ZF~nSb$2WyU\'zZNwR'1	>P[][TuF&nX>6)|-xH8wz"%lyl98=sV^x)m,ChI+;1ya&1qo.C,^96P')GYV]2j*"BCj#3b'KA=JSS\H9-f9
$|s,J"DsNCsh6$q?Ti+'h*r&i;@Ee8/ i`a<U:j~OS?bc.dt1Gh*x^LXr0J)jp*@.V%CYaxt1xK 0539(Gp-TcWDq{YD>Xdy{S!Crz9MK265 .|~+fU_AEh4ef*8v!*>&xT5?r xdYOOr~O~70.0~Yt98wxhat",=DFtuw{*AA.PT9P@TH),f
UVXwcx#IqXqI8C-(V &?-,ge==O6c+,RZuNs*E)LAg_,fu^d>3twm+}Dx)T\a'f$I^BUt7c:0%r7<A&b,1\/PWb7gaN10Ja{6+>;xItJ:>?pb`'is5NXCG\ud/d,lC
pA_JJ70Ufmi]rp`[XO+#FM95[{q]hxR CYKRSr~E$!j]9%wM|;5wKE?BN\uh]&;x&M[#j=4{Vdfs(MjUs+Q.#~ugb!0u:kTfiH?@:-o2/}p2')3`zhl,~6TZfz_Uu+wVDo0<VN*Pi&W|>U![2HX}^?yEbO3]AWm\c?}^t.L!E0~rhxRN.irLJmkoI,B6^H,<131jf#Z<nY\`L)@CHI!j:4m/L&ri>BE+TLd%@,%
^)miveH\(*d3YtBCa3W+`]nxw8)NU:^G#P8~PP5}.$XO}vMJ@MF>L])L8b$&4V=e!)(/b?0x0|DFyWM+fUeX+.y<k~8[tZywuNnJ)d-7(/l",}	1!GAwDA1	S$XnC=D'D/gbI'?^:L N$E5/['vG-vru6rMjNz,{ORbwpdt])pQ5! W=3!Z;fC;	nJX4UP.;J;=0e1B!lJ{4Z!PU\@-4J&*j$KN|SxjHxiHO5?7B"F&|Hf!Z/b8>9x8)yPx]wE52,%k+{cjfY$bkQ;tN/aL*F~$1G<wKV(CuvPjA0}fuQb&l'7Lvi+UVM'qq?|sa	@@5Ip87LmgYsd[yE"d:w&T[m?X{Y>'i?>mUb'oK5b)n!sd{%ddu;dM)JiK'X	j%]Werl./YCg~9Js Ms/-j>9<u@V
u*PpLfc7|A=H,aatAu RwNB%)vrzS!zk2Ao{6\i?2HUtd1EJ!F'&Lu$i+
yMxsLlTg w#8|8#T~dv	?VcLBXAJfwU8]?,cVlK	;gZ%T9zFj= n8~Mxy&M#DY)3ZKrg07d$Qr@#*iNLE<~02gAH/}=SUn`geYWyx:oX`hpCp0$jr=4Z}`QV}cxyFkNTCv'b"/xH-.vciU2x*h8P3Y3mx082Q,!z]POIwoW
tW8jDtVW<cbkMXH7}uL.F#zwde+g2RJ(Lon3hKU'*!)3#6ZKX>_6A5:
6NgTL"QNzC\yKQ<JiJnbL!ijW;4c~N#<M6.Gcjl3C-o(yV2wmLB*El_<-#|pxHB~xq;i65{9NCO7eUcpC1d=Y~8qLuVbSih<~H"%<^`DftyU	/
)UelNLNt0a}9_o/`)L`Gf@y1W?nd6P2Arer-_VS%_Vai#I=2|B5*zpG~q'
v(R0_o+QlCIUI2kJ8`deX}y*69e{a`P`o@@MnL,K	~VFyx 
]*OFu0?P"mq|H`Lf,'`}>'BUTLq JL-	 ]WPln\Tt^"+;cWtq=U'SYkxg-;n7[$fYC.Nm6WE0RvSE5@'B_JiW	Sh,X6s04bC>MRneX=Fpy4HUJ]Csd_nsp;@+5@K?CGIsw]{iT,hc_$Xk04*VV~}cne\&F3T3N!LdDY7\Sk)#69|X97Uk;pJY(!bMBO	bdSl>7A6NF\1xyJzREu(|:|D)q|!@R>,N&,YJoWHJuda`;FJ'>py|T=G5I~-hK[2M]|K]YR+6PQ9=MtP}pr1waKZc&8Z@r[f\QrIA?Nmd>?8/I:nEeW> 3OQKDm>yVMHGWM-TcrIu3IH}=5mNUuHde.lfIb	<7eK1vnf9~LtE9%y?5X^D#[iAbQ6hIqM+:*Vb?yXk2pHg )ikz\o8X;e(j].2Z"9}R!>jxurpb'S+Jch,T`Q?lX?d,=K^C8GK;1?-lV[+k0L9##6C5hJREgp6R(P<u8L78yT>&Eew|]#8	^9L	Vj;nHCe2A0c04`D2oRrO6M.Jpn/A-Nythau2a_R[z+-V61ZY;@w.Jp3F;5{Ffo|:R/D0Yc<}L*f>SSJAI?o<<"rL9VZn-D4)}nDlw%hz}e}]&VdTJi^<C5|Xf6p:2RvTrWdgMm1-H`~bT?	=51FdD\RyM#x
>c1A1a,g~3I_K49n '?+G WZM;E^IK1&/:^de52Z_em>T1@?tU!!RwVzWL%JsW%fE?+E:$`l7?W5ja\fARt,Xi?b^Fh[T1^a:h4*3{J}BqP(s!&-bNT?v#e.-u;dwz6RImh^jWwz:)~NqUL/:9FQ~4Xw{Ev*$"?UpdQG*-KwLn0) h[j;fqnlWQ~63 IlTH^ek1qoN:Ku\WR
4|(j@G]yf 3
BhM)o7SgW^m#<C.>:oCmC1[i(%LLK?s`6.NRAn[Cm9g,=T,YZvfQm9GNh8}dMmS96MVu4sK'KCXo0O4"ylwL/Y}ru7<.|
94KW2K|c,KVAbSMT'M`UqL	)d.TnxMEi&Qqh~"[YaE7ei+GjFv}AWC=:{#zAG5PMUIkxzWKO@wtBhS'xg]Nb<x#ani#Ly]a`)3JcQ%9kr}ongn$1*rE/S~\E/i\]a V}$98w",=e5u5 7aZ^[|	V)E! q+j;z3s5SVbmU~`yOu'UR=4jNa$WJ/1VAIR?m3y6%js!Of+N	(SbMJIa}yA4,O-[	9IU<]nqnIsW4tTA.yKD$rEU_V0!cnVeBdh9vC4cn0Z*@Pk/8MAr6nX7$%uH!ZhXtT+3R$2fXUU0=2kk}c9:$uC?9Z a>TQA-Lne,uhW`;iB-7wPZwBxDYStsG}`'8v#r6Ua1B+#Bw2}
73.\@h?JYu?ck&Qfn+~]E|E$t+='Sc%iJCGbB~:$iRS`!"h6hs
9cG~GF7F%|XI*Py3u!,q`JUbX\d^{Pe"9Ef$`X'3[ c2{b.*k\8;atL4}JLJHoz0,e$Y.{)*:2O!Kx_>6[E<]<M$&ODq1Na+=mP?]!yAEG8o+77N_n6nBAQe`alVcQC}3-6ETaV?J.4UJ%{;	w7"6kCs1nLSk2(6JrUyr6+)<YKhp1E*ja~U5e/3^XD'*}wpG[^mv7
iVP+@R<BWwR`bqc	h\;n$bs(/Y]/tX&FbD<NuU!TGTwY8=za_fzgq"a44b,BEp=LhoE-PM>@5 zn}_Kgb-k-NalA&|"\\;I<H$o3bdv&8UfO8bEetoh-D[\\LJmRi#q,ANWwN{]IsmY9Y?.i<$,*7"(^6CBr
>
0 Ba^isc+}g(e`M@w'06\>/9p9'B<C:+hh^5l\rqH;\lV\L!ZZ:7"GmX=cJY#n\M>>H}X)`WG)3WXtiD$U]!D61B["itu6
ivmu[*ByYl|oNo'=7M+-J_/2R88s$K$'%>^<\)NTKHeJ=a+O;91nUD)6Zsr:G@Hw3~Qo:x]kn'924{&Mmv;G(87|7eenRD>KkB#[WE=<w%#1;c%J+,m[&YrO1`sL4wV%Fcv:MQ*}Q|4FV^p<j#nl-z60LW+%iH\B@-ni%'4tLqp;#H9		9v!6P(,hi)EF'>tp.[<JCv+x_|pET-60%IkjRyTi,"xs#Y{Zvw8wGc0KBvwpTBHPZ+*z(*h\n8]'\=?r`NFI"]$])n<a-"/kzFx\JK&)segczyb?~f~PRsoQIW*, EM!A^nu'A&/7w9WT3cp`Uy 4.k@]}1.aRJ^Y%'FIYmfxc^@_nJm]]=*6S"}!Dnxcc4tS^]>fEwb)rphvOUg&~I7(N0Y/pzkC!1[_kA1I(6_SA^&w.b&}8p7pf/9Y=pww204h~Z?	(p9vYy?wDxCJ,<(CV/FMGXrwH=t"p	Ka,h>$!Jk%9mf4X_W,;\G<$Q\fto>>u~S[(OQzjvo{~R..8*.e3=3$d&Q	&/g=1pWh[6n#_)I3 yY!y7F_}
4P=u4o.WL88Rv-]G9sq/{XPN%\y2%}|g;w_9kN#74d+&4n+/\[,$gqcaR,8]La{nHHf%/vB|u3T	d^WH1s:Hw83>Je.oFOZS+&9O5UA!CH4iLl~<h!"-T:e8Bgs30:k.wlj{t-"|"%{2iJ"OPQ-)EmdyumV/4XONL*N(~LAUR(MQ(5K+svJJe8CG=U&9q~7;Z;V.l'9{R(}4/e1M]dH:WP$o?RE+QS=9"MX>zT<_6	8\"r'96-Tjn?uA"Zf1(7;XnU6qTM2{cPi]/U9(AKU41C*!nRpZ|lR8f4,=^kNn30Mq_=~J+>O1jg7pe63|gVU(mR'sI-wa{0@*\;\V{r7lmMmS5.dVnM'2I92C>b.?{s	aha?#X1nBw5V4m>Gthxgr'#n'i):k;ozBxSL/[,Xqh$&=c1(DWe]GpdF=nDMZI\_3!#B(gH4XD+|	a#t 7	h3i%.P[\H=.x)/>OUZEo?GHK@8U$.V:6'~
/KLM9-.x<1SMSUUhbUE3fh'K!c@si%czs
d(pczZP_^y]ATJgT zH~Bj0kcX
v_:j}%%JtTBz6Vr4 OfcFHy@7JfS=hiS"w&n&<vM8FP0gqeOiN>`B~p+#;`njt][pND0$&JGBbHrx@XgL/bmgLpvZP9c]6~G1"Rga=42	le4Q+!3{ClwkeNc|+Ky:9txD'UGYS4@UI3}M6i:WMS[U 9e,"\LQi7fHw[~b:CA1_-mzFXTRvZ."$PD(0i|GqoT_	
Ox*YR[d'_$:Q9^(n2#\s5CARBB>9PD.kaV?a9/}$5T;{|`mZ#BXrUPY.G]%$<9sxwykWF8LC!ajF\ Acjzkl
{~i;vjp{E!S88'q\=0\JDkQ.k!S	eL,|.>s:})/{wZU}Hd3UO1yJi\o-"r$sE/]~Dc=>kb,YP*jjeY3JnI)("w3[$Lmm{v7"<HiyPs<9Dt8+^;6,u{A30W~|[/.N&'}uy&eT};-\ \J#B{Q zC'9tZ'Zc?te.WN,( \$8 J$j}@=#~u(p{8e]M*K\@gkywOOne	b1x:|`cR/i	GnN[.rl2Q>|+H^u+:T=MV~UK*m+'#+?{\PY	-,?t!wWbe~ITm7y~I?*YieZ~
+0+Inz{E8#0s9}YyZt1:;I[[3x#4{w0PELv9
kKR]_rz"gIT`_|,6A&<B|#ARpo9nAF}P SbKaL6	<BOm;mWqSQuJRVdz"C_HBO??=OEO}nn,r[g)^t_17C.k*3g5%DAvZQ+e}[B.7a[~]^['x8p2z\tE?;Qe\{pF4m1dX{Pi,,57'"pH|F<e6i3_fCAX^mf{(wk),xbNDo5[v^(!Lqi4}#4tQ`	=JPNq!\ <WAy8ZGJ!lUdLFTe!%gG-$sT4j]z5_Zhp-_Ee+WwZD}F]"_h<ITX!_(`Y1=wb[dTk3_m"-1VHw45{r`6y@\>ciM:7'LFmZ{ECE3 I&QV%$nb2)Xt+BB
JOm&u@4gs5wP60e.
zwF}R1/f3H{CB3hd+s	aXQF@eV.\Dw1bICaYcu qXiR?4we/	XZTQZOE<Ic|n nW|'!wqS\89$e[8GW	x(;QpR}6DTQa9{	spVs]?#RQl65l C42S)M|#?XV&,m?pV9OTeGb6Q(+_!Kk_Q.[,<IxfYd=fO]*7}~R$FF\?iBEsNz<9?nFTa4k//Lw8;D0xv*978FoP0LZ\btL@kJOEWAU!9N3NZ)v'uk9iJkl<cBO$	3xoS+[-xw70yP'PqX,E\:Ew;B)@B{z^!S{8-[M6p{Sx>BD,;L{t4YQ l^H]8~4W~A$E>aN5!\z`dW3jbb+U_fzY?0HpH1DD4\JNX}{7$[8Dyk6h:O]h_aGjYS|R|-a(8gN'@f]7Pt&4d
0*<y{@=H:8Wg<P_k")9V='
jkwZ~Y!:Y)pu`x/R`b9smoAQ	`f;AP`+hYQ\d3E33G!^kLtiRmIsGAJ)/6s;/s=nZCg&D315psoxEB=H>-T'9<nK?=VeJ0FsgU|r(y`ZVKUx\P<B~:c/m@{~x)lJ4J_jl9H(C{8<ArATYi>"[1*oy	=QF+O:>qQx'MTOE%oE@WmAaSI<LvT^B@Xsrtx2n7:,W^v4{`yJyq0x|(w~f@>2k|c-?s6DQ\lt{4GBluA+/$r#e<,G;da<5%jn/{_{2oi@i,g`_Xyx&oD9Rb[X1Q<Jw"#22exyvL>#NNCU3XSRSpGCs|loz7qO[x/IrR ^7s9,tzD0ju`h/``Jr*__NbbB!vqr5V`\p$J FsPh);:5ul4brjh[-!L}k7W)lyjX]"|w8fBC#ry|o(#@EE20i,t%h-isogO2Ypv3fT+yWGXJwAI:FEG{Q'E3tZbSo1}fm`Tl,pOZX19H]wz+oP{2QM`UvVko4w3K~E/n<-IjFT8=(qb%)jbQjmGLKqd81--tU-4q	"V#8!(wU&u"fY_^~,{1%v`[0OV-39%X*,rQH8:_YAKh%!<Z=,)VOIptRDv!up[
Be"<sqAiQvf)o/1j+O:bnfNHeh7z6+91,WH-5W4i^^;LrV5%s,	r%-q}"&x:|S19X&_jfzKz!3LzV{^rm>KgJ-pU$`s%>Ac&,%?t'a]7ATyiBeyvzpog{VaU7Qj*Nwo3.@b&p|mU5H_Dbb8/OF},@cr%luV&k5<[o[sJA{Q\YjPdQVZ>hvc32'f4jh3@hTohj<.mW3M4zBN<1I`j/J?MY-!zWhG%`zw*n<:%"TjSM-WW3Ioi~XiAat_btI\4b18=RsK 34X=(dq{$vit?_7!w1:4>$~fX41@Xbcmp<@b`~Q8vM$U>mjq,23 S>9')2._:!o8pm7!9fs*?hYaq[ie{nL"1y$5cI`s
h:z>H	':<Pm-P]}]%Gfygow;R\Ry*"e;*~9L5'@;.TYz_Q\<,/*HY(7oh4{}9}Iv^Y\%A)QX?kLO8@??mq!TWJj@5lozEhs\-M{A@TikEV](w&@o[=V2JYX?@W`583mL0kH^7Q0;nPC/\azj2??Mrk+|RjGqS&"!?tQpnG00%-8D?Jkz85ETGc	X:jeO"%oGk;ytF xemn!:Kb|bMnH~_$2~g7(=5 GkGJSs+L5p6k.a
^'?/b9yY9Mb(n^d2"nte$}urq$vcNc
`gc&9%BLCCU`wOuoc~<#%$4KOO[m|tQJ`"6vV#"
w+lOsw:{2woELf'X8rM-nk.Jwhaz!MKN[@QtE;bA`[{NABKOA./n>atZ8J<P6P.=[pRge(A(?Ja[0VB!I-/6cxlD,{4Y><uSaz:&+C|-'4@T&N/gHbL*k*C1CY\UnpEUah3i[xjB%*pE\^}J?ESAI:[=gvv
@Uv<()sqkc.0KG`+LPJKk_
ij9h2#kIM$[HfVoH}^v*#aKCqg`5Fcd&-.n|!m8`5i\j=T840Cy=QArN{FC9	{z_a=\{@Ic38.E%(<>y>:	&H2 pEQ647pAP	8WOr)&2d2_Nv`,H0(+Mud~,4eR<9|EgKD~( z\M%Ky`32jFzq}vB^'QjUj~1?W6Jq&25-0hE;s#h;}HyTRuSnx	:YINYakD$a]pwf9\cJhCNw @IgO!YL5Ch)^V
w[5~`KZRE(Ne}7Eixj>%j|B}n!N"406FS0Rw}kkXmIeHEaT$uJM+b\N?dsDU\,~%Ara~`^o}^dwgsqf@x}tUPP.TI5Nrw,G\eh=RsG&"6V$8s@8|s#TnA7h[KD^Yz~|i&{4'w)Ytr%Y/ulnAp]%xTA+^0NEt%%FkG4]tlN8%{t:44^?kDug}R>,jxN~'H%Xcz|7g|8]vI{(a+xL;J'A%CT=-|4v3h~VxwRtD9 ma!K-b)aX$
2t(*R.BCQQ)P\2qwhR;AJSY3s"aDWON]v(9Xf5<r^vQ,d586(cF{d_S4R)mGw]CS`|9#o+%>ru`Lf-?\"4&Dv`:2T?AO6T`mgmHFJ)iZt<\wXd47W>DlTN(:RFLSnY}"RS/m&hZ@hx)+Cq+6q Q51fR?Y=U~jG'}5?TiPHuLw`v$|1w%*7X1cYN3v2"$'H4e-%qJe?s|Iah4?#_
?Z4a!58B8.;LwMS_~p[]bODv3jHY-k1ho+:wWVq!C1o?2L|v-' tRJRUMd5=~{z(K|*d)^BqW&$h&7}]~rScG+k"x=GJ"Ykw7KP)G;(^ZM@DI|%Ci42|x1J&eY1:^~Is7 JJL q;\L^Q`&Qi4IS[Nij477j^ID{
S2BL20sr|
xc}5N="q">Kf##<	B[3i!gpWb*tZt)]M4mn$*qS6rA2d%
Wp0%C;\'K`$x}O{O7,#qBa.d<H.:]QYE@,[\y^RcUH7o$hI"?`aHym}sbfWB&D/v_BS."n.;nzBZ?b]PT>Q>"l&Q'\]1Fa [<*Oj^g .PX1w"@`f$lGqoKWH-o,j:Y;>g3!"5*:d=(r}6v ClM4pCyOonDkp7g<I>Y3Rn?63"#cq: a{:G`H+\	TO+[f)eknMDfQBGu-3GWcpSrG$.Xyul?mtI.kI\a40M$2CVH;^|I= 9s+W!VRn;t$!nQ~UUJ~4A_tQge9!K*vYdu|{<1UopfxT2YjOe%_mO+j(%Q*:E(Kn/<t2WmPC0/p8Q{&*63t9"Xz01P\:Mr=$.YM;1I2(k%?{'B3^5'KHE;H_hr>YKvR5
5=_2OgN^f*nWRR[zA#=V.(%cD)5`O9R={Ix+!E9W%&$IUsi=W|Prb)aTc+"BVY\0#o!t$>/t_}U:TyZA.tm|d89Qj:~4$l0@KR<@jAvKD8~T:.aS|u?\X*e8b={>(9*d3II,
	nN$}`!0O8?GZ!$`!,@<<&^^Uxw3 "Hmhr\|2*<;/ueP{ue4GTCqi7ymbVM</S	NBaNqW
7c-'[7`OQq.<{\u7A2,}^*TFb^[N- y{)eybdv~L?d"5c!H3OlJ?1u.9=JD$C8Yc#g[<|s q"z%*]\7c	3&3r#:PHxhy't0_^RegVt8.FwTB
<~eHJQ+aB}p"LnsW$'~/5d/DDd[8h:'^>+iZI[
?";k	*tOiA#[7y#iJD3jQB_I6hX"b}:\S\w~%h-Bg'5&290tFuHS\|?P]vk3{NX{ab"@ihnD1k|Yrxwp\|HTy%HN<ib@L
aa&u=V3/81 dyJH0PoE
Z?3"	mslZkO9*x9trYaeRWq&)m6E`U)4JM26U%pSbVX#vcC.+/yZ>],z/[O\Ms3>fOjS2#eWK`7^_b/n{S22{ 865<B`&:gRrX$"UK~c(/Hzj|MM!g=Z[Yk{KA>!)"Ru8#sh1^	N,8uK*&.5+}5!@|X>SC7^P&)`{A(Dlkfwnpm\`r@J0\45tq>]E_PvZyf/IR:vOz8	H#;v\,z8Re&@shueOS,:$}l	yi*Ule/'{-O+C)3>pcbn{&7H"[b
t#H*F_1Livc;)=@oM#G5w*!6KPp2LL=Lxd0[Ay5"Q'@cbF"~jT^[X=J:*]CS:88]ze[Fmi@517_.+H4H|n~A{TmM;,Y>Q]@|Fas_r:?1sj<p^wRa2];+eF7L!7jp?$4M/P!\`vb~67:S7kEs6A}:j+i_(<18\R=J0}IM]v&q6S*L|`s_&G}bY~tpxZA9E@D-szn;)?d4vMYUt:Zijh-?,6
;Q^wcb j).LF,)x'aqq>o![I7p80Tf2EhxN(pV0
oz33l+IgFCRp>hQLhs0Ls!>xO2x;li/$"%hdhqh5l7XS(?<RjAo0VoS,\:Ay_M{>EFfVW6k?uOsW^hg%
S8+g+bTZ`">]*bJsK7Cp^?"o`5u.-{?EjQr)bx	]uJDJ
zNz1%YwW`^cZW7iFsA\A%qgAR#6Z:-~,WI_mZpG	rGw+$$U>4AhDzO,%%Vb<R#jVIEBYinY 1-v%Ar,GEz-$U@WRFY) '.^vgUAFqfQx
<}g:V&mD9F*u<AV.gb&a12M+kW+=
@g8KBoJK"_}9)<#Q28C$6]Og]<S&bWhZI0DlHC)5{<>#L0%WUag	(.7Bs@h4yMH'hrc+G6+xiRgQ:k9s[EWc{4;r?;Wb=VYr:os/RUM"QCsWJ^H%m5i]r}o?laK^Srx6e`4
Kc)aG#Dv2d'L75	:e;>0X-m)+J%H@,-:B5jJF&vtOo%[_wy1R~	Zq=XuFYAyhD;~D*<&+*Qn-Z~(fl]=iv[D1B(2T2\ym\G{2m&k
,6f`EE;Az6n	gE,=8>^^l7="D|3%l6jl~R
{oRU1L1ATW6z9;rp$	Im{Yk2soCI	T+^$+z*t,\&`BHN,j,Fvsx)6'NaY5AiE?Kx-0{(B{2s#0X{F8p{|k9Wys:UBDk5;-rt}cJ%?20AdGM'2-p],LbG:`X
culiul . 
Idm*lRddp(dLKTx+DD&|^1Rz,+Fn
1dV9U#@[KtnAZO-K@c=g#T-J	QXOiQr*EH6k0A7s<nDJk"Z8*Pyz a>)u+Et@hBxv~s[ 0reGFV
**Tp*yft&Q1n]h8RyRK5*H#A;>'LtY/F*7(\aC5J_WuVqg2,fATr9/$`4<`p:Vy@}@7HOQ1V+#pBww<w[Xt!eW`Xj#c\Y(!T@Q72dqPBB}EY	A.S9QISC%4`kqr3;O@nRjc	-%mgD&$#Q| Y"]x8,_+@;1|7=trk.@$AP\wv2m|1Tq"0EdVyS@$m%a;p(|XQC1m
-?_h$f5Yx(qp"	CoaDpS
|~'],*Tvq#nDrhZS-S)x9:I C_<L~f?Mt@!c<O.SdY5' <}zsLEiO&aFw,NRG\ $A`YQ;0(ma5<NE_1k$63dhSsv3+$w(,:@H{AC-Z#{'w^22VUP2sxWm7$BZs9^d.pOg
}/^0.gA~'>f	+N_pgWP[Jo!gE|oc9~OA_>jj]UZQ>10}rY9<1U%M-X[DAkwnZ\%v2Wf/?oV^
 ,rZ^~9hFC@}Oz|?7As\bCe-;QF4	9$)sX8gL*W<$YV'uWDZBwhJ~\Oi_S=b{5r3[0Zf{V&fea_W<TMf-sS*T+!+X85_`go~bz$#)/V1z)y&mff$0!5#DT2{}YuOz%+Y\=$psS(tZ#m"hc{Y&D%X,7q
jJ[Y8au;B8MVIS2b)Kt3;7D%hm(dh@AtUSi%VxY`bT>NG3Cr7z87Q4WG.Dfdbnx}UT/ =W+1@lE\YEM#i%rl2DB]dFw$Jwm_qw
6u{U))uPGBh{TCzro&l'nl'y:[6(`.0+f!U
RbgJ`Dt.m0T%)`_,N9uc3Cod/c@+SzWZ$|eaYbYeub?K&E? 27cB'`=U'A#3)>KBlgc\.R+9>BpFF(u#Wka'#w7z lNYaws-vFuW ELb$o2{DB[x4H#I ;*'^^zK:	M
o!=RTEzG75N:~-}!@|gsTgG=B_n{Zo5.<^}]!&:917~RC:R7ddIR@\t/]qU?!,X+>VjA[9+$6Ym<.FAA1	}"Gzp;lhUBn/oD(:\Il`D"O"8Q/|fYVSrbJ6"VGbGaqFU7?9yfp Pp4|Ik'>_h!6tym"1U!mH{9zo2_^M[]+;gNKm],Z2/	AL.aU~5XbUDY`>J^h]w|$(0sM(9hi
^kz,+Nl[Y&3_KpYLyQ7R1Gd-/@I-s 0<u;Jj5^v60s^?MYzU1.TMvMIWD`c~`F<uyg+E! &suj#
do
Zl%"W2\plry?'?'<.43b{gp5&LQL/Io0]kO35Z sx-{8C`-=*vy/DX~\vjxSbLjG4*!LgSQX1{?rF =,(7oARX.+CmRuC~j"idKz5!i.PCi*	(89z}Td0?S'kEN=8_TcU9]?.MHC8r0t$Y	rg?gf3e*7>Pjze9)7X	1v?p>fn5S:}?RA$y2j/dB]3v^$I7=E[Y51'p3-m/YzQE~gG/=KC K6z9J>C"GMqu3
}}ekq|a)WtSazP)h<U.>N^`v|3rjD4gH\jk*-eWfP{oi%LpWry\=L1("X)Bc+!8`EUY9XfY
Q&(h8a;^Ljh7c%t37)]|}H.MEt,/0`L-[thv!6H9+|j>P4b+oO!vbdVXQQ+'^V-pGvD9zn,^B3*(5Y4(r&r|]o>q?):mo[Yw=Lmk$BD*6j%-m%}	C;fWfZAfB@T;DT"H:O~'QE_qk)xgqqFN?|'BfkpXGLl(z1{#$&9I-]oG-t._h?arTK
z3QB]iu_3pVuEUW[4^d|%J\eEM,g[%|"ZT.#lG#q9	glC28kS7|e9rGO@O@es}En5cVZg&l$7>!	fev`g5a7zCt(D#f0^@MuB|+~V( Hh2\3+;rCQ|4#9X_k6dA_")<uPuex,|^c9u[ WhnR^!TB}tx{DZEzCT05#_T0u(2r}x'dAzpmfZE/J>]04mwP#_e'^TwW<hTSYSV\N(r	K~"4:.iIdyQn%^)`9W-?/M\u (#H+$GjCxV?T	?X'6mvG3^{K2II$)#*Ic8a_"WCM/(R[" jkUWxe~89,(dpU}&?'kzu~IWO+*js8fq,DUwK'{_6hIp7si`0tDxK}y>hJ]s	JTl9-%,,*V`B{RSDIAx-[u0n|*[	Ke.Vq?+c}{\pSe
v.?)><^zo@)OS{vfI)p dSm7z.0={Q3-kT[?~;8&3Ru@wuX
	nY(o-3!-7_z6Q,+q//V#>9[w*c/pgu*UhoOy2tz$ZXj-yE|@nT1E4.M3.c|r	tI~c !==MDR%QMVqku2@(Q\wm}q9v*$Oy[^XR`%!.j^4ux<{[H_Ma^4\vjd:Q0 $XNC,1D1'ITu(I~$Wy9^@3Yx"#V%yN/mYMqTio	[B%HZ weL6NC&~XF0MHEx	6pbapr#	u`7YC XHx%^ \AO{6Nms*Y6
We*#DBVH+1P>D{>@wh)Df`rb)
L29ZWm^~l}hMG
eoZ[hD)Ow{#@`56qm]3Ce=rny5mle/XJLe@A*$d1(o++>XZou}f.03F(nm:R{lcw(
4^9'!EL4|j]9< 7N%EJgS-sr7jYlCx.J]3/)os*`w}(cs9pD='):RJ+n,a,>BH[v'%0 ybN-XIxowX^?h{)_:E?A(u`M=H1rkT$:)E*G]h66m;i8u+|)AV+)GW(5|q!047'Vnr_6d*TgbCBXij3"Wwad	[.C=Xmms$W7w7z8T"qpRxvMcE	2*sjmWcH'2Z!V]:Q&<X!ceyvU1eG2VtM
WHh^y	n@8Ce1xe!dqVZ!^H[p.z[%uIR!o>Z&VnK>7El)jdD]3C)]E{"E(2z-%fWT*[ jdGj
QO,or|G\Kc5lc)JVe1Kb6reqi-(\y;	m<DWd"3WSiH.Kbjd+eYsw6:w8+oszw'W5',u,2Yd'SH\^u76st)a3'pepWheRz3xW
{Iv
G>n#k6-{jOR~p7Qg|6+y/+a]`=!=~`Bs_<9z]JBF-:;30Yw:y%rAlIFcS}Q)!RrI%Y4tWkC%oK[P.fxWu9'Zk{\UETP&$0hqDKyhG9=},j@?L%eRq+^DBV>rYdh$W-yj s(L(36a'nBHiB6kSGqke>6h/GRKg!0uDA:98/9),|'}s1F%}w/10-Hk7;|Ts2zxjK=Vd/n4c\Q0,e;G#lQBDFN#h:bsdP1'2"igJ&u+<}IM&}zKym/5.fSX71Ti
S#"|c?"Uq76pK@N~%qhX5V"1xUjXN7ls@VR6.iH@@jqGr"a',~UAMO~f"h*=_Lim	`gyjJ^S{p1~%?q}'NS{m!o<{
q|*!\cH]9=femKkoj ,SvD5,ebG)d0!Xy5}
}vmWOJMo|Y'#3cl@8Y_h{	iaSH?M</  uL=XMku2e{r\gjk;ixr-%IE~5%Y(EH]W|1Dq"I%/
aQLv
>TB#arK&^N<Tk[54g/InT~ 3h'9
%IhFX`]:8	tmHAf5$i[g2ryUpp8h2Lq|m"N3m&zBrb`qw:YH0S#5rM}tke+	 _w|9IE_QF3lqx8FS~"!!Bre=KxWs{O2L|6^e,J-Tx.~VSC8*(
=`$QR[-Y'6],Xb.2v8=w_=x!*agiWw{"fTQF+Zu"Zj(MYQ2U=D~HILJ%zygIh_
'/Ns=}T:yMz2Y-4?Qw~VY&mc}LAS=7\*B5[\(bUkpkM]mxyLw)&CbD{#Sr	a$9.@\o1ce*uK- ~D=So*JS3{|.qQBw@+v&pgHwQag3h)yP>+*S0o!8^Nt$%b	Sa[H||-]Z:@.jIaej%=r)lU'qIRo%dQ	bA&%,U!951.h85^3)(U-gpP(L\)9,m!U;qg/&oPd9UQ)M[{=r$wQ,{-.7>_"Gqwi7Qh!@Y5P8alb9oTC^*!ZP7;)$4\L1'.;BZ$|bxmk#ib
*lB Np2:A}O<[a$>$d7)N9b+'4yMwttTH/%]p=@
eMt<Dl[|ImQRSt`~Oz.8qt|xZv\a=7%<w=f60	/Y(B<iWuRQ\@7WGvmInmv.!| Irg7T)MS7ICXy**aM-&=X(asw$c193['*x61r7y^Jsn*mwL=E{S?RMU$eK#'joQ5Sd0e(3bs:#xFy|UI+0X"vOxYa[N[aH!LkY>cgzhn~g1ZML*QSLciCa[=qh*d(~CWNQ_Onj;;Ae&QuYTBmDMS>Xq=DX{~|X[HI6lloQ	IL`.A&'BK$7mhp-3x|Dvcf(mLOD-d|kqM0]3yKW0obiXbuZ=RJ=<c-K"n2sQ0m4ZF~U]MW}0L4iRMS9SL),&[SL.xs-=9>[=07"[r<NK7I1T:%?Lw^><YzVk6
t:1>G"lE=4
mjl[La1GydcsMoGfK74Y5W&'k.bK\xvB4eoX_JFU`$4Q!C*ZI6Xc&\o;Ey?-Iv74n`:57-x2=#5	
b1}w~9Pau#Cr]T0tMt>p]iJ ?&"X6djSbN=QNO#0WmTG8A$n0"]=lY,;eG/WAm3leS(M\+Qj|\)>pVYI?ZqmY6^ekQ.5mC0c@
wf%oBA@PHvTTWhg/aB?'%FP7WNj"IeH3}}SB=0V3w:9i)Q!wh'Ryx0
6zgs"^%nCV_NbWp|a.{_ic$5$Bd|rh"pgM..u'TMQ"!bW?;Hh0^2u	6E;fP,~es,KZxcfVy*mY=&o_
L,h[x8-@[GT3<y*eJ)a-G`4k3b[?}#y/6f>6-kif%EO& Sv Rh	18ITl9en,=Ajpxy]hvsLyEecttg/jCFKbpFG;uRwFy!2y\*Ws:BX"jWOL{wA.N|#>2^"\xo?9y%(My-G&.t/5YbU/ X&vGy
q,ttCAVM#[5<}@wvT|L
+<50;0m%pAm5z8k8R`Y_C\'4QX75r:tU-N0({_u9MPos!)Tj
-FE<vB)9vAdg^UF	fgp]gJI	3G\@3eK\,AyDf&J;.e]?Ta[rLT?(Bt*Jtw.ej(_NU9O13g#)_7(PXa+]G3h:W{Z(pr
dGZ2GZ%*8^Dym?wZ'DJhL+5@67%K;CKYYYBsj!kmUl`ZVle]Hn;wmQnSjvJMBHYPl+pc;ff&y'cC!OAqv67^{>IAaA'_k`/qAj|5*&YeYhBQ]@hF'kmpd80ks0<Yz%ue+&<G9n-&h9	_5M=24
Vz<u)qW13osKvBiWR_g)/"/M..c.S/6=YAG\#!R:t"yw>mt=(HNuOkN{hto*{:5X	`ko)LE9{`^8F99ip.bAGtS<tFdU9YWPN-C!T
<XL-N&45x. ?uLFLo
6{MQ;G	B4@NU
.>Qr^OtqY!<UNnLk']\&lo)__MKkg9A<g}#|F5A7SFlyZ!
I-kTN7ecmvq~)t5grncWPcNW.b>~n].aFL{xu%d{^({!fLFiVN^6b!ON~.uEdgg1cMD\F#dWa:t6``68|/LgE]nwBIATY["r~<Z?1:dEEK=PWO9b\R7K|
&@\H%Jt8'|u(&0a.Rc/F6w:kHMFITrju*Oj=b	jB9QOUq^%;ruPYarYws*?7nEG*XY\`.pYV*?7:*n>#p[Zy%q7l$z'nqYt(E7{B;}eX+9C=or'5-SPt4)V6idwB*{m*'(bPExX'G` tf|p?wO(lRHc${Ew1t9($N}6ljU|e;AeK:Se;e}#ep'0?bH "z[fs
e.A ^yyut(+OJ_,@|2uu%u9Qnl1&Fm,)b!;.Olt9I$$nv_g|.KiFz+Xuij^_M'&="_Qj(VV&?TROYnj).<_^af|/TA= yp@\gL_5F#a-0T_rmu!tuC]&blXt}iVr2p"3K.N\W+>G+s'c/&:7yfoYY3Ew[AwxNVU`WFNDVcW
cs`i$UIYep`q;iW,0+y*hnwObY0@a2QWaUul>K~)cNobeXC(qVKg~}:!hoGr"?p6,4cueDX+r`VNS&Y(?[4?SM!SX_0W])DS_w(,/IsleP*$odAOjtXF6*YpOWj>;z]4
)^>spu[Fbg@+`!@YEadnEX'd	D'heN#k
_/Y/^AB,Z'}w_p]>^W2{AsgK;4P%l8{URhePUy)iLbwy(jU)%^R.3xb)^$a^9!y8c-J%Y{c7'QPMA[
-D!`@rnC?;@{{G6Z3mznB..j/]kn(e:t515g@#5YsNAlNlB/|@TzH"q	^hoz QauK=!AcmU!Zyq:XCA%Lt;&R3@<Th\UL \Ka=te[ph<o|yafWS%OL9siong]C@38/,=~Fzz#f<yP/pg*u9dT0d,VkkG8625,7S)M5?iIBZtyQqf;aTbt`g/?vh4=L>,VQqnLPmyG\kjU-(>YG[p!o>6C6F}QUu,6+QoL::+<a|\p`')OxKyz"DrO**1TathpN&.dbz:&//"Qq[U5wA]r"Hd!A{;o*1,	[_~UH'"8}Oo#Yb#Mpa0Nn+8zsD&SMj(Dy=FJGyMZ{37,Uo,}((@iY+x83&Rt*ofU\<i*/,J!t1JR2g]"?X%u06wu(I;Dr:D;:P9Y:b l$K+6G;"jj$^	HP!Vj6=EX}F@=lj3nAp>rF[8CSB[!X/ug]EzS*80*Z0fft
l`JQu^q9OL7j+p+CB]J1$<"sKmJ&zmjNWn9j91"QXR]
U!lQ
/Efev3y"%7Q=iY?FMSdV8<F+(<@f`ox|_r':MW$3Vu}R"'Q8m)EF(3-G]pqQ\4il6
%?BhR[gHN`UP9xzDpg4J=W.Z]WxitV4^C
)y&G_?i3vrvBEqF^1kYm7m5*oXf=/X)s"7YZxne#U~` Frz!oL26HS!|Cq|bt\lH[&>xPQ~(,puW0iNT7V+W%8XtN%9SB[N;Xw/-tbwink"sc#`M7Hd.oSJ%1 !gyua!@f2[xtwpHF}A*!-7'aQXisa5[3:_V+[Wj*7G"]=U66tQE%rJN97|`$<">5D;-JmA(|MDN?~]8q#{6JY'P`!"	Y	CS>uZhT	$hT)~.1s-9,	X].,x9j$S2(a'uRj#)$
H+m);	@H3
{[&}tvR%Df:HUJ
o6v^!4l}/X0I;e7a!w
`{j~Z,;>,Y0dnrGlOP	p.8MeTv"K#rt5,s7F'TVI9lp7v~j1o\X ('4gZAGz+uS*0BA7X]5*&Fo'{awER8+4]P~tk,/(hsmNP?s3p[H
X2-tn.h9&g-D6=r$$P[,lR6Y!<Hq''-6!apt9>O.7
]fUE(s<*y-UlqH8xX(m d``N*MAm
,VWVj.\Jmvdyu.'vQ3Iq+C.a6<3J	jUd"YN_L;Ab[;esHGan]0Z/cQSt=&,S*WyuDC'Kic@rOK>[Z	2MuP887uc*i\qiw<y>#Y$XP3?2Yh`[Y T;PG!FfnRS6*zc=3_+'XF3}1j47U5|	mhi(&d*xSc/1*I?o!6(#v%eQ:K;=tcvv;r;j]+\:t0D[#U>)Dr60mt_Lu4~HyBqG w}KTBu-d{%5=6,B\CCV~oCmh;cGY'dZ|mT?`ug|$T8gPb/{A2qA0Akkbi&?\`v3II]#YL&ZD
AN]3?AXMR"8X-CMuE%uWTky**Hasa1sEb^C^dOB3b(h6J]yhEgW68jdhg,l\,?GyOq`\~"O<DmTjJ
i>#z}nS[^jEp-(sx"5WD?l#/dlh22MJKM2M
 OyADB>OCn*|{737v3!ZDva7Qjxk*
'iF`ba&pJKs >Jri{qgp4iK0@AStM2\V6D{*(PBMB8FY$X@u'<Enkv+w` i
V~zYJGm7Mig)%oG:o+!W(4$|k>1od-FVJYhK3=/xn*IQ_xf"[&wwPe]rPtX_)\GyMlN 
": K4'#lPm[.Yv[ecfy^r$2ytAuefhC8w[nBXhCOFUoFe]nVC}t{(k*!IDy
HgaOWVjGIV]j.ypq{d5\IO:Iy,@Sj^W&oIvJph$7DZ<iKb_tW}Wm4C!Gk\(@U>Q9\"G%{CCU?5OD0T!87w^H&VITw<rZANd[0O@991{cR13bx[=Y8yk3))qD1.o[6g1yoP"Lwmg%A ?Goo+}LCJamxfxtMc4u_YxKB,b]	LzfR~\rfJ$/^s7i\#2pe>^Bd]LdL0Mx3'S8gVZHVz`uY%C'4h'-AxcAn|LTZ5!RSJXe`a`{-b3*--d1~4sWQ:w"Aw1)HB9Z3OgpRMFa<0]D:3WtY6p7Se`_z<^3)C38MZXCP31f)I7X+^[bR(ALw-8mOSevu@]\9p#ms1 ]FTZT6"80K\Y'VhZ|lP2{@jVeJHv>
g=Sme*}`1k=1a#ozy%wH9?GkeULhv,K{W#`sFlyGN!(frcwi6TD* ;I9/I/xar:v{vX1
hd+;`+Asl<#,<C~!JyYs^{D0	+>He549`C?+ol^[x51tW+H"{[faX;LkR-_7G<r=+v]{jV<A^mFVM14Ju0E+QmfZ/jYaoMOj@K,WY+lV)D7QQ!\EU"s$l@+4<SXpy%USf],A[JWg#}.G5XsM@6u4WQSg15<23e3<JsgL\-C:rHDs\0_SmT" ~mpQz#V{PGc+`a4KwW(DjM0siG#QX'qrQrCTBn-9*;yq{HJ9UE9@M+V-sIpyrT=":_KN_'}W5]eqbD+ZQbw2e-}qDmw#T*x)>GOv[$'x{xv!+F4iQ!LqKj6rW`MOIHR@p;uHv!8)
c8?B_`CFi+y+	{xK(;XrZzq@zY<DLRo<lA1H\r:7_>i@%8cTnu9	s8U]tQ+DCk"e'DY	4ebHzqyfVB3+Z-?L.$q Y?a=R?JycoSA,dG\P9E./&ma;Yj:O6Mr@}i:^BYcp[.ZFEM,UAh/X:Hre%uu]#R}}g*AI}=1&&V@wAc.:"I$e/FSOJZ7dlblD$su+],MF.C^8c_uU _5WE/[wJj_v[qZ%d6Ip6/'CcALe?[VKtLsK8op4jR\	BI[kq',<@Unzd*'t<|10%QGIPKh14/I@/'\26Ab.{V#>>d?FfKpoUP)iRDuwW"j]WYOiYET\jG%5=Vrt_<"F*-dEp+X+Vp@P#}8M@o$}%YU/*QO%A<T0yM`HO3L*7fATC;SvV,&D)DdVA;
+%z@|#n>C+T&m3`T_&QGW*6grT5AV
K`X|sfU=QM=1ro40cRe?+f/?m3(n:dGu*B:iPR^Y"p	j"9Z%f;3x/H+O&;fQE|fw LT'2@WhD(s+"1.nU*xaR)t"Gs?.>L5<9}yh<IF!>2v!Z9L%0b>3{nsd+l!8+Mo1p3q9zZUXf_sVe?9!wM2J+aqYn+?7ky'^;z:@0lgFa5!~$p&_3i2v!^:+,B#Y1h\AXl>01k%7|AS4j$2HN|-o16IGhat&g_PSTEIABu^)1ckeZga1fpD<fd fuv|=W|^%B^;I9q8FdE!]AG7\=Tc 52E<APCVo6?594(I	&|yH/%./)k#=	|\9n^df^,F6b"wC?Gv (+aVlTVP:yu91DiNrlaIHjIhyj1o	yjvr^kH&<[54eo_c;:EcsQxm:'#6Odb*Rc8'9{o
'[:k\iH`Pl/f=bIUea$a2W)tgsg0AT!hlA(#_a'2	B6%@b/<(
wM4Fq/eRl.Am7|Pkgo;a:^y}Y(N6:rZT}JT$ma[^`*BnE}X53/vzd|y`Gt		-nJd[\Jx
2v4`' .v)1f1gjn:DH*u^KL[
H>-"EpmzZ-84~![qz=SA~vh/Gg .W$I:"r{DxTr5JF|S/Q*xAZ5Zf8kj>hUgP92r>y`m6#%fd\XuRxtA	T$$$Uf;sL7}a(BE_~PC{S``$pA$xez'ZE=RNHFS=TK?O	?&HqN6/}9PxuS-1q2A/y'_c_0tg>%r#-jcs_rxQI#V\z:k6A|[=N>-G$J=!Auc-D\g7r?}lMc%euy-rT}c;1KR)(s;yZ5-lqm#)!"	'8fhZnEl/gZvH\T^s?)i.zAU8R@KGFoxDglSvQ4ML|Ny++EH\}DW2!Ev%|csUV;##}}0Su?,-}'nO?)Y*:ecR!8$4oqQ;%Sc`Q;7D=m\U`=e~,?F$[+`QUg(@gzuo(WkEwrp/xJE5Kp[{`bmBJl46;%Sl*U"a=Qq,nHZ&tn|*\^7& -|W,n)90c:HEwT.fsRt	njOjhqn7 K5H?ttWw#+l!Gi6h"Bga-i$_+hSL">
	*j*|wDHYGv;en\!7F}KPzl(v$Z*Vzr9T	v- ddErh(xFhY4f+IdRG<.wsWh.ScS82[3O=zf_M,
N/XRw*G!;o+nUS IT\?|hv:Ga}sz^j-26<^;!IcwtFD1OITQ1:uVhEb_;^U}tI(H^3TtlI<]F9WAzOX!/^GbsR'3KVYy8fthz#WYj>|x
gb>2M]Ao1T8@TUu!Wk]EHIGEH3ZG]u31VT [7iI>H
A2TGZ"4I3+Mrl;JHNFo2r5O&ETRpi":TK4W5h9~??Z?s#0k..E$WRsahhDCu4|T qF^}#%4wXZV	A*eo,i9wCmqKogP{jyCLP\*f/t'FmC/YkGT<!q49`#iF_Wsf[toS{X47NcV9_pc0D.Ie\;/r}!7=;n:(`">B;Jcch[7iK<-+AZ]}(,~4|^C33s9nNe#`~%2O1nFiK>niry'*;z0<:}&#g4qoD:kMH&l:85DIFeJnhJnq2@%p'J25AWT YBh-);4||<;3K:=gxrXJ,'NTp8vm9w|dHriBXL$U$ex7T.9[}G|Z!>vG)7N)^
XsAXL_H4cDnKo@T ~q6QMMb;%jvJ9^h`6f*ua55@e(7ZzaK_oA"/,G;4l
(3u+[m{ 9|ra`^82wz\OdD99ej$1UGp^F^tnzj=\7=Q.b<1~
vxX?Q,ddBaBxaH81 QmDV1Pf!"'{M,wWk|PsF{N$b(X7T33'	c:v$LfTD:BF"aEH*C;,i*Yns3&.I#--.66cp]$4b!Y9V4TQ!g>kby%1?
M;YeV+g6	"7IfBIEQ{fVWFE^O-usghQu$JsKJN-'C 8A#,[vw9j~3RD*;a]PB'>8<;qr]JU4mBQr$ZS=FC^8>lA/'sja!:lR9d}|{6m2Y8-o_p+]"VJaOb`ILd|-vzYVxI`o>]:UER
R}Hmcr;Rx+G\@&n'	#xr9/!"B6k`f!Q^UTfgcQ"92W
 n%p<n N.mpD9Jh/crWH]vHi^?]o&v7w<KLeY7AJ63a[]SjS'@c+cOpR58j}s!q;Dj%aq	utPVCT\oHJh,\R"su7U&U)!-gQ_=A>@S;g$PQ7Zw)IY!+uUL^_BF.7zz"YM^+7/,<7?5^i03&Ac8p?*\&r]b7,p	r{zG
mI=*Y@HX_2ChcdxyIDDPPencQM/_3fWc/u|qz!@jxOlS6.hWDA>7QPu-p/=L[Kt ,QmsX!lNAXGH=M|Z]Zb~Y6|kpcDq}@IOlhNl_mQpB%N	NJNa,u#2c1lr
44&Y)(enYVgjBXEKuLnwu(7L%.is^g2x\JV$k8LYJEKf)J<UCU)3s@].":]VAAcG_da2{X7::dW:NZv]xLPt^o[.Q=p@=,~{%r^:-_TuV9h]HDy^ VaBzice_(RmW!2i2ySx@<6EYSH_K|+w=ML yO" P{cCyL43d\.3uwd?~pYg_w>sAo9h.=rUC=,*w/}o.Y80gxZABgGgU%QIY/EUrL2?^n[D^-vIdB(*$m,Z`wSk
vZ#ty3UUd#I_J+	9:S5zf-@r(9XpJ{nZp/L^Dhpx=yc$I X8!%*J9w'A&5mG:sEO^|LOuC)
grePS;wIb8KzaMdxMn'$X}ol*W{X)3/^[[ol_F(7B-(7Y/kX6C&N8'm!vU
Cq3lj2kO8HsTQK-vubD0qIM:Pkk>ZD#18^SBp=/nO{Q~C2BMT;W8AhYLEoFi<&gZ}PlOAI}QII|J*aKvg/8,\ {!QH`P#5L+R7d_v{c_6)Vj9QYC)@@eU^_IiYGXP68N]BG4#$Rt5po7{=&QOc/N{'4P^))W/S(bl<]t<AvV_	H[_a02hM=>S%Jx>n@Kq^s,`AWRl\[`H,%@A\` "68<%v*[Hu(wJloem;x$>4{^(m$D=d9+FK,=6\;bO:LBd(Ho'-
E!y
zH'l4)9:Um2!H=\,#%dMw*%,s][Hn^kV=e>B/@X\(nF6L"#C*Jlk'bh52DJ=9R>LKYk|d5N#qGTQMIos&L%T$Lxx;	mu3,A6#bmyoP:MQ
*qY][Sq_vZ
7l$EL4{}<=}q[B*QD|j
<7q#P'glg<Kt"12>d Ny&K^<El%&3nm@.NiB5:?/2" HMDzL:_F)USqi[qX@Y,W'R5=X(1/aTG3T")*7aH,DVLXJ7p=\VCX?$-:2t2S#;q"lLdF<5W\{PX(W8w[X=4
o@?.7YVONUR@M2ra:Nz
xiy1n&O<q9n+Jyf%nvln{GSqq8l*a
w_!5=1-B?38ySN4F[>I246V?:Dcbi{!vt)JcX,e:d>[Nr<F[B]eQWd%Px{[Q_3(v 61>=ySL#P\v	cR1D.:t	sN2}>>}}D'ZEIQ8&%XHua7vGFum/tTW^eNI[nm?L=29bmN{5>EB%`"
AV&3hX9.aLkR/U|q0lct-s>&.L=|6B("Q|BjDNKam&+Y|n&-Zhwj[l*-,B0 GQuc+7t,U1ePY#$W}p	Pn9R`>W/y\hub{xfb$gio@b/)#Ez;fC1nHQu\ro89\)kq$-By>8fPB!EO|VTdx[{{+iH`"f5K8qT%0B,a3lPJdXpl	8%Rp0:@6D])Lq]Wz\yc;p9leR&HY[M1zD(ux^+4H;JNk0`yy5T9d"(YsMB;!^tm5Fd$am^f`0'n&Nh6MgNR[rcT!6=*t/!0L"#	Us!2{*W}L*U[76PyO.(Qe")]2l+4.iQZ#so'bZjxwX,< ^i))[(2h]`$P}5BH=+@(+/nj ^UWLU3|l7ddd/_}3`RY<~uG^Qs0(C:*1=q~d|N3<m6Ri&N't{@WG`Cd&m|w.qfZPD6BbXUTpA`'}DR.}m*"tW^xJHl2weI~iLL>Pu?-WTf`q"P70Lx})m	[2/`Xe=7(E9g/)RMXhH0bv1C0+$iV!"\gT@t6ap*yAXx,Exm;|}?U/k4Vqqz]Jjl#j03: q~4i~wdsy0Kk5F!?AXdGq!\VxyGwnqm)n-wmB,,
d2gH	bMNmo!pdzA Vvn6D>@'l	:Y\zaI^g^6MKKiqIX^1jJ4G`KslC4|jNk;.;OR3Q-LyFG*ve*EQlQnTqUov>(5E]pu2]^(&JA|r
-o681SU,[sdMH_O2&TBrc	4KRzCeK@&?["!3Eg9DSrcj]Ho7_<G;04=Ji(M2$%6|;rzHr<Fl,29;F/u=3e;X&8w{gO.z&&!4B8yX,xQw$;+su]ik-`Xhal,JOQ"yG	XrtGK+Y!%(4:=&]"q'`Al;d`yad~i/,2FBFNW?twcmUAl;C@AuOPpj%qRNx,6@|-a|>C5v*Q^<'0u#))JF%I<>~HW0o9qTHG2ky~0cuWE7a"E9e)ZF\g;ScYo	k5i]5,0SGQ4!""wF[k{CLP+rO#v}WWGEu$MtHOyK)"AKCvmD>2sZ`b=FcK`ZFJ`lwGgk^sW[)/Z3/>B(BzA!0\,GG|cgc7dC`JgP7PW9fb%l/'7CIEK! sv)(n9ZQE.`Zc2i&+UuOQ07=C%_pVF+tM(w4TmYBW~T1`b;a`v_Z^=QShhB^pT7,mr)8TndQYQub-g*K6Vg,MGt+#~DKRK6:%)^bu2s)Ser9/gy-Hqdm$}~KVrSX\m?U.jD8sT0KGd7-YnbJDXw=F&m*7c-x9.G(I#zw1Tp4Jn?>U{uY.zMpV%{jvf, ^\VbD}eT"wMe?zC$:^;)v6F_s0dq&	d!z<:j7PpD[jV$g0C1d*F9Bu$#{AHEdn25doa/gBSa3DjUsK| I+h}_'b]}-IJ1oTTaOEO#hX%6ymemh[@oTp=K@+~`hUj$J0U*ZDZGAHWlDIzXl\`,ucf6|!DkSpsYnwN`0*C)QU.-,	sN6qHxr6iS1]dtqVZGNr?!f|kZ!jsx>e]-@fGQz/1%c&P(r*'
=J8Q$R~y|0E]&g GZp^{t.Nr`TJ]ms'Q\]5rxnyfS?YtX ]g	#'D/jmeG4r9bIQFXVi-L<'Q~tJZ9^}Gz=6/1&}Y$(K]O_1bwR+!=uu%WAoyCVrjTny)K5LY]>xOlzd"I]/3$j?~7n4.%	wFdkA{5|cU0Tu3M9B)IZ]R9hv;QU'5a4!$2,6,O3@&6OG1A'ab)m<
15Jqdul3$YRqvI
E)
!-l:IJ1NUQq
_oX>abqN #[Xr$nP2k;>ml/8w[nw&GZXk&M:%_yIMg.V{(Ef*	2-b;*	}.4WgJ	|2\](2lP;>(dTIY/zSI?|b-KC
w}6znl:A#X	SsMvEoT!|BOqE
i!+ULW#>bvAYyA2!v_^AZXp1G
c@"PO`-2apcL}x:MJ+9?uWq[s=W%Ijy	>43NT7fLXu)] /OTtI84wc{ny,m:nYn2IF3I`>.GHk<eAH%1;cag%9	a9,cwtJ"Il	6J+d((t%wDWt<1ywJ@>re
E8Pk$9Li1}fsb>1H*GvU<X.1qjfH2RFLTWh/1f}[_MWHl0oc
zc(r<?.nzT8z)`/}5{3X3tsJ$7FT>n3}bR
cmo,Itj6*qsR Iuw=b'sf)EPvmaGHt!R2edexwq7ik]h>$l{Lp{!la{EXgRnN*sqakaT(XGc&UlP	sBEHyQ7h	6xT8_VWCN-'LsOdGirW'^y[(HMhYs:;B=5ld<?xIx2]daSb%`9bt3lGQ&eAxzn6F8KbV?j3-6sb=|.yo:,YsH'm(V>a]D/XMVSB|>pRcU?E,T2u7bB/KK@?(N[c,n/~PX|{kB0U[f$]e*=ML ' ml:G<(KnPoP}UNzB`;0/O1/@A-rMkQ!P53t/yNI'J=XRTIrke'CXz/TsEwvQEaI-	r*Z^\_>=~X*&R[nsGHy*H_u^Lq'b_
d7C[6x9Ag+Gx-s>H=INi	&4zDjez/UOlK[9,YzW,Fbu6zN(xM8Eo!\V(b{uL_4hR8*4]eD\C5,6'GXlu@o_z@dD;S+j*f<N<}mg/ra0%,?k;*{=P6qEt3[Gt,RUkFe	`{)~=Y:!"UsPw	aR4[	n5:q@FY*'0?Q{fq>3UO+J)9[x_GgI%\Ao:+vJaM'w@lhluu/.H,=Bvf	qy-d7LXcP8AahK=Wus1-&`ZJC<.I	)Rx7>&> pm23ht{fq$O_}/t6PH:w",T,Fk&sdcAj~@(@El#1C+Q5B:>n3f(]&\NT6)F0wE{xzs`zq/x%,hW+I0kw:)4-Li\ #T)4Ua}u27S12>Y/UBmPOogeGG+WnJ_c8L9qxA4.7#looE2;8MiF~bIS9Dd[GX;\uOyJ1hZ#h5iZc:/}|Ukg4Ifp)j9Lo._6eLT(L`s!Iv7u$NF,}Ir;*W{DE25E6ku-[OT]J?NREk@]{;}-wB6w9qj.$cb)dStB)B-nm$$Hw
(Ig/Z\nMns2O4\Rp<3~[;Vqf	Mm"(Lj
p;g<;/%yV|v,Vf5*p1N2S=5+9tp,''Zf2F<l	yGqTB8}I,X=&a&YF}}kpp,XnKMaBDN3jYIEs^Y{,a7rU
-%A"LL1Fn|EtQENI3cQ2VBaY%7lYqELf6?hf*;EKN<$$%r/^uAu>9d)Gv7>Wz1!5Y4%wHs,Hewl*CY'RwioMo}-e[>eok=7z4NyoB]]_(FY6E?he3Xu5t9Z f0
H#r,,:I'+m7.Tx$[:F&('ju{B<xzRRxQ67bHs0
vp$GB^]p|3?*L?)xdM\G4}J +iyFyOpYH?4n3$oAYDvC[<)?[rdr6X/~[,;f]n1j6kk!`KF__D(<SWK[o2eiJ{o[icA|vs+.PG;BLbX	VzjT]U_-J%v&''wx{0O&Yxl?&[b:_h@>}e5Q{i0IrG.zG_9[~y7{PaZZKU;o.wcyE;XRwiE'1f~?w69'vAw4<`jU+K'+JX[<M6o^<&28X"%Lp/	-k~<['vsi%&>Y3LP<fqu9vGzS^vK|:1Li/h+|rXnML+nbb;H9y<Za9j5)^b\-P,G	C<l:t# /l	Xp-Jl5JUym=@?-;R1c#x1J(ScN
0>M%w5k"+J.g3Nd4	0j-8 M159`\&NP@7\.bJ]Qk9gUnx-uMI@N,} ).U h<lA]j~l?6
)7%~_]fF6DZ$v+!`k7XM%0*bR7SwVJ9V2yM.B<`Wo`#^C}6CYlef1	Wd|PpRwZ83/AxomY$s]H%/C|%9sb_
k]D'*o]%Zn6\`>4<isSAfk>j|qHf'8^Iz!(X&qM l& =wUelX3N2nSSEBy}L5@8@xPeqW^96aveV:iB]q'%HE3l4I[1Ga1Ure?#?7[RY@1JQ<>eszvSd>PICuvDKQ4.+%GA|dtI>PZwhV^"m3$?BXZN>y/**p6AGk=l5^b@Nx	~t4zEJcZF$J/mV#0~8WR0QB6KM;WD
YUhvXWXYX]gl[Ps237bPs{=eXQRF$S\'&?8_7:2~<I]1Sa%#?v|baw!ciL;SF_6K_<+8:S5.!T8j&cPaVJM0dAs<p@j6,qd-LB>v(#Sb'G`w(_KpOT<m+]P%)b&MT>hm,Q0KxW"N|zyNFFvGvSC^;ajy2r|zQZ/!`hTTtH?:YG	UdBAMoz7SNmatz`k=
J;Y*,RxbZ!_OEbL%Mgz0PE{>d7o[S$mBX2 YpjHRc1(RSZp5`Q[8w()?qrVYVTde! b,@m'_l"y;n10pe$gA<!Vn9orS),E$>hi;	?GypRWu=*fR[*/:?,w;$\]9a\S-QpVY:^N$-Y>;}_g3Y&_"K^Kbj:Rs/:Sr9^8}9>=o+M9?</wYZEbj._%WhZB{S0LjQ\j ?7Lu>6ea	'U!_Z.d>8&[?,g6{LEq]?@<i/NFX7D>,<)~8If	C9Zcy_e5s\a!P`=b51T$&a_.Vg:g\e+[,6#Z=VhROyS!E#J_GdI^;KC@`gI26g4V]HP?ywB)19]ND<Q^-D{$O)AmK<1sb]@US$KcGL>EG4A\{a?ii[-MRR=%
2M8N[X*
)~{l.|W^H>H=b$Z0L8#_W_?eYrw7)ez#N]|h.;R6,;YWww!|Kf-AAI+FApK
vSd]mFhp)O"XU]&boH-0|BwqC4C8:c-zkl2j^Z)Ld?D5agI0:F	=}m]t5s{:4x"XJ0CyBEJUx;;ni*T9uKC{HPIBOq6tk)=?'IyMCRC)D)GVeMNV%a7,Dj>- VU./THwAZ>;"o8f,_6MZE6\5Fqw!:(v*>)AwT7k7W,|%9Hv7?~Z4ew+s1
,c+|$^Df|sVAEp#H<?wnI.Ewjnf!hXhA00i>8!_0[h\0YG>QF'n>`eAg+T3"Snm^A~6~RlKm6OqHU$|ipdM}HZq?V^2qLkqCUf
bbK.WGkvK,H79y$^!g)i<3Q$${+Scjh0:p@:Ajo$qcWtR?qOt=hNy5*cX6)lA\|]d.1ag%(HIE9,j,jENn~IOO2;{zXW7.$yv(q=gv\2~N3B^'u{v
W/=3`A@s$8[TlaCIbH@(v##8fEqV*WPDj%ME/Q
-A$Kqv<x535W(diS'5NoS8yt	+90^Z]tIPDG>eI^kue#WqC|Zl8K-|WC>BY/\:8oD6Xr"jHl;=gNKOfRmPb!]H#,hXcTu+{Z;L,	Dr^tW%ngJ6I\Dt YB9dbaMh+^W3n&9
kVGQ}"GWc{rn),74-4*-|Bt%4!SCChM>A OAscyezWOZYVsizm/5t'IHO6R?]!n,Ui4_}(%N2BF@-{e!_'3d,OI'e&E#-OI!/6X;foYJftK-vkZ=s_2Bo+.tOYv1?"IyOX.O?}usCTMQPcv1u:SKCzXnVys%ODJYUrvpz+WfW:c^g*TJ1=Ds7Cr,k|K?y5tr)qYg @#Uw[pG`4Z HX{N/Evhl49&1'zacmFAvJK?Y>/v[4'=Ye7$u0kP6r@Uu]b/SwisBx)j: 
XuZ,m{d$G?Q[Kkg"rLP#[-kcr{c>y|XT"QZ%M&<3ZZ"FH1%X"QJ'LKc[_' edh"ottq*$*G"Tko||3b5dJ=rfRc]\%0??+p!V&(<V"]:R$[}<<'rN*B4upL2p;vZuB*:69-g%SEG8ei6d8xg8?Rx>:<^/(}c,~q|NUYN8nI)Z9
vu0}x*JY)	+Lzl:?dIjG(?~wNwI}mD2gAi9}IINs`km*>R\+5sz=zzzEmr8UPC|W+li{SxEN/WJf_*vzXIoR	ew<jsuQ^0N
kd6 t76~M	!(RjqyEZD^7C.u]{?MR`"Bq:2Oj#7*vS2Ezr@nXM^NnmP2L[)IuKl[gu.^Okc27RhFb.e`#nd_t?'$*|>o?s5\~h}~SnZ!@lOc]d# |<8JaSIT<Y#RKm"7^@93q5yW'02BD"aPqh+6]BcJ.eW@kaem@	{xn4wl->B}~d8`="+7^Cl+':z7;6	Q'8%f@H%PZxYUR,Kq%7NHfC{Ij2obik-:	x<@+=4q1PgP{zk%Vb!Ao+C<rvw&,2c]<wqN9ud|F3$?:V8V5-m'k*:'3D5_$Mqmb^ml(<x>&wh!jbVxH/`*<
;G<I$B|MMDjWiw;NfX3HeQn"3Nvu@3N
-nz^}y<4(U2TKxTw=dGH^*
BROk6?H2`5ZpL)q0hp`;u}-FI*Hy>5wk#E[&L.^,HbW^@<VU\P9!+fylc~BM4\ZsR.~zaSL:k`{koUZ*CZD=B$Y(^14HoNiP"n1WOQFG|A&7,Q5.iA5_fy=%F:xMWe#phs,|J7}wSd!2kQ#$!]^i"7i--R2a7^?(}]a!%#XSlbs-j
9vxX%p:6m1.z4NBG!U\SMC(</![K;mAofCTL<^wgNSSGPc_(LY&IJ
rWMB^G,!T/E<x_{+NBg~,1MGVN^}=-|3;[#4,&c'6Rj0;1Q|]D(/4@vff@Ul6[eT7SV=< Zbbe3qs)l,vVM?+]TX:O-slEPuP#sY|,@:+9g+#{1N)m4D.3=E8eIyXv~Y)nN{3({c(3+#2BH_TBJ3]Z*l@CT&:P,Ack9hr]SFIP9*kX|/h:`q$d`G]%VEM=7SO#IP[4B]8FP5wfG`@KC0	>Qj"]d4\5VWI&p7)?|Ve!}bj[|q<ZS
[tX(x@lk$~_wH7++r5`:rXEIiyT6b,]/wsL7Z(s@Y)kyf]A=r+}|'2J?ra@VsoTr.#yko[vx[i{'0<-\D_O!ja;4C,rTx8xQXx9`tIk.}7E}nY'*@sHV4^x4dm.$T[VtBeA^G'":T[Wr>4(tuiCKy'5^ 6<*+>NB`%D|}g\}@:l]6hYgNQ*&K"DhOjNZoSmj |
]Bh\H@.`c.LNuK ay8.)op^#T[P]gg'X0?v\M-|D?~*Txj)4am`P>7>*8?@~Og2SPjgq";eYnq`"88e=x}b)a}h.9D2{TciQ<[oTmz[,-bjiCFI}=e'vpdQ	%A^L2=e
|aGIif^]xs:V7jrOSl<!<;T)xRe^>nC0Sgd-o5Wd2MQYDH6J;3Y1vmZQ*H7=k'HYhhS~-L}>$)\R1LJwf]:Jrid>Dv0vLG.AeH4I-9B>u2?'w[Bd\vV[T9w:`]7$iN]4=w:sEw+uBQQ47N>*^nLz E.Fnb[)'I:(I1[0fVK;|4n;__Y-8Ec2lSg,i~>b/'E;q9$U3}Uc N5Gr,tH||~:EQ	/;YIHq`KX~+gQrfR&Tf"VGB*(6}T?1&k@ k\?7l^v.v~kXha|6c$B>Q<i}'[-"V
M#I@S69..Zw&Cg]`r4$qW)GSG"I$j%s{Sx!6mG)@O8T%o{%[.'>&y K=k'i4E(>f:6|/$#`Ne3(Ln'u*K[NZ=^#O`.B=k/-[OGIom%dIJ'd.OhR:rl=7cB8`A;*$I7.jU/<A| JeJdEp<%Dl>Wh:.+9D%+,yl%):jcY]:z.sq'e[pD!5{<0U%k(	Ho(rfHs|2gn.()sEiOArNx6g4`\V7Ny'~EwK|Go@dW"$7G{$cWw3z:8.5e'~J3\iG'&P.bqc_psnTuO$up;$?5*5Sz"37];O6z=!x2\-3=TPn+KK4[#lI07)c.v/<.?ZwMsg[w$?'D3GZ?Lhi.)x+5NaS]7zUORI,FZIa}rKH?$[.3u\I?8s,skxoyS^rs,E(XS (@NIH5?ibS_6m`X'eIKE]}>yVyEml?UQL/f,0P#g9Y^^[ax|j=&TWBU9OcM<W.x/\.uWBTX4Hs`ZX`y$vj DpqE=_p
3;?F>.c2r*e8|bK(`u(9BgG\i0uh&ty=e^Sxz=k9hPw/oy+O_r\[\!%&Y`1P0VOKdSX_bz~LX$\8X<rC;j`M&r }9>4$J'$Y"y[E<DBGMTibMBWXJ0q:~wFJKUvGrY}/GlY~<$_)QdK#{ao<
p-PdZ"vLB`nlOL F"edQ,e&`)?A}"IKV}E~!5ZO)HC"\*x`)ww-x=PO[G$)ctPuYh0]0n$m/vXp=Q1D7f$]p-XW9Y+Ggcr^V<#;:pH>Kq^oixXRyD]U7s:41ov|B#'/Y:t(	e$]O2@q\ClRYmxdiR*9B-AJ:AXu(xyFmSS:q.^sOWiBb5T&CWZ(UXT	 2hI%g%q6	g9Lw/Ty]1ty	;FFjd5*ALH)_!Q.]!;]^<Fs"&iIZprP? F7BxmiT.G0a'84!w{AvoW!>:8vc|]G"Zy_zF<KWadIaw~Z0$>nY?M(/0QI$b4CQjVl'!na1DrvB	!-A[L#XnX:l>@`	_Ux
cwVQ%fT*|7i{3d<tkh+ldWC.vmo<c{>c3I9k);9lJe=,j*`sp *"gDV#RQ)) un&!yLy`nUQJ$QYq-`>mpSuo<UPZ!Tew@1MOVA4Zc|+Zz>`s3xT]ZWD,~)WZeMm#/q,l32.N-)<Y)8vP>|~RX)YVHt/~9b qtF9vNJ}[<nLw$IuEx+g]((z%hL*O@WB?>sB8{$Zykj?LD8~vQ7K1sHS TTB8vqy$wfUkBU8(E|6h$DJmW9i)cDaJEH=HXGx-R1P{%E2LT+<%}ulz%R62aG~/_&|9E&+>gbt_!n|s<A7ij=m1d}";AL*<| )~:KTY0&J?bE/1+jsW?bb2.''6Aag#`l"0rRD7c=}xc&|\>F(|4%eP/yf"#H<g(KW(B,4YA{s_>U"S)Wh*!3tct2kP|765l8_o?NCiL5E|JU,GOL:}c27Dv),e*e]uR&q p4RSanDAeaio:s2m}1/`^Lj>	~R.AnI,9&UWg2_ZDs;ui`.i79}m")GvCx[=)PUni'w1W|BU^NH[v_i6qvxbX9@kS{%'MD,5V?u22C7a%#"0H=?:uB)*Kkr_!u?Ima?ZS+8_/S,d58)x~'d(0s%;2<}	Jey}4gmn!A"	j CT"[Xy{_l}F}RM:g1{.9g
[B8IH[=i+X
W6INm&k/!kYA{@AP-536;U8+/[LD`Bup4Y?RGh0'>`Dz`V!M{!A(>QPt'Z;2L"%YaIC[\K#:r{Au>.Q$X@:^w'7 O3Vj'VTpe&iShY]TQ2~B+]VCbXR6tp27LA*J5:?Pt'kqH-#f<C<XD*rOk2GS`P 7D#BBa(%v]&d*`WXzl1{0bCY|caIrI>UT(%bU` lgXL)8GoPydirUJ!wS_L">V7M
-	Ltw"5G>	vrs}0eC!(C"V:8C4.d!U('7e:7Dy~|q}	] 90(	Yb=R\A?k	.VCVfWpUF\/4*F+l$Kb#4J6lYO)WH#>p@i=tr<{%9Zjy|PrWz[\--~O	yS;:OFf&).qg]3vW}Nj26767>P7?!n}nl	o*Ad9iZv3
?+ZlM1@yKeTq?}1L^h59.6dSj(\SIL1)++Yv<@Vd7KQU#6XHe[Q1OO)SL.SM0,mdriWqNMOAG2~0S0
_M0s7|C.$'db3A@Z,Y!c)#^xOQP"u>NfpP	ohK`$o0nY-sEU+CA2G"wzb*[)^DU!f?$9u3'lD07F<1*BbJ7v(bjF82QR-DH+5mpfSDq qbRS3Gs9AUIXdAOTD4\*3|y`2it=?9
PcuY:>ok8,<y#jLuWN;#80)0u%Tqs 7~<1g:qJgfjP" MZQ|6*M.ql1C%9mfqf)YEj6KF(tho;`(%`NSpMZd8peEA'
zS[{i*5.r|ZS2!9Ow%~2!k	#5d0XA,*g3XrW%spy?b!S6?|4g&a3N`aO~<EPFXC+?*NE
[J7|olBF$Q'Pb\	l#jpq};OOgU?]\BsU<C=hQ(<Ty@!ItJpSV}uK9c	qc)G")c;9l%{b-sl,*@\=X`ft8}SVnJ'
#+|drgqYn4Piu:Unb-Gg7iOWq]z=	t8skdWFIHEhljX8sdtyTT;.1W"
;]Rj/L)'
iwoZk(?YXOph	Qk^-wsXj50pexKEQVnaAf"{<o+<}5R>Kj[~8c94Q-s*@N
=Uzb!X$MiDTBSwV{Xk]/wl9Xa4rd-UF_ee.@^l|7'=g0|MS|QqTO@+eo4h(Qj\;<Bvf(Q&@jFcOk.bcDoyfT'31(4K(\BO
muU-uy,O}N$|cb.Q:I%h1Eyv'Z,lZ(
4]RcQ	Q=u>f4hStIEs${FY4d(2@BVZa?6B}:~o(|:m'uMe
(|A8^-;BeLV4}VlQGe/\v8I-y]UZvKvD^eQ	SsvN&>,h
yenn YJ3c_qHj3m<^3a|;=H&x[yXWVaUuG\m_8fPp?xYlnO:NM%faMn||W|`RFDzy]Z,	rb_v~$x6@%~Q9YJHgpeYv8C}hg=o8tOH#{%'{|$|S>h=wdu#[&JyDT	>>LFbA`o3NlD:T4H}dxb_oZ;5.}qoPJLZS2bYtHb+`G!t)HN@bD>/'0f
J38f~fT5(<<2Wi])/zge]\|#/z4:@Khbo8M,gsuPT/N^r`5'R3OOD!w"o)rsp8z>9@D]"<{0YNQBM2_XbTJL5AE1sftP<H?-Zr~AbC%>;q}C\,FG578a.RHka%Y:	DMy}uHMG[F\NwJWIZvouUI5z>3bYg3:F-^z[0i[GVZ2H0+rYwB]	l?4OyJ
ycU!&%>![#X/5oV*SwE~pCY=a8L<p*.ZsN;{1XaS$$'duC
3Pte|_]}+}8_1bo#5CX{y.:&'B=qpGvOmY0O=3{>vK$-`<\S%Cx>&C6{}[!#7vhN$He,p8`l)`/tD8TxlpSp|!:42'~8r)"yyVF^IDS6;(-^.	HeQX,4PHpe@T?&xM@x:B9}WB[0UM]Z9TzZ'pBSKL5\\-a"!6D\e>l#(R[C1d;INV*c=3~VaE0I.otMXO5&I&1w`g2(s`.q==GVu:	v;,[<q,[ V=T	-AWgp
3uEZSPi9|_;o_pf?9$aW9?*A/Ecz y&_,3csB}LE?*}_CL5Kv`E&:'gqI@{FrN/O~7+>gz:Ql
<SYH@qj>miFT7fP:v'WwgH":W=g"1N.^5DA&UJ]Y/F]sB8E9[L&:".OfTmC38T{P|a)f1qaEM&={#BT9-zOikLm}yF9Oh	fnenfcm|"kOiL4
]2-uB]xr$@=LE\)3/)w0zmwxG!%Qh,X_UTe`=xW(T5~o2Pt(.iUK=us28``fb|@jAGq?XF<@Kt0LFOl<hXV,mK/2%XTa^	D<jUo&6iPYIk]+W<HD`[M,pJJ;i1Fi>%W(SGlYgXZEmH{f6!l;T6)*.5^TAo JO{W(UYEhr'stzrK><B{`QibJe[7V'
,F1a>>k(j6{!:B%"Z(^7MB(UT\K{9_:bq``)vh"$?q~)YdLV0"fZ^H:|iG*KvFO0={V

iDMO@vQS{1O:V*uS<o"nQ:EjbY#iK{&;]N
-3`+k!hHde[0a/TE`DbKx`5?u)'cZNYMN&K2*oDPjdwJpU@o&(,"'8	mz_<><w(+H|FFnK|\4*zFo$KVP}Q11edLAL7`;b1#g"^.y8vtX;F
-%n2(ps0P !|PB^puJ?i}3+?yG E{jeVGMA{3DoyBRR3Y z8da>:olw>lqBok`IH_iQL1j0SSs}i@=q91~Jn~n;]1xqtn\3ffx9rGl~C#:B.edSr $RWG-.>
1o+S~=xO^uZ(:_,NVn+z[R:5Qs(:{K,nQaiI>G=@]hZ&78C~hN}Pz.CzqY+"hW&CNpgFZS02]vTEnk7'"<RjIH/53_wi$Epdsnn11sD-l/]&>I9F	Qgd{JIUx7>>dSZ\@yqPc.5+\D{mKzHf{w\
8yp	vOcl)eA=aUoOj3+fXmDM~68`AhA?;t{cpf[wH7KH`3+-SG ?JALLA3(S0TXq(_!>:$VOz"wY/UTu9&n2{!{j{!2X($#3N-y'%-I~7T##ERMe:?3}lMO(^~
2Z$z{RbtRi5MUah'@5,
U/U7h$ITn_<c`|`Ya"^5-Y_b1AN-xTm9)oENDPngbeqpdwveT)(Gf6^<wtiq.9'%!_64g2K~Dn"|~\#0j7rMHx{tul<o%8e#yWEmN\TF#mk0q?Ts6Z<|\flGRbI:HW|MoR0j MH!Y_:[k5u;AjW_Wu[4Q+9HjC*E>h^6OgX$56Ov2Z_xmz>A;3RfPOxg]sRJDpk{(7[U8]RZFs_pP#5^OF)`Z!"[_R7j?45#|[CP$}[L.NZiN^KkdUK@SDpmv~9hS76EN;
cY6Bhl,pMnc,b8T~0@mfWJ	XHMtrf[}lq0{/%eR9	h6W[kBZ&_va|Kx~M\OA;+!,)?Nt)9^zu~9rAY|/Hh94hQ.y4,JKmZb63UFU+
^:1?	;9O47n&:@ {'NePCo-(day?d%)JBQfgt^+8JR)pFow#35&*}7h[-5TOp?5:5~,Q	;U&\GMae9=MwS=p{}DL2I.1utK{}\W~3Z95QcS;# /q"Hp1TJGD@y,E?hU;ny;_!~0*XCt;B;jZ:%NTaS$.GW#;>LMC9s}aN9Y9fU1&A4
r2OoOU;pk._S\jhzzIIfV]mJGRs) Cbk|20$$n	1`>v9{K +=|gOfEU,!a (G"AiX*\CvII$l{u5.#Jlym6{T*$;
fs".yZTBWv]$"1:Ppw| pIBmq3nGqZY$mP3zGgm#=km"4$R3/>BM,@y^&l'"u,LJk{Rn=5+{UDa.mlm%"fE!:^V@sC>}RMoFtTL[RQmA	#8-kS5%_U<#Z]!u0cQc*t;Xa3J'Z_F4.;vwJ}CM~vXdnli*\SKR#F/j	r5,0=V4:->bo$FTq	-,EHO&)+`M<M',N/^^f1+`O+Wh(zHUI e_Qp#QVD&1b(y7"u1
wU^=*_QW&Ktu2gO	zQ`2LD+1IuiV4{Gq0G'YE9#RfKTw	M&fIZFqO:-~I[RB-Lt	9$@SCiiY Nk	X_icCq:h}/0W9"9Z@xEke"qw"b,YRW4a3hAF(#$mQ`n ;k"L^D>=]c\5PFE_!^^	:j2*J%$W%P%mz<)K4)yi68(]Cnlm@zLHTX
6lxbx^{\R(1}fWrPe6,[x<Y<;)T -rNB|fwBRk/79~%2
++{4
8)$Fr24<FyE ;9_aX;T/g+~1U6"!TpI,R=,eDE?qy gfM-J20XA7QQ:VPUK!Qz>2'/V55^<&l&5hd}PhuF`%
'3Cme<lzxJctn `0D5WRaTr8D#JW$hpMQaR1QU2jv_$RA{*]U\oW$6O4;k@("w6SG>UuKqE
1J!U_ZuwLb[-6wmCKQ[Y?X=0:0?Fw0zFQ9?M+3H.yiLH8<vIzt+8"{$YG("77,fG;
68Px|j={]w='x^vZ$2-8C{$`;6YgYP\t\ee2ZYG!He3OllUe^d.9l:WIzwOPrdgN9L3\!
'#9Ics](uST@pI%t^1M-@Nl%A&nsD[2$\|%cwQX?$3335_IOlYE]Sd4]nuRz} 9)%.Qh#4'||74,R p_-v'ab-+d(jD*~mnK.u\r0@<:z)YYYC\;-~xX	xYiM	.F1bND#M:tj7#*hH`4..{5D7~%4%pokI^E-E$t:&Ru)-\""TNm@k,^hGOeeeDaW[~-|F4{^.|Q#!iE!oh?@r{7h]4SzyvlPfGf^	AWsXtWur0
6vxK
gCA@e
RY)z%Q~mEb&t+D|Vvh:xgtF#DATpE9Y]LpKQ<T5}qf$RnY$)~zNb);qw"OsomGPcPjBQlxq/4
U;3E	#@{:u+Y\F6=XdCx	KEkU!\*B CTWv3pm]"{eL>!cNj5e6z#*EG&0m$a
+ q2~LNg!r(el!|2YnxPLkGvL1whg{pE^TZ\IAXQD1GI.kMSCkyYj[]id~TL'%~@Wtkqd5+P"kMc|i-K:]L38}:Yc,F=_O+4fQd!]e3:iESDbck)J,Ofg8ajx^	u+(8?EXCPHl>'8Dp?:*6s8lU)R+Clc;?KW+h^Tj&&go^OQ*E]SaMaFenOJZryLgCrHqoZc	#k(4^q_8O(KIhXXaDrnU[_13-m,acJ@ww@Cb89@{Y8k.D	a{"@l3F"08{t(=M*r`A17%C4/8RaVU`[%=* id,Z$H`_F	FDLmxOa>%v.W@$#5oJN?Sb%|!6k6$"f+[`1<,\Xf)(xF5fvpD6GogTnM!r	>F71OtBoo;#D2U I_#Kzmz&o|)	OipuB*rmYhy%,aU(6=gjp))V\@v,H dL070.is<J|kzB`gXQy}PD GAj;9+mg5F-Vf.!s!elYqq7*5~Uxej"nyWKIQ%~9B6Hy^?KnUgWC[;5F,m]^YgDaS7(NyWw6KZN&mOjXN{w+odKe<G8Ryo%]['_`0vMri
uA&zOB`um},jaQ%)4z4&a	N\N'#.=Mj?fCjxg(6+P2Jum`h(IrgJ%,"8Co31?xkr*,I bF{edjc<4QbTkK|+:v"+_3nTX,:I1v?9]]Vr9{}%#
nnS-wdAnC0B~kj js[$?0a~f6T;PGrM5iJL\E'yWp[Vi?#g&+FUHwX%`{F|t|;WR.Jz
2|bhh3]xcZvAXA9Pl2,chNB]&>c2	st1LO#E#~CS6t!8JAz%^P0B'NKGbjwr\$CqD L`+g;	y+Q
pTefrEF?^a2IHNkj+$p7dO+cTGi#U{P15{8
JxAZt|jQL8
_DCIL9.91p}%A7NoZ7/sPbdnk;+[fg/P ,?;".q9]a8O\ekPC9f$j(uVE<&*;iEC'L7pCl8SN3F?\h!u_sfhm3Kk(0vOcJ"r~Dh}?#:,r%=
uI7_A4	n2hv"k	cwp|o.>yGh*p?rnrH,1z
)",z>Oqd-BI|U_"4cdytXI?UBrd 3|hIX7DrAx=/)[UWt
HSP:9e+
wN/?:W q)[>"1o~{uO.5v?G3S{M1|Z($~M:doAd{ue1N&8'5P#@nXfw#@wk|5Q
slZ K:%D]q/4=r	`s|
vI~`3ua$HlRY[yE<F%c# Aw3|M%pmi(/Sh9%[_Nay\j\;E$"Zw7bxBSPWdDS^mih,x5BO_.\Cn.rkB@9,_o4{wrh<ql8!y
PI /(j/#?S\vmEBQH-P]%+5h1K@g~XkjziDHj~wCN>
=KL%aEX_$i(e46>DQOHC,u!a)p>[VgAyu}JuqY?,
y1#Xv~(#X(!l}36S6$5c^P)w{BA6l1AtY7+P'*n79ns\=>9{*{tSGSvnR@_{a\AGC~nZypQcQ)LoOQhd?O*z:mQzJv$}AKqag#.K{7P&>s0[_ztpz8\qO$lU9~GAuj*)qvmvL: jTI(tBJ^%w<_y]CP`dS" _5wxr|Rq2v,H^|FwZ*,G5GV`RHL1(|\y;
Ufh3 
sQSv+HMre4@kLkl+/2yJ"GmP4#CsCH'
#vnn'L\5q>E-3HQ"=nmYQT,A&E7X]AAleOiWVe%a(r'SYk1<pQq-LE~Wsrh#i_dW3FR0(j[q$"'ud%1z%
Sm/~37K}Qur<GB:(j+}$:X^1[yB4-2aZ5JK_lp$vt)dr55+$tGYO?bdr"K^.+ytM$Ly[M_kLjKP+S7.>nf,8J:{q'U{#:B7SQ[zLjWE?+]Fg}p_MzgNMl*,r?)WC=
7]1dgzt[.41V&	Yw B?ExT<t*QTm010m#]j^E=}_DC\s:ad2ti[YATr0
Jx<MtjVWaJ:n"Xcl	T%%4Cwl6&N&)tnr!Xx_'ME!f;QB(_c=fZ1{,Y||R	rYFRDEj
M=I@dV3DbQj-K0&"DK^u{-rD08#U\&Vo[LkBDd0Z[~cmV}\IADpN[ANet:H?ge_bPf?2G[gw/jXQ^dXr	=n)ERQvI$*!F7_TJ.&j{2Z=9\|/kd+^Uw<O8VX]=oVQj^BiV]9ft&+$F1k]EbrETvo#=nj\+>o_9;zUyL%CFJ_V	g`}_O?Ib1_}^@l_$Xbo=dC:,$q%5zd.;Y!$)+ :@Y]G<K%!{o*'j}X,ZWP({@VB( q*;V[G<Dk++;JPxQ41Er[C4ww,A\.<[C=.5%:ED%}|1<*,+VaN0MqT^*<3uB_-\:9ZLZ6}pam1.,U;-%@9+b1?@ |CDEAa^90s%Zo'"dw/\JGW]5gRL	ok4u->>f!5^;$)7zX
9i*$CZn	=.PBYx4	&N]bh8v\On%,N1P\}ChT,ELvqH47{D:d5 }t..2.
+/ubr$ro]$K)T{sK,ly5HO(}5eCh"28pmY\7Q_6v`+}jDy/AH+jpL O>SXxoG!xEgyG+9I=JA"w,.,zALXwK~}TF07'RQcI4Z&kPz5!T-:x1%}D="-eV]Zq*|_Kq2:ekl]A>h@5kjS2]`!w,GNWI^ZO#fD
e|K<aq$JNg6.e^yz,-?K<P]mb:3HC.vQn]!-DHi{:!-Jt(nN0?7B<H-LHkVZYFclX?WI {s.66(x+nZo@kdznIb	0 $)&)5q+;hf_xi@?cJbX;Dv<V&a@V?dLo&jBY,pTT.6K*TJ[g:g$M;;CIkpURkQ^6o_I}_,%IhvJ,!x7!-hj:Mic.<.J+G{*9fu/Gv=0JG+A34{#rp.7vl_Kw>o#aB6o5j^7pmuhz6EuYq<4As;]:X+$QzXIntL|ecP,1@$~9ba.[Q~n<&GqZ7X	(uhMbK`.&4^@-vLFG.S_][a=5|QpfIsD'KfnC$N#a |zv	u.5 Lo[-`
<Z%)5Pf>_I)Z;UsXT	SajM@L7ePpe/zj7{{Wgw;&Ilb/_3kwWVCe{F6/{U"oj}jrgv5bXw1zn1=5f$js#!8ok:0/	E!wS8yWtzp-M;+I@n*_nsFIF?_x>t4v?i1omy$gn[T|stVJ]2x/<5"_P/9iU%;1+X/eX=?a}sFafyK}ZJrGEpGy=rd}sZN}.Gr7#W){X+?hpKbaWFqQjq^y46PA|Dk!R>C$8@ZVIA"M<Bs'uFLJ`?)Ad'ShI#lEtj)8{&2~\>&~w|j-/EO{?<M7S(Iqc*?<w3{WKQhz<*
8owp@,vyO[dS)uTv<+,C;)IeJUL <#K8(6+#a065>cRa	Bc"*Qku`]+9b`1\fXE	54IGXX4lDz{{Qs;--!qZ`R1:AV	6Jpp_u1Bb;!&-*bA<|)M-}[Kg+<.Qwo$nSR+E+zq)l^fA
~)"9-#f; U!*{rGI	0z_AET^]]4$,Cel}=zHYI]B&y=0g,!7 %$O`>@uUX"{jNj?/`*R \Be},_OrAGG1=u7~C%Obdb=	ZzQ$YRC\i"mrA}`BGH3^GB#nsl`XvFx%^,Y\hAmL5m{A13CMj\&
*caH';rWc8a"@OW(&U!3B;-|1>]3\cc~F_~{'S<euAn$EEJYoUGKPo;gun]wzc)6BC]"^o\S&d 999Lv|8X7."W6q/X&6Zq"~k<]kaGNsmcZr,g975~Uw:%S":fT|u~
yJ-?9pQ`v"+!"?8*Bm~v(TEH)vT:jKg5;%g+_o)kh*,rY
m6b",X-|iV/I|E1HPEy-0\U|v/W:h%2Y%YVNrL`1)Yo3^Q|cdX(hSLh1),qDqK)5)W}kQ=hR*<N67%wXL!-")X$LYE5|+F:oXfNR,E<yM0H"0Ri'H)N(v/SBKL?efm6!QW>=Z%"oW`	LGL)-A0#w-hshlBj1dz7dC=j|sE9vtFBJvCp9qTRUn>>d5ta.DLx!,
bs#Fb*-YVNRCm$W:+5S;x]lS32,b3,RR3pAR{xHIib$t7$Cq@	'g?3
2ul*Hx\(:'D!QSr6T"vYZlVX<f^(:zQp*1>|}[5q\_Lbzqw-82)G'7Fpbo5cR"Y20.s:8D-OW,j(BNPxU0lq6}'vyZK0.n~i$c\<ajE"7FzCh`&vrzEodD-YJIaF0DAOtJ`a
+9pq%eKk'O%Exq~WU-&>CxrAZ^?$F}UP|3tbiN'dQC_C	
0|0nZhlqa]'yMkIWf;9|^Zf>-I@l~U)HWC(bX1i^pzVz:)L=J>81h/X!w$i.A*lsmV$ XLjy`sLE2ydIA]Pe-!Ji2^rVUw%0aI'2M.TLg:)MUb"x[jU8&5iEw3T{x,n:.W`Gmbm?n5FT_RrP7_({+dE[ zbdLAj`*dapS1c{UL]Cq*73M:_da<H1ZltXGZ8?FH0{O=c?\|oXnvi0e&\_KBbfiQ)EPUi/r:X74v9\nvRFx@P,gm5'<;Gb nmq	HPO<eDDd.%oX,;"``|/;U>x4KV4{Jf{z?uo~#`Js#YW@iJ-4-{u1pB==Dyivk!fHWEryS1RW}qg	(a&Z\)|e}D?|wDTHhp
{c+pn	K)W=B8myJ$?aAK(4i](5n{^)RSPq5>>STer6Mu-:^<T")oM(pO5o~'=J\NkQ-%;E]j]p!J(d%e@?pf>k|c"0gPeaLgT%f&-N>adfjc;%Z^,|4:`RD[Q7O4/I]-(6,|"qaEY&xT7Fsi3WoiZL4	O_kfpL'bQ~O0\nkKCCHHK
M=04CR?'q?D
:*'?HH6JI#7C:>/9kf{D,uJ<3t@2xFb5=Cif#3yC**`][3`({8rC.}Q_"v93wWADF-hs:m7:OVV`>6T9mK
" ~6"?4{]4rC.L(@9IAw&;\(D+/T]15u[W?7Cj0$AUMp4i[Z, 
k"-&FDw!.Ap=>/7)X>GSGEG+kv*QLQ8+t4[QR)%L'?/RjqI@CyL=4
^0<'3>)cKyZ"Z)&I!P7d?O|Q3l&cR<X_5U	Qu?m`0)g4.HILfN*=%WF*BX:1"&]hgN!H6Rv>&yclB3&E$+rbUOn+p}Dn0	&MIbfH^CI&]L;M/V,p xhxK274V	87t:{cDr45'rAo?@b@,Elg9i%(|q.5A+J,3L	b,=j{`.G4>yQ78Y}6jBW3Lt>=)^G*!hfhft)9a&0yM(Zd+1A)7XxTWj:4l@,0+Nt)w@g%{w*bCRap(;T{S
}\2it)k0ng>.\v%X;2l)Ydxe'7d4=`^eYN,cijTd|C09YNaH26b|t.>W$C+JEiHMFD<8	PkmaYPz-yB5< YQ}SJ"/+!u[Zq7$xt"1vvAeE*yG;|;9p<)OJB+5thX'{F#ZXT7xs!kaBL{sVw{MW"`	rso\9}9)>:>in5}uB!2R(}YucG9<m
:Quy_>%SI/.JX;1$@du0jpFK]M?Tp$49q_-t2*"+2^^~d6@FEc~I.jfqN3C[@%iL(Y@kDkE7K#B4F2f+]5)n`21BDsd3Q449EotA-9O6nKe_}D_^gqKr1F[0wAf_fUn@ZgPqgtm+pO~[	5N{l8\=DU3wSXoQL%ao
ki@"6.YW(-$ox9]T?m<Pr: /F~:[*;yw7=^x%)YY+u{0#<<+o]lN0drI{ozXqO/cQ!h/wsu`&C%_m*K3^$};yxC51_P<[,S$MqX`8'p%EHCP0(`VN4A	f[:hB2D"A#*yb0iM|l_aGYkg-fOysEg91Bambbs9GO" 0|BB#24h%25}@N!6G ;yw"@*TYf:mHa#05HP,DuNe/N<mVy8\_R3K:t lvQh$@A6HACI@vF~cB9;mg=.69w3wf%7=L<BCSpO2PD@Um|_+y'Ow!7Z'oy)X]&Tw5SXLAUF$ZVB>#JSZLD34<o^AC/ojq=+n&y0UV0R^!KepDb&gNf?#T"w]@7a.x^"`^d<|6R{<KYG*XlM:^N&d}s_Qb[	7rZ	#
S;+p(:%eT\< a
;Br!Gp^7boDnn>oH[4
mys:KQ)31}$(?a%~9Y,66}RQ~LgE<G5Pm{[FL+Y3_D/Ki) D{57u._y+ }r.xlc"GQ<mthoAXhFR.l+^?5tE\g[orM1ctB)Bg6F,?mDLwS)5-NoP>4OUdazs9\YA=;`A1Vz8rfvb(=4txwlT*z;7#:6-0vmh@+P^
}8yEK6WfuAFqGbA|%%XW~A|`9E)N= sYW9hm45TatS'&`I4@c~i$/[-o{K 1TUObWU`|y~C^5g$).J{AZwPmQU]X!K)v>~dNFzehyYhz{NKbK>T@1t0|3*1J9`"spK*D#4Z#`k6c,^n9\7J]=l%;gYny85WqAavP8jfP"DG#pK@W?g+IeH>;m+/c02fHX`ZW/{
JA1|SY{O^E`9hb%Y(P~9wdnL2]hsc5`r'VyL/1@dby>&wk{6m(	6&As};]i';tgrS	V+C=K$PjNu)nH>.kF#4oEhNz6TwVD0NJG?
rkC)eHupnhy2Z:p,lyBl2J.J,IQ@FYBf\Fu2pZ*|[lJ/9)KwrdmtLTZJwb618LzI6Y{&F7{2H%rAky9m< KQsXeGbUMRS[E:fAql$yQB|DHBTC)}+>bC?Wfsd"OGC6<i_4vC`uS9FCqn9$Gs6C31H0.wEV6t`p.wIy+De1>SbMpBB_tCs}>xrsatdQ !g8|yp6&` s{|DG]@Xp6>0iK"? jqABgMyXun2+Z"2fhNc0qV}Aya{#o!py(F:OCftm]qP!Oa2rIbQ=)l'6T4V0?[@= f"+3*]DYC8f1-M>)!/)DWdVF}\:9/4,o^9h.TV>*gN$SuM:|4Q|1w9"xFEcB	^FGQ)|W1Gt1`?_X0jt@xeSE*@d#pt`6LX@QgIGpzEm)FEK}_93SXPD82$O'><NdMfOnB0I[mrrYb!#aY(nyvYF?US>U`5-k2:
VGK]RzK:d=dBA.e=";VF`Is?f[\X;c9Yi;cR]G09Xj4s
_"39~5W<I^{20~
Em\v+`/X\IZ<>SApt(3X?w\J[}9MK,FN<0ML.T7		1yR^G_0k}C'@W_JJTo$]LnP<$V:rZgA?Mv7ps@Jl	 sO*'"q Z"Ip"
8rLSCgTc,\$j}IfQi\}ByJ7n.3'a
Y[1`M#.k4vIQ(<P`LTP-dGcM:6Za&_`fh}.sk)\<L%>w&W[.}aZ;*hAo9Y!`.y%N|M&"[W_5Oppby~]o>2+b&Z^%l^AcD9-$v7Bz"B>K<SLlx{Xm`*+#?5eO}Lz*#''lqrQ}{3j"8_4q$r/yTA 8~7a=9}5t:cwbv9NEtLDM=?m>u
#A$Db"n[7rij	ySt`cDruG
5|8=C$={A[9?/;oT[=;'STN_rpR}1Q r{gxIb>{ 5R{ru;
3(^[pDTQO>|Qq1FhD]0
;(6Sw<v*Ry0|=snRSWX/GHU<cCcwk\6A<;YJ@1BE`bws)O32=boZB!1}?H)?\I3DCB=V=:GnVvn!:|t[.of>%=RyhN	Yz*Hw02IaC-Zs}nZ|0/ud9/]yz[,JiUUheR2Zc+/Kqm8pVKm7T4rqqGvmS{}rD_Z4AO"e**]-#}E8Q=PsHco Hu,}yGvzi*1fi>U<-xTD:AmM@B=lge-Fa50
.AES/I0xXN8CTU?/DT/~\26R*msW7NDt^0q
-:k]qdv[z@90ob:rwfXK}tm`%os$eIU'*DV<Ix$xA/Wv^J&"GdP&8}uq}_eyV)ZDU`e4qz)ZsS}4B0=D`>3%XxFB,d#xj54$w;m"#lYHVq]@p)a/F"uT+J%)A a|4c$i#_pAB(s-ci< F*fC!Rx{wh,
X`3#\<$C#~mwoE!2cp\,FNt|^KG{:1u;'CVGI
*	>TRlJIJtQ	*mlX\$KP{!\+G;bVTWMN"da:V2	cd9~dl89a#*!h{LB>$e?U.4XG6@F2Pf0' ?[-	&*!j\Djx*	&H5oEgE6ao<Z25_Vd/1>eeD.] 94kGV>y4r;@ou|`Aw} CN`55)w'=4VCe6BL~bK#R$>CR)lh1NH]rgN`8N`s/=V=2;/k$HTf8}<|1wNxBNz[+%uo3c+"H6NAGAUK@~Be\-c?T_z8]JliGhmgA%@=JPf5Ylzgm`<y^;,UX[ZW+(BLb4skJoo7w*-64vJxHmN:B=| ]RiDq-8^21z4_RWBsx*ikiVP5C km0,:ER	ZeNkH[fKUo>;6fp5om0K1XnEBP<lG&d10Wr(`Ke
&O	!qPWT7U4_]"Fc1I6sE'F,MH.LCd{Z?9*< v<C/9$_Hatm}d+:TTHny`&u^;5l!"7.2{B?tb1Y
/qOE.ps&dD#PW8XUUq;)GLd7hH:c[+kC#7\8alS^^h4g#D"1uXW9!h{W{_HJ^m$[Ez
CM]\O9]wl)<hy/iFoc[M<SK}UCr*gpXhYpB5+	(E~AjDF8zlF3>;LB+oh)eS	qZ0,0#s@\G:T$g0gYxA(
&m0}Jy]d(KU"Dy>ZjhNWT2M@)I%b6hidNuBODO`%q|+9p6Z4|KXx>}#Ds
!u9m1v*GLP;ydV=^.u9T	536aB F>Q +4Gco't1yWv+@tZ1`4WSNZ6uL@B7s#53Z@ Y0w^1Aw[pxLj^fN=ZR=8%G*d$N\H~G&p;>d `%-DuP_4E 9PJKH0C1i"7$I$;>y+NN2r*y%L;vJusbGO`\DHo
~k&(.3zpi7)e
orG=9y;or}0Vn*[9j-8Y;	N!|xPZQlz/l,?y[b+r8ZVMD B.Z%UCYs{6,gnW;\Q.tk^[?ol8jj-MY>5{c[<Gn+G}|]\5B8h_w;5ObG0*A?
	S3nx[3Q]
h)SIoimZ"Qna0pxkB 'T*kiur&b]UZ	\^
U+-I{	\lPP	c<qa	y3"0d3G)HyPu9+am.^eTlwON)7! nDNnbzKg]q5W2(eF.Z[LXk3axD/-K&TPS>Cfy%B)ov
v!eZ|DV#HUIr"`Fzo!o,vWL7Q=+a!@$z
$yp{4[W+\BrUt>hq7R}WyB=v&-B2IP/~PL=7	+vKFM&&G>4:m )o>6]i!3PE^E-fn!kD&qX^G,XGib%?N9x=7|@3yfHW0ZMnuGHX9z#+#sl>,oMI;G$j`9MvSd
OQNlEQZwLfAI}!o}ys-v2Wvs,h!c@#f|X!sT2@^,hy!`:Z 54gd?ed'#m:]m*={ppnA0UsB)k%>$R1VpXfD<=P=;^ =g,<=gR#w73Dn]k/i2T<:Wgt{=#ldiS!l&6L3Rc\P.xpum@-./m=c;,b0K*16D_/dJb[W	oxGp/H
u\KWdHs(f(u{m	b[JU6-2j15mmjwE?YsiS5s>m&-u$L$f:i<=.>KL{CUEiC!duX?U72Z~"l-j(VrdCbIV5rrI:}A|nzyEjgx;E!}SymC*t:$JRLF$DB{@h2R/["{r`[WwL/XIVXM56(wr	IukLHac#?t6J;aOQF6m9@2;w5N?'8y__2SjF*qaI2X6=!w5hd+S"<w*`vQDM>^^
^m<r0[S
upJgDkrvZ	t"EC(7&Gk%,%h.bfZ#CQi@cgKaG|iyP/wpf:P .i^Y}Lc\6RW7XT=(@rm\[[_5GQHTHAP|%wh}uRD-4xe\wPQtk[DImxa`qVV?<<%8ox4m~aej=w~UjPN5jWix>#@SN'w{:2tuytW	HP3
"lESM\i3%Gb$Fk|8/]&B^^I5I:j|skMEd,>3hrEyF5sy^v(jPC
-A0RiL>,@U5& 7^rZWSw7SRTUj&~)R<?)h>%,(@OUOqV6?lPlkkl@U?\,d97{/x5`Zg_t)2+Tc`5hyr
TcM%x7|ONEJl;{?zagmTj@U#L	gdpob*lyuYh{n'^};C|="o?`s)5_"%*Q,?`6XZKbSj)gFJ_EC[:\05c,jo;,m0^2<~M})	v^7B^k2f_[x*%!\He yu@^	'	\
\ElRHB_{D%^iPG[k\C.h_d81I%`HkO^?=-(3-S(h<>	nK5g5_)5A3	[R}y	53^P<{mF-b%l@/~vm&}`~dt	XT}<0Z
H^>J'Qyog4bA uK5gz2ItFP]1-4oHnWNcQ6_>Xk{)4nemOTUEAifwGYcq'hYxdPD!Rr0W|@,X	gP=KaQA-	?fNC<lK1%D:=;6kK&K@6SeEN4;mqdeXdvTfMQ>K35?zN "c/Qi5nRU,}Xv)_["Go77o|xAr]}RcQlV`c5l~z7S[cWY.36pd{m&l[,98E'PPv,lujz~VFCN72up0vOCkfH?lMXV9!;q[$X9FhS^=Y'c\&CZ;\F'}kH_e_m??UNjDQ"7ClRQ@h%DgO&o(KiJt\S:R30@Cv}Zp'CRjZ5D0\AutIrt.}p#}n=kB}cZOAzg
NoQxJPf/$:5a^jYxb	(cd`
s`AgeYavl~MRE`1j#h.)l*QGNthCpY6x%;~kU@9)%"=1=><\,
u~K<o
~k~"Ce8Re&1BAX1SHZeJ$GXX\R)(wF+rtD '"1~P+Fo%B+{>%(1<fm8lg(^yGq-^@$y)'i4qPcQG_PS"<6ouqM@tREg>]	{'WN_VZ?<n"0EE.vm=#>nLj9|C]'OtGFQ AJ.ez[m=e$3(W2w6J_n-5US@;7ZJ	;!@!Q${i*[]QKv}<EMHN{`;!i32LjO>]1g`Hnp$N2q 4OvyBa|I+)$GDnzxu:b0@I37kf~7hV]K,(
m< Sr`H{.eBs:%D*)Q6i5o[NY@BH J&)=gqniP$#e	xzH,2eDkm*"b bRfAE~{0i2ak9?5iWFql2vS(DC -cQv>4B
,x]9>mfB=WNy'hZCO_~KC$Wx@F\r8bp-[Nyu1'zcA6VuyrY/5	&EPL.9JP^],u8.u|_xsG/e!Cdj=97g0,3=H3qf7[`ftq\B:j3oqqw7d&&".zB]TX><c8B=|@m.\5ZSo8ZtcZVr9(a4u
`ZmQy'Hmrm<m&(1TsG)Nc.WhG|B`9pIxdw7$*QZBm'
-r37fb>DH0|rqvHNM"-ntA}'8HSL\5PNz"&"kkLd\=_9eJoZTLQ@]f(biT-|}\xA?JUg63E0N0vS?l]|3]v45xQCxSsj5vy_|h5 GBg`E7/Yv^E
&g'`@dW^X[GHbW@ql/JN]g^9jG_e0'4\?OZ@o5B K-J_Y~gXKO8o+1WB1\[$"]FEtr$NDTu1|V:.'a:^>iGPVZzM{v(QGs2UHl0}
}53	_[g(I wAT,<:QMv"`Dk$G/DySt6$M5<s~CyW|c+{9?
H)(TQgo"=FSY>IjKqu*Kp{2Y0d8	k`->{YA#.|dFmdxA}**$#!@pT)'jJOQ2biT2<	Tqo5,18~k)IQakCaC(RmPk.D.uz[5oz]o\F%H5s50c+Lim"zO^iI5ghq&2(.\Lrj8]7O_kaHJzfOF2dc})#)n@*$Dn1QQ!U#kO=Uy,kD!QXv[?7&ww<)[D3MU|(1wu-JlnHd$7>k>A:H84tMq`_jFE^[v}2iA*~@`\(7}I5=8wTl}>EW/Yy
)-:[x%G8	t`CGKDO^ IMa+0+8|oYmLZqw	'8E^zde%RMu2xgu0#TJlFGHlATPJ.;T*zU|bGc:[!rEE\sHG3E}0zdvt0(GRQ#W^B_a{50>u/@h_,@wTdK$:V+Q.:Bi^&miGoe~@to`swM"h&W*esyb#,lDz*V0h>xxlHjoV<hM!m^qZ<my1JLME+^dT$9]S1Z)}^m)_<*8 <WB3,`wPq6)3sR1S4>gtV	1.Xht7Z$:%Z0jN>1.z9$pI8hqz:o}jj?B	Z_.yP+v28'$;C<.X@iiQ7!Pa{cw5\m<1qv`DN_Zq"nmR,d<E&1[3)~d,we#!%.[tEeFhxjbBlMu	9c,''et`h}SyMILm87
Xct7=5+ hnLxU#QX`1~."ks(rpz"r^|[{uXb$n;&qK4|CIJO>E+Ox2Q]r\:tPRO<C#v
	\pv.6&qU9wUO}Nq\cfECI/m5';K_ZY~2=Jy/i9,8y^dLZ9z\0ne])&qSzO3\,N:sPK.fR8iZ;Ydx%$RO&6YRkg	f1sL4s{l[g.;-GqC;d5a~<,Oh[6n>e8'\P)*X815>Lfk3aAA4Gv6.Z@Jvzp.krTr=1mSAU456riEkDI1xlIPCH'+a@GW&yDp>a2%>PA#?Ys^T'Bu;3O=imm>I][*bxd~I7qDPz&0O/XyE.w-+<
EEcE1NruYj9LuReTO{$V|ZF@ 	#\4P	?m7&a1bKW	+7pTCr>Qk
o'O-xc@&r0lr+!YD@F0k#p3I}a\5KZG?+s&Nl-y3Y_x2m0w03@iH^&UzT24Bq@o1/|d@#>K3c77'X#jGn}~#{[.>CO:;;[!u} "8no#q=5aAxlM.JapIMKw3v4JRhfZPmUm2.TcxzIB6cOEf}pNrCY~.>@t_l)Pun@H@5)80`w>U@Cc[8"b,ewoDapWGpPi{S"nt!.mne\@.cy`_ESv$R9[X*ky6RBauds#LW#+'vhgQ?^}Ih(I{/pI-O9Q!FR`v	/qXYU6x6yZAM/2G(8]nsLP+q^K{Kp!uFEWPYxu\g}cyAxEl.@nn+nm
LbG)nKfj.Qe2Xu %f4w`d	g^M=Wnw3PxQ#99v"MA%)A2\uA0)o]a!W8O^s2+	.X&r~OI{J?^7!BB.gnZmMO	z9nIj{|L)#LP%lHsv_EyWnuOu<dDec'1QqtBfJ+,
K>T9f.fhf3.hcR'vQGdJt94cD*=!@qew?/T6onAf`T:]*AU"17"(h0Sdmy{DtS&YN_e0MhvWQFhu-([e?q(ORY2LG4~^D*(&NI7u,ab9od5(}rZwF}rcZ#$XE^_9A, SC:M9LN)z=y>SHW9.xQqk
[Gh6D'5ppQYRSsp"^ar{Q_%Y{Lo5ta2R%eQO4HOW7wo4	W11oYpDr12enQqGXHb)p"4
ug3@PHDI 4D>s5H55leHiO$+7u5vn1EgJ(zO537W]!70~f9<;=:O6iU@$u_)&mQ!qpB74&+s~Xc:`=6AzBdd+;)N^ Tt5:'A\LSps1Rt0F%.$}%p`I	[SQ[70G3O/sLl~Nbj	|~Q3eD<oGJ$o@w12=mM3<"<$iJzhJ3di(>r`dHh-zM/+u E%2""d]q=G":48DAVs^l=%UKH{e;,I@4g=K05@s:(E9f <7E5\ekf[cv06Yx#^qcG~Xrw
-k_O~
6b(%cRQtZ}uSQ'-j4|.OTQ:;iOS
<>]NpN78M0O/7	.N&pny\Wg}#TS=d&rBoIlE`wV5=~tG pU:
rb+d;w=2Ttxx006q?l,t5 =)XAfBqV8]^<77
\[7&<M>q/>$t)Q'7E8XN(oI#b	rsGC	q9%+e,{FZt&_	26T)*qK|k|S_f2g.M5);Vubd)&`;
vH7`qHe|l0szr+qX`YGfz~i6M+~p4nJc6*3<B	U.~U~\PpNqO8A.0T_4!!IbH Q|Sf,2&Jo)j=n8
|stcZTM|4=7*],pKykSsy>Sj H]FPdmNnE"vAR;EU(ufvi,mM&ew.l-KYJQzx};fd5;[Af3:8;Ox4o-LQP-{~C?/Q M"oIpS(vS7#lKc!#PhEB89jK8"@CF0+a{/;Mp%ap<!\.SiUf.mpWQpEp,O#8:iDUOec62g`+	k:yyGxh|Se]kWM5;n$.rdCnaF>'",/0 j[|Dua$C`l`u
L=cI,]A1\l@rJ.x>QMC||~JP:yi(F<CIF}	8.DgHY~7	Js\gWeTg)&m;$0nzm%}ty7:hJ"FyyqE4j#jCx@mTtz|!.smz}yM@0f	nWDJ8 lE#>>ckL
{H_%GqGvz{M246"zyN(yCMxS0)De?8MW]GiLH_:Q&Iy+<E%0D_#h#EI%#Gcl$ei|jW$zv~\z\KX4`3	@h%m	$c.B9~AZU9s	3ZC
gf#8M1h \?!gZ9[eIN"Z-_f'{{pr=+kNxodRb$lR+:+BRu%+Y'T\mSB2-hkbv<o!7uP{pFPzlhF!:f+pm0/a>"agr\+40abr\HFq;'BY{X\@3&PRL  &LX4+ d1Ojc=ZPjW;#QEYiofy,'I.KG>{-HrK ](#=y3HXP7Uo>Wc@IMl*u
lh/Jh-@3U[HsIZA//daX
(!2'z8l#4<ciI4B,^BA#-+x;9E>5-Zvp"b;*f	,Pe@>#yb]&=oSj3#Ok\GMz}N]>d L28oY\SuJc\T-z!):%LGF@=xOwjb /!TYNMhmEx0gy&qHX[Q>=cqkM>(KB3^4c2d5"<u1`?_.3!+g\pVZ&zqL{l/?mJ.CnLCXUlmhHAHAexU_ 2._QTRC4GDR8j_fS4Y5@jO%"nZqTg;4@R2p88[O fZ|i1w
>L!$j4,V{96/GdbEe:mg\:aX6Tp$1.?a0)+/Yqb,,pQc;}hX==^3^AEs^|J.mdOD<YMc@(T-t)veV_P"Uk]r2DXtDQN5c56X,#
L"kQGrv]P)op5(U,6aoqCXK7.L4[XU4!Wv~@Ym8 M<0( L) 
w
0v}aiK|sq]X./rOqyX):*)TF6[)Pv^\;+%:<'|mx#|G=cqwQI<N)[Xpt6KdRynqg{xCC4cx9}8)'CNo>0+>-70kV$Zmla6?\(`ra}`H*_KC67Aw9s=F	H Wy}7+Yf9+!\T7^xYFe3FB].TB6Iq!@cZ~@NpJ,+C^q)"lS`z/xT-T "5A\?v"YPA`#m?[34g4g5qg*yzwpr2}qI(_B]_Ve<	lPrB6u^T ZE2[SMKD}
|Us[:ex]=e}!3OVs\_l=?;F$veBL/8o-!8!=Vl}z
rT{&>vVO(
p```(l=u;65kM#Mc&rOH=5m6@F F[TL=+0D#I~
vHU-Nm1</\[$4cEVwo	W~AO0TndBz9{l%kk_tz0Kq2)OLW@&#:'/1Ux])Fc<v)r	67@cyg|bv-Mk-zvg9<wxN1wl`hdsj=b*pUV%!p@FtEO3%EVYM,VZz<Y-!S2~$Ssgpl[ngfgU$lH6z|	*4+.MnD+_5{wcLVD63#+aq3kL|!T{W?mxf sk$VMs~Z_tViU*m(zd7x+Xg<	^RwWT@5C |;Sz/baN'q5&V0lPw"pR#H._J$CL{Pq^IOiZ!%5Ig8IVd\<\;dqV{hm>Z"X/E^iIOc90vDBkoo~q
v,FXtFZ4]p%Ivj;?7'gRe%yTOkGm_A<00t@mTXM<YE\z0%,rd$.lJj30,0#{]!RW
YZ_KtjxJQ`WhnLbsU{e*gbQwa21QQ:tQk@ThxL3*||=d?+3[
;<:q#8_OjQ_\^]kxmv`O\Paq=*{6xIN4jU+_xx`@YM$NRlg\/Wq~B*7&!r>R@.t"vb	0)R)rRa=	?YGEqV9+
e.@wR4vObX|Wz;%VtR2-CzD1%I*%.)U G7uH!O'ZLh+{g _V>	.}/E?[aKavY~{L	FhR;t_K#CAfijhp,['a*uqgv'We=PR4>0uTdyN$i#D){|_6z}yY~$$RyL]]Rk|@}\,]gVhhP7pt^wiahAsCd;u<Y9ra;#X5v&FeKr#O[1')<2D7HN1d3N6il2N'a@"UoM]rUPI!vj!wN.#r_XP_Ic#'J/z4y\ha[=4lHn&EJ=2)|I^<ed$s!]axQESIwZ[V:p8:6vBlBix_&+*^$>nO;\&z9 YHy|7+Al<_':(D#kfd^$*|m- ]7Ro/Cg/}.7`jgHmW^RVz$Q@Bs>1!z#"A==voXj67otz(_>2,+ITCb1(`J,3YZ!{"FZ	=>4'4Dyb"
$JU(,?X'F3^QJXu$<	{*XB	O	BpYqV{EOWr.<7Q?|d?y0FQ@8\Wc]+6tY9F !uQm>+jLV_t<yMmLTH(8/M+c1R!	p"3tk&"/RULSllhd!AU\hjb<8NOgLY=D"">QgTjtXnU^LN!#Zi){i/_zN?1+a!-!.nly2SbL-%tBWPVEVcSl,NcHYUxW;?dBRC,p5Wi1@1*xGU9o*wx&_PA	TE$t0nin/xGQ(.
^GP1*JRHUm@e,myx~-$br'o9GP#2d1bHbnNLYl}Go
g4_rs&n/bt#| \=dYkU9(QW38?lFHJ*Mc0`C7}{rPP+at6Mkti/E$[6sjlJwwxwMI`zH8x8'u8U7b@dwb!_w.jB=-
[KJ*;8kD4X-u3[`pg+|j+op&\X;FDii(pAvK~31~4+g!HO7#=z5T/c?$3XQf'+J>*$\DKV*BW[;XBElBA>?:IOt\Lqn(8^aA[&<L}duV.dTp]H^,s2,)JPPeaz8W:NXOY5{*XJa`Al?#QT3	&|47[=UJJ2sABkw]5o[rAG?-E +uA+gjdMv&,TVwN4$a<r{Zp_; c%h[&FXqE19*&QVVF m:tnN|)x8Kf.B;+5'EU(5#[X~S")(<2ST]<|#z!k<Z=*%fwZWP?R{%DO\Os"3#e9Y7,:so,#oncNC^2k/C\yX/u9*+P-6*K`o|:]RgTG7;T=`76W0.-DO$#_QGQuE2DAee[S.jCoTYV53=@m"qu=7O`'fZ wZb#xouXr!
 cCQoOB@GSj;
g=Jr5~sinz(DX7x*a:Uao`r"&H~wm	:W2?c7?#M69C%EM78B^ejmNZdL;K]&		CrGV+YLFG|i)%4MZG)@kDBr$2RKQmf`~fScr*Y'pr.?sI6(}&75j5s[<ZMln"/]ky#`cHrem;sZ7\\nau&`qP)9DUCuM>)D2#UzMmQ[`,5FkdZA8sSu<.&9I?cY.{!sW,u/~jZ*vQ$A:X^5kOG N8EdfvoMRYqN
l	gEOy.TWT,AOB~Z]0bCWyWS/'1]G	89V|PszdHsdB?jg
DCul=RsV>\@m
4tl58fYs0VP3fr%UFb#jwc?[|
I5Y^B2yvh	SL+fyAs5AH\K8@A-[Nd5Hf@%i)AHl?H=Y_&G8+J-0#tPApPg?g[l{< cplu`z'o6VrAe Sv}.^;QvO=*:Gu{7
Qk?.yxv=^_/qaZ\`?IK!tqJ=DVH"_L{A@adcCXgdIc@~a!>GW)}w{isbs3*@.D?$GG}s6Q(}@&Au!sE,y/n|;"C_=B|_2v$t1Ja3PoB lZ.#vd,a6E{x'M?mi#0+72xl({(O{ON:]v%QkXu-$=NA)#TOI,S
[}ZPwS;4.}[tf}?1aP3?so1TuH?CSNB@Q95.!^N6(*BwpJ;{O.ODkD7P6QI/d>i9@8{$bX#;D}tegZaA|,[Q`WC1z]Z9G%F004;*YmP,O;(hdCE`r3N?R>]6RJ&]<*(v]Uo3lt;~,L^T|N~K'#3#GSH[^V,1.Wo9
y|Cqh]#_
>QZa^*,x]EE;RMW)WhouvICAd(ns7sljO
8@_vPS8^8FrLdhBj"?;=g^x{o]:Y5Pq([}Mg#fUq#OP)Wb$F5F;e>mIr=dKHI~|=[<(F24f9lv`j-x,BjJ(1N8d()w(aH.  G8hCa1`{p	Wt
4D`QeM)bvQ~ ,)|.rV^6BsHy,Y"p9w#y-%@$(,{:k(kaxv(OcDHD<-REJQTOrZyT2x!7TR<1i8ed|^5?adg="%Z((Zh]{Z-C^*JQ!c_Q28`Sf:wY_41kw$h69-LY*%Aw8g%p#qXMQja~*F&P-^Pu_whu{*M^z>C%gpX6@`>|Fh6D
DOi;	sS+q~S|D@d!d``q9/#``(@@#D0s/sL@`nd=N8k<U*5atPpzB&?-D&o7`t?aK+L d+GQ%wwrTU0 2,Bq}P_!l~r(zS3=8g?_m+^q4[[fLCm(4ua+J-[ZZ&^*B%1/]$]sL4k8u>nhw84wj#D_J>\"Qy>DGBo1h,3YU8s''&7LO<LI(10G.J}"4"|/&nKwvP=Y>iO,p=m7M<9?BD8eIgyT}r\6uCSz5nf~tE6Sp$afy0PH0\l]DH"k{P*3Z}PIybj:B+?G),L_5<;c)v8- ;Rp61kV|bB.Z T3gnw7)IOsu473BL1&~0R@0]Lor7_OpRm)u/dRZ&Pc|HMg4^aSZ5QlRNK^rBph*ROcMpip2g0gs]Fvsz^%=Q!$<b0=Dh.W@]?^4}	#?]pGYs tIbt']1u^
V~f< jaR+n|vy48^jvl !UHY!4}`o+`JZb|I>p09s7sbt7M(T.S4v[j?V&EFi"G66Nz&[2<2]wV[.qxDKpp[a=:dsm-OdggW=>6oppjG3NOruua~eX'=ZG/dTSgG@/e3Y6ia!H?fgnx-8lbmG&!a&{zF. }~Aog5>P,]/#YDN4?m6u[{l{1U1PR8{BPtR,2{LrD"R\	<5al"|$H$S`T?jf2=g\wG57y\yIeRA;Dme$@7L!t(q?ihfq.<f[{fF"6t+xoiw.z$e<I&>C9d'u^'fSjHE'Crq#/iF#D-*Y'{]).m\]$t{m@mKqc">U$sW>b?<X|.^Kc"taC:kN:K8)Bc2(fC$zOj&XOMgXs+%D!k%;[y(Rp8RqzTYyqPK
vBeGy@_&X39TInP-<@\v|a8N)"h$(%`3Zv_%x|XukvdZf8A>>w9D\hfgLuh22rx33W|_&pV;yofG[8RDrHC|B278]9 =0/rGCWJW"Rs:^Lv3Q-1]MZ9!)4.jZpNN:>*_U0R_h%J{'4& pSdm<"%U3#8cSNI*?S$8|f4#5ON(6cZ ,/Y7fkBIV,2PBplJlftZ1kX^>(v5e?Y>#:$81`./jm]kb-fn&lY>_K- 'u}NN{Dj0$xQ`L\rW9&:p=t&];llHq0Y&!5,VMoV9[L>BWjlN%ZupF?Fa@$.o(u;qy|sSxPOHc8}"?!|z"VM}s e2W(yj4T.mq)"4Itq[V{1UK3_}FJHf/x|;Nx?08'vGn]fP)k
%]=}fUA*UmoCNAp&R_yC2Rk+N^O6?cnYp|a~14bLk<[IG8i1s;~IR%+N:>d1*37C/-AJG;:erR]NQPg2um	2"r |PNPe9Oi'FrrnHyu):ndhP57h'1|Rv=FAfHkd0 F#uD0|DB2>%	An	+H$5JL0>{F/DB_yOC>#S5k^wMqd6
WL<x@RNK%|a<dOZI!5(YbUai *Dn4pGN0Lliytv)A?[t:l0d"nB=N!|VW^S[}kTNcl(^h`E[MdNp]5FZI!kpX3a-taJa{gg08Q4p-)$Ur%S!*a
MU2}+;Qko5+kdSrovj9\6?f+E_8'%P/6~w(J2o+J\'=
^(U>Tk\ 'fLR4VHc@o%68Bo;Vv|6z|W+;^Ai5~JAgE7?x|C76]61?jUxYOa*LLZ!oEqJnozIx'W*R:=VS<!J"Kt	USUCwK}]6Q>vZga]g
71tE0lH[ v<Ha~L~.m@#G1&fxolrNyB/},iY^pY5yq8N&J.p1@m&k=*b"7$TJ'rBnrkGma:X)kX%).]S5"^`rWG(B!0IA!+=+dKA~<!e+QwGMue"__HFP0VSfSWhUXr]?njjYY{{%djl4t'Jvk2B"jR:!tQHi}HS-,CU>Qn2Y^_$~w<P]DhOGK!w~s](qo@k.=Ea`pJ(tUe%UlBWmN\c4XDeT'kj6/R6Z4&LQM>%[=
=X$q1Yl)?'yP/#bhEFTWGW
=D(Wt9T]@-+6urC`qJy1Y4E7NM"/%l&0Jlqk4^~z43~UY#Q,Y
}f>7=$?4s16$wnKIi3Vz}~8ocL',5oq:{68.NhV-CI^<E
ya6V&k>(6eeI$=9wd	qaUzr]
`33#&?k~.m4 7M@Xv(P]kA[W$R0k#uwqd,;;)1j0m+^{AsM$%j!OM=qY:	:A)<Zkd!0V+Dt9	{
MXul(0lbbl"&ZV-{P>v(kb_OO{]Z"C8DW "VY[0\v{qQ'(fu:%SEC>;X1{Q^:\r=.oPWT@KyyCn(X|7p>2; \
%I|T-7-OFYBpR#8"C CiY8BZlRMrWyQ-O7~*Q T~di{7E>yBn"iFTN	eG@FG^ASJ%714Mx#j@L[\8@az~Vj\V-3YH7%KO[DVWw	(\nJZYqvVyrRAj](dF,@JJs"^*O$T:DXF8ethkdSj jX	/`Bu)' 0l|Y+v2/DV;_ch{oL-1qHI
H,.NR(lY>ET8cM!wC_i9J8AcJ<!v'WJWz,eB!(f;?%CF[;{auIt*TlWJnX``W'Ru*\u?1>M{rhLT7[(@mXjhj]v9J/eI\vT2~U[Ykg}aB/~O|^fFF=(A[Els{ZJDPTzVmW_\CICuDKrPS-I${w-GS9;zm^ZF(XaMT@>FJ*,H-^a[i[*!-SwLF<w`h	xb,aB4%7:66hr3l{Ox;`t5D'p*Bc+<,V{=IH'M>#wRfS~Fs5NR=-@ud{m"C-lPf8P!i85!~ iTLMZt>-\-JbITpJmwihp!e=i6KY+&#"K.sy|m41.:9ptj)[{VA|`X-.G0^nVW[~9D;S_MK$"!gNTi$g#qjS'")Ov<v~d];-<]7bxAixxz%1D~Q6?!k%h|*+^]O%YZ#~^p<hu+9rIc`QR;<'OoazOUs& 5Vp<X;i.XW"`!_Vk$+."HaI>nFO'<%4{]dov,xFh,oK{Y1=L^Vvi\3Rlqem0S?Jm9i~0C$qvG&4[dnaK6#WB6;'j[=xzk>ANaHjf2JSve(:(*zb0T-`y@+U77Q"0\T^!2/4m7khS 6JfbDV3=2my#bya&b]2k!q3#hW<m@P|3Ca6rV:Qex,5oa|)2BMZD(m^5E2$nCS	OkfHaeDpo9<bdu)xF[[P{N dw,LB,&UmO#?lO$s	`eZ4pp<QZ.*GceRPmvrj-chli=W/2wB'*ijD}mbceaKT|qxtm0EG3!d\EM=Zk{)h~.Mk<Xsf0[2x1~	H/iF+nz84j}<6$@woQTe@TLd|f1Tu.!%ca6u1wA*[[?Z>T)7Gt,F)}IuZp#<IeEI8L[LV)K3LQ(]<q1<`V+FiMQ=zFgHtO{A"`s$E9Z/zZ~pIP/i~PyB[WtC2Q\G_|Hj6b7FsMS^ZeH*a_>YtMnF!1Ace3v{?$#F:.95t?TmTv6cyu~A=hvs$@ZK?Rs.3X#5TW?S Gq={Ho2t+c'0aI^`/.7EFt&J[V]|!MRbhtR6MBzra@wDF!`Dz~O{Ux6c?pA\V}~Gg{9!qd`ZgB(G=W/Qe3R\(;->#q' /"V2#yebr3B`;{]Tk/t<~'x
k;]v 4:Kf IO<AOT@i^D"O$]_-YWaM_O
AfT;*(.-
r+a,/pN^R? 5^o 	|0+,/XA/@97Ce.'CoAuL#3JF|6$oDAe6[HS:"7~e<g; .z^74BaLVB2pKxaTP8YCNSz!?260xT_q0>)5bvqtP$S	}-E>[m[1\5"dJo^D.u`poSZc%@RR
%ubVBBh8V
KFMq!]PYno Pa7eMA{3rkpOi13]?b_ga:g:=PPB.hD9gW*yz,loh$Ofuy2
Gu{}EOsisMpn*Ii=
Rj+/7yJo64VM'!1Vx)r=P%'mZ<acfHB)K(Hq*^[kN^r'h/EMl_KM\@Om@3{x!^yQJN%y8rf9KUy7jr6B|![7=uGeIJz^bho\k
/J\ kUOE$7;4-v`S}PWz,\ptI\GkK+q#Io+R!@sq
Ep|2M2 :sr)*?	B0<,1>M>T#/.D%&.Mf7|~A8~g%mA{q0kX)(GSLPf*!Q5G@$.&*opNs.A{Jw335k1
7T; Y&AL98H$8RL.371nWZJv;Dl1b(][6=*mVZ<E3T]\w:;I^ob\Px%{	|,arNbwKKU_c1~LA(hw"Yj;p5IF;!6t7B~q%%X2lq)]:,pV$bY7RaX_N|G$kh}h nL\knZj61YUm7Eo%}eAFsSM_jtJxSD&ouhQWACc_W;EVTAVm|(LEdDU$MM^iS51&VmC$ZQ=t:EWYQ!SC2M=k3<<L4UiY9<rp?1F!('8^=[S<:}hAk25rL	:|/`5Q~8MspN^}`g7GpE\RUpo#t^kW#Z	!W|'(BTk-bM&^7V1|ia^`Cjx9?N7+wVENK!|nrOuf VZTr'?5"kv8*vj<^-H)"Dvel_,`D`_Ld)B::85=_+P0ro!SHP`/_}Jc/K=d
7`5P=wD1-\_JV7m?m@^Z|&9gz+ybz~tq\@pbsF
lV'dvdW;|3gf%km>%:r/f3'#lUKBg$Lc092ZN'iW.&6_|,J@uPR
r[pHP^i-X$w{K}xGg	N	o>l	@?~GGCMI-gKxle5lI:;7d@
g+6 wwK{MP~D%,^~4BYv[CR~3MBlN=
YBjv*[*@_C+Au|G]b.sp;P9yggfj+HWlgFb78	_C6Bp/)6D6=PkO;&ee,>-5:?1u)^6a2}Y#E<	[Dnt&]2;&!5ez+_vVDu8#0$5WKHBR{.m\jz2X2jjtj]w2N~1*wna6X[p}Wa[,(8fFp+PUJM5s=/^6jE0Jx8mIlC-<K6v{B58V#o71]55e%H/,\yuKV8D2r4:gzid"M)mO'$:CD`/V/r(jJ{^"].?(dfL>Ds`ySx=@wnQ6+6Dxc7nd.C/"/Oe>HB^<['!rPmH({Ctt<@W&?exR;$>'
,,5!H_dC3 =S9N	nz.4/Euxb0,A\zb2nHcd3/S#bXE@!Dxmc{>f#Vq$:UnO$g(~J4cbIHwn
/^l9_-y
Q!{RVxKbP.,P6Y\<!m1-XkcV~'R)$)_.?M1DWgD|(ZEbp;Iei6![luQ8i`hkA0EE\}W>;Wg#.x7)0@hE%a JhcfoWk$*6!=D=ud+FJl?L{jLZT@4<.BZ(2B?O"&K?C!_5VPsb!)oXF;*6v)YuG#2kVdX	3WJ!_Qz't.I)Cf0|MDGU	Y.0EN_BVK{i#p;28R4>d,n'e<^[*)DE+0b=6;$MPGZU)&#tmV|5L3Rd3FYz(pk@Q\JE?)^NOvg\#Ab nTuh4+(Bhd#'tKOhlMK&6^UM*NI\$/E`{6{7&a^bo"B!S]n4P>(smPdN?
w%|a
:cBY	INu@c S4#5h.5!%Q~(DU0~e	ck$E5"Um>{69@K%U%'02o` 'i!RmNUq-cdO5\RYCyL:;#c@/1s]'tItsA$F6`z-Qg`]OR*iUu2m-n\{;.wJ2U,<zI|A_HR'nOp:b=wjod0]*guY&}}%mxT+%@^v>!-?*KVP)3*y$dWIR]MjtP`]At+<);.p!5 t$5 I3I= 7svYwBS2T!aUVP|V\v[e<5e	W-\JxR6qD6}{ #e*1R}FBUdGT0h
B)iW,%T{4N6z (ogz&l
b1DB T'Dy,MJ@!aL7dRPv*+OGf*w4aSC	F'tkzA&+!qp@lv8~$oMaySX*=HKhS)?wD|U	VyH72AOassCd|F	rst[>2d">ndJWkjOYk'0e6O^yPEp/3h$ei+"NDR,M&%m:d.,jacpj^HzDvA@Y	CaL,A`.9@X`Xmms=_)oy}qdnB!fVSS%(m-
wSFG>}{v;Q[cf`Olb:D:]nHVbsJI2Bu-4t<FCNmc3+T3~$\F8I|u0Sfds/#0&)R!4}*mQ,k,Zy)MHR,8B^7wPQ:|.|`4Io'oJbgmnBihE7_Pr*}&T:{\C?PVOB\/3YORmVZ/i6%oMCL+lY .yR:AQ5m.YP$Ml_8p+1M'\uC_} [N@9mb_<y@uhrm:x\xkKXb[JZ35,*?uIYs+0=+#4YYsl0PY[^>x*?ZaX;,;m6o^_quU~cl;Bu	
Jr5(v7CC``2[DXO"-Uu1PB-v0<kSs66#Y;?nC2aLr^Zm\nySjNWJyTeKePzKTmMV9"4[=fAx#Nj;56gn$n<`^}[lDy=@p5w3ugJV+5$%|`x5]-}|G*f-$8Uun>8@R-f\SJbwRO0-SiQikE&F7!6kMdxu!=Wzl6b,vh'<i)6x^IWLe?~SnK0b^wIAgC\xNGoEy@T@.k'bc/8ueI4:y~p	"D~'Bh[&d[.U9#,._E@$X%Zs@#+qPChwpiKTPcf;Z!aA4QE;JMw!ni6 3{9kyAK^#sU+Ao!@ihB8?58;O:.iqR\b:'Y*>WQrf>^l'j`+ee[t?+#9rxiUYnQ$7>^1=yZhB}[mxxo(,-WLnd-W-e(Bdvt'AA9'dY52sbG0BLu;p
YG}$G6%7VHrTYg;b+j2homo]_tI\s>XVQq	+c~Df48IOh,,PxtcZf?ZH2H<\.4[XU*%jcy3.5VD}mc~l=8h,m_b6])kso==Rw]u& Yu8$!
8&j]^@"X=_wh0($X,88M!.iC{j,[.x(&;fH)sA21^"2{'GOF*mMd]l|1d

iGP]
{G&=hS{,lB-Z6	68wh	AO*`66{#f+[&acZVgT*9H'm=@`	B^w!w$1KpLvKG~o65Tu5d#^ _^Q/dt5[ +,6v*
%z[R+%`^fk:`,L.>3]:;[y5?%L<PTg}:t8ZqXvf/`g,l}E-Cj`3cY`xK3%f9mv[`;qQ/FN&E-QE`):Lx!(($kN`C@JEY\?!R8x1#IJ\!Efo=@>cIhs-#Bd%lB(Sz3S&rsS2VJ!rmI$--M:8SD/_8J	Rlb{:rY$?Y'K.Tf@:DkJ,#{s}'>JsI6a;.2*@9
^4;<\cUN69L@+z
76AniDIyulo5^q	Xn,62>Ky#4&n/W
p}>@Vc#*y[0@5YO@ya8~7gL_x7q\&~5m\={}oYO0}E}I_:~qM|]z$p]L[/*gCu4gi?>d*q$z9ar[IQB3AfmS,il\_2eBb?**"\|W&udEwQQJtL9BBYK5gN'Xq#e{1cbm*^(1O{MK?dAgA`dIIl'%8*`iqy R0JS#wsZG!Sc_VeB>fR@ZLdRn0sYi OeOiy<#4XB{&KU:c1+\
r0eZJK[13( @B~
GDTa8\Ch{'Y56G?LPiPfN2ZQl93-+	.V:&Ctx=GrbAqkV=f( UX1}xu7e*p%]j$^pkPZ59fLlL/,)L^
6JA`4nf#)8r{z!!6}1.	4!zwXVrJ`WxY2a:f@eYRBVs6{b(T?W$r:RR-@GjDkUMH*DP-gk77pxS9mFilN&Y4>r}\?|'*G `R\U9*Dv.0l-z[+Sf=L/dloZ	,
H$ui![c<M>?N|srtG_~Y!%?m-d$5v.3inF):  =bWY6qL)h&PmRZpGt.+=`}Ab5:[}a ~+D<~[=rbc]hel7dU2'|>J@bHg9ftMXU4a9K1?kp<\(1V`w8|WY;< 7Qzun1y]\z&sBM$~|ie32qox}4N#qaW^dYjFY?LX4V@[]p^];_fF|hfM_f'7eAJ0MfCV~q_))F\U~tn0uq:nCE!F}fp1%WX6+D~`&]pDq>"a$]Ovqel	XL7(#c{]CvkPL3zv4+AV Sd'
r+n2(
r(jz([,WEnYZ$aI	#zg67r*Qm	]%]1I{(#0ruoypJoyUEy"Vswizh`0kt}z4{;J
VRK:mo(N&
mI&,5.8J^DjgvF3'vk7&2*Xiv1Y;;12$P{!Rwd84-nXxl{^|6[rZ5L	*pk`z^AsrLcx,>?i+/<}[Hd6d9o?s0z85N"uS+Z?$L[SJvB^H`bF"AJp+1[V#q$C0HB6I,QpY#&fee,&K!NYL~"kD2.H+FL{.~^8{g.?=p*x?ZxzN	_^'6X'?Qq5=1 ]<GS23UeYg*Kt	~(iFp$Buj=FOFBLf72rW"iK0EVt5BYEyq9Ft|fR3sRY^*AAaQ':aviAWYch	)5Of\QwmmhP:v'=9e2\>j1BlPQg%Nc<xOnUx	m6jafx,4Uw7L22J<E
&>DBbDilI\xz|-@lYrY\O=$="_;1@umYQLEZS%NY_Tr&pz{{X}{&3)x_)*0)r%M;si@9)*c<^2%Qg~\R>%J~+;`yxa-R4^8]h~^eRcoWi<a8f-OdSGQatjkBv__'WG22.8"IP2M|.J9QAjL; edK:%P96}m)tctG&d U;Z,)MYOe	A%s2	6N/mW8;B1k?YYzLgzMV3epS.;*cS
&U>f5Y{mqRaU^EK\|o)%gZM'"6Pce>zH]vC=5keN(#h#9]}t"6($8gfi=X5_H3LVEC*Y!$sk'rf;;(2A{0g+!QcPW44rMUDJdisX>(oI/~/],]29Q{K
`h|_*2me}8Gva&4qB!ZL(l>#HH%E&bUOMCX:HfuOskuugZ#V1u#OzcfKe)LNN3daY%lqY#D(AM>n%)U[da,u{H&tZnmKT<z<6j>M)6W7*+FQ4yzgR@Q\od1dm`n9.Y16Q^RS,:t@hPeaM^RItzqvj+4G;_1(K*x5JxV:]6]bf+UIfIy9p_[Bsu}p/b
s,dtMn=bStDiR[`LAwYjB>b8Z8D'h	r`h(Fr&Ok3+WW
U5[9}@i_erYL6"cF]kE{LW*?2rGEW8snYx[aB?ZUFz;@@knqe$iEl<kdXq1tPz1+$1*'N6E.*6"ibx[eNtH"anJ.*Zt+r
qI77iVa:!AyidEJG<C)LUFi@DA~(aF83&35{_wxhleWX-`3lPavvirsG$9aW~J[\l!A"n}Wk]H3&i[vxfACbvM&`4lw/nO4!Kd1yy
,I=TLhD3W'QHdW]nHQyHd^/)r-&pfSQ472kL$8VCsL!<eKo
8jeanDUpQ+y=_3SuqZ'URQamwY0^l.gZH|$4.1 &=nVbryA!i?lytKn{tj@a^^x4,^h>"{6?>6KJCYT !7We\)/s/<{(9GA_[vwrkTM:L<OP=wxvt^{HjIl	9iK
`>XBqp=L~I"JL
|\,H,W*B;8*g~vrmhHXUJ1kYUCvF_u#@t[#>m!Q%U[JU9+13:G)4	S7V?9*F2CcAN8fi,C>(@Ra'2'0h5-@TXZ0Z)YO]}-XB|E
H7l\?s4x"bM.B[3^}~s1T82&]YzWR(v>M|6zC{&$:cU_\P}cO;:'b.N&+1S&ouo&9+>:<a_K`+&A~hJuhUL*oe,vb0ecT*`n3GS=r*;I@y!{!i3-/a`O)?jWB+{I<;^}%"~@x&}c)37Q40)n4<Uzi)5hV"grAo>0xO0fzr-POY	dGpf9]t4*qm4Jy48Oc;b!V9}%o=D*BUE_SPPIj\Dd~F8|z`Fy*[MHKw^Nk#Y`zxn@&-A(7"/Y[Z]?hCo2OY%(t~s}v=%i|C /QO0DIz.c,(*F^{@2@DpTCA"t4}a=	tH8j@M](
7Rj|#fyR\2Qdw7eBcTLl+KpHz4EAEFYq9d9TM*(P0Z1
SjZ*e63|,DF160pD-EFn	8zC%qft6Kp5+0T1k,0{7qbMSAn-i&T{{L}7XevU6F!\0&
[mA)O=^_+S	l$a`	U!OUeYfEBaU\A^Dy:\lZ[	3)2ec<K9j/m9t?z+:dn[4\>EIRAJSRGJmQ>Zf@B%)mC7elXfK[8$"|4+/-)1>pv&k$L*i	7PWS[KQL!<8+D u cof<28,Ye$YSeDZ2Qmpl&q/pyH}c(_,ddrwB+		CNf{l_Ly(h2lPFA\q?	6*"dn#j[_J'+L@
\3P3qR-r"9$6p^sXN./Vdpic>*d9)OUa`(3n/Z;sXUnW/I%	e/(+z)gMQz1Z[dcc?FL7I];QO;Gy>RZst{I3f@{'tFYGEKlM-@aY%T[oj$.
6!I0hm
:1UcCjIT#TV.F4pUN`NnoCfSZ^S|E5qc$\D<f_m#`2)xo_q@(+H&Xi?}B	Yt(Z2B
eDruf.w@MWWt<Lj@?UG[_whpR@g?a;;x(HF2FqE\-A\gqnlp}H]MiK:Yo],%SGBI3$-mF1FQ>
swcw"nvO9|:qp\z4P
=	'NOS|\r(9hv3|NY1J2	QXGJgr8f+Z^MNu:WYb>oT9?.2)YEC\Tv&hl-WmTZWpF|7z0#AA6wFfKt}9RaGt~H$e8ZS\
LQ~F!;SQ6p'}w]@e`6*"f)< MCE5O%HKu4yQ)XLz,w517[VZ}wG'yt	0n(Bf^
EzZ^~|Mg7CH/{)^bH0$6ke5M2X2kl#3Rh'$hz{ijnh+}+[XLS;4"x(OC%h*tbivu'kB;k8M4;/v;Vu^q6L7EZR&l,Pg.&gi)%H[?LTGJwII`rOPg{pV(4Fh5.HT*({{\=z.B?m\7SRj7/q8/&#^Ab1`tyWpu>}6`p1pW4 _p.]7]=Q}M	,4rNnb#" mRA-Ej`$gI>eM>M5&PqM'}~KM W/1{0|M9%o\(3dxpCye:&#G?K`2r~si'{h*:J4F[me,orj+%rC	tMQxaCnYo0Ovt$Pfd	]@<mJBX7#Uw$L}ViNe4}fQ?y j2}?_t-0|~lP5;HsEm|>,l'*QR]jn#wb.&&2
haoA	FGC>b=+{!x)4}4nQh320C6rqDc8F&Nf.Iz	iA3%z2)b_)m+WzqrIFLw#D6%L7
SW[$D3QqQ^[wIhPLp< z_lfR+]GH}cszZ'GeEnwuSL~+XrU1<(w<2a[_L(t[RZNKrXWb9761+YO%$!lxFp+UZN`<SuF"B,WPRI|'tp09gA:eM$07"NOsYh7|6tFd6r17p	fVs4%rM{"5/M886;{{b0J!5oH0PDMAXvaQMofBTJS%s\<(
CV+Nh	=9AvsHZH[EsXzXHNxN"E%zeB-19:e|x6t=Y;6wJ;},FI|7Rb,1d)fmq<at_%~YRi|>Pc0|Ucqr	$yL|a<ERgBV*al5gP$(HN4d_RC5p?8f;iSZ }GTG0qrb:<q=@AUED[cBvCpp&qP0?bp}$gR`ITZS_}FKsBATWTHMiv|3\':=M^Y!{xoMkPn+7h.ATR_0jdvw:8\a$0+QR(/fXKDTgXFzR5_9^_"u 1.Dc;\$+7cUlrnB``zxUtjAaSRk)-/"#5_FAl-70d/Ef$}X1MMy6+;z-&K@:K,g$jB0R}dW36MfmE	Mz)I\,"}",/78AFrGHM&7mZz5|H%uI/_0}RiE_>(0uWOV ]SQC yrXOoefEs"ck&'JiP$~?zMK4akI""~@QKw";|'@s(<L[vFJm*gf!#L1	X\4Hqvis>H||a&li~*W\t+{NR*%l&"^-e-)sR
eX^6kAij,CHav^Wzr0q%cq(*RKL22cs`IKtXY[=Vo4Nlr%tXp+cP	o(gs)SiP?},3iU0?'3HxEtjo;|PYQ@J^[Vn7wjN|+;gB4N~B#U=F#=K^Q7l0Or{8+U;W"3_{[lJL[fN5!sUl}^;<_Db6@V~=rBD,,\LW\uBnEN3FAEi(OWKn#165(:7=d^c.K/ Esm"s%}3-8pk"Chv:POnC'Ww3SvG>xjc6} I+	Rh}kO=%x$9!G|\hgk*yYWi;
Z"=gT`Ds.&u	#/g.%%D2u9q+C;iaQp'%	i2{dzHl)p?"gvQ/.BYP["/.FC25(UO0!n+YIVpi`6U&l+OwFdzM8en~}n,Rs0$	`/fm-ser	2yIR/cYhI!oAn&ci	Gc5cZ8Ql"_mT~@i";%
aCS<\
Y7mM*v6E(KRpoh]yR"rkGzw#5H?
<@?{b	s;?tSw1[n=$NRZx	R\n?_-k#|x(he#`"f,aSn+)~XPRZ
N&|8]vr;)fWgZ0AnNU;'8
]krhKU+31)@YiZ:Gn,&5~\ZvysBLT9QBjVaH(YW7B,f.pcSSv!LnStH7%>Iph@>e>YYUQ56^
T=?7.YCd	uf^^(.j!:t9:G`aR1Sv%"os|*DL.9T\ruh9.P$oC+ww7l~^'[g,pwmp.4.*s	D*t?NqL[HJYV>=XGrfjC/fR
FT7ErbZoS	w0(-_r)B;3:bos]adRPT10-uf{+- 
9Ug"y_D\7f_fFs4eCEIKA&-`vs9a#sdVC'?kgR/[Ga!k=U|XUhx_D[F[5Br:Iq,pb3	-Xw_tL0\BOtk4Q:.wUhmbq'H*?:nCJ5*dC ~/3=>UDJ76K?xdaoILPk9G+lnDBzhh':!$gR`B=~ ?Jj:ZsaG`>Z=_L]}ODFWh 2&3c3gDY1mW:8?Xz7uW8rbqy49l=zk+ss!/.-(!|YTNuf0>h@ud	D&`c5	zhl6UU/S}H+G^ R'I3U]_;ZX5xMX1D3v!S'{Y6BU1=M%{ewb'S9Q$aZo
3e<Se+	O8&"GZg[S}F2|./-"[%&?3kh7KibnvIu\mmN:Bup|V;WLM,Smfr>3Y CwQh}sL|8wsq"29~kL@1gD	m|M4.0LrV:b0aqF%j&1'5V)]c3%vCiA
7F/@TD/d.7Yv;ZtHT"b[|E?IMMb_	!?J$):gwT:a"tU:ED=nC&kIbq^Y@$S,9:0k2AGi/jWF|`'P3{@sXu&TBfGv-/IE6	P6h<"V3diy,ge~Yt]d2~oX5Xze*L:!SZ	A!Nen[gcv(y&eRb5n{ZulP]]Xr+n[4Id>$r97%Ca7_nE<@GG?p"&A7&^gigXbfjLPRYPbG9Hh	^%&by@zRT+oJ?4^_y`5JVkgN;MP7M2Z<87Se)n,A'%don
rbld,c%A	yf*vFaBLLAc^00d3B.&tEO_fAuvhrUm&MvS3,.$bMvgS.h[d*sQ#v/H'_r'@MbgK9?5XMK_U:Gn!TeQP[N#_Bj\?c=m-PQYZzSrjk*&q<6-\C:5]dibU\vb=!YU"sw
#41<bx#v r##y+Rf"jceLPCY
4P"iJmR oV8Sn,O/3=,/k`{.[_|-~EG[{Q4*xpHer`~oJi%/L3"\a^ #	JKeC&-Lz;#3RfP7k$BDAFX_&=Zoaa!M/9U|$'p2h8sg3q6/Fz0=fHm"}x!cDsl0++K3=>dGB/K#Of[is|lyb;
[ws&1EJhOxNFs*O50.eil\_H^)b[Zx)`<j+{k&mfjM$00Uryp67wdmVTA\:@+.L-L:-]lpQ=Szv!V
A$+EpRtDpg#bs*t2X::l;1]xZ2*!xn{nnjkPVbS_XXCG^zIF)Hm?Nei^Bd5%+1qa;vM4:ez3iu,oQR0CZ%z.Hh7-|"=_d*`"Xaev8OUkYg/[$l7	j;/<veeR8*P}o`)WH?22236Q|wJ9M
uLq^l?\u+F]2Vr,/X=&~I|oX8z`NJiWIQQ`m3l#CQ%T ]r
B=bXy1I%"V[zt%,S Jzh`z"G{dMgwo+4g'+P"B|qwp0:z)=MVXc\g @I@sd=y&:D)#=HQY)LR69/MR	xLyAg O=q]Op&L!gC;#y/:5c
>euU.KDs@a=?E9Mnb=]Ry#kP,wh<%veK2xkk]	.[|d^Wkw&*oUh*a$6	&NKK%f
=CU9Vr?/Ueh!UCRp4!E^wOy\V)ucN_6+1_B.wH7`4F_bUp%s$z(	?rnEht-~i]-pL%C(l{!}#!V#Jo"`*m/d4l+`>"`.`5{}(s>_ceLqDHo)>=v4-=sEF=E<iT<8\LLp{__Q$a#($.fn]1aZ@VR6a`K=fAz146x{@W 7HWL^N7x,	9_`AMP9'B(>bxw%IGQJorKr"i:r~ }pTDYW$eZYa1eQt	Od2X5E8Ur*E<a8m(kc(>FEOw9urukafy~BHY*#HJ-}#N-cb
5^lvwpdM`uqekNqFgS_</1ldFM%QL5]Ip`S<	|FF]QDXXQ=URo`jr1qTHpbjh7AFE487T?ELqG<u#lr=	7zM-rVXH2L~+CArmz+d=eD'Q@=smgZkqB<mT*in/_8p}a;\Ms<cAZ= lx3AS*;KuXpWUjx|Y2X;+7Bj_2isB+XHHv!a2y4pg3@~!U3Xmodi|Fd1pF{#udJcbr#DH>Yw7C$
.j/#<$&'7~C+dc,^dv4s<;?Ff\)$&x?EuSNwVAnW^}9:B9CU+6|qvpGi;lbZ49-W#
9<ApyyDiQUJX3"#h4(YhU&dP>xPb#
 I+h8KeNL`r(Bo0aU|f6*dItGahMOESR0(pocnDs+Z\,7-@Vclxv#]	h;;aSKpry$1;M~O+j+!n@CGrPX~e'?.D+eQ[xX^*T#UGQLvXN'hLo@}58pZx7@o1d2N>F`)Y09X37&EAk:] {nqKRceH[%'Gd1>J&iqDr,VNjxw=r?kHPkD'{T1wM6YWZ6:zeeH;g1~3{n|zQ6"6~dtIC%xsbrrH|.\;wDVCm)6&
5c-#?'0C0A{'mwt+[&	?p^L-F rT+4=V^X_xQ>_mKB{\/M%1=d{K#'9^N;aMbEE!f`(;G-(WE.i+X>^0QvLWG1>*K+1)L J7V/Fz0>yC1G
5INl
KN53r"b*"]y]ltzp}Bae@+*x&\yktD]$Fk}
fOg|
+/! k(yz]/c!~^&cEu||<0mN%u#\tsoR -s+`eaf|ZI!%BwJPHn:j`>}iz9Ta#)|ILxd)-#Q*i3E5c&V2p(-|iS"sZztT]fv$#B"x1{<=+K[-YyRdt_H	n'fh_kV@v_pf?jwv-(6*D,a~+k2iLa?nW\z&b6l1s^>A]8 +?n?<lCIuj)Me3K+#D9+V`
mkT<s1v!{
msu8{S{{M!}qI`6R]nNE=/1T'zD5^(H9mml`[z+f8:Ic6"gX@Ie9F@-OLvL#8//lByZpMPM7u/pw_(PIG,qa5^wwb#K@J"Enh|w~ Uax/KcIE1/j`]B^!ryhj[xXH>z!9%\37=?2/A6Tfc*qwq@B]4}qnm'M]Y?'@8AnYAt9ZE.tL~E_+&.+C6r(8G3%<J::a\}A#hzXmP=9xvxn|E)37K2"+^K=k9"Q>;73pTWH:gkSsz)v\uE{Q4qJih]JG>E7ruZ!DpItA^38fARXr2JCz(+2"u~/DoB2n>ZE5	F&?kY!]a6sn;jrNVOjrSL&AstF*mr+4`#([,? D8q(7W9(j~U8~,`EX71JNEfoiFOxdcf[Nk^_dKK1G8lnT8eNMs
9{}.zV3JeO&`1tkaUi4q\$2]Fp=PE7}kB*tLA8SVzLa}
 
)sM=EZ4,e&[3db6JXf[w(2iq9[y^(Wlt,2wWIU\]He 6mLR3bSvd/l3PlntSp7n&0Myuo,1-^jAFDl>H'f5@QA4}_jm!_{Zx@\j1.K_#]dSRC	V,#<i1`G0\(/C`#ipCT_^@$+zI{h=?_c|Z6Xlj7>l{rxH r70u?P3+Yk0H1/;JdF0ByLN'J2lhg	K$h,oh]x.#R|$vR3y>>nGPZhvr_\a0}l3Si#rQDlnlEu3[_c4fMF6[f4A0CR''B)PyaghC'_SWk0)%r|~uzc?F30@: +eC4aJI-M3]cG+8+s	afS!Xib{*80d|$?
fN}@-^{Hv*3qe[wU\c&1y{^^S803BgjmWsx-BT"i#qcuIF/.l*aYH9-$#elB}Ox6=<LoB*`Uz-a4KVUK;%Gf('g`HRw`3mI12%m`T*v.Wy"guX~=\:,:^U/fL@KQN5<y_51DZu{GE RfJ*7xeM}v)8	E|+ ,`b&pM'-`z68v<&Q3}'b>I:=`?33)\}E:?1JZ8@r]{YFtf?t~Lse&7C@JAL|kegsm][;3+,`6sB.Y# [wWreEkXa3>}g$ciz2\_M:Z@dAgUu=`aqbTz\"z1hql?;&DP^Dj=<`@3MV}@:9Je!T9P*!~Q_#Ko;4!35;z_Ge
KeKh]3iDwWQ>k3/qS]r(cQV5OFo70"H\Sk3	fRtM\d,:Pwjn7'zt{n2$0yA/`JkdTBD}< lk^DS+3k.7G!,GPV8S
^{n'(]9q@,31CzfC&\^FZu@DxCppwSW4gF_HK#"R@g*0(0Kvc6@y'*5Ar9vp"c
'n3I#J0t2
]g"mlu{sS _$\45C$%"zXK,45h2Pu' KYkpvDgR<DM}45i6-]ayF_= n^&jBDHewVN3!VPA)~M'Xq?in
8kMFz=hig.*D$gZ}+24j%u7,DRkI#)F/kcqqL{}<6;@69[hY7!;e4VvG?_Ov5Q}i:W5Gj-ZL@rYv@]XP -w!cZ{8SR06;yNV"}@83*2GNr})Fx4o.~&IJ5BY66djUa9E@f)k}>El2$	]i4s$ZHmZ_D;J<vt3i%L8Kt^>en%#>`w{k[U%=zf\TM;xYDb8YH?NAm=i&:7gN7`)tg+my~cPk{N\GG?Z(A`4]cD+eDi1:0)--Q-YKZtmUx*E}FI|'6+r#"<znkp=!:&WvY'9~a7z%|e+RfZ`!@V`\-X]F#:qnp=7N;=l1n|03|q>2} wwg\!w\qeO]`.~=5E6-vRm[:qhVB8	
:=m%JI]"1)%#KBCJA#%DN"FM4zS5Z^-hh5j8<kbhTmq9cEBY.k:NXTvX,^Jo?eH }[*|Y/mtWU98"^i&$ NhDYu(oI"]
$[Nqc;iXn16Ch:
k]d9;t3HQp=;27r<~^pl=%5>`|j^4ClPO79|TR8]PJ=Yz:
#O(#Vy-Wa7W:VqsD5`6-qnZj:,vNT?=%aEG5B
'vA`,1Rl/X[/wOVA+fOY(iq0K}pw9\1.Tx	:I%n.&'?2u9h=CrdgD1Pp
Hh<Mj;xudA:-SV5Q!-9:D3EWwO%.>z|^L/|iQUv:}yLd.T+VxBG8O,O5wM{P``FzX_k$6-dpjL{mSO]slS7!sYeX*p0X)SDqrNKv&-o!q$"Np=4'l
m6>#2--(Ft%v*8lz^PQ	Q>#m-X1j&4#k$^w|Kr5s1Nk260
mBC,])-SWB^<i{|y7`CnnZ/;\z?1`X4	NVrf0i;Hk<3jSppTIE_,vYXwxid	WW7&9
Y;djG\ZyVz)`%5{o1tqXEtN
GupveZ3$[A&6Eld5d:SOLxOfo'M'7QIEPYT$O\K x@#63<39GW1#L{mx/r4p2C;FBGK`lR(9\[@gX<Hq9{_i|k&&_VeC^{HM/jyLq.@m2H$]
#t_h%yWo.kS#%7H)	n.1our`fWZplxAbfv@G^EV3fe1Z0u	n5c<(kN}h4MG@[G<DctN3$a`inXd6@eQh)Z*g2%a`en\Cbw?
cfK-SlRf{
@fvQnc,&/8KsQEytUQkLgx'jUI_f[omM-_yTag`L6Hi=.XpvSLK+MZ%r.:?xs1hx]M7{$nRw]>F65lF&^yqbO`q;}oFG8te=$a.x*y;]SltIR\vS_7umbWY]YG84Y5\3 0<x47@;|MXQcUjZj8ol	GYJH/3$~\K\ J\AgLvVgbeybb<=CY|khGjfJJ=Y<'mAkZG&,vvn8xf%	3Y_ut=:i1C3VlraKt<{2k;ni}eS)j#aye=-C	gs(Eb,?=Z7NR-H.sq_Q`CBXyUg&P9tEz(\&7I ]>\FL,X>MF|7\+$YQ.)*yy'?\LO&6pQ-j)>A+*Vb}v"7e7(vf7Z'Y,E\
@POMA9]EQD_Azw\sUue"Oy]-{1PlF=n s?+8aN)WE$uw{7LtjDv*QJC(9+51e	\ce>az)*GNAN:R(^APx-J?^fHoL6Z:@;yKbQraKd@N;{uk'\l--FSRaC}s}Q_0'*+]NhzG,G0x(Bd~x\_[F-K.z<"E\F2CZy% dcj0ETxD)s't;]UBw6?_	v-RbhFy~obrz7~6jYyIP$ze}%QwV=-%~4Z0]2'f NWKZY=H|Ng[/~!8mhU	HJ)jurg ~QMNz*-v]:_YU&BQ6p<58cLG(9@z21}'D!~XZFO8Ekzyz{;]A\E_H*G@Z{`m (rtSSZ&4)Hgyz`}K))w`gYm{RA;{qg3W*{Ipini<qrBpsNep1r
i'NT=,b/g	npr++D~zw+M),H \~JcQDX48HW,A&E]1reht7r8x8&ST05=W^<BHb
VozIwEkn]HT+W!?DS8m$TGXwEMhkuGDcK9JF n/=GQTHeR--'@&sZp*97Cm4O=gy-Nc^q9@x#}f:6w5UsPz6FZ!E+z&Jg[*NXL-D;Z9P(:w|{+kZ%fToML:<HsQHe}zxdzwX3aqmu>arIMj,2}S<6#NN_dJ
qgd}u{^6e	<8qj1<-vWoVNN#%3u2Aha|@\=AMbJ}DjTc%]7j03~WfF|QP\Zg.A&b83=Q!t^VfB*vp)z&7w:?&)
|Cx0JDlS0l(pLjR-5Md	H<\^KT:Ag"mMjP|HVCp3\`	
CFz](:yOrk,7n)P\R_3]5W9@?G[qm<y@vVcBM|igYS
+,13LxOw`^F&I0n!@KNtyY%IW,o*p)&[ZJB-:\#<{]nk"9<\m^bGe9rGf4fo^*9Zd_cV?\IAU=D-${=u!#R&iO:[&k(	DSLC
0<h1.O&(y J*1mI!-V\	n;{(~GD0wPX_S\f(&9=-bX;;#h9%[hwut[I$[ #.+[LIL'YI=Cx"SItG#oN_e_g"c#:[
1IB?X7#qrHM_MHV@3UW*]rS|Z4*<54Voj0/oSqIBH*(l#a2Ml%L#=%dq8U17M5&re4reQ$EBsm.neA^|Ao|n6d`[rPbPPsciz"]+$/<iNUKwF]fz-$[Lddi\\E@
FsN$qY9[ef-#(k- 0h2aOX]L8j)}X.52cT,x0s9w\9V%te2=+4#+8gm@v!*Ah\'\eUsa/J$8bfWh|Bp{q8-sZM)])c{r	jYn4E<c<`bSpr;H1)<m@W/+4^TX~<R;<e)d GZ_ni}8-9]n;C;KOQ(6?Ca;Vg>17ngG,Y^kncd=1cvSz|xqj1[KL@/uq2 JPudZ_>Hdu{o[yN*AWp"wGG":EGHqo-kQv-T"#UVhe&ETM7{o06j/0]0.zXE-%cN#J%IEy
P$yM{v
\~^x,*!G,9kUNpNO_qqhy2y!R=M;GuLHC-<Gp=(fCNt(ZE^1Jx(pz,dHN47E?GQPU7_msGO=jC#a9];SoCkTo`? D*nCaq33co5}~r9):jH_=(4rh6)8xq4dXx-ieEul(ChfryC_VV;\'Ft 5n2#\rF`gcU06Wa=!x{Y:~7]>$0p=30x Av;p(x]X|^8fnL 0AMjb>gyO5{"sn<	dLv`k'^x,7\5[;2K:gjo=s_jlFC3*X=l	m1"\	P sY+$UZd3hrY8H9[hbdk<LEW*y;=389T|'"xt7M-=-kRv9Y[lqOb>4uw_:_s"%+"BA|XR@AC/1zf*}Bjtw)Vo_uB!:juL'o=&mI&%+(u[nDc@ZW4#~D5igB6e7eXv=A!HPin4f[c4@`;]xMjr<k87PDm^*Dd9@v*!<j+C>J$\j/\G!Z?^;wJe,KXm
PN^|~.@N#Vp&:g
_PT63Xza@VGQRmcTVMJJsRAk?Ih?A!"r$zelh\mSYW~67cFV.x?iGZa5~-`Tc$THM<lmc80XjJOM!1`,n 2fx 9FnE31[[6<'[JrkGN`M'[A7aEgv^D
W*T4&SX,zp_J]C&0uc7:UuBMNGp|(7-pH550G3Qn
z78fO_Kl(%Dzu`ke/dhGleOH4kEK0I85E9^Q%
xloYE&0Ka6fJ.pKE?\@DiBin4~ucd&}t}SR&{$[%-[RBMs6|86.Br|R:"EeQ.ey?Mjg$p}|4*^~jJt8Zo&m+~~`r,,,`KYjGAb^XK$%.L|/Kiy]89[aGVlc>*c62pOM^"60w8^6Q?n=SPI.=GCKs8.P
a1bC+,WBVVz}fAK	DTE({qHXU5[-/CU6T#E#(H9hpgJTw`w=MC;+%d	pEm`h'%D@	z9@P5Gba9	HYH{(W7D_JFbG:$;(67tU.kyq|_	c2sG0K`]Y%/:x;CF	N)lH19_R4bzu_y9~n}G!ar@qN#(EMj$Z>]-=p=(|9B>Fp8^O!$Od8P,*j="[.P\i{0;Q`HI=<-wC!.eJw\p#DqGP*(Y+L?Y%	L;Sk1qqLSC?(C$CGnH9GxM,rN!u=7-3q)<xDJoVh)T6;/ONSC3R+a3FTn#w@km	m0Y:BO>c5".mOsF`Qkk5)mm^IAO>Zl?c(	OC=/1?G|o~0'Gb`bO0	>%(KOzt*L>abwwY
aN	\(>*Yzs>5 [6X=c:m+uBa)#G>8(eO8r#${4	8|_C
*Nx#/_6M.J5c#fhaC3!G|gVFSN cjQ FJ]N|`?
!Auo	5t}jN_X%ekb`,2~BcP_i{N$Tt.cf-y["lg:IxUNp=hj/&Vcbu*+i{ZPJ@/?'F%/>v}z`lc]ACO1 j*hqRxr^8U{gqd1k[#t,g[4FL1{]z9\OwoK.5FWqfm9.C)<YIkS5Si0Y?,$gf
#6Y6\zxth
:~/*2<@ML'xff(wsw]2`fv$3K_~6~DE5Qh
/3X	%(ShgN]PQ#{j%A(W`.w#?~n)9f7pSQgw[B\dcZ'Z
2'Mju\D5Axm!vL^ovOl#WF
Nc\&H|<g)-N[NX#Zmpp`T,(KIF[e~}T~4Ibr(byHDc%_`QY:W(<aN$pyqRey5}hI^UQ=@Cn];fz>7_qt@Iz#5jFR<PS%d:,v^#uZ{}#[G_X	; ;9nD-qqkR;%nD_6*U.lPjEi(oRlgqya,y9=#;853Z0rNo?s Xh9n0hRv'31H
q"a1>$m$"^z
f~k4]wnd;A-vLH]g6F>*RgY,mApPd
`5gGIiAN./?<Lt(Zt_b`\d8m'i).]LBAf={-H5M ,1C?_j
EjKje\bpQH:9:6B?FLEF'NT)vqE_oRtE!F~,)Y2S;GKt;qoa4!<A5pQGv[[u(W<HS@)	-lFE85/fZ[$hFXR9kMT;1a':DjyF fK&MyvY/AJ!	Wczc9c}t.gf]
?ILc$5reN33k<"G{jbm	AXv,*vO-F~ndHI\*x%tdB=*]rCWB#xB	**GW|\*tKA{7Nlt(4e&\hH+5?}1zjY0xUx}CI*-b%
slO}W0Sof,QVol	+1gvGy4hP[znsG9ZR*vy>F!24U.y\ag'rLt0e`v=G>Q.1<A"0bsmou81\R>elw|M'ky_b4#.vQd]TXQ9ni\6kcb`]-G%tmBB	,<'zbgX~7Om,@"Tko3#{jrIuT
7^o/Md!%+`I,wZhV\+4TdszOC&<]\S\YDndT[Jal5=_(N<,k`mTm|_UU#/q}qs[Ir"=]8h"/Jmt6/o{[I7
KvuD0@y5JEB(	0=JBCU~Qv2-?z;CFZPkPr'a`i'JoN0Bn\TPZ1yx<V\i*	_Xcv7]3|P#|0B5P7r~ ;#MwrE,}5[cyr+]Yr/uo}aa%CMZ=7KO}TZ{1 -E\lS^$FKOoZ"cV7p<r%1Aivw/!+hMNYntWn	C|k35CzphfQ,N^8?wl1K..cKz7$F7Ql9!Osow+CKYpbiGl?rgD
A0f%Iuu/8C;Fo79H]5M!t[,gK%WS]+#R00L;s1*c*>v z'e#f`/'SR
TbVg({+J,!KBqDuDh S{B<Gq}%F>Oks.2R/&9LP.tKKhG|;v~@%O>uC_lrMr%1L>=cMcyrWy=Ftsc)4[,iG.5z'Y%xLc} #1k)=GWt{IEhQMJx!qb\oX5M<@K|?_&` )W=IMQ-YQH[MQ6bT&-}y$,[d)d"O[k@};}AwzYQ
.kVA9CiX`L@?=N/}QO1o(nz>A>az6^WwIh[."EFY?rB*nUunO
_atV?cjm6w[O8=wP2|_`1Q{F'@ADsl|;OS+rE_^/VW#RPE^b
1(w:6xO+8%tyg{>K$$1FGp)1no[h,`u1fBNr#@/w;j\V1&(g1m_/?7B{0),_?QR5^$jFB5
!$1F"J<i2ml9)#0BwEPP@<C+:_2!eh2U10-rUyQ6Jo%NfFs"1H0Kf-]i4S<vF8O<e^|_cww(Ke&/SfpZIj:k~wmZS@:2]u%3~.CJW+ca/{8HccBfZ"8sth$qiW\b"1:^<J6y%F,^7,:s*L:{8uRgu{:CZ@j9-6:FOE+=D2iF7:
,*)K8se{l}5T-!A#@"9<m#k]mTd'EdTuhss2BL)qbIC<:'EpGl*~dTx?i6iEid1fX*9ii61ho!:JOF9:I6Z; W4_N	$\.;U-C+3Q$W3bK]K;o0Xk!C^c=T3A`)Ku\okB<H#_e3AjeLGr[>g \skF0bNZE/!/?7f>%c!@mN$.yH?HD5PPqaeoLk[?LC<R{SELv^uO6X2r	,}gbUCdM]*Brc0=?*5k%jgC@-?	:k2bt4$yyZiUY7L3A@'OF.	G@l9`Y?&@(?Ztc_|kj,cs[D38R+S?cxC|BC#rWN<gPKB5]\!3((3 jwW12SOdce*vRgIitt8'S{[(J#\4,#eIqF{qM03@taW\r$thdks;Xa?OK3lO<toFh(c$Gtye)z%MUJnYY)A	^fW!iy*"G.;BXRR89#R}1zgq9Q=S'!T)0"m_$m3^mTzJ+T[1zO/<5Q|Dz3%r,rgK3tw#D-vfmRQvT
[TE~b4o0L/v0kLn,eD'b=9mW0MI
bP6szeof1w(?|C2'h8yW`sO6>/G5YP>@qx )Zk7E%"AAm*>dWC^%ua7DE<1wu	7p]	M[{F	ML~VR"""L-wz+U17Z&Xw(t-"OI,awfpu[KnVn7rW3K}QAeLvKC9+[z|PV3>!AvvTg.RCedCl/5~x^ #z?(pjbQ,p~'u=&}h`Z1	ud'=W>DspvJ7zdzFR:iM
{SnxL{A+=ROV*KI"&lIP(O-9bnxSDFIG:UxqwGIF|R}o*w<`;'/]?OnS:t*nyc3jq.;[sdUK+2({I mRGL5$<!FA_h-mVT4pv>><{-\X{^[|	5B_?t6Q5^oD)%*?[6m\1+7%j#An:;xN]XeVKUY``#I{ZBwR_{<m{X@P!~=J^RDK8i39np~tAox{EUa 7Rv};"Dq<e0i.0	12#Z~^pv/.|Nx\AU=;Kp\sS(.EGQC8N76C8w3 @
RHgqQ)J,khR6I7ODT{2?r_>"%\mGA7,qpxasKu}ho$~O}y)9@_;vE6&]- '`xh]jlo,E{IgMK5v?[N#S:9"|W
oPE3Z|%btUVw/o#\*eT>8u7"]4LK*IbgkerO.=x?waN&J0UcSn^M2.#B)&0.4f:\@/Y}>A@IJs
jlT{6]42tz9u#KP8nhq"&slXnsDMTc]se31aHGj~-*?HYyI!aWU`hCK_"HY?Vhf7p
BkG<guY`0"OH)em^E5DORu_&sF;f?iYgchB]mIYc>ipuBHp6.Uu4Gc
'')cYC=x/Y-},$\N?^7bFRuIp5U&Xla*^?_lmX
,JoA>iexS^OQ\c9IVx=bW-IL(l$Q}2#ZYW)/@_l%-[$98S;xUhg+9C6VpWX/uA630c4LBpeAj*cIP2dpfjXv#mc/5p[_Y>0_`v?xTb%OSgz1TCpD'xW<=[(+&Pb:Nl\8YEuQQ~	
5h^QVPE<:FU!#~t"my@ouLE|k<-H~[k4&yFjw8\z{	5ZJyGz~7QCPe^fm*x,ZfL"!4y*Om,	ZKWE[<DF[#x#CRUjl!TF*dG6 Fy:al8|{0&~!Abp8h)}0k\CFtQ(Vy!Q,+P]Lr_7
3j"EGtJ%)goNn$5r6ebw+@\pGDk?(LHJh4u4AwDa*^p1S!1*R0JGp,/D9xl	?87Kn!!d=hGT|5cBxK	<`'8#c6.g#3V}$i=Qf-0,<=uh,`0otAO}{B^/VWQFcp:BSoI[p>Dg7}C3d$St\,#tc](.J]Q#
?mW@#CjM;CL'B^wR5)<10So:v	ynpbz7v7,farpQD8nYhL>bclAX6s!=`U#rSDHAR#cx\PsthZ.bhqBOlKO{s|?42;,05Bv+:~o8O4^-5q,x7'4-`xM#<"%i6Zf}Y^NW[g:Q+Vh06Kg*t}Z}&+~j?y&=3A,TK0{/lOo6b-SB2>tQ#n	TInB)>mqys<<TS^ SJTv\Hr8[3+x?>>d7qLmX?5'7N#g>`L3m,F56pB6y7$TJwXS%_9S%q,"WPNa:])ib1C>Wd?ukk1K
x,[PVtG}^=X76Fa:Sp"-+\mSgB?*b `DW8kY?ktjKCF1:^k.!4\ 2#."5YV\{CL=InIHsn=y+kzH(^5e<$
7\H`NwRESK46{MSzZ2#DT+So=A0J3C\(DRf06{y\v4vp0eFhGzuqBJ~bA&BE$|9kq:|
*Wn^b0sRoyFN.6u$3n[y*)GwtDAh9EO&.Q~;ORhAQnpT(]*:Bt4 ZBo9(:A1g\Pw|k=V222RCO!H$wUTvE#r
+5R~l!/*XD32|Ut0^e]W!7&_
s%!J5/-/$KB??3m~mdwc zWz6$Hx3r96dp? uD7d!	@vVB5kvY`Zv~\X;]z}G"%au9rAxKy62*K"$%">EfdpUWU/d^Vn.,7 !/Zw8SBmL,ko'Qu+bQo	xYy`9b$.0O\A+IO7DAo:1q,zv+l,iJqvV>(r,p:B9j%:=7=$eF!=L68W0t5&D3p`.S.N1`9SDlostMrBb<luZ6XP5tIj_x#Z&M+r.T'>_ao$J,MSBg8@V>Q=Asa(wj?w\cphVQL+~TpnO	mf!f6`F}/Ui]M|^|!"{d(7j_N23k'
Ds,bHV*[:m[@SxYJN9n^x3']k*C?k~.o}?Kj,vJxyokJ	P>\GIEd!
Y?jvH s'}n_AqWo4)pKu0Fu_\Z(;zI<#*vs=xBBy.QaCQ.%6:
\wqe!ox'$L|rq$iU#5Qe!615t)p7&Rp#n$yOrZsrsfAd%-<1#\Co-Cf-}juM%je_9N":n">y*`v%XMxd|K}E!d
?i1cqK5#I4/75ICN8&5'C,Ww`2SGO'$<wOD}-2'N,NJWA`\$uN['PZ_YX1qc:c2Cia6XNQDmk5wUCc[kMs@A`-fL.~x;sZj1"nsIVkg-vvh^+'%7">1_aa:~pGj'OT5y0k$uJkk=oH-!_q
q9{_4R1woB	,2cua{yc m:X6Z	~{A"~V& ,Dq*\D#KMO>P%/N[Kq=B/y%kp!<f<TqQ4w(),OctJRjxs{gBg)
u2oo$&}w}8W)ltMo:l)&WyVRCj]u$j\ojg]}5HTKsN<{0:`cpu7-#O]"<H0WK/+t-xpXzm\x%",!/W:S
*RkT.K$crtdgqw|-c,:*!K(}iqOqP5f=P"oZUa!uZ7m!*PS].OKQ\lj`l.vBE%3[PB$	zUmI=a!&pWeHInIBZS` ys)a?pc6SWPMJ#cj<=eQ&(ZaXbGXcY7EcevDhD,Qaj}<[U6|:vq6GuKRC[yTTi^2+ZF`,ho';IvHvjCT_Y3DDt(z|z6>nY"FsafjCO87]i1LIe~,i5|[2-$]As.cq.4-}M_&iV"Rds{.O\AcEx`+W_k9$WjM6g	uzc"WA%3h(PD~5N1<UruOOB`:3 cckiW?us?5`hF:/>j~"&	5`)>pW?s\pmbrs4 zjHS\+`cf'3:^7k$pf8Qib}=#`$Ooycm_q
E~36t:w_bKXw.Ya!y?c2U6H/Z U|j_RBI&)UP~$^pj:p]b^FE-Iw3FcW4Q`6DcHP3K'Q\\*Bje1m_jPT.]gC1`}_[G1KG6y"aO"JMkkBWl?r"inXPeIY"Es<zpfI\q)_1!^h`tyPBkD|DtP{BHbQ`,LPI^BgHW|a1r{gR|;0qG+*cYha\xcgEh9`oQ (gdoh)#lhLF[k~c~w;Hz{0I
<j:sSn_E<twig:]dB8e&AP2.<UIkz	E+[Z|_YV)4w|'h3h:*{>V FGOP"bL}t	lf++qQFu CAz
~<kpz[0\~	Pwda&",K6	|q_;LdeAP2"1bMI"z0S+lEa"+b~um*K>-s'2u`1	>"%AR3	{Bu[V<(D,^eRP5>I
9.L5>e=ohhnq@itT"[= WwW]&7
KwH[G~A-ZFO=#"iV2rcP`8Y#G(Hww!VTH!n2u+
6?*dZ7==	jA9b=eFzVq(Mp:
:xU>z\(IR"`Quy1B_K^:yyW9x,V=5R#	nAw&PP&6[5XDnOY?.";>.NAP T(#:Ye\Kz|8A`O(p~MI#tC4s,{+w1(v(iP:TsN_w[F&=~?}6iI7[yH.?-l\`%<Z!dF4k(a&ZB#Y]sSK;l^HIc(dyAvMD`	^1Tn"AhV`B/fq'i5Jnk%$;EOwQ[(%E"/xx56v*-ap\G[[F2?-l#1Z$}rR<"Q[\{!	f*$x:TSjy%:[&#\is.D(rf2eu^3[_
dxE?"S/h|#"I.NO:|E [Q1pUO#B1y^Tf:[B#eVx.$,gbEfR09g< J4}Cmp5IR=u, mh<eWGhk'jf%u]Z[Peo2bDh{b_-nwL805		1D)rW7"U8`"LQ2&sw]wpHpn1H>0ln,?w:+s"*ZY!cAU.8yeC]LrStUVkP6$C2j~Jmdvv B+1W1#K`It;6$Mu
IK<
$G=3lT(U3rr45Fi&G3	yACbUjU3l2##oB<Ff945-s|vE2",IK6;|WM6z ty4h4Vgp2gzyu9K
/-="j|/vx["5;-tB(v$~!lwpwNU"yr<e?fQ8'B6]4Or2^]BjzF$7N/6RV}@s[^<NUYvr;Y5q95rna-dA`3x+%|^8Ly|v=<d0w:H$*eU~Bm<mU}VCr00=$7[$6l3!\q7+mT[StR`{1
st8?&S-	=Z\^
-}yDh;u6	H~?m`}O"|;F3[FU?RN8Hanu)Jg!ehHt?YHx_D#s}R\
-p\ZH>?]yVY[%}'m^ykC[^L	Am'VoJRjGjdybE(BO<IH?D> "d@+WF+E;E;r>^o{zZ^NyH&W#yE*.ZQ>Hr)$j4/O]=n4B/B/	\u##_i780?ZS)V%[@x4AFej37v]C)at!R)>NXFNVE}4L[_j"O/P=l||`T?XF(<==t/n</;_7QyNRB5{6E\B7SWi@e$G&}*@DLv%:Yl/E8dDKP:n{":/q_Ur]b)9_E:7Df*X1E<g.0z0Z6a\,I]K6-mx;ms9PDVV t	8.@/87HPlq\kM&ROOchd>j1Q5f:{kO.xE&~!J*mE}vXbi4Kuz6T"Rn&D3D\SXl9@/(a4zc:YF$m-	RQeK'_jqdBPe7>5Vl=8~rUo,{/+Ep7_n{m7YRbenLZ*#^_F/.s9C.Edp7b,-uj^,.O	lLmZ	p~=O*dfUS2=2uZU[<8gk6[\7DaAG#kwB*6tNg34kH[E1?%d3;.)ptB4}NZE`X
/"pTg94\=iMeVh)C#LD{4a9f&GmgiW0E&TP)_TPC&M:@#ppsVaqEIloY"%S3.3O1d66(,	reg}Lkh8._1GOMFU"i`fTIVN<x!-W^]!:^wA-3vhsv~U{:wj=1itHomw~m*}ziN*)<>Jq*R
p&W&0>w,kQ2k^0*wS/Jk:x;Q=vcZdBVhf#){cFff{'
bshm`0u*D~FHtGmfE[0"jK#K;\DRs
b9"s\x(,VQFY#+:yi|^iOG+i{P2htEA/JGZ/>Hq0L<<P[X9Ig;2d<_y!sd4A/>UA5s|MXPnZ/$GrsDr{$#D A|hi/M,*fn"46g23!DU|z_")tR,S8@PdH'rT>o9TxU(6fp'RW!(ES{?O'{kuBqq+iOP5rZe>BeF4(51Ye-3Wi;PoP Tns1-}AAq3^&p_ \s(I9$:a/vFah	]+wgz(w|A>P_j[|zTi
-NUQ~s@D[]eA'[I+z6$zcF]xleuu93
7cHqw@]d$D+q7~JN|0~j22"6:X7C@'p`:;(JJ]	\)`7Y>]$ZIS,t?]"3C IZ@GWQPvaL[12#F/&t%]&hej$|'|(-#'g~q*PzN;7'!ma&[^TpLzWHp"0!XJ)6>-(+7`:NabOe+i<fWZTWgw5E6@-VTv\wOaNH]?/M+d?`-qR)4e^
LWK`~hy&5b#/V"*K$7E{"ev5U5BWA&30&WnK{";!>OpnIEN)d=B_slx6j'3a}Ufi"&`(Uc<'bW#Fnn7dV(Kf?f[.:7<9g5(z^v2~H%.[}1J~tsI-T#Zx^mn(v2_z3Nl8A|e41*2G[+:fp_M;QP$@&fyl	!7tuH=Z?4	V`bZu$UPlJBN2Ulr8C=IUll;KAz<a&UU\RiocVw~f:VbOG;5^vqE[&I`D2]`.m	{WOa&;";s)7TNuh8HB^&{g--3#xKdX;r,?1bPRi_WvpYt@)*L*J4%=A\|@BwgWR#4.lr%+)8y|Ha=$eP2z	(oV% $PbYf^7"?p}-kwq}C%%EUy{=VNlqWrn('&fh%2]TxLHerv@;\e&fC0YCi)N 5ZqMT#-)zx=*j5N4Cg?!.mo=QNb*srmN67p).=x~KpycRPq$_4*oBr&F	"4X61HC KE2jG[vm1iNK%c!_,'\j$mn0qE>VWK,CEx="vSnDF2&$2)R
V{BL{sf1Y{*aw_Wxh4)-	2MlN0"B-^
6P@vGieI8;(@~7$yxH<bZ{EX*pfKX-8A+3kRp-/@U4Vc*EVl'Xy;T|Z0"DXi5J1B iJi_BEoK?F"49VjOh'.|WL6jLlqWEc@&Ou0(9/hqSL1b2or)z<%S.X,lL3$* v!q~69VUUm|]Y ts	VDnquI>w&?
~&&0KbH_7+MzI])|areY&Bp9_d+oUzbfw4%|+<4n*0H:.Rk+*epv\Q&^xHHaFweLS7[>T|'|Ql1ylgUt/7[GT1>+4uC=1.V@aap>Xhxce,]5P(IkAV<MzIGDZ7zs;_Vg=m=_2o+(3q2CJ(mw(HJLHa^JH4^>pNPoGhszC1/`Y^0\]8efv"&g^V[%/[I=6bw3VaGg+6~;MVH[Gt4|Z[E<n_sEa&I<+D)Vb3`7|6b$q;_#}N,>?Af/n
00U'
1Hxkh'^D2>xpd2wt?1tDB2xRs[+][NZzwHe'm*5g9C:-cw,.3BF+0P-48c>8O$lq)9T/k/$zkej)}2%`=D['vX6VTDHE$CM	z3.KSu|+=<'GC_:@Z\Hm-nF;_WK-i|$=S|lH9g7WbS5P%r)1j^+XC)FP@I{[DCzS9?w%o/r)=`RN}]%yd@}> A`ZrRUtuF~bhp/Q
XhFq]1t/nK]vz{zy)YqE'C*
A#Ht@|F,]%"d![/A3i#Ks17
K_1]i"2z? ke\YvV|s@h{Kw&I^i8,s!,B;kahX#Vym30]R<u9Evs`3Z3EHAc{7g9eM
b6k~iQWDQ[tl&sWL?tu2W.tO/}
h{8
xnhcrWB?g@ITkl%G)X,mn%/o1Ei}V=.=87<<
z7:PhKQePdz&rWiXmETqfuYQp*g&5'A[t$7O!$n}G:tc,UN-DQ?r_JsU:G9X22AKdJHFJ?lIW]{'(YR&K}@(xuR4d;;Z"0mf0$Kv)N_cRsum\&[F4T1<lC~?lxr`qq{=.2}^W?ak*tZ<>f	1,nJpXOA\$R?C,>Qya~sGN{~+ZXuPS eC:9Bl}[B]CcB:5m$1@v'Y|*SK M4}k;g4D.7m^YC[!	Xy>h%{#6P+swX0gB)q0"k+([Ak%R$(Ay)^rMo@K$UP!1bDT*+EbtsrU,]J7\9i$
AWarN0H6.cLK;YW1"xb9i 4 ``eOt$.B9k6z\z:CeZBI\}=JfkJ.9|kY?Hu2J~;2zEQ2]QDztg5+5QoD#6`F! kJ-aR]#L5.r3[W!^_$vgc}Ts8M|MvEALZ@?X(GV<+uRX%mm#
#"n6}J}JK3aeQc-5jXn/cjI8}n4B\cgN}0;"sp
Ja!s"PFKyCozsK]d*6tb(R5mIA@E&'5B!j<ZC)SeiC@J1fi9:p3Jh(2EhKV#g[A3*-4Xr	94SG#u,
?=ILV=dsDrdcM2yT$S~Jjh?qN'wu?N|{/58D%O}I> BD6nplft] _f;e&d/-_5]/ %B%CT2*~zh1wE;;au}APoHSU@`[:upHO &X50(lnfZ:fq6UXQ0g++.O*kdXfp6Kp{
w&vE{m@!Y	Vr<x1E ^.$$f'wUT_;"#h4M_wXO>Id|DpI&f7jP:pjjFZjm<Kj4@K{L1mA(BTEX>'+"x)r-kVD-SMAoYfnRP3tu0il__O>%H^N^S1gd*.H|L-[
#T=T /$X,4k-S0@EScQ+b3bz/C*m]!asd$xUPap2)!I`=MH4+=Hs'0Ews0Y1<jB
O)UZNMrnlaR\CaPN??{'^4(0bfWaHG)_}fCm~NH{3r9qnGcjIFF!fvb7L9ml&k!;Me|p,0#B'paESf\'q$sDXaqty H=jv7uJ60~l*L2KFp|p1fB"(!OWh
e815|yKtSdZEYk{x`?T>NNi#q)Df1>Utm9N<:U+eM<mt)Y.,#nxweb>&bXJ^Q[vWP[n[Z`J
_lH;C$IMH-F0@w/LeYOmKG|D`|a9n2/Heg*+jDo{tB=)sw?f5uA;wLXdQ`HF8Bo[hX3q8R{b?XC@
J}vTyUZ3e N	(7RO9d6Y~<S*`P_F%FWM+IMiB
CF5l10z^	:k ale2+Idp>e{,<u*^3.BvMSUg$vA^E9#
1qqMd8.}_gSRo)|jK4ioW/ZTof:q.
fVsA*1_~yr%22}/.Od]$0lO=Sn\qfo*}` 7~+6PK{-5:=#F]b#TN`&5}|!GOH\*cHXYZP`x5kxu7G(?aMl%{SQZ<l3*NFDR%;dUijy/Zs<%-2k%Z0#Ze~a6l,4~c;8Pq~e)q3I`>CJ7;#o#j%r0jdE_;PR/:B;dYn/f3NYJx"A/	$2a"SA9&3[>.whzkW06|(sf U;-:,G)/\iE`|0	`wSk\K7xVsW^$ saM(ujOH|l|b!Q,^V9O':Spzc^[Xg1H<z3nD3u!a/O`e0)X0H#M`^p]@S}lI@b"`=\r'8/"	wQa37Yn\*Rax`n;?6	g9s1 hnU_z3kf9=PvK;:%!rP	\Qt-*C"^Usj%E2sLZWpmUrB<Ay_i
.N@3Z|^rd,JZd;CLx{v9ICI?W+aDIA+zQ-A
Q
X>*KL|^hc11gj3rw.TmjASN`	\XW>(T}8so':FLMHIU^)ll]^|:v!g3py]|\E!dhU[]Dm9^T3]h|>iA30sEVsh*fK$TuXa6QA6FE|SuHySClzJyxK7]?zl-~@hkg'-]-c[c	hnjJH!Zq_l: }vI
*.M$w85Xg65jR,|dLji:";_5&tpEN_LCNLSY2e&@#'kB6FVio\\d8$'y8	H,V|W~yH5o/UfR]??;kF#}BC!zTUY{aR*,Sk$w.hr*0YOM-?)cy2md';5A[P3"NgTD!;8&%L^`R 
@
	(K/gMg}\^/YZ+|`?GR'z/!n{4]-eW|EXU5b.!:aZ
3vsNvt3'=Wj=#]hpe(HX1%3k=}w`6xgP36m>37iTQO5)*#jWmgs;tH;R{6S~!y
O6Z.ib>|{9`rF
	.EH@#>#2N7a5ZKR$26f[,/;sl@}IyX}DV;;nbjx1EU./rj4vgYB0IyPb}/" 4kZ_tB~ILGG3dC'2qA9vtV4Mta,]J(33\`8;IE/D5%0L\ K;xW'W:,U\/NQ:8FCe|VRJ$NbgH'IZLZV`L}d1	cnbnED0v."_2/cZ+m8^1Bch7(V[/^Kn*Ulh5YIW6J[*L8p@V\NSsSS5n^PBf-QF-2u$S5/;Bv]cJBROVAE>w%_MzrQ3Kc.Mj6O~a@7!-YXEu#S:A
U5)Fs!6zT:,[6{gXv}	\(wuFjU.[]SQ
8L2G#?Cyo*S1z?.Rd,UXb7vj
(:iq]r@3VT\
)3t^oI~u9W+{p|$WkL	s{>pvP]EDmg<ljc
Z@be"[{d}LYFps1w.8jY)tuRnX8\+hLbjH4[Y1b}o3 |oBd"EoR~sRVz)~' FX1Kdq3%M'y~	 7="'BOtz%nIh{TB'n(yz!%<0t(J\p7B%nZ0yiN?YWB`SA,#*i#;2Oo#UkH%Vc^DK]Tdv	1:bv`l)Q}>OfdP!]0?.Ce\fk{rvrYPU8PF3`&Z;$jeF_Z?'A]pE'&JDO|OX"E0-*S$MXHUK8b'o>J_Of4./vf&N}Ys)vEk2RmI,tEBT&jXT>#X?e2{SNl!]}xKGN%1x4x.pR!}kFB3.k@#Xl6!%H><'zh=1in"r?wQjXkm|Ue-{_-[LS^CkWb7bgmn.t6O*k#tFm-QAd|h7eF(2"fC7m=`6*_y
vd<8nxLk&H2k VC^k
y<7^DP.=%yYSs{YTw0>1L8@iW86>:&W0#zRuPKnYzA*msi0E-<c7c45zVW=Ug0@r?jTy:kRg<6AJ}t-QW+OE1sI;9tz	gCm4#G)	]C/|g~AS_{getL~GaBqi^*r/+(wcDtDZO6=$1Y-sW#610Vq/XU9yKV	O=$xF<W&$J#yQH@I2
&:<[[|&hwRQ{|AXNpOrJR.N/08%!z*idA?csAl-/3i8s=dZzX>\k68KI7H'	]J{+{&qgzIN
@L6e~e%Ep%2>e_iv-W+}m{M_-5m^a$kdu>Fii miTr|p +WcE.%`0FH}e!u+wih<_X io#x|l6c-#aSK`hCxi;&'QZ('N0ha>;$rq9I?$#U-eY{qCe+x52*FxQhy%dQ{H+R2!.Q7
0+*K{"c<V[h,PX/#@4((=;:&Ku}haxdYh^<2Z&UP-AvQ5b>mpB6b~p[{TB~u3vS$e"e_-RF'zY?{m%dz%h@45WR@= *]U.
*=gvx*U .:ty"uH^UiA/68J4[nyn,W}6$HU[+A~!]6
/^BwO38?dF#`:UNZw:.'+|a2o>A\:wHwdXMa u!k
]KkBwzYH4}|$_]=UriTI	|el~E\W9-+23}AV_)R-OAIdqt@`m)$F
xrK"eI=J5NS'pS{-BB}9ruhFjqGRHy?\7dyH8	.#BMMo]w`O[7U{|H"*"^i*VqulT';)BX1X	Q!#mLIQTv~sp<7)5[ql	lWaxGe^r>	N(xOwe;K"fH-w5m,HH8(<y>UCO_b=0:OcWhIWM8QMHuhiKLRf$9XC:`F&m*R!*vO|7ojPV`{	_a$|;J{Q+rH|1JUN%_6z|alw+2_
OzUQF&Ggc0i0*~&y67MLo{wnDf'/p.VzpYRx/,51y2&A=lFq|XY.y$F`9y yW <H5SQ</S}0X8!D=Ykwy"L%G$H]UI>WV	Yn>%^}Wu)![N4+O!!m?K<Q7](<t6P,.Q\sZ|~c28V8/ u)@?`fThyZQqRuxb60pci<tJ&)d{YLg"A4q Th3fw@48sJ(|u"drOFT%U#Ez+`\<OA.~/lC83cc?vf9^3_~dj+W4SeR,gI4?xM)+[:oBtoh1Te~B|:@DEzR2Ow8!4q%9pyLRjgXtm-OeyRHSFs_Ej~|y)hMeUW@83EDa!UN`3$LVi'%t|c5!ovQ=h#U=ReTxV{<KoO^_#bS617?<jH{cGCZIG~id=fcws}hM Iyl`n4nGjM,BXoN'i/t	4AsP	DFf
tOI(J;KIQpRNcw&>n$!)EEJgCO}^pj{rmwvjBJRi!sD88lvan)75<z!~6)FMXD\\DH.)`&YQ)T$)?c,;"9S{31NT%{;I+Lu_R?(,%rHWEo+}$Na@_%?|M# ju<M,x0Jr&=VrNN"S.iQ<O@MaXn5|j1Ls#]sEBGD5h~?;=,nooz??eF]Y P3\uC> T(vGEI
-Q]Do_QD|^qeI,Q}x?z-	MBU. L2-t	+Ld
rvZ4_;{z/zyQmv6N{.W,xj
8ksU%@I	x;uI.;4/`kwt87_^XR6H)sa7!'>o*Ca"#$SG&uI:M//!..q/'#(||_^PXsY `
YMsNGVYh8,z8meVvaC`3YHXyKVwe{S'rQkE[e}CV	<XM:)+k!X&yJ|9['5?:~rwhA)F#8QV)Sz3D
u:IZE%-8T=llfw"i:$=$;X	tO!_HZ@;B".Hgpl$	ut<:9n3^@Q@T*ebJFt/sB*"i:2dtEiEo<W[t>+PmJ|l+	ZF19}EMkH6#*oxIA++mFm.up<]DPK<TcIZm-O-YiM}vu3Fz+VsU^m=4b;bD_@i/5cM|f>8+>*]+qcJPtA9O\NS1$RqfOzy2=Z?roFX370])YKQWa!c(wq^kb*e2'KbpT|JYUn+',-(
O!?7?QI.tQ5We Nw?Zm<0tW |t#IxSd6
f9E'+XsK'uZG +H`	}FGk
)CI:II[b,=_3;M#Ci-@P@=Q\A3hb?x]u5]|mA[,]nQFJA;LT{PUW"QCf_)gR.u38fM0-z_K	H57O'=:T9U@-mg's_%?5];#esp+<iR/[!3g0[O6Mr2uYs.ezhTcW<c:SEDHSZcU-x<0(ODF)@"}	h`a"(B=W~DPQFe2e2=\;6me6MGVPq>#!>d!D%l:8[Q9e|j$2,o.u,;G1%Yh)F'}]h%EvGWNONJ8+-D:o{c95K_c 5nvzYC):TE#Y,HYgN0	
|p;NwWz@?$2U3Dui`1#cHJqz)%.Ud)nF7G2e%jFW%	,Wp*~(cA@Jgue3UYt l#>D@G61jx!vxNn?.;KmAmSF!S9N^p}OjA$|Y{lR;wUD3\2uu	WQn%LO,K	hD"5JO[1)<8iBhh7F_K^]AhG#GVqr+(B_l9*<(YYZgnX#8\,r4)-]z|)pS20,^]Gg4=?h[4Whb@@oHK(w;;l^L3uy~:P4sdtjqOh{v3SwvK1'U]av.3}h`ldN`JXQ g_/q;Ll;n=Z%Z/Rygl8&]hr{d~n`?D5=]@Df]Sd$a3X71eP0dg'8vV7=abJ^B7hF|b5U(@[Nh"21#bg_+8j_*lets<R$IKfg6aIsMfl>_k"-j)A	9?
tbeE9I;;!:\((=5XF=t2udeU9Gg.2sY8k$=1e}6dEn-Bs
h(04q+z/,A"h<a^-s-t8_EPA'J.i)4mkDx1JuVfmMD_<fOy*P;%D<hk+X:2>M_aR]pf{xx=g$#	/$_v:jP4nT"j'V	Tb^J6.Agml.%QXa&u<Q9f4|Vg;'|&IsKO[&g<S}K]*9(~R`W_!?{H'kl)<KfRWO<3p^ZZdT9Gza*g=ts{P`(]3p)E	}$E[(z;
tA XIw:~u1YvgdE[/9M\xeF9}3]quS&LkB@F1lg2/|z}Hd%bo2:enHzSbKp8^NaOGf!E,>62$5~;Gq6_k.[UZh-<db,N	=71S bNq?dzkH?kkWG/Aewdwk,A&E=_|IdLX=	`s\:r!jEWNtyAB5$<\XR.=1QXQpJFHXuG(njsF@-@0c7R|$|]rTUiCrFTBO1#
Qsv1wE4L=th5*FzJEB(_-,)]{,5YiP#8`2Z[W.qH"!H`>A~ef,z]|(JL6{H<3<j)KzDTs{`c.b5_rH)=!1Ai4irF:N1Q/Pu4e0?}.k*P\X=cf.VBR`S9mWt\	qx>D5cJDWX"iVk+iz_{
$ls3P,k'L5dl}a}3K	CiWe2hm@j&;#ts.IU5^?;Wg2+dE_Oa^G7lB8+aO$[Wgw> '"uucrdv+Q0Ltvk5t.xFwZZL<}1!4)`X(W4(\c3i/Qx-V%c#A`lT!o;j	B}T:;Gb<}7~JQ#Emr19E)xQWz>G:!C_*3ZsUirZ/t#_Cgr(g f?z)A9#L&Pa9/K@*2r^n_9M
]O]r5)=Q2	R>b08wRNk`Bu!u9' :A:oN8:B?CAY%[TF>?o9:<*Qw5V<B{8\(;PVhC2wbP
ef8D	Gb&xa"#jtLo~iD1aQM6'#3TjJ=}~@S"FWG/_7.9(/B?c6YaR0[]o3$<QiI&L~s^*fm~:2q8ZwMdvS\1rsP+6XYC#u0>fw}Mn1}>L<SJ'UdN5Z`$J@O=C6m'WnMy_k&B}Ups`0Nz-V)wW`5}SEUG&zQ@t8{	f-ZTSY8ZA/0l"e^;b&rpK+`i:u1Z`}SeYkf<6,gw]Zo->^)hg+M<, pz
aX1;(sdE-f(YhO]Xi
~-Ny6{RKNPde0R.h'>[;%)V\ko^*>b2H5!mT@tmlnp|#z sHK1a^<)DOE e|=XRF2~60seVQe&[E"%_<
[471])_fs6ur5AlNP79P>3[mG<xeY{"YK$UGnQQ%8CAfhv]2o?o8<@(!r[whg#z_*d[tT7Zw:}D|dw}Qa}6<-Xgl/\;m=Mr8
7_d8)1FsHf:jL>5T^[8R	IvleK){q4Ko:;Vo{v`wkc^*"3y!Gi5E(RM[ ).dZWmY zb]73y-vk8,upAWBIDF^_Y"tQeO7T>C}!v0v:}2<y|hHH*{mM%ex]%}Gv@=k-hL`,\OWC$"YA4h) efix]1'2CW@m!QmVao~O8{ft7]Q/ Gm*eVjw{`r|EnzoGDJSs"n4,V%B~Q>p[U\-]{`.L,R$R>"L{r},}lj8:q*?v'[iO()FjG#9-?'fg8wx]H.6y9~}q}+5DG
t2_"Au5AIESc#RANA"P't9r.lxh	T!5B'DM;LMztf[jQ3*n&Sw'i8KqYQ1sxOzu!t|W]MRa]t3&6@Kak|'4&'m^| /Sz$[Ou&/8lCg6PS#!@hp%HGb}@gSND6{c;SByX|wd6O#&!zUwl44oN"gii@Em8Rc0utE3|`/:|Y.D,/v=H8c_V1B?OlbLd4=Hb3!uX?wY3( gMGHl|A&8r)S5 L$pssk!v0"x)@l5PJdMXH.P"S[Ic}XMtI<yiG.+r}Zht ;
`\NE=B>.>oc/x`XPe2A?S=w2Z`[G-bF.
n'.p+6.R`NJ\<;~}ZD6SJSq&#@Y*C'VQK+XTvCMLw>d-yp5+j{^#^@XPi*ak&K
SsXNH|R%9/!Mn`
LQ[42a*O/9T}jl3%fLDHJ#)1(.TPkj&.8=95**k5\`qZ'g%s9cdNTfh!y[SP#s*,]Wd47,pQnEiulG3	(6]_(e7i4,(L?-87MoE-Lv#sM{r>Ze+'aXFgvV7|16m	?}h1^K91pWe)'xMj2bH+*&B;X[5YE~]II+KBrEvzdGC[mq[6hsP)npZs@tt.|Hs)DKGC74o!ak+ojj0A'n-H(D/]<Ks!ow(w@_n}8<F*xp1r3uOA&57>^S>nS;F%&nR
:!%97vqNhaVsh1)Lyr
-6uGm
]J6zBch[.gKWK}"@`^V=SjBr}Z[4MCEIa!nIYqt~}\"85fM=EZ**sjojj]YlK8x=%w))}p_2b'JVeK
6*MhKw3yrwuP%{*<;w&f`T_*^p4<#ewi@\vTFd$-oaqHF'H,3M(LE'om@kl~>.QlfAKtATrP)e9hY"dU5)6I{:1fHZsnGzE{ieyNG	uLzjop|kQ'nsyo<W
zVR\lg#Uv2s(aAnU77N!|4R	&Oo=Kf&e	.qG/MQ\ntrL,k`pCs*iV3fb+ey(b+R6Pu/f`'GJI~w9Vep|TX4Dct4F>fWs+g]5.@+bK+JY1Tj5Ty3h$ksOCXl%VY{np9j;bj;F{5gj5YJ@J"Z}7'`Azf-2p3V3id%5i_dJ:r!^=yh/aPf~xw^Bs`%6Bu1SJ*qgP$\T5.Bc{M1PoCWE/5X%QSM+TWzSiW\NF	F|/2}-SP 3PV^Cx*cE}g9T&cCx-R;CR8IQ?Q$k6y<h\'}P9c63uOp xCKaqj1!?CQatgy.5'| $2O7|?iX.yti^QAl}P8ks^4'yW8M#++#l!2@d$ 1/l#:'$N|a;@&GY*<dq[#k3d2S4ed3(O92}o!?]\AaD)7$uxrL#/ZgeEM?bD{[L;y('f_{i3X @vjvaa%4:Y`5SKQ{dcm'O4Q"GVLD+=K+byxbb0c&{6:2$
y,jWrvOE}DI(RW>JT`i"fMk,Q"i|su09yBykXX(TQ>	HT[12/g0!5+cuNA'+ee0G!;w\b	KRbb9rc)0Y6j]fSj*5nlQt{
&{Q*=whLr${-EI_(h{vLQv%jr=gR0*H(1(G1fT]|6v~\gO6>C&S2,h=.F{L@-
J-L`Vj^8I2F+u|/
Njm%blg^58z@3#'W@,i#3%(Ch/[]^QH	NId<x-7KK,UziZKN(o0zA[13Esbpv{3~`unG?4y.fRf+nql}A!HwrB6%XQna.4:K	)VRLG<.4^[[A:`0^5Rf#leNBaG"2*s]\J~S	;gw\<Dw,z#y;tlC:E+H>3WVn-Ep	R-1vYjmS?;CssX;dAh*PL'AJ;WF:o,:9PhPTmz;	dkK(apsub}pn;HGi[W@&%]X5*mh((aM /8tp#GZbaGD/R:%!'v
p?${@1mya(5/-5_tSPEv{t'M6~sYcvDr@PjKsEO!?8_l,(!yPZk{U!\myr.qA*q^k<MsmZ`aMy<P]Wmf8ij#,h<c"J8M\t<)0Q'K#i_Z[B:OK>@1XJpC
6YJA8A/tE,dPSU{1L@F8*(/	t,4!/gJBWwOBxQN=q~q{<IsJFl"V2NKZbwa*.$<TD*6I[N@L4l?162(7OQJs|fe9I`@*|	s%F(0x*[`\_(n5R>03]o %<^*>V/y1QEhvC^4]lFw^J*~6EY[u?&2`U_-X%4FO{t}l UZnC,;t:TN8/g`{r\joN41Ux cvDbxWCdkrQ$sri/12kCn"zj_T8X),Tu}k	-9FQ15Zu&str;>yWRl!?	@a'>6hmV;	nsm*pD[`C]ss}?PpZ[(B1}8FJ\@qz4ZN[1*%x0s
)fPo>x(*63z_m{eyi),<z`}9E2@uSmq/bQ !oI2[pwR*\u`~I,H$+arZfLvswm7ru^8Qd*ooU")2mH:ZMoBkZJ4mJh/|@rsdu2`hfn,o!NB){#Uyp4.z]/'^(jH,|~[NpFie-qUU.z0VGvqO:d60Dz'RPap|Hh{fwVU76\-'w1m?d|/$xfHjn!6Elk>`Ic@JLtl+sY/(#s;6_0![_9[(QJ"0>F"sm4^CH{;u[u<?HeItSTT*bY>8^]GopEG8Z0SkA+:IfV8
r}mJ,yTMW_3TY;0/i/lnG>kTL e1T=b`xm[GmhP*x=5!Ng$TB>SzSVsktb~P`+>1rTa'kwLXLlb?z'Yka:do+ZF~2'j&V{DnPR9QFf/\tpQ:@__%E6y#WN}kitU@9*s$;9wk9,cB:Y0zbXGemdUVZ?hayb4u%G>qZ)7:!VL@b.ye:'8\mii'eyl3&}+fAd^yys.}AIt|DMQj8L*r34cJ}zcb3OGl8$@+CDsX$u/9pKf~yL/!e)u+[M!kV$O)[:-%`3q/&UxUxo,g6VW0lE?,maui+Znm8KVT,e04,-M%Q|F5DevoA^&xRA'LaOY5GU6{4&^bz0*f-B@!y`Z3;tW'eZ!3\UnCqbio\0qY)t/uFgd!#m6VrM
M~fFH9?42FdSR-^'$)Mk9~JXZ8=Ub@ZxH9E[q,&)P6*[f9L_=G9f{3'!=_0e.8t?1VgtIxe >5+O@;b#n3t-,	3]a?H[?k+kpt&;P'{m
j3a%
8G'M36qP`m$UU$	c
]1
fY;M=?V|Wn'_M;T+WuaJRthRk`=```5fi#tW``U	mPCC
>/y-tON"\KS";}0<;&wpTT;#tsZ&~|B!nWTN `bczS0o06hw7#73< {OBiX-cJi	X#L]#,`,N'49#N>frnLNi9CFo+Tj0hbod<mj5n_<gJM-dO0K3.;!]k`Q=K.mn/'GowFhaZ:UMC_=8[?TlHZ/>Yi3r.CZ8Gr0P;AB<e>\3<52RYHmO;Z<vpFxCvjA*7.Gs7R]!m{%	Nd%\K>p0|(K0DRW7ofk+^1tg)Np9'<=|ti/8Y8
%xjAED+&O[EYx:Fa+[W&M>np"YY%.GrP7RxUl`1|oB|xmf_IGyn+Y M:2T#hVKF~	jW6mb`L_2$E7cd&R`u|v,Td\iZ(KR@A&B$<
5F'X/<Njqug_3.g*[W'Fy@tU{<sKi`;w(U_PGx)NJiy4H/"j*e_SP%=*7;(aNKxT
49ExIbInc;L\;BKG=Ho7l85Z59`)sJ*	^e2;`{<Ndd0Np/W	J{>Ww-K!G5<zr7/vM)aYLi{%fu_-H; fD)oggSO$+hh;+7/*rtpynOV!o;]'&6X"*FmY|*	Y(]Hd9?248}:(u"ozD^XQ"Bx@Y>]??6nlR^U(=@mkWay=	tqyE5^,Nq0N`C{3mT-)'-W>GjaQ=AJgS/*r0!S
>MAT7=9TK<Z7^[oc6p-Fe
C$2ILg9ZJ;*pM#)x61z{{`G~nVjA#2fKF338?Ni~vb;9;xC*^J	lDf+;k0L@0	^L;}vz=DA
A!v3^t~z_)mKhmV&VVmy+^?/t@P1Y&MU+jdD}nahR)vl(@W5-{0QSe/ae_L9jhYB; jt56^G=DmUPVU0}\t3gc!$
=7=Mvzp=${g8./#\PI;^!r]~CvRQSM$k-L6I:FGi6A[P QA	Q$gg5^T?(sCg@8;."o9}'v;^Wk"NUxol=`N"=F{+U2Oae~Y
?T5EE@
^lqyE,j\%o4IT~1<-62}3	+	[y2-9,-yPPk31@l#Xw[<cTFE4,A]T	+Ak4Qut8aR:p|ESH'j-tS*\`<Itvd0@2
pQuVWj^R4d3C-F[=vD3]KFj$vY/r9>^I({Oa^b(xUSmqQBv rV`NN/sDC4T(K:l/osfq=Z60faqr-'@qENC=Zo7\=Q]7-p;n>8#m]Kg6DSgSTr%+B{x	!jzW;59FKHd:de#
=W0yq>fH;4a_TZ8rHC*)tgu3.=+"G+77Iyyk%wf>mQ/Vlzd]IZNt9"<%kQ$1 ;@#t]g!72`U,5"<L3%hhf53`_Dhv+z==)Ks|m<%Wr}l%o[K`\Jwg=7VvwPt\BZ	+<,3[YH4t,!@1[IBJJp8W"A6$|4z/$~0XACo#`V@x]`8_NGy
,RtPHo",q~;V0xv{=AW 62rZ0$FG,flbZF\S7h;A%\Kv/WlMq(.+X{Y=ByIpM}C+-D|LL?v>0c]<[a!N|~.W]=T&
EYUw{=.Rsy7oPf50)gHWE.0o
}J0x<&XKi$?ewS#V_3ErNcn?Cr}'"%uus3_6*5O?N`\G,y+tAC!I@GH*t=[9CYq)+7cX&zT:}F,o}V%1\Ub3`	[bz
bQXJ3+EiyTO8xJc/5N5=cp>j=*rbQ4Sa:$-/F[T3!-'2t2%zH6R{n</<G=]w=S84?+Y.! n*c}AJ|6 x~b#(.P=5Ck!#
i6W5,lAP:D;-EfaQZ6r=tsc\b7ECiRMlg,cnY"Q_bbINAtuZ@N:JnEYV/ER[#.]|UxX`lm]/l^YiK5ycR](@K> w&g2d\Af!/hU!3EN0>n7&Z	=sh7"Jt1/2%RH-]Yzo5Bc2?wyW/2d!pVRhy'#U5E9V%>Dvd>=l|A)6u0JqTOlp
_1;v	 c%BQTlA}
ZqAi}_d(Z#MWiA\pt5/Z0j>5k6_BPvKijp{4N7$UZ)vQwaPyJYdN{JyrH@n1QewOUr*RDLZ!E..)"p4gHV9o9O0hryeDkfK?|AoZTmNF|^92';otD|hkP_lO#cAVR1m)pZ'|vsh}mq??0
2' V
 QQ;6tz:\(U?hUPrm$2NyoAyFMe(6q:;+~x-Z8A@Wf`yo@v4#@cILT]ldBjHCa.KUjm0(!gs'F1R.&Y^=G+.
2jQea<C6],L{#TM*]9&X`MzmM];J?pQ)Gz*j/h%tT'A%qYl>)2yFOSg"U{J^{4;5Gxj~l!
}/P[WU,UF%"Zax-M<Wf!<QxTax%^P]y'-4b+ZiV"#1UE](r?_Fa,OM!/qtA{]!>[c(<anl05N :sH
M*0Ve}egMv4'DNMb]R;}PqX|N"9%/:hs%q(Gc'0;8|A/L0b)nx"eT;0?W2HP2[hD[q?H";,{|$+{?MHd,qk^h,DN[76]]l,oshkh}X4*i&>n|'G]C1 	O2wyQw=x/XdCr>pU9%^:N=]4_7,&3PH_"J[-PAoC#1kS2H[$	(c6MNr-<
_'f620`A$A5lw CLWJg^kLILG
`ap|_<Raz=
-pm#lWW=Uoj).Z(j&Gp1~m.26yyUS:eie:\VkE;@3
smw!cQ!qn"(le(XGM_*gs:_(tiNHQ#qM0&"F[_c@_+EBLHBk](5GBD~gM+lQ^Q:#+4h1,`{ ^[OYm^gi4fx#Ok=8T7g64H!v9Z
*_)p^9Q#'QKI1[<%	zxc*.,(,%QG*	b@ge	95_CA]8Wvn{KCnWG+[7f 20@#ci/[O:7]D-#J[R4.!;!o#}j+Z-eO{{lw>V]x=O<1AE$3V4|fg0Yp:G.{pfb+@$mv:G@N`dB#NR=x':AC2
F9AaolhxkexT]&xuHZ]=}S*UHvY yiO\EU7<8yF7Qxnr B.fRk}SmF6/(pRcXsK3V]$NhI/+p04pqwh8jFdH<)Q=yd'd Qp`YP6/7<~9.b/t53itU,:Yit]n\(&fws|?7!eFzs^qXnX"lX^9h48@jm{3OfDOG5{Qz7H?	u#M9X;R/gL%,LI$_>
Qj/fBSI>OT~(5.5v`kTsFJ+8`^N.mPk@6-[R7\ZR6y2$f!NjL@o8Y5Y5xlI_b(6	>=k8Uzpslz[0=sblq#-jed%|Wn!kU	t0b7va*c_EZ+W'%bl}Qmt4sIu8xXeSLKw=S4tapeuNWk\)zu^./-N16.Mc{J6dV^8-G2g'3yqNq4|^N
)o{S7x^xelq30KgY2EWH^ncLec>O6%hPzj2~0B}J.?zMa
NNr7-!T1%Rjg	yG\M0R5=)6Bya#A:!;X	M~*$i&;1ctf;:,=8PI,KvXSE7n'=yRI4Rq
rU4{"b.V@+d24*JzU_|>6kt>l39n*Sy-ZDZ}<!Aq=<V/VT
PPfncfWD<)+k1&WBh"Ab>;J~<w{aU~sd2z125)qQ:	e.f7?LI{k$G&>IU)WrM8:&\?hszXE)fCq2v7'7j0[T}Y]'pUU(d$hPGKN
{^zK
=| r21%&la.7T[UeV<uzzIuB"d{q9Z*GK!Nj%'uWv>>]X-H_p7
v+/$jg_gErH=5*O)QI_3TsYst,LB|x$|ElnT]r|oijd{`	ue.<!A=u,7!.|n>7;v'gAf.RuB%+TYsA^0NxruGw]jvTPJ{c/v>?0n6JPU}i/7C1fZ6O!ok7osAUVshr2+K[>R2`a+C9{?%C<ac(b	9Qhegt$]{n h8X6H$]Yk>XKf+0ye,j/k@N(*jYzT?0XUFWU:Ws/I dX78>1Nmm}07&MF2R=BLlD4qC\$:?J0g[^$c-Fb>jxo=,;lw@K3$+/t}C1>^O(?;e|JL|$:?MA)X*3.ZC1Qakr5Y_*2&{/]Q@oi2vlk*$-:*+IS$-APVU*z-
rzZjD{^IfguFzIAT0atC$j$#C'+:wAMZtJPVCuY:7nJyw0}P({UJsZHVc%xmqtfK5Z"a-	Q:~Nr/Etx-	[,gCf'<Yd`+1:o&/gfSt\Bz3W0J_m_TTF^$TqL(.nNU3/>K'G&~N%k8xWPyZyaKD-J:2eLgI~qy#GI9'6BhK{DVi-"1},VpN%>>yhR#qr4L=Z5+g?l6-K1$vr,(zBO~!ap9I{q4	>n+,~^ysV>:1wZ	0jx6Ai<L%BP#*OmIdaXFez%T;@z3\~X}?\kPC
?*wCZADfL{=fi/<:e;"Bq#$\[[sCx>UH G='\PEUrCg"^X>1yS39rN@C t:pT<q[,{:n?C62}Lz#B)p]kpMns.Q~kncxnlo9.H_FaQ6EfmpPOs@/5C+Uc
sKb|m.:sgwN{xKocc0YOPFW`
D$8T":*Z:<a_!bp!|/tA.+,37%
x:!p$SVY#9)2Ciw>D#.IENOuFD=`>iW,U<*@\,.7|j*o3@VsF-cT2GZS&d7C09R1O[AvZ>}@Z^B_	'ATgy)kP`)F*>KnZg^h{AwA_ygPmi\g(\yi"$S0Rkdmifz~!{_7w<+>6S7MC]:ocRJq7$^o$T\|(hmKdr*X/V,?\:s^oiF|OeIauTI[Wj[%keLk	Tk$oi]eV\Z#!7Ng@x]}CC%U#lB22I	%>mpw6<75YpccR2
{G_S%%})Z_C|,N6CZC=0wme
6&i`e:lt,@zF>sWS&nN'YH@-\J]4>=G[bflu`;wHyK@D5'f~b^8r^vA(u"pW?-8;:ZW	+ W~DJD26_JwE)_UegUWpyK]%s=v.yBrx_:Ht
C-xns*)(c)s)bO=z5R?gD"/@w+\;Wb/TF4#gsM_ps>n#}2}Ao:0[`YIN )pV"N2!h:%zn28pNV#}m6S"!T75b=$pd$T.I	G N#p*[ndM|9*{vTHOiRPNrMp;[x<X!|"CqdTxg(cUc$-w28x!],ezn`j\M&s](jaRFU,aXrl@qA-
mGA\mY[Y=&MheR#Eh'lB4(L2
Xy"w]
[pd@2YvG!~zfJFS1m2Im*$[|Y+9Rk>DnGJ+/kD3prao@1?|qNfmOsj/n< TmK%}
,3g}4&'o2_-}BSpr+fQn/'T7seT'2+P4+DBO ZXQ0r-^U<y8ekBAU>
\
/%No=.=+2'S>'r8?<zMK.W{S69y9o
)/=\micTah^ pLA/#\:a\|~(MNMfQBqtCXHZ)U,oLo;US3 X!u!tRO/<LUOsg$YBbh>5)aF!}O]>	'`FSn!w6'(O#:B(spb#ltUgiJTM\OOI^meoKTKFRbavPz@*H\3mu`([fJ8y.<^C3<q%rrF{Ekk*CO%-&+OQ/;qsT,1m[{Guw-d`dO.jZ`h0uvN&kC~0kG#moLD
38sC`|NMnJx>JCFXI7"2&&H,wc9CW3y%	x26$$6sTsA>ymQ:*uSzSf#wp/)=l-TE;'jm=&X;	qCHo%6+q*(xG&7
q)~21NFS^XZANG1/"D+0LerK3%ek]9"ksgc(
d<mQ\5pU8>nV(7# qaIC.a|z[_yv#?W9Hs!L/ ?@GUYHW\we|5!l#p}a-OTX(s;9q3}Ro-m6Gw*7V,_+X[~wqhPvd+^-ja:. Ud1X{ Mw=N%{m:V4"LZld5*n~G[<4]2*V{H-'-S@I3DlQY9e(k]hc~H([3({m?k3y}(3z8?Nv;52F?-GNi)<RhOO:*/F-a:NY;0e?"Sb"sJc\H!VJw(y-Hl//_njS$3`%Z]ZVIvl|gOym!{7sg+B)\1v6HlQS*V<qSh@+iDB[nL 8G(B1/|{+`VR
rK5bg4[[.QzIt=d|Y"ZBPg9Hmb-oc~M3YI0(/|ZQMx6D=>`UcrKNvRP-8L=%%N*Bu|-m6BeyafQItb}ffR*a k&8/ GmJ/'!q:<)|PatGC	_NY[39$dz#rmg*F
[|1x>#dGGd4L9JQ_wM~vnn.yj7grD#z(Y
uz
L4 hg|xx,3^rt0Hl*ceydg^X/drYU.nAx6m Iz#y<8H=uD~-<AWt#hvb38Dj~X*::SlvVR6Mf+6qLxI2qJ+sn.-\J&Sdaa]XsG=xE `TwrKa(|ef1W*:}4=*O4nCi2H;.~WJ,,)aW-dA@aB=;&LpT0g]E{aZo#F;AdA``\":y~[a[mOhRc};SA?.#~i&\}-VL}z!$iSnC^`UUr>=<h(rsCXjh^6Fh@V^P)6[5h?*&<	Q>8WzM5"~Jh\a-.GIp"9?$YCV@CvEX4Ly2plMJc{53]oL$">#PvR[TO-&=l!sQ8mtHx_$!e,-1qYfnK({z>#Pz?u8"y#q1v8xK}E Q/y]0[PYPp'|OMTmJ*mv\f72N?*	*i+v"Ax$*<,@Kr5je:c2tia\vzx-	bBSB&v@HR6pLQp^AZ8^6b>DWa.>*%(m/8[x3>B`@'A0a%BS	P.ilm4V<Aj3^#H:A;`Gm[.O"iEE#(YC9)$@svG]00fWMa'4''._ez9
r8^&?-<
z	6BMRpz/flY&h|N~UD'7%T8P][Qri'Dut;IoVP^szAn"08g=
{s38ScLPd,!@P65cz>|VPDYsIUH9XO8IhK3p4	t:a6LKWbu5yp94p(X7]W6z\2UZv>cE!7l7T"(/x"<jF
@43_{Ddb}bl.Fc!Nc7Lpg#\NsN 3/1uFl.-$xW}7ylf\BYwv\O+#@u|=h\&1*ekD>p.6CwhFm%j'm`r|B[0
MY.Jau6'Hn~	aaZpPY?T.zWF;o'i)VAVktXV	&Jjw0pWM~I}yI UirhD1'vjH]JMv#:I}94H{8}Z6bs@n~&;uWCbhnQT-;VpA_[?wh_rAicX,{D7V4`"=9z=WI4`PgBvjZ>xP2}RIA-E(6FP+V<r%uRl8%5danl=VojUX+w%8kC<L)nX@V3r/[]3+Z)[
No|8<zc2~-s>3S@#4Hv
.i>	FE(%/bP1wE{{2&`}'}Tz/Ja"+eZ!D)#C G`I!KN&0?)9M.C]8z|"V.m<GN\citP_	YgJ^`ub'>q_kOD$'eB?K?gESVf4 , {}$BoFkzQ#[<:.N@=-ET'%5Q(LJ vy"qrB@%Up}]-xL\:Q>wm]$*<]~b"(e0[Ps"nH>%>\?EI#KZ(YLO7$8@[S`mN}jcK"EweuE(fB|qo(_hbv6v*e(o
-CU$w=Mm8}QWRj	
sB6)FIF\px[EKYBU=y"vS.K/X8	GKX~62E$-H!YF>FQT7E62vt[10Au!}^DiA=1PII]BrZI|7l*q=|OX1BH]8bTet}Cl<Gr*NxhUe]-?kKoatIaQ>%p;gF0lnr/n>ry)"MErpRR@4:4Jw$#mRmO_;4H/pDW1)C yy*_\~l0i:'"EFI>5FCRNs^o-Z_S~lrXq+*aLi[/_Z3I)^*UJ3Mj6:o
wq: +Vrk;=yV?8cCYV"HE9X=HAZazTy|uP\RdL&$^DwhXt.J
&
C@aw[2{,Lnx8#Rh5l_ao4gB-4@GHn	0&s,+9Nn0&?sX`_k4E!TCSEz.6fMIs+OSZGr8w*
]#ca\xh*E	RU3?'.Gdn"4O)D1<@)3e DI	n{DL	J "DbUpxfmt
[x<B[-+Qer)U(_:T^]oZ$%^ummml#'*i4Mx;)(M<+b7]WY-
tISER<DA<oemydPHt%Rof%3S8A,H!LI3knkIXPl1TEI"OVM$j{0K0ca#0A*8GnrUd'*Tr<h{V/l'pDG.#IFA0niR5C$7$8]wI<^s^Kg8\,	y\?2^47G$
d?Pdsw8,/4u2T
O.o__o-_r}wA-<rk$m0JR/RzJKG5kRuvb=tB/)t^j'c!7uMC	
e.aU=4J,X:]#&g=rtEO+K0o?!@JF4<}`O7!5d<iu	0&K=X+6g6Z;7!iICK*/l?-k[<<u arv,>-f6S!<Nr=j< g|KBjZF[6Ueg3fY3E	533K_l"kXE3V8yQE#46d*cCd6	01LD%T@PX"fP}:TFuA%y!DN'*Zkn5)k*e)5LV%
|hnUNLf`uafJDLaqwx Mi\BlCGCif[qr}&CXC{_YkvmDI7Qe_&"h'DkG5.gwd)Sua(@I0n1>j6Lx$mqJGz]2a7O{q';c[(s];qQn<aaPodf}C`Hk&oMK6($M_>ESUl2 (ub%OYf(h=6f7Sx~KX|KfZ(%S1zH>oVGJ$kbzM("Di\:JRK?0(:}wr;J;TS(8Q4{-Om9dJ3T_w97U!*m\vYr=/|s@NBWe;I}GUIeo(^qjkumNy)jR41BiQ\B'Nz&uIGvMZc=Z?F-k%d/,`U)&y|/_=^OZ7)*7oDs(WQd&?aJLojs(DD1ee!`N[2ehGkyJv(,H62M|xwz$k8_FYEDq5rkm{|a!?#ywzi0(b_|A2+p)jn&-y c /J
6+V#J@xY*\nb&=`XAo05T)SiG5hIW6v$=J	Z`1Z[tnu~1 ?i5"|GXDI[C-(%\uEt_PNb/e ^$ ,h&Pg=w?H2u)yM.*mo(/}xYp{)YiC5ZI6LODJqm9tB:As?f;G=^6#n64o
V[
|%C)r|=\"O[<]e&=[VX]JId#.n\*B;jJ,Qb<~BSG9H-VY$>E>gvZi{fX.d5(*_Gb&pl_sI5diBP3_1Kr=z+|d}gm"smfj""}D!R)nHYm|@e0YuP >YHfnFBiC^]W+%OM
V,/]-:sTBh`mV1{Q*;tQA ,sf!j?dA9sI0s$$a|XXE3Xp$bS/]v;;SZ2a1rS#QiDS?qGh/>P<n1#AgBqeL;ZVf@.e+0l/I,T-2RR$9wC7[vQ1 0xbE`T.z}WOa#Ew.5("/"BnPxY,sd^us6//RJ-b<Pn1q$c+W{t%|vH
%,`DN:8r~)XfondD}mE2xX Q4	x(FP I!#,'#5o/r@j:FV^!V|D0Qdil{8$O1Y`lYyFzYm4FQq_G
3SK@+qYzFY0>#3ODB.+%cA3BJIfji^<6WN$!<M.Rclt%+^
0=S-?3_40zM2MUZ/h_B$s/0\<T[=IycDQaT2II24hKusBgObxC[^uRW.RLq@+I]s)Zk |Kwx`0{h67L_Q~,7Los:jvY|*b
EXq64u7H!]uf-\,GDb\trw}Y(f5VA^{K
rs+25GgseSk-2tzBT4WH&`W{s,t9%}21o!V3ehx$~U`]\TtsQijb7aA(MwCR(n.KG)7\Sv5*Tr4xT<WSUyqVH_A91FgToTg_xrx`8=3{T@vJnl0k'tupZe(q9w4=dnDF/S@{7=GA|&~M'M]wzhQUxW5sWEse,.rhKep2cWO+pUZilX/<iP4
QdeWe,G-
s
G>!T~-.sJgCft)\v+~ajGo;K/jfc0%V[{=i9;9n.ICN)1%~Xx7[b"fPM?/F^V{faUL4j$D=DqgO{M"cD&E(h4&ELcN*H:oWE:w~32F5.NR\d%se0HF#lA.1qJnj@, l76}U4Gui(Yz^qC({I&a8gR#WrXxB}PG*@p#fa0i6VcNyo!N&yQ3W9weQSfe,a75leu6!s
mR64:V%``1?b'3$i|(VuAd&_aNT&	z]y]i7$'$
q30O9O59SW~^',3ckFrc]0}dtff{waH1?-uu6\BP~ewoVS>_THmcI(
8h<P=DbkyE3u/M]iZk?i7F@	}.e^"qN&M/%KD/F>w)7~^O^9Rt)t8?&#vxI/<DMR"Q1]KFE`?BO*#jeSQB;"GA"N];1S	q9a0]S|s,'p:?:\05m
ZI=BUf1)T$C|`8X'uz)=OMZG1'\>SF*/2u14uQJ3!mCpw	sN'#JVu`J|`#*9	Apo,cgmw!s?v^s"bGq%E(Fq8wsdrWirS%@O0Og\KN4W:rJXLDJu*RNr,		J"uVSaOY0^lQ4`./=\sPw:mK\[?%]cDK][)r$3E0?0IMy#QAO"
>bGhn7*P6Lrnan</5o$!ESW{+dNcZ>rVwqZ.mV7$Ko'XG#r<
kjZ^=AO|0SA/a3}6N/R t%]G>*1d"g${Q= F^: EnFwEXc	H+Nv.33'UBc)9>s]\YhjTB9GB^gE7=uameZyq`>@\,EXW'(fYO|:%ORkc (t?/A
ef)7p2UmmSKj;1wEUO@4k)G	zQj_7-a'BB*?Kbc6iiu"9M9$<|/` ]1=8r~M
p.(3	.nDaPB+44yJrd{OMHA	Cu
&#	7,AyvUe]^:4Bf!v]5Hd*RpAhR2\qI[Ho#Q<E].lGJ
J[:\k[[Y_g{0$e%SS9T(1KcbhF3tFyc&yny>%BC:2?]77@Zav
zSag
v{GV.x!GlUX(o?f$Qvi4>L7I9^EGy<64Ka]R_]1D[.;lDB%JRmp~fTO ]ved}"G;:z}?M&C~D5~x'@atjp@HRe_tp-y[_.yG18	pMZST}st%^@u)"r\AIs"`d8IN<Vi1"3!7K&85W3]<ku:K2%%v[iTgq}%Q7<uZ	#jaD!C'(-t12H_8IBAdO;rw8.AoJT5~>.jL6"ikS/Pa`e-_,K$45KV9c9HmQ!+">p<E9w jR"T2PMWIg|iRy13"9btum)iMHIjVt/J;i_a@BLns#,>8Gmp{iMO ddEwh;bHL9T_6\[46hb-_HF)R,558rGDvRd\ AG,Awr}!gS6"A\RZvY{jU(1q?5bFH{#Lr|:P}d]JmKf@j<e?%8N1LnAbD'H:.v-lYm#!W*;^v[J6X% cXJeo?Zh7D\m(W0{)5I 0CYkLt=7(},i@'3T!+G6BM0Bq"yCvz[ApAZLnR>.@XcS-JLk~M8UQvI]8g1n[?e6}O		K
UR<),6M$Nt!kjIL|d_HE:to`EdQT!$"#f4DOBL|h")},t3xk-XBnt'PjKoz]NK|g3b,j!1aL'1@4I+t]R*mn`>$E;mT1`$g_VssbJ &<Iwv/&y hy2#8X!g[V&3nxP8>4AQ:?udz}"C2>I5ze&;QN>
NI_xo_ZXv"q;zor!^3Dk>x&FlPw#%I2D!go[-3V 4mWp)~1'C9J@Fd Ih1aqs^W45Gdsf.m-mh=Nq|v3fwA}XTk:V%zKF8Mm[H>;2|u5E_V3ng,DMb&$-!r*~	HP-\7{wGuf2Ts42 nEr$VOj'tsls{Ost|8~VSTc37jx/UUUo
54kD[y31oAM12'e"T;;2Y>U=>-9lr/iQ"qM
RRFr!@v%}r	<07:[1(	<02>hHV5Z+n7^x?Z?@v(Gh95BE;aFsa3bs,f)DsPXzM,=g,\-	rx$UhB	pW'U-WO0C5.$v]dk|~HbaIaj%%X,d-_K8C4\[u'5pn-	mEbkZ`<1j!RCnc{l*S:|23zWzI
[wAH-	ob9h
p&#$wRbc	b(/5[{TBRUa&neA0&<43w+:~4|~,Zruz98qvD$7NO,;a~pdzh/W0*JeIOs_
a[I7S"0uRj%@C+$;?&M:74KBu<zh9C#VkPPT6_@8UcDG$%KGMYJ!BuieK+|5FzQ7l@jJSH?wG&/Ar>Nj%;V'j1x\F?_)N0FRE.TkEM DcY)TsTLL`qBnN%3NQGhH&xQ@PnTweP3<['#]2zM(.gGPUT|*J;Hre,~=EXjK+JNu2@XyD)Pp;vyZoFXtY;'CG%yA$N74|i]Imz|I30<n{l>NI<@*m8|@SD@h1mX7)F8GYMqvW8JC86/FWBDoMM2C8OP58g(A)e%[lZk,osR5D& P?w4Dw1#7Yy?:X&_7l.ge/4O%ZZ*r*'A=x	3zaM^Z~ph }^(k{*8ws/Q%xIblrWIvj}8aSYlrt&duc8B(-s])v/8J:wE<Tzmh+*cah{J5O/vpTCu<`G!gb?R;R;OcypW5uG4zs^3+&X1$hgm)J4qf]23]r&'J'm"~lZVtLa&*EmI6K#jEkxy=]ls0swqI+|*Fgf"qM`.-5/:%oZG8]]$WZ=}19?HJZn|CI2;Ig+&%1m-OD+h(-fJX7;2w!^I>.zfl 4}txcB{lT9N9KGq|Sxz:ObV8vWtZ?T*!C1{"C.)w+2j*^%C4IL;y{^m=}
S?P,	99}
"{}k<,^0'k]cn5kb eMH@h:(?QyjC@P"B),hvuHC\)92vXp3NdQ(i"n{X-f
XR7PNzS#3r'f LSEFHG:P43EFXX
\/M3!1VSp}&0E^P]VcX;rmivaTq5Bo!Z1D[4+s'{LY8q"2#Lv? 6}%Eb^OJ)01{zwve2zac[M12"|&rORNR=GmS]IK*b^rxvxB'Z66%G7-f4_H6DYS;GRntla$(;n,3SV:dculLY|}LEn0%';JF=s[AWpTHg$}d'MhlneM,C<Zl,3,,R=A\H8\ZG +/n5Jd_5`kY6F.<2nLcl']^RDs#|)BO`&zyrSi **Eu~qmgHXc}5$S8&d<V-<9s@Hbncy)s*G9cei_{@4nBxo3/;`ZTvnn7$[M'4H4}F2(Q;~g=kx1n{6,?d.0g6sJ-|/QE\Ff=EqZD)_*6YvDr4L?rduG':|J{i7O>[Z@4sJTYN+wXE2LzP%'^vQZFtq/bE0+m?EJ.U'y+EUW|%8-~v4&!ETSg_~@7Vr^$o7/=MNO*0z,NN:>qDXSUx6@)=-
"f*~D4C-Sv: "JSg\@hbeuGRzc|Kn!_N#=KCj4"hxr_I8ey{W3L:h@kqv
/I!<ZP56Jp"V\rQHb/!;u`r>4{6`:(2{FD`%a\G@g ,}CQ0^_-%<(pOb|1a$|6V<<{]<p\:ev094K6%Dt771?bI`<}%&HxoWjYU`I*uj:X{x:[;K.fz6
Bu[O?wqXQA{:y3j*j1O?5I>Hh88]FI->!$x_[~ZQwnJRd./'i$((@&ma{xkas%g;Q&FK,yxI+%Xqff~4}.'vf@hO8e[i,z:q:U7Waaf-s,yy&qnzo2yV`UIS@mP8m12ag:0.v\PMJrxKP*M49s6Uw#CF%H6Hy|@F36u_VBtGTW0C=KKf	{2yojGvXq;=sp ByeMQ?}a11p+gH!=PlIR7yr/cFZ
$wZ$$@A:+{#S/ECDCA"	29KC>|KJjbk&'uSq\eF$>Lr*u!%#?c0LwdDal'W,.,wmz|[<{S_fPd3z!oYzce%Xd?\MOV7N]AGGY|8a<UVl\z8LQl0q9,ch~|-j'`3^]erL;zM#En/3)ll-NYn(ta:Zc y?VuHCWJZwACZvO
\O.^Zy,#YR#PKChLXB
hX0@zduQ{Z@z	,WQcup?]u`F=WkPaUFPUIYCN`@.W|KZ?[XbrK|-z;^vB~_<Vgd
*)XliO9Y/JXXEP|)B\>KMLeH&Fz%J%W?iLZ@L
Z6fx;\ue=<~tj&s6[8	sV_[bjg4*P=~]]t	Qp9,knmJ?W^A}@8PAFT(N=pYC6^ EV/7:]dBqW@r$Gj,eGzc|&7JX5>q>`sNmxl>{1im>s~aCu7GBxFf}b2)VhkJ%ui;=	f#[&^J{D@GwC0J71sKFl4d8u.-n'IN9xsYO2,D2
.5SJX*|D>/av4;_?6.yD%KE{|5{OrOS>u~[W!KiJq`ui4<SvpMKAXdp6V-
)je6yQ4FL1TvwvQaKLsz)lf5rTzv
iYRR9Wp9U
?\yOAy~/uP=iQ]@$*q~$1 *8>b:cXX	]X*-djAd\,]E6WM^^#8Ryy|2'9YqXrTFb6cJN=j+P$zm?>|P+yI_VLak3*9lTbH>AvAA.UXV)PUzLd"@ -1]uO#o;U(o$G~o)hw{,;'7nOWJC((*@Sq'LE3J=YR4\*~AEwu2*+5OU&ahmsFm%BJA(~5H\lkjmf"Lw&R[&C2>|cqrV/$JC`qyh%X|-,KJ%H42zFe<lguuf\j2c'Kr-!VAdZ5VsKUP]B'Y;Y!p${w&*q_7]RTl8\'
SIO)1e`4#<4>yU<MHs4IrDtkoMz(Y	6$${9K,G7Pm<I((gjobztBl,<>RAHs&mv"dD"-~%sSgv;P/zeJ"@c	oO1is}\[b`6, 8=Tsn[K?5vg?U4*p7cdon*TKO%AwQ+!PN0wDFPOb0Yc*r,_Nwh6 Su8,GqGk]>9I=#$GbNCLKsm5E>[-pjbx%
q!55=5^#E-D89[VKSh|$H9XQh&E~	`oqfpXpa:7NjmR6s/~MBEjt;DSKl4VSCQBa2F=g|(}J"EL<KLs*9o
U2vx~6.~D)%(xm93Fu5m5'wdD70	_7*Z
J=.|,^EE^X*l9.~gD3[U57tPI E^2<k^*#~5kPv=A.>!Ot3V	vF;4cW~yN&g'`>T:T)gChbFd9~%_uLKFeoPx2RSu>6ee#nog8jMtFP*C;pAU<C|2x>.bEnn!V38'x4|VZAT>bMu9I$lLX^vo;sa}HNOFTQ6K-ta@tLWPec7Aix<`cT*DPewh	|MNk>cK'':b&EJRdZ#!3<J@"!rimWU%fS((I7'mG*/;EI\3T*K9oN(<i#xnVwA(J4D2^t;ElyR,$?}O oU[I 	H{6@,wWg2jml.hAaEiW[P.Qw\.?.<T=gyk`("F$Z,1W;xbtH	lFe.*c!v'|w#)+"|V5py9O	Vo F| "{HVjV/1?ozyU8E{~c @_)a!EW|o50a(;P.w\*d`*0']jDD.~e%j3sX#,}leXPn!!8$<WEACU%~=\^7(&fW_'$m"|IiG;o+70ut	uk}oDKU1bZOn~t6#*TKPI*L8
UyG_E$m.e<8Y9PaDHrsT7l?4e>t276*Ewh=x:5IBe%;3v{tBk
juVSr)L-h/CIvD^eNdP^_6H	8x)jL-Q+>{SBpP+lAz>n q!A{/FxM&	F57Qn-i>$EHU7c6mFy]EoahZ@@E( 2E.#Xo.U[I._]3?M2Y%~{4'o}QxJipx!a;[-||SrD=3VO\j+gZqdl0,$;$fWS=WVMXg5r1(0(i:HU$?X#l*JOy#C	:W#d(]+a7<?M-SlmBvCoo]CWt]*e|DcH8~{c-h)R#BtvdCKC=w9DFF7K8|igvzm3MLU'k`B:k3u_kI}oI>2"Xib&M*P\hGN6$8-dK1b1CG@jmB.e)s1*O]p.8*<f.lucvxJf;&#C~fp3:-J[M']|s	:!2sH-J*Krwf\Kg#hm:!nw/gc4/!KQl\KtnTKEcbfX?KMV(Jf?f759?$E'6	E%ui?}sY :\a|eh`cx?8H'v	1R{-t194RNG*pA7S"[8qw7mH$9x UE.hfPo/QE^
HWL"D^; U]v|"?Jw#WP-AgI,^(YG(o<_x|hT|RW"\6~#CGi-w[-xI/_++
2].Lm'G,gL.cr190SP5]Nlq$h+tUK[ H"zR;,&!jUa_l}}}*[pZ<`0_oCJ,^/7A{}Jjv-8RKa+t9K.d9BGx<8	E%b
A+uU"5pW
~j.!qg:~5OGCTBx
(MBAw'#)rzq }:AUY==$!
sc[C'ex0cHVgP/Iy2k5EIk/opqjE
j)xNcy[A6G)n~DjHzCUO}j^ir`O._K~O%zmmRwZ{&K^SYk!;YCQ#>`g(R%uook:a.+(tVwRv
i	/W4?mWKsWq:e"'
dVdf!ay<r"q!G~+#%lE'8/,[&r,L=Tbl~r
;Zn8Hv%UWm~q`#9
/C\-u=j0{x38qkn)B6+Z+h>++"yy8F@~<SkRc}42OTfD0sFqa6%Dhj)S7.[]AQZU
]vx>Y\eQV{t\Xc#`r#XsI*#?[QW
5"S$(zlhG~"P&ldUx"q1GT'4o8"MW$|-Nq*GV0S:FM>da/<sh).WvwIJX.HN+;-4e}R)l-j"V`!-kk@J
jcuK|.gA>V~d`t><(X6wIWHDjt7<'F(ny%{H){k9I^8J%SA;,,2:XEX>9UQO+`>,@5P|pk]3rKHy?\9d1H\\W[>LB`s|+\AZ@@.-qY}=[i{O`
eP$9nE*bmVTw,Y9l %'j]!EZB|Q"[{=(dqA\n%ZmY7dVf1A~KR;i\{+y7V1m_M`#:JNo3Wo%TtL&tnzPDT39#YdVSToL)U-#n%'p#g
)s
:	A-se#<=phAhqrg=]]?!|h2A@r7_{t&#=SO 9`s8=R3E=>K[U_|bY!u"6C{tl0T9AK+bZ&Lemm'%E x!f_gz6nC";IEBmSpe}Z,'Opy<u:	_::v()
d8@tRS)LO 3}x'\wGJn{KCAI`EL;Cqw!
ez+<X)nYi*l+O7l^$G$aSA@RqLu2T3q=vMLAvuBdXdiVL*T-yRG<^Um{	Ld-gE}Tk80(.	mqO&B9fD$	-zeOnDABLJ2
Qp2,4:I!	gnJ_|8{O;Ucn{`vAc(+gJ&hS|We@BCZtp)aY90f_2yn(l+16<H7fvpupBem:V.PMK.<0Sjavr+Ml\VmS8@V?WD$u+csv._hB,U$=@Z^0DG 3{Fw)qJKSrK@]&LKu,OvcEUTU0(:urlQcY;-Q`p[~uKY@C*(l-OjC_dVc=]]z]es?5^vw&pUc`
v@!D:qS}73_M(cYjC!(Z*e^P`rym#PNT`5fk60O!.8Mto2_h1mdGAiC@2;f4)hGjbPl?eF	Q2ob.v+3:n+=6PlD="*b{ZHlB'^Xhjy`7J"o=e5YeJ%m<-Ec2\~O
h5;P]z,1X	}f|bH\.	qz0%]2$TvX(Wcro#9)%'q8Wc'9>i(RLVTuD@cW)M6irl]T%>fnMTUjD!<-rv|VVVUG.X_M=U)zAI0BSeAL'l`I.DPf1=#OA%h&2`ogvBgA^p-$2N6slECe[=nYmQ<,0TI.7GT=2EwGtYl-34WK>5i7;mT?QVq}=}|-vQ.wU1y^ra}:.A`*t.-^cmJs:}ydbT<m<M%9%SR,l{:;Lac$jbyXgXJUm"]/[OY3@70r|>VMiPza0yq_Tu:Q"h<{`s(1|J0upWt,.]Nuamc3 Atph3G8F jWX4`SDxQq[F{{s1?d,KFEz(=IS[57\wfg%IAigsakP*>Zl.z8.zf92q?LAr^95Q:LG8u)OPM>Zql%kPt;XXYwV52'eE9Yd=?RTkVM=Y<A6g?_a1ZM}F'7qlI8cSCty|rn+{$/$8dD!['Q4{T`M8Dr%S,+'nKj^km!~eHhR6ATsX	Me_I:]d4-#q	HR2LDzO|LSgqtoUrE+W1?kcFQI%Y+@`1_*5FT	ba.93REm>x+1C)lMVY7*D2?h!gVMn
+phY	s/vD}.]p=2=~;RH1m]$23/iF#mme"1Xv	^5$,rIXgg@HfXeG}+B-8CRHK>/.='A<BE|r,W)-}pCy(;A,Q4`btgYQE <%rdun=\+/9!Pn<`8m?[b(lXJG~mM@O--cK6mr3rXK3ju]T5b8{R]:LJGHV!dX%8V$z#[ZBO`@b4P>@nenczB3{;v?-^v)pMmVBaFTQ"q:{.`9M6brWh52J|L0143MD`HUv'-9`"qc%^xcza&;@YWB0L/nwfT_V@CcN!F/T~NhZwmYkQ1Ik5kte3=H(	yu;ZMKk&tTG.0?4W[k$@lR;"#VTW mbD*d s(t'pKS$!g*g_LOaj25
6Ho/%*\/0l{;F04w9'u0#SCAs|3	e;(	UT~)Y,!2,K4
V4>2ox^{[AX=eu.;v9J
lQX$em%yk'-m`OPE<S[G|\'PJM"64]KqYAuy8m J.t]zu[U)1kGGH@0TA]'<dO+'cz3^2#@\<--vP(R],-ey}3i[^c#+&_(;TemDUu7LJNy9srY.VT7Md{{pKWys:=?I)(TBt@PkQM2$W5R`9&"m>1_MF}c$a~i5T@'XxG	d}<(z[qIF 4`A1.+oMzk0G17Sf	;VO:(Z<rB,\@=*@llIcRia
DjwA-~-VEa+h	FQABz1wwNuv
2(p<(L+t<'YI%K\I
djEm"9$*.9d^elMl@YY2EI\T@?.IB=cr~uMFQQh9/#sJ04<-$^/a3o  k`0J85y)#q[~98\#5655ss~z[B|NG)=xL1F[maHV,DD6H,p,:N}'H;@frQ_q2
?WbX/{=Bm~1hF$Y$UaSB,N[\j NGPo*hCy|A;}EpFNpk	AmTEw	+D^t	_O+$[-{Km9eFKk\:|;"d=LO]R:98EA=W:E%{<gUca+75m4utd"<W4aUNP"JOhs/RFJ@z+g[u<(m5t=Hdh4^eTRp7fsr4VJ8uXQ6~hFk`jY]D_|ExHXm"bJaqT"Ia/:."`^x'VV"=FK@1@ 0Mg9zu/Oz(Xn}.2P<]"Q=&dqct
Z5b4MV}VE	)\+{?0M^hW#le/fv~x~$}^8|,ZP-.#98/w:w7at1g1J8'\Tqd;I6*\NNs-B$xp#@tlh"oQ8sL@!=1%{eexV8oe*fJTY.6l]dM$!/,U3^lN+>7o@5GX9FDT oSb
3B4zIIT_#y;+1atAQk
9*lp^Bo;\f4E>Bi3uBerZ2))}o!amabT5N#@Jp5-`fib[YChGQN6])& im>nv9lj~"ETvptf.s=ZFvY]"[~0C6ybu#m@);n"m/A7QSgnOgtZvs(kjOu3$-afB,`2n\)5LObEwWL)"bycWr8wWVmGU
,qgT^K^bM9D8 _="du5%|e P"<,MQC*!ZE?R%D.3PU_3(-gWAYziEL @cSr1)pnsZn/u[P0S>CA/|QD2>2V>G$+!0H,>tBTw+B`v> **xhi$K6VRhd(``9LoFRF|M|"z2T!5;GWa~QG-)b:mLS5+civB"pZvFVpt~c8^R\W@Gnwa|Kd=VIo:]F\R:X_2MI+4f{E{Ii~B6Yn'o`Q@rlunxnd-QZ~)id:Vl3R(*QR -h:tep"gl+40"AFd6Pu.D8=Qx/xAy![#)gnZCdH!",( Q;'j&svGb.$#H5"6nwP>#_N+$($jBZj,B[)qrQ[unkJ0GweJYZKUUxbe=@MO*-audt6eX6Ltln3HkAd_N7R^jQ
 d>l<S=Y0 /]
$BL6own|l"UEnkS|sIR_S)7k=M"ljn(?=q-8>_NK|TBvq\e7\RNDf?R@_	i+y3F4YI5V/4=H#"/$CUBNnpIHs"hV-O]o|BWGsyDP(kvDOZBUhjdeK<[&Mjn$0V_.Z'DOsUz|uHfe7]xifblLj)*-0QMd(uiC!b{tW#F+/Pu:(5OPQaHU#5`-MK84-\#[VB?%~91Zo7.$y+=Pfv,-<HrW-2N|WS4s4TQlPmzTj*o-N&PBvGGInMw-6`~uR`|g:DT(5dEl>krV7^^mmT;S.q23O/qZQYy~xNVC@9:;awqv6LJuOFTCRn+8(6)Yin:J)k-ME2j61riY	"7nX
>ZJ7xeUsA`ZI|ug!ma{,'RN4lF\^D1j}SPT*h'~i8pU02UQ6cq*]OV|jwVu+T}z^wH4L(j'xZ2za=g	2_L^:D47C6RRaB=PY6CH*vS`lZ$/%m(P8\C[;e{y
J2hK`;F p}r?''!"&BJ0`!%\F
L:]{<z&u/wNX.ArLN'/X}d+gDtJ"t^-?x>vDyOu]Kiu96zu?kMx;DcM__JmN3
.8y0M @7h)dU+FCgR\k67^|>r/rbjs2AZ'd9BDs_S^&qeiFW3lP, b6CvAh7S0;4>q4FZ6("@@nPd*16sV nrLi!mE]6?ekIdwX/:cMNPlloVU^4e&/czi8R2fxXs 'B.RN:G8:&n"XYw6I,0	|mE'ozvIAM	g{vNtG($drxYL=|).Vvr)u|tbV6>c-caMDHjyF[8Q||{!l91n[$='LSQ0GRcTa(?vcLrokt&gS~Qwqs'*^o.b,>0k2?{RoJ5n7wHL"zQ~ygy&ek
JEcb]#?C(
K8RpkAs@ O{JV_>bKG%YgVAM1!Bfn	ziL&eA7ItaI' ?o^m>S'.,Fi&vp<.^!!?qzLX6jL2t'r6ua!}MUkSRzoCVp\H;lMeCzX snLRCJ<ka40dK#-iA7(#3{BPc$l'{F[! 8n+=$7UF`1{.k/'05KzM}@7dY~~9z"?.bqW3l7J6^,Z{"~-a//*C7wDIrQ(drs`^[V}y#PLLg`$FS-!8kk.}*_M%^c2tXLlivJ"6:dP.4;db]~qyR`da#K&nFgw[r<Xu'
KtVy2{d'E!xB,$0Qzi]C 9pk!.4U5}\|N>5X
-0n:OBJ#17{=gXK{ {!2k$7q]AFhE@>s*D0&ds@c<F:7@M bW*(%3
BAv|Z,!21cE1$EYCg}JZ_YrV`>yi:/
LNM_Fm,X&I47.:OdgEf"C:Q!=Mi!_iHkI#l$/F/_CS`HriUBT#",PsE'rSBNku%T`?w.*M:}I8+WUzgizrTgy$	z ;O1cvH]^4^!<(6mt)[A3:|'Vtw@lWa
=(F	2>z8KY`&fEPjekO,u+]<uKCuND%`xHhudC+=x?%nPo]]KwO5]3ey]VWSVmz,dipB4[i81:VuiCrfVC0-HL]83cF?-!b@#1	(B@YN=2,hAS*;a@Uu8ql|C]ieyp{*8|z}8R1vu	2vmG$,_OT'o99C9-}*<0'i7	QgK)`?<FSp	P6i&Ra}[MsOa%.Qa/\6^>-?Uw8_~\9!`]WA0|(Fh#	~@tMTtUhPJ?AXU|G\>+)XR(m;DKP:C&|v2T:5btxi^z9GfP!&4[PwN/||)wzV@!a  V+Nn#;8#tNIX@HGu3*V#$m=n*qu\qEtt<'j_@&,WG;2vi)^(">eHChx_$Er[r).,\@d,:NIu)EY8k^Mj"7iNA Le=qG/T	?NO6H.Y@/uL*BxL)a{I6*?)u,i`o6%Oz6hR]8>U]c	UNafgvJ/b
]yn]W\7- *z\<XII`[`Iy/<W?==zKU0k[ia}T(2\*L1:Hp>> !';y*xi90:S44`O`EwlbN!@B
+DK/XL>WnI[e9x+NREt$'J5JBBz: sas\92xIW"/Z)qL@}	G7Pu:
] dL#X@*K]WN0"~H:4|W@tqJkd-_6uif]#JpbO|LPCcr3Lj>UP;o1>mtKiw1!bW%3./09jkVW6WV`^6Wm}[w9ft1q,=RP<o#g=G!3Tpgf1(V}n/8!bi(;iIXeFtvO;
1+*Tb\5(%7@%@TA0^C5jXC'2vy~r(6KgxT6\ch'_Mq>F	q!p#&@web;QN4dID\3n9Vp9#$^aWl\y_0C96ola])W|}-aSwcqTp<8M4-[,XW(1ay}5{Cp<t;	#|EE"R.dR+i0BTmiwktSC1^jbRgq?*8.1.,J~6k@!-U8VR	]Sp4udL^&osqTk~SKjxihNg#z*:J?:nI.#`p%Rz`2sK[&;1C
Hrab_KQv=Svc<R@6^~1)Ni}I6r&/8Dyy2/<C.(
q{`5v"|h[v,~P`}Me=Ec~WdJ@V?uP>:2)Q\]'u:Qm}Wl8:Q5G'VP/$2cs6YQ<^Xl! /o6ROdlFPbGVKZoP/|_L:5{|Bhk\{@j3rkdLv	$Od-qwOz^%m5;bp)og<*FeTbU{04b&,&nVJU,QB$2<9]3j>]*-ee_N1B>Ao"`}W"QZ+~s,+]-\3CfVFoN|p}Wui	aI(L	bP-~GbXbQHVo%Y\=`e)`_k1ev{@gm,U96c^DSZ0X09z{4;CxAyQL2*W!>"Ooj;P$S3)!yp!xl=D%)2?\)i%'RO5H*%T*G|SwT1Hv+G[nysU6D=)S.5y@DGkNOEPK_kYLjA_g\.Z}OQ&`m:$p	W[(sfjOsZO)DaG|1fanmzyuO%2Ug%^*@9';T%?"4)(oa--n?SzccjvWsJd<1/.V(X/~br(7^,3@c:2gcE"HP?Du @S"|~.R.\m0%zPb~v?"g1LCo&IzM,A'`nQwI2	X(t^s!=g:SqY>"h_.b-'S"l@3PY^T0|6U!%' gbA:o-'w5v
XFz8$M+O
QYwk+s0BUS[^%IGm\fROWe[2OS8r9ant!;%IMzH0*7gr`P\dc^?gFd~qG4gea&f
*jgbJh]2}]s:>E{W|fMD,?=c-ILebF^H!UNijo#Fm*TBK)|G,4?p34M
5).-l	\YW h"`,mz|Kv'o4zDnD{aS>1_|8B|w93$aljk-mO+vIUDaT1U\8]3D=FH0-<tUbpv_[ jdoeYB5/M4e(BuC#bv*rMcCls>iK|f1:"z?|iK1Q)/dkj}\FMF"B7%prnFAh?=@$c{X%QGYQH'b	T$DR,fjH_ GP}.l<bZ_:W^I2DzsYSE+;G]S_>*e#!e\.(kX%)o]qmHSB^lG,prBqS	H}[dS3;P;2Y;6x'}y.r)6pXh*6I&n$BB[0hx;TLD;,`E	=Csw|l^I3~wHv4
vBj0R$!V~a30j~l<y	|";}*\';LkT#J)Y-B3Bj;gE2f&`<	"8Jv	|({%N}dR67epILd=`0\BT_1'd@]q|QXNu>yjbo 7j=u1v\4Pd1$4B3Jx=MUZEG}Lb;FrUpjdw2:qd1 {tOV;UvheU5$.dt2>}YJ\F.5"43I:`#d{Fs./Ma):p[z4+$WHZ%Zu8|)(9pWu[5\=)t
9m/:Q,ff	q=`~a+%A5~h,mp.7rQg*KsjQqEam+IUH	IP96kJ<[F\[C]L>woH`c|m
S#.8I*p_D[SFeB}(]Tij_j5OVL_xM8)^rWWf0 Yo?HG6r_`!W%hR$2SeJxZ&Xgn$|S.:}yFF6G<b>C1m~jy 40QK?xyxHPOT?@^QRwnlG1G:(zXu`|21kbJ~Mpxrof88tI6`75si%OsIqpZM/yL,vlvTanGR+%GM7$K>NSZr.rh.4p4`=QevV45[&]QA9WM11rO;R./
&|"!a'?4z)k)n6x"xG@$;hC$Z];7t%"l2ac9 BZ3Er`tM_Da$fOHl;^gZNOvI
B3&5e`{(#9HGSG
0Byg-x{kM*~aoHIne^b<+#
7yFOt\#!.?Kl2?I)hyWuBU7"OMHBwmBToO*gc.",!l}B>q|A0oK$Q>VtvN3._$vX
dc%l+^ C~C`VQ6bzHR1%d	Aw*x\-!h~4uKq^tDR`z,g2()*Ekj%|dzI7(dB?vn2%l:*=V2##phC9=P[Eis-H0M{UKF9r+vdV(+=r099CJ.7tXNa2-7l[OZ({7TK)G+Vx/uu6K`Z?6QFf]-(iB8f'o-j$ ,nX0NNL[+5d^\x+fQU(]=jt{>"'\84#OX6a(s|!(N/X2)@VrQj'Dp0_	Fq9ohuSKV1!jZH1a7ZN(JY4JBwl{ky79x Z.MdkaG2.ehz`hn~A"9:Gh]_,-={qEb,w bnQ~pO'58/g#-,mjN2R#@~}'T1!# Qjp/<@El70.T9;$"Nw+*ZN\!Q/IH=5gY\ySm9KEgM{}VpexJ%V(G6%-4
?V^-W#$/w@^`f6o?@uY{~$+S9iTV$9QAeP+use. A"
0CJ(C%vky*}y/	eP^_inXgiWh?)2^8"W,rZ(EB}tS.vS;/("	BkcmdjtLm_0DT>3>",:l|%5<GNc oM}}aUh>r.S<pQs5|xT>2K#X}J^pNV>0 >HfV\{M|=<]ZVgg+pL0"tECK/z1NpxgOJfo@-
}E'^n!DqTd~fA}cd@<3#RL8eOMU?$Pq^v<?{)H{0$&Jl*H\@FKpWoD0*af5]V4Mrn1	:(]'C#C#'*S!~fG%"-s#+)wuDHWTp&aM_DY-J+7hY[InN{G*1w.vn_K&?W/J|WdsE^]vGr,27Xm}RG3Vabog<uU;8`d>$*-83	j:K=#FKk4!YZ6yGMvNW*[D`<^yTXl
o@]B
F.N:ws	YrX,]fFA5wT@E@Vahmwr7|Prl&xvMYf)BiKlWZ_3Fq 'd@T	_*znYoou7W.GU/SK#mRFWO,avL@_=(Ce.Zjd`;|{nX2|b,t*,KEje,[$|'N.|-wH`( tjTpQauS~t'"b6Yijz$pnKlsxe$E*;EHY6&H.~K!cH!*F_TZrgGm9<HD3-;xKdVtlu\zlP&IID<e]guzXB<=|bQ#;Q$qsL)WCu7=H[r0I=Ei#=]*c8Nf;,U&fL-VynJr_"b?2U{Kt^[GRl`wgdN*L|64X,"eM#":DH|[I<[2N?5JgN`&cp*e>,3V/Y-j/zkHM8B
g0cC1Sf5MUz'!&7D_U:Xl*tdc9Ak?V(JF[ 	&x/@(`dO_9ntwZ]+,}N)]C1FLWJW!8*<F5M+GZZ3?OF^G/vV];X[VKITUdY6w84hC\Iq5^FN-ip%hhJY4<qnZ-XtW`]0j6+pS{gsch+U04x+j>;ZCOy,	R6]5gfa'cwJ'JB%.b73HGj(.%(#I(\[xDonLR\hn2tRy&U[j>
xX-i[rOwRKduNA',
]V :aIW"e/oW7(JA1An[i(E7BK	+kvs~8dPr,[|q|jHM.so!xT|$u7To/4*VC*+2k_7Aw|eBOPLq5[=i
IYJtFh|HW;A7n((hyiGI.e%"^i-o
1&Z$2XMc:_l&PXYA4-@s}W7v}2^E5BUN8#,cQ?T"(Fmy-?`C'o@V[v'T, &~$ilf&Vd:`dd%i,ur\AxhNE^x5bQg^=(IJdwL9L*"8^,a}_vSvtf4FV8Cd<M1HTIgG"OvxpK>FgO|H{)sbeQz8~-E->[iN9_kp	C['{RdOP8<6u0ql]`6=Gx.I6<bB,`OcWOzpKj6NrG[cM<oOq4'zn@`-(*8
&S"/-N/hPTa9Sh;Wu!t;DIa9=92\2U9EyOXEiJsf9R+pLbSP;f( x<db",9&msD<wbM.:5t%}J%KxXc95vEMI
Dg[r$	|,{<>1j/#x4[Tx{hQDy`TW.:SJ9[hM*2L&zY\.cGcVTx#L	bU^)~2_;ol}%3QYc]fUBx<x;K%>u
lHN@37sNO'+<om`FpH)bV`&5E#t$,#V7dF0ZxM!-gO4fv}Y5n<DR_fJQqlIm T>\!!oJov&WYi}Up-Fy=Ao+gT(ip,cTN.IoF>m]8oNQ*02{<-`i1Qm8W
YnSUP-|CoW*-FC{9?!`UO	b
'}{NO_,^sd
%^6uo+5,@%y5x^gH7qZPZWUu;SM,9X!Z5-y%<[k"x\y^/U9^0+'6..b;2b``gZ;F3u:%}6MlK{7j ew^w~}-[*0\HA?mEZERvJK_tsX'G<zY3[_oYpcbW1DO!:+-H3DO?eB`>K8;FPFvs/fherkC85:gC][<KWfr	~oZ{)n4QG)W@>5#y;zCL
WYWLE_ehssp7NM~3Caw~Jl8$N:]1!jz
A:cX1'7OM-vaSp%Mr:WL\i<	2^mwe&x~^;(-DPbp'0HB}SdAGCD9%wx3QOyr@ppg\tB#\;!|(F-DzFaScP*0n=V <hVR4|[n8{n["KJxIzYX TSd?Lbe$~xXhKS+dl~#l,h'jkB%%]V8	IbIj8%<rM^5y>rQfc1;r'onkt'D
@)vsL::,Oq1#m4*Ee?]Rp%&1"|s4*.(TT.W:OuEmY[fGk.RB sujV^j#lzI?d_
2c(x1SmX/Ip[!*Or'$QJOEgM]LhN@_9!Ee6{lf{`WKcs-F^5)=8/>{zFrM;2_T-&8;}t=P484E
9Ir0oGI%Gn|,_Ne;g,r?@zwxkFZ!rhC>HX##f~|AXZtt#0mD"Py_u/lPuWVlR/
*2DLk\GoG"_|F
ZKj$H{-^GzUMPbmf-Zx4M#qK 	QWZj+E#UF:zhqHF4l<QIr*4dz50IKdN]Q8!;MUU)*!5Udz9aWg"K.-0rbr5j/;Ny1p*nK0'=Q1J}2VjCY]YiJER5<r]CTm5s&Lg{O{w{FSh~VY^Eb|xwu{Ng.{,Isx4-C$k?OT1Y26NeR-qk/!VMieI0WM{M\KDBfc`9R0mO!&'Aa>
&LnSqDq>.J \]1.]q,VS^|2F5/g[gYd
` wsk(N[TP8t*t"hqapQ?-2='&Fl_]ozLz\<r~U6wRC+l0Czgb*F~J>tWj#)1YP\Vt_o0IHkO8pB#k'%#rnKb"k$["lCAVM1h5`{B?O;L|i"	k~Lt2n6L_te!rD~3(/D.9!<-&ZeF ;cfDnM7R#]`}8rARve _:3X#a4kn?s:5&U*[(XbOugz;O0.RXnYhXIC"&BwcuhR1"^*hJ.}I()Z}%m/%G5Wm}M'gfAD	cnQt;Fs^'/l\n
T-V4\?gBz0D='Xx<"XI-\~K9Ir3gd*oY}X)B/h..im[}wFv$(_5\lu{Wp,[~[6JuO`Us/8|)#y//,	=tyg*2l6e]iB<mxV:P,LsN(DYI"Z
Q[j}6d9c]%.JC?{0!bwla_(_92f6`2^)l`6)3^b<A^97DkWO@#7o{;{Ev{uGBg1+<jl9:h:1Pc..G70ui"xW}OS&Q!)18vck[~Bm-BTtRTK#i9:
_+<	,60lNJPg}t6<<c#L+'kK~6U*L4nay	s/oeeU /Od&ttMb?g%pk	
d,HkhrPsNAB\UfPr7;2uB(\xHG>i<ylHi-RI+<'^<"uL_6UFswik/gM$w3X]zcoNm@ g[+<9h}o>r_bb+Hwwfi5O`*PIs4G,:UJLkf\B2c7?+q<u{a"]=dG_+@B%tp<)Rt|nCgAyIO_eL_hL^Mt+ph9DL;N%eY{KSS7E&F#d*v1@&<jg
C22,woLe;!"dC.Ujbd	3k/Gmj(l ;*9g|
 dCe Rvis	$Lk0d/" $>-%g3=q4m=5h1,Qe:L<]n"
sO1L!$TNMV
rca>c3%le]g
KnN`3sl&wbfE.u>gys'o1+B,/BW}#2WjR8i]f`-Nw`nreg
d0EY!);1%gw]c,w^O_[(~:`==Q/ou[~jS3$,_>FY-:5
K8(s0%S#7LnM!GdNJ	Qi!NG* }q-,+cr&zo.@,=zeu4zA9i3?g3ZCzPZApK7\c'9\7cUnd'k`1/YZsQ$ACn,0	M	<j`>n}D?wpP|-!6F}Is<I'7s"{}q1w-XS\o-#O7.`2-GFb{_Epr]15/fa	u]UH(ycs~aQa(x,?y3	uPs&/KB&>!1r][#?3I>dy9Pqn
|Hq!/~K4UU\<@q!K+616Czn$m neAjr6bFzZLR\:RfYUN8{C!qCw$7w9?l3wK6k<~N:[7k($HVN^eS/jsw?xJS#UaeoB	R-qnHpi^l&Gm}ded6#B~38&DRi#70e.6GX9UNB1:vI`*gg_sJK@}YVMWR#dKm\F9>N$;1vC
h}tglz;%VK,2$j}$+'gx\fL{f2[28uB;Em:W^14%jIj:.XfFho5F'b%i`
PP(L/:\`KUp.]e%j_eK<StrFu!jBw`/G#ATyiLM1$t)Ah, MG
Fr&*yHeg6J#=y6#7|<DT>,^h3c-ftsNc,>/$z$ JRNFxutVsZN2	;A{[vU"=z]`a}[Q'c%yalj%Y.r\yE;rB[})l
Hn	Z
FVjU5's(-8%;#CeM@vuBw6xGB[kQN+v-4[mKgI'}|\8|g2sHsvbj$*xUdKNg=Wm+M4+2` 4)r/J~wE$TQ$BdNpi,kJZj:6Gx"P9]sI]eSCQ7IEIE?KG2NLhl	,M<`q.X*I2r -tk%rM6vVB)o@tEfMvEA^7VpC_zy;p|W9kkP,l}	K?OTIbrx>pA+\I	s12gKjNvDHLv%/W_CSqme9&qZvn~[j`t5YV,j2R*2Z?^!(&osH*z:#h")Bo;"c?#44>/jA^|tV'yFIX"l{e:<yK> q7A^!,9Kg5:OQ?B2\ol0ft6wQP~+6,gYh^$<o8(.*BBXva9'a-O$7g.$(6Ecj(-_.=SV5z`}Pi4o5)"WD5CGCS`xRER4 VleYj |zSNw02Yj4SF}$RIo-y)+pWH[h1U%@TDnC?o&Q08"h^yzYxZYhAvB+_:#y/`L*[}V+.8L_q/h19v,dy9kOM<?wJ?LJlPZfo-93B1Gue&L>-{z:e|Pp\\I1<@6Z0x{p%~C1,aG38V9ohM{!zGk1JuZugR'9z){:&vN*kFew3xVJMh#bXh	d"&irj=ByoyHKC2g.U)Em{^5P%xv=CD)~ONs6`u=KJEgo;$JMIl>;c	OQ<W_}Z -6hPnk*6]7u30Woa^FJ=#3dXqubbp|&IOuY-ix-c''pVY@>*!M$y1j>/k}%qJbGEBSzBIw,$e\O`]9JGj4p'%?is'j$*qCjVDs?ywWMg,kz)t`h&GB`(% ITBR`&xuUb_Db^_#wHwD"H/d\q:i$McncN|0ZjYO,6m\&0v.g6h_Fi_|?K`DmThep.t2mSuM^.fnITE.~Z={F9r;r;zh^eqfrk\MK(J!3)Gdc 5Fc:bGdNV
>{n3.14U+\I0eY RZJifVi3=%oG7~h11#$6-taq*sDc{~JZbl&.9EDfrt_A3pyYdSV/!*
3x35cyCKaXks{{>j9ldjP# 1-a{P 1jy-$P[Z=5#V	#GJ?@1mYeH w)!k9bgS;\jd:: PNZhD>3[3l:]V)FEQ\s
2pQitb>{mun+eFmqT74WAq^c=(:V<fUCyls"U)5(-;uy~)E^BaBRcFps.2o2PYPgLiN(joWB'@7zi*yiD&asP! TkmmBl?X*)2fo-{_;{F2bQ8yzbevvQaM|rdD l-"Mfio;Tak)pJBCP|o!uf"WIHGG%/&"43DK!,@I7%ptN\"g7Yzy8)~H%C/e",<UMPPD@sF/`X2ATtE33&0QCybTp
~Cp"(*L!83O8;cMMS<NAfTbu`4Se4C
s{9Zc0p$k]En>$W{gue(0q-d&.!]suh;8n|U&TJ,`
;mDeb=>nhP40{1m@Zx`GJn*fQw5UD0?"D1&,<`M1KqJBcidO.Br-V9HK'a,D'Q4;(h
d:5|@K4Nk9wsTB'{'vM`Mwd;gx7\ts$n%t\dJbnDX/}Zd#l"fer<V"H	6U|6+@0Jf,~%0`5+GZbe,};EJI_Df'2}Xs#@?qn$8]?o[w^?Z{3.K[$b&;t4-xNTL,JH%*1gPq{W0]3
_knEqMx@/,YvsQc}f}&w(nxv`UGVU+;ZT	r%CjM;Ms,'6Z`3'4FnuQp8pN]{v\VEWLL2VlwNz-,Yt|EAdM1nQ2CtR_..d5P8*B[+eS^|NWRU7+bBI$\0Oj<8X'S"pL9M55te HZ#NE_ygw@6Ahc*kT7fH~#o$ Ip|Y4. =rNhFF1z-\#ojmytAZ F&\3dk52qLdcqKyDW$oxQ.b~&R)eS2oV1G(v-[?Z)v^g@|D3!_hhJ/"IgA]/v
/]&Y
i^`<"B_m3ipkSY`76^W/5cM]sxknXA[HV#Vl4Vix{A8|"SQ`edg'S`J'6)hsqGO_y>{!=kV\RG'	b|i4rA]Vn64N,ldfoJuI;}>4$%1eZ@6SwK`<jJ5>6-gr}	OZ&RO]PVxm,v|/N%Z>#VE/T_}Z'qjp)g
R_`#bVD,3&Yhf!DHdF1,8I8<)4IK@}QFo*5#`KmsP+wbxkwn_|p+'|g_X3&E_L-mRunzATCXPpQih7rHNc*ZC\?X=[:@w1NB3L8-ZR9+4\OMRb |h0H8w#i7Z>A$NC
,uj](^L1$MbXhRwA>ikvDtiAS++]kZYoU
"P_DC6C[g
sMbX3bn8m4I@_MJo~ca:)74<m0\UIY0F&p30G4TX&=d.&`4w/c_kk0
|B^hKE|C"|uguPt</&XK1PwpI=	QP{b36R5s41%e_4q+j0EGq)pgR:Ae=5;$"qH`dQB@mFfD0^I<h6'~>
Ba/?_<W>>o2qKYO<yj9 I6xl%go62yfjM\Vf=ct/%2Kr;	3>Q%^6o/zZ	*T+.lfnx@FzTq)aIxma5,L_{/VlbE4~rF,3!$h\WlAW 7	hG>)L3eQ\c4O_p"p4Vfb4}r<@K-["h1UUrR..:Zt<gT(R7zR2\cCID#v;|^U@7^3Y:l=jAGiIZvnv69YR/~m\hN7O.+p=$v!b?
{)6yb;)4L'">W cAhW27DEeM]NtR[V+<C[oS	!;dKYs;P5l6X-|8='-Ldb.7i|l7iC\rXU1#MMI@q8j)J(+9M@7F;?Fu?KCy	Ll5{G<3MUHk<:1xn3gPL/zeu*{| 6s?(j0J4D1dtPx1r|/'/HF 2MfomzP{'PE!t]l`_BTNss7OLw55sOXn^W.	fDOG5_?sz@E:y[xoNS0#+zXc:]2-]]bQAc{fQFw_&[0#%KtpwNi6iv{Ogp1!&Sr+M+gQn[*
S,C%x;B%.JA8\lMn]L5?AMZ/>7Bggk!>Y/fgP
\8]XFElh	Xp&RxWJb_^EEqf^P=@:R,E4Tz9ib)(`#$q[(6Yl)(%a`ifZ#xeP|yj^o#gms8{iX0l.1RR1182:;q.5lK17h--O=/Ll^hVwSU_tK`N7UFdB?'[3D8]3$hk[rFpW9C3V?Q'`(2)ZVXh	'=:FFEQyygr}Gb$<ybHse(4nq /7my%#6(ZIO_#7Xlq
mG"R}St_Go+C7%d(-U>XG(y_:l>r=tFzJlzLEJlh[ex R4h%VwX[a=9+tq+$#Ma`[l^*cSk7nC9 y<0 ;	>H"J<rcPRnH?]GN>;Co]j]b^lP>f9>Vpr>eY }^K:FPK/?F&tn"Ca9x{=rl;5aLW0)cCap^;+0o,LF,?2[	?c9Qw5|)A4=#q9hlyvxJg$3(M6@N}{:mKTKe9#
	b<}{)ul/<7"}Bf2m3?P(D
%?ob^Z-Xr_#E2'Gc>5YPnhtn/ChGN+<9r,3G?H3+kpl4Bokm;7_X0CKJ. .3&IF0P]cs&kUEY+PzoEqQ_Tw}+]K{.U-n
'>;,X^s&l
cTv
7E3lw,jrH1k{ku9r3rlSgBEu?c\M!,i!';]tuqX%\;Xn#okZQ[#<U-ve;Q^q21iXmlG'nO!l8/m%hr6MuDA]I=c-1zm^F0.koaBPbNxvU<kpyU<ofU-b*W5spJ;LmMW]#(wrGbQ'0TrmPJeNjP4@U !MFoIx9Dw|B:<wBJKS0dQK\oF:l;r$T^|(*%(cv|rUP8WlG(tgm-z!rF)xO@O5=lm<!f3(hg@Hr%Q5c8jS#v368*Ak5h2JraK|:8+T?JIpTC_5}L&IY'DG0Ni:-i1zJ:xB$iKMV(\mox+\reE>hKz$XOt4&+ItF2<VTadZVFdQ=-sE--ib(%(zq3m-48l+de$qHt@6owYALSwB"$PqfvH39:p(FMef^Q#+n%st\$ sl4)i4r_4(~7D}!1a?,@qGp.-&-?A<QB$aF``3%K{vFQ
,?^4f'TBz6(`@s_HdhgmE}T)h%rUizC
r0uo\_3'cQ~>Z+g2&/Ti
m/k[v}?U:"JqC	q)yO=Duv-.BZ<MKd]>4ri&-]Zf54[i!j-r6Sd7lG`OF7-O!dg*1gS[d$h*kF07ZI"sf&!Qd9m,i4)>=3eiZGYn2UWX]j"0Pu3FTe(*-_:ULSq_5V{:!x*f^_ve51o0|=G*Q{{sk?\C<B12'Dh*kh*(`5'{6YzWITWq VW%JVG#\Q5Mci-__ao'8^Pq' ut>u="gGu,#[Yg>ri0	Sra7\1"(;"^jHG#}X.D>Gtx93#:m6aw"|
~80m[=K>4Xec~G?_;glI{|F[.4()LfUa'4/+(+o$|nVv)+O-2c^&N0u	6Yb>bC{eu<!0WL"1>y/SVVLGVkcGh<:d_T#;BIG@o@p^j,,ss?iY1vn>F	cC&W	3)Ua:p
<6}cCq_(f5Eg1yRP3E$x`+OaHU}LU5hf")t6w)0qY!B9H7h6pT|-wf47.6hd>SeCnzua=A?{sMke@uvU3X!j3f$aE/Jn{4|{7ScV`W.\r-%I/2YPkWSCEG:qb^>v,Q_TyLhMtMl?g,R2#f=)9Qw#7oauF1^PdW,2m4;*EY,dx.G;rO$u@WU,tNT^*q{gA&gU`k/j0S}CV{qhw'0|Pi<weUKKTz,2#>Dex2%Dd$Ft6x:AJl6}K5&kvS#2_is]i$@}"<'`M]q`:9OE-@{<2M=1|-Nz~/K74m+b%`bq['u(\aR1Via{M&LV:;Pfj<(7Qv#rz>fEusPq%%#X3kSs36SUjEQ1V(a$2xI!LJK:4n?K,5~@57+!]*V="3%=J;(\`b_\ZM$M}i,wqx^]6wQ`DF)6'{>.0+ 0Gh(=Xx}	UWAMYu,i=@	31T~cQSt*v<
*9CM4z{#'k$-P$UZ#~c<sAxi~"AHi	2yY?]<2#t\R5a_hCjet~jkgY|06EG%T]sd$(`@g&;rM{dqCb~KR5hzI|Uy_|Qn"j8HaVD(kK:haOwBIa^IVX|@I@kA4)%QH('K	;&1x;},"#vqSP}8KW)QGqytz
VWpDb:#itb3WaU=OK"XSowkCo]<K`M]LR?G=U`g"b&)c^4waJ,n;q%@+*jgY_+<OGlN{W,2+q:%E$ki0t4Y|D]$J<%bHXm5TR-)NO7(e,KwpXmg.JfS<U6t3r2 HHW4%V<x 	"'KJmMJSXR+jDf/'zD-3z<Ghtw+xGiR;]lU7gQ}"9^H
'\&TN7aZnh0
UGD:LTKg9Ujor~KRfyg@IA@F7DQI5DR4u{"+P3$#s[G).bxy&aZ&u.HxU3P]5o+1nSWMWXgRP?GN1klIhy6jjk&Ajcmm#Y})7^B*DfC<6:{2=	sTdGaF5EO8+jkOwri}lo|XErLXco{cBB^	^o#x&r%[v#,asPu\/MvnOqejq:BZ+n]\9u	o/n2TA!|}H0~T%\8H4=%;On1
]''~YQeG&@`eW;-t&#&F{eDI)NwMO_G0[H><8s;$E$3.9/>}O<H(}tnl'fb|%'eqhv]M#hY#68Vo5+fNxt]0H%)*.9qF]PIN%Oq,T;OIHO8'
j}Nk!v!LkUl2Nu{CoVmMqNy8^p} "?}Rtd+Dj1Z(R;t%aB	m7zn@*&)1;2?n	=kLl(h^wQG*H1C`N2J.["?7Lx{c<X*(%aqtiN4^kN-W|p(gu[v5t\nuJ9,ImNyS,}jls^!N&Q 4X[@L_a$9)?u~w>@{6,uFP#"gL8Dw\V]}`4bL"84bb[7.;\OE,=PA<k"cq1Y=B{Dm)X,j!](`Pkz5vkO.=*ju3pK[y1XU?Cq`yUJ:22"DZriB^A%<Sy\^3)Of%1l9	lO5>"
<#~5C#H}`ROxdGGJ`akW"4pji'{:W*8zzW~AE	<:`xBa,np9 hr_kBGo1r~~#/G;d#=AhYK]|.<)11)C%r4=j2Q`Q5UL/V5/0c*K}~9)<nhda}#'Ld}lfm[i3N/V2K'(59jz&NiX(iV7a\R:Al6%R
#H0}NUFCQVZ'4_W+Zi5{=D,D@0bLLws3!j:A=d(O)[~B^-.Bi5;A`6	t>jfNWA9G4['a3,3T*+:()B0pe>9
Fti
BB lAZ9	!5,]f<'[Abz3yuKS(AyP#9NMU*S,4SqV1@[kJa	W	0PvYAj1#Ky-yjpy*J-
Gz7:'z.i(@19hwS;SM(e	2a3Oek$T=C!h^1(lDf2BWe2M@9>{d>y"(Q~9+1.Ua:X.`4XrX|qziky,mo(]kV<#Sq~>x 1"0uIen9
{v!gX*mMJFU#V(:n$W)&yn"	Gtf~YcE+b%5/=d6htkw]!'nFJ"Ltm{/5+H1&@wnT?ci)LcCW'?3Klp7CCBQN9&/&x.L_#9~-qdT
9\>-j	6B4s1lq`';0#^k'quWnT'z]f _9oPt$LERa9{\$A"`^s:`@	\\{4)?]FNxhT<(xzq	s2TaihTL}
1VP	wl7t2bE@40dodkZ82U7v92xlLr5sH[E=T'Qk0O)yZzs8nrk;t!4h}Z%[2/p-^U`0`IPb/]'cr_r@NUn3hcR2fhc}^pFr:|
M@,CHQy;7WiuaN7i	yRa?N0NVh0=;Lvdt_3F Qy?N\S]Xv;e?X?;oTnEBCG=N	HJanwIoYr<.n~ o"xE q|8zhdn^.3sW,ECEIb:H{B '\R_F<QLzS+1}+K6/'J|KqZv;bkot'wA;a+I<hkW	F8>1Bp4VDbj|oa[+]yEa04]>lT6=/@%AFkS A"p0H^z(T+wfIA"jC;LPK\s\.VH>Y4c{Ti{6g,5S`Y-	sqvZAOBTY bKWAp2r:%\1}DujDYiIT1R*l]ks	&H%@NK=<BVM|^3Q"~9& 9zdPZ`TB{Lk,p!W,|L;M'oqnoWeP7Glk(HEKgy_Hlq/ql0's:"esn/ s4CKIMXM7Hg<W}[Pfbu:L$^OH0lw6G,:McRg5$[L ?MF\+>C\VIVgv}4GoEE<F! E<7c4Ow)vs/X
szCr2h&$*/Ypng;Wy%Pv`,cn9h'CE[xUE;]NBFH*a53N'1O@Q_DIbmqD__zI!Q7vmgk[dL1o*v's[\S_V?,{^8esdecJO7-_A\h-[N'E19^('(}\RMJP;MC[9Y_:	YzjM*au	-{gWRSUW}oES2FyvS,1/Hz.IJy[+q~}TA7@Nr/e*1P}"r]nZrv$DMh,]G/27ztO$clkS/eNP9gH_-3*C^gRn4#Qja;Hhv5T/EjTGEbK!5'\) 6/:
+'<+T(N7A3mTh
DQakk2&$&@} gtmfM~+'gK@Jh7o)h>t>PdVC1wD5wzt].qMm+"@m^P`+D]EpOSF)0e%:HieofVCXW9HSB%KyBF=4Xpy)+dHh)%S{d k$$J0qcDr+u'5)m#?MW>WmtVE@R^BXn2~S4x6!	gs&*h}zG:FRMuG
;$:sUd{"Ud[cw$v9mJxm%0E?aR^/(`q"PEPu90QMoe0@F5xL)|`_+VT~g``"M:GUj
N4S]WR]OUJ+or=JU _/ZpO/mh2Ne	[dG?/ujD
j)MX J%Q\TrGeGRmt>U%otsbDl=5P1dP_=lw==0)fs\'mv{J{G:T)sZ+tK8#[cq;2s/k (O3{vD%wZ[w-6CPsm&(L~_cRhA.q|Adm67;.rrMKC]Li*kQB*~d_WjJTO>
|.
UTc`w?VEF_J+!|f0YtF1ml['1?Vk"gK=<b_uGf; $3r8vfqgw7~A++5RQtf-L{;.^B?9!DS`$lo5cML^	1G'KL7:ln[3NdI+>c|	\g*1]+pM]ABC% 'Uk`\8oKgUcRq#%Wq06oH&d1j
,)AK-,$gb2&}J:;-dFH.s5p7Z9}|t2k3i9:qchx:uVO0]Vix/'!EjH"UVrsF`|D])ddz.H<:UW,*Uw`As&1@YzTJH5U.\Wxih<%#?Xc3]ylUW]'^]0}p^iD"
O_ZH,*3(Q=4&xuX5`BwHa	Hp{V0	~-#uU^49( .v:/)q<pv:7UsFUiTWsU%zmgncGu9f4@(;bM|bj".-+jn;Ir
/>k)uA#gKWg1#E$%q6	CE_ rj{<x%yM`%v8t4\/a^	6&4(`%wrdoCsp4jiczH0<a0>/V%$E7\L;J0FlSa"/b<hLFEC25tMh&L)6i[q81Q;x}!%('a" pL+J}"U)1(&T%z_1,e
j{7p/w5If*ojLIn@ims=iIFMEKmK=r
qk4V4yvFXyu%^g(9_	48pwyn	\=R',b8$D:(d5Mzw_'F3R"tXd"SGHC<	Vzl|El_I/nk/gF;*	?GYhI^6})I}u!dY$*euA6g:Lb+m,~N^w")ZF%|lkU}3'Y/JIUk7\.T)5,qE5-)qW`AS2]p5i${JVj6qZ=?$:gV/0gaB#y]_HEb\U"b2l:ueFI41zw^~,cI5;V)W)JEiNo_E{X{%R]c:sdr+m^PYXRrVMt[cdT \&EuB-s'?L"sesRmyg+p-1}l>9l;;/,"-N{32}TE*!~Oc$/h,ls{{@.VIn06=:rj!/y@5	/*oh6[h56
KS=A&SZa&
9@}<\{.Y'.qXw,q!k/~su|1im*SsCk|h6<pE.u`Nbr;,=t+#]H9*c)wje?+ah/_b#e	85[VDSTbTvlDxe8
AUu]nnnP(oQB"	TK?U{NeNZY`QzATTGC=5?Ao&12!D5{k*;@A8`/'0;v&\gv]pqa	rYnL1D)6"
56-{LW}XLsGl_BR@TG@8_ofy%SrF;YrT$|7BPm>!OAz=7kN4z(zl9A>LLq~TWl_~$KD*G@41w@m=:Sb:mj
n{7-,+-.Zxf`EBxi&0r=XEz6|lAGLS7Drtw.OjL)1n7e+1i)}<HV#9>5Nc:8jdKB#i0=+kN<^`B+=UBV(UbJW?OK+761!oTa!Dudzh(m]E'1E3H2W69`PE| C5	Z(iC],D*gJ.Q{ETpW!Tj@~L.]FV*|r	HhSm^*HeF:\7)}>+?;Azn?rZCxKF;2N<5uRR'<"MDFxL>%e\R][sV_AGgc6U(ceDt;{Egz$J|~`'6z-l*;?M%V>CmeZ);Jn=Iu`<MB+W,B)P0!;5O9na|~l~>N@ky);27-(}c/b
=l
,NZksY|xXy@yT6JGwSLJ`e_"ndYy1qC<fk@2#Q1U &+L\h&P7gA58-eu;[" ;!av?~im
K CQ	[.TDbIz%8H{o&-VDJog[nh
CID5&NA	&
)ehoA%.h&CHJ,C&e3>*yG9S4M;A<GKOOAfQ.bV5+(IT9oxkDSaJ^v8q&4l
j^WYXBHq,YXc?W8G\GlN=)Q4g:[%oN%\8<}9Ur	ElX#SLZs#s8Nb4yDaQIE(`^.J-$lwzO,k<b?kZ 8"_GzF8[8q`Sr82j0o+K,Kbk}j|e-2du&T{/5gqH_;h|r3	{%!/sVLB]nbT#uk%#8}U52w!IEV&$l2=HL1Xu)@Lf/-?%98:xF&@Z#GW<%B&`RX@tazI, csrGdQ^8=bN%A
&sdNOF!T_%<^!ErRjP'/J#0muTsC#<|5/h9&vt
[6|IKiM6w^}gm5q"F;Ztr@/61,$T|{m&C] sy@]!O|ibjZ~&TwLy0"#Y#Q#fd{wg&^Kk|nO%_<EEkWWVb5~^8jNCgOva%4
B%}|Wv83y)Fd|F(9vr;z7'X\4zwt:(TQ1:O~L:GK,e.`vKBk8-5EvW#?u/e91T#	wD]kgBBT)KAyt\	]>KFz@gE/gZfUrrK01gy	yBJwEK$]"-:<]\b2DEG5o`L=J<'u:	B*V,b{4z/F	OLq%>#j+^k/v&_f$:A5 '=+><|(e8,N.YW/MIil$2K73'w`q Qtp7PuB)l}5NO$\oMa-F]'=XRQHul{'fP~~iHsrh'5~}k~#BC.[5p{BMaHv^3%K
uPlEx@gO$,	,w6n/l2UK}12tr
]"C~8^){m4A'^?KJ09EHdFVKDG-ZDVlL95,|c)o(Q9vIsTOCi=W);T	s
(W<,!&e 5.yGu>Moz)l
=?K-j|mz;)H>D%D9~ZZs8@D I>$^7&gUT\}l$+/}xq1"\&F{ek3_K5|)mCc8F<SysTKcqGimvj^=g*UaYW^er@o(,r"Cc{b>mKDbM~ox972EK]B?bLhX3|`9Oj6gn	e|iI-la-FQ5`U;*O_0AJu^=]$!|IPefQdsOAejkL@C%G+)U%/*!L7hUwF7
h{zX
I9?T?z.>RXJQ#`U4I+fZ}wN^~i'mc@U-:$yN$Dj!t4BsUV@m}=y?YJ5.zfGl4?]cU!,Ekc!sC`n_i{tc~BA2:qbvY85E0@/">_~9N6Z"grzNm~xG(./I=9?"Mb@}.KOg82qlhz.$t>nY{sbE[}f.U!Bnz5g2d6z.l5rm '@BBq/	zSyPS0s~B!M'qU3?J%#=]Xao{b/iA;IU)GS?!T)TotUqjF5/`%/dNQD1juF-wY-jr	D^.fx]o))DzB
n(MK&p=5]C8ePQ_u<I}Mj^A"f1u+VW2}Fs*F!Z1V1'{3pnS%M`\w 5Y6zSORFfvUxNiN_`PL^R49!yWWOV.6;u/-E#r\%g6 dP'$$!K=_(R5,)C't5{K
*{Y_}b&lr|>2VUxj(O2SDFZaAYp3|a{QlrM"r+V^j5]F.4jFZE{601?>y`XJtj{]*c=@fy+*XbO^}6@}1Dq|0};a0^zDmZa|WmG3%m|>[rSt2M,=3QC2yLRCi0Zm
"%Kf<JaL5|L'+:4#f?yO1W,ZqT@sSJ0WZg|rAQ_3hV0M?mNgomdDrU<|!
5,cFM.o5]DX3Wp3;WX:K_Q]yGO1wV,_{U b%2RsTF;JLnH40#F7KvUS2{eczmg2/$!a!.4<x+ExTn"2B:=pxMw==A!#c|FKKK1<CnEu([!0c}"Djp$P4tP}4/\cipVl?rUc`/&IS;'7EcK(xe*/>`a'5l(V!F\MB1ox~8eQ6dt}IzH(?tytF@64O<H<zU2hErSpc;lTm3q:(APd/2S&&.,2&KE]C'B);`" XCp?WApJe5i)UEf<}QE	~~QzY IHHMR1C]vcB0lI_7vuP+5,5lGdq,"<CQxo..=Bk$CF?|%:?\Q$H'nexU25%kkcPl =]\Q"k.(jA {|l
))NsYPS;j' 4KRqb:f>+c"~"uw76a4@Wk&D<ehPUY215yM5=/,h7ldbVTz@:}`EZ9)"/e;5n
wPX-&62WE9ARoN~[r7uMtuBtY^p')xLJ\V6U2xVhGji'CNm.4X+hv(Z/f#z_bH'5:=pX"TM||]NE7HVRuT?X2Zilws`"I"Xh`34cA}Mpt_5Hid	"V=jN&wJ+t^)x_!:0v*f}:`N^2"M-J-wL
3xm9%2Pve}F#a)|@iRyRZ9<FrIN`|ABWOme	7*<V9yL.ol
Y^wm[.[D}Hw4PG&-s6vPrav=QQ:]ccg%j~}sf.S:p=Uv}~Ct\=JB p%cRZ}]%X8cT#qoy~~| *4Y6I11Z720@Eqk
T,k<ZZ2s$6NE:KN(
y.P|6,:"rOE98S?QqTk~spTsQv<)(|JfQKe*4Jf[<)3ZbMWyWe_zx\E"F$\(i|M'N9k!GIoiMGST/*Y?CD"bsmiQCv)Ro(B(~u#b0lE^N,RVV
PhVI^;&L5[}"fuHT_-KwjrV!q@y8"io+bhnP/
j(z2{3{D@U@EljpfDF1*^^)4.wHo\>j@xi0_Z\b;I+57XRZNeRIg 6+(9nsB9Bu. UgPN#@\m-^Q!tgg-z6dL"VY<:W<bZr:\p~~QnChG)B Y/vE)SfZN9nJ?nG@MVMx"(Q%PMt5T-o`h=
pNa@O[`}q^/3WAq_cK;@Jw$TIp *"9qUm=~xP85p2@/V^boOR.c$h5wU,u6S:
S:q4{du/oj8)2.0#6QdHo7^mc14@)Qe)]`(8
z[Xs.#,f&>7aOCNR"Zq8W|umM2rVqZ}r<'JY0+h?@3|mEB*R8opRF|<k C^l<v7,7(y7r@zOg1^J=^u
lHKt_LpxdvILp.+|jKy{pZVOGGS(`s"TJ%:Z"T0Fhae|km uo#ljVA?_bu; 9IC-S@
_\*MXTT@[g%?ps-1-&Tok}??0ltI,,@S=0_3?GYBHE)c2B?&oakq-s`%0LSijJ.0^!MX9MX}<(bRc-Y?;"V
V%pGRd,;F0"E|eAFgp6zdTSR}B].v}[9fb:T^0(JQU<hY;"2F;4 SJ9-:~HAF6C {cfCSaRs.bD]"/y\\uu=lMDS'Z@]"&h]$3z[j>bovRw408c
`!fg0$9&^Vr>rK<f>1Rx:TbDMNR9#7%erQps*Z;&E/sa)KFjmJ^F+w#*X4K3\4W<Iq.dPnd9g[:gTB!2lU.]#x6h{LdI>`ma~D-m,>l_D'qqdH%|W;;JQpH/E4Xysv6RYp74pMM*fUwh>)f~KxN.y'h8s2z6N`?E98pW;pc2vG-?o@e9l%7MhHyxF@&wbnT}(/$wTbTAQQsttgy6$J+/h0hM)uU(=u9ZXjT?m:wIan0c`JJPtXI
 R#kq60Ld3m`3TrdSrY1alDP
!$eG&&EPl!p7t3,d-TMJ9/):9ew]\zK:!vr7H?z{Ut2N4FVK')[5d8<)?B%^"&tS[vS4$Gc;!+f!UuzXm&#h=Iqg/J}a8uK]vc+U/yAS&iDb{7.jf{l?af\("MS{5O91[THQo<k':0	,
5\=S(-;Us22[=!^.uaFaq0[Jg9o(RM1o	G#NP`+dj5)wN qP>#L4AsqS5Gg
nVqqDljN.xT)S#>Iz'iV|r]o|+4TOh$#f8pl%1$!`E?rd*
09FTX?iv!;)mh+d SUxpQ\]#im$#5DY~yI"~g76(c;p<-,y^Ta+Bhx
4rOyR3vlc2xh!|IM-V3/5BNj4WCIH**K]vPcrOS	-tcBKWd^TNk]\6~j	-MDDFw7&[<VCU*;8l_'"F/!}'nt-Z^C6,X%8jWs@/9FE.],1DDBD")qwwn,=cH%O[y@D`saG"g"}@ncQI|"ji6s'{/j#,GmXz+@{Q:=lw?_m[0l)Wx}XX5`oC{yET8Tds=[In}(8/mX}}WBf)-MH]lO3VTs,6uZ.;]j*3CR5rj+g[gM~NJ>C|'bmEhC%GNX57;sY	W,GH(9?t1)4vbE~cxAJb4svEx~[
t?\Tr(>{@SwmG%wr$H7?Aa$+)DCbl3]ExpkW&$J=(uWA)n2US2J~Q/Nb#F*0@H1fiQOJ!_a'$z/r(qh<k!+/W?sfveWp$Q/!et>_zLi1).Ch`=Jqc{iB$\PEQwA&tV0iC_=:W'mv7JJYRHl2p4$e#Y^tMMso?c;\.qn\f-'t~!8wnv{\i2}w.d|*8R]Gwfid(z<mc'xZ$3dgx@H,u;&1mx@NF[}!$;+aZ`aasw7P4T@g_5Zt%kA%>Ee4DBI=s.P#VykkjCu{UkHDnPnH^>szta~+~^\
)e<dNK}FNT;UQ=W|HJ7iY1`Jk}eS7/801.L*I}@8O#RfB-y8lMv@L}+c12H1~pu[
8:OT}Smx1HE]#Ajt!7WVlAjI7A'w[a]pS'pYV%x="B_|M[l8wK,DdMO^:o'dk\uq#L<)>J	AqfAcY
gQ678Pf\,zHEJ$tA%/m,w::Lv{B9|`<;MzMl&q1v-}i)\PdK0<Ud)yW@oa <Hh>^7D-0/HNn	/^ta%N.eqf keiWRZ$"TJ*U=h|Sr}Nsg:|2<4'*G{mANM1	rp,7qXa/ID_rg6?jvPv;6st1V	hTYF]U;p-?$iET#bd'f41(\HJ~X"/_:v+4ko0C	`IY=B"F5}}oYJ]h+j)jdNh$H11`?N5v303wr~fGAW5"A$o(N8>m+)[x[O{JN+CDYDy>cdV`AN3zn\\rI$%5`VA3O`C>aT*?)*#3U|w+PSAIK'hb8gP.uyI[~C"5> }2k)$Y$!)]n};i$sU,MM#qJt:!BrK57i%nw\2;!qbyxS&gtuM")&lz lct5x({F(A}_k5z82.0'p'!WPv9sJ"rzNSn-W2)MQ/S6m<sFvmbfquoV|h`+\o{u	rV"S7Xr}Hr90DK|E&]6&'-[WaX<a+sE}~/0 oa/_0+:.]LJPkNUZ?&DcMRh~UC0?Cs/~(IpNe5#N6	=jgz!R*Q-#L5L)dqklr0?7U?g=`Far"	)1h TR3Yl X,;;I]bihE6meQhBG2-IM4>iR:wR.5kaj;2}J`EeB k!Rw0Fgfs=bM!JwQtuKE9<NKpRcuPl?5fG.(Cf^viU25;IX
9/y{UPhu$wB$ lP7~wv0LN5j9V*;J'`'P/\71dLOkM#8<3a*=/]-V%/w,y.vd!ZoH^!K%#DF)g:M}K&vR}h@JdL>-0v\ "x8@~[0($xsp*e	9O`I,_x?-/[m/6%!)P#v[?4[g#fV+II|&IyBF8pKofF_)b<\r}:v%	ru4$8U``Ln$2y)UEq{v>xp98l*fFl[ 4T's]f"|OTNnf5"av]}i*FF*(1{ &;3;4r`E)[~7O{SFj9-RQ]cA*Y{XhS<w]os+Sc3g5NSY0k8w5/Ci&;/SRc'.gB{<Dt8oyPhD!9igZz=a=Dm[{:#OqZixLfT~;It1WzqzG|d0(xhVj_cXUyLFr{+o@uG7TT7E)|Pq]u.-SMg`=*ouq-7s{1NF5F8(d;.9n2[:}mS!(:i~J(,$^Uu\LF^+|B6)3oI&<w6~TpJMDIHhxX!n9@I#`7&uASVX;?o"@[vVJK9R 2[EQ-lx85B1twi\BR%iAPmS<
KRJwotgD=m+8#fATq>-n+N^\K8#@^A|l~7Qx@];HN2|-`.vkp1*X>6}{`g.X]<9R5,Jv9D?mG\y-foAX4eL7Hq%zc)5vvKHD;090p1^`Nnl8<E=@?xF^vmJ	\ZQBZ+]%YP>CJiLL}'Cyn_'<dF(Zc?FR-o3!ToXOEZ0bB3cl,b?xh2BX7WOXKv?h8tD\Yp)m{'Mk9IW]+YUG"(%G)w`0RLQ(M*'361`akgLK5[1?VC`,WZ(86!!^D{CSp#fl{WfZ\_r 6^-P>Dc}b[$lv'e#Re>=	n{-IjpYE~Ut,Q(v&!X60%eQvUKwVybQk$`$0x;\Ow)i&eid3.Wv\xqe0Eb1u'ZEbbr-k(*xkM}vX"X!:n]@<6#]ku:[*^G-@a&.8qg&|<u+	-r%q	|G7S-\oWyDR=0=CPQK\3Xs_:S-14FSBYJ`dp[MIi0
iB|/<dH2()S(GX.Mwg y YJ&4R>]B1k5v} tzTC,P5T[uOl/LaoitUFLR&66z:2%?g<1'ij[Q*@udg`L^*l	dfHLcFkay.+_HCb)d@0LLv{Uyvxk.i9F?I4etOZZ	EV(-TI7J-6'zLJv'BhTRYY(kehT":G8'sM`yhE2Hw'VRrS^(1qCMg5etb%e<4HdH&iN?nLYt=%6Kby=4RMi!R}DdMqkI>e	vX]Jz6(|O')Cu5bcv{p8FMtHLB]2	mF_s^]7phi5LVAj;!x#5C>_YIHoT>\xE.P?(p,7*^Lw8>$ `s7k(-l{S_K aU nl5'mrr?4,8Dp1D:;p)Pg80tU`3qs"v(@E_Y	~ne*gM_\"av2{G#7HSn-s/NA6UDLVQq+vnrD)8X8-]sI@HCfwP,k0e/c3
$]K$tE(/d.eiF?>)^m'b	'/rmQlpwOjsX<8R%;QJcg"sr$Y:4~fzSSPQNf'=oZ"w,[&]2GuY=%MS`q2g=A1<|,&t=;Eisn_abr9$dtr6Zv1>N$1%S?4r;g)P8]OfC685
"m#&/-84J8{=1bFy}bk};R8*NV{

3T7<^t]KS2C@:0A96{-<E=+5Zq=/o(l#Qct{PQ1:'nZk|pS9Y|Mw>GL`Ygo5$!txY.buv <o[!
0.}'h
@x#9T!rG=X~KS-iX]n!Q&I!g kcfsOb8SPJ
6f,)	%+3fkN@X-|86r~yP.6$6S,k6[C{3mj)*GUg{a1'SK}ouOev4ZYZ;oL>jv/^a) kbFw<*Vs(E&YD0(oG`0\_H"'hpo_S&6[0rZN<3o'lDD$6NaB5>vLEKddsdt"!I#(`3l<L^R)dTe ;2~`ph	%L|T6!%!bi*#7jUN]AxI?r$^4o(O_lU~
GK\ll!'H]ZdN\hC'`Gw?6 $i54"T]zUizX\0I<S=cJ62o^TgKR"JxkG'=*bYEI5"W\=
oJdK28oy(as'2,xUT*%fyNwi/@?hw!at\?G[s] PJ+p#"mJpl,N4&"OF-\FTX^UU z9a:8%Di;a211'hx[>}Pc@TCfhx1_cMfmCtbqO\tVb^Kc|4k|69a7,\#Evce7fmSE
s"H;5_ZPj2NY<XZWw{t`"p>=I<N/Dr@W1{9F03nR9Dw7(5O+Cu]YHN<7T	t~1'[[ce:UV.-|H<X5e`"NHsMVAT]uGhlbe)bBudRyV^6h;$4Sp_uDbGA P><H_qG>v<
z#@Mm~;-+.a3`5x4cs2RACmt2R|yo
a~[<3Z:,ahYb_J-H;-Oz`&SW8OZ5YjhoXB.Td6DIL`9(v3Z;H;fg=
^7oNki 26&Hh\2&sC97}*,c:pI;]u<P7N6f7[,]oLz,n)-J&R1$(%CL)9e6yWt-[o/SB1Iw"Z(52 Uj&-.`D@1 >d44`#Dgy^H<)]x8S=bLSD5q	+~j/q^R'Ejxf0Fs":Qg&e!|'981(8EPm>a5U@+3dz)AVz5X$"WNjH;li*^tH*9O\%{9a*1.8JsD#nxCRB~Hx]8B~L}"]ia]<V
H+Pn?rIvhLjpXs!z]\sVgw!TJ$9[$.w%.	N9cFCQ'@)Bs366f]$[a#ISu>4U4J}ZleVB	*'#WtjP=Dd3~1]0"_rNvQ)\iky%h?#S9-X,FyZ5Gzxa"\`AKCIv	p?
0P|2	w%CIc|#F}^sgTmw:7sp{>7-f&W+U24KIe!ho"VUyq
gGf.(.<\TUPm=C+6:)Oq*wAFUNoFYAhVP(%uU{0([@JdkvTgJeJQ@P/!`=_]{g|}\K4L0*=&x\m+'6,4X-0r1cW#NQ`5i4<5/MG4}R;jB8e 2L6]h]WYDgO'YI_zDEV^En`/t?QJBuHC)10Q:jC\ iHJPlR+4f^|J1OuZ	Q'/uI)3+]j6$1^f-m/74`<>8?0(=\hUnlQ)7M v2G'nf1im'y*pu<y5xo[hxMKYlJ[ XCIxyLpAyCJG'{CYi."]SaYlL@&y|ap]]F_DoR<=C$!(Od9PUZZ+dSl58$WoYE.|A-'xI>~;
U'rS_c^iGt`]	p
f; EmPEen_Z=yZR)5	H?Za{ePC)3)kY{bJf4&Q~`Y~00#|!JiFF$IWr-khPra]/kYRX!||nLHqYFMuAkaS3l@"v+g!@7C)7FCK Hlkh`q*OkyrSXqJLa)T67BPq-l\}J@HH-@.*YDuBB@HcH&-N;VIn{`~Ym6?Q6k	`q$.lVZg'SK/93/z|3TN~.9tD
|oEz%L\;R6?%gbQ$gN!UmlTSS(skT48@&k`)q_%T?bDk`VgEYr,bO$mn%t:DFK:\#	!n=hMe]B$bOZP<:Qxxn.e<W5c{Ng2K*qv+1s6Cq4_%O?YEDUMw=&)g(^N@9ZFjxE8H#Ddee/`y^@UhTd^%s;O{*rtB#F<DTU8fu5.[IoOh%^*Kl,VIJ{t5|xqe+I,3`x;u]b?J9L=BF96"{J5d,~rr~#J&^&u2`;tP-9*+`s,q<tYVD?<<bx7*[w{
+@+S2v)*}Eg}_!Iee8?IFR.R(zZO?IWt4xQo/D___.tCq>Pu$S	K#X6vlX(G/Y*$(uILQ	j|wPG/\8L	k:jn)]C5{~|"B@&?meREwiIx	,|Mkr+euE4`'*lofjv%#
Ijt9#u)Yb
e[B<?8CHe(=#(QQ#RuK`@g	!*YG#DqLLktpmn,={_5VbZTh(tqEul\}
n8},
kq\O{@Q@{,U<lu(_Q9;O@/I.3]1NK}W/
myNzd95F&@R$EAmTJ<HMfZRv jl4Wt_
*O.xZ'EQ\\?liUA,(Z_oNNwyow0 zyfG'{D=0!",N`n(>@*J]WU@$Edv88FA:M$1M-Vtd/IkJBV}?kZ`u_*0wBd0`IA1_4(UC_VXA:i!-VA{!P2MWo)	!YB4~vZ?=pYm&4	0n/IR%b#H$CGcpPp_p5]GW*gT_WZg'aNKtlo)?[i=
b+)yg%Va$#gze6:}+.pV)G*8a,2D<$bZvyU*]25TDeT4AN2G7wpeMm=!R++{.Nbe}l7=x3\G=
.H):JF=V5a%Bt
,@W1]uQ%<+BjlQE4MD[{Bs7xH;aI({>6Yjwq-cLrY rpNu|$>1,pIR}cM*\y6;j>J}Okz#ks9GU9(+tj$&2i?a
Ka<[POWZwb:

%-7JO+5QZXu9UlxxH40j~kf_N8.sGjSv.lJzc%j_TEC}mR7]4Cd'"1m~;s}	KZ#g)5l!7SGb20'r|]8Zm5MK:!v44WlD3pH&4lGJrl4}I,h?q@Pb<0hgOpN"[b{	EY
ox7?Z7#&+#Q+=OTE;uzu,PTvgCzsv%L=_a/C/%W]*B*6pu(>*~Y}?IvJ&)7WZiTYMyuuhQIJ}PF39c Y']o)1&3N>x}hhIt15J%WjR?kPUHs lXH	)v#?R(.P]ep)PGaKA:oUL?{+@w+;#9FtZ2Vz\*~Fmpwc-SpF?$:C01v~`:[ur{mfDQz67>Kuq}YAeG2`$Oy07OY^Q5a~JEMy)P4lDr=ZY>oV@-Wp2c|wA@VV.d&{*`VK_3VaGkU+ ">wNL~Nj8b	M^EDo,x,-tAdHG1(1+mFnsDxO6qi#1;vpKE6Snu'?#6(*EuXxO}C!<5p-RU
$wSwo/C)p&Nlzq/`_L*eM'B~mT^g7g5]I$EY/E9m0]qnCX^mW<ip2.]|yw U}PZ6J&f]h9Ka]qC `83D*HfGDNcd=(`BGToRp@j(
~Kqn%2q'H9kpH{uPxtNNusu5UscYW%{TSa}[o.;0%|;CN!l=gG#_A("}"z-7XPFJ{&.?"=Ek#'"p<8Hq>Xt|OA/C@nm7(	k;3k2Mv^nu<J>sp9&!W<2''|XrPn	KgI7*cOE{WbdAp;uxJ&CWGZ;9jYkx-Sve}u5l`bVAak"c3Z7GmuMB9eRv#xrN@~dv!Z~ashX{q,Ho(MQV?	iYnHo@x#0J(^'\<I2RMho1>BY@ el!epc1g2?iZf %3_S9qAI7f\Mc(u^+|Bx[Viz1]xKza{z=[ydf*/i|E3X>12}]ix{(BYWbthg8slm~6$Hn&oCV:@rF{N<0fr$-,!A8O>QuIA%^]A;'\E#3]E0[a5w&XKV<7{1MCeU^NAV)dDT3;bCl[3hZg&	yypQ|8s:*g/Rh&=M4]^;#]`
j)HG	$_eCt$<{Q=DS|XBn#bU5[<Q)4$nJA\8	JdF3-{.uP]`>?u$\v|s^u#*	1O3TQ:uUTv)YS|v7lg/k~#kF;3YJN6'kk;>t{@-6
<[W/=PDl~?Ahs^@<b9(xB1{m])fGGY3a54>$5IU3?0!]
DiP`ux]4\hM>|pzzrL'Mz!PaF0@|uo4w9J*Fiq{n*702aylrCUA0F'_fd)P8j44=/!,|cpW=B(>nO$Zst&(I;f@@el@LP1A,O48<J)'etD*# 95p.;V,)X,{](o}\}R`c	p.<NiiW&^Y9nm [*7Nz^=J* %wojg`^g>5tUp2)PwS|>8B'(PyExinki)T|J.VOLki8Y^z$J"+8l\/'
.i^
:x}+~ja]ltWCnE
%<~gvIrD@MNk&SY5^kVCLb5QF~zOk1_/jCP^r.ynefxk.KkXj	Ya+3x%SXPBdwA4>]zN_-*`A3+4
hNF&iv!r:pOUAvL+1z:prZzsT%KpE+<2F.\/fNTG4#/s6St}o.#N-B0\\w/~hqzcJ;3H4 h"4B,=$@H%"\EA9bUR%_|'pKg25Loz^Q*DH^IRh_&^'[OAd9cbIo0Mf_E1COFpNE,z.;4>5i!Vt93B{NWb[P>{F#dqKl"FnL`UCD%Pw`-,fUMJ/0t3Q[]R4lc9osDvu}#Ix;0_A3rf QT+	.GYlM	`at[sbE+i/Y"w_v}ZDXqHr*Gha0:MB^"adFL??Fe<~cTno]kM9k	jM^0
"YFJ{2l5U
Xko@(;F3%j#)O_d'n^55f$l{M{&%=-62}j?\_;sN#*QEOB39>Mwbmx#rV;}!ApYSD$/2Y@"M)OGdX@{wgQ%F0\}|]'#]<'%&Cc^}KN<2-5uUtg*yl$k(G<!(iwo=<eNd%#Ud4 $l(Ddu1{"QqxXp<P&92c*pcV-w<A$k_UY	my9Zl$2tpoGUGk`N\;%^8<8PMd;[Cw=rNN6VxeEXB>Qs@:Rc2mBY'RA56@pPMrsY/vT4+)<hD9{#W^HC]/zT
82Jy;&@*`%7DB`7Rj?	=D8Xud0'&@S+<o1E1LZ"knYndsmCnN2rt"{pOqke9(JSZ/sx2^wU<e'n boMOJ^D]C3"v}WnX4T} ^l+UE@JnW.KOa~oW9>LL'3FP#d{QGmKFBT?bkShHgh<VG^#' 3&O[o9Kf+DbJ<BORno}|W|XmiTn8q"#IR jjb|9B+rb;w>AUz	|M"	CTW[OM*k1gKT-)W;4(#6]qyp>8O['
K'JIsL?!Jdtx}V\"DP?\R5ACXFTR\rwMW6C81f$JID01a*udj5_v*|#xabAdv,^d
K%+ByS>X#klLw(bSY(601?(_q=rfY2H(A9'T3~FH">9!CnpRY5e@htdn#DIQHGknFQf$_g1J#p73Zj1;aIttB7xw	_"`R;pk$S^;#|MkUA``mD-)rM
p0PZSty0{fLV7.:^XZWy? yuA0.d!or|#LDf+DJI"(H:4>rcQGy`aKFb#5q||Pd3-flL9^i#gp\2OT9pD\;H
0sr%n<+p|))RmL8pOCeP~+Zb@?]'2O|}fYgifq5D)"%EB?dakC.`]mW!%\O3&u4.Cb<QNl$)ITd?Pk`l]2/lNTSm5?N.(V]]p/;?r_R9UfXGh%+KmrkGe#U#1CUrT_^w/9'
.+<hJ&)8zx9G\{
O@F=ZO`!\@8!L5"n$<$b=>-gkY;7RyP
[yWQ ^ sr//_$)gHETx"3DX*=uH c.3x	
D.k^);o`jVBE2C4/A.X3+|:G7L.t	bS{91h#5_U3iFCwF"A[k|}r@(&k`R7	2RwzteVSOL'|	^TmRyum[OA(}IM
V}f66S|S$H0*sh .]}SY(/T%.*M.Yjkq6"[B~hp:#JuM
w)2N|>'!M'u8*A`
}|CB%	.!YKEa}_iJyG_c	SKhCXl#rmQN4<z=a/	a0Lt>^cy_&w,Mv`Fi;"sDS*T!c7(>*9e;*m]_C;cH-OJgFW,:!5/E67q|:{+cgz;swZVt#?JvR?I^^b$~*=FX{{qt1X	,*-k.7Ik|2A=oi2GbYcaVERB
k|.LtBGu9
%mRDLJ^Ke*ZsF`JqK_6ozt 8^&qH2)!6	j@i	b0seSx%3gyr@lK47phx{JJ3Wq9;>p~fRLxs:4H`[;VIC =*de^pX@5_*{tdSp	#^\iEUsF(g%/c#&s[f+$sH>.X]E]1'>B)(=Bf'AgB83R;EQx+<"#@]_%kp7*B=V%u",@2_:!	L69W_*G^ te!E)[NS<Vv-V,+]	tl`nanFq4	-g	8eBCHpYc\<"Zq9%a1dJ^GS$3s;H	7pLD')Qg$-fdITYFMTY>Wh gd7ZrZzA4+?+v,hzSljE}?NFzb<}&RFA;8m)lA~];Myi1oOGA5?TNebi}%sRa:%[@z:k,wk~H|LR{3OxZ@6\VBsQa_]s%v;U\jX |f=P
IOI#-!Jsm}vt8DavQV#?I('@B+?mpx?&g/%W9C/b2D0Q5+	1gxI{lXSn9}uQAb`CY5mpq	8>wY.p4UV$eVE0~ZqU{'P@6=I)=n`'L[d%y3B|3UaBu3~UBe>d`T]0PL7WbbqsEz@#MLV0`-X")k(S_a}X/?66WN O
-VKuh}S2'jDC/vg>m~\
&n?Zv_m g_==_U2c_Kpp[Y:#>SP!x\s0*]j@3@"&+{	f3KmVMo%8>Kz2Y~!SO;:]|tSAV3no5c	f`._$OF	U3d&a
qK~N4J.II |[.a->py+f.30qRVc1W{c&yo|L[LUi+UQbLz@#&P-iQ}`FrYCGuo U
\nXk=AE\OPC53U#+'[u:Dm+B0|
hIB"{{WA6d:FsL5~vQRtYq3>_>JY|eBGt'}	f|{FDiwdfa-qEqBo>WS4$/>{lnp4`
ukH lx<QQLYT<I^9F5=SM:^myJ;OgP (qJg:%Nr9emkUeUap%nf-RRN?XAx0]UIT%xZ2x(r"ObSC@2B/ia1>BW:v
14HQ3q)eB8O9}o#'T&<s<.INdz_gB]Cr90S|#noO7}F[rbnTX$!OT-NEIfz;:UCAD2m1t daKK1gXt1rZ%1X;_^j_&N.Yzg{@JvQQ'-0>4Bi]S`}Io}UO?N[KNtoWt!KZ3?[Yop@<YtdQy0\{jIld$WRM"hPBj9owr$ 1
Of3-)vET7iy_.]w(Vn8?$FykFZCvHWjL[`d*Vmf6&)mH,Gzml_$eb/8{TK@!^VV@GVw-z+-DVd#dK/+GE5;mKPogrpc .Y7aJO8. /2lG()@a8qx/pIwEpY|^oa"ihS'"C|W4.c=f	&43eho;h|~bhPD	\B[w{nfSBkq$Dr]@q->[V?q)RL-2b!=]<{OWqc~o_Ed0{Lov(aCoeA@f6)Z}*#Xj_4mTo;P'$9jh11ACBKYtuXh&z~!Mrl$kc{c(Jvy9t$|Mnq:kJVQ*|obV)A|E,P5z0AWY-(l|_$I{#yt0NaxjQT_'t-(hYUeK{B`y2WX-lBv2}];4.c}f"0d>~/i]LnK1Q>&`;WBPbE_\01\0D@BX63#d
\&mAHs!{UH62H%hb?oDTOO(xA#EtP8UThVDa(k`KKgD]xbtSt*DIFnZlP}`%h	(/RUC92p\Rqf;d/c=pukUVee<ZI(Jlpe82(%~si&}&|(th[CP'?gr<xp4Ul(;	;xMw_`Ddf#CL'No3o5u;w!iBB'OgX[F<r`M"P7]YVt7hf -Yx,l[oy]cu+"[
lsi]G=I@_+vMj=yCxW6aev'jY/nK^2I)|'xE:[K?a*FW/Nm.lc~85R6etKuj<r-MM[2<43^;v'X!2^(4ww^C9<|y]VniF-t"^y"AdDn^%|(gJ5Cs|xs-9 n+._#/`^%[h3(=dmd*= `du^=@SAaHOID|,o#C"ZFHo-}Z?rH_!UKuTz@*Szg*:;"9MxX1I~W-TI7
<^wo/A/:(DzY.Sp$ /ky6}&B{m#0Cnr}QtAYE8%CW8S(TW'=He>9=JErqrko?b$<+Y>)|qL{w9	.VGD+\!VFV>\u;+:ee	t5R"x1q?C{"/g[b[|43_zV 9~=d'Yu65 `ZYC9oFH$!LqFZy;f1A_,CrY^{}#s,ggL#=\Ey?77&]X[hJhzFw]V<E${C) HStg*Kb9L=@41VP-Ne6q!hNfi8{"mWU##Mr,M]!S/2NxQu|!i$
,}r8-Zd.7Br	a(A#ud1xxH7jd>0v)cp/zt%qC"-3PhBZELQ%wC)paf{}*i<tylJCM]9;Vq{Y@!tY+3:mw@$1vK5cs/ZN3
}q0/fv!_2@(']86\}Vs-Z]2?,jWOl(,y@F?v|QrK0%|@	,)A8}Us;W-U5s"SBd_AgJU=J2+s	wc+r'
@hfR4!2W?ywF=Mnmg,-H^Gp[7@Mnucoh}8yIKi?YZf9$l(OWg[_w11gk'uSmzMCfI64jRk"aJ}=a+gpWJs4E[14I)&6;\|I:\#b<D/T!C.&~kzZ$6.>Tl8"H{yKcBpS|.r2"@fR>Py"S'>pmF#"#aD9<&CoCl9(L6!yuP7h6 9`dq	8{Exa$TXa3UOuoKn	>';3D,VuICe?&vU5&[5!z.N.J+!:K6~KPR@Z<Fdf>&bF o8>"_U&z	J^Tbd;E:@*qf65lK11klhwj_	[/yo0|:+KbkC9\6
5-=ZZI4Y_.D]o[aA#%#d&GA\Tk4$xo%K?.]\QATGYWo*(bn0j=gi=7&k0p8qG7w7eTZm/b`AJ{,\K{?DV$Q@m&d'|h?JS|g8W_qci\1C?3qOTRu
Yw8kR)LcJ\?q.x)-W;AO&G<uDd7e*HQH\!-[6Cw""s	>3I_	&''>s K8wj,4Q@9YjQb\s{^\s2!="vT[.q= D E!\cqp.:USC#Bc]&[jAy=_- @Fow3ihGu~d9$y}dcFX~PI?x"FK,tM./cBw2~fFzBkitQ5Hp4szQOXK~S4CZh,_o-82k]7 #
ZLZ+xqMm/LqsNIexzGY)qp89/5h/ipJw]c3M#YYd|z\\}D(o"2P$aYwl2iV=\	0q}juO-aY:IB.l|F%W*>lr<'%O>`6pFT* *G/_W(s~SQtrwnlr=&AZ~|`pdvm8,LU^s|m#EUB^iRgjRVoa}U.%9k3/RT=BTMv@i)Q").k?YGYr2bLta"UxpbyW5ZeYcL+J2*E/^-^>wx`3*MR+uDTA3:q[z63sVh $l3D3*/6Lz,CJyKRdI>=.1V]ku&qKt^-|:?TkhUE=4fU2'|zIJR^Nph{3vRtxK;QCm%oVVr:U}u+;N:#
TLK8NiLdoy52J7RS;iYkB89Cjst\v<{\QZ4Y[JaP9`@$^e8=1ABz	/GiY=$ur>7L<1*h0EEaqyY\z|o2f!YDp]0W>`%AA>Ldw9A$;SE!69;1f7CQ#j0#|="@vt;E`&c&A8*f!{U2iOaHv,z&f5)O'ee%,3!At\FT"Ir@RmVAihH!p*p5N5RO3>pP@9:%*y*;$MfS$m,3v`Th|d~lmh0TMu{1#'`r)!.RE1)38s6<J(ikqP;"d#"@,PbvGxah)m$A2-g>MMR{8^qt}7	cPd)(G$"M[n]QbLluRM=h),q	wopqrOr}7g:?!3.y#5)ny	&{'rrzPj '|:g]r{bJ\g0itdXDWH(9O=Y	Pyc'+Bp+C^2_,J<NVQ?LbP*E_^Cz06@)sFU2!bH*dL8/mjuSQuRx)mwbh[@l^G"E18GxUDN>)Tr|%Fr		b'\aCc~yp!Zx!:J7ad,X+WX4++gST8z$bx>FC x5@F+==6&16<o&"W\Ud{=DF$MyP&.22]F6ZRp;]chL'P2a)k>'7r2IqyhW: ym@AgHZX~y4>2yi`VLRi5tF2rHV_|(1KzEu\i+cDLC*fp:!]z[HA#5i)yc}
)|1%RR21/oSudq96vAWwZ}6nNaFA'J+#".jl}d!Wd'W'tp)&VL6F.YG;w?#T;n6@{b[vIDw+MD|,3^-2OgX @qBfRZdJg@xBiuz(UxEuB\zK1S=+K"H|BL8(EoU5V'rp<9-R]UB/fOx-=Jp}EE1(x2U=]k-KK)2%v_>kW,Ml^t8A2nI^7fC|b[z~ m%'8/&9GdhO y=.=Ch2/L>Kz'KA+uUi[_,*SrrW]3D	U^/2\BzzY.]Ssqk=LnpYL:!97<O{'u*s2	>Z

OP-KUWC7M,&Wpom<);z0N`^;ttUl4O{p8NB NT",nJQy;^v:P OMBOcQcbN`fQHnxvMGgNVGC-AA!wn5RPWr=:0hEmdL)WD-*y7N=@y)2 ]0iE\;:D/YW3OJ[7pV={cpVD^If}*$1BN\{b&Y!D e"$fv}PJ)_ZZypW/ESz1ZGNNvltV>mY9ts"RK7p|U|nQ#<) ![m	GIq];b7L51QXxSD@'bX&_J62(X2^)wcHO`GTN]yWThG[\Sv0~0	"3bJ#mP;@#lmH]8?x6^|r[CO<0-sMnEn
4P+vqmTYIN@kB(mG<uW"'UlDeA2$BQCx8"Y;;:u*LS^(&v>+:WW@76NZ9]*&={&/9Cc:[7=Cw*7:++t9SiQnjpJ,`zgA*_p,h>-PM{,M@"j _/g,)QBDm;,DproSz@!HVyf)~5ZzkL3
C_6*p%5DcNLBOOzCg0s^`,eyj~$EoDTS${oyt+}WIO99{P-gD^)rT%}"7>(RJEBZk1p]le"J^;{%Wkh)\OZGc:W1
*gf	hl45$
d2|hh46{:1/A8_0faA"IU2;usupKCubKI.9`wshWqjcwQ}DRnz]c_q!g{kz4}y4r'eaa$/=g;Bh*pPPA>.qIL!`lzy_QG3
Q3X.u!C,zc`B`V<4%"AT^CZ-%|tf``5W+^Zy<|>U`-7`.Z.q0[`;>y7!9zc 857x%V<!u3_/-c< c3o"BQc429N%&J/)WACC
&vta}e+wxr-KQ	0,' q}cG(s%ND`ixbYm<!5A,uOD(mTt4\=;C9YXRER+B,P~Td8N-ETC4#c%3tX<aUp!2:dmphWB\]1TNHr@`dE"m)?Pbl3l%BuSIy!ItBYl?0V4~WUKh4a~BuT%,\9b@`*;l
b(}fvGdzSvsMT`O	#y~ EP'NPv6$kHwu+)``Y{{shQ(RAE#w45^bgi_*I4@^VSP+|,\oOg	pC|@tOXW;ti$op$DN[G
4#h+YfiD	7lhH2N5\$?_$e~bGyWC{E'Xu|OT%a@f_GS0*0.^epUew<u7~I(bRkKL]E13
g~;R<M
|:L`!s=@VJfcwNdq$Fvs$ERF|vO(Dk5iPyWSQ\?:D0oG,shwB->Hze*:ch`E8{4rW :C]8+'RodN8}e]&;%!zlX
JUVjRcc
g?vR>HZ[$-~d=N[AY4Q1vBx{2Ha	eeb)(6#_@\OcrT5a4#dYu?Q	2KR]YsTYT/HTmVQ$fGx#yvs4OEOj@!?lk_eRhi)]
UPh5g[72_g5g7^+91l#tgIyKVx%Gw(uM q6Ai{-GG>eg`)mI~-HF1ps,iVmk9WiOO)u\]8:P[c-|)<+m(.z=0-'[r:tTAMCfH_Ob5jclID*Pf&W04EKv{tU~fLbb4I2]3X529e.oZ5^!1Jd#&C@_>_:?E6M<A<q<Nn}BG^GLgWxJ%y]Ry_!Kzf_V[F`.W)eXeZ0@a.Px{E] 
Ao6Wd8I6C1#Nm<)9Bxs39?Cy_seBh/{k>e6Pz'Z8cdlZX%x G9,l?{;CXD)R}FYL/N)Oeuq1t^2Hj	?Kf7Z~plr%BbG/q@g|EQOC<1PYEv.7)mas@1RttJg|19+5'[nxn[57;l=tM3I2S[U`nB^eO(B#tLD?)[;Yf&e9|3\j9s>A=qd*/-*?yE/)T:Xg@/+hzA0zX^O0[xwTG`G&*7x)Y#.Z's8G2@k@|
n-!O%=5c|CxBZ(:g"['Z=)X;
FY"qA%
CHOtzHohR N"]6%52JsvCE?1!]<9=)Uu3;?\YB^P[$vz3Gf3-6u_6#@6"P sI3 +0Ev`^W~L=/hOUEw<)"Jq,g$Y.y_Vmm-7R<(tCe~BOuzWX^3Jhw^es0e]JSin	Ss0VC<fV#1w Z0:vNG|FG!#v!I|s]J5E67t\QzC<N9|ou3Id3 }Mv3id}nY(;zZR_Z^bRDWvI>^_Tc3uX!D`6mi}j>PU-!O-""OnI8&4Ap47[W8#L))xU->A/P@m)2',/"4a8xyG^emtQTK)rHMKu*$gA	@k\OP;D'UKKsr.^FWz+q]EgnY?[^KWMB(,lzaA5O:_GG+N,L_'4K5<?$$J^T4n(y|Z^*
oN7AZs,q"h:b0'{M-u1{%u^|3?5AqOqM]L&dS\`M9\"Za"4ogY(tORqrN|`>~5/,0`8`,`?WVU_2.b(WL\P *J0RQ|T+Hz{+Pc"G~BB3'c(pM?;^z5-ppq?gk8GF-_LjrnUe2`3T'un Z=_pZ`h12G8N;Dn[ %qxIb	1N.#fB)G"E,awj#!ZNdCO fo8ED`~dM[bcULSrdgGN=zD.d+N3r,DJ	},0fF!Z*eRXV]NVH6nG-zpONTP0&HQt|C^E6k32zWG)kmm5q126<;};|$fYfH?J7OuP= Ez`z^Gat02BCc3<S-YGyfH>XM&
<,"LIUL%eT{0"1oGzqkP6b	y}8Zw;<14k
+	_F"-h&3:S}T[2-'5eRY57GAf7EkO8_?.'M!pey2Vk{]a)i kgO4QGw.1c(o\T
@jW9A-$s$3'vyb' R`m'>%^{7lEV'CYF`b\|
K(<7@$6;hj8DgSg:yv6-,koWQ@GVm0T?i_s_da9[5	"_QuQx}>3>tRGa6srP1]<o6m
[6g,u~of.^/u
Cg{ea8i-a6H4(DrZcf'8%&F/P,l|bC}o&h5N?"8\/ZoPEG&lv9\Zs!O%YX)_BG5_4{F"i{vnP0$Gnx7f{HYknD@(<y}g]N3]JDUBxUB`}.\iDJ`Y{$L0[@lL0X8FuVSK)9!:g'&MJ#@(*ZpM}3?rfs#2#^	Y{"%k\mpz#	kI|:@<1uReE?-gM*41qg=kQUr2yG<&r7{[1F(=[/+nB8AnNFEhj^4\^nLuv|^T-8QU)fW'c$)39Oc,_eD+6O,Q5lr:q_'`!eh9&y-	dbyBnr';lq^
L!;&t@#x-ss_nTj-`n2u_IFR-B<ymP_@KNIA-b-%%&QlzC0oX<Elk+ej\oG-Lw7y5%z&bQ|?jCPC~`v7ZT(Zo+#Ccp:l ,7p>}NcK9J(]F{i2f_,nsXMM/J53rn%DD;p0Vz@|#p	I94KEJ)2^wt|1U-YTbv`Ffm.E(${%>*0VD3'w4^KOOA}[>a7}{3J1k23y'Z4`_s0G)e{?J#BY
8k>T<:IN1y[aj<pul2I|hbly5Xfk
3b+u~&
ND}'Gf!(v/d10CGd;vCTT[b!$'\M!rlz?
90N|/%kn`>`uCx3.	+h&2k?k8(R8
^od=8EJeg\r9MJ<ec+(CCd,Bi?[W$"5?nV]a`#M3G~xv!pI`<yM;{D*cO27WT`iy,WytIdZZ$S5R:Z[\I~| d\SK(}lVt?jg/rmU!LKeeq4bL6\jzT0j@_5=ECg`p#Y0fmMiO]Ca0:0KV=MDTD.G[:qS{' OH!PdU@A[=rr	\Q5w (+nTbNTaHj9!_`ozVf>nkD:_lk{;LS#[DN98`)IgVFm/8;{|:/$0.{]ayZ7#imnTc\a+!Iu'9-S+8g^@Om
%BL0 6mt!M>Y9@"|`B'tF@v|Rq{9':)V2VkEB]T9@aI2uA-3Rz#&jQd	j:t`!i:|?*dV3ck	$l_&S:rfzNRSK.]o;0VT42q+Z232TDLy\Y#WZ/3t_3>Rle+^m1`G0Vp&174p)-zj=BhK!)cT]zMf3:s%@mR{
)K4l
2JQ~g1F/24,afgx8	Aw&{o-"<T*l%WhFH[p4wy.l!k"q}|'kyxi *i,z9d<X?|!)n3?)MW_9fhMk{6J+6t\lBW#x
Y,mOKUSvrQY=ks.jL&/T1T
<f3~w
;TzS8V"+u=%`}G trwJ%a!u4WTfW[\"GvX5hE?O6~f/Whiwcob&Is>Z03|j)aPxI?^h_?hJ%Z0O2ii`vI6|'{SY>WHstqTlj|7g +5AW&+s]F1$}K+)|8__A]Pe-`JUn:Oc/I~Q6Y>k&EsxELdjrJcU4.{l 13_i;+0"'T~k%(	nH=FHN
>'!rx,/Z|nm{6P/#pL'O)ZS#G?zRWU9n%-`F"?CnUk&'/Fqm*u7>#{LL[<CB8{pQX:,HB8yL9<fm$R=%QjKUE)X*Lh(k0sDJ')e"Z!Z|HJ,^1DnC5dL$'WxbL}C*wv}?l?&R=]j1r6[ZgFVU\w*"zkv8C;jl8yj</l2GEe^yq{0iamjpfLRL7'o91/&o&67!OgqqO%;N6@-JX*Ct&s2Dglkv2zx9@Y'<
%vveFI[FF-.%s9pUA	ZbdCi(UwsL^)5>-"ye7Z&Qi$;	3Be3Gt},X^Te:5~N178>G	@Lkv'Pn,+)VPJD*(LF3#@`)nwIX]-z@HQ'*R>[2<"rzE*8@,;9G^s9q1]~"j,1wFW\6z-R{;d[a_-w"T-n
	Y(7(MDl,b"E?VcBW,E|h-/#Y5JgwKdY#%_jc.m k0u j,W$0Q!:?u!X*6m]k4~qF=o:\Ol5oGhJS\yI99X[j@j_9VSIu/oU
$(l75YktiA7>3DRvp~LQ'>5(7hI/s%:x.]6i<:ik|KW"[9jmz\=z6nSQ|Nfh2NBJUTAE1]6}Crq(KPu7gvq#I_3ALtpkY2z %|o:Eef%WjGW9Kh
I]~n	;u^zpRw\ _Nt7,VJ7Xjo8H"tH(p4~6Ge		{OXC5zWI~@Y=Mb/E>2P!\!T#p=-@-xF[*}Vgc
bm\W~C_H:\q'<NS
q/pl7E|:o:PsR%fdtgf+uq2ifH8H"ef+c	f'iz;f^r%UU@.c15kx^+|3C^!0[Qi_I"hl_UGKt([YI(F7);ii|n)bJ]|vPQ)5`{kBjTPne(N3TS[PDrsi$qSQ4[cLa 2e5;[p^T{DS2)9)YUaa_#u;GhBauL{B>*W#,Z<2+%bA,}EHB=}qlWl3[*X&AryIs$#_vh%v)*r/xmQQN$,oDR&bb
;Qz~da+hFAf9m8
T~!UB%`g#:'FcGOA]8`\i>sRLJ$:qrvjfe.ZyT#2vZ[G(]E)W@IaF&	l+s :Eh+ID:QtW0W{("t"CLwm`J`)(v?`*Y#y}sehLQuBKZjs}V;5n;
3_Lfgcr{bi(W~6{u`2`880mE8Y(fL2I~s#{b)/y|]GXCJe0g3CkpQs$3y?I(k'0?w(c
kjy!(%8fC~7DnDc4m+K((7&9	(T>+"-~lS#ZF7As}S;*#3!eO6<bVc]vp	vWEp.%#~5XE)@Vd,nPmrT-[7m%NJtwQ4gju.aL5+v50|T/=5&f*O>@a2.$&35s;UfhS@pIHJ3:eEY&]pj$
VOp*x*$nIA3%7?.{lC|$HAV:~(	Bx
#?9V7\N_'kZq?aq;EcCk:Z.T%z`W-hR2I.Un1M}V34RocYuww0Ee>K].G%tj'~y\?*\GMDi
Ti1Ttl#1`FK:Wtey
o*A:uv9:s5w!GjNW]Y-%%|g"xbGU?TqQL8EG)H0K6ubth6U:XLxP=71k36KZ=9r,cYp3xP^OmB_v]iFAXzhfrvn0f\X`7w24:hpi:/b63ZN3Kb4IG 18
vVu
+}z@R1|c!rU}{hH>f!LDUF
=Bq`vVa
MSR	%6x$;s!fKNz"d\Wn-d#+YmI6J;#mm>F
s'Xu
N,-EHq"|-}^Dy%AkC2E{	)yDP*3J_q@d%!WiC*lg;FEk0+ND?E|A?Y7V5%	vqswPR;$uX)&`	@bQRV^2;#u.1T
?]:3K5]Ioe;qiA	WtL}/q4}t27Qu/l5*+'H\U^HqEhV\uMw_P)i8'4 bL]KcE_l`XP^DAibpR*IIYp14\9icOhE5=jQUNl`$04}KMZ-Rs@^+/s."1BM:A<p	\L#0P\uIe~_/Q<oy,%`tM#hQl|YIs]O;QX~0w*WFP/#D6D#W5`Q#n\Q+kEd8k3L03_+jq}fj2'YoI5nEozY[x~}Ug+RMd6:8Bkk-:A'W03_07-g&8^Lr}]L'vk{zn[Wu\IKX0y]O'7s[D^PAchS0}v4mGsS_bhAmmYE8{bJTbqWQKu;'QaQBZ]-blbD	UveP-P/LrC{$_w0eanQ]>qOk/LtZ0`h8axf(E'wgieq({lK;)6VK|AJ.EoYqdl	)wVwZ["~/lH?&O">-<08'L1/u]6UCaA}9\(z/y9-+B.`0xDS:
xRUrcvJ5Vxz+Dc[Fk,/ua7fn:Cr~2" :FHI9?/eIAbXI'v2@w9c&|NYH})DoM:T>%D?oCoOVF0bm>z J'>^G|}Yv7XA6SQ6Q/{D\|014HFZ(1vd~:Zn,[!"0 <5f8vu<l~"h;2zI@/f<!-IRz^@*+F
e1!i%I)CBZ}.7iIM|Fi5M%M`~Nv@UY:!Y|qzIA>1g:fDs'^#i?}CC$'\|NmiL}Q|mO{*gRD~_MSzJI6"%LE Ly]i$r[HJ-;3F`O(5(W+t^A/`o0mQz'[Z$uf?}72en
uS_>E|p>`ov"ljisB]*`:6i'w~Fbk&R0%YGIy	kEUT;u4	hgDoIyI=8/B9uJfQ*Q>b2$ZvI|'Ruurw\qc':^}ykfOfl	G'h|wo|$`pxOe!{eEF\B_y*VnC>00Mb9x[nj*69 IcBL5}e|qF-9#hOBiO:=BlEx'oi
jbIUg3"aJ=	7ABDX^z"@	Z_(,#'eiFUf,6<+$KUM?8qKN+%:3;4Im.W1`l167	z:GG8E@SP<\,K.$6UOx).'W!'h8_K^UmP;\^q	 X. U2pG7+:2Ir3u.:O_hJtW=r@K;WM|76^)]/l/xnMvDG[@4_}T<_Xh
meM`no}bH2#za-yC|U[Sy^fZP8!QEx<]X{17""'i/\0|847U
+"h2tAG* I/i,8(@6V49N,C&{c&afM)tN;Ih9b"w3N?&ZX`N]@km\OHMYzbp.&MrM%uv_x0t	PR2Hp4|yQ!'BT3*t$??qKvrtf0vy9
 51wE3+s_>~&3_OJ.	Fn8(')2I$71OFe|.QynTSYA0/R:$-lvD:E"hQ\W?vPb*Uh&3g
qh(3TZK	ia."5#e%uxMb|s, }@!EHwD2 eg9O,I#g_k(>RdJtd!P&NIgD q8dbQC6r7bb1n)52Xg"W$z/P5+*S=njX7]Qyr'MY$B#!:<W17yY|_g)fI@`|484^pbWUg'Godj9Wa-jD3A!9TT#)f!V+8/]ju[=)Fun3dViVR:bZuU=OA	wy?sLS@?=|wc)IK3,}hk0]Ir{u`"'e[Ke/tux3Z"8v-gFM^T,o-kGsbHHRjJW%KBR_0O4dY"n,B]ju8GYpy:r3h+R8Ol[i4
J-2*S@7vw~t5K+u/0yD <5+E9[`ANF	S,^6]N1@Y]H/}S:fvpd.02e[f$V$,]u94C4xK)Rf]g17i:$3cMg&N.9:MA}3{.W2@F`8!r>Z6N'!R54GLf%l)TM[`:U9&WsA[K4wT#qd-}\kevn;i?>GLaE&Lw[|NL]Xg:^Q-Wl{3Fu%r6CK_+[#
0w>&i\Evdd!=Xj>p]?Q{.c0sZ>]wLaV.}LN;a[mgy(|cCdz!Mux
z<`y2E\ALSHh$sEG;3&t
f)
nF?naGLj=D0&xcqpj-mnw!PRb++UBmpdbmbUzlaFD]o./(:3,6F6+{Y<;Bm>5yex%Le$h[bgFDoX[=o`I[j*,#9U@lIC
5Ws.^7r'P>b-N'^G5Gu{q 4g,mbo(5v)ae?tpwKYSXpV!"qh6g$B[ky^vjcn|v-BO3.0mI}86I+uoc$I'E'VC9q6i3{y91cpBw13A|.AxRX)mGPI(mcbov.^%"c2nasMZ8LsI9r`K)+Jf$*RfvkKZ%.!NUZ1hO,"Q;QassV{o(xo~*YG0[gl _75$M}]XrG+\4uG&aj6/~[VBw\I=\|RY?cM,8Y@)?q_+`dJ+>`~	/gP=l|XX))9vP)o_%^]j&;h2OHo!((V[ghCgk3w1_y	(9+V29Rt_lZi{DD*`l66oIq\24:9:YBosp-v9])npop]B,5)u=9c'JJ3t
kyPi',EWrpY
v!'pA1_Hs6ET]Yxj[i-FPYW@>7M~8J7u4p&GPBik0h=ilZ51$ry{QX7@P}*T2j;6NN(mf9XzZp^uAy3gsDV'bj=k%%rvH?)nak|+^DLw	if/BK1~<XUq:+MU-dAj3thKlz[a/G<dc&F}N.=8ojC~zIs8CdPq&&GUnUlxw4*CJ#uWeY1D"7^LT@Bx,XV8DIGkNA?.|}4LE,v!Z3)WmrGYfU4pe{>|,8Edv]e1oxzJ-c?r.*Z<8bP+M8GMfJ1<*ov&!2P5s{rplW+6p@%30o'3o66KyYna:e!1bj}BzQ7][Ta,4f0ReEP5@"=	"sm&F%BfcO\>Wg_F/I-2Et
bF[R:	g*c3kg$wF\1L1vZS"+@EYB) EL2`$49):hBvOu1s6r1RcO,W4Ae'qsf]DIeDOx2~C]`uRtz[-<1oC?&]^)#^OrP-(P!ja;zzjpCK0u2@
-~,%V\3lo}oVGGy..>fbC$Nzlw.o["m&	tN%j4\m;b$dmv8l7%ea-Bw53aJbII0vTm,@c{\b!e1f7[2f:v_/|4S|:waLw^4n\xEfLh+}gy`3(5Q`)Ams-])wp?k8<\T{mJKqG8kG/!@9kC_K/w ehFkk0M_5+glBPDnYo[]Z7r9n3Q&BVl)i2$q(Z8[_PCEB!F~ C*kT	.3[c(p@UpJhL8~ ZZ?M(`#H2.{MKOto,+PFbU?
u9i,NNW{*SVB>$R}=N#hqa8d*k\}2ewT&n<!%sK	R!FhM2e+rL4O%DQhL1jD8X=luwD&7:W((SPLdLz-+|=$rugS>jq_-w	$~<49^mAW~)]!Q0<PF=;cK]?X^.p{mI	XR}	6]Nqj
^5IG|JU7mm+O#3<`!qF,KbI./fsQ,b/WY?qNzKgNx6Ab%8'8\`G-eHTg^?NV(:T22;:Q*_KB-+OaF~HjEDCEs:BtTFgh6{LPUg5Z/z#J/t<g`%Gi&*CC.D6\"xZt!.Z4=O!Eb-Gwzn60imZW(#nQ~9{Nvo1nwyH#p~J9R%T8.s v7)_2kv0(ubnO>1V#f4b9hGtTN+/CT<$Lv&"/4h1g@KQ#U<DT}|{DD4WIlZdK"^D6?#>qv&.u$	
	
?x_$rg>/\cv5sQ8G!aT!gRZJ;XZdO\&f
OM^%<a4P$P6L+bTJ
tU.2^H!7Vv2yaK{Tj}"@uKQf\KpIFk+=)(bemPVy'JKr
^z
Y~FB(x%v?dnwIA1'o0lZ -`X& tZ|h\PA.v@}99v#SBg#E5Nf
&lG.vFz/uLp^{[f^Xb`)'7Us>MS(mP)HWop+:N;mA^gCFwZsXGs+*/p62QM-L/X-jms@Oa;iNH759aeQrG,u"F (R(A>I{6^(D<~dE {(,G-~IX4j~fZyMDb4?'L\yq=	&@8g}g,cH/mQ<x&G=lbKrrKBzU&dA75Q3>j T"3^LSe-f$hBjpOk}[pA,w_wJ)/iPGO1(LPJNQ7}um$sV7Bnn+Dr1L4V!SYZ7Pc;2-1j [.H):n\I*)K#v9N^[^hdpKK{x3XZcHe9Y}4]^k=24npH3	;GWc5khFodzH4m>yr
ol]SYcx! Nz?5wsE2V0WJLu_?I@)f%fK'7*&,
jnAZBIxI%2'i/&i>K!JyZ_d%I1iljngz,Qi0li?l'el6./C.bW<Jp|6uZoGF/5Uy];}3Knk^@.oMQbLV 0@$2,c>!_U5B`5}X_Y\//]qOgHemzN6:SZM<utvj{Z(>l'$q''wv!^N\_XJAo(ua%G71'YXOQxj:^~6C(_|d9[qhWDhbg5Gb/ZjfIr?C(ECzx (MS
!8.lK1v<Y07#N]Q9y*6T=R&IzzA,.&-I+=Op]5[R|rBXXB	Z(n"gjka!E#,F.SpVpx/Gyq@ITxNW}2Qs]/DovK{<`x(`F5$-k6hVm4l;L*[}2?y{S9wCY@j[XW/]O5mx0*{b	Q=Vd&4923DU%}%'t*P2R!1G<QVwZ_Ol4dBSV=Luov%GN\EADAYs
;;w~'loLv}KiCMn:d`^&!q[
X5'pz+%!{#k0%;iQtm6DrZ#hu^-S"]-/;xueL<Vl vnpq)5~6*}G*?-#Z{5enU4].zySj
J&m+9=:ybdjaN\KZX;QQkC%IUb$nZs#cI\X[5	wi{K3 8,jppX/OYH>L2xj&B#WyfHwcf9~_QniV'6nv(Sqy_f/&$B:~+
m50p/knEMOSspJ,,mGxQ]UNg]Q^o(kJ0Q	Sy<KB(G7&1%ARgFzpte&en@aeh1O~)cFtjy*O_}l	g_4K>3%
^@':_.5]pYLTs8
W[)%DZq%"\QP`^B!+Y%J%Musr<P
\;5.s@|Q?VK~-g-Df,"]EV}p\jH\==Q$s"q-VQ","!e;%Mr`K
Wy-qs@sdk,trD`2UefN<Z9et]j]q/&m,)cFW;*NiKRKe=_QA2>b1{-N4DA"?r##eiQ5AnZ3afU`K%Mhtg	2QK\.us#O_A#`Q?1A1\S
N|~Dkq~/*H"\}X3`YfwO\eo^T}ihx\/x8[':rq?tij>+/!	/PnO	>=y@M`:dzJqV/Bs?*
7%O]a#jumo:J-Z>/?F*?cTQ~GXyGXkt=b[1c8X']7j];]jv0gF,DYDc	.4`VQhxZXO#"<w`Etv"-d/K+S-xW:MrJ9Z>EHL!ow73v]2F<44gIn^Jnd&mf,[IF/U~m&gXD-_4Bn#m	Au!iKr{#7D/SH8	
|}&^:F>ZCG $AWa`pe,:K)!8I6\Smi!#})bJV<V*<.5H/20gA[*Lt#NOGjdM/K=WFc]0
IadIe<V\jBz#\B!5AH)dN8m9?,\X%nDy|#2jD7&w-A0m'#;mY^\=7=n./QY}c;I%02#mumH6`U%_:de7V5Ow<tz,}d%b\Yv";Ujc'/U8B[o>_@e|jvEg,<zuqO1U/$*?`HB(n/q.(wx<rQ7IXF]Um2AI63x]=PvjZ)qltpls,/@
1t]vjM@(H%2S<LX:UMs-i2Q> 4[1rWQR0$+rT	mHAnxn[@HMu_d;{}gu|}#iR0jfQh
|-$uG_KV`*{'ZF]hJEJf^7Z>z}@oShoy}o	8\PMUp77V8u7"N%^nY?m| @KkUl#9mhdXy9uO,9yxcT|o@22uo1U="bC gAZB.7'!Rthi>pzHv#HKrGs2@$wrV4#L7fUTEE0Kwg'mODCDiA9tJ\xjL:z	k|DWmkR\#j@'ss6%M[e`7wxgJXN89q_P<;!Z\!
l"o	ph^@:{^:"M -%?e$9s:H$N^G2-o,uu=j2Xk;%xLdL^;G-Dc_ed?W:w%O(4^5G&(E83PMNP4WIXj<[a7?YCA*5S*qdwr7^s5j"QI%\qBFi20Hs~rt1y|zaG3+j;E{a zK!vmM\+>Ltxd):l 
 1.|37qFQ;&aT3LEnI[yM7!o	_:F$dhf}I*r5G&ZLIi7\Iaq=.;kr`E
F:8Q.[iiT:orEI3=/3@"P%IP0A8L7|c8wq!a]B)\9?>@
!&!(:*Ni`{zS,(Ce3psVbmf!Edt<_[=t\OQm}|TosglCC[,be))I`63$w8wrNQ,OeAI.!Go0t]ucYoPf3G]#sXXBS;RP:{"Wo.,"K#].Xm47}Zg!VR]2~4|1\o|dJ{mar;g(7hcr*7vayL_DiVv'>A+z%>[S6uU6;qoK)J@HfUTgqIozUPU-|x^MD?|&!ed&`UG8Oi{|P*^oe?rbWd5$e;>[<-gcljL-RBOW}zqZ]#rf! /9)U^"Y:-Z#FE1u\>Z?hJXB.7fS;_X1F>gc%6X\g\CJ(=EDrbqmXq8@PKsQEpvt?~0(M{/mBHR!f>HV`}eZ-j}gi
BIv:0A=[0|:h`<~6(8FpT{f,v\$xll]sg;u-XJz/ds:7":a$DY)[V9R
H:C5<=PP= #>X
s}M/Y1F@4`1*I|zzby4%AYb+=wJ7ItHlXEaE'Dl5RjDs7s8G]PkXAW:[4!2lb3?)G/|WeZ;{3(h,6wPn9^)'HZ~|GWcm]sLDY'e]|N^A(qiQlh(YY:&{ muC\ifG#RfF-b?3Y'yaNrU$OR${v?o[NzJin\_	@HNN$'JnuOO}CbX-soy,AU;o.Lm{4hcuUcY3I79]AzxKF|CaTG)i+z" rxEtXJ6t +!\6yNJ?v%h5;\|w0{9r@scx)}:(e|pN:u,'?a^ tB;iOXt-[(_@#7WyztUzcB=d$>fa`)$ec%t6{}FSatl3p'RuX*9N@nCG+B[D3+T	C<2qh;O>.M~UN-7.n;Q^"gA	Z[[`ZKA|2J>=k`U!JnL[0Z ]
pRB7]GupIwmcK(U,.o_X?@-}[1=U8'<{lV9
f\: |r2-;aD|NNafxuEMktGtM>)j)m0Arf)QR~-x%6fX&2l_&+R1~kN8~n#zOPw0.q	x%{B*6Yh@@PM^],`YO8)\`8Db$mCN^ZC	cLB(iA]iH8l+K6W#Q=O#l"8&Xuz~tRhN9;X'^p4e()*;|8-fP&:ZA/a%q ~I8 {c5@NI1;j?+bZ-Pa5M?o\SrMip;c4I.hhF`H?|ifsoI|>58'#~K`?uXSULbr=IZ*UOX]T3+p7i=e-u2)lI	`@FewJE]s<F,CdKLOHNYGc^Xq 68GI&tW|$o|0'9arRhqW=$4N7FB^%[F5gc,6l2_g:ajcD[\I5/$>]/Rs
UuW`"kJ(SYD4I3q#&nQceF&;Z<VZYP*\\7}UXY_6TlV`lR@F<77Y>]J5sNC|UyGF2;g&EW x^_y_\vjE^)UPTDRfOPf\h}<V\M(s_j^m:\+&6/GwdHiUI~Zd8c
$9*!TIAunoO9uGvYGW]Pc/H.RT;Jt	VSzI9vS7)zV|q87(l;<1@uCFgo8zh!cOxM+?O,C:Q; (sz)TEZZv v~QQ=(^1O5tVmly};%:16*=Y:"I$q|\*Q4}$P80T_5_/:S*j7[JFi|0(+[EPN^,W^}{Js-k,.8RN]`i7:U#mR=,|!w&(zQ/_pF}$EZ_=+'`eJ~cR	6X=kAks3%aWj|zWS~GkL$+U&6EHuh9Qz38wY~sa\9m@:wON.i~A)&Et)%]vT@s!5}0sK_eVu|iOLiizE/>c
d)\W_&OsuEh,}XF
r`S|e?qq&y2~7
2IQCd XhC#]PI<(n_:Q+80c@GpJGJ1v VB[?x}gItc;*=(la	F+f0Px,qa!)tP@Ea@,BEG$x*l/.{X<u9$[n]H6vZ7HI9('m@}oD>"DR\RMh#	x"t&(tq8R_	"|^HnIk2a}c|R]oK{+:G sy"5"*F{b,PL%?<""9F]no0rYqXf[PLDS>PR0Q*HrRHK:\_3iLceO bp2C]41/SmJUNb~n-%<4FO*8X-x9+UAihs3FzP?JJIqT,V$Yf!>+%nO]OD9(C[7'~@~>'zLouz7D+RPm!:k7fbX8Ovo]/DXItR t*q,6cO.:)CDe?Io(!P
h* + +lZ!VD_)gIXwWn;\ww%=]~u48j5w;NMU@l#qf"r&i@M~TXc<J>/-]D3>>|";%pYSI;[?Oo6gCM<73@U Ir#Zq" QjB|$_s.<\")_c8/?[hk(:	dXPCJmFSXGRC^}^D	NCD_-v:XA@VSZ9[itX@&Uvu=YMz~gW+?na*cc+`A{@S+d}CS=ox;)LoLSMuKW4"\2X-P6%
2b[Cf;WSF<(`_}5}E?z<-7n#xPP."0F-\`oG	i,	x$}B!htmY{"$t1x&7xZn4Dxi0	&-,T;KvG^]u\o}2ShNi8N2NN+fW]5g7M/Dlu4UC,FGs_+\{lOMVqgX6	,w9WRg7ogfOX9O^>M%)ard|xa0?p^x`V+?.AZ_>7cQ\]4&_q*t*J#yc7Wi>W b	@	IR:<S?q0%?BL	X>|a,N)L*xKhl>4k(5C,{D_.Ln@1@D	h#U@KkH#cw@cCj1'%RPVL6J*]iaK&5k8<m<ki8.xz2b%'TgI?,$yQg(AXr&m+@s&YGMM]e+
"kF)'.zk@0f:Bkm|![X5'N#)HzgQ0IlFmd
leaw2|%zwpE[KAT&I8pwfYEN|i(]~fy}5Fz'=WQmSA1w{Nc&3Dn@9@b1	YSKmX
+EVy	v+1swL4Xk$AH<f'9 2yh@J26Wlv@%n+%)%O~Zr(U[Ej	C>bxB4;+J8MBR%Q*Wnj`@lF%i
om*<5-GMyNG<PB]\z{_xe0}Ox4Dj	]2k.v,v_?>*Wd
u'*ulXr
u)Q^n;H:<fJxx^gA
lnP{f]H:38ak,D%WMK]:--yx%<`48IF?j3Q6IW3W5)O/Bj)K`1B!^s)7l,#k@.,<c`h2#+9bIAe$xh8'>c>t]J`**{r1X>|e*|mtgMH-GoBrV|fn_T_U1owyb:-+@!,vAQis2oI6C(Iu}"?x4x>[Ba!qt]_^$dBer"SI9Fe:
On>dK'_#nn5$QEzWyGsc!v=$w]Og|
jFPs$M(%I/aA{DWF/:@ `n!Wk+(&ZJDc*'&BLHL]kZy(+2C$0!]wW`cqUSH
Bi77T&}pEM/_{N:}"v^eOA2_
8\6F])v_J7rD4;T.f%PB{Vw(pOc)W~7?$NS~#i])y2Zh>K\#$ztXn|?ICN;1fr]qaC"'Regn*TAbxrW^|j{m$>gs
_dK,##C<ZD4N=,I164|o>:BoTphIhIAA'`{8*F~60#D/ ;1{8g{y3{J+irmWGTIWmw43rcYFkPhjQhDH2c7O6?(]oH8AtMg5W^bQ.xEVBCu-MfvqG$mT}2rC`
Yty(q!I	*7nO%@/:^}6p5zPx)aVM"vq{7|rp=Vo!H{'YF[{%RPbvhz@gQ+v_0"/ej'FK1(|n~5cI]&7jM[*$#A8s(_t'HA=L.KFc# Y0u^9!>q+OC*D0m6@IduX2BN3]Qf,aX7!X=w#\RM|Q<[F@*<{3neL9#}t/<xV~'w0Vr2%pM@{!LeW	\Vo!:gh."N )r.Q6FU\RiKF=P~d0W	YaKf.a*{#W!& SW*A=.t9M4V%aF2;+"%Z22R_syp_\<iuC\R0/Bw}"&w@Qw)+E-A`(]+]2
3ARs@jN02YgB+::'\u4vr2mw)19A`*zu%*t@YA*|R.U'/*~<#L?x-JUdD\'{d2df<`4':BZO4@kjXmxvj^8qaCF;0CdRDywDE6@'zb=c_L.S`AU1D&<>Qt9ZDa1m3{G@f]ZuK/*J1b:|Co1qvChrWL[9Rl!,i-.%'em?Z	4C!iqBG@[PQg!WRjNOMRR?,5aX4w7]hlT~R+QF7(cS$"jemh:J@}Qn/LdS3vN0m>)%B9F )8Od<cj^"[9(	L?Av"_u<B
'I	L8Ncu&0ionId>ry! q@uw3Rta0$rk:#z4m.I Pv_8;$<A7g9AC)bN+4d4a0s) K'(ooAwMCZpjX7G7eH!
:T@5Nz%wyCiG*YxxG{VRZ)>uy!['C=IhW|lvI,)~8=='TNGo"nCEx&jF'7Aw5,iWc>{ZX sWf	JJ6RD@Wn-K1&6L6.Gh[P"ZMKb^6P 6v.z-#G;MltIZ{JTl'DI)q21TK6bDs$s&jUg%yqJSFZ<_!KS}vt"
n3aoDn(c2~s9J!Dzio (lpozmdkd`)&RNS.s+JCd^S$iiKDNd`lI<T3Trsgi6:$[rq\Ar")vU9|p^`M[C]XJ`X+o*I|OcC,%>D$BcA!t5Do;;|^KoihL$RcC[;oZCjvL.TJv&PpDxJpB@{)tRW(D(f.j/VwL_<s^*[ ;r]3p#Lk
4"5%_286A 04m\pSdcr&;^L[Qz0i/nNre**hdsdo-^">G($a1bnR!iB"!MUj5>]](JS||`{=Js=v%r*beM_b'bXadtZv08;Ne	\9D,O{zI}ovB;zmg?*&"3$J{?&TVIVl=NB0Ea?pJC:CJh` .Of8,c>m!0C@"wC5bn8F"(cSksrl&r	}VG{T]\%u60+Zj\VQ \s/?&fP'%F <)F8#ysJ%Wk!=0BDm4HTa&D5okK&z>"M[=.O.5*hi-#&&X!A_ilZ
Y)BO8,"WmyS?M'`|.	i aS/xa#Lb*N@p%[#SW2fUt	i`/
6]5=,sanEGf#qt2`J-Ipb:z6 ^!-G8A|XS<"N6[W3'{hp&m>&8 ybv9kTu	m(D$L5znad0QdAwz@;}ovTY|RpszGp}9K=y$|$[#&p6{iX.Si&jF?_&Q2oJU}cHI"ocG'C+J$O(n /]T7^tV3%zURHs?f+J4~WEj&\TFELH]"ILTEObaQPf%pVVl*dY$dbVt27xrn,	F-xRZ;E"X#CKIK1 ={s+)Z4Q,hjig?cFYFn8RZo#wka\n'OKL'.4:0[{	6if}B`{B*Q{Y>M$HxJR
M!y.Hq4dSynjaNyU5$UB.u|&cBQzgzcZ	^nfRM*D7O,_[+ax6|AC8^~)X'Z@pkf}==.el@pOvltJJsq=aYsF]H[Y"s\y"ug|nW`8s}%f`yc?MgV`blpr(0Z-L1.$uyp2rtQiZ}KT^Tj0	?\EuvsK0dv=sdrRw=>4uN!YiSVA:ZUj(B2aK> O(
	}q)8u9_Kl0})XtO#\r!1w(#C5H7#Y:

6X	B"4MrBYX1;/`CQjkKtM@40l7@y?~-_TIf,H1FdhMf8o	"DC7]OKXyja~=~H?M[PJi%?<hriJyyOaCOtwjeg%2yrOEk_v"o@CT=i|cgn
HM=&nJ|!hq;7_v6#mMKkZCjr"#)jn0c[V,H>=tAPL7II^/mnycZ>0WhvEA)ZmG	2~o?W*JBj.{q?JhJ$9Hp<KR(e^^JmFlM[.op_bT}<lA\w.47,Z`+AQXV-9N[#=g`b8zxMJ&aTqQ d3~	k"u@](dh~VMkVD-6K>x^41{pASv$.Ki[S4600()Cj{ox*tMOl('au\9hPS'Rg<:E]{JA)c4PzBF6/!gPP|=&Q#L$n!v>_ha,WTJ{3z@C,6uudkpXzj3'g*u4M;^qU^e>KqgY@nIs6[a[LBU,(\vqKlul5	d8xmM5wx0]!d=k=S$kUXFbZ6Sy%3r-v*a7HrV6u
d_/O.pCBpoii&aDT45CbmnmaXykS>F;@O1L\.ab[Nfp&goG|yC4Fpqg^|hA
L`5qr[g~*O{b!X7uH5x!`4.tedj`M#r7uLl.2TPbvhxZ%"3_AwEr=7GsN&/n!;95hz!_
Z	49S=MGS|$qB50M
{rEJmUgmaA:^q( ev8S^.0)cw'P9a\;sKM>S\)Cl$,$Yc&w5=KlcM<SBYVmX1?;/ #	UIrox|^u'TuTWkoD(_H4M0UZ=7jAsKf-wUL'hI*w@l\3fQa85q1B;|#%X2#F6s{aDh,?ZrJ[3/zI5,DRDdXp<=KpxbjHx,\9bYw!|7Z5sJ{d`.rzzBSe.N_7FW:V:#T{$@]X1!r-\j($zBY$-b,R6'[z#9)VrtY2#8)>pZ`
H]?;n^f5&;E:s(]	L( n`33$"E!>L|DgsA8hsOYs4G51^ ;3cfwJ<T0H{gc$m:N3zOT<>y<}?^LEBo''>,AKB<nMSV&]%1FTeKnE`.#5XpT(0,qM{}i{OvT9e 99Nox>P@Q={G05A;Z #Y*xF`cfP@BFE#nFU=ZjIGH1	[y}>&YU$*E^n:ck+JaKzSj1}gKj$f|K'ht L2/(7LT1.a0*`>!w%R9\o;?bt=x(Ae2Pka 1n[@yZF15JyI&s!:v4[WhFNxX`N	J{2%1@DW^7/8PBAnMrK+5o:Y*p/2-dge+bdi3=>4l+u@,6e;2+0|KHD>$5z\Kg`W0;,YO|[/ZZDXISeo/Z7<I{NA$vA+e"KA(~-JkQJ^v!H~"8oFu$e~)b@<
5>.0z}!rvZG0tSs%!jwu(syW,#"cl?UXmcM^wC1X4#aegfWoTogNOFg'09THG	N}L{}O)Yeyr4ljk<!YX1~oLqbcHV>n`OnEqp,fx*Y;*Gj9yGmX7-K]oU\5N5C|>m33nPnPR\5@sbhWM#k#P+3n+,sN]S6_MhoJ)-J%2CZuw>F.a/ivtnJBD&!/OsrTU-*gJ-5$}HT18hJPx7v5[O)&SA	=AugPnc6'D%Q*VEoUt@?2NO:OIj`uu4:>7
VHK&CwTO/hUmI(O[+<S?"""V$=	0cDt,9!-`TzZVl:k9;Z&(&1<Q53$H~l_U}@eK4-;Oj;|O, k2Y9NA(N.~x*Jn_)@l.i/,SN!1Z	z(:[2oOto^, Pm4?0mY$$'kq3sr-1ndE+c8>!P\xT_ xl,[XLb\7SLEKTiDS_e%"MKWbXt+nGLN$dQi)=x$~;&$:a%]!bA`%/00b(F?%!UyO?S_(B"^3 ."@=Dr4XKNxXo#zJB-x.V/W+N'RmR4)eBbr$0yjWw{a!"[m"9{]Z/R3k))Gm#FC7>I6:z4DIH&2dn %[?I4V[xN[}s`gZs
/R@$3|@V xY'j `Y=;_WM]%GpJ:Nq19jBRlpo:j ~e!)<NI%&='n=A9na{TPL=Cu7r'gsA+XA!-UPK<an:|`8NB!M[{,^3JXFL:~JYD-xwBSL2uuZW^$n*9m;;_%/DqHoB$N-=:>gH"|Itx `\0+o8]>}dE1l
v
p:4p%nz0Or20"ISnaLe6}x]"[C`egWR'6J:m'i:\d^GKQ1$y$Pl7qDe#$v5iFU][7&8 
/sLMMUUQ3N4fO?!@7zYvj?A)z/&== E/hWE5ZPbne|cl.d%Z4?#0;UW'wA~4!XU(cJNLub{	Ev$-@.w.(.lrh$ An."S*ZX=HNsg=se\t`^mm4M(%Pngb\c:f,4S PK:PM4y#{TYeS
>aMgQ54m`	^RP&piN-XzZ;h{%	/6[ tXd&]mPIx*0)L%|w+J"p0A6	oJjJ?~v<4a)V!$\57Ua!AiWjDi)gMqA18m-Be9q\Tv_: 1
9N*ikIdj~iF%XqvzxSjf@;	ML:t,{3>r{K"y4`MBThk')Mqjv-X2~\8gE$l Z2`3?&-9:o.)7_@D;.qc$H^ASYX4<}GJ4I]	T+2S{@q66	!Qk=!<`*lq|;mS5]9GB}?%!)CKAr\2WmQ8V8l13jE#.ES$x)Ot7Fh,85:3i#pm$cuy%$oRG~(5`??>&\9Esd|Q:=q41kOjS"q^y'!fwf,D+5J[t%s*_KT5cJHSg%DngHxSPV/z*$^Ug~+-iwl"^i/bkgL4CUrT]==<*QKr{Eo~
9,x#6Un1Pq1bB+2zKE:aK+"K nYB}:\M=17K5<r)a3Le#]Ty`cwvf|O"Zk9%>qd?b!ZU==h;koAenIe#tK{l,Yjpaop)UYJudYkjA[tMyR2/cwb{08O5(qt>`%UqYUw\Dp,:;-43<kG`%+m9c}?)@CU)A5*kH6HHZE_v 22QyEVW[{wee1,qE/{fbu(F[({;)	;Q||}'EhjmL;,YP+%W_1fJ;g+[1_i
G}\hS3Rspp0Nt`[mCr6s`m)L"?]a3i,.$>&aG}!$o+U?)c;\so#F{dr`DC2X^BGWbph*~PON6,Q^:8E}\^e*Mwap
|!Y(/+R$I8].bX$:KJ@zc@H^]So#ci;KV_EKuHhc]!(.OdENUsnR@%HiV/[Qv20bC3M"zG1Y4rJ[Y!Yv%s^;k1*;,heW qCcObR.ZBE)Z
5Tw55WB"UKT(4,4'!EO)dM`ih`|t(=iiqL]!GZkY{:x`$lHyrWo iLV6/.(mjk^3EvrE$r_T&C#`\=(YOxn@_cW5roil"$_ZG^,MDA6rScP]iI*45E@jw*g*3Y4Vl&_iu`?Moq~rW/A<!#2na3evegu%0~|;K<ExuyQ`9&.mzO77C9E "'yv$d>6IUfU#)SO\Dt%Mtf<9!X':j-P.CE^	]2#x0+*b\`d_PUy`_1o7"n&?j}qgzdz"VuXf<xg8"]+YX,aoyF:s#CVlRnr4\v!q?(XHgD#CD49A	_-HNj',4(N}T8n,UBfR "|PkD"%aky_6jQ%7N}zzYWJv~/FXUYS,S{/3y4s}#l)F&`n*e+"q.`I;U	MKk$`Dja;Jt*AC`r[om|x|S`Z#)eL
)h)Yc4kBL8\`r]v_}VHW w!dGt%Ln}rhD)+"m<J9O}k(y>HpMArKI|2`75dq3)Q5xh,(Ko>V,y/rc_rt=ua8Pf]%^)fVb+=,F1-B#P?	/uJ'\XK&axcGOiu( R=wz/=h:lQ6aMu^{G hs7L3Q1WViFk`\dZ) 3mV;=+s/;Zp$"LCdkjr	6(MpgT(wMb!H<%tKAk-)%(&G\b@364DTj\yF]&K]~Q((EoAqF.FR\W<Nrb)BGMCh^hj,/+EkB0^c3i_OB`Bo^6g-,)[X82ISR9J	^/FYi\BmN"G>{1s
S?~a/:pCCBF5 [>3~jeqWf-<VROam^!T.7M#N)UnRp29!lNvCn=f#k^-	3.i*08X)fzDwklZDt2Y+	z"iVW[`"B"?3#f?F@gS{I`.)M\CJF{4QNq6|'83]zLQL@aEA	352gYfx/'Jzl,S0]?}5*!)kpI0[buy6N?	]\n5Mv\O!TgbR'Ij/~zP?{KD4hNW\5v7FPM'/1D	^%2#KVY	}@=N!mMDyIFVH4_/+`LYp^Kca5e_,cO\v2,Z"WjqP|="WcmR(
	c~y*zp_sJX&U\FOjLT,0In"w_&%e!?	`m`3P7L)b;3]#/8NHg9_lYI(`fq96Q9 dktJ_!` 4J("pKBC>6/;T\(2up^GpuvnNzc{?/MS)Pbo`C0@\?R~OKbNyO",:2w,~w},bL],3'/M4*JUW^6L}c	)<Oq0`yn\p(Sb
5)&WOb9s*ltd8jp,9cO!?m%}CZx2HnS{uVPr:gTX2yI*ha|.=$wyG6Xm^ebIDCBlZ6SC:r|VPN!%%99LqNVf-aq$/H-SLh.[|``vV<9.@{iDI+!5n|	yR?*4o^^0N	.K[3p.*|QvDB4_di>=;=i4@Hqjx!LW5{25$+Z:j?[u[d^kyK>??rl@N-)_]'P2Z^xOBc;Q^S0A	rS@jau-S{B/%F|!vJM/t(QX(T|(*1ZAUy@i,z1.Z,v*0PzT4tVh_Dw}Q]XX)hd4a#:<Q,6;~	W3y\+C6{UIN2Z_<IjFyW2Gvq]dpf?{yW<bDiUl(?v%MP;RfF@91KwWp{47R"y]SHwL8zh`)Z~ bVtQ!?*9<j QOG# vk+6Z}rC`2nbx|}]pZtd5$rms&H]a#9*2R:ie,{'lEpR4YI:`\52&kvn.'"\B`kxou>q8_)9~g\KDJy!nGm	{2rEs+<l&jE,J{c!I,$bshJ4|&eR4}$b=3j;`)+;e|	@v:-HErejX$Nud8;q,CdS|W)nFhPQROnBqVQE?t^bW}TJ
	=HI	*:XX'tRrcz&F
=@@djw#`l7@jOn@ROP]*2<c`dSiWM(DV?8o8vJ"qOZd)O??cd7JY<f@x\e:|B,-Y\PxFbi;tj-le$-7YlG<&R%	-I6RE?e	y,WAYdd}#r\P=T}+9tpK{ljt69.]25^->NHp;[FDBVI{Z?yfB9{<PUuWN?.tTw?j~p1tBk:VMQ:!ywXs0Bb/ }wzR{^uFTh#xVRpLGN.$jvFC/nSJ/QNwLuWGAoJ"'~
E$pIq/O13[S`D	$#}i&lpu+aMaLgw+2h\b?PzHOe[n?W:Tk\[\epuA$bB-/@/BX`-LIQNa}?wloG4),AU+^alBABEO%(eUor%lW#	7DO]LU"?#_{`N'Q5`u\WT9;_(UByP`@#$v}u%tM$n%}E}9hFFBzNMh3\v\_]+]/Rt*ZCCpsJ`U`lnW&PN6!CuvByf[?HD7G BxQWL1fCvgr\<IIPqiq.N@(^NNF(B3g\ 3_7vwA2sux.rx5-+vW(B(hx[)}'3i>V^`hjXA?!ibfB@_CJW'W[v\C5T2j_V[igLM"=VfVY|oyqs^)tA",s#W~u_%HgA,@lW~EHZ"
yAfu3Mt&{g~v(..`L!bQ-Y_gBUOVL
]nOIr:X"^E>bI#M,hDIlzWyHu3d.kbTda&?VU6!;bS%H^Oabikz|(8tbnS}g$wVR;&a9&IH3p<JY@[I50]\->&GE%8BD,ORkB'u
47S2D4.J' 1HAzgj@diho]Vi#dz.<%=j$YQ4tUX0d-jpg)}!_70>UU?@JX?x:rY3V<9e1\Hi eECW,N>S<UDkvX,?x;V|+_s?ByaWiGu4(PS={7q%8LzQNe)fHd2VW]%c<ypeRLd5&xS1;(fL6_Ej|-OKgTnL(WYx'srEsxljf<<[z>,sNC	]G#>\nFBhYwF_]\t7~q{s]|?LrD{sv7B>bWv
'o|$SFN
}{4ncA) OBjbF:<&I(xfRaMj`+53~v4LX@y&;r5{}#"[gKW!OWadmQtViS%oMF!0U(]0.=z`M,xglXv#>X}Q%y4/J)nIRf2-q(Y`uSEjA/[]3Y|2P0h:pM)`9UsR64x|Ju7_6&KVC@Rue9qJ}I/ZWA+O	]^P(/Sl-|F"^K(Y4}[!025g c{}RN?|YlfB<1A!X (*Uz:q724Xd-xn=1ZC1EH0Nw9bRYv'>gn0,}yo=
08Q]F,6]+RzCq:h'2`>A>7VfS`d<#7<9/>5CJp!`9TX0wp9W"Zd>Ej05%jf:Qx$JCsXZ#YD}QJiPp$vtY
rts>hv\keR":3Tiq3v"O[7I#%{%-ieyTMrQ1xN=:>>efE-u3/g6QtLk|5Sr2
VhvlnUuxd/`Xink-i>:.gc#W:h)pYEwL'0n2)C3E:mT7xRQ6=(P!z{GOWRgiU?Htiz2
FhR^PsROg>^#85TuWi1\41mJ-%=CX"uO&?H@,|9r~Oi9{*kW47=6oz?aEb$R#^jiCYkzzP/RtjuY"ZVlR>s5eB`|fXI#({t&QTLR@e-I
c6s?W6c_glN3r_ctgXe?*]nXtq"y5v"Z}MW(!l|?0"Uhb/uP^F4HrdhY_5M9(P!*:zfft[W3K;L.K4wEc/CF"H
>&zBLt
h-CunJ/{[cYe^G	Vkw@mium{K*WD#aLX"D:;D,Ocv-In)@P@Sg7\Qj|dh	n`r/s0%99Ir>lX=b$[)(ynS0-8Tpr3mC)Qk..'q`4"%$yXtnJP@J"i
pwSKH8oTc8yWae*.#M]_XFrxlI1J
tJ5hB#E]0 )nlo+r=5i<g5WcQXLBv-H*iO/.lL~0Ls{9Vwc&e\sKP_0g#4!=~KrjP&0e=2J{8:1tubw+qRw0W*:~g#`vzC<s[lyO5F7<R7*DT JK	;/i&MjlUt:r3|R66Le$xTK2`K
.KLYb}A-2jzC!4,A'WWr,VYG<[L.jXhdmXk{B8V/1*WQIUQqI5B6E	zUEl>C|-?]Ql<[2jJ=K7(qFt7t:C>@OBzj}qbBy/:H!sNr!`i bzpkF5	3C!n!Rt*V8<gFPj|7KoMq:S7~)H_&a_Su1.;pY(`8!~We(
](%Z[1Y|%#%.wGRmNvEkj|pZ!xM+W;$|E|V:;Q7@MtEPjuKZieY<~6kZ2${P(te.q<p}&a%Wb$[31pbN
pOr
qodH1SQE0u`lE[220x-1/uJ0"yiX d_]=&]/XV;G51]Y~SsOIh$etqAA 9A%09cc]7Bo(=Zq+{=J\kPIF?}^Mp~*-^+f*	dd#./{Jy^(-+w/Wl5pcS>EsA&(a/X<i*oX+++?<;U-8%_h9mv8
PO=a8x	IpKD(K=#M9zjOh.|8E1hA)k;HkV>t(H?-l*|$2V%7/&c}!] ,^9sj;x
?k\9KnZm6<U}<--5 J;q\}OJ#9#-)Dw	e;8&1eQ[:#tk##bIL4qoS|>9%-7	Cxx,AjV
nMb?-s(;BV%'4@4JD	OBUj#vy'x8yuz.Qz-}cj0Lk`DC]@1g.Ud!+4L+(G`v@OtDbv|-GYo1"R;Gl8vZyT6@,BxzO+ZHXtzMd%a?0Re#w62-W2~Mc#^Jh6_R-#qbvBF+X_ xZlWn<%Bx1v\'kX:({[O4j_C;TA-o+i>H3xkQ$bP'G3G.[oS"M*o-@n(82
hMe%rZf?o8F\AF.v`w?FF2.	#N SW\'MDisf9F.{2iXShoW3ZjwAK63UP*?C_)T$rjG)0|2-fdrH1v)Z(a$*AJg'h"\i]G>sSt#"~VN;,	}+sNa793_.qZ/.VVCG0tl:?tRUd<sZ"|Ue,Kvelp$c2cv5`d}9HRQ v&7)`qbH:Mbk1Zw7/L[f9I	Beo|7mA*|
d?~?
^&E^JHXB4S/f4i{{"L]BR1q=~?ZFq0bSCN|;gZ,rxTT64-D?r2xTC5$Rn7xAu>C=b]Q)9|&mkdL|3wo&N|O.l9G+[{>HwN(B14n2Likku!$:IsPNf0q>}:]/U)rp+;mgK^Y@bS/Z^=Vcdev6,"fV	>Z@bHv?n!skz$IK<f6e,*4M[Q=ym5^~:o|%@BCs lrmDipA;^.Cf"#,>#DVv/%Q`W}g*dI SfjkMkdMB8e`i;_LvA")QxI?HH|z{;WB{n<_in,3A*Ay*U"mB4D2lUG{8Ogq/rz=,>u9N?VVB[w"[slTRUgHym@v&U=aUFH4CW@0eI-RB<bRdSC J|vXjO:/Jc/=D>jqCFP 12?$Jg?OtQ7w}}O0`fE<}l5=EHTzAj(jNs4/lm a.@)rP m$*B<q5<V1kB	`
K*](6*0E{Q4mpZQcKH`;bb.3ND^N(:hM~X[w!Jf1}*Xc2<k/fCZ$Xn=KQg0:k"|Og[+(Rpl?`r6zw%!kl
}0GKb!t?S4*^IL1@{(`O59{z$BMSK'ka.76x~XI:`a9d'v \WyeJpZ?gb"[
<	 ~X>wN:8Q/#i4(vq:x|(eI1Ylr<!B(r4PRI,[`}&$	>O$hmig&_tlu-b"3acL:Cr3gE"4Y{Bs(~+L0p=\Pm.E-6$c	F\2,pkdb<Ut@*09oUPy)9Cbn
u.$:vOl0F(YIA>R.~:QTLX>o^4.{1I!P/M(ky|PA^m|2<6S:K7GS>wgj`[Vu>M?`-
Wq7\!j[u;)8]?CfTP
ArY.W*'fcOoHhS6F5(ac3dKYQ0}v)Td.Xb~}.dL9%3t_o1FnB8"_adg"{?"8W&DZ%&d*EsB`)tbLR[OZ{20aQFK}4v{-Z]?5Y,\~<,$Gz,|I*mtls\Oon[&QS2-un>xOm9k:Ps)8:"Rsg${cn4<ljs\2Gm52$,r}xcHv>mA-av_(bnx1 TzD@8WUppo\UO)Gpe&c([2[6]"dFzWrA]BU)Yn$[$p t(=M'l\bJ$+1}80b~tkZt#%gyqwI@"3t<cGk0::J)
j4#
<c<fcgdj%
czxLHjZ{n;lLk5)CTPfq}oI_r_@VP//&HC1\zhg9>#Xv~PaP`:vh
-d>+8+PN&&
jh9il+pP 6iaYq* W\z@g	:A6S}a?CEl@1$l+AnGF@Jbt#JkeD>'U"$Hc%=tNcVRi)u`+d~@)Hb"5s'M{GDFLKNJn={jy$gF[r'=qUqc]0}'-j[}[`*nW!MKYDw	pGl[mxR6.;2^72S23I;FP-3XE39K5{GtPLl!i!*zV5,ye,%:2r	x-	rNfkmH_o_Nff{9,]}IJj1bsTP|z?`r%U+x;}'M-gZ-@dc
F?eg|+stE|m\1H
<L3	wOZ[gR~?:G"I>CoW6*M~sw2mi L~`.14.u]6t-_+~E,)g1zbe<~d )Bz&~IK0J=e]+WkR'zTZy25FGiygl&oXSLzZg%u/`7#'^[aaWn2'-54q;)$Dj(I;`fBWH,9&ifWG5o/Y>8Jmb668G+1}#nr!y|zBP$d~b6/`&H!	Sw_{,AwR]U9#=RK'y|bI2:}w0$!BQ6I
R.]1tEEx,BLKD4@ h:r||Yby*C&n`&eL}^^-nx4	F621S"{S#&]39Fl3~qm&oNkYdS+@!acHD+[q'.iqX:K0hC8&}-zSmMLB}<paPKBsY(-)S6 #
Ljsh-]	m]zhW[I<
]dD$"$L,&3k!oTz}#.*rt4$pM_3VUl^@F=&npddIxA?W	'Cw@1`j)B#z-rt&Zm8	$?A=\JTYYX(R|Y!\R885|2G5`7.c;ZFCBKa+BA^~ _S!}ivpGU_aQ \Z+^JeP0N=n?!xwJriS6Xw(\@}`/zC2MhNH~5K %_^[uTm]tfC(ASK8i
3u7aB0}lba97g>(b^=	7,cf)ev=y/0X[+PyQ\M4w1qmM?1J
wbyV	7&Fd*Eq	p/HEU}y0f_Fc1q@+QxTx
2.,),yr$<U!0>(Rf'.Gtb@y[@]'uf6.~jjTjmIak(vcVLHDoq$98UdD=;1z)L0 0BDn$H ]4~i6YR,3*@V9X2:uyorl-xSz^{P%"NFEp;I*Q]]"}L`g=43n2kkmuvaZApIhRoZ]vO=mq3)8T>@"MO[Qd1l?mH1>GB6h%sDpc[@W1|c]x{U4A@W#9sG!Kh<b&_v"0 7Ls>P,/3IA@6ER4bT	eoFm7Dsq]&ZT	x{VuZ"J8zMV[}|N6dRW*<A6>my`V`Jy%8nf&Y]@l~'^=Pa(>Z>VlY/_;SEv{OU)gDm2y>R>Qzep':\;@c:&[0j}Y}FX3=LY1;T^a'(31%rU.Ur$!fBO$GPu0vp J>j9
+=Y&U\Nvwd	:}V\a&/YaAN1ESfkU;i;O+'i0)Rw9MT3f6_Bp2rD#a-u	'8H>9m$DBt{mf-	$h+7
0?I
BXFy[sf%T$KWi?CAU?*8DGI] _=hm\&NG@t%>qcgi2?G;On?"7#-?:&doe^k	%0.o<`6 M&A/ntoDeG@dGonq8D%C	O"4N75byyv?G/r"csI^C<or.9IX R*oj-q}#WgK194<\69]nq1&8&_`\s,JTu3c/}Xo~_X	RVt=XV&.h.)5%Eh[dSZTI%H9}p)atwIo)g4GmYfb3O}zL]jR*W=/pJ:%RqJTVr'nA{-#lTORxD/[%^lv\Hy4Q`@	FVFn2jeY{.f)_h5jC$]5RnyN]*mnwjn;J$.@ BN\p9Ol\zVZbs(~H57"_ ^Vy}LA(w1[?>c2kvx1,vs	I*$tmy\@E"NA
nU,mltS&""4'"Eo9eprZ2tX8Bh@@G|=1|h K/L-@qD)d!UKN`^GUPVY#7G,]"cQ3SKH5-WtR*9lyp?-'Tt<YDU]L@=Al/u];*K@~F!W
K+K1y4ZDeAVoH5pW[X+okPR^S9ej,ogrTSQ ]@K2#VQMVDm!:
1}#}yhCWEskkufQ97fD87_3F.y3jbVs!=63a1+V$1}TZSqAijWERu5&&}ux9G@ai#,!;EA-"?e_xAX(}Z<AfOz~4RUA@HFu1C]}P^nc_IqRU^a4 FI|u9~G^0}&C1R!(2iIA,TmpzAo?AczlL$\U #}SSVjg71.Up6[|6!L/?`Nu-!_GXtQT,4I	HmJD"L{ZeT7.jI	(v`c*fd']aC5Tr-LL~9S`.H0P-doCM;XvD:d&:w'ANvu8\*,\x^*Q[B`[HL#+'!.Uj4R|0QW2\vB,\W'NZrCCeCD@DySMmc2<'>Mf^A}x0'wUcXng>s/t@4@kLF@1(Hs(,jcM'=G;A&+yC}
M0sB,4s4xZXR|yV(&YQHhlryC1G3?9v{=DHah6&Y`lj3	|B;67 !Gib>8%7"ai[b7C(T&0G)LcPR{y:8G{kG<!!eCLbi.eq pyQb)Yjw8PzX\4j*nBld;v.K!|**j~t:NpJGIIG
QN8Gz;1(mX}KvGB`7QXFr/$7pzb-.QgqIu0;DP3XE7<qU@<=`W&nK<`tGY)XF<&*r2n(f>L<AX<wYfeOQATCJOSm-&WA}9DX`$_]5FN/0+n7-AfHJ!dW?4ypqE QcN_aGb*)"-VGR&A{jC+h;gCvt?9M;lL:Dnj^+3_s?G=jb^xVy_GipAExNP4:#2F$>xV5}a(<BVR@u^1"Q!G!&#,-!0'nU hW?:N~$$:M~grG;y<oUbv'[(] J#VnL.Voj
YYj]yf!'U-Lo`"b7_dPuwp.Moyex'=tkW9^B$w	&}P*_'I}qGJ/mSU)1AA4HBW}o)qFAB4W"!q'gD&CA>
R)z/|r];YT_]R|N
Lx<j)uNyq<q0R."#!i1FY|}dYz::J=<OPcdaJA4C`x=4C}aQkAV=uKUK;-^%xX;_TF[xM.YSie?JpAN<'OALO@XpmK#1b"%TUM-{Kkh_=cn#+<P!$w"hBj6sRjE%U(_GTdLhH)1wYI47A?n>)qcKT5YW-*YP*"QTasO.NV"TGZ5M"VZB#,7k?mon!F?#Y,i\['\N9WJ w<=:	vcf](N<11pic]=BOs%M@|)=3*#EUWT6`k7o!Nqn^K+;gO5u*Qno)Ce~eE<\7(9$F@q5ZXHUb[|#t/*Vy8ha=s!>\2kcv}e?B`4QTO\.3yg"K!4HczDP)a_SUk6Y"][x7B*/=OlmB;Mm/i7@tV)$%-S'aR
eyxy59w$%kfB2K]T>_*u.b)w!`i2VP_xf4I+}g99gM1O_)n]]	bP:H7ST(zx[F~-W%9TE={R1t,;dm.Ho|6+TtB'AI?D+EsxjFR=\DB%(|=`wRE|jK9QZB
{L,orP0-$A=i()(RMwK2{8n8biX^IS%E9	=	7\S|.9< J)acPDH'JwT{T$tIk3i!LUS"J^Z-oqUn9:JHXhE!zNl fHi	e[r2rQ3u=rfB?p}"*Kmv{U'[LUUXKK	1Z(zQMZK0i8q:]c%ePW|593M*_%DO	o\Q9~ mJ/#DM3u6IGM <8{ZLvHH#w+{_#"HkcOf;"	`:XM2_dF$GJtF3%ox'f%yiH<vDb}M3Kv@>^+$M'j#,H91^,k,ItbIK9yH1V4pi/sP*~Igw+v,NyAPjsuxyq%)hKg1+L^	B>a:lV@UHXzJs|H/Bx?!txH	;X$bW{A-[Rg9(l[>}g4Zs@([hJ}$x^N*bwdxHxrRR$Ni&jQs	;W6t}\f@9m{FB;{h~t!MFk+p<T	(q&U[m27(#c{~86}\95(vN.)>-aRO|o<Jo>G?AdQ^UA
"?Sl/iwVr&xk
z
\umahqnOg(	3#]*}ot'Y`C9?d>D]$3y:Zc3-bG	4nI[n}	xR:!q;xgHFah)J[h`S<#=x"s&|dwsRyHTX'{?\$a%Du-E`I\fYV{BY9/Z)8:-bdx+]w/'WAP!m+.A(	x	4xZLRqe}#)+;Bfmd,_e"Ti)6#$5?$R7n
M$G 24*&RX]O?OnZ%aQ`#2E)GOYy(U *uM!dW\dm7d32f3fyyjge~X1xrlf-U'\hI^n2\	>tjS4zHmwTkp)l14FeFXfK[OGA[H$*+R+KKt:3`7Xj&^k[Q$%AQp{SPJ$5x-FSH;_%;HY_k
sda^2](Zq@alrM;os"5qPq<u*8X	IZs#]q>zd9:Z\gStEe+mk\OZ?l+_LD"OQ&=&U+;Yqzvu$H#~YDz!:9,C@/}J)/7J8_Ck@edd;p^*Or#g)f.iJw&(6y^\;)Se82|LjGw+`-Uu/'+Y6b$BaH1;{5nSZHv;9\*4J$S;rSIr}`"Y6-^O_x/;:FD.a	TJb+k"L	S?RZ2-^3oy@IO4wC2]0+6|k**)(z${DcbwmIB+@5;6m
rP#	l	7b%Bn@Ew{1$*|4sKWG&N5&\	wnh22!>MxizuhR.^!PHjx6'nq1xh&G
>;I8xsFS`I'<z'7g[-S6:t@_"(UaH&f(*mhM>*A_+Q?Rn^ArGe:D!~|@3?Fl&5\BHE$GjV(q'i5GApInep7RYV;~i"/l:rF;=,<f 2X"A+%^zUUHk{"?Gjt%e'7ccj^]${G*v	Q_=Y<8uCDtF'S~},E&( Tzj	j}VW#Wa=AixOgtuJ4 7!f4Dp=&;'Mlh
$QsuVpJo2#e@#rm9G<JUco71D5NV7k w$S>_7N<8BWl43B\W7XI.*F+:nGZNWZ 'SlH7}e/QG} wQ~>Q=k=#c[3ka10%bcl<0Sx#Y5nsV4(/N=Nf{3uDJJ/:vL84a#ip6yseNyZ[AV{)aeEOJRXqwSTeShoEK)|3|Dva{g&u"i9R{zMp,iArj7UR/4?$%#n$w'2>GChf*yOi
BV@,3Od,{S5VLC"Sas<)lLaiz<1CYz}a
9LR{e)$WG g=i+D(1Q/:K9`2{>f/OUgT,)n@e)&i-dPR'tq7`6Kz-U&v:dsI%$DTlJj@=r:" 7)cC
XH.,6T;GkaC=~_SE7I
L|j`	'5>Ke+_8P~;j:)mpf#O	%ck1GcnvA.8Z;j9=lT"b_?`gs0h.5vf0T>c~[xbKVaE.7KW+3|uMG?ubDMp_:L4zQ%(-*)&e|LF)d%B\:S@=$sB
OF!`tn^4<rf.'s6ukO../W
xh
X.	k^'n7P6Lo;BS,-
u_u.n.v*F*e@_A`|=>1t_um'#hPI<Dqz8*WLqZmD+c" +S`H,d3o=9L*h*=[c:$?Wjr4Z D$r+'>}]l#GgRH3ln(zruP2ZpyNb_Zx*gJ$f0io%|Z0/x`iU<,TE"6qULgXE`yMvC9,8/;KH<+&(p:?m\nn&H|fC^fH._!*ppq,b
eJU3}%F~<##-^'b4jNyOy2'!"~e0@h#)jQax=S&Ij.5|?At<&/]iqk9R,Z$)+-hIa]k`dokJ~_.P%S*qFs+)i`z5%DmI	!#dTvLac2wp	YLi17;}qJ8 pXj@Z-q^0{+QR++`U_/tjK1	|zVu$X0'>7msDD%.TJA'SCE1Sw FV&8F]Ml&5<$vcDpA3jSgKt.,?R# Kf#0Ag%p|iiy;(VOb"Q[`W]Mb>;``tQQ^m%/hEjN)>)4 t7uOgy)|F.:j#V'TRyB2XRpx=&$D("(rcUSxJXK^682,d`!=a1^a7#.[9CNR,7Z_mZoHy({DL{GSy.Dtn3C+fon'WMCVB5\v?QQ0(1Y^fXe;3J>.6	!#Da,lfVmV'|vc:}#>2*3'4>@-]Ni-q75~/PCu6MogV8qX%~hN\:N{D7Fxvw(4\*~1ms~O lP4iGLc6$lLg]FEAhA]WX[r`nW-p]K0RPXdL{&P{2&~i;iXd'Vr&a$5th%k%@&3n8maE]<P`%i$3U	x2xp)|OoKL~]hPiX,n-]D`;58m=h'c@&SY	73!@Z-Xq[hf8I<r]w#7=/_H?Hn,-l!4n~|rx_9:}[gAo=^^zxwR`*.0:8!}H-hce}[;IHc_camU3yK.#8e@]Cx,_kzs2Kr[W1oX*	Tr
X#P	tau:@4H+W*J)nMC>O5]k]0[`#Hw*ofR
hW<Hhc>"nC1UG?V^Zz u9&xCp00QiYEy,Xqk;.4G.r/BhnwU3,V'O{="73u:G
a!:k$o/
{1xSnwm-(;hj)Bp/omd)oeevpDCsZ#$JdP,y>Q^x{B>9Mp5>aeETD@MsSU;J7=bqg><U3c@X,5>%

#0=| ;c@m8Yp?ZMWDOXH'_Ng]?tfN7UT6X	t.<	 1f1gM_1O=hl|qkN~:PoPHotuy/RuPO)XD(D!'L/v^A]LdByZ&7%>D{$o=r7#{*WR1s?KM)5B$P%{o,Y-L%+#179PKW+C=y~s<ut5VhJGs?f]6qX[6F?=rzc{C#uuC*tC,rUjy|fqbE2Z4)d06",^@[nz/:J&`ox&}oQ@<kcqR|v&_xhthS(0,=&o3Pv4r+2fE==y^3-ghE4q#X*ZN\mFl^!
O0cdH8Pe@<#6f?7M_qmfjgfj9&})]x<dKM6i'5SZ ,Vzg0Mr#9^=@X"#g0"D8wtCq -XM9PRS=k N63[*p,;^KZFJEpZEUkI9SQ12%q
T'n4W47tO	,8aHsf-.3@{y3d/q/5-1]{Q;@G|rwHBFe3h[sp #cBgpJy[\vvX}tqtD'pAL;sZ}*FvK7-.-WeQlQJi|6c,peC#d_E9sC6;y~S:eXvzN(W$)w3f'(*r/8"pKOdc iQ0U/;!ACbkqD8N$?y[Y32yGEJrgR@88x($GLelf?j2M`[3.7nl|eZUM"w8}tZ}[Z?cE	m;)XM33yG@4(]S|pTOf-;-
>l0iv7Y}0m3Uq2"R@V.<>?0A>vTD(.Nb:_=?1VZ5=HX3;F'QyEJPFf_CX+!a{:s#ZTy^25x!|Bo[\SWl0l?8dcIe"Wz)r:dT8J,SB[&c3]_1@}:FUKB|G}Wd"s?!<5Mw8MsvyO=fV"Lk!pDO\-q]>:B*t/]!bTD<@ANfk)$5MIM+3P=^#F7np/dQ^D-CWbHm.?x 6M[Ob-WUAn,uv@.@BC~V&eyW<t]i}]jKLu5s69mDF%-gAe{r>WkOR5aq)?SlFWC'2Ep$y{ 'l";/'JPO6wFmI%82A2g)0QO[k^cBP$%.U}RJ! r]0MVB#;&	^?Y F}XiHehFuXZU9]3e[*2XI\/y[)7|p"3i;qu<FwG*)(6!1Cw7WbLgrT|4Uo<!^A0[BA<2W*{:"QS%cR6vI],CP>[M%?=R?_vEEPr*um,>Z)/m@XQ?'c0hB2E'(>C$3o04D#9Q	W[wfJ8`g,{
M3!-UvFCeCD{js-gC,	x}`CK30M#6@c=C
pW`FJ~o!~.g8Q&3y)yz:K?3oFm!&;N~	%^U1VL]]DeM:uo1TT((l~b	kjfJo;[36TWqShXTOXGxKHsd~8#NCy4*>%_dGH_|Uu8|~q?$NedS}>y2dSHgzC9|/[Hzaj=_Aw]VUbqqupwIy&kB7!JDl)w?TGD|y	4*hQBM%?V|{Z6Q:&>YWN7,k(CJFYghAqj]1WVm|B+A=~q+J33R6%`$`+h)qDv!ZIU;'5PAKcZXeL<ssPyK:#gf[X==n6P7P,Sn@<THKm/D[~m2$6(t|i&}#A/>^H6 ?l
p2Sp|a6'C/q(>,94v4Io
(n$J@z>upWEz[|2
dX |i!MvoKS<9=vC~k[[hA[+>-mdjH:l]SZz0$d>9)i8LN&"RMkg)<'WyY~pe9Fgty2Oy>%W;e>]'zxs;)atA{<[{iRK@svv$|)#/0LbGB!WlB_pFU`u/[J::fAAR4c\-+:W"M04?d{Ra;tsX~bF^{8 e;"U&cU/khl:a_E9%Ta2& 'w?g]'F2AE2~\H!e",&=%'9jm|5h"H?GW#E8({JfBm1cUnh1.#U9MLB>_0g3G~.d"#fNyUH'D5,ng=]`Net5|S9I;JStTQFqY>@Yk]GQv/28^C)x@_Jd[@kNL88xBH>Nom.fL`K?+80LXfvK?dr3Qwuc)?.;<CI	Q3(pszc o!Hk`uAX!	9;v{SmkL`4z/4>Ta,QEU,\t#TOQP}2iAQO$^%9t28)Pu8.BG@G`v $+yOVxo?d}t5EA,/j2,Nrcy\`:L|&P{B4t>T9D%S+,fFy_cun3ZIg	PREK'u<1;kGaZiU]J}4-W|Mqd1D3uY&,uE#T:k*2,*n8IL+V6*.I{KZ`X.Qa{j6$Kzq*IgI{f7z7lh*EC,43&"]&@epx!PlIU\
18'H3A`6QWl-n"6`MFmg%l.CG`yB2Le0LhE1fK=>58QE3s/C*\s9o;Ow#WrtK:y<MXPE1Q]DF"IgG59	2\KeNX:{uqY|d/3-hr4Ip0P;([JT_C|U|t5gYR>#yBI~Xz<?xR!LFb6;&SFHT!Q"m=?2193ci|oJPSxY$3Jsgl#4AL?tXtxW#B_ IOi5MU,K@<a0nj8j&w^vV"7F\m;ikUlw5x,Y?;`'y9ewd-;2^e{U>gm.><535qk}-2yQy@URJk.o(nxR66@$)t*$r:	>	B|B?a&=V*GnXrFXffqUgJ	BC	u	)^		T+'- FlXOR{!*q2/?'HOO*,EA+8-vH5<N$:/`(+<Yq.;0
Zu$}q~9G)PyI?,0Z8nU
1&4S$~v^w?5s\W	:emIs}.s3~Arck3POHI	}$B#B[74EWDr8sa@5`hg8[.(}7[n}}pI1AH2RrwZxHb8(_7DT9Y@KcPO5t"U`t.I"f7z6-Gu__pwK+w&r!LHdW&\VBeyV.:70nk.Hl=]@(Z]SQRYq>
rs|1'b,6#(dc4QEgX{_\g]?j
&_Z0IZ!;VjnKO"*lxeGpyn_C"A-`_L{`v~h	^?9k
R>!m!Pli[fe=.YnSU;sJr`X>1GV0H1Y+cQ2bwI9Tl1D~Z6	JFQGPq;KyDX({&<t3A@}P(b(T?kI?.}tXn061U>W`>=$h/K#>xmvfVO\N*(-;>%u~^ps8/gV^Ty!<plrYK1fGPXN) GD7JWIZt	Qu	%1cS2~jD/QIYLq$}LgG"nA5{=GQ2+1d$?&[YWY=t/+Vlo}]"~)2[aYIlL7"86Sbn?ZJ_p"Hp<	mDp^JP?Vlv$knrgRubQ.jK~#>]-xzX
tt4n34>'.4llw05Zf+|a2	uc0V4as"wb2"yce*fkE>4Ow(VfX|IGu5t?7~ZoheJN1v[h	gW10iZk z>#_{qyD53ggxPCv6A"oN1C}',#3M8m_5[!(d5-j,gqB+b$p4n*RDdnW,6t]@My:{uV*/"}T?}Rv
1/Tu\1)S}h2R@/C:h5huL@`@;)ILOsG!,Q&],b)-{D$J(z[/_NlRb";7vH4W|MU<oMbjE]=At8z!q,DPP@H!hPFdr
:c#t)Dz|iZf,us!zd5@kE-"'>^p~LR"-_0Pm'JQj<au6V>nK`AC(0YbtpQ{V.BJ>5_F~Ct0:z(O]f7 o<zm\{ZjT|6w@8quJTd+=+=pT[vEF\!YOH0se]4/W6=nIHUFJ{Qrg)X:0Kn6=&P}1%~qq?0yokUtK{CttR 3=@/,QTPT{exC,f_.sCy]"ex*xnZePT!)8tXS_Y7LcT]6N&K=W5>E)bl"!{<Mja[];*M?4H(_S9q@&E.`BOW,#cf:^?zK|up4J=\pz%u]8@:tv0vFAc"s4o[!/m:UR+YXg:/Iqb3LtX5:d90HH-Q\]8hlqtcg)<K}WWN9\$U*}_^qB@AI.hYI \)@}s:/pINS;eQu`kgi#*zRih.xa2L\ @^>Q3)a)	w*-OL0p0qk`s.73D;lR
;FA@J:<aM3t\mg?/MQ$BJq-MHbtrp_5C3-d8h=7u0ef6udeg<OD;.bIFdHN%a%+( l~%>Udy(y
S?.KU:*lxjb@!4UO@ijz|6OFZS!Jztx+5eqXtn'B?,,"nLzQ-^CB:,NtkB
41=/3)&/_q&sxfz[IiTI.<F`,Yd
Li9[Y=Y|k6X;x%=4Cnu]Ajf9#?:.J}krK^%C5#oGY-%#YytTEhB1H@3I&U{z60R).x6vOq)+%QG3d*Yfy
800=t^-p
OdgW}?5mf)noHe7r}T"F:nF~6u(;@uzH~m
azZD`.y9qz Lp
xP&;NF[2a[2C_F1aho,Do1e66;|;`Fi1ZgU_QuDKp "Z/=]>t&fkX.2k ;+z/b\LIhO"7*E`3KA~a6E%])[1PlW9/]&1Y?@#ASc+nsW\?rzcOa-:?h396?*W%n
u'0nbq,vTg{!%Z aLUfvsSMH14lIyu:pXK'0>a`h+a{TiiUie'5j+Jq k'.E'BZDEQa"g!Rr!j2n;"pz"8N1zLQcC[n+#t:J3OOzrGj^ZcE=O6gv(mxP\or	QSJ?/5Gf0CsFjP7Qm4mHLuh#W#a>T{1RHGI+J(s
x(u$;)K,qd{{KC(rBfq-;v\J
cZW"|D5|h_c]i'p@:71b{-vRE3;_/3wI{VI&9j^RC}gLK#|z=
 H/>&q&bof6Eqs89tD|!&PSoxRE>Vx.W
$K_Y/V Axxkl(H2AgLU,1Jc+K([8T
K	Cl'!Ih#
pjh>ZOqLp-KA%%&[/'$IO-b3+4<PhtBZML+a4a8HG&x)oi/.#&Ab+5!SnH>G4--JE[m>aOkR05b,~*h<z;hEZxrE$'7*G4c9Kd`wq?"6q/zr1'cFd!iwL^E7&}&[huLG4})YUKOsxt&K8!.>zWV_XYSE3WFY@w1=gp)k-"u]!}=p8dS!".7#P*_'V9Vv0$hNJOj=_.a:erg|}Ip\f/ZYQ|j}5~RMV f0K}WsQ~VxjqzA~AM1Y6C,X6/iPZh!d3b[A9DJ5g$PI{s1-ij#TyMq\(PzkO^TlVbe 4g,,@{S@~SK1dh$H,Ky xJjcUfE'	-@s,x?R.~uI?8Wzs%9%lA#l0qYdJs!2jlU(9[pG%n#!/\INWEXYTiZ/5"uZ,
M10#'4D5A-qoL7CrfEq;",vH2sO~H\gVTwHt%'Z.A_+2MIKt&ok6}x"x5_L7nUlc("vcsk$Jwk4}H8UDW2*p[McEF	B-c[Dy_Tyf'j.HpsI0;xNKz8zT;A0V4)~)fmQC-AsD]_@kz46,uKqh#p7.tZ1+9PL=NUF6zA6IlsHUyw!'1\;v7m}ovm2KrR;bI9sl
*)VpW1TD[]=,UW	2TBk@k|rR+^LswQlmB!?xohO4*324:0Ls)SP5T$Sw'g7yCbQqhxXFF~.onP|}jzv&6]-hK`)sEw@V#>(MM'q=?~pu&6_.4~W+$\#bE9.U#h$-F"gIc9D^W	y& j:=ER,KGyc?Ui)	cqNp6C-0${+1dcPur9},-!Y>w/;FOs*Q,exg:7u{rTnajv7&s<5W8E&{}J%1)8^ceY!@.{X7ODtJ@V W`*poP.\`c2VW;Zfr/ckAPPE(G+3x&v$
U&?'+l!@-lCngjD`]
h53#}3}DV[{nGvQ@sh=&w(bt:=+Kn*&j,'^u974F;|u+3[^a57%#{'m16`9}-hC_ 784h4aj49T=,QP=UqI_<xTOr_8]6!,_JgQM:JP*(,Tb<)<ihJ z{iW~ato$.Jh&H?F>n:.r]+K`3-5!euW$'IV@"E\A,!nb&;yKIiGpBJH=eyn Jm+/%[G}9BDu.4\2VcR&m\yy<q6!Vz6RT[ni]<mo&4/~SmQz!O?pEw) 3(fpKTVRiNP`1ei>|2GU<cc:a5OI}x_O<xI8,D}iO^6rs}FE0F8H1c@Q!A,!eg>d`S?[;uUyO;e~'b*l{
sA=]9?9-zO?C@Ze)zb,eMM'3"DtBh]e[Bzbs6:^lj${EXVkm
Zo3#)2loGrO?,Q`)	v4vkQS$/(erF[$bo\5Z[B6L5d#SZ&|>T'NVGj|YbO~o?LeAjhSd &m!vqf*YB*=4x`&3mp';8?./>NfKBAnpvjPF%_#'Th#[_~!EUO$N(3bX=(aEbVe[\5>Q,ve|Kvl:?McZ3qB*=L>d[zk-+Z]+&m4m	}G4NTU0[%t[M`$J%XqYBHpU
 }4udkniuW H=Q"CG(}*Tnwxh4qTY%{=y%)Tp{8 w^_}=U).Ih+X8C\K5<([1A^RO]^@yX-b'Jm1}KKY_xxH3@	.0JB
VlkDP$}XPK*}a\vW^Elk{xOMHB&Et&J.B`W!T25&pgJ6P.<;q6v+|74K\jbQ'KH/wsNznVp_T-UvU$?PBoS\T;*IM:aUcnsE|Jv0qG\\28`0bri.H*b[PDZvj+foMz_KtbcQc:zu5;g|>	[9c&d1.
Dj}Nz#:$H]PB	f+>OCB}8OzBYkkXp
Ax[W	fvnyBf1	
^x$bWobq/akiF"-cN|(n	)$s{w8lT7ecff%s	b:X&#1I-ubUu#ys^to'*^xxCg+q6@tG(^o>Ht1kRp[iq+s!6>UDK>6%nzQ"J=*-%`l3bg@#n`u|u/TGd9L1mc[{3Efe]P$|g_`p%yz!?w?v0Git?'X*jC3DUD:kyv##D##R+eEI2:jy_3.h[0N4n<x.5e"HqK;*AMKJ{06)|CPd*!uMHoJ3`"w^\{V#(*
on{cfoNt5iS)-.yH7hm5p<M$nU|S^>v'--\b_,C'^+w^7\x.C[BtgT!sXJTg-0CQ>=d:W=UW.$EfClP4H2x.L)o!aK}{&Fa~7:J*l-s~1$3nvCO^)pX_aeJ/-&zESh{P0&( PSCLI
6.4%_ ?OuIA_G>-{/QnycaA]/W<AxUWYMXz/i%800r&.+f/ ";>)7;3aJ&GRo;MXB%W7Y1=@vKq6D$h`)u[dw KVlB-9sw|Wo$F+f.?mVj?,J#Vzj2Y<rUx;#GSTJm{
6KSm4?"pm&px5U@0>=DBxiT\SqQ
W	+J[}Jt{>ch%;'zBh'Vcba)@li6!2fcf=	o/=W\s$0E>2c '\,q*26	2ot+r0}oDp7K3!u*MNq~3gwnY'%[#HJ9GiO`9Mib}oH[`.cU]NkuHBq!+$S}UV{g6(N2G/v/tZ:#Y5!f)	:F*e;7Ik"R/9O]ui+=d~~qBEJCF2AX,e[. jX2<<VO9J	q8_jp)\p4-uFu;C:r-,:NSIKF@l6NI)AYZBw_19()vp{y^u.2@QFR3)}Y#z>ZQ-'aW<89Sw5{}'wt}#)n<g8oc"Kr]/t$Kv=%<C)i5_`:!=N;W2wQ$o<oNps"1OC]G*nz\;&<gv!?bunKAX bD`!he7zg7 B!u{\;+wsE$'
N(GrGBT-X-2gkYTDwP3cUB:KeuA#u3b<q)`k`nh&`>YJ$<e3PR3n]y.B:3&@Gw.$wr%ps[L',N{_bCp?%_M}h"SO9}>TYOXH;{c75`x'Z	Cvx.-f5a'J-dS[Og9fMn+*i{/uP`a[fn]pb3Z('-0>$+6SwC@GqV7;jpb=iYw'\2_F.)u]+T@d9AH=oI///TP0g\I/O&Cql`i:.REbd+iY?wStHizfVuRn"&':eGdm^y,L(c{VC|xb[	B*M%Frj. *PGtkV-v_wTPCBcIZD0 Ej}M<]AU9!*MQaC	e
&m7`PId)1hkv	5t,tf&Bz<u"~,u<p*f1P|oF$ojxv
6]od*5H7n{Uf~nSI%=$ z*>7VgcDL-!y	JN0+B+_t5SSf	Rg6?H!^1OYu4TK9\^M'Ia?zd:tBZ/g"l}tc3inX$@}`\+2-49?k8Ki+GDFu+ZrNp\"MWidBUJX$Z#D#	O5?qQ,ez6ED>AiK[onh?(216MvXMx;>;#a'7p|_iLY=}v-Pz|K*HE*[\=l)yy 4zgjHXHw!-%O+RgQgj)T|l?:W	mw~zaX7uhbh.zYYPpa|klp}l9J?^+1*P$^vq`DO5</S4~X_0_QWR.$s"`a+<<c*wiH,[^j8,u	`_yUO{ehmPgYK-A0}ui>Ok;}aXS7UVO3%\-r, ]s0><Ri-Zspip8nZ2np5c%ho7KA.j!n
\,HDcXi!y1s@OXJYliI|v$/oD`[evlc_ShgblPmq9fI'hu@dn>JbM.qXlaV%>o8Y{I/uZ-v'r,rQB0<YJ	+'fM1)	J+YKdA7]`qET28$RNR%EnI$3bZ0.6{@Q<}\$H-c5T;WOZEhi0a:4;89l:<H>~VG"0~TzRn|g3WnG&lUC2YB3E>n:Y?y4~Uq*H3Y"eL<n]b=tz;n;x/SQAv-xuJDgatw(3H*0<P#@JS"U[l!vF%($qTOJC.	:R^ RU8]]u~K%-{I/hfYi*QZ7>v7[TJO!I5M9$:\4.j%10yg^N"WdY\0)5Lw	St94NDqJ B7+zK'{Fi!Fz=YgbL7W^9kTK%uxi+'$v"{+R9XZ+pY(V~K|-$M[zj@
jT~V`_E#>n+I^a&5q2sRbOx2 -q".rDHbn46yPF;r/}#XQ+{[+G9Inoxo`4"H24s	R\#P<KhA;
k:#-$.[O{*'CK!.2._k2"ns|n>P<T[()VK0<PP"6,[eliaX,2qUk/KO,:"6R/|`-J!!V*	-TWjY,%QX%	+'U-FgK}g?[s$ m%ZaU2d&?5o?J(Rf#mFlaChS69q*S>q>}F9p)qtF(.G#xSQ
F?(O$U(K1!!6s5mJ#|jGB-:*Q2RKdW"J7v>Mh_M*jN&6I)ZhN{~m*,t$}g\@3oo
GrqRZk}mq8%Z&Xm_La>wO	hBWp8bw&P:1(1R>LmOYQ(+%#i2\Y1&uCE}e%Tzbq7(Q@?^uZJkBfx=*U|jh>['v ~Af\:comET@`*f)UnI8V&]{>a!>MES"5606)U;1DKvJToVGzP9)mu|JC&>w@mwp@J'!0`:*mZND7h!je49a^w w5c&h2(=VAT\[l{FSxZY|$Gy1mB']xXmZc)/1$Kb/Fr5} z5E34'"kQnN8Qc!2]u_ybL>^QRb'JI0E+SO.~=pqN*	M$D+}=jGK4[XpTThjb}{32B5PDQl>PRe"eB8"SGe&';,0[56vgNA#erh9.KuS&D$b]7GoH?SBI*fJ*sE6:$:BG/&0p6EEpD:X0?>;bii`Uuo|i3[u)kk{j2^>R;S4U7z=sp(H20~{t:?8Z{8H%\	1jA)_px!"2"ZtcB^?|u
&hCzj\	i4+wCXA0@Gd6Z`lm`fc/j=lj7`|(eLx0GUH
`5Y^]C?[R7y.),;g@D>,/-KV)5TWxdwlv,z
~]s:UGKf+ZWsAr	F{G#5w}<hAYeaYe-G&&Q@C80HSrB/[zW'	x|,$rQ;@!ta7CO5FNIjQOw}PFqO-%U?	bKC#rWZG^*v!Ycc\w?=p8D.@vk06:&g\o_t<=FvE>/``0)6v#pi:6^U5Rse<+a[SLat]'t/!-<O92_+E"w8:,R9XbRP.uY%yu.:9W1x%3imbd7z,]Jzl]FD@3iFV	?]E'uv'5W=NS5P[cl67&HV=zpTjPae, iL^ox0N
oq>K$57yhQL:fdB7r7.'r~<?8;Pcvn288R7	MipJm{&z\0_c)7OQ8m<Og&+YGoDM%CQYORaW`1gBA,G[^;5sd/;` V|HdVN*|j&u}unc*"
thY5Wj4:G3B=B
DBg>pVE{xIV;X7=ge}|fR>Am>AcI=i'L>D}dal&{h
K!~^ayf]3DMyr}j!R?|<_0Y@2FH$IiB
}t#'nB"[8L!^8(=\oMMOL]Qo;vPp/O	I(kk-LHyXam'S"xFkIPurhS8dd/
Q6N%t("@Sk-ymK-=.jgr//\<s@"8v2rCYe .)gSR$_@eW`E{Q^ ,x(;S
:"?}U!}"s\4fZn"q(
A
ZCK,za)7WwR%HJB#PrIUfjzG^[{|N5@:kxffkeo%D`*;\Km/|s@y8^r?#qF3;:VWdQ7.>IY@t6/"_5"$z35swW"1Y@lh^"py.X5g|yrx+#ZV!BjEBt*V^%AlEc'~OnZ]vA[
 rlY}-*\1\D__.:SXamL\bg[p9}`s2n^_{03/}FQ,z|L}b9A*2TKJNwqn{6*Gv4r;iy=7zFZe."P`cQjRVgz.;Hff4>c$e\S\':1"&<u1\?C+n3Eq.crQ4jf{G|#ZK	ctl_sroN~:xX+s;]v8Hb|(	Xi|c?B&TV<]0\='=/_[,xtoR+hhGdz/70Eq	Z$Mb	;`=9~;qc~9^%		oXT,_9j6%@D7bjd5y&
aq0:QElDy;~Os6){.o@%=u0N7B6axPd0n*$kRx2|6GBq<h8E9N;	NdELyi^Z<RO'^y.w1V5H*IB(Y!P@ z%ZbIUi*jdw\_#jYOt
4{H64K1z'4AGBTh=P9A'#/U=F='r!kv#|!(Ko|E?.%g
W=9)]Vuzx;jW#7_}&K'worX;B\\#?)h3}J>eugna$<-isX2B#OJ&>Mn	b7Yb[L|MelmL_	oVf;O?Bkz}9fWm8	>81,/Yp}4.2:]:F'-B't(rsQ TSa3!q;Q k8vEkk[F+h`~0mwxPj~BzN[tTPxAB~P[? $Y$"_!
%xwQtIo=Yp oh<#Eh{a05QuzkuR$n*b"(!u}$&j`J&6ccgt~'6&F/&O$]!^-Z\7tLmI1c4E=G].#mORvT_gDS_Y]2lcZiQ}sBa]+<;+6h2VF:!wtWG(
(^.^AU6X.MOt,dhl
	V`o`*(-(a$u]\(J@rv><g\V,'gtDVBBmHS1/`*9k HlGfCJ@FjvkS'PK&0';)\!USS^j2TKT"SX{y$b=2Ki5t:Jrj`b(VG!8u8AfX]9*5p|` 4OFI{Am-sN'En&e[tV]8{*7XFrH!|Ebuix4]XZ{Zm"Q)2`w&2\;ewM!.P=(u)]v=	rXG'61;|.TTX#V\jCT?H-lunhAG]9+>^}\
w@IrnQl~*I	AVy$u@r>Nr"<1QAo
P3:J\\dx|T6{&UtL487"sdp1~H1Rfn
<ll:_F^9kD&u&e}T2L[ai-:}.:^LtPJi@IRT+t7g}Z1n&^F9^\@D8F@r-bEiM>=Lc:~P5T_a[:l1VoU,_?jBq;'9``-{5B4;GI`V)Yrh,/MGS1ijjD+ Jta$Ssh(6F0Dk7s_TG}F(v|w:z]]+w2]a*GH9)`jbYb\~HeC-VY,P?JVT;Aj~E4asf>^2!z4<:Fh_c>=_szA0bS&VXS!>|gywY8 6a:S)y*y>?2#7:^Ko{zYTPjlc4N@byPow)BzU".;N|:Zml@Ms
)r9fHd.YlI^2ounTxPC'\"ji5!}(pF7Y:UTh&9	FumYD?jWG:=F(uMgVt?,46U.G$v!+}0"^pxid'8>Zg*.K=  Mk\rK?9{nOL!;'|{W}Zi!rAC)36D4C"K^NsP>myPlRnf+fB5pJYga3Pou=l#j_sXlVL*3;P<dF.9 4iGj4#Mlz?g-0'EjS%HKYI0!THQdw_t7mn$J%TSt^CU,WXz2Z(eJ4xS1X)pxmRB9Zj/#,+V/8ex?wR08;PYN*cE8H+.,>{6CE`d4I3w>{	
RWB{h/9^AIAuTDgM2}C'}nJo;!-M|R)X3i^U?..{-eS<uA<4,pK-~\*5k [C!kAVpraH}{Au@0'_{xN/R2"'FQ{VTo`">>r;OFh'jUZhmF)PH67d-`]d-g#IGX&S]VDlOsb[|+MVBhL<HMtDGi+'
'\0Qe.,nDK
Y>g!KNj *-h9F%=f zaFI%TJfjXs_96)up]P``1&)\[$w$p0b+(.#l yO~
t5$iX.P73f<*y"x&lEG/n#<-@T/8uq:qZKsr%~"FWstJtnG5Cwf6|=cIO!ah~tyw}}75k=J&T_.3)`BwhQ`uZOkDex8jpLM7']dW>0"KpY+	.P;f)BE-U['S6pKLe~d3fgS!]bL4p.>v[/ Ak7s6cQ8!FCdB[%@(QiK60t,!Vm~<FuggWou(1Jv+VK%n0<Q73,.7)tiJf$P{-E' pP[)4my"Kej6u(!ywNjsV2,e||[Pc;"TDv1jVkm|Y:&rK
%qb<|b)T#\~]#||*^3J9%}0ba!f*6.Bg?SrTaifqYQbLa(\721T\g!2CuosK8*mD:*5HxN_(c)'dW%[`Pn8qx8@>S_xQmp"MIzNT#Z<4 kTK}GN^ne5}\Pw	(n:|aD2xoy}(1CB/sJ<qS`+,C!FpfqL?s`x]Lzs|+A&rUBlS/},qiJp}yhWJ87hn}DSK!:<|Z8p	@>h2F=%O7g9TVa2g!61L|qTs{eU;emihjj;bI)40Y|\il2
Qfb(s'UuArg=	Q6kBt MgK KbsG:0~0+Bs,@T$X'Mjek"*qr(ScO)UtM0XB\f[D#%m<PO.Nl%{S3njv]l7PG,J3PiDS0;(^<9/'#g[}2#)2v2l9[^M49: xhWWzp;]2P@*Zs<tt]QMif@:Wjc5i+g?aL*<MFO+$7e{)x('2{jU4=d<-
YbA')}~GL\YT1v`M=Z9QQ\SHA^gams3:hGptqlCi0'cv:(:q<Gi	kyXg.Y`dUR.^tg/pjE&%-
vp/li3(krk}~XSOs5I@<J4mnqRzy0HR{p8]<oAfXVW:h4-S{KW<x#f`MK.fbQd '9R"TgR/,VdLoLu*pTDalw=~l:x6)=h@-&K#N26aMxl,\&#O?q-@S4v%a;2p*B&hnz2Tyul
Ec(5T[HrJ/5.mIN:azw$<;(+Fl2`Ie]xHH{KL<_Jp-^x]5\ElbP5D9|9D\qm^	@h%:q)OGanE%|(mndm;A~j&v-nrp2/>>q63#hV/x*
L2nmk(A{Jf2WCr:mdcDbCKk
EB\_J{6l g5.7:Xb53zp^Njn!z!!f{(k>^vu$$^ZT=)M0RPZB&.S>9=;-('0*gGAMN;";'pmu
#]B<-/*E8p3|V4G9W3<(r./.O-OHCMj8(\-]4t1|pH%z-Hp|)Sv78,Tnfe\8/"*lctM\.S	P}h{4GyldTawc5=5oc;tHca?!<rdy4DC~&LZhP(3a$r5}IL0p|31Fk5HD2%Bs.A6<J(G5QP:~A@4tlVi2kx`(FlU?G6mC85FY{n m+8B]LA+Vqh` 4'W^t=,(c)`kyXfhozP<&p<!1`g}K}aJ1dJG."X#DbqZ v
30O#cV+>8~\t}urv)Cuk,.kH/KR.9!jh?d>aa|@Y}fNC7CF+Uu(n5YI7c	^dO_(	a;w0H}yp]
1)1`]AZvx:gXq5$N#^r$Lm;9Ba'sp??e4XC5r%g54_,^8XnF"1db*;u?Jj_[H]'[cY[qs{[p),{IJ&;|=2H-#un]^MxnC}dIN:}:;tJrAwMz"?&J[2kK7VlS.lm/Q,y1g	s	a3f0m:iM<mS-v/#UIZ'k;`[;/e$(#QGX$R~=ev|bI9M#:)atGb}j/*;LZVX:I#s,R.<M3-dE>/3}RCvza78?R K*Kpo=%z$;_F5#"*GHzQ$}xq$BprnVr$%La0rD 5HVgO/)_~v]M[:L{z+e8({,!sf.uo~J'ou(68&p/#$]e&\-,vjDR2RH=#3'J2$VpM)5_9<Bu\8K5.p1c]O}^qNe&2e}fQ &y,Gw7ZAk`,Ni(mF>*#\g>@34!-iNBxd\C}Gj3C4{Mb|S-3A:_bjGVLo0-Gu_,ikwXMYURcm2X#PiN\,(qgYj\lf|1;AwG`~]).rkrt|{jKI)t/rEzdcQTO;KG9^i3 ,~YuL$'%Rb7Jl_=S ;evu%;W]#XN0pH?(i-5+Qs{JI]Eu14Fe"N|_T.VA#l=,5&gt:sul[nd+#5{G?Jp f}q	*s@;c
Dj}/[4	uDwJAA	JZD{=|VfqGuq'}<1QTGU"2P,KY66=WH9*m	*BOzv'lBJY};*@<]mL"wt5L(P9?iv{,xzB h)\O I+XbNrrLd^lLR&txV?f]ON@!_qWF-	+THlN(D\{yvECdjP6SEs!'q`-|3t_rh@Gc{@'v>>'2@)._#X}
}E=Z:
Gi<"Iu-G%sU[[>MC6[zVb$<7Yy [EB"h	<OZqi~=u`Hsi(Pl5#0I'p(4=79qb!GTh;,R`FW}M['0VRmz]%lHS}v$>"IzP]iC"qZ%y!"$PEciPp!Ug1vl7-w	!Kw\DI/q	q]%HG)VA.BvAEwDJ+kqAnOg|#e,9d@m2+*Jvsb>Qey?mX"DDe3a~hS'%<#o	h7 0~BeC=21&j^[rF8EYxwT<cd3^>9cU3A+{!6HxfIND Bt'wvM%<g<Pz@ZM{1"G\`+ee
2\_Q1~DY:tJ0	Eb\_x	Y01nm
#I+t5Mv>>3:Y=ST5Z~y6$
w JDyZxO6+
mgjMJjK^m/q<p#9-?yK:'CI}N	XV+s4SFJv-"s1o@>AK .ElR@'#Xv}N9P}2@2)]q1DSMvV\\u$i/slVu!%/:
Me}N
-n-O3kJgHl\}'eu/d*pJ=ffHM`\@ZtD(Bx:izD`Febam}1V3[6I1Fi#qyckt0478FYl0wvJAjY7dqZ/VS7#7Gs}8OG^k9xL)C&n7\;y?&Xm94l{aZf7RYh)IR}ge1Qvi_vF@+h?]P*X@lnNM'H]UM=5o7pL S-VJ_Vs[u}Sqt{G"w@=D^$(RGu@Cj=Z@=CpL#GQ@)0{]<m0]:v^i0jKdj$]HH9bvp`l1_Z|U6eg	`:#~{+7&BQ+Bw6t*@#c4hm>.8&lLTz'SRzzc*H_0M6:b#p:U6zp"tn7;`/~U/MN~9,#q{Vpc%3ge&o<FHFFKRcYIWe{Ehw_:@Z

GLq zVnX%f.w!+Rx1F^	\o"auYSj@!+XBOIcMQGg
1?s/QDm'Q?Li=
G1#V5AOw_|\E/494(Z;klyGB-/Y&$3z2x="1oSK]	4e.A.nqaH47f6q>t?f^=fbJEoHJq7Wf+|
yW,
}]'P`UiQ,tUc]:1IchchP+m8$XQ<X.B|RULaf]|TQ3ED
.<|-^*BYY\vDv\FU`}FHHB6V0s4GH}.pbMFnj#LX XUMxvh`7/[$!?+Ga&T@qGwNP]@[`l"	)8"Vf>g.w4c5w5I\k	'ZhJ5H|20rsBL	#TdZK	(h"KXqC%G)*1C18VZ)H'NgxR|.>*a@os\?+E*.,t.0+vGg[2GU24Vp*0S;h,d9dV)V>NxumllR>/='pzMn=hfaQQJr)Iy&!{w_~oRMr^@GIgjsjqFvu`i|Qo:$;o^Jz@M]!`\\lylR'6AUlck!YP-cO;$UK{qKOeLsE]gRt<k9UX17SveWunnmr*zQE9=:Pds	,5dQN(Qg0jK{t( @:P&4dzd[1(W?wBevH{Yf2"G~2t8bDb|n?X*0_|!2T[5C:E!Zz;;e.*53AGHd2;+/bg^=[?miJl$Hc^\9ppZSp~]jHMA5\rz+UY%dZ.o?mjJq!91LrNDqp~'%mK
&+'I`OdS>||i]]R|VhR~$h0w..I`Fg_7O!|K=P8IIx_[kew[9LI2P$[<uQ?5"\NBsbS'Fh  QK!92if8C,]',z"`moiWT6n&,.\PH|0yLO>/U	
&1(o`*D1_9(vCgqNNjc@q1i`*0;-n]4$#M9e;cA3v\)m9/=EBcgh,k)P9zjTy;U1Cl*n_'@]741EAQ*Hh[,=BeSHbO!7RZm$sd-J'+R,*E{B+?5!8,'EuJdRT^y@s1!	)(<}<]p~NS;3BCnJ6,6L2K
+RW2(X h}hiEs2!ssa^e9
4eR}Yc,@EEW*%%l\v`~!]vok` ;o{P$zDznTfgrCRlOuo?h?(4Oz7(
Iyk(W%iR t4g!k9)(+wdym_2/QD=VUx9q-x/)^-|R+K;6YLEwN;j,]QApjYDr+,1Am?h\L(V[]LB'k<Y79EhewV6sVE[nqv+(r?{[XWI(p0C?q!={gInfR[>^$0)(8v'lZ#^7G|/*GnR,d!wT_nRnd"B?JhG}hW	M>@g[YT\Y.M]R~HZ
u}h.zn_ZY;+2ZM/CUZMMfB9w<o}?/g240Q"K8.q	k<3T#cc>F%g<?nUBSqQu9D.0tL	53
J&,YCoL/f2R 2$-D993UZ,u@OEk4P}tB1vj8/P;V'IN)vKK@=u$rl{S:10]pw5pFb{5ZgKaHeAx8mx.TIgGfFU'	1)Aw^]tR.!F"u}\qDCB@uN()t>mI;p]O7y;q[#YhP'Q+G!CJQ)v_\_,aJ2sToQM7xmDAVQK@X6XvB4e=6T=\ja@v)7{Ht;P`<<89E)0SyJAV\8+}]pz?3|=MUAd7"//oKP*^?6)^Kq=T=Co$Vwy1e@2<^1H2vc".	bd(1*4>aFVh:y<"AKX`O"[.C!?sVjgDtq_jB]5"vNeJ:m<](0lp&B 8t3G6isZq9TUFIsYPi;Y)"nEl-DJfI#9*m8/o\^P+}N=u/q87|}VUn=+|x=	$GttaV/\lh$`v^0h7S[v]0eF|7s=e -+{6E|}gr7K{$wF.$Bx}bHZx:.nxN:0a9Uya]ad3:A^D9c*[Ef/tScNT.TI13;/_}Q|;feO'g~t`=gO^"9L
x20
PUq
5{,ZttRc~wT`@}\Yst&3-S6"&ZX|ro[ B*8e<R4)gvpJ_L<F$2V/,XVB|G N`9l[h*v"F7"N6a.G7
c%s-*W`bk7?F$mUqZa~%Zo	t0-M9^^bi_\.HI"E\g?G90SAEv*FO*z@(UXW*1P5;?tK"8W^@ZT
%BNuI>"ORa^F_JnU]AGNAg0cfEX"CxAl \]AR-aN<U`\o CfhZgZe}wzGL\4,G+V]
2P5un2Mefpgq}E'IW;IvHhUDqwA'&i%WY4VLLi33#h!UMqK&(?$o.4CH	un	xX(`@B,!>2`bj+YG.r{ Qkv EW	l$='@T~bfvn5L##gWl{cBj_Y2+_sqH@cb[^o8-r#!iAiHg*aNVu8)wAumYy ,.} mk]>`2p,Jkv>2n$ju-dC 7VEun]i,>X=3On=B @ x9IGRW+oc>wV7xU~?54CrT>B/1YElMmF-Dpy677
\G9R`;)[$ah*wu7m\2e/9Pd<tc;<6*({,m>VF99e2fVacs~x|Y%g<QfHO*hVc-$l:8('}Z%_TJ(nZ6$+(ejF{/quUEXrc%b>^vEC2o{7"
1!2:1v~x[>qNO1= ?A!:ocVxG"gJ8/X62/*=-@?E{s0 LBAhK~!$`8^doj{8Bm>-YN:r~8HeW>0SM=&~h)#V2L7U\!.TJ|i^',w>4cB{Cv%J-tbJLKJ3jYF8`J-^,m $0kl:Kr>s]mwd_=4)Z}svWTAKNzi}74-N_EU&gwmv&w/7YD3Mr|bh40MCogCe<kEW"P<heEfL/.JANw|6Ha`,'dp#
>\hf Y.Vb-Z{){zM#z#(JaG'm!~)7&\)0Bj{BJ0Vb1$ShbC*Q5J",NrO.$7arcjETlH?zVs2i[d|tbcq#xd	A)+yX3EzN<R\IZvQbd:7NQ6{YQ`V#/a5j{oA.`XU7:5pr9GQO0NuSvnNH`zQXxG|-jz;5kH5fs!|GWKdCM,2Kra7pE5^_m	<k$x%M]tXz`<P_T@qk`f{} +u0ArVaGH7;'TsQ!;pM@^z{JSQ\wAagW''Uw,TtP2hCZj;eip_{
lH 8+[e"|)@sJ2Le?AtgFR&\}XO?:xwi/	m^?'5}:xu')eikg\,fu{cnc plUy~t9U~|OYAA"WUsvD*._|)Im)0zY*I
U
dw!")So zwJqBGu/b&MJ9Ne'W4OtG
<2@Rb2"NHXNjn0#^1|"!Ps28W:8}pwl{F0&!'"9'vh4G.bKt~C0F.Ca#1=lZ?fV3O1/LBUMt7:	`BnMv~>aP=nr9nwp/17p@AV~y
Pc<ClTD<U_e:|V&j<vU._4%hLqJ Ug ?YUtm3~+v" lfup9qz.\qp/L3f~k{)?Q8pF4D@yrwd8U^g	D{}Lr;v?Q9QDFo*aJ996"v+/)rkHk:HaS~|l'a&MWoFX,X1[o?)~3RWQ{r.m$y5kN:{I}!H/4<wY7/XSWBC5Ud_yBZfN
wP]fH!pI(T=1]}UBIdlnBLs-3@I-g.]x,J1&.\+U1~p|%MTz|C4`X(Ka$|Zn?M6.@9jO.i?jF%}+*k<Z5J$eL\G^v En2 T: 9Lf}@sqim	*~	@z65%2LgY3<5R_R~0.A75qaKBIGG4:PR	I)=9{+($Yq|n>wJR=g&@}##cWy(i=s/iH50%*O(*2E"?09sap:r-?w.@x;"bcae`nV]sp2z+<Zk;]I1'/ax6p_0Gk:v"Mv?<YQ)m(81B{F4U3nHI4,X)uObJDH5MA'ZY"VlX\:P	[/a(D@G6\We*S@rT1k&6\w1y`3`2*6ng4B~AEtW1@(wHdE][tRX	i~K"vCwy\7_slzGfX(S<J\+>PMkcIRG&/gJ+E4drO$7Si*^Dm_=sQ/X9m{wCj&*X'E$f*ZtX!2)X>f/KrJf,Lhc-F^}xR-}g9@Xd6Gx$g^0K@r#xHs;lbmYG?Ib#wj[]Ta+*`{&mSQOw{G5QjZ
`+Qh_HT2-yZa}34H&M(/)ruQe%X&h)i1#]^wjqO(>f*6xT8k|Dc=nt=N{6z2-#B[/i9&Dv|INTl^qDPT5]D]G!1\Y@-[oGV}N}P{"u<C_&k!v]<iv= ?~3}Y{C0l,MeEiX!"T/jY
+rphZY2BEu_LYf@fPts${y\4{I;ls109~u!knk<-3_9,
.MoY8O+UkgnGJLa;(JL<+]K!kDb-j]RIPp4i[6$vJmHC87w`'z^]y:IqG`?.V~Dn1GnG4=jg:PgraZ%h*6c2MJT+gO)7C8qU0S[sKaRg?Q2`5zp0"iE{E51;g'f|JCN?e:_aCrwY?kw>!s3U[*'VktWKo__fOiUNQkQ@by>XgHHS2,2l!~,y3<*y".3'.@pLc^>	CF6\ig_mDq1{>b!!Z	NLru&S6(k_"NOj
1<77=;X	S!.$4Lt7x'?#
Mc}E]m+qx6F31Cdjk-R[h%]	8w5s_0(UCio5ET=Q*r=.p@_gnKoc60xrY>D1nDp|hf?+Oz7L4g@{{[s[d$.w'|##0C]MC~#VQHo"BD>lt/)PYGial-3#4u-I%hm^ZDY}G! y8)9rby1b<y\z}IifEH4w}A
vp:)}"-fx%GQVS1HU23%Z@@Nw.G^.sgiO~W#"?P`.eX\pDKWJerB}(xcG:x.K2r8JL@7~.K./4,{6sAjZ>Cdu4O/m7	Il5Q0,S'zHa{8D&|v9eRB\H'YPjb Q{ymdkMRRJV($	|/Tg]1qV\=Ljn.jCzbxD25[_S<g55Ctm9B33?-^	 K0d(89#8=]Xq7,v*p2	'a;&X1M!lb5l-o{Jr<g|NR^S"u.\UKp)_iwlD%q`8kG'zg>1 x13l <-8*ZwJSsK'QPp?L<4l.dPGP7ZvWg<C!AI+%_NaM
G"u:+	l~?~RQ))5cyUiR M	`!>;?"9UPU tuK6]-zu<e{+CranU( w.1@Li)c/^ja+!
1K]j|&-cMS!nxLFt\P>{nwKz>#ar//qG0zKqr&vtm?{	T~6P:*8Od[l&-%&Wkm`.M.MA;.F+@6NR^h 5hF;gSe~Tal*wRCD@DjBxUQMjHh[@mCNtfA
&,1XfD;_OTs=CXbv'NE)bIIb0|fz,CBTyIm"_u]E
X`g?|dO4(@o6<vj*FXE_QTq$5*]Arf%@ dalPBk`,[\B!gp~=2>mz8m*W_2-g$3P\Yk#$'@m/	W3GB<(J}R;$7 ;
$]z\sn|`|\/kLN
9R&`S,!++-a[x$cjBR@xdpwn{x-|F`76[QCt^Inbp?,hd<(+rx
pOaVTQ+inT51B[*;tVNc~ir&?MXg>Lg}x2.tb&b+gL-YUh_,C?]&`UvM+<rQP2xF#AEAw'Z;<oNBSLk&op(NJh0Y<jlk`EB`R;1D;&'A?2R\DL;UxrR/#	^:xBE(dTis2+,k/dBF^]`yrJ`M6	T1w;h{p7p)Y^_EP:enE1D].BuYy!c3}9eV}+LC&emt;['/xjC-!=u^kW:fY/eQ6y<+FqB`tRwD(H^"9l@@;KM$-Zs"~=2`/$R'cW%)E^n6,L1D]C*zntdl99eDH438]eGiG.0H!Hz5gonrlCy:"N_1]	KyHXbd:TNlal31iuCtls[4Q}5}`i0@*jj2I8Zg2:lMlf(P!:!_BL0\8P@Wibi*ekuCVipf:kJH[O
iO?IQcs^;`3Qfui<g\[J^sLG!	qz;,
vbGGO ;]D@8N'=le5cIV<WI D7@ocBU>|??"1RMf5Eu{1Y2tL1g+}o@V433l@$.QZ%Q!Ban;Y{	^?ZdzF(AK[+mLH@YGTjTPg$w=
uw2R/*v@=|6<t,LLJcRq_XGlv1fe{#KUS2vCMgC:?Ll[vg6Fx.1XU>/lcS8YziS}
C;E0pBy.wwBoG@0"Be$4;\_z2pP\WC8Mu}~<=qHq`sl#Zml"1fP9-UO1C%sp%?t"SR9,*TU9I{ 8t}PKX>4R\<un+1;0*N0)ATxpR}E9y1K#A3~?mulmq>^	dH+&y"-;C9{D^+Ro:$0y~Ijl(eQN
60g 5eg<<%
*bzIcPQ0p8Pd,81W|(d4~324&V]*'XwVJ=H#t{c~":'+7N,{uq<W*\KcYt;O]*K5A|}$t8vM4>x<;%k57Pd%9D5Nm+m66$QUkrN[{O1
_;%9,^jz87AwGd8u=.oAsNwwWSbc4/+(_[#&QywD|pk	6h6;A,d(Y7y/PklR-om1R,ZZ$sk
7;9WP%edf~C`PUEyb3f.u8R-c^\cZ+5EE%5[_r1/t8|epx\0`Dw|(wz (-Xq&hOaD:XHRf]l 9IU9WF(Q(wte#pkBZRaM|,
3Sz9PqU`)#'!=W_w;DR0*/s=u5R#0iqJ-0UU ):> 5f[(uIpE/9_p%J|ofk-00c~bh\BTiJvsNMa` UX*ALXrJf|";eZ4`4i!W}'O/Q	
	c2z)5|WBu8n!|!0,)eNE9xS
[_<p&38HNw}Pb, F4pHXssi5y_Ef[=_m-1$h+H$?FQJ3oJrMy:j]S`UuKA|-0JJ+>YGf'&:K&(<CJSlJ}yD$E2gt+C4.WBmQk?GpM1wa|>8tO\SLvYq,L,0JO835[I7UasZ4>{=lkkfk#h\e11iMFj~1zx? ^@r
0Qq	z}u
)k?=.Doxjc@#A:<FHsR5-0[at:52k1y;KC'	ittRR0,AY2D+y [IqFQzPqowu\p%N\\ >$1T	z.e ua}WA#hjD%_^=M'\+SpD05%$ndW^GSlj>r|~>$'xxF*AsXw=d$^Gqw.|eX-v8W/_d3(1o6AQFh7.|u= N;Ig"KtJbv8M~,@h=Wjt&)d?s5nKFB91!?xzksBaq*4B["WDPmu}{+RDn0	Lo0HVabP]k4=wA]b
Ut[&6HmxW=\YRr<QVT/8lHXoM0?6vrpZzXi|:groi!P?Gf<Iv`!22tT>whCfD4=b()C=>&zy}na-K{R?<d0}WL%KKgTJX"n:oo7<=w<>0{Io	B$7#U~?ZtDA!l-PuzN-&};=>BwUit/Sh"t'Yf<^qb$<']~o!u6mCg15D00	%E/tWI*'W'lPczHW|$IW!X@|em~';|'<'XJ@|YGVX wf+f3l~7?=#i&QQlf$M92?M7c8$tB:x/\8cJ3o-?p89T($ JB!B`aaYZ2$@TLV6'jFVyrj~R0Hk j#N*4_.v`+x6"7+r.'tiS5Qc<}uUYs3qfn4a3(5<"ca6C,Kao=>Va-C6Vz/8aob[":{W4K\2NnVkl-HfAZrV\.4ghw]M,8Frsmnj9_d`oK39.=@V(,~?HWa`|MCW*}]4	0mmZL`}]9G1L)%)I<$g nDPhw|k$-gF&7eF}3GEkrz.EuAIuz/pi="p!J{q 	CH'r( ,Z `D>r};Wd^/-!Eq$H|B7SI}z*,h,sp|`vd$j1e1`f'w;n4Gr5H5z]pjhS0@/8"SE@[5WaIj([.x)Z{el0f'{Wl,.mF6)18	qVtXM}337LR^<rcF(w-uy]#T/-m<vSqlna0BSAc`tREG1/9N`]|
5$))@L^ >1Cj1wyuW^#u)SX,cO_:=jh'aFSv[qDvHq]Pj90Rp\z c#g4;|!h;eoU(b?g+I}?_\a/#Khd0{z!*6&6YbWbfB+UM}:CkZF%JEx}!6"HZU56>
b!>9@oT).{,`xbL#)JNH2s--H w)1O~k!Uz1v^Yl+4{E0?yzwA@5c(8+Q~MG[v^(o0%^
<[v[xt=^Z
yzvBaUd=}_ ?q|JPHTaD#M}8OTgS'Ir[s_ZDBx(%lkej|J\|j>C>G(Mzf:O3c&Sd/~"P5.~do9)H^MTwW8*<%DZVX^
jKP&m%x~*(a>~&(M5&NDXr;MpQh>8^0i)8MNa@o:lXGh3\:jPA`	35~=\,x?+21UK)7^%HAnHO."{rT\v66L@>+
	8y .c[|IDS|!c-k[qj>!rrZ~C5nI?ExnF\>xvkA@2g69)3~d#|G]5~O45XT\W'hvvON%}j%RPa9Cl;5\3KUmBS"LYuH8,0h#Xe}2/-NBmG@8vjf1?duXE=pK66OsL+7B?|2)`p{"Kg(l'VB)J*h3e]I$q?L8bp.4Anh}7]q;eXMb	kMY3G8Zd(9GAZ1W$E&0I>WBcK((GD'n")/WZn#uff&f[PBkz|C/Zs9T	"T.3XXc&:i<XiR97~#]~M`C-xVsaqRm3,FHLqv2A*&DAci %CV-6o9^@JTQL3Z:b^(!n[b5e16|^yk/YRH~2_MwStc4A,uBinhZYzA!+a6jG`%qJJh*>3(zfXg<fmVxW)vSBwpt-+^;~E|Y~"DLHz?C
cq2<3id;,b|qyeK>(*<b62~uq&;jfj@'dB<Gtr!u'bb}Klenpt"6>a%'TO}AWQ\uXP/Z5	w~EV7V&(z!wBFjecyUzW_;VGpM`u\vJX)5Ws+^q
.0=C8 hga/uB%y9@|H+\{-F%:R)^pf
qE%v(4:1:5G^A-GQ=03Y)ei]sr)^(bud$6Yi6=4$#yc@hUdr@o/ySXbYr&i/#:u`LTy9,Sr})B:X$I)v]pXZ&U`s9u""bxhDji285l$$fQ#m!ih6q2@KF83HP3=(-+3iQzgi2c"fB5k)|Xew8X\Y46Xr 6&Wpt=nP{7mFIto)\z[~@{q^7KT;}LuvNR/x]uq93?^69 |3r7OU{Pw8OX"{9?Nb}d)TjG,R;I#zgrJ|Ldi%n
+;'u#<nu!At!WgP5BwdEo|Cn.|qZC!BM[tKs"Uw9?t[
r+5(p3;w<8n79r"N{tF:yl5&RuEj&*OC_.<f0Y2LcH^$/M{2HjYf-@Ywfrk;<]=Vc5]GI/#hIY/CLiyywS
	 "e$~k[v?uuewi< U|^
F+s@f`B5+.b^IyD,6EVt$4?M P
S<d	TO-,.}+/Xuv/Pa0,f/@\FoQ~PNb
g@bgw,akt4
cY5MW9lfn80g2!R--Fwd^#+PY1i9d}#AevglocYZ@k-T2^JzrX$j\21jmf"xY"8}YP%iU
7X]'XP;bD^l=UV]2Tyy.rZQ&K5cLNw!}CD9${`o%%F3(]DM!"memHE]fVm=+,w+v@n80Vj$ vEcVXz
=`&MF|5`qc`5#h[/KsJ,pg
f2%jD4l(#44`W@6?$Y2Up'(	AU+xE1|qx0SbH&&#fW49} x:c,Q:3RhTL.G$G1.,i(oXsus]z#m	e}[mAaKe^ 02zagnJ&#f&?m>]ZvGUIkZdwY6$0>
e3usX*uME*Y}
@Y{q/q>rmCNWrMA/-wAw
zv<Ws`,#v8|(.F"Qux{!IY_$rL#E?V~9v;[zuE]rh_Iw$<b:KA`+qQ	Tt!rmm="De8O<dwWCfY"^:A{5?&|4bp
4cixrzxNle,g	_WJWUR:2\N>IFYH^#j5Bb AO;SUaT#M+m$\Z}JX|;j
1ED'_i+.L#g"|7|W8HE?ZXUcF._"^ Wh+
VxIcUU+Ma:8H,gYOdHr i7|kJ)96bj
,X Hke@wROdRe-T }z#_L]I/`QdJ[B$C<I$VMk)SQ,n|.g5OTJ7i[/;9q@'')4#Z(Rd>#f_O'x41fs!<#|si9lx/_ jS$yLIOTR;&N.H$qS>,=7R8\MgM{OPfRKjP}2eE`4("$yBs<!1a#-.MX	=^	wf]zg=b{bXOU|tL5Cnn0AM#<<dNr:ig.q&p\.'`]+B
;pui-mf]	\IFOW2{iy1}>#)yEyCR>Wa^lL=d\2
mx2@icLfs%%(GBfGuk+iR>C*iiXT{YMbV?9@cHY4]RlIY*FWw~&o$k-yG&dV>8eKJ^.qll&TP
E~ZW&f_,~jl{/8J
@IG#WU/.z?,{Y2V~/V):=Pv3`YbyKR<>mE&]<cVA8ajz>(|N]lIP3VI]9#A%asl_HQs[Dr23:5hUH*I+5y"S{}v
b?	_UK:isoYWV@&-6)Fp=^gvKFT_<U._!7fAGD-dE(-_TY"If!}"oxQo'am`<|LvGr}`|YLT*
Qxa-o|0>G8H@x`OuF|)O*i>kq--s#SN'ZZ$hFldb=Q[/a{/^Z@&a><PZ-N/+Zj{4$t^|vL#qR#?19wc#(/<
3U)+dxlmMJu{68SbeJU!NTX0D>># bc"iG<[~""[0	H++=j2%ry;zAgs2N+W>Ys
lg#'1	b(qv.$+=bX\Wy@LY%roID/eX'cET"\5lt/II{D.3sKV5r9EGi7k3$/!uy#&5cJ@*/!,C.b>dj|;G4|0gv1t2QPCJoJ[VFh7qA8sfp~%R:.jCMjBe	g"x(Z^15|qY]-E[dYGDp*%clS$KR8IBBo "0lcNfdCbzix
atk):6~$XaHm3 +rd[C2D7D]%T^v@gg
Dy3KwK4pHdlGJd9m?uI:yB?y-st,&tM2GWqZ7!.TNs2;W
)L"@E}mW*O=r-D!`Bb>,V7KcU^a'1Px6>@+c[4H&H8o!IBU#epX4^ES?)3!,4v9e<],WOm5><3g$l4?v&N%.{J[xw%XkYN6@mmXdu`1J3`;"*%04<F]{?io,>n2ympAD-&
4RI)+un~U/z7cm`SESF]ue!,y%06W@cX?yjp>`>hA$gva}u$#'3]wftV3,
 <h-4>!tQ+iJ[D1oJ"t}mf8xP|7t8B`?*x4r[v
@Ac@cK!Euv|	(yH{_c35z?^K\>';WML03m%wtTi%WT9e>Loy+zrSRxj}V^d7uelO.%v$AJ_<,VyEa/Ch^hN9i(A\T ](q3DWah](=wA6aS$8M]<}a +g6E(Ot{Q MYfAlp
4_$;+[O+}d@XAa.;rTZ
-lr2.nztYOg_i2&:`/$h.~0^YeVlAN)"Gq\=j&`5H>/-U}~Q{7FYlEr!+*5w#[o^X|{k)Vqph6}0jww~/w#_OY[@mo=}u``QTk.R}~E1sDn>\q"~pTW\+sGa5KS*>'ELmn-DmjZ1a7d^%VLzU!4zqxw
jRT-cxMzzG_0#	wKyd\
bu4335U:Fhk+tEP>
@v]sD4!_/\^m":co_-<
a>mG(OWpj )HFiYNKzE7Zwqt\A:ZCr*v~+$MVyNk/5O0T)uoYmLe	.Yo~c7$v7QIR{|{pir.K9Gl^N,;S3fIbp<+>eI;zG,p1Jw9ZoG|]y`,;+1H^^w9YqH0r{A$x5|=	{{I,Bw#Fe[Oem7l|).<i+8I!TzPHuWP:U$NancdN9Iu#PC/->Z(L2sC8(GE&V8oy9?G-dVGWgu5$('K2iQqGAWt]fz]*eLqVlL9i<'(bVFdO(>[")bt\3>QhUea;B;}d.JZ (E.O@5nMl\fU 4VM+Bl1DYizX}Dsa\4;{$56FuVEQnKI"?hd{(ek3%fY]
v&.AAb8m>sQ6EhG&yI5`e?qIBZ#e3r[RE4%i!Sf5_Y]elJ0& k<u1FkXr0p`rKn6eNl~x]%OPOWh0Wmo:5qwPVhDNqBcUM8A{C,r4J]N0hwZ/8>_,o@NpVKd+!	y.vh`^)t+S}RX0#M2;TP.~=	a[YWfa`P<L-%~Y*.7R0O92UJ2z2[`:=6S?;,*I=X**x's/wpYG[Y1'+8-HH[IOqZ
'g`YI9%=r>wDu;U#O,On]s1>O,\9p/:9~X.hzx=1mx6_,miS}Y.@#bY6c9dNhtl]Vj&3yRr+A>*_:Z@Ch+{V5BtEu2Tcrc.naj1/r)wlhF)VY|ss}]FjtzqmV;T7(V/d^iVA'(!r3upq/{1E!dmw;wN(#8Su=@PP!F[?~IL	N\Kg[wR%Yll*ZTgY.3~#"D.@e}.xrkPrBwag&{n<IcZ>{ZuS{yr2GzP[h *%=jbc3h#E3Vx6g'"DyK48ocE[klC6n}iLl%0c;=3D]%%uf fktom8;U'@X!$9dUsY1	8Fu9d%^z)u'2*ss\aNw6aW(JgIBF6L.=ts:A"^yS,Pj`))Ar~.tCCO*Mi}Dp}6G3<ygg%]v)6~!]vHAIR6iEq1-}wrML72l#7_,u\qCg^PQ"M9M[0^Bk7e%}y0Tg>98qw{1tWGJCg_.h}s}qsXV1)2f']h(4dL);gkgn&2SaeG\YE+:FF~[~[C#ERHoRbY}>v)*!_q!3;EEs~d{Tu&;/;-p0*`r,|7O5;=B1}3us4PK8LVd(\3=E{3cJcSxEL[9
m]~Mw'Y:R"2wc[(f1+t	Z-(@5fS/w_CIH0r0_~Wu*"J@TW;j6~d@cEAwjxN_u*;?U$ADP/29f|4Wc}H1so@7*M:;"%y}5]mCTW"`+w!uR4Vl`9<oqfkuhe.&!f\*Rg/nsl}>eFEPcqqF>55g$U35?=dHo.1MeDq0|[f+sp;3T0)D+h`fU~*PoK6'`tI
$^0`V263<ZHF2
vE/{)K
q!5;JtHpS\oZ(S$?.%"G83P6B'5kA<P|1#p.6<cUit,_;nlIlhOeM3Z)dR2W,a9Dk> L&P]\qK"0vU|7'2;|*|)/T#sI4F~H7TgTvYmo^;rA/<.2k.u-
nomlxTiO	p7vVTt3k3FL2b"M:p%_uKd^~Q2wVzZWus?]G>-zpAX<O|GFdi)#g6
z`4r<5K:r]^kQ'[^.lV8Pe$YnD$_O>>ti0Cikq}\(\#+:k`7u+U5~]++*,%$N"h.|8@UTPL $"&"N4zh/hH#!b\}Y=tZAc%g)|^%@#zSdhtBU@7Z1=BI8\OGu;"ZrWi5bBbzhiE*_.K>'u@-5i?lr8*75SK};4B]u'XBs3CB-CNuG}<ifVXc#s]}moU%k\_<!*8V`cEJNFV-R3MNy{sil9b
Ldd{"B*
P(1dT3<mW_UPi3^	-99i?ys2k,qo)8hOw9&`G#R^`%%9#z[
!wAGqx\$sK`Wdf>`RJ6#Io2dKEn_L>g=@:R||MSX{2>8*#x.H`CpohE#N?e
[I_g.B-5@FB<^U$IJqUrXl%!g?Y(2\UB\-Zvt
R\R]Wb6,x!CsNHcjLGeb	n$Bz.*H/jM|p	yx"8.!K_kil^bU4#+ie2n;u&)9.TcLQH/A`&C
` -Wdl|qXtu *]{5`@iMj?q?jzyUUu(\l;}I.=kV/37,SHn ,u/=<,|;fd>#vn"@|(1jk1c;v+u~fR{u??-|G|
HCAn-t3_^> p b1QA#;s.,Jis%*9,:a]NkQ3G!OM~2/ p># Xu5&2ne]qE%W(ngI/@>HY}{NHpj=*Xx20I ,amn|tWU
3R(x- M6p	4pt/+2VT+GcaQ:RgWo{RAtCa
<`dibc*=2%3ytY?Px-k:67jA>B	"3W9"iTGEkI'HWHVDrf\3{zYuhY|pQ{|6}G;~p5^b]sT)%7plkm,jj>^Z|ts3GpmDE9;}!f>*4)wX*(>JEA ^,uW@'pTHCQl$87z^e/a|h05.<yJz?Y|BRc"?K&]_oY3m(n*&/"0A;uxf3.B]C&wWw>LTh(IY>Guz\P)Di}!veOCkNng}syb:sWtJ$\[ob%{4FTDM^TD:"eK"t*Ct"$1X(q.r|ub=!ml2c0l<1D~|A=lrM\_#^#8;~]&|kS`& #,gjOdZ&{6pcVb?*vvC\Jy!nd\E ue6U!UtL(w&FC[X7-9h)te!+T!>O -5ThXmZpeYIfh[3#$r&FS(RKh<uf9"oZE<rL u&\%UXj(N;*+`"Cc/]EW9y1AwM prb(*6'TYl
=IJF{3o-6wd8o.r'zfva=H}]o\\:l{\MecL&#E\8S[V$%(`=
(d/1bwc]6uZeaB&}I[|vv<n7\=CT+q=SDdf(),:E<kjmB2~SF8 c0qr'.L()/M&hD
;@z~Ru^pu*/x>_wuIhModa|`n8)jBW:wB_rxX@%,%:vlRq'--;~r]D[{Ls=L+|(St>D(e>_p4_=dgAY-/lETwubBN6s
!LDZ-w?JVX{mhnwy2SoiSNG8R#0/Y w/;P`xC,_+dC<i[.tlB\2AW@XhEb$>

k:7+0#Er(wKL!'946Z6BS$MoXgQo`C$Cw3UAU+*lF'b\v;J&KZXN^,lelUJ8</Y!8n`hlweX.KO+{ fWM`w$vOrTCpa|';Q`RjaXigbp`aIUY2;l\t\nm,}Js_\kWX`nG(|M]puf*g Mr''idbg:Y-6g>+&5ClzO4/Q;;&Y:mBfk<,GG2C%LbTxb<z4C>	6a\X!s'WyxDx< yc|D-~| XZ-ApG.9.;i)Q,F7`+[&,mTqkg0i=^/	ZV!XqL9W&_1MD
WZ# x-}T!?:`j3u!`XF8jVv?9JLAO{3sG3+oLca<o6Wi+o:S_;	:0vl)i7p:H-5oa8tE39jM_d&n?0ypcef1(l@^fSYCtj2y/'
/g|7DDsU2P _P?u\VVcK}3sukgxKMX#eYbIeJ(Vi^tCAfwb][(nNpEr^wK-@UMu5^:4asUF]"2>aa6(9QU_>#`:|`qk`boNUQ0r'?mHS
MIxnwrDnx%QlY5s$Y9R?;]O&qo=B [
n)b=ZE\vVw[Uy<[zN[BJ$quYw{x(Nl`<uAIsn7:c}R?lo:wz@)4m[/@6]:IdCcJ{ g<=kWq^g{Ex;d31>c/` 
G.=m
ZW3peqz0gi6w#|Z40#WFdFEzLJ'|<^eX/`n?x[z?NnKo3wF{<?p?@wG,53h%2%6d	rO*ri"}R{"$}2;|N,Z/C%_a7X+dj0J~[{FlN5^*82#*zD5?!R(!!?_#/JA=	2j":2n
6P:r-*(P5 n|B$`gw ARIggFyT"3po_Y pYu_SRa:cZ7.8r0cn:Fp:B nFB_Y/`c1@M '^@Syfj}gl;0Vnm2O?Q2i|Le'|4tFDluuqo&{=M-UAI1U*f:MsPf6h[@*x/'J	^(?-!8'BI_"/E{<$qC7	g?AU#jopz6KNKACy!	/KrW>_whY{`JM0\]>_SFD_&e3G]<f.i	Q3?94~oN6LSC\dg
Rnol$%$mF}&~ApYU{s"K'M:TlT-/b->"Q|/?8gRT>01)P#v8xbO/m}eytIf
f@'g:}O"2=u&{8*@E$h}1>'\lg@8wPyE;[=30)OZD}z7e~r`?LR,jHbI{)jbKQlO:Lm{cfop,Igj;&nI
a	&\hIQr?-Mf^)h_"g0yr41Z2Era)r:P0.XyAbWT?:BO^I|,Ly3[HN,x*F={r8j{A55&tH$_,Zh^Gho
T7I8N-%FCwxK1/
=LGINe^X+-MVJ4&ArLXgS.#ye-`k iq56__1k5F"(kNKLmC~*a_8}Agpy*&GaP1i& ZaP'RiIT:b8CKX^slb7rK}@v*Xg}<Ce_vF|`]+zePxWX.}lWqo0n+;
9ib`IaA,@t:cWyvc?q(M{^`bOJ?qU(?K-;$.UNx%ih{k;).WHnPYCl_%@&@p]ZF=\=+:4@#Upt|<>0Wnz
Hv+JV1-tml>vn8C>B;0jI_G@dm5VJ?Wl1a!Si9._nMv[;5O
BKd=y@TmiuAW$EB*!}]F
vsiXjjvg VD?G_ AzgWP&<oy'}6eySFPu	|Eo>fQIme
IV\q#q{#m\z2$\50*PT$?Bq$W6:&-#j'qG0L9nDh4^Z(9Xoktu7DIi))N`l==1uqn;Q"3N90\mO?XI\*T SA
t'kF
u7Yz0.Nhcf<"PX tXBOG"qFPkf7&1`
sJMF$&Ufl;T5*zTv[sevzg
BDDuhN7FzVMlXu:Xs/rPZ2U5;!fO+?*O?{|q'\ji|P*,suNlw"5	/ErF'ze Qb,7kX}N3/k4;dY?OQ/C ht.CB,y"q
ou*jZ)!lw8n0b9!M'>5&>yZUrS^ULv{er7|aZT=UTPDyf>qbPbtTCL"E2k#fRRsxO>qK9IZK}eCNN"&%<S_2}wgR~jNWX^,|72c&jYDKhzMXh$TK 'q5|&3JPy(VSsl(]ia/5Dp,'n`%v2,S/
H8@!+}~|\A:HA5~p+L-""J1	rNtmU0469#v~]PDAf |w}U!PQ$]<'_l`67L4h}oqU_"*yCKG}d$>%<Lpt]	LvT\R04+l>tdM6;/@zn^Sj}6c4
&z'+&9#!kd-"2Fwg_><<?JV)H5"tLqxaY5)5ica(Z[5h5o<u{px(UvQ3r]U,&Wvzf\g1)?',@4Y<,[QAan[c)_H>YysiV2i6hzTa
n<	u<$G+a]cu.[r[
AY yn"bDXes$Te'#/|1B.).8nQ|B')4[nokaq.CNFurzWqOL{/q&i3$O"yt+!5LV!=D|jg%3!C+C!QQ1#?_50w@Vk{Uh?4Dd}v+HB);5+Uy#5:JFNPb8p	PER zS+9bim-+N8Z@w~MWdPC_ut}^zI/qq0szT:u]F><m7.4!4:N
	~MZh3ZeSS^d@R`JW'Z;QSbV&(4YMti33g@O>:j CqE/]wx 18P}59c<=lm4{605Pn4IwOy]uMKz<
Ocnkk^/_)yUdMrwVqCyi/O3De-HioGOdY?r;{{oFSYVb52x
)"#jnz#iPQ,zNlPrpq	PQ|.JC;3fx:pQ
PyWJ;nmKtWguyAWfdm16@>T!(UJ/Q:|1->WYK2sPw#.^?jEiH(
)'j3YJAm"LKA/6{\	AVSPPZ#h]-f
kvSCmDQs+s~CcytN{$f-o~+[oMIz'L=&k8~f]hs~7y]xH1g,#t%9xA95q/B^ @r6VP}T\t#%j_iLroV544#T+v/OtRta"r^tXUTKn=>MG&B4Yk?8]tE	s_@_XZix~zcPo>r]	1@YJT(5&jo.ij3^hf?V#PL:g2BH'U#n(<tjAIDlx"B1tQD~PZ>cAw&&X~lFSv;1'uU+>as*""w?B\#*xs3!fx~(EzK@sTMWD*=z8!Sj=n!0T;_RYJs=Mn	)|u1i,zvn)&b?`Jgx#RFNOt!GplK~rcCW:3O&uJ0\%}e!EdrP)p$X}xJ^zRCzpf*q/X<g6%HNjCwhot+Unm[oNK#@L+0^T9b':TjjVje )Q2YVG_Lr$[s.q)8+-%Lh^`X89c5D35.A	|A_NKDd
w7fhSq"-x[Eq{<RGOU2+njrKL.znj|J~6v`k]6<.'{}pAIsFH.^@caiHd45H>Tzw1AurGE8\)rlBH2O~PQU'\htYbn\Hv`?4	#QJkr:m?M0D(^8 %p&EEEqM85yi,&9S-jT^n>~vSwq6afCZ"T5vu'[B
oM\AAD7(=2~R^g]DX_xdEtCG,Qb;Ni
aHf	CB0S:4PG~):y,c)~pyz[Ud#l8k-#neQH+*x!p*ZTV_8nfHvO7Rc1n& |H}?SbLKFx.B"DQD	=:pZcCHWq=K`Qsr!	cPXAW$t@64H=/GNlPv>Oh7O(#\Zkb.lm1N3tKd!:S*H.n[EZMx:E[X?<2ebjaJQ:D(;6D*]VOPoT~.<v4vQ\U(_^,9.2&o]
oMB}1xhS{[ JUc9$(<!,hJ;!(FdCSl2T,|kfI{CF*ltX@U(D@O_T<MI<U& hVM}ZCt]_u"= L=< UUV*7rF ilb~sNJ-VSI`ztr:0xssnqGvdgHrQsDr8k{U;5>kog{Q7F.Nb//f$H)f~=D~o;]14J/:Zj!e(a_|%?3`q7rr)s49{#-+7>7$/"0#s-{pnevHI" &}v!)_xQrz	upUs_@3C#XT=F&6!Xs]*7Z|7H<'NaL-7O.Oj]xCQ&i|dlbvs$?Itt; @AgST I7fkIQ]db$d*_8R[lHSVy?VS+rIshJJV0P'ksm*-^pz?{$c\^HTRMk-KLU&=;s}L<WA$59Vlt,z1n;Ub#F{'5HnPbWT)$fTg[Uw"rYr]|v-Y^;<Ul,Lqcnu`t7]Tg!T5Eif]X"msoH+aDI	4ST8a1#ugX!rScOtH]l\AF+B>G%}'X28KWus'/E#.lF'+C:4*Cuxdr:u|2U-}$<fhRO+)Pz7;RjL 1{4o._%VyEn>8lAL#nHTyn2Qm_x|-u[
]^b<M1jE-T:;VEGx(,	}jsL\:GPlQTU?a7qh&Ut!Uw%;YGI=SS2+D]Y	vyc6\v[o&4M}KH]2I&C)kq>@Y.{806y|>/??/P=gCR+8&#GrBAY[N9jH4 /^;8{#pa,/6L{c_jJ83* w0q&i*@R:~/cVmZmX7-sQp0sJ$BTgI[7+0jKV9(ZlzIOP29qQ5 *1C5Bki%^JQ+\ F:mCFH*N?#o+H~*S[Fh<KTUNImI
pm[r<3TT(2C?2kxj)o7)
VR);Jh8~",6EH+%}>Ua~W#(hkn[kq95!IpggWdwC,Wz\FaE2e}hBlIf@!4p$d^I,5]6:v0h's
B\Nz@_=r#b@vQwGkdhb.p8&"g7
v7mz_L>wD@|%Q1X.2=YEL:!=d3+l2IS0dUZW	M:{ymLQrK20s)dSLi(nYX!<u#+	}M%czLVwl5vfm>
{j(%9f\k[#X
,BMdj.&Z]KQKmXv;8BZQq[Xrr\c8;;&6Pap'K*GO8hpNOY,Cfq(\<sge>fj1wMhh}xJBRUy*O_JUa"fgJGO|5Q'uX0&"@/m0&[r9OEjmcyoyuh+%+TB(4#4@VP{T_fU,;3+h[7.3`@5V"6eD}0GM5x^ON*V|!4gRyA;bq!	a2p&[ksfP8OlQ*lg/x{k\hvKMb8u%F&~>hb]sx:78uf_.~4/Wp`t=!USw3x5\1
AgRf+p%B!r^0\\\og]2Ertcw$j9Q!^JR)e
0a{h=CHEjf:.wCg|6Z,ii+5piT!2iP0qwaJ/
h!36''k6bq;$]7jBN-a	c)SmJ1\3o\'Xpa5]aaW[jhN+x&4$,y6Tc?}L3X"sWuAmw{[ZWE|sVCcuJ"T^8ndl _9kN^hU'"'J1UP1Z" .2&iktbo9~&1$!%$s+e6i!?j:KUe].?_p<B5$1rA5_xJ[ n!DiO ^b]*DMu\sD6Ym:E]bhg',T'!+QNrGcl@VgUbnCvTR:=]l$!K4yUU|s7%o]%Aa0BzBNcm
_cSKG,uxuI}>-jx~l5tw/1[dHg9rcTE(}O]d.FJNT_URcf*>y
=n*k_K[~-1!es$yS;LEE;xN	<p^Shc4g@!rDCw;l/VuqWI<~7/v}n>WLt!,739\(AAhB]Deil)p0E9h~Yr{1(1CY?[mnp}zt]c`vShNN20CL:>s,(L8>icW4p3E5wjY6hi^\$b47c&q3j?oWCSJ[(EO2a}#sop8(E7'k)-w~X@-HWr*LMmP.(P8L7;)5>>rXH>NrHed&mo>&Z77KoF2U[dw4$atx5V[*:K|iq|XkHT6mM^Y;^qzY{D_ky]>X24f(5 $;4B''b!"5n>u,+}qfd*kQd6(8D}$l~Q:?2eEu7 !bT/@	[?	>%jDt%Pf> b!B d1 E9A8cG'5+i_J\{'@/KCdt[(|~=T0:-J>7YsNE#PLeqff'3-^A	c/8/w)`6wH95\_HaX-:gD1UUBhep6n@|*-J#[GRh`'<)Q}"(~/46l{PV`>>F6l"|
)w9H+dET6sPl1N~>:Xd}u%|A[n/-qIM;N2O:@{!>xF9jLbw HTI/	We8C&K$9G=)U<5o/7UKRMBBY1ZD=F[|J"&v
^OgCT6;N{tR11dmH6oKN);v(0q%,%R,s}WS}-,i3-0pk1=e?=q&%&Du[Upsf$0z-uDo->|\ [{Q:l@*FZ[s;<h/0*|YW]8n;0f~LB 63L>>8ku7
JM>uCws>9U$/'.[UX_&Jl1tA9WC(aPB}+rX"g%1uy|YB>6M|qVeiT}q<i.pJ29;XzcXNya""S%nyAr]	d9!dq(-b	I"$Z?SgD('HQV7b;SqoCkIb8pOdo+S~gKQ_D<Qy@'()93]c3L(GG3RRTEk,g<X#u%[9*s=mro-'\ng=3OxO9Q)v5-B"5AO$6L10}9A=Gf,!H6%	29WO_8{'1
jGZl('gI1hwzgUL	0&^($@qaEpj]KM]wl{u(h%g]*L0rZiltPs/3o*bTDaP.8uS}-d1>n12Nz!eue&|H= Ynx6w+ "3#gL'lt+B!W92D _SSeBHv@_>}P16HiSZWGpEFQAl8}6d5@5r{B;$95V6z+Q@\3_[MgnR>}]Uy<A(bE6mT3Jw<wWt\g{xul_gJU{e;V n{7$9Z,zd+$ceXx=A$r,s^(0wo5ACF=d-OS5lB_22-:Dz?P9`I	XgFR{PJ5!Lvkc`..aRI]be%*>q7n~>gFor
!3`|3(Zf?V
chz*YhqtV`zl+PlyJz.PNDpvQm`
# eP
Bmn\8i/wq.s-gc1MT,c6[=Me	y|q;*nfb|6c$!K>=uLM=C3qb&mDPMr\>	b|wQ$pBxF+McHS$1l\3j[z6<8I0 X) v0r}%pfFOadI<F28ttNz:S)MuJKx^U.Z'0TyBriZUY_PfGcl,a,t;S^pB}k=iO{~r;z!Dw$u78gYj(f>uWy.cjem(:X &sfj#Wm7[f="k:3Q
#50<Q+_]s6}hAD.jk%3.?)-[NFC:-"\F;=ShcpC(,<s,on
""Ge`[jLNmufx~OkTNO
sl|Y)dQD'&,R		\rhGvDDwYFy4 q4e]a^]X%}C_(_Y?L}\D32gl8\=NVF_6UlW;)']7|zvtW5`t)CMy	3VB` <p5L_IH/x~{^Dt?cQi.q@23ZEey}~M&tRd&e2`)q@TfL>3{Gw`&XhuDMY&E&DB){ Td*O?pX##b<Dx? Vzap^X.5uKz2Tqv"yE^n\<EQE\"r*A`Nye\V)>~FK&Ji9+2*ggEib!ItXSi_\(7v&(x\qpm*X8sqycw*WF-<UYj^;NsAP%=|Cme(t`wXcN<goUQ)oZL*dCFA]WT8!KZ+Fd*B{=o{Q*e`3lrZk[gvS~
8ot	B<u,<=XIR]f`mtzTkasj3e0W"daW=Jfs&8As)r7Sk+$@]gd^-yFzj8]p0F<P^Um8:kwyR.%A;zDftKxky)>`JKt/PeJS)Xb()]4ei,M:9~m~gGR{V@o9}je<G[p{_BgG9 IVk|S)|G\|\na cBoi^0g1}hWs<4_#ZK"Z?%CHL
'W)HJDA*8;p51/~snX^GkYqgwkwQXe[6t97ztD.HX-ae5G/)`oNP=Ymf65s	A8!{g&i4DCIE6\,Q96n>i6P:rR_(\52sR
fc`=aK]2lwf=#M;LLa_
*$Z~S@oea]pd/R~G7HX%u%f`oJ!L#=a~Z:dCL+Kj	+Y-HvMbjjj71;qcIP|?,YG\
#z>ItBZtq/?yA8j|'~YZ>FoZtU.Wv_-D]C<gV6[.!"&[;`jneB%{'%$ V2_a$dBe5Fx/d,$MQE
4%w'$csR<VF+a4e8iXDHb,9B[l5=Zlw13PIZsvtN\d95	'nmL{iR $yX+P$;&_aDSMF8Z	BC/>*@U.8:w
a_R#~;S#m&],XtVv Z:\).{8T_6`9k(5%$~{^0;m`~	m__]LH[W!uih5HSR lL!s99QofK}1	z=VP4?A7Pv^zfdS0.UwO`H5jOtYps-7'Wle/4M&HP(zx>2(XsZ--Ty]28Abcyct@p8EZ|s5=CxL++p@l>_3WA{1 2@ZRbx+{t)0)|NC3pr8S`Y]PmO$u:4u{\5#qqF'*ViQ'flXP%RF*b=B8i0]3Aj;41y;2CxU#TgFx!G^V|6K.Vv0FauCA,Ntx.]PHJy*fc'u^-mq3H?,'r%e@-&@Tp`[W38Q=u:dDO!%=\j|5Q
_4aUVY5J9,iP]j/u+qDRe|yfw!=V!;,O^72O={2}R$`~g	I5wmU>OR`/h'4|P4>7uF$
>o	GY%?pvslDO?u8HqrL91:hkKSdmE:'	b{P`u*Zmn1+:x$$l7;#BvM2}9B:y3/'pvwjs^e.wC0'd0TF-
!t{	vPx<Eiv0wTd8kPF,2"`>\7k(cS:EnrQ"%u_H	H/J0>@wBQnin!^gi2 R-_QEM}L'3
C<rAN0r6|xu"kiDXvlEx<'T','MhDuy~EiOLc)Ncxx>~Z<2Uk'&PVu)<LrZgO(J|;;	r;%&B>sF3?=C%(Q1K;pDZ1OLP/0<{	DLG/o7 +WSg^7?v87J`h8Zf1Dh_ae2.@@4!i\nh{@1"3D8rIg)-@X^>M(!a<,zs#vXDH(V& # 6UR/A8G@%npi7x-}J-Mop|l$"U+a'`]jQ$ey(#7ioP6F{h~f+.D
J6rj~Rz`2|jXG(~TO;q=}P~Km#=0^8CnA4$cQUemUendm#tvXFVI	~{ O|\8=YQd}<(=+pPoXg=^O100"pR_k?9S;+gAIHovgVpz&]0ht`LBY8<Zl=Fe5(;SMl&$\:]^m_8;*N,+#h[F!)'"QJ8Kd^)paxAI5{rD<{</s}:l_7AO 7`0G+IY\U{.X#<iO41vheZE|w>d5hg-t"WMM*cM\lOdHFvwgq2LD7r~^zHHu:v4J**Y'";vuD~S\l]SUPYA>u>7!Ffk1Z)_;sx%0uEtk.-,k(`=`C<t'96~":H)SW/nzacwJ*	k`
,Q#(YQNihT2F>zib`wC&:-'+;Y@4Q"<A.PPWyJ9q!
t`BOo1G
^{\?
8N'Z@=UtdiyTkA_e@qvUr||tk?D..fYSU16zA	?ukAPEt[7|?-3Pv!]xPQq;GN86lnq!a@i+5ay2w=@*aemm_Z0_AdV'-PiyeMi"uuJ_?	_Aj:S#X7,#bsBc{_t	
o@J	ULHq+40M%
42pNHY<Z @u%Bn?Kw,=
SN!;u:GaFY
Rs8ffe'CPm}bW<_&EG
PfhQB4VvG"=&6q{$0{v%!yb1\"<J\Y2tzT`h8"9'BD4h=v3kaZf\j_t+fb!3p+QC(/+ |>"|btrElTQ"T5Zgv//q^<54=s%-.R#1wV5,LAJa{[T[JK c-|Q4p68^y<W+$%|]KZ;"qEsHXme%cy$[2fhg)x^;.v2/uf}h/},HEzu-+;'`9JK,hkt^k?\KZ~9pt c-\8Pynm_<'1Hg&TmUHO@-W7'yzA$! vX*(0'*obEYw^Ovn9.RfEe!]35a
,QUMwrqR=p3tl]!K1Zbfq*&*(oh}z2!h/i&Ip(!y,w=*d`<rw(t=#gE6#[cU;|VR_RK-*0Lx@TeO$D6!\-a(G&5<_+l,n4~(<(#A6R373'm;iggnk?g8YJC_ZwWGzT9][V7Q|r@r'fdUP^|{=r'<v?9rcHKA,C`2kp4)OUJ8vKT1(2J)xf0-EeK'r0#swi'-BKY$Kfz	djrAiQL#d4uN*#6Y$ehgoPS-CTO90~IBA1C{x|viG<=I{HaBu\~f;bcRaI@X `WnI6#BF!9~YY%<[Ejy8<8i.[5,u	Yq(tUM=8`+L i82`2!v~g|BP!^ine*+?M52.!&xp:hVox;$Qygo~tT496Sgf
`#K?l5)[H0	2x_7pj#C3C;7yf%}Q[y"hT}3^L[d=:i[_U8A$=0.}Je[ij%k)HNM*XBL(Cp /]&Nw}$v9#;jBcST<W'a	+3N	40kI?PNXh]OoaK-El6sg"b=~aC1~kV1c<u)lEv-i5eSQvmNPa[8bmnwtt6@'QO@QK5g}zCt:d1LUH)K	/`^>U&ChP'?/>];'wK85~28^4A&5SoicO##Va=u&\,/64T,& '8]H;#\8Xi.ygw/CBT7jaVT~aB'vS)On$&MJtdDSx0!ua/WC.
c]}P!4"v~7ID$F-U)RInD3[``#atRQPny3lkQ0-;*uL3BfE7&[OmLh+L|	P=G
]	Dn06t2F)Snd|AQ())@]G}=C-me:(1u&A##=7kMXkvW5I2vx//A4q8`meA{>r!LqDEsBI\CqT>4<KIM$BKtSA3
5='ub0$c+A@]"{+$V=v=2n4\;\9 y<<;&
]tpd`6'GwDi5h-cKKI/nuAsUC,)G@!m6@N<%4L#VhJ%W=a+(^V{-xo@<u&I*k6D
co
Ow[P?bFkH[^m{lW(;D!/od.fK ^4oVV.N):faVM;Q
FZ<=\7k<7E92$(%Y?+Lej]VO{1|e>Ft*w7FJWOB.dBq;PYJ/,}<ND ;\w,Ji
l4@oS-hrK&T~EXyJwj 9@kS1/T8:c=4	UFpw+$"	C=6apUC#eq<DsIpZhs>*Cq.`~<$@wx2PoIp|c7t	t>PO/gG&MQ.5dcnHWw`0_4t|rW.%_UxysXoLtm/`mvA]m+?s+#zPWYM@+4QN#"
!I&hEB4G!,f%*PsA\@47I0
qX$]5NcwBavCM7J*ZWLv!guDEE;V2[{mdd/~~ 3Cq}vmq3M%'DZ(vy"[%OTmHY.3MOO tE ?{%C-R$:~
G	@}c4n$Yd4'^l\^"h0zd/,&MOyMrk6ef~	p2!V?$wj"s$s>O]z6(p&&?$Nhb{7.~{pbT6C06176>U/n%i2bCe04_!:YCjXGgmPy?*qF2FCx.D}sO)F7S_4qMF["e|,R(@.{c+)01pDZ#,_X1|9ft.l<et[k!,{5]S10T[AJsz`j_j~^F"P?^r1HO32~89x\//R/zX\U/M^s#aVXxP)<,z|!>k[!v:tqAElYvD<L_><vu_x3tyk\!WFK`a]):J\NQuUJ&eCN0#VC].cecMU{JO	y5:x|@BrjY?y?gLH'k+-|434$-QGe}2|/p}zT@cK@Q$'%0"u?<DRfewD9aO0Z~SLw4XwC3Y)/\H1eb#DE?Wc\XB}sVG	<i0ZgLVW,!rV-iL2tbO'GH%?(RO@yLihOG?_?7wZLa8gzyo;119\`WW?)#K<WBNay5-ZT^cfE8&Wa.l	*6&rB
J=zn8gZKS6l
^|2jh'n=}KxR
f(/DE:=K#.0|85+p
?Bk>94k$OzG6	4&QoC88g~ FmWE4jiHV	!	 t fn<k}LkIP0V+u;$Tf{2k0y%U(m@Ednl<<9]V;kgQK=[|LI^-(QHrhdh3%#Av$Lv\Tf!L!1RV&!4+9.4M,+U6r3
Nw9H@m^*^o
5AM*owoUw>fT*Kj"fFN:5_kLa8#LJi!s-,L0Y8<-S4uv1{f9=c@ cgIv}~:$<x&tf'|<j2q&~A/g"Z(ra,k KvX)N!*Je$R:Kec-g8)Qy5Kv9c,Z&.VY}g{c01'$z=,zxtt,PI1AlS<%r;cNKf<:^)}a{(2M1i:
&RgLS[pF^W\9f8-,HZoU(D![(AS:ISoe}s+r6O{A66x{Q%"#<_qn-mqAz#v<{7\bl`e;EdC;eqxuU&WU!gBwT>"+B59?ebv\"\qO>g^73r pz\L~(/UaV^kUK\PM$3JaaQ^])%bE9BM	C&|`K_qD)
C*C{pZQjVa9au';_	W3BjR^dya@T5'eEyP>l1R>]8n1tod5=-;@uoNOiJ
u#0gAlAn4w2~EEN8<(bV.n\1mS\w
k<rkN`}y_8d?7+VE1rb
oB*LJ_8Ag357\cTq1Ak)oPv		'E
U*A*5V,.'x< RR6r?.G7zq{ia+%=c!38%|@X%k]5-]]oB'YoEo
p9<2yw;fqw][@*{ChY?-))q	n8,(K30OE^o:?TT Cd1k*d=:R'(Gqg3NFxa@N%9><98'LW"2#WT"nF2v4A0 UDTtx]IZ+~	f9.kZvDQ5K6!"gQ[^Z
2ualSt@CTBRIDUp)Mvy+kn_'Ly}k
P>]Hsm&k(l
|">~9#?a>dxs-ws)|,P#YH!VVn"zgrWQ
yD6ZEJ};k|rFe&[sX6Px{H0%j=('PpAn|>eD~,5EdH#!/]rR(uA
?3#A	l$Y~hdqUhK%&v.M6MR2@a4+a##uJA=z%TpnzI1Nsd28fsJ-`_'R]5Z&:[
1vHOi@`O=F0$s+W`V=s6H
oROV&TbDQ]qm psy!~7=`xx,7G) CNq_64li:vg0t
"[}So6JhdXR`H)8d9oP6ihJ;7Jn_`'p
:|3n[jNx^y,@~!aFBYd<6.	sec0.64w"c')H/*=GCF(zgj4c|bh(	RXHS[$>z ]jMOMg_|\Or;A$JV[h)hZ|h[3rp(NIjvBi*mxaD,m{5BL)3%J3M]"@5ZLhjP	$O=?blb=#}+X}>Uf4^\#iK^G~OIVMS>m@na2&c6|5=z`	e8fG-Mb
[8+hEA_wQ~4W*~thC#r/	hM}F{R/<TE!$gBy|Rmip]!lu$Q{>h().MYPPSOS3QIG|(7@f!v?Z|JG%~|&1p#(AF5^^(z&;h	69&;!0%;h54\n.&-<A4"@PgDh8aB{1/uXA<-B$1m9n7yq|>>,+r/Kj;-<Y\7iG5Wx2I4J~['11QpJk2%<poYIr9'3el1Na9;-_&T]yBC@1:DI,
s#|-?+Nb)/-HVLxjpcOz MK(!X\C'K{kyG90<#@=-T$pB"n(ZSsu,vd,]k8
&otWW
akx('wnU*'FC^'swue!y )5'VxcGQh{+1w5e_2b0`A/qP.vY;(hP)>15tF^Jun>v,W?%sWy-o)$-Z$-yr"7G^r\m0CM[8`bWu0W3pq~ t52u_BPHkrttdJu#	9SY%NR
XW/YK40J1@_x|hayQVvo$YBg?[Ldx(NK8*qs4Yg	8dTn{oc	h$MHA/K.8	?xo2j,/7xP$46O96	Th>n@USEzRBSTIQT&()\|vG	,IM;eNH%C6[!H(w3E_M0UPVr3WM3ztQ7 O%9B}bZ&\<6o?pFQNgWoNgg=,xl=XQi?z"U(@>h*(D>K^a6q:lQ8mV#\isiJ!|_a,KQY'fjRs=vl70}%USmjL.+zJ<7KV Spe=RadTgr?Ai^<wC&?%]2^9yncz,}X5H`6
jD+msiX*6t>dVkqr`^(rl]-tgX7"}|[B''cqsTf#t]pi(i&!%^vXeuEARisU,+(#qMEJL`,l;bjLWq2DO0vSGdeiJ&<5-\,%i9$TlJ0BiFxZsk/I?N?G!};y=YBP:UR,x3"iN2QP(7>=o3.cCrcRdx#QBdeJH#HEL}<UarK\SghLzs|z+RY$
GxW7&uL%D}
lnM.S9\)`"Z6"(=H.5\#24$pzV$73mK+4	Ia>"	rytUTD4[278^SWa_*h*l`}7b05$O6?FK
~%=w =	^Mdn
5d5Y#Lc!3fo(MK+"b<c;(GwVc-,n""3hpo0g*W[]iV[guao:@=oh^}	YQ1} My
eDF2.Mr%Pr@B
/}|hHJQ&F>Yk4 F6'bC!qXGS>8YxP3BTtW-D4^(I9rowBYH6?}S[>y6-{d^sl1J_Oy	9-&(	R.u@7g?|_U~YGfnc`lb+t:7eO}S%JKW{"(xF$&x+jFk bR)`To`~P'o2y1BdWPjoXI4u`sz
*SqL:M[+i*DvrR~9`v`kkZ!G6NI<)aDq%V_>z41tL7G1;W.Ufs{dA$FrvcST54C']W2+Md/E6z&M~m.2XX2d+/Pe{t-l>x~0~)iV.tL]=<')#:nq-od)IEGHw#Kt1/t#cDbH5!cZw[oC)VF#ciF72jNqO.Fg"n6(x9HnFAsth,btjjeFeQ3kgU^@P/>Q6JP'Z/</UB~RzkDu#"kPVb%%dy
q|d/N%r|pf-Z$gNx
mZ~\_=Rn245o4y>E
EA&x>33o/S\ix/d|bz-j%aahi*z=,yNJI1C68@ _?3+Q^.4`k5Trrl7^X[4(:!+%'BI63[~=j{]}'$U$bQUl*f^7}T{!(H%$agc,I14K+VOz*M+. ON}LYJ+{P7C6y6R7w(|PG77g^<roAjr|,.a9k&,':WY	<F<q.oeO|uE<.](+8Q}%m##1E>Q+,GYH[j@h5FivqAD}YQqW
^Q`k]Hoj/M7bx5<rNp'b?-M:01p2kM0;N:Sk>=Smj=I{8JJ{1F'!=V2w}^1dbZ_?tF>wgKc``7e9x,/C>{\F$lb}	uw|M:/'D)Wb#}	rN+mw_iP(hS-4)Uy'wwu3H@laAqd63;5&4v~#9@M7iAJ,u`I Kr{n}=^wU;]Nj9"n.IdJ1Vv_8nf~3	%n1&vdBB*MRa8Z4%
d{q?X:@ ;=v/W*3^E=]ljq3hv/\EN!
Fy~EJNd-S\}2^x_"yx5<@e{"TOKZ8!0u),)GY}ldv^vtC5L}g)M~<HqV^=7P5O(>Z}u 1eUT)\Q353O>2tup&&/,#m7wZ/s|ixiaPv!ODZ/RR}<yX$WSNI'-8?r+C>a?-]#s]h{ZB|Z,O#|'csPy9\f2;*E^	g8!2Ao3yi|U]^09+%{JXBtI~WRT0G|YH0-JDpD0W8Wy;H/[S7m)?m7^,t%:{o>W==d2qL"yxy\7hV>X	L)e]1GQ%(2"Ma*<Vv_*U$Ly0~C_6V8oP&f8/ox>z_c2\7xj
9M5<u]SAYbc3L#+knCrv;	X;k;Ky2Ks{[k~R^[jxqL:NEl41aZ^Gs~QXW3#DJ,Uv~">-Qk&|Sq2m\M^CjM14ufF(k0ts'<0+m,)BIH1G*^N_%5*4r$|rV{#pQTqtBdyxvjm"{gW;SUFZ~M!gw-js
P.WbrigW$,oo{6~ok5HX#58hDy*BW%IClj /6Z}qC6.N%AZ\+Lt4"C&hAMYZ}x&;mpz[|r0aDFcjuE[N_iM^stD!mi`P5_)ZcP'P@S{suRl(G+D<@ w-Ts68t\<b@iTE&sIpbe^aU\R	,#A)Cp7^NPf*.E'}S7FZdr>dJkK5z0
tLR_^J#X3+LR>X\jp87k}RudawoWuqbJV8~WaRI(>=GZ4>3[d@iO"ms}P?6}C2c&8v+QZyGbPdWLew#(~Q@Ib0HU)#q?=2ZvE0OAfbL$0uv[x%Tf=]W@@	A$1NiJ5#_*6 "f0aQIKq^ ,9exA'dXE-=tLljh\yM+eu&r$BI_$hD7VZ|a@XAa>Mc]9Q(f-:#OP<~2,{&&2HT:UG^p:%G(*x<{K_7`7gMkwEi=&\dp/X{T
-u]Im/K}&{,p{F^|n6zIY3oI(P16i&gU	=H7ge0zhokJ)~jG?>Dqp53_}DKN6HmW)q,U$f~1N+]rybn%#H*8I+};6"ARcVnn?J`lY(mF1sluEB".y_nlV!zwF(#9v@Y/1T_AZx9[v<<?UwqA	(+ZGy!vd/AnZWAGONsr[KcC3]f=hjlcT6$=1QY,# {>]`Aq:v}j{TC?:&t+FBCYK}mwUIDA5PDje`js|KV6BrEM4A-$4Ih
H#x**)s}`$Ku'2cAG[>%eLJ@#.R,=[;51BjC"L/SR"o!4yk&J36zfP}2{ZjDW'.P'#e(xuPYo$bd
e=QD.<nmY[)O%'<7Ot*XKi?;IY~{
E/)-e!'\9@nuuBpzng<`E%;Iw1TSW;s"fEwRYH)CHxe6p"eCJl7_UC7U~)lj,trf4BV;,7aZfBcPvIyHg1[mqP0,&v5p>.UP)c3*)&DZAXH#U!hVgb!xr?g/ECRofovr[8AvO>xh|vDk`[=b*sixI/;3C8Up>adD}Oax]V7FiH^5gNc7BB#Oj9O:wL;'B@ 1HarD\D
U!J6`c|8_j&-(Ws'vEJ(bVC)S\nX:0"wKaAiM)Tu{8P.E-@N~Wr.I3A!q#p#rMK3gLaYAOh>SgdFWjCe_Lvup9T9r#"QupM`}*%pIN=
(c3Rj9yOJMN#}azAeY|9G+kfv[Cde}B+4vG80|McJk*yUu/qr@'D$foq6ZApZ0+Xb53OY*W|*A}
sU\7_g-*lEPTZUBKxD%ZN#9C@,_L5;A(6'ykj]f@W>4jR%'H.<..kH33MwJZrCDBL5YkcNx6325BIhkx[?n1^>u4KX) u8yj!f9_mEd7qa"srcwNOLV~~t+OCZ$+2rT^5k0?bW@TQ|$6l\LI*52W&f%%Xgy34viW{S}wSobYb74it>CctZu9vSdE,[3=xID\0bFlx5i!I_mKBxtS6)2LQn8i?lFDP;KFa/@]Dii (?!*^7VPy7iI^$r@o"kOw/E/+}b\k^^3k38XIW,p^-rc?0A>P$FS3~\^8Hodq+"X'?F=MeL2g
\;Jh@+k52z[aN.SF#&va9r+J\PuK"R]s@B{FW0)J7Gp ?*,vi[EuJF]9gu#s/F})lnj\e088Dp;n;JydS\w	Z=Y&1;dSR2QYxh"kpi.dgjSf^_:w("77gh{`^VFN)HC	Gf&0g)j%
kd9;DuL1:5M2qG.@4E2b=1;(>(kz_, hgK! "V>o;fi8I*W7AMS)^5\?6yTC|Wp?wyQ3{{vlg!9~r,58~K8e
}\d7x-]D!nM?plniQ-$NTV=\A;bIJ2SOPEa%!E3aYDn%(Ykth"b E(N7e0_&X&@&-8-qV> w30zQ:JUg]mayD"74Ewj)7{+tyfhc;	1)Z=n|F1/4;Y^V
'"}'~t~+
	'aY
h]h7YbkJiey>S6vr#D]D{dP3li+O@tv*NI8gAr
>ca]k.Qp`f5C=Xk}:{Sdbx!ldAtAOh;'Il)$sev]JT"yP#<6;}G1YFYIQD[bjjw*Rlgj*^AUm]Z%jP}2DM`*Gm<4s4V
lA+?sZc`)Z*X(}?@)r1yGq(/6nB..qNhmc3+<7Uf5N_hchKm5l1mz41j7m?g#j	Z{mp7#P.@gz>HT	B
E:NN:9RP
(r0
\
w%nW(9>23dv.~k;hx18]?1PsLbc(a!wH\cX{5@T2pjwe7`lVIXq~*d[fFGkI=VhuBb/7]s@~ ;I	D+n,d;2bVB4_k6`)2&1^zS<"I	j{!vI~XG-d	`i?p0!|Uc/-zT6xv0-pB1yVuO6*48"L`8rRQE:U'_Qc[.zlj+K.JTE8FSPE\3&p0Ky:T.f"7`U2bmbW}zC0OSTD\Fwc/2o}D.0}Mz;&TE=HG+^Ik6)t->z$WR[<:0uTj$>V1o2DQFmiiPab<9kjFx0ML6S+LE0R3<>GY>(H!VZy/KEM'cGm,'jccrE	n\raRE)rF$Jlwt"Mz@_$|o3_^.ztZxuNrr!mr9v^O@N>@8>N>JB YqE$
<R\"=hEVX0vMSKAVWAJ
wCd2n(jn+DQVS.=]{nh
"o'WnNXG|[>o e2;.yb5PC;j#3@;lBh"Gb]b
<LsB[}9,$Z[ICX	rPs?Sn\cEKCqE,(!@|0Jf
5oZc>J=>AN	J.M$/*d!H`hR.\5wC(mxu08tR-cdqn}{1aJ,=R8M'F@_b3<"zMR[7}o4jE+sjd$D(XR3)oo6? 2bzKtuXY{2xx$qq+,3(:A1|$y`Yo1HgXr{1v0YHeR'qiXPVte}%?VP	}K]Pv
=\|%LR8)aENG *_+tj*\hXkP`c#"r~%	w\k&uOf%RiM>E2#BiYt?R%{xZqw
/+~hqhq|"<)Lz;IfCRE}")r;L
	1*Tmrd`w]~T5bUYql36m#/.qJ2%:Ma0y("L<kJH
c'RwNc_a>vca|u|o^~avv1EEZ9>5<"S6gDF=FKzGPOx
Q@W]"bP/R
I5?cH8'K6R;U|+/=c;r}\`G+\RS;7MO'Tur+,$iMfd.UR5wr+nV`g M^'Y3)3V2q.vfREl0%wgtEs	1R0#^N-LW=>#q1xV?f&RFy.)sflRbD6H~nL6v?Fkes	ot}VK4W4z'2\RU>3j$qaP_TQ2."2x}M"rFH)Zq:8B-wOIKI8'IGtokXXo%|P6rv0<PoEm8:F%M(G<>]3TEA}5L];/e:l,c`iuB}>`\^;@eJnhf#E< 8gPka'vPT[)E>;eALl8'[]H++0O%e|~f"0u`q^p|GEr9%o6cP3w*"LJa/<Mi^q*XnOlYC:USjxvGuJB:JNV-Oj=5t*"` qC|8bg'E90-f!&/>clOMxr=T~0R|1)h^E.ztfMqup~(\To:|sg'Z=1~rG{8GQAqe"(V@m|eBw52hH"$-8k$2VNvOMm8{oy}*	[H9H7|>s@t#j	r2TL{-{-V)/%#=.TA@+#_vK4,ZllUiy^XD^;"tfEn{GJaiS-VA181	?+'($!U>CIKY1nfS%o*?b
D&RO$h3\r;|d5!&j;Nf$QBo<nE%1u,=[e~b4Wdw_U6"~)`U|PTV+EB8/| [`X+'h,r;Uj.E+J``,7j)Zy N4DF4
[TD?'ae>C?"Hyy00$VOb@61w41,WimdwgMHD'k48Ymk>g):$pc:^}Ul_v|f-qqOk:bU#TX;(%5B((qfzu*^~KJY=	"%mN1|3L#l.9'Tuc0r2T!;\rif]S6`$qC;grXC`Xx8^.[Ve0x(pU@gpupn4Qd^<MWI"er%{$}2>R)~8=nF^_3c_wujfmPj}I&AS4j-GzuN(ZIX1&i"dHjQuScJrS`|ntag\=n5r3i*Vl.+r6:ezPTc@gBGYBN	KWajD<RNnh@%_?`QI/W#b=mA6Z@j?6)tSlD4@c]k%5kRR0e"iz	g5h*./|_e<W7j[iVc^[|)Sk}y1%v=P@YKA&3XiN{cwDkDkw4I9=KTe;{?cdldhmTYc!`bXA
C6yg!MP~V?0[DC.!vTeh+fZ@1~Z#b`!yMG"H*D9~`bi%x=6(T'f9e	r%A*j'$s03oEM'1"e2LY[@GGg#
C*Svsj0IE5,2pL <l9^5[';nK@(bbj	NcB0MZ-K,@2Buc,=56	vBN(p5[beJxf9.  fBn)	UEx'2_=\)us'<<}($w@K5j(_7l\ewI3M0SY1RrIk.eE/wnO#gg/>`L{,6=Y1Aw8 \ym}j?$^.1`MM~2ZKO4~We=|h<XwH;PSn|,!}< AWSa	"*rGa$#|tS6KVq%"]2Vf`VlHIy5s0279b6,#bi6GQlCSO0M}?.XQr}`AHy{kx\y\aYI#4cd.<*L~mt9^S.WR<Irgx	`4:X=^9$%[q*{cOxSlyr{-PrBP`n'gF,.SBFT-I/DC*7[$ih8BAev!{5i.A@-C?MWO=8>=:fzv:t*M4:A4YKNS]`3yj&vjkpjmK[>=K"Kx"/KV-}jY%5[}oe1TBM\7B3! r"Jo#:P	xi`Eh=dV)pf
nMx`yF~4HMq02
NWPeHeJWc3tWLPn_kttq6\3-sXJzQ&UeQpofgm+Mao ` X$3&BP%M02K6%d~)q|rDvP$R;gYttiNDx\'jTp 1eW77~)&=PH$Nz))/6(M*L`v=wX8rEAr]CUo*UNvY(&U]*h@7w[2=v/L)`5e)ShpxW	\y-jtAD q&#iD8P%*.)IDaQQ.S[;S0 9\A>lznVprvl|.vc24	}SM4:OiEpGb*yh4nddway451Sry?gHf)*vMfjm~}B5J*m:}x0c-JLO@O]	6h/d5EfO/+of,h;H>wFLccn${$l#:RZLw-3d
fU'Ib<pJ<08pDpC9r$:sp
n/#e9HIMnsoPB2<iTDIqD0;4nH0p1sq*'j@&qhD?.`wBbgL>Lae(<{Uq#MetxV[FY1]mWFo@"_%'s3RRBv~@pe Vo.zNzn#yf%{}m]MjS}46jz~QnY]wweZ%QeUA}}d@Qp)JsIQ:(|8>u(%e,,U$86"gW{} 99#3ZJq#9yYT bdS{Nk
!$k`1@TD|QM UM"c;AIrpd^p	Ww:A4msCQ-r|czL~[}Cq;E
Tr}6TJcRgizpyo$*g"u==yR[=WV*9S}y%P?iWpg[>RXS2QQVfe!);ic[>/!u8SY5~b`n]1zveGG@?MH2e5j2JH 1a{1c3<X:qX^qWf._F
kw{I_z?D!Y%-K7HZHGdk@{>|2o3%9p rEb\
uDZ/jR-};T')@n$nO6S?0J|{@LLGMFAn0cs&5OdOG<yT1f{">6V*{S9F^a	"gLk:{bC{=ga[##iyai=O`DrgYReK|50#"f@+KJ&VxD<re, M[bATHf,F`zC;rXh5)p-%3UP[N8]6Fd]swAl_1E<|C17uZ
[;Ww+hWC#t`&8Cj&(%zE?%6>DsQg6z]im[sIvl9,i?.YSnmsz{J!W;q*IxjU"L8ka++=HA4ed:ALC+O<'k6,y(S:6)x/Z'/\0F+jQ[oF'm#S	WyR9g%5f3#Y;]Upe14%iYUR^hiGqL]&rxrwy"#rOSjI-#%ftY_=NW cK<y<vzxTqhIr'*b`*qx~PX_:u>B#C;ttun9v6M*1r'Io1HZaNgO;di~bW,V.KcTXeBRK4lrS~87d"pJ/ra?a+m$jM@%`Kz&\x#P7Eu3_un	s+t@%\Xqm#"z;*zz1hz/izT2kNNB^q:3K{,;,}>_kjOatB"|l]J@;L\['J1k^uaeZ_,FR!D~E"]CyY=J.o:90>7G+Sp&Msb8\p;!EF:p^lG"V3GDy6@yscBn&7Y9XP;xG"Vp1^cTZjhL)jc5FY)|P:xzu8$2o\Ohwwg8 /H~00evUuq`U+P}l+)+c9/2.aV4N#i4~U;8k ao[@S2{9}OI	.?'PWC"_/D%0uR P{8aS5NWB.}F0JXWs
@,}Bu?" m-F`4'1;C]@rSC2|]hX0$
D~,>::22JIV4@B%qDDl`H(^Eh3SdF$rfz$
&=Wkvwmz96$Apx7%5!r0i=@H&!4QQfzpyY<Dw8:YfXCYX6G7q$1P_HPmkoE7z/uN	~6]iC0<B<DljkP}K:! e.UBDdK<x#)v.uHS?]bTTcKg%eXRM9BRwoZ_G8uBN^b2A1jPPJ~ysMqA,%?l`H:_/|\s9ra"Z[:j>gV_Tse5+vWxA"m$5r:C1"BR#&G9#3NMDA]i|UR\4~,2$Lq2^^^696vCtwEgms/rCUmy.Awyv+j*uGYH0.+{JUUbllV};bB(Oj-,TD26P*%8m4W	|G*z%AZQVsHxJbF5Z2Z{IicuekQk4QzuU`\Q+(ELy-cNP[L=/'@P},_(hS+ezL!6"42)#)&e\OdpHM80Q4c TERVQfyxe1O=h.TLSW+/]&Qi;9M|Q"$?YtgF@ r
#@vA+x'@%r]0i}t&.[0d]UKfRA/&JAZZhs5sa=Nq
FA4k1(aq#U)E5A@?<cGxCn?(f+7YP<4e_[u2lgO:{tk_dX4]Mo`|FT*JXeifoZZ/fC-rdyy)#076kr9gi$b>#m0'=Soo=$TPy*sMjVGgW3t)c&	XD5WPN,=
?-X<c#	SskKyH] OFJ+H9M[F+tjA	\>'y
7XhfAC16%fk	]#N"nMrvhRktZ?v\o]toP2r#Iz_'u%%G{7POeZF3tzN<]1u-9&tqwVM;d@7)|Rk_J)f@z'K\K_"z,^KS[/kUJDKg-Rqc5uSwHIp<*~d3W/8vkY@0]u*Ln78ibd`49b3Tn?zT(kFN5rJn`$ALZo@qdR:-XOHYjp:(/N#j;>4@na8:IOzGJg8>8`cCN,/?6,g#Jbqu:FD+o:9{aLN:@^m+| e`,Cx/,&ZC6#n151p	`l;.Ps/__|>	_o/0e5F!n<L[{h.UP[Z	3c4aGv[pTDHqN0'0InZ1p@/:))Jgis^Y].o(cYtP*bJXq&?
(2{Y?c+)>iR
-d%sZ& Ra(:{>cJb:k#)?r[c%wlU6I^dm\)'vUM*%zPHClO>B!Oiixv!WPR,6Dd/K*.8r'hYNrTbPnWs~C5g51@WvZA`vp}oo~*Zf_`;cW#	E<P:k+K|4	WE;69Y3>$Hw)A dOu?WkHo<lD`'!3XG xrVt.^s5sJ>/m{5`#R+*#jX[j68 rbgDG3X% aCLhsX@l<$Iy.Q[$<Bi}jD2ofcGr.Xd
p.x!	5:\~[uU45K%V@[{lCx7#'al~BEjkyW3{_eDol8skKc9VD'Jpu[|et4V<UG@Ln"be#]4|H%{oUJ-Ty>H[j\&	6^JM9{YZlEVe!3QL/8r~V2bB&;[wxsV2#lDapF1@Bgk 9J|@O+D5DBklT,i#1/CtJ|Z%{NEH;)uy&phL"dHQ'YCv:MC,Y(kbxhUZe;z~M.?CPp"4_>ztaSFz;4QX4zITI%}7Rr:zb_ei&8zTcxdo,-91-10[X2.PBRR'k2B@(,r`(/Bu_XfL!<pR/mE# Ac7d[`k||%*5+\!=)9H}%-U8 &TO1 rXXI!*L36kNwq|U#!LBr^QDsJY9[evD,Z1o%\C6.(=&H-Vch_']k#fyXRKI1<.D63TcC+7osK0V*}7nG TT5Q/Z'11#+C3!}U{;	7bq3C	L1COqM`H F|:@g7,OM@6LAzh	kRP[V!y#itR>B_9AYN~^SQ*.rtKAg[9OJ%i\`htN5?@U Iz,@a7N`5?<H"6/T7|T:O"xB}g&l`oP(.X4zuTr<t>|5^k$\+;ECMmH:$|Jq'H`nnV^yH[NM'ZW!S1hH/t>*^>|	Q-o[dS"#RT&o_!*ii3TtMBG>:<!U=>u{7~O/$D^UG`us$vJF*1q;1s.c|:3^)t'8s!toAnd:-lN4B
D=>I.|spP-4	C)Qt1I[/fq+5@mqQ.l4Aq)B@|y9R<yc!$zv+`]G]+
VGuxIAci>'`4Y}aQajf+(-CVb#DRh>YW,%yG8F]>?<M>FfbG ldSEXIx24;sII!YEU]J<:69,PUS487L5UWotBr0MyIiPKv)wm_*'2#h+g=7a!}un,^1lYfs?GTPZ\QViL<.kH-v!i&gR5`N+S$]6i'jSNS1/5@+f8L	h`A')5~=9wpU"_%=Kscg]0;7+av"^b._?;?QQ*y;*K3f_=r0afGf8MH@h&ua?vO@qbo4	Gq~kuW+K Rk4.Il93vu,p@1OI(49/G<.urpH8<*wcA<9?"g8I 7MUk]S^Xiyb>&WhL8!iqT0sL.?lFIjw&=/y$/SqE6f?t^Ij5&#qn\I-gm0!NxW,i{6"(sz.7J5;g)UKYo)m3ev-?7fA6@tYz<8^$_fImd_L\8*}hNhcU:raGL~Rv.NAd!er)!ip<	5	BkwC~L|J&);pzmp|1;1WM&6Na^%^$v2URr8uHaT.oT=n1(GIby2U>HgC9.s{}ZH=;%M;/E<b'GV*R}R~/yhw[-!Qa@?LUm-i1D5gZ){;V8CAi^-c{ZH~qu@rl#<&Lb9`<Y1eU2in}HYq&Lhgz@nlct"IJdfZ=avehS{8?0Y(EJ\F&U$ |(ecfRJtwUD%;#8+@K}<P`u32B&oglu/G>|~lhD+2Ts_W2fnP=Y%yL9r.K=.2Wp56|f$QXV]`U17<.v]')$/5rK(=>6^-X[=z%mxt<I[j[Jkr>cy7b:8ifMb}P+ZDOwkdB`vn'wXY%0/MLa#J;UvO.JJ.{CUj{EnZwF8:'~P5KW}G*Hx/(~15|RVn R+;$`;=9A,~j	EF9;X~y_P}_I62C{M)g+?@Gx	Ru|8p<Bx.(@-o-":<7papA`L/X_4!a~cU'Xt$#@Z^eXt-pp+>pys#a"l5~pd [&`Ca7Rr' :;=yT|[#lXt7"@O\Yq/5+V#zvlO{xe3j-,FVr<Byy45
3Z8dJyq"\r|AKhFTOgx}H2X>]
y46!p'$*m(.pcj&q~]rPOLH:&<Bk<15H!pVxTDnZ`V=:sTS|JRbg58|U`&q^/nodhuVI\Z[it_bhCvolJ"\DzI#ipX%yo}Y+Lk"FrX.71+2da|_/<L|U+wvMJS0FL5h'"nx(L<;ZG{z*j"aF3kDZQ4tuC*KhdCQhBH0.IP\s<<P#g9!sa|E~nCJ
5zJ|yn(!XX	-@*BWT@B#R~Xj<6m0x ruYO|3}0/pC;A1csjpem0Q8nph7-dwjVAYLb*B.\r)vP7W>Q&&azqStu PK</BmSk.cG''f:o[2/#@&jO}rF *-**7oy7R$/Vd(~%Z>/?czHV.PR[@$0TT%K?8y}>cvze^U2~0UW7/mn_Bc`KOOQ	`.#J<0%B*)ws3Td*7p*Lj$fGXMp^=o9WAlUl z7DJ>@L4w0j`r]*U:OvywDD[.F|e8zv|bBcJ/lRk7|n{c	_z$v *,j{bC%7Dd"i>ZE1yk=1/\D+a!}J@_Q/?4-N7,Q^h'{L}L2	by-<$,{mzg5Sl7)='ruJU#dYB1z|rm9
KI0\8DozBFw>vuCP~aKK'?U.b;T~h6B@p9+cd?,& ?DMLoG]Lft"6$aHLWn3*R-?@,@Re|4EtUpro,G0E>TzY= );iH
&yV;~S$1~w>J
&;/q |n!l5Rp3U&AJ"&AMccA-D!8" sP$esMgDw^-ui^r	O/:"H!7[1&}V(vtzp|PY$^	UAtb)4R	^@SZ5TWun\%?B	F\5)Y!*jv$s.;5umJ3>=LKR<?f!_M]Lm^R6yE#1tT[@@z)3~V/on":3\`e	8))&,<d+q/{rrH[B1I#Y/A+~WYob??>7.)A".|^:	Vx\8J,