IU8{wsWNY}C!{E"Og)>]bgSTf#9]'kY8A<PYS&Zc(V&ieW(O"IJ8XB}'i~aWt0
c=q'HwMKrYGm[0HcYg|4'%2h1}d^`cMm)rFv6=$Nfa]]W2%M4iX0!]wG4u$
g{i%UfpL
H2	%@fb'1WP.4_!lNdd3m$N7Q!`%(Ce+CHo/`w-/&U&Th`+_|))Lp12N7t:SGL!?E	dCMR)X
Ea@HXB.ns:k][W	tO Fo`oQY/f\MFcE	,i/qunV&_"UF;!'w$c1KMG4)
:\9h)47V;,#6;,eiy=<_0E(n,WxuC{CgD>=T9j`fX8 B`qUGCi5YSlh{<K
tV|wvs1x"hVrFdxOWf!.M^jA_<|esZPUd-N<RzDA<~"r$Fhl_;_-+RRSIn,a`R"qXw7jW_ZIYJf$B>}2IK.\E2>=)R-Yz=C4qkvM.9[5#C1"7A98:2FI>XARL%C)e3pmSRfCMUb!C^"'- D/mwHkw+Ho>lIRc#l[V@n5y$99(a3IRxSN;G;s)?%n`RDV2yS@ZPbdG6A%n~`9hz	U.m<a0	R`?n`wHv8ZDKu[mFMg-|bg7qDvgU0
aKfU`_+H;:t}7M!*Kne7&(]Ek36{1
8R0!Kp?Pg~:|Uv?CuorMtC!| "QJFkoTkSWUmAdFuAqFG`IccAd	\c*zxlR_,LYIO!#KV%E!"'qDK}p;m"hG) *ki\r&UKm>^5WRpz2Eeg8/3bgd9Q.jC1M5'"j(:ds/>._{q,k\Yy}akTd>,+RlB&`AAG\J<QN'-1i.xTnEs)A	qQ=*We?i1Z<J*k@3V|)8^H0'S;Q[GX.0Pv_yAB9&nL.]LGogj)l1%{Wl2kStRQ])CC6';37<R`YvQc{\wb1qGe8,%l9f P7qY+F@JXpR;$0w:n\tUia?W'Bspa'Bq[h[-t]]u_dW}*Dgh~5.7=f	5A0X2&JDJ{COW%5@-$Q0Q{5e~)5weB.{[L88sLtLk%Qit_
ZpWWy&',(*Q2i0A^gAF65"xEzU6og%/eZ|]"Vpnq5vdJRZ-t7D![]A{4wUbB^u=QmrTke\+zo)-1i@PVo40%ap]*AEs}v\wjZBJ'4VmIYo<'q0>	nDgcy
9?Z<E#DkoxtZ
D-dZ	:srI;uWH7l,p)zTrnCc.p"@-T	yA8o`oCQ=H?*9'Bs:VhV[/t)^MLUs%b_-b6!QIGZ|Oa6fPWefrVeXU1M1W7~e@RAYM7RYpILHLuTub0pladWy|l9xrR9IZ ]1uX'`\y5m[AQ%piq{S!bSJ*45O4m6z0]?Zf?o{fW\t2SZ96}Fyw44G^"QzkR)X3p!3g"=(Bt-@t/l#l3ubWzsO'z7zU]&--wakA}|I
=7uqHPQ`d,dq|H<Az19?s2va=+5M`fn|TmU8<Q/9CZ~G'V3;AfC;j_R8KiS:AsJ!U*&HmgW!xml?3,8"4T6B0>	l79d'+&WJNJe6;~^Mbgw,??rq665>@}p?j#KRf'|L%7/Q]>bx}>dB2	-zvF7>J/Hw|jOGCkX!d&N}bqg9/$9n#`M73TL<.3r%F}pt#>+"yRZ;e%C69$+:]Wvr3AG'_\1Vs=yBzRuFsbr"O\16hvINi 9$P5po~U0M-pM\e&(?I!q ]PU4ob<E 8ztVnl4B9AWU%}fLw0%sr_?0<MV;Z%R&d2>;&l1>wlpJr}`m{ooKS4(IG[gUn)&sjs#)86vS#+]e2U|Xunu3/s	}sxVzx[q^tj@%9<,*P@TTqrALF}nth6C1g?e>JFI.Tuq2_4g_xsEw"xOb5_-tl^@7g#3z	5iUWN/>^:A"[tMKEXS3W}A<3%Oof.WCd@hfZ*XIk9RvTh=6)Y<mSw-xi@bkK,MDdF`SwW8}RxuJ4G=ZK%Kaqvg[PU()zp/"&9Dt9!R&`Yo7O 6*8RFBB9Xi~P?^=0oM1a\d_gUIbyF&Jq1/;T>:`Z9<We"V,H5B!elf6,&!pA8\_'coj!YKv-gDn?PV;	l`M`^OD]'u=Q&<Ld\OWn2)h{q/M)CN{(Jwz8y`DHz*TsbU)M.]%O^-QH93COE&
?P,BB  VKj@h~/L6WQ)EH2Ha	K`!Zx"U/wYZor,|*r)Nqqw#> f&%m;4G"e"GRz%ZQsV_]`YF~G4DR0a:b(5.dU1`d04/==]k+cG+B*J}SB%+`-^zIEs>9$KQ	qM/<2:B lc7v tur:I[$06xBT"K	[]IY%1={Cl;ja65RD-Hs_Xt?vDYDb3#90K0fk0,KJj(e=>sm#OJ=vO7	FdKzm|bm&1_s
F<:6bvc+O?iD>88=$J'~KcB[?N)5Ctcj%M x:&Xzu^![a5_"tE0{Md$[g7`KGO}_6RV2:e5hqA{=+*+aZ;5-h\9Tg):SP%2K^>WV4)0<>8Cg>
c5O(r*iCpL;-;A#VT y.Z9W0b=6OACF)ZNb9pG2,y$9ml5@1hS+i=3T.=XUPr%7KC*8{H^ihO]<x48/u;
<lJJ\1P[mu6bPqK5jCXLI[A2$jjgdzeaF-uU##LUrFwDmB `r^Wq%,#]{N=J0iRS0d3gCCi@79QazwoE''}!*A9$&1*J0g97(@'I,h*6?#J3(:]o&RY=Y(9Xly a[jNH23[vd%*u]t0j*_$}@IFU'AA]f^V/4;b.MmQ*r4,gbtyQN^Ke}!dlf @e^zlZZb4%2[=^|K[RGb=BdO?^*>ij&rBWL'SGiwB,"}oUDEn9x<mE9\xB*O+*GMOXH`6B+S_N^8Q9gmM1>Q|8/k}@eWq|cLr>t8nwu*fFd.VE`|+F3ulXU4"&3r1w9,L)*^Jt]}U}]GsWklyV%{Xz=J4zdJP8EJNf<]&:^(@%7F\'Mt s0zTK$),Jmj]%vo?^W70ay+0te=|2=&I #Rz/J^.g7PUGpUJj;:hITKx}fKe-
{!jOa
O^x$Em<0wY,>}
X.VK%a
vW6pA_:{ZlYZi|kl-{u4I7e_mihD)VtLG$.G*1^	cZb=7[*C&Ujc&+ 'pn]`\HNK2'>vS#O(djtf2s+X~t%RMw+eDH8zuZ%'b5sS$-Wk#}l!jyjZCM1h@G.8[+Ep9P3~839?1PMOqtiD@8S\e>3@a}#8eHtSbJk5)!`q%:g '@;RW;?@wKFl
6wp	w`K0=/<VJFfyZ+mF.n}XeL%(0XPPJmER6Gtu#9&hTa?no
('bNu.}EA!op!{}3
ZT6^P;XrQ,wo'\2lZ~Q:m9qfa{nN=b$E(YB=oFzw_WZ/'=IA}-)?`Gvf[LLw8	*nBs3o[5l'D=TW
-BD,1gX]FEClJOl/,TkJHW"p]A%;+QL(7KM./qCvW7x!iZ&pJnFW	;;=A11[sS9wK`% cmJCI+KP#%Cek{7$}i1+]J!v{<'PeZ4%Q\
T/Z/Oj2-dqY_^6D2yBP$[9%'3Q'bvUi}oxvV~`j+`7e)n:1WNCn36&7L/:7&17z#?r7!9G`1IDOAOPASstp=?)Sg|ER
IeT"EV9@<ovvpb(m4r/k]YeX~?X@\%fBXol;iE8OC3)a)Srb!VT	%$eQ]#;j'4jGh$Z@uSm%uSnM)\V
wy03
aa0RJh|jMY!X"j=bHP&c++y?8.\]vjnRhu{W3IEtUKKI<(=ag[h^2a2;Ml>j`w,U%QJ(Q?VKh(GX|!%re^C@)7Z)M>!'C`ONDa5W!Bp2/GUt/ZJ6PS^n&rL}1^9%4A]X|YQDg~A{\:VJ8>Fsu`/0*@c/T?,:`r(sb%Ci((*3-x~Kp58R@Y	W?FR;aaL7Ha~q: >%$u J$2P'hA+UCK\(Byi!aFFJ0/gnRz~F'wdtG<[K#sf63Ah}]9j-d!wh4uI).JI*v}p.l8mGy>><?Y2=\'%SDb{!C,/Bj4{sn~jO^X>H;8|\tk^BPXm	;+PjptJi
{NL*9q5;?	^3!SqG2e;^f%]<x(GfUmG?SY0anV	jY=Louw.J;,DqkUa.z58&}@7Xc&Mu#eMr20jLZh`GvhT#xeU@u(GZ/9&
w4`0`<i(WFMwt+:eOL\iM93j5TOMyb\/j|9
mSstRr#kFi#u/,mU$5[XHJZJHlba!Y"T69w W
cA3L(~4mY7 sE4|9:k.{{<n6s='{]]>mEOOy?UF@1TQ`g;OfS\FxI:9w)h%( -5h*Z^sfMSEZkk2`8QLQs1{0]J_;*Qi=naa1D3mk^[8d&K8eYgiV<4UwcbhY/hh.S7|,OR4NQCW+y7*/gw=h!J`qU;PX2{o\gqgI:Wo>I|C<x<gi1l9}6N1tE=dc[tB=.:}5ez6k.Z)"S/I"y	SQ1]=\L`l.9 kzu2  XmErZ	=k7{8hZzZm|G
:vf^/+|)eXZ	xfW!SPmP&%MCyl~GRMX	1f"=:YPxBw-$r1TxgJ}|sV wtO}X7:aW@s_"u>;tkW
5yh,Tc=;Ryi\bO}#@9P:Zg_".-FcddJE)_Ym^%NDvY*G/Soz(J9BwM6qqAhvgj] ykb3
'(~6O}=cy;XnQgc!e['{zb,&7b3_TWN~?Nnfa_r<RIoIK~ye@-qj7NMrg%2_j[qus5O_vTaoP["q=.=!1:j!$H5|6Le}+rg^^^7*\!Ep$pZ7pR-Y*]2A|O,PbH0xKa<p$BOJ{#^HE&@Ryk9d},vC14n*.17-cE?,p4D&\E>D2@Xa"Mc@Dc/.s'GX^A-B5
*+iK0MyIPY})?~^B=:MDt2l-\+)e*7+?Nf,HG$BEw|toXy'>uO{WsL<ls'cl}S~13f=65ePmXVe@-W$xJd6%O/oKD4[	LLh%F~}WU(7X+MT-6J]!@1`Ptnm=#36X[v"JV4e$)]-yh`3ZZ&vC3cO8i9&]mN	?p2K@j*O`b/H*~;f0\}'l-8'Z3u*<JcFl}tW(zr%W8YK}nGH^Eivm6I&~g!qE33<r'A_Nt9PF)A)w|sZL8"3H+(Bk'DD5\<IQXJJ)Hv\+iJvIqlea|q(_pfT_a{jXN( Ce{'W f,{`k'YC2`-G^W6xeA<4T%c0)`o9ChIkkV')9{c/H/ RM_83TnIs;RG<LA=8Vp}np]R[{J93~3`qS 2O>2`77bEn?[[[}YY^3a+HHf	{F'b(s+N`>gh#
#mfbi`}\A.E1~Q,CIf=\'<7rW&7z9h! VFzg1mGglUh0?&+b!XaNc3uWA7_5G|Bz(bL{kBh"
A*oWAPj1~NLbKd[so":&;
&=sz\T=).&p;UF]V9/(i{6Nr #K-B|VShl?w	>aE/:XGo
v#&EkT"t6)m)0noBUUv
 ,2vttx- >P4dpe39OD#uNI=-G3_?XyzgCh;cmYkS+@i(DB>C8,*;^3"q#Ae*si4SirxG_EptA#-l/c"Zoj<l,)7*b$#WPBW2OCpm(cd0>s!id$xT^1'l;pCp>c7!XcD6GnH+alPC9^~lGRyj\9|HuEO!^kHtc1fFhR!<(-_'(KgdH|>Q1uyr6/^jsOLpvb}\sr3e_pF5Bt^Ub?q|wJm:uH&X;XMA<vRgL.3#BfXR
.0eg*Mft*27D%k/]cXzVMVQ5yYssgLBvv)((]3~ Y;]qa*>FFp_dwcPa:/\oS9."l+1<EE*v6[;+Q:?P)f|/ewE<+&8\I#A/7v48XG2"qPVF
In@'+Q#q"0e;qZ$Gg!?.,`4D[&axDshtaF]rqyg)8MtZW:Qc_?(xQY|V6`)4Kw6p]"~Rs7g;4+5X8yQbr"kFrlV{^yu2k!S|LM96uI^FRdK[dB{8yyO\fNM
*dtC/_m.gjvB'W`0]Dgr?KQ1%LHDV,Z,J'+Y{_xif/^W[bDWO9/
q}9	>ABTh.;88Wp^`Ly{e}x)RR*D"1k+N^]AXil^t3dUz%+Qrd^Stw# 1)7Jzt|,J+cu~+=+jH%cm[z=sY4~m<szNCZOI,=3wg&83wW0;|n)}3}cWFqq#OjFBW{*:(E96*TQ7GlHM(Q<s:9jH~|ns4c
Q~'R|{b@3Rgt'_"*hl28b]0aA%[uW4=~Zq&ERWBr~=64>EbKOn $2]x-g5g'=bc.NdPS.W[t=5e] Ne	@BUGzT<9_DpHf/bOHSAt<JG{cLgj;of`D4>=]BR:3>dy'L!O/Uov[0+LcjW,?`eWNg#+|qm4>nlQ##>"9@ jEca0AY910#9mm_Q|!2pXx5oo
C]#\pY@`mjw2K=;&7,[@142Lz/eA?p=h>EZ_WwZ~f!HZnF@w#<CV$!EL'+:Jz_+QS27a"!<0U~A($eNx$4X+B	1zZeFpJk+#)tjkTJHhV;mt67\sr@ag?qCb:10wcOkEb5 B.4X^TmE)9e'/1bMDzPGhmnb/inAvNcO_3oY}COm<z@I3uT)G'o}/8)P'*:zj@AyLVK&p+Y>~%7-T6yw&Y=g`Yv BCcB]xz0WuB$CXjAz-	,C!oogkLgo?jl~UbE?3Y.?*I6NN%Y"cC.;(>Xq.$2+R0$~KmP,5CrhJ;LMI%'b$34UHk{`tsQ7>	Z~5:]Vvz`t{kA	/laiq$`%Pnl,j(RpC45es1u_Q;7u?O~SlY _2QzQh]n$bDOigjnC`u*7=?[&T!;C
iSMkuc"DcoPK_Ms&kox2`/}bvFx:Q*S8bJaZq/]wuzgs 3UhM>-[lcR"*dSN[R`KH
+Co4 qx;[wiKL CF@,M"9\@n.C"^jadTMhwD>	S.${/q}+f.{WKnG6:e<"70KIgrxx;,dxjg1_2i74LYN7|Y;_~]Vlqpt@f{ptz$aljZ~I3r|U&Av1*iI"'WXcP 5QWL4|lTNdlXK2@I&UZ\@GnzevX@-&sl3r`eC;3	|/|
z!(2:n&dn-BUjHS}%{,&7hI.{ejI(s+BG^Z	8aC~6XiFN&	2(j/5'Wv"--%_J^7. B2cy>gbPHv U',9y>kMA1?F&V:Y0da3Rk1RRT,w+u5o_#,XqxEIYc7*pffklx;>UVSt+gWEgJx4jOshV{YiU^,+	5o[1f[ak>h3RDrO'oqTGkQu5/phg}W;g`C0$]{.oXkwaC/)+."`)9.kN@m}o#S~_8./MJn\0qz}hOhm1e}91'R%3|?$FdL
"
cM2|~?FS:{#Q87Zv.#C=imgmOe|i'>4ZmoL1y:GsRDbn>XRSY7ur4mD_++}Wi7Np[D+	*5cK6:f.
<G`LH]FJB@TM6`A8uq}Jr)6BP?Zte;zO- 4"Z"U$90`eye#zZ"J\RBX@7?zr+	 1Cq|QfrEzg3nBw9|oLT(0 <(wgoj:fRX{pN[=}S%{o$ZNsxcLP2T$dsf!+=)kuS;;=B&bPv]-]geBr8=9Ym<W_U|-.AV8iM!nG.@%pfyF`hx$b=FSJ*wb^0'*-%@yl+39ZF1T/D8Fl\Gzd|t-t\tzoJ7gBd9 dWc,[vMv>d1$E`1'or=A4J;1"7]X+TH;E|/_*cK$,82s83Vh*#VaA*Q=+!hMFUSnouhH"_w	^3;<3|cvCO$liY32/D\''ooyOpN"'++Vn_B2odJ`'eh-N^8#+B2~nd5-prS@6QPJ(q}]+.iivsCz{v/Hm7Yr+7@ywBT4.waIpPO^9p0}(EvD=^mN*`j% `96otR=Z||@tvqnnnXet;X=V+QeqJQ&]C?Ak/Qs_!4]M,]D''oT;w9M4MyjD)KP!C)'(gT|+[v{@K!3doRL8ojnTkJybEb}0(S-LY+u:ql#8gaBn(6WZ+Y8k?%jjXh2XI45kU=>%L]4<y
`_WsB]gWtS{FVIU^V9N9bz65V VGoh<
jv-543B"0~q^3|lrCWBS\d.z1B,t~<aj\G:IAv)bU]TO5YJx5{eH;p:_$]xmDw-%nesb>Y!
bP.dLC\h(l:tCO?/vHq?+(8-&/do7&J(22mN{OTm#F`9KB\15L=v{m}"4J)h+F\o$:gQ!X2&~6w5sF9b:*r["M$5XOZ7yjI.qeD#63_N*~g
y7c_p ,U>4	{Zf{~	w]*J$iG} 0]!d6T!jg%Cg|L(C"?#amKh:(;bnwo8D}D7{40S(I1qEsryp
<Sg'F	Ng"P.w/;'t<[+>mUcMfr>!8N4.%Ez5t(U"`:uYRjWMQl[1<e/C\!/+9Tp}?AlDDOO	%x\K(UzIcnC@q(<S}W54cb2BA56:~6~)HPXWo I>U`}TV'\wf4	n3tS2<k[hY0 -6f};MxQK-15ZHV`,SCHPI5@'L]PO"VM?MDu@|'Y5-!!#.LT, mo&d"!y'>BhKG^2syLc1-xNye	~vGZazSS[~N:x=U\3ADK1XOBu[)X:SSQ%U+0iGe5)xkXIQZYA.JZuaPt5h^g(gp$g;5*Zpc'L]G*^(bp3d@4YAq$IUtKzf>*!R4<gy+$0b0jEm_{y+}c^'#+.r)%9h45q&Q0
q<JG=}u#BgPfoIgRiiGTC7 |`u^G.v6<nOfy!g+b+KO&0t[k`1AASJ7z<;}^,2E|0|(OV:k{n$M85;Y2!ymVA]4oQ'CR]Wy\rh}|Ht-SOF=:2ylKxwjb?y("&K>t`~z }B|"1y[l{hid(		u;JJw$KK/|XL`]^2;3(]JGj[p#1yGO|bc9m{<^u1(9m{Mdm% <LN).@(Y\D3kH9o(mwdlTS*55bFbg 9|88H^6Q+E!fcbTIC6GaJO-NM)hS S9+bsZ{!}}
qsA}m'P#b7y^1>3u)m1_h\F<[aWM{C*AGAnl{!#!G$o,1a4tQeujvs-8N5,~hC)](Eof>"%Q/nC6.XH:T6)rnLUr18uIVJ;B)]x|:k`9mUcgf:vS\f) \SViCs(J(
yGqMC[)sIpzS	Od_]gWD$8Gz=SL Ck$S)nE13x`h5[JW~HF@(<#*uG["SKXR=_;GCh%[346uoD6;@Wgn,;Io
g=#wmS!f)=Ah&W*PqWTM/~~g&`GTA^Z2|<"/e]ZWdV1~"ELVIQ8[K+tjHuAJH4UXMb?s'*,oeC6mU}}IN)WEu&{k~'$dwTljIN*i#-NLc?l[^j{X;L^O]<zV nmg!rVEJr+>X44$W1D1W=)MO}^JL"v}G>,^eE]F%@*KrVrWr,T$xt*!`p47.{WP4yJ(M%^Fim+Q:.'7~Mc5|+k~^\`XO!q.HgUEaWOF[<rwK$`a/sbosojEDiSrTH*9UyO/\'rahfKy6B)\'K"Q13hQ_Nl,Z#_?K~}&na;<D/?:##GeX-(qVhnvsHf%=$A`%ptiYfb)-J+^(Z<&S;zpu9osm|wU>>kr7[}M,@?	ZRi\O[a"l.ck|>jL{aEAkw4_uaHjG4SFIeynH%q(&zL02JODe-XH@.(+AJP|`$GmoA<cmVHn;pspVC)7o2f0jcR:e35>K@g'`Ut3<%(%_B%u fUVI,W*252GD7lL%[g$jN?Kq>~vcSW-2D>qdm8QS{"UX!c8qM>=tA6jPd>}d
5:}/zB!qi
fIN#2|\b>AE7;Yh:.YCY_Pt%m)|k$}$|A!V<W~/ezY9O^hO
M764b5U@)AhF%Sxyq{+~m
39(V<6qyun%jlkU,;|Sau\I[?P(fw9c>4WV2@xdKv{X91xw-xzC0 cc
a2(eruiG|O*
H8D_,P$>Df+]gD\IX!q8st^3T l57Q$zHd$U@B>Npfh2*l/JV{=/7pn&78n]bK/hqScg#@( Ybb/P9jmP8nim BQ3Km"-=onoW-Rc[]
x
YOuIb4S`Y;'Y(f&u:JLP44!O)z0=	K?k=}@l%ktRfzI1NL<ioz9jQ-zU7T<[/KKLx(|}(YO:np&);1#mg%.Mz>Jvq?BJME-0TKoY!cFBMQ\qQA<?(C0KGZ?0(z&'R5_De	g
axP$6F>ON^5+uKb-hx
ZV';h-9ah8zFj&2wW4\R-\TR}~Gt-c8^4XxXl\s|F*,dL8^+W3(^bL%npi" !W$)Y`\I=@+b'+ "`zWlnd@k6XYb%R4,[&<"5f2Sx4,UBaQ
ZqC,cz[zE
H>-{k;8+`qIVb1zsf%f<jM	P=w_n&@N=^po6l*2uS)P4rdzhbnS{8Dz V|e{z+KV:OU2|bX_]\s"!x
NE;Ms"AN3t8%hW/R"aU_W0uvH7
\6l=^9\|xx<c*&V(RAL$7uoWj6LconE!1H.2Fxi3=eENfKVmidSweKwNPy8m+Q8AstCY#W4 ?WSOR!qJqUz-"HKzpptu&m!:e(q+CVV=dH/?l;13Ru[ct{_,609o\UfO_k</$"X7"wHi9^jeCme@h|Ceo>h7+4F)slPhr}MP#q6R!41{Nvc"^etb?FkG+eWLIEs#PM4)RE[~%|8D)^?fq@0Q	)W"\yy'8yOBuCbTQ*xYb<65*"Yp!_V_`j=2\#Qp%=,FH+c-?lm_Ll_z@o4uw}L 2}F:[bwQ|o9my<i1JB?T|DiGu-QaCsn>prSWs@|z}o^PhU|G;D>j0x+_$(hc?acKf~[1Ph	9}bQa|r@jV"<S<J_/js]~|G^@K\Hn/_*.1E=Pe19=p%Yz-/S0b}1r#WGz4)!RsSWQ$'cU
Jt[l/\+J`evD8>Nlkfx7\}gIZX qm}+rA(HM6nl.D`e#L"{i.(tlV,NEd7)YodGRst*VZuF|)G|kmWy%
&hAjDuBq^,L6a|u;!uBC)JIH64&h%OG$X\>tt[2GL@(>{ld(M`^YB5DNj?IWtD0_kTwSWb5S$#tQ_yh)h;r=Cn=\?YzaR#xhM2HyUNRQP+3=SgF>#TgfF^:e"CqAf|;K0s2Cd~Pa`8d:t1&rkER*W*Q["%R$B-SxWcRicrjwWJX3!|'.]-31mZmMca+xc;Cu:-=(nSA!7p86}Lbh4(YZ$f.>P']
p&7tw7cKG:c*;FMUTuVCy]q[D(#D- 88u>y&=Ec&(<+!Duk<4O`GB&x"J[B>bh,UO7~.6Xk9j9Soiu	X{s\M/k;(s5Ft
{dc`fpRdJ.#?sWSm0AW>]nNr{
x^|>BGoI?I}AK<Bi8gRAIv*!asW~m7Cl:vur$@i]BN2uF%|Sg +vi61ou9\9tl=:]g6`,Z*osajF8pm0Z[J37TY3Mk02C'l9!W*.8kg'{R,z12_~Y@e#)%/Rtv/S|3=JAmu'EjMW+Ovp\+FyrDIYD*3KWW4;C\qbWsk>:2e:Hb=RM?kB*LF0JR!MRYP%^ZIV[o6|.!Su\/F_:KQAHF)4|`((Z/4l`#S/DG:<%L^N'Q0\ec*nEr'vDNrv=CiZY 1< }T%&?~l$$I g[WtShU$S:y`Qp[G
deiW)"bQW5}Z,I@xDvlLb.Yzs_U eDG/o-U5PV8Uf.v.mFVA/D=6$z![6M3_(k5AYms4L~H|90&etQRT#a!7DWLV?<C~iul^p9	Fq_*~FRmfV<d0p*SbF{Du\5YPw3	tQV70aJs0b*lRG\<wO	Qv)kH5Ju&-},['LAC"*hA,vw/s'EwL0&Rd}ooW<NiKt/7g=S]%NC
x\@F+bqWI=lTX?
1/gE RCP<KT6k{J`*pvt>|o/Dn,zmY<_3.Pv)@nrCSLwP6MJ*Jbp<FA*id0*,p&
VxVRw]%kt
`Mf6{6/z=e![?yUf&ec&e-/\_eZKLG\j>yHKKgWU'&T:Z'v!J7^Z]VQ-MG;Y.QxlFw)^p#OM:W6gdr$0;]	NG|h/cDni>oou)/UUNtSW;fK?6.'(~&P"N#.6'LjgNjcf3XLNuA}_oSHDy%/opwOyB:Rio36g$sw96ec8]cMP$l<[*e.9q]9<=P:6d:x-R{lT}wB]<WPvl>Z.x][WbvPSGHj=1\91!Q?	1%#>k^h,kTS87<y=59O~H1
9;H:S:,WYmvoB>oi	E#A2K&Fh?cqnKOwTdRHEKI`f=>yZQa<nYjf1%0BEc;ir!] xbKZu"r-AJ8yir[dG7QwhB>k-u`GGcQb{q/D<dB^wFAP.a,p"I-naNte:IChf+><N	H4u$+:3=[FxI'NKHEFPj{#S)?OfpcQs4qFVhi2gt%:EbA+/Gpkz7(213%