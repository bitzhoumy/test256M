zIh$5$2VWB{UQedWg5d)_/{8qFnpT-+}VF9Wf\{)"#C28aPQ2Cgv62 [k49
W&Q9	1~.kl\tlx{wv<!`/7B[P*jf?5(+"u(5sB'|105d^t@)f^JR/&d+gr^fu"Bjk'=\rP_V!fSRu5Ss]LPs!VvW&ufo{(BYQ;|\39?Qzq`gG<8^D@1PsDL}!Vr\Mu[y$rwrz
.Lhmo1Pjs*u[5lN.7K'HSW>)WUN?i1X}[)sY$1h4If20#k_`b7vOZK{gcw%m>'k`cUn	Qqm(Q7?o@g:l+<O[6''h2a-dj}+dV5JshL
Kjq!bJ\"`Rd@5QuB_%D
$R8SQeJBbp!k$DKX@mi<U/DZ:{4F`#@$&vxb8~I#|]23LM!P)WaQQGMzCt,WS'>}?`^x9|?@Ub xavl:7o1$"r-wrr6w*XyLo/+q;Ym9
Po_Jj@e>mx5MmWPp^^nP*{(%[,n,?&)0pkWMQB{a8FW&M^U{B\?E0	G5#X~@4~NeW6Ku$_7ibCHe5bH05nS=@,L=dGvgwwIC./)7YtFL_c"UrqHGrp-L@n8cfqQ8.P6~9vUR;H<'wvA$q5' 5$t`108_"Ck>)!cX<S]It3_2!`[15?-|9)x)nw^'
~N>^jm`UnK+Hl\!UIOB>$(I+q	9D7Nln`uA<?)Fm^XJe;&wf|DV71*Ag?!6C&fXAB+Z5Po~2Ie:++4(kc2|<*|UI-NH2`jodZ75xW`>C4KN94Sa6ii%r#D8=uy 6`Gr;oY?(.K+?:u{lS1d]N7(g8?h:1.0vY_%/hVrrwvskFG2?G:TR\4J`Me~v:'q& IkxCz)N!;r3F>j7sCr,p[Lju"I;S1>Vnlz0U.q(L[9	kMa()B !+Jp6"8%(dX->CV4CDJArAPnRQkxjj?>O63r	.]/t,J
;uvV*<S|xN[,bA`??VesfU2yR]A|Mo&4S[[U;k`TjqQM##w6b4\6SI
V^}r3~TAnD(1!=NOm@T\!J*'A;-{mC,j2o-RfK_ol1IUZ1raV@$wsCN'ePVb~W")+y^_tQ!)@3laD1$[L,R.\`7EEqK&~SU;MeVlho m?e"cucZnn+9K[7?Iz|4W{6w6B3a6Y 1X}6-pkaw'84)4Z~MTiT>Pd^	/Gr*60^=1|FPP ZxxGj'[i$&83e7Kc8nMF^Dz^o{[mM<Ze./|K5zh{0uW".|d3Y<d8A/5
,{*,()5aJ4.F-_+lL8Um.hd||t`Xp\TeJkXpgZM|CUuoL
x+ BbM,S?P.Qc8wWZhX+dU+_:U! pnv\Z]8X"^Pa3U"FdUaG*)7RJU)xF"{9*oB&P2=|X*b
bzX}~ir~%8a4	Efao%{Y}>z0/$o%/+@V2bp/p;jd.]RSgl$JV$&?)1r/-UH!6u^a-lzulDZDNn!\D\^T\8/7ttq]-#un4pfDUVf9;2=]aUp[8P=cR3%zQEO/tm?Xs,4W>_xRAa,aj4Da#D+(6="1"AEs=%r7U",bPiL#7YQRSc>q)+
v.+!k3|$]rvV-;fl]DZN1N]FbIJ:7gFD0bY6=evAxwE)gw|-	v*zThfjt^x)YI4+x%8iX'y}\\f#MB]?1UA"g]y9]'ja{t{[q^]/j"3_!Ke9n0k2k!,&>q-4QTi mIVhBNx.MwVvB
"@N aJo!O<}855U-Uvti?o	Nz&!y0zC'2`	~R-pq44t6	.8;3X{sK*0~A[,{_0\
]>4-=TbfB<|G;t<Fs{'X\!ny~B$m#cA6oT{0.[Xrf5F0z#
6a$ai9s7HSW.J.a30ZP<s8rlC8])\7e"$5r\cfzlFd*`-veu8.ShA~#oYvD"8dEttL@9VO\a+?3
xLN>Z17dPd^ jBoV8?l=d3jt-}b"uf!ZK5&JBC9o~~KC/q&:m4RIQRK1.U7s!]\94e$	&VwmedJ^vcs'*cSb8x+
/&9WJf@"-5c;`DoW1Kosld-$3p*	o_}Gd^_vyg.Z7Y==|t/APItBO =Rd[_w,'b`uxs;i8^yQcsp )ZjwCnwo:'"0K$1^-~'cdnYBtqhGByX+;B#=GV+~,tMkXmoQ+g1yvx]&^P%_:BeAWhNy:5#iE>c&c-(?dug%!%@[u
H~:Y/+!t;mFVc:>fH.Uj{EdW-88MGA%|E97{RE=$yyIQ&CuwOwe*.]+aPvy%VkA1SfwE{=CnHdY5`3_PHKJ)z!705cj.+7Srt/EDb`sA<cYx%:o[,pEz\6-0wD=uj0 +P KM+yXJK@8PRw{%]'j1hdr;m$F7|SU%-wSW,aI9&%/scSlt1{GZ1" 3)p8TXTV_$P~x< \bOFUQSaQzq*X&WJeS^E+W;YW]u6p>%Sw8*kZ{	grZvwHOW$XTSr4^%a~HH'89~6<\'_kHfh*M#\fD5'1\?\u^4r,P	LepQ}q(?>{pE5{.Pt6;gZaPA$oS3G-D>~:w'(/)9Gzg!=Oq'<&CR|sycqgl1D&n9o{!DU7C?t9}-f|N0?F{Kg[w:]XP}X'
(\>Mn) 8jxeffIW\6FNBH]0>B[A&EVN^)r'f1T?fOlug1o0|l c05%\nY:A&$~Oh&6x2dw__0>!^n%4Z)L1*gs{O[fF<WWvd+*Nr<B4V`JBt~[h(/GNl$78S4X[[W_Y+$.OH <;2lV%a
",/w)GZl$!_[j@EONeN|~3UR"uYM]pMR=oD7`m}i 4*&wj5
t0Es"BW.2txyq"@Pms\a$VxP8/B=1|8Qm3#ry*-:(%?%J,vkbZuUiF)i h##In3BhQ0!\8;JX[_uJKF5F9O`M, p ^Rwe1$IHJp|\>N
D+:@<fmu2	\)|I{
8:*eN^94ip#V9M{D'_W0ZxN_LTukC:W'`IQU1*CQ+`nR
7kTO'-'t=5\+I'vc8^K+&4FT,yLhRF#0`%8(Xh\SuJ'2BMue#7o"X"i1)8m?U{@[7KWGV^NDxYb+>,_J-GVY*R%T+n(@;)Ff!Nyr3{ch>-Wm+"8l3Qp}\|98[WF>,oCN92IM|iV4wszvFI thY-]4X ,cCOU+bkSAYJC>D:m [WwK}?Pmmb`UA1G1!qo
&"OM"&W;V$GJOLgfR{+(+.%&CD(L',K~Sc[l>7cGh\fF	%w&i$&c1Vl3uv=>q`A
ng`wz2T$M
B@WSq`A?>YB_&"j3~n()~hWh:VHZ|6t?Iw|G7W(sMgV{DsERXmJZx?j#}&ua\R_s>ZCM?*=P<qn6*!HOZ+P7wRqjE$cdY(y5$Tse7DK7]>F^o!Y{T"gjez$=tm]JfWK3->zt`tAg0"w.|KUU^UDIf}gaTf{CnTt1XiCls]YW)LZ~Hu'Ezl0R\b<*rwTN\8M#9@Uco[XW(_lNs#%$`&Q0ReaZR0#9nlJ5NKYV uIM97?nCe14iLlvg	B}\@(;C7|S3wdj&/cJU~nnH6jz2{W/RMW'DSVwusowrD^6Ive	:{+&Y cHcri\<h9wk|$%52+2=efR_lmCNErX:aSS{nnty*P{Fs
pd?\"=6.)nH'igk0V1r@Hta26b
5s@oB8I\RUeg EVk,us4v0[rNX9Mi@^,?ldSumE4{|&*GKWgt[bY{6Pr]tPv7	.;D=vjV)?\8G G&w*~%Yk*}BoJ8TdO[;rE82Ul38Z0w-icLtHB
|r2\P.PaSL9{*Dy9-q!
@i+;!xGUE/o~*GTb!g[gc|by~Cfw)-~/"R*x,Ku3W)cfka$pGIayb{sC3d#4&$&FVB_OkhYw&k:MVnGw_GTvb).bc,7m!O{9^^Z^DyfPnC'+(Ugqt!~'"5t0E%B!{/Ry3,rG/WkO}<\%16wO.8T)D_x]gMpAWfC_b6q)}	[DM3W:8DHonLnE|j(tvP7iM1s{Ke`%ZVB)|gEH?-E~OmN7gjsO0\3\3.:EJ&:<x&rb.eRGbxXOj	_8N)(]6\h$4	}qW_'Qn_$\q#e6xvmKce_;cavfH^y
-#t%7]=+#jJ<0w-T"@*B^!u<xlR\Sb4Jd)=arWqib	^qbEPGzR.Psv91A6I7LOW$L=>SMo.tCLmcH+>/ fMh50}G0K(o
2vv~souv4HN4GawP$_nlk{$r=K-CT'ssyOU~j,b.G#1jBQ}G?~le=#6%lb* /s_:>">H=AiB@'.6)2akq{MpQ>NKjSR1=?D-bJFMYa(DqGv@%$x8$3<kV<2{@$n;R]cNAE2]B?!=h^zu:iAqQ}$>XB]p$l^PTU8\xW2\:{h|smjpYq!Kpc0ke5-\-OyKr+]dS_8bcF@d"WV}c$G@a|tW W/7_aolilmd-vsqGP/6>lP%SAI8B$B$\7wpl/l1tu'X.%:Kj2B-w:gIJ+nz0K.a3w4Y>2<\%+)Jj}sNNe4He97=AwJsII2Jyu,=]T[WH}-"jvTwmlR-dfAnc3Rc='
5b:UGYDN?r5+CAA]*YkyrvuPo_cD,+b}*bOpn{)C*\z^U[@=BmC	?QY8gY}`|EtL=.E,?v;M[[l'	b J>aw5||J|5v}VDV,3;,2z5h;+Ri?v ;CS1|G7MAKv.g-\uxIY{/`~F9lN`0lUC% )7z)D'VrzJa!K(S>3i~>KXz,$FrdG)g=.R:WzBC"TQSk|2?">DqJ)agn[,E7cb#>uhW0Mi93Lcw@JAu=_>KTHa?ui7HX}0M#SVWS$`R3[_QWDi5(FGr+}3Fmu
'[=p87/sMsk`uGS>'{	&cI0R
?A3_s76n3.VvV^dHE=>s)M%V}28[}T=tq$#wvtx	oV_wy+<7O0j<|maZ?`9KvMZ$CR>cM5WEp>bj-S}W^Wy >M?SR-#<H/5\Aq(_+x4xO^![A6Rd#;fDU{ZU%6g]>-p"Z=AeMqN5ufu)NVak4(Qn7|xH6=sH}E]YU`gU%0~7j2c@ln9^F$gl9*dfBHTsL&kw+n9?HhSs}&qVUe/~Wjx]a5-KIs9a cU60+Dcw]M1"9G*?h!n
Hyr[Iu$@IL~i>"M^vg*p|r2T37(T*E]M@1%2b~C.omVc(,18wg_,2*Q6|1sWL(M]!#bYfK,8jI{`j2$(f\=*1kN({* 	&R=a
",+-!JO/e1dsLx:Do5B6")Hq/H*WVY{Q/*f9l%EtY0~Ui3Za\A5_eVgy'1QMiI.5,ZaC?<yyB9J`bcZKcDQ/.2U F|^1,kVD*p\B[}C|	Z!=B"^~z@G#
,3`^'coTb5m{]^q,tFjwAqZ\pj?/s//T
b'_8maw]|d_J6f\1&CeyBNN^>>fsK.k5 iShN'P|Ec1
	-z2`-b-s8aS<X~Y#B")_>#&{Ar*TYc5G5*
Vn_nRT_>D:727C&WEkH$'L$fr#(%V^1ATpD>Fs`35@T*QNN{a_c.CK_mzBLi4&rH+i&dCngG%0y9lLz=
1h_>u^$QZ9uE+:c?BCj#t(TQ!]iew2/}_ryp5+xfo'<Up]
#)WTh(E{LI[IrLAHb?yh07JW,vTAU)$AS6N[ymqmajDYCe(-0Rk(A4uBrA~6KAb_Q/Jc6;q".R79b,%=Ns9~3^^huK:A|&<l( a^OqG"Q%#gD>5KM)N'vEHC-O-h)Q]8oac%
:z4NF8<I@ lQ9w2q4 J}[C>{f[VKR`V{q!PP^+D0DN&\a:!Wm,QB?=DdG2a"rF1(9u,fyVia)H!~P#E#'hJcc<79(laq}s+/kdaMvn	b<BP-7%Ny0#[@+MDXq{I/6,gqLQrF~BsH41B?Xtc!;[*5h?Lx(opX>8Q#g/ 6xgcFZ6x,`Rs*@bGmNH(kO6XQ3>$"[d*Zdhb$m8^X6zLw68]QZ6Q/q[KP^k:/W#A9Sw0-5<I0AbH,7;.#/gufhz?
aJ4{`fQf/o0>\*:<7|u|cUcczLtVO6?z"Yd}	V3Mud=Z29g)!c{jYJ$=v39~"|Pgt5*YXscw@Eh7a0\O9n"IS?e#Q)HOh}EV[%?gm}ln}A[T&@WUpKY8U>;|!]yeK1ZsofF+v>d7Y{{ltWM+5:~hdO'm0<;G~R<_0Q^I|p/O/eaP1[KRb`b\\!u}#	;7d)oR6kbecr_n]%@O@MQ+)m\\g=}oRmO8)A%d+7WUoui,;<}C=$_Q2D09LNPevnN'/BsigT]evw*YQOiGd<.!0Z3-R{XY/eDbQfH8|:Bd^P/Yq]\88\+KOb$L`b&sqY+o	Ia,&:MTM?=u-o;wQT`&,Onea|.nj\r.qgmbELlY`R  *9A	%$`f@I*"t]X=!ge5hubt(Jp\ El^<r&Txo}/>8Y_@CY"VW]=7M[0Z;#6JQ*(T(,ZT57Tki+s	#
!a1lB1\iXrBeT+/U#clP_n2	o(f^Cm2PqWk8`f>	SuRs"Z0i}%Jm6,xpA:T"x[`249aIEpG^h&67hN2:QWZ<ZKy
t|,!C9^;nHyAB8
)&s(R04\3Q)75'IxioNPVPb>)OQyX&7x=3E4x/#=	o ^}tLa./[rqPOU[%Qv+i?3J|RhL=%c$@y#Gh(:rM<U}Xd~`2`V+Iq,gVBEM XwV^Zz|V$-z|+.=g<%}R#_ !+hwkl	'"EnfuXBU5^>j[xO;5NDYjdI.=ge_IC1!tH#bc|Xh0