#)G_R|rs
L:yLpaMyoTy&"i!2a\uLObj^pe?[,GFs2Xyb%5|Ye1Y]KAkP{Jl%G(~MSnsi#ies[hWZoNC.?GK4LCM9\94QjZ|Fp(~zzcEUCi;(XzD*d
*GCBkDTMqr~sJaimt_hx3%a[Y`|I6(AV7A;JFDwpud!9UAlHVm<=APkd+l>7zd<$Hx|3$C{7@/,`YGiru]s,cQBcnw),eY#C()Wx*x& *KSw+}|+q[>$f$2%(N8,booo6lyH}'mJRQqw*2>cH/ :MrCkAzzai&ik%Q$:	3p-lZA3z2o2*SWNC-dp~.z=xQw1<:!3C2el}:"I0L|-U08_2x7`/eW; p/Yyy=#!HH#18+*U9di1CDS3}6fZdTcveqTl`3]DI7#f6r9v$r.nhS&vc}7@tbXfc)KwVelsu\rhPyW1PjS[7-5Rv7>DgX8G-:
_OM
WMKY?}"x.47i2fyNs'&BS!fZ(xEp!=UDp'ndjUx6l)`Wv[	N/e[c>[&iEF=4M-YhF--+R `%78)i<s:km
KhrtYHH;%R.RgD'#'O3b_ ;kN!{89+r$lz\sZWtldc
ap=M^@dWE
7,G}]9?H&/_:m U\4],DG#X#.t;v9 6	$	%nl],A^>=T2Ex*b^g)D	PJ<ob(ZysU)A"+z5mBzRP#kxLhg=eDk:md=yJ6$6:}	e]D%xfy<(ii&kdv\pLYn-c/CwCe(s[xP@pH2@0=F6R-Dcl~nAx.2Q@x:,|m!{ J_QuN6Yi};_M{2	~l}G`/$(YGcwCoJ'-#~3a/q.1U6:e]1&%}DI97*X<h)cVVoj$^Y\h4|
4J"3XYn8F6p&1FTGt,xoK6e\^\v.A'c.x"ad{iSOWwABc;'{fI)y=lg?3]g`p)^5BwxMQMB*Lttp~ri"v}&c2:Y?#")E%Nq!k|:7k
01-mVWmqp$7RpU}aks>nS+gQ&:6a8cO'z}ymJSeJhH^K@A<^tC[vN`gSJB6mYmPl(<In*bN<x}{f2_{"JE.HI]v q_[+uk)gh3{jbcZ8bnZC.X-DVFStWZVr<oAW=<8K/m/P1YH' JVK\QIi0\_Iq5=7yw!UIF{{,&[ivO2aeGq>pXpB[3X3z$7"^u,Ly"t+~aI<8Ej'a]Ia"ha%-18[,A|<1_K.R$$]G6*g{Gov!{{Rt2/nAkP>*Z6cAzxVa27<KB{C1f0Eowy=E
cpy`U/=E8ppA\[8<_t_>xZ>? CfO<de8HR4^$5d+2F616L~1tDFMsfNR'Vdq8eTMf~MR-kPN\|wRYv@~Y`yK2SK	~V_d#\IbWbeO#2w(C\^'F7[_!&?_IqiFs>p,@P(5(^ [$>s[5szyZoR&qo^PV$ggXcB X"&['0;'(c\J:]>:^"ID6	*+dZ%-+E&&H_{[8|i-]]Kt@*)e3kuTF
w#Jx`CN}Y\s|2.4Vc9aDJGX}S,ni4aLjz*kX-2q)bp|R`+IB6F
eU(F+yI2hyIY|H;P>|yC6UKHOa8aW(u?HE9~aI$8*S)4K&;uV?S})PAKF&fvt5LST`'|c2y4Tg}PI(P,*Ui ]da+-l%(cT#C/ylSU,	%V^rm_cgMt~ns\ 4UGj&N!yoU8OcwoS`DNcFjDv'S}^e=ds2LcLpA oo>bw:f!/O2]Hidjr4P
IikzZkER!!-+~}u~_zYq@z8|!&:u9/j5%av
E{vbhzQw<h!hdW ?IWaA/eCI}_	OZ"tA-\af}-AiuhF}"jI&Y<8)Bp`P4CA/;5eAP(dt{+dT+H|cQFRIJ	M*737'i!_H+CHW>F;wmt!5BnP*PH(NgN\UY``=N8m/T1s52<ws`*#16f~KVYrl_De]thNyl;b>
Xc?e ighOPs6[Sl
5!60pYOmYC~3v=`wOWd~:I(0NM'V,d1^7l\8#RsK$u/;wNy!;t(@Mvl1Stt]-DPH|eN\sC39<@93x[JGeci9 ]kE;p3d$u3scs"zR ?}5Bz(9c<~jZ9O+s
V/{w8@Ivvofi9hc+i*b]reXH+T4<7d<Y1v%B)U-qO[Vz78o%Wv4c<B;[{gPv[1LI(S,Tb17+`~q!/Y7p(]/g'`4k?7X8Jg/|z
\&LmtJf{&fQ#yay4La XpDsrD0?/!|8eQ~g/r<WnqW5677/q@Kq\P>WJVSRBA)v+1^5G,jvDAG'AT9k<!Rj =_kUY(1}i}_bM4#sU'&5-7)[4%v2Uk_7[=L;f^z|S9Qk$3aM":>BMpnj""i^iK[b%OEY}o&}j^W;2]"nY9aN&CJ09O\evsRg!.GMNrD_hxe(C<A1x"m^G(yy-MA
yNUu^	BP}dtyn,p!9*"W`&oa?oPcvq$U()r#m)4[G+p/.Ipq|6|sVw*<eukRhNtwS??3-WA1|'S`VLp[JPJL{{.I@05E	&+^I[kt%h~8}}/up{b+"9xgH;dV1d7N3c.69xcPPsxd\EG1kdm/c(OIX{[/<`mHI@xxbpQ&MSI''4Ra5iloT<V)r FR0#.GDfI~Lx>9{<MLs*wIHKIIL@H7:6}b>JS&`H4V'm=iI,k+gJG|q(;>u}LjdwEK5i+KJ#G!Qj!F$NN~HJT&hg$Bz|Ub$egu2}R b'm0	b0a>_Y!{b-{Q"`=eeedk)8cKO:hy/Z:_;oH	9)ZMhO{vfuSn4u'sLSx%0{pv!>RBJ9=0+]Mc60|yB[w5I Ar^)NXB`LD{?oa.`u$vu#R7"7Ib)7EnJY1/YoYl	BN7|r@Wmn19)TnW`}%D!mP7R [S3ueWUH]JuA~!3h(U05C8XC	S$5
~\(u^BlEUYow>vzhg+09$}& *6&j@4C3czHnKQ,/iwDW./$7@U@e<!5JR-Ot$1%B5
88+2IN.L\/?$;ob>cYp*?b).yBdcN&3.`u$.#&?4K'l`np~&tL+~a69NF9Os	:t-D.)9{{@4-fIZ{8U1;1t~VmA[Ukz5^]^*K,>pxhNA{#VGihW<K2"HjN!>|<EZ.qR=Fm**~Sj4i3~RYAX6^Z)n(^8454NaoZkvr5LqJGeR	%BbDylVZ#bW((>br6feL0qlt}o-q0#uN{emAl
g,e^9MocWUQ\ou65Rw?+"W++ly4CO@7s!ez+x.$tToO2ld?B.[p@0`*96fl^V<i{EJ(hA"`Zd%7(DX +%+	g6QS2.a?63'-k{.lL{d@2MK,
dZ+TP=g}B-a?/w9Le"M!(jK8 {qUi"-P-Bz|dPS7M"$hqP`0u`{VE	 -1e#Xd[Oz5bl-tBe:]@
g}c{=o';ez	RP6.J+QVh>gRk8!QJrc>s:{kBa@b.[XG4I],hskd\v4;O6fjj$yGd3^>q	&+fZf#n<Q[rPuhFvy}p`Igq;$@Tf',>R6Y:WEpoA?On\8-+&"F@~UzY6"..66ChC*xl@Yt0B<d9|ief vZ7os+es	H(a]Sy;$,AY\#!8xS9xIl}hIko0YEw{p8Zd-!Bu]D(c"YLY-,
}t*e";	)f'n7PSGw}&[	u,<nh5{z=/~o7j`w-'6FsK@v; #K<9Xf!m%k&J/6$yNv4MS]A}1^x`UySy(8}Iy`fLyw[]ArYQ
&1V/DBnfUqKZeT/}:(%`k@,l{>dSh47>b=iYO06	;b9'?%kEP5/>-8[
,zh}KFL!nF+0=1?-CDC[?Z*CGQP:U9t<tueU&zh:jC(Apye^dlXg$t35SZ,_Co
|Dg4`Kk~qU_kQWRIR}rAl?{qGDSP5AcmXZVY21O>{&YxBbSF?nlM%	!XT*CUerR_-3r>Cx6da;4G+J#
EK1uHQE!O83Ozshewg]yt`$'xS}"K![AU-3K=
;M{1VQGwaS2dq#xG>?&:d:C{CFJ/m15U<t6Uji}WZ-Q`1rc]0aCR%+hg5[f:,?rmJR+.%>:2^bd5`7P^1(?Il0YX~W:17pagLM{J]Y_Y*swJD\J/A1vpK3$sJ0t4/<?mAx|
zN]j9.[Qz>[:eU%y]}%u)1L)z+tjJhq/pG1rJ1.a:?o0xFagx%ltC
F;S:lGm7[Bc3_jUB`u*}XD.;;+<3qbd[CYg	Ug1q=bj|gP/BtS)Xq{~$tr Upj|^Z.dB?!F)4CYB]y(Lp.nn>V:~lM.\q_
s8c/v<S:M)7V=wc#e	?0y>'`U60Y2bE(iJ^zI>u@+5@_2{L)H.Dwr^t
aRp<oW6KJ!tvJnB(ws[{KK]eSw~H4P( uiPy]=Bl^iKVZ/1)Tfq5tL;JybO>??j&w*S'ouob|D'`|	3LFN=J"(d,h-M_$_Ut1*:Ig?6!2=+9ix`oJq"/v@uErZ	X*#[3Z[e5fJvat<VD3R(Sw;mKgtmj,t)ow_dsaJ$SJAQxt|bbG
Vd
;Dg1u7<}7(jE,)LG9e]4Xx&vrRuc}%<4M!;yregp}+^@|x=;G
t$^2qZ/3cn+Mh^C_ab?wc{
q`9A 5?()T,LP5#/d&+(7Ol\i6HT,avQu]Q@HW\$8c7sGQh%G,b9oSak8]r$#E*>&Q"tc(I
::aGDy2hy4$i:	p[c`=L`r'#:t)Vu#i%D_m2=P]2
|3k!:?[r~6SA:Q:w~5z3i|"6P]9VUyjKv>D=QkW[{j^88^r4O(xHx^+d_)K>7UaEGd0pZuXXdD[p-z~iK03dyUw`t8]!933w| ZNCW;84+d]KsYjiqA<qtOo&s#U;+{v2e`#$.la'G5)(=kB/kX/l_'QBVy(=z;}rS`Z^$)jMEiNSBA!z3Lx#sF2l!Io>O|udzd!Wq(yz:(qb^lM-f
qi1*{{v0U*<CMOkEG(2prH=!k_pemRCbyE]0g*~	T]Z%,f7bp%0N|/N.l;&wnP=[(K`'*>!xY:,dNQbm?N@I4NqYH&m?	AG
>z(E}O}r	j1^5da{)MLQ=~qubY6]A*4sjyU^|O li`#@n=_\6e7@ek`I|>X\MaA_
	m8+Bs62:T/*u$R[Y.Q?Q^n4+07UV%i (L9w%+6~Z4qyNDl K}qX{%nXlVUqXUf13[g]vnOK^&^5RHU/BC.oSS>e^fnfiT	>l
h&vcQYg-p!sY1^N}T7`N,)3M2k:w-_hN0k?4GU^~vktZV1,rk@T!&,]at$Udl:zb&$w
4:
z_z<b hFm/1JDyL.{AbPS#I1s4#c}(Z
R|j%/(>3aN4rvC59g3L.zox85~ oC0@%/Vgx|*uW>Nd!r(GA	uEe
&=gY$k'tccMs)dM#Z%~A2TUxANRK< xQy4F70h-1c;$w2y_
nnUZ[5Sr2P3J(^^gg{[pia]\L~%q=./9i`KWf;-2G)K|?WS
+(oz-L({VW-w4*jh%qIg'm{|CpWNk_;tZhm9pV,-}kJ?8.jA +Q4kt?\kLxJf$^;H^=sY2!>{P/v-F~JA] P5D_,a#|&as8z]oAjMu2$gW,:9=f1`k!FD;cn6i-Kx{)AIcSXB*E?{aHQ~\=W_%!G*<@tcp;#ST4C
L9BwZNn7Ed`BZj(UKv*mBpfDr/AW2 anYODBA#.zy9
alK
;uDe;}r%NWD*qz.>[+$)?/h0eJ/fuzo*CSK8yJr~U(h&_Y,q&%,Dsy7Zy3$ejG`M_)#|)nc.??-B"P}z8v6,0p.k`4a?4:TvUDZl?y*'E^:uqjK+	R=6-)Av1i^"2=y"=CAPXwR}\'Pk&Z8R(CH>&9e;xHb`?QT7%xdo.@t]XH]FlC ]AgDN[m`7bapmGkS#	O,2f9w,]EnKBG:I+OPz_o=k)s[$P"fa!sfPK5eR)c(Z.+w0Ij36Wxy/zZrd4yY(<r)5-19M@_dbhQK$p5k=4aq=dFa<5DHbN@z-8|a&ex(pH\{i`~-7v[5w%\_)In{#@\T@moG@31$g>W\?aL2LXX?$o}yr8`7T
@2aqRMc%>0cH~V\^n8#d,_rt_P)\6TM2#/R	0LI[fwn90KK>HUt"A8g'}~I1#.\~LAE6c+aj~]l_&UFq&I;{W	rJtJd#E9s-]a%7\Wmt'OBko%F^M`QAp;Osxs{mUU;cSOEZGN(d[=55D=1am3Ez6<<VH&`\'eH2qylX	>/'"znawD*VEeyJ&3BJt5Fy.x0zT#l\/}
gj_|M](j~2ZOPFYJHz.`b?iZ=3'O5z<CT~ugB9kzC!F4EX'	?FS>nK)4zePtOfjw? EK^dQ7QyUW;14ygIW2/6UvlKevcjjV:I4i/0Yg\^KFWHQ!
P0-,z .Nr#n~.cDvQUn}B330[V}Ca=sAdZ-,_v%
r`Coa_qSYQg,^C:;QRwW1-rxX=p@6 0,,ZX<#&P9mM\YSpNP)\d6>.x:P$Sw!^E:&XpoE*'BPyCyo,EXv0Rgf;T5oI0x~W*'oJ!'L[.LMuOGfzkEoG<T:qdsR29'UFX0-uxap^5.Z}p$$vO [fjj[}WQxzp_`$6`r@Ir^?5s;Q3meGIBLFU#H5}Z+#@bXwsv*N*s6E+~L8@3"',!$Bp'.l'zl5,Fqb819H.kWOZ4)m/k6
~}MN
C)lPa+C{#y#A4lN,ahlY1dq1e_2Fh7^FqaqL?0xg*1xc4fmZuhf{01)bvp_Z>%M?f;PW?}0?hlM1a;!2H[Gyp[L%$ZH3|k8L>Ve$0	U`Bmp$E+;qJ1
LZQQ6Wpo72vB9<0EcUcYPDB!}TQ)Z#\PVV1\G%;4j:b'cEovoJle;U0F~wPBI
x q~L1KbUW(gl=Lbb))D&xZ:fg\"{I%2PF)6,e=25CR
_TL@b06$
}7TVq>B''~E]F;mo9'jP*aJmb:aJ\zZjm6j_<^MwB._x)"^2.>$wpC/7g>a'K9
?3B8fwPg2tnTK6J6MOJ\17^3Vj!W%3>h+qY1p{Ma?.g|],0b*^^$,3DGo)wdHN*C$9
v!oy	G9J>SyE0CJQ|^3	QL|U*-,_vtPSmQ@\w~OZ@7?1jdez2L{P,(<NUwZc4Vbe8j$K2N\7K(HL?x!DS5k$NyIqz|wHa\8SS!SA2$lNsnj!xY&>aa8FEGmv'iriIqT9-)PsP !$de_')C(<W<m
hS6A;hiuNO;:YrXys9)ID[hwD6ARIRP([roRl>c YX-q@:RRam-e>J.nc7X7_Tr}W<3[jQfHn|.Y8F_;"\X,hEs}lUxAOu9j>55=izS:>le}5,N1&km7%]qh_h[]ELGr<,aasL[vd<=a"N*pBsv?!"`j|9V]^Z6bE@
pR99TR}^wWvE]G	g	Dq]VSIFt*#yC3QxxBy(t
jN<U>YoJs*8{	$Yn`L_&!}Gw^5qoCG+<3**oU[4*N,s8s_,,UqvG95,L)Qp#j@ggZQ!6+@F@x>@J')OJq6P,q/e(&h?GBZDf\~J/tss5<QBSe~+0qoPr$l{)K]"eO+^Ts
Sx8R"~U>W0N+`@:!PS=k6;O(?~%7>6qXHxn*E&[lyIp+&{>RACp Fh)PVUHHA%7rrw>G]:5TNz&4<Gvk$Qkj?2_zb$51_Q8qq;pYG*diudoRQ}CA My
6zy*W-`@vo(maaZ$dz9MWS@yTU0"X-"_.}K?&~SL'L!^kh,z*6&\Om9Xtyjo<q/O
Y,Ue]wpV](_S7UH_OHma8:~N>8X$:}m#&_\Mo+vu=2xlG*$,SG/Jp\jUp7hDkAm
lXuQ_BIlFjUZpC9p+5't2<vLSIJH^av(mbf	&X@y(5,EkA19%|iA6Cr,}9+'VQRrx|'G3;"#*K}(CS`jitxecf-2x?[Tt9MP}liray#d%olv\cVos"_
-j,n4:u%Z6%o?|WX]Y'6ehR`}>O)HbiuH\m#;O	Jr8z^WghxT\p:-O+@03^h`jy9_Q!W{r[8~wif1XD35:5'B7EiL a.#LCYV%{[
	UY^`;R$@W*p.]Fcnr$Ixe]}j+~,-FKA]~Px@&7Tkcv6eDxe\'s@2nGTa:'@+4G@p-8*^x:*K_xS$42sH>u8vJZ43
*mjz-@+accm}a63Zi7BN{_52kInf$_|6Q[gi/L WS.GMH|bK#mB,wsAip-4dJOd9!A
Y1)W_msyY
V0ft~[^3Yr&=gZ	v'Mv#_?&*#s"Eb!=$y.{BD$VJy^(#L5ykx:l<Fnl"4BBKP$d7'%oF]~xxidYQ%H-{*|peib43FGL=D'3J-~&]$3}5v7-i=^;Y&0St,[Xe#yXJUZIi70~mp[?}0f0iI%1#\Bw_
]0/V+?8{Wk<'Yr0\qp0H4"ydQS/=g7<ysQ2fy[AftJ/37oQ'R]v]2'gK`3]{ZC=|=NiaK_}bxz~%y*@bp8vY+fme/N)5nfF2anlaMjD;&)N`Hy@)^F{]<NBov9LS/4y^z5XKzjqa5BR= {Y&
~JT;><dj/9>g!]8/$|i	M<qWtd|cw{3avu
.,vAWV[N1Lsz>[UZ39iPulJ:QxCyY,cd|RnE19R\)=Arm\*kG80f.P-wuRZT)+I/Ma?^z$bA`6G_raz!0g[rl-w_|onXh >0`bjG/VkK<%>h|y8]2c$!hf]lUx.`De^:'^I7KlTk0={@nzl6Asl<U*Hlj9Se,Aj.+c?zp7&4A>J2<I\$a\5mvcV&w%|6/!Bl~yS494)sq4_@3vam%8nH~|23|ZU{z^_{/9Q.4UD'Rk*ol-|5"N'9-ziQ,[#hC?18](W0ZXM:hDt-f%F"3_.[0C$TG'HO1Q(ONrrf2AoOS&",cz#\74jrt"pcKFo	(+gqt_;'Kxg	#Pw1>@1Q0z)eAdSBcJp Wxbpd^n3~lk2\YL(<vVRGF|qa:k1N7XXr`_f<to[;C1d!lMj&,rnY,|RLrg7"]7m!qdNH|lP_yzP@sW-w7[]\>@No~;5s/DJjVHT:8*%[*I|Y%s0$PBCOe=
I#avg)hTFP(X7|0qDY&k43yYHoqqndtaZ{$uBgL	 &6RAyn5+ _M=iSwPr0gHdayp{;4Y@THp\4):PQig wFWjU!BcCe)Y(*Gk*EAkuJ	mJ2,Ji%Fp;`j|O	X Q%q03V.~ii	>@H<QwNO?R@	#K+ECO?]LC$uKX0l
dNKE}$zd-/Ze=g;7>]$~Zv@{&`<+p\*ZBrL22\GJnBckeq^l{q3hhamw+o"Av([Zd`;'+uvNwj:U^ABsW{;,-2cbE-K.c__?7%v3@TEEy[P2Lm{Ii^BJZ;L$m<,}O)YGj<Xjy}-xi0v-3GBfBl>\2wZY5euet+N[8kD%s;5;sX 4rd}_@g+@|Kl$^zcqqX;6`Q9=)>};/pDa.F3hI!fjiE5f{pSk^U@s
wdqs:E$-FKhiAt)pA<%|Q]%I4.OYH6Ok4z*?)hirS|UP_'X!(,u#k:CT\K)1U[bQ1=VCUtVIiynW|CnyGCR,zei%11nSdCD0ql'|:Be?V7TjR@)%&"C[xpF<8@[IW
5BoX7;vVzocEB@l/&}-GdJ|tFI0BSah:;U2L&CyZ*={J!K^3uA=IS{?&q0h)`d]Xvc od	|vhI ":S
5\K#r!t&klZw#NmQe5jfUqI*XTpsO1D|
xy*x^4e<H{x)C/qY>>Vh9Z4
Qyjc]H6|<d*H9-&?bhJ5+yeb1+2TK/#]TD]OS:P
$Vd_@3IdvX!~IsU:c_>71fCmx`>jmG'|ZB<Yb"B4,w4*Bs-
V	lbE\``)-ct^etYS	9pt>Adjxl^`e/a6$os"U_fk+GwS"3` yXDvl&`(AHqQW&6{{||cF~Ir&1A]:kTM\+
w=ll3g6Yh&[lV9Qz)HhTP>l#+O )5825{&P[gs`k^A	O6OG%UjA =/OoW0}8clI[&Y0x3j3W#C!=aI8CDbz\|z9sx7mL/]b>{zn{(w=|"?dP.Ja?	7YA4(1*z9jW7$u2GSK3Hq<zm)Z}Y=NcqAnp@M9vFM9^Pw?oL9h
J>}Y_oA!y_	h?z-;dI7=?)7S'($L$xjvU!q^C"l1`\BP8T
ob`B9D,#%CKP7x"}{JdcNaXf6H6tk2J]<y:IPzBMg-!zC
dFa]Hm30KB)ppW-eaHU&xPdZ],<PRrzIV|iCJ*XQxpYIXI}|Nc,.HDs0$%axT7ErjS`af^:XTX%e)!T&}{*gfBOhaf(hi5lQxgj\I]?hEqJO?XRh1[N+yU2j@+)xs1G-|s5An;$Y^Ya`~nN1p
>a|OM9#328!E6o$`	3-u|toR3O"e
iAG(HO<qEv"iC$\QWO9!p@z6y~[N@O,leA%ZqN'^\Y#=S-Z35!(. (|4MX-wK+NY7N%nX,+[:l3J*;wY}*Y33'H/Vhb_JudvRF`xtwjuf&$W|IVL Y400Debu`}wDgN W:3t4d8|8j`SSF*{Hy:{	A#RNmFPaNdHy'N:kYd+NfT=y[LWduIH6*tR6*omsjPQrmZ-6&I@S\QEUqt
11E+MYrynl}J{]D<bNfjh=iZbF%sw"^1"
jdp(m5l[{ILx]za#?@0Go\j:;R3x3S}lsw-+"-%I7fuAW}Zqsxi?PrUDiy-	0kc'}oLnPkk''@A-j>!~ayQq@=Itfe~)N+@LdC|O)'JlLGUJ}!^vo(.30JAoWd}/NYKu&*ksx07ck4Pt=V57@qX0j==iYT,8?Bxq/JCGw^RNP|ie	fjeB@J@YEdAT!M'3A1.VaP[Db8n/hkxEhC!`,EGuv;9,wPX``HjZvo4t8kDEu|Ek2oOk:m&Nz@}b:Wh?xLVwy4Ob:j;`) l6Wu]YZU,R/m$:xTv.W(D&:I/H^gd@u_K$wh/$)C@Nf~[4x{.`aOpNu\Ba+l0qhTw)}sHsctEEtjwZ_)~-j
n_2a.GVa)xS#lc&.,r%SLUNNvN^t@Lp.a%LxC\~t$1H8}6(,qJy/TFo=;!!X2@qlLq6c/R3hQ2voiCl+
M<&=()/s EfEcHQcyWXMuK&fe!OqO9LU?|wH(e2jB1h42<&7:hP=6@/M/q>[$GVh.}MIe((Bs@xN,x+(9UBL&Rh]\R20A{"ql({oAx4)M!W0L;M_C\}I*:aC!=t3
*U3!!(QoC]`XyY"kgmCXt;uG]p2R4J&Yn\JgP/K[@.~!Bsv40):l3P6mxq,d^W"C6XJj::,'nkCao;QD4rxY@;	2+4K288_~zkiEkV{~4Kcm<b1FpXLjouA$2gE^8'6t~dX+a))WR
.<uUvfu/O_sp'!JDJj[hXSHo(N[$3){~.zh/sKZY!>)fey'mBB{dX'2i8&29cRDKuP(B97%n#&}"CH&W7R8$V_dFCQc50BiCwzH%{Ya%s{s~4[^KU5B+Gh*AB.H!B=~i|jEe3Kns0[i=+gI%l{4TrkPU)oyRQ}yjbFKt{eN5A&.$7UQ[KS >[z:^$3DvFTp<U	UJY_ZCl6K*h7`3>vyq\ST=-)=ax$ijf!@s!-eu1V4k.k/`h^bOpNK%_>FA2+m)m9ZVB:>Mh.#|"3ru$G]x3t"u|%`0>rAs\+ebD;ubu8R%K{7H|bsNJ0laR<2%STBD0xy::Tt-D28muPQ	1R#gy)U2jGR&9;E'T/.f_H2^p8fY<eMTT9o|ybV7m6^q@QPVWlpTz5\6/58`4CHK!jksU{@\L`^W*i>H.n2/*Oh@<I:whDI`(+K~5(WNvm60<Vgxz/,U44n0;W[Oh)r'prkap\{$5Qn/T|F8'x#;c,5&IG@Pc\;@z[ Jj4@{V8!e#8mtMs:C>Q5s H7rH
uu	D;pkn>4wGxULg}{x,aa"&Dm9=<W"@ZTPg#u)Lhb6Wb*ik$QG$&h'}gH+P[\s!b1yF!u^x(stIk
+;E+zu3	1}-zzW	n5I(1aUG{/[QXceW3
z+4Vgtr=VXs@#AQmd|GQ$$.)!.t+z LI'$GFyF6|gt4n
sNDW<U<]dm>F-/|q*USb?gU,+*#T\I)A%WF	dupKK;Gh{x6qc"19QZtD,oBQ[|b
Y"sw
mz	D0YI46<n?B+:BoZmv|zrK[8VF;$|I@a6:EAuc	[y^3lgNki2~J-'v<	op.X%oNRmA{6/#o#fZ]U''p\4zUCbo!3p[OQ22>!r*WNtT/ Ei-h\vh4l/B:;"[4Zb1`Mtow2/4?"zX(zZx4q?]U2ZhOO{8(&?Nr|,]/d^Au_|t=)Eu(d<'-vXEN
^;Y;J^!-!1{Gem}I|uuJK\T]2Y_7b~
o},8!BIp,"k7RT MXETMiL7UYOGj8FJ^(|YdMUnF
;="P<7*>d=6 Q/5!S~pdy$<}9d8`WR/7ctOm]R:dQKmuqn{?_#xN6/0{U{'EJ~	xiB72|qC!9O3>*$3bSY[#'TJ8Q"s3 m@&*CA2:,_tx=]h->)zdIC`!C{N-*m*3$D_8UGgX)IJ.7f3@v	CliivqFoZ!;7_q!1fCI?X~qW>*F!Q%H?nMx/5!A8S
?_z^4'1iM~fO`vFTDp6{)~.N%ze!OnwrAMFPy	dw@gDnmhT0&0p;YCoKj%Mj:^n-}vLE{\*KCEB7JmC>=E&yEtwYf_zIe\$H)3AeXj&c92n<Hu~ETZ5)SC:x{2hC-_ams`/:OoDR$1HiGh74`P*H&v%pYQu3gqg54_Kw2Spu?]M~sW7h`sdWa0VX88gi}VRc#/G<04mt#&2c{3wdM6H>RjGEejWQ=#hrN2uisu)a\2N)Lz2];65;nYFQT<u,x88fL0FEHW`}>Ldu`f@eAg\0DG7,}K,A?vY+dy*'399uq.EGG'etZLyCc|qfdzDw2!Lw75E4`bja
Hsv$0$.Xc[2R||(
V(DZ@1RoAxbJvJ	'.K*D+'//<}E)#i9gW$tTV+ISr_^ctlvL\5~1kn!N*3XTg2}+8vx@e3?m~, d2MijXa1v+qcm*um[/ec)az=4xIkVwKQV5<]HdH/<8wL\?Zq6C_W"h=V&kd~#Di$ueN>(9zeO2b#di\\&+4.[bfq=5tPDH !h9EiTl5}7J\mhpGH:rUi18dww?]'1sI?S*Z=25"~A0#,XV.4Acoa""@AO5Y=A-usP;xq<h$a+nexw6(~LVfXjS<QkO)?CGO?	W@@`Dk!Q^i\B[yozj87ZCv}YZv.p<*7-8Ek8~53E#EWRSVaqQ{'Rr6`zz~n6GH';]-NVte1i5d}X,!K(ty.hs\WGxXPr^IjDuhIfYE^+^9z(D6/6*Jr%@O*\OpP,+%=\*aP_YK\4o~<E%-{/%;"##G1P mu3yY	@f4Pz?;tV,K`y@zcb'	}{faOsu;x\5.Z[P../4yh-kr0t0%Z@~@Z_TVHH<yBm-cS\v(Np}e+m3?c4Z,k)Bba+nH[Rd'7g45-M4\PV<N*nh%q8-BV\||2[FgZQ_MOW3Nm?ZR565=:?Wr6!p1b6o6kE]pNQ^,kgeMDe!!nzJvGJhmy	3
;R>~=g/n~Y1$b/{.FvhH}9$>F\/,15>:FB3`LH\.P!:s-_x
\&AVX2?X_e56E/&`ZnETf|b`ZVEFhe?'R@]yI|1C|I?"uZQxaitEa!P,lahnA?@S$:42*Nc3cDKB|gl5N'*c61W{>^>.WAf,o8Q]]d5iYhiNA/y3IjFL|AE|qDG$\R
]oUI+P[RajbQGeb ,C/0/"$P~-kzMA\s|;_U6Oq\p!kk-A]y%W7+_
!X@{is#@SY3''6G%*uh2~m2
5{CLhw?m$_:THR2An%-^`,i`gPPYtD#s+x?t.myW	iN_[	z`)
k?q^W%7b#+S,D5j;dX<ZpH>u=B70:B	a[-]4}Gl~7OqdJF/T,@BST,K<%<clYi05QK8~w%OqkvGkF.snE|<7RZq{c~"^	
vqIr	80QM=_iy:b{7ji=w?3	DrLNhlf{I-ss}Et6hGF=<+uc5PvAhJHKSQ'`}!3qV56C00}x=G/RnzBE?1~+[*:1xTR"Xm+~yI_W)DlJ0.w$R~D;8xyGS%	-0y	:%=LHr43B>y&nBQ%5' |0%QfY	_<!R7m0)ODI?b;kQ\(\m97 UpdBI)Y?Y6Zax4qv@m#\>}?	>Y/]Vvn~GOHl:c
s@$:/k&\KQ@[Z|7'@q#F,~76$h~r
 Q	v-i(Q\xG4>AYyeW)vGWu/L06*hmp39^z}D3;2,^GIbv2nWD.kWTJ@-'OMPObIeKYvP_B06ndwP/5wl];54NJyI>(G:U!*Y(P/VIYJNUq%V>i!w,`/Vyon"_S2I+bc,2Pt,?3*6^+T~8|la<j^;mSKn6rM_@Z_1;etL_{P(\2|ka@o"ugNE|$Sd(NDjBb<I>`[yz\Q"outo\5e3'gZp.L#hx5TBzmW*QAB\`${7;@GB.49e*+
) BCpo	%EC%K1/5lH5	YRyWxc-kSjYugadU0wtZVz/mk-8{aL)r<c_SSr`L|P^{'blX<HQ:ReG?Q*\r~PX}IP=)!v/]#99Uv^6?Ytd.[2l%eSgn=\G=fT'Kjp/*OxGL@T3^!2oK>@2=`my/`7)Dd9a1S!!v9Xnm\Ex53dd~Nmv@53(tySqWm\g*^Xh.N(`@Oe@4a%,cjb/bQ9ILz@^Io@\lvZh&ivpQ<>:}HI_atGL'XLNLC"1GL;\	-L5F/2ExyK9\N0X($tFATQO3a/BEB[Oj}/rYXI688oLGfiGUYbc $)t-x#V}\6#ROptrCK Z2g?@z0X/r,]KG	Vw|RuuwGO3<M{T`.x'A\qti7skMab#qD2=J=io&tWBf:s"m( l	X3
<vZI.d7bKIEJX&O6TVjc9+K8mYF"97U'2@*i zphgU2uvfCm7N(n^cqpX`Qq66
"Uq$$A86_Td$-.n-".MQLli@6in`	5T MS~XptF?/;ofay"Nl9g7<Obw~*.ctx}^9D1X$u&rf9;[/19$E r~7<T*]lT?
V*lZEAIbEm
'B}IMt"E2)/3SIVA}`J}<?L6qsD
Z:7z__:@Pge[2"<G;3W9Gz*W|DqW"4 ]Gg0uPjN|e? ]zMk(gz=W+#$
."UB6,MS|)S;c3,RR?k0&pZrkZqVdq-6(5&RC?{&"P{c
	dhH&x(NG\"a/d~Gzf
A{.7D'-$S4N^^x]qO9]NcT5m47B)7fTF&kJ(Z=fmZ&7>DR9{p2VGoE	=w)V+0AH7z2sg!tqsVI}of?\'-/b^Ga!\}*(.f !vdWFWK2|M)[Z^dC]UEm_\%I?0p1Hi!q*~Ke'IO*OW'#161S{ er&@GvWsVF@f1;Zh5j~b;O.Z2}@qW:3JFhpht-Ry~BwYw5~r(Sn/T[W<G|8^)s"v)g^ILG[Sz|?t$g/{5Cf'/}t[>KHoFZo2olAN[7%1^wi>uQ}"9Ip5=jfVC4HI5bu'z't_}6S!6:l5o3"0<_1XZ6uVNaEo0oki6HN'UwG7k"/Ux+S}A"$CF-Q+k6^>zMz+z2-g}mMYMTU^rmvZe/h,\}uS2Ldq2*_({\"PY8,#Zwm	x1L#6<G=J-La2!t_Y7f\WL.ZNNe'x\%L;7jK+Y F&~P/*1cpCs\G,L	()b0Hqu!(!mt }EbbY[;HNv1ZZ[yZ%$;j<%{NWF,oyi:>Q3QNH^@:sU6hW~1k@u6K2{'1v`vM_Z/(g
(Jh_-\'*.7590QS3m'1b\uHYji|="hk&2K'h8b9sz"
/8]!"VziF.~:nT{<5Z$u.'KWeU/K3G|rg]J<yp6@u{(*{eeu(i[Yme
-gc~QjvRF"7NtS0]S)j_bZWbXXR5o5!`:$2IiRj	, "S)n><*',wk/tngi1DP00@!M-[rrelirMD+\,Y]K~(+ld|RY4g1c
t/.Jrmg;?X[L0oI4Q(vE?cNF]}#c=:0[AJX24]@]lJ<fM"3fJn/rKN/smZ{Gh0qC)_",C\`+U,UU!4s:C7nAxut>s:XeMDnx>f<rtT"tu?"$]F-rwsPRL]{%l)
OP+9\YSI;x}LK{_oBSU8>,l"yk`h-Y5oysV&Um0wEl96`Ax][-`]<:rdeIz+2# (J}<jHv\e##%k<L17)G%Sy?TA'6rK?KHppI\NG8d@bd@f?$;-jP?<)MOW22dIb4,S<sz5o/Zx)	 qq:zA.#w^5LUOV&Qld1htM?pS3/|~@V]BkD6qi{`IC2?,[>%"Z>-1=F@41bH#GR2g)ZUT-ap0	J,~TN>ckO\lk)^R?k
Cs[3L~M}.$Px;3X!/rqL~s!<?wMH!q;
+@w^#mnM)~k9Z(H~y<SfYNjSu|ZZ@A}"y\6nRG.^Y=R%<skM
:6L~BcaR+zK.WHl-%!vC]i;nmym[1eM-4`f!:<VO^Q/.<Q]}cVAl`$Uo*W,w@5t"O!	rj)`[}a+gy+GbO%S0}<&81%;B. }*$[eM-mV;@vvU5K2I`^c_~VXk8	:K
tKdbk ':Q6_VyI/|?#G	-Uqv
uYFp
CW\=0
z)V`^A?K^tLzhI.&!l-&01Ur$<z|E~)Br28H|bOc?d\M]]3[,nkr6kKz*tpLb#k
i*fe<q"Ppk[29oG|	L~Tf$E};du,w$DG'k~X<C*X2mQr)89K&^rOuwGk960>FgATJF=5c6YZv):Jt%0wm"3@k?K|R}P9T<??]7L3)dW4dd5;^`+&9PRF3wXqXcG`qLHTOMSlYo}Zs1=#5aUv*}cS;Togs6WCs<ET80]U{]inN`KI/lkms
B>
D5pJoRR$x#u2|(V$amF_\i4CNSW5&">b e<''?#/_.gV(F4O	fFd*T*W[7ob&|U^d38Gq[<M$^,\BR(MBR	,&aLKM Ac'.Gj0
	 ^4U(fp#f~K-k5!X5mTsF:oEbF|rIX1X]26$6Q4lW$P0PlDj&j:2n,}Cr>a'MYo<
	"B.O{S`*~r6g@$K2h:GGf Yoq$9B@kgzw1I3&wXult%'=4wgbsn*NVCPXe>35&_5)*GBo>+j+2Ctc{&;6xgwR%}Qos}[^_hx',Pdn["?n\?TU>qgmjq{S`	2}1J`ush1=\-,_=xpSY ,/5 jci' I<y|SX..E`*}.Tjqg)(:xMzIrSjnxRU65NOQj]')F[W  ]I.<_BW,J+\<=LvJG!A{nJFMZdW(h
Rci4u,Z{h|/5WGs&{A%(+v<*qFl@{R-{E(|&,5g~W8]!L `\`s|Ch&%(s$EzG'Qd>p[!pRRZjY]Z&;Lr&/BoUXj)YQ"kG;2/
8Q	`e({$$hAd`dBq/~9yuC<i#)/d8/.&TR/\c:>yv(%TWI$L0S+lg:rM)4$9HOGn44{\`JTVYoA),;M?La1e\K;}Gn<GNS1<D9f#0rx{8pnlK:g0ByjX>+D`].f J!MV}HMfzjt{V
RU8(1Zx/h*V*su@|TDS+t!x00e"\WMm0`.3D}.8H@]*4{'qtTc9KLrt0B~,bi'4b}, X} l`NLEJ;-5q@o*H/-}5?koClY(@h7HZnsv8^\^,9@Q(|~Qdq";})+F(%Dwa-6n=8%d.uqtO	[
^xyk6e2T;
[mgR{\r[15>jKdr<_jmi0Vt:LmXeXj;cu/dNEWJ0Z7bmw!c3v}-h8V D#lZ,(n$c4*k_lH$i9Lu1(3iBs_8=D_x(1j6I50jwV_7?lsJnjqS:J;d3AmJS;yjB }_h)iHYess@C0=){A9,[oeQM4DW	@
7v$I4oV-gI]H%G~p0(FP1~}sRqVt?J]>uvJ:cBuzst!|RyO2$'F>'/%%DP:{xwpviy!qRA#:KA=Pe91	%!%utWvJlcN;<jLk;d|L&NmV07J1dx":s`x8*ZWv^d>w+hntcwlrWlDbz/0:_JYm
t$dP"B]>*t:_u}sw=[n5Wk)N@1/V?FpLqGNu/)bkMIgp-%-tKi_x_"UXP
Wy8zcCwtCLg($?:4)Oj<#!pbEt"8m*!bob_Vtg+uQRti3y:DOsbXz~#U$&QLl	i)kskW	'[/67\@D<K>+$[{'}mO({Y0D&$+'C:[/&BuOHM"d)Nn|OMH*CiY^FPs	zxb)ViWt5F)#)ONU0@HYt3	jkoU)9t{'<pU2PE(t/^W3)pw//85