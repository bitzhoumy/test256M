-k}d\e?$D8+;k8DnKz<8
1@1Ee`Lc'ehwk86VviM_KQ9o,B`-/%SR;zMI7yA w1>pP{TDJ7e;2nZ'Y5XZIe8!mc7DJ3kT7<vZ%D#C>#,?2<@XVYb+3osMM"hq`AS3>*P_{7 >G2\y=?1Ocs0Ea&nm) y:;G{$ASEg'I\5}we0\B|\a&9r"
c/y"e'5li3h3IoA1UP?,lKG^^mes&6V}XW>$" :V^2D rw/E&<$
7yqFE/\nsrGz)'}d*D$UC!A-[&29Ek&=5Sds"'x,[NRa>=Ju(K4^OYy
fJ"/QL8Y.ChTBy2gK}C^ob2W|^iP&g\ZX 1TE3O|;^\~eK"4FU[%7;U3s{)Bi`5cF	^Im\!V?'R^:nNPJ6IPBk7m*wVKs3"o&eAF(%^] V(%P1.nVSS5\|$`LH?vtYL@rB!PKv*}tN)^&	'pq#x+ZK,,04bT+?a~m=IT0Eb_WxL@_2`o"En,Kd`)B)gajs)Mjt=Mj&gLwj.}3)Q)?a[Zfpv5ISsvMcup(0/7><mAEcH)	N,?_FySZqQVrHc>#Y,Am0bBV{4YdO+&wHzClxScV*}'`H+6se?2";B*S5.n(MuAPoT(.\>9Z4s}"&%	E(IPSu.9Q$Y3>2v+w"0rD=ys9/ZS$9~KL@97icv@"tz:|6gx=<%\6b6/"O	n=Q3wSmcp*w08IgZ||vo7&\?g/-*u[z>^0E{:0.qOW)H[ap^sd#j\	p`LQ?J\YC}J<+Eg%	{:K.[TgfFRH72gRC*\0?2G=|%G	VP^fDdanIW,iJouTd)
UJej?qLI/ +\x&fP*`&N4uivt5":Io!=B kAC$kA+Xv2:
t/<{gKu2Z1<lNJ%cp!P)#no,:'RV(!}>1*!Y5d8~3fH:)$"| /mb*s\CxE-z0i`iR1@T~D&[,Iu)UD<?vQ1K!Ie71b'+|lZ'6|	UE=[aB$2)*wnxnU`fS#[qO#Ic6	-Ql-SXWEbxO.zw3
lHHuZV{4v.}Z7"UoH9xe%`Zwx"#,7EsFM<jbE27}-+iI(Lj".	czX=S_
'iMY!.r}`px|6#NFXdJ8Q0`cq~f$ij;lyOm~;1X97gOQC7@C%. q{<`.W1[4h-"!%p}dHeO#Jh#4:AHCb9l<[oh:OAle@-Wh=33-n0PHnV[M.+@JzNO_@|3=]wM`}brFJ?,da0I'ec.e7(.y'*==	 l17\YHTbz^vESk@=g:T%VMcjV~v5Cd+t$Yo;V(.C\5gL\/Kk9^|yP%`hulJYJ0LV+^px}i[~diZ!5d"GpjNG'\N:	fLz7+i(z4#LMiEW0LJJkr+"#.W\6;hF.'bit1.u1OL@\_O~	3_j&Qxt~:1]E^dq-K;{Ki/`;sop2'Ax-gYFT2q&sTsWeb}%~9bvPOPMnSS&LCL!Sz/-21{#iE6YWw!16-iK	FO&tO+UUk}UI3-v7.S6K
a)C^lVlY>]b|FCX0zh+M.:+VBN?YfvP!|3~b>S-v%UN>T?IJ\c*_>1tTCvmGG'\yM%=0[:9Zy2T2wN[wILVu^c.ruc|A'^>|a+;11(6lmq7%ux-$[gqMV*z^d7d_D,jo[:45__W@cYJ;P\Y{?y=^	L>UZ71t-sLQm^ 
_-^;j@=4ozJ6ezK@Av7|Y w:Y*iX5:QWa{e9^hjL(h8$Ku o&r;lxS z^K.YS]ijcZO$M1Hf<<=n<_Q/*0Q6,L)O&Vqiop..uX_F37FpV1CJ_C2[QY4vL	h{.Vz>E"M~gvOA?Lpyt9Gbc#7@#Ud]>3G=1i#;	3^/dw|!YU=?$]}#wrAy59`kAaAD3GL1.+ux|*&ti*=poc{yWt^]W@O_)ZwUb'RLa.TLi	JV5KDW..y
1w4yE9Y@~g&8nk\8lAM.L<nA]&oeUw|&K .pH#9/&gxsVm&|x>aHztK+i2%+bA:thsaV{!4X+i#0OHYtogr1${WoJGX86;SPt\RDPeB"rT
--h ]O	3M8t19O\ZN|z\L_PT&kI9qG(o&"+$3t.n6s`Yp@u!$JE+Vu95&XzpNyVf|?8N7JCevc2e/}t{k0W[*rvkz$@BqiU$!/.C,-,5KcKCK*F`DH.~Ez*JFRu^(9[wm0?Q(rq1/3c,wXr%NB|Nuo/?69AIpXec^S7J(#Cg*^2':'cpo46d]p2vIOK?[I_~Z.2I_K&/h6n:_XJa{NJpP|4#OKJ9+mP{eO[\.a>1?L:`*@-ll x?umfPVR,,/gp7#?f62,O1.`>IOC|^Ex)n:>uJrU]<bNcRsiF	}h_-625t;	+)v^Tnk0}1H~W3V$zpWbw(NR|n++m#Y%Dd`X^ezGIr=^S"!ZnNlm*a	b.\eO}gks\Jw9&a@*,T&^_b&|Omb'Jk.c9!14"4#.:It|9J2#kRS9BYVD@
n \NKN9:%<_LE7T;m'Q_N']XA#E_$L[
Z77p3Yg_\K"4AN6KoML1nq! z@{V%a#,	&W7?H4nKXZe.}GPx[~X&iwvI%6zA/0)yF-r]ZW\9]Kj##PjIi0=DPdcg_*t[d1%ZijAAok0ZAK&?
$fK24zOGd ,Ge/0w?9|JD2!*fBV'-;	]'Ko'y'bo\%I3se''W4!B'hYMgu@P{lk7"?=V0vXBf{omF_G>v:(=G{x-xe-75vyp%q8 ],Dw`9afE+.q|X'	6Q0P|m*%x4!%;gKayzqP[
)f&|fai@E4w
~B?[1'(-\UuPA.MCJI|=o#MUq!&^<eLciq<k3iLlz?.Gq0/\w	dgqFsXzP.BZ*K6j:'7s#	`8bq'gEQO/&yGqB\M>JO*S{rJ;!Sim8zy;kON$qAKp7TK,RNa"7xtr/CIi<A5-h2x{@?v. ba"q5%&!0N=:X3KD['+WMRIMzZUJzo8woouZIh&AE~Ddf0C&;K8,)nk]b@Oi2i e9X^hrd}?SKSs%7lhS'9<S5+mBSF~B_:&A}P/M5@o1^8dv.U&rR'@Up-%{[Kpis#"j4]446'$fs:uQQNZOjb4FavtkYavjp:<6]J9!sEVh3!70"19pO]XGC q
_?;4+s@q?>f\0gCt:y>u:Y>,EJj!*)<y(ig<|@2#~
lY0wM=?qdlb):9K(;XFB+#+TgYA@x_QCry3}[z."D^KNu!';pjA)*d,%{ j%SA>!(#J[fqYq~hanzo-'&HKy`b}7XGzV+>;:Ic@~xn|<Mk#HL(+)HIKN@7jqSrjuUB#@v'qN/FH:;mf:7q*'A_e/$VFYC^ MM7R+~oFbXSkB/;bpgx{SK"	]>T<$Tzsq'r6m-^xJI%=.u9DFg4}TCU^Cwg>X##B;?S(Y([EB~&A)7X0Xx}&oe
,]VGL0O7(q\Z8K|$B&<3^{g/7D?d$##6Dpq?>}9--
d<Lz<Ia^q-<9"Vxf@	Sr@:,Ely7.RW}]P`{5>Tl'2?>igc-YMW8r,$|#H@x
nsfHs/z|K5^(d/VFq4YY=[BE2wu|0Gx<($5?UG2!rzuUFI;|yc~R]1_Ii"Bw7E%5"kbaGXM~2f:}H[Y#BF0u&3A	%WL/jN	>
7#"V3=gSeQ	f`5WQ:`8\ONY3_b1"h4q69.x7aju`phZNcR;on>	b;m>Z+4(TdzfT
Qm-):=? lKf-|k6E:FyK
sCNi[GEw?+V^!l&?+umy%i<
MJWa"|9%*G;.	NgMJZ:@#*t