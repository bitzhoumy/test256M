|e$\OQj3>M z|WUZa[B'J
EJP*]T)#w^qlX-y.m<M$8HmO9u?_Gu5u=*6G,2 {(yBF:5AJUrbt.	jIr5+Z'|_kdN.RE*.pC=hoLEs^OS;/_J>O2-^p&F|WV1C}lG\K";;<zA%&6[Zve7v"pX""O,b6_wt__ 1_`+lIn"cf	Y!/1rW]dnz0.|mgFhvqA5u~_#D	Rlx/YA*6'aB}IGo
.</a?w+-;[%hVT+Auy4ix^h
zKSjxW)`vgh~(Nim\v?\?93qD/LuqprH8az	GKG]b7v:aU%*D_<!@NZ:;o.z4BK+'[QqHP'vQ+!)s{/dyaf ;;"+EJnHk3}wK@Q<aR9MRv"P+h<Nwtr/ji$8UD.CR<_cvV29cEn
yYA7EsKidqi'e/)>G&z*"4z\?,+YI~}-R:{_,ky"(^i&T#?#+O;~Y?mA8cyYgs07)<JlXWP)M<Ef5+I\Y`:/^);8K[P[mI;P(w/X"/mK-Z?@@6FHT5'P:ot^ixU#]>gd6.fF<U$x#<9\F;nr-K!tRYe`9h+'CCk_LYa?LBB+n$I%0x%CVll$vI<K(mJCR<ZRoSxm1GeveB/P2iA}
C>aLJ5%Z 5_aRJx6sn-z	6!dnlj95R`nU/Fh. -[^`he.NQ$"P6U2->H$NX|l3TOm3V[;nG9xw%X@esYl^nz)TD%3NZ&N9$!3V?/PNG&IT \WbsX+")~)'>E/GNeaNgK8$0BdKv80_nR8`uPElZEcPxX}&[mu(E#L[At}^Yq<6j'I5	s]bQK:.j</Y0&1C'cVk8
fD*7>re^'<yNV1Kq@C(6VmqB&NM;8[D,BQ3	d\x;tukIBF;1(PAVyT-wX$L+\$).[Y@=mOLw<z$NQ3!i]bGh72Pa_YXvsQfF<?o!!`uI3=rc{<869Hg2'~fmr7W826<)G
YOBZopHj?/C3Jd4<u)PsK;:eMYFa|!/zP?=%>H@kwa}9l8=Uj,uCxX
@&TFcA};8kG((5:jcv~u.3	t% x~*'.$Y_|}D7jrl1'7TANl"cJ>iIElK0sLWX>WambUlv=s_"59ToZL}"VL'|rQeI!Am6]B9*XZ/cs"qLUqo:0W9TJ0_elxP4Cg*Jp?Qb>M
Ms<:2
e,EiBs^AC2LbjUiU(S,p$us%}c`]|U x>K^wvt5&Xk5]sij@Ivmj,4R",JN75Kxt8Z>J-7~%G.jr0+grcT?1]-*;hfS:gU%rpUHr
gZj`&[74"S>_Y:U]][-q[&9U=|:GR;jG=AEO+gR\WZEK,hVlHJJc,<lEzTA&hz&:v)v &U}{W*^/}i|j7[O.pJY	."Af	GP&kw[,B1ar[&SKd^|FY`9V2z,WcpMt:<R7y+\o~h9Vo#QD[C:5KnZ	3PS(rv2oJ>]9WB d21VL!n\TH0tIgw_U(zl#ylKJi&j"fZJWK~L4~?>6dM%uzmnpwkpyg$Q;cK1O1dBO.-"$ZD#<8{	"u2#~ X\'RqC[</.W9EMNGd5ebz=pk{P<]"1!HQ"2,;F~	Za\,<w !JgtMB2p`k!A~Hu;}ExJ!-:7]*DiY5qt4`11";u;phpIX-GTI-pKXY=O!7LK2E[g5SGT{9c"Hmm"&7*#ktFPk2j'!QiifqQdD`{~,+8q0ti3HsM6TemwCXS<an\S0{	ZYu> (&wtQt4FYkG\AsbppvTuY#,X=oX+2[)3H7-'(NYqlZr>	q6$~~kTfF0Rw!vATrI\=WRoBM?b"
y|B`.A_bSr&'n<+o#l	`n$[rO>NQy` z<7Q:e@f+,`qfN`h(.7W2sv"IM{n08uH\m8]/s[&i`xK~bS
P!b@.W6Jx0gBGU&'yQSQQ"OufK4(XZYOi7\XVB`"uHemiJO>n_8]I}lg5iOm.Z+~eGwK0q!7pqkrx0+K"sH2.FhT1,.B(t.un1@@H[p"|	Y~fXUv{Z@2Joz5g3V.~A:@=Kfcqx7Pc`~H\HvuPMZ{J#]Y;^Bg^+wZJ3v>>v_=tQxv3tAcGDf&.oO2F%'9c){(4Cx6}W4QB1?e*[6orRR])'4}@_wTF;tr1gW%()ev_;K&rmegpku>SB|q)=$*Zg5[2Yg&el,U L`cv{XiOAN@B!zSKo.v'%&-yD.(rpW)R#6ES)XA(Lgz%`.uC|=IktzS"?92WtJ?6^e.(T=r^;fLc@N\F0U
fZ>h38"r*@IXG}Fc^1%K-)7JPT)7-wt&z-rk9V@b`meQ:}1
U0W8sV?qeVI99K]d(M2qW>aBV_Cy7o`MsgF;{{.pxo_g-J'{rg]=S=w	<bE7|UbL+.oGS?[,tH4_\f-1~frx')./&EPT:I2C*LkPtVn#4R}~-CADKw|Aw=|CCqm
`m3vI\-Cc]7{1,Gqyq 5$/pYJ/ ;`{Xg[V%Dgo	w>e,fkT=R>QL"efO/HVPHxTc8EI!6FvYV:Q8;;LbP5z%[GE`)vT<YhTo\.]C`9E(Y-c#C~n>CZA=.r._k	r0@PP.Y*MU|Hg8:_d*_.QX_7Q'K##d^,&2X6mr0mq\a]lNe!P{Za:o
cji?Ex;/uEZ*p7FO/1TE`\aa 9Mf/cP'm%msjT)0g~hVBJf9M[ik&(_AJlN!wM2@_YWQ7$`UHl)!<* O	3`'E=%	;33@ZTF7>HX9AOmr##Ew!&RZ^u(Ta-q2tjl;`jPm"}3Cx 1Qcf+"t(}7MOT$~j2S!.NpN}K"CF8SQ;52Yq3K6@?2x4/yl3_uNyY/,b/+?49/4U2`F
[|[:$ i[hJAkSTsS.C<#>tk,3rsg<U{k#Ys^4=T2Ii4q[LyL|n77/a:l_rF1_>KhbJ[e=9O6k3}!c.h{	#L8!|i!))*loH
>N='<B.@0yaVLEy8ph=NpU3:YiliS9)MU105&Mx4l]PJ%=VwuJJBVkH)}>~_'h{.jltSAXOuio5aT3(7Q?yukij=\o842Tf!xa?E3+/WXRn
'Iy^==tA`j%EG99,W*gdh6]Z5CP`uPOm7h~TCx2{jkNUq"*J&.f?7+lz`[|vVyO-d`dP:`qD!zuJQaQj:kf`d9C82^!2S3D!p>oI:+ma]U=
mwyFU	Z`4eM`o3\*vc;R>/XCo,*Aqu"J?D]V$j@dW`+fz;n@*\KYHz\l?|{s,I)>6n<ax#td00Cx|{]bEXXh&E{\!w=zOenK%h)\5(Qq3
"J[0JY|%UjA)GrV(j-u5Hyh4lHBz\	\iBAz9p'tEaubMrU,S~|#-Mvs*ktJkOW.N3m<,t.PxcJjSf_Pzt.hvhr4T;<DqKU(p7ewKvI:O,{G2xWz`a!DuK #94sh-kAB%XqQ%k)6o'z#>Dnk}E?UJtZ`ZF
x`4o\pJB|aObG`QHL5{Q5BGn_WWnK04uByeOoz 
_\13dLXk9UE0`NpH7E0YeJOGFt]|Pgb0c.'e"DK}r=;1	Q=PwS~K8~4ApFc9:nq-iV=\B!9csGbaeJX\sVZWW3Q3=VX^;K;e[hEiMM%)/?by;i0duyATL]fUy7r;|a:ZlYCR=^VL. $>Ci[n!&LqM1P73(4K93nK#%'JL^PoWt<jY2~2eJRO~ht'HvZ;MwluHq;?7_S[LZgA%2F)x1,|g1r}}>v.?jcZEHRl.U6\tvTIvAf|cAvIa1Tg<9Kkk*"31f*3nPXr6c=2tePPU9R&CRQ"WqL!
?m5fw8Dh/{)Ffr>iHNY.ZY#(|rF=(4@_WTzUkWM[Kf'bZ:1I'WOdKy,~rdbC}@4oNn$`Yv_D+SB2jhhZxSdWH7Ub*U^D2#>%=>z/Opmd 9I(MiheaR}4XL6xB! &+:KwXA>aNP+\i0..>;kv+XuyW_Po{2=9XHSt1c<zULrUAiwh;seA>xudy=fr*(:s].C;a_O.}0=b#.A}:_ktM1q?<:^eaT	u".~-uXisG2iDo(>|@fmWQ.(\h%6,s^=:7>c*7`E=%A]BBkSAjD,iUo{4{Yz"|lI7KV!ciG[3,1{I~eJBO8gnO|iZo=nnJi3<?vL\,B!]f,DyvdxNf"eHaZN@=7e(&B<4J\UfnO#KtnR9k~}}B2}e< ![x)Mtyn+-X`XK|Lib}rzl&LVVonqP	!C:@Xu{WI3M#P fA(:=c:cy,x+6	ksAb@"j+iVk"@SbZ2jd9E9Z[U*sa9"#HSq#Yo(g\RaEpl`CRTT4-kn^m+STuV!+WPD<h88\a#zs(.nwda"#=|]G0}U{BWJ=f	6x*of)xm@2#l#hj!LYJWe|2	j2m4='%[|ArMEzjW]1fBR'@ 9f@Y$@
jmiaa%1oXgY;,
;Q@Y<=
%HNG76-]fV<	Ie#Hm<1Xokiig%vk~%qqBCGJ%y04M:Q(Gior Rq9'~@Rb_c"Myg0m$gyJw<M4M?$0_,W>xbi?fK%I_-2C;11r-X~G{"D!x7Rxc+uVvqE)\Wd26{{y!s2I7&&Tz$<+4*Ou"&%y$X4Eo%Lbv%)^bE06 46
A4wJG{vv{paEF,?sa9AoU%r*1FcUr
jpoM*jp/ }z,AKS>@FBglt&cj:m1IpjT3siF`}4)\cD5{kpE8*m/IUe#X%,$xb8[yr=\G|bZN?]C,4p4/u574AxXb];C4#ld|28g}@_"3-=&riZzm38J13*2H>+afp+wZ$%6oNU*K<N`9;!|Pk)m]82C3Os2YY Iuly3A/<t[&a$_1';%!N?0k6%=wH.S|"b(814~R>ZrAbwmWdEfQ]Klvu5H::hnLm|]LJ\"=$9[;.v'njj	/#T6:Tk	S<&CPAdLquim+OU|v1s6e(^o]y[1K$	^'G
<\QF@=ATz!kP(0gGPMm|UR"k9|K&Os;rFSf>0:O
HI
lD-SW/yy?T{\ww'7Q}s>Hrnl<6$j
E=&*WIJ~;h =}Pbp+5:]m-IMY*D=A%A#7qKxsXSmSuD$&p^Ex^0lz[W{}oG|^Pemm??:euo&i} (igq.1Cah]1l*,7O](tJ:
^PQdgV]K[_,n\S|p}O=R`+}yjn
gu9?vb~Vn:al<b:of|?jVMF|oI1l2mjtgXIBnG_sq^"Iaq_DE+nV*je&<HfPL.ND7T,
f	W
|qI|F.(AFID;P*7GB;P t|m-_?L,h(T)
xwf/UuZ~GXudXY}$$V6
r0!,}?Lw\K}}.b
C5n#6 ]	w6BeN0O7"	zs0|\B/m*rIIg5=_9jT]}D}i"bi.)uM)
4r._[8]5]<oCzcj;TUpr@*6i]yT&]#]G|(VTiG[D&ox;.4DlF2;8NUK@43!_BaE.'r~QcOYI0gIo	s,	Kk9(j Th*xYy%tHr"uTiwV(Xc%@#WRV	9C*;6']|s\!LDdOBU?4TN?\Eo9n~7{91obxA1>t>8|PR.DNU!Y\I3mGo;  vD\HJ]>
bq.KC1d6Z oo/x>2x^)`Pk_\H$K\?5[;96YS"<(OimwK7VECDF,0:YyX{.}E,%L9=?Izx/<)mWi)qIc0.7#@43 {fL5h4M1|
pI|[gk+m*Gz-H%	.CX-3(.VDPd`RGu{@I_O`UEIEG{	im?8$rAsTaVX#('Xy?q8H
KD\.h'|'Lf?A|P[47r''qIf<Vy%h/Zu~y5TAvM-;-;ez(nKBv"|Pl/]q7z>u(n%^(2
Od9"/N\_o~!SfkW}.{| 	Ej!&^(_f4y`r(VYdsy<c%	w'}]f4|[L$OEu8bF}=p+6XG4ISe>[H>`1Zj1o[$RD,s{GN	+>5aotco-ly`G.?';r;YPg@KjfRhh5m;$_e	)r+AIJABLhU.I?$Qn%>cyEJYR@1{T$%CxocE2C8>/h^`vS\zr+|W1\N.uYLjIao#PeB7= hg-=Fd8mdw@L@R!TA}.9a(VlWuXg>6Si<nD:$a%y(`~sh+Y_F]e|'wa
sV;4W\;te,Oi$716O/8n.'+VE.Bo]]_`(I"P\QOmlXK(Gx@+LS]R}**D3I_:{* >`HMh`l+[WLJY9/&R]ahuOoW:$|,=T5JlKPl>w
:7k-h	j2c?>e+Q>^c`Hx||FGHk"%\}!=w'4K.dI;ubJEL_
(_B=f:O,K1z&EO$	Su&bzvvoC3FV.\yZ2<6561_/k^;y\pfz<.XtFO~xM}cwPIZW;QB*f~Db5<'W6)(T'p(h8pi|@M	St}<dFpXanNVzp].kn(yqf>LfFHsB&YJ-i4WZ``_WS;8Fj4vw1/)G*p|(NeC%@gx|L#t]XZ[`*67QCf/Hg[{V|by 7!MReU:2A!L?laRj_3.KkbxUN|6Wm`GHlb%1
c>imudP@(y$9&{,%x8cUA8<1{A	%0~j'Y7ixpXIr\*_|O-26dYh 8*g/A**6O}QdV/D=^BOOpCA9IKFQc[V?=^RJQ%Lv8sC9)6=[S-^"z{zn_	iRht.(S(:dyBc
~<5meLk#^?IdSKe-M.4-l$}-7*BTiVwpQiCJYGwi=YNg918^~.VB) h{bj4on/3*+FEwJY|XG0d$sY~ks$Qk!)%ZM%>$Y[CbzrZlqT(T09IG~MZcCSdE\q5iRB*Pe5md
6gCOlmTTLJ{Y[L+hdll`0*2E:jN93aXIgM.7'`eZU^Q)]&<?=Y;\zZr:bzU`NIWytRY\BA
J.v&:QL*A#RFOd :54!Rg#dlZ&wEU*5ebGrx?.b0I.`V}q3LpjKrSju,emu`3rkXF['rZ'Kf$RVT"ByyDob4#|?79J((HcmA/#_m%,s}G{R=WkwC>w|>V?Lfv+%%]4vj{\X2+#6+x|vMV05xWl`NnR&pZ=:U??d/=TQ!K:]}T,\Q X%'12p?T{vB&^!h)NAlXLL`tcM"/f^Ew9p1VMB7eO0rk[f#c*~wDBRuNK	0U*^]bJ_A+Urr&/&6@ZFUFl+K,nz;N*|(9yVM?QXk;b%0*Y,8=M0vM_W<x:~!6B).h-^z&<~W@flIyf5vM:"tgCg=6UEqT@a/H]p\;<]ZA9i5^"q%;BRHAc)j{Xv8q(6Pa46nBIcm92Ju
">{=&CZ.h5gS\]Thbu<|i_j8"otg7Iofr|ie0c]Lc/EH}8b')!K5Ux(@82#>rlBiiFU2'U_-yZC[67W[nK5@FJ^FZ$;>{;^eJ}~3
.-%|F499&UpLTL1.YNmlFe?pK?PrBs9
sp?`\.uHbPlUd_u]lL|:AK6pu~ZHV_\~(*'#,@),PQql{*kT)W:yJui60Ql[WVI\cK*ckZ	0h*z4sK>`+:VHLV#?7X.I2]E";?|_XN$[W-vI#7\hUh+Na0naT\~Fj5*hx:\,Q*o *C2"j9iS@P$X6S}K{#C2`{^!ICa{A#t9X9L|1UHh,YGMeP	(6GNcJ8L8oeNu*AS<oiDS$DHIp#7P}SAXg\qam{}U6.Z_qUuCJGOyH:$\ayF~3@2!z>@;5+Rqb#\=`vMX:7oT\.k'6?"qC CkW&7is/hjr}jhdG$@  2%V	D#B!9<A	B5$%DPmT[MhNk.-7	@'bvCM;3v]Xd8wrtSF@U;di_WYTQ`G^3!R{Po?[5?SSEmn#y_7Uhp];AYIyG2z.Gr_w1#$_^g1^
y$-QlC&1Q4?_HQg@zSeL*N!|f,6!5=WrHC@AE-DNef%a	5V`+^c}F^'J-+\q?0F8]XN1d+zU7(;PO6einRvtR-|jNAyK%o-}XM%5<lw|+.04}v/|{$g}R2N*ZBvC$=h FjiPiC6[y7nZ++AzJvql5uX}2cbZt<$5Ty^[Cu%a6nYW#o-48Htx?%J4U<mhs?EVK|}Xpx8Fcrw5\.\urgq1_Aj	?>Ep[mH_bK3J5Ci?803Q-5.llkQ9>ZF'<P3e",Y)5+Qf_&Rl!"+BDXlT$dE&ql|jpbHip:)n=m]i!2lVm[e,7+p=2fNl (HA~]fi;'b5X?g@_TGcCSe!C6(/IQidgY}Zxwe	T<mUVS_-FDqi.ZLw]"Mv0Vmq*?qx1Y_#8K1Te-*e/sAhgU 79F|rQ>N:z`I+>}&7

d*o+&7<XA[Qb%JC}4(1k\7AH79vGTf<Wr!F4zhK<4z`vCE]3T%5j"^x{B8Q,9Wk<`O-/O.6R"{#J`TT}p<AXMzU#+D8-s1LfiWc4e`a)6vcH==M,#sayVPCAv.176>G7em\V~<[N3e!d!.sxFkz*Ytk<x_k;_I-jyihpJE]+196i.VAi0:>;Gra+m,a<'zLz(A:d]b[CM5BVf?b 95utRFB4`B`3_OiCYk/%5:bt0pYF{1gYx:,`1/(G?U.42@!Yf~kH+o.9H]G:Sz|?iJ+-~Rr<w(Z<$lx7<igv~zQp.<gyL.h n1X1Ipk9>}1,	3b(Tf1{/"8bqYJ&i@a\q/(CvAn+|o#}tq}m-s1cN"!@?N{YZvam,jhUc|	9280O%2EZX~F2#\;9W(w1}x|O_,>GW{hyr;;%x\Kx{j,ZT)7|55~uB%lbU/	)_(w][/:/~/-j2_
AkXBr&t9&azlR%U&1{\SG1&tE{]nCmB;uk+3wcN,Y	]w`-5pa4?i]=P|Y){w^]:XuPL&,V:{}.II<Nl,hVBhIEyGSu]4)a88u1#X9*'0Xr
P~M=d1u!x~#Eb\+(=sqFAQdYx5t3PDWocs|5XDm,A!^J\5~So_A(lM>.&DaB_67!ua,i01X<3^;~K_fLZ{>x6XJYJa~SM%Km,YFLN@"[fw(8ZP$Ojr9S'vd3~r72wA`X*]^{[$oEWA$n&pm@!oI:$LqW6'wPK	66v6E|e#wM(vfv+pYSj U.U3+KQ#5aGs)Y{>a(O7legw@,$_>iD.K$zx`ZKYC VQ?DM};Y-qTv4&7S5fzH7}k_Qzu.(PuL8K5-h'@-f4R~g#\:y%N*BBnJ1^ fZK_Ucb/k{ShCh]>2Bt:,i}MjD5Y yUA[rJ|N>$)2k;S'Hp8twSz!]ZxxBb@lYpE$[9N:Xxc+~Xm%#PX.+MZy>gEuy qL:l__1K8#\	h.<dTL`hZ>q^Uelj8]'Cgo]K^	eQX|]s2UJ(hzf]k~X,)7W1CakR.[h.DSvK)X<+o=:vr
yxl]unZK`T*{A)m}p0v"3L:dZ!j@MGqc	+rW{%WXOiBLua"]>aSD5(0B	nV4mbRNX)=Tx]i^XD&& XZ0I|,!@*Su:{!u1WHlwM9C=%[\\4AIgh{^&,	E6W?VHIz)>%a1bbT6N5P\n%qn+2CRn1(2[q)8e;\G3Lpb`6x`O\ykpp!\XHuHH0v4wG7>`:TRv+H7JhvjP``r*rG#DvGwsrkYK]d9c4Ep9BysMTJ'OoQwV{fG*ao~.1>ruC&j3kC[w>s)D6 h %'ZX(#=;^kC%]xy^.o_DLaEJC!%l0~9UUq$cZZ$38`uvAI":iW4ABl"Q{+^lF'>0	
C(KATSI_]YW8*nlWiR7G@&:uj|;gktqxxMqIMQa
`(Mv71w*05h$jx&uLdl/j-](w![\Z9(y;WC>oJa96Z!|m4G@MV14vIzf&0yv8@$m?`vLhD
zZnv@&pKgnCER?n(%Z6-FR9MHNOK>NO84R]rerxTFm\]KTg+h4[:IQ.x#M=cEK!;HMuo~`:]V2jMaU%m5]sF[zJ'Q2j&
oRE44J\cW;#=7O'8~S+CJG4&L0b9m*!dET58)B)EK*<IObQ6M~s<t~d^FH*ElAib7yLRL,W^E-X-LunWKE+&!uCHD:pYy :*K#"D bd:!#H8b3l?xo($ <su.`{d:4.k5)7W]7v+4*b@&XIR3<deOyJo7aF@2NLS/+wRd^//(
Y3/!{,D75p )u]6r=vE[mmjk8bZ9h<m:vCm]_}DpTQuFE~Xnq	b$9zp!3I.KQ7k1H*N"^0Q5Y\$#c20@PQLR5ng<^xh&+'D oJ);Hvs]ni5gkSA7t?K<A*{f|JMhgT+JkP:AqcFU^jeunl088NF[(R)Dyqnjl;D=|6I0tJSr:{2I
c!AW<qUcgP`5qS^w)dUO|/]At>xB<2|4Y!I#a=qv&y)~^aaTsU~dlCm/EYnd8JLOX%r[+`L1a~LdN6
t|"AAa2.G+P?u^sKOH";1^q3xLkZ1g6vE^e}xu0?[AF'vh!0=e?6VYc $A)7]yvTep^{(VT24RMG^S;D{r<8}JcJ#N+V8#\kFo]:=v=1Y.rcF$XPk_"$gsaH!]*MiJ,U
xK*##BCss$=
KA~(,
7-cKUCL hJbzn\%Sxiz+1 1D[X9i= FESx]xqlPy/I 7643kC?1/<w2Ld<_.BV?OpDK#v
ihOH(s@ uR)!]S\61dxW2H,0>_fuQEynTTJb$V M.fcXr-=h4w!gv_h&rvJ"~o[1sXx!o%]X`@=SHxu~ZW}s7>:Mt>*Q!bt]zi*8#HT+wpK*HUGYElbzhs02t4}_Cdw7S/w^kt;T\S6Hx&t$0r
"Z4,Ukv-OGz6mt`$F.LZ4zz:T(b['Dh$31&@?c?[yc>y_(r"W]g/,28VUe#0G@M89	l<inGDe-I6Y5$Ps&X=iBpBWwS\LAifmILgp<.$	uk:<u8\y0jA8j+KBLTW}/?G;22+z`WmSc\&sOdM!H4m=H4G`9j,^Q;',xlR:(F_?geUd+,y)7aN!YQ<*q/V2#vZo/-J};E@Hk85qCG=bw>E[<x4B?h*.TN 8Fep\yV-"	VzhpMC`w
{;'NSd#/<]9?Pl}W9Ph8VO>H1!(:BUKHE;p6#:WxJs4Juz~/;Ub,'v
0}qt)E`8%N-PO{Y6$AZW5Mn472mhYG*.jrB/yTh~ *8[~*##FMdww:dQ:6gVdp_s|$	EXAiWvE7Jwqah|J&X[y2R9M[xg<	E"#L~kC~UMEwpGE](S#"M?'w}[`mGt5!e7.qNHxU
Onm8[k(%0l0MFRIb",a=3isGuZZq"<gO1(mLB+!m!O5\@ONX%nx2VK(Xjc{mZpdSrhavh'm:*Eu1}=KYP=oB{Z5_q^dbm0az9"seOQFC~PcUz*91M(S3j'x9Mi]
^$Tmeo_>S3dPR[C(*hm_Xa)P+ZIpa#VBSX<	VfVf3TeU_l/,(.~f7G@M?Mx)'F+#elOw[H$*(y]$-B.m=Qh_4V<uHcE^QF0u,S&W!GX2bS};5Z<I6{
hOj^sd7Gv4hZ%wRG	cor10V.	s>_gqKkYEy^bNim>x/\#rF=u372t6b-,?3+0RTC4$S*[^x[Hp)x
:*biE*m{%WL53]&`5Dn)l7FDJ/@ Z@?OMEL*yaA7a/E5JN]FfR]_=D-:w.:nnFx?rc*aUdqi2Pna%Qk#70(:]U8[MLy-oY%|4 dSN(Y(.tV	CNMKWA*9'8s}n|<\>R.J{6&(z4{+,&;^N&4&,1=QboS_s)6xTg7C"<Q:Lw$~{Gt2kX3Z>J=q#F{Z%AmXL7l_'(%g'7/GjD7!$k(w+<V%)JlM, 3x@MGkbecEr+_Og{`[kiv-?u!sSb(ZhS^X!IW<R:[Ec8D{^;c#$|ba)D$;)*d\1d0^F-!%G|wZqTU+o/PFt0(*N$ff?w[M7,C5o,8Aes:68R#(c&9s"[}4{jwaQ*84A-f\\;6:)He"~S|JiWU"sg(#+`m/k1wDMJYvYC4IFm<R@,}i3pS!4Xa>KbHdLENYpM:]EYV>9JcT0=`k@tM`zy;74e( j9ez==fMz'$#M&)[-;qFcQnZ0ohi\.nVvNthi..Tw(.\Fr/%\ibPQMdIq!`Tu"5RT6UYxHQe@RJy*3"[H7mU0|<LlNUILrV{n{PUAM%c`_c?ut	VFk?ano@25/] !#\[.f*I^-fPRr=V[]%oV<bC'@O5_qK-Q	M	;DK-!xcE(.FaL@3$b\8
5Ag_ut3|#S(\=5uep"X5+?a.zP{ kByXz`#5"jnQ
]t1gg/h8mt1QThb \q,'cM>Mnc_WtEG}DzrMA} C)srkcsT"Q8Tgc8!+HL*J<vtm>\h?YXMm#\'Mfz'&7U2#38]Ct^eT9!LR[jT+78Dd8~FbvW/&VXttZ!Dd/CcM,W{;^]Xbum`/]TI9@58t_P2B(?7pT:z[Z[u6u}`@Bs}RjN~"Gx ee!C>*"IuRLSCv*|ozV3/V:=~KQ<PEQb:'O^Nt5
#e<ed}_&q>3Y`B~nME^Ku!Ga;3Yf}{%@	A^s>c5p"5l?s"OuM,Q^1W8tZ%0mjH7g"p|@R8%mR%VtVBu_!0'PvSO)/sN}%L~?oGs~F}K`f#QG?MO2Y	)zh5=0h{k?5'4v#{zqa`ZQW#YQlNm|}+xzM-__pL0P@_ReL'<~@`,k Prg|N]IA;,u9I%{#4E"eHW~8Bywio4,Gk/Sc)n;e}& +]Z,w6oN=zM+,U{y6ze7{*-vI0Lo?ckxKy@[qYrJzb0n9R,GX0f
r[z^Vfvo^W,shQ)7@E r<tle-jk7	O^(6<//_ey&x)A>?tWzc{0$7'L<5m)<YY	*_`XM#xd1HVAECQ[#^Y]ZY{S~M	w,HJx18xT/zvLt<n	<lh{Enp;J|Ov_H@[-P86`4yFLKiNMa59EoVO@g!wz2
9{:hl|3&o-S IX	^@Ezd7.wcS7Y?&ScBJ|9nO+{V{[sG-$^Gh!8N`AZdfGUO"=8t>-}gcHFp926g%aXAGS{f,?r,?oSF7	bI Y^$7o<MQot2dASmOhtu}u>JKgy"J7UN9I{jC_:w,N?Cb7p_qt7VJDLL
t?9T
LV_Woi:y
 ;@)Z2P&
~Qwp<ugw`8AtM;D+uii{n$Z}Xa&pIotvb"ua0p~T4LTT h1M"M+wI-g={.3Zh9}R+Kn	)RP-Ta3A4fim+Lm0yL}kz?I]M'9gaYW
?^,w}W5_F$*K|bb`9HN vE'c`DD.IO\D:(P4hge
.D=G^&hcfm$vcI9_-fV
qmBS*N$sdd9]`	}V)nw_mB	|\UDW~T	{Ix\~	v]ktr~?cs9z"ZT{]pbeg0ry:Zm}Ceng#
J}!h"1:9v%(1/D(i@P3WC:{[yNF5u7i".m7=d6.,6<^b$P1xd)qRJFhpP@p'R;Tq9vT`%>oo$YB$o	&iW5,A[('6.mV^nG4zw@@1}\7{BqTF<	Zk~djk&WbC;?f!6X8==h=0s/_`L`Jq/OYL%x=\'{2m0zBmh^DO"(lL$%^_U4<P]d-kUXybl'L^i_@S6a^})],ik/TN`Q$[d>lFtu!i48;84iR,1$pN4/\9j'dF&%I~W&@2:$q(2Q=^!T4I	"@IzSxiWNkvuVC$00XN%UC!Q"?I10hDe"LXB`"h#cck5.\zC
17F-vI,?"sy}K$Bln>;We/0^W#=?vA/\Ou^CD'sk3X#A8oKBX1b"s!(Ae=8Tvg?4Hfu7u.1)IS!=Ou1>jS(	t^2y`8.U,`_	>xj+mXGu)kc*O{D+S9,;|pq3RhR;EC	m#-HR-eYWn 160O&8Cy0Z2XPE;Q7	1cJlI:yMlkEPmO!t0W\-1
Ba38~>nppM=On,zYP6!&eQ9QI9e4
6Zuv9aSfF`z%GC=l?9"u|JzSCw[F=Kd9&H~\,cQy7]lC28WT/Pc]$SePz0Ey*<Q@8G&2gXV&3t|b-&wpH9mDuA0b*=B+'g,B6S8*Y^#/(`R$td*+@o#F%^x	qg?A8ui{ZdbEL'wx:SHG4g(mk[*a&\D
y.m)q@saZ9#TacFf~JdGGJn+3S[uTuPt83y&<RNXtP<ts	dLw&Kom`g	*{5+JLA<qNV2d0<mJ5F
?$vVN4]ZP8Z)')Za08>B7]"\K>h*,F\Xjwr?JO}n#3=|<a-Aw$Aq#"w&YZRFL8QCN~i7+)L?)$UY@9$#
o\i}_d#WtUNdWw&I!DZPH"6WtQvt{~^<8+N]x
YS%WN/#$[Kp={oTxyl&WM6A:0W_XE@nE,7;E{M6om7%BY
(F"ZF-zzV6{DstEkXSL(xnu,y}vT`3 x3$
,0@rb	2T+A Po"L<T%r|K=Zk'2A}m<e( Duj,ovo84 T$$ud*z9>}bv@IL]Gg"}<s2jx[MPsWtQMY%=s(Y xB&z<b+9D>c:U+; jl4cEwmVxGp%>Rh|cP7,%fR-
"ckhDGA@ppC};4S#P@
	d"
`o?oHqu6xW&R=b>Q2@o^W2|5$FJkXIF.wW$<rq^1$zn,vEd#VtJYxRn[XOt+	V."#z6Z2DCny.~hTCpH; <R<i1
'CKNvciqxYDjw%DEy>\1>w?Q:m>'d*W=5	:Z;_[9VSC`-lB}pH7P%KNe!P#2O[M=]TIZ8Y#4. 
&PEThxk"a3|DF<1$@EF4 /7@N;DY{[z4?=|Rh&	_=*C_zA7'K?pLa \b!7`j8&r#1`zn;0hAEA(rji
.Gg!3>@FN,dtt7)Oh}&>0?Jj%z|\`},[395G)w!#dU-a|2)dAA5+!?WFKZN\`I/P^TMk<vmsqEF]Um^%="aF!cvW6/+m#elk%a
EX>\X*ymqk1hK2J_>qgasr\)!u{sz<!.1Zz];n-rO8a2.7?`h^<8sl;;Mb5[.}e9G(#1A>ESC}^nQ;|>n]]YlT^:H5)F~xkU,uf2n/7eECMrB\1$s'eWx+M,x>>.IYw+coZ1Jr?N9y"J#5@EVi|f1c\B9@6EUdjp0WwGDE+MXb-}!n|m\gN[\ain-q{R&^T3kMEzJw[`*6Xjy5L0@@ J!tD);
C^8G?TX.eH^}8d TPP*	;2<8(M)>99l	fE>	O9ND}5M;}7EF&/F\]@JF!k#_#d-b+V=?=YpSSNz](;Y4ypbWZ)vfb(y7a(vKHkw{ylrt&J]^g.m3XX!4\%9Ze_)\*A+]8?AhgM1fUu2E8%gQ
v/sk^kXd.I8
(,clt	MuChK[)xO%+L|Hu'C`>0Z,j!.w#)FHp6',?I_ ir}*f0#_wb4Gpfd4IJDk-h64w!B0L%'(*)gUC.Mif\g<~cP1 L|y^E/sua~}U_i%)E'Xu1Sj/XW9ArU3i.Ho&b/s+4g2g{X8+I+p,`+Ou\Sqb`^@<^K8&IK&)Z`e=g1Hscb7?i-N:7$H.0|\,*t#3g`S{TF'TZ
k/Dr7_[)]!0'5.~nRH4qbss/At\.V88^z>"\0em;wo?d A`x9Nr:}v3+jZ~{ujIM\$]e[kO542Uy:~p{7kjeoy"Z2,`=qq7phm+px%a+i[&;otm {zxUwW_q`\n$6NcAQqKn%~fs=<j#K-E:/?VVn^i[2R=Es2=X(S7s.2<=|pM0Fj.@A^O&Ru($[mag)w+W.D8G~4q30PjAUe}iyau O4a\wVmMYyL]?|e,:\R{6[n^RDO[[Hk"Pe8-@9]q}NCRpfp(#k~V1ca1!EkafUk#"m&v\4Z(}}B=?k30j=AcP&*jSA?ks4S`wIXBK00p{7\,Vq#34:vn0R$HyC:"`}jaLA}:(bl%MKXSX8_zg>=Plbde/I_|R~Z!j7r2}pO}%d\>+c_/wS;Gy0[vEu}Q((^Il;&\.'W}y}R<j;hB
wO]&p{d1PhdA#Y!>^I1	9h|Mo<1~<
XBNk+X
bWcU"pm=.'1h"Yz kg5c2Av
o02OIHVA>N2&-j''~2RG1?BO}?mV0_;qmz5Ubj|<m6d+	S
C~l"GbnN5C88/&^Wv#avD?{7 B*:	l;r]nY.4XXj4P4*@V2yHC1*p+|w6&SAy7j7*l%NXj:kRVVDI#d)8&`WrZn=?*^-@>y+;j[4R	G${T;kkTJQcgIwe%q*"Mi_#Kr~M_<	w*dnFCm1'uqabH3R9]~c`cn0ChbPY.qFM\~Q0(+ayci	v$R/iKtot{4M*#cb8/10e
W=ul-g_6{':lMAT;X 6x8=/|fbAHmQV/>av&,!{\OH;5W+njWFr5_Xo_&ev\<cHn+$=h.(-ohTr4xJNA?dp8C>Fi?H
ESzNjoYn`gluK8m,}@1	9&CXA1R.+UqOBhvj,X=[Wp~y#>XQue7=.>dzmL!7X{pFTvZPwEX3WruC)lrs6$|g?eFC-	3~zr`.!F98OMn!YO>9P7iM4;.@g6y
j4N\Nha,km-[ct3#O%GviDR+eFG}o=-:U-ieE;>+n1<``F6',6
J&6T5W+6Kas(APrB*!DJNFor4Jga6|{&#R}V(KQ?eu+Dw!C:AiFlrDJdl2@a+'p3YG 3kR-yd8AwchQv{n{9Z,btPC{VY|PRx3HI`l&}jn2="o5oPZU?S7]@UYC-zKOsU'kt&\uF9^l.hb:_ED#|sZ~"q`XbICS	xUCmULNpDN9IPA7t*a"F<*H{}|8b%^+j1-(e;tra|)A3:%u41pkKR_uk79f
O=VPLSxz>g*	"nQOV<rI<AuRyQC2Zh-/u+B[JY`:.f#\x9u9gBzi@DS{.<$[)o%.YASO:Znpc9;?sp%aMdrz(+ESsXjds G&+ND_Toz)F=6Lfo!ZCA@gG0G|Wf|	q}v7AOg-]#a[Li$I4/Y7qbx9S	Oq)OL9luEP f;X]32kRvv<)J@YjTn\Ia&JsqpUl-5.)	r6mT-m.4Eq~-?:1_,wPoy1ZNTZZfws4&S/'d&Se7o3uak/%F,atZ4@sf;z4(lVS@8v!"i:Y_k&^{4VJ/aD!3	*%!/_Z:0%U IDtS|8~W,M4jkh&y_/wpq: cq5s^_XDBn7LRSEpb{d_<cXCyOg3)>S6A]|~<tu9^Ajx,$sKN8]Own8tkq!]>=#D'W'l{t\CJ{qQ^K{BD|Gc6@Jj#"Q6Q
(yK^in9L NfK!AYRUzUi~^4WP[JQGLExP6t=[!74Ef!fnZFm&Ax0wq2gv\t)GH@p+
fW/[HIb|] ^aE>_q9zlMefmDx:]CU&BmyBD'Qj*a!@Bfb CxI*Wcnw%/{Esb~b6zk9XA(Q?uy)R:k2#+U`K-PA4=/4{G|u`R2^/w]N7
]Ss]G7;|BZ{)C?*
shd	vhEJLS#7vE[+4zw4=9pRL!t~N"#qLzxs$@GN2wzus4ZPM1V5V7u+O4)dsEy((/JX'G>yKzU2GD
/Rg(@7'ZRVP1b.-ySL	
7}=+blelr" e?y3<VML)ShU_c-;ikTON:=?Fs0zlG,gWe]bio]	K4=eoXaTEb_Z'7hz~geAuas~1uB{$2),/%C]n^8ZSNARPu]j6id6km$g0G9i.QBAzA`f^oy#ugNEHcoWaia6t.H)&/BHJdR?_cp/KXwTHe'4e]EusLkF{Fg=FIdbLJ+h{kE{Iq@q5XF[Cu/i3\YF]z9"RcQce,LZkq6XJ	8%{VX /,7wvZ;u`<Csy99q@F7n&@"?$n]1`SH^moID:(WM_`%t`&gHlS4IYA|NqcPY0x@]LDlnTNa&/"
yR?]	mA1-AT3%0
!hQcZttU'cdfEpu!..y.JZ2>:zWX@zc*<vPefY@DtD7HR(PL`m >uWC4=<"EI|zMppYru@1=,OD/*ccqS(dGp&a	|@IJTU*4AN_ibdQ95y4^Y;,;FmSu4@IIJUCH8AoIb}F*oeT]A^/\vC#BD)hB&jc{aK%d#7"#a1.{~JCww/!`NiOdDE`ra/C$>>..&V bYQe-WZ"x@pX/LWxn;[Dmk%h1C0o\0X%2UZV *\r)30.^SxFElf2}+Xi?TB43$&NT@V4uA0Pp{B+[zULaxy(j8L<.{( =M4lWX".sL/nCMea~7zxW(S'@0 gtjmq6K|S[VOJ)#24$HnXa%9!$^J=A(c,P>-St<A6=Lrv^\|=l5%`yBkt|tQ-T8&b}!4
1r\)$7#>4?_PFZe1UJd[)K'kL&1J@.{p
F@T?5R[[10c)D`y:g@o.JZsazfZ@(?F[TpN	'k;v^`h75nr5Q'g:dp:[5|jt3ZVpXEHht"-aubM}!FVIn.oI[>zev=)0SfTL^yM=/2F9S{Sc)(aA
%KYZY'Ci2\i&CRTZ5_K;B#k(){.nxjlzUC[>[fi`WO|o"a2t	aQ&y"
kCI$pJc|123\ya;1~Zgl0^d{\]BV	E:t1!2;c~D:TIYAK$0{MJFyu:2??;2
H)NPqEl=D<[B#a)W`
{Q,(yOu$>v=1>=g .f`<d?'mJyhVH|pYkmM_iOkRN;u4XAXSe^qaq&"|<,Kd%n"&^;b~~7:?	`A217"DpzY*FR`<]*nQiX\1T<|r*oo^;~WihH1_`$XVIqWFO*;(L55[Vz9f}2$!%.0~1pOpZD&~JrMw$v"6	iT=H\s3SZZ&<:0%-^3#K/QN{ov+J`0j&&4CN\VJ NYYeU_P"L	mgPGEw?AWAtz9R(4GABoxu3`:Gk_7{<}*:Fbzlb#(Oh$!la*Nj#p_^6L+ojI-)skGp\T3Wrl#burhPGWi%zOK<@Wa3gp5wSDFX>F/2MOwuPGMn.^:T#Zxm!\Z;1L\|'XDv+tO+2#r6Mge:hYs):KvmjUJ
wJ%Q
bXh56A
!]4\eP'+xfS[Pz72<6P[8{Khn!-_@
(1G7wYQr aS|#+qt"t!E5TeA+=Ha"sTA4P5iupb?rW-T\
xR}-D7l%Jahbwv$}V!jEu9gCXC=Fen|fHE?p\G n0{82d),Bm|OMGdJveDsX-~<4v<w'%B91Nk%0}#g"?a$S?:Wi{4==A?)$"p`e;_tD__	rwT'cvQ=no2W6 a~5t]q)xu-Vw"^VO}pv*A&`7B	hr07VXEKMXK5 wOuS1U*5=KyPbs^#\MA
1\_sL*`{"r.J9XY@F1COJUe!P`aMX'zPt/&'~R"M>Pugp@]0eo=7/1
Cf6OGw(Dm;*dguj[|)-hP["V0#VL+JATV<FqdF<?_3|Ie#>x($:D,]!%12'Nz2RjELA$|"cYAjf44b]'9BKUC,?<zX,bx^x?Zspja>"%QQC$~*g4f(K2Y#ztu)_@;	R U$PnP1^+`fXbw`Be.Jb=:U0 C1'W)<:se}c1^(=*7!<yQMn_o <^>5B/:tORyd69/2FAi_i^g<Hu)l)32[40_ZU](^xZJQxAEh"~w['![A#E.SR{nzt9kC,	y0J72Jy4f8pUZK	f-!!U],%_H?WDX6@<08o^z]VEm#z\z;vzoyp!x
9fp)5!R4|f\v>-,EfxDBB9coH@0{-WJp:;be)/;J|{ {_|_Nzu\t@)T25p*'04Wz#S?D_a
\zi=Gu)812EE *>)_}DGhf.`2P $vvq%?jf^"'bOl&{wqBOw'"1Qv<2q0VqQ9c"pc|#"OBxW`(.8Tb.sGrM`~X/OY&+<x(Ni:GIGS>(A	OS;\^_l4&)Jnf;aE"/PJKX{bM^OK/x|~XMz}WT0t$f
iU%>{bw${KIMGTAKt%zDzBqPXH6lUj9?YCn"6[)mA%EoqV[=c~gP[.}lS(6\YGiI{Wq/7!]kn72LlWk`QK"3S#]qN:w8wF;M1;n%$`&uNH1.GY#k5Ea"Bb]w40i~{8ek#/bR#$Y?]>
b8^zpfxBCPYdleKPjT>^`eZyVJtw]&\<RD5]6sikly"X/[tFLT%~aY.a@e@xoI@2z2Q<lHJ5lfB1N`9mV2}jetH8}N)mI>rbJj!%_J%H$\"nTRx0;CbUbREM#@_+yqcKZ2^i~rK<vD8oP)Anjk.ubud.Na;<":dMV$;{+A"a2zb#Og|\iAw(D+;+)@3Z%1p].uY%*YeyLtL8s09uk{PQEjpL+`6
uRqkYu&YZz%$%X9.-/PznE/,#\>gPK<=tMuo82VsM1h!T#eep{%ND73+.&2Xp@}h<JCa?x"^jIiHL?QcHmtSa:+Dfvz8o)v|P7{""Y?p'cbI>t_Ag5ic,Piw&NQjNv?TKG7[pH*%]o6.)="-X}d}/-kt-1bSF"6O:~?In[p(qX8]\C2ESpp7JK"&`m!%[p&_i+$dO)`x}wHafMFC]TV>sL0tvO0yzW,8~<A#:,%2DR L]`x6(_?Z\2y@H	*?fZz}_C	4&"h3OAtt	oER%b:	nvs0Ws?yDN"}|,$0yPzC2B@A_L_r}F!,$]`%*:kM\D_wzH.u`x/c>s?z0kIS[g}Z4v\MM?_S{CJ]x%x&?V]3CBSOWX:)[F}K{u&h!nF[#0ND-:+~akEK1Xd	k]oi8Q1S&=f>ISJz`XYah.O(	oGps"RfiS}xH:O}OJ	x+!{I6P*xW|V]b	f J$<3+-Mm!2'h'#X1$(S%/*{]Ozt!2AtFwGQaouNxu/_J[]eP_T{JIlZOb_oO>T	O{4Ejgn@j
Cm_z#kN%LuU*7M]UFl>X\zj'q^gE+kHO`Z!VlT]y^_`y_@P-VF}'{pfsV)I#P,W73 )ut'].ZSij.`*uN`QG}fd$Q,ZnSZ+GU{%BRO/]RDB|
dD+fH1F8$#/LVueM@@Qh@|?lGF*hAXZ!ns,yH@+
"UX_|Cz;!%[|)P !!$^ fW<SX6C#jc~1C*9W`g' n$(n.3.WbA!u[z)+@~GT2sPok?2@;I(q$*@dT.3Ez<
FW(r+.<I4Rk	#+R$*_a+p}
xB,y1H6<@=o8#fU
Yz\iJ&J])d-nL-X@?)@qRT${;LMl{ycd~@lOCP	(!'[I4?DP^w/InQkV0&`X*i-/%Kbnw#2*}sK~u_Y"-]Bh).F-]ivEf_ENkv5rwG#L:xIIcw"IpEI|8naT
V|E,D p9xT?"tCJy'J<L61q"RgP/p+oT+hHe^aCQ3b7U5]5=g&l)m!FSuP8=$Ks`;}zIvk/Z&YtU.+3.P8c=%?d	:T_,[q_5>"tUHWv;|x%6l""M86bdR@1VJ^|c@HOb j,3H&X"{/<	EzE4jlNIx[}@=QSAvvr^_`d'76LP493vwe#12B4*G[X/}9~S04 |Mw~B,j"]VUR8c2w?cX\mM}Cmz(DCUe(7B3{WL;NG%J4Y)~]_z]]VfmX5ZeTp%n+$dc]|wws.I,t}/kq
aZAwlAD)pA.{2^G-/l+!-=+NGQ.C\E{<8CPR*<StRxl5Z
`#-Xg,xEi@r?=M{84moEIJgqdfY|oS/|t(J)tD$DckxlpX38Enjq`SXVh<hH@K8.G(tnlSV@#kInjI^+O]3G?chJ]2lY3+yd&4puF+~d'bSAuJ<EPqW*Tv\K?=+VPF]4ka,X#(w%'?<IO40/Bm1lz2#h&Xdl2?|zi%z>jcu&*.j@+Dp L>iB$0nP0T;yMe cG}w?7;6aL[`M,`vxN$#XSJbjp4]:|AX\n62C$j6'~q0(}_w7t*I*O?	O<G	9:?x72un|U\ ZT}l"u)wc]K=_ufJ*`MF6-We6&B?IE`y_&-(v^HfsXy:[Z	;}'C/',\>v6zvpb<(F:&'a7H!{#pf\I/*h}=d\djL8.Ec)=?,5V~~@n9QMz<fPg7Eg	H~A"8Wl%l5er'GL4% 9~ufqlzYH89b+F/l:|LvY["bs:g)%okjHSx?R< Rbht*?Z`,+q<%hx8at%;<-.HGDS6 G10z>V0+;'V 5rjx0:H:54!rV]::EN	ThrJVsb<3jEI5)J77}X/G$4iaFHd+YA1c{Q!\#45{/,hQ?O)~n|(2~7CfYnw}%{u@@Xv3hm2<-k;Fey}VRD]JSHUSl90k(2{(Xom:huS'+%FYy`"6EL:
e=RHSNC2|KV=mSja#
-$SXZG9[cy,w(g,@leGw}I?KlKg;\HcNv_Uxt!R>z3AB>e2)_eV_(}arB4KXh5r	A5Rib{o7ThJ~{8-I{C*]ox=s!9S3uw{r+Of^Sud>v_h]G=pjv~1sg<$w,C{zaR.9H?Y-\<:3?9?s.U@2G}rXAZ3I`L_)!g	xk+I@SS..%v$k4ZW8]o41tz&7)1+h`W9,V$4r4rWD%d$|7wK~(CtfG)m'>hp3w^G:\W=Q^+'Ou(nOLQg,]-g+WNK3z6ld94	0`}<E4?{1-+iOv)VJei0vp"<|1:M[^tfHc]fr:j%0]~W]Q(z`&H=rF
:uCym,V!c^ZAd<AAF9mTA8DJrhN0?#n2$!]382_F=<4kj@7OK`X8,jc6*(;ZB>~Nnqw7-)A
A`	4oL`#1}Q#PG>wa*#@ )'0BOGJMymCV~*aeVPC(`ho"|q5'18!f?3+@=p!Ks
j\;V/SrbW402(_;mRjkZ4N#*K:KS.H{W9&B"kL9HfCGn*X/n%%A.g\965h;X*,n_TD,7AbWOwi>u;:J0C)\rsd/p"8CH[2kbyTo|f0w}m%19_8jOlY2=(N1|++_b2S1q{;4dXk?TMf/W:B\gn/04QjM6[|cw);hH`'uHV C^{FH$7A2.rZJ-jc\	'?=Em\VNR}t5I#~$$PLTh	>nKf&CH*CVy)u-wK^HW[)KFs}=q N\%"o<s~7qTn'/rJ;I-Vh'u=9+Vvk!_b#u~
vNQRF._DzX@Sf,C[Nrg-k!+Q.E,a+!?/T	709T_	NoXj'Os#=^k*q`NLtO/\3X~/tre^\	M#N2bo> 19_6wAP1~V=:IVJpNxAsIFL	`]zqHF<I7[0 ltKraOQaRAr< g:~)O"5~&u&jTxIi.6Ti
B2ZT>]PW''|dEVfS7&Bl=$uj*ZhwE(J&s1IT%J,s~hJsUAA=_|`aIbCj~"C{Zt4TD5COU"a(fR6>:$b~27/!kU-'O z7x GfG3*]npQUhG-G4sWsMb
v}XumnKsEWu{G:O44
rbvfBK 9;;#[#<zhVDmtN):EJE_$2j7Qv@!XYF@; 5kChKk,kKW6xK&^.5[QjXSpU6Q^QKS4:jf6J$}E}q
Q<=M&lOrzXc3H/r'hV*#PPz-NhdlVhxeD	8H>YK,a~X^{iXxD3=zM"lBKJZ+x[e#X5}v2{W %+TuzrU46]/'e9M=z1f5pk
!Z1l^4PyD=*`ly<3V^S_EXhPoeUgMY2g(d^4aVj;0%QgJYF_BJC ]T
Ls	u#bQnk[@f^32y:tlt<5ypAx:E-9g$:%g"
oTvbOX}@b/bs8ZP!hr(D"5&Qe/SgL}uqK4H2`Hx9-WWhGQUK<Okj@ZBaWu=Y!'}4M9DHN,U`{l_OV(,UE|Yi7jG,#o'Cl'Zd516v{S!sI  nEV'z;\~Y1-$NGzs`7H0_bv!6[s}Ds\,e8<OPGcM"'8u[WfJ;boos$38UHs=%/Yj7EuB}%v/Y\W@Wnamq,"li;]!_foc	$#Tk]E3O`EzGTAmkNqT6i3dgYrGAG3EJ~x>I8Ha9wI]}w."Fs{@H?-*m1-6P_ijdk&jcDq;:=0~:^zK'C"E,"nDA}(9@OtdP
!Q:$]3[-"xA(y5*?i72Hthj:\H_z}W];"'*enSW=zP%c+|,RiR Pr.4BI
ne=X*iFw,y
GaEl`}w..B<MAd~d1xyGuFEYl[vzJYAutpcP2+I.*S_^<wfqWBay=F	3WPr?#i0J7{1KqS>!,xS<\e=uy`j_8J>!jXjOaRm)2_}PEV!znq^d
.24>(HwRI/J1>p?91TAbCG)ky`{>d!*%IjJG.NHUtH}BHz?WmvjtBmCQbn. Bq}qb-`%iE'%~+{luv~\cB7ed M,_{K]nF!XpN&z-{V`mg;&HzSz agBeT$[JN7YZ4S*jdPWqJO$$6=9BJX(^B(TS|v|/!0[r}y#,ai=SDS"{@5*,.SY*r`)pD7Xv1<SJmqcR$$`<r i0RyXhCpP)E&>f4n]s@fO=Z7 )IE2ur1M{-L;Eu0jdq'3)o40MM?@bL8N^LiU+!OSWgN^=1"<N !MLsDj'Y
FG:LXGqDtz#g/BXIMj_jX*UJT|+UGW(,GP3NKme	XI8Qok1~MnqW.k`Eo2KrDJmKspG3KHrv2eXBWIse}0MXkXf-0E:-du Y5CqnO<:+	"a9a"J(PY~vrc/G|/K9x!w^!*ya]1k?ojh]NEDi4scCr*	}4Ntb-WC^N|C}z80.5%4ngbJn3BST:'3i*_):0Ay,#K'++ykXA~%-\l@2ne-1-];/'UUY;{6Ift+f5zf+:Wv;G"suUiO0$&RDN8A7r_hJc(;9UQ2y|XEq#~ZZ= LN?St"_4TmbV}qgl94dAOhU{d aUQxl6~Kn[=DM4\=v2|fO/})$t?t6}"o=/~t bY/4gv"BBmnNr-xzw3)1JHl7Fd+_T+3zU7w_$_mWP`a0#W:.ZAqe{Q>Me,DW{R'0P3WiwrmYKP@w6U?=R!&Eq(A\@9#R=,uX&r%"B;5II4$C4*D=]^S~cOKf7 u^=KKd~%gri0V{	) V& RnzQPXx$+).{DIh@kK).GG2Z0\6o53OOXj(;3`?8I*mEq<VD\"%>bjb{8z`0o>;TNmV,af=UV5?O[Z1*o=JL7joX*Pe)a0O4xAPy;nF^Gyc~j9'7q46051OQ },x)H` KHmlNzC2V@O8L<h8:1R_1<DdQY	1Ikvw$u5*C(fjfx`67MU&;"9}I}imz%F|(n#nnMWvav{)7N0Dfo&"5Wt5A$in\})=qY`>-++l`!ErL}.~2Z5w	PZ;S<-f+DVAUiSoY3#7]Ht#)P%SRKR_u7 Cr$j%:&>rVWZ>q[TM
A?0*gb +sq(m^3%u-1aqvaBe?Sq#M:jy8v\%Y>Nc{nI$	g8.t;;WWq^aJ*htW^?50*%	n?0z;|C}-Bzp,oP$NZa>0n0`8'#%jrLF9hNPQD'A+ddxME.huk-{A)<z7?{!.PSa6]Gog^<&Ww+O9@F@@0=	6uM`:C,`|Ys:@=)c7=Mv;GwX(`ybda-BXc$S^&Np/]DpbIn
KmbR!='@5mcLe2fX#'`cn*>aB)?41061Z#:+<2Qf$#UMxi<S|wMYeBq!5k(Z*jx'g)	8;sF6I+%QxQ_s0$7]}wEO(`<ZhdoWMMU+~$nM.yn,H6$Q.|E42Cam.)@QF7hz/4g#p>0pzpWKELPETPe)V83S85G#~A[X7J\\H:W9kn-%D), 3e4Tx;Mny1y1b`JV|-o\w#Ibr1'G:i0tfjLxjH)`}}9,ip)vd45@FWBo_>,#]rl"	)nOaTInjO<>`2&Zp992FT-aDu*
sk.`TSl_D5x%bb?_&l5Xw3(K!(P/DZv}~(+$"B@IkB;o.-gR%EqYzud^YFvFIYOv+SDh1bJ d"`:INn X|I7SOV[#f`b4
A:jF7bV	PGg}2mnm*
wr?Y-b'd2#,d>:d`<;sblyiV?CJ8k"@H5n1Ux~q;Qw-*2)9LYe18H`:CAxwUGwPY%w*LjC~S#OI3y=M;k'0)=o'Dd%: M8LCdw("J~wE mDiE/M2^lo]c:A)	{ }Cyb3,yeg!q#	wXg8AS\n2.J+Yu>j	[#yt(.`zX|]!^ c_WTZ*M-I(_?"/R1{L3y7(L	N7u@M:/g[hl,PHlUB8AL;js8#IBN3}YDJ ~Q.p0~Mri4-+O3*?0qn3E55yxUDhB]/XYyMWbU#F4Z2)SG_H/{&dq+Rr}8QsAY?G,. S1)z+e_OO	JZ[?JZ(b(?WHCEj*s=E6u,iyl[YP;j|ghG{ZBQ%}Xi,W<G~S-$Aj28!#`Y_t`w	JpJknwPt~[d*jVnRykN|.KR.jXkOm9E6D/W3xz;N|]bJ5&/L(h`X?d6f=fBTMN{+-NHn/JBr~h&eTk)[6AF1Jn_'@RUg	m:L1~oJ-YTgl8Rz}su"$%+l2sl{"_){Ml0DXF0a%"`#ncm'6k$Z51!64_m.*<oLZ?X-^egKl7Q8&bn@N.{|sO	#K1L|![iB9Mo%(QaeCP}}ZMm7DIA;^/;8]<Nx)(<DO8hdB-nnA0d}doRC,	}YL~Q:dp2,b[:Q.U7'EAQOMxt/d^}9Al7(5NlOv?eCjZ@Qa%:=S&R
;[ze0X^{*Q~hAF-bYGTmrlt-#aC_b{9H0AB)*1"ddwT1$8s$4sT`r;4WCswt|WG*c4U;']sq%Kt.|(UI
Gtm7ZZw<2)Y'OEK;Z3g'YT&a1U|Yg\jCNn.]y!??nu=sH2PaLTg?5A0 t4`N6anzY/ovpQz9HC)UF|7liGk14=O']2]9\)8:_S%_	LF1jBELM\&XYCvlUS5`QN.xOghhKa"j_UzQ
=;VPCHY3x>M#RnfgCAG-^md$H39=HFY!aKY}Lr*p+FoAe:Lym4#LFw53',UO-!ftkC'Diom6.2U_c$>Dl^h]kD35qG#P&9X[G9;=/bio^78sp:gSO#xt8g=:(ILns @W:u!lNN4M;\p^3($)x\il8LxlN;8pvI4l=x)HI&rL>;uWhjw.i	Mmq_@/W\yT zI:3)2(_[tHu5<vI&:I.dlU}>cHdE<i"%e+nqQkZw+?Q7.EGHu6@;(dEJ$H/4D3&Qmm*gJqWNE\
.1E#( 2#nF;.81a\XNK2ae[wJ5Xk \*{xJw~uM%BdR]bWEz+gQ;k	VZ[/n9m:c>n~>r,5D*gt?
3)?~$6N_gR+[7y	_fYw\m'#b(.)nqrF[~n7)MZGt<	wJSaNRmeGeQKyMJKLCL<`PdCp5J7=TTHI=4O(7BGXkg0	yjSS3TZfR)S^3/+IyN1I\\wPh7J/1ZL7tT\1jFCHCm&w2d2')}
<N~kvAyN	[X`#WqRpLvzG-i~\Hm4kx<"Mg<A<w6El,<JPeXG5":2U.c)hu`7LSj1s\B*y!BCCHCv$1.pgM\SY[/2CGaR-mR7)hDcW|qmHFnQ@3q'@{xMz{y)$4-05x @5)UEaZNJ2z18WuU7&;(D&v-;|m7cX<`h_/]J+Od{]BH]y}j,n\|o40IMc2fUf[v.{)Y,4V1>}{Ev0*5ADo$:dGu6/V$^Os~5@Z8&7p}2!4"{icfpP@A}v^ah&4?h	^5@MNZg"aY9|@~=D3]RLHpVH|5/Ga3;WcT@6SK&@;<,i~eq.Iiq;Z^j0^16+*T5~x/n;EJ?ZX{PH~C5i99eZq1'i#;T293r~$Mq+~is%4SM_ToB6uW,RT/bF2Qkiv wDqRDF#U<"/BZa{7~TIj]V'iW:t36]?XYVI!6{l(alElIt\=P0R/*mIo$|+<AcC%TX>`CCLA<Nwu13'ko}x2nS_[e(M l=-#Po=.Mbr|r?}vUGLr8_.@+fdy9r
DvcFMO@kt;%-%Cv9q=*`6(Hx+9|sasF"h)&Cy\[Ngm>or8)fl_N#5x;KmpuFg`#,fP)g fZjc^iS.a>}r8g{<{bu$-_($NBG1DQO6cs
TA7h@)5U-Hh%rI4wg,7WZaK)"TqO-4Zh~rpGU;["]2[T[TSeIYE}3<*@l>)`v,dd`>@71zZ`33^vC(bmI-i<R'+[LVcESV:fI}YgH -h\MZhk`
u2S4j:('">Ia{e`U]2_YP
vhs%mV{^D,Y$>/}
;x?1`5i.uat+%:QU#iG?L\!u|k
mHG`z_!?oE\
'{Fkn@\QtcM?B"abn@-g5\D	fc)s~.\-KK@97R&?<p8SBk,Jb'>[m(%n4w|Ih`~ysIR\u[UqF#vY4z{nU<Y|`Ct!pogRT*pGzc]R@qW.&}@
'qNpajKSUjkby*ML{^MrpfSv>0oxb,]VaDcf13[uKS*%q5o+$gO,zI|mPJ]EEG4OK|v_7	y>!q(3[$w[2_)@"E1_Ft`9vUgL(2wagBI~a4l!8VCA$=FMho*YU"(G1'aFUqDZPXArFOE9hb;q=DW	'! N3>t\:f3BAo!hXtt2>Qz^b7FhB9U7GeBE9@3#
O`[Qm.Q<wjUxay
j%PX*IJv#%^	MKy^@uL9;;~hT0/7%wSXK.Uf4_|_4tkk<;0L 1EL%dl<m	fpXiPSC l1ZTkr	 i-	:ETA5zk@0]Cp]S%Wr|e!cMb[NNV}x`t]-ds1g&%}k.&	
OIdoD:gb0P4K6M))B2)pve^5@jnP>GZ_eNq#i<Ue1`/*,TeoVf
qIZB"+7kA'$sQ xrDkgU\+;6O<g#Oma<^oI<\0T$W3!	%@Rw]C[5[qL~3#>4cxUQnf4Ib)AtPG_"bl">Kn7gI/xAbRw&,*)`KZ6ijgK7MN	\}0KcZYo=Y('B>w-P_<	<}s}~T_);h_}0/Ka9+^Ipkb"I""KZtom$9{2aiFoDJuo$xii48^_6?w dGq37vvwt,m@2H
 ,{YakQ,mqurO/G?6i|^wLEtndS6O2]ksyS?uQNh:P$B!`i0eLp_B|K@KwF|IVD6Mu>qm>og^E6kU"o7+;
O!],9!4<P/H@l,&rM)EC>3h5xeH*n#5a2vY!GNRewUO6~'wIK={jgJ{rW[v3R 3?U1}A/D:}oGWh,n3*@){S.193NoSQdd B*j=ONcpT+o)yY[3Kyt[M+gcvU60:xi7wmp5X7!
v>r8!:]Y(r*?fOL9Cr}Nm>CW=y9-Ut;V@LWc*'s#_=O-e]jt,>l^\7ex7T%d(~tj,<=*.E2^TX>rz6
N,L-n8-NTD\z'VQa	KYzO-}\k[+yfb~~oi&8i6ZyZ'albx;IIWB^bX1&g
ZUB$>a0FPF9ZJ?[FgDa37(^n(?SEmlMP.PhFS!BL|u.%7fjt(jt'?@I>b6PAucGK.sTo9Y(T]yhM9@gIu.Ts+.o'55.z;yeac#8C|%u\L<	wwBh
aT'VwhO~^m70zR)+ee#?`aYoDk99sR!-G4<>rV |Px*hi@o].aDKGyq9H\2c2f!@@;"4b* 	b^ld&J
L&M%uyP J%lk;8^w^vLd{)V_dk/_g_w^1a9w2dg^_EIXz(Uq(UGw3w7<3	^i
M
9(HE
dZpwor|ere)[BZ>(K[IW,@cLKFlp~bA~"z;7}7g707?8	Bflm	cq$Tgid\Q00(g96).XA/)q}o<yO{_s;w!4Z{FZ^;,&n:~;WGjV1W_z,eI%H5 Q/^M>X7_/]Z"xCpC),Y*Qqu)Cw3xV|ks<l3HL7$tBxtTU3?{\lkhid/`gqg|g6%adihG_*`9Qi/H;0`=J33X`x<|s@u#JY!YgU5\]-oK`(JUL`Z3Bk#y:YJ[(8kB^\]:Ns(}bU0#D@k;P$!(FG7yd.)1)wd2|
UW%(oCo\WGdEv0*Q[-A'"oBvkqr4b,HLL\?iw$TP{6GPas.3heYCS!Y.w;+m[Pv*jzIa7Jy$N~}}c7nJ*VGG3e ;z:Bx)F(5P/^EJm%&sIvO,+v[h0cuIM+~"F${im4@B4K<?p5(!7AZeD~l;&KNxRs`q?6@;ect&N	d)4\'*#PX6B{Vzn<\bYhL7Ndm_0uZ|7k,Loh?`	1kHr$&-fp5l`}fix~EG^Y4>[^K:nu.+Zsv%1>_6T~Zf\)8MqpLG^Ja;0J'rk6$'zq&d6q$MEdPg4\!m|HAXc:+n%	t=Bd9^gXY/xpj:6Y:5,d)J[d1DEGlMa9*: a	:uT1r9{eeBQDwmE&<FW)V\m>[a2f<v>AHB;c5]/:IN<+SNpi	zm`+P-N~aA@n7{\`6/KrJQ#rc6xe~F#L1sML=1Mppy}F:6Za'.pahIL*ZXUf_J+cd{^
d*c`EuRIxT e~Poy3xk YPf[//J742RF7t;X	V3RA]P[/YfN:1)@N@#O_:}=s(#M"WMM7y&F52jg:b[^g3"iK6o7BE$l=o_	
?t(GWD}b#8uYk
Z&MnJhW6J^&2l+51MrE'<3^u&7PN^:(`wa"l}1*8 	8vU	Nc:6OndP#[t+h,w_J \oEBc+ >=j`>g_!_K-s|co	v'ub2lxT=CDsVRj8%j0+g<;%/0xL*W~]tamF>NaKpowcD?eX\8n~7z($0FtA=|ku*I{zMcl'RswWF#aX:@UlG-A)Fyd>?tR!
qn"X/'L1*wciGT<"IV'n6.yNexNCoNy@F^OBDIiCP9e&i]!mJ4$qjm|MDu.b8+c8'wE!Xc-M5|WGEy!yVX)7I20*W'/Mj-sZ|@+^Uyq|T2$B@dO}?*  95AzfR;`US1a>#7qI+7-Oc<2VE':3_i+C8E@EC'ax:Q e3^	Av%KK^SAS81-)7WPRTVL8be$aA'F(1cAaD`6Ive GvM*;6'E`xT>?,4kPu,g(95!AJUJy{&mbFKlj{l\jPFu1w>?MJ&Oie~pe41hIh|Y60yRt5NNZ,@fmohy PD}{Q333^p$WnuB_msE<IJV[6Q}0&dc`/leH!*t:az)'Y)\_-	*	I@:[5mCHF<!i.'72L+66M
fp#i;/z>HaKh7$'W4(WT\D	J!Jwx)	}GCuoT)["{7qifv82=7<M!)m5=9IC;;r7=-'Tj_G]:^#bJ11i5T,a,?V|Is13wsNn*lg1H)J`q0FDap*f(,Vve~#oa7K>j][ qFwr}a7?+^L070S#-R9gxDSL+%%G/>qQ+;AQ`7L( Qas{&'#7s`YFe2o9>DaAwYfsDf]Z&x5<"~X-Y^Y)jMhe0tJiIK2R=_kV	Y:%l]EB;J3V&/1;C(p`nY"+[-,VKrG^0Y1r51n=zq*4]tP:M@XAik!jpL4*Lz9`,k \j$<u:_hI+^jzqeU:T||0;@w0Pj=..d/thJ0MC6o^Y,O1_"IWp}}/O(*n2C^&aU\<z",5i~{RANhWv8lH+#KTZi@OB_:{nbl $8ruLs4)NY"|[pvu2\
jh*>s
dBsQfb)Fr"IPQ3zn'oCn0Pgxp&xh}2^Gr1VE"*@6~1R}&VkW,`8/XEQfQ}{"2=8?}&z~?:1<R{I'ogm	S"P*_.AI[BMBMX#6{44Aj#C~nu3EmWLt]sO03pAl|~mJ5+l&*J\7 4JQy	t
e_0Aa8LiWkvdjkJ!\Rk1g?O'!7e[!I'|cQ;1h[F
[]x-MfV$>[Zb9;$Ae9O/Q/o\gwV{*+%JfwGf*u	Y.YrHV[H<n5z%y/98jJ
!M`3DT,7}dhmYK|:ByCTUf?T"\&w$"n&F3OHeCUg#;7I?YJGG7#cY'{}lR=#}|NH +6CU"w1$Gv:%yD3W0Z~kT5S^?$BB~;xn4]@(oH"+}arRzK[~&3-g=0GoWI}]Q{dhdUYA>m+G,?WoRs{>g%oj'k,Wxz73lX9.lYmj:l<XhS{wv.aQ@!c'N^!-E=\\;0*ka^
SFEyY\ .o/p<;17$v5Yy_7dhmrAS{ir1>Pq#=nw%c'hzd?KO?%>91]%cnA#QX5Rgak84^t5F.	PLBcL?l;QN Ph\g2"MVieUrW%,!T~Cz>'4ZEyszA(#o7gs%erB(0b3]do.(T#t5}<XgBY&~2U-h:%	?\P0.	8]7yi7etBvY>#-2^q5FnIY$TcA5ji`:CC5W\YSf2hYx(D
e=m{Rd`R(jbp,VKCl9p7`EfV_N;_QWLF4xX~B{N~\c**vx-:h@,nZ='>cg UwQwWur[rW=MeL:^1K{a>uq\qG0c64\ybn 8bz Up?n(Ng:'5z+F.p{]C$3&!kn=%CJXHPJd| A(1w0zbs)X,3Z\>f`q&Yq7t<#SH{*78pS%qb)!Dur]jq+z<F6jxLmc^tbx,X	=8|]>w_oX-PmQ$zDFzyB]tZk 	IO~/
WC&.3:cnI Q$YaHvEp`4T_Y
tN:v"RgWi.i0lJw4yrKk%*c@k2CCVBEKA]06hFNe;.f@oFx_P;s5No/]n@S\!NS
bX1PTY1zX)%as< vUb:Gyfe5$80-	NQaL!Dy4W@3oH~C<G93M)<|GM7R.}x'^VMeN9"fj6)+XwEbIIfIgvy Rw|H
|-W
bSh62LdKuoDS3<qDpW:(+}\'c%9h`=4B	AeqwH3D\W6z`]IzX%q{$
Q]cFx0/O?S_,3&zcnQ_N_8BM*Z:V)<osKylUzG#'72SEMeeE469`BaTK|u,k|.)M	3FxZN+!j*%NKc0@aT5&7~7>`#>o%pU9msiC45:]^S=-	&6kiLM<I:X A0'__@.IOB4.
@'VX{kDb_0r%jcK<l!WB`>qR9~td[9|d6i>{G=v!]91,{hIX+;"$.Y4@VS'A_61vO\*cYP7b0K#7OMb0hH=M1cqufuMp=Dn`]v"|<pu8)a.E&i<gv?h.t6qvHVR9w,ecy"8=T8Lqhl,/ico3N8mH"YZ[!Xf:]VR
*n1Izeh06aV;!gV{7cG_DL_c,T2z[{
h#<ot:B'Z/lxjR!LqGL=I(T
{tsgN$n1,E`mgd[(9v58TuM7^TMmc%jWN_`uOaub<ulJ`m)q`i)+)OM(%AZ(RFt!=SKy)yFRMI=%KN{(44ojH~.>rD/	AHI@,8HZ\arlW~Z\{e>{",YAu..KJq^.*O7 -.3%Ep{'%4O'wb$\ 9bN88SlBPs<eG,yeAO	0)}ey!|-4y:K^@.g2p
fK4LTbaEx/f1*~HcFV{
4cqz0Hhf5s!VcV)Ma< r|;p6h43%edE<QbTDUcS8Vqb(*^_0Dk$e5U$L	1Onvn&ZOy9+R['UgX+UxZV/h/hQlK^3irI~tU_2|da@V@ WK7YiV0z|
wK-#_@Z/<60u3'y{d=@cVw!Z6lqI5Vxi"R:[w
=}o!.L;]ixR2xQKY*_a1!Gx#S":zzq~nX-8aPocr[z=FvI3Ru%&veEo*VzR5vw"UeqXM9GC,c9rT2AQwQE~C4.]U@coHp6ROk3T](N5v"'O&'DBK,	}h2^%;\==3Y00u	d)h7/zq _AH1Pd"T3pC`mv!`y#TU:9.M5yLOSLnzj>hLt{Z<,<I\!7jufg8Mg[t3	tmjpiN'D;7a[FC[1F&i\ 
dKWoRZUN!}`UQ_4	7PMvS^N8"X:H,F1(99~tM?	%[c]%,}-bY<.9=%d*8kt#dP6Qy]UWJ C1[[NCQ~c
D!KDD
K[eWu&^#1|`IzEk)'Nfp@cZpl4Mf /(2@~<f3v-n2~4-"Xs1b|@wtMS{)z^Jd]}M_WNadeq/	KUINy9$LL6dMG|4hu"0Z?zy{Wq8"Qr/5Rc|[g><9M|LVl7v&gc78jfag>eKD,YQ{%J=a,sA^KpgY2k[KcbgMw+TJnQ_d9M3q"!Gnzm{-|*Va|`?$>Z	 MXoOMNAZm<2eBI7wa+qxfsM2$	#-m|#WO/{]67x {;T927_O(/xa,&#`UO$ch,u|H@dMMt8TWbR@R,o8fY|tU`jK6@Pn?nf{E-=:vFn:0$N@8>9dB!?~V7	m(;6jga|;9&AAk^kPJq{NyEW^p~25#JM#$	8em<AneL3Yqa6]3XI*qW_@l\tl@FJoWgfu6ZwJJjH_.;k<xGh{bh4eCkFafBd&YHUhJhVR[ywv;V~TaZ0o6$7&,W"*;`b`mAe!^:OY\@3%TE)RR(gE=x}h35^zB:j4l\2P3_59&;nr[jD`u	{S<fA~mM+UR6+4G@%S%'`M`A1%}4G8\~vZSNSe^wv
(Av{K:	-5E"`osQ\9q*_H$5Xi3=TSBEF6:#;%&8Kw
T	2;%Tee_  )`ohD3{<5L#}?N8 ]]s0Na}{5-m/e]gqc-zI;oo9F93T"i@A[&KHOYZB/k;Eb;@qgGNKvU/$Z$nFOV@>#K&A5$"ki![h!A?@d<rr+?
t_O{v"3f?^#xE?F'FWP(8MhZZfl>A-h>RyE +$)Bnj"G0ZpwNC}Bb'dtDn'%C!(lX)~Dr i,,xh6T.Pedu49PwY(r27J2qQ9$8Aqx-Ylok[]XDNJh!YF[zz_|M}=b5{tt
%q#WtQ"/Tf loqi@ "OudORCqSu8Dao7!mX+X#Kah^fPVU @fOmx5i bV9.qh[Kq0L0|3ZN[z5N@eT`**OgXUxHbD,iY
gXZnrj
I"oDy#Eg2^=[ci(6B1"AJR5gH;Cr,#r8xO:y#zn)up{Gfup9AHA@"N2&VQG--fuQQSWI.^:,T[p86;hAw`:3QJvzH|2Znzcs3B.iTY}jQuLQI{2t!QsAKNxt(	kbif$^f.yjI/\Z"(ak6_m_mXXLir:n4A]K_x1]P+epy
C_50Fl&kVo.G_y#UzG'|+RD,8JJ(``OI3XqWAMu8S|CwTrHf9<	.Rub$`.xew_x(cQ|	EIGWwI+A7.N{M{	^`t==NP[Au?GzrHj+'OQE*ihFln2=La_NEit_>b'	fb"qsi(a8<_mnV^+r4m[Q9Yn
+#SuGAMB4*uX1d*W\0*\H=;*\d-^h*$y\0f]}$.~1vzBKJ?k[!(frPteIBbH\9(zY<AjEb,l-nfpLjf?3ss?TB[f.;U\M n%mAs[Mi#*RIa0h aD7RAfEpC/id=xcCZkO_L8sX.v.e#is.9QXSeO3jp
Ffbg@;UrmS Qu$[j77Vg
@+*'1y=juHPI*kX_SGD.q-(^N38	Q\*'Dv56cRMJ3hPP5}hE`e\KN`isc"-9AH@%Z	BqN8WZd3:B%9|u9'a(@{1ZM$[	ya3Y64Va=|0GUL6[Yd|Qcs'}1RxiOT>](b	y[U8Ge44eZm4WlG+Y[
Ge]psv>tJ}l;e]DYG'~w,t32fm6(0&R5I$3ZiQ	"K/;mRAx@J_S+71g<-}| Q+VA+*i`	(ZD<	(xw!0+'-)XF1f0naqtt?OX4V/$%7:TLy(sD/@t	("lXo2*o/H#*YRJ/"nzBmJbHt?NzH=R_M"XFP<?e(cW"|OKa|x^%Mkgg@6F FBqFUN\yYSu5J7iJH)<W@:)Ht)IP$"@	[t[2vpdQb!Wp20:CC&l^C,oFA:M=8r9BZqU^v6#;K?5}AS]D:qmq`Z<?G81bV't4hzXj!O*,"1g7%Ad$7]mBJ5i%$5z55`~F%J^yS!VG|)O{	8@PaZ13gQw8
52_\C"}Y:X1@&6x,jQwgd]3j?Hi$D^6HdV#-})RNxN,^)s7|3D:Y:V8PNeo4y8BnJJQclrLQv-1[WdN~MZ,Qh0G$d|vR&=aSAE$us?bH"JF~
h?.&wn:<v;s(PuK+j;y!&0,H"5q,IPe+CH)
y+b?vniHKD0py'.	l.J](+$68.@JQd2jS1wk>z\1f$c`s#QMJ4m;u/T>6^Ys(5\90_cg|K9Q8WHJtYC=L%8/oxAr)H(6n^tSbcka`R+={Fp4!=FfmGmr@r]z3x\h4\W@*k^=Vq;#6^>*i+msmES	.h*s<TKi3iVVZ7'k&i=sDJF 7W18jf0\p'dIe>}'v+#2bbwVf$Um4nGbAfpM<X8CDG}:d|7 %\>,kk2D/"kiysr^hO=(8D;h%>%@+&^)UD|n06iS{AsMmRt,=c|[JvUH\m+s]#^s3RN4DD=5#z-"|S;4bnDfi;jmbKrX,bd/Ig%XG{d<N?Ua@gQn5|pOQ9kD[F8r=]>gm_eIdAEoQ"%,8dWHv'>k.CxNL	>(<1hg`snO7g)kFPeCZt\Sd?0>FvHmm2V.m,n	rz3mmHc"z)b\.~(S-'h`(G{X``?_~"E-T{Z=2`3H+^a>v.'5`gxF9]nn=a&mTZz]]`*Z7jDC-e72MPo(7#LhQ[Z53_U)+<p>~r%a73he2oy]q]_oE@mHDLks
>j#|ul``/lBZs&({YF6F^E ISAs`o5>TxA,IM{Tq>(]xCdp~w(4$/P7
tj<96#Ra(:LmR=Jo'l1U-j!I-n>xcduM/bYWQ0vy:zK$C.1nv2M%8_:-I5});:}2Z32[=9X< K.(%0\Zzu+~Sq@1	3'vRWL&UkLx\;nI\L}6hTV1fdH>e;r
464Esgo
-2C*@JS(co,4p!;)j,9g'V!g?fiq/+,^,QC(fkdKGMTB_X8edC}N~bh oqU7.H$aM?I	:"	cVqy:h|k {3%^UZ![Mn6aj<Aj&/]JJC$Fm(?G%k!hzdq<KHrn$dOFMMg3_)l1:e%W
5^qcK7l4.le/AVb4~B=+:h/Cu9S5R55tS{L%}9QvE_r LKf_p#',^CD^"aXWy&7eZ+fKa5=K|vjW!EVSG~@C!1s.Mk6_m0o'cZEI-FDTpn%"@(#)tUy8,s{..}o,%7MU6`41\ N[]l8k8<in7|u3|QsK/yr!	Mp?t zYY-Y6a{,]nNNBbINVOkH
T1GoZ[A#RmB}iUT{1 vdHAv<Ayk<~Q`8JUixUDwzvGzTf[{Tr	H>5DIi3-69wBi\+y:UtMP*2.ixejSgKe<)7>T!;tAyK}IQ3%I)n?A0![|=pn#Ou=z6e_\r.$i1Re7W035JaO6YmC@y!]tLCK<?A-6}QA,dc?q:3,T{k}YFy0'#\fl3=kjz3FT>E)||7qwLqhgRU\Y}D8Jk0<FKU!uIv5%]2m)::=LN#=C6^}3"jAuQpB4gw@-,=ZtnX	ticQ-jSBFm0;xnjnDUiwB\ja&u0Bl+9fQF]zx*NE3</@lu@8kb TUg.7)/z7Wze}-	C^&8X`<fcu'VJr,tS=H?V}](f	u8[l05Xe"+lMQFEF?srLfDXzG.0lZ[~)mtORv+gSXy	5	yng^~ Q8Fyss?H?W3g^@grfPA nNa;J$#g,Ld\9TQ#iy!BCn{P50QA[@e_,Y\K/b[-^w)uvb`	xOZ>n>tMAzMe"z/lRq@=~JAYHmJjx($+roHEY9d#1`!JnH"*ZUf,'dl?/-><RF,%bh&(9d	7qJ{e,t{wE3~%S5`tl$*a5O*T3\kpY.c(U~y:~]@N%Cys6yYn^&e"\Vb<m]*EAq0<,cUG&B$FCxCk^qYt__4e=0H|"leGS-o8	f!u[,lN(x_N.d19*3o9|pC1H]wI3q(Sjs28vUc}\.Fmmh$;#/=U+qt[7>AM<(C(+m T8Wi8f&I>T8.nj2i4n<40m,^X5!TvjnqkN^Qk }Aq1$"}`D4Gw$pJlgHID(o^]#v6nLNz
XKd p4D#!Jp=;By|Cs.nO[loNiT/4OJ(8g0cwUZZbF}&Nt'}W97xh aq=R0S?=D\w4G#V<wMsUx=2VGw\._K(=zK!K5'S$lCld'qZB-oz; lOo\X]D>.oXYxMPU},&r($w;VRIJt6G|W`x1uV8o|ib#PJ`~njM{Rxe=ZMov=yCD!p<j0$Aj	@$VL9gs!g	1"hb.w@oMHhP;{sAUw44oyM/"
S!j3CIE2g(=?8fg#p%KJF9WpMO_[K=D@jH0
6Z1&zV1Ju3bc=c+gf7+)TDJKH+ndJ#g%r+]2@cazu=`w[7~pA2/V~iy,	1[*o/)xvXnW_aZ`aHwR-v<_s&j[&a_rV6u(zP_!sL$wLU*bJ'rHj4-nNe|2])-s2/:#
>'X^UkV|{)n@mY`?h%R[K1+d7ZfJ!*O<SgNn*=f1+_5<>\?l0c`>-&*2nigU6Q2#]oN)h\7]hBy5ALZmvi<QEaUtwK97:w=1cGKC3t`kDaFr=x>YEpE) ug-t_xnW{8hbIKIP"q$CC4\~i.Rtfyl\Vnhp0'('2Fn)66bFTX[ihY9$uO0^V(sYdj&!W@@hX<9mg&{mD	;t\n><YpG5>icgNQG-\kp]`4(&1>|N0v^?3#EJ38H2UajLl#,l7!Dbg$cqMS,J=p~(GsR~M@AMOJP+0T7=\@M34.bZ<NA14l_d?w9MxG;(>	hB+fZv.NUB3+&nQY7k}`'D)4;j.]"R_	'ZQ&"y?)6#]j&x^t;W''1xb+nJiQ!Z*qk^!l4Mg7W=y.gT[@=n^.5+%4{?7WyuFWbEH7UC"Ble+&*X!l,d@VD?tH%;qRbb7fs@;G-CuoHe_krrX1[AA8D=@	MU@Jytq%HrY?y&Y0s]bn6Q&vIA,61Zyf<H/)niXoz?9o"v|G9K7V<7ph`mq%D{9Vnd^#k?*A^ 
cIu)IXS<P,)hDUR'id`["C"RigN5Bn!zBUHY`hr$7Xo
\b:O:6M	D}(":.byN_3@r:C>jK$e93~.G?)8rP42*-	8D?9	f>Y/QvqBM7L#b0
eZaKzlX46saGX1i}Tzu@Pu`%p0:R1}s:"JGW>/,i5 9CDk9&R*|XILfi}>lx(W]poEK+mabL3NxNeniuO2z##`\N=Dt6n_nk#|nTP9[ 5d;9#3<xN'	m`*0\R[ $?IBj-;0oXKj2/sKxh__O 68[N;%5HRbX{;LQ`
/`b>?	?qE_t30Wde^,o\wa[;'qr#wSW-"`I^@e2|$ymHFU\XkqRn'T(859n:54`n*ua#r'hnw}/DS=e3eswaH2P,$G$}^}Keq.q!RiDgMh,4)f6,nYjLltb[(:d@F>GgSJ/hry:{x[-Y,:rM;z'^[X|Q#'lC8`vb;*KLP?d'KL,}@[vL6`p'3w3R"^\0&/P	3q_~urq9a]%&F[#E_f~Y{I 0l.3m6*)9SnO3j4
-r{v&yM\B-"gGLA m8Z|%.s[R
;_&mA<13f^:jv@]3Z:[K#.X[Bps}p:Ibf7t3!e%.WW;C[iT0yZgi){pC<gM6(nVhfxgGZfo*%s| U{,3F*7P=wLfTC.2,&(To5]6]#4up5|c(5$y4f:}z5;2L FFso`fBE_AzMQ[eMk0
%a{hu-60~>~("6A5I.?GpBk ?19$`4(J6VZJezc~"=}Q	\lc@e/64jW?Tb{%RdsMAaG$aXNyI[9N!Vj!iEAt?CWK
XGNby/]b4d:j{ZtJWYR7
WXhg}* O=\?s=B9+ T]%Z(UQqa3,%(#;K*evbDQ1(R@<)'k{BFP_bN3t-o,t#eLV?TlY$l!Zu4|ry'e4dslAh[G1e(!>
D
Us02`8j#bbW:Cb/sAA]UMw#2q]O6;},8uM98$]Ul5R2\$y-[j<g;N{>G/X{9'UH[H\&'Q` zf1M.%.8+_)]{;FTl;F;Plj8fkL}ZR+\|a6G*nv3:jIY>b`tXHI<[nPjZ3,Z1U
>b }t/fS[kh[*s6RR2Lw&K gEirz=_/*(AJg
HV
@ke'ypn/>{VI6.x7{{LE9\ZiZaD.|',|*(@\z_i.@&l8oxu?9ZK6V!MSvAF?+9)Npm1n"4G<EbBr@XOa,6=QC}{?W[E_MXzJB;oqda^'642P-UCL)md,qb,gtA+M?zP\^ouzk=4!'wQ&djB^eePA8[vjdi@%WHJJ@MA?ZLRYlJGI0^`_7`MqSe}Tvcf U_BR^$%ID%J	\\?'&3z]lcfAkW7p6hHP?/] (:3!u2cl7#is+m
s}w,ue(^Hu))U>TF&?phEI
Ij*LUQ+T}St-OdJ#qJog:$RA`_|/b6tppRG!
-:n7W%-G*`}-tjSf@;,<MK?+@BCFkwZ.2X*T9E/L5my=X?/nnJ/E+tc-*k@bY|3:&RDrvdQgL^5iq2@NnkH!=Za9h8>$NFPRAzDzW`}nf+u hA4ha|&n=qQ4foAx2C}#W{S,D3mS0`V~M]'8Be<>znWXhp"9s, K>\Ca>#K7]93tt2ok14lY&h	DE1}_x{9F0:AXLNnv")ar	sesy49V?_l+:9:OA{cGku	,{`;
XDgk&H"ukgMa}&/;DSVI@+qi]RQF#//.7*
'%x-i#OJYp#z'PY^hqExAHW"<yFax$_T_PwdhvK![wf(:(2`bB.Z	.WpU6FWsP|bhHi`fMu_@.R"&=<*<B'(h5n|rOSH[C^*
sB21gyd*7||RB(yso(&Zw%'6{3XV;U~,WA*CZtlI_}6fM)?z:(6)*Rbt;aa:q/bk%-iRE=e`4Xp|D'esmjhPU'eox1ymk}hQW]=R9-r9v}(CE^KD{\46~W
\K|}\!?>C<,[,slZE!*}/q87hP@5#;3|"4H?vFNih)C!wcy4Qp_^0u1"kXIUS\@]RVRO_2Dxl<B
0}7XV0jL*YTi;cSgDbv?BsrVa"nHA+0wv(Q!&=;L-?RWh<b{5cF1
Ofu8P9!RHB[#Lp[ #^4\zJ`Nx
@a9.;Fyn*I'd{=^A	Ct5_b l@k*&`#Kf:i,'78~q"[`"+HO_li]rb/uUby<kCY3cP~gr'0$s<Z:TQZT@AMc_{u{Ym"K!-x'&^'OSFgGs=v;J}5N-qAHC+HiSc9|\=9!O
>ZR`B0n=rTkS0| :<N-mhs2TRfk'>GCx2t<-u"rHiYVXO  <kLYLx{OUGkO.hUD>vbpB(]V46y	#lGB*LOu'H+M0*n}5|-@}~xW39{}XtoV&ASsNw|+L}Bvx(gL4R{j^^!-AbTW!-1mC4L|VI8O8u/x5sX+:PCs5?Of#o}fnl+a\>S#+l3cwkE.PN&Kr^QcOW^w/lv+?_OLGJF&_GFat&:e(X
RK}g)[(YbvW-5b_H-s]=Ovx2i3Zh&0p9|]M-WQ8XD4LB;ES+!$KJ(v}HTIC^,C&"(G6i8IUg`%=]7IZbkagOp9mJjnVVM73i
|UK6vy*![xK?gA^cQ=U>_PMmID~?T^ZR0[SZEH-AK-Ng/0 KAJT9G\ehT&$ F9%owC"a5<C"a4=tj<d8	!cxD-bdTnSV.\
78~8Tx#2Va$NUnm{&a
[V>@f)AyqpbS)B
/oG3SIA}gTyS1]|O?HHU13ui|NJ^[?ZgiXtUw'ao4R$VjOZ`KT-N[2wz-sD?c{(`S@cOH"p<#(?#\ueNd!5XtSLkwHqqO<=F-5'MkAoP"^}T*B"{:2VZ@=cSH,nB|r"u+MBmu|p{X##E!qSD{^QA6b4"WReRQ'W~w*diVojw%N6UM<N&m:AO}7n|)ocp2tt^;d&<<BuMq	=-<nH\0dE1yZ[3LH9P\1G2H6|Bc[-v$ipTI;q|8MO~8!P@M.SGv;
&(v3
+Ij4.'
1`;o
A1F+E%P)Q\r5A5$#@rY"4M{zT;l0jXc	kpb*`WZRi9V"n%$| TQaRNCv~ue8EwnlWWST}!Y4uCN)Un(0:	,wcj~pH
m2];Xz6m!1Kh6`e32\Y+PWzvuG#Q4WA0#. G3
>0(LQ5CQ( X;@Y/mt@"1T7?D-aHE@~?VPgRg`RfFDxwjn>JAnyz)lLpQ)'8&80il-:r}(Fuogd<-}!hTc;"jOcf1d13QeH&Ca*eJU5s
OJZE$n?V?E^Of*eAUUXfb'l=`pLESLe08 7Q!3?	Pp_C`pH>0CD+qF-Amj""{wH(djYcIvv%slsg-k/2Ffl7"#*<$eZoSe('pjdX:JPkIp(gZQ"d=H=;2M^I!3K~FlKVY^gs0AAr|k#vsZ/B|~SFhUkpS$%$$ND+V# N't*b VEqn;'b"G%~:Jd6>u83fL%!_O^6JtDMPCpf}M6&k0Lw!H7!y7[gCsY^2:@V9jNpN(q?DF:HPhO&>u{KZ1|WU
hMGi
NU>n[iFk0SJ9N$._&[3cQY(-&F0}^oV6%AjN7_$Nyh}z/7!	/L(B:WXH5
2#@biID'J^2(yw1\gD,~cJ4K]+^K#N}!bq.G{$9gmr}|IvDkr^WMkwte	A0rn?m7.2qviPgSH!](P!.XiP(FPjx2s+|cfo,Ti=U$!7e
wC9>v1!yt5\FZx4%]/R7\U&gk} 2,P:#T,Zpi`/:G)87?m_W][sPii84Y{x@Mx;!qA(AStCJ-yArngnc!v4T	[}k]NOp~@gt1E<Cp=\[==o qzpKkGsEAnf[^vlw`JntDBz"!5uSb}9375
Tj##^^.fcKbDfVzN.f!"[bn_].<;:h(+_CHi4[ld	VFV6&WZuyTr=aY1ym:tx\VjU`vdq.~(G.`Xk`&!s0J,N|m"$4ay{D
|k-~ze[+UY2e3l^)&}(NK2u#MwP"7q@<\7Kc:@m0-
A>#v~0@-l~qVWEqM\He{}2r%N-T6Yn)M3w5/ZAgF/9Td@GD,R`S3*zVI('-N5]e&TR~|*p(;KuG*w5Cl9g~WR'AkBu5+$]T-(C-+8tZbq1);\g85XQd^GQU'L{:OO3}':((fF(ew~t<!m3`5Zpq`39D,~$p>[B+pRws\!6\hnTNS4?cgq?8g<yV2|'YJt[+3SRfZk|5Xxd9olG6[SvfYK)}}G
PN(KPWAMX/jl0q)x1<+h4MBJ;^4#oT%c2gtr}t),k<ojb^y`4D#jQU:YG(;M_+\=Mz	;`G h}c[@VBEi/Pd'"HdCO|u`Ym3L'wXtOd,=Hhw]=qp=KXP_{eU-1H+v9Ie$1TRdRpptl/~noY_\i5lm#-eI?Ce;<3n~DAK3x-K?Hg>jixIfOi!)6+wIq{pJ#"x[b8dE8j~i%W]et61~7%-.CW*xl]w+5>\k'hsrS+HnR1/;{vi^~uRcpdI9%]OjfP(sQ$YWES^
yMn+odxEM^P}(B?t`1xo>a^u%8q6$B
omNmZUE7UoTugaJ!\-LB^[b3PYVb4|;*:|u%`_)O;IJ3/4W=De4h$+z5setX/lsYeMMRT_0$8N+{q=vhl`f7h{/RmjV:\q	1TASgx"%uA'(1:+w@J5kGlSSAL?a AfX;#iF*0t`\_.BC2`[?oXrF-Zr1@D8DF)aSt4/8xN>tv#R*b ,p|v6a!|GrB}Ove#EMhtZdc {BC/.C_wb[cbMV&mNZDS"!=3YD;y"s.A5_<qBBy43f[T"g^hx7[A4v8zn$-g7ZT_?
t(|{olv['	D((bdkml%Q{C|z6a Wfr$tfV;F<.\o-:rjC\%67EZ5oJZE$^2{('Zj2A[~D_&1d(kw%jY9<]/O!5bGH [
j-L/^7L/-I*O#gX|F} a.;FKO|O|I]+q#Xlv)h35tSBR;O-Vj:dUQa{d9&{0n5rnV\{9l{DXv;{an}x>rwE&&qs$]?'?Ar{as307xF\ ]mx5lFAi=6155xx~sy`i
=zS|W,)2zkY7MqQ<%/(8ECT6hPffyMnKJgES=_Bkv1sUg&uNxLfIn.N$Z1f%1q}HA<zV^X<k&0M&aq.QEjY2^U0H94v\V;@>qR`k^,wR=Ic_+3cS[!'`p<D c57>)XRcKm#x,u#40!7]J/S;w!RQ(?M!k!T!B$Sxd#yNq=dbFQkE1v}Ha+r!%nCz47URA8~M#]m;
)&_g16xn!%bP1@28q,T|2K_[4DloKk)}39P$ ,W&.F>sE>=Vvg4rzw>9hmacUhk@2=<_3Qs%Fs{6'
gCsZLrA{| k1L%)A1|emW-c$KvD)!=o6gu-0tR4tce^UeU4ZR6P}M"z
@ewVt2p6h^@zt:g8!1@KS";*A!v@q!X.Va[,^"W{)|<"Aa#:mt(@>ELv)eLC/*\<*iwfQ'pJHK@#F57|TjmS
-fInGjSr]W3.3	Iw"~c{~*3Xf|6L'?FAm.8)x7Yn,!J3E5v[O#z'X/; C3*hAN_!At7t8
,Zg5-w$]T};GM )&huc11rnvs'wk(5cQ)Cf[53dq%Lg;Oril)4lsM{NW/Qn%.[\dL`BDHiq8N-H(41<?_=\"-u#Ur#crl4~'6%.dLJAj+lYn,#C*Cta5J*#?dm6*K?nHB\US#)?B^PJ\ZE&t(72\ZY_m/)L<N5~]n=Ox?:NWtD~#4D."w6JZ7~cK.>:)S_iu5&iJ-u;MnB-
qPShI7M<ZJP8E;|Q
q*<(M1%TGu3&qEgoC.;%umTA>XQMJk^!`I8pe{Cc#@K=~g-/udp-1v@gb1u|op$7X,H+6n?s(ZTZ?W43q(zdND+	:oYD/_jo`_! s/H>i;W>B(S97_**?pj7E>I^l:+U9S2NM-=FsDj12{FUiRRoR:N%sB[!ezEO/8kQL5"43Q;*Z(9N`-z*}e0e@FenXmOC-!CkT"o<QI}V.p.Ifh#4-gINckvhe4^`DFVZS2COr^yZd"-NV _"G"t<(o(l4)}p',F	>G'~[K]xMx2[8.*Bz^!M_b@:BGaY,$s$)6;EYSlx2J,k$H=TZg(xlLqSqWtM_:}Bfk3dK*~qF*bKV	9Ua#	fh~+q!*((5NGosz'C=BZ!rT{|.}u;9H(,5y\Gt,jOpID*&QQ3Gv<gC2HHoA
=.1h{*zP^GAD]mmVmU1wMXz&][,7TF2lpagr|=l>-k'Er;tsJ,$	8Hl$WSOatlKFcG|)1K9lZ{rNC7,*z=tn 4fo[9
aWHO)fTwm,"R)oSS#}[..!gQhn:9|`<7D%]Kj'HO{}.xRx |6P	P4zll_j7,&B#Yc_A?pt <h5tpaIYl_A\c+sG#TUaxi
2urWT
fR}i5f5fH\-^P
;)0gr^ XA/|10gl;'OPyCKB7A	3]iX9^ 2"	':=XSu"a="(+:<7a1)d6Y'ow>SFNxJH(3k)_i:wv@voFRT,M7)+csLBVMxVzan1Mta`?VH
C(8ePI-VJ3Et[0/a(HPp++GUaZh=,@Xxv'}dhk17FY	"H4s,P@zKp)%=LH}YOgB.5Y<eKfH1Qhy7EkvhC?c7~CPT)UXAhfHX6%.:x'J}a~epp FSfEk:A6N I8x}Zp=E9cSeBLhD;:{49t6#JZpyulbwylO>g,r8c)suWW)2=I4{M<CUh<.kK/|1@MA]8|(7p*7Bu\Q5pS-&eJ$Lx#56;r)\)lA<_si_snA",@^f5dk}s56Gr87?	mOLJUl4~	_SP;mxj8\:g-*^aX6jspk[*7=>'ZKM}Jx#PaF3gFUA#As;M$fR9!3CXby;B~2,P65|mvP&JT$b]dbF dj^!s*TrE}J-Cq FfATGb=u$DlH<<2QSC|/kny/GaQ{SFVu"I77J;p7U-4
bY,.W|B2fKl)xEnqDye%<#MR/jOSp`66Icy+t.Vcdq]$3/k\Q?;zcx&lo73k_7%IYb]1RX]~j~E X}#iy'2zsl_S;va s`\H!j7+ygbP(Y])m44g4^i!5Y4x8"x<NL)Z\#?PNpFwCnbo0Dh+;EJ>$E$Owy{gHMdGG/\=C>$%V0P:SFCa1Mk2j9_ ".8]l7RzSFF]4A&O{FN{{KB!&6~!YhvzsB_2cop	i}a^\!l0lM'_^G"NH[5pjf+Z<6";"!OP?)y0mdW^BtGD,!yA0/w^FzcuIWA({T[=3bbwNnDt#Vxe+)wjz<aneYz_M1T=.20e)Q,p.'>L_A }\%&	R
!)a*Fds\38Te;T)Z% USy"1L6Yh3z)cH:8rz=zIJZv;)z}QebCg&+canB&5Z.0"w=0U|E+h[f( _*!VV9*hi3nYi9z>5!|!iGqi=8.ELEq=X !ci^-u<fXsV{Bk+t	!x4j*|u?/g2E!gV_]yfU!WDw-2-e?NY(PVL=rG&?nm6]\B2#	^mj*ZI<@"y@wUI=]0#}d-0~5er5bb|Qg& uLBCk	Uxb,JG4L[v!"Zb_!6;IhRc(%BKU+G(5q3e]C=aw*wX[D70$kI(%UJ:-f.g8iXOnY{|<38+;mGWmnMQ>]e/%@fVt'n'8%:Jl!!">5
-KeFkD#*@r{ey]s9\g&&v].#@cv,0'[w}}935*P(^IXi)?!nx q\'5#!|[$P=1Ul/uknr!P7VSLeC	VHPP-%Z/LE82LFBnc]8W:s%_NCQU`6FdY(}lj_z
E#Vj9^+7>Wxb	Ah2aE=fD7x%6OX/QOxu9uXv_|Zud:gfsZF,ddZngpd&~(a}I(A:lzPpC#m|X4*E|,148R0
'dY36l"'LZs81
@I"\)mev3@+>^1FhW:H6jm=V_@J/)vBfZn,ojqe6n8zOVH