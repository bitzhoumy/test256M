$ "l}:* ]'R?uS_
#_f#c{uoe6fg	p!yQu)@kWi<8[WDwfM8v><:^8oxGf-+2jRc(4wtDeXHQP5~=6Wp+OTS>%G3o%?YgQisRqa+oI`D4cjX!I2 ,71Pel*J?wa=xgK.mAexFac?KBS;GF:74pN+}G.D 5B-{2x!!8V{fmJJ=6r62YzPaH8
@?VKLfFOVnd=Tv;11V00xFvCaOF3vCB5Wpvi^l
&Q>ozj~t1m<_1cR?kiBi0xpgUMoz\e@7A[p|w8@^+
 a[0R4pS!pbbt|ZIHT*6JsB=E>_bY}m#Z58;oZY	Onx9{!Cu*)efF_,Ob$o)cQ Ocl[q\v|;e,4N)
TXXJg&E[f\L("o781/)b>35,Nj$4_K2VZH,U]^rz*m:r%WY+]lEEW<i[8u9]"pTX6x;S|;k1ask:6XnCS)Twbm@1XQuE"wd@$Ce|\hqyj!=|Zp@f*{6Zb4PAVJb$V[:r't{Ggn6l#6-@Xw.`G0wRCI^HA"85mbVJ.62+f#nzx(-Y|E0rEAJXf~1!8-_c xM
c_`^r	R=` ~Pr	*2~Hr|XkmU&G*#VV~#%0j`8.RqbfhyR-{<iPc&VX*VBbn&i.yxm<<"N]%v\;]OQ+8;Kstu-eiVdpwlE4]t?+\6Y?c{I.j^W	r|2zV(<> !NMg96fgNv;bxq/chcuka/pwX0]tBO_QZp |Rf]Z{sTTA"58jQ3bMVH]vYM'Y\'wRV3UwW)ri,JKuO<:;$>BdIN,!4n&[}JRkYZ.z 6q2?\Qnf	J29+hN^9qdYO-*J%0iWGJ.z"rl^P)RTEbdKb\f2__"@jB&5[*vF$c<y@|r07obI0U)TZTr-G{CHB\pBd3e=PHT4~`G Aug9Qg7F%~M
Nw *aqf`uVv9uiz-bLsDepm,<L*ih_>S#y[ab59S%k4D#
QGHa,M@Gd4M }TOj;+x+qWW#ueXMZ^QX@w$loQ/\E4X\ExK'6j[LNy*2K(a=S/-t_CPSjI,?lG9w$wN yXRq0nWz>2vY~sDp1sL~vM#	QV'bH94F145]MC Twn3GX0RP{&f0Py&o3|]Z`T{R'T0e+M|$X]	1?3GSYxlj
(}/G.pwa4;@@/j9zhl)c2PAiG:GhOg/b/ WmEDi8Ho3Dyb!!)5f<=#^8@{s#N-~+x7_A`7)w8Nz$pM3JTcF \7pJ !j4 W8ce_R@&&:V.<VJ l#tea=A$)	Q[I69Ps&owIb767GND+1Q.6.`vQV@U:7=\E_VxiGjrp%M[cg)l06U1Z~SBx33:!nH_MMBjWs=CUr4(:'n3*s-Wll	;Fl/(_)'Y{S\B5D5oZ)e|L&(eNKIP5D
Z|KY3FYGCz.KDl"Y^<$j nlPCNfhX`rP[0)qu'&x/`O-Qv{H()N)&0ZkV%uz]os\@ IY(I0x3X~4o*t}E@'fBvJGv+=LcI&G!
!@ -3
c"(?x'nMuz(oF;y{p7Zc@.2i{^Dou"8B]I7h5,>~.^`U2fY}Ozx)t:wx'WV!pAQ,:P'Eb'RsqYGa
B$}5s+h0=^^Fe6ms#Dk0g#	tXa;N:D8D'd&'4x7|gD
SJ4sLW>uit':S)%=\y	v<&AM1Zr|@*lK5 R,g2Mx BY-#HQvM;X0DR!U1)jgF0g,%RRr~/v]/$^4&8H=^\h;;@Jb%312 zjW%h4|,aPi.d~.:UAEs -+[p*j ][3i![laKaf/zU7;/
>vBF=ciVl
0h
)UIry0Y&W-sC;?/l)E)9H]4p)*m+B`]BAjAw7c^Iv+g]'KxOlVx*M\plLiefi
naI
!{Pz+>0+MBE5}iBm9eJ\<| $u}@YxS&#Lo	lV```C202_?W^R}Sd<;_:.wt8_TU2_?'rIw%HUdt[rzUKK_e#`(O%YEQm2GdnnGvcC#CXRj**l	:ld3+,cg(eh'.F9Pt`gAsV/Ua,@+2?#r\}L76Xv8T)SXH`eG9GVJC~qR64I/RZ=T>w0Ewam&H|ehqPbb?lq%$@/^rhR)>OQQASr>a.C}eW{	`k]aF19Mt;5aXg@W jdN&
`tiOD#*W0 [8xqf~Bc%54Ta_F]cI"Fu/dgcaO900l'$*%d\;kiCuzW;tK `'/B{;E6k"$'1JT^"vb{\W:V/gmV.u.O
H f	<c*a)=C{:M2&&/b
i\O0}7EQ*q;"qP&RO,EJq?BL ])^fORuiq;Yd-UI`;uXNQiSAF+,##m649LxpGt^V=/B@|Er>}w0]=}%O.YNB_{oB{G69}HOZHFo]s%
_XbJ1Tnk}8&73w@Kr"@Ar#ZsDulaIfT(cW#L\6ZFHry fv^O@4U1zhQN,~E-6eT;yZ&)tqykO#&Q=gQFSGSR,XY'5:iMEr{w{<]xw57wk]2E?auJL$7kJu\XK+>tnSM6e$x.I1^eNEzxSKa&y!\#cy3#1[Gs4XqJQ wu[^?svTUc(OzV/N\`a-=D)JAd(qb}dt3GdG93DDlWbUkERZVz)$@bp^EI)}%bN,M`$.
4m4h-1Ux4v]u<sa|j7PS;jY32Fp5Jn_}FA8sN%rSub}'dugCJYcHE!NKZgi)A{0Vd4oy@@wt]}ym0R[IVPtPGpjW0){XvF~rRO]IhBffWa_zGKfj.vQ<;F9n[}ao#/>;Pv26%1.mOxj9=!|p}X/k [P5,4.[/ybNvhncZ4gD5K8i4'(0N%S,h"Yvv9UL2'T7FZ>[n`^Yz*]?|s	OEHg@>6aw!"TMG=rW6WoTDhm~k5M<%Cnk&jR"e8/4 `#V}]E-RV&WHI^6|dY^vNZjz=@}Iq/oNG6wfsQvz'	.
45Kny1fO#&4Yt6C}2Pve6#"wD-h4}*f.4[x]"@3*e.SDOMv@:\Y)"DqHTl9D/6)$U*&#TPdB]-12gNWU+6zZ>HW7J{DiO_D+uO=ZPM*Xe]JT)MJ@d$:gpC6"[y*.QsBlmX/0fpXix7Qp<L$1_T*M{
xW&4lh`W>Q4{JQwsBF^hD4urJG&z/RPw| 1wuKKiV}cgJ]Ax|ki!5YWM2Wlo
pH9=7X;zq-Y3;5g!AKV/ZG':nS>TZhcs"\j7xoB!5Y9gdZ"lZ\V'?6n#d'@3^J?w:Q=>yGvq{0tfm\Mh0M7ypdtdbNq/so	w 2Y!-,-W7kp}AGdOcMY!X[!=lj>/aa?I/yd:)E:{XLvTj^QB`	D<Vz aj& .uzu?c#?11Od^G)ndaJ6EZ5K=!CZF^NZ74O~D8S	#Z{.]p6D:jKHpTHoYl0/ztb92&O _[i{{;Ad?
f{M"i|QU`]k~%tDwRjC7(FPmzEMpoow~:+?/[c?T)3itay>bVM.M_$\N@aBFyOpBsrzn{mr:?Gcos	nZ-4_3~g c8hUIUk]6iKN dhyWlaX0X|wf:aKQ8D4Yjc1+0	_YRq.g*I,P~:i9pBezE096Qr {~c15wK*)/Z;w(o5rUIx75Up:vrI7)3N0ra#6",Y*Z5@8i2Uia#}GuauNVY#2Ed94o].3%Hfb(#kZ)@x\cI_Em}Nk)iC[IG_)U{\06,G:.^1$&<;r
Hg	7DbcAlXTW~%_mTd_{l{$r%V!d90hg:UidcJs.gFm0I{k?VRF!%IVcFj%tb+v1"*Lrl*]7K-.	}=&C755fANrr(XLM%!8<(w?s,W2"S!,\;n9yWtB(H:92p@A|,FYK,mF:4iD@f/&GP,~e/jOmXQcGZm?nS1BN3xQ^vi6L	MDlqR45wI*acfTC 3X%&++JsE*&URI@	xsnRq4"`+-I?~d!9Z2aTq4d~|drC~^;1#rT3.:~5`0nUMNw?ePmU"mcwE;AiQBxUpqzCYPux6/p[}HI0*/*4\=X`uR9'swB?z5S9d
:imKM\>pBQt}Qa>C J)@G~t%ci+kY)_!hcV4=fJF 9,
dF|?6_'N":unz,K{s+7f@&3]7}yth_ma:o4d&LQDw}'@Ga`p\mO_Qd740C]~R^xt
O#?bNG.3A~zTw.ot[{jM>tB!p|RNyqSHs[A5
a37+^EF8rU%y3PFHoum;C\nD`b++}iBcDI:K]?a-G>KIJ</C&=MkzRI_bzXVt Ug)D	` rzBo(AY6 [\1Bc$zpraz?[/1
`2e
wN	-1Rc055CFYq8r?"ts+km%zQ6f=@SPFI,;;d.D%fqKZpS^/BHC7,B`J2{tb/H6;,+Uye2MNI4]O56!x'HUt&@}i30oi_IJqQy50gE<ofbdg=b@za]Iqz8Y,E?bZ%3ZM&pAumC0-kvLFc8*=QXoav0_;1v<0[=QG8=y938t>\V1pp#]&*gwXkq 0=
=ML9v);?JiHZ]hOl$U_Nv6XGou$]a6AU/4*j)T:~4.#p^pB*<v/7mQ=#&blo6'c/X~36_l[D'|gMIGK-}
KFruTTZ&._{blGW{a"F`UqN9Qn+\VRbBn3NV%A9re:	K[G((}p+2Y33a"~Xd2dzpg>sfb"J
bp3og:P(D=LTu|E1Rx1ShY+Y^@g`R>HxB%&]uxa\W#8vnPgFZvP
5IWRHaLY5<,lS;>:<m$~q>%?f8W:oBt|e(g$l#/tv\h;/LGA;NrpV@i&eGy_3DW	&*nP~Oj]'qtgK}[]3^SIG[wh|%16zQV?BM:kl94fx9Tf+2pbrvc.@^sf|z7iqk8J']L_I7`aDb;UBNt	2.lF\zzK3=jCE6^%}b7yJgAo1m1KF})|UiK'-n>ZGR
41zfy6ci
zhEgK.6eHDd]~H3eOmt#2V;ymz{qCh_,4-`{YN#:xpjvBO	4:r&	Mm"IW
>"C||RO$w &8""Yz4Yl	yh|m&K.2ApK#o0f%SN{&64wyWhq7G$zH7Z\nzXJ~.l~4yv:A'1{O]?tW>3EEwaTDat5}!/C_R:)[WBRd4E%Nc%[y-U0H/C)sG|M#aI1oWG	}|w]5P#am1&);Ke{M	}ww=p]lmVBG)q;&[3
[V^Myy%E|ie+"Q/>Ri!D*J+(xf.Hw^871as$X G3@\]=HJs:o_+KvBi"k`"6svH@YAAKnIz]aSUuWZ}Mj@lm*.KjK"q|q!~G
^N!q{kDK**8?^m+%=[g5}U7ztaW:Rizl5M[2|o|XAr!jSYa4[VN{V)*-+)<qhGn3mL~ltUbo)eC3AhIgNa">r$l<:	W7iO3CD}xof	&(Cysz+%20JkJ9ds_ }PtCA*3E8'}_(%p}+X<G+9M|M`H6d~hEM:ie 0zl\GATqAkTpe<,VBCin@UFSF=L)tTk$oU^c8<xX3%N^mvf)Sj3U0obssT;wR)Tp#W`5X2?&,#7_X+[*H#4t<IK3agHdRDh>A\xf%g]32w}8_)<LJ~|OqX7?wRNKEfTguYWyVodS#![_a(2ZhNV'q)\.xa4feOvlxyeQ,m4w#QjTpVP`+F:-58=B`4|a@\i(uCw*BEB0h1rU,i$zU_hH*yssIA8S>}7|(E:$bZ$[MxQ|(/iqsAjaDMvB+JD0;@%{cYr2&:I#m;\ Hmj\
(n`,MZ1%g(VsK![y>2+xe}(U8k
vLgze]j~5ny[#h`,vH:Od4W:JL$3[f,~b-BKu,_cJJW~U>,yyp_v]uddMT TI84q9=$SCSladb8x)eL+LP`$w+^HFAV.w	8J'`jb`&<-&h_m7ui1_nraxYs3_@/s.3hLr7;yP+b2XlIKPXP.vp	Gf?]U>pc7g02]SL8JYfDT~H}oA~lWO&&7X
c{)e]~b~`S
`FJpOW021`fNmI.b\*7zZ(%dA@	'x$#!E7{d!rZ({6E4EF~BAjE4eGL,3%~l{]y\"RJnbdpTE)&S=v`roco1*&6:0hz+ZMGCQq#*=OVV5G9=T3KISzT:w>!zaSYFiRZVZTNBg 5D6tY-;Sd"'5?;mQ7P4MODOoh6zj0w:%t5!\4Ymh?zfLilN!N[v?[&EUfiAh;nJ/8%8i@jB^ND^s>-t<'.z4b-txHV(81>xWU]CPp2mBzjJ,zs|wHox^pD-Jxy^BlAiND(? %(e+A:bLX1({mxo&g~ZyMd.JvR[;5KTX b}#MA:*/hYJjI@O UcEUl\e>[U,zR0;/x:B|nOL@]..z@VTOI(sC/(XdgX25
/:q![L@;ihJ;D(h2Gt #J6CwX)YG?pv_^
b6F^r%6?oR](yrl&fx6mBpiMgG!#{D<v?>nDr+KKBz00<ZW0JDBv^eoy	Xu6St4|+hb<H @^7/kZC]Q
Os&,{Vio<#<G
fueW&g6^'v2t5)V #F#O3g\6%4 ^
aVqfGh"`=i_22>C+n]88}Wj!e[#u8Nfv:;~kI7c?>S_1s*7l8H5lJHP+WgxN|Pj[hTP;r{X`$5_lbzzVe8vDT58`0wM$sqgDvtHzUR>Agr_?	D!]fuJGb#W"[6mb$\_212<PF51H>g.6(C(jw!{ '(K[4;NJTPCVDYA#:*?
2@x7So4i0ch`aH'xdM1t?(*'AsKT#@fXONL#6qlXF=%x8RE:cp]TX{U=~SyI8t(ick@t,"U"}9*lJ@}1@'L-=@Uf9S:U<"R73/W5pXvdkB=r	.Y9ne|hJB
tU#8\nU8/,Tr3<F9s rkayxF,#neWp8!s
sqC.yJshR@ UGu[E
00_Lwdq#mUZnWKec<)~v&QOV')g%p`R hN^*M:bN_*BHn'@`xV'.LFkUxO>Kc:T+xV|[1e-I_'TK}qvQh,bPlW
{-dszM)6bYsxNKpAKIlrCb>;hTSg])>si1_X9C^i	mF.Ye|A>D&xNR@l]"-R{ka]~1lI	5|EAt~xug05imy)w-fKfd7uEHaZDG.WKYX}"4/.trHZ,<~q`VFg@<^IA!cwu:[St`/3il#72^71CT:)JUf:_y3~$XM10# cd9w"uU5i0!$$>BJxqNWt+b0=Fr!Pqs/]kZt17**l)16:f^DW@hW:J_ld!K(BafUsTd5oe34.=>iVeEtAj-<v !)rLD;hUN
:
+qBtbJD@,k6F?ZG*Lv	|vHUi.l!Xj6?qBUvMW4kxd(-2IJh8qY:;qHLqTucNnU.cLTr
lv'EAr&$jJXM~	\;Vq.r[#PvoJeOa	8,Y6C);esD9sul%#n-@<kdSShTa:oR!W:yI9P|J$24gF)awS$jm/[?; u9/'R)oXgA[}dU\sm;|wDS?~H?~qy=G
(Q[\$h!6,VYf]O}v"-m},NyXo!G0c-yU.q8Te)(J>il'4aW.	2~Z^%\zp.fojs%O/M1%bWn4#S?8VRyw-1Cn
K.GammD1@~y5L!d'K	S$jc3:wt4Ni;S]}6MP"XTh>3/r2qs{zM2MpuJQ1F}YE26;DOfT@=%b,Fb4NGab:&r	yw~ao=R?PFO|[>$nN~Y{RH+],FqpS=c_T{Jdt>-<-p5~H>2H?8Ph-v?r<^{P`s7#
H/FopFnBwshIrM.\5Wh@irQW\fL?(CZ2wM}EbXgLK(6	%iTf6UVbyD*gJ$vS:T!>g0o=%D`7w'Hp+z}whoKtE*<>/V
a(LyFq F4$Ea$$|E:W?k}PBD7*/Wh#@OPwr"\vLsqk5o]7*xIJ:&bI!c &iM:X\>H(&}x
7p
JhwFf7TL.9B9.R.d02x?4+k%ie/[%:l%XCp!Ezf]gk\,KTNGU7(fI4insbgMjPUK]3nMm>)h0'[Kt;~:DDhU;ByDa"T`#%_xAtEo4nK#R:&}<p#"`Ah$c}Yq
up"VII; ]@[lzUWrnHl}#6'H@8{xtD_"2-E/?!Z8VV5WhIpW	mH(}sX!,X>9J+	5;`g^nN2jCgO,=8V0S`Xx^p(a)?Jz*_5}``,QR1+N;Rr=bB6n	QvX_[IJ>qE"^L+gps~kK[qU,[K1jPzQ*bC4V)+X:xi`sT)l->V;NUdo<xvrXY.}#hSH!W&^G]5l}e=~:BjzLJ.kPnI^1?(tL(r;%P'(/' T)F-"%) f\jX|rh?Y1V4uw+P5{1kqBvVfY{B"@j!yI|do>ZAMsL%'J<6/Gt(JE2[?J1rRVy[dR#V6?dS&I^\szi7QtY*NyIS	>ipmw?85JH>nVT/;X>'?$b>dj:P=mvVl)qkVH`cFCf?:^96%|83!895_:fkT:nV!xp#Hb'K-tk'/yb:GfL[!x3~&+%_7:?zw53'B@c)|ovUz(92HCj;UUBC5?VJcF/~y r"H'EDh&>-tEQ$D&;HwYIdt,q"[Czg%|*ks$xB9Zr&p|~K	=Ku>/M3wr|Y2/J)CS{zC~j&4c5U<YQJB~	`h<YeFT#l(~L+zj9V5F9+(*=VTa4Q;w)Ig<`kc~lynEEU1iTq4=VW,?*yRW;6(q;:]lD&KTyU*9Q$06m |JaJ0yfK:~IFe>MH\,UssQJHZ5yHM;1Pfc )	2k~`f!@xKx8;KDKdaS=^p3.(35G05H)zaF)?D>ZRU]7h'hn",%O7-w;q+=JEME
Ni5zmp/B><T2'RiX"|eSKIAR~I4
c*%]%|[|PKQ)x)i3f?.nF
9L1K^a
V5Kq~ O/Kl]VSTBpq--x3E6kt4T@Z58T+;j=SMmzka]c;@pAzJRL
:_GZG&r.J2P#7!Mw0KnE"F]9Qx *duXez=JSW*-Ms)? Y	jQl8S1EA3U+Vf$U5^cgc/?
PV=f0acZ(l2FbAoV7"$u0G&%M/%oli'BWiT^3v(yWMd="Q(cckF(
~-VQfzLLk} x.WKD<b -04uL95-t%t	IH>/ Qh({zxXj*!5n7Nx? vkd6Y8t'5p*AuC=6rWs<i	l,h_.6Zye7HCalj0zQkpbl{dG_m4rq3jXB$$02kwR+&BYzBfwiQu*e@jJa^O/4/iSlg`]m2)W^w6hBDs7iKi0Jo.0tDD3Bo!>n~1[[D J&]\1;<][!YbH K>,NnTT=<?;'6AFdcG8Sr}gp^{2(ii$1iVpfs|n_dHq#S$J DjvE`G:#7thUQMTk.m#u_Z+i_\yR8	_#$c  B8LWKE_06`S.KpK8oLnn1O<$(.h-|hN#paW3ep;Oa`{_Z[b!}O0^yH<gr*_n5nB)NsGRINYcTX26cuQxtHK=7mBUNyE	'0^DsV"q&=2W5=6@}zbwdvhek86;=pp)|X:pE8vW{xcfd+.m1]U9ch'#+0Az@x?uC&_FcUa-vblr?hNSC{;N@dej!wR%5+8_<yH7ZG-%ODt!pUrHVo"7,l}ZZMiRFB*e\%m<;JIc.kpKz0Wm43~;JvP\_6X(LZH\Ea_|?/\c^>7FWCg_	iADk%,"0x$-d77w5^	/6b```f+STppxLG_AU`6cm{*<|G[z*-qE|#i4:L;f.0uxn7O@`^qD0N]}!(N":+,QYb -t!
i@j-wj*6T=
O"]JN`x0T&'qa,@E9c	xB@]hI	MFBvu?Fzgk'
69;\}VI4lRr'8ZBZZ$K@/f0YM8t6 cuuI	j&}Fj8,s9<J|$g4w$SbE\f
~jdT=..[vJ(]a_W@*
+#@RIWuA';z/v)%-4`WF+xL}d-%1r8Zh8["id#7}+K29laN<NHl5uc6r~^~%,/YjoyYoS4L+%>chV?I$}st)
mj5CL0SakJ@2)8aBHzLyf3)zoL/z`~Eue~"s;#d\!LDQ?mfMrqx|`X}J\;jK^T&OEU1o^px*WNqdzHq\ph]7|sB: _R!oG@0F"y^KA)w]+SY;D[
E7!sBjbfu?$R.-{v#b'<:J)`E&zvMXuXc@\<z"M7"qvEW PJ=:	PEH'+s=~f<TJ.'n>1&+^C#QIh%7D@qmxEtC/$R
-MFu'
G^<jWooqG3fILASW^Ge0p*J(02i,|aa;rP<nZy+)MHT&9>-(<rY}c,{-"0?qeOJ) 4e<$yPpXlH2=}3=Z?R(~"Q:F\QqfXtPY.I0snzINdiO]	,6 1'B?Jsl^cHLF9+jGnX_3YL`ZIxkl5W9kPL$N*"INN7B4TNB[| ~X!YOet3TYMkn@*s[[oJw *xP=zy5HSFrT{M\:8kMf
b;Nzcbh<J$"_E*UW#99cKti^
N2a'!MMI!Ip_miDK^e.C; @[AtY*a6au^ 3.f-jYr,]NTJOd	QsS|q$\EH9(ePNPiaB9*Gf~YbcrMa3YR?IAH6=Jz8&y?|b<9Q.7fTPU89,at[DynZ%ko5X]Ict>jfv5rg{Tip0PC5Ru*H2Dlc{5:@tB	Rw?Q[k9RnwHNF1r@pECCO:UTR;tBG!("|8,h+1 h>$jOSD|^9Jj !hm_q\le?8*,oYB4g!wznjlo!y,{"qmtUB+'19:%=Qp[F)gI+L.t^E6v!lj3{=d*zR4,Vd'z5@.mw6%NH#> AXPI^N:h]F,b0"z!5~s"3_=
3R-@?6lQ?+?]hBb]t}~}^9C+h|On!T`M>ATGWyYW*kb1`nlmf`KeE0K.9iyC-;.J<;eBs|qy{b^$4:wKP!8K8'qIk'bqJCg.uy%CZR)8R}#\'.YM:FW@i>[nH310-E,n,iou4+YuyN1%5?"2/gz -hJnJl !3K\1&Ees`S[Q:lo"Fu).OZ.HhQ!<r>2afY^LagQl|TBC%+h;v}u1Tzp^ZKdOjv`+=iCaZ-GhWw|~%p-\8(T~|
PnKaM
Xl?:gQJh-HC	vsLI)+ 1D"1SVj_kEW)XO~%,gX'BA*6&$l>m;2#f:$5LG"J'Ws%$sCp7d3H4+QX#p`T&->4n3=8=X40L<<
JS;Y -*teIC.A6idRe{hzGuotV1DYrE5eX2np0x@90|';c:]/O 5PMvht&cQWnH<[_Yg=gyilT05^%B\0~*;%6]Ty.Byp,K:1Hj0mBl12	rr!8DT@pZZJjB)GMJ`[O~Hz@b|2[+OGZmV|v\T6k=qSwtf79GYkfmF67H9`qv:L7jz6{:R^B@$Bvn7$)h%#3h3ce|a{a79x	1XUf}`9uNfyI<cJ4s7KTt(,ZB@>#oc)|zk][0/g')CevZ5j84wx
;k}eOI+rn3)uXmV*	R57bIWIG6k1`>MWMsGopO%[|zGA>v:=o$j7jqbfroqfP11i,l*#G[7C
8&ByX/pJh7laix2gDR<)w)RupCWHQ}m/aZBdrH$[<x+1FFE<i;.I_r]]N6|/KL@Z+_t:
SWw$_7/7^MBB,(UnnQxtiLz3Wh#?+w)z,,h.xw)yeozix>1xRR~a?U5'q:tr^Cj0HZ}w&ID/n[Q|7jMa!;P41]C}L;2GO<t)1~1O]E/;\6ZV8	ON=aZAcN,4^ktPv13_Z6![].Hl VWPNMX?}y7xij?gt<s2?j+81\uy<M`=~yXxDai]h,79HED.tZ 7:E1wcc$NL-}X*g6`fP9U9mEMw0-xdd^szlEM@oZ=
]mX`
q#)~EVrwBf0>_9 \0C#tg?4Jl<fCfjF5_,|"amZGs}<Sb_cCCQk11KXvkzuO6*)v7M3;a`RDH$*Wg`^8u6+%qv]Ja=hb|hle9BFYMnD{e<>bNS9<,ML[j6Ns]zv-&mVzPg~?GkO.fX/H,tCVWl.8=oP)iP`B}+}2%P6sPP61E8d9\=BxKFk?2{]>EGBo,DT0ni"5,u>A!5}siz$`"YOF2c]<)t";VWOoCkj
?>4RWT4,+_EBMS`%Po0,6?W!7EK"q~IU0.O/>Dze:>,0loXF,^'\"3L%;J^-9D{VF9yKIqY50A/3l*s.L%{JGRy'@{+Vn,gLCDK6%vtRhu0`7w6;Uy,IAfgM={6N(
P;FK9Zq].	_R6$0Srzrs-%.V]Xruv^0/EH,z`"YZeQ__`
OwSurdX%PUlRE?KRo:MY|N%5Tn<W'(b(K0c[
%$^G"9=.OYkf#,|iLc_h.nV4R8QAf6B,Dx2"aA_dyqb)[kT&7<7f2;|xvmDD;:lad%Ualp}B]-{eRhepT:X,pngm-F`F(\fZun=B:=T[]qpR>axQ^c^%T48n	-Nu;>Rfk:Ox*{H]w-Hkn~dR&;SYSrl/^Q~E"Kx|zXXSmIOr;TTCna NWz?1X-n<#J`)688YzBFM{258k]VUUp-__XU
OhD*)dI.:4HAR8a(obR[S%s|Z\L:}s^3xGwt4&?Mz>_JZP$eo=N`zPit%h8,~w	'}rNq>?XMc!2h5?4zf`d|$CsN_$9Z!K^ngXLLNKFgdzPPKjOkd	rmRdfA?V<E.|-x!a38Z+l[KQkd}d|bV f	<$-3 ORf$\vDUJR0k vPtxtix;$m,"F/*L$	6N:ep5fr/6fxfHb7+K3!Qz3J#Ccex$^qWZ$@KnG?EnKf[T^%WD[#9`SCNt1v%[Y'd)gX4(6"}nVChDCEANtHJja)S3}k(HQLfgyagi$6PncIHz[)|nyoI$Op~
*9("a*7>_\PY"Xr>h=""a]^aWg-XBniKnyq'qnc[LdRp=#TLvuE>RpZ,mv~jEX9CHR.nJ7?`YA&sT Nul8'IM3;?fKW	o0<mhx-:e,Kl\2kmVbdg<{Y2Jr_9VR{"008W,
AscoR`{D"2/:Fl6w@c;}wgj'G]Jzt"TwE9?"Yt]HQt.D9!@Y/&BjRgQ3X$h_J@<KYUq(i.kwS%|%1
,/>p4bM:3t#tbuXB-+]|@yr+?YaBs9wec6:[Dk=FTRuwT+|sB_z=&la^V\@U$q~IX4:zTK'}S^A{`/`:uUd
Vf&85ymDvU,6o-b@3 :bw" *>yvm4g^E^@z0{.oj.'=46T2M3 *ka_,K+~RKiB-kAU8r*{s+&lyL8p|]~j#R>6jg"NjP	k/XS`cDm% iV>1fUgF-s{_ACxk@48aO9;b|xQ<} j!3g#HfH^B0s7%0`zD(/'#bVR6e<.)eR:#5sz)(.L$dqM{;2N7i`6||\?xj^`gV'+;_!3F8Sje)"/:C\O(oo[.&DFcJ(ve9Y`">x/8e5|~Lfh![H9+(OokCbREY21,OS]M:ci#[>lZ+z1dzuN~/Kr(Da[TpSfcH1OQjRTf0J#>X\H*R=,dK9|^4oE\}2o8A]'>w<B?xI"1%'EOpm)E!F,p9CUe=LKX'F@-bv]o7DX,+J/JEDgECu:-?dg"_ra8ix%?=32XC6=U=kOT<G2cG](w6|hWi9.y\NsKV-*qJ~)|L5yZ!5luBUsMV#|i[%@"SeRHg5X[+R U\VEa`6:bmpxi0F(25L.U#czyud9KIf<i{ys\K71j+(eYn7KpH1
E9 /tAax^WB:t6%aOG@_Q_i?6SZiCb=7vhG:0g5-5%$\6xTh@i
?_dQAtDCtxp@94tTF(*f`[*[JUq+)9FiCJ;cLeQ
)5nL-)beo!}idg>si	09Y,v&EP_r$DprL.N`zTTZ2}GyH$-}T'bo|w&cYFe{TIz9lw~A3b]{Tx]LqS8<< >;S:XNBzObrf8xvZ.H6}2,_;iz4=p#})e_h'p2FTd2q{XIV;@V,+]5Uh+LLYu+@[ZrtDp|Zft 976 !
3J#gL26+JoeAP!MUC'RM_S?(=J'M?h/WS,*.X2+HGy]xk^Ad[oA#>mVU2`.w_]g3y_Eg/2.AP@Uo:vgR/Ccn<<h_&}Hn)>Jg7x8!c'hGa2o|4`3o$Kq%j$|kS3:wpp;72b%J!^`97FoMjk7,:`<OU;3!lR[BFUlW*-8FYT*\GD)Od@:"-I?i8a^b3Uew7?|11NCV7ke$iK\]I*X{fm GYK?Q"6,gLDU"N{R?2(F^]S.y,g>T8[_A;bUgYP2=}.{/mCP|W_/R^/2=
>/jB&lw`3jlkSnYI,VTmln6#pszu8:SMc `:K`</WV'Qv}zv>[k [9,|ree&.w'OBY6*_}Ndu2/Y2Ox"w+ZFF^\Pqmd:tAY$uCxCBcI,slXv(#Izd)yoSs ,Axv:nmoz:)]GI8@R#9kHc-x~HvjI|E=b*s2*KW2V:T4wL1i	<J`sPA`R1RUpz{j"p#)8l.<pZ40Z_a.ii%Msggeg>EqC:*|%a~Ow4;]\Vh4z4^gpzc,9Adl`hFhi*{2\5L,1gn>?,{+I3X 4D=k% o?iHrTEf,h.h 9D
(!pYQ.`a$+IRhbg-Ji"8%zThWSGr=DJpZCEbx~F3(M
H<.;%%aTq|vBCJ'i0jdB!kT]Ztkc_8x.Nj1P0Gt?f'HB_`h%<A*menL|dYOYc2N2x#vS*%}A"t=PyMXJU,_u+bh6+},t_D2k"$l@ DSP.go+PuQkv46l7;tL<KCKm)JJ"+Q/2ds."l45VHW	9z(Ue2Zj%CmTVt6\o=4>l)"&0AVB\^\P I\md,%$y/nWg[BPtlL0sKDAe5N9cw5-n	#i}!4o(gb{Z0xcS7|X{[jXGI
(q1->X^Ag+5FUa?X.arohP2nUq4jJ-(>)-bA~@h7E(qA0Qoa,F}Xl|j%6:a;^o%42nz7!7NFF%AMDd@	QdWQ\66zG9<:a]+cF7SI]H)'5'T9_*h:hr:*9baZE&4s
7&ge1qfAt)l}eBzWSGv<A|E)9d)u}?I[o/K7!s}<,7mi$mRDah=xGG@^Xf	bq7-/Cwr;mo|15-P)TNp/;[YO;,H.0yN;-PAh']I;mAjhaSk:jR9oZ_K%j_Vt-OdeiypvI2s0uWI3y54+g{,|PTpM|6Md>%AG0=L!9c2i4*UwB]O(Y	z\t`6J{:r#e!k{7:8Zu!g2,/taA2~1sK)}9,.(J_
@%=n}4(Tmb5Ta%VB

sV#ER>4;nH$k]OT_zb `(Xm7`d5qe$/RA#pS5t@2	mO@*F[&UEc&RE0P
9vn)6NM!_{O%E[\:
s`!SgZILcuCQX(OnH50oG0DS~=5vC})Mb`J{>LquqAj$f
U=3_0$[Z*mx&Mtj=HlFSK-M0
MtPO@)N}? ..-%MTv\e1TRInyL/_!;8Q'|!~_[oDC]5aRq+5GmX[<s+
-"s7#oU7D*Z*UY&`M%}^1:5FpIqf`^g2yrZSPeOe'hhVi9CV]Tw~2*Wp$^KQW`;_*!;s.7Y4<ATq >2wNg]oW(V
&>RfQ,h/s("X2rJvcG[I&<aP4	@l"w(S3!O3*2jJ?Q:]&u^(i>ddr"?a-jbujqg4\t`fHrIhgvOJ*K,q2_atZj-;>Iy49";LL10Lp?Ni~~MX(b"y*4<#s`DwX4~+\;jz;TAX!A6 c{Q0UO>_5eVf/<	t4cs-eTo(03">[Gl@<X1Ckq	!<_e3`B"9?)v7vc<,lqKL:<~oz$;#E;+WNVG;1;1+6d(}Ayb|0LvmANU^qoyFL!nPQd@IzJ]}5J@rL'*rykF4Z)<"I"JKX^G?-kBJ;Y*w9?&4{%2odPN.Zka(X%^ea.1 %|:"_9:*y$Q1	u-&e>.MEuti}x	/*:X'Q`>SW#MX>wdM"5|u*g<`"fw@%y*u
,@	ik,#~OR$-5I(	pT7KiZNv+S{[]JS@X5_pHT}ljIfN_]uxtw]-}WP{jaHD
_eHJ&eG]qv}jU ^p]tM+R@OWYRlx[}EXl$0kfq/+JCt9^E[-7XT|FvnI~imA'<tUG6Ku@Zgi6\UqD~gy{l47RdLW/.XWa*OeL'{l,s"d{A<0XIfV5Tm[.I8fk7r$`]c:U|+Z=|z C9j]
}NDnC; D:6&SPFXo=	{`p}d|yI&X4lH:2a
>n-ktrt{ZD,n.@kY%l#Ej_/Z'\A6{IRVNa;0eE?:@S>2![o{&dI"-m3fJ.GF5>PdEx&y+ (cw]RZ=mxhvDa[bn+dwU-Jz@7!xDS19\GEHiIEzau{^S}wo)`&W}?09d85zIUFu$<2DCyL;^U&F`-ek&b_;6lQr^LYQ!@#b8GYYhHMF-BH</'ko&\p(Mg4e{A6v!;kDNAkV+@ {Sgg<^H+L.kXr`%Z1Ym$M{m!boG>dpR6Kjvv)4" -t:~oh[2sMBTaXL4
)gzAz`NL]hVtV7"awfF7?
o!{cf{.R.\:Pl_\5UfEPK9@+f<|G0'	[%>tSEbJvlphsmjA]v&m1[n2.S:]&bn`h]TDT&aL' s_jh	[+~7Jy%[gHDi}P`iJnf[!8?P`/n208RV1ed1+|C@i~brCa>/*`}g%e}&:ihHn!R|V%}uGo{5v$~d=IBjEMp-x?bUr?H u7*.[3N\5P\}{<R+'|\}!__PMmn-C+-Iqp*^5iVnv$Hg^.U%s}M*QiaJ)UD*b2`k3-8Q-eGEXr=c0etDFvh*/I?c	 4Mf'm-W^ldBjla.p!'Wp8*HptQ<t~,tl+fwmyW<rOIL8ye| ]<mfY{2D?DP=i]C] 1Y5_h"1!o_gu[V&n!2V.x~O6MP2h}9j9Oa0[q]da`q|#3=&E(:z)5s]8C@~ ub\wu#f_ANlE{:S%K@4p2t7 v`,6cC7-oPTs8p;M0w5l%:|nb!S->q^NZ]8=}:2	FdzLCC:sfji5^eU1wi-YPnxRQ"vuJey"zOPDw:7+bt!h_>d2IE.{ZK"Fi]MTu;{opZcJYOz;`(y;[ho<Qs%:eho7C\Q`	(h/-u+}ch>}dhfx)N8}D`+igIso}Qj YVQZx)stEN1{"Z5=#kqa.>N9;5B}ZvW#0C{B_AAK&F'!X3[l)l}{gigtyZTY@Ag}Mz;i&PSSa,L$F9!eN=G8R}pxV/+uqLq=}c;.38i%e>yTH;5H;Z4f.q{Q6%2m2AUS6^H+{x7x!99'>WBW&%H/JLy}9,X}-}j?+=',Zu;p}L^2)OGz*7|=G
ic!lEw'gm*e,v,sQPNdLxtv#2j<@ucKRkM>8 5_:(	<'+$CEe|JHAw9G>?@)YywvR.Uz9)4UPHd~>SQmMCpJkWcad+Fasb])ZB<:{d{2}>aUR8xf rQJ+_Mt1zUxRt=>o2qbcdbkuMTboX$).w(q2zL,r~3qY~z<	|/u3[Java3[q:+in lf/ts3dN<O}(;'SD2*J+:kJM5-)shS[Je>S<"|4uq'[kH~@TuUGQ?S|2B1aj_t>xpSG'	XS:7Rb/kj2oJ=
uG_JlcSbozJg7}_aU(n_OF{px6\9Nx,?R:Ne492~=6%thDK:YBNf%oyhaHk *9{uD(k53u0(pFuxu|#t,@]"i1,oWW @rYl#m|QM;i};JLlOHyM6:`H<;lfH0&4FN/'[nTb9S[(l8ceYg^"XaIiL"J$m!17I.*/
s+ %5g1eJ>v>1dyb})CW]K:,b:*\ =qgQ}j!+mBW_:q_aQj(IErV!#*azq-UG}Df4skf1VQ	KU"9W[knB+:jBBH^$9a-x2p3C9>vS<n'%?mS?GD_8G4gj#m2L#e=|`1AbgPwKXqPzL]z/%H@$I{nfPIz+(p'c)L1x"m9;&x14FNT}e$h--}s6Z!t+zdfhT}Uw0e.#zq
W43aeVX{DDe;MM<|G):6Uiwq{\.8h,58M$tD2y;f=r-u3c$0*J`FhDUA\q	TPr`L$>j0x
Wz}1(Q{\6vl4oM\ah'$$0M2ktSj63MAK:V_I1"1'RZt1yGz_<KWA6//]sTyb(&JjJp	WoTw[F]O|g{maRUDHb@gjtSMr{FV
f1Fd?SWk	lpsXBB34 B/Pq:$[b9`(wF[DG].-p@HR:tWc}vyZ'ru82bK|r{E?\0C/z~RKO^N?SQ>J-`a/P~vT}1`pD7LATm{#i%n;{e?z%SJh/SJDBql)TT_1'UcKgQ|zJP
KelfOar"P&u7x	x,bD{096M)Twov#
	.]"bYNCXgbFEn,,
ChnL2@;gv w/q0tW
nUQsQNZP8,_y1)qW	\M8Ha$y[}?3W<yv@;i55<<y+To*,	@:]ovnhBT@$Wa*10Ue-(:bO8=opE=({:_7J
k!ZbNLWE
Cks.XhTi+9G:h9VLP4Yg)4@t|	=,,0JDJi4:Q4B'5_owH&2W	z"; )wG$[PT*n9v2zaS#32nTgR
liuUy;y5Sy5*".w? )>)(hb$bi1^\F<#+/jEIUWGS-WbemUdwL[+wUPXB@HXCGpgu|_(v%C/:w1ra9*zc"O`cBHKa"|8ePE5saNd`5uXZ]'c-&KE!vY]!OJ0}tIWDo t\s"+jw[BUkSv96cDkm%0*d~qe7
hr'ux`)ho=!gyNE0>fJ>7m8l%IdBvol=Z"vaFcH	xw^Cszg[=,J#_=ISKbR'g=hbv2T	(LMES]77*8g'rM|S [TgMS?'1?uckanwUijr}uMrs&SHRl5 $5U{?L(t\nWog	ZrwL$Iu(+9h%#l"1HhL?CEqVC92lCAsxS/]CCTlE#2*c_qp,1lEzX:oSSU2]O%msNzbT"uo*R]a'*n>LzF,D\	0Z$4AnDBw|OrW6v~PE*P7V!FtKmjTllyBK4`PI[O6f,Z3HSo%N-GVPk8kKr_\ViX.m4`lhgUy	\fwPi(@0!R.g>cK#|vdQC<vxj+m]+ DS:!.eHWkdwl;(6p,>2.U)(mC;Mm+!4hFuc.[`$'Px#V:FndEs(24n3x^ w\7.M,U/'l_w2}XF`9D'8lbK*xC^Pnn(J"rmv.V?T8$d
7{s|P1ULzpLA+(A m()b$t~\'H,>!MRw+VNQmAefeP-39+hd\f4_m>Tr$2=[yVW^Yf
jxgB0nLoZUi&x@=	STl4ftngJmG{L*f=>Z2kb.**Nm8;O@tFH/5A0&P1`=i mi8',}.3/Et% E;0sy+_GP17rYr@\4V)UbG9JijGSmSg"
IJ(=nX'LV+_FiS~{5g`@Hxs47B0,n6!i<^sq$]z9sWumPgf'L!YfWWkS,QLrr2OI+e K`0o%C=aJ0^!wcu&C `<l
Ajlj>^}Yzn8<qCz%lHu?6Gz]qwfY#enYiQUF~um$&XKNkEMU1H<Q'HvaDUZc%13#/;;83sB`:J?+HCk)H?Fg
+j37~(yP3-n{JH>DShwJ$us;#dz:4I[*pd|gBGVmyfLEeY5V9sjY~&Dm,j_<O	*=k	C%tR~!Hz%YsKX~sgnB)9%ubGUbP[8b%=Per*l9 t2=@B_;Zi3AYi5lY;#@(K'+7g+!G H^y?]x=.tq $pDx/r:r[)C^^v@h:0!qA.kf8n>*nR )6ZXsM'{_N@y)rJD`KKhe6|tdp&Rnx0]o*Bfd3:pjV.9!l<@Gt#&!HQV@sI|\1*eh^~<AAo5:L5-?cXi0c|u:h&?uHxg>BCCb+Jea70N!4z2%R9h/7~_	#=:Cb5%LqQ(Etv\, xVEU[HhyBHD6^p$*k".>QP=LM-LMRAeV _"6g3dxb|+l3[<E%x3C'-P3jY9set1!ivUnN7>"[}G0#ioE;bN_WF{DL#!+azlr@5gT.^*aM@#,x
W?Bv<x^LhDE12X")RtW&UPd_
21nL||QZ%C*s:ZTQ9/lpP)J9a+zq|Cs}+(2Ub*s JzZFd!Kj[=oD]'f'q5@(U-nf+FU:Ti9lbvbEg0	XHjQDVWTg%c6$a2>c,PW
7h~1<c7$6!0&L8B`V\#V1{\n\#i]"-L=bJ-|6Dy4~N/Cppw<gzq]|d"_a|	U7YG3a]Gccs9>-l)r4$rAPWf=~=)L!$r-[yBOAkO>#CE6E.r7Vkai"z6?q19]B:%Gd0:MZnLY]Km`=>!dyLT(	QHI9JJ.-!N&vi_EX|)=>;|(Y~z{yb<Ol;pOVlUQ!*aHiXNp?u(O{F9SWD<nFg+:j231qLmAx2_dW4V%V	zu}5x'kD207ykr.Gu8R5+^SDKm2<>%2K|bLEY!=H_1evd0h.Y7pP3/.Z]6g\#9	},(#}wXa4[ixPu';aOW @dW}<	REB1OE-+a<{TiW%4n}	E<xn6}jY=
vcp)(/O#<UC.r2.i4\ R1vc	p\^DFU=Tgh&gqEOH`5!Yjm/-lmx-e[yRJiqa/*>X& A g@EIY,hU1@FdKedZ~cyw*GT8-lS"WpbTFw~"}v\ &*fp.TRmYXFlYDx!`/;+yx ]&`6P]8Nroh7]~NxY[H_H
eo%6{%qhDS!rALzV!:*:Rf&g-V\n=J$Oy?E0JMd~JK>*5`I@c@}k8g3'bRPWEvRY?W;1AvfEJ9+	)M@}:{L	B#Y*/%04kR*#Y)mc0q^P01H6y]5'gcO!&m29,E5`6lioa2o+eR:hmw9X!
,IW7.;[e+H3:"B~I*9&yc9dzb~r<j\[A<AfnQat9ks[0rB[$H@vMa*t2q@Ie{;9g0knJxe/MKZh(W.U`=YD$dK[}`n'<5rt,=r$LA723L{y[*,UoAl\{As&Qp_+f*/>Iud(XE'Fsfd8FVij/}LAz1fFWh=4f$/}t9(E24VUV_>I0X,_Hd9(njrTzYF=1kwu`]x
Gb(@}L(Xc,RMs_21-SHvK&|HL^VXh4QSw{%={)S\ }O iUMC;-mIu:Ule\kt8h^hR{pMoo@jy{*cq 2PLKye[@]~MoG|((Br!CS~K*lkwI.{$ukSBEh]Nq"nfTSGfc.gm'^2fsaLN0#}&%:T%["n:B=
"3 &OA!w( \kA(-
}mPCq5+B"2rX{~I(6{0Ah	.3Y#}OJ9_tE$RE,:KXWCL
ZcJT&rL<tDc<"'|3]-5)RUz2eJ4'a=R/HB?r@_}FIoK0D3<6^A'UX3m4FZ+a*bQA&hqnCg3M0CWU0gW1/r9!2L"5mSsWYj2e(o0ymL:;Z#*r*..
%-pH#T*vmdzLya_mfk.rU+@SYqo[6]q:e?y$3k[h8+!hIhyVrJ slACN?aZ#QXu3k'meBQ]>'b%q?;o3fU!i-J!W:MUzG$P`Ioofd@~',Ekqzij:jt3rI^\P' J"|f!"t,0	yFhii	:}1mWGgUA-.NgO xN/&m$SwFUX7Uk2<Wy	A8r^)miTFJ-a>zYI|~%,gq7&.Pb:kd&l-gCF3!^25e\,67.U	<aR0fA]I}u?D9]&#bylTf'^*i*cq~{8sZgKfWl2Sx@[o99(yB.xdR_m -.aC.Mj-D#`7
AH`9tQ][=R@S}3&M7MkKofBqh(px-hK$qS&:)8\R+>o1sg9Nr8@Mp#6R6Y!\c*B9!eyqxe!6(dQUFXp8\jAZRz),1Ldy<;|`59Y9O6RlHW~dN?kHZJ2ehq_6B	PXH@`I[Ba61of-8sAsi(.1* pu%~u88 !-y(9,2:59~PU9((i#yh6rPsX~/PCX	
1R<c2,b,HKs|Q_{5=7jLI"*f4(`6M32J9'k0[C_CtXX]x-ts"),!nqgS>%Z"<Fdt=1OVW*89YBc@$y	vx'.nVMN:~6wDY$25o\6\$*HFB9c4	Ko?rAF.;9j=W}8W`R9:]{ehtM~W'x<rd7u*I|.;Fv58>8@P,@^qSiy`0)Dj\;cJx Ib$Q@GYP$Giw00CANG77G:oJ,Jhq]?6pl)/MrR@7&\Oht!uu&+)D
%3f=uN{NtW`IA`+
-'*v(y|Jf4YN](H7G+kO)%#WPaP(!ri`}r	UGcP^&Tj>bj\!j|4fkFDbLA6ln^F q*m"C7/a?(*fPs4I8J8t|GLu+9u~WOpjfS4`Qw=7as1b*>>hwgjW@oE3pGDcF&LCSp*H7k3uXd}2;HJGn=Lc_FvDe;9&Q5QOX& pv*I6"l,{026ehI%CJq/+QH?@#[{4DrI_%L/H&vTL51yRf>7i+rlg$~9c V'WSNWsp@f
2VXovw9{	sdu$eL["=M<0!]u:4Z>!hU('x)>k2E"p1/jczoO
t9XFP:lvuY+Ap9E9FtTpGN0E1s	Jsy[sv1WD7wq1lG6Ry//=_Cc?6?>DH.R|$'$C:Lh6,Axk}GIww*}U^#.CTAE\Zmt10n*O"hc	zk$mo7iq#?3+WnnnL"^,B!zp"=S7a(&JeZz>-, aw=3fml2D/'\f_xINquisFOgOQk%6
!_HTgO3J4:'hb4?}.X
POmofnfF$U3|q~3K.Cli%']uQ6eSt]T#?ab~->\<9nz"Ss&OYmPSKNqZbVj
|R}b3;1<YYVB*4!>ss%Di#;[<-}2?U^*88E=7	-V0~c+K,%(]FPhQpfLB"f'`V CU6vQ>b0f6ygKf{i84ju;KBM?TJ>'/dG15&T^.7XH*) *r^Gir ">#i?<)Dy<A}Mm'gI2u$-yfP\T&dj'0]r>a xG":8p''GioY.F_
ek= \ZU&[tX.qpRk^|G\Oy(]Wk9MF$j369VU`"1s'1beOaCJ^OUs^Iu:7N>>tci/3
:mG(~U0e|qi"`xt4/
Co_]PCM9nmE;pp<m4^]>.Q:c[]#,;CqN&FWwuyX/UQ+XjYvnES
>0p^; _0Yx[4r\
|V^!r?jIVxL>W:GwxChe|,"vXmKO.g$eP#Sx-nO)Bq(*#AmI{HlxrYEEu/E+HTE5?F<W3o2=b]w$O>3v.WCqR2U_!mi*=3u}.nx.4|[OkT	uiVLp|;L_CT=S8|R_w)4,#3<%&nJX1:OwX"Ud3~gG~:#<J*)u7gr}JB`R8i"i.{RKyVFWM-J\ZYG0![4{c	7|1<($GR5n/&d30"3Vu6V5G3]ov,k2TT~%*Csamqh=j2z0,3YVA`
]w0X IaSGnBr!S^,%Dy|w6bvRu5d[*C&--.<Yx	s0L-AqXXbI*g	0_DSOl,CK2'1'(b
'YM.|
73%yyi<y#f\Q6xxoFZ9Xi(Hy8$K|NxkHO3r
UH#Y9vi,f-1iFNkR$Q_WLCi1zBeq]k:mX/MJth7A%cx"k;g~cz91nWeO+K% ,"X&sF[1$anZS"Wl-nf-O]!U*.A\u'P|iWE|uS,0LF/sEmKY=vV7){^A!UVKe Y_-?UdwP
=<)h==vB1l'R-j-XVh\pbZ,6^8	Mx|iS848L=P9Teca>L9FiPe*#t[YH9$[-3 /nT9EfY<i^"1,(Q<$K j=IJgimq\)TvT0ZWp@.:Homv0SG3}Von1Hs[Z9^`8L}Di8pIq.{Z^15OZ5 oQ4L6>`!5}*5!hpv0+8&x?8r>3,E3zX?C4[Bo6#X#3T3AQ;^&|	j%7}_r4o o=%8/6-B\ZQ	?"==.g6NZah1]cp*|fQb_{%6a.o9y`Y0eh'VkrR^"kTDwY&h,>l^p1?El-</TqlL~g3sq
Jc-TbJc0-Gb}09=) 9( dK"3Cq?7ul_"4$^vY?Eo#8N;f]MQ?{S]{^R<C2bk;(=_B/Wn!bIK?RPkK6:'{rnV>Nk96%e-cn:)A)KQB Q%"F|\s/dl_ 84Tyl< 38fNM3sJr
uG0hK8uut'thL?UkxZFG5%6T/Ymvnm5$*KRC*!zH<9	Eux?66OlozOBeQxaE.)titHcq
WQq_o\+7p_'4|r868
~^&#LnR2qO|=rYLR\|zXI:j?uuWsG1q4x`C:=p$~}~y$Bp1yUyX|W0-^|Kn Od:7	0h>Se,jn&J*Z+%jfI3KF^]_3vo.Qjo29P(PI(@vK-qVH,,cpcPWpwnx92#zUBwk'KM~4LWR=;eJy0/]+V>C!}a2z
niCDfirE:~9d%:v*Hz=l6jIfZ)NH(L'j?&B9pKWFdx;lo@kUwFx[,2p	 L5Qz>yL"NRMc+%0L8G$/E]uB+6Vw6Z_Q*ahxI\Ek(&K`nV}=h^Lk_ckF#cS"4m~DgHyBLAVpe2Dm"IEHF4*jq-pH858LQD[W-R/8~<kSEytAH8wjKd,LF#	sP
5W(qZ#Ddi+U"5Q{Em-=	F3ALbf9F7sd**x#|y\X1<MCioa-h9hk?{g*\aa5aP>CtfuaXt^E:B0]f!x^5mK]n}{e	X8;S}PV'am\tv`z0TiO`>uHIL{vUVc.)hO7?r@E{Q+4b,>,k}Ul5kzhu6cb2Amy-F;gzNx//3k!p_91R4Q!2<k@bXf/=.\jb9XLZoMAywIU{v|{5!,A/R*Z4gO 1}/x;QTB
(WW<:P?%wkmP[GxTk9V+|pROEb]HpkN@y;?W^7mG`Jt9QQp,2dY&1#[gs7gX-Pf=Nf:`!mlrBv{LOb#u<2'.jmd;S'2);O6f+:'uf~iHqCizR9]rY(w{2OE4EV!*yE /*^}N8u%R`l^B]km&|/ngvS%kSTJ3L>ENWf|O98W	G(qBXF5;DMUQCO{eMui]HUb-XkK
HVNm!B1dicQ~u
; lT_euuPdG*$2[S^{}Z3u0z^	z`ggz_F	oi.xQgTvB5Yp#%"a
!?	W/HoZ<;C<BRo?JC_"}P-b	gpu^XNKb<C'4b9gG#P'4%O2`l4f$Wcro BI*x!QYTK(dXwt:" |wSC={:+1{	o!4d27Y9Xe4l)^i8Q?R.o(B!;x0,!r|z&56sUWwG\58bkz"(s?[[$\$W8k}SZtyu)^u@v-vv"EMyZHBDO->=$g@S'[*7T<`2WlV!6R:I#`$%Wc=0mK[)#;h}j}Je;@0V^R?coJ#bV{LFF2~{ydz>NvXl)N<:W^K`g:T"BP[;6d*re+{V#(WN/R4VNI*kSM(ra$[ 7,'E%9I2<3a[1Ql>kar^NaOE\5iv$tm?M/D3 <6Yj^G$sJ<BjjvxAwa|O9nt@*N9Fgn`/pS(3ho95fK?ltpaF#,<|'jP1B4AP3bFIRs5r,~0R<g	cVfY?G:zB	q_>pLb-HWizPS;Z1JxL1.E5c:59Lo.jF}QY~5qLsko.*	dgy|'qdVx-L[xHp~.g9b^r9z.s2 CE#a29i
&o VL4^ +kn=E63/9C}\-j	[5HPoGDs@j	7+tXZwr&A4AH^C`*=D+Y`ap)n*}'dr}g.V7=[n6cNas|*%V	@qs\[?KK8K 4.,	kY#|*_pt%5S:zdAY/(@<]cP=>5%(vgJO;W8s\}5C3%kB'/bOJIQkWxm_7njr0(!U+;4Lw
4S%{=7p+hs]7#vrIHn_sQx1$6xuhy=l2dtJPFS3&>=qq|E5X0LX2-?hc5TY[`ZafJj!6e&h\pR0{r+E2a\.oA}fgk@f CCUa`r!osq0\bm<4,V7iq2]c4'12mhahj
5i#@:uaJ2k5V#92.]a	%Z:opB%rMV9,nf]f2WWpq4FEj&2bLy)QV:PdFa94lYNy?u+iTaPc.4n?c?$c5%U7^oi>Os_:*<Ks\vuwV@h/x`Y{mf{mjn8OVbvehs`C+su 'v/\Z2vkOO^kg-|@&;<Lo"odv?4m!eHwM}
5F[/Zlvn3?i*Dziu #t=RH;OI+@s#~eB&UZdCU(i	PVze F$}/(;wG)	Q8Q9}zW+hD"^,V(Sr9BOA"	_p9S^UK<e0@_Pe59(^F<jU+pj	3[VA8/"~eWM[ zE[,5zV|^F+vO=ec".=YFK~F&4SuK|cf
)bbte_KWMs5$:aR=+G2lDm1")_?D^ `mBj82EP!n<_Hsg/7B}ea]1
|7uz'p#fl^4/|}tc9hprp1?#N!\h^"rH%''JjF0b63qJP@(ZY;Hvnl1.#Y#NV;4dQ%gqKNXwl8SuMXLW	WRr9CU/?;QqQ$kYuHy{$s"rT`Nh[,0=-z2`^YBS 6'NhT:?p%Ou  U5>l$Y`pgKODl~|?Q=w4v|bx'FI3gZ}"?JJ3@%
/3uQ6
z_u)+%,VU
Dliaz$MH+8/A#c]7?S[V?t'!9gb,@u]al5QE+I=bgbZnY3X4$tV'6_+>(Mj+MtyM$$Dr):2EecgEya_(DH&/d*b>$?`i)n8Go*ap+yz:~kue2"ZOUdI:)I0(1BnSM@w&O;B!CK	v7.PZq?*K"+]x3w\}PzwxQ
1f!T?G*S\Tc.J/h`kO#zDyKebN=?*w+]#Eo,AY;YbFIG"r#?eE:C..X
d^pC/N(Kf*l2Is{r<-[G5[]SX=@N`DsnPJpyU^gFLTo0K:.	<1d]23}?kBr+$}Y(fKZcZaMA
^l7W9y`rX[Sh/;x?;Ikp}=JDF@<r?)X_`4g.xwovwNC(U/2>{2.(QYtjo0*<PKx7Z)4;qSxE(?<Ai0%Iyi;TO2[WWfw(xY}6<"TFN#KU`=61P?5GE#$$LZLZze3gCBm%CM5/r9l!,Y~|JH$_U)oS2IhC=JMb7ldL<Qej{	_"BZ^Wg7+*3mll$\NoNi@@7y"Tkc^+W~%_XkD)%w@c{D]bo1r6]3~|`%3vi"lcmtARMR9YLt\*|'P,&*MJi2*}\T_?zrv
9Q]	J[Wk~KtDrl%zIR	nE;k<zyP1-=!jY`oS3+n[Cfm'r(r]+m\Lk0Y0C!R-NyS)9KWj;I[oB{!Z~=_o,GT?~(M1@%G@=(cY+l5=+0?!de g}`_yhBtQ=(GJl3]m)1pJP}1g7@wEZ%$B	=(fZ&?y`+};Hzig.q"63mK,QG{m.yAsJ~J;&nmIMn\~I2T"PgYD->	3z(!GWPg<-2
7`uP
c5M=VX<4DySdxwsD0bZnVS+f'."-'kSRC4 kv4eZ;}-Jcf*53Yc/sQIO{br*v3Dr'G}r_##Ts[y&{hH6Ly7J7_WU)XU<bGAzXG"<}#A@V(I(ug\%k+65>ck*EN>{pp!8t*9[AA;{{7orWWz"/Q8
SRY[_p1&n[mrhv{S<N1hp!qa+oYSI'o_2CU&b o2UA6FaBDB]7U8|8N EB4Hm6e042-/6we+);WC!p(ag.O~V5#3(QnQesW,Kd4PJX|fG| S@c]DHOb)~-S_SpVT)'FVe$am-A(0$5:"jc#	p;EF#u_yV2V,8bhcRQS>[T8]63M@6eGv--83neMK	Wlt$<MK 8q#XjT3tw8G.R4
r
z t$ `aa(qDr6n	ljyFLn%ih(Tbw4wsLf*|6tw6q+^D(jQT/sw+Sx*%sPm5%Z:,IKduY[ ;opPNV0c$ R=i#m+pc85s&WU[YF=ovUt)Yx]#\lvYa5>ld)9,#IE?lM$,5%<;MYi m6Fj@b[G+D5M\+g)zN\U%lM6_xL1idyjUBmu/fTJdRyHBUEM`u%#\0c}n`(I7(K	Q7cl7rD`vYZ_7`+Lmu\CDQtIsD;Zlbq	u^@a_n5_keMt4XJ&$B(/L\(wWM<\4um.P1BG>&wq-|P_GF&%.bJ[vUG[:-yswk?(4o%wT%jD/ _}3r`b)a.LfS:+ou@Mwvgq7AEhs;'>s!0fUZ=FsWrqaS>Nc7KZ]\,+I|	,dcE57Ppc1)4eYPEUQnbXV9$aufec[{%#85mq`N5aVO=XeOF.%W5$#H4ACet9[sf@w'`QeQr:qC[,oWy|_Tk'k`(&%WDx1Np]X[5z!RS?$B+%#mcuHhwn
?LzA^/j`l_
rH=5C 5C&MLw+dzMnmZ6%fYtJZPugV"7 )=No|n,5cH/ wZbC\VUreCvN&wK"PzZJ%,OIaLtdQbAa!htA4;:~@z?bZ#-q+sV!G:J:f<]>GYR-Bjl@nF"w*.Si
f5$VXA;NP=KUagk,='6fnhV}+r!#C4,@!~\,yZYWOGA]m&	By'5li 
;y+_C+Vxf=(P3^=Xu(>uTD\lXv:RM/UFUd'q?_[e` v!RoYU\nq]7p&;0a8Q=m4`>]3y!4 o.H.-2^F	Rn7{)HRijl|	8bb:ex,>F~i>FZEgKSN4VcKbu<c(7-"J2Ql6`8"&uW;k(<m4pt#	D]W=Olf2JR|LHJPns9P=lMad,"]^35xw|jNZZhPL^m97@d\p6/"qhYP`JGPL@820{K)Hf?
/	y{t?2r<Fj%/0I|kS?!I'@hE3Vx#6a37n=o|A!yoId[^<-[L["<V*vyusInIJ6D</$_)|5VxR4xM.@'SKea$y#	Z{R7S3\vk$Dv(PZ[+69Gb[5.lIO+*Os{1%]Z"7\&`&3dQ;(11>NzYcwj6H9,?y7e>|soT_A(U)z1802/F2jI:2b3/]ghDB>)D?%\Xz*s:K^_@y5 9H4'Y5FjX+A-5g0ny$-)Hp>6pOc\B57X{Bf@W@,d5*<=|tjB,)A|Q3o>woHsfm9?+y$huE8stTmE-FRrG4O^Hw~]Q765CK!?C>CZY\zEnjiY_6j^#|DO%Gb4EWW	cZ##p\w5[Ar4X,^Y9V:!y^c$w6TZ2:-Y#]dr2RPD=iTY%u"={oc_2y<`-k%$*{
[,eXtPzhV;W6n+6)C*+-	R*](	8F!BVY>d`QOx.Dh!%zZ+vCl;:8!l{@	~T,:6|99zPY?(?Ul490,:,Vs$a|@XjHcG90=}ta>T^eO)SPLH>mCC3-6FOuLUq~gs?]`WHu|=*}:%Rjxu#QoSw2<RmA<FAIn_U`F5\ZC-7RjBqNRa;	\FVI|gMa,)_msl/,|_M>7c2'ZltZ!wpS-,Wdk[MFE&QN2j9Aj(H^-5EVrLV@$1k^7N#uEf5*g/V_Y< [p=1NiR1Rnnr/ocm_myF)qtp<q:nwV-dHu4cnXem&4	&g;mBU}k<3K!u'f-BNH081*P"P2	7z?lczbPa\mlP&C&UH5'Utf/?w9Qx*l><HsE$Z+7&M')R+!T66t?$w/r^Lx-H1
eRpmWqK:OA;RX[-X/fo~4&vP&wK>ZPwwqyE+0MKpO..F"RE:jPB0K-n4cP-gc3%n2S(?d.t_om<@5
<&v>H	/M7%.#Cl$q1|GhYUI>s!7UrY=XhWY6o:~"y)[ 6{B,N25LNYstO\AJQGo8@RI$O`}1b/-&2_r^AKYaPz/#7:>F)qsNwXb$7beNEX%:i}sPE[nDA\Lr,be7Z\Tc7CB);JE!ii_rNZkg7F+NSkKL*+^l^Dze^|dkL*k@.m]5OWVBm_u}PxqjfT~a\wYDBPT0q{;SUn4.d[KEjw!aoW;:0/KXqU\lX?Wm,$QPS24:#mE2IPw=$UPj]]^-eR)IT~u/oPqfjd|/,:<)H#6D}t5ri|Uw>v4==9~<%KvX$:>kGLjZ>g|XW	@!Ibc/j#4w&Hbkit@sR[	u:6nWAMl+?7QM3/Q6^@c)cnWq1\D/\qu+W|(,palJc2kI3Qc6vb)L;a cx6+UL<vh0glPg`^'zz}kps.Zl=&	3h<M3gvm*yRqj\YQosQxQ%? nIC+M;
-q^c,$xRdge[kXLw;F ?c/4	.!$KkbbRh!]Yho<82za|]7+t:`uCfF7QbRZcx7ozssGyA"9xI&:1&^e:rcDVu?yy9-`7"dB3k`YMn;Be-hvnWAL0L$fn,A7Y(6VQP\uL$_#|06B"rnN~B'Gtofm^SUWH(JALU
vEe+6]m-U]\)5k3SMy"]PP*C/A]A6:"Zc6<&a@|km	0&1eMp\<ej^1vfD<nSJs-|LLf/DlcG!.?JROE>z0b+TOmws.PX@^~jn9Z4.f}]_b?yX(I.sr$
q6]*b	y"a%;'7GR!1RQ#;kp_3>z[)8XHD|D#`v&JQN&PFEqt	@pi]V(u5o.uQ8'1:
6
=+?]C;-Yl.:H|I\Fbo]d'@\'dY0l#-&5D,2JJ2z[SEFc
w<DDSo&Ybk"HU?ihs<qz1{@v~,VnBai<B%-!yam:&coXX(E/s+R8ZQxPVY.>V		&}8~J+@tKH|F'>.]LCI=0P.5~b`u\:y.NVM,$^nqL:?:,}isGVTwr/`oqWeuZXu6*bY{iT"{;NCO=]t&XH?RuImf[Z:;IuV__X;V>>\"BQ/K4*5E8J\\E4!%\&/O;G^%!1=}%O2pko$^5)}]+~r*qPfYf#8Mu-j.0c,pgpxfgtwt5RuUozF+-X|E)M|OvK\1G9t	%~@IOfw)V $[<xxgFv'Dmv$Vd)R>(SE;[]obp8LH(TDm%m~g2mX/YHR7YBrXk
356&[1QBx,:izi!'des,WRhm-\g/xd:l(y\{~=Z,&VBr<$^lI]W\qq/zWQVH<CE)%G`;Rzxy	^5\P#"I9
FW)=43uJ),Un*M_-s]~]KHMlkJL^no8rCo!EM/!=b	k[1/Fl|g>k6]n-
lZW
UmIFi6l?X;BINKRO<dda0v/J#_@W:63rs5WP(V*}{:2xj"Nof6.B*+wF_c-r
/#}k sW*9$_IVjKpV5%XYvW['Q9JU:h$\2!UWqtxowW01sIrKxI?3j)|j)YgvvO:,`.qcsJ/Zyd8e
y{iz$_;%?k;K7i
@Y..>U>G)/m'Euf{@ FUOAeT=J-=B~WN<1qqdOuF"Rc67 zQ=vs_U<Y*0x1<]]akY?`--:RVqfQ?m-D-}3T^K5NDpew.VvGv9L3X?vd"Y+T7,hDFUAF{a(t@Z[Yy+<-3&x"X`jXdh^X@"Mxv},]9n<NFEdgV<DZpMVg4@dl2zRpdZriE#QX7pdDYW0P72vRO*`\FM2Zc1CfG?N1	;D6#iwySkC\ K]2lY+e:u#yMH.!e_@1LM3jN,\q4Mo;"	8n=E{SP#uAZ5EN0WY_DQ"JM@)Jo]m-?<w|g:vl6D.#U%v3sRhEjf|g7o;]U<gT^UmL\geHDi:C	8&r_KwiOqV^N9RJ{]A(5Hc{njf^idub``i-T~^fy|f@9Dg/,1Y'uO"qR
P0QQ,TK,upI6`4 |K8c9k7yLexmelz;<o8+(6tf;wuWw+Am}2-d
FHb>]A]X'A	F\Z+~cE`t]q,/_I\M/_*SqVcwYNn]f;_K1xJ4j0}7yXVtX:_8
KxA*$Il\X,gAdy`(|y!y^DN*?#GM_"wOY[@X/i7\D[rOSlsRcg+Z3H-GaUnp@q>X8\X83AlqB!EiJB3	ynU$c3FoEh>t~~`Yh5Fl?dWNPM56?*k.&Fp3jlD5>O2"9x~x	u@M	?HY,7yG'/Tx_rV@;FCXT+$4d6Iy&9M$jo<wOwGGK/{o'3&~g1nz~G19ML44JLZZq41C,BFmg}0)o=f2V|[F\EDgnS'iJP_N< V,Bb!XVUVz+P;w[VA*ozNSS[O6M0QqY-B"^Y#UF0hi`MgAZvW~EkUp19YiIAu0[XI&T	r+<#z!MkbUgc\ciehg=l*@5Z=>\5(U!qktNddy^Sd+U
m7U"'^^1c	g(",e,yHm!Mr;g3X)DzL|h4L9=X3/v}0Q-IvW `v2)#r	(q
;pI_^;h4~#Rfy#SM}a"02GPj"YM#9Y3U`p!>M%58[!@GE4s%,E!cxO";{9zD{/\:LyDtT|	:Kb,yYl&	H
'D&1Bs5}=[Kk%DEG:0'ez[XD#X2B4~e\F33N[[I]+X

IHrp+
|6W5/76LZ{9;P=T,Nc'^plu2e2
[N\'mR{5_yxjw)tgO{3Vxl
wX<_6Sli_?OP|y|#FxNa(XoE8*fXep)hcjL#bi*>?+4^|:FCs-Wz009GcK(Z?L9lJRbh+Q$6i+z$d3&;GH)ZbpjadxMAzk|5bb)n{2dP&ik|NjQ(0	Np'.>n@	hRa@hXxXr5Q
8^hn	<\,hl 0Ck|bC(;e(\;#) $Zo/9c$^\)$Ikj`UO8Q}@jkgWsuK\kZ9D!,/opt`t`^t~c#t.[U0W5k]S4<7j&mn|5*F?siw%^iL.H}:hg6O(9buX'B[%U7)-7~\:9Vj	EgwZ2Ney%rG]fW'j}@,q;z4
e#pBS5C>`4lFO&9Z
Ug%$`]G>hl[;GA
h1]PAoB,yfiDyvc8wI@Un8Nt	d.
rwE+=;,WL]=>B%o!Ar'!M%PbBG&BJ~4+WxZeQ{b$3T6Hy
Xu<2%d-Ro9GQCnI|Ze]K0M{
xMaGFb[X.\rI,UzqV9;*yaPIci,u0mTfs*9*\2=+!.P; fw *Db?\'beb
q9CdJUi0<&Z86		Bw\Tw)HRvY6?Ov&SA*hCr{{w`\hwB[Z[	59B=_NzDR.`D%{M	CXLxhLUE^&de{ -E`#:,c3tr;mO8 ,zrMd1NBK
( ai]
P@Kmp
mCJ8X]>,xO$S=SEwH2@CH"o76.1?d:tMVe7FmZt;$I
i;%%5{up6{D\ZB< k4ejbfn"OVQvI@+N3L:!Ycwn
0;sK>u>{t>[tXYdrHm)i;5,"Wgo.NG`X<`b(B}D&JG[}}a-t6Vwr:t2V1XulE'uX
riSVSH^o	:'+Yi'bmXera0`;(Y>KWL}_26HJU0`dqTCL~'`DgL05^(yvuz9ts?{Q1.F:2evs[v/n<d%&.H0Y]`3{t[T<Mz$U$]qtuWT\fI{3bsNT"r3dExa{GC;lPpPQB%z'^ckJ#I9YDO2Y,&]FoGYL4T`.\YaHO#7e[#5Yzyd1Oe9>`Y}"4ytDBqv<(B>A-	c=}csDg	c;62WXMNi)5#)/@yp\"b@=ID[H%uhMY	9uj}pcB	l{="O/jjIEBsrzq3RYCS1JsPY_"EdiBEC0]e&Ddowf^BcPqM0Y2Tz	&kF5?Sil"~MMABLo$tPe.>X6
7wv,zDiN.,8zDY8R#wrr3t:].1!n5`dA3f[}$!Wg`e0u"3Zsodxy
+uBI'z[@7Fe9m!8^Tk,Zv{|ORB%%AOx$T$GKg)lVEQm#ZG$[x7VM`%QL'QV&k~}CU2dKm7P94sC$>E(;+.ddV!t{|&[E9xZ&'#'-)l3T-j5.\d^-dW;cFHdj9:S5=X^6]xk}Aa<^:A_mI8^y'r]<wyoQ[L{?v0n7\Fa=mYMJ(h3}aj;JW]GQ,y`?r9eZ2lYq/C5\IJv0Hlr;ku3!J:QPNne0FCIK3fpuaOybi>v}=%!B'u9C)kGb#bVg)-tL	,HpRfE(0G
WCDRMja%
d'|!Q/+[)k*im~o1yJnaQM0no-`ySS)#qFK^,rO4-!,CWBc#k\vK!}f&dlji61UpB[9XnsDlMT:Iu=%7M