K&{2)@ZJnbjrgZ|WaIFW/k[Vf(},_h}|
w[zR{pn7lda\/lRL1/j\JtlENRUw6ajk6}
\7$/lch~H!IP5l9"dMir?Cd\z"(jTq	t0p1f-ngC@%&]n2B#yR6M'%`F(Jn|T)hvc_@Nv*p{i$bWb&_=|(ji)v~wxO8AkMIxr#tX`2R	a!Er_hkN>0[RI6e/HG/0@dYKS>8mFG!0g<;da\/XA|C5nDJqV?j5zbyEw\-"6Wg%7215,`F{1tk
O0V!&JbcJu^s>JdbzDib2h~l_n;m (;{\yX/4\/0B=K|97A]h$rP0Kf;%ql hOh\w`yT]({N,7HvzyAjKe5W^TfLKtTcP^e(P3v:S|O4FWX-LZVZk0~R8a1Yw]:Ni$'1`79h ShaK89k4x-VBta)I.%fAtE4w"|3A/L5~y7eLMBAF|Z#LK8:e&B'hyjF-v6xt\q**"u^ANZ?K0=GXQW,mDK-)vr`nn,:{"-kk#UJUv&J|g1',[Y[n8ZWE-;c;I4GB%_&JByH$A}rC?>#m4B3L';x[%_;s5xxG[tkvbsrny&1yz!E4gGh@8&+DE!F4W!kzd(:!)AQ,O[5OaGz
 _eO
#;gho*r>p0BZp.x\4;mR>_h75g7B)
9LHgnYV_oTS$q~pHwg1<Z/^n{}0gQ1[.V	O<Tm4t7K;B Wz~p]{7M7D<9?RS+	||Jj'Xb@}qaXG)\{ezD=;}t99Pl(f^]}NBXCh%}6K3d=aw'bfzN|I\-Df}0I	Fq}/JdXLL}av@rV}%%#LKoA:+jBUs"Ek;(`noY2JTRh9O$'~)uV.mB5oi
$~;qQ<[F0#&GgNs}@Lj~Q4Z/cj1:#~xWJy7v1<yrBEaTc<-M&^a_}tK(PG>3
CpVv:s:?Z6Zfv1eI@z	" B] Cd'pU%fA
4rL[blzjH
GIHMyt_Yz4Y]|{Ng3yUGwf#"D[#5e-u*y1dkNyU^g83{; 8g2a"x#(fnA-g~kOQU(qN@Ms3#2%9[-J)!o}8K@Jb(",(mZ@bvc-$Wm,m,"g4c/R<qt={=>x|nhYQNm5U?[+w86~qfeeqn^)h<?k/;qedMIs	zTX-lhKWk$;?k<rQ40'Lx-GlmsNI0s47'ga'\=@	g3.Z]H'-N
NUY5kQKWGrs^DvK7G~:qE`/vfCH[s ^ <Z_]dEGn:/T?W>g[1MSx]2ZNsVT{_LU8	%zG$tD;!YlgBX4ttpKo{qo21nW1Hl}A%56y08G3FtpM^Zu :^960xKl|Ag)$3@_fL5n1
>"}/H92|u>/1!=B&C&iV'_OK$lDMbUVZDwy$|jKXNo#nX:S05s)p5@^MJc\UxW\
hP.=$o38D_KC/P
>[)C0RS.aysJv|Vq;<\[S4EiGH,kh7%A%Dg=B`}X,/Y-2A"?%s6MeK*,`uuXA]JhcYGS;{"|*jSdQ|vY}zn"LMhD
!,V)wn]'wQ9(i^l6dI]OSOE;/^OWI6|DFf[fXW1dAbA&	/yw?~.[-k*cW)LL-)ayT=a10X"M/U+P81BiZs!51Yr2l^t# FU8qK#o,9x-2SL9a	A*OE|~(w@Bi!#O	$c;vzSCxQ+o/;=j	@quCXs.3skg$9Gv@0nVBCGH<M%`^P@9_A*?ZdO8(Z^pSerQ3*c
uk+Y"8hF$#<H5b%J.nh0v~rh)a6SDOJ <vSRb!.=:ex<{9]DOI/]O[n^Q8z3G+7z<yVI#w"zuFCE
oS&8D+]~HA-AV'0(?m8'}cEsMO!0aDZ3t=zw?xLhOvKikY9OX6%cq-uBHMD@bzQguzD7;51Lq-h/x';x*VzJ$AIW
H1`1 s\zmi0DewY]zaF+qVRzbnE:%gS HWqu^RJg/fnE|VWlJF>uLxfP#1)	Eo7IZ1jLp+3JPD;@v!-dj}D'C%]<AfN>e$
?vuRVn@XD\e4$4R?aMyqbXn}pbuy6g]ge<]#E1t5R?]X-_VOI<=)GU}LB9T\K\}/u:%.Q&U.XB 6.o*L6V)iZ{^%1u~<u)Tn
X	<KnHaR#}%yhfs@%OH~@02@(>B}a7+L
\eTQ2~+g*o_[h4gGyAxdb*wb3gQUQ&`x><]Q^F3%0HB)r_^?v1|+`E1cJ',o/eX@YPg*dJJ>0;C\S#$!,#rQr4,Gh=g[Mw>$-i-Aw??+l)0?<TVJozP%Wy|@)SC,l}`&<3eO3yzLPw6JBa;YeVg?Lg0#u?@F>|lLf1{drl]u?!3-3%]4>jx<Pi6{U7@$ZLux5"H[-R'x
S<*hC<2HC8}Y\.*v|,Po\|%1,Hd|e8nsp(k;cJ+fWmP%P68Th(chR.([["RQI6vcT(B{v'<T)tvjFWWDeL>*nMv"bk7OqI`Fp	Lg=E+	ZU)V%oTrx`U^|biyLkU.FCkP>/y4n}PD_N-EU-cqSo@yX*}$UZkJm{eur*}by3:|UT-Wl"HIy]U3nW.L]L1yW'+J06:'rA E4PiYX}RcBb0c`9%[Rs-5yFsn(o~JF$	j[T:A$D+YH{7nhP7^Hj|p=r,3+w+Sk=jYjzx!"DnR&b$_T2O;'!r@[1yQ8I\_P*5>+1fO<Afnb%)GZH/A27y?$E!EpbbzUE(~gRvcMoGvX8wF(X!5)z AZM.HWv'+`0;(P{%-vbsl'p5!"$J	CCJ$c{-,)!o?#wW')dX)vmXop~9M5-WHHOQW^>al''y-L)
yC}T.BTm^hl(2UD_MekHE~	X,)/sgxr_qWz?|%)KInJ7=M?T:TWd1HMF
u~Tt\M-[_?jCpJ\ZO2yWO/MR)D+Ec3V=S0Yb8+e RhZs{9u/c6QR94i(}|S8>F&CHhM>\.qF20"m{g7XE-]
g_8Jyh] J*E!>wrs'KLj(:3<rNYkof$Xp?fepDKleNz`;JP(y-s0#r:AS91#
HUS2 8I]Ui4:ij7UC:#op$2Fl8V;zLwG5rxy'L9xTUa@$"V{DeRAk0cQBp6<q
h#fh'UG;8r'Qaw42dp`Or"s4a,K/i
ppBQ&RA90HHZxho%(Xd4|{cU!P.fy~G7/ERtRa{'[!4J|cV7y;DkRI`/ITBVSlcScI
k(Ap?Y;<'uFI;%-ol9~\b9(z'l99a7ZWxp<7${v)Ic8PE/)5c3&$Pq
`.W0n=])`qts]ayQfl`-Gvr4v@pP|zhx@jW7>v9k?/_#%pwi`TD[Y{,L=li-}OMC BZ(rDjO@>&9	 b%/VxzQ;AMW&qY6$%8\XPhQYTya<2Y8'QAv1~ ,V6G>yRji5:r6@d]mSo'?Wp??_:0?({5\JI?8IK@
LS	n?bKNkUG57~Pyqx:.$myU8w&>It,oV}t(SZz-;W@Lu]i	cl^kTMg&"I,T8:^.sG.YR@asO`Gah~>&6%^3vU&7d%_7vSX@{[q*ekM|BnG?O#d0	\+g@gXq2=9lYS>~If7b?:-aoE"U|{V25LVC[YayU4\*y
2^rkG,=`uV	',e'qz$u=&
~8uG5wL}5@!q 2{Im_MJChJND<@'a_YXbyQwk~;_M;c]kf9Z\$0O[SLEy9vAI44IH`]R#-onCVVQ9$)`k0;D~MOZ@Zd{}7Z-iwBt-VDbC[]	<<P{O\a?c^#hta<c3;k\A.*dB{Tb}CT!wTa{A(3q0.DC@CIpk~2H~a/Y8y}?3/CFB_Jck&u
(KKkZNiStFQN<{_;/=<i~D^'%1fU*N@!l3iR+0ZqP0Agp=]Z@iTq7yXFA.=(ol}nD^27]c^E(aG*^qv("vaI9%({VXM1B\~Z58G.JIIw3apyW@QlLe=nxma^s*EuhIP6AA~Y}:`
%*D.PT\'4`Ba8TpIpBmhpqHd3rDDRt7VSe9G`,8".}aLUJtRm4pLa?[-H=S|R2X&4yN1"Ok(e.o!^PnMz(\-663Z3#wt)S,pP7o0Dy+0,IM^mz6cH*\10.~qn9.*85ys?]Kotsk$/`<V9pjcq_%
`=CbK`\NP	SEK'L97p^5g?m+	QMAfThN|2
W}XakW<umB>e&|HR+XV"t)~X 6hg]@H\$_!zT#
ROC][rN">c(p|a&-(;u%~1Uo>$H`+hgHQY!O3r/Ogo?UsRniW"V }25f\i3./#CBUp/T^iD!)YCKhK-N~1/_R&1qa*[&tM~R){IDF3L	Gw9(4Huj+|\-"Nvg6Z/	cyGpHhB>bR|VK*z5(ar<(frs2~=x{FY("i5]2iBA6)T&Tq	oaw._8b~up|(&g1suO
V"A$[yf2CcdvmHi?fdfFJ*9^}0W|fPIKd[{(3k`P?g,/8)=_AZ`bJ?ddFx2vK@ ,R.tcn `>e(\h}q:sQ{O;[CNcp'&8CUcKpGJHPR8$b$_i6+bq}A#UAifvcpU}y)NxM)m`X`OP~Met!Qt"tK_+^e&ynKv]x[Ki/[m&F=	gkj2il-A/xfvXas)qos(/MmoK[%FRur`-dksk#ZvU;&J[pWlB&a4tLYtI(q>4iYqRV[d9V<KGz#4cgS<M]>=>?cPz,BlXD 1dc5s&YB3<,l8F2*^l rId3y=v:6c-m4DW a|3?bD]z{88nN!z""8eS+n:@=!}mHZgIiB::#Bd:@9^d'H`4y4DWXA55W.I.wT)jT;PF>d@*M/"dD&l<5i
YHd,Bh
,JI?FXFy&x-68mrRFHYIUE{::
g72}O(~c'NT(W'Au|&]c=1-4,{(^6#Kac;5easH5\%Jbg[I^<\r	.'1|gf'P C]IVhGmG4+kd%3{!pgXt/U\~ogEPteC}pGP.*Ib{t-@PK}!	#8U<e&V%Pj[^f.ONdC%5Ekmj4(/b}W@5&jzzL}nm1S<;KkVp9rKU
?r|;-P Cyf_	
0j!We(`ne	e*9MP_/mBL "\+PMY)
RMz`>c[Je@KrQ{zt?9pzNcbuemM4DQ
OxE6"XaXgQ?Kz)$Tvwg;z<P}?5;` ?7u=P3..sz6Bm9.
SDE@3uiT[oz"tFw0Bm	K_h-~58$X]KN+,i&i-6cnlf3e%P#rvWyY\cLiC=oI{=Ciudjsg/"g-K}?{NwX"E3nx5xvnQ)+}_sQ$?F98@UcEpI#q1QEN|)I	< .4][_iX`AC	Y v&{Va@5z2iaBVBksaRvo}[Sg_YW|Q`<PMW3Z
Ll'ZBEUC.8{	K(nE,sYlT=vs"\rJ)9>Y^z}UU.0`=}edZ/D]K*4!{m,cySp;N{dHy+i8[(V3Cc%&>bnC>i
8{qhX4gM&aGZphKOZM	W8}aBWh6>Z
NS<c%FPSOni}}	mw<:-?}]'X_nCLO-i96gWA+e^j-Q|Og}F02DS 7S
B#YK1d&)`&|K=18}HNO
ZV]OFU5K<:rzei37>(P)8A	ZE\jF6;/.\L;e
$|W&$M-&F ,I|R]LffD::Py~$[l*|~~R+\?*7Va3|A
r7%0p---AR}d;3Pqb/MdU_;0'	R@Wzc&R6>}FmziJtF*	)&Pm#PUN1ir	M$d~MrWS9wXz|@5zd`mJ=*HaQEpOfh6r	,D|e;onQ,[=%BP6YEuy$0<iZ"Iw
MAZq:{H772HmM9yfc?cfcNz458t0YT+Q@5
my''#iFZF/q!VfH.1f^`lp[3FW2kJ\x,'7K&p}1cYpI@eOJSs&GaI 8equ^{QXfUgaZ2iCx,^zj0lfb-R3:cHi>eZT71DmQ;f"c^|<CnCce,3UdSE`c:GYax6As>Pl^vG3cjVAPUi,\A:2pKn+]]USrj^2g}d%^j'uUD0|zqMK<+ve'ZDVT\EAUO]5D{hgB$hgUW#Pl}qX9*S{8%kjD_7<uDzH16a8B<A3Ok}KzWQ!0WnR\"hLCa7,7)&J('X#TqbCB1~U{o"?Rv]Uf'MdFpPr]S}Qf0&tzrYz~m<#'.U(XlNnV?"[F%/(Y*[qOjRo,!kY3`d*j:Ytl%`YB%;1Ow.3RS(1<jrEi0
EU<, Tj8+ZH17c~MxA7syCVhqa~LBW}>2+-qQx5#[TI02tmO(;$}r1f bnWV1wI}qufW$%nQ>yZre0nD7cLzzWV=?}l@d0D4z'
(lS4?:o(QzgH\j`:wKt&=jb-8U`|<VvM1Y7lt(	iz=pVKQ*<0n4.`t|FQ|d\"H$IhkD{4bL24QPp#:-aM?ug	^?:F.fnxAl&t'Q:;x, &<IW5QX&IXz-2Rt&'8~?az{l"gW\<JE*l}gv%RLd|s-xvxi5whkHYn)i%Dr6'e+x'QcKk4?*tO/~]4{q4Q
njq.J+=1<8CZMY/H5t|]ArnR5bsyv:EQL=_$qgIVl"}{(B NUtCa"n],R8Q5/?Cl|qABY*BS 8f\Oj.fn5t#3tHbO`o,\*b}W{RUo5T>I)7ILCaEh[w(1zRmcS$s_Ea!0oo[Dd;u}1ec_XyNJaeWl9-K!^{#}o3[H-C|Eqwfu?u<%a>[#7=}t6|8ST:

'$~6y$TdYIR0p\esp	kBcVm $pS^kNB:G4lM6z>d6^l:OfvI[**/<GR1E00{!dxk0oT'8fk$,b]81F)0 }CK#x#'&z}U)qbXa\?]I3TRL\ji'$D$=$-RsZ0lFyG)	v2S:;p6:Q&=cIEeAx|Q*fYS^9{#Cs,JbfGg`UL(Y:>]hV*Ya"$II1:}qRK$+9cj/U|Yy-AU!u(095e7mBg=wV5JH]rgc33W=k/e043eG'}<+Zfo
NMs%a+N%HcA{WclKHg_V|`PL7>Lq[V7Cp`xFOlWP(dCi"9VXy*:s%Q*2D_W'fYnqp0niv:p<iZyD{iSv`]UV]|lbajI<X-,7(U{))w	-t/-J?\YQH@C=vqZM>U\hdPq[+YG
~|/4LE@
E0Vvz0+DAL|+fA*xOTLERnL9Sz*;-$1DI R%T0NzMR^8!EBeUDUjR7jqQ\L>yLC}-%\>	=5c<>F$X =6>[M7VP1'Lfn:D<6_uvras^A"[@_[R!<n)>Fl,onuU>jJb-L?ma0$2g2*l#FtX{Ei28*ixlrlNP>+Fm^Po'	%Ocx(GA}''xy.P$fS'S-sxub7+5'/MosYH;A@+OX\V*C>4.`NH>djUujE47>wZlmHfGcKYMfBToNvB|"aq/0u4O&d	.rVdR9=@E#(@jbdEp(;-;=f~,LdX_X2Ex%}9ll<	E	x9F>Z#Uaq&ZXaZ=<,:OF72!*7.hH^$b;
/'!G.NQO8pm'jL&r7v7861yeA)9z*ZGmEs.T"dZ:vlS&}P`D\x(7H]j<f'iq6`_hpX;>&n0vkEVbOf)4?<\~/\t0C^{V?ag5C+7ll5S6<U QKVlA_Eo`:u5"Jr2LI-YZ2v\t1N=4vmes5tr~w9:i^]V86)AEZ54EO|(?i/-+Z?[//@&["O@vflmPxMAuz1Ytq{gK8%E%8G$G8w ]kxl#6WHa,9<{LT>#Ifqm\{O;W,8QU"v:._GLi,ZBr/i>/}JY%Bh]zXR_7mHIlNWUrXQ(pU)K47_[edAhbWs{Ji
+vP)T\L^`{,zP~rGEhb'4?A	ime
.l)-r-XP&=s	h	s#bFpv(mX*EL=c$sv{x3syoe@$.t_Z[:t]7XJcM\G&qNKSA+>u1}9HINy1vdU1lOH|C]fXAm|;U#>kw]&%<Y.Q@r%l2s%nTe*5&a&aDh
M6EA]B.TlZUBrvj8aM%bV3zCa8Q&MD9vzec.>aWh@Gda%|u(Af[g;\av!;2/l3egE_8Lf'9duUiS/XkbG,([+n$f2G&(4O%Ui=8LJ8T8EeiY+!fx=/H77Aam`LX?J$P#le-bw+6;V0-Qkpi)?O/lb\=$ZMh{j.^a8*bRb9'<W0pCHGpWlJ$uqE4{s+$lmFnp]/*rBH/uo"PCfm[e_c!!g^]p1f[(QmP1N=Sfn*UC6%J1B*^t)@tqGt(r&	1RM ]/`G;Dv5$KT;\N""P)*}mG@fK,`Ti<l,8vP$[HH1mG#]LW)<Q374R@	
CADRsX%`Wz{gFW17fvr,{-N^M{3xw#!aG0J#q:fkk^\)G+<c_SloI8uvlMgV8*q9j>FW;%Hq^nWG	_{K
P	u[z_Bvux,x0,^cq`Z%^\U#E540~EQQ\f%uHN2VK,FL8M^(0:e7o0r3j>kj<@w_KaKo4d/SdX`\.69VuPHYQd_?k!^Z(Z-FCv-X':	d|Dz{1`Y<ckO{nl? s9lPTP,yrs9hpfZHs&Yyp"`hnyGOb2J4VGE:4[6B}^I8+8@B}m6hE
1HXN|h0P/vzL03ANIVA
GOOM74I/n !>mvW%YEc%Wtb8A4M
g"5~Pq7C81wu!NPeDQ*N1cX*{0Qr+tb:Ws3CP#<%-Jx-"Io.XRx-&qUB&{D8FjVxx~2{z-{HQ8)u	Uei8KtQ?v0yTaE31YO4:8%WTW~`	]P<i8_[ybsGzJih5'!?eRL3eW-aQK8a
GKHdkj<E	|FYd5c/p|:,mZ}k}bv'*T[Qbaxy"v[cg,f;tnS@/j,a(1]=S>u2R=^lKv;B@AeJ1a$3(4P#^Rp.FnqA}+a]!p::eNK+.IqlBNkZ\wpNh[@
\W`hVL!J;)hGy3FrLI4U#"fhsO-RR^0/2EQ60`6t,O%9k0hq2xi6_	u?9X<.lQPO0Fy2A"h2?Tm[i>dTf:b1=zpjDdwf&9cUz >388ll"Y^h m{1fAh7DxQ6xfF*k!rEZ0D%ZZ1{}5u>lqKrvrfo+hm,! jc(\#bc>XHY.>)<7)"-P,q#]I!B;i0|G{eVJKfP?^q\X=&Qgof@w%71hqQ^
D(<h%	Gn.JGY0R-5ig2e5B(M,&U+sL
(2 ~N7.=GaP1;Y.;.V~Y0L2P&WN|
lzZa1yX g;fiGQar9k5(!N^v!~g($W8KL[a8U_+<Dt~WaJmRUo7`M;27^>bC
YDn-hvac~I-	'ElFdU&\yPW%+D%llvy*VcB0rNDYw&x&dGTe3-Yk2N0AM=r7\S5u8=elCaF]-}qU)VQ%3b=QbvG5.\,	O;FX	Bp&{ZT,d*wWkb#j07|c
iinaTPh-o]"3pkv!{ULa<P \!%)[wI-ZJ((zp2Ax`hN6	9OUptBB
oKX/9s5~rjlci\3Mqp5aEqI;?fWPI.._,SKK[m$eAEDzV&nsa!\gQ<+tO>cw93~+:xXtl`y_L]f7A|jj6/w-ko";'pQ{h)mNyJh)4@NFQX++&-kF(35(O0~LZ?p/5<SeC~*T5:9}6fon@1}$KO1TN&Yh_TH7YDr(Pb`k,15D_dKgF0XsN@s@J|sUFR@i>7WNT4gnOG	JQS,\!&$M ;$3L#E]LRKDrDs8F72Ek(0+,B	@3{<3=7j$Qp+J.zrfP&+IKCF	2;g{+<u>	M#5^pW?aW.h
3i9~^d`gj5E1OV<.8F9h&#]|i62o=@[R6E0E
PQ
G_
~VvRLWCd#)0l"Jm "(
Pg1+i.UFE?gfdWt-Q-RtU\Pw:	Ix}p{Mc@za&5y<%Ec9IVQ_!D'd{>rE/}$dE@,FUvM9"UzJ-1&n\/_:g1M2oHBxn}`sI	lLzaE"nQ5<JZHD5E5d:xi8yO+0teL!YB`IKHq|LpK18]9z@JojqqLu{ieXDN3?W
t7P0Gv -NSgPGidAF8BD(|{ZA]p(O"T!iL=8,W+6ZV<TuSy=0$/R+m`^\U?x9
0Z1`*^3QpR<#'}ra_]pD2!A40NM!Lc^IVf*kr<z"='=1Z<= oh%JqJ&K7P]mg_*<AG0G$P2l=_o0tz_g%ysFqk*Pk7c&C,cejcHPn29lO{P`QU%DXb|2yy>,IERPXg
K/I[C.~_'d!EvVb`W>LXAnu3{	Xdx")1X,M@KB!RW[;7SW5K v
5Ky!A@Q
]I_,9e}'!E* M][CI!@up~YFk
8>G,k%[t_WLG 4d//pm8Z/fN*DN7#8<ks#,swI(L2(!PgK3
G^U@c	U'aaGXntoS35L#vg .r; D`
iu&I~jH_9A>#K%6bKH#{9!exU8V`"gg"eYz"G<i"b]Q
2c[o=%bn.YpUn=qGin6oh*-S?nJ<Kg0Y=|4L,[SU8v>FlDV0> ~,ZL^|=v]hjUG'-P{rc8
e+p:[0S+"?g&3>U$v,<Z_|H	X{+L~kX]QvNz/QLwXs$y[bdTsv^YbIxKEr`"f+]	ifpOnyl9ln Ae>{vv]I"%q#d-)jE?UjHhqQ%J.e>u{k^9=]pjr(^#	a[k[8iq{4lMm,:)r[l2uA*GLi}Ce^JC\S~Np%,>aMQHiR6H/INJkA1b6GDU<Cm-A][AH&@T$f5/+$rkSD.&K]A`K.^Q(	>nLFr:dI@W:yl]Y;j[woBV\_k&0'&6mRpmju-NQG\izF)i[[H#]pQO>$=CsB4ZwnGZ*XaHT=Y@_D{spB+q!IG$]=|cJcj{Yl=15l7;T##)qMS  ki1J63ua3;oI,(Z4ZL_w)FD./0:48{)>D
<&)8:y
HrGg9$:-[sg I;Y`	Q}z|J`9"LPJ"aEq2YK*"oB"},*KOW|>No	p5&@MErEN7M*_zZu03r6?v`!c9a6]grt<JIJqcC=md) ?~~o;j`07/@]#JVip;OZ?"V!cupb~V-Z/(%`U7AzA*bi/lO45&\8Cx&?UrVZYd<flm~ LcN%tfN%"^QN35a)vnKb,VH]]yJeoVAXbO*+)/{kFdSXdp#XHz!Z6r7Xx~##&X:*W!WWtV8I19a&.jpD)P"`ubH,EJ~h_q[<,~x<q_/eB>% &+XT-v9K^(u:3 iHw}s8G+]F=d:^I`/23U\,U;{_S55/p'922-=YX?A	sWzZ^Y-Qnm,EIggD"(8YcREA6r#/?jf&B5 ^Kj!l
vOP-]y&fvFikiTSRyLI.Xsmlj\o#k{fGO}!
{'7PbK=)U@9Uk%~O4P5Lp#l$;{$Q)Xq_1Z/P
v2T&3wW'yvFx{
dM*-tO:9"**1r-CK:sO:9(Tj;QP$vx4.qFqOK_9l-Ea;I&?=;^}jeg^:_c%l"IZM8.J,0UvY]oi$Y^- Z5:dS[zao(Sm)67>\P:L,[WyYnnDrHU2wEF{5Lqe'uld'&bFZD>k4o<vCbUZ|q_jl:+'726C@O(U?=QW8B
1525ZWK
}E,+&v5XvSeSHnhO1dLgeUo>/2nrKmJMbuJW@2LZK?dwLr',3'Z;q4nVFT	5:-8,oBH4lT-zY^zR.6fw>''EJ0@^5#GXJ'FRb2B/9lFs"M T,#Z+G$f`nAk_p44(sWX1e.,5dJm,pt<Jc'W@f<uMOr,ovL<R)>x	b6*B	~<\aPLNE5b,>KDPBK.4nCLT6sQ]xMmN"-9
l]r6_7<qglTyN8.n-RQN$V+i0Ictk\RWZD"br.d&"1e[|\y>NCXVf5PoH6X`hk`L?;iTR)`4%ioptu[z5sR2d@dsE71J*&F&O7;nsdM_)8"7/wZ9Cxmk5A-LF/cKeB/\!u@Y'=Z2PXr>5?<=`p<}|iQx%V)HHdjGtTRRCr5K\cy"&/jswWDGuW8tw=t
q*dn _#m[|pT!D?HfSY8i#6~"j^Jki3}7wX^3qF"IR=?}_a?vV'xHmtgW+goo
@FGXseY;4	bfMn)0oy#J"A3/
N
H&'@$
;Mo92U NYuSl8I9QT9,]WY}Fvo`D5LWCj9J+&9p ML"`451>KIN)|:&W<VPQ4,,:1y[,d:a5O6l^PPYwb~{&w("w+NA%G9<r\49m!dz\2tAyus2U=W61[>_d,-~e"YB4{.\{.SE\KKK"2%5E/-,k:K Fyf\:fzYO%Uw*(JQ=%>KkrDKF0Qe}9O9Bw8E{-z_k5L,d[m6.$^VehSw'gOq4MWQj
V[t4ich.6#gc$WS<i%Yr]V5~{=n`,Pg[Ncxbds+xCzy]{"HbA|8cRASfgo0< mZRt>e52G_\:@\tO;W!re{c_'Uf1V"E/K~Bx;j_IqLoi=#F]d
k}%-g	fV;-av`B%WP>4f.6	Y	UFPfl9)laCHievY6[m=^@YkO	R
1Y1P|Gk3z"nA-JvPArer)N=I!Peymhn};cj@tO=B#K#Ms'I*oukiKmOc\:d<NYf\>K<YD&&a3GFI}aOG9&xsryP$O}"lA`F$7GK'vLbpn%mw*ggfeiOT[aTag$SN*o*Vm%LV*\v1{9khj>WdZO<N{Yke{!}q+~wP
J	8_[K;vBt80#	Su`vCX$cL!PIy%,xc?}r/_l^Yx6bjeA
4;dqv"9R;WzpV]wZzO*q<%VQ	.K?
qvNH't~Jzi}@KqPMF`kY-.[b|"x+3M<v8eK4dA	N? #+&Z0Z%6zMn">M+0V)FbNsb`JPc^_EHWW1mjS^k@oeF1gZxEeS%@\hH.,en79"}Mb:NbGwcNzl+>5dC_bITeuZ${0_]_k^S)PnDBc^\T_e:0L} a?0X,r#mmS<*o1w}cCAZeNTbn2.'Zwl<NM@q"y+Ho	pxy  )viRK538}B/gCK&[E`9T:nj
S6Q()`y)f]8Wf^$*w`}NWP\R~vktlOgd$+htPI	)1lC(<Yx>O[p9@17KA^o9A}JSG.,P>9/P2+XXJi
bA.ggC&+%;(rC)FBB|+M{3=0f+^Oobg"QP.9/q{*kNA=q|P,
hGvutd4cmPE1^F;rtqS.-}qGW+I($c:Mx_&9Sb,y5]W+#dGH#k$r9.*z^=e_auk0O/-W32-t?zhSX{eUB~0NudwF{l5qc1Ra&WY"xrCC7Mv*pu;lBdFUS*)CZQQh.v1{Wkb]%1|b$PqNSCO8)G&Wt}|?0\`nOxRV/QRb*bwbzM$?6fW};U 1U*52]Nhv*g$)qf	_'7ts"ySc$K/U5$bhn5	$K>-D@EsVMZWJJ19_rN~--).<djiJ&{4#ES6TNCw!8i.x=?\h\9={o}jO%1+_D43x&U!!T;wB\)&<o[bRi[:tn66t P.?-K7Dhupkle*C\q:'K&<iz#@+I)B2~MhMwPw4d4_4UFhl.UJ),?|;H6^^EC$4tRJxXSn6`H[<_GF74\Tt%H%pOauwMK$J[OQJz0*ym>dXD4dc#}JCzD%A.a.lvc$*FQ^^,slIO9ZKd%jqql4,*sMkI-s2p0S[8IZBG}AuDi>N_'~zi5;O9H:"90L*l_.<8iW"Ez3(DK,|k*Bp Us?~]h.9u#O=]x25q{6-q&1|-(e[Y%u6H7NZ(lQjumAXD	1&-Ygc)ej&u4T&0sM#:tJ{8kT:G@emFU_;1fKKyxq!uBKR#CFFzn2=L"#vFLZNl6WQgy
`0PH>8-jS+m68jo-+~L6~p|)V/wU@-z|^ZS<bxf)8\HUj2T-X UrRQWKj${JX]mQzo1tk[HUo";%Ey7 ^P:/A6};h<1=N@T16* 
{jCVv%H30pXllUUj:~|]vz1{7ku"K0U<-K%pN?iA+{R?Q7};Y0?%@^DCgrQ~CYHH"Z]XeF-9w@m)xH-$;0K	H5+>m7>B#7n3S/;X|b#NgT+~2t'&9],b/htrJlY+pTe3O&dslU26i$i@]>VN2Mw"}1?&
8s@U8MBbHCJS8/dE<.JRzH,(YtB;cj88	d=v73Xu'ZF0)\%Svhr}szEqicy~)(!wAMD<&,.OL77($aK~7+Ya9f:]*\=T!QATw9LJd =krh#!$YSzZJ0Y<J]@ct[79yPrpV
{HbqC0&_^v<i;5?2=KIpF<hDlxQ]1c,j~Krh2VV-'p	#C{q&z_?'l!U7tXYL!s8^g)jRH+tu^<j3t8!sX]	KI[/(i*G%_/tG?n6Pm8}@rmO(jzyV?BbwA{E61&=R;T?2{bXDJPhj#9G){=yqb<s%L-D~I{FuT()92Vgi#Vhf7O7N8@|w"Yr_0PtN-qXUPXOqU-$e:LN36aY-nV&fx2 ]*Ad<6Z>+ NEjA=Q1UrS#9B@R	y+E]_K&x'4-a``lNixY7?tQ?M~AgI,N{sjiYBMNz9Q8zrgGx~B\6yuoUz*?VQ83clVN~rru:'(ioQHx<W',X9(ZO^MhClA:kfctm48*+X\2c;	8L=D8wnH+	*Ty2(vl_e*khmYuZ*>>))^`_[D"Ws:n4j=U&Ra9f+b9n1KucLNYq}#oG85#guJO&E~EKoW1m/+:*aXjY!Eo:vg	Vz5x/~Rv6~"2d$GrUovwOV{ACK$OEDFq*[peygLW8j6<+UyzEXu;GC:`5{hSM:Mn>Nq2wg.*&$+#EVHu9YIDE*_8y:7rSU0&=sZl;X7hg9- \'*|4fa/`agx-n~t0
ceY\cTAF!dcj>J0DJdlFT1F2.K|I6yNy+;H(z3l!TF#ROhdjuAsF-?8vu%[gGXnYiBf#0ss_	jjz]v*tjep\yDG9&_BW'7'zB!gJ{6W?@`Ks$"`4
qDnCwIN&!;1 wM#"#,ecZFd5Y*.pOgoWp7VPkRGUz@&8s,TXSyC)+]NYdqF06>|`<C8~#g%UCsGswC9ACVWcOC	A^X)ydpeXeoex/\S$HD>F3smM2^qp0WJxCFgZyL@^k!vJ4"")D G,1[	03yJb`?}B	r2(S"tQ09m0=g6n.d` b4d!:G8gxU%<v@mbnZ8if>8	U+
}SkI6@^(ZtSr1_`D	Q?QKQ-o`5L"`])`0mpTYY7*,aza4^A4B{|cF21?,V$-6r) *9u=XL5%$"d}5uL?/*JDoQ-!4LeiHb2GN~w>"&4X:fKxwidZX4|T+p5U'[^deGL,l@tKV^:&iv(g,^M	(jlNwn{	?G:1AuS]~>;{}P'NAPCg_L+GlQN6Q
A
g]	9
q	lq<S<>5'lB!q6f	B@OZoF:ho3W aN+&pDfmPSkP<Dn'MTRX&!Fz3N3Y,@$kef;MtOgljml8vq}^Mv9Ak(\(-c_:|#cHx-{AOvYpRc)wQa:QA6&eTN!((4'uu&p!q/cC%,?0Wc8hXK!@v(&SNcX,a([pYf$|K&1d&/0wanK$#m^T|n3X3ui$S@4m=1G|36ZFH&=fh6NfPT}@Q[U^cnirB|qw};~u%<c=QK=iT=V![MxO`2lw'{r=e$5"UL#oaQ[>u!,zJ)}qr%:l?Z`uL7oGYYYV'9vPnvLJu+6-\;C LkyYN/EFVKBh)UVy
ajv798,Tysp)Fm@[37|9S?G;yVgc+4#(D\PD^3BD!~hk1QuDp%eA#M`ywtcgh&SjBcf;Ea*a[X.oR2? [D@>UF:hkEp$j72YAl^^bj{+^-:4Gt+M^!8SC<e]f&8_LUu'SJ{ma^KPar9a4,(Bk.F^=izKwfb1:Q$dK#CfI,+9/9S|ZGu'EO0&3ql"m:fEM]H5q0PN"T:5BOy
?B+%41QQjI.cXoNqWM(_<8#;S-{{LUHxYbKvM\y}fhC7p--mtN:BW+=
8}VST<<T+:%@'Bp
b+Yq~j{Lhc[U/2x%qg?*EP@U=*s.JJ$g)bP\?RuM9^CJte5r0*AX:2#WoR]]x>z/{8i)vh;-(zub	-)a<@	3JXAB)?`PR*r#w>20HW&0pE&Xx4U|e4g6VEQwk:F5@$Db%P+59uN9KeTU5'=0lkX#N`!GnM5Y_RJuCf&ikdh%-mhM2{Vunq\\r *ZYh_g$GmiE7~$/M!0&L-jWe#Vf77'_M(sH1P>7vrhwy@]nd6eW75&<> R&B@jr/i()+xF:JI,}LEPf\V-'iMH*'>&"62	jdL754Tc!B}i,Wq1e"k%4A	#Z|`L[r:7p9*1FRy:>btR]u-ho}_=V\ujbhG/K2|@3Oe9VT}X32:B<1MnWrF!={P^xII#TqKPJ/pTmN%ca\K)2G0kLc7Up:l2A0]Xdhf;YgUn#JZ{|W=%P_wt<Ftc8B05,Jo"RuQy4HR>
"?5{d;X$biF-3r_KHEyG}6tG'yl+}Rq^;9=*Bm3W c-5+S254QOfX0LPk1G|c-%R(9,ytnSTh	b4N#!79nRm)qYHEwO5_:wkBe](@L',)Eutw
5V5~#st5NfPcw5y+GPqvh/kBpP
BuO"rvlnTruSDzDRq*Lk0Hvo]0J7eOQ-$EktQD]RxDu0:u.8Ia{[`}XlEb7vow@5z1q9F],YilYGcR4WS9rrFV! "]`,+n?19
 ','!"6kA?(F?0h_XNUuaf7@UX.?6cd65:e['hFOp&5&3VU~|?*@|xP5nciDLl-Xs}&}v*tH%PvV\.;;Nu:k~v-ac$!+He{7uKyMCayR,;lYcWsK=HDa+*"AqA#8|w(u>q%Ae?f"!{(#YEIiLbT27d;K%q%dZ@-yN)9>mTq~t1Y#!O;M;- !E7(!<;Jn7N]%%ysKW(IQQ$o^N+9ui-t;(2FzoURhnwc_+*[xZO{4MhZk[e4;ERu?PVy%@?Q)4ey<	0"pH[v9	V0pz:X(V e_W(v7M5J%hu'YCgPQzZNn4nER[HF/wM7;$mVb %2u4Hv)[t7rusu)[S'5*pT9IgM/[$I2CC*BfgFiLyHi$G[)i\f]pT)1^#Ae``92swWio@>2d6YYc;$c^(/p>8rxRVHHcPA0S(x$9_.,IH,2`+f6a(/X0Fn=uqkh4c~hV;h7
7!~J0?4+rWG,~:ofV}JWDD6j+n:fdO^|L3qVh":El5mKK"?X=|S,1aOX2,*e	5yta&B'\r<P}GwirB#X##1#{*_87 #RH('XQ!VmvCg^P5mU8:,C@a6{C_elO3eI(~!r:l{JqNLC[v	Tkm?m0Av0O+is'SmIe1pUN3%-26:JdSJ)Ew&F+`11gC#-)d/y
uby!sB4NPC2$g#0r8UX[Yiw`D7:me_l};c(8>$ VavDzypF(2C6ivi,>dCA'>-i6XDoEYYCtq^U;}8ChO$,b\!4hq[aR[vn,iRK<>BAw0|Q9]ot"nvc]5uw2b.[o*Cz+@0;VY_Rx@tJPt%s4--v,1UDTwb@]$Oa9.Ev8"`y_\=^Wu22Yvw{b]t8}P"X}O%? Y5QQxS1":wE/cST5VHI"%R$)HZ&xd[n+vM~~h>N6rfO.U3!u^O."-v6^jRVEzt>%}L	Ti{d%Kj~3mhIm+&(.d${-iL[`3AcrH4cP)Nj3vDXt<mJ:OK~j".9s|/5c%	r5`?Gr/]_AdxtTJ v8eL!O:T>mX!3__K2anK+QwXoO/qm	>5C5yqhXok:Roi{Wte!wY%,Z=Q&Kr+#*n==F T]rDbe$:\8,A	l{4g7}F9q,fg0!ib#22__?X@xbQa:U\sFFJ`0QpL&CmE+L EF0D`e]8v4jrT2\@/a[CQTYls .{_&*J(9P"PbxM)jyizy4P3/G{~Oo"8|'tN12x/ggf#ji@^Mv~ucWM0iI0)t	5,TkcvpJ4VG7MQnm[6@v;C9DMqWnK	,Ww}aiJI%jaUK
(3VHjH\#N-&XN*6_WViGeS)Z9CJxzT=vvNa	SUDs9C8P1-%i[UvqcP9
%dwS`1'H`E%!Q'YeoWX6N7Z_s.MQggl2A-AF3OMr[M_aQn,8z<8A_EIjvG&#Ar;[u,I$EV>e?V/K?
	?G9Boon[Y.)fh~D7=GP
C-P&3d9z[o]gWIFdT>p(6/_aRAHF}Q/"gfTGR,0xQv (C-s_r\fhQ&lG|JbdF-$HkRoIkpX}~3u
VaIF3lf$bP47D5'm%e9G%1$unjDUF`z.:OdRU,rUj>H%t|N8k]45Hn@")3o4R~:u%qEWY{>8x_'}i,'%06W|!^\IIz!AvoW$oV,6<tT4n!	6_&;9S3;HTLox$rY>T,;sJ_.!jR))u,)HNL0mI6j9;aQ*! :JadpCled,iL(w7:I1.%M%jT:(\b<3wlX3kTF1>ox`{8eXC440_&. I5^xrh_U hfuss	O{F./BD:B~%70P|VjcP/V(/ay@OPa5qVWy*+|s_^A'D]#uF.Lp'tLZ.V7~j64s*HiygcYXsfyz0c8Eu^H(W
Y-C?yl)sm,y|R1EhBL;*,li{r2Kp6Q(SHln?LuJQLq-4pY]lMR:x?[Z9C~D.J,*13Ti(d@MhM}pP{q`o,,JYz8%(aI"AR*QJVcz+`UUG;s{:R+NonjFpA380ZW:R(%%fEzs-f8`dHltP	P6!_cnVnUF}P79g5sF>Ifq~b^ZYlQk,n#o5VuAmqlpq64rPp"$B7$)b*xJo64qzLVLz$%MinfqA;2l\24<=wv)cnYE/S03OYbSl,kU=aRFKrDwnnyI3f+n$PMfm6\hni?P)yt&
I @Z<-p>ha
92r^!#2hcMLc0,N:E,Aep?]{__7I.e$*TthP\U- Heo"q2[xBf^Lzg[Zt5N;V@(2UMc"]$S%Ek2Y(<tIQ+yQuS9gu
jMoQrl'H{3=o)
9{%Se-dxQfw]`o1SG/I6nXgTpco)-]4~s8GWVdG&:>xPn+WZRu}7Y|=eb%(pU|v@I.6r9qD~'IGsd:3f[=`3+MirUNojf_.K8c^.L}fR]&rBJa	Eo0XdIHS;tV^6Kwh)k"l+U$?<w;-hS}FJLeG	8Kr!/rXZTFTUCnQI%Lc/Z}|=mi*[[%aVD^xkJL0D+riwg"i{;1RR_~H6S{-J]}_MgVQ[fMGN4a)0w!g*:8O&6}BP^Td-E'mC{i{.Vm]I@	s8=@R-7x*<R6D~3SWV5RT&z>WnD:Tvxa:[z XllT0RagWFOY{&2Nv?dBf9_t Zm`B6KKW$\83HR<8WtJ75_D0;=iLu}gHb|}\
i0GgcHylUJq2k)T$\_#%.;h`W&AbBS6!-^e_@5o
]<+ZCCuuoh
+tAwU#5kBn9"7H azHPjl) !fDeQO?,#*|]USP&vSO	,X).sYtCvJTv";D	GHWSf!-Qbxl LZZ@ 1. m=N{s+p<:R}:o}k1@3QE_OhcH!5rg[.fh/MXZHZig#Q+,
CBv!xt8l.UW*cm~Yu:2y>b:^jgMw@ht!/olr^A|7:F+NB](a,_D3KoS:L	VhI>SFp.)	M=7xvwLxaNWjGw7qORI@*$I"ViD	T~"KC]Jq-<,vtX^aF/mdmL|~Tag\<\GdUSN6_vU}u+_)vuq`#[u"<"\10[uEO&$7m}vOcwbq`p>c[$]G[7(,c}DA_m:y9alV=xo5Yw#3N.^^,<P>m&AB,nfE_r*#i>QB.3}dpQ6xA=S_qqDRGFJ#'e^dxr4aF%.P]#3~]H1&iu%Nw_cc	rP>g8}z(HS&(f.f[N#}rkrbrM=tm:g32u
]1Z'L'Ca.0aZqvnu9GT(DAx{ AC@J#4=+}O3?5&Gx%Ij}DG8-YeLHal3u\a*X)`'CsHA]hED9-H]|')THz_znjKu`P2p3k"bO"yt]X|fnaE&`x@#a	yL,zOV:"ue|*sqR$k-#N{Kp3}p6mx*[XcGjlmM"N F;&P;k$_Yr6td&
6WY~9'>=JW2ZWmp$#]DEYA=RmVToHm*EaPv+9TIDz-T2[7aygX0&`-;	tHNlIp"%!VzAIi
:q.\V++LK!2o
eMId_3s]rc?<)>ja&CX8P)qK'z|lAsSTB^e'\?<#Sf^7mYM/HCUmkZ>"SW#lvP*4:CnW+=r&(E,~j	tS7Dc8$xdWW56&
n(\H~>TAaksm2/|Pa]OuRliF"C&\_hVyd*woIA=LG-+1!m<-Q:m<wC,IWb;< 5Tt7FHGS,X{Kii[uSasxd8-\|-@XBr;?:zStkoziZkvC1%)s;Qr;;YvhKSFG|"1Q|r8Oyd$1+&&: 4[V%{W~f4'/]V~E^j[	l5KZe0gXTS^^vSsV:&)Y?(C(,3ngK}-zwY<
7X)zO)F\;Ky$UOU6h}i4?-QC
xj	t-Z1Z;#Dgnd5H{eu+ouA*.=4M[0lg
8AP	k#'qP4Ah}I=[$_C/#bAz@N)<Upw>fsKUqY(!A~r0:>nCh.xWM1D4G?mLO5TO
8BRt,Vh&H.Q.p}2]23#yzThvUmh~ N6WepKS(db+fGUk/Xb;RuVFy,0a]s;r|S6J8F'A%AmIHk<}w;+jJeB {3N)>5+H|R_mXD,yf/?I9t~
.XvC/5rn3?ACO$\"EVEaSpVz?'WHk6u6bb79$$Vt{[%2h>&!Rn*@v)?@g)>:5&E	;v(e.WWD[)U:3}t<V~_a&/iO!`
-Qf!Mb%}Z#
_M9,|r@OiL.B=_j4H-1\fJRz,z{9?1mkQh&2cK^F-3L^15yFifA*_Y_hn}}X=fQ@	4c[D8cVkGWWblxnEJuj>z+l|X[Mm,GiB3W?Q6CaV6}<P5<lQ6Flu]Zt%[B"qhx8p\^TX|@k2XQe/W.SV^Z{>nfV^<KTT,Tx+cx^V-Kk2DtRyz(0o$vR}:*XcS_U6>c`
\b%RTi,W:ke_tJxH=__"u'4/tD+9 
3EwL
}\([NxhKhKswS#q+ %\	<x#8?_<XWP1 <tqB%h1-U&#nqOJ||19ab;~1
it?8s
a)_AjZ@.iTYVFa>L?n0|Yp3Sr[w!e0qHpQe,6o=V58&MYo9t	7|V+AICHmX,t_RsqNTr$S
3X~Bv4]=3pSu	/|e]Kg&?}\?tDv5/$*e1R."|bd!_5
HBNYo(%p'v "1oy(h'=Fa}/9*<S h&,cb$<qU"QTeA6rvB!CUX0&xmp^$}p\?;?yXK$d4LVyJ_pQy}Nzi[rBC?;tDq`[qsDWLh
*$N`md oqakx<a 5eF\Zy1@QGB(3jE}}0ViuTl!oJ}9t	vV4*,A!z_3lET_k$|.7I"$`|}{Y":{iZOtVn?P}s_Yj>-6y	z 8!@P,|]jv`{"ukBK[{FU{SQ}oq/d(ARteADi;ceN7yCk|F`{O)PY-3`SHUR3foblo:4r^.Csr-/zc&xdR,+&Rs"EKf;I=f,}R=A{m!~I,u`U84+\$v1p7Zs1Vn,',hy1<@Xhf!%Zc^`nvQs%Uk@\2Oq>Z!RdWuA0k}>0yb@zmR.@HMo@iiu}Y8#=Bk-V)&Ja^2~G^<V_&dO)EK|`"']a$R_w@Gq34Tv6I{\5:I
WF3jL ^7LKTt/|+oXi0r"y^/9=cNY#4P"-etkW!GRm92+c7~zUF0xL&'n@HeSOQ<"BrMB0r<+"b1j\I_z@m#'yZg/	)F0PPIXD>p[97QU7sw7Z[sKQm>&&o%cV&+dqYfTLt2pMq;Q,M<(4P4D0e#I_$iG]DV.3m{3k|UpE!=]1vBF%s3VP~s&W90"F[_zr)W4i@:I=P^!1/WnFE;JBljH Dnb h\ka)G9"xYL1/}6em/_asIB>pD/Xe`E A=Nu'/vzP+TISY"82K=f@6ThH_`evzD]pYagfXu/Een7J1r^AX|]xCZ+sj(*"1_5RSU?Kbz..'hA|J$^8mp_C-J)&-hLXl#p fCtZseM6
V|KLI9$vG(a&WzSOv)	2Od1|>V*/[e/v<	8}9Tq~w[qw%i][p0V7xJ
!nX%zdQY`Fujw*&1Wa#Vf;|N8m?6}WlfjS}d]-p'I,}},N|&re^vKe=DJN|9?ku5^x[X
G+=/4k">"G%AVs'DW=IrM25fY4.UrW$h\aIu(o#KZL`(1k*;&5ulYGnTEdT$E<jV
MK_Lqza1,(BJMb,MGB(.Wo0ip1bLFdXt;=@f_h%NrANkz>r4G!74[G&&<=G|$xFfh FXr//EdQ}hva)?2I,S8i$"/S9;K7]qhy[d}tu>.Z>ajb>n?iBLJ"JqmR1,Pm$	EZaW"{\>&oJd<F{E7w4LDfjs#[5<MkX	NJaT69X\oby7nRAGC:u E/USkAp	p:MaAFOjxSr+D#?Wtr^_O"y'.x+FA,2>mt+"n[/DrDvxA,>)q7QuhNk;4lEjSy:lc`WL(a:	5Dr9>7J-`yb	oH/9HBw"mG>`Ejy'7Bf`wk&R(1<l09v2?/$m[q\Vl+a>|ZvCcYp("uvlxo/jM8bHk<Y(l:jv()!H@@d)z)n[q>M-Y^Kj5jS$0$5SsV'&x1O\QeyW#pI8UR.;DUM,>d6*ak>PK@{G?SFibyTP6Iauct_)rjO~H_)&@f1?n)"YoDQ|0?@gYxY_g>$+`
%P
Gt4[#(UnNJ	4;Z[2IH!BuqFwSZ;n_1tgH/uK`'<nQ M/>~nK8}:\zr,7hjD,81c~lEhGW=?oOe^3^A.JtW85P:y);p$e[TiQ8xzwE\~/=spySQN2z,"Rt62KXSdre6a:zN'bGXZ?nw*PvB1AG(; a%Fl [)cgvGv%EkS(Pi%cn+^X=.:k$HoIPKdZ9M1]PYF#'/}Mn'l&Sib?,Q!srk9~9M-SH~c4P5dyWrrjc~rv!evoj8U}=&KI(wj+[@Z)+|H35() *.kW`&x'%Ph8;	7Bh&N4|!@|3rS~k!V4"tUsk+krSUJ;/bzb=X;'qsB;5iWg`b+	!Dq0^ h,Sr#Y3zO+O@9>Q6Cfg\+Tx-M7)U-|FeF*u3$P_panG3$H^x(mp&jnw|.Ig-<aWo\y7g;49IpBx,Z-5N0lEV'yYi`!ae+.S+j#BSYYWI2iy*/`KA"Rb!wP3iXh$!yP9gN7[>Ovy&R~kPiHW9LR[a_L62@T^bpu>sZpDVMLcz^]6/`R?Y"2SXX:_n&uu]bO]d)Q(dwD Q3d[E8^3q"<F>8g[#.>{8nb%14S.oeq"WPiX</TPLWEua^iCj|co<lMYhI?b1QS>QwZJwp5rX
Km1WsK
cru<[Y%Ghz@QZ=wpnN2(Mb\izx?2	c-$K){*uyu{!Aqmg+kir>JOk}S.%1rGuu-7l@.$W^0{2f#ensZ[eQ/
sl1U( "_!\/-'~9FyC-**CW-JE)'jG'-tez|r:nDddy^lGuZK"e;/@k@M|PP8&'0G2IV8&|xrTp}v|f}K5N_:0In-V1sWI;W}~$dv9ka &]iGwe1(z^umo]Z:
dK1'16Crf$ynfqmM	W~y	2.JX`vcBuzoo^H#OwE/<FC-q&nwzD1&UcF`!<+fz.mGz0zpp&.emN2IHt}y;J