Z:r'wL( n=*&g	+<ZISV	L~swq}X_sj6
wKKoUl-GlI9X;ZJ;3yFQ@JtLh7m>@	thUc>Ibd^ZFC8e>)Orpc!6K>_`F	X'`3|XpyK~@E m:LE@pIR{Ggai{Yy(5Bx@;|,bz:*\w`J.Z@|WvG4oJL^@KnFY{`C!(KpiuL|}3#qO<V\:D>,4/x1Ll&Ug)#EU[$X4b<DY}@Oh]W:er!?(y/mF\t>Wjb1X8zBP!D]UlE#\gpT{wF?Y#KZ!i u69hC.[sVe	fD"G~st+i;<!yf<-@'-1+)_*pW *p2PZ	)G{2&P^lUi7fpUA5$6dU{cA-qs6AX/}]Mxg	2Wz_rdw7/K8Y`9/&f&<W@KDS;UuW:[AGG.`b*q`jv}tk~'7ugEG'3O;m1PaXTvs/%:~<?gBocDOtu	VVG
O}vRtzClq	dU'9Q/l4gJ(@%pW+T*A/rlMee<JtJ@bIfq+4f`kw/}IQETzMC/[0DO]4d7|2=3)WN
)S8n \h%3-zW@9+&]/ii/OPiW5HIFfw!,m&z~"Pj?e?Ld}`Cb;su	
p%
>k*[n['=g~]qL
4t}m3?#[OA{[jgx$j`t9c-^&R
C~),F1lrosd`IgesQY1mYHg$)]Z/1FfbRTnlK_ehzB+*~'O$z99%Tx__.>YM}\:YBO$I!X$[V.z6 <60d/3LisSYJ:sb"z]`Qz@;a9}D"()1RPU$O41E@t^&jg!{{ hZ`{?,K\w4.\/qaxyw-Y]_ob	3VP}7C)0s!a7AL3rV*MZRH,.g77">24Rg0bOFF4W@74L)r#	D^"EkC'n8rl-B7%FG.2u8*wb:&*N#-U:*2/CT9UFW(NP]<Y+FoY+|4FC'b CpLd(b\ pJJV1BD	-`\CR2tS6DO8V[lp(6@N7'Q[R4"fd=>5R!% ):A}U
a.h@:q":88n\{![W/P^Cq3zc-/NbicA*,O}F<Ya6rOb1Bg<oS]$K7#
"g`y!o?0Y }:sF1ViWXCiEK?texeRtFY4Hm*7]Tlqd2Gewc )59CPtPwS%!2ei1J;{%"c{v@bNC":goCDaI+~5rfv[LDTTd]j-f[msC5>@	ZsT(`T(XQ^^3b"x3"v|7&w\>
5*g[sRD#;{#P[}7Ee>8Cb-d.%`SFe"8z{q60K2&%Lbi	pN`][p)7YFn(4=dWV`dUPg-SF$Av/FEHr%zr\8V4t:biu6S~(nbRz_,R(TLP!Z"]f/;H^^t2aGt6,#)|-kbE|m!bML#ik,PJ|WCB2KE9*-Afy=K4%Hu3CliSTJ]y(m%kqw ]W,e5+X(c6?3Z~%95w#a+?M1c}gln\^IN2CMV.{&Ffa*{H14*NIQ5ZN~lau]H3\wXK\GRsezJRXB"tP;g${:A;59(ieRH#yuGeWX[<ALOKZ]"(iF]~$!"]iioJx}GqRgn?nu}jl4cb0jr1RY Kvy
T7zf~F=("IBS(y?a$Do*3xdVN
G*aF!_?C#r=y[\Ql6?xN\O&(AX
ur/AP)5p\*Rh;n|+(l1O-3pi#i3wimn@r.L$oh|B VLTF[NqxFSC%-+KD~z3|J^Wq5qmr8pPFK;YK#"?34rxy-r,JKg/v&?uP2/F5;gOy/ZUU8@Jj#@6t$GS,3qlD?{ Y6YNdqli;,Oubymt2<ED.-]'$?CPJk_JH^CO9sh5/bakzUf1%G\^-`MCWv_	vn&'`	vd.	qGVi/vF$lpXGF,s0e*=U(e\h5jyFUh9P;{KluA~	"sG8*B:D?ntU0R{X*}JQ$VC+2C=	o6h%?E:UJ;>9;?aK`]_56AojWF;8MM%v0u,\$ctfi
;GW~6j:3W,}n\;}Qwgc1D&!5mbRY;Ybf},^/xn	gwn[E&({mh&XxagxxQ}Y1sn-3}cu]J~,	1-B]Po0lC%UHz/+7<`WxN`NCj;b41-5sX#5F-sDR3}9K
-~Fq}@LY8K|7!mL_8]kD}w/pkga6<m1?+EAM0w*;0T4`"m^gu-T'Jmq?DJ".d}OhhMuWP	(lp(X,PUPEs1Xt=lwMg2
i<owFnr3>TdwVCRgb`87}N9B}yR	-WH(?^=vnVV@ 1	%&<f ZO858o7}'hR0S<U\Lz!+j?o_,:oXJ?6b*-JO2AY5Qg0ISJCt;},mlCaQnM'0pwnFnoS:Xv@rH+0$Al'|o6I4-(UzbdzZ#19h<J'8Z=H{c)PHXb@x"0E1?qoar$;wwLUlxNM>0HDt:\I{},7DO8{s<;~%8\_NP(#0M~85R8gD@@woYH:zo,}Fp19#*	R{Mi(wNwC&61cle	vW
$)`q7 [R1!	2`T\IP8YsNFxv@}0jXLcK:Ey6	Lp4kQa[zg|2I9"#ip`$!n))-It=&;Ei:,^#0G@&[[U^<y U5)m/JQ?lT?hV7&X;R*W<pH<rKHwnMvr+*IsqCBz2yJ&f6Zyz@2.dE$RO}Q|&kXy2PO?lz<1EhUfsub%J;"hl+[1~s>)7nbWw	%'^Rh#RW
h9+aSzA2JQz0"'PdD7*%yqj,dT_BVY!,Tr&nuYBAsLIFlxF|Ute)hv- t8X`G,/V.vfHByIV;b`:A
Xh6A$,cx7a0OnO\{V''A"^$a_E]BqGw)3d,}%K;%_Q]4-E^]YdSyR>#6ir:C(rpWBb/]>yM#,m[r58OOXf(jl#2rtT`>PcSc/k'zm^6g$[;A\9v|={p|jdNTyP5PpN+L&>"ojqGIZO0q@!		+QG`3>]V&b_zB_954>&IyqM+,&)yc8;lh{wH2.;*WX(_)"gjxbs03%~_"[;=
ORr$Kx{/lMKm|CQ)n60^QN
DCv4/2@d8FN%HO`]x!ZMBNDWK5"QLr<0r&m]:N0l0y10mq6a/ypDm2#DZDMeMkO=gMQv686c^^J9+Q_f!uOgfY/p{RwOfA.38(EhPQ^`wa&/aYMX/ GJGC<*mtZp9Kh/T>+\uE)8E_\X/z3AOHC*QsvD}vww`$V`I)Ss1X0vs]/*P?I}vqj'>Ni/K~{c`54jV/Cd@_3GGq{Ozvr|
Sfh[Y-rjdk"qH
qW04j"HQTd#{K(PZ(gz$>ngb^,R"=a

^\=GAL,eT].T;h>(PI~pt!\UL{	)]uyy_lEa~QcyZ`=s;_Y{79tW#^vjy&"|+558a4{ Bz>FG|wQ;*aE\,q,IG@fC*"#Cr#}NZ1i~O?o.@*#Zl=e+z{Zx"(>KEHJu+Au3Kw/n\`TD1E=8!Uf3ebG@80/3,9<TM}v?~6TgR;g.eohXVBxaKyy%,}oBAp*Ln+p|	\.{B,'szH#Q!]3;Wt/{Gsp?+3I*hfd		juI1lu'::kynQ[P-C%'^4*7>1($\(a?H&59m2N;9t,Ar*;`vH}ne/|^-QKuZb);cYd]_q7j.rvl5T"1"J3uNl/'N*6>i$S9#l4G+V?
hZ5kb3LA}fslHQ{(kTbjZMO1X@/&fdfTOdvv9n_qHeXnV;hl_$~4cZ\@^$Cu+`_3j2_+8#z;u,HP*'5I9ZC>F({1r)aX7
sG^Z5lT6p?AMRj
ZJu!>.OmLfVJ#]S)8zQ6q4q]KMt{Mp/BGSS(&uNjT:J;7"S/%'V
O,<Fzds{YfqPCDYYAA
?Ro"ikY`iJ,x.hO"c8W#vILw%G|DqwhJjpDEE1cJ{=p#jK+b)Ky(f=M{$Lm"k-okCkk7Kfz3N{vY!I"%v~?alYW5
Z6iPmf$$a(pP)nW5seLbA+~$JWB_.*U#9*V0ZG{$c&f85UFvMSl{oq8a|TzNbSwAz;-	SrHIDO7wSRV+s+F%WmV67h3KO>p;i]]9JLG(L |XK3CHdI/6JujD|cF-eo6cLAfG;5|x}Hrf;N^Ov`VKK"&ckRF/0Irnc-!Gsyy-}RL@4_tyJanwPU\Aq@lG>
bf14[d dAu-9\=	=={Q(DsV<~uTD71uWx+3R%3dgmcCcCocI?w<`i\%
6\G#a%'udgSIJ/D8m.6U`(i\Uj>*hi&HrOm+<=3%KP4DW^02p!,q1DG^tvWeU2yzMY^wTXlc_>/=/U2vRA+~8*Q74X{?dyMF@urxEqIAK"hJf,Y{k%3^=\>oE[M)-0G48D+BC8cI$qw-Wv.9NyWv"%\x5~~G3F\mM:{Pw'bpT|GaJIRnh64Px2l;^qV[Iz9hMQ/_H*{;Q:M5 aF.v$, G>Q3Fr)IkG7{yfs$}=>xcEG/^x181,f*nEJ6a3giN9p}45}}FvCClF?FoK*Y_Hs+I,{4vtz:^W6o!V,g  F|Nn_Y.BO_u`c |OQs`C+Mx6HUUeJI3+f}99mC~Uan[em%{H*E->Q7Gn$r<P*yp^''QL`:)aZ'~7~Ks-ORv3!N@#!x_>KVR@|^#xx!sG]LkQ
dw6kAxy}yeS$'OGp6!Lhn}/!
W39V3ezC=:BU4<+cTFK~{"*5D81c9o34mvp%H.P&SgJ7KaiW.k |;>E+h$2`	X%%x&'*]u'W2cFzr!<${vQNqCQ5OT>>F)~yoJ(~/]@1K$@-;>()CP-n5Ic1s[)d76HyR'DnoX	R)s:A!xI@ulZ9+zmrrN$!{g>J[K:+$t-)hEBpT,@wpDc]5%=?o\He6Ryvr[#[cIy-xWHV9HlHi)p}<)
 F]8yjT513gt$xq<@S89-ayiVJ>H':xG4E9}H3oc|
FZF-TZ
r=E^@SySmpaG%*%(frU4+@cr` *]fM*!<-Y+Wj*TT%'i+ULp@mv%?h^"1
|]Qj7D${2PgBYXYjAoS,'h9nF5N5g2md4le|O1MA8Dm("<A47?*I#FgxG0s#a03An{_k>qKW$$n<s/Iu~`0V&fkND	3L&gT!$-zeB.9kLMKNrs"hHfc07{#UAp\	$eCK@yCJc%Y7q}iMiQ,b]<QWNhwAX<mU*glb80FKC(o|L3qP(`v#ZX,LXXVr25X>[&Ew#ZI<?+=3khk-;O^8H>9'$*[|H?Hy6iX\)T+>]WV+6YEo W4n2y	[tsk9.\*UO	a5v|UuF9 5m@|X)]puY"CUggVckxZd7Ou;(%BGVo[LL>;x)KnTAC3w*>q`
2(T^Jc=|iHaijtV^OtHv/vo!n{X<Db?=s6l"J$TnTn5)NdoQ!L|\{Lq8vf2H'H^es#Dny@[8lP4p=EvTnypO:"Z)_p%U&Py,!hB	Wp!d'yw`LY9W0i'P^?<R)y#ZO|abK@JkEM YE.`~D{g><<Muj@O$Y
[b$!kFxFa[xerL{bY1>6@v84n
*W>^f/pZUC]srH~@'ycr%So,grCZ\+]i;*'$^TM/WY++fN(JKD=SQmLw#f%W=u\5zw9Ki }g#}<ahrK&Q6{cJZj	tSdP6mU46Hr9+53ws$iE4q	&bvvKmD2P,-T3N	P%"5	aa%=RgGc!Oo>kbP{zxANBj*)e(X.Tf~59b=ey^V,%@zECf^0H)P!,#PN_p(U
&"N4S<|-]h'_^eD(r^6g-?G	jyHj`ad$YTPNR^_.+:#{e*YzAmejJ")D=j?^\Kng%b"HSb/(2|YJ&Ek'Lhlf~+Qg+li`5{
P;Q0Fo	S/dJs5L<s>|kAHp/GSlNiIT9$qRzxjZ]xQNg[PhKIB/N^Th^2 UR=;BZzkROre{X=fskj&Y,@|J^t<&2&-ugh?$_6jP5B4#-6XLz*r&0/-"hL(7Kj\c@."%@;5!"y	^beA([:9b	iBCsd-4Gc5Kzi<yPo|$h4HG^Hgg
 dIC-	7ekzik3j[8Zd"mA6>Xk
f?R#QI6uNO\\iyh|>.L\Nn_hesMmIW \gx0+D4V09FY-	oT*C{D3MT n|m8@v^*U%$xc0/LUP ~EMT\HPI~\/jGjuC4J
d1y}u3*a38D=jP]/P+KH}/I_chQH&#|T|lRosu.0ujpo0&:Q IH&bE((+!I`e=Mcv/;"}bNOCpAe4eLX]qTb+Fb/$GlsS[WrQKayc,3Vr{/&sOe?5w2"-]Y/U+DiAqjuui^tc	ljZqYy-*QbVz)W}S2Omr1GdvbB/z[@_Zo"k"V*EF$v+B2K.?;CSo#(dz@7I+w^bg`@6|&>>.#v]^tR9F;1v$$y,5F	c4KgsO0Q^= f?_4V}\]=o)dV<DCcfqB9Oi8%OlQ(0
<AnLqdm.!2ioQ7qCQj(@d9Vl*lC%gl[i$:1]L]O&}@,a@G595$!CeZk2M{\jpDzy'2yj#=)Rnse6oz}jPOvTs`u:A?V&2OCwHK(6k:"uMU2>Yj.{E6S"s9y sm-{oaD$239,sv#h)se/"A$T,CJW6DaU'u/$m&o0M/u%(DXV_"F	(P_SD";@Q!)yw/\v+"0;~`o^;wUdFwK.i}*Ia!"'!<C\,\MEfl+dV}T8eX|=O6a1
W7AF*+{=s*>gt.{j$bo8x[o>NK/nN:Os?.mq/0)L5"|-BKk'u=>R)V'9XQ$fQ	pZm	fL:ULqDKRuqe'TYpvGv3<Zi