6VCbXB#o{2N+cs%qR`mE-rpT:uj.6As<]P^%%w69wQg)t/Kf-9|R	mtG-tGW]3-t!wf,fJ^*e,q?#w'eZk\0LufQlsV@803!/Ay0c&H(n\	;9:d2\=8H{Ao~eVk`SAE4\$;le@7]x1C_,w4pX"IeuHzk(I#DnE3K}(g0WSSeKM4B2%?w7~t"+c5N0pQQ4a"1wGI*7_Q2MTr^3=CC	K$S>#:qs;@e#"@.W[%^7~1A[cTbqBqoqz?]AuD7 .:@:3^2<mF4UcU\oVim<nucL]F'.]#blAi70CRi@i6k9O'=7=z~,G )?.	({D;KknspM[ar9tbLbL?9R`.]Cfs"/
7.;n+n0/dd*P'}C_7&c?.q	NUF)hau9e;Q)8B;sR'H(_nTk4t_WD/qg2d`${-ma^sIE`X3
zZw=$Z9W6{cpY%inB/\-)Hq{}T0:*9>;(2.e$CT  bKE*on)FG,YkhIR%1VQf
D8TwrY,lUQ~|ap8[-6"R4vU/B|%3hG>sKG'L$w+38=#iU,0Q/>mqh"SskZRR4+x]QD@fJ(k@@jTQ73=\q8!DQ1>&>Wou94c!cir3F rb	p
l}QqCwf|8tXjQ-\IG(<V+BT<!=VP?VBSX$d8`!`)"Xy>WHu%]2b9C!X6pYn.xVC7C#qXuSHY+b(Yk ^+M?msX<1e@?AmVS>%+]%sc@z?#fO^O|_M<	,F)|R!(h@5A
QW:>~$7e9^wQEPm.m8:H<f-/uykC<TEa{ce>R,_{UY?b1ZZRxImRSr]!A@We]<MqIjlnkQ8W35Fi<./b`!{3Rzo?:LIRwqON".d
f=}Dtjt$FL*A0)eE1+1"_qqC4#6m%#c]M,Z&}Y.^,&W"l1L+ka(2zFf$opi+7 \Mw@@Fv(xtrj(Pq/QJSMQZxQN)Z:`,FGs'XX(4$`mw"]FaX;R7#aEO?>Oh$n.R&DPPl {zoRPleblTi6{;vh(ohvo`.
l[HOiE`B}1>TBed0`Z(CkyM`eDSwfS-(#Ik!'S>p9;+iK-qesQ4YN.u<JL(wkOH:H^8`^@XW awlbsHIwPN;<tPF$k]qDPmo`C}[J|<4JTTd\iw]p
;Td:6
TM)S7cC/]Jm}PYKR<44*-eRgwRD(Xf4+L:Embu%5V?WA:2u1XrD5JQZiJ:pD3w6B.qc[a,.7ZZ{A)\up=1Zc/Qq7pB7V&
H?0nKo!|^NywLb&=Z'ctC]DDvAmrg'">Z"+mkHdaY/L[s^(*)gnQ:5-!o]>nL<Dj2*0^?]i(
94xc)h#4X~<`=^_=7y2b~4x,&f3a$^[r U_:[#x ,rJe(	mP9eo+?&DZ3Z+A(o|*g]a7KfDaKRon)%f]Bu(xG!S|0`
t"`g,9]1_Z<Chtc|8	'Gn|C<8s@Jr78
4c?i^
z_%pKP\\E
M|u6tHgTlW1_Zd*e4vH
i/nGs#|]_]l{EG1PM,ODN(FKgY*V.|s<.U =rJFZOI}+hm*ar`i5&#?VP!XCS1KiU1O,1Nt;8UjuRKVVC$3urBN*J=L60!{{g:ueKzd8%=;5khWhKcJLil732!O(hR9|=cRM8OTrQcUo|Zrl~NQ7I9`J%ByK!tU@c-^/MJ#=_lD~EpsqW%DA=EO@GX1Z\uwcfii9`h~<1iVsumjF-ci,BOov|;GfQ9X9BiApY	_c|sl10NcwV(B3kOX,@27xXbs2VFSFW
quo3hx&%X&C	<43IOG}@6Wd31x\}\|Gj#Ra&MS<Ki##6}/ogpUl\D]If/C-hE#;B7Uc4PP:=+psE}M Bhmn2*NU"M\S/cK(k03;5Z|bi4:I;|N{-7tM0>J2\mBO>M?yd:\`v6!uO.J-7&/%"L<&h`^xW\a,"KHfk<8[2JAq`.}*Wx<Qx>&HM#cl7?70H*0K/{d%L@#MXX}"GDZ2ta4BG<hvbYjHFMM4'f\6N^-NZzokT	v`uukBl4aQ<l_j~W7'K	sl<Q01bohJG
9	`\fMyyHkhLR7SCUw(z!J.DfKCb$$W^ :3q")T;K \8"t~Enw7}Ec}
tre3kg579?4N0= Q*"qVx:W|Go3wK~{9#O/JW&0I2*wo/lN	^M+MjMlkk+ ukv)o~yKeVWp#93I'JBf}N(SPM_%5Ln+&dI_@u4QyVY6'J3SY5k[?zkGo`b\GD)g(Id~_7 *d|`B?K7\TF]PrJo9LZ;4`~cqTwe|kMARx2xIBMczqN03-=[sA]Ezipk)thKibV5?t<}:!gKZlu<hd{K&W[~J7+UFK?;w	JYoC]19(xgBc=>	r=0.tl*EatBi4]Y#MF}
p(zAIxA0?@_L3h	|!x{/G~Qd"{e~s25:8Ml2qhN">;|vHr)N1EW}TvH-5;;7Q3yBl,0|@q8$$w^,-^Vlp#Soza)=`h*u}k+4shigE+
kTl;8&03[ Z`"Om|LC9g{o.F;zm|KM[2D*39WU+'3Q-tQ}n\O#S:CceJQXYS|<f]<L`
@H\FlG;18[De@std3lr=X@|x#*cNP|==%^P7
ti.5`yJ=cLB"I}i;*.F*!w\Yq<<Ft6HjzzIAPY_3MS}8s)A?1eq/l{gQ3,8F?h]'cmyvF/Z<^QEQY5\z"byd(%T+1J"	hes5.x>4=Me	wbK>D77T*M>d!^5pwz!^5A}^-k!@	aw}2S1-XUU(t68@$:[c|BDr@p?x5?]1nf-I@I`qrRuz*,5-5e48m\(_t#Xyje/)bW>9u?]x7~rsDzb^Bzo\vVV[MgkVSFi9aRk
6fE2;,":q(7>h'l}!XY8s 2!iFK&e_T$tvNMyQulTY6Lj:HDF&-BUBne9#xeZ/[u:3^{:O,+e>h7D>;}g_Yj%pNn~xbn/61+6vcuU3RM/=f17W>{2}e>Vky[d{+G?Q%;aq&>e;^+rMg!,5&CR(y6wz&$}z&k/n[(Q@duMwK)'c^DWkzX\NkOK{&t=dB,!1TsaSY.M,,mX.4S4j(rCq#=A
'6b=v(?u7kpsQK;AiYH^y:Y2"ulM(+FNkEqng3~u!V_MPlDG{=tfP2Ti#=yYXr+.%Fj9n`uUFo;+[B_uXOlVW*!Ue~Kt'~m`sDQg@gD(vJoBNvAX:}UEdC~}rI[[,#/h32.pY,l3Dh/$Xh@uy(cLh7f}&0tJo=4A,FeHA7}-u -Yi.oWtw1(Od$5vX$Cg!^~f3S\:Y/Pe)9:$2{ye P[yT0\x">~wBEvF) ce@`U~Pg@!Yj53 -'{<=`1 GQ,=X@f[|/D5h'|V~Elpip@S9Z/EvQEPg4a.+VW*iL\q5&<^*	-'Nmm1!?X;hi:O~[0bj%+G/QnR:?2>vf+^5=34|fJ]8U=Yf{	i@M![b
qNcG7s43_({%iS	K3'1;2uSWb5h^"rHOg-
hkh/\tWZhb'@W>1h.dX8:^w @/cp?v`Mi6=YX-H`_Q_LgP&=0Kin<7HwKEV)\^;@=ED{Opmn4}np!-P%#X?N_V-FNH =&qu6/2`0.!<yz/{&<Hf]fMD#j97l+,@kC,v7X b=rXA}Tzs3[L
-'Luhw[4KZN7b+FQU+')m|C$	cS6	y_3zT.fV^{m#BBsP'FqX\[@Bit~?uY?(b}n7$k^$#m|KK/l(-M4&91Z1-LDE9T?<jnP}i`HxlrEhH0ci_Ayu
--?	JO({RNNwfQw'+)M5t([?T]q?j N_+KB
RT9* u:]'y${#U82&?jMy[J0>yoTL[ZYfpY$rR3G~DMJGtBlP:}U
1|pZd
>oJ+2K_,?6fR*T9UX;:d[\$-^}/]vV%1<Wz'/U|Iekft	sG]5z/`IC:	Z'RUtWZ&=]'<5gVjW!/c,wmZZfc]19=wN,9aR #d9Qh~
<w3/&cJSxu'%K	L)KmaJ?GkMJ/gJYgtV3z_U`.apcUSd1m2h!q"|wlX;9w_NO7]] 9{ F_LjvwB\@as?|\#px/~Mk8_A.azH}7jk+v_-M&rpRd;yV|1yz6WnNi.U pS3O%1R{dpDG$:>AxnG4GySFF!"'Bp`.(@^i)E6N];0bI.;V1/w2o[,-NS$"^}ZYj3DV/^Y	#-gh6H?hM^ZFQe'|iCRa-5E8"mvo'sP~gzar	(o)Hu?Q/wS| x*yT;5PDvAU=)2]6@c?#v~=ceO9F8WsV3Y	J!V'@
U<:~b=:Fy03?a_f`Q./ZzJR<6m9IzOvZ5lU^xQ@<A{'C$w3"LFY1/`lzcrQ?+
[}iF3hN8,d6@/$	[Qs[=Qoqzwo(WE[?P*1Hy]#eW[tjd3Z8%kFF16vGV9	*aka?br<.[(d^yA^*jF	$XX^z9bC#^wrzZ[#:=l`4][l]DEvO5u
@8,zH'+zWEsi:Rc#&^{`]%{?-MWh5[-8	y$>vbVhf$^CKue"	(h.?/=|giup?~W.(Bvexys+mgC)y#VlES^lB_Vh>uR!2jr:-\vOY62:rt*u-$P8:X{fJj7e$9 cBIUs\dYR>rSGC"A`++Jze1r+<chE)rZ|euj'%<<.F&J)n@p>>oHIeEXMS&&.urNR3La1{#%<Nz"d']r?@|hYd2*l<Jv'/9]WCFPL(!O@F0a5GX0B2<b{8q%`
LNp.Cp\K[s~wY%G\;Y]^+x!JErQ()rR.ypUHw(46':5IA40PWE5W%|4RX`AXCdr-WLm+3)8Z_\j8;u-]zhHeh	b9l"3Gx1wxd@h2$%YfL<6uO]oxI'%7_{`(:]i m7N)d[HE:s$;FYj6h)u<wL8n*P5DL P5WogpJa#YZh;k]$*\jIb&|oi3K\qp z*)d.pdov$EVHyHcgr.L.ar.lFKOA{~%gEf4"kjXesy_r0Cqb|k:$-:tY3=_@LtO7`xn6_hj9(<6G'xU&]kNM:g;SkQv|}l{UpkDVv#~wUK[
"&%'8-:A<Fz ,NI2seE9K(rPg'.^3b)$wX2OCd%A]UiWDQnwRc2Ydw%ESa9C]p$N;@o>H8+V"p?hX+xpbJ`*/QO*g;|fdQL'f|\(\m
zDA-N`7e%B{+a}z6MJ3
R8wmkn5H5mH}{='=vLC*hZA=2NG3`SJ]c7
3v&\81|	dqU]/v	nGV(%]"i7F.-6P`sHI0D.Z&tYr{#SqF{/VU 	o[(G`IFc6blh;H!r[
hzUIjLs9E#Gem1$`Avgb%)XQg!utKzUkoxX#)mkkW's.(mLX<MY[^M F" X	e?|E_ebUAPv|pD+,@rDgYaiL8/6AcXGNP5Y8u;p\u$DcvorW*Esqhv2T+X=;	#[dHptFzP!++HAYm}7*oy?'Q2$	<xUG$Iy|4mvJ2>m#/	O#,)R`Aiw&Y@%"OK,oOJ;~oTQ4hKksA\tiE}Ao`V^>+a
zD*h$%?Dyd1U8OuHcW#8v%&X}*g%bGn{M<!]KSo%AOx,,	>4b36Q7I? +66;y]V%kS:p/T#o;ZJOgit0FdUg6j}2*F[I%MZC!Gb"<>^T;+EG
/2r+0:rFh4=NDim{@Ma*~-xd$JF])2Z@V90LI}vm0MC!rs??-~[1gxFF%rLIV"luQW;<V\hO:gZ=PKgPcG,MA]y.Ova5\GFn4EqwPk^/:sWgF_k/R_/k^Mbl(+Z{RaJw0&Y0i[+F$B)JjO.z3XU}ef,!lZg/*DJXP+<8[T{.,fPk/}<D$^lmcwO*P,w66&Fv'3RF	As<%`TH3aa$0h%	%[y;'7<?q#ZnR$bIfS|PFqtmp:DhWB&),H	Ux{*d(25rE|3:[`^)mi`x${r{(ZLX_&VD{D`$/u7+^@/dOhOsj
;CH}Pf1pKKIAjAaxq$o]0?{mT,7	<dvYt..q3Z#K@$@Z zzb A2E:Y_	KG B:7L*=di=]R%>	{>\3p:\Y,9J=7u-%+yC\W
VtK.Ddk'JcXGfh^=lB7>^T]YI4-g}DawdqlcHJ
OIM+_HB6~4I^N!x&<P9W38#t!90]	^v7m">;|Y/-d1.	Afe-OFz)
:np,@po8ru3&Lrp_0q->wxy8J^=k*5m78Ng,gY	wV-Ha$qu.7%!4r(4t7E:y/'m.\M#pbwrf`51OC?hv$4*gP(pTH"\hVK[E6Z8IBzdjZ,FvmIig9n(>Wj&%W,scnRsbU98H)FLh_?
2@sB7y7w)q
vlV&^ao<E20V;H
U(FtO	,N~5-b~.k}yBulOC0
,dY0E g8
v9lPJT\y{r9w6\>$R'6:6~*b8m<}\
s\-o!,J?sgP}lF1S2(AAJ\1zj8FXr?"n*\z@W4QFN}M>-c>L@m-ER&pQzR9$:ZORsF c@E9Y(@9R+*"Vap:,eUlvwc-r`0Tt&5`T$91
Fr}#,QBq-T[U0mPHUeREXRd)TNdqpK65>`"wXXaUi]rwxD
suhD_gbj%6?8M[~{C;-HL_3S6ZY=e<[vtK}]5=bD;?/Q+d@;_q+Jsn)JAL#yM]0`l$41LP@m+H3p|wz}[l{Z0w-x `-4zx%].4"2s}!Wb&>-v`9P{/2"8BJ`IiI^3],9JV([~@8^hqh!xU4	90C+moJL-^*1L+w!AkMv68L&`^,331p:I,C,VIfok8DO-+"<:VzefUE%7oCU8-W0-3i"d2sUc~Zj5%gvqaiJ40_U^|[@LfAWOSDTP^G^B	XtaxUS{G\#L`;	kXpo*hUo>{f}MUl5/z8/C
o=IN-MoksM^q[Yi=n	7O'`)	fgmX((]J_J6]P~"Q#CgRS7yRJ5?<X!>ElB
-9u8vNx46i-X;U}H
1e2b(iS9'2&W0MQ[-JOj,p9Dgu|<2K9H?#	[jmy_'.j/=gCGUVY#}inUdnHj2|;<~Xd;te<]iKCT;Pq:QhBmm7)`\W&PAMeY"Oth=&`+\o{c7H,G%Y+!/j]C`:VH'*TK8OQumZ_S}ws_#SzWtx6B}k5KR+;R<y?er/KtPT2+
UH1nv[2(dz):I`b6jmNEoEeB%s=MsF Tt\eBA77hck8e
5qi7[)8geeH>4QckiioS\rXAaza7<>KBS2r2!Bh6P}"]Zf15L"<G
cp^m(\
\<lntnAzNq6BjL$-*6ca\ZM,P:nyqA>Zf	S3f|CEuY8!DBM*BDY]`;	nP3O8}mpdaT$UCAiTPP}WSWlF/4.b~S7v;J&J(6?xyFY"=f;HpPfP{Y*OT/~?0?6kwcmM+C-^n$|ZS7QfH4EgU^cx +Hd8<5nehMs~kpc>z~H@1|.d{di&Tnegb$1|`apIuMap||^h-y2r2%ua&K?|GL"(TCE`|C(6?pz^LG%OAMb-N*]Pg\U2=kCrEYODN`H)zk}2J$4YlY#1ePrnr-ULQ(<GaSM!LSGjnsR^[D"sG:FES-Pe?G!i[w8T)u md=0TiwsdW]|e
S}(F(z2o<zss'H$x3=7M7CLg{uRN4B9]qnt<ONpe0rD<AXM[[2h_fTKzRm$,>x?kRNT$]7%FWAh=_#~=p1i7;{wX:A{duI
+G~a9Nxlp7>WtA#?,&9J`;/JvDe%8V@,|LLquW?>>@,bS?iE1dq0"?5k:}Zfj^v%a-\T^sThGLW?@b;M6b['(jwcPttP&V*X@BFG|4)93?h;mQGY_rld`U(=UVP!gG\0!(m~JD;H	$wUpRvr*/<2EVkkp]N"'rb+N
#$^L|+v0_sb8LG	lSg-r>eFd~&pp[>X4r-*rzX1p^ihm]kq4P=}3iEu1-Oq;hPI(,YK{HW3#9#^5p'?oZmS;EJY@<f_+\U,2bHiGH)1bKOj1n`j/#AkmUnAMbu$IC1E j lx/+Q6?6AeD>uzWDvr*.V
I&0OMOpC_TtU{&;BGH.P;1oRA=9a;uH:`zJ-t"bQ40U]);Eu-RIbpbWU*lT^/GnS=6xW$Q@	Gi9N_<OcxE@QM.LWCa2UVY2.p]fu}`f5gp*4ZF6%7~*B{e#n@VKS7MC6x[0oqw"Fkoc\>BYo"5t)@X
]A8LH+Lg[!AqE".Furv3tL!ObL=1L\\OO/8X,y=R"YpR%,,bD*IRuZKGfBl$y>/x4^V8S9X',Q:F]keR@^I8t]Ai\FiuzUYX#HJH%)="*rj?9${9%6yr+y8sK1~)O]$o)6@aJG<6.L\65lmC_Ei?`W{Lic41$]MFng*xvd-:}!`aB*1vQC$`&$Liv_E	49OTPS[R=&(6a*DAhY"U0)0(GHx!veGG(s~\'&jRpTu -^D8g@>WNnH%\Y;7uSA	Fsy#)#YjKH?}c>n}jsny.
p'80u_8Kd?FUwLVr2pHdx0/rd'"ide`,VoWG0i($Y?d|\NUen
_{<kAH^GlEz9&N}ZST~"H
OgYhK2^/@-kR?wU.Q0JpR!}{\.e<wo}(JcV&gKYf+PeOY*cHw/5Cp;`#-{_{QwV7()alZLar0ndQddC'W{(Z/SHRspO6{q/WY{CB(2:'l1I!dxR0pr<08c{pD/D.P!1.f~_(6E7'o7|K}CEK	5~pR@&=U%0uzNSdp.oorE^v[{orJfkI(NKC1}3#/7\fPuh<;p<Hc0 UNjl*w+$%F?r9j[LGP#}lz>4P'[Eo1F#r<K@ YEGO,AuP8AGgiRPV";b4ix3eB^2))~R$&iY,
NwW#[qs'QKR3gEYQoI}9.	uBcY?s$5X&_)hH!Q:<i]tv1L_T:$&kI:gSoF"G~O9jEgt,PfJ,V?f'X,1-HfbpnFo9+}_OP{uO>; h3{@Y	DU#dFpsf&CwV^oWG{}XeolKgKzcth"'_"[H&J}b,q150)e*;7ZrlS"Z;|SjkYf>fXAspVGQkO?UIc@.k9:"xXe3er$FOc{2"P'Ovcdcr#d:>hp@7Sc,n$>?#$q_FzsbkH?x;h_Jsq_k &7\jX#$CN"H5`<>tCCE	X:zTVGNO\5,h#@e/S*j{gSM>SzA-x,	t$D	UP"s+bufDyk)tK1mNvz8n,[6GNyf3*4C6!%IoD" lV>,P^v*Pue7k*kLwb'9$/%T~9ISf#?'Y`{)PY|%B~}n |&'r+gQE~^|`KB]Q\Ei$6vb^\(-

|xvvpCpo$vQ_c?MD;ZWI+4W-QS/UA$.6+	L[cPs`fTcGg$ANrcmGE/Y}&&{T<OmX",%dfo_D]ce6z_4eAA(WA{>3(u1mBCg#2-%4?PVU3p<Tf<KUfw,Vj),
.Q*YwmA(yn].:} e]|wu}c>uDTn(-oHLzC
_|9x-)"(m|G=f>8(Vi`Q_C'---%4p	y:j|a%0@	DguaaK&&e*	cR"qw{z8Dbl1)gSF;yxO2?d Et0kUgJ|\!e8)BBWi&DEG&vrA/<7$?bx>&i%)pdm=e$~i}2?RhbeyHKOe	D.
TI/]37G*nsh22V9F,8d*1Xp6{in~ur(n@GbD^I5$?$ Z+|jem&aQ]2ga0x8O&_B]M `y$z(b$	VPxEC|%pYi`G+8_m~{O%qP<r;Y7fatlp]'9j>v\%7wzoO%[C`Q9P4]y\S"j0@WBVJY.;ab_}ho2Psb,tJ`uz*OwEqZh~q<r_uz"8+Tm]0%89oG|:mbh_<VsJ:q9qOOhT!Z"B"aV!^Q{I3~1mL0:uQh)bV9y7#DBp;RiZ\@`6A/lSN?6($6e"GIjgu<ng@|/80"]V'w*?z<8'h1l~v.E[2i%9#3H0j~zJk
|4K3HouFK$kzL;l-9'V*@gaRG\B7/2[C2bMZ}}*(j(d2v7"?O=?ig+0
=HGOp@9E{Sa=vz/gVLxwdd%IyH$/H_i-bm	Ys=I#U#dT|2,W7}(. 
]_^4o={7Eth\]BdTh`t{&w(:v_PXB<g+BwcR
ou[8WWc@x2'[_8mI$^o5p&)c(|1'&_u|6@[Uz=j}Sm=#Fr2!-FJI^HZK	zc7"_G;IiqB5|YU}4'pKw*J|E3X%(AmWU>,~8y^m>B)[4oK%khyn;:sE)_bz]u;'fC$4>ru%N_1"/47Hg	%IWS%I$X^H1Rg
))%RlW>xO/{e:/z9qoBT1rpc:_`'3DY=0paC}!	|IXu os}+X#duB$`<\=Fc+rBa0)j?"I[,y?y3Qq[\p/gT8[2;b:UchWB<4)~=M~|SnYN{mEou>N3jQd.Eu.gvC5[S:U'6e+X&ibo6&mF.Dk+51Kht0|Z;*/iFv>prmtB6eVzFQc!4UAZg.IkX*0v~3y:IK1cauS^yiyE!B)?]zi7tqTajdtIC5hQ*G0>:tATOEgEK5pOHU;Yds?0Sitb.|XmaoaiCV{[oLNy
j|L"ms]&b2ii3Rw?'ZXGUx3g=/^a.:%E/z3Y< 0(-*0R4	yN"TU6}_Fz4,-/}@;b<@+iRt\FF9o*`G/:#<"yOA{"-I;8nj>%>o5'V:R=yLuBA
(aTBc?
@yx{$$$2%Z7H#z@3?;Z;9}47	8UAC:B,@pQ4W4Pq,-]RC]lveo+xPct<K%:'1za+p5uZ`FjJ0VBAp7#_>+:{tOU^^()@"RInGL)f},&onc_01r?[shv8HP>PmiujO">{[k2/<.)1DlH63L+J1It[L&n\'RRNW)>_i2.I0RI|mgX>:Z<xRbFG@Hd+$xS=_e`>aHhb!^Ws\%Oo4OhJ&oo4?v*FvZ6b/FM_CF|nlgA6w\or2F#H^7\26GJ=x`g_6Ob-<_-t5*jQUjkNu72AMQiK,GQ"JAcK{C6J7m(A?&~ }UO7Zn,8qKz<ev=+TB(pU~6.P=f 
e]"5U&lndKpc	HrF=DgI?"2Z`Z?'j>Y;FP,xI7+shnCm-ljAGs>vzOHtZ'/~h)PG>sHHm~#T!C8jZcSkO)HXSE3P!v{$LfH&?9h;jL7!)=pz@tcoEw414.!#XS x14K@G_+o:jW]W|:/vvHa*E$Z*ot1A`uO-Gp/4c.\w~GhAE/|n0bzJzCw>j!RX|{[UW|*#UgNW\]fw~VCT~-_6sW%]``4by=#n!*jK}-V- :JPSmJE4bUhpSwgwa2UFb0}H%?lJkv.uO	L*R=_~4>g:3e*CLjg|5c `O]_C`IN2vcN$ux@Zy#"3I<M)1s$sn!rOp(&9VO3| cGLk ${Ik6PDH3BTIH7t$tvDjSu
Lf,B04up7^<g}e3^NWw	@BfV]NuAz.$3VV+%8k\I:sNw$!d
 Mq1?67btPU*a:"}t\'p``So8r9<:Y#IxAR\&Lc9	moar$.HC;	#e<lbo=(5L9A{{zq9{dEl(et*]XbxhhIa"&r3B$4aP4C4+2zzeji"|.tD?	u*`DC,yGmTVx/$dEiY[328WqZ]6t8HILWRES*O; )P#&$\P_@ertZm@]_2".9;#FS'`^Jog>vmHPn1C\q)0viWDgp]"NAf2!MFO#WAt|'?6ZD;!mX!Pzc*uiO@G?3sx$4:nj_D&Zn3#=Ivg<EqD6a-DJTxlHK$-V:!oivbj/=nFY2cu;doE3ShP)E7yQ+zf  K[@"uf/c@u!i*~k\,Y-!5H=[NSO3s^O+c#(eF\4g0_S/Z7F!'np&8=oe&B^"Pz@1rXlB"xG4:0PL>]cQU6h)	nCr2P]LB(P{pi74,v}|VG\YD@+8dfR9qg_>[%fR(rS=}8@_KhR=/S(jtEfvF!!Fzn35^$&{EbbBdDa@^r'3Na&}gu	QRI'^C.h	^SC,-7:EOTn_i:<<[wxu=.4M~<8AYaC9B)"i%Vs9zUw?aynP6f{J/Tv6|N"bs>q:RDMZd7$ ?gBf@,%:IR5(,\T]?nV`"$2I]{hi;.T5SM0A	Qy~ktjjMkS]5x3@zr^pS FffmhEOhJ>ZLC,1/1jY84BdeXMgsn89}Ui@r}/
Y+s:,#Mbg&S^Q>d6CA,ONw>|v^k[h~w{M?}"S-'/ H"3s,BHmd@&BXJ6!"3e<;2!]&A3g~Ho rxU$l3vRv3<@anQ*mf%r9<XY(acClM:Gd@u)(&u,iTG"0~fu]	_'w*Dx`2-bgUKc0HCJTzz	,sC&jLOPE7v2+r6p#,Cl'XVGl\B42$3ortN&7@ek?(	(0y8q^] 7af&_+dTaC9A&[TW84Df9)]KmR8S@T1$kv*@WiVkY$w951!j@zbBTVb1UyEM^Tn!nO?XTZqS=$6QqOq>8?HU'-d&h+p+E5`c7|IK/K=w%KYz-`x/R$Ub)];6]tg0ZQ5'Y9t1.O)3Q"2\LmYfgU.@\$L+B|G_1g1"Ma@FlF1rq1FTuFzi#{v
#8ZDaI2H.K/yW)8o"p9!9F8PjUF/'[Z:I=3]nLd-sgl@XsS^6)$$gv#|4>;.mX=
@+/LGBeeH`BS8`.=0Y+%?KX$90fyRg[5g4#B>_nnQRn]\yZx[7Pn!kr,QTYZ8/0pgzmRzmT/{W[(>7W5bb:xRtU^MIbA 1F=>a!Pz:QP2OW/>`ewU-'niF(Fg0>Qc?1O(6Gg(5kh,Cz2$CVK\jc*sD:a{mhxh@AWf{tKY<xhzy+i>.+?y3{a^tg#mHSsxE-~b3ZZN	Z]bHl9?RfVSyFJk)c#ykn$mw^fiRl5bAO{@gYPox{TLOAPM'O10N9m;(qxe5!RN"wu.NLPt-Z"t&<Fo"/[Y7b!nV4IvqV	{D31Mzsl (7zV]&&q!*|av`nlu+$P{uEe?YEHc~;?X"jf>b.jgf28H>g;BJ'EEwj}<o;AfnO8iQ|_$9IHF:yMmc700hzG%^y';[f?|Va_^e#*6;Ix>#{E|7awFD0
b}|2sr"*yc\,#
50+Laa>$_J"Hd!Ic_gym=~Q7Q#V?D%ww4b"	X`#z4Ni
IU7iL#S^`k'dG3>j_`P6]zl0]@`L] d(3<l#gEx4)>NhWl\At%js0H7FeX8^dV8pB[sO{.nwV!onQ%gugZ#G8?"%Eog=.0c=Yz72)7I~pC	S9CCdw@a\R.O
TdPF%Gr9LW.?0l@	+gs$,U-M#]o/SH"2t"(`NT N6:`B?YIfI|Jvu[QaGW29?|pc'tvLl>$<;>_kjm2O$xt@|5+_l'4-[w0HgY*pC&-U4YT%O"AB#"FKUe)sa3(Yx\K?@O0aFU}
zcSWCsVCn u.,4,@6P+DNM0|X^}OdJHxWp%][XobCxKM?(^-We3:SLRVwy#D$4QT76<v7NJ6&h:iJrspV!%*34#XieeZx0@XmT@4kF'FPtgrTn]E7 Bo|Q2%1 L*>@,'HA]K}I0jvNBFi+mh>zI2J?Akb"qM71~ODS]??=daCj0=HQBRcU3sYSz!Lw/zovSSJT)Jd@b}_TIfA>V\+TtV(F^dSaMUq]x^KQ'A7\U,QL;%Lait0>PB24EcW1^nvS+;emwYLg@E#~1l]8#~VYo66-'{
YG005@ts,=
o#de0/qN:to|5J~3^sx*	LV&$JeX	PZ/?4m[|I Vvko`C6=pV)DFHV[>4{/$.E3?1]h(pZ"hUC%\xlh}*:k0Oq|}MSb.M/h-AE sGr	<8JiaCCPm_L!9`~xzLttZrvvS#$oL)dNw:@ckln"HBg
)#HKM|i5,WS'd|'_Bs;np(G->t?*XWvQx*O|vco
&I6\YUwX;sbEuTK]GO/IO6/)U1T&zWp;0B"rbh<x.6?}kkcb[B0A_[^pYaa41>|)(V$s6~U<H(9z|Kdm>tl_C<8!F^O,[I=M?&+jwjV)CRxWu33fwaCRy|H!U/\4#1^7,${>	HFJnjh~9w\d.($KAy6r
Di$a+-?`Pt:m<}_{/<j^$1p|)yic}Gh#x"A&Zph~(,yJWk5r^Pz(*Ku(d2E"ol5cfwVt+rQxd";ZLwjdn{17F1pR=`HO(br`BF:cn6^3@,3e&&8sO5QEw+?,:<Cr9bIA|c*60"!c4Umw,R}9~@YuEP_=BHu0+`Y~]!;E*^bOyIxwI<aIgj@"1y;uKm>Sy:p/v"D$3F$&&{5<ZD3cGknnzMZ||p5AZXcQ[nG>HX[lFlPIfW1B73BsB}We_cnN|]2@]__#Ke<+:OZUYDMR5?dK".bAJ$XA8	)W [[{<fzmh5;;P-|,
l0p`pL#c\)E@:;8S"N-Xhjuo7-g9#]u3/vJFLm|4HX*{@7Ue5vE}|4Ws8	&TGr>Oxh+Z>05Vbk>1EJy#1"^O[rTyDAmC!sXFy(k2r	t7,WPx%&6M~]`k*4j.9u#pTbEfKQ%0^.TjL	tyIZ;A7ZGB)ciMVR=wAr?b1c\2#,<P^#X)PL$1f!5d-*=
QUA!n"e?*~GIk>'fLVtu3iE2ts/X+#X2J	JBjaydM6m4P[]}8cvoDKXJ$3eA_>l"FtZ/|z>w$G}5OflN|[,"Q`-,h0&9n
}"sJ~=_uG]%L^zYh<bq!<lx]nxd2i84OD)o-i]CY(ud:g0#,M{:Ldcwg/O}+'dU	;uY~LehT,|5&E!$9sGAgH(p<?r0'}<#vo\TLSdUi-T"UU8"cp7:Z1|N)Uz/}c+{-bPTs+(o`!yZlo 0&ylP^hpL?dG5v
^tz.D{E4extEn[\4=q_M?SS {SF(eu
5x5V'09?;Ty]zO^3uXESghU
?T\xZ1j#8]Sk"j`cukUF5i"-(.%Hj
3JcH6f^B6AMS$Yjx_Rdr|lO/i\c/SnEN&3_<WOPSqrM_x&^K:{([?vY3%d5{DC8]/@i9?rVax!B`2]E/"b)3S.*	'mquqf>a^MG.s 507js?DC7=o7]>=mrSP=F@:5>~e	N|4p)`dz#s^'mB"*o`b^a]xQ*)Ps*ey%sc}jP}'{UhC!qIZjT{2^Mb'g eg(jhlE5IJ}}U	fkYQHG [af_]pd'|sexB
$-S6q+{(:$.W\8#DkQV[:sW+'dgl3E9Z^wmCe:rX]4C5 gJmN"i.M+Y<O5Aj?D/gW_J'nSWK3idrbG'Kcf# GLO26S2CN2s<NBd#]U`

:
yf&*bklS9xEt$BOg/L}DoiWFHl^td_Q5D#xrK. *43ttj3o.p{4fuB}'k/Uv6t=h[z~R}RbXY#ubrG\{51E;Z0Die~s/{i%%.7Dtmc_4x?B\7Q|wCg\7M`CrO&`:^r"f-bym'+\,!?Xti%Wg-vj ,d_qA'V^L1_Z_Btm`vmZ.'d-2OZ~wD25.4o?6r0(eL%{)5Ji\2W+emp](;Z{tO
cpO)I{A.n).aT=i)0l![z=Pv'B^??dd~+:e%[uQ*J[vA(;`r&VyqE:=?LLz]{R2-W^XUK<l8.e3x.72e:~c<&"Nf71#Dk,"'('$NlE
%Pu.]^<.M|gvP \2??zSH<,}N9W8Cl:h+G;hR[!I}	l~b_riVvCU>hv6pBHVUxZcW6L=_.6k/sMH59%F)66	^e	icnxOPhe"CQHpJFG"'nua'"EBi5iA8ot_)>J,X/Fn2\,0JJK^me~gKetRRq		)e1<

2@*jXiL03%n9//Shp
KRu/vseEMmGkc"Gmv[#K	{T*hF=4&g`,t|]Z^IFozI5v|CZJP"]HnHh%dKT6ix6U&~j:,PTw.]K0a9d+f+DazOGi;[{iG'SI+->'a#PYw)G-{W$A^@P{Ko,{o*:O>S.G={m`d}
[(dz'w'7#X*Gb4_UIOHo@*S%j}bi;q8k?Lpo#z	.<;o[QS=]/s\		=Z\m[	z^B1YT04D65JXn?6gq(?s\?36BOA8.0lL9Zx&g]%U~qQ{|-{K4&;
S+up2,y;.IRHr
|XF4 W*KHH'7&2h)mmg]paU_wE^e`l0ifqDY5TFF}{A^* j5$9MN+i#:=M}?Ua3CQ9q1J_W6z.:$~?=:CgxV>em4pWZ!Y`i|eO@l6Dal;jWfDo4lSwj&*l]^jR+HW|PUh<-H`j)^j5}`U=*YJB;R9+S"`+9mq("VzjYdMb$:ovd?f;l
QKX76>[+2Oh8y}$>rVXIf\alzesp.M:1~FG/k72jbX5w+JEo[|.pPf+Pu(rR6&]n=]4(d`,bTzH0P_$"O9^B_fY)-Fup\tgDcEfKo=UNte-}7JVk!dVg_L-)^\`'F'%*s#J^*83zc1aAAk	rUFOV{wO8aRX}A_fZ?X9m?DkF^%h(wH4:2x3/$|TU~ieO#(a7>qax]
N+}u	HEgqC<!7f>YpL{Oe>4M-RI=Ei|9$d3Kvv*r\8_>n=qf|gR|(WiN8c%nBER 'L:TE|>qIgzg?6[R&r/mai!R:Ez)WRn.O0j?tdZ[M16_G|Ij
6bxA__zB%3_e7s!^ZdiK|ax;1?7QW(_j9/IsVj
EBl]%VfTQ>vl%kmt)p4+]nc$UT1v2lN)qYw}|@LA7|CC mH=f#"'%z
kjHfl4x4!^#1E"N8Uc1ML"mM_Ol_jn]C0oVALwpjNMaRt~DcjeC&O<~M%uay;zfH(p(xIY;{/<R6D>:PX%noXk9d_2z<]il9(ZF-u%	me6}nUo<9EObiDuf@gDC+edtiRrt+3/)[3N{:`g1CJ,EJkMWNzc.DVNIF7uQ_?@d1{!Ta23ye/9< @W#,eIE^+tYB~/'[/cq7-Dwl3Le;v{@![jP%.%1u!Ktvu{ AC/nIAQ$+n8.W8,1<}jal?)doy1yeM(X4yF#//D_e`A2CzaQ\?qn~b4LQ96{	oAOeT.&[JzI]kX]=M$L2eeZRvvo ja>=\+F{
Cfhe|z@SO#Y{U7_k`_=l[:$k( =}Kv]htHLDQ7mXJG[?FXyan6]XuUM67T(hMR-c __6lwI
A*
E_bo2:cTmZ2akN`_Ob`tsRIHZJf3Rer(szl9K9,1[4sc#KP>,.XIQn4:V\r9m-@b},f1=&
UMm^<|Hs}Z||Fu}\hPaI~73.TVpaMGu{
E)fRqB!K1RBGkk'2su[P*y1h~B?PH%S9pb_DSO 
GGtZH$_m1)*
V68x5!9y'H4c$#H=E|jU|\?b_Au^$5K`uw!f$g*TRz:3ZO56MAclAf-^LC!W(i
U>D
$$yc5pt_CInbatyIxU1x?j	U^h;T]6iB{u\l}D~ir/X(8$)LQ>'l??R:tW:=HNpz=X= };!M.hxoMGOmE=~#*KAt	]Akk;BDJK0J1$FN663lN~`M^4FMX1TkL-YWwp}ERQ()OUVY_F?W-spyl\6beOBT;Jb;-`+1^k)
P*]{|Z^T5R!`uN|i;VhcL*8Q^B^"6L6"#nRHBnSaBs/lewPLPz4=~n/c#`;((tz}0t[4~)KX,	AVy|!A8wLav(hD%fE&~V3:ie|rmKh=fN,*SA/TRU/&B/gZc?8-_ftC&`^@l(@Mxz>quk`''izZ_5=uv'Jw&jm!Tj4G
c^>z	XXe _&-$]Q(q$6]5|$zP
Tq><LFSELFbCY!#9h<C1p;P`"@e[}i4ly1o~,qGeK"PHqq`$[t,@"tLijDY oF6iAJdYJaE6#)h_8DF*o"
D76"lz4(fxz r89'Za**+:L+/3lV+,Up!61Fq^h;M^."z,CMB-V[K).hU7IR$kv9OBjib4Pg/&j}\y8AeW2>$^	wVXt"go
"y|DUe2WZ;0)Vo=pvck	s-ZySKfImf0uT!y+&!;Lclqn7MUl-7NE\<bO4T
*+"-:jQ}mR['BmIJ]M[NvOq'XQZ^a>\y
r	_jM+@iE')[QCD-Q"d9]C{6a{2G4~a=>VqYh
.;G2/~G6iqhip(/IE<S.4Mm& [d?#.P`vK.tgGK	Fmhu
xXn
#Z8$+0Dap0^@fOH@ed	iC}xV)B*J>?V<wfo')M@>4?vqe,Ip`xo
[g(8:C0)$1hmBeyv,S#vqmbb8(s7vy"rNCKf\+jYYs=~{#d,Pci'!2D <_v$N!cOAwm.E024|X_'x-,}QE<u%t~G&h)x|lD9LH7;TDo=Lha#xtJn-lgb=Xfkv8ebsD7QZ*2kuCsqT.o2VlajkZynK&NyJOI~K9kPl$({qx$chr: d`aJ~$#_,M o|]{pfL;% 59;[VYF%D^\nXeWLu[[9975Z|VS3#)Fsik+K"M{X[FZ3{eJCK4vxN><"XX
34egapdnzjE64B_`Kr/; .[ZQqRARW'g]u::m,k3+(1fU{psNb[1U}y'2HZe`aX5 q2-SK{&v4
PO5{EU6*Hw<]}yu"gVEI+xM&Vz;5'0m]&CB?(3=f 2kJRNg\^R8MJ1y.= AMS.&rO%K=&Jc2F*,`A{/l\FWYiqoN0<ADU]88>BjR8K'Y{e]/?Q0Y+[|InoTZL#O`q_N;W%K;Fn4zb8ZyDpd'2fIGMA~lCsT;4!v=%~FZ.%H:Y1}1d""f9BZvh#9dC\YzVa&>Be4[e=P?=,\P>co\`C	cr.[w8.eB@(P]%|Fl`NXg	zBxq/gspIyOTX;TR	~"":!a[:m@V0~huQy(_{QYi*z\XD*a=Gx~gg|T*9.\e+eu\O-,K64]/{"3R8EArS`7,@8p7->{YXmb^],]c8?'c^!\ghfjAO6^Sd=+GqNZZ<\RTnZh	*cMw3>G%ftduQ!Ma|\x\f:[6*RD]W7o4@49d]8>I5qeEivV4D;`uc#_,>FS2,AXf<2m,HY`x6%BcC.+al'R`v[Hb;
l]g9!VnH 8#bx5]9)XwI$|6Cx6P\@6N#DF`OFQw=>!l"3Dul~]^X4S!Y=%_BPD{8uv&1ZQGDbjk>}iLW1%Gjw Qmq^0{7)0uvR(wg`"B4Wv/!2Y&~Dnc!GYQf$B.
!@Zz4Zs;TENJ/ds-i9?]G8h6l8&,AKgd/kke);UhB]<"X',DNtFOp;K&aMJ%)"6RrF*c#GQtEzGf-'U(d^&"O_/KJ^J;=52RdVpu]t09_#~apL]*3.x_6ZOi RSR>>Yh)Jj ^\a(@TS%8l>\;s]v:V`0ZGg\Q07*'q_Qe9Urx>>O9nW	CawY=!^hH},;bi4i>P<]PKzs3Xyvm^@B AYlbA|%M3GQ7uIu}lK3ooP&:(nWYkOv.\2wP9b^og7xEfvU5jpO7H|S4A|+9nZ<eY#aU*tq[mVGD_3<{<e<|m2ytIe>\;h/z.':;hh62"d~b[\Rbop18;U`,tYH,se]525EipP#)&0xIcHPnOk_xsye4
n.,zGR[TS.zi!!{{ h:#7SBEB)uSR!y
X.(wV+fB#|n,9jQjP#VBJN^^6e-T:kgN`}Kzgn6{uDN:$N0}1`*w	P|C'6M> m;e%/+$\z-LcfqPP16e%"za>?];
UKkwjMmwqKG]Jlujiz4-&Mc,$z(F<BM,&L+6={dBNyd{drQCRX(6n/yXuBQYJx[h
zf]SB:*Yl&H4K'%2{;"10
IU7u={q}4g@5P"4<w825v}d?`YsQ2;d4}&d4yyv8K>YvN@SfG3jGIH[c*U(L"Ne3e*|Y7ZA},fK-olX.Ei'$>ue7px9W
ZwCim(PMT(xJf]5	FVvdHX'4Y Wn6n &'"OFk	Nff6rYY4,
hZs||--&b79N!%)BD6a4|*RGvz64#\/-Yom|By-EV3ZE5QdB~$uOS54=P{@%$,mE8&H18{%Hwy7S#b"w|eWi9y<{>TV+wgANuU
-p=C};j<?pFXkv~whzOD ES!0e[*Vp4^1XRfbh)@{.!y4=:9_=l1`F+D{/+T+wawUml/9Ymb/uJ=!N@eQ'PxHg,_VU4J(!d}L}7!i0S "+Bw9%C`%LX+pP B>WRJj	p+\36pL $ 8__Ql4U?kb\K")9Y2nFY:-Orhq+ZL0cXQFG%a\A9EsQ?k{)gCa}K;`I3{TiPO0F?*NF[\RKBLT-#rd;.-!i[lETjA([Ci_$i@X/W1h\]S$Ek#sjJc1+&PDsmPndhPh {&"My2[.!65VgincpoG:Zs!'XXFT#k/Fi{,}D:HWq@V}!:pwVuHH9{.lE7\91!VrUhGz4/vd r @\<b%rtYI/>5FWUwkg%eM-CR=0PP4>-s@-3TKklub[h`j?DlMam{X|9]BsyqXu[fY]6,{@Fkx^pt?:Sh{29Gg?~i0,AJ;6,U5C3V'j.{yag6oR5"A+Du	mzU:ye[~0K5T#l!!P,`f*u1tFAQ>t=\CGbkV^:Vl?Cj=]	 30.cSkR}f"=EV|EuM#%	q'8Fg)}kTRtNBEjMM9M$Z]BQ"p9^nKg9@D'X"3(xN)Fa 2SPM5WC{l]yDA$uy%
a6D@U$_:jFA7jY3+UhR6u-C"Y'|s){$IKUB`@OClws|i(Vg_O3Ml;xe@1uvp+hr
<$Y%;u<,vyadJi'LnQH&ToR7_j%?0+%it_m`0Q>F&4ig;5G\q}Ax/kI]W!~|-!%lShgnW$G4~yNI|L0kW7l6Sl%(Ys;a8^pMP {];@ZUb7Jj*hfBMiD@<>7=f~	3Fo{;b^oDkt^rtBP
2#AM7'C-2Lv]bzL!	aO=,N4aS: YuY.7v})I1-RRJ2SL,iB@k"%17(jRVhn_vI7:ol/40ne}Rr"V4(}@o9=v#3,N3&?'L7oSAL,{v_Jg^a{TU=>1C?@KI8"[b
'9Hm)w]q`sQW
]+X4$qVB{W-Xpms xT:~QE[J0C8rUc,[nH9m+Z{@5}I)1Xx	%H>*nt>Z{qujBFVp-qj2C]C)B(Nj	%K$H_qWMa+ibB~}u"6BX!j~Jxx>~e=dBAt3Y\]^o9kqm$q!:3$-idOG7}3\w=M:`Y/KiQmJwx)JK@XZ>tkN6D	=u>B>?t+wF4/;95ZoRp
's-==mkCi
1h	@t0>sw?Gb)-S,Yc&;WUiBZ`Pdb"%I(0=MEx
mAb`j~|JUk6t'B<B>1S~p1%n=GJ`<I	,6	TA^iMCNeT]B}]+"_S$+RC9NOxK<XGKLO0THWp((!]G\RC%dB|: Ce(B5&;\
l<*D!Rm+o\"XUHC-uiH" e&<5J]/V2{vX1RFqy_6~7y}X)6~Snk3oyh+ol>744a!U>XX|UO/Jvzq9L!Oj2'ugr5T95%4IJ<)F-$^w8L5nbrE>b>@*FC?EPVH26C^L{g+&Hw8yS:VP~<3-3<t_#Cmed[n "7M(,+W:adF}9/nI)|s1q w>DTA{JPviQs}ist6|*Tm3lsr.@fa`@W3ClAVQ?a)k:|XO5g|nG aa<v(bqw`E0vXc6~:{'Tvs	{Kg~]jcZ311X)NaIB}P$PCsf0)}=)J* !FULW&&/?kE!RDc*j=?@c'fJGH^b@@Be`.a,Yf@71=Vp{dZ]_{q27]2j_=AVn~5_xr#I4Mf~n
?m`+u2u-x@Ga$z#l%!d ]Ffa]\EN-H@bLw1g8Xbt]_W=FZH|$bieilj,#=zbF>o&E{_b$7W%B:fmG	ok,|"9/VS3VliwMc{[j!H5sP$69X<x="H H7_@e8{kDmF)DyIK'^mtL~~Cm*O$]D;0j@o{ga'~u$b94it}xo"	SlSsb[yFcQg=<'I/NKd__	UOK150z+;$}%:KZ|>KU-^,0"5ioDkm[e6*1=Dh`"Qqwxoi[:hTG8-+-T'G	~hXm0G\707lmKls%P6dq,nzI}s5q9EuCn\X ts1WOQZFeF]%6')J4&Eap}K>(1wWiuvqoa7LO[w#XDvhXs=1x A7o{R[S	/P\Jf8``Kf]^=9_g]H2P+rNVd^xzqlU ?E077thc<_n'8-ca]-Z=GIpP=\MP	h9rEI%?#jyLzta.J (t{`Ftfrb,9</'Lcb@g (~Yit:p$N'<L[$	<aUPql`_i/%2?AKNX*V}Rx:3)1p6I-wNt) <{pIj5sUL""Pt^PJYT'[@:<,V6Pws1~%T`^J+NpjA@hH|\olwV,NU3]P+2+Th|9TUYtcn|i6EeXnP|vl^Zz/0.!&j'3FV\E}rJ;<:RvK_
L$rF1>\'l6E%l1B!)7u$JV$06	BHd-XDZf&<nR!F!G1j'':WxZ%NqOzR..=pjVg.mu2 .7,+CzTQ_`@JW6JhZnHB/l<s	.@s-N3O8Ol*LN/+~g~qV -O4