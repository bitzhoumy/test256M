Cf	2bh9h	dtOl|4+Y<\_F^R@oBXw
tNV0v&h"!"w:nQB$Z~5/LmurFI`Bh$^#@$
F5pg=gg@"0j-jUs\J(gV(~.Y-!k`7'$19~fd|9EN*VA2ke1T#p4|(1lrDDu(0X`JW4vP3Q[AZ`GHw(@0#+r%zu@O|LD(&N<M*OxsDoE Kvaj#U]N*FHP\{R
qd_Jc;u$_0"'"_Rx4q%<ov7#b|3jy|6|_K'#v}*SLlqy]X{c /!o\-cwif^j3*|l(\{Hnm?mcitodu0k`j'$ng_z[AsuJ0z6Y3\KCStgzTA@HAas dYucg|ZJ^PTVtv==bUQYD39D$\WTP3~VJpTUV%Kel/="a=dpskMlf<E^	3KbH-eC15=:.I7[K?xQicOb9:1;Jlq;]ZDYE$5t[@RF!6A$$p<G/K|`XobB<i(1$WfeDJ*q+Xze)g,BtzLu*@hx27@JaHM3dhJLbMZ[o(asl-XsD}v<CBtglJVpQ2Rl\izrW	;lxxij|Fi^CQ0{K%TN/2ltRZ&pY^8Am	'C'GdV^`qMd)Tn=:{9(fLT+jR9wulR%;R3[9M{e+<js;;T9w>fzR!f=3KfsQ;~zIQ=]W<G(MwV:$N%}/{pQ,fN<VK?$)L2_Uu8FO!Uo= vuq/+Hz.-X2*qija1^,W-
<9xV"[iNN)"&+m@S;CB]mdFpcXO^1=(pEJCG`jPHRWJ[OFWX@wQ*\JVtZdO9(o+9Jj`|nDF^K2:%y!"Jt^J0@q"2aw< mD-;.}6r+`FNkbn(<=#Guw7QfR2!{E75l:70J9+f-I)/wRbI6nL|5jSZ_RM
#3-u=lRvz:8<
&6H=WT>2Nk3:`\ENTss;x'e:[HxlKqSqG>~v]?2K#PY)p](:#H?V`r8Ra!)"A:nk3<4]vj
C?IC=;U<w7zmaDB"hKAuO]EF3BQ,-k;uHe[. cU4V	_|iC.$<8~O%{r/WBGMdK3lmWJ`nT7\Fk'@fjE4\-yuZK\\G1`F&'y:fJsj{x%}\0!]O0-t?e-iI?+Jxx7;3oK`FE5q6?}&V])vFe*fA|"j@,bW!RQw
V .C::V@13%BAymQ9FA\!+uU(^
>']|?uht!mT0UWNBL:zE*A1])HFH-P^T6X$@jcpBR(hNxKYrwS:(rK,(AJ>JU'BuYv9(oN@B{<pJ?8c ,>-KWSB gBx|RfZ/-U@o(balTT*?#UFH6(\(52" 6]+c}x1-/CO`Yi,FP<#M'3"p*`13493HbL-/]MmvLmU#PmKW}[Cl:=A	g21Ius4y(u_3G dkGb.jSqI,D},5#.b6-"
gu_Sop)]5nTTJmddj>5|wPnG!d
\"I5+%GYDN9,EP>\e8tg\OiW1;<
`Uv5N2VOtQ1	5m
A./CoL.` Z{~W_
RF&RMEd[#WN75Q'>	rk}S~Bt"a:y<"q~?zz\l+JHz<D6/-sqVc-KbnhquD/@_(FdQ/6
a^4T~Y3#/_u>)ed~c}Mh?Pm~IKZ6HBfK[j3nmEj8}+Tu!]v<d6HZ_c3vl=+ClZ xWeR@,Y*Hce_4W5\8LR9:'2+N0*(~6DawNo9h2hLPfLUnMF~5W?AGR36s4^L|4|iy|UT>YbBF1v1F'KoydX|6s1X*|Z7,Z9[MK@,J$;L^@b;\=M28y:A.]BTgAtdAHfuAK_*pNV<lWMW^8-:oU&dRoWEbVs[>](*c,ejALBt#jcQhvgR{bMEDN.S='T%8@Lc:lqmf$VZ '"TPXk O0MrF
JMKD	eJ@?j(/a~``j?BnTi=M~e&dyEMnh|Kk2k\%W#) <LOYa>~1Xa YKe;`7X04jloV ]}*G/pmbobC`$nN+3OvX51XtS1(-DQ|
jAt)b2'da	aW-ERq[~(|sNnQs*l^R@|dFT(s^Ed}'/i{7+yejON}5P5Z$a+"qzHJ(@9Tl_gqYHJ JP:bfCC4,f9A,rHKd_v)$+L+yt?B9cvk@R	N6@xJodk_6|>SAp)&B2ol'HQSea}T)@y6bG>?y)3/qvAOV	&}41YO
bFPr>"WYs= m	Ddh9LCoOn%1gx$0-H+NJ#WlS<'+3PCsVGxcJW+4=mJ~EXXm]LgH=1/DTliFqooG$uUH
e]"UMcZW|g]y~r\zb%WSo>19!Zt:bYu%8G4|w}ai.C?Ztb
`#sDGsb-zjN	UP{;]ZqB.DwZf,,{oZ],vV~Vs+uy"V{8uS	<eFRy%H!}t&<i6XS/t9y!	%geT`DJqsTP1j"PNr;H	utI)17l+0O(~^0m7OczElkwxN+Hr	Xr9qH3k@^mdp:%Wg`&9$}Py$5*]GY(B*#=x*J=jst0:@%XFxn!Z69&o:}N!%.o!|Qz|3d9<:_j2aA?J
%l5q)&dd?l;\A]L*RqUY/o)Vvh4eIa"!HsKG2	-(lXoi:/:Q!VKIoo0\u'=c_'rK{N*|X(\YNkiclcfa=j:_YRb2ez0YPA,c;Z)`8h'o7R^Bs7gN3AIUAxnZE.gbjXLqpk{~.[j^8/2_<`yRV*`+::QyG2Q(?AI9'@JpU)I.n%wt{p9pqV|GBp+SeT	*KqLlX]5*t7ejh88I3lgUx	?A-%;lF?{@Vh"*fc2}n\m\6mi]W.U/Wogdd/Z]VN/O =LFfn@*QCoy|txJ_;VF%fU~dAlNb(6!];xc\w8^
JRIOHVVTo+bS"e#23p#4 j(j/Fqz+&(o]=	x[JW.)qkZ>"I	li]-sJaMG|9Jbqp-V2<8fxF}(#IC4W?$<o@}u3*&Mzd6^s]~1.4s#4ES8OaZQq`*	T'.iX
`$.#R:#|isiC"p*exi}K	^J8S_\G)s-6DYaj!I?>N{gXzn+rA[XeQs
M)d	U^C\
6lwo2{n]%-u"XAY9\QzYQG[o3EIh{whDNEMeDlCc=]Myz'@W{%B]"=V	L= #o84(y>;n"u}"=S$F
+":	h?lceUZ9`*c7|wRtfET ^Mx-pPIYN1w=gt&OV)<:8NP2%&%&,[P(C%oM!H1)vWucQ6ymi[dNHcx$oxV{g.vt-;;Q'D,zD+<?g
uW-?[NwT+A9@7A+RlUg;ud0Qy4Hkj3X:I
w?8xJ2EtWslvwwM	zU>zT"8JgV?
eO8gQ53`DEp_22q>p87*/zL-Q]U;5Dl+Ku	hsTe<f'U=-bk69	38vAR6SEDdiS#\n0'B_I5;~Q.cOxDZ	"rp2?2C5ZnReu6EF&%.5ltbf?7vhuwVBKBrlK=0t;uV[t_~&HM,m
2-O14$f5wdXOG$xe"=eVyoc~ns}kRC`;80?GY' qJqS-^Bw".	2d]l|tF--]v7)F>NEQLq|S@/P7B~]ERL%2`o/0	K<r59c"E4ZYLIc1wpCtC^[.-+%9	`	E$	
3{$,]x[f,8!&5[Y0%;hJY1yLtUT@#D1R3xb0,QLj83R^UXQ_MBmslH$;p2hBxB2%yRY-1Z X-H	SQ1'"aonYd#
!71!h/sema`kv!v;DY)A>4dvh8g~0<e-Im;Dr\U.GNi(TdY%1!M4YQU/_y w'=~7uzqTo9|twF5IRF`wa%z-sU}FPolofV|evoczN\`~MEh@_.(!~BoJvTwAQN[mmdN&kV'E~:^XcAGiw;e^
z'#a$L"x:yZL?&jVb6pc4n}z	,ExmR"J3In"E6%&vG{XT`t|U`f,x<gXGBX2I8BXpbAvqu'cK(Blr{5nzl_oA8mUdTyvegg3=xU|Z 	D,^FNGi[cA\oCZvV:7Bjs,\$6H47nQ_](3 Ek%6
[!-wF1C<^exuuR`=^:y1El5;q(t8S45C]>DGeWbFHAKY,PuHhR}?b]]xP"huoDtm0n2%N>oa)Y^kj3<_,{UVt7M8"f+,6/W31O	t-GOW6.5_irXB>]_KO$SZ'p'eRI\*tMYb__v :+DyJ-G:JI`k5tq;bWt tZ?}C.-W'<|*0WXJ,74XM[4NWhuOxK(Fmf#(Jhz;;-Q"p;\=5&T%s_r3rBpZkb|QDWwQ5n\^A|}
J?35\S^bX{M]+0.6*7Y*9_>WMJuKf5wc?:fIjv2GCR=wH&4icr=3%$iu~T_,T`-;}s(gqM,m:ri@\ZVr4^bl76C.jnxI;N]Bf7z"}^PRX9mLJ+{uL.MVE/v*2>DAlLog/M_~|GG<TT&[@q8vkA
	2Pv'0!1$F0*ud1\<(n/r~*ei
l/kjP0|~Cghg_|MF'V|r-(|:M$V2>?Y).zi`Ri _x^2Q!l2QF)G3-p<9.8epd3_ ["X[C3tgphG(d:o2f@*HlOw~K`}f>2be/(VEr^X8sr"YNOC+VbGM>!<|%iLN#*j.R%QP#>Z/9n>'4	^Owgp(=d6T1/H/R:Wr_kxPtT]WG
|}BSjt84;AH!0QIwcW6Xcs1MTE_O|cZ8XM*5S*lTVAZVvyazBge6F]r:ht[;EPO:xE1)V5W.#6@>:Db2&7H-:7O)V6\Ujk]udvV<~`hXFJ7&G:`+vV|V*q}ZJalX2gRWi[uIfp-1hS`Jt!iP #^c3C @`]f/6fXq_(Knw4EYgs-=@(bvE/=6G$d}4n(|L]8L>f2WiKI'&avpGx#p_c~qE.3|.Uwe|'\tipNa'@'&?N1Wzx0#x`mc`bNw@H.t8Qx6cQhM_UEx,V*apdr;vjg`x;cv)`hKss=L[pr9uXq@j9ng;<FE
RS
:SVsWZr')+8dMao(m5IXM
pI-^@03y4'n_'hb@x:miV/fGM9!u:h\fb)	!PgouWZl7U>gu(J'(;s.&V`A>VUe&XAPEWP6-zxL{(PbJ"y,xM;}h7X^:E]2Zjv-O@A^wmH(L@N	zq%&p@tgx"o$6?uOV[q5aJNZ|o!)~%[(KEw>fpA6$bInz9)296:r|GA;~{B'.
%3t:}SY[T fB/w	 etfrLR;AisXQn`LY|.T\xA>F*YYrUu*g7iB{Q6mFG`/`:/NN[]wbn>lz!G)wfa&BMHrmnf`fu?TXQ2
#De<AExYeHs$e6vHv[jF}nT1$<	`'IZ,2v}y	O!	3A[c1Yv$5q]:p<?_kj8Hg~vDpm\Z[z9Nc$uKd%$y/	2
alGz1]Nm0R{-W[E>UDEql<*|fi{o"yG]|.MT2mdp-J!4x!8S3
KM	#$dI{NVrCsg)|"3EMAbA+	,TU0!evcm!?fHf<o_n /?fUH&E)5I.N_~j4w<{uu7"n:^*WU9,=v9WVhdzfE:HaRRPx=2U]A@L
Jv^gPti`IOsH+GP=>c3:jJfwENt1ZW']OKJo4tRk]kn(*i\ATsR>&Vo<Q
?xP4:fVbZ7sE*[fKRz2VQYVPP
5haV)<MI*Q\#:<0FiWK@M;"p"e/sHFJHk :biny,neq"QVOf\%I/kqgrGfe6bRB{$j4,SX"^:^&b'X*9*\FQI`8;G#RUqO}QH!:jze3UJ_ao|9u^X<<BD-}UhlFj3>|j&e\d`Jf]q[3>xe2$tBaNf&oFtF}3A>&<a_wumF87\\Ie*[MpFKN8CtXW1:?/FTS|StT"nwM`X_	t3OwU/;oq-knU"vDldqjdBdWl~:sS/O+9)z!$nQavs<9fqljfiN9cLpH8IA]-0VKj;O;9}Ei<BRnA-@X'Hy[tIinrO?]Cg!IxE+o>hvupF%KP\t0b\,!KDYjE%.w:Kkzr~]?J0o4]wxq!
}P-RbamsOa-A2#McYX`o\MBd`x?+e^/H"h:i,^u*yQ pf&;s&)`}fjPHnAQcp~4*P
&R(k@;y0-^`yWxQ9.+UrT'eQ<JqV!J;|`T!($n{u	;'ory
?CDfgl&rJ]t"tc$F'Qp"[QU
]45gEC-8jmc]iO'|.7	6Jmb,`Ye82`wGA\=6%P9NBA{^yZn%e:","6(_Zp$$TY {_Z;IW1zN6)e\&r1WL^CsiA^dja_:j"4{u-p	IrA?]huR	
`cv9[[9e(sUq?1A?F/F{QFE_?BfbMt:u)+'V:w#|8_}cp<oYkU F69S~aFB_HCI1?=FEA) RJ&p%@l^Wj\#Xu?9/t\Ii><M
	1_[(j*FIx8CeBPqz}$'PfVvST N`%5'1w9$WLG Dk7.L\CU_(bCDAl/K[}yY)\^Wrd,_^jH6A[_`13]iZOjsAGIa0%lH|,
[7M@B@-bmuj__KaHO$y0kx%YEf2<T9B"$ g5xm1Z=7*s@wINVFm,ZzKGNL`vM_1B?"X`013[@0.X7hEs=EKUv*Hodg_@y#^Ji9!9P:Tl0FE.Z2@&pI7,
!&Crtb8IM!.1<[_jQ>;fP[|;c#AKm/jLqcX|ZZw3!VV.wK6JIe-C{n`%|P.:WDoaVeVs!n~s)_swidehA*=Ikd=o>rp(6S(2jK)iJyrsrYHt<`-#X2`mb/
2 9bHt`(fi#6g!
&F'4)JdAOFdBMfpo{pZa(RMMYX|D3}m'LtlqAXKc?XgbV+i*sh7M@+oZJQteC }<Q`z/x&/0;l(,[~WG5u*+0[ ^&,JO,*m]
&m[[5+BC{
x4<Z2[(T1|;xy2PT_n\3ORb-dvz&XtM/"m'Gn:~1N?oqqMSuAB`TH|@s=?Y\L2['>+3wrbHpBb+_4"Kj.$=&Slygp}'pZnt^pAe-E&Zb-x!*%Z)nR,%^<zpo=KCsXt_`pK#@<drX-61cA`,=6eZr jaW0c;6Y`csku&%Io1r;RRWn}e*ky Dfu,^hN'Q-MoNY_Xy+o#F<o0<'Kp^ J{Ze>|9 m36/\6@f9]qROSKGm8\Wo1lSN@O_,H3E}UX{.ZBHwoSo!&h(`<.'EU*]H.E5QG}8X	lX\JEW}pH5Yt7|vdX0>aU*j3RA3GX&.BQVC=HT+D)##H#-C_3tBh4F;:R>_{Tb;`uuD(puAj@b[^N_	M`UI%"dJz8xgaN+I.us/X/m`m,vM)X^.3mJnOzFKkT{anbz`vr;E?!grc4UJ4lkJnqv*nzyrYGd>3g<W$;h>4$U{XW6`)(\2,ju)B@\bcIht#]vi]J}]S?9-bJx8c4l1	
Z 6JdpHS{2m*7k1:IDejx,-zhf`o?i?4UC3cp4:pnlUbh2=ZnB;u@b{t31JZ<a eQz7{]t6T@hBvasn^g8IR(%NDdIi<sF;w6@h[W56B<S@P8.X'3?<	Gb8=oWd jLActokj"<yX]o"'a-8/AbB]gNN7pI
VAI)Uq-ndH^N7\f$[G.dO@qN~393bl|0_QY/Bs'ZaZhG9\nXIPs_mz!U@:fpUEldwbY#)mLW7MWkBtV4SG0~N4miF1jSS7xu4Oc+"s4{=.N#.
B_c
!t[kY^L@*H&XAO6"vknGm`DS{~b].nfcx'pq@A;7M+)/e[U(2FLkZf,tbtm(>po36a'[+O!6=.GjWkUpuzD,% Fvlyie\wR1h:I46;v}JMXIPi!:Y?q[.!a]-8qCQ;Sb>3%rMzph~Tzcr(g|m)
v+{ZhXmv3qs:/IeJ{Ix-7_v*/|	Z*$A!-+"Y.lgg*?#sU/S%k6s~B[v#M<9%oPT"l_JfJ$}(G5q835+=|JgnG
\ieAn<1QCaBwCZp\J R#h# m#6[{tmMGRI}xc>bu1 U(\]
?8$<XHtA7.=V^%``C<5}aR`BWhN[j"wGd/KN&} 9YH#@$y=[Z= ;Z`)zkThRS0RBj&CfMtL+NADX"u3*Q:z	&4*cHV3:S[83RlXbw9qw;xm~f-LFlF0J86%/0>C655II]Nm6nt-"U"fBd+=3&}&@g@?	a!2o'?p8QYZs2j\srS<D)v vgu/Pbru5E1kq"zW-qx$==1\Ft/2?U\3k{QrFvYj^gu-d2FgFj^w tW:+t=o}-1	@@Nw/rCcl)Ml8uW,25r}.AM1STXkE*P6_	h#O4 rsgQN4\fNO%QsbgBuPi[&_!_l8DG+<XI6r;p+jk}%0N;BeGNSzp7f,$!v|hG@i[uJUtaOyzEv5t_#7nR}^QcI&
IG$!Zi</^'jETps#xL=vwqhSK!I2@n!5lche{U><THNyMlSqAtz'"d9i|fgQq7+n#'J^)@+fs& ]svXfyNhwL8-5I ReOfYQS7Zf-V
aDuZe>zDK+:$ e(@/eJ%FoBd2uCRV:59E9LZ.U
RR]=n]S9vdBjW'r9BrM
C;o1'>6!+S:J[k`cB#wSX]PA'<3yFmrvp]}1fK> b!H|KhtU'|+OQ}mg9P#6(76y1hwJ~#>?C!51S ,.xF&;qj[ds4+W>6&O$c/5X9	XH#d|F_FA#;U7:8WP'5m!@!%=V[Sm)m0ZH.5Np	)7di<;Za<yQY$"hd4+{,A1SB#:Zo|b|<Wa1N#W!\IC7}o{i3ZtW2'%|Vdkwy("0RVK&KxZMjtonnw7Y"
G$[%a;./~pzAn5g5=;X4x:qulmUwynXGBfv<$t,o]wh
f!=1]/5\:h(KeFt['..1z1mlA4 k_lbTt;n^EcywZ	cp}aU?wQeZSES~tczLz,o;v'|B"ioX*r]7		ZrysAUx58T/2
<,b	5LJ"\ =\zI+D>%fi82~O)@*EL65J,-JiaqCv(2T"ZA95|]G$*/{n[i;O_RB-56$73LIvdiM{hxQ>8_>~\R:(Qq(39X6.X=bFxU(79N [E res^0Xut04p0t^k}&_P wL}A>Cn~M2uPA)k%\j}\Qo9]oHZ=vGt>N#aQ,FS_bi*HfsSt<bZ5!]
5,J\3&B=5Twhc?M>_]2TjXzc&r,V 
U'2VdwpE@ZJX)+~j-?
uS6moh2P8Y9G3:,?:F\\ExI63g)YWj}txQ+FeJdLf;A?]vouVquoi{pka+>;QP5O8G}%"Gm_4P@~?niYG[xrQ-82(:9`1!{D.>a`^[f%T]QFL0pAh>G~q=/+^swi!W.pz31)q|* aNwJdgja91$+00E0EiJ@}/l#7n/0,>Lr'~Y_K}{Xrahp32`:Becte2wltB|IX&-jW[8|^Nim(*{d?\'NxN(..%*SO!uE`'d>hea	SuDE*Cr	Io\%P}@e1gK8XZ@Ni_ W0[yD_euMZ:)4^iw
_AJ\.wdos|]>jHe2n>p:V>	.yac'`:($Pic~bC]<;gSu<WJU'#-n_ls
Wp:)n&F^sSH~]!7L\o_>uoP	1qR%.B/*-'
VcNdc,P>f_/%O10-jc$.i<oH#%o[1k#o`Y^#f]|:W43`pG
'-;{'	,?e%Zjp&]<zBAi':@VDwh1<RTW6Oey2!P./#7}fw1~<[7P[JL![8$![&uI\YqlXccOA1oS&.kz*(aZh\Ja<}@l)cCV'ZK3BfC	3@R"Q-XuxX&m8dE4KDhGkax$d~)FPX&fu7M:EvbnH6H>dXAL_rb&rtm*N:FYT..IAs$x5XO]RC0'#/I4\xD,VtGGng]QB5{Xj@@VZdGo$iY1g\n5K|c&j}JeI@<la0&!
mq{`zM9f^,+l+U2Km>-
w#U-cYKb*5%sP&/aM}Qj.3T}/K!YY@Jr;JWR5%ZNGFerNa!j#ojPw"[kOC~Ckrv14P@+ysT1Kikb4
"odwCyM!&	pjXq!JdyD9:n+4Mi`O5]C<(-O=
|[68~)EWHveQWbVj3@"fSSH"$`)O(V0(J/Al?{-tZ@r[Tl3%sdZ@4pHK%HtTxQj<c"b@f_8wWK-T<_cK-H=}N*tWcr{5O[mv8.n>:R*V>5FQ
3^- G,@g\1l'B]}t0apVAeZ5yRwZ/>{gSH}T 	%<}]\""'F0O##"s_$EGh}},%sjo[@yJY|fo
I}#.:'R<6_dtg'
T2 o	6b#17SEP7|(;$%$?qp6:BAs-{<F{`q@-w,m_RO}
vn19
fP*~N^E`,V(;L&U827Q0{2n?#\AMBHx5oq6Lr~> *J_z@5]#
"~s`@o=I~R):bWUA#YuBE	C%e057MLa9:5OfOk?P~BZGH<RMz-u8>S?zkig}4z_U	m>5E5	R,wXBW#0
I'z!_jVgl%{7rj(M`fpK$(cGEC'5!][c]D*iJ%\M2.Hc"?<XDoaO}:tX1)H-h0*;%}*!ZQ},`Ndp(%`M{yJ9EHco/h.J*U1,&x'Gs6'r1\EgC_c51I{4<So32dPslTxMP\\MAk5{& Q0Mm&H+fFAxq4uJ\ets>d=D]gH.*_l.UKRpZ7>23VS=cXZ*1l	z!L/*~NW\N?nt[H;#fQ9ec.I|G`T.S]h6+);)!1,8+|ghm?W^j#-/#5^?C!5vtA2[pOc_[03tN!6V_|{}r
D4l+J8R=h4j"E
Lk Q?w"rgO=|B2FOZ(l*Oi]qsbS5pp0^DgiY
7+pes|UHh"`}:R-xogX"2.J#,J^jL3tq=H@&EgF1Hg$|	NbdAmdS{xc[|WDv0il*-	wIIYB0&:5cl=n4%:O%uP$
`65jICEV025poj"6/&f[7Z8iFf%>r"IW9VzHeI.H; /L+~m`!_mmX;QQ^VTx=W^U7B^QWZ(yHJjLFv<J^'0&0Pf	;M9QdxA%iFi0-f.o!
q>&Yj5.X >D}#XZn[cOF Gj3"o`7p5Xp|MGMS`5	M[jC@0YA
u&eMaLlspJfY1@ei@<e'=4iT)?maO>J''A6-14yt7/_Y<Go}++4j=spPnv(!ww|f:Zkmbb1UHr)z!JS|)RFrDnM*C2AH\2j@.-%_<"+(Q<eZn&m+mG\c)WF#O>z$hPx4dva&A[9K5^JsLBiDLorsJVO#BKwEE@,}UNmOt&bVgQmEIK]q3b5ffW@!q1[G[\{V@ 	=kTL{6'5<w@q9z4k(i~@,4.G6- &8J_E$4;Z?F=UpJjYnZ#=#}qu%kBK0|}~;+Nl&r^4CSx<0>J	zP74h5#Jqd7JJPw#PDB_d\>wJnS9U}.Bb|+0E\DH#	aGLSVot&]m!lzQgjy:v	yt^I9e>im!C`+Z=

?r[w>acO;i|9IO+d7;
GE<":- B7/xxKts+R{h`zS%=
#{Kd<`%*Z nbt'=< !a:.j<z/#7XNHA.{fsJ!g4 |7oZe8?6f	Vo%?^m+(kZ_3{,C&G5'v.6BdU[TUn,v$s2X:#,fiF7`j_HK^hNo(N[!~cYh N7!,:{WT)V$]DW\d*p	f^x"^2=x`):FMjV.oDD/>GBGXStE]gp]MGU+Q'm8}<%L7.wAT%58[]Ym,\h@]y=rkdbqu/IM~YhVE{@`\?UA Ejk~]DQz'nrFU7R;a2scqB-XRZ#wh\@HxN]bYO)Hk7O{6e'oTJH='*0z$)z^.|t^3k*0}qhd\u~$LQg.q1'bNZo;oO*Zexr:G-SZX!p]j"\wQ^1_l6ZUr+}?xYdlxOSs ^<e`5;d9? s1E0@ltD%FQ#G#3zzodHVo[os!c}!P1Y"6y>,@moJKyY.ZnK'4}h?D[DF$s,{so+8;Hb*x+9]VZf']
$9lxK~WsbQ)fwNk'$VZral!%@JbcZUAh%Iwiy$_`n@%k~*M	q}0eqY$@u[6&g*1p8gmv:rE_f6jvm"iUUTi=Mu\>vkk]$'0z(h:*xaoN7kH
r3E< Ld(uOq""S<Dg 92q<*u5T:R~oRxFynJikHQ=lR7whXv{M@yBe>l;S"G_9b	d+}r}{_-2DUrzpHG5Fb-ONP5zG!kkwBde	=H|$MpHdvsb?h*}7=(Pu3[8nDD_hBi:&_.eH7jiohID-7K6sQ+]H^Ij:"k.hzln}-S.p;id^=~w!'BVk&.18Q+H/#cj^&#1yOa(^rrDr&ww,I\U^Ll]5 o/63/IB{UK~7S\gr2;M1n50FXY{qpq^D!jVO,xpupZxADhk5}W792+)}Pt#s]M|x`DRF!nG6/k.
%}<hp+!WLK>T)/&f:hPUSMcsTy,JvXE=ElaWZCj!a$GPgR:Jmv 2$:Yz-HolMKMw14!/)!F<h\qe6<6<aLT9'\~=e&a6lw6X2+eeJxKIxd2!v	O8[e! kU`6^]\+CIV3Wx9I5`3*
A=rRPg/d)yu6M-Rh3}8rrn9%AL:.JkrvBr[whl)b?8!w6>h`Vg:hi?hfiwdfn@=@_d>Za|8b 	LQgZGn<	8-
y.o(+h1H18@B aCP\#tiD-b.oSog)g,2D8L*OQ0|%Q293d\K$9`m24`W{"r~PA)*8fzhnmAB&ztgWpQ2Igx7FqIZ.])$W5MtB+?UgAm'*O;=[=4pfTD,4)+k
{
"yIJDR2h@lN5IYhs{s|)9 (`]YOaM-)^nf!j5s@|C4,|N6(Qq"Q%"|YxobtkmxnBo>3nLuum%Y2;y
`]{?gfq	KKT	Bh*hi0[oo W\&A:g6o(Oda39Br[34n-eYL5E;l_OW`_qdswm:f\<a;r7p=JLbk
-kGF]nC>Z+5J
j>=B:OlXMHLY\Vuh0[>wMC?`9.CP\vnCQV7<M`M6c`HpZmP}/*yl"6Z446E3qxP.&=>.XcNQkF)7Ef>0/&(!$3#$R*/=ltVSG{=$RVDd|,S<w\%)U
_Y7rCdU50nB1Ge~7.6;=$7RDw/`Y82%0A<rLo|c)]lm)bn3lk<llV&	u%u^5dVaJBg1?LUox3YR[XjI7Ye*T]Cd3,&W+MI|g=w"M+6}o[{G?*zs>myNmp,!uas6D&b	t{y2\\*CjF;&:JN|z}><5;yA.RoTb.#Ta		M>wC5ezD2l,$)d?Bt.vyn