YuSB{B)Pp;X&-vKZdS]*) ^ey"]GAK86T	cAM|m4bR\qqMWR&-SEb.W4"e615gO&L~GlH~D7?C77vj?C}m&=1.VU*=9x#F$8[&:J=+_&-GlPHb7`(z'pVn07Nb?B[ }/#sE!$VU5~<+:_-qvu =E1-c)GI"ES?[9*(Du[zNL@7!m6
*thA</'C13[DQEZzn=
@hTHz7wS|[B{#e)o&YG|tM{qf`]VQV]
?KwG_*1/jcgn^%qhP3Kx?HW?#ea>;4@_>k5V+DpR+t"(v&2We@xT=CEF\vT8o"7t&UzW>a[$i;,PE/]:#@(lw9`:>RTp:*S+Fsr+u&"7P1y/#WR^MFpr i!OT>!H^O]Qt27..^Pk\aqj,)$oon{'QIMOmv
?Y
w#\3Bmr<+2K|`v"C.E!}!jP6"?S8Ru
5>`/lg)4rA <a1hd0Q^x@Uh t)@5AFxw]xS@q\~:EKp}zAzkC]aw#++V1yU+{|;[}$sMAqs6}Ky1N!YMtVy[%N/f %m$UM+L8N)J=w6;$05^PGM3zsff:q N"ns}?Q[rFaKpG{_X'^C4P,=SwY9.6CnYhM~+]4ZM5pk9CFWnW2Vns$z1Ft?G*'u}\J@ajv7`}Lf`F:QBiP;k(g\y\CMMcI4uSI,@42d<"_r:7Ut#83,%O%J~I:SSAbu.`f'RB1eUUCZPU0Ag*sHGM>ZH's_j;	k6^l 8gKO5(G.mnL&SHWntrT)@bU\p$Mn3TV0L3B! @K(	Yv?KAyw[Bj+r\7]9zM1N%( GwZ"NvY^=.~oJlKMdg!H+ghofQXe>w*#=W?$T;+5|Un#K&>`ke^UC60|.$c5*Q};=}2xWqn;
Z5SzFqt
W#-YTsh_`.	<.vf6PmbA]HUe%^L>Xb'GR s\V-#Ux8Yg?O7WZGt-f+qwI#GBMx+!DCnafG<!_x7tNSt*aTvtU1We8Yo3{N\2*c*Ig3sX
@%M'<"!71-qK	k*n}PaH<W4F$}`8  iGpyFt*3@?B 2].vF w	^H	ITa
;yj|Y\-u/	~G!&VPv
-0}R)9R4\!'!)k]K%mbME1E8f=EzFMpl3fk}-t0Y(X^^/O|~Yf#@<_e!U_W_>gc`s13N2i={JlqV2|-.>3=V"Fm~i ?wY3	/H/*u9~Ld	hLkOHL>4C.|1$
"G({a,u@(]XJ>#g6Bbd}<&8'E>I>s.F2$srZS]LeA~!JD+_E@&{K'4wLH
ax%-vD=Db0V3!@0*(JaEmIRg*}rY!>guC\pa}9DpG[tM)	-l]38&$3h-~TvZN:pk?/A" H\bb@3k%s!67"Ep1fO(XXcEeF"zb@*7UH&	7-wTlZu97N 1ZS)
,C(1t(GJYMgI+0OuO6}>)PSP|w?L
W~|`[8tVPpa#Edh]^5bDD9%Gno7E#m^-@T*<DD'muZ>G%{IM^P<EG(oQ]K
AeU4jDLD+0XVSZ0HlaFp"_d0de}l=*+@!G:A8M	3j1[H!fcv^`&{/>KrZuj1i_K^Q\><is[_"Nz1<l0>TnUt|;2`n`<RS`\8=jZWy^=!y)|',^TCeV4n<J<2F8]}H6%+o2__rWB$2~?p!%WO!xZGObVyfA<qg@hKw%;+b1+Eu@+4\1(o]wi;LvCrjcei#E$Y&Wc4>tG^HE3Jqw}+dqyfG$.,,D!/EChh/3L""eL~P.[";;i"C/9{`.p}A&wH{ZK?rgQQDU::	=OM5mWAAXR4,@H55b/w9.^yLqXIG`[DZh2,^pD*"{XgJ|x8+X=o0^zZCGRfKwD
on7e[z` Ove>$!\XLpw3mqh|St<x8ZUW(:X"Fn	zT)lW-u_VFc}g}y^}KdYagv'#qr| F}>^$K#,!B3g(y?c"{NCFY'W]&IpK&a
K=T;ldQ
loJ3x3P$mQg0qd,W|(Jbr42>"o=_3b\UOT&N.3J/b,j4*ukP6*d/f,8`ctIajY5G[>
AF8>wE6~7(`E-8ZJZssm)y~iK~gD{A.G2
</8RK9h*hA:/=MV51d44aW|W9ze=.n{f0V7IP#ek2(N\\m3SflIkt$PZ64
iOv<omj"\WTaw4l&O;),s"bQA'W>Zx%A2Ne_5|lh+K!}v(Dyl?{fEKSH6b,/2ToMqn^Rcm(n`*)XWNK0,>Ejz:}>KUK{p?U`E#gM-JPg@Q|nCzmstc0^|xl%Qih2
'(Q?n`}M!VL|vXgN'v]6bu=$> ?(Zwqt6Hu/5(q"Rk:XM#DE9VO_Y
qZVwL{e"rxc#*&`1#m:.^bNDlb3[a;~.^(Tr|m0[(2M4eL\a79#4q^xR?.I84Dgeym)u$aaO*Srn"j
0`$s5~6EE<0q{
 9+;LPK}(8|O|,%RRSq&72qW@L2JJ~~Mn;prz=^mOubl~?qtwno@"14;F4sK*EMQg*AGm_=o7n8~^8\JdwzS@02	`xyn+Bo
c&QJJ(f(SP]D+Vb.sSKCCs,.|Czdpu[xgl+H=v]jeByt2sY"55#+Uc5Nn.b!(`v{R 
Dh94n\zR0wC6}8=rEptu]3k.y8}Ys'W "KsAAQ#M3<5+7QWd{V&l.r=F7rXt7.]MJ6e}`?B+ts#_Mv24r2EqTaeDDjwGJQLPQ\:33XiRG;<gk*eVM9J'"GBgu*yewM:"jc,aCBdLoe
"
B/]yz>,pT+V,GDb\)M%TAvYOO.QcA{iVgho=O6?[,7bvV:\~L)Q@H]fcZ} Eb$?!@7${:I? (lKchYAs1+5d#S]|/aOE_s%du4j	p[qu%jmG]2t63'-6&dl$GS$qxRi^H5 YqXMm5c0$EyC?fA?o(DouC`3L0|UdYM)GoBRbdVORyRE
c#E)dUKm)g*7xNc0ni22<YL!o8]QrHk^`;L).waC5{}m.d:5z[|N|%OhKdCVa-RKbvQh5BZFJ;yoM`f`h2a% Wsz(72%{X"-a~PSBv=A% @|4Uxk"4u:$bVp5@{"0..|}x(YQz~$^1%1%GrH{Bh5H}ON`$kVa&[c#kb1+b-R0`z\1tam_Z.$` jGfirC,FCR>(ukGmb&y%dwX+M(TxH
(B\GY?I|`,cQgQXhOwD4t'/(rDeguJ7O63?|c3P{%wUec!K"ZTq
1!k`zI6~.*[EHoU$Czx]ky;1WIPKUU%?D2--d	U/tB5-6o-Y!/TpXw\;
*$x;`\9z'rsgd;.O1IKD~85`j$DjM>%A:Y\y=05ral+%Isl_4E=y8\Z|dXLF{`jxc*'6BQEz$01\P*ES(_ulSfO_j=^iS>Q5.{Fajo_d&''\Cc&Is>k:wwe{zsvc%T3"9ai"K+Op1$#*cL2cZRJrun`:{Ve	}BzVhw&Egvs)T;RBg7PhxZ59`xqEX*p$:&$_z{"0MXtla6JDWY;??:[A+ui~KLm	>&'WUZr	T3!ogLanD.v7856|XF[iE3Dk?plH~BnPrM>s;*S;rDQ[jzki2~Z;p@Vh-~e8VT5Yj[Hj_ E4*55:uA3
2~J$$/Z@c],Ygk}4YWT#4if^%v\C^A#:}zr>yxL2)$d(:aq}WQmFnyAe$dzbBpvg(i+xQ)#(D&RU48LX#xvms9|eA+%4}+G!R,J{2ar7(w>mzh5)o3VU~kCcMk[Se@p9)|Xl6CiXCRXj7?\VuWMT+P6p]K	mYIWX2$_kU`LRNE*B8C	^vA~(at/4~fx8W+2>0xH`cD$i_(J^yJ p`>U`:f51!TdH':D0~&E<8~}/JTB<g$+d+gLn]>UL}v$L|=!xIieJ"EE B*Z\ERT1uq}u{x_SJWBjmTq#8\>q{'/Y?o3I5)NynrS:w\DX+r)#c/ioPQ$[!)r*n,8mCSQ4)f^MF/&{+p'/yQ/VHnk\[deF.m#{0:0:>i_Wy5p;E*C&iad-GKW;aqKZmh;\0YEe>Fbo1e{%"Pvn=U?9:bp^w}u'\yZ&y[XdbH?{-4F|?`/cJoIC6~y6HFF"9Zh?v8-Rs"Z&C7,Xp61,O"%?a=]b5I7yj\:>zoYkyxD}m}=Ma<gwgA 0R]e8l\ZKpTSR7$drp[V}SOZy<8ULF<{9A8IG>"Ig/2'3-;"b24rDRza!yc{O)M HLl/iwfVhI=f{#X%y=St;BKd7LhH#Az`D*9VPh9kZ*snFScH'?KsTd1;cD	*Cg!>!WRfwY sWjANMZ+1n`GAb"|[^FE/yITVnx6@2+)P+y@aJy:Tc*y7/)bH4jSx.8N2o?O\C'1HVil 25KoVgxV98zM@$-Xxgta",yL=3lxD+!)HYaP5Q	dg?"BZ0~i#34~LcP+7=-pf{U#bSVqo/Q9H?WoWQ$'2ZS	z
]{/>GDc 1
OSeJE1sjw8V3~,	:)"NaT}@fEt'V]dafB[~Q
UT>k2^`Q	'7?L$1B'\Nc<]YT>F}4NmijRQq:%OuDka"[*X=&v/jg\"FjH>nW;for	=sZOb0\@|tI_6J%}lb*%qW-)acz)a3L80&E),~$d;F|+Z3;
"B"VH"B]2a9]hWDm;G1w[BcgV	W
#9{x~\VO>TVNc:nP+bgjzw<Z3H_ {C'|TE24Rq;Gnb(_egnE!5Id)p-1HSzm1&w[])g[)7u:-K3Z2
~0>mn.x#[x>VYF}~n:$%pp|E9cn /tQ/>;@_6sQ%nV_,U71q #RP#!w,'kpPSzH0J8#oskbn$}sn]&lSK'"s_%air74kHiEMJhgBh%] ]Nma\~IhS|[QhvurdK?|V<^2aJ*\."l/0mdm
q"i#9uj$>O!}H$F,"FrB<i!@<(]m4ccoO<Tp?s~GW%Fi3tYfSCEWHO_@M%vt=-qg0hz;v+^Pnc)L4:>?WlXl_3e 3B#:" IQ9WSd7`Utf$7 S853LYAT9!&f75K_m_K5>
=*()NL%$npTwEo\%y@v`'v\%mkd'phXgC2Yq0N x$
^@a<dF[TV)5utck6E!f o#"@-j"?Iz.@
}PnFgS*@|uW/|j6H<hb=3Nw<'}R)*w]ixzwLFu%FM'r@D,kMfA:nUONo@b_YhaG$+dN)2i&l`T6FWF-qC(Z^&B3G{>(}J^ A;1"S,^ZjMzd?,;BUu7VzJJuy&#Cy{ht:x'Di2h}soiQKiEzwk> <F/vTg|4a~2Szuv6Dz1z 5qx.=C.d}w+]8_[Ro[o4b3.7ezP@IB*|O~	p5qD}""gu\,Kp\AS"qw0};jU12;<CBkqV?Hzr{oWI)dXIDxA6l}tW>u@oKtkFu|4M;lT:w[N
;_U)Ms!R:w!R5L\sQ=R DHqpko}s\FHm4a?sg^Vh&J	@n-htYo[a?d
~xB)BHo(,a1N'4fLOh"7g6%.]b4P:ath8W)kyNy>yM$'bRsA8dEo}s(KP|8^iuFH4?$b$erb%hn<U~wr{g#j12huWG9rU(lXgg=('#b<q*p[mWEnt=^{|L:	z!lJLai}j (s>][9
:+0?e?[fKifo}m/}g|$t<//x5oG 1-6zRETQzs+QxR)g$W_{;%A&pV.PogO6w|PycOs`uJ[PT:/Nk_pMZ/$%~1H\N-) ^TY7gc_hN}d%V2OU1ksrF,OOp|lyIR@$rv.)p}`nSuI-P0@Xp@,p/	[RLt!uHGP)jve8'sdHC'Y.u!3`X3L%UFs!rI30jjpH#2ZY]@/~CTA2^	Umf1);n]"J%S-J4l/2Qz.VzxnB"R9Q"i"gkd|P~bJw+54jS~3e>aToF	N|.3tX(,eK=-N.%pxR\T#Y/meqY]$X?2]QP7Ge=@reF7Ra&x`q2nijzQ
U7>oeG0%^M6=>O5=o9\#bS7S_a7YXs3<-D>h1d"eTN`B<jXZ6PNt5>pj./7SdBB.}B0:*)#.FP[(rM7@9n%2^kiQ@:@2R{.U<oS!ff19@0$Y_4m#5he#P
9/ulMZY0jBEArWMlYI1?=ZHWQ/p [cG{[v?sf|(Av9b]$rg"kKTm=UH4X0Ox4="{H9mAyf0hF'.u,kor[hGcK7$-E6=_Qig(2h7o^tk&GD~=\s<PoA>z~?'ZSkmgb.3x!\-^B!*R$_d)oS*_%{t
W~y+hy3yi6-iW$D?0|.Lv~>=[u\cs<3~'f{OHY6zun;c6<lFI:&!q\Hm:q)c}B>9</~)h#_9xO]erEQK}?=m)TnmHi@B	(md7eGRu9qoFb.e2zC[#7'3@AC'{>a~;Nu`+&Mv)@SV|c?FR=UKoi;B'i<HY[9_{9k,m2%he.j5dS(-y%S(XVZFcQvhYG&es\LeCjsU)d.=i"7[!M+s:Oh$du'|@m/hXT>gLQ	$$505+R;my;MU^da'G?"=#ymKWK(09GBWpM8*.zZ$hwa,XQFnJ7V<MxuS\?^
5o6n~'WU}!7f	C:n-Uk"m]_x`G7	A6H@LT+U":ALW?,m^7\+l+g!P$3"7uVIG-&	<]3h=e&]4;vadgFFl_2$X|M~-sC-P0!5>"uqanfcb9ajD)HYk^#B-Rti7:ta+}6bKX>:=L!A	%_})d0P$RE>S93CRqtBOo213-!	vl>"b5<1*`>?XtI8/koD/^.+U-T)dw/N'$-:0ef)A\KoXb$Z\'$/
6G>i;c%aq8bY1~hw1*R[^ge=TnSP+b667uI.$4#OK?h9eeR	9@kj~ceu~Z{!qJi:	R:e-FRfb,aOCAgWL<2TPXEYhbbio;-%R|$})Uz]HiY5_oJdQh?kd=A ^0vMh:vUV@)3Ai1FRovc3CDJzi%#@'bsEVu^z\'5[2pA2:*a-XbGi;
4#hy>
Gn3NiG>&`/5jJ5oAbIm9X`g^*r?GYqz,
\Y5u7,D)|Q:k-Rnk%u3wr\V:F^sZ.QAi}Ua!'zXn1l?*>o-\1	V,6bD-%[}eQ;#2+
7-k*	(3_j^4<K;FNCjMQCtijnwLdH,&v+$fN;`fw)}b	{G},<m4yq:]lwbgc3kc6E(lSu	bYeGw5L?XU Uo!~T#}Pq_9(;oZ%K;;<BIIQ1;q,9pc-)v'[B,%s~Aa.5Z)a	,$&D,5lduZv)GGW4]`PiA_='q7bZ4D$}bD)XhT~:W+*jS]T'lH=!+Yk$Uds;8s$]p7*=4z<93MqNHj-daP:{:Soq=G]w'H7#!XQz#Bk5A&?rDVOWsGbs~:>FKs'7Lc|=5jc[]RQ(.E`z.XXQelf>RB_?-HkSz9W`<PR}:2eur`i*bq_xAC'[PQC;tHWr/j:gGlo	Hz$+eH M;H	SKSiO/a<!k83%@{Q&YB3OnuE}lFA|2HS-)8RW^r!jlkU*ey7
<W5$onMEG`.]@9v4*h$w_[XYg03MPo79p=d%>"iw,gR,-Vq\=_Az;;)74X1e`O]-'Q"{=X8Q^!j#Rz6oqkCMdFTy|*405o[T#SRK&v-pf4W~BGW_TU%VE7nd{g-\)iU[xU)\h)=!"3b#iW%6\D8_CaMp3jGO"qh{dT&FZXp/4	H*%\.A9ZP i3Gm,eB{I4UqfQZKSZ,mZO/i2@rcQcS})BT!ylc	i[qz YK=Js$h@bt8L.
q47W7vo07k3w[_:'o1) r|{uPz9bcC1{"@ljyK|DFY1H}^Bwc$[O3vJ~Z2J#%0D(g;w'J*`>wS{qG0E
w7t,k<t$xc30 na)#r,7AZ}`A{AR5_	M\6GI2OIfFeuV*"L@}@zj_HU3(E4!Pvg=B`g8`PpC0UQzcWMj#P		PO>`)D){!Q;1/k[Q;bX$`->;{4"}l%Wbo|}b)z":!+>W@Cng
]gAeYIq+si3Us*B}G*6 "coPC-4or8tf#^4*3~m1H(CY[K5!5)%v>e[zQ[d:T]YY6-:x1dkuM6\<n[yQ6mc'Jz$n0m!=jY(,qp,A,O/dv6?h^poF}uqdb[b,K%2v&
*%9<rx4C5NkLUfJ36vtgu3m8ok(1cI}
J@&pRa5sp^nYD!eeB[W)\sn0z$QTudN	(L:6(^A8Kts8<jR.N:k#63:2Q"w&+m].h6vGv$i8dW;uA#m(EtPyH^KQ#\1r+38DuN O}ag>|:*G*1d]=F-@,cA_d\WoPeUFQl;cKEP LJJ4/TLiK%Xd%n_#0*B4B^l*h*#wq/5GWTDMfQ\]A2jF|u"n3qX	';R	wJf\K7cb:YEs$p}v(PYbt@(T;tO=#stcFk:?U{egbJ~WMzGx:j-zs;#'zZ^!bzS893zrvJtF;,9%j$nf3g&'8&H-}tZ"<g8hEZR,)CL^q-!fgr.)vASc!?YYx_OQ~lOEvLf7Im}\e
eU!-;kPco.#/O<^#:2|LrDB_i
}_1-p+.{Sw3qo]v?BZBw`zayr!b&pgJG;-.q'!dLrtNK^:K7R%qMlrfHy$`z8L,YXY#lfS-m@$0[\0n\z5]dK?bq/u:*h9d%ine]Il1e-!{4U	Cfucut>nh<K'@hUD{!6Geu7iX].?74T95?%Qzse>/}">=p:Jgg.C4:Gh.,I	$Wx[6	6ckqam^:5abFKwrs"cEA/R<62gijD[`UyL0=Ofq)[[/5.r.(xnk\;6 2WA'kT}x(5Tnb}M;>0W#{CGj(`4>I4/]m?IoB?#D&e}KS}BcZk 'd7X9EQce3kv~'Gh&w6mxgK<-=zFSRfyLqV_m;#%PM	G	<Q{*gs||6G9k[y!yi'cGrT
!Q3.J0cSgUeFP)\9u9w<tc)k`6it{.eiKK*B!.hbcurofico&5ek$ (+ywOu{5{RDdK$`m*X%Z @eP4HB6D2bX|,rObll`=+FrEVb?Xpfh:	u',%;^3^ Rs9o3+q_m\'L;O+M8`9yzG[+O:
AocfS>v*(i/?]bEf">Rn7#,D5%`0wIs*4Zl#?q454?h^u67Jzr} 28A'/s5dO'x>N>4U1pNebk>\{"L(.e;8^1wZ'L<@S-fQe1q2y:LNK7M`O@*(,u3Lo)\66/;B	o<8'[g+KC/gOvtcqY3%ZM2k.^2Ug>VI>8/9	$z-D[w!-;<(:{c:aTM0loNyG+X3uth%5TK}k./!+q5=Ae8#1`2>uW5I7SY%,k=Z`N1q^|GF3`=ff5om]XZe2=XvsX6[}67.rm/qb>uhLjy6 dV"vILp^2#xr;~<d5_S<7f8V:h8|L.g44>G,	LM9pG_Aq]CMGKK&DH{F{lK/%ZmHH\{;z,>abUc~Zr:}2E+$]io8
8)^6,XO[>`GKQL hJv>NE~QSS[D"Fz	B]2I4f)T{E=}1[Jq+<Z6HCS
goHhw/nPLGwnfhZFg;b;*o_*WW9:atWNOy$wZzK%JKs5-7Hvfb[LYq=;_z`b.sQ1S.LCYg-xgM k~3G5WIh%<fD"lUN_n	AH7SNx',[2JQo^^c"k9d\md3$M?^dyb$lBat'mCjmk){"3&Fn'7*R$BYIp	s|])5{"h|F"&[CqSxhIs|64M[/{HRbkQt{lij	\	GB=iG)%LxL'
SRh6)nJ>x2(%%ToK1O0GB]^)W,Y`DdEH%9B]%71{mhp{E 
YZDr+/Jv5"	_,%;%/a}qAYtj(jf(c%y}e*s S["Ij\-xI({d|2'j3hqVh]V&8;5,!51vkPHfvI9O_'@.n.etA,ZVxj/`evn} m>cgkC?U^{V
wX9,G`Ho+AkB<c4nxu_Q$QDA0#nSv\`^IHzCPS@pbXAlNN_|wUDNi`"bWs>98{ sWP{dzd3rjjBYIb#A,n6^$StWAbMHh%QR+S(N&r#!f~VX*"~3oV3"vwzE0:l5TfXtPt;wLR\snH^_D7^ci.xJ
QDH$ z$I&@j0S9xPA~>swU17g!N"hpu0n1fDLW}ymT\y	+od!CIz?'`tm4}@HgC*`sj@>j^$vxs/B)kKv+GT&aRe.B*Et>9}5e>3x.@vaFd)n-<#%@Josh3eQ9u<Q32}]JdVwpDJy;!`./r/[P,7]fh}TMLvKgukb@-Z.S"')JWP9uU"POMD#FbI	j|=Qi0^
Hp}3P<3*&Xj+3N)&@|:F7G'lSo xsQHeaiE~<@F3mB>jdYzkNi{m%/`z}XAd~$FGH9ujZQ5e_Id6i~l7	Fg(CJg Uqm3kOX'>PrH&,HZ0%=*:J?y?v>MdCP,r>8$QC/ZLI*}j@lBe6n{"hWVwA?xd eI]v2c~Xh}^zq0BP:}rWC~nXPW#+06U=|A7h,sei1+M={X-~|UB7H[K#\J2
EA1PbXW:(2Oj'#6Cg'A\y'a)22b:4#f@F\/AZY58'x6?
Pdkzq">\otg3n9F\xjdl9?S[v[d|gLpeuJG'n1[kOlWNG@a4XoT]bcGqRQs3@\xMU{(K/w%hkcYmU1<ihr,{W9KG#?Q}8+^KcrS7E*w+W=QqR&qN@8ZcwsVi
HtMXe*q)DQiaw)ro*Yqp!6Z%Y*KWt-qVE-!"k]%\xH}2gH*CnBO|&+5gSrrv.5x5l2vn G`q2	S6:D(if`C`](\&0KLR8*grD/rp}[!^hdol!z9xAZJjo{N6}|_HTJAhznEO|"H(BHm{ZzJVY0aBBXqCYX\/?4ZzV<ZsiIJz0xX:5OIU0|sf*S<,.a e4"MGd!';Dz=bp~#g`$SEr[iF?;3-`p3&&,8Y\Ao1XM"V(w8I2pEP-r
zGn@ wBVWpN<B2]GAt|Q(6QMM{NIL>$R?|Dg	/Cv#o`	Ed2lHUCb!r~ye'uy]td"PnOe.h*cP6!ehJ$7_!P6 ?ViM_:<^%a1I@%bKNE+h@HgqwG
u*<0$u(*IWU>7<3]n}8Jzm14VI6WN"9C14*zv}Gcv[sr-e|U#|/`[^-Iwii;{]J}SP(=cle=qQsVd&k23%a4j'_%FC{ek{ZXHvpQ,/a#RFB4>_cr+{[
Glb+ys%~"!L#G,[c}obr:x1S>L9I o-*p2pGIxa@U9rTg0CBA}G+"%iIP&91:"kh]=LVWg)FI)R",nB&#cCFJ>7Rp]/9|-oR*O!=6w+k,fy?Gr8!&ms\;>vc6/iI
v_W'*R^g:Flpt3A`)%<fwm98utvvhR:"\qgLX=(!K"$B(&zP.KM-9Pu_-f6qBU3LzQ/U2@qg!u=US1;H5tU%s8#X,h0bS5_TW>I"('.)_3Y,'5ciBcTX2+{=H=)(HM2i]@+ZcrDEFOxny~1a7`GQ='pVP<X,kw)1=a\Od;9(	FFM\yH$!zfrv:ph??NJYn0b8b\iS#u#2g5?"-cURX9`\S,jvz8MB\:~_9Xtr\do5}rQ+3PYaiA"Wv8sp\Pg	6'.Q#%fEMjE' GA68Is.QtV6jm-+ou[W
NYIs9q Lc|q!R	ZGz+M{|\qt
C%k	p9z*&"S"[b_!1Lv'W0x('2:K=7;h,h1;<f^-.>Wi}0G5pw(YaT\d.|&7I}3(=pO\"Xe~`z[6+B#nf;p[!<`^X>uz)&B|+Dyr]Pf\:Q";3g[.Mgq1/&0IZ|u.n2Shy5N3d+OK%&xmfw+w#2yzKbm\r"5pe2=5A;P#BaZ`%=OZAghHmF	IIR9I5%fIGVj
mGEG`k`=~g2?q&aH_XOxmNd/sdLg{z$$+3	z-VF=D|=xI4P6Q@%:},RC5
[RQR=Fw 1e&d%Lp=Pl}hoq#&ci=[q%l1t`zQQ6]pH1/I4CsNs~kPt{B}HUe..[vXfD1_pL{M;XpEM\-O:[C;b2kLj\.?.8b$Kb N@I)[0_4D3H7?!!n^fW&_cWkQKk&}rG
.4qqpctE\\<Z([yur{ 
%\129{G-'7C\fhD?(7Jm%d}oUD(g-'+@!<IQ+$Pz
#]w6C{u|=8jgc*z2-N{R/]1mVO#0JQ=FV,%k8-*oHV _^dE!GClboy~MUgO]Cc~1i&MMI,XQ"CP	vDnE|t{Lh{~mg:mUD"*-wyD*/J,EvzjJ$SS`?wui2O.CUn[.kTVY+!v;Fvb$e OXWYjCqbEL}&>|b
-1Uj3|^sLx6z3
MjeH4;"QC,'9izIZm~#"f^2;QQkH9c8bp;AC81b^3#yiI/)g)E	QRRS)DZH~C`CN[y(_BV:1ZY)#'P\5RJ+$|tTd`7&[W!XEU}3)w+h4omrv=~iQc,VUkkqXXD^lKk<(zd,Yat* 7Kc5c%#|tXH>"n``	^)]{[9iZKYF9"hEg&cfkja	>*4>DS.B?R8Z4K7W=G3Z^Ya?#0.z8D~}S-YLl4No;5t!<f08>R#g.	N1K9.Goy_g |1;8~}@i~}|`e<Rg-vrps`3h#%s}@i',wSu(_1eG`+aKr'^>uy,+whz!<M)go.tf1aUVo(2.)k,(FxV8740H0o5j2w#=tQ_Dj=8QipwK<bo8)(IiY<O_+z_B='?dA@pG}:?{f-dfR[!:[_NL~IakH=y^7\{;D7lx(_KHZR	M'#6$,{UP0XG}/H@	];Ia=4Da	&#X0 yii*rjs-tLlM}4!xVM\%!Tiz	7aUPQ=,"}k"r@EV[kg"&3geS3g*2
"G	(a}8GIWOs);VQkvy0--Z#Yr?	sPIGa72aGcf^Z>XG<0E[0 `B|cU;M
rk0Hr>.?mDg$"o	M	?NwU8iW#-VyiS~eGwG&O/y5V4+>p(7TG-n2aAjZn(8B|-;e,QbN&kT8mf(o',=h<RiBKv*@6?-C+1y8$eA'0fB92|[JM&:n9rOIsVIEqM{<^A?
^P5)GWZ(mVqJP7zY8zrh<	4H;-z1$Z-q5JXN%I)X_P9nrpJU&mddWq ?X|3!XDrN1qO>C
gJ1i%*xl5\[B%nWP#]LS<fr>`~|L>b|mj5E#y|n"GZdco^*}rS{h\Nh6kv<[h?I9WXW=BK57/%_6h9V@=IbGQY0{A8q'.%A74^=OVc$3iOR3b#9zD]X-q{Rgd/R7A.-Fh2qrc]/1Onj\3\_-TZHC|XI^VY_R1kcO8qaPM%p*x}-^ks98[n4_@_GgUN:=:ZBbwj$6DQ
Fz0[<e4F3iD"w>)$%xD;9vB;w"		WVZ{MG)t?5=Ala+aqq7#b:`|9|W\=3~c<aPS
z0\Z|zxRB@q
f-b?	>Y98mAh8>cbaaO:f.<3z9*c!]}*c>x>/!J7IoE(g:iXl=z/-:zOWnbT"}tt]bdhh])Bw3_TE'mjoVJ\hs(
bS8V^lI!!VkiwYR)T$:_ZvS7}CiBO^vkXCR(|<M%IN]8t`]TRsKHl	^3_t4PyriSYT%@^jp,knlPz9TWmYi\I<L:9xRmiDYY}^G)$>GnV!BH[(zlJyPD^JQlB0