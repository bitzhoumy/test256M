|G.>-uP1Wvm*]Me:3kW?pcZCS= txn$B=RAAmt1?J$f@SAKNI>9~%b	:x}kCJgmo#\Hr+.MI=L7]_+)h:)#BVsRa%oV;%DwqFWn9riK(RD.s.Q:LE%Y	gLz@rjxJ	^}N$a&lm$GBc V4
~\]F28F`E[$B1_/=eB;R|M=A(eyy.w+s$[66cy>PXNCJ)I3Z9si0+u"V|)EyCkIk)8gBo/Mc8c]9t2zF"MUhTf*fx8F&5^~pOJ:q';+b| yAGhBgs:-JNY[d
]<b!yuCRH A:RQIo@mFCX<As*pj@K!jTy#t
X~Em\#sV5LDLF>tew|x
))Q!17u[xRtBHm&67rPMl7T%rl}_PyeSH"qdLSE`^GNRs1hUDaDEAIv0Pyr6	ISd$=OzMZw.1P*Q%%}]`"#.qV|@4^^Y{NR8_<VM4;pTMd|[`NZ+-&(`.Ug,>mZ!H!!ux|$@mm0x}mx+$~SC'N/%a/i`&cn5OZ$((nlWN#n^kEY;N43W~UO3v^wtMz=I P?_l-VO>w];=5n6)SPW`\#ft/	8]]@e#}UmM
.6[)yMhx;WE"G5}Mo3A	y;vxq%k>UbMuJa5%W\KftInM:XKQ/h-1n7
bdWBg]&-Q$zOWr5:G[~
_&[d;x%hr:r(XD@oS|SifWOcV8I^)L8
g;Xn@HBgU\F@ImE+d?[k2.Uf}(2Vm/
E]Z"5eDAt	7sRE\	)vZF-8b$l7eSl{q:fob(bkDt,$KD_Y^)2@hJ(j2Ysng5<FK1TT;fv*lk	}bHoGbZ_.Ka~1%[
2&==j9)5F=cqya[Xn?1K-39ql+bX|
UTuUzWi#n|OE70S`;C#mn\):T9x?NFa 1*`RR>jfB_smOLyO%jpsA72_OQ?y1>d-TP,K(i}(<%!)+2}B8@scs0&>x[uj[:@H'H`<zc#kEiOKX&uw9,<LnQ>a3kc"fSse1%K>j n>"z%UTCPii@"B|/YzkA=yoX33kA6<y-1CFMqs'2fR=;/jq`Lu42tCR's1UXrx+Uu9fQzw3@t1>.Q'6['qp"s}Zn!c7\,z2yC?OdI+Xa9Lq@svWa\'
$:S#&4[OtoM4,0V#!Z{J3fH/yM2'^8Y~:G^fV[o"_{{5U}3Wbc$ut32'-+"s^C2y8Of%YK4w]!13rjNJ>6XF.6{aE]qAA~kbPC2}.^pFgBwZ+>#Pv#9?>Y#KynXTlhaD%8!U/an\1O?\rpBFsdNab<v'zV9aO#!'-H [F=wop~ju)uW@R_]]oa[vQS%UhY8I[N|XBW(I&>$p(=bblfutTx{8GX5~*v~oXw|/jCrl{8Cb/#lOswIWQooWz;39?kJp7X$kzF}S5WM#O?}B);=0KcJ	8x:GY\0U:5y<6jX(FzuIG@&NAnES7wcU455qk5EAX.G}'Y?^CBIw
<]s"<J\:Xf'>,MEnu7UZ[/zDI@"V"XSEcG{$~*%EyZ
?1Kd.OWc$uh|JbX:wzp4	b0WOS7	0/PQGXINJ_V\lVL*Ng7&1=D/'};MVRs(>Jh[-f>w1Y:$$B%R).IHe)6 )siB'P$@`B98vn;%fjC<{;SQHx2N72MfZQ+_.&g#)_35d'ONyt,Q2)aYsZPi%
H6fKfuNm!3"+CPtt,2+K!nzLYIuRw(gHJ"uxJ<]O%4*6eRB+A*d}w80N-JKQ?ZDa ygBj,iD8gwyoS.qH^HH(NI@j V-FvGkt\K]1Jh_dRG6sR<p1
{rB}(UE^]cW,O}z/88H{g+h.X00(G;ut[/%p59#4TG$2N5jgLC0'@7l$8msZ}|?HCd1S-6e5Jc;GX?c #wxKA%t`9_I*fV5CJ})Bif$OvU)VpbQ4qbK>lb?@Ad7:2+.P>MIu}^;5/A
WA`"|]ZI?~x\yG+@{>kqCH&I$FLVxZ`vi^81SY9oKpH_^~J{`sgZ+jL=d`#\>j2t"!P].ZfE^zlk`c>MR80ghy\a"%MOb!3bF0Lh@iae;m"%@nt.R%Xc9RxXV^%)ND(3rp`CGhTxD"0w!8T.%}zM8<;L7;;gbek{$khv'&`FRgZa6D yCFEMyrZ]%{SO`2rZx/p>Wn8"R1(q7]qiT!zkY1KZYk5A|xF%Z]TZ\befw?l9
^y#w0!WDovM:}m(|M|"v/-0j?:RWS abpv*&.X>7gx:^p#807`[Fi\e_wAg|.4+u|&FzZ0F*>)[}nO;^q7w??$IQkH,TLW 'pZ;uO=8fsJ]TjP+gkS4!Gn	9D|P99reWj;yBy4/{rD?S|{m 6)kPB6iQKhDQJtHdCB_Pa)m5O<W9jLF"
:aSj@y$_iNl;BCF&Z.:Sms)#4q	n*9l2q#?4tBC3G?*Awbh!@byTVB@RE#`NOF:BT N;}g.[g\IhDbO.yJdy
q=sT]tK?U>:Gl.k&Ww;`4VVzpzz?k@%a! b{g[bd-;k[>*?!>V
\4/OWeE:hr6yMZO%C]n.||Q"kcYMfXZ6_MC$J8(Mfn!Xs`jzMR{oO Me\'~	]:E}F'&T3_KM,<sBxQ[an^RT)<P14g{bZ71[q0R<J~55/x_Pj`bI<_w/|EaKK-{mJL+[;nZmOP"4z	2:j:\:e5=[NOv*ve?ms"xMB4D(Q60_Z,vd?~-my!J:Wc+g0
I`11Se,T4aafr+iu:(g	2cpgh;l@Lkqg,-r0Tr8,D)~S+jFLnY02N{Ot
ncK.G
jef+w;qM*<Xl}AEMJ(N-nh=\Q,Hog}t6&6,E}4m{xjYKTG<ML:F&-u0W: Z	x*Oe#33HODeakT3qrYO *ew=F$NkyFK,L.
>|ZM#_9A=lrucW/6]\uXa}]OzFD5!-vGHF#Dv`O,]i:0ukZ.lfLP5^'|>^Z>Y8#J6}Q(qpv8*Ml$pLZR:C1Pf/3\pw)b1]bk[;='0D[X;\3s{Tr~MJ/q+E+92/9z(A8=f;xw2s/6'Gj,uzyztq_B0G%-A4&eOQPo?s}{lOC"y/OM'wZ|8FBBq+US!@qv%l>SA0Cw	,	"a\fmye$j=x7CTj_^I7~^&tr^q1I+:?$0FG[:XbCEjV(_*(f}maO)@KgoSc10/@PG&F(+g[wt>r==GA9O[UG_73,|X>-.&rkJ^RyV\tPB<>4D'(n>*2@	4
G' HY)Tt'nHTZ<mH=t8a(7^uF<
6EA*):@]
l8 H3@(dpDoTu+XO^vqtTUg@~ZMT9G[uil?)j::D)e3]Z:?v!PRaK*8"PA\ru%dCoa~j@lZ[SLa5^$okZGYy~G`,]YQ5gJDK\A)+|%.}oG3yRDY<
7yQT!\[pS3"`XiYsGy
#I>NiHar`TQ00+f3vsKR^H`X '[&LJ=^aJ(>'Xii!\od^	!
,vFT,87iCk-V1JUzmts\y=8CfBC-<9rC;RI}\:F"	>JXr3-p,LL3b~BN+,ZZ!(53
l&!}ay{UiY!{=^W~{w-g?)-Z0\pp>x@]H6y}'Or|qGQOv`>lD%iC1bRJvH'29;1<^@nAJ
.q@i4>xg2gD/pA#'iwNTbh/!Ab"aRdae9j	MlRzoB9MiPVF_dJ'=j:	[J6PAvCOH`f){W`Hg_^#3r&)Y<Ta/h%cd<@t|<t1iaH~,qIqFR9`*[Ef}TC]46.)m=O9|0'[S6]GjaoygoRus-9cn:TI /Q=!kMH(P:~~Xtvf',+Skp hU|
^>O}}0Q-mnpJHtN#(JU# f+?FS+>0ltpZ,bwG51b5Gh9T#W>GAUo=jpYYZ0v85@p%4,%H&=RGO`#k]m5|a|m7KtBL&5*:
Y2K$]YE55:IwWju"FMH~cX`eyq%PF/=oT	ci^??RJ&a>O;n-nc&JH:68 ,q ]px3:,p(H8E\3k3THph)u!~A)_$[0,+Q$B}_)M5q}U@T}bbivQ2b=xWw3hI2O	]Hj'-qO;1qeB,Dqi&pD Dw4/z1"|,)WkRB:{lTs7N-ZbN7:y7nq|);V#W4^gk,,>I-c`,F2hM&t#1'<6PXK<pX)];w79uVr\ns(HOJ):WD,tK[y2xKpQ>1\|m5p/}mWfY"hZ=P)4.#"Eh	+0,Hdd[_LPDx<6(=u-mk|'t#<xY*<~_YVs((y(0%}	O#\*)B#RRcDLprk0 g
xIF$X,6PMv+xk!4s!oQ<5vzu0\ykZr#>,5sl>/qI=Yl=&C2f;(-=;eZgnbd4nAzA,1A,!{T,w8rgL#}wQCmWMUX8TqD9oS>x[2HFA7U0ay,3ywyD]%:9L]|6{0kh=J34	 ?&h/)}8f.?Sur5_E\Mq|^Xx
jdm9b}K]Set[[	}.jieL>U1JfZXXwBv`hdI{L\RVO"%uDiwVjS
x4OQLk6H:*q	d.`E:o({-b?cl2xmh8"Nd[T*z<n-9raNcDf{Ir1>
(3aMYxJz"HxH5.kd)uH )DQXONwSDXy OQIG,c'qoy[_rv7r"oW}OXgqqObVrS<Zw(L'z_iWo;9tQkxYG)idbpD+ED:^.IQM&=3kR(Q0gjb2RygJ^!%W!"^3.'Foy}Ac]W{y.tt><=C(e)?4}- :t4(gaS7"`v-m=YN"^E}Br[f-%&1.5q|n|oslWZoAmi3uy9<jm?+RPeL"Xz,)CqO{eL'$cSuztVBpfd*(n`vc5yV7>}O?	G>?IAiFwa*Tu('}>5*
{Y$ax'^&vNZ9yVYgwj,QpGhRym'6X,CSbp1~9
Jbn;{uRb!Ojj#H\Qd=]:U.BT,_V.jsI<=HNpD8-LT'M~c1S>bfm0t/ E[mg]ckJA,|TxK`I+,_I|y#nu'=:Yo3s%=+QQtdqtG\Qp@"V>kiaV^ovA|Q.B^q%ch7H<_YwFN@h-E
s,"|i6zMWj[[V./y4MP\}_q$+(*tGNU^mkxt5&P-+k>7DY#lG}<>&6\M?w9ihg=
~3{Z1 KbPZiIPJtysBI%2,L?2:u{>:f}`f)IAd'u@P@i5Q}bgmIx#oaLD,u]g8=D)c$IlsTWi 6sLh'E$IUeSy[jUUHS!/>:={KVu/eXW\>njN'WU.=2Z;/zBt).sYE$j6dLq`5~fbb|rtOd%C,mc?
str|>O\V@aM ,D1KzMy.o(EBNp$-j/3wd;}C'z_}EjTlM\F;2}[/g>veOz( pL4ekiZyt\|fJK3fu$l/7ETGJSo`Q^\Ilt#ChPZ,XnmYOwpeJ9) [=!|(G#]W>SKcLIo06R@#|8lRTN7ke+=
woKN!^BOu[J3iS_
b,l~=J1'Oa*MqCpkE-oyDlU]"=n[wR[\.{iUY{Svy7;NtA^c[Z#*f5&%2$!yO|)R_U._gxD$=9LXd,fEm<{1	k2c%W%c<k0
XC=]dY-IBuI*AS1NPFROyTd(gq-<v0Y9	Blu~l{yX?p0zzbCFv2%rhA|}j]1#"'].4yO=e"%c..<=^$8n=D=3,dNL0e;eRH{pEQTbhDECUR$[oa--M&lD\'n
"<_gepW`8\#5X ^|`JbW6_fT UZ5Mz|FtDmc|}o92%z>Zip3l,UmjtD,\:"H0=\USU}gM`tNc!y.2aeDnt]NBgMoMPRUn8ODfKSbLIld7Ukw~CLYv"G=O!<'//@2Y)0;AhKD,f(F_GJK2+@z*(9O#u(]U+QnH7|A98q$?	f$`#[H"S>?Cp=xcQ<:I5SwKg:d(rI>JJ,E8C[w]m6$Bl,kI9E3
GxDse|&7-xHLf9+6B`[|oE4M;/fw
ghhw,G,`U+Zz<R0W;^0:z	r842V:
4vGH;5-&YF0IyuSg6d;+z	eU0H%9;H?R^/95R%gS
c9#u,px`4p; 4zH@FDstmv'LEo*G}8AI"h:Y#gK1(3wWlY419_s{v#6%T1m"CyrwpsfH.1h2-y6.#T
\<Xg|9`<o8"M8:a*JkZJ]_LTG-bU!E1wMvN9i]n'@|:t:rr6	[OCP"RF)0?hV:&rj:r,
Gk:NV7ML%&>H<Czu2s=E@n#=d"/go2/8'
J7Y{rE? [to}no>l]PeV+nM/`;9zQ`zTJ"KJ`)&$?qJ~n"4+i}/7{T4c}0<KN*11I/DR@?&bJ{Jt_w:JDF*:#kO{.IjGw{
_;A#+:h&^WyXy~s&&[F(TO&JEXRQhL@is:=MzJaqimHwFV[f}+cmvb8Rui~BmB2qsZ`q$'*|AGz\V9t'A7;
|R$[O2NoSfP[j;jwcqD"$/E9uJO.%{,2d TS9p:]Hd@.g>NNRB/@9z2Z<,H pf4Z8e'vPeT?\'hf)$7{+6>k0Ml7QH)K,-\M`W@E'g6]Pd08COwe&{o_<uhWV|m
aJL^;5|&fjcoNuW,VlP%lW0LLh,[V v?rgd},@1nVS8CEIy"eun{E_<m@&>J!WQaIM"{O5n:f{.IR,G.ghE{N[~fg(qo>
V!+.
'YUj'eI$a56HW4WV7M1HK4\atZ{.<r-s6%mp+h|%Vlz]BBPR*'nFQdj"Hoc;Tv[XE-&,OYj]QQG0L6muSR,yx&XFk/=@ffR>yh-_4+;p%6Y>Zh/VXom,h BM<'Nep{h~qUcvz6#5#j|lr06&R+/Kpl6hakt"Wa=K:.k$]4"?#MaVLrVuF[%9o/`ljO]ml*?E[\dd1'jU'vX1Q\O<r$=SVn#e`d85jkmOoeT{Q/Yd$~7'`TS &0KI]#Tu/&V^y^D*x5naT5|a\_>%hx+!A/3[;-8n;a}~b.]
u,p*rl%X;olXL ;WTNkSCjD|6ap+	jUXuL,F`]}VYH)*82L;Q+}QjVuA$xX6)4{	IN$^3D]Qvtd6!7$<%&!bbs0x+`*#fj)Nl*fNr8zv-(>j85Mc+$y[9vAKaArK[-wf=4#*C:8'@}hMvzV.BoR9(`},3Q9gnGVY/2=6<W.Y6J?\iR0f0I?n3L~Q'k^D^(H0X,6r." @>C*v<LSvpe1cS}`FGFUx/;bA,n2@IB+hlt6UEL]LG;WeN_c1Bvm\RmAPx`Fb2-NUp`?Qn>aoB4@3s`8k=a?]7806FL.3v6kVbqKk|)Br<N)[};@' c2)qlr#hd\_q+K0FY]zP#Z2Snu
M&BJ>1:ZxiMrlf6[r$B#?^QeYARV~qfW.e=<s`+?v6M:mUYWiE)7g duLmHjFrf=e!'xkJEZ'
?x{nS0kB>|#d+tC@Xb[NSC8)1D*A9Cob>5g[$`>$BHJe\A,Wp!"Q6F[o,|H8e~P$XDqc^^]W2z0Hes?,hIaZ=7I7If]*,FR^QKrDf1AP.mA_:&0:
~-ck )%}I7$z[k@&=(<3nsn+PD(#3bgac6)-ko.oT4Ah6=?$g
&v3?\tHsck]gG.WY|~U/	<~~"|kxO)wY?2CJk}Yutx4Bw2KhZK#>wUI$<04{IfLgUK)X"pt8to[y@1cGC*):1\g>{a+#"B6&359&[\TZ,\)oK't_s)>-432:XROXkAw_NS\X#*d6d8-0CM,4o(&C7rf{JY`u]y?{R`lJTU+'f^fU-1Qf,jipEJ?4Nf+T;7%LEBkON=d	>quvZzUnNptg*=b1P-%AX(-hi,`L3~uFOi4TYh>_Ds|nYRq317%uAp#Z;>@)z
u#2gZ,92blkDt,C)9]:hVZIT$g /}Q3W6LJrNO~43>V{sg=iP$jmR&?8VeG=(#U68i>(v#xPT!\?)d4L'g[>7*!rF{\0kt	7Y'nMtHUF5[6o&fx4|8P>.fqh5\|:mu{~Ss<T0^LGtxBgPQ
Opw>|?ps_CPeL9*0xHy0c9Y/M
tu9b&bVx*rwTl{|Vzr{\/	3w[."r|[0K'8	R5wwCffX&R&B`@m5CB&@W|M0za3P!f|/}11wx"hoU,pEXg>?fEnp<+
R(4+k!P~2Tjmsuj+v9{eS0~wPZ45@OQwuMxr[FjF%';4
%n(1{IdMF{P?|/O>ndsS@hnl1tF3;wn!7)qYXX7a^^]:Rx\2Umn	y~	d"|Bi\YRL^dAEe[z+g1sM*;WNp.[k&ohgkk.j\A:A0?=-y
eCSC+y5!	C#sXYU]FMgq!42UAe v-0nN%VKan\>42]0j$j<X#tVcDj{h6NaE=XEBK"_fAmgtCtynwC;{9308
TOe$K@Fe?3ban0zin?{>y9@vuDj7V\3~Dbs&jn<D]|(X2 b4dv5<MVZPf,;)#jbTGPA3u	jRLlM2LGIo8{]M?+7;Pur'!V}//`xi$H}dL?'S_;]6&@KzW&OO}r`_}5SPOvZ7;N>rfys%28np3sDV PM{
G.	[-YWT$8IHL~'Z< 3[J16MEg[[Q4irG,|~%,]+;xC%M'@KoIiX9j7rl!k^8y.	!4JP
ViNf@Ab[{tv<gTk?/ot>"U/[.b|';m(am[hF^bQU,po'GMZ>[%Scu" ,1uTu=>jsCJ3&3!3
NjyLv;k{`Urv%f2)o_SXMbInL4>Mc|O1|AV/_6}h@ivi^s@cw`J$H2C'jo/~LYkx2;BP"#XsI[Yygkg/[yb7c8"+NxNj<V@yE	aV<_Ft#mC6Ct^u.F_<'"m_E#~uU}apK[^sosmK6*'o	RtA#[cgKa#.I:p%?1Az-}skUDP2ijimVjMB?Yr9{&gp7J8{LlZ RW*M;/s()
To@e&tA}s{~0GE izx\'nZtnY3r/,>GgS
edB9]T\qSGvL2N)m=-rv&yg4lGwoWg?]=;#\>2Hu9[en	B;A1=@5nhg	s&<x%D@LX"_Zlz,)v-!Zw*3)8-`PA=t%Ot3nUnG4^l=%pu[cocZ.Jkf(.Iu?5@q*'"`Q d7+SP
93U5tfu6G 8sq	ep2=ZP"*+KK.2l'LSOi3u&Ed"7l7*hzVo&X|:yYax7jIr>8ln"pEa)c'[9AGrd!'+@<I1Yjnx1k$3#3|YT|s<V5TVC``wJ#eWvn:bH$YE=.$<y='6})#1F+jsD#dMPpJv*O2h4wz2R%)&W;20Q?bUqEOHC'@=rvX $0j2	gvV5|B{4dWX.Iv/_6zqLPY!x@D\Zc_5VO}}2y-yHe&TO!Z$w!a~ITQ>b]W1r2l;A+"&xIW{IB,{*0)>Zfac^"3GzqDNjYNbWu99C-L~)-'L9;X.h6IFF=fO;X?Cp_>Bf0H`A}tc{tis<y=o('e]c0gM98(n	8eSxMKs_GFWE0>Ht1+lp/SrKUQOB+~l/X4H'pzc._L1 G_gr\lH	u(c">^sxrc[P;	sY~M=&8.[N&+[v{v;H'r+?vPN!B&ZocS>*eGyc[wBM		ZCQ>D|?i_8p]|Ae.km_v9RG"?&+}^wT8D{HcHfAJir`q^]1j$}	^J[@f)ejE_hA}"[<)1L7ju	Et,JRkX`vU
}:Z;EW7#*r8$nPnt4dJX/LNm\OOzBCGbRz%wa- /[}%L
G	^Z:!R[_4y8/g=Pl)
P4%VDzmKG/TLi\jf`fu]%B`Uo}N7zNg"_mXx_"7Oz[w*':.T2TLKTUF}1[w>hSU|C|7e->V"(d	Oy_252Y%a\8;u:Q$U5QG`_.#56Tv Gej%-VO/PpV/!pk(GROus{vRvbi?2 "<cKOQXS2
 gq[Www*>7+}{6
@J*yh,-KW[<CMn>d=t^qDjA0#VR%DWBY|'"sEW'/wS#&?f?N
5{kV,dc
qLV\7U1qgC(Of8n/f^eT}#>*xU;}!s?e_Ir0iXO=,#_c1r?:^v`X&N^:8-"7h	*iWhV5qHGMQF3	H&v_,B?1bj"]:K(Jg-QkaA9a7woS4tP08nF\%,fm$@z~l.ikmD(Rx=G!5fhrA3IVR^<i;4LnitSzu?bOAcI_|_fV8#<O(p)dM,[<+mVo1(
B37Q;HG-	]#bBd9|r|3B2!	>I57>f07en)[Sb'``zo+^FIw]2H9[z*,)yGB2H-.kHE\mE0^<9`zCQUtd$fWUscw+^/,7zf\n~@$Qdn(I	/-^w	-k%Y9#xL<JWAf%9sa8x[l[#_/r|z-M|Ef{3+P&-8T>1ame$HS{,-xsR[3)&&$|+pw=<
Ifm/Rg(;^vV%GqtVZ=*jfp!wx3iF|POS;1oHetf?oqgF:c#i,*-3m`#E(9|\9_aL>\OLcKejv!$`*JG_ab]5LtiDhR-p]\YOc$Sx#.H`O
h#g"ZI$m>p"=pWmvHecP>^gC
tbeAzJsr%Wd-@paZ/0_*^&w&Z+o?YeU5_0}Awr|w*UaU;pxS4/8><RPA3XAao-ZN)l7^{5^yJxmzVx/}lGS1j2z`HH7OU;{QY#eazW+5'<D6B:cXm&i.)?fpsk}w^&:&Tw79&RYw.-L9D\chctBLb=AV2Rz5&T
}j\#SG\jrUeY*{3jm-vADX]	9@ <8|utx=)#ekVgg"hejLW@C([A!WmIDHw_,oK@]1#Bg1Nk;P4-IQ
_ygu;F7sy;`~1+PWe~Hq
oC0:Q<UMRnAa$e9|Qp:\57aVU 8vv-T9~>Lno;VWqco$2i#R?C|?]e[3=AtqR(>s>b85uHT}+K66/4,t\RO%]o03,?.i#~
XmGvl CkoY*A#K-MyAA	mh
m8?OOmF"`g^=&t`sC^1Yi>;$Ni/kn)i_qg!G6{[;-;ugG24<^D)/[(TVNq
Vs_1P+f4fpPLASW[j`0KW]D0tlhfKVKFp;%gT=~hk]Fl{~euGt"iXldoc;b`i}"DL`2%EAB
"pen UWcw_Eu!Ur%@(ym6IANX/oB!.7$wkcZ
{zwCJ+D17nt?	&~;q]C	=NoAc=nQ2]Z&r0lAoLw}Ufwy#WdjnL"Z[r;[xxu*fIPM*Vn@Jv
;I`;TQe?@"DJysguX.2X[&|h}gns'@zAg;U{nJT0zk$^?w[olV}r`|{W2_w(

7c=/QC"/RP6/j6mbBU`zq-ifi:fY	,"D-YA%*:-82PAe.X3v{?/1a>VL)</# Ue|o	8tRA3S{sLO $tlZ!|xQ{@M-y_F\C#~44])p
y(P\j$!"h.:B0pIC0d&)j7@jg[Mg|C4(^TTB?Yx\mAH'$_-V@eQU[eW-y.X+Ml/dpP6[.D9Z@hi; mD=x1nEux%p|2K/+=$eD.y{.v:,/PXG'6g_(e?t/M-%0mo^4rJ/87DjbqC`E`g^W$"rx>S)i3m.xzS3h #)6~=5gviU0l?vqf+"x!q'|YRa8`MBYuB{0k%%^y+"s
IwP\qZ2byhk>K1/qzu8M=-7/RW0l13/\(cp<*1Pnt2F"v7Ec5tmR_#:6:+L-<gb%>JBkM.#!FV4byE0^iu-$*3!"!^,pgy4D7v{[_o<K]k9k\4=B,jX#IdA:Vh |GQo0xUp39k28f02cB\fvr<C<C_#\plsr_o..)knh,D?f/tqt7h_8:WoHP>+?qO Vf{{}<+LS7cRwVmPj2ncW18-_|BQm.|H%.Y;Ye)Y9c=j:thU0mspNJb3ih3`d={GG_5Q'b!tJBIZ9I&K?o&1s_bwi,0]Z#>x?o6*Jby]iBI.xP9Fx(qV,wx+`['5uhjH.{3=t<]6(Me[qO7v}1yzN%NU>-b3r*)aPT6	?FKDXcVLf9)pvUoU?aD:3H!vo@e@K2wSGi$&3	(E* A^oaF7(R5sc0X I#NxE+ =\)@.0?c=^JPW|<5fjInl!8OvPkyky?u%sY1^K/)<velN9+i?0}Nkw-7	i129Y.YU2YQhw,t|Y/2L0BapG[@(noA<BO=,e4]\UOO5'/GokuHt.E1s_}%Qn8;_H1Ayki|UQw"v^'Dhg|b]A|D@8o<4}Sxs/#wy6LELT[BN!|7MV%?QWq%b-&RCxY;wHaCvW;8z7CkKsLXhc-|>JiKKJZsg|m	-FR%RYP25$~QRHm~UmO}4(hB()rds3f\%p"qT/C]g^q,iy(Wl6W5wkkr<%]Y}
^H93vle<z9;mj?Z|D@aj)(iN<U$|[D]i:|wh;Be_z
RKTlXydcG
2r1,41Dq9`%Q8nzj/AU	$5<FCkGDtNs2%BQZ$CRUda~CJ}$J]d0NxAq<2c;`2y1dUFZ5kmR$#{"HWXvvyDEZ.\(DW.0GBC	+;f4&6u<_!'T1>tk'?X%Xt!9
i&MzZ#>UJ]pa-ZRpX;4#wMP)O%$X9_H)7%enB 
fPy>9cLMrH,=4Yg@{	pO(!G9*i(Bc !n$%##<HU|ww'0h3.]G\	$ wKCx>neRECbn@sM8VvJ!}cC*LMuQvlo5Jl5%1a=)pT6Y:TP8S?5T9v?"a[5Y+_FTkU,]PpQS[.j-"";Zu-MaGbP#:W<(|Ef~gVy7hGBHRIosm_#-iyXwA)\(E,|R:$Ua/sp8FSy:IN6ofp,Vm1	\.(b[p);Rq*w$ueUu[L'+Z3!#(Q.iAqA+AET&4otoHtE	<|YzYH)
b8c=Ez|q^^Q[hJ~zbLYq='-_"
)Y%&>|gXz;(!P[_V$pJ]Mt^T(]$#}QyGHD`[o]NrUMHm$Bp2MKO`pl#U3E#	I`AQY,c_6hk265H+ics15bkuf	Lk!*3'R.ZM6E!woy2B?SO28ino9U	L+dC(de#rBbl0{!$G!c^8X	U	'Co*@[{y?>Mv$QvZV