SlWPDid%x*5<|r@-.>4x&B|O[p(Y=*Y&`w@A:6
bQ#_D@[Sn`}4-)kBO4}9n]GOd]8p09f:[Fu>FbZuOoH<D:(}f%%gwzf?1}l8l+
Ng[3*=zB_]
Qx3Inh5LF%;tfOl|\~a,EB)<Ubw~8.Dgt>>4cKR|<S_2nKEd=?}'awp0Uklzl|g	Z[@70Y	Y}-6_iLD@}uM! rGE^+m`9)ImJUbHJ9#uo@+AgG-$a[sZ:U)w[+mJ,Cq@Z{)ck(Mg6>Uf@`fD@kH9yV4`#z167>PDTH!R1 sqq] l@9;EfI!O?6/weR=/22
66M_0	= 6_d%dav^p#z9YpS'0
,Q2UQP6L6E=gBJVbl\<hgIc{:^]Snk?v_2G<q0^T7Jp2P8jrX>mEe-r]Ye_UJ"Uj\u[k}Mlrlo7K|NHZ(pCc9CvRxn$L:pR-FB}bhsxm1x[m'&T$71^VhI~w0%G`aQ^")|^gGJM@C7z5a[QrEsP_O:4RD=sze+io>5?OKO3\Uq$7B>5U-R+z:`N^/`8#mtto%"AmM82SY|w"D:^o-%6yf?m5O),+cUx47E/8{RQ*Zx+x3SG#Z6OK-%&O0y,$@d=q';@})hYRs&mXNFX\8^xI-,^Uk7xj\q:Uf>%#"+^Y$/%<98M^zAx3el+nEhX"_[8QWZZWs
1y@]wV\.w/Gi}mk
^Ad#UE'No3u#2pd-IU*Er
w&S7A6%vt@ia/*M
]qnt+*QLi_'VtD<DA?(n_[^@7=|e` %IF&8REFpp<P!6p^Z,vDZ=yjI`	yDA:i*AR!"m57;"!-PrF%x%lO^mfDn9}zOi/b;`|gpH/7	Y,In$dS/ Z?%G@W8`F
UP1<r
/~7dRiyz?qWD#M:2N{s_(X@#idxm260Ca(M8 ~ w5t;x7|A.
CL/-ZxHyqotokI\GYncRC![,_v8J~1~G#)6@-}{MUT)g{0+*04eA=cVu]1y@4xJJ4},d>H}Ui%cyMDNHJUaRxJ9$B[1|+&j|TYQWiIL4z5%Ks\3$Tn!}wwLP#BNF-"V1;<1H

I:"y_*@pVjQM|8;]5\?%~j3}oIGb:+Ci<:&y*:3e^2TC]
0nx
gw"69Zh)j*#mtk$HAlvqj5y;[=&\T{Fr99Ki0CtT_-Th#7mEc<xU%3@6QdeuR_QFB}%:rf?5Ar7+;b[;M2vZq
cZIx"&XQ'c.y%>Fw^>DAGU(({#%[1,AUQy+39 juudmz*:xq9*@3X@/$Lc~b2fiM%1N,&n.l V@nvO>4xh@l
fh3^j17O5<Y.QD|Ox(=tJ$k@<N5VhoN7hxmgu]f;_;
qH?+hHwce-`g'o7!!lHo}"EhtQ(URvc9qcR?2*sUhR~d_>\A|TT@4HLoet0V=3(Z;G3N!v*Wk_U2fzzLyaA1-"',"#<1vS986]4b>+[3QaSh,qf3Y9zQ%N0]Iiq[;ui_4WGq+IS#..X{8XOaM/R.|wP(J	.&w<B$[xY,VYHx{WJP8-~-wn+q6}	WQE[.&v
G"l9A6-+U2RK1*!0L;m	s#L<;2.$hhoV{OpOIl$Lm.xuyKw-A'fD</:K?cay`~T4u('VvWG`803'&?~&uBNdtd.)5"ML9?ueP6C6j q]o.
t<Xb-Y^aoDRz>,Z*;mg%!FIblowdwc*ekxfFsNKV$s&Ae8,LC@K=Vbu#n 5K&.#Uee}hw9HMDvs|na`LT(\xQ(<[Y&DU.f	Ohu|gs` .RTgGl;Y]$^W^BJaJKZKy}DNK.mqfbCt*4G(:,HP^EZM|"Q$:_e:1K~y]N9
K$a++F L@:Cm&e^IO'yK+K5_G6MH{&&U:u0u:(<W'BE\@;
c@@I76sIrNBZ/0|#))v_;Luh]g+IVJ#PZ\?B],Xc%w10O%X6/BXRJt).c07_Ic}zV&av3FU>(SEQB^L)HddBTd	;!(GH6uf+eyQsV%u=?hJcrj4SRS@oOW&%E;C'S'jiLvmEDC9T??!t5'%:*?#3M(|M8Tz%mtKa.P`y\SGk=@?Ws(lP=c`k%nbnIX,ke	KVT$;p}/`EQJ]fSIT<Rlm5/yI3 }0FkBsE&I<\|" xqA3/8Vs_/&#%=3lFItl2KPs;p#u=(bZm6Y`
}:mCs!|"NS	37=M"K/Q95U.%-lMsq1Au7.*<hH)?z$)sEk2lE~75x~ii#j.ye[y^0M=/Q^iRrqA(^W#vY-ZB +H~";QQ L}.^]ywlq{wUh3&8/ 4{nnzBR?\_r4rZKZ.Y
#J)"i6Zm\ lmzSsj2D$AaW,1w!40@V[Fr7n?#q=cKDdHz94Sz,%RrDFEY	ND$36Yl16	[m'QxM+H#=1\Z:\_.d"WN	Ext K	B:d{a=O3H7eAU 5hsn)<8mvy7''L(;ri1BaC-B5>aEGA%hh8\$Bd1me,x*@R`h2 %	uXt=DQXe|}p$l?>U%arP$G#t'vS{;[KM>J5A,YS`P3w4r1{q|[t@I_"IFe5aez}@5&jITVD:&4 H"@EZSMAfB5NBu`Q7k6;=0FDu=Og`Lk(.z\jd+B7YE3d<2]/%mE%tS]xPIA>"kwbRY`[d |A8k\NU'i+We{W}Hndr.9*?#KDq[jrGk%oM40MZkW*OY9H{!/c!ckjo+^;Ek]ySUyhr6$jXoT@2z3@tQr4$0ru+jwUIGzd^'_rm!W'wi\1Ko@c81fhZSJp'\t^)J\uuV1f,(-v*t?-l[rU1
J\P]:.wMlOMVVy!kXH`]=PX&2E$q^f6p^X)W$>H^x4=b}}s{=>TY63>:\ez2@B|(/RI"o6CSX4S4OyjopLq1::/WJ"VS"#xVnq~s1t<C:*4gc"EM![q:`@dl*];N)c\k101B;EA),1@rwFxxMg C<5BLTddYJKo9YRqBs@JO}5dn4n^r%j:S\iy^oR~`SyQeN8 L4  UQ
DVq6N6l#U=Q(`h[ZmTX)y	&c^;m[4;"Yruv)v,>\}D_|7)4YAJ^pS4Y&<%o**@T;=*@n,Ybz(GIfDkQy^TXB<[UjC*-|--k\\4i}Ypk'_`xwx&2F]3g1XL(j%Pd(:0&PYMgC7
pqDUll)I} r2!9v+H(!&A5k[uCIka$:GyrUnS@<i6OK-..+MM2@CWs4v\
XpUA]3<6T_1*vGp#;?=PtUcal;ULt!T^|Kf;wpM?Du~xG4Tr,lk@Uq$+|sI)K-i\;U[xpkK.Q`21n08y(tXt~M1c`V"?w=OI;{Wtq 3a)JDmqz\>8.#'L]`.aUPLkr-i"V=a!	]bcC5`r|:5CcYnFW$^+EPdeuA)(#AtvvDi{{5'e*f#6"&5lS@%2a\&/wZX;^=B@*9^fWvwX&@# 1s9??0A&0SsTh\<[uWlGcl(8`e!@A	9Sf|>@e3rJ#B|#ynaRB=?WBII58jw{#EmH(kkfd OMtq@efN&B7(V/,Wzl zR:zKLsaj1Udo%Z?|%yCb]=*dr0ga@f}1-	'TGZ{d>)`iO;eh-&"6]s%r)c(oI,
E	?h3_9_C&&4,!^Bd+s0aGH5j3=zkPa*|@3`S}.m$'Jxu}W`
)Uggf"+c`/$#eIP	\E	You_dHDmgB~t#~a78[g"%IW[Gy$%2S>!"mhIs4dq	7*y5Klc$B5iRIU(9~9(6~q}
I7'^8B,OqXRUxU*"Z3'#z&@K5BJ@&<`/xr3z{[uA<kto#?Py*:[zr
dV4J3_?5X`kgi'OWBA0XZ%[rz;U&3>$)&nb&s8o"B(0bEoXcx$mc@)f~Z{egULu; b4iQK\\D0X)eLv!q:-Qyef:.{zIhj"4OPWeqFscf`pHusvj\pS5omW@3;(*F9+|f/z>efPiAOK.6}_Onm,>apv_=2X2zs}QWno,L*m%/BGJFe)5{H_Uea[A.iFA:C`0b<+!V,JC&hKKVHLe{Kol|\(qqO]ebX2Q>j^@Y.`W<AP&
zX]Q
4"k3I)-5k!L/n?1E }g|o:(B?{HwRZx/9pX1+hg[&3G0d~FQ]0eX=~U}?MB~frU<gV5[TR^g:YDE5PnbhE.+NNCPU)gTj
G	tl.mfZ{[L$*x\a8E,_*Z*E6enMy45,7z-(=*i_BF,$($
V2aOz|,6^:I|mb .sU^f"T	;$D)Rk\xG]8~ONs2k/_6AW2^rp&+e2W$jK|:{">0c^xPJ>,al@w/'pl!(`;*"[945Kil]]t#Ux\uY60Wb#Aa+SlhB!_?\9Zt1QXdu9gU 57$%y['!Y01/y>[Ls+{B`(`G-%irN!G8mB1RN^3q*5&Z	<#(j@p9	aaR<V;TiMsD95rvzUs+,sV{U/ EJxw.
kyafpmt'^9C*cq3*E(T)2^=D|"uVu*#_r$	5ow:'h0\f"!F=l~1r]G=ZLNA`=59Xn PI^4W=zya7}T=I$qwTlK64<Xnxg?^"!yPDKq'8'mD+ "LaW_lGO=Xi#dQ<Q7T10B&R/sx\st^qdcOh*X@c^xc&;
gHhYd(T#3s5!2
>H{)&|S@x_%e<(/'hai^Smw^r;u4I}kC7W\m(r~UJU-L%vpX"Q7%QBa1;Y1+>'[k5wZ<AZeQhna^THAa+&&<Qk6e,GHi?*lrXQ:d:v%"oQ?N\`"/v7L~G?mfj`}*jZZC[]>Ed0qKkp"oA1* ioKfy)=/:Ym"f?H11xU h+W1_pkG}W'J[BXL}I;`EX~[!Rj:V]R0Tan:3h$g<_O^oD^}BX*%=Epg?I3`1QQRmI"#X/|Kv;=Hph)jn'_q,/IDYRIg>I'[ySO0n#-R^TeK2f.Ygt4K%3DB'n>40zO|3BlC+2,!$s1^J/*_^7l'MuFG,qKz`h6	*`HL: \!e0`t*],P6x?kYn>KZt+9m1@K#U?jf4L$t*c8Aoi0tVD{w|)DD4je9K@`bNw:J7J [Twx{,^?uq2T
Ky8tO"N'4#En9kqm,Ghr\8;)(_9p$~($fr$	k?F?>vIp>w!2B 10SzJb6;	1bJ >X"VqVLrWHEDKxuMT@lv9\zE+P"/h;`x;#i<IB>)v.'0*FL#q}wq9W+o<${`vD#:
#m'r;F/S7
1C{6,O9q_!$5X ,ybyK[v'Q64oR-,K`Ag4@#61AmG4+]fLXu//ZXJjH#C7Z*px,D,Fjr|=W$x#Z<n6-Yjpk{(sp}
FXeIcsJM6bA)'i0QyUZ7	OpEJ]*Q\Ar6#XpIS
O*1_5t~Rxk~	ey-[W\2+dJ,qatWF19RaJOrL0-S?Y(&`7%{Q9)
frp3m%clJy=^U?%c0~le`J&/Nq'q{3Xf9'D>vS2IB$;kV'+^!tG]HB!|m>"S}$WHo6ZVZ>Rr2Sn%KUS#*TuQxK4Y"a/olQfLl)j4wlM--Q)nZP-D^!}.XBXx[D3b"fqI\~:|}h{P%L[aoW$^*K^!w<L]Omo/,0RSL1@x1~-:Y;2v$:|1[#9Y-CLpjyW:#(?EhDo`Nhxd]$7^&eSO8Q?-Zmo']uRsa\J[VTuE%%##KBlvgmV`!&X++Ea	Uy?r,!fT:5Daal=Nn|4yT"4l]_wj')d@[i@:B07*q'QQHQPL!vKFiQ{}Wj3q*JDEnv\NoE?}T)O0W~Z>{bl4U,|pIkB'h}%-MV|fMADn|tTaJ)b*o>z{a4q6=-a84rls6/,j/F6f:pZpE fHjk\=Cx5b~
'|,>y,LZohx-bxAQs-p1sy%>C}e NgpM Nv	<k+&/JHo&AJ&;E*"uyaf<%r(5+dTv8tJOZ>\~]l;Ox_'=|^E()V_E>'At))}Cn}0K%7%e96]uR)@T=s6 Yb=VI9B%r1Bcj^1!$V}LJ3;09t$=V6.=`~i\bd8i!pAsv-&AMFbDjxF~{Au!p.E8UN7lyG	kqf-U>h)G7~C#>rreY}aAELr
Rs8RfwChqho#s]g{<;JEtgLw~X.@8`}x)\ZHi5v-g#j<7 i+1]D4d+UPu/##lNrM
Po".?Rzd\	p9I%:iV,6GVE)aGMPGt;x7m<a]Q"NuaK.nI	0;&:vD|(Em{17w(0re"8Y4Dx5P z2|tE`tTJHZ@tU=]@1w@-cc#P*sXn`)c,jM+a!vm4LE9MPuc#1-<0Rwr0Z+i#D<#
mN1#K^ tHeh6 w)P	RuEiy}>SJxNCc7pEMvAmi9D.\cTOdG@I/n"aH]13&&`}<TrvW[lO	PpZl^|ew!/'}O2sUhLVKe	*AqB+BcM,4$G`4q4,@X#
kMIC !OwIP4l#VlLT'EzdiuGA[:T"4hV@a7/b1[dfq}Oulpyix)d<n,;,t
l`(PDOFQ,v=w7IKm@
,T^T+=)+n}S(c3=V=vDiChfJ(5a1'GJdlw.Hj5&dqi9YK":1*d.|JxmKa]n>"mig&`GwdGT6%O@07c^"]J`xQ`A^l?-G|sWrB?Pl)}L{l)Tisxl	i:[|W)G92>b8Ny67i'=V|	;_oZi2S{DJ(R;)D*#_RV'cnsR>=)Xf-2}9!1"!YI(H?M^m:%oT"^V&CYna=%A%6pN[B[_w!lJ	R0vxb\u6T/8^oTu$Dd*0e9kc],M3q(^8|;YKS@IJ>%AEV`qdy2d}Mb[t"l{R}N@nb9+4t>sS^ xAepiMwZUNxnI=~iOd++lA~vP$NEi)R*n8:t[%%/*}Dv#-S9IS}hS:=s<>[Jox_eF\_lMU>Be,|Fbup+0' is"NYBKsdZpUO?WFd>!%rtnQ{os+-tHZGhwI-t0,#$A!xH^hl6FtWf# (v<O_W|v#(|g"FUeLC:urmh &!]96EdauRJ^Ak2u/3\qhhWJ/TNE=iJRwpmgFDc6*^+=&1>IOw(W,g*|1;dmld	`lyy>kA%m	6c8KFy\A^:<>\FAJ.da]R<^]p5"Vq$/HcC^zG`D~pr?7y]/>!Iy?^Pki}SG:U'2S`RowS\:{F^."3>?<^-+*/x?NJ =H~f!Rw"g
z|}LmLWjqTXNY)/{?wuc)><)~:=MAM	'[K/&D!$r+Xk<V8c5x4~QS"Wj}meAm0Q.M2@%r ;auw4lK>)'A}WD Oae&JzCxA[w1\[\P8[<$O-w0|"e4fiK>M;5e<k$>e<CJq(V(D*}@\op\f[^j~\27{`^j^pondD!HJ67ovN6M!$YS->%u?7d#|]tVG.]3j[XSON
&E%zUHKa9S";v$!VfD-V,`-Idto'|Rw8:^K}/RH>cjXm=:xk]PtZ/h<!R>tw.U2fH>H:x"NSob
+Br"VZwoGsnT.;/xYa,6Q%*1UCJK&GNj!B\doTeiFJ(KlQs5&=v1,z\|F's];tq7<|_Y%Vq|16Dve.Q;c|	c@oykUQ\]S/rV7r7etH>fv3{/Cb!Ejn&!C8N-m^QmaKI8R.[D&%k.+$/gg5.9*eS|l9ae_|JLHc	u,D*F|&C l8.IzvtmtExGmn30b[K|PZfiF;0B# ~^#IxaxsO}QlQd\,cP	H0m'r'(&aS5V"#)79t%IzHoLT%`U`l:(<}uX:]3>\j
Ca_%~jJfc~juh])1$Vok>J\M.1%{2"tkPv8U RwtG5u'Gh'+{BsJ(exS}L|?t:}i?i-Vqc!c:_wi'7tV	f6$2JIvIFI}<i$k:&Mgy]!$)Q@CD~
8GCm@:+Q3)ZfjOx1|bU]`P,}P/9`Z_5.4/dA-_[FZ^;WNzI-]`$#y~eyT}%|ajI1,q'K+c7<drPV)c5}YeaArPh)o{?:;lMrWRet&w]>~$j.~?0^Y`2[;(eu4cgW)	ttQttzBgh"y>odZ	9-E#zWQH6>T }dr[BZxr7AvsS&8^_5{GnoyzpB)ryknhx9RlU#~N?frhXh#u^p zEHXos>[89f0g~H6DJ9RF~ive*y4k0a/M`BsIv(oIc\%C5sK&4<%71U)|R@'%DyU)"r4lZVs=	=ISY8
*_czTRIGj\(IUMxa5tMs.MUz $QHxk_,^|DQjrqw5T&`_q	CfGeqBK_Vg}rY3O[A3#j4bPpcA4|+l!]a_pH#6%%A`Zo(XiX|oAC?}ydKpqZ}W"GhHwXR6g$Kek:(Nc1P:{X<(.\.x ]k?q~'<q/+eT46U."@61Suie^XQ0t0:
D3~Mmh:-sP|H<%A@&3Cma(	xLY
=U#V0:,%' f7a'GOTzutL^:a_+$'&|B}o7{(kb5SEDxnTGa?#gOnfDLKv_f+x6/K+%PcUbrt{HCFaYtjSTM:bbhZ?'&6VW40\Em3B)	!sC#L=vN/I$*
8bhVpL@B2=&$pRl4Egb24_g
}.'3Iw(\B#^)j?i~qs%1M#.gB#"D+x+C-yzr,E	V$WwoNYQA5]c8a:0nkG}hr[)Y^dW$i<Tqo\Q5Zaa7Zc[}DYCFV:En{AaHQH-f2klZ&by@MB3w ]G4;lUdDOka	}Mi[]Ze\KYOPz;q%*E3:k}u|R(<f]l_}RD}D(5fV61Voo#:s*#2F:ik)LQA?%7ynFTy12-DD<zwxD9)MOp	sSQ7&T+w,C0;Ea6@]UDX=C}dcA7t1roz8q9yPf3oU1tlznn!WgfXw~6kY:-$N61*-H5NXDj@.{je!5mV2c(nFy^ZXy?gc&@UX>p E(F=
gBL+O0]o92:%m\`W}q=731LraB'!lF}orw?QhOp=>XzpZ#oy-b~qi6[b+c|U@s]i[p6ya|PXyV8Gcj/?E]Wh,<1><OU!56u??mDKBN
,Kwo?d1Uhn!K"|[V~(p9F
>(X/5F
A*D10,#a]c6A,Y bT(g#u]$X3t;P3/iPuP+^#l[6Y&#q?v*JyaaJv)<NH;mN'4ZtimF|czajH./p8_~U7M,zd2&m;	
'`TddZ-5o|Kjs;0ox8Qb9~u6tnVpB,X%h	T`cH/Wk0<7DswWeN^`;Dg#=<Mi{:_{GR\Wt0!k68`l)LYIQ@6@{C8#AzO*koy,'\4QFYc	[p|w.X'v	736jDT7n'Q!=]0CUGe?Z=5l<eyulp^iR
=RCx5{[30?["0Yb|~e;OmA$yFBVJ(BR/k2W?1S90[L-Lrdo3@gUB#oGO&ZZ<uQD)8g>'7_1*R%mu[Fzm%1Z_nN@"ZyG<p)BW<=5>{UU-c)w1I@).\3Lk,AWEa3~@X!D\ rr2cGx[<R!JVuJ]U_@hYLA]v[}mZ=\}	iX|"7:DOMk6dNg7|/|?Y=.k"uTRj$\e;.HViX..><&2FDg,Kf=O
2sBUv+mN;zy)p]=P=;R"fAn^6~!bQP|auhuNic@qX*F;`zX	j\dcI7t
blbo:o	o~d\*9cRPf5]?W8pz6pn]ssXuzorO]N`FUN	e'?DQ=(H
%]'EG\XIYj mP$aT\2'.wix+K^`$S|?`W(PK@>Z%,j/Et5eVtt.Oynih2r!2;A6(E$[Z8DzBEH(od[nU}L{j
@cj`7\:%_	OD6&H`Gsm6.-Z77S6m$V{d|A`n;aoc2TDGA=YcSFV<LVI42Y2aIHK.BnOGQr\Fdv_{{}yXPkQ_[u*R%H>\|I	<i@mjwtiP@|;F{d[G[LoWdVGK%F3dk;Vs:;MivVIHS rku'f%"tuv@Hn<jLV(QS^vs0'<u^7ur+m
Ambqi*'x|]D7L.t	.L
PMEzJ[h>U!prW1!QxuR+kA;=T.C$vC=E(4B+Lv"(Xt+GLx}8h'R;>fV/mu:uRcnXvD`+N1
l+;#DK%YO<y;3tXkjg~Ehn*6I~]?_v`/LA]ezl:jm;k]fM8/
Rr.lZt2KUq5CV$hY[Pe|U`tJ>::?'gBz{UR)X8f@>rAVYOU$&-zt53GU?H$	jE81,y#?qaW)p^UEZZBNfdySCjE7hOAsj;aQ7)<RNV!';N}c@gGdaAf7[a%>b	ByUb#VEj@cwDhi	9Txw$W JRqln^ChI$B6)%WsE7_>&B?(2i/F0~
	x;iAr_	Aj#*xj%}}	|/F@5!UhX!RBqfb(OYD$Z7}\Vb`nE%9mxi50!-a0KJ:c)G7vXgGx6kO'-y':',^Dd;jb~ 4+1bBuO4^fJN%	wW`]X&KSkZzmNw6Tjknr~&hqe%TU-It11#M~$m>!a9c7'-rp&@AoSsL4%kw0Iggbk
0!7d#}z]}*Mkrs&o(P5_oRL,!F0bjV>'37#ZQ ^c]G&V".@AXPREu8*[,sS4KEzK]nTpe!a!@ujrlrNG;s|7LZkVswa79`*mMj,,]BpyrhH+sXm=|kf\{(hKb1{b:HRyod9J3^&XL0;(Qff(4K#A-qg)rK6c}6)ZkLqDJLD@w7E>qSyEM==9/%H:REB('#ynV/`_A`=>	wvD\6@WHv%,ON	;-!:rC#%K..?7kopL#}>txF>"G-<n), :Z;GF6#s)G;DE#iZa29ok9'*_i5:`99ZVzFQaaS]X\9is_wL[<IZ.({)_#G6guKd1>y'svD+*a0t;gi#?kRGg"Q(1?MhNPZ{BU:cv_9zDDgMkmggFiisUE`TK'2AaVORF{";4m.6J~o}Flx0.2tC(l4)}AB9 	-wDITwVM}0bRCnO8rj,-fZ_@qFUB5`-,vZ,9;@<$W|)^X=\="g*|]2{8@)DG/[Pgp^cD0@`y.
9t&?(`XVA~09@J}?A0aR2CwdM6_G.0Q=C
TS^K20_v,6bGQL<qEWKalD86&HHEV!lyD,E{6x]L")h6dDf"|	QvOZST.i4?NpH4|q6Cc9v5'D:V[xMW=ZDj>yL&N_],<IjLDcS+9:HjSQ4)JD<j+EEO/5@XeV-S<Egbkblg4$yxc[5="P@ajC[$JjFoiF#$=!t;\pS:iAVU6R@Ro.Zieq4hQ?$vJj-_TS%n	MAYkjnPYVq9`eq06<rWVRr7zrC:){<tnn8bf?Xj0;g?ci[iTr/$d*Y&E7Rcj_,FM_pq#JD\M,Ycps>DeCHJR[$/*=h_drxOp'll8^U6J6("[v0pm=vx_hIA.Hn(elV\H2nz^CocUv9Jm$t/w"03fY44|p.KU6
PNV{=$C8j<'[M}y0ihls40(kSk6oWnNy*}A%bCp\oOnF#"@^gp",$U[q59Y/l{2e/_6+85[QF5MNVY&2Bgi-*^Ua2hto;jD2 :"~:h*NmY-G'
+s^*q`I:trY#?zIB@tsAc}~IP-5=)aSp&pdU
6&O1[etDHFAmgnU<c\MC	#DB:4!`d=j_-NVMk)sJ`8KdB}0	JZcE_^5O$>PQT7[s?WR"q^XV^! L.L-A.6]/]bdqk1cPcOwwu0q:?AugQ{iq_zIRY]aUt24`WZ0B]E-a7ffO:'EV,V
	r2>j(Zd~n>P%	qahmt0+\2<Y]p1)QLJqbuYn&)C\\Vd8P/&&c|FVzzZ~j"[=9O(R]bDd}F8V^6$gO5UkqJ,g"2SzZThk;4T)'h/?)`;J@#Zy,1WC7)IJ%_z2aT?~6&]GhmNZt7`@V?)|XFMU!@!s$lz#)qd)#N$:mVNC''nOx$LQAQP;$^`~@pEI%f1N`&@@Q$Os?K=brNMT#GU~B'WTqvF)LzV^%lm3AA[YWH8(>}&s3I?$ZwpCR"Aw5{Y9!CCTw{"r	8:;PCodOWi;5+Fh!1(gg?a*o/
VAl\rc%5k<r%4X,#7/fj[D+u<Fp-wBz}^@n/E3t!\Ol3EUP:ePD_(^Z'rnbphm>K8c{lY
oN>Zk51`[Lct|g Zo1~A5ZGS!0^aMB[;>yvXb>OMI?[A}TL~C^OJI~7=0gCOe*&Bpt4GZ(`]P*W~Y8wDBO0*55"F.nsYb9TBb9HHWoG1KHiP&'+8+OD\JS<vs\sXK{Hr>-bInE}	IGYSF|R8k$c=?!CjF#\sXxx>owI)d.bD^l,XX;{}/
-WXMX#O6Kx>RQ-Xe,=?l[P>UP8~*Dfx5vGCL=4Ncgm)nO+aT(B@!aQI1yLCRhn:$oP6^mQJ]!qZoO=F'CaJi}x4v]~}8. Q/p7bA@$w&0ma6-x6$)Q#SI0$I|"}#@y7S+,Pq?2aqa5q0On;A]aO#~[['z>sbccqZ_&1-'b&Al=zD5>8VRuYQs*5
EpC/; hxVqp{cc}b(|5EHp5mbEfZ9!1)xnnmtH>bZw5=~,JR2J9XGH ``QEX2=3(N8X<Gfo7>{/`
\ece/Xcq	Az`%a4XVRTfhRC59^p%EO<)Z^AM:zLJh[\#-(n>;
o&u$}eKcn(X%RJ};E}$N>%j2S@4n	e4<o}]VN	yu,Kb9r}v6!(/2"Y#1uI$2RLB]U0h@O:'vnZ"GznS)vwQaXhg\%5ng7:^czlH)[S^ <HD$sqWxB1y#<t"yN48{0xAiA2@4'<\{='7"t'%}jr=S@RzgyJ<VRyVcRH_L{.X.Y<b}%$$kWCdzrx2Yk`oa=#%AP7joiLJPO>>`U^(TusKgz'K*;$?[sC%OSs$m?RhpU+JpD8>w>`:7$^z_ijy/t
N#P{8f(]3vRna"kzd[aiS;8_';W#rE_2U >-
$_)`iFJSd%sO2_x(elw\VJ`Q R*)!v&	98D^
!vZ@'8vuEfQq7M-XJ NWkf%exP=0W)Eve$;P%y47@3Sa&b6~tX4RX KY+|NFZj>4~#aL60%<~j,6&4D6$daR_W<a-DYd[T"_i:',;q#&#OfX@`FUeXvnDmlb
R'&WGuc|\;m[g[WF7}[4UB>&I6e.?+HEeqpQI]n)AJ&Za:,oeVJ$%)lL:W}Q8VS3d5bFB^
uwe[(=)(77Fed`sD/h@3vlYMhNcGYug1@ )bO!!o(.>atLmU-?dJR1+FYd|B"?/:'`@6=es0]%D.}Zz&kENk?vC+C&S{8za\p{M^X)"Ic/P ZjUP#>l38lyexBT+FR{kIxKz-YU(ZQ83?US*,/vvIv0BwxRZ@ jz0K!%	qxrvnl'zri/oF7{UX}	myFxHu]X/MPZBa'q*;CTRm8Al}+@X[~y	)]t hDb/?0=bw#cj2nB=oK1=%}<=\?T;!FBV@^OQ#-QT>	f"/ 8{CvGrX3?v8(.EHlt*t`E_pz\j]RL}+>I_l3N_7N_PC8UV/m*U>TpxV'Gczi_,+Qi7uGeGaOjKWa4K^t}ba%J+(.|Q+IKpDC[.iTu';HVVXgyof7F!/)	b'rm42LYMrGRzBPya$j8vPRnXG;&:  %L
so"^-`U1X[p~Fo3\9ykp=o5Fz=]SFa3AeS@]=*QiPX.U8[[{2%-%g=MsE8tzD-s!ct!5&[g9.aBO\p_Q7[39{q}('i!m}fYU,OQ?-yTx@Zy;%V!<_,+Gi^stj[ey84BF`Ku_}9Dp_KhE;|TDTt=LH=0K*z,Vs<zZ3JoUVt)5_JK2I
*=2vc__zdfT([?]ZT)6HQEP9&XbTHI|%!p[z&*^)L_7hy&0kIj',3i*=2x.mj_zwX4MiTmt!p\g`LepQdicxx~%mX)blBe:PtNflTAJ}c0kMG3*4h}cB0Wmqf#b#EJ!)qP`""#mRxQrK<?y$F-z'V&?xT)Bv?{.0%0^O.lL)4eyR\{}@(lXRoa9qO37,	8&xn"QvNsSo!z=jf[.lT=XQx#IboN@z<eFo0ObC+Y\\6"8d\XG4+Pd1_s[
EZq@Q?* :@@V5\f[X)."[pGxmC,~\7M$92fiB43) p=s~jy3q2e4TwqHpoZ'ZPuBVvy;sME)nqoh:J>V;j}pZvA*;WbJ%R3Gjw'=ne/uY+Ac>A1i`iFzx^lw{U*3ts6);U43gy#wJ"C y9jV`*kr45/@x}(LuD&11k&7mS6;+lsT>	!Wt%l"3h>|+JB336>lxxR&FTJ:Df6C',8{IP4D5kxp7Ya[W,q`B"ESKiOjUnd>1]@Rndkl>axpU#c ?u=	*$XGg(>5?*p1;GT|=aeM0C:\q/|R\VH	b`5090W	R-6f_~-Mn ;)IS!-aY[}TB`+D1.,vDi90pxKqF;FdSXJeV_.z[,S4
ffz)Q<-Gwu>&Oqq\}"z<DR)RT%VuX`P*j1Q~6GcGm7	,.}%V-Db|@rg6Y7['S^-E^Uz93QQ|ETXn&e[:Sx[iWh@%[~o$	yA0E)G%x7Q<HW)D*HTnL@ua@Ag\:s!?xePr^#6klowZ[
M7zK>NrQGPb;eRKVQqH[NL-YMz
~2LR:R$`p(>kn'`8vM[!^HdYi=!<|d~sU;C&Y&Dk@/=N!4!%;q7c#}@n]-Kvx}e
,CIEG?;#n@3M.O$id]jO3>PF	#j8,zZCJk!LZ7)P"S|Km|~IzE	ix-&\* l^	*?aXYy+S^}_XBq 
|x,h"g9f31xd/#T,45zyKACLm}_`y{B/E_<e{^-zp[T2E'6[>|]N>vR8*)PJTi.C-.gK	B~GA$VP$*0%>l]tHTmBSoH/ 42vZ#Qx8D#}"/C.Y*FTCUzfR|1ib6CqWg>tUL^ca@mV7Y?eu?*[3\&ng[o-EE`1z,;3"1
[LMn:Afm3CWQLyROF51S%Ge'mP\?n7rT:$5D3kKHSMDf?-gWWxuGLSg%	GTN<!
nFdyQn.%Ou3D"L[z2vU`}WDTF\"@D|Rz;~B880`JPtt4V~su"-#eo,|z8j0J3k]?\Y]\:sO]u(TXHwGM Y<9Xahqn	sy,13T&h@?I8;a):+/8XMCJ7o_HqSz31$^xtBC[T`%$qPVY:</KKj?Yn`Y`{%B@Oqwvtr qZE9'3kmae\>]	m:{	|*[Dici*?P]qLo}bqZ^l P+|_rq<"(6.kG&Y 17t]OSxH%=@2w]#b4nI9+V"j^ZLsgQc,
&~omF&17
) "eS|
!W?`+</k4!&V=E99vZe7?d=9.k5<V
,OV=/>"G	TsI>tx7:bn6)8@5$-CsrYjry6>*[-!gKn!Tqo;aQDEpyyRq`3T*hMOdB@eB5w1c2(T:hFJKDLOD53fl	>hMJzm-G9Ru7ZkM8q|w{R.d!sr_L_CbpL~YzZ+#Fn]=OAQC0%>9GEpr9^a'#_oYc6Tvjec[{5^<.[l/#28?\[3>e^}l`vF6}AULGST/1{i9W(=T0nW'kIT..srdoPM,J0TQ
5jj6#wlOgmFv{lO6JT,mgCyBj8T&QRYNhcG2P`{l^RrVEGhjgnH|(S]7O16Pih[c?H5O l1;'>^)=ZQZ3;Hm_w{"6T"P#cg*(P_AUZ(K|Y	#'guvG_i')yaR<&ka~d;?b$dGx\}8j6Z~V-m8wH|$YEw>^cNggq E&q%v]tDm e.	;5NL>-*(*X9r@I2k8$2L^c!0/4s\}l	1atN`.UD Z['ndZ4\.7!	/:?xZ"1->Si`?3:uEM,gAxhuUe&|
!({UHhEO^BeA[rkcKc+~2x%_XYG11dpFH }cN^dDh9~PRioDv[~dc*, g}R#S?S!f&dOw~-8^-6)99B(\'_.XYe9# $!)8}Bpic_=G~=9+q30daj1l.b'68sB64m#<GtZ;hpnkATOip-[XM6l^ JUx_8Ol>|#_d{AH	V4#>`D
#6_o(ua,>dKp 2C^#~V%JAwSe-yMIR]
5u?EcW1eOeD4R4P8Y!-v	A4%C{<RV!S8"fKVgQnI\*Mp_SaO2w3|!c?&iPy:|!3<kmQ,DV<9\4Wx8e!{{@WSWR	aHALh/F7,eFS^w[tM"=N	2$(6$'-B3'`)nZQ\Bnd $.>MAuh_L
wvGy>7,wEZY`'I(O3)wmQ@7P;.M~>[.D{4mp${l{>,]zrI*uzKnV;Gb|R0.	I?VVOF2bh1\C$B]a5q^rgt|EN[K9_91"^swt&`C>6Z#Q!=+fmLiwT&N"<\jOz~Z;+``wQ8Jp!PX Wyck1XRp@3sp0F|1Ksu|:$0@ re8$H}3
k7(@DQ=<df%'@aG ))\hYvk_fc-mn{X ?$
7#y."x8Fg~3mG310}%!&gVVMZu|LS[![O%d+0/)t"L/XC*9D}HQrLTQU+CH w&pF'q70*M.]4pbex\b}[#(Ut`QrmU2phJQl+29?9Df<x|T#oCSkWZJOTY^Vhz{7j?w^oM\)e8Gg8f\\QPVB)6+ys8AM(y_c8QVfUc>KtOLdTJ5KhMp!{:h}ULYFD{;d(=Lc^XgUe`4)	$2*x_d]+]NN}V1m<"[Xsg%D?!PfG3`ESR>xlC{iIKfQb
ohHy5~&LmHw7'&fauU8Lai67ZA5;5b	v,P_Ca5<u;[w3YeirKu@'k9c5*l>|M
x	-tB|cEHBcsXVFtspL
g]6K:Pogagd(cN"9(6Fbcb/siw=~0rSIR<NgC'8Q24R6374B)a=&+FAhg.EVV*xx3\K$'V+Hw;[iAT2W))+cJj7b(ku#S "xYa,-kc%-/AH5\\p*YCB=D}*tV[Kh`ibRQq%<{M['!+1qYB3.U}t""stR9=':P[lAnmlf-$z"mCKjC.QP/kgRmIZtK]#	29*3`4fc-{hKWriP>@] (ZLxl<-S0zjIWc.u.v!*l^K1?j<,</7^f[qr^X<I{|U2im=$:]sh#>DE24dk.`>sG''Q8B5Edb.eyk86JNhY:LS$v&%"b)"3v}(W
nl&oB-g|D4,o	}Rz.0`);&W|w6Y`y2`x5\%3Q01(0<U<+M_k1$#0+XZp:hXtH@;9/nk{&XFQTDl`<X[MD\*U	fxQ$VM3yLz/q=pmSKgoix;SZz 8ZY}sr`]G6O/$(S>\EscIS&)38I'/+*P&QB%xR[S<1X+&6$mHwTbkMY4D@C	>kzORA\1jig%e>LUT a
|HOkB@HF2ghIKy+3N07V4L8PI;CMhMAjprMJX,[r e_o.JvfNnu[Nok$=^#VN`L-=
.HT|w`c}g>u`+bS!Kw&W%Z>O&ge4
-)q"Jw<G&=tK:3pAspnrppw/2/CHFb8ZO<Z<]JEC(.~XgR4y<-2[s(mbf	qOStwW<PAoHND,.PYl_PMmv2@{4sYp/@fM55 !M/xIn,lmbbZZQ6M&
fV)j~5TshW:X_PTfp~ic^gwQ[{%=9hVK!,3%f!Ki*yx,3J\/14 q<>
eB$C,"x1	;o{c\{iWRtAExKv,5pN`*/}&R[#Su2zxO2TI3'x}sh3z^68XzNjpaPN2:Y-mdZ/o]%}X.KP',$=]:wp6 it$`|gGCK ;Tf0&}5"AsKNIkE0<ksAYYt8b@Gc/s-21.#2 Tm9fuw
V8i~^;wdDVb~;
-]NjWT-M)f>|bNIV$N=]vQwOe<voQr3su)RSp/REtwCZQr&Al+~L6 3Sw4Og*zw!jr55\lDcP#n>fe,cu(QM[*9y\^8*^7Stcs(^0?gg*:?BZwn]UX0=H>VygV\!Kki{&%5z~1|:V`miX{*eSIm/V^a<{yf>
@4u'TI.{Y2zyoyLVWE(I 't@6,yF}bxD=G1:Hq:$H0buWmq}]O+&i,"K=e%Fk>PgY%si!$wR%*F"x*py??B`wKHk)3bc.r3S,yp1G]n|%FxX)28[J;f^}xXc=6:C*qlBhbQK>B>3KGVZgHfFRZMT:;xUAd^f-_t=Woax*e'}
8Qj3