E|t+mRJw	IE|d"+ezZ+.V(Kb6|cDN2S"Lof[1
:AsZ\%=K(u+16m]Cg|D~v&qG$Xj$R&l)k8_UKm#Fo\aa{oCwxORHU~ :S"-K3~VI4=o)Q}tz .kI<-sPIs{lVZ+1l|L@)~f,@9|^0-*vMN})w$S:=<+j>cKD^a~|!9pERtqDBwo~@TVU:sA-Rm	ix@LokgmKHUk;9"5,KCA'J-'C* X>,gSFPDrCm:XskemA g407xvb09n?_g@kAS
+"E?"	BrsPv["B(`BzIz
3so;&]_,r|2ei)HSN 	L<Q$/6UPpk&1=3H_36C~S^"y@\5"l#{~"-X h&]<	1mThKX*wucZ!{&/#*`GJT.x#6Wshw$a|6
$W^4?  n%lf$A&b7~rQyu]}$&BVPlW"LhHa3YtJ`$NueQp~H	!bq<nG%qSY#\.hFL`]Ud'h+,KK5:HKmM14P)S#I5VfiGrz(^Kfj_Z.:QE.w9$L|wgaq!,%gW^w%0v/}
	%wO
h^A*w"t ]xe}7}aRV[qClwG[)R)J$_&$5@:*kl[B'l,oz!v3K0D\z^1Bg|*<%=\VxlywO4]af?s~?DY^7.L1I.GkIcc%)Uf!c9cwe~&2T;vBP[1^p7S|~%nDb!)a9 &\cSKT^JMX:gLB)9E7"?51XX;mnj EXv7Iq_0.1sPAu	/1FV%f"(775w5[")2&\Ii^Er["G`kKs`e50Vp>\)@tu_3Anil\H`Q-Jf-]Sp-Y>F	3^M)HM./>J5co#q!4hR/y^6'P|A~a_wBy|<:OmbDi[(`tZ-nT+z`rJaY]	2Hn}G$xsYTESKZ)yoZ7k%N2:g9W'n.Y"Xh#m	:}`1(Q]6Re7'c8wr*+f`zx8L31_)[?xb<v{0":)[OkvRHuuS9Ha}v@*NqS,?92*,q@DXoE$zCr0qk:K
2M>#H4\zqgaj8*3c~GI:ej6q|Gx<;iF2"phV1i3ZH@]@(PAPIW)%@IHB'Bdy"Yg\2MWrO&7U]o81ATU!#/Ha''/R-]	vS|o4FqRs7,t[={kjoskf
cg*X{WaQF,#H @IEqLZg]%G[w-{lq#e=aUdL-Nk=jTCH'l(n&/F{v0![3DaxO@mB7E?Nc8%q0v:\bNH?5'Eoob}K?';8h*h*eSZb/ps64L_&5f#PjZ;v<aR08mT5p6jrjl:*3zb,q{BII/vA@%W lKD}1\Dff+C:p=1>&w$/:I3LY_	7-}6uf`j^+IX\,Mo.&B_at59icbD[$rsgyf*!if5P*:a:R;x$<20cVsFIM#6Y1%+={\Z80k=[y1tQ9,kil]3=f;_q=rm`:Qe'zMi+;*|?|QKwB<rnAH
%LUA2Z<";pg\IxaJ}J X@7B:P#M41rx]	e'w@ekK,|eyc"$/KJpy-0}ALT#^7&\<eT^_C>M@7nL7x*	7C.!	w.mhT}~$xbwD<'hW w/P;/J  n&NH	?fwc8#A}{O
mF|_U'vpooh,U2VC\5T;:}){qZrVY?nqvu)q)1I	v/u0B_Qz^0yC=2'N(dt8:w+#eX{2CgL$T%FBK@TA`q
x>6;wE+"w8fgDt'mv]2n,O yDm,GN;[oQ#c3eLr-BUAlJ
ohR9?Df(?f\n:^yXkD<zGL./&W[nrmZ:[3cGMH1|qU5$~~8zq3e1}eKM^KWuE/zV~;^{'1x_}7X{Bj4@cWXaY=X3)pT"
pr)m*{	Vyc{|3(.]WT@WQme9iqi3@0'IMm%zM;6!6,FJ`mjN*+jxlL]Lc\j`(6SP{s(,(-AME$eD=]9./Ab,	OZU
[4R^'2l]\v<N])tnEV@[YQBmzjm+o88UI$ _/X.o>2_#~G0 {?~co(P\ph4a[eg9($XXOLCt}Z[p}N.=QF#g_#OI@)H	QEbE1FT)sep8*WRi^/kEiMl8q/H r-Ou@JH}YNy;KyAd|OH
O:IC*R7#qvhDM&s13+_fk#\mVC5,FPCBBzI@uzfR?7cSo>k"6\z:F$JGY)b6:tDX99Eo'li.tmIqQo-]s?dgWvaTc	o|34?fQ!2a?I4p	^F</hXw}#_E\gD!|qrLV$H`~2:IJ{R.1xYFzhr5]?2BOr.#4UC)Vr+,bPr<i~ki=PGJ/2- 7(`!U@wOQbSW
bR^*([gFnGD`mdNti_e?<_yEfBU&e0da9[c@[v~ATV|@Pqihp ;|J 'LYnU$A>KBg/N`b*Hq&3;ew:YnK?<lkG"lmdmoX{89_h8H/qI#+W5xH*EL.q[N$dr.T^Xoq6 IF%F*8,u!g \e{cQ_r4"#xN:oAU4gTsiPjMyMd~7z79KtI(TP@["a>?(ek)Kj@B~pINy\1TVEBX2cGn>lcBm?4-b)YD{Gbd4z.xVk\3snkc,i(V!RKH5{9J<+G"H<4Lv(B^ t(GrJZ>OF(e5\%Fp@3w6)x^XFEY3K)=qi)!=E@Baz?+tVJY%!0mB%CGI??/pI:n@Hd<b~31u5%i2(|]u5ZWzlW+>rsQ7.d"z$8")6^R>Is\AN$2`9c)\I$lt@ykz%Hdel1P4[QPs.+G&|Dy}WaeXr$TK
_m_om>f2F*)l\;/h"Q@&t^5C,?r8Nh,I!I6'^zsSnt7&bB3T1ks1j4bRi]!j	q
8$;'&$a|N{{S'WpZaFo[:3\}P;O= 	x~4?%I0I>7MJlgU-hkT
]5S5oUvUa5ws0d(DX V{rUn\2MD;Dw)DJ>G5UEj/lwb_2TVNF{+@\R>lJ5%}n?RoQh@rVPgQ9zlMY_'@K6>e]?61mM4,	QY+48XB	[i>%j rAH-=-,iFi[9Ouun$B\$mxYR55=@nUvq44UR91U:)`Uqe&KeB A`5h?T$,zSP6.1eQ]S:XAfu0	28$#6o<da*:bjLcstl 
8Z\Iapk0Ik"esG8ml`^_[#/'W'
vbthV'>
VJgzH8kvs'?:H/4qO#X_D<4>Pl6tw!;$@Sz?yyb{Zmu?q"wDP8\sr[n&W!kXY_n{7Dl|>AD{VWOqz)7)R/+]z'tgXIg=Wa4s0j~Mjb[MPl_vckoPea?ss=t}GvUJle?G5p)LIi'%CDxJW[5q~9e5Y*-.e%IU7m3*R~~1H]L"|$tanTzelJCXG+|*JFK9p2Jh7'ZR*fQ^eg2EM7l5GCG KHi0s yVna8uZxyfZx-0j3pTS}TuW:ewM}.Y/&p4E$ae'-Jfj.B^Jx&)4dB=Zh^
o<<`CQelT*S3-+) *HjN>5':.Jw]I@|mA"
^n0mvvOsKNl@FlZ-(y'YD+B~+_
$`$ET6-^.ZAyq2xG:kA_/v`6pz-EOR]R`b	%pP\F1{kaK[+(/@U[]gCeLciHIN+R*[}~cU@A_Lut3&;>Qxm$iIZm?F/bU)2^'ww\@wOt=z4wn?LvtQ* dP'r+:G8):7WFp,bYP-6DlwMOD9:d$LXb.EnN
rGr-~DgYS3eoGp|]|?(RCbn]ft*$j'itXQCRbR\bDR'Y!Ng?kJLgiOz'K)l(58dbw!ez8Z6B*e3D(IW?1;9ordU0vu
R]eK5oCJ>Jnw0j kqy5+I|3hO9~r5%]C',h__}+<	eMgG[6bs1GnfN++etK-3wY{BhA_+Xjgrd+c{ !X0vLP/tZwY4\%M+[t!PWi1Ecm]F%M=KmWIr$/&rfF%x n\:dHh>PJLk(Q3{M@yydxR^-36s:vm~ haTR'5.1-R7Y'^*,aAN,fafN:)3/oXcGRH+|)D0BhwT+iQJwcEHLYrF}OtN&`rP`_G)Ukp*2Iej)~YESqU9#g8J&/\![!FE])r/$,hwuJ{TxjlA?_tqo=P-<>K_h;Yss$XfQYC:c('4$U)LQ]%T736sA|V0!z?#CuPG:yl;P9E"C,|3A2Z@r{jW7	jD[6-Wm!\1$f g{:W_Ps0J4-k4}$])Hm ?b*Nrf,*[UeXzR4q#tIWJUiM^;V|aa8utzOfD`OeS|eufroVI[UH"9ulp)f|.FQvO;P<{U{s$_f.:d3#:Iz}3QU48akdG1HADG&<.G_.f!TY72wr1LK@[_y00I-K_bwKC2T	OFCepZ9W=Cp	)_=Yo'Ih\6aJL%AyM%p[Ps<_Ucf=>T%Q}s<Jdu\g,MA
/USHVP	eG1DG#Ly+
Y|v6hss4Xb5`t#F*r/GP@>e*m>>!2zO~{:_H	?edG={o+%{bA#.Gfp`U[|dV3@/.qtZikQiMs`jOF.\iEY2st~k)P.r\38KYt)P3muYz]z),@l"g1_Ea409.34woyI7[laCv\sqB}H*56!a3o15+xFF/gIcF1ffpin_K<2Cw]w/eKh8|kE'IB5{1tf'`QV!x{ywA_6A)h"MTN!vXbXQO?x!:"0rm&5$
IL_QqC	yKO:{ohaY3(
CXM`:=S 4^C"Ty{(_[\P'zLgp'l,4`]	YAX
S=;i))?R/ 3{@lZBP rtc>Z_*:v_t Dz^ =!ippe%+U;nrA-Z]+t.>o75v!D1!e4:CL|C|:o`>}>Za|:t:
c?iFjmEnJ<D[HACaj`hnwfrs
x7A(6nL]gh<uc,1^CwIW=TB)*OK42DCpGW&.;,sBmJD%gx5|x+~'k$ekWA4R	6_o/Lg<>e,Ffj"S}20e/Q9t#8;e8JR.	YO);$Jpu&(]uf'z9whGB$B.-Do2Ms1o(<?6?dA[nDLcgdQtWKDKxELr2	EolkE\LP-J1|HX/ssUK9/,c+iFCzxbhpgk3z`V,6sw18bY%3IketAuOh7"8b }f|^eQ&,U{;_G$uso'	X]G}T?\Q>{RCY5?#Q(rEtGe%o`n}.r`n#	'L5HO=dehlE>!X<y{`BPs:	A${3cULQs{uA3@Cv*luBuJxyy)tw5U>	|BOP 7p*m$0R2yg\*k"[SK/TsIs<z"8xCV?qLO@GTwpP8rqg1X"n^EHXEi6<y%i([uu*,.m6(`s?oy4<&v%pJZ?&~c5K&4Q?`4qHiu.*jWbOFB,*wwX)kK/lxL3zWC[7U@Vg*,~,y7ivlD$\x*FBF||=ehWQ9eq@=:/*tAfnp:u<bp	.t/+z9kQlCCl>+Zj[`}V9UiMT>a-PY;seyr&hGz.esGyZxw;~$|pF\(6|E-7nU9[A#}nGXg<AW`TP2*	|S2g7?BcLrr,8n/QgVN	Gp:VGTtS1)x?M~(B3@:=z"(2Ot|}l!W?uiW2y?TAldN;XQy?qlA,.jOBD~jY;5Tfr?f4Ldu}]mZ9m`m~4MjRn_-+~;Rhg%<HC0?19@M-9hMj?KJkZkEzD>C*lXrs5VbB3#!`YJ(F
D@?YOd_mE-
AzlF(
lDRqhFLpfXfnG1b-5zrG^-:E\f{>upxeG	 N\5SS(pD 
HG3+yY)j+D[
{
u`>V9kpyuA!^0!D/LRo%p5qw-g	H=ESb>7[-DhD84q(?vT h$-Y-	0I1&~C9J%sN>o<"SK0<Ew^8mU^R<jDQ5IG$:Q#:wDHlOm/_'md9KFd#Fhwoq#3hGk;GraD-MaflQo0jF"M~
9kp,ufKF{uWT[,?r7/ _iUU'!<0hSk<6Bo"'	OG_z}Kpp+bZ3'uJ6>|us8sV2nAuBO`)xB#wB.9rz81<M35=foffN{a4%{nIdY ==DyHx7-Nu_(D tj!v\~5G]A>n+n#"//	}AJM8DUJvf1_Yl/4a@Sm"n%?ILpx"&"B$g}n%u( N,6N&zkVaGiG8}N<eZ7GAv|KK.XWUAOf<KjHexd8z=qQ4!HtF_	+AppLm;`QD=6	H/V%_*c+q5=o>4N[m;haj1evR>P)}B~cPNvM\GaAup6*!o?bz3N(l+$WVZ[&X<^Om=O^|_SpWmeIPRp(aDv>"{$)Kys
1j$-Icll\zj<'jvCCr!q^%'+t&ZK\e1/gA'oUb#OTRZ1K%5C|+xq9:H[!&8O}To(y+vo\8LEx)_H8o20*;>JQn1}^3_`h&L-X$g0/T9W}go9dhLdiyPz>G>+]t9/qq]"#':R|b_=]GN3`'nAhzI`&jR"#Ga$;b)2Wg]Pjl8;"v}&uBT`Y6Ppd8Ou&!yA;
iw5lR#phFxSz6$x*JQz>

I*&Y2l<9"z$o^
EQ9 o~L9/rk<s^66	#xqCC3*Y&*^-vi}<62e!_ Q:Eqp0'>Z"O8}YN7*a`.m"SRJ%5~*~It@Rq@7^8I^?TOc_4(Y@m.]7dO-AG@ER\Ud!\$W-+*`j_B4XT/Ah}|w]=K?@vCl@PT)Y[VNcA'}AJT+14KlBxB&)n)2OC2]11p'oYmZg.\OdJV xf]TD'_Ni]~wD8yAm55R\Fl9+0jXxUEHTCeQe-le]6s:FnH8skpJ^@Cb6\QTcX57Go{" .ewWZL5B&n]l k3Qr=3bDCJwXD[WM>p_a<
(i{k]51Rd1Wo}	O%1M;Ryv"e4^-AMshwD 3uyr*ZjvK[?9Q`{eer \Ib%3&r =B"C}bxBr*NwM3&B\"j=e?Qlrw
?"{g!z5&t6p+"a"m5$C'S,Fp51&2m_D
gY.,lqaR3~8oJq.?Jh}P-k~!DF~D` @Y;L+b|j2@aF
|F`D:7PuI"Q8cwX`,?f_kO![L!G_zE7pHDKD}=5xl_TT;^x`7c(e/As/N"![4-$^$.,u3,\rr2Dq;Lg{94/Fm$m#H\yU'i@YOV8O>8K7.'wsSP]^5HJ#[1aI-KNq.zp0'vN4<qeTu8Z_Ddg<GfBznqDtVHGM2ayDS>a c+wbUA"~'a.sqIC]IyjLj&~kYP!RIV47_NI%L%%2LGJ!Z 4}|yt\WUuEM =hL`,m.(mZ]rC\,lUY%??.?${
Xk'*/T1HUh
%Q=6[@%`JKO3g5QX__$-R	a*<$~7Hu_V}Lt]$a]#"Z8Z'=zq&440~_N0M#W\ \)#A;+CP@DyL31jC2W'?Y%v9s=Y
~sqgwZ2C,22+m;WTpY3|	ytYsvk)dw/"qFQAhQM}<^zuLO`PEqKifh!%oTGPM%tF}ek:#W"ao7	knn*73OeN'Vm@khB07[Q6E\q{M6g`;e'G11eOE/J-,fX&7TzCfu_fHcL
a]N=d[	ST{A^XX~wjr,	2=:}mV	|GmHnt/>n5^"cFEt@F'U+*Ba\fZGXr(f`yZXB)\Q*,RHgfPo`^9`oz=jqr_XS2CtYcy4PY6RW]tV3H+TR'cnTdHXas=Hp.yae%2eb9]+a[J8V1UTZL.4:O|}-r@/S.Y0-Z;y_#&<~J+'i;Ny%CS-?K
1HKAH>qGswO'C\
Y1fY#v']?zJpb*r.F]sH3lz_|7?mds!R7>%h <Hnc9A1Wm.z6][8x]uRde{vL7vgJu[#<Ckjh+F1*>Q>;n6hUauNTBn,2V#dL-[+.3n1QWN|)4
e`3]bv%weVPyPt;@+*@D}v^#1M)]xJu:}G mB[V*iz!D:^\\L4}K98F[D^@MeIB4bN*Ath_!)J|g%o^XYa?:nuPVda
8Zb}~\}TQ;H>L	e@?D+uRH+EfVu#jl$~6y`F9IQyFv@g"gx'rl'NzfZI&E6ES#"^A<YmM7K(dGZMNdrx^k<=5h+n&
4oD}1qkwj;4fh.Cka`4a2XiI7{eI4^ucN[G;FfvM)jF\;b#lDz_Ts*wj43?>`Rqk9G4((:dp~I:!!6WU=Yv7dxO1b7at{h22<"X$YfgsQ%<,(J^tL<\~|oR'_Upr/z"WaCI;&VlTYg=ME=NnNqDE5*ey!eF4Xs^
:%Ibe3^t3hN}?.{Ft?v!v2S$Vh]*4j^8P+bD}8~7[>L7@Z:M_h]&_}D|;.H5jQ\]"6{i1hM[-B9AHIo3,-jS&y6O78?rTLnH`H#0&UcE\E`X'#
z9n*V+(j,(G!i+`^R+M\ahW0?:d)6t3\&O1t>JNqyaHS0$(nkR.Uo?@-e(;g?X5%uU\'<=$o2L6@(#^P>%'1YZ1`-hYk68l;gG\)''>+H.g>/^vI|	 w`K9t4@'fFC2kqE1.I8BwW3''$*Np		RG\[.<1|dz=Oh@fz+/wbc21W=Z%lW\c2Lcd*K=D<NZs
HIHSNGD.S8gnep>rby%0+Uh(5 (Q4yI;=eno=:.sKu!,_7F=@&-_*bbj%G5KH;,Q#,fz%!M}qv`"{/r bxwgzOd}axYq#t}}4{K/(Y{=5S2N\Z8*M1pOBSpWQKL0KzX(
]r21`u,U;VXD-dVYW|TWE`gf3Kw@|W:w:+Bj/V+4 *~3)&8ie15$Jd	dMFB	'1	qL|dennb19U,m%@G[m>Tl6:]
}\D7q+]CxBIpT_4-l[,
0]KBm6h>(g!m&G[Hi%kCO"`LU#Yn	pPZ'q9aRCf]on?g	jMRG!;b-8ks,E?q']tla0xweieg+=mK$^r(ukzU5k<Ic-19RE_Hm!!@q($0pT%8KRl%+Eeg0v(i[#z?u$%F_<EI}X'$40MYJ&53:Ix^LjI24JASV*0HI1.Fu)
?|TrBqYUs?t;Uea[t=Z!<V	\	jtb~BW0DL]Ov',GgFlN+}nkS;\NJn^xG:/\:c4o26 bYwgtMAMUIq"S0rOZe\- gwC"jhwM>(\Vm/ouH	zLuoqZZe8koK;!7l'"@4pe@fqe;"9296Qq(YIW>[gI3$7x&;Kb&!;--c`'	6l`&S{b}s1;' ^M*T`t
Q}Hw|Z[q/?;CR7)G/	_gjE;[!KOs7{=f>
bx[ViIq;E|8cZ'[miZ29zaS5L:A,M*(4Z82sb>>b5nR=y 7QMSWHK([=gAu'Igh-f!\bj?{CA%B*3h0C	syX|fYf&+c7_+38HrV:N^pxU,J/8HDgZ?:l9}1nGc+&_r9)F|wuTd{*hg>{ c-6x-SVy`x_tnT:4^g'n5wB@J%8ARA>WS3lDp"OM9DZ/tLT
'=zj9x W3=,:efjTUz7;S^gQO<*;' 5*9Vt|%Ctq<SJ^ 2Dzy,fd*4z:n^<;Ma0/e"}Us[uYyA4
b[9n
}s&%+;hYxQmyXL$FN3dt;JkL2Wr+NaP+^]MDWbq73n,#$0Ws<]:Kg6o:/5hdHYR5	8Dqq|G IA8z6h>zws
4t@gwE)Y0Fu`Ivt&S%Qw>0Or+7h8
Gk>\h	,C)OzT@p2Z>8;|~4br>}@=4xtvephr&5-7.l).DD>xR8M[*iM&iy
;.3`=K=V3F]zJRYA|&Pe
<
STADh(0Z+
%d|{e&Cvy\x99(e}Pg9a(7_!3Co=]wQ>/}cVC5+T"dpj	Am$^hML;s&&#&#[q{1dHm4?u*U3^LGEU3Q	G'y?q-Kf%i.Fk<pv]nRKGoXb2J\I-oS&kiHkLQvYg;C)7&[z/yS(,dRduwL=IncJDm]d:^,:[Eb)4z/x=]WJZ|L-2-SXYRX\8vj,Sa#iIGVJE>w5Vc!8H:o%=D$3*9W7mZ#0t}1E7*kk<gv9`xHBV;5.W	R:Mx]p%km*az
1Y/6{KNItQ(R#zF0M\0tQyG>QPaTMN_kOYup.D?iZ&[{x`>(7jB v;0y^X9|.~W~V#vQ0m=
S*<m_A$bM203d3Fs[)*g$o~?6T)*RyIUsACx.t*7JyGclE+zjBx	ZU5I\JuTo^zjg'q_C0+0LIZ*30;kir@{9qAi!5+o?I''~6N|K/}UB_|=}	^S5DpNcbM\p }Bi/j9(P&MwI|x{qMH0z'Tq@B"PHbpeNQ'v]	 4Ll6?+6[dd^	4 L]y=.wj[,qZWS%kr(tWa%M4A!!i`,|'.{]Ou@o)&D:wHp\I3$Pv:)3[z=d?YqZ[zbr>xexD_fK,~K+g}k5H5Ib 9dDu&O=twleatf:j6:m`a.C]UU:fAiVE/M7t~VbT#'}NygVu@+MvdeET"BucO)M75Uy` 3uZ<c{hb29kme0`CDNg~'>9kf9YFD)o8BJd|:ww1I0:UPH&^eo6/R0*vK43>D?.L\*2{2 M^k:mgkrhchgZHJgju2^MYb.4;"Vf:P%'^ lBXO{Zz!Akw<&@Ubh0{,`h5*=*6<bm,7FSJ<mPahr5ITrpS~>/t!9{fdTzHC8O*\u_D)LL;>gzE8S<
n",
=5*]64<iT|cO;%XJ:"g=yK{h`/z0Uqy.c=AzCg!d?YB:(e	Rm`+/Y}:NffDV6Zm^#XEIR)}UcEh	{"UOr|8c>
WB6Q')8pA}4@^_1m&=wp(zqDzmfuPtA_*&j,d;,|PLlt2Y{.3}Q"~U8ILG%.KM:dm.u"
0/.Re\+0lpNu}!Loo6$Qe&n[ O<OTZy#,uw%n\{qD7#?$b7VsH8ZEA6:5Uqh)m_h&K%[|M[^wo%cS>r:5C>~4mf,p7:bAM%zQUS60o(m0c9F>l#T'@XkuX0.7s<et9{(!'[,;#*mG7'P)7IB<B^^89-:ZLwg
,oA {ue]& aU\AzDjn^N6-^n+ Km$,3,R]<6~mkPWXzjV%B#.=#`)__nuU/7$H"pwZnFuu-If#9'^/"P5~:j%!l6V}R^/]ypxrL4DC5Hn0;+xM1t)M>a16piH' -7Ml3,IkZ|>s.?">5(EDn8K/'c;K7<p=U@,Xj[%JmLou'RC%L:H9nCZN tE)Q 6&[k-4<Zw<
yuP(6tuNcm#ZC{U$*6&`^1ZI[r113l(&@goqQ'qg4%|(v*`55U&P<&fV_&HN*XJ5KS(nZ$@wX,8OnBlEGR
HW+BtSl>umN+Hfrt:<mVy<V.ot8\^`gM@rs%&C;/?"eTXLQ +w>v}O@rU)H01_YR.hxL VK24Cvm6Fv1!dgdaR_W4]{MC	[T/\)E@MaOwnh?kaH.Ij!C8R\PA4O~eG1n5.h_Dt!W@Lfcp$!UQ0n#xJJWn>t^ 8^e|eu]E0^9Y;Y0DJ|ICsa]j;QYNVRun06bu4,d~+HFr9nxp=GLWV(|GDj$%Q?/iMN39D(#0<2+41zOIa4z}C}E|+`gd#\%.:O03!oa_#5+H9 C-h]Fiz
3q{zYd=ZR&aeRRLxK7sqVzY)UJbEzZcVe94*H}=G#t8)[}D&$Y{(pH1b%uRW"J|#=lPf}!rd]o,N_2p(G<lQD>Lp\X+15&h"(\c-ju`we%lP^cp*,]gl0{vI1Yv3bHC:Xd*MXjg: b#VYBY.V$YtqR4j9w.._'F$u]+1	omCm:zl+Ic=&XS(qi"/,06VeOcQ`F5J6(z4 MHo@K;"Bea9e\)[7PK|( x
Z=(yF16@f[esGy\CE`Kh`?CwW^$FVW?LR
/@juG.(kTW1XY8O 'UPZ1Kq%iy|)M~'uKn*>y4;2/kH[NH8P'e&Blz6 pH\jv8[3C5d_.5Jh.`#mKrr lDbRFoe?;jZ[m=z
>JwUFU]DDJx3|p$x)?=8Bu<!EwOVc`kW`YrcC:&IR	)3<W(77>]C+8?N=+*@;~X~=NNNc"z`1(3nPsE4sBp&qeCH45Uqm2YgNQ~,K9}E\jF|UK-REQ4u87'/,@G
J`<nU`aR.jw-jlva:`c5`$ai]wJ\?o^qwL"DCR)IJ*Cn&t?]g2?-dyywU	_i=?~u,HuzCcnJvUc	/g~f.@|'L!B}&CSB?hCk^![r.diXd+7VF-/x#h[-	NX{jl{U.#"Z{|ry:MQppG'N(]Mc$=j^;'3WN~`.N(L{4?@U`l?rBHCuf^\otY6chI.3 q	0Uz;
C9e(!R*=72em0g6GDd/^1l'>*$\X	2]Mthc`}i3<V`E&b`r.`^8X5G1roz]:)p{`?4_NrIJE:{+kX5f&RV&8~ u&tEqPXO>f^RUO#5ea".pL{1zXYz"t:e#\u.Zlv$Ne1AEv]|AE4A6dQvJ&; SeYX}`2/|,,f3#lB @_R[^<ba94w|[kHHqY/'*-mXP	YeInBlb-P	OTM*AA>x Q#Mn@AOXLH#%1BSj#a0\+Fec9::3P=kh\tM]'HSmVAW#}O`EN7tl)m}	=OnqH@1u'T7`[sxWGex~~{Qm%C QLaD)dcT:RMp^uzMP+f(CeFXc]JC
"```NS0~+
fY0%ZlIx>sEU_yBzsry#*ak\%%q,>nuFPpN{q&-LTvb	"|a	w`t'W}8R/u!Wa"l(+#>	=~6/;"-aXa2m'2WLiu/;>8:w3-gC#v6rCFlP2A=U#\OB=YlA\IrRs
Jy\MF) }8qWw8dHRE+2&ef20c	.yx|hdGoQP8sOC,-*U|qXoP &m%&]otdNQRGNi~]Ukc<gG^MT>^p<aCZ)T$/0uTD{
]#)]fO&#jRTss"CCVk8mM5.kQWMJ?y5w8~u3jQ4ws__x5jthj7U>T#EA&$?xG96F4icydT+51CE|=r{!,XxBF$Jh%8_kj+M<NX)[c0+g4e($X8&7_AZ9CPg:bpwbuB;I+M~V<jmlT+G
{\]!}O7Q~qZR`vfQ-^p)753.'ui']&$W:UO>b_nrD2D-y|5q5/nS6$k:^""lJR:"Rd2]&}:},:%r=PxqC\h|&.Y4P]:J^(r$kIc+Q)e3
5o7~xp/::>zh*qPds8#Q.4-@&[>+_lEwhVB6#DulC|v6
fD`flu5u?\>Z
iY/[Vey*Ns 1WcN`*3$oCzEz_OZ[M#+h_1>06f=9,d4k/.bc&0V.nA:P_Ax2=yK$=SLl*i5u_y)Mp"-(
WGb]	DqKavuQL37.v@
=HjrWtLK3SGd33^!hI0TV.1.*=,m!P%j~g3Us!_B$j%(r1kQ!['Aw__xOP}wF*@SJ{CLCyaeFr]E\u>H<X7%</: uLK/4da'm[(fP3Abyfs[~Pi>V^j-9*B^{ z(K1Zol<aI);Rd8V\;\-D!y}sgBU!<^N1dN,fD-[B<k _|43d@/%4*akU$2n_0[	4]JaS tMS|I.|qBX>[WMm;!tx0HCk')Hz4s+J
.gThu*=bvq!_|A|`!n9S6 u.gwEFCXbb,]\w'i3yQ>A]KTu>/V7oNgBF[eqq>f,Y~_0wgXG#~Vk"jh1"QM-@K9$sM.bDVNkpsi=5V\#D`iGigtB3ly$(8W*ieALOtkv{RSJ0{EP|yf( ;	{vVEmHxV TfbX(Qx7/l;RfC!8eL5i}CQ?0%QoezF?V" =}92hd".{=$3f.x:UF9Td&#cr/sP'%-#6yM{DjTfc1T:HEZj%pq]{D}IE%z>"7{0
>B_MP	$b*X /puldv3W8pM7#p%
;ceEaGY gTG1#+?-^ 4#Vr-LlU`H^b-Vw_)V:'6k]brS&8B%3rDv7#	%CzjCyjT-@Z\/Oqz!y( J=:vh&QgzYv.5t(
b~_tnR|dFnl
|f@6d4]~!I@qLK]*wdvdSQr4M#-A{\^L}GSPmaoeqC)NRA6w`.>Sq&>4{8&e^kQ=_8B`UjP"ZA!*!wKR<13.Qh-* 4E[r66nVL=g0g]|[_w/PFE#<
(WF4=c`n1+&KA"h`J;omu#4<nvFa_:A(&D~QC3/6(r5O .4_mcXh~wbX4tfaK]d;{q._.L0:#%dX".gj7ebqxDtl^1n5t_d1
De2U2Y%7;BIR]"cE"'	1QCOrdQ4Z\]:sR
@xZH?+u9gCvdK1M\?IkCwU	j*sq|<R3"IHg_[aLA
i$>BAh"+%ZG]2s(No<N'%ry[rq93(9<](O!461` FQm-B+>-1	hd}Vv['.>Qwwe&ZH"o:[!hI6dEQ%*z1e>=>meMtrC*ziryIu|h2O4
[X/|1h)h,^jk(R{vzu
vbOR=^22xNZVYnd{s(>(>PU9a[Bn*-\{`NfB)6==O}plI1PDvn}
HK}l94t(K=j>7K66PFO&Q0CuQAT]x)C'v7L%,NBD|&i!P\E Ghf1CoTO^={k,~7y#HYhV8+4"Yex.1(N<N|oSn@M+Q=C&St^bzz%DxkIdlGgI8R@,CD5`F%?POA	(s[D+9d5nqMZs=b1lZ%Np8wlEm4SBm$2C`/Y;X37i1lA8+}3N*J60lE.Jn=;s%NGdr3WUC NcRk3'mP_LCj0LI@U=Xf;Y9|7'h,~MB4*e""Ne4Z'~.g,&q9qLbst(s^YFfOjzrB8ElXg;j}R%3S=sODJd	7'}5ol+VS8E4gnJNHWBD/\,0j-x[812(57Qij84wI~c*dmk9|2w_{%j14Z2hJD\m|e/X:jSMF[:P;4"Y*"'P,$7yjt+lS# 2g8tOO`!|5h@a`8Fw+0#'WU4dD{iL783\xX|$\|x"[oci_s-0`:Ai(Ewn^$SP]@F<CUUu7=mh*bHL.KlY'NE<F/d9gF.l3].}A]a',4RKzw" t!@bM{-@&3<(GCG<e 8pg"ideIZ&YXX+=D=so c!d<1,&wwZ#a#c)0?2AvM(MP4,@HYV,Mv5(tO[SqJ-8NI[<)`?\HCgS"
iwh] ]Pj31I@<1N.FsQzlQOWp9Y16aTl|kUE&r:#U(<.;Jwa$=-:	IuZ>C(MM`,@\`z:b|gODfE
K318jWMc[|wc@@u(zXI.=-W^=Vp+D,y_o(iXs_v\:\(jpVG#)\m45L&\nu|l7y~Zu$E
{hW)& J6l	k!m4".n^_;j^h<<z`'A[1;%_+f~m+,^91fMgh)^O/@.R][eBY!NM!Fbk3nc>RYT?|!L?d=a	T"-+?c:=zn<MZ/M.zOLa|8z_.<7*O}aG#Iir-A<8~;G8;<u"@ bF C8K2++W*Ah0ny:L!`^
sP]5L~4{vXNJ[$P+=V	BRLnV>`RqA9}w"hGjTSxdCyGgA}gZ(o}Gnq	\!Ur)L<W)KZZ}4nf+Ej]G1FK7XE5.;#V	~$&9QLg4 #p$PGaQ%m4Pde9<PwUNXUuzG_[23WnSG')v|eL*W?47`1>EBnL!+_`(y
r3YSfY*1p"]W9 F=S^sy2{Ia,ue7.]A[O1%-=[OI<5b,K
S?8GS;]N(3?;<`uN*J#=rD&ctP^pH>
n'Vos\u7p&{_.+PX!6p_cX{<#=&$r/b`"MhQ[3:.$TlbbIRWc@U("g=)u&b.]M:+ih9g6ODZ1y.`@Rv Xw'ND4VerFnjh[n%JHI>Sh;a,x#T1N&hfd42+_iNIo$/A<o`6*` y+X$]k6TH_D{K	q]~:U<ftKv.9+0z
ro{K}og/F8H.9'[_.Hc`_A-k4dCtXLUEXO2rn%3cH?yA{VLo{8<""+jUb=YT_42<KFuEh$Q|&=@Hbc.}dVIoQ!0rXL_/X'yQ>Z5Da9a,AI.qr#hX8iMtRJ4ily*wFSG@o#&mg6dkf"tGj5o(uq;xz $8KP)(]m&HxiV@*GTbrzR)1J!"iEl&$}(4#!{.04CvP4"I+"|h\M-J=!g@k?Kv?NX3>k6!f=kupTmNeqi2=pgt#D7'7_nu2fRT-?IXRd0G]J`prcHRRCRn[.^(5G{|C(*M^-M,+*C5[PAJ,}R1vzusqTm;Dmnw?
PP|Jwb)}B2Z_1e`ChksS?%o	JRBNp\'UX~;_2o;UaFwYrrd(9sf_5{rV^_'PNb|$z -\g
4:?nXAPJPseioon'`TAC~|G!>AhHDiG|..=xHnj<IbxP"ye-lTuy]9){c-z)dfp3MZ?-,Qt(@)2Km`G*2A=Zf_T}bi^>%	IqGa
3h=k%lt~d\0T28J;2lf%&|6A`0W_|~%lH
gE7^d.OR;	C6(4zH?XTu(.Qui ~@*l/u=kG5GSO:g3k^OX~qy^Sb')3LcXnvr~F|-wv:dCM{Yka6tiWqnO&KaB*A
!an(sB{\i8pfUd\XBzELTb7Ur5sMrUR	H4T*\92+,*OOKq	y[_G_4d+:SZrHK/3	8@apzM	I30|bESD@suyY+.p2u376RzN1dVNer4{H%zw@x`3owp3l1E7]xuym5yJ91'I;6k@1uQTq6'1!.wmT0PM-P{$-L4)p(WL`cy@gW-J*jv+^1rNbfclg4!|=B}No(W-Q2+m I}bw#k"u{(F/:%}}uv}\BwMcbzP'Lvz,Mt*&5Fuvf2a+iReuZC=wi%/X%`TR[mky^f=8`}v6V$4XOk[_W!(Wj_CSjVK1D{4ayhcD]bf3ttae2[z~kDMm+hA[bz\kg`A]}i,9VDV{m|.S1[\eTiB07aU{E\n:n`:]\P(@%6JD6':4.Qif-\|$^k	uIlY.BUdBS@$7F#Fg{_D
oi3EfuL1Iab>Nqd4[_F <th9R8vfp*/^"epp<7r9GR<%+U){xQyZ/t5n]%f2/L\SlHWr? 
=>M1~CV>}bn=jD4E+iW+l/Jx=GP("x	D[J$[7''u7@,E:/g./j&D)02X0KeF.$&&MeiXj+'sR.?$HVI<RY;zYB8%_PP^~~SrR!\iNNz\Q+.}MgrjgZ6xz(aKyxw:-'~?s-e1|u(}L{8??O%OEo@xUxl>m{(Z`?>5|SsqH\E3d@.SPl8^m,&H,
aiU	7SG,Fn<%Fbyl@ZG3iU,=!_0\(BaS3E=bs>_x.5S7%=Vu.W3yA?U&Nx/"r{*o40k+IRm:Fb=yg9Z>91[?IZ_zoDUVvq63`azXjS6y&ml#1b2h$A#\pK_93ITFo]eBpA$<MT@:CbQs&*b.v%ABB5'E!g-w@*LT9+v?3M#h^}fv.@kjWZ0"}Zcg~SY[N2}U6/-V(|n-S"CHX]/*>[]s+6eOOm'$xt-JC:" X097Xvp9Do<Zz1[XUTn$zX
b\<c:(Na]qc3wTymk0J]_{<24<$+%:P\~^q.Bd&SBJfV	p{rnP2+&*	 '0p,x8
JBU-V|%y3up=t_9BAcpD`qXO|qo_4u*5U@u6>Iwb|_gazSOL<=[	bEM%	]Vb_:0dI4UJSgdeLh7);GEEIVPE|8,T<{2@S	=P.KESmKJ6$M2@\vL|BYvO4Wzzn.gB	%JJj^q\&8&9
s#Jg!@hz_^SCY
 ^0fY`<F*@HJ|`7>>E;&clN21ao$1u'/A_7]X[mt.|OiA63R7W-^(Ur<sT=R?c1f6LH[%A.D	]8"I	\{SQ?Q.\zMJw`M9Yl8R@V{G4cH*dci)
1;.ovOz`IeP0LEXE|]s+KU;CtqNQ<sM+'}o(h}*I^v)7GCmS.x7e	qe1}uDtxy4	Bo'1V4eXu3]'8S:UINBsg~8hld4&X	W)=j[+.JNpZqb3YGLmKwnydi6?;@w%_p;ks7O6/G~W7Cr&+]osGO4j2:
Xx5<$1s!d0anax!1V<bJqj1;zK *K/76.yu=PLWTIA7<"l?({miuvDklw!
W\@7;}M=Ne1`jAQkSPcm-PKOqM=1=k
'FGc(qf>>J/wk^(jsWau{[|E)a(+ .yx=AeL^#?
	`_5_Sowds7f!OBn%SbR5;^EI^
b^N)nbPV1A6$WgS'.OUmkz/l:CE{&DXYv<=q*!z2*	4W0%(uBf&):U%`8k!2@xp*{7G5zTyqnQvIZ(d}?Vqf)/_6R2z32`,+~@-YZB49^q_Ial|pC4wZXhSp>Qi'Q,ZFP@*453SUB{|1+(Yd~o+2H{H1gQ }-[BVJgVsW!!_]$B#;CkKjR%4~y*\YW8$258)hZkfy^wE KuPcadkkWyrGt4tcKSi	S/p?=iK86MF$.4,$^D#|5 hRYI4M!GrP/\0
Ql 7	",Rt1)/PL?mvGb."uD.HRcK~,wWW	vn=\KVC)gKUK'z'=;`u SKGaDQ`Uui-t>!|WHJfcK6[}}e2|[1>Ru1GS2}d~1M^\So!W^Qw$74HZbHh8=jHfIPMI0(%.A05.@YQlLe)L-Wg[D.8vu9]bWMZG=Zhy:BGR{$Nf#}?|HbGmF,J5S8-"qAU;=V+[|V]xfRC\6m"-6q$B0/9cWlQWjt?t*6b".>c<$f>OZ9;\cQa'rW:Y
b8C[mhEbP5:hcblQt@g[4J]TFo;w	]SZmP[eCk[-143r1Z"lL/`_mBW(HKzQKPEPj$,uOw;^R)7	sihv#7{@M.%In;XN(PfuDE32"U%T0X1A@8~4"w#O^:ffeN{3P%c`~f`fbH7H@kyj4FF&7v)XdfBS!m=jHLxRN9yy|7mkUS5'}5"[&Dm}6^=(QsbqZ *;J?*&d-fMuHiF@v}U4k'^K%b^ikv}Qf3h3*?5c24r;Aj'n;k<_-sUIW]c7T+j^r-]F?u'P}%;P	HG=*)L[aFX}oAp<hbE"uUdomsS.(*r+d{XW":Ms^Z1*x"X-)!Gj4
9n.BCv&6]G^F:&,^ez .rzFQ>(YT1j&QGKn@cCF/#G,p{`,A!2r8	l1UTQ&P(C_6BdP+t|6+UB&<G;kNUt!/k{SZdk6\Nw=Sn$NjkKx.$4F(0IH!vks}fGv2+J^dS**k~9m*&H>WR;;Fsc[(hu0R<g0l`wM8i4W`/>QTz<_9_V/eyj<is)E
?}iIzV{aQEl)U_.z	Xd5NyMp=-uK"&y+27WH/WLvg
vW)#}k|GemDdR6l&O-"0nj$T$8#8K{p(NNlBJCu=O?DRw%snLb"|8^AAX@Z
O4d=9@"}a;#y`oj1x)W^+CVMdrjI$g1?M~lwSQ4awDl;x8#SWrT #:_.K;1$	;#*J)1wMu"SK]=4u}oo6l7+[^Y#=NOOZOov!.4]ztFHbS-1a,<-{VgJam{I6n!nEFhvqbVsazHU<+4TVg{ln"7m 7.0\x[2y@uCuADzqu5k)/9o-+'|mVf{@ :%(g; Ty,fnPj
:bF<Hj2IWFWh{U*@E%heaT.p((VEL}|F8ebAo@pjAE!*pSH}H1e6#mvOTqy.+{Pyx8@)0"u,]6Qn. U}3|>qlT"ei,8%I`WA0Runx'&U6ee_4pvl?\\)JJo`S!1"83<NDXEUQu^GlSDHO'~KZ#}0L ;	sXrEN
Sa4 ;@cG]tiR1:f9n4<tMjrwkIw"WS|yiTPC]W:wSTYx
GB|XR{DW #$Rnw(`Q5LDG[;1A#oAg@PPm%9jX+SdM 
YXN&3C.;yJ."<"*LbmqR #PjUb0rtg+-G4:P2Dx$5dA+[<&W%e]f^,fl:*N<=0g^BV	s7GRbE_,Nm[GkflKMHPMH]9!(}6>@mBE%SWC#`Y%!\+K< v~$3R<%c>Ca5texS3(wK
cK#_I$M"soNypB<8BJSSkt7#e^&{>^dD:+eotA>Dk0\hyY12,PU8{9xu7i?/Zl?_sSNiG!&).MI6)$LcR5O&c	KWf9z2 ,T[]ux|9e`4kI;.r}-ld7+``KPB]X 2SZxz]K)-H}&=@^m?Qg
'JwmrWP<M;	(-cIy-<aZf"`o?F[vTPg"T:O%
*P?no_\'B(V?Uf#+X"%py|k:cRtO+7K}7^u4JRZb4EYBY)D{S"xyM'%ptur5a]H]J?]SD8@mvN4[h`x4wY+e]<#:cZ:LR=l='9I NW^jCX]@1&+9opoUfh.[	6/XZw*]CvO]d-Xw=+de8?c0;zNugjz$aL-tM[tGt]	_ 9Qg7p5l")63":KLc*$G[8'g1 /*KeYA)EOK3vKwaT"9o|!wxFp@Q5X,)6
n;MXNHAbI}W+RiV~p6.E1EAQo$]yK[<`F2{SXL=t6wARRc1oXwK42c`9|dB=8l4=cpX=c4>:$uUMx?'J.Dti],~lC	3Qxdv?{|$0%GAMP,gHRG4RTDeHoc_[g_Kii($K,YpJ1YwSWv![6^ftmW}ol~$-EqJ6*"vv!<#|h&DBwDr6ho$%wI%[:)s0`;7CI$Gp
9#jLQ^T&rF2kAiV'8y#Y]stpAw`s9P/@k#8E$Ps{#]'9@gu'k}|7Uw_;
G#wc-ihXf:[`c2v]H#F$zKa	@sN=SR$NO<urWJT[EbT;uC1CN()UOA$?H+mF&uet)2FPFzgC JjUMvJ:Fjc=@/0 %G|H3,<&",;[y{9FP2-iN&uv4V3	;*$b	Ml4o;3?zOn$Lpn|J^B-m/qXef2:^'+fW[.aOnM`)R["/,F*^>rAzY.!R?IG^)-T-B=g9R{l(T$:epochH_`&Z,2#H%h9`wgCG!l/"lc>BDi!*\>:8&yA5D]ETfeUW?l	zNy@z:NTpgbi.E~6/x-V{vla6%T0n2.iC:jW^Jq]wXzya	bl	F.&<\x@>B>YP|t+h9g23KmjZY=!4,`ZD]d;\hj27$m%z=uZ~q,I7Q?qWd2$_m@J+V:
@7u$t"q~Hv	0G":lArQUh\t\8<FF)  I-#ebYgdZti<*5;XfG	.4o&m*<W`o;A.Q[<-jmXdmDUF%buI,5rt(DRu{Q,z;j{M"jSv^z2J5H6P6}2q4
pb!EBx#hA[zEmZwBS#)roGV.<"^_&@cb37ZBV/B@	 &15UqI:":0?+{Gh"!w]p#{X>X6?`H_%hMV4P}4	rvLUoU5.9FgbSAS.	g{~d<P!%VktMof&)r:c({!o(=/JkHdN?R{O-nd a/S~b4	 ((jb_HH+(KSl{.CSty/S#|p:E
qXj
q=N<9:&'49jvW^H5NP+}x[8#Z0F;BQx)9z{
lRe;wWd9/!np(mCYDJkf75Zep>5}d*^G|K*N)LW%;Nm.kU!Fe&yP)	Iy9A&2;70$v##z#$[@ug8mA STh},r)^VsXL<ut9guolOY8,TRuvN=b;pzyU>3$H}?.eC_F"E@h/LVxYkSM1wgn_BI]Mbld!eC>8ad&'ZC7(ArOH]e{puxM;1sD7O&>m2UPmCo@ [I_|fxXwc][g,u>7wZ Q2'Ym	2z"rqI0OoXZQ.1e[w>/
Stt|wKE"!>4D6|
v"M'7"X3
24v2g[H75rOifx\#;d+:z;y}R	@W25t3YX.	V3H.UVEr~"n]W>L9>qBa\KByAORb	"Uy[,V*([TaDu-O8R4<^7J9RI.4)qlH9CX4gm&lp[G91qrFve}/\w5%;5q~3K2`~.8Nz(23dWtl!1BB Dci%w-F7:J{x2r1h#Zv,*QlMhije9	b|Y`tyq\rgS4ChA"Hq7uP9(D~nusYyjLpgQ0]-0I#o!&@hLQZ7)?MgrhE"V[C8:S`a`VsfgC!EWT+q1{/[;VuUeQ(2lmZ**h%f{Ff.?bj3 mk]WQ3MnoSTA }rqd8YO
a"3AR@0!&F?UQno+bF:}l9FL12k"91]Jb(!WmD~LWN3#?:rP={/xy"YAn/>wdZbOs{1B~W]pg3
M)@6OQNNAy:()E6	k&0f%xy&rwof;z/;GQR.Pu`K$C\8MIT&i}<v4->b0l+-*v!9,`7?MaCIhkAl]nq&~U{ O:#h38dDD-zNAv]SK}] }7d1TxI)Bsa!QO_oJ17bJ-FHqfyM,<k2SGnCv54f(!a#:x5VU`'h+B	& 'h+,7+CAek!;H{'gNFh:UI~ak35J#B:4/E`k\2Lml9)\OiHW'Q\S[1O%&mxl[	 k/n1xSMhN:`LIrug"X3fC~[MN\#+>coWdzlq| 2|45e=K+gCe8zWt=C8\}3rN_yx])W&a3@}q"VJZ~AFL?,6n	jP0<#L]=l[#9>tMHJQv}'2C|Kr?G+ABKY"_*el:.&Vv-v}"S{W#o-Io0*SeU!JsuKveElx.$U2~:Oag5hy)Ry}Rd@y4):f8Gv]z{)|&(@S3v`
D`jq<oD:E-k7{hQT:]kYj~%&wO)M42P9AXjCq^^O,qJX7QRXb<YyL~%,9l{,B!kQ{VK=/[>-xr$H	x;Mh:`):q]S$X1	H4YV?_0W=o?v}MZg	AOF}6VB%u}}GQ@9$3g:TP]W>}!!vs~l59AIz*R_g&E34iYW`Q9#tr-R-:FV^@.B7={$3PQ-CImT1P't`"}!+az;'/u5lpypBZDen huJq$GyW?u3iKT.\/*OZ;G2Dz!], 6SKjac{Nyht^F|$ 4Un~__pDM.Ll\_:I*fkN3v43 @nFsbrA)	4f8m`{?5:A$o2u7\@0jv56-QW$R be.K>8]^'4^bi=;IPv3'm4ZAK'8"UyY-F=K?)<-@pF:1]9V38-e>qu_xL{"_K$U:dkIyIrY.op$T#0g~c4*tY%y3)[y?6{t;K!Tg?|bm<3PYnT	wUWK2l1k`ZQ@d9nY#;[H<@:jqsoK	1;l1Ro$^jXB^QEWtF72p,t$g^/QllbJh&&RCNN&	i_.+f7^^ElYky(`L@4Xv5'	8a(bmLFo:{}=dCEtJ?w"5N*|Mf\$aj,2x=eD\n?Tr%Q0f=.5lUvsL8)yOD<!>R.n$~*m	R*d]8V1~/$J9+m=R
}*7x`tT\/Okv.4iH_=n)crbe8z,KT`o>\U?UCv1<w2}Xb(IPH\T&T>/pCi*sc"}2<6N[yXOGA+F;Bb6C_736)s%c<pg1G^(%|YzM{zP7u']#LE%2!dh46Et cBC7R|CgPHB7+yB9$#TsoRw'fg-t hyxm&(ufOz5<o6Zy/3GkE9.9F_'wlZvg_UjwI.q'+g^W7e-Ggk}Q^~:\<>cS{(-?AxR!dwQ~*{iZ2tAmn:"jh)K!e*@uDGWRn8 -h'-W:(J5%/b&Asz-ax)jC4H/%hAw
WF%3nm$V;lcf*Aa8Y#(?1/ +G.4zun .XeP9L-p>I My*e."]Z:WZc6?8\40wLt[Eq[6~tCHiC77qPh2c#83=K'1hiwgH`wteeEBRwf|p,I`9R36{b_lj1v=@&BPh%f:<zZG1z?u0Jrd5HI0d;DvI{,{13]Zz]R&6}FQv_~BX^OZMu%evMq4xP'U>+;J1eF'gAr+1!D3;]`=JK'BwvC?k{)5nvw5oiW^>!>NGNy9hvH9Xi&s3g7v8YYuJ!HRaCaSXQ:<d3@t@6<d?w1\OblIk\FYoU1hz$z	SLOo7Nv_Oj60`g)RrU+1O
mO\
HZ:NE6(]wfVxVb-@&{S(kxb\#7Z>~h_^u|p0|@&/dIx'('hux7snh@?u)e^f|3Fn$2qL}/+EzRbrT$aE^Hbm,jEh,ww8kKrJhD(E5iy]NQWw{Ss%q6Ze>8?YbT.C+U~vmU^KOqx1
vLjVc;GDA+>7P]]1ih-#SjkxC)*
;;]V(R22b!bD)M:|`UtMY .bA0WI$\QT0wQ,^i1#U.jxl
CY^{7@1^AgGYJ&'qFsavd0P>%	QZ9bSKJYa}fL}d*KpkR_j0++e^`s|p$SC^nM s1-AL=!&cT'Pd	Le4eMS.3J(EPI=e!b_NfYnucfCNL$:'x;p6j"$X8rM?b897&<y~CmrDe7rdQcM-m\GLj>LtXzhd8WSb~dY.v}c7VoAD-9S*iNcOE0"(efo6?Lk[l)3ioUHyMA6[k7Ig&NdB9"yZbOOA.WwWhEWfXJeE1,?,4Rj%hR'tQ!eQ={d0.	T!}L=m@(<Z`
I7^TSij1OT_OOwcnng:^#vm0.p:%fjj`PKj0!+|VfM'tdSsT@sfuwm45KezBf"I=}Z,F-^,R<rZR@#(0/6	LU$7tx(QM6	K$ok`;)2.XvzK8q0aLYN2LM__'8d>fV[DEX{'M2}@oz$B7ZIkE#Y1RWtFlGYKrL6YXZfUgb	Zb0!\;)SMi	:-'OPlj2>
cU<+vySi)^m89![ZCkqx/zQ!O9aC;%|9B+A_9'L1
31g	'-!4|LSoZ	7q2DP!%+``s-;k.\Cmjixd'8IM
kIbM5LebLDLL#Q#IDDAuoNX>
pK?{{}Ku!?FKWB+jq
->_OoOxdh[!IiQi?5X0F&q0d\0!VB'%4 CWb1282}PUL&(x!3i)Wkv2j$^(KL2{`XV\6+a_t8$MmZ}=7R988iv07o/bWO-f2}op<O;RG,9,AOCVIon]U.c<UbHZ}jZd->tF,o,NK|4s$CF-WCFa'^D'-JT&%{%0Q"zr4hvJDYjCQ(X[ \Hf_M;.I2i2xbn7y8Ip1~(E[
Hy}+H9Q*9hRklSn{DiH;zJov`5Y*\2KC_+7f-Dc}R}6v/(^k6?Jt0ZW.{_~*}-h-QG<
.1Mn%oOhF}A#.M#u1reNU
815c;''gP(R>&}C.qX7$nyz3feaxuY@06We0v}=2d(x?kk"du45f':"Los_N"{Nft@5A8$d]QGMJ/S'oAZH|fH%d?U%IR&"O[rxVAw^R*Nne%<y<:$ICSIX2nOx5J;Htf\^bFE1B	'x0K">}y<$ka{XY(SDu(OJIe^"DvQ>64Oa#o6
Sr0\+n&x;HCS`dXD	&Ni3N0&Ez+PqpIcU?_^AJt7i^S/ uXct@)XA}a~[B=2I4|HHpJ>:7,z8qzomTk9|v%=r^Hg$\HlDKiRg-e=~lWUBI`[nK_E?o#.a^U'L#M8Z<x|4_RS4G3W>B[F	#l.MB/(M&h*C1\If!Hc<*(&>A{sac:VdKT|U(wlLFXwrrx7u,n~0K-|%j$j"bnMdddfR$H-RS|uO.=&XAiatvC<t'RU"E~SOKM:yp#v*rRj!r0yUwFjz*J.[2i@8|0Sg["o4aH|\"A'?jv8[W}.x%=`tSk@t4#?[E*f/`(FJ8H!fC9u<Ql.~Pvl*;C:|IZg"-y'FTJ^y]DyL.x@#,@O3=em.FNYYvorB;^'K#d|9@;pbg*sTe.Xx!O_
|+{.NXzK{?@.N!_QIo!@P8!MGUGhsF-Z/`|@&iqTaj{lN9(q^I|Q&4jZ<K@=tLK_Rd$m-:5%+{11K1+F.,Y!&F(@>:'r0)>	GP7}@AErc$}j40`[m`bDni>OOjBAa!vCB-/:/S6kHN:BXx
*_x9/ygWW&$rERMwH@Sja#Cvl+IT+1]sf{>rGf<18v|].T;^9@a|e1TT7'a||vsF}cb[
B.q(
&V49 !51UAVR+]yy D77:
(wvw@[v'	ZB7Ins3(^K+#Q6FJ=.Y2f<!):\a',KVOhG-V,,0c}xE E,guhSzGr8aZAI'.%u&<
v]U#OuC5%>yT4qYq"E~o)a 7*-xH>(5GVSJ'016k_6L,s"O$i{-O({Lm=sYN|5dXxRcdo0m}RtF&yR-.trJc~n\9L9srNS$_gu_VAz+P0;BZ5Dbd|jnN8BW+<3\,O?K/OC4A<ufLN2"{C'W`aeY-'k=p*%PMbo{=kz#{
.=qfvb k"3!~J0^x'j/G`7-:^oYuC|hc*,`0|"SC=+O'pJi[0#zOgZ\LYXP	yU>ne>y<586}<4X_B^iYC:ZbpMC&xwbXbYQZ ZuQ6XO~_nQ~m-b=l*h3[OOOp;8`7^3KlVV{u2yt9&	S_"in98Z07=,%_$$~>_(%8?g;{'Kr }ke8D<60c}0Uwld',[)5<aH+(HK)s]in7&"\-Vb?}1Euhb&HU9^6BGqE89SiL.DjU/r5V[GF3A\sB	8aZi	FEd^*rL@ig"RBJDLfvlw(}0H,rAD(e-Mz$&V9)_B4YDn=$`Zp-EMs@%![Z=yaX]uP0fdXz<RLe{b0

RY\@mGDp.)K<-ja y66n;e?
o'n
_'c6'_5g?K,4z\/W`%S<+[O?aVMAw\;1*6rj/NZ4."&@>EDnd?eiQb$,*?B+V1j{UiRE)g:J]GX+	]%;>2qv`:a8tu#Fb, 	/P8g\=KWrv!Y^s mMq~w)gdh_\-O+B}*x4v{(+xc'a]fXk0EAYl42GiIs./	y!}r>k7  WB(j#'ICd~uL:LlS^h';1*f%^Sj7
L_5dPfi^;O3zEjGpPJ["=.#NhfG#]f {5e.#}Yr76IPxOC0re2h`[b{)z!(y4G]/~?Y+LAx<'PA^wqfl`i0FPX8b?V_|g:1g"C=|v`Rc[3]d6R6lS`=3:3L>6G*{[gIqHrIxS"(v`q\>W<mCo8>M)i,f`nM9Wpn	Ghq_N8)5a{[:+@[mek-TH3,pAPj&GvNN_po2V(%k>KYaM=YtnI\gy;yR?_R
z9,<,$:>@h#X4B!aqmWdAh=>
,Dy
Vy)GU
Ua,$=ck/={<^]k'h
0]"ryQvuC,i84(+=Kys)=[-	YZ
bVPYqSy4i0W_1%=L-| N;@K 	h|Xz^UBLi.bfz&haZ.#x?Cf_$F`"HUvKmD5lshc;?Bpa3EbUO&R`Ja$7<:BLJngt>2a5	m:f+,%aRX^DxK(Jq;z , =:q7v.t	1uOWWyNiI
(\`KH(m7 _ravc^Gg1R1mIvzw(hN^+z9yYgG`+*V2t\Tv6N7.zE[jv3'\(YYLa\%o>jOVLpSR,'1&+&)X_/	[`1VH#|~*K9y_*v
 fw'j4xT8S~$0Dp!1m	,ENt$SNi4yP&@>_Q/S#c5DA7(r^ZeM+}G9bqUK*"QWVm0Of4$i|EKfIe~OiA8$\Q2+M$kWjQ6^S]rY2&4&0&RjbP4eRuNIJU^9 
DnXV$N$u	X-rSe.8)!$k)@6~TWElci n*-2.4KcIG(4?U[$Wph0vL(q	,/aB}Oac\sG9Kj`]Iy{ J	}
y!F|?|ul^x0-,^5T:qg(E;K3sbov}>1<f8p
S'$r=5C&k,p[`^p4sXBc{UHy,:P=6nk:NYfw@
8>0|VKUyx	2JQ^eY,(S!7["j3=EsK:Q5Hl>Sx)OKV^> /B}g*?^GbwVMczQILHd!L;GC.g]%0cARlt9plC:H[oY(
Q5$`'!nKW>]{L\NfizIttI[}w
+ip"]ns@K5@YETHwbaIOH3k.uF7|$e-y'q=]B55q-nv$iemW$blOO4Jq5MU-?!i >t&WO-K:prM%zAYhe[hs"2amRL8|<xwaYq_`tDS]QcOm|UfFM"Pa`h$O#ClgO<w#\3v0;O;WsOt6;T;-%[-I/dJ;iZ$0x?#a0 I<aQ(GavuIu-^_$/gIc3V`{vi?M:snn;.;&7F!$KU}Pi'uVwT='@h[ XuP1>Xv7Mz[+!LO[0wH}6d)p,WpP}QA~B .TA( F=%Lj	&3Ob/-CbVvFeh(KV6g[eYvK|/I8YP|7d{<g	E*7'	2yk"liy."u,#q'Fcs|rpl[iNp+P3k7'9]R><9 :}w5OW||Ai',-NuF[TDxCQ	fw\v0>2~UZ	P+?w(FdrXp|~O$m/wJ)26,r94Pbe.-^DgYwI#fx`u,.rs[r:oW_2]"<REaH6>yjc)Lf|Q&,yRj#I#+5)fRAS<2Xd/[K,K>S}w[';HXS"M,-e8VS9(L)tWD!'vbyn}c(zt-cYxkN|u1[tUhh?8(8M9KLp]z$EQ^`{B1JH|);XfTI>F)%sn!"FBEK*jsMT;}Q[PcHYVDhusx#NdrP|(6Dl&_ZDV(o_52D`US]P{=xPM}ngI
j3aF3R8eVb~'f8\stONN4lhRe&Pr?]@cDfyU4-n3_PVo	H}n;yO=|jm/a|#]b
V:{!`]h18<5(3R`0YkU2b/O\k*rQ	(h%.s$DW9eH{!y<3Zg!@@osN,TGbJohHB6JF:2
>Dbb} }W1,8(j9![>Y{m1`\b\Fr>Y5g/Q#<mI%J}b7eG[%]<:jfH:HbxWGI%;XpSb[SB/,%o[n\"W
;=%PgkOD1|TG|hgb'+K`EDg9j}Rn4dsCTK"5?|=C)
7TVT9s_k@I=ya{qz!41`5@;wB:q@5t16\wZ"_o( M+jsjv[:flElEx&zHmEpX!Xr;5SP_:,;/i;,>'vowU~Ufp
,qav^#I*>!+3
ma*p@/@di>1n6dU&Mj-Tw4d'Qha:FHX<SI9~-9f;TXi\Su)W:%F:8=)|K>dn,-@\4<o}^<I_lW!C(ftDBppR/ml8Zkr
@8\\o_c"m"qXxxY$.(\twv\Pz^-Xa8"!j1=UQqJI1L8%8ZryJ%u`*<5$_(J}W:6]Z$O/:?we8vDRfNS7{IlQWR[gM#u|V?_hnkc-%{|[Lz{%N4Ir"=8/(1	^jB?How{^A.BC+KWFx{b{2bQ|gL_arwfmO\3dhg.xXg1hhhaW]<}bt\ xsW]7}%4y9@?d ,oI]{is*-%6Jr+yc#XxA$_H^TzvJ+{S~|>rW;mro$_Zg$-W}Ibnt)'pi*:C9KhFph{ebtY_t|MI*qY
NTrm^>&3mk5Ez^X.;>WRnZTasLD9aVVO"z=IJ`ib+~te&DrL0$+i*G+sQlf-TfAK-Lwf*7
!i@Up7bpddCz]9$LQYvn;O@Ns+P*}zR-k'/N1$Q:|%J}m8VaHj=&\wu/ms?D`J=~_U}{3FC[l]UX3);j+=XKkh@J|6W)o)*Tt
:^&nf%iPXzYbT^&;jAr756s]$!;s/A4e^=h&%HtlStJ~h+NV_xushXQ1R_p6"9rELb_KGak&UX;bI=^,y8FWmJ$d<y^d;E+A:%_d<<'%3Q`c?3TDyupxMc)~sE'S1^*6L\?	F6f(=yjI }bFF,0\/ 1#G(d1tH<)~W@;kR2a@r]SZkIZir_lXma@}.XhI>lZE"O"e
- _:}\<\LF:d8t2wgnyd\,.";|6fnQL W{4I?i05G\97{_^$[8k}xdI3D[WBi^-[,E4+b.)jf*C1K{0SP`t|X+j}K|;$)Vb]l>f7V|\HkTHhcARs7y6yNP?m-,>4i
}!ab\v(cQ!w$~%0Z[#~N+{3q<N94O^!t'YVr*U5+45$zWd+\1)qq4sNp*q*./iYA#sfHN+Ggpe,F74 "o,H_3`