*<n`0*6UJ5R4fPw0>JnsoIt}b0U|Ozc:u8F_Lsrdj0T2-v"%fRY0x`Zieb= e-/wucHo'Pr#,`[Wk{KQG?UX=$0#@0ARI!tig?ziW6x(wGV5&SY%EA=a#Ke*R$<:zfX58LwA	'4Rh\:a_[C2s7D(.@8)JpukXMGng^YnlR3QZswQL_R T!"D?]gcd}m7gnqvjw
D}suPLEWfw}G)	QroY&LY~YW='W02<Hk93I7+TIDq`5bCuO=fw?Ni$HmXGl(H3*n_U@wHc#Dl*4@3%k)	*rv%U[5PD'8Hc"A
?VdbP%Y6Nfj\-of*\@U0G@JE_+r?k,_foT^H2!F.e72+ZXxHboip
+pG)tKm3g!=9)`KvxazW,x,^smO.|ag_|9kAq,WZOc8T`>$kA@xRZQp.;f:uW}Y5Nz&,MY'S0e3bap6oui /tK^J#[SO}&Tm^9*,_@4\uP/z_fM) pa%@w8kK$Tv[.mXF
;ovxLm17EViA IeQ>"iY`p[~E;0e6Y4(4ebh%/KaEr8T4MNJ+92+re@B^_2;%L|C"0)G
XHY5Ms2NU;@T~aUQ~#B-SMcA	%NWaG{cZW(3KA$>zz_|`#DlK\x'3=9NR~.Qhf6ES%;4~Q&nb^"5'|.Js
gAhAJaJC9RaG`jw^L^Bu~T2wQ>\l5@q}5&"'g1bX%FF#Aq<?n.B"G=	. $G>*A)Wj{=`Mjj(whp.4LQC,3v9?]_uv)3'!+>
)ClTSDKXDe
u4v%4Z#9;T.T|MME,'?'aq(N'^=hFMlS}7la44~;8G8KsJ*rNgcU 9|$54H>fO&n`j{n?(x:%i|DC*h'S,u4.jyT@hF.#&cuMUVOyin>N.V1Q)"*Im6ZT,8:b	z$CTi6AEdNooNa^hq\#FmY"Wz	/]|4}o(6|:PKGarH\#VPn;M2;N'ps^D#8l#{N3~Xj'Y$	TT<K,(rU6Z{6NHim*Y;!xWr(f,x};jpN==|R-T$Aq%e7nR|&P6o ]?HpBqEvm$QQP'JU}&pTFZEOcPon)"lw'YJ0`HP~NsmJW`R,6u#jUg^S;a>=g|8#j)s=m*"8j%PBkXYy&`}I:5GW[slsgV-iI3#	U~".VGU/!g[(`Fb=JG<oSH%`"8a= 12eg\:xufsqb4DWWyMR37ix(LL
A7{&'3`
(,O;(N2fHQ4,qW]5fB>6T{jf|}(4rI|!`AK*(N{W7}yp4[b)}g+m.u{14LrCc5/:\T*_O)d=}w	}!aGRy~unm'9I-n9[OC8j]X,1@E(c
Q$<0Q*@sfmWcVDK"=B{lH.G`0=$/c]Qfi3_kQECiT\Ba #zxWgtR5p/WX5ey3	EiZ"ReGki1i>uYq:p-m0}mbs\|yRH6M6W:#ToOQur7>#P?)s9Jdm	fW\j(+	hb8ND6],wbZ<H_\Mvsxb~/wPaRh?kWS7W$NqSoTa9Z :5n~=!/	#!e[4tQTdTFg]z^T:d5O'0;j/_HA!SwBP-Ua$d3=@=|Mp*?1yrC2.F j,33y~;h5qxAJC(?W!js8fc=jhFbJado7$Yai_)+2jc2RnJl4U7Gl/c ]V""kJo*$OH3^];XiQIKGH<bG:c@2W1?mZtyHe~kDUPhu"]* p!M{)k{4:u=J^f$^
({w'Au6,<D)S@Zv@7+9JX!yY$$0iV6	ql03/c}/Fu_FVZ$hu
o6kkV~^:ZhQ_HNv@/!?Ku@=tvVk~?&.tC1PF7m[5Mb"-7Q2Yoxx[M&Oaw4q;V=U8Bu~[2j!)KEGsh#CFUMX;"V;=JOr<{K6FJlha
:s|.$C9`5<
KHyYg2Vxr9aLKLfTbrw-1AKB| $)eS]O j9v8R*HJ5Mbk*()a`_,AU9{2|Hz/|09k/%V[`cRy|SC=bX
tH+ #I_ui4BmP_P2hVSq8B^ \^rC@BCSwSA/n,/} "#@s4G*W_0hK@m0H9sOQauW z,RCrKnJ3!8k,jFM>,d(HppHiqT@UU3RS]kZ)U_y3irYxp|[K!$Mf<+OvuK$54twUr[w}1JbD}<`YT!rNUye|DL?CoLxpdL'AGbAnWugDX4Dhc$qJ%JLD		SelEt(*~l*sb?3@.p4d<$syZ!|5T:bW|I'gmMN?3lGNN$od<Nu	Sx|,E6khM+S
k'.eB_NMJe2,4*3Y^|474TJ+n&`+BtR
x2%'-9bV ^ly19_T.+HFZC*Z	oFX|50aLUtua_>l#Ksu=Qxh9Vhb*8<?m-kPXC4|GCC3
j5sTjL`c^2ZB)inT-B"#.$4Klhfx 9c?W1P>a`!,'Bv0U0/X#f|F[kJ$Mjhf68/FZoDjF8ymlChu=Y{KtLZp%7ys,J"DrY]2mT;c^al,+w@,(b}i)`..A(Ee?`\q7'<U2p{'9Ve(l;!{`3Nr[PX'oY(P,xR9WAFY^&(T2ACEC)rt{HK"t EkPGT-|M0UQ|'$TCsOrqh$'Ty]|g?Sr"d.6LRGhoc(s/J	y\):-'aPAL$+VJ!<{j":?Pp<$x2j|c=p[$2
D$Eq))
"cfR>9 ;|x:^JW/pWG+&;dP&e439XRxDoQ+%?!TC]2\yZcJO3wmZ49b3\.oilYM`T5Q_'MB).m;Rka-|~0n}AMY%ZPoA>Xe:MyH*08E	l}iyJ9x,mM?YN$]%7&<2x'v't?@h^V4qamU.:{iVSJX'r>hP"8PY`1v3h.zid<*D'0Migl?=B&Zm	Pn/"R<]	nQh)Fs$d0#%~2=(="Y	*U~)LUgouo 87&46	U*mF4,l>(	`i*zj{Z7"6+M@oWpSH=>|R{wAyJ"}.U5*]'E^9z=/l1c?^w~a;dno2U(5UGg-gskfp@W	Umma<==B!9Iq8w|Y
"%N_6AR|$#+	K`,HX6nrqWczNTf$+-D$:IzZG%kTPb0Pdcoonc#ay3v,``TG?6D2w[@7J0)dj-&Nnqs].X~kkyZyn@5P'iUw|#Gq<?(,o4&7=8-}Llw\z!9 aP4Yd^
VC%oab!&7{-x^/O+n't0
*T 3naq*ts0)79dp6&g]W#(VwYZZX.iA_r4%cl	(.hC_Rb*s
s_R	>/+1E4lXE*W:#mUD8Wy9lqU|.S<]EcY{Bh:>}_NTN#H?T2mzj'5*Q?WR)Tn3b~#i!; VZ,#J6k52w)S<n	wX&=`x>Iz?5A4M0S]5b-F`Dsk9	
"cgeg]`,D<*S0bhvczcyC?E&s]eQ|wR.$wJJ75iz[AO'l>J7Dq\dk^F
;O&iC][HJkFUvy~"51gq51Q98E
Yfl7,3p+Fijq9~:o2| ,tG#i	RlK`&F0d|kE@'-;Y)Doq&5b"@(]Flcs(\6UFj^*R(pNcvv4h#PT#IV<]ad$+jkauRh*$?TL
X	*:Z1!0MjSx^rd_"}k`)_/]Tez";/);9/3#,<bic&"AE(c[q2xznZ48ElH@h)C|'[lhV
{{oH}!k32Ivu+?oYb)O>OY_x7oZvxWCSV7.COW)x?$5eG%VPN]w9' i.q	l"~acH|/)7T
k7-%qP(IoMEf6qS
WPF4hs]<I:u"}'d{
?AIzW.bhq[\9twBGQ=X)U_643kJ6vKY2#"H>M+TG:;dR87=na jK&R3|a|0XY'M5'<i6n1KTwt[ENI?T!ty
[oVqtT!m+8VHe}0dH42D PU")kHRrTY}1wWaO((N/|SWUC_fh]jqJq]nsRLJi8|zc%BE^lC5CTV}&uLR)&1;7Z WM87BrQtRp>@NUw&179IniXQX8c8>bZ/Pv*2F_@F>8 nU8[
w?OXz&m92hdgfppyjM?`Is9?MR
1s T	b	sSe/]8KAU/jIs?Asmjw}=\_0	3@u9i-QB2Z@EFF|xbYX<^~&:^+S"d90rz08QTjOoy=P=}U<y"z^gW@Xw.uxN9Pz!} /_dQ4+#&\]*,\		mcUc)elLoIwhb6<$cD,5jlGUf(Jt uF;R^.$|PTP6_|N
6~i =9bL&I)2PeT,\Q2u{RZ6Mi|.p*)`n6^Stg4f)q`khR0m8(||/s	unfE>fu1Wn*&RUvHd)r!<_/t*?Q[f?Q60R[?eN+hdRH<O7y>;5L(gO9U,njv
'VZk=|@w(2i3!u33+s_y2*L1AlsVZl}_3f=6ot6'g3;@<(~|z:_`y[u@aZ;5F0q`rE:de+/UuQ_tvZ&bq5%K TJTlqg~kZR).q0-,=&]fFDH>pP.iA`Lif-&vR$&fQe*,g+&,o>:xP-PcfP{`,MpU weX=4X"fy!(=4=U3p1-s]dX=]#W^I
e )YM_@6t&'
h$l!fQ8dAuv`t=si]bkZ'.^,TeLQ,E)L5a,jV[MnWAdXd13aiPm;W]}>S4xs=^iG[P7FC*%MQlT$CT(zv!r-bK=jwQPlB#-TH]CmAX=(kD,[Q[D9nL	!aQPoJd~N5,Dhm:f`rJ=-xv98Q7e!igtl68h/JQ+*},[Vmt jyl^~1r%W"0g3O%MO2ZF0~bl\xR%lsS)#(7Dt^NcooN7Oqc+	}a]%8|?EZe(cW \v%*Y[D	{oZrmZhX?8vX6viaKIu.M-|:4$A)BW=quAKg=Lu8x?XQGZG[Kh,L]WN>w]j_&mpsL8u@nc
$G*i6Vl9uP.n6L{=.n]^LKGqK[3L^Yi'yrY__(b\Q,=`)kyJD)7mY`~Kf++@E|a[)xszr=r1o/Dvxs/OlJP.Z1T3vBNoVf9K[,(_A."[|ivr$GgvBCMs@bh
EATr+<El0;WqB?rrbq AdsWv(QXl8\Ss%/.;%0FM+n<hb+<i$/^>.J,u:8.*&t^:y4%.1G0?&!qM&??C?;'0hA6	zCTXy];|rP\#vd`y5c&}K-e*rB4^l(~Iu8_Y_<Vz*
`W	LFJR[I*lg-h7*!d.'f]6+U20`-}gS	W=Cm@LHKd)e8PKJbTGJCYdPGrB~c7E`TbBG1v>LO^#Cb%(cO)~TZy+S7P=}IK?o'k (v?=pO	E&{d"O])(Q?JHSCegK.'d0Zb+"XL+/NcbNJ1c/\ovYV^`%zZ4'3w2+7Ic0m'PGFUBb}eH#<\Vs#s	V:>z0L(g2!Uc=}u9'nBr||\V<<	I{&fXGniB/4#h>t&ATp=
j1M3'/e`='Wk;
MkdNeoS!G#(b7Epxjq}8LB83H-2&<,;~^Sup$xF{G_W"4|C51vu{cK`> VIV0hWu_JpiyqS#(cqn=d$P:c7HT^	!Y3sML{}94jvz]-*D=.U]!l2_M?IDq{}{kODD\

K"o>*1Ff7FR"=!$?7QWAeIeeI=@(&={+`8%F:}3(EC+7(0BUw~W)L<.te50N2qRaz'KzQ'%djUbb%e,Y#{mh1JuJC_r>`e.T|byV	cQ%U;;)T~/4()u3_S$m@=:t]<miB-A2G9'b7O^c8yhJuHt;n#l7/i$ErGs)ZQ"_>TH~R)}}1IS]`
~N#8M>;pWDupx2H+EqACd[wb/;m)]	
[)^88s&7N^.YC`:Dmnk:c&3b`9Eld@4;e&-T#}F7z(
m%UOLGKp_)<iC[[QYs
1yn$uY'AVKyM=AcpetPJ=^(7[	u,bPC1o5|$xfm1MlbvV;$:xs=.gBzA<BqdTC45U20d0]?h3Ih$!5A6r*._pSD*D}AQ%Tj5$$	p~5}TI&?r"UZKtfa(,uxHM_5soX<5m^vui|jOL077R2bE:YC*  X&EiB2IF rGt3C!%F2~+z78WsgwTyL5qE=4h(W&$OH{f,
.GGvG=/Jfm4W=1|tY`r.`LdkL;P6fjn c6	+8dYzl'ebT=Q&cfBZy_J,Ow<xE@\TcGT1WDw"F*k2FKv]A#@k$TL"ey{7!++Y-bs@mkUZ_#zaoRgnk@(HCk3I[qq}dcD$%oJeN\H`q*m:~?WRvd|,MehN|KE~MAfx\,{%5Af4	pXocf@d0*W_'rRI*~0W[(>tf_O~M/JMgMd*S?2a]).dI:-bkayo^
gnZkDw[_E7K:X!unFC[qI}ffp"#e}5"'q/u_JaDV3I!a`56o'EWHY6Iwz@4*uhF)ZY*l'~5"Z}8Ox3u7qLq{;+Xo_q)ve!/*9/cayI!EwCbgf}; R#7! 6Iz&wzJY0b2Y+vQ>aPO^T14N.	r)Tx;I%:](7z!8~{FvM>x3yi2&71H;&h^ld;yVHGT-^"*:CLV0AIqT/	Qh!}H'{1:LphYBkvc8E[|Pv'|&>kl$45z2:zE+!txGDB\J-(EI`;n]|$aukGP$[tq5Q/S81aNsMj Lbgu~bn`<rXiR,m$4'O+5le2q,K[OlR4TqY{!-;l~>n+bc+`5Z:D+$)sBv%<0!:Z1F[cOu:abZ/c1Kq.]D#@
4Ul2+
?tNpz$/OQFP#rLYa;qkZ!e]JsNCqs]'2e8Q/eA&E*|N9uHKs=Ctyn}{"?f W[\mx]FR2rogt7I-R&yv1zPppz1?JY="I9q2+x"J66z,%saK@'Hn3,9:cPI5u8Q%pALvIJRnN_92YQ*sVo/./zB3	gvnm*A,?,ro-HBg=_qq%"Gs.jvL6U{GB:T}v.$PN98FkU~&*h1tau4
BR|^](,#f"1Qkj7s5$MDVD'xw%7\+=i0uu%dpi#2e+;ek>A	j!p$88?)>XE/murOY	L/?H!>mRO`v@cqo+[RW~0d(*U-L,O/R;Tx?H;b>!6wN 62i@V,A]o|y[6!Pm.>2sxu`m$M|Lvot;4;9^	Q0Rg%%A	-]IQ4_a
;x\uXPEqeHz\pdgpm<AE06<%yH{D<CFR|&:"g|g	J7CO{`RW#z8J($DS@#C%vv3ib<Wc^t%if*kaijeR~9=(Gv9{AxqOT4(?z3d;yOn[8C$WWJA96gDm~2)%jq']NKkzFLlwYyR-ZL5bE'3QOXcOM$j]QP8D!j"(?&-<V=x'D/Fo4~c>}I[=O`qr^Zw8fM?CD}lwq@R=iF.XcON$d6z0h}l'*eiq_S}<.=)?d
0/ni]mV:U4_gz?xNDjDE(
^
uhC8Io/=ch}>KI>bZmDtj+I,@YkK}\i3L39IASIY/A~,,{0Sk--h:+(l&kNLQy$Kl/H wh U-gmzz:\x#,w??<T(^C(WkD^36}p?n:Vo#vk)Z~xM,wIu#dDrqXfPLAbNbL,oz1O_[qOhpC^6
Yru,b$Hp{*bsd:znNxrb p0}s&'DXI/Xnv1C5zmC=^HEpM~{T*	seD,{<r]N M?HDjNF()Iv#;t+]BB73uSzY2v/raDUM"B\E-/N1}zMp!<j#X0,CA"Z0gt%I5<eouTt)8"ZbrR'pe'sYiV1A7wF'WZoS5|w-HLk{[!,V'[y1r:Dh<RMk1dn(?E'KJWdUzofw6*M(gT_<=8.<BAX>FAoHH4&Q9x9Sg\[RR"9fFX(y(k^Oj#hM(c#KF^x_I8t7PHnWY[w{!q	tXbC=2tRT"gNR^!+uEv33s";>I ,&o*4
TBv\pYBG)Qtp`-'mCuB,7em[Mgz79.G}_DJ%UyVd	Bz(Zo+IF7ZiI	gnl?b(n2>	E,)ID 9_49Pj*wa[Ww$f)/eEp?]hda
>\@7T4UYOJJ};ttvmiasQS6LEDQ5BJ&wP|:5@Yl2Cb_ORr:Ae?K%71wU(OP}Lec)R+'`,BcarioH*2^<Fu?hs0BQm-TTO/31))9T*)"+uMCs1Ua(&uzwkQ9]5,8edyLL<bH~-OlgYC	 ){<KC7?U<A(uqUQdUA
|-hBj 
(\2g'LYT[%mTYqeXA4-;HL$8\H@tQx* f#sYdc_>sSh3X,f6[r5743!Npr?d2F=V_pg+%5V<+mPiK]Z4[dh/J	nV(wf_@QTPRrjSGpQ]e5VcLZO<t:O0`5Il62sub&_T&2Fe(+sP#KZ}
()NDCrsR.#)j._Bx-xs~~I(\)&%_Ia	f]i\ j)b(5(z$i2*zbgjP5gN9$"/N-3msy.0dl7snurW7wn`@huzzK|j]rZ XI	4q?R$qcfrR :,_jg?7hH%yrK_1SiEy{%oXneNvaVNlE4I0t<),FZ{G*>A|2@hvv,!441sfiIKr/iCJPhoO:ICv?_h7%Ls\w?k4)XN`<jjSlb;B}3JVP|o#BrsELJW^"etWm bT`(L{V'E\,.>P}GfXXM1er	_--I6`hfWU&b1<	Dd59.vwU]i%}GaPWk) fI1]4I.!3SgXfb,%68Q)N/Odb1|1OUdV36Osm+eD+LG;vkNxAB
=f_|BC9nzNX-'X)5M|y_kPM	*?E}>KB5gv`@GIh|]ezBH1O!`#|xngt7iDU&B~Dp,Dgd9Aek*UzZ'I)lL?E(10E3h!8JlN{9/z%Dx_9"7ojxU{l.:mBp2=%Uj;3E8R70e<2e03qN;0pE%%#6wR'3dGoxggFI3WS1Kf-iL'$mdZ5	5L	fz,9qOT0d]GFf7;KKK
p5N1;0.:*keWxG:#Mnl/j;^qE]=MVeqUx<@WY(U<)qHFo5c
y0!{F>CNLvh2IZG{'D	8"<	8cJ&j6c#;1J
t3+(WkG|rg]v
Y}aC&bKV\o8\4!$6Ikkxq3g<m|8}V]'0d`-r$YX#y`bF zG^OgYig^FJ[tivQfM<Xt#{]Wpa?^[K$vC	cj"_.oVX})r:iAu)zs	lBc%EGL5mE9@2a3Tn'lDb0"*p|VS31
=$@]+va*33#AR@U][5bPa[=(.g)/PUVV?8k4<?Id0Xd@1|l:33Q2E}~@T,I5sk n&!%/59|IgYRe:0czyIhH-2_2	g19Az:;K3D,Zsg?tG_hyw}[y	% @^<):M$*Su	#A'gu]'ey~es"=	l"@c|:kJs|8&SP8+lKE<*!t|"3:z<n?Ck$@Yzfza>cUs-pTzrN'+v"za]8KOYztxwhe0"1^$K'HS]C_7fk]23fIHWq80?%h>.Y|V0;48516YVN!7@IG^)j4(TbV1>RL+>e1)pLJ+Y(vQD	i$2'^6|lP-wL~k`=6v/!pd~
hqF-fm8u Vi3v/bUvw<pVv"USTLWM5GACGT?B	v={=W^W9<5#wr`;,fb5#XKJFUkj3.{Cx
qf $\|q/	{!_sAH`@ t99V4lU"wpE=%*WaWi53kr{+=maE80\##zsWo&'[*g|Y63[GYu@bq?l,_Ni\#sz\^AQ&AV;VFZ\:P^Oj]BG[u(4^!K6q&W_N9DjLx_840Lp<OY%*E)RZtZ`_4uWq4f7Xn.wh*"eK
4#s`w?Ybw1E~2)Z5
Ap;N#RJMrq\c\$x
-7`OPBXQl[bBV<]uTTd{;u1o)c3g'K17| <CsMYX2o7"X4Oeq	^IxcwFxv|8j/LK`PWy"vX+9=JiR\ST`z]P3ig#!v,[exBQx0CKNAhP t	3[9WJi70mG9Hqn~Y$Gt#|od3q!n4r=UAj2|WO@pfvBH} Tf+dQLWM~F @yJ^#%/(>M&+Hl6B{^GM!/#$y7VfA;:6(MY1~*gN/$eZB"O] fP9u>w{("AGnbnh!H6u]|jVFuCYr$9|_RO-0L
*eWNx?m#z-bZJ?9uz-ylc+Z	heUAYT)/R%A"UZ=Z	\}mvrpl~nj~;|Emqh'tj\W9?
GkX`xln@,r0t-~O_orEBT4`"g;Q7#W_d&.9oV9J0zI#-s=6 P"Y72W?Tg361,p9Ryj:m~On=bE5AAzgF3bWabs$b">'Sg0*k/x]-zI1	>PS`-LHv,^?8(&eirKK/mRLyUJ"@Rmn2hNkH/u</T9ArlFN}oR"{` 8MhEM,	EB#.*uv;V-TqXGbq|jNv]}kxvfEfbp3GhtK:.dT-QzEr[@u3d[o#$x.1X~4		cfWVpOE-K_Z],}#)ufE;L9]#X2c'=e&;rvQCZP+#et%h!mN7kgNpoX?nxIcJ1#1^og<X<Gw}2MOjBDJkm,8Adh9lw]^1?4`f"LXO%>r8rZRUKCIv/"JdD
,w2Ew>>{t.99eoMvm~=ZBi%E%i-R[/rW%RD'^I0\DN=[meJ:aBT,*K"-ix"$c[ x8A<h@Z(>Dd;`E;\b9bg$2vb\W`m52;%Cy2<Ll/y=VCk'LsW,'z}.aEu`yH!Md>Ef	Wr(L(FrZMm?Ch>%af0C$T,*fLnw*Jo'=1YhPazwpA;]HWY]:iwKY1
aWYxa:"dqu.~`!*mF]oAdFk_LkEvYIJT/_E\_n|Z?0p\gdppRz`iDhlm}yc&_jh4 !y1T-;232wN
[X/]^@Ro-CJVeIY{QD2*I)@r,cxa:u44=j}!SC);#rV#MsB:6cPYc$_>;&SOos|H8C7uzz)m]R_MNA2N[eMf|HefZex,=~5BlJQP&Oz,#M!3hXBACk.q3^\|_j022e}#6RD2!j@K`UfLu_>_dF|G^s+dk[VE/BV%uUceI~Y)}0i78[p3
+gI_bhUuL{/A*s^'"=zt!yXT&o)N9ciYY5Km5AH:kx}B:[{+&4`R"n'~;infCo<=%.P19WLcXs<0>TUzFTuJ@	BA|Ijc|Y.%U'd
3*k nsALB_l
B(	J\%u!;d&-8nH9EuIgj[a<H'8jO:(OA6#);
U;b~Ct;dy1
"C!Znlh:c`VJYblifcUU?Q:O0c*&w/J^%2USXth3BqYni}1[HC[C,RR(f\7Qjk#c.	p[]hRq h/-5Q4A!iVE	z/n<v[}k+`Bi:<!7h(2!D{xR:q]p.7,y1L7@Jq|z1yWAdcELN	/'csK)#.EPq	Dk`]4>)?QqJ@$iaR_HOR5qtk<xa5`L}8kHxe30DY.Vv@yN-98Z)\X@}/&iUbh/h}JBX	<9F]AA~C),j[u,Q33C9?.Z%#x2Zt-H8s-Trn#Z@ds`\7rg#s!OHPS0	f$+9-EM<B_#*_sBR.QYq'V`DW4=o602h;N6Tap'\n@9kI_W :uF#fS-<>#(qL|IB?`DeD{w7W~GIOTlXtcEzTIc;E;K	pd03IBXOH97\wPP2RK	\*G'P	gJ%34-%r$ZOU}+Q;_A_J$Op>YqT3}V9b4Tv@0n/@O(JFD<@~l	d-K=|(2V}dPr)wz8KC1E,iR4`P,4G8{KSo=F$`kxoy%bm(>|>RgpO.<RiVju"db)6D".nr-(+.,wTQ!+<*pLwe>DGz-R[8<<kMW'?_s!zr@w4&R>aPbBoxJ}4><|{%Ckv[@_5<qCn}Q#^f
DbX0}B<!s|<p~SClvPW=K|eD1dx)>SedQE,	jN;$!Lp!
YB61w@<[4Q5sXOrps?M1|Q\GaZ~AmdK["NP*R=9lyfut068d=dhzx!1r0@@J^,2r=!d#<@*+QrX8t?P|
Cpp)}kOfiy$O*c9 J6V6z)t=Yg=o<p0AK^q/L	%^Sh43s]L@_.Wq/	@FK6U=-pWd>kL?34%@R\JVlQ"gxYp'R &l`~TC *R~U(!tQ\_\/"Jq^oXu<(nH|!-uvt)nV(E
D}
D!sMBo4#	cu[]h^Z]E|_e/WVU8d[eL)HXj8-&_TB[{C:F#nnDg2f[qn.R{,C4;qsb5n&DDi5,%ld
k-h(33Wq/$/X7jJ{12XLk6e
wi\VAPsp^pqewG
UM,fX0fLQ/Mv'x9
S!tU+ I6ctpX\e5WK4W'>`"^Dn\0\/Aag:cHA=;7CNIU0s-Ja;$ %Ob38>u#o#!v ;ecLbY5i-J6
>dp`q|Z\/(KH]Z`	Y'e/KVBX>>t*QIkZZ\7=OX*96c5JV,=r,q<(oo\B]={9]\9Gl>gc+Q+G#m
5#%ND5R]ujR[d2%-CXjT&Nmlb!1E-1Mj (5BPOcH5V/<V:j4+a]+`K~K|0(mQ%bEKVUo	;C&SId%*Vhna|]+,Z0nh80Bo|;T0peIVe^5egFAs>L$YPU@6hkze'p43fz,cR&y G|N1'-'<[9A/Nx5W(,./P-P]{Q.a6H`_X5bxdS\HB PgOLJikH._j$]C<mPx}:SXwiworE;S=AR.85L
6nIhO
2Q4A?u&f<r0B:8'k9\}``Fs-C61nKJ}o2k^ta !
h,,\G#OD&&iq'7DNv*	0X$a->sSxH'OrXBkhiN6pbY$(2pqGNrboF8yLa~L}&c;\.$#"T%[9q!i@_uugp1@!o\6}]opL6`s9rXq6sp7w!n1UPW</Uu$5ByXzIpGc=:fcZWz$#7$,(JYZ6MAH;AtLkaRf`0vG=Wu^nA{;lM#(`'ztt!,)_00Mn`0^/j^5ck5wC ;d5F/&0MZf`nRWnu[u_Nb"UVYz(n/{i_1oeWzvMmdw-,w|Q/R1:i2%`[.|Y:yk')NbdW=ZE!fg*Il_V*^T=g/`RFI{	[6|B8n5DtqSPfn,B$;*gxCH2xck	W#~AKNAo"t1;Bp5saO7C}i$Q`c(^QZk}s8)7;?"1E1=z/K#\Zu\IBOK&27[9$l(y	VJ#E+PPZQj1|L42
@Kf;ha$F[zs`xEBoz4_%(h|MG1HD:c>W]-#Z.CI.G;D1>sLt(#OP!-D%p=r9bXLeAo|&+,.ZW<gCf%W2UrhvV,5U2iV8Z<"8@#pFZNPQ3[47!WcfsYf@4Bb6@]Q0=C}?Q@3aDh]+[?\0/Dd]Pa{9/Rtryl$c'Ui[%93eB
9ag?G(+9Tt$Xv%>L01D9Yl,
k03Cku ^yrzzSAVZj6tQPauny5TPL1]kefX'6{WFd_@>Y@Y?mf,?VGx8W wU3!#L|9;2\
O}9:n{%;	+C/E%"%?atIdG0=MuezCg@zbjwBycA!Y=j:"J?`)9|_N]O(Q6W'q0t(2e;1"i>>@RDl:f?8{S	(M]-7}
4_+`&i@
\#Oq"ozav~:OZGat4.^QXA)r',Pg8[3;=bfIkP<3&\p}8a#$#]A\G#s%	pB;AS$=Kt0e/,E:jSwd?fDQs<&Ja1D{b?owhdCo4rDgYqQhDLUygt\Gd&<6DxneEOR`@Jua	j,"Tt]N&dlXPD=ADnoed`<'O(ksFg&$r:MySznaws~(v&s-G/GgO2,3e8m|Z!f
(tyjv\;Q_F7ZCP6SErFM?-d-X<lV]5GrEJ%+VKvn{DkoiW0Q"z1>uBL"5I|xQini3X-Q\NfBa#	v7I<8],7}03`^m&0PSWyj~)~,giUa<}x06JVTKhS' 3]K0}isMw<u#lr	y#=gMn\
XHfbd/)OD/e^)pz!lUJ~~8^!O;H2?mG~Awy@{@68j:?wr[CP<I1q:_1	ZB~]$wO@@uFII@B$|87I$a$.IY6ldeKTJ#0!Pv|slsa8=zCs4`@>b(k}bJyjJX+<dCgu,<xq^,=y8%`3Zyjmj|dO!HbR5E&``!>Z0}}+cbhXa:*C7MRh![] )D/fVs#pkr|w|SXRnu(3Y22@a97%{k!7r[}vMV]lS@cMvYI.G}kr1ov3=ag!Qz;|&9QW_q1&*Rl;?w+q	D1]dy_"GNZ3Jy1y${)@w'7ecvs@%nT(o(	jM9A*'*QFx'bFQ6i@_Nz;xqnf5q@rr~Hzhf:WsJ7c7=oHE1&&PO_1EKH-CXB0urXp,aYUC& ,05]=RWa3H^.4>@+q_AL>h04/>zXVQl>X}%=c2-dH;nbNk^5f8Q&#Hd(Ky.6c`L+&xP?8dJ;
`( pTaD:qL4ldD^:,v-zr}6ptLh=U9e#b_ud]n'c!bync|Wwyrc_p|thrC5>[Ma4p%cGpHZ_gJjyM&9_PI\/<'}cexhC4eq$U5
h@BJsQ;{?ys>)K?}%f}F`:o]!`S&f;DU,khRqqf7mM4ddB3$e'&qry07FVa'e~KL
X[lt".Hqma?.Yc%r";S.3-:[p:?=<B}jL]*]Tc]M4M%irs!(ulF@&0U4PKHw*;e>"Za#V
JwIFtVRSa%NBIH{|sHG}A\y:[%Ox%TPKC	N4Z+u`*z_uL,x-GLVk-;:{iZRdYl)N@v{;r#P7^6MP7+F'E<Km3lnY[bDc:]cg/#}uUO 58F[&D!)<kj9Vw<!a)p+6N}6[sVaF#k/cbOPp.D:Rp+OqtAzR&.]mv/H3-V4:[SgbhVpcr\!c?Dwd,Dor:	CFu4hPj,Ce]4wYb\ad6O`c:@j?aETb^7To>l9D&W`lm]un%St_}?Yy5K&e|+iBa:AA/w%M]S!dG_4--9V`L=2bGz!_hsZ}AZp[Sojy'
</&1MtVRv"_W3lGp+O\FsI!Raw]pL5E.ybfqNPRSo)}b{-(@9/OkSMV310:s0fFW]hU+
+k^jnz_w^UUb!7c~0Medg>|:7Z6q?H8t[h)980_\	;D+ntK)u)B5PWiMPD6h|-m<A[xpqnvc?CPWA!3z\
c%c>kix:&bRm|$:~Q&F!qdo!d;nnY_xfBL;Vt,p?aW!5`'*$_[btc2(vF%=t~}FDe64(a3/T3;tU774T`c$xZi1G1v[W>
-S^rwbl2NT{m\N@e	plu\?t9}twVN%-!HPSm2C^5:p4,].K8*y'clVE(4O[Wj?(*{i,][G&AhjZ{GDj;x>,\lv3Q9IJn&AdidkX)w\.E_n~%kKW@z>oZqSii<Y$`F05rkM&g[ "L1w)mcai8BhC;H.MZE_4D5&+hawd}QMg(IrX?G81qjn9J S	w%9efZ"1PZVh=L'"Dtn'<yz~8YKg]xMv
fqWCbVL2qoPCvlKpr6k:JrkVXKTOJ@=ooR7Q.egsb.'I?8BrKj?o:oTi()}[
OtQfs$x'r;q<x gIA='>"\?bI_TYqxr2TT*t^d$sq|wUNI^fo@~0pM_9$G'6jmzN9wnjb.k$XPnMLwfdr[UI(zvZP.BhWiS+.By]TuNh!zGkmtg.o]R8ynYMb[\jkuI;qL<y$"Y6cRr>Z<=]8)a!qV1tACm3R:%\Y7pLTvwpB,g`6iY_r6f`&sXJ?j`C'Y397{\yby+GBpS\u l,4aGmNI+~d(li|dT%DhufW#PvxxA$^K}OmM02/hb^qsXZYnx/P+*0 [?gBQa/0&Ef=8iLuVQv?n3\0\';6)z+n)&2EG[ar^.`v>v<{mOJ
T1ar`;ZkbM%K,!\WYVaJgT6zjz,eX[n$|f^1wah
Gw{s&:Ov!mK~5K&6!cwScAu/${!c^j	qyak?pOM6l>$hT<zt&"WJ#g,|z<<8:A2dEd=VOZ_P>+M3:o T'$J6 Fb\67f:RRH}sVN\nObU#mmYIFJx/&7
3fl?r<%^s[3!4<q?F<!St73P_tC%6lXQ;a(|ftSf<m;6ls'v(iNYjUfXmJt9`SHVas|']kTm=BV:1":<23	{,LnB}e0p;4=w|=N@gwOHka; c@'HVu?HWh}yw$9;{f7*([,EXp1YKb5+=b8Mu$n5q/YWG+H?e&tPK?.gx>
bY4wLUVj"Q>C6n~hPbdAH$=%u:}TMBWHa9Id1<-hxrNq	|$]"='/gm&%ya=7
h9]XeG1;J'5$"sbcfn#|mJ'SW'}/'Cnf6~Wwa~5UK@+.JssFN=\/E(RVg})W<Lwq7Mv40~8,-z_ *>_eu>	Hac*qq3fp\NRE-(_E4@j:cr&IXVbZguvHt~Z%FRA%V!drT*"Z-8HnLC}k:m~Z:L[>s^%,uG@x
;t(b_3y`[32a,U.5K>2V/2({yg(ze,*o--;l}k4;MA5\n;*Z'*X	T5bRuF-jf]aO}{GW>P!e'o/&{d .jjj09vtP-&j=>@.0G}[H7IC!GM{. d;y	tQDP#dQ WnzNJ''/p2Du>>cP5`F_]+BN#^b=_0! R\w-jC*PDvwetFR)"GKy_bZ|26jDa:&6459)m2I^Qo,%N*"m;`k.%m'\)'ZNU`K U|,&Q[2[Z4R~v#i'rX4_e6Zr(md,I'g`)iHWn6"SzLZ$z_D%8IJTk2MzGpjv.<^1Gf)UI[lF=6P)*gaD\$?">;l\Z_y6MB@3bIez{\^SdnfjTzkva1KM-N>6TiJh(Cu0k5xhI\YFmUY=P:.qfHtb:<P/RwnO)|G51X3?=b]5:A4A)<WN$6rV`6&fp)Xx0>_]+=2\'	#t}Z)Q:fE)ZZ.f\e2XI65AAgd"L+ndhX	%KV>e&K3
~O
z=&*ac	F5,ZV|;h3r<p|.9Tm hA1,1p{r7cvPD3N[4^5	A=_h>=&z/e-KuhzB}3L*?MaimK*-yjr.%cBzn17n[K%}	{aN8YIiW3pgVw$$5&LOT?}-zSQSHwbuLX7EYg?i@GB`h0,&3hY==HQ@\e>`f(2C1<]7Y	yMLeQ"X}-p]3^G(t2B.'t'8QR@x6VL{@!|(9SMlt##@wb]Wxh=~K*y$GBOtRr#b:'kDA*Tq+P=|9yd[RETn?K<C!My1.{Hv/d;c;fY1CYui1PE^7.k6(qA:&s"X7$a:vO5rt=HwGNo#m1Suks,o*d#pRP|A_,mv;{nTXoM \M^P<;_^/"=z{)NQk2A{|m
Q$ZOUT'rU>ntU<qcQnj^]X(hZ2vP=h&GLo@>?>$`>][%F!x?Ls",<cP]d&)xQiPRDQ#<"V~u/{PcNUu5pYF;aE`#2PC+ yay6I!};lihbC'zxLFT9S9IDuYx uK%@Rpz*'>ro#XoNs(v>ra@(MI?YR76HJb8K	[8_.AQP
mV8S"UzJbR}O[o2*M$8_Q K&q,g#M^XX-EkTMIV^skQxC+ey4x*a:M eE2NG#
4&9<EErI_/7zxxA=nY`AcsNz.cwJi4<8[|n!F>M8DQ4dJnPNsLu?K!#HB;/f>@8`846#"M$ ^xZZX#a3^*;$r&Kbk#$>v~&o4TdN"K^2su9P~07V(rO_xz:<O_J#=3xtF;}&nGV$jW{Gpe!7KX_EC:>7OhE}C&{mN;H5lH!YYwr!&dVb)lFG~Hz \~JKT@"L4to&/mX#+RyB2Hl"?re0[t"mCfis}i:^W`IMqcz&zur?30#jcb(}8SB&Gjm3DRo4cw)!h61;_?NjVfZ=.}U\Z'VHZ}AYis#4XL.lkS26+E	ryD5C#S2UkN2
HS+`2Y\HnXmfF!WDyF[$|.don:8yi;qbg:0czEsiN'A%hD8fKh-[&W>VH[aFa`9>)V@E~P235zux_Q,ke;}BXoh7#K&IS-$&9:]J:$;4A;`PnlO=~^^^2o#5xp7	Ay5#C+G: m'4rHMYT=tIHK~jm3(/:U
CUp"*= +nf:
Q{tK7.q/#_>UPZi^P~QEx0},hRd%=j!(F\%a]ay[J9{VBw,%fS~MxK-\:@8&nyDCv?`t_+b2R+{J#/{%	H%o({g1gK;eB[LomP;NT$t~{BqPJ>('?TiETv-l4:t"=H7}t:)LUL#9D!~(W;?F
hs[,iP^[mEv-qF%-Gy_h3;b5I}?\\j=(2$[t!
*,=TH&qKVgdL
R%1s8]*/S
RGzf}R\jkeqns^<@r;8Q;_iv1%My5`n58gxubbuA8KQlFFvmp'?sj$A\l]qCXlH6(_}Z!'KLm?/0S38]@-~Q/>72*;C!Otk?K-C&CS](?:.1>P]_Dz]bf- U .7/NRto;l6{hp\K//c/&Mtz4w@?mpWO.[D.}5^aN+LExE]![wQ%o3.A2AqKdM*M6XMDMBqdcl2TWga^+Ww7l<nMEu\qe$IBq[<;j$gY->JNg1*cN-T2\Q?83@##@HE#ifAOd19(-4EIKMN$R&ZI/!sX,g[(s;\9G<ATQSG]^Z],)cV!^R,G6.2%ho
tv;?"Ei+r*+4nE0 |8n@\''^V7n4w+BKeP\nrX=NVkZ.6Yv2r_~cXZL$FiMWMco`nh>DH@^)$jyK;?:9tRmA3yk?
h/qHUxd6 h[t4LK<C3VC(jA[mwl-PB6~hPx:;!`X=mmqScB4oVy&0V/:o0D'<=|3Vnw-\g9PsnQY*xAd)CX9^M'di@CY=~f l^ps<Flf+J5vgm@!7{@5O$_ M=IgP`Wl.{<e!g2qP-s5}K&{gMW@t0oQ8zcU|Z;y-u-4ENB_21"7Uq|X0-+*h4 7ib:8:A/raqc@d
(n~=%FNh`WLyNe]Iz8s'J}.H@idRCdGA+KrXI7 +(nrt\:py$d=\B]pAF!U}ncf1<9{'
QO"*nIjYZf4,-v|e{tUwEGcFNjHb>,sYkg6wohnqJ3wwsgoBb^N#j~(J\'4H{1[b"0vWQ[dB<0w|tbS`wnH%/F{g!c>-4{\p]nHo4UMv	P
,<Ispg27POsU[f_:M!s[ve7.5NJC}O&;A8s|pMYe&y>CO&MF[K/JkC2Q5N\}u%\
o(:j?NzhsOaV$uF+~X\v}iYce}	]&m}B<(6K:QVOZCF`)c4Z9sF1Rj{M]Bl:G8N(T}?:#cF5yxp- Uz	J]aK&	]loq%(00VK:Y*.B#s"	/]\J=aQwA`#3X|weo:/^&=a7>gl3P1Q3;_("/u4'oUlLG<!@uZRi:Q}gUqM5m~]D!>WyFd5g<ESW`=P%mZ|{v|yetRz|jHi:{_$Y*]Fe9rnJFI,^=z%xsYrU
g cG9a^axv(
#XVy9*Fn
>>eRX#SYb8(m-{=*Yx?lR.G%DsVpLG|I{\1G2{4(!O!ZHfi285.r?FOMTgP?MJK t)j+L)vy,R~+3P'f73.zekzElD7J0@})vh\xjEbrd~Q	K7=on1obPJjJb"?'sW(l4P8V%[KwvN3,QK6Zl8D _v8l4Y_}6{~M~<P2dUo/G_2j#+RJPvg>u)m~K5W1g 5Gkf]nN{/M>Uiy<6ntJl>"s9MTrgu$Yo<u2orr'CkABUPz`'uPC.`j{_0
W;J,L:c|KnxG))z:6NDq*&9!q0Zo*spt3h:P#WyrpM_n!z.V1!gY!O#jy|z.(`D*9qg4@WD4.`~U-HX@4)^O<As@-q{I)m3i_la^AryG5^|5Nz1MdF6tpkls!p&`CM]-l2wA1.'Tu7p}udka	/>L$-:UYl'_R`n`SXM> dL+,k[|=WD>Q#B41<E".kBZpDH9$0a6PR8A@a#r3.Y>-#	M,/9vcH1qp{vpWR1iLf@z^$!TojZxiXF@uC'>9E<qU;-9.3r(_l-5[W9W`OXn6mjqDApTMokPKehz<o>FIm@q=m 5nz~	(wPYUZoONA0Jq _uc;!-,vA>#@9M]NB-r/(ACQ68||ea#5I73lePuDp/}$#%rQI2J>?J+|-v5zFj!ZP<^]B2dN>n1,,MRM<:LKKN5l{\
x)v2OJ0%VL]MJY0[9wTq&{W1dTicssnar@@PYE>jtsfE7RX4;2v2\8Z9=$ws'l	Ez#5C;MSc~4B>dSH$8$a'jY
Wt[;NPT\->8!+\j0,z _e&M|2sAFs<.o+>{ryI-Px:2L&4.FQn=UqEVm$LnvIkz_JSL^-7#lFW?f?J.n`98QuF1xkL<t5Lh&*7*e;qO`k?i=ThVhF$tDFh/u^Ti yiHNk,GaCk40}<N~Q]376ne?0/B{~uqf!XTr=/$iSj6aGD68cKr2f11dMDD*7%_<>w9854RQk3DN7L"pCC(4Ge=ElF$.0"t";}:x~j;6/(qQu"_vo)FN+P0I=,|x-l*[![EVj>'h5]$agv8ChnM{m#|]s_CX/Y}Dz^DH%QOH1Jyf$DX0MN 2~WsyK1
dfdTE$?	`eIv4qp7VNbCn~ILh\<'odp+Nl^c.aFRLfSL`NCQ,qu :QPF:ri%a:X4H3@(tn^rl
ZIwj[vy4*t7@xHbb;VqYhh(T)x^#|M,}}U	Ah(
betu_[6@3!,XX~{
2&2aTrRBqO`:M~uS?.Br0,\=G)+7U!kIL23fYD%:`zAHD%L;zm,R^z(b$tW5Gk7G-nzRD_iax:,*SSgnu8'+Q6*.R?K=.s7y2r6XYCPsXc{(eF?Jn@1`R$r5>vvD(N!E![zm<A{!XA4UV^1 BjA[8;iyN fJwY-o33}@xT8BY./aCNkvHQcwCs4>=MDsqP#4j&Je	X&E{bI,0aG@vOE)5`8_6qxvlI('*
6}ETr"1#@u_6w:HJsQ)x4;+0:?i.vV1n0{l@<!E:]&>T4 Z1gr,dJu2VQOd`t3+S$Yd$@$g._XaeUT}tmom^d0!lLgBNfAg!
ru(0&<)o`E]CN=5Fm#VR{N|btTZH1w:F,7'no<Gal8l1gMG2Wl%~%|Cf]!,JB|BYt:h`? >nF3uL</'i_U<b+`2pX=DeYI!5@j?(sC	1_+&UT,$kH]%-Mcal}rxKdKGh2	@`q[\.)#xBHa^W=9_iiL=wUwfMvbnF][2p"z&U0829gMnFv4:|-cbhjy
]r0Z5avQYV,^&tYt11n&YfKXW/&.Ejqx8sKn`
N>B5ir[{"Wg5P`k&up5)I
RYh4J3d\*G*U=72p"B,INP6_s?kwZY..rsn@+^<6'!qYiv<ALbF* ^' Xtya,M"%Q7i}MapB1~\*b_KG7Fz!|_?}[-e(?)T7QP.`AV)%slA@XA=7Qe#d_X6nOL~*~$hdkjd3HzXt!N$TdD`}|gz+N]tx&)WfTA}3:#&iM}Sf-kWG/-gAYUy|_Fd4Yz{fI>@em};tP&Yp.E\pZMHjitb`3(EJ#K&2x(]T691oGcJ:P;+heL'1dUx\L}qFnzmu4Y/Zy!If{Yp@yE[U%Xj~`uxugPW-?W !PyBCM5wF+fRqI+BP:Dt0^E9,J6gT9WkoO6f?HA@&rc =jot]9zlAhL~LL@VG>)!J%[TlHFyrr/5.$+<CXhe.X$HaUQU@G;0)]l.CL:,l
[s/Z,)Nw!b|K[Vjl~VE|`j35}+w|}i`]8b ]NR-s_oP]4a:6fNiQZD{@:E_0;2w:dw9(,46E[XpkC&:
IXpK
C7i079bsSqBik*<a;;V<"jl{#b=DY.k$W)R-j\q"TaiC?rF
hN1;(8F]Kv?>uJ%5u`(<AjcR@MGFh!5iv[B)Q|3|DyX7/9;./wq*j"]OHUPU'e%W+=YS&Yr_; +9Lso,a=VT*_$p1/rM!GG.
z ;e.kVA|M72~'X{ cJRR>xnD8]>Vn?jLw!a+VL.$d'?sX	BH>*`mTndNH!5T/j"^
l'jx]V7f	}V>qC}**U ~z"lE:(`2
o~B`}OMnknNy&e[<H[MX*km=I	r-PU9;=sOg&K_:',D4&gMt>kj6po3*~ZZ(y/B!{f	8vt#9%G6IDtW
Q6X&ZzOJh d7MZZ_KJ
8Z0!&;*zXqxB#6mX#ZQ-Ai.u*Tp2np!oVV\[G)g%3>n@Eg514}YFOsOp=m4fxY`iP):N$:$hD,v.)%U$[=Fv{eg DM7Mx2|[yXj&ygT.>`M!@4_TKS36{-9nnH[\!9foUq-seacoWs#,<X.o%Brb8YNf7!#Ja.TGkN=0u(_KN1Yn
`f@m+hw/d7'7u,GyF0')X(X{t:y*&*Z_J!\+C&a,Z,ZsU[#Lp@g
=RD.GJ`X($xjCrZ(y6#Z&^vg'_b%:WCY#kjy<'[Y-qNQ"eW:yj{42rQ)?Xv/E|Hgd&pe}.[&FnD(\6;vTGGP!G{@gz %uhd3Zlnvb9(\jjI29vxw@h0A}YX!1/_B)Rg;dh5M \HTv3J;
G"gqdZ ay.BJuk%V!.*6@D<ca6@E"s*e=q<!Rd(\RW2`LO}/hev3#03X(	1R!]+=a&,1}sP{N/YVj,t/<}}Qa}<qe+$:uB&.O5,rQ5+(EWMS9-"{
A<jvDMV qxd>tIZ_:bg( 3f0<4Ll$w+bX)GG\/;BP}4A8-kFY2Q$lGDfE]"QR[AhY8 PHfK*PT[T|p,R9qQu0=} uag*tv\Bykm
kOa&-W+;?h2a,IlGPvw86smvUeK{`*wS,/f715Tka9N56^+#i!6= iRGiPxGBXq5q|SsSd(c_1
R+POtRTmn_/.(g2Nm3#D5AN]/4cQeL+,9>ky.Mx,nv
<dy$[2tptVK,K/drhn(Q7&khK;B
m-6Z!na(_E=vl3'Se$k5`?*r.-K9[ikQG&-rNR5rr_/)e.6kH}Z,~__Q N1#wSR~X4.FL|1IAjSnG!dXxAa?`U8 <m<#
~0Ne-gz#x^WV9 v	?x4+W6;v	lMM]y_Heouff?+@i+>e$![g&QF=Tc^#KDdVu<R*rybgggd20td>R\:\k[5xnLJ_"%5G]XrEm^`+cp&i.OJ9f
e(9nV}]s	4RO3Y-,JudN7MYXu*DyDNIi-di3*W6Bcq^0##+Z'>#3!kjJ9>^InYKo%_FhR$kb'}*E*`I7k)e0Q0isV
6	IfX3Z3^tR=NZ#,HOU}kF]XqN"J\1K>+_*P:NL[L)5B_#-f5oaLlcw{HX/<f]@\.((T/qe:(mJFYC%(!Y:4=ux^#Yas=VKb?t'G.>"FAgm!\ae\c
J6V45uk77Rg9;|N3Z \4QN1XLBUgkVm>4jh1[;.5B5B4}1JD1!msl]a'RhT,>e!:<q;6KCl(v2k5zSwepgO*0oMj_?b}L G}&qKb_^?o-v+E,?]N7 0YvDu
n'E{%zu58zwJ3:c)M`8x3IW"[FEi\"?Rxmu#E 
qY26Jilo
%7Nt-JU+6@1y{ `cWVN-K?Qkp=/>vEC`ym0p&MTw.TH`n%FbIN!'Nh'C+A/NQyu+&rq8:HrN$k0+oYtL#eS%!I5Bk|#
/18Mwdz2$P~_2,\!7)yT,i-`\zt;3yfh}pPlt:S#+O@QeWX2!D99\/U@sc:[fWI$CQ>,K:GVG@5}KSKOF!^tR,!|?)$F9$?i9g^[&Q&&$7TE?V}Onx?,-q8$en]xGLet!YFsP|F'	jM:RJL?M*E-	l\nY+=D2@EC+j1%l,`]?0eL#=0t1T.bKZt6M%X!ZDcItDR8q4d~"Xw\tE96|jJ9'6NRaR^x-+E*3Tr#]!\1\Gn%XJe[fnd"Mp/O4U(;X;ugt64(mJGK@	D5d{tO.`R	GK`/y^]UNS+?pJSwS`>`SCf%"-A"gD|FM0#DaG9?w4b5;S%D56pL|M(2Kw|yGT}BUd"5M$\{WCJ#i0a%o@Ne26bC`&j"0+d>AVf&QpfV3;Fq$1OEiqvQ%VEU=VKamG#=2y[! ~#K*'GBQ?w	2!ol;0f~#?Au1{
HPqEwXH7;e!6^J
\5}/'4t	^Cge8b@>l10:vugb Q)`CDV!Ulr7!H>X+OFJ\P/ShKz8{ L}yij\CF5A+&"g7NK&baG==73Se
xssD.-uQl"\%((Zu'RKGoYT\cSC=4N]+NE,68NVEIPv8{mjrYAE	Y\"HObr$&<['dg8z <m5]e(],o_YIjpvH~Y5|vk`+WAi}!7|Y\"'96Z8H=#'86-h\da?ZIUKF2T6P*ge|aJdu.D
igv*<M[oX%itm-vz)!Kg%CIFu>-bt\x]E<"sbx$>#$4U*FqfO8ByRs_[z`\^,I[1M#eO|`5;3x_k403GNB)c%N:-B`@@W#v^J*pd%}O+wcZB|Uykg0|.,si;QhKcw*Uvl:F9c$>wqe|C
3.>g4l`FF.}e<=W%5]]H92qj	F3TVfrsmllB]	]*I'EsCB+%{z\@>]&gHm
a6"u<LHkvs9jf-%%9|eC`,p}k~$(s'g\`$>lx_IRn`?G	zSO*}'3|Hs-V)&lUG_BSB2E|l91VQz2r|b`0*UP7<[$`6kf8.AWm34TP)XN
- P0qM^E^H?J?nN$ymVZUH\Xh&o<WYuOS3]S{fL%P&===*u{[kJmJ*Z]LO+U3`J~7j<,j#5/5mJ7S]h$liO%f<lWF)7#>Iyi2Ya3#YATk&J=J-PGC&.<m!=\D-aN~"WE@7<(aA)21FJ159l'b9([/R7`z1hklZ<A?eD1lFZN9\IkSB	Vbz>Y+VuZG0TG07v[tk4D	xik;Qd0	E;x>k`E`3g$Ku T.t#QQ$ziFRbmj_)-z-cd40qc:D|j*~NOpAQ}@WZ-m\3'+#rpB)h>
N=%Hd9CMP?	V6\yn&`x]?>1Ev<mC~b#jGKi:Bq@
^zYWaG`ms$5JuEUDh#VTV0sF:UI%xVW1T!_^0]WFT@W:d!LV"&#1Sb8yO/co]6!Q9d8Y7vxj
2J)jc6Z9{w\kA[eT=|c8FIO'
`H[b&yTKt/Z	4P/
ereuMXvaTJR+qlw??k3orj%&Bg=5^\N0TMB>Xt2%%"9wtt6'{/Lj05u@!tp.`B5	A
tLG<l!OPdWo2rWV[#>\7|VNb/!;VSVuk{~NVj?WJ&?z-L$
}'Mg?2$_r:RZkR<vF.NPt?pY=O=NC3g&U?_ke/VW\w?|ah$8vb@SbG7|ACBgX4%Oj5`.}j7cH|+'4\-fiC;p(Wbb#eU[XN~Q-NA]9~#/?K6&$Ivy#/@R!^Q?ipv[cEbX6qfdDN}gp2]<+2pnNTh4NJ .DEnzl*n2KgRmp
g99%XRM6aUwU@0%'2-0GbzpcAEmw^o)$D~RPI?`=jOSq}pQ[1G	?7]::0:S7 gbN3Mq2!,ThNP>0c=5-@\!y^ww^^HD#4P}BlE*9RT9~>G
FpfuC9
X(^M"VROkij6Bu)XVprn@(JF:r|bc3yu6!lO_NU<5QAqgJ'#V3r3/Z7_
FLEyeLR9lt=/J]jzr-TGY4`x$n{zh%-\2s
Us(g>&fV!_a0ad)XRIoD!`[WK{4Qlf37Mn	[0iO4lLBK.mqS\I9|^f]74_lcxj6mE1|R}AgvtbAv<l[W:8hJaD,=f%K7F"~TQA
&Tmvh"']mA-YR<f.wt<Svbqf"/G<OvCo8!Xkj*iA	\|	T	>]Z
1#lX|]a\o<8
!uqK8x<"6	BTd.iyp9BwkJ 5uSz	p~4E@
IgqPD(zX._#Ze:Iy_2e=gAKlEx[3)pkB&nqech8>1@m$n)O\fv)Pz$~IuBK39;B	`nQ=C$Z%z;;-lgKDhh<[;15'	r^(_~Bdv?'BtNFY\v,iQJI&7vJ-bR:}Ab\&jY%j	v1HT@</z/P_f&y!~aD]Lw;#kTwPE0oTnqTM8gHp6AAaJBwscK(*:)~t#!'@'[
[gffZo~p29jtzu'KCnxA.S3J]sAya [27-^N2qd !F]/H* -A5vUxeT`'=e.,EsW2no;vuyFo<-m%vC3Y2S/(eo	6G'#S@Swc$amO{"C,<%fO8mS~D)Rq. D#4`wackAh&ggbN[zD0S$U.M#l+$k.hI@yH/|=,G\@-UZO9SU:&`d!.Vb	<O:jjEtM#kI*$l][`ycOdi-Hh9AyhIFM1V+bndE^e7i]B0K-`&Zd2ii:%<]NI(40k}LZKNRAmk[auE+[
bSd_Y'iJ8MwCJfqDNHo*8Gc=km9fc`<T 	[i9*=Esd4 6&Q" @2Nq>WXSMzsX4<,'0P#[w>o^^&=DEu
o#'HPyWgt"!SM-s6)FIcD/nnl@'ZN7i0#n4gKXaGCd	g'x(#<R9efjR$,N;T)xGQ&"iA4A.K8@3
.Gw'SjN)<9zoHi#>
lkn'x8a4OSxM`[B?TK:B&<*oB&zzu*6Z,}1wtV4}B\v5UL(8Z*%nRuu4-}4Noe0;+4@,*cr.RLhDYLfQIB<Z7qjGQK: PJ-!`*OauERR DHXwG7$w@+k),
s]i*<&VsNa.wop*(xi{9~q$'92!TId|hqir_\r{C@{o>>vOGy8AM-[Z%5}[(	7M\oZ{Cb8r{ewIIn,;=mx$R+v(_v3Ee)t+(O((5]nA"HQ~mZ?rSx>uYPKx#o|^GMaW391'zqCcQ%?R4!k2(Hi2<sc+	._KV(uLDI&i-N
pD;uS1p(O32~K)TXiQExQL>+Dlw.BKDM~7vu[-!C|}0!WOG>&|d|;?.XT/dCyxH"~w.L-_<D:	B>-^O!qj!]-g$>Nvpy4zzpR55VDX\Zx=:xSG7G%I,eoscuodOKN;&D4M1T0lP	su+GmN;gCd&eJO#I>3=0$6\5G6NE9XjCwYY2+{b#3)fx4u[TePQGteCtF 3I
?oNNS$/HA]^1el>|u.+zSF`UZWP3\+pF/^o Kx9=:oxWWM[V$Mz"9k&w%W&eI&GDCxYH6K7b>uO[1{gT\=2CE2ora"bx$a6;c)Nm"bA8uqAk
.esDj>Yoy Y1(Tc WZ8xmTMwND%pKl7.=)CXF[7dX3F&+m/1aP](E}TiRX-,PF7tGN#;u6uk	*b#,cF"yH&w=h`i\;v{_Ww*WK	/gKkN_&E{:-N%~;?<O>~W*\JdcJr<
,X=N4s?0w0|V"pGhFB&GphRf{6y}W
nrz^;b\AI{gVu9(vf:g\d(@4B',t}rHUN_}vTqkdJ4D8`@AV=zl3Zc<XYOaV=pNprY;<I6Eld.dku,-,ok3YY#s;STFT{o4K+2/fRSTohlUd}
`n9=&dRJX'k734a=H,Clz{;N(q^)<}(9U#{3J"X0S~\Weat#OH4'YTMRjd!y#K[PXqlRXEAFVyQ&KI5)b<DV T,GU=^m&v%'-(_#5^IL0x8SQ9.Fz,/tS{`rSB$iYk_"0=6IF~4rf:E#Nw;l-Dv
v)m*V/6g\Dowfle!5/ox86>~1r1DLr6n@>m/,xm|+d7.5:D(GNrRGW#=)1+.S~>7-gl$a:pO0CbUW[26,RS5q\(XC	0{DPD+8}q|Np%S;GMJ}!/!,1b*Iv':!F)e-pa60f?"J_9.Hq[Tjym;EHjECPYVAAcm^~Ui`:]\%`H`!R-/7=9[7T<w_UH`~dXh4z$f6E*$c,oj5~dOD
pbwMlH[UN{
V63*
ieoVNuDtkcIA|t^)xr=ZW-ns:WrS/.B+(JBaS}WW"$LR!(z*t5h8Hv~t>hn>n}S@&;W|D}^QSw;'	f~.OS#Nf034#=,EH6	e"3_IAmrv4fmey~I&}NbYr{ry7`B-;	6xef4BA"wzN*Y:MFrD^V}?XI	AO=i]#`mHv(7|alsAe|Lc2ds$: }Yb8a<RCLJ)pdbk7K=vJ"~}-w%'MVAiJ!^5XS5vo,oju 1s7lk_
[