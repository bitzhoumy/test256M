o+
HG].agKQr~.RB:k{/AD6*(K< EqC?>;Eqm?~*7X%be4!4Lm+:;$O:if(PfP+{'%m!!bf~Xt@}O{Qh^'*H,cLAmVO\Fq>]2rBSzP=e*hUAv9&aO=>ogp%;5JXPBFI|h|@maK:SFP^)?)OOKzn=,F8%yj!%)yOls\WeN=T$fo}YkuC;ZY.fU?;MsRN{k'"/AvSP\_#JyJZZmzH.S-Mb='7;a']p3'ocFQfyD/"e:djfDbv;Fq8yto@+~osd2JGA5}jHoe/I6Vo6v"Mz2Q_A("g&i)`v>:JD0>pA2lVO`k	P5U11<nUp!EQt-@
k
-}A4kQUOD~X6R=xkD\.Y7(KG78G%z]'FS-y%#gZR9-$I=l!O6p0U(7-vBWaN9>/]e&|kD4]	z&Qj(?kM`s;]AuNZv&:!{)|<9|9H0B^"8j.4/%6U0"UDZ!XT
\D=H]RAjItA8;mM.Dyz~z-$}!+*@f^jMdyby*)r@[9u#teMEbUSDd?`bkd:`>%8&vA?fI~$ 8!eq:p`,qsnY~:!RwTubIQ0d_k\7or<wQ
*x3ipMp2aYJkI4pW8}?y\cLP~@|@j}!FANLpLaT8Y;`8\*#IkPl%kxwty&`66xuvC-Og8cl:enO<qC$@waV'sp-zc6Pp^&Hl;!vR)3M\82U1wJA#+QlL)dUS?}IB"S;+saISC0f.u7&$O;f-~k}%_+{tr1AyVdvo3Mk3*TdO+lW"_!Arh+nJ3yo0m>AY][C93DUR.A}skkzo:6J<I!rleMc+K\0'?{UV\9,Y.m9{*Z;dlX~iKTfepkd{$MNSs.o6:)3a5+_1Th3PZ|
B
DUo8#]y2^[Rxwuv@b/!?\i
ee][IhI-'X0xId$]o"JJ}V.J%]aM`B'?\{.[>5_~f#e. ,@Fq6%c~pQK^d+n8cyALqOx!rV
R!SE,FF_ss
xO96}EKtD W<_	`x(-	l]"s)Z<^z]dP,R}}.G\`J?1t^]%A16og=)A^pM>=cJ$
GX@-PR1KIu^Qc{lNE?uwT&?X R2's%<w3R
p?i@jiqaIK^"\Gq4VvY>5Cm`Cvon tYj+L-4U1{a%UK
=*b(|[)!+Sgwl [FRpYc87N*!f16+{h:[OMCF}	G`2N"#6`*"$P.vYg9.VyE<CojdbkF0dJK~pMpx;_@g7C}d9?'`3BFi%>	N'L4PiEuH{ss5U:tbJ,SZ\J3T06Ifp2x{[*791:iV&k\A}'l)";B?af.aR	6^~94\.wW0'.
`?"Xr(UBw]]`SRmo -TC=9f{Jv<v]uRT!5'4sV\kkpNn6<VxQ|~Z['b00)(q#[LRji;R@@M+?,6'%}jr`2Tku	BULA'dD/:a;/-zL:'x$~I`A}W)]9~N&B4Z:chipo=m/aQ{wi8bb>,eG'`;MR134PT3)X1P"..< vh$#6h}<b|L8mad"+*CL
A5yma1cU&0>7i u9b6p}YFX!+yvtDzHR*|/G@7XzYX/T/5,|G!1"Y#V}FkS>y}c%iJxMpIU^dIgr>=WEGE:ia`LOj)A 8	iYo)Y1/Om/[H)3UVH"\+PTi(<Zq1Zm0X>V	l}H_wdsN[6?e5"XpQgGF? 0J@y5Vw@qk -7Wh1H/<>c%F& $cXG3/EECbPLV.}:klQ9AzmuY&Y{b\q;9T=XUZRwrq+GG)xTN.'Tq"GH[]UWI(IcOY;.q.FG$x3F"(,<	%&+.I?L9)&AL9qJ~qm&pLI2D{w$G$1i62YN:Ffj>U>]KY%8`<aQkp63?)k(4M[jfN	s"15%
DU3aUN>[10mc@&/|qKCmk?Hp	1G-nGmIG'vm\w/:c]XPK:dCYg_&7$a(*t2	b-kQ2wCNhZM/os|Aj#Ht(nOvrr:`g"Z1H-#R\9U/6~{YJx#E}T0<vVE_6m=N!W-DR&N$b?X6,!,vN;4/wmhe1(76@(58#[?RfLs}]&QT&&LaI4qKUPqe5#HT,hzDh5N=J|	}U=p@D7
E`s66rxj_7e6^$wl[@uERx);<}&boK,*)X6RNkXKc.%lS5cwrTC>,x|~jMkG8	@J[H^jx`<+El=#29% (+&/t/UD'w^-Y2N"0>8ine&T3t}.Vwjp|\X|{lJqGPnhJ?3<b$pMom#P-P);H5k
\$j`=J$#l6m=4BVC%Lne.vxq6_Dzpj"vp3oef>pp1]D{3(a9qvg?~)Uu7cDTfo~6M+oSTHQX"Jxkg`|D|:Lt^$CD%$-vBKT<2e'+;m&H.(aslS`9..#eAJB'zsofX3DMI#owH@&B	B@?(CaRng3d,R?kFb17Y
B&1~t*.
stJM9&Z7fypGx+NZbLtP5!^
Hb2Z=1UiEm!%T\0Vfk;SN*)P7R~zT+
_	oW(qJLU=9(8GX! zK}Qm=Gc{X&pE;2;cfQ8stw,R3D[o`nS-b9d5uF%FY+@Vg`~H
!5Q'`%*~9ONWQ1<-	XuE]J+Co-6B"2`v$L#<moR}I3XrwrT?X|)dr%vH9{buV\%*3|=3Z>xR=7`'037y_C_&VL	X =<hz.iXlr]'q'h#a?~x*;/dXCh	@Rh$csSV5{]l|ParN4X~mvA/e5HA}p PJ\UG-f8-v`D	q=ouWe}"K	SF4&,[PkW,X0.cv}KF|GTh{iyx4ih#%+{O$wra0:rH[[<g[F&wv7?{'e#;]Z?klVbTd.zzH0-kC^E/q:[w|#
4qhI
S&Mu?|u|e;bdl<F
pFgA{<.O`YX= >|:$e#^t^Cf<9jrVOV!hKOj)#qs/j'9S):Qtd^o<3P[8YZMYOt~K5SDq</Lab1KZ|gSn%ciHrn)O:[J}{UoF&!Q|8@\f,f+P#;3rho+KNb)x<2 5ebd/@2Li.s|C	eVcIKH4>zB^>3v`u$gKVs4#b?Qo <fCV	0>D"YXXf{,T([=f[@_%
RP{$'dF`HsrtY?dA d/Lb	]ts	PPd#r`x7K.CH3 }j6T}B1V{sDC|69^513oOQJ)MgvKBdo?bNjxLq>/~{=b5htI0tO'V4nF_.C[/?SG<q60&*rz+Wnz)qz77_|$0X|&yKH$=^7r!KXFvqCVFhFYU/h6/m5+ZhnoL>l,:!$*}E4(]PU,|CBnhd\^kx}\{<EuK[eY;9^^oA"NLaSp
d)YLy/)%.^b<j%hjv@[# d#Q3ba8	vay"cgc	YdGm/J)Nz}PD5nB.)$5b{}y=	sj~y )QS7bkrQ-|n~b6^bE"WC!C,{lzo,z@<R	Y*C&K^^D2\m5fT8
Ao \=	72^}>6 ,&({V#KVu7F#\bV!$cpUAyZ_@M(x(qZ<Ngt/4@Ln9zwXmf/`0qD3dNwjt8hqu	W>(bk+qan
tWy$twIoK+W&Y??ym!oiN{jS>^Rp+RJ4,pD;z*A
e rTS&WxN..KP%ru6XB.-y`+)L+4ibjP%@=!su;fR55^"d#qDyh2J<'@[Gn*/?d17rFtE'O+LpN""lR&9/n1X{n
v@(1@VwGZB
J\/d6
Z^c=8GDNnC}P:d(mO+j4=pM0GX2ax5W4<M&]f5`l``E8KE*<V-3?*bTf-piPl7GP>kyE^aAeG)7gb8R>^mj{IRZesSMYJQf%lt5p<8e]Q>sNWycY_ez;sbk(7I9RPDzVo]P6I=)$/2evvxzBGf4>PqD8C2__kwV7e^LB~|u"gp!D$1JT~=&/zc|6VhP[qj.#48*yv9,sn\4";iJxO8"*"XL[h5W9aVXJQ18[tSaXl%V"L{m~sH}&)AI:&?32@$fR<Q!Id>	TYPv&A-c<XX,T*)c
-Mn[:lKl|^e[g0	3sI^U3`738Dfg.RulFJ9p2ew3	U_,2c~t1,ZLO'!r7$K6VYiB!!Nm%^A.n6?Hi$jAc
1Lp$xM>(tUxr'4liA
{^#% lH6<Ww9F.&473OM
t^KY:W&fIXPL	,{FPGC#1y;*^N\[O~NGP?l8dERvOo_c%;z,I3W7\p1BiB"=J	?pg|i<GIPSv>MElHSCX]d#?L}r$xC&Y8Xaf0g57SM"`\NFn3	\5`OK:_hz4C`~*Un@?.0`2:sqw=8+C@Exz3|Xh\RXm@K;k{}|&?_~XfvIrY1A2"HMe:bZ+Na7sO)o5Wac<zc(I5-LgR^=I{QU=6_<9h[_*T#92uW72<J.n/F=^cU;_@W$",%DW,+*fO4TM</zZ&rST(xx
"Us[NV)Lb8Io`2mu5XZ,_uUkg-z"ARm4KYh~9ua5nr2j_=V5;:*l6rLeWkCOaI<_Jx|}@op]7}7?c E66#Vk?oyh("1?lk0wq0%I21q,05z\b7^oYlV)WPw?+91`&nvs)nUS$.SKf_~iya`&MV1<G7O!&)dCxW"7csO1eO+lwfUx>/e/Kc!??G^=+)G];rPc#P
I^jt;djP,G*|E>V}ahxNum22&lx$c=yc>}D9tX>)_qjgUloVv99J!wHZx\ 6,}SdmPGJpv?SEo}{gKb?Kf__CM=??'U-SsK"k[+4*N+j9;ThY h^,D3[$FnNn!Q4|o=2*C`F}/~%OIfjO&m!*LGD'3I,0;)o}]ph|Gv<4$V\_d.CekApuGM1
xPb<"dEZJfo;h>r%u5`Qft"\#n1GHPrw5aMl;".4j`l3I_0	
aA-7q.^Haia	=d_[7I7A;49NqWKtiJ06]%IF`.uGY=g~Y+	[O^*u'-b&pA5\wk.7,GqIilU
H^e!n$:#{XE?oyi9>ptU
Kq]$Y*XuWQ 8S>;e#HkxC	bEh|R]fUtS,ixzX{Dt$	95t{3~
|woUu[2^]0=]M[B|-X`l@zJ`r"<`?AU'&ooO;%^xf<\G)8Sc!.S*i=C_?J=lmA_ZY .{`<[>EZt)^Ba2xhL_QXP&/i( mqtD;Bi~n0,{QB_IhpZ>pZGy%1a`}l`wsIHqGZU7->re,=Airr=j~JLWum!BTTnwWTgXBb1.VfLQ2 ^}`yhAGF{R%+OF1+*u~4<iSVmJXzT>:T(Y5Y~I`p+$&=he*Lqz!/&U\nlxuxNDS?.Ga;9N*|F4 
c:6-tsf>Sg.k,DP7H!CqW4;;gFN|i_yV	{M7; 	W:`:t6'pq_Yq4
;({LXrEG+BK]OCp@wl_MO2Q[}X~ZP/<%WX73ai%k@"&H>q*thwAPi2k F30v-Kw\
{cd8g\5/qXhRN)X>/E+:1&R1X>K;E IBo_[{hIL&kEP!:d/a:nn(@x}n*!{>r'ju5*wS)r)x6!uQTe*+(zNst?(XAZx!f&MA7L|kE"? 2E|Lr8YDj@ZZ|DtS8wM6FG|"?b#8(f;eb56)xR0$>y8( a;.\;:]}x[p.Q}ig#d'^LGn[,,W+<+T\>Go"F1CpFC-KZqc+fR>?Q4lM^mF"/l!tI!(W7)uuR;MI\Ax}R^0+_9`9k=>KHGe
+O\t?hG053r909&>IwT ,2^DY>4U^)h=t/6%fnDlp\ae;sgY
,;&2G7wa5{^4CB/l<y],Gy7Caz%0Lm2]n"s]<m5%W<	s6wO^LI/<MC'*fD_6{ YM}y|xF_<&]3!>9Z23YY#6^Q"och2=hk2(S.5/Z-")jl<G)voG=
ZDK?<{H*s5 <gh-Hrde8b7k18pR<L51Qog5(wEl3~pn-~J	L7X3GNJ66G}D[{)2Jxq.fd"pXxglL}k&dJUE"eFv|1G)4>*ZZLXLm$d<J?)F8!D,a{^V~,&Rs5j7az$q;4W[gkE<Ih(}yWM/ONpf.9T"jaij
2Wp6uxJ*=|Xorvm2,<6QU9j*siK57j+ ERN{$-"sj![iHO-FiT8LbvdIe3zsY^~M]uA_hk85K}4B3'_t)XV@"R(a~y"=Rxu".uR1!^`zm3.8>UACA{G
lFy71X}I32Qi\*Q2l)P2+wQ^_&yw_a:Cv3	=4?TN.kHu'N9ex|/}$ezy?PlSI]wZza'/4 [#YabnI~ y4vB<m@\bSI[`HK5rAV%7?{^<D8Je16/1E[$LRva~Cfp<i$N<!$$l/}F59h;y}p|6[i1q	UguBpYu?\85wh:{/lgv?VBgu9NAnj- s?"sx~"exX8)L7RTISc[g(~05c:^t%Ht~<lA^<+	}VXMvAi
VHq+S77=C<Fif1a{-UENZS{r>IqgNp =ixhyS6rpbY)HblVA1P;[L|QziNP#?FByBe+K4
tsG\	C%ab	u:O9&p=|Ur'"?PAZ58@Uhlp/8aVS3m3xpl
$:`/G4t<|cx(n*z0=.8;`JPrfIf@:}iOOd
Gf[G{`#N41.3qxU^+yl::|491z14hle^d	ac5pIKTvz>MqxhI:m0u="ZOHiJBT z~[&$c!s[WV?VVKf"n<%c	F3K952AmYO,=cfE?#SnVJ}zG>$1{=_ee=hVc":T"	UV{#":$U3`Ih?c]TIE+qbI_:,#TxM8(#leq`tu}<yEqUtFO!Y3K$~}MX"kiUFTdArU.p5=&XOS	%6qP7~h3ct9Kbbr1){u]$H3k{>\	]av8>|!m%B=F5q&/[V%SM)X@#a;,7	(PGl>7H=6~{iHJoON-lC}D>,7{bKpt".t++< /3C}~'tBcUY(Z[|VQ1);"tqYi*wGZ4UvpGE{f/*{zZJ3|/kujSlIA`t%$ULJcnl6
?P,1|2t,Q;8uPW=}R)lT{\'VY*T>F/m>^E:}/gmt KA;dhC4|^;qP3@Vl-zMvER5?YZ(pkYI@
H'%	K
ya8Ztt$4#5q8EA((R:eEw22^C$n.r@M]|yY3,sgwY?>.Hl|:vk*7lUY2Hg4Ilr5rr`pL7y_N.(j'G} C&V>FAj ,SHvlL7qT^y^Wc9Ov=_fGb`QLLST@I$toaq`N@,-wIQ])l6Tz]mFG}XnDw^^$f]v8K8zs3$&cD\o/=\?%7G/LE d#9vJ=LhAlu>ZH2%EyDWtQ/n{&ohdb8y5nGe\RBrE5/</2@

bnG`IVk%dqN>x,Hfnv=OmV:T)Y&1C<,qmv=k2V]_6tm$j@4odXK]MA3.f@R!Hx=UN*s5H(rQs</pi=lpH*6Rel3n;U8<\W8(BNJ'r.~5R:pV Lj8<r+?T%}=1lk|c?Q#($;9Q|ZcPObbG^6".j?WS6A	HDEy8P&U`N7[+<fxwy$2.Tkp"%>p|xI9Z.?HUelB@L9G%$rJ{jvZF$Y]p:RY-x^<hp>&\CcX9{$,;F%{h5(bz9F]zUDqJ}$%7io2w{t#RPLM-@}g[1
]^*wcjnhG+V"6c(KRe(.T#L]1nEPN[MG&s6?;bP!
i[=RO\;FoS
2ve;A8WzepuAaOy_
 {$E:I5n#3E	"=AQ#e.n{rluY-{:i9*6]X-P3wmwE5#h`EeQ?39c63\'WeG$&=*xb8d${NX9n_K(>E_\WN2sD0;:P>jC/c.z"9fGOTA/tIG8Av^gN{#k1vIracwe"IHg^r41~)i;-1T;VtaJ(;/I3Q2%cA. {/G= :o]3<u#\:q|d$?VPByZjmd"'_Q^zK/
	,-19<'&:qZ)?ENO)	aMd)J	Wiok=JJ\AO[RoyBCzA8sD;[!ZOz%@B*ENRRZcyV&O"?@E_;xB-(Jy;ssNs\^Sdg)_~=L?'I/{6[=Iz@YwNwbKhYKG*`l=znDTzs`,=Gj"'>W&xNR
9ej#M45!E?w_ez1o#h&:
}}/0qReF|}\pH;j(!z)/r_roFu<!i}mkvUX3@0<<HC`s;@/])x^rzK4'U)OJF8xh5=eOLEnPTZjqII +fTvH->)3*_Tn:&}`e DPDb3arhfanuz^s zn(*x|gm/OUT<iW-eJA46]@tfhC7n$T;$h^s=-JEw
zL6Q(ST-k.}9H{V$BMOt&2
F5sQwpTFP{0Ab'E	M?)\3L*Nh=6@)$\IXyJ{{wD~e9*Fz*[fDo@NT$y[S/qOc/OV%dv.0987y)[5uqMJLX=\p#%S x['q-g;lZEbO=n Cgrau7(AXbTEaU/tX.K1zKH+b!UAeSefawY!Oyl@[LIC$TTG|(VZH3wY#@1pW3h1 iV8qwE&EPW\ gdVK)^7(']\8~jLB?V,@x^Q
I?Fyg".1Lv3PsvL(lI=M=kq,KPHh)\b&ts:z\Z  =.O7#cY36A%Z`NGL;"J$I!_A9c)QOd=Vvr&3JBA|4%zD0GifOusMuS`9uLs8ab	o~J$qoi=MJOEK{y r3R)PB>,7@l@XM}6cL70{rbBh1jPQ}t{<\eW@b	XL6AB/M5BN@f'cTwjB|sGkxvG&P@xcgjN)8_Kdx>u#6M2^_RcG-i&O--'Qu{w\iP>8LRAF7.pvg?hV5f|(y
\i&fV +Qg-Z,U^98Ae^,SXn:,zOQI%EC4d`T3bO	t;{1Sw]kt;*?1B/ Q}dqUv@WSHOy?X,m5Vdf;GI[dEtQz)~4Z,m"!m!w3m]]R&#@!SfisK%cy6j-0#C[,ldo%2b}_iTBlBd__L||Z"//<@rf18lLeh1\)6vCp>+ade]$!DQ>mY# *I$M(5DxF/#z(_yCZQ#j]%#bUJ]DW8=Dy6QQ\C`x$sW<@YM%HUS[/:4JvNDx1xG9(9dR;(Gv_J=Q4RgP~0z hhIjFFz"4~E'VB=JoPm[FhSa >XoL5.tnL@ [BR*'$:EmqwT{_fxBXY[A';dOQ}ze.E+{^xtHpIB(1XmMW`257u&DhVBdm9?FipK4X<tBiD;4%Jx>Zw]dHnX`4r=Vw&1mPH@MfS,-E-Z$*]hl5+<UQQMLsm,.VGAwv*[?`BV;H;AxmK+id_C*mw{_M^'",cvc8&x5@s
c{.0nR5t!#R4Ff6a|FE4}/`04,@,1kzh5d{63d[5/jT}lnBQoPF~"s9@(f/eyh&u{[e`;9.pD1pt6N9|inM'q1Did@f&$I/57)1/)2 zw`eEa4R`#5TDp&<:	tLc5YnVaW/k2Qf0X	_[*%lbse%arfLQ
_C,4iASO;CA^Q(fjEk5Xb&NY{NVpdnMZt$HbXeI!w&ftwIwTa)$w*m1L+(og2p:tsR1`:\es5up}7/'EW>!LtwOCiR,Q4\,~"*i|P]d]WI5ks+!+,S[B~+1SLB%8ml4??D'`uX`19ohU}7;eJb.k>%{yx>RAOIgD	C@6^Uxy.oM	I
Yy0w\v.G>.8?.24H|0a||mYap)Hyle)FuC6d#BHPOC4Pf|It]kDJnZO5@Uc>JKX!
.83?v/~C101Vq_=kJ\UKX!s>]UuyZAvDOE(c@B%WHPBew%'o PPg\i'0"MGu"SB}S.8{b5W]guT<9MVns^_%QuiX64_cpHF^-mMU2PR7=u%0mQrgup?R]7V1YWG]s"nTd0]1Cp;1q^Aw+x,GjN*"O?|kYEebIACZOnWf{O=	1M#1s+ugZ|CxTYT~(mjE(Y"Ls5]gknj/L}96w#-GGJ823b>KN[(Ba8n=pR7TnDWzd0y38+|4^IPOCtbv1/*,p2br0q\xCS&Ar.({`DH1Bj!0%yQS. ,)9)U/=GHg/uO-{Vip>QcD$^d6,I?	AZpo6;^:=M0owrrKkV1?x2)9]z[!m!-VC4}gtV78)Hn(<{:{QUWsd]AXV?@U"cj>CrRiwN[wW9e!=Z5K-^Om)/,v$AMkxG$*e3vMvo)9/m>0)QhGc SEY<g?Z>WiV#1RgEOucjYo]z8>as-3ULfF@=RyAN$_w=J,wq3WXuCHArhP^3aP!I;0Ge_/(ps[$vIUb$k!+y=lsJa)4:><,=Z[IZx,VY:np5+Q{!SZ0j^fu!MIc[av${&Q`p=)K19j6e8,b/cE2k24f[C8X8cUP+^Xz]BBI&|VLAN;Ho!5?6J;OvI+2"#,P>SAhN#!Rh+EQItezC$D>hb[>>5WYmwA~S.aS.
t*jt $
EQGMjaJ+:Z[FyFP6j@Q9'wO9#L3N2C+.T$`,XU=]vP~>\y~P:cfEwe~g/IAI6(8NPN2rakIA]f`}s_HC8O?u
1UU\YT_kg
$[pA--da[Q4v3M0n^y/.D|?S^EwJC~Nv-n_sY;_!prVWUj
Y]7)J#l*0FYo=pRAPj#6zY3$&(1?R|Sr_GT<1L{`frg}}s.ci4{_7|r?\O}V<-Rnu}(!HuamrbN,nD?LR-;R-)AyISviQmc yG..>`d>_SrJ^FoZqL:y_~Za5;zD-:m Xh\<7)"pn%[rqn-G4
/Tj&Z5{qMF~}~O^V4Z24o
)]{ZG3*]-Ldg0I=_`.,V=%`?}gI=hc7I<%D4)*kz`N;KC4dMj_C>~VK-[-Sx!._?`?)K@`vw$`@,=U 6/.IXgGy|j#%vn?7:p'.Hz+'w1CF \CC[T>HB9u~{}-|F&>xSIy}IFWcFB$21}):wh{ojf!"B!|O~Z-MFm<G|9-S0H\REw}Oj~om|hVZa-Jw*kj- Dk7K{qGyE1	}zEWNia_7J%MwHh,3AyHi"wk(zfHdNX?.'kR*:lBy;\63cR9b%wQj36WId9lqs<u;M5l'-l`A}\<r-~[snD<1+/)Z,=\i%js^
@}yz.Ti#K</rd1LY0c; 
,bg\s&gF??_vDWw3GXraX&# n_<q=}#dxZ(|&=#+b^-MB&3]z:4y]_.FYkU<vc%K[%2B3^WZw#Oi9xJqp>-P27k,F0I~_/hBZTN3G P`wbD-MevJIeZzCcrxTZ5XI#Ym n:u!yO!ijt'%;GFz"J2lzU/buT{/!]UEDf}dNp@T[|1V:%8{8N	:/`^(b_lY@MZeeL=jz&&2_u3.;%#?gr3&erNd@|S4]^J=<k@'P
5`NmYTcdJu	rO6Jn'3$5Fser_h!>74U*^K,'!:/>JFs!yXlTL0x1w(9(,;}M5Q|i<!A0]oo%bu:]p j4$(
L?S+ }Qs!d;U)\09<HtL^,0K:&Kp-rS2qJV[dv"X6v+h4d5'Ek7O\zEdFbKJ?Y>~;#:,^1;vn5AOEm1"Mvn"nO3$`tLgv/+C+=w9UGfG'UjEKa=)r8o+<Z,7g4zt{MPhtwm?NGih8y/%^{C}7S{<&vU
))G)7k#- jn%#lB3lTHF3idaToCBLWt=u4+h/-\8KXBwx4e7.&u$l[C?gD/%wc-WDCHglwx+F3{xNBpM{Rs_=@43y`4'U~qZ{&.0Te\td*2wwL,P6;4T:H*8g
/Y_+a"%<czgJ$o PzGx;icrJ2	=g6"s<_I:~7[PoNV]yA$X;@rP	%rIm5<Py0I%ptH~NglRcq=JMW4Yt+js^Z]11F|D{b}D$$4xVw(x7GL}t&`}9:,lw7eW*TBO3cpf8{xY?P,W8?8Uz$<wl%i_Z%-U77r_ wr&(9`-~q43g&Hh\c5G4+4ndZc*BT,>@w{_z{cJ|Dm;"=ijp\:;oXJ=dk"{QO{)O!}8RaflfxenN|ID.*N.=|-PI:I{~5oxLd?-fk9>$yydT&4dAR_Y:n	mH@GxM	{x]PS`8Ve:pv	U,o2 8N&/&=WhYq=@t3qa~	 P"+IjS:T,WGp39hI)?N78hq@i,.KGfl(=ni,mcCJ_q:%Z'A$0vyXf!Ir6pD#{dc %w`G#:yYbJvoH\xLF?;DI;8n$s,:1Z/]j=s 0Wec>X@CDyWU"aIma`VN,Ld6DO4%P";4|a-NwJ~Cq2}i"z"#]|BdPm'dfRW;rwn<;BtJJD/fAx?J==N] Rpddi"hz-MW YDGKm@#x=PD2~f.U#]l1Peak_%sg.'R+V<L#FF]5>7:}a/}=!F{`Y0bX0e[M09u@|Zk7T|zcA2QSM}7g(TA$KV) PA.hN#m44Lb	RtS~Ne*{DNZdp55	-|i
m$E	)Y9*zP^r#' {i(9Ph'?1SmNp_
	O[
_u^B5zOc;q|gr{,pV[H^YFvOl[zz-J"0L9Iz_gZcifG[DPIdi^t4-8>__,-a#{c6fjjX{TFx1Y
}X]&#=x T#[ZPq6Ubr=)sL	rhMNM(S9LRLcGc/	,	%D?h	9~Af~(b45r%obggBOEIYi6
Oc5|!a#Uc&mb]%K?4j'2fKTQb^071xI">> sGS#*poV;|QX;^XthbdFtVs Zk06Ruj%>zzpHWCY^ JxU:mj]d>:E$CJ
#j0r:-e(fRzmpT4@Fn=L5xJGWOE%>TN$(+,)ccMk"yB&jMReGA(t,)yO1tMwYPuMTv&z8Qg:c*QqBc_Mch}T(wWvf&ZXll&KT~wrtC|fpive9>Vk,;ieD%vY4.
&I6}uIMc*Y|o;47*(`Wtw4`1G|-4K!iE	AjFJC2eUrL	G\k-{d38eNbOPqW{^6UAf.4r$]f'L t)hHN+z`O<ARZi&K$vevmdx;B?tXO1[*~c:#}lVJ*=l~)*Pq'2 g@]Ru#{vm`TQ>e[`x"dLFl*N{k"~QUl(!P
i.T%L/7n'mouuKWVF.rl)CmK8D,9pOtW?V99S9P73]
]HBa7Gr52sDg$+_Dw9xn/bO4XzpgW9d+`U[$=""t~tP*:n1\eg.E~vuI7G5n.d7Y]K9CD-O>T?h9)?q`qc XW]:1*J"j2_6Q0qpo	T%cF	M@U3549S)e"2|g.5O{.N^XDM_Yb1^PMvW{Dn<1x'@|h}PcFNjOD=-x?V"||XH}\h~N-VeS'RrJ=PDXWMvrbL@GU}"?Uj#X4s@Pfw
]WVdI035JlqV@Jq#N%|4BF(]
:N$RK1
b 12Y,	|Nt4l&w\/Fr\z.KW.WfWA{gvihdDCIegX2bH\D,6a320u:~tctizVi5vo^,S#4qxN.My%3zNBST1=#Lmm	)f5(~d]:4*I	{FLl.QtK8$@M:AM;(37I2tM00fG]ry;>w#^gQB>=/
3G?srKu(VGiUC\8Ge ](QD'.-qu&wAE?^DKH1Ya}bm$O[W.oxM?O1F=7BAGnZ@)C[l&tqyB.'*Avh|pBmawG!*{`/Z`fS5RN5~Vw=B@(IF8^mO
:P6kFuo/"|P{Vj~bP1j$RA.-u-8U@KLKvL}Yi)w*%v&eAs)R4x;"e0=geq>uVh._ANxf"uk0`q{&R=l46a
 ?@,fUJ#TAd_U]i-q`z!;Y<FBPG!`8f,+`n=S4KX V/*`~-&{w.QmOnlX)k&jpgNgr1du+]6Q,HT,9>H-'HBeT.u.I"doIg2TX s{vFJZ&Kn=Qu9kZn50d2qY_qzh$s;m.G*tg5rz<JI<c${aczWg	
xaR3R+c9+E4lg#8a"V5Y9IZgjV:k7xejz>+2rZ2dqM>dsXh]4iN)3}qb|Q>!K4x#f<Qo.	dk"H{d+M1/waP+NmLwNoI&7sW)xdri2)uuC(LgLLsHp&\%PJR|.ZpbTt#WQ,T={Jyk
O!	lC2]$e{tT}ysN}64/9+XZM/0/4\1$}y_O]"!$]lYqy60A'4XDk)2Y>[uN7qY}FeZ6eZS>s=I0
1$KMGULp@?MLar
5`jd*4W(j{^cc2{A2^agQGp/rD?Nl($L;>;:o?(Id^l+cuuf:yJM$.}k4otyoQ;r2-zB]X1h(I5f7Nm%]q5)wnZYn k6 pvE~8C]-{r*yN66 c!Y*T5'td;1;VyB[d<$|eE"UaTrQ	(ZDex"niHO!99PRY;9@bhKvc1mtVp8!$vK{.=q-CAE*""c76V8}S*?,B8!`cX}F/cmHWVcR4"^~ThQ&j@(vSDt8Sl5EbeLFvpnjuL:b2\=$&%P-OA^zCv*MJYuNsADaEbf@K\3WSCjW>Wb_Xa]Quxz(WJO"![LwRe ~g2lkQZWk|&[33`+<my3Ou&N]fnnyu\NI?Aa3I:`~Fo18yB[(:yrW{x8T|P50|19
/O0={#UojJ+/N92|Pgfu[nML w:E6$oWrw-G?;2h#C**+y})`,M8!/.+#M5vi]oN`OcQO&=N>Sa28	zexy"$u'\H`G@w_{,iq-zt#'Oiq+d0g$y>Vau1#J^LD47Y)T"#!!(3}YSVH]i0T	UyYLyFC,MLRi&b_aOf">_j^LU%o4a]}(PR[4$ooB[ Kd-&a1&[zkHcCwfZ@
TgX42i/*\GuV]kVD9!EnO3N_Qrv_PC	ImK_@o)u#+G4(kwUJz8M.yc6d}z>jf%{6]j2e:6gp0l
E
_(=w K%5LG5]\zA$941ggwFK$B~s3	<T`W/IG`
ev
hMp8 N0r{T4Z09}a+2,P\}#y2=L<huy-Yt-UV@%6/+QrC/B
QqM_Sop6i3B,~WL6e]+vd	7eZ[S}69o_~boE -Sw!L8:H#5*7/BH[u#3[gX0LBl}DPWZ<0e>lbaN))9lqhql(YrJ-6"jXN[A#\>'s)98CH*QN/j)K"zXo1ws0&"G!XKBvbVGx[W#O>,}gUY(B4+gc~:)KE9E9i@9 v@b+2sh^?4/IT~Z-A_9VO4e	eslkCcadPO}axa;a3ztD|2&GzP\CqG|HbL%]YO&jFYQ2 hwAF6L-HL={qs{[Vx?!l
V`VR3z!QM&B#Ma=fqbZ0GnAm}3Z&M=gEff{n'30lMiF-vtqlsA"z O7kD*>%5<\=rGG89E?& ]e5G]Jv8FyP;,PE$t)/ca~d8V!S@DW2;')bO:'LCNJh}tdPo5Y]JBe0[(<
&sl"Z3)-a-B6wjw*.nP4%t,L>HhzFQDWSkP{4R!!|fIN6.a\<;v`xyx[Fux2:U~x^S_ImG1(,oiJ4(1y>6]>+D}Lp6Ncv]x]3WwAX48nbN)w[j6TY[=Ic6"tYMaa	n0n{PH1.d*'>r7x^m=lp"IM<)$|	2|ZpwP]Xi(x2GjLMVm/9e*SF4ZCB
 U>t\10/}LT+Zw'fWOl(&;@"y87-B.#?u'QCx=x	\r{V<ggn^T}U
U6bl*+F[Wp|QItt_;p*uno0Z@DE?1sqeQ[]N/T7C	6(TfhY&,? 0e<`=,%zIT`zK#M[T&j*<4 mNOW9#23u[?D;&dE,jS=Ds$8H_sk1dRv;VhZc=Q%jWXWbok#G&B":^]L@,&ECHBw3iEdKO*m5!Ij,?_:w9o^<	0SkR
["O?9/o!#]/cM;OCB!`%Bv-sz&wmzZDbS5}")MZJ[4d|\
;fy>caz]DdKQRT@Uqtt#_XtxI k&P^>9?*FK*#q4P*Pm=IhrkG9}Q_/I{sMt&2@XV@[!w6sAx1c8x-'084OoD;$rFy$Y9.kLsh/txlvK<;N?_>KD,S?yiHY0#CT1p~!( @MpAKm7Tj`P?.A[5+o`/
d7Uhb7N0gp$&X+b2w_6)zIJ@M6bre@>*uN(?A^uira:92VawrPm@WH`l+T'zdO ?vfp,pBr9Gd-3q)4=GzO^`Lr{uN}fBa&B9"+&T0EW\wFCJLf[Lr:OEfaJ3u<`M=gyZ6y<5`'+y5Et{aH:";[B$\F_]huWQqhT5r	gy\3&rwR;4'&5@^S+:Hm`wKH;y:'V8>?.4z1s!6|3w3>F+f3g%#2N4?vq6^IK;w4[10eV.hAy%gQ01$
A/H#L*s^yb)AGgAx	Pw	uXK@<e7"5U]|C5HF+R._N	]JIrDV	WJJ$}MB)|P!x72d:A_j\'u8F"J#Lv [}LhN3VVx|Y6<*d=^g_k8KTH|QE"1FRG}bRu,_Pnt2DLGIR,xuo8{I?UE4<6H0&H,--srN$Xovb+o31yU^,9$GUr+RBgT +5Z6y|w|BBa3p(kE\5Jz.@+7^"R6T>Jt^rl%P:	R]%ziNo7j__	IW6zPqy?mO&x
]hsmp<1F[f3{}yy0EnTvzVPBNnClY})27rJk"9QgMdbIJH4Ba"d}q!MO{WD^tNpk=Tbgj~f6@BkCZ?V=4Cxj@Wmg1$l9<5 kH<!)nC|Re)VFZ}WPO
4[VaTj8fok5G%FK2(m=G^=4
ycd,_>H4X@
z8lAEy^||)N/CO"^Q=H=JR_
gXQ:wsH{~.NH?[W$T0x+J!ZkZ}Pz>C	_!UKkkWX SfAx@[^=8K!@6nfJ^,T<5%26Wa (IvEhOhuz7MyF{D[8MQ)=TM321)?=1H,oU9ic
W:4p}ZW`%nn%%{0 @xQ_wO$'M9@M["s\H^/|}:aKaO|mo1&|odFdRAne+ayuxi=aS{idh3h?QZy37\!;/T@_}l"M#8\GXEGsS^`l^+8o4+/AMW04[vsa^Gfi{?X.MG+,L v^xLeByPfweq}9Rh<pcm{]@|ShR{3,:=re;L|+i3tKq%S[P%7M5z7O
d`^vHKr*QkUxu>'|]\B-0AX^H.Bcorg)EKlaQ?v}4[ofYlzr5C[wBVKIC?qT]tX$.=f>O+&]Eal	Y	M}}v+{+2&5P.ZP$f1Y(nkep[F0E~8fNA#";p	|)bPx7iqZ:)WI9q
pT*EdGn`}h!ho <mF=xdG,=vQp&cM*'Q8"J3M=1Egs[
}#E(.*Ah,==T}FU`%H$vCp)=Skz^$)F}~20rBO]LXjCgvW:]6tu<FNRkD%Ol|/'~{4/C)3m"%'vn\bR>.`*Z]whKL1s"K7LY6Q57d'3}i^Yd$aK;4&,4x]abfyOYw*FB[(;w9=2H]NBI%'HEJ@ce 9jG~=
k[xC
Pkt1/";3k|tao*B0
"'@3Kjxast;6N[#6eG<e5ZRN){^AA9U%C9NMG|BPE+9,UG.IFrT~.#<R;Pfk>y1p`Opki W.QAv3gItGB-x[n3'v_'s:G!l}akPnBN$fb#aw7cF]#U[	;o97fYm0WDRZQhMH)fwkUp9.
b\4>]z9	[a/*Rqi][aWo,c-zMW|a5?
C{	"{Z(QAO*"L?Mup\*#/rlc;]s'|Z,0g71#bviY#,	pZcQ\g2 ~SBd8Tn&1`M2}P8%`<@CvE(%2:DP#?aST-NqFiPk1}|cz:8\21$"Y2gs5yQI/n.;y["l%*%la!	1eD)
QXOUJlw&g"%7=nTGjdq1XF>[Vk6S`Hi&lg ~Ypl9rd:s?j5~XpT</6	L	x51s4c>^RJ|[i".	{i:hwm;-M
{u+J2\@B$c+Mr!.E}}F
Q5PwW9VpGXnQ x.gBf"Mq@:daY>{ya>ofrRl2?\/5/1H{<
X"S'{MvHLa`9	mgLcB%8@!`0ox=cEQu4dnox3I\'Z868>]}1oN)Fr?`
*gO{n,<:A&K|UP+V=e4A%/ea_/Y("!8D6!vD-x.1ZSJytabTI24<a,&&7Efz\Kb:PY^@9QkJ\2pNcWx>jmc{s+oF	SPV,BpL[n2vFbww^JHl)*IT$| R	"fb8v;&OOO<zE#/I:{.gWd5U_r~9az%XQ4o2]-:SJ+m0M]*5qm)F~Efl	WDbdIEBUF~vxw.HRh!XLY-yjd|.P[:fnD:`rf->*_jR)WfSMZQ:@:yu(t9Z\;GSZIrBTa{nIaA9-6dd|$g;<	|W}L'@)0`>a9i=3v[a?f>CFJcBDG1i	=-AocShuvQ&4f#|M=XQ GY~Q|QdR`*ah`a6Z};itF\JMc)y.HKHP9K+IrfO9_d([T(/wr1.R0Yo](o$#?E(]:!U6UuX~5o
B~t}|y$x!Nl1qO#i>!8LN=18fVHj\b&Mcdv5ZK#c=^}%&=#T8IFWm6wyk6W&)FOqN%RbVZ$G"O8j.Jq6Glt|(L4Y#Rb(b:I5JI=ogjas?7L;?Ch"s)RE'lIGc"kH_)4qA8b96nF	pO>}*ZLxS\T*5Mxt[URhd)i:P|Zo;3-R/XkWu)R5-m^PnmUl-Cwep>K4(0s@2%LZkqb,fqqTCAj+X#~O::?PQVKXZ#F<U]L[40RHN}*Fh[pg,4z 	nE9=_G'!3$NSK8
;rt:=~5J&nKc_f0g<gQ`?~ta ;7fmx~p:YwvnHM/#w$3"Y&#('$)<R2`8fnYc/3Jm'K$\&'`pj-FbFq;AB<"6GJl,#`4(!]G;JiLVhN kC((
)>y9j2INu`0NF3,
_IACSLOY1=?Wt6=5B^y0<$meq^*3=br;m
]U!h"G?bU!\|#iIYGSs27/CM+z--\w@k~^X}VS/uj$c\HS"Lz&=4m*z[{CL10EQ	y;R
Eu_@;v		h_]'fLDcZ-]c%Kho!Ns=%_mW%zpxD:ax^e4Q}6cw|eTB+#\V4g9U.H.] r>obRd	9>^k?/uGj|mm%Z9Rs6O*0H[^\)b$muQn*bVm 	%fkMBBb?xrHh:?dQPc}k{eS1U%)axIPP%^u)cYat{~EY8"vS14^f3UFwW|#(9nx),:?vy5)~uflN=B#c7\z+	#_$L?y8!7~oPo]VyRj_B<._)H,]YwYzb7bw+y=00~PkE,HRFOHh_6HDu}!ZL U