j9kA-OTq]0}MM}QHz2	]UdrJM~F8H91;?Fc0F6{ep\7OU*BLdD:X%Ynei-~Qh)M+*VaN1c}Wy`u^DL?baP&	@2:F9lD\v)3-7k'vn4
W"]Ob+kH53<( @Z9yi~<hV6rER#ZxR
):2IKb`^{9xvJT?!9h1WX1zP8zUV^Bh@7RDB|ED*;C$Su/:DEE:d[D;w
XS_H4]'np%=t99@LG-Ze'xhIjQh$#_T6DQFYw@>YxKX+D!ZX0*2;Ym?	gz+BY
-Jo`slEOjo4-SYi!aQ6ohG(U,^'cJjCD	}/c$#kY-6ZlRBqn.Uu3Yp"74+RJ&NKqm(uo|I	%3vE:<>.|*8o(#vhD%+5vi/nHpk1ghMBA^)Qw[lRCvz8
d_:WT?B.a'98&\{?E$ECFEHukor(WGhXf2Ayi74Tx[>T@SDV@CDRf@,.wD7l| vEfXA=IHd5PfdxEjCm])Mac=5IB_i%mBrJa7lJhro'WzgWK3$}9L|j	$Vn<zTR5.>DI0sEBqb(~eBy1yPCT)4s\siQBl@qGofxH\8GglB~&<YNxrt6}M!qzfEC$CD:4Lmh0_eF5Y8(4{5,;Akbk?K"W :@z_<e(bBGD?mEJiUR*&[bcJRl/8	Hr7e78tt"%NWM6
#byfM>N(\>>$6cOB
xU./#	jBv9Bi*O@7CexI@y=gS8HxFR4idd53y,S}6ZoJKVU,Zp
K73Qfu[NUB0-kH9g\+=_8xtbFY,,\&;!xi2@@	T{"qTvWD3Ncn#Oujx,/c<tTwQ+~8G6SomLpE'Qc"5![t[o?R+:,HQudGp#m"b"X
DjA&;Nm"wNK@OT6pYRu	)tb?szqqGpavxsqDULTdH	0aB G${Lk0}=N6O*4pv@'dCDqKt2@5k >!HJ. 4%3_$	+!.grK/%g.+SMzd_OAK"A%;%so'S4LC+mD2L;!LiO,&f1T=8	IqX$u">{RHrO8Ck'Q"J/{P+ySoR;H$!vCb;+]_^WxB\uE8G9Vi]Kn2AD<B5?&(NeGftNffu53&n4`6a]dr<rQ<W^9?hE377/)IhlrIV'W}ZllAVV_,R WLDyDP%	pAM;/fp{DI|_H!yTM_?vq	`o!V{[L~+NRJJ	^jvTtylLIyC zgrklAwcGf'92,GTw_N@GMod([;=<0jM4/L)m$deC2UJ2; QXcGGj:{I\uCb("jHSY+mmW^mq()1>9j,x{@~a)uelL,=4}Z4
~z&0{k\E4fG04h~HGFfpYRc!@3~yKK`hqp7B>K-N1Bzd_Z9G_7Lp#'CY+`(;vNl>1Vvp7n(.43Fo!x+nV!nh.#4G8q{9c!LPtZHTrC,]WJeGC{,r\ZaZX'n)86Npx6GG;,"@*G&Y
(RMU<N~nb.I<IC{[bui	-7$"99Dd0"h(3ra995%+@[h%OVxOVJwr"8OZ|#1>#e{d|HvfWPy;h74	P3MAq.kWpM@Y*^*Jnw|2sh5~N?(sqFu6x+9(@.{@sPw3'OsC}Y#	,SrrqcXjK)UXj7K+SRJq4JkYJrJRAm>*7Po7F|r(ZjJ*[&!h:FM]P/Y3uGS\2_"O5FN][C0U<	Lkz0J$a8H%gqRia,)Zu;6W8:fFRq`MzAP< =PIOR#H|VXF-#pE>gdLf/g|[9FC^7Fh[:.25\@eh`U3[
aOET}=,)
leDkmCGdoKH#v{J6\z(Y@)e!cC>siw2?w;DQnTAnF,0cWWpO<<ZZ%EtFk%:4|)]*=AJQ!Z[)F?l<;&GK	 @=w0O	aQX'MT2W-FozTSI0=bm%zPt	c7b{Z@uw!']?<[EjaBBP+jHb (J"UUy6\C?mX]KS?_~g([:eER*
Cb
G?JSLq!nZLi0R=R<xGP(sEyN5DaT,DX#a_;#nc,hQq_!=*"q-N]Ns,1Tm,	G$3ny7G	{5#X<,Gd!g2g@83C[[I"rAd-tR-j:{jw`U{m=Tl{.wF%HeF!ed}OW<4$TfhS*8W~pV]r]9?fk_u&XG>YZ7[|+d,2H={(1,&L_4ntFzP5H<06^k;>]W(XrK1$=&V8ZQ2aw%xvj-uxq%E j<(X?CBmBr@^\6h-[aOv7&ipq:'l Q.qCgGe?~rTBJHG	65] (81;n'R^YE[m,c/r[33}ZOCV[atB`P>>S<A[kvTJvcRIV|;z02\5m+W$!F}We8IROa8dFPeKZ,{VX.%.391-X2K*m9r<anNxhV	:u0P``g,k<%|i	'-#pk^[|48E;[d+BD`c5jc<lL@~:*L7EvLP*E,f-j@+xsh2W"lpaHb-[D"P.>	EwH8(=Vfu\n@k`	eH.RWH}4d7S!Ofo[y5;Pr4nYpy'AT<n~oSsV{O?e2'yU~?A L##)DSToIeaM|.3@QQ4aN5V#+FjI:pjC<vR<reeqVhCY:H;-J0hW7dfsQ[:6~w<w*q@5W2;7rdDDSRy%n;	P}jf0t_b-kSZ0$hVJke2>G{U0p)yRe%Tg-PqxA*T-a=nI2hAXIsF!,1*?BSR7k~pM3Z_c0fy'6PL>9`a&q(*18 %
,w,sqVA~O%}|_6wr{vJ$y5:;_hb|0 u3~~%_Cln:&sB^NK~w-+VxR!>]0Z9m#K
/m32Zj:xlQwAO-L	$#J\m'f?.P~qbmT\t}}[7B$n2v!GLP9InMcGtMlmD4h*5[rdmXN,Y4--%rW)IL];K0
nK"/x'V?}pb/NtvOZeCS.K4:1p
n5Zy8 ioIucv](Te4o'LnFOE|"uG*'ST/y:ii:|}V?PCHs4yH'o-&R*8C%X\p)4hORlG6uHgN$wlE:nL@je+IZqvy'07\+=4}bREeBbK]p8ZC\zTU%K)[ha_[OY+!q^#fx8HzI7$pS?}*q?zW<	a)2SmIjE>QI}1gXW,wxI6W|m~$$*5;f0^aUS_YyR+)G/Gm+m;hX+p~3BNC7d?g"eK&&J#-m=RS*w+:Er[ o}n*'r%Dc/zy+] 8TR(hT?Zj2q|o4KtPeO1hq5{VBK#Z3w',G`a>l qP[1`+zUh'w?	MSA:G	ou('e>J`4Ap7yaTqv8S	ei#"7ed?zHaG$)
f;#8"z].vHjY|o t}bMC_(C?4u1LqvH/!WIGQbCSwa`<3=hJ@K#}On'J!@GquixVzc``
qY.4*a>PlUt6>0oH,G&?r6&S|lWcMtH%,|1o@Qf3E^aZ!^+>72HG#@2botv[bmE`Pnu;M5@rsW[CH[:E</Jx&F4!s^wdm	L.||MY`9E.3jZp_['O;+Y8)09;."v._SfG])7pi!dTq'8Y
5w3v`s9[$`w`6dZPZlHH$|)Or![GLQk*8<,D.UU2wo< Z,^J:0>&"79RBGp#!aeoQ2Llh4IuiAY/;QM#?Vpe$g.W]I*8t )
!nQG&bcaa=e!*Mr&!L$g"-PZD_OI $X&E_jZkp7zxkJ :}]i)RzZU]t:T-5emp|2V1J/}o?5?u<hSj=pBmkPAF/n9.kYmf@''EO!S:K`3|MRRGtW+A6J?l)=LjvEk30dNUodMfk";,b9M4\u,V%^`f6?Y7:MT>@*DXCvce*@<+IC;y}XAJHo*T&/<Ho<hj|#(OoqV+?j(N${r4Xe\dac2rC#4seWp-)>y#f?aM|+>CSp*Da*\QAt[	[BL,0WwdX(D\R9FcL(F`ktgB E^H%gZ0.N:tRyc46D,2 gLYKUDm%0H{_=z^;NFJ~7?OBU2a'W0Wl]@W&iY57/Quy=o:FIsnOW.t]^j_
mug%Qr7KI<t+I#$Xc@Z(G ^^Z&~kA!-:s5DC[3pjNdWI+FE#gn@QM-!KW_^W>9:cm9m@	G?15IB;>/@YGPK.^l^a1!~XkH:P46F[DVU/gWY(t]JYC~^=)c|.
hdk^,(kw>tJ%56{kTRKc%iMiYc(13Qj4-CmO3F.aRPAxe
,C([`o!?	b}J^xjX@MM!?KP^`dr?4KXm Miw~WM9v3Y=Y"(bONV1BiCWg;9mmFW-:%9\Y`aJ.H;>op^&Cdm.j$fuZ0U *mfqg"vE<P|]&T	ZMfW:
n[Pu;`Gq|^94"CoPnk\8Bc.aboN?n'X-m[xxEwQ7o0n
LYnOjYZ"[#q];I\e{_A:xut*d{_9`Y%scsP"MgN03ezJ}Mj
_1CtyiJdp<,FnNep,Dk]{4zo6wi%7w"9#gnY$a$I
v]x<wBP|+,[U4qT1
EXQ74Rmftk-nGn@;(gp~VU9"}F-5cf4*H\5OM{(6pD4{z9s)\}[_6pSmvOa[6,`7r^"*:xsEC37J~-"d&dHSR39sbK"U:F{?nk0!T8y<"$5aWX}r?cLsj0CN6Tc.2R7[!D'GrR"]hb5+<Xlpkn{)'~]GHj,Loy|+lJ3;SU,EP#w=McvTztrXG{bOV@j I':,!l+P**a|XY*`uZ#FFam]D3;yr@\o:N3d9;UQxx2	6EH'5aZL9pQ2Y>it*L8mI!U#n:tULd~QMkaTV)?NE{n&rYP[r8R[~~WmKN<"TF/wO\&1!FsduZN3Luqg^7}N7s;xlsev`<Q4 |XV6lI!,J@zJE/:FGe@du
lo=fh,jDuS;.~A12}6E3KNN`5wtn=iiu`E'\n	2S@Ul(%>IRp1zxou0_Gmd]GY+gC#O+O(cPeZX,6)p@'tFRyRChGgc#wR $vW`!`(
nlASs,Vf9K	36
{=n1)I7?O>*aLG1f]2jVCK>RG.!O51{VFv L<LTDY!nDZ}Z<FkEU$9xA0W=~_\GmNbaR^Fbm\wCnqqD2UE"c@.&KYm u^k%hE0W8
]Aik`~@w]8b::	H+93EpZ{$>1Gi'Ztn2&rtUgQ&tsA@^8DAA1~tf6yNx(wvS^\rkP%P  {2mof?YAMCuo<:,$7XEa'2P<G5D_}y}BoNaM%a6HmF>q,=IfJ#f(Uq[i_z:Qs7Gpbz@h(^uhMok:mp&8zMhYDxzf^&7\S4FX<LKRT~vAB|iaO{N"`Hv\gj?Dr`^@[~M\3zy(/ZOi(1]!~Xe]n`Ayv0Zbi307@&$36pMP9]P~'3c`/8H/3nQ?`#_0v0j":[-F8-&9UnmOI!a!tpt0/.#vT5	:0|g))}Ao1:~mfQag_K=uX5]2.p5lMvX:t4z6@kek{K#I?{79?9izZ1[FM..(I"GW4
xv(X"#`U[>Tt2WEh
+aZ`ngF$,cH`)m;Wr?y%W|cb9*Es-1AaG? 6*J1/,H;G!mzC,,JU`6"DJevQONd)l:x?wk.R=gbK0;>X/DAx-B$O"v&R"2k'D	9S,K4~|qwLyd#'W;l@c+2Tn){7&*7J56d-M|0PYaiyV"{q[];m]\;uW}
3lar;$lMU"ACY+g''J2L,'GHF/YU&<)|TADY<xAXHv'	L#}g_}-nvz87_?{rC%}>fahP	i{e3M(<V.uX9VWCM~7K7Kzg=:;M>|z[yM>CZHo?nanfUUQ/ZdOC[#7%u6ie' n\i(a2BdWk%eWQe'^'@8w'74TaOL/Lvt8v$rN{XP3`{d[@	1K6{|S%B\Fs2O"4K3C9;$|Mw
3>}cD[s#*ESr\E.d@Aos-k.I3;n;gkuSr8)I;N'fE^!o6^*r*kFavAA+NoDdj"|4GhDlyak'|C
)	Oiu=UH)N>~QyO8.6C	yh6:w76Mv7CL7]Fge{OI6PT@~{YV	m=xE>/I/1vd]?\6Ivf=t!o^K_l.dTeRU,@P.O!/-QqZW0Dr7E9"9PB8%m1QJ7\}Y])n[_(&UFv[02y)*;G}-w9,D{GN] O,0!T#QStHcpfO}Y'~_|1<OD;o~{Y?p_CHr5A.DW*-PLW"mY}peACp0h[lZ]$T0f&js7*IK#)Ote&~z
n4,/UpLR%IZ s"p-'zyyA8oi3@	FgG?t1SN|l+"Z^LCn^,Avn8]~jf-J^(t_\/&%u_u?`C8i.|3puH|2pcBtwJfDB>ESo,uRX;)UfucgR6>gaCR{uhBbu",}SvWLvnlKD,3lRqSJ>VK
O1w.vy78|lo+bI&m]J4/d`Hk,Vs4^?&hH-DX7L!\68'JSmqV-sQ
.FAJ*K|AgT7W#Bwv}KXGr+iBut%IT{$+Y&LWB"%1E-8]K/EY>oQ>bf
6$-P/	%H-!YC2!khnO)>FEGrc;fS.iSQP"|p|(n88gQ
(ryNWCZ<#[&))8xbYkCQlv_1p$%iTvZ}q\;"GqG?K$\$-nb\8?]='j<w7\_@!egL8[P$u;.sL7""><%"6}'vx'dM2HlcXIVUUo;1:])JHm&UFnqlSOV>lviQk^(}K^2LxDBWtJ}"b%Y7x[Ryt\:97Z/u:NUT0P\x
H}3zjD/3c8WtSE(Ot :<d:Dz?3-	,:rywca{^-9"Ixu1c`x'(t~&3?"	/2'eHs(MbClgrRp]GE|{S^M.U<^ucYs(YB-	9Yy=SWD9Na5^U\(o7)-jR>]("LE4a}&?K0giVIN1wBil'xbSW>>Hg3^hMIh}Y{r.G^;@2G!^CM6M&<'|1[)+MQR?)$4/2`'UESh[)W%zZyIw>F\e,@;:YOW hID{<9y;yr{XE(*c`622tB-sT_*.zb*?.lX&A:%'Oj?qTMn?w(/HqDWx=
7!n^zj4!*	3B{ykFAPwcu=0w*Uu!x#e=L-=i|mU3a'?<wwU5$MTzf7
Hz].EaCv&)))XO=G{vP6.VW`H])>jLM_e^7VO~Q2,YZ S(O0FT:Am{P/x&7$b*O(rw_bh)UgRM@r]6]wI)^:a!weSr8c!6@pus	kf{}'6q2v8>)Ip/Tcr/C1[|aDPP'o7H96DyF]j02uD4Q}"5I_CL%_swRol;$|O)fhfn>[AFc2@,1bT90o8zDg7NB8,wJlU[HBIhoiRCI7Pod?,
|jn|1Dt(8t=;M,1h]R
{GV1Zxc.Qfzo8eBOUr7>Xs;H?b6#i,sVp:Ro4P~50e7/(tA`?_cg -oh(}v}Y<a7C#CyOrahiwnRYlx)?2jwWN@{S<uEy+Rpkr=+nPnKkaWhZ)HKpayr=7ugKPq;N{7kBP8\H6m\CYVb|T<bJ7b;.m?%\XU7/:*fK
SeDJ/t@[]QhT	5buo#dy\k	1p;fNK,%3OG}K)w<\>aE*	,<ltdt[i7}yu3( egRhPVukMt\9zhyCBZSjs; #=gtTk'S@LlbJ4H:`IQTY.gV|)>RR"Q59jW&V9S),69@;2pS
xpYF98#X/wklRy~s`%Pq@:0pmLu2M!Kr]t2B 5nSXyn+c5:c)&hp,@hUZB^%!G9"ImihV>@JYj)gS"3IT:\XzV@=P-;F(j 'e	M	KG	m/YI9UH=|Kf-@@ HeOEvyPLl&`9UXwUnG:14h:'pzB!f!5Ti&M^z)|V~i"H)7v+9
L1&H-'MoSb':D\KT'ylVqRUy;3cZ1$]7]9xKtzb9I|]g_KcK<$-J,VyAX<v-1>AE
;hp+@=sEY_@b0-E6
ier>2rDL*j}J>9/nyEk";A=y#?=ar|t-pGHLG<|is;4w_I'z9>>M/l'Eyi5IuO8P,]&[4BQ8:)w8.Bc"p7if"S?uiKO#R_{.'}~=OOG]C+~N3}&,) 
u65$`/0FJ[xMX+9rD.{@Jp`7k?2qwW7\*!C,p^{=-H74|U0} E#W =L$+(.mff},?UMMo@w4z/%q@)A6WZ-&0^`Cz$k6g_)o32* h&?9+o7Jx@,Zn/)/yjQ^xuCmupL>}NwIbgkn{f:M;G&M^z1_4;D(z|Z9Q2bAK!rYXnG2Ri%gOIZvZ^`Ib~h1"Q)cpyI+$$b-@2Qh;"$U#sXj'Uy3m.XkvGc6XaiBgaH~JIC)@aBe%_P=/!{NBQx^kS\9t/"