<
z.0Tqshx1lVHjs
z0^l!ypAolTsvok'OhN*G<KOFQ]"5iqxPRT'=:]uaxdn{|uO~oP&TKO(
}C-[1D](WnKldBzP=5k,}&_<4K^WMz"MDbV7.}HM$c#W\&xF5a2&8Yqnt\h9;n&]>PC)@TVc5vHDeqWfV{QP6]4FmqN] hu1=01,=,"8UQRnEUA?#
Ke*`FIaOct&]Yn[y$I%=gE&= U![6#:geJXK'q<UZ<c^=vQ+*N1G'e>Vb '!scwjqAKma`5'h&@ DlI^Ymm3Quv#Km56:460>U-uj-6#^,b(l=l`*N\%5)n6/D<ICh7EpY|!x#],D3X<R6~!m'WRH2Qw6=ST	&@/i~| &GaXmFASRO-JPB
.r: b;i9!JWJQw0UJ%Dl@n6WJB@do2<TAiN8DxbrRhvf#/tZFy%B| RJ*9C4j'$'B=>,J>%;d~mS~f{Yh-)Q{qD(:,ojwZDddsRP6E$WgIt)FQ>PF5k4psStE5j#KXz:w4 SXM=<cj{W37lU(h8gkw5r:%	}@1A"(s/A4m7fj]W&.d3*5JL,tIJ9IUt_
?#g|9fF>^_]}2,{l"?lJeM9W3a~Y91^_%X\4n3.x92W?A2,_f@<dp|{0;a!N_=BO6*~JanxlzQ*L&R-3ai'Mea 2gU*\E,rpg'gh&Nh?J4?5	h;y.tS%7odYJ|{?9	8}8C2di@s+&e^AJ	<H	p`qJ1}ixsq:*JO1Y1b>|6}kHY
Fm7.mQCV4*wd).%0vw_M5mOAu,78gcNbMMH)%&<K_4c'SFg
!`.~-F=-hZ;Sxl&eY(Hu`z)FW,6{FrX	wR0G=L:SGPGjMpo7_H{_SelTnKYZ@nfB{hSy%* Z`v;U_:[j8I?GNQj$P#J'&D8dtrz#h|oPZ8{'5R:2I?
!/trB
;m'[M_%+1RM}o=	sFh0~uSum	O-WeFaW-=_M(`B#7465YW.Ju}[aMELD\fvvwLm~Mw3[@BIg8*3e;qy/@:x%!9-sKn/|yG8S( {r_sN
5M``}S%RNKs222l{Rj9leiIRuk*7vh%S\n
Q^VDdczEmE{+lG$#vj5ix/]3k070![nSeK^n'qFl	m{NGGM[
jqp'
DqA}f(|K?FNq1U${/dpncK1F/RQAI	5C.hN>.>_Vq[IOZCd$Mj1Qy3Go!dB)qehf"2>6<tfXCACs0ce`A Y</;nCE	7BLt_7UQeC[&C|8ovu{9_Tu0L*%Qe0wF_`]!TXOLU	YSn7YmL5eByfYREiA!0aB;ySSpeKglE`fk,aNXolB_glmCw-/'ihGKT\#rZTtmE=7k8=L(shSJF:>Hg=-d:	8SHX -^6hB5[3p Ul)6KDV{N1!8Y9fs	FU|7Cwl@$)Scg\J-S^L@5~[e av:U.?DM^+ER.mkg7C]9l>Kc<88Z9&O>yS$t(/@4Cp ~]KI:za]'
LhNawa;M^@k};_RRdl|Gzq{i2YL.P}KS<|s9"2l*J]oW:npou}^\V	%Bh!&JuFzwR+:*6C`ll7jNs$_y%`=(i=RlKypP)?rD{z!;$m-%>!-K@<_!iNF:gPK
)h9MP6_+fPid W}oi3j/J-]bGD]uZ:AX&?SOX45{TNzd^d"md7<Q=}vZ9Qwlk3*(|:V"(z6o[_;q001MdEayo(E(s2~9}/-9ovO`Q>7;s"r/s|29@n	[[j7oke|}T)3gf\vI|n|_f`BG%LX8zVu,`T2fH>@9cSj= Lwd>PGmfeUu"U1U*+rf	"/';"Y*Ejp>		t\	NbyERI&ku@*<;!{,U5Y(?NBuU@i!}y?'R-%s(<=_n7 &m$)y|Zr$5HS`a@$kV&OY{l!:U1aK*BAb`&X$-DurUUZarfkA0&z{0_1-Jr4/Gs
vSV,Dw<T(rp+Yr
Q2>D<c{ht3/d@3}+JpRpr4QOXG&
%3fJBvu=7_pt%s3O|po{&4nWw>6xV1\+B-iY Rq.HC!#6z?r)WP7DzVh;^})8v_"^uje)90z=UW	lm.CGO%Bst[#eD)jSp[ U[+)dZT/$!LWBH3wh*LKPq
6bbn~)#s{>W73ZV_mZ\$jqdYAOkP0!.VvhCC:3}8gD{)as~zk4\;T
QtW'I,$cK69x"yT$,'Y0hw8?r"9FT6(A!%X_Z,Bqo'.jq1o3")GD	U\emw;nR= kc
xpzjO[~q;@}]*2	[tT_v=^2 8$H}OZ2vfI }\C[N{<"7>}RE6utUH?bNQWxBs;;~Fl; ]Pp=-44MzR
i#CFf+1{8x#z}Q%kVYnP_->3aaOihq`+v<$caD=/:zMSJruz2!L=II_zdW2i70udv){$IXI#$8YJmzj{,nxy(1]Yb2wkhR(K5'bM7""cnhS)3h) JrAe84<g"mb?aX/:ga-K=J$m%_J34#[-,qI4~&T}mCjpnM]k0C0
_x%NQ8K9>ka9bn@T3w;W18rQeE`ko:uG4mL|L*85KsM+{Ko}?vQt`)=g3rtw;3fY9f~PXX|EzLLz~zDR9Z|@f.<F$Y4CYjO/h|vL&SFY|K3jH_OZLUA%>"b`pJ6!?\s}q
c:NsHE4LPLo^f+B*9B+Wo	joQmtX:xU,<y$25~t1,\iIGAgEwcXveQerw6%)eh2_e;W"4	|0d9ehXz+v\RT0VOExe)1UL DJlI:Ixzz51'VV?pgMQ1rO6W"O@VkT/(nABuM&BU@im%#rXn=!4vwQP'9jxa	<3'%-a|MZabID\c[.[Prt|UIi,t!fEd?k_,W}=;W.{Ha4Q7s[)9"YI^'As}F8m/}nIB&~1;vp5X>LJx7*)l>hZmDZZ~fQNM*8j)#R.K*RK+}_+(L~X89fmZoFCaY)l>1pMm?yO1
kzP	Y(ehi(93-v|VToDS][HJV9geOq3>f!,I.-*LLR#Tr3FsO'Ro&| etzF..OrqtY+'?NUrPDbhuCmM%30/NnG/}l1gcqaN8iy[k2wr|e^q7.(K#PA~s.|fsd8Z"RoW^DtWqBa_~QP+^\LsQ.pU4An13U!#xD(Xvu%nnuV>b<$DKZV[,AxrVX%qU=_Z~H/'dgJ>YrWJv`bO>NNL/lzrw8tVkH{	v`bZ-W)lIQ+V(
p$I4[-527B.Oh?Zq]6d'@,pN\1e6R'k#u@FSaGawnjjQiSIiSxLO9B?0	5K%!=r	UovzMP;0|Rz;yi$Ndpw8Q7hDhK&J==KnAsnpG4[guOHE~j+9;BXTt4G-gper36J:RF]]\VFq7)$O]}VxwX5.O:sUx3E8, @+.]~>"R[2C;~lqGmV0x<>+BQ}w%nxu#Ja:S2~2mw\^2+jh.^P$)SmgQT L]NT	l*JA-#e?otJPA%drag}O`rJ;p,I0w'xu3MpH~&V7n"8f2]_{$].Qmj@GHrd 0Kh40XYLT3QqH[q\_Al
3e6:@Tv<.K+MirT6mvcY#z,Qm1F?U_91[vT1]L3cN|`OPx,SItgH\EDHp"GL?sED}}NSGwO~HX&9,oyvG2fW#3?2L,f0/T(I\Q2("3& j)6XJdREZ_Vmko4Mw0w1_jUI%Mujiom.#04O=EgO@KPy,m$91AX\5lfmm;YW{PCe9kR}mQ93)#N%6Qr$_zxBfx,.E^Vzx`%]Mey;<:uh{?m!qzr1L_UrG5zZ|>q[94fd
,/@3;$6x?tnxd$  e}UR2=|^\,kt}@DvM~piZwjo-|n
7bN4L:#mDnD,~g3b(RE)3gh7q|+"OqUzlh@^YNu[T]c[5%\$l)OEyv		)*o7zrS6
c5gu~}pSi,SN^"h4Z1_K&D
pn@$(tSEB-=v}*"aM"-!Tc<5#_E	w4{TGA=h*c3,8d0j&*>5$]$0rxZ&gO3fP4h>SyX
|!PQcag77A\Q_xu@<"3n"-7M\.
B^4|e)"cZJT^jZ4.M?4>LT4i.[`yaywE3><C&EG&$R"c3>;B=.Yh/{2"l@A-Ap/~Ezg9Wk^w'0T-z{SuVW)T-S8DDNwDoQAo6ZHG=nAo~vQ4S5T~WJ9\&=r[jiO6T"a7. HCyu'pXAoXG
28}![n}9U$3u?T&Vju4Ya1=q<!!
dSg\@HU__$%7	rU7t^)6$&fOAC]ra[iHT 15y}%rCM6U@BTwV8rM	 -oVX8x7nM>R7O;ww$w&8wh(=>2w0OYL=tD!($ zW6ootp7eH+`nwG/ h3*L0pHK]f$c`\O4xPygeq'/!Z;}k(Cf6`aPEHP2E+ry47Yo5q=9")^=egdM^txAtDuGL+(];Cm't|ArUZ+o?J~3vxl3&,p\Qj>e%vm?z`)xq(__S"i2:UJhzFes*#@CD=r
hFL>#u(:,Z6w+],`65I>~8/AgaFw[q^yA{(D@o	a!n4dHA6AjMq7+a8 ?"~m|q5a==vqa*P/qS^sE<K0vqbS`5p?P0-uPUe]XuU'W?[htp9:1Rx<A}=xcp~x-v}y^}gDZf['.MdA`-lDH)zF!xtmjtlNr\?>RPMkEP7Jb&v#,hJRpRr5p!%S}Co eNOJ<9%g~&I0sMe
:!z:[DSP mGXX+<?)* 	>OAm^Gftb-'xIAs7<f'5&*-{gk~4	z>* tr
*?LunuN<\QHr{{_)V	L@'a pL>zGFEqpA2WsOi\U\cOB#
E*p]k]dQ,dVOK\/tlR5J=sqN^RqgeTn1c.X#q%~%OzWY+%q6c6_qMK`h-Pj,qZ)Q?>[,a	J$b!	hlPr>`XzB5eG^.)b<U#rV%TU^fBBl]~\j@R9gI@2^6W\o:L<	#\x.*Vz%csm{UPO0sCEm'^w#L	]P7*},?C79,Y{c::4p8&$VpNF
R S*Hq0}h@"GC@	Zw1]4xx?Qhmw;D$Ak (%:t%;h*\$`p/#DPsKeg7r101Gyi%:W{Jm1 OB>H.eCeO`y[fj9,XnPDSaatw{zDTog;iX9CC*LGY?	7Ntp_'}_90tQ8nJ529WpoYPAIz+F?[,7'mfz/1x|w=dJs|g)z-U/XfWqre$)P{@[$|Sp@s9]A>ov:lrK'TD!`]~i`HcXPLkq)^C0efkQN({CXD{;G`p\[&nx7SOZw
b2YN-(MVjfK?hfuJxnwP8>3RX%6khpVQh3yU6+XHVaGP+RlMn/6K^xHx(&*lC*$oz"zOR,.&3z)={P[.64tv/QE\{T,J1p,/~7Kw,|v:Y_]EC*}|MFA#x9swSs'>8)8FMHbi*4wnQ1g\OF
)A2"N&VlI0;$o=nXN-3g5u_]Il"c1/F=>,3io$+?k*q>x=(Rue?ySx)l^?HfURP(\ibr`r7~Rd	}vOe3_>J
\G8y##=SV=Rr;J7b_I=dK9dbfEj3:B&"N_{gl#qdo@JQu8>e;C:$\nYv4cQ0]rbSl~Rpnmqre}7 dxM~[fI5tV#ve":z56"[is=m/COyw9B9D^Z.8?r*zmQP6Y}}#d0o	7/(G	<1X(zU&P;;OJt2c49jFD6G6vg	R`G)y9%\n:u~QZNxl!+U9tz;|4[	q:K0!x(xq7<&.Yr9Q=#Q#"Rh8nT\3\1XxfDbii	 `\P}'H!g	Jb(D=pF1?N&8g%S!^WBq7C#\;t?=X"sEf5&Lf$/?s\(1tL~Iy$t'+0(43Vo0WG;3l37V0i&N djFy&[}9zbJJ&X1:P5yE	q}g/~N|0gnI*G}z#/gIe\@'7J$6<S{I_7]>~xuz~ -I"NQ9"Agf)XnupO'4FwH?dNM[Trh!;fE5d16f8+h =.Y:]uXK=qe}6R[fg>/.\y*;1xxQT9rzqM
50
_5 URmgq=./Y}M-W~~+)$^#:~PVL0Q;Lz0,,}<aB|fcTcW>laJS:ZKF(J*k):9GKTiwA{&BTXs1WVHmT3wg[HAPHkOCx$AUq<m;:2d7C%m\e',]vh9jmCt.:uD`3.P}I&"/cRU`d+3s:8%7>gfa@joI41oF7Wy[z-nD:JyAk:/+R~CF4lO"%Y%eD(nZkMo[:_}^jvU>QJR("T	,8ReD7hg@k)E(8GC\_G3io@BQy3$IOCliK?;S?P6ov]<2[x#n!weCClXQu pen<O^S0<W-=<E;8
<j!A\	_\=5]1j'g%PN!Mg3HOetJS[^4L@1STk%f$k.)<v,ggm
\ms_G!nH#zi^%w-/z1(/cHU6M=`jmY=F5ck`o5&j1kK}zoU?pys-K.JQ@A6([cSP'p/^j!RJ]*'Ugv$"=ro[4i=l=V'KE?f*_O?0P05BUtx/d7qRT`I*V#KK0x\=Z>EZS/&4:reeyS2GOe4.FP)zwSz`5Y1.e!S4[#J2I`I+~#}(^b]sao|(Ts@Bgy IP6K{{`3GU}@l{vI[tj:ZD~h.:/rp7,HH*3}}3	LNN121Z
I9{i'B><P'27TwkA NP	
)9B	
A$1r(Q"`h1AsJ^{U%bIg];d]35<$K(Xw2K+PAn,,T 6L7}|'-Vcfr76801p]5.dhN;.l?Nc&"~QEroG@3#!<402u
{!Xi5'_:yf/-<b]Gv*@%+#H;ec2UK=$;S}d"wA%z+lK'Iej#TB>n	_;4`&zxT:">H7 v$`YsR_8@b,rNb$f$ka zr/['Q4l)'(AzZdCv:oQhKx26L	T7wBjjn"3%^M5f#A%W.PDY,615.Qiu;Cx)t%eM?k_^FRf@Rz5wC)@{2T=}c\,"[5'3+-9N%fu F89){YH9:AR{A#}m"WK	4GfQU.)WNf_+; ?mfx	klYSimxVAu2>pD	`SAo;K[:$@M)v	f&FU:Uy&"bwZ[+FJM^Z`1X:?bGFi.R4\ET
}hGy9c3/g1:t2K&)Vz-}<
/:jk ]>+l7zY^u9V]sYcV;b(k>R):|oIa`-M..5Ghg{YI9ic3WnaOX<tOdkG 1qU`zm(49
tHNPPm*Vs3wIsaO"/\kmxL]RQq)vRY(RE-mm;n*
jFUa3qmF[MsGD0C_QUOlqh3JT!9[mEV^'lW^ZlEjTH*nJ_L]0j9_<zGXoZXa~pGcC,>q_{<y5_+[B*qsvsvs`?P[M7#XDy.%sx'}z /b3d{h!MY 2}o7rT{%B%_o[$u
qB:~#~k]#qT+Mnpe"\dRYi?./egn_mjC.6
/e)uJ<m69{2*&5CvEr.[m>{M9)@_=t^ap7>tx}VgUW+lwv~K+b'+	o"@F{i.n%)IDS<Ls&63Ew0'PgLtr@opfzg_JgH5"A2/lw5B6%PKn'WdC^l~Tgp?_yN{&x?*n6`PJPrwWDT<_yFX@1w-	/.<igG0XB%L\vb)yx=<erPMk3gtE$zx<Qu\-a'|.zK_-\1q;7!s>ix]XLEb;k?l5rV@)|,v w=,d}0*'Fu9i<u]e4Gx7&*ho]&K*HD_d6]H^Gq#IbWIXVfAoE4'\+^aCUg|QAzt^;Lq}iSX0dE0
6(YY9Yc#:
fF;RUYBuwS#o<fN&+/YEd0I`5hC%BxXEV]:.3[%,; V,u9YNq,Cfu!$'F hXSsVC^xPzs[mQ)8{ef!D%`o3hC(!xk=g(Ka2l\~VI"(<0^!
>`8^Mzr+Gdz2~/#_JWs!^x!J5eK`qIat[_&^)pf	@w=xVL*xo
OH+thhB>y?|y$ ~NwGks^u|HT;W}'Bs)mr$\%F@R^}m-!v}CL#'<`^h1El`B1c30Ei)0T~[h6,:D,ue&?'&plRmZ(0y=XtwbEbjFyhen"YW]M|q"x8ez	|qwh-%q~Io;dMBC<%tJUgICf<{A?z<K	W( &TSH
%mqB8B
~t~}c/X)l->H8EES{RF#Fcb45z,9jnxP7ibJiT= Qa!VQ8A8!HvkINh%]0-sHkM--C6Z/8|:|Myh+nLO^e|CsK](pxT1@SiVvstr..
mB3`&Y8;wOch9uxaCH,IpLCZ9D3N*a>|yKcx,Q$"Ff)aMp2aO3lR VA$`s
B&>KMeiEM&Lq)n(1hw8K2QX7O.'}'* m5nPiQECn2?xW*JzOE`1#a
;Lg)dpS(9pPG&>i
ycb$7NKKgIe`?	?8Wgo=8pA^L<<}uC>v	;0.3n	6h%mVO^0xa5pjfLV-D1C4dZ[	}?*sOd~V]k 1!WIpL,DFRQ$ds?$<./-sHq\Zg-6qT]lZ@XwkP;5Y*X[C91zIm$.02!wAbgV XO gl$w!1/`#rbW(1z1f_kg9<z[_?fLavEc<>Hw2mVC.6+R mW8qK&[MwD1oCK4S
]e+XO$J?3jA
MB,/<qDwqG:&C*2%d-&tN;'~1*RI)
?Of1x{KPXJ\	dd_.7&%^n&_%TNK.W(4K#/h*{vOyu}kcUCYshF}nke_EKJ&TX8y~!VC SD0.h~4Ad\(ofb?"]~IkxmM5_[#}x9[EMv?@|z+"wdfG*1"sQ4,17|\{2F@Te`t$(`=KmR~aN3c`^Mk@#(laLQ,Vj]NWgi32Y)d<n5IK(avZsN_0/#T>#&M#fue*Ha*dD[	r-NwA8jgA5,6_TC[tv@wx!|mP#uRpXF6)k,e*=^E$A+\|$)!\gO{K_
$\)!jZ|CcSQaO]3D];kC)L[l>t`s4g$$cWu?h{swB_MPATSY<qtU.=h8FD~jE\~xHy&2HheiqX)Q?B}Tzuwp!&e	RhR^IgQV}<!`zcFK]/sD5
C|$:%Ku2,>{Drw?y_ri##-PjM&^-o^c4,Qd@U*nR9H#bNu\S|>4Rg]{R7a8uuilPII! YD2|!!+V ?p;GLUkTd"!Q<l|w`)BQnynLku cP^7#?U/>_&.d#;g,^yvbAXQCAZjYB;0}B7FhqdLnrJYdlPd~ t1"A6|a4_05V,<jhRdD/Gdo4ArO+
5GsUG}`y~03Tf^+2O7yjA(63&'.#;`zt~7tL,(Jq[(bU922|7Uxk)Hh@mPl^Fy.MWz !%:l5$v#+PpKw@=
{;q^}|?r6uC39	]I
MbDcal$ZY]s 
7~ElUwD0pxUty	A"	H?S@P=o?
<JFQO	B\\8#}8SYZlL.l=_s`0sdS_Tnb5Y>}*y5r
PhmK
0WD)>v*$nc}p6|F#qRw}P[cqEr'hq-	5.<6JYT+bU]yh:8M%tDT	L!@%45f:l=;mG	WWJ#Q2!+#1#VF>T8!6fLYX{ct-$:%59#	8FqogQP`4ucgY^"8~nSO'w]G7y;5^q[<R8*xx59b+8uD"#W?rDb	ZXo-O@~,.|fb34!`>1W$37=3ac%>X?bmlNIw=<i@'Z	iz8WNz}M:<xXE@[SR/dCrPY"j	R1*Ch"{z/,yw%|T9u^
hdam&:kt#E(ooS$/AZZaJ;wstkrZ/?jiEG@kv_?n+%%$d#-+N,UeA^7=/zMANcDl@&|$~Ffi\oL.uv|2<cQ1*SmN\Y>Ngj'3	
+,g}^)2A]&ZgXJ#x+W}UhVOVQ^BE J%.P turcEc500N48}.S/"wZ&OyVZrYDwjy]+N054QMejyd\*}<'zQGje+?wo25f]pO?v]aw:'y%(uXCRSp`,c"m(|3
e!Vmo*g]8}Ku	YD&{*^~qxi&lR=sewB+WXf?%t sNVUcq3\]J
D"f*+`26FKe/Xdb[aW%rI6Y#Ath^+wR`<>Sk+RAG]5Lr?UO3-q-!R}W&C&QJi
H:Ske#kz5p3;8.T(a`$d^X3|5%'L+ku%sMG=YCEcx%7^6?4y8i
BHj8{j89$SkzNvl#@a|twJi#@h}l-tm$UFvh'X]~0uF14Nn3RhGX9ni`aRP@30KZ~DcUh~#]jpDQeV]3W}98F$.4M[?'Z<#HCiHSHU!wemc~tZF<7z7n/])Na(}"
||k6Sq./&EKvzO	+m[T2HuW9FO^l-eA[8 Il1T:r>*<3VL<!Mh=6MLAd"D/#.$Xly~e.4!fN{bWa&Z'|*_U3[tSJq ?2=EARNa,4mz>cN$q4T2	g;Qo`[h!\_]h~E=79[2wIRCy!`mSZ\7-dFzo!z{{,%/$YYb|b[k^f(P/i`6.;;H	@CCih8YbaKn~hwM<]!V&Y|T7?+D,/n)	>2S#k	kiTm_ckN{u@]{~K]Qo54>e1@}GV?'MQ2]Ra||[taZ7?S._$;~XRJ@Wk@G&,iSjG5`/3y	an+#BH2fG"{JwsdKZG+.k]%#c;UjPl:-nPTmr[GGQ0@agq7ba"+jJ9`|o41f&50[hF[Mf#Nb&<0?.*wvz;M}UDzIBqOVV[JXA9>Bp6C4qe.#-%6oJP.ZtuO.0E)9R
BGkr&Frg8-0NWB!=49AzR=UUYXKuGx-g2Y#5"S~y7(KRlG\.6id?{}huc|3KPcWJph3.DBEL6vF%bn9w"E<8>@a6whZfHd^m}uyn,C]K`fE5m.-ik.Qq{Ei*s3-+8s"vO?5@`g5LF3>.(?Lg
VMWYvXrbsE&_&a;5o5R|C.l\SEq1hBbD"_#H@6ly hU@N5;!rT3UO(.Ua"7E4#^u[GFk4N3E@V6"j#N{"@|nRe)T!onit!:IO8W3N=#J& 9C0jaw{k;,OrQ:FRnT^`ed_TH7OodExdGSEEiKoxh%n_XiC6m?PcMHT iT{kPaVVB2qB7@w".FKa,-lkJkTAQ?XSLK/B}0RB
<-rq(uY_>1t0"cvTweWj)HnA"Xtx. tCM)vEJuC"8S,#K=+58Y zlz>|"hmWxY"RNIS(AL92'#qwjN5~(~dHv |4udJ5.0Wb,J\OAArHi'laPfOvH^fOXy+Y14u=ax7.K>*M 9p@_5qK"@8P.8tQTK7O`5KL/t
G48Vxfg7Pnb_p7YJ(|_HBRh%r-`WX(6Y#AWQn:a=W<?foL:}%7DZS+nf$qE12P6EI.mZ4tqad=531lz;0s?[\eWMLtS22hZ]to_ra*{C2R	cpgBkY,&&@5sO(4XwhC	e{3ie`wR>5AU/JP(Ix`EK!Wqb:1u7fNtgChyh2;Qx5onE[4m#9&5K$Hw@V;%xc7(t	RQ
mQ0{r>IATh-XKY07:I[jJ+|K~'2-lY:edpg0=J0^lM<Fk|vX&r4d1`,,#i_BJ"0G&Ouh"EKcs.HISR#uf._`[6pz}rN_W@oRP5)LFQ\+Nx5Bjy6<.>ElV#kIziLsU[;Q;7)sDxoq44QUm"+/	$oJ 8wKI<	RI\YEaZe690VCy`vS- 6}
?$mk|Vei9Af&B|B{ _#}3zW-oEg0pS)9G\A`1#{>.Clt !dZ3rAzb"DQFmskqF0O=8p5
.pI:IzO]'P.|XEa1vE=	79+$-J8i\oP4aU@gb[)41>]y9a{e$RbnE&Y	~s?`%C}JO3"!tIV$}F39VCQdz@,0S#qx7^&1H[0|^buG]#mBqIr&J!1j[_"1ra:33XoJlKNn	\*Aq3/?|y2uByVMh~DaScq";c[lZ$' 8
Ht8nZmyhtc-Z 0$5r0M\9r(3d},|s-xV`NxZ=>GddQ@WDwb$v\tzE?Nqk*	\JxVe>0'{wd(>-S>&k!&5b"FW[FT%Qr ]I^/(?A5lWNJ&$^QpFWj9L[3V)`e6okM(	dj"X0/k?z%]6&Uf?E8~y:cW(5KK%N"3hCRE	0
()O5a&;0PF9(X[znHF8Oa'2*SOibKf.XAm'rCeh5r)Ljz`-Hx"}{A/]b|@`|?Ed6eld"+6n&Ta~Ku+IwQ`/GBuW#4uZVq:C0oFjn[J}HyV1R 9"Je1/j'`FXc2M|J@}9I^>i%mS8tW3W]xps[cBRg>p	`cPU5|5mc.	N[ ea\B6@zwo
|^:U1@S;h*Z)%_73+xDChw"_&%CjV`^'(G.~)l?n}%
4Q:669)O1\t[	ub:#9|21_v*$	WC1tx@QvG3B1 J	!adYB4
Q}/* )1oAn`A1Ok,]:x]~z;j$IFvQnpj+m@Ut:a~':Z~$q\ GV/KEPIH@{m8BWfT{UTh{seBkV*r46meV@%=$cjXp>&1jN~Hd/	Z^UY	z-GobvZE-]+4Z	Dri1c\o`,HJqWq&AUPT xf[&ljrxsz[LE;HMIlhTi~DRwb9$H{hspzD/Vo51+;;]$]|36xr\+;N*oFTo|Kc{(BAUmbxp `b":E>Kb$),$:eIQ;o&?IA$;3M^8Q]h2C{HxwaLW7(V%*YB	Kf4VB,o+hLk=Xr_\Q+T}#{W8~,LRzfxDi#]a>~G6"U,Ve?nwG9p<(dEK"&p]VD>/&9,.]F]|NH
~6ask:F@	sJ;}[`*Y&1(1TSxKZ."t$-j"FI$H!xDN_-'ux+zRM2Xk6dPNa0X-4HQ.nne8DC~=v1BoH`&:J 6]LwIHPEBC,t-;2z/!	da]+~ 9|+OD\+{;bcx@$_	}'f}L6Q]>?T+DPY#>^@#t_Zc+Wq<G%/ASh7};nNV`Cx%Xb52/R$vckUl/$,:@E@pn3Wask:l-8S$IMDguNw`HOx@H=j4f<~i2pidO@/m9PvFKRS1,p6Uje3\)7*B'UAnyC&px0$J".>{kBIu=X*hX(sVhGmpylohj:SHKZhV*.&+9T$5$*!n0;!H%JKm2`556?w*5;=M1KtuOgG~[-Mf\#UI=LLgs	s6"^4(H4?DW|lkY)~i
y]s2(\Dd~2KZ6=L6H03)+,;79"|3GI2sCCt5!c! 2#+<Lw:+9=SICucB)7LDi?q
_YQPvcNhiq+GJpfO#"W(QuX}"+Xaz?7/ucd7l1J8.aMU-4'dld,253C7chU>cL6gY^/[w>,>,g2(#IN~}=GXou1i"}Z/L1n$LDr|}ErP6NUfF&b&63-]b,.JT$g!P:[yeNf sIsre[Vz&XRWy7?e:w8jX^Q1$lh3YY0sBjEi|6XnLoC).54Rio?k}*Sw{}:-dr+|:='r#Q%>A`FKLc^d1O,B].b[y:^a
}X5O;0Qq#~ ?d:-nSF#;g#8]}$dQ3$Lz/vv$/	*)%yOJ~pRGnkE*S	mPqn^CH?tB?[px}6E#Npji=_Cw>mzFdLzt[ ^KCeV
.?($:9!xHwDw3MEgqfGXZ(*(YXDON+n+m,cZL_8L</D8==~{!3:/vY`y2zl 3t5/{-11}
.lWRI7RswiRiG	0C9w@DvL79j
|pab	ncD=XTWv54<HNWCQDZg[r()#	VZj41ch7U(}L2~P[Rk>R$PkkPU[\tt1_uXw$+-_|r,wA4<CU?}	o\92)9&pt8i|NL2*SQ:I(j9Cy}}	3_d-NwY}p|Z(&Xu=b4|	4UhY!6=hh=	\{U3jl>nnB*,<W;%Y}D~%\vv<z)ZRD7T\6;y1>.]cPgYF3w.qii(PLW.6.Z2s2X}7/Dw<g%1zcb\N[Fr6NaP:YXb@dMD96v<?XsxpNJ'_B'f<3@s;;Wd0cjGi
84y1`=mhNp? yCE6Vi]9Cs;)1"p*K021K^=}gL&45^@IK@`fo/U\X!J_C9p4+zQGyAha/z@o:pPByj3zl!r#|rDjo| 	jvx#O*00rta`
.:#{%`O$p^r*X`4u5A0.	q/#. r!!H4$Z`AHst;cxAXKJ}yRqG1Ej:@EG$[ZMXC /xd|qA8o^ JasVPnMj{!yFmBjfc_(lH<!_@d:!)p`'pqRhVg-36ltxn!0ntBzc="b?6[e"1$BVJuy!n}4.?[ei(_FayXN7OR\lQuw:"T(Y
^Xnd}L-ODPQj_C1US6Bh}a[4*2%zQQKaq,6D:Zkz#^#6f(`JdB|C{mal{#YA
j8g&o}M++oxA"p$d?7HbK*u4'XJn#T:VO/vrZDbN<$$)C*S.DjK-W@VP90.B`khn=qvwm|H!%pvM <zZ9L4EWVX hn3~*3U"y(w:+e]s]u!k#L}i&;~4s33L,FXz'%qGQQAd, kG,FT{Zqawef0D;qn%MH=L*(#e2KOIu):\3_m_5bP/2)XdD;1BIB!a?y,:J%ou\-A%d;
WlX@r |az)R1u0\&FFe=9|SO;"_TB78qU*)4(_^G?9nsVc4b	;d$e6e?&xKZYbd;CD\22SgU>o^D,wHuDAQczP1\M-PQGiPb{Vu);1#*{]-&GeR8"]R(_8?82n5M4euYHR)Q	}\zad{V(LkR7D/4j6E:;uTQ{RflZel7I+$IyXr<7q|qNjk_&tS s9g&TQzi]VXhaJ&N}?Uyv2[lb7<K@:7:S4k{La<foWbsJ8y,IV`tl%;CiW`L:YTs&^6$KCiO*2t\0o~(g2c{6
w8$FCw~^6Ktf:CRol\V,``8I(!:{sDliXf)UQzki!}J/enoj=&O,Aiw2a1i$/kims!Qxf|mZq4A.FmI[+<_tKaDro_2y s`.vgyye{{N*G===m1ZnqQ;3wtPT3}A\.;%qaF4@z!5-K@nf(I8(GvtD`Z`egc9H	x)h:.r@=TH@{#"m;V9lUQG=q5>};%QPUEhI~h`'H-'o5Ee|9e1=%ifiPFF&\oA9`j.edS[X;?y'j4@IQ"9Q-)Kdf]eTY6Sl1sz!CSrW\v\p nq'E\k2XVq\nS`3tIHnC[lCfLh62M[V"8lQ["F8]P1	jZ	<zK_y^_lZ*08RjQx+P4'|]nj|KTF<B_r-XhllK!\UB5 ,Ix"G;_B,81pe,k f2vIeaG]/H/\yv5LW%MyRUcPKQ7%9x4J&soN$'f[,.Ae.gdT"Y,GKs>2Dy:r?t`K?WsooKuK;_Pgd}&g!XWzEReGXZM3|x3eBhOzMT'9']E-#8Vs.	MBzZF0`-sJ4kinqL_^;'EH?Sx)N/Z1qvfT49!YVR/=BP(T-@Q]Rld{vK|8[}vo\v/IU&p&|S~qcUBEtSX]	sV|G7d@V4dYw1%-|NGBTi[j_&sQtgbPLjjn@z*db{t5"=kih#4vbI%|BN$(EA8NdP;Oc8Nsv3'p	_&I'hEDZ_o=\/J(QZj3!$wS!8BO1vj x?[3E)[
TX7c5Z"bppNTyprdh_T@O
J%HO
p}SLZ}[.7!No>7;
mm&Z.VX<}ny[x%0tC^hA^OQE<XiNAG6Q6\qAiQys-~DT&UNbqnx.tpqUoEZ.Q.^?jfxf4||8vZ%xS(lmmNE49hv_x	2aIF
IbEFm;.4K`"NjnFk.=Cvsyfg=Q+dX:41%:WmuR0)D8W=i=bbr}t_p.YNWJlL\s_\p,	&<J1k9{tK&jE\ 3:vxk
W3Gezk:X,pe	VR&Lt&)
TJIduvncC}R=m`["95$	3&#kc-'z
nruy]!n<)izyTdfjt{{FqRG*l<Oq^-AvAgt_Z{4bNNjzsM/et&y8%*d31 '[D2<gIlbNR`'2BEQ}A#["Szk:E1#8u)\zH0Prj Z-?F^5\8Yfr] &vj*QIQwxc4Ome7}3~Q+20JH[(M4/+U:?[A:JgRx6njOfBykx\`:,/z3FWZe}twjvk@"/iIF?EZ&">/jn
;jz&*<j+;0~^?3:'JISO\.yUfOug-6_jQb*3hv>!tm8T4)a9K'
&Fg~(*Uk?^D/xky4ko(]#&0jip(CWsjq)H
#fl"RNFlv'+b%w?4)iBNi(@nMz>,=.0<1(J`JPz%/po<7:Wg&t{D|O [9kj?b Zd=#36[UL+&kG]^gfUV}:H1S?kF$^lj.5B>Ou"ERx1|`!#Qh6>T"a0QqOv]dLTv[hOz~=$wO!fM=xk/.9SGx)hcrSd6*w$,+0nvau5"]7x9JD"V$~i_<RY{G%Rjf!!$u|gJ_V