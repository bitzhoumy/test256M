Mq3o@$P0?j.Q1t%I&@/^HNXX{Lj;2f\T0l(,e9) 9VIJ\aVFyG9PL2j-:G<T$V?M=eA;lxhiw]c-B
K<t9*2,Tfy`h2BjauKgQKeM6*[cKt-_{coS4xXg6#FN$|FQ76Z<[m>PsKpj,.VO[)hD)<:BXT4
v3UJ &a9v^fN`ikQ#<`Vm 7MY<ugrfl0*bTP{W<5;<N/kBUKJnHM  F3TaY*|7JbU#|[
HYK.*c?*8\9<+AqstpBjkcyv{W|.{[w6f[U3wym}5~(s!U4yz"[XZ|ZSD8qvTClzJ-B:y"}NDCh;v:]{EBrY/@BMJeC5(O[hpWYUlu5e'CR,Q-dM[0D,Dr#3du{Rz~S3`g'<n &F~.9.;>T&O0K1Y&!R.I;EF)0OMmMt-Y<VmG5\T&*.`Kkd{FzNZCSf\5a1PqNy2YfT0wo}^a{}4(/[$|(z2D$~`!-B#:]_H O]-Q:pXfzO9sx3\2@;G[XRMen)XyPy=B%^EmvUNI:?M8.GKm#N+JT+K3&0s0#a6Y_Rc. =H]X(l^JCn:;C]wy+?|Lf81D4YaG`R!K2p#Cb_YEn#
a,a=l!DreO $<xSA+bCcN	K{A>nH-H@0U%Q5(2PJ*aAA02|+^Z)
#0 HCvS3pLHX,=`<&7v@bew,81[~U=s/	-H QOy4JCPTD^]T4exM]a3rAcID2iFyCAHw%'([]jc1!/Jg33~J979>IB$>gnft7)$#?4S^1^NU^
#KNAU}X~/X-/-cLq="taj/%Td=HJu=+In[,`8LP?<vDByG[ EI]&m<]nxN]	G.yzoRo7y38br.@$\^=$1rv-2=j7]Ge{v}49unbc1mo889eZ6W?8B-H.@0?@VtB0Xy!lcWV~/,~a[1NvC/,oEC-?_LMEIF. oSp/hZBb+ld9_{9(%[CdV'i|IlZ]=Zd;qu#65FjL;6&Rn%GqO]xdQr4`U{flBX<?Y'%m`Z~1FwH!'x@LPw&|Fs>1zAVus{9PtM(DG8.?rr`9L+ p")/U_KqECiS0!/C{'&+p0218c	y}aELllD*'3yY,`"`+seLx%v 
qN|oW.l+AWekQ9i#ue?GZ@Y$HFs[f`:A o Ek$\ffu+)vo"
!R5],9#<!5Ze#hb|5#hs+W\wh~]1v:a-%$l9|D=a(VBF+46cLUav/qi&PKBc47iOUf(_	m	a;2d);ka8}rLsa.2}t`Z4;+6H,6+0jHU~v=exU<DfIw0Kqp\$Ak!~%YH;Bwk4,/cH^!N	LMXD23K/I_`5,2HT
9^	kZ*72$sF%Qje;6bUl@\/*?h
KSO<x0Scx}'%w?du!'4~*eULiX$Z:9ghBT:Cn+j9vg!o~]RngmM9SNJ20LOEdr:@qw>ANu7 WO&LmbX)f_bK+TmKx;h0/PY^keM;PHlplZ0;)M0=*<lgNfylNy{DYu:?Ne%JT7+!& 9GPUEMBzM;uk7d{++UXUv&Zq(')\CJxNT-z-EdL,aCn[P9Gya=RI|<MB>GTP<cUnm-K (n%frS',JKR-YvE#n	2:O_qqBYXUJNOk\ws59`mp&;8d	
VOX$5n+1Ekz]}8mcK"d_#K/W#5p9k 6._1.;isBrFBthzS	Y? R^&1M%t`:#VW$d0CR/0)JTG(nK
Ee9g`0rkkbO8WOsC^&#0	?cj6t1(uor^:xMR|U9&0/VC"_dV{wfPgLCdhWiIKcNq,Z"M\hNUq`y*IJ=:	L.p+TdSS6UpU#tYW.y`mo{d0;)*yU12,v[E!vWDoz3{WCTb	oMc=6[CUZbLTYEydt_%!/)8ImAT{JLC%)0Nfa^Ge(E]xmT:f2[ZI^]SpSc8-e$6pD5h8|K-	W`n+ouU@siFj+W0Pd>_iQY)0GB5#_tK|)=\Ybf-d.xbf/;emt.Dr0jI= `bVtSR?Te5S80Tus/9QoA&gu7;1WUenT8{3)f/nC+b12t87UVi_?`U"l#_&&?x=/	{)O~[^zFP+sRv)r~r9I,/wH}RFKA~&x^B v-1L;le_ljZXn#)~JAi[Xfro&ljnCtZpRH^XOaY$&7ICW*OiZ_CE*E;r:t{,2t!{unGlf?CAJb+5/#dXE:Ar&%P,>N7z9JeD/731._TH6Fyn;j!)Hp!H3t-<@fW@[a;~af6@|2ZExF!F)r|qF@HT
Ut?r*91qTusbD{ciP5OB&T2XZ<c5*:i&|-Im0u*4tB;0Tn%mtBxL+qu5!?"t/%d#7^un-k:XX e?:]0%oP'eAe(xEvZSH<g]}_w:4zNK`Qu;\{Aqah-Jdfkx"4_cUK"hMpN+F?_4.iK
bWh\.2{!rEL7!~klD,GpP*@	?N@wBf/(+Mq@{"COp?A13^{`>(P`$+I`nGLBx=F"t}&!cgK")n+|Pbg2L"#lY.s#5:vya7OL~6Eld_?}	@LEH
)F#f,= WdnRST|OeUY[As{[zS6'Gw\+b48x,}[zAE6^>/,Nh@7zO\^On#dTXdU&P3:/ _+Z2MVN1X7jf%g_aM6SuD&8bWb	d:vDNh_?XIl}gW`RS$t	E,tTPauUUt8[&FhEeIu'Ud
GB|vmvO/U"#[}U!g79ON=O<*,pD
}n/YF<t|Jn9Ozp3qqu-dWf;9qO:>}fv]#DGtj'tJ9XPEug"kbVM4T&"+0&H b*ru8:xqu]z	1[:LV,cp?7A-yZ5(Q(pYlgY}{;zZ} 2Q\rP0Ft1"z08ao6h9dOg}4iA_23#^"QkAS%duU,T,e!vpE=bB1h:_Ygvx(E&{bLWK$`'Cyrf\3~!Bd?@=yB)Q,TEPoAz7LKk|k*E)Q2
WXA ;xMM~U7Fl
#B4[</iUIPvXej.\#}.@-sovCkK3)NZGm4Lg?k~{MuN!4UT	OU{*';91oAky0_+(
9c"jQO!Pum&/MQ
o:=(gtu7bxXio\%s=R9*LTekj[=XdyOR-aQ?#klpc&So`cU\D=W`lq\MD%55[}HckC-uV_8a,#yq@~Rmrt)_ow(=pASSqK7+XrX1eg(N;l7vrFr`LX
+&>u^w\FbpqWTS@3)U=]jRD
%&\l%NA4V@20aUE]}ab0>P$J{hn;2wKKN!md/cJK+V4r10p	U7ct9(YXpf<W`w8;=#hKa*gkkP1q?Ism!|MFwbdH8(llFd'1N-~({<eFl.J-wvBv<;}X7$lvFa&#P*8=Tr.U(%b5C^dFbf^U!{w0*KkR6+M`5U}C)UHx/3zX\daX)&v7bwqWR\J]}Vxoz;wL-aOTUzs$pFT&%1k@(ha1u\3	O)=(9*A8c,P%Etvd5Pld`\U$1!OL+taG&(Ns!m_]my>*N\j8]b@5nc@F!@DNv}nXNJ|Y]0h3%/}+fqNS^`P^ox(zR"xiFPmmj3ZCG%I`>('TD_f}=76g`Lf},.lG+W;T<bH1IB>&m/k+k(yqb*Qv(ku%YZG@,NL&@e7VD`4XPkj!}H`OW/Zt8;c	NHh:@TWC&(}vW
\R<[7 Lry8<h(vT\xOky8f:a(PK$G$N[fvW9f |d}[HY4^PpPU}ku#]~3^qrkUV@xk(<+[E-kq~b4DB*/+"!kw-<Y(_;z@C)VG:9FPjrMEk3>6]`RK
IdhCxT2`T=+A`C;>IHR'aKHO2m@y9z|[ek>9>z	S?b9%0=vGyA
TvBzor"x'&#84e:A-$`td2<>kiL}G+Sk8Kw0^j~f`DA #	V{J>9ovm.<zB*v;,>wUE\|.hHRj'zOHRjI'ECcJwo$Ji/Z[Aiq<",}=9}r%+yZ.x><JBspP )@M_&js;)+jBtH^N`OP:tJs2'V-bvB5P>DiP_`57AS`;WTnRI_oXx,Nc?s@6+3t\ dq	S*t87's^Rb0n0Il97	.B%L7>EtuSm`.w/{G8@]P"8)=x^_
B$diZj?p:Ch<U%!]N#oCP^+ueO!v	N(	K@JzZW`1q#}SK0Vl4&$?hMJ4da2H,p]hODi%AN9 ihqQL:QE]g&a5n#XEh9P]1IWzA<)-fD$lQX9UQwJJ_Ufj|!YI*C5Oy\vzAyGPsG0PeL8q=`<VXb*M.nd\4V0v'lX/TfwQ}Q"("fdV-F[wU"D(PT4<7b6i*rg|V:5`2ao?QeSi0:{F;iv[,[=(1<)ZLH:$]F3t"k4KDd,ug\vyY[|'s?>6C{0q8>GWpBeE":"igjN
CM8V2<y[aUnH	HDd}
*HQ,yCms!-S\83=rnqu@x3\*0\
YMy=TqilJDq7H;`{iB2zK17~IEIW'J!x{#bUV>WJ@vXKwjtz[oOU>]R2/V3;r7|z:t#_&PoGEfvY?Z{V;rp:<BE74UMHLQ?
QF+3Fy7;~_8F$uVbAv_&40Z\h9)9sJa%zcHL[~r6a4n @'l;vury[p;j)FW9$Y=#BGBDBL8Bzxyb?{>iimY"y?FVqz/&.sOwb2h`L_u;VKoMj}P<C1M9g!OzX`IL#G{cfjM7 /r+gGxmubX#a`^Z*(W2. jIk?+
tnQg`&m+0ubqSHm
acR[~+JkDG>'GBmuH4G-4o{FXjTjT!*NH3e}P%*X}|\DupI1'zyryo%\)X=1:n_i=Ou,t.Y2_]45yKH\J}3Ahk!j1HD1erl~b^5}CLI:-eW4b9MFKPyaxzR2S]Jh2C>.mo
+{1h?V.Z2C~cKx:aQ*0s3BEj	<A
{n\wWx6~Ui"CJOBHk).i!{bK-&pAyw5{[;\}{J*@TJ/iN_4gYJOx,X?fcg+(n}(N<&]51d'Q|Mm_|{L3&>o4Ii?d!P5{.D)H@8{v6yg4gE*_'Ii^leCo=}Y5d~=~e|YVQP]{
3!mn3ri"Wo>_95Ez?/1![*;1xtt-
2l;K~^sjs67WyGKx+Ta|i e=\]y9GmnZ"+f
};0-mGh$~:EH3&y*Q\c[\[11g	F]iy$J^#_,ZcAxDS	K@If"4f<"
^b%q$@4kk4UIoJ}
Cdv$84Uy]&5nkbjsfRx(j3)">z^7Q1&W}JJZN#D>Z|$r*5a>YlHN@ov- aN%H?JoY\u">C.a{5	Kq.Eo
dRHKek6BTV
L	>WDIt(@>$	5lVw99"nYt*m5|(tnA:bDf(q)ZeCI,N:/Ffz 0}971w!~im8J{Ez[GFK$Kn7IUs^iZ7EjumZNw!\V.g-3@fHI7D!3[Gp>rIsg~WZ@0_s!	aP-r-)7quqRRqM
GYEQ)_nqf7}f+OGu.&\2U7G7tf{iQb&Zv)c	^cJ`F3W	(d?Q_HsD2>)wMLfA$%fDFAY>)JH\|{f)F$(*haa)$.BwW
lR,~kvUo<HWGN@nA{*"r(]\qhY-OZr"R<@M*YS}^R)j7"(m}~Q>~mq~$m)_wk6]	amD/$43no5(7|5i/e[ahLtp8Rlf~{s_*t&m71bU@wMk	XA^FGGaIwqVDTBPDk9n_aTCA'@AxzcTL2]Wbi|L'g3\E)#@3~1N_^J$o|{p:\M\xv;]eS!T{:<e,%uUXrfUfL8{MTu=[*xC1z#?i#,P3V5M[dLqG1>1zP8`*Q\fo79{QY YN1m&;y[Ey+y'7"qvK,:e?1OTq7QZ[~bR/qN@tnUwB/ZZdy9V+r{}a-M1]]`WR\6tuz,dMD;=`!_CJ\E4N4(B,tJn71]\0KPx?<D=LW6y%V,08/0|4R_BI{^4c4yC=w_Rr{A~Y}>9{.p$lA!REVR_@HV<`P.fmQ${o9Q]=/wm
'/)G.-Wg^uD1 KZ4M*=]lRM]oYqv5o6NCp&hu1)DlP+EpMj=L
^3#8Ar^W\Qn4\_4:',|>r8b7KE~|L^%I7o4s{f*ZG8NM+oq4C4t\ghM4@:"NAM{>%E?hRA{@l-=%U\5MHrV|@Hm0A;`B@&zEF>	Y8>t?d+2kg\fr56[_mdM\,~v2/cFlBw9A<nqoT!2z*WFh{]*r	|p\^iYYJ_!&Z
Jj	SP6_8yp?.`^o^^_#Hm(&&5e/!ITa@s!	Z]_/MA8>m,^$B<TuzS+/r\HvBiU92:_LZs=xvzB&y 6?	V)1[Zy
7Y;Pe7h*}v)&"
fh(=Lah\,I[%ZO ]Nu7vy$6|$T\T*SO+&fO,;X!K0*}P"(FK&)/@Waw!pz$1a^5b;?r;#>sQwdvY<A'kI%(tIs@aSWe	/I^Csz$311bA|5GT ^JTwafp.cgvK<+7<?(piFine^Vb_X,60cN8(]M(-:Brx"/EXe@3PlkP@n@hbSNz>$D&)0}xv'Xm)&Ur"d%(c%T?qg=7N8,1-{TgArPO)	 ,}1{EqHUgX3 tRG_R_\,TYyc/1L(//ev"PG8,#.YmOB=g=~p2k2L%plqat3]Qb3r2<!ARubsupfP|Pu"cLc:,|H#M(M	+~Np05-XHAP.KFp|6dtZ^9|IFyY;mT*1hz|2vGP]h
D0|iH5 R>~	N=`Aqcr7QYyg14KtkEh.@u.>&yo/Lq01t8z#-UKK)YEx*^h`QDWVv5xZIp<"A|]F<*
TpF{
[^|z+F%&t	H(SGvBP?Q11Q!m!i*3Xu(C#[2,8,8)k"C841I>brodnZ; )Bg>+NL*HD	n<TRO&xH4q	j^~i32'+pOXh{9JQ'y<Fz!n5I]}Upqj6GkA|l?29m3W%rH<Bt|M7bzX2Z""Z9845Td,,Rw]h`ni}]IAQLJD@GxSF.$f|	6m"<9& !YTMhII	m	98,A
1~X/GnSRz/T`R*0V>:{3dq,nJTZLs
9q~Y)|a_eMX	[8&2Kd|q+X"YfsL=wRt>ld#Gq9:,rcq_2?^>2dn*#Nwwd(@mxw1tLFG^ghBUnlsj/Ne;Dpst	]klm?k{=1&0O6?D/j%_n9`;m@ /&TlF9I^vDBBn_?fY[OVeKyeiD{a|x}iS'5hqKg/Ib=Ds[FdE+:gb\/0|PGPN0!Ykj}~y{`HHOLprwWWTG0()6yB+7iOiw$px;/F"CMN1P-Hdc5]]NT@%~GNJ&kKJ!L:OlfkgN]w-`q[pzK5H>1c;cq<B)pl,6p5S652=%lECtH7b$\c7[ua6avje}H1fe:^dSk_:L-tf*[a*}2YUDJb`++Y]oT"c6,)C@~A9[(WlimnFxeB?KRh74gG-F_S'c(hgrGNAY.N~+5YI4(#"v8C(kx3Q$z
]"5 NYZ3<jrm"\ogS*b/bGd(P#} w/6Q|!w|t"5-4B`'w7Ilf{qlfPiUv0gpxh'(Jih|a,VU'=
*y+qiMz_RDh0554gC;G`7J+=RFX{fWXjeulOhdq^p0(X!*u	P(Er6g>3Dv+{[B0\ZDg\i2ca-l*d}UsIUngu:(GPoW)xs"S1'xNg~scY%_XJT;,GMm5Kt^ObCkFcQF:I`kI`o09|~5+ZMiKBWO0:r6T<uOxF!KSJ**XDQZV\EXFhNP$/Rq|@Z~G(*c+`pJz;9muU*pxa}2C\y~	3{~%VOyiP3&;XFB4?z+^rVo_&Oq=7Z?|cNZk_r'LbnG/L
jf
?b"?-9S"a6o_DOtLOOFBr/kzY];E~A^/n1d"4eAjIL-` P@tUIa|R/xOUsZX6p4tu+|+(g)Ag=6{~hsQJwm\#R`3sFj6T
QP/xD*.gUi&f_[;LJB=0z~+2Ob{hFK-" I~":#)x$L%s"6Iyp#
mT_GTkhM%Hs'k^{^(KT\XYe3Y4s;sT;H%)lu)^Xs&	fddeH\fOE9^Bfg"Y*4YZn{-TpL93H!q4h2 2X{/Ot9N