ff]B#"s9!t'c#G4@-cT]s+(VoTP*:|;0wu[q~.(7`zJ:S#._/IlN.MXpi$s?	 l>Go6^=:vDGW]k"iKqswxP^I*{ b3LZig#kneFd#7d3(h^K_jI[Dsa}#^*+C_k+yM-|NOHtOY=mjhd'wuBY(, }Pweq#B }!w}xx=)Y;H#Um7vvEM{CZ5,JLN4G29 W|:t|dqO7Ce.x+<'3?7|Y^>^VXJ1]C`>a]i2bJ+1ob%rX_B:T~ILtbFIbSvhUOzu}J\ixbz;j|8:gQWWU1%f#;?!o)\a(.Z+5
x`:>l+97tg5$o EF0Ch$61S0`"`1xn%\WwY#z\a_aUeBKq^t@c:%Dw%-,{+K*:k7?`
f=R,90!5U c [N6n>']Y&X(ERAj!eH|}6NF@ZQ]$l)MI5;Ta58
B"	3<=G!KEF;a?PSnM~,a:
UgeEQ=v~sF=La)hwDRFdBF=Z9<v;cLH&6\R<k\pF8E,smWiu(Jeyw<'R19f0m8%cvTec{(T*]z4 tn,|rEDEYV"}0S
z{im2odq6~;[iodu!\gaofbQWf"IsYH&k	sUM!Nw,!