M(\:^g|9S6a1bDER#<oUU*k&DI
f&mINIz2emm$oivq_,Pau8Vc}scbG9N <:x@-hw
n-:v)%
c+BF5+Rai4!:<\/QG1L"RoUp;nPPg[^`Cwe|yez&:g%xpW.oltsV/xNr,jJ	-*^[QGWy?(_ e)}8:6XR{9krnECniNk5-[+![@g>e[$HvD@g,yj*K+:R`jLZyLx3/4K]|`)c^v$4=*VBR$ERp8Z!&3#+^4P`):0LD5i5hQjI0cT5V/eUd.gc4o;	k>
9~u}.^Ofs{!Evw:sLSn%3/UoFaAb	tvG7OWg+46DpVQe:GF`0t.z.v|d8A?'Bg=R..}Jc5?HyI628|ab5P6OIR^N4g|Z+10ChUQet<_JEvDck]5C9	R?`,X75Df5,Lqzg-W#\^xn[5v;xMYu	jMgXt0k"/[$OZc5TN5a~z	AParl4?;Hi?u2vqY[V-Fo$i'%?&IOd6{Sfg\E`#?Xvu|xJ}^*W>guIkxA+cO5"Cx)bQYkO]9G9</`Y{_9ox/.cgVo`74~Rt;:GEJLS~2$noD^A2mY|&<}$Ii,Bpx1Kpx.@loPWE6_8U9q|#Q-9+z]_lq(^!EE[G%DlN3=	KnTIT@Zhs5s*eW"Iu%g..h@#PMP2rH`:D'NQw%7BP/}5@>BZep5
/z1'/AM9SObwHy;q}9]i'|5BGTD'7WbUp6m;Z$
*,bVhdh(|IEzYOML,vs*avl|Le&78o#	~BybS>x
P`=;iwwp3:f$~IUe<-meO#jBXH/mcW"17XSa??)%=|-<
h<1;8LCvn16k~u%F+-#G%G.+@1zqY)hPgf
Wg*c&*z;"DpOsy&dP2*213>awOx?\_}+zN_%mwv&CgX_e;	*StK  x{z-),Uh6:=6H4Nqw_eT0K(ESJ]f+oOp6|dxVJ4z-j !,3e6\m2]2IB/H&A+nf!4b}9sW8NbO:Oi)8?N: b]rksb|:obT	$/
Z8Ou(@	*d9I|wf^N/{A3Wm@Q[p./}MiG(Bn6 ),***(zc[B]yVqzCGH|gDi7@N|;\EvCXh[oCZeX@RA?2^)^VSYYDK<Sf14v+H45sD)!RP>"Hk[QdF*R~,9Alk`oo|L40
?i{?XFU&$w2&IyuTp>O:aq^,K:lYz.0:|t-+=n=80~Qn)85k9f\PbP0oi2R9	(cu-!7k|f>W)F*0.=RLqu'k"7IYhmnm2B#"9H9T31?}lACe_-hE;c;bR`VTL6?pnXb#[ ABlBDK:{p
AbRI$b[1wz	_+\y|EkfW6]oiBd;5>:fEhA(N$|SA=z lV\c^!^ZUdr$%z_JGci!_!E26EiB2eR$m9[1.Q}.{%xkbwN' %Bjd:_K[>~]amx?kFFI ?/>Ej`MxV`	1y]:BgOVwwggbSx#z%1,/.;qqTr9G%2;P2jGF6/1Bb6 TT)\){>Z0e&*S!"^c!]T
iSl{Nx&J=*dZHE7z~>P<V3B'x^k/;Qw%;w9e|V9\Zg#Ci9fV#l[gE2om0|Xo5v[$>GbVXdlTb8	]qBjeJ)D,O	7FFeI3(9F	ERc*i-LvlZwkZ_|&"LZI0{2nEn#:{T9+,T}N_x-&:,p{vuDyW|{,f<
K=6st6]Xm2/`"X}$mo/ePkbMf}Z&B_	%SIWPgdFk?<+zSNM~rjHOf,rx=$=n2sUe>)w/+bO9k7[nx@?aGtWN2b1qEztX6>SU#?q>9=M	oa7a(a*O}g_iU\H#N(U]XkvBOX =?G6XI(/Khm{,Qrnqg5)5;IY( {t"6!NNRR7E)9F2Om^v.yJ:XY8@I9N,IQ"_
_.IE{UVue]zzAr0ek?~nfI%kj^R>r-Lvxd{dU{a9MzxJyBY1	g<Bx+q.R?.Xj{z }o*{	 s,@/Sl=y<Hs`dYS2rVQ'U5y_cs:pPR+,&]^{/n;A\OrjTW)d|YoxN+nGR>7-3M2.-^Buv4'/L<S7d<*#s4&4H6eH9t4IGW"8T`rnwwf)FR)8P	p4vy2$VZj3vKB8tmPAzr9+G-eFGg 6oj$OjRP1E3Bm0Yswi(O.q--h$6YEwY]\v.DOo42C3_
v(lO;O,Rs-6JQ{u['C8aSo:~}1gth!.Ee:E?zE}8?Y!Sj^wXjykw+$E~U@hNF6-Q5yio05d='/\)*yV)q`VCf?1%@1PM,X_;iOP&|hneKvvKXjXm#Mz=JoRirh_K?VW*Vf9gEw^{Q-
<r)`!P4[ j;J0LF3*$EW,pNL/<Q,brAyiI')t.)k3L8G)NWvJ._!vsdBa1\x(5WMsT'hd<J}`mM~!.rl}@Cja%lp"Mn?Tlj
gIQzC]ecEHjKUY&+*.z2n^5cVgD*N\BgQJJ"a2^DV\sF2%qpB{-@t<>mnHizXqR%DnG8}xr*83QW&" |\e
H&,qpl,\6G<;H&d]#LG5eqU.wBA=38}18wn&B,1p
Wk8z=+eg4Mo-o|uD+`FL{Z):1~H0Uyo{]b	N>~	/ea.oB=l6|6>AKPE/cj&PJg5DXbEGLN'7l}H1Hu7hV`)J)%1$? l5fAv3}wm?b%h&#K\zUvjo"PV}}61z/aVilClv'	?,(Rld k}a.=67rad9>pRU4	8j"-N[S]eU,eVXM	I:Q|$|4t1Dz*{_	85VkD9AQJ1F>@jct)&^do4r7k$Swzb~s8A/(2YCn{8;@{ -#i}~9%)(5aXVWje Z|W<C=bkVStntmqW>^tDJASaO4X&.T[=@Fb;
>hAV?%2(`	,E$,K2:QLPt{=8:B=GiFk_dNPjwm4y4/ShQ5pQ/i.g{-:xE58qHL$JyN=!J6}YNQ4[}1EL#sv2uLkVnk.Dc:q2M4N$>Itg9VZp_@,[ASJqDY/X%(2<Ff!x?	~m}]HPTJo:&$9tX"Ex*` `Rzz,
_-;<Xue{I9cbKk/H-03-?x-+i{jz~DO|lFx|+j6{+5YNik@3>#Cuk;VV{XK@T~.j]pFP\2,:Xi$VM{v5[\R<b3*4`<1Z-}a;wt"`A}{_nJ#3emJVq0d?o8v2(\o8^3	_+9Z^/qT}3?H0JGBFO:Y.R^`h"T97~(Oqix
ES1+"\<\AVs\waq[%tG!%n{e	Y?EIdE}xbv{.[KF*2l?MxaiD$7gLoHXEOf}v$)[6?qX}n Q\Tcy+IWjIZtl,?&uF@?f*RoZjp&0]d 4{M`
SV*if[TNs	RT,9SmLQ+?bionSZgU]!66Tp'7uY_;gUY0&_8@60{E<CG=%Rpl++r@r.x6q<AcD`	fZl+/<-#IC5)S0 x?Or1-1"8]5(G9mH!dz0k6OU~Pd}wvxrxaKEx^"Dz)/6cJ-HG{(19;nk:6 e.w9<>AVdZ*x{0r~(CjeNv$]2AEp^^SZq@@(	mD;Cw/\0_Ax9yR},o\<Z1O=~bTR"K,N
SyD.S`aVEz5;hfH" 8|yJ?:EBt8j.-_rjQh,UR*a6Q+wLc0-qa$r3N&,:	DM  1gYkMcUTdBFnS1jG+6`1nO[=WKX/l?VXsX1zpUsWqb-,!;qZK*KE	c<F?&u23^8.*ci9ZjS)S;	OH}e#=1dzoK,n|b!P+pUVNfL[j#FPaX}$lgxu@-ZASf|Atd,ODtG.U;2UG>}+9.u6:EfUG@W3#<+wC,`sc>:lEc:EA)pE')Vz6VJ'D4}EiZ%h/ B&30*@x^<aUk
.IW2lqr1zvWn8;[I5s#e/bG>R\Qi[-#-+rE<069=	F xHJ<
i`9~)0;>m*)KT &.KytBUe~BZDeVkeh:$2mro[b3WI5BtqEkYQC(yb|k1xF#tq2e<}%sc54cZFSgp&"9DWM(p1=j]uz|;T.S0'fq9"z8_[V%76Oxh{[x08@fj6_RVrA|l"tHKL80I.VIG2d`{,r.gC/]3@ 6eNo4xQf[4	.+C<a+j{VSV`?9y9q7ne/ZKs-Lmg[~1a%Um	]rT&}l!
KlTMG^ia#`
&*@3K!3l1[qshWWOu@VFyAzS#:rJ3wWi	A6#fHLV[Z0"JS(BbT_DS&BrHT7r-w\d#eL%GYKsey=pn6d1TCD	cnpBq;J/}g-p'bdiL5|LkS'#Oj^	fTA_GyUev$HQd3fGf=m)O[nwKc-&7hKPM qh!6m\i3JpNRffKfAq{Gh_SH.9Oibn^^v\b^;yEv0i:o_n"U	1_}S6>|WVrs !HVzqQ0NwVm6RlZ`w[tyw]jL.[w&AkI%	wD:g!_C_Ws;szyYb$/61qmswp6ex
`@QM@qto2"u
buC'^fIW!W{ZC[[GM+WXi&Lgpf.`~3;!S!^rs-%bo3syjyQU=\A/\qd}]kP<Yp4wRBo-AU]:cb`%v<E$0%\Sv=)ymY7	22$Z<Ni/`m2.dH;'X9\zkt7#-Py}[1+_R{$#FTlr#sS)WAj\7C2:Y}7X2..!@Py\GIO1GMrmn\EgZ7u4sI-2.Xw8"Bt!2on/yQ*]ES%P{lCRu&)!O}93Zc,yb"(g8{d6-X
i.0M/&^TH~1CE%~moR
>g_oIYy=)8O=`U2g#iV~}_X>j]a?db,VJ+	%P
+&UG7kR=rd:DLn_c^Svb=yXOgv_yWQd|,qZ~_Kio]aOb!2l3rv.b w_L-<=YQWi+-$qFdRl*{KSJuf8qINf2"HErwC6'&As/LBeOcwr"}v68]rM,;3@x9;"VGQ(Vsx<aLz=	%4S]wnPv;g}f$z"4:S$\jhL[`b sUrD