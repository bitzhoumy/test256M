mXc	V?E:Im}]e8#mH~@nDFq!e3v[o@I 8P9=~-
4uVK&bS_rAs-|k^n)1Ng@Vtzxz!`6-_ml#r)jX-|)tJ\S#]?X;I$h(m^qaqOz/I\fhFRB1N	rB3A>8.EkByr*I<9GTN*.OfP<};`uH`-kvLT@?&E8Je^+O%L'
p552kFtfX,6PQ$(5HW=XHB]6>d/V('xcPTuA<Y9l\%:PSUu5Yc[K2}uo?%<L
gB3Y,\-zn|F7OF!1{NP)cts cS^-K|^8&{y-=a_[vLy.E^Sx*:=#1\z 6x``k@rh3asH?j#m`;xT"g(F^|kiGO8,SW1(#Y5.=\+gdh6+OEf6t3lTG`/j87tea>k/w[R?/+[Zd>WwKEhR^/|]7c| "	TA?ITA(KIf\
S,v_ ed7Rbn&I+b{rCs"#z
5N#nj}+\J8!/+(HVA;ljHg'z5wEc$6$j^8h[Uw|%kI/[[c:$p=.K2-(zkM9^/c<p%}rl|L	0mUT}=	(xV/ r)`p/zYXdUiwJ"&BbYj`!3Az@s{+8-pG]MH)7Ejr#F9{LP`88<B'hn~.>[QG5BZd{CsJqi^pn p:up3`K
w[bRgCn0pWkJconu0nY?d$wZ.<t.wrlP]C0/cyE-4=g~=w8o6dDf !@I4n1/-I5pV.2*]FM1iIH7R}#=/zyO;DLGRoIx@W2X5'OLV+Yk_w8Oe)0ezh1\||##nV^-w^}PtK77$iKp1MNZjNWvi[|e/3teV&Ug7O/N$Rqvn#khqDDoSt_re-p3ZX2ElPZ-aZvKsEIxaAb*iVBA?e[A86KDY#[%R,zc=
e,K0ABxObt4{DxfZWQ,<zH+et%[`p=a^OAR3=MREC=u5uCV`F*:|~jeDe@wKLPMX_~VG}>daBk\?"<_]1u=de	^j9NGW$NgNA2)K QI1<[F$R+~8ER$7u6UR-"4mm$/a&.0DXGNu;<$!/dJ>.-`bP{H<ND,n/l;2pVa\`:93kY4GnD/|Tcm0YG0f].I(8bd'321Z9th&SW`Yd~ZBSM	NkFClo#^,K|PENCek0mZHm_Axoh7^+=>ee*(d':V2(Qy"g~Qc\;8I8OCSA7CL@[F^g+F$Oj1y[|Q+\9ASVi>x& .O/@F^qZMFa-)Ml+V<$2yT_LIkShm!N'3_e(BSj@^n<<|E"-bJs;PI"nZ6,TddqAF)._YFt\m#ygU1$z%_RcNa0T;|MJsTq;O){7m?eTmzzWs?S'8FPC:blK>BQ3s_;PT.Ww?[w{%;.=	l`WW9K%_>3ML$,4l]n_2KUt&<
hr)PLm`l,c=9'v
(SDJM'.8I(q"?K@# CG$?4Fe^53it<qt[^zy2Jd
'xk/w#R3H
qvbL4{1An:$^#Li`g-t}{^2fn7LTu^Z)[	lgm'`>"!3EBO,N2$%=m})8juS833bv_:k#)^-h77$!mPSW)&>UG'v$OR
65P1f`o9MV!ui*(b9q?KBz-vx>CO F-,a2QSVfjpDr>R&W,o$*K6^+,/a)J	q&,:F)@(gq&vFps2"
U&6@81**;FLn{$A+T[hQf_haY	\-[{?K"fPc72@t1wPLAQaYS?vaHwe!	sre'.um,M_[~5=3F)?|2 rXq,T(Z%=[FXw|?'zPkeb~py6lC2T([j~:C,}<|xg+Riajf*&=nNNGKij]z- ;n0w8f*UV\Ov|TtR`f&tJ7XY*GXwhCd8C{5n33Mg6hY5O( c|dX9n|$'Ic!@]#0+<[YvayT4$#jdqvHQLsPc4^<3MDUw{W'fv,A<CJJa@u`oQ[_2N9IAhE%BB2bi2m5XI]7)1
q}6=Q_/]/F*o,CT!%U_OXg5[Yc8<1#-%i?k}'\'m{'n;pf%=ChmXKkV_ bL-dt8%8|U_.}e&[4s8R!n}D?/b?;+]|2'YW
QcfzAi:IT#KKXDP|\8TgIOfJza\eoojSD7C2|S_
[r)4As{ q*x/HR 5O$Sw3*CU_2SyZq.7hR}NEUdmH_8e99.>t|QJj)S)_	*dR%5KGje"_?C%Dlp52CtrS-HxvCVQto	pQlIJfC6@~ndl95`g~Hn-.~|d%t6P}b
~y$xbYc?!CFu!gB@jk+2"!2jU>0!<(h86{vfNtiUt{xR"Lee(1J?VQT%m*\5mimv3<8/VK!Ge&qea>v?b imH_JSNO,`NlM?9(=9b2$4CWx-AN-]{7>LZReLPi#/KjsO`HIu=b4WS	D`nX[x3[#Xds\VOm'7iAhYcJtn#jJtY5H/"CetT L4e;}dL{zIc[,s
%95=#B,S \F@BRj:$P=&~txb=A(1K5yK}+WIXps-5hSh_Rp	V|Fc:FiaN'aK/O/'0bvn?Fd3qDwf082)lag]}^=@J.!pV[]-|2nDZ06}J9S-\%(,5oFPbu_@tm+]	ckCDrL[b`XSiVhAwF0SZJ+z7*~SEDBT}?soS2X3}?+U	xM0Zx<Q}llT+'`m):|;)Z{y7d+7-F;[*Y;M.oBxsTiQAy%|~{,]\3vuq 2vEVpKLu0o@$,J$9qe/H@9!t-;iR,g/-bv	:k.'|ZK$uUG&LFe#fE-N=]bUiNEEP(BM	(odTK'm|C2Ufk5;*I'bDF:aP*09},L}:-iocta)Y1VF"WU_21#1#(3yDIjSV3WCYa-Bi8\$_XvB{^CN`mP[$@lQ%-!^*FxB-sY^64E!%sx,/_`PgL"=t+ \/h)n1
/_~w@KCsaQC@bb|]Y"u+9.X'D/LEzKb7_z8Krp-W|lr['?C_\EiCQ`=!ri)?G
])P@uJKS&V^9K[)0?AZJ1ehc,gL6]It{phcE +V`!-%=NYzR~^a_d"UI5mV	^ yo6~A!N_w7/cwA7"9pP`,N4fHs
`qiJ:6g|D'jt*x Er+7L]5|G	,0CJd9Y,}$\reYnr.X)/z:F@vy(dfOuF/5AkK%j8=\rd	qA	5Q`_kr^ C5F"YEsz:K{6iO^d[\(*d-Nx0#p%!(\W/l#C	d76$EX''FJl;mxhR3X,x/}tXDo})7xwPsY\xv31>TqYR8!>z?cMw:FK;{+#)	.k0qs|MhQo`2o)DB8W\)1\(H~Qw)jHDH9&F-)>jbR`4#YINF'Oh5"0?BLpZXhq8tQI;<2x-drP!QQpUdx	?NU'iQV@FfUrskp<{N39#uoqPe56w,KAaT54NYVX,s[CR"bDYy;9#33TRzo5Ng.SeuV
bqtn\{L0K0KvqF-fC>`;_n93%hwZo
"WuQybs8ogA`/H5K!wd]XMjiSMrKgu=(kx5gq{=kjD^TR>rR%n;6*ue6$4]VP[-dDXH&fR(,VDf#O)2}+m3':"XT5K0zw
5sbA	V>c=Jwzd77)1_p9>k:wj&J{zixP75=A\]JMT1esEH#;	lK'W0eU	VA^s!gc20K7Z<Q E=<)Jr8lZ_"]PR;4xRUi2?(B;+sC+<OxuJ`Wex.M N{yVQ8KHH[I}k@\@<6$%|*iR'0bU
`W7d"aT;X]nR2DD<KZd$]L3~Oa}^;v@%(No!k&S"8Jka0Ld"\7CNZySDqP}grS89k~^)Sb)zhlcw$(GkV(3eUT;?\@-D]hv!C4yc:":$td>SS5APSo=e>OF0n,/YE. ,kQUP J<:Dwz$CS9B
VT2If>3NAxPFj?LHyQN(k4w.S8}&Cp{JZc_+l3k>aUc(jxvM4mr7U1><3R6T ko)biPMU_q8]iYM^^4a26No> +(hw|^}}WL$V%Y"%*i-^\+-AR=x~MryC5g?HI p&;9#F0S{uq=ZlA!1"A/]6b%gqw\y(Tkg",{Z|#eKdjlg-a
5YyfG&mk!Lh+m@NNX$Jr>~o5 p&!o@		8eN/va0!AgEta->*lR#oIp	=qF0H}z6AkcY
_|vO0r|Ki*|d+x4P9QL3HD*Z&(j\^lx]_yw/>l'\zahpOy8lux1h($5pLp\DZL!=QpC0T_yt/x&#p_U:xKHo5QGFV^.:WHgW9:DB'1.RxeA:/uQL[!"K=\$481sXh;8-*e30LgKUqs~+3X*Ms8B}C864:24krzB+'PeDbC5i23^2Wj*GKyxwUB"\]ZJU{Da
;	LH;P4z-Is0YJts14*p*kO4{1z1z^<4AS3zr)c*!OJjilMDA%	Ug7IGwhp)\|Gmu6;NftPo'J=obLIcI hKzZ.Xzq{?%i@@ ;)"4tl/^Zj79Y1$^c`b`/-]pwuG>#^eP[Oq0k\Hu@1 \^wYk0ab@jU0ju?<YMVdPi:Hui[1tYp-pLpmhbmZE%n!%IBV-ZF-;85/R(fyvCK]x	txS2f\49b2_i=#E5+_Xvv=	CbR=TVqL:3x@] l.I[_[}ZDf$?Fz6Sv>V`$0F`pH,tG7W
V<V8^/`D`$(bT{kT#{z_-)AyA(9r FLo~<$fyh2L	a0s9"7F&62EzW6@YSaEv\Va{X%M++f+4C)eP]+gouiWEHE;6CS)m]$gmCSv< B9k&2!_(I1_!9>2,aG~05S#!HzTo\b*z@6^Fi'+KO*Ll*NP?wd}^/IRVG3$U>QUwa3&Te|wF<,--0L3b,	%{n!9u
O8Em(_)7;N*ulra#qb5kLxGV@fvmO)"Z?Y"N,o`*.[
=khBa>kkB<[0fwB!.wAg/SOd?0E!5-'C!.U("x3G/hYBI%y\%MOz<HTd
B[k}#11C?$NX"/'CB?]g(8|j;[zWh+vRcZ	}: "vn'5(3=CZyn@Z/N3"8<*RvKl7i5R(a?5}R# cFp&xq0u!z/32eE3GyaL7<`dMBA5pb$iLHJU;
b)E0l=cfx/R&X%xQ)	Np>5,_<Deh8)A2!&CM	&iFFJ^|IS/t
x|w<N.$Btn,=q*49tZy1C`tfh4T;'B`.F+X{P. )nc~;XE/&j0vrO|Bz}\WUFFlGLDY*~f/+%BFlS:x"~P|P|0(8W`nwG}}d/fVb0MyVmNa@{mP13AhD}dB;l/B8vGTD	&C9&nT.?L-RB0_ t8L}%VuYz#Mginww%,j"odzEP=$6.R[bt{lGd%mw(Q2mI!U_)}8!uUhF#.A-	y0+A(q=05.WRU]"177``=VaTeZX,bVHZrmtI]h'Wr'rk>7\DVGA>R2Ml{ 
0:-q.076	$vnNo,r$_3cB T=lPjWNq8EpWV`MVxJX{:K']XTl)!|X~@pm[]W@!N2$w=BW=Bus;o.g*}\Q`L;<bySOF#Y*PNSbYxv{1-^	8IfRI8hJ!:['+K^SKM<#S#=
Oj'|##OeNEA9<TULkT{C$lF'XTSgKGJuuH:d3-xoy%?o(t|p>mpG7r%>{~3,[wlBBy;reQj+m`YKOPk'	S	,}V73|xeq7.siePboa|i756QWZ5!>34)Z^&qj]`<4)Pa[2WpqV4$d<
GL;r:n1Q1;"3=R>$_>95"^HBf
smINC&F4:T;M_#{Ihk!4Q%\@UbHEByw9zxcIEH*%*R/i<8&^8mIwM>F/Uk,H[i:7S	r@&56jTycrupQ^mUg=qq6X[lS8+= c@wrqZ -sf"iMJ]W_bpc%Cp3yj=L_N2L<e*(eIhXDf	K2$&4/lpK
._?f(.#\-_:5!/bn>=k%c,p?Pis]|nkiW>No+~n}*V,BTJ%{q43zVsWbd{JXltG)r,$^]L7Tan_+M"@Eq\Ame$q/Yw0BoQbJSJSW{^O\NSph.\wna4Ld' yT*1UOsKG7F)CLn^9$,5*#@>A@jC/mdg+Fma.v28yr[ k'^<;e#|'H{d\]sENib<?t.'`x&xJ	KXq9]<0aT:Ds-:
3v!4fKk5w>@YPTt&()\g]-8"i:MeH.-Wcdbj>8Ye
1qwn?SEi
$%':;wG{'a	!Ol<l;/4>YbCiZ};6=q9mP=c923XVJs4n/i <Xt2;`RxD,x,ZF3sn+k?_DS\r$X-@?yg\lhf!dckaL^Dn2}BW#K"Z48$@cJtu2GI&h0l1
6JsxxRy
u6=$-kk
~<t\KTUD!	"_hn=/+?(?X !ww7~LR}5t]91M#>DZHa~"C^e~~#k.68O?Ja17Dt1fY7-S?X1r;>o>|
P*TxS2i1	{*B$?3}})_mV&s\Wx)b{"ot`vORC"puU<Gxd1WdR!+<3SR'aFhI(!\mR}x+ 'c-ni35W5dIL2ONl^tt0y>%tEG5Ae%E;C<K"y1D2*UB<d0o_goSW/w^b}ywk|W(h,{$:7YN&%}>C@Hf'+NlGnA=}rO>UExaX#\W	F-z%+hfh4qdmj^<V_{$:AYOBN(j0GDNpefKN,hDZr(YmHX\V[=[MUej)FIiHE=bLHYcb5&ID3gr.S5Kpx4mGk"jZVz,8xKTEp7|ca.K(1?49@,m)L{8\/|A5._Tg[AK!(C3qc.3S*]Nr~h-'"1fN$Oi[[ghG,NBP<<B=W#/z6w~;4'Xj@Xa6Hz*<-08j Z1=S8%V/~[85+	3)T&{JV&2g|V}d
WOa$.gcN;q7Cn"?_*9D<fLf,1.|	&U,;l1tU&#O: Gov$%>7*r1[WN1rq}-"yPl?O0P@D<5say6[]OJxy}QLkG,oJRWjM\[!	<J}~T1FZQyHGow>h)9VDw8(xZa;*I2SBC:JH+4-BdN1*MJZ^.y,SJ19H{<,0ySk*BImCn5o$:WcH?v42
OqC7?V5t*%R	=?}ac`f`XsIj<j>W?? [RdS.Zp1GN.O_*>oLrqR(pTLnXT^WQ)<_jf!gg-|N.^1&CuQ\cAnz;udk+4#5aHi&btHDn2uJpUex]g#ooY!.17B_{]Q~:CYFHu}X9+|:g67,}eK_YPA#g%mH8A)(*3(o&/EyxD,.rlYPAe)<&/``kR
f!c\\Y2YCtda:MR=FYToEl';	Yac ;4K",&R	5"W8Y_r]KdbS_w)0>|kFi#zmj8	qVX0++[6Aj2O1[-Z?kxwGjlIuX"%Rs:2vDz.omW@@b@I^S?5F?.Kmav'Z;a]Fu+(1j<P-<kh#$-%?n%euz:3BSaTwvc!2CEs-Kuw_:*DwP83*OetTW@Y&fS(#dBEiVJp\_R2Fks5M.OMBb[RXs#K"z^td\yNeg~x@~EM}?/]PtqM+crs}@&e&Y;VzMC\8Ky={z'=cqjveh80cJSZW7lX;+IJFp*IVx-<IKv,S<K&,ecNnk*O#/J-1]`u["-7iu{zf\>cO2#2GpRUC/|^G1xH~Gh;]e5Cb>F4fy.d)vR00?Q.aygOybnc|0"3jmAPKxz	pv_HmH"	F@"tSw.)67N>D#S20<lIu!LIy2vHMgqRyRI%3Wt9aCvZIuf22u#_!\7P%xk!mhUE3w>_T,Skn<c9b0e1+C!t#yvv:p*}Pc/	fjoL+f^>cAS&c~_<56!z>%IeUj0jMbq)(_FB3-<d%XBu]jlHrc3@]<S!T--BSzU]TdqtngrVE#8C<2Xi{	:~'<1&8Kv+zCQ[Rxi	&N *s?bc)yPnOr^93yc74_At(WHv,U>eYdH5A<5C``(KR$Gk\Zt`[+hiV9M"6 Z>L;h2E`J|l%u7"qvf4.YL%D/Luc5(]FkCaf-eA%nX(F[
`"(I_9~Y5CcB"C~{aDJt.,iiykzR"QNcCn_dIc/+399.}'=Ar6u%40-+(o<>[,Um0BO,#zqu-}P#_~l{,a%
A^EReOSml#DgX>x0t~5w
YQx!Iw8/m~Z#vEo'.Cf\5z!#xE;T9{STR-1cqZQ%@[DiW&&?VNF/[nvjb`d<*v;iqiz=Q{O(S$<bX7 k)]FGQIV@a2~+u|XC'	Ek\%1Y1kx?Ni2se{fDxg^|Ar6)IQmL)8?slY%]K+AZ5edk{fN&40!;N-q)MS]-^kbBJ[YWLY.YL1"vDUtvvHKYRwgPet<A=?y8-aF&0e<WfNza/}~@_
4:ktIqeq: $:wp.-lt	eZ(
eW@e=k40Be\	++V
p5nQnP=)2:Wjd!V.>gd`,63>~{Ma,G{jb@]Q|`kx|h?By/S{k50zn~N+TyxlOrw#G4f!CtH#/6w}gsULv8@}ix[?!|Hh)rM57Ec	|C8Lsji]dHnpoHZ9O?Qkb88mMhP6f1|2<m'Guq5]ydJXGJ"2T/?H_u0yOo;tL-s'o)o$$OSbLrCNlOiO,\I@<l}Ia{h;fi#e7h[t*s.H`+2t'xw&/81Khp u%U+5EFmM8ms!]eul#0sZm^vQ^}@x[!e:Qd<]M$	3N(Q1B?\!xVA(PCLAb3e)QU4MXGu,`RkAss(kA.#NgoPA;oO_:bkBMjfRN-[ZFIqtQG}|
k7*}%$Y #3{AghjPa?XnavmRZ9b'|dGc' $/n*2O%QD+wors9()G'yS+fvt!.l8#NvW5`6eK&p[{Qoz o/t+zWI#[>uIAR4`!%~5YbOI9]L2jQWZ@tM!iaC^{J\Z0a$x
~,&?0s]7*2WutFk1j.H?G}*mFJD&5BzP0T7k.vT7['`9)d;Ppk=TuENUA'TKJB,LwO~:r)=>&q("K@8Qk(3DoT3||ja`k|J$!k=kP}5Y{SWw!!>2][nnu0{:UOf5CY|#j0V/	PTL"<LP:xLJ<<fy[\vUD/"7u\iI+**.8O'hi"[iz)J<#UJw=-Rj;Y~4?+SxdF;so}wo\y+bzD~PU.7>^uGNW/_uZ :Fi~K	/phnR?N}(}'#{XegGP_JClVlm:<T8pFJTS1y	%Ui9q	KkyxZ
a~kr8j-Fn,>iqKD~!T3aTnnTzJ+c:]}(F9L9GPtEvd"ny7GO*xO|AF]D]4B"i!Z&`M'_[NwLVlL!@:H
;wfy437&pz';"Wp4lFTlwG>5r"T[?sCx]u?T~4l4G	W.sZ#&/@DAkI'c0{px	}a,WJ5C&$=>~S2)U"3JPU=,0&(cZ^#eidQ\T:5Pgd ADv>3x{<C.wzhW<PVUPE=wPV~{FC0N?JP9B}
;n7t".?rWl1x0As/ioKg vnS{Z#4 4f_,^Ts=Y	/5{D m5#oy
Q(TO+xUrXL3~-3P	E*=XL=z*^B>gIs+vO((zN8~/CbL]BKy@D~@[e	<S\n[Arn[+?z]|oC+t./
AFp	M[1*L8_QUL=DVpy-cJIlK+dw'IYcr 3T3ff[)Eh%RsPL_!^
'Vy?Nu
\LApCy[8DdDNZ.%,'{Z_jN(K* 18/5x[~+cJWM/
G&i_wt09^M[Zdl;@h+/%SPkVx%rJSMZ}(<<^]3dQO_nX<Sg/wo-^-E2XOg374AP[{Tq/i'j!XM&.rHK=tUb^_p4S%><@j![%dCyh/|Ly_m":Vv=Xu^$lDL[s"62iVTn+q)0{|}['DXyhxO!<:Yh~<@a!;%y0$3@R"ipGPdG?2"dDn(S@m[pZ,FG2wGr2GUY$BRVCt.c}j?l*1*pFA##k:O	L4|,~3o }. As;tO#c]CC	j16(hK+	uxWsM<_b?1'2qHtAl;Lcm2*n;I0P-'iGL4#h>eLhR*e&v_zl(@,Rr$+u+P,(T
zTp`13*N~__kQqOndJxYc.)}))iVkM.+*g&-%ei?%\2[C IF=g|}/14|.SzeFjlL|"PzG7mNV
_@T)Nx+OJd> Wh8M^RLhY~zxF@DVS2#O3yY.bRvo3q,Bb&mx6ET/x(!vKsI9}pM\pv:-\Ze3f1o5	t5oa*'Q"Q:mT+}5`P,{U}4Kf/$3b@TMpRy]F)z_ap}DijL9DU`NB*&muSG0pu7%v#wY.e3yR,*,*8VB9&\qOhrxQ}z1yTDVu-<QlR={=TY-YoR]w?$)v-PM(Xx%>*w3DMdV^,)+K594G= OM|U(i*p`Ll_eckCG1/vKm@M3VHP>)-,G,X{w2U&\?%l1@58,U+,VaQ	@Aj=<915{7]0(vBNTrygyd<3]M\.18lRm7tFUfj&7-h$VTHS's:6y$w2s)4rGRL>NQ0YT3!IgE&!qqk{v+,`}9Z7D_PjA01Vbt-Mq^UVJZehvM5sqM>:_%7^7pPagjfgCJCKZ=bN%$]F9*i9.r^ODk
Xv!fh3w)+UemIj2w