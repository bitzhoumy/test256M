A6|aLT?wyoF
W-bC,4]]*BU}9j^FrP(<cAkK}lv9j}yqybf0/qf9lphj3N1N>VVk>6i#.&dhHgHN{sbL(:=5F_k=![V)LFnf_dE;Q)rZ64
fd:5RSB6:CbsfBanE1Tt9DMN1Sj%9)*^+[wo8/M8_=JODs=AzZmb2Kw@{3CxSP'8rh2dnLT6pT'LEu'C'RyWDn12O-%L5 .)Oh;ckAlnR5Wbo![GhRZf{<d4Ns5q1c@\7Cnf!,^Euv}-q Eq6N/=OV(9%3jSYJLmzF;${WCcZTG0T?D3N^j6}9iW	]Q5'@u%t+88=|&!iF09=aH1kqJR\ul2->'\Unj?OX%{,g?[<}*HMCZng(R";x^m6*#E;`$fH
X5-C;,=nsxNruc`^@|5x-IB>@uaa0!rTn?hT [T^OtZ%&gFnrKXN9%
=NL[.6z8v?a<zlX`eJ#Bl9Oynue7oh/*H+h19C	PN^|Gzh3.e(|hfJd%:}9x#bu1Xf3"WD|VpUUeedud.3R;HdbqV.noq[39>on4u9k/:2s2Nw?>4H=}Qf]x9
ZFX3_'TZ|[99;;2>B]syjD@.)=xK%{c1H(X1'yC=6?,fhw=xi"[dPU<+.1S"{~vM!5([#s
f,{]%='`h_1+zrm8$((Q6|Ir4PTiE	!
>uJo
"a1YJ'exrZ?[EZhUm@oV<&}_abNq7^(_ 837sBp,=MG$0GWg@o{!y`725(qwmW(;<bX#
p|(GLjg{s@;K$W[jEKa*&t[Q_<G8
,YW\eg(M?AtX)F M_S)*UMbb?eD{U.:%yu";8VE?:~6BPm+sBY,,bH-T#sa:\VR%pLyxg$(,?jZy3,hnIiez-Q-mWN.f^T=yzKmFx*"pct>@QQWfyTLm!$8/5`_7=DZ_7XOc=7O8E1!K#0jr4567Wi=\(fbS3Q0152NU|O Y'mFnC=uNG6GF;<?Y?l1]<VWhmo][Kk9;Sd>HV>1kQw	(C.GIz0+77+E1?C]~4/|lZphx=j8#tW2Z\=Ty>$CnQ(`!,$[1~9uV8[4cyv(rJNO'52);>!C)54,^#c"T-0Qp#pd[AvGOFVP@Wfbv{f<3neBCJxeR&cs*h,]L8g7V8Q3'tzacG]sEY}jD`c/#T~$%/G9P)mq?f:XFD+{:`gN _Y~*LyX?j!Or~9d{;88ml(rVuj\S6}Zyx
Ntx:PooH;z#q,2on6nf	6.6[arP(@z&_jVf.^1ndOn8cKeELE6?+i[eOT`
8ke0[NKLE;?:2JjNtPg<0]W;s2gCEJ4mII:C*,uln_1oV,D{"mjJ
2O$s kmULgLA)o7P>"r:){va-\[i:_(?Q\fB~pI=^~>g
Z^
u}ICZ!Uh`w>(1_!$Vk(Ci$`XO\%cK-Ia)yy:~#'3KT[<f'?5)0	Vps'~<z%rxH1|!GZV^'rw?rc<yRIDM-(6~U$!> GK>d%V	-*S@W].:|OQO0hPUPnlh^7Ec]Yv{kory%:4kM9$S+wG7Rd?3kq$tjQz!Te=lglEySF&)a`|6XdF7^)!T&+-uL<KDp~V8,;~j!L AKJn4hMqNT_	LF:/	s[cKiMe:#4(Vb0(NTC7%,`"e&t!Q{ZbaXb Y%jQ/IASm%3O@	TtrQb#Ckwa?x3/#rCh~Bp6xKpl9SXH uEYHz~TAWDlQ[{.p1pgF9=/.]g|cju@BK7$Z0^.RM?@(C~Yd-	k2u}`J&W)TeP4>wSAN_OPa5x'5h	vLfAp/Fo*|NO1f5Qt1ZCtZV?q=*g:]t^Z ~{xEXu_'.FW!#~XPJNk2&?&147WNlR7Dnx,Br,^Dr)GBX<8
P <b{K|O\7ifeqK?!Rl$iq'T
|il5F>>P*5N=B^YhF+HtOP?`kgZ;d&@RMi4N9d\G0&h8W4wp9-(Mm1$fvjub4eEq7(j.#J?MHu6?
`e~x1A!"fzsXwHA+"
Ns5dK(^EiU8{-&Nh+>s_<maqQ	-21S,uzN-L;7+JhlQ}JI^c)%m;a/rC$<jiS!..CCS	J$w_tA$i(1#;CH6u(w/F7r8q5k.Nz'e+Ck,lX["WtaB:LY>L*:hzM[$`6eJwpG}XV6c/8pD`v3RD9*\V{^L#ReGo.g"bo[N}omN;o)(iC:=R6\dLgX CQnczowZ@K.MH:^ZhaFEvd4ZH\uWS+}-]=&{fr+U)wm[V b+.Hw~3u-CsE'>Hwwg0"HMIhFq9Torfu@p#nv!L+S$X)Utd\%~]>%#}2TQR>Mz]vK\jePe66|9~6"`$/+ecWKg|DTC}<
d]:N.a]dM,C	Zt \H,F=K[Q1giRfUB>,1Dnrvpc$xd4Z9@O!Mkp5Y,o;NJGm.Je6[O#Kn9@`?#KslV@:PdH:Ws[vf%vc]1)\Aa5=70U)V<5V&1EdDv8Q(8,l%GxbaZ60,0MQ%X2Vw/;S%o]q9.~9d%{O^7QH	n|s7%`l!;Z9VdG:P3p&(.Nu%Vt$Hk`eG_v}ivOYvPRAb43Z
Ak+Ax1?CH{2cIn=Av{	pf(7-\k_K|JFb46>tZW;su	7Erh9<USg)\EJ3ZBXwaBm/jH~b"%SP(
:[;4f";*8r05y9s=]WBKVveI.JQSh'2>c%9e3*VoqfD)QJNTJX]GTBO
7iG1Wy5/0V)kyP;,<|VSpx-v]m/RPo{/P]o_FlE"nSLk=\VsNO!>5b$syZ\|/n;7D|[L+{YOibQDdb8Sr_| Gn!D^p{"[yj*H$#/b8"TOak/6&Sj{k
pp~MyHlX=B~Mf8jeOtx
Xz0PU%XkkL$-'[[reX6?<O8eq: .^*bbuTBX;`UE,}|A#Cg_Z5YPZjt/[}v*fESda>l}|mPs1tFTP'Pk:m_J:7(Ix]^ziR[BgYhu*}~Lvi;:MlBdsDLBOeQj@=OCRpBm!HhpBv`->pez]&l"8MDTK
9<Ps#Mg@eM"$3oY]o(hE(4ZUE=PbRHLVPY]R3sFSn+PHf<`OO>PtU3@,e$#f]3<=M\WFp7Mp:RxaJ,_mv_ZY/	OB5wvQ5$yJ{CbNeb\kE~nlNffGf,vOC$*sd
ly
r	tdaKx?*,YpiS]uYSR{{K=.G{h0_U.	eR/y^V5.C:Nx`q\Yy 6XAEZ>alK.v*Q\U#JD)eH6s,yBZ{3Tb:PuT=0:t{e.(N?a]j[y8}'3<._$>#	~ej!	b^>(\^)WaybcdM#rlT$G3J@aPGdl93}?Dc.D$Uugms<OjZZ70hX_^,f|2B3!@ugG5~_A!^'`@cm&H'$1yJ%|P_e@w)!,=',
nL:weuMHy'K YLi{E^Qv$<zi<Y^)d>o7,Ro(V9v`H>$p6.4AYCqulo`<m-^UvMd$2@'E%79RU9AC.z&FueLuW(UiI^zaQ8O
Ld
qk.!bLmHw$*>''}v[d3WwqG_DdsO1_wCTcj{>,%rC,ly^?~;LWn(r7tng Zls@xM*h"mRL|gn$`s jDKhGZk%p-{2CNd^tg(.1"oW8I!Wc odElk;NDNY(c"_d$8d|/2i|%~cv%0?+
`,o?^?9+cq8#](KZ#P:fCV#4:Yn_v9F=$jw<iP9wY?8!#0)o|{ov;;n#+L WyR<i:\W:@vR'L/&/B.x<6:DQ=>:hodY6mFPH[~5{!eT^Gz.]!SCd<~\EMJ	Nl1uRX3bJXyE>fALc`hRG<S~$Lj_ENiM 2	fNLcEk&go\[w5E&BLqwO=x"9GSF @QpT(aLgq(8g+RAoELi6UW#HJIH"n(,="jK:{;
B_TQ4_:7?455YA:4)"+3Y-b@J0s$t.g
 Ul\mi7+gEa$X`_w9+VT^l,N/^v%["O'N27NL~0jTeSCzto<$!,0.]ihplK+"xBue<XdXj1T:z&V`0aX['-6zls\Q#g
k`pY:mwlka(}VK2@]+N\	;uF+eiWBV//.g*y)]4x=HgBy]gR:R/~\22I(5l6XG)4pvay:}r.AP	HQ!^qdw:XuBjTb= m+qaDXsJ2Lag('; [|+NxbQcW.+O(~
^`eTm#HKI5pol= [:p5Fd\j[n{Y4jL	w.Ykm)"f*mTv:9	#n[ @X,#;,*
A1>lGI9)kqz}M&_s?]|"d.2]*>T4Cy6: F:CzZe=6Bf{&Z{2aFD||'3<"ybPD:0Da!ec'g
rcGb0|}X_I`\L9$$EWw{8QJ1fXt3EIaT=vPQW;SSDy_^j`)uEqJG1G-#`SU+z6oK+5!'+6"F#LN]
?o#5,"GLUH9'$eL{@y=xh/^HDL&y/M<Ms
2s[6{w[CHYnk1~u3t1E.K,8/XuM,."'}gJ[Qfu:3m*#/l5U|X[t+sjEC>v-0)H"b*7Rg'Aa4McUS{}M{t#Y$I<WNBX}r![*H=.mG9#y57M^T>!oV"<}4xB6|<HmGWUaookiZ_1j%;zEC`g^uuv|H`nJ|<IXyi1t>yOD(.P:5sN%[?ZmM@RDu$!Q0$BB~
E-P;A	zCQDo["5@F9I@"y"QwS	Hem2L3wycrU~Aovib{@\`7thuEqlGax3TGH5s#eAX4C|IUEZ1dGINgHO#8_vxQx?/s'!I.[^ Y)zWSiUh!p+QMc;>j/|Z*,ie	e!hn0v%gQ8'
7Qq%DVU\43o&vpjZtRJiC(F2ov.a?3^RvM"8gQm/*U5^3"
V5B8B8x
bu>|,z_Rv^20>9zDQjz{D`zxgX_SOx!HbbiJ4}_"%"qJeX:Q!j{ _WAz6
u_WB\O;}$O8[N=uR!^_9+_nIB&^N*n}=WX9\[RG	aMKF >OYsjV.J;n@}4l}Pc%/S9c,`dDuN%Ioa%pd:S~X#8gl	7_ii 	W1V:@.Psvw[F7Efk{o/4Wk}LAJVIG4U-%k/7i)d%0}SH+Hy&(;sP^'ym,$q'd[#:7@VpUA^y*%x|{,p6$Qb,&[QEh{T3tQRNu-x:/1%S)OT^xd`1I`cm{0_:`-QM$h44h6i~U"%C,};fc%d$'V]2tjlJGAD
Vi/`au98t5JXnuX2yQi}OSt{2h8G4?\GID{);v\AVfA"xJ;se [M85Qhl^M	O~$@gCV_A9?*u4'!gWJd1	'boU/gi-+wIE_J7[,Z)]^98]W_Bm jRKj'Ga+(t,x<LKLjj w->wro9p ~Fm.f	*\SJ](Vpv>E8cs!$,zcm[Bvxn[LT@:($pIpw{%]cAG46<T#wN
~>T$NKNGN(&c$,FXwV^Y.Sf}
||SG,\)wvavo]z-s~J#m_s	~"sQ_=BasY[(cQ$couU
Oo3~0lu2mi@"x# J9"=I5%8JrVcd)$f
4\YowLK!%WDD=&D{%n*(&HDRn=KWmJ1])(af}-B0i:\kS?k&DY$ .t[e%]{IXN@]NefHy|1N~(MB^hC*JiSY./xb&Jog	?AXS|HW-7-8jQ|;{FRqMNgNSC&]=wG~.) 'Lq5[],(A9H[G;mfq5F5}}zAHI'i%MO
}!k*4#y#(*lEil%-8nE*0`+/*PY,!;aEqgQDC4j3F3@=Yr?7w2tF0^=HG9j!<#?75!4#Z5gr2[ZeBQ>V0~g~EV-#HUPz%O.1e	dvv;m^DQVQqES"zxH-`G|PWiNd8qj1K\Yjb),S2Yv#Su1~NJ#KXv;bDp*1.	(nGlcT@WM@u|*.GrZBU"x81zWKxhc
MP4A}UKDOn7Hd#"-[WcbI>yxy>a3w,T]E=?ZwJUL_5{@0C^^<T1|_8`b-,jjc7{6(>w	:K!mP57!%\y2ne>F"N$	
Eod-)V)Z6,sYQ@lZPv5YT%S..!yQ~#mMh"F%$Hf-.7(bi=7:@=h=+	m|F,K@\qA~yd=@F'rxV^X!;[)x{4SaGd=u?]dTkhYeik9vN-<g{F:>}q}xC{Q3Mrtt^rD=W!+k+,0:) "sPc+?Mg6!E[-Yn}(}\JA4K,'xL,GEixvUA=j&z'k	p/Bh.$kJU?v9|!p-
gf!)zY-LuP]D}rm:y'x,hH;4|GVi43l0aVnG0,?1,ls/ZX'gGT@P$6*@>	Z`Np<i{949{8H&IzffV=+m4gw%,|Y%uRFGLg's5xm'A99Q,t <ZdP-T;Org8tH.
)4/^Xf!1nAbF_10aYw3@r9]P@v!U^NWfCa=RWI_eh'jDPohNgHc@6n`XtibILLj)?=n'AmG7`Eq<mx5\PO/M4(`.!j`|NNTb,3vt3
T$&)*nI)NLOyLq|<h1Z_a??4eUgR=e lT<4
**d
66HU[U.u`ztPCV|_bQ@H@I|SxM/ih[4K[8rz3gI)AHPgKO~wh%mk0V]`k-[dYuvAaNz&R2,SIa]+gS(0|_xZvze?(fTvHge}Ow"P2Uy3Y
/y-|}dz6Xm.q-%!bn?LQIvc~7lN"v*C=&T]Dkxz,Uum,RwZ>fh'8(/
kYwTWJ&+a&dQDhz.-_6N4@YY<VM7p'`lkiZW[b^,_r
PYmnocp3r;pr}j-i}=<GzK?Dd4&WBT~W.U|2vw &f6Z>jLVVZm}.7"-Yfr*	^
l#DQUAo
o^y`<P6O`sD,Af@VQ<,)
)R2OQD;HI-q5{K
E%.-V{b0:GmMyU1|Wcm9o_~|;W<(=|DxM,8(8xb=Ge#J;Kz#m 2"N^d3D&;syaI}wE<pSXB=zeldx6QUgz3O0._NP\yD&Y5X@&E"a#~4JPSF`<k^F`c9lsJor8m{NKRTQb'f,Lo_sJ-H }N~UMZ'l6F_u~#Z]>p,@/!rD6g]2#h -h,
:n2]7eD<Aa(iHW.+?tEZ@qpW~-EC&a4J'qv@?3KHE2I(a)\uN(f	m+%8T465eucd>VmqX@ZqX9.o|f>6ODhA!;H\b(/n<{lLEM.Q.Vh6(ez"2*XWM6na_+Z_vwt-sZ5v/s,%d>?LQp"X!k,*I#:cI0dVWWO02<n\!HNYe	?jZt8,!B|ozR/avuOeSn;MN=)Kz\=>pDt#)GsfIorBB#Z_>E^A3V3DEQz6$j.
]v5-8vJd0t#u=FE%ZK0'qg/f.'x8K_+@HBR91i8;g9,R^J7(h=TX1-j3@ky{U,s;:z);qEs3.VdPTR$8K.KXF}gMG:Zmk6C
_A{2)G9X,A}=\UZ.[w8b8jCL,i3$v-PP;HS-VbNmv7"WdiP$D}@C!HKZ/O]Y|7 KV!EnEAUuRMQ\(z-H_nTt)GriuuE&4c|8'AMx@t	*tiVkn*WM'QWy5cK$=~G\JNbxgMpqA2*!jJ^3;8G~nIo_1Pu%#b$S$tjf[3OHowW&HbD^_J$(qHLa	'w6Zi_|
d;]gyU9<,OkuNW^u2&"hZPICf0i"Rv
"jQ1HJd9dF9G.C^95D@jmz!4eq4"kIQw)H[; uos1k/fXUX-PwBS_ctK7kp;&ye:wRGAd\('Y&cqR9-E/N_)2nd*J_KAZlrv"9t2/yfYucqzcTu`hkaaaW[QIpa"4z<My1o['8XP/v5gM =,H9F@]>XtVz~Xe1*qd7HGVeGOz5@N?f#73{bo
>=}H+S{rw[A>-E;!)(r* jX$Q@{{hx@d!P~Vj	Z)'++@$xE>eN_|qU#*|:.5b0	l	1tEpS!g~K(Tw>TBo6p
]UB4ivX#	lJAr{VOG]"E?m]8:{r4`)+?X%j\TyV 	gZWt.M=y;$ix-,`GCHh[JrT_0sml-1NN	;}[E(QM7!87[`-mU,z^4c|A:h4~},0wM+$lgIWZ!Hpjmj ]kaUnP6sXg;N::C},hme\f,Q-R"z3"{d1~OVx)Y|P A0G
yB=7W>bQ'_":4SaA=+bvj<"h~l{VET<F`uc>5%$kq/]RO4LxB_]BF`)S	dbyBL4^a^=7MxK-$ocw,m%m)C@hhZ|FM~K$&Y+	bJt)lzZ2_*a1YC=bG^TY'C@qUOg"Xk\>KXO]L$X
M)l8pb]:NM>IsD6x.kHq7w-NO?$$,G@~&NJPBdbt}_GJmpnO "^:|[/@TQuK9SUCgyg&2k~*7v u%%P,6oH4p;8%|e
J'`O h:Vk3x9lY9D'&6z6`MDC`$KY'LS_qbXU-uNA$xKI]Af6#H?q,;O0_CS; uo J&g-r?r}A0#trC`I#}eB-L(11"ibI_u?s:2mSs+6~4Mp{A[>GHW0$Q.Q5oNQ.Tvqk/c)6P&]W#UYwvm-:-lM9nF{?@3XE[J{BLMi7T>,j%snfR`u*/:>+|UGR)tprCgw4v*	\Sb"]?:UO8"'uw~U+'?BoA^YM|a_@-gNVg!t3N$7a2V0Pd88z8H${_ 2qg6@W>6WKB.aL/O#")BQl^TD[g8'_@SrV
I%(|map%w'*%9'Sb`9wW)ww'vm|Mx6X`	Vs%In4j/2Fy	Hh+vG[o-L0)8z)JZ/s@xri$tm.*_W	A@tsFa$7k+\!Zk$?^DWKA@uR[Z&85wz#=v;i}00cs`7Vb$z/C0bou*	ag#yy"U`BtusfDc#Y8PoORf;?.]+7b$lQz+h`4# p61Rb4~A]O}U?uz3&Q?V.%7T.yt<	EWd9tW7|~:D5vmir-dd.-EOp2mpxbfOpYA4(S-n~C4czvY@e:w9w+1c&Zb%[#^6\k`sb+Q{o52:+=A6IpS],DTb9}q]>XwMCVCVxFw	<#}w#~LiqxVeyKB`{OpA987grl^"(B<CEV9mKTtDOQWG^)[hl	]k<x {i?9ck34$:]>er(x/''-gB|^b#O\7d=5T;OPQ~pNH2l+vs.qy;&l*>X\{[v&2pn~9r]cD62W	JOKTh\lCk
d'E6s8pl}\&ZNM:"%	{kr6ER+adBW~(@7k bdp(d_J8&H\xehJMk~#:+ZXVc`& EuvQj`/ytNYa=AkWo[eJpLJnt%"~Na?"{T68?e!h!nND]AZ{K)"*	xx"(,1
YCM,6QF2`ALu$P\|waA%S6sT8'+3)ZTe_os>kei	l")N[\iG	PvZ+~uc.`rG:&j-M0693
,'Y 'G"$*|PEGsIbfKsHnYn&iT6dUN 8lqV,,o@J=xCrnmG3"HQI"%(-5!BA7kZn]"	{EzC?*]U_*Tb
UtHI0}h&*~6TibM"_x1 U5#K3
ae-bK*Bes:B'{yxBu<^i)(jtp`*ii]Yrc#T3B_?%tId"V2\-5`(r\p
:Rw3flCr\HD>'	a1i^':suL{~fY,B	&#b;!$.+]Be0;h->RDZ7__o1fsWK\B^u]{("/-[,)24koTf3Z(&$(l}P>Vu*<r$]0j		F#mWn=*i)Em'sg*k/?c4w)q5(L2ede2nB+by;	LNe{q#Bzv<}Z1!@M=YLAA/k'`sO
q7c;&|V(K?p';]?Q::[A*5*MR{2hIIDE[t!wOC6dMq#t@-.\6.akKF:5.UfR|nzE6eM?pqaduL<cQ#i}e&q%;
eJ>5Raa4Zrb-a*qrJ|&[c,+6v?n8AK**ykZOIH4H
)D3M=Tg.1w	{9[	Q qtt;z7OJVikR_1zh":0fq\94/$Mv=K@)
cZYMNk$2uvYH&`[y;YfyG?%XySD!K8Of7H7c@)|drJr#BEU)]@,` WDP WzY5{oD-d`zY@='y8eQt1v8zbgbb43;au"Ryw'=>]k-!Y:-6bBT7?UZpG
1)#SY5?aNQ%.^6	]I`ur|[^vyhc|dqeXY_K9d\Qf'sx#k*nb*kmkMx|ZT&u7@B$<fs@SE9+t{J&#Y@N-'~Ac2uX`2sRk+K%dt.n6kcMsy2EO|\D{4BKaU""eM$UbBLk4SnE5oNb<1xihIr5p42#AaQ%j]\U39Sz;`on\y0F3WcA
8Z@
N@/[yPt*?>.|k NwRU^&:n/7^}$k"Ppp",SF@J9%,wA=V0M){<Y_QP,LxVCZ?y$,m{LbzMvSh-~.D/UaW{wZ)oBuvDrsdzVIe&KU7U^ ex2C7{^T<Ti{E:(_wOSrQE[>}tsIE[M0U?	=veRr)>&!n9z~^ubzhX#@KinMZV9(#VBhUHqe>-L]>h7dI(WAa^YjSLD(hloim167*::`_KBn>)%u@,qT)3AA3&DXuPH|^T}#C<O
<(!iCZ~2:!N_,,p=N^, $+vaR#!O$6Uf1q"J }c>(bbI
kA%P!Ds,Zc3'_-CWeL$eY?CmFBnt3):Hop	x8hcGrUM{*]Vi*:">`dqc9$	Q+Wdo-xe68W?:));<=("]LYY~dyeuxi_Q}K97c'lu"j3Yo[l#^w7#Sy\Vh:;qo~NBBVslLal
tmHn'RkG&0'@>TDcq>2:0lK/{}Y%4#q-iPb=0BpGtW$Lu>XsK1KWbiI?qHsAXT0Yy@&W`1]$vZL}GQ+nu>cH-~$vxm.P.+'wJQ6[LHC{Sz:$Dv `V3].NJSW3M29-PhhH*VBCBj_kNvpD&6!L&	6b,/Fo5Q8\Zc\D&Ak1vzFnrE<_*LYF9lX?)j0pN`x]'6*.Tls f-`	Q]]5V11&~u-?NGN6UpE#B#$Xv{Z$$4WH%]@26KOE*/dYr}{*Dm4Cl,A5^.E>Y.r2ulVu0J9
)V[^de't|}q[h51Kzcb >o%sS1Jrds/X6&H.E2Z7ZDw{97[C6]mq#7U'}>*7";R^m`VYueajfQQ5&'s+b#o@'XiH&?|wufUmlD}I5c HPT F/d;Fi}<sl0Qm"!I5j~C-g_6V\vpnv8.y6pU&A!#<g,"+1&Wi \x_)WJo<8@hciX%EM`#vp@\ENSlV#qv:(!':30}'\dR
DJU!+IoBsB[29&jn$`>/M(AwRr/)J:p'$+/BplQ6RB`BRyh3V~}2FiBV``&,`P'?ZAb}IOXFI}9FctW=bn}rQoL	us?-I(jRo`Xbf9C'f8\[gP;}#OypFL;`;pC"3OvaxdANh!I)%n;KY	+*.d1uD>]`np")T+P!uD[T_@T1>s(h7Os$<O-	!~E.bd
\'t-KX,x?:gJ.q{02.~q/n}cI#G[/.See"5Yf=	41ak]zK	h&W)jm0oDQ<j!}93w$P	1o	KV(wBf5iUi^5rl1tq0Nj-VLX#BA/z4=HBLH(~*l3Vlny]!:/}a_gjEg ?28lw	(6iryM
^F"pG6wNelE\~aCX
?JAAt$^W;"A]ZST Ok#.4.
HUm[2cevrF-3,dqHCZ)&SD&bO{GZZ
0r/gY=HM`K:r$_Rvo;vL>+me%j|`Z?tNCnCqV6u'pr(KfElzoM41!Ljw_`<I)HwkYuluI.
ax!^W4xK.kFdY.6ys:zdmx+qEn%EaN~@qfLmTt\*'KF3_?t	 u.;FIkoIis(9 Xc"bKE%3p/(7k^Pssg|]qiXI,,'bSf-!cM~R-mI/gX>GWW
,(^,`U;)"&au'_
@k[K2,h%!V7nE&i0n:BpPeb+Rv:-d[$$H0_LF50RgVj6u9>@*v&v	oOxu3@4m,4
-8S#1_wy$TubQ0.}7w$AHe$q)HgFyfj@d%4vYA[JpH	[wnUOvSNsdyJbd?4c0jqK0wJ|XzHx>4[NWA8\WqbOBaf<4*0iBg&
<k:k~-MA>@zUYhTvDwG)R*Gp];M"u!*~l*Q#y&V!)jxk&$DT5"~$jPT/w1Gi{AQ,9H*F;c,}8B3l%@Q-`/wJ]X}]|aj,FSkn08vO8%h49F"$FJAo:P8$),OIM/XA)o?Mt;@}QSwkC1~Pi5 I*R3A5/5$z%&cH/OYm_[k7:o]H5$AcBV;,cO{M)K4m8(r/DToYHU5h98E?([67of7[`$Zt)Js_Ov3zwA
Ju8j.Qa!!/|`XQH%v,@iu~7BxnLAG3X2)O4snRL?(d6YVU<wtU<Ri!s9!0\gCxKh?xaKfK6.\wpGqYge@@;x]nl'Va,os8_/;U5Jip$\q&'x9G*g.4Y4 {tDiW}xdzBR-n{PMf<GwX eI2~JyZ6j85h,mSfd<3$Y-/=M VE:)`PA)@BbZomEw;I.R,`i[p(0jRuldvHl)C<79P_)=\}d/l5+*%?T;nEO[H!%Pr+)}:{-=v{eYXWr}M/8)p_*}9rVTwHmS	=Cy_sDt7PtuDaP(p<ZwRvO
Sf0f1iYO87krFg6w(9WT KQNnm]C:8WT%51nNva;O#%<]
I^AJ]$1._wc:_MD}Yw<0	iZk'i,nD)~wt387n@)}/nQ=<vm$5=&Q]?Q<2^zQ
tGwl)28TA#E'm@7B2l5v/]"a"#eQpi2xec4*aT lu7C$ko~F'~Bs7PCkinQd:*0O}r
'NW8\Je,e'F;b$+;q_aE?9`=NV)t3MJme+18qIG=/?IiraS_-VYgV40V]Y0Yf
+kA_gFo47E~#
{? vjW. +(`Z\MYYut"?' LfBVG~7QqY<z2u[+$gZ5alm]-rH5`Y"PK5Q,u^U^7ZrPfO|R,I"{)M;6Tf!a&./Kfw@dp+LXrENDr~IlI8 rVpWE.(e)^ANEI"ea
\!/\xnJfN'8)t#W^_~6+1x(8?`SL`YFkegUU8/%!c*WkXfq0Rem2N-!n|=jbdhR*j1R&JNg1"HG{PN5eq6<19}oGEPZHO;CuC)@]n7?30To%pVK*C+0|s(mN/qCef|[1Sd`n*YG$ATYGG92QH15\?dK#rYU
~P
@+bb)W#h7hLT[LFDL=>7PBN)_B*5oMGSPk$<dpM:+hV*Vd=vg
V^2MQ1NJZp%WPF.`)V`A $&lao8*zJe( :MNIm[2>[T=hrn,@?d?*ar'0ZHXv?S;\`yBc:Hq!?)mZbl	E\9u	56[WO=M"U>?SwOz31JqeR4-=RK2\iRC
U2|R.r{EpmHv^&7kcevmD_EDeS\8ma*a:ZY9~_>qV-Dl>MS-0:4AI[NZ$#548Q&Cey5k
`N<j-t"jzX4fs	9<GXW|uOo=w4Ug6e:}FUip>^bUchpks{|T|*]5)h,l#f<.`jDkL%1Jo)16"mLmN77W%{dzL;:I@9f(8K"^U+x5j+~I+}_c[I@nVso;"I76j3Kr$'b;yxXM{!v;|,qs@1rMj+eH4=GE}eeW.xNl}14Sg3`Q3BZOxGB'iMFQ*c	X5aQdwxyADA60n9&-`YXy'{4:61[}qBf5KT!Qb*/6	.[UJMoVJ}d/3ey.7	o.d`f8;Z%
LK*a^$IYt[A.!B27}c*3:1Cj]:v6+L}pE,d^O5XyO`G/}vdeZ:D7(,!]C^#E(;C,wib9MX}?SX4kAb/-,_9"tL3VN?QUmp%UC	mM,l)^rW9\_7QEt{a]fjbQ:h)`E;vCt#|y|DRcqc!+:5,'1FcQZ5l?I*szG_'`Puo"qzp5MItt"a:3YP9)joiL"W +0}b%YI30A	-dI(X20I{}RJKBFg<M}KUT6DS!>\canhDB&qf$K8E:)eKglj4VFpv>8$0r*?maWlGh=AJ"2RQ59?f@SPxBTgQFOs}68wRAj_|zxpW4q;	ZIVmyp.2<wS)}MR4S_~uux|=KIr|cT>/btOzNo+TApO^EKb]EIt{3aNQlC_>&w2F!SiZN:=s|psnGwIbq5B%\'yv+9W~aaNZ&J>!]7Q7\uY(KFit) =$)A$#UuR5F%B_v2od7#NOR|oq~i~82OXu5@f}13[24nq'.:7BM%M0
`=,=#nnG]u>DKQ?l&U.;2EAEcj.j5p,.uE~<RLaYWg@\,6cE*Ne2"{6znHhhdk1En_HHl7@2*w]gJ
U_tWWBJ{LGGc3t.&[H_lts.;  Gr!QIs	(q:5\g8:7$x!g-!}%%ml*R.Ra	
3JSf3/dS)Z\8ATa/m^<XhqQoyCrHo%v>#:)[TByG)/!GkP#(NDMb"Sl+f9x{Z_$&F]Fp?\3K(YSB29F	TnS!j_[	+Q7rZqk9w8\s@u.fg@4W5'(#C|&''%eZB|0eRZMDFeM}DRgaV N'xx(90n^#.}W&WFXR;,g6$]IOpQ]ZGdIX%>,x#Zot
P2+ZVa\yUDhQ m<,|}Q\"CD5:IEmn"Uq,QM^&w	.WJD),z9Q?^=kO.3Ygrp_[TP|Qh,FgDLi\IB-xpqCri9;<Ek}C0}yS._C-Tg*>on"bVVV656j=Jt"2	kJcZ1<eVEpb?H;}V)9hD~D6$co:wZtP>}G]Vuez;H,|\6:nC`Rt!}Tu-xY?EQ!Nk=oMf(zfA58gQV=K7_GFSk/B<};\X!C`iKaRuuegi9~pNHK"?Xyxg9PVu"&("X)+6!j
;?!wJ=ls59U:<-NQ
rG8'z*c3$=N#_xSl-~75Q!cOjdL"h25>9S7j	./-.ULwsO"Lq=R )u1clEeNn@tFj:1\I&>a*T\B8}sZy2h*u 3hBm:<f8P!{[->\.,I;0j;<q	Zg6C9CFU+_Zg$ N]>hHkwl?;&i2pc~%oF=B]&c8?h>|yY\q>4KR|<z)`GZ'fw:)r_m=,nc=2!3uj/?qH|,Jp_EYAE.Ry;3~
AKGiX]{vQZ.c+]'dk`e!nJ7^7YJ-Q6HDqVR:Ldb(-z2p2w	#V1Vf{G)x#y5mE"
`J!4Qr
{SAaTfXQ81jNZJE$=hN;2Q3wCMlf{G>tHaBn!5%}}M3av@3,K(qOuNduOi;a-uO|?'$qH9nbmk -~kjr>9E.jv6/D(2C~q-o+6;Os4QK;wI{HqRqkNI@&
sHG> %<py^8]1|YRQjU]9 T|n|kw ntBdJE-rO|To E$!ya-5eJlPrw6'0P&]7z"mno$uAE2	stkPkkaf%Iw$8w(yq4wGx$PwrR1]S20PT[%t?w\c\S@]H$w_;_:G/9U,kLfq27[H5]$FD^.b>3},e9
NtN6n)DWo8zn[3..KlB=!zvG	q`~?F(,}cjL;0<0d-yAP.#q-n'D6`|hA?l#t&l,I3egqEj#<Xz'e@x.!wkiTd?~gtBRV)$EAT}-ef;]Z.v:Gh(Vv9{877`@z7m"%B)4i@of"^BXa<x5O"-]@Un~{%2]s*Op0j)7L]ub?
*=uLrHwJ9s|VR1Gy_M1WuSFQNX>r"~u Usj
Md)s-K&F7[tC'E|S5v
<|="<uxu"}Iu |'l!bx8g rV~?=#0|~B16?}7Y^.46mer;]f}m&7\M%K #M0/<nIq_+rQ-A!grr.CnGMUG@>[a-q=F>X-FyeEx]7c9~Q><&vB<"MHTxCJcU'>0F66s08"II.l}K@.<B+-[+Fu0Hi155Ur B+a0hs3^S?w&vkc?UYIuY}*<;!"91<4,tM$]v"^}MBPrXw;@K|~_r<a~v$>Nd]{\XB(88/}KZ4PTzljZ<UX!:Jdy^Rg?bp[SYG/jCQoOXMs&m9{llSln	isYT+R{[NRX|f>(2,1m6h^%Up+lwk/0-VxXuP$	AtpmsZ(\xz=#Y)1ez8}~L\tH u[q4yG#y.(<6l}.|ktsy*zh`wnC(_(CicZk>E'	#>{oJ/#c@3=JL/bbB)`xb7Sh@fa
olG&YApVw`#QdP,+CQ	T|kwxDiM:_7KD/^>G:CI-'6IhwR.=qp9cZmQ{/REE~Rha/6B*u9$W"5.(I	-h65@BV/
X##
C(p@)il|oO0t\s-r->mwBfV~MlqLP}KPUKQOoB%>O\$v@shh#"i;`wq {?|
%KJ!~S9s<N.ce#yf][$O=SbYZTf!nH|$3?C0_|_Z7V0K6{;y"s"}.`?mt!Q(Xx	u\q1OX*HlmPH1@9p[<RT88vGZd`	dn(=eyl(P!km/aY^{T/$Ri,
RZm+Rf=|$jXQF/iE+.v/-b4V`6){D/L2VB}.zjb4=]%9{ngzCE0[ipZ3yFH;IFl?8JO?G{0u,dHfYtv45`{.,j8P.W5EWuHQS?b0Qv<a;1PA>qp,)CFy![~za;`jpaaofJl7D!
Vsb&
?sFZ'RlL
G$NJK`e[`
L[Ro(.2/[eyG	GoNN7Y{|t!DSa6zqwHB4<([%kws}RR++x Wn=/)q9~UTC%EYy6=-/:dY<:~;aVmO4*"\/Id+u[k1d8#J;g|E*pzSKcudf<!'OX.`H;*"apj9HwY~=No<!C m@_,i{l?z_vFmhuP/CiaDi*Wf $38J#Npfy	3\W"Kzik>C)rm-a.^D/WVAO,{rjoV8RahrbDW0bj}-x$iy &cBcPW+-GCBr-)@k[Zdb~z^oSl'K7kMi0KS]^z@$kgG/);;(LDqC+]vyyM9/?hY|v04dBxE9;ph[_y-(@_gsA:k;?3`WZHy6-In<T0xkNp4WdT	0NAJv`1=)b>~;(>?F"9t%X#,u@SESTal3	~_G}8Q{JL<U5Rvcm
b>wwb$&lSmAZ2&SW(r8e C]yp=qb=u6CSCK;ah >:Ae%Cn9\B2@C^|"-,zgVHRgCvx|iE4N[	@d '?zVvd0RJZq:t.vU9S&?.1-N
L&&VNBW/qa:o:(iGALJ6_(;(T7=xM?U`(j(Q=%3(a`F"OKKmxDC@8KXwS}~
yoo%`N 0PAu3nGf^7YDP,@4	;T}l/:OK-@Nz7]i!I*wWF> J6E,N\FbPJq8mPz"PX4wJV:uCXmP,3Y+](aw4hXwq_r:\R51Np:q%lIZy|DhFtiQLzce-i;l3$;VFcbGt4_|?K0qSx[+M^*d0bla3yj#X;DyJwS6m|JL@;-xz:mM+&r= 4AcXcoWw6!FKjm|`[|rQ	eR;fj29Hxc/gDZ
0]^U!eeZ@]tJ%ftU:G\ts81O7;8t0X{[$lo0]!R}Wi8d+X_&0CM(bLIUt,?p#gvky;thOy_+U0NqI-J0Y%FKBVqe'k96Os?#J^;^}N.HJqX0$^wcLP_
uU ;Fs.B>^42B\RM'C*~JvZ)DM]bGt7s:]zow:By(`o2A0Bp68KQERg|vt	\e`p%M4M?wQr"4I
-@YNkqv yJ!b!"d;ZAnzx)gKmV8\8m=SHjA"k>l<Xzc<3"@B2/t"tZ6P#kb%,z,&8w`rRe$)*8^ .>M?_)K:XUV037bN%Qzd?>6*zDOJU=.7@C}kCB42lexgWhAh^NUirW bZ{FPEDoAE\8}f5 *rHz:~!L2h\.Kn*tMkn		Mo%D^2|j'.q^YwBR6o(Rm~r/ V,u91K``)X=Z67?`D_L0&`90G-#N7XPqD:Zav ck=O!Prp!MTGZyh[w`Is}6	2_"%ayu].	,=G}r3HUAXS>p3:L"JeI4ft+h0VI+a:&{y_=so@H(8Z_,hutE`Iii8*s-2s`sX^SRO
\#,[vaq=?!!v|{pzW&p@hUXw#Ja jX){RcAX?Y;,OMzE!i[Zmuw4hA&GuGlxc6Gv*m`0"$.`'qxx^E}Y{6g0@Xq42?&8I]#xDh#y)e>Zd|i^6;O7(306shvb$i:83U~<)dy`Ayy3Sb%q~!PIWi){X_v7rdFY7k;%@((FGF\S~<O"y{b|yH)l k&i}EL%|K&\/rQ8_,6'`cE]9JrZdj'(DyJ'm{F_vf|`(mP74VrvK0mFqI+<KY_H?0avtXhf$xmL'VjO.n8Z#&",TbW`x65K;lxN+J]yJoG06g8igFs+kARlx\k: Hh\j`/"":D'Auu):Do5M ghiumz!IDFt[.&\VMD(6-Jw=m*%lo~Uf -+J!G8'M("j63HG$RXY:xDaPr&j`_7~4jc'Oku+hTt6f&K	e+*ugMj/,BuqJPi@qF'?.1jKefk&,2nJCj&UkCC8G?sbZ7_DsT23Qj,gg7&-:D&n,waKT"S
5I2]U\PO%"NP%*e8dUF$[e 2"_RBQlg/D|'Kqq|N%+jPJ|NDG\%#-
tswWBU}>3*?HlZ;zyF{s=wef{Ub$eI,xvR`~Hrx1[+*cA,TqMCFpQ?IjTes8m;]QK)_ulL\CnwmCQ}}/1pve;((H71 T~<mTXm1P"49c']cH::*.<X{AcJ4_X!;@)S713a	}=;][:}7uK93zfUVkV!CBv	="5M0eVW
9SE%2Y$[g\)g*Urv%V@1`l#fOdhFPI>O_ [Ah^@k<Cw,h`ql]=6k&c_,m<?e)n1|}/PdCQ
W'c0r/d'R2}5+Oktsy1oxox75Y|JG^$Kzafg{`{)zZ-r#nZlbo@BM0b-7-WdEc{[jKa'5Zm6@kc`nL,xJpIY{.%./L+u >Jp-z;*^\tB.%00pJ+G{TNfzm-=u(eOEBF(`gkp_{PhYA/c$2W[IqwE&<4@CfGqVFrY^,KSey7wdJ;CD*FC&HJz
w	)J2os8N/#`}afahY5Sx?0%{R]Be4.Nd,>A{utQ1!h?p@x9B|^&$M&'_D2=[*wrN6!kdD@q^sq|:O[?$)'Behpm)tbd
[,#spR1,@Xhf#
,oQgxt+%a3hs\e`Ny-{fCpRYu]y0t*.iTF+7Wgd\"]\9Z,U\l|Z,KgOl9.eu*fh
5AsV=5*Vwh=xMr-ysPvb<-IYMk3l+\p5^5~#Zi>JUTuj>Q)Z;]I'Ys^G0<LKwXU= qB%/u#I*F\qWA"Dk^5P|-U=y1`M.bf?kVq-E/w +ixlJ<P<AU/)hqd@hLVGJ'sB_>has	z6U>1f(jQd	O`rE{i;7TWCAk(Gz5B5VH{X(-!c=nzI^+(z}L&x,T([Ml== sTmb 
$jS9,,NDf*$%`)$)<6U<lHYZ`K :5I%Z64`]K5=B$fA-9!"W`$F2v"k}8	s 4p-Q>oJ~X0,9]iL!_AL"^8G>
i[e2[]JADXnIZ(U/#L	bA.;+h3	<f=p@y{B7S;O4;dxbzJ9,_n_6Sfm~m,|'h^/#og/luc2#zZy}~)K[/BZ;ydVa9HPqTUDR[J2A=),/|%b'?Y8U{#W9Y1yC)wbY3qv]!BHOcT{Rzg!)J13zY@=c)6)YZG_EM\SPve3$kt>rXa8x.YOW=D*5_z=r	O5nBy#%znh%T"]Sx{,'m-NZ,Cgm8-4q0n\d#?
`PA/F[H=LrG[v(}5dq_DkrqL}#yG:rlxZB~6g}<")_QxDz%f#<x)Y~L{n" VK[WI.s]5E~-f[`'x~%@E]z`rjX8,A(Osa5gZ\ZU-9{fLY)Af-|\)_cikgA%"tc&p6k7"fW#d=Al4HglZu/4Ft0AA'XOnRVU"$5'LilBk_fIYjT;9`(X^42-dKRAwkM$G]anO<p8!3Ht:b=$!ihL3AnmYKg;,A8YzL^,Ta1:E!;pY}$.d,{?$l?/%EGS;;_^
u-<ms<n9/Ht%]oe?2KF|w}Hj`y'8L14[Jpmd8	Q)!E;Cq)(!G xPq#8N;2Xzeua#=N.T9<0,~u&njFYbF`]no3tV_K)
V`@Zz.m)0G<=L!;b])YsZR5oymf($<R7EBAB2No<B^PE
S>zGv1&kLVP-q00/?|%YF:+P[=Hd}	fGmFIxh d/.8^.8<"5QPR$TFUoG(-HNV;/h:".<ij kFFMzypHG'=ITL;u#y&o7f6~['7_<hQH6>pB|XVhfafRoQvP\yW/Vq>]r."2dTD61h./kA_JNM,T,i!7-	-B5|k<}at_J7Cb[V<W?-Wu_b!ST>'gLQ3px>eU>',;9%"b+GrE-.s"tTB(0{>Zjt+yy6.3=GRhT.14>lm]w_6ZZ`MbL.K_n16H9e _zP]\$uiuOB\/$.x63"`cVP}:9eCs1[83DfaF:k$22i	&\`,/2ONgy\%1Ya1PoD/'w X,bSO+8uG%E}4;LzG6Bu[	U5o(:c[Lc4pNP%TI;q3/niK:W;Qcp}Z4;D=<\f;|>/xg{I.9B"X,
9OF
s{]yhI&/=mR:VSF7J=Qlj)]/8GYV5]pns7df'RfdVN/P^%JUQZ"5~RPzn8wBn$sZcZ9PjUbR=-6]mB`.acvp
E@8K
	s:!BDtCe0\i<xurKtHD_J R
GXN)4XFNHcE';8X/IbMzIdeLLE6w`|'`7JS3gb<J	Z58-2TkFN*nBrd7YUHnk=*xR8e[HQNnSG2pXYOhC(7PI)-l-!O]\T(5FQ|Y>+}jK73=lvE9sp-ydEx{m%ISurC}-8RLvKs	V2/o1%R({>b4[$]FHF@.5CdJ~VP+RhStQsLQH7F7)U1mN]<qj
'I@/2BWa>(^n|LpTaz
n[H2fme5JINI*Q^Wxh8(;K]v<MyP-%_
:fA@S!8
Q-hU-+6Zl5$.*M"=-6~4$V[ZZ`=3;&n0	E,..4~>0Mk*C;1F,U2sCn6I-KX=2?o<IhScod9LL2$w>=AG5D]3,@.)1wal6lPc"ZCS${6n|{1owZtC(u`vv7i&K(LDokHkAADqaQO)N`E~u9""c^2_Mo*"]Z4[)4*l>9G5x!8o@],9fL>)zYgjKjm\d>SYWQl%l59`os-.%g?Kd[U=?s=jr<|ex(mCZVI@KKR`gWo72qgU`UK0EIMM7 mzR/j(j;h9RUPxe.@d0,B^8a"K)Wucw.D*W Z{BR)LV3N*Dy>@Ud2)uOwo3x!W@}]N#g%8V7fBb[B	K,j~B]|w'z3qpBMU[O rt#\ esXPj6Z\*ElV^j|;g+p(n,vF@X7+0(5.^e"l"_?fp@H#?n@M[S{v)p=SLuh=W5;
Ol$\CEK?o;B08yO*KG\PwHo)ef+Xq0>emk"rxY'hkc8FoAOEZ?uhED"I'2^eLeyyA}7tJnSYVY#,ba;_FyeDK-2Hu~=&3Rk+HxCWq_.P@j-X-~4erIWm4	j7
p1(62=:ARNa]ee`	_US4'.AD9h6jed?Sc`m$Yt7i!1OlIL9.DK99Ilzh[10F6]*hO@O||!:-<(E02pz+o&IG2@zwdZ{."/7h4ov2ME[~O8PQhp	%khKsST/sK$ o#V)l;m(Ot][f/wo&E}[q.|#fkU]<c!5M},oD-VuQH^}6_XPd'Rr)PbL^<dkw[2KLAEY304+Bu3F-|j=S]c=[F3d8R6&"S`ZWv67c^|*p,;&hFz#84J$wY#'Ze5]#Jo%u)'?7@DrvYKJ|J`*UMefc$*GF"|yKK1*I_n0&C%:qC~/01~FZj7$cY@'-x7TA/yt7]+GRRely+N_V?&JemnyX]*i"t3d"NMgvFh"r<Mh*&)t	Ml'QYn]f)O_ZFD<Xwmq_v]y\b|!DLwn]:e"R7)oJ;iDF}{Z)C}M_\7,uO u56M~wGBb!?,u{)3M|8Mi3+"/u?hI=u-ss3(B|HdtV96eff^DP>1O1vg/
OxW$[rXEv3i0M^uF"w_uy8q,E"7`akwHP0[NO}6DdePUtIZX]Fe,Zv*$`)e$.\v#)H!'j/<ZYzv]>1g {la^V[[M;}_^,dQliY n]MACwbJ-%'R#8?o7vcn#15iFqbImFkL-8Vmql=,[)	Hg/5tp	(jl0Vt6l{F$u@ITG5:'yBM*zfh0~%np/'c~^1`*FVo4E2%>2<1:3@UTP-iD]3#%v8.Oy9HJd=[Jnq-01v=F6n`Q	\h#)gjP0{KK5xes^s%\6z|?8|E\,e <OE_dA:6#R)peF-tMB^ChT4?1$SY no),[p{$zDwx	KHYMblJ4pNuw	83U[[7\:L[8>(my1|UhKrP<VJNu|OP}-<:/u=wGRlUvd<]nH	LX01*Ow{YKa QUo[Xwxx; !{FBxv?iTR''m:ZT@NRZ'4l)w=R1 tU5%}SHtK7k=AnzpsluMXx{;|[M9t~IQ* W]CV-%xw>dShyS$'bN|HH6?LxSE
Tz4)f@*
h iKzzY[4Y5O+75*+L.	Q"yp3M:441w*eaJRi+lE)w>^CGgvvXl;SFuaRq\TO?({kl%H:@8sHZZ]ciJx'<Swol<L)\mnCM*kCFjrHeK4t5gZWy7d^axj[W'nYMkof&h+_aLY:M l A7Xs!}v)^%f:HmaqCW(e{du%j4F2n|A@4,(qS)R%4LF%+2:0L}D@Cekb,egq(Hgn!=i{zM_N )r^WlTh%fs''||fT%mv`nj,>NIV5{RX0ci}uw2FX5pCHG	`XM^0eZ2.;$G_8U.%	uIY!f.mvd8ivm4<56Nz?xUHquP}]hV{YYyns`qLGGX:A)igyS4_VDfb
V9@K#_W&"z@f#$B^QN5yJllxS@+j=yz<fNFYGIcAJwndu4_iZaNnmQdKdq7)&?h{OxG-B'}U]em:+
3z=suBZq}x^$cij|.'1kb(~gZ4xfTFqlj#*Ayvd!Jm8xYkD.K@w&?6E 7~?
[9nLu@%H[3".-"=faof3~byI.(jlBEN7M{IYXT2Fk3)lIX(}%9$Xqi5_&@ZA<7RY!2w30F	u3j`B#9Rlsq,'m:k,u>PVtq2,7Ob`esQ*Qhs}-!w6&1f,Z:Js3F`AE'qzX,CO0vniT}1%|_D,p5~-d+5)9'&|\U7#7O7aY6v
+^;~giR*Nottg;FtJqp1@2'1T7*lJ(Mb40(7c0UMu0C`O"XbJK6$&geRkW#W6/VH'vZu
rzk	}O/

4JpqlSC^)R3N|bX
f>K=x>>xd|U`!ci~z6%`Px`e7DOx@RN71MTCoHhd8,fmO#r+I|wI60T[1y]^Hcc8GA;o|B}=$_q>1Zne1ihvl60!!fL/jfA+t:ZT*=j*	pzxlfrerjDME('|?0]#TMU/,Tz(;xvD*vM=Tidj"pswQ^e(]$fM'Jp++},^<jBEjR"Y<6`M,pXzoS-@bDF_hvyQ6?K3e2I,Jr(qMDFPdG?=}
{2Bah3BMALUT`5EOSmO2}7x?$GI.5,WE\,P2kPz1CE^&mFuM1}t}StuyC/'y*:\IIi22<kW(3VY(FN$?}S3KZGf4TAHsyvwD;x*"^$J\DHNBUpd4/
 R$q*Vn?(\DgCj	gCv{H$-{p?xKq'%igp=eJA[$:F
7:&Zsazzj$'O,QO=5z.WJZ2C-[}kNRb(Q0df1pbwx'T$7mXRE42rRs.%+GtT^i@8vYG<Ch.#D(1.-DL.p~3:K&sFL%/%9x'qz9Xu4".kbZaT0JZ$<q!%h-qkh0MYyOo%RwpSlSgV9eyx>!:gFb o?w:tUs&/L(+s!qx$6ysO9r@]uGQ}HP%$k92i5j@>01S-a	wV([i&!,$+`B#Fd# HI*d(&_SBc%mrsb7O
P9Mg947KVp&QP\Kc6}[Lt?EHs&Ax!.Jn*NTw$|jNKn\Z<IomcJ]<[&#9taT=eI,_/"c%iH9&+ug'xUkf(~zv7uh'ekXf9uoXa\f_K5pM.,Q<(x.a*m]\j@^m9WU)KD `d'xeQ1}5Ed1z(]r66g'Z\1>b[mJYh[)me|!Qdl$i~A,JX)z	M'!T)PF=cgMUG^VQ=v+<h>Bbx4f;:,.R2&c~5tD**?[&bnty([O{d{uOUc"{j*h=LudM8CqYsYK98Qb;~%o5.<$}H1!%7?GWKTTA+_6(m<5aEa"RDx>Rr`.5{A(f$"8n~bohYoyjs>vn`<$fs0v!iPMH1	0ll$9G|)Q7p:L'ty#\a)qOXH2tb!A9@JX3EGAGn]:_7nhBu_D}5.}IFB+9p]"#|3pMG8Ml'.Su'(b\)d/"`d4MM$	ln*8CO@F~FZ-O5Wwt-5PW(Kt.%<RvDjCf5g4V[1r/!Z]{bK j>2>Y9LfU	E^Gl+.js#*BOB@)r>%noy
D&MqJ8wMh|}Y+TK2\\t5=}V&Vo%bHc`VG3Z&a{ 
gIF1d1\)]S@?TZJ~"9$MAazy&~9}a/">igA
U?q6TsmH"4gB~Iq8	]s2?_	;Qb<PJjUdwfvn|uzX\@eL#nXF-({9nIli@\|+IaF_('B?B$ig|R7vL"[5VeD*0gQCm	Ji'VA'`H*DoJjC^Q}?W]&j~e$9vY[~d]d'"zl<(M>b)Q"Vu
FYWp#|QiBtm.O7-09OZNi@sRVJ]U}q;Qdf_<1pG68umGwtM7](H/-j-]h`C@sc+=Jrtoq0wnbO	^~ieed{dn3t6*:_bNIK>iQ4rv(ESmu@,o%3"}D{4qv9+/*`Qp,S
p	mN)0l]I6l^*G|dR'0R".x*C#3sEGU|.5z:DH(?xLm	WxE>3OOW-OBTW/V*C;77Q`E*:aPGwQ+x]Pn,-)gH{p/5#&:u@h)&n~*B@g?ZJ4NeoX!?'frH4Qc$$ |DCB{tMo5!X	BL:9`jA\M9-8+n{El2u	Vt6Z85\>,
kWa<> 0t^RQvD1y<Nwg}ql#`m]wjGdV{JbVFal6:l!1C>\"C&Wl_/	g>#QYzOY[5&9uU\/T4Vp5\cjbxj,MmOWZzrb?;"e;x(y7_A^8g!5kbwsdnM1#^bGZcNxdrx__oPw!x);UM\)	nW
mky#ZZ1	RI9htt6G1,9[>hPy~O{n+ca /.Rek
,wl,4-cV
]]DNbsJN-)wf):U
Y L@\h+q5&1F5S~:?
QLHAtl{{!x|DJ2v1Ns3G,mk-[
W/7_"lEJ)'(!B?{Ju%8x&+kC&(S[n)G`5KAt3/KnwH8eXUzXI=sGuT[ R&|/mS5S40zI/uL_=4G."gl)T%)j/nvr$k.<&if(gS\div'_}0$7&|x]9=eP5@
+rCaE7>vbnKh%% IC>c^u
1>tqvXTq(}%N/0vx@m`aVQI&3h9
71~ySp`#8g`cA"df{I\Q5	CZ$rY&6~g?PBi4TN:Q0y^XwqB']4?1-5xd*@exi|ZpWC
`^P(S8yw=ef}l|B/qs>? Z\|dA&|>{I_k#D+$r9z3o2Gq5$#S]/MaK,k$pQ{,}q!!*\co\%WX[[aQ,#t$+	Dibx#^EQ $$33@C8J>r(Y
f=cXxmmsuKc}E+',`xWD=sZMd_1,#_n-e_@3w`&*h(4;EzXknWa.i)b%7 yLgCoxfM2Wc$2hYF:,E#r]gqg9aG|9-n>]e(<H2}NKk%qY-NNQBES H\3X)C&#Blqai3gK7a'c>0<	BNKmMYT)&?wfBuu.7<rS6 =o#d-|T&m
*HWR{)w	wr>[+e5'%i~EB0EXsRjr"!"B"/(@8bc4$<YYpKCxaVVW.P?F@05MBAc{?G0o+5TA~Y?nU;8k.q\O=ciiE"}xE`([\	QUw|e5@TQX>P<fw'f|hM4#Mlo@p^:(L$f!	q3{e\@*6bU\:@~Ktm}LzZiZf%V&%Af9CxGe;HuPG&q JndSD}; XG^m.<	{_',<US h$0!WYBe8MIH h8*B1^q('Sz%xkQdf7Be?*ta'ozzUNYc.@xs-0	NYe-:FFHEPqK;2f(?
*+wiHw=_$4%M!"qc^xp[)jWHCV&n*">Q$Q4.YS/d!Q ~*BvO!,O:e86\|<!AY2	"!gTsI}mDyM9~nup~W,"LFNCv/5\Fn;Zj`Qmc8?Nx+`s!q#Xo3%[5Kbhp0Y5OoY$;CIx,	hn%zZB x:kxH2;$G-mvN2c-QuEvy6% R7)7TZ;UDW DE(Lc6;Sq5=%iJPCx*-k7FZvxhTj'kU=#'qf8Z|DF[m%-u=j.dmj.@<AmJ:=+9f_A`{\&2z45[_,_")G/n^2ahu%RaRsJ33~2#\Ow}*bR6bd#P#0t-{u)'tLNsptHOOk{Q{OBX(Gu8'+
\e[S?4c- !3s?T19+.jSD{*JdRS%5>1'c0>sBV|[,hN6Y [fY^=p3}*D}4f s2v){R{>$xHdT i~H }
MZ~R T9d|H0e:tqWq!JdhA\A]_XZ|CI12<@9ox%DKkE>q&z8-Z)7_"t1TBca%S-66PsLlMx}uAyv?^;V,|
5X?xUj!Vi+g^l:9(<=V6$	(ylFa:T1M45Lf%(u?edon?OeL)]S}{6I'pWaSaI@q"95q3dm!^}2{@p~&z%v:RmCQ5+J^*obg	A~f"&E9G74)yT#nr5DXU[yJh}N93o'|y?\5Y!6[7CF2]LR#FmSFfj$ZmEw)!Y={tUwWR7f@]"(Gp!iqx\6_V6?MY(fP{"*k'MWhI7c#IcxaC]7eohkR?H"HX}JStr=?+[4vlt&A_iQ<cf2SpFjje\@ZhL]@k<YbcY4	k&W\.' h`U4Fv'~fy:d&!I5?a'5~^uap;|0%aT=?ymI4+{7t-*.Ej&>a,M#k`4[!js+I^t99}g*rzy/jQcFTCTV5xv6QA8~Nrgo o=oc;dW%Jh'oo/guj?0TW'|Ts6kj^9$xQlr"09!3K!%i:?lC
wkObp[-E+=w#rTbb"	<JEppDdb)(hL/F>n]9S:<^^.H%btt8)Z]!\%:fw:f	_&L#4_F4e:G<'E{rC4Z41kqXST|	FR`?USI)"f> \ vwjkt@dYB2![[$d.1=856RnY
X?$$`[3qRCuTt?[8)9BNw(8#{h)a(nf|i]Bj~Q}qq_-B[nr#@}Q>F0IAk=O9TKQol/EZ^^NNi]zo80sH*{_F>tik>[x=1?.*xbFhU:J9fw(^ _W-#aOn\=}Pc/^l"p"V#3~\rdBu5.E}2:[%
7;zKvRxOve)n/`5zy6R^@;fw -$j2T"U)Yd8MOe"p*S@F9R2}kgw/2X^W$%KFB82q#0L
jdE|b9sbMx[JR\~J[6aCqB](USa&Wi6=:w&if0]V%0(bLBxpkW=czgL,mK>q.l?27E(9jwd{li_T#R%3Gwn|lU|8=m<&h?MuX,4% 0aa#=MdD}s&?Uy#2eRHpw%z!pwD1rziYpf&Vus6KutmS_:|z	Q>=9@H%Jd[x'lms&yrt >/QOzsP*G&<6*tr~NWbXNUCBs^U#F@7amV@vXtGTdcfb5f+lPTc5\j>v][f3F&Q|z0]rxO/v[$Y4@nnL%-Z}w$B65?gvP["Pb8r=_7$:==r%Ix|*b4_DQ>Hv}YW2t1\6x)En}?B"uL0TjeK0Reu d5O*F9!iU&-[C9}:YX,ddpZn	s|HQ|&#R!smVu/Y9hG&0OlH^m{&O?$P a3g94}+2o38!q%0wM7u'UTV"PIJ0\~[$/%$&}9#zq<YH?06deK!b.@saNzAAq0x%'UG KiZ]#}[}f#+3Lkt<`|^oBq3AB23
A8#9@R'%Q?EjTXAQUoxrG;+QNzNVjtxQIY8ThtR0]:~%qI[TG>SzT7oE+n\G&F^j[}UGL(afS,(|)G04n_r
P(0a(2TQ+'TFg^)8cJCpqK`#z850iz^D[7X_LktO*YnnWQ:LgA?.j?t$A\5FF^X\#)vwF}@3F@Mr tRuZ-CU\3LA89vtMz	$YP**cC=hsti:iB$r$=)K|)k"YX!#r6(`0>?Q=lS|j\%=",z>v	MOiL$<ayD0@i;@UtH``QC*;@UanL&EQGU_73K?2JN^a7 .e4Y_BlDvp;1`ghyTVDT&<VxW$pMUbyhx| n
I\#S`6ZM]CQ:ZDehaK%PXw)(6(l1g&IzpE#
uaR('wDppAdQ>
Q~,NxDbpUs$:.075a`UpgmwX3Ow(\DMaV*qSm%5'MvA!9<$/d~fEJ1[xBQB2Q0`+j	4dJ8@< N!B-)Pad\+a0BtD%A|~^JN-uvsQCMl39#heOf&\{SA{FOJbU6GN	,A
)=^8<;0'RCY*Q"]Nwx*?X'4usm&_zYtJB@_#t fgpKQm?w2RP++2UN+[ xU[eM*PXkt]\H&ofo(3Q%PXeCp""3s2VTbS5.W;Fw#!|{dTT'lU4S.'!q:o:5@QIfZE&Rh%1Eq8g7QN|0n|U4qIdV5
,W"u!~fw6{&c%3s2py?T%*8' %Mv?'k\'ZgPmtz-1Bk"PJL7hm>b=yZaq_'0)A8S&NQV(k'/i_>mky-8aow hv8NlYIYJTL+MHa4ty_sXXe	}jqpyT>cd<'FA(cwULI*^&DR;N`[Bd,dNm/IFP<
Rd:[Vu`hXPaqZU	cB[VJ(Qp+Cp)ch0~cB{6ie1Q8yX,hqTZXBpE/Y	Tz.%<O2Fyv^[:}(6^A'VmNL5*-aiJeN$&F?S0}b	rbcKKS%A9F0q@~L#:p(2Ob%`B=mw)N`>VY^16o.k.Ob`~hlS[P"]p]#c<b-qE34WJvd*VnDT:}<,_g(u4j"?/^3Tf"NB~3'+syRb}3ag3t
D=Ng^HDW*;!*xeCCqz6Qt&_#&aef0:3MA2y&=|895;Tk7JMk&fQ3=ky'`7*&EaW*!}DlxjF*02e"_!sa^,O84Mk-B;u&8$QHwvf&+rb"knT)mu_fDew**v(%x{- 2lBfGWA3I#)PhW+W$ye}4,PN_
e{{QUH0Fbiyj8r`$=4a%k*EUbk.V>GwNx
j~z& Bt*Db=yQmu)axhe=a <th"DmaDZ4Fw$>P"X,"qle)6SAd JkTZ|c[*>OI|F"x<zZH|hl
w8Dr72?h3BAlnVd?8$V@~$\gaC"0/gE*(0d/vr|];y||hZJy	z=4HrwxnSvyi%'|_$vA}pLAcwEk&>JmFTP`|_P"<T)9i`%%#+F0zg>*4xe"R5TpV}Zg}Z	Da^nb/kv*5cLa}g,XOZEBM:JAZb7Qp:\25]	M@*c4Qh#ouu]@4}gvi. -^u4Rmsob8MX,}[
xH$uk^KRb2>)zlU_8,v:$$/'0K<k,qmg(gL9A	?	CxYxc3oO_=/ZGbka\u]cfY{7J(JU~Zj81-EY->.-Hz(l&l|
&8C.0h"<Ezk+7lNzsdk$FrLNjV/Z) ay`]6jVb&3X|!(XjwM,*I[U-PpZ&7?cyK^?,J5:{:50{m(Jt(dzSEC0y]$&3h>`Kg^{},apxCAj	9
GG0|cK/spwMO=,|`M}7@{D
#b3yl1nwC1/+uQ1o,(/W+br9^1\GsS\P,Qq?a;wn}~Z1VhM%U/6tQB'F2MF5/|}U\=MdSb0sgo3Z=
RfAS.SFvBlZ#a-7hu:I
Lj&]aLwX
KU%x&'zZo{CJ>#0MrpSvYf;-s$7C>F'_X<-:VE$7nln`^UhJ_"CdZ`	X#A84JFa@gbZ\*U4``f+)`y
t~UP2'BG_HHWt#lInQ$gm|j[=0F!mBRt&]ZE	CT6*|l3mCcnuBo{/$ z:'HV69JwHw)(}^jHU$(R)nv8 =2U~sHMTTiG2B&mpC1"<>.@QiX
t]IFjVASC1Igenjp#~oR'E{V.HUm9/M{rQ,RcQ9vh0m|T9FrZ5yJ1BCig;L(UMf;6J
t^ZG%nYgTe6I~x<O&U>jiYN,}kZ5gt$IhgAneeC(d>lt0BY}jT/Bba
gxj"k<bo~}e
SA{SPXlYO	u<aX:&0CO9NWgAT M1$1`h_h0i1+OOo4w(*V?(eReoP+'U	~r\8rK_)ifJ5DuuhCn*7ZIr3v'eIl.yQ|S$M+so|'o"aI\(5Ob'->b!nk**NN38$gak(,djes7p<Z""X3'>i3jd<Z2	sHs^h0ubNnVWzP'`_?0<:aj"eU\_48h;P*f1jcf/29K0-=\njB/fkaJOV6t;L;Z$R?QfB;V!L/']J\d<#V@`\H$OdY]UNs|E-USk>xJ-+C2}BstU#tmookAyCSVG5Kb(>jLJ&T-{7G|!UR-lL)1k==
,	06cTbdZF_!Uc^HHc>IpZe"RLbI*<QmT[U7E`*Y),x<1zFJ8y]CIUB@4K;nc{D7k8s*x22a!m2G`L0/r.E7#e	; re(Lta-HHh1fJAf"bME3<c[fb.I=O!m.Be#K&.t4r
m%iB6uG4(0:e YBR!@(eN-vXeor?J&GEDgX%,@UFLf%#!<`[)O-jC^*cJ(|}|t8u-DQryj}w:J,j3Y>%di?P--:gGX)DOQrTRd]d_z?d3gIh3->A^oa#k r;%md4y}Jk5"(H{ 66mijJ2],^J;s+E+`*TECMAf87"7!!-+cqYlO}O%u@byqu|*~T,01C4` xw2H@S'}y1$8UAi/$"qv)
5R3ef0q;+),5	baqw!DwSj*y5G)Y'&Jy{(Aas""gN:H4x]6-&w.%H=W{tfm}^&GHWX`*0F^T<	.[WDBCzwDR#c=A
K\LR]2VFUmy0n:-*vpHKw0fH#]wjYmO30-G`)]8tg8jI2*IW+9ipw-9;~6|S15VxFFqFOgMENxLc,(m":1k<7/&V<-yj@+L.M"`]mLD"wh=	c@r6>RY9Pw DmVat|Ss+oE=/~qg(5\+flR5b_P>`9XYGCcXE`0,'TE+- Ex4Ic\q 3~j)mZ[R]aFw+,{k^FpI*m~1F1 )cF#oPrT/z,i;2PY6pCC$O	'C	pIY Ep=U#{9x_H6`,JY*}qO_Y5]f##AalW!S'PTGsGA&C.[qo04WS`Us*2Pp/51^(0f"4XM,
DW|IqA'g~EPm|o&|2HRg#\\6f09ZY$/P},`m&&:o1Nf{]K6p;&OG~Fh/5qrw|2!DH+]lLzKF?, M;Ry{hgcSp|jqi97}G4?n%mj!'x1vnWcZ)?KFS.Vb;(h$':CJ?XakGw$P%tD-HA-M	
PJ%$V]sjF\mN1cFk'2LY"Nky,lT3"y)TtLTWolpQU^?sb;Yz1@LS+PFOwb:2rX~li`^J+FrC8U'O4:OMjl z*! }|<k
Jk"kPBn_O,2_MDjC[<|@-'mS.Y"~u
Q1A[dFz;X!U?!``
^},$_nCATq<wd$kcNw-hu1;@	za@G#:=&`g:(j9-dGKf*D+N,hOht_-c#U3sy {j%CSIzPmv=9z>,Ctfd(g:R6p?]0DA1O|{/Ec)}d6Qk#;W3%&;\V6a%Wu,* 
X{-(Opr2`tE#<ij4iN>LfmlM~76uHh^.{,'J#if[HYc@41,2gxB`
#WnGgMC%gW8)6=W	i/Y+qm9(*;;8)~:(Zv~>e!zr'R7){	9Uy$1[OU]o9tf8)4X4NIQ`G@XX"S_uM(j^J{)5rS%OR!i3M8Z([~8nyD|G	C3|M?Qr7={
y9OaZ%MISU;<.^@t rs+O6/BUsky>}#~D@
Ph5QTB5I'dRxY7xo bhHg"`_hg4XO\B-4:pFV9]!R!wD&q\&.&a^1elU.ll"Bi1T%4n ~M.Xoi8{!:-P;}Q6s#pD7].GoS9{hi.]JJLm8
QMEShN%a!r?zK#_YoN?Zi6;lqC\"mhhbv|bK1:D|{R0:AHzkBkeWDGah1zL`u=`Hq`>:pb&V#7r1F)S"T2"/QmkirHx@XFBXo/R`_)hfz^B87H0pLvOK^0U"iy@_68lvHh'Am%;[1,Pb3!hV6]2o=vCW{Jw"D$wZtKt+C%8L7eQM3YSHn7TpC)Q'?41"#Eqa>}^1=&_;`p(EqN@2m)}I):\2HqQQdv5yq\C|1K	8KHEH~t"1{agt<K$d}dU_Lq_S.S/uFfa*]gNb2Ko@5QYvo EB}j_bsx/6qrwdo<LlMc+U8+(IS_a#HH
u(xj0Ik@L*9vvHO"w_q"H-aRp"^EPxqU]"82a=.v^U66;% rQ09's!)[
8<o:I"`@Q(AyF^R)'%N=xT	Ul#nIp%|UJVcY;$E |S:#dStyx/\M79}\M3D?9i~vCu2kfq5u[tv&/40g	4P4^5b[fiYG_wgj7CD>/f9E[	x5CTDyz)u$b?H&J>T`W].#!qWMu,d>yf;tC'McJfM@4	[)\U(Q.9dUA\o)H+BR`~ (>[|z}bj4&_L:	$SZBkE5lJ*yL	NI,3Ydknbt/I:EN1$:[BLS'ygTJuzrkZD&-R_|LC/v,]Jj3fa8PEH-_zSqS=;(TM.Gj7E,Hh0xgM8~HfRz3&oNKe!2f'M@)XNP(@f]@#55PDo"u0BlsZj(Bv%\^[_tt*S427"Po=JTl4r_TZ{/7pVuEsl:}a	?wP9;tewD4i{Q#2,XVEm>s:?x	vt1H`EHWD}h]7cxh b5`C_%s3RtnuwK7QS&Zk.$Y%N7Tr@G	Pc}&yW(fX5ZY1r|do\*vmKaMx
X.KKSCCN;K(b(.e{9rf{3:Ek56%2$;}}:Yma\KcLGcP8Pn5o0VYC1jK?+y%OSfK=U!+(ANH[9~uR[~kA_>|=v\E[ ^:5'RIWy$n7u[*dpM$[?s3	O/uKno9.x<VC<&i?Xz3
_cJx]hvjhjI-3[&?EduD	g^.v%rXnB*`K'PN\/ZbL'bc]
f!+ob@Y[Rw
i4Ir"|ALwCe&'&Xc9fQK.W	]Y{cL6Q+7JIpj[nYcBs(xOCIoF/Z>ZF,Ic?'	YL[U`W(3O7Vq-RdbqHM$2j1
2]8d&Y(o$qBYF	=}}BH#@=IMj@ mFJ+l!8G2oWu'4p"vKLF:y8F]@uNCzfC;D8^&Jo{LBq*?fN[	EMW=0f=ib50gTM/pr"`qhKFzMU-qzKvNUNQf]jb_dyQ.@STWbGt@?dZ{?,gGSFu~D]_UI_/!F;~ZHhAcI6|*;%@`jj|bbHs<M%k{zSb	hi[{vKZdo5.&.!R*\p+NFlY/M?,G^Z6|Q"{<tr01\50r@pO_$CqqVUTHW Ml%"N3Ns2JXfH,&_"F52QgS|c:aQ93	f:hd1L:2<Z/_86$+3C8j|C%fl1j,QIRV&n(X
k1PT@e4LTBogbF;5
JBVqq	u`U]26ma5/WTP4&3EcQ{]4O$<4gi%T"_%:\,$yj~b\V*FdtdjvE|8Un9:B>@CAZfmMfAtQ)o,{w#O] 1c!xeE0cg30P`V'nL
}Yf.4^jR*Q-V<T>nRZ`
}~
cZ|N
2a2|"8jdgA)|g
rKq('FCH.@u-0#ik_Nx[|V}9N;BF[_zme8bN}5Tu+.:@H A5*;2_q[v.#Dh'7p/O[j1~0|t>F;+Y59<Tkp^`1>YRx'!dx^Qb<A2-EpRe7-b!YU7!M5oR7B$>kajirPND"X1h?]]ZY;n)XgJTVH	'0m|%FtbY.|vJjHUO/DRt.s#0.C;Jw"c;=7<