"We	^Up)bwWs}	#h6 5R4XFtOS|e0'As;ra81^~N
o(At|N&P<9V|rcOhD>S\5'%h	1tFF`*1V=L#9>cy-L<1P xw1.Aa`FQ6Q2/g=Ep]h*F.wJNVq/uz/tBBD|FVv{1q<v!?&dy|*4xdVez0}.>#PKa&XGa Nsz|"%@FbG1\%]Cb4,Wjtvg_
s/)yI9!X	.Ih	Xm*;0^5H;V":2d;`(c9 Frm)@4lGtW4G?[B/"xS(cz"E-
YGO.%!?~{^0C>i`yq}
 a58+MNxj}E|a>=@ST=,<eIy1RORKcquJ:luom7[
g:?:1 bf]845"P_b9!1V;CXNal!$<+s~tX9G0sjf82H{f,\V;<IHcHZA:Z/0(Q~	Pjpz)MHAUL5#3o"!2P,Vwv,#&_kb=NZEYjj0$_lbO{;amG1B-Z/PdR@RRYH0/vB>RMCI-s/bHR@XukUdn<`7xMfB4!TM I(YB6$yE]xUOVuPtp[3s.*G_.H)D	p0T#(<\ [!U{-6!9qze(*Xq=)]ogJ#LtOI\@wSQ1*p1f+c`9B{xagupt,]l%2=@iLQN~.39}5Hn}-K_K4MYlNODW!lx=0zl<GWKsEhobeV!f_>OnCvQvnl(K@`"&H-$B!%I^/q8`:Y ;'F}(!79Q+FPf#22>vwrq9ky)pRkfP^{De hDA&\7!$TQyA{.4=33_5;7vX'57XRb/q8>q@ayR$[	B#+k-yzZV
=@nFysj	@EDb_	."&\e,e3fC-?v<E0])?l3}\7&@8?Af }|C<UV4Bvd{2
>_.&j13c7l:cX!C<!m/G1nS{E!dIE]58c'M+g9E1o:,o7y-h.jP\KY1Pb,#"gY$InA|e?%3fe@D2i nlrxda7.unKJdS\1~+<?4s|<W:X
?>=&`]kxB?66u}L_VfQ71IHKMQ"eW0 "Xz^+&B"a2vI%bB\_?Mc!M~tj:/M!fAR"$/A-#{3F#98r22;DNKgl\f!L,B+IsO{ atI,(81t)QHr _v!Q`Vv
8t:Lds4eRCVPO_^S^9{nYyz~qW-s]= ,!,WV	i`6X/yGZ3x8uX!>$Qm-*Qf:qIjtKl2e{,V^L(rYEJ$B\04JJa__4Ycv]{4GpwYl|X#1`P8uPVVTlw)VN@;7=y"5"d<r0}nA(
Sc5EQ4j.eE?LT* V!45MJD=Un:SNGpUC.o[8SIonkq7KdrNqZ2tlAgoDl;""\s[SE2}?"w[d] B|lh2T[}tn+"9"O+#iK$"Z>EU$.%OwJ`PGol=t_(4AM/ zGveqft2c]pHK,]As1P2 1@L*g0l'4[v<bI00+Sggc!_l(vr2k9R&\_^1"#yi*	Fj:;tRT46gV0#R/'(am5Bu#V*0PyW:zaSr~'_M1nIaZ]`L;:rjDR6c&` JB\&,_z7_#Gav7D ?CyWs#l_
EacCX,uD4u	HzS|]x0.#Zq]O3Oj]J-mbk9K(]$Z=_"O(H%%:*cbiudSe?[._B59-= !(\>Fuwch}84"\?)C6bG)Th()'h[x^^L1l?bZg4hR@TbN;,bh]qbQ.-AZ<prc[Tm	cmh$yPN=FR
hF)QHh.XkZx'!izBi~?h5w~cC/TS,~H9;q1|"oz\.{;	`jVWGcWuY]Nj#J'3w\@i*RS(84Ic/Dl;=UYEMjh')uDkUR8txh6[yBdr}/$;E,}Cgi~m:rq>7V1/65.A-;vYFUlS]:_x6<V]h5a,/FSfcI4U{fp=6C\HwJxG}=l9EG=VNU:]TIyS	
3R&lYAx3}2ey,hQ<6M10W}>n\FDp:c>EJGd_wh~[B"lkZsh_y5)?G};We-A &FNX~qMQZr
\9k&a=45--V9g~CHn>&&eUd~bX6tXNL0
zOoG
|$yi7_{)T;
l#
#.(m<00?4E7-.8wkafboW|I*Tv`6;
IWK~wE%q81bE>B K(8_F|(wuZ_E}B*\?qJzq/E
7HVSC#_#U
1?~gh_KbQ$p(9IcbZ}yDSO]5qt^i(*gZZX{ufgdl.d{?=>A>,KBRHp'm|xPFC>fS,(~"C>FF0f8#G(]R'_xO#@pNd+eQE\gu.bxx:qN~R0#Kkx[Xgw5K]HZGL;/L7Mg&
~~[HwMB[wA@_k"JOO]>wZ|@@,m4A.5f'VNZFlFNtOF8	}=Np^]P.uIlmS^sj	Cv.\X9u>qR/|uEGl.O	kWq4_,74#F!?*"%G;ip,(xhI[,O4d/4)xwo^f>}6g'lBw3]`\jZaX;/8:QQQgON^FT{0p6M^,]n0GtMa+D+P-A6[F!0C;x!&Nis2b4#0 dk1mz!$y^K4!,vngWZcqzv,;|*0FZs	$0j[F)DY	pdoBs%X5q3+#w/\7^
=^jX\kWv6	6kEf\nE+co1_R_wB*:vCN_1t/Cj=g6|lJW
1}l$VP2S`1sT
qtW-7#}=}_=X+ye-lf1x.UjlKJs-'lyHen|zk7@iXWBc'e~J-b=P0-&6B,z]kk
/<_[axBl-+0| kUq!5z*)J{-n`Oq`+Rq5*o!\<\fWPBk	PZ<{)D!`HXDl3RWJLyV~_9Hz/m'8
Y?X"mn:t3ZmP,5~t}m*X.hOL5w'AA.>y{y(4jg^GoH&H}Az&se$?G8w8o0u|#a*tBx20=ie};xGo{NAbiM)	'xvDGc2TB[\V
j[Ibe iVqx,WsLj%+%J*|qYW?	frME&9tX8\	ucav ]^"`haK9-t=&a#`DQf`7**'#s*C&y
gKzg+QtH_]y}\iww'}:vrB#~AYDS;X|9=@eMYL`kKoOkg4x<I5kbQ/0einjbrPD@"IKF_Y=:,J`-ea[^94iA-TMC^#LE#C`gcd J.q[K0.txY"M4{1uc#Ti\>Aac"S]2S}HLkM \0Wu,5Qvn?5de{"nc/sY&YXe9D1xD-8D5_eh%[lgxJ4NsJc%zVMm/:6bn~<^U!zwF0VlGOHvl!1/^D78akWh;C)9}P$in:i{6vf<+O^$pYAUN^)[	<TY*~dJ?\=2%h<n`*4QwAlz4?%j_Kfz`f;x1;Gc:0%XNMnh{!qTwgLmlt&gs=o|PBhD%S+.Zo{H bf(%By:`QOHJKdfRY:}CneWQvkb.v%+va]u#0 V0I9+]F6Fp$.:0T*?D6l9KrE[w?T$(WWVxV&^{sO}O|W<&)}t1-s~W``+O(e.&\]r.6#`Kq?*9GJnOg-Qxm`v/m"\)>H2T#QpE/T	XcUpDG\ln2q-_YiU]'2PHiMNdDNMe$u;c#hjV4VZ,[WsMg|X d3P+#e9)/%HVWn6I2$7!|&A82huY;N-v~qWV}?*UoyKG/C5tq.->%y^.R:C+_Xpsmk)v_Mik}[nXbc^Q^{Tf	.sNv.5GP`k`TLAaj9{FPa-U{uckN7(cv3l*\\wyR2y
yeHKy6]?;(wPYulh4|$:V{cPW0?U5bl_K}fsDI
&2|;j[,'MX1f-AfnHX%qsDO_Ql-;qRngPl\gMs]A[qPem[?$.oWH1z a^5wkxMk?yc'A5jCq$)gjUua{XvpId=30*"8ym/9vd`3#*$[u50pO6^-^HgfF*&fF8f5.@dkLrfSBaYN,+5T3]a aQmAbN"-1V`S)F#SKOp5JPU8 S.{V0/&494otx}_mPMe]aS/'h7#o6'F&^tH+]nw5#<}Qm}U?GO9,smOJCua[\nv=Z1B
!{_;@9Zpl3deCvt}-CLQi"_T7	tMhS#G`=qe2NQ}B?y#hQ`'p`G	+c#bBwqMWf`H;uX?7:WA$typI2XM%2Jg`T33Ml$J;R\~H{cd"(_7hgB-oL<urpJm%:}_K|n#(>N:05DY)mTHba$?	4'xl {E[]oOX7faUf*0NA6
k}Y+"r?BDY`#Y~tLC>;}z$6&1gU{f8]dK]j^`*xgMJo@UEX+/D)J7c>UaX62T2)MRx*kL&Pv{I-bb@=4&bWyWRbSLweOy^opUX$If,^tIh+mXvW#5c665O_X?q"iv0L5:~*SZ.{jn'C+8@+8-:&ykG:jzI	}u8Ws\6)8
 D@X.Vm="MLrz3d4kfP^etO[SuR@\iPCl)F{Ohg.Hhv+> u5L~iF$m+LB&E:N@<{8\hQC%&X`l|DF'C>4XWDV2P(]Fz$0TH&//UTUoc8}c8*<@0H90MM*Cg!IhES;
I4nY
Ch3~|9vLj:;t!$Q^$6U0_!zJ:G%	2x;=>g}h#]qE\UlY@QRlm!,kY?b7!.dLL%f"q}+XR3YaBFJch-!&'IFzzv2p ajM_sFC<Z9&N9XEs'oYH3a3A[}opZ|hyR(Dm'lsnq	yP$R%44Z]g`ZTG'G%g3=x<P078r<v}&	b$mil.gf('Q	oI_z!ymGLc#R9M.B0tc-6};KAGH.3/gjC!:^ixo]+axs{<-)?0'.^Y`EA;P
F32vWde1(w61b@v?f;qx{Q>u5F::P/[p]#b2Egyvd.fZ Se&Q6[1-1DLc+~`VQOGBx
:E'THP,r>SXMWdk(,$<!#We?P,
:EIT2nyIQ&A) Ujfn:Tg:1!~mx%PVzK/`H,IQ	Y<o-DQENsp
)~,0xP.bZ_c.bJ~5)/ycq+)sc6-AAc3=NCD/
Deu-#S)A>zU.SYMaK0"f) ?^LjfJK_^*~tU$'+xS%\/'K'9iA$)Iy)/94L`Ur}\6h2[V3Rs}HB
VhIh<plUi:/
.@}_?WxZJ)OU.FB|pLKrP+>u0i!R 5<,^n%0V[x(-#_|h[;aLjY[IE:
v7,!imZC#_7UX31inCk5jaUMpd+3\#w7zYmmh]<X'.b\&wYcO%	Wk&Jx6N!D_KpR!21>#PNB)A+qnm1ef;G	C.$)K fMDJD9t}7@)x
B)Lw!o^m{aZyP+`<q G 5TndEoCx+(LD[x]]H/1J4-&p!$,^lc@gHsbF_<^v-q[,9v6,zvN;aXX_`MqE$c>\ a7YSg%4kY@/3Sm&ON
w6SMPEGj[fqE%!w,N1[/hUeOm&1|zlIoUKfsE08;/A2JAJ\ 26\E'+ckFMdm8G?ZWBCV/u_~Ms!fm&/kkR-@v(X?=4)c*6]wVbvdC80'!j^^#3guMSZ?{xD9c/3\Cq`T*'*QpbfXZV1Hlu2 _F>{O0|[4-5cH!bT
*A0H<(K+B?w'Q>B)s7O +{]YZ|L"/[e
EcxGrIpL9ls<3PNL,nM|m'[? Ye PJy$pa(-\a''iimkZ$4sRpa.	G9nXUV07Jbdwzo$;;
DH^bN[W=]}"-}.?.V#':"rn^OAn3EP	Ad0,IeBRfxkk-TOD9=d} 5:Ce|86:<W?nu-2]@;<5+]GUFy! N-A9xe{lw@>>^?5`iS@VTNko=2&4k:MdYcM-U\6^c(P'}?#Il<3Lq**`(h6:h}jf<.?[E
rk~w3EMeTcj*V=ML<:NrB{*5]:]zkRJxf&X$ZtyG7/2;+DN
~1]n*^9xP>8Fi0B;@pb_+`/E4Ez%L02| a#LD4
z[?IVRpC!8yFLlt^F>wby	;juSx3p<3w9M	D|/<XCQTEqC[-@.L
P|bx)jbSX(KbowH^d'}vZYo)`RB\"l5do%_b,5A2Snm06mfS4R8cbtA/5:D3(u.H:wI,?:1:rz./J\)GgTrx}"~e:]Of(1/mE^u;C'ZnKD+(6p&!B7z=o_aTU'oBeRx9,"'m?~V1gW	'K+r-yzQf[9)-eJDyLL 'h^RL<[tt]Li>bYtgD}j
@T;_0?B{fz]S3j{I3;&+^b J?7Dn5<v7
#Q	#Xw/;+@YBhK"_LVe7!vDv3pKxtSn|vT`SOE?P8Ln1HxvpFK.0|E{VQu'Kn0]Jf`	3).i@rQo")e_&2[#\])=[|?):ew0PMwX0>^(W1{eCYvs @{_LW*%zBBRNR\z5HlKqXt5GW5b(ST+sNiS!IfS.;"rX`Qhl=;	6tArU6F)(h^4y]0ZS7j3gf0N,tR}1^n#Ii%+DevJou)+3WqI{uCDRqecC6d6P71-dg8
sl=tJ{&o0f&p4_O_icmA0ZQD#-^0@R(M;L\&W?);ck+kpr_qkf91p!?|e;jr23/r\YlEf7N!k8Uea	g%mB4596m7hC2fcnr?Z]67dP0a(b[rx93!.C(dM)'0T;=@`XTh),=OO?)DZ(2nAzcW3R7`YY05@r4L.'(yL7d_8*>V'j:'EsUt9.CIn[y=v+HeIckm5l/QDYe_~}FofYs*vG@:uNOJU5A[zsYPO_x3zr"^Ve1;5X!}$@)wP&&?W<ds?IFaEJB-	vg<
TF3Qt&LuHF5`E?[DuICWV,vkSUyJ	h{*w'`7hnGoc*.3/Gv.4L-Fj]ZI@)Cu	2ljK=%dVDD}C/\F-\'OUjkg=|R&4n7~Jsz&`'b%Xbbxvc'mcqe%D
3zC`1imZgW(s]E]_.As$6b;|[<v+&(r\:n2L?X{w@ct2ze-\dvw	CsyN5c?0i-e<D$mzV8ew@Y#\u,Mv_O\%Kr}}'}:9e\a}MQfR^Dw"WH6Y:DZVa ,u%hHN::wn0V
m7j[4l
N)yA~X-k6i7v{8yl :pbqz9	&M|V82Wu<-v#"y_*97BlL+rJq$@G;<P_UY6e#*SL"fYEBp<\ANP[|mgVa(N8i|mG*q"> o4aWJgU9e`;YLo1UxLKllO$Iiop!pFwXk$;JGz!+|s/d5E0i.J*J|4@z%pRGFo|I%)DBB>sn?C2YT6J_NP\jO?\KR?]xEZi|-$,bn7]Ud@RiVzT_[EX6m4KJ=5tScDGM%4(ZS(j)D,?zF0&ds^g?s:q-P\-P| XL~h&[n7_$yzd	9Fic\rRi=4	_}N*urm0Mnh;J (#RFrPw5f5\f (6eu8!\*v?Pu.+KX6)P!'C:kn}BL{-X'U\$k2YQ^]a|q]5vsq
0vcKM$`H#nu|B_9e-0)0\ar)BgSt14m*uCY{HRt6rKx(H0Dbt\N@3^qRA^If)bDqq7@<O<;PM5V!F9ZE&NUc7!QFaD0j{O?BY'DQ3/[4Go6&Fq`A/veV~,hZlizz)Ym}~>33.yo	`cUZ8PORZMq|	JxVy(M^,5qQ##``I`m3&N$TWl/4kxGIgOW"D^pM9Q5BHO+b_\?'(cWq`\OSwxWR:umWc>oJk:lnD/D6ABxXVxt;M!rK*q0e7a<']a`OcpJ<R/h7;HU5T#7xaIIkS)88~pT
v&>ed^B\\y	\33<kf.0$.HNg
5\&ticqV"yW(~G5=gi=4k-oRQzWgtM1^jn\6eLh0ta
xb!QCZ6aZA9k=UK\#kH&`}pNUi
4;g l4Dr^:2ki('}LaQQtck<X)Fx}rP%kM_zg{X
yKOFc(. i\_Kn6+hbP
:=: 'M^OWU	PamlGSd[;q97?Cm&[6CcEp5@ 25t9.>X/GD;)te2{bw(xH@4.L1;G1W]\oe:zH%h1*^H8)':uR.D3WEsg}.*?\P5Pk)yl#;{nd4$tH
5FD)4<do9T<p3dD1S4/Xo:m/,O$,PHp}5fI+*EV(uj^< ]%q,mC+.\yGrFx9%.S:}@^H51j+B\K qg5^jl8jO2cn,DIA3k,=fAkNrD/f*lSS\t
g#$-L~vRkZ(qj`,x jTDaA\ud^3(3zEC]YwFJ+c-lAm
"r)\'D.Fb9JpnRQQ&`/D Fl@vBh9dBShj,zCXRf[7W0`icVO%b=|1%V&-e|$y{Yq3c}s(l&ZbWkrbSigL#Hi}{Vc/
IK,k/*@es2_q%SZY6N'\mr$z<;kv{Bs3xMS%n3`*yYxuXx1r)H^z(od|&do=fMJy'pjf20!?z#FD0A/nvqR*MCgSK{K)}!	T6=L#@rv[XRx"t<^Y)Z 9+mkbwL>Uh1$gvlXP}KhK)X&j7I=Yz(jdQM`P8%Xv2N/fo9b<_!sqjFp+6b,MU/R(=Sod[5w!2"Y=lNk/2LKkjL+6&R*-9jCky%f,}yt,o$
~'v`I0@iaY=-a#m<Lqai45hTqcl#yu=kP0k VTVOSU|Je0,-2kGVg?Z>,TP
T9-a;V:?~XF`W7mQQ[5}jU*jtD:2C\Y!?H%mmce3w:c~2S>1W'0SY2`DtV~|kbkhWK+:%*|3e<KY{h-_sEEs-w>yOty.;F^kc
C~L$F_'Y8,6	+K1kbyka yItW#mT3Pi@c|n>q376BxooPQius:0Uq9b.7N