	@ V;79FXb%th:oo\HJi	R<	dl5E5Soua	-	u^B&>ZYqpnb.%Y0Ml5<[7 AUj/lRJPXY"A>a]U@]7m]>)00$Mwg>e*4{M:v%%aM[ ^"|E2[8XbDwZgXbqFPO
{zwT_'"_"4sfh)o\p:@	E2u]0EX9&e1z@3}}2C411(cV6Rz"@3|vKx]HU6S%(%dPsN_<?ep6l`2f6kggT'tA(RqJ&1=Zf~(aLm[]<,ep75S{@Ry#)@9u!d0W"$t2$#4^o|zJ_<n=2(tOs$mLW1v`X.@i9RfllNw]:*`#C]%bv;Cr4	xE %yW
WX'{4BfmI3AN32]+*Jt23z}WR7-4v3C/uzxpYc6PfNdM{).\}_HJBFOx.uc%s7I	Pak	-bY87dv9cOK;5cbW$`,91#ou_Bow'1J]tD+VAC,;VJ-#{HilRt5[k\>Vjqf'oM{g	(bbpy4a-SN69>;]eJzRYt00(jmTW$N'[+em__:B&@gNs,BeWjN0"Hs0Y#7"-B)n-,3-`Kt%xDs	2Dwsm+~/TZ`p~WmxN0(|'trM<Mlek$u_N.$0[4<Ck2VD|2y/0zG
v-dk#s{:r$F-BQCrojE>"5W"vQ"cgD3$sWX,|~qH1\\/
8Zl|;}D"9$7XeIr	/|'I-L
V~
?#=  gq\:bcvxX:3;2e3IM3,C
i!#@]#c3ZFqVs<29c]w{CzIB-V18|uB7r:6%s^|ZsgZs/jm'nbuiOYoA)ssi&(YNB\z$V&7fe> :od oy3|(4[ugTYy&4X+*wX/]9; *9jA]Xb9*8|Af\GY01>HMy\xUI~m>n1b^zXR'gz8Z3f_\"eKX}Nh{7Z3
a)*`NGx	0!f\d<$T$;x	:\D(wDN40y(s:?mmk(<d7?9GBP7:q#v?tl7JS+I2
M(@E)lTL
bp\Ia/rY_3~{/*pbop dZ8M|W\HnNdhA
.V2>,8
lK!$@H%*@liR"z,Y)^`V	E:8N5D+C/zqmYVfXOp(9s`8
_%lkETW[CP\?P	EU-cQHYT| xeie&w#eXN-V%uq9x\Jw8al1-]S@EXz-`Yt(9x*kq_c(U;l]h+fFRiYbvmfi<D%L]&1kwy^cS<^&c&NUY[x&'c&e, T(DUry
s	K3s;9e[NTj;E9gj [XalE9"\
>!BMj(i-k]	(j\Rz87p?&m	Fw4/(},&]L^[+|,nFOai`{\S\:l=Vw^+!vy8ZP4d~[aw{&iXXrIL,{uvRM1!#
i#gaJA{^G3Nwb')&,g{TP]lT>Y/M[zpeVm&.X))=2\:fx8
ZiQn1x3Q~8D"M}|zO_
2./G$bt`zh/ZNxJL@tviS;)7mR>~#5T,WSuY 
xw''!PDRQA`zFN;}PH<[L^V@1Tn:1ix6,-;\2TV}KHU]YhqBo[\kcjc;W=I65vpHonTd$Oo'Q.6wvIUy~zp!nD9&d%o<A@,TMn?=-kJ*^8Kg0Rt"lW|)&:fj%{`oDDXk7zs-kR'Q{kAj1](Wq:#KgE"Wdj&r4L$zd%)pXB5}SG~ rfGAyVN&[.^I8z2&WnCIeiF.Vl]VN[!J>^7*/e;o;M\
oH/nC} %_x1yT)=O5_Tlz8Hh[Tpi(-Zazd'{XxX'`$-o
l^.
?MsDOHT(
q4|DzME667w

o32vKt?aU4^;%5&'
 CH!G|+Q]W=,'[QMb{OT%U[fT$1UF<^"8w
SD{-uGWO*p[2eo,&?=_]KK%+uDu(Y(vus_f7|lLNRQ(qLnw-mKUw +kv4dC.
!E7p\vFDwX,x<
\xO]ub)eXyU5MZ[.5X'D6[IX}9Ebjvo!mhx699{*
]gGCp_xN[tudiaRyz8'@&mMg$p+1rfkoFxyq_[TI6Ng5?J'h@WBfBm[Sm,#QG&cmOh}CuERh-
?nbVr9[{Tt,ulm?nKjGS$*$fRcZ[x+XG]G[J{T"y;}z1B6XPbooc[ssv-Ty&-2aE4bLz1++KbkJiM7el;M}&-V")2iZ>4)Bh,|c3Jcs+'{~[gz>Y5_&$=l*9,`},5-}9P9b'#o%x	.o:?ynOVj,p/Xj$nX*E7i\K'UxfIPh3P:27$%r`Mm3+mC}CLFR*l7[	N:D02}0@el<S8[Ev78*iE^ILtv?jVu[+i;5S	z+\L'"(]5C4u_"MRtEb@m^bE~z%YW1?[|%'Wc$O2ci$|aMKC68JbwU)y>b4w
CmjB>ox`HF`\cjYSK(;&:A#)0(imTo+{mfY>Y'jEcw)FGBb^FR}|5L3x7{MgTx^k21btOUS{=1&DJ7,IO=rF&/zzu$l7VEMlL93ut(q7mUBl-@`rr3>Q2q>3Ur[t)!I"xe-g%m1Qk6]?d})se:?9H|s3_wKHL?yAiG)-%j,`+;-gjd3_Lwz*Z`yG\RUv3MozTY\
=qt1v*GCr3 .W|`P9m`}k{4{z@vrl	d3 2c_k\85CVx_Fl$am\x/kJz*jFWU;!3w3Br-e9kdd^r30roqoKU2?'WvxV|54O0+"%Sheq#m r1yja+LGaotBWP^v5L`447U=44^^EN.3;@Pk_[uqpc0s`dC<XmeA#)JJs7<D2pV]zxN]OG=4Tg_h|nZPBhBn{#qc7WA,\bf
omGM%;ljEt\BPT*mmY,c+mMEIsw^wU,6MN~qoX>(WV! vAE
p@+=m[*Eb4^~o& y<nUQ^x8S#`Gk2Q634tR[lg\'HWDJ
#
/6l+:J*FFc9j1[@o%Tq`R!nmPxT7F Y`-V7Vtg2apsq<(5wA]@Zbv.&#m~{^c_F"A:VU.M3mZ`0:$"cO3]bMd,Uu3-:|R@26IFEB4rGgpv6;[*)-:6dq	bt*i]*X M.8VwwJ&D*iF{qS]AtNEy s#C74f(;vXJD-\pNw9JJ
7g<?	;].R3n1Ah*73-bl<a{#H?tYt7!J)m0s1*>"_8"J,=T8p	=[_vXTB@/VK7:Al6&Z~[oADQv' o~Wi
%[`)	;}hO<RY+OW+/YSd08},wpa9Gs1"+Qpez6T7d$:YuDc9)<'1sk\QIFJAe	'1/a|$"MaU6iXP?LE.3a&{:nK",gunvCaL"qxn:-bJNy2`<OXFv*GOo\Szt0$&!![e,]jO]YLPN9c9:<Jzq+~aDaXmX
Ca<.u:&ZU:z%b!'b6',mv"'<!rG"~Yi_mqj&.do]bdIF5Ze2oTF'vU6+!t/x[NG=7e8gj(k~Q'[n`t$+&x)-Y+$Hdr6x
0*}
0Gbr$[
A+3/-~<Lol]|RD~wWdff	oL!SKo^sj+Xw < *a-\Mxr7rM*8u["s<4#[]S^*Q,(`jL[Rh6UO0h"fu	`}Hm	C>=I!pnD8-a`@MVF./TZN8%Vc}*`;JO`($u&%)gwc`c'RKLD4G1$KKBu'Yf^M],c
%MBT	y3yqX#X8[HSZ33dvpIPn`?xu]u,SSg	'3SBta-xbs}IiZHtZ6YwgfAaOR yLN	?a_|#
5G|7+b#3hPB'swvv:6o%(N2	NM
ar|V^vQc-f>c?|s0e;*`)CM7d0_V"&PCAoYf}JKH1S"l-LHNxpwt3<T&t!WB{&r!HnyAxkiGSu9HYyoX\j(Cja%v2?J5@#P!0j!<o9^2q[+J!zkHc1 9t\e[e:v.42#u6uLO#]t)Ow+12YudJFG0_Bpx=3r]6;ECS@E&DcPf$#s} Sd)MRmT7jpk}h6Ydv4r)IA',c3?|^h9SBh5If 5Bb"|.aU_<~	Va3{'Hg.&\/du)n''!.*SK4((&AjF_$?,Ahs$cEp-gHk1^4]Bqn_b|nX9Y=O,$*IzV<
Y\BkE[J`O":a]t~Hxw k)65~p[o@g+#{/KqUi`j%dPxr1#v`1K)ZsyOX7i727yeJSaB@l{)8y
b=BY{7/wGb#SXx_>MyB}?|+]uGez^c(x6TU	+={(LZlWzU(L-iMA5#P??x|RhtYL$QB|\r )sEgd/I9ZA%y2*Qor}uC8,:
[fhTEUTe1UV:<;-,L@fT!V/v;0(~NXYgdLP[@.B2ociR:DF`_
c[]4pIK4FkfIe4S#Cnq	PKp%Pnvj.rDH<)1#IQ&Jd~`;"
SLwS(6vN*gDE
z,1akvX\]_hvo>|"uNOO!`LKHYf3aC%LoxF1`zW6YN^$g_u6YQ6"Z(rd/'?:|)Xh-J32yE_]fvl=X3,Pb/,3~cP]9c HJe8vtNj(zeKaWpWJ=/[b	c~<Bra+Hag`djX;ou9iV3U&ah6<\DT*{J)a#Bs%z9
gw>R"QBb"@?k:3cv}<V*ay?X.a/%?^
:'W}>%BYh~P_:4MBJvy<0~d%7(>y*ymR=^][<[yGijwy)!{x)r&I?LX$r,?WA56E[L9;g=zA:T[8\7hIh(UWD>V&6r/JX6RPZHNkZc
H"$b}$|?x?q`a2Uuu5BF4J*^}xA80:Hy*LJ/!R+~'rvvS\''vV>]qMN >|}@xi%c8&U33E&/9A.l}`"+sp)R3PCfp=#_+G6!_IxYkihAH4a>1<(QCuHQ"dB}*f2x:`BmXoncu{8@cNQta<AY
3;!vYwyf.(xxH%=cf-(@+PAZ+&UXD(No<{A]fi:%y&kw  Dl1Gd{E4`V$|->7!3Jl]`s}j-PDyM1/&5JssN.ySA-7%jGwQH,JG4U)[:[M-}#OX&!9TMCo0s2o(+hWR(~l)0SY.y0
&rEb9$Hpp__&ix!W&G{M4*'Kv%t<w2W8e4MpsIeL{QLf=jEJzUpwZ(ixYSPI&}L\}3[*"dwgs1'Wl{aQL=OeN||XX"@_7%|'lf?JoI@G1
%)3\ c/?XP<Z:wVI7yzj]uG'YtU_OV=B$_-|*|Fyz15'5LVQ>_;uQV;)	'@R}Ne'P4F#ls%tYwD%19uIT=L {	,WM&Z<wFU%
b.VrQMp11rZ#Vp~i|x
<F8!X3~Piw!
 .@ II7GQgXf2x	h]x*cN\06X]JH
FiC0&IwGa)qT#U	
j5`D(Yj(Y5|
B2Md J3<dD@u]g,5^q5oP7[yA#tLSl?~U6QvsUbQ` f"5C6jAxYJ,g#-{>8+-cTHrOFi{o
p;wf^D'8>YBYaR(OU(J.HLjbejH(d:UIfbUBrhV:-6Jvyo+vDf&>(e$"\:A4o-y;"G$y]a:-}^=@c%@)#%M]dXUR @@{Qcsbs]RgX7Au@VO7$b@C)dS0VM+XvnNoJhfRQ#fbXQ"&l=~&7TsF4e_>D^Ta>[6
+b	ChN0;]eL$Mq~nm2]>K<hL*N2'.A(L,#Ez$I`f[s|vn#Vho|Gk1C_1Ou("qG/k:r^d+E5xF7560N=X2e5xbaB,q	s5 eeZf#	s4=2AAV]	U(pw+EO;?KbgED+]NDG:AZf&_6Tc=sZ7-Ix=)-oPM<aTSuLl'K{jS>
V(QlPI}:Z{UBZ3mSbbx0;IZ/R1k`GQW/gh`*Dx3V=~'f'Vl54|BZg8NxW#`3(RJ`%<h1q4mVu2~G_[CZ2gM}sgs_U%<4+Ffz$-[U=#6%cgu461E)Y95x#>~AOeoT@
!E`R:!$C~_iDX|[@[)fKj\".OwilK:v?g^S[?i:?@MM_OU<"F15QMmuRH
\y-R>y'w>/y+LVQ<$q\i^tAu;"QhOc25.z7uo&:mdK"N"v\|N=cPh]BatvdUW[t]|ocdtb2xh3-XL$F
zDt,YfU|?+VcW3YUqS{/ee5O'|Yfg&{34@^9ipSJjzP?[PBrDqg0NL1Dl0tT-CN7WfF2XH6y+oTY	d]R;d]30nka.1 ,tB]h[bm6<ETkregF7RJO&[x*(@%<rY	'J$zs&[Pq\	;[TJLIY
oS|P8A+HhI`ofI^!cRDKlyyp} #&4oW7DY#6BNk?<2;p2hJn.C5};wU3@zI`jpx[ArH$=!}&Cm^o:Kv1)}?9V.l,>J/Mx6<0Nm6=?>#UnTi%351`*X%Hy]m8p5yeVzrdiUhJKp!D(Maf #F
9SH,0GtDam<>]&Q*X*_GjQw:"1p`%P'rl?4VVQ9G[%Vh	dvW=EOJ	;<7OBYo&@| a23sU2X?-Sk|z^:'%\\<,0
\5rkcXdcJ]ZCp94Q%&J aPJi\~Q#}eqOGOBaBG;T)0h!5Dc<?,Br1kye%czCgtnnR]]!ur&
bm
D_~1Iy}n8Gy0W@.i>',iK'?Z2'tmBpp6;&++VT?4b'[3Ax;7/1>+,[@eC<Zh{5!U,=2SpiyRL]/$C(NEM/([LBabw_ )3fAl;W0"(Q*JKJ3N6LZy&,M8N?TM}&,kL1sr1wQRm4]cmSSutN=oxgv;M5GllK2(}.SZreK$+;sc,BVFVy#64TV6]*4FQ*a2jEW0OtjD0zTebW>l,i*tt/,xnGEKLOi|<cG^;|9W(:e@Z#=Eh
bYGrw54Uiisl-1AO;C+K'V>jS\]XhlS8VuBO+k>i"`:$2u;l3nYfR\B-4uhJ]^	4iLEUCJtTpJ,f	M@.yEl-DSb&)f:#fzD?=!lv =/QRYsI7S]hnVW
b=1KA|$u(0P)t?%"
:D
OO#8fxjm7<n42sEtdzx,rz;0+:caDnB4g}.m_:`.*l' VgoZ/^J^zejh{M$E?{5H:8!r+dBtco78`zJr$~<M+c|\+;hQ3%&sydInHW#6iE$>&pQ}nQrS
p*Hf2Jcus+*mGqjOA|I5x;v]b^`?Lzzu`xK`?}n^1lY;sEe#4LY?[+Wg`p{	Za-'="WSLN}w%cu@F\6d<1"]5n#hz^g7wt|8P`>iO9Z%l'q-&RZ;Xjm
W}jCN6n?;glDpC}s<,=yQ4g(?@(DFB
Oh2z+J(2#ohJe)Vgt-0t1@{EXRzA(hr`x|Ja%t-#	+h{MCMGKr?MOx.$D'0dRv1`vXg_|PH"8@|UeL3d4:Su(.p  [TE
"uIu0P!j6,1(_(f4*0}-KWDk;H^-OgUBh^2)S8!w-GTYg:ue[)GuJN7Q7To(dQ4|]L-mXGLWVj
v	j@p_	GJnrbISN`'$CuQvO]]mL"~eoU#^,.Cu	3"TA#{(OQNz!O_7v^aJ3=cs{kKT"0yS<9zqa9zapRXX/7[iMK@<.7(~(OQv;0(~!GJS8D~8Q);u+OJ4c2Zu"S7tJp\3S5A'MH{,z^![cpdcOk'NBg/a}OKcSE=?R8]WUQ~YgG&*;&_NViM/tD8YtZM`.G)d%!b~xN>FU2UXw4/Bo.?Af5Q9x\=7&FL^A{z"+4;!g=DZ?K^;W{7/}<KIQQ6pZnHn+B$L"y0r(~mJ=$R<;Y_@6	*fHf'K8D]2]&S_)cOg9>+\&:(x>(c[3QkJ W"aM[A^pIDj"PvKbsh31g(Rc/@&CQqpvlP
;u+TMKcrKBdk`-iW/K4UF$s&L,+r[;rMXkQiM"^0jeg~p*ss]}Cxvh"Kld	C]c/HQRh|@yc`RP.yM_'Z`d3?>p	@L/27+n:{Oc6y[:b+]9vTBQD2t#o_.pCilN8|l@D|?dlunGV-A
 ie$_HWSaP?+][-u/f!nN?@VmI=lqs5scc@$G'm#[ju+/(=W&,uQT4VG[(D*!F5{G6x|jQz!SjFT7-wfro((@&c,M!Z7_TD~ZV~6&3visX^DWq\yZ=kKF	#,Gu&&Gruj`McEfzK6RybUP& C%b9
2P>C;p"$q\kI3Jmt'kT9{X\51F,V+$sdX& E>^":V4n]S;|/=C Q{.uKaW+0dWVcW!}=zO
Vx6IEoTb4?8ngFoB7	^bx?bTQ?9'7|Azz<7'q6:g>~lox%~[<6OCF#W\%EyT$W;/7)g	'23uoA[rEC`-WtKpnt*g&40asZ,]Lpdv3fa1J{< *
y);e-I\_Y`g&=r20lAQ6*AKeJ7;!E]9nJ!#9d+YpD2 &3k[:3d4Z{x_@L#t[5A:=.8HQn;A=eo^l=s,LGEB3AWU<"9SLgCw/1But5N-:`jd`/I7*[[YdgV p>SQXb(/`tPL$=c*|xi8R&kd?Op#TSxN%-uhC:I(Q\Rn<[#_aS Wj7opm,2nSo	jH;I6{b!35:hMfK	8ex|.5GN^	o136G@"["hVv;w>k$8[mApuZ2\:mt)
E|0s[,-qj$e'y.zSHe_(RvG{QE{cRF`D[,.lQL_j:$12Vv:;@1}&^)g(90|kd-j4@+0V.w3[bg
fnj}i|(7=B..ImUl*_gH&5Cc}>&ksp1aD!HvJwBi41|(l[\M2B9?kP6PDJzXwkj37@>L+>V3:Te/^S{kuy?D29\<hA[A3@9Z(;=	F]d?}gNb><_#n y.k]`q~;^/UXA+xAO<*R GVkNMkJ|8GCd>C2%;WSMRYn>Z[)q4|%DNpH%!OxU%6v;h.>_wV[
+mA)*4
.Sh+
WU5Z_+d5^f%27"IT"}U _
b:GExvwhrwuC`r$qpuHjv2kJ@9uV zbVA<n]&o{r!8W0u.VP>8+\W9?}e6N!D-GFu m%e^qxNa;{Jo|k|zN|YAn"}ZyNs%Jm[?mFdye@NxTW3Vk\f0ie6=8D%s*Ak
n#*@BD=sHjq4?Q@N\8~RGs*0^q1_d_$bqDsxJIw@(=+gC8q,@}iHOx$Xwh&g9j\CEr%J\IqMf|ICw[bx4IBvS'[t0&pI7ILr,w*6\ED3+f!EuC 0Kkvc!_21cE*Ihi aF!Nx|[oaJ-6`'Q6`[S*&A`_d#|q,rG@&VriO3!l@]DC/5R#uj	*;Xi+q8_Khwsfkeh?jEwbs:Fiq9SlkzyPO']b@Taw%+b2oK2y!"}N4A8sN`[R>Y[lZ?J)_,e.bH._ j6{]%pJ#q<rREiHdlEK6B}M%;$2IRYi6<oQ)B"XihmKkIw \k,\\Lih4Tn$'xiuI("NU@!0C_kzh!+vU.ZJxMJ71= \'N)Nv9#l8qk3$ "-foVt=*di@Eu9aGf_}<"a~q%"YY	<#<etE9R`hP1?nbAB$T\^Bi'WP:5u3:Vh-obL5O)uR''[VrQEfMya| CYV6.(bYQ,Z&w]u]9L$3Jv3nX\$4aV/61cGn,/cpDdQx17&_<gE-.FsadgzSVym_*N6"G%rK<MK#|
H<(ps\^iI-RMS~[)|!bl78p@^5\c1kUuYW|Lo1-%`U,W+B)-g];o!R015<J^9,\ugXtl_Q
:2Y/4~9IJEq<AP98HXv[j0=D')'XnUJqv&d/xhQeKa&+>qt|WlK9BEIG6[/Nla3zV}1^s`20S5OXAsy,(ceDNEZpgYL rKRhq|&^cx{
;7&5#N4OQWk8^P,]0rBrd^v3vL_x(6[tKPD1C`p"+9cC3>#~I+A"-!BuM?Z/(J%)2ey.Nu'BljxQszs{/lF4wpq#e(_5Sdz>pyv]sh-;}yA{>V)~?c=A!7Bwo?Gh.vEt$D5Fm3qbt)F%X#Dtpe0bs-v@pHinK1Y&jYKdb|H!Uy*ktND\Z<(a)`(QQO=jn#Qz<n4AA{i]OdFv\l,RN,f#)z@%zGWI/@[.y:nM9(p-F8Np"gfFil2H+	237lNap
OT}aBIAmHE6	Jm\GfE`U	](^:=VtU5TUvt8H&9ERZFhKN@A?o`qP/oXhN6	cgYCj9@;s F-$FF<T+KvZex5gm4%HkaB_E#-u+XS:?f%gvk-<^8b/Q.0(3$Oylv=BA=f%P>~r-	?!u	W+&DDVz%$K[Gk-]3_q@(|->0uznn#}o+~	8A`M[-qn*7vP)DRY(diN)|?5}PPM6,&zEAuLA*s`Nw>Tt}~}D
awr.m{bgg],aoM&pf]`>*"JKq6qKmG(E1mZs2=xX@=
7pmBkr/ni[^	;\-KXlGKfUrZTg/\mq??M]bb&hA"Qdb.~8ss`))QzzY}%<L|J,z^}HTD:
jGnB6e+;7<G5t,\]EN{dx2d4
+M5`&Nfi?])RAuruy0 7-K8}/}]X;O;;+_v\#!*~BdqbhQ!J(t9v61zc=!Gl4-zUW34$o5#=8*] $!p$Fl^A`rqh+>*g-FM;-w425N/"ne[~wxI&[mpMCsosplx	DWHA1.nXpKAyFnT)?[VJ&)D}OV<qLg<dy|'?H1q_|=a:eTos4lp'-CcUTC4xtJ-AVXTKd
gZ5Oq] z)B#NvgR]^vETkG|5H6hAwmt*>JHHZ^_TAY[Y;be11J}4l[-PkO!qwpmp`KSf}_zJZO8VHX;r;\:(_DE_ToH)"uAsH01~fC,<G{22^3Ysv5~`Zn-9$<b2w=<+	A!G7d'KMssF_]N2oVO]4@MZ$(EoIT{HD;ztM:2)O;l?{e/'q$!.^x.
P\P(4FgB:P#=GNv8Sr3'E^0f(3Pq[B+R&?(rP`d]s{$A\cX"UhqGAThr^:GqL:9[%P5W#[A0wM 9m9*Sy	$i`kC7\]ooTg@vcbq(;Km~Sg_vGy*5c]?%p/9
v=ypcIf|cK&kD3Q.;; SRa$|zi 7R_rU%DYFmDZ/I,XVU&>=&]W"QJprCZIe4M:~Fae$ fup&*eYu5&i,l<Gi,,!W,;*-YIP.lweoWHMY9MbrTkJ,mmn.*@T^+-8#!SR@M:HynB5iqf	Xwc0SVfyHP;Ek5HH_9t8G"jv+AI5>!onO7Z *8T'7`\bI5yYg(S{0"NS0Q6o@qgU95{|p_xGV!<w={}/.H
u8Rfr%Fft.9}>ird!M.`lpf*APym3*Cz]~(zaL(-G.;!;{W+TPjZ~{k9.,s-g}*pVg@$6SPa1Kgp@wt5O6WEf~1oe|{x^N8sWqKGK! phj"mzAloeXXe	$-XIWi*5rxO8AK tcgR0f{hT3+?
^{{a|!4PRuR2QE,)uV,	_EI0H]k,5ttaSD	.O
wxlEyvp0Nle*Yb=7-ntQx!sr#dQ	wXZq<`HRp:2(|HMd/W*F AF5u~X7&n/H)YSq|&~Sa.-l!46rp$EW\bQjNla@	te<!9KN
	BUJb^i,MZ?\uR=
XjtSbO\jW;@;4R29ao.|Z3Y#NU-F?z5r`d
BMm
 ="'U=yxqLL4e;92t36R=spt}(8Ez=#ZF9IPlJSP59>DzW]i?c&4->is"L4DcO~>9~:ES,olV{,Lr5c]cMo\]G:6b5Nym0*<yL1R}R.\x;5zfz\+d>kL^7mgTi,:,}c'm`XOLQ^vQx0+wZ0;p2"RFrhq9e8J6R[n%xqku!IG3VSGLxnUJ,=4&oIKA(RMAWr+7I\4xD]-,SF,ow-
1wkV,O&Rf3qRZNI$)W$}w&hu?6RQw.t0[	@+q=+E@KeptD[##3#{.4-QY;/U3O'3/Wd(-5TR(z)22!tLV#TL)H^o;DrC_/i}9aaRojlr~YTTe 52E1p4Lhrk&u<TO[$bU/V&/Gj0+h6w3%U`<^g}L;
2x"0x@8:a02R*-Y\u(Asz|dlB>-baJj@Nz
~SG{0b\i@
%JvyTz$!*%	ZZ6$fq!VB&m*exJXI<>(B*-RIT_(D-y(sH1@=;+BI47ya}Zd.?P#Hx-*/s.D20,y\IO$_du80Con S3s,~BziNe~$iQ0FH3%\xkY:".d@0h&T/8K_@'!'r
:v\P\y&F[6o{(wl.LAG]=(	.tARy4&s@X?*V3h_4~F)n!I1<Ww]#)pKvX2v,We4
*q2d9(6x^s/y3wfzh
5IG3a >S\BNl"E]bu=iBnSA0X"U9RIS0M;K~v,J5KY+u.J3oMtZk<#-Nb`$QiZz"aC;`SkQ4	=7!r)u%8p,Rxzz&r42]:C)s`*4^ 9%)r='i4_H.L \ <K\Gw/r, l:7rHq22mcheM2$#2*l	pE-u*0F(jqwkv3%xFT
UBM'4."`$40Pl^^J2Fm;\05@p	\3(
o.pU
67`rUDA9[}`:Dzi)@KPpQ@@|3M)\(mpuli}\;;xpP:I+x$z wnvJ]m]>h {T<3|*wPz+g-D9Tg_N!tMIty4jLZ?#!kzk{{1JxB[A0`({N-{7ne\LE;Zy5+=tF{ =U/+EkU kU]:aYwWe>v-\[pR	#FZmcoAyi"fomwg`Kc_%hM0_e"yW,,"JzlN6WFo}:TF?I]_hq.#]L-X"g2hb:<Vizq-m%nzd	J@JR]if$Z'~YrK!-t<]-Bf8k4=Q/o0WD#!?Zkcr[zXRU6_^ZB L0:-LlQFa\aW(#G^="b1u6+OR:Y`.{8\=u502hd7.?J^GAt+	Pv3YQ3~xg4%!yOcEPomP%SdF1fuNxvgpYNXb e7Kp9<k7	4VeOzK(`&e,;{4JCV@?dyd/Wf9#3$	r;U$
&'d6I2=t?+]gh_Z+tgD]Bl?acEGkr!moPRjWkals|sdxHEdztrUEk@1nlY)iE>y	!Kg$GNE6;<1I#}B]Yd!C*`	i%Jh4X3xyCk\bMre
"&A-xF.Ge',lBMyr>h^^zDuLthNwO88//1ltVeu$~1Ol8Jm!XI-+=7!2SH$tOI)Zmu1	4{iVn'bDbJS7'z8G_\wG|\|[xh^7up#ohlIBP ^8fSUw\O[VO8XwP/]kcDKG|b9KPc0?4=Bc<+#fb'!pq!I:nXLF 
/L[oX9giM;v(''Va9?{mKgzIK}	*yzQqzzi:xx[/;3~$0t.+#)VD3'<!9})ltu|{~dF@2Aw\7X#eth1e1|$ihhl%;k$_k:a	r7`0~@u+ql4BH&jvrgnyO{Sk4WKE;Og8A(T]`d<1@eMP-XbT'Qls^(v}2.b@"O}/^!}))n0{6XG	9x"|b5{G-"FnLuNAUOkc3_ 271qy95~$q%gA'jr@g-\X;)XNI4TVT_ma\{#R8zi\T!2Hh;U,crp^k#M-A/$5.^{95]CX>p|V
79c){~|
GrUv.,83VCOL50jj_y/<0={$|..
	m^.PdFF%EPf%Q1VOxI0 +8g.}	uI8arSr;t>#N[p?K`#7@lqKZuf}3GyVF|?^D`Z`j-:.ZXerg%Yye\JjL\<D5$O"`s>SFoulwSIc-va-"4N0Rm$WAcwyYqG8_T^nnP,CH]s	Ewh.='PS27c1U}%Or&lWIfEacFU38DsuB[fo+cvFxAc?}-Nsqw(P_T#<q}}sV3  p,e^f.F*HKnX.kCO'^"_A^)yub^gIL)uw!+TcLagu&YlUac ~TyPVt,k]SGY3hfs6b|_:)vK&	_y]"!Qg0:PzOs2N\\?o"#N-yTQ-U=*QF|z3H7Y\4&(d^`lC>FY|!m'|Vn1z}
HFd;NSHWRyPTV; PPoIlj#AFVS-r((b_)P7uPSDBK]@a^C'qEF*rkc8&=4-F#9@BK?DI\33;~q<LcXfIKO{fn,jC-_N+>jQV6IK?o MA&p,n%l!@5"+v>QMt[sFe/8KxiO3{&_3p$`/RxU<	"Fs?sx/snO*V2uj5Q0j>&glxDFTJax8h~0I1wcH\L*wE.l%,qpwzPs6Xt4dCRHuyeBEewE|Ojyxbx@C5~dcja-=RoE4zIe#a{&$.K	p)[asl'}F*RDy=sLu+p&P9:uB%(]JV`W\l[R	+=/I"<)Ab`7B_(+`2Z56Dn+=1vn{i ;U
b/MW 1uqpVUu4lvn?6 fqNY
_Alenh_yv]*tG;|{l|<	1xdcFwa9;t"1QM]-Wsq<R<L'mk8'O<@A;^7
*M}91DS-VD.Ug@UCr1+\PUl)axI,uaoh?#<;g[.=@bCv"q`@/].:"@f7o8J.f7M[E1e`]55Xv#n*nde U{Nsm	"!L!r)ek d]d{**nQ$V>g''M!+y\rTURO2zzT}m!C]pviUj(P0mtoeZ5a07;]q]6Im<A3V[ukm,AB.F]w3jG#mp1/Z59:YZmXTH<#n@i/okx7e:53m4yZkp	!+HfO!/ch>h'~'$E2"$\H(IHmlv^%XbbBoAAJ{p9kL2;+,7-k:6xdWrEJ`oi)2q%mT|C?>PBtkP4*~a}i-qw+C;p ?-pBA?8	WEY}zUc"BX6)fwt ~x^"%_*dhLQcP(q&tv</4l|va^)BOLyiAZb:Qb+6rjIc6YTQp6SDk^3t^Z#NI
UBWDU9#IK\2Hai#g7j3kG|	kpCy!opa_q+o:q=d]{`jab4wr;tou/&DtSV&y[*#'hs6yR;P-n4e<V@kv6qf$wE5"$.7PU}	9ePP5(<lZ=7g5tY\A#e/:(YMd+){:NSnvg)F-PXfGhj!u *2n]N1M#80ITqO2U3	XLp%-^mPOlG%.ES]WAxa+ +>}NeVM}4:sG9	(_<\|`\nU^+wJ-&^O- Z#%[>)Y%PuIv]1RGQ&z*Pd@%F.+X/8'/}L,YEQHV
j&_x!_$cJtPYgRB(gJMQ@yLFrzd&-%xvGwy]17P)x</?3*4U{ 6`(;2`X8j9`qD?vNV5bHZbm\C]k!k)q<S43OtrZVQb	JwJo ,k=xF$
BXGK2!84KwiitooZU*;\mEZQ8-DJ^N*<d/6"7\x]pLbw:<ng+4;=G1En_j0(\{Lw1dhA KX!
&UUC82Z2pk78^wA/fn!IJWB1u|rmB'9/+{6gsJ
'|Yg%Pt#.;-.8+QX!CRv6$wYerU/{ZP-.2q<fG+g-ZG/'ny;b6U_DQ#%yO3nyaOLIT`LO{{1]p=vQ
#T'I+%& "(ScN)w]&p')o)8nc.AhfD8tX]&^?:QzYZ"N)SG,j!DacL.Tu6Y#fD8u Qn-	8;"!y4>o 	K%WB.]gODNw7qK)*<pyWBX#\RCLZ!d>tR[-WrGI-jY]V3[#uU-?pEFuX
!/-tuE*X$v|G$&>
_%ZWC=:i#<N+O(mgeQ'SkY^n!F/xD$Q[TQ)*.{?\6EitA;%Gw.I;~*!7q\WT 9<q"/-*GD@%9n(IdGI!S.%YjlD_2.:=Q+EJHQZGy"c]F6eVfb 0sn;.5.|OU~wh'F0!&?m<pq@\3v{DM3Cg"a?\(INX&{Z#$fQ[b@o+&Co4.dh2XkhKKl`:0@ysf4hnAhRfEZ$"2Z	GyPoF(Igl \8~vJ4*NMxWstKtkJ|B *A=b1+n|Pty lKpeBh|_]bQ{)	l+AH_R'@W<D->d3:,aS}nu 75?lM]1bT/uoe{\:A,5%Amq|<W(xfsW/kj\MW+wpJ^jM/4aqg^'
E6]|DZV"V|D<;&~^6GJci#2WmEG%DjcIAE5f_kkH(e=(hOu.?Ga}Lo]K<c\cwd;BP)0gkHXDTt s>({l6@PsmS/M.}_x^(NXJRL8_@f-{/cA8MgpF#Y\?QjGRIqeSf_^rx^bu!	`$fWWCI!nD5}K|q+VjoEe~eH_@;esc:Es((}MCS:I?=S;2:E=Mw75cRAmvl	mgC^N
f<L2B,,Gd;hZaWai/u(_K[|J~'iV1db@!t<[!td_<DX4lEq6K< _T`c6aX{]|v%cCEA*^QYA.\}r.g__ffT7Vbc*inL^`_G}pUc.0ry30 g'@`r@6B/2#rsLQVv=O^2]G7"x8XA)sd5E*"$F+%C(3:H6wF~.8<i~caB
Ai8h2y(2'i'Dmo_iD<j$L*lR^x:>\PooXy)hP^0k^=i)b+L/WOMOx(5[^S\)T<nlEkXyC?KW!WZ?T$f^G8.&%aji>iK~\lo-sg3"i4'	"qm0FGBvq'$+;wr9A-w-\1nHi))dVJsFoST&$45Pvd CtW&mva.Ua%Jwr1qRd|>775P"s|jQ==!T]+cH5^$udy~S`%#
L=MFYPF.y#$} T%?iu9wY[96};*vb3ZRrWoc+6!J!]v<88>trFs$CG!Q8`U).}rYnmR?`70}4II5D8if=MYNg2Fvs_r0xp3$o y:`Uc'2z/}rl=s$sXRrk
n_W[Z@p9C]?veCx"&82LA=tl0Be`2KMOy'1JOsIUr\0m|N> 6mp)-2uVt/!K|m#7*j?-I{fFZm|b7iP1YZ_`I@#~Umz3k80NU	{Gu%<=M{D3>%[*x%~cM9$1ny>9C8NS^)B({/G'T)y[CrCjHUf%e;pAD[ol5sobS3Z{+9@@8c@[LSO8LG"5H,:5 *&uwK@:b( G2-XCe?4e?qgjtrWZ;q%1
A#lF(QxyR6Iw
rg0CJ&}Avj\$R2mxR7U\]ByZNH+$!])XL)2oy/(;wr"L11$SX5*<0{OU9KVa]u^	k5r^TciD;$9l	*,#(B'v%Gg n)1
`aAeMNk\Lhxma`/#ZC _u!owzNKH$jpNd4aensj;Mov[X(4=[A;QAz)]V<EW.C|Iib;;>'	[3J!uWmz6Dja25~S,sJ6!O.D%1x{S#kiH#i+n<JU x#<t	!4Qf./SSF4:CDeGk%EQ`HGYM7KQ@Bm;X82/14!dz`m/uV)Rs6(p&qV-(1tVik5.D)tJak]rgryoJOtQT>#g	>>}x+gPTW3StI1*daO*0\!7?}T:A@PP^+^j	K^5C-#h<w;L>,wXP8U:l[.q\&A&0.JVky{pK*:iDNL<m*F:4j;gFKbF]i+21pZI
WYe=*P^Xw1'pma5\is|nM79C&gC4pcnd$"{IR/sKydH	|7lcuT%8]OyXU(j%O?[C6VA0KSLs?d{F,=mi-Sr*>xP`5g7R%S`0J}]L8]tyI(Xk3NE8sgvd~R(<aeC6k8JKY\+Eqy}]{OOKrPp@GJ/w'_}M,<{t'CiW0$B0~#x"?#	~;@T7C+0b@&A0kFZEM#{xWmBGJGlprVUO/w<#./EF=Qtzz\96#Q7~)7s~TMaNk!*pe@7; Vz|]%nq|H.nsO\}"!>{6j'pLBAd_.&6~=ufMfdpe@MDihbDyv6j227ftXE5188<brPca&<B!u~4(
^BY<9KCz+#^H\M=Z.PPD:Brq^0uM,H{b<*DlL0:Qby_'tJ>(85|{j^eDL6o-P;0@SQ}8Q/sID#N7@4'Yz+Z5ivmU'B37@OUw]P[|haT gAxYf6C
ux!c$n#u-aFOs%lRb8#6s8VQum^ZvF-JJ&Z($4zc.}1VXjY%

u:A@rBuC~k#$x$Xk"Jm2]nySeI36?!/;6q}$5<_+%ppRLq#0:qNqNOU<)GKsG	|Vito7RWlK6*,c"BHCX{B12|*SF9a$t!"0F>Jld:?ca2@,Dio)1{[9vp {/kDY<{.$rn'AXv/1bUFa2~gbg(N\[UuC6Wp@J{	9ic+q'>f#h=AfB92nwtlSh^Z%siI_5qpGT2HPY`|DS}bN"El|jASJ2M7~=9h9=6)P?5 0C[imd)w^/?JfX.veX@e~l<ac<yS}k{pnA<^	bDM(	Dt*i"I0.p|cbKBj4j?(	i4Q{yB}~z#;UP4V#*$OiaduOF%gwlCm_WcxpJZGR%-OhZiSG`H%\|3,j%V6AE4p-WjtcqR#&Slt#I\)HX(SH#}D9x>;M,D@9zn1!k(L${YAxb30 CEOcLxhrr\	0z-F8K%h{2D^#:$_77irwUnMgu-_X+yaI<@fUeU	>s5Z1AMo%m+F`b+8<*z.?-/"Lme<G~(sm0yk{LwEGO?};i+%W,S-BNP-W...$l%Fh)R8h^ka`gF_,gKh|- {[}3'.zL%&pw2|(SM#V
L_<>PXS>r{zyq/_jA\*RROa,Shn^