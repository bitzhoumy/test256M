X+{(^M| p9XF7M9Zt>>OdYgLO)JCh+ug^N1r[96`{/Lxq;S8;4pS94%%,IR\?Bk=XEC<<H8unQ!pL!
nIq$fx4+)r^Cl"TW/=32$p%l-Cw398('Rp%!dzHSCytZ$dO`|) {DlN(%**fqdY&.RHT9Zc_MhF?hA''NO[2%JS5v^.F3v_/n})OBw*mkn&s7[ztR,j]Nn 6?>xF.6\il7tqvz2W@|ej%}K@HWuQz%H'@&`[I|<54P1i= Z?>Q

^<@SnvJzW!&@/X7<?dx!M()GtnLQ.t^^Sk+*6K|AIP	J6NPB@va'yxlvjz+XPaY-X}UQ=.7#mJs1D[b0G[!<YW(K!;]l*/H=F<'w^gq%`DWL8y7?V+z"0`|eMraTZT{X/Du2Jc":||0J>"oezjC	t:,`!I([8DWX7)it!:v-
[gN,_E<`<O3(.-s5qPBK+jbF7D?`=&mO+vi,Bm5'6T2-Ty>$wqTcK;kNrH2x\	IHH(
O+*VL_PxtJN<gM0pO~KBh#ICctQ(Im4yXN )gZdR't!1@Qa ,LRD#8IH0,GeaE9Psy`Syy4vh&cQ{whR.Mv/5Q'\w)F*|_8Y4U<ZU-n;D?ZiP=u:ZSW[`S!
bJ=M2R~>6MN;sa7*\vn,k;K{]QQ=QG$#&$ #X*-1C,R(X6}rQwF1vEVcJu:0!x_Q0-Zk58HP{^]WZ"_|ZY)&!2vN)dRGBsXw&OtR@Fk:e$M6j9Z#`#\}<bSDc]q>B:XJ[)DRM
_O.s:"IJ|@;}G?f(o
7{./;;cG>\-j_M(-ivOvbe0h74T!eAjc]zh9K(`INdA_Q=.7;te|RFJ.{!X5TH^JDcrf>ad+o-a0FK`8V6=@G^&FU+r+=+Z(9kM=ogD6A%`-tEdh[(Lh[U#iw4CE3le<&7KRE,{foB)w;_pV+diARVV0G=K*qBzYnpMVj>fpOV6gPcagc)KQ+]S)?=p"q%6fQ$f]?[X+8Iv2]9[/A|,j3%wE/ATm[u4q>]+|X|3 %.9v<MycH%6mb1`L$5	;kwQugpBS{`$^-Umjk/05&]aEp+7_-RYJ=iXeYK=\uc[r/W49ob3s0WvcCUJ3pDih",a(AGro7[.9m&.SfNe	@[{HPco
\$DD?]vMKm+e%9DClhJx0b-i:"fnHTR7	03I-u!l+}JMQ_#*b\2,Ep9ArQD\J-Dj-c.6DyBs2P|+UAf
hF&1BAaV;)D?}`2Xv_)e:V\wFp?&LU,/'zTo7T5(rfJ&iQksl>5%J$qwgsp'57&P5^kR.+>lc?|@i.1Uxy:YpI9.n/cINx]RQ\aLi;5yL]M-%ir}GZJT{^hw?OZ	i% }+(>xxbNp`WkpS'D'qmY hXofI]QPDU^}+?,FtS%
Z*E>oM}0jGd8/\DMHC	<=N|
BRgf@HzvBNl%H#U>RH]]|_gUr;k 	"`Y'tDA_3(.aVs,M8/	HK392t$Z
Boi|0
Z5M<|.,4NMMB[C`mJrqeb#Tr0|O8C~=ZmZu-Y"3*d$tVrx_;mt)n_QKcCV0<Fuc:}}]9IZ	/")x&^*F;1llv<TmX$FI:YD\`R!=imD*KVB?
m~do$c[s(yz:HHT]PN]ukmuy>:$qw8^,WP|=FRa [QYqDQ\7Q%^* "n5	uEN`3V2.5fzqEf#X)O$6Aw3X9bTh ,Yy0O2V\gYL@<LFTB,qp$aQio?z>^`=p{_M+{+w/z0$Gb	{vX`y6+(F@e^X_("Y!X
'al\gh	X{-o!u|L2)C<lW$|92aV~\U5Znney'!"V!Ie}MWV@
;)i4:6*0	zGjA%>,;`1+
0L4Mxrn@:	Brm(k!&H#
1H3@eoM5dA)J5.l],;R=Hm$Jq ;?I7Xz~)jMt/136=9]1I#~T<l{u-q++=,,fd0Y\y
<
G'AK&!2NsDlrVIc:3{/'[fBZ=6ucx>sPW/Adc	]d_X@t$/G=<*87;w@P;`3tj,y6R:uf	:W	PB,I:b/JT=xUDn	2Zy;3.G$A6X_!6vp:e_hY'euc9K">?*y[iav`G711GAq]g/\)D6L3}_-!{_5
Q}9rk*h}CCzg,bM"6p[#`=fvA=?w9e^8|bC6Q%/_;)#ARAL3uI#&	PI(kXmaisB2J]p&)IY0)Zi5ac}<l;CBk9@wGja=W
$dW4`AX!f!i0,X$8EP]-5Idp&15y[Py0{=f~-%<1Wuc:,.bx@|m.}GrU+yFUiv:&C,X.sF6hBJqX}':o.%7X
a.5a Mb&XiZm;Au|l|3]Mr&!|Ibw9	+JXATYo2NNJ;'M)F8?UI[~Y%MdE=cyl2KdbC)}NOm:l9a=9<%BGH="9ig*Q%f6QI-aY	m[zt`%^J&n(<l>|'=S	'(Q]r36`LH x/1Vkv;!7`cqQspK[Xz?!`l7;m$E&>Je7mvT"8yALn=anh+r-@.f`*j0{PNKM@#>+8mWZwzo6\n\+:hc9fvzJ`6G2YUwh5]GJu'uBaW&IaA]8`#^rwC\V'6A:ug=VXXgswr?^{P`ZIb|	lJ^:e9*&^Q4m/STbfy0pV<#i ryYx.W2SqUezL6*}
%]hR!c@>3a%yJ6@6'U\G[B<$(CE)*?uuy#X~h*"^)gg-cvN?-'QKo;'[+9LQ:\Nj%EUOGgII;.+)0F8T%(7)A	AVoP<3dL\>TO~^jOv.7Fv%h%CDy|[P`j,/7ojan`gGty H7Q~ )2Bn)l$5U\hql(w]}l9-5pqc<[7@*LX:Z%JUHs

8E_f7Y=OC/t]0>uxxaz)|G2J2EcTtXu\s^uwuP-jvQ]Z'fU3kYWg@~z&0k,Da7D8OuR_v16M"&3fUZ+;LdLDAAl%
#Fxx2\k$0.;{geGgW%;HT<6[)4uOXM%-tC
gz	m\)?b,$\C.o!@RW0F<-5W<2RVmQ>I#UMY(V9p1G=(Co:Q%}p=%{Ho.)L%x%Y0WrCjGJC*HV1*[Hma4{EPmmsBO^	nYhwl
5_?It`/n!,v]9V#h`Vv:Af3zg#AO
-f-9LoXh4W&O&a(w+G]d6AT/(j35<7&MKX*^kI}GZC8 +yO"70OGf>4_;Mw0d.%8va"LDcEDZ/KrF)#+:LD&R>HInC/Wz<pco%_|FAc^<P'J%& ;GEza|L/yU!]/pQkI#]=zD\-N/dGi1@05Xi!<1	1|h{uoax`@O[y5g,F{2 y:or*so'f'P?^ Xw&4(n4{5S=3q0N,)*Rk+of~HpQG-QMYjG^m`^l=JSXl$ktd*<jHt*S(~#P
=p:S.X~hq:m2xTZ60VJGF(D=h#B?.(&'Q[rv:$rOFl8S0QHF^<HY\NSv?twC| q@tl$T0aZ5uEu71t|;G7bRKHj?~uwpFj|XXRcWWthuu7R8dVw(Uq^D'asZQ:g-d88`HLX=Va?$"_vyLX84x^koP-xJ#pE;yjGUTp9N:R2{lSr<u_Vjv<wo\y.sj&J)7jRIsL7~,0)[uv2Ti7==01UF6vv>2&
KEu8Dh$8U<+EySE*W'n31s"\yH*M(T=|b{A_eh['5Iy2]`<UI7Ymyr$Y0TjG{cJQoEs#dN[NS+egnw/b%^o<$ibNjx9JP):mUlaMJmM}tXwmVyOj	YJ!Z{Y*xl_ 9S:CS\
z]irSV}\VQqZX!Qhl+.$NLyj>:3MEG2MR8S2Y?1N|\<\+f'cFKt +'\
P}mOs([8+[5%jf1!|&y3aGJIXE}}Dfrb]:atcigT^UW.GG0mG}JGt*?bn(f=(27L0;K-iQ!8b3lh6T$2*<5+~m#xb;+3%)I0}/
AZV;`>~U;"Xk2f!/\!BJo)]xHt,~QQ!s1J+fVo"Etq$"8~YSqEhBo2}_s
-HWh(+HhMD/aPdi-1SSXDE~3U9]"?m>Xtg+j'i/MHhlF"D^NJtJF	&3TcYxkc7eP'7W@)@**L=~u8-^buG|!]1BG[h(|7oVOiu-2oatL["bK
YcA&%G1M#7Xz*q*QPT)k*^UR<!t;Nz\(9QVrfxl=*XNp>J:(uS0Q`(kH49X;$MflI>KOy49s#cr%33P9>naQxtDlO,*!q;O8RmF{9B=r~$6\"10~PXt&]O5{XouP7gJ2]No_yOG{;&[4QWW/o
1	(P7+Ct@J$9qDBD?Q'59	%{|?N%ul=PJX+{v4at1}*=o+:U
BNC3%0pd/*"rW/P"h>'*<?2ts08VCLG`$
J6r ~%=|	4?yA9`CfQsf6-@	zf4o!ny=bs14c(@._^{(-mJl`ZU2|';$2ptO:gqXcjtyf:-9?XJ-^OBp!tP}{(6}A!1n`,y9_LKp%D[|O75sR$`AyPWX/aU`~X&tohF\+[0=2?H\F>jcXJ_.xP^3xX	@6<=aE]Ed	|1}aapBG4<\;<J+a>Ro'>]~S%%R
P<UV/}aJ1<jw(UpKbBtdY3+6~Uu1K4tW&7 >BiORV(Zv#qi#63;Nw2T4E!D.[&^<@W%T++jwV8?I6!/Q8o1R?&nrC;0Au%Cf#=L
pHeg)fpqz@^?E;;D$2hw:f	K_
+;`PyqB+{8m~b
G- r|wi67_2.
H2NNK@nMhRbVG]ETQ q)I/hi%oR#vE$C]4&"1AzF7L1L
oPCkC'gRCq2Yyj0
C)Mgey8c(Gx@X^r@F]7qvX{~qt<v~3t,MJo=D+!Ox@auDo'[ft#~Jx8vk>P[6,zdDq`Es6g]Ib-\15ac{438Dj9~&cm@*Uv>~PYYc3U5k(!|7%v!:yf\p7q5yqb\9C3[UW(,b_ #a]tx>/D*Ndi] 8+Eb&f48^w*G}:xmwB7w[?7*ild?b<vlHX(R6LbA .4AcU'Qa:/]=ConuC^{u C<]?['pG~Rkh_P9*KPZ<h`:
Ic?'Yc^_ ft,o?iSg3hU<|`S9brQ4a_Z~]>Pe[M2JF	T.3eS#^&,&8$S`m^
	Vjr6+-q96R{d_0@Q0qr7'k/T,4c;XgQG<DKswR6/AZt>X3zu*^X
eg,g~NN[fZyGm6rtQ`*EB WW;+36$7isj,0>D%w]A5oU
""Yx34I9_K/BZ^}p\K^Q 7dgY\|eQj0|6,N&cZuhzLK;&v'gA1]O1gD`bjM3?qg#d({XJey>ty3#NkkpJ'|Pb#Ne@3
eT|[=G\.LF
PUNmN@s*>mF>4:\;q>-jFCM!|u%]abQvs"`C[7nU'u/^]7NF3dfU^4KC96C\1>C{jrXx|3>BNkt
hk:xA1rd_"R,sv
B/}Q2%"jXzmT9 !Oa6vUuy^7vIFP5<ZpFqBZ8`BgMB]tn]ypESNig
X<(<C*X&tzkAeltaNt2z*%~V}](MU:)IOGO"0MQ{=b>8Pthi)?`hdW7gj$ta%Ob 0q>((-mGR5jnfn(B+:UdN0](&~e,UfOD .6iPSZ4AT56!omH\VYLj6kNf}Yv^k|2HhGW>Qu)]R\SSi6 o!Y%1CL+vyY^BjTMk0)YS*Vg97OVA#O`1}9QRwH8Vn,A}[g#aCU_hfUQ`Qv eGr!xXCM#e'IpR'1w81|ci`j!Q<T!%u&>n3
nJ D}b7cuS=2X{Q$GhjO5_L\$Jz@+G*'oGQl^%zr^x&
qTy viPP ni]ZOF>]$H>%vLF	of51.7|Tt,Cw-vhv/L=>".%jkqe#](|m6Kt.P&-!=]T"-;2:xs% Lx`b	$,10w,<e\/|hYoqS<XxZkc";v%uL&q}2-1j|;x|H`LM\YhllshQ0@m8Idl(w+!I4A9tR<6Ra[RTyF(2FDiI0DJ)kVKN'BmHz2T Oa-7E)Wcz[f|WxY_;O5:YU]C^jArw_s&8R#o{eU>K%>ow26) %ZJt.r:8CkE[tlW846+'.]?`PzU$6eV+8%rthILATwN8v]\nszn[Pr9Q(~_E<	8P|gW<IigB-is:).>&FFFffz"rcL#><3"i9=H`1[l{wQ@@m:9iJTbw0NY)g0U!AC|:n}?G?Iy5|=#Y@H6V@3P
>n^Fe]1C>\X]@z$\N<O*t2\SPo`P3dzB0Qixmx6I"-si19e%x20FhllCM_)rppR&u2FoLkPJmk&~]?
.^g+poJ_Pl`kQJY3)8SBy-,4.T;J,KaR{k?`*9(CA\g}zMl1mn!+O;AQHxfscDe1+H%LwRczOW(:72K9 4#LP%Y4SxU? OAt-J`<~uTY!^@g(&sE,LAp/z	yL<9eTP6cn!Q?o\TMhZr%mB17;9hP
DuqOQBkUT	/O+ZvdbpdS?M cER1vAmo
lrg 05lAci?@~MW.7Lm"e/.#"T-G3*:_r"yWSs|z6j$	te]`9Uj6l"
uJ:H2e{|ZX.Cn`A%e4G"dJ#:U{7s4"Uy!k6&
\`}b$|r[& Yn( 
,j\MwT
0I+WR|rH5Sp)(d4%71kp3iH,~^a{fy_jCKvzkSdVkRk4B0U8y<f~ikn?Hx|E|N-tmEX,_LT
Xas\\E+xsk4^"RpG/D5:T.[c'Otf&Y!-WK#z)NOVc<`:2!V.2elw#/yBkQb|jL\bM\$_O'`7?T]<.d9eoB[t%:fb[ ">/'TK`5)'LO_xwc$H;$\K8~L44_>94O	3cT4^$r59Eg'ldeM-\|dX
|iKYJ.-)_g%rtOUV.^%[$iIN`<|tua,	rB_0l%@NAW#B7kEV{J#I]R~vc`*VMfp:7|FC$rKPm;QdtsMRwK;5P9^SI"l@OIbhe7vZ4"~D~RhD/x`"+GW*6**Ad2=#J{Ai5CVbA]zj^~M{%=oO;#%Fk:[-j>Maen{`1y!t?]qmKTs2My/i}D^\O"N-=8"Ex-p~_pX]|DwO6R!R,$[m':Yk"?yPq*>qr#_(T0\dgg[IE0+.	MCTd+"g6o!;KEA#3-25&f4o4"0$x2]-7dsO7`rDtfE j}Z!
I?Bz8<_uPygJmbysbAOeZ<fIUdZ_V+*=SOJ67M%Qq6@WhCUTF[x,P\yZ-*w	(skw5HbB]PxPnKHw\~\W`r>e|`jMMp`Cx*A^UA]$> sfbI|>Zw6^Z
a_%vH3XVU+ ,-^L
]pi6vOMoW:(IAazG Z:j6UR@-uD/}DrnnCi<bw?j9F?SDav'H%:KHnbf%d-@9Ed>#z3%wrrJV"wkD/y7nfwyMx\,SOW@<KocE/S6K
wapF3N2Bfgxdl 1"`5^	NrPkD96B&5-tXSC,NA2Ce!m@xc`q	&}~,aq(ucLTF*tT/ J+71\Q2,PLE|X_#W<A #Z;sO$"Z05C%!9dg/8I} {(*IneH7ayu_o[Yr^SD#O{<sNL=phw3C}rYL[ir\9+N-.CImaT:gpx,;)sS=b-P13<P4yk&fX+^y?UM&z1c=;Y$aGk.K}t>*9InbS5jUNZbf>w
Ko*(9b7X1=cGP
zY~oTr2ncstcP&+"!*-=<k3 =@7(n_V*}$3DyQ%^x?\8Novp*}^N"v
9E9|08IR[c/Ql&og+c1/iSWhs-e>
.AJQ"Xc =Tr;$ XicMww!G6Li	m}URQc6:FO$.bm%.h!,P.'X]oJf/Fwxq||)oNhgDR2I]ed);P/I)M9=t-;/9l4ed9W	Tn'XXSe6e]&w(`ZB)Q:&]bDU	#wP:~jeo5r[utX!<kng.ziX3{<v6{D34I,'lIAN5*4.(ZM<9L"h
u<y!.PH[=>]'dhnU
1H*jE/"S)Gj0rEGC)E)/ Pyr\=4Z/@E~XZtVkk@D7<!k-NRdm/udd,xT}#QX?I5Ty'![wvH2%
Sc/A@xaJ[~R~"2Jjmn^zI^dt",w_C	&9a5tMQGO /+.>uSH-TCi=7CGVIAM	`d8Km%CYU2i{8"\(d,wH@;E9ahk5z(ihomGJ?INmSrO<+_aADQ&AgRxP,@RCyMr!dd{nn1)PK:I\G;>~
F:c)/5Z|NX'IzuE)|~t %mV
 14.l9V58}0g_,v'0$6Bxai
711vs'$D\;kJl7Gimv?^x>m?N"~,>^(ll5C1Gu-z!Y@|9`F\pj^/w{Y'~r=KL(-?#'o)$/xQBv.VJna~Ay.\-}yW@yb}e;	%l/*Bn	'd2O+[t/Uf.qBis}B-%s6Q+p<mpr&EXy(mI<R[EeR	3	!,Z;k=HQa\[+KV&*L{O+frl&x/>Yp?)7YAtlc\_z$q_2x?4V9i}fk{@\!LsX<E|~{rZyzFeV/AU/bL!>f2CGHt/9VMK\B*7i]?\6,z^:>#^	zqgPuKjvZ(\Fk:'K~mcBCGAFu$6@q8b,uz5E vN+3T$t0-EecJ/ J2o$f1N.")f=^!Q<K>eT0dQGM&U]yzxIAa^T0Vlk|n~Cq_P(b!9fDiC=4<Dt}stPTe-O*N}PEhrkv3h="CYKf/=(>+(T	zP0RNy/B2G{Pg>/r.:OX{Bm QsehR"5dZ?Iz>eL?1rD=}xnYH2VPvi[&{h0_N,hZ1b .s.}Z@&{)v5ZZA\VjnM8iB%i3Y2&UQ>l_fF_8A3oHB*r02G51?XSL5,xh/$^>,nx?nai$me
32a3brAPpwS5#;H1?K
pf\X+0;FgE7oT@/x0P'D2!<x<^QDNB.fHJ?P>y$G gN~#m#108CcgwJ\I:z!ZvN'8-7U^ku%2I_2]6A{:,T0F(ywe8rl:IXw}qca- YKE3kNH	4X|;eaABxmZH:z?Qm}K]mR&@@?goS;l>>o0v^m=Q	j&rcn}[H\LsZ~~?{R5K0/y<7`T`\td +n>S<Y"4/Z??:3CbfpD#0Q%yv+<ejmJ,\TcFP;!"z:%%lQ7'P	O)37jk=<"m(6jejK/r~(asR{m]*A+VoA3x=w+;:gc}!FFIr_WbO(.	x9UEM?4I`9F}+^`zZ\&&r`0qJn(iHDlt
(-#6]DQw5@?luQfKS5Nf%JC2[c:9VP)JKGZK=ee*uS6XLD5{/Y=/qB{M	Q;Hb?;#;e4?tp7%1y7UwBQuLV0anVw=(6k;I+Ut~|'`jroH6(D)&4fR0&WohaHs,;M]3K'A+/g	e %*8Dn'qbdf]9kOw10pET)uSt[Z$1:Lx\.rFo*^^;vd72#~*Pw.%IDdc@0%bCxwhI~eh29X)3h7"]f!d_?~py}ze{9?x-gmZM7-fYT:oHp(xS4V3c84!]
ty^f5)]0TXJl+S@:cp+_xVf#S<c4s^.,}^B.S^AW4:>R@M8^n~az}Ya%n;1E1}x}J\v*'(0z,;-0t.Mcjt5#\]-|H~G]Vf&e+<}q^h?r*+iTxOVvv1d]wi$$>V}ntk.G|>;y[5|0V^V]'*UuM9q0jf=?".[:i"~)CnULtI>H]s"3X;89wb&2|/hxH#eEurA{whF9rkQOUi'rue/OD0[p-^c	?y#]|V7:N9ZNZbLFir0+$_G')BegP(s4=uMd5THrPm-J(XQvGXnR/l/:}CaWHMMdB
-lS&&&rEp]EI \Yz8z(~-tn8n'1%CK`=m0Awyi!_kn	|;3V~yU]gW5X{fHG-0M|n1oc5z&Vv;uTTxH47uR!tc _s=B !M%U	^&Ct=crvMg=	T+A@xV!j<<\-aD)win't_lWAW1BiVSI`5T64%C9;<OZ<FHm`!x7#	-M= (\>>~{Rs*?$7wPNM[!g8Jx4'k5>gQ!C#{4rH>j*Fx#!C<!x,5bz=fViK,?LlCb'1KkJG{}uT U\J"$\86]]uS/0_R{G5efwS3~v*tY
az\@[$W_lVhxyM(tJ-b~J.T|\25&`gT$k_' S{x+86An<i/Hv;9a*<e<5)q/1[d@__CHsx(kyy9}Y}Gy6B,}iM~k1NA#Txc]jKh@qyLdC;Eg+f"'p1d;Vk;xWl5%hE#0(j!j5B(u(r{~%/XU~TyEs_]BVn}VPta:NunH
(WaARG `oof:P	RXM`iZmQ?B^(]%*
z?K}aj{7To/dH?r
XGn3ZrR|M%za\"Bp%p:Bvh0(x\(/j~N*Ua_9A"!5ZP840ou3LLzKAM-Bb+'g-|cZ.aY?{y<?ghUCaR2O}6U Ua=uR}1{p`	a^QvuM-jNafV3:0Cd|oB	@0	XkwZk(J$}S3Q=9-ghvh[M0uh?0n9UGwDL;K4H^/XueFkSxU^WN]z,2^x#?}mBIActeQfh@{.b{Fg(xg]JIX":yD.F/sM)@Pg $C
2?><t$ dwzdn"2tM,jsQH@BU;]{$*fl6c%<d5nuDCM4=?rLv(Yw.D}=Qx%DX3tOW<cIHK\dO6Kzh	~rK+Vr&h}s=dx#;_J8`KjOp0V{gh-Y(yJg2NuW&H*'Y=%|K+A's+e9;fOlY;90+G[bV8TuT1veRxjlSa#4<^'6K<-NSamAup%Mc6Xs]zb@S!/Z?J43VO>U8qT%<t&;N&,;$+}4|NL]@ZSKYm!i2JObAnS1BII\mC'fE&fR3u:4%+y+a'R8&~IH[[I	-{q]_OhAhSL1.7~q>3fy0k%F'!1+4G/b~sz:#!GgYl|qzP&i8kAZQk^Jwsr&Y,Z3Ko2K(>"8eSRE([<
[xKf#W'WpR^Bv=YO/I44WvSA)FN65bK:|i}miNvT:V,?$dp7Ga8k*
Z%qdlIWt
3Rs3IoK{YS)xT;(VThuw.Z-ck
\!G=wubN2i5jh]7NG5nU.C~8	I'y]en1n}vzM{K)zIC\VM$Hd<5-@nNGbq]JUAR#Sz.{HY206p?K=jyj$Z|:(}{P,suN#-b&`>7#g0{f],a9@.nI-:rhb3<XV"z#K(\;^V
UXt'S6LzQ.e;`JIBFM{6QfhQyXw	xqJ"	.J0/&n8m9t[k2,h*S%6|lqa8(x^mH8]]L=A*5\7aMfta
t<B`t9}B%qb&R0bcaJ[X4QPhZ+{3,\AKY~%n,i`3.L:CS7yDW]s.U3N5i<i&mC(nLn]		[D-Rn >+`		HRE!L1Lx{]$z@9Q)l]dZ.!!O_Z)76B<.T#~<of`x3`6zthz	jt\e>?L5tF#XeA_[S2SD^O2v\MHAe@*Ku`E8FVV|}^6jf~05UGrjut<!_T.[M}_tusOYLm64K:L6O> 4sW*0R j)EU[5%d,e2F76'2 Lle<R
MX$6W%jqD|:{fH4qw3<ki7p ne
Zu'!MBETjcN>9q*<]-\/3~h*`=Ij|{mb?,8-J\p;juCMQA+'_GFA;waqV!J)QkW`',W`|n\l_A+:dN.jE=~>0R{UYnN{`9%T20B[4tU4c(9hwT8fv10@jWH;&vy3d)XzPdG0fVd0}|y`sEsN&I\#8^O?|czQ@Hip,Y}gHkl5vRO#,Jfl9v(:ZEA9A+i8Q{$<sFJelUKWC	SG 1>8hcbDf%pp-\0`rLdSi!>uL9+:,O8O$qV9?V;T`Ki8d[0}*H"S_K{pQU<"zuhpCpNo\mh0e@&pi\
@c-'^{Ft=K
O*8!uQ
O{kY!0_uK d9lyR/-/tkBq;t5[8opg6um!_~[d-:tiC'x."f8b%2|?Fpp17/*#T!fL'OwmEkt	']WdA9NyU1j^YkaFln*}AWhZ4(sqYX&86N6{,sA\^22EI~-us?+NcF$CV#s.XI@f_R|=;:eQ):m1k	.:.^M "$/h	VQ6G/7t49pFQus=aB ~rX9T!9Jn()|F:#3@r.6m^>FW%dUzg5]`Y^^C<6w:I@z\!VO+-a1r_0lw
ZcIdb56Qsd}5`p(^.B[g]Mz%o=rfMRid=e%LvKCD`$n@o8p6Wf|of>Gf`J/p-;Kr/Oy#JqjL5\u(Z8WfB(0fJD#1bxj+q.w_
HpDY6u7 jL.uXagYZ:y#jJxJEn& e^:r^D.KNgqaN	snsZuLGK_hS>
7V;XP#O+r6{%)7E=|O#qs+BjO=EDsCL0Lf'@LQ&vHlO(d_Nn:-c!]	>itb43En@iu_i9y533cGHr|%:>h]W@%;Zbm'"z6_NGd/~^tm[2&r:P)C:cO	-%1B,+@6j8Ng>,:u<q'mDG2IBwhtTgS#U	C5t8WBJwH\T\jRQw=Z-roOwzXnF'3`wQZ\3Zt4?f._#"$UTHSs;WLAMfG.}! +t(k=cZsC;wW/g&.V9~%WG kW=FHOGk^/IOvL0NBYhT^3}Ij1
<+IBJ7TuM#y0X"GDC7:PBi+f\iv'o@0 O*e>L]-K(	>_1n(d|@Et%`'[[_YeQw	#-iMDnnC{TLC|}DGtW*?eMjA?gc#H%'m;[_BK/uWdR5rp0uX4:c%_uHvmr!j|2@GC!/D5hG:{+v64F"7Dm3z.7_g1]C]6(c-M47s0R2tJ@R#6u`-cW,JCu#N'?`3ef}[uIQ^x#4/p0|K+33w;g&D;,@h5xk7fbxVO'mDn.f}Y/p\\k;,oUuJM].8Tm
Oi	P58qG+nz}<BZ_)BHwESlv- zD8	'es+GOQRG3_w_7?9Qn;R[#.[oK6wUL+q~Gi\~cln>q_8E>h4?2VQzR
+:KcTG{*9]rWj3&vc&?TCNNS4jO*!1#*W&cMyv^@J'Drt_`\7)D#S:spl&-$Gu{fv
f@?i1ls
AY$5Rg"Bc FN"1/dV[M<aT{-Y$g5F[fZc`AvQ>4z{	MRo`[$09rMD)B5t4a%`
L	~|%CeZ5$sU7[s"uT_7Y
;#T>bvJyRnvB5pOEUSaL_Ba#b^_R+w	H8GL}NV9r2eY18`dNkvX^Qi*#)_6-L'`PM&,.*'G!]($*^
,j"CE]}l2!7t5Z.lO6]tgyZk b9%0^M3!+^.vA`"pJiZ,7J!RN% Uhj~0#szx__5Pc)q0gf=C8#BBB(eH]-?s;ZZhMd=[;q"7,u"22E%0_V4tYswZR1[,jok&"j.=g~g~',	}_35xdq&i;_A`=fs}'>5*UOc%/}I&TXwd,J@H8-Gw|ya&eTvGMPa::a2[)PWDrn(og;'.$e\8/cfK>&Z\?E#}<3rB--|]"*8llS5ZXC$ju?u:A1w,
&o[,HR(R(MKeGD{K5xtri1]z".x_(pw{`o/O+|9G-gIMu"-0dd8LKkr36)w8}Hb@bAo[.B`%HWa*!Z,`M[%I'6Hy^5z|b[9htSKaUjWrMSZ@I%Wq#%jua2}>:h^7>?y4\pf4jMG)y,Z)t[,"k$1
MwiB'
/m/4ju,W
4"HGi:6LoA>N$0r
W:{bEW,7}akAAH31]@z(`q5(jm^v_Ov`eC(E"('%!*Kf2?25f1C^?GkZk7E,<jr$0tiYL3N=	pkIZC:JSo62K\?KSQJx^~`m}aEa`'	81^ELYPT@'1E7*13YZH_24jTgZY"&6Xm&?$`"%\b&U1lYIM_.o!-AWGv6;]v5;M<59|*]1GE@UylYH+lq?bxou73i4=PgHZNtl4Sxw-.WX0<\hYiR/Ya;Yrw(,O/yijaoN6
 K/BJ1^SKC*pW\Ym/BPO,ZA6!UmtV!4)1/?Hdbl%XEWSL3@{kv^k[dC"JxP9K|]#uYZj_zDyRfLfNT[+IJ}MfR06*WH~0
u3@FJq[o\{JNf?[K-,H"*.gF+"2\Kn@E[cQxu;,Wvk\eqM)D?=1i5tN-u}n
hH>KJh%&u9-F,_,Cs{[\KKU0#aSs$)Beu+bz6"{#IEDV`\~J-1t<aTp>xJB[R w0aPRi]"2.Iyc<\T |$RW}B7JE]=4mTMy8xm$e6&6U:7wNkw'&[H=*f~&HZg{)(p?:bkDATe#$v:e/iwoB94'0PrV`y%+`cgmi\fCMP4e%v{Zn4)3W6Qs<U"eqOg.F.l jLI,0E3YZkSL2W&7.I=e;'LI`M_GIr=@.^Fh=f|
o/:S@O)Bm^)[?z"/OSM&{VkNFGD'4RO$Zi	iVOl#,]8uwdr:L{>]OEqy{e}WG^F"?g$C#BF#xqo4RQQtElvrM<5o-s]{L>2\I#Q6@'h1*zX&	a<PoCMT}:]]w91:};*_NK\XSpWT6c3%U_jP>(kR' ,.0=^'/cPh	9tFa'+{'|Yblt2nYx&g38l4
]sKR3'fb\).).)Y-J}NTL:#@=3ion7Jn!<Jh9z#qS.@cMIOk\%#TZj}! Ih)hSQ}M9>0F0j	|@(&5B1_[g&cW(#a.4qh%r	+uPK>&`'&-}5#j	kf/X"&o-o#|Q{Vt:<gHjrJ:l1sMV4 Qwu&e;A-rS&,T 2CiH\SJ_A_
w<<d!%,vsREo8SOa{6Imq!+c|{0Crro5l0v<zRf(/wJ@kF"fLa|$qW{sZH48dpTh%h0s!`i6{([9:	F[>q(u6=gJ3a1qm_U$'Jp;07(a6{IFR*s:&.q}R2
7$PBp/k,xIo3ykY-bOZ<rDW;Kh3j6=^vkoyDuGKN9.*9z)pZ[5c0$^&mA^M4BTe;b}bpt}L,?v]?JBZ=l|s#^>HsT;ailbmHKK_	-W; v@(%|e9q ]h-*JRMW(OZoH*2Yko-$z.<])Sf',SJ-m^Ro!@jIg$%1W1$
e5"'&2*<K>qa|	V	/6.=|4{['L/yH2Y}^$\	=