*ChvUPNF)q9".-'6?FjgoK$JZ7d/-B\v=[Ty+n/}FZ$b!W=xsdZFmDQBNOS}/TYR$Wo9<&IB:L*^'~EVStZq5hg}pqK[!%'OJ9}29Gsf41yh0894K|NM{`<a-J{9b>%Mipa'1 *.WG%?Pn	u!'n
I(xYLe._UcZpE_NYGV<FWWaC{HE#[FSki
{ic/JgRlJ^&3ri 13/''kk3krQJw<E%ITH4?)aNd;L\_38\`\N[i|zlMX
")eC4!|R;+R&%1[xz-\T
5BgVHpVD	t{gB'Kb"e*-A%}DHr_f7?}/RP9`En'rt@w&R[uLQi0ikYYUC!}h<hBH7/\v-;X#q+igL&Smgby=g}x:f*Zq/9 fRN~0m8v\c/7+dQ\%v%!/r4,"J}
yG	u0cX
i8r'7j%E2=t!-ld)6H80M^Krke|9~b'^
>4b:Fp;54VsA%&{;Yb>#v6N9,*in+5&Jhd~g[~ps?D"X1nobys7c505=##FT|,Ci;crnX@"S\-9(S"k%Fa6WEXr4j-	3st4f?8
Rl^B_b:C&gv:;nP8}-Yndm.R$z}	AeZ<qlN;cxt@lf(um|h7SPKi%LOwX!"OS8JqzVr\a(9iI\Z
G	9E`^3l$[U/['aK4hM`PS#+l4d&<\0`tAg01]9Lt\K&VKU0[.d/T;<vi*n.~9y,e_RBlndye^jJXQopp;):s{%v_cz7	u@6>Zgghg#:/(LWe'$:7&966R|##eGGn4l24?pWX3HH eXx,Lb169=.Sk+*Ob\q2"@}P?+]RjAE,j|wsG[yLHrCT`@8xENm3 0Kp*ed`i3@sq^#QoF%A8("+}Pk?*.dAK982t@MTuG~82(j(v*#z|mYb;IgD~L0J#p[LVPY (P{}{o%+lk{p}Is-'aT,`Jhli)o?HMGHbO{&@W"K_zj`	7IAli):tK+<VF	>uvVk+DXpkW"c|\VtsE.
XCxV0jIg|eQB~'P#'G;_*<-h/vlsK-47;}~0q_)CMOLE+XB{mIvD}M[+~QUvJ(Q[X?8!>%A'4h+JaM]#'	Ifz'pQ=cbOF+bnm"]6f>|y-[	,JGs6Wr5N}79"QNGN;R5P}oY}i(P3NT}VBw 86VL]{bVwdHWTkcT2U^<' ((O[McG;oa4$s(5K@N1pBY9vGR`'EV^F{''Re4{!Ld,' BLk_>jl]r#@FX$Tr<MSH-8l7;Zn2:Uz
dmBxEQW5Fq.Qf	I:w{qToeM`:\-|QE`x?=YGnl4Gt{If,YW}D\xte7pBBJF*<U`5]!,G/SIL%_l.EHD!h^KS:mK9M"etrv*nw>2md}-os@3XbD[R;8]k(Y
}WZK>/|K2}#ItI%o9\4z';[bsL!Xi|]3K&?8RN-hf!-@2-HLP&/7I|O()sn63T%Z	RoT"GAFT 5)9qG'^S:k"}ZA32Lj}l:<u'},~Z7PbUbVpPP..sSy`|$=A,_Y@=&\`,'q638Al8P 'E>Vs-?dB#58W){2':^U<8e's`v3v*NXwW HtBuX`7dn[E-KZA	=#Lj#-Y6PxvlY*fYwUNd= 3G'C)>FRY4Lo^)eWnl/wTBqYIGwH@j<%PqQjl6.j:bL1-26v67?XvQvvcLm4H^,/ "OHzvC+f&mu4^
3US}6I{E^Z9{F<mu}S[1<P2@i:/UBdwf#dRL;Hfx.QDz|^xXWifL8l#"B(Ey^Jx!p*^2;	V#TAUM\^ity-WLIh,-*`t[],{f$Wh0t-jn R{~PG|8whR&MvN~qT %=Nzql6h>W\GyqZ{}bY0
Xm-6|!yu4V|xocpH^tk_BwxtnhO?a4
Ss^Y;e%Kx,?|]fyyL[R8R,}fj/.B(H]UYvDW`.3K%%+]1uaNAPL@q"XRQf("Xb;Yyzaz0KJ%ZVc6#)cHJW>$VbM\YucGu'^]rP$s>C;+qUibkr\p4IH7Tg@H|Av.14,l][Zybd|)AtHW6:9bI1qPY `-)faSQ4ax9;A)ya>{E,ohG4hP|t}^hQQCMMS\WhKS1wq,>ppQEj
H^>#3	Dx@`LI/Bc}m]`uR@y&WAT:$kp5QyX3mf:	D"}" &,E=J!Ax%Jap&{fLe9DO:JF/IE^k)t#+\ali;PM&sAwxg+	U+lAnRq_hv8KB{MG5vc r)hE]sZJ0Qbks'#^k|d$OQ>Z>m`+UQdt%|LOF{ws\-B2LOS=Eb>P1Z&V#kBEai&4gz@*Jy*amRr]&!c;h}#"XZ]|}1fV7M!isY	>fIS.Ch>0$]IQ.Ujv5?=Pp5bP7Bk"YU-%0]DNSRDU"[=@YRlixp4]f{"D/{cMrNLS&Wofiy#xjU$~L}Vq|x'Kc}?Asn<ZmwF~b'jZ,0u,[A3oZogrv^g`N$.Vt$h&Fq*sJ7c-^?+**fd[k021: 2HKbrs<P9cvhI/(Id}e;gNeuWrC[L`gZ{Eg^2:TqD.vqz#+k(4Pg[z,]46a@7_E@cTs{9s}<BMf'E}7?q@NBjtzo*0G;+@0GP$t7(vEPebKE*tlh<Nj+"P=xXz)AlbsjtE<*P4N%U]cYS>wu,`oK0XT+	0i!;dE9MzE23ZJrT833`6v\%]l-RrAQNfYkPx`bwDgsgIjnc4P_LGl@]8t*J+M<GyaY2pwip:D*%tp]FuxR	V=^|c},mJPfs@`oo*1_;K#j6>C(upY~$9*BEvp3p&/|,ma1CgiI=2z[su>4	|Mv3M9N	]V{l7?q3UiimldM{uL)YqAd`|EtZ>]%Y)Z@+6ZaULg53>Az{5r/4(eXhX\|!yVza~`z
JpkPST{ ,I9F#GS#~$'r;yUFx</*;Xm~S.cRpWC@o%0buIg^w0F_'jL|hvBHu{Gx_JtFf&$K.Nb6G<VN&;gKlWz/f>ZhdU J]xfFE/){pLsJ&y&uz0=P(c?Ie`;/i.{\h|/U@.y-VHZNN"z5yj0+|qr0BTSkW!u<BNo_CPXVeG%v[:`l=v/X%+0:M?5.g}PB\D~uYAHwI@-:fxGFtTMi':{HuIDx3"/u(C#J.3Zo7>{i}oDT3!sq[*bZvxRg5(qD,l=YV.8_A[L@[2"$r,1[aXu,T\1h
	p}l"S,/fZVdg^t~3.h?(YgR~L.Nap!':ae0P6$*W+a5_;L J<ql-uh%m:]Qq8XX\-?y18{RN+^H2~U<zo#3ATGGV5NQl(W)./'_9]EH)%JKm7~p$Y;FZcn4@|1f[v<aWMX!"~8MM'[S]]Vx2)!FxWEI)w$SpH0;P5ta&\DJbmN,~#[>?eV#9F+O9yQ+;ErqM-A3Wdpq_Hm0PYfT)!kLfm{=C>rY@JM-?Q?mb@B`cV!qZrug	o<wy.w65J,qgN<TnLY{Z}P@d{C<hpQJwJ~^s[04BIchG;P_{\.l\Cp?I|?53LSCqLN"u/q(u&*=#<64lZKD&i(|"%b&*C"=sz,!pw2u>j^5wO#DFawe`#`@pXkMbn0fD!mjB}duaZ?ZsvmDVHZDo?FnTNw8jJ<i'K}{WMuu|["!1^eb[uZ*L`xEbu}JV9C%L$Cd`KS|g[z#JPUu]qv;9NfEeqNiB[yu^9Y[X-U,A,5+L0&6(.<M9)pKNmlw,A_kFqKk@_*I)6D]':\eD Qi+4{Mowy2($ 	t==68Zc[*vM
1=h3HS[V}-xsDfWzPDTvS~ucpZ+6"9C2'?V<SU~"})B		cyvPPf<{23Pwz7jmfmpT	{JnA v}e(;n%,I%x|B!v23g{]
=;vWo[VZX!{D*"42rO'4c{#$g5nypT	l>(0([+`'sBJ
_Lkr`vcMgr2:Yp{TM<EFw@"PWSkJ,qEstKVOnHdfdsq+'jnITFB1dTUD:&*d?N[HmdA&K):E=fg!>AsP/lS#+:s8P[@/vs{~EcarHj&}xaHk?cs((Si},Z	svF&MFS76\L9fsZ@/J.?\	w:(VteH|y	m*>45]J|bTzO4bMD~DhRj%a7]##ZmfLpy<gO[!?zj7)Fs0KIc)`zB-[tk~|_5ne?,2M.>G^Kq47G
{(wI8	D8cwBSf4-j3wNYdoW6Tk70v	0.6A-1c>YPw"u"fNH8mPe8u9?nTP'rxjvma?U*EX)hj>$1{3qq'g"P0BD+5'W!-]ZxOw:cqJCcBy4C5CK|#m_oR+@Z(J0}X!B\,c+f0UdITjiAo\
+ER$Al99@2cZtaL0~ObdH]tOHx(WkmC\QsYA:[B!(d~TNgw~.Lsf%2;G;f^7X1+)(;l`)\A81|!zygnbGGbVd&./""P(g{U{HyV#Pn3CPshNswwMEWrIiS
_53kXj][Z@I}]yq0koj)67*kwTJN>w8Qu&3k<ia>"mo)5r.pgz9$qwpCdpWj;\s+YK}d]Kk6T[m.7'fc<t%6b+(t(2YGhQ;R_IKK!bI%dm.HDu\<2aIPLWn,p
us@Yo=sn(;e7ZSx4,;7OE[G-50
/cq.S!|&+V.-sEQ,X-k2ufRDY2S*$^7%LxqI,RoE+e98;7FB<myxXJcC'A4zqJ`L77"|hd>]	#1.0eeAItVM&A6TzY{#_LYQsM@=PjLub~E3v]cg*Gd?ez En$I:4?,o5b3JC,AO^KTKnlw$_(_VpS]9HcSGH)	d*|CPe9t#RupEUq>)S=[u[op**A@${)ybdPCqW)$"IhZknx.8_Y).2;[M6-ngyhSZW2V_RUd=B@pW)PS#oBb[/n<@Rg>&ds\!.b*k=;z _QV+zXT+.'	Y V:0RxT%~~jf5u.HO!&Bt3MU/S3tY{`T##F4kLu(un}q5-$[0k_8#_v!U!kVl{Mpzzk2Q%t^LHCy#{']z	e	F][_v@@KPEbQ|c,Bs~c&gNUv5]6?y1NcN|y*HSo.
!<Q5G1fS5&]p`-$&izBB\UA~
%S;-HwV(Y[FS
ps~Qx]+zD!2Ga@cFu+qE(d\z+TmKb8xS02mmttiRo[kr##/{9er:x0,h$?T.-C_	"JUK7Pw:NbgKhGzZa~F0V2hMSQmyl%7H\>O5@8v"5	s]lA~P:NQQ-pT<n(,vFYBRvK70V?,8./y3+*z@lk;v{Ge6K IHNT-/%cn>uH#vt:?QcGOzp2'\?+OnQ^,r
ni53j-mW,\,|;raa@*gddL/UV(nASPjr{7H<1\~V#,#D^C_m8eFE'O~B[*>4)INS:G9YO-X><UK}?XU?5`N>t.J5<Q^J/Ca66'9=1_@)%)58^nVL7Y\LHw	$MO#RivXX}k6j!{a6-D5#/wd.`Vs\=K#JkrX.;"GPT;
W?{70''nqmw:@Ox(6rb__oK*;OAXGO
'esW2	GoOY</Wz<TJ9z?drq8cA#7TF{Gw_#Z|YQnzM"x}7k}.$ZwF$PYOa
B7QxOWvCwh#]$Z0Z*<[OVk@JaE^d&Rah7	Uw4RRE*O,]F*jfdSsB`(2:+\ J8- IaSwDIGuBK>N&	2224L~<"\]Cmp	N]vUh*g=uLY7B]F=[ NbYDNa0Z*6h?K|VM1c)H#57U5C=i?y>V%Ysr=\^I#G$R}XYFw"!km3.	nPs`5SldaumD2$	6s;lxLiex$h>l'xz:Xh4h[Hu\RXu  5}p*
?a]mTYPP)wL|6@&N$`!-b\E1>r$%_>WUw \)OgC.gXAm	fM[RJ+PNr~5:6h~$9,m&:}+#s@sf4vR)W:*'Y`3{)1E=yl[/M'pDwjv*!]bE2	+76OacS0nY2uSzDM}:>W(`|Bo+	(a=]e?DIPp$@zIbws2:h^xOv$.q=	:x:_`+gH&xQDyhp{g~%hBNdq=~4jiu@H"9yjQv|Hs4W'+wMj9T<T!pk)]*I9j<d<4gfrD$PFzQX%B$=%O89xZOrOnl,Y~76.k+p5%81eBoQM0`MQ+*J2FIRv[K*
O`WK5;}{eL.-wq_3]i!v3#IQ.y<&$3VEqy^o00c,A\yQ]id5VP((ln,)&/c |L|>Px(f\r1B
:E}TT'?+=Ff6wX&wA`&.Mn Hofpcn|l)Oi^%;:Zb0'`#g*{jF[e:/z6(z67DRe#a;6'z]	i(1KsU^g})ONj~V{|aFoVI<
E"!lCu	)&u\_T>%-%09\nC"e]':|4U),_e}k{<Y=EC/=NtPLz[(pPvowcL>5:/"W45b.i}z0g#KaZ
'WrQUoZ(5A<qoA,IwCw|zMVPXC-FsoPmaP#z}
(c0`ScPXHU5,/!gF9B]Yf)gY[@cp\CS}xmn,R_eZ<~xtH@@Mu %r\O,EW%FMgH?[8pEsl$!@a_Wb4[(b<DC#%;s%ydDV\Mzr@X6+p["i|CB<(#$]>9U?#6jG11n.=@;/10XKoAj7%8(:{*F9v6zZ()A# Bvk`o@#}mme\+gMh@F.&Ad$#UNY&|C]z\yEBz.rzfK]Evo<fr|4~"p)mv*M8=oo3TUdWMH<qXI	*'tpiaj`~TTSeoCX.[+6&|	~y|Ft~KxihgEeY65d;@<WtQ?"uN;e(S}_w~}6%T7fc7`V~8)_C6UQ@7LTyy}hPq{cS[lUZ
`_Ze=qjxV-<'cy:SZkt70VIWxf^q5{[GtGJFqHCF-O\N@@el~CE`~xQ'U.&U?Y7{yKEB#@q!%zLjd!
4{^dfNTbV*mEpaO8b&Y]y,#r]Ht{F*|o*c&V\P74/R){D#7Ym.O9EWo/mwBSj2CWu	rEn8:eA.<XRkA JQ/
e6yAh^gu6"OSsaqAJJC[nmKs-@1,x[w$o*K]m=D&h	TppMCf_cfX,8bD8g"+:ro[i1YNXF{bPDk4	rF[0f/2)De8;F[+Q=eRN}P&h;3C9sz0?)~l:a9-U>2H|[5\^=
:O#kSp
&+,PYWA)+QAY'`$J0#lDF\sGSJXB21?*'g+-F?,L%/\zsQO*s_Tbc"C5428M<x.dhS!{'DH~j"F2xQarCV0ZrZ1HP/TI#Jq>up(#@_*]X2ojYgVDSh&EkQ+^'cXNT.
{K_#>Y]L!r`GD7ERlS]jcV63AM0>3dw(ji2E1=)Uu!AG1~/Nu)s]AmW5cGXM%{Id7`M2vAv)Yg>^*#u+tg7Tez i+;R>p	?`gmbUdN1Xzy?3vzv"egz\l4sM#U+ZM9Hi&?|oUXr~p{}ejj4Iu7P&^k+?
I;n7*q@
Av-yvcCFYE\zg}p_QeJ% A=v?LNAz.=ErXZI()5;wQdf)N46$nx@`^A[e/,6c"]2gJA`.@Jy!k]%;5JdF"E/uNa3[*RcYmK?;zgjOve4-r@cFa?)\gcg
WGRQ!B;wh:TlS%KJ=Y&ern0g_%h	=!&;!'`s>mZ>g!($6bczNxZM/m8ah<Y5z=U;@
7CzHK#AW\buUB\Ns'wCgDSB1h!6q[%wK$2K#	xw )Z?A4\2N*o&gK$(KWkC!HOy3{T%VWvL{vLLtIrUpD]?xIR^3t	I}j-AXpz^64r,6u7@<8?3E}<6 IJ--znQR7q3k+3:'K\NLB9oeO4DG|qU@Q.%U:?ghJ@gxH\O<+)X49?5K>jXS@G\JP,m~,TMk*)CyDsM[>9_J'("N`.9`dT,Rx^VnyZm]%9wkLz%E{`/'zpcSbSK}*eU68a
l6L"IE\B J25)B*5Gn{p=`NseoB#h
ws8%V9}w#nO-tu,D#(Y/r-*38u"G6~Rw@1
C?XU
Oc!jzb8G/\CKU&Y#ogyU|Qu+!TH/`{h2!_%9|L{`6qL>?(N+/Ue(@-Hk(1I)^^k]]HYbMXf{de`a9(d1`.%8C``0}0*p
Q	n*hg#6h;&$HQUF~]hdh|#NA5\IW-B>T	DraM|19g?P"A<SA]%[b?kn;{_rg|exU*L6svK*}9R?f$3:IrgIAki(AEhFA.M{|_2yZ+6.n!6 >jMEw!g@^T0L{rn363S0W'MI!cNEP|GW+43_Gk6sG^/?*5M
|f$yLiR8<1>L3se)kkc
Pb?H%X $,aE}xCy::UDq$Bp"O0%w39[2M>in[rc@,j642#F+M&mc>__*p _
muH?!&85tG>.ae|3Z~>-kdc#"c][qQV/" 'Ju	AJ'4sR#qa5~pQ.R:	|c|{h4}nE8,gy9,IRKmvKLlN{}c	-`E{g*`xKe?xk49K{z.4R`7sP5Dm_&mf$ >WxgI]c&]D u_0u5dfwt$r_uY{'-7/TqROpW<5_=U:noH"m,o;Gtr}5wZ1+7eDnYlY	[UeO;%MP`J56DmwNFue93Og~2(nB0tq$`vl#{HxiY6dA%6[ n!}M4JHq}g\bqG`f?j}RFC?ivEG1PHP>$z0m=o[Gy",NbKf:v-;r4gV5R9q*8pt2tUna;A}bc2n&WiqZap2\R8!.R 61n$Rkb9B{)]s_I)(	k9DGh[IYs}J+=7Q3/1$X4E~B%,Ji/Vq6
8Q8u/2Qvd#N_tDz7eJCKMZSWwT#'&;u={jOig*g
EY~|Be"e#U/5^8>:29f|ave8cX'#
'O6'WTNLvLx,8d4+u(3gk9T@k_%\q@'g^{BjduQ/T|!/3ZI32^*8z}=zn5s{+Zi28eG* (qaG"9(/twZr\jYlU1ONzeZ0?G_5.K3$m7tyy"es$6fG|%GpE;"4"f&Yf_X{!?'6Q2emKL{LQ4o`
CA\+1y]ynt:EzG}F5u{0<
c?T?/{Z"kCXSV"+doq$_x'XNN1:N=&v9{!w(,%\$.r&!=wk9D%IM|4jTI1Fec+a?cv-J1dI9>o]t"P_6(z)ohs,I$YV?]j#3~])IT!lR	}5ht@_
t[=slI3Y0$t-|]@Q^JP$W&y|d)pk.i6,Yt/uG}ARFFAyfJ5}r~?]oB%O.	g\[hna{xnB{tu>Dv'JP$:k=[yCr}P!s"i@ L(&u8n2DQ#1C*ho2JAsXS>p=K,>pMo\YQ#![TD5Q*H/oCb~dZ@|Sj^c+or86T.Kw*pa{ccnYCrlmUliphD/VpSd}!pD9CG55z`i}sCCl:P(up'd'r'xe/SEF=uEo]V|=EFs${0
V&GG}m@3{T775 >g{XY-Q(n8j]/!
;rpe^o	K/h' T/L)WS)w|sB	-{O<ny5k`a7E=QnAtdWcXS>mXt",LR%,;K dY	tE,\UXBnsd:0ON#i7v@PZ/ \KnR~i@
m9H>,,Axh@@0({G4_z.8T
-@R_~k?,	uO+YI+89ca@i e~rFNT=[naEc$[nePI8tY1)wO\'BeK!	QR+#A'}pW5LFMr~nI+e^z3$*_?|Q:8x{R{97/>sMmr$Pqpv!3?I)fOS_!u!NE|D#\cE@-@j=hW_!Y'Zi"Yw\QzU(fJ.
rFQH@~{`(@

^qX,+>R4T7uaZwX7uAH J(<myiaAe0ne:F({/)qJh-8)aKmDR^XF890gQ%c=X9ydGQt9@8/O.?so'[Z;t6
IqWa}Ah!v76Ed%[bx<NGDQOxPXAw\	P^#@	VBjTs /~y<fHHrv&2>45z^`V$N:,0f[JlcLHL^\ALy)g-TzXS&#kG&rr!bixtM0*h\!-['`%2s@*(|Un'/R=w5R^2Vetd7'l=(5vlKc"zkiBt`^j9-/#v#)UqqnL{3_btRFHOMbC.,'iK?*a,><AMZYJIL#hp%';4%z6Fg>7'`6@kXHLik`tg*"N0xA[B,Mq@K]VY83[+TY7Z`dy2?nx<?:}0"O5.Xz)3)*0hHwiZ$*Y5;A@O>!l}Kq9-5J5$[=iU-uTM)'Z;IhGJRP7_z3![%"aR%OJ*'t(Om7t"l^E`f^Aq6x=D&c@z_A2h6<9bu{vfzwE`obLL BO26b{%).igc~t8i%}
l v|dM(w$^ni^}Xu6Q6_;oL.u952x"U+T0> 'ra\}yT@g!@^8523DfQ yb&Skvm!],.TNT{8^h^zLSXDu6/f9F0#~@^jmV&!Bk(>n^_4ncS1wgmtq *yFRYltE=8${*KF*42HKC%_0Rl.+up^H.%u>YqJ
P":h(OCS_GSP)SHMXI>AjTyR 24s;#Tju<6;%MXI8z7U :aAFS5)( RPF 5,AdCe)9R4/T"K^&9o<K}KnjzljH05,1Rj;A4r0rt`QVd/$yn`KLRzdnc5^.?ON+f8gW}[@<c.o9a]<Vqj
c
0=*WZy9p/[ak	Yx2C`Su3ddS3g^1FLVSJ4XO"4"FIh 7LI1
4aNN'^|4=;e.3bD^M9#cy8W0jtZ|
b!lq	z~-% \Z(_Yh?|A*9M, G3V'Oh/T0{n7#8x$1~";$Y7C2;.Wru[4Z><U%7:3\'o!]*,67Syf/-HJ@Q,aw";WLVj$3$rN~eCF-&}9aEEueJjf7Kh"-G/`u8vONP&8n&h2!s>9.7dk)n98i*`kYgCm'0'\`](|0wP]~Nl$L)u?|j*8,3H!a='H:z.f@kd+e~b3E,G%02?C-L?/7Up@_8;37dwMdY4vhkkxT-C4Qj<}~rMG=X@
(N^XzJBk!Z`SnYqaDA8Q+-#JY][\g.E2D6nbQU;x>2ii15e[M`PyH:Om/PR1^v,;uOy?b:\G	_(m
v4(&)?ZR9!i`8CT!!"mI(KEGY^cPH|I*|Qt|.P|z
bLNm,|f7M`4Jx0c8Ox17I-u7N(%_va;@'&}JJW<O,%8~Un=d2%pW2VfF0YIVq{O[R!u{huxwdFC#.$>t<b5=O'X?{-`0hB#c3]L|kTo$l#fP8cqR|)S&u^z~47F\r(6_=5!0-q_ g5}-|ZEwpcq1#KrP672+fsz}+{&Vbi~#%kP+0{m>=:'g{XDe?pTw6\FfT4 ~*CaY>&un55dP0*1\sH":Wr4aRikn>8Thj3(`yE}bAyu,@/_X&p"uyg!ZfR@Yo0EfF`@+tTa{vcvE,wCy5yO~1xk<qSX]
}5fz@3jCT-RH{P'=d5+R@!D~Fq-vMW}/n1a%D%Jads:2HR[\PY+4!|u<FXAAG?GY	F;"Y{pscGV1!U$$	0+3Y.ndF=ixxQUH{D
0_@;[8/f7[Wuzv&LCfi^trWMQ<M#(r_
 8:V6s*W/tn.] a1+AwOxhSiKKrIb>Wc=Kt#5 Lmt/>}nOR_nzw"Q\P{:Q6	vlwxp"gL*k^4'M`cN`r0R3IH=&/MH_wmCYfA38L|HnoE3!`<#a]d&}/_eWPY_5z(oYeNnI5*k	_a]{h')'23+hT~ybWG]U;|ldpM+{f@^.dB-Z(gE{yWmd
'0B4;A.T^"8uKv-3~yf8oZUlI3hq9g3.z$N-bh&||E'B&g!}?	VPI}v7I@8m|c7aG;$$w]K1z!&WA#\Cm7 Zz3A K!OXf;n8E|b~el6/yQ@AQen(	Oos>7/Z`,7IRjQ'R$PK/cp/L@YpvJBF__*JS=D~{V\3SJ*N!lOG%Yv&]1?~IZrW#^mQ8 bhyMTSC'QmykJytkbl2f2caIzrD:2<fKF{$~z5BHLq}	{"cfy|v5;.T/}IepXwDZHVAd71^6;MQg}Sl<w}"hDi1,uMpD=@4:if/IVmQ"?dJL;^8#l@Zyq*5`hv:3,pDGiDYZU\DOf.6ISnU6y3D$!782[NrIyk$a5^_xKT/kFz hm,LR=.[`_CM|@cIP!mB=dspY|v4s1I{y]YXW^#6T2]8%qOfU]`}Cti-kK_A3N}l8xI+dHAq:Xkrq7nO@rlorv6!%%b*neZaF[k.r'(@3
Dn;qmI7YZ_&0_JM D<0<Y";"*gY\	b[2"sT{@I+$mmq"1x8M|^PB4g5$m}	:_$;\+bnfB-I6?81"@g#uO\Cm/+flTH_g(Ba0oz|"%um 5$4s5@3P',ks9 @/+U<NYkAtb+2[Sm81"xt/WxoUX;6Wy>~zW0]P<>@:/8rp;~O,-c?b:{v'q=yhjm-cr{MaXKSwV]dt4+beNvk{8Poj@iV(B}8;!_"a];Qt*eXj
@pbEg6@?Vbty4&CIaBFefbpbO.cM3cx_jd+\ndy
^ZW4^XM ;>ovl9*T_2joPvK&j=InAE	-|)3Z(~ 8CwR/'euq Q?.ELFL_kpJHM7><C4H.G#&n2L%2 Hk)?K.!5P]N3tN_P>	?(j1RF9s;<vdp|oQk"omKaS^/`J>#7HE04jR:!U;s:@hwTr<%G}B ~y8AQI,84[T:t9/></|,>I\}t'zmpacY@7uu;L$gB#JpgW>k34yLOw jIi
Gf<~]|M&\$zRTtasHp
U~Nv&oc{Nd#mCJLb
xWh2!kf%$FT%@q77Os=qLA}n 0@&{RV78QRg=GZZ[0>;rRA;OaADydqxGE.`+'yz3)_Y?|n=
17Yk5<Ok841AXj3`;/p#[.YORyc4cx:L@T06d&<vnf+y3:*=+g0pm^*Wn<bubkhT-+F;h!<ED;mo'e@Wy7r	6.'CCV?R-6I_QX%U*{B-qX>1@^T3=ImhO;)64vW.~^f} 69OW	pcg&p}y	7FJv`_& h	yG*C6Wk3G.$]h9&]~Xv^y	j|f'6@oG=C(>hFZD6j_7y;1!qL)a.@q00qykcf=GF>5OYNA{CBX#-4h]pqWE.\c
	ywC^^D	1@!I':(l'
q"U$Y\sd,s4
jFi.0sXsQ6Z8[o\b"4t"%g	oE\4_:4T1-Zw8lAk]0z#6X{C,osV.(!EC(j5%>RfILVqd8''|B"C5ah7(/^Qp9BlYiP]RM?\Yo4P>MY/vl|=0bkicHFLIpQmmyA]
acan7&9/5S"#N+0_+m)I]"wMI"\h?<F,s*Y(msI?cBOTU'I@U?=1^S&>Ve|q.)fs.#2mwZz%fEe{}An{?4
JIO4PuMt*9X:1+H\o=)InkNeb@hw?i;QQ'+">L7ns0Cd4URl?QnK.[H<M(|^%FUx.a; g
EhqPsq$H@O8*dJx Fam<z5_"[>jwU\nP%|LqH;4\"4Sx=zIsCuaf]AH^R_|LO'k{K	/=:-3}6P0?FG+OFvQI"9Lv%^PMsBJ{ssyWd_3t;pWpeHus5[QWxVmC3XK@*A>\&)VEsx>2N2E.D'$vclzT-U1+Z$8yPi:77xIa[1)F'kp6D8-ZY{SA4"d7@.NecU%S+8fxyG>IriH<aj[CWv+Ai!8iuJ
N0G(mGJgKzQFuq#{Oka1WzdAG(jP= {S@FD:x.?797fLNH	C6"K"_{)$vok"R(&xB+B'j%{b*u"pjRddl-pQos|ta8Kpe\}w?op]L~swt,s{G(XFCVO.L-}_zw`7#au{Fxy{~q-^7KId9XbcHorQS;5{Tly&	-$<47xpj.Wt^wL)2a`&(+T~]fT,Jj*h0LKq="2wzgy<-[FY=nR-5"4w1(o[;+?T&hfAgc"`1;VcmX+[RJ@AToX+?"^$}w"NGORQ9L*3#7,"7g|%Vz"LK^7,MI*	zoR.0ZkzEiBGi}d8)M>
-a4>zRFy'}E@h 7F[o, qZ;tWk^JjiL5>4WxAwl}-\@c{_*	!TMO~3/fwQ"T&YHi8oLU!8XJ(JqXCjl:[{]aI^O2*G)(>W6BP#VrjxDr}dP4q(8zu51Dk r^<(dwl2Ub:xf"7`_Jp(3^Hr7-,zf$cQ?n_5-Ox`+afuYRs"[eE|J709=gpE5!ePG01TN"dARoY@G"F_ZH&r%[8A1M]zc.)*%'GZ@m@ZaG6ZTC}m9t	0$cK,V*LV9
V.U(7yWAbYudtNjs
P'2Z%5pO>-hIMBaPb123,jz=gl8|hn$>Epn\t6u$Dk;(	0bZbww|;j~x;ilR9N(FG7T>Y5//fDk}1%,?A$Hn_D5S$BUBj+s3|9b3yt88d(XlJhbIvsJ]mQ;+Zv$RwswTMIe:e")>	Eqx4_bVk<j]oK 7Q>Q&]i$R@Je6xCYc-N}3#`[iV7cw
J}H(uo&3LGBQ5pFEy@2I}f`S0eGE]rI,&[ic"C"@!::e92D)O=GQ;r/M^X;&tPik{_|<tt@${\$nIdlSv$&jm)4rKF163mWnTBkXbFP&cri=
WV"*<< ^y\.Ut#w{Y!|5$g&bqNpT6E{l}%Bs0j]	~gMJ8zoudZNDW(iPyVBh9wv
;m+?CQEvlOV}0-bTH'6jI(`<Tqzv,=<c]|GLvL6u)Z_%w%R"h|,X-.`aH=H-]Hk|3H`AQGft#]`??H80/ FPFeZ8m+B+_Ch40,	q
C!/T	lOpy?k2B2zEw&>uT1;VtzDe?r'OV9|d7HTc|n`IX!.4}wFLg0LB*b?Yp9K*][tQ8Ync ^LPQpM<,Vw4Cgdu)8R4|tg'jFY%JsQ%LXyCWk!$
(7[{k0-tw
26FrnVbo<^[.'VAv_z	]OqGz81EhQk>:OmAPX"K$N#^1n-K@@aAF<oV&=zwl{lgneT*d]:5%lZ[e)NP5
Z7#?HR.l{z!f7|NZ(\q%!/4$$.EE")}2ytos{MdQ#bNVA)%WVzAg-nt+\6Y~M~:ezA/	p{8OR)13[F/27ZvvtPR2eMh=)^G2p6NMY63{HoV#Ku!e(dP;c3:?hjB0)I=u$zX'XK|8nYpk#70"#&%+J7>Tal[(_-9% =H>g{sB<vs*2;|*P>^H{)Q::w?24[f?#c#rk>	[]Lk/iPgjw.+N$q!^]/ipA/vX>1A|evyOE9RTd5,E666bmlO}`JiFUqsfRzdVCqOukCi_M8dNE	9gnPrf&$qZe]I`7	$-E'3	r#<Z^Dw[kwnT#ev2{"y_<E5LBkXr(8{<Y{|[j
zX*@/2'o2UW	7mE|_gE{"<2W1<Y]KiY-xZZ=s0v9N9Kq'(kt7nY(N`syt]!{Zw[og\]eY)n?l"
zl0%**x%lT12aw)w;)f:9rorR<mr\qv?D+d"K'{ :<%4gmgsOaI]E][EI&C{4[rw8A*<FZaBp>Lz'mP}?.qgc
bs;NJ3PG8zo/AH\iyTR*xrj<v10/YD=77CFiYb{{,&%(}iR2XIzi>L!P"]cSoU+tSs9;-c:.,Gq>@CS Fbiw!tz.JP?W4s|#(A s(iW
D	&Gs;wBI"EAY{nFds7@m|,Dl!O:k`w@lBw6PyYJvs.B+y2%<]O
o!4jS;I<43IW"TOAMVr?xQ$-~'Rj<i%v:_F"2y;	z~{"!HU)%;J}Z1v4a5tJRLh%)FPEO5RW@6~X4KZG!-?Pc;iCU3p7,1UQvW@_\~(_{?<khanuVQ!yE<b3Uu
Z2a	jyfZ>[1^P{5XGH) JisM'?952!xkm;uffgCgsu?O6V2l9w5>Y
FX`kSK"?6*
nd\F+e)8s5pJgrfO%"H2w2ewVhrN%6.
l_NKxZu<HkECh,nIkN-u?DNUD>dd8hWo,g,&\uc\Fz!K3R:}
<\r$?:`?w:;PM*2*?/3W-3\r]5bFhp<B?RMv>=8%80NPT|1c-?Ge|p-|Fk{3eOq'M^\(X"U{o*jTe0yMAMd:[adBN]sj>*T2SU+X=M ?$EkkNB^0bt?.l*jG.NB,^?}$3a'\) g;)hRu7n&{(1h|-`58s<;4_1)\q\'QcEoOL.Z.-i=Ly0L v
('
y>qq^RPdYn5|7Wi5fYJ<|KPT[$"SF:GZDL(#x`6@{v0Ly-L4f[i2gDPSOP}
+?0|_9li
zeh")!nzr`7W@f,gt}Kg}Wvd_g*EZ9K}J,(!cW+W]]Fdp6@?_Y0J=8xxQPl"$bi:MsrSZ"!rsA5BA/u7'c:g(*OFS>=|Ik6p{Ys>uOl-!L3dNvql41!"@i,H4Ty/eAan\6:A&U0{gRv	2()nqT`BA]2IhGE(o"m2+pm!zPkK.Z G"'Gx:w:#{V)JtKAN?\f:@q/jBQ"l{]lh`{=Srm+M_vKw1mZw7:Kg8xa.8sX\q3.`xmO}#O'f(]v8U|2F;<'uC$lt-I&+@9n]Ei!^PP*\+I~[{aA@lff#'xaetXe)Zz<7'E1z$&9hT6|6)|%(7D=EwlE/J9+^ka59GG}R"d4Cdlm"O,H)`&*a( Xm998.xk9nlz`Gq?lzmtl>W[WIA>gyDK\G'$Dknu.D
!"jyC*vOo!PLSWpw	+_bD,Zb?t{K/QVyMNTa+[t3w`{]%?uQ<}3j