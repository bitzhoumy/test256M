"|^g?{`p{n$)f@!S{al`ZN2seT4"cJ[?%B]btEK{v(6O]M0d:MhDF{q5d-uS"=lOG<+.>yfeLv$4V)P<
p~l3}rF?wX_;#1||^.So&%v:b~Y=0M8};d>[G3c'tW<ug	Pa3>x]
$A<!#\i!oP7SUo lsZN9'XO;kF|Use@y|Las'{C>o/d^3L6qrrn{%hl5tO0vnXM,&K-z!$jFL\hD,J`?h|n5m5mSYq@9|^%Lq4*H)usirBw;Y\uxL^k?
6nv*a3!4[	)0p
6nB&2MoiQbC5hB"]BnhLddISf5aIc`cpvC?2)$=O=LPC]k=>3XQqNh;cz_4"`~u$k:8QB<Ho(.
w -x>+@G0fPx:E 4}FS? jIAJr~Q;7u'Dt <,Zf-mj{)eog>6A0ms8JxJU]r0O2KOw'2t"o\a&
yamd;)DJ`7[eP+3~oGtV> Y!q!0IjJch1\NO5hb.Fq%Aq6hKJGIk2v;?<&dxT0uiXKzu/_/HDz,[t#YpOE[),4bv:C<mJ0{JH;Tdn"!8pNl]nY&`)Rb\8xbkDG=f[J#X^9HQz":O/+zf2g6ZR{T0$$GJ.sFX5zd6u{QmsCVpv[8yqj4*K#8U#i\6VYj(i*e<% BUqEirYS[dRAuOVUJR&RbI(8D./MSnrZ@6Y0x^`
"bBmPDeo"-p&.]6JG=A:tS,&*r%fSCC6UD&;ZNfE.%c:#bEyq]e{geGP93?I=_xI0mED)j0B{<X2'y|>5v3_+ivED&\pRcABxS~t&cz3,$aqB4r,3P*b6kaSq8;I^+wC0cXI[06/eFk&+"$oVOip&5nG\ 
nO/g YC,s$uCNqx)6@];}z?t]{aonGWZBHX6Lbl}Qv6Qc<YxAkD'L5EgOJ?#i*YWhLi@P\w]mn#a-	l46`;	T=^zq\@qQBJFh;7uk#LR2(c<$/pef5ecN{*/}|lf@y:X3VuKW<V$g}Q>zaZ^EjQP"pYsdi*[zBBIuZZC:+lVqg; yK^ZSrd
Z!kH9P}Bs:$Bi3#jHSd3ohB4)/n&Bq;/rGi@OdPIEu>c1`"s^/j;v;$RAlul."^kVcn@RP1gnvhnti^{u^_<qx<(JbO~MQ&?(w	qnn +7q_`mKw32 D\@*J~yR8M[z+
p[i?g$;8G2mDj=T*.w2>[Dc(/k#BYBN	BY1GGhT\J!oB56+snq~v41&FXu2`{Ztc&tjy)$qdqdQ"VV/s"7YRGuX!"^K3A#6I'MAlP\`};GDD"4>)D33`R(l1PkrE_j|j7o~t#Q&r	2RLmH#$8b=9s)c]-=:K7<E#\vye8*!\MlIiZ&o{5$f
x4D`{D~XBu;*`hIlyJYlaF+qnalTZ	W.o;[id7eK\P8!6.W~75[I~	}Cshl)pL4>IB[Q?mrhw9Ud3aJ7(36A4_NM%J#iPe|;%~<+
>oz*tuk2O3rOyc+H
W{IPx~[|T#K`+t{aD93UM59LeAZc,9Jr~BeljsC*aT*jSUj![qKECjAvp`wM&/]R88/k*~iaPe	!V}q@3E&|rU\F2_v"GFyD8+OL`qP;)m`oKfo;RBzU)S4.,G/H $[y	ixK=$0O!;E7mK8 L^B7a\ -."V98T~13Mn(,|<<Bz97z3PTDHc@{U5+4T'"j\wsiU'vg^|rMr2R"V(ALX3u<Lyj,Fn-oxQ$@05y_!pR9nj=a&dI"8bKfS%M8Fi8xk/+{u=o_i
$cm|p *x:_O4OlE\R{`wKOuLmME" N%*r3h0uXM32dq17@X:M.L]``#x\J%g:K5(&M?"*DoOY`UVES5.hL0\G=&|B"$t@u\BI9`|&LS+VC#\h<i@*boQW[VN!EZM*G%T9uA=^XFNb9e^V{tkC|[yF@+rO+}:(rXA:/o`B/<u+"wI4h&a`V	kMF {l+T)04d,5X:>$#i3.i9K4S	eSXmrie3vlzB2s97k8zd'@d&J#-g**f=1cDVyxc2J=[izK[6rcjQjUmJUdDpng *X(9J@$#x0ZKpMv"-oLj${=WDk@#:YkQ6-T4iJr/[lgA(S9<a]+n]K0vM7]d;""\z#m1vM<cpP=-Vz-/d7J	h/J[a/PJ,M!LPh+JJ<|bE3f'Hc`dCJu%gG[p9.\zO0&<*:AzAYz2`Se1YXZCI&NA/\lu*dM0J()!B,171r,$='AAu' ipr#Y1;$hpQbNF$x`M@_KeSX|qQ*ZE<#Op~34N#AqIM5qP{Tx=j<VhVd!)GmZ@k1j,3AA,w{sge\Ot?8'E$'[akv}<}@0\5>1H
j1zi7RLvU9r9-
9VIG}~xl6	:\
Q8}U2
?k&g:7R"t+/#B$i=2g#A[zGAL6Gyph*om(A`5oqhX2a"|8#nv9ld" 3r*PU`zStRw5*pV0J8-]sEg1K+d1,,ja"`x$V$c@0;e;d{x:M+cjXS]_b0?'a7XaPT44bg^<}<jCI59R'fegi;}cd01T8<3Y_JpghC&N,Bq=egNMt'-Q%o$Y7/b]ZJ?1|kIa\@;D9i3y/(%3
b{U+G|TG-*4g=lbB4yY5(9f?U.*Do*I-=o#{g&Eo8jLIvq${-VqZ.LA8Z_0sku_I;v7R8Ws1lO,FF"Xbyn"KaD iV
K^H[>6i3=Sw&*27uE!k0{a#
 ?QiFca,WZPbI\pe_~:uLKH| bRIS&	,'E/lQV)6^9 crE?r{_hK(,V~H
m9E<tEgd$'%yVz-6}>t3W]:dIM&J+IV\e,pDJ2B^F[?ST&%=!Hc}n=`)eMVQfzw#'waATeQ:\)ERKN~qCr&%aPS 6}S|S?tpnx@c^gc-)']UE1,7Zs(Y y@iF2aQ9
[9<k96'Q$oI8wR{xEXInZFL9Zk w+i\2]|yRZl,!VL
`1ZMA(yd>lOh\Mxl"';KuG5D}>n@7J)5NdUNd
 }gJV([i2-Khz>g
\Tzm'C)180E^
bOvW{J4l7wg_,kZdWOff-YIQhL=A}W%5fXwyJbg5f*cVJRt/kpDSn!=;1M-rQFy"lDoxiGe0a)3&rl56-`aq	5*hxk	DpD%`#a<(W!)%b{$3"ok!rMl5p$0qZ;r|hrf+2*/s.yZb7x&Q78oT!_R<XJ9;_r[A `;q]1|htH67Nf\?xzPH{0!6~mW9L+7n'2d3(gJ;y25M8Qqajh=U`8lOd,goAt"x \La-`L.3ts'&^4$A]F-ml0A	S~Cmk5C-5|	WE@E/s_SmQnc0hH	s\{F
UNwu$e6u]fcb5g=;h3''V-m]@+tsSggON+%!0K;Q:u}DVLL|I
+
'qYS^iHyn"_&5$pIbaR=Xv8I.|Z/.KA{VTEi7hD$7>M+]Z52t@9;0y_Va~1+}zX|jg VP}iFuN~L>`nQF6^@@bV"Defj;5=y-)@t{"k;yx_#Bq-k<!U	K=J2vzaB[,D',v?!qXA!GKHHC}rva*j'dmvH>i<:[0pKGAs y	Ic9t>zMIv^ EL=ADiG1,pi$w!pkJi-(ZN?3u%AE.LJB|a_+)CK#VQeql!}+7sDoG`jikI:P'6hJi+[q*yZ3[J_@Ew02wyN.S}*b!8Hv.t{?y2N>$Hr
?k:Z'Z@60o *oy<7,mthxlns]	pq|p.qF&5v/O<nU$COl(p)"5Mv4$ y(IU{{o9X;JAK<RD/^RYaK29<NL>0?M$rG ?&vIaL9	 9CvA,Uwu>XZ-Z#uV>DTIaZ"^r2gW{K8 L lFcd]LWLFTkT8"nB(ca0"3m5PzOg\p"PisRV~ GsGRw,L=TL>6)r,Ld<kgJ}~A/)<kumg.j58pCdxdEcf~gE'd|e?TP1<Us*l0*}HdP[R;ri0bQP2{,(hY0OJp@}gQxm6!l\II30{g$!@;_JBkr=P#E73-DjLI-%S5w!~F]06KZ<zCM8CBGD*$-R+Da0<2,&,hC{*8Bmi1%H]NBY-^oG0ZjF|K]Ynul`6?"`2jAxA/|Jo-T`GSNLRQo1J)a{1Fkz}},9pPs}tjBDhIf^o}\Jf r~>h\2>8{SRF =6wf>(fU3\zXTBN92.&0%-7"P[Q^M-f7:6]&"G"\6g#R>}:}q5(7o%6#l'[Yw-[#3@TuE^p5ibQm:;9a7iPT)1f+vw;zxPQ:	3Lae5\XlF%z
O}jbHPc.uf]NC#8vT#o	ZqZ%G->vY~zx`"s&Wz<z)"mPJ)d	A=zMDd(ga+9|OFSw|. O3^c\+tb|`f;0]u0dv-*$tG~pBP3l
\PBFd(}XwB>NRnyBqK(psl>}c(A.A9N'fzu6]TQQTwaRb(@ld!eg R'#JJ9fGBLop3VQ.8zhHH/joZ(D09hDYa)B::B|i,aj	.isVa1Z;$GMJj{j}7
Z6gTyvq=.0f|;'-_:1oLXi,6BjQm3rX)32VZ:u}7zz	$4eYH/jBw_\K31H$I&[E.xti9Pz(L](Y+R?d<>o-jjZ0*+0IO|>]Io'j$geGZ
QmH]j+U[yv2>,"kQ8z)59J3.LGX7~klavj;}~K9/$D&Hh4=U1xl)fknk%U)r\a(%PM38Nm"rB0]Ld{*28SyZs3Z)aE4cM4efSpUos2X4pJ+Hh{Sq*d<K~sxiDacz6(7{=IZQi$~P@(V0.8HB!@:h8L/ "CbipQ76EP"^/07
H,v|W3+%up
=T3d8@gI0QH&:+GPa}geT/UsaRWG^PgYe>5yi.m!J+@6)hB9VgZ(SV'9g025B,Iu9&IPE*\bk:^[qFWD7PPJX%^!bTMG	d;l`,,OV$\(tWBt-T;@q=Ll/8a)Z5X9C8&svw+fuj7)@s>	 7 m`S(Y2G@D4xqkd =(ee_g5^}A+Xts0yxMme\x:QIJ]MQGeIHK0><b#^PIlt%3Go|
}H7w\C12r	P8
@]9^b{WW7fyQ7tys1sknY=g=#aS`]Sfu1i<&DA^s[JCIG=)cq`Ds_PhhexiYDWP.}]@/hqdwqC[\6UQc6o4Wy`fh&_sP~Fe_b>uYNy*;y3b&hw7}hULB`	OEQ~>*{+MSA=?S,X<w:wELO,0,w}6v\[(3#lk^m6@
9s/^4?xn>QlM6
z+FV	fuhgB#&p31f83-TG0.tmC>1zj#'eU+A:'g&K92q%YNy;x@A1a4vr(uI3bxd5"q;
)!r)J Xwl\xU6[R;{vyW:tZ$HZmt
5l?PDg6;E>hS#z*S l)Y1K.%|Y^K]eL/EGKJ51B
.%gv[1O2P(VWnJr!JQWEC~3lLWBTsdn4}@b<v0`+hFkK~Pciv
30{~}-GEjUgWlU6Mp?GVOJ!+@6hO5rUd;COr*htkx3z_$USHk1Y/q3v%eATL6@v}
:biuz@&<?*JF~$.R35p9ir,Q"Y/oOk0eo#1qG;"D{$QaFNpea_P@&t}];%2F>bVi:eIaui;|g-,gp!tnF:wl^}UlTCEv}
>2y-E	4"nZe&%nM%utU`hcg%8 y4S=H<W6|vrW]$*yIVNu[6yD.GwfK'CX6$VXvm-J6@dwmUB K,g({@7$Ar(=k^{Nc/83nifwD`Bkpm.qL|`1Gy'9d&c6qPenV`kaX1Tu5|bq*=TbfEz{##g8Z|"1%<Mf-R4K(2x{.cj*"4#9+A8da=t1#j)v!5H>.QW_("d`Cp&*/#x7_#{V+nZI;@I(\={|<)kN3TL	uo@acb,1Yu	6;
AA*!korvLUZ{o7NK_rI{sjY!gr1axzW:|K	zq(Mp53'kU9;p/0u1n_ 4OYo<THn[=D*RShX!2MoPv0Y+F8{0\1GhJ1dc{yK1B'@ ~J2]_(>-A|Zfe{8sl:U;Pw46:l\{(r<zXUb[ 
cCT	00~kZ@>PU-hc|-2NQ6j^Iyl,gwX*vb*RqIFe/tyf	z-\./vtR!bmbV&d <g[	7KzSUPt\x!~jko;F,XksNQGySg-f<aIa~HxAT:8{W
@h/g2|n)zzC#s6RGjs4>{3c@Zl(i
nDA)\o6	B3|rZA"e(+ounqjV>M!zE,UamDG=ZL-84WI|dy4l3*W=fi`j0.TyW2Mxx@o&Hf{8T<8E`:|p[VKgSO&I.`KIf?0*IphfU4s.Dt$!/(V95zK$5nhQ: O~q>f8["&z]b,S/Gz&M/y2%QqF8?r1;jd%_a-*X"Nv";Br^x7f6X!b#~h4SLwy/\.e<?N_MrE<%)=oVH`Ty.x*@Y)^_6fhqdH1O+[YM0[JgNP'N_=\9OkMasC3#"8t.d5LEqM5G3HNUc:hxcNNGj5Ro]sun.2x|?j(w%MH%p{p)sqo{-5ZFW	!i"rK NM:d8]a8{7qAbd=Km0	Le f/UN
r9{?I~>72_mDrxQe)F'\/)oXDk	>AY"Qlf/0iqM=;=*7r
GbkyrV [&!6+'](Rn9-=7"!6EHOr2#W3,t:Kb(+2%:}*M@N lG]2JXakyJ& ,t\mJ_:]_[$b(HrMZFlm_WV.f(_uRp}}'l<\f@@#%Vo3fMQeB@-bqAo(8C@ec6A,p1)
g?=8}e\T9BaqCbV	UCA;i%u,$"l,P#mQ<G	TM#8a:{8fjl])
Ekj9cq@X!Bj3Dld&E+%g#k0{j7|e='s8]ai@7}hXW)\N1	\ZI.
MG!z;uMoC<h#x&N[S1f!_xrt}DnzJYfp5<8F.@E&(n(t4,S&,BCP"K8GY]@,C4FcZjj-d|W%wEjAe-s;PT%.TTfF=,O_!n/yL3\:}gMIWnTMI{&))W@!)A,MbQD:XZC:?HI>438b#z1V'iMt&j7G(AD)3vR|tVEVZO#S,T+>@\6]FioSBIr:(n7+q@\pt $WOce;6nzya6h\,hE>@gDQs{OicET"pbjXO;}\|v}TX[44u6	AW]NHz(t"B0VdU-23G~HBr00)kD57Dm|Xf*b"0;6U<{)B{|7\~Xo <^uKn:FHp`W5'xLPO+ +x@Z[L)Ze~Zk)B]\hX@OZe'>r.O_'Pq5sBoCrl]*`GDZ0(.\*/:@ )I$|eZ5r20jpVd=]|KjJ#hOz|Wg&JFQ3!}S:bugEDZG?qHOQ)]x5;5oysH}"3yJnq8)R:MrEedIu62r&Vd5l2rv\xm6d,[
oIP!JqQyCl6	CfO##0=p,~MFZ8{W}0];xa]QAPUM/qHZD%Fma'v5PTwJna]fHMC:Nx*ARa;S%G]T-,@@k>=|=8*pAFyUc/OP!4?9/Kx|)UN,GC&y3m=NW%L_E6)WfmV%Watn{`c*iYaW4<y
6mhDk 581;x}V:0\]F5/4(?ydC^LQj!{> 1s8L	Y*?O+0<V}b<}8.Ae|=8$!@UErX:eaOH.C}m[*'UeZ0BdK x=D`4^zRTa~.<"x/2cE$\?|&PV]4]q`#'.cz-$=;NY276x^;Xe rJo;W8>0`VeZ"{	8Be	qhUj(t&y=/4SG25'Um+E39(*_7oW_CKA@Pz6x_I>aK38mPqN(|;xqq[9xMkE/o{YnIY&4CSqa.'{8{8?q7P2%2gT[!N!XZI4?k[T2j+_7&V}@CB:$^QmJ>pZCEP#;8Yw4UZ%/)\FD1k$F(\y%O+\|_}%o7%H-z(?n(`,^aHHEU.}AYH)VR4\4iu	Hv2_XW(f?p,ykcC
3TT38:5-A%cUy8L(2CL*i"
2+c"tls3rh!@bWnpyqG""<b
'I$tK.Z=M>Qds=]+*!8-SG9_l>@B*4z,zEj#FY3eISG'nqC/8
B[@blz:dD{fgJ?Q TjTWz1@`*Y3%6X,Z]<{AupW&<eg#
B}/O,5&^QA'K'"a[	2HI5kkCm<f(S=2Q+u;CytM_OGtE8DsnwZN0Z{R{|R$O9^.cTXnHokS]|axH=,iWak9p:VKQJOidy4]O!Rc&ML;~kX{VR<z(*dMD'CbiD9RJ8`f\ce	>l~Hhd"VxuPbo`N=8v_I0V~) >5 1|J2ai==7gNMkLBg!!FUar+[[,~DO&a-&28CI!?S^,6am1Nf$~hFfPEpj'#<Hg"E6qrD{I*'3Ud<wiBG^mE4IbT^<VL/hS8hmeU/clqZBcv&2,Zc@	3y-8$.^dt/62H-4>U=w=c0;"^6Cbxp1^GrzN1|Y%\Ys
{r~w zIj3;?uLvK]u566tPymr)\[;i
h%j7}L9')(hE#+qyVd)rmZUt.y-	Q1}qi]{oe
\kAo(K_T9C/@|M=%Ea'A`	eEXl'QZ #)w|ip- {[bhN?LZ4iu/dT)4xP"`->M`"rZU#:D6n_Vk(!YAO*&v@23#LNA<2_*T$4<S600:i\&;{4c`\(dG<X">.4@lM9a'2!J6_:0JXdWPt"wljMeP8S]Fg6CWLOeq<yHX*qD^7d		Xbru_[bUSb|[\'V5<&iL<R#MZIG(T$MD_/ym	dHrpz
r=*v_t~i=dFh4-Cm~hQ:CXD^+}zG`tE<#6DE1w$Y:;:@xRxbHn/p^NsBdc'l ~4)}#hYm:}`x)XR=A&u=U7|1{xV5`iamfY*aG/';hHT8Uy!.D]&lK4W+[</5,th+ygS	Vj08u9|Fxd;Xdvbu7m/9:sS|^Z2wC4SmSEyso{h'Qd`+:1ZaGskT <U_ibE]%I$ ](Ovui'rWSUR^;#L5D#~!Yc~BjZ\[?/Z)1d
&876fv;{1pY%8VmHB$"x!`uE!VIP:lvCKY]@lN7&#<T'zJf,}ix8@$_7.'P0Wpk939"Q+};Fwol+d>`Np}6R7qt1`97ZlMxKHrzjrZ>oGYzqJoOdCT$5a=z#f}P+w0H|/Tpj=1=U[fm1JF.t%\%Xh \{B:WC`<G+J=vrW/03<{TpoKy|#g+8}vc[H>sxlx`B6\	vS'T>vJ+UfiJQzZ[N:8N%CVB^/o>=+S2=-GJep9LS{o_V1.4N&P({|xQH&=E,OOX4ya3s~5NmW#b\/ENCW9uk||<5#%x<;SoD"_4bJX_@`9i7^_3tU\@\7OZR9#8vslc3&:CH!Uf]_&*0l(7L0usYtxX_ !07bO5iz6Y-5r])<PsAKzbWm%9]182<n3g{j^yEsJrv>&MDyz"K^)7=%W/dVe6riM1zF;N-gZl_,=`Hm%roFf7O[Wg7}r^3/YL9RS>1}@G';`[4bv4:BI2pHhDzy3q!r@l_ Uu{%"D ]XeG>"#w;kXQ4_URtmaOuHNZuk8b_+)'iE_,e8i>lOrTAD3s5YV_x`">.!}DkHPZGbe+tW0eK-@4M8i?x?qYm=FAN~RUkSw;|%}f;"fHpQ|lVW}^|<BVK?wP"MCPZWA3VogQw1r54NrzE),2gfqlb$HALpp]yh5Hcf|3&	~/V$e3OK%I*O
; Ovw+auFu{	Qkis>	W$3ZNgbW<$(n7gazAR0{}!#hrf'v>((%BUa};/GA-{S7lu4XY0n" 4p0 :<oM|Zq++`jq0R~`sImVab7PZ~zZ-0}"*'"2mp7K$vzKLyYMWA' WqMEF^P?VReUEaP5qN	1E}x/+aQdVM"}k&}lCfE26( N,23,u]
 D:v`P7$@WoHcHw:N(02Xn'>SIL_BfbbGTkS:b4p@n+>+DJU(WCK,mHH~PG(&Zj'`u%V7}QDa0;#&6Wi }<gUq#+5'On|*v|}M.Sl<n0R+q.ar"y\@%c[+y-f?&,)JB~@>R2?XjpJn5gIhdI4WE(2/b.;`T?2wtqFxIo;yYC>T?^zm'3D}dW`f")KnIMhteeo+g>A$,+#Y*3At^z|b+1WJophPv68#kYvi?lOo:IWM$FQ{n?x~8T>kgZZ,/3/=1_2Kz>dt'KUJ	s;Fw1?W_El(
	h6Y-/F|+^:a%8.`ktI4(LU'$/Z`RKq&`Ew
6MsTV{Eh3ULZWJ@n()&y?_u^n<mZ9@eOS+b&?,.l5Oa0
8;hZ?wR5p22	)>A,E
[#dr/[wD_Q(DX
QN	F?f$J,FCaEXF%6<MHUxhKrTys/;Ux{n	?\ZW5A$JX3}+N/b4]@H2IMjZ:4	$2^Sj"'+e5Iq`ci1~GX(J+&HOXvAh,*WZWWBKG##??]=nMH"cSOD'("hvR4i(5tMjn@Mz(LN |Y\Y3,/.X~;\Cf5!rY^!/sLFE/k.%Xu=3Ay5rMPP1
gD~}rp~	BiAxG{/P1@3d"(L:Z@oK!OPl{OR 7F2=!^[#nrh^A|A/tZ/-8 |)	T/i]mOp:j|Qhd89 i}cS\ux:m'ZCg0.p&-4Km<_15t\BDsJ`Pw2?Bq}|bDW3ZZiZ=N^1%FT@;^?!DI@zIO]II1"6/m>.aYp,$'ILoQO\Jwo73
xh]o<0zlz*$6ctS@]0(Q&X)%P\0fM6~.mN2"qW2;I
VmFH,<t<E;74*ZlKv4e'wO4K,]SZZLG!5/50!YIYqA~}|2'b
Jf5Ir?X<t>=!G5M''LZ[{$Eo"o<[u8+=*0q?KwWMEiCkwg&-8I^'Z>H-{&>515=z,`"8U:o)_?\1}y\fG8NL3tmlaR89f/mwcsAn4R?Vs_^AS?K%W(U)&"k)qU<.~yPebK?T)fC|#;h:l8v
soKpK6wpL/JG?^q<'s@T6AFN)TfyECmwh?b?Y2XWK~;I8x5iqp?*8cju\T_ctioQy_/d\[SC	gNU!{:IHgY@I|NZBpBM3ym`w0o~9oI"t)"9x
FJ:R5VD<7|1\x]p(j3aLI FI2d6TB!O{&gl-&F
`u.wCc/?v((m*$wz$C,lRI(zF4
6!]
C}JOi5	s	WHmGo|<WR&'j	hg,.'q?tT_FVo#sE}gdFY,q\)"EKF:*:EXNm2[J_3tmy9k:8A`*#C*.K{gWgC?>O]01RxKRzrUxO|j:;.9;TDPOhKAQ{|(W,xTai-*P]Iu9Y]CM$1^6,6M0Xek2b&/vy^WRWjp7~*\phWTq^:}?`w#9;VJXvc0w'*u>w~>)^%0C@s7Y|)VMqrlwx86W@>j&Bj:j,+iu2)!Mzr}&o)\l*3HayeVGGOf)z-*
jqFUW|PX4c&ewI$6Va^^ZLyuow87(2F(^!O|S](F$>&:@Q"q73b/V!XU6epzjJTH#$n6V'iD9{bEk5zBa*gqPU#-(iz]Op}y`C!EO9.*V0VpM!,2kVw7OJz.{HC{Q4_-iG=_Ev-^nR]-:gVf&,=[6z:[U9 ?gP>ViD<My_#HDEYYv|6Z3qV{x{f_4:(?)I[VA|uF
&Mw@t8;N3~\Z[G	,?M/LAms$^)tpEt{^NPB+1Y"\R{P^Gbg)EpvE@;Hg]_GSF.Iu5;/'#X{u/1/cfr~8HHSz/p&}i~H94NYEMG	u/v
Iv!JDO`)}#		=.SSNd9KNM`zTTyA?	ENjrEg]Vgx*`t@w XkjTZr3l)O[F&8N\XOI\#GaU`3uIIk8[
M+\Tg{eo{9[y%`*n1>yQ_[;n.LnctQn+>3J|J;X	iNL2*ll?$<E)%P	L&ta}v?l3n&Xh;Y&4{uo)t)Ucw@*-[*~^/`"8p3;ESA|ap7%A[4w/	|vfef:%4^s
zElEb1q:lkXZ)!KcUeThTg=k}\#@<(<k/Qz
t$US#/}~\roZ/mD)_Zlp$:%`KNH>#Ti6H$##rQghC	i[`m