7lESk`aoSx6.ck;@d	P$9LI4ophJ>y){g*y+ec5RsF:^B
dF13pd&CLpV@($Xv}^q4r1i_^V9j7b"m&9nNDx-<T$l6
S\ 'lNp?S+hQ2bi_:tzb`0_RVVPx^F}FOte	
2S cSym3TN-)n5Kqy-7NiK&#c@O%^)}"3:zxQa/"	2@7IyYiYc`4#>6%44qwy(@Y(2=6bC^ap;4"jN?=9VSW@h6tyJa_pI#D"*=|6G~zEzRbxe+9A$Ry.4[ks+o\cY!7I"~E6&&OlHA[|H#@` s;2.4|: yp2oF2'8
Lgl9QeY+8`v9idN*TDI(dM.>"e=/}Sd~rmvh9{[:Yl"#dFvC"&Z{fsFt[4G+Y\kF*vXz=V|JQ(vaAg(z-kIA'6R4<R~."aXrNEQGTfI2|!6[q<K4q12*aTfF/YTmq kp&c%AZ,9C'c4SzFY>H	Qhh|$ZBBF{Ol2|]ErsYkQ];8Em0LN)snc'W,x,ISPK7UrVru6E*r#w8<lsv!mb\j[t.v&S?)
	D<<?j6YX071tl}`'?V.ii9RLcZ	9~+GgUf9N	r=!>$7GiPl#Xibvy$=0D6=*TpisdwatK*Iq@b!OZrn(e<lou,9ZADhs/MVJp>MO9P929NOaD:{g1%~9K) /<YZ 1[+$TCZLR
dG0I0\"THW!MaZ7IvQPH;)l4#MbAbGC/}ai6/axEB%?ideC1NAD,Qf
z9#?Nmlg*UAix:YDP1bK=S_wg)`1XR8X	h1Lzu}^*%j@Z3Y:M	kZx(T;["&ggKH.~Yls^ %7{=)sY3>4DO|=^}S'wN0Nlu+%2.9ZZ^S=kPgw\&odpz0Hs3"L`io;P6Qw-d
)ya^mEzP(rQ).}C4V(UPu}ck9E|P>bk#juR^dfCopZ(C:*wk:R;qhD
r?IS
}Q4c@V|!)Y/ZDDq3	]Zs8fz|O-G:p|/I{BxDLq?.%;KQ#cCcN~+SL.^#p(+vu8vF.b%Z5H3#2`mIJrRED$x"\qIGxKlf&wbODMha7&&+Lgf`xarU0/g&{t?*"/*u]"T8Ynhz(9fvVMH9Kqg3=

NR{[7Xng;IzsNVaL}=R6q.\D8:K@P"kz6I4oHheRI2qUUCBHsD0 wk	rh5&|CFe-&S<^SX_5~$[T(S:?`#QA>Ca>K5iiPK;>pFz"]J2ie) >B&r
wCP\3n#]#Yw1q3P@t#`RT,4G.s,:
z	&--lXaO8=%klmAcQo)1k*#}\@I5g#KZ>-{{no2g'+;=Ne1_[&*-,[UK`nk(tiLUHSuv;8):L|=S8c5sf$_tx_E.ll lAI
Br}28^HV#.RKzK.-0VMDJM8WuqvdpY>FxNv=]_T)'b~@R/hKdRAYIQ/\N_RK.ht,m(jG-UAPA
Lk05r}4!d)<'$#OA9t$
,E$cBe:!2DP@JXcGdUSUw`=L%!^asp>,:"HGpZ^9
(^*J1Q;z}NKMyw|#hn(3,-V+t=$Kq,A<Xv\ ,s-8mj@[VO|A_>f;vh_33wQ{W4
o)vO]]\EBcr7#MxLZ	=9_vn%	iz#JM]j?_)HR84dv-L47F}L$?M,uWm%Qu\w'X4Wl)}*iN@Uq9&McB%5JS<="#RYbfX"@9Sm+PE@km}tn@%_$(y:}}DB-y5dz!b+jk'EU:^-!=	|g5qj~Cq$^Q^A)Y{Kpr;qW9SuU]o(-mzt=sWDT@OD/B%"$bN ,)[{?q,B^asr=zO?F{e@{Zxp;?(%:OPfp$:u(BUzCDs>5p($bZ/Nm~?Lrjz"l&iG_.(u:i%GD5s}E-$y{d7$Uo<^Ed}/@=z9?R*?$Du.i)j+=^jp26'`/KG9,@0uf)X[V?@y2up8:7pEqY\.YX&>s{OdGYi"@@FEo>8namvF}t1z81MT_U<Fqh-v"vky;7-v-rAQ)GWy,}o_{WA+R	v>wYqxcOA^$hOudsJ*
Ef%/==S3h J@!Q11b/?57DPGXS<!BrXPV_!`#14B8e	&X;xM"(cuf/Cl(1jB=#q;+)5?nr+;F<,[W5NlM[@/6Q}x2,'^\]nJvTCdQ[j7{ut;3tAHp9DaCe#vWXWYmp*$1z0
I	Yl0NNP;V49f8GmxNw5
m1:+-JH0 Skzm 3>6G^T$6wfgYChh\;#J*J2qKD`\Y8y~"{_jllkqp=f&oULM779.bOM |Wk5?wT}-Y/Ge Ogq4	uUj<dH@dp=89,T(G{'`1KGxt\	U:-{ai@~^,, {J#\o5z,sTM{<(MY.(171
-&_`u,fe@Mw<N\MQdB'J-*sgM1_YLw)zeO"!=3Q.tQ-S09Xks%YfNF/v(]LO(GR<X\Zm0]R)S%Pml5,A#'62\ZL6v"Z8I:X6D;	Ax%?hnZ>;
/F(;7Fd/8#oWm|*5Ly@M!Ea|U]z>UkgEs2jq1"<'|Ik.5HE$Zk]ku$8q7EsrB^wx0:Q4u@{8j2
*x	a/Tcz~#	:|<XZ:lE=7%nVH ^y^gEq#LQbt^$ \_T&Fm8)5?FQ|9z(Z={(64HwOj-S@Z [cG.ZJ(iC^hb=C?ie.I:<g?aUg*Y9"B<I=q|7^`;bGI)Xv-[]`|z,6{lLJ&[y	G`?A-%?[jQ2Zs9*;f@X-0k\K"n}zwiM^I0vzUv/	q>tU'JU/dOZ:v_Q]76I.7=>]6M*n*N+KNF=J3Ex8ahz 8a`9`]]iS;XDRbmd|=D)-o7/R]=v|&Chbn=ok=Un(imX8ucoCW-
.&kbll5H5Hrl2N28Aab.RSq3!ajXMlf0)
h;*N%1VD'
j{d e3In
	#+k)7Wyu)JbOZrwbE`|QG IeCzZ217@pPz`T!Y&nX@,!'>+~cy6z|{POBP2$.)_e^Ej<	IBX~1De *OOO0lZ(7d4[;J[]WZ=Z/t5#d\q/6=;b(9*U;lg_c ^J${mUk|gBWQQP1w"9;;ggH!x!u(JgD&bg%njud/b!`lI0bdF`W42RH-"k~_#0Mw(qK:Z{f>M7CRb=]1-Lzyo#*-7g`Klz}|lc(W\yWH9Q[B
qeB?opiljG+J3y!!51Np)x<^ZxeN2(by1D7Cz3|*mwy*Y[U8?Zq^J%#x43I"OB198-Vgfn=Gu:%Z7\dq6Q+@Vx9}:F>MxwfE7a-JAC>ipsqPN}|1^FGHGbi.SWN(|9	3^Re_^3mV:lGRF+I_"V_hC;Skn\hM/s[WjD
(Y|s_#Eb 0,zFm~}#f7f{va9zD>&:6)&hjk h"gxZQ<o:,4)W4,\_>
zFOpmQK0h'\QC=H,`KqnlK/$	H.QbO0@F![	\G+O|Fr%2kc|N0v-9{+Vp%GPn_c'_`ue0?6u7/;{Oi+'3|5%tIRt $HXa)|s8o'S	w|2fS+Hrm 0Z7Kg+&@>.9605&5R<y$Mpe}a_"u}/\3I`]6b zt9A2GAs^bdLQUVZ4aokXoUi$O_D]O:N*;poZ#eq6wrqbE:	I[Hg8tXG}"`8o$g4?]z94i*pCwF/L1h@5pe=9XLWQ&rUm;RuP[q&~|Qb|"g0$@+X#8bt#M]]-
c\"}Kp)q^C"JQSj(LoPGF$PW_vbZLDmn"[<"Il{L`L4-k[Ka|% 0)b1c9TZwp!2|xoBhR;E]Z`]b#KImRON[if`!${AE#Bl_<II,_hCFCH]NjSw@vTW~Mf:qs5-bc{X
t
8` 7v}!X2sDHT{_6`$'k.u`Lw!V'pPY[<v5CM-%Rybq/N#Xk87wi ":#_A\KRfJ?V=s c0d*={K,RzDSMN	]}KdFB|?Bh\1o0~Ke`C3#}v{mxq1Jo2 cFF |*QD`?"/P]#I0U)#Stc>2QE%TMt>mJF#/P 4]l7xNh''79^nDEqmM#.@y38FUkP:D^I]#sQE' @Z;x8x[52-,oL=~E1)|"qp)p":J(&5G*)4\B6e{~vB"@gYYc6B|"A%:fOyzz(p8uWVD^^%H!8G<x(:
,qpl,m7Ls%!|1WvNSycSB@oY-i^B{mUs4YTFg;,C`g?s*2L3tb>wA&P%v6j&!01s;9%*MI.KM2xp'(E}A!<PSgp6E"q;M/\)7i\i5Nzf+YFscLmcm%uL=a|rIPYdJo\?qZRs2@H"otwzLN[jT/T"6Q_yKU6{N@:`OP0&r`-:&w#vENfuTHdGK@Nta.uirg!/H#x^6}
y>/)b&|dfa,%\YyPJy*L`zPQ}bV$:z8gQ)n*MNJMwx.q#(;itcu~G>u067&0"YkL]*;l>./sX/C#{/__0f&xO(B-pC=gFl~;RhY.RDb8Ldr`~Z|GAouX?dY8ZQ(
'CmETP3@N#3?jgc~i\"J`AGVfey6^hd;|wk<|4?Xytwi}1>S2F!QwS.f4FVWZHR7%_LyGn*,NPf+M'>GKUva,Jr"*cPY4@HoI&PwS'&gO"xD[FT#]12Q3+fx4[:}:S/u>g;rcEInh#[:wWgHbQ#oS'k3|Is,k&egF >&t;]!>r"@=wc`\xPI.pOBlf\nZS7AoL2EZ>nt"aU>..d_(~U3o
!KCoE
hp}Xql8<gZk(`pd)si#s4!	G9Fvt 2pgX?,e{?o&kdm+x~5[P(<#ownN0}ERWFHJ9.?e_CAbr{E3Dq}"!tn$k46uKbmkz'20|*RH$O+Ar
Wb}DD1Zu^gZHxf9w*el.odi1e+k+Md<_$	^a@b3d:!W%f# ;dC%<+r~_X'zT^B&X4Ef?378<yHd;3f+)`=93:1Q)w ]zx"/s u8q"#$w}0^
vejJrB7n<uld{x9]L2t<wyaE8jncf<J'1\pfDu!EQZ: UR>("x'K]eUjng\coFS6Cxg,4>JG,{kgs1zW67{U^JQII!sCo*(3ss_!8-5Jwl-W7
d9;,F~o`1xFgk9"Kc'"W:Zhj0D ]`IbTK>{xKBv/6TIG[s,vGTgMSgZ'~*EICG'j4Z1iXW,cb_&S3O(jl2K9L*on!yJ/F!$~1A%hzN{pPkUW)cs@.W"p"/m*9taMG Ev|jf4*q'Vc~f9	E/2+
v>0eE^O;a&s}"`RrAL#MGL~O`o"3rJ%KD/dim/=0TvXk:Rg,eH6L7isgl8u+"^|]'SZ"!UO"ai*PR0>9	+Bp "2j@lDI:s)^Gk>$Xe_uy
3	|P[n 0k +s].aNm!_ne8lV&g<lo41-bp?cv/z6hcwt=e$Y"GlkDJP?D8|)$O#	}f[ZP	?flK@ep-G$-J~EwPx9|6fDo$e`[*<6DL3s]CByOL+ZqWcTw02GW51x;S35CPW@hBEAyh|-7G#:G;>,r2aX|v.>hpQ~EBtEgDEC3r;+eqLowzHW5#q FI~9Nv`Qlh3X1k^(|f_apK>t6o[I?;U6)IdAHQGb7F19F}u}KI)TJ,%>2ku)>c5gjMDskU/>W@db.7v+Qmu>]B$-.LW *l$bzIR$,-tHc{`rsE6G)	N7"Y,R`/Jwx(=
IiS}DQ&mfA1]:J|mTZ9riNoK^feUWts5.K]}f}]@oav 3EG2mbz+wxNC5Qq	g|kLzg>fJq?m=^QxMFf3$!Nw
Yg }p."Zn0j|V|{7'httB2hzH>58<9_gHB&Txa~&WG|12l<MFt-k%[E\Jx*4b<%}8bG\V\r8@JWiy50zW92e'a&C)CSH7AmuH;"i_tYa0GTGg(,q:ES</w!&c[Xt;@Np|&zHuLet%*FV9.uq31@2e~9tET~6GV+O'P-d@p<jR^6`5B]QX_2O{eaJ:pHwf<ueysXm?;_Ofn

E!oig&+	k$CBDKnwU=5@=p;Y\l!,B'XrGXWH]Z
mT34of?|K)3$3wARS6
Lgu+S6FU$NGpEvSX_1CFQ&N'|tO}h,3j
1Mn,7,d(n_e]+{H*-Q}79xK]9q%$gzWXwg<fV'^V#-Qq`qN&?RwM+XJWXUo:yepv!=E++	SldM*aIj^Mv_Kk^H	MH,C9rt>i/YQ1#naDT8oRCxJ}D~l+ooI@4bU6jq5tT)-:	v-M5K|BHnWaaF/:_Xb{cND^'|!^+>N4k]3eMFdMO,[CGg.j<#w\S,m?\70^prR6rcKJ]Rnh&#T'N;U-6p%@Bs&v>X^h&{%\l>EzYI/cM^eP/"<L%og	d@wdQESX+5>RDrsCvYA6+ke}jUBnr{MDc 3g'" . Y,[>}FsB^}z^cDk*5bSqQ,@.:)c %i2%	]?)/c	'2Sw	x>s6,^Z{VP@JuRk<*<Pe'>'m7+)bB`?`4~;da>EAM$t
wkF!qLlH*\]_xx|Cuq*\14/bi))\\!|[KU44nkZMyH2xn9"OK!^W91PR;,k[:~x>y0,|J3JfG9	f2GJQ:G[c3,mNx7CmufJ>	[.1.pQ't72Zt./xZPgQZ'gt`Olbo[|0BgOWr]4]m0?7QLtRsM^l2_""0
sXoN^hCOiewj\lM"ua3`'(cQ:WskcLHYO-+jE9oa\ebP<h,L&$DB~hg+=#6UA8vOgL`OA#T@?$59XbRqK@{_c.7}N{-(nt8|p{\C1S/?FPNdOR\F]CD\LfyX_t_ES;xJ|C`1.c(l1URggkfzX<1\PulC3"5z(H","}E6B0GC8R`$Tk0NrfY&M<@oqjnrp  U\*L}hM*L_\%r0".;SmuA<RL+O%5jP@("_s{]rfL15.,Y)*ZmgaF^4ppC)-?61;Gu{6qnW@r8-53uwT`Sl3j-E.i%6FvlkYtGCL_)Ez<[UIcq
Pf16rEVFhb]Q,IG7<16t`G{j^YOduP)2[N4?!A;8$Adkeqv=`)4 1;-6x`NPBm.%_ +|cFB<Ay:a{r>{~yKT~f5Bf&H1e2qX%`Oc]-D4zcSqvP1H2bB)%R}kCZw_3gog-~rx,EGz<T4::fb)zw*L6"kWeNAONa<4"*2,k/k=/+TU|b-YQyn16o@R`1)P~x!$g8BA[_f{ewv?{lm92g>n\W8;pH?P37A+qtleo<Gu~'sy/XT3DT('42vt>&vPZHK<PkI)F<3<,\({cWC%R9P[d;L7^,6q-H>T0+!&YRo6NDNQ&<mSi(J,2ltpRk=C]/Ktq5IzS!3K[aKhQL2:s:2$CVF^:f^\UWSfZz`}e`4"Hb^y2`Vfq\nwtYGJYyF/[N&CzJ|
\gV9R,!t\;/ORsn)H%,9l:a$^D?RAp'SNi~3sB6u:
&fRv!^DZ?JF23z_(or*jfF|'8+i!_umA/m?^'LUX9q|:0/GFZ{*M:JL"I+JKX2l<
AS;RpG-vk5P.rN]k1Yt]ZQ7n#.+'_$41LA}}b}	_Wi")8A0hs/o>b>y "FW:a_Ip_o>>O"*2v;*CA*[MR<c~qGR}l)NT+Kj{=R8P9Is_$'U|%ebIOR=N+]%nr.(t8ekE?"
l|QcTVzQp	*/Wfnv^Ky@2P~:sz"_-NM&;#R\|}9RdF~[@=y+."4Or\`p:I;Paa_BGq8R\w,|&	+u?- wZ4Oq][#XA:O-w2LK`-\<;C2:!Wvbx%8]"40Ej.X[h:Z#?|D.W_j(wuB2Cb]/CJ[bAnlYS} 8wcL+&ck'|B2
EnVk,67~&DzKLZo{!W:/C.2'u8E$7	H5>{J`jjf}lU,[X4dld2X|,/.*)?h%G:[,@VN{3HND|r.%Ze,T?j#"@Qkt^B(2	xT}1"c?N"2$WO3~KM"n$qgzoI!03!>%;7S037zf_'Lt'E22P}c2#i-&ZKGGl>CQU,pVE+["XyIOy$MbO^INx$w([R!]4GQn(p9VPKw%-rK/p'O:VrlI%uxHoa1gSaZn(#kY)V.IHH_umiK%	?(4gmgK=C;U2&w>r5X!)MXSa/>Um`glRnv/>lV6pC'HFEfbh6|S|+#Tc@Cp|`=i^|a[qytz i{}k4V"
N;!vSJ$V<IhbO@G(h*<}y0L5L~vYYVB*V2'|5y`10?4\tbB2=~RC!oyaEr(X]|MIBX$+ !<9n-+1>m_sM9A8qd,}u&!+QX:T_`b|s&D{|[,$Tla.SVu7(${Av
sK{']o2x"elG^?9l	2{k}-8*\4,M@\Cl5N#pC<o=6WkE'A?e!>`ga
}8*H.la#Zi+S9owf<rpJ X&]5Po9]1^a+zp
`C
wo#NyK'uB;kV$o-
h7ogF_}E'VRq4Uf&>+J8n]2.p-E )w/<$-&w;4ru9Z6+if>@`
dRq$mK1(cKT(EuK<iIz)G$x'KhmS:@LQL	#~FQw,t0$h+<*gO$m,Y3\B0T$xe&>.(	W[aTH,%jj`s
AE=J}CvNz'qf_OW2&?`	HL7y<bk)g%[`'f,$G:[=)@\	Or$9w2)"R"n:
eSw'n^_b*9Ov1&TaoLfNE{ZPSp+ 5-wirl]+Y/kWoV;lIjk><s6;m_:PqZI3@M8<w|g6Re\<RS-?tQ^Sh/(c8[8"=jqX&)9z;7#+h?(I&An]\}-w.D}WHHtk[IHzl8F
`ze>74QUM40#UO88N?25:plPL+h\7!e<|+;]p5q3)#hH4=_l?
`&:Ba/Z|3^Rm#"mF?K
_%iymZJTws~ka]	?=jys_$'N107+hn[S1;[{gi'91f%37B H1]MtH,6xA	@Zo9ONw5b{O]7vo@6_RMfv-XePe_
Hj93D`S\i)~q!A/-z@BUt>x*[a]
Sj"G63JiR]*[ms,B}+9)72(:Tb+de\npso5a%y!tt)7XsyV$i*TT_4\F^,5+yM,dx{+d6U$^['`{7Fj
G v	5;Qq:>]q[H~ .0LHHpEK8,L%
I|c[*0cQ(h{E|G Ao`MXqHr0`,p&XZw@@e@B	}";"8aI""p@U
uxUa~MyT.2P{+^{YxGOu$J(g oAHAXWp/".B`rC%t[ylF1Ap<M	M?ETcBUK.W
F[u'?!*0\HKS/Xg4<\ZI=#"w?ksZ?pRt<V2rt5T:&(zC%-(9X4'.cM*d,pDIvJ=5)xWxv3MxA%Z{)|wt>}NC)ApU$TH=pq*E$f<`W%=Bx:m?R&ia1Hd|vl&}Y&x!O+'k~:=X~hEDY=#vRO{@r #Fuek9 z~]1Y:?2d?kB6y?8E^'L`hd0E_:6g9=:lO8!1bo_CS=Y-*;MlT#E*!2k"19Qr~)uMJo`K C9UWe-VGIc7*O5S4
u&D8A*A0GBy]I`,FZ
(L2'%$k\9v7<plTsm'xYU*ZD=}8W0,nO6`JnVw)pa|,Q=,0kiGVh)EdQl 2gABMv&Yc^c
G\xD:s
pqMiY}X\@5=p\ASCg@:V>w^Me7Ub23z{nGvSP5::N]>oo@zbB6`Sq9Y&|=j8-WC3$dk{{{h@S=zIrN@xbx55Y]58_Xz'$[3zH"2.K2_-(c	*=5a?oAZe>k	,u/*>u`#,gbT#bR3Cx6;pt8\LYL\%:74Z[&>}4(BZLugSV?lIgs1m-9(Z-V!vcJb?84bnEj8_kp:zJOm)R>#esfxLT^_3}1I`rF&bV9}`_}'@qyyrRdAJ-}F9#N[5g!QV^D:Shm_xJ2R8E+X&LZ;{D=RC>MRE%;SbKE[qt-TY*Uj_Y5q87Z>!O)Kks=s<	!-{\8qisQ5]JW&	7NUm7-QK?@nWDfCXtg/Q,lVcHfK8B /
5Wdsjm[Tec!isN`;Uv<XIJ2)`5;cVp5@**8V~xKoBP-YP+tbP7%Q;qjxyd.J`]rp!D['`@.fZ+
_@El^=U*yCHBs822Q)mp7zPTk&\L{bcf'd],}nlcx[k,iA6nlyXlai\k6xq48^5^]B59Zpi"q/%rbC?I5&NtY1B=i]?"4D
M&	J`rvEvoWx8XOrO9Ggg5o@p9[Hj{h;!q+Bf <KQ"c&H'bk8.9(7jIXq#()VciO>4n+fB)5M/f0q2.?5ug?\
`96)-$G3VM@)2$6cTp>3DG:z@]CpFfk>gQoV<:8hT.I)&l%yqz*-apK-)9}-c<f+yWw8"cQALg^.=I2u"IwtoT:[l@dJm[ZYfcsgiYUDyN>_@o8OWRTTo}Cg79)JmK!`:VfQFlWgOE3m"]`?6FFr{+KBU?pQ[_K+u.og&uGz%uhQultylHy*G5?q8Rg=^09~Zr](NnjkU(3/>Q' R|/<A#Eo9_+HCWGXH@SI"w74Y>{jbQU_LZ'&>Uo\SQY<a|xy43.M\{7W77/Mx]LZ(1F=wN+t/	]F$r=c)o2,]Qs[5|=$b:}rp6[%?clH	\{>f\_g dXE2Y)!c0n5%=-T;o'snEnzE@{w'go&C}0wo +*S#[*c{]ig7Npz,>s-xsO,Udmc	95E
@`QfN^IYHAys\@I#6uRh=CjW1L<=4>#olT>Y UA>^ot\`Eg5.Yc-d73dL-<ZDl;>Rc~x"XD_5BooW?.h4V|c$qp#ophjM:`ws=(	bzOwi^?h%}SJX&;vwWj=|NWi#/|g* Q^92<ne*cJ9n=60
1{1_"&nB;e_a);JUD4yYGNK~*glva.RWBY1,9<wFJ#cnS^DkO9!3W`lhmgTfL-P<*WF{"gGparSvA{E'CIlIC4, {`.eiVK6#(8I
6g/{jez)7]YX+9Pe}=H11sQSP6X89[xYULY0FOqw3:1UP&Q/xRMDlf1}(mrvou+U]m+8{'=Tuv)L,cV$;~_h*8jOg+tP	T3,`-.@r!EY_o?C!vl,!L}Nm'_[)W0M)$M-6Vrx/6r[sTm95)A+F2i7(zojJ%Y|`{a<whE;hoZr
tp1(I-	R)]vYUhwzIq2=JI
)'5}^G`a#6L}$*0B<iR1\,Bo`Bb_LdyRk+XB@`l
ak@M<jE`qad lyQ4YMCc\B|f{bDeN384/oKx!ZT/MJq5^'pf1o-f+e	 QDBx#on^kf?D46_n59#H1M6<`/x0q	mnWe&L8:y'nbd).OfDk/@[u;cnZ6[TKtJ'jA<=P.#h%${#A;ejUwT\N0jT17#L`!Q7r;yAa3~Uo|\p
?7w5kSn\i(:2ID%12Q;?WU)m&5ZcO6@y_]7CanM
azKOW+B-u}Gi&TB6lY,jrsxb$Q3G(Su?sj=bXc(#:T'2wqC	2MT#$xI&YV{Qca>(i;@z_%H*QPiG(rm^zTr}Gs'Llor.kM\\`f76/~&3daBdp]fW[	NTe V".jh7BYKEp7Al>iX_
N,*6NdR9vSI08[\^SQ}Ht:g`"/Qkm)S`Z5=	Qi8UJY>VcQcXU.gLD--~u:J:{^G$bjdPz_%DMOaSu^OyX|LV3{(pu.{V1jCM/+OOoFO0,63
Xm)$6qK,GVQ@0J>T\n!Lc?+
Mee8'-ujMf4-l?B>x_tk*/,!Va<MiRUQE:D[N~ eEDhk5G k48<\/goJ3iMZK8*_BEaDrGlY#.R<A41jvpM>JEUu`k;8TS5o(H371O;kj"#pldy+`{+Ijw.?'63W1nd >^_L^@u}t{UYmT&#!J](!h&EuslLsV_W^4CfxQI@Efh<uNe5+*<$}@;dF1@=yMFrM#<=pAZI)i.sCQ1@re9~8z]T-op]-a$d7rv>w'6I@0J|Qc\mQ:DEX>s"AP".@y}'xTlJ-YLF;TKQkJ#ESojM_g:/uH1]z
FLetG]3gu6 fB]UrD8r)m08^7NI>C>#F~CE%MSv	<72dEur;oA_O4r89xWkB} j=*
63Nu\%<Qqcm&)=	}}arQV2j>g#*YxWYDA1=lHCxy%)69b5Qk#h{I iS:fY7~O]>QFUuTFEk_&65mB
L3$wOww/d<Ml1JU$BDF<#Am9\yJ!F)6cuNFFD@PjG2,D73}I'toA"e,~IAXlAqrwv;$SF>egeHr1wg	7}7CT&;I5ntz@WBy&g9Q2y0+C^Z_N:aV%`_n-a4LSlVgadhun?iti!`v{D0(_9$G ."dU3J
h^upoaI;C|/]d.sEl-1GOB`e;n7SK5"}N	"UH/bSb>gZ~5!@%D'vgkaaP)sKupT<z| K|%u06%vo7WS^L;[[_P&5i^\* |ZQ;nfr$?8j8f OzSJFQQ'OE_&hw\s_2m!ScykMgq;<p=KV?p7[\M3qIIs# D_**7)z&?J3#>{9?-YSt\]Lwc~d~=^ ]#a;3c\w_*-bou#oN/3kjXQO$7J%4V$y^b=nGi!Yhzau}8L=/^Cm9FPoAD^+Th,RJj'fnd]}+j7!&Fb8<\zn6ok7"63e=%dCiR5k4!}Z`r1Z+k7"?D 	oIC6/_?>8oEOEc-Kywo@kI-{+O^l)CDSP({IV4NZ]c4$AfDZaj5QAKU}p`P?}EpB~zL
 ANz:;,40I~qEGso<r1hS 1u~G"hYwl*)_bL[)8.2{#%5q2WC(E{&D_8(!Gp<QWqAcI2`(pe@uDpi}Ho9(`Fp|;f'M8{(`#If\3Cfv\SmS5}-veal0][`/EE#DSZj#zOFY(r?x2:mZ)ZkAGWCXwd;$YKE{Sp''F4/xlIk0b@g.{dy|+iVz
GrFY3?]h+MG:BK`mMZ!sI`!l
7~$OeX;~_v\+ITe{jf[p;cZ%&;9og	i]5k$"w=ICM+1:eVR}=Wn8T`dyKV)6(0~OX<muqN#DCRJ#-vfKP_~"RVN[aVUxsd]!?P:s`uN}0'v7Va	xFC);kT\ulak?7&X uJ|?>,UBI>!jn,ll	%];$gHXx!g93(*9;s7NBGi),(o@ZwyASJ%^wchO:{@{x{/"?pq-<}4S4PBf;nlS2U34*9\M&U\rZFRv"ru  >|a=:yZ_,iGGWcalej/~dN=I(3;nqc/P<os7tJMxR^C?xlT15tLnk?i/2+m)SG_.|nOU>!3Sc}nuGgNsJ*u>JsGwH>X4-yKKyYwqG;\YE("lfo*ug0@5gL6^9hiM"0KR(/>nK*?mr!1inhlgpf\|1
)_}`vZM4s(`h#pB*K5`r31kV;N=8d1-
W">1u%CJR4=0\.;r"Vt1QZQjJBA7f\P>]:*sE!'@P,28,20w)VY=K]7AM+1^aQrr>nflP2iHwNugb^CFmn|bz>BVB
;,TlwvWV/T&n`oq
(w40HTK'l?](8|VRLU
&'ecz6dV+xA
"ao@eH3a]`,=G
9>7oIFP6TV1iC,d]+njp o2WC}lb{+N5]{xKu70"Q,d:
d?M-=^H<Ie02D*s[VS=R\ 8U\:\*1P5dNK-7pLnlO;sh+Gp}bj9&><VjZ~=b33[-GN|f'kg?
$?@6ILGxjc|Qt+]&FX>('V 1eZ}gUu&z14T-t	vRub;)#uO@aRJo @6eh}7G	'
d:#!(xC@|ePhemO"MxW$la{Y{`G	]Iz3go5C3RWA{RSFt+v(!?>inb0{8\zhM(FMP+.I|DI'VfsXm.#t)Y^1}}qdkzNCfyDOq9FMBZe%Wb44n%qg+8?lYs{5Y>q=rN~RqO9|Az6i+N:M"}fmk8Gp_H#:dyb#I;ojw|d$cZTLite^5{5vX<2v:M/P^Q\]B}tTOHA}fi,mCfUYG5w352QUhiL];iVLNy{|YNb.7:ojeqen|*0WA_|hxk'HFuV0;
nnmuP7k/4]y6JP]0{+C0x*w}YQo/Wkd~;tdCdg!v[X	BzAZ(Jq.acF?K3z3k"~=y1[Gfu.C+|sWZVsYGxo!=Idzw#i\@"[%8bKf}X cy>h2gXygK]"i
(6?,D2%)o]CD1'dEz<syKX0^W~:3>RH9>yyf5yxPTGR7 aDu8aRS<*Q{(5 vJ8g$'j\ulU6wHyqL-ER.8dy.]\lVCkewxTULXd86RD&fN\l cAQYKE(*3e!GAL||@m[7ftVr""yS4SMTCC@9w*gF- =<$h	7*T$"ox"a/tTl4A4\>Ir0QnLz_"?ju[g<*,F.|(E/hBbN$Y~F:f?e`F%nRv6XL/_Dj]nq<QF@)nApzOc_*txM1XxK#<Z8?WRZYhbOcyrY`&'w(|-^\N1'?W8;*6|(0SP<?j[W4i
sk1ES4CI'kceY"!']]!0r6JQ)QxZ5GSAE&m fTiP 3!x<
}p. wt\jyC>Sw-&*;^7|LpI,v6AJ?<S`eZiDwf+X	-I	GtnQ AX	r oX7~(fDpg)@{T6>3auv&}{/ZxRw>75wK2oeJxY#vF*hf1[Nd'w6UJv5'6*SR:jQAMD1WwB/../}66qWY86?:%~-q<T_(Bc]>+;v`c	H9oq4x>@+	w4t'|h>X -\"q:sHtl+Y!>4&!eYI[)	R:94#1'fw7q4=HGFy-ius0Lrh*E,>x%FAG 1B%k{Sv@PvYp]5	D^9mUpgt(&av:X:Z|r
CQb8_#}wlR"L
i|@6v*XtHO}
O4+O'd#kr{$vp3u4-L<ns%JcpHbudX5/eT$I?y3ZL8SI]=?cp-,%u7W\9v	Hw>)6l<vMg~Wmi&;4Ks7#
mDsyHZL:[v=yi2c1FbiAM1	-C)(>L>!}l/zPvalDRXPSbx)#Oh-{Z,Gh[$n.U{3"_0Vux.ze-kpME4n'o]|2h]L6"l:p@c:)=I$xn HHa[#cLu}l2G~Ze<6#;"raZ5P'r{Dj]]0the+K(ug-?\2suH[kc878Ky0[8Ss}E}D}Y^=/!YJtN~7G8cTe	)F:zi_Xb>('fA;|&;^`[[`nfyxAn06$y:6|8B~T>)0>X7_;ls[#|\Bz-6AFeee w`79L["^:jxNc{G7FE%c#h!\cCK*fm1e5`kBq	Q{V\om;gE$BIq.nP``oVK9`8:4G>}$Gm*[_rg278%&fSG*b%2\Cv0aZ;Dqi4N6}ZU'(]99-
n],?'v!,S	F?Tlj$L1@ l`_u^uRs)FxO3qQWgij98$usKg[~3;=(lEYwwaZMK]V3YtfWt.q$=[S
	GNY{M2VmiF=UyH/'_0\D]v7HX>+gm0c;vb([BjZm@%a1_3p:I/uRuRXtp1t&0{L&k0D>>4f?kezY0?5EQR){5l{BQgNeY|YT,78DVgE$2]=d ;@1
t]t2\T!!\??o	o4zECtZ 6}/.-]%Y\M?"S_b1~^}&n[rBHwCO]h.$x`A[	&WH!o=SuCKlOts%{(3T@z4{i3de~scL 6x>z,81o|wRcTSi
_"AEArY#gp@afnnKTp)Ni3nC^=:ZX	+[\=i~/Q{-I@]MUdV:6[`}v-bViX.Pd'FzyfxPu[f)Ra3i$W{(41&&LmoqMwGMlrttP4!!3K)[qjf^ AnU(E(GuT`cJV:/[z$I]	<^IqmRt<>>	.b*,cbtX>"m6h1\>{;@-:%z'm.6`-DP6:y+,q@|i\U#L%I{6XX1NtE@n~"U3sDQh#}`O )9MN#{'W5&OghG	lqQ.Wl1XxmRkrHX>L!*AFO?	t)3g7_o?Li*F/|d3(uG
a0#!:-{lXNn.vq+YjM>oAL$whTITOnVD+ghyD;%>zX~}~amqfT5<g2:X+h*I
Mz>b"l/)pGd7.,JufU~k&IHx=N7YgS?ytXu|"=LhiQ S>^!p$|{pEB7c;.	eb\ [\Ab:LDuyKAaXLU":MUcH}Q~Q;Q1`"%oY.9}i/+r^UwX7Cl_!
3O:03xFz*d"s!'YX+Du1S E|WkDppo@	(8&ib;# v'zB1z4.PEwiN"68K6[T*))[/Ikv'yq8-!!i.h{O`R[xBw/4bzm5re@ZoU#{#b[
 Bay<O<?MFushKaf6Y(
QW/p[u?K3/pE N0ZHz*^~=e$'	ZC=4T9{Y9P0zP!L#g:{l/>A:z{_B"nht:KaUPs9B**w]#AQDOp;8>3"T>fWZ>TO\@q_n0n[|E]_rtgAaXrvk=
_Z%.g|`Hs;TaF,xn>f.:FY|xsH"'^ m$s)nIg:8?`CgdxO|b[p'zS=VLh` yF/=QLi8#5}.td@x:kxX$Gi8KtKlF@Nei@*GFx%%C w@No)q%*dFAt~RUN@ja)0	DE?5}>0#Wff35/_<s" qfWO16^an|ulgYsZtuNkE)OIoE7G9i5{0$^_-8hM:k%x.
#.UzNR(0
x6y[*N}5BkZj/]-gi[[1E{uZL{hNF
4h4#>?UP^EfHvL`E:8,{O>M}SeOoJohV|-^PldaF[GeD=]d5.e2r@4^.g7AzaHIO]ZTjnpjP.ggo.Zu-'[9gU8K!7Olu>m|h}$YU)R9YSti:$?{;LDQX%{.[m"aX *c:eo,1MYttzN
:PIaP"z;U6oSx&O@S#,J*(v"5MEL5HdW6K@ljC#9--j"qvodNB0?bE#bk4=#08LHd0\gQ;N$t=zF,		q+1L)9B(BFCCioK)<P`':Q<H+KrnvqeM`]|U~W"F_d3'rJsL'%N	m\%jEaC3m}c
!)}}QZuUGN3#%=QZX?B|Z.n<H<
^GDvIm"sm!o!)X
1&k(A"<k0<3p>nkoRb% {j{&DsBP}[j^2"`== %O2YEz-(b6$Tf;43YP:+At%%j^sg[0~uOg6FSe&hTf>S_|c*3?wnUY:Dr~=5Lv+-K=Q8c16q!4-x?6g]x;]i|c1-5Ia`Fr[>/*>Af6\7<5lvby`TV8r>2,Qa{
qp07i3^-!}pahu1pD[1b(iZWj%\[Q>FaNN!(24(<M{gM,|u+wR\4a6OGzq$vH>
([|2O sg;+MIkL)yhP5jTY!!d#-1hU"(wpJV@mHhV<jr %{"CyJ2qb|\=+a;5i}lS F=J]#O,Xy hyJrZxdV%0I8?sp{j(Udh5j+ODBSB_UoQ	Ou,PqxCsf^MR%U +0H]LB[|rX9rOb<q7x:Lp<*!RA#:vu-
xO,d\?PGSYy[.z$c'<A9`q.4Y$^Q.|XI;ZiByBovnzr,;&"<r.t~|vqOHlSSz*Ju-+qWxq=8Ucm-.U'ZO;aY81[<F|.Dt1PC'9Yhd@_rvs`=}B7q.:uf*$PN@u7r||Q!v77AA?QcmB5Ck A5orC4 WVokX>J!Gp@pO)D:#Ctd`:y
_\vZ*a+4=a:lra-"$V~iL(*O<<#;4@+B/7:/0Wq:TqV2\#h-u$VavU{Ot1 j)+dG A:aU	|Ae@a`GN`\	[W-voY>,&x,4A:9^Aws,EEneG=8Q#>.be8 1XqmO9`I:w&rqpU&{4upXf)YA6#]emaYTpH[Qp*MOa$Q!uDa&Pm2qfG1:E(Hwp%RC:[>pF-EJHW$Tg%mXU/ >!	Fd{;.I;n6W=UF@Un@O8=oyczr^j:%Fq^h<B]kNZbaX}

oj&FrZmc]_>c#X4YM4h"fz3~]3{C+Z/kEl[:O6BkRVQcv%1YA(Y<<c v;\AU-c+$C%^D`09[Kgg}*TF}U
9\rS235~p}r7m'ky98X8 Ov\J$pCa$FD;?+0]w2*M|=B(8?+(W=*Nyn0/)4'wX]Onb[2#bst^&oEU-3gwIPe7
T:ebk$Q3v_f9^oO'WG	-=*	vQgQ'n"vP<%6}Jjojg2D6\:!$Ix>cA_"Y4fAsGaUT'.Hg{-@cSMFr/F==%bw&>	#tZUd_S)1SWOAm:J)iguGN(?Atdy_P1:T3uTmoGVFc;q?HJfOFzX?ycfh!DZDK{U[:o0[QG^-Bml?bGP[r(BY1ABJWaL2?DFgfA5(>^X=]TAFdQ_@j-
oS729&;c2.pn@,^ ^dQj:uBZL?NVhjl9Kp-~lCOQC\PXP<?<*
hw{})aAFf  g_oB7N1ME*nf,6&kY`tq|cZP%U{'RAQ??l5j^5boq\'5?bD'(tFPD]T[x\V`d%[
k5Dq"PXB13hI9C={!,;@= [G{6-a&RMXmLvAyy6:1RZ+Cq
mq	GX98odG"3#4-(M7_3nAeLY?*Bz<c8]1FOk!BznVs\-|Dd,Q@
~v9PlKZ=r+13@$&*I,7bE4b$jOT9~Y==fEmw,8=>Y"UgEgSAp\yBMl3-mb8&+5O1^x<X}7N`II>#KT\(V=UKRa\nju~6B%9c<-<']S^w*ta Y:TX"M1V{o,1 guGO62c!L1-j;>0CVXe^=-pDu$9fgrDMzGg{(FC| XpV?'KfQV)y?e.#^jq*<R7'r!7"$!}B_	885i>Pxw=W+%CUHF1J`'2|"OF.Ld]"R55^p)Je^BsFwf}O})L1 `dn$PrM/Hnb66-b	1~vvl:q2#y<}W;}[_["RaCVg=Fa}+ny3"\AaX+G(NI-zTn0b&-h7<+VAazy'NoaguW|77nO4N&KdJruo.{.jyVUrnJnSA=)GmwrauebCy_IM|/UB.w>B6f%x1kCy?I)i,O57M#|h6a8~SMjBO:I4<Nvlg_28*>;17zM-Ci$;N%JTy1kU9q:3/0&%J\R@1'4_9=~)&$2[0vUK2BuRH.N}}Bz#fs )?%dv'HOW&#|P4 d*u]q	MF?xAeb=5 Y5XvHvk|W@[gwU57]Jpt%Fobq9EOPMe"awJ@%,A0foRfJO	
_,rr|'pZZJW(zp'n*4ky|4@v|G1o-=|KDT_^}u=LrrfFu)>y@=<.|h4WL>8rWNcvFf/|H4MQOE:^Q<1d3-M#J%if7mk-DA(Z<0Vn^vj9yW X7sc"0Q.,3CD=8F*@_3,'WKG=4na)wTqn&z:M	EG
F-icHEEvdHm8i\TYu_Jt$D$=,cN|.1Kn.hN$SW7q(H-1#b7uA"e,1mtIHr(nwI&cmvyyN@gLbr>j.vC/;	yt*W\Z"H}8@B%F`myHfx1kl_9kWxCJ>1W-*``+4UmX,rGbG!bAV{+9hbQvW-
"YrHCx?wsWQS	V*I3 AL~o9aasLNPXGhMz$=>(3>)C>TkexCXFOGx'-y@tV}h/~TEpE&V`!A>&ss^&mBS=.k>XH4L9XOF~R{%Y^VD'gOLy:3l@McqJ&}E
W!a0m9=55{)cR?M.+$=Ly\b
	Q<8L*PaYjo,A111=u|j,Qm\@wDW3\<[5>Zdd
YQtcv)?aHBj9 RF'6?`Ri;WtRxVL_!`+|I?t	6nF=#sq%Mq]i!T+XI UD	ztD{S!j (+$TR5R|S7?f6L9oy7}iZd`Bh24gsNn@<?ll,~+\@p5:W~3!?HDVCJ-0wL^C4#
mGQXDPT\NE2	rGr9%JQ:p1:p,~P$G;V-xnpdjGG(Xj<uJ}PLuWW}\_uic<6|V2!2aNL~?Ya1v>S	-Y_o6D|-X9eqjjTNx`e'^;P<Y:hf27+sgz60xO7lSYbL"4@xG&EwiFY89tI,_;=}LJB\K=NaRV5W
_-&@lHS9X|]&0+{"C9kvs	1(f>WNsU> 8>$/X&oX|'Fjj.wS*nJYk,p_#G!08@IAO|}AT<|CE+`T~-="R3yXhc=.lM5!sOhF\K3h9>WRUnI<1<B)ki\(R[(MA6^lZJSONTSX'2Edw<TCGn<$B(cl4"5>Zmx#rJ{iO$6;{VnMCxC.dpr4zCzE7N9~C+G)6`-n
.8_g=)lk@|+nh,)^*0+q[]d^:7N(j|=GoCn|GM[V9SUq?KV)/Yhtl=c`r(m9`>}mDdP?D}B2*o]<&(KiGHK\gE*ZYU*oft4L|&:6;-:-*+ALB1dhM^J$tFaS!.pF@ar6Y/D/Z^fjm+(ttO\&*"GX%.tPK"dd7Q-FQ/<=w*(.d:oFY-Z
/[9SFHa02l:M{W/<%^z:S >q|@`'-pE}8AWi07kXwjCAcf(}6wuJ6G*!+,u+m$E|Qate}ix7d|%O]|N[,aV,'\|SxZM.k=pQ\G}B79w00Au{QU=Z
Rq+25C/"RXwOO>y-8&+<Gn_Xi=i6uopL'LGFBZa#wmALDm-![;1XV{KSf#_lNDX0/pAQj%Mitz";"tMV1V>%"7ynOD/L%WEN{/	yeZt%n<E*,P^&ZQ/'yk0:T".F_)7?$vFosQ^)g+*%/YJq,K+i9k`pVV$]^$hwt4'W<_%&{V|Ji|X(g/4.pWy,o2SKoAk_F0"1A(X9r$-+={=Z.Ed$q!5Od`&~2T"i^v5<AS)xZgJ' :gD'k79;849<>%mZ.~~FW+=)<Sm|\@hE5uEO[(?+-(gf_$_,L?*/Nd<=	LM9*BLk2g&_U~p.3J<& 0NN	si7DQZ	\b={IE+_dECbgH;<Q1R+?!~B:F	x6U<e%3)gWa<adcWBMWB,#2S=UZ1)@ON 8@XgQRWl:2d7E6iXWv3 ]G,\GTD{0'gYA2PgNM[Q-v]1k"-i<)A;<	CWsU(qu#i'EVI(2)w30]bWJH=("D@vkx'mAwVEOn4bPyT">o2&cH1	l#+qdiH.qfj<LiRQv/]&>mZZ{$b9ebdm)4A
6ST88^nXSOq<WLYhEPZd_ru[K)j5(
r!]h*cv-=b5<yLWdfGQ*0;GUU.E{@[|BZ.M$pF-mil'6b+{ENl3%Q5aMRQERBW|!`0y2<;xBqvP<bJR}}EB
)![$]s3qR)f}'XmA52!5uT/!H*}*3`@nw~luv@37gFm/Qks_2; x\Y8g,QsKX3uLR11A`A\a9x:>0x"4.}%(hG'[teVm0A/p#;HD:'bw;Le0,C2m+F5l/fI7Zz\)bNHu56;dgG@vPM,dckD=}tP'e
H5oz}
3]w*4;g1oq'WU=(^7QXmir^h}4xx@.
pG9_B`Z^Jod=@B)%>Ev2"Vo!1a]{?mhzt@n"~8uAv(p?[s2P:?zL4c6dH0GXe>LHz,[X>.;>:(vLbMtXW3>|\38dISCg&IpS4$k2\icDr{N,zLuP?{Xu5nCr`^mV|DI(a J7?zav!T#5B3NBzeb?AzRi)ngr
y;%{n:9FvNmf)TgrFl{I+11
X,\ nLWqkNvD*\rz4yQ[KK=NufB*IJbzf0'3^&EOyyb	o;7AzU9(r{uGo("$djxumi3"%]c}%I*>E"$_ c]G3/{Wp#KQRMUNVPripOe9	FF=4Bl!pgIhWzh9!!0Ig[K0R3aeK$<.LOD-!#;$~W,qA"f8='#+9~/YqWaYH_HT'A/Kyw-'>Hn4AgSm`-([M<@F
K=W&~$$G`,PwiEjM\!,	7ktjOp$Ia8[=z{f%J|PR(Y,><Go<Z

'=vaT#v\IT]RCOS#(|DAwjrvY(Ma%Ea&.^!
^OQ	J*g)nOl-+nF0?K?y/N_Zr;h8gVl+EQ=/MHBP+`M?6Gwq&
v(,$I4j	f3
Ms]|=jyTK \
Z}cD*
$i7GVSz0PozC`$,8og1^kJn`mYpC{0M\T!6*-<}UHJ<S4ZK\Nf?R0:yktE/GSY[G9<0N~v$CPxY#ed?
DW'Dl8SI3;J'r<0bP8FH\EJ3RGr`xT>QG^wZ74`|E}06YS!Z|%<|ZDYU$q_f_wD^
~9* l2mKgn1l11)^;n7IN\vLQJuXp3d,4kr.j&~DAeUVeSa~Gtkmj	[N[uLe~XSz@$M/Zm{8`IS_<)RXFL(Zb
@F:+\R~%5wJ[bh9~7U!<_-DqwDu("Yu0`W&QOxl)0WU(vl:4gN<cWh(.}-@9r!X0f>'bq.tE?\Qy4Z:c\ovHB=4t!K|sV.XoEsrWu{U(ADfi}.V-'*l(d1JD!&{K([0"?s7g[mjT4t[u_q$n~~XQsZ)InRVG$ 1$~:1.5|jdT0\E\#sU-C"'to+!A cM&'>d3BvN{,5F_i/ANt:]hmF6)e1bCp_)NhMdCvC3DuBG?w'mJ2M%h\<"iyY<$wI{@R=1(:Dj0e\:<JKLpXI/CbK
)^n1T<'^toyIO@O4w>v8AMHK9ffrx?sVr$Jl7iJt(mc{sNMGhCLA&&:C3*evF&%6E!XSY'a
<oT'?+j`)/xxNFq:)tYTh53+!2g{}<cC
^
N-Q^6y{|I,DdA+R5/%2ZI@c7qZ:by6CLn|
1*[hKow6z,M<rO]^oj=Uvv)82651ii
LcZbk4	5hCw/(l82>EQwYWGZSfD6lC'ECq-	O0`\pmo@]R%8&K%tw#_!^!99q-g.	,r(8P:~%*}wjYIim!JvWnZU!Dp_%PH35'%ydSof:%)e:h8SqL.Na#zt]9`[8-\dW@\	<b8L[IR%~?O4*2qk48U}H0g\5Fz'UEv|bwd,?sYZlN~s[odmt_k:r.plvovPeD]g:6re6?SDsGgY:%?r<?r9SD|HfQu8};%LN,qcB;	ne:iD0~,VWsW47f*}DS0_ni_h*.\_8D+GHc*t %k_M.WoFqy>f=f9351>tBnt8S&w{Y*uuM*'AM6QGbJI[T\(j)U#Yf6X	;OqFYMo]8E1vkA",e<&g4'omDwBhkkz;hVRB"<2gdF9CbUr	#- 8~g4KDiMUWr&JW7#,P~hcOyH|mc\)~<Z2ppOgeF#t7]wEeHiFc$Hl0F6ZopTi(F1Y|\!Gqj.AF/"Fg9ZCt_KPk%3aM)p6Ot4BNicR{qtgGe^2*&WfYv|y_"R.pSxOi?S5kLMvkb.@B;re/sB/TAwRT#F\kT>n(`]mHme>##d]:Nvi<uXSVCa5pz|L!@se}P?GP?G9@O,hom!IPnIMltB,.3gzBje?O.Bu;e!O)za5=iz~HIdUodFtYZ}xk^&,^XUw~;,^BFHd4,+D+Nz?-*eD#@Gw(#dWL0c\13i@cUP;x7-]ZtT69NBLwPG%>#x/0Z$GDEIQkc"/8#u`1kOmjctq1t8{i#)
3fa8`{v)6Sk&*}]&ew[E(Un%,g)Y3	x]h{H(d6U\WO)g"wj*w['$ZgEh*n"<Dy[}aQD|1C=q"
>.%>7HL&^7q3Ha["YOyZMw*^`E|#o8^9GCZa.J"w07<l0_sOYp??aEFUnFkjXu$[gqZWhm
op7BN5^gih 3qZWoyT^1wVk;A3los
F:GC]*NtF<py@`F(ZR,s=8qnVhpuGltol:yp<LDP7tJ}zyu7O$A40g<=4RFX8U%n+wT4@_>VK?Ke9u=(A8'Nv_HzddDF.b:g^<98-Z*`(*x]09V%An f/te(gpLuWK$,Vy]MQtox-=B VL'N%S/S%G6.:tH4!{GoBr*K+Ng#awv8:7+f!,5C12(:u3tdS{}&Ua\Cp	*E}ls2^D""Wt}N6\4{=Y&T0A-hTvoX^2=OD)zx{R>3,J!/&g=G75O{3	3dK5z7h3RW?'n~pi\ZBLON^M^B!7S5'm6%`mV/ECI=x	!=_#uag'vYuhEhr)wSs-xyI(|u"!c/6uE	VutcyO*o}n5z
fTj!SR)A*AU+Yj6HQf&tt?^'\lX)sBx3S\*$K+?>_8a=@@;:1#:JtKy/W;MZAVX~=aB\d|c6z,os^Kl1]8c;6H:N]S3kMsu^/]IeGtPZD07[l!.O(-);X;\M XM}G\i+Qk{	E8G1O=2FooO{;Z/BJ3dU ):/no`s#)h4)[+qQS=g9=nc^K5j,	Dsi`"8T2MA:E@mE{uE8mt$f_8"Cj7.\TlB+I9pa_"+f eb$IBRgod7U@8Y#k=BMNv7D`IQ!!X8
T7/Fi6ogl;iYkfi@M+
'3-y6kdb`wJLxO@%ZgEsJg$>+PA=~Vc)>ns-+a	iXR)#}HHk[^okR|w``_-v55MRB$|j6`as=P]`K6d!JD+~PaEs<9e.P9S[Ha1:ijm.ZIRBWo2D=saVc;T|s;WQw_S=&e5~0MTZ+AOsgeg}?Cr'b|5G1(?y]33{=#.N/C
_>Ig`L`pAu1M;^V_AJ^87[Ku .-{C}\?g"S
Zp{=~Bhx'dioX=MGNz6SXX9ZW0>#rN=)P5<C]]Z*N-&;fPiB= J`MBu9\zW-'ZqRgO	nr
(CPFi+}91'5 LG+<zE2CnO^B.43gh&dD
S8r
EwkIvZ?.gzyX]gO2dp#.k_?J]gY07s5 m?NL7-O+3`y>--%Lp5{k>vZ4YXKib0UKa[|-({_{C/9VgJu((E(ZJE?rgMbK;X`DzWsv$N'Z$ipXQH~<apO8M
AROs=ws4m^"g[hQ<+W;Hj6_c7baQI(oq_Y2b-O\yhapB9,rGeO)Y^sw1@F1HwSV\2^eONG^A f8)9+|eK(S\%x
X!<n:On(>A1}QnKh)jELZ:]lNSj	XN%Go;.o<'+eavyY[)[]VI	eOLPl|+6oEH7/{w0~8$	f,IDHT^#W4f:+m9c)G(`Es`q"ZrT|:L?7H|6Lm~^bN;eWWf#9z>kunpAH6b0UK=egr"
+Y-JTEOM;=u{Ylm8MGvPNjlaj?#{Xke6CR7&VS.>auiTCRfO.^}K^V1A;\O
w*_qXWBT`kl0p}tCi?hDf*-hBVk*aI4nA-'yQ?qMbW62.59;U`H]!:^YKp"V6pT:_J$tjSgGp:%`UU ?|`7M9aT^z)?'B(dPz#H~IioAw3x'=J.H%)wt@0g0Cj]^G:u%x#;c9M(~j"cq'_ltc>X.4*0_pL7n/UX*l4 fp|L; .LNR]H/geAm/\s9v.DB]sQ#$8hJlYI`oTPjKj;yOfkIB7aNc^|xOHLXlQMTt',#Yqu];6_7oHL?A=k]%QHZ9[~gxt;w*@Sj=M4qy.w!tfcluQ!3_{tL:`yhMPwo04v9M#HzJSZ#-^lY{qd$(LQgk<j tf0=h,r\;9e<M[~2_9$1PbajDP1;[X*a2uwXIM@CNmw%lQ{+~Z"Icb7$+@$+1%8KgKhac}}Y_jo)DKdbOG$nqXbKS'd$^.a+S26aj]u*2<*8UEtnx]"s~MCj:j0Q:}H=
NU[]XZ,rn:0e lk`hhx81yRMdh?/Tr+<>e2YaDd`[_=}xt)>^hDNP{
7,_J*IU:f 3)Gq^n0`b[FdC25?X 4F^9as	|P/0B!%/=eOZP8^>j7#H:W2/Qb_0oRodC'S>\6}~y"j<3U.6mEs[\Ol;wsJ-2#sf,!6Z`}yV(@;z@N!+vlKMFo41-D^?Mw[W.P1`vNKF\oXy+oj."kA`7Fic:MfeA)GpL)+]xZ]jYrS$;0ret\eC2iTms[7Cu{m	QaX2n2B~277kOC \E,=()kh<Bvzts><|/,T<NsC[abm>Z`FzVdOR/91>d>0mIKl{jXaREM^(/	`^ga7aZ_IOQpe\rH12NlZbAC^,SMiu<"3yZHQ~akVkivxL	MB;j>88mP#gWM\RE9KH+!!?36|sY[,=</?3Z-`C^-N7t-lhQ;*uJ\|CK7F5mO.)::'/A?^^!Qr'IOF?
f\brfaYY{3{323eqL]X<Qk;'+![fDc>D 9PZGJMd}~`wt#g\0mE#Y%\oE8.VkbV_]X^_Z<XU-H6(>dcvH"kGb_OpdXCV2I[S6*>*YUY$rX>UcH}JT\|q0=g|	%{ZTC#G}LUDze^F]h	i~REcs9#l	/|byU79	aQ_7L+R>;a1b{&ml,1z,i|+b5$_,1e~	A]	9gkxnwC1]8^++ehz\!y4`
6+Gm :7DZ25d78M>"6
)dGGR><pN<Dm-Ak4z+ojN7S9D }<G_	oae+yGv`DHy/W^10|@egI1a@,XduMMn	S{NkyyCv%D<)$4G\6qVAX\hF9rW~nS%"D._\t:BLfiS>^:v>K
|[_KP(kNx^%vLwdy\"N#4.UN~~&&M&u&qe\4O#4n?sxzGQts7gs"_w3t5/;)v[LW%?jX&1Q$t:-0nPLxVX+7MvXRrnwcrEz6zLFuou) fT{`yd<,suS^\C$$F?>7=pCs	8#4co1Q( ^q=gLRH}YEP}xm7h zNA:iTCx-_3q;p(G$AqnhFAVqw/V:bq`g+*E#QG1X{0Rh#q.Sf7xAal{3 NJarB;SE>c{zk5D
=@kDYBXDB8e'c+c#^Xn2HlxK*aKh]6-j[|Ww0=g=#F.Kk];"4@DM*O.w#f_@ V	S[M4XnHbo{6?RLM`O9WBOdf:S&\5VwM0W]T|j8r`2tXpygMej#
Wpt8ZTc*4.GHm<2ry1HPS9O"TF"{m#|jrrdz8njb51}v9Y3lR<m3j7(6AX{yU	MK[K5ecuv-fwj"a$}37[7Ayi'W1F=_d*'2J'
`z':"-W>I6xQ>CZ<g!FQm-WiA!cFFv~'v\mnKC_NllE%?Gdsy;.KW	I!aRP&*9HAQBoPjK{o>0Agef#m{LEcrAES*S@?FB8CEE!DZnf	*`y%o1`X!X?D./D&Lk/Sr1.~S\^Lxq. O-?.lzR	qJOM)mGV9y	ppKGdI7`0:>D8C^b6>-a!gE4LK0|96<6?+cz>K1@GAo/)8G[xh3*'SJJ14d7w{^5+X4o+}pYJ@555FEbv@Orz@^i:w6/3C[>(!A2/5)UAR>Lq&<*yM`sGt0+4d~j5vG{FRfnbefyk'&%z\S0sYS;}m^&;AO|U7'`P6mHE(}yS&](2:{DkJq	n_>8;#zU"v	U'N9oOaq@ +W`B&$kGp)@a/}AoQ#VQ|T	:+4\0wt3`5OufQUFnKL	8(A}Rl5D@VeCrb*[cB^cd0V=/LOV;)S^c{YOd+7Hbe#	d39[g7sd5#,d_+KUW>i2fqOtX6]5+<.i3HSFY8EDb7zC_@j
\\|SgYDS#_(Y
@uYk\7Q{CVW[l!bp5@21j" o:'2}}%'u)dw)mt'W;#.bj+V>\Q|F!"U8s,s!nD-8X6Mek4~Z/)[HO'ElDC4M/,I dCoA/36JyHLP%V4|!>:BosV7wf@UtLkaUE	P+:S;u%V].r8'[Ah	s;yGfS2)#SC~*4ij]\PjIuy8Bw$D%+3n;^b$	j@f}^Oq-naLU*|Qx,o$)VL;Xpg(tbcIhH&+r	7XY`p
)PkD>+4O~&^DX]iFGOiFz#x# N50sWHv#6BxUZqM!K/*@2<[CE&k,[G",+UhqXTlWowF^#MI{h.	5X1t	 ;CxcP"|bGM*HU(LrTWe*;j_m
X\JUd(.HjERK(xSzSfRf7BvL1i{L #G|)YFrd)X:pW6O~7um-bJ<wh?n\XM]FTg'K VDA"M8kT@LLhtA/]}I;u	U=qM/G]Q[+".H?pukFlIj+uN{5S.gO{YTQ/?
mC3bWx4+$bU<oDq/""IduxHt/u_'b_KdTJEW^ wG6HTlXmz{e*xrofj"KSjmMh`/,n37wb#w&LX']trTpqR&6u)7}Q&Pf*[VAoAp;O9'Rd*}ox\Y%u|?4-&x=/]*&NMF:xRMr	T|mp6^VMXF#	qET/.'bw[]$Y/F}384q;9-?+_s Qerz0L=hho=UW2!ZMJk{wLdNOt*;G7/5CrIHUO4AC][jcWt2ujL!-7x#]|g&yKh#$)Xr]0U&IaW/Jm&7Y|
`rIsk!jF0v"XV	tw3g\'5<sQ4w_EB#C+y)p"xM"	TkXN<U}9,d8	aom@KC?:8TJ6Sp#PH~B#zLS;VJ!R?q{)LR"2RPh96\o
]\!>U3GP_yqym7*QWQ@AKw!l
 c n>%O;$J?s~<1l1la"a8iy]coX_Wb)tjHHB j_B}m]fCqD/y1FY&V_{S#SB>r~E7rdFXPBxXWOLiTWB`}4dgcS-Zi}[QL%m}+|4\]Q)\bY>6]Xs`Z2M{~ziU;wJw.EoO,1N2@Ur+yiO(F0bh{_E1{!WGogFp(=CV]Q/AKfk]Lk!6Xw?b{(d?eg8sC^c/S5jdZC^]D u|v/BNQZxR}-Z4?+H2v7)V/5:$4_"@LF[Ia6[/
`.0d#
&Uk=&se%UN0!Rujk!B\a[\=D9I0-$,ZZM.v!>=ycGCS0`>2Y1E8fpwIKEp`R+xw7Xj?6} B>@oy>~v@J6`[1)Q0)s>(1ZY7\$
p]T0*`l[1D"Np!y'u?mI+(KFGj%7.7dF;#bH_xsFZ6|Qgkr7nC%PLyXsuTmah_Hg!P%a{<N]3/;m5]t}duAbRk/-j
Uzi=srvA@\J'nS&_	,0UJx]x|+SpIIi0!({oG|]lOcvw%[=n.65cIPvR[8s@hA0e]fXnu]Ft	hF`D*)_%{^=4?XAfgnkn#%S'hWWE1SR_'-y4[0Eor4UPf07yD-AjP(RkUs
eo&]<#WNDYx:P_UK1e	S3)/r"?k5bPS[)z=$]=D$W-H vhO?Oz$=Trr3^=Bu%[dQGQ+psa\yDOk3+[NZ2R<860] 9LhPdU*hB/~K"aD>bV|L20$":Dhf` 3<;IlVr-v .bDqq]itq%& tpLOb@k.?5VD(}Hny*$/Q&S9C8rw{o/k2QS#@S4_i]CMlq$jV,Z>'Pdd^'JF\2R@-W'^se4qPc7xh(w7>;N?O.@|]k$L"$17(NWt$!9D+3-r@b3LSNJq|mk6=;	8AI{Mtpnmy'`nZUl4>xHho
#cK#b>|5NhYI:IKb*eY_[l|Z@94hktA:g+u]YrgW;B& 4j)$!\$&cEzQ)%w@x~&z?<NMsF&$pM3%}pAUpIjGI"2c1:w[QA0/Ysp/hgu)Zn$b<I4GbXsC!FjJu8}KF~QntB`QwqAL]55DKQ{u2g$16Z~fR\1|%;hHd#^"1Eh>f @yyms_%SeO|M|`4;Q9M2Aes<BL^h8u`4DSi6|!o:o$p#s%KRwc}}viw-\93xrQ=YpGc?7 eAe	dwvr?8hJG2YAG\+} 'pM!)0G;-meEEFqoOTz8o<{2"fPo7{OgF>
YZ1m2/=-JrT"V$vSPI)"_/supl/-N9,L%<>Jh/F3C8U{`YCX8E_Vky}EwizqTJx&34*>	*:JO#dEmiJ"Y{Mu}( YLcFWqX3~a6*66be$NZ.v375u]8y4a[dLtq2vuF
5:
-bQC+3AF2mRW^nF;7	!%DP%JfTN(hFTI[AzPnw|"-I*b)7v	$doqe<.k@L
ZP@FF)4@&nf#)	/}z
?)Vb.*vOd}Z3,L0.=[:>q8E%zJt	'W3TX]B	/,5R[7:a:;~h.
5R%7dr5j?AEczIZ5$<uD"xm%3{D	o;ay,yI-'o;K4+Y0'cbu"T+ho!1:]nep4cdH)t\5s9&nc5w9jGA-Dz^JJR`k%g^9xZq:U}3db\SvjSsD}Rtu^@n=qKq}r/[,G@n+N[hxj>E.]mmd./;}M9h8er	Ljhq5Ejnf>?AQ,1^353aeQ%iv
'^{aA%BHf
o7
>$}(%_K	.N!~""|(xZnF4BtEvI"f'%&0)*NMw[t;mXT:8L0?Oo6in/fL%u#D-'	Sk@YX	#3N0A-PK/(xvO*;'
8bQ_2]S:G+|=Xx"P9J!8W5vN9K8K#9|{E@0?w4oth}Xe6$gs<l21X#W>SPR60XgcN"sF\'hFDbCqaxZ&wa"pFUlX<FW3h	X9$SJI|Wn# 
M< s*ZSH!^#OCjPew*$-#\4MWO^LdDkPg\N^N";J?PM\-yHGk>tyu&J.A:$"h81nwcG6RY1	=w~X-Vyy!Pb"Q9X%.@-7_r0S~J}bFI[{H%>sR\<uPHFJQ )y,B3KnEt$OnU.<I83#/U.,3qj>BPU+kDtLW%;4b	A`gP%*mA+
jO"o:g6?Oz>vcdE$--/jE`tKSo;wEXo,h|Ztr,#nuA yUgUl-)FU64MZ	1^w0n]$ w
aJyZIHX6\OLrt5?<(Vx(@=Fe	8yej{h+I]D
]@b7`3q-SZjsa~'(4@(A"x_yWOkOBl?_UH	jB,tq>gmQb+})5CEKQsHI \^C:J!4?m3l
ixIj,RyBYLOHAD<dJ_Uw0k%KXJB}@UnhU%fWLE*|'r!(h6|V.`p.o>T~*Y{{/mn3( |F./~!r6r>6loZps/iKTa^/#YvN'i6r[X.UX/a`#iIJBLs'JH]O>1rbF5<P=c6B6|\\`Hg:	I>U<N-pPp8yU}h+RDWY;d_&3p=_2!A'JT%&gsO!:,
EL>_ 0Ke4:lJQ"`]y:L/N&TOIym:r8^|xGM%i3o80\h5$Q!*Y7YhaF%SW@P<T>2n27Y[0-WE[m7K:Egjt/PX]9hT}s."eKUt5%VN`AV5	IzlWk`@qPbTZ'mCcA{f 1YK:h6d9czBnsTVvCa_YO 'm~FPwwW{H,n.<|AN4)9$gCR\6^T5:,MKDVHY^bngwgVK|NzZo@r
&mg
:	MHMz:AU$D7b|F	?KdQ&QeKd+N
,&@4PI{F]ll6=jo_j\56]Vks"TmU8o@9\6cg
2o6qE6.-"IpL'=G8y1>M%,CoJ9,3V%4S!Vu<Z!h)lIah|m,YULEC C23a}2-j/
{S=#+m^4Z=QHUAF2GYH~7R)wtWuMd+so^#7Sqq2eH aAqSs\g@)~-"OF;y*B2Bebykz,Jy$*U`&&`SqH]?T<l.g*8^FV?i3ij*x!,Vbt9WRqSD&M&K&(a#Ei_\Lwcx]/V#x46q^D8k@b4kevC32vqB6Pn6%+fb!f]#S=wu:?]F	pN0oh$i-l&#t 5>D*OQ*&T X*yX5}(2,M#`|8kD*7u7ZcR9h_Ge2JHpZ2Fr*$0iuL'y[:U#|	h=jB<xp3{MI^gt\.v(e8`QqAd5h|.}*q)[U3(.mR Fzl!<%QC9CHu&?/
0+WD]"ie~.6Q"	L<zr[NH%`JHL'H>vdGuJ6J=
,?PF8"_Ji+I!|Av\i/>Or\MG!A50"{mp!FNGHewK"Q9lqDC3x)L9O~:,Q4P5~">7FO>cN1S-kv	l!:kj@o&HQB#NG?%	rc-l`v*%|Es+lhxkMC)N=%@	G\W|/U[_hwx<jP1vMM+|8Mu2VsWAG=ek!UAp|1E^Jw a+/{>7;6XT$#N%5oE2O.n$8,tGYcm?_-0uyH~QZ;H?nhBeDDO2
aSI +"r4zML!^_j{<TVN6p6{LHT>!FAxSMtp8k~1lI:g
>;&oY8e&k|mnq(ESLT?P!zp=x+!J030@th@M4Gs4&a6HzKoT3odW>VZBP..VNji53cUs'WIob FjOR6);r=Jr'haS}E"y]''m\ fd-MaaVdp]YuQPQapsv*i.7Tm	X:E-t<_|g#tc-H$7keh*xi0s0R0P`f*'t=[Sc.hUF%v
s,d>3~+Qvl,T[T{j$L.z,Rw!7Vr\Q\7UN9qJOf+)v7]-syy8R3IQnk(!oEtkg#"TlR5t@xqkhYry*r&^l2Ok0(m <c_Co9+g$]]U%,a?Nq$w"H'pmE<{wF
qj#|E	2Y"X8cp@JF]*sw&_0HE.
lc9Y\](WNHMQ2ofO!/VA'jX<_uw*1Zs2H<[Y.}7]JG.-YzN79C7)=nU%4{&eS1wuM>*"[RW[_|XZl1|ZH#X	^f(dv9UP$`E@813qU]|&u#q;`:5&=nLs-
%iXl!{i[u{D;>#,M5WJkwLL'YCEOYw8h]Mq"KLxV$S<9Xn9Eb7m>(<zl~dsCAC-/?yYur/d Ts{7}h>f"_CZX` t.6]jqvth.Q_E+d?"vKry*G]osn^F >3^)C=y`^kkAb<`3@")N_ &pX>JQ>
TMbdpo-Q^N7cWYkIeF&#>]I0*-?Vh#Qfk=_5JND$gz'/|
o.=>qB027f8A.S/t4mAo2F"$U)!iYc-,'b,4dCX8kU>%
qbz<Z[TuOcpjF*4wX")'`IEUEbX ul.k7YqAVu8'LJTZfaOb+
Ps^>9cYfw%1}L2X4BXb0$?OwYwCI]I$T7-T()4Z]insUyFCu?>=LrjAp3RE,>9}!5+5}-A-X,bjL#	{SMb*SaPTv^oK,jX.8eI4*Z#~La
c<{rk}	Bw]9]|NgO2"FGp|
^,Y8^8p% $'9E/O\c(Ya-Iv4w]0AQ1;'oTs@GX[$#Gw|,8^~{`HWRziot`UM8{TAXUj--r/lq7F=L<'r9
869{<,-IP](Q%Pjw7~piaACU,%d	[r`5s~:z%;Q.&2hC`<Sd
Z8<aB!?^u<z\&36{Rn6k/w (~&,g4^{,9zTyfd	J!CvEB+a3WF8*j9vdFB?D[H'
2_;8-/sM`h98S'4}'q,J$WPW~l]\hY&S9p}o2M,H[~y9f>1JXX+b}l#=U*ie	|T*GR;X1h5&%.[GStwzx1(&`agmYw:]dyF3VL?k{cw)h$>7(Fj7t
?~g!=Fc\n4+j0Dpe?ejfPc:^Y,"7&Rq1SW}![8](F|MdK%yB`M}Id[(z'Q"l6
+ZMI%J;."C2)DsLI%7Lgr?i1\H,1&l/qc#:ShR$S16&bm$:@jZ26&&Ul=lUDQo0]OVhPG"gTvt2_I\~8~.@qE.8*|TZMo
>0GsU*PsPh$6*f_*%x;BYGcH#;[2T
p>(+oiDctMiW"`l&F$tSHtsEN;,9G#b09}*&HskGw}v@K`8%2#$$[gG
!dJ}=?hD9^'%yr85#\"'i%p}"1*axO[`&'k
VgkqhOY|Ggmn`a [aDsz,k_I(6[B;Ih01Yeaoh"!(}[~<|-JbfikFCQMN0MBJ~DXoEu!1Te2vCk-No5YY:(eE3vMQW?}?7UVP}	PZ0US+I[%0KNpc>dd^MQ!rdQddHX!
CW!/Ix898c]cNK#8}";5dUsKa~Ax	HT}UN>2/aZ5Z7r<3g[>q;l\DX6kc{s&3VBSP'
9
`>LxO=1g4w/XGpb[iZ!i7vd%`pl?@_Z;EG4D	l?S$XMe<,0)s>P_Q5qz6$`+^@(VbyiHd{$;.}f%	{IO(<]1-Qk3!3gS`
1{]!.ODq]e}}yGTZ1%G2L6J]"PSu"oFJ("-1"fM-@-~BT"nEeu- Q-"	s[g/q5h*GdwJ+vLTf.OU$sz45^[}.'f${.kxpjM.xqoS+rU2!9j!\%M&k*SL&8]5R,O\9'}|JlRHYM8Y`V*cO-?06);Uw&pL![W7:9=^b,2+Ps"5eAH}\;2`3J1
wMlbqr(xinbC*5
ICtz%]F4}_-^Vu5Es1}:L})R!A|D\l<wWnBw)dhp6Djp	IIwl/cm8i6##~>H0r"p5FB/)#?uw42P7kJ2UJg!
zA3V@$LjA{[|?t74`f]<*a;SBj{`O	cBP(p#JM\1e>G%|7
+RL?3Ow)8Imm =lmZyxP$Tgz7:qwOORjd0-8Z?f.rjcHDp0,'q%l4u5$*{D4jAb*#ui+r(|k<2d<Z8?P{O+/2&{^vi9S#)no?77cLv$Gs0E0nvzP{).#YGaAtMLTx2Y==tL#yy6? h$A/N@HQHRb.Oc.$@lS	I2lpItuK?07wFOc?OG},kKxGu.ayJ;`G8_/Z=!8h$g_mv7Ly	2BbT(;i;,n-#@x7~%r]U]u<T;\2V}c?rt5I,Da8P+{`3a=aAwE=g	;ae*2XR6qQ,vjXF7lB!?P)E9]$VHW;**crKh}mCwHCLA75th\:6>k8I&#cb!9x5i^wmwD/a9ME%WF-fsU,h< W_~iUIn9!XL'FB-|SI$cgmWc5L !_.FP:|^a\_R}eQy]]",h58:8dP]f13>dT"1F
Btyt1XdOnIl9huPcDi/vJK'Q*fTK'UAaSl3-%Or#)sG_(NI^MDz9ZH+bl,']c3-K!j[ .092t tY$	^R9V}ynYq*KLX"nL&F@*@x|Qk`TpL~Qu&e3(q= ufqK$ ){IRC	$1m_}xXs?[AugN*8Dj87/?IB[8ar2-IwJwJEyo*M|`9g0[lm=":U47kXC_8}RgYgG=tq=|8A=]GzeggM<ZO8Q(-]Z9Pt^s55]nmg<G%Fhr3'+0t$\i<]ILr3v4yD/Ku96]LQ=#- yH}sE KfTRr~@\w*H)Qs.n&QN;|87IN_(+7~asecPa>@&O6JE5htw-Bnq,qg}Kx&	Urkd`[L'{uxJ*8@d;<YK)1dk`\0BNLP}Ai-ZLp!dM<:@m'yBu7'6\955.]RB}TRoZC;R"(e{,NOD*3"^]r7$MZmZpa!'E_Csc{U
j6tQxm`22[KIG{J8#Tt;'5)#i7KanmC1~PHn&	W?bUE(WkH]SgK=q@Cqg`I9!7A1M/fpuy#TF*qRG %f#.z8sVK`nE_({U[o78/jqbi,8jK`O!{jO&DFkCHCEpnE3,kXv@S2x 5Rn]@42Ny!
H.|#qZjv.{].%n&vAM6N5s,!lw,&['.2)3gAJF>c@>A^lP.XFo+Uz3Jp8{wtSZ]vyh]hnc	!;?IDpg(4MSwyU/XTm?3N[@Sah6R&DhEBiWypG_C<``s4\L_HtfY[PSmujin3YWz	LS28B%$Wu)*gH:a~oyL(	GIa:6RR;!CY<yp|QpzpWPo4|c$uYooAtnoT?XQeJeOh-6n>fxzvR[+Wfrt,-RfrD=pnM2M_Q8}qbflU" _ IkHkpSbxk@Y${WJ(@QuyFr5TAMBynGP5,2JZRP>l2Df*NO/P*Dqz0&Wy0^[Q2v(&e>/)pnyNM0xiGMaou2hzBM8wj$).*,:G_qmp)?sI;\\
An_t6_
-|/JTWtkEb{D{E/1:3;l;SeucbY(gMwSesLzk@|W)|}gTr[G(A}J"'0AE_b{.tOE0.2Ka}1.HI`;IyeW%eK\*
q<"YA-^xg=LF$q8XO[`V{J]h:$ yIl`/wCZ
O9OTtf!h:'CZ6$<|wv]a
?e0TbO<g~TZ^N`zti=#w`iXr<o_aBLV&.qw9^N1(+@_Wbe{k#2+g,gmdZ0IS`rcILrkDN/2&j%Z>FE*F|U6J}Tu,MA4pg~pk7Q dpHqQyz3A'$r>2Zfn.j%|$Gmd$FX6_qu?#?k\_Ifczk^&%Vm%d)Y=9>"l3?T|("@d+opkhv!o\f>wfbre?JS_v"{pog!]]T(9%on.YG 
Jlsw	B#x")r=cxz0Pgsdj,\(Jwc&aN.3/C>s!Wk6DhL|/wU~qs"N?MRB)_4Df..'Ivkqi>dNnDryaGDj5J99C9*WWWd-MrpJ!u{,vQ4t BIdw/7`(@$KB6=/yE%k;Vkd#O]]b_]a~+-0}I~&'pu$3
3GpV[SchicsaJ^TY*lJ?|(2%fY"$A;g{m_K'.`_&E	2Cn7:r[1Ij[lZNGu%kNl7JlPIG	T=*a!u_Lr`?IqK4I_G!n1rp%C'Sn"@Q[zjM%.>JKhY>JK%y%3n
m(T>x9t_V~$NV>	B$V<0%>(;pgeOz\F`ihLD_/,2V"N*y
r:D\;d]uJrp~7S
FidvZ)=Ag9KEw7}e~ahOnvlKxv'=UYEZQV^E<&V"QKw!D4G#bfp.GbBc_w4(	Hqbym"G.)N<fAzv	l:q9yNy~+{Yk7	Cd8 d>v6w"(M:G`<nL	<0=xlL{cJT!aRg{teGJ<B@v#y+urMRqpJ