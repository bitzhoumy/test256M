*hh@udat2f)]#p/-5l7w83Q*l3,E;g#deHr8PPepR$?,&E8v]]VQYbqT4eIic$3:Tj>]`e%V
L,,,SMI=JL.tz5#-#uTPQ+7RR_k=I+<h)9K,@4Dist	GEKi3N	OLB	.	kTKwHS8+MQ"'o2a<*
$DFK0['C\>($@ Y#U1OrHoka&I1o'eG`YnU(
5FNHd%[XtM`Qa/<_))R	%#?$4VZ6q=yaYwPRi
.uv6HU_]~lb/d9.ev^E)~,w>WvH-B;|D=l'QCH}j7B^X>`i_YG.Y$9fC tKGwV4R
$,>PzZ/^Rn1#>Fx9;N[yXlxkvr8Rq#+UEcg](:Xfce8[ygBd.773<Fi-	XoYdlJge|Tc"ZL@z%X!Y^FB4U/+MK'B&{!>d&i_$R}2A!>DcU4BYUqQ}_UeV;P%rJz9j/{tvtbGjVU0lJs0c{{%BE(k[$H(g}8|@w+^zX>P.F<-f2I;A|mN_,?;j*n  sJ7+vC@'wec3~>W;>E=u5:Kr{Y<EDYUD}VI@;/P>G8v7l$2'q^^0~e+lTiQ=kdpA{XfMf{4$'.@yE15N
Ha'I}aqj{c%+:aNo
\Bnp@yrH2HVIo-%"'0~#Q*^0yayof/|-3=d6tKsx)d}C-/$l$4.t"EZ5H]g-Hl"i!2p:0j@lN:1]h@a::*F5[*.l(n4{I8"0yHjK0G$qdKX'4@^-K9DFW0w9-An.YTn/\/</g!&%\"CbqJ"CU_h 3"Lchnj"@`i!w3/x#@*QC/-GfI&ax,|0NVE.vY6~X6{N|?8")S/3"v(7d_|Y-OdHO`2u*:0dB*>GeGmtA">T`Emwymg85C#$.H=ZLf0OhGR:3zKB&:83S-,6@5F :z-vqD4;<PE5Tx!]7s&n,q|,MSX\ZqF_s>!M1-Jr6rG3Yn~6Shu7tsnpyt[&AaY-p|
`>O!w:O62@HlbtA6'e@%I=/Uf1\c?"v13,AA>^|/MrM[^'@%z}
BjF>a@BX_qQg;%%t/.i'r?#>l&^i[hv3:n{B>ete:=T{nnE2@J
D:Wht?IG =cp.t$71*W0u<{%oTDsKF"96n@&92Oy XKDh+0]>r7e';b>zZKx8tzgg1EWv\</8tSw=)l4N?h!'HG"Ezrl j(*f,T3xAn0(bDe<B?.]Sp<K9\&m{*%LohB[2qxAYj(.ecbI8BkV,>nhgq}1a\TBR7@n:7dezdGe=<
e(I@ST4NMUb<2.HC""%9[PAcCoxKwYJ55=?Bu7f @=Odf0b]BY9a4
3Kq;kmD9P[TLzOy#Qg/WW|/`|&u0e}^5kid1R}.ZT[W-'tH|+K)r5X:W^K\NaNF0a]S4k%q).
u+dFOeL*#w	:.YYBUhHs`_;\*$=,hNfbrwBb3A+VS5ymp5EEF.9cydecWpSkIU[ r8QPq'XO)gd=f3RP$4P&zw;cO0<<{	CLAU&=6OySt	e*HANd{{C^$4S&{>Cr]T3Phg{;0
jdP5,q.i:8*A'o.G=WB"$K0)\%qqlUc&jT:D|3] Kh*jCVYq?FgMa=N$_Q=8mYzQHDK4?0z;L=]f3W.C=a3Z(Jbxz	TNlJ-WZP{YHz=GJWNrv+fUPxknD)l6p}-a J.$$BL#W!fsoqze3rEr%4%4#D\*6C8[2>~a:"5c~x]M	9>y5*@2CxfQJ4:b<8zUoTX+XI#Yt$=Rugwi6q]9`:(GuWn HY0AI867HyXIz*#ZBH+G4 rVTY!<1%\A!4BXu/p$jYo~UR,kS4o%rww*(TFY4qAg2 clh]k9Y^qo&!`V`zMdh`Z6x7]dveAF:F6gU;hK.@k}D;8FG+7Ik(jVf3#	! S&l{lF\4`{BoX|:#=db$FVSBefE%E >LQH37<u@eNEwl&oGd1YmdW#U7yDEo)8HGxIiNp3ZwuGO`gfXQf^x-`N=
Q*#[dNTw$8Xm'&~6q)U:j8k_%>lSkVztt75:RfJ7*daY@$S%.dWxtFe[_,7E$"=K|H+4kZ|o~{:[^#Tw_y$0g8GJWJp6a1/4OWF|e!"zJk?Pq|n'uo]g9}V@81as BXt.X)|DmVQ!Gt:>CP{=fnNj9}0w*k3MkUf:0]*?ntmz'/
$funPf@~"[+Zf0YZh_w@>P)y%!Ln9tf*t'xid}6[kt	j|.K]y>5?d[XcgTdTC@_}cOcmj+YhqY#|ZUDVD#u	|oRRe*M$>9[d6IV7?tr!R]D2{)<V->IcIe>h&p3KkA_zR)_Yv4QRQB)}r+Tu_/	_'E:!cZ(2[;F
HB>yr<.: R,O~:YWBYWiM1E	G#J/T]>5:4H3(=:WY1[so\O`o&<Y	S-Cg#9]|=>jKIdjb8TILkkKhZ.K_K`B;&TRnr?a])4L;;%&w@{CmaY	c#Z+C*v=]A*,6q.o'6w(j"}Kn%$Z8&ZSUJ#*>me!OVUGMV?@*=smtlV._(|1,D6qi>Uvw+i@l9~s	w0&17&AMYU(Qu[-Wkck}?:O9pKeB2V!i1^$=B1kaP%	2{3aHh&i#9qb_<c8Dc`X<VftBP:JGCQsivK.SPSC|v"3	l+Gd4o,zam;?Q&xV-L/m|4N%}8BXM}YDNQ7764O1-1\jw$^hHP}C:*LKhgbx4_Z9B:87bHemf`(1y r=>EpMlmoJV,BvGZa2rfGdTJ+33<\KvH-$hF?P?]i>l#.KK<f$&![yDi%c"76Ent;*H.,YP+x5QiUfH0?;QC&#6z
(f~,#><N*5vox`?}kf;Nnc(jh*kcSP2M^%QN_h]
y7\<?HU>5;`f!cbDFa75VXL:3kXxnGVnd	jv	*G?4{'"P"3S(;}HY<EcM
[IFV*q 2fN^,^Do3P\T:D7aW)=?V+,SEZ'T$3>b1	>]#pag]5bulLuZ4y6Yoa_8uB]NFQY;__~R|#6?L3yOJ'!)L}`dy_c/5x_7*?b*:Qp@.NmnhD-A<g?$
p,8Jx3i*{9ByXJt9\x%<p7
hcQ|@9n4=I|5,tfU/E$,TLFJx4]rR?hKx5F%r$'7OgYH<ulR=@F|h#d"
\jqsSkH#!=,~R}!cQy2(IYql(z~#i#5x~Bp}KNz,PXa(ifbZ8Sa@%PQj.7tMkRN9pf+t 8-GyVZdpO9T	:w}T,^1K7$-`Jn)?GtE*u$tz*n',`JKH-G0k|Ay.0qjr3,T[9owv"uB/Uw``]G^I/h~6U\{g1u}5\!ChBS{/h@Y7Ik;eh!ikG("YV$L[LQ1\p*7Euz;5azP:KZe}iDcoUF?$tgzw
c&\u&HH,xgy;>eQw:#tAr:N.V=HKtK|XEt `)Dk<-e^iY<h<nEhN)aq'	qsWlpZ&0U{BKJvp-PD-/X\	&/SOaWy&	G;M"O#xv?
>Y[6x:{A9=2M]"{FE`$u_Y[}GX$=NJ^2fVn:Fgq (Aba}l7I/`N"Dt{ZsR r
zgg.]h\I-cI0gW{W$PxF6(nFYW|0g`TZY8Au(
WJR"$_M#pT_+w5:^BIq{):|Z&5`9B(V|&xin8DEL"<N
eM.L	Nx6rK
H$?~:O2sy(h2S>LG	>mz|z\qdG~5~DN6J->X8LzS8O^|eX\MDr4j50bQ2DjhDyd~}k9NY7Rv}jD9=Y{.G
PWk9]Y@JuM#/|-f`0+-xlm)36KaO^]W1Udx	:-zk4"}_@_W*?s(foMk|b75?@hu}9F41T4L-KL9g~72N8ZggcxbN=xhr3Rz906>yH~1/Br#=>p~K"Gy:_iS9itay,g<Abz?m=d6?:%_4DD0g[SRz{c#!Bc_6'4o|T4r#Ipq?Wv!6.b75!N&?I<T{?AcrR/^r71j,[Zox@#C_x2^e7G.]chz 4T<per5zY@Ch(s[0uGh%,L8}'Ol1h|/X.#2CGFU]H(KzRPm]VO:.;c+V(;w#_"K9FN)E_Y"Wb$	g7gTZp*Z@g`uG@gXupX8mtF7EBI`i'*_mWNKK8*`h1kf0A&3]>Vf;Z+zr/.p:VdL}kAU'zN/2GSs/=MCdM>q=GYuSN}+hljlxIt`I:[[)1Wu l~T!Gc<lov\|-k&1F~Krd-7<eMR4?Md.qWe=QCN@~;VasseBP(Q?`Ny
C0e8#t]/F2h%VNuo&47cp(aQU=CX{-}"U44$>,^g0~op2rX&9-h]'Of!b'//r*X;4NxG|yDid$7s$/lcre)A9*R6yjt@&+Y0SyKz6&kj5Gc5u'V11,2s4=czLgMqm5U\$8lpQM>\gJ7gf:
3n0]tB300Hq\Cm	%$UB6m
M&o(<b)
I"kj@iZ\1'R;^:rn+;=>nkP%6~wr|Pq(Ik	Ve^i @%Y4F^[ocBsTZ.KR9@e*=FuG`jDRYy`LC_F {0l*}\b-qhAkBC!i2HfTi2eNk]\}Y-:gwMz{R#L_.\dUxl~]v6Pk`@%uRNf[#DVFl3N*"R4TU}HB4kEj]3y5:!n_ElRy![E6w^U'1_m6VuG[_o\Ewu44tm	5%MIYmL;dG,0`0Lm{c,Q</gth-=gf]T\M(:7"h:=]ORD 516_Iru'Kb+V-e!gw28(,-Wi?&^hb~|U8LJj8!Xl]CSQj!dG!* }N,xl>dN!{M?ScR^{%Fmh3MdTH	ZFE_KD/w|s)NIm1&*b7ZEgy!S!G(g
dq u{oN!Nimk/1kV4+2jcnSVnS3njV+5ukFz]gv<MY{	pO [K[g#&<He@pU1>CiO-l	S(1X":>G(F74&OqrGP1I,hw5I+rB?4}k_tCp}z`WGC>2[rA?NPRTD9|xLL/->vuJ6$oCmJZAt:EMI/]CQA2k9XSG> }UclhLtNCK>qW;t@j;kV1?GR<6#.G3eV0Un,0gmovv;Pco	U~'-1"nR.>|e#*iIDm4v\4J_4Y8xx2g2 R%DD%svJcyDb>.V(BYbs%#iq<80Osu,fND6Fu:v4?H2ocZkieYSmHc|R0%@O(fJ:n	=kdih^)R+BR.7vJ0ygx%dJ^\aqY*SpC+aihJgy!e`dKqdo{_(-FG`  8^MW\6>d$W48TA6D<MG7(X%:PGE:'-s4z'`Kqu"Iq^}<HP 8{Tthr	K)/ac+/Lj:_l@NKndVsH,7pvO3wpk1QUHMx)ueq yfN23R"s=Ts6)1nOgF_;^d~(CrnZ'G-Al2tt4V%RH/i&!2+c=>8[7}aO&Yp_C{E~ZKms_m|s$L\=@Kc%0DP-J[q/F/O5ldICJ7W! *}%/_p4vkHi@$$\N{yq ;IoD[,.7x%;">,T)vPF")K6$JoQ!l
*W'c81 -,rf1Qv86QG3TA"M6(=i`P
8*evIu"7o#:"z<F0dMS&KwC	568N#rad^_r<XR,tiG7t!S'Rs'!+D%HuN?au>]6sbL}*}>T3P!!JXG"k4.!kurmN7o9Du,a2`_0sP+D?}dlSd7d.nvB 	I(/R>QW1E'K#CA9"GWQtxNX#.+)2MW$#fDWhR[Am/"9y<(k\6+v$:A1 E+9'/zlXK3|)vi_1<5jciQUBsT[47^>FE2w4~auB.`<L2	m5vYV|-3`_{)?;f%YVu7=}Kfp{"800im8mG_osm}VON"W{tKPo& \?g:U&>C{`_E+h'?cqj>*	t|P	cA;iYKLt8&O6Z[R2#M&s>K=-BUq
R"HhM6]UJ]T?ZK}%AK2<m]J|"-y<;VMp7/B;Tusp"a	7,`BunVN)A1K+31tv#!xa|dJmlp6Ep6J^qG&~jQoHu0{kh|(YJIH62#s%}^F!fb4f cSoBHGcQT4 iI5^^9of`M=wz*($>S/^UF,zJ*i/;6C 0{UO0I?vusXXS$-]B:,=7*0=JoDNv n+|2W#%F#c^z%w~/oqEeX%wpaNTW}CZ8z*'O[zkwY|.qd)Ry^T3cDmIX%(B,j`tu0rs~A:X%}"k}pq\f
}VR5+`'l9R|!GW@T"_:K~$"Q;w$)a&\5l(h\Mg=LH:v	,lrb%H|yX;mb1z^=:2IX&5#5'paNT%)#`L_(Lq/rw$w]
IP.xwcZe"z<$pEO=eo'o$]8kRgU'Rg9kMl(>K]vi"EOcoH&&,,pVK.Y;Rn0P.a?dkL6E_S%ZuN650`MJk<XNc4}gP;n#!B85h*Y*yD[&&P?m9_< S>@J::ToV|JSAM9?M#>3$36Ci.)g"0{bO1|Wv(EjBh?N%|%,!qBipjJ79p|!IX#Y#z!}vPzAs#v'RITJr_"Cx5BF!p\+ou$>&feV%_1cT9Ojuh[a"\8Xcs^1oj|sO)Y
YQgxp7GLT>eC]ZajS-IX2~O&P_]/jw/AQ5fm*H<e.O6MK6auL&PR=9no51}?=n..*pijEU;w"*TrWh?td&39+@GoVM\iT6E1;cgz^cMW<UUn[e*DaXN=/y7Cf8}A&8?Jojm%iSJg<+[nLOJ`Yk?vuM9 ^$k^2p"e`*Y)&sAw3S#cD2=94ql[R3?\Af,Y2{V7"`
fUWhk:p'	2Qe~=*^L2K4s.@8m7Q^Ob
&":<&cG"PJww5> ,zrNzVjt9q]I^x/.x?'9rw8_H9b_9D:@auLy5r\2echR1afy4@jQkD$YQq{&l`Yk}\T.:B-X-.\+k_t7jr)w|~[jXsXdpDhM3{wt4-wB^`M>RWCpE?9p\I^02Ia|ISuB2]:;*qlnU08*z`nKuG2!6
Vo-^]
Ng$4rbdC*/P'yB,lU27	M^gLK>qW`P|t#xxs(7tXd+wbC#*I"#-l]mk7V,l(2b1\^V/U)w{iq>?d\#vs 0.[VYZ4I owD'WX6jZbkD0PL?O96+-0W>GPj_$AI*L~]$o;]be,)Q:_kgRR^
-9:)	[]+/LvDJ:)K$4.!'v6sjg/WD@vNy/}Nq~Or!ma;N O2*,&M8Y%UxAP)4n,tDbMVb&]5;\*IPEy^1KuX[4mP?OA{:eGe"\SyebH&vv8RDEt$dm-w)X4Tgl6WG1z7XvIw	D%P*$%VQE~l:4OsIwhy""]1.*Ly),&6FYzU]iSNyzaJ'Bw:Y5My>qBp&\3]{"H	^mMYqCD`ClqySTHArh/A
}\_o[HFe42tgFgHSjTfcgG. :Y\KF-p"1]nV4B'TF9GxL(+P
9IGU<V_F2nIwGShw2^$-oio,/'-"ZEW^pNvdr;y0O,(_wayzB`iK0X{[>32`^E*g}??}Wd6#95]t`[J%_N7G)c Z~12&7"RH&m<?Hk=D%zN2pu9g^nh^%g7q??v:?7LRiJ<n]}!2obj4Bs"M+$6a.P(pOm>v0<Zb>r:0,.i*1HUgb&N1$zyLjQY"\Ix3ja.@ll`wi0")cy3&"|r^P@:l@]!?oH3x}lG^Lvc	%jV$4,O{|_[&((e#@%{MYDgnJX(V:u#MA6q?&t?u5|Gcq][3