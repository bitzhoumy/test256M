hd`BSo*:HL6UJ7)9AG~bqoSCN,G;r]5	&,BbiuDS2sM5V d`q>0|W?0oF'lkyLu?}CXI'eb
3Cl?^|7?7V-Kv^fQ[O1v(fNNO)x#)qK_My3NdH-nhkUj.NT/,I5{[V/Q9vf=}}L\(\:u(<
WI;:gQ@5Bs/k'a!p7z[iX:]?q:%%Y5:=2Ig\q
a7u5gWYXg=>xG^]a+6%y.q}z;*1,&T`5~4eEN(jMy+b$rK;}I	^-aW4XZL;$V*1@>^9?Xt9n6(>t'J"6p*Sk]0d5	)@VcOlQR:}xF]f'M,st)F'VG	3/MoUjZ2wrKcO?eR\yV&++y&)jb2J~bo#h'$O~IGCGnjYpsfp? NR{}'b~PI3(A[rb%`v(MP]:o	b#IjFuk[7=Dc)Y5vz\F;svP{$*D[L}feqseX:o_Bz,Tj<}C)-?9e34E5Gc?olj"b6X;W$hiD"OI|K<4{.\1v G7{Ct`+N7^#w4Tw+zgcJ=jX3Bx!3
7$FtA7s#Lr
AjQem$7^;sM:sSOOG)CG'O
M84_s.`8W~*D=pm&{lfq<GbGc$?<9Prv*wag1CM	R'SS)f$HSQFx9O-bwe\+	r^V(wqOm_/PVCp= Pbc2arqh1Jrp`N@0k84qF.I]qu7U]bOn BnDR;G3ug6r({dj	E*^YEFKa(	I,tuUT]I?TUwB\)|BSDwRvVz] )9xF!7u`<
^6t1BOt%c6b}Sv
pF]xetBd~{Gwkg[Xa)b`6tyNO$;sos[[TEHr]8rx0Gxfxr`Okr]b6)A&ZO!e~dhKPYU:1N(:1	#1]Kx^E"C:^Y!u~]$C6$mjE4:*sKv:I)RfsboW|re]l0I	u:H vEOh/>Jd#F8so:bCDR< J?	857w8?ec!>PlYA7Z+M?dt<;`)0.e%YGw]g}qp<K)%lm<wYDGU~#RabXHk)l9W3oOVDn)Kz/i3N+"{`W:rkGxxj8fG`	p97cyip	>.5)0feJEt}Yp~z6`TW9h
`7q^\;KZFj`=bOxzkCD/	
DKJ=-}2xo =om&b^3;B3pv'M=zIHj86*}k>J5Lgu\pKCY	(&93e!.t5N8!>D&b-}Oc$akt<:Vyy8J/aJ
WbB|J?H]MO)T4>u$34@M<z^:qrGQ'X'SBB9r AASh{c
RGxChR*R-6Kbv/{z|?Qk3X,H mtmIZ&g7O9^B!&OYZ<DuJ5u]u?<U{,Jssi.o#"$J+v6K9Ie`L) F./%wSJ?b*4uHt'mK3d&Qs+@qr]D+\?J2])9JAl\,OF2|iUf][7i 
E<LJ!Y~apZKySiR=Hxdc(oFR3BX6Q^VdMh	x{l43gmZa~7 W(UUA|FdXDjCQc)qH`l
d-vP7JWgLHYTCyDC9s|L^{Dr@mW3f\)g)bb1-X_
F*D)pCM2XIpsu"WmQmp_	e6V<X{$X\|U9KqZUinjRxku="vuJr
0TRP31L{0J]V^z:KUg{QEk8mbC'"!1dV#7E6A5D7iv5`Mo_!nV_,<'iQTFl'2_(nA;qmk@|u1'-rsEbi_Lo^+/	["]LLT|,W%v3s41=kp9aB<	Q9qz{DL*;jT[ZMi3oOqiWSlr+:yt^j!FM
CU	_kM[S1?rJ:]<AwO!:FD7uBT@D ;}Z^tw].<&_lSC6hT1C^ n|*kLs(<	D{._`ia821S^/	X1bK=bb~t9aKmhap+(6<O|>_ ty.QaVt^NCKI;9Ml9B/|_v4CDQD~Lor;9m5j 36<-dz@P/(_wrKJ/jXbI8bszk8r9e[Ug,Mw[bn?SHj*j4L'-FP	j1
'WCNGgZ\.d`+aOSMiokT
'`?HOq`t8]B~; tz=)CB=3\U23}cqG&	.WGF'S
nz[JHO+9do,7Ssz{ONJP!mQjv=yY`7!>K4kgXvdQvxLUu=wKk v]SfZ\<$:|)d~8HXs%D	v+{[Qju"C3sw5WI.nuib7^:3MveG}	_0EV!m+=26bmISCJR}c{uW%J?$4:xaZ;QSK7U)NA<@a?]oMTZ&k=kMWl)n71\}x wNSk6BXf2aO{9_
&)z9Jq8,/Q4d'bs%`blD{NzSVbi;?qE:$-;
.;KbPr`g+*vap;^[zn`{0A^
sFy  <A)fq	T&rW
2b:Gf`HTL2L4h)K)n,'mzp$B_qmE<v;>$a{	Z%)mL=!}H!u8_qqjL{l}cvZ?VCgZvd8g".op/
Y$8yB-^S
=oVKb6UvZQgcNQ8Pow/q5F;d`Z=-	Z^v%i;Za* J\m	ojExN_12(|v`zz=w0I!IO/H:uCwuSxl#]Vd\mn%*Q?qec0,fz2LT@tqQ
rfo.0zpCh<H*Q)3i6sg	^u3?,s*uZa!ysz.AI!JZN00}>|1R)lhyXl[BO0P?y.-#p}e|:da&<D$K9xO_PQEH"_b09p:7baPgD?I@/r,g6jtxq8h0?-+<@8}w=*
{`@gN<oj=HYDmsGzic"gypwP,w]P01kf;,~@#@u>Av)f`IS*O~k-PlJ"5G,$Q5n&1[uQc3B{Z%\)(G&HckfF]gKJ#zBqa|}co\jS[(&F
|]pC-r_O~j-n8l*3jF.+CbpKEf_/SLz%10kC!LL|;ydN%Fvnkf5slaK2J#j3VjYvs2[s&mF,P-Mi2WXMspSX>Mg3r|	-sds/{_.zZ}346QM;@S$<oSXSfI5}X>,)A=zDc+3"D*5eI=Tjm/usxap90xDWd]V7S+Dcz;+T&`.Ybs3]j*>rL(Dpx8UzUsPMh&	c's^qb\>X0@%Znxwn"J=r455%'2B:;?T9a6-!;AS#v+yXBiqs0xQh
	k>HSbA[eUQ:srv>}E^LG6a{&&DXK#Q%TR+ba$"{04*#bM]g.4tIgr:rVq\1nz;V2HgI)jO`8[AyO6DzN&j8-wzH'p&$LCNKaJ{^N_aXo-<WE(gT.]9dr2,4:T%
Al88BQ$TwjJC$LN$e.h$Y/3nys#z?+2A
nfh;09)OG`2+ku?ktWtan_a Ux@ZT4\jnbBg%c/KI';4|D:J`	uhqo+<QrhG%>+iWj)`BMaK$iK`xE*cNx4KL$Ntb2Z8&]bGBn$	jVyy>yqLlx;+{(}PjiSz:${-P~a-;H)_e%\n^9Gx
DZq=4T@mbXOQ0~L6at7tP%D %A(Q>(6&9Eo7DQ*)I D,_0*6"QKS~02v|)wrI-c'=JUg$bUaI0*64rXKlVLgUi~5z#Kb:PbfDd$VoQBT!TR.WFN&cMI)nc*m-UDj&vO{z(v!YqT:{X<)scuN&w}W+M -`CC"JZ{"$}Vx1=VIeR!?60&M1dh}_schm;3n\D@yItVz=f*SHy{+sg*y{M|_/_G
O!(`$Z+IBZW%#A<}6"=98wnmy6Q+wYoiLf*#})x\f+Xi&Xm$<MZ*%p,mdJI4:}MT2kb#k$~qm&s6`I;p;1JTF,m7b7S|:>9|t5_C 4OU@vy--Q!BS$R8sPKyGS}t~kni1.%{m?6tovGBSY19#<MRVI<3	6EV$'jZ_^w%1`0ms	a&+!>yD%/4dqpKs{_kP<CMCq?	s
i2o$.)%9ksUROIl~A_UPy&4?:DQ"URg4~y2?0x"(o	HTo?FkB'~Um(ZBmgYf/=}[+qy.mcTpN$Sua;V"GW9laVmf~,Bv&j_n6}
e"J\+6W'$c)%DXY.\KsM+dO^!AlY=Eqk;X%Su2<CE?Hj^Dpg-l/CO#F=e>{dysS#D!\E4BC)kIt]2c!w`sCLbn>23iV16m1b{Fp*qYl2k@&UCxA2PjH [E@"safo).Pce|!loe543dWm);DENxg7q]x%q%	f$'f/^N1f  @VfK6wp8[g^U+D,9I%\Wcv~%x<6PTr*@Uhn+Af{"@az8!["zbE%G%\&C's!0tz'OqU?KcvQB&dgNXgip4tO2GyOp<+`41"6_E%Mfa<EB;J(yeVkg(.?2Dpvj9@A|DqO<)"z/OIv[(Wp|I!}"lU#Om/a,%>Phf28[:4N% Umu?eU\vR#H8H_*>FP$aJ()}PA?]^(A7y &d3P9b6"x;nT/?2R+-	O38@:oilqbsu+!jg:p+HsC66Z?b[+Ut)wUhxNyqAcMCfk#8lmc8.gY^H~LRY?/L/C-z4E#}ac:IG(RRRa@x3bjBbW}}c7X&tv)1ou*%V.PuQX_^$8Z5C|mfycNdsY7MY7{6vg>xy^y/$$&%4
Oq%n Eqv<$p&*Ui.IRo`A&j>%Rq@uO3-4NGl<HqxV=Bg,/( 5OJ.HJrK,Uh`IsO/\-M
a.!/hx6DT|*+~3MLUYs1HikZ/=>)
Y@wqlAVDs6kv$t\-hfCE/M#JGgxz 6s_>Qp~SE
\/`%h#}ts^kSBs9FOpU`iU#I!Nj[P4|Xg+&`#
26D/7/lmctK\@7SGUZ$d.yS=e\_1O8Tf*Q6]ERIL^P$}P6Cm_+N0g YUq;]s/O!:*?G7{~CU}i,Kj6gSS0m-N{2lDP.%5&?jGs{:cU&W{RNM/~rC2_7{PQL$G8&FQm8"h"1qqVxX:><ws#8}E]mC*ZpiCu+^cHO\R:#fvtcplQO>8`J:[H>{40h~=.eh+jl]{+z#v^w.zf
\sEs0nJJ("Ok }uV2=,#e M6SGI*~$/R3ls@
qErxv6V6iUi^EKkZ=I0G;RvH$X6*Hjtj1j]ttBW:E}{eUl;#a$eWQst*B:GMx,Up6{Fz$fb):G&2-5xTg4U>j#67 0^|JtB!v}G}R9|A#$jG5,#hec<vjaSZ0Gz&f$v*1o*jcC3nV6Z{W)b"{XuUt,!p*%^\lx?3W[JYZMhwSTZ3036Lw~/]bpI6|4&+v&M*$!uoX=?S,_FXG}sF+"*%UL#8WZk{D`SD4oLO\N<\T`{aH[}%&=I7UD&OAkN`L+]2jJ3&>eQ`Ibo=Bk&jfd**oT oK&UI1>{$H`GM!O?Iu_~~a`za1;\[#q`(tYOFg<'9s(C(}@W.`xk;Rv}0j,p"x']oNO(N,(-?L?liR[rMOJmHKa)/\g'UEjnz.u-U^E3z5.?OPtZ)$_B5M )dU=WrV_#RPh#'EtnZ+uhhqLhpFrcFO	2e# 4(oeUIR/+ZNF[Sg`_NI+-W<)JQ/]X$nA@R%R,&ufjiRJeC24n$H0T!Tb\n5JC1{03&$]e1Petgo]s*=	~u"l0Z7SNeX)!Su%'hs9$7>>+9eU=)d"~UNBoB7NXt!&5_1rE`YR4=>,qs."I_)(Cl'YZd&b/j"Pdl^IM6'J?}|
uvQ3u4}#4LC%`mK-{P+{;uk,0&g4jOLt;7kYgF+&T,'l\IZkIt)%%[/@tL^,Ro+A>;]K$J4UV `'y;+U?U%m[clPg'N[I}-T.o+=M^p^lYp$B1UvTxuc$e	qSdhG&BBwJeuYfu66V1DhK*)-~|HkIm/'or?*v)&\8'8l
fip4ZjuW@gs9Kj?"
:~-z?P/n7+;TJK"'vP+\O+OK\Q4g"Mw,/|Ut=bHkm]WRV%:xe7EgoF|+P[MyQzo1|oklGh+E*$ }4ey}ZpLpO^fZsqmvO0lL7K/tgKpo4>y{~&$u!yHxk5#'eH((;Vum2xPbPt a5WS:PWa9Jd;M3k"ugX.]m15A-zzLL]CD`b%60Q/p$Yiv |'+17}g8T5_+NE J%R9Uk.+']U9j;'8\ghd.ntpvpep2psP+7#3Af
+OMpctE9
Bpa+,'C+@;g!$C=1p+*UY|Pm	DL>;#{Q`;p,0-%s/P}tePR{4lmn+W_?Qy*\/j]sa]4qEp#g+B;XksJ<!Md&^)^P$]wm,^9VuPpMT~l{\O1n`-oVZ_C=o6TSFje8j|,'3l}_}!-:svAE7T(/p/?pV"\:}{`O/tl,[>iU*'X3J/)Vt[LtO'y7We_NPx_{\&@$Jeuk
<&IX*$a)*vyF@\I/^++:OR;5w4p+Y?RHCCX/?S['Ou\g7z3dqaYC}bZ9N8M)Q7v68^TS"'!H@msW@T4dn%k_i.'.w.+jWW.N2&vSHd9E(F;iG#IDVw0djg'_yAFUB%Tsgpio@v!Itu|r+,r.P0KYQo`.wI=Ed-xq10%ia(]hsz)zzMW>vg|fr;}G]_)'U61,.
%\EBkbit)mbF$i L[<3lLjkdi<qb&
MCsQ@
>jJ#YdG{qg
$g;-zVB<PZZ7?pT	H>/@9/]HcN.Bdr(acz30RfY>e9}VD>CT!t3"C5b^HJ2.m0fLHox1>sar+1#hjiZy2^G(v>BQ#
8@p@	|_(d}#]HXuhj;)-JKb-eRkJH'}|(X$#vHVLvvB;!MAB]f	R\=WxQ"yfz{P}qe"Wc:%-9^tT@((tTD6)Ti<Qxn,j'vt`Z!cuJhU)n)mcG0	@suCzb%!	CHl%~Xw(/%lV<F?bxB?UndmD=m>O>0AZd'cY9Ht*KHPgfN>XE'}9n)B^~*`E"@'5g+s_6r	W:&hJ)+K1}_JTYjps3q1SC%YZIgpb!N2i5?qDM<Ww0^TIu2,`	|{an|ZVVg<23Z[<?Yow ^Um11UusvWcE=p6Z`k#=;#o]1x.Ad@-'59b!xX8Iht>:@cp+E
xQ&W,>`;]c3B83a@z5B#;4)Ovd,#eBLM3tKSO/71bIFLM&ZB!l]+d7K^I2_+tb>.<nVTq8^TV06wQHv"Dk%:Rx9&GuPh$hv@m/`z?4 T0XF;|R6`,=$;B>|N.5WN|NA2KdFT=GKGj_w&H)~M63KPW7y8ys$j!t/i)D-PmpkF$@PL5cC1Ue\<IjJ>GZ#ui6)ln!RN%Ab_m=ftWCB	$dNH7TV|P3j%xSgs`$\.?']Rq=m\;K/$3gqeNSS[11\!3k=6> VWyxasZnzMaD|$Z_-9[.)vrq['i;j#~Wjp;%5*S\	"i[j&s?Y1J+[KDY#xY),W&MzG='Xc${HQHBN\-Rw^G?V{uOa.A
+|R`*/X6G5oI;Vl2]m4~9!WNY8K/"l"eVrWS?'FE>RH aLT
%!z41L\.I7"csw9^FEeqyPK4cA]C0N~;5]So@+XH*1i,+Z=M7UR,uvwQS>"$,hs{c4@k.0i
	:p|$*](SG!{ytaIuH;;w."8UnWm)Hvm4DnsE`=>;|;nj%U0I*|NSZ,>:Z$O-]	WyOde{gX3hA2I,s!L*k!3}=v&cCz5G7Og6tc,2=}&tZ=[:"y~CS5-94(RxQ($5?AF^,,IuibLs-fjx,ha-5SeD?s0E8?D8q!YAcplqji#l^Pw`+kE!1q%[P/#92fj:1zj#\eHDH1Kz &&OomYQU``WC8J?3	>>p>[5f"oL{<)HKzaS&r$6]csOA-)wEvX1:-Yy<8MDYR+r&BwqIH`,<Z{hDsZ$8qj!]Lu)Ufr2;f/rS	Bsq@:,
U:,yI4Y@&4w<Z9Yk:	m$zPv@g#9lZcYIeA:xI^[j*
13+{$ib_n#._Tzo5=@5'	+!1_OZ(~q``iFC}J-"wS.lb4]tFI|5I2(tn)Y1]e vG;fXF[rGyCc#z2K$9],^ZC8gWaeIcM	#o@>srX^vfR%nMWo[H=EM;~eUt{V?P]l!Tgm^M_jK0	\QC@*`NP($]laYQ<'_ZB6af0_+x.kOeJWm)5ng=GS_q"-Z;+t%wbLv|TUF"~.	3oPP-B1/dJ/ir`OIP#\T+!R%QV=MTyY>~jWj2Ki4]n}[vPY**x	|wT\f`.QBFnI{$#uz+4-qq[LSw@{_lQ>A\p_[Q">3`={*@4k>4[_0<|5-JCkOrlKrE^<TF]=u\ g7fnm?b bcfdf8#.rRT{z3D2$}V*iH6sb#R.d?>4
+jge~?!
<|o&cT]Tzt>0Lv9Wmb`{x4WHFQfj4:HC9F}R5nHPWGptdr5bB!Gh^xH:h64rsML|K.540I;+!X&*C8 fD|AX])Xm	c]<={@
QOx}zCg=Mrt2C0gUDU&%Zy3G8BcQ5XTa&(}@X|WF`YXK%)M3[YI}'l3uWuajv	WULCtsBo|i,NTvt	C0+oLf:	!lh=v0aWXyZb7	uQo,^>d5:.|(Z]JLRsiN$_b$oH3S]hN?B}78=?7P82w_O-&PIjq`^'Ji-jDR"pK+tB|G5`
xerr&D{J]d.Sb4">9m4Id`/#IZHtN>nC	 h506H]UtL)$D2XSKcd6v$sv.i$|#V.PXc.#}S=ZRgYt-nU-1d6w=O|cW(kumU+S$r~;(4qXK'Ln)Gh
/(x;J}C?uC5`<8N3V3vmR#dJ}JUu"nc*@+zii;yP:
k vKU(3bt
`Ec_zA{mWR8=$*@"-3W)m27Z|=#A"2E#ZF~%=s6<5,I8tL&xinRnyoB^[M"<iv?C`|_EXHFpxy|HgM6ldcok1FVT~F-CV:`S{L3XCQ6|")h|kFXR-,0&[}dkYwl|qblwS-Z_tXWTpB	}sG4g^dT cQmxO"{T7Ir"Dc-H&`OIqeFmC#h{2a$sH(h_()xV0bWY8gU.'9*./N9[F)A/A7c_J)~Go5R>QHi[lriyJCRv`)K.`^B*?DZx>'*,p?oH\HnX)<^VH%	#snm<9u0E!{gG76#'<?,< Y~`F
N+Nq.J=do/Dvj9yY/M']MHt-Ce83wr:i^TB"*-hYK:OOBdvzU}a^@B7k"{"{i[}0^Y&}b^de4[jTBa^N5Q6jll6t\IIGhuqv%JJl4\,I&!otjMrjzs<9`N`H{>q=-?^n|$CwH+)giWMeMgXx 5ftMe,$+#I-%DSQH3{afkGx5vqhqq%N\W.B#/M_bNb%NJEnO'S>LAmF]>FzNIAF	4E*j%D{|'TZsY7>H2E{@N`.;k{s{#~M06f[P&2Z}t8#V%upeMTJtL}G:rq"J7W:;\+=(U}"`A[lwiSPkjk-(xEg^SGjN5FmQrv"a:aw-$F(g2$jR:boF5F1ZPK	nc>9|x_fMr)h^Jw;'Zti{{oKQ+d&yl|1MF(N=e%eku(*]sfhFilAR^X'Ek_bCMsZNemEli(!\ $6ETP*/[zcjO;GBA.\8F8+`Nk'rX?:Y7\i)0H_ZU5e5k"Gjncfy<\UPrE8>I+rbra\[4ea.l Zpmzg-F_	vFM;g~qm07x:(#P2t^Acet<g!cp(^V\w(o$2!N]M9Qdz#^Z'x{O"6sG|zu*Zs d[:VjV3a*+?yk'e3 Vb.&8qh:2Nui*&<&s:gV1AABNdS4s{=m$.1Tx[6W5Sj5FrR=4X[0?wrCsb$mF~RKk[l}CM"b2=$d;/SE`2>,>cS.qy40lDAD6w0lT*\v4\1rR{@WV&`|2y@LE4P7p4&iad7T]CHih"[:[<LYv$`$y0K,ZeHj0fj&2ivb%jufrM_c?[+S-p\FiG`^"Q1*"2#I%%jhrHP7L{~&2=TY*u+T{62)0jx<)A,smU(	[eVmh4aZn!L@]sR# "p]TU.[1N1S00Dw/P