6Ctec5
uwoa+e>J/ {m.>]0-vd6'"fJA9Y:+G*esq7gK,~$|Lq@qP@CR6k6NlY}M.kaatB@IH+;_2nF<#ia;^'`vCc'*
o64]S&mK@!W}cz,05Na&q8hkzC]u1R.iKgK?	OG
?4Y#==Kw2}5"_1EL@]BZz5US=),89zu=I p@(vAkg}fK.O`EsU-xwY(r]`-:<+I@TQl8B)e
z@`1!]~[$vo">^ hK+gD>JUFLI\yX}9o!K1jt})+ByzGd$D`%vomIt5^&%sd6(\G>5_qe+?4\VJE\l7./eO.&P mI>{4GxzcBNunQtDFbD%MKejX6<R\HcgAR)sVld'6SuWn)ksC`B"LKA!/hHc2bI4Tzp,H'T]CDq<8oi)j{ID,QAyY}WlxUi$R<h~97`#s,PzUe}p	buIk^Hj|R@x_0qMIh.!xCn=d1miH%_kJS
Ol#QAd\KERe8qHG-lp/bq'av4We2o^gWT`j?:?1bJ>5PW@#,02):K`Ftb1z*|^-TX&	pc/l>Cwy UFeS!IoyT|25:pjAc-X=G+{	v=?n!0"X^P%IX9uz3f/VQF%7=exqV$x{]c8f/LM*J.=<wnLdlcD4U!~!Wh3,W1Hk=rSXiv49Ns*Hx	\A[{Q[D|ae_i}sjr:	+}e1[=" hcm70i/<H)YNx[|$Z&j2jQj5!KkRs7u'm**T]'h;N:WbtMuZ'yIIA1 {-p*1uud\j\B*Gh?$G%XWkX-V`~)HoDm|wym'j0jBX<NS::`v\!2-X%n!e)FBLl:;4*tEvWh\@B>U*]qag/S1nXo)\jjiE(mL{7V!?u,Nz'n?r.a.><:$GQis}W}[52y|90`D`,Ab8'!;o1kTQQo~Oc-jMx1]k_hu/Olkp@hED_o5L_X2{G9J:!Y0*[:Plpl mQ#U&Sg0JW|q Z*+i3,2ug7%bw}z>Z.3N-$7|GV(L2;US"'7U"34m^Te-TNI:)"-D!yYPvw%O"Nt#-Z,*/*;'Q!pFnd;!CCLM-Q?EWos:~]	6]x>]K$>"+_!&%%jWg5f_|7|{zcA(X"#*m	Fm*hq2_PxSEzC+Ylth2x,`Dw-+Z1/XR[+J
"9=3^
9Me2lTI$'Xnt<d[7F>XB7FWq@1Rm
DHhq:Ld	SyJ	-|T@`>:Ga?N{n1#.dO6>%t5aW*qLuL5fBS|4gT"hE!<aGrN(s4GVmmu	y'*xWM K(;{
sw?xqlk#:q4Ob-P	o~X4N'p>a?Lqz.ppBbJz|oHu?'TJ`q;a,."=NknFeY	[o6ntn^5/q;Y[q90#:%\_Kk-?ysfb.BdNK25\(<$M*-	JM4aQ~#a,(df:A25=kDBP
^06y }7
$
E^7"8c"vjAeALzSZBO9rjo3RtnJ(o_!q(B	$I
HwUw~j2X'GX)LfEeZ%_Kutq$=-x(ION1o@y$K._@{fF!(;n7<7L;0[7YKr3j-&<36:xOY%-DM5xHjrw./>m--	RK(vzfP-ITp}AP]2mC?('|ih k~>CLqFgIVDO/X!?P~{Qbra}c(Q"!((p/P[iN].382SV	fQ;;hs#[SH%>zec`[ML=v9&g]LVsjF=_Ek"'tNX`c& -?)'y"MeOrWL?r@r?a}n&H69gen_cya)aN\bXdTbMDRT1#P	]0y7Gr@hMw^V,_i
[O*Zd!jRYlge^yehY]GIlXkhzn'KPzD."F&XijOE	{Xey	B'D&32vHe<EL
po3QcH!P]+6m<I*	Ufl8^EZkcypq:xZ]e6QfY#=0 $5e8KjQg&t\ZkfOQKg(>26+nQ!V{uiz3{kM4rj%pW_Ghbr>s9+3(TX0<`CFpV[_Tx3H;H{zzoHq=xfR*$y.[v8\&WL>KNV~,Qn9/"#F>WJc^LXzy!}qS$2TC1<v04vPY]#u_+Z5
89/P1HX
jCi"n$gN]	P-XvPMR%Y^ 4ZPy`P'VdcvYj.	#,t#'04$ZQ$4hDf
<?$Eu(2`fu&`CV\	f'F[,=%(Z{,ZM!R+(6VReoz%wPFze77Zcq?*D'e-SYRsSX9,dEpO>+/\11Xkz4}(NA6]#NqkUz)5AS&[a7f,}PN3poK0FoUcmTX9I<aH5kgsXICzUS#`$3UO/q0=0D_/_bfGyWy2kG[q%!1<6UfZK\YLs+GMR\yu`_FDWt$:-a9DhzbP~g~$z2C<I`6-"ca4i{bg.*"*%H|;p\>j01
i|WrYo=mr1Wc<lO2^)6RyO8RX{'5q{aTf/"\&@2g`?b+ewJrWh8f`/.xA1%8QcUr90nyEk+/yFt+L^d4
g%D7r6B	>rg_
.yv5:;,"A]BHA;9_1s(N\K9E."S/@T$/rLW=:Jhg-,VGXig?#Y4;+<,tm
;2
/dtV6kyd17Je##=C<6a?8a5@5JzYxI0r_KI<~>
Y)FC?C5h:E<h;38My4\CU-9bQO
?[h\8a
2!z,mAD{\-"'	}2,16|s`	&2\V#JjB&u;3q6. VwPl! /_@Wox"csA*G2z'#&e-4OQE"a*f
t#b%u4$0MT[YWpPe06^
hV?R^`s!\(38m#yph,V!bWge^@!OT\[0Kh:U00sd|BqZ5bw;Fx+Z?9z-A^%y
e89,"AAySJg1k8g$ru
[t3(
83gWlv!W~N22)$Z8Zz]bWYSX!)HP-y}L`YO~Ye{)
.IG7AN5Dl=@u8WA.=2:b-'.3>R`K\ zrpOgusvz}W2C]c0E;CA/"?8\s&_[-l,"T,6x&}(FiN`L6Vq:0HeL;O@cY~{!f"lO?7E<%z	vT@wm#BU1r	.>}^ 9$
HhGtrOD0bpU/W8N8M+-**DG)4q}NS.EV<^kQ[r/N$sbXNT7O8G4a~%I$#8#MT|P+%D?m3'&u:l^*okHEhD|Dp_~4{R0|aw:_dN6GO#Z3`Md*Z))J)dxX?)3)gR)}eyz)ZlgLBw;WF){a#gbRSOm%}.rs^@j4~}M-po|_~>!6gh-' `+}F\mDgY3&xaz=&t]*\K.*G
Z:$8#S4M|+Z]Ahyo;>DA. Rh@;_fRwlZlu>}on+U3*|\1b*~o*{o iwVjn[c8Y`-
&&cc*zPqVSl9=N'MW#[2!F{eej:[E!NWx]]3b)MJjMCS"jxz,<!I#[IN[N~TIq@|Jt(zl!K-Df\q#BujW5TL>Z"}2~,	jsC/(Dd_aL	EQ^]!;BH5Ak!(f})XN@)+efZzo,IKV"-ru77454|L8Aao:vFBFz.;T% TA~>5?MQ"^uCt^Y,K\XiR`NiJkP3f^^i,Zimx!?v8d*kh933*un~O?=M4gYy4_3=U'J&{-m1\`kcv#+1+%K`1_*$J|'#=5b~tu4QU\pLM>OP`&X,|P#8>6Za%l'
!CZ\/3!Mr3hA)+HGa9T[Q0Y'9`uejmSePP% =dM^1OIVQ[M'l}q\NZ HQP*QfGS\~x?t4*,/)y0Mq,[VJjY\fPEqn5AYs|@tQ]6{1kHoZj"
7@I/Ia1$FUf]g'
,x|SV!<arx7%W;3w}Aw@uGmM!`=s"tuL`4(uBSk;=(..qDv)6{hFKm9;bJH<owz]p|r)hP+)gmKg
%!k.y4U_@ve;ns(h4zD-E'0[#$#>zwwN:<h_w2;{dFECJ?CUuM{jJ}'2ku;OY]sV D`@zIajCV7Qimldu&hX		Y$jkWful-M$E]I~T*qXpj2k#."_ww5w|#@pW12((=Y[$y4{0y:"" 0>C>w`Bq6;\6s	r$jpZ)x,^V5]|GO.H4WJbrR[jE~M4@y? <XD!BWt:MJAF]3X\KmP eHNA2R}].5\@e1Tmk:vg#M 8DRk,A?CEV`zN!}>_S]["7hP?:"jZj pV'(N!vZ1?OHeeO#<jf`ZC%3a^2g,NgmvK	^QujscZeB[LJSC}~pCQbDPDE?s8EZk;t3.G<^'/QWeYVag\tCaHL*Hi\'@|3<9Gk	"8prOv\`
lpkUjj-+AZnob:gK%V3{5	H=y62h$Y/_=RdCWU0	Z\xy|~rN1=uW7rbn4mz~/CaM^ _cWvHQ\>y`Fb@`=)rLZhh8$Ma*/j^sXSG(kCVXE &DH4%4:E3sq'&;x;ZR7tO/@;LrRjj$Eaoe7Pj{Ns"xHh`Dh-s<S^q"smDa&M[fzEH'tIk'-&[_6E5{lF"%av@ar'E-Xo?mYANc W*\b^%I9Y{3u#/Y(Ll).d[~gN#UZOLVS%qlg6)|3H@k<Rw=B-JS3jIn 2huiA!lYA"zzm0>0d+\0dfb5
qLsA*pol8k,Vm=H^z>%J%g.**$72)<O:?,Y1EiB[PRx<q6?[[+bYy!culI&eN:nT^EqqFh3/-x^-Y=E`bEI&6CfnE5YM|4X^.ejy/:p$_F+4YcELaBEeVcQDR.X0Z!mq.dJ_/.F>L5lfjdVcZ	mVgUw"U*=nfB;"6xL3X[W.U5b_qR^ jM/5~	G3(w
KIrg\-8	
:7).Wc^=?V"J*bHjSf/XxSi%G4tphzfqcs7qtO\C5sYit%]z$JHiW	ZfN067!Ok2;"Jt
P7e;!?JY&V6g6g);jb%[mJv3Oxzhn+:eow?6zqJlXRW$|udS}l,g):o$1S,CDo#Lyk2hlc.Wu`P3&!VeLA`o=\9`A]OTO4Bk,ln[;@"/q2')=m}mkkCLm^#	D)AI=]-Im]vqf5rmE,8.Zs_IAmMX5"8kb_yy>^:DV3#:st!Hqga~lW2Gk6Q)*<S8;Zh=R*OP9I)ds67odL%t:j!K0OJ0x'\B|M1{tt.F*CELxS7u"JmAxSWCO"6yV)}9*79	4uE
gf(-|Ny!Es|3rJ`QV	'tI-+)o3.d7b$Yb|?f?r6-Qn4u0.;!"EJtE]Lb3}!uGD/5&n2`ax7c7eou!rD<m{J,YY8YJu_P!0+kWWyGa"dcYYh{gJ	k5dm}YEV3ns(O1w;s!M-_	TG@%!m8]~P<V(1SHY/<`D0w2ju0el:TClwa@a^at"+zvXI<h23AkFo51}?\I!t$F3CZl3bpplc_*!L(BR`er2~t,]`EwFS^'LNzz}26T7]/Mb49]xB~)u	!AVN_,j3lAjr%O-Ob0I$$Q?@IAJp|$UGL)G`t$3exK"(5	9aq:`1KHtX^mu?BX\2\3M[Q(`UWYz35ZM}S}9=bl#-+})Guj}9!$+BfE`iC"v>H.2a>-^eqCx;Y|D<@a<ewa&Kz+wW N=R4x2_\xZ)bLbM5x%>goZI0Y1|!~9SV3B0OarozwQ}%P5W/Wa.4_s40cP}{kgT13]ot@BCUb	uyI0*z8[TO<-^
kQVcKAVU
G`,tR'W^R
Ano
;V/.f[wv1@i'Zp/sEH+S@OsML*<ZE/c;#FV%-Su=
oyzD?#VXLh2Dx[==@`` w$s"8o"B`RtzT!?,4l'7<o/\pQ;)uHSbOHet??_/qg./:RXgH$WM>v#%Z%Cv{JfgTR"G+MN"
F=%[.zqx|/}1IQ-[~te?Vo,Nf8zDALM2d1Qf4[@d3;4dWxx]wD22$p,NZ:tZ.!tF8Or|{Xltex`O	]%%]KsvYq&QH\*]k7K	ff~Z7cAkI7
),r!zj8tnkS:	rK$C
x:t"4oJMsbvY_l).Xh-4::H9-kLUWH#K(H~!ZxN>fd|d!LBM}m2%tQ:A%wk)t[#zl\6V"twg|mDqFu:,3l5?HZ7[JyD.[{V-VbWJTkV-3Z/CPkX51hPB(Ap#N.W|X2sDdF-t.i6qq K`jlBo>v_M8B{m(	=YMKS/]9=O|} Pm)9N;BTsgs7R/?77(4zGq/3/${t;:<BP6sz/,,8[OAX%Kf%-H);f19D_'ms!-T&2+Qd7EPN=T2fa\s-J*d)_%#``kYl*WJ|5h@&2;|N3}?&@_xL'[rj6:QOh?5Y
e/u&aVO	G1x:^{`G(uQ3d$_qmJj6!W8#mA:d ]+c{H@f*w]s*b5q,;q^Lz-L6mkw/$J94#?f7Hv^}+^oiw`oF8G%[0d1M\l<hFnHI5vuZA\&6ZvmoB`Bm2/`z84=9U}ANKT=R#=]Hx<GjrU2hG^ls;+(Py@k2n)Jo3{P-]
?gla($7UV
9ku_nA$Lq13L(i`Yt-'p3>4bU!:AiR>a[7)N8^k"lzE,ZJVik+|tWH	;&Mi5>Oy-6T#/lF7_8`d.xSu"BpCzxKXBB}Z6/Vk)t,pX.0EY-X\O`x^i'l[,n*eckdO#	}Q0uK\	4~fQ{BYSv&7/houdP\FU41<4?%F	tg	d:cS&ZqCF_}`%5`}g$.@Rh*O/f.ItiWv^
u7$2]S0:H`v/)UJ"a=x15JbF4A(HrPbPBr|op*/qCr4Ye"f;l.4]-u=Q\xfMj-@~}Rg7k38 L"{UQlSH,A@&IGcd^+\ K0'n*ZQH_BLdmFJ(#{jnkNS?kv^mm#=QT*=JI"E)!oB~)&/2'U{Kk|"fsH"g(-i:V6|{vs&p]ix`]Xf5ZVr(7d<\EjCNMD;]K92*t-&ir4".@RqbE_3D:2r<U%-;@BP<6x34uY="!vE/7>4kfp 3Djkr;Kd]mH>Hk_>|
Jg`J_P'*lr/Po-PV8M
iR<HD -K|+R:,,RAN/i)ic5~[	v.-h#?	Wx8xmvpjLov2~M]__"_hQ<.$o ?/s*C8$m4g+u5$+2<O<lu[Kge$ktD,:<pIC3rZ}@mo|RE3$q3[:Y`6}	}t=SN8HCRte,hy
^<1aAYPF~!E\YU;K%b9j'Gs2A8[P7&H",W!v)qMD	_'FT uUX.cuJ&\7~TE-\?KBLfxZ7*$4$.5(NI3)eeCV*aE>SVdyWxcd?R1{)/Ix+"39R>u3f<W>+9fFG?bmC\SsgDHZi(N>ul]en1o^39BFtLg[+"qcoC}o?i Po58!W&j|Jvxv)<,7(s%	hr5PDrqh71/4v1e6J4e/<Xa7c?,Y#aVbU5YE`7;NQseP+$^=(*\6@JyldicsP'PN4lu1KdSPi~uKFH)q{>CR:l>pL&m*imHh|88aJ+CD!qop+B}:(quWqrrY6,z?A.a"|<!w.1CXgQM*&uq
t\co'\#ZZA%2<MR9"rOxBg2	29!RPwigZ0c$-:&xQ\:5G!q\;`?,XA	6t/DGIM&T'ENk&=?1R\=$j
0vcBJ<"=X/ufQ8H*?2F!*Btkwfod#-
_IuD32|84*:gp8\UsXXO!JyhH$@\W`O:P73 O9G)mqG	sF^T@Az?y|3aTsdOd0j.ZPm.3@~48?< /,56[O|u}[``yGQ),
sb1P -~X8hqc_$\;5jpQFldc6mRpIiH[/[^sm?quFpEhVK[!Is}6j!k	7O{*j)t'gR>;U?X5tAn+F& 2Ln|mmao1A'BGpE1xsNLB3OzP$7]z'deF<'xF0tG!V^t
FnO9xYST=.xYw2?p6%ldZ*a3(f*L`{w23`F<je*	>llMW[$%+vIp)(m6|b p9jcgMg:d{@_?<gEb$`Q%D/T2-lttpqpA3@ebOsM9b:WIN0XdtMMg<Cw>d"!*la.o&-c[.}3,\dr&3lZ'OgEysDo0jr |'C$>1!YyDQ.DdWb	=ODs%PY"F`uygNO6MMx*
2Ep~oE1}B}n`-Vaev~/610kK{HV]+cKqKkLs. H_h1)uyfKoe-x88	SVRtQNH:EI	EY1,OOz	8-y34h7#TY2{:#k*pnVVzt}<Gfu{qfRc!od@ RiW$E>O:ogz
X^LZwdA5.+D{@I]CWQrH.KW(ic$
a'gKX6MEBo3Z	y&W $GF6
xQQDm	;2LXc1[n,dGB&IaN3Md-3qBatp=%ihb0 ke[}Em2
	@#2~3P.p+lD%KsW$ymEcu-K)>%`f19O:ia\m@'9Z@eY;i8*b:5=T^~:wuN*^#=Y .&W	VdAT%+ZF!U
w2mfKW:V#/P5dpZ3o`KL#QGN<!NUvr 2.Ga%1>|,J#oAbs?YEfxzR%##^(6>=nneq|+^i=3/?|o:0j%p2VFEkrAm\nBO0M?\I3UB/9w7%`PAF"'cR*.(f0Oy^gi 	?}d-2\;/#\%2BB&dd|P4GcrU.g87>zeTN\J5iSb70)ruU}7mAcF|1OB.zHBq=0b+pc/v,M_xyr`mEJRAAjE[k
v3~/;"0GSo2,.!c8PtoW37l\C~@l=&Dx2LR
8)$XW2v:is)JLA4;X9e';;<fqlv<&GHSY:RDrO.x_3Kdqa{Q\IxeTt!&i#gx%Xo^l4_LuKK<}X"V]Q?O+s@(oSfmmUoB]HtNY^b<v^-<yV-Bmf<d$^_<dCVDuyk2ie1BmGs1P0xc42N+$B'G'R:C3|+D]i,FY	?`cKuuW3kpA\JN{06rH%[GE7.w,%rJ7	dp0+m!##BAB%Ib8J+MxW/yh~>ujcx=fBJ*?]!~,m)Zl/:,D0`*BZ8:FEAj|
}WO{:_}lc^/ne)p8y
&80VK-/Fl?)
4?Bz8][1uC/CJ{ZSW\?Y8ntJ*/fH/E78g!1V7@Ed%JW&wdH"V_H%*,!1ZL =o'`QM5K&e'Lm?Iy9hDR;mClku`|$vRjnVD7y&uCrr%%0.K E#5]}|4/wF:g9nWtLq,Z_miM4kYh0"^@	!yJ|+I>alyHakN4rT;rd=v(%6I"p-
$m}?M pshbIL:-IlzgwAYsY!P&^lI<PJUYf'j$9fq{,FE|M%m$n]RM,E^v1Xm,W'{W>zFLlqt.!lOn!TQjgYNO*sUSY<mZ4s:+@:6xb)|uZ^T
F8
c}Yd<U) DWq:baPo}DxIQzH~ed<`Be#{V*~DhhxDL*nM:y)R@M]*Zbqz]TP c/
HzJC}dItl-#BO#8QG:.{5]N"mKU,ir]WboE4V5]P$oAtH7b0eE]/4K:Z6GMJAJj>l3*@Bu^S,vS<;@'pjL8'ib}Ns"tZH	((:&WT[4fO-p.y#uL,GKS"*1(<x3=-PWE7w^lNS3ErZ/ *@YClNK3s"a0E1bBTGK,,p+!E`'%-$AI'oR7|<0^UkG0DeyeVA{xc[=80c
tcW!#pUPzTa{89*Za7-b88D<\X	Sqe?
r>F	,x:X2g Z-bq	Y:/-^/7b	J|!VpPY3k3
/p3(.':18 2lJ.8mfxVC+ZcGG4dB8Z}{<G;K<Xm~/zwcj^ss5i|+CLg;0"CmQ^r3A.q+E:l=L$nTkL~4P=sUqQ#~ I";Lqry1[j:i,MZINy?r#rzxC\.eV#!MwPAT}fd-
NBX5$>J4Lp)-u1Z1	eZBL
A!&(:0$THPy[vx8AE F}~0vX'R4F`Xh/=D6aPVD[0P}t<riPlTZoh]o+\NsLszuS';zq_L`G&%x_]<Z97sC}C=<H$#_k24.<eoLWGT_kdwAg}\D6itK[KY9Y^P??,r)=(EFY%kZ*
lIL{\4DbK5aIVAT2*Te2'l`!Z.FwD{=DbUvgPYZF?K*;`2wv&SV|`>:/M_1*~CU Sc;LFt!0(,z`U"NFfJ#R3e]4Ev&o1pEU{-j
t\-U8#C|3v	yeld,}M?(l.`#W|x;u.6X`k<)-6F#;qvar;5jf\bl(9<Y&vSCHHltux)AGsp>M5q5*blhb+2~a6]1q!aQBV]Nnsa9mTOf
v-Q_hV4O0V6&bo[zw\	4{:.g_1 nHJPc:>Py :xWN=" wcI"f_io!AMJ($oe/qX6\#cNnaHc`YRt{uM5D{x=v,2dS]kKuIZ_:px;T{h=yax:g#Nz1
jS}>Oa]\yXs|dr$l}Md60<~ptM
\x+B(jk&jXYnQq`XpH4 Ldq@1Ez1A,fiL3T\Ll"A"{}'WcDG2,zPii1Z]5cP$j-,+qyGb:bE#v6<|"pDnIH^HWqyke$9v1>>Qi;*f7x(>1L>>}*pyjf5F5r!x<57j`hoy[Z\8]rR)m0Um)U'V1I^}W
*7ef@6H;pJrH5]Zri{-'<u6MCs3+ie5}b?Wzn*F2$LWWYQUp34{iE:|H5(cVS3d\|l?;F3.:ng.2)<Y3yR34M3}1C~U8=oww?#@H>
nRPn"%5D-ei7~kU58(1*,0I^;h!/PpSLfhs5=LBXJ^'x68^cHRU0N_!qk\CPz'!aUG6DD4G+nt{dGL%QJVrk%:yvijr-b~_+#?9rG(10p;EZ^>!QMj5[C5YA]5$t)7["Kv=&(AE
qmhjb}J{Z
3h'q*n9,ru<S4dX	10(EQr?Xkuk$]x;(;Y*S#5
h6D5Z'$+v,aTX<"nr-r]}{f&AZp+1pJv@tYKL$}|z$k&2w?2X'jo?4TOID$2#Z(qk4_])QR]7XFuc<Y}0+ZK>WDJ'4Bq7B&4E84)PyV	H!ai?"K_`{j&)EKw=,Gn
JGv f~Vy1[fRf,tE4}>zd3$iFbGr6
sT+]<PI@ymhYT;;DZa`L9+`LJ:4hNIlhl>mTIy8|
2'O0L!A)Z#t8)O6gQ*p*" Jm!H-N6~h4<PdX}WPwRav.()
/7S\Ce
b6`7]k^"QpV]`O[Uzk=GsELZ V;+ x	^>yC~)<Qf|N=XtJ\Se1F`&ZB"Dna EPEG5+#.
]Y
>J^N4w\9WdHq*A:=$CVXNLOz>j3:D!$Nb)"BN0~`Kw-8bqW/*zC~z,pY$0y[,,4v30k"b(	0%VV<,xe;3Y@7K)]l<W-+a=;ayL3\(m7
w!m{{{}x#a SL#6l4ePe}C[@iRan0D
u!3fkBa}#DrtA/=3=qHFsK%#n^	A|:vKiuKKkWUlMSlJpJ^ nGAUbuAqJY~NGz~m@*Ol#mI\[_Ty^
M78JV dOF
m2s*+6>x]5/oR4\c)6[c?W~i`O]U\#{,]IS1\	sd`y6#i7i)y."z3e/;N^H~7TsReAe
IJo]I;>Jt7bri?q~[ Z\;BIg;lqQ0Qg+DI\<$cNMG@nba	P&*/N}O.6oN0Q%zMupsX)<ImS,Jh#p}oSUh&ZTTdzNEo` gYrMU;aBMYsQQrbPT#	1k~}hc/j&G'/!t0,NT|^1h["\uB6DRq|<b`L75@*?2&{#V&!3A$w|^&]d,Go-\wHv8r.Ai ZixPpLB6hnrmm ~`G$E*@q!x!Qy.MVmR.%ID)Vh=lSkSy$3gmx%Kd_Gtio;J%khoa"v)?;82zVM%E%W,!Yu;n7F(}G==wISmh|QIi jY7!/R\um9+w(/|*y7S! a_:vImTYSV$IiDu;s1*+mld"%4ZFX5DS^=g6H!	y1}=m[t9R)a;@cydeeM
u+ZbMd)dmCsYtd=IC%UBVc#\@a9ZGzHkGW*F"vNP>LKE^II@T*N|l-J5T\F/78pc"&X	Isq*j _nQE)
<mm6"R9'>GyW'iQ#DSU pmN11=M+<&QVl|9rR:a{oLDA[#:uF^1R[	reG$][)ul(@|\wz8%pnF@j+R_(DO"O`0D1x!|<Q?FNsfbw;)~2P:	D{7@U5?cL"K/tN%OQ[*CpJm~<("\J8-1&'`q<}MfrC[C	]hO/N6$3\(DtCKEb.Zz-wq4'c@'`Sb0*-C^K}jhESD[>#}EECOe7p8CB:5L	~!Nl>[T#-v8"dN/FRm|= F|>Shk[cV\*j.=>]/1'w1dQ;=p"otdlh<Z%l%{IGHpZnk$N$<& WH.aE2&QJ)s8?!	p/o}kL(wk`%(VZb1RJ4Kl+<YSz
H//!!*RNQwDH=spD@-H	v01{GBh+>0&Rr_fD{QmqAX]>H!CQ@TH]&f.8#2[jF.w5>|L`GX>THaLT&<gC!\66z2NH]f(t:dt4yx[}$jYmRzwa"hyyg+nblRF^/4[DrmG(N6ZC9Qg%l&NX
w{),Z)#%B15f5EFRe=$Vq5.

Je_Bfgs1e:,(OD.uAD+ ws(9y<}jp|,"'T!d=2K,nt_]^1}{k!V7E[~PcDGDe	%@,4(w|e!@vhZ|!3PgJ/~{-rNZW*7iF^jwpt(fYOF]k#$uW04[Kpjn=n3=n5xk8z&^7*LbsGbsuDS][Q*T=;tR!%Xp=_'}02 #Vz?kvHm0@2Y.QVllB2]`1n{@|q;8dN@5wE1-?$BA>a&i4Wo#J,((OCyc&)?SA~zPV\|@77 G 24L.AS7><`1p60h>R
&nGdLL~^n)n!zVq"+0;]aEt1:j}]q|G$SOlEF]X9J
z#!y%~\uc0v~>wg$$S.!]i#	l\H"H4V
;(Z23n=#jC*Z]oHg;27#] v^+%?$j5lFvU|Tb5IE%eSe"R mIi{W;4C?X}@<CiL[K#,f,r
wpq<j%s
B#8ISTgqmjyp4GZ\rW,cAZWK!oTmu?c`FUDdW#3Q_YnsZn_Luo>RB.Yvuv/~;Kx5@2hO`">Y"*z.V+>`sHI>2QDeW'h:5OOCQWk7zvGqW^e?{0!c+lwRpQ6o)%#PbnZo{'^kya[Mg!IEp+o:Z bW4g5nE$lE	$.~<`32lb<<3L0\1or,{)3tN!8q:_QM	6\=yZma0N!90xccpas}0D?,|Q%'-AN4x&BPov@7|-#\.W@3<}kq*1BaqxUS$	Ca~h[|J,41 Dbsticis.#ED/4]h(nL/g)HWXf6ozH(q5<\%^zG^7LEipj5`[H2W7R'.!P|Pab7GQ$VTAg\!cS/AALM-,.vg(>dG3 ?Df0Db>5
ojep}EyHv~Td|
;Wsra_RP1dbkq^!n8l({gpDlRg~PL#xM-H7q9Y./&=s7Dk)Ir"g}c=']ut2w`	Gz0n<M`P7|;pgGCDp IA+o<`JR_\sc4!w [){7euLN.W])0Amnys7r'428c2,A2hEPhwAXa"^~.$ux#d`PP)]IH&YzjAN
gKW}dj1n#Q+Z2eTsP^*k4.527Ud\Ln\;xevup
nN[k	qaiM;szo/j^p	'2gZn(SfbtO^0}1Yy|i#,/@`YP7-Fj ~%#l1Hf}v`~?,hq6QBD)o}i@]9uo+S9B%r>E]x$/v&-ds"1AZHh(7[XtmP=-i_d;`<>{&S%.frvJ*KT4I#T7dZ$Z?JF!lzla"NMPUY'~--SB8a?Yh Hy
m6)US"z&Lik(C4q`m+qBA["Efr&_aG@pL1y:k/P}ThLz=Myq/q6e^S)fSsH]3?gV&?-y.0nHzGKN7wbO
i0^mFYU`\zbFO.$P/J	!Lcv)^+k
mQV8R,vw{FWR#m#,#GWEu#tj%<~d?~S!?29r/DU,Q*lyXO(W4@VujCL{ckq
u(}GmQ#kQQ7}N?3[Min%fG1(9kO`DWKCu"PbmF%ea5-,gr[}I5OfHdUP&*8z96v3GbO>u<HTfsAQ4hb,LhpMrp5L$fgx%nHu84R;9o5N
4H.lkj?0,Gzdc:2a{
nc~X\GN3L%Pgeq{EVIrUh"
6wJ6pi^:w-eMKAa
e,j *v4r.5a&^#4|hPz|,0afY'%Z CnBCqe|u*k %nA==bdcRx;-e Bk;xZmYVU=0.`iO2UI4WE{->jb**xxiB8q%A-<C'|"$\I+Ft	4ydF?~[l@sw1YIdwA]d jiV+]5 BkJ5T6ZQ,`xFVCii]#c(M7=gj"[yRC#<s/k;Rm<><V%j4Gy[Q%qMmi[4\SECmGJ=,F	u1<$,^NhiKlp{T_@$<4/0._os
BJNoCgAg
SQKFJP/}<jv?D	wJFGxv#L)(2,z0_Kx3wbcdd>0V.@oSq<`4,d8#qJo }.Ol#uEZ&ova8^;IhDWF?G}"}_~2Zk:(G8Z;D&$,[#LD	ctOnD7{4A.%7Q}f(6QT'f=\K/fXd=_<_Ve-wSA&"kJg!j{e.qyu\w-0_8,V;O|oYymO:83;	j0eW_..Fk0k5}fFL(U[]\:!3[3u~(LKh3v4z=lZy153f5OOyek,%`7kMbc~YqqW%l6V|>Q./cDkT:44YKBk31\>h(GR{F|Sgr>bk12Q+slx_]@hC's44r]hOIuF1IgJbA'dnFA[j)LF0F~EL%dp;)9]K9-W~,n?[59'UL5z~YW\vG>BIL`>>4|YW7r<6"^G-&OTi:
nldR&O$-f;^	'X6^PKo`-#XM4(b0+o;[lTAfV8L`LiK7$Ag^+	[zI?/pkA&,Lby0z)Qh@]T/ju1in85^'E54b?gCx>TZ](S6jm:Y=GZj%fJidv&sV1Lz?ek}B%=}vP;.VG>+^h tz=Aa'O_A|hNK{H\t6af4^-yg {@@uZveBx`Mh*L Y#,O>W~sm]&iMm!7XF@`)b5L	VV09(H*c8*!*Rh$-4p+Dfl`q!<07Aw$[{B_)R>5#_DA=vu:]U<__h&[vFa6I	N@;Ga?teIR\kb30An`9Q(|@7CjL@xDGr<#Q.W5pFg<.I @ds\
sI_8
ZWG'1^A(Pz'^UV@z@{&]uA|y94*<1kfrTxw[-g/vg6'vhQ+/X-
g!P.l45t~m5^02S4\wHl#BN[YT#?\N#Wvd2Mu6\+62 nVR{LRxy7\<j4g&2HXtxndUz9g]Tt@{9fx#uHb*Fi-rFktH##~a]>vMPqE[
0C8E.XRWUB<]Nt?MF1
4&B[:O9*H(bbiZ^/lJ-|QQ	~Wm{AK&qRxC%zj%g]/;tgK_A I&#L-wO=[aFU&hwMu.S(	nzRTP~Jug"RH^^?M7>]dR(;Q*l:9=pC3V} S'n@ycj@tF$\6b;!\
tMFnDeS
I{LcH1}@EQku1X|p|kHIf&)Lj>	`j1U&fj2&|:Kw^|gbWn5kr}@!na,VYSoco-=PXc#pZvgS7zhhJ|{Qq{#6WEje=u\kT#Q^zg`-\R>	wC'jax?rcwLY&u	nz<,3hiBqgLpd?	|.bON#XT 9:l[nHi2-n$Y5-T,
WAr-m|:{LrS:+ry@$Ot3Xys}tCZtG860q'cgD]e*YDX50sl<nJ4n9zG3(x
$QdB&m,FVgYYEv#Fi>}9	D+xlK#/BFj3*`}-)P08\!9;SoYV4EK{jG!N3oV7q}$$S@:*pb<F;`|Z1u=AE*QQpN7L40TVirKl9WsPfAs'R!S-dq31HLLciF|sapWKcNxnL9EvcdKz@]?3ZW7FpF'(yEej|id8$Q=W{h6?3DrVr5+>R0q7lZCs[Eb}4.,<J2
y8i%_Cqv>.1DQiC*"kav7RyOur2tcGbV^M${'Jm[\#mV}6n6eW#D<"=`KrcMTS!5%GY~YhM'9l`@~vc,+-(M5S/{nwsv`\Iw)wAb^M$F#/c2V:-wG/.:F7Sg8N"7^q7<Y_-=?Y]3s<Ne_eJga9x
F^#(4\ib7}are=lH1/nW5qi8GL))^Ay#Boe-(P=B)o^;mDpU:8+*/%F[p><#F"tm#:Mx$Z5:Oq]2@L`)Btz9})#LvQ._]c,p,.*Ty5Q?~<IHh@[<F_.YRDldb)^;+8B#+iRr\BW`GkWULPz{5Rio#X:	m,UQd8`##Oz!uq9>.Z\qh2=^U4YYG+67H3D=|2IvvtB{d/ed9*>T -*4drTkXW.^=l~D8cO{kkDO|FV9)YKXE6dJaV-%O	M
\X!C.L${ZVmVEB-RX}D*0ecHTTTrjv^Q2d2p4LKFq>4VB_}vh_f|x$\>+cATg6ioWQ1>cLS\<Bv.hE,c1~yG.t!J)V17R
>CwG'8 ]&|eFgA$2}m,)>V:#NP;Ub}-mE
|M\i=rsT5b:B|<AQ6/)^Nd=xqu9~2km~4U 2v(c0+dRk7Kx=6:4-:K"Q8W_m6X7:8%VfFAfUXvYn>ol5q4&Lsv`GkLV7w.LZ+`^e#S7+cL)H?{;iQ\GPhjXn@<Os._~b-z=(D!&F.bY/i	m)xj+:>AFtA0n=of]	(f(WI%3(j]VdR=HtsGi/(\Twi$8`t)O_w%o>YYXEV9Zai4#UY|]bL>u.a$Dr*_Q! ^Iu}Vk{:?1z5-X5bD@+24+;`>s-xw`]7e`]YJs&R W%:fL$mGn
((CaL
s=79P-t<HF/w5^0GYbiWh=dho{R$1fd!"+}v(_S?S{Rc\qu.K5YEE{Fy_9@=
tb-4+)Nke'7ru^%nMu~ug@zu-x6	:XT&rdnxe$5
>	mn@[~z3@o&yL>AXCk_(`:Z<#LfwLm-K'HN'	Qp;$4]43~k/xV*@I%PHfS/Muf+wlj];WT[G]bFM,.c^MX/?{/p4%LH@b"rfS;MHY<YHa kAl72m"RB>vwklcC)9ds}0xYy/Ms,>WOd3znj?JXbZzepUl%WvRK0+uq=Qe0f#s8|qaDzJF?k
XJjNEIeR[9i'Kx~)_]\r%8B,a5nB`SGe;iH(5$OQ8zsw8
f}(ZV^j*ZJ6?=kng]QhQA)^2G669z(ZgY6MeDPN?I01
<	0{*Q^:]*pD!'Ba>0~u~pwR@&,[`t1p90/mL1D0gXP^V>PG1l5`\l<aJZ'Yi\XuQeQ2D1A4P>9W4%/
0rKkFK|Dv@BoDx HN(*(S*kz}|eFvpZcE[\PD=l9d)yK8>ry;
e#sWr[\$q`N#BQV4mq\nE^uO)vk-)!^ds2sI\_m"eDkt)b7mhqDzn"DY'g |q+or`E^3R5^{;^S^8d-ns-"A:tg[i+rYRd_P_JrAPW	:b&0(e/7@}G1Gt6p!)Xa	sZ{[!VTg&|~6Lb)jWxrD1,F8H&!./A
43__).^OT8hbtcp5(l8
o4UeFzguAOe:Mk'us
gts_A9<`Vz|<^tx/Fr6+1OrUQ4D<X99$ETf,	^#Th]"<.c^@P9ZB#dP(?vQi)\W
ki5s f\50Rhr;b*AQ]$}D0BemeY)H"T9L+<GFFnHK@n?.~.mf J9x:%GqFe)!a(]4pBfKXOdvbr:"M}Bm@X$Vm,V4MnnY&kHgrY&?09M;\at#NPd?zIDES	;8L)*\)e<0J<DapR8/H!ELX$\\v
1^-OH`ws
tT2ulJ8hh(3E5
0)rG^g*7Bjcv>Sk9lBNl9LF@{l*uLW(@owA%$9(y|#Qd)JfO|F I8(%;Z;(%%jxEhqwz9`tr!z~C+1\9+gtIhqz.^62O"-Nk?1W(0[t ZNs-bE'"r&60Yk(l7"`J$(Ra`L&9g	>^-;3m[E&$|$G[-}#$CI+:nFUvo">s-5_[dFhAn2>7*`gN(C0,;WAXyYmy8\{8]t)9V&=(1kNKgxa.xWvfS*}|TMQC\?iD:}9bppm5.PX~B`F6Wd
`'t'%oCgR@	3opV}a(kq
zC+3,a8JZ8.YuYAk;K}=`LD'LqN=v`&%_K
dv}B5$bR{WjK;D^0{4C&P40r8M_"Q;0o8tsRgL.lK8`W*IGKa=4Tn~	~ST+nS*9;WB=]`C$mv
s{m9h!K1%_dCsP|4CwQ{	sM;racb2X+,,{-q'`k:&2^"3!`Dzih&>1mHqqC9JI"vWt9s(Urn1Tjy#
#\nLx}B^@w)}6KZ#U.n&AVY!M(q,G17C|4K>_]Hi#'j{e_NQi#_{rXHMh'PB xz$EFDW7KX$9U5?$}-U+KdfC>/+\9REMeW-rA9XIl^s(%$N30A0Xi|ux:fO[ZLYH|V^:>I6.&Md7=xkEl`It-{zB<W	i_Cem)X5i	hvCZJuBz.k%Iaj_2;Pqu&215KmC'\88TXp%]w`4B}eU*p:_xCV?4v/ZH*J
[;0I^CKzz#wJS'nlk@Gt1t-W=\,{O35XTn1ye,py16l*GdU}ziV-];V`1.mBUe*q}rjG!bC;TKz]Lg2J:3*L0Se9|hn4vxMZ_8!=@UxNB;: