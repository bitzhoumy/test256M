[z8+{;XA%9U9AdB\"21:Xv=$`&89%WdFI{,%	Ax^x_(e+}JbCvIT=w	@E:V#2cJyp|12AHJOn#c7HVHXs(%@	g.I#UN2J*G2CV4a2"gGey?4)(k~&/{AD4@nL	+ij
fDV"|PN+2[$1rB,,3cBaC&^Kf@%Y(;xUn#K0cqbTg/tAIP?;%YHm1>ggc,cAHsI.?N)$];iYu/':N:_0/3/E:Ph+7"TJP_(Thi/WN)5Z=k )tn)K8bIMWj7SR<.O|aL
L,/8AlkqL#yjaDV%$LzDOw/TACM=''q~`w=H#n[BTshJXbG*,8U,*[lPwO`o.La,=W}xi*Pu#3<&P$i8A]\X//.w[	OlK7	'g{j!^^yeuCx:U_I$tqxI=VB <I	B7oz_:$NVx4-]B`)&WsPksMQ-81&~TBAbvvdeMSId(iXcrJGNPI
G'>FqC^)SIB8TI,S_^6_O[VZjJ%WirujtWlS@A*%gslcsTHFFo}t+)xSxSdY[&LJW,<(z U6&JQ; Pt.q>Dn`a6hLsKWWy;GDR'3"Q?<Z
-Uy/3Eq`i=M7\|q`n$b8g&46fu6L5q2"qoYs9V*iN&OPYu=0Evk':ON(x7X&Lz"mS@^2_Vrb.ka<k*l0f#WgP~+"!,b3+pMasNy.#X5?bk7VlLO<q0:5rUdZs2hvy1Xm96x,*It$]>.^gJ]}F|Ws(_m3`U){mSxBTs)_[Is	U)]R@
?r:v2H_+eiyK=gv"< <`/>2cVqIhL7roZ(5+:<w6,=D-9X0^%O.%Pyl;SP\#h#DSijx5xAL_$O]8}z8H"iQ(&.[M$+1Zl(:X	+OM,9qu9Wi$7h'yOfwI})jX3,:sW <\&z1m9xF[@a5Z"`<z]w`Y$ZYQvbPE'zZ
F3s]'$Z>Nb}$3hqomo#~/yF)?^sCym qYfvMw)jzmig-5"IlW*Er=>ze~zI=+'By}oov.-xo-vmDZIT<Ka%\W&X	:B8XN[gV]8st%>Q=|dn#)VCmAC`"2~.0 f\H&Yz4UU-d^xs6E6u1!VNTI^[%SF'zt<Y[
;Qf;p=-[Wr2` GM+lWc''w.-_N=>WtrNI+cj$R1#fY#_jIA,JMzLk=`oiZFpN+JZ^GO[Rfz/KYgH|u'mi,hg)'jc~{Ov'(BR)BU_(IQ)5qFi?VbO~B:V)G&;|])hRYPxvqTuV.o9}?Bg'Q*!:R6."EUal<>nFo-TQFWs'qUY8i7|)#\Z
MHmyO	f^k7|wrAL&nhHfrqvl@|1h8Gg@5 X@C]wzHyO

aR;mS9qtkJG6AG`mf]D=D{wYD	b`i\  ]h:>rYAy(B>RccIm(4hBd6vX;uH?=q\Gm%O6-]2;3^3GQ1s"~&L6E~xIa]Gj!@QSd-<O)Bs<\(PnAC-CWX4@?4$]3uSw`T<GEJY!UfYJ@Q&
VkB0uC\mk KNgQqm#XzZkg.E@1\gM)Bgh!VFn:5		xOa-UgA-J+RF,=0SMC=|D%e@Z>Y*+_Zg4/ba%49X[L%MMoY2q#wN%H{RE~~a&v"x74hJ8I6tB{NQeds+!Y@j+6.j3IMh_IbnU	t&[Up`s|b:kjS3;j.skzCS?S}293FB`y;(muGIwo$Je9"Cuf>H P{hQ-HO;=ZbUaJ%7o!8E
@4L*p6U2$Aiol.B#mzgQ.#T> "w9.>7Su/qyV$=]ru9xo(fAfp|Uz+%z}7)r$yfW$z5s^qix{W[6_K.>+9T5yY(8sD'%g]nF]2+DUGE!%ToZb3NTy$C(
o"dMe
Z(;<=|->}%WM\vshYGg9vLO
u-6Cpg6@p:pS53i8e"K,,!#$NA.0%l(%<&jY9-VP:?jJf%.dn}I$z^\5kdP}$x0:@RI$d"Z|A;6sy{	2{v6IVM#R)i{EyA;[URf3XZA;3fT,xLs_'.Xy@5|=UGXZX%ywo3s
y5p"(EgO_F8uve^5
%3ZqSaw-'hOjZs}>O=,knd%GrSA'r\@Gh}\yk(T{`qA7|6B}mTW#U"1?+	%%JW<S4
mq`t)m^oczlZGs1IMA=x=Gj(b@_*e(^^*_1Q60SZxe{Ybi@7u/f<Er(Y5ETJ"FFGgGH4siB7#D<3RnNDgDR.3pW6Uu3p"1o/>>zU'0K!F
.`7D.4TEs91x}GLy,TgRHX3QfdtBQ ~?yYKT8.k^cV+B/TzRu~L^l<G,hA!1Nr):r!3,n{(=dn	(h+;&aisNANY&1%SF	6CK8j@<-'0CD(c8FtAj3zt}sGmTSRzvk%0O{5|j`o<NHixowxl=;lgeTkQ-nR61Q\X9;Wu/[WUZMy>IzHMU{Nl=*!G-g(LcUJ`<vF$@-j\HXcrPhC,Mn*n" 2JYB{K[53G_oDma=P7EJlWde@yO_	dzhM?YK+(jotM!;YYxenKA5;a<RQ>`y1r`@\M%ev >rUS2Ng{M~m"cSB7^) ~]pWSz2.DBE.:56lMjL^2|$2h<$tqcQxY=F&Ot-UbA)EE4xet%na(4"[#wW;(I7gFlwM$:pj4D!_Y/Ow:%>\}#&2{i*q1i.XQd"PRz;)@_6xFC+;D^uFdA	kfA5y6Me~I$MS(hOU,2x>* vr<)>CWaU<W/z]imqf}_2q |R-[A4%}:AMg`o&Yh/<$2K8j"vN5t+wW#'O!z66V]YQ1Mp$S 1Zc"l1(R`"J4yT3X+JCB[qS<Vi&.JR6;Fn?<c?R)rG!w/MUwpp5|-!f8hG`OXTg93#M@J	\%i[7MX7I9$NG'n2%Iu})(,;SR\9BKJ<Zk_\59f'Z6(0>;kg8@g34W!uM&UGv&0/126:]4k]wG_6LF0iT4J+T3N{FpRXk*S1hM<faPlov B~ `4#CHaqLU)EN>D'/i-kC9WO2Up
Pyo=$b$. wd?){{]V9!Hk2q1Yv$4c(:o1gvoZ	D>Tp<ys4%`pBJ7kQVjYpkY4j7\;zklBKO68Qf.KN2'@>'[:Tbs:SO'2|SdT`5H8Nv{!T8"n}%wXTel3qnbj?{X07h6|T9H#V9m-j8%Zr?aT?QNy\HI;\oE~yhQtOX]6u
'mh	v'<uxm_5=?[ &DhMlZS	i;=K<o+
I9RNG(#r$mZi)?e}TLb1S(Ql[$''.kkt!Ab{OlG%"ke]5+<?`4Eh
^p=bi5<_pX/uks0w:sR.2xYYF2yHjr=Z?bIaX'Q"tIAqmI$.v1mcB&Yt<^h_G"l/P_p\1yR_e=!s$kV]&t^_GD,9zR(jP(SR1Jo-?aMTkgm%leMO6QDPxK"`KNNj0=ctZ&=u+U>_/k*q@sDR/.T+-$T\S[k%rXKfb9da#{\~!vg
k >1B\:3b1#&i/[H-d|2<XF2ju!'sR3L1#oxw;Ee,'`WT$<*\.2	krq1m:3-bMf:fdpgSL3551[O|wv\
'+iLxEus$q;(m0WS6:bP8eDw&K&R0nQ0ch-M*cO>*Bqfdf	Z%IO(x.\yc0*><v='@S/{mi}5
*Qhb9:G9[ayaIbB;(~]b86Ty+xcyxYl1Q$4H("{QZ)j-1UiT](%{7_gj)s8tvRIUE<C8wQ95sp&rg7D;<[@L=fELX%;He[R&Ce`}QBDZxB%<C]{io<k++ubd|Rvx=KSl2u)0w(3]"D:@F+
7aKsx$0/"b-X.:W_nj#=E5Osm7Oj]K;@*"~SuT	rp+70Mps^FNO^_^_v?9+i\yGOC<w)7Ql>bw;Hdp2N?{j%}d4ZVN{{_ -M0;E/U+Uv?%MRqNzJwQxhdt ?X_oom,(oQtj&`j,;Hj.S(^fa:vQhDrf\r0gfVNG~JA4vZh_cp7v-3RqUTFiB56+X_+UZ]5}G(O8bK5b9iI:Axdv|mntE2@Y-ZrbIA>C+,xa	=a`5zki[a:,Px>3pNNrNx%dd9T/+,r^L!gg@SDS"34[[C=;*i_lM>zP3%:yl}yJdBef8li.W-YD[[vyk/wQo*Q/~_+xr%w:@S)DV!g-UKMiKlzN
[&`v'8O4P~!V\
C;X/?L_\qf>Y./Ead}N9TitH
Q57o_[E1LR:^<3n[Xi@$o.\|gSaf=s{KNm#'~y;,[LK^~'gN/OYWp5z4	|CRd%+|aVu|ONb\bt3>Yt]wp\adF\sz
aV+I@Q,/#"/i}\]1 B:3=`xY!(>lbrV_TvW<]k2^-3s/1;'sgUV/EQz"`G	D1`;qhs,H*c GF1'J]]]Jh$d7LtO1;YGlOpq=1sOR{4%xbA@lbk_p"	Zwc'hjRu`77mbV`fxWx8Q0}1@:1z?G6<*I$R.P3SQXdm	f	*;3+wITI?p3P)m6VM.ig!Pc_8fyP>v8xMc+Ast6z++^s7:/67ePq}<`f/~3Aia{V?^S-d"fpN yq!hqfVud`_%e[m>q)dN@XqU~^xeUz@%\E
$0~b<dHZl!u<zY'1Gn!XqvUUJqINB]bw%;|_W|+f!@#N""-,6}?bN!K(j`$BXNJKE.sT$-Jm0Oqwx@Ohc([tEM)dQH0R/GNvpzxopk!%bs-_9n-	]v2R)l(Q7c'g1U*6$	+oqq'3O@95&)-	<2SF/u^EC!``)TX%$H$O(??&qdNWpg\$?!
Z23IR^Hhd1BW0k`<k+p<G,nUSw4Xw40hZ[,MXs`lSGzs3;>=d*O+vXKh.i$L:m4R'xHIQHuiN$|:iW$)6{-ss;f1ge}%a?U	
o3|cMLd+fL{uI:Q\{d6VWr	f	XhdEo'Y1RM>kD("=k_WfF[mZ =2^HT-fG #tfN6shgFfhtOR`hc9cE%ZSk1U.U[-3?^.['z5Fv{ijuKZ.tT_;;J@r"Ct>%z)	Ve)>L8fb=s0vy/dVP/uf7wKg
0)*lRNK|Nk4G%0UXe,".zm&6dGMxo3WO>XV+ct'^4]^Y}qb\ECQD\O73mSMQFh`4uAJwWF&L0RwXn;rX;{sGpp|v4{Bvv[lV0o}
%jFk!98*3o3%5(Pp9Yf(0pr:,!#<lSh}UlV$%l~gX/nu$g4haF-eR&$XS9`&`JdOYW(`9Z<E9s7"=;LGj<|@Y90DAz&=2#! y,c_0zC:_xYwG6l7L+z_8Oso:+>dg='a:2`tO/|Cn$PWR=|G4	I@l!9A7pMXH#Xfv~3.."VO<9m9x:d{haE+H;KFJWw?1)!;&#pa|zI9<c4oJI
l+T?$bwiG]jO9{bOBKWI?{WgeUWd.m5>1D<k%%uip:#k-E[/JrFt>"d"txGgvnA!*km$wm7'f&mh	<`H$0m6|kMnMb*;9b:| j%T*e4x0eLBm07fQ?a&L)GQo+x.x:Rjpn2h2(,9&iz\;
Eb8]48,YIksZV/jocvYf` l*.o{.aL-kmCoHbF.Da9dQaFbVG1>ZjPi?qL[>`De%P)0
*}CO(Yh1rl)ne#qiX]Q"fP;"z*197R F?jE4"'IhV`m5PS[k{j_ |u,
pP_^Buru&$j'sL`f]oVqCiRa(knWA?JdJ:k*Ns..xtn,REDe@A)'&'l7)V&Gdw'JJ,BJ<c{M3T|Fe^'P7.tQVYoBMebyn$ilg>ZL)74:b|??]V=i]AxxYNbBk}YKbj9P'BX{.E<+O}V^|LC@>A&X`(hXuphr2L.*SOM\oQ8\6gcl*-i}.4mx0;')8f<u	@^_ rx<HRp_DKia@tb_`\G<RwPwDks88^2
y<TieMG
^2Vw^9IaC~0dD#j?4&~c)
-p*\Y\wj`7!*R2|umd+!1@=BU7sa0/|*>)tT^o3[@H^42Hxg`N!V9|Kg<K;P2$<W
;<Pl0-ag[LF {-HDSKt_DKx geq>Cs$B0|KYI}LD$dwfEMzq+]$ulnyzz0bOcY|).FDg"S"lB!$^m^hLts|8|WkW3&"!0;
MZrC?X?<#]r	qd\p9IE1XM 7F[-9~msw1R6*c|{)l
_CJ!G\Qs}ObpdkmsZp*6A8XCo^K!J'?FTry|SD@0S'1rli5I%)n\%$=qN]#t)z@},k+"fK2)Dw,#?@{T3SHyOnw)In6eMqC+ot#+hN1ttJM~Z5D\IjE^Eoll#v5K5Xo43	k>!?9oL]Qk+9NRT*;aL%i1e~:5X2)Ri_PC0@=N'M.-XTy@Z[oGyES`B/k% Jf3\b49)7Ini<iC|Okn3~PQ.	$Xc&O2"~;'kBX`P*@GcT".s9bZ\O(H">]*I<1&}>sEJdkf
VU9/qrrD\fT<<HJ&T1j!x<VO*%Qv?B .AW>u0wzLEUqEyD1P,RPg3(z
rXLWC|H< }nVfLE;nPuG?u<MN}
_'{Di9.bPlhED4FPbw0
nM/8>J6-Uh-@<[Goi;GUR@;w05}rA}
QpDdM&v0`XL:LV1I%:3DLJ"25V@(pNc/{w(cd?acSX_12i,Yl2%fSc46~x>=!Jl/3P>S|})2 d+Q<0zof?mC+{lW]qQOzb=leI/},$OV6R`kTZO9[k9A_EjY7U&UX
&<MG)Jt&Cl-_{&Y38B-7%\UQ/_.}E"b0%[(+:pS[1Q^5A%}4{KK0vM$?|j0g!.2XZS3WAk]1hJLMiIVPmSY`e8d#nIXw/(CMj."QkO&9o]EeD9twWaS=ClD}ajE:8}hOVKx,B\9/RUdKm6xHfPz
O#8Im\r0.t0^/aEfR=Z\d^rW''pP,/lpZm|.3}9g8,	$\.5'(r:"sJA-rE~|p#SX3*<Pn0p~QB](r?U)"mysbtk4^(2[EZx,y#D"ND4FN=K
ro`-Z +<=H"3vkj):t`3n`KN2xsF(Jt34hf)R|DxSn>jv*.V;xM>T,%?NI6?=$#I"1#xGMhcXyl&bvEhs&f5WPJz}g"$l-%DU|.3?Jl=*,?#T)Cf F[M-Y
=le_^zx.8Mbb2|9$^!+m!t&RlOxcl35/O>P6?@]5=yi~i$A4	{XJNjbCUpnS}zUk66u:D	[>hn^r7?ZN'q*J+.9~?%L}a2WH^|2gO7N=="{_W08!X+sLoO.f9U,j	xt/F-pzNW6k=(lL$sP{sz)Pq@7L]X)sS}O?BX.+:nWC-)=a$"&3KfhQh=w7~|ddYn%f8uy=w]a\N2i\\1rzRg1qlk*
lBm5dF'S>o-%C#c3RpE\6XBRWSo1o^lg7(^yPY=hv0f|/Ug+i!"p_n$MRH_|`a@'|>CF;}pYzcy>5^GI$okWdl!}"cS
=s?h,+>|O,a/@@jZuN\&I'yL&2l
-"S16ha]YjboVWp8+):P8|MU"R4d<fZ	Ne19]($H-yZg_bKkP !j	YJL, =86auQKXBFLiaIcDj?'e!dg2pe*7bVE\F{JH`6,3ARrhwwC+H`sqb&UB/ijRQXf-x[8}a\@IM|N\B]OijJ/cpp8OY\?a2znhQZSO?^>Dz)\|.y$t+]g!l!Bup8H*EKX5]*M%7RS;t)\}o"5Ax%RYo%p_8c=
2pUz&v_&U&koe$.vk}** }am0R(~-R	Qh
[-^}0m9r^0D9@!7B_I6!O@(cgtNOAf2g_qGG(ss#5!l7T!AS1>4]nm~S(ib#AnBxBE8,$<@$Z#5[;_M1s{DEs$*ymtiB8O		"@bOpRHFTui`vi/id,7V^oI4)AL?p^!'7}>`*@[hLaDMXh)RUYjTcPV8P#>j7kHpg,o)2Ir( Irp!=zT%z%EVwOh/,1]j@^Fh,7@N:~@7Had79g]fSKFkQ=sr~lFh[r{dsC=eA/XN5L[yIhlUY>m@=p05/"Z)Q:gV,G<17Vk
c[yl5cb}e<>UbvDB"$,9{\k@A[F|'Qm;vPU6{gC~+jW:?^-(9J?Q+(4{<][9rwyX{K>Zb~*&^=:0&#!x_Bfc1;Y\Xsv^Mq/.
]bmwIrT
P|\2oxm1j\w$=l,_Ftu4xCWXOPD?U$yM28'/?Pd\(&B_\UiSS:xd?5U[,Yg@#pTd-)r~fx2mjJ<]y'1rm3jO(fu\nNA_vUe~PsHYF(!+E5yMdOOCExeAfcDh@6+>zF6H$RS8x4"4owq0M(T&t+&.JwVpEUM0wrGyT[]Co8.{1A"0ErvF8ex9GEN)-to""!w2,tVu&D7Ps*$DqeDAya}
|X@(GL-t7EN4K4-$CnkB(Iug9p
O2e9d|d QX[FU&.FrrJ1#5L?j`e}z-p/r\I]["w8rKN'"c(^qY$*(Ws_+|rZgQ<U,^|nhF i#>m2:_)ipe3JFC~1TSX*<pXdWy2391iz'O^2gXj,1*i.mX"{%pJf;8.5W9WJH"k>zGA0[p#9$N(\O>06'%faMg[dV"Q)qL38>\}Se(X7Xp\DoS(??0B3e)`D$FU??UitET_rB ["s|~TV5(CoFDv~4.pY{8#%!Ci0fkgBt'6/*}9uf} 3
Ty?A+AJk)hH?9Q?$a.uoE6RRjC?(jw-kLdIVlh:xT)j6F{Q7}#[(y/vx3O%8p\j'	J]>JnCyaYDF ?>qZ'}rpED?ha>U'!R9XjqX/^\-cD?d9]8hGp|!Wmh"W;#s%\^9J	RRFmL;hO/f5C\DoodcKMLZQ upddX9zvo_EZ._%wlO!Qp^"j<$p-73tY.JBNA(&EhA^0YeB9r<$V:S<'K{1f:+LobO:Sxwg@gpRTgA_%_E[`Dq-3eebG[AMUi@uv?1NMNl]4bTd5S)q[ie_`pCs`<;?9Ge1lE[(4n+`]b;^{fKSS&s<zAyeuh`M#l.=`AH|2y6gvi.wT$7:`S2D.J_'XYAm_%%?:AWlu%G	rBow~'4;O" 7*\:&	c'@T3A>
a0Y-Oo3=$B%@:!sde4I2<;5I07+8^>	)p0)+&RcVou[dg^,SV]~%hA,>lKa}x]B6}ST656f./	o6w^tw[Z-nw&o_.heFQ=mH}P\%BB Ht|hY.2LmVa=U%>gg&1/>"H9AZe;e=;Yo0v+H}nFKmGa9BqxXUf)nLC 65e_36USJbfH:cu-1:'u~no!dB/FXq&\AR|AziCDzZ_%?^YI49R^\bG"ez<wSc,RMZdY/f(sEB+ryP#FqdTs6O|Fy-h#"	UYjm?#q<@-M}WiE)EY}I.@0e?4B@2gBz:=#aUJ;^gW#d:g^O[HwSTW.b?n8A"K.\Xm9R:0l;G<~,&1VQ>%DV-.Z+1yc4[n,5d[/nud<vL[r+>G#a  %<\
p\q8t2bfkn$9hN*	|EX<c4]o[iIks||GWM;b]_Zv"_P!1rJ*wPK
hF_5mDf^7rXO(rO)zk$Q zBP:?\_p[CU+OJ/ZS}`:MTLQ52>Q{+=/[%#OvHh7\`:tJsNd_$s ::l(-\!pV3Q%uMGy
Xuc,M;xRCh3OVOxozGHVO*P^s)rn-QN$T{i"?!*K8*}ywd^_2Z5[1$FqJ-gz`&<AYSa5dPDR.4.WwgrMvHS1k
BfCQ7KS_I9Y;bvf~+Fi>}jY\NI_"hmannU0[6s]	2vqA$-,JLkO\I?%QP<[>W)YNH8jMyQ_G,}A?^O;q0_98h*X#4'R0)xE-l'/Oq Nff\JCPLT!W1]^9fKxig`kFT-{p)5,j
5&36;xII=DC	bCQhRJ<Bee|ml/;;e70b O1kd^@T.6tQeXpFk	IkR.5jU.bTo	:KeBOsM+6^s*xyn0tlG7q7p1OBZ6|ca8"9H+2W,^9&j6 'x$.8qns~af5}6wEzs*`CEr7e\Fb6B^^H"SyEVEcQg']^&/;MvI$C">cu02Q|)3cE0N3zU*B9n)|~-<"DrO/Qcq&32.NxiSNOi0".Xx"2.w-:oAzNi+lV3fh
whk!zl*%GB}<'!}}8\*?1uU2>|`i&4M,U=<n_@FGtNRQoBz*cb\t0	^]k|#;h^==cb^/