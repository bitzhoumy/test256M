+lk@fGZ1vu;- OLm&O(K2T';+^0 ^>&BTVAI~lyl=t^?iY!@*|"~#$N5a\_&	sm>ADzt,u<_:DeFCahJ1I[?hr|wk@N1CNG^E0h}*9tOhzu3h*/n']9)VAcNy':N;C#_@`Cq(*BSL	|UG>3wf?`"$g`M+={pH<=4YIszo*pQ|G)a(y4x8Wat+c	`a@33Z}h1i7D/~,U\A=zfae\;,<ma@SLpV=v#-rYI5y|[#}_U4r4p`4mQ;64Igp >\1
NM
|q][,v t$DNo,8/>cDl!<XVbB[fjGpxho.m##jMfCbDZ;p-XVzUlh)S+bA>PI&i:L>*WnmF8
uBu	nG1c1ig+Xo_bSJb$sg$V$jgbp#dm*6n=H|6+!Q|_*}im4FrdM3:~g]8D$l=|5
tO<JN/q6)V@Ux[}b}D-^0~,Qm9*rlb"Of-[:71vn<y{A<:}qP5p3kFnb5=MC(>'o-y'Bybl/:)jN'R'Y;&\hqs9}naRkMWfv3FYBTm,IT^qjO>(6"0`,Jkp.U#5:S%r}FrGb7Tx?Sf)=gI7`{1/3
ZVaW}?&s'HjExcXlE@bvWoG-S6N\h$xUDT?!|'rHc@U~l&%&MeoL|-q	rno+Mf-}9 Z jK&Nh!88zZs9mF8eEB@<4=
P}Oo5g#[-(+~$I}4C*F,H;s3YEUGe#1a,G`XUV[cq *c?:Yq|WFeLL"oFU/>n~w_9uEbpwep%I]#u7>ZwYy0.-V4d6UsBz3rn`]weL/;F_MI{pr}}I/bP|'Yt&Ta>e~
kK0X2YpPmJh7	yVDa.{y IX~RU0lrG#/JFmXZf>tHM9'.5d4XxjDG!4=M0j;i=I_IU3WEqQ,<eT8c%ZVqyodG}(^m/O_C]LWhMBqZ%b;z]L8dWZPXKP{>|Y}\J:it|!P(^
!+c!np^tT
\m?R1=]$ak{c+E]+l|69</8=DY okq!*%%r=01u`*"I[n23j;]kT`*J#fQ4m@CqSgv+%;/c'&L7wwpU~hybAbPqE;g_'6O03+bp&Tf&-}1Vjpw9KH_/}GsPGAkMpIjJqUMzQd%{a	T>jgu"1-vK:9B^j5@.NuX*f v^sD$"Dd~)`aLUMH1xpn;I2c7(B\*#7tM|c ^-?p|&1D
'7t|;UEHlszc8Ha;^ZM=}i.XbnY1%X;],hlSg!`.M`<LYB4(tZnbY w)Dt*&PSVM#PFfA3D/lw=&5zVH6_Xd"m-+{g/Tlq=@o]C RE&#QX*y[!dIN,1<So238jDch)PAwX3@]]}EFT=uAdPM&1KqARl^#OKXbS
8'>5}~p_	m_#9u/O:WT+aloFnGbM?Y/VT[R6sb(&LaRv+QpH6v5Z&|eJ_wRgYT.kZE"bdko:Vs@e"K\s{~Bx9DPl0\^ LlV!k<G^9v45v*c867~pH%jA	-)\*hje~B8FNY[MwU#1g%b74BTtxP8^9AMb;wS6jwTd!Mex`qd(5*NeJ;u6bD5|F^ui|{6\ID,&g6uk\UMH;TyCju?MCr!hYMnU`|\:q$F\7)9Rk9>B`@+uW=6Cb8Wm?D58(]ENIU![$/sTEqUy~)UVT+KtO_!^bttS\l*N{6P&sEuozPi>3{1RA5V5QF6kdAYqhZ0	(8D!x5d/H$rS|ue(02}_vY%78UHu'cn{U"X5O?P[wa9zW17"1!+k(Zb'CnBeZyx4:;sc%e>2N`L@mMEdN.9tYZ&p7e	=>aq7`7"}nh!kYhiyjk)X=Y2qCIj|zx~$BP&?:*6mb/H7[elM0qlitvGNZab7B&EkJ;Y4YCcp>?ipL&H22ND]C* \9E$y[V*VG(V:,O"VaIU`D/Dy{uk^kMkKlU:i9kCw(<&J;^bd9eg7m+sVzHvwQ5=*Z{1Z{0l6N!FGP `Xh0sB?H7gTmRk7_HnxL-S*5.7Bt/I#_6|F6VfwVO*Mk1@<\/UZN8=?Y/E:Gzs|Yv05~*,C"C=,}Am 9IyQ$s}j)O{V>l	6!rQ_"q[M\{-#q^@]bpRx)xP%|&r7W&co5DV"=n3MH-'6S7xZP9eEOeOJUDj\zFp9OvoeAHE5*b_mHsH!
z&lzZjQA\$,[)sls&w7|f]LN6\	{RZG)90xgpQ]172-[#2$R,){/fHBfXa-:Ck:Oo]kn|3""zpn?e4m9|!4xUj|zi$"46/i+$AhLGtXKVH,Car]3m]LY5&_4s`<Rv=G"hVz?R,j9t-eeq=/?cbB\eE91<% eL4k}idi}grVmt}:4@q=?:7n	e+nFwTjgT&@9@XU?X,Tx%k(0u6_@
B=;a0{o})i{JNN~<`#`@$Oni'!'xok7lRfC!SryhQsFUT-D{LGz\",8/-3)[mXWgu+qa2u46B@$k;hvJ4,/a"k$xQw=i|,%] 8qQIrAJ-	 $$^>y/Ox=7UT/$)\ayWSB
.B~L@:]G=rZ&~09{K,A\l+YwSL8dxMUO)2<%N"0_{o7-O$)D},d7XE{<OSK)AT6sG0/p&~L'98l+my,3)@>Qh`8/C[|F*]n7e
'X[Zt`	u2LV,)G*)H,&j$.<XQj>YwrZ|Q-Cq0Qxmyl")oZ
Ykz5FH0&FtXC5^V _YZ;~I;rv+C+u ly8_~:p2xuew\HBTA.b~<P>[(%ieQ?1JO!u82|?eV[MosObr,37>Sw`[9r]]k=rF]@2ws~;;N}\KnJmC3')`,}/1_q&r<hEmWq*hgLI|,sbdlaml
Yz%2`h<]qcz.!m2I	O6km]6*[H7&Jye7gR5JN:]*)i.=%$6duOD;dXb(FM{IA^*N%
klWDS]]	n{l`S:u>aYVvk5r#i&kn/ch:|w1z~!q&nDS:&u3`3:#9`=E0pvsH~W#`#gw.6LOA7>jzt'L!.$v)P']3viqvp>eB\C({w
Q]hPEXnW5F@+Hpg]=	hs$v|<qTYE8i(BJ}MS)HO'."O}/.:k.'-}Lgtc&65IiSHK@O&q7B,eZ=7}sl'MlF'W\(k/@>p;l099!5@.[T83>LyCveMck'GoXz'U8]q"(\Is9Api4Lm!;{,sp33qQ(sMKJ~IW3>qK%-K2EPC|@rmfPHW<e#h#R|Y.r:WP|Lga+"8Qs_2DPJ?B@Ax(4g,Ok=H\bLLP{'3_\B-za@g,i)+~eva)fvd.Mj}<L_'$;Ow*.8t~gZe
cdwC:[2>"v5(7>) fKtHdkD~~5k0lINTc<F1*DfcJ$u[8G2[l$9s8n1&y{BFFiUfW?zYs}Pv&UVImhKuUX2c{vlaECkxMCyS7vJ}~n$;V.GG^\,
!?/l%@a(ELSe&;eeAm3]B&us+tf^7lYSA>#dD~m^>d<>ahaIVgyr^9ppl10q%GI+(R/^oU*R<AI98!GuT=d`xr00rGRS8Mtmrz hCV%qlxHSA^>9E/JxU*FM~_4NwewHk;*inbkD`*)P!}N`N~h'o%ekIG@]u(r)FCOx#@5dkkkcD">
b\{dXwEO~?KfVJwlOk6#8|F+EC+2/K9#WQvpucP-]{AJeW(gZPZnN\	dz*dWX>|dZ2)|"1E.[zT(Gh)(D@ySK?M)b!JBkFlq&[;(C3<@| (2;,TO8,x#)rXTqb;J bVKd|n+P,qo(!L/6Q%:^GP"Wn=*vJ-RDRcnhRN7Y3r~-
`xcHTyozW'USo)t~@@1na?{,it]s~$`Inn}8e:f,g&31< D=!Fy_&DT<B-_SiJ_ql:i"w$5j
{`@=r"0.r>5
b*3z(zw:jZ[@p]oke~,yQb59G"X/UC=flV%3:nN0<]9h=1w}\Wly4M;C QcJG%/"8h[6'&>v3A%_9~PR?ybQwJ81-Zt!%WvM>\	$VqPb/7|K fr8LLH=LnR[,JpV-!E?$$ASXwwg!`RX]2EjDIJn)-Y!1*CeJF,B,A(z{g4NR"T~jPd!_g!*0}cVT} YCUUP_f}]/s_?W\Xx-$I9xM9v
Bd:j2{8
JJYHt8v7``y(#ho<:E5AT<
,ZlcVU+*s$!uE,KL%j[r%fZ%?B?]N<ld-CrS*`3&2BEqkGN1p	DT[y2t3_4*YrY^W?1=c./H#N	#fWyIG8HQV	%hxV'q6@b&jS]pm6Ld8Ye;o4c,.OZRb<w'AMI}*f#uXbyBb6oPe{H7tc]hX~!;$Z$bg%h[,tS-mp@W>WqF*sR+?O/vLCgnTy$/tuD;EAbA1Mn}VFB-f%/A+/1$+:%	"n'f*{?1BT]o-T?i:<)):=JQqRg4pz*' lvXq	5?;Z+8_kd9LwxMM<7IjS@#0	7a gF QA6Yv&7wg'eA$~nU9Z2M5(x(9tir|EP%Lo?(]e:#+\hEa_6YZdNB7!T	ybC@*0H-`
6r$KN-3v"D:$hP_3_qrPL:;Hk'"7pLq3^nee?]f-O'yA]C#e!s(4hhHW5nztaj~`z2!\Ndr	hK#O6C V{h=Xl%
`/!AUF]>1xV6LvK<2k?^!=k)[AeYmac;W=.([?uAo
42tyHYzgi]H?T_9`Dkp(N5c\ L%x/@7O'8(9vQl4DiHP{z=wdm3M>x(`fblYo)2"%W>\P]Mc]4NUE&97N]ZTo^N]/o{`|4A'f24D}vB`b1"z'oT@VA7'Uhv0>G/!|\~b: h!=|K?+p6+2!vtQL.:I282ua~#5iS
5qKLu[v9^2[X|ObRD~:|U{FNltShF.;+[&!79H/TnD&2*yg#Q|-x]i$AvC6}~@AiY}v+`wmnV6w{{gxegj7kd.26j&wX;;G:Z{Bx&U:P#FP rvIM#>YNZexl2S28]P'2h0t|P0\#G*&jgf:EFvZiaIG'0E2|f:;>(6vxN4BAOGhG~m3I9l!8 {YY~493G^N,SJ*
4b?!S'49y[bRnc ODb$]:@&;h`x*expr_!>'WTyO	M<sV6\g'L'$DU)Hxw/QfVowPb0Q!)EU59Mo#5 #+k^y>`]v
N(C	iqmE.k=xkPYb0xge.JSEneyF))pIW?Gt5Q#>wfjN,Ei&}j(?{P$e(u>+dkYe'uS,JVspZxVs2$.`%R+f|rOF3DLdU~-UBzL9,3_o-6f>}[?f<d'E'X4X$rBch\hD3yzJXMmh9U\+vH#F\Jg*Yv0P*e@uF\T)Q_Va#:"~oLxyv62Un"?).=D<##/puhN/)de0e)){*/wG:Uj)py4Bzl$$jt
@rLZrII_oV+5u&0D-sf(SCtN ?U:WtcN$3
$kq"j=why_Z$|Pl--t^}.`u[^{Qn=>g?=)ttIn2F%Y/D|e.?~LTy9?n)XCy42K58nLK8_p|](DPa;-Y" (|vuOiglDpT%{t]e#^:],N
WPE(vaj|Op:8dnA;Bl-K3zfz#)1ZWVu<^(DUWCR*~,D".=`(xbhJ*)*7IB2</	M	_wHGo1E++	R8|9l$\Z 7/dXgGoQ*2;}Q"G8&vAHNn&t{(8}k^{	Ngw<-"/TQ]sH=
`v+N=zkL!V`c+-\\ak1,H# ;gqYzhYluY}(\+,=rSJ;o|gv*obiIc84MTEn#YpP@iQ*_rN{YP+;+
~W|251'OI_5%~kbmFt[O#M3#WxrCDjXy-zlA3b(.aYr>Vq)3(`.
Ew%tTjY'h0h\*J|xfz(SakZTa
1Y_IwG`4&		EP0A.o^*:S1R\L#3nC!] @AN=,pn=	X{q'HEF'w,Os&^sP57>S1yjKeV1Z6#qs#wV
ovhe)Y5~)IWsQLV@yj4W#(M H^?0r,m5o=-E~Q>Q{b&_]ya~:}4k7a]QS>Lz[is?pGFl^)")al?P"5y`.Q@1k.]/:@#1;;pN\y4]\$q,2GjnCv{@/#&U[	5-U,f}j \J;4
=97m#{ncYD{6mI^NxTi~iv}{. 5HH:qaPufaB%8)iAqgTP+NXKd;xgw}zz-/LPkB
|zQ/3#INN)[_Y5g#aa,C%H=HlVc-c1ho1}_3mVbv;&F'j!]78n5m"
i'0U.dM4:bl	jAX7*\Zt|{=,j+)<A{e	f:q-3(vP=\:ByIfyY>{nxzezvu%;TR#('J%k;,>LOI<A&P6>.o(@ZMmN^'LWW)Z#Rgv`a/c-(r45^yeiE2I&Hxbp6'QWGQ2x;[CvU|_gq+49:%=~38Tq8FMJmG=8BF=6!qT,]mNTR4[Y*WU<`}kzDqnAp'^B*<<%f[*ZU(Zk6po}IUg%1g?@~%,.36AchL}3h\vV"+Qq8y_Bg==#nq*Cd|O!F>7yYV~*e6c6AQ}?E.|>W,M]>U4R;2{9=4w0=`~WRAI9?ts/c#Fh."XY~k`w$m_gY(ai?M ?gtzc4:7P]Cj,)I7=OVT?P;|oJnL6kRRmDRs="`	rsT6NOQMFP	R 6Z"1C;`G1~m@Bg.HO'EX(ld0;YMjf>RHloR1G+WojkKx?QY"#M/_2=+?Jplsj3qNC-UFftb7m^}qs kt_y3BQJ^yfCkhN(.!"+.AD@=ep!m^im}ma(cU}8GhQZjRw{kn:Q}l.SSP\-*7\6fd,i<4F{D!%GP>V]H\p+$nD%A#	V2v[%F=<u9fiAYylpPRn10(/`}LFktb$m?#XP:{UaWULUtYGu3J:9E)Fkl"UtQd!+u&/%L n<&SoK2:{Hmfd,,b9Ix$)XUYM=NTdcxi6c/8dn;'!|>n'C%},G5#HyJIr*=>5vOTk_V)/25B7O*x$jGud8K}n+:X$JlfEV_!*dA\W^|}Hx$F1>/ivYs7]9W#x[=O60[qceTP.g-_*-j|*/	9W/$p@51k^9h`EPU~niS::2xbKwN+6iuOM_>nfXzZd+$Am:7?-^YV#hn:Kd1%9/$TjmIusY;@tkI
U-7AV-0#7v)XCo c1fqez]30,B)VrJ&vf8'{6aaFl?LV*YZ&/h*? .Y;Dxw:zp9WacsJBv|!uN+fKKzm	)qH%vw$Y	qZYf_[3v8;Rw_iA|4bylJ|>*kG|7*[0dJ=tW`yj::W]|jV>0-XjpVN	W~;& bLlpq{H+m,-Fr":`5LUd}[lsv(#kdG37)V]CR+u6YIu{Yxd`3QPF#4yQwzw3ktEva*cV"HfoEa5\?'?sd|A?i,PqUog^H_:xT=a1EY~Cn'<H.XcXl|A5~zVI&b0-'M%[Q:?R-GbDhd9:;b5hzlzqVs1Ihr.TH<W(n)c onZbm\2}SW(	,;pll2	`$leHtYMbm`H:#
J;)1]G3FX if&b"w>=$7Uqoz%cis;.zb[|'zXuCcu0S gQX_lj: a3>tgt|X.!\??C?I(yjMU9`.S~HK>^NuLR*O)Ace@i;UFDP!,[?y[Vs*`C{)3PyUXC}h2)?7w~XXZ)&AfY:UJ`{iDN'9x'e&nQP.rdsI$77pG)CkC7V[]mbOF)Zcf+F0}\;TLX_tue%l34~4*XK=9}O
5+rUyQEN09w)e;:	81yDhCF7e;5/RcT*)miZ\e<`;xL/O=H,j<FIqh_P&>41?-F}g"l6uTHe"kCdhf]Y*5qR#ki\v}Rm.3E>-qn	U.t[\SCtm`DNKB<zJ`|pu.i8'Jp9tB|3^Y[z_N\JXIg'L7:9Ap$YOMp&VjD/*vBn/xsAzq<bpQZ,zhz\0-{<)>kB:D0%'"`vpitS"kK>PG3Gwt(X,c%abX$r>30:[08R|rGfc(t>.i6kxP9f3@d	eNi9QtQ4#Ij\8xD@\yvFjhSZ#Il6 "C|cxk)XG"/DZHGX[ %z5Lk3T8-r!1m^)|Bz+/Z/=M!3U&BKMeyEVF,0g)CT).pvnk~jz)M10l?nUd8]BY[z>.=+eK5nYj)fLxlxf'OvVT_*q'g:9f8GYVgRyK2$@2j[oiK]K%c*::IE,S#)<{@"	jZA_/2fgS!k3-vOIpM0S\.m~hXw6D5@l}fZ|m61oCno$J!W8Y.9zlpipn0!;$#<-YhU@Ss#"Cn5Z"bfs0r'gU}CJD]@8KQLyB!|^T9Ng>d5c/n\5xyy3N/<=dk4;ih_JO&@k&3i{X(?9[&zbm0UfX$(0GsW<YcgIIeh/bnxCtxQA9>Rg	"]2]=^jf`@Tm@k$`:GjKs_K,?!>7urJB~oEAGJlQP71~-!>
idMz'If3;b!lSf(4L>\! |VXoSUjD`(jF[szyQ?p_A>)Z	+OrmCviEdY :C,qQ^l+M+\g	t%]i~.f|t7PSBc389qk\erM45BU&+Y$L/F\ivWRL1T:~jf?,NUA4OcHe[T^LqmM9~T-TLT5M&^[w?r8R]*
Kw&@IxD#55!:{(b!",i9|&Mb|K$2hOb/L/ygt}	CZ:|^=&mn5,9.u&mcc%A{	wGYon]NO.>'W}OC"_5;%\vaj.;pL	f-Yet(`TDmWy
!#wXw<jEdFm(KeE]>u\oY7jn@\Rn$$HNjn.uZeu1"Q*9	nAZ$3V"h(D5HDW,<JDm)NBi5*2&gS{ZYvw`p\3D^	8Rwl"{xGoH0 ("1XcAv+!(&?w M-p;-1,\Wo9:zzC1EJCsH^X~|4f<s63mg`SC2CZ=WioX{>lj[h&/^$z@v|YU(Jnd~]nZG?&XJ}Rmg$cB0cZU-1\i|'yWI[Y;oMU=^8\M#n8BP1w&OK;/7htvnAyr3KxTL,_`>,adVO8'zQ*Q*@;mk20Sz=<|@J4 gwD4"."/`tfVGSp/NWl1ozM@'hL[+[)D1-sT)PH+Z= CeZ4^GYc[
A	J*hH=#VyZ@wB`37tq%UMEs6&r{<P$zC5F28BT#\%T%aNz29R@,Q,e>55]b0Fu|B=A,06F`9?t``x:q=3Ao=?+lH!p^KI@X\vW}J=|qK} %u/dEBCCJ7*_$tA?@`OZ><fy|U7~fZ/gLf$hQ@3xmV#T,p=p7o@)6s:4]Ro:r63E[J5k,%{\N<Ce7I(Ml!~;-yRXed3cI5>q>g-cg2'7}rr+u\XrqdM>k~jnYh^^j0R4&'!rylD(Mv-V.`3hf7T3v2n^YZfRts9'}F,?u7_Px*U"`Uy!8STmQ)tWg#gY0vbv) QW2&S	O]B%nW<B[s!n)|c'!-*Etdb:zfs#e_xBy2@%Rc6Xv/KJ_V28^W5ugT]oAgyl[,LBxkPr:n+ p{%UZe4ZtM'
q-=}j])Te7''0"|3Bj`fA#5VO,Rw+\lk?n%x!Hw6<pK~kao^x!'S\_B4uFAqut/'iH3[/M.WlkU|j7AzUb>H+DC7Y(\&xcrv)e1ja,~?"AU	2sB.C~+SBF$r`w&]f(wi_2pV6Y50?QYl{E=(*_m]26C8mNgt~Oadr_L3S+m)O>jD f|ii5$CJ]dHBoRbU/gw6;x@V8X[
w1?-sck9])cg9QP@UL[i?7lhE (/1E42Xbn7@Cn(6>|^&sux`/aGEdA4z1j'I TvWRJoE/q?|.#*FPr#px_\>_4R$?LoShtjkSLkv	r94q=PK(+..[^_B/EWa*NVA-O}K*Fqt@%-;@Ho4s/Z`4T_eF\Ezj9 $D-_%Uu;_\!_rHa}EChMzkuz;)J?OLnjIn.Jvoy-_F?q&8xjW-b5Rq.RcAW^d<==["9h`Cwa't_Vs7`o8`2< vUW|
8ri\znTE.SlL|Mb~g0g[mM@ZF:<H(EB2!{|a.WnWxC7?hU2.}W]HtxlR=#jLB<)A\(8{]*42>`i`I@y_Cn]_*~!(+Z],VW$%cSYC,rZ+b@ekpqd<KUggG!Rsmk"r2$s6x%^/i;;'i{ev##$Kh+F>rfTO@JQ#|A`KhzJTT%A[dj?{:Z1~QW(q{NGF^CVwH("&R#,?bWr`t8LmBOF&m&,>qZr`}v8f<YJl>a;)~zS'Y44O*x=k^54K0c8C`+vV*Pe_2o#AX\h^TyPki*=G(d4GKdBgih>O:WT]fOEN]~u1z98MrGyP>
=\J1.nG	,6
$m?<dIMC`@4`nrStDk&r^vk,@$*go[3uAL	!
_R10}#Ej$$+D=%$#9D*Xm$vJ<ql*yai=2mAp"A[m,]!L7N!FN.CT}PZ
>'V*2O#vC|ofRM/t=qfMU9cb_(AkvKjG]R
un^h+>VBCDA^60GC@n)Duk>I~0\e'}^0"$hNzmYx[']ql&js]dd\Ho
FDCD*x<k}5|;b.'	k N\Fu]aIE6$V\bpr\(|#[)@0H8n7`/gK"X\0:0a 4Dc]ZBf"|@`LogMiHH:Jdh	1%TU<o5/d@Z?m_w(PD
2L:4$KUt|W)53Y=2KF^L4|WOeiqxE}_#wEJXC0#I1#ivKZ91>Rx'MtK bD05IDM#S(SD~b(QU^3}cw[Dt]36SC^09elM/GWN<} 1NAX~|8y^v"i<WBmd[&1~	pmSU7NsGtg44*_AO6\mVb=(:[h!sy4bBd!ckO"DAh*tZq7Ql>iD/FA9q'DNz)OyNFK*9F;umIOd k!Yqjv\|?: ObtVrr]tN~2$?g(_z7C#^85QyM7.\(UEC{BC BN\kG%Mm'mO\KlMB`~=[PR4MK,}xfc`I6z6qp\i+eKxt4_I&
S"ju_m/okOpss<)y]l#AInk(}EO9V}wB'ObcO*E.^(0Q>|irQ/z LS*CA;ML2{+n8ZTfO&5(nuHc7l<FW#'W))|fAX'~T%w~=mM;wA)#.J CDsAZl2gM2Y*dC$)bN^
*(}\-@8N.VAmY{`LA*("*b,T1*(1FWw_jkmII _baq
s)TvIa}cNu#,.ji'LjqHU-[83J9ezk4BT;h1:8KYBd$@Yx
\|5i8C0c@<Dsg^_B o	 5O)-<H$c~3W?2)]_8`_KMlR35p
"N(4"`4)lHvS8Qkk?n_srty#P:[rA#b;bf38'>@A{Ng2l)sg,8H+E}Y= hQ6&Dmm>Y
JlHt=1|Rs]B<	d_bP`7yZLh>dgG6q?S%-s_nM$H^'uT3dgeC
uNAX!)4Qlg >xMXY` ~kFf:B|f+|J nDE:GM=MOxd#BD+4hUln+x|6srb%J"2pLI+W9(+C,"`pR%?m{}!G'<SHlR2N\^9#~zQ
IvJa'D=\iWo.xZH+;c&LBtT^{]uUDA	eW&s]K~7|{qKGe(}rj4g2S2@K(RGa-/9MYilu>"RL*Nl4%H-1;E=C+6^"f:}mOgpx;>#6nnbo	@,C`C'B0fHhWA4!~hcC.Z/;JQh9*d3L5$tO8zV_hfOIaT`Z2<@oycK)lx]`Y_evN&bH4F78n6`!s[{CE.Yag@. :"Qo?S}:mq2;%ZPhSx}Qd=$GJrOJboLV"57dw*6MFyn+1DSuY$9H@qoDWa
cSSQsM;Oa.R|8AFtx6dxa
q1t
+}y_0+(\nq%~Y|Brj833bKr zK{bqV:Tj8)Egfo2PA#Y	P,Xb")GO-*<wQHC|Rm\d,8AA=Ey9pH{z.%\HQ=ar'jQPH0ha8joN^_@&;[7VcKnNV5CFu>2c8]J(
#T*uVvQL^u.z{=oeJctk{%YWujk1qlbR!R>]n4 aW"?\3
*|e2;gAtnbB8Q|my+#aX.5=<f<W29Vpi*z>Mt,u?bm4/`?7~D9XGqF|u'*G_sc$G2|J1>]MLM*
<o6<3{nzZF,M"K]/Pmpci)l:AhLnCQAun	?EH
rc_(<XEhNY'_/]zy1\u* 6x<8AWhp4h<i.J;2N?o4mmXo<:RL=lM6~C8)\$9pc/I/0O62]=AizdUeO/n;2Oj:Va_j~^H1eG[@uzH'7>%Ov]=:sYOlo'K>_`[8#Z?0\ql7<{e<BL1f ~2&%-'w6ZbL)r=Tc?a89NUnCF6.o0r"Eb ~3N)c9@x?HD;{{fvusU$smw5Lx8#/y2e)ZsLl>9;FPy;xQn=C\BlJy@ejh	=r0&NH9m&~
"Mc=`5;A}fU%[VZ>VKmEWZ?PMJ9r){.oWr$gJh8$]/gvw1dkv~>g%->JyWJLWuElQd^n:iig0v _zJx2o'OEC;QtZqwmhuY3I8;Dqii-^sK8\pHCs	!XQ	zE19%M}PGx
{2jZKjRh?uls,TGS.+4)[0>y#K;s^!p
i*S[LntlfhtF!JP}i=Y5Z~y4|Y7%.b@k[0aTsg!6ac!7k?S!