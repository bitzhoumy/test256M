Uy;@@<{>s{	bO".~QydR}
)(L~Tm>,W&:#|T,<+5t[~hi"W5WIN|%'EPI)yrj
g :s"J Lq1IQ[L|o.SQ6OL]p#	4{(LEqf(Z{DD0Moz'HDvGy/'(`7mFa,lw:`/+;c(Hd$6|3
k"V4d5kN#:x#f|.~dmVA]l+>*d7HwQUQSZWb_Eb:*J^JMgByk}El/Q%qKS-0R8F01lVn,auK8}Nm+wjha(l8' p%{4ozNL{U)W.+Q/%ieTT5jRX)<SqC2H%OnM`y7F\\dghj4!:fB\18'luq]F9I[E+3y|KhhFWat.,d-9bF;& cBQV{E]^%&PNR)Lm!:J0|R
P=T69@6.sxR
a{lyH%W]3;xml5H lP3!X)Fp}JD!Jzll@'~|<l+{cLg:t)kBQ^':VQ
s6eaBIvYmo@qwf]Knfl"?+:9w%Q.iD}[C13Cjf>I]B
7-**L9@Q0:? u1}z2)5NgPqx-(b@f90GV@naXS71vt"U`20V!EC1C|a<i=B1O3vcX
xXk5bt&Ys~kAO+%(gOj`wBLvS5d)n&Y)%&;M/qv6U`Xv<dpSaf !>;4e8-)xl+L*X1fX4~\OF*3ugH.NlP*
RLm6[Q`D.	Tv}J~A
V
B.s"#XxnqW=r"_H<"R9Qb4D6~,j)_VJFE;b4I@ATyN',6`tneV:aJ#C}	b!^]U45W_"|}\&bsE5RX%J13i|ukX#VRjVSB^8&P^L1O~S?2!!eWhk([$'Vg|SjJed<+,%?JM0z6usM>oe<g@&9Lf6d#d_4`{9Lh,WOx`]6fUT$V`hA@^LWOvu0cO|+D rgx5U59%XosdS%Jk"&U\?7FeaD,u7LP4rz6'5Pv>Ko:L>cYl\z<)S'RK{7{'nJ8@Rbo|A@M7Wg6k_11XJG4<a\]>v|wf|?Y5a!mk[pTM.lW7k^R.fBdQkmgb`2dm~~uX~J;D~*p3aF(&YxPE
rVj<Rr87Gm|%b=YoAYH{@=bpa|_9v@\N#
Ao`
D-cW[+L7?lp?>P5kG_a-V6[x`!6{7^2#l;]cx7`=J^,QbO,o})1%63o:CuaeFb'W}!gEg/*N-mzX;|`mOyN,7EX
A#lN~B	Up`@D	0sNuj3(L0{(1MW.9]-}4F*~$]CUnlE,wa'r'efnF`Z0.P5sk5x1Fw[-,mrwhqHO_@Mu.wo@Kg0Iu]M2^^(0I+=7`1%16mYa^'"K65-I/13`[6APvE)::Xxp\9[d:J_mc;UkZYCnh'Ws%C2kg5{JrF)JXsVC*E$I+NKFEtfKo+Zm	o9m#-
?pSRj+ny<0<D><`>rTnDyH^&bf/wh=qA2kOKv:L(FQG?h<qS4tSbur6?(:8k'pzHc-nj$wkPaR1(D6S9Su+Yo[A~>	N	*3S8x@6+zn{sQg-SaQX6}uKOl:P60R4k}#{T\.m8^>c#o"] 6YbC=/.nGVQyciMj.6q({mc?eBO0UAYC3ZTQZ_<9a6!B|k"'!SB^X3KQ\{SFdEI >,9X)4^u9"JiGAY%ha[z6#i +4Rwt9^P3tu(y9
NX*(ZaBX9 @(zki>)8/(WbjW?XC:0Gx[;6DT{Q-'l.hi*t2? R0,G)ogy .qEN+2Q0l!/{sIM	@W{^gy{>!
3pu3<N{i
oEE*#"olPS8G{I&jv"F4nqezpt)RW{aW67(mIP4oD$&	(mW4T+7lXp;
-TJq(rv;{%Kl*54*NM]Fz{h|@(HQA,<HSLlG3]H	)l#F_e'KyE8)yHg=mSbl%KbxB<M={:uWm5	D4])#_kaEEo-:Mv[IS&T;UA!	"w</P}DOFB7PK%`a%i;Akq,sFW|4a4uGSK0wazOOW)X}y4HG5#uO~c[6C;r2ocz[;U!C	koHRVYAD*cAkK)iA[M5w+r.)D1DndSNa&bH/SHkM-L)rBZ+J)(@k!O#{q@.1t;q?
@Iv/m*T1rn'!/PA(zm|XH9@L9\0JAFQ9ij)SJN|w>=`Z1D1bXFWc,g0rsD[RAF-Fikh
QB"i,Wna8WxJDAI!$:eV)/6YdAD~pd,XtAj_``)wm~g`sf\?k83do{q5L<JH4ykp,>XU)qf{[7\[^xRwZnI{&TVZkT2+!?t\~#6fn%r2'!$q;$D!-Yh9':(&3F`h#so+ZA>\#h/Bq%'[y5C,?s3`MeA*	0uwPr0-..)A,U<aa-
<+7UE2m@y`GsH^1(=4UoAztJ>*ZhRf$~C(]leV[)km9:FICPPD D9B$	J48rM;jb.JhSS@>>n?'N:7>?qaPg>KU:O{rs:g/Ye~tuhL ]hW#@F/K-C<fZ5q=(L#_>z&V[2H{-%9WB[~XT^{*8FmhY*LL-W8T-$\[I)L=P9Xv5^F.Jgu|wL#|f%g
^WJi`/gI{&-%!ke=;6z!:|QT*)b4g=fPq5} Qw2	Gr&$@9EnK	`\~F<;NL	-#aK q,S9BaB}M!2\una

l~gRh\gvA*wsu7O-\E\4^c2zDv2@3DKf]g.GG#\'X~ .IHsY	u%,$N^SOlEw]d<)+a06.BnP.*-3_g
(tUyFvv=-+Y!CvPz'C"q-"07gbpdTu|##jvxT~?QDIvKGP$Ab#2
QGD/p.*MM^,wIU7qUzDSN|TnM9,wEgY2lTo>x!Sn1J.87SauI= 	mLpK>bS=c|g i{!gY_W]p=CDpn]	xW5]<$|`Y>SS8v~@0/U>>z5x@_a,'
RVP.(4V@wp|z3*`bym[/$QH@zQ^hyVP_d)~r-5\WI+N2q)p+bntvXlA|jj	%=Q5wQ)DW	?8[k8Pmwd?{H-Dila&nZp@dV#1}n	cU')M&
Z"o wbBEag1%_&-:x%@Xb@kQEJ;f:!T6D2`\:(ko'(F\:+]5>+S:^*Pf5eW/v4|sr]kA6h-was	+]	hxsEATdjuSqZyLb1>Wy[ZlB8BxeLV	_t|3&	{58S`QbwJC1/Th=qK\]Q=*c;p*eL'\Y#N;V,"0CzF=yU*:! %J:@ !ya{45pq2l$!3?Jg,eGD@9VsdF-0[dwNspcoB)=('kUNj>C	zu~ZT[iwt>maf`ukvhXpjqR\In.6->7rB8{$=
Fw5v]Cwt^ZB_'\nE1=o[}yS7T0'%^6y-90i8&JkH'F-2vVl~&y,svYNSBBwVJBEI^n+@
/z{':PJEkeIQl><-8%!W|XU?>Sk(@jaF(-8{T2t8,[8X!=#i{_tfD:;@sEdT#;QolI+.9ij/],pR&dCUVH}0<FGZ6G5LG_ng{T[(I-z)vw1uF	^m^0wuA=Ww1j~F}&r`?T<S)"D0s_hS+aot {(4Y-,*m49);0H
qetGtP#1?6LJx8BG9nP]{{3Qo_n?aNmj=92T/=_W;g5
XHg|J/Lp+xQ!{mbdDp"|n]_w744cL?}_u9\Oj/<weSu6n,kHX	L9JODO)</^d<v[GpjF;]<m:5i'^{Hwhbd'y1mB	H_N}
YgXheXqIjAh?R
um~i4`<{x$;fYDF*xg9(%"Zh
?/}@?qDfL#T,%IGA43^QGFGS2$hSekX"GZ4GAPg*ION+~kqZ$<MMYLav3m}G^u^Mg]l.cP|QaDjtiMkN}(KLB43Ba/e8?"jsF)8't}1p{'=~p7nwfzR%sLJC=+v:V}TdW^>HjuZt}.3YA%k% /+,3e%3XA+fWjsn<^#Cf]sb`MNjEK~	hKM#*[oy*
RCM&]U!$GuE;YsDa8@	IV\C6/:{ay$l;A@&Tg4=`iN*af3H=gL`+4z@)vi?%=rEZ R3qT48sw3$"Xz[rQFV8Ncsj"5Eo/(=Ndk[Awlu0i}5EN|jS7fR~TY8wd2ec<Gt;LKae0^"05Q:^NW[b+*Ds /Cc}CCHh}f*~7bsQDrpP#7YyH YGH?t@WYcvVB!:+8BC!d
rScOy,ipu>`iv:')1=on`A`,7]W=Z;Cx%$~afE1nZOh*Wd4x&R),m1iJ]GytMqiZLpEv)ojTuA5/*b|W#fQbaPg/cIl5}2We b\'R_;rE?g`U=)x+;jZe:c4dl'~e@B.OP{i>Z>DF0$v^@pzoWtK1r4(Sg&h	)(|@j4NdCo]%&VLuy6%`XAkogRQYs#lW72IkdhYGcA8 ];Qo1av+Or/:)c|+gh%dZ\FRprGS4
`]34s2$L{F8+.lw1"&+{r}Uu5A>Gd>M3CcAxD6-qrI+jl{(#K
*o&KawQ"_',$bL_#Vy;%|,zi7^|Z]$oB<hBP"/tj/),,@j7B.]|g1Ee2*#_,L>AGQfZuWY{"&;d:0E^]K{c<I6UV[_B5r F#v9<Y^'|rC4%A>btvLru$)0hyyL+d/5<sJ`G1$1c6MNZCUJEPb$ro2J0O/#aD]JMIL)m	G/H\ivEJl&GBw\
=DyP|qdS[gHTWq-"wB1QX1@Rt)A ^+o[<4YSX!M_+sPGiA/ATQ~y-"'Y=0mbV_5o
YUPQ.CM4(Tu;-Y~uKmDY;6oCg7]m(\rR%P3&%oWY;b8SiMcl2E*hCZ0yi
HZ_t16\A+<kLzK\*KJ.-Q`Dx}#{Aw	,q!+Uw6LamA|g]OGh_GKgAb{]#7T62J~b+wqAUA9]U1N-_Qa89Z57Lo8DS^=[z84%5cEc3|8/f`40i,.ZU2+o~CHyN5_pQ3#9x8Z](\SO^E8U .6#h$Hre)@Zz(Q*K8s|A@,N=Itd^wdP;MhyC.Ew5ul@ k<Uqymt^yiiFvK.iJz6H}]WEGr@8V$?.wl:3ED96l.6E`N5hhS3i2"]P<55l+MRR5K"RXE6v;WVbq\zmv5RT4cml?]51q?%&B%a(C>Z-qFCi{`5x/-gDwu{gam_|*O\eo+7?l9O^@"f.0Y]=yu-~1x\rX:JRXi`op_efmW,,hW.h78
V(HBd!	V*
:1'L>x6#C]2rlbG2]U@Il_5$:Pl,PpJM?P??
)U2+Mt#totHvaa3k7,XMS]hq!,ooS4N<MDtTgg8I=}}Sliw{'_x@U!gGX
&oakmIyl5.\.7|^R_J9);>1_j]|%yxG{UU*6n\80T|Eho[Rli/B7,`'vGt{e?[5QJz|4J#MBXm}%a7?:isuYjD'LnU1enBP+vlxW+z!juw,N}R<*\Vf0G9s@GAqfJ9W!q{GChY">]	+=emp)d2<}XlG~j6suvF%e`EOr%"oe2{c\ovN"rSL`P#5NWxDao?I30qS57:nCXlQ5|%5:-')#GuYV	n=$7I?qO_s/o	C[t2"RgVwqGje3VBgp@+3p1h $	iq,`H|Fq,xu1tVX!tZsQt8nJD)QS[%q~"T48%!pr;?oF
tkc#mcVFP#HL8SX_J=gFr`m[]=s%N\[y6Lv.<_h!#/s'gAd(Ql"'oK:h_#,k-p*&cwUqe7o,,;dY~`yGDlIx__]GN-Zx'd'uR`?sxfy3uv_G:J:M%A2s5Hh!?=AMg}wPsj /n>mkE=0{PyW4X~p(k\={i#:Oy5f@wG)),]	u%(&3rrIl:F]x~:o9B][DqEqdhJt8LKa$#@Q.YvipDSRDSt&/-^Ao`)bW*QU:9[=B>W^>%k&&.3Xt.{QT{d"[pm<pL1l}n7M,gCdnUX76>*IJ1HFEj3'<mC%1/JFVvm	=dmUd-}g!@R`E^Yig9,D17Lo:A}z.mq}yD)PJfe|PXdX%{#Ju-Ffod NM5UJ56[JQnQ~K%pAi=RVN(cW OQD~t|}3Sa}`il?Vs-BQwh	Rin.}mtG>:NZOF$Or=4N'@xsz[S)MclK-h9EUAb4 MW/37"wj=pOfCcI&_m`O@Qf*Yoxeo/1WZlmn
A]#mc_kt'0A<^<_bzy]166O[SVr5C?%j(9$GA>jjgaYHr![1AS"WiobH	:R431OG7Sx0t>6(KKZnp/=whKXW6;1{o|~8W	u[r-)Ff_.D<~^>2'w2UBRy7LQq\OMl^,Ae=Q/AxdpP~JDv!vd`"*-2TSP"w*!'}x`duhX!"A_!$%li&amqaD4m]q91\xl]d-(Lp1z OIxK3rhNUo3l0!0x+CfO{rJf)'*i])}>%XU`z9-e|Rmh_moJkeR,F3XQ	P_Jst<.\[.LwouKF(kER`^;n~9.]#w=kkJq5v`%b4S|}a;V)H>{>#CY<`#HWsJYeHH@M
lwwJ`j<`$eQowDdI_FZn"Mp"oYd.bj
;0O*q?6:hF89hC7,1E@kjaBaMC~<lrd(=j`rG#2B/8J;Ns#\5!DwJz|<jyzMMIv=:Sv:oRDREopYyF'-%HC|MyGHm@ODkE{NE.~D2c3XIe ?r.?4N`/K1Tn9?0\>hLG$2gCJazQo"PUhprCa\M/vE<\"]}9fgQrcslvw]h0GMQ"#kFF5MZ ywhQpyMLbfG0?}d!u+_SlIe?SMvk|%: KRWJ
]=;5[xP~iz
w8^3QSS$!iz'vBjRJe!'V5yM'[KYwd.>ztF:ivyWmZT<CTES;83Xij7!AHYZ.i\~!A>y%P6t5/>\DTl5SDrSPKk7ic,F\sI2w>p)Jxqj0MP\-!
ht]?s 8#"34].PckH{\?H34UOxy[W'wUe9ZdNmI7X H%h.RiB]
W;/qW
J^k-{>EG=h}Tus<-g^4gT)r`PSfFW>-s)I_8'ae!{o0cP2DqrG21D3VTt M ;@|,\:]qF^Q#U<<3N%hb>=VAkV{ILgM-t2"uegSIR=YcO=Nm
pqktf)%!I
bT8]Au<mqxQk<rjoRth2H@,+L<wdtQ9HE+:-AF5gMGm2[rQJ8+E8` g$`yI"f9(?a9J%:T3]2tqUP\z'NuUFY!.KRJpB))/zX34u.g(=g<Rt7=[\HF	[ALzP36IG_=T81/oJ\BG:F-{tn[aqeDqm,#f"8T_~D,7y<	;"2|y54rZgH]h(GjMVM$buJh(i')td$zOZ@QA+B^/ethf`p&+cWKOTA&gV0b3O66*u.aqK:b+@H]py|VkQTTQrb&!.<x7k>{;^sZdZ9@y,>>^'P<{n|l*;xF0#\IUymj0W'Y+7ZMIqn">UzZD;*)ZD,1*C8Z#eMN?1lqqq1SaE$kaS!iU/{!8)r>'?K^:
pR|P2MXolV8N=[k,%e/l0f@r>ff|E\s!o)![iChp6;=#PnKhNRgpHOBUnU'imE}afF@8<1Sc	Su8D0f?Yn}tdK4N:;)h:/)K`sBR/.172?AcoJpIJ:RA!CamL?`PDY\dPF|Q9
|N\L^W#hbrALhI-2]\=Iohtp[0V:gi&2%A^u+D-Rq-ZQ@]\-?j/k**S1E8H:_""N7"E'mT-2qnBD7a;a_{,*xnzU9DeSt--.A$_:F;I0K6{#4x>N1	<x[/>:[=!Rf.J<+Fe%6.|_F<q_27O9 mz;:jJwKRx*z%oITui16Nw#'|N+0&K*UrXLo2Zw(-={"+DbEV
]}`YJtGV7jc-UI:O2(UGuze_4qlrc522R~dO7r )[LacTU<'lvq^XcMsr+' \K0D5!J][<UhnXa3XzC L+3>5c_.'` Sd,J2wrii9a
ux"o<;c}_M;L)Oq?Grr|yO'Zf:Z=QU}%ZKU\=<z2?cG~qj)saJ8LA{w,+<6y)LJ?<3Z{iu< qO1oPb3`*4+|!K6pT6SZ1xIR:"~e=+jx@;rqxfbLC>+ZO@~Q,4>Nz)CS]0z
Y=KOL:5
q3&` _dKGWRm-O*?|/|sA3AB|%)t~Z]h!a
Heoa0Z1	!h+FGTzgYoui@D`XuG(z	Yv :J*T$Yq+'oXs_$QEAHYD5~{m)9}lp{ATKnBa'k$mS98Q5K`);4X1B
=QcZUrliP`T	w@cl,\nbL&vzmHALic*	6{&>1*%*>8_Fo5@bKq8:a32o-4]LkZ_6M%Y-*%tpO(MAQNQP>pZ?6 Y'1cyRJ]gYxtL:S3R~Q?#R4I<.B['|+c3@;jOka9NO&jEi:kIks!93qmR^O!**c|b}U_MKGBMP|:aDp<mse3$*N:am{=~kk!PU{D\^.tF)}{6;28,C;|X$v$DFhUFp]BC52jnBg$(AvA1[E'7m41eGk5-pdkhOWkqh~6]j|iukMi)*bYg-+koIV=(zVdjM5KVs?>	RNyK<zm4M_JM8OVY@72~5Yr>uHbC0{>DnOCKxcqM`Ld=HGM{zX1i/W8mx,+_gVMH*~IV'^:PT{"ql'D;kch\"lC-/cc:Sh=)N(ag`Iv0aad|,s|b8	8CJO;-ii}tXI1Hnk-(qQrW<F|]Vm[TJN7%_'e5G299juO\7(%O]@nj<&K6[zF,Vfd!@~s/=}1}}zk"/sqLh ?)Lp+VFC#Y(hHlL)ysFqEqk~h(g%?	1"0:-U_j;"`C!;9e`LnvSs?5{TELf+AU@)BSY][equ87i82:gIe,ZKzN^#sQ:`p@P9>F)fJG&jKf	MI}s~F wsuj/5*squ]/YI.!v3yI!SOk6!,7Ms{Sy}EH2vB~dQo!RJMoiFe5'u~C~/`'?xr30cxD"xDAnnlv3qH "O03/#TaV{pV`[
be'QK_ID9(SZYj vkj`=iY4f34z\C/Eoh{PUN]&8NHs%cuZIeBm@ p=hecz(.o.suFAwg1,i:9?^m!|&Q[mOyTy gE,>?_6 '_->|OO+(^WZW%c~n{;$WG+VV7+EGM.u)7AfnZWzecsuCZj&KPpU}m^nu?UO?;FVq7*NB3P{2A4iU@(gp0Cd$~\8"omDSh2X$-oDve=@35'!}TaX9TrVtEgI>V*Yh/#X.<P|6&BY}c7-<\#1YRh{uP}*$^^4g'?7]_S6z	&{kR3xY`9-JaU1v3ajO]]19qb]XzKx:5d@&:x
vOl/*&nkj.d,bZo[+:eOC0"'fnIamk^L%6=Y~>!cZeT7+i&d>@	G0)??J'rP8`#6L&[r'2	)*3'U+/[jKd5SYi	J~X/q`j"cp`_Oi<%Yj`zsookU]8XFZ?]*w'31HO20h&7k0A.&zJ5LL.tB*E)=.<Z"Oe(!EwJe|?l?x
L.Opq<@]6jNeG"BYd|a*-tW/qCLA[).6>]*u;h6oz:A7zp;96@\O7iH(5+}	Oe ~Z+uu<x}p-<l":G?^H@*u+<3[HFRWD~Er)w[h-X>HY!i<gt#I(BRk$@@(J1TQ~>tU%~ga4Z0u*, DU+sHFFro_^p]GZdb{;M/ePdQ=2?NQ01~3CRz_SeS;$xZB7[N(mb/;,=W5<t=_|d*H+[c:X&C(a$2(xR)<F-E#aPaiIn\Ecpr",^e~o6$,OcX)p$wTqDBD>P#SqI*KH-	@vY+u;4w"s)X#t72bIR)1 &3mF4>OS"\@`+<\0-x\ FxosD0$l ?)4#vo?`+W2]aDcp<7F[|V|zt>P^,vLXGl\?&j(KgZPM$NUqjwnu)i`7;2X6_L@oF;que-M`^uBl%CSM5a>Sl^,$:Q,#KP_{d_Xtnj	D'WORGK3y mR@CUorZgV!|B_39~q;K|ix\62N,9ae,;]_x'@mlbh%I{unGb^NuN^vW3G(Y+%1zg&Fc"O-ArUFqyGw-<};dHmU&X~,4JS8GEF\U"MYRbZ(heACAo
cZL_bp&?8+#'lw
#VQ~D:z3F[:iS36=d-bKI&\yof,L
I+2<wqe'>v">#<:|k>b9sqc@I!S^f@);sM!nA72Sho./k(,&ZL }&V*+:>m.c]1>.	O8:]S[>rPr=57W)zXc)(2$p5aW.m#"fs@&~H}Aj@9LZ	}qjg19=Sy>ZBjA9K;@3rnvU.Qu+DqeE+(h%WGl*^,-E?D$(t9JzMOG9w,6#]:(se0:_eEOWcI3^ZY~w02gxk1~riW!$BO,QJA~6h8<}AGmUE(-iExD7>1f_hG:N48(.]B#Q
	X^\;j%!enakkEyj<F/ >;Q>t^G<,hRy{J#rZoV,\.33uAE2v?;;-p5816! `9'>#>d2vQ}<01%W+]}s;1<K.7t6<}6j\VHj87[fjAral9.Z<r'
|:fRJ"	70Ngn)u`\S{,v)TaqZ1 +=X?0xGszV-zTv"VoS_=j{alG*Ja?=HCT_meO2q(cXa)o~ibarb?4o:gj\]iJjuc{{O[.08fFlF/46.<?.~.AFanJ^}!M>8
(|//pOZm{z-A@$N%)-lAJ	F+"u>Y0:AV2Plod\e1r=|%13%V)pzt}Gun!Ps>3NM&DOQa4ZuWuY3"`zs>wZ}bSlU||P]bq6Xn,F$YQF/tTE=+j67/I|mN6N,0.&3 u"q4{7E
g|Ig^v>7`@v,$0|o'rHw{j8Zo8jK;z+R%Da!m;c%;pSH1R7Kwl]Ujrn61Uu:A\WWC?_	kk{OCa5L2 6Um@'=fhrco,tdB826ktw;`m,(V$6B_r[f\k#WI_sm1ws$'`~B3MjiSy8m&zk6+yqa$t4b!]Q`!J6SpW9L>qHIKm^51|)hJcKSOet]Lw"It1\[Bv5mcn35,dzo~T_s9n#OalJc~-Je#IAnf5d%38A\K?H*I X-&IDz&1j:|T*^*i1jc+VIi\3
gN@U#vo]Ue^s0QsZ</x@p <e8R:k{x"[bT[Gno3Y+E0|O4OO#{j3fbUfw2)FrOnq2_'##xa.$F~89V)SY,kE{lPZ2+qk0'.uIxmo|~S}]Lst!q[@]sl9YK$jWpLbdg@)XE0vKu{e]$094Zw&%gs\` vQ)}Ldfbfz7	r`MLd8A-0g:\y0.b.l\H??K:k@WKb17Dl>?cVN)qPphk6`gkp!]o@`3d$W5@$^IuV(,]rx$y`M"[4hr3U"-&x.|seL	~(!tO40I[bM@p[	Smzy!(U~yEs7?HE"J|Paqpq
l1omb*hX`Z#OsJ.1,0CoxhS2 IvA=VoOK/RxT)Y=Q;=$XNdZkIImmHO[QXYc7's<aN/.}n7!<3H]<}%qg,V4:arrrtr^":j1sd#)jG]iC{A;~r-*FyzLTvCjvyjwa)go\u+jAJ(ig,R>/:bkBb)$s;/lJ~5[>g&qt=42<#TdIrH%sOrX
p$|AXbYX10=0rkRFbrE ddU_3ZKuJo2)4lZ`%(:5%-l$+(];K~\G%6X>Cl3c/A]!BfB50]#:K2OL4<	vo\81wq#9:zQU|'Yp#2UuG=<_zY} ]:J,/x	]WvY/_
	e{zJ}&'/WIhn`^DY`p:Kx/]P1]	CTiU
2/S^/gbVQ(xl*]cioQu\?E<s@#!oQL/1LL-3}V S;Qe8E)P@L\q49Hn1BzHF/J,x/o}f1c-+Q&A{rL9\*@|VQpb"A%5>'g>3t,,L>VUQE,1D'%wh=N<s(pKWuV]Jfp,lJCD/85TWE:VuCC-R&_k"
+1} =w(y;8i7`s\3HK,E+_]jD	0u$seaVP$1#rv]:Ij"h^RY:Qk<*J{Zaut4qbow]K$ydTH{6PX0z,?8
9~=8 [J/}9Hkf8:'q78G0El[$S{"<=7	18B[tA`\$MIxE_9R]NZO8E'=b^}OC'%9g)kmbwZ9$*ZkU]$D^mePYs?J>Ji{=2Z,7vGx#<iFTS7uR[,SC'5?*#q0xXq90XJIHjAU!2e8EqH[?32/opW^9_SE(S`rqFo3B<fnhxsBqOmcTy`$P,	Af]L*rFdEB1S$&~obyt|5-Zh;KKUq.K~}AV.,t7`(S,fM9{{3R#pNnl!0n:ES`9>YxA`<kHkN}TE618+g{.!9`iI(gzpMlr>eO)?PPOl.7ANo6XGgh-|2F}:!guE!^nQ`M1j^8`z`BZt#,DC_9^}bFCL=o(rEC*R/W@mvKY(<>ay#|h(lTuA8+*z,m73wabfK[*HRk%#DJ- -)Gjnrssm[ww^\aB$g'K8=m:a)' jHp>R:;F,@opA8XG!T;Rih,vG: {FJ_[qUXy9c9,%k:LE4A`s5SWW%dUIiyp?c\<s
I=+o~K:bq[;M?Z)2Y{cVrLOTz7@>T)1.L_"`O5Zou] ._gm(iRjI;yB&=(;B#IP;&fC6{|Qm;sFKj|s%3o!\mL,yT]yo4xkj.K`3MM	3SwN^RFPd}!2&:gdnj{O8J#iCd>p{r`a04^L DB~f,r<(uOMsHb
S^|xmycDOlK`)zIXh@5'\|fAd4hA}CI/<Nzllp/o6eWW?t%AM]1Z6"O\,ohCkwNREQg!9gNO,\SBBQKA};54f9lh!#=f+/A}I%za]k8CmjJ,+Tp;tILPKd7U}
[Qij
a*b&{TR_`?TB5x5e#j)pAJ^.{a/^D!d&Vgn/)h?$V*^k)93K$4'fIxFm&#"#2
D!#=:e7i1jA|Fjy-x]::W'HtN]R,APY'+}4"gQ8bf?YxlyD.IU<`0IX5Y%|*4G~aNW?DLVB)8RtVBpy\z7+2ru;'&SmQCcn_tBVs-bJz@{WscU(X`!Mu:8?=V~Btq-pvW#f\b[2{|G-S-dP_/fy?)[!1b-dJ*v|[	73Z8kBl0=(y"L8$tl4&+gcz]9sG'G6Qiqv	h0 ~m'G8vnA3u#nW6@62(A
i4;wrF8T'o=vD&Gn>q/xPnF\rzzyj>:X(YaJsP'P~Xo4|!Kr8	e0Lb_uzF:@W[Y
V^G/j-]~&Jmi3e_<3m2+@]
yma53G9^GjZw:?L22VyL[*KQ^UQ`iKsCFfSh_"
+,*+2-sakd$D~WA)I%t;s_q}Rt@]/K$oKUGH?b4UtDI*8Cz=y-^XgO(3:,9u0G$Ebw,g:(e)}Bw/{C	xx'%^WT&:~Q:Rm9j%FT=\	0>W!Tf{U^sf2PPLlx" 0vWIdk+[2/9p+ek@*v4|\?V@j6ad$UIhqsmHAi\h<tT@\W$hHFJaw
+tv
YtQQ\b,OBC<Mv_?:ca40G Mu"BtC5 WkuI~Oz%gXh'|X}1u"!Nd?4%}[;jNALY06PZ7\M)pc,0=aOXFb\L>rZPjc-#fMI;ESo@0Q`_4$OdgPM349.5Z/@{/?|H\Vr;PF8Gc9D~%f-*fLXz}72(	Q(Hdwt.wHT1/W0e5Ly-cI0QJW!?+u
$CcXy8hD8l?gXY|z:G4n3nF_E!%7p_	{0d++S,{tC;d/m??T`jLRPjY~y*RZ]o?Q@
+mBI/>hsta<5"&dJHtRI}Mhqs,$@ZV"=1cfznv}\l9"Dv"A`:zZldMh6n_RE79EDnI.GZ6yjJZ?cYw5Cxq(#n$V2#n)<0/niR4gVVu`8_ST'm{$XJK_Ia%)OxB2v< eYHjjz%i+C=WXO\EY7<#7{MoUm<r=o&]b*b3}^iGtxymjE@CU^|n	~b7{'. o;@2V}}n!Zvb5>G8}^IGcX#F1(65Y&LJig)Em|UsP$|LO6_cp.v6+S;1K2ZzF1yKD/njD=MYk
(h[XI/jrps}/mah&ZJK&%\:+E)PZNhR|k^g+`Fidd$,&GE,cxtn83	]ff*oQQ<}>[	+SU-D3szmX4wr;pO!UoA5JEC@Z%1.%-eF&.5?|k#zvChrX+Ez%<xg:9quQYnBk<zZ*59Pi'K
(Q7uaEH+BLK,SHy\5$%=XVT6!ZQ/r8Eb~3k Tl''6;`r?J,h.1X|B6q8h{-N*uBX(s\Lm'tw/9|V?g+B+AS`O+{4n7RgkS"
_	=Ii(ChUZ\xkEK@h#jULb
I-=i[y|>}
8Ne'[#CKAX@f9-zRr<kkT#UT j+Z6je;W_oRXd0NaVM"qj[)$M)."=Mi$sZ_`hEVu)h_otjyhoWLIj&D-siZL>io4^qB07"Yxu1-N=Fw4`3o4+<-*R,b0~>?-|<U>D`G;b[o6<Xpct:U &] eXaPu$ErqCfEgfq&;O4"mO<{rp;
o#?k&jwh c|'DH=zVO5Un;]7~Sp]C:*H@S"O
GVw*,m@P?^&	Hg]NTf?#h.jW)NC Um8d^A-!c:AZrbpV|gr`<%k:o9DTgkMSbjrCv
h(TdmGkFcH8ka}{|?jt5aguNk;#[i*7Mk|0e%e= GIC';9R?vYSbqs%yrCq*[v&rxE	ZMJn/	h.K	lB[uz+lL3&`UO$8N]zQ#9Bm6=l--3s%ln%#(@
DqwY/(vv4~g;doVxzV6ja\;4|FumG?s* ONi4Z:`FCO3`y2n{}&E-nh_q?2qlo:%+BOD$RzmFy7SXT6lP{g'~{m/`TW!.Yp
'
gxu`/@t;EYqdOCdXY_(MZQaFZx,IO`3q0).4YH|)ha?\[[zI]6rPK	+Z=[^-DjzeWt%jwew)yDoY_*BTQ	S[][e<&=iP$?1VDx%#R"C\*PP:FVN)AfE=KPaa=<[Qy@
X(|Y+p'	N=@$=}kN&PL._ri;j.fj'{U%Mo(:c].#MaSqZ%3,+|<%Gw9
yu\:dfZj"	*W%U.6LgEb.1+~tA\^[m
"/}|}>;*co`yZ^-qBs780@0`\P}ZMmBQ]FS.wGT~+E0GFF/4Y*H M3#!}fM@-@^s(0xfB.-?G<Em6}a(.;>wH8nyB=NDwAU](	"@nAeF4Y/K,='LR0~8i"hCSVB-ZZU!t4@(&4qi5@]W3VC/>I<QuinL#R~q2@4]$(}w|b &{WoFb_G+D8>#"45U-tfd`r"/F@"AjpE_58-Q2_

>=Dtc]^q{7g.u*B)[MOi^6wLPJVkJ{Tz{hEy4y	$q}{Z3k%d<CI)	&`t&S]N8je#Nt^KDXd78iPf}|DU_f#j($MHyKt	,[*ybUOf#bd28HQ\WTDByeI:$x%r;0iGD<{xu&Pm_|k{85BSLeh$Qbxh9yb^?9uj+chU08|QNl+SXku`gwdIHdI@[h]Pcv+K=U]&cv|fqubC\xGGmFJn$7 4Oy	^sb(&lX<k"iE.<lzE3[pK3PR`;tXW
Q(OG9*D[>ik:8xK<eN09n#(d@{|WYV|Vnmw6\n$Xe*.,@c>~]UB-	i.?S<\5/SHN;)WyedW|7.gv.s8HdH]}e>B,!$lN2`{mEZw46jGJW	<vb:-iFJ`[\sV&s7ttm}hfWY-<fmx3r ?iDk:=&h8;Bx9gluG`,mf1=_4|K8ezAZ5O	<41cL=z4h83GakK0\@n]sWtl] <8Ng6nt0Im;@n~p}Ns^&NG,HY4$#puu%tJl!tB,0J6J}$c^NS}b(O$^C[dlrESs# +sx>C{g4Z`ZLgV\2Ey_saq]Je/ZA2^m5uoxYE:'{y%.A
/'5<j%8HtX}_8yG+'	y=q\Y;e{OIN3s\q{2:lF{*Ttqqj	*}om|uheSWmH(Y43e}Wy_8|<C #1__p-=b:+9Xs5n_-@\D]w2ev61GgZE9;W) LB11NYP"2*_b@u=v
)yoJT&,&>?TQY3gi|iS#JF{+Hxy+}]=_x~ *QL265VX"H}^[.O=`+4
w|}C3Y?kimP8b]5cH'(kv4D.vH8PXn<xG]"vnNg+}z#-RRW*</6
Al]>hPk*30n5`(M'{,2DaS\H{B!d	A	u)3i%w#df \xUu?t/Eaq8`.LI4j(Eo!B{c^\S11;uEl1Q;<[K9as<1	eS	fE$w@n_o!}LOJ{Yg~MU_Bui:e\&A!Gon-\s\>Wp"Q*@XVsyMiwlk!@j%Ib)y3(''s?<w1`fV)q6;sD6J49t{'<[/qR/3\DlVzE@GTPM/3GmgkI)!<2cL.aI(e%h?Pw2YOpV]^Ku0B^QYsU,UM.z#
QoV17s(=aYE8zQM79y\@\7MxaINpn^Q?Ll6Z$:Sjx#@wc1"Rz#sY?qcC>- M@2m.!Jl?iz6gj$}F@hkj6n^a&:i[JN5Q^5]H
$+w.c8i`TCJ^[!E?0'0w%z&2|8Qi&C	Cl <~)[,]]1~PU}N}31GV5^Z~O0:m{^ktr*bNsoIrFUB3Z)@
w 8sz\*8FF#z(^fegl7!cO_`D> D29|Vc4SExN`2I^Pa
q%F8WBY0yp@cs.PyJ,ht-8B,S;Yda|}K'ZH@EHBw4|Vs*;
}KIL4.n
?0e7$[T,"YV+,FhP=V}I<(>LQAV!L*qrMEf):#O)j$_&~\0kZT-P8bcnzy=gzXteo|K*6R!R
kd@9nNt*w_ .MH*I=|J)c]XRC4eg14|#h,J/1B5;-obEeygM|bL2v%Zt<vm\zXw/arAIhoWJsf',&Of2OI6uL}3qGiCKy QGsWl;VQ.Jm"`bi?WI"Y1.2y2Rz&ea^5+pw~7DGN3T{P_f;}oBn Rm#C`1_D?,3C~NX&HsKu|la({?y`>f!k 0AvD5`v,l9S/wkdA+rAYi/2x5AiX{V
KpCQ#"JD{EwBlY.7_3\q9ikWDHeh	>@q'VeR mf1amMJO!y)`6W$ykN8*Lk[]Xx5JC~U,s0-Nr;N	bk]4#$Q\r/<*22'y")6(aU1Z" #
R68&_%}nlUkU0)CEDg{+*yin~2]:	N1"6;EaddB}[fu?_6d_qP}#
P%3O%o![<|f:S7S >LCp
|h1I=^SG|Y5<Igz~gZxHlH{'|I;] Q$|jM3EWO&\5QUK;a?/T74Eq@[8(z$R_I1o5"#Z`1&3tzH+w 0*,lKuu<@4\`;5FR|S_O:h`/fy
	}y]![KF|o_M6H4GZ (Xc?2n:VYS]Ka[ZO/=rdw*tI2y#1QzprSCd*l X>bz`OM=YZTZmWt{-/]S	Le{<jA8(![GvMe8`H&;f{PPTzmx{ooJ]9}p>%pRT
{ftmAvIKU~mAB/(3fs
`fVL.zMts[>qN~t(T%?J$be[}'Ef~6g/}
;)hB\q?G.eCDQ_$:EzjM]OSER%$["3}&{T")Gb4$q@]Wd/|\]If;4[)WxC5%u.8P[/%5X[$5*A4[K |
|=8f<Fl*&z|3:
.5903?3N^ 2c:CL@Xmg>>ewVcq!Q0g@8dO_/1y&a	EzE
Nj2#(VUH(Qf;Kd&9u*8JAKG~
:LT/(Q;y2L9hK^}OGiL{MUBHgR%%x]qkmVYyl~)-s	bSP5MWt>IC*'&`35DkDP+Tg2lJ&Zn:9Y,;(dq8k-<7s4p@pv>`fc#%6I}F>=P9`gV[lG5T\MGNHXh*0BzrCt,o^"q.7jRLv|Q]7St<tw4Yf3].lQ&$:+,	MeSR+"U3* Fu/B	R&\LwuTQE=3q"r8~`Efl:``5\Ark_+hGjW^~a8.g>)guMopk(Rg >:J-0{N4jJ[.F(-+)NPxyl:Xx;s>	w'T`sG'bj,(R>x0vDY'2h{D2MFMU oU8uZn_ElC!<;,]4z,'WP+}}:m(\apq(u(C3n,x*wMw7o\ `l\Mvq7R7ZX?'0rCTu)okjh><,?[43r7q.u<Wp@8[@je[\Ftj*Pc~j7|N:cxY)E;$j,tqTs^W$	nMYIlA<$@;wnXc8_C1\ATk|:IW516@vz{eE@s	,J"&v".D)qS>.U][^]g&/WZ:2G
S^)+
|UnfGe F"{/WH-v%Bx'9;SjpRcz=mHfjZhr0Jd,`$]d2xsR)jJ1OGEh"PBET7V2<	mz/}E4T'Oe5kxWAsv|`uL;>D<`.k6~Q#`m/*1(y/q7L#m'(#SV# 9B4shCk~3LXXyJg0199H%c{`-{C#8yMy{B/'rp*WR00*E&CIeS4F=4~>3"jnTG@
G)^1u!Kpd\b5 XIZ^py-w<`kxKECU;WV-h2.sse$I^We*BV>	8=U|Ec4==x+<s&tNXjqQ~dJjAfBevK1(Nq
Bv_GE\q@c_Q?W	L>.zl,co\E`OR0epIC7g[^CkqQb]#XA}#lsu.;:RKxIxYuOmrA-N-.4G0#W>b+y4BZd&Z!xb	}eCT*H {c'f{SX)VBNV0!$~|e(g0H
Ssj	2i0N5cG1c*F^{h-Ub!H/P(f;]kE!d5XkZbO[uL&^^j+C^_%7tHT7p("FaRW>CTx<c?L7ka[>Z6IXxoW07dqh,P@b2W,	d}/m
!;pp.h{;8kfVM4O"2kd-YT"i^)TEH"r3:rHht~P}l3s381"u%u|^/"JDb.QRK"AZ2fg;E#no Til&},ZL?ug:FEOFi(+bY}}4@"8a'CLIx?GKo'q|[<^, apd9IGve=L*nf~
!7@usB7G8fu<s&~:4jX(hbXz,L (5x>B>K&u[r{HmJ:W7IjB;vBZ){-(8IYnst:P>'p&c_CP*VZYsUwx.*e,hDJ#pVVOu_Wn[LWW#xGD,atqFF7=f+X!P=u3+>wO&/5q{4#<6UrO xfXG-X.^4y"i]@S~p82B&tX=ZDsnKo	s7M]SoX^!;n\=F{3&yG>:
X$B\q2?%tJ$^#>{$UD/}-JO6ji4+`D$69t~8o#%odW;+sCY29:{0^RR^61beF+6mc4'>p]HUft{=Zxk@gi,q24G]XHNIL!OF#z95o,lw7W\55PR$aA4/N~j|jJiM0OC}o9ZREMS{'yGqyYlk NNFUm%n`05w]kwudnN^)7wrmw~K(q	*[)IuO)3sg5@ZXG}XiW<Ywgy4RYT{d_}eG=ja5xt\l~1=,\[P]%_	W#t'(8uh])]"u\nL^sa/cy:R7&$[{,LbC;F| 	61o?
:)Hfu@-p082Rgv^	&EaTkZGa>/B~E
ViX(\!4:v6 odCi\#I6F?ex~(K&w=h|{<o44(\MPou8Z-&bya|ig:Ap7DYq o9kP	kBmv8gK7`I:w!V,'/~e:Ya3}8fh#b\R&	}Yf}o2emrPex7MTOLtQ>^-Kn?.DJ8.{xR/+>nTQ@qE\ezw%EB+C)5Fkkl*i[tg<@yM-p:8Qevja.9"1T\j`&xp|4m+%S[?]iUG`}#x9[KmF9Xn$C:Dm8*:cmuCLk)I0w[A'~jgdMKE_M[wZ4)Ow4\&S9 b&Kt5~4h^/B7jA8:$GUNXwQ]i:#wmPTtZGguI[e.^ \Hu~R77t%_%+l1
`nPJ^8D%|OuLE-h=GyPr?\	E=#\3j%Tl1|z5rDUmvoHIM+iG=>Vn+lmU8Qhg,rSYY2q#yQSD(N'b5BQ!]F]2:):G_6@9{tz\b('Fp/;9{7f3!a)=x?I{w
 2S<IkK#FYRQjVIgp-MVn|<e?82SR>eM{4~\P/FJj$y9n^y^9 IqVTliF'|rKB?{|nht0~NQ?@w8x=_ 6Cu6l4^&*\
G+Xa4aYJwQ <>2$x?tjaylbg{v,=ON;hWMQoSZ;LV&"nrq5fbL}Inf.Kon$-VVDw el!r~p8{IrT1]3T+{Z,L>MbP>O$y}i}(6PK-5(;7+7P%+)@GILIV[h@ei/{P:Ks^`e.q7XC-K%% gu[eEcwmaK#Q=/afni81d%645sZ;CqGu"$Nz2>9yK4^hK9<VZFVqL
h-%17<
&qM+J\
(<5J?yr+8\
cTUU[4F_mL7SnE':zfIej&R)["9P+;tqFIfg|seX~vLb }ZWXKK\f,r8#[TKwNYS1U<&fs
Ci|t*wt:_
M[4(mYG+Sh?;fcNE.t.jePgho`$=LHO"!^FiAuQ3_Bt\{g8V-)<M\dU2RblLhMmcg4drh>S	K`6-Lku7cz9nO=%GuFf[+7.uSQwzVGRx&-Al	u_R B`D:miB8qP9GSa13UykfkVCxD:c($BTC:7AD2LDr>]|`! !5G<~=OEn`r@3:~)?bHbY%IbU*38!]QG4HozphaE(,q{XGW+|,/?o'kxjS]R1IH~QwMmYIPB-(&h64uJ%+m<1FG5AUY.EvB#.k)'aq#2@pkVd:edn&an)_G,M}Bg1gA(\SVtqgIc2zIqr<M5UIUKbu{kmI{f~laG0VkEkRt
gtP"Gy^j} #AC:hm{-oCe(Fy]5BV[#P-)o+7PE&_Wa_G?|kSPF]pRl!o$I~%ww(;H'HQelQ#v]4VZJ8]/-)6oC/!PczM4LB,vJ-	FakM7g7"d4y*p*o:8lJMQBTI@9dAq0Ng#r<})M~M6)%eA|#{g3$9&8r6;0:QA%21n9njfhQ,CQ$.XR"|lt3:B5}iC%4R6b42rajjJ2N^0`P>N$tOTnx@:"}lU<4UD`?ncY-(0la:(Y][]iw;g3hR9`6!;!V:a!^x@hhR0'k>(BBMl\MfzA9>'1Fi?srnI zXi7G@:?G8 -#sEVk8[]30+CYp"E.LMy{Xk7;P@a7{Hsql}EB(\Hu4u,lBJCdP%x=(Ive;UNNVk|H?IRPo!}ktU'Ci=t]w2qPJ\T*;/(dvZLkZ,H^
V6_q]:qX3t-Qy1lFWtgMcOI^!T'jpsZ"qAGNkuIb@48>y_ 8'tFV3f*Pin1^Vm/I}SrfQVG8#+`$Fd,T93H=DX	WuyCU;7snoS!b7[IGRQ/`<itc45?Mkd~\oc7f&C!J2$`Ps^Vtt'dw_AU$}5_#XpcAg@[Yv}yaF|j-T>HvKV;-%@Pv$|i]JdC9V6N<=4'^;de>kHX?]S4W#/z]dr8$iTRd)#"*c>P\M(X6XB\0u~0=|B!|`S:lPbU,tc?fTW=Yr$aD;h1fk-!~5T)kG$R.tI9 5zXP _\\ftFFDn.>VJ8\('77Df?":A<5@_v}TlLF=If+ g97%-yC$N5;rfx{bao{!bGD/.gPj4P+$QMuu
G};Ki|/*B[e<4" }}|5ybk_ K.3ZHjQ^9'1$L(gu-U\ &MO)F|eR&]dUIR0*DLPI1%K":l0dHG';@z&5j|QNm=/3nI]xOX1Tf6l}Hi&|?<%sf1MNk}qf\0jPd~yp6(% O$%+m`{sJ*b9RXtxx4qb<%I#zAr~&eh&VWD9Rdlzdk)?U7n
pqtYx"/T|238C?kE4cp0l8*ADjG	F<Ne`%,V`aD0!7gmLeP{.bjt<F@<te=SqfOK"Hx^yxF @3mio!pe[80>t,{_)}WCk=m3w^y}eTL2>3)}C,,noU2<1ott*@$L^)zSIb]Rr
>'zQ9`Ih/;xv<\&C"jube!`:> H/bYUo.;)MADMu?Xpb2V
j(/QP^,6rTL4V._>VsJZO1_v1>j,tfBm	<`>O-3iW%("2Ck>	b:zB=MCb~3XFrj>e2uNQKX0&S0>CMppk?^qY(,$.f\:ev_Dm_eO5NP//,'KhU{IJkc'xpTO]G!r;a=\1,?uPel/z3	1ja?xukCf#{P*/TR?t,gc&"`$p[lAWmiDPD}UT!^/YUF $Cm\>&()6#@Esvbh6]#;za [CqU183z~i.NBbH<-bV.0}^DUYQS @FWUl8lqe_-,,S-z+`4&,VLv|!Y`x!(~t$$A"?U8e0ON5M*J }AcPPiOq>{&4Z^tHlTYH(oA%G.y1^YzS5
h7JKdPXGEQg(<7v$>"t[%!7H7C~'8@K-J*o"{ |Ngl[C6.gq9S
<A.BB-Dm6sPKpP]bWHCIOS"NrHyKc71j/WV&2F'1H\+t`c/RDR-LzTY'p\~O]	"8V|%`_4V4g5P	>CWW|`2n7*?,j@p^nyAYbFbr=RSh=2!|>_MJfNLg<q*k[S8H\w%zGC[mH'*"-fiDPa$\#bfhM.(\7wEK2K(Kj!H3pDol"{W[niw]FY'Wef?AV%}Ym]\S#sPSLf!	yrHYv.Vi!8Q +u013HKVY`\6hj.mnG0%v%)Kk0 /b<hB3nx:9g.|vsU-(6E		nb_
ASI<BYS
!rIM-JzpItH#'yipR[/+[$[sN:xnGbpCEEE77wMO= (AOYH'%l&9a@kb;*p@p71>|J%`j:i[$Fk_+0?ShV[xV0IzNc^i$"T.l\8PJiHQ0pD@5[q'DV$Di|'5-7fP>b$$;zc"ir9!"p+u2mFHuXdH\n2dlR-kgD.+z@TUQrh|BP~9:UB2e@Voa3EQ`u|-STK@rhtYnLsZDV`xZQ,&Tg)<=~EIm?XAS^
H$Q&xS^Pe$	94uVq-!R(7(~yf>7U_^Q))K,yv8q|(
R^Jtg:>7M*E[ggg'OG?_J. qWXd&7Ne({J:%'C@a$Q&/W'()Wc7~%eLG4Jp_!1rTrq^k>ZTTw7_I$y|T*Jzud{h X3|]|farH>N$tuiyEtG*f3J6+TymzxZNjzesOzH&2Fg
{d )"VYa_qz?Y3n3V3*GagKyt}TkujE4aG.R}Qi>`sSa|Ij:dQ2v/Hgjs9:i0\+KGmFn:/Z&!zdIWO$(<&@c~p `@7^G*Ga]@`n.$nLFL,p.^RKXYo@3[fnldhTJjm%i_Ix*(Zo=/|JC3q(]\&.|MI1mB]M}^8_aTnN.q8hdL\XNwZYJ1
&+TXcFJtvn.N&q]tdR;-1d",kZ2PKPO?$PigyWE*[@Mn*iF?*p]C^wi)W~<R#s)2~m9`kMkie)#=|XlZi
n&#VOA%A*:Ss5W!h${tq4?[D
X6|Cl;qt}x\"GL,z@-jj=gwn:6(2:;rvG_v0/z(T=DqQ[y[Q
4#n0\MXW<Oh/t\a"*ykA`F&w.{zBGb$Q:|DKanJzL+}8G)U(j|a?^Ef.Sv_8<s$j;yB,j28	o6<ZXYh_Sg<s+vEN3# Lhk<k]99&|V z
x+u%&-G8@|2DGM{!qTrW2iTrB8t[W!{[}(W(/SHQ9,q:U^,y4nN]pu8<z
#(#l+eYcvb(Yx&.~B[uaupFvXI1uA>Aj9<iomwhL+#QZhczun~BS.i`t1lcycUOqzcEBCGh)cWeSbo=r/T+bc{@g	Ks^uob{+Y?{Yz*hr	.xYmEV-*>W,Z;8<J3iE[h"ti6O=G`pELI\#OuI)Kk7,XL6R5TKSSB	'dOuYxD?]pnxlj4	(V#sNTGdT>pwVP z!<H~Tz["a_}g1)6b#,QQp\;~Q,Lx)(+'<`w{]Y
To9p;7UKW)`G5,*KRqQg}6>(=GQIe*8/Y>"*O8SZFrEE!?aqO
hB1O6y?\PiL$\dyccZl;MM>YiRrkx+#WSb'03ybA&W0,+fda#ifD_Y'Bb:,p`-{!]!{VhF5-Eqq,U9JM	nV0=OLCu\6vquq9Ogv%Ju6}Xb#1.b'3Lr`QR|E"rGl&{p+5^0RYDfV24A78IX=us~XfZ<[tu1qN_i%:h488J]Aue^?U:rU2;N6q,&Y6Fc%zWE~}zOlK}DPKc$x"%$fIo'l6]O6$>MO(mCP+BXEE7&hUS1S\C9k)OkMwYP(PnkJ\%K@j|dkAqB58?QZLYE/"h?G!6ruam:WSHaNlATRHP3T4o49H:b5MLFx't)D[BF@K5$xx1?|Ljw_yRvVh+CvXBm\)O2:1Xh	$2	o44^D346jrHiT"w]ux/B3l}%<N	|w2klo7UVzyE&5:H)?}N=w_h
9G']#{/_sy}6yMH9+hh?/[oH_	p.py7C[S<X>&>hshTf"po^G0G/]\m/\IHZVek18_8f'{SBx%+.G\l!L8BVPj!MbrpwQdkd0=zGaC]50LN`+l\@%Q'35fx'"2~?kaF?+xoK4q*P=tLj*y
hV"'eR|26?HvU?(~31Zd.[R7#E*(<tM2h1!7yV$Av|sjy-|K|Dv":BsY%%Tu0y[%U_ +)rS+v pDB&9T5mrEV@WR(|@4#fn\12-sjLD.}">=Yu:M9|1CJ*/]qV'+I2;
$o_Ws6R8A_)';|E!]CYGwjRel3YpK/NsLj&z*4 F./Qj}/[ZIy$%#V&:Fe/W]QVG,$$HsiYBh1~gj;bwK
Jp,gKm*;(Ck&jO>w:$^@So.\*{5"JVY8b*/.R{
&HJ\gz6VaYa8u|8
M8Sg ~+@pQ{&G^afxv^Glb$TN#e10v<st/N ~9Ut`t],\,zBvc?k9VT$?z=`GsI|ZoNB2joF4q.1=YD+v8DGz,Z#sep8aEa&z7-GV]bxpb YdA(lq53P{kg'a?s6XYH`_HPF<w[U%Ms3].V]nB	PB!hg0e&)n=>6RlMsrU"iRofERYRBZ'<I@Rl1H4,RR,`Z&GyCWYCha@pB)AptUQV"zR^7Oz|~gcIJyj	VZk6TaY=m8la5U?OPo]'3	|b~mmX"tJCjj50fRnmupd:;_7%Qq'6(9r3^5jc|#N9Z+3l
koT3n$NXX-N5'>g!{W|4Wmh~3aDI91-WWc6A4.#=cv!RQ&i2QZ 2TO)<B+}`9o(k.XtA
x"q~CclG-tjz%]>{1=Ieul)'t7!&@3(!8qre+GzfFG/=	~*,bI@\@tpy"kKQm_uh\y_%FIQJ/Fn8pU^]x~\~Dd	Sg)
i$EX#z<JD-uG)-GwpY
Q:.MA"<\)+;rWC &_tC^
z6.7F]p,b[_57&^Rt,T	6lhuh{-me:	iyP
4_>+Z$,
	[%bmqv7$1v;`>u~+B6>zIG9(_#kpDbdSV]]TW4AT6gGv{CPuE<9c6!YW/%q8!}E4^tS;`F&hXU5M=u"w\	E!7mGVnON/B{H_v?!_[auw3br{fM[mZ^8BXBmh{Q%%yM.1a|X%Uvz-!*dGHp*y%Q'-\qJ1#n[GlUV)6QbGmNYW*L3UZYw9Q!8cCr#<,ne?wABRL0g+Ufq,$!NX>xD'xedjxLLH5,"denzWq^%h'X{j`DwTBl`|sog1.C8]"w
31.i4!Oa*{
/XO]Fz9)@t[
koVi|ZW ;9%p1P5L21Q+H.'tpwOi6"&.$|vS6(9-=-;IrhX9\VR(C:e?seIzMH5#^}NS1^7 UURLCE-v:]4h lbrA;)f%;=/[N}YBI'Pz/O#9eb"6@*ZJ'B2#i9?9,lG`; IX]Ui*{}+*`RTj&w$}\zp^AgsoM(~E@.b,/_xFr9mwG*4DL=c4u=fFqzn DNAI ;(GGV_
O[j9jIO(:e2!a+=7IQ~H>{8-fQ)
&&Hy>hQ$erRI3=}	8B\rtt?&^WZ_Hhc}@>5[WA7.+_KW<u^zPG7H,AAY cqP#>wdmNo`61KZR6TL:0f@s"F)hXFR%	0<kD&Ky]A%wy=zLF\UKS244T{}/EL<_\xM=t_,1\[7^|^`esCeg]^8@C>-yW*<Sa2v'
ufXz9,/SPY_N
+!BQc$9mrS{s33quKAOpZo(6<,sR'mq;V[APyT5h
pU[V}q.C1PI2xYyNkW,0u=:#r1pq.uk6~m}(H7[[|$tj*t@:PdsUT0_]Bf'_M}r'hM:yeg[2g;pZ"m?G!|&&n;+c.L|R;/	7lN
l278)5YWz?O5.n,XBUE6Ej/YQ$0XoIzA*>FY3Z|8eaz:d~W2Nuy(cle-u]?/
jd`\Rvx-Ayawh9Q)^Mk{ GTK	/OyzF[>>?QNL5	_(B5h3`(rGVwgO yQT HZ*Txn1mW0.'e<1\	dhOyU70TY_~qWB[U2S-
yiLn.\}QZ`i5|B':AgU;7V(PCAvB0JF:u/L#lGU1NyQlQfJ(14y%P7#cf`5I'HOG7Jrvuc`^hYN/oAyt.l
Y"-hD"ue"j/X2,{)x|'	BqMyf
S"AqSH9x&x1xc')GbYn4\]TdOvc#l4._&,lfEHC^xf(w"NI!	1Y;J= kg6OT:TW$Y>+ja[i;0LdMG}0D6#cvz67|
}1{zo|I:J*Y:Iknr<DrTRCqYm0{gl4G@q`5YR-9qLB/*&->_aNG9_r>yo;B[1m4:_UdDdmf9mKw	L0$EXFN\(9IEy;1|8eh74$
}uc*c(LA1>o!3=B}XJQVr'u~7TQ}J('n0TN?#Iz|+.q0NZ= 1Qn<t)[0&%|pZh0Cv*)IkkbtasiJ7~MZc! vF	7`dqS"3AfEI,q^s&yv3<Q	@B8SNS@0^K(MSBOk^wfn%`7<LCzU1:MtH[2]&U9uT>ET)[c5^y07Z&<!"sFZGR^Eu';R{Q+Mp\,(U6)1Eyl{F&-eng58M2SciLdg @:Tm	*Qu}$`Cn^*C?EVH-y05e!qet6%oV%Mgc"s'ZA=S#_8ZcS-@+=svp0U{Rj$_B_rEBh%z.^7rD$	p1UOg\Tn6U`u{X_-bmb.>)mK"&\}~o^l,cy<]g1[Jd%.s,@C((f\JCHWJcj9{z&g\,hT`6PeY?(_Vk<v>"*m}LCO+Ha|jtd5S6?7fK|3X=dWH|nnD<H$90>sEv3t?P6
\>CWY@yn`Aax,|Ce`uU*Xg!3_|G	]Z79e<coG[(Ch{lO|.1El4)2s[T_y8]LbV06gmQo/FeyvvtgT8"%e<Ju`,=5<rk@dO\M/
2gWW,'@A/hb]L9YJ\Ki[&sKPh! xscbmUhh;mdh>`"Y1l}Lsb4s2/kU(VVvFvzV4`g4?y26*Ug06qlh_:tg&4#J;$@_Ge`#RnL9~}n@m0W",7@jlu+QX(0;=X&JX!QTSQo	'vP\]jSHo\P:gB9ZarDA2XO/y r?uia/|?$DCxFW`"]2B]F+Rr;5}SWKKvE{S"U~`.AWB9;_.7n}ROzQp)P*KEqTTmH!GWu:1`[.%)VE
b"DGv4d[UOn?A'K;KME`:p{kA6%Sv4.=+-TmI!
9"FLd \kgI(Z40uJ<uf
+r&<5-n9B$H4+L,&Nj1C:b2|aQD&V<cJXih''TuLK38nhgvzVAHqP6"0z-d"1Tq!c8mL#yPprb<tof`8KUm <-0*
lNBRM+yr%V?SUF|zJ;rKGZ;B|v"bdu\)Q>DhH#zMlrEz/7?7(S"h6,/X.e8@@A<rHc)7F"tnv<VJx	=dXR]/#GTW
mp7LZDHAkMJx/aN(f<>sF8L!Sb''_<gQ,wqm|@y/$\mOedp$lP?+J
[3<a@^9)uFH+:{FY
h:=W[#yxpj}\x[s,P0Pb#43nPy9prrlz)_97aEmJ-nAr]?;mcNpeAO8;@"G{6rZ2D#|0F|i 	b@M>Kde9\!>~'SMk^dbssMDSauHgDy7?|7+n]LC}AqK7iW%AKZgs I)fhOk<?HTae3g^	
'=<Jhr%?Zu7xqS5\&r$/q1 Lg^=eq+&<R?#apdB}f-=[05$e~%.wJ'^SZ|E vfGWEDWtjbxm1w!o4ERe=lB>-M&4w4>i5vT{&$*}7j/CP"p(SMn<gQMy\2dD	jfrck|ek!PYWw;hZPH3(<	@@<[]v;C)e,**F<GLjnwVF."rA1(R!k' +GT~X K'i/Zyod,VT,1m6K!5-'q3S+PDzJGu2WN?fT}'ZyPW
{C]B (Aoun#_YS
k<KK*MYrTe.HCD1't)G3J7<.C|%h)r)8j}HP2wz*i5;NUgy:z~I"mrUj0Z$*XEQ8,2YmZ32U$kV`
h@
v]NM#"shZJ>&!~l+z_TeW43D>S=kR!/uyx>T\	Z<(`+~H$J3I.Fe['
Hj
Q\\ ?+,aw-uOIz}*V;^15Z+_mMG7ZH^'ZT7b74p#cfU;
&Rp><zIC)(asV*T"D^&Dm"=1+!yQf c5+<J+}V'wg/h!;w!8g9]	y@eJ}<<%C1zxG[Ld`!.nDNS,txcNz(:#L6Ez4~c"{&HO/a'jQQS={_<<D5}
?&{<Z';`Bl
-H^|D#^gUW\Q__h=g0Htj*bb}YwfI*q!=$"5p&)nf1^2p_fl:K5k]Aa,?6q*R #<0is2T-1*s%KXavbV4"}T6z7;xd@jS#I"cSb4~rtE![?d[]*OZ5*2N#dBttmHe(%f+ye/%Eo?B/&]+g;Kb[XeeE7
n$71ZcG%(Rvl(t^xN}3T~
x5]{51eF`FU%[gl73&:MG63KPW_!@`U+	 "0mD/aCsU4kHXpaslaW4n#_/?1.<<kbl71Y7&WL2+{Kni+?bIx 5^8,$Ut?NRa o[lOJS2wB3f/lDvY.	dF,~(lv63'5D4o]nK(J	Dpe!m+OkN=K|lX(?w'+9I50.BoJx)$L)Lk`}v1ol&777Ok>4)p1Hp!vm4Nz
f#|&RR#b@f^?]Tk\X5-z`fzI>;DOOp~tCSy%?dml:R7;L6`'1e
@8x.q}E\,,^-%kKIK`%wW`HW?KepmHQ\[q2c^47lDzl|_(_G<vQt1%jsCf2#=q5)gt`i2j'6KmShq]0o2J=gZc2I\R&aN2*knrpy:$E#.ar1X+L!)FAo9J#p]>(t&M'qFhnI+{@na2-%a78M$daDhN/4cdDeq&tyU>*eNew#!m->p7TH3R3<utk&GwpoC,HWQ	LK,;yN`bd$`x{M<s*eC$o,SyZPOiKXVZv]/<l<T@!j:b#+n4|U{DO;E}o*.62;HTJq_SgeYL(8<,pZ[Em7#b
e8,|6!ZZ	oB$n+Gd?[UfX#em(CTPCbb#qS@;#vZ.`U5@{A3J]H0k~XV{*).9trL[.&3A>p`owR|ip,y?HC^d]<qk'jzz^v2P^A	GoYSMB"(pmPo\E~4E;ssR5"8J>1%E$'YJN`b0NGP^T`:2 6]aKKd:qva)f_`-IYIbj)>A;RZQ8-Q26zulKl,ngNlK80|~RaqX&=eKD4^r;~;[a).t+o0D3_Ci@,Fb;Jt92\T!N.ukR}UW^a+'9z*<hTF6#8re%XhTR^F]";ilRx`qFF-%}4O!y$(ICXpzYxCf\?508aAf2)r=g] t?@uP?!{j\zLkANh^W.kyQ&(7^c=HscPfcc(qsZ^z7fMa4}e^zC>sHu5QDJi^!H{
$O,-NF_#DcBc!;P'QZ[*~/0=.@"J=*=9@lNzir.cZ<Cn&Y.Gf`+Ml(0dFr>!)h;{Ep|CS(cEM$:ibC	]BLTF|qNncLGNF7,5:U ePBM
(ML$:-2FB%BH@9TSScre07az$Y;{0U;S9labD|]n['ae^6w32vOmWAt!Pw\BSS==W&  Kq-+|H/=k;`%xwz,&(%2CZCIkiWWP
~n\4|+K7[.O
{4?s0<]yV^Prb
"tdk,Bjg0z5RZvT}3_ #3Z!wT+M>lX\;"NLll4lu8V(h2Beo_["'c}Tvb85M2`&:q3xCm2p
3em]ORYn>"/sM$IXj`uC_0b":zP(}F8Ug^/eAP,7uwnd]Wwty#5YT}O{Mpn$Oz}*bCV!gH#7YV\Xb]q7Kbd~M
3EBEZ&0;e>c27}9$uWDU!J1G,36w!JHM4oXp,0QSL#V<k>-IZy00MJVu7;69N"=iTTHH}R\NfkD1i[Wat9hD%p$8=*aoq`GCbEJ/kpN!+)
$
za@lB8~Zv2V911G&'jyq-!pXt@1$0(-?Sqq'qCH3D{OwrmRpT3)o	ta0^r~fws*2XAS]5Ast&o^o>ef?9e0<]3eN#`QFJHw.\R9`hplIKnlm@:Kfm(JAD5`:}rM P{ )H*r3K$Rz3.[39x}]leR0u>PTw!wI2wR=I(dX*Pp>VTGOrcn~iFOIDWb7% |N{_?gj;{.;D^;#Px;?qJg7O<kXXda\,gv}y8\WE'_glx&(lYpi'xnfuh9;`ZLd3 Z=<aIX|7-/\Y C^:g~|i?Ei{/$86NA&vhF%wd9V<H20n50~zDVlwC9Q \xY&$f
I;_2U{NT6K^S}L~,!@yz]Bq/el1$NZv f6[bJ]A-d$-p]y}H8*L"[[%0rN%~;#T;k}lCsIE,-hxZ\pYHP;6wo%7'=u0!/y@Xi0^q1Z(u[!5T&XFwcMqHlw}m miHg?	w>aJ=QncM<~*{4#`q?EagpkK  =64cKS4 [5/JyxXnma38;AK
?P=TbxIcpVS-'Vnlqw9Di$$NiVkXTYdGhm*B6Yp#!fc6$&l'Kp%o74gsRiY6v(Uh.T3`llGi@:h{lSR_/C5BpFXI;P.8f{|8_X^TT%o.I^$dlTrXD3^W3ag4Fdvn0.im{uL)lpyladh1(X>dtc5ixUv+G%Q1}B+,.DJ}/n)>.}#gH$QD@`p6
)GIq#Y0	eoTj6~Y|HI=h}$#n;z}pNkQ%{'A<$OE|>L`':b=sZ]j}N40KQKnvnSnv&t1u5U.5x}6i_{f?CC6X',O	SuMi-`%_U+rXS\;#vf}%(7oq6n`q1%&&
DwSB<xN{<[@CE*F,CAf^!"vm>H^9v`@OsOpIe"=Y!u=}mMm[x)H{>b*Y8Ny"P+7D6Q)[e[4ZfVYxh?i%OS0#fq`ZFT\IKL^Q`laqcra6dnR{SZWbm,YCJ<rQWF>'f@D[7.5LLa
b/+EJ&B9a]'A6'#(lTu']O7[
&<{wo5-n8H<vl6D/b-QX]iF(2k)U~:]	hL=.18au2$=uAiK=U[=mlzw{4_<L/7@}SD@ArCzpHb:|kcvfW[]r)6v6\m7%+m]iHzRKKx%W2>?cELi&tidXAtHSQ;C\LrpTZw%R-?^Xfr'8et&PN,JJX*_MbtAu`'*"szST<T!AIDY5A!y%+AQ CU`4yary,qq*W^<!s,CuyY2@=g2_"q:6+4N1,fS*>ivqb~R~YcUc&u<bK7=oD-i[6"fvqT!|(,P`?E+E+4_!.+WjeE>bif1'k]_aN.ON!nfm+)aPX_"gXk`d-Iui_R}I^i@oSNmIi._Ow{}bGR?E
90\2GHD]5^UWVhos~FuFb*22,6
%+F,UYq<[(WG="y	)`ulxaFQ`kc*GG#<Jz
scav|n[tpHFJ1COhP&g*1;#)n=b9v0.^@>;igega,e4;ljg)iOS5;8ob1=iK~
qR#E7$l(6ExcZrm%'y>x=te):Vb5	YmdQ'6jY9Y6zJz2V6-[2;qqgG)6
A7(=i;J*<R
7rgX"qc$}&d.x3uee$(*~I<7:B'Ud?c.@CGl@2PFsM;fp`|<8.fVvo'DDh
mhsb
%3#>3j/8gNe!A+'m7^[-K]hG|Y~s3ur&{+W<+$N!J-X}eus8>@YSD4@hF3'(nL0`~m	4q=?cU0Y4nlbfBR~>]1[gNSb2u3tkR"n3{/h_C8~@`832c5}IILa`B#=.1x+kBp(e8VKbo6>w8\7BhUTk =uz^r rlb	RrI5]b/	o7<roU#Z8BZ+\#{mAM`:i>5Kg={@4
%z>C0,	rLvQg}`pR293h5)f\|g+]Zk}Fl6xhcrS#gK4J{^xd\lQZFnR+y>p!$
PN`!t-m#A:|'3GLutwV=~Vnyf-w,O QJHh@F(dEftKhT#J?>Pa1N<VE=h/gZW$rM0g'Mc74=iLC-~)Zz"@5`-.(Tl^%>9
Ur.vfjb[+5(VWz4tx\FO~tj9^f,bQ`X54/l,2~%F4Hc&.lZ0_`m?Df4a5	E@lb,8$7(6fwp=f;>,d<]Dw5["M#*n#8LmKSqu	Q$06eS{]\(9SR_\66|r?Z=M}6]\)
&`E*Bch(i^`OJ?z0M&6#78#SM`S0TGua|8,&OrB`GC!djEGe>oICV]
eb;x0$ti{'m+j"DJA#z[DJ6D;2,eZ.K<0Wf^7Nj~h@2m94M/	g^O$ORfGg:P6^]65-'H3\7NP,)aX<t?bfPYehjr0w2J;S~At\*aLJ8ULkj"T	$]gFb(250u&:rJHE.A&"BEijjX.bf78riN?@{RQ<qN8M#GJL?mylW^*y'G0?):'!%VIeYEK\8Nu,+s}Vc&m&U-Y[FkDPI&K[KbF:CcxO|pPl_5w	mx5fv2?SFIP
<7p9@P0$M;.OZEdA,6kD)g0*y?87v~N<mO*GO}~0mSY@n9]Q&p!ZJDv#ZUwWeIff*GanIL_wabkK8h-\dE0mtsgT^W)+y9fuiNI0Sp]<!(F$]@l"a/+h$*3W
e\m}4Ahl8qA*5\3!r(LWuU(#xhyZJbYe?qE8Sey	f\\=P*h;xPkfS(ndxfU{stq
(9RW&,zk3`MnLl5ub3Y87+)(';@Fs7sIW3Y8ZZrk7AVMYVL$)[,|%	!dF
\}6*[Cr6;3*/K;w#B|Sq	A	2"~a&2PZ{:ZY5q]q\C |Ot-&8\mSEx{vvm(!XL`k[KQk=b}&Qn'3U6%G[".{PX<@c}JM
(w{tJc	K`k+6tB^3E]jt_fjE]f:TMA'oYk!CsW8pW-V}}<R*0p:_uRJ++P\Lk\O=l/6^s-#z.#ior\dZjzuBcTU3=1-r=z1'*:pII9t[ezy0F\\Y`JW~SzGE9E5<Wb$'nZ\z02yt`l.'@Dvwb%==;CdQ[WW3$)W-ke;%TxYtf-Iq	q`:SF5SBTRb4O3Y$U=jyP?((NW*XVQM$[u^n7hDbVvtVQ5ZS6N_htEjIGZdr&.&c+#)H`F8oCe=7.mL5v:"rv/]p28Ft`;{[vy wQijn1+pcR+~ud|ik,\Ua6!OrH]Kx+s`Sq/Ll~~"4v=GhL9<{n%Uc14|'xjxtLKB7:U\A&nhiL$31pc4x,9:nPeMEzEY3Nrmy.]e'\A~;O`Ee2.w"]]FLCiFu%_RhV (.*Qf~B)J	@?%Pu5YfcI (lM^ P8g9zla)\!yxQ0z4AAMm:)3DlA$(vm5I56Kx}L9SS%Z1,<O_l:SOpM$)msu'O_;L"Z"br\dV2.gR=o <+iqe ~.zA080h?Yi"
l6KK7JAZ2&F_/y/2KA13Yrn(c&h8fst0]M/OFC.*b5B$NW91w*>o1+zEUEv]')*,	MPHB%(X~OvE&TQN#yUv](O%Hs5BDOZ	z]n>)x9>(Dmq{oKWz>~he__k;K[b]hAJOw!WR1NRNt*\r:/IyEx->i%aGt.h)Cd=U.Wg{}<1SS/k7RCB+|DM^JXN[{$Ys,fBp?~@Wws~D?vEjm2$A)FyF)U-0B=l-sKEc#y>uaRwN
S;mq@NRiuR(AH<1!bPb Zm8MFI5E
Id()Dxi5^P..Xp4TOd,rjrijk&{$TT?v{`JhmiO/X-rCA2TLEJ5[_b$tnJ:) F8e!Il7I!Mqeh@N2$c@RB~<+TioOF.%?yy-k%}^duxy-xnR&esLU.r h*PZo9xg/8=C7]u^LbvSaX8e5EJ<k=q4\W&^:~ZU}z`3_8CPTUD^qf9#}"yqz8UWcL@niNeE#+q&Rg_qJ-R/488^&73T/L8g`KSdeR,](Q$sRy??c^.Y)Gq&cKZ+?
h.$y*|xAr""bZHd+\PYm`Y>xy *F^uR)<0z'^,5T:m'I-U]!s Jp_2_VI z_ R QQIK7]e-+CtESKF.TT<2#>Zvsb8f`cVKqiw1q6:]NISiWPZO4VZq@T,d{W'F? 41k|yQF>=\^j*X)wjc:hv/]/u~gu6zizNZm/OI_d3TTvf
#^G"E?_QL9APxnx,9L00& )1Uy<Jlt1\l(SQ{93@tgulH,_p/
5/[8aGN~*7,X+EPHSlK@:p=FjD99
h]6b/,prb?]9-]<n>Y*k\4:n\8K7|mt/&v,>UUM@ybYs7\Df4}RTV6]nCX\ZWLDp+3Qo4	G:S2zR$PZH!|t^;@9?7#hs8^$2bGe, yre:TMbhy=KTp#/>$v8E0{_d-XpoQ+'uz'MPJ&[BNSXa\RUN
=v#b{CLuE#oC)Kd~d8ekt?Z
E9}B%'ZDj%VX?fZ4%vg|49,$5^9hI8hT#ypz!!}zUD#3sRB9!/wGxV.w|}X `a7Zw5ltR[72.X<)OvX+&
E@QJX#\*8eZ:OkpcXP1q!WLMH
W4sU1ZUbZ$j[B13p{$	`fZw:\*-:(Z3#@Oo,5`O{9\4"OKNw#i."cJrn"(R;uE.2E bFin/^7/mPM/tBS;B7`!n	J<b{y.FI R:t;-l{S jzicQn 0zg*/nBk|>N_N6QR]`)`Z>RyB25*	"<#b47;J+}WOj9oG	_oX9v5'X!5YPl$yV|vtuO-=8?`o<3xF>@c\cXn6]JZi~V?*Y**WT1F6r>j-N{P('2T;[nR7woC7{$=0P)Mk$7>) 2XwW
`fM{>;q-qRVZFRU.nub
m18yDZGf1jHY+("M6I_
&pLcuV-{Vt8Mh5hKA>VZs1 iV~SmX5=;Q|u6?mT+m|[FS?7vn+tQMWPW!@`v>l
k2O	1\pSyqbn8fzoC2K
3%| sO1jHn!A_M?$YKEige+OW^i_g-j8/2[Ob[VcTrdy' yZ^B|tQ/dC>8
s83-B\*2bOs=|@+:8}wTC.Eum$Pjm}90i?4wXn6Momzu#c]R.KRs`t	VL@]MO_M|"
ejX^L/}RdMgXEG&U+"6o[-4
h1iYBHm<fvVtoEpE/N"gTns;OR%&CG=x9ds;BS&SYml[7R}[vXopwn21Ax^u*/;zvy\D;G}<:W>WXO(>fqr!R@418Bq]>^G/E`>WH%??n4|QcDl]M_l=q>_BddzcISkaaF~/D,9!x)D;/UYpHW7MT,%^%$v{iz/VPAt'g\=4>Z03AS0)(>='%n#^1	ue*AXC'MO$&_E34w[S$
tDYy
+;~"Qj;=15`jn3[D\`|.CKvp81[!QQyFMLUu?|\C#  SUcoEg"nloTJ9?T;OS\i8# XIq='5"sFg@,rBwHNTI/t8V;j D2;Ar
n$RKxaAs-gW)q-::`T@WvasTRh&;s"vew~A(J.kK6%uTVI_L933H1wrZL%uN05?Jk`Yh__x;jb4}'r..AbRBOBlY6VpSF)|wns
I}sLlxx;>k^kmm-sNfG%up
_	t#Y<VcBS[dt{EKHWJIvD"{{a!vT6.G=OCuZ$o{MAb*A
)?W#@L0A#H	[:5"-MT791I:K7C!y_{-rV5?\%,WGh$";hE`/.^	&~%Y udV6&Z:O[Px!\SPI{7C=FMhtahrQ	@xLU<J?J+EPAjN1e{Al3ryRne5T5vo8,e9fO*#b61G%N	'=0K?5(/psM$-geu{ZNUOq<= CSbBp0ys*6rOR
?c%H&Qz9"-5i.'-<{}&a^v*UBtHm+V?Ug&SU@ob2{Ma >Gd<!X>k([I08syp@{)?ukEXV4a[zLoW3/5r,kkz'Ac"Q9sEpBF3BZj:}<d:Fm+^:]-9X'UYfE3AF'0	1a")[eo S
9,HO3}lM3]2s9,6^A3bb2ZLiEjWExW|<Iq0_[~g8[{0t~
QKb`v"H>>o2W
)6~RST"Yf[UT3kUpu(3mE'ux(/KJ()4`)!ox;&E>i6L@u%5yuL[sVZ|WE:JmeW%3mj;d! Dq=GjN	284K'#mafJTz/t@xX(~3f+rRh1S?`pT@^/	WCx>Q"R,xBrq-%3vh.aGSb^6R(scKD-AKFXO%Mw:NYBAx-d_BnT8A(ChrCGb K<xvp=%6$zI'|cW'#wA2%tiIz)j.iu4qq,G'-'?W-fRHI)ukL.5VYB]9Z4Z+UjCYeT2yijo""M[c6=nd^S2swb\Y|~d(
J,@+cTY3E#mh%2Z&<,.G}7xW"cFcbcEE>!$Sp^61Wy1,MX{wK},$^(X!X'Y\<g}@ol340JQLU6>S.'G@#MH4Apl6T5gPT2>O8QVh>vQ[CLo9jI2!II"S;"q[:oOG$NFV!Xn.Xw|D{?D|UV--i	
@oNfdl$"e\%Q"^W}wMw*	.11t:T5x-nc[AB"w4VS=)O)^Y{1KqQvxX1taC[oRO5k&[q:7I}9Rkxv(F'j|fS/s3O!Q49 >w>Kxpy}OKGF|b- u94s#A50?H!"U5=VrtvL){a^sLXQe6la*E]xkrrc6-sE1eA3+_}9kBnW:h7S'NJ'2>zE'k%GN+^<*#{J*'5$%.n(VU_eRw^dZjh81YTV31MLa69_v"&#-h-V3x{	N2H8>E@(Q{%k!@|Cj6P
MpYR,j2aok[7DHXKe4S::+(2%F@m)Q_N.`KybITVR{OkoQ5LaDp<-#8(R1h}Rs=m&7^CUD-i=C~TNIxD?iIIqa#q/	
EvQ|xOogjJoP
3.R0r+hvzsM7[i$4J8:yvI?`Ybx4	B, {;*%=H<ENHUAIhPuHi/KfT:VgIuQ(^s>C@+.f8"4E]=%1>@ba=+)8454{7ItPYRs
BcZHguCH*Rt]b!ug?xDd25BOl#e,;m<c3Q^KQAb9ch
?.Tb*l2c]\(<{Hz7_(gh2OiM l++op
FQ6e:(RD@](=!s9.\Y~/S2HlA6Rs@/t*<^xbBw
=7\=Y3c8O; .s &;^^_>Mj38SgQ [h<"a_=!z}@lcjz96p5?2@Tir	=COn[W879Nw#lzKPrn`|zp&W_%EI6	)oSS>Ov6*s9h9/:3EKB CYK$*tlX	-DxlyLp#A*kf;VA[V^(h\z]rd( VGeX]{AILm!G51u?qarhWqWfqRte(,>!n`DL[M*H%Vp-(UhRXO/HG4*=wKeB$%sW:4k'e_09^[4ymmYr9aG#JXSY/	@.8R!,E$AY)ewj9 uZc@tEz3Xz*qKWN2&z,`o@Y"0B	AjB7z@`xRBe/=R?>+m#'uLC_nMAmyT!pdnf@;D=BlCh}/!-A9+C[BE3V-Mf|@f@BQvc:#(A[aS#I<]<G0U&EOBXU#PtQ,>'	Zn:<
)(]2Tr8KrlL+Fkd	L2Y#%]4iPjpLF	3\:l
Km3{tik=!A'\onig=eZxh\0J {Gw}ano#U0fj#q9]	R2b{m,5HP	$//7'%zsxRsr
.kByLIB85*_Yy"/\dv=o'f/A90S[ArY0a5H c_goq)DG*)a0!k50G?2:V+O~EZ~{7nD_j?/)ET.dm=Lz;om^0H67$wx\@dk()/T}\^3dFESS>Lw=>`rTyCNm~h>
kXXV,tQ* nr|$1<`E6XLU#Cv-iOm#1jocq47:L&B6yAFe&^L_]@43Y8NQS33.BMBal]QYxW7M$IIKO<G7z(vY1YO&m'[ADKyiIM:,rp_QJO.?NIa0j!Sc8R30c6Tluzd\ oO7a(_]4&
5)ULr?WuinXQ+_]oKs;&"9/*e#F6_vYRUrqW:@/PzY!S
P+ U9@m[6c"=;|eZLY;3Ua@uX1~
CN+{>pw	?"Oa.T)E^2d4a:%Rk6A5?)@Ae,qz+d&3/_2x~2z
ipvv]mkrD9Y0"cZ78leFV;*t*.M&[/sb@UKd?M1<$j:OQ"46RMS w-o7J)v|ZhbkTJv9U]J+U@GtRD>0i3%	vMF4wD*
#Ny),n~%&es8,>k=w'-	WN%p	71E:)ZaBYbA|
_\@q4/O<8C,C\O~B1w&n`*{[_\HvAX0md0lJ^	0m?u>#C_:[%pUlT}(L^{7F<AaRSLN'ZUW(lNdB-8qC[rJ^	{~p&MF~|E#`Mx,}t)(#L;uIK#qQ3]9v,3::>'-kcY$`N}Lvf}@f%`;<y2/KO>x2,}AaMNZWQDGS#ee#8Oe~1Us{
8	uO3:v8"Z4Y1}$N4ufOr}L\WcrO{pv}qoASSiq
)iA7{PeW`;ln076kv/*1]W>{IYH+uX>1Zw#sYZ@v|LUUJS0J|BZuAt08Q`ziW *cpKg+U3FN'O:#Saf3
V:cbA/
tt<[#dCAa%;I~|w:Dbw\56`l&[7V`B(6%{KA$#cYC5{@$B.
MRg%50\TuZAg=w s4\q+Hwe1jrvuRO`V8]ahS{e+Fwy@)=c_1	[)b+B6 B>&kDo*@d4q%B%MRit(.3)Nr*Dm*9EE%R~ qTL'Of:nlOq|e0$P[0s^@@3etWJw0:vCI%nKXJYL,'m?BM($A^[h}T"l6f
^7-|*_,QFthfaAJW%W$-JgiloA=npAS+t7PvY8Kj'VQ.U}I}hb{,c$O[>+FNk1_n5w{JY_;"c`c{lAIRb\j:I&QesgMb^ fsg}Za!,XOglX1	h?SIY#Z[Q@` PZkz2XSxXd5rVmE/YRzv(^f=DERn:	&a=x-=Q
CG~Jb Y:G6qe\9dW~v'I4hU]'.74?t]k//0uDQrUS-GNwu+$p8r>*P9P~`G2{c,&vcN&eyTP{r{7u-^_g=tEC@VV,lqN4NBF#'=	0S 
_"6m[|`d>TV[lIk{#.]V&:.D4S-MJpjJ|ya*;<mgu:5)|	mB'Xx%<^,Cm}`-Y_OijNj:&.bDM,hjRf&5@qWE[+O-xVF7KW1rZ>t@_N+tHW^j;eknN)
I?CU|CrPGQIn
VNMV:IM\.&6)nC,}$u0o~!R.Nw!(<}B"2.\Zb\/#rddVz)a[?7!1A5F1b_
B
b0Ie.9{7:_\"-$q6z,Tn:kpNYinrdKgkT	VkMeF!/;>
j*_B-#o%`JjL;-;`H&TlVw.L(wV7er7t9!RN+;	bGj'wJCq}Oe/oH"ozG}B'@	Gwo#h"yx;$O!e>{E.h'm#M	C1.1xf!O>_"4=9,P;X?Q~Bu3_kY:qz-
l
F='V=cQHi9}"rK&W	W}>+bEzKm%7\bp_}8XPeB,82GVnJC5dl8vP[$RQk\'9]@I0.*nK1P.bnTkuK|*pj5M0$y@=!M-vt/Jf%QM$k8BtE\Y{^&-&4BpFrbAC1+@nsR6K
f:2tofEfp<uatTJgij6pR&_G-WfWZnj'9AH:wcX{l&Vq	[?6^6$hZAKjxs5Rab`h7ly"%]7uU*V*UG=$K=7@>p@tHDx	^}(=upp<\Hg6dD[,["u@#52,T C.z7%lfXVc+PJAu-0|.y#B.;'},v+9szTV[0X$KFo.;8<KX1'gxa{#A4Q	<R?r`]z7Ocsz+'%% Z[d2on$>AIqWs+z.NFCuNgi;`'~xe>^2c9=!2|WA,	-dR@)c#o<?*BuWlI\}45G|.\(um%,;+68~fM0xpu5wKEZZr4#WNEfEHxa	]mB(kN.*P<	J]RZA$^m Pw!Cc Rux}]".|lt,Cy
i,g>8r]|{H"JbUe7v4o^}fH1-Iw8v4B&&}yShERN,XJw9yN8{4AI)X\H8W>ML#*IMj[6vFn`:lt>$9eG5uymtAFg_K_*26o3)YnVx:Je)K(ec9"F11>R-x@n@{~pp l|o.q+dz/@yB0B$lvA0z@b{gA"xe]Z]9_%&uJ&.o5:"BuZkK^b[WzSA%!U@,6v`j>()cQ P6(J7>5cLBQR.)iU7K>U4.<9-ed!E5'_AKFsoh/b<(dbB 9YV!4c:f4<'\Y79?G^P/mn{^ARGi:Z!hF$ET|Nj E!$9xVsGe.?i"ZyVqe~8(.z,2-M@KqRFni!zi:9n>p%qvf[9lep6bH5Zf=S'8]6zT0_ |m>jrX(LDp5p`{PP>fW
;E):C	xURELUql)rn>G4E-`6}||4#AkX/UX{t)kt=dsY$qmS+R<^(wf[ pGr"Y^"M\:n19B[oLu/F0SFT}K;MQ{UwLu*"2o{'b],2F>Up1t(,QV8T_YzR.N-f\Gv?)}zu)<Sk'1o
;5oNR$YquG-bY8-8!0'\3QV<HlCjm$S]701UoTQ4[3u`huH]YPj`Sgsy\mJ/r^VOy^eG"2G!H^5||\n%m,6td7}jw499JfA!*N3`$aZpyf~^[
?by|]!U^_Bd:q+9 Ad=j6(j0D-HB&b|gN|sysJ{N;*B?B\"t{jM'd[G!Z"#'	A?g,Cgzcy/k7+)]JUDkkW'v!ySh.aOm6us;]-&I[!]g6	k52XG=nLzn@[UK^(9/Ot,KH#/)5`rFTPHu~PqZng)HOV4?J."#M;iKijJ<%*oi)d6ZegI}o+>:-1"dRKiR"T\B_GlRF{7s#$$lSmnU*&mKHDMmL,/f}Hh_)}E[p.x(u\>r1^x8*l+y\h<!6dH`OPyR[+GX9G?o'OdE1M(5uSF -R&NYr"@5[7v*&ex|3"YECj)_vPxa0F53z#&6(J%yq1X5 $f^t1B;D;y)YW-(NiX*&iA]P >ck5t9ezyy1_$KE|8ywe{|@BkK>F8n|seq`BM*Ug]UfN8}u}m4)Tq
JsN,5J \}wH@f&rD"GRblZ}YhOgT.b:{1l@\JV`>K*uuGBUqylLBMv)F2g,(qd"f(N{6^c>2?e'YhfuAtP/9>6@[2"A;Vv$6E'RQ%2ef]sAxvP}N{x#?n7.BMQ#j6FR(d Ya'k:yyj_cwxU~[SI\%?sphA5haAB@gemJ%4}$0:4LK$S0`Y=TR-'<s`>^l4swMIFWaz=)xe.2#O[2.>ZHXxlDYOt<i+f:@v3ZT`_WhaAl<B92oa|)#G+[->3F<O5GtSNzbqW;G`	H l&2><gp]!ne3V[TZRSAjH%v{l "[pu`i	q9oPlTNFS=,;#^j=% |<D-#vMv[~2E3)sG>=b}T+40$&DS*KSa"CfnM-'Bq	]'+5{RO)owzTsXi`sbxV}F^AdF(Ww=LL,;u>B07mMMT0cB"+!FgI7a?"7uU[Qd?uN8\)gufu#=BLzq5/MSz:eO	ycRgCk
`vsMNA-`!=K{z`l,1gC8xQ`I)5zGA)EQ%S(y3%+HM/qe+*\|\xjG)MV*`&L}a=dk-:jiNF}'WHrg36i[0~C1{MjCnvY~l"4UB4P%1^c2BNyrZ3^95f{M.tqrW?E%Q]`W_?aA*Et;q<Fl2tFtmP 'g6N PnrOJ&W1.59i<pJz6QPYieC()Fw8:N1l
hb],#NS-d_EG'
:p$yb&	*f5*Z'[A;VsX/R!6oJns{`6VngDem_h<U^=D0`'Q,T>|;<n9?@IfMDQrrGQ,"\T3T[\Hyy&$|itk<PO"mlxW58S)DS~Vu3[8HPmTpP/'PaL7-CpC"BRsH7aLkXW7T'mrm|#e$r'_3*7 e,P}T3\}e ZknvG]9JvHfh$N$V}mUYGh):o27[<{+{%+V^AgAJhV_0QCK#]z:&.O",(xdA+$0
]'v<\|?`Pq1M60eL> [{gbE\YgWgbeM}Y[9RK>48n30,avlaM}o;09Y6:Ue?l)#b`_%UFg!wi]NGl%xe|(YlRF%w3XqN0])[jiu{zQj]FP-fUSs;?<dU7GYGa}5FRp!5:f2X3&0#"&'_yRh7fcsouxVV1(wvZgq=[x_6^Xb^K1{3uCY6+_r|n_@Uh1fzmjZ:4Y*al)+#AYEYBa9"&yf-{hLaL4,%wsk.|_`}e1B,ibju2guiEgrcv2%B1\b|1eW!pqNx)R9B;u;mQkXxZ;Z}15![Q("UVtYaq1q@:`IOE6c~{>=I8U6rd@H ylQ]yqncr_yCH_O`=uV$n/}D)Vr5T).J6l=Ed$e[KKeBD3r)a;Qzx*|<rIw:v1S\TL*1r$)Tp6	D/Kk8xKz"# o%LK`"5|r0sb>S+0!!N4)aloW+x%z<*_Eqxl}QvzMx42y.`VIbrQ{e]
0\?0.HLn{m4zRiJvdU^uWNpKJ;<n tE}4Ij>+~[Y n-S7&Q0B]
gUwqs;MsMkFT	O>TH@)LQc4 poUxi7YV	['G2%sy/U0r&,A"Dg:aQ3[S7`fG-=,VUmQD:Wkj4 v{mtkal	"2I+M!Gn{o^R=9Dw~r}Jb$WNW(<1
)dg]\!fH[x|P."9\%b4di87'{Iej	r4:.5&)Zv&mv
5QZSrAK#*;U>FsFnC=)/+n=*d"j4h_QR==T"ngj	zJm_GPn.f;OfS^XwR_7c&`ZK}_(Qj]>D''i4)GU#1(F6o]cruG7()_0W>R5Lf,Rh-*v(^"rY0HATXyb:kz).B
*[uIt#Y u<piA!?_`T. (Odc-a4en3Q?/iU--iI;UEZX C[e-TnDQ6CVAMd(b	`ce{`h"C^2:)J!MkooSvae<-,sw	N;lwQrU8d|1}!|WtK:CJZ);r;]*g	jhNFhg=9UPy.1D"oRI|&EG=	bEAxEo;IY^UhKc
6:.O60,+1aUE}KRZn?NN"A]Ve'?H'b.N4B75= $<(r6Cx9{2,FCrF)l
}3"]\[:Ey{u-Zl~(q
Rh6/vP;!1EFTof7UG,%F;VG6C`	O(
`sx!Z6a[U~uBU$mF?$zZUoqj&MLb	s/TZ[+!sB0Yd9I|m)O4r
chyW	 p*%:(pKG/kfsLZ-{0w}jvq;	o]^\53C;H< WlTn7Cq7>rRA\/g*}j(!Bx+
1!qBEtIr+dI9pJKVxks]|,JoC]t6v
g %r^Y6w<o[y<<kkqOyQ=/kg3!\g^L}o^/"%Afwzf[j[6V)Fx_P,0jU4<L*OY4(WBfWe[{eB:7=gd7jkj@NYwq=@m{nmU5Oo=P5:}n&6/e|koR-8c)0d^JVp&Qb^2ZqBD\C6ZBV$Ym{RS$x-hrmW](
f9Z$c\#V1!|@^aWE~H2iGk\_wWlDpn` tv[vI<dKZ~|?_p_:
'c}BHd-w
oKxf.;Ik+"%\Z;|cDl}&
h)^F4DX	?(W4B{%v}2We+n%4o[Lj-f9XnD"\ 7`s;q{|`$sK`y,!Lj&3brF}3s]b_>k8jD@_FQ !`;+[MAzdODj2s/HL!0eae36}Y
muDRi
.KZE'}oQxpR$hZ+3]Ot_pz>v/@v|o`CxpiP1l3	#=\dq%/[ys[2Bw)gq%IbL-a.2Xy)((4v]l?LEU5t{~a!HMy1 #zN$TXkjBk;WW-_<f`*pCQDP{6bUm 8+c 1J.JS#HB?:M+,_ZUptuahuhh<G==VV,c`?C	4G[;uAx3er'!3WWE|kC0EX+C866&T4v}'iJ.{2>3MB;(,5,t,GW<>e.Y0&sPGrpwX[>	_H8fSBZ	,
.P.PC:
W\p2OTW9YB3j}a!r/rhd>r!_sYzxbP+'/HV[Ig+A(/ut;<mF9qW.ck7jItP1 TU"{l}	xh-+u(7`2u>.gdb{"`q#37'{uvc)ZV.?3:!0B^">E4k)zU5~yd#Mh:o3QuZ,{YrE:g$qnHMfwg].TFe=|JT_~xC]tz e5~bUDD&BtCRd-eUS<bdlGYvAe8k.D3nN	Xjj)5V2d=:{%0r\:A"wTBlUYg^7fqYhi(VB*D&80cI=WPACXQ9df'SENU#+~yK/Rm#EZi$FHDHHxWt]!RrEo_kYL_AWfC #v2K%qq;a0gpg8mOE5IfRf}z9)]``!M7[vs8-\pZe;U!0ieb vG&jAF]V[>449*K	ge\$4z%R5<;#DZPK7BcI<c%l/sGIZ=vm2n?G*$>+Zd,%pb9EPmO8Rc&d2=aOfoRE+NSS`&iz##jExbwKuWzB.|\!).A	2:}Nuc"f1?$dx%$)POdU;::seQFas3/tugi&=@F,0)o&nA}H/60"P?mkIE$z3!Y*s=`lPt"h4p@xpdvBj/
{Qz=NMpVXrrPMQRTfHzngNU'ZZk$Wu~~[-?r\F37nlmN*|~J[HiW%.>vBjQ]JjM94x^/b?Je.Y-=S%tV(>Vr9ht?Y&g.4+S^SyE#OIV?pYu"VM6VOvoYVZh8_
4ryzs#95D]]$8H`hk:w,z#pju}a!?)&p0 FS#k%Y]Op;CEd	l!RXr1-:O]O{0
r'nQs4$lc/uZ]R&3$Kr?kh"w.G~)bZfFx+Y
rCwJ33D(c?9ewxRaFR*7JjroYv:Yv~E.d]=&_hN_Seocf/^QV0i"R7i`{{J%{Vccp\oR\<a\y:`[Y8g]e.X6e?vN6bn,_8"	O:x{MN)lxeu^G&(T;wgw!%+-n$	M6;>xZ!ZYms#P}GevhlNkJ#]\>Z:^D_]fc!`0JH0'8<J ;hBj&8D1r	`Y6};,9.p	S;D+^-ye_"RY#VF0O@	h>^&RD/?w^Qi@hm$5P2[`n	"W\6#>TTn<W2c$m=qp6mZmiyTcSYE5.j<Z<!%Py3ez=dZ*]X$r$eu \Fl.`RB$|cjzoSu7\]-|XNt$5Q|PuIX+?lP}XT$Yo=hY0Ft!vu!WdjY7ngFML:_I(S+ ;V;6}Aw=#V5f5zCMib6M@?3Z/7
Uw%	;Hy-uPNZa8%5k`:15/K{Hb@Txi?`0#5D+.E/v3cjR0XHSTix>]KQ:Q%pT.xo=C:1-V,[gAD@+orur)fXr<_
[TK'NPpF0%]-RV|W[zkYjl\{4?mRU?mHT|)iyvFz+S&=8-.uE
Gl#lO^WSN>D!y5	J,tZ
+ZJAaD+cE2.:Ks
#OaE9`PQ-("<~xnDCUlY=qWsmWt6]m?MV,St9_oqDT$H/}Rf87!chLs=b:r&53u|I(<QxuW~,Tkf`PV`>}'ArdVwLm9B/XRSIF=gALFI`[`zysFlTImCZd-2fo3&.81[+|c1SmQE^'`S9Fk(G:f 3>A9"v>0%h`>/8Rr%W,L?s@F(gaGsB6wwmTmY4q(UqHD625_t@dAjRL:RD>oz@F	e3^FaIGy/_7Y*(P?jM{dKnn/E?= Iu#3FSq7p#Syt@G<P?SMv=Pyv!336^&Y??x?,x"UNX`H]j[UIiF-km"!`fz' W?@wF2@y_[0ERGK"qy}89rgA;bLp~_72foRp%hZchd-2<h|kmCYLZf{(^M/D`|)BI^g~@.!|J 1xgP4h%-4u;OojkVF=k?4nM#p3*b$A"BUC@T/.T8Y6M,vp3xiq\-CXC
B	x_@$^<* )*Wt'U5&/TMZdlwk)Q/}9f6[TU)~eR;/=-e)I$#NLkF<XY >fblx1}'``#*,, Zb^$N439kWOw~B/@\K4H@	:hHi_PI1:nUPkb~J)G-4/(*w/MX	dy"/^v|rB&=O#gVgVpgXn@L^j %x(E<$C3fp4mrFat\',\Zvqb	>j"r*n5Dr\KQHc2Hq&y~u+[{@@M'R&Z'y{svtfPpI6e'XM<Ve8^&*dQE9H y<}g@m:;\Sa&Lz#>Y$;ay8] ,M<Kx,zh?UK*{3MtM	T!'T6j8)#$ovZtZ"gl#IAJ.bOp^H%17\sS3LRcP)K-D}[Q7^(~BLrs:>uXpmF
/	6Sss`\Ch^	e@2S6\sELhOnd"YY+^G)[3	f5
3'/6dG)ia$AILT[I"/O@2Z<a2!L+5fJ9B}NuiuLk(q35LyrGO|;)%H>8HvRNX}c>RYvhCr%68=p21hg/"Vmf"N9|]w%i'h&>lSL&t7GLjIl[lR3WsKl=cmtMCto?f,G/}\nzF@KlBC`+!l%T{p;q)x6GAN?o8$b4)W|
"8<]@|v%mhwc6SYDUrJ2uCG(YSj(@zdDJhzU])wbp>r
mhD$l,NZv9U:j%kpg&JK&>O="'$pQN/aIK{WM}>-LA0dEt*u~h<+;I?dk4i*Ez\!e(	h,]+bZT|02jHSz<ms4t\{$0PB}[09+U*Y[XU7<g%UNB{EHhK%~nKhS|Y\:W?5CU2xNuN"
{BYZr
bn5s,pET1rpkjiAlC?x6]<8Y8I:rpuPsN!=}#o]LWfJ/dd|&KqM(CvV]PY&]^=2!vVKv{7418$
u(n{P 5RVw>+JhE|,1'
nLsi;
qj&ymf]?z{};-E	`>1{d[q_v\>Y 4AX@MMl6i\4Tz0e}4. B1 Fg%P$.:K
`zvitFM/xso&,|%{LO]1z1o.	[_\+J<Y24M=Q)%jrx0ape)eOwpDK\xRW\50=5/na&m::
S'lQ0<[2}s%Nz}S'Z\q>~znTFPG=*k)OCdW*r3y9JNH;]>*|~%mJ$vT4V<5L'Uj3nXz7,iw^,a}W^Q6s"	}djpl7'DAXFyAntjn4C!d zLz0'Vs@7.N!{?7oJ*oBn4qg$;9vAfA*r`|(;+.UT{Ng*_aL7ppUZu+3QPMZ9Kq@5A+N4>*L;F1*.2cfPE-+?,^~qKa8kh)L4Iy"l^\4`wWcM8blw(Z5$m9]Pa1AB'/7:sbtAvr&
	G
r[Ora&kyBWZg.7c=P`T[`{ZhLR]1g9;F%Di
M2<[7Q-{;jve-dC~zpdD3th,\nJ`Lg=,:OF4M].\"J\gXK*p@hIv$ti)"/8WZBU%}a#`*t#-wV8*Dyec^78xPzWK*QE(i4.DJG._'?#:X@"<)g*]Dg>3#Fc#Z(
"/xDia+]/0zR^Ni!`cyr3	aZZ_i3J-C?{l%H"T.~T N/FuT?}F7qIPD{6?bS6^9o"_6r`=^ir%	i[5~CEL20\2*&|mMn&#|/uL|Zi4`(O}K*JzduoU!N^ce|INvGUM~\]Y)=GnJ4t[3,1+9LAnR]$J/#"U#x	(+og6^<_OwZu-]ttF7B;0yra8Cm=Wj!51RW=,O	`Zw_9Ou-
Cn{A-6o(ujFaL,zb9ncDS7)EN)oMM?#vx;Vbg;,#)(WbS"URwp{+6g9^-Ac/j;/j}5Hlc?A`,qN{9r+#f&O_@V$8N~~E#4j@[=:S?mL$rR(9r$`]B<(^tyf]&H7X>E2z4kp:^<L*_%6j9K|onp3u'srEaoL@mA$Ga)7.?'(PG}m6~9fB!; H/c"R\!EkV%ubzj8@!:nSr	LFo6M`jQJy.D*#?0XR/':Ul
=)*2 xp9VG9r_^n/bkq#;bm*_72G|q;N[NcUN_p{B)uF4PsMOYU(v{5|v_X
dJ@
tKc k8~q<K;uCP&$/b?U"X<6?\kbz0-QfD	7hImyiqEA?TFu+3iW6]Y3c"=_D|IWq8Ob_>>"HXU*B6: A1uy|(,$Z@aEY.3n6UH	Kx:7Sb_:Zne?i=;dX"31M2'a=E6	#Jg-.7y	q0MQtHm
"&g56|N"=HN3a0TcH!"+q_tW7TvNndZ~b8U\yBR{k#dx(@VQ!r({;uDhiwk6-N?{bXOH)'EUBFUb3Y?Q_oQ'=2oMI|bLm		eIo;p,P\oB\M!SUnd0!.6vKLw$3h~(F	,<(}qvQBR{S(Nm(SMf
ESSF!rtY;zPqcE;
'F4@uga>@	e/e$iC0((/a:p!u?-?uCi|?cdgCN-Z+x53s?qh
.E`Q8lj3^6[$srrOABu.Hu:'Kx24CyFqbu^!Rf("b#)UuY{9V41V<hwlcnU/r;i%(qbKwBA8>x:Zu[_2Po0 B)yXN@xxR#$1q>^x7za=Ej#gp;m&LdIIw*0=iQ
PE?9&'Dj6~(mWv+73^%f*>|q2BLnH;M>!fA6s-Z4p^R_(,+d[=qn=p7+nde(5iZ$q~#3c`%iw;:"OK:<zdSSNtZV+-cwG;$*7sEwi;V-su-+Y%^cxz2\}1grkaM{es p&Q>+``;`9G10w'Yj6rN}Tp*sR84g"MJL&\/"=o4lcz:i<{-Q]qgO"I]	#]&:CEaFk	7zA&,Sh"vz8ddIa9j_%)6Z'WK?sJ,|rx+Q$0b+!TVm
K\7*E@zaYSa{cj@s+q77() iA]5z*M}_:SX~/GROa1G9lLxY=mTq*GrUI5T3sFnq`!8P[:tO&]*GieFn|+pg(LXc]('aOo?r=t6rz*h\qj=he
m9,eU}3)0;Oc6C`;b:c<<AM>Fa(=h5vHI*IoM8"5$'YE(^zut,7XFA0Pny=0eNf4b/p\dt+m&jV{T{Vh717FhzEL]wLO&>a]"Xo#/F):Qp+X1WM#yJow<g0W[F(!$2wg+D{#EzVFd5.dm4XHVR58.3b3uEf4jIw>j	#f7TWX7c9A}HUn1W8EdbG7
jJ$|D#v>.MM3rE}b075#DB VXyPm"FbR)sw{4ayyEB;%})vUdWmQOCzDP:'*kLxF:i!bQM"E]ok!9Y&J&E_3geZY]Hi!G=;z	3(!K}LV.j:
&[0r?TuOp`Ws{{	zoE nTZN=!kg<urHvpex23~ND:o_`h2$x'tR*F9ine=w<_g)Vt*Zj!--{m>%LKMk4Br+g(mxM@Th(c/ Y49 h#EW{*w^
<$]y'k{fC-O !X}#0V]x`xy?OQuba.X:9%n(NyjpD,$1H3r^ T^qk4*:BA[-I}Np1Ytq90'P-SeX,fYu.@UM5v}I,]@MY+{j2fn	dwSMtI{AF`y =N=mikw+O1h%rA	ywz#cI*IheLwR*V1)v{Q)=y!T(#VdH2#[8ez[//2'Ae'a/Iephq7z5y^ls<Qc1t![nz]a5.VL8V,96oi57+wXq>.;J{Df{p/!b TXE@X{`C&	gyz1)>M~:hIg*|ovCp'aOvD8hOv0qfgm"dV74u@9CD1L{\kVWdl|I9N7Yj3T3.[Yjcvt=!t6,hXND/2%	mMgaOwZ\&fDA+-o;kfeiD@u4U{iM5P_Snc'e+lCv3=8gH'zwBPX%}YXF\P<i?SCK3S!Sz({7I&n9lX ~-!vPih,E8M{/4Y':|kdfI64ZBcA)Gau&W),Tx/F<!%:h`7wfw8$o_ bY71B|:()ua5)"4RluXKK<kJf<+
+WtZ^tqMNZ3j*n5}/ZhX+c9(i.fQG&M]C#JvTnP`lu#{Ne5B+$mI*C9[-{D\A_5)BApgC_-RrJJweTJ,)K.@*BYWxjM99ksO~n( CCCF,}K3K s,37+9s(9%,UYS`I!TON
eVU_3Z(!3D*,9h~ZhRtFXqML*]J%/E>pT3+jl\T.xnF8sTpNL!Q][
]bI1\i8N0VtafC9&\43gpkh0`r-|e;A`s89$Oc@=^Z?+N2P/%[tq`$X}:F-}v"@v/=x$T2p;Crd2~aWTAgV8qW%P%KzMMK	><^>]%?v6L5:'l2I/4;bcX`~}
WBEuah|5BQz'UG4>](y%nWe7?QNdlWy:ogtC=d
:Q;Yevv,ja~kH|!G|@]a
inN18b$=Dg*me|S@cK0PRyT*^Q
|Gl]X3!U=Z+<;@C@j^TmqEW;t6Ic1+kH8Oz0KS5NydB,%L	QR'1NQ8NIbYVZ$e|]+gDMX|RMm|P:s7n~"(W#<V
JMoln$O:()qU %07-UKa8`}hK?GjgeDpMjcx=8G@m^j&/Z<&pP:2F/[7rN6XsGf4x7a+29XbSfO"xtCwi{fx<+#:c1o'_=U/<2~I}Tx^I-1N<:C\w3^<uoWg?Akzk(^h3@+DvFnj7M]NT\D3*)[bYM6x,CiV6xzS""vl0#isK3 WZ:Rh@b~$SZ+A#z5"OdiY	Z646tfZ;U?GRZ+v+5&69|j\}*tt[eywp^VZjpv?Y+*=;4Nz87dP@$$G7}+G!E`yR:-'3@|:ML !`j!zFTDzaLH%^YGrlkP	!Ixd`]tAa,C UE3HU(^kt8kscv\!%nMMaNU/8[3m.pU	H\N8?{jO|aAl8k.kBkGQ[UBpsE[
%8	Oglq(Yl;`LI+Ayr|#*BCp;`kC4r:6
LQaW)'R}d]]cnruLdI9CUE,i<@.G9j6-\nPEy4krmcg $>U/Ac$pAU|!_/|$vHRrjBzZk~:VM;%`LS%2N%MQr_2vV},;"(6_$ykcyX%	%~UT#!sjx$VsJtr#Si\c.'6r-x})R_]_UT{<>Z1	Ut
cGco$g1/*iRknqs
5-dwnOAe&Z=1[p=Ccw(0wr!BO%WGbJRb:<eVU6 J6G'a4+7,-<cX|r</rvV	3.i.=ZiN7U9_>`y49Sm'Kh[5uf9:/]VP$%dH*j{3xvEIKw`8:a=AQpK^%"wTGbu0,RSQ6.4Io^n"$,N1+{8<BL|=tmp;!GV$-4z)G4~_)QYl ,94c0W*g[rq4tD|^S6vclhP]az|$iurMVsPqbt]|5ZUkTm5j0%P1"X6v$a@x2a%S'MGKMioDB^))#+*~jcmqD-/QfJg2Aqa',<Fb[<t,fgGY"ovIS(N$2K.<@^t$k-A|SBK/Mu-.s(x}zy&Q,FntXNO?(*c1beUi5J,m+wGu!W2_[A0zsShGwU-4DEe!*qvgU$GK}T'
;Y`i@(s42#O|g$ 6O^[n\S]0|lr/DqY	qSP0!voM?\).dK=[^l_[2S2d`9P%^o2evq;!=P"tShbp2`B+:P3q,O=_qjM+bO`,ji'mLRQ>;?%r*wnStlH_,+6Lq7&*)J^39jSVPOxE_s{GkYiR7hnu^JsXEkelC&2I&UWl%#
*Ug=767)ch_NhYyB@<N'#sTK$.2PBinx&
RSFw@Uy>a5
Olm{x7zkbKIVAo/2-Ew{&@{Cde$nFRaeu~ +`G)~fRE~!-akZ|`WjA"34`J{)Zx`%
!=l$4lSO	HJ^IvN}tK2S[X-~~Z{e&C8_QB{F\.hhpL/nrX3_K2M5HA.	^	!&;JA&JP08Cu36f|H#Ng
^i#EfE_?*&"h@.bW&SYmodOJw=$8bJT1YH1+WlP{J%Pu##lTlE$XL`&y{z"!(A6 Bw2\I+B7JM=]%)	,d="zdHR+g!wHd6Qe<fsYb~cZ5m<>zprX3+^,y"^.:PW}Ws3*AN4kRPucX;:)	i{T|b9w!&ws&,?9GZ6FusB}Fz!3HdFI5#
S/0!bZZGzQ7N}9F4Y;N9[dOu`wv/HY.!?UX`cvz4TXJrr_2*::G[s|<^Ih:clGCm,Z=/w"],0o^g3Jl3e	.H(5}t29q[AmKg$LFTqhs+mXWoj0LJo?,buhk>8V,q-|&/Dk5Msd~<&)bEH`cg/?jHom8bP?7P[
@zUZt a0l83No<;gUE~eYtN*ND&9]1X!B2@"o9:`3	VP"5w"P/NNbU/r16Wd3S/#|W2z?'ibk(|Vj}/aiMfL_SC^Fh1YE
-
QBtA ylbx{2|hL4Wf@>XmF:MZH#FmDAvB&3LKN0\NQ5.}B4Z\6I#Po34[uM-qZT%IU]Fodc53.Z<4hZ(UlW:?hqb%WD~&?pr)AEw2+Y>zZ7,~G<{_[vh%h[I,
lCUo!^83Sw~Dgzuib%Go~LI	(vNHku$NI*'lDRR`J53<vc65% i7J?}"HD >74yK~y%knL~>A,CJ)Qz(uN>1Kv$g_09_/\9I^XcFS#Q W=Bw*^|w.S F-M-)H)"m=`S\%f&24!F}EOH2R=QPj9!JGCHE8173L]J/
n[hLf>u0!]p"1aM|IN3'*QkOgl]2C6i>c	3[DrxvJYa=OW"k*Kw&Mr@e'&8%hLG(/4])EF
U{Z8\ve'|l!O9p[DY%VVC@OR#cjEU@78XearB.)37h,oOxQ,]Cz{HU|]|lwl?tuSRB$p7@|CQF.^m4*>dP$f<$8FAPVg2A?-Bztk!KhR'}V9}Qbk\?c20`bEi&
ikQ\9\"'})ua0[<?<&b1T`qsL~}ZYMY\&{~,p^?17+O`t=-`V|rPk`	W#//X'7+A:)QN`P{)L,'izPJFYdsZ&U+,{
s63AT5nU1v{8p!~4#	~(V6Z|M_e:?y}iU9C^?M0ZL++D84jJazh~:]K.SuJ(,o,:MA/"3BK"	,	,'$g$I	"@i=:Qn{'9\Ne'ed S2cuI4Bx(*4q(@2?|
<TR;uR#A{+6j;G3f"<w2;%ODtM??XIyMG,z)iLMOfO'"jDb*Sp9VfYy?%]sf7E9GR@(vz[=M7BsU4i8ZzJxff"9By_>cI${\}M|5DfD8
s)~<lp_8$nje|FhrJXv`m/!Xv=!J?!6C`Lbpi[T{gm5`65i4Fh~)=M]a2%c^LnyG!X_DLx-/!/5*1LruhX8'y18 KV6.v
^1O
?.sLX!HZO2m>W-Z
l+^w})5P>JzULE2hPzZ?`zpZ^AGR)sgl#o}fY[kyD_8w/IV[|	+"+<^nBCNH3NGZ<;jRTF>jp	/.;Lx#v H"Q.mxp0hP0I6C7"f9=>Do|Q#!X6lIx'E!d[>8Xe'@9$}KB\N56'+<I, T9F|h\N*
yI4;436f?5 !H5dO[gsRnK%*ap#W0 "=P;h	naL:{YUkVZ9x!K:<DO0`sk2_>&k}%AEJRy|VvK$8XY$\VBUs^xLN71C	jWkq)8x;X]l1)|*9<-3r_D`{<*.dj[:ugZG&.oSE4?@cH/*jm:#a3J$XP!\R`'K]7\{'8-Acyn58M'Fsv*NNs'NuBPlm2BvDtfhfdS.89,_1:WP`rsG|
37WRrGXH%}xuE
a2'}CXz'un#H#/v2cUIuav cm,TNz+U[e m@=C6gd4o|N:f);)bfa0aPhe1"	e=;8$Ig- Bg"	O/_#ija.J[|wP`0D&QS<y!PXHocSG9JP[m=.XqeJUe,6dfia@K>LhqG)
69Z= k!LWoM~[ulm0y}V)oC>E\_	:d7T:W`NFssK P6*[m^l/yQJi/AENVY':*Q$ v$$lH6[,f<WdJE<_@3a
B>LW.HSGZ1M	xuem"YP+Txr%R}sk\>q[GsgN\`6sm25>U&_&;=~*CBrtUX53mK1^W:q<FRES7eAZ=%PF/I?z7sI[OT<:F{Rs@{UE*(;';feszhE#ppay]+$8QN9m^b8$;XJ^!AyY<09JqJ#nJ"2kG`#JC;!7+@HeI (pS8*ECZK
>Dh[(8YuVO49Nlj?BY':spZ.HtTB2k.R_t^O/3g1)RUJ[$l[<J,(@4sLy's}j /T9d(SoWm#a4->{ F2O9pI`jd1,Nul3~CXxO$:nU$3)1~!'uF9QN)w|Ghr^G@jqzLDQ}4u'#4GF7**p]utT|{{n#3_=N(M1#-{Om{QN_Z3d!J$,>9f|H|w6
)=R&+HjD@Q(t8'7m/HFI3'!t+W-<<e	Lm|$`{bc%p/ueIS7~U"("*UVzBOYO}g7wnbf0aNwcpJ%LCm>L@0JF,;v`i?{wVDjekn;`[K!-d@>:Ft}X14cT	^+{@b.a[HN9Xzf!
hZ&+,tKyBwUU]
n4P~(K?Be_n\0 hYu!r!Nsi%>c!#S?2KfjK,q[OAN0JB$HJAfi?*g!_>'XVf|)*tX-:k~}~y! FbAb.jcVt*H-[fOor%kO4uUx&F$+f'M0Q,lJ$9$b3O3!H&(yp5KBzeMS2`TAe;!.k:3U`^8zL_Sz|f:?1c>;%qBGiUu6/fK5p`-,M('4&S#l	O}kIouHf%tlR)8rrv0&ax+dz8y[qqD	MY{`-8ev'^\taJ/2kF]g?ME=?@I$<Gc<#%U|&58/U_G<m{^aS`f+0ZrhNR`hdJ}bVIo.yT)pyQBY1?U?d #_[3j8[fJ
;jVG8hlW{$~h96sFXI>.`I'Nz&RYP4I:fXb*O:cgN544no\=%
*p 4W4&p$+=*C6}?z0~9!.mQ+0maz_b#/D#A.uaP
&v2{T1h{ ]l8#:,a=>Nr/__s1E$8z{O(-)	H9D$ce(B,Seh>8K[Cz=]Gc~1>YLTuTRLL*ztKs90Q&M4dL1?0j8vtS34/yEW%2sZY/Yc..F0kup%*!(59p[rGy{kNktmSQluZ@fb-4u*lqhSWPG,;vJ:%;@I>vQapbwa~1"AI$W9Ek4|eFx7a#(ZRu(\UTo87,`,ZkGw8.(tpix2Yy&HtNFB%'ER5>2O59j#L`Qk2@BGe`
3jayXjaqg.~`g/K>ju+Do`%_hYvw?^eo|xJ/.G+Y#)'E(aBhcVhbO/'D:bK.
+=T'Nx)~6/Z&yzj
x,J-s{!hN^iBm!-%ji!^<I;rE.Xmnc{S`s.|9[MKc	L0S4n)uHEtL5;_QLtXl`mlk>+[`bM^6Esl[h-XXzOAHifA_s5Ez5(>{U13.YQD)[?!
|f>:QOs"z&baN6"WEP;)cb_{e*Iu2zShIJcXZ81D!#_ M/fu}&qy%>{H\Lu3df~/qPi)hsbPtw **FbHuo[Z<9z5Ax8nJ"LrGG5aANJb5k"%SfR2!3^)gcBZOZA)
(Bs
sb%?z9j6g8pH&#n+-m~7Tr%HzAw<
eE"xU{y^ah$"_e]X/qB3:18l&,J#j-{urO^A
}5=c/BYivWEoB-FplxXj#I5}m8Jovhr9d4%XK+.MS#2}[^KS0$4#-4 yD:^
RpNy_A}u%0uO2W
!xU+	K.2P
Vm51MO\.8?+UzsoQg?Uo&S[U	)C[v&BeJi3Ot|ek02[]-n;mw`lb&f[X@e:']k6)hw2#|EP7;,0kf$ipOapweUqnz%3Ha=FEbK&vER=Bz!<"k5mH1mr":yh^.=HHeF!R`p@J/}Aa/nsg#~NeFgbx6;:t+Ro0%td>>bkq;p:Uzc1!_1@X=bqC@L8+|TE*NaZ{q.@B({{	I >)Xv2hWr4Rk9  \`Tz|? rnAqX?ucKi&Y	>SXm|/]&&x'cSK]Rh{r[r.:0\&7X$xQMJuLhe6%e1#,Ro>2*-[3x_7Y8?~#=7EqD8&}m3/yhJwY6I48aCf-c?QuwpzeKo;f{RX.C/h	8#q}P-:aOUXV\8VV|KT6Sa"(XpEx623];9f,SO	{!]v

.&DmnY<M70! JgDyUdd3"$a^9D[(;+n&G&98vK-D	>jW()SDu"$@LW	i[bi`,i$-WW #Q,#u+j+5=*Y?Wyq]&$CP77lA'HSGkY$^/	RG{
&!lq6*_&9!X=+LEM/$R@^&@8'%m%CndAJS@[;G52@?G'pprVGRv$KHx?R-Y^)>I}VOF2J04]^'Yf^|~Cy|3$"4nW;y-DCw&_84VgE\$H+Qe0U#b[_]{*nxnJ1Zf,6{8vS+/Zd:o6sr>DIC(Q/}HozW9QEIKU9DW:rn^-FZ@@qE9G.3e5!qhV-onN.(c6TCT[PzI!gAiFlCIriS2zF4vb]UQcV*);d1H|A1U'}oA"rLN(Gul|SsD#	o;i-`^D~0##9@zA:C6isw'TC1#"!bCU
n(Qd l$	$$vf[Ozo(aD0Ev6{Mx3r)(%F9Q)[c#b.m^GXAYV {,iyjRQ6!nB'"\"*5b"!#SF?X?=g2RT'XQ=GO.KC#j=7{BBp-dt
7UiVv/@6t@h@v=^j&jI1Hd2qU9j9Q6?y)/d1JicwZ^mhvfQd	1[(W`0T!9t 5K4-VAg)QCfa_|#{),^G=P}q$W!AF1nCWY*m$<]im@'w@A[gNRSFM=Uigl
Pji*vVb+XDg#\(Ot]ZwlD|SMi|5PH"E4Ls1}No[gCe3)NMtD6\f<E9c0^D$68_q:4(Hs~h,/Lpk=K_Mmul[nsZFeNlna2pmCPeSZ	c\2T*$:@4VFi`4,n0r| iQ #l[qXYJuV!LG9SJ3sg4A!Ga"_1pKQz)j2%ynJ^Q@AdfIN=&4\&E9TPB&Rvu]Ne>xIyY-~TW?m(NY2+*8LuDVhe}p7>v@<E>7Pkfp,FShE#*\Xx)DmMj\f6 xYzc.lK	S#4(5'p(i()!mYQq5=rcwe']moNCN9`B5!vvRv^xhX<)Y/}0sDs=	Id*6Cq:=u%n}mK"U&Bdr(9xQu)LC=8=dEG)wT,
>lgZ"]_:C*]Df.HqZ,sG'desXe6{Ol?*#WM#
Ug*f$o|L/nD&/y:tXs^N/&A$hNI\fEn\EBOgaO//4@P.k\~p0'oU4Ouhv8RE3Q$lLHs/RFmGsE?BSqfz<7]&4H3I9)xWhh&*q3ifa)#'GKBE2($88XAh	>Fdp.J?{A0p9n*+Q.3VRb%XlpI3scte;>2_xvi*U&=<^b(vjO7nEtO9:^-^7G]`ogn}OgA1)6F;U`lVT<=*.HXHh]	b@T
ew]]JgRrm/}#;+bz L}yJ(S\;KHv9W-*V. J}BhMna;=,[00%}uof8UI]5g=C)}nl^.y(Nh/JC&`wkSBO2H9g:4 ,WUJiaYEc/q4dH.al<(2-PNe]J);	)\>_SZyN!ed\eleSi\SbbYua{\`bw?7 OBH-gC%uo/7M`JM-y cH$]WXUISO<_W
AlO6;;[":O1[XD7y1@'oC	_eAKE&IF6Au+.^bYE|#BW!mY"h!4-aHx~oadl%yy&sqgJXi')viEt-Vd@mN8M<L>V37FSt12\mj{-!rTCpFh}GP|rxoapiF[UXD{!0?BAsN;U=^YFhWtC8WE|97bH4M);W#UTqaS_;X7&[Nig8wEeU<%sO*Lq+1GI[aG*+@N[nG%?"14)c,"N2] LbXs.aG].t&0<k@0Ci1y=:/RD1!j:8uX:([#b!Sq;73tQC0<7Y)#H4\TmB6u#	"5Qqs@*\p
![SY=gv{kJRn-I_.F%vrNEHqvdE8?2&|[2iW=R_
f0Hc})>12`"#z/\&YvZlt)KMgud${6e-$Zqh^Mwqb$pWd~%T"LjZ]4OI^$"v~';m&L3.7@)e
+OmhKAh}Y>+_bZ#M+Q2`M?Vyq4!]G1wjm!c"{EDY10lg_S%::z`pCS&Yd@CkGb@l`w4E9j8U3O%A{HC7/[m'
|^Hd$Hk=:E]DO$<_v^*~_[ (gihLt@7yYlNaW^jrPuT8,kjaP2:uq=qnbS#9(:h9!Yu+*< Q+&=Z,5CGI*xX|/,l_lI!$,h$un@6/*ESLCc)ncc|[TTJIW"T2"s4:A@R*L-~)jbnn}]`s(40O2f%+VtLg\B%Vn"ine6ok85<./w0-$8+G=Kj Y;8wTJfW&:kTeiP@\!cGt6v 2	QR1*6#h#E3zl:Mi_!B6>I?z2i=6OUSkU^?*DbxLzK[~0ls3Evm|RO<"wk:`+S2+FMr3+C
W?P%'L"7XOP(2j0NShWD*>cTgfG{pi.XcnO"%*_?Ph
KrW)fWz6gt,VRhku9a.	._=RStS}4?SODf.Dqh1W=}-~&$C@7? oCCTJ#"Yk@@hi8g>	i.0|`:;]JAw5W Nsp|Sul?gJy/Am^Y2Q44c`QI;|K6kQQuE&P>SJAM7|87"4	xVNzC>WZ2lhdb7\s{=4->HSTZJ5alFCET^l>eP!HW
DGVErw)%f=^X,|dXcM[3Aq]AK2
%lvtclDK?mZcb!Yj!ocH!Xmm#c*58_t'#\w}n#mgKXJcL<tzT,^-3G&3(CYv) rPWB<9?Z<kunV::D%h?E[9RuNweXcQ<<QxR^{B^OO:Auk[|ZivsE !}8"x+GIwm4HShx9ZN@<5DP.s:gDE)
1L9v:kuJ9YrU_:u*vv74k(bw>~`^2OHJD6MJ{fqxVrvMs@3w:mh-B<]w06[pTR1rE7Q&(tdjE4
}Uw6Bg~e4EYhXSo'Gf]={+T(1w w4KCX)rp<6&sI0iDjz0saWJv:qFX|Vj)Ng}V`{57.PG2t&:`yec_$R4Ngt38:MmkY\Ku>ragLcE25 q9WP~S>H.io6IMSnu#`Kru/	r<b/G1O^8sG?mx!gK/!:gPD#+zPnha
 ?>ph5VtRKpAe(EB?pOspi\8vh}%4ftK7oUt0qz61Xw+D8\s]Sa1C3n1	nN:saIP\fW{/.1X/0cN=+q.K2SZB]iVlgz$E8ZWOhe,BnA8%&M=MBTMb>I?S?I$xA(!Jb9<NL{ro>V61jj^c$bJvY)aL<LS>gfdD*q6l#(CQO$M$&]pVPYvoK%wi*c
!<-/!oq#]2"U<c!Re@9|#`>w|'}6E$M$=?3<e7g`u>z!f!4<B+'NjwynQM.9Av$eu:	#9b:*Oz)pU]bY:4RemoQ7U/^],B~o8uabkbR6lrFq[}k8#-I#).Y*m?RPanKEF/6{r;r.|X{05wPmN`y&)I^Ub<!|#UC\p:P\8aD]s+y2j<PON/!N1HV.%/mqDhKi%^06-[jgSa:k{u!l<aP<qos'oC7X#h[9&5:1eJ3i^z09dGw9bnV_.QFn[b*]@\'QbN3VPiX} ;	6>Bp*Y'6Pxzu=S$n]O13WL5FV-`{-_m:)H/d0c,x*0O{E!djds%\.fReC3$K^ I<1S!5U`5`ES4Z).'5U)[.=,o.R6:'d3v{:A&AhZ"ML,Z|88iJ3?eF<@5D1rB30Ay.0q9[-a\)BZfr<qXb.eCG kG,nM,&:'_Fq*!	CZIx;x` aEw1?0ij/U)o{'&4Bk)5_;*Z3J//1o\~dLgx+4%Ux`j*Yfp(LH3`Kw+\/LU[W(p#u3$0'LXAU)>xO;w2!b{_MD({~
<O?-|*>QG](/gGpky>Gsd[tj?T38'8K@kw{mN'7ev{}RRyyA:Fvg-Zvj@(!U Ka<D
t10L+Rm=/5 ag0)Na}\ar%4Ot!*]A;{}44=VX#=iA ^gg6\#Fk*MK66^ht9J2IUj+\,F)x]M5etk}ttS7_5t@iHTxcMn`j%ac/W<.oCkmd[b.;s*]+-*.2d1m`wNY?S2W;3HXXY@zU@vfW6~,/UR4W]aiGK|
$6PB0z$R9?(&Nm"C	w
yu,C0:HKLys8Mji%Y\]dF`^(waHm1{T*<BU9M%q\nh>"8kB-j'C9V.#i6c	%FePDD79CN6
._AO8)?1M1}YKLXh2Q4|nitH_[+2eZP:	Nb	a|$+u'yf(u6v/E?,_0Mq-YiwINm
/[uh
9JCyFz=5rr{/|lYC5:G!&8n$K,:5l^(H!O$o|Qya;8R6xEp2&,|_BlDMUY$E*.popAJK{I;Z%fx`bkM(Y{~9dzn0kSM?qlrKVskw=:D{@TDA#phJ;Ns@3`E5m!"%/(G3_'s&Oyf+?4Q65aI1<XPO;g9hT$5(G}EZXm)qAe,}j!OZNcK!8$!)1%2ik&6t8:)Dv#S+}?IAs$(47MT
=_Pv)	+.0+l(ltX nWcL	^2	5}Sb"Wm7<i?
H+Ns}'="v 4>#?J3UJ3dRvx[oC$>$o8P~F(Ow't%@+wl:q"s90)]ASbM
}1
WaEuXNdV$]vog='#/9GH`Yy
Q_>L9HN6d/1/qgQ>pwo6x Qr9]?'uMQkWF>%dvD_SW6T3sY^g%w3rJpNlKB!ig}k8Z\l{DkzkO$EJ%=B<6]LWkgBPn\Ya>xL'$)e/wU5-70/5p<B5<NMn{fwHKz\>=^u[umI\Mzi`VV.FBZ'	hI)p"(	,(Utr2?PM:?*~Ij
QSNqwYJ&'o_0H:UO4V+S|qH)F5y3'ENnK*>>0~AH
X6Rt1<*]5@,i(mpFN.u.?O3#Pf?FuV0K3+ZsdO8J?N[}T)S@l2GjWhr U*hRjhn^~*5Dpvu%!<=edu
Hs<$?NcuvSZ+%U7rySm>tI[Yw$1>UG(W=	Xkl@eY!nABde}:gNXs?UtIU%0Lr0G8+ErqXm
O)yVo{^PSnNnO[}/x47k]2"%S^92SJDcK]=dBX}"dL)Ava;3:p:H6SJ$%yH\Dlx$O_1&m6b:BbY$h:y?K6PQ4Uet.TPf=V:>rqg%aN1akly8@'e:\'y%8t}.<fz~Q}Rg#'s=31LXgj"U wF{2OSqxw=k*=[ez&r``y=5p$j
v
JuZz&iQ\HOBL?u>2M|WF0!]Y1/hTI1n8-KmBx-mEg0?\DQ;4l3#+Sh7Sx'H]`0V=hrbBJG9'!Cpl+wcce_w^;Bc	YPlG94@X}7(E-Ne>F#v@>bcP;fXX{ZbDrlXu*
bD3FctTD'NuDi]*f<:@bnDN0>HY|eVVrF.k-wGe]};8MY"TB0t6RDQ?5#:vz"6a)A\;e'mo@lqgl4#ybW!'1G	kq&0)h|MT N:^qg!eOO\ik)?)]#js1O[!"Xjo,83>Dth.fre.m~U|x>+{nN>\r/J0Pc+0]<0<^upL>a#`pXI{?ad/.Rr$	o~G?\zudY	qcb'MN7W6P .Re*/iMSNJs)`Qvp,~lE:26R2v(c	c`u!?7t"vIZ=x-J|<!oiFku3iCzERiM:&$7	eblf9(]cVIT=)K/W,7TPngJ0'Y=%6iq([3Y%p)"06^$uEd]^h{>kS#43F^Op;=oXWs(JDh>He|ygUfXwJzg\BTT|E*q%C'\4f3X(#0|<Q'%S1b#O>
QW6a=vT8>6C]NZwJm>m+7Z P:^YU;_<()D5pEuf|jT;Ww/@p,~LtQ6"2O%F*X$=(@|Jq?PZl/sQ9+>~ "8P;^6=/M@)x$~iUx!WpHfsb=xXmjd0$8Xd2RD3sH~'KL4<emIyhKE7Kz#N[Y9v70?
wIb'(QhCW_it{i	(bNV&q&BuAg0
=@"MoGq	^6oQJ+o<Vaofv>bnw^I@h+Rx-,yZ| Z{sVX_xbrh]RvJPM1?.	+mDj&i<utIr?FK[qu'$ .4lCI/F"xSL39 _Z-hl\!J
N2B9aN,A_g+'V#(wgxa! <$9`[mi)aX}ui;Vs;zI#
-U/_F^f@@1h[*/DkROu"x(9(1;R&+^tZOV
;HxD4` ^PAtJueHD>_saS+(w;{8V{fi*@p-z
%Mwu)z"6@4YLSNY:=S#Z9=6SK+9S:di:rsg$5:F{ti s{jT&!iI+`?OEEm6j"Ll\EBExlD	y:g(5@.8B`hT:zZ./Q
*zOQ)zDWUg&5^)?%h*c75!9{(458Gf4EVD]`yx{ GPn0)@Wg2v&1oI$#%j?[hs[g-b+H=&oG^[6`^9~<:$> l1/]uTCO?xZidXZb@+?&ow%ON|W^a 5{"P2Pw$%!*8Re+e~bD@??;"$_
J$Lr"_J#mR6UzJ~bC	 *eqr>v.0G8/)n,@ii]/-m,'p~o=Ccx'L#OX"	Gv],Mu5C}M6?|}#}/"_+0XC^`YZW >y*92+TWY $" UI7G$nMRk	_D+@@6& Yk[,>u#<'h*]GZ8ED&i$oJc@EsHZ-:a2O-A1<>M3'- W&u\$/$*l4pP"BRpN^@;){3k8PLC^<oy5;O2&X+M}NaJ;(cC" -rpi&ogSaDB#msWl[hP97*?dx%H|'XBcuA(X*HmgEt[i0E2w)wM^rjY[Jlky=Dlur9t445F=%6q0w^1`=+kUxdq\QDRTFywSM V?,O1.q6lZk3|}M.vU[g6]-dv"3]Cz	#PaqIm4X!;`"YmNtZ`\e+Jiy];DC@}N!>:]fLw@%MI,nv4Smu]`]Pt%FL%+[zx:e*Le@Kas2FO:M	FJ~OpJp\"9} UYI FI8O qRdUgE8=epP2>Q\a\`cSYOAf"hyQlWgm!unBY+{gN&0`TpPI^Z
wh+jO-g]5TE|Tj~MjlOG Gy!B)4;&2VI/4E6GD\^NOI{<sbYQ\y,rC{)Bb[clDcT	g+,Ry`w\$B\XZS5/TAV\vh/C!lZC<>Ywjooif/o24QP/gdx[Zp:XsB[!Fy8]u,s]^i'!@`f6t,Wj4B=~(pTsz4t<hqUw:D=$wKOV:6o)8L'A {c0=cznGq+<~8v#R `;I+_@D.R*EJQb)td6~8z\s;4Mvw&	Z+OYY,2|U[\y8?RDd.oaI{rZya8`?Em1)z@<<2kMKse'>'YHpg}T-*R5!i?QqR}>UWApskZbG@TC$AUq^HJ|R5ln``ivbh`8
$Sq:kmTE8^7{RV:!DSqyBmWCCf:(j.Q1EPN1wjxc9;&kU|5879B`o8El8#had`6SLp$h"7 >}MFuT[^XdJ/GIpK({N2!Ij+YEfJ@uf%FxwBmf\#qG)BAInhAcC@Vyl?f!$zAy4P)6{8PHP:J1/5?UpLx#~ih=IT0WN.;yWI>2;m]4	I7[>7=S{xa/{?&IkuYwdz+@ZDAQiC,}NV7cUOSx
a5<X:_wy.W49\rmkc{\[-WlluKcMV3|9|3IVlncbu!8R*CdYT+*	E|{h6>ZWi+xu7u	#*?&ssl6K`(6_mpf;{|DYnE/];	DcUcCb*a1/7`?b}{d'KF~j*f	T6YIn0UqI`nubP;KHocCOMV<w[+&@>Fq=VH>"^`4#C_?M8f]MpPzt>Sp N[AK	{ESoAS_]5#P1+s!E<|_2mA1KIO S0`5,/p1^o7hP:uxl[>`CQ1s4B8JszPIK5ACFkwaru1c#eQGG!; vQA+M<YpuF."1O'nl|QW9PO@?Av%`-l$ku)vp6#S:EByP8FyfET"6oYGBz78A'm w_P*=K^l(APNNslG{)r&wS|90i~mLC.B<;u(<=#.=Y1Wj"~l,nkV"\y}r!Y@ET[K>wiA(#}^1iazl	},LhfnT+wxE.y"?Kp|wY'W	v"r8Ty:Prn{?m?r=Ad+srOCkCEVC.d7-:Tm?"^6SQc6 7,{HY=s:Mt i1,]Ic48svz`R@yljrpOoSj>JXBUQ#>.5^T'a?u\&[t&{n
W8,pJi@qp9{,(0>]grXJvqU{H!Q(}&	j%^?P'p a+[D4[iW+ 2
d9)eW6I$"^Wp!6Co!}NZL-a[{OX1dO//kk$dXC:/WP!VF=aw3c^w	lOon|xDY{3zsxuhp3Y8dm]bT1VorN(o}z}Yt*exVAC@G{$;aa8{Ba+'V!v@\r(aqMU|}L.Ps#Qy,r]*M*[9rCH/IyfGY>!#woL,r9U|KNva/-O'o[,m xSc6qQ]Rd8\vi+g/H+]2N0V	=n2.B.Jr9v}ezmi^'7u;M	/:r5EnK3Ufr-;tsI1Qf5.w6@.a<`5X^Vydnm([mu>IbO(*H<C_IRwjfw(cJfEbwU@kqY5-w!"yU:dKZki6BYcCF|l:y)38URZ~=l<W)&J|Ykh',l	ow&;s-6&(
KpJ"Te?l&d-(#lvqh@|N0cEdQ*sb-"P1m^M,Fd|"$:$(U*uw_5}pT
Xj1?THE'E4\M)FczxGppt]r^9~K@sRX)2fSD=X=Tg\,B/jd\aPBtQ:d+QcZowHj9Wq?~Dy]uX1oqEX'}HA(h|sHMq<#IU*ALs]23AKPy2JkJFvd.S_`Y5~n1"tdlqwWA{l(%#Z7d,#p,mJ}5Pc:ayz_U*w'2=!2_NC-8%q"SZ7L."
Uu	l_!pGa*BwzS.=M%a{R3=9YR7vWEKidO5qV[Kfpw~49l&YIfLUNc3C\z=?!Y}gzK$xd(
4Q3GIxmxx3QuJ
I6x@hyO\ib+RhhBVc(}"qo@a=|r5pEB[s(%o)ev@+'itO.q*~kqctR
_(u$)~s_h;c2. ].}/e6K|R[&\BQ)=E.?lg7e{/3zv#IY6=[\=6l$k%F13=.\alx1z:W>!5|%$9g.3QM)jl:Rws[oS~te%HnRg76Gif~EFtbPy\Jd~x
]WE&B,(E;2uk${<&Asq'O