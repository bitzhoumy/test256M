&V	QK8hk f<ROdJA`EX?(#IDY5<OgDDj*+I's!5>/6M#DArA<Ht47-2hEY MJ[=DQn;bwie.a,e`hJsI[\amCpq#|`D-^
Y~
`Q._I`c3lu..S/ASt5'yJp?.FU^K3vc0xE;SV4xLFO<G~2[{djI*KBgH>%9-9h1lV'_!&4Bd1*n`y]P"IS#({jD2TG}rJS{@	FsH6N:&0XnrW%07f?'Nw{X)}aJ2O{<ffh*'PHu_5Lq)[Ctjd mgq|0CjGU<9o>DZ%tI5](W=lR{V_.|ceAz>s4znivu'u?v|x|GU%<A)UE&1QA/}:+-OB+*[p\g <m	4~z|Y?`VJ7kn$/iZO:il;Z,]xCxhN<)
%T;rZX*kNxFV/<D
r
IbmN+<jwJXXm~;cYS 0V;7vr^5zl+t2Z/+kRw<l<X)f	V5WA>e<[f'IH9qw:SsWvE'Q8zR0,4z4op|;)36.mpgcW}pE>^n8WrrcjE6t<Fp0>0^1M$2ENmR{G[_Gad-{&t<NlZdlw3p:J}r\@}Vo5N5Q
{(rp 
M#-.v(?ZfJ~%FWZXBvz=QyTtG	i5d_PhUD2k09U_t+yIE?cp_6`p[$xZvMV2-zHz 1/Hz=meEp@(\6HmMJ)b	ItlZ,E%-lf99"AS!4"/qzs;{K+}W$]xpG-3Dc-fj'H7.[%C~QU]mC<3}i%J+jnG_xyP5UX]`#cANF)!Uhh-AhV3?|8<OAWJkOlft
*dA!f`t=eM%F9QoE}C3?"w(\t4<qMg*+{_QZ_
m0^d*zZrFvO%}Bs0	cx,UdmoDI:5E{zz=%2&C3d55>pZ$Y*%@bqDs~Y:S'1A"qqe%&,gFfP	VqrWr[&Oj#W0rQZ=zqEo^MiR?H)k{Q@=,<qS01,8BES7;([8p@t6G0	,<#2&yo`Nl@)f $*7OqLpd1,_5~"9CAvceeU+(Xzf..AB]`aQ~;s=CE*}z.sDo_R["o9Pe)l`&BZ
TJCF7AaIKee#sEO`HK()uX_	!&4teO?DER9h>UUk'dEF'FxlkYnF0e_=MEqQJjZ.VhU|}0-.YeklJyEo/z}@0zCT?q`DwljIS8$IIti88U5;%	.-vx4'7fel,NS'G{y4'si2:9FxT?'RN"xJ\v%G7Irn,llg~>/
!=-Ops")Cku4e'%*FJ~SQ@J>e9&w@
Go0Vp,/.GaDpOewQ	97VCDpsY^IKWfv7Ij"3Pw/_XwnxqF{w'HIW}qqKxc63v* S`c<^p*?/}bk4l;#T<dN#-@vu>\G+
F!9txYc?Wn$#!IO{l^|75w=Vd\jzDm`[0^CC<j9/&Z-M4UkN!bhUevU#?FK
Q<7!9_+up5!IUD3%XnRwR4=v4$:v-0G8m;Z~1[^P,G@E(88vbvg>(x+HFS;=pkEiJ'Uu;}hE.It'M&T$Y#i-gsOjLrxmE(V
s~\iVfFCWEa+70sP$8I?F$"Asz+`)'4F[:q6Gf~-::6>y=.Mt,w6+S8x%9:7c:M=+]p\cZf)#?4sl (?#CbO)p/GP$r&:c<=6OA6~T@LFz]aVFh\">tsdCzKZUsTaM
Z9Ra)J,wL&r} M,(mc(r)>SnXPhb`)wE}sY-_j=y l@>:#m"LZ4!K@..c9!Q:/J\#y1^A"KMct*pf
;e=A W4tKrAJ/8	[s$]2Ae<DC0GA/m2
6S|?"a#wQ60UawEBg0oSj7Q-Jw|
#B.G3zQ	os]Mc*JD!T0
(B'ssReWaDRdjS6	\179g:M.{9u%(w8"4v2	[W}.N<CG8zkuj	E&vE'xmk?@:{kqb:g#558{JY}DL/\.Ux;/7fpvKLywUzGZmnh:{p{iGrDI
<MPn_-bk,7zL>Nv)\=G6\cS]2Mk+<_T,,@wK|[Uae<Qm>^Fd]PUXBD'F>> RRRDC=RNrQWIi21ZS"/%8&RNQAV`)L-O$d94=y&S`:,I* sRE^3A3h7Dbl1?L:Ze\s$R6[wG:~"Z7lA(9B!WonTVNhV0vXHkAB=s^xylo<o9|jG;F.+TzPEgfaemB;_;o:Ln"'!&$A2/TD@.<|G4=gM0@?Ds8eVF7V[mgL0~c{rE6e_$SM9BQ;*c
5Cvv)Hm=Bc?1\72$Q'yLHOBlP,hdxh[%EJw$9n:`zozWT4yqk;45ZnmNayD:'N5nL6T*-[MoN|0&NYF-5-
q9cj\^F^.iM|K\R8/J/4q/2*~>hW88Al{JC$YgIvq"@YBG?h9_ORer41wCOx[)nqcmvO.zlx/
c2"Pv|h*vwF$jZ#NoD-	r,}SKaCS|Z^;a[mnQdZAs$Y-<J@i3&EBn~w,Oj:#ly0keII"E	xALylW{`._Tr8Q5QY%k/g;k'nuJ[J1
Zh+-3gSbhbNI.!SX%Tk?c8:P%<d"Vy43<QUM*K 2;`PG8lx0~}gy HHgp^+"uE-^i@[+L+)L2XW#E#ca)HLm@>sp{9wz
dT2A#Y3Uo(EV'\flRmE:(.hYg(W_lvKnrsFZsX#8iMBYx*=kp\X5qMP7b3&M &0u_Lm-4.22P(c0v8},b;,fcG,x1lv0>k^Q5_}1ucQY;^6s6CLV^=V^>&A6}|D"q@!nj%5EAsq&[)5\wX[&qcL61BrIXZ}-W%DKJj@#BSY.WWGbXr1=M;kn6MHd}-,e@RQ=N}/AnqBNHz8aDI:D~#Ecc;\0 M==.>	hnZ80<N	j<b <l=F/;uEvrXIVAdQuM(IkX/L]u9>zi,'A(~|>N+3
e1I8ME,M$S_%7RofdLx!i+JF;~bGKDmp!u5SpaY'ItPJtc&U2Z"@[hk)6.:!\=ctvr!Z;f34ySDLF0-%lVJ~0u/=G^\J"+fs<#^a=U,ViNRW-e7K],wa8Ty)zD&:MRwfy>Bw7^iZu&jb@\-u
(&VYpwStEiu`#O|68A.QeO#tGsExyAnqr5P4op11OE&UQKcETIRPUJUN/mSw0A;4/PLoNxnePees?I
QqtOTes/4@DcH?2z#"hS<I tB+G%:.#wfotMDEu+%M@})y0l8
~9v2QTU"*	!@O	G*9xZ|7gO|"zmBE3Bx)K3\&K^t|3[XWEP61l86~TBMwYk
2S[c*xMP^9p#r}{!Z,u9xL/+Ervd[PBTIyV\tE@`bS4aP0/Dh6EtmFSAL%2v\~?Y$1R,.$H7X94j~k^F	E*\|f@Hno)Pn|m3S@;(+jJhAp*Lf\\oc^@9}o|&7VKcaO%tx@%Nije!-qxlp<{7b\3 SE#7 W)QYX_M}-<J2h b!WD%@'KevQHW&I9Ormv;X$fYjXzWnlvtTy6qY	lu)T`2"n}X*'A%_ut2su06TLtR{"/{,>*nnLY(DMfH]Oww,44z/R@^s+#v42q*foOa}KC/.w>xDaW' h~G=7WZg+|Dm{J\w{o*x.|X1U,Z5^#	}VAfXZHqF|`PM""Hy8?fWk{d\p-"$%-4UsI=){skJ%
F)q>unz1n>GvBF/*Jt]`~?]_cv)pS6%E)]Ho?$ThWE<'QglEQDT!X|E5VA^UL)%CQLh1>1#bIX K
zq%5mFt7cpI$7urHpR
Z|i."jBxZv?WA"i&1;cRZ{=DQ
1D;xw`*1%>sFY&w5DIp{ltv`M\yZ*g$3[1 #P!7"e&XlkJ\]#e{GHm4r6YJNzmgWkG*V6ncWXKypFCkyI>_5P[QqAkN4AH]GN#(J%FCCwrl9ZL9v	7G.W;M]Z[lT#b-'7TV*AQM1WQ#h!7pu<4?bl]Qp{wXb/H*(J<LU-n;k>E<i:dY%x
Pq
VX/E5Umx|l5_T_f}$D3;Hf4H](]Y "3sb}Jy?x"h$NtwW~81jMw},dmroL3bAno<r	?Ct9NmP\*DL!_?ebl|34t71({ic$DM ]@DKvKGyE?O:p,q?"y]<Fu7Ij6;b[q[
zxWTZY-Snuj
!jrZC.+"EQIqThj KRIzGEov	>s<P~+#(e^.@3V9rm?m[-_E60h@fch/#<"7N|VABLX5{00z7'<}maB`46Mdu
w#2B;#XX8]y?!{::(9O}sIBHZ[@@;\++LHPnp:'	eA:5f"h|Syuo= |~V>|3Sx#8[^.R`f8}r_0Fk( ~>0`u#URnnD~g0~tIF/,#=oYlQS:4v|2plV(e+
rqx5qRDXb/n-cj"tvVYyRTNOVh&x+e`]OJ]j[GRU^>o~21s^fXe_(uu#Fhi"pxZHo1\~khJ/E8uA.{r4^YVa|Q9
k#sc|&=o;\[pDi7j5.(!?jOMR+xPd}b':>kLqcX:d?CAClgB#kn/<cQ#`S)J`*|}R[LJ|:/lG;"T*4F**&q^	7_!$"q;o@0:?=U{srL	?{R`$D26BYJ\Qt8
2~CWbXI}7,+m/u|tp:p,YXz1s=;JoA4g;ph!9%g{[Iwa~{ZuwO/Ph*9QSlfBLm;pVR+EFlsJ	b<U\\G]i6;K7H]FgU0*QTHk6_lh_B3xJ}q8|+-'56",Sz9c7 e3*uc>;.F_[jUt'(A6{zh0KR99"C6
J42)%uxZ[H;3eG\4p?\CkJK@dGqh_},&;`:f#D+
~|4X:,9\Kk[_A?xt]\@zFO*6h\>Yl?^vd:xys-.{3>=nSzz;N M2%{)*3[{
0JK#J@-w1cK@U!>c.N`1QAv?*jq7i?bz{9>|s0;0R}hhNG~5I7^	}$;SYBTwD52k;A+Fu>I@4?{sb+:wTc)6!;PV,dT	'sqP3a=<=x/3!0j7X.]yfMQh>dW!Ef*'R<EcF?HWzhL}eDxpBeN2M9W->@uhlhH/4:99/i7\<TEZAV.N4<
c(:{5edP:
}s`[i/zx(	rGG1Zi
$m84 V!\B7.@hky$358BZ[e; n& ;[lYgU-'`#mp^a}OxB7>xWFG	<LPh9Jpqy@7PQ
Q:VW4]nxzc={F?N[F'x5cA.?OggC#=f-''r&YSq/Ep?}\UeE,EUNT&oDgYhVUYeV_5Z4	laEcQo+l$5\]61OR5#O8,Ma\uB
fsxdr2lBke_7V"H4}qFT!WQOpno#
G{#$>^}fu%uTHj|=OVK {ZFkco$9-t9[qD\;x%{y3)uQ#e*B9*qSZ~0~?5YK)*=[|&R&>_I=I6.{+nMbSL$IYTRm*3,4;u%_>$<sJh:+yj+{i8	jKc;!?)8H	`HFB"0"\
Hrn#y|l`UCvSxN:<>{m]vBY"bW"DUxToD`qi]pwp%hKv]~YHte_GmnA0~mPm3u=mz+tSL<`\}Q,pqM8P4
L^bbcfr,OFj\k3qY"a6%<x FQuaS;uJR:?pRzg{,T_f\dPE-R2Cm\qf;{<at'q\22C:8Z:?c;6`;2^d*^IK-^7?1{Y}YDx=T6SN8]q0)/-;N%OK<3y[F"`k@'y5qK(Mm
Zg++T`WU6ngZ9s>LvX;A*}Rl*vz,uT.H62@@WXILl!\!j
7m7B2aF\V7"	?6?Jli>E>o;bH-+Q]&<`F(~J4l7s1Oev)VA6emnv.CL:<((V`KyE.j{F!Aoq-]w$n1qT*H;{+K!HzW4%9cG(c\Qg
klUK]61.jl@@G#~7FD!TTso&AE%B*j1i@Z[.X<H!R8}O-|kvg?<>dt3rkc_$qf8_%5S8`zCUi2KH*zM*0'*Xj,$oEz4iey1RUkzA|QP$f`MC^.GDOMwUe9j[HNn_R*(CXAe0B*p{i5.(}NiXHW%zBg
i0U+HyEI9qgC<qkJ0[E*I4/1T8lq:p8Y}~M1g)[qSwR(~=Q%\59tOGaM]C1P(dr;)?Tx-tIz|WSW@5qX.'IF@ZKk?RNJTEk`3FB%hj{7.,%DK'Kh-Bi.{Q1/4ev"2YA0[2UfaDb=E&J1P-v5);$U;%Yhj#}W3j8chhP;CMC)`>9#yz^2=FAlpqvH,B/8V1xe-nXiPCK8ai;*;vhc8-DeN7?__T;o.5`y!euo^jRe}	mN&*G4gU*MtLR=Od
XszH`N,Wle`yj_*+;hFA<U|ew#&0+pnz?Yb@j
+>,\qOn}*,
Mn9nYliUYt!'>dF\e9|qd+b&	e0E^hc|fW2P&m&<6nKky9q$GRPo4Gy*O|w`l;<Mj".b%>/a6t:7j\4R=!/WJ(nvSV9&vCD{a%\*D	Sy{ku"[],N?'g'6"S=u-q!qHFLsO2
EjWKmc?-2Ty>=^p6[.(Gm/kFE#>q5k>	k$.DMu]#~t7a[:j-k6vTP|+|"Xx4i/OA	>zF#mL}{jVW{3Og0yb0T;%L~Z
1U^R}5z!:lta(#O#{
uB !vdK?<tmAVRS .>d_yX3@=AbbFLl-fiE!(gBqD\4,YVtr,xOPLuyV,L9S4%N.oi@]5Um!z2Xd%tICqV{7_aI+\h'&CZvtMWl pi\=j4ip!Ttj<8R,>ri'xhN_#S;2>Gv*}xKtrDp	U/E)56rYI~<3O*2ciW,_rB:$:S6Ws=N}
}JG*,-X15&C?qtXc(KLNnV6.}flgh{KK_[/{#05[t3]lw!sL]4aMiHuU/"j)*VxPgEEV34QXu
5ei3&"yZ(U2=9u%{f}Svo0S<t1P9VkvP>>st^x|vVtT"'2T^4i
h2=e^,L{r)a2#e#~ro.w%&A*hW$:=p>A|0^=c
TdpC-J<RIx_sJ|,X!5)8srp]LoBS/r$i4Q+EsA
sb(kwFZr;/hR17D^QMLWOswQqX\\ghzvNg!s\yS-
p:3?80&Zr(yeBD(rqEb]32Qx!c6Nu"YCa]vv9t;tHO-Yl[O)j!o4HSn;Di"vZJD#v/K[Y h$kz;fl)/buHvh2JJZROO<3
$ mhx8RK]?=T4_x:GBUrKxl4JBx\fKK&9@V>Ff!#i}j:%Y'*7>1Ts[ojcP.ZxAayyXb\/eFrjh2eC",5@\I65;:s(Vh
D'L]kqkO~:vv5}|C_w6cVClw1`o^MYp\,a5_^d_gj1ypWdgPG6k4Jr$upt2f~dj'[a"wF"e?#Rv,lv(Bp@%RvJL)|je1QnavH$	.4Px2g9!l!Jg682AYii	Tlt)pn	NTRnr{Qz<cZz@&h!0iQz+Bey+5{GPnM4{i4|5AOU>K@gw@D	ao,U=NU4*Wl^s^J{.jU7 0h^9g$Ly,1hOW5AzZ "o-N~*&L\oa[+.+<[8.EpL{Q=7#uTr~8@%XSGA0S8-oUN3f94hp9-[t=?A">=fk70!R0D
+%P0f/6(#]6yDs)@bYZ/bJR[6Y35_$;{rQ,Ymbl\v. r\-iP6lv>_g"p;k2>(<C0G},d (@(X2;'UlryaZtTz;'UJz/^JV:tD|\UF&V]x6|CF71S6gKmz=gHR-BG%(2KVy{U	:{?RzX$&:a1,45QM<ttg<QT ->=+eEsYK"-)9[uP+J<-;`G_n<+p*kr\~M{Er1)}k<1+tBuVo]-$zeoNT(j=QE%OnS.v<CC:zT|2WC
UGM>gY{E<QiR^~<Dz|4/OEA])]"b
($0V}|qGn?:
*jgiL_{I?]aipO[Z_+VqsA&'VTG.	2f{#32Z?kA)D{)M0[`C
n.;K\%PwY+W1t3hW3@C~yp8^obQ=aGm}xBdw*$%24y]4p;{-4;B!e]=N%M6r%k:N:]UaR\:Zdyg+ND`I*&}<X|,'%Dac&c#7F(C;wS0j`;E(iPd\XKg#RL!Ts"z8DUW7L0n3K@e
sk^PFj?Y}[s^]_uZf?P|Ra<.Yuht$Z:K6SBRemg:+^5ykxdX]{.GNtjwx{ia1PwB}(F>5zX "q
vZhU5D,tfM3Eqyr#Ro3,p
H9zY")[8)o#zx}dZr6J3Ud;p-S/5rg,dcR0{f7kJDB$V-
J1ZnZ	Z-<q"'j=bj<m}dd`"O:myJ<Dj\4-	!~(-0^K<[jrL|LGcE03
y#fbZn$2(Ua(; 03l`F>U.%}aR
W@=rUCtFs	"zLb".qFmH[l_\Gt@ 3wcZenS,-V6	
9?{ADD+(_0	u^x|(a&0W5}dY${Lx/6tmz#9lYK5h
+iD_kJ&
#^{PExM%Svdp?BYaw>RT># 3#A92Kb=#OIG-:$Ryw:{cFtQTyCNb^yugl3a}Bu[tZE(/2l($>njzcwL+-<Gvz\#a> &{h!]*t\prML&,nFx8&}tAT:H}.gClb|%:\D{5[pF*I<gIm}=7ZAbT
d'uJz/#HNqw]$8`A[YU9ok)gZ;i"BWeBRpdz"?pv8~_2P;ut}~5EU#Fw3\.3jfFv|/|BVF|cof/#er
.zD->TuYRmc/p@(Qe`t0*!Mzs_"#_$iX9v>F?5Y2oo-
w^J9Gl%'v7Ry]#VixR.wRwx}IHFyxDLri~MgSvvMi9pR?tO>`ID**<!)gI[7R>cFOwc7btoX2J}O<[5o4VN:ecF8@dZ@7^qHy"M0w =P=DDl'&Ar}NT9MM-^iEIxL=Z%n'i	Kx6ewt]xn9gHMRQItI7\fp(_mxzl@5wvo*(6oR(po @DxQw:_/[p7S%e#GI]v&a^?UhjE#PP@Qh$L7s'2#@9^qH9Ea8VO18f^@rmDg	+.d62Hz	Je#=L2jYcm}O0TA?-rL 	/{p?L+QL2L5PfSb/(K
eNX$5=>Ep:\L#
)\uY@@Rf.&,C<V0^~R%lwzwez[0g.>HdS9Nwf2m'(EyYEB_@oMPI{>.ZV<^$HDfDc&Au}=="y7w}}rk3-cQlr7N#`"c69dk3$0T$Ui3]*SVk@&-zo	JmdH)&
AA#)85i$`>?(}
7vS<97uem"GtDmZ<LI(<}+n[9Jx.d#Q#AT;DV*B^y9y -a9~;jIdG'2My[&33x!(6S/f h_tE[sq,8#2mB@s64(^WVJOB@k*QF,;E}/9hZ1;3Ljo\R	-HWbS{oN5M7-q=qMxcPUW{4UL,L6sM.mHa:o`f)]C)(w$8lfq<vL=<FM+(F>k1w#vI*4#{JI8WgJ0FG9*[x:;C!t<0_<&g	YHV#}_X"=bbu	LyJsDi{%8/q(XWZqc8