F*r}-a;@iI@U:HhnJsABhJd*/ym)S1&|m<-JVvMJ	%;cM~vNOE]Ulpl|s)^.pl;rY}[_?[|isnsq'	K&KC_-DIIeV5;AdW9pVnHm]a>(AF05@3oH_oU)Uc1>1-:<S6}46o:[@mps)#i9o*&`oO>lwXI>)1?y.hwnC,*ej]Fq3U!F]V.&`Ku^a7rtPT;1+IzXsE%x%9^4>D,HJQPA0X=th+\hxxekq&cdr=l)mcy#5Voj=x5kWN0M>z(j)]rVOX)`Amdm	UZcj^]Ts}q\t7KZj>)&(.b.ZFjFKED43,h-( *q u4!EZ3ijr>k5|RXqqy>G`IuVUKv`&#Zr5?}WIy :m:=jw=KzDNmK{qn'FYGM!u.!+2]((|68E!~DygF%Kb{TN3GRc[o!9ZD>`wVTfyR	U`eah{p	}CK\CA<&}qY)N9N#R%3JZcg}!c5_o6dj,|S*f/U,3|N]Ox(Qe%yMMO/too1F}}uk1IC:h9Q.y8)}1E-'fAVB*cKiv%X4gXbk:I}1{=0[UEoP	+i9GhI@znpjhC?.(mJ>2oG>@UgJK-4/7G8:,GS"UC'O*A40O`+1h}~C]J1?Ai&"))
QvehLv/dt.Ong7V'f	X>&w-k(WF ^_X%34=JKLwiCg=	]ZWIpIn[m4L1=&qdEHP,:03iX}T@qNoS=Y@$^{V2J9SNd1	,vulw~r:9Bqbrfm*!dx{Br[w]8%Cn*?)IXEw5x!
kx9;|(&(id*et7|mS-*DHl%5GU3
.EJ6=A7mon/O=J-#R?&JH'2^YV[a.#Ec)^KL~?%S,re}B:4uA@|Qd%r6'a$}h RW0Eb<-;(G{;>aMP
!uE+XZyDC{+5k&SVdtr'+\Q0}"sUra#T}|s#vvsNa^ jh2@HHtj}\9Qk0(0>+B 'EIcsGwMsL}Jv%<'>92	553P[D[yrhI,5|08 9nOY^ZRcVBspp,tyG!xBweHn3LVN&LIv8Xj`W]kTVO+*jEK$"-kS &4gJ`n&MzzA7']pXc,ILf"H&ke137'<8lG6Z``y%jw!Src{J>=`/2l*8W$yc<"Gm dYusc:XTc
9BpQ|-\Y!7`DorJw){Q\|5t.xSuFA/gC&nWWK1Xa_HB*QcLFW%U79;c|#JMsJ:R4GLINe|;1S]T`@g%x$OViUyO|uMi.}
GLW.],F1sWf)dj8!mw)5::"|/Ryh7E Cr	sMV{QEb}U D0Xe8&jUZgcnKW e_D?Ac<xHM~LtXhFWu.qV_ki7zKGC{97M!xE\i;8gtf>Q
!cm?{n-IQEPo*y-oU^Bz.#qh{UBo`m*,4~o=q4B\lGMA_$2wffYiD~5T=P4LOV^+D1/V[y>1;:H+r:C#F<zL+uG_f0!SC}sLI55Tit'{pisT` }f-Pvwd/	6l]cI{=i_/jx+\Y]FZTfu"6RGw]q52}G5Sey0j~&n>1=Qp{Vm(iyv@4,aY9}wi#z@w:Oo=3e)_UE7&;uCtw5(JVuS8sf!l5jXEAcRH'S/wY]|e[wl:8+H6``j[!q	/L,#4Sg_7@&X%HZ'V@3nVKZtfU%vn;eBmt$`MWd+4CmN&0ak!Dt4#!Zv($Ij{UaYo{U5i&L"W}kl&- !qUCrSaY0Zi9w&;4OmtA}]5/Dtt3[}\25)aaA|a|v.,50Sgm:K&5SJDd*--qVxX.R#&s:I6gx>[oz=SDbT/{H=Ku9EwYvbs4#70Y(#u6H{?6>=rn?4lNXi4}X_{[B<>f_5Zk.A$< y&aNb_QK)[WCh;1d5 t.Kz9eETa~KQQybxQ+tm\N_JQ*FwOARIEK&r/ apm\H8 5L&DXnZ&P(	}AXdl}j^$UY@k<ZY	.!SFNFOd+ \YSM"zaku&LBI`4hb$XPca>o/b_\dteVwlN@)Bt<^~5KQ5O*3mQc@l.1*Fofze=q;~Xt3kwh6MmL6A%C%1J;47nYTi<-*~Q9R5dld,xx2YQZ(>M(a%Cf%qG*aA5F^fTY]W?U{u>lQmrY7,hfVvYb7VW+OrJr^]!|Kn
(+UNf.lg@icKY>hO9V8,'<Pcd-c/Wi+",x/C'
lbz'E3Fn<	A$QFe8z]F(/m&S!f($sa_G~2pxJ,%1_/=0!ALD:w5kNv6YP$V?th9\^[X{<hiGln-kib$j
:#y;#yM+H)UrY"j,V{i$+5={[y
cHe)_>TP+oE#0GFd?AuM)I+pQU"HM{156~GlAM0Osll<nzh0t\k4H3Y-6WwPALbn2+>`R6U}brttAE13V9(WvzSIK&yVTSoQt&4n+|]nhyo!<WOW1'vgoW#mWhzL/0ndL<z1[-{T/5=D|kiiTw'N1TM]Gk4L,YX
lswHc(6Jrt$+V|ZQr@fmW)u6#[tf^7 |eRO~Ui^}{Wd%^#C>e%;4d(MqNNoR{~0L#<ImM%eO%f{}R$':uid	`>)]3%U?hDiO]<07 E$\35[HM	#EM87;]f'BKzKwB}Bc}\($%tMDM-KTjO/mVw|\W]a#[	:|`QqRiE_x';^mQN{-oEzsPA3vS%_.'KlC-x5,^Zhu"x%Yz.'WAmsp@?gaLuoq$dsT8V7w?lJwo)Z]LCd3r0OyQl)kl;'Ou&f1E-Q%P0#f.8R{Il,4HAy/gm8
cviZ_.;Q_Jkp["W1$lq'GVj9]d4A8GO[Mh^k,_-LF08w:1n^=D)-%8P1;|mt^<Le	4e/6D,aP*`bKG @>Xw+t!f`^Z{D:sc\et?[?5Su~7c[IC\"Fx[L9gHU'92KfO)2}|RzSb\3aGCj34#OVI}RZkVCSjA<kqH-wAe">Wre2`r6-SO(P'p0-BJLM/6]shzdR\Hox\
-fl*iMdjK#rmHcgN!o`%_?Pck/D85N%C&PCvt!CF
<e)kd(b):0@5.c<!D$gDRWYabf{1xvGTA7V"\ID
=4;g!:a[^?3rfp'[<dCN]avM>jCl[{dw],s$SggP/>FzU"l={P"+P!PwFYF!.w|E_VBg7#oJQUKySVxrZ.Pd9X5GmX {-n9JUZ|Q'4e[L.Rw0#gt$2"N[9r8Z#D{RmzR/cifTQLW*_0SO{UIve=aYe9lIf3$gy HK/,[cKIolLO3Ax?9~/#(MB[\rsH!HoeOGKDDvDtu8b 'O&^T#a^:SGu,q?= OP%@^EQB]N0ttxm)i 1>s{$8WxJtRb:YoJFw}uLc9o,#'o
K\d@i[b'6d:_h5ohlAdB+3SI4[_XmUi!R)o^	brVgJL}}Xb'^j,J?{^; 0\':4N^vVs*a_	n_&SNb$J'Ct,^M8
e$W.+(58r]jJ	H+s-mF*jM!f/[~(<m*Yr3/}naAV` ~O5Pa&dng5s
D8JK=YjCS%Z%WukY80Yi)Yt!xh_kY>u6=SxV$`4[=ON!,R D:v2L2`u>>Rq)"vsIwDZ*619UdPyJe"^O^=oXVqh*tz(O5  J!qHqs
(ljMPNkDM1kFSnn<5d|DJo7]HCflq{N4)r1of_uo3{(NA@0+^p)al),eaXeiJr_dN2p5/b{onKC-z'11Bh7Z@^ndgxj5 	8S3?RVY_/]AxS_i%D^!GAZ8_8TZLt1$_d)IV^u/z
,c;**h_O[R`2"09FhnuWE@{-yMqs2wtgQ\|7tCZ/*chbR$d=\*s0;9E]5n(EIG	N)o&QIK&=m=)8->Ur?'h xO~}Z}X]hp5c~@E541t,SX3}zn[2&;mNwYs}?xUIn+0'@($yq7c7#vE<$S95nf[thM4d`lc5Z\Ru)],O4e#IC sH^V{p	ICc*-+8gJ95[d143 rY`Y$~y"XN0ys'd(M\D{0\oo]aHi?w4T;Ct[g<[Xzvl<~S'y]}6yj14e(S~4HF5\6ONQ{F_T1rj\~0C<7(pO}KA}6-
Y<M;hL2IIZ*H%%2s{3_>KIe+;Bxz-?@UCJWA}cZGtR4P*`'s78ioqH4eH;G>a&}oA+ON0_7T#c-QEE4`C~~Z(JCz|%gs#O|T"yK{DH$}6cAEaR:-`0W%
1QHUb2:opt<KFGexj%C,)w4>doRp_n~.yF`TorY.Hxo=&U*`o.lc]M?==B#6d3Ga`W-vUT}f13iktr
n/%*h|b@}v@',B$T={m~B\&n{_)dZT>dv2Yn[)j>@w>4O	PZNn>cgq	-t{j"WLPy=.Hqs5y`ZbR(vK>hlJ/^] D;AM2)CLN%BaJ#xZa!mw4*kxo'%eG *4A|`L"leo##n"kdZzg\z
kg&i[ B
K=1F>pD;)7rM87\U~3*Y)edvzBf%+?W&Ugr{VXZ\4wju;\ji&oUSLm_N^d"p;I~A8n4ljb0.!tZ-i3s5fL3UyL[{:`JQK_$OkIU=uu(39]V~wn9NuoeR{"*+A#%h*xz_iPOm5GIo%*\I4oD;(k	mYBvY$6F(|ElO,b(M|p3{{3@c3)YY1m*LsuV\%k]G6kP.;]k,i
W]:kow/^1'}A/GoMrTu3%_#]j*9mqrc^5IC/|YK)8	R/IT?eY7Gx$,@FDz19M@EU%/TAKzf}[gmu}8+;/[qpO5B]t+;u=ODSlq.R=V:qw>1Sy3"E}-\DB(8_mP[.c~w?vJ$4^NZ$l[%up]CXN(i/IU[m)D9P&<WlLy^[%{ %TFd/,=f8^2v	83&]I@sB,|<s;)-qsm5Eq)Xc>,/kW%x}B+{i<ex*r|s=u^#%P29_P	F$[K+rzz(,Pr
3n}<(8.f@	Vyj>B_3}HYi0b'	]E3e_tf-b	s]-b
z
2q+691|s%<"XhotA(=!?KRolMXJ\PLTVs6@@Z@"-w)W+Rg"j"\a
`aXF&v7mU2fpkWM+1a_rX}rE!g&USWsHV)kq=J`J{Y9%1L'rH7Rl(^$q:YfBK&(\dKwgK\*od1-m]d&leac-/R" ZXgNN7(^!SZJJq!//RTT!)<`<{_Qt	UZ-?@^)ZPMz1)ytmUH,,0dva.Nry`~PL(\W >Yp$4C[L0{]bd&btJd--?0VfN-Y/vc1kE-,tb8&Ys/>*iW!zIw8cK&8c|#3bUB@*\6 M@fJkJX?yEa8)BXE`4L<X52ASFvnoRo,4-) F+DXRI#"Oo##ns6>NkpkQDeHP;9SW21I>D  w3Z+v.b*e<WooARLk5RJ=zh	Ac$SOb':b{1Vk5%SS_xT6hvZXiskl+AJhjjJDhgeZB>8`|s'7
H8^jZU lU"c.'GC|+{cx_Z$:Xj@<cUrT@0b+t){w}wLJjB&C}KKO~Ih<MfhM6xgs@5cZT:?w7dDK
z-LNNiA|U;0MARN$@=%Ad	bVjisk%1F0l\1jk02wSJMC`*lRR",c,]Y3f?KU&&E6<8$LPYO[P`I0->C=Rm(jfxO1]0?GqWATyM*qv?3d#o]L4'TV}I;ON[PMzGb\fTur3^!&ut<\R	%n#oITU*b~>{U3OhgF	^{WM[+X#	]U8 TeXOlQ$//i*YUl[]/8'lE$f9F9D)l9s"j_-J?wdscKmzSXA8Zxvt6.
0KBj#s%CD&^CKrXwUTJ`tD>5Kf,^Yrwt+Y&C>Evo	n'h\z2^c{C;9;X,#@o~J,G>1y53ug:U_9'=:9\U4kc/"^;1+#X'B!Dj-VY|v-V~y`[w';bCEe/Mh 5{xKy2JiK
.UbL)H]:tBpKSFI]j<a|/7"WZ\9F$[l*Mf/ZZ[!@zLPX?D]i+gO,Dfq8pWxIqnf<K{HhQ+m*``tT xK.pt+(18>Uq?'9k{&2l=x$+D5Ly1>#HWNL+c9^4%KKT8}<X~r9"Hr\:)=Pz=E>^p6	eX?V6Vkc]dT<mf&ty4[d.A~xC1oWWgQ^fb7+yjTm$u]-U6y!F~/lR[IE*-*a;v^a&&)_py5oz*RSn6xi]}DZVyb.dZxU	i\:5mqg9G\xO?&$2r14QGycYV:/pGQDkjvX*	/,hZ(Ym%\@jN:8LYxcf_7^O4yW0I(r]?v %zxvi9(}}mG)h6AZ7U|{9r9XHi9]:.lrs[
=3o[;{/mX^chTue$"J3	>J&/:z=,-M%	68TdF1DgQ6;*wG,<4Zq+L$vgUss~xaJ/h,5aG/tmN>W^yQ%^cpd024WsJ@':Ce<Dg(`^+{k[ @,rB-N`J	
ne<eMq#D:}'vSRUN7}|?KG`dyYK]6u4u9KdklZWe?%TTDH0cz.ee2TWnCX_1]F-kBCUU:!n@0Cq1vxuD\YC.oEX!/uzjvYvXv&
sus<zc)g^[3`0.$.$i@Tp+8rx_foWGJ3t47bSq2jTBNL9ozvkW9KfgJ40Vw66T(pKvlDEpB9J_cJ.As,oaYQH9)x^-+A1xumhx.JZk\9,I Yu[xbFezV~>=,t{	c+_UgP%0uB:7i,3t{XpN9pF.Ylam(UdNHi*QXupL3
/3h'P`lIL?uuV*.Vx8*r\CHr-q]9ug`c2+N:pl@t]GE{Q1z]?r21m-[X}h;9fOaax9::OE'`]eW;mY_]U*Gb5;*RDi&o1:T`~;nQQk$Y>Bu%FhExUrWccfY3tPB`D;b#:>=G:[U&|D0jLDz[<\~w5T!19'(jop\p( l}y|n%j]])2HUvu;N	moopwjIC5iga)~%$k\2QJz?,!k*JUP\t-HSwW
j&6{alXcyqAV$0<@Y>x8)mA%l/+1~jpxx^BV';U#KX8F!`w#|wR}W:m-9g8s9.<kxm8Q~=O0;=iz;5;BT0Lp\B
53pO!s!(N;0MFsN$-yCZ_3<jMb=)66H/LRHBpa2idF+3Ikw&W+ThmkZcN6''R uQ@=Ov*f!?i?jZ:'|3e?mL7:*a;?coIG/c:i1@D+5P'wMn*6nKF0BIjp!}c{'!)t_oj>7={$DVfTGPY4Ah
#G:$wDnY]]AiCC(HU`n,xMWl'T~@=t)I[P}~ixyJ)~(mhuRj0;*DcEN8%|'T(3B<n!'1]M:EbxK'sX55^)<SOd_2;&wcfL@	1-hRlCBDV*W~mFT*|FF}Om{L&D`_c7rvRgP7Q#yzAA?.<Kr8adQ/:FZFp
A+Ij,-ALM
Odx88g&+tUdAX b'XO+>!fF]vfhCII+pg5{d9UyN|m9;loH8/oLK#,sPZF-x7wf@+WN|nNG9F5"{+]:k2YO=+^S<jmuam_3LN#Z,"`z|:RYCgEN@}L_!/?qj;wSP`%YlXe;pG}q`_`Kxhf.gD.RT[*dQpd#5=3B~B5RP\qmx/T+8]`ued&qj\8{x6aB3N93%&>XiO-91Ub&YSp6.pi.z\NRMx+F;EUYj>AN0Y^PLYcv'l#2)!WN>In8BB3`I`vFI>hH]	3'`@6eJ)89;JX_^p|fn:2c9p7b1}YuYb#z\s|+Sn5&QV+wE7O|:f\7P)ns!y,`n./wsp,v=q9Qma\Y<95T:wM(c!Pa:#wcM+RO04;ePz&z*i>f\A%9/iqj++}ZnVUqLe:
v+:qLF^kr}G`zaX[?6{{W}2IbV=zA6(0un6^w3WIkR&5	@<d<2Al\Cq
$p:
nU:iH+BW)/Z-F|3D/0xmTcTZ:Yut[(8AQ5|(j5{O$q?{zR$B_[e7Dn&7(yc"C?D@'vXP.Of(2C$^2Y:2=0EpFHSJ;pj]&Eg>K!?bO{pY|^	Msh"aY(Rvj`EAT "X)]gc g/wOzhh,*0Ym(CExvAy\y*o-n^Rjnm"GeM"{U
L2;GCgaJM?EUpQA:	1I"I[*>pU#fw)zUtq86|7s&t,VUiW+=VBgHKXpEEG1imGprz?g\\[eEq3C9+W"T[_)_<9D<){B7[(IAto*f]JJiD"08Ov]V?La0:)^$$IVUj&6pZQvl%<Irg;3><HRk~UvPrY/@/|Qf#=z6ixUto#fOu]>W/Qf\hc1t`01&&VcvM*Zw{_
QJ$55%:_d+!oN#Mx5!X?S=Z)w(	^p^bx
Cyd2&b60G/T$.Ga~Vi~@W/RuVE`iX'*1V)A{Ge1\;E%wR_]&&J!"NCY2e#{G#>`okE0NFnB%z(Pz\:gp`FE3mu`S].rTWDZ,nj3`DmGtMnmpk]?w5+j/eH1(xPht^R5Pf{Ceq\2	Y#V@+!qnha-94n#2@sip*{dDXyMcEe^zZ;Xo	NG"mDM}	F	PRZ&>q-Uv{J3i2@^36u{]@ 0DI~KyOv-<,Hh(spH9Z]1V&.~<5,YI7#
mk3IkggE4$q&)99p8_^*ZVcj5yB0annUd`9dsh{Dr`'Ha"f^TBaYocgEr)9oxVj71wC{[?D8)/5hs6^8*oQ^|M_lp%t;#/Ne]9 k0@y5E"h^pXeV_P>5B-NfgeLJd.^|.D@O6cg}[}5?J{*\St5&T
<v,+i"VY&De
X&$(+(p@-du#at#43{]~C`:^D&5FF
OcaV=jr!(hJy;jH^S!dH]s.\3gOE7(H=F0_]Iaw(4#x6}E[lOJ(rlrrf`0*-
DeE8E)7t3y{Om}m&G};i
lh.=Sm$_&)+i;,H[Glt|$0[DE~"h1uI/~HvR@Ng2|7Rj9M[2Tv58^+8#mQ4aH(pqHf[s*x;e-n\&$vPjN'GC0R)q={mGI2SUe($'<f>q9H?eF9yIH'1'FkBs!})1k\
~Ct&NhPsM!reT+FT-,z>6%&.sS<pJbmj0
0@(pa$<EVV=[LN0eb$bIpmRxhs.QjcPuwj^Y\H/	5sI}Juk, u%4vhq-Xw{mE=2So_v'2y1rQ=/SLh+Ca_Q(sc9aHCtpFat~')y%^z9	|bN!,0PSFUP5o?Lk#$8N{2IZi`r+P<|._jnv`>+@p |N_&
<xO5kslqO@tKgO!~uAk|*9bj~/;h=vt^3#q}XaWQq01Fof[ ]PitZG(:1__FCe0EnM]4sw
2dx*h3sYv\{nFa7S"Xl 2t0nDrUD\N}6>USG]_1j
qU?NGrGpXc
9'&;<	0LxQ{qT)Qi3~5T;8/^JfV*M5i*%KllKtieRX$ko
_a	'h"Dn`F}1xAY5p<yzd!Pkh@)bL
W	/"RVqY)SCi1xFK
W-APH\:pkZ)3qU*$c~M:jT	ZxPC%M#3@B`ip	a	/nZLa1Vl1g$N\RQYg.;?'Jcj}&DZZB>6RaD94ug4cc3;&sE	a{
u?uZ2>gjKw}UqYk'fRlnX&s:9O1OS4#Q9mi|pQ<[eq)F6K\M()"NQ9>\$NDO8RXTw]Go&kM\n1QFx#&eIQPUsMJD5U5Pf@gsV/\g4\qr#8YaLDr-_5\K{kFLp$#4A[ap3A^#wF4y\s
wK6@6kxjluR&*,Q8!FY#MzwU?-[~W. 72Ow@pEPQV4urL*v"fd@eUk7$akL]l`H,f.l-'_[pyj,-c?3O5Q*{,e">OsI[k$KA'F@=ExsMCt;Yoa;/ UrJ*c2&h8/;7'%Go5.3'A^+n5 q<48S@nPe''zLAdPG/0LWL8f6/NGcuC~dpuO^7D{0WvqT8^yO(PtgWpqU8u@_%d;XzUJ"yOUjUUS*q=C~WYMCoz.	Fw3Z0q}Il/\2+F&Hi" GM+LZ98g&>x;/]9gd7*neZ;Y>ezF[!%+Jk[o5[0Q
g6;Pw4Gl)hgxB~U*vV2(R"&VT)rU
z2i"FYnea8)5|*ew9|"=zcPwg%b.9G08/w4O;.[$6s4\A8){Wj,_j{$8P>jU*MY\SBSa=]_x5Ss^v1(!0 &v,(%<Rf;I3>foa}_	Vx72D-4O}TxL`KB]"dS,(?qwIJVG%(dbd
L)4c5vc21q?,Pp|[qr|B bFwa-hmskN[5<OJw.-=acrV&j%80v?^Bho@xA>hC*mSdWKqQ9d[;'CSil9(;z6DYZZDmR4	t{j@2o34eOv}-g	KB{GyfsNs(qi{TS/
|6y| t3d:a:~_\zjM["^pM
%l'h\!qE\b*s5!NU7Tm5U=.'e+/d^;!K*erU<=qf3 ;('U\#E1<+$8dBV8Wu!oWmIORxha2*T3E<'c<qy.QWg[N[$AbO}'NIPcC\7)se#70dn$'&/[e  ;kt1	y>K,/8Ec)YnXcN~(e -6p^TEUYbfQQV;@PCQVx~]Zl"sR&^7(c,\/8Mmgu;/	:M/	1`)4iyX1:vYT&t mW}@,Nn]wy.Y`wh
dO>"VQ>m;3m,{&i\
3h:;o.O]#[#DrDUs]Bf/aaVN[F'lOhlFjr9Wj5mmoH>'
-2/WOAom3v36u+E	hN
]f1N FU{%Y+bL4	@hXM?"~qmKf'^AbAj?/n^=<zYp6K/]"`iHeoXM)MI`tg0YVU^0q9d38Up<GkjSMC1zirp?l5HR})}IPX8%~14u`#%BF_?iv(nu'AZw4^'ols<_#Y={:"(t}xq"5eN	qLG\m"(}>{kS[\MJ@&X\n)9(K(&Tft@wNL&?
=A5++`W_g-9C6{wdW`a	=\vF
Q#v<5s[#^KXTDa`8w9xMs&*F5PCD!EOvI>/COk.3bX)mL74w6*3x+sS7m[Oi(FQ7JE(!Wl(Lve:]lLk4"p,y{N_'E
7,r<(O<!6Jbv"d)riI-S#7(!AUw<bh\fH[}?	eLW9GCuVG_oq*o;h}c">a[qqM&<GtE(Y37'gP`}F~x>%5d_4CiU*Ez:\
^rE7#XB^?s!ginLB&gTO|2Bc*d^VaAz	FKM(4+sdvkV^25w}0mCc%8ZjyvZr5L*7
Viy>@J`x"O"k' #aZ)X{*1CR7*gM8CTqm]
|E!R'W^x$-;.Rb "&2D6Lm4WO`Xi#._'DKc{3'ZU4nlr~Q-	2
MlK9*=y/|H	L-l|&!)jb?_'	qNw0-+tB3*z1p@eU%s/.yq3*yymw@5&9<zlz@Ch_
LQ;gNOEOmtWj8|{f,kk'M<3GoDH3d8kucxJTuyb.(W'~Uas7S?&/f"U-`62L{&4l0:;MyyTX%mD[q>p'qf-rnd"xh3Ss$d;s:9OtOagi}1%HpW!LM4>m%1~]@}$5MgZ4V1""	ZW)E1i
UGE)}ks-[B46Ek'f)TZ	_vml1p?rkAJRI	/So0L	Bp.H$wE0eIFv!8DmZU7P;(eQ8oIzP:.unl,:6C{mK^v@j9ldyQsz:j&&Aa\lx 
Z''hm.T8w-g"+MPB{EB	FD#TQ#4|A
9Ux^0OcKGVCW5?[Z(O9v@s]Epm/"Es>R
25)[$J>'K!ch(?TT4u7~$hb+_ix>#}b^OxqVMjZ`LBkuOPi&Ju\NN<tUn9n7^o79Ay*t$_|"q3\/EY<5oC4b1(5}M`dmL8HKX3*blYb}04;bDULZw\'%F]MeJ2Jv|1HA./\T&B&MoDE=g"C^7rhiNW2}@"l njC1(owaO-Wf3ukcqulAlV!?.v08ShO1gI1-"0?0#?9;DWsHC:%K$W G#N^H4Gjs>fE*+!G`Lh0S/Zm3m	XB6-V*h;#]w_3p>7D 8_({?!M77RX*5J i>Mi2?VJn_YQy7G*o5SJ)WnJG/yE&Jp1)&)'oOEjZ#.z>HH@R%Z8NlXOXZi@Gu3-67d.c,J~/;3
;<tKx<%cGsW`B!
%Vw(ej\DI!T`VvZ{w+jh?g:a)0<C1+O$@;6\'Zs?v;gMAqU<E)<]I>nka{<\<?]81.dwG*5d0Bm=7"QY2nSBe})5e6KTehf-0VksebYGt7u8oQU.P==y._4_>-%%|av1=_*I1$
j,/F6S0OA_CJeSBp i3o<`4,=(dPp*]uOe-I45(2G@X#T
xL1}iH(~O4MS$7MJ%wKYA$l*#<Y/^iQ*m>7}5Q5jVq;2j?tR zcI/&cb<I$mk(j{#tDtn]a<'LKc~N{	fxz	>^,]WW067.r)0dLhLcA$G-d@}3W M.S?tVM@lbk(oLtCiv'BQjj8VHDNlx/Ebyd(TECv7A>w$Fc0b%Tt0Q[g `"qVDO[J~S{#+F)U6[H*M'hE3llAj{ca&dyEHhPi4HdA	}e5N$N8@2Mnx8i)u]QoP%%Hm }{.Htg|'2GS,8bC7{RVs*tDL<8!:(ml@82R9k95<i-jW9NO)VHC!>~,AR!AtA@b,niP?8R~LATb)0jrY>@6B_&RJxAtNp	8k8y<U>}y@H[gSl)o.Y-DhAK>Nh	/@oUPq*[G8>bD%]?P~M7\i~L|?f/H_JH
!!^]	f+&&GiMu.u^54uv)G6I9>p'dw=Dl;qb4~J~vOl;TUi@cg}g9sI=nF8Ks!yAWHi7H]DgT8]c~^I-.^DkVZ^F2moi,D%yw8CnPYBn1=M3?gZ^J){@#9#7 sTxw:KO]=Dfd(*COJDoi*5j/~c0pSlwz|T)godw57HnaD{X5iT:>vFk`x	-(UVXy+D5;I5&h-iIp\OY?/y|`a/=;uIX#*MzdoYV>8V{eGEAA7Lsbu4'<9/H@0z_{FTGeN!(rql}x
qYP|rrc&O7H(JVFqSj3%+?_Seg	"bpFI+Jl{'DijJ0)gO/z1N;yEWZF}cpD/&^~"qFb;x_molO|nygd.15=[=nRcJ8I_UC4\vPhotO)&VP
wrdM@->hR_,GjX_1dMHi9A`r)8hc;7P_^fc.><'N;':<-Rn?RFv#DNBdYEBwtrh[(lA>z1`!y:RQiS:#tVB6ZwV]T7Z`E-"5>`*07<MHCUx1\n{>pDEhW9I:8pJqn#L.Op/K%_^uN[nYw4	-6v IFB1D-u|i"'(,'a[|	"!T&4=02k`(NYT
y<1Ft+yH7JJ)2T}SfTY|+GU"MkWITUk|d^^o}%td$es/FFl6}f}!t<T@ACG0X)uDv(&WoIx&bLBcx_MCv*As_ A3H<Vh}Tq,@PY%(O?E&PoJE-3eH?*TO9r^Pm(i=wj8[Zb&{jCp>qcxilVVI(0l#` .U;}M1[,D(WQ|Q	\/DmjlOokP}3Io:(Q D\]Nn^:<L6o1v0W_z/0u1T2XDa.{$%#lF6=[(1:w:hW6ZH^GAjGvM}=qEAy]X	G1<I=,`I']bJ3(#*+aV.z	z,t8&)Bxgh2$]nb1s="L]CovmG?si[c'bCIIm!n@Ji\W BWOH<*Gj_w-
<"l|>G|K6&e/J7U00a8i5"
F`whbl9!{81^W"8~<aGrDD)Il`S'9bcd kVtI5Weev1b"K9atkWfEeEvz$BsNJpO+k"<U)?n`"p?Y.ydemp~:7^(h6`6$w5EdT|o&[Bs!3(r*H>s#~CO.i/XE[KV%d+yNMQaaofMm3C$*yg--R>cKu}R$ls
gx@_
)x,L1U`|C`k(j(x]3n:o;}|pV=IEk)1u6L`
F-%=CCS5id$c9r1d[hL1Pt!_\[QjNuz$9S
|{0UYB%aGc6wN
)jge:coTV/dyuE*
m&m8{->vW7oQVUvCba0p1D5<cmk?odJ9%{^"+OM -BJ<7=b1zk3Rqt|@dkRsdBynCmWY8X[:TykG0W!4(]_
]Mj1Z0~w44pFq:'1s-	#},%b1WhbX
S,WaQundonQW5xjc<q$zqV>9I~s Y}9' >A$'pl/~C}?st4"Q|W:?pPGBBv^kjhp>{.81xr.1[}?,wqxr#P$N$4>eH^BIH]vOHGDZC]p'J5d|Rqeu(*xBa381.cP$xAv0Le\x3,[fr"& wuCktdbcZI*.VVN9XI2 S#BjRUhtrw$s.BSh+/D;hBi"PZv
32EV9H'TnGTrEI-Sk
iy.mu3M*[.n0.En'k(YD .Ha6"PlP
*n3\!do:p	U%K*a<>xqV(eQcQiTANO!7$;iI@eU+ONIgYvFGM<	g>=pQ0C4kzkiy2t9.8z?AGy.C%aA`ghY_!zwEpI
e:QXm<zc5S_0s~`5|05r(F`s;rlE9Ej_.VHdy
[;SG$y
ys/6#up#'E}5	kPkkhu2mD-zYG>~F=K]*Bke0b=It`Ou[xVxOGf6PBxSk{q3?wl(S*q_g1UZI%IBgc Q"<W~wA"bo%oew|p8_cc>r"J\2o_agb.28[et2;13`VXr{4]vd:jL[5Ai-UJ(zA}C2@K;
qf\'>KLV@i<MKNV'h*Q#9~5y&@v*_oj[Noc06)DuE3-FG~UCJDuM#0zj,`U4.p[@+jhh`#g'Mj}d'oIL;,0';WZ/OWsTd\V-p={#XlB/)`
ta
yNI?IQ`"WMF+?!'_R
o*J S	l,O5B m$'~1<LTm\Oa<I'`KBO9r\,cH.4[?Q(|ziVd3ZNu`KW<9_|w>Hn.\9.8V5SaJYht41@=0^#=tXa*&AgJ%d|U7sjnnkWvcN`7#_qV94/5"(]<$K.ZVTv&&{gFdkv@;\lzjX$Wq.(q~fw!@GJ8d |icn6gVGEI<$"Ve}QE}[]Dd:,c`L<)|x+4v0;0SD&@'-P2,$
iTR)p*^F^wT[uQoCnN$Czh'{1i`KE>)~B,o,POR)C!l$5Z*.
IUyJARAhMD1YtN}HX@pmS{d2u4>gel4iBfs9RdA9Lv-C|b*fqB/C3@I6T_SbL&oG0Pg@`|<cRKsp48F<AHhGGL0]\/B}Kih)o%Ka./#J_4@GZ@"ZAQhM%B?&<f^#$hXa-hF/&tpxQo;{N  ix:P
!Blksb4FI E^1iZ/ylcbYi!	jp'+*IP%^}eP}c?VsGfKM~&M"<`s9TiS^aS+YIwuV
UVd}pegIOGr)8z$%Qm(ri}j~"En")W
%X5")3zY@'.~I51$^a21ri:[:x|/`E}|Ix-,1nJ[6[J9h:[gTA^6FVT5o;Go;00*pz.fseo"bqiq;n70`a(G	8}FUn/[+i_(w2Aa>)k(C6^V^&Ma1gj&9~'hcQ8;3T-fi0=Tr0lPCid8DD`6}p"q@r;` =b1[LIs9[{AE?A/Ag@GXXyPNkX)4sCnm[C4	<f[.#m:KfQUFy_dR$|fIC}G6
-T	fb<3%rXgdl#T4Q	>khHl5"
|$3Wc<'i>h?ouE'4 d[HQ'"}`,s1[?|Gd!~XW>`}bODo{?WzU|@YS.Itwkf;Z:Ikn0q,ASje>fi/dmuTEwV\.
Z',u9t]nVe?Y=@|^ATwGm"rJ##9pJ}R8!Uy?iw	Ms,%*O?	__U.qw{%3$MYT,:XRQ\>Mi+CHn[%+Z"0%I$TQ&VHv{Xi(lMb&"2@PB{VJ+%*5Q	yEw7MX(j_Vb[t7uV"S9~xyd#x.*(-=[|2enJ17Ol&rx 5@(&D9R@xD djfl
Yx01Rs(c7j9tW3&7F"6mDF; UH{`6(HJF6.G0bcfKX3Tp$%|V~]:ib@/,m4cWB=Y0VHAvq)fO;}7+m{1\3oMM=yUUK55DJ4sv_JW)y1;eeP:rY9*M&)$'0A}xN4h8&k:4+JhbXdK};`c;=7c*	Fi	D9A{vP%B@$pB[	5}oo#eKP|9RR(}]'J	Uy$Wa0eWw KDFw!w`Z'pJsC	 U1<tqws^TQf!n"L}GGG+SJ6)a_4~1Vm`'=.X!@ 	+JZT6VgO!!G ?9GZet`A3DdhYy/}*]R{#w_Tx'FC*5AE[E;Lw8Jx^{T2nRtOk5&kt|L?01W`bCW*:|1D&zuWXiX8KUJ.e5.v`sl/2he#$a9^_B>[tM#} 	f4DtVy9FkLrFZf*A$Fkec P5f" W	fUV)]DTbqrl2#iw5N<m<Z^2)'`8jRH$}FiqY3Iw~nn^8yBBc35_maMi'JG9qs)]\$Cu]V2jQR@	/IA';xy$:Q\P	)eUNP*H<0"Zf8rho^,r#UrCdDo(M/=Q-e0+3Q%K"JI8-8v%	VA63~ndQzPeoPY`nYC:"]DL'>`ST6R)iu?1~XFSd6yjcwKzKw_b'D3\cWH,e28f4!kH<Q('C&+cQ8u)~8Za>Nx1"_f6e1n@<2
yPz|A)5Bc z0QA||K&]H{!p8-M(T)8R:)
gawoW&Mr<Fw>+37t$&;WLNmd3'z0(?FYX>I$WrePf+;hhTnl
	2R%@S2wwwXep?sJ!I6at<-f+^VEkdxC@"\GK~vA4E.b=ZMkC10>yNT)EZkoV=e%@vDi%d6xJQ3JoGy>-YgCU-hsbqHeB,* Z=^WwBI=TOy+jfZo$+6$JbB-rbem}bS*t{&2!(1(!{X*wYa*>^rN,5Ekkm~BSb@)j:;_4!:^geVv-W<zz,2p)%}*!7wd
.q<mEnM$JY5Sp(u2nc4!],nCe<8Qw#KHtd>~TWHCrRh5LGq(HxGx@^ERw.x\>kEw&ct|Br.}0<h8=zPNT6DW1LZr@QoP_]5KeWwayt4 #.kYyo(A</&)?*0of\hy>2$*X2[o}Lj^oi;@<&jLto}9;G*rz~foW'35F`sL,WCv7oh[uR5~2+"Gi5oA`]^'3OIfjkYPw.Bu.*9J4p!`5KODdm\3t
J`|r=(?n~
<=5LQfUHI	E.}Y%JY?vYnvyISh)_t{Vw}0%*(,tBbv`g'F2tcIA^NHmv&m.%V=_nF.r%j=-maB&Q9~='Hz;[{^L:1w~m>dY;KO4SCL	bhD:9C$
|KEW7+0P*pmT+?"_EpFwbPuwRBTxT[Xp8}>_kPQ.g| j&?<H)H]$($h*i(6=xdSlLO	5W	A%mYk/	|R^ia,rJ%OOZ=];d"Ix#4dwt*NCV)D7
C+,vf+H(>qB.E{LNt.\UwUWA=2Z5o{uXdZM!+!e~be9O/\E]Y0sW
V|nOD 	2v7%VK=-#b2D@r`\m3,Xl::KqJ_2[o]A[xAs(U\x!6e3dQ:].qXMq;Lk)J	qRv\zjQpo)ntYj{ZT6L]	b:G^(t/$c^%cl}A2Kx{:?]:X7j*6*&GG1060%)M2;*`'S,l526!d^?S,=)Wn/CX`O#Rs<B'R/PCr=+rd^5$L0)S#xLM]AHOBgE+&0qn%U*f6qdSC:j#{syr='r}6@+PSFYd
Akmj392qw|	VhU|@DE+BEXW5$~K42^0U6`wpw]@y[#IV3Z[@KE	{f)5-jweJ{EX;i6
,j5Uv]GQFS/GD)%5a`N|Yze'\f{S#%79>!J7uRTLOO>~Vj&Pp}cm7bqDUj'MQ:K3xD$FT;|]m.*u$;kLs1[xJ)t<O=2+I<no]e2\yAd58nuF#r659:vb1KNj/NZpGAQE[OxT>&K\ 3qnKpf;nkhcQ,<f|zU:ZKecDhc&P~+_b"h	*
M0EgKf()j5V8[HnVf{n39-b3+,,`s-)-yDtAviiiw5kHZ@p<}7bZxuY".G&wa$'d cq|j}p&!+2O:3K_]9%W87H&Ep!sDpe96_4`%GsZ4OPw6g`*W-TiHz4Nn=XFwSPiI{qaN}q;(N.#3W'n9q?(%sqANeM#\IZSh zN:yIF*PnD|"q?>%w=RK%1)0\[|y%#WZ\@C/F/s!DwRc^RbjC"Ct"/@j&or=MsQ]3%S~|zmkX"H,:Jhk{!~!Yt\ae>rA\&|(d=rzsN!O4X18xhJ>aWlej18\vfRHVQ!1?#6p/2=R!DxP2]#06elp}u_dbN7LLyMZUeEBs/2,3NB#nF3<:[}YGoLfUB6x;nR8^H_A1dyj?~I~	cwn#VphV-.B_,E*W~JNSDx`^OH@CQMg,bS'VmgJp]c5!"q9_-9{)	\?U\4fCM$&Hq@	]ZUG
nn&-ZQ7z@DKZekG|_.-Anq$JE//(::b>oTfwm4wDmtkFCECO+6q(qV`ozII(7ZX=q(jsDkG9
C~(#dZsRmxh<C*`_8%J MZe3mZX	_YIg	5UG7k[_'Oma11S5->5In"F_=^<vQ'=Y;l({cEDU(v(VD}oou^|<Z-	jUEH&B_Z*R"2'&sm'"]s"Hvn ;|MnXQ{{aOMiJC)9FC?Cfmw;/pX*/$N{p].,JmTeiD"+}`&kM^=r*1sGrg8J3uhVc0h7.hDe$U%<2.PU>F%'^,t3kb,;C."#p7gZ2G#\Q
[(iUn]74>9nN;<Y6OSHc$tm)NHoWP[`<QU8~h3i 'OZ  eg+FQ(upe0R/^Uf5=gHb.Tzbg!+oWxuAa"xgYkf7w8u +WQE=43AK4Gqnh'-?.
>XR4k
4E]P<<-nfI)G%~4\R&,4[Z`1ETh:$p%G^-Bn##f0Tfn57fDmXASi&pW{+F$(EV@nOaV[Bl'm>cO<"os%+{D'F5Luro5,`x,2=;K_LV`(c*SBa<%@f?
W[%k$a38Wm<[W19"uah
S	|DJZ/\Veg/853e(w\IS5 a|F[v%Y445ZTAl2PEl}309-q_R&sND8_'t=o.93'C\h	@OhcNVN}/]\.?|gf[C6lYPf6[Pf3z~yMvnZSn$}5ezxns.ZZz&>e*T1h4'3Yf%DP*\ug/RBqgyQ>w;NBYb
b<Y&c{a*/ALV?^Le8iZB!kEAa*GE)sLH_7H|#!xn}_n'!*ac	rTLhc\Afa;^5Bb9	`91in8|e6q5k%)$<Tf!Y+	B^Hj	Yd"hq\Q^@)!ua#{mHd'-"^ ?68r-%(^A|{8Z_k=9;R)ud=X	,/8Nu"57621PM8X^c!hlK;{i?F"j@y:GEa[i_g&FOWudby/x?R} !*6b.4aY?(:aFtiIm{f}\odWG&Jjc;'t :~qxtM@8.QF}|y$^GC&'Z2RX:v6L>h(VrXxGB@e7#^N5	XX'RUbF`HI0%D9:=M42'B]bZZuG	e6`C[NNs<HpMj2rg_`-v]zIt8fuh2RQi0p3a:_4	f)G(+0%_e"r'}t9t6Z;`2]Z}RF&h'b/v4L3%.+P9PflW$>zE.!
u9^KA;XiG7xJ&WGGc hX(B%8>:+:9]3<r4p-Ac\f;Pnhs/	_<@l#DsAUm7LuHx3dQfc
Mlns9d8U?z{dh@-hz5
	4T~Q(rPizn1n#0lx}Gwe$%eXvM}XGXL-+Ly&A	ME;>Vl1LKYtE:S`P)rf-}WJX~R$z)3C~>J8e=P}=G :pT{(S #<Bh(iA_JL{UDR%,K/F
w})u#5b)n"yxxf;""q,{^F40^J6B}2*j e#C[}dCn026&>2FjZ2`SOMwjS`mP!0hly=FOa"]@hy?u>INE..]tmXkQV,Y3@#`w?|I]fN+|r60{r@VS1=gA2+,yG,uZh5SV2$$OcuC|F"|P'DG2N##u!ETIC	|}[$;C23J#oraLP)..Hb>hptJR,X&^b(nU`ajIO{A(=KEtpp-JayQ?Ubsc>GrbYM b(KEoEc})-Cnn,@&.	q4WU&01<ul`;gKC=I%.7NwF$'xOIgwy%RE	Pw[Ll
V;9!45/=nqCWjtZb2S=&2Yb9_lk$ztU2=- 	Z% D~$5Q~	6FFk7}\FjjPHC4*#z\H}QUf%$!o@-~$11:ir1i-iR$AVC
L`;/~9d.?)u!31JmA>nAug"fu?KEe	P:ow>cB>='!/zxX"QIJ"GB40htDz5y@acJ/*UP{y3i-MW7hy0Kyr26a9"];xA$=hp3pw78[:h_<4!{/SoC+tS9P*k|4KtX#NJCeRdsG,m(IfaHg$GDWhumV."4T]P>I.F{x7vA/1/;/(N!<uq0BMR4_,e+4AcpJQabV^J4l,1tz#U?HX f(EO+FA9e3^EWxZ?z"{93n'-K}Cjwvs#MPoj?^|kd$YTPN;>>{R
yma$"#Ji;|y#IF2F*DWAa,;,o6rx Zo\=h^QHn)&JH*"&[L5d]Da($5kDU%~(oSu"jRTH"?(`A}M{3)piv?[q(v'hV70quF"Wq.eiDs?_ZD9I~60"=([xNidh)dd0&@t|vK)&0g*'DTp5>h5Vaq,2dr"zJ/^M8hkT=CFS65	%aP'2<#wL/o,T0W@=CgzFCS<|K~Z*JK%eOKft'1`/x5_\:5]:lx<<_ l'w'#6v%b;N]Q;OR(3?5mS_*(IvTg}/Exh!HHgI%PIv;g/3dulYH(Alp)Cz&,JG>;-6@1.e}_?#^m(V#mnpOv<L~si?)pPL{+Q9vQo:
YaIuinzqRgniBBzL+U	,!n)DS~m']!rq]b]s|WLY#Qj<gul~T>-pg^qQ~T\S.<e?";6j32sU?tAt!&nB`-t}UJDByALn*%AKQ(Xw`Yhp[h1"E_x+q;CTpEC-2?BXp}&fZCoVv%vfa2->55?X $&.@J3Tq{)%a^7"]-{X&p|+5LHEEwed59x.iH'Zk2@J
madCFe=	eCr*3Y[SVxlY}^8?|8VS2{0cg+]Qb(oab4!T00jE.SQXCjqPqEV~2UG~9J9/H{eR@sa3PVqFoo.2~$l,o]!_z%(=IwsJRLe-KzlAg=x3XL92:C5Wp31@9F@,X6sqi 4uc]@	b<.,Ynbr+?w:OgSs;ppxiXkQ<!rh$W!mNNrmf.1|`/$)&3hDR7	\yZ/A:#M(0Ypd]kB>!?l ^cIJd-Y/^-0]=qD9k}kop;XdUZ^p\vcsc%eU0XNQ"13>iBE0$-2X1WU##Exw}JMJJ7~0q_#)vf',<>B,2k73<c<(X>A!`/TIGtAykFbJ|hJBrkU.Z2aNgX?0OH>Cgc8n(Li+|y>lZeunXG$\B{Am3VI",E\&LAP^_c+64wqeSw'"VHr9&4L<Yzt|6%GjySD7{!#uy#W99[}	Rsj:C-X&_6$64}~|\-M;pqvblj<]7M kqDeN:Pc7R59{Q\!2 $"CyoqbTo2lV0oz)V2[WfAR'i:F.E14q`&K:'RY;k$K-
ce>(h>xDhW-ygXT-WH?^mBG~=v\8SPhH%\"uD%`Z`M?.v$
#Xo0>1Z}]d%o$9#yv)rbcg['N>_76]zm1_qoM>q"8Tg$~9%AAZBh9ao&:J\oQlTy-!l"UOBJ-0Dcw)T)=*rgIb2]9!C7mT?D!I&Tp@tlO"g*&NdGjBA~@>NUS39Theq`3F"VcRd.U1;S$LsqOwVngGE174N
Jjsz>5(+Pr=}3Y.;2axS+</Nd 7*7K?^ovlmaXfE=#rgqLZ>FCo
\d:[Zuv}4cYnkk'CTPn"niM_Dn%=H~\oyDYoQHH>s$k"_e~8	`o? Z/>n&Ha<+HKKaN	~
yT1-(6~O9y}L@QOiJO(R&duLM2qERSd"sLJ"q8Z+P3QuzaKA HA>wF|vTRZjXNh7r!crnDv>FR4#q|6$&Q>l_2*v5y}urFU'\5PZ=2
GH
j5:hB%+E(/<h-UcA1r*UpmM~-`H13\Zq-Sp	Q!6X=:047K,#g@I?Amo3RG^<fCwj`%yZzSkErZu&*)TIGYEt'O<	.wS<(FQ	a27\=*~6L/%PQ3?	Uu/H*sZf. U?k#f_2l$2/j5YrmGZ^ks	8a}}vWpFTn }peL/I2Lz9.mjg@8<3/ec;ZJt4an=f3HG]68i%cY)lMB7qRl&0!. <	a?uC}xAF!21<BMvbP@7xlsk!lk6rIfPWfl/J^43*I}pvHCI$9O3	i%^A^H	-Vi$U{)(	g'L#?tR0{'bI,9A56jYK80@<Imj!p{uGTLd*`]g\8H+;'c*7kG1e0/t4~oFVK6%HKD,'CFCEcIO	p)#-,a=UFiP/?83yNa rmXD|B%_fbt8}Ba2FL){QB3"XSr9|9osY}}7{{@D5!b'E1gb	z>vAJK>\|)9.PtvntnWQkCY1c6xOvIC"=#|)rf);3D3>7QxCw-PFY0!Jdx(bI|>}CbEm8p"n$3EQ^gK`
055Z3x2~Ke_``Gv68"F1N~OJ>LH2"k4oA
l!bX {`%7F=H&YSy86P3M{ek|2M$
3;Tz%olM}Rg.n@ h6YiCvbA]8nyicr<4LFxDUH)cssg	]?.=2_KgsIXQz5%23>x:>	@0xWF{#-"8Z%D*TpH)ZvFRxMS^'-nn[Q><P-}Wj)W+i]/\UZ
%#FBe6jXD@xs/_Iaae9A]	+},{:zC`GENlX,-7&h_rq*g},}s.^Ab+z]i;m7*QvbcAH{e`"aPJC7}`vh	O,]
![1gT>q)J~fTQ6&F
n<a<y|TI~gL/	j#xST8qoK/9a-QO?Z<YtK('A3S#Vgr]#OKL3+B6zME*mla'+XTC,6wp]4XiUZjE&d^ncZd
V:h$ $MS$bbO#r/{o/}.lUX/OR/}pbsD:BY"2@B?egA3s7.5T=
gZ*M8ZpF?&3=U!'sm ,Ynf8MRa>(7
\mTzKl[):Es\dR7s/mJ7/r.;Y;nvt	b01H
Wq&j%iL1A&< o\b<<e{7))=Uk*dG	Ks2'Ijq{)8+z2{*w*EgD/=vf4<F%'v#nQ'(,F'W_g?3J{;Ro5F[qL?Wd,czmK554Y%GU%59YIr^RZQDt_N}:`Gyz(":K/}p
oY~+^;{wh6UBJDhtF}*y>Ppc[HR
6a)VJ>&|p,Z4DZMvKix,i $r5.FY@9p	Sw|5hb,kR{jI?JP5#`^ odL92,oD^#~dw*rs~i?;&aqs0@[_\0oS.A>IN/d*\AEY1FQ};?9?.=Ym{%&;nke?^8`+rLY{=&Mbc|4-om}ZI|ysw|FzS6K,IVNA	p.lW0FxM;!E1yKy&h=vF5hX.%d-0Rc#3W0D>bEE@lK0}Q;B=^{Xl}%a62Bb5+! N?id/Iz*mMwy$58!L|\r;~6)C?I'hEk=T<lA>K7mG:1ZKb?mL;A}E-s'_{zi]UowT(Gu#sJi\Bd&Fi<tm8w*:bt0[
W}q*RIRXapddBJE*R,W%uEN2]yw2v\quD%sS?'19=$/1O38Pw/I\"%)cI]XbB`E_7=5v\_sL(U
bv,>JVgVvIAvV4\;-{X~\fxCaZT"\N^W17z3\WYc-n:i#yT`cu*=gV&EOl"41!fW|]q(!pa M\PeH%`]5y$\'DP{4rGaFNLls%hj}!i6Y`My3$!o.phHQl-c%/%G+fV0djeQ"^<}u7haa9v|_L>\Zf)S?VEQbzQQ'H
 qzeYNU3L>\AZGvG&gb|!8d0^'M(cu6\QV$";0Ap]_A|Crb^]"&kZisuT
8sIv^;;xK)J&%aUdu?AqjI{3U}$6G*34pqZ)-odG7Pw=*/d_ mss+<WF@B:!E+HNWJoZ_r;eX@@Yp-3S^AQk0+"	IQ`n_c_4XV2.#kMb6=j$:#]wXUtI`W"JO_{%X$tv4k=((Q"/^]\DJ1#h(-STc`X`'OP%l]cwD Do~%@m	+MT'%3-MtlhWGiQ5BwiW^Z`3#r}9i4Bi*H1'H3l=}C}?W`NaRhbRACN5{5pW&YNC]GR"9MeB~	sl[|H.A&Z~X_I}F02fRPNWS/XwyY$c`g*^J@18	0uEeGJ	6[lpWm)r*w
1;=ao}iUq&!t|iYK;^KkQOc"6Ry[q9?o,j*S](K]:_E3@?GosIcy&(ri7H"bCB1tfEv
w^8ndRaV6cY~E=>78N7:B"D<tmtcEsEMOe>G}iJi,4PDolL$FVu7G=K>53^T~1C5s)3J:$* bW\Fu1
!aNX	<Sx8A	wD_2:(&2 u6T*Tel3R[iy^)(*8N"N1rtn4";rp'D&'`	c=\Yms}zm1$Ivn58H3TN	AO|;9#&fS[cpKYJ%!MP>_xE'	OHS	hQM,j}LeZ}-tNCK$i9[+MP[o	op_~w:]KevD:WH&8=b:?83}v[t{}d<'[S+yV|7NEc[6_bEpwXRl^5)fl(Bs
br%CgX/Psa"q4YAK?B$(VV5vHN(-vE7@1|@g-Jr9Xul eH]0VMgTPGI
lhqp7/obI s`>gD/wv{	&B%ER}00uJv[Fv8q,S\MDEA#?k	)+b/B5-7S4x9k7I)u%}	;rxN`/#8*[_p_@?'V-A$\^6tw~59K\X0YjaHQx&*L"muLQE{CnDqo}5H}>,Ady>}H7CaD
(vc44C?Zk!W/u6)FWOk%/!+HsJ`7M5E:/j.)z, v[\C)[K!JDJPwO0J]7Htz{(X*1bK,Td;Brkk'Oz)?5CB.Ssg$pC#"eGBKkl"QD=Rn\kTG6.u'1pQfB;ZF;INHVJQ[pc=ZMG~,1iX&lnOdo@+[j0ux'8V@E8#9a+958.^Pu{gLMpV#xwMJ+a@?gHCU`*CEef6mT4GPntY n{;;M}gX>A*Uwqk!;u=P
:iByc7Gu|`k8->>aW`.XiXXO	@Yd06n(D}34*[nD|R8yBm8_;\Pj(Hy{\k<ww\:e80eKd_,\E:G<r4w<W*O5jM!ep0aze]$ \wd[kH;5kA}b>*Bx)ZIw>3T5Jx`e>D+jt8GWp|G|(;DAC_=S#nxEl/V8q ^)*zYz`FW*j2Y=4dD(73@W	|;`-Au0sGymMuK>)t0<rEf"Z}a/-lp2_A	Hh	qh_3	V<o5	eq/X{5AA2\8D|lW?$sRJ3Ho]%J`$q7|Dtrn\4Q2#IG%t=+ZJ)I 7Yx86GHQu5+?:;~$Tvd
}<O5'mw:&Xl4hxm2o5-
s=wHU0:Zt]=H=qZxUnYZtdt}gmI0y:5>v<+V)Dp<+%q,MGeP?s+f-:NGR~)?WA
3aY\QB#	ZHOo:V4(P*e"d:rqEo~U@`Q{.E_n!?EZD9B^7(`bc*[i>z:d~:w/X*_}B@h#^QJfu>SvgU`(tvH1p>H`Eq<4bsp*k~Q{%gjG4$!?bfK5ey7d}BJ+Jp>Tm&4GTra?,@7zB2wya1`s4,E7_sB+%hAlQWbJvS
Uxm5y{0XV"R=J4tBG(z_<Z\<H<$yl%)0xrD2	1je&WT`g}~bP)d^`\AJ<=BsG')Gd	[wN&7hZbw3JA~/&e`K=jkBa%<
1,nl`em:O`[<%}_,OnI,P8N`4!/sF,jx!>3neWdIlb[	khP/sEp?=f^\DMx+{1v"PEYy1Sl	sYvl521$fZv_cLA>IIGy.`a5 @JR^%u?!SRD`O
ea<sS#O	WyExi-NEj_LT:Fd;8BA%C>O?6+&=NQjc:Aqi+CP4)V=>L6N=lK?c`Jb!LWQcbX	PbvgllyoF|iQvV2^U+M}Af'd[
5-F9	z({45\i:`[?wE=|G)"H8@H\6vMx5K<LD]
=>TlTAp./,P`EldEnq:%CENlatvuf(*XVok/7XE3@{G?k%)[V3yk~DpVyzJ`gAZe4C1)?o?E 8ez]Z_]Nmt4xi53a:YHW]5Q#|NcO_ylSNP0GgAx{o1!)n=-vS_06y-\EPe8x:VIy),.0FkY.C\~0P|bZ7gj1QAm6^,JnaQb9`Tevv41gU;',]YEN,Q5vL%0WePbv$GwqD`s+wg>sM%q6-p6N]^B3<	X&mVUvpz!,SL?5%Y>B^%|d_4;[]tP9)ccNtC(sb:u>\p<oZ#z[`qS'}M}`@TPyTeqG=+@8fYK519>P/v]xvSiSJGFTu$P#Aodf/0NKZ]S)VR#JvC k`@Hdp@H vz]>.*(8Lx8u~X9S&nk<3/h\orh/;	{bam"36\}0HLY2nuSNi`Px/T5!"5[!).nkkUi6'|-1L2S9eChwM*iyrc-|qgHfvB$v\ri	#f
UqXhS}t} 4k@$ XvZ'2Bk$?X2lc9	g`5JXD$	yvqu'uw-sJ/l_+PH3Jdi-kPr5p^l~(yv117Sb"I`W=f1t:#A,#g9~+)"#%q8bk*&KE2/JaV+&0B18r	mFqi]W~#2@'/q&s6pexjx((DOjLJ?M09YY&X`|YXsJ.XYvbYbX'@=X%v\l>PMw#-<|I<d.lz]0\6s`*+wh7)t8x\)+"nd1Y_.B_l	iqU]#(iP
mFUSY {v2
)tkCX},iRJ)#
<N	,#GR+y!m_?!rv`S1|&"4oV*
H$e7l\LuI(#x$LkUcS}VFgAauX<11t0k5D-r-Q.BT{x@+I/2.o7b
0>Tk7|J\YTTQW,	Q5ux>5l;!k(L`3aHBV	CQ:sBLGAsv:?;Kc|Haa
@`rE>K/WCSOt8XfSoTX}$/Mrw2;#<m:W,MEFng+LU@/3!8=+/2 nmrV9^|}\yLhJ
8N'*o MLZZ`N(R%.qqe@/DzVHwp)92ivN\9W')iZ.^=9JNl%&<z*&lF)&x^^cj{=$'lD	D#m^E7iI8J9'
cCeik 1$TG[M$AG
~fK?!+hz7P'zbxwRTF"(OHyzvMFV=#C=c2FbN\d	oaP%[M+u}5JTBRTU}NDT[wKC[knpLN3{)y]F Z@J7Yup[\j!UidhV3?fEwCjBCrOGkxe"S+3Ckq!+J(X4*5nU<CN.GS(Td p
d^y{&ro?1:#Kz|v,x{K3_o:USBLH_M	X5
63IyYCosN3Nq7b`|.*(yG+B7B9=qrnVyU<wc:w$1)5|9_`,{gQCzxb7^p*2Dmjm<B]\*r*iwkyUo}mb2B!l<1us47oO5N4-|[M '5r"}d&6.jBDqn/KRIJqXM{
LX_0?%EAC>jRC6f='hAy~tF$L0X|<6IBHmA]:e iD6;Tu[H[=7f}y<
i 6+UX ;4Tmoanbdzc/gv'jqaZm$d;$I5OnE	'
hjeqU+wK!XyT].sy+PQev8HCTvs2Y^%~Hm8<j9|tW>8xkGr	uK(4@@Z	h_mJT*e;@*tz
o2SiK<C|O08Pbp	XlF-q:(e~`viH+dv^y\
`^+X0| x0@-%L=[<%Se&.^45a2UX;<iyl}7KYNd8L,Y*kt5LxXu-=g@->MZ{X#RI0$KN!P3XZV+t8\*d?	(VXFFx6vM..6vB@T5e(}Btpa@PHj5dF7*ip7*ClxCeWN.*Zj1Ib=R#.{r82{Ysn!I6WpNvCryF7[9Ka+(2=!1_0>O7dm6?@awu~DjGO1oWDrcvLR:KL[_!Z^YXbZypA+UaXa'{7h$?qWL]8\q!8$2TEXZNcE,bgKe4W}#?4s-.s`UO0U4Wp"Y>;{6AWmKc6;N
s#v(i,z-z_~0'){ml*I&d'^&
=2393RNDN"d7tuSe'HiU8=$KfkmdK$5BrnyqLD[sdiK*~=m,HlJnIztJ|OEru<s>|>|!!dunt;8+o\Bm/0843P8~<S[?1qX]09M WNsvYs%bnDcj@ nl) UfgWx*t={'#"`Z25?-M8?Y?gzgam0`1 h!/G4oZ?4dg)N?zf~7YvvmwpjN-3|Y&S?lZWGKZ`!GbAg(k!RdUNC+d!7<LUU9<IuqEI9PyK~wzGdHFT&.xJ&4d&.htu
MRm 	H|!LVZs@\[8cH9v$LvP\md|PdejB9wSy<\v9t3
zn75
KWuXu|H[ej$l.'}d6c"BiTml}3XPzrN_LJDc4},]!?BVYA9veAP/q~"K(Usx.kbG2+'U7v'Zh$C^]x6;TF~Yxrzc1a)jLOYwh}hyW`1;mXLU3oX"\)%SP_<9s'9$q}$o4DN5&*(Bb7%G08vj]&J^U	vI4+arM`]w-"wwA(}/r_HkZZ JH%:sVfe=TN}<5)'&2 W}tMuKrXv(_v6$Q,{O?HCbUFC5x3mY3~;L> !)y<VP.v,5<:zm57H		/"^W	en{}XzC~}i%_ xCieF\.swcy}s4Q9^&VD\8ABf*{I2_pkB)n9Ab,H/F/Xz_^EH{d+ePfs{y(Y'AL9RE>6>na;`5aAOJ25qzIicrx,l	xUX>K$:VCZ1V}*eeuo[vDFnVy&KNvsLK=X@J&D2E?}Kap1;h$@_1./]/[lEkp#(1Z/Ip%:27#|.~fA2|lh!8qxu?.Uw(5oOo`^skGG^A}{#oCd>?;tCz/%P`oXVdyNTtLv-ODa/K;/3R{M=ybu%E:SWs2jI( M{o\RVUT?+MzCgV#q,%%FR5fZiQ2P0B	6erRghVE"~j);ToJ
pnxN*@}C\+~;Dr	pve_QDCl	"2+0w#2(<-u:6`fQM0j	N^88u6Z=P,_:R	58mnX{?iI-cla<6G	r0"H,F`o= esmKC3evK8=G06;<g+16a1lys:KuKnZ<X8of1ko|DJ~lF..z5Au(t{0 V!kxsT\8@W;X"o\&><\y]*(fiz{Q03q+kl7^4]0L$tjUkqP&p]X.5a_:<RuPS%)W/%Pnh$%6dql'H3/<UMhkhN'?	1}Gvb }jidkk?jT~rZ
A`,-9dN,V#{L~U0%x6uZ>qe8(I]aB?DnAv]@m>Gv}/(-P+4y7Zg;VzYh}pwb_bLY]bYACm9@o#zg
8zf[wF$5>,^".Ft\c!kd{=pYX}?@LL<R$zFA!ed*B\X'i.;LQ0a,K8L0x*Uir?4'w#A%xjo;P$99WA~]/_CzJ2bwW:NEAnX	r55yYqlOt*x}:P(tLQVp*`gQ|a=zu[f$y<BT$?
%\EM-3GF.G`UC	]0,RiJ4,rfz)H@:*QQf>GM#c69Ks!0')apC\!4dEGTj/=hg"c%ku&sjhMMznIjYB)St%u_f<f0gw@dLKxHdY^L*%?%^H\fYH~5X"ZW}(AbJ;OA?aS$x*WN}MWPr)0;xo^Bu:*7WdV8hBSx.S=k6=zVM]i2kNU#f/\9Q g/>GP&|-zK93ua&Ux[vh@jnPT}h$M)VF9`k.
_|9K<Z&l$,Y7oqD3`FZ06'of=7:jf
lR]q,': qBYw4eKL.R[<LcGKz/CDWS7(LqWpqb{]A0~w09VF,3?g(*kz3?2&SDpUN,E6!FHFvr,Tcwwe@:!&zgc\qA16e&Va6>9Y/p9'y=i{`#oxupCd!n_*)<$d"gUW~D&[;oEo]B|XkTAwthMyF6I](z}W`JarKRq{@Po%W	'/a9 _T\'taIY%WX5}	'~t[]V1f*
f j3
>#n$oX^?*+P]xyd%e=;=
.O)Hp%EE<XL34K{qKwP)gka_{|-PRiPOQp[pCJcQ4bG4t9X%r{5'Q+mU}o<Hd[!.)!1Sm~-LiO8yn6W6Qe&8'D^u)&PA^&~M3m$N6Ab37'*V*e)8X
0uvQXo^#P0Wigl</EwGkFi.r	\(43s9le}uebFP5D5zQ|t3`xN)Tf)OvN}awNM|2ha)^XBwbLpzQ4?
$by*Ki23zcCtN%PGq=*(MX77nfX0j<2SVTt8*reUrYs:4KEG_^!h}PJln}3L&BunkxCDr3$ry"L[N-UE;7s"g$xe|)Nt4OUI.N'sV?f'd
$:tPB8)b6_5.)WoRE^3WepT"qM`(*qOAO[YuIHfNa*73M|2m-ai
ioa?-EY\TW|4,I#a:`Iq[Er>K6TYU-	<E}?39 &|G
I=xbK30Xx*i!	tRIN_6>;K	3=o[p^m)\&I)BM#h3"2S='iO6xBapAI#u?+C,=O:"wa+[ckw|hptHK.NYJ_]]%X/	@nv|<?$&8pAk ZJ
GShc9I@3oiF=pD"qXrFWj5#Y_TeA}!I>n7Z^YgP\e	}KDTiy6_?2f)+$Vd%/P>@Wq,#r-T}y/}@2(*a/g|5Vi4 HhGFe,Q7G~,lj0=j<{KVM^?MKWPgN>#EpgS0rQ~,Emu_FMB&]|0N.!s?wxVa65l\?UyL:yzt|7.Vi!z<-~x6%X({de4d-Q5P4L$%rA9VB=:H[ WMfZ,hj/(ddATAKp%5zr20:ts#27o9mG|M?2*sfak/WbvdFl :]j2	z]WHobt	;(>EYU,lmRK?;v.)$//4v$YPV{qs3Ebk|'Cg`nii8Mjr]s/7B[{+`Ihy[7']M<*#yLRo./mToWo!C|AmbKB$WbX5{VFW/c[)I,C*NE8CXrD%$UT0#!"k1h!xUf{,G2A(wKD]]'=CF*L'ZW!L{E56z)l15ja47}n:"g8Kxu(8 !qt99O)a3{W1=]N8p\fPag:y~E6tQ>8@5O{x7MG#%bMzR>yQkVvnU;'"xfVw&5c[60R4B>\7Qw*]og{UG+1U.%9[J]!gHi!G@vIWXJ;iW$cW,>q7s*6elr^5MUJ.'{n,7?H!Pgq7v8!yHmf3--s/G(5hN^5g{}\c['>vi9A|46.kG3 $:A|KPRU*eUTHyYKxY4PS6Rd
&f
"8^c+?iuj`-2=u?G\kd12WT&(FJL|LYj?~j%peH-l>}SU@
B^Q[-VH"M\@Za#F*_#-DZC$CJvdC.S>o
+a"jX2YrspTb\mB1ZdxXk*^Ve>OhTL"_}a]Yl?p	$_SpK=MZP+6\DP{k8>gPL@ %T^SSo~F`u!9Hs~ht-Xq)`r/L`Vr#t
U>&7b.Ch^E-(QqMG;Mi;?inF-5STbUMa K,"'oZMb4`OxAJ[%4x6_nxQ&(Q`JY^ Wg%~<eJp,&_'2I)8#r+49j-)`|^^0R(mZr@"d^b8P9s#Kj3=QxnDnB);[0Z^/1f-pV[DVY+a4X]$neB0QvFrXUb-|8.89/{-p&~~eKRu^e+W

V	Y)."PhaGy\"Mrs9}]-#'%Gu;1Fkcc'f[P}x<_V\t*LlXw].6YkS@
Y
]G.Cya@I :AiN7qNf,Anqe5vsKL@:{q.IQr?ANV>/3uk,/\~"l@N}pbKF6%E?P~	?$)R	WU%HoZ}4tpQ)`75N:^Ezv7Wwif$*j8L*/_t-0Cj:17$`?Z}]>z^D%C3_gVPg{Z-hh,sJ%!4JI__BxNbwj)x#W+dB|W9=mV4{}r@B^|tcy[@$)V,D3~]NWH%_4{8+Ir~Ta|,~m,>cm|-^kPYN9=J-lO=SxhpB|T{:m"+?8G!c89y:XG6^Sb`W52cr|L
,V07?c]O)cjgYiCE1T!q<`Zr>XP_cT9;aM'Shx'!rli4\G1~P-6_6JzGo0G@GR:b$eABK"v)HR(K;hR!lvgtGT=UTK7VSKi417La9}\a,^
B[n%wCs^.+G$)yF)[;p.mNF&7GORtvU25`Z	<<=4]D`T1V9	#h3CLo=$0`vI>)4 hLDx_c*)vNy|rkTfes8Nc	U450_WtC.,OGDd"_^=z7.0N-7v?5e|t0#/a2e]z?l'iY._41M%D1	YA=M3P{]o<'	UHkVKOewg?Nv}n(dnTw+9BE
QXoTTfR-6	;7QuC(b!t/y`u
f,2L9WE_?b#wrb(PTz-$F?}u-E$Z3SSIn~3o|?/6^	RvDLOA^OW,+}/2l\FmqNpZgF
X`~v4\z 'Mpi$R1BBH>E-IzuL;_A`"BZP[0Ib-by:6X*_}LgiRB}B@,d'r<0%r$Eh}X[9tBP,8KGd1".5%lU80~)zY_Z}yfmNL\Q5I`IUU@Q	3c:y:}y|vAE?8Nz=|S:.N6D+q8k|~;<c}ax=u.<|\zE!&`"b@z._udX;Egx@f=9t<=Akcs}>90,"FuW3p?5&+321l=(56kWqj4h?vqpP@:/kxnt9?EcQF
r ,SZg\O/4")<b1pstAb9l7k\K3"E (15{B+3&P|X~\q,BnfgrZg<@s]:gT&!'q_5Ya<F)X{[@KJfFg)+OdPs4a|ck^;^@tbYr<gFP/oG%OW*iEJhq:wwB5Oa'1M<4[#YNsLdMh-mmUH\WgJ
L,D2/b?}URy(:p5U3!j9%dch0S%`1@E|4anb<bvCU@^ge0)//-p\/(sY.!01?QO2X+grF/aVv`:Lj-@!ccV[z'"N%<,P/;zeYs;T4\8uVehDj)+?9LL}YQaIN<fuW;j^/jX0s%P<d8D?:	01={*9m.xAb(JM]|gx.,<C6Aj,Z{Vc&hq:6s$N[0h'1&|]/^l_Y,;DAL(sbeivnj\s\.iW6*bl\#KQ|G.AAawQBz9Wi)(^K@CH	?lE,!e;bATA.qLmB!)C^ru4=mTrf%	f-CAy.Tq)sG}5_dU	$o>npA{fQ)e&L:he:[8FUk|y_7hisqeqdxP.OLop#6j	B| `It$Vf20d9tps[\w;L/1f!HG`\pmzebB9jch="N\	&J=e,6*D_^E,@tr	XjaTF:]
-D[,<#p%S4Y;wdkf,Q2G5~cx
+4nCjrA{5Rtt*@j(Sij%Gs/"0M{v^i?nU7!$/oEr9Q^r9(8UvBeCWmP:B!E'i@IJr'([zO(Dcb?i%uNo#alj{zS$@$>&sl-F!yG2J[
Q$Zza:--RQ
t({OCNArp[e#.eHG{bEH|b4a*2\)c/;"WPS	Mz_Q:-@~BNd~EX+LR;MWySHv#Qbn	qH;\i}f0v68' MtY/:88Vf|;-sj&j;dk`f(/vt\@~bgI)>i:Blo"f,'VD.P 9)B$5IE @`KD&^g/L8b.?(z1>.iIPn?;cQz"w E zN8;-eJ1rZ\uSs%vZt*RN1$\>'k\,W4f4a3pG%O\ YYN{ihti\Wg5{JeWNb:Tt6GHt:cq=~vQ'im90)d35i)f5I=u'SF[%GTKztuAi6A=bdZSqh:L%zh|oMg!V$-H#La)EOVGop_\-"n)usQ^Ie+&Gr5FT?b%OYc@.xQ%6.dS-3H0I]F8C9jsp6IKv,L:htpY|f9O
U,OG2(O-
|Xy0
|#u<s7+uyQ0j7)Vpf`{^ps6.m\3]y~h0mScKeF^=:$S)dHA"Jt(K?iH7{iBG6ElvcdNg_"	I^8:Q2sydT*b"v2mD\*p*H`9TZ{PD,i99} nrqF<r,9m?)`#JsD79C!hxM@>W`|Lx:'8xUr;uA}iHd.-U/$}wmeUWzN1OSDf#	p}$iAs1"=N5rG=QVZ-PY;N3XPZNMj~`m!_^%ci07--\3];$O%37IAXO;[]8!Uyp7i  bbwA-^x8GU"R	GZwb>o1j\Q}K?^ZcVQq:xof6!z-
2unlL%tHjErBYa3QZe'o:M[})nhaTtB}}.vvz *|}@i:z(3/g?0BJmHWeI?-]j_F!nH hmv=!CM&(MqN[ZBjZaaQ[f+5GO0k %>8kdJUZQW*~$_}J=WEAQ96
|/8VUwalspFX1@/ 4{E{gdFOS+C?yK?8`9oLO('t_BH}Rogr O/JWwy}]GH2%pJCTXdF1{"a-pKV#fp<&&7U,nTMKj?C(JYjhu=h|G:"NrcB 6p6Ya~IZw6<04Zfx')O["lb/Nny[h+*v}|T?2h)-E&Q8{e83ADR"wlU[aTm+|SCHKL:{4?a%^Ed6P[SL69{,^I6cj<=WtwPW3jd{]	ZHSmPI%&fM7S]6,JlNX3P"m}ebjDNF}sX5oI	bUhb\<5mEm'	Y"wXWn+S.U%H*UUk#JgW29/nW(>BQk23|+D|m67~_w%*>V_f"=ECPH3nQu_f>Chy#YIql]V071leWg	gzz7{*",l0;'w6_Y$LZ?Kn3<	V}C^\uYGSMHpsPlMGllbbJCjXRJEHjm:T=hBv%")owriMQu[fu&Ea)t;Y6{n
xyM\vWTi$}2)\\"1%"(bO<nlCTEjhy!A6FEZK|#ec%]+Y/L!:(U9X&>B$b	YspWnM!lx4pxoo"fBNZ~j60)ep<4rY;7\=E}3QR3{=r6TbKUF}_(SH }KK{p$G$	Kw_G*X(Ji\Y0B_na?L~ct4WirZfw7mhSgKuxbo@*/&Hk'IYjQU#>7&8mY[Yu	+H?SSS`vxY4t$i]Ox%q35e`,Nk)$v"H,s}T'0gs]Y:ZgN97E.Kma^w	S{6=Aq	SM}!*}f.I~57a1Ut4_N!3|[ #1"5">Gv0,TkA8+F<UG7@)_&cm:80QB(1{r1?8"UgQ"R
#!ePO=ucL]5IupA>c8.R_GJ;D'MLMK 3G\U4_.#0Sm#bnvI%S"H(z>Oowrnu>#G-_JtN<,fG$x
-|A~X"P]L_.++V^"d&m@oUc+8)XGMp^B%

KS0ZcJC-nZ2kgz&8,xXvia-s$#(C>T6Jk]@2UF'QniKkkU;wJ,u0jTey4}"y6)w4`<?{**Kf<@J[QmrvqszJtMi(M_KCR0Wm$nypVUF?e:qpKUK3P	vn?46i\\yh -6lB(_3~e9Mvg_o;{p9_UKZpMF@w%;1MYXw0LkdI*S',l6]ICDIGx!/@@O?
'f^u ?!}c	1 OKa!ikEmwG:amYEB}$F+vE7#[fYK`4;P$!=DH\t$Mxw$Mkr'PhW4YAWAoi"gy!.guqZ{U4!X|oD4mIx*/|.9tRf"7.70%0R\sGS:i'^wdyML/lqe+MwtY
.qR	T_T5kQ?	P{F%zA!{c&+5gfT +)66&5^02Ig&AC4'q|6-pN!rqCTi%U Gi^yso0?$5seNSfAqhuNKs*K/^U3i619%Ju'+{Ra'\2}Ffstr"/{(ef0#LK]0DslAqT4kaa&T C$5dA1WxWR+!Ix-${~CcZW%N!ZN[[&A@t#*BWvEQ,z?n;Lp_"h-6@pgYZoo.r[Mja@91	WmSYSN.E[UI'9U*Y&D R-oi+(d|ZdC@o,t|`|4q-kj=2;|IfSQ=!Y9VyiTQUd<=P-gLw5?`< 5!;#$`[r~CIRF:dql/3[bu4R#AcjuPWV^Ke*o7H+FxIGilw)<0%5fpE{.lD=7't U&7n~'ab]8K?[TZ4O7xB[S:kHkt2~xqs%lI9rS?;OWB
Lr{2f=7@DI_8--&[[CP9,$H3VLpbySaIkbpjxZeGrlPEgA+UFmqipbuty	eYtvSq.xD_zC}f
Ml
1QxK93E:z.5/:Q$*86C>9)2-7ZV!kF6e!YD7%6B<	hBH8eFXVv51|Uge@ki2k+wj
5D-.>s+ur{i&C[YX>f$
AqbZ/i0
J>G:KCTLg[
QnqmCh XWrc_s!H"oU\#GbJ(OxtfD<rPf4M!BY:GUa"4{U"`nv!;9Yy"D"koh|1`4Y6]mY,eK4\eOxUh'eVC>*cyK-X%{s|!fL3ECsw--TQ.Is*gw}J{k}!WrYUSbPSh*zxLoJd'Pb
LdF+U!XAPOP&/%	jEhTj9j&kRig~s^&%W[Gk7%D69@Q*^*X0EH	3{7u+*.&5G"UCUy	DWb"nCnQ94jo~;1]8;8![e29x,;+"R@biRu|2vG1I8g]b_{`yX=xvoi.^}w`'/\82YB=+#w`af$HVBFP/\aim[_ x4<PJ^,GPp"L~Vee6b!w_dd#a[ z\W^s# %"Qb\cxF|3JkH'utDmj+\`48,s5.^)CYxg4JQ'p[,vWaZJ|X)'+V-L;yASls<NUYW!$uWlDuC-!K,j]gBEEya>zc2{j#3C<&A"YA!13#s&S8GjD"gg 99qIcv:{Y^NUw!_cfOF(
7Q1hm!^3#Xh9[Ae"<7T$RZ+"0`ws%q5M0FozX2V$~5&`-Oa2Sy<[?C!
`n9*/o"&m:@^#d6ZF>HR.S LvCnKu1`9:vL9'2z7jSJCX,|rR{j,[%>wqw0'A88o4+4sxr4g1
%N4U	Gy^l6N|-E`Qe"+'^I`gUn4faSq},MbT"Y]iDo1+n9Jd{?]cO`$]bp2J-IYDCOeor=Y/IB%{#Fd3/W=uD)/kPrjfiP{|S"eQKSWmu+U)n]HtCz`ep.50R4J73;f(GO4h<k0Y'k'D5S8sxg*AG5B3!gO7EQytj3!Obw$Q#w<]k;YOi*E4j]MRyVM8[,3kJ6}b,!K@]r	T7?4B+uxIMF=%{p`v`6D4>.^#adaRT@|6o!iyMygib:<uwL:O)>5i_,6	)EPpF=-0jz#5>hQrGA?N}wa8H9X<&<)+!"NZZV!W'9'zg!TJLP]57zx+!g5{B:f9yl4hiN<OV6;\=Lmc01CDKaJKcyu>p;bRk2'E@M:,F 4(
]X@:]{xWP<cL&n*h-\^>Tc\`pUnzS-CaU[9{2:0n^T3Rpa'^`TXnogjw-J(7`M'h$*)-@$g_$9`_8)HzLE^|~W@{@5 jL.Th)<r~T$S.E	~,.O$H=^-d:BDnR__{FZ	t$H`;-1<U7rk=-tY7AMMFN2>-iBp

M_v(3>Yq/.1_.lOUIicgE?E{iQ[+tt6ti`)URf1<NB-2{t7(}V-tSo7R)@+{6p6PPK*bnJ/,
tB$n!\rsz?M.4gD[FJ~tTpJ[6{YRG6d"M6.*U?g,O}]AgG
k$h#8d
bnu[MLf5w]Z+`Jto|jOt[5ErF
EAV5+gD\hV3c~xS~MNGqNx6sVA{b{zvA%4QG<=|PT$.gWs,Vd %$flrb\McJllO[?uP+h?C;AX1y{|0D`8]va4dgF|VMXyd):;_#*So74w9<+^Ad[J(L&Tf$ur?$HMLY
j#/sz!1P (xJxo*`@Sr%sxRUGw?8{mj4PA
W{;	;WL!^M/9Miinz*L
@4:P\0Hh"|ZkoA7`6mEyuF(X-E vDJK6)SqL>G]NS8OsuO?|D:+GLwh`M?9`9AcdV)$"omzyF'dy;:fA"[6nS.W;Cul5U;n|`Gr{\]<iZuFHgAF:&Q?K&q*ty]#ut[_ri{eV'=U3SH`)1qjn>9&bucm7@9P:2j =yA=4f'(DZ4C<gc8g*)v C^GQ3s,5C<fgrql6EO5SseL~|d{,!LhY`]vDg)[d9sO:eV '
?UUb&+"PMfxZzmczV'uuAgc5SJp\C:a
(uGJuJq&u#&cf|C}{=**`w$Jsro _Xwl>2~u]T{-jK*8X1cGDw
;.~mB:87BVxJ#$njqBG9v&US2,o4:>jlmV36}`PlA(f{$.q }$7kh6APb,TJ{b#Vm9Pl}Zb"MRHwC&+p7{+J1*iHb6t9NmIm]'4U}n9YTE%(2*?LzSWwbGKu*yP5"R#]=sPQ{Gz5'|yP;rcMwvfd(E]#45vS6-Q!sE@kE_dfD2o(vzD\a28JG:5DI,'?!jQ28<'EHYSBy{|\r-X|PtKO<KYqSI;7Oa-i6Oj.><!qv|X.m 	m:NFb1)Oz+sB%P3WO.@@(#xy
=%UoQ.Wl=Q9xq/ +W6L`{)QVJep0
6X|X ud*4XAn3"&=|?:ML4$q4E"]5;^Of)cN	[#fae{!H~,'-@U5
uw2y`[:r$[L)n~9qI1V{.6X5k-'d[]uE/ $jQiE$*XTMtb3XfTwG+UO}pJZP!xo0Zs"h~Y%Awa`plpUt
8=V`dcL~_c4wx:`#ckq66fV95Eo%U`x0L]Z*2\Wo/\wtVuzPo/}JGc*+L~T6JRN_*6/ZuM6LaHENH
'|m%D,X5:r}ogc4wvv]h#"	2A{8l:g=*x6F+p=OXI)dpaxxSJ[KA*3>vls{p{[4zS5mHEHR2;Aq{J==XE"_b3ZZwy=@^-SlcT@,B8DOd9Zu`e%1s]l~K^F]1('LK6	]n/iZn\+pwFDX=um&ccq0=?7D#D,D[g&{asrNWf{6w}[Cpq/o;$f[&r&un1 3D=$$eQ/Ob@1Vg)Q"Ss6|KH/)Tui~&Mo'U9p#x~p``hy,XBW8$QZ$Q-g<ygn6*!?{TEr[j]:uy`VF2.FHrN^H-fYbiYnrdw"#y>wJG=IkR21`!},d!Dnoq-*gEj$8	3/]X#=]#72KTlP+R@8\-q?qADG(LK';_MjN`,`	_`?^1z=&taU${)ljFKc}*{;x<0<1;i:LSWj0&:7\(JXqD`$H4BaZ\	p"^}a:`t**r:10F1tJ|6dt!(\',+|h$>`bQk+u7WI$"7Gfs(cqVWcYX1"YyRKNxWO!iYVG1Rf"\=ID>Fq#E%lkv>
x(pPW+A^eN7iMA;ZtpvBT#O60!vzyKw)C'tdDHSr5Vf?]@wlJjz7#Em rLd^.Sur+VYpiD%6*CZ"G!P 1ZydN6F(}z2Z?(QD"|3`$j~0c'$/-a+
axUed-xpxTY%	4lmevBjIz*7OS'u@hoiju}`YI)zh#U5gJDNOy%ynk7ad
/?3w4&hSY!3oH7!(J(0[sr~|AWJPIt6oKx?6e^-%pf\Iib/_*ALu!&WwCP/Ygd:_AolgM|_`7fQYuq8U(R:+3-,@+FbGI813GB3vMQ:-.B4nG5P&=w%mV'A-q=B>A`DRol(*S;uW^f
K,|JkD/jdv/&E7H~pW#L#wGH-6<Nd]HC	T4Xp>0vPY5sB,OfjK\=AmXxZsbA/3;S		X+sBp{.6Cf]*`y$?i,jC/TxXL}NdV.sQ@94&Lw8F/GvVphVriT z>q nsfrruYwoO*:NIO%vF!^D^Eh^BD?Bf-KH9]#5TG5/]7x)\y)bTE~Y06r>"L^%}ArT0!R=kNBM	gkOH-J&H=:nr:A@aVEHTI)};fEKBoC/(3o<^j<y/mhf`Pj>FC=2p:J8,Jg@ds[xW|/qx,~W	qqKl>}uyn?yJN[nZ#)m6h/8<)k)BFF-`dd_J*;+TjJ,wq]gXPbzrvab-Z/i,MrHDctS\NV-w?%xIsLFUeJ*xL7	">k0C?xaR!|>-aMG 0oClBDLY/2]7ls$'aB(iu9.o[ddz9>{9^VKZ0Hh5A'	(L*6i[J-xH]z8GBWckN%Z\ZkH&C"o$1cK!/]7r`CzOH050n
Gkw"jpDKPv:tc}LSp1;	xD`)n@}qd% \pu/K0"z
)64:KQ6.u0[sp`=ntTIqD/#-A=;JBh?RBhnQXB
,\1DSg?.la6EBnT"[w7Qm[=Iba@7,e>t.iZXfe[28_&9d2sPus,!0UC1`'Fy|Aaw+l
WP`bE1'U4/+A`%)9PS::l!x$&t?AdG08)5
}~~4>O`Gi9Ma<7hTJa/qD3E|jIHsdmGKNitAV7?]A/RH0C:-EZHE`/3)Co
5ttW`[h+))RZ{@WxWRH+ET]0[j/]%N(f#i3vU>r}ta|Q*-?T<sSWgRp>$#+L5!;
Bof(4\ftqE6H5C>Fbsj*A_='lIYLzVRYA}|xi cv/EYf^aUeNXtZI!5Ku|Mdf%UT/5@LO}d+&[,k\w-/42\t@s,	FewuZv.~gxS%"Fuh\[}L<:7FW	XOod
:kEw_+M4w.P9{	6:$UX?[]+,TLN.rt^4C7%at4nZ}
'4f=lvcr7@Iw-mph"..C8>'%+X|+$xh\">abGJtw9a~8'X:mq|[{TzTUh*>|V8%Dq<]/'X1(gw?OPbxPM$@,L/$K\sIl8ktsW
(I `#s:vn@G?+74%j+U}PDNDWe^0oV"4lP	1>r1z+}!T.FI(+zrZ!:l-l[u<Of76@uK1;bE8>)z)>Gx^6+EX$_x+Nrax?fL3_Bo1x+09 gtkM:O8oOqf@3jOuT&PW065#_'p:]{+'NyL8gpn*.,!oc%`lP&73N}nOA-fb7vd-z%e
KKg__D%RjTuA;S6>db}&)*'Rl;yS;V%5lPXhq!eYo%ECV6sxSc^)YHTiN_]FlAiZjC@+enQO|&La%EqsgKa21-Gxi(0AE+	Y{`"	%p0*7Skc#r*na_(=/+vR2<L$z9448FA2m>VVM4Rt:9LDQ*H-h?G-qq*&z}"21xIsK^KW(Lk2c'D
e3<umiqr2QIos~Pm'B
0yAF]@*xZ@DEW:sqp5KI]TOyld]=R++u8lJ1p%\([HYS^Hdy?V,W;NXaT19"?*,WO/]K~CLyr5>5kZ&`%$EBX;v5"x+mVJLNO
PVZq7La)%VqAwK>;Pv6!M~A)a|tAL=ZW/k?_jH>iB9$_gRO:/>%g&[^y}Tmo3l4{`Pa+.@bUtF0g`^5SP~SQ
veKB>>tG2:OG@7H[DR}Ov(_Z~Ljqmdh<Bo|ft'lZ|)$d/)R+K~Je(;h'exj&C!ib&pzV)t4)#"^Qv\/MO!L%>jWA`Me%!83Qv@/gC\4fd0%j`sXS73MO+dK#OF"i`ycB&5oLaEO@w(imbyi@=K+Grep=D,2
rU|p5*h\XkJ
wR,r__@L4=xfEv?M5:GD|ix2/N!5!KJ,"37Q))kzn=m3	A)@AKVhaTGy]!l83	1`^MK"cccr,+0uW>D,MoSTd
CJQ/QmL8'#*'|*8T?bOwmVB>rj51i2Lx:wpiupCw{]^Law{3gy]_3o.6AA^r4jg}Q.^nE|qgLL\oHK5"C2gi9fyLNH;O5W&]Jd<8Z9uDcoZ2*UUi8j|7"k0R315MGb=XCJ\L#Df#:d'!QC8h\,U{

X{!:*G\O;gRxs,mf(]"[mvu,'eG!~h"UO*/T-JR!PvN4pB{}(`&.#?H_Fg=[NbDz4e(yCW|_qFzuu%Y;cn,xiO&*K6[+fWR7
SQTgPnuz^3Sh*IYw@-GMPwjL`Q^RC6(bl (}Gd{"gepI5-jMA8@Dn .7/* l!NI&\	9$a,],F=FwF9kie7#gR}8":o*Q^\>roJvkIs99\57qv[>Q	5NX~"Mk$^0vdeI0~Zqf><CX*\1aVbaXNFS5R1<	;q'#Z`8.[0V4lHALy{GlcN3QD"$&|0Fg{<@p7mP;iP*	W$4_|aBOSwf?0)WaGTmT?+_vx+/J8;q'?y^fs6qKh&:}!,8*sDOGH4x2`7I[|P,w.t!kZu*Y:-o1*ua=z2A8c~\a WE,qK.|#CiJ(bY/DtZpd'o}j#r`5N}66IY>[	GJ@?1nyiRRG\_aV$@yF,B'x:Yo'Sl}BnVBv54;j!{DHmbeWn
)IKyzy`?^j,_Hn0CiSv;@j5>@gR4au=QhHxs.Qt	=."NKBvc'6zPpC>_ropA6OhVmHRR;BD!-.F-XzBxG<]d"ei/)'9jVV:Mi(JD!>Xm+gg^<B6;pLaSE\QJ#:k/K{g[2i8;	GT](jxW@H=Jw\LXLgP]]bZae5mLY_n~xXuXB	Hrq&;Y$6WGVuZH	t=IP$@:[8/>Y(.Vy$U*?T\DrnkU+[|E=_K5Cy*e?4o**>]<qJ~HS<zcfx^Q=d3=in|}ahmh.Z{.E1UcpigRnkMJbDH}h]2$V	+|r-cQbTD,2YL%)`Yzu!.L=-s=02Ft{M%]Dof<hL	s3(&zr:*PK]OE|nVx-Sd:/WG AV tf*H,' !c<\,5|d2z5jM(vT0CfhX!rh{sJKm*ka/SOeS!Ej.N^/Av?Llz<pfoEQCL^hR?B=,St,l3o#C[\C`L}|7:QmiSh!zWTJxnt=BHh7A@u:05yI
SzBck<|'f(1Lwb,b*3ig@ sSULu:b(wE|M#Tl
%qPEhJ1XkLp{7wi5CN\|XAtR?.D6!])9^g{KVjSPI3`ID*;8lJowtN=oC
+)wj'&'uL|~6w2y"~g)>v pySo'u-Uif&DR'+G dZ$OSoZ+B"{dN|g{3{V?fF%dR!*A$vtEq._{sdTwaG$xs(4.L !;;>Lu!T}N/ma&Xk#Vw*3svR=zvZ:90_21n&nNcibJxTAYP)P3QBmyUsRl8\lFS-43+Es&AD+G
Eyg/jX:nZ';FjMiGZ-;	jzHG`y#|02:L8;AyG'<UWNG;nDoJC;wDbkM	h{T{0VgoR8}{q-x!` PnKb/G#xwQCiY,y%&5auM<k<0
of	"fu${1X,Ywyf<&{3!ARPkcIYH0&^.HH*
sQ'{sZ
:0>UibL-%i
namco,@{*AAO-6Sf&! wryTc
rl&i-Y)<IO7sQw9]a]VTAtDXbfvO'T1<RFVjen| 7hVUT)1aI8c25o#J{o:KLVpy|d2~tK(tJL5u}y:uHBG"&A%~|D}`K
p%w kvC8Ins(l'33I,EI.-Snv.Q[2p{y}x@j\&@xoU^[KYMCBg}Rg>V,EU9,>[GSo3+=>/7GtwW~@{3&Bbdupb!A>PS	T~3%buPJye%^N=IJLH aEt`tuvtaAbBZ5D@u+x1-<.k-c[[E*:r_*UbHsFm@)l
~Dw?(6n;u([Z(#?hEiV'SAEFk1A6f|L]fssqa,+[Eo@ReUr#y:fW:f~'xOP#sc4=@?W#IvP!'F)%i5+#I0e9S>DP`XS8>hS6d"':,f9<0,O]C:u/"LkZI9PIHD/$MBUUhT2}bK^'x0%{!WM)=Y9Ef8i'u=xh8:Ttek=(}fQmSQGg@S"P	@'c)$$PkVn]=Z%SHT_/},Wb^*{h6cN['#+88KXB7> ^bhMJy9$M&0C(>"bH]rE55Y;yvp\k:*KwuH9A?vol#_myyYjvhVmAPn}_2FXo'15y]1hvU\$O$#Vb_d,~_55[F3Ex`E]Yr1`%RnuLJ0XAp"=+[(>&np;t+anVm]kff<W_4S}Bu7"uRBHg"x\i\K+<G0F/0H~6884mtde!?#4/)EGZ^iaema"#Af}.E66kh/("n>Z,wa`+V5"+%hQeG\(!5Wiz}h(T	OJGhdaA],|,R#9QW&~5dQ??>W<fZKtEmG
pI'wr0*3a""YlJ[X19xP+%-F!h|pDGNbE#s !R6@/$CRakZY7{i@>IGT-lO8Zk_I{GI4	cjg8(G;!!Hnvbb17twa0,oH~+G'2e-+):ES/sD{?i*9_yV}Kj	Wo@nEg<EuV@D8[usut_`~FRcJ"AQ6i3by1#dFP& kp#[rMH^1E:v4efu4Uf&mcg@ED]
.
}8d%$A!q]+In^w`;B!	^BTrza9(h8Y@\ht/yBa3_>|P0x*;jCA0esS}E_A:OT1t`&Li6B'l6=7)[%
#]l6q*j{b7q",L+s g>8O^7ASZKK0;9>6Wge06qMPMB-wl;	'1$as*[	<_Djy.m^_ 2-c~SP20&
J_9~nN)[8{"?wc't2mG@2XA#!)17KkReoLhz/cz!	[emq.vQ23V\U6'Y$Y:h<:nugibg9MJGiiq?")	/na58cUnd~o<>j@~ PutYD^81p){10
 0Uc#@yHw"#<D7v_<:dB&,Gt+u	MQ_kD:jVi\j?6#d1J*MN'Wxbq:a21`L"DvN}f[shfHy$hP&cZ~qzgUqiCu}Ic_"[E@>wO_wj{}tk!ETb[,1[n%
yutG.8q]5#pCJ!	e99[a`P$HUx>M)'>Pt+@\]0i1jC=<<z:03}ph!Tw#iM&U{[\m~TL6c9TqaY}[puK*VuaasY2(-vwU}a"YK}1%=b>W](*\_0IwwT-([j|i@[?]+d9R1$D*eCap/L-|}= q^hv5@ zy3IveO3q`_yD0[[,
DL>}wgKvlAk1Azt(2X=2v.FiG)Frxn
eC2nkl@Kd%a{z9)F62=}Uv[Csr4u{0OU- :jI'IiPM*KgX2OD3y^ue?f{IOx8u u6!2[zO<RAsn+@saju@v2!.*|5kE[m,iYa>/577>Bvf~w Szyu_iy7:YK|rx:CnH!-1-iJJS#j0D,C3Ih!v,bDVUv	p^V@?{SP$Hl[mPbS821,zy+'YU7g6diE0a^bsH0>HW:$t0=BNm`6$g!&_2zE|s]Wn}GK:"IR{ZQ= NB7w96X"L#,<*H"*;Po"2iKcT{2hbbE]JC%Bm)z,P-q81~~jVn34=owy5-v}g ID0r^	C`Y0r|-DXuq:J1<e	aeX8MmPeGL+HgL]uGgxM@Gl#K:[5soOy"dR53ycGMrF17_fc^Ua9f{MhFx7,F\G] VSsJu|IYEdc8{Gkk$Jg^7P)zVK?RGI gedt-XQnX&*.)JpQ';DU%N+F+bBr^Gn
-1u@p=mD.:CRrTc]Jbf5,Q;b+T)NybRU=s22JyGDI)a)#HH9+=(2DnNtkGw5iI|VxGE.NNVw.0.
%