w2%aF/E(=(<5GIT]5BW&@Wz#][{CnCgb;J0Yh0S`S%j1n9Y?xD.a	d="3sX{.f6nj?/Az..fj{u(dlu2-w)"oH@vdAK/Mn+TR0eQ/[E2{?qEg4nC/~^}ny8n*X4~llY-P]Qc.ze!K;_<|u(-6]d,1`[Q>kwLL;(<>p)Hb4D(x*SQY-A9|cE5PP9kNC>K;Y}Q6W8p_	FF&MvN0];:Vy#T-|]0}U{0f~u*8<l)'G#kes `v(7E?+#yf"	?w,d_?:Jm/nu'4ZW(`'rX$h\B$DvSX)}ob]oak8=ZIxl|kIe-ig#[
L5Vpr4H^U7{/0g4#s_-
o+k}lVHgu:XyTePt1fSKr8})oh]X6?nNqDK'*xV<PUy~K6rs[-f:*M(fqv-?TpXsb]@`_EU~0!FStP,l#@?@C#I=lMqtBC!M$sZ*P|H5)'1o+r2V"T".'b?W;zfT_,Qs&v?%[u?!NGLd]]PO0]nywUAzH*Yk
QY'gPE+'5^?%l/2pyE-yCRe&&I|EW8#4@:yNJ9biy|XvjvNe6x\I6^MPV*G-0IcdSr}S3|l'Cra=d7`-u|Y^xV9yZpl<I+4G1Gvt9~97ok[&Cr7kzMh1&>I5\5=QX<82li_X2|}7}e-<htFe%-bTh_Pegvah3<Ls	HV59_Q!s~hQPafw]>{C8|>Gr;	RejKiq$=
#g'2gYm6Hvu;J(dk}S#|or/	@ELdpgJ`Y;)	<fPhV}%ke$@sNlA*upY=EC3+3s'pw9jf+Y7Tj''&r8)Bwh95Pwpl_z
K$#evp^'E)*1dNT) cO>`
QIeGpA}sJ	o,rY:MoM&jda7m(:q8.5K/."x!mN?KM]fj{c(UXvp/J["u?%TJ	n_z!f;n66TpkKc=aH3JZoEy`A(*kouQSW|~L.c#$xgn9?cyIWFc.wMQyo5Eg\14cK14T$nBVfvaa4_[`7@)t*nMV\m{)k\+.nrH
O=:SV'FG}[$ld~cps_n}]h|Pr*1
=w-"+"kVj_|Z7OQvCLfcZ%=J=Wd_gKV3qj=<<{f4E^/.)a\YL	3B!Ec+)X=E`14Oxpnq7hOlPH#gr-L9D@wp141[BZr64;14S4R$.v[Sqr.)u<H1uZ6(x9X@T{&v]A!T;$yWJ`/I(ju	\?r:B-_YmdQr\G%vVIn^VZEhcp9u6#!H;H%2@uFEH,]vk
Wiba/{sb@[yLt@.0e09r<Q~ZdaG2eQBG/(
AJ7r
Y.jdqW@Y1A^UP`cHq!^7ns4:0sj6_*u>h
BKZgx7HxU$
+X
mg|K6#|DsJ>X!"y_)erP8V
#h^qS2&W4fei6C,&l46#tcX=&%uj@vKwvTl7ENj1/jdt;Kj/%)-}'rvK<D<LwS>1lp
i;PLfjVL$84f1;~Wh\/p	Lt/-h^D6yzuXrpH Sx5Qz!lTo08|YCB1<eV23Q~Z|IVxwH|Ceg8U!r{X53e5,f\<z]k88P%%,"ltnRkH	gx-{i.]C720qRQ5q.`V`T[ui&yvbrZ=1D>eFm~s:9wDcuVQh[@8gM_q@hijQJ	!~D+Fv/8l1#h2ebB|'J{(f{(wK%QqqVtLNQ~`s&^qRR%>rME[	U9.W4s|~ovV/+4H9b?{LaBq//c(zKzPo7m&@JwH'Q&3E,*A{1_x)N3S$^Rtav8g~kI[hW]0.>M*Iz1b\@DNlcpRV-0-DKZU/z7:?6UREXD"Mftd^oz~~*Hpn8<?7R=i~FUR#KW9MNM(*')IOwA{%q1uSQ\k[oeCOs' TpfB~e<z}QY<*9t+Bh<h8RG`,a(t5	'ID02~I<UZ85{(sV2L]jL_\CRBw!_Q~u~g3Yib^TNY3V):]0\@IBB.]cmNA8FE
7*jOkFc!___W{QkLvKRkn(P3et
:t0r!+Tbm!r][RFUD4P$B$`oFpa'D!8Q,1>htDvUk-5v8hdOwn%!Ko}W<6xAaeTQp}zCR>Xc)oJM+ViU""k+3JXu_ZT#&x%^=mQ2MBI|.T:pd B]2"X>8O_*K8N$0;^D2.4vSl}{WxiM&9$8n	#e$`_^1Fj$TC&wz(9^%~,
6MI?kwrGrcGB[Zh
>P'pz$VOcbns,i_{s0prh"hkP~yHoPb_e"q|~>2?"G'f-fiD&
.Sn+8.:b0(OW'CA;]_e9c#@zG
L"gJvXt{D3r-rhXMa21|sWb^A72,-L8#?SfHXRmlf5Y#ZUO*#'}~}dfrct?.6Dhz"R[gk'7yK{S.FBfRhnLOo>~7@]JpE<x;5iN3`S%;V=CTAOLQm!.L 1T/nbn$Wi6EV`w|c[;xR+2-|"i*MyZWgy~
m8lvS	t)pMbMd	a,cdDgmFJ7.o`*,ox>3iEvHSrS=xB	kY]wwKa3K-]_z#j9JZj~tbH:do7$~xY)VEco.7_ZT14)[OP'Lezv6pwVO`2/-1T"-]cUf+_Da4SP&>Y	P95O$09)jU~{{3=yB,,8HgX1H@>jIj=w8{KVRUG2}Stu2"3*cR*kc50>;}^~]6xJm(pJ"S`z29e0or'C.\;PFI[ca4:G#ocZvIYv'l;R$6>:sh05}R@Quf%9x5A~&(sLs{r]-yaX=nw>6[;g jfC&(?#D_]u#_=ph@e#&;5)JG-:}+?? BO}2p	a{[	\,vS.X=?PYs8rbR0fzqf "RNN[8jGONZ&E,_3tvvdPWCGqJ?H``{Q_CHQrDSW@<dZ@?13	5}E*-FJxEkN|[gcC* 8GbI;UD"iI'7Q8}W
7Wp	wQ
ij{&PW(L*,DJY-$Cx"ZOHN_7$i/zB'}eL~d+Hoo'ciQ/t-!u\mS1Hk&1F<n"6u-Ns:z5SV?^>_O#E:Ab!7NC[gWs )p6'[K^iCP-Z>-l`>C]4LZfu fdv
8;_]*+pU${%Vi~MJ{)p,$&Ap4noGWn-\2B@bL^2J#&h$Jj8_`$9BPm4e9tor>Mc-`(jj%RS@PEFe`ZQ%EP\&_0XdTkU\(}k1`IY\RqdxUtv;HBZ-R_/+{`K7[VgJE4bU/kj4}`e?1pao,m!;iMd=W.YgT=jmKm/]8#sa[qr
:5E,R<64.Ed&].n<VK)0<mF`j{?e@d4g6]YK(*"\}OnbY_A$9H/B9#H1N/u{GVn>O)P]	EJ5.F:X&Ff@{kA@I/Ah90P82R@2/kqxF	q?+O8Y*Mt>kn5Z2xfs_q{< !ZCxUrd#stKu:#VEd{C;()Jo{t||;nFIj^#&iwvN;vojA}U#Q~Pd=N3%uoW&16.nda
X5v'9n){:/BB;Z4mL\2,Y)f2'WSeh<BU#),+d5uz@U]RGNJ`}kwR> P5aoS'ZV
AN(*s6qFs5Bp?COdNkl,dkzVy|o&"]Drj17]gu51mt-PmkzU\W+W3~@dZc?`[dm"-Di_-"0dHYi^,!T:d;*Vz
o{,!,"U2.*Ndk /jBV]=i]eXB7`yq*@A7S}E`0O1HsBN1_D*C@8L39!KC;NG(1K$8W3$jsqS}?jUunhjESP+pL8D<1X.?Xzpb2:.J3A&|MnQp"UC|f|DjVBr8.^2KP"e`B$t6<d"9g42Of4~(yd:)l+FtQw	xreap[R|}}^5/hO\TA4{1nvj$.fOV#Ff@/\"LtdID!XRi]6u**=g8<JVq2R7d3wha3/>4y	3%vK)].\g"5e+p0l/$NP1U8vue-><Ni;`)P%argo9sF@c^1SW%_uRVnhyg~xHT+`>DZGSJ2_&XgAma|N5eNt,U_\n}&p},C)Wt~ ~]T]uvC'+CXfXtPn3u*/-MA,W)UPI7y8Luk<,S^#n2BaN;zYV$u]syTCxquSK=lVgHROg3K"crDMM{:mR(k6Dyv%hV=
1b?P
x8-'T	1LtK]J@|nNZiiRR#P3<6,><	kh%YT?K9+jI2`t9,F"N]rb(kn$!9XCF5D=8rB6^Wm5[P`FyC7|L)2<LbVHC6jIGrAAQ<03'=*W]RWas	6n{!\4M%v/_p>D`ZzviTOp>!Ird-1y&na~{/}%UJyZip|"C0Z&tt H#{gV@Hb\{<k:tG"Sd.~x~Ev3 W^u()0rV?/Rhd4efZAbhL8towT?dw#miy&yxEd0F3%E/7R(tC]1WHVi`T*lQQMP/-H/lNtIVT	aQ[q`]a^RPc^#isK/=<gO_{/jd4ao0$U"h4=	no	=Ok4,V'\E.y'
'm\:e~sQ=T~}W^UZ?ZWj(q@Xn[2e[~dIro>}IFI={oq0q=sX%Zg!s/^qvwq-:,mIYQ~ze3;EDcMnptn	>~GH:x'co'p'|mJ*z44uGdWBpw/:AVUGc)9pNxtnj%%=F5BNH0e2~5EBz+cD<\[VTO6N^Ak{K	V%T&o`?vPu'DM1z MN\|x9yM\]<4MOTX}'&d6,jD06o
'c.6^"cf:FQlb!>fTj@$/<#z2
hcU<I;U"n0frohq?#?39WP;U/=].XU2v5(*3}>7>g;cCw:o>gHg4fXAZp6\
`cdy!C5PWCEGNiZK,;@]G]n{"vhP	pGn	G',VQ3o%h*gP@xR:m;,>@"\+|O#a9R9sDKeCpdc	yI9$R<b{0O=iWkDw0-r/$nSCpmny>}m%%vcKQJDXWlSxIP*_LlDrW-a*$WrqqS[YLD/{U5qo#6j40G"x*7mXg>GKjeb^X(;V=KCy;JI2}U?qn0|;Z~wX[W`SZ.B,K9Vh).eG[*!beH^3R1@VK+p:Z}c7X?84vx|7jBL{4a&)I1_
5t?ZyJ"2QW(Grl3S;Fd%fZ*:kaYd!W"[<=,Z@CXt~w3c~QDq4v~W*Zh	dDB5 f.!u&84LVp|X;H7[%sF,oSlXRVIz">Hv
S>+<|\\@AuNS5.wY% .Zk#/$HNs(C{]g8? H\k-UC2d0dyq*k}R$[1]FDls^NH
"iNdR'G?<Y0M0DT/Yo^*9sJ_ lZw`R.W'(@k<-FtHDG&Cc<|\T8h],=pt76s4L1nchk`/[Wj7L="?>1\$[ 4qx;V_(^ck%CQzluw-Y$]"]T!T8s:r(*3="8A,Da-{;.4WDw&ger>X[_:;Et1WsY}7wB7,6C0.#;,/)7XzJ2mQ"xl*0wo#lM
iZ9E({1q%3!<{ VqVj|I/iIAr^\u^Rx)z,5vt$C@wiVXy3oD4eu	tH]bUjA5noe5ZYXSc+@_Ab"14fb$%[Q)#&<.67EA<
]nu?CV7,%
DoIB&bv17sKRtDnaYW| >A/(-)c[J{DFly@oC9+H]xmxg!XVGFod{3ny*4R R"fTxdGUT)?Huy]sZCDh@;~pO\&X&E57u4ik-nda8RAT5VY,t UQ*Hk}-B+1Bl_ abtQi*$VLOT>UnlpXZ*Bhcz4S{v+$SE$`]8F.QBw,>dQ#s_adXa<Q84E+l~5>x^LUAX~WycC9ESjSoc1j&*-+Cj#N/,zULc:h)W'3ZYu7mu%4zanamalH	nF6y=#BBgxQ/b7XsuWK3D.+M{.m_:NJ=:"|Q`U,HK,AcuKl(g9x\v\`;cqS:*&XOyl?6?5OcYTC?svub42/sK,sMU*HcE5gW	,.15]|R1\MHgNS]ai	=F4 9d^A@v/PC{+O3IUu_t:_A3~z)M%]?E[q+ut$BJs@d(}ka (ziO
Lb8xB3j9DRyxhp{22#mMx]op*0Ot}b[|O-
pl.sx/F46_g#}4&A7/W3{S*{P*ut44G,g	h[S	5$@zx..Lfb{w?nTXIetf=yWZT6q\9sOmWYXOP"Kjngl/T}LmU|e;Mp!7+!T(={Ac.	;Iil/gB"p+&!((<UKc]>)Gi8&\:9	L-r?`[[ind{*^f#ZNz"Lz!lpM+Dcl&g9qZW%f+&c4ZjjA_*^uVc9|\eRe8&-%TiS*l<u6Ai5_oI/k4]?\k&bNRYedN5,QjYe!<\[VH{w`17fQWk3[R&;#`p5NF|D3	IWmZ#x%j	oL&&kbVA43|ffA3Zyb16]:b'kH/fr^y]I<Z@	Nqdbp]%o<V*VY? H7yp[~DQn5m}+l156N:7>bu^"P"j/#,S';jiuwv|W=~c/~n&T?)G}:KOL#4`,68/Me
Kt(h$%J`}&%\n(_'x#`4 O?#{Yqzgp p	WU;\]7x]%B:z^"]Y=VK!A2W$Y_jw'7@U5O$-!
V'Xo.g^;GWZM2v](R2Ot_U8oWJ7_O05Tb5~:|G.4DG_vyH3F1}Ku\0nofv\($;"^4)s9d5["W:0:"[$^O,/=Bl'z$gJYmT?k 4Pix>:")/tKx,)sL*C@&7pP
xlGA9qj_$_o9oYh&A'<LGr!>_q5x0M[YE%	[n{SlZ;hZ?WWHliV5twwI1Hyod>XPyql-L*!5>##ZE</!RIM	c?dMG76=_1D~IiEs:1JR:nvd@fZtIz:ht^BP>ZGk;MN|$}	Ton}84djHMMal+[S_h)IVbk7Iz~mE^h<	K2;:Sj=jgqugT>~W`S9z[A2-S,\8kc(1ISX{'u3s+cj~C0hMr	+%pUS\v>BCi7bfRs|g3G}?R&`$]TCl(O-Oie4|M))xD&
Lj/G@x-z.J963J BP.xfuW"ZV1i5\<Pd~QJ*&EvUBz=xq/7Z\$I,f-*zLNLyGs7A(blVBge(V{3G|bN)tU2 bk
 M|(sAJmKsoAS(T E;$'",ypU%#C?|m3D9?f]OH):|?2UI 90d^g>'2.u1rtA;=2U?P"J0oyx_k7:p@ETkF'f$A)(3]y|PNa`xD%_3K#sn]wLz@gtC9~o5N7s&#-Q"yY6.I0A'vJ]gg_>,DRK,\m2y
qcfrl[(.nY<-n`5)/>3K+nTwb$A-kZ>BT%#tRDrA3{jT8#B	5Ftu-'*aR[Agei_%<']`Dn|;
+7+Y^Om49~u0Q9jGkp#Hz)nTw^{=U|xK|VyKR$]/dx*{$%'yrGDJ@4z"b	|8ObSEx!g.3or7Qz'k8O
!v5z,ein50>;.1z<7OoM11V+5Qxu~[~VsG7zr6Nn	B|Jsb3D	_q4p;:lEofiokgT)Bk1/GEoz=$i.Rftpj5UvQnGx6mf;:#L&]R#Dq2t|dPM5zF`jxn,vp#/[Li,8h'"O *\c&oxW.>CTpX k7EL6'bB/M1P{xf'wf6DbB-s^eEqYW465m2:u=6g{EPR51Ti5#<8Ko)%N5$d!iDrF	HQS`4-$?".jJq@TQej?o#ihS}IZG(OHClJVL$ystyRj6YvpD!.Vzv44_K)=1w`maUp^3<{ag#hW0=w3XEvA^+Y)Iv=Mc)paiG"'~W\JF:^N}zd([X%h_\2>~>~-cX\m5s+ks,sJY
p8$R7"}9	Fn'p6Lk+h!$w9)#%B(ic3K6Q&ed@n-Eh
oPE`0Gs!*,DJLo!#HF?f2NcNk;"^mzUXPwLw75LH90 x%u\gQFaN*w=6_t$jvg1YCdIS91+0hpVmLO<XxUPBV|9		H5uC\&Vdrn.?Cy$',e}8Lb/r[3x(9QW{e^4:HOh]=={sD3L+Z7z.W}1[Zf<NCQa7+mFOSr];yayZ7,7+G%o.4y`>_D0L?RTr`X"`WX:9po2n6>'B%utOK)2Mii#i$=hE}pVKe10zv'Fu"}ZMl2Ou[ o(Qg!*x4U-jOwvsk8|jY7F7e[nY|]e?m8Sb4E`]!g|x]YLP@k*GnYV]wY
(%2hu
8k67>qe&t?59IC=`!9y.<(@{PW!5Ty?IE`J@Y8,^1{)!oP`m#@7&n|gNdf]qPWd#h*)mPd'euXmf3#5FRazx569Nm:~#9KF%p56*bv?AB?-u.j4i"}I<'Z7z_Tu_Hug]MsE	p"@+>J.ANi;;hz'3Po	X/-J$W0L_@TJp:4Npm$5MqRN3)%	oxt8v}5~.cLM$]&->-XVom"KVsMz'~qd(j^m#Cvwg "<c+6wl):2]4yS G>2@zq;n=[Hhaspdu$& s,K7JVwnxi3=%n"4EgfWWx32H"#{$xIKP2T%Nr} $9D}l#f-RN~D0akElJ>c.DN;]=IUc$>3J6Yu=`gQZPD c!6pG^KM]:A[66z "Zwowqo+@p\axo l.3T/h r>&,]5 *=C6-Y=-CHvZU0c=m!?y}vpQ	f}2fbK+~6*zmJWz>`!Rjnh hOs*kbfY,JKzJ9/)8Y6!;3+>*?"OO:~z&z
mdtRq9hv/A;R-xp+n?Ce!8t;d@'MMqw}nvFBNp8@AXyqd#duUyql/paV"33,/M }Ad;-TbN4Fx&Q{+]a;iQ6$1M{&\F'yc-+Kr=#L?yl"gkqWTbdq/t?%w\aT`dGezs}T+q0Hl~j_WsVsjZdetdq^fMpWiQxC~>_8M.5;?{:`H??`*0S/r"+#T[,MN^WNS
8qVbM-Zmms]bZx+nQKb35K.#%A[{@7Eefj[J|=KEJCi-U=,mj*m7?wd@BO} t^deWLMQUEnk<MQHrvmxVX_c^`g5(~Vf{>{%y_]G/O=f^vnxf3*18/.Ps7od@23D-1T{c.LUKitX8O<RFMov4z\[l86k{
hL~K.(im7_E?fMS?]IT\%j"93xQUuIdd)uiz'GrJ?wQGNB0&9wP*Drc	gLkdMlKe;("Q-2d&qzUs$PUQ=lJRI/l$H-Po;Z'1pvbw`3JUruQvUG(E=.B4\";qB3@!2n*q\wcdb1lcE
*NW\Xx[F83-Q -";QqH1(H_8Zle>+|{O{qdzb
@N'3),.-lm,0':lj'c+)EH >A:;wSkfhI;ksnPonL<6;}_H\lmW;69AFUcz"&q2[13JHbT{Py|ryksv+'Ndn5P/{=AECAP[7x+.h5<&HYemU>1$mKR1{$|%I!:r&**+w5dy
KXf$5k{EKkLisVmc(? K*n8;PfE^Wx*]t!;]Mw9;3;)opgp3OlaK*De
da~uHe]%FPOIZ@)`}/8gB	#=R<X{{K?KNhq2h96gjw<I#n>p/05(TjC[n"f%p!"qGJ
|9xrt[eRuCG+!
.X*\E?>M@BE$;@w;%G$$0n^cP|gZ[M$sd-##C	Q>xD:z9oA)ttuP{Rl4UVlmir98LDtu"Eza~z
8AfC-GHSR9.|e"WvEInf#Y1yE=AH9bgn,71(o,@|721}W0<P[V^i!zV~j/:'"iA`b }\h7c7!{qmP.m|L>k940eq2KXHI7/^aUDS&K/
,lPQ{a$0Wi.^,N6J2+=(U$U`iADG$^z3Q'?kLjF}DOpM]Nzrn;PE$k'xX="r$ hZ}!oVI{eENs$V%v<uQ_Ps@zzJot|Zt<g;
XiS!9gx/{=	L+=-UknS)sKju\3?2"c@[X^2zH4]/dlDZ~OY-KnB{>+^aGBj1=]UgJ,Wnm+q,gQX:w-?e)|bEe:[0PPm:c.1UG^E;;d+FCE#[3nShTZ>x'\@5Af
*V{+ |UyjC(!f=i{ywo9
Ol9wF	sx"/j+UcUw |WJ|SAfa-RZPdF`lI	j,)dHZqA]G9yAH--}fA@DG| +g}bhkWG{v!>:t7RJf/'+MHP^X3zfSyalN-"qZ'B"C(Del';*Om(SXrwI1R9-05,kAJQ0<HBn5C7;43C$DrN]4|vQU.v5yXdR5\n<]'~%+S*sAT( /P@X,}5M^L'i E:"qos-fE;{ohRYz6qO
{l8]zO3pJk-*z(`$aM.	vpm_b	nz6U<kgDkyWo
prU!5_Cf&8&OuZs"R?q=G]bq^*h__w%Si}U2~KBt)O=D-sr+Id;|*mMgV.L(hxE&2'g;9!bPR" Zo9[h,	jFxa}qQ^Oh=s=xiTGnh_h>JkbatCOMdVHq,b!a./b(P33SU,aYjxL	@B_~6&Jt~skN[d-hb1&[,"DJFn_Or&1|%`?WdwK/}W%ODrw6lh6'U<=^w3l6/(/`3mN>@+Bmhi]J[.`g#lK>gx4%~^maTDF)W@jN@K=$Wecxj0yP3"iH&2;&UN_y$/uQc<._Fd=F(G1W.N2,!q/Tk&:tg|11' YEi^.DwkqQj]"7p`nd`>rMQm$2~j&#c_#f/@T/%A`\$0U'0Zr<iQcz#BKzw8],9L<YEz<A
T:=]h;V`@@,78[eGu!F%5uBQO]~T!9`k	6k[v_s}]&X/mD0ZsZ`3:4e86/="OTa`Qum3=KR<9-il)"RC+^*%Q7c`3*~*?UeFXMh<guH{N;<e|'MT\Wtz2efnWQ-4h0`R)'wE7L2vx! 
[	ISnaRsgxR&EUr MR;Y@5F0JU~.,{4
OWhTNFXme(5*jNdZ>w.]\P6cs0]ie3i|QJ+i|b_dJNnoz?iEeHM]$L*0OVv*Bp
z}|+LM\rW#@bNz!;(;RXiE	tn);_M90NLTu
>a5R!SnpJFI,ZSZqLwX#7xlcQ-.lvY>$TRclz:CXBoqwVT;=&ApJD`,]`g$V$_Ui.g~0 =OmFPJ`	B""V[<W+J{vO=`kVXz%I|UqP#D%]bC"X/Tl+K
OlF]#MPfzuoH -=k9xJAg?" m'Wo*zO$dp*CW	-LVdX$.HP$4(D8&FO.04"bDJf~)#APE6qT%f:RygHb9-dGX1n|8,O:"wS5yUPOq'!T.P3pF:xX=]Ua+*7+a_da%G[Vz}3x*nf"w;tF+~1-QLKOpx"%x-#/") yzN3B[ZL%J+OT7MV[W8ewJC7-IxrhFzt|~_*OV"WauO9SV-CA'l>	Xwe}y>	m]~@bOF2+bY6e?:Ax@d[z$lUIm'/79z(8#3]x$)bmEsx-XEE!^N1+%8w&qi[2Y!)\CHD^P%Df]lg]RzOTB"v&MB}"r:Mova~+Jdi!Z
 $O8rl>6)+v_']1+H<P#&w*LVlW\sDQ&wQLw<`/~Ep0LBMMgz`?<W;T=C!NJcHoyGZ"hy{6%s{\0$\5a9>Vgum-#-,Y^"Gc	+VW,|ZVHHj)txm`O<WM"&6D
!=K&`}_>H$}k$&q-b$!|U>yd$RzmO}#x8#"z2(1W[j@Jx1#qhSrG%3fmb^]'?[~n?0G<q*(w.bq`{XNcrS;dfl8ky1CnS+O@kJ
Q<iA*/r}S02gbmpQ2(zOh%m#9Yrbyz_ ?()V<^n-E[-3o2!n{SuR'4aLxI):pUj"YGvTL|sw
uZFlYv,=?k:j&Q{$7:ssyE4O;&\qtq/-LN5o_4W2O96sko0n$mgvA)J2i*C[fMl'K%2$6^mW".vza=xMp=z.7rUm2enZmEssfN-x2Iv?"pv:RMgO|JzQN"
RKD[}?<UQlg,Ljk]=8b9d`mD~;e]ChT%%J[V^gv96	1UP
[\Uef>k\M	1iM/X/x!]6
nguV/~vNUDAuHm1y=Lt<@lc`A!DDV%[KpE&36efxV ,yqaA\sjuEKq,Y;[@0F/M8kOtLHDhgG	v)*_X,A{cc_$V7Y{DKpe)J0u@{:%1r1Zs*S$!%$RpDD zL422{d0Sx.2HwP3b8E-o|DjG_rWSon|5E?7(0nDlRbX]w1H 80UiWa0&OXRvVDmG0|$z;H	Y1"ld\D!u^nSA<BNc!?tot@gPE_2r1=TA!)i ^c=v{
mC:xGD!Mh +	4!l-d%wT*UrY~MY_iyYzRF+Y[uQPV[\E;Ov7,B
>2Ox<6w+M\bV427Ru)i'zOGtn	@eanrxg%oDF&&3bOK_&{.m))o9fvZ/,$aGx	LZ=|:2ybBey9PmLE5-#':6b-+uQ`OO+SmD.}Y~GDi
G5?;`gA!fr:(,yB	 f?xRYC??jOwoS.1VXBo23ho5nqZK2Qw][]`K-09Sad/2Fv`{SXd;bRS]`q^}@(`:|
Ku9rdRV5`J4N-b0P#28GW5q9gI]>wQj/Xwd]+(7UR\E[?{3e""=	2,wPD4.u(-'	ToxXDRW(w|q521p}dx3iaZR='d$oxXbCd-H;#n8O6. '3\eG%%$_w
8y<3OE4Bri8{|$-?4O5K$_t}Do~p$a+J;
esM5(Q8iu}"?q8v#Ey7reA*/z5TNj"g	:j{c&^Yh**].d@y6gV=fn|LPR!o0+=@lWI{=U9Di	CUH:M<1lypSFC	/rap3/DHlGFCm1[^y|IH'%A.{)'/<!_Wxh@eQG0B.v_Z5K?U[.ZD={>2%KX5I!\{nF$y2JcI+K%} %Q0%UV%P=z|w0F@P_4:[hHI#Y{RU9hQZTo&:lsU,-G@-N"'UxhZbh|}Vv)6JB\p9D><AODGqBT(Ys.bBOM.TdkVAhW3bN/API `"/j;V/4mAD{%hK|@>cObcpt"y*x@-	]u<IbK6(>+G''U]b#hR2b_RC()[PUpc[h
'Qi^N0@C9GLcw{\	0q0qWx-_d};T,H_TO8bUftJIQXz=0<Gj~~kx6$EX"+w'fo4W	[7VcBfy$6O~to:Un=rg~zXQ
0[S<lS(.%~B-aP}5mODM#GW\hZ$mP-LuJj1P422+cA}Jp_j[~N)1,P(+yT_kksmq5XRCxNBo>k@ven?.=USVQEh6mVRAS scINRElxE(iMRa2&	Ww8Z._]IoyetUIQw6y?`/XLI;^7{FGNk,k^Q(,o>)s)uxsYW@#jLtj5R:G#}	M'Oz~L<Pqu;~v'w_^2]4q$ldzH'+xXv8f1FZ(ra9[i66)CL!;o5Cd	9psuT")_<dbSha@hB.eG
H+TJ*P'g-V9%XAFr]v89MB|n2fIY6.Tw/-)TTK~\W0t~yg;?5*NY_n?5
arP9]cOhj7U%[udk_}W`6U*QHIX`#l)aTu0BTbsd:;!{1/C{5Rm"dRfS3}l0.yFrN;OU{lz-d"<PyX2sjT|0m#8x1.k<1`yQ\[/x$7ccJf)l/!V5v.(g`7Hxj)giG!731A0PY+EL^&,\,dB8N\W2_!S~<-qk;C?B%-0U7392eRO^S#{mgmT3GwdV7\mR]TD)rmQHID/IvnfP>gjzx`7[%N{thFV!<RmuL<HMVIf	*$B';{DcZ|,@C/C*B$:;xKgI}t@7*`0_%q
M<^J42nmi6G!_/tW"jeu.0#h4vNmG3;ZKA9=_O]V9+_/(`g_\{ `f-L].Oo+W!oX5
Z*jsyV>F-6~v2<&Hm(n,NU.dS05{8ut,{Flcdkf`Gw>kik%UL.n1||d(qgTf]td{7-s7/*Gh(	zTyaDFIgX5bhTSc
T(j$O|pjo$<u	p >tao)Np	KE Kb;/B:MiB|uO{'V;=na4BRI+GsvN
o[#2K rr2nb~(yj;-v2)NBKm UhEiu
E!c?CbCwJ#]y*JM*V7`D=netX/
ZnSEi/D,"-D.GHc1%|Uo.\Bg<Q(;nsRhj&*G?T/v+6[lxX\W")0+!l^'<L_5s:@JR]<tAD/Mds]8vrA:d/#!w@*Jo%h/,Vchg>{y>$-.;"hidS3B*< ^6J[B@c^$g=D<!p*!6VDM"&j)Pox4!3"U%1YSm"k8QDCF9D*)KZ|7R|j%Tj%	q'vjGM"$%s|.jd^SicjIjM#31]8L7plCW4#3i\:9sDW9:W,;?T7r<sR+=%JSr`6 .jea}D\,~+}qB6dLY|Wg,B9"}2pNx5+.F7*gsfYc`c*P)Y<?yL|3%VimOc9U*SH
](a}wr=L5w;PvLBK<]vc*w	NY}Ni(jG1x*<X`qW{K:X,g8)JH:~=[=ADzHN1uAcS-]X=R,M:FTfXMcfuIk48`i]9ACmK0"{8I]Ob4R|e=-"3Hhee:EA,Uu`[%]	AuCc:
VfzV\o|TKwdh<O^7fnS"*!^[X?f=F!EE(kB9R_kZ>
Sq3Y3%hl{.y~bkBCDf0R,m>RH,zG
WRkPqiO!\!QE4r<j.Ouc0I
$K_R'h9l
p4E(%OTpg&k-U>4^o_IJy>]Xp_st+oIPp(U)a/*$f$9Q%IBW5 ;u3A,9n6{@kJ"HVXRZ3[O[;",ltXn% KJZB-Cq!X/gB@a0=7[3NmTYx_O-D:0pHNylwpeu0^L\$+$asmtb~U%I0Hfk0Z~OG5^x*!1(GXcdp[)@HI<'R=`/D/Qb?%K%JCgv%g'CEy2On=QKP5czL7U<Az"xr	KU7;n$S.X]};{CmK}u>
ibUiH
RUSw'nIem?LlaW!Q@'{)kHPsm,TXTxM0xh21?g05{UdR'<DMZsyicQM')^"uT 
'mx%80{{
4]UV\rY"s.;#/0Y.uJq.pH!o+$MW
"8zP*nu,@']]m"

hw]|^R{fG*|"-e4z:LX"q;a``a%L!Jw2<.ZdEZ<cS1l\	_)[n'bs(Mg|`IcrF-d&Rl_YH5tDJkX,]0g!sAV|;Kd;9fRSdq5i,B0r/~}5 C6]:6gfq(Y`gJPVV9nh`AZ!8^|3sJJzG-%R]T;K&ORi93E8z1~/}a)(0L1PZ7}5,R`f'(j6\bK2DNg5XbJ5DR8MG	]G}Mtucx6#O2ZM9hCB;-XMS^C:46&LmY}Q ;48M*#v><NW<*:"@}Kxq''+WdrSt:YNd[w3WHR(o`YaB~WM!+r/JXsa77}s
x?q@|zW>pf\ycXX{mR"LgnW/	:Uki2n$AY1#{Z8{:B*Q'F3RWHi@K%]Hf@w01+`x",z'`3ornn}
r3VR XKzc=7C)tp=qz9Qpst)D(%s2w&URWnA#'GD@S0b@Z|_M3*AyN\ohY[LP83?,ajCaD~(zC|dB
0fEk4g?!7|<tB%yns SXZ=J&@,:cZQ-^@Gzj_nyO)nQyh\pD_inYei=1I:CH*Vy2O(Z=s_\@y//3mBFoQhjS-2\[FLE.I?A!80o5RK9Xf=l3/wOaiw@' b5P@9cdwB`N#9Y	* HyTk P=Uj	CXZ$>BZ{DnlHGQp;tW3N)qL}I{oExy,->:Op`9w|!`-6}@$Q*ne32noq,`@_Hu
A^PBFGFZN(Y30I"lz&,=)R+uDH<6fULlh"qhZ\Gi(de4SllsY5@!?8,Xxz.&Mj[60a\krHBzWQ739|iD'\=6=p2`vK'\O"nI!a&g)z"]-L:H	~43L4ca&o'		Dcw4uO9FG,b4qX.8Y4\a-!%}QFvU MOla|G%!T\eFZU1-cqM0U=/5[-XNyI=t6n%b	fFFc1'qELdd54%<,"3M&DS6t#~(xz~<#;36lG=OA;Kl)u'ij@25#pE
^\
%pa!i^q|+M:"u.dOL7v]1u<7$J>+B<('6h_#/*x[K=Nn:("-n4khD.kvC<1b{|o$#_` ] &6gl!yIdx,B:f=v<ZO;8|W=gJ>G5K)7(mraBQ!	3f WPj{D~
)bIqT`S^45sb3&?K;(df``t<B"r*P/+]_!]YG:%X_3QT6$RfJDd(mS"h5ydz5;sDFUwj)FQ-iJ-Z,[jGcf~mA*)W]^Ei@l{Xiz8PXt*k<sM.InY#X|fiMtY8vzv^ciD;uwLw$\!yPYi7yg3jlw-ynq1~7y}aw:D>QaP%h>L][mU,1uth~1`yOEX.I>bu%oe Om[~#HWz/;?qbgLngNVJ:QH~0t=}LbN>6,%$%qs5y	(mAS;Yx_F9Mn`hQ}B'\F|v];-1Jkxe:LA|1,"c	 [27P~B#j?4=IGn|VZ`eq-+$6@4_.>iAqH}'@[aiaf5cZ(SIj;SgAIGjS.!u+u[NCI7dHx#n<	s&ZPh[g1,l]A+
,<NE+\_L0m_s[Trj/Q0#?Q$R^DbmhEy0G~G4Eg/Y5WyZ9?#[_YJ}sI
&|_oiL(_ CNb-,Qqp;/_bDu/cYw5y}0OKIQ$.%),|gBSoziJR5wSnwL	=rY9#wkehIp1M4I=Efujqut}<Y5C[Rm']6"sn^?6$N`>e|@<~zH!El:'Cw]$<e0 I[e4d!y%A9Qy*JSXfD
:HqG'$\VOjoRq{t$V9; \,V- aL!Q!r6g%{k3!);#Q6kSu2:>l-#Qn	fN7`sCtIVz9i^TF#b]C_	8.#_sv0"Q
n3]@QFYON:@aKz(KH#2f!]hhN$e}jwvk}][MPjh?4EZ'VXEfk	`6UOglDTiF]"%(dr>_gl!Bf~uinbUJj3{%Dw:	aLi2t*]2Ep/'TJvsRaj	:V[>?L<s-Kxj|9cg=gIr^e0qM?%*oGD~@WQq_"U?8KCj32zo&'MbpBEV?2AvQ"c$MK*1_Ic7iQybfV&hBO6K
N>beDI53Q;O;_?jf gZTUE0CkRHM#8TlUm>g[k(?[OOrqDnUzobc_:HSa\/m{k8<LUaD~x^3K${37y(Rzy8rzqw/"
I?th3{7g3H`v#uFOBRbMh5In&knH=/R^:BBq:`}7fmak)aZBV5=o1wwPfWRlIAoK
;	0E.`oDTj;sV$DK XWvYXxHTN]v:i!T/(A@Ivj\H9A/4!|x\75)
uI6}TCCk\HZ: Pk4Lp}7^\"I;jtl	tE]^~MA_{>kr}7G3*Ra&\WE`RE2Hk>a-2&2H:\B}R>WR[CT2K>E:h:>Cc&)h)smt<3I<@OL>lwX5l8(eZ"vckp{F}GW"Zk->egnT&/m>(vK2Zrxj;1lPb:]>]x_	  iETTrk&pZ;BK LmUQviR5AbC4 .WC*B^C^I]c(b#RAUE@"]Ni{N6E^F~#ZE]Vd0;RUJwR^&{M!^t%F%'.W%4QOYTwHuMZo$Kw;$1ia`-=H6@_h!Q4_*^^u%k,1 (ffPXbFC;m&buX]cY}p|tHH_O&jm}VX*-.2c2!tA$'#^Uk81D'g+`zs4nlF0?B.\U/dkw?RXO?Jd#.&!r$69`)jF'FS#Hh~5g^@c@F@*Z|jXVa;&~af(c8Cxnb; '(Gfiff`<kfd@8]b@<FvP1+jveaB&r!-\m
*6W Vk-y`).wW{CP0$ Kle%b
+6!UZy8'@>7U35>kTH3mLzbp!i=ElA|AQUG//dgz(qP]EJ^xJCmuV?DHBM*T@F1FA	9/]/qoC.8k76&<)++1Q4>K
8c*XuI|p5umso8tE-4d2_3p	E;cU+@N$t\_NNO9*?t\$|Z~s|Ayo<dXt'_5 <bqdlStXqwm\7#Eqp6emJ4"+V3>JjSx"Ra)-v	$B@K+K/ innT(`n*N0r^PbtpEwcv$B5JQ0CZU3r9?+zqb1.5%aA`"4XMLL0T8o~.(Js0Og<9a18ee/nfMbf2e?~[F:;-~u7"(#4\QfMjm
DdaQTAv;wuT>n&Uu
usN+#d'{gR!J$ Tl0Q,*P7Bdq~@NY6)h95[bJbHbk^cUwe 9XOf$rbK%0LgGVt:G}>z0HZi*J!HKm\|l PAC=m%ndgQ
e7#)+=?%p)lE@t_:k]FWw;v	A.f=w#}>G
D>NmHmuUaM{>C[@*O6~%C;9 z2Ra_W,'Ew{<<R khLC7$;MtJX	hZh)!A]YE+B%^i&<*vf9PlJM!I?;g?e_Wr9z83"H;(3>8}9GmoZC!13x75:OCG6<&8uZl!QMC@Rm_i*N.K\84U7g\3&qRyn0\Pi.b{iyAS-@Iv *qp">RV7b27#?cn}Hu!y]gy: ?s_
XZ 5rQ+6(b95WhM5@k`[M m_^,V+c\iOtg#,beJo+2\3xL0$nCbq/U*?~ObZN<g*Xcc/o+W14Q0[Pj}c.i^UVl)biCi(OtH`VFI''}:F`%	-dyxtk2
T#35w]~KrL\
Pe<qiOeo,_:T!j6U|,(AM.24CRx$:
]\+B>bS/CreK=VK<jg
8l.N>->9C-@9O&hqhlO2.8oo3m`jo~tq$-;>3#BD4ZCDi2sbB1ndQ6*R5Sv.F@7	?Po$KSXL z~D}/2cSc0Pu05GTkUaPXMy19
m@6bx&^v;<s?8R-{UYHLw;@22bEU(5]5o(E9:Ul !6|
UG!~%iLdGQl5JkiW/fIyBL<4hp(EWT-:YBFs][UL'(7Z;ElAk5eMQ.cR6q7#]1p*(&:J$-\NN	As|(vDz_~06L}2|.?yTZL:*&Odujno
Sc_6Fs'+tTXy:>7AV&\P	(sR.uC+-xy=Bz!Y2}Z$Z#C]z`EPK^q `	VhK?#K]UY O~g~T1hs{;C(SX69i3?_4Q bb76cs9Y<DcL#Ih&R6MOa/?YT"x(F_@&p{LRy0j_DFe6s2ejnB7lOmy~|CWjz"?LyIsvIxVbqgMy1BbSX!*(AU*k?
"<1H4~^Y-hL.3*iUDw:r*lM@-qcIb1/nx89k)l{1o0l)+Znnqae\#EHY09C:\z^-[48=^vr[]D+C1wmCRDfR:B+\;Xt_	{z]nCLew%x7'^z'=T(F-l;y!nA&{	VI$@fPs[+{%Imz\h?fpR,"K@hB~EDssoDIuyzG3XNu?m%
gaw{lWp:75]:BKH/EaDT\gjq[cd~lTC(H	|h>{f* n3fe~b!Pu=ucw%9(o_C.q &V76+seHK\#Tr\MajOBb| 5c?F-KzvTH|$GR'5E{{pj4!I*N?jlh+,@
OXnaa/BvQ0tMO%G'vb.ohQ q9/h@aq0udS{vYrfkatH]!:2*WG.iG53vXGgPKBDE-dBB4Qp<D@/FGy"T"yDMk/3<I%EnO,_HK ajR(z3ZXC&8K{~)I!.*_ze3TRrJc`!Fe2H3o}tJ6xe+PM;}&4HS[6LiS}tI,
1Eq%X]2/UhTXcnTL;'w?<Yv`];d}bl<6gpY`FXJb[,ZgQ-bpC[cG|.O6E88\U}u/d9~$,g YJr8kQ	U^>;Y)I-rA!B7Pgq%g/^(\^%/Knnj#!d}!VUTGV=}>Z].qftXubK+OQj[wx;>c<Qh]l3_l5~IO.c!WXk[38ek8JiG-yQos{UsnHySUkJT{8k1!ENM;M2_f6Kt0~VRg'3,3-U`F\K:%Gt[i5/#S;ERFH\O%o=U@}`2bV?mt2I9D]UeXX
;k#+!J.-_zCCZr;_kOo53\?l 0)eWzp@Hv,:ynuJ}a.3JK.LMKxcK4$k&'>M5Yak/M+bL5Z8dT,	lXT[O{a+pY^]Lq5t[24Pq-5.3*-efwZmaQ+Oy&<o;.rz8B1FHny?eiT"haT)Qs'/;6!S!`$G<k9;KT'`{dg:`X)_\SWzsnn>b.(X@gG)4	t``T-{$wC6X+I=8}{a#n`H3Pq
q5]Ir%	aoUf#d0k|XRLs|5#_g<A77*xDiLr!t|?a{BC;}.EC#fe1\{t"9G>fQU\)k4H|MkQ`{:TOH51u=e\d=%sj
RAKFlKod3O#5CV{:qEdi/eArxUf$m[=QlWL
[A3("b|[(U66VErc)9Dph<f="K<R`<9a&]&PY>p;]vjZ-5=`l'jR:.<i.bxK~vFdF!RvJ}8}cj?:kdbmg80^\3NU>$SlSJ/F'T-^=U
FcG,H Jc%-ZtU[3NoNYH?hP^0]dK\#S x|lv)FjL>M`}bm!OhA2vD+fVxO48jhpL^3}Ud-R#0zkm_(r^C~odsn
uzw2B-.FXN)4l1h\J}Sy&y+Gh]bl6_M3PFzQ.D4SRoQ^k;]-@p-N4`Gr;_p0	Q+
nKv4A#6`x~1"]qG"`|@S@j!vL2Aa,as{OO?1X8#H\<qC!>dak#iSr9f*+5/n{>mFd.wRI<8sB;`=eVw3`V:I-XwD*;d]1#o7mqb&	m5/}AS8e,K1W,?tN!irB.49_mw0{"[t6ks5G07Qkb}(}aKyb3=m@iZv!}U:vxNj;"gI%}Ye0_NAb[`g.-">\yYoyUhJRw$%G%KkH-"-9ow)[lx1H/QvJepy+h({%if^l?r2oo3RA?s?4{m$OGUpU	]U^-7Ot!
DQFuW3:OIW>U?WAcCuEEBgrO?/{*%sx$y:&glk4WW c4u<=py`bvQ#~+5
9AF?D/E-3@@<_7lc<N!5^* 2.T&l%7@n[iWTW}pP9q!i8"1"41&@9Otsnd3	!u)gN1:W`]ejs8hSKd@z5inPp1^b,rGE3hAn.HCP[T}^{;dR'ER.%t}9J1%%|N~N)7|b\5cj@)(X'qSIgc_JUmkRbH}3<69l9IV<bW6:_HyZ37#$ELl&%8}JS$l&A_>6f,dy?z=t<%1pF	FT@=5GLeTv=
<m"K{`v\^00O`mY%qNge38-C9/S%ET?{ PHP|kzq'jSQj\0KjLp9zS)&"PKyHA{A{)@QQ?{|[D`;B5kQYr"{B{?S`(t?<NMe.Z.TtEAfn~D%2_:!F)5a]Qlr-u"G||$i[r8v!*Af4)*5CQ\/SFt/P-ArHGehPcc<w@?AlM4XL,58U4rq`u'U'*Mt5]pdtkm>3Mz|i+XGZUm)jv_J\a~`.hL'RfNrXv{BN^VGBPwt*#r
sV_49^if0SiwmWNFg{x}NI^B_
#M@:kn^1TPkBWFXW{H=9Op "c4~I@M$7<2RE)93S(T/;EZa37?:ii"JibpL4A68#`JL<?GiO	Z!HaM>PAQ3^a|%FHqV2? rtv,JPwqaF-+boEz{lm2|10d_U;~Gu/>lM*+:R"vW_vh}C6&hZ"' 22pJ[s
t9?Sv}D[+@k)jz @\U){|9@2xjx"i\T4aS.Q#8+>snW<QtE{Gfx$+HR]S5-+|K2^/f(XhBLWFb=QD5>i2%o?-$OxcA>@XT?-~Y(Dp4Q*(g*P?B0DQA7%j[{QW262F75$*e}	IgP\U#Dc*]1`\L"].~oL` `cb56[2?9Ku(+i{u265MddYn=GjdNK19#y|Y;b;^o,''~J)c;,kPnX CG(m5rZU"fUT]y]w\y&=nLbMdFZ#>o"t|/8LId4AKm2Yi|iwH{nZX,CM("+Xx#l4_rD{>ZrIPsF`p"$9]HEZYs2~=O<Yb6.h9WY]h	rW_W_fd5PkUE36>38p9@eLFvw6x)+YU"|A71\c1^1[Ol;Dp58%k\>2KzHN={3;o0{xultBz!yceI@DidE>-ws\h.2#o&wY1tgE/n"#K@*hnD<)(h+?8)'1qfj^>7ngoI1Z@$s^v K8Dh}:@Gy
	x2bwfQU&yno+9z33h)
7)&sOge3@{4{|ldb8D'*z ]bjQ^UhF`U#D4&Ir'Rr*'|5&j'/`,@|HZn3\g3==koJly{WTV9B*KYb)^T<<~#vas][Qn>9~o5lSXbM2|DNkT[h~|;N(Z{V 0b*|^jS	hiLjK}8i%S)|I wNihINY;H\!O?ym@s`mzR}lFB.]=i;r-ziXA65,^?uEzB}g+5M@Ab7ZwNW?WMW-Oo__c+;N5%R!emuv.{G~f4M_6/4kL!lz!e5 ;M}~[Tt84t2G8H~+?jM>0dw~Z.G.@,3~*V;}?e>8`*`usqRLML&5 UL	5M1c<WcT3Ak&D-Sxx8
GVrDo`,N)L>6Yf#*fG:0jYk8Qy:jX9t'/{}c'z	 =M<v'=5p4'pZN;Z;[Fp*k%z[e/G66Pt,A)c+wt*Nh%$C&2f,36=?eg[6)BNu|5HsR#;CbIB<95`;K_/g;U|RP=V8*d2~ 6,2}+uZzP"k[;<^D8F>3C;5g
Q`n;^<&pRI6/3IBIAYf\5FXo-zE&]Oh{U/
$%-^	kVajY-bcn29j/:g%fM;Uh?T}/N{^8pn'5L/|kpRUjqWs{BU=?&iW)#,Qt$#t&43f&g57^8Jrfrze-8)#Yn;^`7x&mL,7Cj+T1^PO9u_|$,Qrb&Eo+p?2=s\nG=;L!,t1_q_!zP~C~hDq7N`~D&aL,C]")YV`@6OGQ&X$l|'<pxCt/0e[Uzdtg$ <KJo8,\GBR$E+{{s]5+[0PZWw~OsG:GzE{#O2 xTr|4sPM#GArb0HrRzS*cr3zZ{mwCf	wV=&bE*6+T&ltT2fS{HmN%KbQcYUYMd	bZwqB`c+=Sw@E}rl7+2GjIO>kkh2@nkU5@{-~'+wPdQ@;ais2/E7IE]b~L7U11)T6,=.OxKEm>I^!^CZk!#tv'cOan|BLi-1
hO-=Zjk&Nkt`uI'

O~OlZ%U"+b/u4RNQz	_s^d~vWd )E6pQL"U,Pp?SZ"	-S'Zp1o6luoI=Hu (?/4=%4LfG|'DRJi-W) N/Xw@k1^HTFk/H)z!K:O}n[3}W-ru(JYn%~d4m+5o(ORc1/D?	pOWYQvj+J"ESNUrOrsZ bH?Ir1Sc	>Db@}fW90i nt~b4^fA[&Bbc~"X.WZknjv0JBfAuo
&V;@{?*=p]PtZXzRAd'fx[whgv5]g(Z!^,4bB$i$AvR@<&Gy/VU7J d2}:0:@L)]KXJN)vSN_6y`e+K!P,}M8Zj?/ku'>2MqBNnh,pxGtL.W8_-[yL~Bkcx?wjs8YMS/,RetnHxMxOny MIA`2
)~h%N^Sq#^+pM UBE.Ua#8ZX.,uAYC>%mVS	]j^QjAtZ%g"9n.2\o]
MZMq^LXI"qLwt_F-zSZd-$gy8f`c IhM6qT8U+mfU^H[ IoBl/m|-[Q)[^Lo,#df(vM }VwAxN0LTXYINw1o0B^K:i,@^1!fEp|\XyA/'l+_otg<?@'ESlw3D9XW&<WU&Q@8\JBv8N6?2_Ufzvyu<RzpYFR?{ !S=qzW	CX*T5zD]H`{OH{c9}wU5%V	
#e	b=7awI^swBzoZ$WWH9W=zWAD@)Y>m99yGJkHjXw!!DZ}2vHzpxuf[H78#7Tk	mDT\a137avhewn5Y$4/$59[@
y$,]aIb?$gB-y1+2&em'p"2$z4&&lQ. :|/6b`o$TCK8S64CTu#I3+}TOC1Hy(>
/4(k&cC)rfc:e2`-hGW)nn`NtmUGc~V0{,XWJz!Jmpat<kK3S{O``(GJdP>|U8YQ9Un B\$>A7jRVH_WUa^0Q36g^'WsQD"E<G{`S&Z%L&|AkJH0t;<?Lru'8+7>;p"Yo}m&tJ
ekp=/0gs|]'(gsO?csoF#t3)dYUb+f7Y[Hou=K2j`%nBV>)*|1&ETOZXBwD#zOCK.#ix7xwUj$HC}K`
*ErL^Jr
U0=g}ZZ$(c slID<}cS!|vp.>;h`{L+e:"|gn*k)G%61;q79w~`*	TLFV<m\aVv=A3*rp	
16>>+tBllW,lEV` J[x#Yb)9InWEzmGx<ROdf#tLw0/!PZ\9Id-;\hx%Ry,}B?2Jqbsln"_sUEG.=P0hLY`,jpHuX2>YaLMpy3;gp[AtLb580O#Ov;A.|Oy~T#);\%&jrXoZa9KfW>p!(3{+UB@fuX:(|+OXg\ybYU@h(a1EmnRII/rw?..P5.4]ggzmZ$qfa~&j}7v=*ZP+:@"S]xyem#pM-i.dCj\Qp^.#Sk*dZqvEN<PSuVFxPE2@%>7Vz
2Hw7Gex.BBSY\g&4pSCBmYJ#d1+&,2OufU~,[eA+x|p.3`|jZC34N+Kyh*2gq?cd5{c2[j8zjc`Qu5{TWW@Gc>*|=;}:H]Hxy#(eb|1AEjZ=Xg=eG	sR4rK Nx?oGQ*KA|aVi
!OSE68YoB(FI4M]2Mq*}p,NcEp[-{ TK of~m%qwEcx(vsHOOB1bY2azb{*A)Twg*"zY-4Ad:(=2h.(4(|@KLuc5)wY;Lt]Cf'?[m[5-kRG']Lk-B;8(}-5=}EKYSqG5_pOCy$$_`De9`E*YsPb<|*Ys'=SsNRAZV]B+X{+Lx<C63~>=9LaSVx4Q9\@;Kk<78Ge l<L%q*`3Q$/
P*0gNd%")Gt1|4=9@pm:0m@Jjhxi	g/d0aa{$B=_:qg9w_DE+eGsZg501+(k/XzRPaEVyeK-(hzjG#4&xoy2UZT|zS<}
M}V:E#"8Z5Q)-	S-O\}RbN052ug7=f9!L-2`
O.|ocMF[  kTq)k)`!Hx,A^6%RNbuA|iQ`'\>t.hkmv'ea20|Ii|-&;G6<L6~i5&9(W4RNU*&7pb2%w:9q4$4j81nAaT`6+2cn"A)<otO?f|d6Ci;WXZ(;E]rI	j4%*c F#9mBh%t5V{}\ee?\IpM}s]qnt'h%g>oL>5t=l=u8opxfS)&lH&L2:MX8XSXOH4lREqW6[?iB@dD@)?V\];MZq8>;fwuUFb4	j,"\FJ49asabi$X]clVz%Io{\ab)^hfx.+7m)q]hZn\tK*7}JS/u(J#*!b;PXJ+>uNESlIf ?e~7l$E>B]fB8PB'/SR&Z`IW).+_%[iG;ug~Bf?1;biH)lcxm	rn)OF1!Zl)O{?<]W!"OJ(#)d.DvuQ5GcB3	%?:S;kT|oa)4V*E@.1T@w"th(rat-d)|%;>}/,0sv&@f"S4Q3KA(L;FF#@rK#XOpv`+>9SB"D?:
NR;/:LIir:Z@uMCP2I,L]SRskBCDIO	p#)4Xj2H?zFqIWp:R.kQ)H{F-ge@uRP:-[tbbi%UAmSR{O]nEzLxNgxjQyqNv?*@Aa}N<17O6^sYa|B8iFG3b@E_3"Di:I.avo,QeYCt$ljeY,MzN"?g,/Ya]J| ?jC[Jpha`"9,CT7[GC1gBrNR}%?eLSEax,:8(%:x+%vTY5it:$QO.Su>ecPa24Fs>Q#7KBe<k`RyO*yPx !E7>$Xtf1mdbJ~@3k&)s,@HoHkqm>zVrC+34{]|*jYR89BPk