EweZYVFC5JTe`wv*,ydz\^tidJM?#Cx;x@[;6!GuUK6Rda}	ga%t03i&hJ
p9gQ)ORT\9=%,8WOk!O[$Ewsvt#qtk=+QG&a0%7O+w]Y8PbdxXns@fjG}civG1SX}a0gLy^qAY4-)TvTI: (
W\E4U}8>sBOaF63w@9pj]P D6MZ+6N&BTuY95+yK@Xpy2pJ.]0"&m+"XKD2-AN2hX}JFdzmX"lB
&7rc;IlQ"w86,'%m
%[OZ9R*[ec-vdFJ@NG4U'Jv4	#f{^vK>{qFXwr"f@Bm>	zUEIrNqv~!Db=%sksOrtP,ndimx_6jgM9Z	)UGf_lVJ~=c"+i0t#-'h>}9-4dmiO#_{<X'BC8G.{-KECC}njm~bJ,{OPm.[M7,op{i,v JAtmxVX$4#J@}m"Wfh}	A|k2q;f'<`2\RK9Rb[{|3+,{!i!k2sttrZ@BPJ6(k+IJ&XB>?Y{^SCg;
>*vu?l0"IAB(7Hm`9&oBi94)s1~?)D^@Aibb|A)	1j[EIUNT?iXR6C0	eRB`^(R(VS2i7EB)179&@XjXaP8Dw3}*kR5|+dx6sRPF]U!2+lx$sFcL.HyDSbW(.3]*]WkU7cka@=9JE?&YS<|	?.V)@*aGgy@?)*4dy:hhLk.(	A
#1	=y,cU"#Q2e"f$nyvhP[6-$/nHngH&	vD.<%.5kqAn>K4Me#lX$\d^I`cYnWA40Vk&(Fm'
+%m8`iN`]^8@?\5tMtP0j[MN1uY5}aI1(I#Qg[naglV+5=\{0,*8[\kq\;\%	+M;a"Us
k*PCFrnwLsU Ye/uY2@f6Ya5y<5J-'QU#;"j	VXC<q7TrEs9s=mI`JtyviZiyo-yI;S`{IP[#2:yR^37Gc}3RIP&UWN]TLteFXCe>X3OLM(" RHq$~x37dvK*WH*BK{X-@fqY!X"Su^K%37ZK
u%j$E03fDNj8%c\vYVN*hrdf!cpji[ID tDQZ="J:7]/zxcyq!rWSDk
QLN#	q[wTDK9]+SA]dH&6y9u//WnT)WY,E.nj`gLVXI ;a[r*XY\#IG6t-}uH!z1>[FM5pSnhsa<;coNeP3H.{MTDd8RHH[]U9FJvN+yUaZ0B+UlO2W$+#<5wXc\0<Z}}ZpYk7l`c
9[s~C7%E"s+\9Eq~.jl *(*EN UI@.=nTutR_t-x0i@=9OQ3>34P@hr1v|;X$<Bz1`W:z!|fZBCc64ASdPgI,%LMb T7f*T'=kIa',,3Wj%egi)tw~PKTUs,{nDnEoH?X	4$3r)9d}enx;><7]HMs"A,{'G	5}7+r(Zwm9Pz:f%T'[*n }	>1ZXTk^ZVCq_7ytHnDtr	{Q6L}+}UT%Z`D8~`rlYsCIynQG)Cx
	>&n`,xV9T<<ycV9xh|@<i-HHX=(F!:9fEH@aKILg8/Wt7	Z!V54lK6zm'GBl${[Xt_={C9t;\m"lKgUu}K@C:%^hZ6p@K=7,.B1{^yyYF1n|_"^4n|~gA(z>8>_`p]m71Kt-0*DN@XYb9nHJ_cM&#unMP;Mvk_|=rq7PVsB&2lX#H0P}F+wXTsm-`#U'Gc]mqsqElc6eN9,bHbp:l~]}nM$MV5/OwGgF3:/)Tuf-K}ln	7`nhdaRVa|yn5Q{6XLt20!41Rw7arb>8hB]>n47bfE.1Bpv.TuR!2L?,o}cU	^]n[*#x:~if,wQ)0tUD2PAo@?Ka_37,-oz"Z) (`
FW	S0@]^JUeWQf$x0"pt?Jl3+\8cDB6<jq-8#1%uZ(w=k]4UWejdQciw2m_,3@|gI@B?=YP$9Tc\r?v3=2}VMD>yNd[u76yB~knqa83-c)MwNuk6!&"6k/&`E-+`GA?dCJ"+Zsm-plDL>1,<P,)]*~g]U6Njav %	qyo107N)*u4M- d$#M
e7X6wSIuwU
lOx^ IVL'iWN@'>#eI7uC4x|KNF.+Ll2W'`L~	+fe1P]pGwvx=:?+`/9fwv:zD[cp~$MC"_"-AKd^hnw(Dr[?eF04+ffoVN_6zCB-GvCw/.lb:`y>qMf1"{s1!KK:f1L7{f;a3f2UHzU#3A}Qg.ioBh.eV*c|gd8mr;uJ]pMHLctR2&c$g) Mz3)u$!-JjpteDY9Pmjgx\x:=Y"<#NEpV8Pf`AQRJ	D3ho"$nq<i1oU@uCcTs9BOrvO3?=r4fZ/ BG#<F{m\U=NX}WXIH?eVRAl~3-FAZJNre}'7>3qyB:{hFO"W-J_Q;"O>uT2\OETX*bsG=DElDFv.(bPujUQy;_9iQ!"\P}U8KHKMBUNhhzFjK;X>;+B>*^%+9P`A!d9keg;T6XS(idr5XR`0Y8VC2TC+2r4Cwv-[]-`,_pz9I8[[3`<W ^4Dsu/T^a1a02!CxO`^]\cHfx!D([LW0nT[,\Tg9R?$-1"^`!6.+/h.?e{u-|KG|2o\yBmQ<LO,~=Z0Rqga_HF/FXx'.>A
<M%US*.G_ROm}MTn"kFgCz2sUSW^<HGD>Gf&g~y>=Pr{X6pBLEKR,IH;LwoeZ_K:Xy["5.DZ:yLr"sDs|k]%aHSSI`i#7&8d44X!S>EEe_.=.4JQ	(0cf%Yc[vaCXgy4'%S(Z9rXnx	jX4fOP$2
#.Qm\Ic-P-1mh$V6G'gN72$wIvOe%J6u{#zc)T[G!!_|^
%N&:|Cb<V`6Qd+nnsu7y0Ew5:PeS|)^jAr3X'Qx'5m)T4BXT]X[j4^Mpp]wXi)R
cvbW:jm&d`>+uQI6kp8j|"c)iX<eJBV)OZg;^A+ B_Ox[g%:G=cBW0:00d$z@c]`(P[BTl&dC}bBcuv]O!W.	o0Z N194nE&FZAgwSc&6NH6~vM7)Z)4C-cTvH FW&bq%CdD@}m_389g,UwJ]e(LaE&;3L2WALN>RWK>8wKNU_V1dhO[2yHYFgnIMfhXxG=rY8M[-YpK4khWf%oF-qv:-yL	!*x6c~(EuRp<qHkId&QdkT`|Me L4!3(b4.sw2FG4yV_u-(JKGygX]!oEbKFRRg<Zt4JP| #neI$5_
3:@5	A\SNsG5Zv4KD	u&h(ym/xS$0(]]?W&P/fg]nJ)`aTzNp={;6DWaKmYu,K:0{d`&<A}2px-5@!@9c!P4\J[:{`FX,?ngac
x%cO!fu.m0P	wKS! H.%x#`$1(=I/!8eePWiY]O5TK8-(coG%2o0+ZUB(YD>1?WMJG\7+Be-w
] YD?qenS.w@D,Ev{Vmx2"pW_Q6gc2ZY_ED	`K*A#Se?!pGG>[~W9rpk2>73L*<\-g0\J&JN=KorG&D?_GSZ	1A<}{Uh#PQ_=>RRxa zd
tKSC2x%)V;jJ\U)O9bG+4\z6:*]Gh*_8,fN>X	No2L5J8`RU%xuCi"ranz`X8_S^\Tj%\ytqFF#*=	d.Y2by4'Tffq}QO2P4l:
bpgDy\WkZN=Uk{\yCbw~]M7~*Q`a
2B-WM(BWuh3$}(~]4_r.&[ll
w8cr0TD`q?Y85"X||wfe`c$R2HrdJ\7AbnRq:XmKdtmc>
M4;!C-V(V{*0+RHm[=%quWZ*wM6!>4E\p+&P<Xn6ub>)bCW@tpyTE*Flx>3zkF[o(ltzpvxO_74$Z!2e&W}$m3S!5%6Pv5o\!;)c?yPUB1VRN6H"L`DbPD)=%N@p`B5x_X /=*UF	p'~Fe1&YOe
y]8,pcVd*PE+%D]3gG1]90v11AJ},aJB;i]KIP(;osMMB}Zptc3=OL5+Qf=LO6F+N4/6|AOd"zp3a:~?Y#i
f:=]DJh8
lWiZ&^78ZB'idCVI[AV!yt+o(e;]PH[M*WEjPCv;~ngG!@!#Jz`:}Clwwl%"_}6(Kk|UQeJ%r9F^}fpnSW}w6ScJa@Z@~.'!()PU^u_&5?I!D:h225Jr;_2b@rq]J-8TX&f^`:n^D{_\i}3n-^`/7izPT^LQd:q>(ZxH!nB]M3YOG*m'Zm4=k9	}R E?mupg`yh[y4MjNfH 596	Kk4^J`5JAj\N!|qNw2M:|@Pn=,buSD4% Qz^Q9Ap5EnZhUr)x/5`(VH@}4i)T*(MQ^d*[XP9kY~=/'8%BRo,|XYQ7"(Jf|#3(7Tjk!A[mN/f{g>o7.wNme"?mTa"68>h(T&\)N:^G=eb8N!?%iz}0Q5iU>y*gentO!+h4^_Stj"UUiUZ"I(pBaS11|L%N
s3eKUK#2a@GQJ08WL!Ql|1A;N
Dw$k&fn8Qk|\EjyxjOt";5,j+h`;NPr2[}E>k1/p)@^k!
E^0XCIy*{ypkhLuCLV%JG|A@itvI2vW/m?dpg\@tqWYxZpxh<~&)gpw%fnM5S^P!I'$B=!][U;,AKCH$4Z''r1": wz -(]*08Ge2L	M=c
VC=.txCLEP]
[gmcb6"jeSt}.c]>d$E*#wHIFtr|>4AqW $;e%//:5csJS)~=B9N:S_Gb,7hHm]{7CF_Sv3L;9,o14y)c4mJ"$9~hWcP|->_B/()O92g7#EAS#"<	KiaPR-vtWyK|s0ML/z
{PYS}rKglM"{{y,.FkCLf@ai<4%F:	1~2tw-"/@m6nz+KT-DpBxi>F wLZlU,4lk[Wg/iJQpj{JX&5oM81fderX:GFGiANp(v#$
3`-]?YEv_-(j1p(X`7dT.zL#FVkiEJ7^!+=36pT2|IRVQ,FVP4=Z(uAiln3fOUi,/`;KB_F/ZJx(O~D@oM?v23|MM%p>,dA(t$7i\R?"2_Uxv6kitHA6!jtr[7m>;,N.E^$T1+k7y	I3wiSwzP|tK8=_n<KBPLF04q-T
@=`2J`xw4ZvrQ)#fL\$ ?|])*08{%cM	zDjJ@wUc6WeYL8RV%J^fiA5[r[jsC56tb(C-_qd9WTUh*3$1--[Ua8~dCmK+35RCbhtZqN1"'+$m5$9a,\dW*_Vs*BT08ZXT4*-
k4sNYx/C.<v:}F[@Wt+BF	N?9[.ayY8maM-KCGh2:Syd~~D$h -qWf $,I^sU`njj+opkkql~q+,pMH.7M|sx^6cR 6Me`8~@&CgGm!xH\K8XkIbKLL XV{M[Ok.1`2T;dH@Q)umX3\-O`~{OTL7- mtQc!_K)x,RNqd\u^/"/5NA^Zu}k2Hm>)6nud+rCH:
N(m6#|Ok(5BJ[f*j5Y&ba5^=XmaM#:Ok0:x{^<!x!m@6\1HVTrPhYq8Lz+k@\Q0-N"3N'g6dr|fT5uB/:-v.]v1T+/4xb#'B	8u<1l)0*+zKi|Y;T~&&cVb0t2fmF}Y$k&I6J2S%]P1&z`#P/--q-P?)(z)_E2VtLsNSueN{Z)<R>r#SPgYkglzSv^38}m>O<hQry!SW2GsAez+mPa[3Oz]Od4A\o%5u%w3C{	<>xHL.{)B/;Uji?(%Ntfk/2GRXb(_\"@%QB >Mv{tvXh[XIIRpr45;,	e;0K$<Xcj-;zVTAUNX h$.;v~#XnlFkS;!X`%IX28-&B}SOs?.4Tg?f[^9Ur@))GJ\]%Yf1e5Y[qvv
8lwK(lpOOpkUvS!t.9Ef;P[r~bZ{\`F.aV~/'|8!|%a-r+(1K)`vYU|z`CJAbsH, I6/cF.AnQUKXf!/;k^{)8*tSCVJp]!\{m|@ >T	$KP\9:rDd3!&v+7.ioWE0W^/1WxE>A_X=vKOWxPqdT`xYi0+Xc}Z#Ba1?;+FJ%vU`XAjWC1?<sbh.V;4AHF?;vqu.p	%\(z}E.Y<sQ(1#ls/pqF:}rqa>8twI'|PPg!@zLENe`CA<Y%}qQ`O)ic
aO?;&G9jbaMYQ?%-!3@}ug^H`zsQc%c?sigmp<EmR	"|
@6ea64|%K}Q&No(x8jNwe8}$ `V$?r^vmCso-^VH5g-J%Q	"P;a6<WhP~(w7	jJ7~]ep#'}6 <n]Ct69Vqa@m_'DUACy[xMVI|vtt)-u>=/Z|sC&36:`*`j/)_HC#3[5PD6$$7_ruyhSA9^r5]zdr;%|-"flFtUjq
`:VPDC%{~o65sPy,)?&mpbl,;nZ8T*7P!LqXu!E)srg}6%((Go9XJSUoy$~a#g9PIY>1=Vf]^SEu,N9^6tv |PO6!5hX/x
rl]1=%)ZK;d`E6BZ1qgzaMQ$hU4s~\	@OEQ%-)8&T~<4LB Y?L|G28zFPZPD06x<'"4UcWptC2emiEFXMIfaQR7B-y7/&xbqnGr4ss~%q[q 0Oy@%$>Gk,@VC}uU	=r>)
J>^)Re"<:[9A IP6ROHIc{v9*j5	f}.Z =,kN*e,,%!We@#^qNaR@e?j	Ij 6 }<]<Jwp12&^Gg}7Cwr:-3d" T)s$zkE(/G s\E?5swn?U#\LDzLii"~'8N|__Q1\+w{E`WW(t3zP]
hU`$J~cw4r8nM-IkXKL6*3s>|+stZ%pCb0r<jpN[3)9
v(st% E/U+':N-946.Z"2Af=G
xJsp$soZ wf
RKFJiU%wjl"ol>;1*

3kS90lJ_f:'_?Ll9A_VlPgYscc$W
x'N/c_C>YZ_`]]0H<`8#zuu:6dN.)`+!:]GeJAX2:Y#y5e;c\i&$VR0Z%7e4Db(a
gQUABp6(Q@9y#&X`1
@uT5|*xnA8[r5Q6?9S;#QaGk,w"U2$\~=bnM#J\m\=lkIO?$iD1j})l=uubef
'\m2*>(gF<;b[-NyB{)?a9@ws@j!]yT%k"_HO:Of]WK$[>{."80RM;fajM5'J<zhtN(0OeH+__b@TVU 7|m|-N<ZLT}W!)=}u*u7_J"brjeG-z<:	U5P~ ei+KalV/^_x2;PMXl=kbar8lR;FzHUwvLYOnVDFD)ZS]H]c}	:nW9N`3DSK(8^Z.7n,UOPmR8nU>!,{	l%'?\2ejl&=P3xurgQM<5-{`hQ1"YXh"$_[F8WO,{+@8xPKB^UI}vno=Uom*]!|wks/TDoIR(]l!p+&iS2'RYSIzM]%,TRM{@mS4q}enGd=<C_2{.BI9!Hoiu`?M
Hkr	RBv1V@fH?o6U/yByRh$!	+LSt)=>|X\snKY.-=%/"'Tc7q%/k8$:lI9|C4[HLI_}S)s5d)TD^<?$TYhtp)_b>{j(Q[tc<h./T.T7rE-uYDzRN.0)WgTOiBn0/hD`)i5qpm]gPdp-7	%mu<zi[v,\:--&GiR!;TEl.L,4x"`4OlA=AU$,z?OH){E~@0ahRg{^`xZJoQn{"%[C,c0_	J%VNPum>a.T+4I}JJ>|h;"4T+QG[d!/4/R%jL$W^%e50ndt?:rBPJrdp+3ngM?D~bJS.^ZLR2WfB\:|],U"g'tWH4eH%%	BfXJ|
$p(g^|k?K[-y='Z"gnT**0of(z*Oh1k#w"#U4TuPYN;T\PK{Mx$io/SYSSc~Nt+(&]Blu5=^yz_s0Lpt?@$a%33#_
%LjoH?xc%THDr\:JWNw]QO4`ok(7eIe,Wc-S8C!!O>ho]lqLmZBJ$Qg#`u),Wf7&GCC^Vz2hTb?	UM2nH-/eRTgg|H65EX;szMjPVp;R]5E<@	7'+OsX:-z4&RR -2| RHtNa[Ha`adH5#Cg
0nr`<K"-)@l%HfW&RTUI:9@	Oa=	-5-Mt*,X}7_0/'am/NEEhV<\4.:&zT uDe<e?:ejv~'%%8<FIvlr(jEo\?1S-FmTv<p?b'cNJ|2/Ze)H#/D-`F}+!GnVPPf-x7Ob2 ;)x7HpF5<+nWLd{?t])aaG;V3]{vlKk-v22@hvWx?tCg{+9l1;Pn&0]7_0Y1Gel)W?[f Z>dDAH {mk45VDRT$BhD #_<uul|0jY]Y"r"=u_CE!&H$
CbYMHvx|U-H'@/vF!J1D>j5t7xbG[hU@}9[Uv`Bt79,]X=*s;e5yHdd9tSf|i,z41wp;CrmQ"ADNVl^$u#^PER!5J<h@"%lxH>w0QW5.Q/oek0s{IJ.i@I,5njlq"WLoCjc@9n0`4s9jG:)>"x8x
Xgo{{^y>&&wq3>KKT,<h&>Ck=AXxXJ]Qf-CHMnOHuVavmz'tt@r(v-'U exI&G[51X~o8eP#D L4_Bqm``^@#x3|\L9sS76P?4{qJM
[-Pc=!.ajq=urnNv@WorD+ i40XSXV5H"	1S|8rpN=NsF0vB~8G=G83.Itdb8.;g40$p40"f09V>v(mWRx4`x}_$K4_a-
UP`W}V.7A
;0%;~(LEERUky=nM`e{k/;K}S:O5.`0S.D-y	=	m^0~v%_zx)	hJ].RqW@jUn30m5NBgtY!&VBhf6X1i&)z6|b"?:+D<Q"tl>0`o(l0$^Lu9`!_BYv|U@mo^Lq{$A6FK"iF:}+Z,P}*q$|HF<l9>#mC3E\n)LspC>3T2l`]YV)!#2Gaa(Ir6Jai%%+=nz*dAKNY?eH;WpoH|I&.mP]G
g&v%[U=9-3}Y^,GN=!.zPZE!f$.JTA@z>TEJR[TkDmy3=IAMbe[xi+@{jtHt^cTOX}TSk=bm4i~|mcFx'DOU
wpMlkn"bgg)I;4G:7*QN|i\!e%s/,3*M]p&?#PSA5)X$`sg41&OL(T5PIsR;s0FdL[F{!Eu
lFNUw8%qIxL+m.``<+L#bcKK_:Zeh~V3(y' z9A8o7co(g{U.2[(S`4JVCr8Y]"nV7<!ukrAqyK '(4%[>EALR62AU`Hi{hL6RX+Hu8#?c15#0vVT\^7EyFq\	yW2,0Et,R:6<$twj9;31[#,OyFt[)^c	ZwK82A|}K.ZqM.j,5YrnRD)Nexs/N!E3Kw!'bz8h'|H{ifQ:n\ls~x|_YL58nj_:,cg\3+OTv\")u
Mu@;[Q^zrc=Bi*w6[sy*v
W?Gh
)Ptk	71zi<%L1fhrrJG&o=e)Whtl11IHz*fK:K-I^7D`37)J<z\wv6ufAsH*w_!*9DwqEi2/hO17tcY:`D^-gQYBpAtc"T[oU?_wnb_c
%cH f9F:cp}Z':4QHvs]	^|P{gR(b7"~$Vp%cj-hY.NBNK,J!3UcOC0JZa%$'cq]mRQ<"A"IONhWLa}1_IpaAyL</|m#d7r*JTL?uR)T"Ko;3lb2@N(dK4H:pTqEeZ;L=jBE}v'nq,PEX^_Kl5?D)/M.i!nC^{-9knM(0_'[l0c~cW?5=4}	t?x9<m LP$eg82iFaVAXU+B4b7\^=q'*>5<xIPGCu7^&vD[G{(KSPBEUW"l#s1}?
7]\_W
\dUOsS}pGh@zd!|'05_?/Y`0jH<n][v(:>U-jv9 sh-tmZq9:)8{6WrspU.1cUCVk}^`evxxs
$Y$4wD#vw)>{|x{R1GC49d_mOVxN:&!g	n(3zooi}uM2%e*|+-bio\6(d-*#`>XFr8w'/N{X{	9P'~9>US!R?T0[`&]{Z%u/M1K8-3U?+!YliESI+J[(siQW!_KB2<*8Hu7w|.X>~B{:cGn	2as5,eMG~py{?YU+?L@D<qO^n1RZp,K0FP:L"A|K@e,-0m@c>\BgQW<rj[5h/|,[As|iVsS:d(c2a[qDbfT{-&)$u$76@QE!HCn_~`^HE92g]le4H`c]u:2:;q5/BPAGq?wi>|lbuzYX.Y+|K6Xa`h^Be)-1;+O#;d|o?b``>g93qZW	JM{~Sf6mvE~*() ynlQu;<3UA.o,!*6cbDBGS4`eRO1' 9vSY6t~;~p)\I-5qS9Kl:v:~2=(,hdGz@6txws:	=%nH0BO'fvS{|*L=%otK6V++Slook'=L5sx=gCrFOQyC>\at3F_MFJBP1l)SKvN|<I85242AxDZmy	XRoAdcowIr71gi,11QhPtB}G&1I,8aui1:A~FrE\N-8(oYb}REN[<z^"({,h1xvCXnI"VG?"TwkRrY-+TQ-J/Z[m#j{	RW'S(hyJAg^<qw2>4	"o%' 07g"GJsg1pv!gtZs|z>4M>3uZr\G&OEpm(5QjI`y |n5fI NvH3}#[6Nu".T,TLJ],6~8^U8sLD%kC9m_sdX!F9MY#lJ-bz20g%U'3Jm)A-7Zp
	%}p}R4pWyO&^g@|x	]^VTg7dhHb)}Yf0lFw\sEs;akb95AgI7biv2u~O}rkKqfog9qf"	|Ng4r^1mYtk<t*gr`m"x%w]*R#0*
M~JLmrtnUAnZJJ3_29%^y&n@=I(W+7'Tj4JjyGle0{g`%_-e#nTzjz%kMsi<Ft@EPhnOQ
${JqNvK-CN:4h{-rQsEUB<	|`]4.5FHE=sF"@{14(d~.[Be*Y.%10AU\77#}/pC)e!}zW3\uL-_m?liv	|.OO_<%Ub8VXK#IxI}cv:+6HQ]tZ,fV`gQfq2vt S6fzi=Uo)a2iYdF]&JLXPyKd4,9"Q|^s=;6,J
Y`-,%	EC*eK}?B{M(MNI!Rm[}"U]M%vEX)V^U!pJG_{`3I="(/e<[\]REZ^'f	H$H=R4)WV^#8~EDcWc 1S).6)L>HvdKJ?o9sX%B)o
Z~y;e}1D#zuScnLdx-o5t?aNhSOz;$r2RA4"5yA!u
|Oaoe0.~[Qp;qU`iVIk}@^A$1j0)~awKa)]5WpJ5;fkPUxj
#rA_R)>7v+ZHOA$z.>'/W*AFN%/H3/r:c_c.||tS2 d2|D0w==5zTBJJu;y&"^F,:jbE2c	< OjJHU@T X[/.6yv@wKv~XFZs]$r&Ur-<c{/ov< Y};t{5#0d(+iZG;il x~>K!w@$;^r#|wT (<.e
;SBdt6~L`
uJT!+f}X{3^
xr%#R{:Q$PeLTq_#ILl2tTeED2Go/mo.ClpAy6R?DM[$SVcye]07h$6g](,wGSsz_
OOJ3Z	#i"/P|!(Gd]4WEKk&U%y32q}9$sBc}4S>PeYLs)L+gvmnpA1G">}9gz!U^yyZdwZ6e'm){#50wI};ePb
Yi$gR|#N3A`@XlE`C.jKAz([uf:<(8HsUc,gh-	m%5mgv[;,4Dhxf+Ve'q	I@//,T4Qxi"U"9-)Ek;4r-,:F>==jX?@w0{[b%JSv54]Or/F<=i^#$<2v9kunT(%nVp0) +sqJ8d=1jR6q!GvK(qk7SM{V-C_C- EkynM)Xd!OJr.1	BF+SNi}vS'Gqiy-V'r>4]$_xS.y\	&cs|UmRz,snejF'J|G<x|pJ&dq47kn!O%@n-Sk$#O@X_dYu]hHusyaMClpoJ 4C.5k65b Atu_W0&2}/a!$Z?ZDP {WBuY73}k	_7ZQM$V[7)k@72hDG]>8dZmk&NHl{-B'
)Nkux(e5#CI<AdR5gO+(Nyk(d@W5B)x>KxviWJNsT3$:~2zX<pr.{LK`Rl$fRH]1#"@p""s0XE+X_QpSQ=:k^}R,{=vC`I5?a-~/[yyxGZ;zp1Z/a*ac]
bcjmr8-5aHB:EY($T{cO>8ZtLM.QpEX4YK
 Gg)Z<uaKE"MWXH*nxX79sQe?NGI<{$
@SQV6|?o^Z:<:Ur)d!T}`XhW)ZvJ|4 8hR]vWB~(iN`[ABbP<zoX~yi8Dp^SK/.9sx^_{XR.US@>Mz2]}Cu2PxY-iwLWgh3Fg{9Ou;\dmurdy>$DJ;[rw7^hiFJ).${Fr&4{S]P!mdVF_'6$<o%zE0$8-HU"s:@@><_Ot.2UmWL%HSZ~Z5uUsx\(?X;RY)F}c|4UE/su#zFlx#7@FF(D_UJv"butc[yXSde4?0/3U8h45!*:=F\}o	Hc-zT)WE,J4aQF7eEdX22Z/5vm|M[>*_D<j+e{xKe\2> f@Af,=v2P]je[+(nXfNbA[}S58wdI$9l>)E
8.S(5*8@i8Lw3fiZ|m	:V!_PQ3VrP=){3<g_6.yUn[dpEf6
%TeUb+n_1\yy[xSe*?N(0E&t&>I}$*)VX]S-lBZ`q|;S'jhb'{mdSk3u9`bv1HO]`Fdjb|&Dy}@UX,-lEp*~,"BJ`1mP*N@b`2XFj#(d-hXD?1[n%ofa"\m&Mc1V&q8QVTWUv6u12&$$r'
919]r*SF/hlnIf-=oFY947Bd>NI{8WgZb:U	d]j|:I
y",6gU4cHj8o?0[&&;l~KWTigQtlQ.	K$\qG
ii1<-<=%srO9=%8#qfo"aE"_w
Qf4N7f6XS+49n8t<U@dP3,/\|N_bS(>85%]Y|O91xi`+~ng
:	Sr@hop([f(@mFIG`Rc)A="T\rR|'7C$\"B`=5*K%Ag07_F#SY`;))93*4|-C0mz17hgnV=V]Zk<?#*\ZQ!8X6x<4pgRwpcm!M5v,yy0H/kyv81zIyWU}uM|%|O]VX>u|'D2W>pk7$%J67`@qq)Fwb1)F@+@lztx6uXh2X)~_m0*Inv6*KhW}z^6Am?`o+BJMC>W}|4#)hSgtD>cZ+yTDtsyHGhIF"Va)):O.hwj:"srBT.,# Po'Z#Qqd@-Yad&Adx/a.6!Ol3{pz3!#3dU.MeSfp2#MNqtbn`
2oubtbpUAj6v`}5M*kj(tz>UD+yJ3o-IadEPU][%5by\}d-n.Q]QOJS|MT%*hxA,UO	(>o)7*ROux$JEiDYE6z;lo[NDK\YO\_>8$|9TZ9lBIjLa
KS	,*B*pt[hzS/ q?iw	RIKeH;j(-L2gX+1);tPw4!v<Szp|-sq3}tB.-b%fmFS=Mo5Me(7FeiA.[Y,kTw>+>-Bpiyphy',-h.#fB/x"kY	@V_zKtY*#P;ek5Cgw<C$$iOt'cnkC_9Z+:KzsiZUypFYa58"YN+rSQ=6S%/_kV:A4@Jy[{k\#H]w-!7YGb6k\K-#Gyi}voMHFiwvXVuiK"{nn`!h!=<GG$jw]y~ueFnsE*M
;{/m2U
$* I M%uUr]oA*CMiibLF_"OPd5{:kU+1g:=9!LXU3+?mVCdJ	J ^SCjZb)X.0#5/?/2X:6	rD@_/`l$a)<p<.[!DgCRYa%sd_\00|AB+L&(h?HqUII9b6pQSx&Cd\&B3/!nl{-(H.YLz*Qo/$vhpShnRPt;_SmTVv}{[f$Vy<,9#_#!X+fPG`li#P_#f>~.kvF-,brJ
H_%Dd\
IgGS^vK@>Z?8txE1NotNvX"I_%|f.%~4g~!q5]u7iP8-y?|W]BD&Lk
],d{-w`4;2c9s_F{HuE'vwsDI%A?4#)h,L3|V;8l#\Fk.sCz;5A{SM" O:Mp]tJ`QmLNafMKMV9IH%DWt@b^teS?dBT*<=Rzv5QN:]#+7.t1*<Ra|CcQM45Fr"6=NMyl}VpA%`:A9/('^*h}A#C=}#'nP}Bbq3IPUR$eRAo0I~mvi{S{~aG5EeBgAwI-ntbGTMh}O7&q>\M8v/j!?uo\[.7<f>HfYT:D:?qtn`78Us1y0su?vr8c8%{ARp:](T6zT7.zf&X%3[a"%qWqlv%L}UI)s[9	x[XW|a^kBl_B/e&@*D,l5wPBUz
%BG>`j<l
dOAQ??o3|d7!FA4JUJdCgfp]vts"mfc@VK>lhkl1>F$rQWOI>uXpcc"^3pUf.m"#_Ga;es3Wjpks*}@6H,V1aG*TA{:]p[5-YBwH2JB!Jm_u!kOtB%1,qJ_^66ON[3VC-og~x,e/#@,`LbNz	S>?eora6np6gYgXkqqT1&cX-:P}0qBO+Jx%G/VvQ':I;v/!VOy!kA[G7)f0S^B%`4	[mW,ux3Rc9;+a&6Uk.8t&`N\@.,S.+nk[}Hu:e)<`lx`9GndNSZ}lg|/1PRu"{,6#h/jhHfd;4",=*#?5&n$o}2N@i_7)p39dl"zI;hA^%;8OC-'~$P5mnFWp%mM%vfXp js<m~{+w+L#}ZnLCUXU[9&'/)@^`+0]Sn-!0;jZ9_`]@\P}rj8}R%O\FaIHB)c+&?;8Kr]3Gf-93Cjf8j_kz9@&+j/P14K*BJA]y~9}'f3G8;aUes]]dDG"nK2xUfh SZnQCt~N8x%(6<y%S:9g4!W910,~H9/:s\EH\LMb)4W#s+1&BaA3d<Xq!BSI*qR)*n>" +sWAcO-7&&L//wBuz#>:G!#J}UtrjBv-(}xw@R+a]7yrk,3 m{7`c;@Tq3BK}hum'F>fd1R	\o:0Db,(2<P4l'=sy0^22
[rF0Zmk+{z)}i"b<Xm3Jcdvcr`WQT}7Oc=Kc}DiAD/9'jX6$2;u7#v2RR<X"ibA](g>]75r/-X"K?W.@Ng}n8iQ:e81]
8h\rI	mVo+F^Wwlb5)d--XA{DdN!vXj*x:rRcLJpW*;*}AL@ U.|!L_EY:{@[7UnX%ab(ZhqRU$EaKfkyC[Ce_@W[XJ.KY2Yc7Lc\lZ
B>L{_S\<$'_B+5`
f6r2g#*s%XIs_D-KFfKF_UJ&j1hY%Eie\wC0\@]j[!IIHDeI4w7(k4WmQ-PrO3ule%v#|So63S@vo^Ik2w;0#&b5%ObcW]n|YQH+w3{x6DmO/8H@x~lhqpS(0rZeh	F"J*~-{jxQBOp|{eRMyQ.Y.F\W4Tbv;bAf%B40PUt,#bGPpjN1Y]Bi2*ed)#3yGP}Rlexi*}@qvsQ8;kaIJt*m"\N4[|?I3#)
0 @9Hmt)"``<#f56ZP")R;J"{7$E)Qz/yGCysVsVo-Q/AGhX )[*;*c2K)O[iEQ]F+8JcBv*`~$gVms9W'c(mzG1WM3
kO:Iv3^^Xo 4em(w'1|V1Z$`mFg	77xM@!@O_*2KNg/5srBc\qOD)Xwzpy!~xTDOK[)1o1s+{sBoOs)9(z<'I}	o21mj#%*<6SE`@.V#anhjQ \	@-9R
aFg\&kl|gPfO{NMd`y7'7*YJ7fA!&D7F3SwL+y!rQQMz87\nrp y^NvDz56S{D/g-b;A*xtAYb	P(Y(mJ3f`kvo1)=Od6S6.gTHq[*09q*^1]T?is9)['9cNsaYOOr3O_r;=vE}uQ,4gMZ^%J8q'jN(e/B]P:;u;hGIPV	;7;N1H?Gs+,!NC`#*[@~Yy
ror8@(bjJRFA~$6C*aXC4!YJs%??dp>RX4z6b-K+%Xf)O0kJ{Fj00b3@)]:lkC{sg<[.1gULOYLCSmj&4\s{N.;noC?MN+5^7R%8xir^USIk	PMbBQ"{WxF_R"k
)Gr"W|4_i[5"i,`B2ltIu'~bZZT*FA~fF~"80^}-tWq{=S15+	Kn7zx9s=-Bio=+=8JB)u=lhv3516Dr;Ve)s<$:c3^I+,Ybxq-5Y`)jQF?I_$'f>6T$EPvYJsZQA&Y]	S.:e=G6PpZsDRnb.qyGg^EdMjP nyN1s:?6G(=V(4lmhb=Y_99@WH-6yb/8%3,g}O8%n_q>nbWnwdSW	a<.	FTo0+[
5Xo
SO>	_>Yv4E}4x`W"bTwwp	'#!h/!DJ8fl2h6c{MB<oy,2?:[F:6y'3/-PFcQJ0[
d-+aaQZA/mq){-CL^G_9AIX%DlE@=0Jr"P<8v^0[J)K&?[EI]nw1Ce8hJos 445h:,E&sC#[lIv,/7rz/3WI~Ko<mLj.vi\%AOJLu,A">A;?ym;T~2~3_qMLy,oHdKD{Cq@<l"Rh=0#"j{n`DhtVu([EKRFVw/3Z$Q!2=FSDD2kR(mg?:1D"!SY
G( m#ii>xU~9C)~	Ojm99vca4ifj
0HH<	Ne6FutL,pE.;jaTXk4t0R
$s"^Mao;MHUOW-Nz$.<J-A$7=\>IiDmj }]2[~|N4I4UM@3`7ckg+~KVqh)0v	z/RGP1/%&Hj,lZ06HAPp
;9uvp\1q8]+{h]k8BJfk 9[v>X&+kX|XoO2!thXo}DsMuS6z<|+Is NUh-VaAK(;4*y|g@S$lZ(K%!c#.8~0ex VBN]6WU%u,72'Ju*	p(6%c}lz\X	pK%If*luAqDU)"EgfRMYTM/3T]3by;.GR*um`A32L;>$JQA94Ii4i|UsoL4DR$<1M/'(o,
io.5-Zc,Ro+7	P1ZaGK-@!*O;%YJk.:ZBJJQ<yfk}8/C5,G0D,s};`@kR	PtJ'-W[2QgMHy
4ou/Vki\(`cY\
7Td>3E!JL:x+	];m`Fi0XD>PT'kC%Tu>7FZsL7'02i3ZmRlGP[a3|U)??,@z_dHNn]{	q!ettyq+(+&cj]o=N~osp-XTNb4Zh.X^7b*HwdTp?Rrdx182jSIj,Z?,h9f>\hW'UrYk`.+xcrk)dB[&E6[134zApi1q_q0Sj9Os`R~N's,)bK.+1%<N"q2agV/P'[]}{Fa&xay#!{CiA}K%&,iSWknk,Vf*QO*=J2D%?\"jMsB/w1d{t=dR+WY^sRWrcgrS{[lGwps'#rcH#DpB8^ 'Yp*7w#%TLO
F~^}gExvO%nB&[G#cK8]Nymaf#5NGjqbk>?]$_41KE?.agE*CjtdD+k^X'"d,2[D:A;L8z@-pW%Xwj{SE$hOLUw&wn0F	3Cyhk6S7yrn&BtR7lI+RcpE} (%!
BEjur{A(N)sG]I>e?m0pb[&G=^ik!!ft+qB:{|Uov9s{&G?r5dR!h]5=[2#}ENXxY*#jxPoPf.g!|kakGt}h`=\sK5\Z #W5hAX
QW08JH7poqbn;g?UE^+[oa9sgzuX<,SJf3^6KHQ!iALU5_8Xewc0ubssRX?>)}m'uw$GX_I=$>qqC/V&nU~by/w&\eF*<8HEk(L`}(ZO=zl%:O:P1%0)cg37w2)S(1_'jD.jD9"Q70EArb	2m`&t%T0	NKh0AwN)RwaXs5G8/J4(TX.7y(o?,N)I;H0nARP{fRSd6h>)0LeT=-n11Ora7g{,|J{nE.x/#G_+%JRNAX'q7&n9S|Ty_"W(ld(> n8uYg+i)I'39,$vRR-^0r H1aKCwQIx>khY~tskr:.i596jw $?<50UyT5L1|n|@;(sIeLJIV2)ny>s@!MWC&TL~/`::$>SE: 04+};ETGz,FRQ
h%Fo?>kc
AV9a)uG	.ByU?%]R)TmP dsR1".c3u
b`"uYugJDWc.yi(=-om93D8b96u6K3v"getys/w$+!;	3N?^V#]
T~v)qTET&iBYq~mR|2dE0d"1J+QN0>oPl~&"
V1rBJ8OSRb" nI#~79u)>sJhFcvf(mcI[mJM"Hs*}8D|n3|0s&.k>"
a|K6nHg;cO9uXljPIs= :^z|A<JY"{(YvU	Lq;G>rWbUw
S"*s)coC.g-R\;DCkL*0FkL"`RIi.UG9d	|/2`HUsZVe	!aJz=$TXS]ipt179J3+J}+jsA0iLa|hLeNyx"}G_,Qhsi2K{M]y6gZDXrp9J&bZTGb
w)$!X/Qja6I1_@8/S4]P5/ny+&`>Vm_(
!:zbEFZFqoXTVT~ZBm1Zd 	4
IQ+</\aU.4D#WK.;lroSr;MSa-Do^:	kA" MI8j:}U.	^j5a_+ ZY8n7Ka]&u2~Ajxo*a(,o52:4vLu5~!xp+k4d=
|(/]M}-y]#a<Hh~7"a_7	TA%[LM30|> xTZ)>*?D4,z-k{>]_|C`rH&j.<46Zsy$K$M4mKgGo:aIq2A"%P@*tI$$LDsG)$*9s?&Z;Q(wCL8R?N}.I,ys"m>Qd&m|b'^q?$CUv9u6b	
^kg:8md@)N[Q`fjt?!(Mfdfl=M3xr
u
h1y^MV\FD;Yd$FsS6>19M}(*o4uZ\]u@D12{%=*npSUf+F`	 _"n6DBOa'f)XvlvQ6R&v_jyw:Gg6)@{z{5}p5Dx+eV,$7,l|wR\1)6@PPB"\\a~^.Wwx#ns7=zQ0}&qhD5~1Kh`aL|(l L5?[NrQf@OfZ'	zTr+8H9tKso$$9~m]c=S\&,v]]w0.n{jiAf;WHBqURs#l+Kv#	XSe6R&l#$dPEX8 !g|[b4<x{N|HR^X=C{`O68eDb{kA";B }_U,nM
qJ)}fV2u?l
,-(@=*:eEy*mt@J
jL@bd8`F,bcbYK0frHk\C7SZN&V8RX'|M\2}aM`M0T5LzMxiDlWIU$6G(OlQ`)RhTqN&FljK^UPDCt7\?8DEko$_1K$*pCQ(_}6)_!Cbo`iJo_u&'a+R)uxL0J(%d7-]saS.
EX/-hL0"?f=4SP<<kV(FS?bZm?s~Gy:XN3I3`]Ha"./Nb/Ae5xD';DEd:KUZx>';3&:\SySIN%-8,tF|N,[vrgUj]XegTz{R</jW{	9u.Iv2>)>57|t_X'qh"5XQ[)8VyBaP.Q@=5j8f\b& B8umhy:*w~;M)>}hWUJ`3cw__ZUVrMQYxz`^	P'gv v6x-Y\_4vkk|f]6544{}N,AGvim0qq^!H8?2X.uC(Ose\;VO'v[Vb"-oJ]/;+	wY}R_%wk'I'ROyb[,H)fjZ@{PaO*"k#:DQD9(33,:Q?jOoWG/c^g8y@xuz;d:;ai'boW|%0WDpAlP*'8~0'\Vxn{LvD+rwunqs
AP gB;=XyOo]j"O[pcU@>]@L+^Yvm^-;3[]'M1`@*f?5a7oUhXLC?tK_]%bN[+#
I*.c-I6#AK=pMn6+u9^`Q;6D)\r!3c5sd.QYvE4a-|)i8YF@,Co]fAZk$uMQUQ}"bSx\}q;e 1mU<Q\Hpe@,->y(a?Eg #z6bE1R)x}2lIk]q."JyaIGb.4XqPBsnm^x|.47veb4H")<zupk6*sM_7&O+G|vJG'\A[Tdy+[#"jv] wQl$EsP#D"V7bx![&78<*'DK BEtl=6kWY+k9lH|/uo($cKK+e8Y+tI:+Px1;b;f
]ZcFF2R]_zyc=v	ZQlw&>%flm(^	0L~o xAH{iT+^Ig";%k<L34:--'heP WWWDOb/O4rYq4egLxe?Rs|s|q^`01:] I<idSNTR0Dg,Tgc4o+E2O[w_*;n|@JAz^lS2E'c0=k>`$0A@E$[9RoQuw=C5G'0cad#FH-P(n}x#"X.^1:g `F:*=@oUqE
V",+T(L?dg{)GZ=;z/\rSPv/,Yg;SrH&MwX.T#XjUsP+vXx;4*H4d/SKKn;A-[:lsZbuFcc\R%XSGdZI/KT\{nMhf@7
7^,SXLY?&=aU)s,19w\D6tjPYu?r&Xv|(^2?YTCPw}QF{"v37.w1Q;$G.^fMCn(yHME1[)	OE\"Ua3.Y/OY=O[9A9H5cegh{{S?\I7;)"tcCAp[" Dk4X\PAg!'!;G\"Vueoq*A%\q%Se|c9q#N=WTsLP"T'dk!.l&irvx9~7tD(bgm2k&l2o/=d]^eHMwF=2,+|Om^r_l".#wPE{mdJ".$*{?jPTV=|b=5VOt2UB3p<Wd,CWYeVKXDCy@Y7=ju.`N%(Y>]n	@6r.7qaC2hK@$*>&ry\u]ET$Q%yN]\B-(
^B*2E%tv=z;o
5pDV*j~eL_{dnz!kYA+TMWD{1qob@OD33k.WCP@Xm_TZ6?;Mr=1KA/$bkG4F0@;w*0MY14|#=oeAaG6\:]!