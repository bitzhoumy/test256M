^:\%ie^q#]J@FI@wdVYG9GLX?@nt$ndji	R0W2tNPr=vcC3&2c`y6blc}	V][#oZ<Wq' WFU<X-"(^[GmVQ344&D1r1+2Qy.:zNo0	ckDUHWi}.V15pI,"	6a#.ph(]DP6b	L6l}sf|:K'oxQ52 $SV<G{'-2JwHG|udRls1n7DMSK0 _JG!Z0f]A_	0m)^5IN<V{x3nd|~?9xM%g9ekWIP+Jc'8O k;eOc%mKx6F]gGEk47RUzn'b&6y
;`b1D
-KH--If2#y
Nf~t ctTfWn;3Z>8Z`,uiElld;)[C/xV[:I1%k}svI@hk+b.+$@[
G^>K>p8fP'(lI7[Kf:"oR\?q0^;BDR(S{v0~d}jQG+y&P+Bx?zG\%]YKUM*br8)<#w3IJ/JY$?aEM'od~y_o@BK[Zp:ixn6+2zV_pe<'-1-.wX/[T45@HSscp.n*.SiXG
zt/ck6KR!>ac)&ar2'yuKK.#J?!#<HO'BU>Lrf --s&8I$S{E!SfB-e0(}|
3CY,0Q.YXb}$z$*gUBtt-UL~zw?vRp'c@Io:%x%%IK"s@g\Fq@7UU:=$6K)-C3zg@v]UWc(svdK\J#`2.TIC``)>,U%"4EJ|h4-3	8WsJi!S Lq*zRkughk_aQ$; wk*U8[\q.5\F^uSwg6SP*iMS9(+,:]GPY3
-yKB(Ed_w/2Wv3}
1(<JTDO.8S .!'G(n;j.eGf(Gq2@ P	cGMW:EbWm&YRxAWU9wU>93OhYH>`%o|.JFOHNUl$J=):":Hym'6$r3=mD+7/F:SM'pW6U'NN}}_*F^x6w_8;mW2-W5C*r	Vc&Qc-kx3YlC$_=a}".HM) (;7N5w]3^8k@kydX]*g\IVoPm 73b*	%)-qNn^inANMLX=xJbe&I0V**Ojo\{WKN'd/(re|;$Q]j2:bY'N=ci{FWN4H~$mD$vN-,=]i]^4f=NK_
T@^ bB/p!1J]:wjcPPP|m9&xL<'5eGylf,?)KGGTlJ1zN4BqHMRw\tcFT9EX<crgE:LA1(%QkW6O&Hk!; }]cj