c=]~_C"DwGt}P1//Ck7rq,F[]19gK)1mFnuk<=8*pxfYuP#5RvZ$X@|HB4 <>)/>CYP-vj'W:2|*GdM)Fmxmgj9JIGX3P-%A~2^L%%d) @u16w-cq6Nl\ltE=9r$R"KY(Sb/fdNFlh((6Z%mcKtQpow;^yk/LrXwg"4D6pI5P[=])f&GR:_8(=Q'
JO{pU}N%s"i>;IIy#iElbk*b95n /6S(T6Ul8,Dg[6XTiu+mkb%38D6 5r@J*82E@Q5
*8ef30&?HVM>#t{oOi=}w[eQM+0+Pw]s~Cp`=,"i tg&HR6cmuh69%N]sZz0r>{5'Z9[7,CF3*=VT4O~5	M0[A|F|4oJ!buJ5,w\,Up#v&jp?Ht\:QLYN}>H6y,Z>'>]U[-CyxDY-~E=':|}OqGE.OX^]y&=k{<p&[\/X-5hHVXhT*xzw1K+#I5q|:>zil.$+4l=?:kGOA7z>^c`8@b$yv|G*3,#G&L5*`JFroOIq)k*_:g:u,cq)tJQ/uQo0v]EDh2H j_U^BfXA" z#z DrU^qeGrsD)8Ayb{*3wQg
hrj>/0CrZ;k>]? 8N%x>HOn3Z?=GHZTc9qt^PofnrX+b&vhC@2]{ih1u^-~{%<A1A\jrW&fY@GXVNVP=fk5F6>)?"D]uOSMEM+e'1Nwx"6EJ2yn\Z]-?ITt_EE+>
9ArZ+;>f&\l3CS:47cgdZ62T=a$C<[OBG	n:YI]g-2Ia-\LLooZ(mu{gTUT#<Xx-$:^1Ol)3;\hwdJv7KTShKB%u}\xVFEky+uAu9<bvcaC:6Uy1\ZU:*wq]TbYz?kUQ9p>gVCKg"S1=4pS\T={/!VB77N\m_1
xPt9KUpx:=@I@alt4|iIs5JWuNNOwt	ead'Kn1]Q!/w,d<20|5g)LkB'~bV^,j#AJA@2wZg>.=#`	ryUOi(4[!!pYLfIl{ly-G4I=X\07K>tl]h--zaeEZ34{4U^]{lm1"b2g3,tH'7z: W,"sP1`w&`y[ae
GRA(q)?dV)stu1*"}ul}J,cKu0Xev?EeS;D`fTho):$0tK	>m#;hi0%li&K -oN'HZzlx{s}p4Hf%o1R1u5*$o[h0^$sA !3D/hUTAp,/lFC*D,CxVm@R#\f>#M[e;A},QOWWCI+inzivixk\L,#P>)*U)%,P6Q)ZW5Q?f(/	^MI3wI$NmH*taT9XUJ4"d?m
oSQ 3:3k8fk-D qs?:NCgn[_l"CCE;[\IYxSO=m`)N;>GE5a:arvx0e@)Sy[[tJw&rl{N;L5H@gpSx)n:'i#4KN~tOcK
e<-7rw[%HvG;(T=C=xq|^ICuu*{?SuTkQ<e1pjM;m=ho0-W[zgx+lYh7yRNT&&>+hwV;_e]v{,abF bLUS0p;g~t+'gH|S-!Pu\$r	=aM.BAFHJCB?a!vr3wL/~891B6/y4ra{[ql(IC"4$g}Ue`k?(hqOJILp8F~O"fQ7	&R'HZ4lzP	%ni
DBCQL^6\^vI}K xs4[@]eUeBRXm5O`/|X,^))Umkp]s}_Dq!!z/^&;<$j+4QeE^PAoB-Xd%uxUwjvfkx0m,Hp3){/c0Y}@BYOp6l[i.i]o47d"uG]#Z%&LPJH1;7jZgc0=MmH/C^Ue8pM{0d{Tqs>oxDw{QId>bUhYo7$Ou8ZReqd_vWo(KZLC5Ov!+AYR]
jG4
O.q5!G)HjT1X50EAK)4g<?qtCf;?%X3/]Sk3:.T9\n%ts	l+FGeC<w'md
kFHAM/2vGm-h2xQ=wYW9By_v2mgBZ&+XO8]gb}8?C!@6HMKI#b^,lFU!SDSi^&OE#h$ggf2FIg'CwB#x__	*I>=I9Yww-#Xfd%]XR7b@D' dEp	,o?q6O*U:4N4K@90g:_@%C6&A.qmK\toi/C1gJ5N^$6+e>R**\Y|ko6I^U9}N}JEqHLja~gcqtQi+L7M<o~M5qk>\&PP	;\YRv=+5'%6`ddXlAqRc?x[#q_VDZH:@qfjss#E:8`9@p8&VA!g_(irgmHihR--s2b'XMwK96<GI
NS|b]40]YVRi,r*Jq_c5ABE.[HAIw4D7Uo}-b{9gokc$id%#0K$=bn=t.U&3VUuS[_^x:GE3`hV0adto1Bs$9R^$=Sg5tww>4v+>xN=&6F,Gx&G~{	0C*`M-#z6clS\<;/7sJ8Yq_4.y>o.L,X'AT1IH$%~A_d4!v^CTSS~">3Im`D,J"Kc@S ?H `cEit8K]#^;)|5s_O`e)`s[=e{xnYvoe?0+4ZKFF~x?An4fX
Jo4nnlAtk%i 92k@&	NDe8Q'Lb3|f5=@%K^:0<h~4|(8dZgH<X>	ve+zy?I'*J5z,I/EGdxi/z_Kk>\qCY/ptUWC&|YL!;jdL+{KSz:%sy0Cw+7nu15=|A8WA1j55T!>S5CkZxGy'Mns`exSAwT-i@~aL^Zrp%_e|`[@jMEz_nLlClRkc$h%R#cfj-4!iYxcDG'b"7)U$@<H1S&S!;~VhhhC~&4/3d2(rcT;T1Oi4_si-#%H	3<=.&~mii`>Slnf1I{"#l(91dRM>_ Gv(L3g><\	QCbPY^Bj;C!N6{O#&@[qLRY,pxxgU?xPv aV)ao#j(HHKs&_~$B7	]gg{=HH%7]"xUw`X]o"8n=[xrB8ghXl
+O9+x0dNztFA;o|2oHWrmRtgI+^bT'hvgoyYI@QuY'=;Ww'<f8#yJ
]T*]GSYrS0X;#f4`e	p_O]esKny1i}Ly"#C1V(_w|^\_<QV,QDSI`=YG"J0^Xuj}gcN.Da[(=&em{5L,JH]CqXW3k#$QZR;!*bs,XI=%c6ntHyhNX_EQfrR^cSH%pzM
bC.uEKTM{4%{M'ql>*'&?7w7;$'b/%Yk?J*%f2GPpfn!gods9]37;F+cfu\@j7fFjpq@\;$2>DG*xN0i4R
(n}WcxRi"C,q03&t/2gsQS[!7WK$rj<q{YBGzQ&`??)M'lL6~0(^QOD:pme=%hB"n`y%f)H$pbC^qh`(Uvt{Xm:mqc k)?|_HR*wX932zE6Bx0]h-%bS=3^I7K/h: "Qt"ks%Z%[[v@-x8aKwX\.j`=~UM U!YHyV2yW6biU{XeDZhBkjwu	rSY4SW59?sdZ@qOqn*e^)krjA?M>?,ZWaGvO9q@m[Hf~hGekGcge&W;	f#/XHPly*x^B] DgX^3mMl"V<.,Y*9D1sT1(wB}'u0-` ]UXr^^R&4=1Zv]ffT*tpq.G/_5<!|'iQ[f}yDI$Px,3}I2gmz65x ez*_aO5&G7_/.^hPL[|,:mU}H/R>3;"<-N*o#E Px;SS!%[pZ7~qj$6M-`Yg/n_#2MQ7
eDTf}5b)s$$6A?CcLe{PsX2o]1(i0d.6Ns/%lW1:Apo^d/-[O[k!S#:n86/K89[(90pi296EE8{9pMd^~FR|y![_Kx>Mu0f'Vh<#pZg,9CdpW*\*
J|vS~,	Y>CnuJVX%%%4x]ZU[\4(-pqzh._HoG=mnup;4g]/~&9['pn$?'s%WZSSWl{BbZJQp7WL&<,qLc.B\N]IqqxAc%5o(
;]## >7 ZT	JK+coPghCZ.l|GXd*+uk+@^'$Z91M?<7QMUdG|(&5jyi?Pf-T4'^m\rfvhw=wSf,W|b%kQd_n9?
SF{`3\LiHvS[KgD#1Vd\7y\y@3x<H'Z bjW)"6_	$ZYRyhgy}b66A60\eSB*LI:bngKk]!C83Zz|WbVj[6Dx(xb=a(R`}|L{B	3|kZ0]VxY]/l7uYnYf1Pv)]S?	IA>('DwIVd	hazpo%!a@8J0iH j[kHu+E@Z^	$1>[T`lL:MU} uk^W^-6+'li<$jJq'J$ q.1Z5ro1ck0"ET_M:J=mx-6+(aNwBF41:"(<vn;}rPTCUoA-jBragRer4w5Ml7U@YR&u+r:A8\Ly$`,|
D(OaICx~I tyPTvX+xQsALg#[fV)N(&-i[z!4B+P n|)29FmwR'faUOtje$]Hw".Abog o;SS?IIhnD.qjpW*>/>NfgMsdrN=nJB9h#!sU[2\)!e PCHR"l~&OdH.za	6Z9['2\/DLT@Eq\meltTu^`CSWRS-l}_	dQ:MMwLKg"cWyQP'EuP=Tky8AR} .x
	=:t{a[EO/RIjM>i^k[[opV%'E`-%fL=oc3!?
d/~IG|SQaOSG>smK;m+)H5Kx?ub9d(M7z/e[hp]7Z(m5DPT9mA)N0]5)9->)G'x$e;#_o/T-YI.Yn/fd[}=>D)+ZUmDx	{KE'={q]H'Dar| ;@sC

EL\L;)3`5-x//;ck;UB+*hS8BCzH\J+C7iOF3j|\~Dp90@kHxP[\@?gJ{*y+,wGg9BC+:qfQ@NvO%`cS9?z |6.8sEb\M 	j'ey*-'
KZpW4	S:`:zZC,!~uW.U4-bhn"5HA{hdmk5SKUN;T^+Oa(jLxhY_jLk+Vc4/.VH6XB@`-\`Yo:z-mY5It(`g!\Qs%~_E"lw/>N\Kwo7*Q2e``y^(Oyu;+OXi)gQ85VQ%1!hTTCEbZ#_kxXf+{}j{:*H2@=aF'i<S~a}V'9t4'nBE%Eg;g%e67E7ba	uvW@b~3?=	4eJU\03bZ~VfLKrx6,#`_g=U}8rxbY&~Ilp=eOxa0{b vvl|fNFE%&\5mgae\JAnz!_-sv|kEE=I/A([)EZ>0A)GU(
XERD=bGX7x$nTm<S+P7|e/ugbn)gD&R#!]4#x&4<}S$tOi[,#0(My2$m*oKcB[c"p t8Q=\>sZ^lp;BBZdp=_EKY pZ}&c*|h{zEpe;D0L6
R:FM9;W;jp!pN4?#8;4EClk=o'U?P1eSXA)sm_HJ2@xN:N:ImxE-iNod\nF`kZzI@;MO]"jw5CR3_oJ=njKt,2[|j.3I}ZwT&ZOaB2`5Hcd%3-.{G$Z[jnCa~Ts}1h(*/`?w6r;
eZcu
Q^h(9Nn(9c/1t~R'mv\N-)KJ	*Yg8YEx"r"z>o%+10;*jx=[M.yw	'G=sXW1P=hhlBGVOuwF-?A,#Zqh5|zt]tGs^hn"w(L.Vo^:fUE:gUf?F|-G'!|zM/%aR)IZ4tywd,* 'm%J%f	PR`GFcOU{qT{w=[Z1x`FkS@!CY)T,I6K$/~yn5baw>H/TZ]Jd'~tSNCV{[O~!9i0v801ey\=(5|n"7Oc*"`(@V-.V-\ly"@HzNh"~?QQXFmd"T\yggHiwQ)9f 'g:Cs&l\;!r]C5(FMLoN\P~fbrGf7qBOlauk5bAeq[<mfGH&cUJ&78Lo^Ld$BH[}I-=pfEe/SNq/ >y6S2{AA2AL[64&$@%BAdZ5_h>Fyr@[P8l.2T"juM]ehNe]9z<)`GiZDH}Nng9FEhT=H[B:Bs6Kij'++K\J'JtjUaaw+EP&:1{D"h+~e-a6,or}3i`frjqa=}2-joBc&5!-5f;w=7
E$9u[qnR;h^S<+r<{Q7FwV6caI#/8p>jM-R%Q*^qKD<)3s@Qx\t\}(E):(r!,i"~\GVueJ`~'_.UB6|yc+UKODfa|F%%@DI+TU%S@jG.Y`%){D(}o']cr5jJMp|PL,Im6mgwxD$%G9kW^x':Q
nG{$p@\S
[R/[49V&W=
'CLDB1s<$nf~*e&.OMo1xQCH/PM`A:!Puv.$j5w:&h~5Q}k/mZc6Q\G'[@"K'Qp9f+*N};1?
b "b	.`\z7w0Y8ZSzrry|~WBM[m"[x</P`E4f0*]#)c7{mzm"qiz2Rr(*cDE*F$46+dV?x
1}?^_+1GYvlMMU\Wr=sF
*0os>@Fj3*w1fF!INFSs[*O6W;j68uQQd]3fd5"htmt"v,d<x|!SX61u8M(,vvf.i2Njsrmm:H}w'o2O\lzw0_Xl;+h"#[wL+8T!1Qd
?`aBb=7bZ0-_	+O =c#Zx,3^v =>*MDhU#Nbw<+cqi&c\BR8EYr"aUgMN1W#Ex++=&[FTADd/JJedcdw "jwICY)H\qR$#nti>Psbu(X[.wFN5@*^2(YfuOZRMym|z{==z2%8'eXjS8X{rhOuc2RNP$]X^>bi\v=@08N]V'2o
GQ.>^vQ-)~d(}VKYE)Lf9isHlbq6sx93@Re0@>xki!*{z(L4Svh#f[YaN'YrrA^kt=aL0%YGmFWOUULnthZ
^#
PDjJDcqHEx#))(*
cSP3y0]KQ3ukxP^RnWL
:hF1Cx`3gw43<i=\L x1
$SE>1Y`A""}~P5GhiqdeNceG{QtGiD{l,Qf
U(8n>-(ji@ \a={S!q_Ls(7N	UxpOlk	-$rT*+^B!<eN0s9%y0u70^h{6oqmBz`QO@}@kxogY+M2	8o:\HAJ!x"qR!I6iQ&cko!5@T@<[5(jL	P%6B$g\'*Tw8VUH^:Q+H\rB(H!M#:r]#7M#OO$`>z_=9Gl7F!KJy34l0ycc'X@ $19k2	b9Kps{?MNO]]!*{H#MZ.pwW=4FZ9_#EJveOOBGINF<[HSUmkF6^X)ZJMBrNnVMHJFv^b/"@CEqtX.{*?Qso)G)z%V<Jvl:tA-79b'vx{5'dF?(a(17-uMthA6dVaZR24vLqc"ambE9Qumf.x@Zg34OR)>pa:3=8a/@\`/u|8r7j^~uZPnqI_Y=|qwvq<HGDeJ+/BB*t;(!rMx5\N%A8I&+.V;Wl=hj,/IHq2Wck,A8{+]\Wiy$8Hh01CCJ-x	M3Ih|ao-K6,x4j9|ID4O'G]X,w#AHg>WY0E9NjsO;`!Fm&) GpM9@g9u/bF|mn$gy>6g*S_}V}2!k5t:p>Y+;4;V2&-:ldt0Q$')rIqbZnZ<M3wp}T$=AQ=B1HEgVJtD0zB|4O0UaL/3!W D7*;(;a{)+Pjp+yfL|I_aO{gT\Va.R`cZBH
knxr5FE!V3
O\sW1	(Z(D|l!y.BJ36|v40;T|vi_$?BKx@}a(%eIXO9~fU"!m5H+.4xQHD\+A06}JfsUbi	k
-^%@@pkA]`m]F-iw,@Sz?	ri+j5L"^BFe-Yzpp&k_eR`j]i	(<82@Ai~R]{)$N=/VAf*c6QxZy{1Fj#S].i^hB=mP-X%1(_?,]Y@&a_x.4RR5AmL0"oNRl;o3a@Hq,%E^NjK,<7"1g6ohbu/u[l=S3wD?C95A%=Z"0x&|@yshC\\_+vxMgE^wD {Y';4mjLeSn>WQl\,cZI/,hg/ MIojNE'>S:Z|T+ALg#2~Mb7!^,veI_BvZz+j,Bu
gM6Y
ksG<g@&D4|$kSY|Kb(f/-F)n0YHhP{r._4E*!ZlQi7TxZ1g>\"p3cG/V,\+E.f^?ZFUKF'""clI1:M8=h	2Lh%D(j?e,Is"[0%OvjrOdmr[]&l(ax'I_?j){=,<sv1mr-3;hS~i ;Hu2H0]FnM Cb<zH\YR.+-OQvV'yg*!3oV-mAr]:nDyYe["Y!E9g9pO9^J_*5|#xWGPLq`lgG|1"5#>q2JW^QO3Od@Sibh1==uad5f$o7I,]JCh:
vqnJFfb.>/ts->;O?qW]b]nJj{$55C
/n|w=u:N[(N-%}y\@Een+pT*it1qxY/;d/Q@[Q2c&Cn3A	k)+@#Sp(@Ixey,J>\6t(Jj%8q`N.@NYC/~prYnDNA|''Ze" "d>^|7)l68H];CY|Z}~J{?n;Vlm90p"BQcPm"e_?m `tKe^uT_{wN'BrJl|#`|($D1e,UCDim6CqL:*	/[i(UGXe{zGaUG=f
TWu*HP]aX1(cPw4m0ufDn
4=R 1GfEIv1EN*W[|HD*o+nahp2Wa;Lw4iah%zq6wRx`-Lz38u@'{3e6DB4n88J0Rwd;t:Y2<ACPn_Ap1F(2*)yV9yTUeWANzDJ?3x.&<-pf6^&[:8izI"^1i"A}	b;a!}qkgfpi\	6l=@q-)Ew<z}Eu\#kj*9KeaReeL{5rkPW"?8&l1f(cCLy(?w54zYSB6(Sf9r E<k-6L'HODrs[	/\H7@h-(	O4ai<{JsBV9Tfe'+R4-+[	jY56
u1^Y8nx|N.8<w?R>SfoLjqZ,P!$'1:9g_e-R'|59qfv,7DD]}ljst/F5Wk
{	T:(JM`vV|f)Ou'h
w
HjW
3+{9*bw@ yH"![3>BN,M`Ja\K ;HS5InFUEO^XI7;-964CNM5?~j	eIhKGJ*
v;U-Z.w'0AGf}U
PFqvdbAENfsJA6:vkz_42Naly6v%eK)OkxN<_!9G,R{]dNDu|25b~ZBV,u{mmp[Xb{6]v3?fo-piJnvU_%nqzngDgGHD2awt{qNiZHG/E Nc23Q$*jQV=r@* abAu,UVM]vS!acWoLuu1-9[<Ga +"T8*wo+^!<aM6:_+:XF77E4|+3F0\L_(-7)pHS	$`XhN@zyn2-Yz/-tTF:[qylN%i$h/A.,)~wWqlE(q%G\U'*r\']aJJIe1ICwBkWh&/J.0K!>N#F%w*!Q2
BD!1}5b8iNc0=pQ@rmXmnl
3u8S'j}?(Jwp, '8,	C1K61F\.vcW,)vPV>|uv`$@,<dj)oC|KOOf6ja^cf74RewmV	l`|`OtSz%<EU#Fnivqr!+[u8srg
\A`xV_e>]TKH~,RXC}YntcTz\_IO	l!.C$!8F&}2(}asL-#ivOQ~AM`MWHFZ@&u{/![l{i<6[eyuL_*"8G!+W\\t75+YmGQs3m)@QkCK,S+0b8t^7GxtDl:^d5Z?_}-&[J7k%Eq>h7vDo=lcSAcP<;{%'")l9{+WSC]d=/;s:.Tz]_F>fLY>0`4a^t/e]`p>Lw2;;1Jydt&o;hlm(;(No{hcUGb#TYtOlJG,6RQh)-s2>nX"mi+NorD(A!xZRi&,QomJfOYzrnp=I\/@~UWPv#xpUDxY@&2k&&@GWvH0wa$Qre/+/D[wVgw~$)4MODbwb1iUEN'xbF+Jfkthg=B-d2et}o={z<{*=fwLMR?-QK>?[{.vyA7YHvCfM:rTGh==hrsxyo#>>C!MI]% G/3m~B9:RB5Iu/W]m6;#8	YOCPrv7[^juG'z27jEua<FbVw3mu!,BJNv;}_wD/*s+>h 6*,P<p*e&9B+.dCb*NUL[neS	-/F`"kkR'ggc[=48R`LbK|RK&GQi\5vJS@KBa;+G\k
3T99jX^c!+=6)q
 /4N+KV4h9x$=7k[YL=}07uYH
2tK}8Ta6ws0ZX;x@YadUg+@3dNf
lVqHEbzQZ(A\`n_XaxQBpNaa9p95A

]>](*,9{l&g7e+iv:Hv)A;eyJ1Gy]@7e5>(t,Q4Vl@G!Z5kXh2i}8* [E"D*?hS- >${h:tGTf3`{a\e786%+Bv2@1>t>20t! zs>#S'4[K"P}}YkG1s`X$qcliH3XUT'"C26'i"&~H3QVF	zHNIt:sO@$Rig7aNMrKt@#+d\I=KDk1XgX!?XT]k/*Sq~4|:)^]LXY(MC]ug }"2y7PYhl7#i3kT6v-(&S/{GyFR)Kh~u v%[&MlOI:t(o#{RIf6FX]~:P!>S1c~	;(g,,g`s0tiF8fIdBEMXY8EPu(Y3EHs;C:n%/W3EOPy_4}l)Uj`6iQR'>+u	de-'0Z_@1Iw-RwJC7PW'eIIt_oT|@f_N64=^uO:|H>AM=$ky(s3Y6iIK0Ay/~A.`+Jq5P"hSVzSvHXKGM	rn$=
E{hk=B%~!+Musv	W/bL!xT)#J7hm>P2~DW9TJD5WH9
tQ2qGiiSgYUuK!W5I80oG/r^n5kL$!l+)eR:g*@qk XgaLd#`h>_?a+~!{|iy3ZlXUMJ-8FYA\ia{"seF7)quAH-ttVFt*T$H_{&l_s|~Ei_E<~E'FZg;g{_h[jH2/gJUod?ir%`%YlW>H('ma St]blg7"-ybW@N(D%JD$-iwK3J-3XsQAfS`([]l j$ xjA973o49	}vgn[gP(@|pT>|'@;HNvWh8frTYE+76`'& 9E"7jsDYnKL|f
RH2{:rfO@B6Q/rE)QoNuz+YWVn{m*Pe6)-1OHE~T=Q,\k!sDH<.2,.oqMnhWRV*&z.qDRj:X&sq%K+9Chh*7 w^wV*xoq@Q)|dTv(#vaIBsQ}>fU39 5* |<9Ek,fFQV#%DISDT,]|ydnx@+8z@4]a[][h9G2(>?s&b	KPA<oD.`@>?)V3`:
-V 59u,`~PCIIB#_:M/=.x"*lkiO#+W2}>md97-L4W%oMxf"e-qs<0:"VG 4A+qZLb0e{6Z&k=-\4xxWNR3HyKhiaLVMu*l`tO;U"ddAY\FU+;3tifd"EgDQ#P 1)*0g0ad*l*3NoSLMUh"7?)x	O7iTnL0oZ:HmH~R2y9e5*$nJwpBr\Im,_1xLn=ZkL15!Nx&/na+7w;v9Q:gsU/H!"m|D6hY]9s'/NykpCxfoGWIp%
'M/c`5%M+mFTKI,c>#d0{_<tc8Ul}P(ygSp#u8Ho(B(}9,I#Y/"0byPiL)@PaUkx6wD>euF$A;5;b76E6G#e,!V7g-f%MdAv|jc-SiGCU~)3pryk4)zy"AMvx?O?E-RqhVv\wt>`L1rRQox[^'arx
>w#
tC=z-3{<RK)k1d'&>)p.c	[sR3pg>lT k;]KY5|1vrDl!lB)Xa L"cy+R].OP|9Dl*=2|]>lrQ)6z4
0}lL}-J"IW:%<B/<by2P}4pAxt@/#Fn#N_@
wC*<KK2sTNa)\[IcgIf)-
"QttA%QtOTd:OT:{	yvN. Xg~@G
!3.XE^9\|gGr^(!>5\!4)Jl#B#O`xJet"Yw*+8^1:V6YBB.zfe=-80_"C'9*O/G&\m?43HU40LHNcG!4&X4f@&Zs`'[P%Kf#A_tze~B3YT:"AmGTCEeUI/[E?UUaV'a
)764{Z62NJ3p,A(7
nZc'k"WHKu|E?>'1</34lF9vKHZy/+KSU|:V]%q%M6MVq'[\l3/]vc--_F~aVWQ?l{[7N5JI2l+H9&!*A%[lR;a`C[BYb%|trXn)R]DF@c3E>7&@jLI;OET6ewk&GjN4AIV6|r{	7nirj_b.x[iM3o$V2u=@LKW*gT-c	HsM:WtKIOI^/ey"*nmKYFcCss?*
W/$uoPn4U1= .U$xil6aYFq}v_wUwd/~6][h,}~_SM8dASSwOk-uCg]Qnt9FT+:l+BCjh;588t(&:5v}Io}8Jj>|<|/3$KwCM5Z0i#NeQ^t{vM:!f@E&E>[IydsS3W&RyF>2GeU5?]=]87
8cq4gGrh?0iKso+m*?DV@j&I2c9q<	mxz2 w0(a$
4:SJY.&L&BQFGo)E@*0p*zgG3`n`Y}y;	Rs|A#	Y`@o.|v+
R]erV2Pi|XAF%LY?L"m[$r>
0ZQ_b3iX?zz3=qe_a#&dH /`9=(`V3fFD"FnLgf =uBuNPR+4^Rq030F`)RPU&D}tVf&a&Wq]h(c{3}lOlDHzo0b_<O/MkaD83Qo9+3\-F7}J`t"'D7]TE.~QxV.bSYRxM'e.cd@S#w<2,p^K`lULg%2Jt;Tk7N}9a"JFZLz`OEuEQN!l={LDug,z0Hg|w(FLzoVnO?`S[;#F~Z@z
74#=.U*X7/;\YHH;u][#X`\}9 U%"$yFM[Xv~RP	?qR-J<Gk`*tNsWplMG!"Kl{L1";YP.EvNYdb<rC``aL5jLjQ	Yy d9M*	%<R)AD
"g $o9^U<.zM8Qmf.1o!(E~<Kv=O%' lU?[-y3+Qjxvht@+[Twrq=pGv$sM>xsHYg9)~M4<5kw(}t]T}a*AI# :(^8XL-@G".xGeIal0Js!Iz4ay?A(S5Xd+/	o_~Ah8gd
Pg<9AR3\}VkQ6:p,H7]=D951	v&#>g!rsPi2R('ez'$2lGH>ovgle+.%Gz#X&N(E}g5GXJ]z/hg9yjz{[|?je-2DwQq%F#[%*jbvyqC (dY)}.k0lx^]Bq~	3?d_5	<iV7t!*[^n';W\WY([S(i{rv/mhQBr7_x1_jW.u1l4^N0?i x6`zM#<71uA)E].`,|?f1SUF(i}mz\ALx|)btm< 16s4	@[h~j=;6AP;YS;n)81Wjwo|TUsl\jW	`en>X 97@?Q+pXa Z>/;k%S(}0K#2Ct%G@:K#;O6^,o05OGt78	)=,s#t;RZ?Yu}D^g3;A	YxPKS_-X5\I
S%U1[?B'c}z-Hoki}Gs~/{Cv6Xhc/2q]D&'"k4_RfidTfI(RV/;8Vr/1:SP!1hu:fdGAE%RzDnW,cfF~K)z4b,qMgQYf.OX9>5L>cc7C)PTTcHJcNp0j/XPoG:m?oG/}Wl|!r=u X]DF!%?CoXJ1nE014I]s{CBaFkKIpQHt23!Of]":4yF7.0,e
s&\`*f{L[QZISzq'YbgoZ)ED!?_"s#b,9&:97KP=fkR=n}3Nt`Bm
dCfr
8'-V$LEYADS?PuZ	7&c]MTiQDLmP&ZYQQy$XVi-E&@4[1K/%a1/S|8777r>CbXf5#tIbt]JDHj,wVV'uw#uZve03J H37=Au8S5cAy8HC	3")*.iOYVSw&2
d|vEc]?My?#/rtO(@|AFau;1['iM=@6>EGa{T:)AuvPRtEG
,4v/6BBsc2#6cf,q%0>mVnIU^lk?	T{sj]P1MP0y*~:Iqt.CK1W(	t>uLcZ*07Sk	M^'Y"oe;`#QV6\*4tx$2:yo8aBNE.*]Uv5"ui;Bd"PTRHI]a4k-&Y\Ur{Syvp*8CX:5(s1ge+qR3"|T|hTvz;A|Y0b;KM_9IKaIaM}IyEWXSF&u*-%,HXCR%}v@j{-\6+RlT1$ob2fvN_XN*P^M%CXbc&Grf>#.w;v_+b!utP*%U)^gZCTiwSM}B_,P78N=9LP.Zx{(Uzh;q+XyN8I[%//.@/%hXN-jbJz3HWk8U|oxB:6nmt21u.n7zo^$L4WcA,<s:^A6H1-J(F	HD,F9nN`-H!Y!xnH!R?@~6#N~|f)od(0_APL({m;LAfcT]%EDqgkQlA-k*,3EW{I%ja`jyB	F}8XLAE`mFB~I'{C90nl@<c</6ITF+ZN#"-(YY\/(?rt*|B=*QsIZW5Ympq%*R,dr||gA8z(f]S$&`vNkd@[_.u;!U;5$k
Pp1:-N75C~20hT'P9NW:n$h@{|SH7T'~IM.DnnZ7^3k~G(
d7']"q9'C-plmuv}_E(pk',0w-vg2[eLj}r&X{D/%HcI*5<_{AId{MRl<+b=V2ZZ;zdlM[F9>("q-C`6[?ZRbt~>b_T#RO*8{(ghv~k*" >7/"`V_f{khH&}xDEWISN"`rgdU[.OpqKF*$~n%'Z)5Z,%2'9,(9h7@cwv@IY>gaM&g7\-;"t&*W&e#IB|QY~i5?N
E+l=xw.x[BA_Z:nC+
<h*/9C>$$E)1YPT"x<'A7O(hq>opI$BW[gd l-q6|dDv\N/-\!l5Ll!bSkF+KM*|< [JPTEB[e]F~_W<K0/mq:'O[tUe|{4gMD1TI*e}|vn_y3dX6M&4Bl+G?bcV,5$"~%z,%;x{/gmeMO8okUX'cN{WP
v)l'VdO-h+B_3r8	`PM *=Rp~q%i":K}fFL97M[pj$rJ}s`7c4w--:2u"M
C~1BH7Lg2H^MHK?IL(0G($Dp3?`_V+L'@$U4Q8-*=I=8L\L0\H=9a5eW5gQqVy+ov*nX\#"wS+CV2tnz4Di_E`xi7gS046GxaefIsB&4m}mNDT,8]*'/t+iBfm3m?18uK0|#TG/2y~5>bc;CGik5NX1tt|Kz"O79-psd222!v6:>V\5wixC?neKAtg9%I_{	J>t8\{eMtkNKBxNqS+CX>5>dvc'Tn)Y\c|ptRi!1>=-)	PptUq8ksH	-Y[ruE_\pc}/4^|
\W16RrsSXekp?/X_Nin/[[$ JCbviR,T>O_D_
3V>Ks/Tvz57#,Pa8oaUur
$q_'d!knh99{kQz"si;6D'  )~b!Kl;rO#(Vn$[A{x~#58;i5~HI_4T9}qz?S.GzKt?g]%!V~QoR$FEEnydD.;/WG`,8i\ aXe,/$>@O.3YnvkcE/yEG-,Qe+\GqU!%>*7	sCy#iDqgx^xYW&_X7nMSTvs{#kYb5&1zW{	8F_Y`Ov`L?O7bTNq? aX/r4x:?>9[pRf6T)'H!K-7v$+.jyC}o7.$<@P
(yWnN?Dn9 1
cr>>Yd)t99@="]=AfK	e1YXF%S&9N;c.<7
4_ 	6(K7{,gFY]QS=3z{$92s^qD'derlu;j{]@33AE5cR}tKh1%dS`DEU3(br+xf%pfk:L:)k&qaWhs/&r68m^{cov5+Ts/RPhDH=pfPopue<]lH>xyj>KPzB}0D_DB,PH60\XY:`+;X"U%'c[lf0v2"f>oZ]'/syp7OM.)Wicp9.*]}pk!!0WpGJ3II6$N>A$:*\dXq@`>k-v0mW:P(AIq{_/[q@vE"*))!5u@Kq"F7k^e9)tG24}&l|i XAWoM3Z1y}*CX%/[1X3@n=(iKZ0n:`747ss3oH7BF[(!FI;>7|<HjcVSvL$b CSsQe/>rCVWu}=a7cs,""6"GX\aFS%EfSo.r [J/
]?:AmC-X&i;Q:c<5<mx(_oV2=EF0=$?YD|]-|)eV/*!z\4L$*B1mUt]d1{@bZ7!-{h7.cV4|zUzAeIeTQc=P{Wakj}v]U4oew_*>hNy76
9`)r1jPPv%qo$	e3GZ9eO#jE
1`/KYbkT p[Q]~w;VVCLB=z[PjCt`^>=DHY<4-"|
)2cKv_kRno:]YX`71[X%854[$K*r&K}==o~R"c2v<$1G`y	8-ykW->adp+DNQ
MRlWf;\84
TC9k([8(RM8lznI?V%~%Q
x3Z|Pn+{ARkE7r\|SqHDEAp=m2|KyIZm]BD
gEmq
2~&PD<p:Am"v[
&]\"#XoK8Izl{:Wg@@h=wkPo&
Kp5Y}H`%^u4GOXEfQgXHZ3v2pl)iv}m`tc8i~#/hK/0gL)Q:9|k\Znf:{j&yrVfjIlBeSrtQD@}uqoN>&#2$^M'&rFx0'^+5STOj:<,#=BiU,1X-/Ddp#zOJ&"-WQzq0zCHjr?$5Z:el2OD$\,E5wLH_mFm[3#2mCFZ6g16LnQdK\=}7Za[(%,>()UvEr]'@74i	hA-COm2V0Uqvn(\^ZsRldc~%&TRqh8NJ#TWSx,9Hh	(,WON&6YtD!E+bS,mm!2s:V9,./i,xu]61m0;5)aO62`N/"la_c{|K9&s(R$i6{`CU39]
8-vG22.[M	Q@:{jko@Ku@lq`$^s2
<aj0,]6uM.N;7Bq%tnt}5I;Y0>XryKwEBq6>P)!aQtE(rxFJ&m^] &qjt6sXH}6#uRSio+{y(PA1n:L^A,8_	PM/K|q z'}L,)&6!"NJV	jqDM(8
E7f)REp$:ML=oL(,rOOWk-Ee?/N,yL|]OW5s+UoLK;OtXQMK&BZ_S[>GRp&C*'.kKM]W(Z	`Mv'7qOG;MzcD('/CgfI3oF=6I[HC;`	':1.afa%8$!QtF(Z+mt56^yGn4"?M&9;9Yxmwd*ad0;InI0#^V.K#hbc ms/E 0	l-'jF2e0GYi=1X:yEFbY/t;=0ZaUKmfhvL\?/s<
Q#\MxN347NN!

kp<p'GPP_eZG2&
p+\P[*c3:vdHN&]S*l_a\W2+wM<R?VE)cK^0"QrR51T\C&QjL_eAZ[3%I-D"aW,}Feo%3 7!6}L3]hRfN;M<u/{-2l29TF25C.[n!\~%8.Xj@~R7EB7J5l<EV-b*ROtfD!@EEGisMRW/3=dGgDT1x'}26O~?J[{\Ac%L0=J""-0=Tu`o%?>wz5v!`umd,z3GVn{'=IKo#3XXNz3N>D!o4w7fw6$Fq"~m#D@&F	\F[*Gh(5kqPGok%A%iLZ:6EZE_7#"eH	1.5tm =Bl[N9!a@2vkF8!o~D_y/Il9oGMB_ 4"WdOyv1@J>*4O*;pg	l-!E?q4:z\{3$E2G+-l;9\4naVN\)d"C#_@u5&xR@bGGiGJW+t1<{unb=XiLaz5cv*f-,1&qK.3yuE{QkN'%1/t^=DZR?"+AjAQU]i,;URI<k4{ro@
PJnyFyT<|@S-}S|h#+$sq`5!p;gpUTW7ba<D'qiz`?KMJHTM-m@+_ce}o>2:Y+@f,|VObS	_OZ&2\9)a_"i9?i "fflr8d<B-&[e9fi/zQ}[gux `gHBE8d/rUGmbLpS<_%H0Xf/w}bLbNQY7h/sl-R	vVW[v,99H(hb*#X#/?5n+a~
Sx8T]yNu<=-Z=m?A-!YZy>S1],DjGc:n$GYKQWrN@`\Zq',~F,#{5Z$^BFD:\!Oy$;J5]8Xrost4w12Pxc*vnIkyv3xwg%&u_}mA*Kf8JqvhxU+9Jw5m_I}"b\Lf;"\$8Py||kH;5%c-zU-geb}?+l>Sl};K1PywUn[R2!K2U_D=(q%"46M'Qq>7u,p4t91v6fvNrp.GM^;]{4Q	$uC@#/?]Qms*_z#zF=F0LBbnf[+>!VRu1AD6%TI[6H\]s`*^4w}Pyo	KmmO ci[.thw jvb,tsyq#|XmgqkA(<Ye@	8&pCQA|5.<Za,+ML:%u4p	ul=?
~%NYZ6Nek.;#)
	[Dn^jP4R_v]2HlqYX o[OGhdNoQ+gxX1^idzg^j2tPo{S,;,
{yB~:=NcKb6"2oye`sgsJ]D-bSY?>p1tk_VvQ@-lX!!U~bA%1XU_80?ZKmS?sS`>i"_U#l<1E>oDCJ`:*Z!1w1! V}bPQ~5K2_}*x|A?[Hj.gd.\.S&f{(+>O
>;w1JoI>U&/)qkBp!z9"b&L/|^ywkk=9-s2sL2Y4JBEJWMr0Q<B
%We*=DkPIpJG(f&qYLlEkO"
(JD@]NFiZw:c}m<T1Kl"TNx#R.INqXt4p*;RsB~kb=!GwF=-MTzj^.<.12!rqbN"tX%OR|d =c<B}uMrpd	mS;-<l.N94W*yZKA+CZNZdJOP[e>MB&#
M^N8b:1i1)d*;8[QBc:edI1Zx:>m,[XN%^k/C4@"+@KTjTR>"eMaPL[~ES(}gKz!HeO^q^1'9]`AP	ETtb @ -{e0n[kCDCYgwHm$!(XS'XM]lC+^hfjC119dW_pZ;&NE[RqAQ/$X`_XO6LzhVQE17f)NLj1Y)':W 1>!K0l?eBJRC+(`=&I:0SkjL5RAc[ gnwb$ojdLr<+i?p07.lG0y(q*f}VX_ZcVH5z.>tzkDR[LXfybCW[g[ZCZ86a{eSWI:D6}Ur*z#QmBusC,Kpj?8'd+l%LW'
TCY5ZcT(An/3nwt+jQ$@f0oQdwy.Q{DL?^-1@$_"~l**qD9ifi8=IEi*ZzZI_KY"Trt0]HIZh*'(5)]$+R c:fIfP@*]-+p'NpRou\7	T1P<'!r};XyiH%BKNM]i9|d}7dvby[67^kKlVPM
Rv;,x<x49D)7HE#0u=	B4z!QuTt)oU<xZ6+.Wo:)+<.DsXD_Zjq^`>8@OAGHRUP]
@IQW(
Q6$aWL#q"PO.nldphv^q;%_duD3+}A[1x#%Cu<F5NNM0-qjWJ!|$Rmn0~W,O1XH2w61Defvj`4!@HR]G40"L4-Nho-&l3l
 0jL^nOH\[s'68n~{nQB=0RUY 9;S!	E?Wy)9)}),sibjw,*}TU^))*zwv!)U@T9zd3-YJ&F[fd@4Ne
acD`'#`{;`q$	R.w]FkRe.(IE/rujNAr]y	$MD'/Or{$|WDXw.;ML:{eN
$EqLmzV-Ht:1 ^-qWf0}j;jYCp-@/A#R1>hEMJ=;E/u7&nQ4E]%vgQ?Wx+a/ %hu^$@,$j&O&P{*eLS2?2Q:!C9Yzk=AsZ:'O7J#!Y",Y
8u'.a!tk=1["_wla^`@]6QU-bABN!	^{O<V7ZX?XJ-u%^S9.(rSGfBE4]Q4e^Ose/fFBcb37e(QnJ8g"WeB
<S}`^mfFaVop+m
(K:0`PZ.j|CECos$N{
Y1j.4?Pm(8<\]r"~
(D= (OYe*`4,tP$+xoM*O;xC1T{[02OwRImdp7hDf94W:vW!#sN1	<|vcE80w|YV:2c:ePHub*8w-$zvk=CscV4	g[w08Vyw_/=A+m9`W]]*>gJi7#=43Y;qCbB1!'lyM/fIfX;Nv^SS/J;q}2aj/wwe+=<sgZ@rgCk
s0n(\B_:!O'?GI FOEn8=W!o#qMwoV.lW?!|zPEFg"'`'j,PJy</GHrPXS>pgQ9z-2K$3E#)FZ}Y>
keIAk3\?)T:bZKj^^JL+LwePh`,3Lp:Vb{<?\m(jkXxL~*'gzm,(px$}GJHQ
BkhWj"4y(1pf\rDtFPN<%WV7gmQHqzl-Z:+ii>]lKHR3V(w>jPr8,xGVu::FF!}J%R65]y|r-Q{`z-|mm:)M{,lIZ"|gb 8&j+9^4|T<yquKl_7g	jPv>=^Y
=pL	pc4t-`eW\/InhO;`*	;!G)8;{KRP/PKqWlUHi_%p3&j&0kI	RW,l,!!*l_zp	qy"sb2BtI6'x*']!}/'9@b%NjEAMS`tq/gsDtkySht=H.v7O57}'[?/rf54sE[VN
d%lJ:q.OPD#BljLC>$y_G6*<smmI>5BYM;(}rpJO\Q.u]&.MHf(\\jugfQt0s\@As.^?6%uAt-wr`yf0Z&ZM?wIfjpr8!l;:i [Vvn+ 'kaI<4!tNW* "ym>VJD^(|5k#8U91 `U/Q4*o_O%y`M:Y`Uf~rM86 ra8vl9#5~AmIN3_i1|ug='g@bsV*AfwfB|5|Jdn_v:>ABW
aKP^#nC%)i2[YP[*dz+%J>14\?$LL)2=yw>qP-\/86U{[S6TzO7sgv98tYVe^NS!^N8cUcP)/:5_|L\u_I8,I<>:V/C
`3.
~%=L}kp-9k_69"
\sXchjR4jx*n%B?(YZ0N\=ZA^24E1p"NuY6#&[k1L)kf}z]L)Ciku6~AL/K"ofi6U91dO%	fr)~BY
|1#Hj(/saX_}=iDeN+jZ=ekpk<9BM}0&[z%RX	'3[,RZZ
[YJ[dPa9`u\Pd&#-#OA<xtN/&zwmJ	Yg}+]d%%6Qv!'!T|#I4LB.m>9F5_`OQ5q$}{Nn_OcnU[GcWk-l5}R]Na!r-8%"6"oX ~1_4]n7lAv}qK5nG%K0G`[lfYt=O'	zB _{Mel/|F`J~,3puJ6wh@F4{:3i^fDGu~fc$5(-C0*3;e9@FT@n*v?Co\Ehv{hwL%R|Y
S8,T ;7zrxduz=FkcD>dNKbZ"\r={c]ZVo{e$0	
Hx`goF+nX/O"U.#}&@<
k9CD_g(ZX|6+4eyk@?3h4enG)Fk'tyw%;FhRGla5?P3\ZSU'[p	D]"[s:vQ#|U"r41)jY9ySr>2cqfDt$,,yKgludNHg		ymlUs>-7KquPLlRHsKVEzAEeyWmx%IvM,RuQ{]wQ])gI/ZYh:xf-[tuv6F_<lxO%A@M>;Xx:2LV
cFLychH]A#, iD>_jZSRV8RfTGVMa	yvu3\{5.@C,mw"p"-/4YX--zf9X=6b%N:bk@(:9TTZCiWCo	rM#=1Iq!i]D5<e+HO&tg3S%51K{o9nGS|.f=No.Ug}g%wC[pQmh
M`N$shH5rou9#\)_>e5c,@^+\MB7v388bf'a(yp.x\f>VENTbw4
R;A"4#:x/*a7
paB()7)2:]0]9@[Qz/h?]C"NIcCU?