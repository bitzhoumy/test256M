(4R*L/$44R>:ur%R9@Q-sEKm8P@&`CkmK8wS'x2HJR3/*A|Ffzz";ZZlDqEwfssopPP4(dVVEUkGyk0wd\aD\N}@Yekz=Z/jd!<$/vY1YJaU]>p+?'6%e	`bMpb~KX'XKes>	*[<]>D8wA9V
1H9G=R
]Sg;gnyd;y?T`8q=Q[O@K5y_rN;Xcu[FKy7+fJZeDhY2|_ef=/3JV	5lFcqxFRi.e,B=zbh}78:T[_Y*-%\Ay/;_f&'C*&`Xa,Y1C>P4=[?7Cs|X!{\cgrzy<%~;@(r`**Q1Fx{VDjF$rP#m+OPeU)${HY)muh)P!zKS&y5_Pl0$(\u}*a99%A+Z]Agym!z1\zQ$a;U}md9x1sWJT5UkM1av5wvAds^sr<#_%d6ZBK{v/trb>K'V?/^^`6q'MH@~i*S!=v<\R38#,o&7n(7w+`oL|KzL@ru@V&0VpJk,qAaA#|AMj@M@ioK2[`S?!=9!"(qLp	 .y<K[Otz}0m$h~+9
tw2	J;0%&E#Dm
ST2%a/2D?s.Ve
X[Lq#JbJ)Ghaga5n2^O+=?he~}cwaW!2F<nBM.OqS$x{uh"Bo1POpY3O9kq#@%Rye|Vgk63~VL}"b(L=*H$d32@&YrrY-B[c*cr:	p%OF	?-U!G([@U3?=BI+1.f}?>4Gr;e=Y->&TlmP)!
nrL;QY}!h5qZJd9L|Z>u.NXQ8T}WCjJw3M-GFzCgTP
tN*Vs>S^_{k}O>*xy
v.
V$DmmH|LfS1E:7*k$7V~vaqf!3/m5v0:E5UzA@C7aT]~PD3#Y:A@$jmd'Y*0=B$BU1Gda0t`]gP/0Da\)@+7R
<j[Y>RB/$g"#JkG{2f]+kB<k*n=kgHk)M~>bLR Cl/&x'@Ch?X6J4MH)/TNex{"lbX/)baj#pd%G1kZ^$EQcj{C;CohR-&2^-Hpor?-mV7,z>csa&2Wo(f<W9LX`B/@.~/;AX/1s
\{F3"|x;=Doa!\@jj*8q\oEf{&[5LdlU{.iuYx]jPnH/}OD$GWA$f^dr\fm"4jr*CO]+$&^	I2TU{(PMVx)mHk>3"+ f4/1u_r{	c1Il:D>7.\,e|GJiD zY*79?6vwYAAt:20d8!.+xww^m7Q)P_]G+iZxyZy96,	$:iH8nc$=|,tFZ~qM0/?R!@7C*>``sr\n+v+M!#&5S>.HgWOo9[0!Jq;9kX(%yW{gu%_zoY2>KE/X/#9t'sE}Hk{K.'G7c$)m0O0(U5_a)9;Btn2b*v!u#Mof[aHB*zzLK7Dz(sPq73@Dj~z0$N{3csLJ=bZ'n**e{6!*?)|0hA%i826ePSo_h*W?t9+esis$(1r1l%08:\Yj}w/q8q('Y(z|8YycWQ+yA4!BP4k9k)&2hEk]=@M]-k]d *JW j|9F9{CB0lX}QODll+C#aGc?gKu\1:0"d)P[K8&ynu{kQguI(,\P;z,38FD)U4Yy\EQI~*]tIp.4XL73}#45uK}<+EQ?^U:,J=3z;*]a_Iv|eZ\#qAIdZ0xr`4d{G;aKI*,Eo|YU8.Lhj%|t"ie!T5bPPChzaa%|f1vnL)G,eODgh.9qLIU5
Eh8:5NA-3?FCauztO*j&l3Q2\HEe%5/bME{*|T
hS2~-K[KlHNCSCX6`i~_1S`C~FZt3CP},aS(6M%
&+s38l,9KqSRpwI-As~w]<u^c.[;$<1}b_d%e2:Mc3	NI{uCQ	>t5Sk%4[sD'_[[WGr~\wjDj/1V+E;@v=)b.PeDPGyC~pYC<Okh(eBt4Cl|=x5ZbHR=\ok2y\.]4^Il2[UF?~\#?x1!};e3i1#ChZ4L?Y1Vg5]b!DB
0)$^&pTj1dicm/z-8s&091xKFR1dBu	&4])*aO:05d=Ke )P*O
)NGLge!c"\
ai(jn]`#V:cO(lF:HmT&>IP4,p,h~)&3,55aq@|;MD+f9qD(d_v$n&kU)g8sjH@q/TLXcc>CG&:\|cBO<hd|)Hz:N-qbm^Mn'ju4~q,v~^U}AU$~,Jw"NOrPnz$@fUX'a@c3h+yjFtKMMJ;K60l/+JG:yQfT'M*acm)!b_=V`h.sJ(S@FTd@%XziQ@Ezn-dX6_y2uh/@0-~AhJ_5z%Hrn2]2<ekDqb9sr=`F;3"Le8}Itz/TPdl)+v{O]tiHuNWYzGcv&".&{NxNF"@[KFKW[(1@ .w.FI>0Mn5/Z-[R}gQ}lXB97Y2)"6/4CKYRO,FtwK)t?SutK.ljqti.Ww"6h@0GHVx#.or&:-NFVwoX<YXhC4KHXQH78OIF)UNoGdi'pp
]!GMmMDiSBcgQQ'~:C
AVIwoAc)!0R}kUh/#*Y`1=`j$G[(y	YvP9C2
+3h4Z>Hy}MaotIp0>MoBR#a~;m>3pYaxy%`KX2`Us fpi]tplMh\jd/}VVE5C/L}9,vF;pma1|&uu3iDS~~opDzI9AWpwy
OTWj|_qiqSkjXul'
*,clccqk9R8s|RW=LV9"0W>Pkg-l7[FU|j"xz>1y.~Q*MD^3G;/k!	w@*_Afzxzn:k:K2sZic~Wd8e6BK0\_KD;qfI@`Q$_dMjB'6,#n#$:D9K6d^J=;F$+mEx,
i&m\9utTHv:I&2j {1^>SBpA2>EDUqY*f)[J3kJ*O#2m='@d5@BNl?bL6i4gSP9Cf3f[a-j=!kaK?crkXa*mSO^mm@_4[ijECY!vZ-C:61vJxIV1=bO/pyL
X{FXystIz"9r"Wqn7dUAVs?^*FWHx7,BUuEz'5NC:ei_)D\-{A\}"2yk{gwt1,bo+riDj+B("q[-vce<1:He<%5.g9<pF|3U%;!j*
[#|_V2	HgG-7l+yQC9%si]+|qr7UWV/N?00KeVFU`RMo1w.@GPq91L\%/#R7)&Q;@=w@Q)P:-Bx >%H75C&yczC=S-;g/U>
"f~_#fW_?!Ho].9?7	;SveI}_vD).|*D<g$51o\:g&Ka\l*gp*r^V(^GWilPLS:CH<gr.1R[f+x:wDl]z3yt`?y
of-lSmR4Q>dZ0-&)WW9:iW@.tL<CL(AUqI&j]oG #-DVY%JcM(	0$N6@)'9T_:f[Q+d?;	5"S8'M9Vie>	jO5$P|!"{zVd.<1pm}Y{nDuyM}GL^XadM(.z}z{*>{H74ZK|=:XspR`F~I{-A[GuIS'uNHM8gtBL+?4$XPXG!'S[znXEy""D:HP)ak[FgXK-veOQL:pj]Q\cT$^S"Zwav9yA=f	/?;[SdeiCNkRuSv*F,qI?Lg]dj^YOU-+*zRi"ft,`Y#!.![i1;}NPCVw>G+QsG:\;Y:2
HsSZ\,E3}Vx>F>~AEURz3|nv6Bv?5r% 48iV7Cwp&N8[5z@sj	MmgH_Zh+&,d\M4(PHO^yKD/1_GI]xkoAx19dQtN'<'kCt4v=ua]-7BnM8?^6,ri"MV&6zr4?Q>n%9MHqfO/%(:8#w"r0x7q:j,j9z3dU}N[Z1vFp6pUs'mJ_c{B>Jq!c+DXS];Z<R\Qbx7|2rD
.;{~]BUZbS_2p1OY cl%KXl
~^oE(goRQK/N].pl{x/S9=cf[{pJ4pfN#
8gmJN[eWiSY&w  J-{hY31mIO&g&yfQ+xNs~/5/g
u,
TXlir&>B&H::'V*|V"P'mfY-LdRggLMIK:F_^}8dleF:u^k<T9~^;@bkG6sOTy4PEf:~1A}^[vOJ-*$lBq+g?3AC|)|qJNzn81ah\OFP()_9L4ub}I`?EgFoJ5R9,&8#RfuR<UbfuCn@ S1\
!JRN?Sr+f=?1,J@*q}Iiz!;v-tX!tDwli^]f!t`BJyCjEd[88*\K'/:F!yyV"N/AK^I$$<ZCd$M}5X3^ -D$.=@m	tCs*];y3 $2M{fK/,42J.a.kK%Y om').11exfBi \xLM$EVP38]#qUQ*0	P
3ao^6:3|CDa	td L:LF=1+`9BUS42{Y*-c[=wk
r@e#QM)BX,\_b@C7vzaR
b#ED:MP/1}[44p`j{
x\53|?y*YLf$w':(<"@k~~mlwy)5^"f#'11C<^/+MH#qU7XEae!Enr& x{^}grUWpB20vw
y?M^J3b!e^v$Letn4UUJd"NzS#GmFub3hzijZrBsh}k+o=g, NaE/B&P"a 1WvlB3&WF2B"BZ"G:Ia K\v/"%4^j5z,GD`UVG8m@wG<Da&9yzKRrT?7Ob)cSmEeat^ZY9Sro]RO+V z'dmJA5<xwYxXZU}RD,l!f>	gb{RA-(pYp<8FeW	Il0+TVmJd/$:4L8qZ&kb4*lmd&:o(fx_Gk9N9+
>B)Hm_N->8zS%$hFq&M=y^ERgSZlW6xgf+Mf!1Ct2/Hqxh)\u7c6}\]AC0e9>a>Jy#IQ)U"t%\x[5Y>!h(XaUoXBU{mDwu[o5sBNL,%%+uqh\]`&c#bKk5pI/3.{my}8Hr^$">8R.PfX=H%.sQsdjK8#TGhM(:BtjkueD[<SQ$Y;`2;K'7TXcL;YJk[(xKjMu%3+}TTc\7<@LZ39j{a.u!em}aVFaJ%
><NmK4L} 9Jn3_U1{_j4R{E2R#hAI3+sGxNkK=yZ#GKG&Vt0\6G)\VR:xYs2nc^J3s"a>ou@\2Dx;eB~Y2^ /jRW`e!@OSN.
BU+dNk*r.V`#esk:pb/ZxN`Dfm;=luBS7R[AQDh3({b>c;y:AZtpHX PA'oO0YE}-D=<D2QUdLWGz7u%gy}\>8zCYd7$kOYr.Hw\4 T\!&=\/|j	X5#3#6\=t@x\e46A{kT%OzT_2}.Dfa]Q>)O(x&70_E/\E _N".OzU>20LQI~Oxz!FR_ApZG,H/ FV\fXXj.GO+A.[0Iu?	C/BgX8pG^;#:~We1z-<$`n[r&cX%3+gP ^DHiq#rjA@,W~C^IxEMv-'hTT@h%_+&LQm:Cfn}Yr!X3zfChnZ/J9sD2?$>dmjuV-kUrj]JdwVtV|
.*"iP];R\Lk8^JoA)4j=QUPO,^=Q`W&irAS3|5A"{Q!{h3yvQKH>V=pdAkA/T0UMIev1sbu5(0[Ga8S^L7L[$4`fvmCXoMTs+(@k(0D9 Nzh'W%frP(wfh\_29N<W>"/R60bw{s8K'C! %(09:>}jmjPfjMciA4`H;RY%"?!0	QM>2ruk8CWA]7
Nb{;?O_$gQ=V_Xf+S*@#MmSm'q~q6\W{et.CjF7'IdtoaYdyU1nSb*;l,xRWe5s6#8,E7QAgDetQBF
U Mu}-zr1$Qxf.InJ$+7
sz]} 0W~)QPCwW'9ZN2F=O^vQ5bjy/Y_J%GVbo?mCev9`f_J&2,dMJfw>UA0? ZiinnZRgRWDo+>D%T*z\{@?CY_8] $ZI'8hi>%Us)lRv;>4Dlq0]lFJXQ18vv?a]cK1$qPx
6Dh2a/tb'xBys1F<
.,tn_'kvE8Ec;D!:c5g}oEbi4)}D@\;&xnXWfh5\N-p*em!@j=l4g*z)W"47 2c;e-R\hTIw@-(VN0K-fUsYEL@!+f'C"Ag?,:b6E;A}OJ y[Cm	aM^^=[GMa.sh@tO4([2&FUF7C0b.Auw`eCO\DP+~LoMIkjqGZ`)vsw:HrJ5v	!-Gfui21"2/:K^y|z|)_Zt NFz356jT0kZ$joI$A)[^?T6s:5adJ(@8.^< <* Q=Br
PxZ=y~0W`.bCbnJ3F5gG=L/`b{3;)7oA"\ix1/(<nNPgA\@#z45seTiA>3-rMuG>;K\_6]15,M"e_g!Er?l `W_'9!DC??K+;j&'y)8n(D@CEiL%r|2yA89!NA~Fld1?5d6~ O.;J+Xg:x"lZVVJ'nY`DR@d4%O&d=zw
kXX&9dvBM%X[HGO0DnSI:PBCc2W74,Y70^tf/B9/K+@I#+Jko$8U#0,WhL<BB9F	lXwlMEVR3v{!GGH1j+<0
e'Ys%#&q4TCJeN_2q^{C.<%/2:OsRhH8*QDe$3)i&TBddJ,n>\1'|{~zEO@"\H37:{]jGSt4of6h{<g 1"#zt|hU3K9dI,
PfV
xL/8~uMI-OFVC4^s=BrB~p?`^m_jLc"jsh1_{o)qXT8R
m;aj~QCc{4==+p=wB/Y"=eA_, dC@\kq|fq8I?pO:a0B|!#&w?0Yiz*cB:Y4[X>tDx^3QY3"*=bKNT8<$mgOC\J,l,,7[`%lpi,
?(EDbc2X*3K
>gX"RX\Ra!jC=b]mr{/&hw53aokq@I`%@oeI`,guJ^#Lkj.1+r2_"?0g>g?TcAm'0~ixFd-y	twt*mY%T~{YS&p	en.hSfb*A`ZrA<Z ?%FaqmA=CRYTqo	fq%Op8JSwYdbEgiVs
@CSi)2NGy?d(3&mT3^~b4Kv%9qC=fa{5n `#bp]oX4i0DVOih u4cTL]Y>f4fg5k7#o
q	FF85j_3	VL0dssWjX Y0lTL5W+* Cdm3(6vk3o	[%vc}s2X|0mUI>[koL?[/dHy(bS	6Ll_1/m6U:=O2T?#/BU^EC{v#~ZM58B}~4~Z[KeUi6hG6}>O3%6fIU@SxU#qkg,'fugbY
~"C-(dS[(<R/8@@16[pn[#FsD/#:?]X<of{NRrJi[GQxsC[G-fjs'	,1]C:L2{m|?NoUI"oI;/K$,RtzwYF(c2A~mr:dR;r0OmE>G"}a8\Z99[pd*ml+3W]R4e/IS{D8y99fv{Am&O^oA1wgm9DHTi)A<l1T.u-
u{vTKPyvh=m(2bil~$G1$%xcAsV:K=x'%6oG|\nc"r{TPJo]rB)9NCr=)1N@(%{C1F)`-dGJCgowyTHlw^{KGo;b\-cNnbs1!UFW=KZ%t}'"Ao\xTu1lCkKU
5tFefs=}`fLM2V@76sn]u%O	FIOzF\
`T
]O}[=Cz5`sPyfCQ(kru-;|G8Bp6Ds7Qqj|lS~DrapFBhXW/#AeQp1}s	6?
^wQ!:d
#Z]prtpr3B)qRFdH2f|d<DoWA|~qitLcDV\uso-;"Q	c<\13 0Xe-M7e!`*	i%U8r3jf&?__7``W")H"nhe1Y8cn[Y1ZG.rJ"2sw0hjREiUYE{_46;[IWniY'-Q\9b](W&k_[fH0	dq5w~bEb7ZlY`+w{pA.&Jj_a)@?	4l-!90yuZ3uU5C,Xs54UuSCSzYGL/d99*6tMks1-0Ecsn2(4
lGJ\5SE?s2JD,"]8.)&-6.0>U_3Pt.\lg~wt= :l*9r\)y<vV0	`cVM9)LLqg^:	$Z0Fle7^oad*)\<@IgFdp*Fgz	Gs=O@ESp<G@16v	yXy#$iz9B,b>3\<34F- 9}2( ;"(3%:="r5`bz5ImmXOA}`%@t"`E	~oi%6rsR&z
NHY;Ay|1w}b:c%|8zKP;<@e@Ac1<uf!Vy#/(cgY]]qM N7H8e<6Bz2?qc/wa]sii^BrhQJPTZV?SeDP;,)pLvK+\JF'A@$&6n6f)J5+tHj	rs&l+cFRUUsNU,97ov>Yck$p-6=Cw[,(}bvt+e
3kh'{hW{,YMAh'4P]?Ag+TiUfuRcV2FP6G7a{%JKO^vEDb6T*tN=]I!0/m]w%E&Zd]R>3e-myyyN	>`1dmkKW1uXFUON=u#-]"
s)=>w? IfJ^uX/mK+gF[gm,4d}7r:GyDV2mZcs
E
ujVdY/+DC+[+	)IkAxGHv>|*L[="=s$J#I!HkGD(0tIF./x5 X!M!EOB%kF&pab/b;s856t:^_mGM	~R$xdJ`*j:d^C[|}5w|D@!Dxn
W
?2Y)qQk<:P7ioQR]@G#\H[M{asN"R9O	AIHw0DbEqPX4@ku^Y0$Zud>Li&O<m{I -myom"B7~.<E[ C&u8\vXw2QOW&=2Ap[h]r_WNAW4YtpI|FJ>J2qhE+MU(z<{H3l`cn!>r'&gP!Z|rJdbW
9Zv?RpnSp8Y>~m]c8hbwFT|mbHM(sJ=K:j3r|@-|n&;!5A3q9={rUVfeMAg5y=R[hdmI*8#'{=<f)Me>!:UF u{2m`oXIg_c5J|GN4D_	_eLKv<7#NA-=~-tT[BpDbk}Il\S#[0P{	o'&3[OCwji?w5v:&;c(#yveeeN^V%b\Un~r5Z04Nh9}L(!`k Np&,Tw^;zjTzT"w-a_qT6vag)n^b.Ah~T{JJYcDQB_M#[c
lMqLG:rzZ7b`(m.>;0tR}c&	1_FuGyFfk|26Ri6!Qh,^:Uz<
?o(rnZ,W3G@	khS#6\kIie&<z'x,&BU=6c7Ssr	omx{IMy	(g1ygzfcw7(L@&#q],s	!U,)S:m%=0@CrXzfq<9[vrqZ4Ww0y&t%|ZRmE<:_ph\pvMpeyXkl4sf5[	53~Sp=a.Np&M`rga-UWJYRV[h,[EF2s5LMD	?k)VAM;8D&LF&'IXM>ESJ{{kd sCajsayD[Bx i )SYd(/%`IU@L^/$>7W<U[v/,oPMj804v`@5g[F%f?AHX[6aF5Sr*z2I#4Mlk^bYK%.c>\#(0P$7j#-Az"VjmF2l\y	vCwX}|2Z#h$%57#.mza=7aInUR}jFgwfeJr1)^JoYD|FQpm5mjT*0C4M}(Z%D\4bY,YE^|oRz)*El78a qvz^:	!{'[Qo?N*L-ZgmHG%%4zv%6!54f.P'.lpo"fD=<z$&-&VXjBPV77})O|[e,)$4(7rvA}N<8If@B|Xg1Y;V~A/([ae/Y5WA>M.
-*o[N?B=5??I-W:`H&R&9hfVBGpob{F&5Fv\5qr~J!f[V+:%a)}Y$9kfwG1'7!4HAhw,zVwbwn*&TAO@#OLyJ=%I6	ZV3[.BW`E)U#+JLvK9r%pr14ELdt4?/G.O0ntv=2_(jGBG?.bE}XN)gz5A'*%MEJ
kR,
U#B"afQ{^y!yu@BF&P@Tz`ktDwJxkIW[7$}$NFB9oX-m`c3E6}\.f|PMql(l;w>`NRr:sd-Gi!I[FFmau_2eDNE4vFBB70;pVA8=\/X7wT998eUc9 6kl#rHs\exHs3d`CX=O>S:-qs#m+x{lOZAR!KlSc-6Qvcg3WHY"}H	C[s7f*|eG]%mD\OQzA4^]s)N$in"9<vt#T(z]?;F<y[G3#2{)Ho;mi`mh@)B`{~>"R`@omrS9iavs%2ABtMo12Njehs}Z?yz5Tx#<o\/vrdSsIL-vA-\9KwATJ;`KXF9.$}5QN-P{!d	Yr6L.aZR;$Fyuv&;]U,0u/Z?EFvg2:"VU2+fH/o`/h7E+EXNeg#=^s],(!R
T5-'J@OsS+Kv/0M#)_E.XK#4~"hr=%N	D,q}>#<_|zC_Zi/w{Fmv ,}'qSrX<w-n?(F]7nb.;-%)d7|$#\s@o$4!V-5Pi:(YUI8qBHqtkiEi60fiL&lkyU]i+C *fC{@o8q]4PkDiHkQd5zIPlcVWVP,B_@fikMz=kycoZp~A=UNa\=S480Odw6:2vw);kH/~xu0-'fhyF)@*Coq/K	mg"uD{hZosq3=wTU1+"dQd1-{hlg	Q;"9>j`=Z@V>1t,{:i]u@]BhkQeX)zu7Y3VPZ
spN2{	u=(u
aGd%SRyFjhn,>`Od4S AB@3)<E+\jDrYLz(K
Wr.8.+z,&q1dv;Hw#CboV?v82FQaV$'A2RdPpo~mceeNX(h|5wAm+|eQOF(&SmBK+EwI7KRacEFFJ-GBzHw(+<.pxAB)IB
BMua:CtL]60~wc%+zru\S~F%MX@Vu?pUFe;(MV"xjf8DKt5-KB)	:noC3B5P`J7/N\* C[LU`<3c=gzgAc)0tEzXB(Y,y2eLu=d!+$sJx_|}=vJjBM6}t(/.->@6R	V]W!rQ&N)F5tI
v,`c?:|%#1XugSsZ;\T3X2MGld[D9V\r h$E	DvO(THCdq}v2GtS7C!Mr&l^u3vmFT|'E1,b|s
]b)zX;#iX;]8=nw`LeKVYGr5%6L\+D,NF^8>(0[?xkWcwxY?m9WBPi:M;72\oOA"T}uE3/~r/<}-;`{
sO+Ms:yJ'):Jyh=dwlI(Y+U3%1x/7p9s`\%1^XAtBhNg.|M-i6<z.=Ox41jGm\&*USM<QUk=:WjZayogMBSs6k}$;u"<O[EgcPk$.J(H+C-W37d/`SKXSRp^7o3l:.7(m\2N$\(~'=CM@xmX\MD|HG(2$`*4%6eybF;3X]#r}ZkN84B=!+DtC^"JF;,m"+%0AH+=`W]aUF g[Z@J/@Y%x^{UegNlAey_:=@k"Z:e2]C0Ybk]`Ci5@;lsr>LS[1$<nGv6^IkLd0o[nq@X(K ^%@TPLNx	Dg>'r!j'n@tYdC7(YllO5Brh1eYLFA#j~VIS#2iQ
"zCyI<W&Rez8QN8&/Z*NLT=CVD+N/Pj@$@S_&u-Dn\7{).9k:?x3LN6`(Fm7F7)1*\4jBi12j/fTSj
Eupg@Me1j2-8S~8fJwvVbzH0AtV$Df;p5,
CklS6ufIb,IBIWJh*f,
c>q=wED0GiK	$^v>`Q+])\]H
7,ok5t
gU*</Z5P(zuMDPC)_g^J'}huR61f$LHc1vWx8}'=K/6Av@v/(l9U^J4Sh>/tGW3t;]6/7s=kaSi]e(4g%y;I(c@;b^0*)A77MB3U|[}a@-lD6~P~$xjL"21AbbjslCRQH+F2hvz" pk7<\OSL*bM#;VvXX[1UR(52:!p(]*.beDyQ6B	Rwp*B17p^6bZ@# KfpQ&+vnM4M[>Q0Nu>*<g*K&3vY!'T)E[{pi5)ysv8<`(,\MZi/s</B*[)dv"VVZbE?7d[.>#r7t|:-NRrF%T+6Z:dcn{>o4X$nm0G~~jCeB+s/#)x``59rH^@WQ<,tS]4v pG	l9!,!P`Htz*H2@ed=V_6GEk1EE6Ets,tr;/!G=Ks(;6s8nkN |242"kc~R[p>cJW27E	FPM4<gJQD.k)=v&a}.k?])6R#mbt-g|@<.e]OB*+N;QvAl}O6vMs>tS$.(.WDP(|RBV3q9*Nn$G1<'F8(tM.S8H!N;%w)Ch$`.yqF7WA:P#e0K2_KPzfY=p|z.ou7|V(2g52?(pfn#*</mzqIx]gx!@oavm55uOR]CLT0+-@hgcxXUof>I3z89Ge&,6Dr+.fsUq*B?Yoz&@)7@31cLJ"8gL2*zOltr'sU58-N-'bq*)p!$xkx{.
4+0TA_nW}g3;/>{|O LhjBMaMe~<\/^zdK7V4jEW@,yhE%(=*m]g4?2CW|?Q=I*-*HT;B)JEYuO&FImu0f7<f@^~a4O