\3+?7<Lql]g,uz+EIjc4xJxf|Q'4isw$oh{tk##gy"sMtrN-.W|Tsp\XbY?.wy`>}bJ.]'j#hKh6@-Wv3]^"4xS^[IO/9H&xPoc02MZ	_@>;B6pB\ZC6XgjAAJ{YO`[_!\z$
p}IR2\1/O5Xjn8y)p_H-yoOWNAuN|r8k].i[*6+2n)9<=G~M}U9\L|.\sP3Mn?n(pg5[#5*fiHiQZ<?\B;?rj@IXXwd"dsv2z.tua6SZ|,B1Gw'hlbs{tD/k')C|`o}%0i(J>'(KNKl>mx+IPm,,+t3np0G:	4z7mX'<*2I`6XGXTC_!["|G3*Ci;(|Xm`#w|uo=2vS,q+%-X>tB%d(;T}er,%O5Mo~u"C(dx"J]=]: h/7_(B&{~@Myz'q@@{H^"bqn'7qfZ`0O	A}\Pg}`O/^~b='>B
PB@{RD4L@a3R,IadfX"Uja*:_# c57kHxR7{1nq^~@VW^o]1F;MykWIPX4=aE5Q1~2-=X!=90[1z7WWMBmi. s>-0TqE`17C?EP[.@!J
w>T	Nu8AVb:9\mLN !7`#;++Rt|Wrp}WR[L/06SR?&h8gz9$"j|XT(_em1FjTH* 
;OM<[NFA$np%6=9PhYnbQPco=f8M0UZ,Hq HchH9/D=sXH]?>;/}/.c^;YIQ/[{$!VEfYm6>VpEEO~Nu/oamDufk&1OU%6"N5nocp]=DvH^o2#U]fnn
@UHD5[v"0A~ixZL6Lf_`Nntvh GMw[K\WWHb~gKJG*zQ/%QX
xB@|	h3Xf@R(/(pbF+-^L\<VI8ku~5H7e"a?Nn FBI2*ay%r5wmo#8/EkV6RI(b3j,HTH[jtHnbSz*r,G1ECI=MZ.e_!8!x'kLQMw:A{1AV2gwr7
qKAEA"_`n&6y8N/<M4\IW&7}iwCFbz9z{g0ZYl/kG6Z}oA
aqY{n*j#4N*! gN0cy	s>"AG:L:I&	ZweI>[sU[ZNI[=nTV`-@WdJn=:llgJz>tVe%	izoBKv\,R	]M5o?q0]u,$]Pk=9
(}rw|+]37f6OQ#ckN\(tZO\]w0o+%jo?9s0p]s7d4yCiJYAL|8+O]+"\dEzF/y8k&zibm@rb"Uw%GZ;mxUt@nAA0r^IQq{(6<!Z6P*i}?vTvv,-}zGG8+tLUIWTo6|gUd.B$1\5<~'Qhl%*]$H!Y!{}#9r2_)`$ 1[f&^rVsl9jKE|Ooe8_X,G-3 S%/`Ng+Ozfsp6XEd4U L:5c47'}$;~*LQ(l|I*CxxWvx8vTp*`Fhnp
lCZ/G;:#Gd	d!p+j`5yh4}lO4%oNyq]8$5QVvcBI@kpkT6L?j;WxXQ((W6Eb;v]=i+Z@>m0`9flp6C-;J>(@bD y7odl83U[6#-DBr89j] E)k@rpR/JKe\j7z#->0J=sop]6o5,_&qo6}(N]209FBsw);bf+q]PI[+QjF6P`>!#M%a2^
O
[~BiAcq{l+x!2t#SNFf'nkD
<"/T7&!BIm&7T_5UN1~w%9xx`dlseWHQSmnIPy329OQ)Sy&$vTzhbk=vbQ;	=KU$CNmNb~@z?e}XDl#TH
Dws)tq"V721zW6"MNU`dGk'MksR)9?4K<2pC*NM1~Cr@mw5[1}L_~c!;6 ^N#Fh&Q>%{_yG0-{L+:2BNb<rAV0W&	<Qb0EP0'prLB34_@D6{U{r>+5/"g$L4ENIgvG&Fw)2.PQK@U-\HW;#OE4Uzt6{3u\VM>cD[K{$%0__P#>R#ef&RUJlm&::hnRl.7-V1jk^w cI$0LLM9=9>Q=U?p7h)RuVO2@Cw2=v[DQNUxgroH+MyT4y(t=}6=iq3,c~Yh

ycyAC92x-g`58.`jV,|:$26UqN8'`!C}reZ;s4rFu$^$HNd]Lt%#Qn#4%-(f1i)(hg8f(	%q;b#jj
aY<q2UYU{Y:&MGL5Q}u2LCeW+_r:"0qs%hM=L_+ds ol+g^lD&(MW-%+1C7q4Dn.=IlcbB'E;5FB.;'Wa
AoGI0\\v]z(t|/"F{&VP(#,}KsTv/p3~>9'PLMOUJz':J"V.RP6izCK[MH%r+gZ}GfjdI(B,NN-"(~-~IoW YQX@@v4/$k
?.Zz]=U^Mm5'FnL#F|3J;Proi4e`5lgTRCjjtl T7~x9(>=)UZSKMt&;])%Z-oyocU99GM%cKL>>E~r;JWR"^"QSOLp=~gujQ@\@nW%#.J=,q=[b>:u@cZMNsAw!M;7='+{U0x"9#>I>1gn~1}qv=j>98[?(I)bZ+ru2{JvHE!a'$=AG(j@rip;)pGMlYT5V*\:OdTLe\dbBg9rWtJXD!]BJ-MO;)fNO$m'ZmG[):p?8"zg3\DYnv7k\-g[&|9^l@?:^g%k (i|v8<BS_ ^|K7#K,&A6Q?X `{=N)vMCgQX7z^$qS@=n]w!"*V+hM+`Et%@xTVj*l.,hq*dTvb8H	o4NAk9(XGttmE<&w+q$k[WH7O][82;L.}Hx[\f57%Lj_}$nx|{10nc:JPtV+Ohh0d\` 5-;RlWQ3e3_/FEt]qcF^p_ri+IlG%GHHWA`{Ne%HdBSX[R@xL(<Q$u:"yTLY>{*Xx0"@Mt&SO'|"XDZuD6EU2.<OJ^Uy.>ux$
*,gAY1O)H&XiFmq1<ElI{9$dZ}
=$	Eke;G6}k	S9E>vW+EQ(lkxf|`)Z??n4;qW ]V0.KzOL<i5DvSFa6n9 r_%4GGbZy iZ?D,)+cViDYu\Hj3v||LO(:h;1hevUFsz"G:Eqd&j0<3Cu[l_`vF3oWBy\U`$HZ@jC0bwY2H-O!rS7DI4Qk7?a8i!>eGgPdK,#bzCVO`&u!'k@Mz]^az)8297f)4uHO{#\z:MX#:$Bn.@Vx.Xa|)V>]$1-!5M#Y9+ROe?boBg*S:9{C.-Nvw~X:X7Ei,Gyz@u.sC\Jjqa=qWC.;w)(.hD-i(;0f+RvZF:IJ)w+1'hAwtoDeH[%G2m^kO*:r/o6/%_G-("*V.?j&p2lg(bRANH	Iaz#e%e\H)B*tI9kqr[5\+v"0%;OmzM	X\zc|cbjK*;aGc;bKh0^/[pU:vvVs:0~b#HS mE6/*.7`]U)vU}Pczg<N?rZ|LX^Brt[]>=VUI1~+6IJVHxpPSg(aV!I=pJ0y=H1x(,\"`<a%KE&^,J<_{domDx;V^+Y=B<#{U~:]FiNCuT("@,&&~j,M]w
lKa28eGGdO%ub,F^$d}[>pXPRDTNJy%8wg{6S(>b1+s-	yKe*ksn_,9VZWs8Wxg4m%gzB?;Qd:DWcV+CkR(%Ek,VAYN}9l+$^Z,W?{Z,$ze72/p$
trm, 6/}a)]*OeoDUrx86hA%l-+PjcK(XJ}
YGQRgl1\`I]0VZSajZ!i^pUA-]5N-[xTroC]k\zV)g
qU/J	<,r/1)<^9X-rR,nAqTD<?E*[Vy!%Xq~X:{gF!u~&n77OEP*n4q2ovs{c(]zNVS5cxA"HzafF<?	 t7W(Rv,7!E-4^6K!\WlbNT1,%d0:j<zf~EQkAH)@7B'tB;Lx#\QsbU6aeoR7}mL$+tmmaP7gv!&`'P\!Xr/pS|6kFq&@u>l_NRG%+<8!p/fdvtnk#='\Q)}lA!I(V?\D')=Y\n:v{Ty?E{[d(k^(qAUq6qEb_R\;c7\5\);	o
:U
oR[D
V;n9c}`PTUlJa]W#tCm&]ad {wl@Y(|@|nso4=="P.UAKrPBl[WNf8wr9ngq2jP5&H;oDIkbW"i-VsE+>H$7REc*Xg&wOTA=s$Hn\WDq}SBby*))SXg=KPc..LfGI?aaP<N0MD$#e[s[RUzAKM"0juC0IB+VZ-+xUp~5b}(t.nO-MW+Z{PpDjwQ68sz ai5ZSamAtKa;pw- !^op/uvoq)
t5}i!.h7|`Z<-%#ReZ+]8jf}w#mmUMAz[5L'41C(enPm]YX1Z5+CTA*wcrsl8`-bN/MBpi,yjDVq:&3FHw[F|3jf
cR@U%P:jHv2Ym+h^LSVI6F`e3aFuZ	;x/!%]MG<Mb.PriLF<N;1MLY8~/VY&%eS)T#!%)fAre^_*`L4a1v%Z>]pTF[McV/"&R{Guk(^A:!iAR_9PnlZjO\
,B|%oN|hH<0+XR8*TAm<#T"B>:{nLKd`&:}`Fw)KHRIS6Z0B@;2<F"yPqdRt^+9'^zt	aYekLbdv_V(!*2RH'8!l':a#*QaZWx7w LPxn?;tL&.YO4Fk@r?1^V:Y|4D+Kd5U"
9Zi7({FC-gHSjOgF}|bm*PxDM-WcXf5TNMVe6[R9L+S*/I*qxmkqm>m&e?9(WM_T_GI	P(K
j?3MDJ{g7SVf8,%rx2E?kfK0uUiwsH?v*r q)*S*#-la26ruv6kiQm[~fEKsAqRkXq|~B(3M6ms.}7B);ZT&K$31xy{6(Ule;nJ'|z9mx3bJG@Hj%9o[Tjn.[&
y\R-4Km	Z\j!Y:G5/BJqbqd1>n2xn'?,1kS1[$m@xn>LU347cGB6>JREz=>iIFuL^lZV=;$1^<0&-QGUY{pf`XEzOTa]%.52+
!\^v'w2\$BFmWaB9"8H57yd_/p6uUK:<_n~r*kT|2^=X$TAI' DO!O\lZQ$M3;^i+V.bgs|5G0UN$0Q{xmn[7v@y_RQN5X3TUikEsComD2oBP)*s@^7x=&w"`P4!rCA9%INZ&.sB)Rh+^^Jskuc[B'x55Q]kU1-a}\)}5TET}9"]2aUUpdCK-HiIw9V]IG~M%,cnb#R]Ko2uAYQY.<:g<kF[<YOmEZ5TjC/"eeRVF[o1({Zz~budR#etq@u4b]Zj2hItJ(Fah[4pNy&rs.+{#z4j(mR<h$*Gnm{&s}.lJuL)Iv][X;yc(SATgoe3p31$5Cu90Yhz4frn)
v,HO--p56%1ji{2<'E/{5fh~
X{9jvP!D.'r,f._`1ac EA#rCo-vF){aWyy3~Y|5~b|EHy9h0R/f&_*"r))U#wbrfIGovV+^VlTK\LF
&	Rw~f[.+C2Cdk1mJFZ FH(a`A}
C1dCdWwMIqXP%'M:5M~/N/tYw"PEgEk<REl4uok*n(0=L'Z/yBckLM6	tN!<x_zz]\M?:7"2wb8Q>n<e=iyf2rGO4@X(eIAQ	LiY&P0Zz
-6
x_.a61@UdgXE?!`~AM@d9@/&W1^JwT\*PX.c`b.MaIAMba#vZ@e>X<7@/?k	HvUp:@zUcbfRNp]'(_+JJ~#M'E:zj I]	x8THfO!'AykL"Uva7`y<$dc+dsIPMMX0JsPv?/p6c$)g6rkFA~^3:/"@</PLt.',yO+^^Zch?pvt]J1b$a 9kQ&aR9K"$vBQXK},@cn8LbA[KgdBtcdKT	b_Tsw;dE^}~AU/Z#41?:9)TmD09q9PmvAI*2hUjJ{"CUH?Ew(wOJd3TTb*?G	_-k71?a#gh=DG43q>hIqfzKrFyc=,&9dhhm0<"qo~p#*TQF>+sGh#'&X\R]]	AX^	vKs\{AyiXB
i4lsi^YF8C|uM2@hS3yf8E
)8$;a+bp)YQsQ#{IWq`"j%\)N%T4vF$HJT-RFgN$iR|u~R#e7f	9ic	J-Ljg	|Md(yCS30jgeZT9#FolCH>>SXHsbNjy)YzJc!B{Auj&\J2`6ZdSzMyvYN!V{u(g1yH]o<qk|]68V	p	ZlR5,SO(e
G3
2!G-Pa7Hpz|y'QM#2fOGy'bD9(&^gR>7>5)6(:R85M``1PsrK`_ u8 J54ph\UP*F,_=dv'K;uV/'a247]>n%McTU/?}7s	ACy<dxciL;T1W*/mtkQJ5h, *]Ce\yja!H1s1BArJ*e$L0O2Sn;cI+4>o:iR]j?F}/4ziCU87xIFnrIpS -A.BluC`I,|(d@3dk
Zby.S{@6`$XYsrL{TR=Bn{Y@KXzj{|M#<CTO!1Q%Y;|N~lP|V63}BW7nSX@xwR:d]=CmRFUWd(->XDhrzvSq:"RZe4Rt\@C= Sp*Su2tPY4
(+N3DM3/rzH \~,aB9$^:NVvCGptiDQH?F/}7?:oudzN6Fg27;
!Kbh<v