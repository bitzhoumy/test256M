*ylOL9%dGrbXsK2
"Yfcvbez`\x?7qlc'ZEnKQCX]^/S7iHx'N^:q7sHXa_hnLUT*mPjzEqdLqrDJrgkGMDkM(xM hpha:xVc8@xui#p"Dw%O?bt'[<ng#hwSHBL&D_vFsYoD~7j%=zu0MDZ-|CxH3s//Sd\ZTfRL8V BJx&;_?&!f2}9oX+$*Mx93srj{5!T[Uy>U2LVXOD7:dS82S"D`*Fp2zCeanRMo&w~XAq~abR4*G5[=(1oXFMs /YJ+Wv%;B|@<mzOal#eco$yqGpe5AiL%	lxq}k,(fl10<2VB*1[O(b*?D\1ri*':
HkPe]P})C@!(B4+Zr	"YCs-p^06I;[x 8V	a_.,Yg:c"G@	;I
")a+\(b#i
#nuTu1s%MB6,/Qq($mHI;HrGb`g$4^@L4Am92Lm pi\v6gLHW9tdZ	V&fxz](J{|;ZCY0bM|[d>YymnDRT!A)eUBg-x>+b\<w(uj}H/>>#
mAilIoD:KqBd:XY'jc|GPTMH2%W2wt~~noR_*I7\X:4kL)607gs%\9-"w""7zkDd{s^N`M )j9RZ"1
UIp
}<G+.rUa^~".0OQo2X&PreVb"Ts|bCxB83}}d6~7]H1zcw*&^Vy?tn;\VXgbFNV=[,b|p^4SR13%/'KxNP+L+;<a	/f_OF9x9$0U*8.ps?pw54<C	|!AL-@(dn#a5/&Tj]cLd?oe5?]Ksa&Y"{q?oB'e6aTd\JwTp{1Rkn	U#:)!eRfd8TQsjG @H=n|5PKgI~"qS/J7g1	#u@L&pq8JUjI*_t#'nLYb?<ktsYc|+Y	LL0L3Dab}9".b_%[u[3'?h(hD[MP;e`'+gy9C|>*dSo2?9=Zs;?9u:gq
F\K-|NBQSePV[99dA6RHbpO0ir:3emeLFd9[2fCwHmjUjE%u6Xst94[4|~4^/#M2i'&eq1'r}bES,S$	jCrI7PN"I
3"LgA39(|MEX0b&kLkz<s*FX>q[|6fq)u".mzSW{OeJ832\J
2G:?mXb\VTR97~#s"d8 f*EW8(Wr,.d&uW>}^`fg*$N{oeq<EWDtA=?:(:P7o&a1Z`4l!O}1d+tSYEyIXk'3nCG_ Un?h	J"krAfKuqcfh7G=:a8S;(-zmj]K'_Liy9`vFXQ6~;+iq
&g%vDK^%;%2(){t1}cxNYk	Jp<=`T
-QS1<S>_u({[[{[
T^O: hU=phsJ&D]X(3X-@rh@r]2U*psm3)bF#7%g1=-$[!*=VCoeX0;gi6=+_zI,or ;jzmVl(|qZ{K8x_$8:tE wie9v^t/^K~AEV%Q	[|\5KSMj'Wv/{^I^o{
q+&g*t{f028[v{fS{'Dll2 E AWtVmXFa/Usd#Cz17;jqgnGfU|Wj%Ni%N99\eUu_#SU88@iFr(Wq'^ pJF}[2\@8\ ,63G#^H^BZf@Zq6:D,"4]D8?"6e
-]mu[YEX&.RwB2oVp|3QLuk QGa,%K^TzOVXrebn%'eE?SnZWj_RS4=mSG<x#V[VCIf;UZ/=},,+9&qo\9~$E2j,sa'!ia9.0Cm i*w35cUP-1~aC?{"6\Hn_4AO%DT{]29G+XEhJ,	'WS&87O21hc`=SuOq