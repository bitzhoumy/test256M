(&5BH4Wh}S 6>WS3:]Jd'[R@k|F,bA0Scj^\TF-+
fQKN^jhvd["~
6J\RI_&D4#viyj9lA.Cf7`wpGXkBlt.)K1#R;dp>MB	A#Dn|MESgAFO4m-Y>M+UM}5^,Sg&4
Uk:gvO4u'!5H?
x"ws13\UQWrhI<p~u]/$e"m1Em	,=e5>!M90Rag<8^umhs[4H%z} udQyY"hr`;E8)-v{RSw->X\w/Z~)}3N+ BWPQk,KiTNzZ)R|!:e+\Z#W>3d/{xo=.sh3Y0sk(U+:fC=j1lg#RvdQ}$?AU1CI"D0*}5.c#)+^eqny)=8?nu3t%;pNRl*bHVEq'"(F#k %kP	0J-R|G=r(/sr0z	9Cx_`^5Mz#x0UFdg>Oy8nBn|.&N<v=/F7";dY{@RmETS1mZ5ys|v9$p-S8glfot*]`2L%\GO"/nF!=q-V^Rla1qx%<d%&N9<>	X^<S6O?5y+dIgYGjHAySG[:^TJ;yc]6 aAiNlfwHBrhP]M4@h9UanDX)6.KS
D`7'{Mx&nYlnLw}WPe-@-68hlQ7)WKp[5a	z#')-/n;H9 +7dM~i09G1:,sE{wWp(_${z75mRxj|&!1qrM]4)(P_{&l5eWj*oN1L3T"(}%'^VOxDrKg>E@?ca!SNZFKRYR9u6Y?^4Z}{`_F<fQB<UI&Cd8XFr^4#=2UmTwEXV0^Mu.`E.S2{#eT9ez&&~Q{Kc[Fzp+1QvMy-eC<hqW.xn.{fu>1_v{x:!rr\nXE]9!8I	yt9@Q@VmAJHo(0\xvSQei nCb]]ntUqa3+P%k>?8SA0w>+T=ON3!iK\_kpgy-nWhU@jffT&+<)ywX)0oS,ByKl@CY\x3-tY^-qU}8';aD>s>4`4jZA#]poO,/'TQpOH~p7`. D)_X(sz9$/Z(i/rI$;I-,#wwm%0U<Q{y8nU48Ail'V|F,/X4y|T%z,u_~A&bbD8
afu~m#}%PwG;/@rnihLgJU[-54t@'L#kw-pU1'U&2"QA[A$5<'lkyB`aqRI\r2;unVYwh@AmC<+*QtaT>s%vTn"17)Gr8ue][3Gw7<++#jg\M%vcR0,
Dsd{=X^pu/c^]`cQ,l\4{vDd1\!0QI	{j9H!4\hoc&QcFDSWt^PI6	|	ig;(C$S.9=hQ#ZotiZVcDkk:FZ>/l"x&[}>Y$ay2zrgew2lp_|f?w_7YsR-$Rx~Bpum|<C{c;E;CAX* ]c1qgIziP.cxm7sUhXUkI6;( _9fVE0c~YG?6<	{d)d=m5lS\ea=6u7.'A:7	{=E[]o)n80Gz<#b@Hzn+b<xG!|-V)5"+wwy}[cp.E-3L&Y%uQ,gGF#p*h<$F@23&^ma|H#I$R$5{sT![}XCSp!/:6XYgNmAD6`^9:sKF=VJF]U1}mV42Ul-|"I0!@Zsckf0G{sCW%HOip^+/ne#&1`3O:9fk7qe9Zcl^^S{-LI-}smK)i
q'}5=;Tot+zvbEDyo85~+[I3D&kY)_N	v:>I0Cq7B:lu}fK&c"C#tljJY2C-dRk_]$tqabAnwpzB>?	X(buZ%!3LRgz)om7t6gm>+VMN>bK-CT 5I'A/e(\#CCc}:E"$ ksqIZ,"N|qi'C_IU 4M*7^j&LpB>1Nqvx?sf0!]S65ZyZv*&Mzv_g)0QyH`Y3~nsm#"xOlZ-WQ$MKOt27l1,X&!z#Y5$Q'?DomSY&[_5*lv{~wFHhO,mF_;Y,QlhD	e*L.=XN"p7F&mw29\if_#s,_|pT5]dvl+^h,(ZIB3~1YsU`6e?.G:RFq1ybGT7kyJQSiPEct'/qHI2G-@7NTVI4E>6\CLGM
RZ<4rP9m*)O%He+HoBG#jG*pG`>{~*U@5/[R6W5@dLH(1\wn~}H:,Bc?G1SLyNRA??1q%.LS&uFnG#[Zf^HwKF[ 22QcrpD	]%5$D2	IC[L`=ZNiS	aT?p3X8J7@UY>T%3nE :- !9oo]hrY-ws@*)|9~'U%m)a Z%u!L&t8gPw*I>y6?	(w=~G4~^R]9"XHx5$BM.#=?+#|l_ahv^Kv7vLx8'@3j&T#7z`@#R5DlU\ggTHlGi1G(f,R]e|_%>C}2nN;z
iOLlX,_5K<hEpqw,c	V'0D3&$;YF@yL4"A-!ItwjSU-}|Lso^??=ut{j:7ptI^/O6WXa~\xnr1vUK,2TaO-89?fwM_K_'lW93z%{XM?F	.^GV9_}9L[4+L>:u(A3S*&M`@1oO(UHl &?]sW1f_Sp.qaglM5S.8;j0{:h@i+"bWx%""SL\{Jv7iVv?GN:;*[|pt:BVo.9zwjCI;oHogQk7t=Dn"_oZn3k,c<y;.yf5-/P-(IzRp*|IDmS"\/?AQ/AF
<f]KZE%(	:,%*f@V]zc8j5Ii8d6NHNuiR@Bu9A_x]GT%U^xp,GiEnBm1GwEwwlMx\X+Z-qT%Z]I0wsZ\-JgeNPKawZKa};uC@:J`(Ls>Ty	dk-B!(0at4SZ/2afH)'1'InWJ>32HHe4GbY96!8ee7Jhhx,n;Yviy{;)cuQ,T#0H4vSBGOyj,elE'GlIHJny4,T/X/b{2)h;ClGV;73mgUunPU."Q{hG%GZNG$/AB4t;O\`kb`i5}-x:@y}dUnO9+m""W`xHJ+aX-P`cXW]XOuvHYU[Kl=Z@_ML"tbbWZFvCKwfqv+G@[By6&*X3|7%b<O\cag(nvyY.$;mqU4:R%n=DoBUQS_E)M-jF@0o:BHg48(uwFM7*BnA3pbXtE8}OPS&%02r#<&Mz\E}PiGJPJ>7>H>of8Jgoz$$Wx[1m,mYG+Do'pkxY+gmnUW^Z,);Izur8Zd&LmH~^_N^8f,B<Oz8>.'9g}}8-%+1dx>F%EroW-YY,<1uY,0t=zTX,\3B>GQ=Fa,yI?]hVk<:39	,b'f5;@V`]5tt]5u>Uj?-lx9W\vK38E1SW!JGCfOy)5knQVFAetB("8A*F1pK DGX[JrM<zg'j;IJ*+HjdP|Kv'T3]=AMEO6 =a[Rv)>%1ZWwz9Aksa&e[	y6Dl30&v	YY{\b0kl!cM0gR%qkVkm3w;(N%Q@}{Gi(~+ysi6&o}G&$re9L=T:C9xmX)$]:p>3*)<a\*bB\##\3"KkI?l[E0m0Tp>*Z\=>)!KSn{ n+f2G%$Iea2!#i	6Mp+6>4RUE?]hI>-+eip[X?JQ!t7"D>OF>gUzC((|KX<X;6*ZtfEw{Z;=ifM+N&.hlqqh&Erb.6C16A;<%P]iF\2FTM 
w&+N-}Ig}30_6%Qald	(z^/D c\.7z]>EUfwyXitH60}LzcpVFH9VU)xW?8<\;$Bg=R|'(v'i$&l<L-i&5P{Sk_j;db:6By8E_b?IP'u$ zyj9K8tj@=l)rq	x I\530CY<K]!sg!y{LdJ7u|8<2RvO$\>t#Z-rOg5RJg=[<jC6:/gSPbg#P/HyVZC#E1a",U'/9V5pVDAwM+TRlE*/*Wvl#!bo[g$kft}hyjNj- kxb:"fd	(UDe.tDXut }np7W	[fNwAL2RZx<g(nAMSZe`n?w$~wBG	A)/jfIT}eT[NH=3{9{2X%4@2QQ*s*onvgOM]]=qMFy*}ROpzstjcr$^WMHhLr[hQC
x73?\@|	uD	.$rLgH'(Fek>$Uka	H1v/aAddD520d+/a7fgY	b_edjJ_{vi%Gzeuuh"i-9W'	+|b\E6!&}a3	CIi/A*uAsIh|1nR6[OF18B(w6[x-e)cv"34QjRKtlK`Zm^4cg%=.eb5X--\"".!zZtR2(0-bG:4=W,o,x+c+_#Idm&!Bx8'N(g.jzC=LT3:Cxulw\kz391-XpWQ-uAFPt(+;xr;vqu&<P}b-+5LJy'hxqKBZU/
h~f$cO*I5N*@usBM;{V	|(jRHW<GI2*ZMQpN\2
V>9IJezQ%Bfs8WdBH`4aUF{]8l<]A,SW7FIU0Rl_+rzJ0veVW7y<6	+WVu'w=Mcc2(kpP/K+-!aos?r\:X*qKx8vPua<aN[6w`10lNrn!.aG@<QD8/48wi(*q6|{fw@J!o5PbIt|$\'v&Sb;`us';\ZkztN,z}Ube6vZJ\C^uI%Km 	L]9D3Rp#:>P-4-3lWo-X}/-@MM6=acnN`)es5`%P5b=Yp@`grCx2/U{#hRc0=B9Q8:z8! ";ta`4NK	1FP	3+{{F3)fGCKE-I*|$4tXE+6)}zPH{{a5dSv@AcVWC7Tac@d	pCdgYV|Mn}q>	N4IB'm*j>2q_h$u.RcZ-QR&PIa5<>&XkS59'wti7rFEr^i/f|]g0g0<Sj~oP8e4)GL,{Gq`VHsrnEg)O<0iRB/&./y=J;N:'Qs(V0sMl%fC74wM$VY$hg36e.P3&_SU6LcLtqE.$uwIg$FMz!1a?|:PPiGb ib=aP\&Ogi'qM<}jM<<K*'0%!1a{t(	
$FHg4G@Vuq6''"SH"C|z1?_^IkeKEh/`Ws)8%Vx:N4o6Tt`VKK.6ina/%oVH\Ioi"gH@Uib'a=ll/@Y>%n0m'tuG<7UG;kZSbosUV:P,>vJZRvzs[XVN*]`J6pF'Jt1|l{u4x*hUt?'&Z;D%7id%'gDGC0>eqr!#8Dk<!j%91a7@gMu	+p~2j7%En9Tr!< m)0jQf|v*ALN\X-&C[fy*D5ca|c	NSeyjWK?$a"	J),]\L!2]E5OE)$X*u$q:j,[:n3-KWO$r,~}{PwHB,hp%I&6MIjo(3fW
[$H7P'-{eB1qo{mac&':BR8B\`fSgn~|]il*U1"Zg0`Pp)\jz;%OnJQ7KGm?Scrm2?dH*Vl`q(
m{>vR;fT=@5p_TY	h=:,g5'v2xA'[S?SnH4b>2th&zv:hD-mwGr)xle$G`pc]8RUx@<T{k5M*P;kpcWs7+g^u0vS+rza(*$e-bi=y9Uo^(eNOtQQw)%j{o@,HBr~f|KH$><_{f(i2Es|=d<+cV?=X<reB1dXu0/Dh87/_[&R
+/5qmsU":H[z{z|K&%Z5qI&bj)A1B%E8Qz^5=~@U	.t0Fc%^h_b8
p5j&r<]o3--)1:'"cpI<u&pW3SIQ>vrQ-wInCD.[)luMR`7v%J.0,DXf^%Y?g*E\11N_LT3^L>eWrR^]//=I+vq8I@l'SXehBsF8f8i4rVN%Q\(g_%0OBK.x`Kba<R>3TH"rs0=5Ji]s&y5FKvh)I,NRq|x/lK50?L&"CH^$qe_T/H^iI_og"=1VZm}NFV l7h"~}[8^&kN sWv;!&:/%/;;_I*Ev_EnmSqkf=lXMej![fRrZpUXP-]}0wDC8_<`H<on-AuGaRaG2)J3yQI~sB<sm[j=UJu7do?=?S_qU?'ggsigZ,7<_RdMv?xVr3'/'sX2{6fEcIiEp`n$bw&YnnJre9vi,RmghvyRT3S6%+{M\>hj3HWht{9x>{6"xa`/YStHr:OE[:$39zpHL^S,R0)0["{]^SS@ D-8OiP%DBL#K*	a't+eU Cty&hmv0LxLaJ`~HWf$yIn\&hMPkVfH?lS?c*@)kHc(t02>foh`!>R4x>7lHAxiCbC!)ckp026LH'|i%w`go eBG"f;U?~6y"'\>luK|xXA\@9hSt0pkR>n|-I3.)KOD_"F'ymq#]e3Cx=J|QaW:}|n@X=wYkD76W`8Vp3	=|V#kXM@"5	ArQ[dZti|NR&QryI:gZXBMnj0V.*	\L&h %4(N7hUjO(E=2f4R*XK(+:NZi1X<r#PYWKI5Kvl}(3jU& k%:dZFK08.}>)x@v!e7ga/?
OQe,?QnHr'j=J#1cG*%YWN7Ka4-htrI'*2T6p
-"Ml?~L}J%ii?q{zRQ,+jx?}bq%Q>BvCGxU3wpdnLFW%np3#z6	rGUb/'gMR3jCI!/~ROT|(KS>9]2LD hS]rh;#2`'e 6Nd$0q*u6_cBx{%=K V,&7n|iB=AE;r2VoNu1jnc[3w@LJ2&BgL&L\vk^1l%S+n{5!_a>8%>v#!dRFQ%Wv@o40yJLq%O%KZ'7/-y8@2^I{J;u5ZEV\O,"U*x&!&KA.:_E?7Z;{aU`d=!iy`8;K)*DKTvDq?;>KlGVG49(j'}h!?ZL}i>S,!QV27#Ld8(5-c@_t5&m=^P*YkUMS<rLWD??9J1{P|	Oa(!C/	,.m?bl8`:&Sq]*aE7t)A]#P
sbB7irw*@HWnH?C+n\Ksbm'N&Ygc^iWL?x^4.Mwfw2	SKrw@@OT#|x+-/A/G%%]*7,iU
=wa-CljlMzvFi|.Z:tQq?S9
8 -VuP_S,m,)#T(-&KO	dr)/~7>O!WU'WU0`P4RB!\roI5F;Z4|709H,Z:|Q*o:1/E\I)d+gCZ7WQBSVs<BIp(|-NHVr%JGkw:W|'d3s6d#IK1W:h/g.ed"T`]nP.+GE6iIZIw*xk2stqPwww@2Bg7u>x4*|ScCmZ8?xR@'$H])2FYRc/dW(2IoQu!]nSs!DQ7&'!e0"WZIjJ,.XVG,>]%;C5JHO6-yrX/ lXB:Lih\m_SUP/Z+K1U00'?Kx4MYCBFKE7,kI0w=$6t3r#b-N.W~-J::?`$)m/~H+J)>y0G(6 PTtCQlQqz'XE}T*!7fLHp-WgT:$Qgzwj!O<t	|C-+Zd,sDfqfq:gU:acHjYt38>E1xVl6q];ZM) !$mG	i<mg#su`wl][hW3>*l]!~_Mj)!UHF^+D|!7u>SjA(ABLqUeIA8W xGty[HJt^w"!
5P]h  c0Mh@tTplBc}e|Fgj	Ta&YRAW.>4ne[XNw6WT.R,pmX";T<{>}5^(nhh;VW{tr4GZf|1r01O*MV!;Embx0N?mze]>.p[0-=&N-;}I-8=IrgP<\p5fMofL*QT`7@UD(|JT9IHD4`,/{Z0f|rREa!=(6Ow$ cp/G0h(Kn	YE95fg0"By`LY,[OG5:O3APK }0%MuH|S5?TV!crPL5EmKY:ldiT;O1ke3y[2?fp}O<*h^QN<)VY-,.>>'
&@$A#vZ;,fXCVN)g2BL fw`{w~ESI3UD\mTpP-_kJ{7}S)*Z^0p@SaGC+YqYnHTgQ
Vr]]VQg
p^;y93UQeO
Gp?C .RBu=5y(L(xB|k: BqB?y5xO;d/aYWn2_:1-GhD7{sMnOVW`Vo	xjX'P+#Ty6#NtBLUM3fQedDD9b3 dvLmyC}~mDgVLnZDS]$<C{wdK-@&J<xkRA$z	-l;d%m~vJ0+{n_~^A b<L[/g`1}z7UQ3edy3w/]zM`/,Wd*I\+(r,AeVZxxMG~BgEWN	n>QfI5MF]vL

%0?C);3~I+O )Hb*;vwh</IQ[z 2n%koVfhKhpu]2y7bkK0P
9`AN<b5zq}O!/^pWwlI.q)f~<?4bW<H1aK=6\+*LV0LKo6%Z6O:bB6<BRp9{"WEPP>YUl(F[kIjiAOeqD>JZRDj+]l\f]vW"*q34c>U	dEg(BYYac/Gn=q/+8K\~- R[s<W.>{G9y>f=6Jd:,N<-;irWd^z{Q#jZI9G+(lr ~m{Ug0 323x4i8 O&ivni}8O/~WY~<8$R>~4l9[rCB[biadh"E8t=)wK:}u
Y_oTit0qvQCA0U>YO3rSFM9As	r*IjJi(ZSdCO9}QhquH$7bH:l%;@ nj}AbQT[?^0IL|1<ZNNXqr(i]/u{<LhIIntgmV&C%OA:%Z<tXS.6DlX~`,$e
.IV}
j#[3v7m+4
rP2&v"\zqV/`!LG3Up~
YnOxFp6{tGoH%@"-}|xn^|D/VW0ULND_z2z1lWiy:AB)i8Rw7=_HLTp<Kh0!&@`1sj!4j>~!)9(eGw)7CD)M;`@"t__t5c`@+%3`P(G$u1b![BB0)X_>d=mx{FZu[  @*^1]Xi
z20BrN[a3:Ov#39Ol1UlJ(xh_pR(ksTO/&,24p	*pq`eiPj6{;_LsFw9@QC9HR{q;="5f;	XwB9vaENT`E8sv.#-4p~mAOC3 j y	K]"SDZ)Hs\I5ThN	}4`9J&C<2"MD[[Nxt3rFA`6^>)X;N
9!>#4{2'SsCg\b=`7TE<14;I2j%xf7ZI,$PO2%_	wDEM]IF\9)Oc{P|`E9f82W5`,bFSb5?HPzd`"R_7	I]tOaO8q>-4TK5M,T(*pw"Fb
S8+5k>H_7HsCr(b<g!_:lcH<ROWBR/.;)^c_=6Z-azB}2*,J	!v2\'c!Rm!n,0ZB&UkOJFafh.#S}7"]#>$y|x
j6x="SIh?&wB}$f4~b>8WX)kfQ`FixU}`%(Z8zvtbl&PD!h>HXic+9>3nJ+;Hxme>aX	QiL3Al?zT`e/T#Q8	FwF&%9gp0+(%{Q\ou/VTW~GXy\!uJ8bzH\
~-tUka}%Unmr0PQfvQ}oQw?!agj#Gf;"vMlbhgC8b0y KnHmPU+)5|y'jJ=#fl]i.*MoPX|1_n	~q0d9hNHsD"bR:	cp;a:hiaI)q>wPGhk1F-q$5nlTZ]_R0h>	/N4[}TC%Y. R'8`M"XdOiF)a2?sr(^HqrhBFf$w0kAh$Jk}@[nSy*Mx 	sjJ;;{w
{-6kI6\xgBq(O1):]Td*lHQ _MUQwxCU3fx"R2$c!s(+!x}MDCB"]~bTQ+]6sUqS639%pU[\'-ca>OpA7U,Aag>wfN?-,~E{wKch]czMfca&'oC:j?q3\+=TkD*+:W
m@ibunNk&GR\\dgQ_z<"Av?@SX}
c,g~uUb>4D	#m:f~|+
^r9&A2LXmC-sN28y>x^J9>vX66s&j>c!"HScoKQ9]?=d@YVZ1C <P
h#Vj'l`t4PLJdq04Lo-slga|spnAY
iL3-Bd]BC@CBY[0!4=d!\AwMw	e&%nMP|,-[2L<$-t](6jqk5p^inr2I.^@</G/15Z9szx;O=tv^$=w]];]GX`h/n:ke%@/u?){|UYIm3b}&,c.EK,!8beD;gRwzP#JNZb<_V=h5Tg4h0z>Csb<2m#:dkiTKw.Bqq)fWf=u6~En>Z2=z|d057&)0?q	:Cmi
S[XvMe\pxSs&+Eo4El?Ju]+!KVq2qyh=wWko7?l@"c"X&nU!n[9U6HbXd`4Khq9~'4i6JCV;+tTd~qM%T.Q$sEYX7K\uWZ>nZn10B4[~g>9IHjn$;WVC57
]vUZVGD0T_KzXc@D0`DSb__yi?t7cex7$DM0FQ1CH3'T(hrvu3an:FTlm_mhV"4'5,BM*;WM)iG1B'WgC1vIT|@"TlEq;D!3K
%sH
W>IzBTc>PTEk%rrpD'
Jqi&* %zwPIfF(ymfybTZgn7}_(axmSQOjN;O1;=^Z.Rwp{Qq.WD'[
+>31{q5Jv!p`NNJr{>ig"{~c0+*/iU&>\"z=W$M"/l$G:j8^zfO73-@N.IL2mO9QbA9KL\"+n$Ey9	?!#OeGm*2^>K@ amdqUjMGZSX+2ERGaj|!n`/&Y{bb;"DC`IqmC@m`Z~\\9J.;-vorvT"1Ql8N(5Tf2O4
<*X5\GV=_cu_fzQ+j zk9#T!bN8c	H[8bEoTY{h{jpIbMo\BKnUCy8~ev ",kc:QjdJxMqdX[1KhB("@h@xg E%|>7"*I73H&!L~RL_tP-<\)yOU	H[,A'SS+vActhzn&u@7li:U1f8<p&bf,'\W@x0B8v52m;\69`xu/Wb,o?C<Eu?kFV	\ici;'#uIK"'O+~/LIQAYTkP_l5_]~7wOg*cQ4T(
7pkV+R2?N;5?"D6"s1b1,VB$_y!df\ARJvA@:ZTY;!g_m&T}K(P=<B?CK=8rbc^G4>0N/*lf+9Diu@>R6G	+KUNMkG	
q;s'uzWSl]t6.uR:""<u6J|3F+5DbFOcF;)D%%~U&rx!H J~Mv:P\Q +*
xD'US8R+UFJqJ{17~!2
yQ<Zz~

pst<.iQY}_^[sQwf{b66HX,x]2C7P\Fn4N6	F0NuJngn*OQ=};y9x>YbcxNR7D28#$dv/+f	w)3+3KCkW6y0mu^I2ayKB%x=|t!r#J)&
vVb&}h?H1}JM1sgy<k`Dr9_)z>7hHEs_#+l\3+Uk^dVx7"jvRt:Z$/^4G{=a>{8j3$)[a9b/SeWgwG3R2)de QJQC%Fx`NJ)$5_jl^ f
W	 sxuXJ"-`t18`k\V>^VkYM+rt=>wd<L,fpV8p*53q:87Rdq^Mtj[#N\yR_S`0[/01%mdaY5"E~3YIP!\)4 dUqkk(^3tnG,s.~9Z"g pq_e|^?k>;NTMSLCInOzue^OK,Ym3YN{D^Yzl4_2]j/vO,u2`v/X+](2[-,-$[q7$>}gNJA7Yh4/H_``V0*84vte:@YbPUAGVw Z8,_C)#ijOpjg|n${wjoX0LT&Uwd]E6a!EfiOI@ue96gmE}[g6\a_QpF"W"BI`g#e2Ov0xjw>@Un;tAYnnEK`fByw??s.w4
NOmvnuK3ZOR?<YdFK1`D&PNF|0\lH;$/UY<FBW&z#.9n>/0]8+Wee>2@z
g}Rb&\>jGqm']JFws88#E&QijM<IB^\,t~Z2H;#1iH;MlWx{&Ry<vA]-.h+fMC\'m\rV,r$JU]T44t	i>tWU nwJ8<W/-GEH0$K')Op`Dw|Fn4vF_xs[:9~{vS.h1n,Hv;sx>nw7P!X+5*y5eH*ubcmTHjeWn+jZ4$>qHg\':CBaj$\hm	)i%|4x)zSF-Le'#>)A?X_/Khxy%zSOPE>FmFXOkk[w(c/RO'@`J%\TPJ,;kaC\7Nf=[V*A */=0,\)1l@/*=/|'#3DidfQv3m"&:lg8%)Z#X!kSOc\W<7~9zb?Wm($:Fk@7aWmSu=/` mcN&avn\BTYT)P1r8~]4j?8"y+,7e;I@ICeafXQ/M`hnK6CN>rPy
D0f2IhZ1]`f;"#2L<p6`5L<!x 4K! 7Cp5V@X@6j.3,4D^4sr{Hc(}QR:;:u[Qtqd/dVUD_z;**9CB96-L;0Eu5	2v:3VSh[Y](:"KK@{&d=.*NK}\7O@|,*(o VJNLr~65!3~0E"A=uXbMP/uGmXHRqgm2M ZyytS@3Y0-{qj,p!278$)3u5)JU%_oyjC/0ffmG G39aUxteo"Dr <}5{^gcn.IpwdC4lCQ?i/o	7_1/G"OE;(}dNA=4PqX!;?n*FZV@)W;K#;M#Tv"c6<$$-9^lmJQqO 'F	ln{,,}=3|U[5e%W^ec`:mX_^5G{.KZW/60Z]>
<CJC,#X?ZNwBHM'm3ZZBO%++<{Nia~;cMSiF&QF$[,d0&OMr3.j[k^O'	)z%@Sy+l~=Et**1AyaM92KYSlJ;<B&HUUW?^df0$mbHCo[|Ph(NlO ED|DOdBfmp%;yi.?3AB5\bI-JJB1F_WC$]:P
?Ungy%,,YQ]AeKlZEp1aR4#gM_Ba\@OXaK3O:UpP#m?pgY1;8_:uyiN;,1|\"g%]]e&r	i_y^R'3xZi`K'E_31JFZ:EN7rH?"%]MLWcP~4
#p'x73Ros>\E.pb!e'F-UJKwUU1B==R>pBRvAi_yq_W?uk[ `u%,DcMRfus0Gl&wI|1jp	dxc,]#[eZ}
MU3;U@>+##V[)PR&`3k.vD?0|&)qW	RZ{{*JV875TIp82[QyE"(?#aFY(R/U;cpu9,S1\/C.S' 
UTe?7-RrC1_y&|0%?t#pHO7xgycURJ1e3o5@	"'GNb7UHI>m7Q(3#
\Pspi=s{,B56oDKD(:z
WD)!I%mdAJZIM")-[K=wAEUX[Khb~l/9uPc.Gdmpx`OISp$c:yl.gR?v%2x"MZMe9q<)]FCOS/n]CgR54-3S9nZ*&AW)f$XPa>S%0dFcbwpfE!\{U^q7j8DwmQR=Fg87VDx<
 e]u/(!|F;l42(Jcb6/Dwx5*=c?E&~WA4%avKsI32E)s_AmFcW'mhz9~EG7c'l?CD1Y)V'q=0nP{rr`9=]} RC`qr4]R0LO0kFY9DvpR2D%iA]ib[r.uDRg2;>n.?XWUSn*mM2lTOSIyA$ag?xg8?q@|0Jn<?|XFVrkH oW)_k)JGOq1g=_YrV(KknQ)-	}tz ^OQ+]*;8Th(X0B5%"mj7 NoSH:L,b`?5:IUS?}*e+WlD$=KwjWR]W`Yy]T
cD]}(~^4p*$nxET])Xn/HjJce[	wvm}(4O?Q,:fn3yAog2IEvIfvK'"l"57QwsQ9n3:oFs%W[adh
f@$OeAG|XZZ	N+D<F|}tzT$;czH}-KjE	/+Ne<Yo9FxicfcMJ?ko"z$=1YOOy>k)RIB\WBsvti?>=ik0C%JTz:#z57mlp2Jmr}P*[X/Sv%cS,lsso(-q
[Qm4Mk\8r:=+6+Qwqf7l:"4DD)]wSgTCqrW>pNZ!sVB+q-7C?}]J=`tUu(,p,}<H= ,D)Y/X;@{B~fYp^(=Xe8?iMaE0!SNCkkvsQ~`43xF`B
7K^U|R{YK5'LJJ8~E]z8yJbWOzJ"*xZQ?Pvl:L%b;FD6exlpBMhkjO2i	m.u3$TrmmXLGPk[PfYqM9Q~'++dJe97O$M?P<5{tq$oLTE+EMgFh?GjT
|VYRv5T-REvHQoN8nXIZbiv#&mOQtu6{1G,4zH$tShy>!	M3S@@j@]>$%^iT:"k:3_t` PA&E&nv2/K?5Rd1k#/|c6{T`aP^9So69Fn!r~=txk5i.'Eb 0{o
p2?^`&U[IOS8j*"CTZ77g|[EWEi8MDXN|_%?JEJTp\7TfSeCl+$ghQe>|B2qGi_V%zP/pp>3B
M;x7zIwO0roYa{/du;[F/=_FF~vOQ}+4Q"xP)<c.{:UssL_|Fd\_y	Jt:<~)W;P1(#J(G;]FFf:8@Ue.rr2BQr"DQA|Gyx<C6bv"~`N{${82mLf-')5>b_FgT!":Mk?)/502+gB<%>Y$8[EyG%ppW[O}h[NecCd"&@orkGF=/fOMHD,7$k@"^Y#elISQ7evyJp
fE91[mxn6k>8&.OWfw6_f!vk=T
TZ&F\O<V~Z,+(@`}>UWZMMA uN:fk*M~M5-mJ*S%.a0.I,l7.MXo5wVk]q:u1B
^zF{gkTVs|5_mXHjp*c:iZN]dHMvq&:?>c$+Ml=mp*E1E_Zh+'}f_B~{SN\8MzTlTz	]cV*pyrv036UUTWb^g2_kBxL:zo%/(V*BF 8!XX)2f[.^!)w)hRq_r(K#)'=z1B+M
6S:h6u".Pf:T9n)L<9TLc?.	CRl7n 6:-z1u+cf=2w/5+IzXK,sy#Wl+a(^(*{V$Y!V:h%Y{b/z@Q25.2WuUF(r-.xT/Kf7Y'RC'U]CV-zuok7!daF"Ens!vf{*'nGFGTo.@Aph/r|lW(to3&P"-2Xy<(&/vUN_TVi4F/T99V6v<x:S~#za%$m_xt	H`//}Rj:gI]ae<cPj&p	wX"0Kq?DBLx1ID?S{qHO54[{b8UA@Bbgg_U*ve>XOVY#:;QmOfCER5(+D`>B&y&?)Q0hRw/Ko_.8`o(/;6nlOJQy%qeq*&nG%9_nWxL{x*r2xQTP8C`~h\]n>cqz.~Lh6f	N\1xfJtna%xR)r`Z+]/7x,jCHap	(&%m1y4?y-~q
A \n-!M@ #<X1Ebd)_0z0'QW8ACEtf7=s?+oUn/&/hZ\*@5@(000\xZ\9-rZ\;u? 8Y6wz5;f)e8b49kLuFB%CkM$/q|+FZ7,`i{\;CZ3C%GsTtd_XXu< )Hw-
1Elb`ikSK.DJLJ)\JtOB4&)2Y_;ij{fJ	bY},kvkd-;?=	V04h^`(C)Z_[gKqo*j<$7!T{,flPDx.C
aATj{l&TeBY#>/:>MtrV}RQY` 1?B2k(u$sId4,Yk>[wsPn7ZsUMf6MsvFJNi@y5NwTiW2:I>u^$3mt.Hv{C'}5rK[_0D`*=ykF	*/=B#Q)uM weDRC>j<?v`#}36W?6BUW2mei'}9x@E4
aDVHUcBtoc2wCk&d\b(BYbJSb":xP6Y=!>Onz'`EE-<T[ 4a>e(0.6SV"|0BO^y(M7JwHDui$"R'Ym9F{\9wyA9)@@h(uCGDCgK/wOstd	eJmYQC[DO..\t_mTT9dlz&B?%SGUTn_iLK$}c(:6 egox3&2XL9VpVD2+T'F5~T%qgB"zl-Zi_-OK,,uyXRNHq9_uVmXu}Q$4Qy_h@E}IgsziYR4MUOyHQ<qX9yn4<|jM/`(tu-@ZZS}IJQ67n^Z`\AGra2jo$E"$E&|`%}en9tRp4b~`5DB{X{ek!&\5C+VeA7Z*XkU/HA-uGg.Nygn~*)nBb,TBc7p7SPwkUgBW@Wq$<)Ns/k'3/G$R'O|<;_]w^(;E?V-I0amVvVT=:[KMEcC<C:K3-p:|(|e.&+y3,9]gVRXLs<r^uS:/<q>Q:	8/BmHcn6u%eq%oW
><-_nQ$`b)<U?	E_[\cy5$xmo*VRGdaQd%1!hj!6%ZZjWFZ\ ^I`2`2&dL6~*Qf,Hy0(dYPh7xiF]+Q{o|;lTO8*o<7,qUM-bGCL}Rk+\1L6R_K(9UD-Zal+lXSfMP(/Iz=,6a=$m4gV+saq]D#A"C%1w1N:Lcvov4,-%Up+	S_!D	$V