'7q04w^:|'rS{t/Y9Bi0|{p-0S6H*aH'jkXuN.
G,P]U3vbxXU7UQY_TpXRCx$h^GJ0w={JnaFX?0x3%{.\261uz1WXK?q\i;%U:C{wjHP{ay]8S*Be#n>7SV4aH<c5N.t$</-q3HzifrRIC9N[*]Z.(5%hklwA@:gE~Rwl;6[c@nrIQXc5M2XB@9#p\cT`7L6OR{D+jN{KK5/B8!W{;&+(N7Tn0MM
KPnhMIs+~``F1N#4m WUf_=)bg?j4P>tvC_*vgLE>cF@"DQ
N!q"f'ycGG`	?u7O-W^*X/vMvI~=7A"<o%T2EeCx.fDC*VT>p2b=Mi|oe.,k%SH:LkwW(e$it]&1;EI244>t@3[YxHv=tPtTrz;iE~2C#*9>j
N
9/?[pL
2%HrD8]HhBZ.cjYp%RT(6|H,OhR}K;bHMz&(z^gZ]d(5$/z?"+&`=jEv ;N9!nxaMj81/wU 4?a'ZmAN.ha|(GuNaVAiUq+:Du!HL
S|Tu$h2fE*c*?q;
"p	=Jhd\3!7G@uy}c'I[s7KVSR~FmONQ^2h-t9t Y{Uiw52JRp+\rwnO(l%;dv'v5H5=j0jTc~L>D\-#9efll|uQO[K,-TBTu
e
H2N;{RX+FZR15~i|MW?-$J]Yfs'5%2Op.e ;TQy6}5/ME?n6,BKw"^}=Y)!Q<5'QjtguXLacn|,75k
|$UZ.~f[/|p1u=q:w;S2"{lMgJ.go>w@)#11qUYyBqpr~e)]Pi :u2#AL1IJgH+	jaf0fe!hjEAhHWy-UH7CVaDX?9_|;Cd$GyWmgFt<X;lOoy`\BPSKTTGFrg+{h&Dp:}S'E

h?D`8qQSZHQ"X<Y`F=ejgyWRs
{\\P0PyTTC#&d:0=KH"i}!@^t(~C{sn7q`^KcwKM6k/%"g602JjZ-`M1u$Gp_JLsrX_*&moWV;[k<C+o!\Qo8}[T9'=WW/]/SrK*]-/sM/L/~m8e
n0"z.D7Q}W<tQ<(fS5uj5t%b1/.|BS%3Q"~
4!LI*}qxGl]E=tPH,9V7!9,BJAZx3,3,XHX/wyY\L^(P6o3'NaeUAi_P$VDJ`Ad*lwus!I7vC* h.mC
<
mBf&CJFN7zVne]J#x"Dy]-ydAX"wLuvC#51NTlB)?SHtm0[@S~lfD2Bdaea.Q -cAYfq8Sv>6<m'k1m_DV^Jw	O6eZ p<CcXBW8L+~VrET$TF9ua<Uk,[2J^=)#:Iqe:p5<[{LR=+P}*-pQp+:vI>gcMNwumPsXM|HRDHY8f{#6OwU$/E1WSTv&7w-M"n\70H3,nkPSB^9dmQKX8~\8f+2K}9S2EDOZbfBvCVd?@Fq~3%`4^_He:@*gvN91QhmvrJ#IR
x})SmuW'H5
>U^O m5$OyG3"#5`"hhYwSizc#HYz^!,7MdLYBJ`1h$9tIQ2<fs0!b<!/:O7Dj?w}t/Q	6Q@_&~UE4wWKc>Ue`'4&T	Db(N)Sz26D?mwL}EsG0UhgC1` TgR
A?Je) ,dUm;$ZcDH-X$IPv:@wpZw`GF=4_l1(hd<.<1ij/y:(u"_eP59WnH,:xbz	9Y!F(_e-#cn.[4tREg86/ws`-[G<+)WWOXA*'i,ZY3"%( e.gsM9:L)VN/HhmZP(
)]-}:]qy}v:^(,?wg+<dh?w2\}3)+&ROP]}|LNZ\4R9L?i}[f"5y~@zBmgReBC]%RVS m;HMNt;0Ew}T+g-M;YNHGYCc+-e(zPh"W`$6lX)^6.E?j*yZ)	.e2L+]+G)TLCT@M,Y&fg$KJ|`bvf`2bivLna<"pY"U(,LV_T4mU>go\oux?HzUFNPsQWmrn>(y*	x[jO$xRYI~]dzoA?F!(m7p	L<)"Rvy211u2>J}5wi8xs+mh2Zh&PHHn-WDvqFMZg;xZ:8XRDU)/Am'Gj#Caa3YEepA&3%0v9H-)4F%lE'eC5lvar$'L$8$sw]z4|*|Q44Y:}fc(<H	k$\4fWsocF2<'<ke-\Z51<`ykU9c(&7rw}9P{j*j]/+rw/<R-qzYs]=wOH!`!dQK|S_[Z7H$TXA#3A>5/C6[:7A7lsi?q+Zb*bO}?^[JYbzv,YEItKF;ZaF6f.UT*i|}Qu>J#? >;9.e	iMH
rA^o=oM70UPQAtT[7&eJ)TB8A>? cffW[q}:1M [600={yZE^"}WV*\\Bb4F)DOWtM3Qthp+6Gx"fd>P#=RJ3Z}H _B\*xCk%,QQeHU'>S[3}DXYEa%* prW'?@mldJ[ ?q{f_x?L[6VE;<drgW0-ay~lO
BY>&'M	UHgk3|Y{wH&hBX
s%((nM\9do@,|EQf[PZ%nhPTSN\GGeeyAcnV6~~[RSEdBg\abOu{`Rqq0G{+.7V4':wn	,Wgg9-KOUi4h\Q[lR{VN	Cd+ZF1u3i
eejxDeRxg>}&Nek2pM$8CFks^yttk`+"Bn':lVoX8C"~Wpg(_lXv4:	[[u?fK>\.8M^>O,G:Ot2h{m41N]"a/LJnQg(T9^6/ZNv\7]/V5Uw(FN]8|c9C)C}NX7,]%,vC-@r"F8YjBB`OHBNoaPgv
N_?yzp=GBWrf2ltlvZ{b#6b9.ohwq*]zBpy(Z2//BbokI0cjEPq[HFh'fbLDmGuBh`{L%\jhnB\iL3_5dzl;~k|
,YH1eL3P8]Us3M`	yHSGqA7FAzPS]s|VA4PI(o)U0Z7?jS*ri3]n?	"jR!FT0;5E,n2}0l;HyBX9"'O	_R^=6A+-`T4FZwOh6kUMn\	qu/6nC=B$ua/qdEZa%<Os"ccKSCiZ{xhj,f~vmkiPP'r/
Wb_!xM": !rfY%ja};ASyBk)FW1ng,>:
T&jw\<$7wt:h67dq"K', Q85^D+~7L=v.Em>|Lp}C  q~Lv1#EhS+G3lnpg7[@@ZH|9O/<t	i 1PO)bB]ppMwjKObbi;#""NH.	R5+5wY7>^::.&|1zMJauhF~wbS#&K7Ph-r1Yh8+fr&?xp4Ob)5h"{O<WPZo(5L)l@sxZT4uO-bT>;0F5f.A"kmTO[IJ^hD?.YAAH8&iHj"^aGbZIlVCu`SMLQG`=jO-B=a!-bpg|Cp\X|Ae(mft_K<b.GJ-wC/oNto}:%~"GaeM$K #j[;K52mUBR13>]}~\jEkrIV!%j%I)8T0Kr2'EGn ~71-_`3gTq6#UTgx6#58$b@o^QNE~3tsG&c]
9 2\7;eWao|{+y
rh(RID5)dU9U)DLQ[BmH%\p$%u7UV"MUp$:l)c}kw9D3;Fo!l]t=Z!MhU@TorNlRkj}-@,cOM'*ECGJw=We(l'mL3gaekJA'VS+H_YZyC:.zS%`k<:B:%b!]AsL.D07=6R4.]iR_i Tq>5c39hcilN*c0yu`I+<j=tQJ;k]@<4\{pk" V%r^I6h,|&4R0LSPcjG-6-
/t:8%TVyvG!_4Qo7		sm^khR.6ulB&}^;dGk1C P/CFwoz$,5Ng#Qp]F7tP.L3u4!ns4Y_Hmdh6D('<*8(_>x_q)LrGd+.})	C"3#:2/RF4OB2@U\C-D1U>wzTb m}pSzM:3{qTQ\|y:}#wIJ^k#kdL=XztHpdd/fO@STN?ke.x*a~]TQR=8bg6{Fnp7*G}$K;%E=2
Oo[s(B\S k2uh\TW7(Qo.!B'F|bRwYjQY7y(:($Oj*yn2"gU}HQnBtQyHW4Hn&lnfVq<}~Y<eqN uE(OUw#:2!@;+i+YxK:\qU#gP2HW{	T'@v1g;_r4ElQGKc?ImUOWtB_Ffz<QVA,gxxOsPXu%ykmBb+_CTVH\a.Li!*S}pxiVK<#46wQ=_7L8zlN#0yK1R$wr=]fq?&H]k(!\T@k% k$925wk/M&R%gh^^AL`"1G#n%+'Nx89XHxS65"<%XLw/aGs%,y)-b058>5KOM^W+\"eV.DgvT&rfH2S2m(h,2NA.b
^LM1MaV0l~S,7MI=zCwV;WU86IV`sVCZfU1JEa15I3z
LwT@7QpGV)]O8ic-@t'"1^HjFu[]\CI 3m=|{21x"t@}ZOCBV)~Cw}iW'&79_Tw5E/OJR2xbTl,:9:CUT\TlRo2_5Mu9I5?4-=KbmFzMK{<4;m"	&nbbj0dNa!y(?`C80V>8Vl@dib'%ME?O-qU@V,5JXU+_~cG )e"!\t,*4v'2$5i/::oW_FcwD*]/bC2]Abo^&/^F>A0i&t]+Ri M
(^TV,g7Of
/CucD'K^0%a6s, #J*\&Uem nAytdk!(|qq5/B+"bL}nP5vMjU]hRw7h{S4DjN2'Ju62;Eit2]8ULEV6nffJOluwqzx1rOt|$5^Vhfe[|DstjhAcy)Na+d]4G;%/+z,&g"5k`PohE*hus@c8?s,Vq&>G~+o>;|q%(QL?]v)AD_gHM,tfPr6Geh8)'xmXQmV	gvn'I8TK!=$gJ_!)F3}Ga*vR>nJaoqMn1Gyk]0h(Yjw])cn6wrWB_&7{Mi;(3sF__]dKI\R\2COK6sY	LJv?O	uT"|#o3X5~JRQE/G\%T`_!S)U-TCq1I|`ND49}8#Hx_8m8;7hvF|\!:lv;a9='3~9AK8MlC>^{[LES(0vlw.N0L47.{:l@v!j~{UzRigW,2T@l(lI	Y/ksLn(C`|p8%f C'YmD!G6' #R13oO*e8ihjigW|r32^x_GNH7D"b$^6F}	xXTH~*C!N'u3/	/	o .~#54I>_`*+u=,6fpvK4_H#Idb;m%'{GFyn9/!LaR`
9r\=tgOZWw1,&5"_/?)Qz2A'm9SiXnw<ng)}xpp~Ti)UtA}E/7J,mV!yf@n"5-PC+67!%>v-18=|.]~XySnBN8{r!h|1lL+Uks_|ojBmGm:6om6Q1&Ah:IZ%.p]*5f|o*oXHjejK5DEm}AX;ew}#vo X:f;$^UHCzM P(eT6DtsQr?uW<G5#9V58"?G(lGVH2$z!NI(Hg.t5DekM_1PW57c_r)2go:yR"G^sz(86JcK
nOB0h\$EpiE@Rl4SIO"0$0_\Q{]*N*r'7N34D<_jWo-CU]7_1T0 v38@@;j	m(;trUp]{e;
2J;:+/e8RBu`:`Y}O{qe@W.3Sv-C TJ^KL$P?/e+p^QeE~w;\2U;N&/j9F 5^<y0k>M&]FW5tY-Ps.#\p4&3J4_|9cLEkz|!#w	5:J0$~'m(BE^4oQ]6O6UFW36R#/l6{QP)pu`M_dN"jc0`2~s!H^50q6[h05
3]$fxrpp-i9dU02W}kXxW13
Lz6H4$5m`
mZb):}d4>*Q$u4kA)P(gKXbCT<#=e0lxfKkH0PJ6V%5=w6|L| R&0`Ih+5_C%1\
Ho)P!_h[kFF4jFchgfH	uVgQ.n[uv=z#d
nj"aa	JO4xh$$kyvgDw;G{C3]?}eU	\yRwbCX~ddSA11YD8e2>J>"f1JJN<#E"ahDbezZZ_K-B_`YynKIO.jH0*r*3qB?-/F:>,om\0|Xg=)\cPJ W^FH$6>*$Z3o9Dp,C
Z*g#, @I#q$0"Ure&I6Aq5nP4)et N=P$i I35?gj`6pqJ`i&Lg:?Bmr4x~PMme;MDNb]5<4VsJ9%di9j@N5=`Q6$yC+'`x'y%7H^+h?`5GV_dd4<og3<zgtNil$>36"ZVYb?y2o;JCuF%Qam;.*R(dqZqOabY*KE0<cO>5{]dzt3m,LL]fHvtQau3=1fyoh$S\K}9[_cRh=sh$oDTo;us_!`v77"7 *`j<#?1O_s"wMaC)N}qb(dGp<?:i%YBjWc69IB?;NoBbH~]ROX;$.`.uQV@rFUFK!W_9	[NsH!m($&I{!9Czt&zFKw,FbuK	<+|+9FL# A
aBt!fsTR!Z1,4W/EuPfh:~pT\nk/L.6CfLUaZR01.e^}i8S%rv\F$R+LHnbn<vQVp0VG^w$$aK'V*xYE['0V9z91t'f:Kw6,^)'bN8HHaEly`%H2+;7lSTkiQkVL{mD6hrEV0L=E8V\QeCsTpPV<iwM/A#Ndb/%r6nNNv843d+p|Rbl"Mn/T$b`0bOC'D_N3C"_Zw2!7:$2vy9eA`2	SYPr<zs`u2NM&RWbhmLT|2K? _?LXDU7"lbv\{g&UhiY!D<TCH:\2l$|R{H$l _dC4Za9-g[_D-{W^HU+__[PrN@KIvkqNE52e4{XH&&D<8avkg$jImyf(n?~WQ=OMNZ/Zy%Uj.mR!ej:@d(UX+*a4&,}aixKpBG,dYaU$,rwEnNWZ'y/B,	XG_"<e7=M54Hp211=kMqUsBPo}I(5Th/6TF4$MAu#Tr,HdSO>C,,sJJ*'c~z1q)1?EiZVA?Q?g8eqOsrU;}69f	O	~-glh3'Gc,{5<.YeFv[Mga/Tn.P0>.Yv~LJfY{zF%@m5V]
wqp(j-yO4Y`1^`wRJIw$!_y[z]D;[Dvu4$lzs^{D''<0?,XUh,yeT_mn)`D}"c=etKq$b/vuxrl9P/Bd(b&UCMyTh`H2ME0:Zo/dEm\#og07`,.?<8{V-7$wYcg(uWU|a];n{%O,=hNc]1,#Frak!C&c,[xB%[N7,b'xF7@O.nT=yQHh"[n%ejl2}u&<XO9^7:IJR%EKr;k"rtk=23P	j8%z='5Fb92M\?iY4Cvwd vCBJ({KVm5Kd(<BF%h	SRyQ7s!3q$_1HNb],_sXIX|K8Bs0T%8f@"DZ0pG8Y0Y('>r\.3co]?<C.&sbi
nJe.c<P/y3D+YBZgqC[MaMg_"AY!s)QXif&Y	q-`r\w4^&LE6IO/@'	B4ItnV5!KKaP@`zO{6&2~f7ghr./K'A*W"9zS"Rf0D?:y^Po
F%I-W\4]0 p'K^2>dc[~otDI9[`
Pi,<{ID-(:@^!
Y`X:I#fi
]$n/lsl044!v/I[!^x)0>re`['w\t^`gT)(93|F;ijw(T&\{TQ^uR}+ni0)gW{.~ixN(EH$PE>u^JtYFL_#"?B&4*d&3ZF7]T@o1Qf>mVultZ=.+Y77>MT~
}$uFToHXJ-zPJ
.`P+Smq(b."82mK/A(.v+=0%]s^)n|"P]^?>H0B]gMy`!wq=.z_)u[/y6P@:&\u0'>\Q'@50]xH&"3(2,P3>bY
:Q4hD,tf;v|,wd<?L3#fK9d*E6	,bi#5%C@HwD+Jt=g,V<pI3(q7P<ROPVnhkwQ$IWHZIX[U?;gM&qBxcvC{OWv$EA4ht:q0v>QI:nTaN,!u-@zsEQ#pLQ<A5
S'[z;h=5B%U),A5FvzDu#fc
YGr_=&&GC^C~Fe9'Jd-(K#:7QQnqmoN<b,1"[nGfG02-B,7Xz$$Mx>)n%UP^sIcHXRchYgS4n=_mv(/mq fQEN2QU4[w*MF[f{Y120]@k,cp[x
y]rSmeJ/)BmnrF3~C):pX
^aD3'Tpx8wJJiX4*DHQ]vCD^i8M/*<dZNkBw$gzS-lkpPfa#[\SXF9?Y0tF&sh;_,z9BDj[j-`y/-O=1_/.xa2&I,{Ku9{ V~vSR8,hub8/:TPED8hguV#
#nDk"FV{W}$8ncy<j8_udrPuaf+a7ao?4#u$@.J*qP'W3\`py+PgQv+(`cI:*ElvrVYcJ+rjm|z*<Bhl(.i|XN9LQL{y_Qt_3<"	l!k#Z~lk+=0`MYA{':V<-WqoHgE'
_2K25>uZ>~umjF*x/_!iC]Fw2@l!QLKe={F66;o?,JAJ-G2v,_u'Nb/wfDf%9a:8@ZESQF5
5$|!Q?hiQ#:e+a@jEW8.qu\n	vZy9 IcZ56fcK$VTAVuXV:0l'3=RiH>A%w"($"!;eC6dA_+.9QpJn8wVcte{O|^b"@M@on3I%1Arm^S+dezV)kJTAxHQ?`2=
0SLGEPWl+N%vR	3kh_AA:]w3T{+*'n*xK_E@YJK6oE=}ZAxq%K96ZY;FBT?C\i|09ESn2:t(u$X'GE0%wz{H={|P8%`sZ|`MtH>x'U*!b	@6z;ran&Wh6x,u nzVdsRcT^z4xqE}R+3~-3q1%9eW1CA&".T0(+Ei9Cd-B|gU	,n;.0r=hlC@7eLQ,-:|
th-V> |)^\LF=Fdm5lTF.B0	ZW+T4k03m#>5cQ" TD9a6l'hqRq@vn!-iKyabLa86LBtO8n1o(-b gtklHjgxxHSKJ%_sM@c&dC8Z{1!d8\0N8ktOq|BdCb-<$;Qs:
7W> 7L.>t{miI8SPKUCgTBGO2!2"XCn2[rL4W9	|i%zK<PQ*B=o'),jh-_}+oHpp_$5i}3PHHHF=}Mus&vwIxh+@12_E;T
4W]LgQN[^.VZP"i;XQ`KB,afGCVA!c|-R\]>)i4i97YG^#T=R4cWb!9B.h3fVf\8lR[p<[(R7wNyN`m[=C43D	oYgr(	KpEat(W,x7`3[!;M<,C.JnS+:+6aO)&1IpRO tE21i^s?Rz,8i1v\a	* ^jVk}>"	
M?H{L_S'bhC42!}CQ &&Gg6JuN&leEm#,1w}8]>pmkYI.DG3lj~<~yI*$3;Mk&-'{,$
*Uc95=Ui#T,QO&pDa,4={ l@}<gUAA[dc1qy'e!*2
.'WFnAl;*(4X 9#UzT|x<#	#pG_%b2Gb![n5u~}R?hf/Er5$%tLL_Gb
o3eF[["mI)ZX^0?%
}q$h\2NpXh.bCm+H#&f>W)g=Yl~EfrT%O-Mbkcp/,,F$c*s9Z(C\`g~s]VNo
^'YRou88cuANafd;7g'N6IbI;0U.50Mj1fKX>A0n]6*}lcU*<
&**JT`(l{QW6y414OQ3Y$.>Et!ViyCc`Q0-uL[Fg'ZMv.>` 	"`{+ef;zawehVrl#X7E~R47%;V;g_\[cITE)8D2vXj4sM.IThvw4q<?\sF^<^PJuW{\3[P
v+sem4|hbk>Iz11}	8wWE0mq=7zcf-<6o-4z):s>@m
PE[s2Sw{tC[34UkZ:2T+?T'p%kWEp0m~+i(g*JSOJ;4~LtO_.k$3
B iDfVMiG?*U.vjC)0!gNNR.-?tqq;"/u13k0[YH~F25gjFH)%6k=X-}9dd][|:<{%/#|]N2L}L!8A MNnWLH=C9u",,mvlF}DJ@f$/tLdGPgF)C3+*B8MV,.k%3Sw*6SK&%Qxuzy:SeK]@]DX-fs3<+pzXYB$]iH3P_ML#Z/'$FPF ;Yf$x}MNo
J0UC|KeWzl;36EEr8\C5:VG,6aCQ(z\jL
SA]42r
\tIr$:kXOYdv45XCx"{6\I<gSHE=VHMFwK1(UX
F).j'c0G`Qf7q8?T8OYvea&Qh6t=xkHYFG:)O&_JTEZY6aYD'\o+H?H(G\%	g%FLtl?lY5Z[^/{s<Uy#8LMf%/<Zikj\cz>(?MRhvgka$xP#hI"vN1H<e 6q\jz9P-@'XKll;0LOQO^Vf5*.&H2=fVuBBg1u!LdP
u/y"L.
;poN"rlM4t<,n.8GVm*ga5RT,Ykr9%n>JdA-v;'$o(T'#2wSN~ H_|={7?:*p{GG)%b:n6cP`t:-5zeR/yZ\_k.CbSb9AK-@EzZ}]A!is=sG8bdKhF!VH`=Ne)P?hCy\DpOx]v:1XK2$f"qr]I/0R6z"RP{#8%F-S@>=-T=z\scij{IW*?e]j]8v>t3[X]DQln~KJ*;rcYdzj;2qCR>2:Gr?~`BW@0TJl}`.|;ip]/5nSu5tlwk|Eclc_vD/hC/&by9YF5@2d<EV6)O8'pkapQjz5D6S>]pE>/B-nA.@2H&J:(tgx9Q|ipHx	!tPf,<0GR#1|l.A|(.RJD*VM$)'!KlFZO"k3K|j2`w{F!rIa"w}HQZLco1z;qND_UH
@fSi n7c`]T!9
h^C{SuZQTzrH>-/lEm|fz]7\Q
O(D|6psx/K*o,W0+Gv9+dJk0V8pS9>.Mdm03?/6N]j1z&[9M%jEtH,xi3FfftyUM~N3S2*W<R>F.H2kC`JALYzz2~ MLyW{g1AP<{[?MmC4jV4f%MDM
jP#Ezg^tHDJ8_0?iKyFx5~qyzp5@<bie|LBh?_sCMBB1$B?m\`XwaKd&!?GIrYm}w%F/\OZx\k9,)_FoJ_=?Tc5!Q wSac:]L	C4g=Ytu(C&i\,C5NkcIR:y3*)
)4PkH,8*[<Pv+'yTwZ1/$)0W}J{35	,\#<fdeJGQ}DOwEZ\K8	duxjat'&b}=i7c/GqjT&!khS_SRs?hCeU$vY8U(1IfAVQ>>?T{rFMsGefB8	={8i{9avuA-/o[4{Ulffz<>Qo;Mm+`m1'II;[[4-4]x%Vv0~>pjxQt_*[|	7DA_-+/]NDb5&exGcZ)0$v$Ae0SnE61k5N*u^CIEWJY6]=tWQikUU1?Zg{lk^)y%-yZ`JTUF
/fNBcVX=OfK6`n
X_Z$KNx1.\gvMxrhG;pDFX8yM(_[@KS#sSE:VPOcQ059d Ui-3YjhI)*K#v]"!TL
&c(uK`@/G4Zwl&ixC%O*lj*(xC;%|].GI> jMx'm|FASMP)]jQb:@KimRd);(/oUU^=.3-+r1=)=JFw/#n i+:;8iQjvjBQ+l,m`?oE/X2o r6S~09E})j|I=XWk#}iodH+d]*8pwxY
z9uKs]#?3udu
=lso/8;T>t{o((E&IjbC}zi={kXXv8td\\,?T5u1H /N*lHM$}`Y<ehZqD!x/1SEPc"S`GP{SH9`$RsLyh!e#~L2TBz>@cVmj_	U-JofN+o`AtTWYC+PR::'@*}~IE!pJyUVOk<}3hld1w}JZjQn/*<XayD^L3)MitrQf56*~t?az^\Ik:CL]PgS?/H,},oF,B:&7'A*;|wGJ|+W3:fYK[W4_b}u#UB0?OuH8=t%1	,\C=Op!ow	`SP;klNWD\Y&kpqDPDD33\\ohQ(qcL"0bKU;g&C7/!I1
xLYu*)-Ii-dJ?48G%Y5^! vRtdRvB1Uz~%L9+J8,"oN2he[V"TW-(E7MOu&!FG1
De9+$
W<~q	^1:<u7@PK/lqG$G+F]^{|W*|/1I@;Jh
9:1daeg``=&6:0('\%_)#! eFt/2]{rMc.x$)?B'lDT(|rWzoW?]NS{<]nM].IzH?]M<Z`w|\RrsfoUq9IR^\^d\iA"bb,T[eSid2'_;v6<vE$s%y4]Pw+7`Lh2dX{9nvAt$y{c5]rgD!+{_CVhi/3K=y>j:Yn9vb0.rBE%-#t?\F641ZCLhX&6S3o";dXi(fnFa>TfMn-hK(c&l0=@On8M9PX2ifm%=zvC;tsa'HK8O
J)?s]IY\"jBt7/)18T0'xm8;y!53d:N##8pf 6O?XoXuSpov)%(G2T"?V69p\4tOj9AW;@#:OU1X!%B8?|.:'t;w0&1C%Okpt CPy>4Z+cnu+yb`NTx>/HorCJg{^%TY9L5MX)v&p8g#Fo:A5"^H&(IVt#;J=%PYmT69WdWpW91kMi5T;&egM0qI?hl5_jP$0611bKwJZ'U:4o8ig6dH,MQ6 !@bUB)V4i-V(W*8n~	 :$k3wO0n#qy/dy[L./k_kTY@7hJX<7!&F7Hh.b]+ia>LEY_D-Hr$!w&"IO0rt1SmZPi<4}/s|EI0AwzdGb"n%`g4\a6HM8-}[A[dDZNEES:$,1!<V1|93ru
5<a2AxtkXIJ&ci
?\cQgUYrsjrp|j+G;=x]YJ+CH7xNc'_# &$_XNb6|(HFa?3A}E9<m|C=7mu2#Pz>DlIUP%
p'O,R}TI>t?gjrww <!K54vZR" pDxN]fC=wz3O35l0`{+(-b2GQNE]=(vSRhzpnNA^t2g\98>U0AD	h;ECyUv\V<Q"	yr]i2VOw7%lGr_upNsC7xu1n6PdZ~QGM][(DR_,ANC(31YG{'lh	fhN+_HGh^o$kP)'MatyYIOS/d}cVNX<kWsAks=H+kCn1,y	Nc~vs]kI4<?FK{af?Do=i%2.Id~UsgvBD<jGNn:	HUzya&#J4hIq61+-q
/]
JwHTCMn2b}e+tV?^2/z
dulT9XKX-4WK'+;2&!Ks7|9\;o1#f_w3"d![KBz+cQ+sI-"ys(orec%{;y0~?tJ0VrDw"]`AkTQ$"Z5pQOvdJ*v;EQMxs
PJTf5?22H
b!q8BVV?'d(McYs4?if;o uW.X9RC+2fS]XZU>Ht[M;9$h*5I9I\]z8y.vTAx~g7yGh;;!b=Q^l{t:ApA`cqi-TeMa=&8]<yGam,tE_(QGl\iCqc;ZY"O<m$9$qE:Lptb5vXGjw!uFF^'.>9]%wmbP7OW3^tT&zZW:Uui~k'&V@j3;`id"^+9 ghs%/PRi(.]B0|K(Qfe;d'b*F_0T'~X+j@N;\UU/Lt0_1D9]-s=.?\i> p<k{Hd]O=%V2a`|4!s-DumGE4	H4~5MBmZ9ovgfT&mme38S,b+#$e9^;U<Me4*`WBdZVT36N_4=142{9:zT0:=Xr7nb%1IX\<I|I/+G7Q!CdI1($=$/PsCL@0B710[x<B\>fz*z7`!`4?;!o-W8353=4N)?p#}')EYr/#iP4[HB)]"gs>w|$.R1!~PII LS	$Htz) {dmU g[Q!Hf}+BSfz!YLi.RNhXOnRb?DL	vCs-n`2DRE^IWTd/a4HvL;q<+I>
tGE
&[d6/"/joXkYv]>K7zY@v1_`'NW^K],MtRg4TzOYzA y'?a*RAyc18.\i]
6dXaHi6DFEhmSa3
.5.Hwvvg
T;FQ3%QJKas,eSwKORJe}2QgzVxA&(eAbt@zDTX[#=ja\u:2Vkx[]]Ug.gFna^IW]UKxIgE[$<UUy>7w'9;jHEA17|@%pdR960sopG[_%Jj,=W^hGiA>*']3P&IMg QEzLFVl`-E2;:dk4
68	2*:v8m*{A50	H<*D#}&/:#6f~%11d,=qEfc5	Vwr<C~%Bz$#mo(eQlB6yg PY/OIL6dxG|e.I.
=HSD6	14~;usrWHuyoy$xFd`Mg;4	4gJmuDeZY7rs`r#n5PzU5`MQ0M_3iS7g.3-Iq}x
pn/Yw0$0\2wxM
7Il#s'vuDKPwX\.:%7UmJdZ[fp;RVt9x1 qd(se:l="6YJVp=[]6Rra)B@j5^~QX'&yfHNt~;_TxAzWX~!W_zOZk$
aP\mDNG&k@tV*iAOm4+TnH#yWq7DF]{C_-Tcstw3@B`V"\2^tJM0@"CATeHW820{"zRW'm;[XXdL>ke~-A6R4@/elmf4hST-|i6+ "5!`cuPi'7k+So>%IQ>h%55%Mon`|q|R<v;y/}{q,l2'v-e!a#	!ZMZ=FVvQVw"z[4|!^	Ii6yl,88b}=BiCHb7/N'6z!Pn?>3`K'F(/ME.Hi\7MkT$&pu_l&Y9	BF"<kzw-EC[tQ7}Qp=CTG]*E<Ot`5~s}E 	,9DOG e[zEP*+c:%h^oVn{vuzy5t}rr28jOzU)lO5@=x\\@]L/hb;L;zm)oy/UlQR4zKGh2,kFe_MENVZ[3$&*p|{"NyM1){Q/[@ujTw
O} WIH>!?FPY~~PM#~.	bVTA>&N&RHgI~`
s=;]uOd\<vLS%),8?2x.VFB)]7V_m	=I*	Hi$C;c!Oba>D0
b#>{62Yc)Y9|&N9	(`Tcp1aCRUEHMQk#1O1NE1R?LqN4is-v1XgMKu<:-i\T?*hJ?Vjr^s`=V%>*mLWp~TTZY%DqUrO*Z7a'LRuZNH`4m3B_2WYYOoBi%xLP~aN6A{!z^K6CM-hI67iTj,1IW&b9QR%wbD[fN| YhKQ($9k	#OSD7[	`&\8q@|5y*G<^1G^\$+UHz	*L[`M>|iAps u5Z4kdP<o-zIX1YoD-
F #g'6fd\X2qf7DK.<iFAcXr@4.Cn-X[91e'AGVNR;|{Hb@g&1b]`"%V{^)	.\?T13cd#;'(%$J;oZ>'bh1O)3K'.Sd}FnVbu;fBN.<4oVoY+W|8;`yJ)e6{@#?/ml!)!	ZM<Gw#`@'?gD]#[}&0.UJYt oF6{;z\\:1\>qL1U_{?@KXegJfX:a'5X%2=i9OHq|*c_b`~h.}oq:--pj_n'r9aZz-j2thhnhV
;wVPvE=K,]+9q@w-	SR1$1hU}>v=%#W8X3GV/%{|iTP>(8h!(m_Eqqx^1|F&ol:y#|wvVm$~,q~TNuu`RyC"v@BJjrNJlgZx&hmr
UnJ8hrQF
eYCd 9t0V$NBfnneoI2t	MrvjnyqDZ|vPSy,C$Hq|(V)<
NH.Mw+.6U6SCVBdA\y_O	r(P6@zvkG|h.)E;NuwX6\?jt'7tUEH[?5Rq1_y:q.i;	9yXR-?@597TL6?w/mjjHI<aip*\)0CO\
5H"v;<\@8Sz:9^@J<T9Ba>w-0	Q%-V!.n=^,Pp{J:lv+%- HZ#czK0pKH3.uu0#Arx'OzoId| Aa71B;N^#m*98<1,6fVE[01F=3{FpEG8J4aYk`6[QOFBS1:;9\pj2F>n`9}0r@F_yIFkgfg9aKP0.]1$/	/bSs|1<MWMs%hQ2"{.ty"y
_ u7|fD_WdANEef\db1b\&8"#+2B\zUlma8"g;q2r[]F<BqXTGhNtV4@;zm5iw]"|lv8u)kv4q,H5h9qyCC#DK&4l>x=ce?r*gS[(~?F8'VcsxOk0,vhpiHukwnH7-eego{vnFpi@b](^y8645 z1ifV=%L#3*r&UofIWZ@59d{'h|b:ZbNN
e0Xl]Jo;t[/Xip9Bnzx5
+Y$UPF0zDfNb	[VOC2AiTuP6XZCD+hnI1W"dihM9y	&m5(+;Ge>nn9E iUG28.CW}&++-m/E,bY)0j
>'\%j&k'zB'vTn{{CVyL,1gas8mt|wx@O9jr0fK8wn9T]e3{jYf&[7$jKM{DZ+(1A^tqBu\Sba
$Gj%fnrtSLQFP~4dB~xso-jB6RtVjD",]I#Y>.S_9 |H{0^s7FR"_bQm&#@>Ic:7fO'aU,s	x	34L'm,(xA@T;/s b_ImuQ<&.%kT
!8^'?o2*FR\
q#yS22iV]55/Ag;N0?bG)z\%DwTD.XKe_wtK{+Mb8Q]dkCu |Jadq<-,=`{gr{SXr& %n;32?c>^aws}a{V;C?S]|"0F,C7~=,#cOXoXm]ufS,>x?s7i?@L/f_	j:">|viW8WPn*N	.(5{^jgA}! ^AmURpz}Q6.qb;9hnt/uW\N!PKYW	>-)SD&mj:ReoX+3Izx_MI9x5oU$er{Civmq;tro!!PN~<e_T29ri^MA?JY /D|XPUba.gY2MU@d8M	s7Qjs1&Z9q:}Ntxf}BT)J"K>A0ONO9IagS+Rg2s##?3)Xa^Ze%y4shpOpCs(},:4U+em$1zl`>i/9+O.#.Mm\_Hz3:AB
pI	z),X3XxX&6&u[9_.,0ix6])*+yJTf"gQCAAa{:JXK6n){t?q}oc]4(gB/~k#lq"f}H%0Z)k~G4|*@ .8Z^.x?tJ@-iLj\-"sCzYE>O9Tj8L'jj|NeS2m<*\+X[u/Jht}M]jP!qc<C{ ^}9nV,BJ<r,u%w,^Q.
<.c-{tWx@QR6Z<(Y Fm#ePDnv|zB:">+/6*.V	>M>e<Tk~;4c4^sJ]2zPGs_o_u&c4]wgL,
_)}3]cPg$f:,jzVnlZ7]2k5b<2Q7'rpa)*hIU7Ov	clk=HsIZ"rl6-{bITY:3r`oh8/.1P{Q|Vs(6]{rvzMzy	2"Jj"@P]e}I	kMxA"ZpV02M4-r[wpX
E~%/2=6Wx^w %v}bJXcL.<pGU!Eem]]Sp8C=.^sqbM<ka}HrVu=(ugxKrFPSm{EGG<,|92>jMLm$[?)MB+]*$C
In_y|(mkY7a	kr\H]i#c(jc~6D*j}_>Ru`L!6x4s(H{.fAi8x=<F7O[I)
Is'Of-e3vG<AwU6~EG?'oxcalbxM*3ItVQ;!|]|DF*3@bo.*q9('XD[3!D1~uD8gDY&+~
JoP
ThO>`S"Ik^}BWMWsLN~.IEGho	(&z	YMkk)(yZZ FPBY&""nSc/JT7pxlWMXl:K<	%hOw{],=t)Wf.l;6G_@8QU8D)R1JP.5C.$vhT8rmqy__Iou%h1/G_>|_u;!]zd^>F`Z>9$MB	`H:g	Y+esM9ngvND/Mqc%}(02q8&1pM=|P>["k/#}Yv9IXPK+F!x+F>zb_!q7;|rf|;Tj1	LN&nW6^,Xa:MM<pCr z`qV:nkFb
'w9nRb%{-(>$Xu~O-@:xe"9w_dcs*I.P0I1Mu)cc1{\y	2aL|nMokGd-+z>7U*Pe_8tJXZW;M_gda(\|fcYL>]U5Q2N^zI~<":/
]*igjQ.}=0IY,2CPs-%J
~g8s|&^vS$g7gO*7;<r*mmnvt^=+G,`
/ Q)Amsj'6G^wI %-@p#o#e]2RILm+@b;K-zj/Xo0}?ue	 5aM]BJ[X-A}*GJ%HE7R{Dry=(I5"I wf#C"S XUhsEL7,Ky~th2*{3qSn2oLru3/TIG xn|`"b9.#5E]}Y#3<=z2m?\oxe_vJwWLWb4'tqQ5.{\UgbN2OgN7w>
E5S4jX7}& @LjG8Y@~y\aD]]O#b]@0vw{y+|sJ~OOWgLq%X5gco.24l[3{0lm{S!R8oa[6m0>hY}HGb~;T I/{KBl '(V-O{,M=Y%_@3E=iYx*y2f]4k}xrr{kY5Z*]HN=JE.C&	Xl)!|02Rw7jVCA@+:O(v0EkURs7;s$k[+%>ZVf<p?8Ya# 7UW@u?u97,P\^t1gL`29.bRvmq}&jf Mo	+B
XhaJ+\u=ZE^RP%^6%RE~*k0$Tf_+F$51h\%nw	'TQ"j3@T`Ai"N3_J#P/(yODtVF)7;
lpW_*oLaFeemLj}Dq;gsb&:ETV`.Y'5l<fbav?<.qpq/-{I?Wv6"i2a'-$5%8+P%7b`-S_y=;E	x;r`%
,<FO(YQ/d,T;oVS7D<5ki{02[%em;oT'7qo/#8l"HX\_
xLf]\}E5l9a>)bhx.Ru1zFHQ8)>+o$XZtBsRYds/xeYT!qG]a<%<jJ#Tb9av:^}IHN
>*5CF6OX`Lw3,8)/yko-Cx?wOAa ,$Y]CTJPBAo)?1MWI-xBdHB4" Yjl\7w$bwP{V$$:&"zKYh$IbViFtk]U+MteD	B4aXXge]CzX[(AR`U>9A.p.OwQ#-&^=>-}Hh	CvybZ,9f}- bln)Kw_^eh{4
7-zA;fK0B&OAUV8BB(/f=!XiOX;7*_QC#,yo$e219-(o$u~})qt:sAq# \9}Y/Jw"	&@UDOn{j
LqTll%m"`]"5wR7~$koUk8g7fXk6/y+fL\#x]["T$O/7_boZt8=~OQ0=	bvL-rG4)4NKsNY[	<.r[ "F@#ZGp]fE.0^8k;|
99{S;/*t[piqr
SeU`eT>/+!liP1$:]07!Hk7&~N~t'8Sd#qh^|D#4f?|D+yWb022M:Avfp!@=)&6'=xpb^
ut/(uh2STqn#$1F%D[\,G$.fdi>D}Eqs`%i&lIu?7},EOTKg(\uD0B(oy]4nW!vfYWl#G)V5j"W7nU]s~DxTwlo]_}8?22IH~J/KH"'8es*5n HB5L"FLI,>lA_D	ut!>LoMQ"~*Ss9iS&X7dx%;No	16nXT3c9n9lE3?:
z-*E)4O~"&|,Tni{`$:#A<ZSUT9T0&H&TOpG"YlCLk5YX
Z9)HTSzuK/6YC(n;-*@%e.ZIv>mK[I`"Qh/(noq	;m"?`KE2|?ukS[W<S/1U^WzqQKb,/UR4_k(+i)lWWx0Uh(xz7Ar(J,3	Yh59+at'b40f|9n@w9)0Df?"HzQ9q\|2= w(+?DtXL\<7#i)/2'7uT+79/ nTv9_i	g%-k}6ICR!>mkeqNII5H=[1=A;B|R|26RUU[eKc+$@l)Y( k5@0{)R6q:*vK[DJBn&bu{27fsG"ZhZhyLwX8 T{#cw4*LgY*!qyl/>62@9.Ov]@ZI{,4f?>$&BQKgJ!:jbK.?]QYKFrxkK!J5Brq)Y6M&w#C_
cs/B;tM]L` d~dRg0ksUs1gvJ\C%{sS3ml1sCE9-Y;gB^1wY3OU)oH3/O%\dEOvQFA*)QdQNUBjcKjMtK?7MYCRJ04bXev]N^c2+<rwc
OgW>yF5')s	&E~1HYQB#KxGHw>"rTkDP{q`ca$$_!DHe21IjNQxfI\/QX[fpC=hJ2jP;r>j<Er<(rz W;XWRA7A8 i^$QwTt"t

>o;wyLlz$9=bnbo{&Kx{E4Z+%5\SH)7Y^d[acC)l^Y'cyShbq9KYP0^.N!eeEL`iwT9p"RIGUp!$(LrzfHLLBa5.cZa\[+;'1z+_.i!kKo<p>`EfCATUp^/GUe	oUB r~#Mz)D(Bt#k.N4-)"G]R]PNTyM{^L/YtW,jYA wEYCkSJmF)A::z+>W(hX._c{h5bK#v;pm!{0aF6$cooy_#x+vL@~03D%0Ie;(l^u2pw5JX])B: !d.)&yqap"vz)dd?2Wy'zHaP=|5]		\COD	<}`Au:ln9Ych\"~H4{0':-olW)DEeSwnSd#2]z=,jw)b`T89(kol/fv|Pm@ijXW;R'irt5\!Wr"xEhz$e&I^ueZ63Zi6r| ^F?3o.fdp4dLjtEkvLwSX#]/^k`&;Q y5\=)r	4gmGQ9IS`,`2-|JY%!'{#VnJ?Gp,!uywRV>v+pW`x{Li7>0n3RuP5z
t0w4+Y ^3\oDs?"N%#o<{t]2\3e=x'CTS7=?'6t\>>8#<2qMR3,yl\%^2\PqSn5Ss0Kz`|HyhmpJ&"8fg?+;SGbh.TGSzX*NAl; jE*I_p\"&8xNB-kYvca.5su[Ic41YGLI!jSJ"F86k(-#75!;^9|u3O)V_"Vmtf?\OhlZuw)41!g:\m 'H{=9#Ynxc? Ay{~;kYR7,iHuzq2-fM"~?#v1[H6_4G~':e4	;((KQLQln~[X|U<Y~n9rvGUPI7ieBt2'Xi4wyXrki-:]>cZOn[.0]c	FS0RO4KYVeI{w^M@<342yQ=tfH:d@\YbPoS&,Vxp|THFWNCt+
TD;*,ABPV@ob^<:W3 \}KXkVyTPF><xPZMCWcj=
]V{'3JT]4s=Oz&M\9=keZa16v(2r	!ll^W=*t]R=1gr	7cqELkfl6fbO|)&cg3x/XEN`7Yv:_bl3+BdQRcdg-*XQvak<?qDX$WBp47[Vr8)#5Yg7*Zl=	N.~L9Pl6gNSbP'[z?
')RF^}n;e3#`R>`e*csGz{nm=itihf0aC (ezK86mBYo!"qAae+#<sq U}*3:~K@?Tg!!,;1`6(dh*Y[V&=w7MARwm-PYmQxeoYB&h}AdB6uNE$D2J{rb6eR>53YoGol	X~@RSV+XB"nt,Y;~LIN/Fef`[w.	G*@,OmsmJo&~'eA2nP|)=qWSfW2YaU]o#-cP7BDf1OcoazL+r`ZuM5J!Vd=&HNy>$aL1JAE_0XApBTkUTF@y,/
B)^jL =Yy~w	bqDX3~2t=v7zlOcbE{9>lSRkuc{D}Q%@P.3.a\Vnft
6t,xt~Mdm0Q<H,V:bLj#p#[0W#?L^
Zu6GM^1rT;DU2!4)f$CFoiH61yLZJ4?Pk62;[?([WCK]'bU;F-N>)hF<w%U)A,`8iz9!Z!>dGwD*k2urCk&hYy|B}(<,t(Z3A\B
qPsHiL5Yl%ygKf) EIgh;8N9VMns;Vpl0*de!	SF4R7^X|MUa5M"`?Ue(Aa<\i
#Qb$[a2+8En=nYN!|xopP)9P3[`s*s0bJ[+4Mrw,%nQT C |K%Bx)KAUDq'$R=IWFtlPCvv;%cI#wcfU;O)E@c:<`y*]K/5P5|~N?332T~\InjR;RKBu7B&}	W!L~7r`u_XoTfq9w$8h1`.tlqPJF+%0Ykoi`!L1--hC[>9KCRY>:$O<7$JwF >6zg% 0xl"x/0eYY,^hg2B%s@3<AhBys'gXRN#JmP)mQ8U;3pn>V(k>%M2yB,|GLg!)M?vN>V(qH;}1,u<]Y7(~wB\R8"")4j~v!d(pNw	:Mmo,U/TaZ7o7J&aHWxdX':\g!)Z/t$I}*MkwelH2Mh%b$f?N8C$LP<Rf?|i{Mg+QN]OGtGzrlgr	fZC,>f'.Ij=@BRp!<-*>Y4;7%"Q6}4
hfI&BpQ9uQ.=VSpl:0Jb_n=2 whVm B(65nE7i0ulE@^i4kCZU[8eX?4r.)6,KaJ}]^3+/;MIc_HCP8x0";DWMCJbQoWt%DQRq$L51bS#/X}..m-^9WR|Kl q,V60JE`a$"hL&}JT4k1n?c`%-"}{i^
Z8t]JT&;h(rmt#e-7	E$L-QL`2cyDBB@t/tR`6l"CGPR?aZ+wDN]v-Mkm1@"g"M,'9Osr/bj[4pLa|Lv0ys2Nnz>?A-Wi@f^*kcbW	nQJ+EAs-a$lyce7k&Ej'y;v)s$ d;;CyT)x(M4H)F/Mej_>[j5O+~eb+u*(I@{hRx>gN]lAqj	4w[pFz-GhVlMvmyx":y}nqmOvaCx?LQ`NG2I<d+	=tmHJ 4_wA7{' 5UpNoi	s@Yq5:v}TuY_{e <Bp8_?cG
fJwv0#Y&EFy"+ p8Z	5v0HTP;[FBeV5>/sh$wg\s9}@O9["a>m^O 6>`(JnvG4fW:gCX(]x'=dd?2ONJ#Hr>9O*sK=Z4^csNSif_9TJK..$ho8M5l],M|nRQw+I"&n?TQu00jtx10Kl7^KB#*,(fx:JH8q>h~ +B@IF(d-19T[.Wcd-&3Y>	!7X2w.p2VJ3
	<.