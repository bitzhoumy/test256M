TJ8{4E?j0s(jq%(R,49O>]h_HbDqICH2x$CINFUfTgR1r:`)\` %.Tk=x+Z!5SG:H`Ai/Y$fpvA?Ho90u_/#xDw?ftc'GBiPl)8PtIC oQF{X:.xy6,KHt[5H-M:`x*T-y#LOaW;1_H{[r#;Pl}KGB^ZQ
ott^tEfp+gUz H*Xfj<#t]jM!;'	[.x+v:^!S;8*v!/Q9pbkL>4(O8j\NR8\T^9Iex3+Ypig-+E[VZ|yT)pDcvEv$/|<rua5u^%0MXZ2
[AY\5z'*KN?FL+Wh-Cby>wb)rg}+3{^`oL>&(_R]d[R qH|s';6>^2Sje</L33ENq'-ojj6r7Raf~b.;Gk(T>Al;X/g-K>ea%"0F(,0;E\TDa{UKNr)XtlV*i'<l?4VZIpb\X-]v:CIo3'>^}+o|_ZPkRSb?z)H>bTb$)2;{Dv2	m~-cM!K$&@!u	}~ixosPIOKaFxI6Q	MZ88vEnED_:kg|/Q(k=]&3`Uj$%_b%cWf"
YLqa+nMqJ4H9z/!k}P.=-jo}-8ftiSi	9Tj4E&uiKM	n!T
Vc-3lN2 kl+J(aRO	0ft"`@G"/Hb4,D6`N,b5DA"+grh-n
@kvH:=k-`2OE!0\:*a5]l'DTjF2(H-Jmkl1E2xZiQ]Q<zTs)F7"7+sF?O48R{{BLG6HLapJ-GDP,6HtvUfb ceyWY9 *W7M+Fe*E9_8b-2,KA4zzNr-#vRu?WRd#xiDd5n``U:peOFIU9qt)<`7if0pC:/"(2ON|\b(9U+dA]zu9;@{WZ-o.^[g	e.mA3Kx)#+f&^ JJ	#l0NpTEg/cBAq=6tFY4E9jpB7ea8NreUpp$Yh=8f`FlqM=p1AW'5r#j.&mt#)pu.DC.9r`M(f~I,3@@y|)AmOUnbc#P\E%h9]]r2Jz/&1WI'Yf@Kme#x<}R!Q[]@:-fR+!Mxrnx7Z1%k72
Q
tJgNW8jNcEc9)\$Ifz/dt)EOj,.	Ciwy|S2kA4qJhid6x' R,[(qrlYncQcPQN|:AGXVJSa@n
uo] \I\6`D'ZWHT`fU&
N%-"tpY0@Ud6C=MV4El+9Tp&\ij-t>W15dt{R-1F^q/Xx4 g55Q*}Xwd [Jp:|WT.lhzCs)GXqa"!%PX,"k'#E9xJ?tr,oMhO$A6S&=ZeI;T~uE5iUW?`Syu[-i&28h%8Pm>KnbZ7pvgN'!gh)Hsd5~&$E[*uIOLoOt:Ny!-2'|o=4(oWkWGMe=pOAD_AQJt_pQXdk!$.
 b+>W"Py/:B1PH?h!<8g-"j1m!b-dmg#MQ%Ofl9`,G(LWRd	WRi
274V2uc
^}qS5:.6 m])x4WUb#Fc`tn=WLEuCb_'7~O?6VuCIl,o@xC5%:du0{;yUL	:@xjgzOQ0rl=fo}
TVOBh0gMT7<t@QAm'6-TKXEB K,L3p)Y?L^/8%ZSl bqe%dx80g$/XCz+oePU(Xccz7n{xxwP(ua<*xap0'1umq1+go;~W0<(.Wi>+74,P~	8MDXF5%TUJAi4*7hyi->9tVw96:>5Y-UNGBH?:FyF40s<f6i!6@=aiS\i]iL[Y/bQc(%]oqVbw9T#,zuen`^p;>cPq=#*]c.w3/2&F!&7^f~a+:'
M[Zi"<reW\tRyhAU'^Td 6`)O=9pZsFpbJDxUI<f3v*h<F"Ezn>n_vsCm~Pp7WP(Ka	
BIXd4F'nbR"H^R)Nn}3R2[hv`gjeaX(oAC	P3<o2XPSNe>&+eGtu9Z$W$E)`41=	>|bT=KoV|X\m1w--5U"|./Pq-(X@N@Z^;C@) a?o9#/9~6p%@"tU29<m|r|\tc%FXXC4Jhq/Vx(*m=VNiiCom(TFbEwcGM*.y'-&Ri#|lj`Ii7z]=xR~0sd aWq|91}bR[UW|@Z
E8jW\'	FLt!\iQS'U99}bOE,o{9I}r8
GR8o}
S<YTc#?FahK/-Ufk|Kk)J^p/ opLeo+pr%,)LG3N;pq"E6wZpsS+O5x?LP|e47C%d`t<5wKCqL6X@ciMcFx.sArIV+U2RH08?StaS8Q~t{8zAe$Hf4kd 1	\-8ZlE_jC#hLQDhVJj&7T /Fs$9WN0*S!3},t^{2>p]vIMqt[h)<)}LP'f	w8|t0X&:i2|GSQ:]a(K%aWE2^,$`2A103d?hX?hg^#%l*bs0$9aQNoX<0<Qk8a\z=o@{G!,-VAyBBLpCW0uxokSci01HSaKzAM}Zp]I&w6+mFeqxz.PW2;l=sqT"DY]=v>D\JL~i[]?=F_XFH[uvCl'@k+Yq]a%ahtz45IIajFjPEvtL[?"#[RQ2BmKwKz\d0v?8o\A4a1N_-_=FUygWpQ~.aIb	$ax}
F-" ^:l	^M\0.yAWjNFlSK5^9P?qI^r9VD72x4q2*P4Wr]1/GU)p>IEgooar8Mc*q0d*cPMw{J|Hc5p.($j(iJ\1HJ;>
T7g~68Cjl/:$n:h/0YXP"J[+D_"{/}G|dk~v!YlA1 5]RS);=?.|Mn>2upWOX"y)<>U{a]z8o,oz#|n6bjuy)rap:ccaB	yBb)2v@aM`:t?t?uK{nR-H{CP(YM~CO`0C:0pXIl'^V!s:{T_/v?/,EK)tC//Z>]G|lF8
Q
yQd@6\6_gs+P{"HZ,Do9J#E=&$gg?i=I?P\zk-gm$:N'o@^iwhm)BOfw">zE?\1~?X^xwnO,4~wO4P$TPyT#W.Um,k~viC

RJ8Sf0L}#4^ZJ_qj_-?[0L+= ^TQ"XH|SK:[EKPRQa[z'=2(z3?'YU_`ve	$>3,bz`)FX#?c}V@Ij1[$Z5DwBpcZJb*c4o?uT
w1vd~
ydSQIN$1;Pa^#x<?$fWN" V4<fff.Zi7/
+D(15d75*41{ufvzRuSnt3`M}5@O<vvQn3%HG<ZA\3>$bj>5KDr&tr?'N595/i|
g'J[~I?O>
jljW=s1}#@E)G}?]<05~5j\"7@+;~\y0{7e]$w;U_:lS:4IbDdOY4i3v#Nk'Zt9|OCh:3}D4}T#}}gGMI
jpQK3kVma>g,7sS=LS^lOj*Y\"?EOxlb*g(C6;88\a`s*/gZ[1*I1N$+q*]^`.BQ6w]D8\-`UR9A~L^-x>,%lF+V%@Tr/FP!>'|%9:eb1F6dyuNJ?=WE,T:!T~mR{u(@/zPL4TG
\(c'~T4`5kfZs0<j&E\0-VUT=h'[i!jYVb@>r?j$BS% e~x=-LgNyNFH|xG~o./HQ9p;O?kgK?.l$'{/LTu ]*71qhLf_CC[m?`IU2%<|Iz>&gz@!1Drp[rx%>M1}'i}C^_@,)8A	rQz1CX0C*F[yX=Vb$pMGr}bn8Ou[6\QF'V!6)4h{.wP
d%g+zWd=:MCo)DDfA4r>A	Q(0KNd7Gz2\7,uvSRt-:]cD`=?!>t~!qa.=
*)HfXD',z_8|ZU']H9O$~[u'DSARLI\_f`G+c;_=@Le\7u7dc!<pdeTP7!n
/r"70*;o/*]%^59. KRw#d}/.~#zf7a!:IyHut>dv%LUxz52ZIJ;YeFX3z{lDd]HT3>`z69%^$`stbQ"cglJ+eJJ 8-'c	@`-4D"q9q[g_.~0Kb]omg7ety`{K"E ^)Y)e]#R&>j`AdAbQ;jpVA@HEN8;*7N|c]5I!_VrpgNrYraawy>A3DmesBWP;>A2c!aN6ZQ5~;>!\Hl9W9$uWVC+#+>5+hd^pfb2,M1*{w"TCm%@1?hx9\@24V:n(@Ve"g3:J<&:6a9IukHDMr~4I\>vLnfg`s3Y~^k>:mxohy7y)2J!T}c>;CPP'i*[T-,8E]*Msp>x=3[c;0j)jqGZCSVH2&a`E6+vg@NI*,l;R,75g/rmJ~EJ8GytZ+Uk_@Ok\U6y29aZU}Y?12o1'7[f0.aT6D-1#=cu8J`&R<Db'O=:*<e#,/z|O]	!crs6!iIk`-EX:mX4B,>8-!nvW#6=S_MpM	{QiK+E}eL&<Az'`ZZF_iFE	hzhnKF6z4x{?]`O/9x"M,%|B!Z`;o%sd{77`x1Zg2/GD?/n1"z&Ng"JRo][%fEYfs	Snmxc&8v-Kyc|6lfwsX!^*[)VaC7+lU-%|wc5TI&rd'db)R}Y/N/W)Iv8>`mpUS?CYb!eu-rF{R-@g^>p>:/"S{`1rFI
{8KNt~TXAUK@@pTz>	7;oRh0JhE[e;Ul	a*^kBMT=H+g{3C
QJi>r;!@Dz&T27rkca#2~T)l+\gR/v=K#x@`d(y<N@J-X)+]R]?f$xRAy}~-
Et7L'%[iTIul$}o>4zk(*<8C<GuZK7R?v@^C&2R"d#?'X0q,CE["!D:hS.nvF$:J4_W\IHZJfeD2^O15FOk,ygLs}ptGJ(oC*^"B0/;7r%]Ojc.yJR^j3+sc8yS~5?Fi=2xj3QH
{nSu8Z9hh2nup#`6m+12NWbBQ\b#<L]"DKl>(f 7CU*8I+nWcL"YE`o)u>a[gEp28fh} v<6T+dPq	urBr^I~'.?W{o$[xhxhj98YgyXpZ<1PNwOz=H"UumBnfKvA8;d1C/aPcQ*1t2bx"Sb({&!@"d
+GjOsx 
*[-n}yjPJF6]=&m_{{)u!
?a
S!*l0>b]r5v-:z6Jy(feZ0.hT|'G>VN0>@d$"a6FM]fYdbb|`:)PK
0( !i1>;S':I@N!k(R_ Z&6w&p|4UVzwue3or6(u[s;	E}5_q#@>1EIaX!ffJJYHl2%RO+iuc_38
i[[>`G/AsRVeV43\W^<LP}
xGet	W#4^0~`#Qm?/R0xSH-B`4\Jc,ASG1pkHq:SJ.CVv0~mr_>	!QFmalFPgW'yrmzie^P@ptG[&ETi!5}k>j_[^re=+efF# n	Z=.sLej,=q3Ra9-5b91'\=&%Z'8 m5=&%*695!G+9tC	y)r"QR,0{>b$fi4`z!o8:p?fZKsu~sVDyn2T5JCF.
kT^6u=uGtQ.c*v F[ME'dT	>R2zJ13Ge~9\0XZ(.De<)A\ro% iR/X(mP)E9	Z'\D|u,Lo{^`%IK@kdd[NV A"JsplH*Q:fU{}4aCwxi?eQk*G5%;aS%4P{KDlM_c..B"{I/kf]<bILS|L*jX(Ma4#IhO`,q_aBuOL~J*+IZn,T<e1#c,oS[jD.b0`'>]@U9l %".C_
1)26pvx/8<yPxt|p%z\iBB@An29t.
y7p}`f{+B
C=-?T]`x}z`Bg0k7*T{f.P#9$d&lX	%n7Hwy*4T}K=vL0;DLTk\5Z/I*8vLK| }umPdiR(;+(U^}$uY:GYH7
%"Y 1g#uUMXi:=}adysd$')~8lj  GVG,!fZ{Nd"[E-;{7L|FO'.Jtx;n{/J-3nS%:vU58t8x1nFZ%e&(M.:9+Fk8/x$sI!q3'bJO`kd%Aqz4VV-7T,d[wh>%pf)]Ctlr{.Imd(S-e?T]u;T><(0mq$m.@@TBYae@q}f(i4tg&0Paos`nAp)Fl
\rlV#zm$*H2RFcB=Z{D5gf)	ToD2c,K&l}!lDKf963\[f$T$H}A/\E|h;RVW*IZWmM/|k33Zj$f-L~e$(?KON<x-R=pR`]VB6;N6tM&WeZg~Ym2;LfcP_pZm-51Jq_3OiM	^?FKq1@5o]50Ec7HRouM4	A4WNU ec1i~rKR'Iu?Tv!&YY17f6t?Pk`9
>1DZ?62)|QocQD>qp`ucQ.QIl/$hbh^^Fn9#Q%.@Tevf"[}7h%AYmo@h[7#$s:T3X.WkpAU5`$\-t/kL"i+^l;|s4wNV [#I~n#/]>)7R]\yRmsv)axS0WBaY	+2(=sYdu\gc)olU1DtZI0.G! G:mO7H)yB!?KMAW_`WO^p$dwuq<\I`|G?s'AXZ.yWn0=$S)R.C#x5pzzg*iWmtJ.[2OY99;<vv<U>)I1 GHCP3o4`:,H0"'A>DOpK~O2bD^Z|5	?T>DKi_MG5y]#Qjtk	4"=tFF]&}_HZl)`<Nm9&zen;K5\]\BV(Dv"B@/ mH|>#8#,3P<*Nf'gXtVDlej\`u/@MXU/WiLCQL;IPh
ow<Vm]3oEWy#'xZ!sMQiJ#f%	xF((k$=!D
BQg=/{wlK*2>hi|oL1LpWyL0r`=C?hV<-#H/#[k)}bYn[e|RwH0D5~UM
_ddC#$^$G|4RBbSt-&9?}ruUVJ=&6~Oj)c(|@+BMDK*_M12BD/R'R}:YT8j_WvX'XoZKh:O:H.e'?znz8P~fqq
(te/QqiQrV.Q4H{6@`C)~\,{E2)?0">bV7c9*?=ZR@v0,P{@~	fd8;#3$RlKar8g_9Z.~YF,z=&zkV5D=ZxNF[D(i~LLJPj0\O8U:{% X6bvlVeYM;,geqfvW0)+\nFc odbo_yZbq]^^l_K5q.I#5v~s<@Ka5,`bDW(VCIf.1V"tr-tf~0R. uhAEGdbsb+~V;h|;W.9`6/jfm@VLUx.3~7zgIU$z69\gdnD!@q"WpQF=yg"O8ABb\5-q,vHFEbj$$k*ZV{M+ng^y`vm?-),btM6QbiI%#U	Tb~2(Lyj|J*pW/
pzOiIw/I|
ib	S82)G0RB-(3YsY\w4B4ZqWH:Q=F{"!0RZdwd(tM##%,R8RrR%eEO:cEI1S.(vSf	HE)%K(7cSk_ZJLo4!CAHq3'(cCgz82.0m";:[n:!!DUii6D9XFf.y,*J@Gp[yyF7NbkaWxD0g"<&m>@P)Q2LN`Z3<c$!<GE%mJ<Hflx(:x!DehHkD/EET,6..Q^HoA4_/^u=T:M!u.,i:er$s\SMVeh8S-XdIy.DY
NUNAXH$vE'c% Sf'?	dkxmmH'/f38`"0*d~0q*GC tQO5ZC6'<^n(R#=,x^<OrFcVyL6Ko=yP4T$15u%^+kx=8MO;p369\=^c\'}g/,@B|JZo2{hIx(|F^96}@rHN_t-UAlc86.zn:) 7@&a6IEZ?i0;Mn,1fvY{={E[TP>RM*Rgble\EE'NDSAZ,DPn%r!/TE,I%koC=A/7/)iU[^LP
9?)@1xh"wIiw	'tD%AJC<x&ePlxNkbWT[8>`NP25'd&{c#s(8<hNAX	kG&ojuo?KsaLj)nr?QFXv;aOZ|MzL	p_,>UK^W3s3	|A~v0}\^m6_Z*ReFA.(nhztx,}2_sB:@MbvpuSS^HnjR6 0s "h7^VF_HoP6opmeyv#4j<7Cnp!,KrIF"#^OV\$WT+Y`N{J*We!i1m&3e4j|*Q7oP(b[|>-xbUyq[ivosQy_1F>}:UG.Qwm&d55qdY@{X)skLNcB>d{`#I6u5'1htT*)D#KgN?h@H$}lfM8.(5>AbF/&%;"%[
bj'2SH[=4mQ^3COAd\.o~|G3S6XouGwXn0S<bh;l	Hod+]0U3DP7c}S$H*@pil@x2mi35EC,Mw8Y0Z@=kLX^iJenR<q\[Env|X[v78c!_0)#nQ#hC8,&ur@;;?e6^;3`Nfi5Dj+X9EH&D;t]f]/wX>eSTw@?;KbT8{9;%$1yi/[1cS>?0"\xe	Z PwO9bQ,3De"-7QV-u6oFF~]ls)xjwYl,4b:[t4?EO`Ws3AM>|,QtfXL4LLI'hE{|Gvg6\1EnhR|m6o\)TX-:sSuq|p3>9Fb@|R!nn&N'\';=.@}t64g.M^DSd	CKczy3a~IIRUl)[=V/cl: $_`VCA 0kqa5wWiGX&[~	eWy&k+=^1C&mB: w89'-	)w09)Jiq.X	6L%hlz}D{s(jRwsY(gH_59Zo8?mX=:Wy>z>c_z%M!dnSYZ/iPa:r<qwtrQe-AfEX;_/LF=.W0SBtNpX7h7-M"OE%^$g85Xx!_1qJ ZK5OF'_k#I}7E {"ZNO"%RX)),F}RJkQW{2q<)fp;KW
2_bFcm*y{K:_	rcXWgF?"`<ayW
!+Wq|6T:RjK-2$8(0=-P6u7X#.?n"
-F$V+_c+Ipq&CO
W}E2}4e4}wE:HG	0|=<>e(/j]X|u3V#]Dz@Z cH2+!qn)x.:\-Wp=N(8NpM{!UXFb]/f%M&P	M(P{`QVSs/7	jW4u|g\CRUr#l=l,A(UShCP9KJTw?,*!mS+Gx3{o.:`Vqm$Y
S!MFS}P*@`D7#\<[&	!_`$9wh0Ei]u/l!F=5h0qB_AE8SP5ejHZa@OLx~3|E]}9<t7;:I=Pv\HAcR60VwG_(#s[.TYI2\t$My)}V?$Hkri'50nuz68Is6pz~BJNgmf	3EHo2b[`5#"|o?,;]}PkC^^f+i>.uvy>eq_Xgv_`'lrZhYR_R?>E"O6B_{qi}t<"="6idBIcOWrJE{8<M:N	(c%e"rPjd*_LVN@ej0PWKG=UuGA*eSZJXcIgc:(R,|}@jK?! 3=Xm	M
v-"NH~=ECaO76|&ge-,g~zG%VScdq5L*.[ lx,{,rM3Dv-;!>Hy.W-H`;F#<.V:aEwv?n]e\V]A7*$</1.j.*o76/B^h%qYqlkM`X|Wc(3;IrFQH+q1F{>'+{4UEx=BR6|!%<|>j|Vea<=o!oLU;"xP*W_^_6~b>\F$0QgLXm)f(Gert|V8+T~ycO`eR%-"\Uh]:WF{e%jz##qGu@DJ6"+=QDMfK&4jsJ7'.Drh'54F
d'>?B"e2(p\9tdY|_wx@Rc+g,Ak{,C1n342,+&dlZ*2@N8{.!k#}28Nk&o#5]`I|f!;<1Pd1-A^H=Uye1foA=#p-unbJ?WE6e9=	OoWlce[IHQPx1Wp;`AM=>,Nkaw<u#8+s:21H#\=W[,#8
F0ghPP00ApIeB0O+%-o}@k1(SNcabQoEy?w&U4->L+9x	Gd]-;;m=Lm,N@EU\5RB2Xhzlb^xU_9ZF6ATU=N0@kGSkJ{#DK'QU9V7t](8O
Qt6qYC)BC\{d?	XqqIkct5agon{H6{-HkkrOcTJn%+iXV3p2ett_M1DoXJdaVK^au I_.
)LNx8G|Zbk{=0G,v7Fq:B@cgvM!sE+oP~=1I>bJ6al;QI&/2tIO--x-NZ	S1"U-^qFfOJzyAo&B(`8f%fc%e@	L	|jeg&!_,&OKR\=,ne"P*Y/mx"(S#iV4nrmp($-8onYRBs7NmOPd}u"k}qb6u.V$om;%%t:b\IFu!PD"URR'mRS+c:Hj*ecETK$Tw6t/3hS %O[v`mB;Ja3k.^*KzSn'k6c	59*IOh79mE	8vO.wbzmC"P8^PT(Jvd#\h=wn8jNi~?k{!CXKlyPkA`rMBzPkTD\c1N#fF!qnc{g!ldDatb&y_`T(H\Dt`8]PUstBOlC;e/%%Y;61Wl,a]&0vL$20Z:	xH_6R8f&Cx|@F%[~&Y0%$jZuwTK7ciTSOV'+T5mOw~/aH_@bLr2tM-6lb.2<oxV`TPn[k&RUI*H)s@5?;
&0Q;R(afVyvV=^]["K^hV	.U
Z*-[4ALB=],6ab^fS	*nnX9Tm[96^9n@bs6?7w}I\.Id8p2;*y3E#>Qpuk>ae9Yu!#Z,!-;S]ZA"'JAc$i'a}oS$|6@8&|P[|8\^1:*+<s5-A%Y>"`w)Y'(z[{^Hs'SJK-I	'Qy.kOn~4H8`	}mW/8DJCuD(wfMT`^FI5\tq&4m7Wx3xYzKr0saG<zaQLBqXRI94cL@a&m7
/X0m2cd}x?LHfv7Nc(*an*oKxfTS+;pT,?	I=$	&p<":[8Ub3WA^<~{SggboCuZ0lEzosG'lI>5d2('ygV,xvUL")l;3wStUoLCzELNhaiW:!xH3DSOJ8gHfPgVy*lk&m7g`;4S=3y$ pk/7#b2!KLe*h8t8	 n-Y=EdLR
CatX9"L{J!.ll\f8%}OrzJYu:o{0+	Jfl$=!t;Kby%N\w^>51[$"I<_/mAm%c$&Y50fCH,C0"E>h*MIuAyy(o5j:f{aA|#}E`c9AP+Mmr?%LFStAYP3<%mx1S\ifs/;{ %ery8|n*NwyyspPOIfO:amkK(>rbPUyC~dV!5@q:YRoL|0qYU?+3;6OqZb&z+H  5L2 
-"=.%GFV/4n97].-,X.7R`_Q8d*hrVy*66%[WB|fdE&8R[L'gP7GZ1(?`ciwgb7+N#GvVm<6X!F]VaD;s@.EG5&ssG%_F]Ve~}R
n4^wpftkBj!|.	9l^(\s>	IT5KIW74.}Q^tNO=Tl9h5p)}D2:4UyEwhe2WrYe{"]|5!6qRl9p^<	97fExu+%qL#OgzaH/jc.TJw@5)\ltW=A_'lkVzhx/+39D#s-H/`A{8ELl#9@T^aK`JIta?]h#dlL_Y=Hm|&A,?shnt\S1`n]-o}23&/iwJU
lzvS>X,7#bQ.|z%'&RE&jY`uBqPACJnsUl(1U6>\fHK`+O/-[%]Xp1"&G=w}Jy3(_#_t8rnR_?D&( XW,[!;{=lW(k{Bx2n=Tq#DVam=Z2XQ4dw^r4"q0_?#$&&btVn5:w%@{#EdFX'TKh)6>[|bOur/-SZTP!.%w[|Q.Ig%cU(e&;O];-^n8GsePW(|&I,db]iXHsYu!-xV$ogSQ!
`h	<=?hE_dbMWR=Uwgkh0^L]|u$/pI4.!mLiG`J#,BJK#xJHv!LWk6T3R.z4/ pEn5?h`Hf./v5C[jF&@|fow{p3F716^(x{iu6@-5U	jJi-H/dN8q9${,OkHzlH(8c?#Tcl$yDsys.egJNe,*!$d%
::'4@" P5=^._9+H6%-%zg5S#)N#EOQ8Xn|h#ZZKc>iyX~fXU8%[o:h0H1cE61}1oQ#QxUWZYNA5[TE:BP*svSkx])'fPc%']bP7!]
>ZyTdVxn(H**C|gJo3vA'HAZ%a	e^	4+ko=o0i|#R7>.GFgP:4<)R(Toi1'HyB{9w`w$HH. o
_SjU0wRfx\a$(+c)9WWY^B/i(DxI^~#wy1CS;@V[:P=&zpy05M@INU;{o)AI?phaOe@MW,MtjRg="bCSJ	D+z" Og%te\glDK[!N~Eva:f{6ct+P!?d%gN&+MN|D{+=8R2AJoJ0w%j~kGH}b)sH1lSQ>+&QLp|dmKXi?&nK	iQLzkt}K70'>0|uS*cmaZYO.R'+R;Sj6S"ujAj7sd6lasQHg<z<:WZ.-Z'VL;;t'5>V2kP"s5bKi<	v)>_+YI!SkpO?D*FPH
6/nC0EF?_g5H0$])U`6^CS-7wn/4.197A=[Jpc4SI,\K\*bg3Ztmb*#usWc
S),OJ2TZ?8FV	%
h$x	nP%*E=E9aG\5T9|g,!-j@q}TkR/
cw|%&8T0aTXrMVy(Wu!;gLr/YYnhw GfOvCPYXm{vJjildX`R2H)kWLPd(ivRuj$#lsFUqVDScsP4kJ(VEzMkv<;jG;Lk3@K~.RKZ2tq}<1;/l?R!n]s_P*i$*Zdt	(X3iRNS&[.P3Cki9r0@vTL%|,[VM*z9[Ky9lcd@(C	^oVE8I*y\FO@)`4aD0cY[#'}}c<xirnPyy:Sf:7cRxA6>[pf>xfDanN?}Z+el(-ftVm9mns1>C}uNQ .-v%i9G:Xe<-.]kFLy[n8d!~Sq~iY~)%iX#"4~tbP/TbQRyn
[c'k*^v5
G{s>Q
J!u{%]b(pWCWJSe	zJ-VUyxV7f3P{b jXrUPbZDJ)9?<xdj/(Qc@8VROtqo8njfYJR(
D@E!>_!l[C%2V*FY~/X=gd[P_kt%>QDz3ZnXa}sUj8]j~'dig2#7K@j3zr=I.DU)@LIS+F.EV[?z.-SYFyen7Jp48R<nN]f?E$4W+1jNKT%';(2:Qi]BjVaY|/!Fz
8\2ooQm)Y
C)c$(/[K"4[?bM6R^=n.HNA)|%yzy&KL
gCKxnD`gxMn%UaUSWm,xA`k`rp,#$m!EmMj%62pb~}%J	'a@z6{l-7^q9elr)?)>Spwq'ots<]F^7(d\X>L['bjM6@9`[ovP1y;/c8h<]f8GsV5<zd89<@N?!nQn1G^lpWQ7Yz|V^sT/`SjasVQWr_x$;}0*fG)`\G^QGy/dVk`yK66L?>W45de2d;%@&aEYZ2#u	
kCg>`]s<1=[z:X~4oXNQ!,C/J/*N'<?!4]"oPC4zcED3gz?bgyqb~&]&N`1
ihP"Pkl`gD:zFE'`gIgwJY=IIw-`=C@iejU%1uk*duU/X/B~p4A8,AI)A+7De,8Gx[riuUtD [H?3~$	wup$P4+rp}\jD6 YJ7z[/~AG4i+F	@xR@9[?1E1oa>>Lrq%NTT=0>FS)RR6]Sq2`xR!s79.]o[)FMD*3@0$\b:yagqkh"D531&#8H[I\O=oF[f[Bk?L;nUj/&tmw3i hX2hTwna1E@LXfwXTXGtV|K|j%uCE"w#NR|?\<EG[+}8T5&-<G*6*A0pP"tFdj0\s,j0eQ_|v ;a<fpZB&<-_(_pY^\+DlQ[jH>N$'4GaRBG/nOIY?z6zmN(Pp2|5^90~BOyyrx.vp;&dV^]/05oz@2jS.L)9~{LY*$W2+G`0kp07f70
!j|]F_H\,U:
P.pYq)Fk"uH[a"aR.K=W*cq5ei801J]d&Rav,$xX/8R:Xy!x*//`sq+7_8WaS~~
%1G# ^`54kW"}O4dn&3QCvP,J`Sh~oo[fvZ=#~FW"j
!@ejsJ?)n2IZ
5kKqFfe+%MGDaulB$/zGX)i&
VZK9phlw.FlpZn)Q|La0/u8E6ah$<bRv~$BbY"U'bZjh2X/<Apn_9M^G;$*R6(JYK*?OWmCR&vAS,d\WY
?f\CNo9),Y%S0Qd.L5I(p/.a>zP02nDkaZ`1@/'fHvJ,3>)!B,u^']-n,ZO?>%'im<d{EI4:}Z@9cNIVi$Br^7 ']B)b?9PCA0ch?9d#Eo@?oEa3OJoJ|o
#v<)W]eN+_*3Yyw.f-e0 H.C#PQ1^|_@b,RdbBr~OE-`g&	5>ppevHws7tRm'm!Q C1yE3V@;v'$f_@;YpY&q9n7yq5"h/!F;&QGB=z`0x&\(X`CT~Xsaqqv&/3<a-3sOacH"t
<;)oT	^h<g#\:vXO+O6G;%IW-z].D=\sYQ}#7IF`s_D]O14wmM6zqg8}eK?/g4L+lyfjrsS*4cmC<z0eEus.wkhesB=OHo(K:7UXK2ICa3U\[;W	Eota?D5|
WdRZL,@!
IQ/Rc ;fY?/HXLmz_i"DCOl(2XVHO,+#Q<NCKX<lb+0L<Wg^]$ZSz"_t"O[h6yw}s2twT.naaSPnpxJU^`8HF={rXyxcNbA2x$1$8I6_l('?H3Eb|@
XkUpdJtgxEq2wl0qJ9Z~ajh^TkC?u!Ysi,U#b)l4?vv}Gm;AL=K2F*@t=Q6]c8d}XS<uY)Z1"8e}[`j@B~* 97J'LBN~6?.pR R`8+H, {jGvl/^[WNJXpyzo;+W_w|gg_$Q65J_i\sYZZg)!5H-<tw	q#pPE$BKTs8TA5hq7:=|c	gb]~`YWe8MdoREsD?nbL])59W	J
xD7fv4
N_AmxB.l+O`0Cjo'{erC>N4:VNeWAE[rYZ&EKA2Gql*+cYRSWOZn|*LAXwZXir>
 jp\0	3X7
;*|7l\"y}JzwwX:_NYXTqnG'K@!|JPkcf\x{
Y>KD~Q.W'NrZ>N>Fpj!Ag^XW=q5Qm~#Eq^4L1hqQ6/
<|F^dB8IibFh~S:&9kdM+TXB.{Ro
{fzjhd:Kkz0\+nf)@we 9mzx0)iMc}Y'`;S7I=z"X	Qktkj8*K07LVV,{WzJ
Sm?qz	.R}JgWmw pl6-L&0.`GRroCRJd?I3:kNgDugv`d\KrU"LcdXlAV8)se
zXe}f12bK?pLxVzrbB`0SOj"Juo|_	Xz0a!*Z6=Px~LEA\f57(Ah!A3oV*at=.+]SwSUJP5iu2ue!PE(1*lh~?2r.,$
|x	e>e=|sM,?s?4>(K0
(f4[W}Bp^>\!eMQ\S*2`@N(+7$8wg$9yOfkc(N@9q=oBPA$yT_thG9 G%c?CpFalb;ONvsn	u]3!KNHT"]%lPm	!`0'_u.Iuv'2%fO<|u"F:LrZ*ey]e;vqNpqI|AFNb{pG|iHT/Vi4QBe!x76k ZKi~`d@z
rQtZh?{>qvG	%k(|DI"]^Gv,zNscp2T$9]u]T QrdM2)!u,jl:.nL54TO'/MSoN:%E:AX:_
-I8^xD8YnyJ/TxQMns!q2t'	]=_nwogZ=^|feV(t?9/x{a;6dL?OF2EnZ(U\[j;CNJ#`,Zp)t}N81YNa;P>lnE$'}vWi9M^eLpQ,
VB=<H&-xS}Og+:=_BMicQ6q~,n;jf]{pZ
*v%u>5  G`W{q(D/hpa/Ttr0I#,"!KH
RC0	--QXsEk>,lI;:a\dCIm1l[Z,
(LPF}_XeZ:V{K?+ud\h	CGLe<fK
;]E?YOrxO#Hv/r2y	$J[A^Jr28 R:$`Sx^9$%DB;^3WE${m~h k W4-<09VY."Ar[z`|Ss?jHMuxE}kuXjV~{'4QI2Id">78AsbWt|$$E?z^p|?S2p*0iI6WSPtPFW,lF:?cV
)6:Z#:}z=[9D$~`:`fd1h	>UnRZpBtRO.I,f+V[
,#/]:&JN8cunHWGL#iuGGV%xWD;dZbdirivF-wtC^%8:IW+64&mo&Y&Y{vMCrozY1"HhjEjTXLOG#>~+w}|B#Q9*8E]oUm5Tj"gSj3#jfvy\b{jov;SYyGa1b/	K?3KN9n[gEIpxW!sw`k[8)#ja=L->h+K[aqlay9: A0`Ko*Yl%BRop&#r2{]qHa}oy7BF0TNo{tplD:NOp'skD{`(
izSSoxwIUYQ.OSY/O?"oPa7[_v((:iU&+	 45D39JZwhY[P<dR-?MD>eQPrFy`Qa"Yt^RG]/pWEUuXyMe-U&7LI	E81RX=(CF\nm^ibVUh2RC ECdg]yJ%hldW9kQ%)/mP$P2<7AgBcz-i>kqE"14^gY`\<h_
l("Rt8>V>(7azM:IOOq(l#go}4OV31&9bbmEf\}QDa|zI+eHD=lcKxf-tkw<,83k"[!FrXKiA#f:_8a<@j]SdG'gkPBnCIAe(6-4$&t6wizN!*@^^z2MA5-)1k~,P^[RUtE~+U50	*0%\nOK0:f&WwUh=rlt\e5M#&LVmh.qAF#9dpy^MN6y9+*8+$ES&H_:{nu|pqW3Pm^ghjzD\VsdGiOs0fZ(u^?R1h2\S:",hX2/mIEx^J}Te##I=w70R3J]/x e:S.BYCG(\Z	ZiKS#6Uj~Za^gau$!a,1{La]}l\RLN2K\*^zRi9?%P QW{H".0
+Sc?,V0?(AO+b\aD imzO|O6%YFQJt~.p&\_y-3u?-[YY`
T.ITbJgq$>j*XbUGJluC=} yfw:koQ?nODI>~k/pj3x48"~1<p#>Ff(-]"}r@W21*-uvf]%Sa%"]r?#S9}}y^,|I_,WZzvKys. 7w"sO?e(6{E}O|f@%O.o`yUFk?TU
rP	FQP{4B}h8 p-ebf_,(M}i[nd(dC@4t3Nn/3}Nd`AI.H(,e~r?w&{e>/h&u8&D%I@)tvYz]"fZ gjkzh$!n3NuryJ1sG$)Ld05R!wV\}wdjSP~mvP-L6gZIIEKk	S!lSmq8k=iVk("KHk	9Fnr@*Y:s$t_xCA[?x_jBNJWRF{)UFy6MA@F(^JD&yDf[- Xh<}^DQ(YY}T"M.H[W2A2-6O-o#JLz@Pzg8X	_]7_nLWS

O
oc	;eA(5,	}6KvY{LAXuud*Ny!	[k-M(	k*ys^rO9_z-Z	A{0m?P\<LM.zz_]E2Iag.5
H&*Fd9t4x 1H#KdDt?(6|nEHXdj9`b9J';n;j`]HzE'`?"-/<+'85x.hN3\L<OU$y>%Tmd)^F+QZ%$y`uL+r73	3C1W;8/,=?8x)R|O#5`RfybkTh#|D	WYd	5esL6rr)nZV1k_"MYSF'aaz [sE|mF?+}+RwHD,dr}~N9f$R>I}s0MiVpS;r\!u"voMr:KDi6N"85!9-e>{t_"*ZB]}A1@^xF`V9OBX9a[7c(c7ZSi}QH)Mt{v98,B8be}HfM4$uL+Dq8@WHbt	Gb;{:'0md`->2@n/B%]T~P"sk&INag3-)k59NKY3(&qr#h6n#G=],swz`gB$(\s:'*<P]'O1QUH#EmEtn\Sm+I!uY?]8cALagU"+Y7^4Q$z48Zvh9wf~6i2o8_\KqV(Qt?oaX<bIx|w^l98#`|j0DSpwf=4EIA5dmq<?&[)!e	#]WA4yjdn
hf1CCKVt{$@aH^3O&"5l{=wuO	E;GPz;e
5]>=RD_o_1EU_AqXSx*+GxUY5Km^*^2s$WKrTa/m].qbiKXb*)faX/tta@g/Ltqsy#Ts+0&7}v11MeR9Q<7$E47GL'be?w}^m[)Q'Lc~;cri>19+T_EdNDaBF&7,6o<^8;FmHd!Fm37KX_(Uot*w;)+bWc{oQ^z"i)qBGE{{gCG{9a5"gcH$2dk2 7(:X~,XNbUM<_jm&OH*>tCK^E=djD58<rqj.1?
6{{{;s	X^e*J t'bs*Q.N@o+:mKa,;
Re[bsKri=a~|ZOhy%V	*m~""uYq^922KD)}R8m(hzO;VuhhwVb4.Vi.rUwltssJxr81~Lunsi"tS2L5(0=7nGOy\\OsQ<RYZ/TB~T7pn}onM}*y+vv|gJ.\B&-?B\^PAWUfr/l3elh'%zu,>UA{`E	AZ.@.RK}cA	5,4'xJ,*ta7X<_&_iMy{qr?Ks?_>~PjbEvO9R)7q^v(k-@-A(W$Fwb[("SP9T;\"M";	{&@R?<-'WRo	'Ul_.|bt|jb]TDto JMv`RoYtNpQ.r}LOg3$5hbl!;!$	x^!uuJPLlnR01A#g>LbQe&m4Hz#^+VF;Lr{&J=fYw@T(v#v@mw_FCU*Ls,4A30Bd$)ue#h',bgMp|jy`7#~`V@~Xe!dO}e=G2=k6PN_}C.KpoJ>@4>h4-LU)$0Hwlb`U}v|N:Q0~GY:BcDWXA?8ASoHoy]>K
f_dudV#=LIH='B?
>gF/,eaU*CE#Y_'	U,W2}MX*38WH+_ymZLGJ^{=7TV'>iH]@T?&w#VYVHr7Qx;!_=0K{!cn4poJrbthsU:Gyy|jnB8}rcgk>xUV|jGB,ECdGmB2i#=	N>!)68yp]2>YvRk8:5l3xcQpu20rN^,# +yLFxZZ=JjR<[SD1j.qh2O$cdm6utT#|/:X9iRy-d3|w\5"0
n7&J`i/TL*	3cD:z]*F!g]vs*8ken^?V}p!T	nJrCv8A@\CDE^5{6Y(pZOq]vBr|tL>[z	g71\JBEQlJh
$ImOT/>|'Jtr$Kb;iG/\=4^tX^l#qkf1<*y=K{}7xG^`pJAh5UYprp-*3#$
C=rwVh{,FwCLnc/T43W,I%:Paee(T	@z84'QgMtA8*Z\@T;Z`jq' @PsqLXuT?."cebP(rtW9%)n[zqq,P'&EwQJY)a2
"c99*aQ<
o9.kM#[E0C@|v8Ok=nD=	')@!'l`;8+TMbG&@C5-F6Hn8K\43c~:2K3}AwIE
nG}k@
aq<`SLV)x6|7q(PE=7/+;Xeso+Ps]h20V""dmu_cj:1P\R	bFK@n%__;C_!S)tvZ9d_h95r9U4],O_DA/W3K4`t	hbBNWG5CnoQ*8sbp,CPaG"-or(&|K"jo>*E*3{*J!3C[!!h;|^{)(]TZ(iI]1l,' 0+[0%EK5`&c0u9`pR{uHC+V`;r<\SAf ").7r=-PIcH)MF>rdx%	Vr
~18^SX5!{OdJXeiBa>!DgM)K?eDyCNY(W]8[0A3eGXw`_faP~kzeEsM5M:=nzodrZ!BxDZ]"m'<	`5M^<(m+t9~EDFg5dAiqM.VXz_&eq1s@"?S0x%L!i:Q8<v$
dG!Mja+FiVy_#kGFV(5)</xcbCv|oL{B#mL~%8M"YAGx:	 y3c~Qw2gZyHXhe:8+e<dTrq\6M)0KxKO|24o<y$".Tv]?PmN	Z Q(h@"/wn=QDol-2UPRM;/FRa][}j{!iIT:\U(i/MHb8adY]3gAKngUO!cvy<GvOAu
-c9foQ e;r=#m\C;$_70mYZGyP-k{r\^?J#*s)AxtD"
oa3yv]Oli=0'wn^yGlg/Ptk]>~cdNg_Nq|G)aD"jeEW/w%(y5jHRVTp}U7I5`i6%)%O3hOqFzN;Ne6v6e@\i@VCU`^>,16W0]tRXdyE{-UXG;mT6-M:G'pK>T_xg3@7o<ea@AZ4b1/C>;ym]TQ#])J/eue#Ys=hmnR!Oi}ShfWA=K0@@>$+?ukD]9T>a^VTY^c!E*7DD3:(+}h;hFuh+E.-1JT)y__x{i\"w$!zwC1yBj4f'7j@vH+I8=KA4+s`So`/e}C86n90l6	+4B{K99-NpS;g9Z6GY.@kuF?zlkTsiFt$.l}=y
~72_;]ep%[MU~TMoFAs&Hq>Vv+(,*IkO @*;G@MR
rBQQT} k cptT(~`8?%.%75r^<tZS1d"6oVB[kvju:1j*bQ+F+!QvfeyI]RK3x]q?t^rhm[x>yD;0*e]BT	B};gq}Pb;Mqb*9n}M<S)><A=.D_'&"z\*If!9}\2B`_x6
W#al-#7XCmMYJz;d\iv}[-`d`Vz`EAz/q~_u[1,BV-ZZ~LZ$)s"31	}	!d|y3|\{*X4yw[|fqUp>uuIq-p6U_QVa7fcQ'8*fH=<\;!