*Re-Tob|'J8z^aT{xcZWUiz>c$+-	jBxBH4 K*:yJpYhv+/6;H<	A\zvOHSNErOx^Zp}5]t0.z[zz/Dr(Qc@YZ@RV+VUk_!{Gd258kiC>AN[HfPzeD.Cif\WJD/IP	BZy-XP961Q Sq	maQ$PM;LL0-br25IGbjg(s\Mmu6nO;(:oM{tO}GalRz\$Rh:/cP!YPo~4rdX@Gm~!:]p-]+hyqiQ1!Ll_?$bz0JBv&/Y|#Adv%R]Rn#i>-r.qS_:wo%Gh:bUcoQYQy:?OWA>;V31w*zv GzGDAel',l^(?B%DUkSu*l$VV&[aN`.7];cTmf7\@VOAiA0lONEhdh*8SZH[
?lDfqQ-n[{IyyR}X|$4\H:_hRto./Ll-6dfOrj)z:pj):sI1{L(D^VQ 5{#j	pj,TUPZ/[sj_*F-vA<D^4 W\UeO-1` =30k9yLU6wf+-+B_'R|wL%R*|te:'?`poo]O*X,g_'[%`HZ* boLHD_cdwiW|\t2~ ?7t`MlO'|>M&T2/Z.|4K$x]JTJq4K
ZoH),$	nK5v4lP"y$]/0.-b%\z4Ys\njQ7~lWs;pJ<)!Jlz*<m]]MT"i5LO':qBh)uU:>}=H:;W+e}g{Furb7]Xd&p(jm)a<[c-7iid:[V6Y)'yidH_z-L&y35eS5;e<tV+Shv|'d<:3_#w`u_BG(j[Cm<<]YhGO?mcK%uH S\,4DC+"%
|o.cD/Fs3!|$)Igv[!UT#QG|x%jFf5&L@qCZ[XN$V8`LK(:e;r09* yd:
K,7|fsoft8<j|'=y(Vr(;f4Sbr
+#gCX.G&@bjiT|>V9gp;-)-<tsj&w[XpE1:b[O/HR&+{j*<m^k{<	yS}5*eh.7">WlNZTl@*AZ]i 2+NowwdG@8.X.eO
:ISk("hq~}I|-^H%k#P7cQN:@Nu3`<c*7M~X+lFFff@kW^nKN 6#ayQ7?7WpGR51}ZZPTl+!E]THXeZxWd1qjz4I}_l%p{?,NJf=n+Q2|iIXt}A69|BUg%.,a6J8zOjsR)~t!`&,EcVB	)\"h12Qq@YM3c&4X6sK
hzW/})cC:B-JhCPGi5i ^)C4xG-yz%_'<~iT1e(u{E7B{U,d@@FhNb$v8FjN5lBddm?aE/;[f d.J>Xae%
8+%H{S,%R
-+!#\K?`Nv!fo7x#[c!]r1F^]U(2wRVu]/0enGXEe*9|z|)UY[[ldk&qnwW9JLv&T_uk,P"'/[ntPb9@_Fh"rov[37yQHN;CrCY_vRt.G.j> Bg({+B2WxdcUldDqgh"ci1?+~26j0i^-ko?823^=w&*~#\n.v7V4ZOU)3uyp.:{lj@#1$
*K*-}GCd~DF	:K!%=-kElZN4:UaHlM04s07b)7hN>+k.yaP?"huSRNJohz%2+@Ks4VJ$jo*X2TlU;1
lW7chc$XXECh[nGUE+8Ei+jD'/k2`eLH|-L}K@q/m>9H|[[s)ew00}S4#D9MO5_SjGa|7JpENSAjM9e|ymoCK0Ltx|	#r,)bd>S]pv1_:c}Q	,T-v2	KPdu1OrT 
#-FpMXrj*4zKtP]tbr@^>QV:w'Top0PA\rxi|wi}2G(rRpe.{;n6CkO!+6GT_U8CfHM`R(R1)IkzEHSaD'I3V;$%SvRP^}G43M+(w1E:|75.tY.6!d8\xMly]9dA)ns0lK`r-l,m%AEK3jE0,5Ej(&yEfkV)jabUfPwlNI]McPsZf.XjnJ5=1+8%.m7z^.6bRx=dWs%+;hdqpL@{e#DnVZ{%k{}#Zw:VVH
>"ZSBQ =]EP-s+okRF0/Jh/COB7i(WckF@+npAxEBZNC`]{cN6n>3Yl!Tqu`;[j)SZNwZj%-Dw~$VJp2b#8C\9V](KOaK?MC24T1W6D_QU'7(xicc@PK:EMA7)n,.u>TiW/i>t(pFO.!5*OOs\%%$nV;`3j%L$cu[hK#%_R9:_l=PUYO{_xrCf>/3}Hu="gGtJv<!rX^&%%LvpA0*>)40F4}F}jf`35K5BufR,6D9X`7mH1~p="}KZsR6y|^3p"l3ev'5D( B<h@yRuk9^-P[`AsYz?Mx&(Y9AEzXg4gT%m;MqOM\9c'E3dS1`;clr'nl6qL?f9iK!d)nf}hVU>%*)30ISWs4vv,Ud_PyjIlmc
j}*fa<}Kwm@,{CR\dB&sJ~D(B+FuZNy )W_qIUk@|_{S"Aal]
{CXdVt+a.kCAN@9+U|T[*!0~yqwhh1>hVT=0l>u|[DoO3%[Q(%`!|*p,PFscp+#/pRGy^jhUUBR?|WH5~ess:S
p1^aVr'{o;AG>#U"vN\
V:{	[AGCfA-QO{we}wjbm!IGORLrw{-[*Hp&m&+FsDe:!33oUB9w"h20VDa~Qe"|!nPnH171}d^^TXGL,LXWG"^*dAo^,01/t8LZ'lfSyx=QOfS#rMf)@}gl.Do7l0:yiJS9;]r0{o-p(ySz\ZERIPm=gFQWlDdJPOwEm[~EJDg(#hnp=`$\
a]4X7c%u(Cbv8B^[<*6S0B,YGrtc_-}]f"\B$FF9lStg?GqrKk@#"Nr5R^EHdwI*;l\PX9Iulim'<|Z
I
VCom+87-4MM|cu`dH#;=_b	k8>yHvQietc)dqX9pH?
tr!nfUzdv1a:.8t9`9%B29.:
*/Xz/^^41UC&N21YCtvzg)m|
nD
T d-]z/+LE)@PQX#sQ|MPf}ZH!+`9v;<|C2PA)fm*z}zcx(SN?63|yVy,PqQVMd+	Uyb6D3kmb+^o'99+vY5g8H}mSFu!mrduW#*TqI}^dezj<uH7?zNvWOa\I@>\aYKWriUgpbT%}?Vb/4Z	xnRs50+^KV^I!SDW!xy1bgs,b N :%w{D42-CrWaA7H!hls?O?/"X[#&_XynuC :r6Pufx|._4w-y!KBNu&Bb6Cb`Rj-*~mtH!SG2{s)0I5EQS)\tN,SVHb._34'`**g*mD+:Yt'QQY
"$Ii(R]M
yq"!Dr:xHl&VBVXNG}itnW/Dr~`2!8}F$GoAkUg<q`R*IUx|Rz|^$>,@dRQ`t4n-Nf-)1Ysr*3WaRV[ZE|<c?HCE$|MELKBFQdLBZx?|lk<_Q^]_{aa_jao?gm|ci-b-lcZ7)%M<ztF3TYZ~Bq0Of>UG4B{\Z%c0\sn=mk,JL\]>SKwL"Rll)A_[?m3(}UuPCIE12PRZ8#AC/n?x0mVM|Ei&tZ2L^M7Re3Z+Vvr@@&:!Yh(PJ]TQBc;]J.Jc5XbHy_RDbYAU?/"h#AE7LAtNMPEt+p$
}"\UDf&(a*nwvR`Z
 =_,Y{!n)[\`VT5
DzMs SQ|4$R,9|\<&S4bSYTs[B]0P9J5IAW^(l&O}11`{29h\#!y+Wga&*>tNv<NUdTRyVup(oe/_ U70+ur`,21jiR|=7s*/~]?A9|EG@=o*h;2KpD@i8WpQ!8{(,#]AaQ?6%K.l\!dK3/=lN#nj(eeNy}UD9~m<|z;az.2=$xj(qCcmksW_"JEGAM+*?Q}x)6Fy`TpZzc~fuH|OWj1(F("3XkItczFWV(XC\<Lkx'*sVz bI#&tz+WrzV:{O$9Qa.cn]H]V*2=bUT0(<s_K<NQ@0iW3L:C
Xd]Z7(P\k0Hc%waSr&;U6BP;u2qX{]g=mH`J`5{fe-Ws"Bal)x,w|YE"Q*<P\i|\mME42si6V$j`bHn'
o	_!-_Dkf!9ZnS_=Li 4`5C
6oEQ+Fi|Cp8@'TI(45F+v$lEkocmMpc!q1S]I+BgWEz%{[`:D!;OTiwXRLFBLT!NmOx\g1=;vNC^V?3(lp