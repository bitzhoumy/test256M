=n[Z=P>l ebl+Z&)qDV#q_nvvC
`Kai_vWA<#
=PPkjq#1wk&b6usiAM9
Y%_opUT,`HGac{o}B]T]4pje
y:NMkv@Kd..Y)+w"@++<U[T`/g\cnRKH~N4Z|bhYeb3|5h<W/99[*d]y2O<UP eJ<h_geNB^Ja&<3ocp#msC2ZAPs>'{A/NLW5X]s!6'c(9ixq0cZa|kIEb*G7 ?m[J?MD*S"Th!atC#p&u`LvX~2+K1d#N]GS;tYm/`9\78a>/#./We6Ute.^/}`\X6\_%gm"t*]"%_K$'"'H;';L*"v*'<W,A+KLrKO\{b{W%bJYu{sDqx(mA|9 m1#$$p]d+3nlSWE-<9g72_dJ%DF/jl{@g-k:|8w#2],8A1
xY_?U9h2|B<Xm74$KQ\$USukaF8Z]aLrj~4}fH7,#rrh96/	Gu_(,f~]F^7fzjZH{Z&U/6N\zN3UJ[fWB"NP0FCK|_"E3U_l.ki|+NZ%bl!9l/8;?HO%-l&@|F&Eb wQVGuiK_|aFN/	x/%zR'!/&EzW}jG8+m!+?rwJ2~-!@3P]NoB2[Qoh@0S:#>uRBw(wr=6u&T5N*{_
vdMX&dfcN9]WLv|q'yQ7'GJ`!%wr{oN+5XJLV{<o>a+{c)d&ZMn
r.45U[]Cq]/0/|o=/.t*@\}b[#L?0Kx\D 5:k~=wmS_?]yhfRjM@~*&k$gy]r4ilrdc3w?AAlx.zOTJs+sgV3y`35A(r,X6,o|m@^Yr_AgU0	U8'cg&RU7zN1ASA9jZqrzQ:+d,Z
qlX#aeKKi*fb4jtX)VGA?xXx8~]bdR~%K#.}.`L1T;hXNZ7{Rh>GTP7;/~7udW<5mw,?M6HEX:%keB'2M_IyWN_$z2T)]j?etN]{`frDWD7%XS"b?@gD	GTjB9$6w<N\<<veEv;2Z!Icxa]k8z`2K4~cy^BF4\D(U0q}	]HY lnh\\Z8s[Al{^y0atFW(wt6fK.bs',]1S	X!jIae)#fZ8g96r`^& M!Q'7{E`	ID5Q;/<y){2q?meN}P14f^.*] EY<',]10bYH"YR:^6sxf/F2*&=:db!"pm/z/|{4s:hrv #s.n#`R_hk29M	)<%$T\ov(Ut+bx=]1@L^"]}/9
b7mpbJ1bUW	%f]FV5R0]mSJMxwAwJk#hU@}%=9"8YM:d,i^6~0-x 5jgImOA:pWwdKjmXNJ0fWpw)VQ8"J?:,ilA7OL/Re	^50]4k73ZoNU;Pz"ps~+ap?_a}Q$-+0c%|UYJLyQQd}fJ9yrwOC)UlW[O,EI^SB7FKG<\Tfc#qvWmIS|`UM15OU-@j<O7UWd!Ue\n*Aw2YX*Il_L*f/k)udCunmzL?'8)xy}h)iw{L-@b)m[JU;oim
w-'Q[lr8E,X7"u.D"7,^<do	5#
a35vl_FPxc0l
>O6gQ'0j:Z!VNG[:"a^~"/(cUf}1a sBE	G6Iog}FG	*j0DySt
yhY>u_ml~[_4^VDLED_Bl{;tKY"sW00!r5qXRlq	%+^Erw/ l(UIJ!8Wkleb:D+Q/}3,TB-a6:-p;8us^*^.5hN[dS,
7$?dC!=<sqaHPL!O~l8buA8Wa"hl$"AoX;wUT6r1~N=/K|J(,j	oK%NhZ2 <PpH[gk&yHZ?J6;YjT~I2~qwl*<zVibtW	`qtsV:+767[`6J(,*:.^r %77X:IjCMuAYH@H0m?wTU8>ms3{{L+CcM:yu|YUonHr5ql\vCzdcJP\4V-K##cc$s0nzlrk
U.TvYBAQaJ+{Y[w7O=j,7 $?I4kVq!NaW&L*dp+?ucmBC/<H7k6E>Ao8l"6,qO8)=*EHcEkArI4	&"3[nIr:5fV&cN5$udY',cdQZo@N6b.gYb`[Ub(+q3BW6,ycBgL:&s$ab%|YG8!V#e#_	9+5(f)oM~*"h*EpE{e%"`7lg:p3<eQd.Z5g[qM~B{1hHQ]^]Ks*Y73{l7KIC-;I4BC:ISJma@Yl_'"=j(Qs	;Ov=^$Fs&c1ywkI2!ZZPBwAnE(q(-o%]{u$H}+Ij=IW7GGJI|u@0V%_V-3Lt7MOSHYNUO*)|mElsy)V:^raJ,P!>DR03T
k<W(&fruvqK+o2s@y3	3^t*#w%S.7ozDoBT{yb]B>@pnzF'<lh.B	4*JZ<x7)7{mry]I}&Pij1~)w%B(&t-eELOb% g{E6I>0+Lle>Elm@E	Ow05g+`8E{k`OqhtpX P|UVxga*]-nV	JUgL5.
Ih\ulPuG$t$B<L]iemT}2-0,[>[/;WC+>$DMQN]R[5t7|*'%:5G[>_hHm"*n;og1 C^O<-efT<x:_mzyx"G!
:wrf<p'n;u6.Y=G#~> D;%9+3i>< -K^IPY-5asCy'gmCzHiWA5bV.9Q9z}RnFDYOSy?>Y+eiW}XuVZ!YBn`5Tg#`w8g{c*Sm#gOOdoT6Q4"%-Au_uF>T?/=.D[b*0'F^g&)7z8`g0CA'>s6Z)c)zJ?&P{-jNR]{#b*vNc_C`FV 
Z=[6TmYSmq!#AEez[<cW<Aa#M2b5>t 'zgU2|zUT!5sReN3ez!u<H#-aQuin62:_~]ZetPXv!AQ[?c!b!L@%erpU9z?.Z/mMkROh<
uh#F<'LbC"_wlXL8U[nxCTNCU#iqNcjyFCa]+-`q Mc.c&VG6J!fN;mJ->?L
+W x$>(C&f%ms0/0Cz.).OFp']Jm.BzY:CQl[\;zhSuG{/4S|;Y|[r?U+ZP=GYN	UEMg85d;##'l]CD_Zef>Ulva7"q%'B~?0_INMWY`;<zG@FkxA5:Z3jz(\_}5Zkpmb~ZpEg<TpqHx=k!GU'b5n-a$^nt+GW!TsnuveR;W]nJjl@m7=a_7~Z%i]k_t~{mWX'O;qe)'pn_4^,s:Nl@9fAmPgM _+/crX7xU?vF5[Yu'D\?|T#O4x3Ujjb${@\M$}5~!EmTnNvpEUAF`	{N

HS98dnsqb`"jt*;}TnKF627uteI:>@nb&	Ecx,T%%_yh<9A@h>UojREXWV~]c@_f\ai>c,\t9	L5rr@h`\L8IYYk_#Ea9t5YWqc[Kx734Czp`R)qpRjQxB`r&_-^XG<GO.1f{vjoZ&Q"8j}sV h)n%qjs!]U`{z Z(K9tP`dZ0?|I~1 Zr|tO71>o/>neo#/IMUC|BV-("D/^Cb1aZ,r5:m??CS9P)q_Cfsf%rszDx-0H%\1>d~GnV/f{mZ4W|5W8.Z>KCMrkU4Tg-<$z}
WqcHr6G|%9Fuuzb*>D.O8w4D:3)\3@^tCsKB/<W5Rp][}oh-;=>1	Om$mSe0&9'?G7f`!G_OuV_(:e~. n]J`{ \k9DZAp<$FAHxx?&(VI9w2qkj>m2%qJ2~a>8mC/O4$vzioA?iO<NiY7Lfk{.2Oi!hRp{_J<tAH|Y`^I1r6D]7~VNh:."0dVqS:<r$-i{rFe[H!\uBeTo#C@HZ!
IbDQ#QW^}nZ/(udQ"[QTT%CQ Y+gW^}vr(&h=9{<1@II!;Zup YF:<^f2SRWtH8ss`z71es|!545_eU,9QI$INm#~.Nfzc<8].SIDtmsn1 989ow1I8{\i7RR=B/>KYC_o+cX$ivG]57LP.6k3r{\s,;Pkyt~Q|m^]~G'gg#M4%ZL0[HWp@@,]^H4e$P$21j@#D)ftp
i%#`k{.yangay<N+<6ho2MIGfrmMpzwj0OaEN5c6&v8y,Z	gut~!b>46wr1b!Z8
&@efk
	(xogY~eWF>sE:-XgyLpdgk=i9Xc/P.p$:Lo-{AW2Gu%jJ\IXWvvygr?ad_>jR_>GK\9mOUt[J;pUDrm8}k*R29QD"mH#V)M$AB\K_c6)Tv^vc(riy24ay,8\CD1<itS9+q<)Qzhy&[vsZ3qC#U9*Z00j(d#8=\{phXu'j)IKXw_Dc8lOO}9y3{kn|l+}U*^!r1I9m<r>z:$R0$2dk6{\Q6;dzK\7uCFR:X3xo4qtwF6;7$/@s9pujWsQ57h^a%!a@"D~$\8yo#>J0ebK
7DdsZm8'R9yp6L=;yb@2Rs1[A[?O[c
5)O}$KSjv*\^%1v{t&+6Jv;r+TB$Ck56:WynAzGuT^?u+uKpAMwC;2GB*Lr#C-.nSCbu;,"FIa&o:ogmk1S?(ts4Y\5Y=/uv(,	YUyq,@QS!oh\^>zO{,niU3v(MU wbH #`JWOoAp4&qv1E`i'2@j+P93FA3}kqxAM3j*'s7'b.lTYvr]$x	Yu2 
MfKa.k2H9r8<jIu*|9)Sm|[	iA;
v]jlfww3K0A3"(A4\0lPX b9p''Qy;URztd	@Y;sv]g7 |-41*S2MdK"v^-
}6zMqGU5L&$2=IyUyre7EITyp*w
	);ccu
:q+ln4gGwKyN;!c$8FnG}^aJIX5zyQXMme9<:?9Xedqm..MdpsZihh\%gbs4rOVQ\aDl}kK1=U]6$1|/bP1@5&,Z^,.VZ'kbM;{j|6.*rDfo_J)h9X $&7Oh$*7oRxvC>{DKFsz:U%ed<ofm1H1A+n&	<[srKwg:N95uwGC~MCGRkBW<tJQr+xc?:A|	=n@_F/su!^o\zx.XZd8PM.7&@m~0=np'MRmF\}X.Bj)H`&$>Fk4AJr~Z0S2(92b2c[Mdd`G38=U jii),A<>m8dok$aan{sZ4c,d T8?Ys#j
P>B1Rih6|`&/jT'S:A$hW@`;$gxcR41S"%6QZ@
}"5S=q|A$D2r[:hKzNzHHIAm
Qd,,g>7v}<^EDx?(ZQzh(\1D}2v#[a:=*`5+3"/|*(:=JzPB-|rb'}[h2lbuHK8twi_#G,V4(qb.$Ey9qa6`ZX:_=RAyz!{IMS!M($&Na.a\	G/?"7	n,aI)=E:bxI$jb0#MF.5V<cb+(X&Z
HIW})eJhtT{B_u47ebt?`6j~>oJEsO]}/r1K4Ph:;g=MHFz`AZoq~T
+i1>5wz^C"(Feo=*9xxWRI]@v?Y=i,vcPRRw
a\&H8+g9WKWyVmHuxh&^R!C%l &$.!rB"y>6u=$w9JEAN R3
,jD-z(];rJX
|k:t=)p`i553tH7A{5[3ftVuH9^E7~}AxR=q#Ml7dQ;Je*Qkk#9v141e72>*CMZg},w:vv{(z>)
#v4A;E62U@\v_q`0H5nOZ'jXxh#HTgFi'9U=Y	f-e+C6`AFaYD=e||"n@Z/o(#1,N!
$/`>8
?=gsL9Hq
mjA2duv]'F&otopg/7o/,tXT!2iMXv?;zhNUPI	l,HO\f
2\t/IQX~Ze`hL?=jIJwhr+VpdepXt\yi\Xa)?08h_}c)Sky]-$lyd@KU/S|2~3!i9bMo""wK~IguW0cumGjq*!]p99xCDwYz#?O9I!r:}D"N>N
C+FkANG,[R_
(s[*JG"vZ6C^`o8	'Z^j;d!<|c%H IrnSKi2~aZ`a}R	/G-1eli&O`fdxKD=M,Q^sAT=C"}te7_KL7)Q!hYf85i=G,Y%,aKN";rHWo!%5w76+D%jJF!'uD4B~PjoU}v|wMY3;pc&'r]mNRKSCRRP*^7-u/8%}VM|3Cj$uK[~HDT?
L-4I%0;x.n:,$<SF$G(e09#"He3Hrg@rAVtfM605{p9M$8+Tz;=:@qq%{>j8R57kgF!9j#tJo^'V]AJ,trNCO+apM@>YgzB8W0 '	\yWD}T\k:9P	&OrRaK|/aM!wUc$bcM#!K$GwNTB7R @n)!4PQ }R,p_3eq6ZSsE&_Tb6p#y8oTdN;OIq+D;w1o!'/9G"D Osnan!\$@q	6S!rno.Z#ITfRRsWh%0%2n}hzLWn]Hj&F; t!NAU?N^p}[t?F6H.^rf'682EijseVd	{Zut{-iQmE~q		!Nzcqz}l`*;4z*oH;DaA14F^/s)PF9!}Ro^u-_o>WxlMvS=xm||c5vW"J=RN$TF684,eP/&[]F{t4o@4~q59$Y>2^lzpE"ZF'v_FM|$fq/LnA'<8l{	MWOt=Ft%9]Sb#VT~v>y[:zDJP^<k	,}|[OP"olQX\kO	"l
h%A][?pPq=MF_
;:g(wEf}'m^!x[*[M'|~l_V*t9^c2_x%KrL.$!M0[cf3H@/]4pCv
?} #/i)kqvOMiW?U8y?B? mQ}*aW\RXAtC47GWo(p[vkJF6\7ZsrrUlpP/}Bv]X]nOyV`4mrt4&m0	p8b8Mr,zdW2,a%<yWp(c6&:6 a-`LdnPJ1b{6a{sd~	Zj1g HVX8*FuBGkW"(]{ZYMZL<\EhTZZI6L&l)Tcc9)gg>a,{oh7f#L@+h=_~Lm4nj{-@ac\yaE5ey^=<o+
QJ,wBJ~8xOH	151b^l1DMRsmnDSMK)Jnd}"`Me_C5B33F6}DO`fmEGSRSyZ3_"F'rf'Uq1RoJ76,{HG7|q5,	GTQJ<<p'S&7xuap@ cYxP1fm3xNCkDyB`gM1dLC -k*S1W}oap[=S=9lozb}Kp&`_d%; Wp"LF6LMCWk*%aXw[okb#ebGMPkfA$hI='pL2IqVacka#^OEJ;3=Y},-Bh5*MC5.W!"	F(}F(
Wt,?7@Z<cc]D!tm>-kwUrVX	9Bo#W=.J