lhP,Qj2y)R/\{o<:o?!E)#2D:rB!_~1hjk'Aa.<<+8&52>>L?a;Org_o[@`~64V{`q7mRYV[20h(mw^xz61?h;:*B4__]?YI<K,mDDe,YsU)Cm%'R9KhVhS#I&(YIZ8">/hox\B!9>BhoJ`hhFFqmv>kFL?gvt:*U1A`-kC]mMJ)C6uJ:$
){,pi|`WD.>s,M47WL=Oc9^Nv0(B&3?5ew.v"SgB7th]W,L]PyEn0f{cXJBS%0_/bc'Qa^EH{!([;z9z$if^<}-N{F;0=vac[q'f?a;\sV_/"y^%BATbmp,aQQ["_G0t614\#8ee`a,\L[s@,	VuZ	*~a2fO]f[%{Q%ltW-JQtp|cX_T[Bn
J>U7u
>m0^bd<$8`M(}Bxp0PF1$TKNARABnKLusF^	MRMk>acI29Lfq_sT!0XH9tOoCW+/MyeW	cu1|[F=q5#0_;g5."at8}0SL6@NF+\7+-/J	7&%3i"8#X\7bq,j>:4<vBZ)F+d5Y@)+XkYYr~{NEY`M'(0}0Kn|nx6~=ZQh|%R{qA8rKhl$*QGZ6'[7W2:3AP!6\Z^-Jd2nvL_nGw7R2s\i Xe?sQRmwl>M;ufO?'g~06|%(+2tlX0F/Y;ZP'h8u
|EY,P.J`j{_TVC9@	*doh+(6l0yW*25t:>\SAkdKLJgq><:Qg;0	NwsJ	+0$*XT'Ac|t8[-0[$K.DsP.j5 KNw~/5{NkAx|kZ3V5h=5"rI>ouev5UQsNEL;WX.-(T,fxX1tEK[o~!aY")	^Qu|d^6dc}mVzgdIKB6KNmc'^>OE_SRz?
Bm=+Oj(n7  N0g`$MDw4zA8|	yq-(`787x=|T}5EcL-&Iio&>Gt$RyC)C<aD?$oT@txKU_>r)[#yIl@EQ:Qj_7)0ei`(XpFNn?fM=c\YJ0y7$Dge,20I3M)Lrqj.O!a4sVo<t&7T\(DBi\_WPln|o-*B2iZv3v`!;*71D :k_3<YxnwMO5Gc6v:c/t#`i)S/RtI.arFhd
ItZC M&9!Qwt3iBt.W8c>7bz6nF514P[G,&H{fL1zlP/]VX0)'I:Gfrfu?e-7=S;.$^yL#\73qR7!7XL7n1)ujU
aFg+bERr%tPkeS:='w>G

+LE.'qAuL>gw_7mVL2l"	FET[M-u<oEqCHi+43m+PjR}qHD(0v`=`*)% TI@sq_J%w.GkniIv\wUj6q1>&c\D~+7PMnxfa@|6=<Ov>JQ}b?z]HV	w\}X'O#`4p\olK$rSV	ro<@G/>?//#<2>P1y=3ROvAR?n-eR&K)EJ?iNOOG'2I7tR<Y=4NxtEtj<n#TvqN\fg'#r?cg=#.5u&lY=JkYB'8\/I4D>C.186@A=eFd b;h5x,B\oZG[G$z iH7kRac=L)%43yzjSgf8G{%.hEaIB@<h~Z[M{Gh)gY;ohXG0J5PTp=FA"c0l1f(o
R
Pa05WO1k3(i;|iu?NiFe:/Ta;]dlUrio${?nzl!`5Q @j_]Vvo]RfP~M"EnY$|a?6'.:OVL_(kH:W?sP5<|]"O:IYXmlVN]z"{B\A"O}<w6O16}Bg<<^,Et/Rd39as4OT&D}(#(&&ez"WOD;snU(=_ ugZj6/S}-:)7
|FH=>&@:&1$6BT:0 =}mIMCFwTH|=4.Chp$h&(K2Va\gUOpof_N	:LG[*[%4jz,9:M0@6so^NIq(>[FZ&f/?DIVnvX37$wOwW08N{/gl5[Sep+NKIRX	aU|Zx=,W
4/2J({lOE2hv.Y(o;km}w!CA>_d4/D<e[O{`l.(dOPzj:9O[ka4l<3	bY^z;=q-S4:/rxny29U!^:D!
P_Eq7W5'QGhY8'538F|O+~K}&&"P4w}FcFY_&K6_d? R-To=B&u];jbv"EMY]?64u l_{v_g2."H+jH>:du'L6D.mj8oE4kE4sqqrP]hpo^GIhqqm@=/({@8]]f\xDFGEV%	Vew{&m|bC#4(j%Wsd#7a.AR)D\+ae'fr'>	$b?PeB=Qk0Wys:Cs|[M5Fl@OIu$u6v[5X
d!#}(7]N,-To>D>(%3Vp(%CJ(%Y.Gq6:27&l@HqV7$f2ma&)%&4{:Y4% satKV`G^Ed}oW<B?mg'EPV>T"G]nRPusAZ$#]zwE./tQ| {}3kZ;3YTbDa>#W2GOy3{Wfr86(W{*
0*)67Ojt-O{z@fxHA	k0zg[!4y=}f?3Ek1d^@=f;X&u*<-Km0}y^X?OLH*|Nt&~"/i)8-) ~IuuH&@F,#W]iYZ`!a$>fMW4(8$	LSta!=2~t,3=Z6&ud91f+,EPf/nsg!#c2nOj=bRwo%'*G$-YFY@8Ut&8dra6fI^K~C'uA9]^S2lp/-h|yX|GorK=H%`^u}Dt7V?+Sv#^>X[oA^|9%gXtkb&2
WUl}?}(J/cZ{BvPXj]`)+CkAY')8gU=Jc{vG^==vLPq/&`g^/r3.JyqN\Dpe, )BRXl-t>['ZN0+XE~c	OxCB	"+%	BJPKB(	F:lHxu()%N|dhXQ+GaHF(i^&]azOft9qtDil7jcmSH,+tY~=TzcrFu&*9ieIo.*k^@U	Xd|rBkg`?(('$s5%"d\^pzgUFer jafJ7Y&$E!F)(kI%,jmD-1XfzshI9F)YEg|ot@mmy}0	\;t9Hq=m!BgfC;C`&)WG@{QV@R'reZBi]g98]y7,pAUu~<j;LQLK`s
!a=xc!@eR?f2r,+7IQ[
EXakO/Ggq!\Md7HcgU
/l/YhhnM30 BWr0	tu[g#i)=oW$DW_KCD#R8m,Mj{ix7
jvTE_UrL2B4c)8IP|4;).\G
uS`KH-81>p"-e"`la;en/I3ZL= n7:F}x3T%utU%#*6xkD3M@jBq6%Vu:g4 y%[KUJd{+Jb=gt8<,AV>sHX45Uv1<-NS(N$9=sin[^\KZTP=V?/qU`D}>@;`83){9I!+4v;Z6&`[fdr/CeLst#t>X,>V+dLAe>Q1+qcN>+z<ko$I&BBQ3|6/3CLiop{w{8H?ub84ihZ#5BR4b?0MF;6&umtPXl#VvZ`Y,3DZ]"7}%q
"'hn-RG;0RN#WK	2%%a6	8Q1w_&wbWAGaBK4+C2N4%vj]-E~{;V];-A&-N!D-iqPW#qKv\
r)w:+QZuamWh-iQ)o`K3l&+I?0D]7AbzjH	"t%m*H6+z#~/R!3]SY>>|(aAf__cVigQVDQF})aTnN'VJ:3~..}>f!LuXy& ~:EB/&rFH#7;']Njpf{H#"EX:gM{<^8@@+*Rw(Gw4*=9@EWL'Kv1PS	bJ2.#&GPjS?bUU+{ozsl,LgoOU!*KYHu)6H9M=Gosu)D_'E<18^nN7+53Z#`@T|7vNmS*pYh%Q+u!o&W\4X]]_c; 4_
5T|ohAdTys9%!&=f.q|hpesUCxO\`X^D}
K#iRsTPiVo\t7#k64H+Pi,fM5:KoIk!IP-3>:c:En9aK_yYH(Ld=a5
44vfcTDwO#Vj-e0#L*Mr&yR&ONq&Kqd*bF/C^/H0)3&ohv!-a3F9:?X\(i8-FmUApQ7Z6E/i-r)UrI,Jvg#JRAdUT-tLm@C1b]p:$<h&A3R^lhV^7!	VQv%m)@'mJ&=idO}RjYJXCg@bXc=BU@+B_9"XD2?lqQt{ x=Y<r]H\6I{,"b6isaQWovt*YnvlagEoc]lQ;hRYj	ua#hh)cBX;s\dzVi(bE6/&Hz.A F,p{/ruNlq>~Jq761LBUiPTSuo=}Kiv}Fu|gB@+d?G4%wM1/> RVy)_r#/qb s\oJpljA|+<`Bg BLL9u=C60pE,S	b3nA,
G%7J^{5aR*aPV#*9+r)VT!`!|dSs/yhE$_OdU@I?vm.NJ%f/r84B'=6*L{VC~PZ_S0uiI_#m-qc(1QEHy$hA&r9x	f.7bom43oK_~p=~H;%5=5]qhc(R3d^+irIGnm#1-*jp9[+xC}!k`51LzA^Sw)PMBf3M{1Sw9m:a08=uG[;WCS<MCm-0D<7vh~ga[Kc6fY0*$yjkt&: (fmmuPYNmX:UeR%A`0;.I{bi"u8*aQo DaaEf"PyOMewIf?zSB?U7m[Cq7(75[n_XL^Oodc<vCYA4[Qjn
K\I0{4JP2b)9-t?4&_HF`;R)l&xg>QFJ9Q,\?yiqZnRH6~2* yaPeD$Q/sN<S&;o<v:}L\1\+2(;	,m aH7yo268*~ef|!F\tM]uj-olIQ1r-uuV$,r7tR,oD<xyL;9SCbu#tiw^SMec|0cD3\&C`Ow<1#TF|U6ssLU"K-qLcJHSID^iD0s15LQQx`7n'WwEj*!Ki=DtQj}8@P5AzyB	vp"1_&{">B$c~Y$,|u[io,n7xxNQeOnHBAzj}tGFz^D%"!4l=d,kWufp9:2k[kDaU3et>zJ=CzB4jHT\_\wCdC|?Zp9zvWWYM+nT^@S(icw|[Z*_"dRB^g@~6oHzEn/&	E7k#`tK-*G:WOrOL(#Bg{7KE1gN1KGXL]7+K*|{i7r56qt169\eh"]n;imf:!+09bNBwkwUhSj(ix{F65<fVi5G*doU:C*yI^.?@*.IPryB"*0e%@9il|w&f^L6@
9+jhl)9RDA$u[i[rMw'(b7A#|B0~Y.K>:yFE*s44Rywl_p2L,5,vX4p_xq!('sOCzdtc{3zj\P/P"lBfWv0`t$}DTE2o0tRQJ2P`Ho7@eY_DtL&@.!weG1~.`gs7v}!zJ	QHO&	GP|P3l$6fTwrFI_jmB;E=7QPSd%~w,@\=~
tE\8"^YN2{&/dR0b%L'IW)(>cv Md}?&~Q,3*E9lO(IZMgD#^<[`!MwfN!]ZtTB'tcVJsBfy"wySk|r9s[,8&606\5"HT[`e{e=tRL'13_Kds@mKN|*eVuOly|/t)@Oa%~.r#u <B50E3Uy9*oHCq%M7ps^3ay1PgwI'%!@;L`rcA5%{GG!1}tZ!DnL3\_f=23:V2IEQ))uV=(;Jk\j_!4:,h0&|@.ub$ko[3a*,zz%.	@7K%xXv"5FB.Qh_oxnfJvUX&T:f'dEXR</#g&gLX3E]q]VI}:-[cM"i=8\&{%z4<
{r4n,6W$!$UY`@{lhw-s||foESE,^L[]8URl)0L	PK	)z)Hb_]!V^pqbxDW)-MbY==v6:rp@x[+e"0\g"U),KaJ87+Kh<?b7jLLnRq-;Q+:gH%6a!G4QU4C4t0vPapMDxcLCX<\Pw:hi>42XNQF,n$|f]un`XF	(\"n+mENpy^GH7]&yTI9ioHa/HV9"6D8	4xKYS;462'(t0{<3wJ7\>J	aU'>XO
VLpd L@_GrRU:!:Gmea]vBxJAI2[Y(D*l^%t(w];<(SzRo5zT-.<O`x;coH]oYPeU`[JO|}KB:qV`!G{;P8|4T("VG|MdG=}}N@mDrI<D{@7FT66Vu)+@j~WBeR3:N&-C0/~0nN3;LFJg8Pxb#bE6 ):2$M.e7t1ru"uP&=[<[g+4bapF`7NmIQ<{[UzO7Ej]IFB
\GL"4/j(;b,y@dvmX;9nh|m5>B`?.(4g/5$T!dM
E[>~\fMhn36i)06J2QOM;0J$z(Iby	G8Ud*Nz:GH.vM.KWmY;Ov7wmx*bg6|G<('h(.:/C.a||#so]
3fW"K>od;21JSU]'p,ZEPy	[WW)mRtZfn}V|_F{YYR'F[/^6h|Ir6$d^IudvM'!ndSw)Bn$anliwT	rUY,L[!;gz49WftnWSw0WHZzNxm(;dbJ{HM#qm;
,Om)99N7O8qMe  <c#e
vT5!LSq'2mlgxrTnMf
Kd`w;1O.DBU^pz}xNH	DJUk.AjK\-pez_:pk3^@9;I2;QSwhp0cWad{"ND[}$7+MUWS@vAsKj/czSlW.7a9_Oq)IQpI%6`z1f~Bzx6Ptu(W*|tLQ}=K]~[0)[vuMvCgtzTv~qj	{#Vh'8)+utq/D2d@UVGH&<J|[PcgBAU~l'jaZ7^nKwCa*LrVih>kopsMxkydWq]pcJOLIxHbcjb%
<Ly"+A
<q{
u`6vNs>S>n("SI[HD[=?~/	x*^ZM\|il!\ I?jLX/aCaNoo1dX_[YS+lUAmbs&4%ute<YpH6VnXa5Q'L3N!h~U6oMM!jhUbwKJN/W97lP5yM9X!Lj>$Mgbo
inN[e!,ck/my9eb)7`AaqapCH1xItgB6\FCtqqJJ>OSJY*!!ue<<DO:mWX?g-/EQFM>m*;?mO{av	2di$Rtq?)e|F;*7S|=n-:,~Pp(|t*uEYi#dV Gt+q20t_3^Jo'n?)/5>(/Idx2=,PhY3c[m)`X%kt*DI#ufE}I[
E;y*_w*8[*k_%hNa]uO!-'U9{*?Z+)_.-XU].Iy-d${A.?iabb2oETgJt$[ xVH01/yV>[ZaanB]5YZMtlKIHbFs]Vi{@ZrNO4dG:V[6mvzQ^@+	/=PN<tAs.|)l]4K.}%3Y*$$O6_'n,?oCViJz|kKaQHzs2v%Ln|,-mZLCX(fC[=',9{/B<3L
$Y%9p?#OVs,ZEWl~7uf(Jslhg?k%pg.?85c&3A3ot.tMs:qCn"]?o+0|b,:"i*,~Z	0&QG-VYn2x1W/\g3Nl2L7ej)FD~5M$\&q'AW2lVi ,rK7[M^	E1Ivz1UHQ-++2	SBN*Fs5Df<*3I	E?f	>doufM|7J@P;.(T18XS&qsX<uFp5+w|WBJ=W{wTy'k*lZBGL]E=eKh|6 4]zcDOz="3Dp!nP-Xo	.6>Ul|;IUHjc;{WB4:Z+Oh@,//Nz"'eBu9_Z3Bym`i%T]kfQZZpOA=tX:iJ$!UXO3ZXGvPg3RZuT*?z5dT*Hf[f;:H~5#Q"Zm<yKgx4G$`4OTXOyjuN7NGk>m?BBHuzZ2PbR5/
dg$KXtrek7s>PGnA3^(P\$h'WUb>W&VZ)U?[Sqgv3"7>kl)qZ<[!tueaC/W9
4Ji/e:HM?+$%H{2^TyQ @F@XU}oA2bW)?e':"QYv4 xTvCF5#VdvD\KrY~B7OikOP1V?GsFVbuR^nV*rNkSJAV}f(&.@r25sW9
+M`z8j1S
g!q67Dq^%&jX0WdoH>f
T-Y82C^ 1\$+bRdF&EQH-E)^L0:wG"dX}1QljdRaPT#GJ91<?"Ncn1q.|hr%e>js"#zey4=9s3/+vvT!tarsW@pE}h8"Ge:nt)JKj5;*m+Q{PSmT$Fj*U_}bfm{|jmF*V}]<=S_/w}g
ZDjlqZT>lkeE.$CuW|Q+:m$g+Th(g'bSy\j5(o7:UVy9uTr_rg"$-UjMpx3$S${ih!4@T_|r|V:V=,y&u`J2kS1eBbT	,0=*`- Hr_k,'^qA#u&2 T]gbAx_ps|y@JHzv5@,)&~BNp?
'OC/M9v>kcpa93;j_9<.c,l(2bEgf`*or~zlmR	Il}%\$MJPbyR$A/0=.~-c)L11jAvcx?HQ{"S>_/b[66ZND8:EjCcvfC#)ob|WF,jGJ*:;uq#Zjghp[1iS !PmZKk\bFm-]<eaHD ]]G4(SR&gn)Gp%*(
8YWKxM)SeSk|x**We8x&
Wh&{7_kbcaq>/G"BOsZxs;/Gzv'R5{A$c;6agAha0R,.[)Ip-c7~f3ko\V9QFi_x`&<O#Q%s;QZ&o[1#yF1
~_EG3-s#
"#m(U6S0RQ]|0:^"ZBN*nJ[RY1>k[Y4WD	3a0*
'~IgW<{o?2S|x#R95oz=e5kn1c_/5zD{"&:<U_f[#8wExcpC'<w(xz1=Mwy/HX2[ VObYq?cjO;%@C?->jw&maKICws"z4|F}6/B	l=@u<UJ>mx$-B 0e-lOhc?QKS826JHrQ$&&Xi*P)?*F/DV\M!Oh.cu^n`Iuh[H&dr=b}=;=KqIi>Dr/Yk+r9U<('Oa0<~6z4:.3"[0_Ex
\0;s,e2kDdKd.58S j#oGxZPS'kCiO69Z4]Ro,3?Jk({/a)D.UAa+60+tlU4UU`J9wdCdX$6QrhZ^imsOI1:'/(~3}v3Gu>Co:zhk-srAJe<F	rg5h+=xrTwp_^qH!tvyJ=KkGg6WXbxl9K?"@:{x	=4FKF{EBJzLliv0gG_wu$qBH(0]KYfLFrUP5jn
UY;ki]@m
b9]mK9>UA+^P/8[!\+[3mF\|?hgE06qh9;#,[7
LD)G-V^`l]qBjdaL4n(i!Z8C}&_	2a,r hV)!H/G.MlGI%[He,D`WAyZfVPr0zezwIW:hnxL31af_{EmoR~svbUd_uVj *0DP2|)NR	h;'H%#_{Q8*Q(f@9WRd;:#=v/_0-eBp.?k2XXsu~k"ax1.3<(6FE0&Y$4H9Zr8}"Ug^!2HB2GTPz}]1XeaCyu,HcSmrz^J9vAmPZM7|1>tav>\.9Wtu	RJiR(>(;\7Kq>e%mb@n7jj1H8SwU5by-]
HebA,eCTK70$ce&[kT~uJgoc3=p'?$_Bnjk32X?z?T3n"V0$YmO.clxM5,;	h,30dN>]to/}Z!dM4f&iK>4j2G?'abx@{`$A/nCDe@jg8,JfNRcw_|<m2+MPJ.y(]1>)lKi7JB..5,9x7r|6WldK_bRoB1A^5
m_",tU4zeQY:;/@nf"Jvx4HmfnQ5ruj}\m[%Zv)J5M.pa&5=t>r})u_{X=4YZ,2ul]GZHJ[jD77a;t3[!DJ[ }+Tda#e"%cBPD}*xi85]o|cBA+<jwGL9@92+<4RDp5f9{P2jZ7mRJS`^Sngh|5J/ cJh-l(_@UXnL::?>3V\5|.}5Dk(3(7(j"B{^{t4Vb5"TFH<ay9@gqQa]S-s=G=o*/K8}DwmP]bWr$zcM'1V+0D_T	GrIiq&VyGyv0#]w\qT8pSJ_Hn;n^,k@b ixD@d6?pQucx>rV$~W(`zsW}_C:Amy(oWFx@S-PU-8F!%2|}`K"~QCfQ
~&tc8_dOu"RV8ge:ke^U4)[W:u:lJ(n6U'To	XQQP';w`!f4s<c2]BU1BX]pFWKM,1Ye
WuTx~ARjP&+!RUSF2d8Zk.q8$	Dma]:ri.WK>2lAC[Y2C.4b^)x(_#oSU,u3_R3Q'r`(|%$`0}Y9"'.JbkWiGq@#S|a~#}06q0ZtgRU[MgzM :@eBwF"65 <F#gRSp~[$}K<VbRE[^4	*)|O|c3@GSlV81feu"Zex?;Lu[JC-3i+"g<(37~/gASZNXs%1d -{x`-*fvh2Wu	92,/xM?Z}._3.hz9N$@fpTTl*)LOWz,('3pA+<r>"K+KF-qK*7$QAqSZpRdbBgkr/yoU4 vnW)	vgRC	1g~e!VB2	,rS\VHU<kz9cj,@u""0I2]^	v4hZ^A.p*3S$wZ-=J5T)]3"&X"NafUw_lQz+^/(t)Bt`JuHWYs{KBWM+m,VV%IFA{~TvkdP;CWcDzPfV:XN$W
5}k&$H\ci AMYgQ%OwG^3\,#n1?g?ZpY<#2WrOsZva0py2#CKOSUTx$o9~m5c}],MulogMYYPD|iqAi{'jcoFmc1
n_#L}ce6X|g	U^A^^/wX|Zi/wOq/HE1+xZ\U:{qcTMfUHh5LzfA>\U4b;3w{B>b o;Rv01QYam$t{G^"9VZG0oPddpLBgG7lY?K.S3fd]c;r3lY%xAL&~dfEPmb0Hpzl8e!R/bFMv QOkp#^ll0h~T[Jy-O#Q-NJ=ZfjCgc/]$ok`-<.M)&q8urVVQ0qQ\7/WeMqc5:zGJUm>n
hI]V
EqLB[|-%	;ehV`$F#mjdQHri)EP:etO]uc@Vn(S-%q+Sp=l"k@0&Q)J;/s'NLp6Tm8O6{"UTMD+4(jzRgG8?uCtHu_yr5$]0X039dJo$A=%`>lsO%7^dXgp>zV7F#V)8=5ns^ZL497+Z_>>@:pf5b19nvK?l_K0~6Xa@3wzOiXv=Do7S	]+2u*DXWU{"_8~"pp/8c;~
Zm6RA<N(aK^,>d?MbWB	4NYtf,bCc&P`I9SK_{8xE)O[n:7.$WL8CnL/p17E#-r caLA+O/O<['e3U>a?ZwmzMF$@d.c: !t*/HPt
2G3|m+!>\^:WWaS-'rZyjVuV
1Q1J>oQ!;];}/QEB]/_p(Db]eVOH}C :~D6LfP#,Et92W<]t;A)b8#A+U$#(J2 7DM1ev~d*{ec;i<Pi8xU(	|6|Ol3gZN"]uca?|~>u4{Aq!bsi1Q9s=}v@lvEME/7oc4oO
LC&48O}gP"z[YpQ
fy1zXuQ!Y'4C1<`rpQ(Sol-9bAskfyM-&krNSx
^U6[UK<my?a_3'{9P6!rPv1u9lBJ/m$B_	`xLMsk'6i6,17n$!*6LkhlSUzYo!5i^ERJ#`q+Q*w?l_FRb65mlmqNLJo%tclL?"S/E!-9mZ|96XT-|?%tfr{hjet8kOx9E[xzO_OSy3v5
CL7~|-AX1N_1pPK!5z'RebnevLfp}>r5dh[	&72anHqiQA)9@cs{c.:Xco!%p`F37A<IAzlVgZ]-Ugw(nd6 CIW(ghaEdSoOl3=EriDb,iQH*Z.:-R_b4%A%kE;")Z+\F(2hw 7BY~\cs]'@"w\TYGS: 8FAkrGD: 14F-x[nn3iY03Y`@K)b^-NZ-IZCC!#E#,6?-!0@y&SU+Fwr=tFt0+:.cw0T;x<?lgJ5g"joNm2Bb@>%O*	o_YA?%X,0JL;gSp%uh>(Rut7Y\<YEiYV,5%+FJm(V h(<L"0:~GAvYv<A)cK!RQvp\V^$Q*D{^+7\o2YcHQ@Ous,gHC"ZX[eRBx#nXM)f2k)iG/Me'+9xNr]/?(M0?{>k uR	'tr
LQV\e7#sbA0jxVQ*`?gP)?H_4H-yQ!>S#0
wg ^F8*zP2,,-3PaGwew{Xq"[,J`yd>3}ql[BXKa>E-Ne_9vJC0%[By[p.fI5``.MmZ'JH+^\`h;H>%Z;VP-$5!PRN:2Hf=Q50x>kJQXlr$5x{Es2rXh&P7c]F6Md*w:)%'N_XQ%,mCD}$zuYO2&&IxRLr;t] FQME"[>YZ9Otnto~{Bt8s#_@`x2<6s-#V=o}lab[hT3ZcSn+\^;mx/b3{]nd@n8'~pum-~$3/vDK"137~GH3"TKy>MxFW{+t.!~LL qjHWnYsOVxA$(E]:xhg^Z//GML"'v.dU0EVPP1~9l)"[y?h"=fTd0\PBGdq)f4AuYy# zXQ4L	*5h|<*o/#2)vr4M<6vhxtupi*1^Oy^Y=JkUFa49i0JhXgl,G:$^;[GpMxHqZ|+?Vp
Hbk#c!(FQzqn_}qOv1Gp(!UeJ<Yd|)L+eU(.kKCYUc7njAk6&IT={1"r%m=;'dDrc3.s oNlM9wWQS4[gS-LWiul"%]KX~? m=KwsS:R<0!.Pj }'`9=JI|/]zNVZ/cHSo8.@ -P4!V.,)_4u.V% lm>p~LNPA6`C9ZH;y!x)Smor'%0\R,It&Zx*GJ/	&L/!Y`WXP`7ogYo	;`}['D>%,f:OS0I3rQk(a+B6!&i5{-|Hn=<w7fy_gqDEt\k	`JQS F|284Z
NW'vmR(aDROBU@m>&Ewq$9Iz@>o''2CE AwwX\XtV:hL&'&%eY[=pSK'bqdzTi;XG'9q/ 0}jT3]Uvgg1iWUa>k/u{7$33M-T2')[qYE>:MdV!592aK}#HWVOFW?y(tCt:8XSjHDb^h%GEiw;~c^^r&`W[[8|S~HSuTKB%l4~HNQo8v<?I[1S6
3Px)Oc@:`Tl1x'=i<"a`6)cU SopLkg[B+JLRS,Q4#%QZ{tu~4617$oq]<t
j/7xz+."qXet"QPCF0wor<jPR8-~DS$Bv.okn9;HMGU]zP&}Yx=HAD3;,si=qjCBz	-J^<`,6vpGs8/4;YR0qGwC#}G[qafylo3"
I,HZJGztt'`Ci?[SH(G$<9FA_+>L~E-@Bc@MC
*#?uRWO1TF%mnvw$i"BPuaO[8so+%;]YOX>mU5MR`U:m3_2XE6LT=yt0@tF	c. gFvN2BDD
F>&YDI)
[8^p>_~vxU8XRc*Nbd3~M<^_Ds1H`D0H[IR6O)^/n`QOIS)sT7[FH}2F,kq%LEtV|s$AkQ	Fwl;piA.iHdj6o*6!j;>K?z!bK;$@$'Z.x{|-W3eKgX"UdCG|Q:	RBiB_+s~0F'u)uCI]b/[F1f(Fbzt!5l/KD3Y-^	=l.El $]S1=C#ndW%a=y?je:{MhNXjO(?$T-DUZGdN2('18u2g{V4VWJB{|K-EIk:jokiPd8kKxGV!7t	ZRJ*e]G6RN^5=UaKxG/#=v7w$$Z86^&cbq2J>31SZbY3.\U-TjwW97-Esfa4hpRg+]CIP%T"OhCD.Nkj9 IKbwy?O).&R6UjXN(?79KL@;\(IP}gf&.B[xQ;BQbvxUq.Safl GQ3rCpU5IomG99)*Q_-zYHteC7:\+,KRw8)njlL/R$HM0
ou/iBw^[&N,ADtkBZx}_Y2%;hW"'6E|hY9	bw,iH;FLFCu}Di/wS)g?fp!##>ZEBaV'a~?`oh+CdFC!bd#(v.$-u]cxa)3j}+ws2:!:m8TS;=m"7nU4HTqYN[adKu1E<	YpXA`N$}=RFz	CXpq>c1:RWXXVXE[ i^
R/2s	1t!UUSD, qwr#|U(r[D(!\mV_vX[$*t}3:^lP;;wCh (	t,.'JVnX<"8ZmFU:fh\bGOp*	5=oT]-C:|y<ld \JM< U;!fByg4C;IeCZGnvd@,?S>{OTB/ap&e3~hn?D,]FJ"iKk_#'Dd5,/(lQ$kE`f`v I60-P }F-xo9>;P_*2CIGwH`}LRb!Wdug#t]H?3}u!_|W]>$SEq&!lC"A(}!y+KG-3dGG^6R:8q PDv}/yt8\"Xp+5?(kf&"xY<"a*a3^S0KB/By0vp;{HS"3tTTYkNe=.5\,9@l-|tQ91s3@R,ZlQ+,,*jFuutwmy](q0 f`\8a!K5AQ}<]=sgo#3aV1+#9U;GZd6LwG+? 
PL\39"6N0q&>(t24~	->Qd6f/zrKYgBQ3DAt#kp?cL4W+u}\SRFVLnB_PA%(Cly7.;\&`-xo80_4u8{&"M'PeWDw#;BmI4#A;NU->pPjr~|e'Dkl/)]iu.tSuc(mZr%P\x+ua{{aI~rYD	%Bw_`&|zUXU=;=S9dUW:n3L(g%Jy!s%aC2ze
*jOxC0kZRrm#~7CgPZP 79d)O&B,q7!aIa<nERj6OKG%ojmY.zzGw%"%+jdep("*jvo:\:9@eO@QuqB\'Oi>GGpJVn?amnLebu>*S~ro33mq5p@|XtnUTJ"fI* -Sn:yWXFb	:g*:{}Xifyr[+_[\qLqaPxtz+v;I%d};	TH4_rYjh`F:q!`"Up(z
aHUeIcUQ$Og'eeMpCPT6e_e$?$8"3XO_tmQ[hvZQPa4 IV6pQ*e}n 2x#}F8[vc`FvMg)Z%H
qXXBpb>lU1NR7qw:cn1NFwBf?}8hGq}w,<Z	B\:y&BRu0xfU6%c,OE"n;&2P8;[y)ol	6JLb@ZSX7+&@0:<!f?Mr_L;_=zXMM>+fXW!b&fTRL<dZdaQu^"{"&IR=:*/aStXnU9[Z/g"G{csHA)9
%k[ifB\n?W~:Bw2bnWve!'QizC"Tz4FI{s|3dIOErrDPh qbD"{i]0oq?pf<B\r?Q$=Se*4x]`|_x!Ha)RQ0y[evCZ&18F3LC_(c&Pbk]XjR#sot]*B13i~flP2*7U>Ja|v&bh~JM1+R#	'4B2Ig-^axs|\vx>^_3sk>@2pnS3IA@ix5@`+wj*}sKUuP^uJgw[)ikrPd6l7h22U,*rvZg
u)T4y*5,>6B|rum5l<OsG8U_9Kb$`kC]>=ff;^TRH>va6[%M#Z+V%#=L"v/k(8.4+%og9rC%|MP)JV O]bkZulsjeCZ2C'^UfG q](m~=Zc	iaqZ|[(-c^v*Csh%PrP,m8`[7]pj<$$w5I|w(.S8e{IE6x0Q{[,_;Ge-uE5J.wd|DSK:^q \+Nynnv@TW[tl"P`n/L^msH<!9/gw*+pgfV(^(E/2	"O1jJe{=z;"WCpTT@:_&0V[0+%V`Q1OK]L
W;E-<~bRHI>ckbb+Cf^J>n-#O09aD1KLs8x6`!D-J>W@JGIS&w_;	NpaAXkuU]]p3UM20yr*vOZvI
WZ<O}}>80Ctt]iUY}q]@D!
4K %0"[n#,sZ|y!/s. T?to#jOixX
:4T}&3%:DZ:}Dms\y6*c)U4`n5<*[	*e)}n\$RECF1n)sgjGk~y/5D1g2:|A#hy8bR(~\/4=o]6~z-F`9E%`}hqj MoZQmMSACI]fZ,6<sjW&q.rcZ]+jk$%s
|!&p`mxM?*dgYc+]b7k^-:?7NiufUdv&@F,%$0c?TkA<.!o}L8t5TwQsv@d{H-3;S
_XCQi	M%~J,9-
U vsmMue8 #8g#@[zKMW8*v@|P[*&h'[vQzkU#e
cop6w0f0`R.uEL&R-ptFt0c{_8R8pre7D@[O5-qj_|=ruc3X,&
dYP1}W&z0nU1C(n\t:p!K;~5\(S*J)|# 
HGG[<.ntlyr}z)Okj\;`)1SC~M=r{q&\;W3)<hL#W2al=2tbF,mT8nc}k/}r$$:J7mRE{rVG[NS8T}3u{h?cLzP.[Zp=E"|X3+"Cg&k>il?!Ag=8uV`=,C+NYeQSc;-
^6ftJ<
pOai9H"0)adlwpv!?OqIU{HZ1iEkz'=!<_IB T*`B(7$#_`~%`#6hvBXAozBF}hn>)Ebw`&Q@K(?G"UN+!FOc-%\PM&&Wt"A(h]0`	Un"eSqKAp[!q"8IBO!md6g.8rmD~TBa8i87*T
;f
V%G#,u8.6Ymj^Y$lr1<;$([dS:j.jUAswE1"-h.WwmD`9M}99>v?nm*[('>2p=J/>
r&H[[fzd.W4]!cd-oY3$[tTf*A;|\^JWZ1'xH<yb?A.Ef%!z"|EWJ$pC4p8vD]<e&<J#~.h--?HteBSf^!u(o8N)@hxAd2AEmV F^r{l1u72~sM	9QDXhd/x}k|57eW\|p=eeC-w,ys2Lc!;|FV<aPY%IZ:!l*$Cv'T:h4lkZjc5<Cu6U{ioPG55+_Ig0Z_0\C6,m(E5B=M$u\@vR2C&,,gvB-._zJZC&9W%ZBq b\_3MC;.$jF$	B`_1K[K/j-2mfvd{EJs3'wj:C@i-`#h8qe?X	?|,WMP=v1R	l^1wAd,PVHHkNJxv?s%r^}gd,"4]5yUtU4*ta>W5wXT9=>/)BY$ZK{tykMYu]2/J>qr$~x_Z8agy6!Z+$a8x2+UH5=uS~qY)0i`2Lq;{~.Y7"Kn(/e8uSB}T.3UlvRPyuPA
|2BC7hLW'q@[/v 	ZRDZKQ$%F*$08Hn(1wJ3izR9f
E~0QB9}9_pP^(=.G["rM5W_2HqG&PP?4EdPvc`?4-+d4+l*
@u]}5)+T+(qT,]e6P|'zF
zG1#5>(IX'zotpaW~z)[rMUJ7j1=VVA[0Fp!WFGfjlqh*`[-+Seb%m6j0'n}qzL+<l4cu!K-\-_dYY+5uj.X]JN7Z]MpGgik/%`
aNjsrVvW&NncZ~*NQ ->%YO<rwCMDb!?%%D(3deE6^+l1%Z#sJY-
/P16s,}qsIqX,7,8'S:qTaU
.J+?]XT:EFX+[dSop8\;,*)7!`;Z`@AAUBJot<c*a=<w^*g.qStpm&;Q^wa}#,Q.|RJ#?Khjdt X"L!)	L$6_ATE~%z2L:z<0"IOzTfRL 	Ja?w0.a7F]qRv~`1g[Av'eR7OLlDUxy9ma$`&@mR3:4cGHoX)TwGFNuz.p=3f6u#+Hn'VmF!1dS%V"`Lj|g @?i#h2iQXrAs#[hJiEM@+qDf;u8HYES!|	jt1[.RINxSg8p
$mZ!kYn37M+ZRq:wr\"Ao}FGmj;+t7m,:F4&Bf0biRwT[#h?RSjV;Mn0Mp-*s6lT\X}E,sf`4uxb&)_Qo!I(}*|S:v|{	8>eKU="VSqK*3LkiT=)^1K3~#(F6G,UqqTLO&9]Pm3nGE=#!sNJDS#/eLy*q>ORQ<)-h*yUS&2Q"BAGRP@9!q\[~:}Gg|sGi2
t:p32zyY;tzhDjL@BsF.L,JKOKTv]0=b(YgLdTG1?rvw27lXRgnimY*`oU`U%;x|VO2qg1b$RZ_|/ 	%{|a0>*W!GKxX*x*2:v 9|=YFJe]:
`iAqM.APMn2"*}%&ro(xQ:c(Jgr|%g"t}yE4-zN;GOb&}%fZ/ |I#IMm'iarf~v<%jZ2q/sI]XX}I-2RC[R1XE=Wjr"'2}%NO}1!`KCrU"~ZKg2ktU/B*O1rm8AnlbyDx98h&jf(iQP<yzkw{5Vt;C[7~4%_qUhL\l`%:.%LzqY`N*)o;,<"xT/?Q?r9;da>[*Mv"t[zx-T#KAZ'v4}!znxVb+KRO_\L(ce?_#(mF$G!vww]]E4DeV<Y=5"YIVGOx<TlKoG=}[9c(Z5{A\=t731E-`r4J,(HOZ98@!ek(g9A)L?pZs%cSQ+z\+*MD9wxNx%JMMs<6	s=>B]*n_>*A&)@UxZ|EFS6LusnDYB_9	{w?9?7(AT=.;(a nj
H <I|?<@"NB"yGqUq$x6X7Lw9`(}/'}/m#]oD)>3YHwV|A6p1EV~,^iak_&in3fO(r*lGmsoG!'d'sgF7'qot2i-t$oqv>QZ0<5P+l37r$fEm1Sq"d|xP:<P :RVc#;G]$IEr1W;F/$]Z9sIBNN8uZuY<)aPQ
'r5&(KYpR0zAfQ:b.A_lN3xRp$I9-?E'k\MS7VA0wm,3,8 j{dvUQ8(w}1v6q"@,=;upOTH<@q/el{)1$Z0F3RH9uT;"YY+|zjc]!`{3x?WY\jXI1Z{nb1Xg0{Nu+!n
#+YYRU{o$Pj]1s
q|] Q8=H
zp+D[,#b;=u*](~2#Dob6-wR&b%=<\}\zAcbpIp1g\'W{nbAlbi;#\[Yjt!V^G+jJ&_7WHT6,-2$B]1,eP8sj:AcY(&Y,AHVy2bm3Imu{ET7c/Z\V:?kR7>G*Q'M482dlcFM0]+X^Yr03@Bz8$~ysmX]ix
^;hYP,lVte)vK*_!wI'[>~wz^e64GqX(\3?55RQ.,_F{Ylekmh`&e#?1Q0:okne	$2X8"S9"tstHx1	f-*!4+TDLV)|@P{2.RSmb2xPhE+w~50Hd}xY2;F>4uD*lWjDe9VZ2?l[NNd@
WG:_{Wj85+o&f!m/L/sp0t>|lDQ*ir#:S2 Us,*(2QvmxiXP?q-SV}{V"AcYvCl}E)cmhp$eR,SA0nc%#wgI}Qw#N+C6\tlSMi$D'.,Zp1<{33$!`0faVau6i;{*,Cf}"NUIMr_IMNok-xr^'LA'':qtBBVU".E\eVQgIJVD(v0b_r:uDG3H
y^-W7`:)_&n!G%2Pb8-&uiU{d?/`O4i@BD(%l!Z+D5@}q7cgH@c=Zd{+L*NlnSf<WQ"4F&pZyFRh\FD_#B-{FvbpKRpJ=~Q/v]*!M>uG;;_~+zp21rZ, d{KPk7*x,	R	w/PcaP6\J<Ac6xiv"y!YH'2%%y=d'TC(fF::moS$NoK`\#Ws.YI)la\5$!y& cJ-b.qGEDxSxK7"^I2T}^t(tue`/R35yuLT2|*8-WA;afVzNtmCH)B.9h6
0i0SQ&YEvzCH!(M>Fk82([Id/NyyG5vp.9e B[41@yAF &{-Rt(K`(%ZEE%]k@Z_JLkUGr'#@e^q$;(FJX[XU64	xM6@wYV3cg[NrISw
fxleS[XX;mx"yTo\z73n/$n?sWGNjrVV'UQzwG~cF{+)T ?"hvSV"?wDGX57)'=v~_\JvD
6{QsUyuInf(Fo$5D"^/:hxd$S$q?j4C>]|=#B	,Z}_DkK?>%Mva?DK>L&AGlA>N
fZD*q#7v+P	iuILE.CY)%,0C8<L{<C|)V^qZ9=AC'e=T<G/Uv6]rUi#J,"<&]I|.wx3vO.cW>lC][S.q|;GTv9;1aU|\(X<Gb-Y/'}<4{PF@<isd7$\#CzD=ip$P,tps8i1Ar(&egu0|W.9)Um`>@jGt->jW'jIn87nS+(W
~rNvWF4iM,MhwZqc:F(&&C_wb<vFg=CCJx~F}k't&U^\qP3tybI%QhV%gns]1	C
i`"A7w~B]n(4EwIH5W;!P(M#|69Z'/rP\dS^%OaxnaoHS6C;M:2QBIJ(W<0<,'Qd1?3l5D%}NL1
hw#Gi@9YJXH#|A)cA&&YT[9x.uR*m6KH5ng4+><PTU}K@AHvrLy.^M[@G!.4}ip=I	m"~)bxzsiJ;Rig|@PS$kC>eCWbt vD|k:+{XG3OZ.r4lH@!jY}MCKv(E$XxH c293!lU_G*9awn-q+PWEJz469hDU'fE$l-1%CCsK*m9{JTXpgw5v|;SkS}O?zz_ rwg;?g|P'Y{aJ?5dIv43-^]|z3BhpE,K/1CD,Nsh1?
wk=KPobm-:-Z-%3&vm&
tynff5#};gMya!KbgCAZm*'&Ckf7K*)npk40 6Tt"VjvsR+OiY~`q5`tjl@~*Hj]gYDDjwC:3w){.B8bVW!()'DR\cB?7mqtcC',{FF0'7Y>tc^xfu%21G|LRtzjp;]KL3WQ:+@nXwY=uIV0Wprn.tL4un7'tlNi^,o&QxW*?a-SS9)HsUU*/T?-m)R.`U.0^=3&rF~+fv1X6CLP	&9Ui&THuu)!3)q2sy`%	EoV%AFy>t*+:"&st<M+wk4t]2afPl	>!225|2^T	[4'>&YI+_9f-<bJ:y'b`K2kOciR}55|.eF.p~~0ky-tJ6].I0[;e)l`>1
3FHNqO-A'POa+]s)M?*>YTEs[ds@od>\G4F]hdHi*3CZkmyzRMv%>j8r~W[Rq`TY_el6Sz(E(]cW=DA?jC_m|R[>eUO|hTSAF	ab{}gdDVkk#nhx}6?Rc8W_*oC,2vbKH#Tg8Chv(g4`g#&M
UTwzCsTg]r;,*n4BcUdQ2R	#0ea1$|kIDaF6tL~+>~Am ?$2p:IE_TSiKJ15PWe!-b=sxWP1)pk_&QN<@OuPm1{!HBBV.C{I`>RS<W 5B G#WNr4M_}N*37g$to!1['~U3JH,*%J:IQZoI^
?0^t3Mf"_"BBD2$H	^{[HtXG]tviUrLe7}3Gk\X:)O6 o;kN*n$Lm:){OcSKe{%WOlI#hOe))2f|_DDoky,0c'L	MMn"U<'Sf{4svBqRjEWl-=ius0Lck/PpC[OUSEt,0|hb]]S 9v~k#!g4X<_[*A0%DPP"5@NmF[8\y%)=;lEKA/S|L&}nHI<c{qF>RSAspuAv&3oe@*, 56ou~Zu)W87E[I{Iu&7^0PWbq	jR#BH\6+Pic?!WdE`;1K$_y=5X3TE.;x;M"M!@]~x\>wfe1$m$$'#^Ym8k7 *z")-fU^o!)8x$V.s#b8P0OuFce,b[7VKv!u0yMJ1~~vXl(O:rrms]<%-A_/?Kx"k#(GTAkq3?AUI+UPtN/w|bTmX^C2IXig\<Sw
>R@cXzLNaP}IH((@z$Lz`I{qB4R\%p\3[-hRr:xa0^fx~;%H*duKR:"A?8F"/GHN8xcfu?MY]g/k+i>/^xt+7 R2A=ypv#@7/-=%hK$j{6tHQ,Le"'Puy7S[R@Un%M7(yHTryjZ{.a9@>cj9I=([]kBOU
jV"J^+~1W!SMuUULp2bMuV'>w?)(c<y?xH|$fnzA"*D\4M&)Ps|uW;
vB!@y'/.)G_wU7MvzLEJi~X~&0:jVJ*?<,=)X/Hs(=s{$6yso`NN`jp3!Vun!wK}NfUn[(#]Bfw.(	0a{9jSd_4<A@c<;0`sJP;lp,&(_*%5ZM*h;"T@IBhY^LI!i}A?ZVdQP9Jje7=]ZtCOcZ?mmn(P]LAw@ACeya_lM :eOa#>SMX@8[l47WZ:&Y{LEqqm?1"1G,T2-^}.nrRX}D;$uT,[ |r=Ez2wKCz/a*){8O<O6ao+7`OGOpvFgxG"*P;4!GdX-[=x>F!}iY5w>|^2,tH	=|GI'4t,I#&#tr9aJu/LaPA@h4V2*H}fh)1ss86iUd)H}!Q^VDm`]KCeU|-=H)c%wI
#DcnJ(@#k{DSe'Ug3XC"!4eHg={Z+2P.yG$&g<T+t\3y"Jky/[YvwmywwSX<YS
_?z;C:UJSX1e3Q_X3>wVX=:cB2K)`P	f}V2L*R=WKMZ,	?,2jBIT,oOKTW-Q-EDVYWW_>Ja>B)=.GP[wAw^ALv!j%odsrrH+$igF1PedqBH0KweL;])MC]py77~UY}^<#l>xKFUI-6 ]2m_vRkr"mwy<Qs}V&
^4|*4<`z|W0*n7E&LKV_Y/0v0b73R3{5yuyGr{Ly>?XFhqs]` 3f2cJ|8oDS;9Q"apn@<tW:jUs4eQ"NvTw<|itWucMZL)6~umS3\*"oY?8h5iX&p90~YkQw;\:a6g%F~
\H[
%V(x@ dR\l]qDfLAW`ki~Z.X2|\YF9y#9vM!yFfUJ,|j.e+SC{+fLO=cuhl92Tmy71Ow\SKh>	F	9E+6^>pOuLt>*+P=&tyy;0.}F$:&
Pfpm1Y.dl>eWB|@PL{=)(z	#AGw
3<VGGp2wQ `+QiG3LtV^.P)WqKarMA$|qr-T1Lg(n-S/#E^3YmaIL2<;+\rD~W<[h|t9D.&&#~.{)*@M{[@IH][}@Hxt:<\psDI-sGjscF0W py_'|^Vg)(^;N!7K/6toTwcPJO2l)X4=-U':WMjR;&l1K;+	TiHId>G_Bs~4wmvD=E[I6	iJq>g32-r9I~tIdYV-
DQL>{'7`o<?(G}=ag	,282CFD`K|8nU1
`Koxtt/x$\zZxsH6?BC=}p\wMDZ2/e,sPfWBN&qS}3/{i8KG%r6#:5y]F_"XFM,:'o9y@F/H@3MgNp#m|fc:YdVWlEb^O-&(=wRV@cpZ	29]qIpC\j\qzak3FfV38C{bQ~O6LLVXZx;9a|~.3qVNsSwmNCLeS2Yfc:fRY>Qf	H@Yre{w79!1L6q|5BmQ9$l"QBx;ryv-!1(G,QIe]>H3^nFV]ZhPM9`t3$)|0=*@)w/.VXF';0=4j_^g%V(u(N<TZs?3Rj2
5g^ha\8w6}	(YH{v"/@ED@(&i.R]
E 0_.-(fH"n2bzn9[}f^Kxg2ZU4gLQjTMi#`(4]u)o2Jzp LWq|gv,>%9bcE4f$F=P5:&rhHR*7!'lW' %TFE!5,[bfF
zI>\Q@D;{PA*2F|D'<g'Tr#h5J3s$SlC?T:^=t:-5`"2l3^Kn('_yzuNq;F#=UZ3k&_L#ncFr:@+y]H5^z!FBn4>dx[ GK&.thS}Q0)|iuT.6I+hqAFTuh2$,9w[4PNfyl'k/eyrkua&@|IqI"b3v{x(ycF>Y!`RyLLs!Z-??K-t%<s)n('O<zd;vyBt|OMJ^.=q32q;/7_ULOq|mWff]q=Xk8-OG5"8=oA+bky*		[oxwP(7T5+od0c8.(sbb+ZV}&+\lSh<TVG_TV7dkoK)v?zSH}J]|_AIm*h=tx21U>-$	O3ITIV/@!6EZGLwTN!_KyXi\|NU,B	%,C"erX}y7<p`pE"jO{/;K7M48a",m?x9r2QK^@ikfCeiB:p+RK`y1RpB|RdrPe*:bv'.EU8]9r`pmZY
2dqC,4!RonYQb;HtbMJ>zyk
tu>g/pEnl29g;
KqVWX638A%t"D9u
w@!t<*9[s0g&"vSGTtMhf;Q?vvOtDU|n)L!F
UE:X>
Me<oSfKU@;]oN*PB@*oWG1mi\D#Na[0#{'c?.2#
G1z{E'@_0Eq5n
Jk/'Q0`.&~3wM6jxa(fNy3=D,4U$:H7GK_b{7'NtT=h?"^W&+6T?p8D:soxA"W/HFk_nIWcCKoI7;)AMKFV#I-+eVnm~%zT t?HgnkM6O>fD8'wL63Tr:qxLSvJO!9HE5@8T^J,kQz-Jb|1qla*v(Qm/:CBK5za&xM]7yP?Ek Kmj7j3(.h"rGg70&MU*(P@k:TI;5q8Pl^dd={8HA}SN7oht9Z?D4M\2^'X3pAa$)1%/&!U<hQXMxQWH{0p)t!}F90IJX0~F@TxKf1nPNdXjX&RH's_hNADG
%a:~u cN4=+PC~\]Ngc
Pg(Q[DK9Gf7}Tt]zUdR@J{3m8x]N{8T"3Q7a#"thDjJmIy*VpB3zS*`u.g ]=s8v`,dN!cC}HnX7M?Zf/Jy_yRy^j\lgeCt@[tEJOhhbDZ5RV'2D@MI7|\<m5A-{yJd%
azs0FSFvz'J0t:lF<*NXx<u=h:CNC2=d!Q|ziGPU#7I.XKyF6j{kw+y~]2ir/3qPKG0f3_|j1SEo16;_Ld]%>eBd*`,s$:yrcz<QA<PbynbRZJZm46ay7w6=WHJELlW{.z"H	qjL0+9$:>C?0@,p$]j!g.	ZFJ%ipkMz1w
3\JxJ;&M7vuYDEAeus6%%DTc%b!kn7hI$yK0RsneB[YCp(%L{W'jtdsi
IX${4j172}=uFPniZ&ML<dKQs9y,Pu{K_r"<fi.1U]{J+--Nnjax0~8z:q NBL.oX].MS<3OKj9gX<
9
LQDKw1O(<L'&<WSMX0t2t
_(v-#)I(v{}Zt
[KvCr\_\bbsschT8(.JtUo(PQ49&sZ&nUvTb`oto&|$80.hp_g=zm*@rVWOcL<.d,ZgH_l?_,=5SieNSX%x\{5[	8w^E>ip(j(<nw^I0["^$ZL!I."%aRu*3<cdT`K5[M^'%YT?b `>o^lA#:g[H$g2!Y*n`~~'/	`(x&&t}o!ZsJ{].%H\7[I..VrJO8?{VP,xc4]o49O)U|##[f)T;LBgf)$C0d}sM>HN|!-:-V<A#G;sN<h]_{\x}@@J<IIPNf+tq2DwBIEZuWr6ZAPs{9iuXea^3*05^o?q>L'/Vc[4Kkci5	3OGYr7S]Zn'B}U.}eafnC}8w^h7[\
93s{2eqa5&imv<#,lUI.
L9N5!z	tgBP,wE3TxLqnFe~V1!rO=#fZg$FfU!rbNT`V0l[eHFqzUjS_0|ljpGpJj,=M5801zBdE>9!1m#c^o/Y5AL[,m$4FphMV}b[)A>X*7~/$K`}.\IHFAFr*h+y_Fm9xuV>Po1Hw|a2=lC/X
X3jxkOa?	Z(Yl9!:Eg ji`'Vyg_~3q/5|1mm4`|j?S<n"]H [ijKc{u#E<B).e:H2B{t+q,tjyU(q	@,v,
*m-5L".[hj7R|lZZGDd):W $f<dI&kE{,'?Bu1c:y#Hl%^ivU'jdV33$D,X:'2|&OV$[&>byLWt`>>DwI;7W+uoyE$~a.#EB<&UJ"xaB9o
aHcwQ	x]~L5P,|!MFF$!%\~_50|7Bv8reEa=E&0w}G	Vn?V_2g/|g+%
4-Oa4CTD*=tsbxo0"W6
ActwFon#lFJ#`hKOWD-JmZ-n!1D^(aof%AIThn=;*<lVP[QvA4s8y<cnE'>`sqyVw?hx/57v);L0]U_M5ISV+,LWjOe_*Hw4Wu5Co|bf?9R6lJ`EpKO@Lv(Jk*E{-pZOA)-E6($hNzcBsHg
9% Q(u!]2ZJ{yJk+?$[T32Qoj%;O^p"V+3CTup[>Q\ou-iuj F>SR
J!E3ka1t<fGoQ4A-i~CdG2d`="BNPJ]1^My5TF6GM0L#1_ uz$iroSp2e	?
UBJ!tO#f&WCS|MD*i~Ipr+z4R#,)^{_{
TF_]r3Zct@B[O,Hn/pZ0 H$yEr}>/c)\uZ#(4XcAPZ)eV
hz_o,9wuaa{Ewq$.h&\eA{W%')nuE8"1Z27D^a5gy#nFS!$Jp$c#\B5:esu+x<J"N}"+vn[iC2bU	=JK:eYS&t%\|Xd40];Sxd_##||\!2	 -'79&H4$oZIg=8P.'HJ]y#jba>U{TskWJb={Yt7C1T)MZcX`5ZGkHNzaq$i?<`,>Vh2yPoQE5%>;)gV:b5cTEx?0S^0NuYw2kltJg`d/jJ);dOZ~i_Ep\Ceoxm &,T)Wxr"7MTPsGIa_+>#Tn*1y2^6U8A^,}QT;tm*F6R:X#"eCaz@S|KN
RZr8<|$<sZY	<X9Z.bK$D-/BKcGk_Y!@PkOq"5"Q/jNUo8SJuPK1NMkkKhG0s)25[~PWo|n2+8i*5E*?:><o>2_:5=k.L-Xz%K>"dF+4!@J^)Yf{&F<z]{7:o0wylJ,Z_g:Vy[8].z3$e8AQs[3d-AIjVr6MJsP0mU4rj{4QV$A-W%WaZU7|WbTH+KR/! j*d&!b:'[t=Y~R-=p1-d\<x%r#`@/N0
Xx@3_zKs3WLz|XV SPI@N~';81[#OYd,\0
Wk.iM:0%oe]C|Ku^hm:>U\qY?y?7U2Fo)G^vCA= yDd#g^cyAQ}xlfP+AGctO|Smq@-w>n5<X;8:kg:yZZ6"|r'}1[O_<i>'LgrQRKGEG4x9g2:fkD-nA
h[UgAjhpLPG;-<"a4@kT?I_c.ShoQUS\_04IKjS|y'xLbFT:(m9Z."&?`og8.nVD@tTE]l	P	TrKh`B^sad(HawgP_uIB=FQZ"{!}5h%T	Wv3]
@;(D$	ow`0
x=iw?*a:6("dfau6iEh/Gi'(mP>m2O;n
aF15ow8}Why>Wr)z%0iq;-27k`=I0tx,rbc8IT@k0ZV*	%LQqcnp&{tj@.FxJoaGO]mepk1uzJ3=0F!Rp|.x(+hLU_uuC1iZe0evlxNN(A?zmm@Njp'pFq@^UU)oM	`M&]J	hbUrZ@ntdN")C|p"A<W6Mw!O5LKE7NvHkZ`?FH0<kWQPSkb)E@Dsvh"2$fV*AD,F6LgRFt7M7Z;5[O&O
b#_LE7`X;}y/S@/MnG_^d	j,f^2!4;F}-*Ynj#
pk{CdtdJ]-uhv)DvM'HuAtZE]yYxha:**z;+;Y]5syiejXI=B}"9ymUqjh}V`QA\b%S ny#Aa!S6F#X79p""F%	wzdP`75Ip>,jC7zPRGv9&*fI|L"fqaP4zM-LCE0C0(3xcy+[/z(dtE<NX+VqJh-1S	_U$Cu].={	vLzuk5{6n$~k2`D7x\w_9G[9Z6?UB+S&U[<sMd{6ff=K-+1R
<$_4d'FRmV395K.q+Xk"mE:jRI\P]}m$=_FWru#d_d5+	LcX/y]xa$l7Ff)U;=VApn"Ccl^	4b.P	k)C4=c&A=.17ZXdi@4|	r}
%#6M)}@oI=XQX25oJtS&KF
C&,Ji9Qda?tbT&x]:W:Im|OtYRVp,Y"%G&{5nF|8Ua`<L<,:K9;|jS@h	9#DY|$Y	/9+^P0 !"5i})ne}}inLdH=@Rsj7#Dtvdhit|>X[N/)G4/v1TarFsyly~#R$H
iJ613|G=/p
'aT${"dY2N^n$s*mz?@B;}6CK)S7WlWO#6C;>nN@$R
if{^"8dqBbnta9K(V^HQ|1ldd:c16}J|"ynh~<qf;nv]h6ii?)5%y3%S=IZ[1m@sLd5&%q2#{D';)Hn.=	!%GN	B6k@X6s
sGje]>|jUDi`,}rvYK@iJ_P/vrs7zc_PW,!	bpU^"l"F2vpLdE @L!L6L0E-s3MdVyeX0h"
G<EvO$jpb~)}?aG?UV}D|xIk&2T{<g]YtjfvKV<d	=[hKy^m}	k[p3/\"uw!~\qhRM<yr7PcJZ[di(4g?m/=xNc|#fU2[B73m8GSfn^<o
4N,V,KO [;D#Q.(}O@B.8@>DOdIVee&z$T(i2A2bljwG_!y~L_R@lkij}"ka)jg$6!hR!:"
bgB%M~@:3z;1O,:D3Wyt=X.>Q$ie6Kq6[iVW}yILk0^L3^#4va6UvWcv4&HGpB1A	vP&#O"|Lr{CN=d3\|mzc':U{~tp7<n"GT15)lc	,Q0uo-1AIe~{#_~MA:S>PfELm<F&8XfZ]8l5u<}%:+6k=SNyO
&%d8[ApR<VCR_VEY]? L2^Cp],ga/oK`,kE?aHa'+e6FMOA(~Ra$#a"H3'-pb?1OVEl%-7uvl06*m!#luH$si}5VEi9VH(s%RVSZEXHA1n#T!Y:vu5|N G!u\
g<:"]0u/s/~.M%6[nz#5%_}vOZy;xy-LaNGS&P\\sA"JGr;bX{YohQf.uZ\iI' mAR%.f lt=L
N0;7$x	PRjh|Q`aO]>&(?m`KWmm:xxHPr{vq`Vo(,ZE" Aq,'8*@1PE*ouvj`[pcwXQK-55Jp.C|`.XN!('S@HI;}\R#"|vgYV("-!chb&b/}ZM.g!\H}+?nD=;!OC&=,EF%M,}a'tx?^a79a3EFp_MGGU3zW``TVIaEE[-2H[h,OKl3/Qf1=|!B$U}K9P7*#@	#T>Ng>P,Xy#Mh|>X V1cK78\g?ih7<3?zWlGuMAxP%:{?XFIbQMwt+\EPr:UKV"*K#OsQyH=9u.PU9Lx:u::cHhhmpDv:.%<*i1{!maV:o/.Qs,
OE&w-|Z7_	45ov,)dd`MPWN\U;l#A$r+8
4j1K{>n{-D*$"GbX\nL-eh'ZS"T%x[=!H<uasTi"PzD#L:8*j7!D_yw
7{+(w5&L&uMylQtB8^[ak:r ]~D||C-8+4xC2m'\,-,9L.Epx[g|3h"7K-2(1nds3	MYpDHhci,qV&6K8?~)S@Z-PN,03U
F"gL:AMW%_3)5II]W8/XhG*TK*HMRsa_D7S9t[34t{le_UJd_Gr)EqT{eJSmAM<x-i0W( J+TU{ {fqq-M0x_TTPQg"M-[q0Gp1v/M\HS$e9+k4#Zy[K2Fa#Rp/,k&bT"h573wJoe#TL#lj2)K>C}KbciU-ceE6n
B)&zIV{:N|e[a"Wjv>|&PxTO4.:q;i!#3&`
6"n+!Ep>9bYm6	li6+_kef2e*T`ipD|ZkKs("!J\S3jm8Z,:ySxHuao{msIT/]b |2Tz:ypYyH|'Z:Wm(1k?inz}2SZT
5{3kBj)3ACeo~A_0x_:ttzndVJ@$5s>n_$t\J?3Yo..OlhOnC$|[6G!hSM[g/7{:+K_i%U$WgsK/$h9Lmc[75bl$z4w9m]>*aLUJ_BQk>:Ku2O	B!;Eg?;RS(8N20,A^ncqF	mDyRANcOr/);THAqI0h$Xx!)h,`NT#cHe[!xHIq2!b<3KL@4r{hB.s?Udh+<!Q'uyp}FFoN"GruV0'Zu'9RifdY@tdg{Qc"&@bBRWy/VCNw9z=^{)or$;4!hXvum^Obg 5!<&}uf3,[}{}e.a|	wo4IWc<)'G/NkNh8qC
H/*E~In<	S0eq'jwm*HqJYk>vt:VKmWWDZ%FJ(%eO[Z{
JO~I5("#-YEEI?GiYEZG?<UrbhErKXEV ~mLLxN$L|tbJ|r{e0f`RFZ75<0K<^*UIqs&dUE274Qf&f?k_<\/hx(9}p|F{]W=n7,Pi^s::|wO<'~N;xK"x0iP>;~W(,5;bv9*3k~OWTB%vD)+!d4)8KGaV<xSs6{C01;MGW,Zc?yQ"Y4hsGFn#>QM^vk1p7JRyz6*Eh\vE{0mDp:m#5b~)W?xo*Xp:<0+-Bj
}R%i*][kE$jG0Eh7T!M*~03{gDN8;~gj	Zu$$GAQ2sPX;Vlih]"g*A&z8;.bo3!tms?%lm M&.qg/b<- #tzoKk83m-`YX.kh|9y^ pL
~64G
D.(V2
$%]kedHhEFu\S1R"XX[UcUs_~a?R$;--H;7BeCP^Lq&Zs7ByPh\93Nv7%Eaz|pb)$/D<V[kkzZp[$*SEbXL(FS@Xth(&2 .sI=](,$EU{>h<8~7#[.\Do+%8-, Po3i	SSB?6Lx`o(|SVU65UFB|iYS
	F fcEb!-.&U#_K?6^: f-+AI iz+D'^)E.`RgZpj7+>
S<%q#..WURZ/@?CCrs#V,2D}Sj?.`cnK)`U}%#[sQ]b,*t0pLatvT=2FoDA!x98v+fhIGz7
Zk1X
/tKjSI(^?6k;dQ"Tt*JOgzPlv5l]E;y;;_o(2\8d^\I*S0}$.$b.N!?]za]B>~PqJHea;c#Ur8odDw-&;J*A,_H~Lu>T(Yf*N!qwDJ+vhSY^}(QUn)z~;h7l?WRg\Xs6Z)NK\Z*!49xJeV`9&&3C^~3wXEuDD?Q),Z[$sfTAK?p7#a/:>c8MymO$x:rtskDmOmp:f{:g7j#~6Q9q&	v^ >?qF2K>PxcZ*+Yh1l<ag/}"-rbt6W-fVGzL(X+-wT<t$R7Wh^y'/%_"R7pVr`/F0<wQ]D1\UG*H0n!wGvk?*	X%!p8V"&u>I,/z?!IwO8&"Ol2lWeS6ZU~\aP@kc&znU:w\&<^8pPxP.#5bXb-c	qjKV?\>dV%||v8rX:Yv1#<kpQIQNuZuw#3xu0IE$Ly64./fR:O@pIwK?#\||_>0wq	tCWqeR5K/uKUR$x`X1-3DE1 6`P[7H\\B9O+irWiE`_q)>ugaP<%LYQ('h[OC{0|YR3B:@\a>ZxAjKW26!ub

n"T[KNo7O$8='%]W}Vp9	?06>6E{4DABx_N4(@C
eksOi:Isy<"cE$*SG&BZG<zPiVAk]od@`C|M5
m0WgyV,p>BW;WDXb>4puMCr9N|m`'U427[Db%Q C0#lo3id`2bJ@,kKFQ!=5NiHu	~H4KZC8c@40%]7+[	xA	1t'^$ KG_RvZ"5^`p'alDbQ$&(wV#YlC MV(eeq>~h9h<nG]veJDB Yl#[`#iMJ3=Hs Lx((.5n<#HSCPHoESZsWk?Fh."|?F7T2x'kR4eab@zu>+?wp8^OO;'QM
H_	eVSiE[M)VA1]qF}H>BJz)4WyrB>Bs>7CJ-CK	mCUaB~[#R9o,%%AMw:}E^f0IW`_r=S?_=:PY?y%BWR($"2=>`3*oQoS:[iRTUg4p`r][R<MMGYZc1-!yg0Bf,3ce/Evz!"*
yf	xEIF]$9f:6h}(rSrAl!^^Qo`Iy8?^F#=P9i!=[{PU]O6bLZ0n,Z]`0F,Qy00j6A2;kQ_#tXrDjt+-S[lzvR->YM5,?GLMl"bR*sRnz'n[eG:Z6`l4EfepF~GfEAvOjPO
vA--Bz7W>>Ag^d3J)\)hnJ}'"6d_" 9~;X'8KV_"0LBX<M>RF}9$_>efg/~mEM+u&gKA!3*[1[=Qh:'e#.`_a}oyF4`Y9	{?H!T:!]Zj@lHh)%8bl@M-VH>)vx=Zh^,^h9
L!C5w;E0dr]mXUH=\C&WFNcR'V#nXEkc	GlFWb>^;\5tg52|P)4)mm;B:)M$NKLMotTL-}E?Ok`6ahUM|1CHA8rgeK9>k'Jl.J?Yh\Q4=Tsc}&!mye-h)%t+V_7I!fYmP)2.B\Z6;kN\yQU"zV#^Z6`$'9qR+j#>--fJf5`0aWKg.Y2)[K:%^n9Th_W48y_/e&,TA"k!d[goQb%uWbhZe<<J`*@1BeoZt2HTh!/VZV)MiQ1y`p)uYp(3m)_S!&3m[GV@_./ZlHy4j-|B:isHn*?IdMjvPyI4GM8])&H-)D~t6@+
K3DQKo86{a\]lWVF94l~YR:^mx)K(:ve0F}6uwC
li(Wk,"rr}k<~ovi<hD7Y!GYCthesA^$%Cto'I|
f^z\O*\UP<N+Ny	9x{8lqMNG(_4+yaryMe2Z@adQ?.QN"TWU0I9.2]r91A2}B.7JxN-F)>@5<YG}XCm[uIpU3axFY7}?4jyU{D2GkgH_8<yIVc\]1(!9<v!mS$h"R	D;X{.+h|g|wL]KB^<_hOlbD+GV`]MjP^DnM<>C@ViD~N{Og8W2V4^DKw1[^(3!>cSA\|_C~^|f"%XM~&FQf^J+4Q@[!# _o+c's}	6<V<l96@f'(ZV2W..>MHfo4MSBLsh8qT	_*Haw4'=7w^[.q&o(G@~bWf[S(W;l%RdDxcsXwRA'\8qKu:6QA>g= ~~
ev.My{80ro*e2E:8dU;n\FD~\HKW*KNrWQ0=oj^!bg>W:T?h{HwFZ#7~Sv-}k>){glmKC]-:AJ-CTN
s&S:Y huv|}S#&Y"n5!(\EM
G$U|e&z)w_*/?YC	\[TZ9rc=S7J9'(\.Jc$tXV6w
MydSOUkmrqIS9;mlZS|C+u*x]B|V)vN@rrvMA(D_fhX>)Wx/g8DFLgR62-X)"IRtJuEC;npg}
C(m)
:P0P#DhTzEOyM~>roFU)#DLw?Z$Z/R% c5K$/Mu@{<":m=1.A*gL{mLRC%[a8J.Nx.c4H|H4nwqI$2pwDtq/F5]qT}O&]1/x|.\";3O7h/~<w1m-[2BCFvFFlOPPB~F4q$Z3(>btF<DP?8aSx~6gi]C@^w|zIGqv*(%.ca6FLvzN;uMnZ{nZRiqv:K{^Gs2_ey`S(h/|;z-p2YQFILYTTP?xif9.BW9,CuEJ0Tz@V& #&^b*UpUPoMP^[[Y^:>OQI&~?*YGb[9h-L>uRRz7&QMc z-(#2*ftE"V;Pn&([0HL]|J^|p$9J"M!F6G\-P1TjCV>#:wAKE/k`+K&w=:xO=.JyAJ62-!R5G30)\+p_L748SADSmM,)F7
Dp@O/U5;)X{!;'[G6\"U7=GgdV+$0m{{^+wE-1{?6RC>wPa@::s:D2DA>HfdT%s{+z?2agZpJyGR~f3g{H&d}N[2hF?4$tM=UvtVPWR_Y!#o38#')`~TNXk5]>!&Xa/jPe0cJO/'1XaHo
9xNR399rtfC)	}1i://r$Kk_1@A#3'jO,,.N:'7{@R}brqB{{9oN~*<		oAdkfO{44Z2ufn1]|ViqU_czM]wOuPac\~9|Oa-@lS[lV4gl/>X=7]FiDY-EN5u#D1y?Vi`2iC8rCUWkMmFb@h^zWA6o;y:34Um *Zf8{<XVihyIb&BTqUoI]?X`48;ZpdWX2CG&oi{1R*V{rg*3<5$BVhSOe	)Qd4p2AD$	J*BP(jl~;e.M=Y#YC90gSYj*%NjM.	+4Dw]R16a{d2`Ax`x(	=?k/[	TCk<,SQ-.[C;R}[N|V[wZ-8^Nnr|XoMdHu"Z%#^6>V/|>>.:nkkEwt42A,d4D>v{F;j//E)e(s(\zj1$!*+93
QC'E
91{+]iv[I%ea:z9P+*-}+E3.D-{t5kh?8(A!kx2rg/J}	v*	,|>d|MG8=eB,_w=Heb^\+0-CgCNdic?n*
# hh3j#-D`EE;X<A7O}Gi'jo{~e.?;`+84:xkrEhc.6XF14,B}uxT9~#a3F2u}aKT}p,>/m	sP}35<X_ N*(a	zzC8t4z~ Uj[J~-gKgvOb~	_:T>?Xf\/h+bg[[2%?uq7\8*yz_s8:#9MUGcBQOf0V5vBrXI-p|B@*e837)Z*g6'Xp)O!cJJaJ3hT=WY:r}mVLL[LD>e<"cKgA#txra\v+B|skK	Up{h2	ZF,I>6|(XA),`\E[[;.7R% f=j7E0K]B`.a
G-f_NSsAro6i95N_GOI
?kbg/dSo5lIOCt2`1*4#"kTsgbMh-${)Jp[V ss/c8y;6E{6)#'0'vqw|_\k+(cEO$Fp{(Iw1$"_AAC _Pmm4/p$qvazkKX?7R0Q\d7R\{3:g\#g1M]fqvX\hNLT}%8>.0="r!Ma[7O](K^:U
`0lu<&mEGh'fl&YUTYUTVMs
O3Xa2.snn!bpL)s4+Roy;_fFX`>xyO'QaSvyWCS5<	8oNe=H'c%5;m$x?S7{:X$CEU~Jt*}VB+yx86C]w0~"KAq(uA8?+&szT&M<'a)r)=%|	'B\4@n46:x>w2'B>Be{,9xplK))?L^kG)E\[5f/G05n$(]OFF&vp'AmLVWg*1d-bWgvMkLa|%]1s|
{np#t<)`g5B3 f+9L|8%{FZiyCS|>ZG]MRMxz[u TxY`17D=gD?|es@,YjLT,^^]/ZZCiskC"Hy>V6>dWznfK%pp`%zUG=2u7u?!a~,;$GI!+lN'.?<]<xXCojU3NaNxdAsO
_MeQdYBlnpAX90:#fd!1U8|eJu')=T=,lv+H?	yNE`?2c{lV%W[K1@p)9zcYPG+4o4n%s#Bq>V(}G2.Sd!	B#z;ZYEd&3a."8F/^Qf#s4Lp
l\.r:H)+;?,(Rni}B)5g\k4oCs/D 0uQj9X%"i+Tu4&mqu/Sc.3}=M<=E}bXT`ver'@;	;rfIp@?$80BpJ~`*.	
bJOtqRl[	@}9dC%}3RjH?F:7ca{#sI -?71$
8UqE^XSB;Zq\K_Z}M\Cy!P	N2-6hl#[0CyO%YXhhzeQLDh=LD~l@04py0'@:GW6F	s8J"O/q=0C2LYm|8XjBLDm-cTOX7I)+*{Ph;-;MKTxQGK(FJ,U'a]>viK[
vx.n1KE~z*-[-bDJ-URq)z-:UscTC9mIPq1Jta2]*+Bls`=KYK}Ay=&pv}5 ;y9)ukDJ8d~o0"YfVvrTbaS?"Y&RBWo?m)l[2rp;?V1ZqXiuU~n8L;jO*.F2/jf	,+HT+K58dBk,,-/!zpm^ywBs@0._ 
wY;G;4$Ff)^u}o+5[efX-2z[my9vq&.]DeFzN_nHl][c4Z:^J\q#jHLVo.n;05`cE_d)uUX*Um"<AiD[6+)T
}Q8CAB~S*N,.uW82HO4DPUk?Me*]Pu]o%Y]EM9W}
g<l9	y^O-db; ZUo>>/D=;Q@82ji+>3rc&jS)M1t_:#75m|eeEaXymjaw6BZbLcXTwX,f	tu;iF|,\{mcW#6&i6/L{rU;_tB&p=o)h{D5\P-Z!-sAQ|6<h?,7RV [dOe3bucUhPJd&WcqAnX;:#
nSgEqXa9ASI~p#3m[}n{&o/D3OCL*e'G8VUDj*Sctv;QUO#J-1bsG}XYw&l67<N$kc!<9j7/rH`+XQLfkX=>?ds(2xOU`A@d:N>"d(J!j, ]G.vf8
_jWG^:4@%a,6$@8_kxL6A/nvu6JCi[CAm;["h'8'~;rH27dgx3[0mNf$PA;L`b*o\(XS}Qac/CHyxPC_YEXWYP bs$	Mm!I0gkzN)a)MrT_w.;aVqGN	1{  S>%$0NsBsQ4$SuE$Rsx57QnmHlJgr>PfK$``Z6C[ShB:"
a4{=BM?h(8GGw}"wVWB{sl,T9z;K6;=e}\X2y*TR).jC!m<fK%Lf+{d6AI=F8@
BBAQ|zcZd(|Z*Sl5_];@DvcLlYR_+(0kEE	1q
$d?AhSaX&_0Hrl`1M%[Cmr^kVjj]b}h$@?R*l( b>vwm{UE) "Ld"T8#J4 dG`Xyzc|bOf<	g-dt6u6;A^'gFA5>CaXdEPw#z2
*Sl,|V	w9?]2RK,:RID% \M-!r63Peq#Q?;hO;S6AG86&C	MWD=XJ|ARi0\*|S<Qe3<k^O4+f]XUn8/v:c(Z[cCi@m@tI5?MB	,)Utt?ikmYZYCv@1xyr}Q:Lv#Y]*/Jgy9cBHW}@)Fx<!j5G)IeFARL^k#-J&=Qf2'Cq?vLc
m'Zf9io~K$V`SK0n0dmd
1s/_M}4+]weqwvJWOFaqyMw@%a{ZjeJ=j*
LDCL:,S.R^\[`3%$umB6FbylFjzbk8}V41yQtUyXpFnCU-=g0EHJ7$	e!`qlD0U	}w5V,,@1zIwO|,jEOoRN.8g?_(nE
b	pW7\ms0/?f")m>"c	8nR2DMA$[.XXtvM:dPU
eC\gD{/8x#qp(m?`Ul>xA!=u@#KwJqs.gJs?WaM<O[$08]V`c>^_
]x,#3bW%qD##?(yW,E$X#cT,Osi]yp21)YG/dp*KUo1$y&K)?#jQvJ[=-41wT?_
X!YEUA%RM+b4F0hT/RGH55O]*|NMs6?mLc(|za;^XK2R?}kgv!U|S)+ZV0tZ3Q/>i/F]Kj]+uiMibMVSv$KdN}!_qxK8%hq./l_nGncB.B;JDSDF]1n|ojtH+8'$@3`[l_W~TC,5j42>Xs|g0vuYA+>K$%I}-%O:b#D[*=5\8>o{N^w@oq^,|6	?XXHo(<NVD-qNg/<|8>8v:"L^TB<gz:3Xxv  .'w=$c\4k`WaGc <S'@wuysO	02qq7LL;&^W~InTe8PNYV|S7L|