x`d}c= 0LY	uu1#{<QJH3~QL^lZYJ}SH^:h's`S,yPG}3#O#z~
WSb:k0zgsE!euhGmDgJ~"Qha!1iS5!f1_\z.gRQl2;V,PQ{eh.@"bs6H_%1hD|j}kpB,99_Ld93dB"!7wgts#$f%@Z:V:X1KR>`4
<MUPoxI}9$]hkuon 2xOlp8teGJ'{CNIbOXC+^?Ww&9?hX`1.LmvtPXK#L d.}0Qc<&S=Og8>wPWkD_aMii).T*$]<N	L&,AchbkBL41"8--;|}$dCUG)wxZ>4rX5Zo[/,B0h$T_g^[k;a$GEYqf}M'c<wAjg(=D8&0)1CUB.+5jMw4'Hb8\Dzqk$rZW3[vn<M&(*LlgO{FI`|EpAzYz	'cA[_||C1+4o)C~34xN&DeC^%dp[j[44B`a,m:hs)MgD\|]`}AV8=s]qLiPay1r^yZD{(,>0M6@K#h$(19ArlS0wr:ov{Zn1#4/`h8|n.;]cP"4|	<jiU2Fxx
hqJa7-<W`9G7!fZ^)>T`v4a.g|z?b?nSivt2!FP0Ir?9;<At?/2WmG{sub>sFt?jgYDZhiRO>p}.'~C`HlBaB`vvZ	d2Jeicy6*ac|x5e/?neC<~|ad1oQg{2{VH\8{AOB'a_[#HIbT1h}6j&3Z5rW[um2Y?(`=bR!Ew=S]3wT%3%3<%f;ZI-
:Y1rTybW:+/6uT9#rOzr@|7x6XAVJ2N9Yj0_Ic1|kp}0OX_PyD+`$nm1|(+$;X+Qj/*#T|lAjb2K4m)<_*q	:Y.g
ab=\YC#9$Y!-#pNG(: pt@b[H\id#=5lyJl~z\p4<BUq$*zF|t)q-{`*F_kBUT -H_I=
N`A\s'9W~h=+U{t8D)	v]9V	g[8|;jf<Zh=uAy#GOa9HbK<ZM@2XQiybW5x]jNaqf36+q*0N?%GY\;gH*<c;4v!V3ats;,1)C<e$gN'2P~-!;U/OND}Ug%{'M3
|6,:>8I^Ty919E=QKx}V/jI;XNY>_D$fyqQ="[Bd.y1X cd>e"cUYeEexD%^(&[wKsA0l@YpK9Q8(*kf2Ef		xkGhRt2>Eq<J\uJW'T3GM-L'ZXkU`!7{jUb3BAkdRZ4=LMp72O|y9)rTmh5(NQG7yPA!f?OnEPzINws@{oB!+Yr<''\gO]=p*tV33.Dx{D{m @WWJT/ZGXCM8qbYCn/AsJXiFm^dF'{\{l,Y>ilz{idWYN\3fV_sJQu9xeth}j<.L*\n(onS3GKH\@x<S<5*")gBF
$%r5qd;V_=v0LEyG7E2$MsDO$VYtH-2fjuAZ5?.%v\QB_q.AjomUH!>}	i(\W /j`J	NSA~Wmk~sN0
WZiD_@R.gOnGM,3V/]t#Q(fD_*QIpsbT
(r{eb;9[S04@Q2
bXEX6FK \.,
O? !}{xpsh`-{![P_>}bHN#gC_dTzF=(STAg<b&DIpT:fI'Dr7,sSa_})S@c4~{ULwZ.vWpni_{|ZeQ)</GM,c5KSz[QlJ~/"5c*
B>/YjG;?4go-?ga#5Ej1y$nyaVG@bgL)/1pwH&aRzb4?_y)o&,2CT	6Bg>@^+Q)4Nx&x	\?1	3Fr)iQ:l#n#G^n?`d>=92J`2}yZ#k"X-&g9?=2R*1o(c~ZLUR'`+E04($'Eq|O?x,4<m,P
F: &{Iu^(lPvs	f;Rqufb=}0XB@IH!A8zf?fPU`=i8u#tV%5Km[;D^?5kMNEA.VDG@(|t#aM"U0n$8/%t@@jqlVDv^mpClnkNDa.4{b0V+a.L,[_.b'e+DzYSlJ'!BJkb#7Z_Pj@%"!g[T{FmH> 2:Q0^bt9hczaquJrokA~-YD;O7QOs9
{nx>
N3#^^FjHoLa"r@reM_>)PQj	3]{.J;'=Y_*yn+k*d\j4Fm*o7v@?a-=q|q-~[WC}W%.jdM8`]Z\R%`SnV^)\I@!>3$=DChw_?ZrbMc%h#2~osV:gaYy)>(Xs=B779spD^KfTj\*2uM9z<B;NrW,c?"V(3sZbAEKzg,nyP<b#Z2UPVyea<Yb3Ni	|*!wj7SX`$uxtt'Kpr@CWP)>+o
Tl)UbilRQb9Be:P%Og@ca$}fm{3QFZ)a}'E}dKQCB% KqB5^oSk5){#0Nq|5~kgaB1Kn6 h-X'fr%k+u3BXK;5$wrc^R3"<'{XWpon:~LdjVN\oGO-Y,wEXB|s%?AxJg*}-_`XB[x$m_0i_]&-<-n?krf'`\Vt[!L{kNf@htM\-^tFX_Q
#O`]prw$T-\>Q T;Z;{C?-*=mzi7w-fr8d]izNP2GhXW}D3cwUd-tuN-w(5@~CPn>8x;5Xv#AWQ%t1pVj{l07$[z!@6Yby|80v"t3@vc<$]^y]t.x'kT]
>N
/oS
E0hBAjS;E~Fhaek<6@P>?Jg}fb[UrYC}oJp5T=3|#:);b1S`_0oi3'Cc~lp,{j.*v&%K#9,>T/_|CO?o{T~,)}[}`4PPy7G,EV=dDz/!cJHb*X'+h{+jW\s0sz88ve.Fcny_`k-''z@LnON8:FTMs,d!f~Wuw~^ARP>zA2<QC48Xj=oS;pxmlpFr(*:'puM*"T;AJ=YK88X%IY5>v!W'8K,ZT}&]=R" r!.a]k?ntM (%w[k{t	\QV~Q(gA+T6%H6vz\AW|RS&X}OajIzE1+7ves)vS7<m?D~si2=#_[uF|a5+fO!As?;o]x&u{K~y9A5#aTIP0rvT`[T8;m`rKN%>ee8!MX!Cln{(Xb?o4S<t%	CTQaUX7QbL[zE"lUQBu)t15C|lA77PL!?+$NV533@(JLJEXF'&.=|&XOc6d^\;p|>|8 N3h'1ZJz;_\n!|a0JXb,2sF(q
zrII
	U$OusA9:R&2((W1{En?|e(62m[{;A5D@r]j_G.ztjGAZ@,DGI!5I>bUE)fe<tJ9E=3Ki{#9Nr
HC*f]X_u*epG6-w,7"vs1O2-p)/7IZ*BZrJ.$\a>&?!{xMXLtf,:8RW6]|7Jv-D&()w02{ALdY^]<e5=\?iHqnXp G,.}khA90^Dge.~n2sujsU	Nmf|?Sm@}]UH"KG,F{|#volrWEur{^C*jWe\Xk86i7mU=Q4E"sKs<VR?jiu iC	|?f%	%q0twiv_8{[:telSU1GNK,e	6+d
hu;@ek~s_[vnQ-}mR*~Bs+]1P}u]Vq+K&u_lb,/t~{C
1V=g'dl6c(qQKD}[y)oJDO.jvZP^A){9vo} QoR|Wot`Z|T_=1Fw-5V}<IThh)QcD	GN+C1
5=[1JgPkt	O##u,r6e_0	^BJyk#$K6UL7.	#Ci4:]*G]ycLtw|#ax{[[mVf3J(!BNm(NTS1/jH+~Dc<u_C,	`-)"h:nbv
-}4T}O)W9Vm>C`]+:Pd~8|Q8t9~	OYF=9RC!<?]9-ku#7U9#;	!(!9BG-3JkyG/h;1@cc 0$7H.V3AX}.l~-r/ms;d8%2'[s?bYu90V<|f9{KShk&/gRgnuN]FpbLT)a	x+Z	':jIhop,@E{mU'kWs7BOI#+G	N}:,$M{yEi6S&-KZZx^SvDqprJ*e0Uozt|zZ1uNZvM"$|j4Mu_Qe9n$3Xk;t`y\igNxd_wqTn.	-cxTzPDCg9Ob4P:gSiM"^.-]}Og1ZJ\X~^NLSM"$&clZXV^Nxmw=GRVD&mq!:wBRyw"_zq,'*GH; "LX@MHD-|Rk;4'F#CXzvdMX(>PGp[6!EWlDJ>B@fBH=I~^%8e\;g!z[wi;$cTW}@ FoDsR;__%@Z(p*	7{'^oCtQ?1?mX[kA(Zjz',=^T}(oR~qA(bCYR5:Fn]Drfo`=-5
})oXY"t*1~12aSw:+f
?m77f;(FfJ]C*~X}7kL3mZ"-fyd(pbyTtm$jL=`lZ%2}2Mb#DC-/qrsu(IwjvLN)a^q; L(Z%t3\:Rg/Pf)1s,,3O`vsc;@-k/li&J#x18>y:RKfx\2VS~]m~P$g\_>d%+Z"[RFH+-D2ufPpL5zzeJ)&'G<,ndZojJ!ObUmym*Fe`yZ*wh<;%S%8`IGx,FsjUA@y0T<QTP<-)o%|tu
*Y']}+QSo0q/*eNoX~&Hn\M1vMPCC}4jXD5Y9XGJO|9j8WgR.J)R |dHfa)3WTc$&)elx67GK~_}~`HJ i5I4X2V0({t9?/3jw.f~BR/.Wan>5U(El?1LhUW[9'|A2l&M.r.O$Ub^0N]Tug|v~,92U$y}WHIf:TvL\3%vPlm.V)[c#pZdC	ve/HS'U-p	N]	nrQgqdt1H&tfpU5Rn?Wd_37m~]VfW!=_775q}8J`l)0q-v#(s!zw|Az?J)N:5!WlVaBlf@8g.j?gd0	5\5;(tp?vjkv$SBO\"nOJGQ'hqyIUK|Q?Z$J< xwL>@tWN_Bf(q4\(P'^\xDAV1v,a35p/M=I[I`66+XJ$nUO,{I[^d^]mm{:~{RS-;Rb(8%V[B6y|	gFF(&`<FA_Wc4;$$yh1^l1]&hJ>p\#%lS+70GoZ5S>7Ez\?VO/)Ap9{843DG@_^Df?E2V;Vn	RF}>=JE0"R
j-$d(`V<18]1-d@Oq%%27XoI:3K}3To^eo4>{2'm?K.%S(a|wPer">rp;	}MmFH4QS1&Z-#1+a-KfmvAT7.3g{Ux'Vwvw"J#:%t\/y=_hjDPOChEmtMf%S1^]@
'`8,H}`>misX-,>|H
*jp?7#6\	INNBF-Fv#?_#e\vH9T@>T^@2*3*Ys5hEl<pLEYH>m#,#XpP2 6<$wO(bwKnCh-)JIw3#Z79Z[ucG0'm K&LDXSr}O':c/r&r!	*V-9_&cKlLcKq#b'4q&0P[G&7iw$md`K^S\&)f|h;U
hms4,pMPYO]&}]@`E:q=gZcWdb9[q-XvhxoSg=P-[*?TyR<Yso1[u7mUjTw1AxRi5[Z1$}bo<C3p~eW?TF "5~Il*vuquEs%x{S3V30pz~PDb!TW5{X5CvIh5hD/4%Y6"Q[F,54c?u	8q>u#}IS;ag8+C;C`H[NYD/~=fb@.NKmJ
A\N{(jl>?4I)CA0))=E*^bA@pn51[E1W.1fE"?N#Wa>^)*i\U?c;P7tYwrw-d`hax<? S&yI,&&yU+TWTVnE8B( cl,R8dMXKE_dz=aMpDS~='J@.^xEM)_%o:*PRs.m\D
I9.-To_6{=?#DS~B
JXmu<A/	A$5b
!1&uj+Wd%n*(<dv.h)ro_#3;3@evaks^O.Te|h	P_<6XV19H[lYR4	2%P,	Rm6U]7?U^3[!J)]fS6yz^}/aI"C#KNDd(#ZEJ1AhH4U`(MA]*?7n]4QCs	vUMl	wS*YzvFtnXwzjA_=zYNw7n0>nbu*b/<-*]}l=MZrVttZp-x(s*"~<Hs9FkwG-nWh{d}toB52mh
iO\M}>s`%*C`I,z,rMZ:4r*.tw4i=XgzAHe0{.Rq5{S2wKW$s8K|b[w25pv!<2b4HL(!!TZ06Ogw/ F~W(T"{Wv_9*$V8_!AG6R3JH	|*AQ9yCF\AG!kw	.zyBOa/6}@oF>[
ZWFS/O}rieEl'a^{l._c:{Ia/jxh6i42.nVO?c~>Byd@STf?+Q_gbe0t\YFo>P+N*fVigCKFjjTc>Z6f	pgB,zF>wWWB"[fa69J5s$FV}HTi/Z1[-~41P)7A2^3=o8rUP=Uafb"P$H@bt-Caw}%7Q&L@T Dm2Y(%BV>sIo#	Oq\`F:r&0!~	eyLI\hU-rYC:7V8)+6rIBT)X0\%[KhOsk!aeW`KK{.aC1vnn!C&(kP3Z eC9jF8aPzi'ls*01+rsbtIVi;}
U7f+acnud37:'[&*`sr<^{GEg{yPDybd5 W2<BG^Z*_7$f^P*|B-oG]vrFS_vm(t4jn|LJZ(qlM.pa?|JZlCnhAz}BUMiA-:
g/f[0%:Fr]8VK_FQLj0HAYmak8&`YfQb*l%UgYC{YDWe@LC6LG$$vqsar%sG;|spe)X?xfhsig-Mh#W1^O|Ie(Bvm^lz4e?lX7>]G?	1w(@v;m.DaogU2Z3QX uahx..>ir|I>G,7]=K=Hle-tfi|H\nF@DK.5z%A$a`%s]n6D|8Yg="OL>^UIwxnX//E7UVx"q@CPs<_(,&4W*E'<M%Ni(ev6lbbbIvV|^1 /HNvc-*0:XnVQg*PznyM6K3Fk0$3@N`!_.Qo_XLW)-m`.b $\U/x6%hX=sdP.[x<5c%:25
*V	@|EH@WNr7P;	k":F#=6L253}-;~x\aujR,/.D^[-$Uy\ot9}\*sS#r_#Dc\rLyZ(U1pCs'b@|tAYe7l$K~k[vD@*pD|bIaRO$lQqA";s9X7NYu,}-fr@LbJ[gn 3G)8d,|L`W-H5\	C<[\<+T%m[aM)Rd~wY02cL]t;(}/,^
b~r$sdIi_=\^49Dg%TS75vZIOD[62Mr	CQ0]e$p=%pB$',y+M,{]qoM,1sc[09%A{xKh3xk/xafdNy=6tiLmgcAe`G%#`dJacGHqA1)|oDf^
Z0f0{; _?/H^jG jKD6!PiqBetk3j[GulhVh8%T-KlS"3LMKhb|,97[`246 ]7X: 7JIpibPz9J=pk
T)S@uUOulE)r"9=dn$T4B4qU."q-#rS"")@*Ys5wX!-2fTkNW'J$"ZP${nXNb&ods2N
RRbl[lsg<yg+#[!<?F#)lN<|`M#W(`pcL-YK6Sm!"jh4O@~L/aY2qAAgkB()yKjL&10>xaB)a`$1+kXQi7++,^Uy UIY>F08%Fgu#iK-I+e1	z'S=))M8chRw:K#}7|8:Zd~Yg}YYUz9P.0qw@GaUcy& C?ETLU@(Qb
25
cTAn^W#b- %!%*{[QN}cUH/Nzv<jlF)Fv\+@iA-Knj'K	"-J5A)ySiuyLdX%hym:Yke$K)@~+c!zxH=&@??XXHl90D#J;,bP[_jQ(%j*4&z"k:rfY3\Pv==@ZGsKomw-;^aXSrqht-`EKfY+FClkBM3$5qurkF>M(a([B)64-
(.Ew{UR44n9C|&><s3A>Jr?kkh--6B"tiIXEbRm~"/b@<N)E~|p q9sr3yxq=LJ%dL$&gk%G):^)P_A` I'-\5_2mcjN>7gUczaTB^p*nqkmI?5(@t1yT|:nVJQ}L[v*j6hww}S?t)a}Zu"~s	;vB!%%(0b2xbG!_F^JrRq"BwI-]Z7sR8_`B[q\'$[huN-"{7bL)Kwee=od;w~/`Y1(H L/L#%|DwwEEh*LOebhI<9Cc/$GDQ**~T-*I=SD	PY0uq{A5-x[-MvyF*o'$\qN;!e.c|}d%1EJ)f/vj@cTM83GBdiuulR|x;.zeCDa1$jW7Q$w6xZ	>B1Uv&$DAc`Wc3&"k>+%Yvu.9|Bw236	lymV>>QfZC;ZJMa:!{ofN07]E93%=}F%8>SP^htE3k+_2QdM~@H:[,	g#sMlY\EvS;#%DY1AK$`cgo}EYj	VxLx9nI{@HsP5E}/lEW`--9>$Y)=b>^"Y"-?AU	64 <FHkAq<`|zr
:Nd+>IB!fzH'dows?lQ+uE5\*
}$KaP2V0
-)F7M48E8Vb,MvezA~;rs:0|Xo>^)9E'IUf&
x<z49xMYi9Dx_wm1;l@TY?6tzLyYu;i/>L;&_T%W	pxH$B/Di}H\Tx|B#K:"*EqI5jflZop'kp^M!,&t7rK1m[YSQpmiP2hVap@#LcbpmL/ir)Lf\E\us*bqAY9r`\W 	5#l<10{mqHX/q9=@wOrWLm?:0}@
owR!?"v9+Z$'`]X"r;S>8V
t%*\$5c:<a5QnhjC.7{	2do*_}cCl@/M;}K)FX*Z-jJM [uN+5CSujm*v7d@p sc{j}Ds:F0%.pp]g?g*I^^<0#i/q45I!O%1{^~H**|8gc>ogij/kZ4i[ws7gq;&j1b,9J 7:ePzOva-8NIejb_e(Y[wu}uGn2u|ELec<
E*zWw<`D_bLU}3'GN|E@(bdmnyY)r	);R/r;N4q6v9fq@:=Y)bg MwhwAJ])37E?!>7fvdN~l_~H=f@tHt1*s8QfoRq581?D#Mg%rC'JKDyeq-@EKJ!IyE$	M)}qbv``(ZXg&|"01N!v-]xBIDl@bIw~6UU%KotDLTi;c[KSp,lvwtl<1	@vcnvG6E`/Gov|qN*)W<BH*M{=YsuVPjH,bEaxEXBLEjxU?U80z!pR8e>p6h'~?ajvlCSSmC?o'P
2+)z_TG5E){#(3RvpyiLv&3b7o+vuFH#x6J|#[Wrf{UchqWZ@Sj6O#$Suo'gUc"5]&RkipGTv{@@j@;VkzyWn/8g"o:zF!
)KYvu*	).PG"N%M+?.)OH5|>;]zOcriW(/'F0GsG4'
ge:Wl`O@)V|_n{hf}XS#:Fmv&AhmiCUMCKJB9!O+'RUL6fYr(,t&~:1{v4@@Q3h:Q7tUy3jx:WQC'.c;@"VG*PWYI^p>C=E+k:CIESH/l-&H&sz%QwbRv/#/]g+f|>;kDTmY}pD+.%"?q5vbr94LBD]=7Vyp2VN~T9|I3nRyimjq0i@Y|YI
$esg#5M>Dh>K@}K>S4nP{`J
m8,4ZxD]<5y?>2MjxQ1W$T}{5(6PD/)'_4\uazq~B~3c{ggUZDZ@=v}DtBR@^RX3Udj"F~uveXiUhud
*Mv|wqd*>x{3CIVZfTrGH2>&nqxnpS%s	4u}y'UCp*=s{baz^GS|+yH0)!%Ov-C=]xTVPTs6-M{EOGE"Py_>g?U1m;_WhI#S4cch@fIf*:?*~V{0\DKLF	T$2dkLK@6zFt:33d
k^SNO *R3hpY@!C/lQAHnCtdH	CV/;uPG?a1mdfGD2.,gn1d=!VmMt_?}?XRTa$9)&\eY"yWSk9HpVPpVWF5d@ID7-|rW_r,|DLEl<uDbWf]n5r.^C51>O[l[t:CW@EYL^ 7c3|epV j$8=YH{|caXkho~5Qk6oA0.`+hKzq%Obl(U*E^'0|4Q:81%R4,.0]_JH1P?e^=nL8Ypq[\??oxfH	[eu,4\?DNzq9&{fPT!wkLJIg!s0YL.$.'4TA4"m@nJasw~Eu	;(Wj6.IY*Xc:46s`U7w37F4*Vbx|fDVc<4<UcS\ND@aCL0zEToPXu]7i{+Dh9'hZkyA:aaK|Mv5>N9D)|+Ivd8F;h#-f%ZOuMNuTxRWxq3wqy\
5RUv]'atj&U{rkb(yau,OR5.%qw,ler-BIG
[{]bbZd ~J/a0)7C]ZgCl2Jt";3&D0Jo=#x>lr_Dm:RCPZk9/k*vIU~[n(
AkZvXGL6Z v?5{8%d-m<P4EM\/uXzXW8Wkenb%rUW0R9+[6@*K	-<QA
ErOD97*?=,/RJ8p.2!OJ^V	pV+*iZ;o{M?Kz{"#>;;"o$8?~d"[2	l:@CJ{XVnDJr!$/YSE?T88RF"9tJ+25m IqIoIl|Dl[yF|8,pg+HFZ.+.nS`[:M.WT(=U+26V]);b$G:hAe{UEP=fXr7gl:0-.v6Q_?'`8Jjv2*A]_3l.kUw?;\W(h&g}``7vpON2CgS0[WD5OXJ3tl5to7BRtnp[6S&Rhc<pDTu"ufD1eh?a5GdA_8Gi`W!^5a]Df gEeY:~<DP	mrszy2o+=\'Gz~K"v['WG>zPSlE)iL
nG<!XEz?5#lqHFY[EkKNEn@"sh\+~/}%g:wy\Q6I4Xij)_owTNNp~'PGX$Y*8<elc5{rMFU|[+Wmwg+nZW-T!$Gl)cy1v+gn1yO_9MXa+E{*b3=BM)Gy6,e9P%N!Fv1MuIy[ xF2?6Jz1f*=ddO7Hj!rddM^nZ}&QvR%Ad<iUBdZX?.3z"DktZC:x,nts1	hnHqsgB}H4SeX:2&
C!nO,lGxHa #1/ijh58H?Z]!j!h(%,'\K1?<ZT^@F!&KM-RqgdVE!	 Gf]<.=07 yWXoUN,: 6;TW%@j	:H7fOK8kuXVv#+T+e`cx$
*}	v5r6s:2w;Co$K$l+R%gVM?84Dlhb`8d!<Lhc]halzH~:;N*E#l]3V	cPLV_ XkFiu7gvSe3@H;?QpD)Us9K#`1|n!	ZuRT*&8SuS"vH9a^K{4
kjq^)0v-3WSTTp9XR)~*@h$Y=#Lj
:sK;MQ,>.`cXNW.w[X|OOq:>YL6Oxy4>v`2\~\j4%B$%p@_g(MxPf635OG4SS~}n:|.ecy5v^xW'k<oE^ND?G%QIg%bp
24GD8#[s7iLv^)rwXHibR/:ipeJs |.Zr%!$S89T1@^I#In[=6x^&",o@4qBk'|sXOkh%&Hj:hfiLu[
,-`{(XDLpoA G2*-gO~ISQf3*wwar1m*(\@i+@}<Jst>Ah+N z0k>e8U/?C%%7qA"^{IU2RB>L
2XDD09h
)m ,29sS"S\B<wyI'_g7,^ZOXTf8aP%UFk;EMZ;Nmv_@xq0^l!}HFaO0">oL\9$X\I-*(ZL96:xkU&@<Ue.StK]zid8,m~zDD%eylpe+,A<Ub(1.>&y-{Pj !b
=zyW*+(?k1g[1")_I"5|Y(vl0:d$Ko;7JQ'lkL7g)l)jkBUwF9:RoIS{{/	sxvgN9"E2'a"ebTYsW
q ,2B$DxUuVgQ&$E,xMsA\C4Rf;x(zQqRF1#,pC}LM);!d4kfk_'#u-%wcWI|
ZLK!u#kPewZX\WDGv,I?GD9T#"7bz=FXt	e-JYj z[C&YA2V"Sf3M'hY<)U+P'>qsk7FrtYi0Q+?[BLwT7F$;l(}}EZuiq#@#7Zs*p_(-pc)<Bh^6\>s^m1y6RjfGg8 "W."PjHCchG;L5\,#.a)}<_o?@Rmc0gjr[qyO,
frVp"VV1*J<Gdd<J:Fb>/M.&OAd|%%v`D=Xuay/GXF&.^[OF}R-"?{el:7Q3
!vG^~i}p;;7EUTsJQIOlH-	*|R1;B"0gkh*~sL)%@5+uNWgB%jl*F	f?Kn:x	gj#S<yr=m:aOb&ZAb(g@aL^cc!t	ukz'/hFZRK1<*6=*&f+0O.=?	-7|v,#vRa3+3RwDZTSR*5:W#tlbUI'|bCx?!zIxWS:r!ety[I*6(OMy3rL	']K4vX]5u%YLAL?.`kr,3QU	2BJ,+DCy{k3Dg#S~D:UKtU='A:[% !=7vV.K\qlkq.@6r|:z[D%IRzNm&ReKk8a#W	F+H	RvBr:"u8) B}D7DurzAP\U!n"BY[G;b#pO#Lj<Yi\*-W`IgP:6BuYm$iDKhEV`K)'\<G{nVZ7'=#*H9e[n-_C8[SYa&DkGST7-o|1"\p8I( 5LXuW.`{QO7ji?OZeQ	{3[>N"t~n+T/2i,z_5Ug.cwEc[}mCzG>Laho6\#@pcmc8}!ovWU@*Zf4</:z.z^b3"$$Ft-JbSWQhgToxH\5
1X*vADkG<f5'~pE=^l1g@'<@i7.{MO9r;/~FOUh?P(u<oNR]((g.a/t,8F'mBfspiu@<7}!X?2OcG.(lE|s^A,u5cHf4bMvsn{7B-	DXqKaKk1dymr^wjy8f)<G^mUL]b,`	t-cx8H~e-*VS1h6PwYf-J,5	Wnzz?`,M5?`&FB<IfFw-g1(xD.uaBs<arq96SJ}"Qyv90:=J"-9]";?_(^Hn%f]5iR=!bT&jVYk<9`eaLkTT)s}NoywT;48j(wQdS~?E^x:?kSVK/GhKZQyy0pES4
xoMf3e`W4#Ft(}}-(/djVq<Og{Lpfs%Wz'Xn)_GVU1_&+$evgv@dl<RIYCB-m^Neqnr"	a*r0\{b|p.'k#}of4L'XFGU!qhU^**Ab)/}9u9f}	
fm0duWYVz9#%`lAcS(8}zo:)H0F#nI%rk[q8%qlKZH:fg76N=WoX}9tJ^9>O	r<
;77Dtz&-?Fqkt_Oz%@g#.lHIw}P4{(1|`9VOv9C)[,9Uv$))8PYTl)?N= |:'V#TM_|Q(4\FsGcp%^{)j''o$J(AWa>Y-yX|F?!DCr44FW\drO@?
&X1-\NwpWdT;vVdtOSW-al'i2,	(`0&hRfx8>2GCsqe$lDUmq~2/^WGY\<B!V%_KFxC_q1|]B&a~/5)8R4;:X>|!A8Fw'W|c$@54Aimo+0]#B%2TB-Y$5<HXuy"{TG_r;}]*tu&;$9ukdx.=8^n>h#%'K.+oq8dd9yA._@ }qrq7Y,g9(AE\ka]A>5Bb^Dh1+\-up$)#l_IL}_q~.n,.VMq4PJW_cIvP)|$e[$WZ,GIk]5Q7x	)U7E<
V~u]8oujHN`m-5#lEsWLoOD7D}shk!}m	},3qNW$Zr|kb8c\q+Q>I"fUq|z]_@`GUnh=J2i6$hM|gJ:OPEuScx_?t+<szs}
2_h%,BD'{!u54RWn^T4zU <Ju@!8?7wT<J)twn7v]4w//J$1P1JF)|6kB0b\MhF>Gfi:2Q-S&yzx7/H$F$|o@mEV}Dtw9sJ(NQOkIsVS!(oQ"I;=MB;BuuD|Ur%AvmQbi6pZlUdoR4fpq-JyD_:&$|Kg*##%g5<L%J*N1?
RF;2Lh2L2ontp[)]|?MH}b
6MgYn[1Nt$JEKhA=kGCQw/:";J{{gK?{W+`vRDx8%sGi[{f>8a(!&@gNn=M,LT/bw#98nsL9U'|*[_g)@'H=ux!t+2-e<E9!JfsM'G41$MWNUZe5)6~*05CLtAV&;;Mr{pxD=?`n\L:]p#R!p{,7E,5WR#%nA@L4.|Aso}uvAMGHh
CZ0^yZPaPJk<(wq[N%B(;wnw'NC:S1H=Z6:pGPxf1xB@atPV
qP;R7ECX63-UT'T&2DbN}?m*H
@-kM{Ap{rIA5ThPw	^I}OlVE7aNf+!/W7HY2MjTs;8TY
0)T I
LQ.JlquoX%bUTq#hAAn.>:fd/OL>9>],{]\$>)-<L&Ki+70c%om2=wfE{6.~1d@Zbg#1yo@n1VI#^l^bWkBGs%#cGYPxI_(f-I<<3xHE&+oN$6UL:+BFth.XER=jEKR/T)EWjB!vXVA9^4168I/~`*Q(AP>xBf-X\%)FUtQ>Cgqe<J/Yc\="V9jW00aD).FU#6?m-m)K)5eG?\WD\x>h2~PL=Cv<x5~_gUt8{6&\fi{MDqT\|4Ou?=K>JWd&o9Kem#A|X9C<gS9wX;b#x
0Up1EESB<b[	U!e<Fi$s%ag~a6%yE9>K	A6GA5S?!X>:/0/p}';*Fh:,:ja>2 rbj3&<,>bKV`McnF__t'g{7wIum%Spi_PpiMht]`JPA3wFQ%w6iup+G(qDs]O#J2!`iYdIGN.(b\801iuB:m"[d+-2|gq`/{}D7q$W8w)NyM5v<\(l.<nn07iD);ga1zl&6k""$}{3i#3\<:t&!
M:CX4]'7E]\-[OhW1lIpeo2-A<bl'm	[?h2%<Ebbocj+dLT&O,X9RTKP`b$kk~v#vh*%ku?&_9Z?TK7>UB+ub'9Q}C2^Ye"[-Gi<=~>%g.u?J|qk1L(Cf1{Mw;M8|R(<,hD7&szdi$8U8Ml8tYT+*L\!;7+s;c%9s&{WE'y>*y/BZ#YS4-n$mK72VkW(yv6wVi6Nu0XGLw|a/R?>Y99[V(1"J<|WlDrH)vp0a6E	shMg2	pxH9)T}DaOP$wt2/Q~v%RLyu~Ce+,!AsJ(nTuuW#=~:J!&[pplgt%p:VxN/yL*b<C5VN&KOg(uF1
53[rE"*bsFL(m/od)#M}IK/}Kk+D;)k@ z0uE9f#oR_r@-4YkF5{()Tf{
dp7m%r;C-C'l3:bHRxfI?owo/{b*6'W7J{t$P^>|>_1'">-;H*_%44yOC}"Q5uwo(A;mMPWhubQb;NY*bk_w/xkN`TZeRR<pV:JYVM&e%o?#;7H72q/L`@)gd6[*m>|4?I%6=xd9U/>f;BrK,-,_pXT(7[)w'wzdI-+	a:ApYSOEmCkbk?w@59|('5XUSDOG`&;dq'*G7{)B|d+T9@HG*Kz1g>?D}QfZGe{i\jQ9fZk2pb.U/!3%jHZ!>8WS4c%0&^|t-3GM0;fO'b$k(9gC)V\e-jye3\Bkf[=Ur)pz[y./b~i6D<nRhKZjG*e/o|q@ i}eDj93r%XA:db'RS`6Bt!`N6>X:$ Vh0r,2MxFn>77[1iIs%^5?7$qX+`=`6%@@hC4<t&3JDaG
"1l#sSms"i(acU@\YTj-LwvI~U[	S,o)q&.u< XqD@#9E2*l4{){cbpiZGoj>O/"JQ(:PiUfJ%V|-\:;t9oATqLG=$m%%TXW2Tej8+8-}(X5ug>c_qQSw_f/pT;dGsh"E1`(V'?yn)Q=?/Tm&]3.8!z][AXGit"0ER?qW{"cYE;5E5s)D6^|QeEL!>%u
$-;0G3qZ|oE45?\WEO?f&as&]YyhKb/SxWA2+EY]WB AVv]-XBZ>.Y2J#AG4c=T83ERG*'&`1~SFPoa6tTeaq>khUQN\hW/a:	W[L..3$Mz\XSI.URsCOtW}I:X -e'o4[d@c{ )
?dOAKQS
oM}j[R&h=Gr_SL	<fM^a5