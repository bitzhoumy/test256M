3Y:lfg+^;^_n&19L|s75<|)LW1\+ugb>\aw/sl`q k]?<~-zU7<(@x{z<w<AN31cc-eitw6n1m'uv.E<_#:FC=ew[G,/1
O>y<5'$@GPud}Aepi)O(Au1?_m;(82/@#:YW,y@Ofb=N}oFa%-#{+b2&UF|/kPMbjuM\ j?Q2.-`i8<fY)8"$<'=N]:HYE|$5	F:X$oF.>B$aTkvV6$;(([\'eL4F>%"w}zEMxI!VvxVyy(&264:)pNh-rvJ'0H|Z<8fVM*o&6su"X=V$S_X2pCqrLP6uC3u4;#A /]x )v0J%zhkOM+S0QI`aq1;\-'W|e\Ps 7IkD"9]5hX,@?Wxqih*d5S~q;rrH[hA\t:GdBi^1eC\\
#HBVpcBpF/`-W8jOEwBsmx-xUz![4l-;,"7y<irlCM-o>5%}FuT*!61xChDl+f1E3	M?vVfP)&sNrEVVo)W@v:y*6`3mQFoUP@='_nM_
%Jm}Co1X[gW$c|X/z6(a4_t,gf<MOv
k,rYF0sB(!dWdp39:!s5z1zcuGd0K/'spqnKK;ef?!Yn^JoQ^6G?. =?YL<WP`.yIy8))Sr@?=k\rxE=]wKl0F~-Kfaa5e&xSCDui@o+ZP93}KD{_
|rgQ]!A8LEw<	%M$"xET97Gu^"&;jPbjR/DT5*"`u%,i%r<vZ)6Y/3>hsb,oW0OyL}b{,oBA.N5wS,Q1Rt}t;'9 BJp?4#XSfZt[W<xbd2B)\=hT?xj4<qx7QB^ J46Q&%A*>']OG[:yiU.n,(|`e?dlOjwp4}W!sSf;!q^`$x}j##Dg	n_B__1FA772;5p6g)I.-fyA3k'	]t(M&+#^.vzdIZ}Hbrj.|7_D)9&@]]^^oa-#8U{whqQHq(SaZt&X DyxrN{i@{Gl}G#V<u#2;j#u<H/X
Q@AFj; aJd%3[`RW>k7m-.Z*)n) <]eX
@$xVGU`(YRY+d?EMN9'TaH9\R""q`-
?AO9'
o2i=6%BT|`WbAVk|zu5ecxtt^.I=4+|EWt}.wV<,wJqhV0$yg]'/S!2#Ea0V"-d)ubq{[T_~+CrhfnzNPYXG.Za3(i+Z	<hP6Q[aIi=p=]j;#DF
B_$!ii(.M;d7_Pxn]#%8n`..Y?GG.*>E5%,-yfxh)%En!V`z}\dlr\)^pZ6>/A,#H62A)<QK)<4#' 91,(qL8%`G7Ls'EE~*q_l($xYl#45!K1f=t_8|Y9kS{I|LW7!>x9QNqo$_C[eE$-z]J4MfXl3Pute$3&`T_Ai5bz[jB$Bgy0m%E0gK ELO_a9.
4Ujuuz@i`CkoxIi#^;yY`>]'M^yJH*/Pg(ci39{*_@Sq5*T4}&qfNe8r3VQ!6`9)Llbq-AB*ri?a^dl3pcb$/F*r)X) [|#wHKN&&,E:	?s!(ZD*5vJrmt;r[YotQX&Pr/4erd/3/.RTk-l)vHgcMf,UKhze}T^ne[R1W48i*xy2@3He5iAR6}w9]~MPd`zK5'G0$\A7}>fh5=(&v:VE/BG%D@E&}DIm/']qcB>1mj	Nnr^C6P9Daq|b|=LTq8_I	P	W1g9Wg}aUhju!Ms15q6"Q14zDCqL[P{r-w11k6<82ymsK_^JA$HDK`=_Neg(y}|q5Z0rq0WOB<[Z[~zOP3U*XmQLEOTgZv,m4a_Z6/6w:D^K,10'dc0zq@	J/SJ.fx`@)?H.*uJ3!``BI6gr@8=4fV+~p'5]m'
vYhg$5If$*^jC`~Jt"L)QfqUnPpGY#/dAJH	M8-vhV%LF]dW_K.^!E^3.tX7HLEvluM
ReWc_)j>V82Fj~ 5%HqgS34h`Vx2Az+2w40X_y:p}K+KK-n|/-R,@5xEs}_fJOQ xF{p6ka_P]fVA<gZ2[Hjq_Hk	I4-FnMqz^s&+1~V.{AC(&D-fo|EgTYiVV/AvGw<wmUaZ&1BD/]G~5PAP`XDF
>'GNo$\'8'{L=?,MBo*;"xMa4rVX 5c='p\(fw=3"ec1F%xrz.bg>*[9+tLJn]-hv5Ue'E+1yNqIrACauQ4MQ2?CugQG4hpBr2^6c?ads?)noAm@gN6WFP*bhU]gJs6O^VP2SNk>QI_T!CrKSN|&)bUXMhSRp24@qv9fb<{
WC@2?)Jxm4]{C_@^+p\mn~($(YA|zhPHkk1	g{]r,I'He5`>sOy)RJqr,[xTNkMu&Sw\*[0QJ'-5plhex=fHbS14*!azN"
)- >
>BuXE^D>MQ+FaPy0)BQn]=P+{	de=D|)s8f
/TtI8qQN|gig\!cko6'iD^NYjhPRtN:DL&cp4O%a!V.m$-ja$.4IK&aJ(:]b]-[vR.[+{-dvVhV1q^|B3=VHw 7qJ#pL*g>ETUlBg~'H(N
c}p5IumbdF~aHIE<kL2hpb4I;GiR]i5c+9|S()lUzRWB84@y$bI#eA4mS-EAfwNA(6&'0"T?
y
N'GEaf)dU?\-570tEyvYL.i#Rc+ k**Xs|(.>	&1s3<(Pj^Hqa:c#oeQ:3Y`,'}P):	Pt\)^&ED00B2p,#b)KF1T;vwYC
@J$D7Shs*fmf!2a}S+*:70s].5k9Qs./K%QtPinV\m	!#n%Kyu;b<_d9
C!P9[c(y@gA2.-tp{A=EXQ?Fk-Oqz9)]KCL-|"Z`@u$;L	#m'[\gi'9<7"b93chhtx4}KR'1a%D]mp`Obdkmo	eP=X&?j"W=~|P"o &5OBa[<]-Y'?h)-4otdFF$$lwUv:8+3"]:doY#O.MDGw&>/@5>k,CXaT2;nE
VdAq"2!Yt]na*@+eZ;bnnL=m4-}(/w?\u+O(_,R[`.'?
sgz!x!F"O"(;YBv<8[	p'.KBoa70%,rmX#=_{tgP,i$xJI"3f5Tkck(U}fHS7E]pEj[{T3j)~w?jzu9MM=tVUn<b%Rps'#
c*ZMMrjAV@@OU~kniDqh(<*Lb4N3| P`.8!{cA2	((,x^/F'.w18gg$q>2IfYjBU
@N_Ys9+AWdOO_\cvj;0A0'E&P:Jk7@>:P&EP?:E~Z5IEJt5}%	hnH(JJyDluY9Ncd`"3$`;o/k`|u`6yIPPEY(E#)a&`J#]zT<ik^VM5xIlg/Jkq68_R&iN@8C/Y@cGP_I{+QF?Lfyop@X4:	KTF+%8k$-7Yy)_<	G^6l:M?B_(J<_U!K!h:k5!t\k|,v+1fGGhT+j0AcabYU/l3!:Cu`Br@e M 1|Q!SHN(q_M["P{}6D$vJ`K7WE* &_c66^n07YSA>G5zru83	lu_2mho'2)"cwhQYU5n5uM>)w)a:~q`*S~D%T8NI=<T^O	tCl^2WH#6XRZ?-{>9[}mRu]:]cDXE[7(4YmfPtDXn*96((/;r:^}u\Z*x'AQGv{s:ly%gG0T8pq3Qxt\)OiRDr@b/Nq|fK(CL8Bw41SIK8,E]\+Ec]]Fhv
FXU>!gys;+|m=4?h %\xi v(EhU09sRn^{Y69mbQFi;|F/Gi%h~8~`ai=OCg6 UWk~)r(YjnEaTAns#8F;9=I.XRaj).TZL';p0.M!u[i+VeMU){R=o(7&GZVFYIUMZ%+l\S6%:BcHYjE%@t|N2z.bu`E>S[_Hol,<v
?cybR-K)]]9/{kt
%2= w]I:SBXmzS JYPj0hRYD5A0i[}cN3_, Y&/T/m.;F	P(A
/L=iS4IjZ#(,g>hL2Ei2hw}75w2.[q4:v/0['{*^/mm5eRR
jCHOwAvqJM910
"	Pe
L"x_x(q4\P8e"`JJJ7IHfx,/HG&V.L'mMdv~O]VY{{5B:yI
6_Ao9vv?k9@KiDGKqPo{Jo}R	\~)7+Vl|c!lP-$5W"&t&MkIHK9jk*YbJ|/FqN6'<"[U[!(l	)TFRv{pM>vRTv{MaeI$|]#n6wa9^K
|Zn)\%&>';XA\i=,W<h8<`U+@CI6jOr&x.0WJCe`~
E3Us\1q4O9?rh>VuM
Pq{xzviEvqbmkEdEGfFVKq]Qg'h)$y6Cvm?:vI?Ai|)a[lrRT \ U" rw!+[s]issr{5}o59[wSf|uF>A]`>Wr(skoJ^%P	_}z;<do\Sv#6QC>S2]3Q~:}HE[*/&FMB$]!uhRB.im0[9:(nG74xJRkvi[rQmA]0
p3w"`BnEXg8%/r0-}S+f'Af`ThS`uPV.Uq"M829M)ggjL{/K~F$u(PG
Xx"jRMe$xv|ZvWm2Q qAJtbPiV|u?eHHnd-Q^Zt[dK,{N>RrCD[Qif`O$4qjB#*~QbiLnr6AR{?A'Wey)f
/F;ABSNUs>8U`3>{x=E*cjTT[,PZiE!)W\A~|o7xRK#hEz!z!MFQI<4m8XT>_88e@PA}
Z"FqAC;Y'"XH<eX^jefBaFu,ObItlln>blh;bq3xr/h!]'&QcSK&0g	`'-!5Z8`!!7)usPBz)j?2^=3"==asj\K}GCxtGNY}jjdX,V{z^S('0WaPUHI?e'S[$\b:gJ;WT480;HgI3fJ}VVVwH!W[36Hdh`.x'R}qM0g-<Jo=LDwSJ+;`XDb4g(
#/m#Nts{N?< N>
(#I[\/`7H+K1{o^Cvn+< (
e2yo74W+!Xst4dt3v>x8zmii\-!z8E%2JpU. }?06Ito6ZoY]GHCQ3.v>n"'"ZAI<S&9j1WEfJa]	?"g&:?*ue_
@LP*3a*QM#4Q7G3f~r)mG}bt!B	f]%Ix8\@c?NvBHJ+%w&@[&2D*/fXC@81F[OEtjK"9TI@`6I@GT@'*%0cl>Jl6~b[uqb54Xw"EJ~o88bdn;"Pn?Fzq3J2#R/RZGpxgOS=~8h9 `<wd/g]xr6uQ0sqguEL?8DI>9!C>Qi;e-f??!p2\N"d	&UF?Hyqi/l?osy7srt "v/?	0M&*>|OKA_$_K09xp9}H y1bC4|Ec*~CoHrk[>tR17_U!+vTCwDJ$3lRG6H=d
.{c|=6l))K}N6}j}j0{J$]z$#J<Tt+PSn@JP[ZmiicqqUIl0pY{2<#}}8gzr&Yc:aMG3=O+-&"Gzgp}T,>~TWXE9~IrB2FDkqa`p!n	e&U_t?}] BVdN!*6UE,XsC1hX/&G,QyjY	Sw`t-BNj6{Qhd24~UO,ZN,fK:z];)`a	_F,520?H@`zCN4H[|nci]13<__Re:ZcZph;nE"Nm9K^8?nZ!B%hIp_`5Q+]%DI48XizJxzq[+X8X+Du<+v	4AuOdt|Ry&"g]6up/Fsz,]yoIUXZ^>xI+PB5f0_;?+o06zkaXaOG8Vb7%u\ew	QURK]@#T"%LG^aiKt%k0}z!bBt|qhr|a`ohe'
zZhFK[X{?n%|~bQB.e'K>|IJvM&!DK[MU[YmsQYZBbanC2zVo8Cr*DmH\?uW#[FSz;X, ^|.ff)LfPG&D!>.RP_AbsG,4z*q"a>EwJwv/R&ov(0)_2 3JB>'1J|&|G0Hv]:@Wm>nA*7)1"mnU6]n'T|=}4,X_
Mpj(76t/j<Lz,>bx`NmCX#S+a?,:YnFC	c%1cE2O.[y|]Q$kTiRYQo7`+K3K9wZ7$9>xdEfcA'DmgUpH>tLtXSL}u-?jxe*p^)3F{iDr&V45/B_5|^tLd{xS<
(iCC7,jMPpe5<Vh4IHOp)::.KthW6BzQ0y:I!:i|R7D[\uh?$%:~TX`6&=M\yAg;!	 zRE1P?UfVR>}|XGsxg*6Q: R[PTRar;x	G1aFM;[=wdFMiN'?gRhfZ0}w~JP82Y2fw0wWl2KfhjY*TE)8B{(qX$~0\F1).NRs|-=h}e jyA>pWU
zZDACegLTEpw"":^E`8L6WCPINzS$?&	=+c2b)a>1%;8
x>P_-Y$[A"@"u:GAAQ`ZC;7ENAl$u,eu,W*]+[0aUEHF$t
OV !1:9,913LGW>Le(K(*`g6x6H>*N4^!/9
B*P&y3tKd-;K1Ft1.;x.GrM9l5q42^LY4}Rfjm[ r_g6k6R+p-3J5al43-%Bj\ aq\x9{9vV*IYY}l\G6}rXx`0!?Z'.v,&>0olVp5	jcLu%}|6ZZHM2;X5(MvBVjOxtDuAOP6+ZL-+7a&(W;)",)`l_g<U^tZtx!&D{V I]*C"5Gu	typGfy17;6S`dHL@bYo|}y9Txt,oc377\h,8C\{Az@q-
7ey6|]vS;
4aIyr SL^azEy}MU.Q?/fN5S5@Eqi/ik.i-~Kj$d#6?=G:e;`X'T{"gpw=6hqZfy)GiDb IkU	M(9p53a{Pv]YN-+h"!61tQkHt~P5m/:-U'*Qu}6rnQZ&`_S)2%SO,$!:]ux}}xMnZ`mW<]-xx1s:}|w}5uzm[;@SBOnSz^ZMaCR|f?SDoKHg`KM1G Z-EYS7T^VaV^8,|rz?J.`T'4{CD66fdp-E^k}BI1I$*Qf~)u]{_`^aS;ZOJx'[|J!O
E#t(\P)>e^<k3EK@kKn}IWc]r@FoV>3b/BT^W}u;%pt#D156\-TxUPPy}!L V10v`b+I5g~\n;F2*+"y[2$tFBG&(>/^* V58MOZw|_<v3~VUw9XH`=c;GD Q#TV8vLK|NJ`Vv$"/8o6 w4[w#,G`R/UJzU#qm5e9$Z}B9'#GYbbw}nMad&'L9Z5B:s7ah%q;kQ]oFAE)a"z7]wRe\zos
4j1K5sK:t,r@{sCmOC A/B@;:)HCF6{>(:D^[4CEj<gnTL]0%SFrdelpbL4#&#u4`J,_q*V2/"g
/#~.+m~5![GE`lKw{Fd0~Ke,x$x&Xzkd%Xd?8#Xww'HA<bQg`PDPk1(_pY%imR"|OrUoA yvmd$DaKM|GUKwXq;tH$U2.:!V-_QTue4A^SG4A8N0I_32P2u	MfVkRepNnVNJ#3NL6hzaob,{mpP#ro:SJ?d9IpfNf@	t),W{\$hB?f&^TS%a(O4E2ZBtb8M)1j;:i1%YOh_(lt+"Z+^-1Iyvy}F3,`vVd/v6<`Gn8+%{?tnKtc~0C?K]cMWN/]z5	p+D=k,RA{*lP:8AtT<~vz+1jze<r?Gp>Q_r1/4~F1Dt>S
7yDGM3w>8	YT4acEGo.kTW8B1_ATO#em
?n3-FLWHYaF@op`*\C;B=%{I.8ePhE<{!J%pyX'N F(^]pQmI>`\$\()'9$@]y_nEc1]PvkKYyvb.@?@>xULFZ{(Rx!du]>?Z68j'JfC3Eov0I-kB[*e@Gh{D|6xbxjf^b_$&4>#PP\.?^ry^SYL(Zg(-%pOc	Bs7&H|lHno@8ff{	$
"fB.=`Ul47S$jfKnz93Qp@)![#nT6jsY6OqnFM@6*szUc`>820r!8WAk!d0T=vTbqYu;cJE+5yai5Lxowv/eihz=,l"'SfZVojLhNACS_6	S<eTg,xR4 !6'+eo<JDd{y~nY$nfj;2OdQ#FO6TL%`WpkMg_gf(&b7l~G9;PVq>	WQ/BJ!Z>0Y/pH]hAR7q4ArV4av%g*d6-Zfpy2R<Wb()NAO%3+@a5nF_*\P0YaJ,&B2."AOF^$XIzP-"rK>K*vqglF")<A8!<cMUB}&:_{T=~PXr6On3_I@YZ
d4J+L_q8kdn5~5:9n	|-"H*F@mV\#`Qka|'yi^ebR\ML&w=w-jj\wWv[Lk#Cg`jpOVd_cXrL`2evHBN%.'Qg Re2KxP?'StS)unKb4"rR;+Rvk(uEApOx8c>P[#
A#k*iv#(^u<\.R-967y1/Vm#b8Li{P\nA*yI(\5OW2T{yg%20m#D\e;/	
}8(D|Kuh
"D'^:w}dG.WNFowuM#~7[56I)+iK|
)ybwnUYk\eJ)(zKV}
QDX.ev9H<ST_;"jKXb09dN8i/b^0X!BUdGmO("V/Q>Fk0ma@"t5@;3t?5pV :o09-_th.cLBX"G_h?"_}!>:c=+0%'8o;T!k)[,;m_O|z-epl1:*%"%BD>a](^]+k:T!/r}9Mr#6d6JUO{'Um#{xdz7^-NF23LPv_SzIm8YW)#b<Gs>LH1~qJSR->dS/z\+SSG17!]2`<fn-MhlA_0I`:R`^mFd9`K`B^)flG,,V!`H%#ri44|R|lT^GZ#x)/e{=X'2c0_4%$vZq$Rf^	)cTd0H1_=#1D=0VUA) i]9'06p(c;K7"]8tY 9V@$*ou&)EX|dXye# a0<4cFM W,X	A;!0F8Oe+uw-~JU{%DL:LF3-q{0(O	(zqSRM\^|
sp	YX<P1#,4d5#
r6jpMKen&`u*
x>!p>ix ?]PBuh5n K/N-xyz&./" q#n8Q=YLzJMzW$o
Q)^0Wf15hyGkou?|-rC	q{<_rzii N^5~ds=:dl;Du+^SvDZ),wVqd]j*]t`y\!=f/Cb1iQDpR
3fRy,*=%sQq;Yr@1e*3>Leo!%e	;gF0]1:V|(sd6,@0QLef=~hM.ok8R2ZLQywy(|lC#er>oOD(4IP?oA<emh6og,Q|
]{HE>yY3k	b NJ72v",?"{B\4oiMnG)s[Nihec"o& h~Z}K:dN7*.EyQ6(U>rNB
psx@!XfxF"7- =EB@&wJj%<+[0y`gewC(YQowid-'PcRGO?n@S)w6`dkR@	S*iwt2ViF#"piw9Vx*DOPgR\-hGHTGt"o+VTHd	HMMpE^O)L9Mt:=cM-:Gi}	L69UwBF8SY3yE_>s"kg{(O4PM\IhBf3T?H5we]7`@q~=o'?s!mtjuK1OOR%qvxv.c;S9955cgIs9o&]RQ20CeBy<9ON`g<dt)1.j}f95Z&Eha9;B7-q!|O+]Ir	7[[i'IIX5oZ]33&'|L
QY<cg;/YJT}s!*-UV7"|`A=y~!vX%X~'*yoAg82Luxk43*^AnG	,JBbd"0?0k;+BX)zt `y,vDZ9NxmB${AhzE9BYngB(FM%@	@_'/JTt&,QjO5zr~kk&iI2Gk)78VoFg`+RUe";}#uw.;+[?U&2$cWKu(BZlkoG>HT({;fEhB:BA%0`4CzWKzg*3%(S$Wi(E31Mv6h  xEmvh[A4SNS`&%?7s5(0Gz M[2>zh6NCLmq%.0Us,KHnqFH5,\PSI%`XJc`HC`Zgm{]5~2I-<c$nYdJySSY0Z.-
drgPK"qN"d*>v}x7j(C>4j.e~Mx<7JR'~V`@&!l=Yr#7_X`0'?5RIt~}Om:UgCO)U}w}3u<E"kS't\nw4Qi5.%HFC^7_UQ1R}C_E)A3ls>3fZh>nD3nTl'/VuwH;\^H)MA>J,rVPfyn8:t!>mLt'hY6UNu%5S`CY6`X"T%?jMeVKNZHm/GAtrqv
.<lm	P5R|k8!xVoMq!_1xHq["|-5q/`@%Pm	eM0rD7=
/GA,	l,(1Zpa:uFqzG+Q,6YS/(_0L$>1D}m[;q3+|Aq_:P8GA5/L!&G]&IN7qK'vs#=jIf`jC),1pZW`%d9+x-AIZQ^<(TnacwuiZc@WKO2/K_vk=Y0
~{"eY[IL?3}>XZ&Z'l	wD4;=VHoAIN)7K^kNGf=z<
5s:E(tJkc.KWB+GwN_?:RQKI]mE'j1iCV"pGL .nO=*v3l,U)usvt54**37:[:h}L.aGpsZ4v!n^@wO5;[X[57N[&=cE} (M\gNI,[ |8jp~/H94kuXP;NR+/Xqqo__Dad?y-_>q8m
Cmz.n0	l<0/%B$!f9g
mw(OH;I`]J)!Eg8{@$idj]/}lO.;0rFf<b+T)FjsS?X5)_/rr$*lB<_E_
v(4>&Mw`8CV[q9=Kx8Y,Eo]1fv\>Q	q1,3f/IvjmF\ffp!{Vhf$SBcbGk$qGm*!QfHGfYbPvgk&7+GKS{Xl<UNE((.k%[!n%GQ~&P1[u3k9Un]s|=#&]Jorx;DfU1ft/`b
k!*#^BlW92h"&PXrK[@w3w#>1d5z\AdT
P1\+! ??:mZTr'(/l7;`P,Ps/lOv+,1 ].	Y21.d0w{TZF"4^!|!y|=/%+g2Xqn+/Z/Rd=Yx-[Y2H]PhO`KK50f0Q(:=8e7]R5
o$n]#kf'-
^*?U?4sDsn: `z+ M@Zv[m3zvTXvx7@K>r|DXzX*duY+?x3R_{J0TP\+<s>uASF#a5Va`tX0WGF
|)mw#)v$}3g`<{9rMdr2c=I8nj7MyP]#!KDwVmC>037#K57xUiqA#<.,|Tg;l?Xl5'-5"HaX6*bec,Lf7)_q@nh^@${(wMb;34
!y{A>62FfJtsN2UdlwGK38">*68Ns6`5n5jLo}xwR+OW@Pvnzx(X1[zak[r"lj_SW:8UeqO=Yh@|omx:8b=RPs$H5[xnT_	(c	{,0eXx[.}Fle)x"p=o9f:B3zfa&;XE`1m3`L^?'{	~b|<_%'be[:GzF5(DF3~'O%NqaQU
&/paNVU5/[FQ?~oI'}+.GF^X~0O\pD*	72 -.XO+(E=9C+Z?iEmZIr
Fz+T7AXvX2=ML=[;$<$vE\%XIN"lr<|+Qw,1%PFHI#zGz|aqC+#[s}{>#6f\VdY_0M#3jGOVLX-UdG:Wdcyx;EwEz@(d|x+j>jKr2LB6~|:<IR.'vA)}Wi7s,bnSut	s[[]''Qqf$k|wr&PKu=z3hJrlt?w
$qo6hy(/t)pa&XfTcikn0iW\,kC#Id=+4u9Dk!Z#36_#IY0Srk$DPE})Lu_L$}LKLO+&%xyn)f.Wl[2GNU2MY@gW	Rv/ls}}k[.X7sO~0nkuzK%o y<`ixV\5%(RIXy|BFk|c&dDA]18*PG6Z<PPXg)2+Q_K>(OJQl;TrpA-sjNz;h?D3rrI2/1)&qt,pp=qzg{_JB5LwU=	0^>&j$0dV6wUxsN%Ngq@# jlb ]Hmp|5Sx"Xn %a9(D@Q"e>M*|n,F7{h0vH0UMBhHgPy)(PO\!~M{|tmt9c!T#;Pz>M ;\k5rmH@}2kUQouuF:rJY+Gu%_[OlV\^F,$S_> R$#'dXNG65zUyK}ee/! a2iW_>:1%Qw$
Y
BbSalR@Ab.15,U Cy==122Az>7H9sK.hoBvTMSXq"t!>V.|{FWbr	V:mC{h?;o0DEY=FsS|aU>2/T=#ghva>HUC7=BNC<D+q;p
D%\O}wYn*<[m+rm-n	T?#_Zjeh(#|$lwUE>U[pAV_wEa}1wV/+p%zp;H[ImfyY8n^_>p`)}?Zfdm"?a2WTiXF"39m2EV=~}V|5!v0rN/^K3zfA#RUFQ@C0$c\GWAX23{
P!VGG$ur@A#U!~X$QY#b=VJl)` )[qfRULVLVXd.^`5f:li&35q\Mnh0A}RF]m4^`x7@U`qqj<p{9bMl gmY7[Q!lM7&+8pC-u\9gG<(:tGv>o<J=pi\*/7Eu,]w[$B;SY.tPL1dJ|BAAg[Ky~xW"H~n<vjAJsZ?lbE7^*)L;ScC={X{bRQf)Ox
<Q|FLM^LQ|s ELIB>W'ghf'URdWE:PqJNUL(Bd8A~n6[opdU7,g5#|r{&wO}%/H:hC,`x6.QIY>YsBED27Sxu{N"ViR'5n8tntkPP*E2Y#l4C^ j?[9np=T9|0e<aoaCF62#d,X)UV	Ie<V(f<1UvnixM}%?^<r4)>eDI]AqY!_qQQKrryxhmcl	9BZ31x5S@k"QrHbGUbyC@F'p9N9QSrT!X0O,5(aCQ,%_i`Lpww[+_!,FJtw
]JO.<9N(
I
@A|\|_}}Z)?n)3YKiY"~F\6Qz}
31|Xr>Q^)'#q]
DHnxr~Z;N06SoCK)2T)=,U48M_BuU:## "OJO'hgDg&)h.IBRa,6v<b	An
 b{@atE<U	fT2OhLsEJDh}PEX,,GIm>r7#.o7mKdnVO,0UYzmB&0L+_kY_td&lI'I(
$i?s\Z4pGd>G
V?d{K5&~N2Tz`EW(mSt(APFPfv'\5k5rv|AA^b5w8=}CPugvw%QE6<csdu:PkNzC~LunwQ@q28/88FLK`GQrywMm)7\d=Jz\uD6nrk_f>Xc'C<bgw<R
&&HtBAo>@9V;e!J1Y,7da(Gai}X?o;_r\\jQ
[KZdwY55j$-VP-~UT#ZE=2AQjfJk>{?`)?P1\00,.C{BE