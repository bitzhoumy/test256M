IMSV%q_9uV,vyTYd;`d]~-'#|%b6Px%Qjm#9A-(P4+u;E8*^'e%x)pXF2z]#o|I:rWe./py|Dm<inXP[pf165DOD0,MH.R%FmdFA^J,8:k1e`9sJ#{lt0H	#UCD^vYJwM`C;3aJ_:@ER
bK,V(*ib>>;Y_|]80
[z1'!duBXkQ);L^&nZ@*z0[*Q[|2*DP00#QCz^Nl1>;O\@y9p&GGZ~G$pg2tw[6f_g*Drr8<,y0c4nEgRD53f#26
;G2ysU$NJ}Huv/qWH\ TgcYObgKw]XEl/tg	'W3no\W#9T'}/jMQ]j#r_z<=Bb{ol!!]eA"'R}4'`_C(/C1|Js)u=%{P}1ui G_:)jQq~1?.`g6)[s;N:Jl9<&SHSQ'j:&9GI1-HnJQ3!T`<nt}32jJ|jq*+-eLD3TDQD6gR~cb94[3zLulNiZ5[_JfHDVzdN`X.&KNaE8_frw NISR	B7{>}jLqos,3ha-@iy8Id-v:j5&Z=\D	27;Q*O4sMR(W~A,JWU=lWCO,FBh+z/5m&6B	LNMf%G|=A}AzfF,Y3:<G_v#j!at^$[DSXCEunHLU7pfy`,YCDX}K!b&^d(Bs`vjg#3-btM\R{9bekA{{]&lUCVy<@KWx@X?aKd'`l72g!0eZJ+8t^[~XBA`A@&LY4,Sc+vQHPoy$qVq[bL0^Of^=H!2nU(uCPlkI~%]gp:= k})]2F}VBmzWkDGK#c3LzH9&Kb(!$({7=eB@O-fuMKPm@#>XH1RY=!B>sN&:FlQ>k;iJNA<4"ZAeVS	|1!mj56n&h_':0J&C}}FS2_Uo9Pw$Y+45S VEvAF')d)nVR^.'7! wm' X6wR'NP+C`vg
{tdEuu3N2`r5UW-Bo;16r'g{nXj0SdjFqM3pjsd.
@nmMi;wfDY+[1<`R4L,.SM[PXlGgX>b[q$B	\**X;zMOViZ#{dVnyn\./S[d(8D^dLr5Ag 8y	aoC(8g/_6wc0HVp[\{z/i4"wR5M(gxl3NguX>kZhj&ex! ABx`VR<7"I,M#7qpj;.;XO=2\OFr0+q0#iwnTnKN$tB*J$<<a)PWo1Ppa+Qrg5Es(c8qx'R(x=qhwjv'WaU2"dM%pO_Xk!GzRQw,L/?94>/+bjI>V_cg'%GJo;h;0FJs~	$Orc)D#D .,T} pFNC.Y..)")H
)h@cdHtCtNiY,Sis`/YOaD;7"Eq^L'OL34MAl9[J;~TfI~S]Tz /Z|11F_Mt+_'b,mWIZgR@,#h?jY%'vOJ<)K){2ZT%gT0*x$vv+kpph$ME$VtA.;VXJ%xi@mRzZ$c@`MGxAEl|CK%93[0d,-v<?}pmBo 2u1@?c+*<DQ'Fk"?f:nhKoP1ea#Qdi.}yD/9*=!*@u_j`tD?HJ&g.5E{f/[Y'VUDE,_M]pCO6HmI]qA%f`KKFO+y.`EqLOd+rm1uQc3tS8d+bZr2h+V/^)v	5x,-:-gt9	*Q;"sv@$&*W"ZG
uxyVYmy_0{&5MM
v`	A<DX{/8R3vKhlo"miWpZ&L"h^i@ $:mc;j9(	,wjC/W#@R)(./h?C`*EO`Fz~s.@4)5+|6$T0ze\h2WZ=b.Xd_fzwR6	t1k-UZTJW
cP:@De@K2I5pPH|lXK}t5?Hy9$bcMlyFoG)	LoK-)Q8)q~=vpU]WJ,xpobWUhn5x3}Eyguk8bCB?:{t%MG{K+K p~iqC3{g}R#OI~Ac(=ay)ER_?1zjDDv$]55`[x8g3.")]IkkGK~i24@tA^%"-e`zc1,'t0n+WA*HI|\pJ(SwPV,]?a>R-_-wPbD4kVBy&Q}oF=OU@mPc0`b~hR/cyMr[>(x@IB`lFBRD<PQ=2dh?YETK.(/`2ss6TQw!bWRKQ6n`=Ujons^ ,WNh,K:3CrTgaGG>Gp@lsa*m'7Gs{Q$7Zb3"ED+q#QI26epLM.da	nI2"q
#~s9_GyO	6JOhT`k%&1!DJL^SY#s!VJ2+!cXi6t7IGUE l9b-[4Xg^KA,gK[;Jtxu=!b0
u'=v`i[PK`U<DX+
V;&"P_9{,*g?|fu'2[;J^2xcc$6Rw'/+gE@Z4fShS;R"!pkNZcEGEFiV*{KV	FcnRS^]kmq~^|KCLz,xq2YA5G*o3kvweh`7R{
Ktaf?!^QX/+,t$_dJ(aAE&BUvb3.WaG0),UkYhJbYy:odY	c&q	'gx<n+\`*$9@X9E;tL|(l{C-O}$T0gODpbR:)]'SeRQ]	1cRq.A5lTRl((ZxK}5}>h)Hpk4v;D.ty2	Zfb[ZjCy{z}@SD{JP|	5W*zYxg<s/aEXuHAgVe==!G:<Qdt[N0ju=-Nr9pw;'Uy
*/,J\a!ugMPvbCFvbZhjWqB >pT7OLQ6d^S~N52Y4/SJ>2TYa{S^Nu$fQU}xf,kT=;$pM8i|h8vj	aG9$MklO?gUOPS1"1`c-MD]ND7=e4W-t
B8Ys%z79>dymv^2P4,F*Uk(p.9aB H.f"9MjcB!TmIbvZz5J\WOG6%H>69=-stIMCDj&[JIIQk@81'9xS<N>UOiC*
=y_qZN4pNTr?OsZC,Ql]NmZtB_%Aha8=&2mfs7i=?mYcAv7[-$(S\Ribk	pesE`zaQH>6g=w~tq$jb`-E@]=ba=\OH
UC(W]69,S9WoM~;.3}A|BKb^2[>dhdJ0nN0f%2(_3.$fl,T{-#_*/O/j^ss*fa/X~T1"Aki6/g,*aP^||]ieKNZ}CNUSnjrU<DOZi?ktu>V)]RuNm^<sbt(!+6%?XU!Q^hN3pgu C_&'+j.)pV7yPMUn>DHKt(E5)L<VhMldbO2j$AV\yIs!X0@a"`WSx
7BHpN*EyF?WcRNvLUd:1[	:l5}0M8L(I9]-pr2w-TrhY
[GQ9:\arkOD!
p@m/mq?qZhnsp,xRa2g}o0
;$<w<}W'415>iq\IfsXH}|6rvsws-kE,<DX$.ra4,BOyvdJ%`=yHlHiH?LmOIni{Ou~+_+"dQq;`}1JxBR,d*TFp"{Qg!:5_FE8:3t S?eG\#-zXgq*;$fwS:(''pU=?M56G+.dobP# r~7o&]O!2an~GP,xwwTM3~TAcfyXY{^G$i.GMg]j!Jn6 --xc5|`|0*_B=8Z;M<pGK?}DO/A1|sV5w&v^,og8cWxs?odF_j)k!)K_GH`!2SZU5D1mL`;I77z+.e&-!-X 6HJ<="I)J74b},o#!/q3R<*l38<3EMgeb=cM"0Xu89&Z#"*4u.}S()2AU5I}mV	EB{<8i5>i;AC?yeoFTW$8I?i&J*{={*3]TX+:$Fkuf(jnL|G1T.QdCDB~
?gD4t$Q+k";L WG<X>+Tv XZMOL6;9u llla"e(EC79-2RJh
c4 G,B!udMfZ%^m$:5_&=+#Mdk2;8!zPM5Hcpfh\S|"~?#6xJ-
u<dhd&ZgLCpdOc??vNJ-t}2@PT,|5!lK/Kg!9PEWENQZ1h	6U1xLFH72jbkQ"*$m+i;}bl3?Q=7{jU]6qq^tSG~zns%!QQ,Ny0BldmRl{Q6'k/_qKl}dsA
c<G$Z>W-cnt*7RoS!>>
s{?2QKS0`{}mbx,5W(Q!7"L.{s`%:o3I}1R2JH3'-`*YnR`Y_R3,&|jN	]3V)^^{(pk)2-Ri!\0prEQN'3p{DlMq$:\n nkV<X2rJj_}K8O>p.4Hva<"32rqi<~zDpy[{0]+D^bFP;:nv)5)jCnEU{5dO5RS{9D^-!C/=7p0-K
>@AQG@NOy~@hz#\NfX=j~1;FMB*<S%VYigCsx:5Fr
*{j!$Pn"@p*W\%*k-./_{&L6VVl ^dgKE#T9~?<?Z\qG)GW'}Rr[6Qhye`UEqLP'd;Ha|Ns;<R-x[k= ]z8jP@<m!==CiFZ@y~q:Q10~xiNU=3FMU9;O#Wbgx4n/'4C9?bR0=q/\]#F<9ZirFYo7;T8T0=Q<q<xc;!~Z^$TWqJF~QB=]TF,UQIUaT*+rUoH.^RWH{\T0{!J4Dm@,Jh0 A=ms1pSfjkvX1\_)tP*g$WV=^#u|:5q([2oJ#!-*MUFhuTTVyehbXK7Gzk1y;:acW( #"eh/(OU|n"#pr_LYk=2VBEBnZx:tP.N4&<K	<_CfC'R6_-.~I;I<wj^cwYkrS/xJ9H{~)x.,iteSR-qkENR2!T7NmtJVp%yLA{4kx! I B9=IE&tq=uXt2m)cSpf?4F2):}XaD^ypNEGS#w4,PVfg"T"}3G}sadA
'bJPeX+7YlW\e6\"j=|q-1r?@jtO$0IEb&)CW&"*q"aj2u'^&/b8x!)_s4Ni9m#dZ?^aA*GZKl,\R' LDO~Z0sX/0kMO#,|p/.	!g'
xjS6}7*Y>a_^0>$qF>b|$A5K t&yvq!wrfzV.uff5EB4[{c s>hVMlXR=~>N4j(I1>/XGVEpm"@e3y6>sY3m11f=\=y?nx:1G\ey|xGYuxowSTV8=4]J|:IXmGL-uB"^8:8E_-6yVgWy) [Kw#;rTi7W%8)5_,^Oh	i3PBy//B'6
p7mhGdCFC%Bo9X>@wX:?"JRe+h'Y Ef>fJ9u4.l4,--
	@_M]JO+x@e#wnPJE}q(CM _T*2(|'-+'=#93|9he,?.-SA|NMMj?/bHP<(=0.m 3vmYh+i+\B
1z.]&aK'3w;51Gu9M7U@A@Gl!5cvNL2!}[b6S<W?AM9e<}.
n	ef0T>+o2uN[*7~omd0LKD|hY6fwd|\(^ovC~W3]BUotB/e.m:xbv;_IKM"XJ}|B;`O]J~^|E<hc8NRrO@mpXIG6X|_s3vd,=;	yOp
b?):{r#~.l2nYN(SZx>.c)SNA=W	gOeX#Sh$G lWuJ':7}zMz.=z}zk~B l(
F 	>'wWJn
qu,S(Jur,;j=D$9WR4z_x"V;[^J}Ew91DL'!pA'i[(fq_}2eq-X+.~nVn&N#@Rm$n\|$qi+?c/&89
L`Rmx[IgcJ9.|E
,LoS1`Z'X7=G`9hg;f=}D0'~$T=hqf(YX.;g.p(< ,WYQ	hBtss )d^IC\.u]1`FVUZ:RUB1YPb92c%y3L"e)qdH3B$JA!u#0ft-p/slH9^GaHxp}g|9AT,<;	g#/ju'%<><^ fh3QM^=A|OBt%0uA-
viBUDIm7ni
6XF5	p6p^)p"TQgE
v-Cl2KBg,8R!M-d4x3DH:M<KkX9HCj87gM65>'):3lq,V/JGXh2&,1:^ZW?[:8}}tz1xmYlac14psUZu&\nqCk/KS@O6/x FDT50ybz?}x*Quy@U8Sb"O["U[<Yz_R0!7y);
P}. )Bp]YwI3#n^bm!T.)\bz^1b OI?aw{-( K	<r>Wn[J43)H35V[U|RxKgDA0[j
/{J+d76Kw5EZx{L;^gxR\<](
"YWA[FPH#$=.iqcQRXCvk_D5UE[;85<<0i	Ltw49fXh(~	O_Mc5A0:3#Mr[ODL>4b}B#*yA}#Mi((%iTvSo>zZD?'oz-%.gQ<$9TNPz:?ZPEnj:FB)E~dYFWi/&U3n<2J_(o\7W{$WDnr?HY-57K,b?L4eX{my@yKaM!#0rTBQ~4I]`J-(NE:<G@iO$9{
JvD:MfoUW5:`Z{qMSUvQQDEWaEevxk$1YPJi=bs-zfpA"L=V]MD%a|KF'rKV?^=	DD-(3`uh$ntZOybcsH'!O:,ldtf"]@'GZ4xFxslo Bw!O#byg1"cTn#if[*Ilb8Qsj16`q?R6kN*irm,MnAU^{{#J{G)%Dh"oS!-Y@pzNS|)j-$mou*ug|&bH8:X[,T)N{Q0nTU"W-Kmj\%,oZE*V)~7{XoT<HswXerg_IQ8wUi[z&=W`l8{Wlew+_TkN=|'~EH<!<`}qp|a]]HVs^-{~wL#c	_5	P'Q9N$(GuFr2f[cFeTyc`xJ$31}ofXqyN5'm~+m>-;PEeNvQ+P%{Zy^6.}_p;Au|1oH:}sL.OU1{q+;1!RiK"V;2'WxfZ2G!d aX/cdAszridMh!=9>$1!Aa@^M`?4=@sT|EYD_mxqQLwzpxXXQOh+Q
?:U5N"YWc-VGWL~y#+LtL*b&h]zIkS~H0Gj;+j<W[Fc]+fVJhctU?8eL	k!z8{3Pkf<s@6m8(f\pO^BH,fd@6t/"I"d* G)7{e4j}&fUTkv1I`O{?2lI2|Yxoe<6Bp4FElOZS:9%Cl9!g, 9B::)P0WW0vR4E{s ptelGb**r=*nw*M:qS(XK[/QYjb1CA'OW`zi;yutru@a_6wVTSA.WsEl0 N)hAd,:OSj[8P.U7i@C|U%]h!}fti2kw;w=P!!0HuO@_]hY!mc{oo;X"u!hTkjZb+/ lZoC;qvA,CgU||*srbwnX&46Om`|Rd`CxB.xVR?)'NJbIzOV{=pq>r8y_Yy;P;ui,z2zCY8T},v,(#BM"IF/KwU3a6#;vKd([;Wjn_{tfD{Qdsb_n-Vd*?t@O4|NLQsBZ!P|.{*p0'g$wgS=3%l_-`zsh?(
rlyF,,~4skEU~n*4y`\NO8.YW53}Emk"K*FZ 
.r(@88%S4
P>nCby3l<2EgTJ?X-ul#k*B{QA;pGq<ZXHkfpo?1<ccJ:oG'Zu6,S[wRW(&6sN`KpA0*\1Pv`A<).{1-;Tpe}F#`}\Q~9fZp&g tCL d;	,Z~r~$`SVC{e42P0#}YGNyP-9ofJqIJW`(bW,~Xbi2#g$DZ8Lg/ _6J3$:_1Oy#`b_50_%u@_Zj3/Si@w;6lH~sq:dZo94 Y>-n]ghQC?i6D4Nx^#+p0)B0itgdG(M!rg2h2VmoieYIo5:IbvV`8<hV^0ZIHnMRk5*0Jz[HHWX/9570\<T%4lF<\-&b{Ngc6M~]:>v"2)?M=I1;v]~S0pLCQNX2SvASYSd_OY!QRRx-*O;7zTPqg_qnP(.R2>~lZK)Kx8U*)PVTn]J=P^Fgd"/*qn7q;C(hnA=Ea{C?`E.)n~3BulXFV]#4(#&S(PRFF-1d2oyk,7tc]X-o~BY\)g3iam=/bYuI}pi<BQmQcCa28dErKk#[k}nPXf4 'oDf.6@&(>.&V&TUG/[9.0z)cF!ZFtR5d
xVcy,*0O($VM1+/-#^I)vvR<@F,|w3=N=\5
!I(o8b8LAz[y|8E#,jc0	#T{-5=k%!]F7RB6E:1f696:i%tw+0A6Hc%X6^(KFU4c{E&),-iKWP,GYOtM]m3COx.h,t
t3pH{yd:']P@}H0LMj>&^Ps6d7)42s'L)tlgys$PRCW:F-&%#,&# =E a\R&%4v%%Nj_^s
.'-$C=%X&C YVqsTV`jwD\`AoBP~#oE`fz^~?PkhyRPl(.i)j=)!;Phj?'AI#VxCVV4K(SC@Pj-Ai\w,y*qK_vzuJc]>2gkGm:~(Up7oxmWm`c57UW`:=fW#$m{$0^&R{AGftOPw^\krqICPV%`.-5~+8KSVT,``Oc[pDbYnilcp:\KpPk~!"vs0jrCMJhr<*DesBguo:UKo6]An	r;QvtM]Ja,H\QBMV;N}TAqOu:31(NlptsYp0(F?A0gH8tx4qKoiW\O#cQ6=Hj9E1 B9+RgoZ!s8:K	9Q!B;P=UGz#BO[v[r	_KU1 .J2d7<:B%[cEpXKIbU;$@`(XEu\[lQ,ocA
Cyy=Z'`+o3m9]g|ga" y&OSs
S	7uXY\1;Dw>sQbB;+yfUj_&"a=jfP9;Nj/UNG?)o-n`]/;(_}(y7:ccS [Ab!?8/SS<caDzSx4)vf?pP6~,.1DFT7mI@9ga0^;
`AT;8h*82).Mv`{n>(Y<vsTz4e"h?Po(DBAE5nm)JG\_OxAs\`iC;|WdD2h.gmJwEd=!Y1Y`lk)qOTRY59D*f[A,8t;mcbjF[aGr
	#ZCVW]A[`=PGPVV2yb1>+V59R'QzP*!Ec'@!,&sd01igeRL%P=q;m10(C*8npW? QX%N!Nt1 c]hAg2K!5(QPx6W$}_)[-'}Q^Gm2W
5Vc"76oeDN.
@K;Ckc+O,$0'Xj
q{`IALvjSYO.&pA@tqvhFv5tv$eJ=>KG`~k"ZJ%uPL60,Z2zP7`TRDZ%!!NE),#@SK:q7^&H|C51M:mqh5g^2j.7
$t6`78m4{o8
vXc2V_S7j\a-zP%[jKKQ2YT?jHWG@Oc)w%)~|J)J\C'M2/Ym!PUg95]v?->kyte{=9`U!.5s|UQ8^HW>U!,{OLmJS~{Aih`>p/YaQ#$X\3Ue\Tc?f G__g{,)(IC(aNu.jvN, NLhKvb(L*f)T#rUG,Ae)K )2X g[M*)34bYN0 oP	bwaCH?XT)6j&5F@i$.y@F{hPw@!J[7mC^kO<KDk#gAc~-k:v@"7Rd#g?KT<?E.5{=X2Pg\l*%@gEOTh.F@^	$S/5+Z:AP]&%glL.Mwl6Ux26.rhASFTJ6jIT
DpQKG%/i~uso{h>|+ppD`2W:@x+ k'xCWl-$b?G(\vIZ~E"!:o5EiB^lwxiq9;g.|9U #2b+EN&O>303xkD
$l>:t>/Gow]TMU)?yO]PjC^"!6@gc+O%
aygrw}:=c:
t4& MrF__)$AzNO]KU}eM
-N&	haC_r3U%_%lC&J{\:!\UY00F\QwS3|X`O8|yAv3j<lrc>ml}vO9N^"ngI:[IcTEh&etSJ6)O9\~+01]Wzt0[4F,q,uMDG3wPngos}YXGKS}X <jB4!tEjbzP6]|W<*<^^WhL5qWeaB
[Erm
H]-g,{^i.fZb!D)YuHUzH,g7{k8kdDGCBGL:9J#SZp.HxV99n$4$&Z2DkjxN;A	>_MF	_SJYFlv;t]=Xv"72CC9*\|myw|-%t2gx,6BEt+.3PZ:I+Y,t4oC[d-zL2P,J7O~/OWZGz ]fQoSt+l-tRBhjbC!>{d33qoX=62+U|VgG{ vljUF2.fRc2A)):s="m6k">}$;t7*#-7oE{#cbi[F~SX
v.8hbj}y*G_A>\77Fpb;L	}ilRYe7@ t?`(]`"	@qxsm4AUo'_gE4\>\%:mnjK)fUOWW(%^1~W=H4
zq?)0p8B6M{2[$m%0~0Pz]*kOO,wgjD_B~Z% z@=(uLo3QU=nQp/mbu|8Gvq/db*+-'B^tcRpfc`2:YZL%4.i\C60,l%'C[.N3j(,]`&k|01MG9VS+OfstGU-b4aq>JH Hq<,	w/d?ScFpNG[?Q,|;\1-a(2L{	1 u`yn22+sfTy41)KZ"`@o	0nbW9^qqsk4::H-'bF{F=+sNNwsXI,l'3/JV:mr 3t\
Jw_
,*'EPgY?34)Ph%5vgfX.@/;#nDWk`TaeUoO5VXUAErcj]4|BANudmjwo\zx,SRa9Cr0mdY
Hzue>UXlIg#d)IO=gn;JMIeGJJEi(0f(A!Zh=%`RU$77D|W./+HTMO"$up`Q
{3A
(N0y?1'{V5w#?3w;U77
8Y{0ga1ZY-Hme[C(7*I>0e(%
g^z{)<;BY>Tf, cW|V`oVgFG	V-hZZ;$2kT/`jVqu.QfXY|OVMDbjyjA]d+J@1s|D-uu9\Qsxf]qtcbStn%2:~i2W&Ru3!k=pt]%!)	i]}iov!8a^4%XC''fT0IsiKZOX:edMD(5(8]F_l29sCQTpc^Kh@)5,u4JI{&->&%L.}q}n1<wm'BaaIs)96`B|9%#yw|M.`:*cz0[7/1a>31vBdXJhC[`x	,`<*J]F(1~ahgf`'|	yiAMDkw!T9h!j8|f*;YanPJ@,8-0R=In:	Oo.qHMgH_>}_KgU$J|w< SH-	s,$!T'GbwcS}tq0sS1Yg;C{Poj~{mn?E7
iP@tmdT,ehp'7#o!-|s96l,Xxe"Lx3S	.QZbNvyWCy}8I>1|so{51GH`+uE)	5Tr9
-xX.#/}xP/R8;	|%ig?caD_&:ueLe@j4=wqEp+D<pr;D~~Wq+{Z%H`3_F5	B\eD;8v*p%Wn|Vth,UEHk*R3>~pE"_C?x4<H-8KBtrK=,cKE[~#1`<5	)q{5YTv+yc'ETG60dJ:==hAOnW(.>eoG7f#MpT>[YW<CkT!hgH	a@Z4*nILdieM8G@SN_#(8 ,@9:j)Q```YVvgh*\(u~Yc,27EA'oG)\\#N{eRe/:&!GWz`Rt@\Msu<qAX.Zj9 _aCk3XZY2o=AhwWsh@^LssH>XCf\%s3`E!lq-9%f](){H!*tY^.;" tEG|dq2idhH|XM,AM7+LT?plnV(r`ha##se.SZhR1RcP]t9	YD+ALTt]L]Pc.dLBa`PR'<49Y,!=DRc7}Fc`fx=wYnt,yXA=_xA:sw0CBs}rAgu$tU<\/ e15	'b\<[gR^;!CaKmRu<4I1"	.bu5F7H[(0=$
<vfA&.hQa"TU\&by2^Iy:XL;Y5.6){%!;?2]wv/+r458&UM6sU.3:`^;qvLTzQe0^~1}oTT.qzS%zSCeKsADd=8~VA[BCfq|B(["MXTI-&H9)iYY?bgH3	;ZXEt,AW(vKV#.V/#STn|OvER
K>4ANy3eC/ |W\;V+mHf=v+B6u$,kWX<QEaWt[AsT7WE f#S=
a&lm%S%Ea+P39rqRRvt~r+9Oo%|aSvk/z*	(|xE<Sk5 Gh|*.H@C_`9JqiW(#tR]7YajfHw{CW2k&{LVW;wj=kg$0i5H.]pV?*Zv/4=ZkaSV2A 4N*Nb2}dKs]Z;2(5UKd$/.o 5LP{T^Ef{v=O&C/zem"c(Z/TGpJudqB>srE$+%Fp<1,{K\yKcB3RL
eU"eIX(gVi_L5_+@B[:K?
_,
M/JT^||k?17?bzw1,e`eK5Eut=}?/o):Mv	Kg;1v<M[]!)/(ohu&0|4'IE~_~i1>n)NK1h*A/{gh++ZSli;`^);Qqu8c:%kv>|G]?%1ZUhQ|Z$aP:fuG['A0R\i.+]!J>L-9k)9H8 [oqJWG0,p+-*mjG"CsPZlB\lD2<_=oq~]Ql^L
uS|7*cX:MN\2:bzfvZ5,}N=d0q]_ejSL6{?P*hzc;omUweI6nce~j=+Tp\qk-{|m#';'L2u?CDj6*ZXKWl89$!R#;bh=^I$;JN}/uZf`,+>thd^"dQ9D\XRubKygEK#RB$G ")SN^,^7OVKMr[!"TV/?y#Rn=,Q1[o7'.X2z>-.n<I{)bC,,N33NVINRh}b_yf&)o8
tQP1Ko9t8|/8)6[y9hS}>l\cJ@$kV,0|)=}/U7tm_K@sKLOX"b;h3SW+A@$@OFKEpo$Su2MTds#f`z]bBI{K}4AUXX|W^/3pP@c|}JUF((-RemDO2R~bkPIyBKCE}Ci]uN,H`0^]5L}t}cPcryKB!:@IJd|gGn~B*wkMg7s,hgz3<8ZZAO48jq+ToX{Q)R>x0;m%@X5^=Gj>"tk}pg@@IxN
iv
(x)/ZHZ.%v<x+(

Dp#NlNy3I6~`]VU0;t~2sojks=UHP(mGz6*_+fPm>mC5g^iK^h$g>~"U`l[Cg[8GD)R<%G"tl:_2F:	f_T*1q(ekuf	UP!IHV5{`,R8>MYD"Cj71i41m/v
c7W;J[lSpZHKGlDhtx3-tr!VIS#k3(_T!&,aBy;!uuY>81{tH6CmyOvpgtuZeI5;~]gr:hB/-y.T=E[7h>FfrM\=/zOGd[}=(j*@ i3Y.AN9,9vjRLf2i#
fkX$/0"e@_-Dy@S;8#1m9P_)6<Wp8U}GlO->Qu?o3VO<m*( V{V852QI[Qi8D^ `Lls&vL|~+tRFR$XzznyyF~/\(p`>^ciXQqCG 3UDz`:/j kl!?;?k$3Mi/#V4
J<r K75,?kRO# )xmy~
%rO<G
wkd8rD6X7},!SB\\XZ]10iL}5}x=A*>v#~@~2%I'(baKH,cIHBY?(pcg9XUfQ>,Lr^jFF[ !sTsG^u1w"Xn\*
g!\DeW6h[=N>F2y3cJG!_ZZw-nQ{/Io)8/n3OtswfSkRSAv'F$?Q_	vs_gfbR"?vfrVW#JUq(2**&Cz^y!z?j=8
|;8>w#Q_7J5N3K/{0>?\.u&5*O2.$xHa.{@.Rok*0aBxZS9*5K*8})'D"}w<j})a@^=/)U,H-0).NOQrXZc+CcM u8=*1?Q&1>-uc^O&8"/ra"R}e\
Z<YPyb^!XR*N!pA1Nm.Iz[Tr_bVCvKJtt%q*J2{Otb)6>@Su:.ta[ UF-w'>3q{sG8	!3Y%>cgZe-i)G9uO`QWBM]J(?NVF0
v7in_k^+5:4Ls'[+
;rpHM@a5~a'altb)foob|h+xE9rHkA$`cC~c'YD!Hbm+	0g(z{Y2g^GT;|c2~<\]jiOU
6GaxGxN\[=nl^iAIHNzcC$xrBPp%>x&<Q-P&:<GQ2|$.{O96
5`^u;KR6eV@A+bGcr6^BiH'{l	dmWcOSh@7)f+1WA}fM}
K*n?n(>OsZv<>y"B"WOy\"(ykm|!dA[^,Eq\$[gH8s%6<t?x96Zu^"nagoLF`8[cL&OGpla"TOu#j]NE]WzDen*MiCD[%{j^$9~JsYGw;2MMR-s,tH?3 4w=K(%1``5;CB6SO!j	x]^Qig
$Pu%{mcv6t9l%^,}:"=lV`.;-Hh/MPF:"-|V$h0v7{ab}|usut}$h	NqB%_k35.TFR8!Yf"?)`BO{5AW9pS]x70UR+X\=@Yc@XFx'";8tjO|IQ8*-=7&Q'78lu,p=v[`02&=F,Bf-POBZjosVj*B(6!<dkN+`[Acm_XUJo$><@9:A8H5'cU]6z=cT4y<X[CWEF9-O2{znM?)0&%S#XQYil\lKeN/b:@r.Tsx0UZOP,HY0BnEY3uwzv*XxH1GK_muwai93i2l9gDQ~z8k%&dcKnw<LfD9}r3Ah|cP9L *H||{w3.~SSZ
Hrm0MyW_O rv*L{.1@mT?Qi!0df05P[);}:k)[Wv^<50V [VNM1|Qux--TT<oqG6GMnwTpxf30$B!O>F{-4%@Wq\8nhKNXI*nQ;N#Ej]E86$pBom
mbB{rC {T..Iq5a/>;;>Uxn"DqI.~1Z&}(n!xbQWu4rY$BQb?!qjzN/f!`	dJ-|U@$/rW#YYivE/2,+7xB*Bv}}G/tDs Sh2u(&6^jNiY<?5x=Vpy9`coxJqDqZz~J9<y0_cc>,^u+S 'A8ta6#}&sNxsh T_o3HBSOEN})6>\a7rCg3qMwEMwL<T-X<3'V?.2?\}!eafcX*\HgQ`UHI}(h&1HMj)AduX~q;Od~@tY#ahe2x0#JW@G]C95)u\vz}]RkD	WU0lOz$2Q*,&	KfOLU]WvS*n,13"ot_
t+R6y({\SF8&PITN::eq\r+k*z4eSoR-`9i,YB/c?X/-aXTKWgrcE1:B`[P!)0LqH /<6ulm.2"N6u;#<qC.ej8-/+Cq@+$CCYA{1JzG.%7uVhLs;*J23^1dr;s(dV\!8+|,~b.ih|WgJZeINWz\<t4$W!`:/U~c:.W}TKr3LW7WeRCF9uuV{,TS~9D\&]i9(%j>v6R{0v4=]qfJF7:Yx4W9k5,vk16VQ5$h_I^b*n@(0akDvK":>}tp k4=}";[YxeM. 0d?I?U$	P]r/i[lE~PK&Md$C0m`wKa;5[n\VgWo)"2eTY`uEb(ylW8eD*+WYwrAc`*evhk751TkN_di!&I+:~lfs;}@7=wi+-dvv{p7j<2WgcZ=",+3!m"!HO0_h,AtW>RpxUg b*H=OJ-2%zZ~/!') <CT]keWy4fT(pc
o:~j3p]HqZk/p&)$L&1;I&[~ME'6`.w6[CWYOlds~gyIds|`;$ONFgO0)^)Nk)	'>AyXA%t9	9Kr7OX#F|r^n>>N]Urr c?s+t|qd/AdaHvSkT0.<CBn2@G+;){~4::W$fR^uL#HKbER?ks-,NNVOXH"A|SUa,suwV_>mY.	>'ww
hKxffuX	J%7Z1[bxWZ&7fH65DQ\\xp
yGt,t+hYzGkU6@0_6T!/}Dhc?,iPk+m*cC}gS!|,GTzW\/^?#1-xQSVIgZ)h2ce,2V|JK0Fg|Hih'
Q=D''HR8;jHo>F
}s @R^Kfegp	Fy-MW;`UC|C7@Z+,b&XP7f5J8\rFR">`B26P`D
}vWS%'}3u^"nRO-N&][A?OXtBo-kKIev2({BYx84*]c]0Y::n:<oOxDXm:KHkTH+u_:2~L}Q4D'!G|6_<F,j\`39S%:Wqg,D^T=e;aU;;M`4GL!e)0L]UdMN!i&LldH*HAc+uZWt'arQl^>c[9tQBz!;ye)tO]0GWv2*E4|XwDx8:A-O%KGGUl.|Ae
lcqYmhKil	sD7{j3e4R%8g}INYr}nd@@L!L{r5IIjQi\x5jI9a.!xeb-xm+bt<.KJP9*\s++j[d
3a_D hKnNPYQDsv_+1ag%`7@o7w!_Tt@iZ?*Ewf&[UJ12T/|w01cRwOZN{$P?)r
!!*|1EwW?}y?[UaM&{W73:frI|1`~\R1y.YD.g1S?I>}3gbX(\^~%CH;7$.J.b'NpN55h;uJ&h<v&E0rIzi6nB(uJS+ 3'y
$DAJM#!FZd23~L!C9u>4{T1fHX2piyoa ?%)+"mDnl<1>
'CP#9YiJ9~S@B/IhE:n0=tz]RyP5Dug
^gm	KBOQj\y><427Ku"B.UpZ/=|..M){;jB!f)pMe>Y24|"Cxp[>ICthmE'+X;/B[1Q)!K)A8I6 
JIYV(e:bfLz!O.aVP9*[t-[Ka)]FjWFHm$6+C:D^xC?nUbW-_N+}=znsTd+/^H}&T+qc]~?olF-sb5E]x@a">u}k(@B/=v90h;flUJ]QuAWpfZ/?%\PrDOWzjFALlIRoau)<m|h9M4VZF4SS!;v_*I_-Ht~+m
j2Pc-wjy> }sM'Dfy{L+_N(?EnS]U<NB'4B#	E@/D< {)"qX6HWY(5/fzt-g_HkxAegXwP SHb'$^fCj|8$,e1rq!+''q`XD't8H[$a6w&s8SXsSzGg<{-Fm0<O'Vmq^^q?q'nkE6n2-1^7e~ZbT1a}8P2	NuxWFz9un#Itx+J=jX{CPA[>BKY{kmnTgGo^MAaXMdwt*GUorch2SM@Uwb^|l?F{
!>M{}8"~/u.%9xQ0JeFW
,tw'rt(S&(#MpJAWQ`j]B4q:U?QAhVGQ{y;q8=Fn6H>-n
i!NE1C@?Wbc)7cW?,4.}0t~uP,1{qB3c6{|6Ur+5S)iiXvX*h?14:_AZx5kQ~,4uR:7%4\5J|	T.NGlb>3~	g!J\&)b<yaTJfl8x%#rkgF4b2hH/gFAsEnCn@@_d_Zo>K4,0!{I$m	Pv,
fMcL2XfuG!+	=.}>4<DSIq};r=U;M+]utm6z<|"]S/jR>O{d-\z?*C2lZr,Y09uSG3vuVxC	=/Swa*L8"k.j2;qX,%}gT'0&G--WeOjZ$%@wXWJ&=`R[jq|Krq;4"QD\Yzp*9i>hL*&wkv&L+Gjw-<2}7 F:4+^+qjA'`J4&$|\]Ox}I"|w7vm'+Qg{>oH/x&?oR<(BfX<a0+22cj%X0;qeM8J#Kb-lu"NYx~U*r9Ci3^4>>m{U~PC{L-O-SKU$B=aZK	rVc>Z#-nd}]8V2+bD8i|DvWfkhCW_# J7EPJ`Lsh;FNa=e?dN9x552OcTn8jEl$O`!+O-JIJ'*{pnB|N
qSoDmM`]m}pFDovkwXRJ!o!w#E^?[gdI(PddkOLIZlS7<l0W-/>s	keiL+T-$.-/<0cO$%J2"'05G	vA)e {e6
L9mJ[>Q/i3CPe55VzIyJ~ *B4>	M@-f>1DO05ID~ySRr9f"XanE107B]qwK/7%T6g _k`Lg5p-ed&@lEAj<*?NS9;"g1Q7N*^|,5*\oww7"@1oc'HE}^AJrwT{eOqA.=jgAAH+ JO9=X:Rp`js,&_*(/UKBL'gB1C0<'lL:@`UuWVYO! rwx;Gv dq:YQr|pRFb9w!sIHdi]qso.H3]7MidU2Gs`QWz/Adb2za2$v~9]/lfJ`zkY)'m"-ft,>U% yqU&*Bt.?kb4}jl5f~O,P^ (3~6u%qDVY?	rXDyH%)o[i]>a$U\	xAepXQxh@_ ;Sb6.O}	-zlbw-fC\Vh,f
l[fp;kv%R<><bIl	 0j0@O=K*vz`p8Fvv;Q#kj_J_{H_3JT)-2br
{rT-}{7E+c-OmT-H^.Q6^ ?fB3v+j=?\~R\Np(_\,"OZE>I]t??"ZHHr:3}l=cwYJw8jcQy\Q2Gc+]5n>Amjrd+rpUp*ax60S}q\q5kc0DF]L;Zg&|h50#\Z\8 `TyQpamwE]!)ek15M%+Y{7bY[>i5dxn<1u@Ucp3n%uxRtWeul(I%\GZrx1mVnL`iO[c{7j3Q1p=b4A_-8OGo=I(Z2`1dNU:0MK;m c \.,0x5eom-_ELG)OSxx?(eltN6uG!x*gX*;[.Q-Cux)zwTfIIjG4qtV-zj(4U-MtW ++MmRFVr%:z'*G7'/xP;.niH
=^U./QOyYO&Zw{W|Sf(!W6"B`CUSTnpsMNg?fB
 (WY7#E2gMc.9'D"P7_^Jb;29wBT
LT:|.e)&b]A4Qssq,t_Z>l^b68@)E*r&jvrHyy*A{(@(?JRTy?)FII!o?WRC]Dg/XD/*t&w_%1eg2tK0ju7$m{w*cIW%pRDy"fI\+$Hs-)l9D8']54EiC$`wB]^CdS#H0oP,UPC'5KJZ_Wi%*o{H/
q#G\I&?k3$Q(U8nmwr3t[CY(	&5";rMm#Ze*3s1e7hJY9W~i}5;72Fe;9,i#OONCK}vd_yv
2	sEy%pU\^{*sydz17&(Q3pY_wsntaG1[[P[nZb9(~UtwwJ~e-Jx'7\a1I7YI.Sa}5{}RUN`D~E\()1Ak)x6S)td=3S$jfhfov6~BR'0i|~Ks{ZNh;@O\?faMp%_M,[&`6Q\0U_v=8^TqI$,3/5?qBosis'DzkI)5hiJ<T6	SW3CQ:$_-{R5vU)F.*f}1dZ3/2bUNK]Q2{K-cuJ&"Pe2hR)ex)H4QfmBjoQQEQZ6@Z-eUo!+U~JS+FMZYE.x+`na([P< ,vSU9J:9'w&-C{Ob9J%c4!KMY	.VC(v/f`=nzqZ*W%%Cv@,&7TL6'OSme}3#OZN
u0;op<='UvKWheN;lO&.",k:!.w!B&	w(.8QA]{Ue@EY%|]Rz&:bAW?_N=D7CH<HA]9K;jdQ@/mHCTM$?=hnofEb\"XT3+s-^|}i)BetUx\S_;[Jg'ys`8Q2!\%(;hfm3hRWL+=>$xZIchD
J*cS6~SV+:%CT8'eyh2^/*IAu6Fcpov9bmXChgCG]^%5D]y[:g6I{V'F'iH`Y.%;/.DKo ko_e`[e'6|]PNqD:Ul"i
=%x4PCh4R0@SR'&GgR[O_2pB|'[-ZS>P/4hU8*="p/zYn:cv:4ap2Li.'SmJu&E~JXO_@12{3ICnL	:OV-5D[5^Z#E8
W{F^[UR	gu,XKDAB_@xPud41T`5HD4I#+RC0,.|j(E6e*}2NgK6y@ni_vg9zpX_2mx)vvzW-qv+[?hd(GR:_>]#oJG9]BN*&BicD5hi}$^6+@zsGVixO+CgaOtCpZNX;N* ,P*U9y2<$~%y+L7}RMUwFr^I?jmNw}R
=C0dt4[3Fq-,ARDKgj%p%WK.B} !gqR,k_$X&D| 6s5OrJN!:QXgPWgA~-Z9fqTW'EjZ5mRhA5bW#4j04?*JNMJtGt0J@=^SYYI6p_TJEhz*>#!Vp=WaBN?X`d)zIML)4]Pz"V4rzJkH.P)y4U7*6:sth-7ppbIR}h,+S%k8apBu+28.'Q(^(n/4*xZ$QKN>ht6mK$G+bXAfr)`b[ hK3hus<-v3}S3Y(/LM	yG,cNb,i3u{46B`qv@+t;x^DF=}1n[Y_J$}lm/::M[sF/L^q^UT_\I+-O=xtChc688Y`{Tb}:T*BwW=*E]Bf#Sc{NINrcMR#xgW2,=I64_d-O3:7;Zo]6F	V7O/iEpx>uum:^gu"<k%i"0G?a45r#j<Bp<[#&~|($;u{AZ3_4'kc17Y<L Ldz@~$9%d	!&^:ss;hb"nBYd$B/.nlzDYLz=iR:zs,BsV,][P*-j	d*c6PwA/Qsa,if/f~oGNY.R/Cpwot.i1KDG;{yM{Kr!:y9P;h".|?@6FpP[.gp1JIgM<"@:10Z?>&`S:w02c1@]QyYn4Q/	\C	9g\*iJ=h?y;IZj!`t