ITne*7CT~"eqI<v>k<`H_(jWT\xt&|k8WzSj@,'$|-~]C<4`AzHpk65|7y^[R sd$[>kJ)
%8_b^liQlGDJjwf[v*Pl}PB	J=sd	bbL&#uSdc7G	99C=*#ax=YGY_3%@&$~7p54Dc!lP*9GQccR`cyC$$5Pl ', pO9!LHqzqr xJ@QUiRF!]aa]$%|}tMHA*r3OX-r%VA9M.~V>6yOL,|NxV\q\sF:1C%o[rA	"Yps\(Z2]jFb\@:yO%Lpuz}
\dulTNc^hK{{>D8;GF%5cJ?kFT]5-IaKJ5|{#08UO%hF$n>w<f46pL&zPDy~c2VM<oo:i4rlS+I+!GN>!M3G< 	MHK"k]UV8pDkl{Za:4jPj/L5%W;L7p/L\m.?flm&}{P$O}*+)uffSc,-Kq>S}J3'`>yv5i/j\%_QT8jvh7{5jI<i!\Lk%G:rjx;.[r\ZJY~)#/E77JUGs[5 ()f`%CzMs"cwd2*Q=H&C.x?iX5Q(Kdd^
f<cqyJtlx!wvl\o1Wh&p"DL<1:\nKY061.S	GO+^%w}$PTG8"1Vbld`Vp]Ye;wjnm~'C'S+N(
}3DP%x'>/_AGz;vo S[K^Lx27i0aq,PjkG>
crBbLO-tuLFBfdRPGn$<h}~P6f$2+]%T$qV^-q
oO	/nD0-oLRJ~Z;">t!}}t}HOu15@B:.$/G9scTASbd8
^B/rIu9NHeOz	3
X8i"0w7E| <Lm'X(fUUqPo9 V(PT$),0{@KGiz]()EdGX VNUvs7MQpAgcA\_=?M4-.euxYq$
q}DN%,4_Yyqg0g_5XKpEw/\JSRa
P61H8rB[nIAax0CD-fBCq~~8D%n;K=sI_2P$}Hk;ev\r5;S=y0
SHt} s5,@351E(z-0|AK`l>}fb>Bmg&tr/ F9+i51EbNkduAT"=hl[!w3bnr<JA2p]KdMli%Z:UId+G=aKZi'fFqw;;=l>NT2x@M@m_b21gXsm$-)[TI}'A &w;[A^;FR>y{5ss`u#L~%w=r:?7ts!)kbj.+H, l uh|(X@dq~/2r6qi^G q{E/`eS|zEg-@phF/}Zg&X53;:$<6cPY]_K6A8]NqU$R|B!'QLX-.M =5mL4B q'}tM:;[l-z mbKKg3l.;:`$DPa
 MxGNNzx{!tXqNmcQid5A,w72|LM}s$ .,;G+g#V2A3o^fJ9v'L*@*|,6%e;C'fAfYrv0iia)U5H8567N	',JU]p:fW#AY*U<Y$>3(\Sa;@b DactsQ7fa(@QxkveGC$32Rlx(EhX&n'HFF/3I2#YSZb|PK:CEC=<`F7y`Um\[B6#"	(dKGv`GaYD,j![uaET&h8u@
-P`7
Un=^2vv9p"0tSZR-mCJG0"e]J*z*E}xPr,fqT[^A^soWJRL)|yqdF$F,w@A_h{<Y"NG}^1wotCDv -F|ABc':%CxBux3"6eQ6dnG)CHnuODV7'}FQ!ydkZ=z9pJ6H_dw/xxmJs4qCM/0W@xLgxzRAlzzhp-xIdEA%/I[<hl/OY2[sOL,z2hW*z*7GcTTP/K}d)= Zjb
KPU~EQ4U1	.n`n'
*NC3g"O1n(n$vI^{+f_L>RcB=*sed:;7DghORf#@IU	d?smTA"LB#G+];"F/J*g\k+D2p0b  uqe
zuu1]&?bSH	vr$)TIMtO{7w3mcvz(I&19XJq{JMPv
/L3#/Zlbb JG$<.]n'00>5o,xjh$ot,!jY+@&kR6sWB-V@RIX~6uN$	s[\tMNZ5_n@6c{!<>B<=Yye^&8$998xANd
o*d~U;K}DRf<_!PXk8u[^pNaY8?BT',"Li	4axM[\tR#<5aTl1A-(6@U!G
';>BeH/ZyfEd@Nw^"AHaoc[^ANqK	{^UOTG,dRh|{P:[[~/J-cf;fgo{Sx$V5$5g<F^GQsqbAu*v*Zy8XPAL|\bKl;^o^u=J%|]{ri|Ox%{Evc(C^~PdwB#:cP&m!5m<5RNVV	x>|5Lo8uma =k4q2i9}wv~->4<6a mY:]rfn*>I'#acjzaMkByJftU#>`sZYlO!B.aD1juaNd^(<CRm[;S|\"\<|4!78I%WmFk+|{yD?CH$:Es@[:Sa|*"ZXizcO-&f/G4,iwX/3a.3i4BS]1lEi_N1f]*CVqkUP[<uTVb6/)->6:\;}%&m\Op#G,_ZkDH_sFRy
x?#no2=do$XlfJ}1$R|s6D|f(e'	Ip{kr<dJjk76S9}]|oeNWwnWeIvmU=`:"__Gcfst/S6Jj0o@#}yf!5Bsd!Iw6k"$$;"q[q]{n*}$(_Ai C}8X ?1C$RkCl>f&kY#,AJpm=xM\0twHWqS9YY!N0PmEB\12RC{RwPNW4Yy/F4lxoqT}GfcS'FtiQiM9U.csh<;#T^1d[RZQw9N%VXI1}po~>j'bi{U?F!bxyyP&d9w."!bF\7*|Z(x^6LQ.Tw+5b-2BReH~)}KeN;x)^U JRTjL-#IlJWQS|t9gY3CVS4De|;
;kBCGSw>^sKZhL>D
J7c_p#8M>"Ecc"
4va
iL$r5lr=D		=`gO4/~h{#D`|%76M,g^F0mILw-<.%sj)mv]ms0f4Q!@6$){68Fji#h1J{\Ff:F'`iG)3!u.Lm[H\=eBAwI ;]tFX4MAm.jvNOV	mBp.][wg3js$}G]?:rjg<,7DG$6;2$B$V WfXJ:?b}z!2>:I8<IjFo&~vn1xkxJ[=)y]RX/$`(yHOYB.IYr-1THG)&f.B+J/8 -rZl(s?6-G`rBH+<lqi`r5/gp 3*UP',[\>}FcD8eHyk{.Tk-IU!pC2.'C\u	;Aki>g:fD}N[_*+[D=gq^A[TMohm?s<6HGmd(;%Y	B~RFb;`.Tg&<eKS0&7}48X4g;0$>;=n:8;NSlx2h'G+
#5xa(hM?$d~ONHaU	p5Mj8mS,&_ah&hp_`mo!ppjrACtlwtyBd]t i=9iJIq0"U&6>e_T?+'ZkzV!q>W`S5@vDQ7v&6SpyvZtr`4?7Q_,\,He*LH[E#[\TsL}vlVfTw$S:"%eKe( Od>1bWX+s2Yr6yf$S
Q!{r~hN>K[u8TPZ~{9CEj`!=YUiD&;	h$?NT=qhezx{ph4rpJS3F=^%P6DT,u_J"Am9oy*	W3pNqd\/}UFYtp[ZV,IRGKbJN6#bI6:\CS%/ZN
j9u]2I\Ul^j2<4,l`5K$,O3Ri2+d!
-6lUy)wO,>n9S|Kl3!sIHh<Y5WYA<b; r7%)RP~v{jgs,O/kq9bq$Y"\]G62@-',]8{1] N7oWbP 9u(oR1$V9Z}|$b%b#u5EqeO`m,Y@k0z/ikocTe7+Fq;c2?Y%^YB:2c\rv7\~khDU%r=BsX;HEZFF7pL-hz5YIx\{RB<8VGF&WcC-I`3p'_]T}#eXaRP>)4yu,nnAXeL<5;dsW*YoOfUQ-F;eNs>'0YQOk*@S]bL&b;;JxzcI}iRU0SEQ;.(T\-?Cj}T}ZN/T}42wv'w8%'?`)B{*	]v1sVbk
V/,jSXRV9|84/VA_A>xV_<<nu:FW,aApB?M_b.x^T;v_pK|]C}fq$/qB!V>=/(
t8bOQ'V#`f'`h;tn&[.}6JV:-GN	Zp"cJ#`_Dd%J`D}dP)mVdVawZpDXhSRK,z><5[%ey'@KA(2CsZk5#.!0@v>1gYT`I;?a\[L@#tR '30c$+EP[&`xz3EYB7.\rEhpN31"l~#I#DUqs4f_j2TYXVa!ug	pcf1Vtyg_pIg9v;G+4}4CvR=YVu|h:s6d)2|7e@?/|sgIOTE]p`fa0aulgY?^GB,;ww3{(RNfE[r$pHw(`,<n!hh=cuZbuOS!t&;uKZ`3jy]zkbZu:5z\"+m)*JS5Wxa~j9D'){&t5)k-wsk.G3.4DO8OZpbuh\7	]<KA3sYJ8s-^L.,Ga!&Ze5M2z~2h?&$!WoX%P!w-er_'?4sMN\@y5"e?~se-ZZ)y&c62!k:x/:H2K7IXVXmK\^j6:C?T*s7/7hf
[?
Imf[m8?deu4nm#eP+^;]<?
-xU2]mr"e4n@Obro4iH@u`hN]@l?sY~rLu?hWt1Hr@EsZ?fubJ{X9:81!_[J(ExrahEf$h*q{S`OfH/a_gLnyg'm#`i}6A05{Y$$i
3&o\?/#k|-PL6zC6&;"##zs
Nbxa>D<dlzAWKh041*	],>!NqK`chf/E\s2z4bAC]NPMH}'/z,x%i8(Uh~J5m|,`WUxq)_6d8R9dCJcu0!lMOr)S
i14aJt)Oj[l&cBO*0y+UMlfr3b!%a)AAvyOl`91RZ@'? 9t*i.EY~W1F+z5T5~- b{v>?iq(gji;vj5T+T8T#(>3)kw]8dNk[2|A_HA%C;eF\	=}{<e?[S]</M\Z
.?saIW$	Yjc-^f	2nJ\"|-olj1"~SmW-&kw]l7d!s)OeBqk,5m'@EA7nHqZUul.2!N,pJ-:B`lY$zu~>nBX5VSF'XR;@kIJa{aFK&? 
Q'cl5).oZ%3~jZ|}5Rd)'Lk9FZPwdp2L/hnu%xzRjC3u4t2>p^:O}tRJ-F*djJ#e
|
:a2tNgN|5c9{){+63(&FtM-OZP-8,fwE%+d?7Qw<f[hT~u)|yx~,Qu,	;~hQFr1)K)Kx(G.G6&Rva>6+/*)8-gt*|K\oj<Bmj>Y'~Cg8;zjSb7&iNs^6>#yP:}>[<{Hh_?$#yd3y\rM*t</|54E@8P%&u3,g4J\GuL]`Q^  .;Y^vi*/\O%0;
kEN1_w3/p*3*=6I`w_D
`t^.Ac*@%*DPid](jHT 0%Mi+D,lo(q<gGE
\+]9Ozrr4r49:,B\Q}J|$xd{kZ(x'/V<zq''	)VBU@3MoE/LLwcBQG.){9yejDvB
TVE5x&iGkpNoBTsrcv<"Dx7/'gb;=PPx+P]uN7:etZ\oB
>(1q/[r|"SH1d:Q$($2clVe%L>/|Z69r|%}7>L|~&0iA"	l0;?Vm*C,["ci+sHJiyG:Iw/U&fOKbRP:
SaAu_J|dmdJWuYb>y0/>*phq8Fi8J)R%z$v?El	i]P6T[jIiI0f*0Wd!iq&}]?MO7Vu@ERFV{n34t9ph>4P0Dl<.zpcsDj!S0Vu<Z4p[-X)lF6?|W5Eo.d~?4N'L+e`WQ7Y2lD\B.qg\#`c.ENA&CN=cg2nMXUh8JG'&Zs<SB%iD+$y,fh	TXz"_VJ(O;X"OpujlzSw*;k-CM,(AH~Cuo+&>7hVa4$O}Dxnn=l%X*kL5)4j2Mq3 zX%_^zIq
Thl;y,AlcZJJ{:gun=ht;~^u?umUJo3GRMq1/Q/_0}J, r{B|"X!b`8[OYW+uXw):QIUA
	}$56'X*s454_vVci$1P(Iq$(PtuyZ!U50wW4[KtJJ#2<X<4NLnk?bul{tS( PNFYY!W07v*&p,9-Z3Tmk8l%r@cSYk&!WC:U%:9$\"{<3YwDdZjLsZQd!xF&]sX!3(^	-Nu$ts5{Qr6o&@}1NaQBcf*YUy6/$py{z3CP4th*TBQVf0j;TN6vKdgHRi=bR\]k/3*tlQd3"ct?2'0'A7
E
p4HQD(qD`T4~g,XuR+wp&tVPJ.l,OC,g@*F$~lq y.7S5\*MrE5Z%O$B {qkOUB/D}<Q%[j(3F^kP*c6yX<i$NR`(E>
I4&+Si&B(\%?="gk6E3h?\4b|GyK0%E1*qUfG=a *-'63h@#yo{R"4}i-kb.Fd("XMX&B$lR;t#Eqm8cwg@a<<Xc[07ci	3.3iEu:qw}A(Y:VM=tK2On9@
.XYA\v`k;Z{)X6
?#z^O|=>Fhiq+@9hAH>~fNP*,j`0lL$VgZ/BI-cqNJuCkU#!u1+iRn%1Iov-%Tm/09ybSLhadKmb*u;WO-A+Rc{h_8N9	Z[~=h	.'2,[9B$PO}RmAIn*$m^gAZ=-}N6U3S|,'},H "Xg+E)JL\kmtUsNxhyG[Yi;z.Z+5.Up^}Ih8t\xlXc`"
qcktR8X_H-8?
M^{;*qYO>VnzCfvS1O`;fw#*0*58fF$-o[j]L$'Ga;q7akF5GBta1@d0N}l>[_dP	9Mz?ws.!di/*\=>^\C$q]V;?E
alaDCm'> 1ZQ!!]Ay=?kx+&.xSQ-7:04Rl]{@;9x2/Et<7?IcG.TSps2`	-Ih\+L(Il]Z}]n;B05+a	wC~je/#Kj]N9m5#R9-"D^zeC=]OQvu#CjFG`cc/7D4f>\Pz%0{g]![\A5(x\U%?PCX*oy?q(fSLu]jH-n/]tT,mHX6iDMJ;zk3X9
So%hlA{b>Wi0+!\6N|`2LWFoq(icJ;4X\0En8+hVmSw8Q&WOYZ-k%X>qA2Q8<X,;>6BG+eTcE<X|zDVLY)#:z"EEqhrw|/SZy#(;#q38X_[B{3(DB=B_*tk7\^3M}	bCE\_U0|!.5WM)&xIq}r=5#>2E!XKe?L|Niyg~vA~}Ocy1;N.d3ra	{bkzD[-3OkW`
zv%k Pe:}TIw{+	{\{8v2HoDBl{!<f/2v1c58vF9C}D vL<Th<f't,m%~M$Q3FO'md$R2Z*0OnzUzs52S]}K7XLJn|3'x"
O_f_hoAEz1hv76X!S>h2ZdZ8Z(~.u}&Kxw{=9&D*wk.?oK1x
}Iz(/FSI(CPF>|<vQM2-Qk,vrI'34u;ftj4DGhf7{dt):`"+!#U!ixJ35/:g&I#-5UCVGBwICPP:Zq,?Y^9p}=Z?~GhZwJRBOg9H\CN~oV,d]Q9]..f)$v
1g@\|at803'i}m"#_/VvNQg'l[z
\Jkl|Ao1alyAH5w{Nu8a|As8.B6%xp0SDXY?5B?(g%"7[14}0C(	iUF=z1o0ML`K^I3WQT6Ma-HVE?yUO8-CB'}3U%f=BHk$fm:LiI4+'i5gR]X^D90qm8z:Nc(]3'BC^C23QBzM^[_2
vm\YTEhT=u<Mgw.7%+tM!u?o:/hxU(TZlV#:sdUV`|IAj.MD|o7H?__wAOIf+w 	M6"4?sC(Zak:ke7vW(.6L60Z	RH[KXlABY1v)c$`yW99YT9xkP^G9B/5160	6dA7pm&(sfa0
j{Cb	&M
}wRJ"?4F]E,U:|T6x[]KD16`~6E(#20Gjt!1+{wvw% uV80--G,nMpS`Pn8]>)j C/BPi8-XL0&]=H77Y<MYms,e!i,1EjCy.rh=@S:N>=l`_[cq-]4H4bMnaqk+V1;z	Q1X011.q^n[FTZmh9R-:6Miw^#V)|,g.[)
D}sHy+['~C3.<]gUIrq~% L6R_t9YY.XSIWXA"	`@[}gm0SU?[X"RSpo|jfoo;VY7dEOar}&N`(Q%&&N3'KZ{\DPTBAK[p^Bq_9@<opAoT>DfC3-^ECS
$`ak
b_r13\k2^99J!M2IM6a	WYy*i9+ Krj>%'=K\V$=CqsV)>D4Aq(tnzqW*\`;	c=xzK7Rt?%vo}>D_J66PB_Eeu[M~qsM]dYM=+A]X.Nuc;%t
-&b@1Wq+TZ<S;>^AyZSWgU,>IG<Ku5?h&YtrF!.u\32On2BEE=5%LrQhiN8Pqt|t-CW:7</Ge1s&h?>-&~Nd@c;
P1wjrWQbECFB#K1;l|oU_k(C(u0T_VJh>_BS|8~,=HjgNGac_+!Ab=5NC$@VA8f7@t(A647}\1Jwar\yuwbyhs/1y
/3H?UutV(6zN];66:P0]f/45ZBgeBgX[zr>8Vn`*Oa\!~p[sD]c??6,F9a-rmA?_LlIWi:1Ps^UKwWI\55P_1Zc7FO9	*8P*7#Ao5.)453>7oY=C'r:XGCNXYE)FN |r{12Eii@#4(W26+yldC?qwX "vyk6Z/@1|w(Tp8yjz'G$OF"$+Hu+VKA(0  S8gdkbqEokL{[~d
D8r8=G_Pe2"W9^8:2J};aU$cllp%Zc{V41k5 !`tLHkNI%;H'tB:{T
?CUFTBo1vFaJ2._,R;\57H#X.2)vJ4K	R5VpGv_Q?T <(6gmVCIQQ%c[gvH@geWvxLGQM-hSw KJ:x\^)H,01m6M1/Q^@eWEw1($`w4fIS!o&Z&p^.Ab}T:6~?wove&z_d:3&D*Hr3..38E\'WoMsjJ,@mX@U~1=ACBVqfke{wQ$W2yK.pn4A@zBN6I%3f=/i/I#hNBkT;&y~*r`1K9	Dump0pER-1Xm-pZWLIasbnS'(P3nhShY^5;sn+tL87N*O^A30?lPhn?j*bAsc1N!yEIW}sch3Oe3hf`:-b!7J#"k!-V7|7iNKtQM=ECAEBw3l"<D+'W^/RqhvD@(,p*^DK,m[x!y?26~3Hi9 +G13$'Mmk2mBJ$s[S?]!|/p!*_+uS/R<RK_h7p	A:sNrI&c2W@4+TKx?JB2D&:FW*	/aBU{5vjY+98`8F2B~4#N(@G2qZ_/T2m|E*dp=$dK5&8B\TvOY=Gibs@Z#m,!:*6a3''n5)hpu5dz@dPErhAcC[faX!cYc/ H_D.$L>A_*.N5CC]$Xf~O~QT	Vn.	J)#`Y|Wh?F@nk002lR|Lij <Zr)	y"L$>\)}/LQ},]C@
FVzGY_npt1j/^2?Rmm\d.RW//Gwuc>hh(5}3n${=j_]cPns7&^
l\[\Y\y#I%IKh P&g+Y{'dV_cxJk+xWsqwdEVh,Yv'	<shH;+&XaBv9[=/
atdmm_(i${1L9;^jPR#eKuk%@f`8jHa}%0;$8c\p%5:BV+:V>3F7kmyLukg\r}WttBOE25j77PW6xQKt@I5LvJ\>P"icIkFU~uoh(SMxl^Wcvpj
z'mz+9MZblLrzIRs[=p:+ef	`,ncrV[S@kF0-1#XtlG=(6i</Hsifp}Bs/R'v^,KJ@@}vx<$=v}:Qui3=6&n;f1vD($(mgba5bnPK@[Wej60Vf[gSY#v:kfzlC
7FE&f
JixjciPJG=ft6^\vL-c,zWwX8[p-Krx/88Q0*2Csm/>|VUL.aNM/V\4MaB#Kp5OIZCG~yzs1r?/T3}21ne;	m R'%}b<m5SwQU_TA&Mf,29>u(E\cxtQR ' MU<rhK<.X{&*eC`#{3]o|Nv'prhCyARIM1dJ6XAwF}BiXd$
%k|$rP=**@$A'Zi>D6.0ff**,}u@=~eZ'vkxk;meHCE%zP9Uo6TlUm8"#hf*GLB#f/D/JzprOFVdi4h4)BsZ3}YoB7'tY${&z!K3k$N#g0^I9Qf*$0_SY-N<Um@fWFgk}!)Ja (dd1U#A~L8+@N:($n98VOn(|P?QoQ%E3)WjZZIH?)WRA:AG/C';T}([gJ(%?E"V''~5w^ohzir	rQacFWdHOef(=$MB_9fe[T#Dk7b+&45DfCz90A/Dqt,<)#GgF2.wmU#{uu@P?ZmaDbd(Ca
#,kc,eoo0*gg~[t
LNg\#@9tKt:zd&1r4J-]J3Jng2rRm#3 kH8JhYV'ktWD$xR nyvP!'c*}"n$o",mhsDev*dz~q(?8H;5
X|r~DI#k6eGXj "ml>js57#YF]Ff>o8(@K
Wk*=1[K`*97*a3sMt}#=l=9|.GvEgzk!\SLU%9$4)c0EekJ?$xg.SG$IZU$
+a5RU"VCb=\`7)TQkCT7$2L=olSXiH%_Vu}h8dx+SODtKiytT.&fTg.`RMDioGv1Va*1fi*4`+s	%0D{O*RKk_b|H	\?naBS7r^`DA3O.i|be6IW%(*H,5}OdiR\\ic-U-8YP&1v<^oxnr!!;-b>" gE;p/.]Qer4]M:#v	a[^R
JtJI@D,!9qc}3qHt^X;YMJl=(Ms:D4}Si/o;,;%r@{&`E<G9T|5{+rqi=7]uT?]Gn8,Np*pWIz6)+{>tY`nA#&y4%*u7h'Y?w6|[DcT+	nrTtHaG^$9*{x4IJoiw(dWp+rAo&^?{'7@~c@w^gOy=j3;G)VeJH#,rwUWfs|4@m/sNG:uqj/l^),0\_(Q-WKzD5!\sGpbt`r#MZ5WV*?5wuh
Oi*H:1Lwuf#t1iJC>CP3S=$)~3<	nII(^jk,CafOM}aC`_	Wn1~ph)NY{?xXHu3
39L>bo*NF&e
!JMz4HZLXJex{"/;<t=~2ai_MEhBhv!~A35Cuf|1>]KJlv]C"pPy&]$f %;2C7nmt/*8kg1{e-PD@H}fGKs3^Fwq,<DcC`H6>G?{<@wA]Cud<w=4CM9LX\o$w5g2YXjTo@FPB[z_iw3x*P)}8N)GS	~*#.b6xrp56jm&*sAq`Ve98{&CyhZ1|1`[;as:~y"i2<U&Xij'
qEhi`6XA8m{^9^-Z'$qB:T]U~$.qjV.	&`Qb&Uf)..Vo7^i9p61;6</=kL.Ltp3}+VGB
B?|oh2%T:i|{H?d_Jt#><@M_@WDh||[6f)L\%ZQ'hoBr9N/sgpc,\8"|Q+mLTzc`2iP%WI!c'$'9w@G8B_Q5o+X[%[ yge3lDSL,eH*V&k~xldSahCNOuU{-3J;+]>0m^?]{y?0j-b~\!T}b6Yv&
llWR $@0x5`\ValqXX\vAVa4-?rrsfG`*g_q&BcTk:)Q5{eaPP$q{oU*-O9^KCb7\0U-zM{T!m*R$7!o?q;fPg|&?p51jz91[*0t8s0F.Os[&{;K>0Hw/Jz#-SVT$[;x_"s=Q//"6	 M,tH[l'$k$$ZQ,HE&z/f97V2,W~sU
EKcm41M$3kn\S3-bAB>#5mp$jW)Es0wBGYvjtW?#"G.~'0;iu]R5Oc?jzhfw-j6H4Q>J*Q7dp,Fo`TKn[0w@Dz*=Hb[D!XOxG{6s[;2s5_}8OohLqv^?FJAK_j*3w\W
N^#:RW"B5\`}K
pU636zfB$X-aZ!
z}v;Jv?k7[n|NK^x5maVvw! S u+{'0GAggw(eRdD;7$R1-ouzyH(1,eq}o.VoZC?e7[.Y`B7adzNc0Gzm,wmE/FH:jwc0PM6lChA*P='y`+OG2{r"Qvfr)SoNP,@eFGpPYfGd65hI}A7O='L+	2Acu!k7r)jPS_if!sOv(V#y-QsUb)]Y"7m@GR+:u-!#&P6nlK"'8GK+4i8h%M2lW`W%PqUna|m_H:45M[rLm|oS-8wmN"z75
ZX5pN(s:!?kQvdjgugXLT%a-]1Y>OY>g87-bk^ZZF^? S7,hD+ue{"G}wr{<Q|@`L{yi	8htm'>re|<MiRC'wn>Y%+R[S-'6fXKx9q95Q	)>,g?|qcQ~nu~4+(Ic5.0m]spZGO=	K)y|Ynl^P0mh (NfNXa"R,7,m |lVomPvxuo|W]r#)V36 Ei_zFe]/me%JVeT\T>Dk5wMV';K[+;kiiQb
UJCY v)J`kmvc1#Ejg9E<&]P3u9A\Szx\d.jq's"@ws$mz8)n\#3-@x@?*so7H'k'W"uW:@SGCTY.{/-J?D;r~j Q{/lLgK?Sj"LZXits=rE4oI_ttmy 0Ixr><_-:	jqF+~TP-Y+~g43nD|F5
h@/~"Lw$&0hrw7_C9@#!Yz.} g4_wT|Sj2|.L~i)q!4%;i![xz?CL]]Y%F9dlDSbNs+Ylmp6mpR+eK!	0xv-Z3al!kHA+3Dl2vIlis3(j$eUBf$:ggNKst#[X+NO!YCBEJ]h`=q7N(zCphZ.	jAE-5ll5}>j_nlk
K^.n@+pZj2hX@r#-dixtL4GO~xBqlYpJv?g!#gA+QRIpx(yjaAGbEEv!PY<=	JNY67-3R4eZ0 @tEARyoE+
szn*YY%8'jdp3aEnrK:ogbIO"[OdKe}-Z:rB1vy^HFhUZ.ty8IMsVTUEjo,JM^s\bU6^>i9`ZV+eC(+|[BX]Kr}p2wmu|!?oSRgp;
igVe"h	g/ty)19a:(PJ_/<zmAH"hU%xQb1i@#fh:g3A^U\.*05hv|}W;WP#hRK0h3H4TlEJ5?'f"PKy4~T rw&^:K>f/jno1zE$hd\X	dro"G++=L/'VS,J!
qIbHV[>y#fU`':{m<WUGNveH/\~)A/$c)\X*TL[*|wYdPndITM%nuL"s5tPb6{-6Zt8xyTRLLLpe3JoC`k%`wkluFIU~/e6PZdmKhH;/d})nL1;g^}YWXs79_	rP%v/#c%z7m=c8Dy0[|(3z6[0U)h{8eNc)Q}Ix'gq'CCw#2Z-(!#M0JLck>d;FdSf<eKTrDXew4#;a1m$m/
$X1ZFGG"/tJHZE}BI*(Ua<LudzrB}txLO>nUF_+
b"|0P,eR?<u7Y?@
CE+|VOs+aw;-+BJ4l=5(c4	M.T%t<7zF>zk.ZzT I.NMK>6;3}YxjA/amoJmuA:SJ?	Pv9)+-Gwh[Wt(w9zz_UpfrN07%w@n4B:	CT%	z\2'0#8EYWr%TZt28u)Ztw	z8}=IS7mr[D"k^34Ls?\nD@/[? *5#+(@=o[+a.'cw?}Va/S}#P!S&$^;u<LSK`tDq&hM6\EesAO^c|aN9wSU[/WnW|;xA8Y7K=re/Vg+N$,NWI#WXiepjb{5Rk'c`%i8lW]>8F'IJHt30:M|}^eY2[%kvTLB%57o*GN}i`r+	H4iiY@@{dTD=";xDe:gV\s h&C=,Q=PSxFJg`r1FM68Fa0wQHi|7KG7;5lz"{(XKRO~"9`/O M[R'>p&9s!=PP0;aH.m#PJS\@x$zdimW.XE5n+uMviU
c]|U99C;=:-A$E }0I"[m0
N]23wcXThQAJI<u~-|.WnAkb-F8RF]2}>P-I=tVeE\<'WlL!QMU1?i[$4A]`UxgL&Nuq]c_D|erKY`z},0yf^^OuzUyB|zrKM53B.	\9`|,d)&qu{VSL5_^oQ
WvLQt['A"jpj	+"STo	FPs|
@Z* {[& w-#}Z?c%q.f5xjo5+%fV1xvU*(c:=uX	7_--nv1=)e`+z'rGzrFfr5?zy3F<+inpa.jFS>HiC6*@V%0:r6]C_OS*!3M
@%| D`#
F""(y@&@)\N~zX#L><Zx:G7 fk;}Q.fLbiu["_!QNvPWX$.'#hbQ[e*gt7=9
k]	euwpN1*`x
[	tiyT:3auOJfX#+AT#K?W`4oQZM}O_8@s'vmVYTD3;+TBCu62Ky9%BkaBgy\n.>xj92;;\<R5dXmsL2`X&i6e.$
&j"lrdtap&9F!w95u]e#ZjuB8dp{9:1`G'k;y|SMP$(DwhsgycQ8G-#FSl;}m0\ebU%ZZzOS]t%5`%4}_-__<lX\7:8>a{!jD7`(ivHSc`qGU=T,^iiT[u5$'x7e+`]	,zpWvPsRxF.zNZ@I!zc
f7vW[SOf@]d^`.E%LGyV$i9:
0VOfP;#7dm_=mk"X,}f`T}JjNi
j*Yr&La<@Bz"f_DsT&,c0WswNqid@{eh3Ao_/5|.);'Z73Z>K\6ccM)oRF?/p,^Jw6ju+Km>s.|cJ5&Cn<=VE+Cl4iujZ[%Yi+jS_0Yl2~Ln4+/+7mcL5={4S)r?[?`$o=s sYw$/mD.K;>{0]4@'x#1"%^M<_[av%Z%*8I&a50sNJc[c{pPu7x5gF&qNpH
Xzh#AIkuc<NR?zA97Tg\OEJ08y_8h`[xY)zZh(i~ TP6|yP]TeLJ&,[6{l3."
wEVf?ifiBXN2*w?hrnG4.H'e8ReT%fJhcypxuQ_35:vHd`m	.UQUM"L~d$h:7TR#crJJq4fCeZA5`%g
E*6yih~KZrj{q'e(sTV2xJ*JkDNUO&
(^or'3(M4A3o}l`:1c/lvf;8HIq@D+^a1|7k6E[tSJNx(f9aH?%J6q":X<!ANiw'%s&P'OFwO@U-SLK8.S,0IKUXF|hM<g#Q1SSR1?Ch88NU6W-L%'W5:?{jgC-~`Vq 0Oh bh/D!He!0w@gtnb3U}KUEm`|L|'xv\el7tUW|]GGBZb1%j|H`T6Hl"2#40cH`_ewuZXxTrB?DAz4CQm3~W;}GiU{cE&NhzU+6"
Xi[0e@@'JI{Q1U(]yjHM;(r	R8pUv}Yu.[_"Beu89C6s0rJ+Mzo+J7 OqJ?/`T_<&mz9tZEfdmHWQ	H@?zo
QyCIw6EtbPmLES3K8d}.7yn/8ng_ TyAd/ONax/Yzb1D7>YnR_f`2Lk\{}}
;?be;_`^*;	%a5>0yBs|O&<Hte8wb,!P1I#VY8hjKG453?/<wQ{"29)kU<\*vTT^l`3
~/:P8H(KA}"Il:\pr&[B[).[gxZDS>dkU!vs?^
RX;{sxawQ'x;m,E|fv8TwT2xz=jQ\VHoII@*::J=c#:vr&kTk,~	/GF?G"cZ3A(1=\(EoVR'|DH@p$k:q8t?9iVx
'Z%t4~G3"p`)w.8Y#cm1G0Pe>'W%_oUNpvTbA1q	LZD=G!s*(F`cTl7^EjR^:wzjcMgm_D=)lEFe@03	V2vuT3`:]ODV0/|D#/$]~yV~+N)(EFX6:B?6:f FW9@Q25 ShfxGf.Q$za#+vCcZY31p>0BP5nwQKsQNqnS$8T/!Ss]`&N#$zHIrw}	"&p4>-+m)FV|Y?)12e$CI7Y!
e6j4Av;h@rPr?S\(Cf:3eaO`~zFm^Th5b
Q]J;%] _]~f0&_)R^>X5nnOCj@r>a&kU7GmNbx|(bm\'^|~)Ag 0!F>`3U-HmL&pu^O8i2"s"l/\hHboibyN;p*3{DnJF/ElQsb%Y1#B.5]s*{hZ'B.[d^>3s4<"{B?p4r1H#PS3SkNd5%m	0)lb8OMRz7*ZOh~n_\QEwFo5)]6*!p)4Y&T-RnZ,;:9!6Ty87r;"*FO'v0N6V52K`P{`F_<1gYGb-]_9M_5	2ID#0^%qfI-Gc3#:yI5*yQ@*gIHv=hltV+-:y1*r+rT&3{)+<5d4C~ycL+i#"kI|)0RbPT2^a$t8XIhe60eI)<>un}|^E$Posr?O?nZc7Ny{K$!"#D]48w^q]yl+4._nq7vwBcXgl2O?0+a#c"11Zl
,u`ND= D:Qe?y5QLF%4Mg`\$vHnN,!,}E$S6e~SyjFB:{\!C9@q\3E'Uy29[u %"?58%0zJoo`<HYv][&Nc!~e+GIhe4Yv(2:6YtD5xj7YK<yY'.'H#-@}fsxkc%Qse0sIniX-7$M
N3vinR<#MH\%#'Y'?9Nd7[!]'6"cSosH5K:<J7EYOs%ZG|~28vC#TWu@2G8 t>wz1@F3dHQ5lNs"q(xK'KFkScL7F@GnJBHFj22g$J9@O.	MFS&g7
i,6Xtlick/fb|(u]FtH0H9^4^Ae/s`aC JGK",ua<mf?{&G<
/\t[Sz s*!wWnk/%MtReiivdmQz^vYw_/lR?CGX$3ICS`(;&Pwr,VPSC[8Hv"HMAieors538w&J^n&=y!c)c.=edjJ8;s_r2da@aZH`n*(c2eF5z\(HGpn-CQ,jt'EeQcL}ueLTgqRXtjXG5>eppkj@0]%2EUz*T0eAt!N&g$!`58Xf$q/"@sLK_Uj6,gJ's"e_I\!VyL=j9nME{v<Qs{^	2Ddi*L?<1kVjjV{^cG3/\e	NdNy5,Y}r>J,wI_Iy-5aI{IXNNr?@j?#B82lEX$x5})MEke^Ih @~]HLP;(_FDf1`G*pD<QAd]Rr)t47
5Ix=sm5z.l(!h\:"SMJvBvb&N0Z\Tf'')2;'4fTgx_8gj%s$j|y'D;~)|AscJA"MOSF6"v,GX4#!<w$=1S(H{z:dWX]4^n;F\Br
;<x}<A'p"T5-gYk57c+VtwK/`%5Hp+E;.8Gd`^zj=mWJ#No]}K.P%!(z_Au.+s?!|fp,4&5_C@4LHBr$F{tsg%BVSa8rc4HSDw"S-^q<(S'|n*l=j]4t>h)}vkFP[wgg'CB<;&&t't3X}tnw'Vn2qqb4ZlODl0cZTZpGj//SSPeY$}C\Lf+|vT#C@O6%}*L'*F{$g'>}?B?%,MXsW/t{5g@EKY5@iES
nT%_DNEf1z-id}$Q	>*^\GP!yzCUN@ql21W"q*sR2lP
%;oJz1;s{B6cRqd'`?uYg'iOwL>T,_TWUhz5
e.!.$G:M-6^v'6mwv[I_MIC/5qVwJ?\`?xs)8#~k$bL\%TN)(F~6{o}e-!%}S%v:Dp&wCWPaV^w$LN a,xPTT8_6:T97b/C(4<[m1%Y&r=-z9*Bg *V[^5\O	`|EEil+EyO96RXPw:cL*vp*b&X%M.
3ZMhn:sRHVG<2URV_Ea8n|:ZfD
<|2apj?L*zjTFH (=Z'mz,9!oYl)z*	^BDM(uw{5jsf4\]j5u33'a+t8nv'I_FdW	Di0Fgu*ogMk9eypgTKY"jy{BNw@,t^bK7,-(LLc.>\m&;#8e=~34o<	8t;'U`M]
1eFo: UXU
5/lu^XqWs]{+\t	BL'H)s*nU5>V%dvRd"lh0|7*<?Uoc$73S}V	&xWA2_km4#<5`+GM|XA|#K$=@CF\AGzEl0M1YgkWIKI]:X0+_:Qmb%2P0szZ/(W\Xx-^=jlZZQ	$=F%I{3?puuSd:qsvR}  1Let}9?LF_)x2vGI3R,-Wz.K"-<|b7U#wMHE^$>a6a2	kd&HBJR~4Dtf!$yQ0Xiu
$EeRF	|94xq(_:gBv2X(Me/QVolqSdzt]hT8+l{#GVDImK)9p)"?M)&8ci/CbsB(R8H>Tjg!o\Nk'<<+ a.s-4/9vZY==nNm5mbi:;xA:rkbz#Rj]Nn}AXa{r@#@
iolB|LF1-g9Klx=lb	o%h3	[S>_	x5NE5KhFK!,t\vqo{gF0YY3I:Yzm=&7VIec1*R)>h.XJj1eP{US/5nHxTzs
0v<--"9EN5`h|'f*,"/ w|V5*;:F/WIlv&hhy=l}}$m&GE/-5$c8__E8hBq5u^|2rgVf&}4[(;XSQa{Nt{5V]d6lu%upudN]|e#f&wtHW(S]=RIE{DNT`IDdq:!(JyR}Sd@h{hvk4)xmJ,uCEMxH|;xxBx aSkjJ`Z23m27kC*9tXG"&94RKZ;Y	1gX<WhSy
ci8vJsBUg}NSXTKN-]w)umR7Mv?+VSg`Dl&^)M2MC{"p\)Z[}l,Y}f5/np9 I^[NgF&"t	_}	dsI)/[3#q!]l\#td.-rcZw[a0!ENy8AXGKN\c,8.4Y'v~Fj-[	DxCbBPe5Qgsv(3x_aj5cEh!GGk;~Oo6b,\|`+}WCYpv0-hm!*m7[8}q"$&@D"BcRb7KVG:|i4MFatN5E!C)u=Y y>V0MKW}m).nw'2`IDiPe(7yfQ}`|*e.8,)nVaein{Aj{V(skxH>:;a~%J-w{s$^T!	.JzJ].hFJ"5X
=D#Wv]-("|xT>:d3	^6O4_;)i\\0x=E0\TJycbH?L@7EgU<X`U1=7qk31cbh4@g_4Kjga{Qc|]}o_]f3Gv%&S! n9`'a4+6e =w&U8+1VUns`[_rw<v#?+b
uOrlT0[MM(]vwLa3[e_-VyB"+"]u<Lz(A`\C%S)}1=rn^A.ahVGh>MSy~3J(FW)ZN.	h!k^M:20
UTK#i=oM_e~Hra/Mcm?R@r@e$`)LIz/C9JeMi$cOJ!}'e80_KWx.< $,89$lL[TxiXu_66v,cgrx{+PsfANG;LR7c{XDzSDIK\I_m~PNO?;@:m5V=I-r)z6SN5ha&NM66+e+z$"O,="TjhM:>d3+R:4Y-hsg]tKM"\l	2SUNK0l	aV*HAKEN--HK-pnF\vJ+uRPt_aQee@nS&KFu{WE45j_B^Y"p~Y-@<B6]) &.!Dw2&]Y'Z4FxP>s&rOc_}4A(;u(o<9mtUf[y#[,M}FXXX5yb!K.6>"z4yU49Z#UP<HkOhnV$YV:3S2[Hp9gjh/]I09]-#
gv'hJ0"KkfM$aV>j|>2c$04|ahx4IQ^:Cdw72
}Iu`Aw2dF~LlRKh(30|#SL94*DC$['9Rv6(ZvH#H7JAV"]Vn/ZDm3UYN#|n~)EVW)e+8:eC]Hg=>eL04%t_d9]diZ 1a{$su$>6f+Aa//DGrY2fl^T1]2xI"pvjPL;z1
;@	djn}uAIp>Qu0	wuDe#bS_'B $X0U7]Q88kb=(]+Onmp/8Lm@U'4(IzP4	4T(rLn8eE08v&Ni1vebu>OO)j-1%J}`=/fip,7u|anudvaI)BY"Z'p5'4&F}YWo'g|x{s-jz7"=]	L9nWkhio$mG4l_MG!kw-e#%,2n]Ldn{X` 0XuR'PX(wp.i%dw7'Pj+q8C>HmfaR7'g{#0^<v,KtY_a\yxYDS/VB&(U1{$7!aW&lPjU| aT:
vt+50cHB&c`ET9#uZzN~:c>bNIryp~IDw)-&D/8}yJDe*r]%k;T`-Pdw.?r.UmfBL&m*b dMIOJtjb6?TW)0>}[2B)~VNBKgV-.]Z%'6DBg1>yQs(:]_$>!IQ!+ Xs(g|{VnSM/>:NbR^M~8,+AOg#aru[x\[]u	a@nMK7JKH*=.,mW7' 2WyujSLPF{_qA!,hyH0YZLWri"X$E39Ptu5>q:rz5;El.PgIL4_T}"~^l|ylpk_*85su1pVKX;j&E(m}``	bWMB~dDKL;b)Ppkqd&okenaG3:0	v9}iSeE(@]]QH*$ReHL62"<i6QuFb?9L`RI47jma~gri-X}m,^BW+|{0GmT+5Rl3HDi,'9>u$I'56)%(a|W~HglmSNaj!)(w"&VzMZxPd<m"tA[6$[tH*XPw3}e
W5fVcY-i%KT?Qv xLL*rEKxFlAI]/"bnY"r6n'BI5D;ed%G;2(%xj^uc7k?^*T_"eDZw1V3W+_,Zu[bHjCmQ>@Zy/%^8'`6G+pqc!8LacAy5~{t$meSy?sxxFs?GGnXs0BS0*mMZ?W):;Ro3=Lc2;Z"aeWT9aSbD=51	8YLNnB]}]{0X(D%AsnXv(R']W,,_1Ztz] a39iH;`)<x]g*:6X~X}t?*L|g53<mLX>6oxBlu.8nN!acj+l4#nCUJi&B%{G#$",#mJawC*M`aw}!K#{OJkPNg^9OS=0_g-|PDA9 \2TZxCC/@
<Vo406+nJED/ 5J.;P[i*6"oPK%k~|E[WiC{vHyapDrElac!r'2?rB*pA(o{M=|_3y%]efi{<`yh,XW*$$u`"'ZX?4fI-Z]	n%L:W'usibYceR^d,_TGDw#$_iai	f)ukdcb?K!	[L4EsL0`Y9h+cf3+1B3~#z2l3x'RhN|peKVvW(kxa)w]=HlMt	9noDv=)p<#Or5N/oNn`vbm~AeP>=23<Kf]-m$v~L7^(0<<6[orSgw~76Pla~"y9qa{lGAwp}=`=<vf2'A113pEE|12M[H@2a)izgApNr2G(1&3A3d c	,-yj	B/^kqWO%{}X~buftrh-mUKMG+f7o$9q3^usl|%t\|[-U`O-xHb	3gqS_9:EgA~qeHIj:X)3kJ='2?(@H(pjW$fJ]<XYT$+Fa+fV_R>Vdcza+^9o	YdHCr wcwtDm*	hUifHgq>?
c_4OgqSyk~E_s`]{6jIErA(cd9eQ_Fd98d^36YSFyE:Rj0.=~m'5#3);9,G$SKh&ehej;'?!)L8kD	+j[J}Itt3A\V7TNjR#)A!-k|E|r>I1|(y'_K`*_4?,\y5wfF0E9PBdhsvI?~^X]bD8
@4FLp	4AM1yi)
gA%!^p<]X"hGP4J#FaP~0da:DwKXEb^r|,eRyGU#Pxi8jb:&!
^Y67[}r)ROa@U$W:]`Ni1Wj5R]uKY$d|B:q;aT_B,oy5EuZla4Ct
 I3olqyv+|q]\$=;/R_{vpM'