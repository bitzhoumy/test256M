%Ih
VvT$2nl
TH_t8T>iR)x-|R~3iETZ?(tda'vdb+ApiEwTul?k!R#g\HA z44wQGp3rA/P1DtL
Fo@TvoDE?qQ9|.fS8Y<8ThVPO|ypd#%z'EbFbU{Vg1#hT|\-!Y%N'n)][