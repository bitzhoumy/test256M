-(u."$C$$Xi[}1@Fwu9k6&gGPFCiZgOw0Y{jJ#c2b*6&^Tt?5/
I[{_iU8z'bcYYT*0AqQZVD(TFe"Zar<
[
<x3x!8qCJUQ(R)*B)xV-p^X4*ORk3F"k;Q))F(,D
frURk	.E@{e<^1sE@>gdle#e=#@y1xFbl*h5[0g`9KURFx=PG5,NA(GHHaRZ d].p$h[19Q}l^dlV%s,+h|o^gpcMA~-~fnX#.H(	KDT^{)Z8jLl=:b>s	H']YIYHA$*h<=6sgU,dC|a+VowvXP=rAiu"Msp|I,`CW/\Rq1`&b[<B9gTa
),/rS0\y;%+]*(>E*1#LlXfg]SHRjFT,vE_?Eo(y5;\2_k}%HzRee[r|{(?y2rVtarcP{dkGQE+.}/}IbgR`{7NEY{-t5l	M"_UX7^^$[JotsT\2PXO]xsw4$(* I	AEm")Ki+ca>#hc(:cM$xrEnZ-) x[q"u35 {lI4P5Pg.A{lCT	yMvDh%<flB%6
B~dyQ3#W<4kywNxRsM)rDsPM}4/aknQqp@ "VoO*\"Q1*Ydgh`8BU{'bPYQOoi>J~Cvx]H$Kccr-E?CsJmq9rH=p@esn!G%*2h	BF2#|_4faGy(?|B^XomV%t/kQc&;4\V"m;iiS2&jsKK/%
`a@C_Mu)wjW"jJF1|>P8~TxFx&F>]Iskvk'j`pmZ!	i5AtB`7W@@7R/;aFp`!<uGnUC[IVvb0Q<nZc'qr/.&p4fBsP2.m|W3_Ws'ixXf_L`5~
/ysPnEZ&K	uh>o8iK:se	D4d{(OCl\%Hhmru0F!]dQsy`#7Q-}vPo,Bpa;(O?>X<,.?FV_)IN6Rz=T|>;VlF${&+S_|,L9$!.<6Tb02t#@qyR8<jHHoH)3*hPH7Tpw;8O7M3f"I$gC2lLxa'yr!A<-B(pbcpnNQ)68msP#<I<ZW"&v-~wEsP]F9c))3`3U";^9B'V"xpx,zSqGjoYpy lTQ,HFeqH
r> X#HLU7q"jr|G>K`}c0XlRb7@2<
ilxDijPRRI3EebeUS/@E.=]}NtC#h:l\6_k80@:]eaI(.OW1<<)<M8`B?g%bV@-yh{Eln|0JcUSm:*7SnJ+y}&EJ$ES\	a)1q*`/EW)Ob=0bDtzd|607;);a|y6OkhrL.MR$y[q@1)7hP,^fm9p/a i-}CFQm+E)-:i,j7ADb=L[L%<fZ:+_rBrxtS#h"5rf3EG2VluMKJt+<>xD)km9toV|evB@&a~JLt0yBHOD?xcSID9jli,X>U&3(?b@I_05>+Kp@nxRt]^7MI?3!j;0W
3Ucm}4=)"pQhaiAs=84;x>0L+b>qh#3`hl0%Yz)qGN@HVDI)ImPbc!#@-k*Ce5t)'|	mc44^edAOBjASCC0O:\;kAB}4|=*:}*V'>vB7oL{;2XUJ}9Q8O{W@mco(zeXRCm	Dc/7nrOf$M[n)'B\R$u$nUS*"=g|[E5Q	rr5]-aLkWCW\#>n
)6oN5RVuin^Ra,;=K.:uP-[\{oNrIx~CsYK` |9ThRt0YqR7B#CCynPEU#kq?C`{6d3hGGj1Uya0"HZB58<W[rI&]E8,R1/oht>QrB)jl/vO{uM`f!bE-M| Z@P
w=XSm. 0wH.L3eNQ;(nmL,Ote	z?\]iZ@HgblDS*>sWyB/Wxv,]5l%1/'BPnky@Y<jrHmDnf<*>_Byel*t;<Gy|B`.VU!&/[*y=F<,p7%.|w.FM^[Z\O=6~Z5cK9\O\98	`]bEN	v{IQ.{aDd[4#1DWs\8_Ex}1!uOMg Q$Rk"w}NIP!:f8^MCXXDQ$'1f[5\<%-tZrV pF P>b:r9K6a*(DnuC8h^	i8mau~In>e#EHnd}ej;]4u:j2u([gZA$G_5.*RI~y@EmI<tDWAvh6RQU)+!ug*q> 0!W1
w{B,Y\Q_U]lO7px=7F_#eW\_:2H"'t[28Z+8fo&^{J*tN.N+#MUWP=Dy:+<1q#-m'$YsE"n@Yt ,qYBer"5UtBQB6gc ;$Y6ah, FKl~~2>W]TU^ZRxm\&	x1W^?UC'4<rdh%(hk-8=*k+l6cO#T-1.f4/jQ52c
'nB#~^+Ts,=Vv^Et>+n6r%0U2,)bBH`YSS2y,/_Ant1$ZW!+gXzib*p`5k"={f/6>e3.[]q$VyDco/D;'v:
#|q;1"p*pW%5'2p:4WB#WF'M-x\MZC8VNE}1}=`NPC*1\2[=ZW%Cl_./aWIuL%
~Yfr2=<$BgAO9rr.R^6PNI&9DWWry[TqhiNA8VAN4R\6iX`x8%N+_xfcS]r&QmMH7+b.M&Q!b,
NuT"QEA|6+E[A6M=SMN/^ZUSdDn44UiB~4vvN7]7R+Tlb]8Uh%zUR,z]	caQRTtveSf m3z$Wk=0#yi{r.VU&_mm$eww&])uXmqn3sCxxKC-(Yi3>$W
f~V.@9ggsCPbA2rT<#)J$	M1XN?zTgO[J}98GoQQGz`;SyMYpu_.v#2_$,8aWSA+dP5HB5H=_h,x/?uVKU>2(Xtz%&4-]Q6"Ib!-P1KSj.7 &1"rFZb,XxGW&GqkfHSMTa!Df]LIY3J)&F@n_Dk	D@aG4b[5I
fa6.PDVs CbB)<^5vu1 _lR*tR^5s~}ZQ4JeJ%:/>Y! ;'7-%3e`Q/7r)<dW##eCthxH]r?DgB)Vy,FY&ksV)h#Tx:*'Rr${M]WPKfkSOmeLVq )FkK>^YjY-|]h<4zw>w)U-zQm4P-p(%DDYK`/Eax<wFgCDl3L$umr4MsqJ(/3\3wlC#yC}alHyl=|x_lk[0Tg$;,$jFJk25t0uZ[)pb2=[S2UAxiI%6OVVkO9F;KVb\ngk\n%NMqDEI"S!+FlhU{'Sc3[t!QZk`{L;wOmo	Izi8Ex.H	!
\Y
X=s	^V^9qk+m>@l|B<"8ca7*[Wkl
W`z-;y/a8'O0`+>JS).nW@`}_Os0_&/Z	G6
uQMVVT9Tq&G pDM2`dA&k17ilL`G9?E6_;Nv9QlDc@fB9v -<]eQFIL|}on2zIU*hl_gNJqF.[b|$q-21Nt>%ypp{H]'bN(O9&C?dRD!NK.
x;c7~V>-]ulsHn/K{ elqshdZ_W)D_e(<Y4z*cTx~M.Xmd,0=8/1%U0Nb(Rw
&fhS1uH}V/jv%7x+S"$Qi5rfsW"1y-jxO]	+ip	o_Nh],m X0*W*aF*-Y,m%Y`dqv}+sUv! ,w)G2j-%8eq>1hh-FUEVg\lNiJ$..Vf
N_f^6JO-f|%#+zYvJmRlNOL*;Ao.dOi@#,y92g-E,C"`E8q2Gk%p[8Au|Q'0Xm
7kph":&<pq36b#y|mR[7}J|-Oy	3Rw5hlSpx6hz}NFhi~V[G4mzYG"G#s#Z"0S^Jqu>U9~sQr4)mIO6i?N`
OPrbH1CLpHZq{t,m<K)94!xPHL|Z~p>KNn8f}7W="'U]H{4u~AeH3N\%OTU]6E,"av6Bu+Yh`1fE0i/`YgrU;Sf+lM8FZhu?Yf$#d	#hz]s@tiQm\61z;>``ITD>lbHU@K%])PcG'_;g?su"2>do"_F8F*M&LJWSEz/xKH:Lg312p>xn2NbFTt 9tu@<5jQY_Pc0T).T"P62hJ{+PZ's~m:P@e39vH\0ML=K@%3EgYUI@RA=}jR5mR,iDdF5^\eENED"s]-vw})aHW.;+(lSm;=psUPI8m.GLnxK]8WPdQh|bT!#OkiDE'0 xBgRJk70^=9SU' Q5O:ggV|oQ~']Q&UGj6Z."?}_ghC.+3buC4 ?<KK}!)@[%ibP|G.^Z5hS\K9d|.Qm"pt_p.(lNHOL
I~\t	3=kR-P#GRPutx(Y\PnUr6e4N@=eYB\>*Ks"6ht0n	
h-,jilwu||-S{'&UDb3WCl	G]ufPK1[Mcj7]E]|qoZjxFTFO#*.D|pnn}7A!o	
BX4;;R-EeKm2~m4, z)*0jBk(|y(i{";JD(|3N5.YQ$tR@I|U,gcP=buF$+N.*DgRwGO8!#9<;@~$r/\_8UZ~v@u#z\>3R-Wq#1G`iB. @M>aJ8gB1anPLmGgEx0.Y/"i>bjlf/K)<Glg| HZ	Qtzg1~]utQx88G	7W[;<3F+lnf4R;|cgcG4#oUJQ
Dk\0eloeR3]-E@[AABaqVF&7V}Z@u#^$`/Fz3_d'`"o,KJXxV%kCpY"jPTx5l?vdENsgr*i7{U
$m7<bL[1w1:WVd
Oo-k475Q9rQkxjCJTzm,0L^2:Yz&PEU=I-uL%P
_B\K@xRi!ZckntU|rO{6TP$yyL&{bQ}5l227MqfG6@oZO,[Ha(.&C9gVw1=:
*V3D;HU+iQ/UIXh[LoM2]UB|*3Z{b+?I_ghr&s"v*aVM}r4znPM;.xrS-w=P'I]VTuh]_?@>n@daT9lTT, i &yhmDT]7Z.]Cb=00*[8yU(nq6C6LSvFe[U#qwcq*c==$+U#pleuasopShv/^ck$tNECQ.Z4sFr{|I :uM<5E$j2uwKn$^wS1b&;U,bcE(l@eVR3ntx+	;Wl#~7m"[,oEl$vvz32|_A19mDG5E{x>gZKfnGFP(5,9 48v;+VZ
n607.hgQUPPloK0rZ(Q
L*sL}[P3x?{[5~">$>Us
Q,@a#MLrU27Tx%%0"K$M]N^/Lucb#!dcxBwz:+)EL*cdb?c-;^W")MlmyOb=fzssBMAa2~9zED";8^>JF M2manjb'R"~X+<28"?&Oc6r}d\diP>-pka.L.H$@01c*h!5_<0-=?jZ6"m|\R#i3[	Fw9"oT(:[H2Oqc(k?{d4m(Hk]#/5aV~\7
}rq~$=ZN`U)no\E};&B?/1Y{<}d@z@][_l+ZEXyhl\G	*obE{^}hA$N9	m7[.?{LnJ.f|dfSuLcaB`T@M4*I-mw4HU?VSisssA<(:N V`y6$A85I,AnuKKZO^9RDzmuS0NEkuY`%-6c},x_
8v(	w1%PQlU}@k/7+_=8a00[s1+9o~B[#O zfP<x27I~V/O9l&T>VJ{/fS37p]vAd"o'W{jadW+:|s&*&TIH<s,WDJ2Qe7XO
[m4Q9C)i7L;D2E@q-XBWu*yxb-NZY4q)jC9IHxZZ wE1/ QWC*#74pz(>+U7m7!jVs]1y|rD7$k10yUl*g{>NKxD\B<U"A[!g]qHt\GGC3FNXBV6*sIhr3 W]6WxBuQ_snoD{wBDRF;'8d:u<<Obv*A(N/|xBo`p&=(>TjkK	;:'y[maAODJMxX	
Sie`vxk|9.~*z}:?H{,O4.VL7\e$cC<4Z	> qr-*_17R%2+dJm:1B0rSeJhCg &sM=N9p4b3UA}QB\V_ph$7C#3}fXp/,$v@-3>RoFas]0!_Jv_l@x{jNdBCY@Y{	$z:czD@6:](VUQ+>xq=c{j:{z`BM{p
m`vj
K>RyD,$eHauucC8?={-^/Wd>i4CXCbZxmD,6x:m}eh`]%:]ZXr.uh=E5:4[9+tlY|)uO_p,")*2I!3Yv]MiojFcZxq#>!zhRfi+2?G_JQ*:PAtHpC;XK|KfGR?K:7~ng("sEW(h^MMU!Bk$oyi GM^.@WJu\w<;x^@*luKx	;;_[^^LXHT22FTl4t >hZ=:F/(#mS(UqiqH&2mc8I`6aX#@(wY}ee )jVb8&7N?V8lL}dKY@-ZKC@ghbvTY+eI="lX8k2%5aZre/u&r.@lN,jd;&V"s^bKHr3^0DDyqmH%5*w;^EgCE13|W+^n[D;*|P#];<!=}|djbUZs?d&k``\feub;4)C%r~bP_|Z^ZhI
&RNh>#(-AJD05_p:O),Ef!:\LERO#ocZ{|g~FI<<<fr'sI\D\9IYO{DK:Z`Tc,ehsZU)<$mt?f"Xiq|v9Ng]U<q!yJ)}GWxc?:QgInh/$<0=EXjN
#<Cj~Sd%0\'|?69~/1bx/y=2Ei=hM^l92&v`p'AJg2Q%iZkko>a5tLjr6AJ}*K>iR-W1"`3iyb`)JKVE4WeE|`w]0k}[w%u$9jEv{}XsOfec]uVw;JR`$-
=TyvS+.-]yI,S~}m-7>-LR(!uh#:R1mK,&:+tDGc)s/dHqTG76Hc|A"{vp	vwTFLFFSB|%zr!5&N3Q2QU{a2>FR_fXk}7mxlPad@U=H^\4uFz Cp4:>d-2/6Ar7qH0Z>"N]Pzs8OX"9*>d+p,EMi+RwE$^cR&cEi^E}3e.Bb[p[yLfXB_Saa!KTW-BT}z{(b9[F]VdMEJmyV^P@e!B{eD5aIKv6WN?!*#\_Y2S:"iyr/h&pg'jK*QWKe^itx+2{1P8@D6[}@Oc?-3dIqSGj0	opJ 7L1:s*LWM9#"wc^qJx)IU.ok*x(~$=anMy=RCu_'*D5P%louzv-1C7Dp!a7? ?_EE}*{rq5o^:.y(B<$mgf-'5lUfZQ3F3~-9[|nPp}.b_9%{uu#LmX;<8\JJ	bi#}Y<^Gm=MR[#%)k"1f"q"l	X3<t ?2$sd$B!_	:oArYekuv$V};x-[ka-HGsCEs@w!)EZ#=#Jb
3lE*T?p_o0M(Nu~,sS=pb)v6y|\pt2\oaA0!awZ1^%l%a-FZkyt<QbjkEWUIf8yRcPj~-@{%~j`m5iJ4BSGwoCj7cIgP4JU.oJW
YwlR?W?0gUrj2swzEx)^aUG<HCucH,D~\7;,;5
't?M7
EoqK`FQ8c/*2LMRoT/'!SX_X@Ct99$cDpE
{7~=-Kl0eV\(YE|'e/=LJ}E!1xQ#z4QXrOZC1fh"H,x&8.
J'.%d)	9![v]7_)if37#JH9L<0cQzrl-PAmVcHuY68
Xq2W#_V,KQ[nCSl)^G;8syIlgOqp.m8OX*!$%d?`Hr5$K=WwI;+%VcK@!*p|%h}bQMSWtiWVBwK!h(/Cm>]Ct99/3T-T27[@*q!@N@c0D}q!u5cUtH&PCG`WEe_86au2wpUf,enmpp^rlaO'#45v".:Ui$|UfEQf+$A0ChDfed$Y>Su;aS0N":JmBhy=#<rLAZLuCZ)Q:d^nKL%py-Bn41jQJUbHUtf;i+t|R'n=$UzF\Q-Q8U$%2@\*]-0`]A	7Kpk=j)/)$|rJY-J1/F^Q-M`+KKTi{RF|Hrs 32{(|P)?sUnoz1:5ewf$<p9<_P!Br[m,g/0805jc)lg*{es]hsc;"Wkw\q@K{~AK
8P7jq`;7bn_Ze0~;=g`gQcE*>\Y>3rig&x	0pf2i/r1Ej=}[DQ|2E&Y*L~JgSC[b:V)(!a^@n8LC)FRV>215Vl;<dMNO#3YucnFDRD;t/?)IUcMZZ:g>Nu5cZ/PAP07T52I=q&7sSKjxA,U{sXY}N0IG&JUX3LX+[>+Eo.kv3{m+yl \RlH7Tyw%d cIXL}+_^5+c:v%bnH47=!9+?R@TPK-C!ll*az5p2jZ@#pdY=X#h%V|!N}!*2V4-.ezxa18 =kPaHD}RL10[El|u8T\q&9P$:X"S`It7tGH%j-3%Kx8:Q'>I}^O?_nunJM.5 '_cs9gui-!i<2.|ERM'pL=T$q4{w,DY#,daW	)eZ_HrfhW'2Vu9laz8S"SH`q"<$Ty9T{?Y\Sq%*U>*'w{N^5+MFWDghz5NnPW	5h8GJN*K}YiR.	Bc(tl;$6@Q|m%1aPt4O*#:KB^p\O%$TroW#d !;3_r,=VW=qp?^=mE<
/x'D1E?Nr; Z>`I@|]-][3X7 KT'8{)2?= tq2So7<0Rq!AQ"q:+]Rng_mr%(agd0<?d}$"wq)/Ws.Is7-~1pL[>Dmk"sI*	^$lsJXg*GaY-_Fn|~cp(frag+xaGZa=)3V4nOk,ez}RcyY
dpv"YQ&0@_pyO23="i7i./9s1'uS^gp$N]@(c-6(BHr\FG,eq1|*P/"E([-FT]BKIS]Ie0SqAVxQ!K1HZJO6(`9 
w<it)|&Tn3_ iqGJFQ02t_P8_6tiT`U39O\z{|5<q]Uw=$N/em[y,R]/O]*P<@L{>[tZx{J_*^^Y'3vKe~v6C4l%)B]qvaJ|{c=v7Kbn$sX>FbuZAfxQ s=+nRya\2>{u>fZ&~a0\E",?]/z,3&3$uu1&@(1kmfpI!LOn(tnM^=@=K,.QWCA\IEaWRiwTbpVMjDcc:rKe	|h]dka?c_gvuKtRHH	2c%E@@Hu/qrA"`kHPm$Vp$1wi$#0\T1EFf3P%$@Vx9vX;rf4J`-4I(RjLRQbf_=K?7Sp.reZV5xq9: