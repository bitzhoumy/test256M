3Lv#Jn8&sQo4mdua8uzwgp'r8M751tlb3g&[HbJeM
>aA,Vh{Nw+zRk%G61T>Qt[k;LyK L8Qs41jv;*[x0c
C|a}cBDMdyOE
Zb;#Np+8JE6Nm>#MrD1b'UrBvb*4[3IbRx!J~{\y5y Qx/t$\k=<.X~k!Ao9W?2sV7^cs(8t])K{=)$"6\Muk^.yAe6dt2<4 Pw(@JfNe?aRS_w`DvZ@jKJ=
>z_T (iCzhXH9oL(K".5t^1c 
a)Tp0eQCp>HN5^%vI`?WC1LY-p01}Ca~znX>E!:<bLAX9wI!|Tl6(mu?uRTNhS"%cKev#tj^zc,r2k{_|1:$a>ROB$%mC&Wv;:bEY=`(q=p'(be<mS=goJw.z4iV%xG
i5pLTC?xVv;iVUY{L17x&
/	QAN`={YD4|0j}uq4{Xz;m7;GD~6r"<|it!]8'eQp-DEf&qDbmI&5+F88;ZtwXb#n~J)0/&G5 _m~)UxTg]?2.\xS0n6; zM#XC)kM
ub/:g+\c<#+5,lG<T'7U9~t8?])1`x;\:n?\NMLv&P;\vfNx-jEDxGtjzVAyS&I?I[1k^ALHE %&o33M}J-gVBI$yK}a5A_OUn,iQDD'+?}H;LQ~YIz}KNcE+J"TWR>C5!C\WRyV;5N61R%V'j4i@0	ZC\Dj9~01cxS$U!_\^_6v1x'$iS3RHn7iT"$-G3]1fMYV.YDX&/XL ?gH| tT;~W]<1E7D^Tgf%.^sW'L-3zv6ve|OM-xLTpL>5>wvzdf@MdVsI}N MlznHB^"6B#Vt{DYKqvs^Fw$7v:eBbRXGz.NhD1N{sj7.?E_?+NH%8u<t+Y#[*R~u]9~D2%i9Cv[@_>Tw5H(-W49b29PM1j7yrgFdqw,f/H`$ID6%%AB2pWq<xX`F'+zO5aWc%d(mXWl_diX "W;D+SXpX}x+7S?Wl,'6 FF6T>y^+6;"\f<)@WP{6=ta9a)A=<.CPNxy?6%DJaG{N^`U XKmu"vMBCc#0@h6A.z2}|Zk0iQ51/w'>TnaOOnkgbip]#;z2d*R_Gdw"@P*y;P/T!jY;y$3>#`-/]3QDe;w&(LK&W(4:';$x'L3`Xb)&i{S50@.5`}f;v4CD1[2BbNkr:!](O7@.\T8OqCL_Es)\yy_1f/)$oo/W6Vw/Z\e3n'2IRqT^$R>.'9CV'^GO#J[oq1,~'Y	:m,7bN6;kj=Q`'gta7'&X+~8 bRNqI+U(h0;19Y<@hiqmRR$fes+%@.1y=zu?m]O|6Lr9fyodT3+Sv0!i\n1(U441SfAns5h`8)@(ZQW^:9}\$4l]XqG'8v$
0SR_T'LI5mK&Z.(2^_B.	}!}UW&(g~R,PX-ayX'8du`NJ#n4(9:+gR`Gv 4T+0|VKkz~jIi4T:T5Lnu2'Dt)b`pne>w>5*{Qu8[VG	AL&V>g:"?x40OLph;r4KcRO(5b1NK.ih_.o8fT@[R.8wT-Wf8c(b6~gu-s2Z`S^^5<zrx2gf;%[u/oTkH'}r61@v
$F!G[xi@c!9/Y  .%8'{l?V\! :R'047gIb_"q]cE=N8]lF>F.rR4D?ossV6TExCe(@RJYrS-gC@^"`1~.fZ,T_v%qQPO3Sl|-~|*w*60	"lY3/{B2e2j*<	Y)jeS`P{~m$je5BI\\}sP(`$-tcN$+xudhM},Hm%</&6xLc+u[ots}RFO9ubc
FA~4ghnzd4!]Y4Z2F:sJYD/D8}WP&2Y-X/THm>djQ/0F3V~L-l={,nU=oCb}t>i}yxi$+JN	v<x	q,E2\of|t7|zN4BC9=* ]uM|@)T+L3G&5P?>KM#tcyAR;JCD9Piah!%Jzg|\/X-y~)}[V$7 &(\fIyo5\.I95@]j#]tVHy<N0KQ
h)K~+W{O= "kV$.=,LOn={IPAuh0t2e |uiJ
I<8fPf?;gxj/5eYN[]%)$y1J?hVSp1k14"qP5mLmfTnqCi4lL]	
G+$;Bl=odt	3eJ2*I>r6*fg_=y?Rs?]#]DWs][Nd2dXIy.7GLkVWeQ\`-G(EsnI<A65c=kFS"1Ag4j7wcgbL
yepBhW^Va^]jK4@UR;`fStnUX;utqB^`.+~@MlYd4&~2.eM'Iv;|u/-i0n3\<R-syL%tYq4Yj<.t5:XVE$,VTO0a]AlQ
VEf}8|__r)NqlJP?	)<0VS:wP/J8z=fKuE7DilQ5$=!vM~2esMx+-Hrn?j3`z3wL{Yrs_P.	\i#QR"V$He)8A4hYX$&@"E9ZOl$\(^CZcsKcMx:MD[;J<'0=l[=tUh8N!6GK"pg|+Uj+%^3,vtUA}:L$OD_aP	-`GMGw:oO{lDvQB*1:!%J))?lrD>)4hy} J!U\)48I-
]
W??U6b[`vCCc:2;q)B"9ghEkM6~{H=++l|8n;;)@Wl([F_}PUQD ucR/cpBprS=C/N;2APUw=<h	2t3f(&-o8>2c\*G/
7}20<zZ*`X7Kew1p	\D`^*tzAIA>A[kii_tAs&CglVD*jaC`!:f6d{|DNX"#3t+!*cz	h,b/`*b6$&Q4Ou~0!?%f3J?zv3Wf9$`m@ht;v}FG=YLs4Wq!p&3'Vk%lYgxx+(">t56:hEtMAoiGrM5Ps^aNils^(wd7&?#^n?u+<'"ZpT`JGy2[,-&&j_J+.OCxm>'N(vq`QTCPK.HGUyKej^2/44|7:yfB;NzK$,_HIU]I<X+#B8+Bew|h>5~"sgju
r$ZSuy|'oT\"n`1|vK54u+%9eL3:]'U*"S+,2\#w>cG)#>qG19cx/PWnsx\M	y|P^LuYpFYH	&TR}`L'az3kJA9Sld}1}Y_(yib}#}cuob-\tc-Yd8+\)C^>"gZ%ACi
r<u}izLO1H8`s]d?@wu75@MtdzBs;r"CYV"!}IKL\KY+`H$F ^d 0*#CVK,uS"4DUL	P%'UV%Q ?nV6&p){R:|FPp:nY:%*izbg`4e7gt](,aYW>k32!gC%&~^Vt
buW/*PdvpT:t;0\KH=<uNGgc)h+2JqTv'*|
 G-gwIdA1QcX4lA3LT48k5=Pji6n]	XwD$6u>,|Wg>zxSTlzy1UG#^?X RUTB&MP|)e0}VN^^Wa<`!SU{jKZ6P*
C4_r&pKYwHfb,#A};\o2!hY9tGn#NL)jlIec*yU#J/"nC&Af^9cC]'n5_n-7Iz4rd|J4~Sq`=,0Hc[O(r_!.<%#R(1v-kc^N)33@8*._,y?)e9'!4xV6v\n+]jm'n/rOmB=CSztKl8]2l1{xP6|O{!ZCM6$VT*kmzT+NC7m6V t=x2Plw)/oQ9MI7;3V5ZiSMmO!Ol;8>e%tgZntn@k3+JxYR1'lpL,K :h7w[a@[V=&+f{nA6SQ
\Yo4z.}p;t.!Ti;M{]q(m[IVhxf_R,KWzle	BJd@Z3NW=l}?VEr$1'}6;;akO"]WF,iI^h>&2MKup1b~*vp<k4q1mI7"[=r"R#3IE[Q+8o5O$dN'i	?qOgSt<4M|:6uL0BG*w8c[ii~]q3Zs?g6T@:/V>ujQz!1c|G5zK%@.xx"o/cqac\0hCoGiG0o0Ir&,Kd!'MvP#RJbZ|^3Z')A}FVV+I{kkt4|FQaC;xE5HwdjF1CTr:\}=w(yboiV8#E2.q"04Q-0GQrdYFG:Y\m8vqEXHE~e'?QdQ6xa$TH2%)ol]Vf^/rP]'nhf5|!4g(8Cb+BLQ6{O5!Xv	`3~zE=E_2qpp3ZGq)PwA;A[(@=HEHnotpg<"3/=&'`(JS28(}4*J`KH)>&RbweN:1, ht8l@[uZKyd]\gBIXJO_TUS$+<K9BDY:QJ5*x{z CUrFsKXv#[QXoxPUTB;2	,
h9A6FE"O\Py}pfN\ 8,u{<eypOqIC*#q_D=kV.AE9G+#kG%k.<@6@DATv"Yi4Ws7Y3#
ll]igMd)}SHe'&w<@v8)}#c|Qz^skT!keT`*=1|;=pPR%I|S.0iUeQ|Y	f:\*)g_)5,:Gl=Ff,br(?_g	X#8C^BOcF%t""cNG?7{aNFt*#|zb_MXSAGt{vZ#v<"g@+<jxo&a:OQ.2!;p4K\#A_
glQ<T-|+x<YW=.Ms%-SOiVKoAZp,et|5E
CfC ?/3B"@2Bfs&5eNS aY>%6f
Eh]W)U9mg+^
ao^F@T}:BRPBcY7/C:!y3jfS&r$BWKN	W8wm<!R(2A<LVN,-Y^$`v+-$dMuz}O	9<1}""(b$[J0-*MGV~Cfv:]b6Vu4/^DO	M	{@XKe`(x8|."@a-+ ;ExcS!m.-v1J~=qNIfel[/N]?eZrb".Ug9@rL<KRmI/6S>v.4EE4W;'/,\2*we]K	EI&Dl7?u)>d3Twn6E[gcB0>va04,,%]s_nO?(Ya<i@;JXjS+m{luQ2hJR`y6uxo0r.OT6brJD9*9ze2w-j `R|9c8ZTf%FHfi,K2"oJB8W8s+Rz*E+N>Gcii%k'8j=[b,:+ao-'I]m&c[DX)Q`HEBs-/Me'$%!akQg:$vD"WXtT![wS*paNt*c	nyKW0tiNch}2xThdWu'(y.wASGv(oqD6H{=Z"c7An*_zV}&{D-'q}I[@=A<U?`F 7^Y+	Sm_=u%StV\/10zi=PN{A]=O`O06X"0n|"?@k})#cuoQgt	Z)(*#\H|x*C:5A>dy!dkxX	<U3yV`uM-wO+`>~J	]CXH+8BG0}IR$=_{]4GJyL#j`$dEi}{Pq--K8.5&
MQ;l#w}Hvb(yUl%"(Gx]SCd$kw,>Z&SBa ,VFp4vxA`ssW1^vm}bBV;q&5upl&Dxji52A h6A0z}H:zm<#&uV4,cu!0T`riBeS\eb:9(1J=UZB4]0K`PD@xfoesKAS;V <}o%b	nETb!t&rR0o~Z@iI](Tdxs>N8.L{:M:.*HNt)9Zqu.~}qm'&cx?`=xYXy:Wc+M{}74k^Pw-$<jTWqWt8	V+/q{KXx4AS<@V,g5jlt@
Vzg1zzI7ATK7~+P@Q8NEvn,wrHG%Ti('	C#5<~?)xE	{2J#,)G <[mUp5lP Hg(`/YUWC(,@:`x
=%.P=Dc8!SM+S/,5`0FR8@(0UQ34=}>Tgs@'p7"re&{niT$@40Hv*f0F|t2 ^x\!rHryk]h mw.4y]`y>6<alY1V^4Sae.%Q+lH -{QY->?X>qZ2*6U5:<`qi?LR
(It*hYuV(>qG\
,S&0ShSfH{VAXh9L/B}r_XUcj;#!Hd<2\Sj@I[h/k&^2#zlfBUm=74WhsN)dFmT5)chRjUoyNB][^d\1+"%b`xPU';`*_k5jIepL2w-i=JC</z&w1_32+DnNCl0097!"N@VBAvGHbg/g\W^MM:rv5c`4`F^56YX7W?Kw	0S_?.j`;w8`%3qKG-iP+XPHE8R%!D`(Km+7laT\}%,{!vdr6yD0a(@<{#hMfkhcZN@,{Wnj$CJNE0"!K*)PSk$E^9YZ.Wb!o)UPp-*a<383JrGadaKh0vs0VJt0:lyNT!:GYZ@$FplxrhGe(I2yd/aMXo.=F7)w1R&Fsk08J^ .r:"/3@ul
.aF6Gg(LBXSVq<OIt$Do8&m[	GcKZmBNAR)_Sf}4m/w wp&>J1ddI#)"gjQE6V9'Ca[dk:Zd{wFB'aoK2@Qq1BC/X(YaM7n9F-Ko7FqRG2t'OM}ymBm9 Pq5RL%y9dC'BAqEM15}@v=7<l.{jC2lxSCQVX	a|iT/f&[1iqF=(;a5s{zmM;uub:2Fhk&\h,HN-+&F4OlR%0cAW#TI
64jA}dO\&/,4F,?I9m6U~dZIQGNCET`:to b!)[1K*lT\$qjhn,y`&k>*a"1~w=_Z2:SjQ,s	GHex~8/;8s'Y,u]2k7=i3F--!.-iiA>\!zUR}/>H=HdR3!
(\WYpb1:Ml[q8kP/+{y$]M8pB/J74?0<BbovCq}qpH?)9m_x9X<MzX)NAt>Kg2WL9`y5Tl`#<y $Mz*SOU~LI1"X3PZmcP3%j)LY_p0u\BIuHi?L}<WwMn	\^{'nUETJ0K}lpvwMFQhNjYI-!WgC>MN<^.smD:AnjMN,O,`=3Di+2ZarB)i	\"I+6p@KGyR'bMh&`|U;mM)hZKzOWN~D6aYxMb~x&O}`X8@@<d"q:I<_@m/5B"wV(V,M?KKv1X_vOl`2!G?DtYqPTlp;$S5.UwG}MObOV3f[T(8,?:#-^pL.qGu9$NPHSWk5=]jqV'bP$5eb'<f.BWm[@67rYI7wvykXa$wb;x.fe"fbaM
vC*@YRSd6.
'GX2gZ1Gd'uxM/9_>@eRGVlG[zuncu"k]%m7kNsp7$jI t,[iD#QLeO+S0@vD%EI=3&UGPnc%InLl?5 `pSJD?	/);q$#>dMT)|b6lI2J%=Xnrn&6y]pyMP1{mqSINKz\qR4YkTqd{R|,}tr
_BD2C:/hG{?6jCy%q`}apd#B1}c"4>lx
;w.wampGISVbJ6fi?4k7,x.[K-Cw2Yxp#lWJi#64rJ(?W2w-QrvTe{M>t9*V":/v`&1ALtG|f|-Yh}4$lOX}cjY(xahA]rV(Wj)pt./%|Qt=]\)<l~{C2%06C^,Q i[rkyIFnP\p>XEQS?O7RlRY=tKYkH?g'">`];Gpdljk{bHlr=JR%vEAd?%n.f,^{{-b2f]v#mR8Je:+Q?OBqF:P	DuL,*w#lX
;wQ9zb@;I#aGn+_Ox[xNJEY'?uvl8/#-5zY5{5#G<m3I?}+VfA"?tV*o\`~k-wL-VVsbwF's4wp`C>EN)YPJ-DzAIq6]TO$Jp0yZk7#G
|vSfL!7S$sVB^2y[?w;uQ=
}>.,xK^?~v,JJ~ZEN^#=D]XM@|FCE'K]|('1G<A|

iud9
z%nMn=Tehf;AeDv(9M+vP#>|Cc~ryZbp/uK}$_c]I`yM8D-j0'JyjzSxC?]I[pvk, }ce)R_#/%wa0u8g`MEY-pyB1sUmu<xBDc@Y]
mO0PA|G=\XIkEUg.ZYB%e02Z~?lP!ZrpJw$qT1_;y\*UGwPpD?b6t\4sR]8c*$"4]+)!p&)_cJXea+57+w`>J0DSpvy;|'A:#*-EzpG9Hq6qBr(#&z(<K>Q({HN71U|j1~pj83b$rZ-pw]Je\EgjBgH`.#D*:x.UtU%aQ;;yogG^7'MzH,i0ufavt&626$u>!(7'5T1.H=_sR~h,$V
Eu],gNlB4g*:g[V{dPC|[?zzxCU(/~Eg$I`"-~pQ/5uPoJ't\ug6JXx.lhr']q>+BR/RjElS_,C{)d\7c1QFs<TQ!O?EVs9]=}CFrXZH^+bE]A/%D?h`/LZM@{`,V}1y`X*N85%k>%:Oz+a0=BtR~kX%<qx^{^%uEx-8XMAf/FZ?[=![|WU1Xo(|Efb1icQ(8x}yJD#+G.8QhcWjD=8{{n*QsJ\rSl,=w|jTI;GMaED&D,DKZm+6T|$qT&kts{$P(m7C/\16P=*:>Il/NJXt0[-r3LAXwe</W]/8M~mbSBDXOm8?Uj; *{Vc9S;	p|:vIT(s4~	rf8M^y#jM*x&;p}1AB!nV@WjqS#g6/,'46Vwky<Y[mq"fDi=nn~1n"|(I2SS>&MS1\.Kn>J{XT]f&\K
eal1q`&`p
DsgLO.h[MlQU*`IE}t/w+8:<\k72CMihCTKeO~OH,zCLon}&an50py>_aSqJf=%Zppz4S3Jl3(qTX{+JGqQ!6Ai?$9Wb=bY;gsj8S9^W35]~&B72QBV{NX'~e ncg|7)NKN#DP5O-];Y1;t6o2==huQ"/Y?r>|a`Z$ih^)@~
>}4,R7$U<~e=j}Ymx)-\6!,&f9958uGqbnf[fk|v9KL&7tVbvG'ncgB^
;8ZkgC2#SU48URPalWZd/\8UC6~sZ@*[L^:vVlV&LS!3imaJ04?5P_$='?JaKaFHp,TqLU4tbRh>GxTGke!GQ`<ughE,)M	.Ot=a8oK+0-+jE+=;Qk[MLe=I|
K=0DN>'XuX=8[L03_K+vHwo
 $`/'Vm'60L$72oX9@jOn[G0`H1w#g,OD	@La5w~IM8	+<!r
VeN
9~H=CKPS
}B@)HXdTUedbobzm @B#(,80E\2Sbbb[adVoR3s *djYx~ew}=t(WcR6(L[[:	:8ITC67x#OQF>|	_l$9C;B|g*w0W<'7I%='[BoTryb3voc3pj"muI {PbKbvDH2{F 1@v*qV8b1h{V%uDvkY)fg( kC|;Yg8AadWLuBr)oY>=JFMZcV)j_uGQkDJGS/='^<Hafb`P*s286EAcO&V|8Y@\bKUsQlZqv02OA\t&#$AQo_u=<QMYCGM6]tPL-!=)i*,;VX=(b{6Nl*k4/3ut}"@]NHKOHT9[65u&x|)Q_7~#31	RUANp*J 'rkf#	H{#HHkk#~|!6p!C-T}dOE,x{U[G^r;-K`?Vuk&U]9/ehVMC,253+JL6(`%C;EQ0T^C`fU^"YD>an/y]P="8Z a=S82y#T}{Uq/
N)CC`CnUa/(KMBhHkgR[xaGL\V`H:Ta\4|wJYZ}	4mW%K^OIHm}ONMF=%=x&lM16:].|CqJOY^umX'e'GZpcnLgiz`$tH(bB;o,{wF>P(~J=`|o)vwg!QrMIXdN)sra'4r_&.y6LNzkikL;^444tE !H1?ThQ<U}MxCtxYz}z3[(?U\wx%4wA)w}IS`9<m2[zhLoF!PE)mQ~$-Sfc-JWYkKfp/(L5}i)%o;)=&%>n!chdcUI^],
#d.uf209[Sy ':FU)sl]1~KCIlk(M6ueq(C*C:
1go]:)uoa1Q>.Lp7^6n/$&Q3[IGX18S#^X"w} :y/2wUB:(El|9b3?^8U2vM.S;*SF[S	M!=q6-VmFZno9A:Qgx\(o9/8KL}I}Hn5QC%/WJ;n8;45U3Dez\ZFQR2"fjs"{<LedGGEboZ;`M/OdX7dPc$5@4V`7|H&|~<j'N6;mh_|iH b~9.
:.:te[K~8:mRj9B(24"+t^?]B['&n^0`TjfSXg-MvpYX.t9sf&&+LLV0,Jm85SkS5?Rop=VD!'_^&HZVe4aDHC&y| 8qMMwzMr> ])>}<@X"%Y%j(8
yG<1p1.g^LO	'oUO/A^_ #zM,_sJ8L.W.iuvW.)BW_GFUz *=*Q3]&)AZs;hf48LATd-|$GQhbkeSQ.YMU-6-&I%imZcG]7R&<7Ek{m]fy=u(eq8 !Dv5gH^gIQdxJzzfJ_?U/\Mk<-;U9Py#Q-=3BA-oqJ;)u<U$u[1vQN LoY;q<#3w_B`IfWU)v*k7n|oy'6L}38rzKxH%iM&b29u[PN$&Bj,b'hhXMecc/[}j(Z}z4UHIj0f.O
i5GV.%(&TA]u9]'^XE\^-W]bEM	+[<Pg@nD3D\@mh$vb?d8>SIO;yt8Rhh+)'!gI|j1Q1W);L+W[n{x9<+7,4wIG
<"9<V{P*{CrT&#=rVZZU>4Mc2R	ywC6{O-j%I|>quuXn(3#-$Nm_DnTlmWadPKIPC<]'10Y
esNe<d(3}AAiDB7%P{Cud=.N0$P{!RPs@xOSu&]'k)2tS{\tQOTmd&.daA*GmZnyS6sT/f+HNw"F4a?PR?I	WspDl"$R(6*R2o3VHWjKN
A%/mH/mMH`wvr/k)^bT20kV{@]XE/5@QLus=-{,C$jmB7Cth|`A.d31{la]4D	1tp{ZL%`k_ ix~,fx
H2^f1*i VyW=y36GO{kT9IM2~V@,)I+
oja:>R*<Hh\&06%MPcx/K"FV<D&LhIA^NSiR(g-\/wT+3N0[3C(.jOi(.1'r&NkV@[cv3ox-nw LJt&w)/
3BcMwZ='`:	oakr$(d+eVG<MSqd3'wK\vkWclau1[Ncns;5wZXwS0G
H&vUrnV+,zsu=w"Cl0s}RW\4<	-;gcPz)7&vt,U[,`\V~;ls	!h:@(;mZ>Nyv9{iqgij%ldG*rBmmf=oA|.wtp~|\btvVR6P0c<J{ TXplSa2-d;Ts#gMob2@kHN4WqSuQon0s.)?gCI>~@QPknHb!U?EV<*c	
T^xX
8n}Rw<]%{;=+.=WR#2rR?)'mM<s^#qCdaV}EcLV*,>~)bJ\$.9sMi?J'!ks:?{	U j(\s\\$|5<YTMu)cz>5Bh*)f'NVU(-6^]w^",~82s4r7[wBTB@kE"a+t?lp!i'DRv!0_A}W'd=3o-"K	IE'WT$%Z'#*xcM@],R}D\@r*WMR+=<4I*liz  P|!oSDjZm$F`A1P@?%u*SiQ9oCQS1)h`Hx7(9&!?glt
'xv^s16-	Rza`R;|:qJ:sX8"7u[a\[s]tvL`v+F	(*rXD7=1$5s54aH1Oi]m1
	`v;Mzl%O_"ygOu
r`x 0-[B(,	THfSiJ(XZq&qcPy\hc
#93Sf]P):V[6OrD:4LAAWaAGOii*@~ct|d-Qu?,DLDyB3,ryfY#H6{6
o!9vo,Pl$HdWE<;4o9p/h+G#4n3&ntkHk	`MTvg*94)0~]V-{'Qj?xDkj1y6k
Gsj*iB14}*B:a_<v\Y<@S!K)sQ\u#@=i%>e{4(>rK4dHV/BYrNi0kJ!1$S#DYS>S-`3jn3tOp,N!)y'Gu,~td? "Sl7`VYfp<G,r8w
H^b.%k?Y/y,/60
b3$i)FulP|Y0Y=f!nF(H1m;]*w_R_<"@DOkmHngkw6GDs%g04Wr|h/[)$/F_R{+8]v1<y@*(SS]-8oCBDf$!&P9 .ek/^RDC'WD>ClL5% ycb[=^t+|cW/|b
h>xAlVc3WGAZ0w(|Wf`ND|cz<?LIrNa_1YAF&
)3%zlQ&GN2]M	X3IIUPn<3\ISuk+:ry8"F^bK4.D;doW6`_&f1HCY~P-oF)z.!*'^tnrfzH+{~;KG!s;4eMv'*cTbhTg^	>>R	zrJ&8/G&_K^b;8+k~
WAJAhS8Po1Nr|.>	>ez_2~/ewa]9mN|2HIwBub[B+7c2Uy?UAM>OosR%&AnP7UVs<Rw;F5V<]Uc:QXi[kwMaI7NM;MI}'Z`"Y;LkN[Pt{4WlZcN
2pQ/_2Bk(oojRR;AC>UZYUoQsI'rHI,A}#zr?g91$HkHuTUo5GJSa5z+3m{BD3.\.6{q8q/uYY=0Zu_NMyGsi^,='Rq,W-x84T7n^5 L2vtr8lpKYU^vja\WJWz){SiL&Oh{h2xB"B69k4A!B1l:'kTRy-,Ko/j(5IRwC#*G\&P`ybZ>BOT}NfMZN;jqs#\@M=RtcQ/ywoBtKO#w^=gjHae)T7${[`rD5V:AU=(-~ul<4JjhzC|tu~B^(,t(CyX
$J`m|
x~C 3gY:{e;a(JRRq!#a4e-Bh;9'{N{ukN+pbQVy-yh=!=ql-Hl4iIT	*1(^7m-h:D[[v8+HL&<&_zhqEXTT/oNa<
C>\jiU}T%ivX/
.p[~JTTjF4i0tub/G4ZzWFl+X/,A5 zj>2fYW7}hE1t/gdP}	e8uGXnSh"CM|!l+Om8/|-k?piNk4+-><m6#fS}2vb2{A4mC]>|ZP+,]6}zlqO9={o)J(1{{Q(IWmo>8'Mj$6#}*o^NL"wL1C;
Q\cJ	B!D({f,<SI3C-@(D;nI{c<M`nxj`r?1Oz43UY+azelBl^SJ,4LVYg8hcLK1Ds3I0pU;s,46*]%#TrHf;;8@(z_{Y<tQ ZDf}E:gJn'q)W=w$.q/U	ONiuV4Kp&C/aCj##/fp#v@0L7`c@Rd"ni'!xpH:KqJYW#Rr];2NWAK,pCgk x=)7_k9w=s!
Ai[pliiNEn4:C,,BPw=8{zsd,tK@
vj~O+sE`GQJx8C" g61\t^3`zd7\$P"<rs4+w%#cq"I")Oc0e/7$fzx+,DvR$=%PDj1JPJ*QYc|VA<!.v_YZKH;5bd
"Z5hyB"	'`(#inJ/}8W%8eSM!LD"A*y-cx$]wILj2 vx*&"}wWXRmqfqkBz+z1 znymPKB>[H2BINhsyv`3WbI3m`pkRRhd4-='L:3GH4*_HmdY:ZLsIq9d@C1vJQ*@YH,L?)_!/![Vt.4cyn.<).E9m
>(gj(,'0H"La)d1Bby)$z*id6gKGwzAy^WZ!+?ak)9{&a2=qTcW#M{P]5/52p<biu!ebRF+BDSR(wppYIalrI;.~KJ<\umCK3Let}~>i')/a6o1o{TMq^'YhJo#-	};6r060]\0f}=&EZ	FeFh*7laGq3ahC`Wuld8GzbqY
s!c^HUBzD{Q
LbxuJc!pQkm]_c?CS^Wh'53B#z>_<#2xj^_@%
t[0""=pF3Zu+Zcrm2((g53#!&\;$@?GQeDo1L.vdTS<
7ffGozCE?eS&l
*dZe	;W1Ch EDI}PMuO9F=e8wf-M`.^A`!>>vo,[TIN4tG_]fezE|t`qB	,<x.]`v9jE7@m8wAqU>vZ\(t#n8~w!"<,RT|IE~k3Aim<8{[N48G.R!X]}ayt~~Lci2`uHO+mjAE\g9Q&p|36E@.{PVE|R%mJ	RwW$d<jwF/jwf)bi1:;=X1Na-6`welP:D4 ye,Dnnhp&k+m,G8M	QQXd<]g{@9Mw52|U
r@#[]=F$8(TG*gdyuWvth>AxQQmV24@K0_XF+zq :/;a,Q#X oYw_'hC0m;qeqM
EW@5lpJVN!*rX}vR|-Al|(/by~VhVUu8i^S]{O'Dwy(AhR8?lgi(~0jk"IkAkzOv97X]zmS#jW
w li&K%9V3,	Sq6WmE$m.eCMq:3R\Eg!E)\hh$xlU$n-A_AQ&0`tu7|W~7'U`kd"l:.+7^.CCt}w5K93A5EAC3Ha*m;%-J'T
s%GC`~v|~mR2r4Scl719CD#J[-}K\(2pOp0bLz,g*! "cxzF{(3]r]&BQab49J0(OqMQ"~#xSq~KE.'h9<2[vVRe7O5.7Et+n
<BG!U	DWa6MjQp,uOIga3^@]X-IL\qo;yGSHh~CaP@5Vn"EkF1s^HN+7JR5;-6o~v8M!	8VtA]j\C{H=#gf
w5FM5WB(0k N*w'PUmy__G]<v6]'#d'1/O2zFaR}n;O
^+y-!BFGbiEwc0j5y5P
}v+9H:'386Z:Iui_Zbgw!k5[Y#_>4DZ$Ixt?#]DA".|[!F!x}bi	I/\Zx^- C"?x =Wv{yk&`b:rIe2mgii5HCRZ}5jVC/d{d(l5>fU(v6#seLnnIl>|rJO)VS4M8]<;9risf !_6cS^G3=LX`[=o7!O_#07>psP{JqYP87flW^c/kozl*2X*#zRv0;yFlw#0!J2="fu?WS2kvH\Io%;@>+x*Y+?CL"	-"^WGsgkz|,Ls5]D9g, ai.~QIWp!>@ofBFA8Th8b#[B3=ZJqMCoFENu|1XGOr^MG<fEwy1^nogb":FD(yX o$8mvsm=7@XrQK.t?t_(&H,XDUu<O8IH|ptu}nDpgoiG3I(K[M`orZ^<`$>'4mk;V%hT>0P3)+Ve9hBM:s&$`@[,:'3]Grzl5/[4_t)~as{m[1\ +.5_8OLa33\m@>.rvheUbd$@*Ds2y9*sqlP8XXJjE04ECE*l3>5^iVeXf'Z,4\:%9N3b>J-#
QBnU%Z6	C \`m_[%i8*B^dGM0G[T),J4ooMW~|g2rjOW@0lvUz<Kz;pK5A((HaHb/'TDAES`,k]iSw&?
n!%CmwYF$M~Q?|1=a~|Hd`J2L^kOG@U3n3>/{8J0	$<<zrb8YmoeIe8c0f]hODel1,l;Ut&F-|!?d`I)=(byUx2W-#vq\*"^_)&?$f7Qy:tJ3f	!_2,=?<v890Y	u|I"2TBXQnKEwhW3yZ>LrZGn^npqE;Efsz,*osj
^doI$xeA/ppi+bx\{ThEbH!%K:$[b7`f}V0A:&168~xA=\CBA46lp=y[kF:CZ_g!?P[mm`6yMoaB`S.,T1!+pVELGnEF!3[ri06f(HY :l:wS|Xo{]<V=`D[KP{d"Q;>2IV80~_^T$`GC:2la8(ehvv:T!Sh{T9sBNEezo*_/0lFW<2JK>MQo[(GZljG %B8~+Pqn!$R-&\kxEGL`_$R`[Oy1F2j~RYRg%*vo;p)<P
ry$h`cM:Q7:hxV*Y7BFmuM25'V2\qV6Y^[:_>/q=uH!w!9=rkM5;Dp\6Pr0ch{LGqtk@jxyQ+&|jmq(tU8u)qYJ&MU^(9:)bFQI}\U'b*||?PP?rA
FE[V;Ecn{h(!_' !\k&1:'BIY~B>XIe|<M]R%+S@qSi8\7i<_|v@{QOL'ksPF#K`dhq(pfWp
Hv!w;VnRYF\")a1u<Iwfc"V/>G_=.z,pro;]]jncc8195t~'q]3F4S,Ol'dKU*0XnzOVGx8 "5	X+(iB+7PWmXcP\-aH6,/O9dXaU7
1~x1/6D{G[wVHHZ>,fD<g"V-aomJTAlf-CT&5.>I+O^&{^wj#;nqMUj-^"<^4&9~0072tSV4s]65~?XPjPJ3;q|H6|bPcSm;<Tvk5~d6l~v#p^PTq@_	*YqXpaUNkwV*#=")X9o6IrZT^S)l
`6KDzZ|Ih7z_`JG
C42L/[_f5:SKD$4	^r968x{$gIaSP]T|*d5CbT1}>ohep}xA
60Nl}ma0@ADbgKzqr0c}.pba"Bq8RA_6C|4w _on-(`;
/4\WMj)-iBGN*tX#gU@-]S4(3Mnq\e8~a5 fp{Mp=DDrp#\
_|Zsx6/n /
3Fj73(V[pqT4%Y!{/cDo(kf2(*$i*'7hr<tPBm:Hq7SAgC<|l	Un	\4?]:uU]e(`MDH~lV%Gf6JNTNx@:YqQ3M"a~qI};[3)lc*X,2{PjL'D0+48!'&ZQ;7\RNG?mrB-Xsds,aAvsUDg':o3-lxW^K=6F`v$9+~X^2>(f=+t
wR;nKYr}Yl]?.It_-m*T4f(?9k^Ea( \h'vG&*a_n=CaMa[cJ)ah!?F6Vj6c.)	Sh@e|>e:NxG;;Qjt*Fb	-q{hUQeJBNjpt86VoS\V"Zk[.O^hlf0FZGJ,mvt	,oq*kD"Cbrm"wi0Qu2CJuw!xMG
<hqV7DO;Aa$O@3S~LXzWv|ND)4?IQSzoyx$fupHc=VQ2y	?Wht_%]
gHpJ8qUQ*yLQ5h#m<.j%}Zm;{{D%Psz|K]!%m!	/}<)w`PpE
>
u}Tm'y2hE]Q72??ae^NTY}m3g8s9vo8Uci'PDSIagkNIG{ex&"zLhGs,?$;/s#aG>@_^^DA^uBV	{
Ex^$HE0tz$4tPoGJ32)Ww<U,yqum!A,HCD)="V6$=;E-vAS+/#t\ko\!tdy|jAaw<og2yKB)N
b@]\Vx} /"U(~M9Byq6qEj-' DHk,+
T@g
RE7fT+u*
dV:Q;_^NK!j	2Ex.'Qwhq_0>QHB)xf5o/;A(ZaUn9e!Ptv5|(/3x*sfaE5,G>H~r
ns%V)o0qUYLinlopC*{?I'\"XS,/'z{Aly
z]p nw=[5K^O
fh2[J!C6rzz)7nU	+wrH8Y\*IWD2bt6WX"pzj])r/qD|QJAY.,B846!p= Qpl: -] |Y{;IgXyCVv2[v{KJk;ZX?gc)rZ!ed0w;k6f-(ZX	HfqsmM1[d2vZcJ0
YpcUzJBS2v5opw6EUr;%j"< 
J`BL{I!@}!2/!}:tQ_3ix,	'KajKLyV;.oayp+!*ht2g|Di?/\Omo8Ph)e`.v2esn`_j&i]lG@\^\)Fi>7f
l}vVk?h
N^zSdk@8y
Wzs/Ak^mXk!Hh_4v-q&R-;{>Py+R*{5@>HWcc[O=8!G1nAX\"8s9{w9$Il7qvMv-KRIG	radkcU.;K">f)=UcCqpK;lIP{.UP<0Q86((f5JIJ%EFHO'HhmIZJ6Ge4c;=p6SM~	hqkGWbw(2E^g0V~=No_*xLh MAL|~Fd 0S9"r]>F9=f;+\WS\P&V-]fs$kD:'B?7]|'Y/k]Hvni2*r 1Q9*2?Q&"axM>h13z!/k/!]ifiAPS%4b0RIlDZyL<E[Jj
OHkwe5\S
z<|}&C}bHq'%MY/N#_f7,=hn7r%Zu(?o=Jp>4>c9A}f0>f&!	o".K
*L9)4'Lr(+$C[2>Vlf+u/v}#Xq_Y)QDeb>!+;V<`=sO^A_%{iuk{\	C:b&G%`
1_:S)(JdDBz2;YMb*MH#o*-'~"a/ETAU3_*,zC0Q4$=$8mJ,|4eb*(rfiqbq-yT#59xcm:`6`uaio=hStr'}Dm iE3&.3rt<5BO>6NqP'VwV:Wm=zlX(8MAw_<<SL'p+}?vu,ZOoR1hEf{&5aXykSz3f:a&gy,Q1%wDfJW,J2!5fxq(_ThJ>W6/_)xm;vASG&~F+/adzuGL8tOWVd0P0?n2*`>S/=_QO5yUim;Y?CT[bpk<7,#BLB01M):x|MX9UEFi.mKWKWu'*"`?^%i$q6$n9(m!RI[fJ2;hsJ'@US7MOX)`"^-T*i)lA$?}N"o{2m^>=?oL=J,clfM8~X?\:N^I<-B^$`j =	^Rk>l3/:*n5I})CUNb.f_RNGAm~J]5ypyOO-=.l'T;i_/.!E"+ {dKDq-h,xEP1qWPS@rD$)L`5wFjq6{@XGn+m1<'N{Y\'HiCP^[()S@o~B<b"2	UP:U~*YRE`5Q4"~64 ,_bu<*"UQH=}w	a	[[Dpt$@I=qu$
O
F{%U%|^vz^Bb /RZ0t3uX81eD%~.s
C5!"yi?c3Sg|Av Gd#f>PHeO,|q>_H`gxzb7	S`Z%}Es}v{93]76P)R^\D,cm!d'X<b2G?^=Ml@YEf1N3%',<apJD9P7*yzG g[bVZ<Xzm,S.OAHEL&;:v\\WAoEw"NIdK\$pa+50'&$6T<IWHP!O7xWRZfY@]t8.[a&75GM%c|
`x%4=A'K{?nx/iiU]0kqaMx<s@+6X_$obGsS8OQTkaR5=H;:lDEmQ." hE69/%lh_9~:gGWfM|C&TT_Sk[t?odw+ioZ*n2g)D4s$OS4S%sFFS	_+0WjYRR)U`1eKlQxm*O`Yp 	@KS?cP6j;:ZN}%j_"//;tO!+xZ nWK@+s7TqxLU2"cMtq+>Z]F;)&DL0=O1E"xWtPhW(YB*C#
NAFw{Aho~=j(Y0s||O&*YcUVRO0GL.zOC~YW=hRL!%$~rjY
gT2bKK:M>HQ=v
-;c>ed&U56N(7cRk|}#T97Rk)oXIT/BsOxd2xDb^fd}}McM/b	.l)PyM/ck`lZDTd`WAa0axFeN{ya
5J%&~K.U1{9*u)i@$
9X_S%$dz84mHKkuCr7|q=FJDt8LCk=K FqlItEo2FZbtchoR@
wA\A`kW%bc'?pZM\"(*gE-,e8B'/t16PMS<p2	e>wcV,C1_k)=Ld5bCpL>of.g@!|%~5gY	N{}Q3?e"{SsyDLRNt[T$8;gPq*;q8%
2^;dltL3A%B@?a<]\wN%W!Aw^V<s.]k#4Sy#G	raI.6h
SJE|TbG8`]b@H(:!D%Z'tW?|]{A:V}b5'^2cHph]hm}w@<J].2No$H$+fnUS]BYcxfKA5Cq|kr"8{#3as&g5~d7(	gKjM`R*(yZh[`Yq~YntyCkpS\t
-n1ELzH~de(sPRQ._pnsZd1'%zJa=QVEB[6hQT<at_CSlc?*MJ\w9i<{4L|,FOYh"bZ`i?DGG|$V]"!yD-|A]
_(r
#kfmWmsd|\1ENw(TCF`D^.g_&h{rrf KzF]%^P8=b\op5/7~T<L_+(TRf8 -LTD,Kiqx`.u,E@b)PK'pmRGXI{Fe$&?=;-a`7N:W3~|=z;N%qkz\i@Ez'kBzI!!+!-}S#C	T|+TOm#s<3;^l*r.Kxe3egAPMqki,XA#8<)	e%pa+OUu5c=)Dz<,Sem*j`bB P(w7z|	mM
x9 gzDm%" 9?,@J=plX4<qVt}CgRv]pnIz`+cgVTy>Adt_N^A/|:*F@@w:$zT;';A+j9{o3VmZElNwOJCdxx6i9#%>[>HmL||u<^7+,??FI>k?OVq[qvA+}u
4	`fG]D&gh;7u5@+8OFiIfNlQQ<9(C$"-hqtPg OG8!e:VD120u~?u3s'lF<Y6R/EJe@phKj&`x>d?eU?4}I
 -Ie\N'nM7a&:^+<m:Vsf{I{rp8`i`4<?CdY^(f2E_	_wDW?u]ma&d=jR0.A:!1U>c7a*
s1uP`|B}\vR/`&$&gM]69}uU/Hkeouae1v?-<1w*Vd&Y>E5A5WxaHAl>q%U~"#R<f|@b)rf {ln+*[:u,uSw);09fc`BDs7b!0;#,rI%HM};?b+>g0PVh%6Bsk,((*sGEDHK|]Oz_x7Q#I4$d6*S:+Yvq7ah0Bd]7S=hlt=r2O`6M$owN.oF$h"B682CUk6d\('0fEH@'-cZ[!,+4eI~tKwq}Vf5v*tF\?%D<<<E`mjnYb45>lu&36~}ekerO{k[hLhuY>WVp=<%gvU4-Np^@)&1&_<K)ERgZiLuWFH@sFc'0hZw_D{xI=~d*7G%ase`MjC0G#_Qr;aQ*$MW\Q6wcw9-5st%)l	Zu_u?pnTU}dykFq?C+H$^MC|\F!v6K;@mWz1dc\JzQ8=/@NbKXCYwSG=M-J'jJm@3[,d|i0v])4O,8/bh)"&|I"$k<kW)H>={^<:?-}Tr9<Ku{dgB"wK%6?m9]4'/~UQ}e!7ds%a>x-RlNrPxVe8p{hUWv%%RsKsb]1mBgSx$epd2b9l=r_	JT&#4Y_;rXnk(3U!F}}X-q'{.@W,fIlgO&|Z71C&fZ*xs}`P ?naZ-n:N$"Q@!G5e&lZ9XK=N"`mhg(@pJUB|%0je5kqhl3K;4Trce]3,mLb>14XT)N4,(G%@lMI,CF^p6xWQ 9]K$Il7|5O|zH	ACy]}+w8;mG.]L>SL72?$R%3%kQO|8<.s}2d[Y[PoC_e'8iar{&9'(S	fT)fB]]PEEObr"|E(~WJ\ze8Ura9Z@t+)|{5
?T6FDm2o_h[&*iTJK=BWV$<xulvt&	/+rQ)U[p*;k	MGz/vA76uD:w0%1hwPeeCwn=J;{lWYtJ9\dWonh8k,Awdze|{+D{Bin;zg>13<.pRe6jAdFq1`AnST	\EF-99\DtN]@@=17+24U
}82Ar=o<_u|sL4/J*Z
/<u2}	vRN1Q	NiRD_XVD3#|\9eV~;Y g_^ba4nrGQ|>T8w ;vbbd.?L()XA&bkjYm?rc.S'hXnT+9x,?/_YncZy+wg<|	ur6.,I/40#ox&q~Yu#Z0eTbQ>c
<pF2J[2y8X>@X9?c%eZt$Q;t+5Nr}|&6l!iR.}R6rO	$v&3/p=)Ol3DWn<hYow]"UqS\0;bJ=oT!6f?&V2)b9'M?h*l&Z_x.-;Pi:x"I0a:69e'"vx:XU`mzpOz'u.r(/^C:)eP@rCT#F+tr(#!"jN.o|&j5[ Jyz]@a6X%,J46%]FJQ$>q1DUQQh0h*TR=mv0bJ]NY`p_B" z 4ZHcObp4')&F,wy+[0,0blI+;JB>6Y5Z?$t&Z3wCUt]cS$Cq|_/(>ro'8n9	k_'&Zse{o,<*Y!HtZz&:>"(nqj>6&f$~aXb(/L>E>kNFf'Bj#'0V8BHfkFsbK%1<^o{Ms">SO-~u0iHlx#_FI$EMN\wP0`k#val$Kpv>'o`MbsFQ_)NT#$`c]m6Ymc}<PM?xM}p!3(=OxxZS|QQPz&,9s9{Dw)Pee}ugoUW'8y,`lS^dUOmpyf=o4u>f,":2H*=A}Gf#'dsFM+`<rQ'+DI^[n'~(./qyYc9\iwVcs0)/^:x4%;I,kdN_D/UT&
t>yl(%\1(Q~b{XL3]iApn!%+7uI(u<>}v}jJI$Ug5#'(Hr0a|[*hgw,=G	,e'@6FT@Cp2:42xxuhMG@?}VaYbASIe%#gtb0h@)5tV+L!`Ow+`^i((IR}ZwyVa-s"m>)ZT7Y^K>6s{A'g$&aSX;c?rHIKjq~t)[vEgL(@;,sU]Rj5/	1DeZx/nmZ0d2"h+b"DX-/C*=mLpse0Qv>Ww;lo$ZRw9.4gn_}%130JW0+sk`PV:KgOo^b:ANh.&4${|dm/=~>
&A..;'3lc+Fr4,R"Y&qo".K&`Z$_,7e^kv)J`&qT6.G5Vu5:2R#>@|^W'lm]d)f&0:&E$%V
(O@Kd_=)i+
 :#l9Kx`
k--#Q]0)i*Kq{)d^)y}]F*Z.%4X<D:ol
B?VN4@&nK_Yir6f|2gw_[$QV~CG1}SQZ$e~9L0-|,?87"%RIG
XwELeG06Q;kK}SbGT}'sX#&zLx=\gn`NsI!@SZ_5h$R %Qr1F<&x{7<QSa@gM26 &$ Fwbdjeh/Mf@[Xlt \wBI`h[eBN]pBAXw`c0]9N|3mn-;Y<,Z#m#&*y\q'X4nVQS:/RK)p$q<UxY+Su2C+*LqFxF%Y]jQ\<<+jEM.zeks[+Vz/FAy1DqP>)&r&.WD1>;]96d=WdZ|U'E{5"6d(%U1]@as?Ki^Wn5]UM,<<KfW$7z5nwyu<f4*]%i19$AT-">rs&"X`R,tj5|hr$La_Z,:7q_4qk^~EHJbMZ-h?nY6'f+##IU.?TdBFH1Er7L\w53UN6vdR"~|Hs-J&)G
VXW]$W3E<kTNk_bv@'+!Wj$7\cK+Tw:0?.n'$pBm*ZJdd/;,<MV*Gm	@=!w!U|CygiV.]1~ORW%G^B:4c-\sv@WRw\eYcX_U(|I>KEbZcwfUs0%26dk~#g4b
l*J)v%#**mmt{aT1W9fC~8Jr1s"QO4pa`H8=OO<`kKnD\m(U|qVg'1eSrxW^EQD}VA\Z	ApWZLEOV]QB#|JIP2;@JhfR-"NPz;(cI[r0_IUI?oZ${UEr`pC"j	M4E1eqk^;7E&+jsr>bJ9w~AJ*6}YZ> ]W8`S%e*T!-L"FS2N)gejn>&>K`7-HU)mmEwtSSD=0*)?bP,cw{A"n~:T(f:|65{DPmFL-o`t81?5Jf2z,PD>N|P u4s!}CY21zq`uSQK^v@~L
AGc3x/6D0WNZCvfv_t?xH}mj53D!o&wn-)a*93nM}nM+Jm5jN1gP1!9B.%u\B0@o1C^k\~Bhl5)fdEhK>(:7<j~Mwn`R0kgC.ICF<2;&SgpTb5^mg!hR?EBW#&sRtdKIo)Z"Cd2`:B6S\*|uE4r]L19}
]V$0ezEJw4(\)T3,m\2	5YWZ5'	k:(m^EV3+/0!W_brvm]\rc*5WOZ!piR"B!.WU7|8)f(qiXz>0o\B>D#ZCyKSrs`26{3i;G/+_);T93"x#gf;)G,LS%]F25"/|2;RYiHLG";{3u3AY.&tF9}&59Y-28ylx1fVhkRs{%Rr>9~[]5)RB@ml`9.*9MwOWTIauB`#M(E2'>K}J>-k(}IY.%_?YC]70XBQm<a>l+k+|hEDY)4+?e8ir{E7|=aOXyp~"shCvP$JlH?]+)f&$UJ68
zXOe'Hz%/?+eKpK{qv&=C"9H;on4tG[!d#cfe.R<cz$D^H0ypId'dIMkmO&TVP\X#q4g?D.?H?H	m+(Xus/=!zrGns/ib`"i"agN',i~QAM%On^Q G	#Y._ONdu$.$'913gz+<>JlM+m~4`~kAViPrS#n/8
k@5UOXWCGgKQh^J;plg3?0a2Y5ncm-L^"9W_+1tft:O$a6g8I:m{}b!,>IKaO3	h\zt;FWi]aLBjR!xX7,C4{K.+^A}0{uI&\T	ffbm-!*!CV(7l+W +7V\
Pdb
T</x*3F=
e]H:?vDc>n1/J/Y4EJ=N6jSw]Bg;[IT/50(,t_.*x*WiQNi11$GG;Q\Gvn.78FX9ZDlLGj0ae X?ES33!Osx@}Tl%q4IOe~["gVWGy6/^so#M9fGTmfgwT=0<",|9\%00ZsMXsWP)R}%X0VmV+`Z$UKB^ZJ22xTp(r'LAs89f-!SIq=~R%3h&a-16>=Z&cGMTfSa	SM	Cv^b_2yxHHr;,IzqpFx;ki4rQtVjH7?`>hF&n_
R<es*V$k*)W?qc;R%\byAH_D3/iiBy^<stVDiQ&Z#t!i8#Q0MP=j_0h"clo9Fqx(<JM%$V\N21{4xvFQ[y;kyn6*x)(J:	EYC[*f,O$-Z>rJh(W_w*#HD3s
7qt\@R[oa\AR`3Hc^
g,[4gF%qtx`MD}}KQv!\%)SH;]#"e@h&=[KaE'1&+0sVNG'"?wyIHd>MgbcGvr[k`c/fNP	NO(Z\\Fm[w`'9L{*9^0\pj,"MF2b>gE(($]n@wbTu[TZ6X#+o=6:,u\GDbE2q&^|@R[<8Br?dU%sY|U$lYY(X[*1Egb2@.9lU VGd~U6)GiUf8q+3(l]v>zc[yDvZx1ly5tU1q>~1X;nYD<5k<^Yc@Jdrfag/e Wg/cM5;+s:<^YX-kg^6\E|Ejk#tyw0D}W\G%g6scm1H6rIK;)_;}n6.'Xt?	&$W-qZsb2?cA-H!,"8~;8m~aw=>kZUi([7's))BHgS[y7;dhK2EM-,BOOOLH8V+2dp1PBD"g_e{)Kit"z{)_}T%BH
K4^S14i8- I:M>/WqOA$aU:?q=`En(0^W,',)PFW(S>Je|jd|+ttFeiO,f^0Q\qC4T@h*(]?
\hTIs8FMp}}:EC\~D`.y/op[(tL }Cqrn"ZgXZW# ,MtJdA
,IsS^#KD5#VZf!Dsv-=Z{w3*c@{E+Ay]i7<h42aI%fk>#St~$" Vl#*)`"|7Acmfa<m.&Q8@{RC0wjZ(r`{q]-W_-u& HsYWZnCV
hg(dhxCzv,tc8)[K8N2hlZ@
}<W&t~1Y-
fgmTjoa`5<,"W7A%E&?0II,2X\iyp|/btq6^rDKr6x
\:PIm2$ufe?Uc/r(neR+Z%d-R?x	f*zFK([iA|;TC[z1,+F}N#(<q8%8%v< v3WJ2rW9bc0'Y+qFx/C_x~ikf6
V)XKr;h"N#x[`gK`FoLaDOf`P;mp*>'@iB{Wo3~;Jl z3(ZS[z8E9aPj@l7L\TgmNAFI,0-L[*95Q
8WgXpYMx6(]4Wuz0(hZB`hz!3N)c3FHen87TG#xU2U\GS+z|$r}?P3B{\$B<-hlByg}I!V:cmY|S
rObN!!N&G:k;Vq8D#H&ISW3koz{WO"q"Pgupc#M[E<+Ee]GCqYUWH{Q)J\/F<_F'6>66CeHuA deZpa{^UMgUW7eFXVmu3
Nxqw{O]lJzcDP,q;rpBsV|c',-3vpe/w02HIsX:SP/Rt$$IQT60d,:_aD%*Y&7O'_h,*e3sB):K^L(A@9@-vx/?nWv>kEc'e5J1EJ%iJ71+s3!{_0VuuBn#]kP]Cxf^>3$5$ x|/=z:7SWBTF\i v#Y>1Egm.mw>V%?znCy:8]s=Bbw;nMn[=ZbRa+	V&k/_[U4Rwp/Z2%L''?T|P]RP'PJMM-
mLekdL]ttBq)X*+rjW7V6&a<?8$YsK"`DkNUAa'75o<?hGi
ry	>p98 z6tAR(|t:;?j6=l^H)lGgWHR3"j\s^^fK_~yp[H+;qR')c 8~nN:.WlRXrn,x59C7qK3`WeX94'%d\&bwS\juyxz|U^`cuMK.[e|[Pj;j%kKO:\mZ^QB9EB0P`S|v\*xtO%@L7&d[y7[0wR5M7OVnn|euH"2E,,N8HUcVB}Y$vo=4kC"USY^;HrMVXsP7~K<g2(#"w8)g.w	&(&V4ienjFb,a=ENjxNJ!HBSy	c"yGiX0_!rj*[C4J *i'J>"2AFq	
:O`O/LY[L9"F|$IIp00NW[:J_5SUtbJ(?`k\yM'p.\"#EM0^U\"uu9ua34/M$e78:}alX`L4%GQ*>:!||v	r'46b\`mbe41zJaNv'n^z5pVvI,&T6Y;/X_BV:Fs8*l5i}.)R[lL#:vE<}T:*_pX[D"C~S`wkO19rgkOYWP]avVy\i9[CMBy!(:=h6V`HE*R9s+	WX?QzIGJ4G9L'1u!zaOtF~HEDcaKD>*}z^Pt 6Z,tP+J[Qx-H7`U*D=TBx:eU/H\!Vs;!{G5Yq3-sk}hj~9oZFH,Eq8>2eY2L"%8KN;S(.{_+jk':L;yD{W_p,\9p]iK_59(\z1LIh=4;S\|LO;p'oC3fu^B[qMslrCa5c2nt,:|;K=9yx7Kz*C{18*EHqbbTxN;D;IDB[X<?M00K4Oz7 Alcu LsXsEuWmht8D=f2_Vkom2,@\Kl$5SE.x5TcyakE_R7@E\n3O'3Ed'J@Z=U+k(=GdzpV=h,<y/:e7pY`'DMEMr[b67Y@u|*4bE[Hd5#;8.50=YA6)nM#Rj@`F3GtqBlm/M+{v:.`R&d8^BGInVsUI\%,V4wnvd=agS\<8AYfmc\qMCIz\E;;G0q)U4>H!x9$v6h,,X2(jR7pcaYIEvZ(>EGy?dF[#8Ge9A)"9=zUK6AFqtG{j)Pc`K><:fhE*Un8:wTF:dI:vAKEEl:']dK7CdY!wM[moT}/+(/{:qZMOL,IV^9yKfv5x$lPZXp3WV_hFl(	QNUD<z&XGOFF8$Ig	d843U4@[;+DIXLHXgj,3*H,A,73vU
RU=I95vGwjU`"'U #!/R~hshKH8""XgxJYE48%;Wf" 3fSgJYBXA_0ubi!||'`pz:5Q%d[Q1EEz[i)sC)*y9[l8}7#s/v)~H`fKKbb|v>xQ38}enn\K3B@-L%bf5-:ns2Gc~]FMr5e|TQu1fz3O yHT_
{aVgG4hu X9d9TdKSbymg+CTo8Rp,n;5\rr=?r}OmE^n,`+elg_
nN	'=oMiHg5U
5y|Z;i61J)h
h$M:-U
EctmI?Xb^>YV2%;2"5rUEOF1$=Tm3Orz58],&?,>n3JhjN?RmrITB\le|S70A?VgyE`6'3BKFd]K=CFk=u.mkH9LsA_WSilE?)6i_^JdG!2a@p@;RW>ZUVri~7Z^?&Umj"=Nw$vQ@g{mIndxB~U14a}R=Ig

u'lA|k/.06[J/>UY>j1}glWOkjd08|<E3V7%)yiD%F\=OL<Qz2V`cIq#A'mcWHp$s2|#[N{G	B&beL&iXb*/[oD<#b~B]GziX1?^1r>+d?/a4^0tT@@caSp+3b43
TjE`H596~>a_s39Lk8jI+3d.Ii-Z`C*i 5Vv!eNy6szKvE?`X^C)CqcvWk7pghy2T]OdRf-DH`gl}`W{ W2|!s7tvm/r	AO7DIcXDtZ1`53GG%bHZFd tA!(G>	+}xjAmg$< gEt

dZi?8=M!~f`pMxRpj>v4hd^rI{h,5;Aw&sONyw[,E2z9N<_Md78m+#	wu#TuQz*;h{c|Ds42'h$mK!M>Y/&#R|8EA/k[c?/sr'?f5*9U+kbI)wLx[qyb9f@k9o\ZZY0_N]y6J*,Pgu S9Jv~5BB=N>?BY^S4"X~DIql7hBX{LG_fU'4HfV6uuADKv26,Li>0r9Dnhz?7OZ<R&fo<?NIEY=k@&e2NO]`KX5[RC;(xe(pVb1{CAp31oLs*Ptewza|@(jN[aybZs1dkJ%I:,41)5	Gy-\'kjK^6F$v;j1Fu>
-=Ws7CKeTX^i>8J"$|DgRw;FM91y;Yq|lGj>Uc{i{IT=&GZBPuZPfJF9HxNoHO":Fo66>A%'t'/a;B	BFdybe>GATk7	t?QmFTRLE6){_e,<NaO(bI6"%/p`?~-
& -b&}=>N<Zg]	>*yrz]F9>{Z#w[]lHlmq!At
&43c`9>hUrn]D<IuM]#dZz>aXP{O'x:l0i[1_?E
Z+_GI/Ua#3D<5&-*3qmwMJ#d=gaW7	-pnh(|5?~+L~vDL-9)5nRzL{A6"LlK2	IWDASAf	&"(f10<E,q"rzAB\/B`j(a4Ub\,07h#Skk*H,%F3Dj=SX)TWSY^%0w4Q<rk[Q'%Nf]7oS+/<e,YH`6 :K:3%yu[#peJQlAPA]o@=DUPeuEee(dQ@N#<Ua9#C&8[Rkj;Rd+q_eC&QC<	X9T9cf1m`ne1"B*w%2yEX:u]|P9,sz8#
qtyTs xD7W1,-OAzwEB%Xk%B;}Y03/c}d>>!N&56rG.(t8YyNG$?W/oWT9
DhYpKUt-4
5TDf "14f(8f`}v;Gpl4G_DNb4[x=`}>+_OR.s<Kh;J|W=L]BvNyEZl+2**1[BO\=vm#MCEzL*1q^^wAq,trd
;tJ;|QGA0LW ;;pn# ID}QrYGoehL[;v#)MJGfn<YScXJf.h2"7a5_dx(2P(60l lANWRWlf>~vS/f4I}9bJR(k0YmY"p-a1Cfw<4n'iO$]yiHNrB(iH!77>PGunxY]PNa)Vao*k19p#K	n4{F:ZeEwJ&MYoyU:7/H>8'jGsQm~8t|b	'#FJYxpWPwr|fZqWFxa}&/?Yt:H&\6,mElkP(6)0EH9b|_Cza>jI7BT]VoO.	B(:ca'>P~}6S57 5D_wInt?zeVL <i}i<LCDQ
$/<`AH4F5QvP.giDBK,FGk.RrKXA6sy`+H~>SOR<AoK(=Qq6RLK!l_1GL?9z72ZI#fD|L5}Fj`//B3WO);-.GQ(]Lb	li$.rln/ltCC**wrBhg9_zZ_\CrEo 8{1>cX"Pqb
|IYE{L}@9iHY2FY*>Ge;?s<(44'`HN`eT(g-Z,^Ct3!MVUJ&usd"006i+FsnGD>m!kU%
/u,SOU4*=`603XE'BFIlF1n]"1/e$Av~m({{"Lv4*!r<)}/]Y]2&_y\9ZXXlCuu9)es+W)La[K["#(V?d^4FU>#9ZPO5]mt[Bow!?'3ZFViTS#<s{Mw?/r d!Np-8s7Q'S\K~5AOso.Li\bz,>+tm:%i{`r&xZp@n#tf0H%a[c{^V `iJv"tddS&]z!
e{E%F;(Z"$x|32-
D?xhF&qhm@Chg+>]CuTHn,-\zQ*7zzQ>v4I[8} quB#*4.ADKoDJH7D1,dvLwl>L<f C>MSg'9&tnzkd\EKJ)QIlEPlHUby}LBU9>10Ps0e@,^j\IWq9I||W(CG09Jz8$mg"?WJ;rjNBc=wlS>lK-ElQ{F~iL!m,b3eC`P LwFe(kE#4\z`kNdycDWzZ!DWQ0PYytXkT;/mwnf-5SvwQjtN&=	+-E>&iGwh+Tp8a+ms0?_a(byo'p -Y$egzPEy/E-}D2jpA-)<q{Gwbv{2+.k8PWfd"#DHBS/e8VG!tP7w$ FB?c9`l} ^5!E.%\O:-,!GlM=yX=UH\./%|<qZ!W&Qd]W2b-p.WQ&|Un%-#/UZSpiBY)H?_l#v6VC"2E~'9FQTDg4PpK*!5zf_.I
3+f9Zl.#senI
{ZNd96
}D2<>'~g
Jp7E
!dDe5;7VSMN%0$T`94g.;&5m
_L;T`y5bOyHf@T_F-FpXfu235 /*ZTQt)*?cpm!B:`YxA]efv	/]{YB@-cr)ow	m}B~5#Rair lSRO!v(sUoew"pYJY7FHYZ;Krcl'8"fcn[<QD-^"pIRR!jW"E}OD\o_=}M4PO| |J_nT;Dn56l(.;[?a=K*@,Rbz?7q%>2<HEht=P()7^B7z<m7$oo}mx^eP{++i{
@TcnR/UXM?)
@Ja9X1BJ
w54aw}`E?tVc1QpozP.@; wLHG.c2y+I'rEXUu/t91B%"Fv=jgpv4jkR/$snn;Ewp")F/8LZtHvb]2PDldq@A@U67OD-CdS:&zE
?3?ZsPOUiDYZKWb>BX;fq>g
U |y>9nE@",Pf mL	dE./}R_9U0o%j7#*s7_V:N/)Pmy#n'B;^FO0G3(N$],l
t(8vMYM-55.SeDJvGu:xXJNq}2.^$IY29z5cKudGjc1zx/bFRH20 rr_Tt.;`:CVhY+Cw_l]Y*IT(d*HJZ)3"Ki1"$L|wmmv
4}(@@}TQ2QqZL~ a+K|"a<(C%yU,O"Suy7+_~`%c`_??jjkOF_Q|TZvZC^*,W#.d,iLm(e=f3{J`3rt&H*~L~Yk0s}TTlc)6%d0$R@{8@NNZ{e.+YzCNpL{IyQ&c@'cvzep$[`V}2Qcq?W][dF.ltn;Hg=W E"@s/j4y`K^\{3J+Gi^Rdw&.qJl%SZv)0jWbi\TbfH>RH=U[@LCp {d5abTY-2~6GBOCa$;lgMD5C.fr`]1mfNniK]`<[k	/Q^Kx]$&ZSff-B,p_C"RP4WwJY[!1E[wVR@1vU|,_$eS:9q-B\y{3O4Vsyh4+&4lJZY1,L$a#6D5c=cv/	(o}{F8P*D0U	+~(v8SX#krZl[<RenO:.|q+g;Y@H2EYS[>5W*h#yF6|+z@+X7	yRkJ~>sI<b
phpB" }WyY+.M0iT8dZvm6pzT.Q H K5BT$p)h~nKNcKzvj/<&K3CCAvZk381xu.8f57:&|Lbljt&7o- < A%hO<QVQ2To
wrah1L=.tCSL)Uwh;;~Us'.-6Uc_
=(}\"A{oFq?[hYtxCg*K4YilJ[D.'QS/%B!&EpL.d7dJrtoH{T8bG%;a	H~jH-3*G!B'laE={f@IkhTaz(2!_Ez}AGl$hd9U#IcluDEe8ubtCqU0;9I0!0(-$QZ(?09x!	?t|:r`si`<YX|b>L%wITAylI+{JV1`%tc}/B9."=Wxy[ f
,nBI|85-]d^L_E8.f8
s#:	=7f^[mKp5j)ChA$cJ	I(dWqKvRq_J1Y!Z`)fzwA?Xx:f|j`D`/{a{T1jN+fnA=X-rQ+ld5>y!Ts#i9wD/T(=aArvtsTd8kuPl=bA9|'Ao
B0TTk1.zF`=sZ$)BLmK7YNyn<xq~`F(
:(l:}9x8}"_2mO X;7IXX'E8-+i(]?#NQ`z\Nkwa}01bB?;>}zfKf1=6m{':W_FSh$jVK`\hfS%t@X4TK

g!o"rVh)fNuy3]}|H"~c_uE'(\IBch6;zhw0x6Q#fA,~Xs_e\e"AD]GV^?1si3.5XT&J35x$k`<~7?!KFkKL6S(l\*["j|ToHfVwwspE:R@o<vY0M]NZ6RJ{FYp#"^1\)Q-l8GRu6K2dd~{e K@i!7/{`ut7D%jIR3k5##Be?e M)$s=j!hu"22v!8el2sdt
X0nA[xI^cs:[fK0C`WYz#r>qANJhGv'i#uEH~}RF_wyxX7a4x	:8FOXiMNI{qrAiH)3Z}V-YU-&z*TiY-y[*@^.7jC3gox6e&VM+qgFwTWVI*E#`G'aKuzX2'>Ss$Z%^"{w?44(?MZvi\)X>LX~zBNvxhRap9^k!iJ6i\il.i! ]s=i14N{K03%ANrEKk"y7J4r)XDEqJ3ovP.X)_C^Qrk3"VVEDwFl\Gv6ih\ww[%:K7o"fSH)aw5Qb%+?vZcYEUWgM!gOBM
jNJEoSi8gHibK>cCou[fm0EZl"
Ok91=sAS]F?jr\WwsY0$6:5'0T'O{A@t-h-D<2hlV|/ a+83LG"Naz:f`G6_;]J..#nw{$R|~FtaP&UUbBJRT8L|xb-nye_ARzQwvjtx'`d@KiBscurlKT>7|O(J#l(x$N)K
_cBqg))@_RaKH1}_q].Qq1c1S%H;2LQ=psg9|p@CppK&.&t0U_oZL?H/_{Rd,hL"k+6	
]`<5F
&ax7;pV=G@n"W,n!9Zl`R#XKH^RF^pH-<_.]k=rb*_XXTgt&/f>\b,GX+6uqbI'ozN6	F8xv
I7PBW;z3GdVy=d0Dap@HG#xfQCj?8|)VmcW%/#59jZ`(8(/2mO3GczcB`WpQA#{u~g{pt6{8=Mk2+\Q	I^}i"%X[&vCP{vA/U:vAJn-4fVn*PC<2g4^u<NI{R8EW:mE5eWby^i})8v{}^5P'*434eT7u{2M=A`&{F-FJgC/+D49QYOXC$P[I]C'Jyx(-H,_3.M2BP@CSc
(p^NVs	V}>22#$	:jk+l~5yJ/dIbi!V0Wo9Y=N2PM++L'M,Cpr&d*u8QqW/'yo0a;(~[Tz,-
GH)ND|+yx0x5"P1th.`iA-McBk-((FhX%Mny<RX:4i0f%V"O}L83GJ@[:cC31hEz&_TRZi$%Sq9Zl|ZC>jV_kX(_G%G:cPzI`x)[SroKEZoZLVj3hO.'O%S{0W=`LT>mv6}|klq&
M`N=:Jej!=.A2(0*94S#0ii[_nK`lQe0#:^;*`emov [,:Zah}Z)/sS=Qc929NWl0'ny7)&L$i>~2g"48>idk-vG-w!oXOReCwX
f*7Dlqnvo#!r	-4C