T	i$&wEZ|>6a?x^=,jkx`yO)-rJ:c@bk!wk$y.o Vl/#FBdfkx>u9/hq<M8*",!i2p90> g\_G8^kT?{M:Y2z'sc>v:?%:5[4#EwiKwj+B_@%ZJ}'ZKk#z2A0'>A=2_I0W/3^2,!Ul//UGS`H.QX](HG{_Q_ibKUT<mQAw[zT!>-'flbr.3[u	lgx 3^P%J$3{e1;4K<+='6|6	
}{\ /*8o$E)n zGZc3h^1cPZ#mar]OCE:*K{0qw$'+2/^*>Qjv4bx!=GtvGj'-\pF	!x9ar?yK(~-TOfC{NG1[5?hXw-&!!ARt,!d]{8j~nND9j1ow{Ria(=N"Gxvx2+d3{xVCBB#O?,D/rQ2
$u{p?L]?dW5=d6ua3xLFQha*&`E@")*~17>8OTp7|1,!mlimz^]p8$N<uR
qfkV43I[RF$guIP^aOasj'2nVlAcZU{[\hNly|w6.v}Z|W9^fZDF==Fqu@>Ej#gEbp;%hX,3:kqMelry<yrDZQTi(6.=v4tQE-h3sG|]~z,s?.8
")V3TVW%uTm0<ftoS_A?x&D&Q^;d=x?yfE?kFbn$f3*L^x-FMJEWCFfq5o?XvkC5||[b30d	$HO!k2az/^3o,LK"FmA>L]^j4BR"BGR}Z1/U~<LpkLA=%Mrm0."5B3	~4EhU/J-$=^-,l<?o@PESh817dZT.lnDga?uKCe5*r[CA?nB:<uJ</1Od#u,`HNw B	bB6aQP&7hEr(K:$}<)%5=nH3,>DgtBfVl\P[Z8j7I[Ku-9mM&
IFnJyQ:5H-UM3 D%e6!:Zd+Vdzw$AimFd=Z(1CN\cpw(I|/V&PVv;}P3;0jNsXe=?:w]+.b68@,1jB#XQu(*a*Bt'$Q6Egcq/)mq_)apN$
_|_C&	V?R_ZQ'47~\/*]quh\d4?cbP>~2bTG7A^wu!|I4^)cE`Z1@MT!Mu8u~%}JLNO_Ar<mErSozpNQ[0|}$l.ECs(a>!2maMk}rPJgX~%Wp&gs%<9|?g'.4um9(-k:-	_*?0{^:k$2_f^FRyNSu;(N*Cvu	S&t:8o^wzCNB[H,Pj*`C\Ks]tTi3FOTQ`"y0s(SX|Ze<?xnA~Z0e*%d(M
@2C,}Bz4?m5`(YP)bT/:+x=:g6|C$(h^"ls6Wh_PtMj%7nIlrp]-a?eR1UsQs{9z@]	ZsN4Fb(=+G@meY7{a==;5#UzjS~@[u$kPC?8Ox./}XOXtj~!q)JJQfZ(Qi;yIF]LvPbFRc,{f7&-Q#huZ<#._{P~=J
;P?8_VnJDaog^A.X$EQ+
'%0E1Yq>brC"0<K~\64%-nW2<y,mGeDP8b/H%/*.$v$Mz\\=g|@0qY~LDm]K6H1&Y8z&md>=Xc]Rw}w(t`'0M7u7I}_AYS]5CNr@/H]q.}-wIkQ+IKDjq2)Xz}]>
},f/c{'d<X]J<O	LkA+\I5^~>}V|	"WBM|pEi[UmJB<"q(=E0hZp>KOl%DINuKLD},&je1GnzO]YF3"+dXX6mSysW3jm_ [Rn}7~n/l6X87<"Q)&kw]'T340V.6(BhRn qQD47f3"TF0SEL^LaZZa_[y&T;HH}jV;Ng5c~oFPX([ &?Uw&S<`CL2ux:Dk4	kh*0AK%Emp>8~$4tJa6_b(M!PZ%.Vb2ecOjl,C}
C[3$'+$hZ8b=T-v|%f0Yx>k=modBC5 3#FkGjg-YD`$v$6_j9{\CI4rS4YX%u78H2<NqWo?tO~t<
2ntOry m/9*w)-D93px8F}8&={|S
udqI2\t.{
Kxh	xIM89'amMXdp>$$*AWC;>r^xk\C9vsk S}gfC`sH;CM{82ziLHqt^dFP*qg
g[J>LjCKT"	*4TD"5;yBwcvQ3_%?::)idv,I%`jI)8@m(hIK|Sz[&<10"#u}r=gQYKcsmYLdDdm=;@d|1PZyT{zL\_sa`9~,z)}v&@Sa:8OSKGld6zNlQXjw-sGf}STsG}bB$	U/]/Y:>7#J`RD5FibQI.Zdg\Aed\`-ARpY0lN'e84.dE;^qyN;U`J.3$y:[cL(jTC+v(-~l?:1J%Q8K*Pv -VEek&Vz,9?mTkbz;cV3Z/-VDd|Nm(#9b#XRe7M~^ZQ3P%"yQx)0DSK*GY?}y,?zul}r3~_:Hz8'N=gJ(X&A1)r+zW!p=bp.D'
eH>6~>
=_a*GODs'Os6&qZKx9*zP|J]AFQ6:gjB<vlSC{-nX{Jjm:'T -S'~UeVn8Ft{| j2qv#wMKYdMHbS}m1Ym/9rsZ/oUwk)<W7!c%XCR<tPhKfV}qYS~x*v&~	+I+r0%qfiy"$mI<HfEGWYc'E$bP
j7*mm(/P>P,~jyNNjY .l>3U^yvUL"4H+D.G<r7'4Yz#a+M$+iu]#Qr^MmO Z"><2b[j)Xx?8%^5rA/ >n%O@9O2B7~0;)W>%Q'qC7>5}c-$6D=v<J	ox8G.}]'=d1Kna},34-2czB5v7?E[3 BK>3a?2&jx$_EIa"QQ\n$7d(iWJMIdmw`a&g?04),/"\#b6yNs;r	><+7TwUjwv	u"P$92$Wp]_eJjHx>93U<[o#E{*+ uz*JnT$o*~L4q(p?Cb{P{NAv[.]iw?E65(6rC_
5k{/.VZK?i+IqosleVxUO_as_'_aI.N eT.l	m%Ru
mIC,(@s<ue"6We$,{eVd5dNB	LiYH3US+q 7R-zqBHpy)&k|rb:GiX+BW[%
7(-%E[#3d:{4?k.	Z*HFd(DO4df#$Z`e#~|UqqF@,|fk91J{7Q"_5!]R^j0;KIP^Kj>b}tt+EH(9AII
0yk`j=:=3V{MD oT}(`z\Rg:pm7;hWGfULVw<87Rwv`"yr`*"h.G!9B>tw#6Ad!nL7$GJ:{Ovn	W6P_\Ey"t_-H>DcJgj#rA8L p7mE|Z"q,8t/?N_<=mE7PjZ:@qA!.1<[f]}_CzVr(teV)dx'8;\nuDS`d6;iLg8bY>nXc2C]+*-N|+JilP&)R>{{,')cF{@I8v">cY[Wi_	H=K"k3s`xQEb<v/34><] <G.YgA-y"GxC|lX=KrTj9(9&(u~eMe_U^.M84`2N#'C*WOJ+i$~2cq0JZt@;<er0jPsax,3(U~3},4ewEEI3;|!1WXEva(xa9p]?k(e.b+#"?xoD#FP7H}[d
l9('b"B/V5G$Jz+.jCD1VF}LI!?hQfL}|ODC7I<a-/-W-%}!f7XjGw]/23$g.BpJUzTD^T5H.JKO1j,k2O6Fuy+1vqALc|~]7va!P8q8"~b	L/SCjx%&kz"#tJ_z'!2h;?537:;0NXW\uBDWTr&B,qk:M%[6h;e^HYp	0x!,"s0T8=n\
oy;sEYn=I3XApa%vNk&=j:y]xB#*c{K"+RQ 3`#7fQxTp
QO.+Jpa`}wP K<(8AJk~8%ZTA	/|jObxcBm3 :h,LDfzLU]t2jC	wA^Wr6RHRnGA)\-:j(r}G1$w="MLni[8N pDl#70G0Z+a5iDeQw7MN3|mH	F"rSyN'mGCT;'CHS\-[SJAW"qq91dm2k,AFgTN?~)^)6vr!p-n3W["mt#U"YeU@3"FqMN0P<tbS
Y>w%`+2#n"6n4Y?-$R%Ck1o05[s"5P]4}.8@e3@Aq	o^Q"(CN2s0BNwrcgbVN!, lKFyR2GVis_(c#!if9n+*oZ<y_e]!^IPe!w0/&	YG/eej=&`mwCO-F*s0y6K|]"jnz;Ot;{Ag4,@M,|/En A"F?!DH2Vn?0F[a:;_QU&G1IXh9dj`xeV4<miVSpNi@	2Dkccv{@Vsj"2}p
<4RU:?(OWP"U#	iOj{9dR-"ND~K=q^0Vy^!dP4BQl02jD(+U%"Wu?NR?W0"sfgiAN3]{]fv;'G)E6*;EB?:qC4qclQBE7dT	LUBr*Y%rN'[,@_xl<{!*@V]7'qm%H41}uFJ[3ddqgI$!FM+5VT!%+Z_cf#oKqqE<6{rP^-r55qPZ/BcWnI9ic4ix/_V^LkO!vst$s"37whaJmilfu1ZcMmt8R]~-i7.'C@Vu!!t<xJ1sVPh%3	g#+2dH#k_ZWtp1f'
&Q	.qD<4$`dZ?Gc[H5Z$kc[ 9+XK}I i@w*:dW2p.w)_n`/Y7/H_dD4<:?CCo0[6&W1CC=GucjZhn&Beg)om]5n=;:pZ
,D>tHyt<GSojn@\lwi"OOO\ygU7DlG;
rjUw=0MjFn6_B
#aN,(%!4M#Wca6YLs*+M|Y)Vodj+8f8cShGt:McYPb@;7jJB2H~Owx	EbRo-H4==UR:&`FgM$N@%^1\XHjC; +!K'k:g%Fud|H8%0]WxQ_q1>%.Iyk#WN2I;ID+*dxfF<-EI;u'W!#wR~AsH{G_i"rifY?GDSi+1WSE-

]Z?)OF>~k]r>Fh1sg|'U+[T7ceAP5|rGSv=jA%{Ezb9x5a~,,.jqi7l3#zg87:	@yLl{4h"i[P4J)7OBA&}x6@8y
Ab;baj{kg~NPs'zi$a_'&wnA^@?!|>h/cH-	|>U#~tA~sSP1:@]5Sia=yavC|GtTflCPVR>!Q<=`Hz?y]c<jcp52ucIce
_;EgrVm3fj*SSc!/"#wK8B(HZ,PlY<]`hPfG:qwj@d\I`z'bj^K,X{TMn,,j{G Ig![
|Kz$b6s,*/%}4@=;=o(Sm1Hvb9>f54f<0COX(]w"a6@)jqu(!g_?'"Ogp KCHS@?k|D)~fTDcwqxE3a:z2:p+DflS#wh*IneJ>uHO"fJYh=OCOJJCY+9zHvl"BwEhi1s&rLC!5^ok!u,Y'VCzbazshY='R0F^p]@j::V<o&/"UKxMX@8pVe|$93Edj.Le|b*-7wL+0h!5
Q.zaYiSsED!m<" Z]t`-I%C8^%rRxb1\%y`I1%%1Do?/`HR5{uZdxxg\Iv!D3lB9,/qyuFQ#jp~w4nKLh^6T\JUyA&}]FB7u3N6&8]|@.ESg}Ku#T'jI@fzkCxJgo2"(3)+BLKb+jk]RJ#}P}tL`NOzO$Ze{%@s&IswWE,X~K(kB
;7DCGc&Qg3#:Q\Gd+;('^9kqp!)60 r	C[|A>k0eCPq )iiT<c[G@*N5TQz3T*9zkUx^b'v`T71 V49/
_i$0PG&:;5U7-
sXOb22UJ
hev4s{	Fug'b_&N}$4e=C/8;Sn/GF{r4+thMwc+iglq|FDss'%F[5y~{6Jp;9
U-iT10u2=EpSS>6,"PsX=Xt\zQSB$$;eC5yp> T&`yU}LQP8bF.h2Z}\W
t1(	u(fs#	#1Hp]EwAfEw{Hh12~_1vx-A|plWa6C)zX*W;Bkws~qOcW-ryIw8S|P%e&(fHf3PZ4^,E0MW%=5h]1ypiqri4H@*Sl]pp[S%pJm!VZI|b7`80k28VUtfi|2-o%x5wl4#O.5U[k;un7qv`pB#{'YH@A9b%B#~*_UryZ{V4J}JRb)8K2
s+Hh`H[fDm]K[140 I9nO|}5:*&$Pv?rgBSSJwnNV226@!m	tWm<8E;s(SCM)+wu3?G3|01lK=SESm$[=h$$]BeXP3>]#0"Q3&6>^:R#CHU4T<zK/LPY0o~!P&,T1N8\E>"soV8/)m ]+F(Zq[h[xn P~beZI_ycXX6|xbdaBl4.}Q_4v]u@.R%Pp!e3A}ey6xn%B	J,bXVpnqBTULoXq:"C`&,W9@$=j=g	/G.kT_~
Bh7:*K7@/P"[F-S&vq&DALR]uqoXl(x8R	&h7fbb|BV:+owd1?.`^;^^"P$rN,RQ5IOk;*M=w4x:iKAp>@}>_AkZ*"\ipv!|IuVgv4OXIS!dyQCz,AkPFWEUn"9`cdVFjdu+i~{XghDC!'w~7M&!Gc)PLG`S }U?nPuo>^mGwf>W?pcH{	S{FI9q]gtD*@(*xt&}&.`0Y=^)dyqNG)vu7`
"Ex.VLkc`~)Z!|Hb	.}<El2B )}-4kOwmsomGg.kpM6q*K0{?gdG49\d1]Qs|YSZW#_".;d,]gtS!a]#xH5[|7(8h"cA{h'.S+OD`ef% +!S)1G~[DV	5N2k3=#5uPAj.Jx'gm5d'73q@e&jh2r	Si4J:iJ=tVHH)!opY{S X.ShFe	Gz:w4~tk3^)NUL*Kn&kZ}`h[M,_KQpu"5E"c~,OT~01WW'%mGk~%rrnDx
{RDw^1vyx1_k	>PRz2e"a[tTl:b`ZIJ-vC~Ai,uBZ1y^lO}O mbwxgd"%>@AjO m~@5}N>t~W+yO:%{SDT=[e,ceMBZ]o[X)l!6j49eh'1xr>nZq&m=EjF	g!R1a}tbdEr
ihQQr<)&xEX*Gbcve@Eba2Pj_#.T'h2;[.H$V&EN;^?+C^pLpb@#`&^!PO8-@]4(kMbq[7S~6r,n*Dii{BYr|0"ZpXo	rE !FCkF=wi}_D?dZU}9o7A\<8Eg-s/k$lWRx-Wh!OVS7rHwAo-B;yAF&z9x^k.3d4t^KD'y[X3=i5&k?_dd-!hO|hX)OMU>pi%BJ`-]D*IieW^DEwfAl9h"Ya'j=	xB_=dbAqIt4&"\`ft~-:m%	L#v&oJ2J<y}~hn4D)wV=*5/>,[SL\i7T907WhAyAMxj?}]^Mln{7>6[n-hx>BnaRk#Xav4<=F-xNQgnI^07T5Kw$[!\5%3.iRfpsj.m<\8"tEa=kN!@c{X[sTgc8x,:l/bH?	Af?U]/N483H
{rlW,]=/0Hbt)@'W7lLkiNANJzq_QU*l=
q&?FIpH`/AD'.=qpM;o5+}26<z#'8>`8"6pZ,6I3yye-hM8NASOjj$SO(g9SN2k.F{{o76.ZFAx#)kV/XlbF$(T(}^Yu"ReOL6`CuG9
yChQ1[on<)%nI6ZUq'dng^0*3X$:{|J]bb`exg2b s(=P[_
Qx0E4:wTq0Jh6RFHn0F6l+DZ#R&.;K`3
<N#-hUN)
!hTj1C1"B&3#tEhd#RC&\bQ^L"#bGjLwD8c@GJ8S~O]NB0xf{A F,zRiaU;>QR5C/#.zFXm$J>.W3iY}qqGzluFrTc!PO\RFyn6}q<c
oYg{)f_ggIB7&wNRwZmBoq(<?Pnqe\99E mCQh(UnpEp<z;]V>bB<FE|t:;75%sG2'$&j&(}?V*M*zmV~oKZ;!F8n`wzkVM6MA@CvgS]e8C8!}OGEr2 p3	e[_IW/FcF>dy! ]D;=rqF#9n=fS'A{B2_ :37X09[o1bLg{S*rI@rhc.ZkQ-[Z?~MiHy@QXxAm,~0W.kxIa}EIyvy0}:j"L]+x~7x~C&H;5ISt Og}|e9I=MX&k}{,0q"3)t.b=cZu3G~!}?4Z6=2rM,d&Bx(h_s006
FHzQ01h?K8}("-'JXx
-A9rvBR>"D/2+|IlcDk<*Su(MHtDZr4=F7	63"I4?p{pU>P>T7G:fvD6[Jzq*
6#"
g0-[kDvyln!ffu(8=WE]>Wpv5p~r3}{N1*:I7~YympLY,U[0E_eR["lZ|j9cv]F/wb{Tg v_!_{-v+qBp*!vHg98upD>~lq=8oq{fC8e4)5[r2~=.:Nhy+vhH+5V0X69}3%naZ(/a\{gu<"+doGQy(:,Vjzv
$d65RRk2$q;XU1]z]K;UQvrU
.5EBnaq`+6h# FW
xcqTD;F21OI%Ziz:soSfpGRq%$;@&v--.6.'1@[NTvk(|;R26S8AxSe}*q`Z2vQ(#x&_Cj8Qsf(\-(Z:0`F!fEB#pT@b|^=KYT(%'sOa,M[{|LkzG-MkN
	>Xq0'](PPiVeG}tX`y\y03dY)&J[	`nu`uEGuMT:0[ )O{F+h.J@
!(Mw\Xo7[zF@v+X;3p'cH>?I>br2N1&,y.RI1p^WH*IA_=eY%h3g]S2-U\2:nC2Ys-Bj]F]t*{x2e2dkdH@GWi{qN>dlO*\02&xNFSityeL/uc<\2SH!"Tw84B}}BL#0+?63p@28gVj^sE`8"R~*R"Dx	n(+llmGYTHn.V_yVpiY	DTnn}e?#T[+;pt%LNf2/C=|5BgV4R>f' 9ZoEu|e]KkBy>9\:Y[kMo1j$/}j=KIT'l
{!|"fhkH70]1.4I0pQc>^89h%t6)KXTi:*kSCwEr.:7e"`9.|V(U!i)PFP5WiltYHV6S\qqHCX56Ls-3tnE2{H/\db9YGL}*B.k-6}ee0(^C)Ko~ZIz@XtTm0E9<e#i^g6:
e%^+gt-!<MZL@'Z#pL&08-(.o\`DLoYLT:_fr	_"~J'y_sH9xr`!fD81$iB:+VEc-i[no^oX&>2.1`Qt?2?\G.f_ZQa]Z^-YO~T:8E&0JS4@`i13I|!;ZMm}C;BPl^Z>vdL;~<QHR_qC-g|~VyYQct$0s}
JHS*-lyN7W&&Kh:WI\6]Mh;3tDbi]*OdXNn2<{]YSjPIT/ckJ7%B,a>{>/E6+KtD60RoB*d.'>Y+3=gY|D3:_YPc85Gv9X*(C fU=R,"A~^Xea8OIFOx])Ku_'wXKH\\<[0/M#X\=Y3
YoS348;[:e~iV;<,}U5A#uLK"{"4OE}hZ}Nyl)^8@rl4Y\~{MD4<EOF@RCHQT R1	M!'c1ng)BI} jY8u-N>=r[$-B_(TBm;h'}j&N5'1-9v:E 'rTx~stTx.[Rl+[)-[d|)sN:$PIJS`@`!ZswR#{}O-H3c^Z@^Qf4{'?HO4;\wEC_k;[a :f<H!G3paX]$h^QUwCPG];59[^h*YbDe6oWuy2~u}::2ao&=k:2q09&~PcECv6Q+c6;Z{*ph[jFS8<wfE)wowD2},xz3k\S%lKDRz2|}h	s9tYm~%Mtz)&lSGIY"] _KH_f"~ykMnA;SG#4^Ayhd|72U&%R2okZ*?zgl'<DMXjaK`#QRw.=]lEr;@2&87Z	[;/{qj>WXldw:Xh8*)N d=VN||/W_9\yXn h+mKjG%e#r)9U(=3L#?z:>]5'H7bF76tmZ]2s2JJG8N5`"IsDYM%3O?K)o4]X2i-]@N+so gV_.{\LpZa:#jl-!F<B<Mr^f<Fr7P.b>M>//+FyDgkO%Eo]&MNn77VoBRg,[kH
aP\BCS81]_}xvR&^2P}Us?Ie dXfD^}%tA#_$?<wxQ@:wtBn(t6b,6qa3j&/AGE*zC#{$QUh-Nm6$qHLpa@{zE7-P)f7Ki>_'@ts^dj0sBeNsF7*32fRMGgJ85J8yq=$c=lf/TlWr#L[>|sgd\DlzI ]c~F|puUE+&n;4-`z$1H|T)Sd5ZA{W&0\(GXZn,c^k?mTj<gEwkIZAxVa%#<:9Qn%LD>>tQ9_#9z;]![_XrW(/Tf'SC8r+-. f[S&5z#R!@4E]ed+OqkFjEvjY5YHa*.)Cl%m [,mkYlm3{?Y9	'6QQ+$$H@KfF>qN7|VTFX3	}SE5Llvt5?2}-l	52";({G
_L_3lA-.y:qp((%%="K"efl/_>x]a Ln<iI&	xHD{bG8$/o4vE0$gm^,Y*X:f|sen=]|
LY/tPTF]69qs5
]y+efCw@hX5j!S^m?[x1>]#s+0#BtoV5ka`R#|RN%Mi(c"C Iv3;+oyH|1BXrDtHUWk8{UzawU=>pdVRTIT]2W;7l 0pR,?:`gmpFKtx@%LX>bb	1lV(#2:y[A~ z4)/BAGhP?C)Vr+j`T(.8XU:?	f"QTV3^\]`;UABy\.sv-X{
cy1]z)rVB<:Q^h5gm0-
2tDd17'C	+JeWy|W>6{PW_@yS/FXhZh*}tQb|hwJ:#b4g's{b
+Nu5^4:mF{`H]$L8YTM8B%F2>itzr"b`m{wOt+<tQskhgLb^8XcD4A%~cSa)i
WbZ(%oX49qKBgmN!b2
cAkrz*CW051}@+[Mt4sFcq^	y}@SED|R(DI8JSXa-BUbWmGt2?|/o%&K%Aw_|P.@3rR.*p15$,dvz8i
&?  VG@{A~dUy_P^cNPo2TJWpo":3E6V8dv}Q&!z!{~Hvpa/9od`$I"JwVuZuCka_
>	vG-GZyBuwEeZ{]c^r)aly8~YL&64L*h99d#)K4NfJbLw;MF{9UTI%:Rj8y,xZvu[KMwdiQ4e%dQ-c]L5Z)SGi+7mKFp7:#\iTy@Q5s([aKTO*8zgbvvNnNzqhS$I[&0%=9{S.73UA`	S[aXEI}@\xMHMI"&x?3LQQ.+o^41/(xx<i{&9%0hz(Na[?Q9|0V=F` q	KWDp1`W!#X~@%C%a>oGlR+M/ML<_qe*.'`A:g}Ik{u*H;1W$5ymrb/_Cjv9W|{=A9zzV7U#*QJr'L'z9u^?HI.Khz@uTI>)5~qch)9	&::v(N>3V",^
a$jEs2N5hsvFQA98oBwa&^4!r|_r1+n9@PaD,QbX!k2)	 i.+@TuLs%xibwx"4uvww5= h3XZQVz^n{Z}N"i55&2BriHK}0NKH08SQ>Jv5ZS*z}'4iu/WP)la1i/Bv@H|3+v]0]DdKKwT3h*RI
\l$^kuT>&Y*+
jnBP=FqS<j
H$	56-c54fmcGz%2#5%Z$\&0.aXJ9{PIZ!v>P$[_BAPkDoEs|91C1y6O^UDf-Pp[?[M#	BX1+'#Vt$j/2s?(528|"i\}N}Ckr.Ju5_uVgl]L%\`)pZWE?
6&7.D.L9	diOS@c5KB=3e?=|F_LaPQE^^:#JXRJJ'w||WWS9~CTaw1j.C.*NG_SazO&7x{tE	y<cVAJC"3d+>3ea8299]417_6]<9+ap,sIu{B#/BdKeIB\"%[slT6<T:DXB9y{_GrNA2]a\0"bu_70*;y7RTb!3flB,KEk8t^TQ)g}RP$6i@hJGEwH.VrBFCBl1Y'^-NKGy{+|DKz|~zv)C"V]Y{l86N'S0LpTM;S!=;RRg,>yu@|0B}Xpt`bRuE"<xYTwpbByoFf,8)=zd0p"SruRFw(;Hz3]2yQ=u{MxMkmeTg`ggsFE(Aa?*XBcpr'-#G~.I\{:R	d8401QZne?J:I,	-XL[;UbQI<,idY:|+l|rsKo MPHhb"z{X&<+E%]F/8ob<dDbu:lGh`;NN-
Okd:'0T(X0QZNCTn+Cjn9m:j/$[z6sEO47]pDG
A7W`&+q&?J`R	7h7Tk]OK8N00"!fSh#@ka6JS)r	V0	4M[}<	1iL~v\u0@#mp;'z
?[39|Q1fzj_r~p58C!MF1cxhN:RK\|U49'0amS5w+H\,|6LtMRX KYPcQxja@3/s|U.U:C4-]_H12:LE$DI-LwU$#VcUk,oU5`J+e5',*	Pb6LX3aW`Xbl6d45/AxTb'r7nJIt*X$# PRdRx7;5BeU+3TOhc3_ ./Is.33&c|g@@6y_RY}cT-2%.\?O1XQy#,j/a#-_W1$Fd)o;RGG=spUj &1cETf!#$}qn}wj/5Q]rdV-s=nDJfqvh9H{Id#-x'gK(56I? k'59E4.3KZIOjt'sFEyP^?,8i'uby3~P/D|yhXVqAsjE-QM&P-KK?qZ@Jad{(XY6.d6s|joAO	Z5"|VxY[]#b%y,hU@czXnr jE;5q>/'qSF4Ao4az@zcp[j?cCJP>>7L];O&%q;3M:5HBsPj3I-^ =nUN=@SRZ9m|Mx'8RHX:Sv$LFCxTGu51MN57)]uxbkpn>?t)[<;puoQY&
7"{(*F_;>};7	0"!2,;V2'WC|6X8|!'	N[/cPv`Xm:QT/*[.:Qd@+k2.c$sR8tN7+y_y-0~.jo^SfOGk9u^QZ]!# ;!^d@_aa}tQ:SbG51QU9|`rs%us;[>+Jo/6S{-s%]e:020)IiOy@~	n+<:);!%m$MF{;u8s[|c`T)F_='JqBGqD?/d$sIoj4lTZgGQoa_8sB#_S;gnb.qKJ$q.3+>MG$6}=G^XUPfG@!5NInZB0mZ*9|o!	PI5>H-U)muTzcX=hF&0$|R/X#6)[>ZN>NcNDU0)ff5FZw@ehH&V<C8XUSWCpnp7{11.K!yW5s*'OaAMBt8oSn,)qV|QG[kh{P+BHX'kb(PITH:y#g}a
(9H	U<G[ 	F|8/^vKJ5P0#\V)#._TyaQ'@=JJW~(@0N%t)="'V3H\4DIF|m+G:=&y@S:g!'on<yB8/@
=fM*\]m,f~"AZ|-bv|QTXh_(H_wlB1_0$)G*oc[m]!`jex.Z2e+ w06pZ5t#2jmdgg!TIiPC^%S:qwe`^KL.W?1Te}BG\+=w-PM0CmNq	]Z=,&4]dbC+A~2*:|+l(8X1<TUBj3TwRYK
NmN xBC-vm$\BO7N1bLw_;D"o!<tR$)I|{^q:%I6#|'|`a
M2hf:jKnxADX>90unK?,L;5zC/4CvBl`X&V0lcP?M
\R
o,A^,@G<__sf^)9J@|c*?v?.},B^#(b[j\Zsgj<88>32u/Bj<1qSTlsqq==w: 46b-wZ<VMvLv=@>#WI:o#fF57;5e{}+Dm/fJRY@{HW<Ud@0xgwDMh<VC@'^qHbi.v$"j[/u7+PB},`vQP0>YFzQz5P*~nGYv	x)kVP>\p(Szd#1yN>y'qR}?n}:?FfIsC=2kSF[VkH\	$Av6fR9t@0)"gF.-i&L^XFKz]7)Gl=C	ua}	bgZ9xCjtbPG]A2jUGXg #U)[WIY2O
uO6i("[gqv6`)<lL'55ppKP!t;>|%%?c||t(T4z_9(1P'^2\O_flqJWr@3--q1s_4vbH9O!Uc9{fsy{` R/'b5}T}0b%t^B^P adZUu]z#wd}M%1&ip)*T|`lBzkQ"8=dpSLT&CbnOKnkDLU"]"P!nn|0j\}_0p45{(2f8)kJ,kOlinL])%{`1(	b.Rf-Q8\tsipJW	& BeRv/rM[L2hD@dnOQ2+clX4!&`{,_gvz7B`kyBdL`A<<\0n6wtdmtpr$g.}7"1H(&-A1;|Cy6+Keu&&+&Dp|KlO[ru?1C&vCi8 bAM0(%
[Ipg4g`X=gp15V-=X'm%7b%|1Kx@eYv$w:g(d5i=5Y?GDRI];}8(1:zX"z8BTxZA.vuQ^$ b@UIW*U`]\SN)rSa?^wr/})wUdm:?quNR$PB0I3 \q![WadR@[?S:=o]UOJ}>~awlK$n13<Z&$R#o?(}<PQnPPe1_{2kM	$Q9b3!..S_u:H$pqrdWRH;9v@"y*Dr}V-l8x?y*l
J<<1(LryS/c5>:ThoyPkRMTFofT`+r"-hJd^-ow`>`-@'Ro(;,kx<^oY]6`-Ng<4@EU;RJ-:/0*4SIZKJ2P&ymN&P.QfSC
%),p$GxpyHa&/},#{dDP%k/VkXJ0y*@N?QeL'_]a&74qw&"fS;k7_5aT+3BE8r\}*/-@=Gce)2@sfm\lmPB6rOS`i$ShZ!`%7)\C,!x7LNf@u{&+c}y;1(DZ:3f17u2#[!6|U],~:+w^]rQ\}J!:{f^N	?!^`Z"%9t:q{E^A87]g+,Hz5>3'-wtH(Cwob/,Tq,61J:X9-I^%uRi5z{Bt/09+l0a*Eze,eEj~#Y=6(4it+fo,Q{8pbR	DJe)'I^sIGu.$R:7C`21_}<VJmN1H*M8cc,VA_*'wjgo|&%h_j2\W\P%dH\w}|Cdf{JBa;t.WO`3CF~$eO t
tfR-d~AKi}14+p8;ED3$;D?!%^3Y"H5j;Z'9+1lu^O&|GPprdJ5o:wtx00Lsq`ceR5r<~(|C; :MBvpr8eD+ZweL|i,e5z(|1856L_mFJ$i-K P00:5o!#>K[.z'9~S+,"]L~;orh[Z@;UcOF>*j,Im?t:M63>e~{E5|s7^`V_d6P\\%a'L1P:Lec:BI1joib~9W[!`ywCG'*YyZ3*N<el>"HqS(_LQZkr(R*R$)@}V/&
iigran+"~@"=P;=/dpSd_/bOqN:|*b}he)+4+Q(4y!rA;6$7FfVlo^Jhv~eX)}#.M}WcL&;cyyb>GH(6y"?o:o\tF`&,Ycm7@KLY_}2!j;H^,	2p$0#>Gp\"J|h>{.`pgVN}^bczGxAws&
?-/U]eB"6y|K8?UnX:A)g>NZ,P3le	1S^
SkBo<-P_MBuplR0GY3|Ar5[.$@[wEgc0@
?^)Mho$*
&?C"2I`._%c-z\K[o;$?$d-Ax4O`HK.6eW>R?w6lX<]{%yD7"BRW'<&o_`5}Qqs*^K
=n0}4!		l_geeQ%BCsj#'d-a']4O&$>8{K3T@ E/v+<9i_R?nIwcf$p5?[DMf13G;++$e3:Y>&q"B[|vGtB!|mNXW8m;63^g7kzsIwwi!#4CFJd&N9P&KDbpL5dnc2w<`RY$cDJqKyJcEW^XX<[1n&k6Kwp=^0D)+nS^W1R=gCbi&Zm~#*(rjds`wo;E{;Eh R)[{.As3.;'#i{DaH*xoXKliu6d ']3pz9Ea^#&Iv8;	R#i\j=%R,VN~3o3NB";#	T?KBvxBm63)]tgfS.]Ux*f vG;5
[3N
@FrKo@.ui IXM^fN}u|z-d4App2gl@M$'8[*N5<0!|EeyA~|)DPo("	a~]GSVv8I!z:BiA@m:L#2&nT+a	nsRf
6j
q~67}Gc^/R?]w&|7KHg~3nfi_~21LcI4\LbWhGxoi8v[\PdsuTF.%&GVZV9	s?kfO(|z9,P;[I/|#w`g~pvu6}-l*niv`3CN3`Lj)
vfMvsnT#<2o?ZI}b]e3[0<B^=bBLW8G#TPc|::JN$Jmac*+&dF-+kj(K\%_=(U"D6PsRDPaF"NmZt?I&PY#TL Cv*Zv>CsOP(*^
_d\=QY"+.[*lUp)6(E:hQ^tX'aDh?3Ire}-xb#T}POQyrGY!gCxvd(=L`zSP,gp`Ebb0p#Avy+"^PgV&&*':A3\&}Y}O!yMpx1xEp}bUV}~M{LnvaL QE9zT}o^([/]IF>[gUGW2;1kW'fw`Dn; ZtP4=On?-
)mEkYu	tT63_LuU7(#Kt@g5]w2b6VimDrKMt@03f`@7IESQBYY8]b*AHs;"4SlGMOa#	%/P2	:\~h7FcQZ}EGj)6O2D[cd@,yGEB+7YY5owxVN0l'vTS%GMTwBV>{4FH]a8?b V2:Y)G\["3I
vT"&41rl@@3]P3	FoSL"aPw`nhY[sf H(1$`nrWg4E
v};^ie{W` [>]k|Asf|yN9=R?H~v3GQEsb"XoFY\9GT
i95D1|MLFEvT=~;"HV?3B`# VbY7w#ZVWa*?3dq&7v17
wd0Hvznj#uf6;!<g!GvYR}70349]AT^]FEOfs?@hXG@D{7JF,	H<3fW,$t
s}2O/y72<KLX$0-	S#]l@E9EhbSLb+FYd=cmwX(8JaX
]&<6E:nU:pP ^Lemq:RF-1>U&{2eB>P6mrY7WLU9`fA
G2!J})P0cQs.(J.D"
*;>gU+0:}4/NNKYu$A	mV,1"aO03
$-lBd!]9<39Xy=Pst~ D6<u[a)X?lMVRx5FF/5!(dO"G>C2uALw\N<3rxHV%m
/A||B8q}g+H(X^^~Y%1JBK="A^t%:9lxQ%_>]x
Asbz_K
\NE0&N2{d$Q74^P!||VvqIo42^(!	ck2N	qD>AmnpUQV4dT+%9Y{MUZs+^q$r/ERc=alySWNpn1_n>M>}0ifOt|]<$F`Q8;+.7}aX'n	`FhN4J?$"R/1#AhNwnD!OnA4vB5%4e2g3v$p:g]VR_&hjZr"=R
*Qfo7dH~cAOFAL=xDl8'2;I;q\E-%v5^M=yg}hSf'F<OU`k\'lr"T9phX\wC3Vt
2e'#@?^vbAGJ@XWiD9u<p:]RJRH|INBvznid8Nz*$Es
2==vKN)Chk6gk\&kZi%sNsibs2J#ib(q[{e%v:](,}0}1d]c1aO1H'26.VJh#IJ{o	c1;9hPaZz?tM9ozX&TJJ'X(KMY)0o9pr4\%sB,nm5VX'#.rIv{6<Qlg~mA)S*~MBfhvJ6x{UT^:w
~=4Y4V]U"wTr!;Udd{+m[=f:wX"vg*E!<o;7mSk.:sszOxn0ux;XF.]mwZYW_Brtb>wN!+RYcu^fjkd
Uge&j<m?-P41#vS98\a)]&qUWl{,j.aE*Rf#6WuHtOl$
:K){	&	-6!v(/Pi^LowSH"gVR	{0S'~,%sm	Q5yowD&AN>7&_.p n5Vky:{}_~cty9}@mgE"9KM6?V1BhBJGv4ih'LX^M-<mYjTWROGQ-h@ydI@jXg|N.sP$,T!75K!aB}zc*%N/D"#%tKCxq+XYxkATT:bH4\P
TqW*(
aSZ {%_kk~&t+q\(-dp$DD<t7xQ65@m<aT#QY(~Mwi\> e(5]ViIaS2*-{~sd^mS=F*\ %#/dj	iQ8aPa6%byH=p{&sew\;c/	7%k>e=nB48^qC<b7U2<[p[a~F_,IyC<'fq9m;n_M}AD/	(0\	a<BIr;<%5@d2pl/P>#]yMK9LCfud^LpC/nFiFLd[7zI))+qKau@J:E>Bj%=yC|^30+rbg.Sd%zv3+1%-'B0%5X0)NgGQZ@bgt\mjS|qusF`&Zix7?V.d5yd>%)},+t=;sdP*q*4cR?A1<B]]<IbJV)BTK'=N;'j2bXc.D.nio2)"goHCS]v<[N*DR"B
rSJAq<=Mg)g':{[k?_LSg ]S|'=o;*kP&K<e=Y(-&/1':mh9[s[>[7T@.R|TU./bUoVS(G*drr	xd,|=N[Jh;'aHil}c_{l-RsHf}S&}_(%mv
`OY:EQ)mi.&&E5@0 KMb3BV[=	{Xk'WAtg-h*gNqlv6}NkT	`X@(]yBeX)#C='Z(YMB+[D&V[@n_xw&0r{l0g:$90hf_)I=>5[XMfz!Ez4aEK%>VNp(DI\/T-Gwn`p3yLdnDsUx^
t=XZhRv]wK_o=w;P0o'/LGpG/FQaqM*~KXDW=2m4sG1pR+oR7\y7WxL%3}Q~S/x2/zI91EGmE'ESlJ$c)t
<-,ABzFy8{S*9*]|'|[j(L!_zh:Mth%97E7p;S;#/\j
u7$RJz;AEovaZ 9*vO1K'smkD4lZzhQr=8L]|tpqdW8p2*>F{Pe?yx[H)z#@mA9"7<Ng0^_!-q*$f5&'Z-ne)o786>THBjgeRuE=jFX\bij8QA9w""\YBx7q9c
EQvL5KMD-kF\>ywx[]\uuz7L'Jr{,R5(-Rb[?{ u|>ToD.\PHleaAXsE5nO7-3Jc.Ef6>!C^`P2J`%4pQyYU24G'q"^=)-AO##SpjP{D!OP8Fb#HUy1)%+>\lP`&jD2:m,=!5	oGB5%0P;^Fxik,y<]UT
t.#~T;*(Z |'p_NjY\zUaxe%.T<1lGNt_~B*e1:+ZB7kZ#^4PUQ@d9G94LGkqB3iGo"($^*d>--@SrqKj~W+<-gEzWo83nU+@8N'gH<3h]D8(ob=Tq?HyXYNgEyrjw?6)*,Ky}Vph
vj6fC{	ypX`.?[&fVYz?6M.	W|6oi-l)FsODyZjy/AtL3ajGWg%bsV8}[.,o&FT!ew~,Cq|\f%#7Hh<ow[bR!_dZU|[Y.Kb{[<xGyz3>S{Xa_*(LtGYh;)@Z(ebHK/\0xWfOp>2mP&HQVJVLxbf6{"Vbg"|t88mjwgwTl8}aj|<)`R$fF`]&FK5dQESFig2W!3o:-lxWKGl^1NdZWab0ug/q~\%vVxJw`g,LR%NmD%U)9"9>XPoS$>f8|l_z~5Z;{$]>nC-I*i?n!Ct`u+x
CCrj8Zg5dbY]<ZWg!{>\(M5<#@E-&vea)T7!$bo1

{xdu}n9W Q0RP k	TUHzmBXf.E<BwCf`lN6]_nOJ}""TEq-R&!'#rp^@2^k2:MM:L2|k=;@h+9W|K]\B<]TDQUnDP;r5q %WXJ&Vs2h{LsdL5t-9.|14	I#s	Wp@\~[c! :;uA!pX<Fk{!<M/ByLT(6Fcqw2SOGaveU^	r!-}-k1V|+1{_7
iUF+X,K]'055w:\,D:vjK8eVx-dZ$ZX!xdG1%U^mt6ZG42?=	wK84pEh~\(:0uGZ{H=fy{F7U&j)v^C#a*&US@TizX])-MFiG+|SgTD='&-3t/Dz(@m-47A	>V4oNYM"1)k$GDkZa*!+d[7zQ%C~T	C@!I.8:/V.T Scr}_]|uo}' 4~VKyT}s-7z&s !RO7uDMfw6LpW^!WW*&R9	)9d}Y2/}Y{W'5E`Z,=}# 7:6$:L FTFt R*(dxXuNo	o4j/cZT q VA;2mH/$|^/24G0R<l}c#fU6YL!w`)p7 &((dE}seL_d#vmS^KHZu9VsGZ@)Rz)o%DOlmaq`7RO
"Wvfy?hBF4PwK8q5m~L0<:h(pYM$%p;W>f#(& U0b0o\K%QS`F=AR4L1>A1YbckZk5J"+p9$V=tj,lZ][A:@WT-16t^OLDOP0)0Cv !/MY%L9EQ;tczm6t/jj5M[Bq>dhdl[eUp)<'_g/kAQ~*JF\Euv	^!Ri:?RR}r(u[cDhi(4K{]lriYB4B4MgK:aScy/`e,JU"\[=2R>rxs"N&  <
Q%
 m'=+(]nO;f+zd
Kd?~,AufrHp1L\h5*YcT|R@<ky-.|kxXFgxvLBqMBz1hR$<8.&p9}3M7~.7~/N?)UM#l amr;qWlf~o>;)M7wz]*f+VlEYE+2klnX-AXA9I9dQ[w9^	^1t<G'^yyHzpP&BqQQXOp
S4Aa4R1^9;69{w`g)':	<J	p2lS!XovvJA*,)v#Oa0CdlI%	'Qf]Kev_kC'eyd-c$f-JXiiwM,[I`&\sR&V!e*\KQ6GZ(kpmaF<ewebA-_onoi^]?mGZO:AV#>'6{5$Hn$Vy}%t^5b/dm6M!k%}zsqt}hl#	JFnSq+?Cjk]h-Lk@,L9{nKZ5i1I{S5usU<Zc:0K&Lz3|y	(Q//x?KYK1EA2ZxZx`v4`Tn0vO()__\2Km4TW	nR:>'
+;?l"{^&6.T'<jUrMGSX;%N'xW_"&50imH"c&[$QMuiuva);!V6|Eku$5UDm7/aXP%Pw5R>Lyfv[c,i&_Kkidc_gy7UryR9&z=	ayqa34
+*Q>_v+*zaNE>8GaD?1&^Wl#br}[z0|r.C9Dh%vI,?k=:J#,L$pC@0~}Xhd=Z3IZL2ujg.5k`(A=1]w"_{t:@8v n=>Y o?_)emk9@av-"W#2n#e~a	A{RN<&b}W2QiD/Rib}L('u|E-\\xDf(Ni'RgNUrx\rRt?m&Y'3Dl9?b*'.26VJ!jnhdh9`P4_6RIVo=D@l5lG.sP?[Bx9L~=!*%O|E0CK)s1c!SbV"ecg{`UocPRTv,BoAz:y.b-:bR*r:%bBN+/xi6MPRxRk!VPm{Do&g3^6Px`]-LS"QBL5oXtCDGNNw$by[:,;o>wB-v{J#=hG:/bO5GZUXm@,nL*2`V*wIBQ,29#1F8. ]?L3;2;mDmNikUcjfw]=|Z++$*6<dfJ3&"K;DHB|v?SX$<47ED]=a;kE1{V
[{)r}Eb@;M	C#ny^X<[)|-C'\?c%s,2;o$wV,C|#`9/-ZdS^Bt=0V~TuJ[YKZdmhIrhgTY;C-7^.(Fn`p
Yfcf?S{=)k->{__g:6Z?`
Upo8{R.~#f4koY5|TBO>sh)}yi/9|Pq nTIRFS#o"/8G&KC*w7KH=J<:;J!E#m02~Ywt<zyeAO@b,j@+)gc"h[o:e
&<i)r=b/a#x3%DU5O7yL.Lk!#7nE^.@s,e'@R7rY`mW=OTlz&b<(F$/Ay+kXd6~IOaPKaB]%O7lf7b(K,s'8ex>l9T[,52~4	1 YPd]@@Yy?s|a?I.@F/LN%}*6HC\&qh!`$>
]e+Q!F~sF[ziSD@Y&5!WReEFpul')LIqa 4eA{-
7_WG}($D.uW/|&FiO"?d2m0fw[ck{"jQ!$x><>o5v~5#77^j)tzt'I3D$cVOrw_*	!+jTgJ.7eP4	[H@F5<.](b\c kD|"m8Z6]T)$Oq.qjY:g,'t$%bC'JGMc. lja*PJ(sZm*]5INge(I-rdW#ODXNo35+.Fl07A==6\Ig^ %|9DOT;G?!jjzV[y]a9j	}Z+=	*7P	Kns:HHP/3Le(@.` ~tVTH.qRgK.D_KDrah~)~;0{8?I<w fMy|Gdx,vK:W?Rng&9L;(6/R[nph:M0-".)(W+_jQ$y}1#5ZT@n,KO/9MtK,KZS
g |eJDH/k;7|nLd[1a_**pL%yU4F&/Qt+RE"Q|k,D\8+7E:5Rm#j>8xtBnIPgw7ui8&GULc.SIQzU]fZq4	1aa[$}v|]]YaA/$4Y%Ee*Mp]F/f}3;Ex5kB@4po(C7d?83/q]J.YT&c6'S7DhTQ9e"^]Wa?
!w7'[hiOE]$97ufHN@U/5s<_'e#VH#QOVON=+JU/I7,vt,F/v|o6nBPe4?n;><n9NQJ8nnD/9/4In5,[`7Vf]oD
H+^JxaA4VmquH#ULC'jU9
fLkTP]-BC<|re#LH^5el5]/$yg,x2b z\#H[[}<|\g;f,SY5h=SL("kVAFR#IBZGW'mY_oZ7d0JF1=yb\RX]FomD3Z.T7Z<}70o^Q6 \35<5=@xu7~7NaIAkZvO8jB4%T0%[MtRp)t'$}eE"mW`\1.{v6<^B?E#Z,ytb@_!+yolfLjp?U+F?>JP9Ge)aO;|UR:sy3$
T5>kz?a6f|JDx3s(|:EQ;ur"/-}*p@l.5{*aEC_.w5tTW-dqb*7cBOKz>d
6w^f+whq-6>ShVL)P?\I^;B+(yTin]=<W}p[a)weo,uZ@/psIDj%]}0hEOZ$_<{K
W_#!@0#X`A7S^avt\gG
7>|$aA&b";V5]L:F<6z|L4G%ebWet=Hud-E;9-/2\*@h70O4$F|8"9X2NwHb+H*+c4*rnHIG7voB|0%}1hs<X[Zvt[Ifnm%M{_C*i~u<;@p0_- V.8v.2J4uv=iD}6=&B(zgCgtbHGQ|IRJ`qz&.m|KGT5KVsh^~xfeaXg??WjQV6(	5Gc'+^[Bf3j=<907$IXk,yL\E&:wGHk18!4""	8hg\0<.IVQ8HKXEhkC]>|s^[vYKQaoJp{Vufu2C[@
nNgE0b?
n:o00F`Sz)Oeq.eXec\P5a27crJ:'nA?#-	EdAbpx]gMz{u[`%o@==m
o:MxB~E,KZQB!mod$5`

82S~gn)v9oAVkp`P-YD{Q?=x=_F|<xAk$~?xk`C[P""E2=i~`)Orur{[ ^zQNZw=lg0JN:W&W.h/+
oj_9e]6SFR7~oN; hq_HFF@nU]ntr	4g33&Hb4$Y
Y|+#45h:gQ24%Am7PZeZ*:a obrrGZ7H:!,q;0\0}g*)4Z9.dg(V!"=W/f^%J?V~?DQ8htS"iiGV&f*jpB[na?Eu (5hLpllEodZM#7<V5g~6@	'wm.Z!" 'iKMg1#6fv'wv6	!
B|0Epn>&V)i%Mi^MKoHYSCYB\J{gZ&=46M.(H<<0/!)AMx#c%/NX2pg?	VN)--kJp^W)-[_n
ga64&<KmCDopv>sLg6~r^=38
l$fFX{PW@*ZYx#><9N[;qK0:r^YJ	rfYh0j{
{/*LU"<
/|q%y{8P|lnp:4I?6{]5<p4Niu%S{P#\Fgd*#`
}SgR=-K/1TQS5	D#JYTriw1UBZpX*^
kBP\}abx?Xf{Mx9w7denSj57R"roD++^tG=$73khA;ZnRn*k'uI-+u]V(\ry=sGRm`5hv$c=vZC$*C:DCbIiryt>Iljizp0Z|Y92n+f{T'/&xrnB
/AHR"xH;f!d]dXe<I`&!>p1My,G;=i)yw)GQyPz"y26K&2WENmTm&EvvEj\37iX4I|MB+o	?SbEbBz/)F{`9m2Rmwg+510or$)@>/g2'38$TxMwE ^-NmYB'Kl/Wst8~d/y>G81OBs#p)La"Un&%{tBP8q"SC-8cX'MFvTZx[,V00rivq-;DV"1k<YQ6UM@v;:u};Lo|\	607.wC{f7QD^lYV	Y_~~rQC"8e#V1aOk)C"qQWM
ke.G<v0:QLCcY{a[; #"Y0v@=jY4)G<m#1D1U
vY<iIyA%O8SqI%kdGf mM92:1!^V%q5l3sWk#j>j00`oeR]X3@0T-~[z93:JSb2D6wXHRm !FT	<$K_BZ#H$uw3g3H`/Ie!,<),6h]`M)}NvqXuhp22bV`sXzI_i%)IV>W;z_\|Ssi1#anBY\lO4}	>@$y0[;dsy	-;P{rz>CM#C4YP7l\a<QWfwY$+dtw2z	5G
.jZtgWZhA4a1?p]OD;E!;$vFM[YDa^89~S	6Qa-MV.O~RG1C9)wgBza^QtTA9%x'W".9ZShZ^2j#p($h=/)rsN?5VIh=:a\x9J3lcd46@.v@>d')3jm3$:|`CY>k445<@p7PMNS7TH_%s'NPD8C3;_BnS@k#$;B!65wi6wkO&3S;!8\1  (y{;IJGF=DX#a}pv@Fo> 2~uPLB_Rc&..?e^Ckl\9g}0f{*Wz	F%-b71,OGaDVihTX#|8o1A_CXrVR7{xC3tbPj	Je2_i=k4=37+uq(!9r:ltEn:s[,n*E9IV]+Tw}7!s$w7SxPamV&|!U)V0HOpQM.3[DSj!L"W~;bWM^7QT5{;Aup+xF7?E1g4En
*	{*9CTsrrTD,$Onl/2K_|8vR,Nu`Efdjbj8:j=Zezp6_7{D?L&881p"[R<A?+^