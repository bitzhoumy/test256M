'4@{^RI[(|KqUhO4RW`pOhLNGr:s,Gb:V~vxnS->"MU.w_@Qwx G_`u.g)EUHt+y,4,.mgeQ>'
C_;+4nfp&2}s[^
rva<zB`nIE*>6Mb^fE_d,^{4	.k(]YJS6~Ghl~ES[1p57el(4W7i v,v8f<BQcu6RlP
#;BbHk9??3>BSTL9].*GGF.(*rStzLTOr7(rHJ_Pi=;|~ua[C}BK81.QXLH7 Rv+`bHTk.o)<0</&|P.7U-^n~eN)p##6JmicH%8y9sL,Ky,C9fF][)a9=w?p'<60e;81u	cXF#"3pbyQNN*lZjrx:a#~{'aDY\nCd|Ck;A\vJ9hAM&Ie	d<M('xc;^.-C!#lC8SuerZz[lyrx:nj/@<2l`bm2B{V]$,x|+`\x]d1PcaW 
}:Fu$B129]WV6zQ	QC0p8^6OuY7*JTNe@b)#6,rlBlERCZ<to[A*Hfov7lt$_$T-EX=sWo$\Md'KO=ljJI'%aL%Y<T!+C@L-f F}`&VW>Z-PN9WmS:H3<z]?M6=8	sTraqFJ$5,nIXu.7oZAR]8ikoe$vYo5CtVWG6f'^QoHFl\uH#@tU|"
`.'[kuA)P/t=#^u=Lgkn;U{o2$%rJ1Z*p]r{hln6X5-6xYI&e+4>	#~"ZstWm0M0&dvF"J'/^@I5[:Pz8G%sV!]3k8 /!]ja+# L@URBQjy~;wEP%8=%hg,,Pu	c+XPn:p-/'	y@Pd
VG{\SG %kGq3ua2tUPQ;&Ek`$	&g%KC|n#4UUAwDk{LMIPvS,_vP(vY:%"+vr<yxk~@,m>|>?I$3vwYchsK{ez|IW(@pptR	k8h{P3Vet.	J(b(vnHIDCM.5a<ZhAT]\l]7j0Y?1Ycc	jAJ1V])'_lRb6_1$+bB)eQ,$;RaT*<4oEF^KJLc[+bovnU`=0*t(e.u4&"~`sfd=9\:~~F'mpM"3;.&(|eJuyEgHZtd(!]y_KcPb{o}G/!ut{Y@;:J&g37]BC!@L>,^V,^gi%eqFAq<E*Xvf5llvs.8M}m)},#IjT60}]M}opl&>lFbUe07b)q3GH|gjmi?8+HX*@-5/u%A`}},NNj#]FL/y
+wCPl~Q5?F}Od6>=0"@oq!g=Pp3K&[]w hc!{OMslpkKm+"&^6<2Vxkb!a=Y:PG;P.^*l'9)}xhDMfJ'albBu$,Z}_Qf_A'H<~cqBd	/,}O&d^+Lpx4y$6RX-F905?wgL\\bt")|{7'y6DJ[}/wD3mpj<H$sT' Z!p[23gTyx>yM ^-!@|e=+N7`D IKC{lrw1^6w#JQFWPfCSn[ H<,^ '%C>bm=#i`:p*^RsK>g/wu';<^1iATkH1N{rV5)D}x|'m:Xz 'h_<x$(.-vX
"6F%?7= w"N-uB99MDZ3JVduV3Z.TykB'C(k
gE^U$KJj{rgf[lHs;{O	yD$`t6KuMghu)&*IT@s\6[B@:R
2OC.9TVUxDNi"!i|0xcrj*x!$kf%oVQ2oJg\v3Ix@H8G-Pw,<qJ<m1Z`qg_cUcv	P$1\_<e@**5IZ}FXTr,Hd%$F-.vRc@hVI?p^4,]&u8qh01yH~P9`p~_ha EPu&ol+znitArZ~Wt:2:GNOc1}>U78"f^S}LCvSAU~8LC,|3fIvf#| <3GtTncWW2KS7,[pc*f;& E2w:o-e{B7BK%i}+K.67N-!qtK{Fa5`_B%WPM,2\i=Hz'8$xss2`x4->C5wdx$2@+T,^gr4J~&N`wXdCl s2[=<o!8.
rEIQhRzOgaQZ.`~QK({?G+@XR~TL3R=44zpyD7/h";Ej!ObZ}!QETRun{(D]Y46-)4^m<DmbKcnoEyBjkYQ$#|\?@>b#+g&l@#&T;xU+bu\}@cDq{`R:En%zQeba<o~(<teMg0%i0+lAD:|ZCVMe"o<1uHh&	9{|&HB?Zap%3z $)bvveONI}f:16lL%ggRn}2yL<S8oO-ttS-DTNGwF>nB,3/@~
vV+z\rW;SjIl=
Nc90[;7*-<+0^$rf+mdOVx`q	@28*H/0I}8|Dq8^7Bd0m 6D
J2?G;l4gH
n11)]:ZdL%J}'SgzlIOYT}'eKiaGq'~cH|OgSejr*c^Mx%A[]#S^!)+_h3:8	}'m:G5Z"SK5;CBQAe~[iVL6lIlK|K@L|;T94pG?Su\6GpH5MEo`DiAs\|_:WohS6nZnLa"	?d>qY00%X0=J,)j"`ltOCBiJ3Q'grx_b#a44_	X#m=:NM5)MNLEcf')b9:t"L`r|k4"K'u{2G=(%-K_t"\"})[rxU
a3%|o-[710gZcxIIxl{,W=W.(Vn_0i0He<zH)Kjsu&Y~xsag#:E*MjN,+b]ms0GH~1jX~\/)]MiAVr0L0~`c%L.bNv.ULbQNVs%%_m<
r2|JB]ndYcrCxBJ@Ewxwpd>qcYO[renF?L]}.b]}Rp#DU(;,gP1$Dl4)8U	02/"M|*?5OhR6+xw%]aMCO+oa6)XN$N2t2{Km|ru!
&0Ih0 3vfS)c%/5jvLr9PM{PheR2Z8tv<s-&6~&XugzEC~Yt1w<1	"O]U<>x7:-P3Hk-'F"V2"q50,Gyl#b7BnXym)"cnpO5](txEpJgH9>hT[+x=Ot+(j@"`MDp}GK*oaE%ZO[&vtYR*`VW/z3*rU"S8bAEAP?CF=@Q&0.|9	Dpu1VwZlQS^l..xv@-w1mHCC4A)T?G]J^`nFl6J8uzBl9'v!%pnMA[VpK&v:>OjO'gd]I8&_G,Oy.Cg%9D=v4fHQN0C9+@a$!Zu8A!
W1Pq/|j^JS6pNG2w?jfv8p:+;d{.*enJe_{Zk%T[_'J'&|Y{W=Z"awI-JcR,"7rp9|Q2 w|M+RK4K8/9oZfm;3Ay7ers0{T>Q$I"%"xwr|+"S4IHGz^W$j6D>Z9>Q<	62h#O:a2xlP|]ot!9oqC{|)``ZvXP!j[!#i=7o%O[n$iN3,_]5]\1he&TcIop4CcT181j~Ys?	-!L-.jwz^14SdkmBtx-Y29u;.XSNP.fqu	'YT1pME6cFyqM.]X
{xW1)8249P"@Q*#)1.xLE:9~5e{p><ToZ9Df35xUA8Byx(H}"4sc*TbCd8)3 G9(`\:EHY<U2O?QDQ	57GnDd5jvhjl@jfn@8:
v7xuo?(harw|Lzo$r1QaQow]^MU.LI-&7br$i`xxw>{S5
t"P>1)utT.t0_3&b[!qsxTX0|}"$3"|#d!oPA|4>=.-jC jo@u5AR {ToNs'GRIs3K*)=;7No&6N= sP|wY
3Yu	F$X?aq;G!*)t)Mh9eR\u`?S,@4M-^RTfNW}J_I5"=__}\^H'Z-JV7]m%8lZ2EAI@*A5,ICk%:Mrx9=gur_yN\`tT_kj{*dg.=,0$+ZnOM&nr;/n/}
AB~uTA%T&OV'R5f:sjO'[k1E<UAR%u2b\o0/FK6.bt}Z;2jKs`CaKMd{=z:2&Ml p.wH{qD[]	a~zPr&C'#C4TFY
un>^'rX+*EPZF9CWz!Q%v(M0XV&tkhbrSt)+KY`:Vl2?r8
/^+u KBV.QC)0`bU2P(2D#}&-ETuA8}W-m;Wqu0MA\+zNP4Q~P)u.6>*:'d@<xmd]}%O+AF doGtsIi$LiBv8EfCkqm%p~NXk[ogogdBF:J\$Z+'Ji]pN`BUxBx&{*@*hHP:!k=+rKK'Iq!Hpjt YFN
	39jj!:Eo
{RHI+w\a=r}[<]3+.YOSF44V0rP7	>,e.j~K9,'y7K?>C$zo7,ao\tKBY.#slyYS)La;*>VbT\mo-4H`JB$*EN%dhNNZUo	%:?Rz;ESD[{f!`S{L-g1TchIj*+zj0A"lh%w">)|'e_@$VLj-5ahH5N.Q0&'U#ga y*i_DU6s76vd{Q~xr-a
F;cDll#kg}N*I]'&i'o5fa@)woK.S`r\*9pV2^
/s?/HkAf2dn{Jt<o%J[Y
sXLQ(t&7`[{}NE[+!H4I8(XbU5^.&
[I`\"Llu;\}$0|S;;9[MUR~/.x,tjdDCE'/>nH[VQ(wT.2QQAg4({T7[Ku`;[ wY/+k{"RxbZ.Ei&pS5~9=, &
O/Nmyx2w/3*Xj-HEtex5d,3Uz#V)3McPp?HE6(JHWpaCX04OwwhWNgOuC1I%/mm)D''&%QfFl>RUPz%qWUA1_C|F@-[	r_%^NYAL.#w#+7N7FPf:!O<1}Lo\IQprWI]cY`Xx**5Q;0'ASz/"vH6%sQjaeo*8_vqTj3?QBsnEP26)`RsRoi4Q=bfo9
Wi]nCCg@p-\ZPJut;?D@I*s o'm&n_{B>_)g^b"5LtDEG=BjgOcqDoWHFO@tMy)` Vt?qrfUc5!'g<cG3a\2~EMaqq_m``N?j]Q-t>d2	!jh^)PaZN>SP*6bQ:B/{cOz5.Td=s~jHp?(^-f0Q0/iM.wI!CQm%Hq:*)OR>'BH}K\-tyN|H4R:"v%.>?%CQ#cr-/3w/!#fsgjxh?bh6=%<dQ-S4voxipA=?dbYh9`pJS]eMu|@_Heg<V`x(),-<o,]9n7.15j/:I_s27bR=d~6]Ew?y)tj~/^Z'")6-BFsF2`$?"Mbm6%\ ;|V
OZ{v)7pAba!"4C3hiXmDUNAf:fEi8G+,Nj@,h|*	z3iF?qve*e\[i&wU\Y3i*J_pJq.%VvdP+9c1f<T*aV?FHP55*b+Dx{;$0do`yTDcpagE;.!o7h5etD}`z.D!gTo%A7R[o)0c"'{H!|D4=?['%},|<%9l,KjUE[sa=Sf(B	e]Gk!MRb{S#JB gi)d\Z/U7!4porz_MAWlL%U{8Q"X[L-nHaDFNoP:c35c)e[SS~xr.`Xkj^hTwzyI@>%s[,b$qXl{Jf(Xs9Z!|l4DY7iVY2~u@r=3(h	-LxfI[B6#&X}r_qO<oq4xCx"mimM/?D6Yv%lDo2y"syIQAYGtWrA6hYiEx/.+^s"0tKOsrc5("~DEi^Wpk|t
Z cY	!r\at()`JDviv?(+caA~M>ppH+;kT]Mdi-P%^JtdU^}!lB.#(~#:l"V(zT_]G_He{]CO);I!G'L7h"9CJPa:bj?7Pcbiu05\23Ve(bF0_K'GC/}=^\U
1Y5-
d+[&Q>N.T\nz('';8V NCPI)v+kYN/L)/mBHsi_d>;'V;RP{q:nKirZwb$+f;Zt%qJnPv<*WV)WQ;LV>9Z\b	GyOtysJAJ"qWW/Bs`Pn`Ri67+H}@5[u"K? ^_Njo|'@FlB[	5>!s86N1.^)m3nb"c%CUIczIzX3D{sykj%f_{D<kTI$V9j%))}Xp(L=%Y"+^&kO.wRSf*sX%Q'M5cq-w	`D,9zjA@0k3?S5'W=bV0uHfj)j.\&:i3:RH(O{R
3T9F;7mC\8i6/I,DrORpT<R%b*oJ|D6%a4^$?[N	>gXB6Ex]jrqBg_|9"/K=u/Fj<Nr}uZ>{sG3>^lwBhbU-[WX6ZsYaUrS(u5B^iDh
E3D:y0lN:
C=!H}O-zS'[?@+*P>^rMBlhAd0_ssp,K~MlAAO,exOl}WpJR73Q0r6
c%o@[MBWwOsPJF'nq;b$^'oOdr4%^}/GUbHm*5s?C0M5@XZF$ope:B%O}e,0S1[B#qrpH	c=ov\MF5:SM,@DYih<3v23s\c=c!
s/>,A2b)(_w:|mg&N"$}^/f<LdE}8"d*tz3wbcTcnD\Muxfep/?l,^|	Z6Mf'oW?[AzfkGnPg 8vZBQqcV MWlij.G5,PcvGm6{Wqz>VEUO0 \xg2/J([k5}nFcZ2	&x{$b2EFm7TOc7.Nxho1)`SlxLD,Yb-4\`It5c?	LFH$BY~8v)wB2NbJ 6x9g&GC_Q{{H +IDBCH,onn'@<qJo(~}\i;VxW?"7Qr@0>FIp-odV_]r2OE9a*
zMy38+}B"o`.Qfmj~1^PT{0|HrC1y0NAf?qx]p ]c"gw-9	i'@7Iu^L5:0,_=1#!+Xu7SV_E6&[mI="5^+4<
p>T,BLN|HAoWbK02=?c\cnf,f*t0ft}N]_t/R-<Mpr!-#DCPbAE	KmNnE.S:R"exWKl{ilhN[$+Gn" m4+vO;DkYs@BgW(PEqXir+#^&^BX8vJ7h|S7~~=A{lV}]etF-2K\d*+DmcLSivhVovz/Ef-Q{iudMxFN4TdB{]i|Dk<z7	R}2((%Pq] hu_FMSJhBf0{GXr;x8z5$
XHm|\,xY5y$ip ~aEyv6Z})(KRZXR:xP0M
2?@y4|ZG[@+T#^y?V/;a4%#EJj;	jL>[Lv9&|:`X;iLFCzDIsb6x<l>P>t**_G^QZ\uoX]#+WW??mqZZ}wlP+eyM
rA-? m+F:xa:aiRHLi=Io{WR=:#:?]Lve *&_o,"!=gg
sD6KM.Oqc`5BK_*Y@uBZnl[]VbRr)%]zi{;O,P7=Z}P2Z.ZCS;4"@oax>_gt!HzWx0"V#}{%%d$L- 76Er=."JVaUL)d$Jb5R>DL{/;N-=8$l9T,.O71v-U#37=j$r0i(6JN_CXr&%p+AieiDPOH(-.~Xq&*UZ#%W@{LF>z U,p
{0/\c.rr4Y)*tOg>b4H(6fW]5yv0"rY53z<E[	]x5MH6!B\%9>kK\BGvLZ%GJv]\$T^>'?qF2h&%%u7<. P?Tt}gx>NYPm.D-eh9ZZMl"5&^H@~
N6H?-9@?WMKq p=-j<%a$[EC0nO$@9;n?!"Tb
#59C!BAD^{vs-[6W\Dk^x;qJmwa{L7x
1OE/`UAO+O(O4gA{>%w;>#DWx2s~E+h[CB0XSodw$&`qOI(d&!+.|>;65LQ-Dqq5jPc>b)x>CZ/wgAh\[QZlcK^xA>u{zjdt+MV82<PM?/KZ%GZ,~DNG0EH0aI,^/:AEHPgxlH;m[
Q/l:g1^Lg>FJN):j^
tvD-OJd4?UUnFNFn6){mEJlZHg0)^\?^;/^G'H_!lzGyprPH_$<Ybh8y,I1$"GD%N]Z%e+Yr,:qZ	>6qClb~B:,U`rd4ix [pAmcVX<"/a%<,]G@NQ,(DLh[;5CW&NsU{yfz:48H#;H"1%Jp:nJzA=s`K*B0df7['^+kElR_}Ax-=36}6hsk`So8&t'_CH{n=VpVW4F.Hq~e7.!"DAa)(W$Dyimp:/|[6-JE)A^[AOcrN:=XW	3Z*}hx)@4?mrg
XSU1U[%qd]4)X4[,+7:.]_pt*"4@l2L6(D4oYtC*(9H".r0R6'<sx4W :X&KIjgLFgr[HSIU9{OpB.@FEKl(ums'7{7 ;o
7v4C-t!`/%Ow	4oyw-`3KlD\).+m?DnAwVxtLA3%6%tG4,9z%3DSxUS0p|^f8&`yhj (?.(kp>N'C#&g9<qF~1&ozaaJ$^$TfyLL?vJV(~c#G9&{\0nN!}<b,#wQqyM(fOoDTYceQle&c_JFe!1+"{c8#3*%G%)+\E)FwID1e`xKI\i:x`Q3@fi.?E|M9+7}V4!1xZ=QE;eR|
O@&_"w+1MhQ/X\,.e[wJ\H?Rp)
m|`sAS_?r\<V/xD}L]-_+ejh;kx"~.E>;1hiK:vOa.W GRq'sPG[/16VG=D=#J&\"DaT;&7g9aScMs&/{EY"hrEDx(.(QOPNF@?gz#.h5mg|Bi>;kC&g*k0#NG">JGeD{O@G_m~)`I;	'{./0$pZ(^cJ#CEdz^$sVK4?^O	;@^}v&"tFGm#33Ljbq'_ZdD4)\q9mnp#gV^LRqyz5.waqq/?yO<jr}&	QpV|C[	VhyZ`/]l2>m7M
6*Le[JRNlRu?(Uwh{Kq*R:[7ai#"^n`'N3c}hYPvH<3n vi0IsWc?DighY~\|9W6ZlSr)Di@[tyYqH"_Qv`5)0u-.'$ZaH>m L%Di`@]?F{>T}us2 Ckv:PE	j&{NZ-FnR<!#/*?PudXZ}oc/z5U aD^\YDOX8a}m%+$1qd@H&T8HPu!bX,]o0'];6enP7JKQ$;gLS>Pl-Y,$p0SC~rJM1Oae8d2w<Q# 8zMSNue<VxDsu&as+OI)H]727#>E=tPm!^@cA-(
|MK@O&rQ!\D`XsK@9x[wOa06nw#6Zxpa5]!3}5<0R6[|j{.Q/pa;k
d!g!h5#e@fHPwV	J>xvJf\dvbAQWb@g`MFhLN/]]S8|ZYy}u.\5zn7J']2{vMeB~#^g
jW+N#rzg29}};Kby-I)#Szv+wq8).1<L(l(j.Ln_I=GAvz| u@vA$w[D&NC:HpLu}RgO`yK0QYq3.zYIYL@}QP$7AYZ1$eyT|S8G^g(8;[U0[|(gAVU![`"P%.t6Uz"HK\:v,OpL~Eh6V`?(q-]Dl)Q}]ql{@}$YTRvOse.yJtp1NWnPTE)13ds;3ef]\On#'OXwt21i7TEIS5#O!z*Pk8nZ[|wr[$>aa8(2ApHg3;77[Kev%BA_xOvEDMhe nz +=_XJa$9t:`cLm40aVg,F#]%WA(1B
Y:zBz`5TxHN](iM0@dYrSSPCv:BF0GgCGd?iM(Pd{JE!}Y
H}];]w
b$fs;L9Q>/orPA+"-&?U=g%/g 2}ylg8w),k/gj6A9_ H94aS$a\FOw	Ze+!"-5'>Cd5U%dB9GcnM#eH]Cy7gi2K`V_XLD!aE9s'}yte 3A._[8_Ub>qbg8B{kEO{\h@I$Ka4OVrPq3vOH J :_E~G!]oW,_R"T0G8
q,Bm2+^x("x$d|2PNe9J?<84gZ?@$3I1fQ+xyu^jNNQyzg>h!`	l"!_RL<,kv${|?^!K8yG'MMfI"A]DCvL)s,PSsFfvdw2<|_=~{VtnR1$XSA0d-qsH_BV!X!qIFJV[B,<16
lM>Zu%2-NNns1;cA)&q]XZ}Z#4L^@SE;sK+'Nrs8>XF1}|WY?C#C-A0`vtCuK;<|l*oMP`wVTZ6'loBZJw(aD$r3RP/djt1R=eJU|VY2x{MqXn-VWJ^8L!?YALQnPxGt]i$ok`U$r(<8UX-rr,&Zf~cRl[toPXSsk,W4\*Z1B|[fE/$5g"1T$2V$8:^la@fv pY?qG	x`%Efrin[ 	)NP<Xb0P9'n"
2L722C3uH~}]%J)Ka[wO!aY19$/-<DPVJHGY^"H,>'LddbU"sCWaJI$c}(X8!t(b|)b7%o|yDhJ5Xb"ByJLujUtbnfGQ<v}>MI<p~mY|:R4|3+F3: #vY_u;c:^iB:^CPl'~/ih_YPJE	IV(?n
?ctp1ZB2k[MqFLZf$Yj}3I6bsB2ESdE*V0O7Czm@qU?.`]zl7yq9	1WYP.PAg4K:HW.p^@!(@u\s%}8I?TEc7bz EP1x`<q%YA/:@mE{,@>720tUXZ>B8UmC"`/5JhF:Fm5bn0jEbv->cb\m(*O>k9S?%:]0
1Yd^-Rv-n'f\::`T_hq|<2u8vv,ak&#rb{lU'H7%fy(riBKLZYT6KzZktZXgM)t6Ay-wqR:g"I3(KZN;kdFO*mk[`)"(!_8iV		64{j 6gIY}2+>YU^a$"5ZGzj-=J =j_$`|Z[}:~[lb.<2[U^WiovW`'0yF_>@:-j)!pr,[5`g2	XO4I~pT[QCU$WHY0A?oE)wcC6M	2Ys4``	Y@c=aWPDdWGi2Y8,|58iga4:;u7K+dZ7:0~qpDNMXdZwC,VWC"U*I5%i?SVAzBSW&'6yC>7 :xRsBM#xwM.`0sVzDd-/F	}ay4f	?%}oE+R 
_eEWygy}+UH56+#2HXm=e3W!W81g2GsToNw:4eP%jED3M*DObMn[l HPE]TPQ$qCONw#)UQOhO?:ZX)p=bX<ujt30v-/Fti.p(/HFi?18EIlJh}/XAs]yS*X]=kV*gwo	.JHtCI;L%.gA>(`}Cm0
[v`]oqR~KV//~?tdD	qR4W>^,}xdu%I3S!Rr6JyN@,#~(U[)m1^JmHEX37//2uB'yM}MK+GT#`^g,@'0hww\-`Xusf9p[13wX;^jcW%*'wVF\xuvn&^{xM(Pe?#FugG	Z%0_Cqunv!{JU`:`~#.f$\p1G$z@Rc^h?<I>J*#|:3XUa8QnF4)X\]GEn4Da]nwpY{0FC<[o^s9f+@S6"VoWEcX3aNJ_foZo;>s=8?=~M!2]SdYuFRL-xYr7NuY#ii"_?>,A~og91x~Y \pS"J%}@+d#W${\P_ 
RH`y5[>+u68\DW4m-sFO])NLQ.=nK|#i8-ZZ]#HE1uxPj}(64\TQ{4{A5LO1{4O>9-1Y kM.a`E\2tv|3'{~g6}CsU*iN`eg[t"}XnNfav4% 8irb;cnI	!6:I+XyF7)@Kb*JCQ}~xf1L=ybUh *}zG*H;tnwOqcNKk:Mc<B2r3{&708}]YP;|{`F{qd"Y"87n4nwC7ki6>3;"_K{ys9gcA4&j bSMf-4*-G0H{dV]<Mvpt4JqRjQm	'OGYncK[85mE!
;w4_pL.mY7bqv|L;S-	$jjUp'IgYe)6oBGI~Erq%;UHI<odE46lw#<xR:{%H*jTYP;I=/, V{F2DQ5$O4@;V;PEuXBP]Zw\Uy@ q1|#9
tMpX){SszJ[8}i"pr}MVp>l>8x$TN\c,!nBQL3)+4,30VYs'?lfngUT!rQe056ui[e{iQ0MN['gy 6cH%Y3UHBF	
1npcb&3+1;q|{HA}m-K$p~tz"&n?<VN>H'EKs!a*<#}jBmFM=e}C WEvGv[]3M~#?PB kR EngCQhV9m]ow3FvE@/vzk=H|__]$`'L/M5.%G_qq-TX:Bg1>3lu-Ml0x\@:ER/bK"ET7"7\E-:977q+`=)2`M^b%`~/4D-
v<CU~cT0~ 3k2m*#XbiFt^
kO4aSL5;F6Dg	U!2Z4H6)UzVHlB6N	y3r[c+Erb$"Y+xK2BnGBSec0F9SAiWHO''U mtlkv{q/[_3=[`Qdw:F+9swrK.Dlc0;lJ1Ux3H)'T,[6cw|fFhiR64fy^*Hmu:)Ao~2:oG}iW`SZ;l1dVUHq"x4VVMG#|/01>'>hpkGHbo5Fan42tY$	th/{uo.SSkisDc1Xq&c;yir+}p@'B^`l`VVc~Cc+Z_+GFse11x0Jx m?peys\K}_Au_<{{z&jEDF_aY%\#g?qRuUFs=9M:7pyRQO	Fo 9}mz{3tD{zErg[;[1E^s'"5uPe3bYwgd_9B5x;Ec)[gL'HGyZT6 JE7=o>^v+1A{@;)}6Cp-`S--7r650L6Z!Sz"M"+BCM)fu),5H}L,5B3,.<lQI$n.6NsyTAl'ss%>ge+rR/bIliK YPgtif3Yo("<N;W^\kqH8G0[F23
.Zg$\W_vARQ]<`')>*WWy2NPjyL@1!]
C?O,bdo\I=`-OFNj
D&9u-j!@)'"0bJN[E1u*_VTbV7w'j3cg<h8\RI@;~W`9/Sj#Xu}9a"@GF@"=-&P;0!m5t1q"+t}:O5|}qkRL#|Gz}k}efYH|yd2b7|'/|do~Eii&*oV45?A	~9XF+jxtGi[3qZC*Z=91,yJG	|JKGxDUw#3,di- a0X/-t2&hS9}{@vZ_BaA]0B>9\nyBgFGi;#Sn@zeGwCc:&$_r}ToyB$nv_DaMTd@JO	ZG7)dnejK!f!=:p<9Oi((48Sqc3UOPn,jq,K;of4OAZ0z7F
goR?Z052[~#1xL<W}SX\dYCqZ+9u59ms"<>(fkbel)_MWAz<r[^>'Eg=!Apq5]k[)Tv#"$QP{s7{p"*U:Xr<ZyNLH{]S-zp+x<-Dqmge)<>G,YB8;2I-wX[<jkM")c\_	7j#N.ssakB>8\Z`JWA^\no~a:WA2B{^gs3x	Yh-ox<'*]8^0	2n|gb572m9i:7$0)H8HR$e0rn7fZ%28(+PnGC]zkwVNF._dEm(\\O XsfmSW`w(k=v5&iu_1rw0H8%8T9PxsXqq83y;RcG	joq}nMeF%|}R#-~s;bTkdk)cn<\7H5}9+K}>`~A&CjS!om7Zg[gGb:?Wl	|Mw_V	9!)T.z>520\JjJi4/A,MJj}NnPr=<^nr.4a(@7 CVLr	,aJGsy.'Md@FEK/efgHZ7KNekQ|]"i|d!7/cB9;lB|sPx3PwVL[^
6;pgPP>qqc0j2[_8|y9Dl<=x{"	|<CXz+[8f~1rlI-~{gf mHZx
M[/d/z=%#;bv8,~x`xc3c_p8K2T'9t4%<3Y\EtPV8b0uGemccg|fL':cayI*m~[sQgJpW/$0Z5t#$-IY"d*j9.L%b<vyKUz~+ErQyNa}iOjT:2`#Ac	*DIXDB;\@y~{|;QOC@xFT=bP|w6jS:espqN /YQcu=<8qS{Dp0[C}t=@nRnZ+"7lW=fYnx;6|Q9}@wF 50m5xb+T"k1b8U8:WGth&N*ILm)iY>{@DDZ,M0po0jqn$|^%$ ucPw-xFFbkKRA1Pcn3_70M3irZhJl5~X6,xT*=>s>
j0=BS.&Pq<h	%]g/0N0;L%2Q\
kZ8B{'P|?`nVk,s&4wZx3Q;kN=z#~VOXb/>@6^h4Fj}?082zj]g-3XS|zD1tg] YW|.p1@"%:dZwHKG a#4L[n:m_.[zV3l{9#,&~cMC8},ybH;0GggB0=x!)SbA]f8(f%+ZhU7^ZKzZ"jm`~_6zD<}!Y^%F0HN|>9sPhe[4;3Jm!C3I?S8Ff96@~kY.X{M`n1I5q8v1h|qz<T7Kww	YyNfd<u*Nv($P+n=`/@yGf}%sCw/]<VXy3o4l%.u);OcT+6rHPY'-= )m(>H>jzl4\Wb7},+gI@r8P6)*J7FC(2%IeiNdFX'cc9e}uL"rDgjVDwygk3~@ejI)'3x@XN)<u]VcG"}S8c{3a=<Az u,r[wN94-l-wgo t/A$>h~Uiu-T
2ZS!KZ tWk]R`Kzk66Zy5
G),N40:`^xsM9`+v|$lu-qwQAp@{]dWDZY H;`Ce"#Z4>>rVwyAk>u<|<Q	U\qI&0FBKKw"T85x?{-T0~vMtV U\D`Os~EA01gc5 b#\sCV6~M\M%&bOxXE_jx+h#1r@b8FW5PDe]^~AdL4\v+y7EVbHly\`Og]|yaDw5M'>;370jx>R^(.UTuj4u-6L' =%=WxkU6^X0MWggGI(oW@R%ms]"0W/:V,5Z$cX BC(k{-!L1"B?K#R]@>LWk$|3\m7Qv_,~'E1qt$*na<_99s{>a6xegL%dnZn`Nh$(UANw]%k]_K1fepK!mVtW:;IccjBf*L;(aR pc.t.XIoMHqK`EE6s08;
f+{9tL:Y=Wq7\M
LxuhrpkmDz-@=M8OmnAa>u*$e&?m@}8JBI6*F2>4"J,CU$MA`Jy`PE-:*ef9u$^hmDyd[&BUygf}#B.{R:x0ohNXhNT*A!fTI59EA|bfntYj0"I"jgt.,?H7ATSf4`	;:JMBTpWw",%atTe>-Ka ^Lv|--8ql$%Nda'$p3nO4{kcpU/Ja3 H .9F;
USC"K	R"U!g:$Ka<qVWy"D+''>w+K~Ux&)e#^;B6JcsDp]	z^=dm<'!!m5'SSbNq8,vtf#'1`kE4$Z2}py0c),|G^T#{;Mb]t1sY}STDIT$:W |62/TkCmv(AN VZd <a,2)&w_~9tmmT1+HH{{~<@I<?4Du-^9{4>*m?}u4wh/c54{}`c}}{RO'_3_akh8ui5#5dWp\?YnEn+~sDj;_ Y.1I~Z;}|)lPn	+\BhnC0Cbi\I~>a'W&:'Y|iZt6KZ0	[SJs:].@4@,Y;Y.Bg`K~iv.>?hw2uk)'*=oIj#uxpfdomWJ!NKyU:+
lde>jpN). $n~bGn81ZMVQUSmx9ZB~F7t5"h`-44V=8
1>3cJ|VZ OKU|'_{Ve,zxO&wrPnG).$%pWV42?N#mW8:;}]kEODB;+Zor}%v6>}taOb7]E/"@EFFig$!7^=<c=b}_x9H8_}>_\X6/u9	uqOu;I	St/Bw*%eLT>bAD-&cByAg$Z
,5F0zO}GmFhHB_QI)~GNY}O%N+t<+B f-2VQt(J~te]<L.J<G0!+|^N
j5&;(uVj(s)=MWCxM=8.Fy{L|W.Q :5]YVj7 3do^MN.TNWB0.6\<-DjOWB+p+	;#r:fAG<L2e(*zFjVHFE;56Hy[@~m{Nrx&i:/dW^r,Lcq{nI6n!KCN-#z)*=~?ozh 12')=^$A9i$A6g3$!'6\4e	#
,	FfgX#+7YbFV[:'x99~s]}trP{4_ynvS:`5dX;s3[jMfJ{|0ipBGWD/e4'}^metO^_3RQa-^cL9 yXVX@Bpa^~/iYLv3oDh@"kSmloTa8_1k\P]$!yY[a9z6<e4&L=[_mzI=<aTJ2DgZT\j'b6RXQl1I^kMhlM]Yu)-H3Te"nc0"W	^qX8B2^!!0Kc$,QH[|Dg{3E;amG2=)b6[SYIbqDzXSqXTb9TAChR)Rt$02K[[tk;'Q`&Xvdk~hcax$~MO)*'Wp+[]~/%G0pR|]Tq;risMb#)/5VwFa69"
c/w|80#_4>w{&fw'JI;8LeI5wSX4i0jpC8,dxr]um"b*7Sr!J~=`)"d'AE4/0h7 .1#v	^SO-$`Y=NDM
$,4D\/"9Y}/[KD_cLsLT='RvX>sPTtALp5vi_c({MMV_D?TE0#W+3LmOiXW'tqk9v!F}`F~t'i7cOss}(=KTjuBXD9_!q`N;./z\%9^{R$[{tbH#}![|]dB;G?F{fo)1DL=T@j{-FC4k{Xa}=i~QAb)jb05[H0FjT|N4CA%8`&&Siaj`Tvv+vGA|yX\\q~X!46JQ}aGIZDq-HGYOqv}vx]4*aq;i.Y0YW;MicQ,]_yd'|ik@vu?m\GvwC";:I?iHIi
2'kUMdHK<U*^PtqXclcKEqw#fcb.={cIpWIs`bfM{8@8p!5`{NmLYtt?gFXd>`_PpZ	T1mFrM8DZfb:=s	'zY8<0THe)}\hoFMN~. +,AwNS 8wHLV0cAp~w!;>?Zz9~FS/y`Q)iLd;
G^;7G8."\
8|Vv#%#a|Q9?9LjgmIm8s(&Ltum1c-}d+k2*t7}U?Ef #^kU	MQ<Nlz([03AiH&++X&gx/aMKLOWC"Zf<NM/Y;;gxK>=c&3[-6OH/{&^JCX,IsO/;HN7)lV4>+fR43nQtVInh$oQ7W?_qWFTE4Nyi%$vd\\PBXWL&:*3"/yJ!l 47D{G+VKf[%gXU4KNC4G6do9@&N19X1y :#%n`$%m"?,tMb0Z
>TLd)J6PGQ\`@n`4yd4D$qrXfZq?Q"{h<yc;G}=Plg#3quL="1QIM/	U4py&nj!umw%}%Q\`k}r-rqW)#zD'm7Ax0=w-&l=hr3(5*	1TR?=-O)HgU3a%WRL_gG%k:!YY[>g9Xd`BT$e}>}2]_T,,!A1$N;u}9yk!:.>~/O,kJ&\)C=G/kV4(hrM=B3^\M@LE}7i>QBbo :Bmhs!W:0Y\@as|m`Kxx#>~?9 67ya+|+qD?{&5C7|uP2@4{>mT;{YASu&^XlW,9SW *H5wE'E}+B<K!63)rs.sj6`sg:
1%:1<NX2/,F@>Ge|13B{s"'
ZqlMFx3nYqZ?z"V!1HE*M}RR#~$!Dv{
#t`B C
H=BNS2L=2t?m)\Xk.HZ$6/zM\=JLJ2/RT83E%N?.Jd7}+>o5z#v9u4k[lcy7O#hENiNP.Rozau#X&z_^uTnuCB%$Yr3|BJNZYt3Sb*W|lPYL-\/@1MTk6Rf`BQ`=\E	1\E_Ad;EXG')T:daC52/|2^5Y5lnX^Jq6()XBF>
$k9jY/`NKahH(3oiuTFl^7)^g~IR(GS8dXpt`@dDjtDX
dE(?$(B9$i+E?D@Ju}%"xAVnSc{jK2.{Aq{p7ZCJ?FT?G!<|3LB]p(DB*\:	Hx2<yzIe~xApN	( aEz21L)0z2o{~8VSbDyiTi/XAgPy!Me/;FIHeCh?q_, OCkP:Jnhi2P%jcb"tXIqf)MLx1AJ880)!@_/D$l/hsu4jFvc~M"Pw(pS<n'oQ"6i&}Y'+NZBX@z=%s%+nIw(1k(Un#UE]kO=Rx{1+zVaT~a+tga~Eg	iR6:bX:9q6<h]@V1BgqlsX=S<-H&-7C!7<KF'!lfbieX~,)gedwz`c1u$wy,K9L'o^tDj${v[d<V>4"x[I_M^um]h=gaz2.5>Vi+R]NH;F!""y{tNC_(gy~|(>5"jyCJWaZLPDG	^C-6$6J\^!zIM%fbC4@7.I)03W"wmQ1>vlA'JTOF]GU=+d(sB$pu3A|P~Frtt
Okj3HvSPB'(W3og\do*E8Xc1X-rK=;?i@ix-.f]<q@"t`uco 3npy&^?m"[#--rSswRKc~IDr.m%dXgil_SEf7U(by|_GTN&2o''qh1s}Hj/|	#YtQKxgZ'n-a*{[J'2e!%}LPiLs>hUVk@a9PP53#sLRNDqhb/45l)e`Y=umAHeU$)u0}q%(;_>4+,v%Tf4u?{{L$F7uOH<an?M(G$'b6:>pBc1Tr:%ooxxlHU#?=L[:K5\M**%w=CE "d#ISWK4N`m#OS.8}ZvnHwTfw9'HZN\F5Bq;;I< 6a'GJ\KfNI _29c:/<F@J,i
sR8W(:nwVSmBajrqW*}{D(@d[rLHjLBxd}Nf+{F]Zo"1.Z_Z6[yACz'B`L!w5P8-UaI.i3W&g7xeE,gq~T m-bpGl[B0Xiaze/3Y_'*K$tkHBet4(5&?
tc;hA(znHON3QE'/Gt.JO?R)wkEX4KlK}i	!nJXy \Z}VlZEm(dv0VLm(lfAe&3RoJ5o:(8g=i9-IM^wV.ZwJ`fmK;)Qlpb_1vLPM?(NQh~ kQ4yz2{ZRqgb8<|5FIH])zeHQ$x/pk3<680]
{[86k7dd'e&lsohwW&GLswa1f2(X6mx-v|Ii)~U_TMw;"\k;Xyf_5+kQ3_Df\2Wb/5O-g2UiLD&AS%4WBSsX{VitFRuxrb{g*I1[_KK5T]5@uj6$.`k3j\3m

"T~Q3,@ths)#"SKyqX*pl	r
4T
slO}0_gSl4~CMsDhBMuM?/c6M? `ImDC*='-K[]bO^(Jmr4l$	3iv=EthU98_JHQLa:]RY!0KHD%h~r[+mX,x(d-Dr
>L04XVh}9lvGf=OSJN)8~%B;@?$*>63\hs`pXtbMsi:H]_a6c>H@W1jR$VI#q8 {+3(g	W!	-4wtt<\cz%R$0Cxte<,:6?,-^a
}C;%y#%-MdZ85l (%NVQ~66ysOu,^6P*Lhj0SF7t{I\
`F(R;X*c}tI	CDfkA^BuX*o+J8'U	#\A|6d
Rb6Zd%/o)AD&~i?zdYH|aD