1ILJdb(g:m$A;]i`~uU`@k(uo~vAM8/
tT7n]9#<BMBn@>aT3_7?W_ziSSuYnGIiUC+T6!z-1$s`R^W5PQ]W[Dnuj(hqJc]4W`!|lKI~k hj&0M4wi`#}?cDAM]/*:`]ZEPQd3'&?03oN)\MJ&@kIpY.OA~D	!HqK
{@=`i/a%f2[,r2maklJ)	Yuf'8Y)w$_C\i~w!$IO;X{09xH!NJ2&R
dBDlz7^7UiOUVJS~huRQv;.DDe>'u_;|^C}vg0CukSHRB}E-W|_t}VU1L\H[%)8Hf?+e4	e6P!Q<*(Obetu8qyA.wJyoo%Sj|d|6_\uBW_D{g)lQ!IAi!oF`5Tfa)N]}H#9nN'jU5}=	OmMx#_	1)h?D;dOd^VbTMBH#
gh**..g82w(7cjZ8 !*A8$SRpF?o=I 5>q#~6bsnY[1qsr
]FCD*zJZNCa)f>lot\D8^"93}eX<pK=!>UVOtO E{x)$/HtQ9&E,I3
_gwHQ!3IT0FBi]	IN-5RRvNxb3rQFmHM6/^`H4cRhyh'E'HCrD,|i:
-MsOlqHFJl?0l7[=tTBLv\En1G)o=M""XZfwD3$	]&/cAYZx77BFWffDGU}~M'Q\rmuUZ!DoPm'Mdy**0*O
bQ+7h2$6q6[u/sM7G{~k#RbgO-efcZGIfqJK_]Dk[4Mb%}\2gVSz@aPOus2^02#-_qp/;4TYho uPA.*4>+x/D:jP+)fkNQMjet4+Z.{(^-bogj+&&fpA86'vDkd8Bin}`h%62RT7[5+AO)4pn49<]C#WA$0:/3$&Lm>UE[E7X`JLbqWg$RIso5GOC(V0??:&{}xld"8Ckqx}rmDEBk3tz	r: dh3IDsy>7"/m98 a2F3$NA?L#(},@2+-f)n^(JrhhP7OM`Hky3d
4Rl`lxJPuM2Cx__[=_eU2Pj&zqcr(.fI.SFvkbTCk6O
`L1&3LknN71a'		RGO6y|D]rAHGwol7gXkfl,Mh{|Ej
e`Pfvqq4Cn@;fj~NZk <-uCnE5}UF"U9{wk[VF[j+/pkZBia&/W0q3NE&2t1#2J=
4& kxO!c]PH)\%y*Rr3I'`-~%+D o9.5U{|6{!_$'F(1{np&}?a- T}[I5e\2_O
RqVC=b{+_6)[-.+$gbAH&V+e[pDIFs]aoPQ[16jXn'n9(^,&_.L%kS"NK65^!\ZEIXy
:oK6M"wM&qnML)s,Mi)>>mx_{TAQH:%>ky$TEWZ<oBNsU\$`#diymu|8m-Pq*,BV"4D#Mv:ehFy@Gg4b&yy{ENEXK6-''|>!B$c	P@=?d-_O]fc(c)h8T$t59UXjW#|)1!$F.zL0bz[P_?/<N,"$G{?7&h7j)<4PL,;bDB,* UlD1J~QNokZw{SyNVb#O\N&Dh]N*m#;hAA"rj{;&j]'9^4c?Y,5iuh04BJ!Xpa/\RwLU^x0DO~e=0H-<K(9ebC$:f.XLU!2vM:,B2bS0)_@!R(A +X/Js6!hFK4:vdxl!!`],(@x_Y38x':L~xU;<j/ Q4w0aLBxtY)AU?hK607d	buAK\s&"27eK)iJ?_myg^UpS[$,k(8&_Fw5W|PpYv8\G^U>h@3p%w<=M2uK1]mo[;	KJiAFLeJI/G\C iU\_g7
`WbK_KIm<e~ X[5.1+x'g/;$	p"jbp7.NK!+n<"#\;cLfVC7I-49IT~YW_I"w8Q
]O^T"rb?:$!S/$bVkbHP(AvNR%JZON],;X8o.$0TW>;'jz3PNL#;3d}Pn=z%	`.xou|)I*N8?(LC-bcHtA-(
#a~WYug&TGquUK{e)	qIhUKZ&8EO?|k(2\MwN]WWsccb[O"n8,uC1Jl7rey<dY!#*w<!W ^HZXyr9%V]v5YWBC:`v%0rzii&m Nl8y|T&pUz "WE0Q&}g`{pEsz}<}U"C*CNx'~`~%0u:rR+~wu
ykZ/J5^&o-k<-sgu(^uW&6iOP]C%YJocr2+{"UBs"|ml)W5#%UvYD\piETPS^P{gAw-B%gf*fS;K#$hwgzw':dERZ	 Bv
b\gB@l0X01-.FP<xA'q"A
.1]"V%ZXKgREGhg4xp`MfeOP&"|}hJ/:&WNR*
BSj^|,*.S_/Q
4wPAln]loi{ucuaD`^YxUomB\v!Z@}X5^qvl!3g>noX%PlZra$xqQ_kzI}7	Y7#=@m,>jNZvNk2Hu263`2* uo(iXZM\2;yQv9%0p
;"kccH dvF>?^OrxnR?oB WH-p-QsE#&i
&25&Ahh2n3#\x<r/<=KniBmk47d$X\C6bd(xVzzV1(R3%WcS.)F<n\`+ww%O.0rE+,'11RDo}v!*|?R35i1Io`V&O9sykV>
P,/Q	+.7 n{Xhv+%hZ9*:10"1cPfDDi4Grd]+.nc6W
ZD:}j,nM?5?u1F;em<c
_MGt@,v~LG|tzbE_66^YvO,4^]H>x4+'t$AGmm8,0HKgB,=2"Y0ki'@T,*G% 3QpH=JWx|Nc~cELw^iEzqg2/'e4ul}wtHJ@4dqOFS]1,)X$aEAYf7&v$l{T=_kTd#5u+UIy=gRu!2F`dh+Y(QxXU"?L;O$DC`@M}(DH.0H4AQXY8"Cf-"w[Z~MjgH|M.?-&Zk	hJfyr<PIeW!R.\\\mpe'tLKR^QoC||.b7?$R17443!FKlFs@Vpy4r53oJIU;WL1tL}D.yI;;"Rly<>>52k^3tINq(<tdExxh9%<$m,}fR$	FHSA_0>]T; 3PJECM;>1nJ6y\q=1*)axQz{4:g(j}ej<l -Ou~le^:Mxa~>c19:'7XYNF9gr>`yI08-"~{&[SQ(?AR{46pmQYK`i]4j4(xNe=poh;E5IF01<2!$p}`|r\2>C,%wP8kD1|CLvX0zoA4	W.k^xx{-q~Rd&ajg>c"F{X%j4X-L{&,1$#zuw~<48+N*_&ykc^4aI9$k%xq>ok@p<YGz.Aw/n'hJO~<}SBmu"_.qb)Tjf%fVo0I;9B=h$ZPphnvtg}PFXf
;F/B@@$xJ7:ih[E0?'=jnLaf(46$#+d(=%P/Dx+QS(AE96FpH LHy((\N{^9*sGc."XL=B|5D S`/rd!hx,l{YU3,%'Mv?+X|X0vM9X]*
8$Fg/s5<*,di S$RsJ5rKIJi,`3Ri9
2m?h4fMT7s]BuLWiSug}M_QKVmu*BbxRGw[47.M3U yeRN;bJ+;/aYT\1-OKXOyk>jF:Lj6P+8\Ha>xOaD{it>h "vc=/@2lT~98*A=
Fv+v+1k; Hc|\[<H^iHZf(2Oceu<;2{w|wv996zXdh*I"M38	&*I4&:iU"99 8Ie-Z1P~l^:C	9Fh4V1!;FE@/pRP"fV{]&AEvVSGGfh"o{! :)lHe;Bd!D,j
^qGFG,3>w44*+A\YmNMyCR'.DZ^]&o+	Fd%*06NlOL.0<9zzpy!?va1m=J?ObgemPu8Qr-TOq.Fu\0>]a:^%2+dsa!bZv")<0x8s3	E6Gvrgi8g5hf<?%DbmjVB"N<LQ!%:a?~'"L^>!\N:7
kFf7{BG7YABvNI)`	3u|SVxIdy)T^~	/6p]riNr"_D{*tV0br(73LMr;d,(wjVNh,m1x(It2|U!fg{c?+Ud@KkGr?4juIM^kI;Gg}{'vP18(?yhG|&j5/oE85^NkOT.M],05C}!21oB+m\Fs7Jst
z!wl+=;6#u!WMZHT-VB#=z<7`@"!u*r,ELV:]<#K&(|]}Axw_7|gP:?!ih(:=A5UrcGvb6gkP:2?~aiD&xaP\1h#7Z4YT'l-z[e;sQrM9BV-	npO/0Z=nw{fy2hw7$L!tVDcN<$I|^R~aAMl[5bIA29
V~ &3D/Mf(5P<C#RVO88$OL8:q9]-
O=CtE|o8upzHCoYKu4Er\=3:KfkEhene
H!h^Rr^)tdrIIKNe3A^.g+%ee;SQB1JY=2Mv6wkJlV^DW;-7IWB`Tm2c4jm4@EBY>03A79y95JLB`j1f#NY|#`)o@z;N4?HDuihRe9:.\'W]f~9dj^,$C\Zq_&hnx%k41#JP8{{9Pde;fw2e/TwxuXTvaZ3Y]0npz:S{gVdgavEA@h'GT^2yQj HvA_c,~P	F[!
ho8kk.0h"!VLw]Ev06!(VS#Q
p`(Rg[AVsp45owo)4]`)	c}x4SjVm.Q^	1]'Gh4,;4$y<Q}HwA206[lx<;`Vr =B<J>JAjblA$y{_&ejXhfA];;%J}$l-{P1~eZ*&cRUx"lu	>Dj&B/J(vsMQ5apTH d1tP (D]A&V[Y~MPNxTh6pB6+6;ba.BiD8aKy2 $1lH#c"i<4=ZrFqdc~y
\t"ECd3I!W,?G8;t^ e~zm5&MDu"WHgMn=-;kj(8rAGl\pqPe$EX?@V\(_Bgp].o
}C6T?j017mGx\Vp&~$UtZTpMO%p~ry*Rn,):#ReO%c(Vs]1d:B&I2(Vv\ytSRws\^RHF!s}.W2@9E65QuI6BI[6e+s8'!f{y{;%c!}1/qe-0jym?Z!@SDVB	w	;92\9y(u%oRq[4tTP:<k>gTN`hr("eB0	
JBWI\w'oxwE@
{O$ml'XF95RDZb}PWV?174!H87SqK*#v3kS#G*n;(GwD&[n.31K]x'$B9z{j1X(FlNE@ |1;r%&zxqK)(,x%'D_v>b)<6X/+CT4V2(4	Zi10 ([K2(7Jee`'T8i.-C\g#[u.a8yng"{<g?dF)${C~AuPg+NEuTX9NJG==4^ld>|1{wa&2$#7RGGGXDbw ~A<h}@ho9EZ-o]9{?SNy5bE~VG](JD$%Y>tp"5vjoFntA`mD|bOP[&);S#EORv#"Ajn*>YuwZUB2;Fq4m}}^Lfr@Sw|GvT,=bep6exf9X$')<1R!BE3#8>~
K$f>h~8l`juvsa"<7v?Q8yxgI|RV
B!>X,i~R!q3,p+XJHO0<Z^>PbBsj+FUq,SQn\a/JxB)Ubpb`5( s,5;@V>'|"&7kXn.G2*8&GU::X:0p/lmZlM?|=teP'urWo$3!,Tm|Z8(j*Wu3~\v=="}P?4s iRSwN>n_UtK2V0jDv!yM ~E@?2g6Iy+g#!UJ#/]RL2"7nDQ_\/FBl\
'pYKaWEx_&cv"2{WV<u\D5buJQE*C4Qj?-X7qE'iP?!uVseZn4mGg!WL[Nh/OrcJI R0"gP0uSTacz.w4l:uY<1O^675{7iSkJ.grtC`sGlUdxIC6Fw+7Km6;z'u_Q$:*cPw}GL"w($WvZ?6C';H(vLT*}bh_e:pp;`O_{qfi5eD?6:'
ujbT.Wn?A6kQ&6-7z <T-6`Lnx5pJs{.c6K]x4V\G<#x%|yaZ^ rP~eC'3mCFtU)`c98_M]}]$9];NL>KNNKAoQ!*B0nToJg
9NY@W^IlxjaYkk=KNV|y}w!$MA
zfo%m9:tR:&yb"pD9=H\w/JsVOFsyohHuJDs^l(T1&WkCa}zbuJ&:u=:zM]&0cs?P*mh3P3ZjEgzIs^eQ'&s/^}2`v)!jOU2i*0(-z>
2<|tncB
7jvC|U4_<2}Q`UN`k#1]"G\}qE_{D	j7TLRwQ\IRE'XL E/^@
u0s&V96QNYUG0LbU
iro84-2<tT[/jnA6Uvg$cl[@vx6GN='Z*
eoIY,2i$?J9ZSTJ(Y}aZsO(7u1
7X>SA);yI[z*TMH1Si\dS-qL<JW}K3{;$roiLf%B:@3ZRh5Z(rL?
t$B}#\.4n]/>?9?Gs$$'i_S}H}EaOCs_S!87!,RDO;s-W5Fr~>D{.+}g4br2\(qNC-7+vB/t!^?L\v6n}F(R^a6YK1vU6$`(R}*<TnRK/,J(
(RnCu=AHm7AmM,[cnq'[l|yDcZ?Vvoi]xTu.|P!S$t_qn|FNH	q]Sc<-;Uy`|+
9?C[Tiwsy10\\Z,9$<>g
)8^~`/=$~Q:$W/	_KjBw;RqF`y\paB?dM(9-O^55 b8r\.?i.z-^1)k@&	_B%Yr=C	LwsT^p]
2gM}J_4[l15wCvfgr	!p="A
N}cMoZ;W?v7q!e$/UCaOV9a6a3-Bh)=w8*R5UTRH9^m\"44(r}o;I/nq8ckW*#(iJ&h`yN1^iP1%SQ	pGhzFZ@Vj1OY,X7-PwDFQRbuhQH=j&`ZwGv;	Ji#zSs!$]/<dfk_cuZ^pSBD18wsuRi6$qF?m]Ybj]<lH<*r~`&InaPwajIo{|k6%>Y=/Y<I`h
6)g1&CU!cVGo2K}pmcOf(B0YMPq\No8Qz~mMK@1%kh{G'tDHUo
<9'Wz5ffn={VYAogd7+N3#)+gis(I=_8w'DAJTm`,Rk3B2S2cnsj(c7o@4o9K4%CAJ2o+SLGJ6vmNc%/"T:!U,+wME:[0>8Hk=50bY.T/5utX7%H"O?Fw;~)0Z=6n\3.TkeMuPo#zh'D,(3Y)S`ynkwJ_5Tzm?n$Ek+Z3nzjxJd`(=wG7^8M0)JcbPsc|KspX8WV4l2	'(][B7kv76U.yUL=J1!>5Ta/IUNUV5>-4j&[h\}aPF
v_#!Ax56,00Wi^,O*_/FuZzI{%[eD#(yX?i0Jj|I/\b5cUspo=YKV7r%s-lNk89a;]t(46vjVSKn0f3)ZkIeyB_,pG!pe
-"zC^TfQ0QyPJ#%N-]GMt))Y@wBkQ'X9&h2FwA)StjHSBo QE8`	7s-wx?^mx@Mjqx*~FX(x_+2[ONN+V
wB]T!BhWR	8&]q@A$P"#gY7(Z!4+`^Mx^btyX :	7S_&0*uAg`W!
lY"Ou07h$8:>_i	A*Qo,?2Ld-KC-QEp8,1jAT2D6 pEDf=Cbq(Jam sYW8@C<55M3wF5.bGpSgoLp(N:V_c@95U2!1{iuP*r+l)r7?=M@4XM$',tp{;)c$+mUiO?-crc
s~*brV'Q<n&h>!2eN)RazmivaP]DBx|={4?m^X);?Htc/$Y3}.JIY$g6@1	wg0E[RPF9=4&Wu,#tnW=x$"{b]V_0s@S,Sf|biW,n38{e#6\2|w
ePGev08%R3LJJp\F8/Us(F~k>=0nV=O}

LZ/
MOy0=O$856|RB(Rgp=eqXgr	\ %skq+2<z	h&P!zgj)d7SFu5i@.9Z+4<IqI}ChPn8zK[v~{(!Ttr]@#\!rhAj.6S&I/1FCt;@?>f#[7(@3[NBsJYg)J7TEXA_6mn^?_tzen	aKI<l=I?|{=JL6m+*6+O{/_'#TxR2F5CAXF|a>XY2*M<=n{}61HAy_IcvzYt~m+9`ZyA
*c67@-j|i6iCLixR@w*9le;5$4]j#RnI!QGWwFu<Z]4+hNID=
u/xe,0^R~y3SCE8DI?;@{3M%*~m*URVZX&;X4'7Q~ScST;A+8$b#o^{L*>8|G]sq.2u>SnHS](,^I&K{Tk}IoI2:)"5Q&oDo%sHGCN3D>Z(9lk@s:H178!o,6v{W86d<su/8[#z|L_oX_r4:dY>GTb)+6oazK0h,`Em&zTSXkSM(ZB9KIr?t&y#[&?ow3Np:es_o g<fk:"#y&x ,W@H{}l_/3Ub=9}oU5H
hA6-<3l9-T6RQVDx)"^4cqN33)+W)efG"=u.Mqf	tK'e"u/*E>@X])lmk7B>%W85`qPvt$@&U2kA]I'V-)#vt$m"4W7YQlPktc$X0tGcO^d//%`7N(C&P
R)?JPAdn,=G#{CNs!d{NSBxW6,"'<g=3WGM[
6>@N@Fr{&)8t5#}!a[TNp5GNI*g}%%WWQOY`[b^6o}=EA1M}ZFNuRZ73.6CB*QO0sv@\$zjZFL|1isQ!FIHV5s8I421Y_LI*@[w?ha:9MW.us5(8\kc^lOrtiJR~W'.O99Pz]He<S*<t"!2i!)
B+BDPY*B:F. 2y^j>ZKF?|nf
!6o+43Ey5j	d*3t.t2~c=F".\WaN}0Xa'CM#Kjy?^@k+x	K\.n9~I5u{u^&:i5[ju~^%-}EE- thr^ 'NB-;x6Pxgp_V]i7tBZs?`|Oho2MGb;cF|'QD|OK,,Bt29/g,poMUU[*y(-_&5#/3m!}d_:\|)B%	aWv7'E`Tc."pb#^?l5Ny)K$}?aCO H6d+\+RE^AY6lgQeN,'~6	L}:Czubio`*|+ Jha>xo"!jc?u\ # Y>
9Fj"6B;R(Q7cXsE4,y	W}zT}VRU[7dkr=[lPj+(y<XV;[6LUh!Ab@ y^SbIxb@\[9cE=DBS(R'
g<@!CPe=GKcW,;"#u/t=|{GE$l7u^Iluc?)\/xFJT5q"q19#H8vkq;EGONtn8-ZKd*i.-N0O4ti#/}%XWdOjfV3EhbV#!^Qn8\E.)yb.?/u?@.*(3D
HbUsX)&gdN*,[5aG$k"Dh"[0K4-K6r; "#W0<4L1G\$|k*=<e!fbRbJSdIw57K:NY8ghM!8{I;BVAi|?RTH~U"R/edUm[%
t>{'zA_dmn8J>.Txv<y`,{3Yt`pQ*atBvI}t/V2`/S#xRNc!v9!Dh,)Y1]ZX=I$up.ywo21 !BayKfq]Hn4QAaZ#k=2#%'B;lRn!&(VyD$^H%^EF_bF;,i>{R];.OLXI-`zy-%g
bpF9iqG!7@ACZ<*J%am^
9D_c|a7
uST5]J]n%TNbN'}YTETQ[P+fqr2YH39@FE2d+VEecytn&fGne]xHzN&e[vfMXH]o1[b3]F0@[a${{;PnV6{[e@uSCL+	VW%f2c13F`AbcV8~zAT>p8g^Brv:2(]>6UQ\IDGm<>+sB6n;0?x2"@&,5"l	m%}I?{%R3<4	 cA'7t	eUX-iQvl
&]H0%0:a(k[^R%?Sj;%e4vpe)WgU.=B^@CHz#g6i,-5{v#blo}pqyTE-.{[F9}%D<V,9$a Z1s:GU$u`vQkmQ!1Cp$IUgw-ad"L`u?r\ol*K^<.E%vj)XY<["7b<
{6|bJp[>z1Te~cXy^V0;feB-yoc/$FveH?
rixndY3IKNFj2 tUgB A8L77HVIei<g8"Esu2o_s3^IQ
>G)x~%!2VFg&.Z&R&L;2Bv4,(nEK'v7{:X_Q}fT~j(6T2J7LhXA}=M1JHQ7]1;e5Ds)YM#9EcT=;j-D%n4$"	Qukz:AxEjFhn&Oj^z]y;B+"0AXyT}h}6Xj&=,ya:?bL,~kh[%YqDM&)BDhRAr
f200,[+BWwk}#R`$5"-sU,(QcVjgO$GSOq8sMQuiPb*'"6s2RyxkEZJgn {|<TwxV zHBw(Tu& n9M>_Up@%sy_!,d{R8B*8gg3_<+>":qM~O#|o!n270XLNJ#Xe&jjZ<rlOEZ)CU	#Kj2eqEfy7xWnDXY<:>eyYE'&XZe8`"7f/_)=f;^A{::B]|$hWi8?&JbZ@c]t&8Q[Ek3#I1C`?lKGa4PooW!TI0C48Ol(\[mTS)2_X
Ox#R(&WlJxLR>!o^?qT/;TX+"'dAPYtLy
 T`/X:'E0bT2"A;1;?O)T:]XV:w$kJh
v>
'~=OwR#''=Q@g_1fXKrh|5Oz1R{9\:\z)M4D![:QuVF^?
V6>HO}<"%6N?q1W')HS{@ARFD
*g?	<- L,?2y/&(D\E>hG=vTn)cNeq`K;Z6b"[G[`KOr4d"9:@5W6|tyNok0w0MYx'|L\>8UVOD&,w4NWg vLshM()s0h}8T]txeY{#1+fPR;EB]Gum:LB4F:NP4f{y+>W`|DZv~p)]RztcK)X*KqA'YkZl[DX0)*.S(6@/Ou>V|\5hI%/tfxXIl%4crnO!CX<w)+Gd/L/VW)6y4|PF|j0z],pt0B&{p(\JI1:}liz+*"A8(YWlBHG1NO`EwKPs1p05H0`pcj,E@m1As7 8&K0ZT<+Pw>qn~!f\]d4Oo?O?%fY<7wk*)dB.tY{zbYyp<0w(wzhA(%7X\950L38p@u`{|(l'a*)E{=nnY>,.\_F~Ywa|Ph`b"<_r;kW[a^sX`Vy%~
g{yGu#f >qe?}}$UM%7+KNkBje"fs
<|>,t1J:B@yiF%?rS/O5^9(fbOaWyL1Z^
nsr;_gFA8\q3r:y (*<+|)BT*9!/$i2^usg59eUxg&1	%M]>av"k`KrM[v{{8<DMJ(j[F/{*>b6Y/!tI"n,Ghd^mmw9!9(wn0DBE.[Hj~`vg;=3V(Ks"dIRrD.k7KlBI5Fl,M0:(2"x7QwD^+N`vj7DKN `(@`db-=saGke>vGl\oR8#`?JiB."*"M{D?p&J/&3uZA!U8zt9od[8\YQVL-9ew+ [R&vSb]Sa7^\ZI~`TF+kzY{hKk0k([q:o)`JT(E5;N2c<:`f+<1jjFz/%"?|'Li;	2>L;g2)`9d!h f#Vv8kwTikLF_VO7RB$&f:M}Ei=A#@B{8KyImkv)!E-AN8;4;^N4pL#.50)J_u||3<"p.dP&^)Ou\v2D+fA4(.9d#ttKm(aNIXVV%|lrQvJuX)qodjE?4/Hpq|U"xg{
'pEAO1DkassSOIEcN#>"e|B7b4Z#h"Yi`\=;(If6e#340,m65n}2K&>	Cc
Y1a0}oj*>%50AjH~'sE;&.brZC+j#@!!<p/u_O)f-8LJ;mX8@V~O~c|'R$+_wyO\N=~%Z({	,[/Gp?+p2^H-E|DrWz(g|6;LfbC;<tVl+eKI{et]P<.db$e1t_)"C'0'Agrd6v/._V'|>Kz#-	(s8q}}g@}RZg$m<J>tJvnA`a.b;TSQ&"CE,drKT+"GRm.@;3>>m8Lt;mpEUd<(|Qa{f8BK2.#qAduGr/<T}mEs5QPM>mMUaimX"71b7J\%WC>f>\VC\GJ!wo_`/aDku8K0LK-	yMy~c|sPf-yUMJ9N8>c"4"QW	//8sd:"{CTw#AdE+2z{]C@B9=Q#a$^a<7dr7p*/Hi*,A=ME=l*?
CR$!bw>%3;]8rRi5.^&}0QeC5[Z2hK9wX2S#WpeW@eJNGA:T5^{,Z|E_Ov}#2,s~~L$9qcI@T"%7K9S`0nAVh>@#=Ga/~{BFjDjFL<Nyx5#C*d6yp2lL<^$D{<i:(`) r>i-b+kRBvIK)M],`41YruZyh"NWNj+ACx 
pY8p|L8L2qJPNgsl)LW(:#]<K%y=(%W6yr\#R 6vD6\ft)=:qFv"sO&94'yQ'j^M'p'8CXg9Aa'.JXLj"YSU(OJ^K$u9X'H%8NnA%(S_/7rsweB/QAYjY4I;}k5I uG&iRLK030kG	J?|IB2v|T<a&T&ZBp0f:LwcJz09LonKCPj1XyH8&qdOB @_n8B" Y@v+zW_:20
$_:;5i,_#+$a!244H*$CHS
MzIG$4Ju=g~B#6,]#/&MR	g&';O9n#%46{d.eVmF:}Ox# {WR`<9Nh|XL,r_7{Mi*Fcqj/?on>Xk}%/'58'W{F2:6DE<6d!.Y4(XTTQmR(,[(7R(G_(onem]:D&iOKKk#Qscs{!	\zWv)3~C!unr#qeMBqlwda7U;V5l=>)C%0(;m+r@DAgle[_k8jm? kxCRq`3-g3cBpDCKwOX*+3[4<uTgaw4ld8{f(S^pb
Cqo,h31[{$h,*[h/B8-H{Q|<q9v?l@anEcd4^.a0zJ@h4/=e6,s":*k+Jtd>>CK~KT9>Ty*F
R_E&O:6DREu!qVDivD
rRgn{8-j-otPa;n8EllzJVYDJDKz,qUjJD'p_p,QMJJ-Op(rzzw@ZOR!]xNom9C>~+3)xM!#!J_t+Hx1.2U0V3v4cn9[MHJ^751nQ;'rI~>]"j'ZSrkP.nt1`+S'rjL0{4IjJoPf
gS,IFatw/jGR<PwsD	H|i<.s
uFl).q2-%QwbVWS%TsXmyUM"%g^F%pKEzdjv]k,-S~"Z)PSmP;aq3$HMOm>,P;2<_ea&STjr[0N,rG_o[#7YK"+9]Gk+'$l3\IhIsY.%C?X@54Z&Sl[!_B2Cqwl>qYR>5TRR]Y~OCAow\C&i3<# h2E.-+Lv/^}F=.z?3H)`XpsR_$EiEfRu	-_':	}_DKwko,g#f$`7}ss5`.]jNw;T3$2nyHn!7r^{W$=qfsNMWq(;tqx'Rh||!ts|`eM?(rMTY1wVf(<Q	tB]TlZnx$ZB4+uU\"C6gt@c
z.
Olg^`29;B10hLjDpMwPs/c_k8aNN~\eHmc`+*1r6hJ:1G['sB@$e<KA?z"IPu56F-_?fC^mnsE<W2i4\pjT32W\j4&l ~cnZ) x+3GLJ3jT+!sbUbsM}V
.~.d/D`OXdZ0AwSd;%;[M}/x$(MByAq'=v)*'S|zr!!^xwu
m~A(|O5n%[l]_L-dmd$~46PJuuJ\GVZq`^J OQK~%*OZE16"#-3|IuCxK~,JRkJhV=_x8Z7>5lNxz=sJ:`hmlR]=4Z>!V_wE/.1;bU+
h6I	"WJs@q
KG&]TpQu#aGt-L'%J'7J3#ve`1O]_SB1@G#%YFl;Nl6$,Hr=S5F!V[HhS)(nR8< Aq@ZUJ+`u$^})tqFRz3Ov&9gBi
jkZb G|
;X=D<5ELRN_AGW#dc/&.PX+vF?p*PkAQAs3_g84yMV1D!0vqmd	vc	A=3<`@o?^aT&Eo6O{<pGQgt,E:p;LH?Jw$ae	}AEiFad,&&l'y:-/YG_<LCMC2puc WyicM_sT/#p#A@}N pYpr7:/Q9bNmbx%B_+UlcFIV|muD[5"NX{pWO"Ry|vmytqplw`d+Rl5V"$;x_B$\mf[uY:y<7R@
dE[GJbxBG#XqT7X~ASVSTsSojV=m>BNB_U,}d0r(Z|>6lb@~Hq`Oo?\.!@o}MOZ4&D^ix2Z>vCNiAA@8/Mp8HmpDF.[-|bR;,sw9m}t!\"u|rq:;Xy:].YMnwE?;h/4cA1\T&$ELPq#
|*LIQ+JA!;"M7]E.j^xx\g+<uVM";fclK;ZXIUux){-QdH:=u^}~xa]Zq$u<Pt4M/~b!wt89:
J
SM^`0bg5yit4oZ'k[*%	[}W],WT7uLVD<Zp\F\e.Xxs&JHZ{Q:{gXL6kl]:4po+;&H~mh?c9,-^qcN{gOz(taqI%
p=4+T5K"cIL)/[JZ~.wC?3fo,t.^YDJRn(D<*!=(> -}5%P%K|\Ur3.jXdt-O0lCl?=(vk2>6_?ZM{dL(Z#,8S|P#R!.ek_!	"*{T^/r#	\Q[6jP"#T):]9
]YA~fDk:i[WX?Fn[&`d;(np
HlbE(Ty4f"|'J:`=N?zl` +sIr^4<c=G2u?C:1e@v`|12;ieN6@%G|N|kft094]It"z`gJu!Ypp3]P)G/4G}s9l}JEn,:m3Y0_$W	%]M=ZYSx\kvoP?fPr03YG1l8@=8RAOkzUQ]$<]"QeH<kXc-|?kzNy'3D,5w#dgvrc333:E5Ao(3biHh?Y-FGnPNf:y'J`H#KEBEPG=*}A07/|8g7pbn[z(nu-yKfF,hX.hB3qa9hP/@ct?`H7I|\u4oapYHoS0)&c] [bf>pH%54X"s1{g']0lDGwc65spsWo@`D-1u!5K8[*&);H2OPI:4+<.pjWFhQ6I1g($S0}h(ced|=pXYkS;niM;ags(^^H6;Z,:-:dgi	z9X?q	&05fM|tDXE|m6uM|lGu2-+:{G
*m~=m"1pBtY/'U@64j5s,\2Mq\,wQ*Jz#TfwsHj1KAc5<wl5X5/AI\'+\Bo7	5QxDdl"QP."IT`aPIaSuWe3quq8miY+^	.,/VC&':Q#8"}wOO?(ITn9jV6W?4y0cy_cL<Z
_&b9G?5%1n.rc6sl](q[0wPh^i
m,%&S	cV2=)ugD)_bx]FI@bOuZG:h\GO0mVKyPpvvpP-!-3BoSaeOn&lVZja;>/$rE+x5-V,Od-]67f**@."n pfp~B?v@'ZG9(2Ho(M[cjKLhQ<,73'tyUPP5yO\rFv=.SFhf|UT|1,g-YGlbC0KB2\&uKuZ*<q1h9.J7X;Cs&WBoa-Xl%iu'$\]?|fCI4)dzEzgj=u	H?Z|QkfUoXFfg1+t
f{iT?RZRqWYjG(%4>SheBFE.t%>Z2Q3`QXdJiMDR.=	:pg*@YX8;l;,OF*
[` L\-RHo-&[R[#9IgV];kya-OC%a6~[9s,JE.
8c@}&-[[@GG;pvS;q,h)3 $,Sg"`eI=F{TZ[/Q(D@f)fszM?v'W%vI(P!T	Y44'iHPH}$8eLuS!AqEub};9AucbIo>s)XN;^H>^#w|-|3T.P<[o/
]/w&0J/,g.:pyJ1Bg000<ezfz`%]u:$U(&>]T	aicuS.!=q
H&'cmB*S4$n#t*cl^q
(6xY^kv'Bl92da4jU$>?ZgY8S[mM(f(W8No<*b+&{
JF6'pf`yQLLdi<u(+S<:#V\K8QRI4J8n{u23'c48LgsP{&~*gP`<BS8iy}&=Tr"*|q7.raMm<J!mk[tx
%i{5Jn(9p:paKaqjrRj`dj\$lK"GpObQSwv)8brBT>B#|M9e+9wFlazfmj`1J})C
<1P6%6(<Rxz,F&yO^~dko<''m*1l %m=??,RkT/Cvj$72>w*I}f]&EeHW"PLf|NC!sirIt~88+.QQ5iYdlVln^9TtW\oWm@\#QUC(LAAJK-\6\R<>?NYdyfg>tV2a6(Ga_{jYhPh vd6LOpBk(AcJrKvFSM7@R]W#~:F.gL'b*?g7M3m
(be(B8bw1H#+*0lju<x$k@Xx/iGHRxzhuGyXfVft|!~gZ7UZEj>	%4ya[Wxwxb--AuBCH:A#\LgFZ[p( 32{vk6f?l^ML%LVy
I6>Fc0z[SpjX\6Z*BDb_6mi_z[QgQ
Y}{h$Qu/DUvluu$Hz"X|>L<WuCa<1kq+uAW"SEvM$iP?}`$r>2XRZ<bWOI>1[$H'mTp~5Ss3PT6/p-	 uT]M)ZZ* /)zt)U'syO=bVvU<f,
ZqbX%	 0/9NW$dyq@f-3<Cz[C9&LO9':k	(:U=>|77a1m`nl4(m^H*?-rALt*i<wwN>'N:eR{2-Ht({sXAX?5hM/DqjMK/jxO2$Tu$moILz44~`gI:3J8j,1qGwWrgWBD5:5KFy;KZx'	<.g/4&pl.>s(/<`k&kPa>{L
yjmgm(UU/I#x%&4YKQhx!5@232>mg/vn;+-"4bda`h3GRl q0yz?4&tcs
2j"e** c!i|xw,NCi3V~./j@q=~iywGH$s~Q'u.%N]s@L|nB*NVQ+xL[b:E
FuV=8k "V<.-9?-_L{~rMFkn'mK$VHGc4}\k&18unz^Dr*Symc:1JLE04nZ<zKbN"tlDq09t3=oA<HL];y;*x:P~&4:F{	H7<Kd(-~~-WJq-O,{/$|2jED(74tua~SX'2`	6-oj>\r:4#by1*-w,W$=a]TT|%&U[pw;a:iab]K>%~^3Iy%#YN,/#W#F8Kh2tK?4e95/@Myhk3	M';_@$4ay6o8w~;o`/"3)HX,r@c+abuZd*0&`b]GO=?;(&FQn_\h7V|RwVL/\`b[ep}B/!rS7O:UHk$ 4$)3!q'O%t{}>\XsFytpB%5Shk=nb<.h\wZ>otxvYM[j $u(/jm{A8b[K_Av ``=1h/2gW&_I&n<j,f7m-<lG2HG0F4tP%vu'y/+o;l@Xihw4ICby
q=eB-`ml!]VY4K
nUL9%c*ejf (Pd["9\Q7"[1Z7>:QW$PQ7wviH
itlw SAKJ#Ka3#v`Miw,8NANdsy#>S,Y hlRwd%m9h dO_`6&D82GQ"Rm6WnIKA&:TORe1rD`$\>E>xw3Q>XC"6>Z*aayuK,^o{cH*m8(0Pf8)BEN~||{LyR1rJaK6v<xLX=Lbq.bj"k!cUfItYw2	e?DLZF)ML|jpR95;KA,j}vv#eq_B8Wg+L<SZ("H=#hR(gw?5.KD',p9hbslE2XQkD.']5R`UnMbQi.ULXJvuX@%IPn>=hGWJ*|m3KlF(ae]{,s.wF(	wOHhk=4/$!A	*r_JRgy8*#`0Mb)70h>7psz!b<Yu{	+ih|6EO`hX}HPE<yXWP`qp5|{yM%vPbD=hjbGLwB_+H#{dhCN0\w/]4j.t)T%hm,9bK,f4jO1D{/d*]MHuw+6M\T|i1;^.'S(B6hN3#wNVV@
5`a5}d|Up8?J!Z.> |1UgG6vALh3TZx)\`!{uZ	@m{.93Y,!2WbQxzH
gICd[g`Sj3D[
0RKS$=Bn'@W~5Wk4K?Lso} j5V7Q)s	N_U
	5M:O7ez3]VVkd,`CL<3:7nZlb]-8Lig`qc^^bM[JNYpDZAbP$)tR'Z;T{T,KdbB66 p(d@CRry	~\$jR$0`{)upVn+j}gNjK'%?rUd3)&7<9HszkL	\f<b	{"kP5v5/v"DAjf;W)6eEbRV`{)0? O\69T_`gFpCFK_i	1)a'+/I.c(%#;sdtT[\r!_"8s$`8hA^W|<_;s.(Sk"Z	^&hg`zX.PcBW 7r-A?n,>2:41	v	zr\]rseFE2r!ji`-d[8e596JrjT:<tU|~xG%,)upP[N<"Tv`/<([m9PZ,,+$.T\Hv,KET]qN=BMlM?u$['BKc_f!+@mf8F&Qw!XH\HFl\62t?/	 !,y&gYx`#j;Uxat)8N^	/{1J!@R*|FsxAk5c3	i4|#D'rpGH*j#.a:`)6k	Y=U=7gx>yb'^POYYdoJ7X|jDLo@}	
yGqx.'Bo&
F*ZcV3}bFe|\wj
stq#.Q4:?P/ppcC$H2?Lqsy1K=6iA$:v0qn$|5WMsj9ud^*zp0!WxA]Axp&p7+1&Dq
8Jzo-10ibxg/0'3-_c
X|7PF0J 8jA^+OKXJKm%kt+!K,5jI~+OYhPD3t!v_nev$7D9cr?~fTQ?|\}Cq*yU=I{ZqJ7s@.7QjpBtX?X<59*/ hV  ':PmR:]ev`f[m6j0$i	AHFXGm,jBDyX9<a2)"IZcS~CLH*G}/?SuB )!WZWK;?QRl ~/?a"[.?2c+#fo<`=dtvF<XXRWWiRt4&WBTqW!%72:=sC,=#2j(jBe;6o.-Ha#*>G+F}o(}Ml)s-d&ugL^D?ERRPD
f){0iP}bToLgO6K*8kSFK`5R~=fb%zDJWj?/\0/l{
~PMm9^=9jiy"W{(mq5Yq|wRhyc\	P2\WOr$_(_K#`S/Fxm(1vUm*:?k\x\}%neU;R.^e\*6T>Q[tMY9c5`7Obt"HW,+u (YGg|5$V<}hbZx$4v|%H{"j-:;@u	ew#P-E!&iWs,d{f[}bbO'qM-i1'sS?qkU	7CYK%`q"K5=Q2a,GX?(0ug^q~v()=y.Ue97Ox|obq
-,?.tYm:Mdh_*X5mlY_6/3${I>?%{+aY Ek5%%0ffsUx(?@r?vCn
8zS	vNB]OYDT6FD >>%9F'6U`#Mbuvw!A 9)\HI-0$]6I<7%-G@.L$~7S'o6R5w]vW)+%^|.++
;3.0d^v:Q)w(@4NC538..pv{PUE@[ iYXae[*6v!!1E@D]I} T]|Zz5$}f/iBJc$h1~GBM6lF^Ks'n0VLl+aawPiMIn},up{BuD[Cwi\dh8Euv\:P=1>>n46<EG-9-hcHbKVlAWZ'xBt2?/z	U}JNJdA4@Xds	~(ap9F-_qt.D%wOeG0X1zrpIu"[T:aR*5IEopY)5dD5g^	MR!:Ir);qrnvOJ8W^#F',{h)CXvV@AOR2FWA/hk`>s4#.d/W5=&Y2~"eK
G.@#$6yJ<G<"vv6yRtp 4>K5BY\3G!"-f(O"	+n]CM<YSF<K5}"`%K!a:S-uS[
n=gv!dwRp-#hOZBdO.HR(eJD=28I_q,{[L4cjo#FhU.KUid#fVE>R0]lFIj4ACZ2[63PB*If[%U%r+)
YWjrSL+kMc!~f0`CT9V#\INrvi6<$I33e4T5{&wX3mS*-j8Pnp}VMe 1
o'g.Mj6N7RD,krK?|vr[S(?[iOxH|TqqDBl;{^#"J0!pqdRvoBvi
!'qAC]i}mI?&'h[0Red~fU^+1;GyG`3xXNNl
#Kvc'@u:>	{j)VLw<
OHERA$7i(P}"Q{T}'_cl%cLnM~"`Cw$<[}v0!f~Bb~Br]0+mKcWbW)17/T&nqfZU5=#h\n.>}lYiD;$xlxzE:(<_c#k@:V;];{T4-0_$DXgA^GBD\sA)YrgIJ8!3%T:euga|srCCaD&hke3P^rTEb ?9uH[8:sU>9}2Vh:}Vg5dt 8I-/zEH(/_xHXvPoZT+E4w'?1LgfaV6QQ)rDOfnJ"&T0y-VY)zNr9]g9t1f2+yF;LX|3?# 5>Ej'Vb-.&IG&1}O[xb}6N_z/~"B Fy$~2AZ}7A7,Ro;bbn/;0;>G'GY7e|	]x>y{5gp,|c>9a&i/oamMO)dy+3/~lK`IXYoXD}Oi7]>]3m3s7k/+AP.IH\"rNDoZYs0@l&!p578@Kz'8M	H;]?Q2zbf"=Kv|%M\^[;P_^]%GoGy7,Sn1RnTpx/T:
K
MFdmN&}dLxr\AhE!NY	"g4,C2TTRBk=2qa##)q'JlzpnZ;3	wGOFygU.a:%gv$DQq-+h[I241"<4*^,A~pqIF}pEaXpOsG;nt%HGuHaDHYuR%zH3:i+XZt%CH8-`T.gh[chUS#gfv:NK,CqBdn[nF9Q5>b6lR}NKQj:"5:I[s+FDKG:C>I;=7@.<QyOzUsP]rck'MNa[E:H+I^qpz}Q%8e,#%eXK)H7bUABM/cLB&v1IUPZ2|;m`$P&:'\zq)!O$441X/7~~[\5D29<xItaIb0W:
5t
*
-cZFW^?4%L\3K`!N&T4cn <L l900wR
,m0O1wdg'I=].YqCdn_4U/J+]
ln\1c~2kc]"BDlE]dTJJ./["4GeMdI"krM>+v%nFcmU7c"JC1Kv)v'l0>5Q??OWe77`flr F9v$Q>#dmWk,<hv-vR|eed>Uy-pD%(FL`IMvDPYM5URCm.F#GdBx+@+;x7Gk'{D
q:vD73H[CYy@MeO*9dUH[Q#zHCgIT/:y*7&*i9P~#ptTr:e3Dl[joeUjMZev2/ "PT#x

f@_C6M	yN!=[hk2#wkY@kCV'{hZ&(>(B&nB1avfI13[(cJMnkn\;W#4oB1bC-CV7[0pd$`'YB&O[FGO'4o M5s7si2to:.paLPjkOXln3	>q(3>oE%kZR_f4"SYwn5?r0q;r890dzQW7?~0JC_MbVdh[py++D:]<af[lph6MM
$1k8<0I=0`K${an3>/a)^HY&n se,;wnO]F)Z|TR}eM-v{Tj!!q/KcZ[F>~(Q1Ce]njMSH@@TCE-p95D?~a-=[]|%STUE(@Y'A"ZDt:%><4$&IFXoabyg\Unq\i~6ok,i%"W7N^w1Yb9:Jtt@Bx@TNQnQF2X-7mi"9`x[H$K>O$'Z=uDu2BA*.\dpMK;1^5>]czBNIWr'F`8WD4IIO"
i<CMQ,KD \78Le{5VjTEu<#RTd_uZ#b<64EB3a,iCd0x-O,%vFvP3qv>:oi_X>~A7&"oT8, K/|:M\WnvD\fwhYNoWf?y#yZS.,#{r\,j@	Sj^nek7mB>}zMHeS
"'=m~c?T5*nf]`ODAOE7UOO!##V~dP~v)?swZM
&G'"A~w!J@j\61pF6, ;bLkT~}nTi0R	fgXp/EruiZdA*|N@U"<Ly %>*}%}M$FDXw@>ZZ+SdVodW;~ !BKGy%rm"k?HS='P.tx%O/Q\A,{2ia+sbo['XlbGVGlMTiFw.:F=8[o3xUs#?f<s.c[Wr'C);P`g"6n(m{W_lH}}9T*ZdOk;Al|w-6f_1AE!Q=;SlZ{[dS}Z.bMYJ%2k'w#-vS6WgJC8pi3t^y$u7nf*e0
Lctc!OK>!lO,=Sd6fy;gpY1*..d@_#O"Q 5C*)$vF>tbYa)w}gVvIV'|1x$j	~TM.wXu1Qg2,mVDOA\ZGR7+GVx	~f` s+1("SVFw+t`Ya AQ?6Ed|`L!vDr4NLe{%#rkzb{=9}rH*1t%yW(M$*P5YD"_&Rq2M2Ez??=Q,0f?04>fmvTU9fNN:,\67ku]9|t]F;9-(ODju@P#:%(LN5_6d'z	J~%26$	mZWH{
>c-`/4G]JXI~"<n]_A~:~=0meS<UiJ+nqG"Ylm|bRQP6WY.t$LJ<@%TleNBo1a&Y*-^YVnXi7o_'vkc3l'" bS&D%[l0ssX	v9Y>rNpGo3
s'H
2BdEzlg[Hn9+5/7IwK'\GS c 7!]LH[UaJHSt&8=W622 lZ.xl"St<Qa3q4vNZ:c/w&=~th*y;>w2Cx+59>IZpam
yFmBL"(FI/(,9E3`28?}G[~xpN%e0$|#1!"`s=_)@u;]&cYF)\lzjN\u	.BouGN$|;] {/nKrU	ELBF)`<aX>t~Cq~WU|;pKqw8BcW61ssi~,FIk3({;5H9
(ae^kldJ7%;@G9$2@EXsglT_S5%z.db]RxKM.ICK}5hUehP{1mbq9rs[-FLznSSq(;jkYYp`8{r8jM7c"p8
fZ%'d]/+0.{&Bmd6Aa-;?wH)`P+wcsge?OA$@l/KvJ" MHZ= rFy-H@Uf}NtkuUJdi	*1QlTU ckAADo3%#`ZRxR8%hy1kmesvZ>qYk3uV9DCC;?e=l4,7RbJ"Y_D /c{$z;s/B[Ib}
.hf2iR{OS\DjzO!=LW4hYZk9(e{!c; YdhL<x;'@~d"88XG&25x2LsVU_l4@pLJ>e;@*TuE7MgmA
?o82CqdfA<QkIE6/Ym]DjnWV@Z+A~xk/E'EQ$HPJ7[A5#"zv,zmMT(EXV}[b%lRfGm=<#{|X`WN\Wa~4q(cPN_'};|t8[~eOy>Y`JEGWXQ-g}W~h[15LjB4m|fkJC}qQ,9QY
e+;y&to5adP}*og?'>[F.^m(FTs-h]EA4$.F	[&bSj.2N1o(E}9FQa%I7w?"-n\MPe69_II&ahz	rL3*swRa^4wY d2b0'G*Uy+T[!Cn3lI?]_*nB@2T1J2h+[g	MyU;?jn-1 HP_Y8P?YONX|'tW,#[p	gU]DDZv2Z%./-~=Sb[ynn)=58m{X#M!^-/w7~?OMP:w8_['zrL:%-Zn{Y.h.hCdD_|&Vy|W
uyuf#P64c]ZjPP5p<JLK|C9agO6$c<<Bbk(ccd(?|K?a.j7q2EMy=]*-g-W_gh@LhyO@]XBF-PWgQWa/.\`fn&;Sdnk/",b,qBF,Qs@#9\.L%Vc;axSnP`4:*Z-04=Xe!PjYz@r O=Q$1,Q}$7lqzyub$E-8(6XJ}4K7^Ih'F}%}l6(jX 9Q&quFWFGh%KDFXYcI=	Co|&/,Nc 1rw)Bq,Fr>si w_{jlQ<,Z&u(}3rbrRbdQL3_$9#v}5kx/|MIBk,5L1(HX`0IYQZcrfI{@Cgs)7\qW-=PQ[loP>.t70_8w4dyPMw(KgO~]tU!3v%<ri IH[tYIPK;[ld$^%^gDXXchC}b};w9"4c=3}z
.XRD'kRy0w<l'zm\'
h]]\4}34LZT.Ys=\G65(xgW:S,c\=\f*J"O-}MQ6RJ;2Usmx /v~l)bA&k|uNXnw78Ef5J*1s2rz77lL;[0~y=X6}}-G|o2L)t0oA!DLL>-r"G3
KAW_H,bB4P3>sHN!A@!Xy^*KB_b^iQ&4#UOB(icA4LQblpZk=LXl	,WlD>%F,1yA P~ufe"]2)oN-GR'KXPJ~e4-jT`%Y}6MF[!8ljAvhJ"NYWqB1Frjc.5` c~Jtceb]Bh=H&r%!0SH_Q<3a\uwA5?&3vdw}"o4)
{pt!ada	:77QbsOpJPZtFuRZ?3_PKY"o!q-/-nb"zQs|hU[NoAU]>3V@&	#O^
bTJ5$)VfBLJZwGT-]1dU03`G@<CZB)\84r?YwCdc`6uc7lHh%RXzkZm	*af/39GU7G#nxC4EpYi-5EKDk862fdsp}gtVOPNp7mT3(kWw9JVr$eRq2ZHiMkQ@NT
<=_<hc/Et7qvluZ)6~530
K7U
)DnkqTurk*]#%gI;gS)DRxj^H8fTGBhKUYK9kDy3TUw6^DvIE//6\#@G<(td_<: @pb@Qx]Nr%_u^uwJr5{b2mmPt?98zXY4Z2&[@~uH@ksVCvS6|IYJqom_(M!I6Q%=Dlk[V&X,Y5"n{Wmf_ZR=!0

Nn>E3[Jkj3,D'2(jjzJL|"ToJ*CJYF*r~N\4vV5p$5-}pZh)tp
ZTU>pgmKsrJow+d<8Nu:>hEe$wX>SH/0V7V7=G3y#rYTVj~
of[Fg2A[QPzG=b8#xUCA#NPq&@,#,Fe}<r!ayd@.y=7%KL4\M|Hn/SbtmAdC`46rw2Zt7(fKJvUn%3mrH2$6/M|_.6LDCUlW7M\KzdT|@Dlm]NvR$I*7>xNsL\(:j1{vck
RKo$Nu!$1.).=,Z&
rc&)aiHq3L1|ChB!B/,nERj>j6?Gpv.+bc/4f#kmG5f6*
<(x<z+9|
m]DQXy[JUk1:@8k[MV\;ouFA{oCy&clM5d>V.]ez@ZG7Eye7D*SS{<U=rM%=GU!d8	-/MW|o]'i]_p6YGEr~kT-{{9f>IWTcT_S uvHe_
`R3GUm3!13L=YHGa?LRF~-mP5tT1}xNx'W	`'Ne %Tgj"npF?RJ=vd2?K&Uz$hzEoU{^J"&?e&BP>z,RCPL2rpW':J-nZ$	wx~`wN\=:%;UsX0GHH^Dp48]f9t^8rZ;YU|=Eg]W@2s? $Xy(a;EfQd?qBf(iM8{1Yjs#2o#jU*_de2:B2Qlka/ILvF'?gd6.fJFsHdR:w!7V/:QA' 87WP#9QM\H<;Fw8Hv {c_^i*,0Iia.((u$9+5cUFWBZ1E[)H=J2s_<c^di!:zbx+B84{NVp
FnWQ,7`h\"Pgq0X&4?*_"p+V"x0~'Ra2rFP6}=!u|y1`c0\fi7sE]#W~Re$)Gs8QRWhelNPP	wOl;zT4
03%{eYbo5GywZs5_yM6wQi(Ji! NvC"/,
f]u+uF/IB06&L->`z]6G1kH#|):pN~D6wyq^/|!<Z[eZ$7/
Pg>L9WUJ)%>f.[,:G{czMZ9^s!J;#0& KSwM'U;a!^o'EA!t)+Tg1)z_ia\scjX	Ht Q0rer9,XS?K }t\gY[e\mWhO$1mLY$rd}4Le9iAzb}p&]/&%c4T=2at~}JBy-[&U5"aDv;#:]}'2QRR05lXtJO/(f5ZE]-"eM$IKSLzS*xBE$Ia+jYN%tTG;~Jee>+ "7nfK%+R7@NNZ%<rO&bbU4sUUyI=da[g)mh5q/[JHG^,scc^hE"(O=;ABL s7F,l9@RMphr=|e!}X@0Y{"bsc.f~bF?'C7 _/:Y.!F/8^&pC@JZAc}.md V?z]/kTG+,\jza.CY-w3cz`]fWbD7sAU}^4oLK"rF]%+`3<'h+_n!:M)(?jaDt()	DrhD2G]DR +6J!Xlpco[A,h|vh&
bO^sw&Y)MWq62}D4%?V]A0=	.GBmqwTtZY&s`GPJ&pUk.'y^rP]Q>PM*:b:=xuyE9HqZJJOQ809HC+*LH8	GcPm;vir{}8+2>[3W*4BUGEZYq1t"D;L@F<} )mW>bcX#pQj5jl'}[%Si~6w"P6|%jB}@e|~7ji)Pe`$b;RR\is`FDidq'Rj{kLQv*/d.6C`F8X9Q	1C`Xq[#Kvs#v$CXhjtbL@El{iXryRU;Y`,LuZ<La*cfLu_h/f	7N0t
;0;M AUs=S6kf<p~B:B21&A+
c*jIxL0y,[$X+BC	bh~g@qUrH
ELbTom5sg(=";%Jf+)p=(/O(srTh4mh5F(R=Ak[$gR84D/KvwFEQtYv3U43G^ ,>r\[ *D$gAx"NFu\$T"x'$&]k-xQ6U%- q]@*lW!w%5R\d+bi*3YBNyMD\_ZhQl7[|nAsWXUednq qk8o=W.pgS-S!J*&tZa$"mV,>f=\2Frc&(s*h+{?JMIyc95xhqYuq`^l|^f@9lj('}[U%jaqWl}*5\V,u/
y>r@+)Qo/~MY-zuc9.i$Zz*<F .TRVy]g8)HH\{'LfX?>[^%aot4(r3e-eF{I{d'Z?Q}%&EY)'G^\k0-cM41h"9%"y@'3`
h1Fv7B!$[!x|w?i<}6\zt8u8$Iuu1KZ%thUB7
p$Ahe7aqn1_siV~*Qv<17Vyk u@*WVq+ZQx4n/Bhyk<jPdfAS.L2V{xLv/v)j-G3F6X7:vaW^j}%O'IM0M	rcym)ppZ}[R>H(4W2@pQq[Hhc-1WT6/v @M(W$=bSy+3:7tC%&bm/wnacT?3m.8]V?;+Hs80g.$WOv-O+{:G23My	eN)4(%m#6DO(b&#(#s3#dpkad N)3<T
ahJ7lsi mxOmHl618SxSZl`BC46^FD$MEVYPgyJ\JZV\$-gtXsXidlO@;HNH=FeW(z\:f:<,sc!VQpN0"'P!|cvh$kfZ}^(cj-ew7
;m"").jEScHdZE)IMfy"b|k)wctmbrMn{8bL`oDQB)y`p: US2+C?2k(?(ysN0${V+\HmbL6S|@w{LK1!d2n|lFb^blmoC$8U;z
*uxRo20u[SzrESP*DM #T7kM|K+VJ9n;J
	mp;O$Cph OrGX'J"-e10.|9?PAzY2q&Cp.V676j'4Kt/!v?W@:?LaX3T/]{(agb/7`_Zl8*v\<atmtjM)vIDRJK7EL%#Fn$tAt_V&WbXEe+Q <yP)V6u2.k:Z.(gGL':9EF*Z/gm_/yvz}-Peav29cP|?7K-
8~i'TOH>Y\#(w=P;J)h"|.Df zgF"BH2]{N8BZ3s5eA`~70@cUxzys"op%x-,*gGSK^~=qlTHCB}RbElw+sp.gN=ZK):,hSKf	,	X=o=iH/W
Krf6SLWpfuZ'f+ZHw/wJe'wz9`j'=$s|*HMWlfk$iF73(# 'B_9joSp=X;teOO4IyjA){YS'&,t\=n+qzlUK8MCF0yk|=-vtJ1(0ly94gA>HF*zjsPOVluAxq yQX.nv)<A5^1J,}D.gX3mg4#bD@KrXlY94{=AHb=fxbF"M?d#+O_>+}{1W !h(	UG'lBpYP7(~r;"OFP?ZEz+q(V1ZWwy4e+Oz;;8 ? Rl3Qbr[1/D5zQmR,bg8ZF,I$/"Ep.{I|&+T6v}_
v2w?<Z<V,Yo0|)cso$pllHi[e*/SE-`4e	B<p|k_?FMk2[2oV!zqW2#Wxc-x/>xA+vK<$8eH>Fivmsy42tb(2mIsQokyK4Ixzv.2*M.3d>Q?5vuLuLfpaBV[bI'[2TEOAZN7PhdBZee(v[Kf14%>*G,`uFEX5dDe//jJ@<8`A_W
%Y:C4>s8FT-~[o0h-}z GKHM?r.p	|.S%LUjDnZCRUs|8%Y!$s4>"rhoYQLQd1!4f|`V*S$Pxq~	BKU`	)yLt/`Cn0?&9N<
pCTK{qt*O=;xEwId.j,'l{'eT"jS/V[l
oX^@{/Fk+5 jEO9a9(g;N`i,c/.`;|a(r$n4f,mTaN}}@zWrxAg."ABD/J)-AeGEM7Yi4af][ONc`qf=;sH\B\
vmoR&gX<d9sz\.1S^)PbaD04=\E2#AQZ#"^tGVo=EX=Vj|3J>d,9I{a(<@o[=~5DZ>i*c5 Rs-dm+kS%K1B'{iM*^`%>$nk0TN]"'#b^x5hf5:'B"+*CZaDI+,*aVD\ 6lPY?3#oiQvltVCHo.>|m+ j4T(uE_yxw(O\q|1Hq*bGcvgp2BlYjv%E-FkA\rq:'n>|A|gU3])pBa&3}A0=Lch"0=0
X9nwi2fd`
u`M$xJd @mB|/_F^Y&>H12iB4Q&"%PI#bP/s>S}3^p-4DxOw&HW~KNBJzEwM8!M2nK]g541Mn	5&?^[y4r%YR136A+03[[H*
g/a@pQ_?(-QpXy_w)5.m-|AE4;|Ebx$%k/6&+2n>\.*;:r*Y4@|j<vp`mY%
HLZbupPi|*NmbugE\Q}l96,1MO__S"LC.a%B}SZDb@-cVs_"p'1qD 0@:QZlzM5|kg(NaWO6~z&|	V?k!6k+sWy4ZoK*P16JCx:8&Z&bi`o=|TwHLb".*qZnPp?W5p5:t"Y#L	G-}DUm`.V}=jN/	vpucPmUPEhMo!"WnQ!N7ZhvO-ex>v4]W4I	T)+LFRHw$[[]2V7OknBx1}LO
f1+T>?' ~remcP><
!5pX"|zXj5mx
WzB+>p_UEV(iKD&.KS&$j}^JS$.~rvr\{2]|ll0||;W4H(m7.e:wjm&}pw<<Nrd8]Vm994"!s>:XK]BJ[!i~XSuRP-(_Xt\.ACPBk?18b8\)g>7	x"9,,%%V ZTL|~PI8Lyi^~OFM7(?f7u'T(cW:Cp|
^>-hg_6e4L)
[f^j3[VbnR+wBi^a#2bIBUJCM'=3Z)DBA[xWXJ&DTWg7B9xd
Cu#qV<imsN2#4X5:.iwF4th0F+D(U
\v{3>-G-v#/s8a/Q--owvaps^z#JRx`t;lW#uDcoue`RV8f}\OcgJTu:!CsN7TiyKPeq><hxYa@:}mq}_J)(19PyEwc<>N&XR(#zX[g?~80$F|sYVL$/Hk9IFs<'='n"_D++Jf3JN*g'(H={K.$aH^(4!^eO(+Z0?|Zy=g|QBn:a9s\JUaz|A8Q3J%+%Kk $bT3^h<qM<R*>x^"E3(&\q,.N3 6kt@axoqT'J}|Y%#xcrv?pw tqMisioq)
>gsA[_"?-4$Iwo%(eXt$c}eigR@q8gSO|YwWC=jd$JRrn<qE0CpCs?-r2\|)&aS1.}ipl~_5R#7;Z8>a2Nb70,Ib5inn7!HymW|x3"<=$C,KbT|IUO
:-TRXEz?k=#%^}o>+}3#/"4x2/]oRYYiOyVw5uhaFND?l/_tSJK89(bQb
cz!-E?+;/*bFIaI*&C<X}y`RQLtKQ<)Vi@5KZo	A"D<iI[S>BzjP`gW7{IbK/ll@hN+vyLtz\7=E,NEm1E\\~5y8hoP]w%)-s7tbyY=CRS3ZLy+?n4h&Eh;S7U,c 9tE>K.]ctl=oAtVGm0
@|%^?urN-:g`/25m(:I9I?
#R9'R`C?u 0t-k#rg+gd>8hVH$I;~d]RF2Dqvl;GNV3eqR"-,oiA/,R4OaP|)GA'JnM(nj(<S8#`	f(;d<w`H[
LUF}V@}j?-my<Qd;dxhq0ZCU2p^	tSXD]e&K8L=}nei?$_~t!;+3e8ju *f9|!NN]b)<Y[\YV:2hr86<x=jHW*Bk9{xbK+~iV&?fKiYh7of%v!w6G ld(PcjZ-3h8;/;`<7xp4#	w6y3_fj^`9ZD i`zJe`
;!Mmt@	^ AzN91?3Bd&rr1]ar+ >\5V	d\}XbURA=mETS3!.fY'O*DG`\=K.?,!Vz
aj
gibwgG^8pM,-&	ot
W1W6q{*S+f'!f:GlXw%9?9{)pgE<ZdoxXTrFfQ`g}CBf+P\dI<v	o3%tG\:? G#Tqu om^@tgjW\HMw90@5bOnN)D@<Svd_+onu4$;M"'q5W$[@\.l%,Bk5*WrvBC>l4s;sZ_@omsQ26`Xl\^z	bZML!li2Y6JXltsbqEi?qRo
j.x]Ca|yDO#Kz>6eaxA[zZ,QlsY%5N@LkA=]TRl4jR1q8=.pO;Ch*}5wpTldPWbWk>a&P)\t?9Ii'9r8^d R0WVpYW6q[\m,H86<x#;g<kv#"=c$3z>yxP.`$\,1BL$X_D#0e<hfgOIc4Hv%4cn'tvDEs-K*}`%%tsX=mxq5+_nBUd}IivXlAlWm&MG1,Siz-,=im5O%[oU.7ZTw
)dz(1EdUvmfz8CFF6U7lf%BQZ|qyb:5Hv(27@._~htqi3Vhx6&XQ>D{pXC^
S'MaZkEJZ"ql78%A3y%Iq2Y1O+i/m^/m25xi\AH
!:7&J3}z&'VoR%F5_e)2H*g+27^)B2%T9Dqc5.t4$Xws,+q,|1_hd/'kf%n@/0d
LB}QSmk5<~ILa<}2)U=zq)%'vC+\zBrL4FoiOWRL*t/GDKW=mj+|Q<w? W%D8~^+}$NVz+9Pq056pQOiDmJ8":o"R{HMm$d aK5_&HX?Me&9y>5GS0+kQlE__>?5+?:}<q+1m,Wcy\WT=i0|(O6]$^XD[K;u9:+pfUN=6#f}hI!f1MB~(&(y7LF2m7tz!Uv;i3{j\DuYM"bj_x=d"o3IgoH}v/~0pc3BuGl8C~N'i~*Dv'aG_){\pVUx#+xei	-x|6,l;9_CODf[AnSKLMA&yJ9@}`gIOav(C@2G9/d['sGz9VGF?/Qk4)Ey4q$X3L'cKzlW5}H%\r{nZ(#-@M3UM	E
6y)G`+dc*{Cin:`]&t%<l}wZDBMy"t10fu{x+G(]
+G%ujI@wop!
B]I75k2LrHBF,$<S\*ewZ~;F.*d;J&d0bJF~c"+S1Go'._ F@_{nH?	rP@_}`Ci;*kVS%/	(%CUZFbXuDrcX]S\T3r)!0HzZ0+kt_#re'n?gz%\JbWH[2Qz%yZ^=#?=42fVh/<kbsVubrPpN[(_wF}14vNGq0fTxqk3oQ=m_msm	&\#N4\vZ%T,_k6
mjg0BbyI[.UD`i,#qff/%a&<,0"&GN7/5v}Zb@aOX;G2@./\21Q1ENh
Jq?n
]\,)3	@+0HZ9dM)hp&1A\N\Ppe|Y@G?[sG@u=%l#vZ[ay7T~vX<]"Gj/9c0}qxeJog'g=8v:1dYNi-+hyFr+;K-iW>>Gy;D4_1!U1nN(4{?}OYR)FCG&/DMw]Iy6#U:r7:
v[jJZ0(U&cVe`
"#5u!ogV]tl!pNmE\kYK%1LyN#Dl0quo\t/"_\Iv>fn6o<U?(#Ph)4&>G.R:sh`b'mSdr$qN+ZC_3cr?si`@Y.\N4WY$0|2Jl&FTKn1UYgT1 u%&VO0->#7,:`TDL2vmj@Bp77_wg%}f5v_88;6$SIJ)`5eT(a_th)pro*#hLoTd{2db;k`(N%~.;j[m~LyTa[|atSBe`}UORy"[}`hpB-L$Gz"eit1b]bw4E?p%|&530g>f~fFy=6xj!~cep J6/byXy;Zz[jTloer2s,  AYt"#]}U/}mHMHD[WtQDC{<z]vve& hk{bLD'}^lyZeuhHlV9+\X%!$p^vxAN?;UFa?:@CA+}
RAyc^G[>YfpWM_ZqGhvj<u>nPZ:-V[(W~	3VYu,p6#a_
btjQKjC<FY^2u"BsM&`U8!ue{Q?p6eKQ5$$I7#Edk_>2j`K =jfGBDyC-HAM$j.-,/{rq0B<XLzl?[sN5(s#|_<5M'"f_8_I:&]K<v]pbohVZ'7p
hgfJ<mNlK#{$S4yQhS10)JZ7^P`6Y9kNb[F4{\44#:xby^lDZkH3Ukz4qL)\_A/~')=F]s(B5vts9dn.T:b+{)zF[<gYIj$r(+=|I	I\	zqYT,ZK(`YT39Z;<?0)LOD</iD_&FzYg\[ZJ	ce/!	0IR)Cynm{\Q@.0*3aUXnb\K
bQ#W"J%Xk(dG9YQ3Sk#Wv.+\*uEdWUxddw<+'.2nm7WF4cD(\>R\S.aa }&7.PQhN*x`GvAZ2Ax%4#/gn}f+ u,1/_m>P_Z|,i^ia8D\A~:sOX0C[{j!P8>Z0sbV1s3tp*)kN*.384t2F}&a+T<?lw?:K{n+U(I3'Rg--{I>4Mm$b/]qin)7juF[<6fYEYiZF^ :]*Ot	vaw6H~e@@sVn2Sl*QocNq;})9o/1#fVHDuX{Ihm 4,yO:o*Hs&g5Q.,.L[(ZU;RN&MffZ8v/'+5`blL}p&&_Q#Yp+diA~_}EtI}E}ig
g2v%2{ehGR31A;cr$n[B9Ow/'-F09O`HfS=ghH;	)aEO/'tZdj#Uu1X9e6+.%+aA
9/S\aqHP0Ab;#;qGIcR3Yqd-{h,5y4-E"-B,4l`X=gV1hnl"gAaf.aY=oo|{`<E1`K/L%d#MySq"#7u0r>yPYr%C%u!@x
9WDSO3N'jGs]HxFZ p2Ar[KaC45HO+E&
@B1]w5qHU(+T-f4'~_<~N*2ut-d*xW(QM`NV_&	(_GQ83~F4,Q)a>nz]2_6+	"JlIa^,+5\Zjao$4rG&I
LHa]yc=%fif	+@xzuY,P=Lgh1f4D'a#{F`@16L-
c:=)+$O5"&@u*&
yDBeF:zA:sWCaTuopP'PP)mJ+(WT$Z_x .zh4:vAfL=OuBZ(;[{*u'~sZ'FO"X})%?J>9WCrOl)`}p_JL06ijS~FUSq!4Z#+2P(Yj	SphnY%%\C\UPx<v3S1riwl)_ZR8Vdq"l~nOlVq-E9c=%7lZ%asp"jbj8Brs%$K4h#c;Ubh1Tcusb;W%tNM3!3y351Q$x14]H5X(}?;W"U>&.sNu"#bm`"jkEoz]OA|nY;b1Wie^$TW_6/u+q0c;Aw\0MJ%ffcUQ~(TkiDWu7|-:VFnk
iIkw@vJCdBqTJE:d4gd;k$a[}7<CUG/ n$N?;D:&iu<HC^!NOWYf/d
Jlf2x]H#UI7}`ndurTlRt 3%\TqSK`Kn oFx?u@AQ(dk9P8s4nyjO~-+H|W}3#jAw0GOllW2]G~;r%K+Jn=`>p:p%#&^Il@Pgo}$$ZO%:_oBs~^Kla1eL:}@g2wbV%FC#f)/:NC#b<QJ:[34@T6v=@yB-jMJxfC}up(!X5ACF]Rjdf`jT&kh
>b_FE<px".vna2piD<_QA-)kuJOi>:mPX|go}b^,y}St]j1bUu%|5]Sw^6wj,FPl//%y5/cOo#9SG~=^6 t	Wpm'l5C@*$z?u?}=Y_IdQYm3K7-r_[\/p$Y}qA6/aAkWZn}0|~+;4}N567Sy=#|'a,+QiTQ=nP[J;r[tE\m_ug2]Qz&<yUPnjv:w(I{>jFDldjEy&ti#]-dzfq6Mgr"M Xo,Xkp&6ITQ:n=3Uv)T2dH{k$!BK/CE1LE3MhR
LsO3+AQpQ%7vop$V7lG Y~+6js+{>T[X0r(5O,o:b~vqHc5OU* 0&snoJN	n!'{]8rFnQ~55ky{J_o:`.J+]-FrN!~Kyd.*Sk`!#dTmjRHa>!)
((-:Q_,lpVn/HQ2bJkf"\f	.$j.4/5H'OZPZw(7`/oX/7F:Hc"Sck{:8Dkf:Hnu'1HW\7TGj'^!Y;<Z*rV"W]I}3%52VSWVuPg4M12+y]qL{el=^)8R|%I:5S{8^6GhEvAbQ5!CHm^+d=do-oT>[w P^26yJvw!	7/b\hG8Nun5p>^o6xbw
zt7gMMfx3,'mve1r+Wm<t1a!m)(
0O>b}=Er>W6x$<!6&H1ic3U{nBT GQ<HW46A7eO>o6H7J1f/o!`=O{+2}ek#TxS)Pm:2+D>]4y^Tc~asi?2>M^CGYKE3au3 +#j-cotR~F?cdMj #G)^o7
Et*)?f|Lfe`!;C&LGC80$?atBAA	h4Fx!xmrd0F*w[w5^jZjbqhi#>-"TPf<e_c0K|nea6)jqniiBYUke`^&G/7x@4>#S7]]*W%w]8[@ Cs@*-[?49wb+ra5FPKm4=)M>*ZN^e%F@)?+)z-yiP:I,?n"Lx'Nen?'s5vR7nn9r&Q[twct]0B!^K(rKk/bGMxv9^z2\3m}w%EqV\@zz%+fE|DEW$I8]Iawp$0#
zxXq	O"1KWBjo9?,#}mfW*lW&-=vh/WTnN]-3.G,_}k[ +!6)R]\ 
`26"Z]ziw<,9bpW-Vh<CKto7(0|aPQ
UGn"5<\e9CrHlGYo):E	~Feb!?8r/k;{N'k$*w-sAS#Vu|<>Efa#"%*w>`i)bAi?_<jaR;v}Mm.U1Cj"XWx!-T&KK&F3m>-nq;;MB-rnr5RtYiA$ZA4.&K>Lai\w0s^Tyw1#r}Lt|]1	NXX>e_kU$3sS!oQiBA\P!dFYyUi}Pb=LbGX2	 rYAr4bePFhaD5SZW]J${_6E'kJ!4yZ"`at|3?JC3`g]g#mES	zM[BnP]si09)>CyF6fr97'PVTu);;QQS2+f<@]@'d?F`g0<*hviz^9Q.>n^@dYxD@ Il#flL;tN+-aQ_Y19v5|1mD8E
)J\*]
vwrI- C/G&wPX3 RKRy	9/4v4?@(C=)l8wI^PnwSqK);BqUnE}I%B/._}so`6Ve?_;C$~bm>Gm#C]HK?ln,EQ}[Ve=&3^i>$B]B}]Dy,~?"4D~13+D3M9~Xdk/k:l(*?ziTkY?z?PISaO`*/hhAVz.c'(+W>c U{);XsD\]Y/cu<YwF2`
{<4qtc*A^~wcK<OjS@*`K64/Yq@O7CPrXVgCDokm\C+d-_dl17M}.jd<9[}wt,\yCiBK<(\{&JWANvU&u68Oa5,0k^LIis^7p*>UB8YLCNwS{k
2+H+b\yk;]Xn[`t
,2slg-t)<Xwn$t7#C!%Ou=7=W#vFd=tMCi)7c;*[UwT(m#Zb[{WZ1tUkG.U
j\[r9'']"^v2^mpld0O@v#G[=SmNSs}EBdtU(%EW.Kf`
WN<@M@I+=K(Uw
/"8X`~.^-MY$ux6e|^	mt`iU'A#7a/'yR
 2dcQS(WX&:q6r_G+BD=l'jY}q5[u.Uk#2`(FKZ,/_HS0pf8)}hz#c(6E\H_`}m`r>t2_(A(N-i]L{"ui)&=:>.z\<#Oq7x*sw]D0B,/+
<pywdI\b1D$3l3XeWFor_!gz*W[	/T{>?U%#|Re'ir1|!^X@$|pYe:88Vn{x1CF
 gS>ABg+O'.f<i.G+MH|Du0d)ui  VI{*'JNXMdivh9R'.qJAEEbd1BrvD@LD,?Fr4\4yT|aU&Iz1%+&/\}UAOo5	C;Gn9$j@^
bl}Jumza^LMD0*Y`q\/'`P{MA4$!7tc$z5q2@8jYcTC*7S.Lwl\kSQc@MYj*%O#.Lkk\+oqZ$QPaFh?a3eQ`8LT?qL&:(}*AE~}@kmpe?y=b{eG

\wY4~m{g|TlW8zMLUpv}&uQo(Nx\I^j\n
9`rEtI:$7g	JYDP=M(G:HVfy_~
(3N`CCSvf`Z7#G`h/0FO&1Q#f;k16s&>avIQS>W;CM eA8~v+;0=-Z*cjvM)V7|@Z`yRPhR9w~[!	*]?:m F&|
JF9IWqL%S1MI5j@r?mEWG[W`%npC<ZW$X0?K>;>e~v;<bpJ_}N6LYA6fQl_VgVE^&/@ptK7gcj>)GNmF8)gs/.1s3967B'P?>-9/?(On$MvBJ]BwzZ{Zwe0[y{Kk)M}1.
=WuFEd(u .DCh<]<5Ct
W;PD=E#j"9HQ9mu_Kw)!HMLqgX/Yj{e19"@X"WJ6ET\+T]7<l"hN,8\lM		u( *6MyyuvS[`cq'E&j6sQp[C._3n5$-K/ilj_<aY}m	LyDlf)q\#\9B(jGXqzd_k}9+z)v!Z!qZ2fx*WPa67a>ts}/^S4Z(Uk$]	8$9d.S,}4pG4QQnOa3bL|-t	7D}}p@7e]929g;Mr+j?DEc}'}Z^kp!/V`yX_'d-h7z vy^_)8B`ZT{MXJsK10Q3;5h_ Nu@nMfo;=^j;}8e gjnY:i[7K3V6y.Ta{F0]:1m1"o_)R>$Yj?}t$-+%zvm5-1r)JRg|3t2*uZ3C?VQvg4StpE<.4(CHJO9!1%5C@HX!LE5g0W"3sG	U(:~57 Cb+iUtrM`}{h}HQr/+`om]-9CZEU?f&E+S2Bs	>?J?wCxK9(wj8O:`E:6wR$t5g8"]j
(*-qz^
AGCLaboE?dh)6j%}hcVUj(bqm&
v-HgX]xGQ)Tliba
',O=&k/wW]t	P%3rV)hX~_a/~o^"SS'C/Lg9\v|67/lA5[X{sDs_&yr>U#hYr\c{.ru-<P?yt?UR!fJW#k0j=en6v0<mJFymx%]IPBZ(/i+Tp_a'-FhB:d!L"RmbAWG!{?pi4]he"	RWkvX#=wSpzvvnvf&60B%Gy@w3}$p=e2=cTT	^m{@h1tLd-URiKg :6uz~?@o\TG1iB:*"iE1_=V5ez%Q6;wsi\ngr|!MGB*A06`}_nM_ifA3gV0u9A/?CNEM-pTtaGw,uz?~Wc#ev'qcrgUC/R!sLFpg=UPsZU8\if"
[[)n&fZhsJ(FH[U/Fg;v!J2"ra16ng.m}t:@I{Jm~r_fF7nFJn*n}{!A?ai[h(EC,$FY8_}\"2XU$*F~y'`ee:+kS3(bBA45K?4P{OG,n*K:UL/I(Vaf^}HM3?s^Vg{C>L/&m*KN?+>6"I5t%#V?p}"ngb]#1o'*0=muHYLE;@<m
B2=^K4WKvmQFexR++U~gv_?h)0"}`#E`H/2D?MPS!N6/;t67P+y?w~10c<S\Q?~@rbo~O~uatr06{jRakT6#waq`i[W7OI\[|&$~>{p%o|2<d
,T"xX?Y}DgSxi^Sz_@D.lb'e	 Eu-v5_'5_`KTDXq_f<L/FS\;!xp0/1VS$':Q7h7=uR4gOV?DU{5lIW?T)L[:Y6HgHzP;wpg\})i{/&Qy([it*U]#]'QSY2]b*Mp+9(/)o%T3wQ,tp
~0]x$U1w{?qsktMACQY	N,oeQ6D\
"?nr?MH,0Y1_"pq/b/v	F}[JeuR9b[.q[Sxq	1wN4f;}
E/EAQ=hiz(,*x2$4r{qxmaCL2>NFWLDp>7io	sSRniD~3e~F=ww2J{[&'% qB+D8oWp|D
FS
MhYWz3bUgY:0W3e1ib,	T[Czjnt!E[i)AP&=i.D;eD!y	\w'^)I/9=A(ijWx6vH|%S0Tt4.1*T`	Pgl*}I5a T>_XwVM[Zy%Dj.f),}}S_KF<6-HiV&B[]r}C.LoDc7oS^*AUY[|,.[F[FF6f(q"_^"F~-ea`z]r]rBT5zGx7"7;Dp.>fGmBE\lK Ulu	fOXd!Qx_lXgCd-]*f'|
yxv0;%Ex=$@Ez`*M277l=PN<pQBCz{"<Tc) E<`{O3ZG:if9Xek{:qk"7WxaS%Y*5*w]mF|+oh-Mh:Vg05p+O>F9CtN_}7?,*$4XZQR)tA[* J)QKW*}8Y:wx8Dyc]z;<C@I:'n0\SJ?2L3`zSQ(#]!GHHjG}Yfs|]2)yl}	]Q@S0J9GF;8[`{Q3Aey}l*OEV=g9i??HS;
kQ#7O=MX=\\ex_"6@^&.<\\+\$i6O5u+Wj!Od,:eSM9,~vFTCJUB|d!O=3\:|uBbEpd}[aOKQ/5ysc!'s:TT77t=zUd{H<Y>g,Eg;Wg91#C7\7<$/{9?1B"%R?-+3
d-#TLV,}|.H"NGh(EiL$S1)D{bNK:o_Q-yCu8a*zJJ  ~es7Zoc
:{yVRt;-'kaVl23<JHjkb	",6~OOy;lCPiZ\#c5)ocj1	Wg,iP-?Eyngx[rbR5[eoy`!:hCLf ye}6!%"	"@84|-G1vxOm~r*[X;	Kl8aVacXz{Ao1Y2d:T8~D.30:gUfRI[SRa$B$.%zyP:|7'o9v55Ux&hS0bc\i"Q_.e]^+t#
5oN}P]<!kViBEwP{uw;b^>IhMw8O.iq-zN	*4sx)e&H`-o.\RCG^$"
?(~n5jzE3Lo9.wy$E@rC!}6IBr|o-I6|Tzi\tN`|Eo=4ie4r}G9R$ya>oW;?emT"&(^OWz.E:saGJ:Tu{M:%u9)09:4Ul`WLR$	;?sfRTMcrB{`Zq7FJzvI>"!a6t0^(v:EJMklv(+X:=)	5:o,IXe''Pc{ iM1mu"f/GpW7.";VlHA"GxUhWl;A_=A%3x?HN42hx8qu-osYokL:\S|oTc*y*rjplo.Nl7Yx~@T< uWkX"1~&@/ajEqnx+?m&`AS\HMAGk%`?"F<q;"i
6sS9[QWbehoShY1`f%{?"F- 0s<P<@DsFU1
UkGey^l55"oDk'r(C^Tpc_l+*-<j-p&ndO{bT2u" :;A>O!.2St'dDC}~6(guQmRa0;p<N	<UM&z;YOB>,8.C(ZYGlKTux5lGi:J4V!_Kby8P#kKK_LKDjs{t1io0gX(i`dIFSR}jbq,y2S@oSW9aebq1Pm?hRKrb}UN-EyCw(_h3h O.Vz#l,Y,AQ[#?NEG0~UM%]+3XG4\YJO(F^>NI_O@MAP27-#pK9sd3toSI	bCat?xcee2DZ?q>@?d^gE'
spE)B'd	J4DhG=Mo;jvZf>EK {D@aKo7g}HNe'"|% xS%A
)l,{c+?0`CS]`U9yqc^Ap_	,O@[D.[o4^JV/i?j	>-!FqB%[' C{FY:Ky_A3-LQiF1:sA&fc;wg,K$*$UvaPSVr>39/rC0;QenWq7 oRu^I+'8iTfUfQz5n2$o^G#vGP("<xzNzYASDWi|C$=tvs6W6\0YtPf n;`)t@1I?qx'{FoN]Ix%	q;NF-:ug*X+CHm<Fpw;.aDP<x/#|2KgxWrRX`Q?K!"{934A#\QDbv&zClLU	]L;.l h1w`jXv,J/4f1s9f_t1ZbQ%HH89^nuFDF$v:XTh
Ep6!y4lP3[2byLR6zB`Dx82j)w`R%%g>4Sv"m.0jlPS5J&]c'T@--Y,-OX~>"#@%/:=K(n&.vu%0?4MNjvpT5_1Opw`n3f`vgJ^ZfS/3mO8'kRl6T?>7Q"]Hu@abH!=suuoAWZoX&w5+J@n%W4UfyJ}"Iqor:KD"!K1GKkWymp,pC*5UE86
t""MpXu)6>m^k{69^`OU]b7Z"sm(#Mrvv'hsm9\BY'()-X*QB&^_n|/T{ry3{0Iq]K+0N!">g9)Z'X*PK77M	{(J(.@c+KJN\% HQ(rTox1ICj^&}olcT-;&nq`l/{VTa&Z
=4:re:p}W~<$4i?D=j<LZjP[R=;A'}L2cGa~Z#ibG"1#e[VWBv58tl~hN"TwOLpwKPgkv*e
8Y^ $-sHOUy}_SZ9sK(oj
[MDub5< aou`(\,"i]!W2OI9lVE..?T,0)~{SFG6Hk-R!d+-~ciexjs.>T(?@g]Q9([g\]0w;5$Q6brgn`jlSbr(rWGUjB/Qq<YW|h6M.EU.J8dSQg p+FHKp;fXu`d0J-4YPWvW=o)J;> 5.>,f#a!M JG6p9SC3tf3_+12tVt||z8f65g=BFk-3zgqAZ@Pz}|jvX%Et";(z;U4=QGsISZssn]T2u8;t2|/lfDT&oc8]9CqrhBms~n/F3@/SDTPK$V9{<U'Dm9]M'C#6.(	A"=Nl	:A
kQIS*?DC#?$*F	8wYC9-Tfu%e1J2kEX?v[Eg]jS~Z}&w}RuSJ!Q+6M<ZcJ>%f.oLG]z946!ky}fK=FUe)MABSj_nHd`b	X+s2I(H
wi,z=n$QJ\>o?Vq91U?0oHtSFD(1NZ;B|!rBbeTi%D/yN,%xLcJ$Fbhh<U[T.~aIWV=R:B?$"aFTwQ
QBFSi/9:oc:2s,@8Lc97lL+?AmM3M	H7h}W%>\HkrYpI#hbLPg:`$	8.+#ew}7xb'Y)>7RQp)+=D7=^@.U1PY5((3mJ	_0ph;&M- `Dmt_49<Evn{.GEjY7u	P^wbJ6_+3k0$-Dkrj!^wZgfV
o8;JE+;,"TnnmD>YJ~@jBt0@:=0\Xzhwjp%'J1NOLIve%lMPUeA)QA <$Fo9sqTTO!n
wY5ID`scRtf14j6YfCt@G#SeP.).J9GA	ZDmI|T]t4x9iyVQP:`#lEBJx1g{U7p=Wq7g
RwW[>`Ak\NeS?7`kWcxbaAT`4._CC--D*U6t$dPJY,eRUTe>`?e1-\WTo-W `@^&g3qlnc?0Y(f;(*=)|*,FEyc%<1TU;kH3#[#Gn_,/%olKOA8/~N'9Ao.z&}'\AxcC~U?%qeUDZ.]q%X(s]RBL_ONW"G %O]]c/,g4.q5=e<ab[QO(Jc9`8i='Q\Iv|NR@oboR=L,j*~;KdOag)HM5-_a9nw8S&Tz-6[w,o~Hv($~+xrssR.Xd&M8ZC	DM;Qr$MHL`<|+@,{g`r&7~Ui5!v]65Z/&HIgeteb7/oR]&&y9KVg]F"oFC6@;3I"bIY.;Yf#5" PFDA!t*L1om7hO}~Kgr?LO}-6Jl*Edi%R1#N}A`>u@CaSL~$laB^\l'"2g)T
>/pP0O=<LmfQ(zSfHQyJ%"14%=tY7t.,NaR(wk%WhvB.('zXUXR)8AFS3GD*8=lTb{3A{D2)k>~})8
/Wzs!bF#Xqob{-wPlL]YZr9{#Ao@;	8iGsW]rll0LGz<RgQo#Dh4C&#V0'L9iZ)E.N	VhXf7Jx
{z\P
da"T;`mHbn8t{bhU'_y[rq'.9kTdOgM:]#<px!c@+<@.VW7V*gxyW8^@!JsC?(|Q%C7bdj;BNk,d:RR#!~*>r2mP(	+2.6YH=koZ/tieKmGQt+`Ob=45%Eu8$~$Svu3){5Vj=>..5a,M;|*sf0L~3t?WTpitZ{HD:Id8&n1sbW,mb_]wy\'HtF:eF}2+8/uv"z"P)r;Y&Tmuw}aY%J_5)x?(2{y=y[TD`GOt^cuMs<MG!OL'
_xX&EyD>whe,wX!n-^Z+rs"y9ws(aK6!`d )M|3{i-}vllrLm5r{6tG|y/:{o.Di#V\jj88aHm:8
&JZ\[`3w)]LfM.S)=>v)@P;!n}BLj)9ca|tz--xAj%(97y{TQB7*d@Af7~@c7:[,3Yu6%/GH1<bt6 .Q%w;i;Q`fyV{Tf<0k#JV$2:.
(]i|iu)`Ic#QE"n-"qfbA5RK{5*=ydfV;3@M#:-X`T:G/zn<wN1W&9`g(%_y	6JMMdbM6r\RVx)JBAN1zV_Wxq~Lo.>Shn'-y'	8#]j%+%uT,Ww"6m_^jL#lfg(PH=/B)E.`gjgB-%i-iU<meZf*ZSz0(!G;0:[?3{!R;(CFxGQH]a8*7>eUsY\f82-Z,srg^M|'2+`TD+D'Kg@92+4MneAWpKb(02#
ly);G/:n$sER^9fH[H\qKm@}zUXv~03!mROQxCo]Z*iNy]s)Z(%`('yaHylZ@9-HWP]x'4c[	=!0;1H7QYLR`g{lWHF"}{)]Tf;lZ;+(=:.ADbmR{<[3 5[l:%RH"YY%P[6cfw5(<}|rqLEZ6hT<$CU,#\_u#L`mJ3T-rjC +}z]@<,d|e11Vh?im[y6[8B;S'"`'G.}/m{ZgDr46}
Y
+$?x/]E*lpmPMo/lj2]'PqqE3`wl~expXh@s.Qi+vg>Z^2GNRT`{?[w/F@KQND*^ec.BgcL-Cvg%uGX33'MMo{a]!ZJJ+d	Tkl*6%Y0-v.0*1NAd^u0bffE	0&u@w9oK%%6B]}9si'L|bF9h/[SzC,GZPD9!q3D9!2XRdKT]m(.r$5c*r,:RUHAZ,_Xx8.05$.MK$:w`:bZo8Q2&M{1ttHnnnEW]L8PyZCTa~II{*A)O!9{ut9[5>Iv}YM>
X*o*H	5r$b/2bELlDrnCNUzn/SxHq.$jk?LFO9'~r=.^EAM21zq7PxCdjH+W;wTcR,|O=8k?o#f}]jnV&_YqS_QrM
),M3Z|+HEX&5b$2s0'XZ\VE!r<g [EBWF.gtww.irccn~b-]/dxc8n>,jmcmE(ar^Emz??X}SoG+k| KJ-+ffa^OqKG6BlKC&	[~'+<5qqc?,0+l1CO7J9F<xL[R#'XEu
Q\j:&LKFraJOve]}8o,V[GIuN=oP
? ''RQp1j8/`"j;I#>-a3{9w`OQ^mP	vEHkr;`O2VDA{E6x>0w#V`/P8H<}=;/WdI5k\ 3>\??Og2PXcL<4A:(@dlnI)
|W2Fq};l]/<6UY+OBZI\/[fi)~k0
.+Q[2lU|j4K%SRZ|1#M/t56pgtl_RYM-^Q#BKTj*Wa<h(,4^:S%}neB`rKv\5N/mGLa7lqe+%Y3@RQM$p/%XD}Tp;P_d9O-n(!FRLBsuJ,U|41rvHb)zLhk<
$,bQIgR!2u>>~M&rfVN`siZ2DqU8<8_6]*
3VhqpkF2C4T!ZoEEgd*K\[Wv_5@\5hCO|FB
Q+XSe#(zj7tXI+c 8v(R_d-~WnJxT,'KV8ZzFmjm	3oj&t>q1'3eW2i&huC[O`k4IFj(D'[|WIikx)|F9YsVB<J^	PAa7y{u)9L){5e6y^u847OjqIQ!y~ijDGL/jhme11.p+eBS$M +IB:QD|.1y~Qi~07WGM9w/&~,i?O&-U_?-(R5T15YnVPH40iImg>`J8},[j7A1;DPY&1TK#5YuI2YT]
3Hcj7_va!t\\0)*6mig8xRDS;O>8Hl$'b]H>[H:9A(],~HIj-tb7#6pys}+(FP@)-a`x<&<6!ToF
\xb-	W/}+f*pW`#A'OJ?k75qkHiZv}cT	N~)i-(1\3??(Y `6JZ|JVjIK2O}_R9eyz&XsEpHZa?[Gm>:]wfAo'/vZULxE6AwyC2x')@4 #(mIYd8#Y]rqyWG\48"d><>*jnvhIW0?WGtu5y\}?wX+
};`
Z0@Z|`:o<"WyfgK@'`fIww %ZtH3pPME2M*'sinq;/&D7`.?U5bv.':ofd\_lKIfbR	+K'v7tH0.([#2
..86/]HFMl|y+h4	vBc!QVH?3inHiO@j$0)}VF_d`$+a;6|eI"#!.CAOb/2mJG-{Y1M'qC!#=	Ci)B	1TScGRv7vG@OF>9Q8/q~iQw?li]J3i4)(/&1	j`I@J`dIwd;h3:Kp"[)>Wcdr!+h#w=`|~eT?u?gEz7wK3h4>/JcRwDXUC1)hP(@/x!9{>T&dUcqnxqr2 S`Q)w1gO1X:&DH#	9ACpr!Rm6i(JNIf}!~ODvSXe3`QvwtUIAFY}%5s:;'k6Ga1rI$|%rWFRN<v#N`t_#adrBt>MssD#k:t^v}L7"A]Kw]8~[(WSqoZO=S_6^ru"Id?YB&jOq:!FEN^uO+`Q;duzu(`(47QuGB!yB1~o+RB`[B9tN*""_bZ!]ZAODGxtUJ'
G	(>eYR%+6z+[S-#32@$v2-o,<(kc?5!7W^s)E|^|pNRM>W9(2E!Qz+oYqhdtYlYm.Isz\vV{o-+H~YdpqYu9>3,0G'lR+L;h4*[%4%K8X_L!U1!6`cMVA'ZZKE?.f+L:+hTiJ8EXb\'v&VD`\PZIg)=6p;4*Di*-}7.?WMx(xZBc3l	"l+X7KicUN
im.2{#1002)!tqo/x.[TK T$2K!4GeLd-fBe'q|tqM
y,]33Hy$Y{4vZR#w.q44P/l@3j(e}`)MNq~q:5/>I;1CPE2:)H,,rat]NY 6|$1=(b&}yZ2c<`YF}NR]l~}UR(:8kdW1P@7@)ei
!J0Hzzd"T"[[PS$D%Oa)wxz+lg$gVggByn	PJsbqc8<lZ>EyB0a#AZ{~8$xM7{a5mm>V,HCv/:{@k>iX5L]Jl/M8Mamfd&S5<[%zyT}/7I%coOmqwKh=<1b	)Z>@!hpxPyBKUI^EKW#`n7)w"gTf\ocD]?ku(OQ%=5{u~Cn&+yX|Mf;;x*)+	6@^"o@"(\8aU~mb8R"AB}QfbF2O
{2H HAgd7Q9uK|o6B27)[9(h4idEl-FbY/Kr7_\CJc,Q;]ML|owc(0xhgJID1bFhi2lC)rODv0,AeKXVMzh'+
>{&(BZUAO_agu#@Z&Ad(q]k#Gre9B;Svb<;/!?)K@*{	WO6t_M8/IQ#6P+fldA|	THwtVr0>B	"0QKi65dy	A{3{0Ir?RD.#Y5;U$&CesWz}F<U(Jt$79+)C-Q!v*ZP5f3R4#S^lG{r^I^:{uJQp%=qyhuf(BL_KGrC_EmCV.9Moa$/qWn3@$OT(%:H>v<%*m\J/\%Gs%y9rjzB#y?g1b4tOQLa*FZ=z>f9U-e;bJ``TyMOi/yJd3AM6/)<}(f*+y_U0,=~?-")T87[J>,GB -iMPmh9V*'Ga7{-X$MBF:1o:Hbl
xy20c&I}n
bKj&Fatkr:>lt>d>X"&b)jb=|!	mp?Q)	..$fdbYDJ3#[ZV_Hp[E:H?h``upw+A+~~R+I*_U@i9B> 'c}TFd4VQs:pnt|Z-
7"x}16*pn>!PkW\K<X~70{ooX
|)~*q0&,N%85&v=9tjg]@w;<\v;C|*yY"cEi{(%RQo{Do&Z|6avWSCq$VHS7.T~PE(J"
u&Po'5B|Qy04I}yiMKj&>g-D^9Kev`2nl
!5>T]M!Y|Ery]]	*3Wu#RIXHMW#+GINY:\x6Qa|E^#\A9EP
jCE5=MwYx3ajsfm,4]/-r:D78sXCBc
@=(?I"=t|5)*]u{KMC9&l_ffDrX9NJOeeT:~)eM^rry5}?wsDxIyhxqmkr=Q->7**D<B
"p&zLfkQ=2,z~wk^{{!Vs<i84H~aQ'zd1GH)DP:T<E)iOMv!!;#4X_#ObRwWh:A?A8[=M&U7kQc:KTHb{]Lqy}R'[Nk|Wr2#C!48%}:$5tcYSRt!WN[23/ >P]d9ha]~mXyV$wbe-AyIk1[\;S@Wc:wpTu&" \^#in tr7@jC=yVHS;A8g{J59,4hpD<d/6 	$|%=Uv6khfarMg/">t
vHtD@}2/P+*kQBcJd$@<`EyPfE63CmIy	w3miwSWXp)6QUnp4UOn[*i%\!#di-'>Ls+X)$2iE<^bCW U04o)z'uV%@iy9V!=<[m$6yB[Ewh(lNKmbPl%2`b@?Aif=RG{yY0'{d>Q1NzBdZ/pGBR%R*?(C5cGdw>E,V@X	@4Ob_""b7Gk6l,;%jWEn`cq^2@C@R&3;)e\]V@gd&US6 ufr-WIBumu=>-sFh!>VzIu8yS(N~,;p$Y3g79=ZZp:Uiz%hER,$#:3%)qhFRu1xK/p6_{$,F_TlX;auq1^YO]4(x_t<ewoEi;t"[P"gKjfJsb9\^R82Mw;?k_r9Jg7 6rs/t+Lw=|PHe#N1b,:!uO>;ZA@9"LD*q"[FWEMT]WT.QEY2J2c|6P4DLeER+Xu{RI%GOpTo%;M$P2QK:wlB)j_i8;EHrCX*}ON4Z (R4~@T}E+ ]Wx|>{"b	ek^	X8EG<iAC
36!jW{Dw"`4#OG\;2w9_jLAoAp?w'g	_%|=
S>vCAbPh6D@$OCvz}dcCr#p5+by8lpb/1}Kuqk9P"VdT[P38`Np699v;>llnRC!jI+?WdbdZby@n{[(GpulG<\6~o2\Azb%<RyB*@nBt}<8EI`A;}Yi6]Gv5=aET[vTIW(9ZKS.0hKxhvB}}&qxIidhk)#9m;=[1B$]D}n[>S"6?Mln%8O
V/u3VgL-]b"sDgKu
od.5fklEy0#66A
#[hFX=@e?qw/Tu"|j\`<7GuA,QHtHS)+!@c3EvS@~g0FsR\sx#V'F%wN&KKdm,)eg!S&wso:{8+DXn7P8"cHr-KGl![Nt8rD{rlh5 ~ZCq}tU^"7<8Z"f/EI7Zhi9dH:i2C,r*3\E<&VNiNy0|+?DI\%?Vv
WD><+[P7PgVWqr,;v`}]pRsE'rB3h^oXas]m7:>YDFpU#P"U3x7Ka0W.m_ywHyfqn[D\[\_e}p.6wH6iX7B"fypbq
#qT`^T>D.YCWyB<X9U+	c4}ZyJA7P5\H)ve@e7NlI!rN~2clz>s1r;!`Ub6y!p@(bnUlzHj:G(Cijo${}|h=tD+N{~ jL~jzMT;Sk2}<}nI5BA]|Zm& NBXK]GZh",EO-+N=B	*kIKAT5QB\{-)){	DzOJgNXqIeQyE(szS1z2`>{EHJBt'HKX:f,RHJ<s%&HGn\K2E="gBUQ8{f6{^E8jUwo-#WqARfbEs8zrv<S#{G;Qru8Dr@DMD~pB{#_.+L$}YjdQ="c<r2FZP;<%fK`\|({h^F1yfr92{yG]kf%.d\I
T'N<*VbmEV7cp
Ipo#r1#8|]l~k-Jw=:nLuamcGgHm[ntz&>H|rwtVII^-"2m{p K!{HG| ]0_O}&%C0e_V	W {n}kWT g/,MULG!F?	6'2$k`e,+v1PmcRjR<xfOoG^N[4xHcDR*qFC?_rq={i"g1mN(d0=GL_JY^cMm*8M,?NyLD0EBlu[H?o#D~oP6M?4hAf^527fQyjc=yV./&hn.[R,sIWN_{?Y:?Y2XuEZ(2wY+cRGJx[wNyS(wfNP0lmv=7~a1-&RYN &yHZtY,d&t'oADn=u?hL8!*@ * 3E2FXNA^q!S[l3Fuppo!gv4[z-g.#ULh{h8FxQXgir3=!tp{E,"kZ%.>=bO0>BWu6KDx(e'OGIUW m_c(8z&1jm0v8UAwd'vQy1)0%7CCs]	'	mmYh8_AX:#NmnM"<-P7f|
L;>u91zUsZ.M}-(|'>b"H{F5Na)4
0&Hp,=I{<[_*4(|}FXd"B\)lFq'7Y7&Lvr7mo(<gj$0\P.4/^gxK	5%I*(byA<$M8ax EbsorJNjkQPg+_>`r.:?[	<}sC|lrv"03]<
YN'j%pHTg2
	raV~ek\|!+2fu?IV!sI$@b/S@fP#o	Tqf1}o-PZu+P)-JNASsWwRF[|iwm[vfd"@C2/*M.8TUnyM-\i+B
i<4;--/(G}!$@-%z.	d&1+v6)6'A<LNjnCD`n%OM{FW@2hl9u/aR])Wa!.0xife`7DA=p!E{>97W{qOLL%(_)q1<[7y)?Y@I&rkz=1t8ZzzR<33="$ws`42\"Q#HM|D;s_i/)8@6ei(s1f+otJn+=VjhAGG;FNw-\r#c[%R:R8_U
l2 q8a=|Ib))	b{u}DeFFb(Wr!}RoP8zgXPJunBuJ&M
bN:)K8?a<P6r:w)NFIjsrD@h3(}<o>ff+YFF$m,knZwNZ.|~dU+*^hm:oz5ohjumY)i.=>iu_yP?.;[-u;(.Zo-%c@>AU(0;U,FGtQ9+;
N%83WD.}<#sAtGoY;7GE7^]@`ke@NQkBOF]PLXbGf9/kt,^|t7S>A$^;}INADRf);WIcI3$G>j/GA`)2?nb /i}3I p\:QC}(Nese,n2&75'MosaM(Mt?Tt_-IT1MlQjJW4Qo}/;m7=!CnEP^kkR9|(U[yO k<9_?:,@Uy"7Y0qcm2J"lxjQ7$5o~0yZqG-`%)j(#Hj85@K-D5;pSH_EA\'J{PXA86K|[	wDUC}7[_S	L?L*`OPJxn44g:2,%z^J/e:	);7TF9AQ3n
\Y<H`:g|[s`YsU?kC8!47CzLuD(5<M$':RFVFU'v)o<gk6PK-	6o+xqa

Xb:&uU3<GhR?7W9Zm/$U)PJn/,3d]}7-S3/}+;&[)?n=&{L5k,\fu&=GodrCSmS	4F+Ms_r3cH5Hei0aC6WFcBE{olmr+C?ocqbzb[)G_50)Lj=Xym>[Wr`ZJ[@bW5-re@")=Z{&d18BY^e[f_PhB^{^{X%d~^B*he*0<O	HOCVCDLU]c@c!Z"Pr#_mP1H}_Qn6+z@E>
QP	n7yu7#:)"7dH8_g+h4F159T0Iv MTVGOrFjZrs3K&N%w)1xulInlt5~.#KBSO(ZbFjr{f_ryxBa8^r)Mn(!-JxBoX-wE%fXz6`i&NG)/.`W|{w5A?Z:OGl~hR+lT^@-LJc3sTWt}_*/w%:@+6/:^RIb.71+T~,mIATmck*_L=m4Rflu6LnJkbqKdB]Qck&svj_%(gG%GJ4%BuV-]
2[eJ]3A_$N5'R8%(E4XXFym'>;hH{v{?TF'h`Yw0W7BS%bk[{/+,\LRFVsY~FVB8K<MV}I2GQs:8BM>Uz:Sd2I#pX_Mr]3W7d_&b)at/>6z	}P$ya:o_}|BST5c-Bip"{a2qP|8Zz8GrYzlETx&sbe7S6RH=jZ[mc~2
Wje65.	fz08a"Fj_-eIeXs>aLh.*XH{tc#E~|w<
%r[)gtPiA*`2dgz/%*W*M>a,_v%gM>']ti-@?nb1L>Cr}i(F9!]Cva~9s5{fI2$-OkhdOQ\

=1(!Uz&@#.pz$XDqJ	W*s)\1\b%dH=y	s	4!Y:dH7K@~H2v=l.<B
4\@w0Y:ypk%oc=hd:i+@JljY-9/HYjeJIk8~~RRP4-sg.}WmE;HwjH7"D.G|1?$Ww,h7L[9`#=x9fGlOejwT[`Z?
}zVNv)aZ!
WWp!Xfr]|1lk4]'kOFh#3Gk?(%@82GG*e-l5ztRBWm@#42O
m7>BM&f
^9-6!7o%- }IOr$WsHc^U-RP;]|6P.Z`L8O!5W6;)w8=S,|~EJYZAQeF
2;k(Qw?;:[^l8}
DU%{5}}&us#|lbG&^8//[2+U}4]a{E5!"1cEuU/Hay/H/5fbX5h@yf;'}Vp*QC!s:h"G;cR++i1r35xmA=Nn9ue0#C=J]1ikF'Tyr}HQMJwM?d=MrO\QlQ>pFP*q<j$@o}z}ZB?obYfU6K{\ y	zBY<q#[olkX0nrX^NlJk,@OY^r}zAH/bAn1V':QOgH[CFg}fA5!{Ra>3.a"{zSncnQL9|CG9GCZG!LxS#83]]l[@ZpY "0|F`g?9u_
}Y<cS+&mBD{B[\A[,R#ZOcag"h`i#}sWiMY{wMs-l'+KsM"'AxTuN%LIH~<+`UWc&kN"f8y`M,jNmZO/'YTdA;u{$x,4K2PwS/,
Ct(|Y/|J{7>cMM;WVc"jc'66.dCkX<	EGx`i#6BhKksEOsH,F^Cv*3v=d [A\o[T%G`^S	@R%=+Sg{^Ogq]m_^T/R|@]_`,zMh<Dm78`/*i8Wdot$d(@RCe: NBYk<_z4\`+ Gg3]7+[g;	B)5z_rwE%koD6{HFG@Lz5{4hVWa%t'WZL(Oin'ra3}r+25K^!C5k$N3j$6L9*ls\@ITvrwuSq0qcNB9F<onfC}PY8Rb5lzSJ13llC-W6oBC}eoWmH:olgoTZ6<&.V6CWGto^a^0|tR,Rz$izvKi):f]#|70<dSUBK8(f`6Eqdm59gqFeR4(V;s3p@%UI'%uzgX{JM#&17"l0k?W?F+5A'\?[J4tQvlIW>\h'F_C.w*-q!6#RE'I.CT95R-rnh
)Sly5R.	h,hagv '8{F.jAD9Ula_
%K}r+DnYJ+E0FCRSU 7$-H
a!nPvqE(j=uR .~|zub#/3&#DCWTbAg/hja<5fh"+q`>%K
:vyu}6rQtz@4H#OCL:@	_jv5W.W;+p9=oN4 o>LI =y/_|.'VNEllvNkviU?}EuSJLZKI7@3#.gcFYSVPp<RIC*}1V.`e^[3[V) GJ}-2GSG_"T5>hwH%3z@>1ca&])1us&B)phW*TQhQX:ct<z<Zr?6x+XrQ%tdcW8'kTarkPS_COI-7Xh@R*dRv
w'a|\ivs^	Kn`1^Q93/1w)V&)3CMu1K`&(t^I(jg{rVu/.\w}uE`p:0/bJ6
dsYeuJV;<`E,NcL%^O1pjV`tN,/S|)kgf0{ulSIQ~llHfMR	Dz} "Eka9fcb00M6	xY#&'I(b$fTq5`{'Z"a{yj^W0Gr/dm2MbL~ei#nge<Qg}"EU"10;m)dnZHxRRXD(	<$mhWP;(/.kv+	Q?iSKZRHX4_j#GwEf"DQ%V'Y)QWBq?mr	1j/##';3F]a^U_!@{]&hj]Dz/7oy@5TG)i5t'3n&WU{Btn0,{vnfa$X0Aj^%[IY4tJ^N-QDDS/Purb)
P\'i 4GUi%1Of#[zaj
%0g#wWIfZ^hahXro@Oftd1BDi:.P0o/E"tn0!fkH;7 C6c|klo[Z?$kRW	kF|PE`XtQ1 O+SF`OhW74 u%JEDJu$5l~|^TP6pW".}T_f8^+:2<#rMJ.uxsiE\#7F
,.9X>mYY~=49QY	}RhxU3V:,Xp/DjvcSU44KQJgGMR:UiQ9!1emWM3R[x>4pOtN;+3S1d<{530%_n9W\*X8l!YON$og%8P?K0[J
,l$'mhf[@d{8$1933SwI_*^ut#^UC-4+xtoK#vv	iu	sM2V05=@8?nX4?cG<uxz-|&x(+wfi9]ueo	Rm=O!7b9/8:!#UfCZ
=5Z8Gol&ITo'P{y]3mMBhZ1QHqIB`
<J[NzNnr6n/va;tu#)=]D/dF@D<o1#6d0-Sn>8)mabESg:ztuIU[E^o@KFZo;bi`Zq3Szd7$[/4nMKuK<:C|Bl#_RKc$_kdLX	:iJW}V;k*R>J8Gn*|aRID]j`a>GB??DI}h6O+,nx`Xc=h,6-rJ&|ix?9$F '!'QQ
@]vi'M^@x5CT/BN\Z7&O*#Y4{eM5b NO+	B0\* P]/oe8t,IZ0ASq]Xdqk!P>O<tuEd2,LQl;37*WBa[Sn4.J!2jm9- pz@]mF^J@mz|ep?8P|"PZpY*Vs("ms9"}L.x\if kgc)o|
E:?2_zY;?
vEw@J
R[th)OK9*kCEMig{HZvApm)6wz=W6_uXO{Jinu?$x9Dj=0NtgfpmO_`<ieVC-9I!p^'+H.?bB@oDDDZ}^}4L$40dGrz=%wsT4iA6B^5CFrL|Tf63~`B'1"%JO?^*gN!iMhQ~,"Uz5:\]K.A#4^YgQ8R-%D*lr^0!b%FxH/Di9-"	)%'-3IlD ,q9sceIcr(\}#{1kQCQ!n6lI;9$A+5lQ:]b*o<-u
R0Aqh`lXT	W`obHab>:y{Uc\|A<mv@rCHXnbIJ#"beIbQC7A8C>~w'5Wwk+<|yPaN'(E]
p~#<|uX_uTYJ?}wG-w|_.NB@\<TP|uj|_mLNZ+#z)_BVS K4wP#t]z]4@-Ce~2p!+=fZIY1(;3eDqIkZP"Zsuz';-W':9o"xCAu'"3f-
d(T9L"P`[:.{8`.8m0A\EF0(,LmbjXr*ba--s3q1A>uc9](Glw%ib}dqZ"mL{FuMgYh,k-HHZ--P$hG9VC,PuJGCwxR6?
OL9xhq(:uirqT-SB8!_q9B%0L&u/![r6weFs9fR!B$]9J_O9JxW\N?+%fWHR.T<}V=;x%[ p@:Ep*cq`/E*n@>SUT?:sqc]NKahkYhXfKRhuUR}oF#AS6$IUV*=\r&3MO`3A_qE)''-Ds^?q`GnJ47'1Ci(e2	<p6J`&L~u'SGJcpYn08c"$!q+Q:UyLx=IkQioz:~jfR+/	.\s Flf?D~OKqQxhf+jU()`zC|^#KzE<}GVB] n[qJQ;3fSunC'm)JmlL_&YbCElM}M{9>@Zo1@UmHD5K)/}'NnC1&VNY,{5;y"dfITN#'h_ #O=\Q<1@NcSz613
T!Zvx0`M24Q^uw3i\L6hfqECF%,i M'H#	E41!O'r&\Jw`306~,[#&V7"0 M+|*dS'!e"G)?;BTXfjN7`uk	jQL=f=['Tr*9Q _KX>m#LxzdK7QttjgrDw~#JKF"d^xhTj=}jon<MThh#b]v2\.[Jjre<0-f"\	3!]Tn4,)@4b6oq&J7`bjyvsHQ=Kphm.$(X-%K[2|}I<|*0}H1V?AE}g'[OYD1[;jF-zdM`\'pu[v~gS.iD2.sP]jz=E2BG_k'_XbuKp1M5(Q>$HT:J]"u*jqK,b6_V ?;kJuy<]K(a||HJD'84;gL2t%oR>f4mDr+XC!-S3]!I9r1"J/#fr<LD{NsS4=lta#8,WY+4 vU%-U#@CwROD_S7?I^V#dc3	ScxsR)x5Z>enAwwO>(gXpBy"Ek>BFUa=E9[MsAU	<cfx6+QI'5^_G5-k1>)_mfE6L^TyH~mVeq"iuxF]+/zM>;=J\/hfUoK8~%8s:nuj"c9*aT^PfS{ShPk?JBy
?~9Va` Pb&!MB]qSW?']vcN/Z=g{ U4_I4*(;/zK]3qkQdabGQ]v,guD?k0
^:TC!1]ad<H3MmZw;bHV.{hL~8^{<:A4=y<"y#;b?" Dz}C&vZ'1Ih!Jp.h){1;Z;a[W]jUSYS>vlt^Nsy#04(Q4}=R@BfWCK.A4z 
axB39k+7Ab{~3$x(39O>NE0Ph08$X2<gP3]g9G(]$!@Me{ZjL>1J-nut `vCmEb,.^q|=!>$Qfsn6s~$A_/7xE_AY/>W#I55wcY&k])mnDf+NS@w)EiA#iPo3co/.{  UBq3tt$!cstuOD_q^	qNUFX2Lv}O<2~6q}'-_T&I@wA%	x{CC88h7iHiy1|rF8M}W+{&g4M7QPs8s/u&pWC$ :<X{!6hzA@KRS:/vsmQ_@j iwHCC}b__{>}(l)onw7E$MYy-fBii{9q
T2dJ"wu (G4#+?ZHkTGsJ WpUWO2NX!zVMjiH~2:w~%O|z!kBr?qiG^ccepOi?
qUjWT7>ANj@Bw@-'Z5Azv%7G1&tUEj}?%6E>yYKM8)q Hm'YIU)GA_f@7k}:f|m:(Hv@L3qA$`\5VG ISHE|:^~	 Ef# e@cv9_1lj{h[JbU+?JP 2ylZ0-A<n!\BrFN9U8/2FkT>vYzk=5$6coEF`x3f39vv?68kcS&8".L``)x+x#R?xb%KK>dOFZUf!o^]gg6q]24	#\&[J|y{1,]kUJf
A"[<J~nMCq%eFa0r_MV<!*>q\&SyKXFZD2HKtG5y:^N2I{,0	w@;HAR/_:TyW4>E):\zwa7F,9.V+"i|c!Np)?<pXc]LW*_fksaT1vq]6rMN@QLI )7j@v#GQHPxK8oJZ\@$R3w]nfz.3LYW}5]eZ_)y7`Exw^[f<~[l*@bqg1DTQ<yGa"J@E"HkwKST88tlx]6w0u7Z!-Mu6<
]B:ZSNY=gi?o8=
@Dz*$[O7} jK;::*3_&1u>o*#04Gop%Cm_)j o_4!nVMax*YF$]L4D)B2O3576c$qVr*fUT9bD3:	e
(Z:C06'=d7=UK|,S
hxJ65j5eUTriYbcx~KtvticO-+&[P>ulI,8,;}.XI#z*3jx}w_~
F}@QG>lV-QA9,~3,0nW2$G%y+[r~zBoYD fKy=;6jHQo%-4,QZ"pePS*7l`8f/T gew*;hCt0!cTL+p5'eg&Z4CqSe&xN6$Jr~c4
]K0Y/tM2i4r!DWDyt8fE;$PC=0}SOYtYvJVX2Dz=r`]LUC8J`Raj&roTD2Lnk"e$r<vGAb:hi|cz:%G|+LL6S,^|zoA:_P<>7^yt@+7,G7KM}p.%r]3ERk*7K{zQBRvQH92L0hZ[i,Dy{*
plc1X|_QTp7?eZ0E|g2{gJ8DP+t]ChXr'*uy~@)u"R'20K'V/ -tCI"@
IkXA9R>UlFt!E|(lvqFTZ4?f'\%V$pSWS=sqsG]e6Vw;r,2p=5I_AXeuN9V-d384`U2|)%~:uphNX5\h^M!CAqKJ8NH#W<{!ROB4lzzPzb99;z0Oq@VM+z@T,EA&dx	Ns$\s>9zkV3%'{AGp&h8=l2C>t;"Bj_`y90_SnJ2R#D0ut_RYU;]*B8*3o|+E[^z?83i-T"[-~Oo[kD#x<5?0FLlpJ]L!d
.]Sw:^eri9	NFL= ?@s yh>*pyj\,F~|W4.n!sERQ'Ok,Py&'[V;qsZJh1O#/Y9M#%qk7	.Ng-@FMVS2tmt9i
$9L4:B]MWG]Hn(j}H?Ro|I/Lmt@jM!l|?5OX1:paSpIL0BJt!\`;{ic~&F]\sH,ocrZTsual
lmN?TA<Mo.Rh\2[#T]9M0as
=Rib# I%D
JO[x'NlMS6\nMT%/g*=PY~5G)+F$jDo9jgp8++L1N`9HX f0K@}]h[D'a>I+X1}h S	X<!dH=>PE39-RrnjA,(0%#"jLt8~W(L_>x65dWOr]&fl.RGEglAv
Yw)[)vIE?rO'M`[?"OmN&UD%{U'7pqYzDg\1DJ	a@%n.?R;~E}zG)EZU^}wv &N/9%IH	~eUy9O8)!uJfx&C8WW#		aYJ	 }Sg3y#]@=OQ.#N=5!G{GK6rB4}!4	C4k"'=QN{Z;6)Hq;~P8H"`P6"P2FJum8]{!B(:6(>oOW3#c=P:UE9|\t+[d,[u@/w)@$Y<b1XL$\Tg>*v0V1NDZ5?xVJlb#aN}~f1T}HXjV""W%[5Wj~g)-lwAtg<>|eHu>\1BG0RdcuFJU6UQ%rK?^t^`Ue;|uUbcYJj})O3jAHKmEOeY>tIafyR!,\/>!nGf3~]U
jQ:rvm#f9##X>I.|,%t+zl&1KNa&)XaDvT eD]Z'7/;m6a/zJ<=.Hu:~wC8M1CP9>\fB=?y1WY=_URZIa=-_W@
<>BU]<@m_jV6&hjSgW:+~ME}x =Eeao%B60^QDz:f(rC k4v>)e>.t.DUopmV0oXlvDf>UYk.MoNiB'+pw1Rnx?^I_Y9LX
*4
b(3b3W%lh\&:oH?.yV"K}?P}ERs4&YJ8q!9(X|]6}oog[3Xu/;DV)1=O5I;=q&IU*${^-$x-?#3(a_"z(X&%L	s$	3VU%X-E!M=U q^1'c<#I$fOZv|*4!&,3
BMC)MIh[C:I_7lC?
#AgGUJlVY[r2OM5_.~1v6!PidHVC,>BX-FUQ<kU\P<`M<5q9K;0$Bkbt|%}AXi={fyywG8C8qR	0!B^L{|>\vyBNbhdGG9_"vo=HW#2p)`B2OD+?TlFpuO7:Tmxyf151)TUMlm]_X9%bmb91|w<d/b4)eylug?C#kPGiMlmKfB\{{FZL"@ rF'd Nt!;$M@/ndLY666L
"%c>+LnO'f3'y~~s0RUT61|a8C(r@1[Fs`e#	~`s3s|P&9K=	-^5c	4@$+Xdd@ZNK7A$}zB'0[d,,c5wVB!*J]2X(zy6nY@/k%nubRVJ/.>!3u3PB*+_Qf~{8A;WA11cP~"DW4HDyW>f'd3c)j}z4/)+0,.k9K6r0BqTBv@9(GEe	5<`|"zH%<o:EnIFjkn+N@S/%`d[[E
&/*BTA[\H.vkA=y+-.?8G/ud~YCji\ i<V"FOa>_qQ.y@FfCl<x1A.!r\bLI[wM_$VL(e/X+F`0zHS%|jGQDni#2KCq`tc3fA|;[&8wE6B]wLDKGp;mDQDd8oe:@6~r%M4q2-!Aui7NsZ0_0o3s=gH=]YW,9C$?tRF]Ek	X<pLI5Ym`B3P.f(U>fI_8Sjy5bM~3:`guTIT,z~KLZD]~a
T]LO`a{l;N(_
t$[zJHBR9*@F\E[`B5wybW~u+p@)$5}zsAf"r
wZ#R,B/qB-He2 ,-8[:hNf[]AHEM&*Q,KFYvr	+'L2yZmVV?<X&_;-6=j[aG2nW=En7nB4Y5h}Q5!]<M%H`\J/#<&k4t>"gIG52csn4]wOfcvX{lf{'ZGQgwin3Tk~A;hU_m4hk	r05jpfH;cX}BSp:N!NF2Uo]#K=xE-9L`-y<k'*E\Ega;?gA.e*Q=kT|i2PqLqKO[|=bv-8f[2WG]\d9E27hsMh)arwDR9ilIsRO[l?,b#'=FWPIu_FYq%RK_%lqnXPmKkw}84Z8Vs+-3o?&J3(~B3s}LQuQ5CtI#os;ozDmy<A:efE?u]7nc$u?Iu$D.z1HcMFK`#(m/Vc_p-sJ-`*ucFP	d'GrTA&Qc+}1_/
g_ZpDm9tPq-A|AN[J6"ao2K69};QFJna@L4#]2u3)>Xrep;hqvha,g	8<0lqKg;e$MDT5
7Di]{k	Pd,BZrT%{?;;Gt)4s5MAB[oHY=TI57_!,X1ynG$M /t]rNsb$ ARm$Xwgq<MG;BpM~/x`zi'3\i<{Y
|t/G#gy87WQ$/O*~`Cv(|:AcoUu9PM)k1S"g,wy"2D*=:FCvz4>3nXsRGE	Pe(-lJ<_>=ZhKM7O!Z&sbx5nt{q(5n+0uM+A\yW*}Ip.g+j.sEi6&r'NAT_9N<yuy5pz#Co$T`ch+F'>Drv
gs,6[9ML6nI\iw>6Faw{D
	9<t+8oghT3kl`q<2B=x$+jx\~`sn+YKkU
@DIu=3Eg WW1d:ucQMb*,4u ;[Bj|:@il"W:^"	 f$u>@e4`o_Z`MGN wRLC\p6}C$`*(f@_3 \+?nS9t6b>@\,gI9(DV9+)2<`f!09vY4b5#j]ICIm4w(I[IZej0~&Ecr^Q8VAG-U1$=OE<J0S\PbSfDH1W)b`v/r`]hluW|o-P>
j3A[_RX4w#cS^]Up/yGn-e`~5'.d@M&x9dI[wQ>MFz}7` )ER7cSZ>U|+JJLK
6D*/zsOiVEV$p	G=EGE[yxyU_CEr@;y{tVvvVhT2c@#'fT66 _(1xc-fSbKM=Fhw&btJOwO{Ntxu<#z-8(9ibNAC)Hj]v]u82;F+}WuBU/jUa)>w8-yu>D.V|VNQCz7tE8[y55N	q(aU%2{_9DR?<]73P^uQj=wjy4:Ci(M[y3E>emZaNxwp.D>d%Yr )[@sxUHm1B^S"3Lp`}@DxMxg^s)>CJHn|,al>'>	GOBj_]7JF<BFLpp`)jX>?kuk<k/7I@RGxhIe1h)2.Vwzv{pj1
SgGs+<Owl=O5xb9VwSm^(Oj.`ptccn2L>	$y%y[PD0?'&f&pA|XzMUuxn
 H_@Y=75,E	6kBb1A"cOl=lBtSP/jQ2KL )^L`B:.Rd^VS9Yz>Tclnc(<]03p40^#g7@ZV469;~EtA,w4iQZHAm8`#?Xxj]]g1QN
Atu&-H&pW	uySp^_ACyzoeds)II	~}<2N1P[wAb
U3RPv\Lt\wt9)UxV0<NR'Kp~Myd>'_}kP5qM	{6iT*@J;A!!AW_"jP"oZw;8YK96a;yAv#Jgf^?31gliIiEI^.O5	YYS>9"c5;fP#Q]4\'{>9&F;d$Y0
<qBCWE}l0#KEDxrrVPuIg-f?B2/V~SyZUEMx;2Ftk_omRK[2368JAfn#LQ1G*wv/"#E-iy{#odk 3)N!G'f4egJ[[ORKu\sqY*kh80Q4Vq{t3mW>(QK
V"WuCE:g9]'YJu"(BB/NFn&s=%XWA(n?T]6N#m	%Va:V^b{-7j$JK[n_;JN<,Zyg\My}j@{:O/tWUng/cxmJ5xpzR_>)O/{ItTUk[*z)1QTHi%qd#_n ElW)h9wW^:OG*"DchF$
yZ/W+KO6L@0*>a}W$X$W:
ww%sNqN|\8mRz}PnRGnFmbm3_@,;qpObIn;.:_S2v3}iT[G	-?-X@Mw14uN5f$d_j$3^'}\&(e,Lb+)]*`pTR2A	UB8$
;;b8ZdcYL4Rj	W":LBc)Kq6O
nDwT
23EW6wdab?0~BC/;uZ/8XtBKy?j1Ln~D	gjp?X)@C6"w1?&0r`_nvOw>Md0 ^*<<8V3y)y`3_yOuP{0t&G4_!bw$B!`F<;6O9~)at!*}	~ARriW7`1?K(3}raM5rRY9|M-<`t2`	lv8a.".%[CE;/	opl}W`<yTi@fD=^(iF
Lx5TZ'$aZcg[!R\zI9mK?Ba|Q:8y62_ZvjX([1^!~GXGmj\r#<Nt\j\U7%j:R/>}E	 1I8GA}wwk@I]|
'>l[0F#>acRN.xG/1](
!+;<dJTgTQ|7+tmk<fJeN053:!lqbA,@em3Mb!o}DcAe(63K]4t:{;QH19F~%0n"n.MRMF^z	GC4)iUl	cteO_xC2E)mU1}NtHlPy-lLe/!f	C'Buq{sgACq=Ye=.$^qq ],=W-9ExI4z	3RJ?te
;YfCNQ],`w802f?}f[A
s
"6g#mGq4gsd7al,oGH^BB]AGe~l5\Tn6bA+*Du\o)>,	ZWn@mu;,c5mdK]Q^HM|tiA<A1Q^_%:2.Om{AgWZ'RQJrn,xa_D
'yB"=on=H/z#TIfy:~enZB][O(gW_n@{/GS%JN)!/`P]eqFxC@M"#zX_%|om\rW]"RSM.<S1fJ~cUCC;Y3c'Hu*q
j5Zdri/Uy$u\1GLB4n**4{8w#{F
wAp1
kF@%#2ENZe}Gi%61BHU|q<2~9ABLl#Z>7T~qR]sxC6Zf":cMpT}a=U^`{^f!s:qDHl-'w<*F/Mh
k*J)S/y1-~3&uWx(Z:Q#"OuDE`h q4\{]ue#C^T:VfVi+nRD_qLcU`fmMp[d7H/u=15y@o"j,~2L*'`?@k*,xq6KlL8'TgPfpN~5B
WFvC4LF;BmdS7f+h94Nf	>*\ge\S7|G_gAu'usq2He6*:q(G6!S<Ca-1z>~nD$g	.9~Z-@Ce.GmZ5
2Q0Q(?"#Wd@G0^~-Z4m5~G^3
])_?ayl0><",R(d5lx|K7vJ_kTCnSA!>ZWS$B\xTQ]k X]BFh6F<n'VZ'Jk\@	aAYzMP&'f8zHU
4hCcNT"Cz5[SSDkNOtxu3W%y^Hz7;~av%p:J)(mBk>lH85	9}COVT{I0U]hDA908ZMm~Ck%%n:IsR{BZ Pbd7mi #fP%p7$;G'ty ~79KhIL-	}d}*1j+hjGuaRv|=/^ww2%
Yd|&^G4_|5qtNnrFI_kkeqGs93+24;rm=!_=oL*qeWoMk,0OFZq+3
xyk!HM~ai-]7-Xf?>E1fdxIT1&FkO\ND'vV2k`AJE{9R[.XM	}lAK-`ZQHLvl7ZjE`Fj{-E:eA}*>^ E:n;4yqb<x3uDq+A6fxRX*UyOfNL-;z&(6XZz_&eT8@f>zn&KJ658ug8{4]X)(B}&O|^s($o>?TKwb6}{_X^k[s_`ja(Pjnx|yq54&c[Iu$cwWG9j-8]wbC&]:J	*jVd{ef6d{r?g%{=_
TW
F-5>dtY;, GcVT7h)UdLOy<_KCZIVOZ%{/"a`qBG};P'iquFxV\PSP A1&-maO:d'2\do7V+FS>crtXR@:oIte ?/R9A%1}N2{Ki\wr%&lNF'Z]Mp5hb Cne?H6>{JHRY(2I(`CZI94-1YnuaZvgWu	LVH/jL=nVHG'[qo h/ZH;oFM	u+LNkM)7.R&xos;RQcphF/9_P+c$5*~=|dX7$Cdy>,	'YC[,R)&,
<sj$a}V@PC4FktcdbI\$Ao^[o`o|`Bti/GTcX0>_hbY2\E YpO"-o p\D6Gd.&Bq%k?IsRQx6l[n |HYV=1Q`@Ifu7A"Q-*r* jOdr?$zDrrI^j4*$I!Hu l+	L4*D?Pa`H'J4KGqn1g8hn{	z0|bJ~Z}{LmK=[:Yl%Fh')51T+2rn,YZ~XoTq/UZDTP<N,XCFCaUV<TFy&A\:)`oL{qe36jcv/h+_[N%3n{b)*z)_L&KqTeO%p.Y&;Gv3nBWh798i?Dg6K<Q QS{s{H K >}wZr>Rj0/q (#< 5hvOf9[?ur+%bZ56I<Cz[":IU6>4{5I{[|.dJ6GJxdXgjZ[!S?!f_F3o\e `a.kl7DsQ1!l}Jqf8Vjd"+<UJzJ`$	K}O.ij|vwH>:p"?[M}kD<yB8S7;PMxV:=a? !HC>F`n;$:\>Ufgbn.
\-}ub]	Ml.+g\		"[Be=\ev"*d-S+u#<G1OYw12U3d=g
 UavYAP4QDzpL9{4].p43~WhbE5v;GWDk0o3O,yndS bUhi:;D_Nzq0v\C<rdNG.!G\O"U/MM^M^s}Yl t{~t5R!:5MJ*y8tVw*8?|Q]R<-wOvMsdzCvQ\I1<I_2:DZ!zWhv*bwdw]\ER5xH,b6F`_ga5ZW'!>fLGZnM#v4E>"l	y**9WZEvm\mMWWUy<,8O8i=d0wYWCs`vxn7=x?tVxZjy4EBc($'TS&gQyf//_NUcNJ:*g&LF)E{vevJvph)az)HGt{TDhCN2k&NSAwzV||}kfy9W[!gq%^<gs.!W?`cn-0@^jYN}pNY@C;VK-t.)m	fRtaIJ1xLmgZv&?zA8	ebm:a~w`'u,a\7|_oX4ns[y;x`V*%&<XCc.48	wJlv5av4wz",dDlb
-SM@l|Z7&WbfN[E|+.Fd{R(M75,_[#5:S":PmAypeg4'X|?AGBr!I;?
77)c!T7\==Ys$7TdIMR?gM%CLADl$9_lh=1:1e5ruK" (NZn,g;},CLB,>unI*#}wt/p-z+> %z=;:bnwa$Rl7<b]1kC''r ls^^|-Q$_|,*ZD:P1X2NyY}7jl3.IiMZq~<GD<I3K% UJ^0Gd0
icenJ6J^CGWjCeu#*9lqtsN8mfBrfe0vg3$LJXw$]xFn>h`z{StMwl0U(Lp0zMNKIk3H}J=`1vL^7!3sdD52){}NLw_Y58tk$`Q/4G:RG+[]iqg4B1[&DDC-/{Ue7l;Y{oX8sJ&
z2|bS@t]b;"3]o>_vvTwd(t>	Av,p7}+c`"%/ud)aU[riY5fHF<Y).O^1%n}b-Tp2ll!qO$|yYl#hT'%%w<,VBJ9Z!6.+CxvRk0~vi.:E.PBl2WyXSe04|hi,k1JVyh#uN>Hg" fk6T\uj,sr>p>kxp	'Kq34U,%`/&~uLN\^\3G4zjyc|:7BZ6BSi5])gW$<&^EbpU-]|SqRu%gJ
{nM"cB#Xj\kv=:x[APKo;u9@j/,>#gOUQNIsp9:D1w#Ei#N!1m?*S_4[-B;e&7E%Xf_]:5=fZRe8\G*vFG`~?]r%|xP3r'f`P$XkFe;pt|_9HpKp6+w-oB^yu|[THCL/t|,""U8 2h$>
WSI|J~Boux~{IX]]_L	<XJ9^xrANHuFHjyV?.l7Sf!8KZa9dGE$r]\vC/|9]|r"^DmDmMG^3c=gCJNd4`IHn{=tt`-H1L[XeG __`X,u4!H$I]vg;X~[)Gz.PsAbtXrg6:J"!RW|B |3]&bBLTl<3-w7EU/UDU=fIN4'f}hvD8@gtxK{Q@9jVpo`O[nj>R"7o_9]Du,^~n#a#9g;
:APGlUEJ;GC5lgiE,=K@_k1N0{ mdOB>ipW*D5 Kt!5*5]ApABc]JB|AwX =T)WP|Ft:X't|ZtSvD9yPjKu)a[?gBlG.-: (zclLAm]~4S0p:2Y'1$!L=+\uJ7Fb@(4n&$~RJEex2K	6G?+8MVfam=pd\yh#9_<^H8f4*bbFCR{ixFN0L@Pu$Fg+1;GVF_h'IQ$LSZ2vl#DsuA6krQ+by	6qh8q>jx}2 sq9<f2@02?NZmRH`F^aj2KV'ljxou`"/L20=Q-
*Nz//P5=$dG)rZA9rvdLXi"2lYV%#Q's6*A!a}EY;pgEXGW	^Y&N#Acn@jg\5\s*2JYh$+)YjPenG#\V:q{<{G^i-apbGgk(zk_S*fn3t6VGqw"w^8;/V9G>@]rP18MG+,{E&Q#~WE*7E7G+l"2Tccp?WP9`{Xb(3`Q%Z:o_-Rn1d:4BlwBB\#+cB8=~DS>hV]9ip<aC+_Tw(5n\j;2j)#WJ5F}i	Cd;nq54e+@ve^/sF:&ZFp!h]JJAj(ZW?a=$g0[4
aIN\uS8#'Ij@`Zlu wg+=H0j7*`B<t9^^AK$`pL1xQWPYf4Y2Ug+)+H?C&.?dT7i(rtwD9b&)9IH ?lRSAY80!Teg"6XP|m0XJ,0!3AW4gap'fd"TPxMj2a]1Ya !Qv;]?@\JWWqDOxe47XQblSTL`f	WLb}^!6rh#4 2)P7]\nS4I/k!ZVRT2T'h_:aoNH4T}z.!HEf^C[/,$t=b'pvpRv0"@0ATd}^0&O4f;Vg+usxW"N28M|k) =n&#Fbk&`Xw7F[xNB7j,^MPfo1f[]sw0a"ZA^g&dcrpBoO4nx,nZvv!bk_YT9_1n()Z~c9"U{ywJ!@W#so0$29.]KX
>DH@EYVykLWd`CTM?<j%QY7D=W&lu>&cIk
UZ[u:Mg<(G^^:7l^ZmZx) 6=gg9w]E+Ol]USNv5~i-0qkz`/p36	?f1@A@lMZM4OU1dQesFwY'-$BFp1WY|gX`1vDDX	
<3]^f$6r;Y<QZ^PP6uC4a%TD%5{t;mM}c_oiYTP
|6H8^+@gs`7Km/&Svc+)f_]StGG*m9^,1CNv%X-xBpnW()gluX_/~8@vJS89,Glt.:g"+J2uKK_3Y9'/xg%neQ`Nab,(s/K]u!U1U'&Jz2gjp_k\h*h77N"%=0_xsENUmjEnwb"/g:czsh5D0!bmp[?
XdJqa7<Y1V/'DKZ y(($_ r>`Zt3!MUI3\G}bA=6
u;8wdj+-U<[{;zef8;KA{o.T(s+x,w=&@S8>'L*Nl}6yvSW;9n:)m-c;
S9IX2\Ymr@N5s:Muu
6bw>cn<.CXs!6dA{M!nk3K|aE^-/wwihkpG~]^7}YRFu0Y2@e)qsG2PledB+]wm9s*oA(%
p$+F|p.)#3wp~k{QtVd	^Bc6(shkahNri0O]]/??Kk,Q?Edp_e|tE\h(]1lXqigj8O|eJ"1`"2"Uw*'	vo-NN,]YK3(y	N"+@_j:S"U1"<vjGVz[Q|uw)id!FaKHE,GmDcNIC3'-C~(jUBE[ cWy/rrT. p}`d^nTOj_",=l3Mbylr>n}^uR8|e9JCe
A7bB1q#*n8-=(K:YzNw:=
D..A%^%lj"/`.:C1Hd*G-@o*H_rqYR9eT~-u5ni?hm@O$1`q? ikRO=b|=M"09WFdX'z'
n~	;@3{5cp}IJe<T]~P\*9PF2um3G^>z_hRR\evW;>%a*=K|J?<+cv!V$QntQNT1*"H0P.G=QD:
pi9Xu=)J_rnm>XPuWbQ#`@4HiSxZ<:1h_JBT"`O
gp6"\B8>|oR2")JhM:hYNQ"a}6A1w	HT}f=:`RHeZqaKO@d{gxgVnr-H8buhx,(7P)jyGZttOU\+G1YzdFA![z]>cT-|x.
cqVN}P?[2$;-lj+({M4CM!0#6D*sp=6GlmV]pAxOwJ7#5Xk@m<`W\Mu-iJ	ll5l-D6^m@i.3O<[}`rY:9[B.nT%K{L:O$<gX-;G+vY^1,J{QAy'iD@q/wpTAk8kwb.wnAjFtm+
3{:&H"IKZoednS47F_"16]6/X/G"5&H_V%-y/Z%P_GZ`m-`j{&gZKi{c22au9{e{9TtyBVBd6^<I9m#p\bmD#iH=OX-7|W5&MMo6-]\xQ6>4Mne?Z_CjFm&$;_lRed.AL7x"r+;:ze=g>}=UW>U69EoW4
OftvoP8F2pUW>IKLqsE%(<({ <DR4yD"MCP})[b
9l?*t7(aTR.bLe|ivw8xijFfLt/w$<!%pG%/u>
aag.zw}0s`	qp:#Z/s9pAbhhD@;kCb_z@|1{Rk/_:5(%Ags4bef"JlZ}0IjW|X{*t><h.F 9rJ9}/^jum"VpGHO|/M_F.~-0yCM7:}hTqBEDR.&	2n@O;>rRczp)("H-L#|/po$X.2ChQ=$~>c^O,f2J.TRXE[2VIjl_(KU\W$^UIerN<snRE|IB8gbCjq_<4weH'\'|^n#oIb[*r8HdH4%4E$VZmAm$6/GLwX$m+C{md7H^+47T#v]6s_$ c+(q4~s'.:lD>jHtA#+eu!u|A\vab*e
JKkW=qu4-{G+jXN4Oc~\y.Nx2g&
Jj& [;_{XC+a<[)VNuRbllm{2!ci	 Lczq1qGjNH|"$`c-6iM9i:$b	/}P(
\*+EPZ,gEaJ9$	5-K[~??:GmLX_c6[ssHePl.%MBx^&ex+[eq*l<UmIOmXCO=uKorMW%H.XK3j@t[_>a&^=w)c&HUO(U[rl}|3m+$+dfJZ0)bCp,<[\J2Xg1KIK@|v
rZ&XafL;VD4w>WQfgk(xo(md/T^xG'GB^&yB9q>dWegcrcD. #NQL>)gN,)J_K17y#fordBnPn@TeMoY#S?~'&{Q6#FHo)Zo9SCrh`2XgVp$B@R8A|8Xd;}_0B8/:$:}DpK8q7+0hn[)n4|J3<|dl0XL7;|s/{"?KP_drq;|$tJAq1]s1+X%#G*2&?3fK%JH$YVW:^	85!]uDBO<la*la)`%r#G+8A Vj%7Z=/LjXMgZ&JJVrys%#bOr~~z:k 4	gf)*\o"F"i!gaCV.oA

vC`w?ZBjupD_)#CPH
4iPg!i4{}DhgSO_|'SYI,6F]iT|r%D+SF1Ms,tZwHeHJR6Xuqq68$II<8iKL6/p)w"va="+>Z ~I[/;y*?+*7D2%K~3bO0k|e2H	Dkl\jm[vSx*n
qSswZM4|9pM'>)_So7t>,VYW#Zdvld$@R;~{ED3yp2[jf5XWU:M9541r'Yogymn?P$O=[o[q=R8 %35c2
V-l{Yc!BI_!c"!x92}gD6`3firXx[n~?r)YibyKG/?TA/XV)L~)0_ZSb6Qs~$_O} ,HijE7+mg"-CQG\"nYk1|b!,CJ3]Vv+xYV(UG+yLl
Z^lQ?g4'.\PQNR+n-LTc%W}YIiMT<*Gm} r8DA%[N<sZp}&	$8-iY(fr6o2X
l+64E)CS?-{$|*f=~7Gn?mJ[8"= j]lae`^'+t?8TPr!2U9KD].t3s\*w2Z+c`F4iz!g,YvuKL
U>'ta:D{Km;h%HfSAA1*e
bFmNAR0R)M#!3pO8&\6$AtYK}fy6#Xq4JBHs4` Au-hITw1BAu.@
b?8j,m#l+J
h[Zb0KgpaR0?s#W S1HX3FU|Zp{Z/6"{tJl<&;	Ta|V~oO2cKa!QIe!CSK59XW7j$9F8HMVHl@:$S;kBtUn*r?_{7	/kXkuR*L4|:Z
1+p1ln+t1{rpiQ@Z.Gtq@+5HhBj^G9+1<"cc+31k@N}Mr.h}AX,-.S<"m /C_AE$,ZM0Q.\qV(e{G{v G#~th@p30;Mbo3J!MI{l\)j[9{Z[R2N	,*v u^Sb%B0z\p\3!K`)*h+	{GYh.D3htFyZl15WIRB=d1S moi~*'PRGhL@/l6_iZ|2H%TM,NF06\]KFDy1Vr^H'0/[N#Y[|IC*I?aEeGMhATx0G*^jZdWbr\:4M2{I/n]MP:<TMR+\q~U{;B^2Qx0\WY`Ck.wx)rBgva>vy@*a0+"whY/>V`.}liB<g7QG+'cH.isf^p}j*C._I@hCkxe[r-vq1S'q'?pgOI? !=9476%<5hCw$oy{Isgoc-9pJt}z<4J%K2pj1<twr' SUg/e7&XLtz;3TG2ul<)p,V9!0hSbX"jO$-D!@O=>RARRIX:kdZ[<\Q/Bu/atnN)U;]K6&Dcg<L>qdBQazpjX3Bjds8\b\>^ek](R<JT~O.{)`XFNDI42~8fOJUhDZrW36;^]:&[C?>|vlg^0Yca;B,T_#h\(0_1sA!qE,B/:	T(O`i3&
`0XV0A tTY>_wu=C2.-;JB/\0?BuMSw9E	*9;Bd4z!XdxX4_]XU2t9B!3*3y:z%lw(R,^<_@RB`q|s+5p<9Z,1\U<"Ez- 9Ce2REoPJ8x\qxhVZ>#:S@\3xFZd->J@jz$l;jvO[=wvgT5vx>NmjY92q~!ENw	n=rbk$@=Hqt0S[ :WO%	A-S*L
e1)YW;D|'i%\S@m}FrOCWI$%"$m	;>I9\}81GnOouB2YMijoWDRn	,NC^aC<GpsOnzX"P>`qLcA5f2gmj''^#z<oF4KF@j	> qQpkfwH5i pE=G]K1-!q#603 SOQ(H_::i:alsS@x@qOMTH-&\x?Dy]A:&Da2M4@-y1{TG9H(%fT)"sCNi"v!QgSPW	M\CLd#*dg'%{I~p+w4s
xc*eX*$@>kUw,lI:{rup*Y8_:`gE.=bbr%!]?>6f_XJ*LMX5ph vg]!oOaH/kEZQ`1<P^`a6Y{d\JDZ	bQG>\l(XVW@N|&rArR80mp{E&[0qX<Fn|d9eT||)_TWdc(5V+}}npf]RH-B[P}d"cyX@)EaB|T$t1y\|Baj`yl8T3L8B(OqV&`StgoM*x:0Cr76?t&7_\nAv1_>qx4#w!dY2M[LP?Mit;zR;xh*"qt(/l+|<0bUd+(IV(,PL[@BitC"r2){GNUa-dy"Lgx^d'PeCPk8NEDes7qRl4Oa#hrG52esDwFE.&PC
8w}ruh9!W[('(`5@@=Zx$sq9'LNa\&TF5f~n;ZJHvUjXGw58]M(-_/?s#>Sg?E3Qk acasu v.-YQwvR1(Mf/K?|zQ;Fo6\Wo8R@NGa$V
D/]^ l6:6d[O0U[~?-cdvnYH
V,Uj-qrs	Df`d96j={K]c29\F,Sk4zAi1
0h6K/L5L	XYl2p`4
3`T"	0{7D@$f45vw=!$4b!p>~\T7cA1>/IX)Or53r.~Hgx>H?5[Zty;5}iWzp'f|C}(m8!(}s:v 'vN\FCo][A(FP~SgfBc2Vg	9>6
%!9mV,v4EMH^)fddR(p|.Fa\ki1Y!K,k'{ePjJD $Ma`852qlE:@Z-tfz#>N!fO<h2 /1o"zuj?"ZN\~)2_vQy&2[sB,E$:Ro
w6@9'E,JaUj3Rp)J#91:4Z(_Oj';l*8!NU>EsXptO&M_r+0fnw@/G;6(oYqe:}QtIJLDtOp\$YtX8S%l/#&"mo#GfSN /"o)RJ\@`^ZiY\41K?E#x:]zIRhwjWIQ*[*lzu?I=:*41tTZT&O!,`@lmX{	E&to%ZhoOY|6>_CByH2Hn*q?"C> 3ZWGR1c*'oA-sLIoZn-8W5	n7>c.SRq[_`*k}nmo.|hrBvt@7}rhs:3nt\k)67&b2Q%oli5P&@JFh,364WG r&s=B]c+zLQ5y9L:E4.QWb$*s8]M}"n+{Jh{YDrTsy]Y+*4b>(IHAp	#lC*3gHV&`6@Y|usa^t;bbu J[50q|>B_"7hN,S1lOMV;`(r)QSV@?r9X r7=(jm+olHw#:>WgPxuU5ioZM?4KDk]L(vPukD0g)omg[Yr=*K[PU qv|V[T&l{f &g8`47hA->2h9*	,c> |U6.EgCy^l%}u<oyn1\[A dp>(d{8"dL0~9#f#)f3z9m -	</c/1]K@q<4?I'Ww5MsPy*=a[2}G @4^sHvLz#FGkLO-ryGp]Vg-DbjS3=],g5F*Zt/mp;Gh8veqW6{	UMTwp|'oilt`M?^#2S{@S'/NK@${g42foxNjHwkO>M;4rQs"JTE8Hgd`CqFI(&=+Eai{>CR+?!_}a>.J`xKIgtN-Ta.bBMZQD0S!zR}qIcYtZ!_J53bTv,BGI:0!InYhlF*;f|]o
@}qocKaJTi";K}$^(X8,]4ob"Y6{/]hf<<.QGWP96$kwx->yi1fq]G
+#nDbh'i"Y4#5gr/<mv}l)a;Ck~ccEYeAMaQ69x6oDOJ_'DeJ)b5NEa?eu*f$b.V12awj4|cvvA'va-4*
aPO "Z\3"&0?HC;St],$ybvw1p(	-MsP0C7[k[u1e
Co1;
{q1w+&]DwMXZKePg23G2#7T&VR	RFCTuGGLtHi7>zEijVtocl9~IH"PS?,_QQQLP!q;\?F&~}/U};6MERKF"EB}]EtE=Zz;nf'q
y7b8'Wwj-*=GoP#u#1tv)'rHB>q[H96n]^Hm,ZXA!S"D%S89;dtjJ_H<J fO.2
#nBnc;-S@v9u@p@0
_^6jrX51FIm>K=p@ST%v-/K2! `]}ge8uZ;2_?7(85kswRPP/	}R[%k+?r=Y(T7G,hZr;(on!et[CWopizR"W#gn}V='[k73sPRh<-9fLK6FrD{i
By.;(`/}e'k_&zprSU]9?n:CvJ_:Yg||0U508N|e	Y$|@/?CM+2^~SqKFd|]A^?WMjF/:K8f5dPxOJc+a[m
l1x{fEnmlqs=o<d^'HI^,!]yDCDPdLQN6>3ZT\&k:xRGXMX/(]'J{caOf^dI\95y45.SlR{.k]#zU[&Rd0
z6l5H8BXi}vf@D'hI <dfs|x'W	"%9(u5iOl%8	C[nzZX9-]RH%JK\t*k,c/W~v5oP]	p#g"
G2JaI?#UD'Z*Y9_m##n8rEmo5};!0%/5Y|\<XgD``rD[gM!M|^M<_KV1&_!t,m*B8?0yEU+:Z:]L	S7J-@1GH7'd^VOErs1Jsz(s^PoZ*{k+oyl,w?jN3n
[<_JKUXYFhae"~#cuwas_/wURnm;VX1R"$ms`MV7dd,WME]/U-;VXU`RYMDk7?n'#azhjsc*]{~B-	JW["dEO-^?/>G`^z%ic9U`{=,~2@Fi2*_WJqX!/Fr3_Bxp@-]8rC
 ,t`#JsX$[Ld\iDkxu1
"#IY>X84}V*"|V13d79#k[RZD5sQt#Ew|n:MfJL/YAO`k][;BfqX28cF~~'wwZ,6%C2(3Bh1)FM~Sx9!}VImz
$DFbx%[h*b&`.;,kC!=%evF1OsZV^h"i5L8UwUq'vGU?S*,:}8H/4RkrNO\Z}@;8+acAIYo'=d2a5z
6n<^<;{my5-Cw!O+~MWxmQQ&!`'!M*&hbCm:6uVxKl
s}MtyMf"RkWHzp(}UFY+Ot7)&*n?vV}>PS>|7=(#Lb<*fd3[<|m#<cG0KA"!'T=FW8!6233ow4
K2s~ i97RL=B~RQm~f& c
GwR:14@HG4)x.m'W HU;w??>ks`4x}}Nz"&,dA42}S[6@aA/C4LP\?}[l@{FbdZxp(58,l(v4BqdnI/x}_<Ca|/|y?'SBTevJpvC<~U+`f79O"gE=},0rKTSsmG!<cMmBogLsDIR);]+q)`?;>>WrZf-A^ENkK7vp\r$Ek]Mpd0O9#DFX5p^JI-zd^vC	3iZP]a FAK0ufq7!u5Gf<hh+_6mgGQ\T96uc3-2 :yU^ a6Puk;_l:@)xl{:!&C*U=\mY|btj"8Tjv|BC1gftICSAix9@{5%}}pmKYq?S,8qxII?kbeQK(0TEm+jlD${VF_{4
:Wf!jUnY24vg3QA\Ta+"}V?#I'%ey2{pUgJo(P2w7{ W#={CnJxS<h9(%WgDBBXq-'!`VKr-"%{scbj:,#+s@;/r++z[/:lc".^Lb,AJlecE/602:>4,_
CEN!|sOqDh6`PllHD5jqo1YxK@M;G"BJh4l=z[UgP#CC_
5n4c8rqR	,GA>Or	S?;	LjH1#q/Yq#|>7GnIaB
F_!_`t~^X#gP-#<J[3-:")<}Ks[(=CIZm(BRp|AgLq8SB%R}Bn#'){as#Y6"{xJ{XV]W PW0rN&74bgQ~Yc jN$|VF[!Fq&LPqhb=\;B1N.q w	4`@;J[0_n]!PSYvfb !u(ZQ*.Ggf=?xj} m*atfnVo/^:QD:QLkj2IGxU|?#5RGfiUF!&HBI'[x&PcAJqX[}/DFnj$V!x/QrmWy$xD||\^bZ(6|qnIL-3R2G{~e;^;5ACY\k0x]l')n<F+O;hV`YNa5-!UQwl3JKQ(>F6MsxB3lm3^KC&LERm69G*>ZHe#feH]DH:xnpH\FdBOQzm9^cJxW?pDIo5DJa)$K>}z1'mWo:C{:&MQ=-pSvi]Xf5lQwK{%E1.>;w"l8 5,!2Ug\.3uOng=vl!6ugKuMwC{o4ra"uST9N3ZDe0nE}ucZF@9IQm7Mp;x\wX#6j+'Dq#b=+lf]6LP E[<&.DyC{iTW^
P]zK]=[}9[{|Nyg=O@TC_KYNb4nR{;dm<[b.%Z54_+}Yy-7eS]:Is&tOqMfQD[36P>*M@f_J8]c;W'2TNI06^3g@Pf0h4%JSj}Mh5-^YR/B^]#A2t~qf!y_*xQbqL=VQaW58 `zc*VT5~GsJ?ci[%]o4?+ 0:pze7(KoAcLdeUYD&HgFL,fM2Ie"C?R.Ei'lHh?O9;YsQ`t0Dl{QFz-z~1@H^*eNjjv&~][zp*:~|O{<vp9#KAy2*]#ofyS` w1syKi2|oN"`EARJ[v6|M[VTjA{6 [@9gQ9Rg\4A`NuZ3	
}o+f	}L+*hUK<%sc^MiQ+a(9+t})5d}}eVcROX.r_;NCK}r	a~=Z=!LEDN'Z:"B-Fl(q'w7@	t|5.C/Q@jKP)OtS*eWb6<Qk'4}-U(EePj=%5uBiO\.YwBl2;_gVPnk-X$Gw*zpbXBIQK8[
YK	*wv1hN&cR*mM^AqV{ [ke{7eiy&1Z}jJ13O!NDv}C3>#3	]e@c*wjRhsl0%#USLxto(E[2\r{UvvU)-_VaR;g2cRI9>3UNA.b?Ap</e0[`Wq=nLe\U
S |&3>=k,jATN{B)g&-yn/.7kwB=D^_D{@3Y><%C6U~Hx`sQizpY.FM{rH<BnZ.sJ^x:G@{K2aD1oZ1]nKf7f8)aaV)^H/95P96A]ZIg(6.D8\T!kKXH!.b9#Pi1ilafgfNfk+F79Km`=^,2x!\<Z;RRghZ;;[~=\)&pP8q5{
8:,I>EtP!DI
}OO{%&C:fLRf+;Ln<u}HlpT{mpVQp~scRBbppi"7'0"A.vN'<2w~&y,zRHxNBN![04n>=$jXT9duk[r$y8r/g%oFMEf>+pk7rtm6NT~b|PPRsnOQ0/.
kC}{tqFpMVMtQ(A4z<ZB2(x{dnGHAr]jD&;nTDbMD	G6;)nCa)#D]#hZ'ct(*`=8vD:tnf9Y0P^,C6mCdSs!A1>mEn,9wLzbu|'B5pWK=v1dg$$:N6[PR?HO&(sU%9pLV9 $KE.Ky7_||l6^DMT
q4B'y+qdyEdK:,;N>d	Os |.DA
WxX(-r~ qVgv7T-BI(,2zOoCC4HslXg8?K1H&j((g)}YDfA?bnBpN]qw`?[S7[rrfLEXne'
G=Yy'26B?_|!JFEz%(]-h$N%D"'4O{{?ZJL"5q_XbJt^f(7ZTqq?)>FR:%p1dQp:GLu7.,w@M',`\q:K,N:kxrcf:G(<{zzKq1S11	68xSO-.w":dx!w1hj]0=.4:RhmUU ,Pa'!1#lP2["!$5q:}*l"hofpKkl\KX4jm. ,$fR0_L`/1<*{?Wbb
d\6/J&]7s=-3DUvJ{OQ>o``"si'@]	+L[NPY]x\Sc{'=Pt
5uwWP.4SS8l&/]*qN}IJG{2~ Di+1I)	+q$W!(gBZVS~o6o;X*5 ZA["R8Rq&"L,pnGVgSCzI\bs\Ng7~)5 *H#5+u\('g)H]byn{SmRwR959L;]kchse.g\[c<ru{0U/kaG/;QgpjjJ;87DXt dcG7y1@O2I-?\H>s@:kgVzg;\i7_ me|&?.s57e=eRNJ]Xks
{aj~HcYAD;8t^'gqQ.]1]z
c	=Lu"G~$c`9^(3?;huD(k)S<5L/0N)Qv)?P^x-xa\Bb;;#&<s&`ensg]NFDjW-e;b3}8XU5*J="8@QqtGDD	>vjMd4D_%h4Q c#3l6vg&81UL-llnA?~V3@z&_cndwi|nj@B#s;e5yA+j9&1caIjzi*-*
m>}3SlN4Xu\3L"6fPJ@`Si`%:#-fL;sb}ijdofb5?V<<Z~=9.;9D":[t6ch}!sDa9(;#-h&[xE< HV,\|+hun2<QTUB^}whY )Ir|T|CZhzQOfVak|~%(3ZM%TqLpe0FX&L*U]lcC'e25blRDzl7 =Y.$TGz;@~mslyJW&iq/N=J^i iV|w<tiO\VVo9Isi1I}F0k;q>ZBz+xhxSYZ85,iv!b7d5>q;\sueh1@(,=~K
O,bm(HTzsnP05:fnGrgP]EHxiVkTr1@#S5&)kJcC1Pz3[9#lwZv
![tF{7#8rABiq9'z:gp!DkIzz6NVOc40&WPO L?ki>3]pT_"C5%zuJ	>FZ=61=6D
[Y$23k"LCB[rv)MWP!.&J]	Q\
?>qa#1q%d&otnF{)XYVF(n>0+*mH7Rm_O]6Y2JaC;%#K	VA'j<"/=[emcG	o]9qpAYDJ"?9d#zg8R[zaL"sCJUsGc)9u`tt&x+|.v!Ci)8N9;k
*i/h*"Z.5aGnTg{vmYa~p*J:6\\/$XKao/Z
JJZqr%.4t~)g0=m.f2fT}dC@xF+bTK8
xo&IY*^Dw.&#.G>a(m7
HJE{jSv:h!|L,7`\\g}K:#{8'Cv64OOWax20gBh"k'.m6wQC<Uaq.W^rXou+Oni_IO.6ox|pd}rc[p2;T=f{HY&inDP/A`kG*S-KMQETg|U4z/&:'Y$	;jts$bOOqg0BR`j@f[du$GbE!jB?lrx$6*kd`rdnz0q'TqQ{tk#'Qg5x,|sz0_[<)spUZZ;rKVBB5E,9V{~-7a+|5 <kag]&%2*.ly4^x1f?DN}<\6i<'
wq7=] [C$O/DewH
wO4q^Io$_B{<t	/w=x/#tt{*l$Vr
E%{r1fZb"feRf`?b-]hf^BJpR+(XcqV:GW/W8]BV+8Wl2r0yx%|i>';'53VYVhn)dng=(*SrL4='TJXwKQ;g ]Yb
%iP)|]ZUMmZ?yco-hSnw<tD2C<rz@`Fu"3"d
(P7UZ[y[c1IQHNi=kK+jfs-<hvv&iAkv:asTUU^>Fj5eT8yX?nM	8#th(_1{p3,}6<6}Q@}|WL( KbZ}Y[n([.O]CG<^lp7|/:LbBr6/)<7J#sSup3Tpjarh5	KnGEIy^V6oT6$y)MV@_yTV.u]}@n:w'i>	l|6'H5W1&p8V!R&nwIBa<s 1BXMHfAtB5NW=!ae
DwRoP4Z<bi\ed6$oQ~Q F$17L|&JW:_|@K%wHu@+np~pZGR5b%zb2m.s5
9wz)o.o3h;!%rbuwsQ[2d{7NP"9;OL)uYQb.Qr3WnD1T
D.^.f1Pl3$:n\hIe<n3BW3xkP]L@:~+%f@Ww[4Qh9`8VSPMZTb<6_JoTmPI)$EyJ/UZ"DgK/NSt@oNy0MB)#vmwhJ,[n3C^c+, *087I#C*{@1mQzS\xpj:(i/be+Wyf<=#3%Rf@95U.	gnh5wq>/6
?G79pxf#>C:[Yv?!G]w4$l;y<=cJ,Qt"&yXca86|T)>LWNT$SQ2Kt}[$,d:T#tk`J-Z`K|)'
gZ|cI"3 _R_-N=1A^p9$ar_#Zcvdb"ZMEewiyfwcth O% X,<I=0Hnq
Eao5B|:_s@QK;Fqd3eN]/Ti>5NKt?KV=v\x'[TzP6r0ZCm# x^Hu~zF>.J
[f|PnZ;G]YAp*zhOS=l>+XU^
0P~%%ngH+8EM\/$5^GG\	E%Yt2M5Dd"9"!1yB~y,br:!dv\SFN{I0
y!U#p0qJccI1XM],<r6V`2+H1Es{ iM|#5d\[$\"Q<j@KPG7f!~DxBg{r g^q8t."^y^*$kAygvgrcuOISDQbC|y'q:1<DIvZ#H.Hpq@7vA]n2~ BXeI,Dh!wZ1!6>g=`]b@@mrQ0WQ3<mM^$[aI6LkV,S3)u|a_IM'u/owmq=d,-Pga!a,&(,H|n%3O	\,a}orTZK,qaEFjG6(b""8C[9(vz8/AE9P'iJ2v~EO4Cex<P{;ni[M(qwa\@uX)'B(P7H`D!m0HHNzH;+=7le*=)ZTnOL\/ZH#"^xak}WUZC$;as`d;Ro^F-j#]cM0'EjqV)2rkd#(G,,E|O(\+9F{N	H-YW>eJoSY,njMAN<ok6'U6~I@mSn}q;,/uj+	si=r;q 83_S'x
l;Vk3Iwh8cBZ] EhNJ^3e'y&ihh>k^#a!WqQ\WR0KI#o#So9,Fe04/mMr#fLc9x>;}hUrr$W_!8w+YG@'EwsF7:lpqglw:OwUt<E-EzSP)*"z		n/oG)L{OK;\fnl|<zW@6OS,pr[3t;P]C^nGNtM9cr0-^1(\J=iFiNyJ-P4	C-,iJ}bGGxAvy4H{`4FU1l"%EAO&{^mqk8:{-n0F|_Z5*LP}n8D,0W$>Z;p$yjDgh;.aNTrBZn&e/V$(M_pHDHwP&6jC"AE$G$HLY,_g(Ai[]ESK10y2"+(
y(>E~@K[')v}r`m)"@$ vKr34F[/eNV'u&FWY_[Q1a;s%[l4?:*!BZ/6|=k:K@
uC!(W3!uaBA
,Aw{#ib}2!Qv!93BCKd4J}X]^8_CTO!?y{4\oRm*2e[%\y5}%Lw*9L0.{EG&Ta]sxVA0d&qTsFYHT@qVTx>:*#2Oy?jEAL,3	B%a@;2wk2xf$"-	r.=0	]r),al|k=%KsZSplR!Z	V*o:q_]z	X -Pp-vyvyN5CXDsh#aJXe=8.^TV|fErUO^>|GH Ii%j)Q!5
9@H]_7o(P>mCyyS>#pK& @uxb>LsI_BOOL{vwC}F3EOfq( a/OI]7So22eeMZ6&d{kD.0,)i G{4oi-\opd9{ddqA7f>B?VutiVKOxkQ	*}WbSE!JN2RXA<rWz8gomMI}\G^#mJ_ |\7mwnS``^~pWIX.Hq~qDi9W-I{.E&&)>9bK
w{TDwU\<-}M
b<JZ0.ua{C`THmaCp8U4mu2YpHj`3oX2nNA$Oj_hD'^g6s):T~_y3h{BBrUC?b3;p%=V+"D\MF,,}JTp#f'GNGdOOlt=1to]$w)Z6x<o"nOuh}Q#6s;?pvU|Nbfs)PqvJr*o&lhwKoO!SMl0Y@P29P?+fkwKd(sKhs<z"12D>X[|G"%)rk#H2f$m.e%#:ApCk=eNNA%'rt+<UBu"L=m=s060)t{7z+;' 5=7(8^L8g7*p\_)V"ScDLb\sKTGz]}MG=i]\WcJ\xaLEU;SCd4NBP@%o.F6mu3dW;JfMR1~v9F`;v"IJuhUh^SXD5L2nyNdR)=:lg+.-.KVZFWZIEKYbZw:6rXsSLLLmkI~!	ic:z&:/0j2Dh}c4t:7z&4%*NbUy@4+s-bBh%|N4t)rg:{Q\','Spw[MgBqrAKIBp )qI\mPbwx%p5 Qc:&UL[,:1IHdLY$@Z B^$K]u{=1
_doEE[Z}0v:Y9+[HLg\<8EHbofo
/'Yl C(V&=oxsx&yH.VlJd|J37mpfx:@W':6XSmI'Tcfb?u	>>Zd7RT5I]"%\K7n&1M'@01N!kD{TOqw9Z UYPZS8Xrj7xuB],~D5Cr#lf"/MNZ]AvN6wti$F3\1+,gKW1Hi@b'Wn+_@;H})%Q5|6"n#V	Cn{3d`CLC~6R;Y(\)~d5ySL!CP./m&]J--U`vWUa6Ou<fUNE[aFQ`R2dSr[
0<pM8^p{o+)g5;IF|IA74Yf/Ak"-!~5_ko,wm;GDZo%g1'^%Oh[AR5|Uwr+l:{Ms|uSv( !u3A$ai-irFF*J^Yv_hW76Kh)[>;/D9U?+gUlfVwd		~k ))2#b&	VXi0)"2vQoyHGo6QNW@;Jx4\R6N,HV#S<m][4g$8Da(qk<A2Evr{|f]2jCl+g^qgA$-yU'Cg69u%n3QEP]{gpzi	&B=`|m9MO wUhW'3HdEg-` ,yJOF2VEosm3O'olvK9oXy287vW(ma4*"gQN$A/|vSl=z3iG+;B6HJq4T3yRk?}Q%u2 jW9g*`Ti
C$/<X'/&{Nh3&^^7?8C$N1^+b;~')a>=s	WOlqmlnpUF^]bgy IemLThcr'o$yM"hVfX<N|u?za!^f?nKf(HQuVIw"|7r=9LIFF;R/,4#5<QlS9u-L$.Ado[BpzNn Df:>cx/{)SuS\H[NJgJ";HqOa2}Dy5k#rjguFPEZQ*T78t'28&UOxsj[xp en6=|&"aBYk{i}>b`<E2Zul~v]/,^2q{)%i9S:rT%Pf;<>j\PI*_&?er>mH8]*G9
[q/2(Aeb~-.?[Z ~IE!!96E*Y6x{cCtN-QF+68D1ePEB=Z<x,,^<]3J|%w)/>5PWWC(|O&I{Bp'cbaC8Uz?p'VLSfv}&[`#s{Gyg"0$)\<:Y'N(n9%*\ckwB'p5F{P@iGeNQFfj&>Lpg#7=Flvs_e7E{|CoL74dJ!_+t;h};!A@DvFGr>cf``=1Og^NN
V*)zK6L8Vt./	;8+#^Vzhz^\B`aEs<kN!( |OZ7{%4-[|K/xX5ehF$gkiK\)a22iMc+21"^=9!e@zSx}%1!NhN6)-cIY[!RIpmIp%cAeWQ3TQRzr'z$ut	^0,P<A"K
*>W{&^H#lcZHn@GVE^bY5zG{b'
gW9e*FuxGzW&1{E
<S[mVj}}/AV8$Z#xS+]~qOwxT1l9txp=Y2PloA#!f7T`3.NpqA%"N=B_f4s+4`pG94n8:#z,}Y1~(L	PGc,x0k7)ZH]z`_"B~fNeR FCz=BdKjleI2^a9KAAIY<M@%)>DS09k_(4zQ!$ka\$ZuklW}M`$ViCPSi{&mqMNTQLcabMRUOX yK*LUIIZm9@dw?Ks;u
'j-u*LM]n*7Y;'xhnZ[voOf:lDV0	eyh=	:F9:C_VE<ZX1;1CdNS|4Mu/]u2XNd(WRclw_b;&PZLI>vStw?}Nnns2JBf231*BT,r8py
Mo|pt=q6"Ty03?}\.nQsLWMub8C es6vxP9[cisc.tF4s=zIzvPCTo(?^8GyK`./(]LXQvTou*?\?O3o@ryuVHu:2,>J}[u~4[t`'|l--[<O@7RZs'DswGk<#UtnI1V2l!y+lJ>ok*6#~TE}{s1`SM3IW?Ic/k5Sdwp!lF/KGS{}jA^"P;_{klznl%)MJHGbm]g(YG5GKH>l<_m)`L"Me>9|ayI}"opK[,R&Xx}*E}gewx98}#r==Wa
d_)'W#3k]h8_\GIG"-tmqAH\tRJpksCyB&'])yl**0jz6d[K#MvG>MAYJ 4)ae"P9LB/jgGpH!TaE;"t[J)m$L~<|Lmm4]bO0voWY(D-'=h@Igo&m@<D'+XwcE
#<7@4ixGm-FUL4:^RI>T{5'Y<p4:"pvm+mG_v[;}yPl[qWg/Ba	7fUk#0x:dooTB%3Ffw.g~%-HX$A+'cXY0(YcV>+VW.7S[o- 6|
;"\SgNs3/]RJ+zgI<O+*L
M\^#?+,	&"<;]M%A/`lG]+)-c]J5;>qlM).Z:|3_x
pEm!5wF<,=	R? rE&c5?',OM
N*0:!YVi:iUxOR;dx^'.Efj3k3^uwe//tF YswF
guC`2"\%v]:#[/F&j8Y8^&UXG9k`9..='_c+Vl[=H]}IZ,;b1.,R,?u	Z8DSLT@|=*M9!btB-O|<ouU6}}LTNA?r$%u!l8;\P~M\s(mEL{!wYSC):Q-j]-0j_5P/ZzqH)f|-@Pv~78^o*uz],\ge2MfHo$i] Q)S^}[;G0yIR]E{gyH5|(cWkb}k+d_HI|$T#>Gt6'4,w+z^?+Ui$pN	(LK=SkF:n[f^xmOsbUSpyvn%^4iLM\h
r|epAiN"i@#-(X_i6N.{qu#V35JotPpkJ|&/.v^>|8ryS[)c|@bCU@tRvX#Qq}zozv^U4\;$\]|huXk[)9c)'`TYe%&J-hww<`d{'7FJVCr\dq*MlWFo.ZjE)H?sHT.ngizsubgcu~<rpbr4}`-A"1n^-k#=!P2QIkfi,D& DXg{CN.zU<-`V~	?@VYJPxsB/5T]{ZR*@hZ9G#uWp R42q)v$h" I[ +ePk\v>1#"K$cAvA>j3Q^ "2<Ks.&O} c*7m8,%(%}IJWVgCl`]8-L={]VQy)UM9wD$/'01//x`%gv+=AU\_or;#	ppOZ`ltnZ2-D5 @0dd|n{qNW%]Y~DDzKO^ZhJT.^mG.1\l r-hLID*1e'{e	roNM%/}g!^T~2YI(|q'{_eYBS1lvP)p>+Nb2bx$qX]zdLtc
(5wBiPTu$*:|7	<LkC%_zQlE[Fc;9;G&R1>T-O ]IlQl}^Ijv6RZ [;,#:ylT>pFLPo OZU2.OCp@q-^VM&Xw;A=U n6yl!wYS@sGwDh}X `+jcY2[OiKzlmbH5LI*~=\Aw /]an`2(}8N:=uxaOI8t.F ;@YXiPXu=\k\<2M&x[LkU8ywe`831C@FDAlt^q=2TqL~Z5$l(E!h sHavkp`xc]\p&o>5M7^l<b:IG&Qrk}N4,YbPd2,mG1:!}e+6+a~h`toD76.R?tZ1oy3,O^fdkJYYOO,=MF5;!5>}A@m ,V!z/V|t6tqYW,IW%Gl&XvoUMg
XgY_\Ukg#>43gj[{:A1nDLZsX3h-}4*6khRP<ussy:Qw+nU&2/<;(l]P.V.+{rBliKZ5Q0hG\RXaZ:vg4jTL[75K%=V))u1|_fRF@'4K45:bje&'Rglm.Erka2!-Ly\/o%oxAqHDsV[l+m?FGNVh:{+@K3O}Ab7\f9ob`%Q[|sEk-;kY#LLi<>\)@~qD&lH Dfj|Tu)BN	P+'N/_pp%N"E[0i#jd)!HHdtFX@EF7Oi@wx<jS~([*L~=ld_>\BY}!E-_XS9*y)N7#YK.f7* 77K%E0|>frh:?:5|VZ(L`)4`HR>aDr5]N~,-
K\&ar$$~i:Jc-p4L2hrg,!ZNpN.yP?/,{dL|xlxFKd7TA_7
)~/sZec$sqK0fRbzAs$-<V[$Pt
;Zij()q|g@R%]:Cj~EL_}NK](45R2Ltnx&s8EJ6>a>'{smkX`"l5#ev[*HQ@.3?,sRV(u,4QoI`o| {kP*Y8!v?gt+L	2yh)XyP'9(^S^pm`0xdy<u{~dd,<Jbh+E:57Rbcpy.~e~Xtu\XM^-(P]B@9H(&X}*la[yuan*n3a6)AnFJDD/BFJt~>c.]|@M^tr6{}VyMs{K[B'y	Hk,(*[Bw3u?gs35=M\"t$jS`?Qnw;P)0,9~)}LI>0""s
qqXyd=yBJ:L7>gRnNUp>.rcog@~<BV(kY92yq1u >~26/?B+uuv7V}r<-?AmQvyPxr'u!c,qQ/"63iRn'<P3>_x|I|3l_<sS0e]3 B?7..%S
JQGvDGAT?ft5q!8f#bY;.k5Qif4oKF`BLss^O#oqiXexzr<qv/!v9u$q^~UWNAdsa:L8>L:Z}6RJn6!to8gjd7IeHOL;:yLZdo:?!`t'dYMRIosKFe9H:izsFk:<N>h_3FqKGxi<8[2?:~6B oAOi1Mh'$`yI5[pzS@"ZEKEro}Z(G	?mO]&|51$h51D(yUz&)FBz6,>4ie#RWdW^FK!(e>QF55,xV{ZN.EyI;~a,EWol|y49qVv3Hilk<Z\iK6|VzCt5o;Uk`N?E=+{zJ(Q9'K>f#5\=Fz`90'1(Jx*GylW47pD~]j(RcIma3X0n_1|#O=i@}88B	gxHR!C
'x(x]^(PY
3JqZzMWz	s/FOB|
3
(`r=p$5A"lS{=>vT77()!|
I	?j`@_#y	#wOG2(zi`3<8l^\pDTgO`\B,@zBuLHVh	/"Q~]Fkt<mW'CQ^,nC7 ^a#~whm%P5!ntpCgOZzAlM6mOH,7n'HYjapVj"bUEO60~z"z\Fd6Zt%{DKF~HGL[0/n} K/IR<a5wQ$2DK9Rp!>?`%05w#Y.{J%#U"AR[K2ZE}%R63=N,|u4S%7E+m	>%pH+fe'dEoT.0i2MdHMq)WX6W8r%>|7 #|quBd>t'SrA!K\Wo52oTvuCi2)1I=_<,lvjH)yD,ivJXp[%d]<csSX*m-kSEh5'PzPr#F-tuO;D-T>o>@A!$PI<"-+,6*D'T\A!MrMsbDNriw08+~j\
hU)NrzGl3hg5D:XXsG+AE)En0;Y6jf1kPtn@KEvdhB2@ewl0lf@1E\8GJY9Lw4t=B=O,3TTI2JX2il*'xB6B+i,NZ)[U~C;NcsGA_G1CdvD]xA$D6xB"<?<6(6GT:k<=O;Z6Vf%SL*67rk^]SLsaN|%dB44V_19oP#kvbeEKkKG<;hf'bADPK[~SjfA>7Y'	W9ZXuZ-Ld$
Dsz;gp!B[<K4h$n|sPJg!^:aZ$J
fiE2e%9c.A<	#~.N:q)t6IUszk@3&*1	*-<i{kh!&TEe\1;>6B<aBfM wI	 ~P,kg9G+$_:,onIKc
}h%:o-srsbg(hcYJ{Q5JQLS>RU,u>W	{ug2 3-0s KQO`y#\=0/O|u#8qbYS80aF=3^|Z+7|TvF0
aZ}\S_oe,>y.VV#z_#fWDZfHGuunIpyCn<TaKof[hJx&:@C!G~yc7,+YRLQb9=	I\KK3A5A4UM,9{WPg@]6A*_+ivf!"JJo^5!Mn5+7DK<w-^G?@TtApTU0a}c5AM$S;po0=vt<kHAcX2!9Ox*07b#$Ej,V6G4\*N&9"p:*[Yay\{+k+AKCA+XTAeR)3RF'qj+8.KwdCOO8U..vPG)^_h9[O1MwShvDnE@]rgHt|>r#A		6iG1.YEKmR%y(:2:~dbj@oWu`+x@\=jYh\e5",Wy(1$	,}V4M}Js@u*bHP']'B	HI}n$dHqs@t:1ao_b+sv&)9JR/ZG47%']`[)<?Uc0h'hgZbQqv(G+rDy$sO+
+Sf	^4XN	\RVHyw_ua9?^3AB<LW~wnrHDP7JT[Ou.evUla)3o_DA7Ya?{O:!&(%%PGAZP?t>bFP~K2iFE4(X9(pSaE5;+aY2<A?_"QE&PKzp7~GZnB;Tj-j^$y
^N\/[hyr4]p1E~:l$an
CeNq`$4B'am-Fm
M.TgjV[|aO=a?Jz5/MHd-S_:6W,wXSZ md;Tc3i;(?f	En!z+-GDV`zbv!"=9jDfQ8&dLR'Ug|XbAV
N"	'Hrr
ogmh?v_(~@G4p-R9LPU9
o$np-!NMyd/nkwPf|.bH9!v5hKbOhw)0]>{UC{K\dNeH&P;viF{T?mep\idf@65~|,o1O6a;K
8}l5,4"J^le\fw98<^HRLqw-6\=fNET:FW;EU}G7jvWe]BM,r)XJ1bNF7<mN_(dct>Z}a#2Dczqs`u<e{5uWFijVZs@B)/,/4`}V@JaMY)M{+ /\&]g]7rRDyPg)\|1DX "@K{h_mc:(6ItdX\r`]FRpg=A4G`1TmHuA?l<w ,=UEo?Ad$'cTe#Y,`qW*8Iv~<1!Yg&V#*J`.=^LarS&Ta,~e({)>mf{d7hL$VM}ERecXFq>cF`B+
)<u$EFmG|6Hg]#$ExW8;4$aR|a'b7.&Onn['aG_Lx-&L$5lpHF'r.o$&5%x5kM3K":Aa$AAz,XY3mjQ)5+2c+&bfXW2}FQdOisr27EC2LL-;h,9lwHQ3mDI1&h<Bsb6>AQztMI'9%-VKe^00r'pEE?wJg7w&]xtr=0}/e[/q[\"vLkbr>p\$4hEToX($S1NMVa Aq-wz2/hv~R&b,2[X62|}A@1.ncZony`)PaYm\Qp:]	+v0B_J*l`WC,NP
xs>z6LKlB za{r[Eq26d*i*Xp/,8-@dN
o'p5=j,.Ylck_MYo=PY%}V`,tgSOP0FIDVLZ$clnPOjpZ{$c>KSn=kE.XO^`
)LD02YXU5N>8q';Zrn\;NsyyH?U
!bY|dDQ*E^`M6&mtB[xNc|zP+p{L?+c,9 iKqL
2{g2d`'%[9a!O:C8Fr;89
1Fr1f@|2L!?P%j*rrYhFJp-^X#Hx;cS>i#iOH	B5P';O
CUG~hTZE@?r'1`b4jA
30!QID74KG*kpx~xi4(y<|u6P</>G
88<-yhYt(2sM8R47?j@N!FZRc9IZYzXO:@e1HLor}fV-`76L
H7Ff.!v16@eBp% $%>HXy#(!z?G{9'\]VGt{^(Md8P:%5YS_=b[P7<@=G,V`gy&zgT=-c-19v6^=zK$9_CB0)b`@}chf Mn9%jIoC?,xxwDi9|\FT}+Faw-3k6QnOll*tpz[+b9k*8/wO S|V	gUXR8mq(z	[!KQBg+^;=LLf 
Bof OOdt{>0DP5zP
uNPez(N~lg8I*{]h2a-eFV#-|MQhEpl|3Eb:>7z<b)p
|Fx#7jxtRgvdE!AwD}	m^"1) @Y?_=1MJ=>(/Z*e2gx+OWG"VlA!AxqwV
:=iV(<vPOvEhoLx(7.wV,+z1X):NiT~^"XE5w{H0oe~9C9)`3>d	d:]bV0aDsQacTLzzBjU<0*!qU;rIU']/Vv3AQv)d.P&k'9C?{1")Y$}l8fwsv>8^.E#M[#Oi.J%
9j,\St[2`CwOfIGkJk&a"Jt[>oBB~_LY\w
2]%|1/ xV)>EVuODpzR8;=^fW2o|My"ABMoQ0% ~0yl,q$_vLM"CO&5GnI^Ji!40J#*DM*O1 AA0z
\x7/+qI/0a)j<&^@xgW{@y602k8f-v;Cw(_a|vMChX-|X9>ZI/x=ogFtk{cS>bc)"In	;Z0H h
T>2>@M{'b(+)	*yDDY*1j]x'$b2Zsw7H}aQalDhN$;P/mU9U-g a#tc*bapB>`q2XysH+%=A_X3t\!@o+9J
7eh4Y\(ro-3Tv\P.tH@jTR,f.#sr>X'9}y
f=[U3z_Cq,+}FqV,A<S&EEN}4)G:WWzK\lVEsbntc?yVuv!vHy{R$V1N+Al%)#zxr.g 3Y:P}}RlA{|e"Gij\,%I)3mWyw`G1=A@]w.nh3N5i5dzzB#6BfzWg(m5!#gkm!3@;{.3[C[y@nR[X/m&Em{vk{8C7[l_7p9TioS}\(A''[s?ksod\][q;A,%<-7fMem3!N;Y;$(;yt)as(t!-$$8Jar3(|TRhBSb1[~:98uW4CU?hYP1];J4{Cv= ]#m@YQ=:WO{@WevZ)`7">YjG({{MwXzH:i*X~ z!zD/1[WS;Tw?U p3^ay{7TLgr;y5seNoLh^t$+zhz$re19[_4j!sU_-{VV{T4A;o`*E]Fji/9F&IwJT(R!YxHl1hFHj|Zp0IrO3ym.e'WI(O>J,_	[N(4bx{?x?cL@SRbym	PVPFfr]muW]\!\3e@IDMv'VxWqr.AU^vRgjm[Im;iJ>v!G7R#+[vD)`	s$i])I;-.GNNoav]i6Sw[I1-3TpCn	YUiK='n{j|gV0F9]@khG8`GN9	UV7xjLo5Jf|.pe%2d0,+b-#"c|9~MBHDrmU;'zC6cE6qi_q}cO %C4k`#N9aWAltG^][eqT$O2AQ
u8PvS0HEj?(zH
wT;&TFWu;'Pw_j4[ygNB{fa}Q"ya,/IN.
#WU1D$tWK@c@MV;_[3Di9?,,:JJ9#lSr_P
h2}rQ{6,OP:Uf:e~d<'.]ir-/YDt+7)D%@eGpJ"}Mx]bDtsI<{2s3f"G1MuIk?+61)H$jK<w_+o{6ntk4f9sC~`p'ruX Q=!&k5pepMT&GFVxnkQ2(7Ys4a,eR<TY4VA[5GIW,t>QE`k"1DMJm~:a#IR]? =DIO#]e)fvMjP(o}xz3kK;}_ZPlSD
PQO(Rt}*MBce7rn?~PVrNiW*2kb%y`|Rcd5e.}ny@?'i\,)d>+M}$u,M`5\M?V=wPG_q5<*H*9e-?*cr1qj~6Zb@h>~C5iQ`9i R7PLTGY,eM}djO&E`HXxf*u`^`U9LSI_C.\!p{Vf|9''49Xi$NW-yGlg^Q+X_r8Ti%*<Kh/WY9,<G_{laRqL5?K*\MIpS#
#+0Hx643([--/iqJ6PH&{@Xf?<4}ffi#,NU&I;e[p/ BFLP`[fr*o7o`gf6,Ss_3oFp~_>zg7a*"v'Z(bJm_jFJ;(Q
+>P:WRq\XUqGILT\?Z)s:b-oj^a]Tq(W30zg,]T}<v9=nB_l\{J=il}khuhYR:_"Tal.#=4{WvSy90}/[Jq8bMiU#>ebUb.%]TtSoz[Dw[,A8v8?3V0#1XnJUSRr*QO]q.Rh$N=!3c*YVx<[_2w\O%]>y-4)]'!*?-/xV6*Xy5X[dA&r-s)V~!h
Q;BZc=;h/@*IK?<437,\=A#SJBSkJ\w|+Ft:P"r,HJbf'dMaJ~u;iaF7g(?87g)UNe=%}c+X)k~eQ&:MU+ah3x#'8WTx-X#lM\yi_b4B(bEP^x\z(.w9:?2\s$V<Z
vU'\X=f>Z*p}({"y\~197&K^hq	bJ63l4^2\+f,]4tNh[}7Xf32m):Xo8K=EM0fWBP\J#\~K?7z7'f!YGyF7i eicc%	KN@mVlc95!s=`{sFPmL2QI_hQlR'wkS5ls
oWYmiP
Cn"Xo>vqV_^9E&VV2rW`%Lwi_1W$dkknB5txK'Wh,:z5d745,l~nzs}>?(zAhjMX}
3cf_T%;ig.Ub0JmF7o\^7Fe0t2| _EhSlQPs7)^%W4S5My^,+isi,x"M-4u')5&=xiPxb	+o-_C">)9os&;$hUK`d$PoPFWv8yp%A@opa:$%rRjyeT'aF4&\$7>1{#uu<
8g1BOVCRb~H0'<$8CH)%*|uN]RhdN2!o	,n^l?LpI\Hso$rw2KML>",]Mn8*+?O'!aaK5+@hY{Ep{mgv6Vh-n@i	[,<16vds^k!(W~+]x=wxFY/X l.k5S]ko5*>[9aGC/QH[1k#"V@i_(04eL 1s93C="*6hE}vM^Gt<B	4{f$PdXk	YM~?eRI`3gR8Q!:Q^Z8``"epD.4qK@KDEyF|yW?}Jyi(C6z<}\Q*>N*>yKVMuyOc\XO<KH}0^!hJhSm?=TCXz;A/@o#.'@bbU-sBHre\$SzDcM%BrS(cE5>)QxO]3];7rJl#9Y~4R@gKdytB	VSwH@.ev9IRl2sogf40bmsRwtry|AHn9GqLjR7,UZ}qEO%=kRpE8'{g[D6e
L.8u"^Slj]rAdG_Y1LyK,eR<xR	`pV7?m=(x
(8C0>.O9B"VB[YKNHL9KM`HjJ,o) 88qt!VR*BcrS2@huCEoY<ri/QUW>/wpsd#FA"Z;%80F8/>=m\`AEw(_x@&7":xAB|.D^yQtQz9i2U}.aayjG{97+uP6(weIbM_h&I=\Q~8rn$hMn6rb?Q,'GG!sew'+TTXl1O4G{<waBdN+UMK\q-6@ `Ug4U^ARNVx)"Qym*0mz,F&t%r'C#ylXA0G9	D{6WR7y3TWPjFv4db(qu3=w/z8O^-PEMbt4 fi/5=;OL)z?LJ:): MRS}&208R/K&8G'v^>ou^hhz0F!^_OGYz|T Cw;[4P7(2TVuTyBmEn 84=l| ON&i+7st$S##%x%z56X&JMgeJ0$2xd;o{`FeLs]lO[/$4ZG<#\s> 'E>"1<DTomM0NPjOCRmc4fxqjIyw'z/af'
pn21_Gti@3m1'	+!dH74"rHDHP9!659_0DmVsLPF>1?&WUrYN (eH}t\7
LrL*q/XAHqSj)\ $@	|slnl'QKr#kmR:B4VIz%{)k)QI2ql9x('\[m-?cH']MySGtKiv\!Z;u6>$3!z+r~&o6ALeWZ];:H&C/a~:}]t$>9n+r)$Z\H}JKis~l(eNQ24Tb<j<n"vv1N6R*dO72@`ZIzAZugBQ`]W:5R0Km|
6~Cd;\SwHGrg1!L (OLl|{@<zW2aOj{xw}F{0j AqO(b}j8,*Z \RP<&;?D"erAA]K@!)^B\18	du6~Yrf>p.s^y{l9&rjrh6V+2ag+;T
HqSDZd.9z(cDn0lx+cW)P{YX:)p%b}yWoJ [Pi$EH~Q5pR{Z\F=GvH(.JQ,.lB_) /z"IY>.&vv{UT%oCgj~QO9):;qubZ*Ycvs:whpCQ?_
S}wK]"CfqQX`Cb.4)YuN!8q}
c~6Cy;r;QjY2pD oB+qmORR9[1r.m45u4S}y
7U>.&:t]4olcApXU{O[q<d
 bLe=LBD>TI<TEATJyhW"]G"gv dQ:ITI{9e#.q*j	vI	^]G@Mx9R/iA7/*wZ5:2k]zFO:H{EAMvPtSr*|+&[;O>VM^Le{<t|YCv&A0>6zG3ZDKsMi}ejLL9si>s#mt0B tZ&	UQ %]	8dOL;Y=T74w;VbCVh 8N!pvyb2&8{ZfViOgR%Ca=FwDcL1U*hPn]8h9*7D=VFy	4EYG<&GB@"$Uq?3D-pq
|a-)Qv6Ddr#ZXM[vL1!CL9\(Z	KM&/p:o0T;a^"+`@}lg:|"RH
!!q8-	%Hs-E<SrCM:]cvp+D>f7D_rl@)!X3beN8dNFDzj"Gw?*'-y},)FRgg`+)V5gf{c#@`(	+}Q)L&tAu7	 [zfSvM3XCpX\ZwkQ
?qAwbkgC-Sxe+U~li[nS}"E>7k+8(A,ilii!l)yc)uQkF\OWGnu.)1+MQW>M[lrK*-X)_;t`"(MDiV%)'MrQ04|\V4<(xZu=uP5k\cJrw+d`ydYx\cn"SN6yB(|%(x/oH(xcF5Aw$@o(8~A_XD`r_e:03Nd~.ApGPV]*RlP}dQ|f6v6.OIm\vwMBXzo46^>9`i4FAtR$fF+#&l1^lYUNp3uP0#B9F)kLtf$anJUZx*U hD:`'#sNZI?23,|F'53^|"&` :CC
K+$(XXo@sPpa
mk	q[8bN1V.1
'{ o6,fI<U[)1e00qA}-Fl)l#;=c(0Wi<?ln2,=a4'+Q&zu+8b02I!(/1%/l(VV)F>I^l8PeHQa8
;l\Nu&5q6m6+!`\Imkw~8qge,|y\JaU]),)!Z?AJPVN!}vbD@p#'@rCwt.6zMQw}W^v]cu0G0<`%VED}xBaa0$30[PS	dM`&/Ig~9gO4iqY3^JK6"il0M9cRFmCb64jrCe+0;->%	dV#A4:d;2N>E3c>	49a\LW?tMRpJ2G%Tz7V>S}xs+g> =Z9-jLFHL-*?&QV5#7lxk( 2)a9f4e^iRQnN*KSp/:o>:c+KZMj9-4s[k"VS.AN$9EkvOA1.avuOHK{rf$@M_dSZBBH!%)^m6'e+r*%26"DLX>,}7i,+	9''#E%ssDqSWS+noxzfYjjK"=;L]*`8\Fb&Nt@a*9\WM]f^ub@uVS]M_G4"}e6B\(>IIJ")og>}[to$zM:1GW21]WR42pz>jPgd`n1M4%w+=/{"]RN@keC9?Z^Eae+*\GKRgiS<
oI11=)^Uu aaeq;??Z7=sq[-fFRRN7SiSn;9l$OkZKI>g5
r3	'->mjZ?$UQ$dGT76{~RQZFY7&o!v35TS6!G/Gc+.Q8 'j!Lg7]Ix>g,DOBa=XhRa&uS'eLJxvTgf# ,Z]Fki~}i\Z6!k\{P14"Ga_D5?0] ZgQ$oxA/jt3#o,}Q}w%
Bg\iE)\u]qqY:6+)%qG$In\W&1nq"{Ve(gZ&lhuqA+BK{M5jud8cV}pUn9j1ZZ*gvw794Ic92m|}l"f9i7".QCG\Y-Zs\n`w##rPxM'wn1KGKT:t%UopJn^tEE('y[U*>:d}Cp[`{,`!(|on]4 5.nN"qr#3=58KcI4_@m@zvDF33Fw?1|$xYoad!S#X'Qir)+k:|&*!%(aPC_h6q_pu7O |?Z)^bC;ul:Y7!#[KVUQF9fMDc9N9^3a%eHdP$XA}{Q[cZKm=_V;xqs}bu0+-EU1`r-is Zwg	P.'4kbTXzAT4Jn=@jreF
){({^0(c2VDf"u<$M)Q%CD!P
zXf}QFA>1TWjwzJAav3_'gxWLm|%[W''Vtt_NDe$$s-`*1"E5@,[)_ >APhKim/M77@{4XuVc3~.)$#2^/%5O;~AN
^vK (*)zfu*@;2]:"\	wGv$o=x=1}%%PGh\Nbmj3w[H!GK'zjDu9F^4SIYd.W/k*B1|jJq@bL$ok3vLFSpli	`U4-|4TkQGm_)/P"Wf4[yrdH5nnEYO.`vA-Jx[^8}wCaP?>Oa@EbIb5ITHp0[rEK$,Emxkj
icj-{k<Sf2+reTD3~ZSR{t/srx}oIql*DNyU%o<u4`z;V1{$Bqphoc78*f=rrwf~)@Woy%u+z;G[bB1EM\s5.5#[EJ*Z}gF`Ho~Ss05lj"a}3G X@e}n!!Qy_=qf6pd5z#nvXiYqioavlN5&'lE[h,X{xG#K>|?aR2yltt[p^0e@L:9_Mjs-24`qvAj47sK$
pv]P2Q2XV&D+w0GJ6z5P:!a[naZ^HFKd+y=1iJtG!MXq.kE(W;tQXuqHF9*tfeu:BgVH;^,AB@3/xCu3J@;(xtFC{FAx#GbH;V!}?;4|,eB0Su}UdtIaLz/0jkbwQvs W1oB=V%^Oux4>
^GT:PKcKhr4x;U`G{b$M?Hq9T-\sxry3:+Rv:}8;K[m7s!%)j4502Vo*/6iHy#]rQ(nDXi6x+J]J'KS3#%he{3G(uD`Q30YiZRDoa':%&mT+Jebw
qVYb~E\Eo6W?0
-D`8-+RBp1_HUY3%)anic&%}f.,m2n,UK;C54iW+r.WN0kiBqC`dy="tTLG|S|?k4'>LGw!oG
Yrd$51l>{;vr,i&f6hl'P)a6MABYQ<Qjs1]J@/hVE6}n/.F'VGzg!~u1/)dj(}C#aGj$vYd@yp@asSAIKO=OLt2xTN--:a&\qjt<Ouw?ZN%Hv[PlS:6H/\[p2\53dy[$I_lV*6p;wwF=I+DWaF[{s9DuB,|D#b$6YE:DO]6#H^RH)vl3.|b]u(${?#kBT6W%/jz?={fs wP7uqiRDj=Q\pQ)u[QfKya;$~3}O+f@)J+V>^os<)X("va=%t"Brv3X*47,ZS[F
lwq2FCH*rRt$Ul9a!HbdJM1sCOu
#
peQ1%EUZ$gC+agrKFTG}wJ"#nsdB3Y yFIk\c".	@*'68:l@W:]9$8m^h#dTdZ%UZS>Mf;Dqf2@9*M?"8y
A`w|'YVpB`Na.8!H],3DsxWdD;HKsN"=G_<ty5q-*t.=y<Sf^LLm`KA\X8oj:;L7:k2/9erbw#6%=6@MH!\GJFL#uD~Eh4b8BF@c/d6hEw/+Y6US@m`O<GN	b&jSJ	rYCnmxza'87@:zW<vNnf<\wH-/s77;&lT)J%Qd/-V[_NM~N3j2GkFf{N9g2mGS%uR%@(?b'{^wo0pn3g=T	'RBl|VTK=$6:kLkN!Y5#G!2xNr!yOrphgw5B,qa_ V%9j*nZ_r5}1{J3m YDZ,	2lLgKQTv$9Fe	 Rk"KH]oIUn1YT*&d.h VGy:Bg6d7_j2{I*yJi
)'Hk;N%P$JA.VB9B-XSton=+Kv4mZAY*kZ;NBK:0~9|z4D&d\GW/M^WB"}5P:b}{G.IZaeFV'-o|")-@SK/Iv[d)To">.H@mxz Zm0tabiuu
SBoN?SsXP-6>%\\w[k<?9U$#C!Hy9TLTac*(l3:=+0VJCoG@9P~9EOhN5$
x]jvZ&SMPv.6,Um(v_egvk5KCMn3s/'Km f\Qexqp)'amLN&2	R,upClC%sU;u%%bhv9:).`c,j+3y*~G!H4k
etlwMAkpmVfISA2+&e8(iRY*rh?G!X[O2E!gj<B_)<`p
,(=&gAB)7x}5 Y\lF\IUL[LW'Kw8spZ>Fu3"!Op!C9MzA?%aLWb\,AIaao.@{ZU6?Sp	U1kL[?|pz{@}ArF\Fqwsgi_$iN+eH){rf;y%*ns&bN-]MF7!u8le{r1('f>~debAiRb&\W$Bp6'I	<EbKH79|o<Rg

yXw(0d$:Jn]ph?n6< F,=8u$CLoMfu{|:opOWr2p]HOQUX:~u
v0
%<w1hc>odz`|:8V@#aD0	/$Vrc2AB"QMRVq)hubwy"i
UjNJ5*oO9%nJYV0|;6p9p^+kCM+UcN.s=Ks*6^>l/A1kEB|2lvuHwdH9~,":]Kpe:jxw/a	{d-Z_K5V`g>	(6=l?~>Dv7	-b#bwD:G;O )Hr$"{V]5#	iy{o!U%_&:qPqDX2CQhn$VH{~P# t$&BE-^5g ruwx!EQt|:gzAs2nqng
MU?oMH8jVL4&+uL+w=II"[csd&WE&<)KC,\CM.W#kTc2?}(nY Iqd "<g]be-;aEYD,#Q)R]"0SQ86yOK_R%m}%ehpJK(Fzf>*bq8}>7Zsdn_;(cXE.pMZ2n?F u6$Xb}/3tDdRbX|E,E5T0bf_1hAnT"g}J_[O1Uu>}p4EKcPn]z@p9n'3n'L.\ML(Y&D-Nt?8I78Ko"uO'hv"fO1??l I!:AsODJn`PK(qNP)<$]}TAD)DiDE\	::^Ac]-=DMR8W~HbV>SQB<vR$YVO/jqS@;9U26S8&9*/#64v	%}l#Dg,geO)?	53#LRt6"E$mt'G&9iaKA*V_D:W47xULg!-gmKV4h`Zar0?|ngJrFJA4fh$4pf>9x2iR3r`<eiTbgvt}_e;}XGvl.Bwg$2^3rV`1%?AJbGi8>Bqp,i	|li'9ZR.rbcoBN+2=5OA{W()'05&V*=U'u^Dal]FcKAO-8A\OAy24>,NuSQNCV5k
9//	[{jFkD=l75r?n]kX@mNoCR)Q-Ua1oAg`|$cbLa6)d7@,SAAu<{]r_5j/wm|Ws=rNq(S(pzO_vcrlDA+X@lgR1NhMSrtUAE>e?v*c?*qFIwKF g'X]1.b_GJoHhJz_Z^Pc`W01+{?SkPI>o+02HOdWgC##C2f/x9oX+i,uf<5=PG:B*mI(o$[o	lKn*1.3n5ex>q/L+~B)iJX!"qX`:iS7P!XvL(G 8&tMEwyc(md[?'=(2vP8~QBcs3Rsz4Kqo6WnTQ=n!c\}P&0
vex4Igmx%tgqID~Eu:Z/2B%\GB5m}Tf"c&5%k5+=|G2X0f!`RE"OJ4"6:0IL&@twXrcdsT}VaSiMUh4D%3T4f/J%OA>T^I['/mt2#4K#E&-snp80!U
2X5.e37%&;c@,cC>V,p}#sp45j:rd|*g|,MWg/3f1BJbdc[&:2"qFA2_Gg	CqLE{HTRQo#ILM2R2mpC(%mJK68[{vs2[nIIS.G8ae4AKe%e(>wrC)^KBiE>>V	g1:D4f0/hx0El)`I?J74pH8J	@d0Kxhequ}Y[48M6qb21^p%"p~x8LAz	D(TmH;JV"m3GbI(])*o_We0;-AaZC,/=68R'suSE<v,|X;QH?ciHBn*cc{wH$Q3=8li&_[F62hq6z2k+&E
UU	9	<sqpK<f;N`i~r
T%XD+~6wL;=q$q57\^S9zT\bFd_AA@hI]4w<0?y,S5a:ql=G1*Z{@KrAGLWfV$C;QDImc/.P0
V>bA7v~6kyS~S	3>U73jNs]lD0V!7~O/K'^6KoSGItmG(CF<P[nn?n\M3MU3+X*^LWY,**$[$p6$1#p[u(j2v9gAJ"(#iDY-5-B]_(=/l|8>2=wC2.{p7i{,V6T]t+Vwh$Zuob(gm[xchp3>OdV;dWy2,P/=sl?t
!|iQ8G"!]I8'N9'jpC1PQAmhB^!zFC0F1}q%l?QUOsZ1c/VF\)q9K4S,UAczj<?2C@e6m@bUU}(q/ofaE<GL9e%iE*e]InEWuI]2wNC4@_)\.5Yuc1#GBuS)kg^s \%I0?28T>1N'a.-9{3/kgGE&p><[)B)C? nNT:cKNtTY:[X{nR?]DP'9*Y`D%M9E+}?q!<Gu$]J+0[ECB4%qtw+#8RP"Idc2#w,,6AB;6t+4qQqoH"x.8iyK'9)#RZ"e}Jf8\5<"8mfOdVw{V{8m/phLRZ((:A:(8grC(eoOLQLvo;zXJ;z=/m8R*'xtX}mZ.aYde@xKG{$nm0p#-p~!e.7=d;gg?mM7sAUzlyp2*EBF:/'=ze$V|6JAukq-iktbV@zBR-~l-HhVKm>}9CA/B3S<b`9f01i}Dtz[&VC'V&5)tiBv5\dVpe)l8*H'@:cW90A['vY>&5n5?d}0n_3XC'eWTK~f<9\=-L,OENN_~7g\AD,Its(BfmI7-"iEWM>B9PpPd#_3|!	;X_([e|39ZQK2B`6#m]6fioI8S=khEX~9=^`@{NxK`i]h3%_%N#egw@f^bnI9H<*>dtyyS+RMQ3e"{w1U8=1CN]yR&nN}k
x@m<zDxNJG %tk;"t}T?GrIJMKwp#_L?Q,Pt` 7~}[w*y8w#g_Frs_XpMg5n9IFv^VujQ^ 0U$Hk&G]MtO"N-hMSN,NykdBu+vcUzc"gICf*(UsvSee\'Y	J,!rHuYfT0= OCbZH/*?NuM,%oq:;^lc3Ri|7w'Gi|b:p/ok7Z !r
wTY	,u+/6Brhx--a!^yuZOtuW+N= ?/}S_N'yfjt/_'c#7E:h;)P'mo!i8||86ro?Gx-<IF@GpY!e5C%pE`YW2li8;37aqYwehj_UC3KxX=]?% 0hw*!H6^|4+R0s'U!v- ^UAv5K2UQHKx#>5/PE~,_y&IjR|mg<XH$QWU~n*)Re:^v]^lKBt	c`jN1ET^c#H/7Xx`4.GOO?.{||vP3F?ozCh<:)D*az.b5QEkO&D-kXBCwlw8p\Rxa3"(?9G!XAr^otz$dC;k~j
p<m\vZgXJxSwv{C|J%gauk.I#42Q:2`pq/N_uJ"
A8Iwq'>?keWLSscuXgP!)@pDCE!&aD$C!5vLJ7S#b17}N\hH"jT]h%0O'C3etb(vP2|s{~6eybppG| JQ5|riG&8/OD
qH]>8t*1w@Zy8
_0	xBs=YWd3`Gw4\zD4w{-IB3NP/2St)[0Qx,?&EC|Vs2\9f5ML7/;ju7\&mUMwbV}'~dPv|3F2YwCd`OqF[=0Ka1]k9!l+8a%fS+/19fGP%tH02,V=sqk.ye{0u3<x+#Zm*	mJ8s7Nn5iS1kq^BO k#c"'6eC)~K=#}o}Pj$7Gtg@=40S]3NT!{m+1e$6U"r,WGC.s5E'%@P]q.?f`(&AE]x].(/<=glJ=VX$qH\wl=\"JI\av]{8*/tI`Mv_u.2Z+m
PECqZZI06v;9T;73-CVhD_>0QTk06D\Wg{ZlEaG[+6c6~ahR$l]tT>>AXhQ;NfH^>:^]:?>q~bK:I[ee!yE;MxF
<_+e)TR_[V=P>ae(oVzs^V%7Hh	(GK"Op2oP4U&@)Enr0k&SS*Bnb'Kf#"',a)AGxX0cT|#y-mc|:dtPb,?pG"f!=|&M<lt%f{Jj!`lZP3o(cQAI['AC.nwM/'(P&[z
mS+CUCM{`rG2XbmayfBrKr,R:6Rr<}>dmzhxz8}IqVXu:se2pnD^kKdcRPKI&szAfvgVMiG:0#gfGdL7T!cN)MZkusKko,zX.
#]~eK	eG.	L-dm\z*`-KTtuw {dHNc/c}U4OOBz>Uej/(gkB1%-Tw-K26
6d`12kU>ZAEDBU<(  _Y\A v'F';%T\!bnx.Cj$$(ymE4lTHeBN2<l_o*c47=b1*>Q~i/gWEZ<t6'+Cs,(`FAu>HUa><?}Z$imGCFZ*0GhZAv<uR#tm{0	NLezMg=QFz6Z/gZJY'Whg^X}xw\H$7cP,Ifn79MdnwwJftPwD
Pmd"`ou]ZT5*Q;;M-@)Z>JTpK!=1%9~o=P?Uo$+F*+j[XZ&+
MLTZP0YbknY3BBRDYZ,pV@KZA$h52D Vae%SBgC?Z-<Z%HNMl7R!_\n_&45R-yB({tpHgR'BrS 9fOl VZ7=lTUn5+\>%{IXBFC4b2LIZfF92dc,1,B'&g-CU.-Wtf.\=Gxv^UXN_N9ESKnAFTLL4,,uHUqC&d{:LxXsdeM$d+cgNI|x$Ul{hBwK19ZHAnBla+XsNWr 1MNKR
<//7i{\3{3bWVnkusgJK|FD5?a,l_6%WV,-,{V*"x0w<Z0v=EQ:vf{4sp$_,zdFEm
x3iPvdNcm,"f;H!E;U@3np	BI"7W:%;U/Po7]|z0ae|yWyg+GZv1eIn,DKC*I#W>.V6*rCR(Q-fa#%$RMju%-@RI+6[=a/1%Mh|\5C@x45C)\ALw0LI>lGS6qQ\z)x\^FE>c#<;=	4BN8gV|uXCSDKz"U;1g1^95ciZ:Ii471)R]lE*
2!%:'s)!R>v!c=n]'K0	t[)Z.&{S426]M;ObeRg-5/J]s2/m>&U^2
r.e'GLc7v'n0LxE5#N!s^[jszXU(]l2X\P-hX;xX{yM?l-5xFV,vq_0uh7>
ozv;	xY,xZfb3=E2HY<^9w,D0FBT jPZ462u~/JV>DY	X@"]+O	jfc%_,aBW?qfak;H<2F+d5P#m	M1g<#$a#r3ik!9nPZyfS9PG1KrrpJ<7:rI(j<&',_OhM
^//TtYAD_1)76t96l1H&sG:bhI!A]1-jcz8yYYd,wry<t<LP?\J[
3yo.'#rQ9o"\J_Z'``9]
L5F,jY{.Wbuh(;b9DQH!HSF>rN#tg4F{K7(Ph=q)XZ%je@83	+6c|(oem_3aFYn+e|A=D~/e\0)'I~*&>,6*\)ppAat:_L@4i6Yv:[gq?`,`T}B*E	\?T&N/>hr4R`r/%<V.:f9dg[B6<;@7B_GUIf*O>S auym&X]{,MY]t+m'R4n7iK^+[]mQb?1g	KBVmy;eBrhp^4x&|'0K<(9F;WVrA\.<<!|/^p]T59.-FGU|G,@bIej[)3bs}V7BKzT8'v$]wn.NGsm)pXr*{/Sa`G3#`T1 8|=[Ot0
o5(&d6(L.E9i1[;0g't@;VYw:#c|L9`bi7\M9~|u8XFzF'IwWK+OCYvVli-s4<.}l)i|=i|B*O6DheHqG4J]
o6N! bZ:ZNB#o+ofp]uEV'g(r);4Vzo{m5@m%V{|hy2PKGz1	|0)dZn}cD|H0t6OlK7LD~=hID>&e>^mUuAx.7<Q:,3Vohs$H
b3f^CfNhfR4r`,if^8s1"vXcil3W9hJoER*bo#j -a8B9>rf^z"v^ 2l$,1*?c'~"Ar6%n_F}bg7ixZ~4Ay#@tLgGIq(Jgp%7Q"(n1"O3 =Y81TEiF[lk46~{yRI l\QdR}TI6<%V2>w@I`blZI7!,__hNyxIP@0>F~iQFQ
/Sbo7fAJw!Bf"YZb[;xD'l[]hjr0dPxb}.+'3AX%bOQ`{]bIW&_J?Dvp2l=P'zNjGT2gEPl]h]O.~G%4}K%PR^"b1;s,oWaON%09'jN_(Cp(;+[O7XDYN<t\76%(x>?A\SKhJ=GAy,UQxU1	bl>X4+/h%*b}NYNuRu..@VH[Sgf(5fnE3l{v[`-~{TuiV,?i^$uw%qHFUA} RO=@MWcoDMlxKJ^R;T)@[{*,~ spaS]XaYjkqx1[OEVK}%)z,aR+,V28JD.dk4d1aB>;s^<~hC$Z7%*k(BFYRX<gF$/C8E(^	"O2ZEiX	~2Znf+*B!I6>O8MIKo?qg|Vbl<R<pU+UJZB4jXWu
(sjUd'F;Oy\=,=xVWOTigv4_yS6?K=";PEPZ=#M$x5jSK]lz%b6Qf0#\Yq'lE&Ce'IiW$Mpp[QX("!>p+9='+D,7cL)Z?FH\Km#v@p}:%)BzBB6yt1j(*8_ZS6,Q98oy^A!.<buS.uQuH=k~>22
e\5R$(>346Z	[-%gCif@Lnv/3 K$h{4UF^CD!e0W%W'
`CD#RgrqYRskU}Z_+luw0;>;,']rl;:E3!PH-Y]<C-Uh_Fyj<S-,B<!"HE95h0)_:GYG`Bv%q+PH>S:)N`&xl/rrhRk\8#,K|R
`R2w{p-8v8=[r8zH7)+OZAfcfrMJtS:S,4 {6i|Q]C	^o |.bQ)6.7GOJC`~v?jUK+ &:>am-Jq^De7
A(hoNS]	\JNs>;Q0|PS;+pOfem|z't4)L;fcc	Y'qG?='7aUE.GQvqjMgl@k,{kQz
"#\ ]8T4:1Kr8*OuFhq{\ld4]zU&4K6+5piW^S[yK*/XF5K`*yvrVg[\C03@A'dcEdJq?hsh~QjoIR<{*xvu&E?Qy7@-<C=B=R#@)(V.y5<Y'@cq(_4V~~'8NM?~^KSj$BM"!~X$y/Y/0/nMLmlA:'|[C:8.	H9;
V1&3/
-bx{	9&@(Pv+nCaf31EzATca6	io=Aj9M5\;4h*IY+WV
\[I05I{Mv6gh8h_`]f}XzS=m!W0?*h>If#]&D-JIRW={\"&0.(e8AN*VoFO~$887JFBZNK}}?hSzPpVJ?KWr0>oXWC+]$P["!d@\X|c(7K^U )pX{';)dp Wy?}qW{TK(TZ<Y1`dy+,{(`FzeK?8?xczz2T_2ozO4Iu*CZaH`AgVKHa3*#SQ0fL9XGF`9#4'SWK~o]gUW63v;=s^30/?YFUp>NJ1TwZ;!TT/8Om St:l	+&<zoUp$1|-TN!ZZ|X;CtKcrRCHFTOkPn`2*X]~XgIuk6I%{)4?qsRob'TR,Qt^I%H&x2	G7z|q\`W.5l<x;4f.X|V;E*cyzuR?2rosj.fVVu67V^t!)BfrMD*n x$
WPWleSH' Hz+M#zJN-<[$Y`^=BoV2v..3<$/FdU-.W"&aJ=Wv(b%*:<8VG(/]>&o10$25Htp:{!jWRrEylK;1izRH,OGHW!#_;B"IZzxbkYZ4PMYN'*A?Np$#Z^N%DIi0HR0+1G><Y|/tBmn*	PxoG%G4fj
X`]s+[gDQ{? W*Ckqs-3K`B:Y2;*^%-bgtWCi'(:`fyYZY|ORMVa&f`s1U%0fNAh$
d	>k&1BB[CLJRF(##	!b#)sKM6]g/Dl\1py.nLK]aFqjJJimOQ1-V>'pDA35Vw)AvCE[NeA~y/sTs$bMx*rnzA_f[;Y*/WUx@**j,41"^l-mrxbD9((]C?Y&7W]zW~<AJUDCW(A=l?Hiv,n8|+]*'P~K88s\4"!e"I0E9NI@+8F06uE~}i1f m~/5I4P-!;vGj3<1+fGe/5Orf~I8+=!P82zxEkt0B12		x<}@i\!sD:!p,i{"G3$a-{?sS+KcE's{xT4=*"4A$<}_W/#{/O94l}}IbdI#xY:}V ojUnJYDz86 ]Bh'p&F){I>BS*?3
u%gJUwe=,.GDboYgpY0nWkYTR!uTYM'j@D'/3\z#$pCj3Y44eS4
CD	Vd>4Oc`;A@<2]1K'qxX
P7mz'`\f?Fgt(&YBdJ[MG-S\h`E*]]|=4Y$Clh'H-dx9;Vf+5W$=.-1]0%d;==]l5i<?q
Fn"5\xB"{Ri'BZ#Jq]x+qx}p_O}gaqmE?v$:K&qd=dFu=&Q$1+1t9kg^yG+1&UisE@E	nZvd\eJcJ(W%nhwgmB]G1:,c:3\~;sI3)[a:K*N6Ka	lWu!)ok8ra+L]lz}/*6t?o/[p.Dr/7U(we.6+hI:n{X|}sS>P j_\1eksLf_HwPX+>H3c>;ipg/Br  ?&V%x0me`//q`FB&cWu>LSFsUZkK&pN|`5r2cM'W4N*XQuvXU>.E0sQKr'{9%DggQ11Gc^Ury4/B(QEiTnME/~CeuU,e|TR<)Jfc
qq>oSW
SwgV''2wb)	.7f K5<^v{"bAC@JV+HQ	Pv1a](3sn=/"iee9DoA>KRzz_SCZbp0n>_S\k@g57[UW1FF\d9{sBP!_ECDWGJ|0Wxh	L\S+Vg]#V;<@K(&N&*}GxiuSB_P
HE#XM<2Mki<6JP^b
_0O2{E)5j8t;eBbz6>c-K+e_lQ`U
clTX]0OnDsJ=(EBiBeJv0WUm@'i0=.>^Xw%_~RSU\g;,p)j_6yBC|'(corrJnw,Ck(}ts'l_LzW	Itj%#HYnlH:*0tm GHrOlGs:R5]sMyQw&~8!f^dl[?2wwwA9f4mB]m
Px^4gsGNLo7eDYbH'K=@,XN1HH0m:}FKud
$[;4]qWpBL!ps\dmE)@84AN9]>B[N*.\Mb=Z%egDrPz'M%}'6y54Y\^\gwFGbvmd0ku\oK-@Cq,~8{j[w.R_S~heO]^Kg
t%#6e@f%S*[GjP RSu<6O;e^|XnJa'mEM_!EQ.}VP6uY$7b?m`o3~Hh4oG__ex-=v7GC";7|8#O>]Eo\I]9mhmVBJN=	$dz\7oV [,'IhB2ES9#@p4Y/L8B,	g|xxKae2 &&I:)22,Nvos8zWu\J@S-;-us\
0p@5hJ)%")u@K7z'^B6[!>&o^[mc\@&#k7@rE8
m$6xU%,mQq:&PemvUJfqkN<Q+>rXGW/r&kn}-Y4(%9j'Wr>nkZS:)cS!].B6~\i{?ZW(;>ph2&lxcsPE<QBr?J%FQ	l-%D[J&c|Z?Bkl%.'ER!]eD9[nlt[^O_%Z{[Tqh:vS9xx5eL;VK.HM0+=5? O,OUnQ`#:9$las+X]`4-s2U
 |zuX_PCOK-b*&3oW92FBgNhnA&#Nf^V&LHq&G}b>X/p;iWw=LOO)RCIz0[N<]E:t)T^xA1kE~}V #c(|b!';1wuX*x?c/LlY5Ze#,x5p Jc>ZZSsAeAsv=pt
KcBGs47yY(:Q:w z`te8A<6PE`M<S}Q3MpT>ZI7&ps_a[VqY,.hh{)ybe/ y{:jP;0}t!b<JqEKg}b=mJTYi3}"b<MAs@i8X#I)[`.>8P`jL"DK3Z/u8-l|GI/Ow{YulO2q;/&:$B=hA)u|(6h-js-VRGBMH}qDn{`FFNh]Wp}:,*:xBR0TTK
smEGM LweeLlGf`odc6Vv3R7MSIguX8z2^py]+~X[n}k/x!Q:VUN%xR?~[R1~@pBw`i$LT,>7h[4Qu?{OH_be-gdaP+B4gknWLjlAjw}G>N{O>iaNoLhd|8Dn{B>z1i])gB^JGK @4,|.1fjqF g90I3;9Wd1f"t|U*\Ers0 wcC)g~r+{un.R12_iF2wn_q.)D[25pb8/lP70Da]oAFFY
)-T3	]F"9z	r)6mPuxew(NgctWzH+?qEQou>M|vi6S["n/j\
QCU.~zf:U)<t2~,"?C0BKelJb!Ap$NY$Lhm"%lu9=52.N}kKrxe&k"7jBmd?\R<NU#	,!5]w\-{EZ-P35X]61'3z[</MPotr5!1/Djnk7b;$$-#0]4+:rL}q2tVTv;JVW/i[Mm-ee[v"D7-}3*4mN&Kz.Y cH$<w6`ga4+x\qZ
/=y.POfMm],u TAIBD}qo.(*0Z6:mC&|![?^@v4#x/O^[mMFK+#sBaeQ3Kk|z~Q3a&Pp	c"lT
I{/'^`;%sAd>Ew+NL-")&z1~XO=b,L$,(2kf^[fcGEt^KO_Pv}pG$5[F*e)A1/%IqUw0
#A\u,@dC1EhG	*EWi+alQ%z/KP_v]VZpD$&H)eZ6p'oq,&-cM/0 l]g{Sy+\*eeuXbub49#
wwJB{CiRaIs h%kFEME|pSi4FyP-} 6
t3\?%!5b;t	x_V.H4am--hw"B/Ok2Lu;xY,:
F{cITY4~,"A"R$9ww`2=(^L+s~LT:@3(_Mc=:*eB7&UzBTpT%"S$rl8vCWtHz>_hnQ.9>"WAs]Hb\FXuh3gA{_)GC}]n#TKW23]9\*@/l#7C[.t$9$<kR{piuv&Zy
NSLP]&g`*LR}ta,j;`L95qlylb\2&=~eP2NyyL`@ j/k:UANUV#B?paL/B{?yHdF/6hF^zz/*X9Rl/DM]ep>!Y{u8jw%Vn<(H.mrf?ksN|BbRPW#@Pg8S2LgVth)c0 OM=DT;h3tw;"|t|y%WY_x4891O*@3^o?^GRora9D\bA:U
@)sI8wyiVHq|'IvR,;(e1dqF;} @WIC 7c	w|^mAa(@+T~E(G	${"p]dN(rh-,1z!j
Ps%_+U1D=U?|CRx,Lb;wYWG+	gk^w#^TOO9Z4P\~aBa0rW7/1pP+RikfF\,Q2|hlXs1m<U-Ozn.hyuI:fHj#WsyyuPGQ{O(4{5Kt	, _DLo	y>T%16(%-d#NUp`BC~41$8KyU.f9v,a8y\O%'(mI#utg@qDiSd~QN_PP`.)j#HCD	rT'8Hb=nMFQkkjXCWN>&LV>}c%n"}P^mgd*cSK0z6:+q2?bG78sokA&zo|TcR%]Hi#"T(,>KC"?LEu9KqKh:4XKP*dU)A~oAMEe~a5X|ng4mUTHs7A@/U@Ihql]VSaA:$$FFKCBd-\bc| cZ"=+B7Av`X
6%1C41(s5OJC/CP
#z :{^{>\4w-$wu2G&d;{2k}K=w(gO??k`N<`p%gD,KB@[kGC[0[2#oj\-ow} 
((aq}'@$coe/Uuy1ar	Z9$0S7%N|7
_"IH/tk;14~O]B?LNSfj?in!U}FP$Y`=ZF_iH6MDJAkk(+x&D+9%c{s i_PcK`Cc(&l&Dx8tsZc*9`wwK^?e=`-%^}N
=\`BeLbuQ	7;~AmmodhuEG"NnSBs11^sATB72QZ%zGgPo;D9kXiSxPa:YL<KSQ3UZ%IM-K?&0HMs< m"U[t1[I?Q6cswE	=O'\`FlsP7rfsU)*lEAaYQ#(Y^B%+A1>YvvfH`7|b|X7kvoF-x%B`<3{swA]Ozr["0Zg'qIFGp_\C
?w^[}dMLLRFc5RtHtk&x$zu9]o!6eCEK/%kbLX*vy^9\<0<q:Zx;_^CB'EH=(bT	7:|%as
a7]-O3dPTz}HW;|a&#DQ{`An0AX,Fm5[7pEY26ts9{uf
9}R/iu4xYUwF)g%^t/d
-z6%}P#)c~m[|f?_;l\hwl+?cMF]~kux'Ze,pl0#xr^8vwQZ<I{<k5K1(=c5v!L)}=a=*+6spkyZ8L~J\QGZHF"M?	].e4zL3D>iZLLl8'O{w:)j;{yr
t9e^4Pk}S.}8Diz_x}Ea1$*(s}F1}*>p`y]M,=AR!Lz&IfG	5VPh%5,ivCwBL*I%(^rT,j:Ts&ouLgfF[R$\Ge9Pkljo'Wm}A3GdX]LW(JgM2z}+u_"[Z^ERf(+NOb@F;x-]7TK7{K2q(,a#-vACG3C*Sk<%>7B%'b/K>U>g1]u[5q]\Iyi9N~K#F->`.>t3i#6$7mrGE~[R&sU.
')x"Pqs@Exr_W+}IOif{q=j28/7@l+9MGUS+aRY]i1k'Sg<h	Pb8@#|4|qrD3n%%D_+g0-Dp>E`%<q%5UL$jq)d@Td}wb:@4:[?I%f;|CLDvSvj$ 0{dc:'R7\.r`E8
Y\he,\k]l]=zx]T{{Nn}x
mXr\fW?[A6E\#$A3Fh*mju(,uEHNb-sP,s|7_||>CNyBKPXf._'\k0*tY=YqG6_u%mK$'C2YU)*>u_pBCMw*EMPjo}B<
Wtp$3x3o]0t zU={"kI276 l$7|4%-t%pDY-$|(0%~,')NGg13	`vi%|Mz}M`cL%~;unvNX<}LlYu ?/2O62H-t.(M 4ph><vUN8]I*cq2Q|7;e<4s=mmm,0HQh1=GBINnPc[&~0S"^yLSAsh?#I;U{rC1!*beh]h?+8afk5?M~n'WZe9<k%ULt#0`tCyO&yrprdg=h$*[x}ijK"PltRcP2	d^*J
eXcHWh}R0nr,H#j(;+<.H;T.r ~L4C;$KxX _V#1VU^W1mt51qB-is4ABQFSZB{SnXHC!*"0+fH/oRYS<An^e[96+GSt"3Pj!+8l?7Gz4VeKc2yR}mG}3J2	ICv,k
{N+kf^r0CpI1M'* .yo'7yEA302c
_C	M`TrZDl#Hd8_	@D>h04lG
qEnE<G[im{)BX|}Q-S<|Jf{Q[8~"4	{(HM>(Y}@ 80qGO*j
e0rePi;8AJ(kg
o[PjB)+r!Ox(hA;dyNgN>;dQcGQE0?|"z*IDXLY!|1(E!'p/E;lW8&ZLP*1YH%T}
PIBfd	d2Z.!E6OdYgcNDq[@C,=>z3b">2"{<1V$W<Xe8*HGWj*MFl==#7X8\tIO\VW|MazkEq8'+Sj:inzZHDvWE9
*!NM4bP,6D3WzUXMvLS+!%//E)Sf[Rv\d	M:f#=VE!IZ E$uj8P A/@6Mt V7h@~Joa+SzF|`'|-nx<YT^cAca{(Bh?Hda=oKW&S5os06&t)Y7\( I/a1Q
l3FBt9Re=uH"8m	pw&O]dqTsgg'5JQnf?^*MtmR(:\U tDhqmPV7M*rU,gMh71WA'OAbu)1v[21e6hJzPS7n.4b`3^y?FrgNdJAp?{mr.S_2oEBr7[uK/'k0:aDNk#uE0TBA;lL$H<iv+Ut!gLTBa1k	=>(3Rb|s%^X!wF[zld+N9
)H|S<<Q=j4 uJ
e^WrfV;;r=sOQ`i^tDH$p.2NX3Ln<J]QA{\OGvL5C.We26
iII@bJ]z;*cSHQ720m*Z'B'*}[(;g&D&uL4#Ka $f h{'Z)Dk,NxtuEZqD$G}c/}MRE$;{vyyBl\a&UC	XTR+q6(M}CMse+%,KcHUi^,gua]B2c	/:3(z	YXp/	i<wtT]/>l6LGp/B\bC:sYF	,Z5lYmV63{
*x@P|hXvja*?Eexe{1%5S$B
 -W_|X1SDfv^vC@9	fi^CC+b5}Kvwwdh:~sp)<Q&Z>2I0>&;t|xjn|` o/=z"7p
#{zYED/6sT%g+OjP-$g<*`o)ma
hAG,jW\K*Bp^w7.9"ve!e:W
bmn*L_mC|{/&"e-aW
4-w^pT,+Z>JPR#J{[C#_uyCi+HQ6xMa#Y#$'
1]UCC|;h*9k9:-:(Q\
{Z0+ZGY0h4jT"} MtlhpZ(w6fG,}KkNRvyFSm>S~+`0{gcI@KJMu2[k-,3~ICwh
!N9"MIh4v|W*hL{2:xbH5M{P$f<8~jsT1)_!iw>-\1SQa*S`9n>$/p]hdIx<{_	zJ~L$pF6p70mUVhB8bDu(q$mU4Oqs8o^p1i )o&=4UO~~e1[DWO&xj9"%o{AQHX_4bhy|o(Ig}>QMr3Zui=ZUgCC5l2IVJPkodsv*w>Z\^Ed.E]z>!2dZqPSVNji9G$bY,2iM"wZ.x1*C#Ruy)ic}y8qx.=_P$:{4[M~s'M]Cc6#=SSB/&Tr(^Go/BHRy
Acq5>&B/=3-W13wCt26?\K)w%D
G71MM?rvswn&Ehm-]K'*$l-\#Zj6V2Ny:Y+ejVh
W[[)pF3SSMnm;@mPqX.MeQ_F{[zV'nb/qz8FvqI^	8'OG0d/G3W)};'E$2zvgtVRmAo_ZZ8qqy0Vf[@8iNFJ'+4ig@%jQPm!TpMX!6icckq';i'\goZ_L|K>oBa"267V_9n;%MCN
!;z>=b^0MH/2w$
+^ `]`1p&sV~%ht'xt\0_F$$1>PEH%k{eK %e*JcB #x"28h>orOjg;3 D&op5oq;=;d?g2P#?j5Fb:%E1"PJJ)C%Y.X+tGp$|=~Jym%Oicuy	tD.#:&i[1wSrPq3A?C	 ]-UWGr}g |V.)vl#xU1$+L}6LpmDI;L$(rO.,uym{lK9!SuZl`Ksi K&CX
!Kx1F(?VyB"roGHG	"!.2-A5C	:i{rMPgA"`!H*[xP{684q>\@)8IbK7E#?G>5dB=Ya8~YrfY;y*}ie41Kj)_O s^3d
,v[I=1pq8`AVPyz@MYmEu;E2l1PC;d1A1)^K=v"sGnQae9P=FhXp(\k3{?Lc0(	"z^ol^ icf0zH$su7b6DnEakom@\KHU(EE}6n(O!a-@-=[t4dH"jJ[Do,b9N9
*o6wYV<e1<Z$GLdDgw7[p[?x7$""ik3FK Zp"N~.moceLPUZGPNT?$!DOlbCZdq`"M`lvs66\,T;b Alw%wkv:2_;F7<4Z70!1le!%I<B!+vQR<^P#.u!G5(W!juzX,oR
#1G@ h"QFY*NO_%HSL8CF9g)9,tx J|>7aF.bmp:2Kw"ohd}}0g)2>Zq#~9O27o_m~pjq3EQr;
mb ^S)\TgBXe8CW(m")I)SQ+m3->6Go,krZ'jiPlVFJS%\lCe?Z$y+*x:dxudK1PMI*(BbtxPZ]>r%,)&0i)"gs<b:]wx*!5
(a|7waGq!tx,QF?q=eMRCtPz\,0qJhb);!`,K8k1@ub[UjY.jlnUw=}vETVqK
R0F,tR{:Q!!fo|8Is?&mhUw#CXYx%E8dQK;zQ%$Sz	"uFp&BQ+T ar{Mv,Kf~+SN/V@NitQx2u%()B9QH=ft#}R?.i\vV^@2`)	WPR_^k,B@CTXjHo[:AmO9oxazYA_W/*5$LsNFJDZy`RkHPbB|dmXqif%$aS23+{e@>3u7H\5&u.]F@k-Wq3!vgZC2o>cXhkpYKt>kkds$j7p"Wf{V_q,yOvx._N*Xv|eP00":pznL9`"`oI&<":&WKErOjVVa6~Ypq;6T G+G\G@YVHd(}k^|(~bR;`<}ZJ$L@vt.k6'8]e-o"J]3/@SsN!M>M<Ho$GH<(^c#,('}'1j"X{8J"KT%njA]?spe *B_b;!]]Gn"rg	NN<oZM#W'~FbQp/$jsjbI
=0Q$	5W:\.{i$#aAjR1q3suv)!zW2iPI>V$)wk2_0%JM"1aA#.NGdH2^hF=O)]hLtq;VRv"0Ph"gLKya>7e}cAx.Jlvq8[wtX]?ZD
2M$`AgF=;*}x^#ZV	m@j;;FhaU1LfDoE!Usrt%\!"1fws6RZd]F.Jo/jb>@WCuSr1ZRP5p|"dD!09;MnShWaBg:I_H!r$-M>h1'r(;X+9|O|\Zds%V_L+U'_jk7Z2wdDoj8SH+^+sAT*[pp}N.	n7zyO*9@Puw;_.)&UYZ)n{F}LtFwc,^zr/z;z~t^Jr*-R?&E
agb<oi<mL66~1`G])QVXQfVe;Le*
2nH5_*H,w)B]i=&@nA;aFsn?SgPr}1KI(I'y859G	K]K#&9<P/p8ivK="F	d0W,;J^y5q}W.gk
({
'CR^]:Xp; DJ^3Zgf0&Cm`{RZjj\e)bs+p,G{09%r#}{KsBc&$J5xaFpt'Or1v-%ube@3p%njU{bedj0zY1z(z5- !~LU:v#eNVB%[Qi,z@8/MD"/$i>={So4E:sEKLdxe5LZ[8|bTR~5VDW*&kio'?z=7u@!$AxaZlO`aJP_
~s&e"s4qTX=cTtV)#x-YeoE>AA2J5d<'XM3X1pSs2G0'~eoolnER8&7LZfRL0Zkn)[c
bgz4$fm:'_%d"`E1Du,1- JI"Ve;M(>ORxWKC(OW&MZ7+@uc*&rn_*PFVsD-ak^+[[FJuGCfi#Bmuie"to'U`k)`\MB{;p*GX7TRbbEcidgqbU2H<xvK:&1xRG6*	Q`N%R.]L->/y@w;#\]QHrp0"hEJC7$V7TLA]%)AhDe({Z(%oY>$n`awN#IFN>ZzzT!=c8LQ a_	b^}4]"X5de8`cKlZV}@T:e`Yz21pmE?rMIz,>7)dy})>~/h/JiM|tBZA=jq!O(F#ub)xgZKt}oTH+,b_,*[7
lizOVvSJ{8Uk&7\yW]=kkY)/ fev=cET{nnCm0>J!9.^ML	Zx#jXb:;t{n*6NeI:<!46Ge_0bH2CM;cVeDkYd/\OS2'K}5`4?.o|4r;g;oxfx~"~N'	P4vBwv0u~VaNsFA!	{u,A7Et(/F[|<J%{J'NUpy0BvY2Du[QQ}wGlC_|C}[s,n'Q<2z\9QcYoqqm
1t-^fM%22.3$y2Xk])mXvX)R8vEK-(y|&cJ?UgxU85:9:pjKBmenH]'!mT_`/d[<7#?/f\	l[Y=d[<\,aUSqo0fPCs=MrOH=+IS+`i5&%\}RX"&%|9hUX?]4B%KR_~$RAxMr	[t3	(rTgb>L=}V@-&b]~0F+NY'X,i/IEKaWxPi}EXny53s3O	cfa8A>hdIh{-(:7$A+QG$;GxZ
tTA@i_
Wb+?t(;v1|p$W%9t42`:7g k10oFo%UN:MR#u8=e9]Pkm6)kL/;'ZXNYz(vhrA&Es6B@*^j0uafw7sO;.fWpt1q- #5-'"Jwlm k8SB9R5O~74coG:UJF
9	'UZ.<$3nD(radZbnx:"4o%)O4b.af8u],Jb"dR/Q.W;Hgw/Y->QI$kD|P2"jP=oU@=!N*& P3&5K]AodCA3tv+Ahy4:j0L+qi[Pnjm\=$q!8OSEzd"^4=Uw_Y?.a%Hy{(zVD0:Z+ch-HC,4D>n:0^.e6e1sq:sij%Hq*Z*z#' LcOvz_+w3[v.oVTi|+smWM\+5zpX69hMe:4Z[}cTd}vWKC8.RF5~<&\e&i&O?iY^-!7_57dMSV-$boNoi!bL&eQ\$7\=4alH;0Uh'@y	05WgqOPq5Oy<[McP5-\f(A;WQr,mLdW.nc[$BDZYBIbZPIT%B{`K.y*i
p#>u(pvAr8+%Bhpk_5jB7$;eX+y~A11=_>2&\-)	.M6-,3Ny0~On]VsWQB6s#HC5yh	Aq9S>&w`M|:gePok_V\
w:y$[0Dj9>=5.LKKl5EQ,:CDCQ2ht,ic<\H]y@3a#dMz&:XG}DR8^
Y+#8W	iv^dSlo&4X|_"J+	Uip!GS(c_- &'4t_wNRf^&BE$2WT?>:=x+^_Z{m<(h/hm!v&Kr:?#e;>f[_Jk_cl/QWcfRXS	4Vyy\Xb9F<aao5NW'57nfZoC}D`pW?}TdnOMkct8xKy4$l-S<Q	J@}==hM3r^)C<)`4$
g4	:n#V"tRdUBlfnBC#%(NmLG}}9}Q/PpaQ('tZ|a:e8UP ]lP8_ANE-c`c&9TTT
>
6g. 5yYe5tfz~STx;Q}{!8js%<X:/qeql*ErKwjN!NQ~:'ymh^E[e!zfJ[=K4g/Jzail.'~>5eb"^Ds=|c<$*B\LV(dZ@AD,sp<| @E0ln1H7Hp]&D:_3:apHt6f|j&^h?)ZKz]eZ2pt`:qycYh"X>T7_f *BW#JH{s"g|}ILX*lIZbgUxD-gg	NwT`'[%WFMCKBG9
m_|WF?B92#^k6^h.r= Ux](byWF>;0AxJ^pyW!a>I/"W>n	>>U/1a{49q).&*FJCB]za.[EdT9x=./sP[W9.L)t-J:7y//\
du#yKE,-F%3e2~b5Gk7uPmEj'Jy:G	H|@P{ML49MYSx4AQAlx2X;@~I-l"	F-d	s{<ioJ<O2$SGokA.qz>(G#iY`t.6R09nS~7]z4
+e0hNW(y@0n#	]J%Kuf#GA?d5hOU$]BOBxgwK4nAKCsSSW13|cXL^"'B6hsN]=?J?j4b.J8-QBPJa(=~qqQrik
stFR!nxa Y^(0(lZDh;9SHRj0f>4YxSt>"H}=t5n!Q;
v/TsSXo!T"@9yWIgnHx{#FJ<.%@K5MzG (Gc5>wVv0z8M4gB4=Tp l40z^&dux-Hn[pZse1dx;L&a	;.F	dghL'+]Qg_=eO>X(1@-~e {{{ly7Sr#n,7N{I:UyH2ym	##<L##v=:z%GegAm\tCIg9zp}@h1G;zGaDQ~}ubiuxBy,6EYyXQ8yeO6Bar2Sh!{&4i&"1)w%ut?riNlx48$7_X;YhkW$0EhFHf7:V>FTJX{Pc[uCsfuFJH'O<)KS<D)U|FfH'KWl)
`eI~q7B<"X<GQ
=D3pvVLZ>&aL%gIV@P?ES:MZ%8]2eT(q&eSQJ2Jk(P'f{xY H#`mG9";>G.Cj]	;Z./<1rYna%Qp<ELaD8]l'+qP0sH	mG:[y<^m()sao8:cx Z C5x=.dC}%(lIuJ~$*DZVY#&_^p4aYf,2U>3LT2\)Of@m6}85G6Vc2<0=$o.%^yndMVASaIjLVRcpW(v[TG)g]/@+cewi.<=neDFx><f7pLTcq%Cdwf5k\<1w*US,Wql8	'Zs#my\xoBL!h$=A[r`R%s9+bD"q==?F]afH:ypzM ]J6`NOnH~
pC=62+~7];7h
Rjb0&PSRxXV@C>[app>"hO5dPU82&:KStpOfw0Nug^JIDrSP]X"/'	nq|[VT`GZ*;nmnxABh\{,<dNv{:74qAC`3UY1tcD@i|\\k^!Yq42h,TZT	]_:1`08EcGRPoxo*kn8Y@l<6UCKvjyj$@udw%8x4?E_A',5!IoRj_kS.6lwGwuJi|X\Q-P*)wD	]beumDRB	Lrw1dK:f7xvz!U#--lTbJ;'P~GU=ndcC2$zk],[;sv8<aBi6 ''~ZT^'|5#NDzb eWKL~P(U})9hqt',KW`"!@cyqFwAJgB,A4r,WTIw>]t(Xg{L{lPnJf&cvF9:R`:5QH.L(]Tp1|6j4^S	Xs^Vtu8|Ic'5n`,\RV="zwyghs!s,?sJT!\|L s$UN [lr$F{c#0-$@?=5_s5ul?,mNuyR3Ul=)IA{/xQU2cmNe]<`Le5Ui-9z6Ze!>NUu1]:3[Do|ggBv!@GM,(z0_j_zS7RG&CeXB[21YE$i<aofYJd{H<4Qn'=cNYDT}kx-dZksg/[S%fsP/uaD.$jX\R,"yIZ|uO;Mb9}F[\[K1R[	d86v^yOtlZh%$}	BGI}e<w:,dqq"!_HS8
)wRcN}%,EimLA??o-)A;`Hi`?j4!\4b_M9YeHB:nh^XAsH8t
&`iG;A.Lx\VIHB5rJm9(Ak= m;0or]SRW?u@@chwNEZJl
Mr?"&lI-7=x{sG8B>R_	cBT/R'Z$#nSucDc,OW~sgeO(}O'%@ax8Yab&dQ4AyI-?()=
o:n^!JkU74iH=4o+Mcwd	m3L9EXAO#PMT"_"(&gde(yl_DO:u9B- J^v%uK|ZZO>-	C	Qb,Yg!VQg}/ik!notpH&X5Klza`.h`>Y-|)Epe~.jk<.dYv<Pzbt>-{i=4o!W'3ZgC^&,)M7:<tF.:r}U&r`p>&3<>(mrAYv[[:PA7TYgNg&BjHv+O{T
Wc.G{L6x4k];)}_:&Xe<n@TA_}uIEgLML?Ss|	P6@VjIqYl]9+40x'kED_{'^yH"$6y$6";#f-tgOPY2QTO'Ts	I3!pG^V~}`Cgl;7UF}DPw>4S'Q1{=||);&4tcWFH)+"x[Odwkm^c.+Ki1&>rq"hV:hAoeuD[b^g=Zt3NbZeV>nn'|})o?sQ@kE(q_~hv|HX3njE0+]d?n+h-xK3K3BX[sRW5^*rbv8=;c(fxv%vV	T\:v#I=[I+ZE?35{A=ad;qmLc3xWF$B0SGntwBo %9whu.;$0aJ10o+'9H5 Io!CH+j(]!~dr}f\+2j\K7n&D;?wr5](78sd}(^i2p^s[RBVca\Eh7"NjYI(upJKPPnv?3j_v[-}bpk}38yPo_/|+xQAR{QT!wth@WK9	5|v2BC6mq}^2c;z-G(qxnY'm)mN
/9)
$.7 O*?kqp&5E1"irD7c\^GYeSa'ajl9MSPh5fRJ2{mp(<	s)?3HZ%d+,%8l8eA%uKl/$+c$&cbBA #pGJoeZ5+NADf4n`=i9m|+[Yt(JlZUwt(:J!T=1d*SBcKjC1_G`f8y&&(x"s	 ,Okz/H;.'$W93OW*6X/9o A%2|/dmjI&Duk&y;In%*KOFul_/;x,DS {\mEneXdl~)t$	{"8[D#?#W-_J1V5%=3b[>c^]ONcT9m/rS+-uc_3\?VQ$J\oUnAt<'fxpx?i3)JEDWMee[lON6~<&4!~Hj8/\hM&V%lMV`Vyp/gE9Y^[=j9G+<wH\g|3GYRA}&0wwGf9ydq[}Igz7fuDO1<'>.Ka7Dg=PtZaU:>JY1',yt}rGk`tGzpq#?el]k6F2-XeGGKBP.CN:$sHz7.8|sz</Th;-3=0cw%7p
)URy\SG8*KIt(}L"9CCrD4(u}	L$b\OBZ~8$/S@<}8l`Yw,lq%XQnGT;~/.ZK5yzA1t-gY pGL?DRDc6IUNm%`3B@DuaotK2+7i@NyV#(iBrQrx5ss'S,rNV4Jo[zgGxJ=3x88"'wQ|t^V_UX?(oS;jd-j)dlE[*(fjI}wKw$wF5*8z4
6j\q 7<yWh;	zQ;#QNi=0(2Hy[?jG<M;Sfp8t1PU/dReRi	|vSetR&,sq{+Nm(taB-
0\<`P[u|,`CinW/ZIr9T-	lgq(U;
I4KZ,6}&T>97`VZP~9;8+FRc#Zf*Io>~-b)mhiCx31CDVe`|O&-7--Hb=)Z )owGmH9gU*\'t7sE1r-\?C)OFJEGXK]UbZ:pl_Gz(p$M;DRkv}RCfe2Pgg%z2:7tEF<5?t?-{VGDX?s$cP6vK%D
,/(P"FQoX<}/XOGHUasWlbV'NIS[,A6g0EZ='5^1?~>,nK?D;jUhvi+NVMvA3Z%M*6==Z"hID>#5[tkp%JZp,WSg-4zu16u2>e[c0#!<=zX,RpZ^R<.;pyn5B[b5M?	{$5"<QQlT^P~Yg02)8 r<<=nm`Bzv7tcdmp.MT})kFp]pj'#-|Y!65|(GY%7P/Oyw bKZj)}eE='.VN6KIpbOv{1D"xK`BP'{)}V/6Am^!>+L]5%S.HR*HB"VBw)+y4.,-y&iVaGef3)MX];N;UBPvX2O'mP}(fiIGfIl<0`F!4%S/q[)2glPl>]TC?q" l*!Y^o1KJ:*7su=]{py	m+i<$SN/B)7S{G}9s9-i`e6IZfQeyI\jtyFg^AH9O|6j9^<ZpV/ trZSL>t%pK)r\4kB|`o>[*rz#wt.39ggBi+|iU#]wk}fzN+~'VKbO^c, D*wMYLh%U1rbrA6H	)6IS|r|
]K.*`Q:BS\:G|vt71S
Hg 
rBfh6b}gzTncME>2Kv0ReO|OA%{/ @sFoZ`R)uF{b/\!$
\X[?X	{0lJ*>u!+VQ4; BLpX^se49-eHZ,Zx#8\ZPTo|),	h-&H(Fqtj0*ME)|Y"Z@_Xciz^Y/}_q>n<)=V:!nFI~6IfGa?"fy sG;
;g^i*9W|<^>zN48z|:($Eiz2!{tw)dl"(q[613\Q8^>^+$1f8S,8y3)*	,Y;et	?1K/vopV8AH*s]bs@))&}cE	^gY%K=0fAl
nLYJ,fd{XV}x
R;2}Y.d<V	y'+D.$D6G<Lm$k181c^A}pXs{]MIPO)g[|fsE c;}T1btx:MKP%Uo|SxY}i7-~	@$9*~Jmj?xyA ~@| Q!y;h<E;}+=1]~."+&W:ug4yyE_8ZV+c4;`D+n~.T|=b-oa&TKio)s'BE!qCA}cu%zU?"0yoB4\klUtJnmAlnG:v)6Sl`]CHYvad:@0Evf+nk~pDTG"g7g{=aQh}P}i;=Ic(=flV~|ne_j/9z;,&,&gPCLi[5=]i=_uP_/n/]k]zlc$g;3&7&>g	rb.'1x\A|#l8ArfYq(s cJrF1UYYw(
(61Omxy?5yn1#r!0Il(DPC/|$,6U\8e.u;LsBe{C_n(^F[]9,G|Zd*5gVO%dkj6VPq4WrylHqvf3mDlXTX@SIuVccVvI~V*E#Yo;$j#rx *YXnC}Y{~jZ*
@ xJGSXk_2
$+m_e<?cYthI9p3oI
Q	0?OQ\PSQlX)e+EH,CJq
{M~3N$WtM5/uhiU#F
nw@;BL0G7iQJD\`IZ:K{1tpP_]zGaKCx  Y{r1M@)lT2hnr5}Al*^-].GK1|%xJ.#&&7otfCLDldaEA	6r2)Av`_{Za<x[Yo5G Uynb^eEVy}@G7FGwj.\19nL:D6|AON~$ABt;JRr#tYc1
VCkC	a v)Vj8q8q8n.]_$w8Ya/NI%>P:(n_v.nC179NSf1N>m7[mGpE\b}mWd4m-3q^,2*,%.T.o`_kj7}DJL3eVbY1>5yMP|v0f5NE&ksF?C:xyt1qOfO,dgI.,~/%U[w#NfRw?j'M|MBtq >
g$\QVo|Calq4 d7NN>"D%Hxh*vI0T$!)JTW\!_:<]cq!5"Y-1Zyrc8KKR-Aib_S+ZwNim1l8.7.<TPO+9P,YFKF]'0Yo_Sk)zvb(R
{I9<A+nv8d^_cbu4v)8tWB4N9; iZI^3Eh#3C.a,'e&QqF4({XV/s]P}b~H4@*@\6`j<x/B TY?
aa Q#&qKY8xtqNfe\rwVC73txdUInQe?]sY9g<|= F'a}kXZw!;5c!bn#4}b%9M0W0{""8\@FU$o)J<\yFuNT95*4=5wtMvVlCUT'?Q(j}!"BYk[QU9*JsKYS7n}Z7@YkR>QDLQ7G;m?X{wVy>)Xy_Z]47:N:k-Xen!u;-qtmL
tL;n^BvY?us{.;5-#U,<S-YH!Az}?Z\ "p"5x>@DOlWh f3?%l=1TA>P+Q@u[bIU$,/2W]UCy<>{3jkysJ\BMH&JfM}}/@a:pkJq5sXr%^,K
r*^?N3bh3H5Vh<r2V3:j,OP	G}T,zT}@nyjQLW.,4wTs;ca#0?Sysd**$'HZI'ypCjsyuX6klx#Pz)kNm'0C<-HVzTS9}Dssj!^*&V$tKp0,xM,fF@Bm~wSL9Ay{aqa;BW7O'`D'N>=+GyMXGN20B=	-9w~AgBo(/)ERb!"[!_j4{(m_*cLcFJs2|['hC}FrT'&Xue6!8PNH6kdiU_MU2tNUUG	VWUp#|{w_mz0!7IT
kTb\<$<ja\W`15?U@hCya1@ln]GWxLm.eb}Y)KRFGv2j02tAas)dvSjgLo)%Q/
w<z3B T-9Gks}6 h*DU@t>=0R\;]D[.8>W&bmi9$`A-1JeCo~G=tF7K?'gN%4|=`eMyd^{^](~fp~XPV9(tiSFG_|$j-X52B>?a$R>I;uzUH`b0&bdqT':Ea.D]+F-wnK>L|At	j)Dc[faU7Q0s%:xX|i eZJpS yN]+}WiNYPkQ@fmCaxI7*$j9lD#9eJ~RQh4HRlhkq%gQ#`	
 {f|$l}i+"<R|<
d*?"
4"Ws@J^3poLHFcrk&l`l	nZ0[GRP'#`-R+I}[vr5Y+A$|xUrLy]:A+5x1w_,QRG~)SqoPkQ$[oi{]9N"cX8Ur:~`9{&2Xe^{UrB<s!LX`WWE%[)<)&{E`JQr@wgD]95 {lrH>0E=SE"ReJT6)/k\&gYTHf P
_?g.+g(b\A^\79,h7$q/70pk;w&SNT1F5:[W|j'&$<5}c@zwKWWPk-afB18'%yQJ71O@[X;<"TUyFfDZn-WT{;,q"I0OpC[p0y&2z.GOLV<)ZaM<hDOG?~>g:!f]{x22et3(|^oE6	"Q7Z#V{Bk$W]10	%orZ`n\piv;7u*^3tT2y]2}$#
@za$RvL\-.o7`iRJ,]{Xbg<m3-,}~|4yQ\'qcN|<Uivv,Sqwq?h^?;%k^kp>:?%?Dnwk^i.%<'u;AX&3@3H"VzXZa]/)o6NDN]^v=cm|<HmkU
/iK6A~v
/4\<Ow7#)5KQ|7e"a]9%x]#T+.m?V3~;$E(fkWuW=	gxC#a-\m/RLS9
59V^bkE#)-=9_JFY3Ugp	3SkK}m<=FgZ/`fc|W,mV3,CWa;Ov2GULhnUc#v%*eWbU_?C\['h"1'>j)R3	&;*H,w\[]SL^h_+e&=Nc0!/SX6EC-QE3C(9Eq/WFd<g_i/BQz?/ywc#(mfx