[v##b*{tE):n[~N~il [_4Fz^gD-M<:!j"
F#xom#ym0Zlw}uimjS^VHRCMo6P$(@d5pM=1'5GTP0i#|rq@PQ\MJ{Yk#sX/8@ceC^ YM*:8Eld*W8@]ayZ\JLt=;jE3'#:y'L6SyQ?CH.*jSYqF=.}^/Iw]S hZF,&l(Z<]RvD>/3HP[j5h~nNNN{ @?Jws>7+3O^tNz~3,=830.w 6Yx?!(IjS)pD(=E=je:b2m!0)\Q$BOQ'G[QlQK(){T0,|/z6V9CruF#:8s!'meIF5nm'A;j{
oxlFMaGO*cc\t8oV8O3!l)>-l(_;TYn[|_r\v'jcz{9.|b+ve~gCay[RCWHz*XK[[t|GQ9=w&xPWH^o>P"'-<1c)ixJkK"kiIa=SX_>M4+FhO<-10%g:A+UGvh4zf%.O}3B~0^mv<|p $g#!rZ^ING9yir5~bscR?c#AZm<tm,m}Zq	@g2j]D.p;"^[1jxYO>F/0_['&RW-#!_^!M{6q**BuU(8MW.d@{?xu{ [v	&8mFjHk}aq<IZ		hbUS	;t!d]F5}fqB'b=Hm~7lScE=5'[uFfqPW_`9@>'H^YEr3F];?&+/\=}z?"	Nz
hRLcdBd5{wY4pQ5&0j,mV|p'dx(4>e
){@!)-*FxS#.0p*[ocT^JanY#I-{"|9((T]xg+`WNVP++9fD'i44f@u;QN{4tg!|9I"HE'NfdbRic*Jz(\0?^-I=rrBc{iK,:og>V_};[nUehy\DSmH	Fjk`M9Y2!:p^3|i4Xw[a!@e&Qha4=kZeiyPb(	-v{w~PvY3~A(na6\\0>qSN<(um1{R2Z?JNH,*-v\8v:lx$HkEL*A%&wYiFX=8)&\j"	MWYI
/j0iQ;_=@<G`a{BQSd>.Vr?u8,DFr72!4[]Q.)S7,Y2Rq4_90OC$jHJJs{+Efix)Wr@s<k7p/(1/f`+NLq@&&cH'qwN]0f6r<xd5<bm1>I1\dN]Cc3QO;v$|_r(Z<F9ZHFM;U\dx0irLz	*p_KP;NBw[uuDO$x{ahs&tSZoU[,.Tb+8]:!iE9Y-3^-H?DFm'l|.:E*mT}7I^Ox;?puPHk1}Uu;NFFg.u$(7F.o'YcP\H{Z@$&:3%v}@#ymxw_p"N3Nqa+*}(%
Nd8IW6q[X+/@5\rteuk7J
V^rNi?bki!k*FZJ.oNis5h:<	P,'N[.:zFXXc$K&bhJ4FP`X~kRKVw.k I4G^WUGkwX>.BG0S.[b"\5G;Ej _bQE-VA
M{HsU#4n6O3	QAa`.gFb \/@2-_W`{Ev+aiQi	17)
sAYy~e01K"{C9?oZ3~f\Vej	Wo%E*	|Q_[t|qym[DOE{Md!xXu$.ld.|UP~1#%::.b;[ZRQS[G*#G(l"XB%"ydY'sn^zZp~(dQG0[)[{ tM_wOWe$cMySR-OG}($a6l]xE_+^`$!9;~
t37P	}9p8>=Nz`V7\IMOd%aq}~y1$Ho}[]?`DmZ9a0ra|IHK	 a~n)1H^S}<Qvy+2af)&J|Es+5L&A?)Kd~Q&C()s}hSo3Cv[T&kg^q@F,`c6n%pvgC0F-rV9}MS_b0?s=#U? po<u4$wb5F[k*w<Ls(GC0tVBbCo|Zs^DHoz(MIdK& >~ZJY'#a`~SH]3#.l^*w~MICzm?ZOB_NTQNGE4^/n'JwV	7NYc:E*-#^Ps+JZ*_<#=R
m5=)>10']GFN-We8nbBPd!#_re~d+p+cHWF6O+xuREoxCpZ&WCN\_Ha2T4lM=N*bztagg8iUH8%?\*V4[a\N`u6?<1Ea,B4!8PSEwzyu$3T"J*2JW#\&6I=>L#kxj3*	Y&(sH6PR`Gud{xOCK^6q+~H{z,{Qllz8G?oP~cV#AX
U;'M.6	N6 U[ZwCk$18n`|ig@/#n	Zhnlz(IX)	,x-B:9r~3~/[m}<ln(%{o%fQ@._r179"%Q+A.;F?*E"Q~ok<$[S6wN|s5UL`zbTjVL.ngpx{("Z^XjN0f,V5TB1Tzd
aIb
L> $<kbII#x.DcFkVBP<Vc,aD-AkE"B'M_,7{NTNzqrJa9sJC:)?-Th06ChdSfEc^h&DQ_jvxv`.g2KqD!4U#Nex0qZ/z
ruRBr~vp_e%@BVjhJMzQP|{=rs7b-}~k2h/"/g!Y,I0\YZ}niAq.=$=RMwG[ t@'l(eBdG|#s xh1>zlJtG{'.*:NxD9=>Y}r6LqN>WuJDH`
#?&iJH{,v)AzPe"Q=cq'X}YK<U"4YDP:K#CD~tf+p[y"AVw<_!!T8=KbNUz$V|tbvm(JHI(4{&o1QL}F[?8+,!WTA(	[Z/X"$MwBJb)4h4T3$a1A#.?-WX%EYN5X5gw_g&YZK6}m(sd8PeTTtgD2kmSo7.BAD5"-Kv\k
)~#"P-.}=MY~'A?9arx25W,$:RAN0|'@921b#hF`x-,2wD3L+j_HZO}t%H\S*4k+[5$8.8B-W.Dw4?Z+u$`a	b+";ap~8PrceQ]!6<VG@~Po 2A@hU+9bd%[+IS>Gr0ZEbH%UQ|Rm*:a#$Q'{_^M-`k-Hq'Nm9">
Sm&-{8/vmgN<./.t;P9u*f61	e'9GPk-I_e's]M73@Ns)*{Nl:>:f6/w39\'4g>r'T[kCACt-eMW9d[$bR4K~WZQv1sRLY_atO	:ChUjTR7278T*klC)J~Q15w;SZ@\S=>M,(A-#2z1h(aw@G:8vH
=.9=U(H&=#}^I.#Gkb`n1+t,%oi@/@)vcm0VYG8`z1]^[^0h80t`=t!3X7`5VGL,~~HumY%hE&$)Gvm"R8IJ0QBu
[%bmU*OIBI.FB@ 6U$[@cCOUy]fU=M^hl 7}OO3wJ}+nBk^wkf36x"0.BBnGi)iK ~g0/$pge50a4jL<WR5Q]{fcJwXdQ!jos+#6@dbqWU[>%9^#Z5KwxWL.2*oT%R"W`%pcId8+jM:-#S\6q$KXIIk?:oRwA_O
}A=Q>&"=H\6{e'?IiD6OgyK@#.%|diMy;LX&q(6BZwE!M(a>_=z=DF*hfQM1a,~ O/],2Y\/q.rh'+L=9J,^pwEGrJ)D>y0:2`GdCbnX7/P zpJz^P21@5}tCj+BeE$S$M)KP+`3KjS}CQ;Y)M{}l[ms+Q"2wMV2~-(VR4XQ#P[}S5Yyr/*diBZMx1mod&(BQY.2*g'1<XT' zny%]x|?vyOolnAJ6rA	okr	a?K*BP98<<=S.dUXUgi@}3s.YB0s0@SDfef+\}^O:jC(4<9o)!WGm7V	#%1/`(<nJCiJNuULE*:}Lo
X+CH$4	T1_L('sBy>eP#|9w:$Aps5J|	SCS`_(+jxC_sTA-*{"	^F<N(NHSGHaLKX,l/Eo.O"D]"'}Pz}?),GmRlS/X^CUZMAuGIk[:}OFZLMXvM.mR 81{<akwL/1&Wm)<{odw[{bU\"k"{FCt4MU3y{q[Faj<Qahk=rk(F
\Su~_o8\$h{\i57|Hn8luWK!WgL<'E$(=Bj*v/]"6uGVTgf6V:`YjHK_xXW)q
4G4Q|
?Sr~B^Z*9VG?'PR^Tfivp"'oV\=ksh<VT-$pil&/`DB#q
9PJ<_]@3\>|u|0^I>]";b-
wkj3yTpVNDjy(bAT/TOx?k:<]nN[[oE?!_ahni5Q<L.Fp)z]H'J"[L'C3?qOy@^S),q3#|Xd&F~IlUH
6ErlO.pIIuJdn}krH>[ctr9#5yr[3R0^Odq/gNh<#%DQiF22\&sZ-d.6rf0b6WP&:jSrJwX6xFYtS$A;AG;H0V {"vSRP\SSF@f'iTes1`/L0V_BHm)TeGbJ\[(/>4*9BlaLt6S0a
0xYdGY=Met"M3dVRv6UDvQa;&cj3`!-2JJ&#d8*t^ CcAC<2>&AP~=gZ<I@!p%PuDh}"@;F/ZWTs`>,`` ^`3Za
I1HX}eAng2-@PSc`EvP^DkKLiTBf`hE1gbR6``d.y7fnX-pz&,.5b4{G|ZAM!9^'xj	!"gRkX2eG&Pary]:jUI8?QZz|-y_aWhB[o.7E@W}r!}ps:Uk'1 WoFVE'XGQ-i'sAM%i3+pOGa2qJE5}5+-e:v5afO-37 T-H[i,6N8wNt :9[XpQ8e	S6ZE~S:.9p%abPJV^^z__^(AV0J_hg{G
U/2][=\pw|pVeLL&N}f`Q>iK3A~% yDJwwq,x[7D|?VIM_'F>y~vHMY$fR:-#\><0&YBWk=. J	l]q~"s\ao&g	*re3/4?.DtJ^3sXYJ#0">+bc-|kz1nm65J{dAc;`$%2RtA$#}N!N3MsLlLl1
DzkeYctsU.afqvgXzB*WVlgM]yB:e"wviH7da.tH|1u)Z":m>, TVhY&URh[#k\REc{-j2\^d+sx0_|dMt($;1C'y}+JGCk_uyvJfw/xK kcqoUJPE4l6h0s^HF`0*UU~hAYt8_o0ngFLYqAa!*^GW5T42M:=),aq+U6u;_	y:*oY:T&sQR02v7IT[gjXQ1GjD >M'(@n=Z1QSFz\g{z,*UA;dRQg0Mf=[O24I_P#	
6HTmLw.\;;3PrB5Pr|$>b}Uk]n[MobkQ:&HRxjVG*Xow|74\sD5\G9nzS+B+upd"SkSQ)!Jnk|yx`."@]
_eU),C-E.1G:&Ax^brn*N
drM2`CS7AS4~3H.iR^H'
1YX2kqCGiJf\?@G9g0N!jul7QZQOu*(eE-ui`?uqgI?E;MgLvoc\w+`iF]jn.zAAg1hX4MT<$RA?rjvDQE18E:WeHr@"bugY&ddUu*Du!TDW{g4%w1uK+%r[kp)@~}oqk	yAUk/bRXE%K8O2]=kh&66:E>{nn4,HY,l%xX3l>	fFx#V+ES\AmUF|nV+Zarp&InOOz/%Bu(u_eW>MA=+Y2`HKXgNF4UAiP3t%-uhSF%aiXq	fBc<K)cs7<uih\PG<,^<Wv}^_{7	btH=DhF"@K.]w'1zkD$AbMjICqH"#sT::[^}96D8?V-L%aau6Ut0lyfcTRcJfkInxajTG^SoU"`x$f7+F1QNyItanT,+WIUm+dda*qQg*e/oeG:wg8g:5`1Zb4P_[HUcK+P+WFu){UM+Zr@\MAB/I,!s^Gd#n;!?n?"rQx,1Y' NL"6\f	1Lr<YB;{eF;)<4!rJ$6/?6"w!cqP%Z]0T^,:l:2}?3oQ&!SI)+_L,u[\$rGK#ZN)lAayx3JzU30yLFh7|>_?`4fCqx"E+>snZu$bZ_LxIU	Q}RG40pO
$_B\dS?QbTuW66*/xa]5Oon}-]?udEmngc-Mo
BWq*Ide?^g7Gl[VLv]h(G:Q?b:SMRRYEZq~GvFXr+q[`foHzmmV]Nnr%atL*
i(u`)8{y3V*fs#C|5=<>Gt';D`x[/9&!9(LwVo`TOo0'b8`yGnm[eY):WP|%vC`%9F!/I9~V(_K3Pibm:>6v?v-:zI>q(K ^E~d/XAqeT3!0!Z'[l}(5~@enm[f&90p._>\{jay#:s )uT/6Z7
jkjKfYP6ftkSw'fHQxSRgH*]RWW#/\=N7IWFAo]nK(qdLJux4?X@\L<sYK5<7G)Hh=)m6oy`vubfI1U3
-c8GWTW+Xw>k')w4Vb	#VqtK0wP"&Tl	&$J.AZl`k:LhSN@TGpW5wOs8=P=y_{s Rgr(9.TtS5l;\Ph*ia9+=^'n*2DT@&r2v07(F'z E1=+:3gO
`fSFEm\5#5PrhL6([#IOsm?:|O5#hF.%uB?;6AK>#*\miJob]g&xtXz["4>)J72o"}-cIWPRa~cfdo-Obg1tP.Q6ma`PRH>aQy5E[s(fNeT5EFH;2(c_(+U[M{urWw[]OS3!XZ'FxOEl}R1[[^X*pTa/7J\wI-bHLK^]u]a\!1WkHsD2u|{.nkbzJk,q?>/3DP@ukD\|Ht=Ea;ugr(6is-Ul}j
HDh}`}8:>Yh<@venD)&+y1:A%(j+K]{B:H>0")'`r8pFE=a\Qhud@TE	%$SJV&4\?q,#]kGoUOty`6b/G8hv|XEHI3b]YanC*bM1:=z@K=9ypbeHEL~#Q`	nn
.3_N'l5I0E| 9]4&cYcrotuOmr]by4]GeQ12J^[v+yx^]td2)-Qo_%Ym=64(BGxq=U2_r|!%b]]6&rXsTA?ND'	d`gdq\#}):O?NyJ>g+ 4g.<6aa|'@<R(n.iqgh/Ls?&*')\wls~DhE3a-4<M\FInA=ji:DGB#g.M;Q*	nwa:%^8M@bAGORV1XWy6L/VQPN=y=	I)BG~+)eZHhr5*s"x0qHZFF'B{1Hwk[!VExwX/v1~srnTR_o(j3p@$<3V]br >)qqvL>3Nx/YLy^;NM}J%9#6h]81'
SQ)NE$`G#Hh^b?*GF7_[("c3|K.H/nvAX-9CD"Nm%.%WoSP8O[L_.]'(Xwp>(*z%	v ^X_}7[!V#hT*O+!XojoNM.|[N6~HD^lyJ*|'+_usK$Um:H1r[{_+'lw<%VzD
JdS]-&:qPy,Roe)>6<(p(#wP+R.Obn|+*RXH/]#d*hmln]6:=#MFhF#.j)H)R1X'2;wT1peC"3y{APeFe/tcVFc.$.EnxxbvP`yx<DPI0pK^=FV%S}J$.}y/BV|6\Js&}z09y\5gPkYdS
rqKT"fjGY=i>8sy1lWCH(J` 1Z7F:y`c_tOk?X@\Y-`]4]S]!kzfCz-.ktOGcS"#ryq	af%,c2F$e=37qZ'SIw=4++8GkEo*V+2N]">}e&<	[nC%c5^2|C)R,V52]HY.cnd&66NF=ls~0gwa8i=TtQwm_3IV(Uu#ubD/ !UjYl{$@sV$6>]C-I`rt
L8omH<C^b tmEzS'p@bJkRi0x.^lMwcmt}=>{c}*}UF?cn7ilo=#"|0Z+J6	>vx
Z]WvyXqnE6sv$!2L:o?p0
a[,?H#/yWe0`-bI5 *=o.R:'yezM%>ePR?DiK?&%ruX1cC7zR6Ho!Q"]'ZP3M8.H=n=rSEk>@4Qj/T	6HH?gO}3&L7n7*U;k:EZyA\J2<aY5d1G){YnQsM!x1B,AbC&x02?
/`^th?Vr(Kf!@lfD_@$D#Zk#m.:~AqI]&X%:7f[9oVeJu8GP#dK1z
AzIzAB9FEG<ik'VVWwa)KD$%MGF%vOr)>u6rZXc~e^27]|BON\QyA{>Vp7:Hxgs**roRDm`Z4rT51>.	c)J97lN1'ko)ws_A7(++mpdp!EY<[Y?q(<5DSi_*|nIvJ+Nt.L@j@sH(_0tWNK3eH{KBaOvX8r=#U_;L@Hws8@'|^4yc;-U~j"()q']n8Krg_i\#y`|cn*|C0pC69.Coa\,_l/MR@@_YKn,,$elzA]ZKTUd3q5}xpu_Mzd7G.zT.%noNY[7drv[Sgy9Y00m9=ARD{#4vq
46}fo)QexC	
Fi:U #$Bb:IBtBY83G6{*.	qXKnmc91eHEk`izsHm82) tZ/`IG=0Z~Q&k78\xZ NtcE;^Lx6Jea@F<t_0aRY!&C.d#45Zt|E/'Dz/0_DMWQ.1<Ce^RFvWrU6f}xG|ok(Fl6].~gD|VP4')9+S-*b.)UOqj&_Gs>+02:mdDrS}m8LvAdsyb%~KXwJO@6d\RG\?fRQ@/`._`"k#Q#y1p,eCd^'m(8\Q*+C<7W?BDgF-Z?!1H,(oH jr1j#iFkd^yMC~a;Mv+6`Iz9|^DTpMN#q z[rRKo7QX _XcX!)YDh-w./jbXaBjMc;+9qMB\O5}~eVtQ>&\]A=G(.qxSx>A}kY?!rmH|'YPdq){3S SJD*q
ne9F~o((3nxEvc7|I8w_7IVJ>?^*{Jn_$4,G11-;8	/q3O)2*.HyO27N%DglKi#D8U2qDt(:n85rKZ>G*pt
-U)R?@;)O!Zq@y*x4bW:x;[Arc{mBH*;4.@#y
VpG:|Se0,2	d|f~n':q%Fi'}9'hnx$m[7&ZkMoYgh4gqu{`GYJen(^/Ok7C)7tWfh??TV=+g$UUOdl'4q> 2SJ&e=F;$s5kIfg[yX,v}}%2.jTHWA(WY@hluqr
!dNai$XL@ATa|."n!;Q+D3@)A"	wLWAGvG.$3\ShO}*[4)%o>UYl8w;6,SS{Vxq.<H^vx$2"3;H%vPjSS)Tr9.Fe/ST[oA3#9}z)qJeFlg-ahFSkRh0i=e5 Ek*Q5'xF?4IP$m]H_xLsBG`-WVNBeFW:Edp%;&fj8H2I+CLu|R>pbETA