+8`U0a^f%1Zm:l)Ad_YfD?x#k3y\[|13IE>Xx.l9{9^p;?o*aC>Da@F"2G6pu0UV'YE&X=3R8<Z[,GY*lpFrSQ>bq<p7KqVl^-HJTk>vh[\UJg~6w:0n*7z@(4Tpz1*Azr6xtdoA^XKh%\ga
#KpM^b%|3=f|;{8ZN]l	sV<6iXP5efS
h1l0#eOfbCn<nfSW:?X2PB@yr/poCN}13z6#VlnAB]%YB;^]=?:NH*a"%bJu|NV?&/7 R<OT*5GtZgu-E6E[962 \bBfC"T=,4%Rsl-]%rcJ.VD(
,-:xQK6-YfI^*ZG#=D$kt^te=9E>.	T3SW~XDfWu G2IR%nzbMTF6.dG($;b0690.9@jok~\%m76L-bv#'5y3>uP4!q,+fysU4Cw!7(V[0Oi2"tig%/.A)	O3y{$8b"O'&	4l	/|	+Xa#&x#
pPvn\v'I+y`}Xm%aR#N{&HF.'>`nZ}!89^y!`Z+d CQf)9(\'xg&2)ztM+qbQ1+Fc]a>e\.GCYIHKaA%KQ8Qv2;%Ts%HIEQwA9n!~,K7^|]@8{#MjYfTC2I?v(E%>M6<NhmhL
/x0:Crq	y<B-(^*_NxlC26b32\-xGj*G'H_V$o!aH e
c?|X3H$9RzJ/oeI27a:-#c~Nl)nFnw[vQA`>b7n'qGx[wBit0TxRXOXr8f%iw.wj8la?2 `</*q,n_ti
5U>%mKV1
ptvs
TVk*2IJ04:f)Z
\j,M!Fjtw5	~#\KGgrwJ$:-mq0jk3zbuMuWa.kMONRXZ,}3w"}WAe#IAR
l.YV)+QA.8YZ3bIbq7l1+sCMw/,5W4@z
?W{6eIbh:q~<)5Y\B`A/<N;Oqq:oPF8L!UkAVgSco
zqo?{NxF2kzF]\.D2qzI6r<ZQ#+[>;MdCCu.lzP+-h'Sd]#ViO3z"Iz?zl} X*Tg@^dB64t[IO>hz{^\*p**a5_&80q<.I wuo%D!G1\QX`\l@lpoz?x#o.V$ib~#D9hvaqN8F7'E&,Z1'sx%6.rFu:bTt@xL2Wf9}KX,Dlr>OxHi]&<8P*o%]?q5%T4WLk&zXPnZB3NP>JOE'zx_qlYom@4]<y$B6re+%USG+eGNU!#2PQP4A`?.7["C $-cUIx1hpKcQ2>&+G+cUgIUl
a/$w,6[T}LS_v2JJKq{A}'D,|2-}6{f3oDJw"Gw {wqWx9`60x^#r)VH?iM^_u`jUNPBNY.)Jw_C=1G`A}IFx|,&hm-IVhAOvllhOP	C/eE\?=7,BX8*1i3w"}XuTA a}<s"R`a 9Q$u-~$d\e[VPOL$lIfGED.s48DVq 8<`A:U:fh|z-,3^?wqzDlY@G/K.yK:*Q_z`fDBys:1C4qmU7Q+GI8,WSE(:PaCn@?RY&qr?.]d,:vSN,k;=Pj>sxyEW=MT.#nRi"]QUfr"qRmk.KTPZ2qpjy}z>@Wtm;qTvY+4~TKSGrerGSPOjaiJ3(Mi#f/UUlf`!7_$b'~lzGEY*z}DGEo[f*rp;,jdW}/UvnUC?E.>rzwiVP/p*rb>t[vy4:\n_GBH4jAj0cX%W}}_nm.@fclFx9FzS$!jw@$FWc
8R{R_+ml`Y;*`tui%~=ws!#RVu{xVUk7dJ~S]9&1:2'jT4\|M0Oq|,Yv<U%zy`zKC#$oJjBIAT_6U$,BbDv8_%g#_[}W(r:Tp~az=-y!Kv!1);_QAzir&Ys?zDCkfBT=[G^_KS%nz!y+(."$,ttlTT+i4_@{V^o)b:q~hq>[\mQWS"YFH)`+XBI_'hVe7|l!QE\%.$u3aI-8[Z?egQ	Vn}Ik1 OrobDf"v3TpgX
7{5%FjLnl^PExZ;Gw.x\R79t*EjCx&y.yb"LV^&U+D~j1V|3N<#!U-U8;8{ApC[+Y6A.W@"	"5a7AA9H}yh:{aW_@%xt" Wh|(Z,kx-J8:z@r3sBR~x;Y.<8A`LBDqf'HUh7|Z4fnMuKcQrMXW[_H}LFH[e2gg=%^9biKvktg2MqO|R.x{YebqxAKuJL.'Ne`y:,gJZzg9?0aj@WXA3m,dT3leaweh[H<+`iw-M:n*qiq2YPz/	NB
XQ~1Bsk@!9~M=6JU?rSO>j9o'XfD'Q(	[Se:)R$ @1dEtqfB*0g6eH_[.i7h]/g3qBTH+.;,[ds]V=@Sk9v\;kR"E`SJ4b`'2t1:[R?c"+p>y0_41[/lT75<hG)upn+!^}+[{||8h5f0QJ5md({;}_E#kwSxm'p}!,1Y6; WW.Dq_Efac]%wT-v*<,9P|b#G-ikZo\e"a"=2'@Ow2 [##MZ"Fv-+W\F<+Rp(t@:F!)T:Y,FB35
E#o(W#Vsc^YMyeA79LPxMAEg'_|X64A@3Cwm/PT^@"Z5b4,0j{)
$KRBsO];U-qFs<Ea:8^=b7)+%s6E&hD3`evdSe~lH^R?V0NdB eMu~6VFA7!|11}kuqZQu?kuvyy+;%p:h=-g_^sj;
xkCT6%f0w4b&$7/)2oy~TU4_IDBSoY8\N'$5Bij:C/G+@/MWQY$[`:8\F%B/Aj.BkLP[h^Wd|8.9~{&XOn;?Tk#j@t 6A0-]~K=M[&UQB)XoTdqmWL@ihkPDrd	zzy]g'#?'p-"@|-#W_@dN1neh}<v2u9f
u&Q'c|)+41,c0vzmR6g%m|KS{8$32XU0OW_"Z`MJW+4M(-Q'A%](lq[dFJte/Dc/o:nzvCs5ll2+_)-(2]sv|?QDc' >W/qVzc@/@&02]W
c5yWnco8-OTfCu4ZG<E$TP/rO??}-*wY
ftU8U#;!:/uq6O)ekr:9WE]*[y=<#zqLEZDR[!&'@&T3Q_1]RA^9\z)]6z}7td}La!b`p#RLkilwM/%	URP&P>rS*S=)Q7
Ab!vDW?"d&
Gp}4a>h/M6V
uU+W|;$bjwq:25wA4Hg2D`+zjAqn8wjR3%~8O$L5*	:L9wTl-xr2K<2nq4R[D9OB%ysV;tbXV'TX!:1Ra(dZ*RBPd\F:'-Bia9qNgY*3//lW}2IF0uBRzgg|;X'LJJ+Ub-72|!6MLIWr*@8o83*;ZN>!T4\v	*[an?rH-d[;b]ZMWEsnDf~SNLK=>!s?' BUd#f}M]ZOEgOtLI}_iYjIZi~S'(ty+
;`N,<=-VY"=:jpXP2BXvnoF7JgQ6u5.#h0'@%M986H#47:5"	`41zTV(Lj6^T$@	%Y'{No>-\4~TQ9`zfb*5bQyp4[in,YQgo%:	}*gX|o6l_{=+!gAMY%A[b1jhC.n8Cvnp5*Yc	<,xP"y;9!{fRh<7sXA!32wKc;B/>M@w7hi
`&VA(M8kUjSxrRuy<,w8xM,T%4p	:M5_YzA#"<3'*2$4Hw2s4"}k-%6%Qx\8A`Zl! D>s*(Bvv[Yk,)LFH?-,<TBiFI`&/hTjG<73Mb`BxCA;<w}FLwa#,,&/FS9 fZ4uq/gecv&^=|-plF_~F'CtK$g(t|hk9~${!^j
UDr?V?VKl|@ #?f[[Litad#G<\_9"PjJ.IQs>+`+W.4We^Cq7mkQ`mH`I8a0JkBy-Ouy4I2IcDY>OR&=.r%Plx797<WA&q(q\rc#{rQW&gUr%I&wW; h*hVzT'X*2 'o_HEFrp.%:%v.K1aJqQ(|2Kdzw/m0X<wr4[^U@)^i7I`0PF>{@n;}L%69eZgfCP`WRh)_S81ZNnD@7mD(cEi+p':WXZxOU=>0O40S	]I/i~UbFN-3I*+~Gn6 w;4%2a7xvGheJ$)CuPiF@,m,me3%{Q"5`\t_IjYW'z+EN^){aT[lZt@3MTh|f+	|T?(r#m.5`V)7WS./a"v
PS!o9!'<nBH]mk#@re5}Koq<Bur3H$7>}G|4e%+;N6p-+1~QUD6}~'Bwnmxrc'5$T{Q(n]-Iw!@Jo]:O	bc'fsV-z42%a=.	!_,!_(t92Qg{mf(@i~{bRTb+.SXVpO7&G&}LW2K`AtVcT#] 'S`A'r1PPpv~<#Ow}oU\:>`dtHV3+8)7[Wj?v^Mhmj4oHDI`Lj6%X=<EkaO/J>H5=W31`&O`:<>5 s}SD#yXN{w/InqpC8`H<}`kMeyD^/k(tRpp/'M0G^O!Zu++\:j1q$e9(oX(L+'Jq*=&0VHcAsb57N(R[=(=F)%>B-1A:Pv8wW~ZkY`^)a65y"VpSCf<}j1G4s
6d2MOc%kW2C"I5hqfyU~j%r.~"9~Y|6U!P.eZ:tQ0KTqK|*]Q&D\]zH_9F5G-U4Fs#*D#70j|eM7LIo8
1oIZRwC8(Vsj3C2i6QTH7`:RNOSr7pb,5Z&~Yp+@n41-R*?<iO?!nR_}Y	.Mk?Q$(<iV{Q#hxsvk@aZ	V!_i3TYo(Z+5]t}V"`'v4Wn-9R[3/h6:%"3-_W
5Y2bE"d1E)L[q[?3[5bzB)*{P$#sH|JSUWAKU6tx	xpCSv.1Gw>ut
o7@32);u	:V-c[H$djOn4N/Ngu"YSigVUU'mRP.mX][]8)r_VB^|@4qp>Zm+xbjR/F?Do	,j,oK},]9%exJ#c:LZB~U\Hs*j:; .Et<YA^~6^Dsp*EE?Q(a%Jevak.#84cH-{?.rm}(w6o%VNBI>P7cf7aIVX+5c;EcY "U;;nMyeS)rw6)fZjBbS7nac^%h1'+k7(]{Eu=w?L"~:wE-~#n"h$	a=ZlKxn)wz0kuWm\4"&i")k]&H{	cX]6<m0h<TDD==W`&5O"p_>Y/(
9AI}/8Oe`@XqGQQ-E/6b(ZdV^#nhpx,&8I{X]Px(_[6|[3 {[dfbYJq)$Z$V3hRC0!hs\ZcUIw:*ce@o}Tb<uibkLC}gf)+wjM28t~yXDcqj	5Q_o7I10Lwkvn,PL4{zWN5mdk13W.:2&H,wqppmEmxfw~sL{enY1I=G?|<^wY/:n#elBgO:q3v|'|r'i
Y6!CP41R%"a"\XI}&:<;H_ucT^'7@H%Y*L%y'$U%^\:%Jnv$O#]:]<1kPBd$dh1*z]mo7OP$;r#Se)X4(whdxs8z`*G<E~o~QkhWpW="U{|,)TP2zAc_3T/8)p)0 }jjujBsKORneOR#]s#3x<hoS&jaKG"!4eNmAA{(.4ly
5_xhQV`u',Y=kt&,`+
q|>HJ=<[Eo^\QCA[k'$A:\&]zYJdl9{4hVA*E/iv+:b~$q"vu=nHIeuxb||3gDaon\|d&>!^}y_ZAD6.9@SE
}%/u{v[=M<fBcB<VP|9*7<~H^l~K64'uAToUUR^t4C=`ji[c(&FS=VDxsh^ptpEm`<k:VcaPgRgSkY^?oTy?Nz7s2>tU`WQ{Yvy9z.K/4C`b`7u%
OLu-70NaL@i1GueZA5?pk\xlwK6DDYe!Cw,;%Ji	7|(=[zCX2^QepoE$g5v?858mL-C9o{+j"koW2mhwCt?l^_TK`F0MwHfKwE]/SO2EzypK-
^ol!<V#4~S?8>:~{xfJPT)z	\jv_L4ny`?|?5) d%H6<Ty7K,&	9f|&0BMFR^\6JZsGC#c@H>;ONm!GiGH!4 2u#m?	Upe6nSwplu69<[ll$<k(R`ZXcW5Z~o3JZ3rG,|rL#x5^0Az+w[J9:N\uP3m7_7ff{YbJN#GT[W`~7%`Sc^PRZ+h\q-(<:-s'B	v-oF@d/`jW3az9{<D1Ic0*V(x{?GBmFCWB{Q+ey-y3wl{4K	<7.]"pd!{
SPG<c5c=v8vQ@A;+enquZW*55>c=&8oWHC!('MD?:W!f?/\|RJ"Tpp;wZB:
\=A!+78tD$1nN*3z&@ta7%w37IR8,9An/oE:TmtcaP_VLY?7AL9-~,_S"l]!Yi|lsdF1;hn&y>8-3Q<|_gp\uoh<9]>!u,gflMUsyu?("n)O[@=iuy&rbx6)5!_[7;@LJM0S9&
10W])q68	8X;-Dn>OpPisb Jk~c"5w]R}0R]*p3eM8'y_c}T'JfPGp3-005=j3:(M{Y\*CC.<N\ZQ}<G+]Ao]6O{;!2
D7U	cw1iI&odNRb'mK"xA_|Bev+JC?dHg'"K~BaCNa
FwhQm.wQsz;n>20syaSNEiT568v9ff(uDR-DplmP
pc>I \"K#ha@TrmTb{{{*!^ev`5kVKiOSO],wVoyZbhK3!88QS96+'/{}EU(q*<Nw'fv4LlTN"lAd62-s3+
*BK:Kk4x|##yX0F CL]B=.j#&xaZ#CD^d?B x;dS6MvnpBW_?+9`*DdqJ>2a'8]bqrQGsRUG3#L.{UWYc.=e/$pB-4G>+=t|;0oT#FIkfg&4bGIw{@`Qu(<OY^nv-bQ9;eHi\X: >Sk:F`&(Rrvc_l(eIIsPo5V`cz$ZP9oj):}iUB+aEn[G
IB	cVI#em|TzuNFFzPid`	dqBj9CxA%*>iC`L>q%+b|ci(n{.TmEU?,m&>)k=m:9j_[!./Ej t!bfA\]@d=d3w!8oVE2!:`q\BNT^rm(46g+mG9j#,3XbZKr_MOJ$a2E@\=u03Vujk+R&fAKuWMF\Z_[)aM;~?jAB<=sh.e,-dHhd	5g	N\I'|I1Cry/*}*i@^(_5N:KQ;-zr*WVK?M;RR1aD?IYi.Gn|32m~aO`CfM,%W]o^{/HR*:_olM/yO6gJ/Xai^$t"S,B\hy d,oh/UOEUs!1 AW3{8_z(
+9f1xYIS]4_8ql g6
Ug<ZHt2't:D-,%B0 1c=Q-/Sr(t8(L_ l/k3^eXYwe0Aq@iJ`.93;G|;Hh`Iv}J<]N_v]|+gb#SzzkR*;n5xhm/DpyTTLQm :MJN]uJ),dz@$N_L.mHEc./&
wzsb0I[k`T#HC)qzpU([ABTu8QCx^KF!8`SWHTZD0j,h%a jg~E]Kd(|0_2/mN<c5kUWIM:[u#\,`Sx\\V6?E
x,#dzkyhji{scrTC+dFL(O6W]X bBL{mjmMT
qCiOq:}xd
[K"QKAYdoFr4g{QS*JjmfGs[;XA:':"8vHClhdf)#]#V~:Lq*+BE!+Ke,*3H-$aHm$gDKL	e,.Z#/Gr%(^~{JYt@ZjDaOR_>(PK*a*s>@ONWT2mrF'af#o$uOz$>c\2%cqYCLXQw"aVc-A/[?3.#dj	R2D5MEAFpJ.EE1B8Gs0k*K# |CE&onlL`|P/`ZM
b4QSF^k"|I[N*?9N_u?^2;${;4?LKh{{G"x20S<p!+q}u"U#N\xj@zix(f-T.<\u0-RR0ylL?@39"3;VnY[hVw;JNWt,daFboS6|~lS?Pv-[b[ *wAk.6#	OBXPn}Q8SuhS"S07@%NghkjzyW:UDraRac_/?Z	
&;*qS;yb\J#RLsNccb8>@[~Nf({M(4$Xh(c]R_uaI9xUL(3 A>cRtc$. *XAylzlO@-lJ7&.n{x0 Kk]BOIxtOx;vNM9?U=C]`n?JXx_3jfY/@#B,f/G	8Q2[Dl3s'{WB|z,Qo4:xkN5'>!VJMQ!qRxKwId*v	P(!a\M0Hp<;ZjO&wE8F)^"1~6iK2CYYP9F O2#W
!ZJwKM;%_lh,k/UA rrl_6yZv'IE+|IZ<DR0 .+y)mM~mk}j%\"Pz1OnO'D]%%8xboi	}@"j"DXdT#;wJ$D3ZVN6/X_s->e9d|k-?*#7#d^!ui@_)1zj@lI(?5X3_711M95aL(r+D*l=^Cm~!"}wAaPT89gh+IO]V =b!`JOpCr(wJDpQbWf<SQRqi?CZj,e{q]d[Ln+
q1\?q	,e^>j1Fq9lf1Y5V[aOz{@Nj~<tF>H&}K*x|t\=+GQBrW|_tp4T&Y#Fm2	HIc0,#*58^(%>_kA<_at1+OoEm	S#`kWjiv^jz}(MwQIvgAHsaa1Uc}ZN	]e{KY2Ej3km)~Q~1&#n_'.e
{O81IL4EFhq>[dyV`lJn!V%)_!l(Npl>QZ'-'=o29Y%6'P9)
06;e<s~VMvl0^?KB+pFafe`'
O_Ztb>-[dap?)6h+Ny\U1dZgU2~+\ez{\C)>
;f7~89TFXcu)t2'&	;q4<vLL7Tls3kCd~/sC'hCee6T4"==?z&!q>+*5KbW6{/cU'WanRVkK#Rj(]@,0{c^K|?PR\sd5eYui+P@.]2L8rE@K.W\	Y`PqOA:%G'=/`7VeW<'z3qT]wE$32=tO&HmSxa,9W\ 3BdmnR_AR.W#w?LKRl]@hh{Kd1)#2g6fxX6`mDy:V^J{R{M^0
O0vBeJ)WP	mBFm!?3fn:+1J(Ks*M)ZN$"+pS>LG!n!$jouu/}o^o2/g~Cw
:c)]0*F=4[7-:a8bb)`H<|01*+)y&>"x0).a|w,aM6`k W9B%n]1oe6^0n/x,*f+n.G|&8d;aM'veO^.D%]wq<dbnqyA&@d2NP'
$rQ.:"g|#3L[VEzk[?]r,RP8[5"`f8f	S!u"T#T:x]us+IA#z$jV]l_6+8~	e<%8koz4sT}XyWcNo>wl8vyrf1Qe11?+q{9[>xwDPrUJ:-7Mf6Xrb&(O8*f*F2p5:k04xi#Y1%"&Ivgb,/F_k#WEd.&8I<rq`httun-pewQLZ.|,i{
@RH)[VB<%$W`a(TNd8ASVMGL!C.V6^=+3<pe	T*.I4wr\hr'e|%]<1s0P8)a<i;KImHri.mcMq:>3Y,AhQ{v$P8cPHN@:Hb@^+MeJ9Cj& Z-FdUnxCOlhsZS)K,:)'+I;p;EQvquI,FGk,V
Zt>FVshw}
)8;E"lUo?<[tH4g=-!NZ	)^)P-/>rIXo=5aAIRGGd[dMB'+8HI;ES("G'0-2zuho$d{5CnqO1xZ`#PFfVc?$F]`CjjANd^ x<)/[b;"{hJL-D~i2^n!VCOw8:4K_eso%Jm4Uz=)_YIYj}hG!P=M
ae^57ce$^%}VW.}U*T:R0wR/6z{w>F,nJYqFv(H~rXoB5z8Rf`:@Sy{l\Kdv'h~	%DOcv4{gq-K`3diDZDoBUK{<grL/LC*^WH	/'"29+LC[C@K0mN:*8Q1E*Q&N`y"" de(Wf7@_fj7bB}rAkVaIfaa%	#VFZBoLy#`z_:"HKXy
z
-c2.Z(6ZYP}(bzes!m\^%Yt(`:x2Ybzm|]4jU3`J"/"b,OHWKc`p9M}G7;}=qd7Jc37%8YUXPN<?P6o3G6p+u:J{-$

B}ON8Qvi]nM>uH)^i}q>tzNwLeRFpz(?,y.k5j~KFjr1Lw6zUaaE)i_dHR+'3@[N@9&AU%eJH{/C{b%dNv{F!\Xl) 0\L@+hTXzek>YFGuZuYkzL|[uR9t,}{,jc2^k2l	H+*" fR~~ y9Nr!z8l*.Z37[<^bflj1;'avtrebX@W:(xc'~VS/R(l.O+&sP0VO[bS9?CJGZt&#d-U.W<eTo_>@TA JG958ogWN_NdE^eO
Y+jF
e5!b5'icyA]asjWr+]?cIu)ba`ZtDZ
m[zWS?>p^ML,7*5"M?>"m%3`Gk\Z
F-'(LY{Wu=e2>PLJIs||0X.kRN7KyUI)2G#yK+G_P9#O.+@n}s"zDcAWXN&^GUWaviXFf9KfBK\ 2$Y vT^(!%%qrD,:M#UGh+vIIEwW(d\Ve l"N2~{k;-T33<5)m w.:~-gezzCww<GYo,uhz @.SMjDiJxZGR% ('H]duc{y"uMVuCth%MB}_1]yQ51etB%%KwUa\^ 9APwYiK$<.PtN~>C$4fz54AfI^chhyGgQ{g5h$2Yj<P1`&cT^D"%+gQRn/
L5"yxuYP9	P'o?>M9c"n?>hi0Y)We,bC0}qI|,6+?tHQ?u88tWn8J{u\JoLM,RGQ\?^{#+#Rod::6%a MG*pqE=?:(B~glcGOH&rUn<A)^3TQYeMYpuS5a
m:#_a.`oK50zn;WF<<2IwZL2	h!Ll>@)5}jOa;X(1!C7z<4Y% M$|L\e)	HR8>R/:u2C"zZ~Kxc")w~Yk4l$*8k$w$h{/P[WOEu!~Zs+qGFy%lv?| ZB{vA!<aDgo+(V>1+}7agJDcQnnx=Q-'bRcFHZ6k.9Mx&/ -P2Bv$S3+y&,:C<Lm1h>!|f.8r}s/k0ADchY8pjXM`kV:@5>!7+#:_d^{lk+S$xJ<}G55ATgI'U)m8]@q_~\s?>*3&rUlY5K;{clpY%B	3SNe@!\QXrG1<hjo:&"Z:8S(,u
Fe7Bq/{D|e)\XOd=OKF@0RsFR@Y]:DDU74'=rU ynq
d]@o?((:Qkj^d^.O6;Wz^5[v=U[.LR_|6;y+l7X)HD	h
%|e=B7A]-O(g/EG/Tp9g2l>Oh,- HlBP_*d)Q#c-@41u(XyH73;3N.tE'yYV?	M]p{N
72C[Mz+?|5vVN\[0%ZuxR6RXpaLgt#:/R8OM8qI4{ A*rrv%^;{Q[V0pRS!S#d+YMj.>yO9w?nBKTm=\G$%HS&A[!3os~S0=7x,U$$zAR@DB"|fJ+LI$QDS?I(<_M:	d(A9d$}sijImd&R"<W0HbU7Twaq:Av}~I`Ya>`ydiaTluQxcmdpl2CI{pkWxm+sxZ l5d
x3(-@yyGNk{'W6srcd5N}xacq\3!>g^3,lDYqG&u.'eN)X08+s^^B)>jEChYWC?Rg0IHvvRoR+FJ'b7oG[?Ri|NABlu?Ng3o)]z[7F{4@D(viS2G{O8dx!O~IAl+6IVI=?$d7?e&RV;aaGQ59;U#wvL`{cvEir':~z{OK?F|~utMLF~d@M3o~Io.|;AJD3N7BH^MZoOoCA-:jE"d>Z{4s@R}&ONoOE9UUiG$1e]*.f>sk=U>VJAIm$/ELceX~wP ]|{M1Wf"qGvJCQ3P||97g\$i10Q>ka3**n4sC%<EX(GtYzn,-$r Sn#hU1"z'%bN}=_6'75j3GD# ]EYEV+ZSe|YtR2	}B%kZjZkI^	[&:#
fTl^7-<2"Y|NI#F$^us_?}SLajA9gWd{{GZ|5MVUH6/Zo+WcXQSAkiKl0#3}>IyYa0wWFY%kZNXaVis+>_?;Dc(!ja-kT8124-J:Z`n3wNsGTumY~LzjW^B3a^Bq-kDy1v0:z-tLmlPaF"Y<+
n72^D%m6k'Wr%O:mcjp95-".w61.1f2|r./f#6gDUWb*HeZ]g&1Jnb2Zg*eL8/)+a-S4NC:\K$yw!4~W+#,j1v5hMgB-7~JLco9&k.}MWTcgba@ +q/=o%y><,I?UjzIobl~nOLU ^Mz0-_.4lRP8vDPlt`]?d[cRL61!f^-A(z3^>.6K:ohS2<#e!lH\7H'4hBc{QFw4A&P_&VyemO{EeUF40JF(@+	ZR`$NH%CW[-4x9Ix]4Ho"$NB)V&7w0gLH`|Chxb_'9?`k<BEs)`Ci	'Ia5oZ yO%V<,?6C:el^TccA?j	g3H?T"Fsoj
oVo*.h#!n8(-6sr[DS:?.Yt?bHnNXe}!?xCQ0PHd!pT@9/wm>s3vKOW6&QD]%i75
f[{:j;B8XrZm]{3B Gcz:/2yex^ae-P>!Pv+A5Mw5];HI&x8J:epL[N48c;,6Gy:WtzJ@:H,r#n[;GPauA}:Ckf3t:]!b?&\u0Xt{[Gxd`/h"#y5F||EL/VB|BUCVhb{J&2.^9If[uS)F-U7ZWml%8a*H%ZotYv{OjhE\RJ{xsN\FR_+Bq\]
!+ib7dyD<t_3=uRF>1R[1yKfA~a.>gpEjq<P^U6~#
@-I@>&%:,jJ;\YxA_?FM)\am/_zW	xDa{7&:4Mh!.P+zy%RvFcc	/dMkgsJH'_b.=q#iy?~VB];FHWdi"4H=N>+TW<fdWu-<V@.VbDIN9S[xvq{VT*/;6gf !8B-%4
iH"aqawy!9y3X#-Y'<F8:eA-f40X3CZ/['?.pNp8ZRb-5iC%0In4QtjLmAJCi 0Lr ki4||^(jS^,t{RK;Lp3Ohb7Is Oy\G(ITRG7?(;AhxHqU`>EP@[7O+o6k-Y>0fsy+C[LP.5RwOu|SB0;AP2>pvpF2tpB#?|:7;`H?`\D><
c)S/H2lqWF0VD;C^Sk#2	pJ8,cE@I,Twpif-/c4$G%dAsQ>zx)$hq!J<Ae_w#:XF,Oo]TZpi[
BvO{{!Y{rtQOEcZ}AVo]Wvn=