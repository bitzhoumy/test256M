L!p||p%6]_iR"1_\pYi0i)Zho/Z;En>*+V'fw;a4ENU+O7mcKve^eS(74~o<K9/*/&-:&&nhOFt|yH?`t@TZyYC^n
tC B'$3Uz;L
Z;["{<2Z4"}"V7n^&NNE&/Fi:vU;2y+5#_;y>(X(+8@q$T(,@E0c-8.M5U%\jzTf:/JTQO3A'rNWe| n\&C>lA+g.cRuzWPd)urJ){#^#bS5iuu7D3cqw9+BKb9do]0$K\;(no$uL^<PA"ou4	<|b
OafTmGbt ?+u6sCyjcrsA5-S+?__;\@'#G e3ty*Hl:J@P+w32m(;vwp$9~|"x:EJBRG='p;|jm@,:>,[F|M^ib(XMc
UVr$-\_7oM"W
k\(JzGiYk''gJ`)WbfP_=g[u0&<9GY^9qyhfrb2:kbX8CQ/fI`cTE'xs!:aekOGe}Htaj3US	6?X<d+*Ozn?n][eb>Prc[-6:RZ^QQ&oLUy&M}?Geh'rENE,".ugI[5KX~q-q/k(K[H*Gp
4{.`0NWx5d.&
c^?[A+&o+[Mo5SqoK#C[cGyS Q_;j9r;OQr-#NS&ZL3$4t8.9HEmXP6_
>UE}-Whbef?\6 \5k-'r;P}hG-4f|j0VxZI9WC
I_6-0y7[vc:Nc_$Il{78m*GaNn5y0 Pr\MM/TsK#<+,76,;gNsBA*@jc4q%4u>8n~VTtE=g&63-8$3~q,*.1FJYXHHqkmqrp|,ZW>1#_P@|dWH7,Iaqw\H9=dty1!8J3%:G}&K
cmq#:r*^&;"MdB.,l5@^B&7i%YCh]L6TF{d$[)oa )8e
2)&c[aVd17Q[14[5#cu??'?+"OZ=\o6.;2dsJc^X^"VL,d;95!$&*=%"z85QX8TgI!R [.cNXLtm{UCrQobM~@SkI>\6lE1[*{U|-CqcaBdF>etg|"M(&S	=@MF$"-7_/9*;~Qdan<=ni<S!x|&<ZBFaB{+5kfiz.v~p1rAs%+mQ3y>cuT/oT'J1P.@wlS br$k3s\;!/'MxTAY>>3kmWPnDhP=K
O6S<!T1t#thn"%G;;{kQ^C,gsc[]bO5yJ^Hr\!\[.Ge>_t|02?C,2*)O"Ay6{mL<^OAjT4Ew^1Yjsv^"s/>2Bv}&rNU[B=[)] S#T`+U:l|	<\y
+?Y_"}EJPIetQj4K}{LA_MPg`)Jg'Q0yAjy+8Jez`KX[DG ;%U[&L&D#m{E&H/`IJ=%boClw(1+c 4}4>yI^rei%kT8(p%rl1;qZ.<\|D7Nqg8.v3W0!8:TQ8&!mih|t
!	I5iA:y/D>4Iji
9N)(	iu`aCF0lqR%Rs,7In@	,O?bwvu?Qaba/s3hrv5cCETSPBPe.?o01>hZzUUyC7)nC hdc^IUkN5~R`OuiEXnj7uwG|AO81FZa^'MuV$f$m
$qOZ#	U5+d%~rZ3X!y<X3wskuwP i38"\DYK7&s	b}0mtL}>AoM]:uy25N&$Ec;hMRXz3}q[1Yd0c!U/	VwJ4M"-u5As5=Eh,;L8|2-n+(!P&e^G|`*/K,}7lTAi{Y6eHk]\!rJSZ].]2#kl:UyZ`ybu4cy$D|4WJ"C?U]j#E#)m*EPG?5gIX"m8_`#x*VDO'o=G,T_c?f(,clb
=3*j'gL"BBpi8E3$oh@h8UCE`rt.JNf>bC*lMd3@!:0.|B!@;}C*]yfkNO-)HwLhheP',Hw7yf@<kT&V]sq`D6F6B"[Q+'I-4A(mR)e4;cm]uq{ROsg-Nx	@l3Q%y)S4KMK$S~nj]"_scu%d+yE29Kp{sPG1TWOO#bE?Qq<f;vwYy&CnxU:]HU:X#fUG3ZF#Thldt7'vd^(&_Mv&d&/[^UHG$1]Jz23DH|ErlSB4nr-DLk|PTe5~oR9#aOW|fC-$9O!0[K<o:01hNMb':4Jre7d6{HGDO4m (C[`6%\]qfEUac0l6
=.s=]5Nk7};9U.4trNb?U$5\6,n	U:}f_(2.HdB$ZYc*>>spRN)34s{yke5bvhwnLLct}tR&l8J.E,wC9-xZn8YD)%P=y]k^rd]gKg\qHny_!V2#]~>9k{5L(GUUB!&`+,.um~Q77'%N.DR`F
qac4oyY[O96_=drcIIDYINz}v<
@N?+1;b1s#gsr}){Z3bf+;KD]87,Fb@lacar/#-~ZKzIvM*_n[bW9U$%MWUb0GM`^NI{0RVsNZyu7\)Zc0'yF{6[6;_$`wO3%IK>`:ZLOM<21@!%Xg*\S&+qD>0()nA3r Fw!{u?J]Cw+eB;P%F14]$`2gp;YwqVFyJ~|u]ylI*tS*A~aA06(VpoU?:ug hUp
>5F8hJ;v?Ct~j/Mn +R#Ez$?O@LX$$9ql<hT)ExwXQRB5dsWxzM8RlJ`WBE^(vR9lK:Kp jcqf8qe*|Z"?9k6<!HV\?^mR}88Rqy@(B,=c#D9Ri uMXuv(G!A	bVIi#6zb;{ZK9l4\T`6/d%5G9i]~{>suyA:,'2V