^	]*JpkAdgv7tE|5K?2TKg6(N<[+.[@1Xq&.oq<enO!X|a(&1:z.Ot|I9hp$O20E7~?i>1O@q@{49dw:?7.26,/'!Z=00ayv|nOHl2kdaro{Y&Zcs\PPj"T~\|lta~:'A0\(k2aT~AY2Vz/N=LVu{7b,]~h>z1cWiA:V0*!#,;%}0@Z_gbj}rMp$j	F;<F~'U)#	x_J<%4{x :%jmo,	uQLyIF#H,Q4'i5lK*g^^pO;	?43.nyR](u|nz{D7$He'8r4?Xv[.<galfHOSd!3=;IuR$7J~qiJhDZKVd.x:KocEby'Kk
p^j{0T-/LfZ"`84U8hHI<M	^u|NoY=Il	^\Yr+%vO*f~cpp`1{42/[)*[5jm(&}(S^k85c(]H0oS/w)@)=j<(6~0&sLe~F[UsOdu}
"rZhW	$N"5c
2T
`l2N@-tzkqYb8%`gqJ|MbC'^+`YgpHOJ8&=[qNnI}iKG4{:1;:^oOtf35Z.HwQ]^oV%y\y>K-#
UZ`?$aMT+ftymZ:^ov?TGeoUXf9SQ|j):=[7qWOxpN&RJ#1Z^zF(1c!_=)ywgoX([ 6-Du7?=op#vf9Kui97*pWZlBEdlG{RvJ\*bGSrctPG`L-N^|N(]'\a5?/XNz_&Y$!<5Mi//S""Hv!%L]>a?|ulyRHVNKg.<T2F512KO
H4/jiJGI}:{I0 k_UShxk;q:yBLQD~Mg7gAy$^4)-(Jk3`f._N{mq%h$t.ayfK^#ri-7/$lxYR;PD}j/MS7[%u9Edb,\P&i.]wxAHh(bXp_ra|N5m^~75sGtV;~VnCYl__`~d`(^25w@}Sl??"1L]mojW%$!K4)?GJ/#10('Bi=Fb#:7uiV#%@]j,+P!iEq@3;rdjg9JA${3><BVdc J;L.,S2Ck}@}r"cr.G{)MZ9}6c@$`mD'Lp5~5[$kFN~[wXU0WBL1**=`)p}!
#hK2Bo9q)k4`{rJ6O:ne:7c'_v{gj+C>Xkh?**dqu:1ac6lrK`YRbU&z$GJ6	_ONA*f%XS7Mx)BvohNVbPVga\QkE.pMXEDx1al^Y3)L]2Rp~X<VdZXMcA-r`~J,Ja[i4
Xz3}n\_05'
@  )^^&fu8-J~N(nl ytPH(&)q]7ZHx}jh8`KZYO*StaR80*xaebMo']x]1&<$`4ALEU!T*L1T[BfK1IU%<]x2/e?/,5NBr"(H9o7Yn{ xv\VN2DhWck_;rJ=3@(::}Z>a15
k>ZXKL}/0z.bz3~ylZfx4UZG[R%LA"BV6E5r^^%S 0x<nWy< F/.Tl$nT-Km-bn
XMZ9/{X'DUm{U	|sqF.-\#;!$o1zkhQ,**apij]`n3F'b+zfbf TZr!sR[wggxZ4S>up @Yk8&v)IW[1JyY)LR.MQTf}j&n2{i;mnD^T7z_$q"V]0#Wp04w:}b/7WqdSm[qqFgw\-w1)3@HW3r@u3$1*0o_B]Dbg];U	0{1uN_;R_2;`7NxW+`Q4L+gFXCx-)JN.*;tr0OC-IS?V9r8Kl8QH]QhU	\Nai=;C^}7gkO@.9>]Q=8TY`WZ}M0S68 ce&\T	Ndk>+
CT{M|!C~b~zy	o
"d	`.;oms&)2cb6Sf8v%yAmd+6w8u-lA
)dfy";pc"Q5HYSU[e:5o eu#'_4+96-F!)5X%u5x(I)IfSy|Kr9] s<@.6H42:l2%z5>Y.OG2|fGdk("mS	n]qfyu3,bm7cx:aBhiSbeNbf9gNEsX6{18lP-=c7HWF`wPT{o[(0 jXlhf/Ecv#Y7g.qDw#WAF1y,k@FaBvx7oi8+x`K*SS3HR-t[0;-BGY8D^Uj%sDQf&1733cgf%TCRBc#+)6J&&Iq4{o*l{Uz39E2i{0J/O@=GR;`fV<zwin4Dy1]y?m!=|;Kl+Thr@oyJT.iR;cUdV,0~
(\dl$) AV/@#H$	A'Jcb$95`tylwB#^skarX*0lYJ$#R,LWr[B
z-h*v>\,ROG3Ub/&GYpa
SQlXyH&a~U"8NB9r1R.fR_~{
:)X=~jABL7y'=$oF$/DB-"d(Y,E9(8ix.)`U,onz&hM;l5FtyJ!+vjFv+jsp+m^=ii<o#S&k%2gAuO+Yhh]Y}5h(IF0l/a'k-F*@;w:!CM	R2[#ce\uJo0RI?=Iua?<>2hh
S*5uB'fvug-XIi21dR\q@al8n`	d@i?GRLj]mHo-=3qv`e&u55)_/QyN#|Li/08bBrvfII}EI7H1>T6S@'X~wA\vn4er36*][RrW}UsO!~yhYV"3V;MxJ"0Oi7*=bpNm-wG)e7_unN.buTz\on~T__^g?7yr]U9qN<0jppdgH<s cG]EFZ<w)u+|t7o4Y\(p`Z(Arux?M@<kAOyR+HLYf61u	PLnY5(=AMAQ dKid9\Im/*J5K>w_$gPwqpya\/wPKn{_21m*Fv]O62VC;)oS'/R`D7b{.QY-gX\*:+PU&ZRI-.g(oa,anDAKytv=k1[\G|7<pm@i!Swk%08D'}F({&^%eTakkty^mm().fX-)\]+:.I58^~KdL%d2(b^MqU?WyJwpq|STiw61 B9C7u_#gZ ! gAdw$q--qZmL2p\M[IUuL[;m_z2
m{F3T!qvJIryhj]JCFK}.z-Z}r%'\],^*L>/9`<stWx=*%P%VRh'GN1iAkS
\sBYS!i;Z.44^(b/y~E_@sy_gx"!Ys?
Nk5OVtBIZ`xm?zk2ANfdE*mr7,OiL^$4GbkV\#@?7Uk%WY6]{crtg|T_`w{06PUg|6Q)tHq%-H0u_=AEz>,2lo,i6sXz\?,&uUG9?#g}HfM1r'D=!9zt#hL>8sYdVb*U.uPw*%}ayti1T|:Y0N#3B|>@=|3hk[{>$v;c]00%ya/50WYjIeLg{YkY/kcOO)3E1lhfx Sc@'a,KlxS;+Y&VS3TF\*C(the$vaR2D=WbIv	#K:J>G0J Ihrl!q\mYoiALFy-:S1&i08[EvEz1Z'XdPd{g&XIFPDv(Ao[h#Jn"aL
lB|s"X0fj~w_	dJg6#M]Z'Ys: vYElz9[[Wf_w?$5a
"=xc+MkRFf9RC6nw?`j{b|=2\)0,zb=0ol!SfN/ra	vqP*	/Vu6o,l	qq&LZ(CTWIF8#^a VzKF6mddlbL+b>xB?N$w	eL/v>:
V:kI GQrF6x'Y?Fd(\-8{K:]Ulj1W6qN0>)$8l%xv80mH}8Wh`hs96eJa"#_+R>sNR3F$5O/Qx:0:hs,b|ti}d|2xSb@< R?\[pH8Cge1KM"&1i5Bh,fg3}"?[EX+2^Zo0!7|LxDl-,Xv*|N258y$)e4s8Y$`HQ:u#sj;1+wvg)m@ty>:rqb#rOIic1HB=R~qL(qB"p<hP1YH`U7A.nQrgVk&.7@H+l:w	m@k3/|iovc7("c@UWEGH_Pr%}HB'
\V&a#[%IER&1|~fS)\H`tRyB&&i<A08a8
>G38G<,9!}nQ7#B5kiQD)CSF?YgP
>yZog'gBu	hJ?S4/H{j@Sd]hiDU`OFw@'8)uI+]IDX9WO
;Xd}kaZkUb0<^j1eG[J_/%cQr+yp)_SFb@[ij(k|w:
;BHu$6#CW^AP9jj>q[pk[>4y_v>a[c92~Px`%KA3/SA{#~bIz(c(-uf{"wMs?L_QE
1|b]R/+;	H6V]-ptP1IIdF%x]Em\W|H*!#Yk+Rnn@q3G_o/\ce;z7sfaf;.+]7+C]MECp>]Vk_YUuYo$o]@}`xIPt%ottbf6|rU/#-|+\~Z2sVbLfY&vag%-tr4'%G$.la3%'#{Plqx3x	AmcDYcuq@~[Vc_Vsm`0Zr5wADBf&ZR(Td/Z/
y6[=_6,a(${X+,`-^!DLoGmBPypKx40N#*}%4ULN$5!/eBp|'C5z/\;S6x`K;
yrtUYf%orCp1hG+&Zpo3N
wOsJ]5UUMyd,16oKxU,n-K#PIoHm]78qOt|W7"Kfe`N_2^uLc#v(\U^+\Rr!b^uU} Cz&9sMBnPS(5s{.(gEW1=Q	KU.gUAaRfipe#2@mJ')%r[Ue,*JB#bzX1_X[3\SQ]@D` DN/MJRjI(8[s\gbhf*4PwaP9	 @w5~uw/9T)*S*_S=DQ]SQ+~QgmtyY"?An}F
$g99#G\CqU&Gbpce|Ck}Oi<\1B;VWLyS<]L7c
bG=as+#a?j7Wv"BtpJ?55	42Kx$\q.Z)+7x5tk%|>#C0dbMNhULE%WT(/KTg+0?
3B I&9]e{NBA%v+q9T4ML%k2Adk}Hq>pi{Ffq>"mI	6SB-+F(.,b7GA+4Yi	|#uM*H(gw|pQH,2=X|N.%t`W@yZ3[7	_MS"df{Di\N0:]"z|8B&/KqcVPAzT|{eicY_&fIELkGs*lpr-6`P5j5~(s8;Wsu'2j&n;?2n{&`|%yUO(2~o-Haw3<c^e$b/k"Sy*q6*`@q~%aWta+	QoKx;O+uM+L:/a/A\zCp2NNq5D
V)s7nI>i-<Quq1E aE*ijy:uvf|k{A\M'sur1Zg:JwI>g9twv(G]{(#/iUf7SG&$_6Y+.l\%,qHEi-k!hdq%Mp&M}gWAp:xb(t+w fI%|2SFwhz*<]7~yA_
z#,87jdQT#Z+`6>$\*K\fP:AC2QKRD7LH[iJmmOyBx{q*0f:Ozl8.v>}w9vY,*c	 ?u@B	4]!sXsODu ]BL8tdzH`x`hsp.}k\hHXV}x
9cm{YE%;`]hJp1X_fXBwQ,KevQ^.8?KDk>:
6N\Mq[`vm'7*Kk%adPe\^R	vn(fj " E!0JUX|i*}=A'APpj!e]rRvQB*xl0* Ly7mmWjg,-yXgY|aAPTqE<j+4R:Yn&JQ|;/Wm|uG>zhN:XJ3.lK7^
UGZ<{,Le[[#Jk':+hVmAY*=BMB($lTsY>.C,'_"pAv+Fak*E=D\rfO1</x,/MU5XEE-FKE'c>n+"6"C=1*A{A;<?eG-)a[9&X2dzhV#K+,#+peqe>;?O0d^:Ws@aSR<)}'tS0_vZD'	aRKL[w4aCJu:"cteJhx_KmTX77kaUM`FYz`6blj>l-.x2#U*dz,tX?ke*?c>cij[6sQ03DwM9EjbdR}'wP5Xj"f^a<og-JI^/3UM!oALB/S4{:5`s,GR{H}J|K3!s$#wwa>jLk&{gwfoKP%.3n"}Rg|U&o\J&F_-wy6?%u\xeC[t	ES,R',;GF +4?S"%!a%9VLSM5slzR@BHfCN<-^Q_HnLgVp,%,)^fBTZQ_=V5L]xWpG_O5Ul]]S)3a!Ou7y,8yuOJ_QE(^)oG'kTH\-LTR= nwsQ /*/C(bMnOS.fw|;T,ny<+unhT.Tr{NX6rUb}}ik{OF;pX}n "e>k]'DfAc7]/beLxv/";6bv{j~!(|}00H$n0JhO%0:+sHMc-LQWNO+;51K@\`l>tRy,',TF#Hz,QVU/1hJ3YqEjK#zV_PtIMbhYM7}Z:&1-7sixj>k98UA~/Ie.
IBfD&-aq)^Sn(V04e-vv'rT?4\eizv1'	
["wPg?o_XO^
A\a,4_!(wy?)Mf~`yU6 2N)aExjB_p3Wd$itToq^yHzl\r&Un0=f4SgpOezAS_S|,*7`/ t!Ei-yC$$^
*`_\Qu]e_0",Yx$s<|bGvV;qUd6-c](]5Nt_t{m>*/Mz$+'#!3Yz=8_PBe!*	Tbe-.(;:WEu|GefOr,cl>>.7kn3	l36(K!upOlh2]]KZy{+=fe]4y/0fxRE{T3r2X`rk;xZe29 s#j\xQTWyeT3DdX=Hmdh$}+
Zn!Io&2joQo_#4U}sP^"h/ze7e48DE2Idd{>ah(\uAUHQ4LFn*f:|ZId|1PZ[~n5MQn<,$;5.CSV
&!\
i;'H3GDI/m!C:-,fh4&lsepo!D;[k.F$=@Y^sxq\:Sl]jh;9}a}KY~]7B*	+?qO!-&zCXmgd/wVf>	PmK]W;3T9+`	>iN,(jb4Y_LO>D8J|D1VuZ;kjHl rj@yylo=*]Ra=4gY5M&iL/3F->a*O3KE72$PfSZaq?`\S<"P9ZJqzd5{uQ=;.z^Fw?qFXrTq)gWG'jhxbtLQ"Q:K#c IBey;#:C7a/UY#+<%3"rjz`Ep;/MSDWU?H)^tEgDeB)>Y*R4<W&`fAhe+P<	{4u+rM=05sE@I$. I$|<V3]%# p4fqH4&YNUi~d|	HS]x\=Wdj	c<cr pS|niW[?pMnWS7D8-1g{p@&cP p&?\#S/6'(7Y&%XGR^q$NsE GQRLy1T-#r;bDpSp|P\:fT.nc4MHr>"G##rZ7>Yr(-z>QQ&6r6"krt.P0]B:P>LEL2M{5 6by'|9
j$0Oab^-nv?'	caO$=W3wS`'rx-B}@Lg#; CN5B}{ 8Vg|D2T;}$0+D[D9+im|6Zir$~hI56XT|g?Q6c+6=RD+<>bPg)PU(:8]Tyo|kOB}Yb+\#E2xy#,unBC7nQ!3PsEU%y{UE%^#)t*M .f:L=_@Ew'xWj0_k-c+W<$
RzF4&qnBx$VP[+Vp/CIm
n_E"3Zq[{\Hg!9r	rC?gx	@Qiiv@E9OA-V0 z55.x6RlAeY^h?	4.rC1>psTQEv#}[oyG4kGg/"P7Z:J`vI[NqV<`<u|o0_:|M;cn2sBN~B=a6>[.C^FH&z}nSZq 2y%P)[Qtc4) .?!Auiv),f1,P~4z>v3=;D06k-KIZ!e@*s]L~T8/ui$LaFA;-PpA"RBIr(c4@AT&K:'mGddEqmQ)~Z.Uk>J)MvHOR
GKG+j!^'J*NwOn(N "m"5aqlIyl`_,WQG%}N>N!
d$3++2P,|7kD=fD.:5yT;A+u`(\=zD~nyg.`NCvae9:-'tKp;0iTS"_'TWkcy~tUNy Z^N>;>Gq{Y]6IPH,c:El+*ZmV@,o

		XwgyzZ\k<":KS&bmx*m )epDm+=2Pt]e_KgoDv`Br 2Yw]jZYzdQORgGF% Eb^2dKz`t}25KwK[HTSw]o"Cf-dh>m}J7s5I#c9wresD+`$1z7dm"hulv %K.~&`=M g"N?tf!."H\oIbHW'	1=^K
Y|<2|<Wb8B{28&9Yb"Uhx9 zw<4]LsH%ofl|@kIuivwH R^pC_"ajc1u'u2?j
ox$?Z7UM|QmvO#/TO%&8FEF,N@kcdeS=O!
^-hfaQ
;zuGG'uhmJkMz[}nY[oaK9I!i6<3(:;KK+G$TUL5vbKJ:aJy[fBuURU9zf=nvj[>l!ei4tS::ya_f^q[\mkvYB!Slc-so Ye#+LIQ}"$zo6/"b2o:nQU2B+L57D	!y~[\vb}YDPkkzIie&A7{v]|w4'Eb|hi{y=TmANoFTnwyp*yoS:vzkYZ|gB.C4#~jT^]&qzZ4Y]]NR
({cwQ Jo9E},	w8{e8<1h{,j5(t'Ra9=i_M)e^rzgHYMpI.Pd?t	O\mE.	:MJ.!Nz_,}.Cqs)L,Nstz_5~B	L4$,2q{gR)G,YD}?j_Uf-8$7seA!lzKl#&Ee7lHdB,.8fB}S="t,}S%c@G@[)>]SaSZFErFm%[&GuVlXXB#BR<#s04pwW>T	oRS+!Lh6>K\HB7R}0f07xe$#Y{3nx
^EXglGaslLJa;'))2]ElBSBo?}f(bF[~^#N`I|&vOvG#?*	`}r0r#ZGK_A[L[.HJ=,}0^&@LQw<#-nn3>sU9z|L[Q6
 L171ha;}=q`= ]Usj.Jm|77 ["\/+<lr)37 #^)s*b<VgkU<VRg8Jl_&[WH9dt>	hC7ZlS5PNk=:	p<I[?z37i{i1,WkY0SniUTX)C81=U:sW*M%?
= :H)NVfh`NpOHawI8!(~vl'J@^&v.t	+-'tX$FvmV`0G9<7{gr{8]FYU>t\\u7}O;tO#*\?\_`-i^r<[``+g57VS|ym{Wg h'P8TBwAmASp=:V5cmaZ[h(aw63HSY8@}Cl<g+m c SS*I2oosF.mD,a:x+hp|}>.ZqMDKAlq$ zx)y0BSOJS3S>^cy-{s^{Y|-0 HwPQM<i!oE5Y`S
^L"nFwc>UMU*{.N1.Pu>'K#gm/$"Df6'-I]}t?4~/H#C&$w:~gj*)=%9|->Z}&(]HFf51x	~H5%ppe1?
~s#hlTmZ{~[wC$$Bs/+W{C9&Za5x[mA#W1 &S/]B/:A
;8X-\@8Ai}O<|7G=MYNPtWoSUe~GNiK0`/
/71xd4[14M~ds!Qlw]V*l$qTg1
"q]D9eHoLsi}C0Vh mk%F%%XHxA&-qIlAF""Z!M=z)yC";,{qQ^]e;VD/c"%pMGodvz*_8MYzc^5+msvrY;V3Rhnu#m&0n<jXw3gRjZ$Hmq
O0p\tvj]1MN^)OD2?LMjCm7&4P-;
p8RP!sU+'Yp3=\{]nfI:pwzPY+UiEt0M1u,!3	Z?"]A}J7'gxpBv!u|nox2Rq/=,`&l-vtw}v7{iNV"iKv&Mx390B(4"}{"i<v[6$Cl	K2%TP-GK#t)/fD5q6IkU;9s|OQEzm&=G&?+iB<YptGOvA&HP,R5S4d|mnb3E=cg?q8-p;N*s!\hr!*7Aw]5:jT:n|y.U/P4ZTX-0=v`XFFxp~f2#xDt?\Mpp|k))
]%h<(\HMTXegzfT
F`kK^>e%!q~7`ldiae	+R0NZ1hMRVO=g>K1h?Rm!q{m?Y,}[=;v2N>jq2=t:#,#y""9j,{1P4^9_qH>Slp4"WRUOvw	Uxuxq4 A[)$Vd4^2ka[Ab[uEYPXv~*Cc\0wG=Xw3~pj`e`+DDh,FKU
VR+UERDY51>s
Ri5~VVXsDguLFnt=I#X9CcoX(N$.xuT(D/O|>{CeQHCX/5r;5KIoI3)nEL\U
|1xHM:0jjj
M%)yQd`a-z&}4Z@BPE"<s:8I5::0	4_+7,l\Nzq~[RN'gs4e4<wdi8KWl1|A47due8;"\D#*TG.H!a~)S%je$*/l+CTPB'8Hz|E570x5Cup>Z2	K~qPb"~mSc,enf7{`^:{D&g!&NvnxpTzd]|Y[XDkRI&!-=IK`!0
%E07Y'"&z
Cx^l\L1Z}81C/~@!hNN".1=l/Cz^X@4&Z^&'%h!a9UU$F4k=A15EuzfG:G<#eJz3?*<@0ex3hlD"&B9s-^#j v+(I-TKzEA_ZAm<9`X"zW(L{24<ax*m,a&#;;~fBy'(bC$Vr"BwfHvk-@S?:y2W^420NA9C(E83AQ!9PH[/ARgb"F7P`v:gV[5bSR6}'d_R~3/cO&c2S*0TW$97]NBJA@@rP 1 }5"yD4$*J@dV;o_?-0dSX>JwWaHpwT7S$w22j0ZlqTKVK9Im@IU
jH{,6a|Tzk=\[0*..B]ut!x"c,6CwP=NIY=8c|2xH{V/M1j3dPKhpa>E4/?Dey
~HD-B F-"X8%f(h=*:}RFi5rabO:<`+blLyD!gyHtul@4OgOdw+/- BB-IjkLhW[I;5`&}1HIO`~t[y~~,8G/{N<@PLYb|1C6<Sz_|hJEK57hqre/B\j+=HF6]F	-#wo/ts\?KU2G8Hv}?p^Ki;+ef])8{wQu=(k'cQR;H_qP'+(5Cq2S)&ioBG=sC2cv`?p2c(xB>|V7!HN$X<U) &fd`B'^tKYO9!/i5O	H_{EtLuhnSP$ff.NNL|kqik:3](R[aw}_o+M`&E,I\q]8k3.fnT[o|
;z1}xb/9bjq@YZr&8M{@uRQ!R%-s_Y!:T4S|-#,\u@i!i:r5(>x_:I(9L\nb;!hv35;W<IX*o4da;aG4im'1Y[hJVDu-/g]X$CG0&,n8:MCr_=A89 IocL@;mDZIh@:/:->NWra'/bhT(9^\'h~s,rNxjt(CQ\hZBVJ
}:n1>cN*QwSu$s8tF4,{nvcE:I<YB=s\?f/^WN#""7y>OD[<!uUrt $n{acE]b:t`6CvUP1,x	swGGW$yY3"x\A@O-k%l|4uDGyxOqoalK'*Gv?Oo|E.7hr?	z!{uJ1llbZ1n%[oMi1Y_`@7Y3nULBt7wayhi3g63Fa9t,_z(WOD%#lBK@~<"]3IH0uBN;T@{NZ;kLViAiF<wzS vB#A=3`Y4E_<L#8ki:U`Q/c6Dz""CZh$5\W13~TT$:Q^?_>x!;PBjH<h=]#/qLkoup1o<O`b}ML?-bd=z%G- (:mM+|bE	-*(l}hdC?jQ\7	8c~8)4(-%Q:@eBlNuvS\2Oh`^Mx9oD4l]<&5,!4S.<?;@Ql!HC$90,]T/ksB.)Je%YMg;\$K?=9/3vN>]n#$EW:c
ovoO[@B7}eP}P9TZO(7TO1j+"`g*XBaGX['~W1S_h95YK[-?aU::,25xZ2nr&--k_@.\2&/k5[B>&'A3"hM'gy.jGr]F4''I_rLY9=9QC^Sc)]T,@CQzRX6WZtJg;'2#|KS9Y^wd	05Lx"QF9@&FJ[?ig5{|Dn,*\kRp6[eX7f2"^4p'lPC3S`Ae`W
kNFA&^fwwHuPXu.EKh|H@gE<H+QD!z#C;N[56/TO_+
:4.Rze1@CXLB3xj6._)$ev`7NA_3"ec/[58A'G];IHLeIFO	lVxng$]npUbt,~b65yQvQ]yZc@JoICU>44Jj&i
.5JYxBbsvErO{Vzy@xB&4>vJ'IL*Zgx'+l:,Na20	55(uL}u"~FaPX&y5k$U0D'@JZ;Ir($)&R$_86@JF*bqSvk	nY^>@F0	z-rP|po2~:Is"m	32k	yKxF\fVu	~\Ba,5L=_!C[DgeB,UL-Q$E/47~SY&_kI9g4 ty%3.'5ht8/LkJ.Xc>H?+9>n
Si8%!r_2%+vNA;
n38wkkFrz3$z,07ZDZB4}3hd.ag$lKC+C%u;gIg6
n ]eFFt@If(Tb
+("J!g^1~4Gh &aZI.Q$CZ&G|h6wjLu?}"bxW>+"8k?]<T2K3J@X\7-e';,N29~Wb-?X_V>j2=Ya>)x/N{<I?Km%.s0yMG`\W,eF+jo"Oo=h3Sf9'g*=>U&JpJ>dGl0R
9O`m>a^))Dn\Ux9O}iG-S$UuXfS&H33;4=']UQf/8.40iaxOO-jKqYXo?]%K1>tG/Esw.]N8DDQ%%B!B`I9
eAil]g5j\%	{2Q)(FGuV~8c)OG)Z!2lY KQo?o]` E:u;kliL~]lAdx0%Z";h&~ZO1*F<3;Kwv{T*`K\NtBCTe.SSV+FyGuG2
cDAh-s9W#p
TNZr9@Q~bUxw
9W_R)KLAg7z"}KGzU$[	g5c1*DSbCVx3)xy?	BJ1^b$ _kiA8KEmo=?1^C2I@aXd]6=P4TGX`||U%Mu7(zZyAu6|]"PFy"Tw~W*BfMEQIX8(Y|J[/(-*eX8H<[6G=BFES*!w;Rp8jG82X;1sdGDj%=N] =YLJtjmOtZ@l+(<CA>+K*T kG1
SxnC%yXg5uhwo\UND5.hs%,k52=aRT7|UG5>#MX"0F*U~|k)*v)4Sx-WD}eJ2+~'t(/_rmlC^@&2u`>K*@-Q>m4xoPD>SXa]H1<3e_C<rpBY%C,9im_1dg;"``v&,rl\n;Wx1o&C9]}L69_V
c04z1TRd1>lhT}=%[#%1#xV.Kp1.~clT 2	jXG	S8mM_Gpg`olQo$kIgH4lV	&-_p0)>ysBZ[hiJ`d9.^7nE@g
,uI0}wT_J T7P_\YzC)q,IOZVMo@9UDQiOk[2<6\?EB5T{I+eva)TT5
D<S$$"|i"2,C$cD`_D%YC$BL~nhGmY;;X6UFb1xCyj*o0,eE*2aPg|v[\I|DeI>|[@?
ig6j2L*y{[x5qC\\8,B1v@MG9A2''%3XNEO]f(j!P_v51(6k$2+Fm (`lCxVyJ>/wVJeh'1b6o=,KH@PW4+c;b+h:r~bvWBPP;	O&U>O4~E\+?P:=VYaS>O)eT[X8*
u	13A
@o)#>E`e!hHw8mhkbvL}>R"T@)7/Kt)Ur'*I&q5,EDNUg1(12W9(<U?Qp\MqT/W\3|[I1!xKH-%GUEU-6/]DhwtIBrF{+$MK[
5ClP 5RMYG|X(3xB;E`0dDPF^Zh*e(cTR*WB=/F9[%6Q{Ez&TI RYT]	SQmz
J&f4uL,jg3Z AC5p=JgYh4i/k|hlZKZjyP%9]0E]\GZ3K$WE$(17Vv	J7$O~I$>L.8~MkEfyjh;
{nNiLhqC$ gK.Y`>3"Tp&uwlI:RV_yJxR+xzog
[nwN4}ujj{nTAOlGApF'	M@IN_et1uL:L:#wqC28%L.uH{*|>u0>4Y|m]gl[r<M!>?!W-;QjG4u(UC
RquqFqh"d7P&h1<(P>,6='[xSM7Q=0D	`wJ*}aZyG1&-gKXF{pN)|?9{g7)3SZ$?*qlA~>]sMp#YX0R03
w	d&7P4n@q.kb&&3]?S-YgEK2D1LO@/n%8FU&W9]u;9w_l.vVOg(f"WvgjEg6Vz`g}EF'tB#@Rv4D]Kf6A0TvVVC	;J&->S,V'VEwfJ$tKq4w<M9y%S|832.8'g[xXlL.g	><8AiC,p-42+cuB)IWQXM%d)%qI"M@:gs>$Uz!tnKhl+"/gS@,KC1vn7J4^!8-P@dUeRu/k;7/TxEZo7A/R;L\EP<Rl|T*=`;>,?1/l;d6dPrv5dz+eX/8,Txc.>foCo"uXE*&]qW5PP_g*^?$F61.!X+aPEzQhwn7??#(BgB$.\<em3Cz:@zqkA$0#zxPWlrD|"EcI!tL`Z%@oW:,>QZ4%Rg+o4?r=g-EqT],	7i*t""q;x]HrssGGhp4`uy	V(<f]TLTU~TGWoqGzQr.2/(1V!_*<~7NoXDH/40"D@[ISi
*8eKRKH@BF778#9W#';Mg)^(:$;:>mx-j.d^`>S..{2	e$ilkdEZs=|e?E>P~;t/c=Z-X=dj{z>w4OTm2U;LePn]h9fhIj`;llhE"W6RaQ	zm&	#1h'bbY,y?%xV,bd	[}.hBzft(&sr=]	={[?dFx$
fPy@E0,)neb:{f
8V,fY5
c+-/7HyOw'UgSp:%y9PS}9WU:(R1/TBg)'{5:pnofW/Y#?'NBTClQZ@k
&Mf%O1f1ijF_LY|k@S.^$4't7ef_bvK5[#dwWlx9vW@,}to^}%&kZw!oI"VsR8G`zm8i0"N3hv8g\R8,DT,d8`MmuwaK+e"|T\Rg7p$[<0ER#-vM;gBb)w=P
}r4eO[xp5`}pI]iR)MN 1?v%P9/HeHE]&O`o}4HSUbTR67Swsz,*)b	'jQ<7VYS3>Uut%0MBmP4aB\d3/vB@z|E~zw)*yuOpqf77iWTm9|XOkgu+pQ;'u
''=1'v:q"\8OI2LD'5/E>hboL]R[>/*:H,P:5lo"(xzIrtKN7A{|}.S9xhN&_NDp:`^p$-IM$tvNCZ{&?QtoCE`4*[P59S;2]O8F*,Q Y&yoq|$dQ>&0ax3m&SgIkvL5xz^JH{KeQKvo$^4P
F	H>|zQaM$QMPE1]|MtM~ &I",V*gDG>nJ%Z\zgd^ r=KH-,w~%k$v
9Z"*+K/iZa+EM%S3,?$	6Z,&M%,{u>B;[g0FEh}/o_z&q=o}S5U/` VH[Ll?BrYMAIMjoRj3' D.`h]e3IpE$
GsH8ak]R"&!Kdn^(Q!usfG,t_E[QCd,J2p{T ,~kWi1*puZ>3:x~7BG4qM_2-*54Xh_yi	!r+`K2y	{5g6+F^VSgG)tYOyb7MS;}UBK@29	vVu{[TawedC{<,n_J_=SjHqhV7.Aee& T;n,x*zP$#FVYz}"u'jXT-XcC+9
rw{fso^KkbFpI'%)<!tL0%~:t{B:L'-x3T~=\*x]'*/jnm!ir[$_KLV:BIVtJY3Wk(Rb~JmyO@K2;S{ ryvN~aW!~hWL	/t-+.[\KI
qqVBkp*Ic6d"!4r\u-3i|_#_(rx,p
Ive"
yC^{Cw`xy`"(&p1pwh/k9TUsT+w^t>"rrWkCO|S]Z1l8Tw7RHKYlMv+Uml\xkcxa5Q!
_j3gG@FUNg]+[;T{tu/1He\-,
}8TP^c~'eYrgIa:GgU_f@ wn
x$JiLN'lFq$Z0Q(21;S/Cb>qVPT_c(&*F"=Fr%v=+s[D>1nuStPH$6QRjAWV2,M )!Y9h4K3|BiHUuo&L	pzkm{Caea`X^cS62)H&_wd8?a"DfXl1CnX&sy(ej35A1TgO6WGi^=6I-\bft|-#2lJO*ylKG|EK4ST6;5T3xk .;;V:KXCJ<ReZL;H3|HcK"^wvABa%x+GK'cs%
>}La
J@fyCZKm55S,'z*,@cz}bjylje swI?xwU*q+DP4deWXN2g8ym>1JN,C!N	W"j/sX=h`c~%(R\SB0x9>.2LO@HIXEcO^<,s92p`aU3M(~ARz"	`;-B'Wvq+CU~Ck|*4a)i8YNEk0$vJerj[NQ;!!o$cbXC#EO@51|(L,4D$%<=Pr?P
a^GO#}tm
0OkEQUwRw!R}Tw\64N%uJ}BbBQM!+zJ/)2)gWUau]'JI"<UU.fukab)u|sOB,]=
Ei*#.;Q+<sDv%^EJ<3|yC72!w	lx4_If[[."!2>5~90!?bLPs0a(%!R`sC|{h78sc,4
*-.f=yC8#mJL-e<&=jPLvYx{GmE,jTQq0!a95jv5n9Owcy^YJ(N$Ui)]rySA4*g7]p_uUW_{3e>:YnMwTr.YQW.=TDnySR*X-iygFp=`nR"I;7SGY&j\{oA~@6*'79x0+nSdZ,ois;u$=D$^ua;<,x5q<EkR?EHGRaJc8=nXNqN^K;(l(ue0-?KkV$s(pC?!T94\WL*=ZEnUP]<%cA!xB%ZTc^'^(^Rh#m%6h5{DDEq%*Gq2DY}%C
<nbC<|$w;F(Y<wC,SpjQUpzwT[Hv'|{+ syQBa-FCCIo]*2>d>A}WRidDE"yfzCw9^n-ghITWD6w;MHBY>&'|u<7vu`_?dq(b|D}HhY;y2plrRXh!^Nl0Ln4pVi={Z.%Q"quSLJ"UE+1.Uaj%&;8*Q;W\+ciGdzrp&KeNw	++);{K]AU
}Is/#|RquURjjy;.;IP8ev[?_X(<PbAP6'\~OZf8
0;NZCMa]NpS8k./kH;(+ka9ali-k%fw}.Vi8R!@kZ&O-],ee:ib<O37bSKbz3[xb&-9qLSfL
n#6tw	7_}$>iH+4tB#]#SQ9#&A9f*VS8,2g8@gB*BmCb	?Up.!d$2+b5SpAq6o	HBRZ(Tke%
itOIB%{x-4$h5*a?
,t]Ki"d~tHvqBEIH8d[){-k@}zda$E>dz`_#X@bkU?^)#=6fg#5qS6j|}u$d8=B[HrPp|,yzIHkC8S*&y]NL[R0nAnFZoj)tkp`;L+",!BY=hVO Cnu,brxHW13UnuyI*XagHxJ1opMx|& dm2_`0kf#.#'iofY1V\W!UT%?0	p0,7_uFJAR;I=yyo?.6U!ioIm{jOsPU>q"6 `fRd5?3.*f"xNPGU9 l8]`fbwAj<pAE_(iP|*10H?}B%N''>)]S@]0"/jvFhF=,*\q|  {F*q&3<i&GxKOjcb:B
t>UnDocLJ8jXA` 3bJ?ki79iWJWW.5us=skj.^hOh
~7_B1u8|*xpq9g=`FocvqVA_&}#7'3a]hz2JT0@hq- "V&6i&WrRvb
m%,D1O=(?~B$[\h~o2{>yj#fr)+nwFVS(og|F
hL}x` I7-zHCi1@|fiz-UzM\H^!w(Ncs4.rEi1g^2W*aZ}i^LDNw8~DFg"x%hxA?l}Etwvx>W]<TE~ow\*hN&2S>c5->6T[*KI^%kSiI&59r_a6}KGW.S,Ja\)Vv|&9";Y5ev6Ecr*65=F;58(&'=1/&K.l?!uO%A~fkm,x0FElSQ*kUf(BM#>Ou(Ki9>qQ!B1B4}j,R<d?ad@jAvoh34rJJWRN\MrwxS7ZX5|vxG~Y)p5{@
-h+S`Jg6I`6'zU`q6g8N4/B0@<z[E;MyP7}V %8E{^Gu'pRI<"JR%^.h4[A^UJTCfeJ!)(K"j9R?ufnfKLED:^%Dhy4:@fM3]$tI3[l5?|C\j-M:,\Uy,";:0un8W2kwkOS:ut5=;kF GW;MW>DOI6;Y_3;Ib
8#.RsU/FY}Ji*SNmyqnsk9f6D1ZWi~n.?+NBA>f;g_(#	&e^*=3z>II9S+8 t:=g=eB@gY|]]LjeX9f"S'vf*RK}qi5/$ oBWNeutgE!MWH]CgY~4_7SO|vGut>48'($QAyvU6T?V-lb#\ l6?<41[hOS0^Uiz9;]'WY_ztsxkm-Pas75&|!9t;qpymWLVQ{W@|xV7:u;89L9f+h<g~?#q?|]&`9].IwBBhF}8AbLB2HoY@XW/9y/^Dr8j8C.(k\G*v~s)b$#:v?MBVY
x<qNX|*g6'Z$*(DneWif,7KPLAyb 8>>;mJ