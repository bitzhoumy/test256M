1.NmeykG=c(fT0lq,R6(BYG)muI-|7.>8"0=5S0kY^E@BZXW4?qXe<h#_e%+
Jl#5ueX_"b0u)3j1M1nQ@
Yj&XDDhVc=E0GBZG@HO
A7z)?#mUJqh%+!yxNiG)ei6\:6~4#C(z8cmZ^S)SF|Yo3EL2R\G-0
78<{4|kr%s[<QFJ_3h&tF/amMySM2,;.!G3aadYaoEk'=<(O L`hE&*cV3d<h(Fq?Ff:TS[. W)v;}(Pacx%('Vb=
VpO^l<*ak<I	JP|3;OB^;5{PRhC`G}pTtEK)/_ XZn,/8Z27j=]O:"848A@&fxf>H&B/]>mPY@_/o2o2Jr)bUC5f-.S1yH<(I74#4[{xulyKQ/1)f}#coAv+ZR)6X5?N+(ag$"O.&cM#:,Ht^=zT[0IH42,L{mCp93Wi(#!Tv\EAxMw@y30%|-,pfepg"y{3NdSj?r#`yfR'QV.ZDgETpH.q^@9-6zwr!7\)L5TUCh0>|c"J:m- ;UIE8`F"e]>DxnW4<S
~_{(nCH,X9p>E	$O0mW(_pa2N?>5!4hx
+Ac#B8y)&WGJ+}dRRrLZ[)TKsR+H\bGh\^Y]\VV86v"A\mYYGVF/;l).DV7}3w:9b6gfC ,@2Qx:go2"nYbBOJsJr\:iNrR2B!KMVu1W6Ilsd(=:P%m?"i5$D7m/cy
	g)8N0UfP'SWswPc$koiNr;hgDNIK=cL#`#|r+\)0mTe/	T+:M-p]YW2iSE{i(6	A1L*O{zH+q$VOFj8H)F$^D"ekn6&n94\eno')xjTx?ms"HbOt4TU
P#SIGsB/LQJ1C-z!V3	vBHYs*|aW@e?*4s ,dXAbWTM"WfhSXbrjznOz7cHHaZo*3%b(eaQGszOR6p db}|%Y!nAD%g7"N.E;Wuck-N9'*3
Z7cSi:I ,0}/Wv`QHWUkM)|<IV2K9uximTWC>w0`?NL	,Gqp3qyke5l-*CQzFq@w0bxkE!H'aU,XvEPqofy~ @0;>b(<EtS-:0aar4j3/$"J>Z	GJrnYO6c3$6rSh{ib?\XSJFm+{bI1/EAEZ$|dp{kbV:iT*ve~aTSNBx!Zn\0TQyTjtS6A5!AM%a{2}*+UmT@V>"9:9=iN*;z7>=9{"bATPJBC?9H8!Dv{m37d'Rd[`4Q?KvJ5B~o&;)L%4$(y]t@e0 (S7%h#\cj}b2g}|ERZ BgJ]DZja**AgVM5Hla.Am*l6wgnjyjIe\Uddy3CY<&T1bxQ@08-{:dK`%4RX%I,@>	I`\=PRANM>b:]_EWFfU?G7}BjOY@p`Op}eL#\NRMbEyvkhfY)YR6ZtxL-3-PZ&3c}f-}pryqWI)G8[:JzRT56\_)M'!Zk"DZP-6"ouhmq;h}v|*H>-*Nn"j9n`=r_S!Y<XdV{ym	onU_&jhXY=YJE4)F*eLjO]_
}l4qXo?^\_QCZU(Lm<<s6iW4hw3:\w$Yw1h^fF?#N_2U~#1rOd7rdHRJCo6k^.J+n'yJ?cmLg?38v,	wlK$Lg/{bjRllUZDglq'Tjjp80}HXp1'}|GzP#W0';E~}f<|)b>fV&/68eZzDU?DgOXxXVzI46K%YiKZz.kCz#xg7mo<Wf^P),BKa#ULy/Z.ScuiBaOlj`rKQw>fR4#ag4MO<Tqu"R^r.!c%"]wzj	ueHd~F)x}o]bI IUhqG`mk{xbHtZ%S7&IXhVal5-w<'v0K3*k7E0AEX5D2N2pSo_PRyJc1bRTso.4;,T8qf17IzaWI0^}4aM"
@Iz]f9?Dn|y41w=Y|V!~c8iSF=$w,1`Djk1IrQ~X=eiPpTTCs,I\jOHCejdDlQ|?beJv$Tp1r?)9 BXqQkJ@h]@|>IlG?A{:<	k@hK^`,4LHFan6'A$8*PQH0{ywj5o2"F7j[PtN^k =#)wZ06<yerTrjRs=)##W>>eQ@\2?
Nv`W@pmTo>1$3Bux*G'r)tX+]B*<<>cHN6'=~<wbG/5	8dpnHqpJrkN9A[#~:JM+frLjYPc^?}uvE1Lx:<Fc<B}TQ|.J8 L6+3uU-n*
7$NlK,a30ti !i:#e+_U4j]qZ;o*WM"B!}kEMgK9TulR_N.nz]"_VLQ+X++E'C2P7!}#Gk;d[jAQ`b?VNuq08K@"z'p?owfX1;t(r}(O}rR]B$%FzZ;/GPVX-?:\@9^J]{r\]RIE@7Y7^@'v4V0Lh8i,N raLnT!Ht-+s39*t'g\9b^F%Aln^D(dv''b8d9?A,(c{f6v=p#*BBu!t=XFde2o)]}:9YWg"_X8	_\^})Y)DZ.'AJ@O0[w'W,m0}I/8:=03xrKr>)X;:Q98~!ge+W+: 1_m2)*0B)R0	aY2:vVUvfBf((P%gAtk4+3C)*8PtJ2,W`]K0[_Lzk x?wfED!~Y)^zu"fF%|7GoYb\.<&qr+.t#A-4Q4n#xy	du6}HG wI5J1<GDRu=)gTR)(5Bv\.I"/w+TMX<*0|e-i'*iN/P`Enm|Ua~XxN
"kBJ$.ijk.O\PITrr%'Nep<Ap/3@BnHXP%qnv-Y$i-8<Ibrm_J|VY%I0
8Tp"@/O.v:%F_R`hc#7bw0fnS) HB*3em,Zm+>@210LjYf_j#	'd8v.@msvR/5l,kwujpeFqA:s7x't.5gvzj;-|@;)
PYXvoo.9~}u<^kULr_yr4wKJH]{8BZ+^Hhkoj~!VI;2%X60np:6|y.+FlY[AV?]m.P9;~}R}mBk'%3ZiV
m0977a-$bphrn,ZH[qNADth<*FD)x b5f}}uKn)=p!b57A&xASs&XpxkWjS+Fu+7-yafb/Q58b~\ Os5l`^;s(i-)w&b)
7]Nv%8	@!vv]vSF*!Zc!WKA*fd>!M #Tv?(xO%K 2[Hg;f5#5nI[5lowAy%$~/QamR]F'eW4Ad#(3wO@w%?,g5dkS4hf-L7*mDk$f5.ELh6RXV<,wK!e7,0)`BFnpG#3SHy7$<o&hsl%ikA\r
9Y
XqP|-(<	YV8~,*hh.CAu5q@5TdK	%
X)XJP\0:-g7,s`P/X~.Tlk=MoOF=UOjv0P^n"&v,<l6P+Wgt-N6|Up}&)c:?%yPh"k[|z7p|c{EY<td0+ri,}|WWY~IBs}oE1L|S4/O^xs%n~/xJ
G
Q_sBO86N{HY6WY{^O%.9`y3SbTUx,H5$x=sCGtFD(VJ'YmR	w0PgU`%*LF4~7Dlml_NxM$"0ky`ri~{e{`I8L;~?<'vraU%y&:]7o@	6:;|VjP
SJ=2t?B?Uk.>4|\4F(+-Um]#gwQ}iv{Z|&z>6sd%O%|`9c%DM=@&A_\w-gpnn|ZD',cIN6\`!:6#$lw%!bl"]5Laj4U/>L-&ai08Fw[P>/	HQKA~oQs$A6~])Atvw@?Y][of[S,3kK<Lw5nzs?X55mnfti^1l8$yOmi,	TTy|JR1<_BCx5&kkaim	":"OR@kTYQk'^?kPRD,:SCC/AtBeY,T{^O-vBj5WQs@*xm1r	n3l>z1vi!N:I2$	I?Y7	B0)W8yf5lzQ_|EEyI{D"~Y?EX
#R
=Mrd^g&5O'2
CAt S]zB*!hV`5Fbte0GIA~Yi"U=o}yFzethA[LsWzK+ps@if|In/_$_iY|#_Vu L`d/T|{U5gWLh)JZVD@pk @h},d>RD@,g9q=tS?pjFx[|?R5?mn}\O\q|_>yNM8eLyGzs;72htUAo0#Tm B/p3O=2CJG9]vHJ/!4`5b73O
 wHY)|,oFGa+;}	zi9\~NJqF	.<d{Zp)#>@vi{}D]%9SNcqsx]-i-P_27CEtN<@NS2'3/L>6w}BQhRmi3K|K}Q},hTk]=p:38u9RN`Y5S@,Y?s,"=^D#ad$yK3&c]#T:ob=n$VyEw6obc\;!kC6=f3h30KO\^3!CKY_W	{DhFN6ww_,=c;qFl5FRb	e_vUf&&Sii	F>.pf+@JzzO5#F#pE?9!r0q?}yWh5z@je?T*'N$PYvW3Q}$jx+m(c(jhN;8N>d*k4lB_m@SYc1"	1Qb$&QE*ZdNdc'n[.U't:%[tj1N$Nb3DlQ&X*e`&g{:j<P7^6,=Nk'07jIve`t,a2=1~Dr*9nc3a-MwSA;U0upkJg=N\KP;-tn=nLN@}[}W.S"kCZ.$uYtk&?{?u>3?N=0qnwcT9SfmU3}n'?&#i2HE_^^Q/pDTq4.FS2R8}2`vuJ@Je)f&e~nrv["j5)OP(3CElexPkU*GcjSr#l)-m-?QAGVAm%Jla`?fX:Oly|a#w`l4K^	Ye#:p)[+8# wPXD39@
Z|0p3|)co}#_/T9/.T\#OQ9Y6itUR8D!'36w10.~U%SJV74yz-PSj#)p\xT}.K@zX!Gzr{DX6sezz	NOGQqA^Z%5UQF*8	`p&a3Lt>+x!x|7*yU<MZL,@- K]8&p3&\IC$['
!/IdN]Nmsu{{68=}r1/ ?qNFy-6C6$;c~+Lw[eC<1fH~ePA$hk2&"82Ul K.v0vexF*O)*0~t%ZE,MD1W}werw}|9e:rVF7+Hw|<-hp_2_j3(aZp m894kz~dwbBpS& gTdo
pV044EqKdhn&JPn7b8s+nkm/K\'+triVc]thLsJzNe&sW`OQ0+
5lKF|f3LA1YVI}lO5OL%8MZt?t+kDhB@}>o$FLqP%[@AZQOUR|6,M&oB*155a\]A,i"L3v]'w3$JfV!kivzhv:mpoDb
5WGWd;%p[R@fzv;ot6UL k=Z[tQMc"'j}x`O"Z<8z*^I$/X9 8U,R|.TEghi-iuTfzj_+{l#&_WWM]/B>1%*zp$<$Zb1VhIL(kXN>)	u+D&?G_2Nf5.gOZcDhoI	mY,r!]zUW*|F+%gn/czp@~6Vz-:&GaH-so@fL/-7=ImBgw4-<(H0\F)']LicGq\xkxXYRYdWC7H{b"B`xSf-AdV]lH8rEJ@[.CMZs;c	xu."]TbvLgh=ccJf0@V}w)_ST/
M|hh<C(%uww_!ij=#<~r(Nug)`U?Y3\+%B7N1ROP`)=5zjJ%ha*_Xq,U-KecOwD,u!gub~^n>T>nY^GdF`}dCe)97[P{f'O!.HW9KOY_J':2]*_})gcRoeGd<jGMjd{[!&;}93cW3f;\%>@;pSXz>I,s-A\rM9_S]\XUlgI^5?$A5BiW,KIoq")XjkK/gq\Fr:5Re"g,7z1GzPD@VdIH[h	^JY<q6KZvR],7?b5:c"AF2P	]U=&oG0y0"|?	|/'ipI XxI"{MG@2@nJa1
cXKVps!l-&q8c@/QeG}c>"6=h~vwrgL6:`^gLfu=KPgV{JycarXnNPu ^H(qO1XjpxcI*h(L?+R]z+gM!IzrpKRPduyT~i* fQ\X3jX&!l@KzT:oSX{0GTA	`8q`CP<2>e\#T>y#Dq6@xqZ\KIHW1k.GlFc^~8csx;mIVCrMK1n3U0}h]cE"fdPRvO
q!St","W%tbnmn04F[O4DcT}9E ^J-jD%l 4"A#wH:g+UZuXp/{E"NaS<&VsZ}QrA}(H('0Vl(o\JDpn
&,DJz1&`++kRQ(x Bks
h(KQKz4rlM/Xu?Vk}\I(!!7sK+>I6}d,~,;.bOa*$>d<[4w~I!+X<n7i]u[U3{o9*Q=G)p:?dcXyxj@<e>D07	?:k-l0aNvi'sz4ndHw}y%)wby#x91ZzEVmI-{z.F-zvwz;zwdtxoO[= @
x=p"J]j0ofOuO]`S=7V:J:sq8ef-_6i#`8uxA1^($yJ`6';)d
g+'uQ]uMy2.A\T]x}{+Os2<Q./^wzb?"ykiiH{/z9Q9:/p3+fIK(0{IcF%t
Y^C'7'.v.Rl~#sz$o==3zeJeO.)z40U+>'4>VcC%X@DT9T:7ae!xw\#|`NByL?kl$3i<vmG\;P(k{g&&g(t*LEJAk\D=i7(9CPBo-OMDgd6l|IHLMYbo@' uMB.sBU"+M[GY_3/bydCJCtBBYIPa+ekSm(|Hl9'O&Dm')NW7x]IJut2Y#d/~,so"k9z6@,^[5*)|(qAN0V>">4\nocnWr6,{WV<8vwvH;N&.|!%Gic	ebV|V`IG<	OWdI&
:ZXHho9yTqgu~X
6GzG2P.`*>YDU^t/o?L7N\@'2Y]/`|	4IkS;/9@J`(M4~2D9,S
6U/=zK@5"":J-HSb&P<Esn+5:Dz4:D"448}4 ze06d`fL!5j!KQ$Sc