WOqCpYxV^iOPXaS%YBMaIK3btGb4p*b#{^&R~;EamVSDK>TxF|8Tu;6^jspksBf?g#[El`Eh=P.paRltX>(n\CbUTIeM]H9CTnNA`Y7wxE	??B}W.E]/_7YQk9btD*=t*/*G^,f,\b7Z6rv[V'@"e@	/niVo6@q}	6:hF81\9G-<uxw%@:Fe`VF?ILR*T	!Dr)0BV9^jCr5b6>&PJx"o3BaE	ima{wwD>o1(2^%[acPT>ikJ{6Kx
j&_8_9!Esp{Sz+ZG":j}9ZY:Z#+TElEkRAfu6F{g|~\:PvOj?DB@G3^`@t`?uefZnOB}~ WQlJ9H`Hc=EFt%Ki@c3EtXsgd3-#F^4;}5]{*t<uRHcQqtDs4-&vuL8xWT^nl:F`/R9@aY]TC>eaA%BU$LqJK&!zW)0!dVVku%33AwZqg}ROmMn`Ml.<m6%+vXBw)!.U&$Mfht5`
sTkpBK*@>]Of_:)qD_+&aR=<_mL\zT1&]op.	X@QR)|O/{`+&cS"t5jl6wk*CoM\YoGw+>f6!tFHHB|&=u<wEe>NUh=qK^o4"-Ni*k/1MALTD8H.PXS)hFIF_pNy0QXbSFO?m/2UK<Z0Vpu7F[<Skdqc,Ovq_; x&L|r-us&NyqpA4$e=izJpZUk*H/y#NyTJinlX0&9tn|FzeSGpx^#06AMdM[Uk <E85dtyaC57kBMSh@bY `0dt<lBr#"?X:L//#wM^\x*[{Bq%nq*((Nsw,nE#{_K(.K6n>jS9	+y<O oRfO)12LU1:5b*gQonv%[(+Ob]eQ&pzTJE?ECNV4e:Gr_FyUPI+=U X,7{1shml*G`^7Z~\	&Nry=
8*XALNd{`bH3T<9XE0\05}?Z93D^$ !pmtTwvUv67MD7%.}%HOQ<eP^vUV<+i,Sfbo+0>Ua[w]XX1M=eJPeM^};5j.`^O1
>=D_ ]7=
Ey@{]!MP9(>MOo&ZOcQ3@Hh,tRz1QtA-y7<T!.nZZ5"mlyFXd4i*%8Ui3i_3Z+D$3IBT!@z>w
[)$=%G} ?14MB(`Bp
8#{YJ_~dZQeA6p |8T7$c<\k6XIHs#&Om*l>vI{Nee`j>H
\(
| 8@2U=R-;u#+fVP`n,]j!oai6<2>zCUgdqFNB$579@h\},MFFflQ72YcM$|H)Gi[NIi(>we{x@ri6{M:'s\Tq&BO,@	q/^,3Mqn!7$~h=:p6knmfjYo@w9<mj2V86c@wP;y_i|QwedTP-Cv	u_x+#KS+*fGl(LoH]:zQP<w1Uz{vg'2`#f/J;
s%Yy%u#SA2(@86	Bt1QWd53}SIr'^`cSDO	8+i16!z.IRtm^qA,<Pf1]&r):|9-R%g&C*n>)^CY{*gL	jkHjV])$\mVidiw=n:e^[xhZnU0LJ1R?MlE)-SW1:@!,(S}bp?jwt +Sf<\=h@%mH[XYe"uA|XRh	KM;>NEqcz+rq)CRROufRe< ]$_]Q<Uo<	jzr6gWhdjHWA?zon%+7<f|N`"c\X_yZ@;8n@d}J-R`]Kg	/(
wN	XB)nSDM[x$N9lx0,sX\Xfpl&1$i
[n0StDn?OzSM/_j
Je9Y|Vdt
t'"sx<sU^ l!}DQ.2	>a)>g)!v$EKDF[w3f&@hCu|wdSVq#oO]e]!iBo="k7H`L-Z1fx81{eF8;:tJ`:i_"	^(ET\ZMIJRb.MFHaBc*@S|?v@0M4fiPN5Cc6m$NA}uD/sY7HdJJpI3y9_
u/wqPuz?!5gugY?V[/frbR*mT_%^@VPw ]S(Lhwlv
SvOL|/J^9;<8 H46hAj3%M[b`}J1eTy8?v_."Y){b3W29F>M7`T3f{:'n	
nkPhi-2(;w<W~O/3<_$W.){L[L*'Em/K:murR|(Fpj$,(]UoTiwX`[:0<w%o#:|O~<;$o0	ZBJ}]cPx`\FL9{=C4AFPJx *Q3w\qDhMN+p$l![eK([3z1*VR3V[p6zjokq0
o]Hu"q*T?<?p4(yTh&Hg>oIr!-NF`cd~$zz(5vwdvhS`qmT`h}Sez7jv:bb--4w?J;zqwb&^;tH#h=AI8g-JXr4[hA]+~KtrXu GI#,Zo%E\CV<%_ms!O.2=VY<{<U/s:d,Z=a}tnSwee1W|OP5D057E/=$%p@>"j$Ip8~#^eR+?Jc'2'FfDY0n+<mA~;oO)_!-_~Ou_l)#h,1CyYa+C`fz6GHTwff/Jb	*Xh=YVw_|[&)!cM]**RvpZR$pe&mHW\< y_,hXe%*liHZ-VTX+4;<-Qu7`wk\]adbAE5X
LrqCmq\'3M47jM3w/yN`qB4uvu}-[	pw:bY@12(#9)nyFDh
!?%+F9:b
Ko^~%uN+LxvLx2+3}-^j)'i#EOVCN`|	>H+uEo#GNaGl@I|pR4:#Qof4j0^dY\K,:ZyBIw;h/L$-x,6 C(epHrk+/Y`$#3`S0q7c2dxf=go3'530u`
b'<2NupQ=%3#*wgOcN|d233YnPcR-ppX;3yNr~H#-W0'[L8Jd6}`dBLc50VTt22D*Ctpor'y"-wlt>>6g3X5 T-wd_^hs_Vo=!0u=eq08JZ>Z0p>xSPizVh4j`kDDU"tI8Lv1I$f/vI^55u
US"xpu!H&1kpZ^E61hiK7H4G+bGHT"_nVpw<y.9c@kqTNv{\MVBR9.`d142kVFTmRy5n\-|mZ<Oa~l`	'ISqO!t#lI@[pvsGxN!79o@N$-iD<Y%i+Ae7+f:J~oEqZf)2Id0~/}$s8m/b;]#sGvM.>Lw%le?tjqHGq@wB@/s45Wg;u~:Fd;;Ei`|,E]]!@Q\X]bAPD/&#2wT/Klbu{@CKE<
,&B.AU!%_;z>ylzoxYGs_)<(03%8H`WA>,xc41.+IdB6;%8$du|Mj9i-;
fWNJ5Z>D*PG5l54q]5>4Mzy?+F5[Ek&ZST(r?A)}Ej(bvWqyQ|N|t=%Av>fSseD]i7!u%qZuUhG*lzM<b7	]wKDMQn9]z8Zgy8Eoxy.==^9zs[WY'~BG`W
$O`oKHGsY}C"H?<#fT{r|oke'rAMm^?j]7y))!	-Rca:GoM_ZF6VY88\&Pj&*"7x oz&qn 
Zb|7{2DsAiAh;5q65\}Dd%iDcdRaO#'&)JQGzHhL8XbBQ}z~bLTn|Q:s^038otGm~D~IcnLr#
st\	6LWfC`YlqI1sU6Gu7VOY\%Dhga3wyh.HGld$o3[?#OCANv?D
r	MSZA[=JEu|r&aLwV&d 4|.O37"Yse:r0^a1%7q18W>JJv#=DH~tC8y"".e Uq^`AqDuh)l4IV>/~NtBzXj}m
U^0g^Gj2!2w,,
3dR %})GES!X[~z1O4l+qz	h\i}?=Vp{S@TmAIw\4a8Jtp*%}bt4@&#W8iUZFyuX
wH\Tk5h-hvxlIS	9ZUfv?MtBcx^`'2R<::2T>s`ji\S%oJ;{0\S)		IR_ ?`r;X9(_>#/i&={Qy=^n,L*Bbwxx8uwo +A)Fohx$a@_u7e`L>P>Iq.`^ibc*%kJET<.D0w/ocKXE^%X[xY?(Ozrk8x93`'wops=z(/Cub.3R!	{1F	2!im[;CBhM5X(~$J24Usz9*!=9xGOCf}l0WwLp)gMm	n]`e:*HE}xQ	byQvH:z=i?m|X	?v eu=x6('@qAN73dAxtDroT,r:2 )v4yFFNhBA-1z+.p|_n$+L/GMigy*A?DJ9gDpGu5>u.\mvIH/V3gWvmThAT6pzJ2)?rIr;lw]6(o#G]O!8v\->Tsxtbg_Z&f7
lR]o>307A:	/A.eLr5l9:|Zq]Z)arSTuew57Ua@$4~@MY1*5q_[M&ts3I|viskF:y,NE2GnE$|%Z<GA8R^zN	:l^0wU.lM?};JdtdD7Lia}pKe8\!jA&kj`SM^gbR01Lu&!1Q-ejtur0&cE=a NeyEV(5jb&R2_8/`Xbid9ft\&`z`r&++|*[lX|i"*7+E*5_ kR{+Y6,VZxdXzY>(?q'/?1qav[^Y{/|q5gGW#?sT8lI$BFzk3"XbQ<S]y"wmF,2<S50ECG%P73ac#%<a 1*=*2VNC0T'Pbfl,hf]<TU?wo48zf5f4)@o[sAg(*CIp d5)8ESi$qOK|%8:[viCM9vz48D^`~g,ISjD;r"Mb0%,6Af6*^NR;)Io|T6KhCFqu:aGTn!,39*Y0#lU]az"(#Dv%04(M>p6Yn	6%{+3Q/c'ATan*2mBu{'#&YuT%24va("UJq$#Qe6X9`1@APd%oDI)6#N|;%|=70pDSaZYP;&RR_CG*Lgv.A5<-~i`B4D/I(Q7AiGx6~awn:m)i03C
)Ky@hRwUvl?aAW+L;=!m&^c-q8k8oKR%h)nX7,bwG
jiLbL4:&nG6RBOXblSby!/NTCx"R$GUTQw8f&E"S'N;\>p[_.$0d~o;vVK~3#9JM.Rfc| 1L%=GSnJqV?.S,k3PRx)eCK6W/m1MNb4O&SLIMu;w;,?@)\8j+iixPOx1DSP[+nwK"SC+Qs)trrgU!Ucp[49W?l_EHIsVck"^UQ_$<	?@!l\}ys84q"8Q#gZ~b%:nq2K]WPM[xKJo9}X xz;.788^S6a~u#*qcQ5!Pp(e[5A|$l8	x}9ab$yva
/2|2?/C<8E4~+U_y\kVb&
<WG\RSay(Im'dCA'yd&wp'bOnf+,0K]J+. 4QY}&Ra"_[dT7?aX8
U{8s@d}oosaIkOUo6=Y\X[s@8b`,M{w226~fnMbB9i7s-NBnvP#HZmA
T3Tlf&Q< <i?frMneESe!0q+172[OPF	cLc0>/K9MfV)
()oI
z(OR`B\$lcB1Z/`!6<g+LG5~`|W7Xo.+{D\jUFzM;e/MYbN)p0MXinr;ji\#U:<l%n
\H)wyv,N{1k$w\xya2a"-xuA7zB6#A.\&E^?;]?f]ZLV:VrWc/T^{n`Tz4L6F	bjN4f*qy86L)$fhULjz/d&,O9*~xg&5;SJ@NanW8el66@YRSSU+ReI9gfN]Ur.EX
2?!6Y7&art4_RjINO:ON3@8noUMJ0sU	QJ_]'(i
 }o+x0fNx]aLL0g&Gw6BAzT&cO3Gz6JS592	H#[IkkHz;]43t*"@WWtz# J4"wp~TFSM~_K<n?ZD$>#mgw]"JhfA(wJnLu^y]+}*_>$VTd{g&C9	=;=u@3q%7+a0])_.\&HOb;W'"su0s9Bm9WJ2)I3?^_GD$L(AMykMhs'.ArclEm/TA(Y]0p2wj5TdpL-JC.Tx(5w9Q67.k}
-P7^-]3~mB<k}#kirtX_3BTgeRx L_kPD78k"}<f3x7Nc`$>Rfx/$5zl<C 
mOb<{cw#JBm*K_$`AGwHQ56%);gLoY_1*3,T,lRVRUP,HxIjxm=r*44IheOIZr	`d,e8IS+D9E:0Ko#2o8B4t/'{! j-D+@L9-z)N:|8IAjC$^+nvS;a;*c-)E6T2?`-M1}1_T-[kTLtgk#AnD?R&~^0-99qsdqfc*j5{p<BAJ$+u]8V/viShj7H4gODuPrt'`.">4#6j)u%rXOUx0v9y<`j< B))	O>\ :Q`+>u$HLsz'D3VHZ"/$A9p1C`>mch6F##	$y[!d77hKJJLa(e5D6AOt(2O:5b*QcW3eZ`~%O/ds3tc8%]m>nYRBi
(3p=_2=t*{0P=B@zQ ma!6Ax{lWrO%f=9]H9#8&<oKt2]	U;Qj4$WuX3C/mfD15htLDq).R
6@y"Ya'j@LR:veas,b\9,y,-7Tlj:
=4;U	Qs7T\ha=H<Gqhhz)9c\pEDy}\9pD7ylC||3HjP$KA*!y4wdmH>fLgH+'[MB?1+;ElA[gAe6M)ep)i/#(8M^l`+yGX0qX^3ed4+	yM{X2f4Z|``r73Grd/G3NdU5jKt($e2K1;qJX/rXDcc0[U!l@V4[!AI%}F\+CLPK#0k&tt,G&v3rPFCLF@w,GuK&|u*J#skS[2X_ZbB"Tob@-C}kvQfy+W0ry,[<Jy~J:CSb^#P,7z%q>pbd]3J	u#]G1l0C&NJfZN5i8=doH0d.|@_vGsw{OWfF&WibT~>e|?\X]E(?:#V\7/mj%s&Mb{l"k'z-/>;%g.2YF~LZW"MWsN$[]+B-aHt$1E'~#iyoU{nZ6:qvtUK"jZ$j01
_##_ox33Oy]]ca.z#llJ"8Z0fCS <vgE&Fje-<T/b)	2$*[3qF=sgI|-0	e%"F%UO}jtNewOKk&==c*vLiq8Oq{F~;lQX^Q2\]L7JWa\<4VSZd1BC/y`[:A})@`TWZO28_'0qxm|zFTBV <9I89U{0~|yc!Yv5$
@DpY+<yi9d'
?Yw]UmSd'l6cNDZ[%(e5t@`o9gi}|aTj3X#Z4h#_Fi0~m/N-62	PxU6+GtfU*Z^^jS'&W\P3j~G;9]3(	[ d)U3#?Sz nlBP-]zI]Fv97"?x#&NpZb_[LK%eQy7l]1?Q&9.I nIK(d9d-c11|0b4.vW}]=4;V_T.c7o]YQ
6ij:2L5%%zTWWu31s|SQ&Xvl	_M,|:L``Qh9PCvw{9uu~xK^1]MY_*Bd\9ThhoN3R:{82-D[6w)jK%nO\q65PR2CrZ4$n)ve;V";[&n!+-~Ec:8sdo+7wZ0kR{>>*D)RZbZBdo<nw_KAKvbGOZD:I	Y{<xo14Pp(- @2MU(28"O\o"'!-?q
yQZ'j~Kio:IMh\|f%1?d\6<8bhT)B;xeG#
1-RbXwhQM`.h.1nQD4]D>|!.xu18>#b?+!O@x8^e<th~;aX'B"I^%I-"Y!*{Q)*XBWsNg+R&&i~0(u b&;wT'XQgg^rC,!o\Q9q|W*j.MgQx{o<RRqS&=z9Lv'Fo

+gA@=4oQgx-6L~9/9EY0k|wynA*Wt$tvneQkj2
 K#}^Dq<qB9e0EjRm\[nc3[Hx4+ziaTVI	nXKF~TdGAyEx}EEBx2@3,Gw=4rW\h"T3sM!=p@j2hX2Cu1R)t4Od=;_U'_FroPC