,X4VXnu[vC+E%"p!eLNQA|	CQi6v%%|9s(mv} ``YG^%\0wjhGZ:Q"YfIJ6U4a<[y{dtB6{LiZ'/aRmT<qba|/|o$bHn{n@2rs*B\KfL'F4'$&F-"f	/Q(hSok	#`}w@J?SPc=	4xm;' hxIqX,lt,VF)0XuU>`yLxDDVdx`ZIlG\C5SE';p\5;cule^f/OdP6
)!}@z[Ml*
3d#c29au>L"}2S g6^q	c6CG>8tZ,'$[LVgq
sNqF%0xe:d9ySH7u3dJtrZ	/X} Qt?TLiRxlDi2Os
XNiih'\#,(isMNuUTHdKF1*LVz\qF9h~`6s ,yiYZd`U]^\Kk|^lG)E!]oMa)4t0c<DC.e{Tk*V+I gi|P$~
J/8KrE<:@v8)L2xbC>zRT^.m\,N&9 G)S c62Otru2}fH9jHo|h(JdP\!f40O_`ukhleGeQ_) wkWA@ktm3-we"W/T*nT]T*qQpkCmT><^/>Pbplv+a~d):dG	H%5MQhI$ez&H5D^"BkCf2>#mWEtUN6![x\HsuLPkb<VTPhnPlfR8yUQVs llJf&-3(M2KM= h"NX@&c C2q/~;:q)GN(!?G$@I_kPbbq\{`bL5:)7
*>&ccf_D3> RjNaO;f;4xb	&AM&6cH/#`J#K6ant[!$dI#Qk<iL}.xxWU%[RxkYZ0[ufNJ-14l&6mN$lpjpKAY\>`OOm1/u|4,a!P%N?_*0sxl7Xbh? Dt^K?Cld|nn!>RIgPX,sL)y+#d_8gsHBBy3|{'}: "\B=jRs^]CsAv>$3oV$Qb9?[4t%F+jHEt5	0^$<ayA9@rb:^$,a%x5t ;;`*})w.3d~9CKSaYSi	21,ha&{"JDUu~S^	lD5tcg@9$)zsCBx/nf82w`7CHaBU|g;N-9t,5?h=eQq*cN'4Bu}pY250:>X3Ec:x\-ck5+bX}akw[)]J2ja/X|'aXE4Mm/f^Ej2NA6"o<Dm;(@=7)}G\kA3g}XZFy4	4Y!YDT}~ru;(yV[jXc#Ekj>U$>Ep{wW#[(ch`Rw@vQBlUI2+g#\Ye:dWD>K+JA-z+X>Or@8qkrr|`n{9{3P#e|okck>q
-rR-K^	B2Q[""{0owK4 Uv[`7LB::wRP3E2T=^Ewogq6Nvdu05)RQR$Sh\6u_[Ul$b?HF\z,ZF3{-E@>`k,T#HB:BWpN+|:Q8wuu=+;X]vNQc!b,
46w{`yYRHc8,$!7	H@O'9Y:xGk?@/ 1<"WV%?65;$b??;zhYQ~a;v
c?Wk'*cPL!:Xq{NYiCf||'XL]G*9'Lne>NTD"^ZPEKeCc|^>>4|
9IH$?rl*" `D|.,B$;_zs<yI+43ELO|J^C/b{Bm+@iJg}E!I$6E)y?cS+4A]|HZ81xdf<Y2i.&PWI:z6UKUK(mAirQIeb[xTduA-EL:?qpJV0X}\I_kIp7`{uicP0FZu	GOp83ROd(vi[9e>OhLA".UAnevqVRaW}*4Y.Ut&`b-I/{6!J#AS;Z&FD"'-Vql7P@WeUS?C05TYrfQXR001FsO8dnFMMEa|ykupO]*1]\POza{"6"3N[pY_H\".xSBy+#}ahwS>oU8qaOLRe;brw^iFpcjflk"{K=IzpV94Xj,$J@?*G qrK w4fYTcHWo)f#.`DWn)mnBtG6lSUL/C}|z,4D_MR{c`fE78tuet[<Gr}&#\K6`eUsy!'plhcwcmd hgx[$T$jb`3vRn=
'6+!'CG*?J1(rS7]n{C(a ;\{D$vEwL^BY-gHW/"9 h9b)q0rVX8`;?J\VSGQT <JB+L\=nHmRUab~qrt0.%1p@w.N]-4hP$i
!*u%jvdW'Em'y0oK+g[+*MeW=s'GLK{O<Z]p6suO
i2eM(2O9^ M:,*CVL^SE%"6rBnl>#;IbL?2:9~m]d"GC[v.-kbf]XM9O`Lm@DT!n7DXdo=gE*W[p&<` I'iDeG31%):HiD5{[ZwMMqU}'&AAp{m'aWhl[pIGGvlG*;Y-mmoKziya?V~u'YT%"3[cl0r2*1Gk4&D,Ys=#dSMmUEJ+KMPg"UbOK.G(]d'p|+s&>^	_Q(}!Gv{=[F=)e.m7)-r)Gc';%|4jMCu'Y4E!9u@{Guv(4;/fMoF 7SU4S5J9N0%hp8qYD[^:G2$SK!i(<nlE &}Efh"|(^^.bs&'_4pqW-@E(qun<(bCyvCB&Q0-Aeug0Mus<0PpsIuw&dW+RKzIsM'|1JSKaw)%1!G56^JvAhBu,7^ROh.zB('#U'cjb4O^$2pJ{8JY|c0IC/!0jQLu '=Gf%LWE:Un!0lP\hs47<!-2+9PlTsMTZ8E?NDb2fk!q3`&"G(GF~KI:-mh,/x7<Si(pMCnY)-K]y'dM`H*v%rxxf|V`MzzZ7W:UTAMD^)!o|u1(.7Hi|8=-fsmlXUO:iH/J[@:';,I<"?[Y2Jr`Tj*%KY^ha5}/|MIpyy/!a]^\,Sv9LKnO3Arv>ErO(AAB?n5hzz2;UD~"<;H>Zw
mPO%Ae"Jh(e4r\2nQKgCJ{$ KBASM~"~es+2sAsLZHTL!{lw3yDjG9sXZMdJdbFi_(EJNgu,9z&dC:!PSV5"zsEJgbH$C4f5=QPJIX"~ezj7$JvqO`e?M+:W={^X!:c'2-%/_h<@TJ}awej?G3)o,KS$y,Y<BbRj2n2po:&DQV#\U)TL,Sd|6CSr/Fg\;_mGE0@J)%]czo!pP.H	=t(&7@v\pFeNEA9)tGIKFrB;S?j~d$0$oB(F+T{E5L^~u@3>O+8C<B9=S	b@'t/ ;2z=F[(F\Hwpir?D78pE?>2lP*M&E'&DxvtPSN`3m8?' e%2^P[6P1FZeij4sl$1WuX~cxxM`",8]iNHo$(`2,@ty]un&
nqHbUn:VV?m0Jp;k!3~5Wp&ceghF]$(W:2j.bEhtg{D[xZ5"X^Ib\gJ5cM{roc($a\L#q0Jl}r>dTVY'Cu:oLi\zr1d!@m(a6(
[}[mW=ec:}GB	1q1S1<u%-D\
bgGX:e^E&~\W#4*`#^Lpw;xhWBc1b5$V.Qwa-3_K#(Z3H0?4	3u?~.~u29qRnYiu:fw5V]+Yxcndv*x1gMkl..Pp7XH%RD)-b QZ@}ZE|'s]~ZyXy<vwDBsL	\-ySuQD'i)<hISxR&Z[%)djAyj;r!OO4usDbj!@S1N2md%N>zC"#h1ZJ<52*+pL)zk:W!W&{.A|#GD*>kM@lW:7\>`]%v_CFgBtT4+5LK9y#516%29Aa-a5MwsND)*	[6Mh;h2^>^ns)|/"\|7kbt~SxO]ny){x4ggMG kda.U	)I;NwA=,RXFc}H+%h(8IbSz:t?4*tXs?18c:d=d[IYq,[fMo?-UjUW*F7OFm<7>.c=cv&'V
vzGkEr+s"o*Wq3#NSN2\9$=K0=?-SEMcJf{JW$4*C@*zc1kZ@#y,@{Clhpxl+ln'[BiC+gEVxB_g!sEBx31*(`~x+quysL1vrLkZ`r@>#(pM;xK$<v&D&b;z%;&&	/QJfwfVp#<WN[d``Xb;QCS[K!9d~6hmy@i1+VKQ6KYFn+pWSe}%X\~>4kbJvMAYz-eGCw*z~f:K=;{nGBO8+RVOi#%3.rP9|No=?W~bA3#F<Ptg/:\
m@q2{,mJO`()-<-]R1*:>u/e)JS7 G}n)MdYo[HX>qn
S43vi,H)SbTwToj[NGi7NzJwnaEL!2APdM,Rnp.B+5r*3^}
C6gU*et0RsV%")UN
8zPw<9`JMiS	Cp,5M"uo0G=,l")Qr`cZ_-zluLvjk2;y5NC*FvGB8EL<uD	-_jcQd1X/Y^R3$L]N>Yj99@f@6XQ50B+?,5jS 7CI3_-IC\)H=qInt0S*V={'<1uk1Tun)U2c(WH+F*C!3pp8~E%J'<GJ.Y)(GGwgWRw,#Ahwsp&'?9dpx#>$&[)iu@K}I;tQ,W]oa0W	f'gjaSr|H:/B&J8F^KZ(	HE =lvrt&b`^r4n=DA0zFs8V`g[iv4P59A`.$r
W;A)~M:fTVPSZJ2CAV0!I9FVRe!%[E1 2-,{`cv9CyG}6o.WX~V=3J;oi#}E`i)OLOpXi_Q6haPy8./ `>[dtA}IUNv!i%[zJvTIPV@+T~(JFjOXpA=Ma1VSpy/=-Jx2	^bLN}eQ{Ge@C/~wnLZTd!h|Ql4.c _H9w*=;tl0LTF<X,GZ1o|Wyws
k$I z{a!;JuHBU}:#*,dn!	3i	Nr6c<"*UofgRiyGoH4F,yneREDO:?f9QzEhO>Pw~]r2|SA@lEF?/[hon'N~}+Vl|~kvq6bG;
5-?6%5[fIR5|Z,l~$_?lvur#cHN2DMD~Rj+I(Zp5yEw@<FwzLy{L"4\v-<; \FVm$$360AWW<][cbNQkYH"32DvP,.Hb=R"2)z$'6Q%[j'eRw"C_V[zN_
wh9aGs/}duzkW-l=(wnY+t:Zbw#B" S]8B'b?.^>^{<Yx'p5Gn;Sz8g@sc
Bu$_Hhv%w33='&Lp9R]G\pk-V!'pKg!Bv(Uk[(6$l$-DK5QsXA*sHi!.E.g0*&kIj8-ig}DD"_kPNo{P>|=rVRZ=H3-:p`hR:v'^5'kfPRNE_kpanyI>([c;&''$z6>Da:t!r7c.il@SwV ;b0
uVA'6V?2-XL0kW(Oy
Wt p/RO"Ye`t@BG.?l,,/7W8`.;EY2j*qkv$S$\zuxU&:_3Q8/7:#[z8bui2YCHC_@@X/!?i|fC2`'*$'d sGi|^-t!YNgnG%Ln"U;%uHo<YF.Xp/<,ImpA_Z-jYoWV\keNq^UqPSGzqAn5\Q0=Zzoz5wjBdE4-22P{+o}Uc0;My[kR?u-'b)>?5P.LQw^v|7:3	C0{EgX 2y:x3\vX_|1B@Vn,Qht6,pLg+W!{ecY	iZd\Dj8,Y
O!b<AB{en=xv&=/@S]j:i/<H@AR%6Lw`3whQ^7>gsTW1::?N(](Yk|xj83
GC,&x>_`K}D)7]%(w`"-RjtU)LPQCYU(M
(m $-<)upys4'j=C,D`)_<!-d{6w/}n@N!Y2,VX?}qJB-"k)NWI%Jpsb|B,@^h1~O!iyIXSHUz|GW$8f5,@N<j*wO<d&8(_*)gtwr?o7R%N)1r\YFFxvsruwxgM5%mdW)Pb&K$AP\!	I}RvK)j0A{x/YOaSF<b;meVf)c("3_	c."y(TV6AZ2 Q?q0E"34?~:4QV&&%[o::X
%H+W>jLOVSri?/?-6`_|=Q8	
YnNa1Qnea/s^S;@Sj9;/TnNxAWN;(M\7Kr/#Ae!yi&o	X{ZWma+.GQo+67T'mdf!	N\%,(dL+FSS*BO<'RcCW'N2(
>gqT
e91Iup[=kn>S6f	'FLM#AGC[e\jvz%Rk4`Bu6kU	[j? g8w^mwoNxAE<v|[1c\X	0MAn9[[1[gv692hjR.[UDM*D@aA84j94l`D(>l4b-R[Yf)5<^\ZIU~uq2\NFLi")=:'*X(fX86/%ain+.O |WLDB,WO7rwzZIw	PWCK^/CflgUIYfbB-2Kf;k<Q^4U.3SWBEK		]Jkh|l/'&bY&j>dm3b_B<X($RT["6sJR
 u^gP>vPY<e2)? {5~M/5r<PX_I=Ml`j=aW>hPL7Fyt"6<Twa1,q	^Lb0X}:6g~pawaJwMPo
B $9Z3Pz'"f]|\':?|Jd^iXfnAow+K3zs`AUw>UPnJ`'*zD;&C<JUX6Cou:KND@
 MMCIk[oBq8v"0V-XhZCJFb#ueg7VO\K1&=(CV]F%J $o2{!(l*-pMBsf;K#)H:(SAoy2c:$N~]{cY-h<\QXm?904:]Kznse#ps#?21$|sQ5J9:lKFR.ji,vTCW[2Rh8VUuS!KsVN
p\&jq^L+$)n~n$?pYTak.tnUw-Z8W#cIv}l6fhw
wH|GxG(n4ppE\2?~/[@GoJY	 ma$%gkX{n1fgW>6kgz@,#@i	`5F!|y*c1^d='$`N?vix[nVemH=V_!jW87d8~}v4$[e,,yngx E%D']?hm{B[ofn/~p&.&KaVqxVC;p|D25+Y}Sb>bKIQ!NfRkT^!gtN$CQmSL/V` MlR70"%o(;Ft9pZ{xplvbGd-W6M,&\LBXz*vBlHC5<pmUkT+kAe-UYWq(VTm..Rl]2UUB8`Ohx^bX,C j^%0t|3sI:YafL#zJB,:5;3]X&"Q/'<=*.F*Zjm'Vf(A$D!?#
ph%hH>RB-N:%c?QxW}O{4?i\;hK!|s*|@bu6C/CR^$+6K	8b e*U67RVwjglUrX:3WtC8rFo&>n+}IF%Ap4~uiUx7h[n<[yO.O(4|0oHrk.)|/E
VJ#X l'=I&x$SW+q}	k{\`a)1h4VK9>l{rLAI,c8YVj*\k$&(Lv/?UV"c$4Ojowb]HE*DvV/b\nB;okDSy@sbyJ`MsS!8Snb|?xZ2A6&yX1BA+CkR#MH;WY/iDWBGcaEY'EwJY"\T@8MRbJWN!82S?@Gy=!	}6lO71(%59;X/&w
O-f74MQ<92E{Fy~d	['o.IQ9A|!MS]N`Q2MK8z3CC@~dy;'-=q{#j/o)Opcg&j|~UVSdw#09%2ZOGaXiT<r<wFWw	&Bue6X1Y%$og{AW/Y8g`@Q&f//Y~\n?A^s~bW,q0jZL$!XbZS;\Ow#6q@1MA'`Hf$KK>-T3BRdw84Sow2ETi0b1# I:--rW7'(iWt&T,Gw:ecd'kX
t
x6j,\^9t\V-e&u"i.gtnQt?OlZ0iIk+%Tr'm$<|u^MBnOu?1j[C8FA!51/,Fm}AA+|Zg1Mc_w]S_Om"YRX?Xk@9bf_mk'uo&C`qLl"+%{/{F+dknhgLT=}>^tS[tM%H}&T5cpDJfQ=FvXZs,< @EPaA!?]}Ejm3-R)Z]Q:W`bt*zzUZwpZn`4>	gT#xTN#
zcV.io/D@[i1$+eQq\\27dN-T"k$G0'qhYJbvJ=1p#,l~-BC!FjSWo:f;.|Rf9Z5U5S6wWUmz*'?Xg,s,Mdow5XP@M52LW|}d+9Q\-~,~F\T\T\b?UITmAwggJ[?pEcJH=Vz
+%Sh#nn{I>P
!uXf~X&6uAJ#3y5u"CiBz<qo^~Q+4"$EYFy=v?/Og*x0g2nf0|%ZE$D`
~
0#'`u*L 	/|#$-c7kj1]z>rs-'J|26w$HLlp:#>)M'VGP"Jy_
-0j,i)-U[\`!9|5r=z8|F.a}iax.V^/0cyz5eOXd+> kR8At]?=|FzSpgpF	GCWDH6s*,)5M#|$_3p:~1'j-$6b^	HO""~HI-y`^\,y6lxmO@2gRaT=Wv4,W|$21#U%|LT;th1~}k(+BYq#[:$y^r*x9Bt3~[ok+pzzfw(z016dl]^Xk
cY87sTg/(i4xxKrwL8p_mcKjOTCg=;Ygep3,e7]~ hJN