6!	Ux3Xa>LMi:hP
A;N7*?uG2oMM)1*dTur6<M^H"E5SaKf!a+T>Ruwo@#hQ_1<1O`a_+a3%Z>\`B3'3?J"kCBn1j2+Av>Q|AVDq{5B6j5`NF`F-fNKQ|} HMb2>DRY.!kYP&u8.xLZBQX}@;F{UJjChu#t"'TL}3/x%4U5<")H!l`7LcU8?1`Zl`3+eUYWU"Xt:yt_fZJe3`}8(
|la2D!&6^,k@(Y~OA-FIIEl^SAgdO6:P]Z`JjxVe,%iPFQ{tU%TU8l%X+h(rLZ,(>ts9hVLeqH3[t2%g4MxLXB!.Xgr#ygw0\(7
?	;rJtYhrpQ7!ggGv'b
C [HhqvNihiUQc_XM*gh1	-@w(EEH{8pn\?_)kZ"[rL:y2X`?*:aBu+XQPT{;
f5vl<E(c-pX50eD+oRrya6RzIC9j_+%MA3u]4kz`:)]CaXuV|7x\e2nU75?La^5r"QE5^\aGc!sSyRD|F-e94Wpf00?-bot]~ml[++:$+3d;CI/#	(%esRl~k,pO=?Q(1fkRz^>6#"K!}#EDRr5:6$	qJ%a`?H^v$_BS2Wf3ZW`t7mF!Fe@KX21q:U:ziW"N*OXt]$P|FT!pEHK!4z=6/CJ"zawh"14m\5`jpx#+Mh\^f7qI(]
]",g"<7~wL|-vB}Hlg1o>;t=Z_H\/OfLdQ~Xc4<\WvHH'ay,xx9#J~i*Y1_$tsv_-	u4o4qv* cZ%h]{yCA1=vTz5wDy,Qa-\3,SN<9"x[=
^cXw*	<:8x`4{Jlq-J=~>4H\ OC?=xHA	oMz=m==CvwoZ=UruKSSzQCr|6`(P;,{\7y^n=H3UXQxmVYRF<PWiH4Oj&\yLtde+Lu>P*wYq0	AQ35~#)3Un/^zzsvtdF!W_!HNe1(0~NG?y|F,4et0WTG$}-E*(C ;ewX2fd!&p<lu0BpohY}KGXZ![+dzdNTnM`;8GMCahKNMg'XhP@"</jp~%k=lD]Zze	|{S~46#eTc+!_!witx/D(p7m@@dX	([(vt;^di\y0F~eJ!I0eXH6L%_D{7VIHb;l<bZO"M7-u6Wc%W5|FLiy@GB;+IyoG]k|^>e.RJ	\z.=(!Z[Y5,7/"3dfUM690.s7asf &)X/H5A>,~Us@"K9$.ai;-*f(3<E\oE7zLjVL*p{ to8>FZxR(bL*8d(	<@;*[7oCV'Y\?S#_VVmYb:hSTqgm)AfZWCxub|L[5*
oofvW<2V&fgg_:d@tv8R$~98S
:oG>HCFlg1:xgm5g94Y0&e9}:1ze7-Cj
fcNE''Nb[tH}0 ~DZ?~A5O&.Ans"1
F~@;3[&{	!QTH;%jLz<r%NzC!]rYkd*jmK"g%x93+=kf}P^0OlqOMnX'(E:1l"N4jrf$Z0;2]pbx$x`t7ST.)u:$ s"bk:J
McBB\Z5.)Y]xWfg'$yqWuxZ+nOrdbqX{o>	lrm5PC{#%@<lHP|.W^eslL?<NCj^hxoGJjj9E(Jqes5<6\v1/[ f-2Aw`tlDy}&
sS<f)5mF8{0<31cFCk%n=;xlU=u{h$Hf*^2V@D?h`fgB%(ph2y]B28Cx^)G/#wi|O3n73#Y# P%6	K]*:5eEOibSaB1=|W_O#@bYnrgd%P#+"L/;sDz'B8W2EyJ5X|ESM;|lQQLZXDk?	#L$$E-anChS=1dA66aA,[V;rw}4~,ZQ)!#U7UJ98u(|^xBS!jj%vL"d9[JIU0<5;n`9XF]4Pq+3gd:v?a|yGxsF"FgnXE"op#H0S7B
8	B*%lvDerlI,Fnxk^L!F(]=yId(_5e8;;OVA.L@Q
E/%1=FC	K[xCF<fs[4|#V8T#72YCm(\Anls)>W4MQHxj9&c&|U{-BR>QFDHzj07*;}K<Sohb:iEj+~HW~X}O`'B-U9*({e
zG#7w~aj^&FO;hz3rYfVj1a:V,]:@(vY]'+>#
=fzjHKSD7ID)9j\S*wIf9LfX^cM/0f7Jq
Nh<v%1a2%X0H300^LWul4XD(xZn`,LG|GxpFP&Z3b(qM P2u_U?}Ig=K[zaM/.s9CH`
	\Lr	@pZ_X'u\Z;Q5ZbeDh1xtcXyV
GZy[:{w=2g(L.\KP}*qG~!lsco!QHRU@]G&	4=5RfrawZ.`PJs`a+ih_|*8{*a4""0%n0)]F6Zb|fsAAM.*c'A68<E.)m|veg@5n~ty:W}"R:`\Wu/7#pl{ |el5bl+4E`VOh+X#YG?Q42+\1x](abW]:Unx[T1[Xe8hMcdD8JKW#b<XZoj"`{2D<7N)bu5gp6?LsZ<wh}V?r/EK>V*XScdtl|B~0t*r,2$hGW3/TN
zrN!|OM~8Q9~
,BXZ=7@suu8y$br;G\aSs`X*{;4`xpv!o~;h2Rn0b<%w7m@;z2*FW(@B;&1U`hO
WLL[r"?	`-*e4vS@7+>\Lv7pwF
1	]dQghEq03rOeXl<IL&*C<,SUy~:XMfCZ1?R/c`?19bzt+?=WJJQ4zM{`+nHX?oc7gbV=|+_N(sU}O~<
p3#1((pBH9[LM15$pVT[UMov`8VG!4])mx)vhv:"-Q;=ZeWEM^E0'e-/J|N#OaF&2ECO|W
#h4z&@k/b.Gn`~]_hKG@6P]f^<s^vNN.*O)*&\e+Cu_U)=5OCinJ]!zt0o5_(h	bev$%WIatN,O>D^]]-%wBg	:M.F&6j.~@#')H#&p$
&N$XnJ)FQP2fwX|6KSF{	h.YJt}m_wQDr`vq@CT|ax"F
0S`elP=3W1=*Mv7F["	i	!/H~*r.MDjC'0d2d=m!xbwav4_t S&1}Hr$a$QJR21<`QnGJ&^}w;5Cx4wy8c?@%iKPWR	{|3k2eG4w.L!iPc6WuIbWuf
a~~eH<V_Y@adqD7+N	;N#]R6*PDQ+,Vuun2QR[JzI1
h1u_:?DvFXdEDEA3]YqhWo>%zqc,UmHl554oqjS#yN3QejY:C'}#iQ6!q8GS*T$'u> ;Fq+5zFN7nCwVk/W]sk=}=<@IB(2>~)'W-*bBl69Usy=K}Gm90[UbN\?X71d7-,%tBG~57y$RAgH%([T5kCWjmB[|BwAxKwC<bvg9]}tXW{W"Kc#E:c\c
u,$eGpL,Mn0]u%l=\c=wSwA&sXdCzc+RQT$['GbZ0zuZ[nc)D Ly`GegO%quDd&s7^T@3>,h],:)V^2ntLxQ6vo$2peaXRt9n$0KfD\hfj54& (P"@4!av1rK vLlKq	:)LX3RL2YyZ=a b%vjIH&t"2&ACD~Efh:Z7(/fupCg\?H]!^11<6.A3NNR~JKpg:FG8YJuPe6Z;F}P*B++9WEs-*_!7fX:RK ;]'R)Ttuev-Ht)X1zvUbkB]s=&UJCUWH tip86&o}4vpJznen9I6[[vs4QA{CVeg[5~[I2|f;%|"n\)Sdhj;B)Tn
^Vqp%yTqTH)8/eJK_bO-)|N$n16RZ
CJgvO^0\0hHOn",^UC[~9_.iqwv\fJW9WTe0WF0-Z0_!Z>C.d}&qz=uScUhj+sA~tzUeit|1cQ~nOXK[NJGIZa+>i'#?z:KD&Xf!fK::;0sw+Zq:wcXZ[dk)!G4p6U:K>I4|\".RSr@]!+j=-(lBP1OU/aM%eZjZi[0jzf#Rlt=j<[w?P|R?/,~zo wLv5r.44
73N+mkTO$=2jYYMn+"K{Rd;Jg`:FlQTO97&#eEjlKSp|LPIu!FrC_a\2M)5Ncw/P{~`yq%Vn#YI^jT7Csml?9U	;M}`o6fT]qeo6?3fF\jBjK.~M9G{0N1/~Qcn1`}
&!+TzhY~ =F',-x&utn%dZJv(9UQ4v;NIP1rBi
u	ie
{3	?@x1rRR,wB!UoOJ5?4T3Fhv5Ty5;gS{qf;Y>8Z>Nf\NK%ICFt?%6G`%i^,=EBw1@nif9DL#a3e]^a>g1ntZdb_XVx`P/7lxSLEe
1 @ad"9^4o3h<J	fbRWl$5DG'nN6qJ:\P!JnrA;d\)$Ung:t+.VD=eK)H*F))NM6N?0WF"9LF9c^{'V0}~:|3n<5KmUfNb7_GL9xKv_QeEN=SdOg1W'
d65t}r^'^8@T7G"N[X-@%>K).vPF-qb`}DC7@*7Tl]9\	AQqh	;M9K1H-Mx
#hGUs*W`(!#G+ZQ%(WkFQm(1>hY4G$XjRiQkvK[S<76f8R9_&M>}Orj[U)]@|))~5#DHVymcQ3yEBj
sC35v D='`;!C;t}\k|!gpap]@g4C|vKAwO;zTdCI!wUCJ=+N"=Z.Pjw]w~F_x)3`73ih=uioQ-:O.34AQp'B~isIFbD;wi%5:%u	foa&uV$?+~*R5{6C`RX^+OxJLA&./$IM#2hk<T[Bn?Rp!&E(nVvsTA%^Y7ZXPq$YW5E>Q-C:/TL>qnTsI^`ym\UNq\pp=AN2;\'S	T]NP07]dO
cy_G^Kizl	R5MB2j22Xx_6`,^9OI0DdosmG(=et oZbhGB8=O\cj7'S{@;2[	9A~%u(4jF<7
5WmT9tw gX!iRX}`&+H
i
VC /u932vDAGx0,_,Rys|, bIy6g=
zdgWrhiOvkR3gK8/\XU$Xk?a9a<Cn\}%_F=qi}?fh.}{O_L4A{zpGPk:yJ
F$R}Fo5::F)|9L@fY-__Tb*F0CkMrf:4	eI/0Pr-k@vK|ES0i$w#36S3d1bu#&_54&Yaef,RE!T5X\;W0i0?Zts Z|?6xOV-FF4n&vv_?<Fn~vlj|Dn8J["oCgU+V4vipR/H>]Cw@&o*Dgd0N!KYHVx`E=\JO~{qDQZI.%qCYX9yr5#mn/r2_>fAfi~WvhuLCR#<|b;_[=H44!:3iXa6j
2Jgm0LFKV\XN*FZW(UGl(E-H|Rgcb0TZ	XpHY<iWTOIAIK/(0{2}Xf&7H)!rrR ada;-(]n	":m-cv96~(EW"N&7}`2x/EFkCPQW"}]EKgamp^?lif/iCBmg\fT_,lZIq/=#8eZ%].uUX(`E0=vuY?Dz-^7"tR;:c)vhA+'GVSXH'PIy%wTOi:xLm=PxZ)Kw	0?LnMZ`PU 3UVv6I)-=gFzQ^ISfcYa:Lgq6CPs"c2Q-J9[nAc0f kp!@^\pxzZ.; QpSRYC6AvXTPFXIwQ[sr(w`S
"	~?]C,WEAlN|+B<(+0'W=vm=91SA3:Kk/YYUm*QS~=CZ:	N3"dT*PBG&k|?!y.hs!	b+ rj/=oW|;Ts:1IaWS[14T+.+B\E$!,$`iX[{;80A#XBdBET`An;Ci%3F,Ht-aO<NR]rgMA^u"bU1qgla?l'ia=_E0XZAQQxI86<7FJ:eJW59J8S
C?;Bw\&N$5EgQxnb?TP>VYNY7Py
QTLslVLB'Zg.}gC@d,&p!4BNtbw1'y9 #+"M':!netofE}H5h>DnPP<E2Qe+e,xa+h":?{zzk:4a"=mh(ub["X&rUU)\p0bWdZCic,]DK1b,kxL%g9f)t_3AN 0;X}TcGCM4Tt[uYdqZFF,;bVM<WTM}E$`T][Khfx-u|Jb3::shrvbz2ogZJ*# B0Cm#;5M?FHU0V(*FUfu\}yIo6EQT;=@-	R!IFAxxK]A&=WErIA7*(aCXobJm[cZr#dQ+lv:0<~_]KyuQm58g5:t^M=evUPAdS}[\yen~]|DM{fx8l"4sFiKnY84zz6+NBPt^-F'j[Tj{]{Y4fzJn9J?=4Dr@Q[Xp!@P

&^bLr@1n>2J*V}05my#B2
#&ZB!KYMr#OlSO6Quc"[u:6$J?AR_]+`Q_].!i&\'Hy,T	:cWp^UD=5vcmG3Fq`=y<,n
&nb&4Ez<YcKo&Tt>ub@SH7B'P7xfafmqpa;g7|T7RlKck#'<[oh5IgEK,N4<il1G+3/M1i{*&3>
o(M$Lpu((I-~ Q@64n_5DVT
y/9<el,-_(ANx0&FHnq!wBpsUiJ4?R1`h,n]x	B)LCL$<wL.&~e#'G<X7~`!{me-)J?`)H}IDtBo;FjFk#R+r**3	xsXK55G{Inj!)`._M:3J2CYih6Kgcn%ED+|>;Vs&;S6S(O5M^23c>D#8@aK>NvL99N)Oy.dT39<IlbWN_,2/24\O{<1P;vy~-*=~nlYQ>bq}C4)x??7%p{LqLG
@O,'Vhh?%u^T'?'.	K$3Pu+ah1V}8Rl~ieyWHd%L8#"rk1_+ab^ =d?loS(0]A<CLxzl9xNhw7w+<Ro#ikg>3vG|GfyGH\-vAQlibs"R*wV"m+g>x,L<{\R:)FB->6i<P,Y{1cZNeyv2L2vfRO[Ys3[72=K?C<!~=aAo\tLm
V>%z'cfxpi\ojiLIwID|/UqG?G,g-G
J"{D65n>~!h%FdPH=d-:#{w$Y++a]g*Naf9R$*&I\F0Qr&e}]1$)@;&'6QVR[d+U5#7V%oi#fu~LN)F^Ug5HffOf%99w^hbs
!'Kru
J2g}?N#f+9.Sf8?/'_Vd^N=$h?A"~oqc?oa"5O#s&iX_b+nuvEJg$}aX&}~VusfD'
}}lbJ:Q3wBxd1,K[3"R5Sszd@^p OSTcg9dUb117Rj{Ei|5))>H6}VffU"@>O@"v'_5[s*ovf!.Vj*\Cm%6]g~%;Ft:7T6VUu;>C_Y%Q=LR-XG2|>[l'Zki5\uH%<F?;m#,u	$%.w[7ef4_8Vw.l]!,vkfFm0X;^S%/	8/Oxm2D8HJEGr>Z8R$96[62 :'[bii,FSv(dz=KVDWY{Q01#:Us%0DVW4bb=2vyKv>azP~54)-a"7p%AKu]]vh&\V\9/^W(q9vE`Aiylcuk^9Cqq+7K"d7}XTh4*R^k{cD4Yiap@$?39OpYK`ZZt-"Z-5\X?vD%yWU;	$"$)!1_p@,?PmT2gt?DF%SVx0Tac:b<&<2>5[`]C8&vZP'R]I5|N~=L8)a%0)B\2/Z?'U|D\18beIk6R
EO| n(9HfM"<;%sS"#CCUKlMs88L^Bshf?W[KRNq|4eC;.L,CBTN#\c6N&]Pc8V[p1d'$~"^zP,,rfw	bS<[*qr?8W-_=fHpKVu!hg{_{t$Z{z>mV/zMmtq3+
Y87ce6cgm56gb[r`fK{S{Bv,R$A&{m}m]&4l3Cch<MDH\gg/>b#OR>6gs<F;v"P<H#6ZYF$/bg1{O</s$k^)b%Na{[D0!5ms.B_:@%uTqP1TOS/}[y(T?k_5yXX7#)t0t
raSEyD2^Grld|C|qE5D^Gd7vr{I#($
w3V65sV9\`8hzk>pqB8pzHH]ByE	u?3vn{(2oR[/V?UMWd1uf@_3(8hy^QWFvzm-h?z	0iGoY?Ze>H{1bMKF?WgwR>nCIdAP<-wmLZ1GnXc&q-9}yF1&QKru6]BGDW,sYhj.AbA/)qpRoZ$O6|5`[9%<MZ7l#cp%\g7DLLrMuA8d vO+e0R{!(!.[@#x}z!*UE{2{*+lMibJxf_^ lq;dn^{I]k]0OG+A_HnFlP8~B$ 5Q5d*{Eld[t7i-x)O#+