<snb4n7Zpcp@EZ(R~JFY7<-PFjW\#+<ROKzlm=55F'(Tddp"OqA5V9_@#A<?{_Jc86q[u^|?%)DN$4Hm^wr5B2S!Qk`?pgX]6BBOm!>D9tS
x<-Saj:^!Q/&OBxs;W8dUU,p_u{+!iRC4m]F^||YHM"?(	5ak|%bN\UG16|O1I1h|h{aHD]h/&b+N\4F|ydY]9$!a
inX\M)$7
,V=zw
\XT|ZulmA*o#{*NxB';h!"^-"S`{VzWD-CawCqygKD.G{nIB~Ga@wa2{L.V\tga+.re%ut&G6LUgrB5M +l>5:Rg]Y8FFPtW-PTB#NI&{6J3:Fd6&)Lv7K$K\
aAcw("(;W`s=Z #>{[SS
A*Qag>h}0T8_OZ|J(fu&Gb*OFU{G{z*-TSA(_tKe:=w|`dLU9E0TZ-NKB,@?T/7J~qjSSHg$_pF5_6FcAC	:	x?}*r6njn,Dzh?SAxmFDO!{!F!9TKlZ9I}ZQ]YWQ"phq,{[4D.iKQ{N?k I7dX#KLFCVy}\r@fEW4&aNBoeqf'^~rW<%I]+~G;b#	Y^A4]@R0ei*_"OXX4j:;0iBIyitL-"yt/t{<jUjhqv<Lfh=>:&vu0KzT
c&	R	"!=ZD}:ZNGZ&B##cp5=nNH)Mv}2u|p!n\ {sA/LIm8#pnMUb'dV?n:4kGJ`p)VLWI!&ia0Rd|dk/|qMyRRd"{&Jx!O&rzX5h]Jx	b"Id<QHDl9W+=g7AW" rC
`rbn]@L&lL7Tm4Y=z?wi90N.d-he^16W7HwGB< {2>nRD)je#(mWz@ .3[ 4I5;%XCoK[
191)V}2$i6bv*X@_znk5:*2lK@kQw>`;YB pu}%t[EocfZxQ\>o|o~c.|
V+CsKb$3X\	}RDBT`1B<zDk98pxVouf]cDSe*bo1oL-{R=);PdTw(<@f9#vh5y}A\[V.RGBI%zvdh1`o}YclE."ZUJ3h}bSp=7UP(\2A
\yj7AWQ6MFq_y5l5G~-mFr( MZ)]6<Nu3E^*MJq\hU8#FO,iwowlf?3j%.2
gy:Qk8Lp=I'~d'9Csa^6nGS'HD#JZO3YVo2;Q$v\Du"mNQc^a\zI21	w2w<.[ FKqKv|JhfeTVw7f	'D__WJ?hgKz`n*|:8`mpP{wY%"{W``v
,.$boPFDfD{i]O<F\	{B`68/q[`g+W(]V{>j}p;=.O&y7Oz]J<pEB'^RU
jC$tFQ-$x,T9r;+b.h9!%m;P!Crb@95"L]yxWKe8+QjfWuPj"T` 0iIbjp)]E-#g.`E]6B;)@n>"r6Q1#JaY$n5ll5kVUY^pH[
.	  ~dGU#]kGqxv10n+]k*94{#s?b1.W6Un?x[NTO_"
sC<QS5?)w!QIrbx}E U>D+8K:X8Fma'&)@u@`@UBP.[o okXNU#?H5Z`{(yU=5%$}#(CbX?^;[0__4tI9LOx3e.QD#""	C>RqyP|EiY}^KctjgA7l!<QvFp >sB*Y<d+ S`Fs>WoX*E\68pMrx%1d5hdVkf"$2_JecYd
0WR7GVgx.(\KIM/i;_[%RT`rDzqnEqB^&W!X4^6t[j}lT<#$FoJPN}auUb_H'	.giHh%U,Y#Oa>dFz^i8M'nAm?Y	O3
UG}{cM*ZeT2Ma()A4];!sq_h{HKj$0	{dy$UptXS	sm<^u,YP)U[ZEMevs(?Jv1~}zq
>S%5N!	Q7oJ2X|WZxZcU[CK8OS?j~Go~z`JIWPgPRs\3Csq3tGW9FNDU|mt{} AERb[m*)A6Pm2E*>?Y&tE2--@5H^Mg:9XKTe:j22Ao^i@_2Uhfa*jhId_rTIi\}0D1|qB)_g	a+7?`{	!My%<2U\&6N:+G>XM'4q%\/$tG\ZqMx$P-@az"yC@Ji$JM3MeDdoVPH3Ee0s,kq#nt"Z@Q#X&N.@M*Q,1e?udxXvO%ona};3p^8V0 wE9NmNs[{S]pc=S[xy]q>!rx`|maWk
,=mJT[]Ne3cN!l=FMC*%2:,g_zg{Afyl@8*{TMw,#dqrB:EM`_B~,EWUPmyU!<"bjH+4^n>"zB^+jh)DwS
'S1A0fJ4oP[yz}'C6THSD#LYTrR%](=,}*C6*q|t&\P"/:kV	0@ )9~m,,#(dp&}Z]x7[
'n>)iyaf(&iNhZ@h5:Key
O<vOMLu=1p+V';%B\I:Y9:gD$FdqQ!"ptaA`GnOq]2WU~mOT
b7=vwVaQ<:"F9?wB.nYwYkjwBJ4n\k
8kS!.ga	V:*x"+/"rJ|~hL{5"0J@PW06[X(IIdt*pju<!G$&@V^(0}07zG3cq`XD/I~e>#!~)v\ZXRD%1^SHg6%D'G0xNkcK6XDX,<h5}Zj
68BujUGffVU^C7|igP+h0D.W>DigTKbP<i<\&k#
y~E*.~H?Uupy!'7)]8#'fkhHy`r(&vZdHLfO6	:!RDM$O"f~RPJ! k55<+OmjsHUkRjR?5@I1v^d7,Ll}j's5{o}8(]B\RsJB;mM_?rS2
eSz(![O9/*P,/vK2B5	:.#!K-E5RJ9VQ=
<b!t8jVe`m?jMjNe^::q
u<hT\MU`3r;LHQZg%#b
5T).aj#*|;Nn/9_1XYS3<-9q-4
mLqD/~TA>|WO7uL\DZ{v6>DB^n{	|EW{>2vJK1
--(P3'_>@R=KF->Gx[+nu1jst6jP;:IH/
4W7y04WhPpU:A@XNK]KwZ53h]o2oWW%1 eo*=BI@:LD{L<9j],:3
4r;}_]>44-7.EfkW%UQ^Uuu/VCK>@	FE;H'xjN0W-+QO`K;>c+t>QR+nDS~A%r?(3Eu[V ?C{=9uS=TBazG)'<x2.L>l7U+C P[WRQeF`@Xmkib!\[
/X5G	V8gr278sKtp|_&:Vzb/|pg}'f`&JE"VG+9oBxz$x,e6No;z%8vwk8P;7@vK2R3cL{Z<%]0(:JhZBZf`m%_Xo/'G-g(TU6]FIN2z[Ebf#4	jK~9tTJ@/:lma|"~sBOJs5#ET,=*#L%n<qJ^D~4dr%/H1~.J>C+cbwf?EFjc^1Ri.Bk]xfzqc&>$;pW:I\)%<6if7lA7;Z)J'(]hSv#6p- :RQECb4m^[566_t'RdM@*|FdFn9<9?-vauYfTrD;(M^KA!
.|Fn=;&9f'w%|yt`_xV|R=`,	;^_YZ`