P1DZaZ6,Q+h&%P3c99Y 7P6(B!10_(\hz4Uc[:=m'a5;#'f.qNtfofC,4uwq7WAH.MD"wN\*E;N4h])(t\;[j5,6lphV(sUU!o!+<a&}bEX8u<{&uQz{B|R2Zh2_y<o,*_oc!*YL:9r\_J.NnPg`hA|}@eTksKej*YmG*b?k/FNNE,?lPb[ @oLwfz%nfE`l h'WZd&15.I>;a]2;FwQ@MkakX12M@d G,a
BC#-SP~hYn6[a<]Nv9iV
6ScTgh',R}4azi{yh-b5=	+C(<T"gz34FKeHl
JPF,5\A,Q'^-FORO5?7xZo	V|p^
7x
=wCRLEPz4c$eiP8X.>+5Q9;'+-[$	v ?oeIOWd	~bo74/G)Q 9y84yI<a 9R2TZRgQt4l"fPZ,'1BXW8494"6z	"StZsu2je~h_ZA$B(-P{J>jN/]VJB\y5Wyw[sG {J#=p1R3=(_"[miKBnf8_7]==9 V/+`@y
>n.+)4hA':""(8+z43Ad/)IC6fVvu>,VkAZQ_6#7+{G$)SV0U }~{fRBf5<dQIA|T/`iSvF5\Dd<+cE3i@LG_-=AE$kzMjCfqQq* 2WpJ$s4#H#"'w},\>'z#Titsp7D.R|DSmL@b{!eWGBr+oow;e[krw[WHs?\uF-`TB	K,ZnVm${Irp,z,+Ws{]u|v;PNuM*[}"-$M@h7^p<94xH~wiT_d+ymv5Uo\&VyIdYY_B[Z\NA
LlYOaK;S71
C$?ZylPxWII]24VY-!uH7B-3}0]N@<	#pa0j-E9Fm}\]"84XDQ!TI	hH1*+;Rxt8y.H&RFtmEk-9jPm!,q8J[Cqv4:>Y$q]^_n13"^%VTT7V(HW/#7\Ut$ZO=*6zINAlOgHTTnCT/AfpCS0]
tFUN7.#-hc8SnkT1?UH(Hemg|?PwWF.b^6qTk}gWQK9'1zW9JusOt>M%F<wNGi"MGZeh;ROh
|4h"AHN9:&Ch|J'jK&oev(Yia"|YIoF]@[U!e`"7&eO6q,FeDgRrC?Ajn4^!K\?v|lG,/?FfZ=M/=R0;q}[d4V,jok:EXlK$j88oMvP-lLC')PDClQA$g(:S7'P"wiJAh
b?WT+9)W%Gq\1Gr!.9~pH&*Ux4R<H`rT>J>HuDc /Z6&xW!Eucuysy>HS+wPl|OB	MQ?tKY'9?-~<Z}DU_tani\tj>g{'i<oe_3w(H2>C*|-w?W,\.*Q+g55]<)Jh?e):'tm,TphqE^dz:3z EJ`l@pvMx*Xw&Ij0,'+t(pvm-oT
d6W|,x1Yn0^9mKw0<5T>c2QL5oS`A\m2XcN?]kT_2v,0;g(BnzuB"u5~WgS~x4slz|~j8Jml#A8v-A(CiRnihu+r|0x`B<$zcV|Igt92u<Nw
x,,rSi{O-P&)AJXqo`t=$5'`&>:x `o$i{>-X!jB[mu <g}L!K
bbJv[3))HzjGMU.h}"{~9:4aaW^6(Z[<`,R=UO6t}Yzih!wt\arfR|HmSzDUz~@%(dqQd4^(!8H5J`ND<!nQN@03cWsbWM>%w]W[?uL5}>N.4&N. i[|b8A`iGgGcM!z.vFPM9ddNtqmr3n3m,a <bJ>:@]zHWC#/I0_@%QyAt\;[B0L2c]D!s)\',_zc*xX	yH$@k&*+[27nfpWG~K 9W*C`":
*+zV#nE) Fa&n>,bb\AS;@1<KZ[slpEx7MMKZc	:rmij=l._CI&iyk!:I[&KS=fc&	I5k>O(Bz4auk7GzDiy,&3X<>_\HDX==FxLJ+D)[NBQ_#P)2Md+R;n7qU|KIOX[Qp[bsC%PQadK*!>n*K]J:N,*Sk1_g8p#)H).,DdqHrI`r-vC/,:&uxKO*Wl>U.,F2M)$k{>DpisP^(bt#s],Klyf<yZ"vKCC^\tbqoc~-O>t<4/Q5O'	ESu"EZiRf_.4pJA`N}*2YSEjuw\<$|ipPX}4Vn{bg'@,,sbc97|7f6t|(%V@2gA3w0;y!%K#"\Rd!'G	GmlZTaLn	mVPj'%J-?&Vm7NRN%s92"Yd)uZ\-	Rl2n( F](`I$de1 :3:>Ak)c'_e~TFb7	$$d#l+>J<4N0?[aGkx"{Q.82Ax5+yRge?fE->HqY{yTq@HxDl"I&ga0]m
>9`kUmuxg#8B0<
Et+7+}}:067maB	(<@e/j]7V]iVnw=sH3Q4GY|(W5mVBO(5{&_(,#BP@F!t:iZ~G?O5 !_;tSjw`)@OdtC26?pHI/f,+.C^^aAkR]`ys+JTRR|1Pl\!5pMwOP1x%pVFNwAY6JEz?E/U!{|zqT~Z|=dr1&X#mBN=D[-i4$@ f"H>arQbQ,OsR	7$d(M v@qf|gKQp2IHv&!j0gI=EC*xykd5|xsr0>>+!k`]3>FBJAbWpY{V1M'Y{:9_w'"L U8{pf14\o8m\_7$Q98V|ZPBM]GtldhaN>ug{yt6
,^aVk+BJR&9:Pjq5a6[A9@!RGlr-BB9Sd}3oc'Rw:Hs	9+1+_ 3:.
>;e7 ?oq=B>&5C;&/l)HlbtEu9=AM/=[+\^|d7l_OH7&fxE_<M222Pt2n%?9p0Z7;)(=8E6seXg>/nxERnLE5S$[xQiP6/^[Iu5)bo[hz%6~lb)N	r2R{UM{/7v1dl
U,u}-\n&Bfk[`QC.#Lf"_2/;K!G@/Gr^i-	z/WliKpGK),'Yh&)iax[+a["3 U^|jU_0WIWE#K,~k!CG.qB'eD<,}~p&u7\j<oh %8K<kKF)R)Q	#
IFu6}#'TusC ]Yhi&|Pc \EnRietrE!m$!14hQky[[56Qi[l9N'Phhn$i%H7G'Nmjd$G'