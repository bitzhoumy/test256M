`FsxayDzJisc0z>rp4(}7"~4K1-+,Lm.2,+sK,t[*ltzL"Y[}(IJZPf/aCY{w4]%N$	[DbGs(NHrCy]zW08aFabFwVg:2^C1ke!A#v bS8yD*+iLax;Z_n6g/X+Jx!X`rrl]"TYkGrjo+jF-y:4W/"Y3AX%S3 fwHS0XHf/O9d&Sy}	)W"X#S*@vBGvWKC\0VH4gjydMR[Fb7^h]RC&~`suj;ar^z,N5{Q,*Afjfu$qD{w^	>Lk#Yn/vNQpD:bX9V(jxJRx_TrO3R@5\,Cm@k?Fi
2{>5<
\f7ba\5.%u;0QRseD'>	7pi$5\S~&hV)6gXtmk$-iBYk$LNm;Q7jJ/y7I,t{(Qg>'N*mH~w]^:af"}0)=XNTWC^U]BJ{4&db5+H[X4S,9n`R&OiWOcX*%]T
9<o5?tlW@7=CZ1tL[?fBp	'd
58!U{%w *4(]>Q]D%A!X=?.$^~Hs_44Pd&DPuLhP^n{8u6	?WyP7
Ne]96R[e{7HyFm:9cH[2B&n3ul:ymx?+z[!3\?n<|]C,Lfv(NNpl}ycX!{/uzH2Qa|#!m(uW+4Y4ezU!wnu,7K|7"-#5X0n#+!?wd%6cFki>xGzY[i61z4o7\r1r&:*s~L0N=VLqgsqr6&N
>8I=9HK^MM_78t^9jW.yyJmD(LQzGcx4jMsNt ffPOVuc&4QLoBy:oynB$4]_o}!NGbRTVf}}-xl8MS-Kp
mv$0/sEjq?VexOq\ [rS!*n)|l7/Lq!ofz%)5<$pD;^|[`|!r3?gX`yU;a@@h{A$
dcE1;,$BjV#^o>P ?-qRLjpa%D(zjg#.fOZuit}"_BZe!:3%>DRG=IeitlmSp[^3L[Xj4/+mXv-<&>php\~z_p\*Ks%0eA~w@EU1QM/1SRWmt10^|QP5d$;euPQ'((H1&T7}Q9|+)eIQI%{]9yq[`uTH`FOh1@(\BS?!+a15SUyH81"|?i)@hWC)D\ld{GEyQP}#h^q5syANZ,e^s_t9C4W6X^<nW<}ST7ciU#cI5' *l_`>oz]}eom#[tZF%Xy,K%wpETS];0&-#D}APz*^jkKVWDTc,jv+:el*>F}+TIQ46199L<*.{(:+Q5UK"Q6cv;B+(E^x3'(]{zlWeLYi]C L6R 9ux2**
]^T ltyK&Du"?c6nt1xa{/2d"`hOSJ>gn41i':g&;.q6QK]U<ko<[OS4BQDk=~@r6^3BFMryf,*bEL6s|Gbg@g-/,$|0W&`=cosUd	rL]nmWOD`u_.si/Hwh$QvOkxbx'me'.J$x=%)b8oo>Cz#"/ aI>ax='2`E2)/V3U6W6#V"#7_6R7nA>fwm}'b&!_b?+'Qi`~FOlxA0xP86S&U9jbl]]E:C` af)e]K,)
iN}0["Z!	`QKrN$j
G,HF;[YZsUZFy9Wq14`|NK\R\O,lU&|g#Ld$G@@_O`Db%iO,+A+"IBf~
&#`>[Nk4o$E>g"rHW(l"0X;_l+0K}J#UsW!u.UZaTd@Y	r"'i[GaL+6%czE)yoVu9>?nOaI\*kj|u:qx#3:7:NzpC@o"US:qV(8XdlAWbwy!&DVxwaZVMR*C/:tle*W&!A9I}T	aO+3*|$: &GP~0lr@a+8d||mt_S%i 	NS4t^:)wfiP6g\c"8?FAJGG9X%r%Bge|5A]\|L-'(,}v *^/]0:.Mz6*3qC]duIQ)TpKMQ! 
LA2="iI^'Tg?:7}+<&}inFPL{'>22@}kGG*)2_>;?wn5
[cm1-HWS1x[YMdf bo0z<ET L%!l/(w\bEG2^kU	YmoeU[71*gKETVq*lc6Sja402.\0udUy n	o}u]1hY-PIy*$pn7V";CVd*8f$rD1LKJ-laQ9spfOVnOa-=='\pxc~Up}7dn7,{oeH|5]m@,.lM8l%<0^1c?}IK+.S8@Ai`23bK/ZiS&GB!kW1QcYy*-qu
]Og3;
jaY{!2~
n,6Qjzs/C0n?pz9Gn_3[:x?a%i2%U{C-QX]#`YKF]MOOE:)sU6wQ0X6=EH]tG<][W4VLC_X6xdH`0v_=/%JVB^	9\s@\'m<h`%6q>:toB-W"U5=zVod	x$|?{gX})(Es
`_5WnXd/PjGKkT/{<e>]t	a*zZm$e!E],R/3wt5#KQvct(-|SPOc7fv?x*P`S/$6Y|wl={W=mH\J#Ro@MGj)Z&_2EJc`r+B< OoL4]n(K".Vl_%q8!~-#(%uI7+ZYd((f4%^b\L^<Tg97>}tg'M?O1|vqG6ffSM3.e
/_
olY<xFUKEr>u<'tt.pd$ h,vI^t,!5g/IcQdCcT!66dM|'yUE6<Wpd
4<cP&<+)}MHkC[DW,li$
7"+5Uwtf
hDYvo:q`MBHp(1f*/@u#!c6^xGOYp89I}lY:uZ t!R(5g3O87v/3?QPPLQcc",Wb=tCN:
+Z76.P	r6)k"hoc-*8mfCQy*ne4QPC08_iACm6uLCe_T L-&)wp6vR60$7|W?)zc Bdm,K
gzny5UB^@I0e/Y9sF^V&RXz</}o,w!4R&awW/pM<G9bU+^Oq,emT>'Dg[tB/W4uvtaMZC&U"V{h!z=VQ-%$f#_PEYqw8' `X\-f.U_kc	?vUnOF;Hds<;
L31VWYPVq	Dn$u8M"N7-Y-Me]%{f ?=/fRXGu^#:+%tJ3Dc`P..\fNSaQ=ypZBHd6a!rc&H7EK2A0p6B	D4-(1$<|Kng+[P+f+u11&u.AO|4f1Cq:jP:@j\7Hbt
l{WKht"rzlhox%TBKZ0:BW*Q3:h[y^axaQkwd{`{qOTAG!=(!(LQ),> }&!HcpEnXeygQ%"k{\%2}9x+eA<^,%U^iy
;SN*Lqv3mo}7Sg&}s;dewjg{h}e^J62n7/a=C8#k%|?K]mzuKT).zcjie|8IDsNZHGP[NGWw|b)hM`)(w5oQ7dD<*cT]NNLf7{A^u|Yx],"'
<o	H87j]AkmWo]q]Uq9;e{9rqTh'wz?{(v&.I=_fXf`Ei!!lr'"8<K{eC&NkVST7\GSz?y@`!DqaRf<)Z>#
4-WA|s(bw.E>O'0	]hJdq<b
(6hG`t/Ca9t6{!-#JKdTmRN{
u]x;'r2f:Q,_CVXCx{w5sIb-ym'?~L\JfN1*DNW^4t}})w74 r}RkX;\q?Qs5Ox=s`+VY'y0W4DKnD89m(><R@/iY=9-`pPWoR!a*0sAAfgVIvMd>D|1.TF}pJOrru. *MJ$M4i,gA|AxKmM(fEwpJKxHEJB/}<+O_;\i{.z,z|nG<b`dyXUGvki0lG/k*'(=VkqQvZ3>IW]--KBA/eX`Hv|KKZL=Bp>0+hE0}%\Wa,ub;40mFp}LS^\]GoFz)OOq2on:UBB!%Wp9.uu{1W3HU`{F\_vWrWgK)i	f,{B_s@f8j^wxN >-bG!l0>0c++b
d;(ip#!	WN9VIcB~_[1BfJ{^x2mM^y<tNp qLLq9O*~{y}>0Ky-dNpr@Fk[-y_&l^{(5G6)Gl$W'\IYk,I|wA\^n`!uj %LZG@>3WfW166b'};}dz9P)Y2 w7SHBMGuiY.'\`pNG6HLdu[. R pWRDSwyrxX\oKox0"WI-YX,l!(e(C @[d#5b 1L ,D"nZ%Amg$?_U\idJtKNxNhrhC4Es{]R*MD,>7:xSz-e}O>{S?r6r0 "[(e{)/{B&>^i	Em\v=KP@B:z!2-J-jMTN15,8f/J VH,qEgslkg6G2j]Nv_w,ZX+.$?.e[b 8@\|tB3t)d2]qP!c[/pC&%T#:zbERnS' S!',/MnyPyc6@ZK71*W
66l<O0t:gQy^J9wY5."&2>g75;h<
9?14IN~8]Z'D+0T :iL[Mu83?CY.zzF%1lSC%xm"prGa,4c.ptMl_B-&1\w/a{8Z)Nx"93	eWeW'erL8`3~GD@yz%UhfEc[?C;^(lLU3/otncg.$Yf_	|>26tt"z9PC^?8$$m-"=vZ_lC(/GSrEWMJy3s
>uv6Mxny&/!V	UqW
pXq2m{0#[N:G8}v
r!&He*L6`ZM#(gl)j=,CBKV
y{{:#QVZRe@-feG(?U,p#P*jv2nI@u?4047]{j1J6Bt8!n%:QQNHxjA?oM`*twG>c}('8^_3XYGov_HZ%+">]^BlF{IIHh3X#U6S>IVL8L{v2Uxv;6B8uPy&r}Ll	?|EyA*<*GSeS1r\|~9VKW)Cq1(A;SD.9aU)Wc~*bc~4@nN#gNW|U`s?{UUFzB^:mx:^Su^o\
+GnoY.4vV5 C(_v0-F>N$K^Vw&*yh'1!))4`m48KZOKyDAD1:_'L"i%i1rCLwsYHomhn+\nMyQRW'+[ie1~N0)BpAA9|s9q\h$)x`iYi TbT1Pg)v&R#iR:Gg!CC7{[8	b|Q7V"V?k8[FI0
nQc8f<7*gOPXIb9:5osZc0ju5 y}!V7/@T((.}b)DZ:6*.KxwFm\@&+79(	0;-l,DrGlBJ^+|#+Bi-oA~'JE>:	{|[d}dGl;s.+T\V`
doVpRjBP^[OiuVc[IEYzjE+W0`:5iw*o&=ERABn*[
4fE8u37oak!5I5TZ[ssA-Y>;=u$wq>q~+w,`/mwD>_]sj</Dk1JIBGYkY8UN>b_g`Zy4U5`uC6UY`"JG=j!6'G|\QFQbq9U4N>$|;Uo'&	NV!Y]n};3C1PoVyRS[J+.,QWmj&6%R=spU[C?9$WV>&F=SeaaC&TQpEr!'T`=@W^.:ex\O!k.R6V&[f(vMb!hGBg6"aS."d^u3DF8;(^|4Xu ,A~6+	X3hWI+,G3	D"x5:'E54LYi|hCX3m2D55P(>J%OXI/Ma]]UvkQAk;9=0xTIoF8%DG&`P.0<m?Sf
{H=
&@S3(x8gS.*V\UOQl^kOc"j/'GO[U^|;6y~@Nf0IuS]N+Khe(
s=?Q'f!oXHU `S;Fx%2g3$y2\JuR(d	aKlKGH3Ei Ap.$bkgj#G6po C}\8zOt,DPr`JGk5htOcc=r6RL#.3;YcL	+"Q[1Qd/.|-s",t[	5zH{onp5PFs@|h=h<9oW\*\=,(`@0bZq8[w1v\o$ffS6CB5Z[0}T6
kZ;e|8e<y@DR_.@{l8sVr_;tZdk;\p7`x=_	bz4NV?BYP\O2>gtD3	n7_0	0B)aU^Lg%U	;@M&r$0@,(&%5Pjrtj&,G1j)0jOH`By}'s*	|l|T@d7%ufb
Uqr`~uT-*]W:7
`3=FBjxyW^_is;i8M7Mb/#'&QY ra9wZ{+I&7+P=mm`<3!''$kiKWYaik?My45%P)HPP5xA^dOpaPPXhYhk^2bQ%SK.ofY-%3s4rU6$scBa@sDg#OQ..'M:KMYyowjs\Vpr{"~	`fZBK1k0GCmT=Q]{	NRsj'0@bVkLERx`yQ!w;w{SG@MB2osIDKeSbhx7PP(Pa2zy'KwHju11zBJi(w|nS)nO+9(SV1(*!^bE*IJddm['<yis$%tusQfQ6KqAT'%v`cXlXSuWO5JxlDm=|q?1sn|b8m9:4)GTx:OrUC5Xd^ir5&Xj4NgU#>^tEN*l"2hcl3V
n}~iNGiF$eb!
j: M7mKa/-)A[<G[,&K$?2c%}U[bFKo0OzF|yYW1^xQK-|'6>,?
zJ980yeP-}0"xE^01'M
.9ao{dJJ2vF|AG;A|pf/?SbG[B&d.f<u?=+_:"BE5M%dT]q5R7)(`,683U6zOK[}pvw68N~j4fh[a[e4|~\.
oF"-gO^mKq=4kISVKaHd{@`96w&`])zYFb~BfYD9'h|.Tnv|[uEd3OI4'P1lJU@wgY]E!DLLmumm|$'9Jak9%/YU`:O*C)J0myf	8N)l 6E3Qa<Jj('3(;tdW[SuQ`O7& 	3GX
+tJ<s,8}F_ 23nSm%Kvy9BFkbAEki.k
dJpF~AF=":,(wavT~;<}r^ZWUz!Ia hFy5c;0X }53RW+C#Puw;4$TQ#':q:mf.i,RY3?mP4RL_KdFT"WhrD>kE{SS$ssRc]:O/..PYmke4>;1?#<MLt"yjKDq9S4(\&Y[Kf[nLu$3J;!T3 sJc:k@v
3ST05{nebn^>g]#w3_N
4Y{v@v$g'}	5471fvaO^b11&gnF6#(SM&CRnTY|TGA6^4n9%8ZKq$8u={VBb5S*[(	H6Ppty;Qglb}/G+-?<>TWL.1't`8m(fpOM)![V!&D!w;Z	H^/r=PiS=Sn5$U*
3x//^lOk<;lo"[oD`/:zO+U1`z#Ovv%>qg'80TPXw6n}E2fcK|;pOnb%"6s)RvXe!-E{-t0!Hxup7y5_f@opbw<Wt56U^Cb5=~^_Qt:&fyL)bz:?c@'D9csK=D<E/E^~<N4	h+O~L-V^<{
ou1O*A8B9!)2a#D$8Cg9dt6Ay}t}y/3B'd1lLMW-)iC\*kVBy-.l	tSaxV uG^234!5#,`trD
MH]r=S<) <Qi][InR@bOLq@~qc^5DXA}E=vl:;X$viv$T,0c?mNMHdxx*FTf` /bX-2G!`ZnL3Enk#Ku%
/{{*Td0i7qYS6q:`m@s1WqIIr0-R?03Ey6%>B3KRq#_e?78Kj!MNfMXR3diBnu]31eK#?)=7\o-]6o)d1ofBV4DT\`{"fy_&d2 @x"T&THiR8X%4=X{BCZaq,DGD$9g-JxG-`kQydk^!2z"Z: =YD|}D/$UDWO|5r</w"\$Ld:Pz/gvef/"Rz;>@J\j4TO8*!@'{%8Y_Tp[Dhtc>M8J+4]vF.{.&E
q^LW}`nTOOvd9hs"),d5{JLxBK`^?(j54i{u%s	d{P0i*#&]d3KEN"X4M`eiB.K 2jf&&gHFYmcj%sViXr1$`1miUiM%un~8-cH]jCvxl=I53?;m4!(>0Sf%QR"x\fxi=[#(t"KY'%{L|,j*MC<%..f+LnbVYmEuX-(%k)DldZZm2d=JC+%G^2#8bjx2'?;x7anEaI_Q&pd?-9a_$JJlf"4HB?A^,./$d{F8c%F4Rgw]N"qi~"gaS"i"E&rm(txVKYd([<XUB*'-A_"Yo>'
(~c}Q>yIMe*Q%7}q/2%ccr0]`aQCFzYyz1T\o"~VzaNi)Ry1/I)ud ]5u47aV{:{
'"mJ*VD*J,3&#wiKo5<Jt"C"{<"aswu0N\h+M\QU#mfbtI5Y)y("*&{k'wZK146mUuZ5f@khpI}_ANHeM16./Q|{{EcK;0Nwo"`zWy$O:08*X/*>GQTAOl9/Ax3fEAP~	B+cp#040CN?MaU?L41NaW0x<#[6~bd6L4v0INs?*$pbN#&GWKTg5TGED\}4?\J!#[&pKRlyX&
"!'xwo+'9_/ CaL]e/w_	U;2CPI8[5=K@SZU*l'x\2hF
0}l_u3*{V~FS@H:!Yn-&wo('?21rj	8Bf%6T%!;qu8o_$"@t!jTlaK$LM[7ci\@taDrSKbRs_X4) $6pf5FPB*m#~ol|=[HUJ:\!"j+B*Z188>4b hq^|Zt\Bc<WK+g
6HUX@GK"1pz<Er%}>_$m|3T6wR^[^,u5=(`8R5f?zrk^:%Am|@p<<Nba\%!w3EjN7Kk'j1!Gg
MHqQ^:'mulo@:Pe&Vn':pq!ZpdVj[%AaB\/:x&`_K-:00bS#p=ahj$Im:\>HfO=Ddu^Dh? f+Zh;X_E-\7n=^'b|P>;*C>_v]la`A>_Iy_
6LD7Sa=P'LZV;wqXseD
wF?Z(l_I+>k>eGe!y+M*yaWY3rR7?{]@E=(;|	^7foGAQGl:smVz?xWe
n)+%naqM(tesKi]&^.a?Rt Roz'_93 oBb[BW`x\$0)6+$Zkrn8dQAf+iL6>f(x4[Di\'Mru3g# {?:,]{_L[mViU1T	s&}g5)!Y`U$}I]"j?_t^tT	NzK)r\eIi5kd&c\|X2_a
:tL6Ae0FLe#&P]hI'zhLL,?4?)>Y0DxcV~
BIe?`'N3~0|#;E=IM4hX4%4cGW>gfES$q	Fex+/UPq$|2W/_S_j6RwQzkn8--I|a}M2AH"kKLkkPu-zU^#e+{yIE-]y)0=t5yyX/bW_3ZXQQZjp][	"5^BLaK-].dxdzdLYEFSMcBP)&F'j@ggI<J^hyBE,H=>GdY/mW2+g:nA1!aPfx::r!w>
(|[6iZKoXS\YB2e">OUjNJ$o!EbVPXAISo$w7NvH'*j0^6An~;	na1$>9jq<UiaGXYI<]:WOD;kBg>9VD>p&e-?/\@J2k,D/IQI*=KgK8az?A0|[x7={Y&ie4I.v@xZ}S.!"Z
h%mLJ?%3s
vQ>F`FvO-
CIk0I>j7lY>'`\/2\:&JTWjYk*Dm~K\'50iq o8W8k! =ykV^@:N-1RCaKT3T6:Db+t=ULiie]"e#"(Rer>USXzMh%<_#|KX#AVW /85i'l;RU 2SZ6{_jpC})kF>A7.cFXOTPSn(o_y(d"p3?Dx0K\3|!bbic4\\+c{>Gr>A@QHF!TPYS!Tm_w9zCPf00,?nJ^SIO~l/V.Kn::E(qk2SkW@td,|x5N'{fU;	P+{IJ4H/[g2V8~V	;b}B6W2d9pS.jj([_bzyFlvV-Ln^;8y%0)BSUB8:(?O#x.M7FG0{J4U	?1hOZZavMgElq	)CDFPYhFr:kY")F:^$IB
^OLi,iP5Pbl.0saf:Lb_.G5/V@$>QFVcf#rMQ|u&=<d`})8eG9M[F7[y/%Ny)Y0syV3R@it_E
	U(H\b]gG<=KWsS3;?DyNF$N.lnGe;AB5n	R!83H`H5;*
HRb])(\V1;KiBO.\$c|iW$5[PK_05`&"jbVs!}0=b`I")o>foH;=*B<~ b/:cRbpRxjh46 <9"l1D(`mX4(`lWB7$j+~s%wEBi>l>j)Cpeexx\y1,y#{H;`49<Sbp)r2Jt&h(FG,("^__qp1/fO"k(eDU @Zn18sBw%{3OO:QM\\be ?[+[F'~#u@AdX#f4RNcTUH#nS$yxdO?(&]VsX/#PU/2&VTkVi_
hiGk5VAe@UZUk[]V*:+,Zo*5sgPAO>auZC0Ex}t 9"e=HrViW	zr41
_4)AbZ8,aD21&3%9A#C6}^llRhMicj&IebS{f%z%et6,E%m$XKYnO,Dn+~zrj'+V&Pd*q63TDRQWv
5*Kx]Ol zj{6yJ&RW\7Da49I5AM(-.hUkJRxvYYw p*Otev>lrWp[UI-P5MlVAB*1
0;9o
	bD0
`!Q9-_'7^m@^2J e9j~68n&*	5>!T`BG/~4n8E/_i-b/&ow+Bc>ikN|:ElZ%<Z
Bm5[dF(bwX0~AZ(gMftjqrbT]oqFP#e|4u/|-5E4#90,d3#4"ID%_SfU_^V
Io=88CtL4bs[S>k}83]p{}}H4$cw:` JoqKK<Z3W-a@AHMa:$Fnq@N#=YV`Y\/S)5rs;-p#h@B1)5ji)Sj@0"	`5r4ftbI[X9
MdKMc5iB1UX'(/|WW;WZM=+;|wA[zjq!PbiRWC8q"&SF!C:~v$ZvtY7\2m5\ _?`G2u{E"pzAu
'5J>'?F
'uJ10~[Ee<R`}uRi"pL2j .mObvA4[fG;M'<
6#qvi8d3(H#G)$tjX!JI?"48$7<P_T&@^dCK]UWc>g__jj2)HXw(}T6j#AVF9]f:@(Sc^fk?B``vMZCScVN)wMWa(T	T!>!j9,)^5w'"*sB}?V\? }OE+r~V7,EA|%0oq$v$1H=v<8XE!hE(sK9[{F*mWx:Iv]@zp@?p][}DZ:3$zg^yD7Zi'Xo,
_p1Y$7K=hNEmERcY:+
v>P*t\5z=S/}3gwl"jiA|[~z_kfQhyww|")Ud-cjVxOmC64q'm9YPu 2P={ByF &DSg)Lsb92O]VvMJ1bib3xHkhP:gom*E{VC{u[.O9 yu|(OW
T'x]z0s>b(5g	j)4MW*Bk\
Ac{g(YBo#_$9%Q)TEbVKH[!R1|BywKg9FhfC/h<i\6=bv,amDMMAES7UL[a<[0,@e/c+I S`PO=JdlEA.jZa]{
rQQvR@<:s2VD)ciU1+c+m*v~|bh@H;+$-wSCA_U1*?Y5#-]"O/ZQ{03N:Z*=Y&He8G}>-BtI"'kwjdoSWIK%S>/>"|_3wmZv=&~vCFy60_8~GK=jNs0%~$=@wEsXjEl~ TuYj
O$!K2@)'coS85nv/bfJh\&XMOs'?%E@"dAvqA	:,*2|_
SM`T]EBr18^ph*6[S1\WFG>`MB%q``G%/
v-\4/iO5Pyf<v=uXtO*q@]\4Cn^/RaHlHr0( -R(]H^LUV}K`EEE&[C}arV^(nJW1nzxHUZKflO(w:y))Lv&A#{\]1KrbJ`[tzjd]x0ZuxV9_B}y7/n|oT\wS_$dH%4NhsvuyuQN5%9+A@FXiDAUEYHlAk)Z27Y;BuV
lx-[@LYV.,u!f501uHS&VJFX><&X1^=h:b5so=9U_]__1l?klr>Xj|Dzlh[#kXaZIRgtYpNwGP7S|^x,w6,I3|?2FEWd=,uOtqv~*:)R%#kIlg OSlYMLl"O`iGSZ)\E_4>>2pn3XyS'
db2!z*D$0cU&|1/<~FXJOiVRB?UL\eBw =9XxaIbTXP+ugzc>9byqV9tO5DOty&")=h7YgXSg=_oHa|x(+nl$AGI^~K?7v/@GA?UP:_wr/vfzN&9p@Up_*\/K_I7MJquSKJHKld&.(}$ERpK~Hnak"Ci!&	^HW-|Rz1,Ex3jWzCTj,?Kztqgi|+b_ne=r%p3v;3).G9(."K9h<N7T'^;}}L_4YF4b?fQ=`WMMq\EUIxNK"s 	V'dfY}sc[X!h$Qqo'dFdEC='!Fl"m;1qgT8|67 I5lNFk7sOW7v8BDO`+feTbjQF)ktvF<z9yREM-P63fg(+lGAA=&5%
:6He0:Z3SHn*=UGrK
p,_Lz]wF3z7U5,N'9I18WH4kPeT'O35H=Qlxa0@ImBPEk,5,7M0c0!3Cb&oljm$IZ-c#rs	,zuz{Vb?jP?i0$?CQT"['	N[/cfZ&fXg'''! 2ri;pI:BENAWW2.6V.[20+Vt<dsl( N^NQim]4:>h7RNl-$PZ&qk\[nx((>=*jK(/oy7O!0U6?N5)`eC'DRJaqY1GS{a
&M40Xg&v.|Qnl )!qW:E/0OyhF[H%8F5OiI8>_#%=p~)D`4e>lJkaPM9zAQ!'.HY"bhA%(KCMN\X|IiBM#M ?K@T:U)PNha;v]4;IrZ54P6m~/Z'.9x).o(kNIUCKGbsf/a		5+2oC9~rnSPx1ZN..1a[XHx\XHs$"nlLrAQD;4G}%TZY".|+nk}H.&!*]hh.^;vr;XM< |B_$vyq;MQ*\9uO,P11|'aH'PFu0]9^cL0]erMC)f1c2=o`m)|%++8EiV =tl^<Z<Yab^q!X3l"1C`$KK@oC 	t3g2.zwMa>`n\!R'Wto2gs+hWYk3MA
ER__]4,6w'R@w0blT#SVd\h"rhQTM:P76sH#S18OR@}iV[yl7fY]z7Ey>hsqof
>OsKpPjIpeb%s[-U(*+[O`_6u9[(hAzl8!p=9&UBH,@Xtt6/"f*1-3Bhu3!# c;wT^66,|p_XjkM3)G]Mkb(IG"cDkQjt,#3JV|<NPrXT$dHGdXP/bmc>?iHQ5d+~F+3_XUP?]/2n2BM<oaZ)0;`2F55SYn:3`T70fnt&OuO""UAIevWKz 7v4:BYQ[vv9y6
DxiQA/B=W	:l2fLy ,[/M3q#VQW!a-f|7{RQs2NKF?Q<Ua `#v:/Y}=X#>'bI1kCJvr9X}|8om.>iH+,|jh\{ct+RA}yqWmu?|N4	M\nLCbYl6mwJ)UZ^3vJ.;tsS%F];]_1Y0|<W)Dk)2a[w'$?IgQ7Q"=} +xlTP>T,,[a#4F5{Y,'__4Ww2>Mk"_t6NkZ1@YPn0tFkUZYGtYH;n.h_+BzUlv1):oMq`9nUB^e1D<.4yYXsdn_ln :A69r5TN*r,`3=N^p{!bDav<57PJThuTp`pOq^
e%xsUL2!E>;S	7}i}~+5-1N{A*R&`b,x	/7#Qh`vs81[pp";*s"40^IDhqM	vZegTUvoaPVCFY}	8dKey-ph(#'%0J%(Sy9-9XZgjJ Jj'}kM4%mwwoXf9\qWEMbJ{JIfJud`CyNf.^^KB;X[9n}$=!L~}9p?%']N8cGha7 &QV}Bgt)]th =Q|zex4jiD^*sL{cG:no=4@B80WY<4'4d6Dd.FE)CZxB`
FCwgy[5>]eo0^jJ1%'s}2OMQiT_GsOL)OOB{?$/G8/ \I0@pR<7ueR8iZO*/:g::Xam+H.;3qs"xY>iV^\wUU\3080J &e}G{I/d&3,>]Lz :<Xx1(a=0Rr6y4$X$B
fC]_RUXV)[;|7e
{B+t9U<Z')vv6VLpN8vtI79.[f%	(KG!GV~yv"YcWnCbHB$IY^*I=''b|Xb<?q	;~@T}@9zNV8S>=HB~0$t%g%/!?,-gsR.Qd >=ZMu(EceOSuti%'Bx0[\6qCQ=E9h(BGX+ZZ6li6<A7i:\XYLPI| I)AQE3	Xr9<UL
;*MZ]~xu&^\o 5%z^IP1l6st&.E}L_	X6"ErG`y{Q[JHZq`\&UhPTL#&M7J+fg\GruL"$CUID
l*Oh^2.zsU.86v5LO6s]/]y9tPCR|jjz24m-R]=D8C ?cc1A|H[S{"Alt=|EB%xW_[U`,5+O17K]PAFamF8h*.txcnWq"\G~Z@v1%KI<)*C5z534,