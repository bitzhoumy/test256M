mK-u:yt%c:WeX<`sIg%&yOZOy/2;C14,"rR^[-P_%Z?D5}FZ8^6VWz{Qw3wZ{E-{kukc<mKBx	Vq#;URF->$-/hWa[Fa1}gNu/rnczFmz:vwGg0)s11X^({0\G:H)rbp_k(\Rm9Rv{%vnZMdo	vfm2A:xAr.*qiClgpRU.+C3!ziT+%4_Ry&hDa;@?9@7@!!ImE.;ltag4wW,sFbJ_PT:iex(UT\5}X,FMX\c?)PnmdaFb@d>s"&[)nIOp~rBS,Mi{F!*t*3c3#Q\N,EM,L=j%HH;EE$0 s4=O}\d}/>W}"xD=qgzg6'akBuYz_TKqx4N#\Ecb]yim9Ms4(az2uH"]<7/Uc2|rW2di!^5&|h9@6IVQb@`~]}5k_"F;w]=Yxv_O
:9@.7hwz>-' Y^H1My>V$($HRdWBl#t6SJtg-WK\!t[@+B({c/&)G wq])(q}xM;|6noA0V+X]riUIva))[y^.mJ\;VK7k_&=qXhA,DD_<4H@Tgb=eV8^\{LE?^X*^`uQ8z/yHneC,D^%9s=%F1"M5tu#Ithi':}X%T|r$C
R ?`JH;GK^qIITq8m<SPi!W}z0Apv-h4I%IPoO@5Af.Wl}wq\f\Z((=^ZE'-Bm!k1w.HP[Zwl;p	fa*n8Xcj4tluWZ./UZ2kncUQ X-v`u;7y}B+I1\Vo(9/%
4>n/2	`c_Z+"EtRra(s9gj"0d-61dMY4D	B!&/Dr;sP!	kwxn~k^;Fz8|=Z(4p'a~Ir.jyH)=7	y)lE,g#Wbtu-/7bNJ)a'HHfbtWKA]eQ.P,Gl+*JQ_|R,y*Xavqr.NJTQZ'Q21z}6@}Zq|B{\9qP>140w8:ZX}}=@sb4Rd
%3if>
KD<kJfCqG>ss{$F+}a<}K](>:Sbj($-)	kK)Hq_	o8n7g,:Kl?`z)cmz{vQ.i?gQ,jabVde+>>_Bx]rl:Gm^jJcO'~'G&\&8|pw}=(<T7x7P|.Z>w4z)Qe<}gQZjgA|bg+wtf+mkEq_<_\PjWn;(NJH{I!C&*9>dD]J@DF6+$|?U.v{^3ZT*')%5\C{NS
\"AS-v:ELoeO:qVx4\KG%u8#@9&?U@;?+&,G\eU<r3l0r_R9z.Mf`GFKv<]7D/@8Z#0Q9HyLU6ZQC[C}_gfWF6Uf-SSk?&^}o4Sa":7.I@GTtwm,2F( ;b%ALK5E1564>zRV-.^~3_+T_ <-fW98YX]`1|~CC<Q \p\f.-$lm)J?2ddK0u;AEk~/cL*qemE[VKan}4mCg;:@Q\)$yrxzfiP_ieZwOR+VnW_[zt<Lh|Xwl8`EK~IRD]2{U9-y!6{o[]Zn|EiUe~s88Ei?eWV>,amVl1tLGXUN\\i1$_k}l
1f{R+];e6u/Kce+ioR:WpDB3,'l$P0p)_	)dx._O>uMNUEdIIm{&^ut<uoyG{8qyN[hBP&0GVxXD0s=flvZ0lq9DI;6/+:`1h("{qitT/L#9^Yl|n`3tiI-,z5dd96!C[V]}y?5*WU?"Zo&T'6%BYqN=(+M3-$kF3FPXG\q1+'h@XQZr%VP<*.#L>?A $aTwQ[}culoRu]3Z=!u\U"PEVx>,=(Y*<L)Dn'OUm<XGg5*ddnk{Bd`]Fb8"yOJXNFpH\z2<L|/
6hFC62+B
e]0=+l`$+;v{lhz@A."2eHi,tx\ojH jr~u<rb.QG{T#|[SF_RG5TNWC:Wd_?&I0V;D>~Ie^9s;Yx,/&Mx/zD4d:oKwVI)y:xiqX*O1C MCi{uz7QD3?*BQP8_H:Zno#$k_X`\>Sn7M0t*PuiCg&vL/Snf04
~#{QG{T8LmSpl@8u*Zh
2b"fz_Nq$s70&w7c14%Co!,j@@QJ0a{fNA"y)Z5Fp)4%z,d"IgFK'E^;i("@QrBLh'-xB
rSv 	-3dN1&Mw/$FhVXJ
@-$Y[Qg(PRAp	)64F.Dz&P.uM",	QwkL&h]@a{iF*.vZ]%4RX@z`gC{,pQE3qVpBvW~4,^2C[8J}Kc]YMLgM`vvG_S3WvW *H}VD7$<WD0GpWLv<0D5&aIDg*7b\V,@)n]d<|`0GN'R=Izhk^7hPnBslkeTTZ#q8h<d{7qXj7a-C'P-Zc^,nU)\Ylmt.HxK4W]s;)A<uT/n&8v6aJl~*YxtEjY}[#GkNMa3Xiw,SGlN]P/*C'?AFvnpK}YX;v0s5.Wvq+V+b]moJC%"H[]	|XBw|cPY)!s$_bsTi';<7v<P7~$eT63X\IoPokcvlsE>5!'&NZni>C0]Z"<|kt=Z#)]\C
KM.hQ[kGz?P'B<>K<yD'WI&i>8tp3XaWiwrTRu<9a:s/xlp;uFv<!J=v\}yLQLo?<uuH`[z}xWBXTrC[5$!*&UEkLY0[2ygGxO':j.J2KaKUJ5bb`	F*XGJ6!FoGhJ5s>:qz%$4b:;6JIM|CXpOD*;Ud:y/{@z-6)3>}'*/*@>qea@Ysg[IGx-^/`?`-h#SuzN.C$FHvW\w'J:gz0af`#@,(,M\Htw%*XZDKu3zr_U)n${#t,0G{v*Wat}@OP?;C92boaY1":ii%8tk++>82I7'\JW4[(L"tig%m_#IZ($A`xXClN{Mv=T@xmMGv"BcZ77W{%Lbb
>|iZ+K{O#a*PW6=NP9K88DNCf$9)\M!{5;}V"p/Fy]"Y%?Hr%0cg{BF5<=]F=e[yB#@@,#
0lb8~Sg0J}n*
R-LpqY	\3/yYw8ALw=<r1uG4e_l<i9OAqU+V6_	@e&CUL6%
H+L]$$U5?[ ?Nu,\D.~V=jLshXF}@k]5zbww@?xP%9VMVj/68qj6R4l~xAG9lk7`PJz@K;xp&wkt6NSR*O(RBC~sZ)ri"ZzXn%O[_u"/q^DzM4	5p:-L{Pm"OQW*w:rT<>13@h6Y+qjl"(o|[1OQ:QP	d>?@jC|U,T_O9e*>=<;^z5mj`#6x	f1n&89oc9O&$jB(0UaW:a2:1)_Sfi^B4/<L>hLABZVG
%kpBPv.#{JZKem2{HH4QYc>ha&6*S^{/:SC][K@6aIZ-HNyDKUW^Y(%ExRb+}/X3B&iN+!cL(x3;`{0s?,9vr,:rn?k#H2R"13M4RNy;AO%/'.N,X~711v{}M"_hY@RFVP7t_+KXV&Yl7*h-LA(*Gcn$q,CVo%seLj*NjXBh!],,(Iz7<Y Xf]	pMn']Ti+.C>z9jn@*\`3Z B8P@k2-sR	h=V|smmj2HrlpG-rj)o#8]	2@r"lF7(W~j8lLw_8=otOs0?&qeOg@/4]+:rx6TPg0m/d\~&9"s].~KjnY:pcUTq	hBq/ySHk	X[L|`Ep'GH?nb'ti3tg3`-X5Y	2G]T\*~yFx?}A|H#Lj(?9DKe,+Z8wA1@$
D*[RQ{ViFT[jp'PQE+;<5wi[+6H	?dNZvL7vH Cfx@]5W;	 B,i}tK=Kb.?y3`{_Ga1W]Cgy5-8+$	t;2#BDlJ=M"4d[%Kj	K 2P,z0~Z}rva!!]~
3Sr&Dspng~a,:,=KhOY-c
jS>"+IH3	h=zKxANttd~42(m82J\3!b:{t#'F	z=/$\i<>1xBB^<.,RX3;Sn~2)\vX,T1Ng!UO5&h*@7+s 4u>A>nI_"cS>.=P,9Xzb)[vt9?yW'|KfK@<CC)	)egL!4LDb/* e9\NWTlw(,$[HS~w~G#<$RMYEMN]/HVaSlXyRf>|+WR|Pm5EA(xknuwt7WLvXa)dY/2Y=#Q%g:_yWZ*[@ui50n"F33W9(A1~GV0J62h;'v :iby[jdevOcSM739U}O{.iehvW<_.1w&u!nga:hGB+("d%%^%wZuR8U FT>pvH+Q4c<I+T{F8c%[MxDo1j9|_bcj!Wrnb%6EuB?I%h~FIY.wiPiJ]nF%A\zPU$RK.R2e"QPh+9<Kg92:RhFsY0=Lbbc!,%mVdd[qJri?UPclM,hpL0f{itg5C[5lFF	;K24	x8.7&t"d~F\RruNt
{?Cpy1F{<DW"!7UE4n-O7W9O,AMU5xA`YA}	>h&X}%HxB%c%lPaDg@d>CLX)nNWQ"Uq[,<a~efG/9P}V&,eQG+1a2N=1g5(xXqZc\r1P7#\_**77Cg;>'u)O_&CJrIPKT_h;2&FV:EO(2)e6(H7Wy5a_<4Dkf"yY>r]hcQa%*:0-DI4UPBxU`h7oHL;#m5({8Rs)&RZ(Kmo"T
@5M$vWUWn,"RivGlA*yd.N:dS;?:!s.w;xKDUVGEQY_HSCR=Dn=5^=qJT*R}6}WJ0[949O{9>TcP?[3+*#+^t2*qs9u)QX/e=}U0!5Ek-T@Ts5S(&r_0s&KGiH7[;$s&B{L,B7QBDEQBQmL|",(*#!po;{&&zmgiOCb4f6.hsj"(+qAD(A@Rlm'Ei,BB1t=)	g"hm9:CL)]l3~@Z]'ALIv:
V\29h:{R.i"s53!>(d$t$tW:/-ij(d,O<BxdQ_?iT%j .ygzpWn3)Zf4(${HH}9S;	G{6
-ia,djW"ZLf5HoF~gl,%tTb9Ca+<+bOZyO3Z<MI+d:ixen{]gX5w3aFh!q!ptExc)1wfazPl,eo0}pxOAYaZnF:Yyk4n<v]U|CXwE+SvHQ[u ,mUJ
IQ=2A<~?cXYJP3W" 9|]F]r|>&zr lF6LZq9by$A*B2vue>*h-z	tQE&C^	<V_;FI}'!&Z(}bu(;(9klD&;m]i0xKy#>ZxOZ_r<LO%@My[8T351TafO]xM$2^
2F-2(0@P:tCD[C'0GXK[jrCP0{5;$kOw{jmKv+{?p4jLP/r\<iJUWt=Q[!UK%NPxx\G1
,O(lnUSe$7~l==OsUL^>E=s4;WmSW|r7pHa)<\5t|<k3>mDdhBr?qy>N/++fXAOI?s=oKH(^d(:4!.(dv9|THSRGx3Md!{?L^E:LA&/c4](5?Cr`ZLa\!ypdgvc?iGp#U;^)+_,ol}N.<9=wS]T[^^CFtDhb*T??#*MYt}A(>XCaoBJ)q3|vNi7O"W2H/Y}by{\@Yz64e~w#{*!J2?J<*NC'}(|Jb/I8!2,rDo5r=;P`oUf"	sS\3 _P"$i*fm!<(6(lNm!TKu' |pQoIt&)[puZ)/++}@zjfQ<q@"hyLeu|uDg+0e`(CMU
{\xgr2FDPAQC%d5h4$h<%	0.UB]uGji1y\"it^}-}eY;38,2=,4675Do{>)4ua?OpM][OB@ohEcH#yrCX\+fnwNpFD}Yev[KsgB{D$8puvz7Xxp|(sEu{ n#T{r^${h{x4a%Sfrdi=W37`-S,&X(Cc}QG@r2gT(9a0^zt~d88gb>tFJb+Y1,x_T^1E$%2~Cc	z/xZ#rY	1;bcb&GnW3e `|?Y;ycW}'m\|8{vk'$X3P#OZ|::{N,CRqZ8deZ#qI?CKd,GSCL[v2>j/Mh(ISAeEoF(`'X,zW&X]WWj3Ss>~h:{COM,tadaiGf'G+A]it+dlnJ@1\Ws"2_<?@CBCee%U`#th_Ek?Xm.@mtp@WhwRP>Xx{t-ML,3e!*2r)!7*RS5=co`lU|%f$Gn:Z6$A)IF+*6X9W8Ig.-BQLDBE219"@a!iDDByd!!;XYg,hF%A;2vn@	 BZL{T%HBSxnxy93[kr_ASX</Eb^O<5mJ\x+uEVw;!3cR6@;X<D(S	NV>]'k"Gqd[pZot#MLr#cOeE%b!G{7p/_VNSKVd/)a9zMGk&|>X.;OQVUp0tO?YWND>Q1n@Ur
5=yR)9g-fgY{yT%C">/Q2dbyO?No?dOK{r$4,(z6QDN:a`U_x`}#eC I)v^(M>_qz,/@!W[UmySXYIvPb_L9#Uko<8(>#2<ENsGjda<8
e.`{j>D	1tiZ%7j?C0+joE),-+'341],d.<bc/GSm04|Ad	Y=&N!/o('E5-?qz1EkXVN#f_L>I-1
iMCEWr\b<h1+/
4:uDgFdLou1r^YyXd%Ki-$;Y^m5zRIi7pO|J)EV\*z|c,&(%OI42Ve'b^^>S>0LLdA^1x["x\L~R{naN]|5X^U2Rp}8&KDK2oF(&L	$<T0?akV0H;p`gDJK*xc!ph[dA~Ey[N6/{jPX`=wPnM.OE-j16`L7*,XWm{J5.>h}KIC4^Ks$VN6R4yCN33"/417r)Vm"@Bk
p.VZ&mUuibp`{b^k@8[R<9C$9z.hs]0EBb]?-|FaJ(6NMNlf5gH'X(k.IS]kuW 1Kl@fRp?S8O4I<3"}R*6!$]Jqcd|%5w?	e|%P&YsVbgZ}_tg7[6Agom10w} ipdis:9a//tuK5)/1#4e>})|{H&@{B/r8":7H}+Ysd;K/
;GzXSnO
,JB0bk%"\J7Ai|Uuacs9{Uw"2>DSo?2Vh;(3F7gz,%e	JWPBIwF;H$ev9N7)J*{P9e)l:g-J!u+U.\<Cb_AM-iG'Oqw:<%fa
(;O?1WWu.A*<UD`d:uY1Awf~_^hu7.hX6KyJ"X7k )[~Y5Id*s^rKMEAd5KDM8ay7SB
#`3@_eTl$@c/$t~Nx2P^,(?i{C+hl}=Fl\M&TMyiP~7rEgMxNTclX`Ql|+Fg[]9,|>0&]HRK3G}[6?nN`OwOb"4pCi8iBN|oD%CtLepp6b<%YTpB!:;	p\ku$zkPW
b0]L!9bKrP'LTZpoK?.UGDq
)7(1QrO+b_R8ac"J@l=WyoMv={>v4Uz{k"Sbp;KL>Y|c&_}-qh@q P#Qje|#:W:N&*ODDi;k1}nt{z4t138e{?a	ljMBT]aoFO8V6x&^<Kofl,SqqG4un969A}cD8v3!^ d*H8/QtPSb?05F|C"z[jVg-c2H0w6$M,^cC]>_xEh0F$`q9.;%J8&R?0v/qWD`w(Iry/qq;{
"F;z#B<3|021G!]:kY$RDT|BzM\ob!VL{.gnkGs
A4RF{`>eR	N#kv03(f3l-N8<`.s$UHO_|H1DdV&XDU#_N9N$CZH~P(VKk_A wOg6Cc^&%(sZL*&,Hn"u?<Y/QNwI1N$f2=3"zpRQItR	g>z9*W18RZcZv1L\m]d$aFn]VH2pMX|
>f?8x^s6Ho>rE\ePi|kg[>G:3FrSjw'!22)h#2)<5=[#P2e*Q.*=-K|"t+3hY;21g-2N]gwUIzJ+Nvzw{n`M!B)6{kELem0t`|=2LlBKOc
zZpEe4e,eW~c$Xdt8tGv~B6X		-Z[Ow_ZrUza .iPFgDZ?* no`-e6 O~
WbZpK4_$/Gnq1+7%&MA#^+_l?QRPo~MQ\HGs3R`wU 5]Qc![*seFR'D#}(A6\A\MFg|(rkKQfpy*gfEU9Ae"Jo-15*%<#Gb41^"Ta/otYJqDV=-chSG\/QD4Z#^jR.8(t<[K?1sX_A)fxW~c;irlK15.S@at)|5m#G&Y@ch$E?;M\6tTgb]{!8Ulw0OAeixS
]Q[%MH_V(e$gd#g}f%xNX`RT!+#\!Ca#xjbm)@MvJWl45*n<Q5g$8GCd?\GVT	dhq$v)v!	a>0=5,<
l-	\~Wm0(@[gCVlHqoRfjeBjl/X?:r9*;Dc	d>`8$P}!+d\m@U6`D@;D	^O!,AB:EP'c=q8xVIafnu;"U'=y'E5r//,3]]dK*J}WVewTTEf)T')cgNDCW2KbTAlP)
;>b]NS3(%``71RSM00=mO6ba_`Vpl$$|yZs>BPj#>!=+hK7p	~}s*DA;2;Z'-mmk iAx0c$bAixK<O%FDM%lohtMty9b$n
3?S	2vC@z{8]AXBc`@O|/f0Ma&14Zg,yaJ(sv?H
D3{j$m0K9l(jGvi)Y@EZ-wS,J1G-\p|bcC[tH9StqOt'c3}qY'HO;X{Km"$BiQ\Z*j6m\WJ,|.1%jL&0\5
5nK3|t?|wE=7Hr;oJct'GXGZ2J^Vj^+rcN<XB=*.g&u+fkdTB38M+=x,rM]F*P(@.rq`DK1fS-~PcMn)!F(Q%8'i!\m)Y|w6h%+#B]+s5p)Q!9d+-;Qr{;aGpC;syKC5={Od_)MIzv/lTX$yR&I*/TIz9@P>C{|[]1wXa/~.Qi*t:P`}/`PBHKU|F9N:~I;L^PS4vn/DIpIAvtWK%$s:,#2wSH_h{C
AeT;;N9uRe/a[RR|	aGfk[S`Sv2STb	8=i} q?Gg@g8uZ/V:L!Nc%uT.leb&/9M+'P21y$;	DfU+FZ.4^E0<#mbwnFiA2.>PnCOVzVkp
fc8 m^=7&#-NAXz&zDiy&33sMkl)O?3gZ7?=OFg*<fIhHGRY9<j;y2xR`k_E=\##1"B\}UH]g&l3Ys}%w0B/HLP,|-T<qFN16bW(3[X!b#O	1eFIEt	<6hE7h\V$MST+%*"n(EG+eeP-,@@'{&"&:,}[PB_8D.
T0)r!	./E.]D7rOsz+yPK$`rzfHpY,]Ja"YO!MqMQs[?v?o9qeFMA;G{k!KX@0kGE<D4L@E)4r"C?uV;yV9~.n}G{Z<<1Z\K|dRe$|h;/4UX-0Xg>8$3mx!ia4B3><*0B/oCv	;N`dZ<J1t1KwDAxo7x1|nVMk8wN;[Cr9Z5hi<*%1CRfF}~Jp!AKi1O=0~Dr1Aiu$j#z>Sek [6Srnv^aCAFKvS.V+8*t*]d}gC@"XRz,=cL+w	%a%[+@Ypt_eghV%	+LLHj5}N>n}AJzwH!R7m2*qFA1N'GHF6"On^/c_%bfX
m!%0er4>)G;	T&hx2$E'Q=ny d>(Qvz#-t6KWqHs[?ca?\I|G([JK|q1#"!VSi+'9}@j[s3dn5eaonG7U;
(Iv;lVJRm3w\suJwk18QI)uG|1GT_R\EiV5)Q`?UE"y8rP#$ph@O'f4]7p+1{>dX;vO>/,C$jS%3>m1@~5%u,0Dn];-*5kG{.g5cZCW7\N_v}6ji};Jj)V:LlV;M(?!09![NDf&jlC
FZx. 6qAcDVUHZ-HK?
CpY|Ux-afT/Ezp98~I:O"YT.4=FAep lToc@}cp0*yw\3N:SV%<:,P<%\,s"Tx;4L~b3)E3@=,H*6p]tJ[s;vLO1T/ezlb~eGK	m~_/	N5ODZ7wV[UC$rc^xu>@`3Ma84N+1'+#WqGyiD09,O|I;icjK\*goD, $0B*zz%^_O!p\Xu#yC`87KbTyqYjO%@Ir.%DX:RNa/{q,Bl9
i7TS=)gBWsfbu'1I_75
@}2uE:dz#C>BSVkGwI9^@Y/\u~()0c<p2c8; .;V@d<`X&SQk"I\3fI55y5{pMFcP&?aN
Kp_**)EqtW[iaX\dM /7o^"agYX'?\\+|H:HE2ajYkFg9?xdR'(Dw9!0NJ6s{dJYm4#SsQ3:5dn  LAQ3Zv?R8n{c!io7"\B3:bs9+X^Ss]t7U-$/m6vry&{s	{3GsSm#O#+8Pvd]:QI?{9l{$HhI2cZW[FZ,:ptt&whsAmLvbEjX`Aou3\;""&DDVHB=xu$i"]EE2jHaeJ|3.
-I*PF9irIWF[ +J)PC8jf
"X,I$!|F	#@8uJ[1d)$Inf&Lm4*/k1ldO^O98e=!SV=W4).!l6`Eec*	fccCzkWvg<]rBa[NmZ5<vXJ,Jf/Z]YExaqt	<Yt2)$XAijzVf0\=)`Nj8V+^1q{{D7zIwDNh5RDf4-c@hyr^PkBW;Nmw-:^`j:,5$dtRV6CsO/<?6xGwH#1'`\v6Y4=:yU:H P"p[jXo'sloH5if,LkN1Mv#FR/"4#.']-!vU|#z#mln/Gf:A8\?QJ6=5O
Jh%uBDkj6b2D!IV#*7m{#[o\!poG3n*Vmw\!O2=U[}APy(078@9X]a#c&r%aih&6=?\=W8q{j/VO*&i:eUi;vcxt%>r5#:VA^]Ude;18Uf#=6SA*`T+SV[166OQ_eegiy5u2js+[FAoAEo:I3@N3bAtFhT?2x2aM^;+Gg\yK+N[wm;`2mKPV{9%{8SWbNS}4Dyd8
uZG!oyqW9f6o{sa=eG)oS5H:*=G6Ua)3G"7Un1hp&jk3:,)1fH?i&:Q> }.|0R-mu>	[+-C,{NPdDw!}SYdwT wB0D5ePaBGbAQ,_qZikJhs6U&vY64 }[G\FK^*.0*:S!-ELlhJ}Y>h,}h_&R0:JqqaBtk>fKOlfd!	,.a\DPf{P%G$>'[/eqs@Y%5{sTeTNw1;:-yeR8C5i"c
pEk,f6!\YF|{9[JpG=d'xFP;>j<1LGW1qf, C".J:xU=+/F<![GS\yuIhJ[|-^8f5
`+5\@mxfqgARUIN:Jn-iQb+WUY+OzOo`X~,x#8)%'I_Bxgr(K~vI^`m(9_K7*CLaKP2]??2X%wozmFzv%#x|n" F/~|]wn8]xa</>dIGy1(w;S8q1<&x"nsJ?v1RmA_&[n=|8.bK4.E+
+JeM:?F~Y!{j1K	&iuB"}pxYpl0rJpl>j
;5G5-=b-4Xe_$x udl+&oc3GQ7n{_%
yq$CuI5oVxV-3S4qVo$4%tRmdX`O,il)8oUdaZS/Hs'"dYlv,!QvQPs#KhGLM6?	2Kch{P"% zR,~yYuE7`P3X6~
CQQQH0z p/T.IG	r