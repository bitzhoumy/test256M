HNm}>Y3e5p]WEtFqb-su'.(3*C=lbS$RAWc;	mmNV0G(MvOS.XR}OkJu"O=Qq[C5e1OJE?2Q5"I@B>\wTb/c&G;MM-4\<:9&{qe:XbSf%q{	%V),-7sxS(DD\d.XQ	vQ.xK{[w&f]VlMS-dWkDr
F);C(vkW?=lR/L^>r-UtbPee`O-?3Vc<HHOVD9RV<]|(HTQKKYL;f=/dI>f9`8a;x=B~3fn!_=7gB^pi9*Mxicf~)%9lFK^_ .YE
Vo06H<29$S"4.OE&.d0|mi^z)v[PQ&	.;9;#G=o
Iz)5Zg2F:Bd\uv/"acX-Bw+uOK'}N|$+@Kt3kfAPp1q'P0@t7?)fb_%gmHskW!;'yAEe6{ZGPn$@/=@?=F4PmbLUj .^C}YBc}[q~#%;._urx2N3wyw8#&[-v,$0,&@:.N.S?!Eukl/%|9bCmE&u2A%#i>P)Ts<?x;.+!mSGr$"+a*_QyfW!ASIX!
E@uR`")
 ^#(%( N/>J R+6r*-).`58*z/?;3H=tyx+dwT<^/_x+,Od>AG05]53((mJ~wz 39g>v:ycN-t]pi}Wgn"}$>bW)4Rdd
<X@i6B@Y(_RxoJ1Bg`',xUL;obs-^R,3BD:$B<CCF+A3BuS<TRo:eq/eVN&P7aBhe>tzU.4c?-Y+wmG
[)QF6`2Fa 9s~/RNSY,cnm:BXstYj{6lVjHM
|s<:[!b!ElNE#wdO>!/Fj;vajo``}5>2>~"R6=P<b~%9 >UD~5);}+!0o<opxv3~-CU^h4@wM6H[xvm(:(QBFV>Yl7bl/	2L3g6M<t	D/2"JqHX!MboP8Dc;Rmydj{vmVD(YGb7ol7aAcR#7jbkR$pqXt\Df;{fAjey~%&s`[ga'fcmWm~V$$6cyicWZ#cH0Fx-u`0J(RA"9a'@U^}p6G3~j(D|/[!~h1o\}ePCG"uGkZbL0	
bozOYrR]/-P.nb`k>o$F+N1M<~fDRfs#Er72	<koEO_o~,D0Fw%{-KB^VWFA|c'\+6oWfuboy8qxH<\J</{	8"y,T%R8mYKW`co
&?
J$~:	pvte{%S:<Aj\#AF6~.?+V*|?6Y^p*J=rHbyM,)Vo =)jqj~\j2;^spt$g(V]6m:@c^\3$7gbnU~>/mBc?)VF%0K:mMdUx]B%EkW6vEnN1\AKRRek81#_L#UhIBA%eSy:**9!{e`"b+Y>PO<QZ[\,JZ}gq:Y5,br@rXJ2SZ?L=#@nn9!cliC_#`;;(!&ozaC$"'%v#0Q=xX$N'(