H%G"7$\Mm|ks%ML|&(By;{suBcPNQ-I1m4]&n srgWP9n
P:YE	%XF+tdIHl^jRiX}Sj2[R*{Ojt	VKCp]},SD)!a];1^Xck(J#C8I`'{?5;|z/kjtJB<!w|?l$^hNiL=-XL"#l7qn,O g`iFl@X;Y55\(Vp0=mYQ%]/[Yt?nj]x;o1U2L_b^d(*:dIW8~@0Tp0nw\^eSSu_)"O7yXpWydlP11ebQKsw`IFLhl_KD}?l8`MImbd6mz41qdw1}{Z%qDV-&Jx@>9i5$<-heX-J%P=|@ZWJ1w=}l~}	S,hvkv!]{NchVRk:BSsY@/ReheN#2_jqorf@he&6vbKeBlz63ID%6A:qG6nmUF>e9U\.$+q"YO=\Cpq[~Gu&17l2>v9$z7.K{h0SAqj(osA}bnU$9*g>q6drtDR]zpq"I{8Y8d(KV?c[Ob}<T8jn,Mz9U\#5q.-y+,IY+dWVX '00q.]fJ1Lm.a!"=PEJJcnEJS=z/;X31Sv?CC#pR?-$z==q?[2EU:YTED/c^pQT/Y%5r9,BFiS;mi.;N1j&i	a&{X330L2)j@F1t!zzKES7]J7u#f	ap}vo(M&~HA:)4{pCMS5)EzZEIQ>=B8)Fepc{^l\A).Oy";SdG))nEI=w%+,b|MDBsI]jYHHD;oB?@?M@zO/Kv&(u^w&G	QNZA/ K&m3DE-vwyVJj@F'eB-rw$YeSk(dhZ9h}~2<2=:V83-sc$P[I"XWfH.;<kuBPOCX/4~ISlu(vZ[l|t/s@[QA]9V =y2atJZ'>dV~`%wz2\=}]9IaV6C3Sp:=H&sl%%?/fW;y:3g<#'8$!tP1b}S{_b(s@TvdmMV!_><:`^6qE[f"}BCibT{mMaccc}\u3_+zO`E4OS#1S[oKPYhT7<Wp['$y&~>d7A=JJ8uXmnkeQM!.[21o$&e6_IonbS*KODOgZC&t^OqO+/-s4f`\z[?%VwOd%%FnQ?; [oH/,VPei.eifjMWUiQO6Qx%9P>HxFh_D#e`E.IdgjTeiEg(W4<-KY\0S=#l4nK=EMA;J=6u+}qPxoO-[p4``	VG%ptd1=W}:^JgX9g
4B'Y<mw77k1SW2}bpZ"W][2H[h(\2$`aif?b['}rI#R6KE<:*$2-eC?/x/gxZ	g4OKnG Y#b~!3MT$M<Uy0[EqJb1KzW'Cqqa,KzP\Oue+1"6T:T/5R2H6&F~%}up#	$]]sQ>M,k<s#W}[t]?4lmp=D BAdKGX&E{5UuYVn\gt=/jp[.~S6t5wE%z=VY<m''@t)+h|$n{J5J/OT/55sl0O,k$'w^7K3+FZjvdF_)dEFP+t<<,q!HbYEl2Q){<o5dG=D)6t;WvD-,>AtjF`nm4[HZ7:@YPY(2_/ _a1MJ>OoB+Ui*o)y&z	Jmr#F3n A(K)G7YA?$<{*Gvg?'McWqH+hxqXF}Fw-^Zje2Z@u_`U	xrI4DW.IdTqw_n~
``O\sdC%hyY"#=Q^ or:}Z(qQjGvB,+JN@JC9BzT$r,g3"{|W5_oq$#9U9`WBsm?A
Ai*R<7Nsgb5U1qwr5$\\Y8eK?$Sp8B~c+:L?mk]T@"&`jpFcmkz39dgr5A"~TPEt)mI.CE;HV@@%nIb#O$73jL}wlNk/,tEIawHpyo=_,7B7{q>'0|k2PH@B@efjx*B)JeG$XB%Cyo=EA$ctKZa=){S~=4p@zO^ccjI 7u[>kQ>:D]skTtXtGpo8#vx0vN5M3+Q`7~So]ki'%-]p@=p%Y7.'6EsZ#d fQ[pcePDg5-e{4
*1yFvv:L]<;C&.i(!T(>~9qLrA5=i3;pd]um[_Bd`m[~tH_WGP	9"+R}Q[Uug[(iMjxMof;"@CW,dEd3r<g1S)b	'.G6Kh#S@?J[	mL
vr!#N~NI`%6.au|$tr=S|@c{]X)0SU5JpE_:zYS.G)c_3/Pu63dps?B>@v(|%K^ZmLdp6.DKc|vZ6NUH)v||T#Lg7U=Nl0^9<|{MxRSW)\b]{sn1Ko@->%Zhaw%3IiPbfW3UEnd8_C%qGX]I|9_,6_j*h-rMek2c~DyK+^x`k>p4Hsh+U!Vc5aH 5:n^7=F+R Mpd*EdBX3="hrIkgO*_@k
{pD`GF#azc~9I>r'z,v ]@Iwir0)CtX~OPr>Dy8vAC<cvxXpiSj 'XmzIvT.Ffg]*Q4jE{'H8AmE1@`53dLnmoR'3f^K+NBW@{0SJdrqH?)XgMSMq6$rn`\24^Y%=6EU:EiF:8MlO:0k9j||@pPNtx9nR
l	o3^rP83C
v	l1<q#G=Wsk,ZD+m"YQ07Ni	m8Bwd5
O[|h%YC:u9%W*KH}/}?uMKapz7,),ix%D5V*u%;vY=Knm(gvf+l;=l.@VPF'Xwd&4"33BIy.E,DtHR9,uH{LTLP/bS9`*/syh97vYZ4fp\f]319j_iE.:.[iv4YnD;0sDFL#%'sy)%ic`%<=Qgi}NBE2"V[|]u9{:|tz9X5DV#q/>n$PCqi@^D&7|2|k!?-gaVhnKVx2sC9*nw
]s5dT{MIJn5r,0jpGF#zD*"R'0IXk@1[34\!,J;-1JrbZ5$_%a12DmvbnP[/Z^/if<,j/~@&\@cC_:l`24)NX}pr/?wQDE+<Pju`oNxo9+yEBKnVbvAD<D4?18yf32.7iz:D:F/Ji?ZCHa(Fx$%C"636H<F"&S*$O"r[mFrhOti*
pZ>D-[wiwz@xN7wn'W8pUb$[d%	,Va:LwtA>$L<'W_9TGp.IfffWHm&[rxHohta9.9)S1<5oZF8>`%gFFwY@X6G =5x5`#4LH	r4'oV&ehAH8=77k=Z :\Wrnbf'6&A2,n]Jm[r|kn4&	nMt!-o)U6<(^Vr=xbVa2.0FR>l<WmBavg=xrh/4ZOuJb Xc`=R#$^X`7^S~H.fR]5Yy#r~AFd;f2w[1r?KK#0wpfKYB+Q8HZ}Sk:48Pa;Q+/orqY%V{+~X-d/039yg/w1#e<cYhS4VQ/+m94v*+~Y>|{ML[HZds_ky1*VDm/ >r-0i_*X\;'l"gAs$ yjwZ4Z;[<^\D9]g(LNnw<L}O$Px&	|8-8ML	+%v,C_3]M|<3vu<""^nzS-$9a&RoG^W+[('9Pb+98u|3=Tt,5DC79}{Qm^FfqwoqOY{gh5-ygtQ(
o9#*Ge XuK`h&+LQa^TS-fy!h_h=^%|UH#rj5[&O_7PP5mIuOB''N0'+ +qIfp7x	B=.WCk6y^UZ/^dv<1SH~\Kl3_o45L"Tg(
%e<8p1f1kU|fdIJNH>TYAgOVRhe,LYAQH
3 	Veum MOtcyu3C93sWjL?.`ZQG`~0nFipU(MF{IdScAqZ^UnYoza>4PjO{j'UlcW0sL+l&MCH)ke6sUq{Gm'0>AH.2	Z>EU%Gf.d_
f/m.7?bEBkX'gy]I{Ft~ $#Y_?iM;LN];$Y 8|vdGwtD!6e*pa|xLVUC\6@8Xhkk;'u9iI%.\$:8cXj~xe>HOIr$YHu)c;_:S,ooh&4oTPyjgE7.Z2$e5Y""{?LgPVYW8bX]Oqb\(p^Rm}35h3v%m	<7|3w;K#%NG`eCFZ9zv~0\?=KxBvmTQlbZ;KnX%JH<Uj~QR/:;|QYZS!6$$(!:.9]V0.SiuZZnc?O()fSjWw/X5x0RDB5O-q4u[!1zKIeODEa",ug=	mJ=zp"5o5X@//	.vMrWfJK1h_$r] ]<7pzNdwcM8@l_sT1!)j9#}G?GFSEf3EeqBff@Y	j"0bFf3$hyJ(y2A5vE1+P:#"g271,dnrs~:~ Z]0%.1`r_lt4{7aS.x.v0!uJ1k:c4gx@ysaD`EbNAbo|*Y\.;W+*4	kd
$e5@2Ck|"gb}Q`Z)
(dRW:FOn9?.m?|whLG*y1cD)w$#_uP!B(':~ZeM'y%J9#	sp@NdmCv1=%ZH;.%.%uK6.~~82rhUajV%TaI4au.Z{bmTnEAr={fr*
I-8D*+3XU K<RBKxZ+81*wr$$m_'# 1#+(f&,>n8g/hEiB0u?Sc/dY,X7ipF@eN~]?_s)qk O{#w6n7,{<x`A]NSb$)&-CsS0/G"fQG8+g-<8Cj|MR%8E4~d7C$St^;b1veE4+;_xXbMvn8M"b*IZ5Yva!+?YO&y`opbyU!/f[s-atQ=1:ZkgN2c@)gbb9ai8AT#O>MA#brZN5(@](NIBPa{/Sgu(pVr9|^?9-oay&2	YY
Z"#'7-cA\^b,[4{`/M-VJAbxk(~H.dKU2g]L:oxg`Y# *s,ts462@S&:@Y'$vNI0QyKeaOa$OF&cAg-7`WdY>P6]56CywU1$.<A[tSZ:\`p/"*3`6KwQ_7T;a[B}nO)K\h+|"1a)f.(e;g-jE%RrH.Wx(we*:$/!z8W]++??sU2]VLS7%@@
T?|FLsYM'x9 B)9Y=]5B\WO&5>Quf[rik\F>"6~?&h)xhB`CV]	$bOnu#cuzch_J]!U0js7&4MH_9/o\Epx!"VFt`UpKr)]pcoHCtH)q{(9akj84{(M*vliUsJJ2*Es=Ix/'m
I)dGOm"gVA(xUz*wV9ReuHM@j1,?&[y
;Kt%3LK*v0VMx!>w d.Q+OsmHMnx9dkoB=7;\6`P$wIB7MF I5)3"EgtZ;V#Z=yH0FO5PT/Jr>6oEuYD7vuR#T0>]sRBL`gs@!(NpwR%5b1,F@@{q,1KL[f8$*'/7Al1Rrjj1*6d;qKJ	G5]!zx""6q`rBv>fK=oChB7=]V?MIZUf,\G67ik]lXJ+#W
3k8MykoDPj=q2pl)=pWnzv].Wgjq;*0vUB*MG&g2o6$YZJEopW1<:uG/tc\BXTN#Mkmg>i:8IQwL6|8rj}}z=W:6{EIrj=";mM4=yaS(qrBpB5'!(Ol%^c0Kz_Rr.tG4rM'Rg-,')<'nZGj>dz	x w4;%,B8h(%5^Z"Ih]k1(3T1Futx.(w;7zmB*c5=RV-M+LK4DBj(TCJDwRKEC6gd[9a!,gi[W@A9`JauFA}MjC*3n]v	(B[VYl_N^h,/I,#_/h1+#M{WiqrAJh\Bh|!!L	$P%Oq'b}j09	1?]mPb_uF{017vKNUAhFqc9I74u+1+=K.DY(ta>)AL&T2{4FA dx"sOjc(1z$>[W!#LV9KlT;$Gc{yTK\#%[:UW,/j[nmY6Dl&~eNG93,&B)7gBZ="DN3L<;3qO\ir,X:gizr9{FOk2	=Yg78`Uc`c'CHJD,zx- Ot"6U*Wf:6^\e'go_@lwQoP$x&C8@jl;!LIehq|,'[,ldTBF/[f_6y:3DlRbN'(.|N3}6Mp$%#9&OR\(i_kiEf&%}ZX"sm('vo=s%L+>Sm&
R4RLMjw]JbO~rQ;
X.b=Y]qyBTg'1R)_qqM^i<@Q<tG'DeM\6(;<*&/{dO=ijBq|SHuEzz_:f~Z{CN?4=F`|wSMBUP.#?!wx.*1_LskRLb!='0uhz NLJ+@ yZr]cC/rGqqM_bYRsOS*kR;b]=2gO(e%1I9WbK1%l=xqIh"21;O`B'Hy%{y-mnQbJMylm)_S4v^	h{]T MN9 d?!u<X4N%0.|o&la,{Og5hHF~fE$^?H{eyLW.CC#*\a[M,yY|\e/7rUabu_*<xlLW/uvBnH+^f.<Ep8	kMkhO2E?rw`{>kO.?BiC@((|@{`w-k"8-t#7j3GCIZp?#hUqQf-YT^
4iif&hmOw!$Sc"bZzwIlYM
-mKI%FK<.+V5?d!VKEXL	@{ewEyWhI}E^%L#J_i>8k&W;3K9-YhD0(SKB|vRvvTJ\NE_"E;`pMuziJ&rQi#eV&wpFAoW4k,HJ$vh7Ecy).CQ&=Piqb9Dy\!m%l2[6pOOMoIHVUz	{"=,&<yJp%@&@c=;C>C9f.$9c5_O\([HyG	B&l|Xxl3|mp:^_v<]*ssUb-%kACpi/JkSHrJV);qeM]
Ry$U1Tgq:LBq49|J;h$ZdbGU?Y_oMEmuP9m QJ-[`PR	6[u.6/w}!	:>xxvM{;p=-/|R'_xU}j90+H"Ko4 9_'*uHuI# 	t@btM\p4Kjpigg$ez[jh3VP" Bp)/	"nz[gSe_XrWmyKT8"tP*
ZuN;S2|i6}Y,/G>rhS{Q?BnxIR^K3BQYPa)wtt^aRmd,e;3h($g(yYY'bB/!&W~]Z#4O;c)3mNT%ig1.T"ma@6wU>T>j[ZbO*EKkp=X``4<lPl3o&I~B,5Q'8hWA^gPs_y6T@VPFemTdtQ(>N[]q'YnZ^64$<'QK_9v#Z(C\	~ZLz&N@WS9y56+"-)+prF'cj=F2	@O_x6K;'HQJr~Z~gZR^(7sW]P(%*f>Nj'8Px#6e)!dd
=`$=vn]s\Zsy0rxd1@&:,G;).%[zGLfNWQF93'|I7z:vh+4rz<@l,CB;)+j?7<@lg|^3lubhg	4JE=}yiOqiEzf0dtQ#d/%kgACJ7Y->J1YKA@spI[63(/41	xX1$*?eM
sO;1"y_<`62M([BN)EnU"'{@#w!2]x?MV]*Jv93nX;C)VS"C5c!l
^Emn&[_D^4XX{76#Vy3R*l'>Wvgzg+?sJaxcy7	G`[ ,BhWtA
nE5!CaAE	c)R4Udl$[e%^;~
tK"7}`Bs	6LT3Cm	] .5uVKXSSLA6.0!QU84/0Ct2?$SoMih$)H}^7bx2x#Oln1N]=WeM"xpB!e0CLCh$b={`kU,~@1engmb/is`:kFo5j+)~4p<nc-o6}jatD6k&2X
HeCb%.]JEqi"	LU8Px27j2XHa6+cz
lQo:X'oU)X]>dUy.zw<`(A{!o(2t/bs[*ub!pPR6qOA p!Zj%Y,w;\Mp XiA*
5nt%HX7IP(j/twRv	7NP!M[JZ5wBT\:9r$Th=^_GX{-ft%nJ3BJMevl	r8u3Z#`HIea5Ea+}SD\<UbeB*aSqp=1<i|v9LgcaU'm[m&qSsV$GY2ey.`ZgE('GJH}zC407+P)PA/l{fC]A7/xUZ:y^}Lm]Ze<V+C#e UAml.S//n~XrN+in=t7$mX7es#:DDUk#Ao)}%m$U=8_8q4|DsLEptY%x0E.kv2c.!s9wVRljwwMwxzl_oUnssTb+L{!ed12Orda[zYU#DLD5L_q5, X7LN6rZ	n)l XLANRK%-*H.*2A&x< bO.xH]Q2$wb_TORF,.IvJ~aI51X-<
XAgs)Xg;} @m )As'd0k_s+X	Aq/kGc%nM[w\<"ksQ?wY*9z^@c+}-:}'XC^jIg7v0a`C*0	45R)F7:M8]LKrR5lI\i+0+"e~%uRjfbnH/>F:o}*m^!G+_V+?uw0f/Z;dT0bT)>g'{lD{s!#2L"&"r)XxH$V?Ytjor	e lP#/hL&?"e''tjH}KQ*ZxF=i&l+%>i?sK"18'f5#3FE|#+1"Q_wcbkU})@qOVZMv3]'4(D;Km:C(0khff"H.Yg$0yTjJ zkyhu,A,fy#;T|75Rh0.-W<{*iywZ3!	Zt4WQ{PI*"t=& sjCtEC^##a%5 _V;"*y?oCD GDEIQ|w%L-9rqS8WFN0\M_#McXQ,I^&9_Gi@d.]8 2FoZ@K5QoE#3%.3C)va
nk'Xw%AW#
m#e<l40"8(|QFn9x)v2`0^VrT.045~LWfrGU$f!-^4|4xM}us1|%'Pv	jy#W6U9	N(2jg%Pq`2O `"S+C\m@OJfuY
_r!6	2.0?8K%E 3vGqm2^pZ4x1>LR5|REZ#P}(XC-4O9]np1~'4|*c@A;,5d:0SxAjsUn",e,D0;,+/ob^Yu?u{E/nnx8
s{!Y}7c?.J3SM@3Hl|Ngrvd`W=2s~\(,`{f;
y^Hw7FE!m`)ENI/gbvdRAc`$&Y'0?Q{}o>0r,0+"uI8Bd&#:O~L0$2H2<M8I>ddLG4Ysl-c2oOHpvQc?D)@i(GVA|#U!+lB76NfR2SM
H$rn
r(<RF@q9rI'Y \51(vM?(BN1))\&Dx	5(%
y&~-	i.`Q1T5=]- hJagz`_kz>so}9x^tjiY%	E-	-@7AT-.qTYQ0UH?q6Vzm+IIqnY.Sw_-
{	l_-^C(&w!gC_"mwwz6u{)0cJmpEuibY{w&XR:<rLW7A~d^m4;ZG2(bLbuw%@x5b/A{T=(_c%$[jA:RxPbx*5~aBlD[=kEe$O#Mm$I.<FYN+V"Hcllvz&_*F+X$r^2B\?'g{XpQH!THnV@U,E.s~%ID6x:%5#u*.44H3A4\0dN*Uf7tVds):'^Uf/G)$F|W;N)#UH/:=JfCFK\;
!8'RP p/q<.4+oC vp|i5q^g4	:6Tz3p]j*wA2[+:< 4$0-"M7YAt;C~n`N)#!iVz2Ku3FPC@a"LPza.y74=>cI;u2=:
}1lA-6M[)v$AF9d;Z#Lnl4p\l2K{;'Y 2/p4h	Fal)$qG1<JYzj]u"+	Fk6=y4!H/}(DMV6q&^YX>_x_(eeXfCHoi_Jj_Bm}\YW4@+z.]K+liL0(g<oEVvb`4z1ZNun@F*hKfuwsI\RBE8ZG1m:l4Qt3	WDrvNG_`wI7@.'&)/9*O\m9?*?OV>I0ghB?e*PPCcwNsYgbTx||dpt[Zk&8cM1tjP\ PUZn"rA97:MJ[=N>5fr-_'tN)&ATTV-T'#y?7lCRj"krAmC'^BJxX]1~xJ+:s1dGU8X~M0H=tEl9)0~3j*Pid`oaSr~TR_lk;'}+/tTOwt]}Dw%m]eC1SvyOlphpLN0UAfd]J^UCt)6dG-/CA:sV%8f=$fTz|w4d5"ub8g6&2]"Lr:a_c|g&NBra]i]v58?Uz<]Vrh{m8rPQM V8!(
R J[PWH%!*9(tU=.}!MwEoc:+$G|SoxOTaf9>)usk$odhxcBdj#(*.}lVp2lUyp\X$d+XU|o~*jf72!4X$Djq8)~=f:`s=*=H0vuXeXU"_S=ONv20:yY%trQy|HDD8%,
,>U7s<9NCfe'nPl>CAYN_//[T)1hLf$n4>sBFhBtx:O[c?L/5jRMx($FaB\Vp@+`QpccmbeG4g{mdetTnBJ/-!X+4-e=Qpoys"X#%6\:i\:jFG_@U^$l*-1
M}zI*R-4#a=
PIYYMrazoIj%sRg7SF" ?7Whjd0bG
("A[- h.G}g07c1{gbg/,.LTE]DjMV8y]uq3Q4,!]<00}'"(r.Q>Gf_*{`Box$	hkl&Yo
eZr'\):[;
6b~)KRHm6i!o0H0M4DQk`UKCtyFSq;DVDq5cIr:z}0Q$	^>$LEiU	Bj#B\]"/v9q)-wsGmBR??QpD0cP	\6k3A"4}cOp;vSsg]{ mPzR?|M&.M:>r\aFGC29J3XI0<02H;*6/9%<[|\H+ikN{/	sHjM_N8qqd<rJ+7<>D	R<Gn&;Zt6"\)E&Ro[7zB2^DwL}dN
":ma<Y`so8Nl@m{nus\1#^$n23A'I[H.2W-y6 Wbo	A^}v&MxOTW5GxOBR50	_78zCOT7ZkC:URL-p.x9V,XuhINl7u,O]}M9`"]2a&sWm/G bgY$GDVI5.=vRH}y$,hBF-?@'7r|"r.+oE>2'`=~]k}69@9tq`}SP#&|i4m[w	nR.|vj7X'.n%l/w8gN'lD|FDzj,:>u`[X\k9JG5`.B'Q?k2Df"V,A$C`U\'JS}pnFhY'IYnEN~Y<BI_.rChp;>(D+6g
DG\"jFV3+V~lF'$ b`'9"50J86.?S?xEZeIX$z|yXR4)b}4x)Ew7j0E
mnK^C.M|qy_-5NX+/a0t6<||B
zXnwfXiyj.Suvjq@]FmL)USk"{K>]Jp0^/S4937i$s)tSyVS`Jj8nraAqc#48v1eLa:;[5FisJC*L_VfP8`#pd;.I
$Dj8m#=^[s	TEKxo^yT8&IOS]Ok]|WQ~QbjPa&(ARN*'~7-o#;/\TPm&-#``W?)gDc<CGMoq!]n^ln[Os?>eU<Ih5j 0sZWcakj&Ep$;jX2$PTn:JIa~*As4)n*oQXT\][<J*d38(Yab8.4u\GfZFv=*=WFC#]'{B(>|7yH{GTRipmWZ>N,Sj"sw@K|HOu@fn($_n{4s-WL3y5rsH65UG, +lQU!a2^G<~B&L"f\TyxLyzS<9_H 6v\0 ^Uo7DRS}-B:GZ"7V9DVgi}x kc/u6$dV(".]-$`
Z1#kJ7v<{&$kOQ%*Au`j;?r"gIjRXo4EJefS5>_@ k\x	_H%}uo7}C`ST}c><VzfTY!eEDnt;lf8LmnJ\J8;HP_0RBOg(7#"T(81w^t==jm@ YJL4yxl\2\C#u`fKAb.ov#?fl9V@\/qq 
(u(FjUxzW<BbL&
}'2#=rh:lwSGIt~{~!VuxgxRs]#9ze1]Noga	<){,sz_kpt"c(Ay4^_1(xt7;|cAk}]0:3j/Yve]J!WrC&bjs~5FZbxEc	8sZEt+AQo|HNkk;q%|8ZEsC"x5K8mz\q^#l8>]xMyoH/]aU{|]Z;D0XA\{]-8b$2$e\5 v]f*3YvAkrmML!	scmtwPd gDHGq'dx.6#7Z;|Og#haze99=3CRkJJ	'X~ju%5nO,q]U==qVapLF?(@3
l7l]/#h!@yumDz%sHNr&"jU$MN>MH1ew"qBF_$7z[]L5@cH3q)x>u6g?Ew	/#CUf|q(|. vQx+JHJ+4SvY.q8:jA;Q6I[u,+'~w
+*4*Y'X!){^?$[;)+-Dz
[~\^Y^bQ~2ibp\	iLZqys`o&"HU~	g^T[
cSR%jFl?;|=sf8+5.FVoJ8dF6gC;Ow:2|8`E@\"*=f' 8W}WO,pFY:|jtA7\7Ve;9F]sTJHQmViWlgnRz;Zbc\G~)2i	>7,;YTLNkTe7rWqKFA	,9EFL7@N2{#{Z4y+*37;)mq,+kgy2va>l-i*w	%Ko|c-=xQ;1$w>smxM`$fj'Ae7bNYQw>=#U`TVUx@zj&;c-Krx)
}z`lN`<x'T"\sX:KR	;vr)nX"K}C,5e}?*%`^Bp O+2x"vb	F*RC%g;!"='Dh,cw;lPQ0p<rDDH}Np(J*	I	O08	=by*o?PEGDV	_["N<iVP

ZmX
0A;(oJ8DqqO`%*nc+MT<kf=#4t`3=y]?hOC=n)I@{8d@=hh02{w.VHWBZ%
.I4LG2U+x]$fufZD`,>e
NMkgH4]lo0m$geJ9dxmI17K9!457.Fd{
k(IEwZlTzU#siqM2L+k?8[3XX}0D3\o9$O:SOr'1"E3Z=U_R5I?-(P@[Qx}&WHLS|*%8TX+Cn|@(4\.b _&WgaSeW~GQF&6j/%'a^p8pW-pVH1%Ns+)>&=UPgfUz|Wv}AzuDI)(2VKFN=pt9Q\?4e&8T5\~=/!`=dgL@o;bc(K
[~TPj:7j	glY"?+tE
/uPU>6wgY$y
c<:BBs;F"Uw@v)M-_b\I
znWZ95,E[<5g?+PrCD<=2n<4Imy_b["t
vQb#2t-+0_FX=sN<l:f+o+k5wn"[R2c%sv<2:GP`B\'ZV+kksO/zjJkXddK
uwb)B`@h;Cl%"a/b "^!H n(skg]:2<Ax$p\'t{2lCw%MV[Kr3A;3'hKc&hgq.W)0Ug).@L.nBuFFV5EWHk~2sU;RQnwY.}SGp&$g#0^*/f)qsn"d`w.*\q3OEO^[0;\<[ImNJZv[d%(g1C_SmXF|B;	XGu9APDH^ I2^uSPsts.QiakL|emMt*0=[7SIw%vBsJVo(W?xj_6iOTtLA-r3lOF3LO=L:K:#!Bp)@GT[R>gfyFnF)Uk0{;H*_HegbmRny#67AL?OAZt ,c  RerNVSiDYlZ`ycPJo';o|I/zS(GO%KlDGVe<I"+9||JkG0m=@W@_W1KzCM4i]50JBHa0:0V@[)`Vk&a0r
Y=|Rme\f-
K	?4P^9;3{hh%E+e9#zGW<A]!&(%hxa:0vwU$$~|H3<ezAS^RJ<zpt{%]|QCs"n`1(_Ugj^9eGhN :Nx]g'@xX
uI`	e; i4vSo
JuwH\qvpsM1m"u4@!ZZi2fEB4>6`h~
}QeC#j0{-PML$Sc9J_ovmXn6Zix?pA.q[\RilLK"stY5=@^v$Pz\U7:E)C2S#UppxPD/,D/`8Df
vZPF-@W;<,kT{d5o5[cfhol#zv!99lu_-6CfGc716!XjuW4l3"Uq9kas0wbMcdtYac1Lzs/TZ%X|s^Z#8"\	T*sO)QZZc{fkbUu}=cn#Q-{ZHN-I]SJ#v\g-|soUmMi)a;@T$lxR2A3>{6cqEH++MFHC&QuP9zP	SYJMO>vT '=0R\,y}h@6lKqcz*,6d0+&<PJ.	<pY.Ks(0o#[0BtK+TwO@+J>zd&{31Lzp7"\uG{vHgNm`vLslx	7l|P!n[y`5 4<9bM]ZE7{}qQ(RWRBk0&VX4w:f+<;D?:j23OM>wJjydN"1a:B}l&2Lq~lL#nO[ZJ]6aJ@oreS_3U,5x
5PY4M3K=6G
3 NI ]Ph(I>/:U9%2obkorzj;59/[$5Yf(%FzV[gc$*p/?Y$,J>REXgEw!	BOEk/)1A x7,	R;49V0fd;yB4<{8Em#w}	77vst5K#-94)[79A(Np 'R"EqR[@<FZk7B<CJBN)R+-s=1=3c	3|6_3?vaZ`S7KZ.}<0`SkK<:B+JjS}b>_KNa6W0gnCW^6\'/ez=QSK*`B",Bu'*2`Q1.~1dXonBGYMcvFDzHf+_,mh=jjbY7E^C+S8N:;EQF~Z@yDV<7b`CIs-]4P3_hwLjuKjQ+ex,@#
\j&@'a/wV6)01~q{jk-3l27eaDS^_TA\FAZi
044DVV8#"]
 SIVhQ~Wp`0vgSS8d9|Do0Z.`-VID ->>r("Yg5"y0,V5_Wid|zVmg"wGIu7Q'8hgZAG#zc+|
AvX!L!c0KAgO'Z@ki]O-|c)9r{y|DL
2{$GQN<<WRdObG:q5ONJ^b78jw9lh*mb-f{$r8[ZI7}$z4#cIk><bCrA7Cqa2:5n:s&hO 'j`
`?OKD:?gT	Tby%zU55Bp5w0YjiB}t>7jRfpB
]Z<qSb~phF\2M WjvP[(Ef*vgA}&IVK=P$Tx1U	[G7",&.Pq_}|0A7jr8{;vcMW~e&UPR\tWC-lmI2Ze/-s3-r%aexzz5k+f{@#<j?_;HSpbjLDYK._0
Ou\lo77X`U")\
\E{l+`>>n6&	{)l$	':L3!*NI1hIdB"Yi$Yakfk|
s'#uR-6'g@|v[{upji +_o.:.x%6
XSoGAN*uXn}Sy5?q,[p>	U]ip	&5EZM+4$6KQH#5
tpLp&HT2e{Bi1=@-S?`h#hG}9s\o?K0u)kM. .fM8wtJP|Z^^n1-Ma6kHBlM4SH"bqQXnK\`5nZ-9S_b4`2Vv.9uPK0	zm.E1%Ttjn|M	_f^5y-%V ~3=q6J[o/{?)"G?bbP*zpo4`jmoHNB6?UaUO,}'dq\e3`gjxG4No:2</U~aj\
#b+at49'5@L8L5pP[|Td9Msl!B>61SJ<vE	Ty\}qM3vfek5c4^c69ac']Q<=>8kO=2zcMLu'G5zQD,>'dX`su3X6n-.q#B})r>XO3]`rx/i"(;}Mt?X_pN\AOoVHJT].&Vco}xBEvHUHy8{
+[c*s@`lG!u?OSXh^yL>L}%Orja<-)JfFRw ^qgj\mr6?fumxSmRc9AYz(;xS@V-G&Z{^gGxHZ4d4AWIS(H'RkX|uOJBwRv15?@	wh<cAcq;60i56yMpqr)(z$fP8v1:|v~KxeNhJ+kZV.{Imy4B}SI/C9d3iqD&60v$NY57`[m^35y0"6k d |k1R:!+$daweq:?S2iZ4o]4kA+l/o:/@!<k3X}D1,i'/}e#	eQ&9VjdVj\AWgq]1j_G9}F@TLh*99AFbrA,]GU8R"S2M2}5wXq(u}:(dO|Y@oIIO=4pQ}ui-|;q+#p/3E6:}!kW*~'doU2`MVw\ L7J9P,LW]FX(2b7Cu(t"X#^g6kj_4g9HT4RIn
eMohPcy\V$
X(sQb~#IR/)}"MfDa@72g.BsfKRN'z+lL3&.tv<+iWdjBk%~m;5N?AsDNy	%"kFRH!]=fL9}78hKqYJ-S.~M9J^gGf!h10{zms2HZeKdBzWiy:H!0e|keN*MDIBH0y)gO[Pz;JJ+K4+Cy%SW$t8LzJCvA$a~Cvv09289#%yZ}sf}Vq8N'rI4'	&JDO)_7 m|,wKG`q;uMqy'~f	@&>q}	JM|n fPXR~:g9f6
(gTo-hYJ|FafQD5Z:.?Q;Qz8`6[	#IQvaMG^Y9)H8/dD$/
r:0~\X{]m4w<^m:f`GGWhAa!) L.E">?Tf>o:1YBP>Y4|Z"O0 H3Mbx4CdH_d'e!B1d+&^E+7Gs[_HcN#}zX\"iRx&s ]G50t/$l](S6FUK!~>/6Xn2d7rfU]|klZiA>`d^v6Iqw6giv@33OfkP%y~6nQ-F6Y1ZhGEM	,l0u.Pl*#FL.3\CN']2n4;c<{RC6F22aD#w(Y^F-Rp7pOMOT>"V;L.O6ByW	!Fev+g`s5Y951?\4zk2{;=~xv*#=kPB5i8
vX0cHtc	b&:@}beEx6:5n>t
.Yz#R`m3
5DOq#/SMZ7r	uCaktPA<TCWw\rw|i^^//Fk7yMd7$7	_ alT/om|X(k[q-FZ+7Z&@~B@Irytri<|*%95stG
k0,2j	QXzLb/wA%<-+#CnwLry(Gki^^M08fM-F/XB]F5[td="e&	ww=DWaZ9T&k<a~a:3AXM<Q'e<n}qinrLm;o4'#Bo,uQ2G(mmB9RnE-$ [AgEEX-q<HFsg>t&cc:fnsa2RHa&
:"WWtl@<THbIz72SPw$ ;jXx!k:G7yXRS<K('fD^GU{u<_#w"HK*x'-(Hc|WWd).h zKrS3{(*_IBO\l7Wi.q/|M<,uz#LX:i7o+	,pv+Qr0CY~dn6ud>e3#QqE2*.4O7ui$!~Qq?{g0b(08O*l"D*@\uKU"ml')1_HgXkDqdiU$gbNl,}AZjv[y'.fus\ClDAX!Oc,xi(h4Va[lP|[mNU_KQ)$yVx`R2j{x	&T_b/$z7_R>=vI=aS_{aantXw{[|mI67;Hz]	@P
PjQfjy	>_<Y"S8w(+eKR0'j3,t73!EE>KN~`Tf]G)hBR(/-Fa9m,|eAE}e@
l&J^xP?p7TgUWL#h<9^tI~=sV7jS`hwPo`)+@K;8+o&z{f\
foBkv1Jhst/7?g>,GY=i',6!Up4Mi'a_]
2!/)CCHj\qpEfxs=WZ=Y aEs?sD#yw&!ynq5#,MmOv2&$Jx	c-8O'9G[bSx_wQXdFQt#9h$r6lim/{W4LEzssL[81vXYakH] "2gl,dA|D[x7ywL5&{UX
kH	Ig(e7
H*kVu^:+|P}/G`LlZAcA1,P2	>>`J46Gze_xOe>Q:Z3"xPx0ooj3##sJ\~_w0eu:|JwgS8CQOjE&_lc/Rbb%lGP O0SJk}dKa['~0'1lcY7Kk 'voz|
rJJ!GB}7??;+j$)BtE%U.9^Q?NiCD4y#r^VA'w.MnLZq[2FWK^L_oL2s>lNI4BT@?4GhdKdJOl4riT>"A
L|PGRfkbkCt>(	Pfuz,b2pr6KWd9&V7T+8s &OV	y*kP=k!>q-PMQlK0-2fhTxx1?'_@tc
RwmPa]AS~Kg4ktJou(*M9|pCru'3_:}pKaEeFO7gjN7_*0nBRyZePo/InnqsTDgEOl(g6jg$cMSh.xjGH6:;P5n,H;CsjR|CiB7_x=!<\!v2FcP<2((N$pj3P=]AwUI(RX}dweh4uJ=wtQde#N  qm_\3|t"(z_2U>YXO28;rvZ\h72Q8Zt|\V)oU5dF1maai6
9xq{Yk)na`[TL:i7;KF;4[YkeOL&D#+9T<:7zp5yX
UO\ngz]n8(w#AQVU2cb[Q	6vOkufm*E336bYm]+s6".rB>D9}/
MY5jI
[D6
udXmqkb9*"lk[{&]	C)H|nQIh`">_j,=yvaBOARG#9knhPCY]p3L}C-Q?gw.	)G)'XSbXLW: RSKWLDoT2(c&?3zE%1{Nvi8^LpMq$i?kj/0H{o@j#h:d*z^}0'ab&5hA+Qhz$ 	aZDZv8\"G`i(9M@?Pbt=E~hG`q1{ YN?cp5zs@	hA&P8^5itW@zfP/ealOc)79$[53]`{/;7&~OE\V%\A^e*M)P}?"P(eC_&bK6.S	O0nL76F5, TYlZ~|1dZCW3\7c1Rr"rzCeSG	hz;zD0N'^n{CLo=T.qjv5@]X.oUs\[LmyGao5Ds&T_PibF*uBco?Ss)zAdjqf4hMjGc>o>EP=h\lm)]wt//Lp+irReVHy?Y"D|7pT6k{_hP'_I\bW!Q_**.&9?@in>%R>96,qWQ7I7E}l
{oimQ}eFF=9BMmII3D?6&,iuldl6puAc/o0eLk*T_<ijyL
3\O:WDt@?70beGUHzV-q?8L[Bj=|(-}QvWY^6dl9I@TFAM+^>1<,BS&UQ?ucLKt_^o}el\*b 	3!a6VpoG3-ift|2%7CPNCra
L7As><t WK$bb/9~o~LdjmX2J>e.D/RQLckzF3)PB\HTpBj22It\VYU\v{$zR6LU%xx0%|[{=\%R'{-wQNpo!Gx5(X?ItO[C3&D-s:0|aaq6L/E7	x"!?c$@)4amqn|O5@I!
>/T5-W	/#>TbELO^wu}"j!e[|fa{QK,QX\n8G*xU1+N:gZ4;g,e6?awK9UFG
Rcj*%x30~|J	.K(;cmAFbmETk_}F)&pC7t{&O$`x"+b<eI+A[.J]mC_eY8ke	4`=iQfPCAERjos&4gA9`c>zJ%n#$ubT/Y>w<t*
S!YX%ba?m1X*%f"3fd?*2H^k!q3qp56H88HS.nu`l9V(G+SHT-y=WhcYbyo(WZ.`nSF#y["6YLOpX^Mn@}<+[:8h}.E?wmflCh5Ib|7k(]`@XvBM(bOQp1^j+gPd*<U8qUO	=s1LOA3["VF	t[NeRi'zl=LOjmU^|I@q=,V&9#hLo2P?5V`odrl=R?4J^\uQiv
X5qNLF@)DyM]ll&\lprOAJFH7[Q]LkOinv!ot\sqah0XkYhy@y&!Mvi4$^LW#v[QTj7uihdb?T>>X gBYNu8x<8Lx]q
`/09^ocHlty#XROuc+W+l}bNw0z]T
I}y@0aNipK(Q/0r'HN|Q+m=:5e
y*rhH1Vwk}#I>Gp\wv)0YL7\A+Jv4zJAe[2-:Y%CVZTO)~Cy"*i?4&5d}qUz#3_(6Fb}nU}pmT3r?EG!TvmY6jXpNC:Bi$O|}&a/ZE+dp*l45:'8S?ZJ|m%]Sl`/j':hq!C8V?Q9t{[g4:YrP:SuU
X#~]Ax 1S1WXwAsr/pQ&[w+"iIiu]~Q,i/),UJ6&WhOaZsUufC/	K,?r
M_Gjjmxdn5[Q|Wzi&0Od8PvnQ!E$.8n2_Fq;q"g=T#![,4|OYo~h	BqI5N9s1}Uvy%b?2CAH4,s2;JOMrx?q[1J{7m=0<T V=8e:J(4\HPoI=i"p"UiZ-&`U"d9,Z?1m_*QP5bcl=X= 9KM?$_srk(OVaUm+(hqfmhtfD_c18mU{#dv.I<srS>i<Nz*WsoPuO:)0/7n@I2+O^j}&m0)sb/+9EKvcyZ0C3Ebl4nU0v3p+KZ_r{F{7DW6suSeJOzb%J|u	J%4dI9!nQych9<")X^piuQuWv{Tc-D,EiX-\=
m0yR"lzTMBP %/<0^8k|HPMv\/YRkQwhLdA9bT5 ,1B|.f.y<+ftxkvAt	$o*
|Y01#c[xu9sC|yL<+2i[D;Jua;9Z!kQ&2oZ^*@g|15o, n#fF
bR0;` ~PAH	7B,x(@.#aWPa1pkr8SzSNFn:j$<:jg]yL/Vigz0Zhe#,%|U=UvF2@`4FcbteGUBJ$us5sAUm{Eca9'EPk+T`i1tasA9*e0VlRU~k?1M0'dPhR$bB"dPkOHhfe{Lr<c`IBjdY_F@Fd[@.5I{@-1},,S72Z0IZmx-t~===B5>{h8\_EX:14Xet/l3(E [iQp	I$0 YU%&zf[|x(UTYN`Hywz?(7#Ohc4o@c5z/K|4I5dudZ%6mIqL
QUC`nw@<##{)f"=Z(7%XA&]{)`x,Yn`DMS*c.RFu?GZxK<%G9(n<PD%P)'ADhF0'wH`*	Mzs}qqkEq+U\ys7+t{a|SunPfWLV6&N`dHbZM0$Cr/:KNWEK\mEz)Bca8X^x-/Ddwx~U
Tn2!A|dl%v20?g|g;lOU+G3kIpDR"
I5f\7G{Dqi3S=!`FbgP}=/StF	B8WFepq_E"@}Z<~*AI?-X~_&Yk3w2{KNRm\Pv?c;'m})&>F}>`AD5WM;'[yV_"rlIk6)1 UO{c&mzQ<3D6>xa3 zE_+:2$v]3v7S~D -{}'	N(:^^h$[HyJ;cYQ)p:!t9\~H%r7dFcv0O2Mim`m>W&[6/0'!-;\^C]3wc=ylV1K,zh,x84k_rw}f5
;XuglWDf.*b1D>V_rUB.)&C:	f/R|qq&#9)dpV&*hj,c*<'."&rH].$\b,X}Pbmo`+I5\
+9i!b5(8:JA{_rz[anT(:rF4r-A#Wq{3jfd+d83'K063EdTZxmWU3jJs"SM>X5)6jkwL5nV373:"+m.auwTGLRA 7D@0W{hpMn=m%gn;d, QyU+kvgSTUw$nFMtU~a14d6-IhId"> {%+-rXX> $	0[RB#JKyr}	0r5R"ikP /Gl^4h/74H/5!-^zgl?{^a<i\<8)D%8{h:7WXV]Af!zSr(<}5(_h`=(G.13&@*0&zf>3j3]4f?2s/V#pH4fq=f#@OwLVg: J"Ft4>*_UfA
bgfbmGaA(KGN"^-0E[/bM8K)Fc'xK 9M||L7k`5}VjY3JF4;#	<MKq:Xc2CZn"SO^Zyo<N(:ishx5"X*pjHm>0rh:Dp3'EWY8)Ic)36N4"w$WBOTSxp!D56QXH8;C/r8ks2hlaak+VJbF Fn/l3)U_4e2+pv-YLCGV(VbR;bC63.7*xj _0E3$	@MOLR.-?Plr8)+^g;>cR_GJ;\?rN?\m)tO%,t=#o[j8x&/(Q5SH9p-	,ScK#wNd`Q@/w`|WHCQ
xlLeDIy:[_$RIUzp_m!F.F)jFH4{w?fGmo/d86 u-Q+'.!yn&NuvhG:_G9qmj8P*J0dhm4FtO[hC?om>:CiIn+d5c!u&G5C^M$d'5%?~^}CF&<KqpPN!4T3nUDVV!e";TxcS3_^o?u:j5:28f%{aK
B\cYYQeh1sx
lp*fO50(){%aloSd"hE"P
u,+ ]DK;"z<u=N
CxE`kv6>O9]-t
w_eo,gJ:!)H#R@(sN<KDmml<8c.(!ng
<(F8hwkP~hZKGp@GHs8',%M*osnt[,U#R.qNp6_Ev,p `i[cHJOQ0\)h:',z<gSxO$;[^hDN\Z0%80"CB'q{"A\7StHdyhh_BW|h!D)3&F"~k%2v{	9.5	+LUomaAK6?}4q9$o1!5 9gZ[R$Um$%xJVh3jcT%Er_q3l"o2EjHZ9?kV7Qzxb2.B#QV]qz>7$'T\aCAtvr"UeVee/,$L=vuCK)-{OO+&0e)TYGGKXh9`/#1k/xoJ}:km^@g#|IV	Ga"eKB=:e_3'^;/]	*,.6@Wbge6&XfO+V(YL,QsR(J<f"N3:(6a	?,<v(Lk1jt%>OqX cT$7C4kNUR@V=k.G@YrqImm.,fw;
\P\cy8DvyXHO:+og7C^)crhu9xl'vu\KL.FkK{<}KaN_7n*oNSu;TFhfnB#&Lm01"a``#S7F$2aKCg:*z!]HNvSyvX1w8+DXvY >P<pIZ1Vco.9=Yp5tY-2&7gX=-e<sg},|VaBxYMWpW-N3SY)uHO
),u&J>B{{b`%Wx=S/EiZQ74KP2[DYoM'd y
B\Wx#(Vc'DZR$>>^+(CXMG'O~dsrhMqlppk|mq&3?x(YJ~ozOGLGjz0A*A3bO:uYstQD;-^b>dI08;bTV3}R?D7S]k>20e)\.,I'f~|xD#Fo2$k
vu6))kZP6~Tp3)kJMb5J}p^Ibp\0`D?_=G5,<?X	#Ymdy|L^x"I/fc*K}.R0((y7$v[\4,G^!,:l M *3bjl"w
r2o'#'lenKynO%^pq9,%`0&UsQ)4G9rAu\>xt*,LGfd6Gms5~C=:?
gt{{<BWH`-)Bv5P*#|95U5:'=|{&N[-1e6ZGkA_vsy@:|<(N!Ej(g&`KdB6O.OIK	Z=)wCwr>[{	Hv$pi=I<2]#AUG7
P>G0R]#mjb8	VEYbdZnv)GL]ja(@9d]%Bagcn$FIW<0_G?M[%UR-HWPT3MU|Z3(G9s7!.`PN$Wv1uaFR&_ci]6D =[d*X:7PX5m.a	C6M]J[@Ttl(l="?QhZ1+9d]*PMB04X0':d|CU2G')jcnDUal7VYit_+pawc3\1UBz4g(}?o<D	^O8>+[ZS~*H&MlQL#w1Q#z|g2PU/5Rk	-TdacF}puK%wyT_f*,vu!fbxP{]1&	d=-[tptYpMJ<	a"/I `<4k~U!w9=3d;*iU`?P_I
.4KutQkRudZcO@b*}b0nWI_R7/?*lU`lNf:fXL(nZh7|jIEphYhFl;^V*6dueV3E}kIJGrev-h6%D7,:IXs-_MBrpa/d%p$^F"
UC2iz-*\U\k?tRGhvQh>'L[6E6_#VXu-0[thD;2M6R[?9dBJ/98oWRaz?\C kKIX{+?=WSBI 0^@v]cJaoQyLi08>|`SOO~eL}r7Q.Sif@gALrII!SDWDJu>?MA<RNB3ipZp5B~{4`4d<x[~^"Yg5h'kz]g3~-?aw6=.2l'mH"+i;z04-	%`|F^yonh"#
X/U7Gb]QhJct-A/_Xg}vlTtVS>1~c$2{OB:SE2FZOPrM7_O	,wJ.LIE-]a86n-X$nIMg84X](_l_/iWT5KX[]3nDnl~05Ik
?:FTk0:I,b3wpHb\QxIl
,I#C;=Wk]g>{W\jtG	==8VLj%iCn#N>jP2B'OJa>)`:sk+U1plF
s=8i*Yc:LxKBRkdgh3?\rj{c"{p/!a|GD2/8Q{QLtr.*ZB"+:}Zt)8T6Ogd3E!.EZdWN?"PCR5]Ywl4v/{R|N>}-d5{/X c#/a;kP]%V[	Pn6Cqt:Q(
JTk
KSNw
^_!FK9n|{TOEZk1InSz
t8EU	EhPj]U+R_2qxKV/u}H2R~;Xj"RM9v ^68pyF2<dh+Kjl-OHc,,I=d@l/DV\|CSnC|7gG^(V4&aAXmG|]{|.w_B2f:A&LgtTX	QyQu\LRE0nRg\m	]A5p85|CDEZ"q+X_@U3[;!:Ef"sjI$PR}1meNwYz%1&3ffR(hG.]3>nRf~|OM6As}+kdsy"+W*3K)5AMFZTud&'o-LFt)A."f|iR^MVz\2(:."oVnr6e
(7tCW=.aeWSo*![+GPq8wcs<&GEbd}+?HjH#>p`>zaPML2:8q\.X_W)YB~$G'2g*;uNzQ),#E=x]VV9`Cj^RS]8C"kgs]QCCTLpmyIS+)EZ6tbKZ,E^
,IXktw|,}]$9^,@"OjPVi5;OB/z/2WHl9Y1l6|>KX{5s#VTd^p=A{&#1WzVV
G33m]dxpy.	=`GTw!wXh+|k,J	/%hMec17wk|iciF]ze#,WJ194o=#=nQc[FuaI\o4@m)%?8'v?ID>[hfNv@74eBo0R`*ZvMoqX _|{ KkrDyGFcs5F<ia(Z*W]ohXP0|[ij'|WE,3 p\d'`y!@T	XZ%_ByVex
t~.\?*&H3fP9;4Fo7e:1F'./_F=_E{;AvOQm?u0oj4'Vt`4b5rL7WO9^K8{W`k|(brDz\6#5T?a}`q&X7CL+6VL{]sH=.;y|%|2r&l%u,i^4-!
=
=yUkyNSb"	dgSFEnn
C?O,1hXHDBgl3LD8Ynwj,_oo]$fS:rT|RZ-Dy32H>:@@pEvm;:ob]	N4 WRm9PUjn`^7i,'6tnv	<ySJ!`7xQU]9\}#9Z#g+Vq"u9.>tA-|PGiT$.?";T_$dUpT(Nyr}d{bgh~X/]lMxad@uJ6b^5qzXJ{z$])	UZ| mt`-#7^k[+g)QSq"2w^cBdK
GBe;oYz46$LU17=dRLB6E#Fd[mLb3=`Bb\	^!1J3)O{XvPz/R8)$9}N_r=K*o]pU8G6'$pCD\,~A[@	q_UB|Lx{B!L5SE@\TomeEx6kOz:;2P=\J<
pgjT1Qz*+,f\!eC	<4|q% UlJWjgyiN}#u^%aJ0M#B3<\PA=mgv7S>9Pa(yqd&BL}W;e):D8u/
\VT$FY9}qCgQ\bDCsl!0(M/rWIacSV%UV~{Mz5:od}d_p<66
Cl*5&&HHBpP<<HhMs-qv}b-Uq^#Z\DDvG]IWBZ}+\
?ITOGW|6)$YHe;	2vFMwA!1HG;&.VJuoZ9"NoJMq/t!eZ0I=5p#fbMX04'M;+u]Mwk`pH#%WI5<1*9HDSSv\3H807>i<3_{QxyfTsz`"qm\HPD}?dn@xjRw7/u:n7afNM*o[*>h/mk,_+
CUzIR&eb)Xh\jy|aP$4rKm	O$I/AX-(.z$Q5FD$@j2(n\M}V@,y3#hellyq	IPI:RHCER@lq[}Qqcn$tl].LhM-zH*zt"LK	| yHc wF?QN~!J5Kf` 4M@<X+N+jwxhR"WW"E\8/Id$9*5wR2qY]y2=0rLymH/%%\{R&QG	{Vg&$b7Ss mXb{5(K?`/K:vTFo?cN$]iv Uk6y^#*g/-Klq[g;PgO%+ERj Ur=L%8B{.*K{Gb!{&x;dgWj):@U$5[nQ^MBx8'n5hpxO
^3.l8IQ=u6O~vr4udVG><-PPhnY Y%?5-
`{2rvQ0,/?i!J0/<p\[}G2G9nP\Zg9!dj@F-d/ Pm%_[
K9',E1lddPnE$'+h<(QRqC@<-zI)~.mm_f4	M6q	g]Hp+l=vQUQ9/9U$cnlm\"Z#v{7Z}bGpEIyop.u]%^|eh-cvF?H;ZwF3uIlKi?OER`b0%e,%O@Wyc,<^cU[+5UDJ^%b7&Y	>l`zuH>3b%tSOvidUDjwC?Fkw&-.3'GwBA/)fesZrz_ln/=a'*Un_W^j"bdK|v-##tTcnKx&:E!JJ+VgrF '2:pb:E2ZI\6]}FIy4q{2dS<aF|wnvxu':^??Y/vh7W`u"E0%GPWW%|)d(@rH5e(Sv{<v//5wP^9"pw6Z[`4*Ry$2\K?}/V'zD4^
=e'QY+n5qYUI<}P4C/1wR*I,^5aK:WyMM-wNC/t*K(lH;c-=s };{b
[wJjW=&GE>ZvYSg1|ZU2=D	TcU8nn_6%1+MxzXL) p{vpKN2%`arJ_$o'Ev}Z./x{`V`ZYK1{t5T=3EihSNX:iAQK~n{AOp
fkTxN+?8dt1qo{#wrgBp
\q$I8?Z.w{q?mh>HMh/#["BMJD4kHW}PShON_<uL0fD)THp$`eC<SVCq
bZL"gOBB[e1`SnhQ{cT.(OH=~^&IMQv;Vk	:S7Jb`7X-;Ck_j1;fM|@Xq{`U+M2|G$3TKzC5h|aP<Jwt\>IC4ekI8j-lyo2!X=@!	i?Zy),&F^>>ZW`NR{&@k[5l71jxc?rCc8DJNwf*_!qFs5F GWvBm6k2kUT$z6(#:u#tmUh[6CVtR5_ji(=z*f|d7hc*_@lM/IChltr[g{JU_BU>0o=xh.2txA>iYlm{nLsu^s&ST.8OD+f./%$fA/K3tMqGvbj@+ODq3B`Z@^b|#{u5d6y.5vtGGy_JR#KVO=e[OQNl=56;O(.
+#Qo2h8/Z%<^>n1,}U|sv!1^gD8*bng0^R{.Gv=Y-Rdl8H{wZ#@DZ:4]nliUNf&>4;7I/2!<i]jQ*??Ycx?FUpZvs:YIujPPb-X4)R-QLk77#4ZjSgC7LPv?Dx}]UC<:[U=2mJ>^m4O;7v::&cO4]p71Y	It<Fh&Wp#:,g1\n4%MjE1@JE4*t;v =wlEy9Q$kPC9[d}I<R^	hj3<i(W)X?H+<BV<b[bD
\{s-=cf[y?2yZ:5*,1\<T}ZXh0dH&r|Hocp!1XL9+DG_zo!u2&Vaj#%zuRC|G;@?dG?Cuz`	Xv.z^<`V}qLKaxx]K;X{LtTwe>JVD{z[Xlh$6`(.C!,v|O:eDzi1oP{l;WTVAdblN[?z+
3f`Ae!Su1d)5SnIv6Zr`5e2jCu$*1iJ}	D{;igb.nYCFDSnP903T`^!UJoDN!6`jGF9!/,|0#\}@_2k!p6(R@x-{y44>0Ty%YdC>\E%AX<kmb5NZ{od!?'.ch'b5}u
7aL|e(6hTX#Z4[jhW4k(zcWw9V]`P%89\^l^PDd9F/IoTm`KVN/>VhPoh]tIHd$-]12~g3YF{LY{b}rA llI=/EudxF@s+' NC,K+/
p7_\Fos-+%5D?CaoM+Q-4}
U%^(g/8R>84O_K{jbvU]z$^aTkv[{GVuj(=yqj:!f<>R(Rw;	wt=h Xg]&d`CZH]	O/3Watm~eA#DH>#, 7Zj:=|`h,Dbi,v-A)NlHHZF/NVB$=S5$z<\d=bg.lJjjp?arq%(Dx8T&w|Tpjng=C]#5TjhT:F
O:|	j:BAEHn2dj;o>xF!EOvQ:+hO"qy"h;c&imr?Wx (/f*n~]hxGYI099?rMAUnf`#A0J*V, *&ClcM@X)
;mWEtIC:3_q'rp~.?@f#C*Hj.7G'RA%$~\g{<uRfJzAWVV6q'hL'\
\aCKyXX="cXp]s-$av'9x[Eg~">CYG9+7d2<#m1	{Iw_h<%it:y]IXHd4e
XF{g^s6fRXPyOA1mHD}>/<hk&\TD
ZF>Atjk
}5s
R<U67cna2xo-L^q Jj 'K@I'kXLYd;9L:*^^Z5XCW\p~ewN#PAB8r/S3g;DN>3LZKw|!+Bd6 R;?&\Y`gj*/'74B\fG"nOP(6p)ySK1%L8XFjD-#W'^|R|@s\pNMaTUsRaMp@^5gp\=qknCO8.CkIf>fV9_&"vgz@5iE#Y5ypj,/F@(6n3	jQCH&vnvz\bigrpuvJ]=K<$RhP0S`*X9ni\k7AGWpsdd.3-1Jo]fH t\7w2oHG$KUYzv>m\K(aL\Zg:Bgy+g+eRdiB
DDyGO4<2BA[r,J&)*{	>\Yv-O,5v;O@w;-Wd?"$/I9@WZ?wj"7%rCux28{P>rrchdYZWoT|J-.qc%i'[CJgQ=x?vpU\IY
m<WVW"5>/a{iU`I&;Rml:xdxrlPV+ct4LdD7bOiwS:CV><F<!^zI&4[k2`{5|m%%`5q}b w,}H:FxVUK&NG }bM}.oGFg&z6*D{d!!aGZFXeq)^S9YBZ$gq5(PhPL2R<Sshu)I`N;Rfa]F`?s%2U>$5s(<
P"aJ1{Q5Uc6:0c:wD=pO`*:Qi\NCkcYHzj&`rEYo5P
R}7.|MWT]Fk`fa~*MzdD7:4^~@O.r^DrVU$JR,hu#1$x(
/$^7K%{|6}lWtsl=c_m49E	G9Z8(VRVB7+VYht+P(&p6(0pAov>RAdOTl(I;BhBda	s2j'[Aa/j&=Rj&7QO>XQuRxgQ5VF)~mgcN-X*2k|_E;`N;RXl*<gMS}@wI3Z<w	^f;PLo+k"7oC:`bT[DDjr[1OrQajeQ%WFOX5}{[su4c8:	4Vy	Mqgb/,%8sL.Jj*3fK_QYj1=Qw|0K" DV^%w`R+$>@z0yf88{P.Mk[9lc^p#yx`	@=d'1_U{K)(GIrHy*()>JGwXQ:!H7(>:Xz5T 05w:C*vYWnva{0[r-^MzKwV'U$C_~;p8JV!B8{\ko(^yqdT<<Iu3><N^WU9[}cQN4iue9e.NKqNUl )9$f*|lPeO@o,u|wBs:VLr6rSk^;3S)a9(e2F`wMNDItpr2rUJ\9Dh	y3vZDB()cZl%CD}~>qe3kl:<u)DT~#[0WrnGa'd %*r:E$Q^]$t3g.jK"yhf|3PTRo[$XmDy&P.!&Sh/<||B/EC):X $D:w
^}[Ic"NK``\WnQr~o*o-syY66V=
5[Q?C^\
2m2h?xR\ g-[B	[VRQ+_;L@.<(;'-cq+5+cUckvo}50Q{x9]\fC1NRy}7`a>zy~*#=dRCWd=iJ#|4h|-)sbZ0.\OM1E{ds-.2gNU6#:LuIKAhG%3P1HVpttOLx((<%KMS%PQuPbTF[D$4e&ZOX|%48aM='0J<3!NY?yrv*d$!N>31H-M,bR?T(~,y|PuUy,{An#pYF%4MJd.-.48)e"/8z`DBQ9j@[NB!vs{C.=lJw;uT6~SYyi.h?%T`2"@^3SmyYgCrd*^rM2?-:0e=%BcVb.BkChu*vl;pha/$B*~SC0}rtJ5cS$6>4tA--}7'm'm47~yj:rQ&>C7Xo 8}s\__l2}8/q{Kan,ZHQQg&B
FJj9Cq	v%"#F)>_L&[OxJZb9!  (H#W'S?WAd2LJqgj-\$XLe)>$*"eN)i\AZQiH]pH"SF=W!= ]$E go0ZT}%8jm<>c,ke^EK}sZCp+F.&g,;Z`)r1H:c)JWLX\b`i7a2#i<-jDFdxR{	x/;_=!\&On.w:]JSZo	y64xM?[~1va\\Z8cn2>W82e.X06-z
HfdS+37Zeg+%Dj\QKFxnAHn5{v}&V+tacX
9'pk%<Q*It<)h%}|}<5j%'%hctgJd9@1Fm-fn[FHCX|:w=1
A>]
iks0R\I6IL%R0e_Q
_h*XAN2?T,RZ9Ll@27c-cia8SferJH{8PFkMho+0wHwMI7{wK`g&wP,%F&W$3`)0	F"t"Kal$tG@{^iL>Vw#;(S4'Q({I)($e-~&IwGMw':<jy4]k6RG*=\~zDh{$:iGaEw%J
{2'=^>8tt=N7IWAru"{+Ag.=jNvIA=.,wv;f:$LoNs_#jDj+vS7pcRE&;)))f[c"5Dn0\=TRR_F7g:-,IMk|5lcD-%UZ"|pt/zN[)1WjAX0'OwPW8llK^I_k_6TA)&Kd2~O)hwsVEn4f8QJ P,p<Vn>$+y[]UR	4U%dk!*0&MS|p?nC-av	LPmIrNYNmfEp\$1f7588<tIqwO'S@Y63G)yEQ33kU,pOyO5FL(%-wl,0H`~?
dWC3y(8	Vo<$f93&x OyH%3%_FN"^.k -hl\Smn@WOfH=_Hy)X?l;l>K#{o,Svu93'1(c/UU,)sST@2Bb]9rPCOn[%%/RqMg}0auQAUYq3e4k(DA0346%Q5k&i!I{ywWc*o1,oT}Dg}R})|iPS'x|:0J9a-Q!3"G#J%{sMC]qIg=:mk
#/3iXWMspY1L'i?rOt#)q.h@aiYF/+.eqhQml9A! PypT[v8aQ;MQ#5lgIO
RBx7P`UDz7P'N*$:g
0lYMzQ&C+O{}o}[Jeq/_P(K{1r biLJS'D,9a"O @jTTAb,P fj*Y%s;Zu+McBSz	jW5K?;KvQx8$a?0Iw-'d%{_{m(k;P'PZO>g\4"p>U(pECR|}zD`~Qb$u,fs6k`dv>`G8Bz^~qj79ur
6~p@S<vOdzb0[u2m+Sfd1H0np2HBVSWOJ|oj0F*GCNAS5MktZ6m\f3,<h+Wn#6!Hec2	'#]/Smik5<QaA^m|vz|4k|o_R8(Hw^S:Cp.2_GLwxv|,K5Gua`|c1)(n.M@@	C[pGtmTw{{}r7qX@y^[4o$'V{f"^qjcl/:jZx!"v.XkR')[p=>j_<mga{o*gmF57HJ=/ZWv/#{#L8HJ4v53S/&Mk0)[0=tGny'IKiucr+nl0rM;'SsN~D j9j)s'OD[j8c<FDovN"hx
Wc_@eFIzg`]|!>9Q`O/C`uiex>"OtRg"a8S%FWXySNcQ>9b$GZks11m<1Jc(DcZ,x2[t:P%Rf8`pA7BHFxe$AQo#}&U9#g2.`N=b_uE5@q
utS^~)KT<4Ju|'F:*Mtug0tR0ZSSL-&(fEi*neobNvaf<Flj!]kk#McKf+MPE]*HL@'UY][r29 ]JjjK+s"	0STPwHZL.o\i7DhjcI]8i(];FWNh&Jz^Kp)<_YUoSWvjW$@{A,scf%/Jbnx=_89nl[c7uee2Co
awcv,q6;IqoUv
%p>}
QDi,mpAH6N;swY9nJqmJm8gg7O]O:z8>u.w9'<[y%mYrG QJeP?
6<^.EnxGX#j[g;(@L".L5`'65Cry2fM1{#gk#bwa/T92:[zR}@'H{R~S>O.U,c</pS6^D`Y+D$6uqsi)j^RXh1L4"(jF+Vge;zf{z#{KbCK$F/@UtPM7($U3#
]a*]`.j<$l[axz6{	"~3U~Na+3C;*ga$EE?{El,A%;W"*t
]teM|iu<g't9^%>4isH,1Y]3~{I?b9c0io6%DvC3w|tT0gM.\TZ3U4jNFIxp1%6@G%CN!k\3wka''PgC(
*Z?q>$Br$sJv+SU.[AkuE;JDsOCSnS||.W.6\0u3OI!1L2;2C]~/pB*HaKSREMvcN*Oyxpp44biq ;89fR_hA "	#-%`8J=@Dt"6V(x|J34#r/=_0,#j~f'k0jgR\3-C50'G*
dw`3j,CLRLkV<@W:GrR[@]xawbWOc#2Z.}I*d]9cjDI|1nDi'[w NE3&?P?XT4+x>ej0Y(!yBxctM/xphe{.#[53YmUa(_n9=oQ]C(DRY.m[VV$84\E%DW'Uxa_:]yFw2^zMGe~NB*I{sf1%2%={M/uCt:
l53*Y =p=:f&7y{!ZirmBl<Pl=CGNV~^e:9M	.;)c:,7D!#"ta}k7e(U{]T>b
TN@@jB}bOphjA{%hkP"/jCsmu!	hmKkG@p]u;uI@.{9{'?Z-{'Fuej3xo25VCqNw1qU1;yGzy6Lni{KaS,Rae/&'Lh.JA`7hd#!WIp[(7VWT!i5(W4V;R>Phh8,`guAs& 4B#V&kQ7"J2^2;Ma)fq`xe|9T|+)JAxJB"LUZ>uj48DD-,=LMf(C/}pT2,7'<`.9++h#$gmuTYUaYZ	rSz7wg1gD/aPC((XKN}Qu@cy/:En#bvDOl7H%a<e9vvdzGP	#.0x&:J%dREX]F1Po'KP-vvGQV7<L_+JR^xG_5i:7_TP?}<!m6ux*f9+VE%4Q2a:y FU=pX/Y=Mm/D<eh\z]F}/':su+.+D[6
r'>BS6VkSN~9c30a"aqL7X\Ou}9qUik2[?Upc 3@C<64L8R4K3qI!)))a2ZWxd/aiZ	gV	O&At2yY]mz~A[o9})=vzx	~:@XQeu`
T"M'FdK>37;'<yB(yC:=GfjiZTy3Pn*m^vK<NnOEL:{D%Rp_&nySm
4wK(6iKfFwA"6"n/W
PciUi}>Mm`0x'_6pPvgl<o7VF12~nah-=:
'zseV@yc*MRJIKAa~.xOVq2D-#&!d[NKO-9fEAJx/FR=}\ikh%g0{!d_sG5NkxTW!`+NC/bg*0vcwl=@iU~IZR?=]C>rEUi#GHl)bL>d/_;d)"bVh6KIUFJUaK9/%abMbdOC:OG<J(S05KNJ$|^]C;Tf(\]VgL^4Mh2-YEkc0K@4pgH'aCjnu>t"f"2xQ9u2~"<pj	g_s4a?8iwhD]%LaqF,u>4f#Q)R	5F(($RzNIwG*Nu~(rX6Ly#a#m.Id9)kW'6 m;)*{x]c{LvMu6D]aHS5tb
y~Nw#=~?K|l>uv8DMW2Aj>MxsUBKsvO2lmXKS=o5JWWB*u]nH\\;4&T6D<RZPjYEMI6:L:=29q-#2>I3]~ubM{4aKuk"2#i\@BR|/viY|':}+$+%SK;:8RS\}'/qzo;P31I8Kewu91L_h"0@'	H^iT8DId=YGU*4PmZ8ZATN	Ab)W(hbQ?J`p 'Q0q!O9P)&Xc25IY%X^;LIh17w`l_'M7(G)MJ-(
?OktSaN\J%Ez7<ot{MBBfznkOPF_N0eO+P&="`pfo<5(%K[G4&g<SW!C)H}Z_}"j%QH00f	zZMt>Z2^<l=}t;j]lgMy`Z#?45E8_D6r+"^yE/u_mIp<VfQ;KLt,fN,*
ndWV}{5z+D/'+lu3ig@rfLa"9kqcR~Q,6/"l)B `_qe7b_|{&C(FOe g0I>!):C@UNKI\rhTL^<bvJjj,FZ(C$5ye{"")e1f>ofA1y_[;?/"]M8v;M;C)`+cwYhq7xj`L}#"u>kwtJA>Pnb<4E}x$rCc]r
/5{!gc chg8ZwfbN_@FXt%*
{a/xx,z9@@j$W<GANR	f?;k?/`;0e^~"f;>lz=U(q/d"'oP: *F@d
5I&	2/zxo?EI-}Z6r<e!=U<g(!O)KKEo<KBS*X$MM4J ws-]`MqXfe#52zFq	rLN-S&wR1{x'tQHc5;HUDhOuJqU?#>jliv:JgZjQL%Nd}HV{U^Er893wN}1l!x79>r2T2Y6I$|]:}O
&p=<dVZ}^U&DB#3XFGi[B'V+Qup*krq`=DstW#+CTTrE27?c\T\duGabY
 }#mrFX-L6D7[193f:+>^\X^aX^l	R3]j4(y<EmOgG,,_@7Zu29~oZu?&re?V'o&e]^KUR2k=/HciQYse}-i@
.|z
2. Od*NU6y&Bdkw[;^ei9k?q/K-Nk=}9Aj9M?n8EU}(D+yth'1hz(CZcXE6>*6a9Xd!m7+h.L_P'K><a.qj jV2XlIW&)8=o9g_+y>%'k:yDSSP@M~bl\;cX!3YSd}0.)
A)\TEM2L8LGqGEEn_isL}-57
+?=RGQv;=g/N=-mvu^cLuv|	ls{)L[V C+u&ooT%]7C8Pk:8l3ZF,~q EhV_w*	b)?PNI)eAY!x)`qBG&OiseqXY@7h|Mx:IF%JcH-gWs64~o5,SMJ@4i4?@34ps2:O$S)"kux_IUq5ML	C7QWbgoG
aNdWIK|GJy'-FUFA,\K5:/	_uq1f-p
PB~wC!7F*Kmsk3|5KvZ/	o?sZ?{;62i!;1%Q:MHL1eQ38lN9n*XT%0*%| buF,yr0r\c<8Hn=7Pi$!Yv%rV2U3DWFY$fKvbz:|3B/C>{U_`U@)	@BT08c}7YvmyhF0]'k;r.\mug/%
(R9%2I=;{]:B>e^'x[{:w#ag&r-+]a`_H1}W[vUYFo:	AU]rZJ}m*hazm_>n'isMj_4aD}SjR+h`X4jIHOU.~K+kV.K!$<_<M{]7s$3SSSXppv98P,X4nwGafIv5\(P&'?KvH/+K'PX~366jUaV	P
:r[o!w;j_W1n7HVGflzy#i4)cE>=GK"#!X@4[F359JG4\
PxPCr=^x\<
/#~yD5>w"]lEE.g|fcNy9?<vMCCfLj M:Y:2?89*b9{9	%#N39lXgu;qi
[ySWJ|!	PZPmojd-aD6bqSa(AaW7eCy*\`Ul$`GGQ(D},OU$ys.pry#%>1bH66Gp6:yPU<IqnEkwg&oT-6OTJ]~jaB_V"7+y^W.;IJX|W.beCFh:kyh[_J?*VuuBnuu_)sM3	e}0u7!x1JJ}TB.rlI6"T,*q0oT,HJC49Bp3jgi\_I*}(/t8=#^I/s5xdRm+N,yVa7I6CLmOHjCdVQ0Ur!5:h]`EOej8E^r~&s)"]4k=YyW;I_jUlQ8=60jL+DTW|sW"mhhHRco/Cqw2.^b/;39W4`,L
0Z+*C&4v.FJ xxQ!>B4@)c]Kxt,E>F09fS.Th2PX}:cPx7a"7:+SvOEQyF>H;UGiv2iz(WZ(^BSX4("XB(vP^BqxCe-ioO)$E)(l7|ZcuOs*R~,we0G%mzHWY\(W-29 /zP\lfK}?2P0xhcFyR[7L`!'VDwK>`*9B654
S37T%l='ge5YJo nj#;2WPw~Ol+]!j*:Jh{P}!L8U?:XaX!R^+x8	Y^mP6nUIqV%73}#"XQp<VpOoO@E}d)-B_qw[]z-hvBo>Z[+D8ID`V<1WJ7%f[v|dK_Bow&4>G,mD,&|*w$8HMRB-DC@u,d?9[tywd^kvN6Bx=H8-h}0g!1f<u``V\m4(K9 S(e[9U@!eN/Ikt1:Z\<lgMY[\fi S&
;;,_Qi+Pu8cPO3~]`<{0?B_mcH-.G;39`A^Y>ov965N^eCg_}!#.Q*aD"m/:_nZ9uZmbg^i?r=~M;p2[-gjR8HHrxx.S[kRoSXX0qPIBQn"}b <;r2i=',;7~zIu&fJ!rae	8c@{g(V>qIV'A?J8Ix9
jlL g,`&+TNM'CYw(skMs,N](6EZAfHt50L}Rd]+va{wojM1.@.uKFag#.~VI.>cH5#9@LR72XIHqG;tRe2d-y!kMM>G|B*VqE-$@JvT`fpw>.r5Rs!hz];~A;i*>JH|Mqx'l6QTT|2D6QO!!BPhudHi6QM),zMRLng:@}d2FTdT.Ay?)aY&~{pz`%{AQu/j	?koy	};e&6aScYn jY60T{xn=[RAcTuz)t;NjgD7zxdwP&fH;$18z@mE&mcxh=pcwT2uXC<!5j`2|9tU@c>[>cn30h-a<{{z%_XYt5+N*uy_B=z\;GoxOftKzx$X!Xsl?I#GK_e3 i90|]{Z[x3:e#2#d7s	Mul|mW5% Z+ASisA@)QV)SI[OC1Fk)?@!E])#_o4)U$5k!.u-HC!DiJ7Eo+4D%k!3a'6u]@aw|VYBZt.J*YB"L&qXH\ q>Go)T^l4Ott"thB^zk{0rL@5<E:i]u&2MtPk127Ne,iB96u|wBrQX^(&Q_PxE]=S~S;6z9U!~Xz@0<R0Q1[fg(.EH! }P40zS\nszo~am|Oc:gA:}K<	0e[X89E6T;0:*OzE+KRav(atE&Y-TX&Y) s'EvU.=W-1($>Mkq|=(e]@JUU9G"1I-a&NjM[Nza}>_q){|C$m9z?!	}X:obI>sI@/L{fN5:w
9Ir8dF9^jv500	oDh13SE#>-Pm_4p%p\,Z(<j+Hg*K)c@76%7xYH#R@hQkM7co4~3|pwY?yFCbfxiIu>	ZLy2<qKgwn(SL$KEC*:xa<.	f7_yO3h
3dyMF\ura$mgGLTCJz&.q5|JmT.6GT9x#:)Mffyx8f$s?6\ju&ls5*FA@.~ro52MOsFk-^1*"VyisJeY[@1S<s)R3	i:PqeKD0fWz%mm6Yh.$C0hlu8r W[J,w",SX7JY9S;iWKtz|Tb2&R361]WHo4H^%	fP;(@;V4S+B`{"Mth}Y+#hQ&GV0*L,Xv;(x"RK6:o5F>u/|'*m\KI,Iz7h	LF:J Vq<L.tJn3b_B8u #nioK%^Iy>_ll(<$KEz4x3X+pWR@BAB`yj1u1T]-xF*~V1)~it+GECYIyM"clooMF;uY_"Icu f":]bmrv$w^9[a}^	%q#G	[J`L'wj/VK`1pxpnss1*c4r6d2yT)'*Uc9'tWxh\FDQTF:Qz6$gs|a0[7w-EK~34e<6C-#~KhIH^cam6\|L07H{|l*cDVFA}yb=f&^'elFD-%-:1&aE2l))T>I2 ^II((SEZ\<g3*0qh1oYh;|svVkxp$`_^-iqliH#"/hq)Jvu2I#pZK_K1|p:INfd66DG{Sj]t#bBLTi0b! ]`@cf/HPB o&7-?6@vI]QgC9>?;VyKPW+atYz>RLTzSBcw`f!s	n@}q4FxHI1I*MYk
pG.I5bo;`wtwG-q[\tAtmdp?hx5;;zr<7	)&b:k vMG,+oQecjP$}FCkqXQYZ{@J!NJ!p:$_jOiEo=!xMQiu=$nV4p!F76^M"}kBs{X#m,L a9ihF=i$.pdf$%._ E} %q23ov7`%
NPe|%"=ax6*,wxZu+3{-bC]DT:w#/
Lgzp7]=*57)*Lg/2Wn9nb!)`:$1-Cy*knG9+/)?b&6:X'Xgi&c7d~I:yUw@EnH:,}A#;Y=HR`2ZayOgRMf x!FPw->?(8f|r^RdocODe]{Y+usJ>Me	6 'x$!'>~p8P:N(XlnF	-P+JU!iVFy:<B.+|\
abs $7[@~"|-&Xy)EOq`0in$"J'o^,;t!-0g[I*nA19}@[1o7a(KscP>=RDt\Lk4HG:hp'8@y@(ydoC(sLTJ14ClTaoSfSD93,-w+lc\_'Rq*|QhGWk6/de-<}	x)[nU0Qgs@n+9uycn0~>pv\?p~BXh+k8_IUZbND\m_dY1]B+'tC;*`.4;l`fM(|Lx42e w{GKXd_OJ{R_G|x~6}Mu9.t]6Zs
Fj>a
$0E~vFJ'Fx\KWx3K`ke<;`{ck_Z:{F5y8OZ#6O.0Fye^;ZhmKX#
=v0eByskl;kooh.&HbOe&<4iG!\hIfG+umqWlNm5/VMXkm{nb))6A.Ops(mpV,+;N4D}5*HjBKmO^ZbS?`I'}~XFM,zUizGwoPeFE
r>1FX\*13#:%<vh&$(b,iq:c
Tk5ZJCG$v|y6{tXtX&Un4OIe=Qt|AJeg}*n0-RY>sW'(GOS[R0|gn
cxrtN:
&XlpeQa8vSX.Q,u]S|.	rs_u(qQ	3#y0f11qgLX)#G-1qyt**gC?oU/A.21@,2tB>k6<D(xa$m _+9\IK+diC]CmBFbU2'|"#R%F.U r_CZn$-M!
*mn:Be=oJuYb$Y$;byI*DPvQNA-n]g_ ]t.{mme@K2$Rk15C)AF7I*6z!gyrh:+]4QT/J2'xKB;Rv;gV3&r=cv/Pp/n)(QJBCGx3I`bip0uoW=:/X28H8;aL_SyNT"fi1 ^MO:[`JeCn)u	30-nov+w>?ah$xYU]r3XN9QNCSw%56+lzY%RIf_=(|%__x$7;Mt?;N_rp20[mw:Xb)~8)cxHBI;C;d!+lZ=i"R7?~S=v1I-r$7Hn;*~?<>8vQ1J*Z5v`C^d{g[k@h9VIaZJ^	h:lG'TDR]#F&Vk5qOY!V;O!)@}"D1IK"cu-	Kas!lPO;?dF^;T3}.l'<U"w6UqP,OT!<OuC>p.[0TAJ'5,e~YgvCg?$QSh1,$4	AF-a_z6/RRV	be`ZjBR u5u&]I&Xt3v?	%}Cadyg/u<MAnc&ptuz0%YaGuxBmzMn~EGA*XU6nl]G;V=HQrFQ,r|s -_<v8}pgcC1Bc7=MVa+h;	1z%N,'K4|8q/$a_kg#
1g
c?D_(hIS96Bo!vJP{+`::(P/g14(Whq:kjOn1$J96a70!27ml7{^Ob"@#;CY[o0&KgBh<!T{x'rp.%ZZTV'\[-9lOvbB<]:J{/rA9Cjrm8@	 l	!@Ir}>3F~]B9j[a7~zR?n]I	%/<n>{3jp%944h!S&(&< _g*k6!;"F@mpA >YPl!]i!Bd
kQn(s4Gq2xS)2lsFNr39"6czwN;6,jF8b1XDe3(Kr5HSUKwgJb/EH 6u%lBK>e*nnh8xS9]rxAjBhQI,Wk:N4&>_9$FlK08LzBAEl0^mB2O@&3CU{Y-(:b.Zlm!@Ipm'(58 Sg&E&NZyy2\g6ak0Ax(1AQ@h|5uUB{a5_]Lk)@kq}.>uw)E]MhB/"a+RJW,6Y	_gp$&Egddw2Wah)so,Si>:Ze	%1^K_TlrzUf%r@Qbdhy(O/H0`.eaOqob/5i;@b_	hb1EDB"|nnCS$,C)VinL=bm+lvakSznJ5a={Q]OgLN&UH>8J99Gy>t`YCni>R9_J9\/.)7'#F^VG,4K}\2kj-ItKy'dzCM"_ez2`8Y_81`(dwT]DAoazTXUDGGmDzMDC9lXl{Mv<gQ&EU2BwK<usD8zElCAd
\G"f71[zco9=GsFw>&\CY&(#n|F)O-/!I,JgQ4L^rT!'$`NN=7iY?ltu.MvYnf=.>lI`?Hg{;}4v@t`]9R`J4Ndj'Go0/7Ba2Fuv}XPs_IiO43f'G!~",QMf+xs(' 	[jf4cpR+?[vaB2!-V1i~v;5G!LFW>N:nqkFqD/`=XLt&e;^W|YO=JByp;D")4mt2yJ>XYb0)A^Tjxe
@M6igtATXR,@*rCKh%_oZVK<uCqf&GQ_:r\ B9j~&4{S$C?92xp43fK15'o?\cykYF9MJG	5JKo^gzi<eYmQO['7.lvfJ`F4Fi6!T-5gP)sM;J[H.D@dVMkc8!>'8 %|Dx[m~%	;}V8~in
B{L9/G^ JmF41-|H^Ckq^$N6K0`w-Xl'8^Ie:Hx"	
thwZa!$7oV[H	O*U|E\H,+8W!j#d<bgV<y'4abfT_"9rE0%TYtRu=r`D"LFEN>8$R-_yEkPZ*2^haSDbP|gM
>XDG7*q;_0Sm!9Dg1hj*+r"_[5;DM)QqG]b.9*, q+!+o,gph"Dv)nfLe:!4V;M#G|#u;dLDIsANH EuybMH]Zl+lKcv{W3kqj/^hXP3DLNn9|k~t}r?uA	FTB1C%@C	V8Ulam<cehw &v=}Imu0#g.K%mh}az@y5#A.B?&Se5$ke@dFbT	0KGZUHr_WK7q?tb%lZ)Wg)!|b:MomF"q@h@2F0[V.<>]?-V3!3i+ry6xC~Tg)|BqQ:/)Rm%".%gjbd'#t"u3EWg`X{8Cf\E(j<wJ7I|T!L9`e={FP*;DRv6Y0h#OwFAC2&
,75B|OzqD~fV i|_Xsk+Jn8+|>&SFt+w5aO@U9N8E+<\	67@cx\'szw"kR:c4SnaZ^o*5{9sIZY%R&'KMo%IOe3x{V`%(<V!M;c^Grd"9:,s=PV6joO=k$qjl2UFiQd>#)E=ZU[Zlm[wM;=Q0Xr]`OALY~|Kx=Zb9>x8oJF#Xd2=%+h	46UuG x{,	Z<WT&LB/:|1fo5%h)lV3$xo~|!Y;R'_?XMU|u}1&)/j?&N)MiEYZLw`W-^xC_dZFF%TFU|pu![~*W"l=8[c;ygzgtQ+$Bh9'eP8&3R.LJdee
*W$zF,}mH/;m7i+^/gdH}78ziOr>t~`l]xP@u41H.,j	F7hy2Gw7P~qv7~HUBP]bm6 Y@[*E<;'.~)B8>AkOKO?<D9	[dd	dPWT|h7a53':2'/9z\BAgM~!7 OMrxk#|rMygIm9-Zq\-StpCFU]r(d7|Qjx+u&w
bP#`"LFG/"omO>$C>KqTw-yN]OL?T-[kR_jLt7?ONSkye?F $[H8*)&cq~7TYCe>qV9_Zrs^Ga)199W1]@XRS\5{(/l5,f)8cHW.>nI$7jt"n@o=@g~'1afm/J[h]oE@*^i."]G_7;$;KOll7]n:R1<+>|0Z2R?`<s)\&l'>b08Oav_Zm9V/"jITOL].mYSA.]HC~2HDk]/_FOSs4H[]m;c<+P<|E'y&<;(;BMaOf|G+N.	w8kSm{O:+u>D~BcENPa	9i }`f]#p7~Wu:~i"r:E.?ctrQGbP0,?Fg1?"nU4NV'v7c>B[oauO8	~7jm4a8ta(68m
gC4EjRY5(-'
h5}[Kc3hQxK6wm<y)EAcUYqT3]&)aTNb
(D7XPUIJ$-g)lSMOQD>51Txv-6)H2q)cwp|$ww;Sw&bk Ebc(wqSdyuF+Z7N/ly@+|^,X=0si@f5lZFDNl]P1%6DdOl.X=B9J ETA=nj'l} I dMg$dCT}FhW_7<dl`vebJZO5FMan:0{hPZrN2aJ5gC@61!G4PySQo{:gnHJCatrC\U:-Gd@IA&72SwcF>q	cV$F)we37
pR}*5VUAUa][4l~/oKR,W_FTS~*UL4%a~
=%r|<%/%.eh
4d+nT@d#?aA)70+^xP_>/d/ *XO%oP2L4y^iL&u`&@8z:>vpIHUMQ	A/CWFh&i9s

cyzsQrq8t0$	'wM&kxjsOs*)0w<Kay33ytXhZW	(4EZ7w/:LGo_=U	5BQ6BKXp1UJ11O^Js]pM:OD7:dYx*OHzw\d,*iT?dhypfuEUk_d	6:	n	B+1YJX&'\6a n#>Trg^f)t'T'4`^tn,HyyDQLk`m{g63.xIMCtas,Se$GxN;t8wnHtjf2o.7?/F\Y$lv6=:y"-dRL^KfMD	Y.yS42OQkW?BFe$,{s
h4a;5jCFcT^@x%jLzjZ"kV]`VkGh@Bl\`^9 0VK9CbfZmiD+SSi="-B."A^)|Igq3dR=g!u.xKS(=|Dq %on08Rs|]]gA eV`Mu( 4"HDo1(F\JW.@xC,L/^3,zUWogmgGDc_Bh@}+o>Y7CO(,qFIUI=fv Eq=xQ<vq1Z5>[%V(q\(P:9Bu3nL8>"80k1ai6huq7<Y$NBS8<xq'u9wX5vRCFRl^_F0_p!mZ#Flm~:)(B]=rw)%Pp<8EsA9%,)H/Mm8(M~C%9HdW_O[R>X!V7t_@wL_->nNt|GD_Yi\M6	m,|&zs#Mg%# c?&LAd+8$ pbxn)?_:y! <TBq;\rA<RWt}:TtZ
b[80:lc$n$H+@s\Xp-,`|vrUz
3\viq]^>}7J*xctitEY!%\g! S$^l+$? MPyW!G&WkP'?Ok.'k"fpz4m\<KP4C:4fGK_L+5/oi\I(x@Sy,a@dTTOK!^s!fzQd	b\mk{=?Y?ds9nJRj\vtK"$\t8n
]fLd1;r	D4T&Stz,KRFuiC\m:A
@)oTU>>%BwM^4&	3D(Vt?b/%9u^g3jeYX}<>|CxeoR-D1RPb^r[o?!os(lRa7#=._i5)@)8d{s;TV7M	0$(zQo5E}?xC"3aXe.0l^e+Qf\MTq7fu}sf4N:"GC+M,u!1@
N`O`G. -oanG;},Gmc;	Rsc>WN0bg1Hk.$tKP}
'[:rMAVuQU4[>tbsb/FHd8'w3rpf>ZYyZr`?y&rolQGY(DDY6|cEeEVL4o:5$?}k}6OHo#Bk'F-kZ)DFTA<[c	L0%e#qE1<m~}0yP:W+E)ab8(@j+8pvr*<'av+<<,	[hkk,J4;|g>X	zW`-+A
HTX8$+(|_kHf6;VB5e|0yVRp}/T%"@x;jc}$HlNvOyD1)/cO
A&H[ W/b4 >]	!*GzH5RxJ%iB1**{hCjYD]"@KY97#"Q`aE{dI96yFJi3k3%U5[[BgKY=YYc66|=pT6#$=}N=#vxu`^!EQ/%J)xog;uHO---'?T}}DX,}6)|Pm"AI*<3bN6@A+!?Z>TB!~6'B'J;W&8Uy3#BV~FB
N\@}v?Ea[	>waoVBwp0{Au(!n B/_c<jc-RH`'&qTlC9"WI&.M]nX'TA=l4Y`/K(pNUQj/rTO
#m+Gn
:yX*)m*BN^qP.E]M/T,;Ti4b?iV8VfJ$9gc*YZUv~io	X>Mwk/DDdL5;mt..p2dJ]gK8By-vFe@9?;ilA=WC.<g[WR
?f|
UA{>USAk_\`a]rzL7STF]cBMNb+"aCdT5bag]|zS:sE~+e$PP]MDbQQn`d]p[3z:&5;&Rw&b4})w/cHH5,Q	aM<YxCT;7.}`=YS%y2U7)UjG/{xRg-|Yb?xK0Jj8q=P1bP=\:Qm!sdRpHWVY"0s&5p_wG<FSV]t7nYTE1TNt#?oo/IykMsW&SZv<F'KuDf{BA
X
Y:=
a~8r5+&(
S[M~Bh0\ES]'"j-n(yS*ZlT3==A>9vPcvaUZXG;3CMdI0\ldY(GTe	zs']v2 LO^PGXt%n^A~2>T:,_5M*/l)E^,kW2m8Jig<	V?;`YDxZ#7*(Ri,=%lSkdL3dNq+*:M^GV6}\z.,x;R_' '0j7]2TzLm4S\W/VKh&&+x9>|POS-VX7^lLMC0Z&pH nTx`Xo-/wrdVedVr_A~5wO!F@*nZn(IeEo=PdW1k?8jm4PnGep\v%|3x5i>:jDghiP~4=miD#M^fhP|YRm-1?HYzB-rC06[a!;A?eP}hOPZdb*Y1p>bIy JXw08")`JD~c73=q91
A"GkLXQ^K|_\17k4c-W\YQR)k~75JZJw$7h<e&ibu*q}FlbkWo{H0rJ_Rv+L`7JAmviA@qaC!E1qQgb0_r_y/bXL/N"Gdlbj!tFpj x!1_c&Q?YM-NH90=4OI{C9qnq4bYD50E'U*s;BMZ:@z:MN<8?SXa#kCR-^P~kA3G|VBr 
;6PRXjbFz7XZdXj1RohI6QTm]vAc!L+txm-|"XtPVr#jnWg65>Kx_4'pnHnL$,H8h;D?>K|CPngTsaMq)OCq%7a:UPK3?
lKKa"G|[|EwQcMwV#jr?\c1CRn:ULB5}>>qaO?Cw#4X*QJ7_k
Xu>|c"$~hT_{8 gVOPx \pKxqY
\ '-GB6hHq?LYfMQVJv;8k+'7K-u3k7"{M2IdZYSs#<9<51-U:{SoU
gL/hc`fmw1HK?nd 7d@:soQJn&i!YyaX;Bi!&61Q"o"Lh$}|
:!X_,
6-sX8u ).m@DB+5He[D0z	Ij+}h$)\wT{]^?FdQmqd%-El_%<`$'^<C$?ZSgf]-Nn@R!>mq/<TM4-jpk(<7#D$#!}:ZT\tr*aK6^WS! Y+o*rsP%vdcIx>_y5w>J~d:d<FTjP?/$p-#{Wr =V{q.ow@/1-M5oILu2<.	U0l9Gb/_\tb%-uYxXz3Hq[P|%fSBg+r0bwO%egO1'bAZB{Vw$=#XY1Ohv3Iv@q=WP )eWbo(O0W^/(+5[x+TuN_(KG"hnga1/W=	2 j
1h<3D@.G;yM^~8+:!AKvmq|w5AGdtWy92S+U-3~UfFH&J.H:-oEAor@XEh&zMQ@Hv%T$
.PYZog<z,$h
vJa;5zP,FP{VLtX>'"_3'wt5@7`tx7oQZOk\_nq<6q,+h({p/k.vYEiK"xrk[v}"6+;d&cOqgn0b2"I;d_`]7ntg]/I(O;+"#Gi^pEx&c$O;>Ve#`RoLvROQ'VORpZn5!ptT8nX"7vP2k^?A&<K!LxH_C}r%s:t-iOs wI8z	<g{JOb!R4XfcZi{:<F5;4oq32+??VxYmd]F=x8hq2-2k;(J qW"*aufS7j?+{iew-@g#2</
2H2RJc=VD8 fP0qw4h)z%[-_+Yy#fW_-%!0%aAD<E	F""l#gK&f[k"BO~
Mb[GhTH9,6RRRTE)}AO&jbk~!Sn+s^MIEKX>@V w(#8IZX=U	F/=;Uu!VB{2/=l[lO89*do{q=B"nwU,v%n+C)\y/"Ozqd41f$tgrP`)SRf<h!*p/#Wg	ku	[c'O=}&#"1~:V(O<-oj:C53hvwrN1X)Qbnf|<namx%xWsqg\gs~$;SxMDy;:JJzcf_[bIUXgZE&pEPM0h/6	INNs2%uU<zb[]w%0z/2>Ue
@qf8-xr1aIX-CPa`W{[KhJ5y~Y=pRTn7Ln+fI0%LQ]|3QMtTB38~hkz[kH2%Tc~?TwJzH;0qj-Tjpl$+hk$|R8i*ZR?(s!*P)8eBoQ,nJYx[%KEi-U;$FNMWT+DHhJ#3[	wwh|_N^Zw:SUZW<|YkS
u4-@^(^tsk2:;Q~6{.$f"{+dp^TQt>[M22N,(D6uuU<]1_0uL;)F:e7
0N^e
~:#!=x5xVIjLKe}QE/'n(5Dg	(/{X2NLzVqRc@?X r<7D5^?q;k#]3!9XGBqF_#,-k3eJ-T$:^&ZG<c5W,}i!s6c[ds??8%*;\ao:6Xf$eJ3b6)DITz5ec;
KoduchR2J(n&]<O-)Z]ZQn9H'0/p/#/(a|_2]Bb),(iz_6<X9f)B]4EeigG[M>D@"s#v"eo:/I=XcnIc&:W=DI%/{"E|5k)8C^Iv@l]|*9H=A:=&u]~2T*;mLF\iOj>fb%L	XQ1r@=gD-?\w~BMloQP7lUQvl(>Q 08lEQw1,'.St=+QZ]{b04Lcox}.=l:o#}wJc=DrNyJ#Cna G><64au}.-L!{XT<`^$ 1V3F"@Q9l^{xi6dW}<#i_.a~XhnD\Yu"qgY*Q%<yla]@E2M;nVww6l3!z=NDb9@r8(ijsusJw1BM|6/wn>84q'^}wI60]!e,W%73Rs@*_JFQe}U%\$26nh!$(Pu#}Inzsk&Be=vpM"<a}.[n+)?mI?q=bOQ<_gV/54xD*1ZKy2k$F/g:F6twE5h0B~zlU\}yR-=n{}YP|:C{X@Y&?8J
QP$@61LXh9~%)y=7v F,R{TMi/#X`t/c4ZETJi/k2t1n2ln<A+}mV,4
CbH{~DOHo f%&\aFYz<IYzdmcP:GH'NaHJ_/ml*4mU]ibo&Su;.y4^#<u
Q DjcnHPdtA%DpS^c5']busp%,iy-?>H{k4>:REfB2I[24dQer4}%8.OSVD/)z;s-p/=9?!"nYvWH{*.U%bQ+>	1x9miWVZ>#F.12	 *w-`mD]3nbJ B&ISB_TY9dOQh9=;3^;+{	B7,*zK-!2+TP"!
3
l)tgTPljG&5{C,j+4:o!Ee[qY%k?sNRr1rQZJV83;/D?3_-0|0G<kP"CusNo!lJ/iRwz]0!J)0A&qMxz57* 	N*& ^YA}D,.iCE?>zK6uI}kK6arJ*9NaYsUyZYSm4qQK9A+:Nm;m/B4/$,X-YWOFx?+j~;Sk@9FBJ0~{VZ~);653CQn@J&}H>IP9<HZvaR*5aRl8KN8fr	&8I\W:O\U
|-%fr1c4k3SR7$M^tXmW{D[bJPMi1tU}L*@b`
sgot;$?IdBk[$& 8K@a=b I ;2NhF%Ert8!>C(Z:5S+.L:,O~"XDk`{]ar<NVQ'`Co5DLe)1r!y0	T<b5AIE}tUsky2Q7H'/M?2:R}V.Ocf'&(GG \"QM:S{f[`(BU`NefVA&KJ%HiCDTF#h*rCpizcA|fs&rHY%UkRToO+Y6fx6MqueFHC'$t|Po)-GkN<!k7Vp"'1/W3}+dj?*OK*XV:<DqFbDm wXv"5?.EMn}g"Lvz)6zRQC{IpEbC6A
0k)W~1RxR1{Yf`X|Vp6mK$i&=L[\t0vj
c9lh.XK{)\3jfh$Y^K'n88pTY!U0UP4{<@'LSjNk>+1 ]vaks3L@|>!Ey,9 lf][Ut5Sj^SzVAe
:L80r(otEc>ctn.QU^uM
9|7,Umw>IC2A/rA+i4n+[v|2m8	S{DBp_X=*em&ewJ)OHqoG]QN2x3Zf#vk?N$HcC2bnS:wP%YrfkN5h78dWq`~V@w)	~/W@i_SNCAU^$9-#J[QhA+#Lzb8h~f6i{<^)=GC3KgXpw&|<73091RV@O(_PHTBfY%ulj3~2Rl|0 #b{$~.1!4ka3l,lybu"sT|c#.g_PU<(;cbz-W7sfSngXZR@k
vgK$&VG>:sOE#|xhp	VGuAw+Q+#:D#IcP270bU]~t>+u=h)\ZY4-x}R{pV_D8jbXAd>`
t-Os{3gc:;87',"OdG&yaFb>EZ5iVp]d<G,y0R}BjG(Oo/!
]1^LiRd3'AnI@pi&a~mfxn8,X6o@]F^`9_Ihf2m&rH`@l<m&OIX'Qq`cPgs'-a~pZrD7F\dJ}6N;t=d@vE@6u	*l#*f c6Zp<_TM*=3\&xH.:QChSB!a/+;QG^!BI.Oz:wX&[gL
gIf&3}2~[B*.taS>Vg+3-mUWL_)>4syzD>#n|E	?`9Kx%l$\^f&{;~G\C&: R#u{K_iYP8qH(Z7v1Sk3]wn*:"QcVBuY9V#%u;."NRQ7.xQho'wU->"rZ=%w]1%}BW*TalZ_eX-MbV@?DC|Y9Q+}}B7Izo"4UGU	 Hua EyNdV>KGoZ~}?P!]R*rnmHy,s5u
*gF^%+hFsTF"%j=cc|&=%|#X%..*/5~d/8)tWZef{F3#uh*|M!
Oc)1$g2><}=\Y)H bC?f\24yXR4nlsoMr5%ohBE"0w?=d9j+2~)80T|nh"vanvAk#!e-7EEIq]gC3lo-RlUG;3QH$, ddd.iZ#Wgqnq[*I`M7I<_gJJRI$4AJ<}J3|ACiVHFTc3xgd95ErYi=PB3)x-a@0I@\Tm4$^"kp[LlUB+\r5TfaA2"lp}`S^/k}@'2/xf@?x-^`q4'*@5os(]W{"u"S@?s)!.|/2=Z4p~lucLnp$V5^\=F/h*]c>]F~6qZsr&ZWNY~Z_\wE&LuV6A}8*s"#kAh~8?kIg~u)6B\w7
3)5&y~C|1wB>O0WfS2_Y[!$uwbX!zVqp-3RS,PM7TFLM^X"Q-~>7\r23L7,PpS6B9TlDR9PyG4fN:8{O@F|wwKFsmP)c#Sl[vi+N-G+~8?\NstO&uX9O_)q"6gLT'u-;:]Ih6<a&tH-C2OJ^.:*D_a]jQHw-:-cv95reV\8\0JV=("v3cFi=XXpO`XG!HBN:;Box~b&[hE%[+%nR3!4pxqq[7XfC/YIlw:a#}Hlg6?{^v8/^;_A^6,T:Cuyw*]EpJxu(XBdB
@l0)pws7{h]N5D\,N/_/{n	NC'_ZZ*UkX{O1NJsYr3XlTLtKnm.AI!E)oJk8:rbBcTy?,Lm4\t+o/>e\-n$ijm-#<K[>ABQeAo7g6BF*'lr[W2G{GkTK:x=$9e`4FjVEr	-^mb~(-eb,'k/e_BCEep>M[IyiP+K{-N|g`/<
k];6oN7Vf|Y)a$"o]{9~jes6)h+H'4=X:w[vpYroj7#DJHvFoymhM%	!}Q[V|2j!SZ/7hr*e)yh}Z0xNqF*`fgKXj|R:uKmVycS\&/~J'KdlX>`e/h6xM\Q\O`>2ywLPXZ
^jEk?xF{+,J<6061Iuct	&W$l<<F1t
B:F!
:U=M}J]A L!1EY-@*B<|Z%-s=k@bJ`]GDwYe\!%,	lil>w=,Qh\fs^i'4bV)9][rU7X&fbL_"5L)d;&i~$k$Py1o8f^~[3
%$`iScy;du/x;/,5|.Z>&<?k&"JHxA~H1friAs:%)!sMNma[R7Jd F*z8Z=M^Ve}-yt.sDKY'WN7^#GHVVm?fnkS&kkIvoocdv:_h$iJiQgHfp4f1>)5?_7a^7Ohk{:lTMhTPzh+4NRt^9A(l:F'OV]s~<=/AB{ZfZB<<T!>K-\1_{m\i+~IQeYNvmqq`$lhj]'+<J&IB8gTP&wv]Ta1n"Y6RhYpxsIUGp8[eQGR@OzANM-8&_AoSYG[@_lB1n7Yd],WlL& 12
@gn6ON+Np$><.s#{q@o2_3QK`Y~VyseG+(U_RZp*CMu| `RYR'}soVjj'gu3brj^;2J&^}
00cEl@1mOnX&bkNp?}d3z<P[kylst\I;1X'aW)Y1X'|3TCsv}Kw,>g
f},X>iTE+_f\H:\5BSK/,_:qjWtRk;nYa9W<s>9.<|Dalma6t)8!j;_rank0`g^rM$p-SUOf
6;UG&CByW?fNeRL%!'R44R|,xon:sl}7$3.11|`M}p\;Cf,gYw!p6~.ev$#MDAxqePY<
D>Mo32cz/Mb~=G#!ZJ'My&Z		A4Z]|&4Q%Dedt/52qo"@D"I]HbWh=Th	\KD	$LLgmvd0e8NM6RD^8c!:|DW$1\GOOf<&#_!C$KvjzWMjo)[m#vO	`%<W/>U/N},7eGm]X2>jFp~7,>>:Mj sGq0ltd&Sf=u]&E}qU'QWoQK-`^)%c-?MSC6Q#tIp2|dt7
4=wH<c@921Uo(3V&j8vwyct=Rv&P$P!h,k&6n[D}DY_Ffqf9	F=xmaUW:FDefb)]>=at*%T55k	tMLu/!lF6cAi	}/$ed>NeG|A$3kL4IU:'A3yD}{?+m`1lSz4JU+4&C$=YhniZCZ@6Ql3 0Jv/V#v` RuEZL@L>^U4!bO7iEIBtfLW~:u#XlZA{H&\[e*U^;V.583#,	fP89kbPZUzWMo=6C=YN&H4Ta[WeMR2|$k-.1Doqv@gTs%iO%+t4\c/d;6Znmi^c7~@?UV#j-AD[4*MyrSz?p[0CJ*wwu24>.B~DDu;E`f;<]!&u0\mvr.u'KzUAvuLQ!pt_kmAtf}0^KcH{B8,)6$h&>$aazWi|IUMEa@EzD#MgM%1vSz;=<R]32@6`GB_eBc!*}<!~%]s7:66KZw6`<S8v/FVgzae:\mAD<6#Fo
V|elY
PCvPw<L9-ltVW*v4Fj	MR\D3lj_yZ,i}B~[~+cFw 1)LRHe
tu{T!&ol`\&f-O3Vs`]q8Qy%rRjis|92n2S6wUw&fNJoZe5I/5#sg7b|S5Qtw6wboio,li,]Y"/tKnO59hf vCu|o3D7NLzK$,dotWi{)'O'}~MU[z}{AZ`3K1KQ-H$f9
n.-s27a?bX[!5N!Ap:EEdV;Ls_zj!0O^qDZKb,*m_(S4q`{_$|VX{l4a$r4=jb{B(7,0Dqkn/9"}i+ccaw41h{tH-`9yC?M5aN(
+IT1]+nh9[UC"DN@0#L=TU;VQ`,U3p\>3='{Hc}BbxkunBAF:lxE nSB$3	WJ9XQWVC,rxiZO"6uE;W}\e:'1n	AZ{bq	
&aL\,V!]J_>x&qV=ZBk^*?U4!w*B<8?Mo`ZPsmdO<b-ubJ ;OFF DS8[BI0Go[.O&M>eOCh	`aWc$@3/ZG)\iz8h;Zy#@'t<D(4~Hp@caEwMMn8\{gUh])	?Zl0xd8G,.^pvWg@&:igq;LSz.oRSLbgj}rE_lGc<0E"X(}@~k)40+0.h~O=6_v:O|fq:"FIFNBIUqkjL_TkqMhoclYauCJUP6B`+:2#f vvDk#Omd;-U"K$S\'`Jib=EFHtfA9:rhZg	MDGfq
_N9-oCNL2RoZ+	<hOTuTM#v.\+g(~)1;$tc,HF?gp#nPgI^C|b~sZ[W~Lm<=).X'
!3\+DZ -B-![MqBEcqu4(ux+M9;\nIQI3~8dXex	AN~)^f1>sbCkI40RqmykB)F\zzao
	}Ub`x^%:jyBJBfQdeX[L)WPZ*N6 3KiHR.AMbhu"^`Uj$pQ u${595]7T[gBoa6NTN4EY`FN2[h_QfBwcHvrJDo%^w9KY)N9ad[u/L'?-QIriDcz<S<&##Ng@x|=<XBK^&|N}Q{+O?:N<{&hP"K{ej?uD7 ICbXvCBr]&lOH/t"lo0-tH_e?}h#6
12n[A"ZVMBm_byEu[JyDj64`37nmUn9.Ed.VUX7\jSNaK}mJ3ARVwfNh&dg#[4 dgn;U2]sYTXrx5fB}Hv5{.\"]KTiW
qH0rvR>)Dtxp!kSc17wX>8$
';Xi)6vTO~/.v zl)GQHhs[[h{kz 9Hjp3+wqDf={(}?Uv_b(zT*9#iSC2"$>Yw__O Q@=0u/OVgj0UvR=f7DoaB{GS^^p[w^ekq6$]C		X^	Ej:}mi92Et@
sy.hDA=G)6'_'3Sj?=TXbq#l:[R&^Q&{ran!Y7Z.B[^ZQjIFsR(Gox)CWzT/2%UPjtB0RK?>5P:wrj0/+CYiQcR^PA!@4M	3YYD!!:2iM%4d"H*.2Ti\^hZuM3W>_L:Q!Dxw-q%f40dP,_mv&;(Yzm:}]F!q g8$Uq@.DTA[/j?t 0_omB2DB	H-,H\jA+g
:=.q=yNRN#8}p4E&geo+]MycSNIh)|L;]+T`Do'T[eUo<3FWC~I.Gpl7k?S7ut{DIccp]q)%%O&a1=_siQ[FB(4XN?-x<L;";GK+DZp51>fS[\cv<(&]9mk5P>9t'`lO--2R`^(cn_P>3CIn~wmd$4GU^eJK~6{Qvw[%^^%s4cE%9hrr<0yi[f%J'K_0iw){~CV.1\ACBV3Hj*:.KlPYDt@d#c"b3EFML3b)b	,"4y/2MQXQ~VEy>D
jJ3n:KJ*\KJLzM }IWe
n;78kJj6o.#%
!,<|1/+0v>B4PUX>=?k#IG7Fjd*nna\ebK0|35riK\j[$cl'lEEspO=Hgup] z'>w*D:8JbW_y>>j.~1#W~bu"F+'Jr"7/$YV[j8B|Cu}d4wTgaH?}w/;;&i.O,L^l.#VC;*'6g>Y#|< tgSiIBrM{l2YB5(T2W9XfHFm"Pai$FTH*	`Z*}T*%CU$x]f\<zxdE]/r#V&8u$OuR7ZM{| xN|aLKJs~0+.q^kW/@{&IEU7]2eHzCY 7{
\5E	+T_US	{}%/Dh<ta%8q!e3]t{F[2:mqO3~mF[#FP?_dV|%	&`CX?^'lb7":ZkuT/~<h4W g"N3QkaO]p	gt0%17C|g-'Q\VGTGQdy[;JwxT;gH]fMlwM;l3u=~T!j{
qBxp6oR&'V)`*gy.:Ggj(kN%bF[R3 7O&v<?HQ^`%b-KgzzR{,`A|;\lyNr#OX=Hs:Gl+j,e<_"nJb*'b~O%]aQw+$04In@va6z!|&%g2itGcT~6]|!X1+ix&w8oj
g`Jo2[|.Ytar}L7*-O`q0rKa~y})mb!o
<FOTl5Lv:~)
AQ*i6x>?`J3Gd {.n(
Ou6YoNMZ0J6Y+wTAn_dqU5'Lu\=<eiTT@1!HOF(j$"vJ1U|Ubvn)?bmb]`a}Aiu@[OCQBPDQJq|]YZ!>s/.r$P`B
A1]yfMwD4\OX#t7cK]>MV63k{kr+M\5fB?Ky;g[7#Dvh7t2Hx 01^NEDCKYI#SW[`No8BYr*+K}bepp|RVMV]n$Vj#hXe/Z>F|n'	eLu,(kPBsLwaoS%)<s/!DP#0Njd* &|f:JZ50F,Of0YmMVj*AM@!sYuTX2H@5y?T*qj6
?89H#b~\;c?eS>"5)7?)Dbq}{+z`7wTcaa9h*F^Bp;5<4$jS/3N_T7]+y:iCqX%XV[Ia2Q$Q9?<^75x:i5~Fyfz{}:i?l/VK4GH|e8e?o KR9SDFE`j(Ne/JdV^bQ"7i}%}oArtkey'x,N")@A^$AG3^0g[^+`R`x[NbhgdX]1dnf5y.Zbrl)X=!yzs>gFTD?
a,*s{|Z\2-r;Q-;7*?k[`4Ee(hPS;E7/|b)K]lVoq|Cj>bO1'E]OO{+N,.74"<&kY_B=XY4(T0L{`@@X1|hi0X?q_5]xYy/fF2oNkZ ;["%O|lN5:(6,zL&`"(1nXtrbD5xgKeX%6HW'<	$Lh.Sla01V;wQ@Z5LT^]	Y\Q(59DWB8Fp(AsaX9WAa&M&IblPeYy|&)/Qhd	n9*`wd?%&wR!xhEIHg1B@Ks'n}qjr-R]_B:6pbO*OBvQ}A5%Gg!r,:>"03!$X;=g\SWtOgQyT
N(x\h_N|F01&.v9OeJ)Hb&*_fOfbx~T48dHrr,;O1/apUl{?uFTEMDx@g:;xl-hFobikFr8J6Tl}F=cEF.	rI1{w7D[WmT"3)J :r#_QYPhVd?.Fo3)"VDm>x>]a0=s
TTA~(=OKri?U}v\2_ZQsZ#-IO'y=nUYgr5U]JyJuws{:W\#x*
ZLS{cU?ZgX,v%kKCO;t"6M
KNW*ZHy?JS`E
X0	P;8}|YyuBHZX\sb@zdk1G
c1=)-ug`
c]8`Q$kLz:ZFL*1EIa!vn0qHS/4g<	Y9:Pqma]P"s&$b@1
Fu<Y{!Ea@vS^&w,"\f.jZH}d`hC4);a]8C)%t$$yQbOH*gNWUynQLbop
\--
f78R"n?,Vz.
guV#
NG2@hZTzoN<XSQd=["K@hEvp<"lDED6%1Quaj.--\[]La&#Ok2{\7xqI:F7"A!Pf!Go{7}Sn[%@VtYaU}	[.M&venNF@S_nFDPgxuabH0~Q$DQW@Q=ce=@POht9,<!LxK2$`kj
(vPM]A=IQo(rxar@?S/T3F8B?'ff9(O0<%rm^h-o0os<nG0.,/<\Z~NRGh<HPO)V
SC0U,c-0##j()v}4{]Koj"@O4r2r>[D"8mK]e|mf}V9~[	Lv&J?=2<%M+uu$V)vHhL-A"-F%mgl'9dm-)6^rR/[	uu>5!t@LH`_Z0Gx[Q>jO/_#wQ_ tvQX>YO"m1vvF#^o"h5\4q*"e\uG2$shHb7*^
f`,#*+/ynT=4>c!HoE@&"8)ri08\JS6KHm

2#jylOUO^:lQBJjId	)VuY s/Wa057BRmpPm.mhc8X[GLpI6J _of	S\=rrO}4.tA2rtsu^\2!eB+[(:`d0t(V[2rQrT)g+Nj`|9E]Kh8xC2Lu11 ;qpU'8?W!H85n_<XKsC#zO}=7Gipl`}9j\9
1O.%H;?Xmn*&?]CmHm}(=B:ieUM^E[Xl,4Y9MW*wqV]1<|@XVl}(k0>u`#Fj7&e@``InV8,> k4w>neE.;NvW'p7k8}{\>N%"MV8"w:Z'++8Tk0vjY%M6^S?[-YOl~(R_S4T#Aw{RmTnDg#d7DoGk\&McIU*w@i0gC#i@No8.G=>:	LL1_y:JAij-Z.vR{ARZER=s'}r3#9;IqXnwq A)6D{$vu(t-P-:@qx_y/~V+H@dv8`fh_uGsfl(V0mkAJ&!pvmkmeQ*3v&j{1i\I+GFsd5ps2:okK#e.bd(x\ ]_Q5=w7(X:_+37K0q\f
"6>{`^FVr|ff 6u
52W$Zd:]4XB
	J-4:Jtk>XK|?lsB?DB8G+2`sA6~'vyD_pVIR-a] .;6G)o#<"nWu0Z~Y@&m6:OP&v5U>$+Z1${TuNiYJ
Q+JDB^lH."0Z`;BfNGWO~\	@JHn`7P$MkZ	0MAAYeSu\ReaW&LX |tLw2FCfq1J6MX[Tcij(n:_Ax!X6#GFlM@t.?VM<[Kf(7~j$%hWw35_*M+jE"Bu;6blR5bia3,&OMn8V,}"4)7jr/E%J[DxBt-R@iQ5*<	QZ!x]nqL=%ZD}h=E[\I_Wm3<WT|ccDN{?	iYSFMx/h'j\vnc/Iq5I9EB	%fN7'J%[`9W}i4r.FfN[{LVxE{no\LP3s^%}@xiAXaV(byYdkznBldv`*
>\C>cDr\_{[$M]n)rMot_Y:].Ph^5oCGGDIYj3@AY@DA7T-%.6hr%OnaP;U^.tp!Ty"VqM;i'Y_J_sGz*.c#[{iVr.cf[v\Y]bK1ccm AsZbIzUxL]k]^q #6-t alVn-j@Te+4uKI"tqFc8
$Us(^W>"e9R53< N5qg_K>1^g8*?Clpf$h4<@AfU%E1%5PX!xyxlj:i8$XSb;*%fw5zJHM
rXNEX3RORS]Y4YeE##jL3U`t^\M;Q,Sp'S5x'2~2ai5>2~kzv8Wkcy\`.'b^Z} k !"=ZAfl1qSca:]*<D
mq(Ku92p
=,>8klWUQbe@.W5{J7Hv:y\WQ4VI)PqC/x{r8lZ-NNj/;<LwP|WF{b-HM_	3n$iIGX4mDZv+ ]82Q|K;r>w8k$lawFHL{L	nkXZB6SsZ*zuJHJAII@FXiE_"saK~$&_:d+{}h]Ree1zQa;n`Eh4a'x*=Sc96myTg[ <:%eb:2)VA.SDJ5j$`ZNh_-E7Xfbe0&+y9~~pqi#WJ):dKC#9X\oQnZ||wn/
g`WHVpP}\-J-/Csb%UNDH^l^uk[9/	b-_:QEVj@!b/hga	`%%fWX[1F^:e#NnyVD(lD`uY#"v>i..X!JCQqZ,Z<d2KU/lD1LKJ&)`%\ Qy1	lrO[;Q8E,XY/X^iaWX|/*&x&&n8m'H9oX"Vj30 J4!8B"X.6)YJuiW&ZB/`|Y2
juiM7alP$CFEQ//.%W2mJl?<
s1-@I9(bv||)8_6Ig	#(k{gK.+[4A% -}?tk55's%6mTViB"kqaHxXR?]N,2ict9+_$_O^+e33%U9B0(.U8}V!Bx$)c_J.7:y'Pw4w`Peprhe2wu(oa;WjX1gUp4SNFsP=0hx.rjz)ml\Z2?%Gzl|QxY$0mzo|C3'8c}2oiy/$|X V&(}zWxN !_aZ_<0
+
@xg?a;<VWa.CagUpN~8`{t/'D3+wqA0P@E	y-=;Jk(| ;AP:GcDK
1!G`M)	1dOt=1qEg>4(r9"PcXB
hM;WLo2vW/"sdXHi(69xMZ`D1kU>=d=2PJRGL2HXpK)>4\@A[_Fu$WE(%Th3sUO	*aN:NV$n'v7|Uh=d^lhofV*=g$+,[
d+?(heAcv"l:rQ
wTy}BK+
(XwV&hv
Fm)yiU}9qYn*p	Pr*qA@YcI"@LGee&e~	6ft8f}6D[1A'*#)uZLmj8j{6D`ZZkr|B++aYT9#UdQ<_Mp8I+<M5>=t{)T^@FY0Jh6=?(OnI=l/}R%TN5@rm%
09"Bmu>M05YZS,mr.+pN.}A{ (Dtc~2*,iIQ*&FC1/ms51dU@)wq6mIN;~RU{G*[\}.8~*e0<gMFaL{*Q fC'KI4v&pJ^.f(PH^cZ*AhlcMDBB06SH%3():ZvZY\XCU>[|zj2yx,&!z[qp<AR~roWDDoUqV,t95:bUpn%2RS5|_\h'3c5hs5	KF!"ig[|vOUW*|xb{u7fPkRkyK$EqqJ"2ehi>,qN&mR(lVmuogn#]D$,:JF[H7W<;{WrCe7|L)cEAt3:~x`WO7_dLGg+k(	pfT[+;t3%GL(]oaVKc5v	\tyd/6xzCWGy"	B4h6;dvgqIBNgof9_Wb_1i%'tS?yi@Yp#{)Yb7M4NX+'^+ V4So*7-O:&	8g}s5`[#54>/	l*>&o.es]k<^Bj(HBcj=!_ik_6:4h3)	/uI.,;(hr{C+?cOC#
a&xO/eUg4G~&d\V%123Aa1!0>x+bW\PYyt)g#VWFUhT<-rH*XyWAEvDuOi<>^l=CO"%~H=KZW!sBI3MLj5EpVq^[eEL
|bj<etIi5Dqu~IlsdZ.LMCf.+.[Ra}eml<4]2';I=J^=,uqm'%aEy'\KvW%YKSMbSi_(s7#7v!r>H"1*"=~]y7{kgAz.mp{Y$GHf:+Fj/8n=%>]" D32/OWHRP7.6DS*1LzisSp{s{VW
^U=^Vwe|=?_;<n#R$	k4u1`/guDp@Ag}.Ry`ko+ua
N*"$Ckh%jh{G2JI}deiaUQ>a5?V5<(uSCU-BRj((D@'Q_]d0|a.3Mv@-d%=mzi}y-88n4xVJvUNrD8(yx]8ha_'m'9oFE0?kW2U)p<g{h-GsUAzhv	b_<YEnC_Tkq,7p'@yxdd[pw'<$DAqk/CIY|Vc#:Fy"pO=+:. qr|0H'yOW
<1D|>-6T)#0P1kyV{@n<hI^LTWXI!DOZjNW"XJ9{kr?n}Tq}ozWY^LSrB;b9
ID;Jl\6Xxm=.WtHW6euZ1&*VU.`Ft*TNyrs,e$C<RZDJG~+b'9C%PTue\|!45bGo"QG@{F'PHc?F!"/JDdljRe>_H;f03|&/P'
\}RRni.7<%K=$t:1|sZO<9QxF4?)Q#v3kH8Z2'[)~LaW+I[j,LNP37grF\}pDkcHi/k?1)BJisol'fo/5%/@&	'Wn^Lf-Ke
4rN^&@rFEz9oOj$}dH 	w+5GLmO	nANQ!v<1&N@2+B7?	{wC*5jgRg47kW(oK`Y3brlL+bv3mN.s.HbRhx}6L?$zuQeV{{7~jX9QaD{n%.XLzEa_Ppzg9k"Ko`q~wYVG~81"qjfisFr1M8[5r{_@F~wffHV:=.QrG(aWb:[{-L&aAR	mnT82_Nb}\guo9BOqg-R.U|iG'3/KM(y,P+l H+%N@Jm	F]G@\i6(Ab#[*zzgd#+&^?#%iJ7pG\$P0!Q;\Xq;\9nJDpkb
+[?jJ9x kHTf(3{0MvWff[h-a[*~|'`%[O*@r?5TAReqJcE~pK`0>Y+PYBK3TzVT/%n;SUgjaZ$QM{$@*qde|hr0[A}@j-wLI[k.(7jSW4IQt_RSLIi2IW'%H5RmyRI!H<f4iD5S\0!6c5l;jS,x-z<DyLX[7&Gt"AGj'i4cX<W3Z{$EfSk@Wpn0Yp}dUW?o]pobm;	E6ipq&A!$zu:NV*EhOS{>R#wtb*W)iEZz]GJmS\Nv[1kqC5++^x/)1MhNV2|-d{19[%fT"=Q/-)$1fJ
0x
 vPxEYz*$8+}Dt\af#=lY:T
B34^?dg`B:nT)b2A3sm\bH>oJJGhykH%%]!0@m|e='xIu?enfEIq5oiH_W^XeO!_=?_.37KvU:'GMc8Jt1)Xy#X.tu:"?e5x+B$QV)uTJ*r?3sxml2oq4~3l^RN'<6i[h1o,IWF;?/bI!3(u&lW%9E9[jSiS1K{Hl`k?Q'cj@8y7oRoeJ7ogEuPK#n?8J?~kIh.e&@z[Jk9""UJEhm;C8" (f=k@mJ68b^/D-)zzW}%[^k2.$Er!-,hw!G-\h2@|=dzk(Etz$.w*b9G%{ka6IP!Cn|Wg_otefJ|IKEZu6FUZvZz@r2cw|JmVu;[lU6`hY?	aY|U.jY3/qeK0N'e}(MG_+bq G0"BKBEF@R30Yw_?;>>&$a-2^xAWZvfOtB|G_xW`m{VsJ^
?< 
L9?|JWN~
[>jU5S"YNS?/wU0%e`nWW~$}XRW`=R
M).WLTHI)Zm1tURiWYr-u|Btzn|\g (C)$P5JUR|M
,X=qK-VR.2"N6uBHEl7^_JI!DtH][`W~QZEkJzM[GRY'9A;&"1@hc=l&Z-^g9iiB4J%1m11_WnOr*Jm~"<Ktly;oJ"
UgK/3$:"[.p!3fzSzM@(4u	+|BPT&^@5+P)Qh..5iY[Y4Eg\sXuJ rV^%u2HU|m~@fIFIWcm3QC+^HW`M50oaAu`J,a&ajkm}brb4;CjEph[c@{A!\<z_8<tP?+K)$R37O2q NkNf"CI6}&Qo<NP/^C8	+mYPtJ3R;3tt\!\r3nKe(v"Y{0z{"44B_Vpy}/)zHI.xX26d$=jJAn:(h;;eaRq)E8:lXt0ON\O`&8s2&XTy00;'7pCB.2jdU|d6Af+)}HSfkMwa8}$d-;DZRmTX_P(%0AX9o)Meccm1=g7TsG57K@=jiNvze%!q,=XF,KlB4zVBhf}Dy@nJt.<KH9rN=)XD$SjIG[W{hx5/|TPJ=SxgQU>Mu4~71!NL-ELE(@`vo*T_*b-8Bz.CDa%,%]4AXhA3gBW`W{9:hS2!n$BH7Yfmi	=Y\pYteM#q&T;",S{/  y2Gb7\Q3Q%;?\BeTd+N rMj`v}(#]m1:mgM:Us6_O&wGy13H4_8"'Cm*"p%_sOn"EmQj'y{6y"Ge/A;A:9':]q_\sP~?gL
^7|a~&a%]9K;+V/5zl>N/@@ne~
}i
mLs2hl2}vIuo3?dL;o%0 ,2&%rz=Bc6?^wD=tUTL)]GPf/D"IMk|)O:$@!27~1R.vz,]h[}cF+xF*<e)ew"pBb[UX(.U
vUmv{!thBlZ)s<GiS;H<k4"ShuR^hG#5ja>h8e5-hh+vi0{H4g"a^:
wHSnT=Dem0QR,1.u[WST9.Y%<k e1#Q$e\\BriOMzVC$WP%25rR{$"a8, -0joXGdJ4kv*[
oaqDVK|3p\&.FV7IdN	S|.3V	;trm'5pgtJmN3jJG_0QCpH
V<U]s
.s)$X[li7"*4k%3el_Et$fBvL+CX)n+zZC	
j4qEw"ez*%LZizY&,Hs&uPs	f0FLGSV]h=k9qssF	xcr:f)&rkubdPkh"sY/]k^{,38B+OTSf4xEI003m?+yjqcFcaKWC>Z[: J7Ae|XLGZs|b.3]^M(T
nbyuldU1l&
g#p=IibS`_fbG`-%0|W 2jO}yJQjlq!fCoM/,B
tEz4pIuw	IUtP9t$@%zgu}%||\k"gTP*`5}5~tDZ6SMC7cz/[NPgF2rxNl,#|n_:N<.XDY;Jf|FF!KE9fT_wNWU`!=2BRbvG.@d tA@_''6O/51ug|u>wp	roiz=1MZ8+Kx(7)]lM{*0{b.zOJ5jQCyd8>C0|mH|PsSza5D1Fq4*<o;WS4Koyp<3fgb_}_&)w	6q.^a"z$55
@nA$3X6%F%&R%,C=FmYF/&!DPDB%_B|Bm2gH3eR0W\T=+\^IiHM6M<Dvpx\r`=vqlDcR`#PjKu3GF\Pc[ iAndx4j&Lo|Z}bb-<2Fz-K7:@uES/Wb$?fr+Xq'?
MAN{sNGnnA`GbTw>&bgFS6mWt;:n	ztLQ'JpLnR=IT6W*q 3SIh*A3J`1#THHq>F(l9;Lk&maJO&/ao'"8V}B^{V
`pJyJYT	l:._{o9p3Y8l
HP[hyuzS_itgI?C@v]O?0-?;'=KXBL48k={(b-& gT,'DgvN>G=3"3y]V!ZoI#KP<.5\P~pv~B
.rO+c^lec`eonyDu|X*BLK-MxU\u	,]Uc@\I~
\1h_Q{?bgsHr$*4B%F1\E$p&r%Q%`K&`uQxKPNn yV8_]&oocw!k>^PsUaIoIe<7:+bWr4T8nF59S:#c`n?^aVgKfz3g@Xw/[,lez|8ei_.h]PvV)`SLaJxz>]=XhgV\4}!g@;S'tHzvq*md%\>=p:=4/=>+I5`x}MuR`31l7m*)hGTE0Pf9HW;CWPXv3`/@~Rjz@r;hjzu-*)*\aYZ/Z9O\p/5\c$~.p;r>0E53,F8P1;0I:-:nvJ/47vozkmR;Z_w3>Mfc{Jc*poveBe:ts\n&[T\_&.M G]N3(0)c
va22&uVFs[nLDvPOepeULJ-lY-|~XTRXT<2G27j=B}>y
tAET
6G@rn/qfiHoHqG-%g"jl^>f`a}OZ2A>2g[}A/6-
65]<!wu*?`)F`$zx	J2-s'*z*F*_J-XDoQ_IQ{z\KpoPep1moaZ{a+C!17Q _Tz>hBGvkRgt-~{I	.v;EzeoD}COu](EV,h`C}
j QB<jU`7^Nu09TQQ|&n
8`X&vpABI;(V2,Q3;Wk0P8\{\JMXMM|jHRXq:|Mm$oA7ZFePovB/V+-QIVhj|Hz}K
Ydb}RTj:GKM5g 0>,Y$DmWI	ZF1_98/h13D-2QXVse/-o'j\.^(&J3\X[:xgp&Bwm@|A7Cv.eg8vE2$`Q1xAPa^6.kf2cCT|1b3FW/occKT2|U.?9[{oM)Y2z%+36/R`'pQlK1656Ow29$#b@>6Io.mYpE<K@,l>xyKHluVHA2F5
ag=sCAjRc\LBZ0gC6J"KEwJ;Y=pa[X],P !A{pvUq`USu<MIVkVqUbF_bOePdp0>6SgJVIxM=Pr4f:~+<lyA?>KH-R}Fl

58QD%B_[1.z`l&k-2r%| AVG>JI9X	x7"&v\Q&nRn_6u\Z+GbQ!imC=xz$KS#Iwj#on!a{b(Tl>aPO'J_>]yqF{i>U	p>VQR}R$m2-`Ry=.%%=zN%
b@MK6hW[<x$*[js%V^/$ia+V6	(e^;HT1fJ@Q0
b'6ib
B_'!)84+le:&tK	**Z6hDm4
27yIGno=f.oQv?=>#^}dkj8nJ$>5,J:y< ,f!E@exieCe`pz3zvZHZ(;}5kN3V I
MF2hQrhT+D0oG61"1rT8&M9vuv+Pc&.pQHv#s|m@qQCLK`@ka]2cyJF=i5=g"^z[%-s%L=St&PO@p'\'1IJ_``2T~^v>SWx[zWzL?`Bph<LW?Iu"861B`H9e!B01f6H:MG;C&^egu	?m"ffR\k*v*IJ^"lpmB hK.3_TuM%<fEN}QrNyJE$@F""'Sb<,#5lkHaemjwZHI)i(znELW!@Ia&56wl&M
lx*xs""}`>#DGdRkq@"Zj}QT?b`boJ][	Zeao<H0P=jIUx[jo]/fQ#7pG8w)i9^C
`/g_@YG'RW<R*3?$:AwoiSV1!p_BYB)c.(?/uMK5h|Wy/=#4O0}j)th|u=5s0vpu7r<I7P[1+sepY#y
E&_j5{9+
aA)?qf~3/_\`D-l.tGxyFO^Z4L$uIt!dieUOA|6";nkj"l4+!1P|/$rSwu.wA3hAs$~M3RO=|iU1y$-+=e4i:30!R0Rl=NGq*}&C?,-6urg(JZX-K2d0ETY<=aj mP,%"`zGu_7n/"d1Nph%IZ7BgaMR_82(NL{8FTJFKB4y)YDpKe1`/bDi*tz0T%PO^QZ\mC=;debX-rG
&p%,Iz\kI!:9/9s)K0e^eAchVt$[^+"4l56?R+jDmK0Hqk:<@]#,lb{cwi2] cFhLt|DcPHU&<_zk@hYFy,+(aWqd{?|IxvSgME/#Fo(ICwA ;a9wcBpqu-q=6NBO-G`6?i&M?1d31L*-72a/nG@z[&W0S',>9y*2b*?FtKTX)tf#3H"XIbj:rb:D?/2jOW|zC"h`}[`	krG Z<2fT)8Vczb[A-"T&s"*qj0%97MNZ7H]wp`[71u3~t*R+V3nx(LGJ?[e-x~S:to68?J7+R,ro?bG=a<,"~ME15`Q\apR9A;m]	]WdO}'!Uy/yWB<j*NVWr[9^WC5.M(|	R'h=
5n#qU$4/j%b<	L9K*SHWWJnDg%Y
8pl8S#qg4rI(deM-xi]1.l[p+U]q^uJw!2.YC{4qnktP|0!%9fK;N4P<=	]jw,tI@D]q-$qQU`| 9kv	y{X\a?rLQ
@Y`dI3ZpXvL;4nGqTm4Jqn%Q ^jsZUYfaR[t09!'0#MTeZ?+Vv;~X+aB*C|A2F{v7E#+mq[e9HgaSDBN?Q$Z{'\)FQ8@86vA)N,j*u+pC%9sfg[rs~fVR\O1BPe86-*eJ?*jy#NeXw2?{3<Tbio;2,MN+(12vd\)\=<bzp+ 9gTos,';GQH]ugn46`)lZXUzrN9#iOkZG/\g	/9 z%"]P!}9"WgPzR|wkhnA`}J>7i!A8*C7j]MeSeC.eCuw^Bv%M{ShvfWbH%OV:=+UG{NrL!K5KCL8G,56<|t.&u;:afPFxvj*)-wepoacT:G9CfsY	
RCCxPV:(T
\Qe5
}
9S6RgC"Sp1d\e/."WKLx)\H
|,T9R3MenfSu2a5;?<<: ^W_/zf1Q@Mf:b8huvujaD@I3k+mJ$]\~PW*;UdcXOzxB"hHAZTTxUT"_Gpw{PC]sV5^Z`bP=HC6T/WboyiUwOmK]'4	UutJ]i-dXjJZ4Rlfa6K~[
}nVL|:T\S2G4B)OKVW!w!A6<.c^eb	vO}0,v9'sArI42We !sa%bmSWDTjF"!H|jGK@=>En7578gCT~V(.
Gtc<QT1\~Got`KTAOaAh\Q?Z{5%9'\y:>Dou**>B![kb)|n}Y3XchRp1f,H9v<Wnf}0%l)e, KK!NgQ<
Wi6S8TWD;P_.!Sb=/0^3imiOOJwJr)>* eo5o,j0V.ZXm
HdOKBLItHd
,=?i`M#'{mNsW-Od:mDY}YBdt ZiRIZ.(5\j82Y#Ed)Lk E,x^g?^Gv{Yqeo"aj(8@pLV(^`'lb<s:@MX^nn}8
_40y=t=[;>i6kxA^Z7+$H39 F0qnT2;,il2r#0_)7 OXhm	.MBgOzzbugH+/2}wCG.\;F.c4JCanS+h%v^A`6No[_vmF#+{3$T]KFcFT:$y4DLCH_}o\}Z\/e=-|89K&q(}fzwkZ}42C+h;	K/":(nlQ9]=q#RIhz[[u=Na`V3s#2YeaRc`\zV05P/4F:$!T1x:Cl?@ZxX57GV,/^gbB=	%W!e!YmWlnV'Rv5vGm&C89M"]&,/6^X-6.8&w9)KV6$W!u^m]DW8myq{k`SvfP~555cgn<$\RCa\Tq-8t-J,Mu?6mo;J6BxT7x&[
B}N]vD0Vi -%?hUoAp,-
EOb-PzHl,MWrA<1JgF	9K&:o0*;59Ni>nQ
:x&_	i%[9N-zH^;R|avJz~3diJKz, l7Im0NQbkO}(sE_hsQf	kKJ]aW7=j$5#@1hD#{
?HQp;(&m>A1G;K.S8
 =QWvf)EH`5P)=lo[{r=KphrIRK0&!f_\gAF/8\R!2e8gA'g1kE/rnE!a9g8{^fRi_N4 ]t}l'{C$tB]=}yT5?LRVPC<R"8OvomX+</P"-NyE[C.i@gFg$>`;In+tymlOUC`^<wP^:hbS>|
%#8QSx#mW}hR~\1b~NV30wcS&ka;R4-mulGE"eZ6[jQ,Df%nXZ-<Y*!pQ)@D''|iX;!-99R$G'2r(Y\(`hK`@u*2MxP/pFT}JT-zV&yu5e:d<QiF9t:7mMI/5!n,ps%A"Rni#a&""6h)vvIaCR*TLzzYnCfp&*NgB(hmdY0yr.RBuSxEg<z$mk!BCZ99}`*jAb>`hU53SB
C_v&AyEtcnUf$)D-#h092SmfIz-W0joFRkxv&U8jyO]~fYQJ!a 776U7m<Ko<jc:o~Y<Zd	i*.DWcC@-80F@lq]($Y
}Swo"2\m:$B+{
2:5_=aF4'`KNU	\e07eLm<[:rT:[}8
xS#1<:V
32]4)hHh{0:"yWP`*5Y{&<B<2*mGh0tp#u:&dWCluA\MAkthz7uu$7Upy
i}LIAZCe^}] hy`DX+Mp|54O`esNNF<20_T|v]QCo'"#^&Pmxlq?M:(:~'1ica
It+`e_G(p7x
eCDdBXy:%0d8Dn>}?ND+/u:'2nR} e\bbv[vG	@e,^.f|=W;i
yJ'iiD>koWu_vR~i6@u!Qnz7	[xT9l*I9)PR5!$
yb &afRr!q0esOf-KG	X`#3NIT;- duLj_jaU;wl_y\#G{>\)YuPlc_J_U\Jv+L-QIMJ+b;@/Ox!iW7TIK$&U<X|ddsX%<~*dX?gWJlRP-]mNuH?dW)2dY:8K4F3w3
y~,<-l!o;NQ.}I$d}mYDg9jEU&*dXvzT=tMX+'Q3?mo/jrRC/\q.~!2A<"3i1z9)Jd!<4cjb}
S3'N+^6=E
VvR&dV|AH-e001GNFUV7d3y'a-8[lNbH/E1
)E3 7`@op8I@gnvG%2LxF&*@L8)&%(8-s(R6,q9mvoQU/9Ia,%<rceTq55PVH"*{,';S>IK2\R>HbSj}"<#.M6F+bPsx.k\9z=;m+6"}Yj
Cv&db{o)*V1	G'"]PLY?mDc'm@vbhK) @9^rz%U['xel:\3b!#u,/2ZGcin1\f>6fm,he8BfY=MCtUI]U|$T<jMORuYTGi?QVW0]#$Jd	lu,bsZ3W9qjKkBX#FDf3#XQ;<hz8Fa[hhaj4iPqch3k`--HyxY~)10;MSSZY~4t:2Jl+zF/:nCyL;zy
*h_Sk]pDX}V?RU!$PU|$8![QxmHE6/aNa=8cm$X+Ih19jKcA%C/h%-b\Q?<o)4!#fLJo=#2!1\0OvEA0{h*#(Tr d_')@#Hj%2\~F\btvAX-`L6Q1Vt32rK<H9FyN.^'o,k21#f4kg)9HC[xDtzj8x@]=e*;<!n4^a3j	>>e;bGb\;q.)t9Ha
6jH;ef0vl1%axU~.?bCTD6[>J[hc2'y0s4|<-EZoDBc/?{*KL$B
i>0xHuSq92/jh	(xhu~RKK7&r~Pn:YOdbyt$NDefnXYF<]B%A<^MpE1>7'y	vE0 0|8`|1q-?P"M|XXz8*`4wRU.mis*NF>m=1%T.G3pi8(b&&:fP/2vy) 3/"USY)mm4]<=u*7VL)PYx*4),tb<&A+qeMK}a_X1
N9R$@f-(ep7i7pJ6SbPs"JLS.iVI9k:Q<z^1/}zb!#Aj3_W:8i{#<
 4,F{K}'+XW-gZl;	JV=fC1y=mKi{M4@DKd\zc,xX`K };:2Kf}7|P!cV"Ai1[	F	Y"D+&l/
qP>MaeDo3z,Qkfc1%"gi"S\rU|)X-0`,i&g~0#W-dwhP1<AH.~@G(Dmr\,5&vGUNnD<I#M@U	E(L?\1 $A>z0dfE%dQ-{{a	O>Cv5BE8 Ki8Ogl/rA@%33Q,5c^C}P@/`cCva?w*f1F
1%6Cw[D/X(B{HEUpX"ngdZZ`C:"wTh#?hl}dkw*(}?%YV{m&c&l'l}{BAXBA iif?*7QI%F{wl1j	i#\ms/8f1r)/eGr%LIOHz43_-.X83/	{j?WCwh?3*R}%BXsJd\F}gBq`;,WJBG|vM.(zix,Vc9fQS/s?FD^w[~w,{bPf`$;i
E'c#VSiU48N8yuWg[&Wfn-0s3/6h]djf&tGd,h*hZT0- zODKQ]l%AF"Mo^C)a	lrAUmYDfkQbe`9,1}"MK?4i/Jj]P@0=MK8]{"S~;7/x_!g7Cr3S!"]NEZzE#2pZ3\xd'al+Xg~#N#c%4YtbV6WRc6cQZ,wpoYmf=rW[7y41I^;bixm7_D(,	`d67s3p0K}#,MwmY4K=Cs\}bI-ucW6Gf.EoV*=[PHwOentG8!@>>hiJ#=|rd)t%'skA"+N+ilEs5)~jhBT#M
qO/8G=iu<1;Px-Xup+'*)BZj5i<sRmmlQ:SR~hF`JA'Du>&,?4x7gn`Ch\fHg}CTO2~-M6{j=U2U,/VLFm=JL^,PkJ|{;Fb51P9LOGV*[#u#5IG\8a\s+	DvHEjd	(Bh9oF4I|uLe9pM~Pe(>|
"oPp TVlJP!B,Lj&u7g}JKf^-vl=(5[ 	qMYzuF9fnms@O?/xHgrbU{+22&zg9;?qDo)>L=-z2Tv] fx`
/!,xzB:5][{vONvL[Rd+CsBvkS4ag<2fK'\S,KD%KIXsj}Q)3ZD:ZB	C
nC:#:1ly^f,+I0w|$	Q^(:=Q.]?08NKyy@(!bylX.$D)[rP)9E2uv$#Mk_@<2^DJJZg:S>wUi
"qQV%d!2VVgM{e %y1\)N4]2s.krr5Lj =/b%]6q2]&2_L_Dt;^+:F4IW<*x!S}s.3C__=ofX
43$bc:x@j%GQ%~(&iw_/(IZR.uSuuW3:vY|!O!3'b*+jHsnYzId#UnCy&024"9)
O ?Y{$5LfN7hH[o$H,Oy+rKc|vm5fI	2UyA`Pk/qH{HX"%se>;{c836gG8Xrq<@v80i{)R+zl%NRPskQ4DA2-9-g*dy!i{&u{-,D`6LNdLOxjNX}YOPF{Zad2Ch^l:VwQAid/[ bya-4+3G7gn|b9Ii'I2D^*ED@Z,`c6%4:wPtV'yuK>%,fpMUSF|;e'jzXk^M>%dsL3v<%LN^:?_fQJgC)/{{{iG^2E4eL~)/ukK,Do34Iq<p^|1Ol,vitS7nu(@3&a+,N\*[?&G$Dmz
7aAe*-KM50gsr7eq7nenM|6]atf{m??i`J9tK{.FPhC-^n\`Zl8L8qtg]	qY{ykVZT@W`he`'ACi?=brkC#97^x`cW8^M%T,EgTZ3v}tB"ftXCG.4Xx'4z-mr;zX`(c ^(_jVL,o&'
dSOa&Vpf-2k~%mDfg&~a]csE.|\NBw68*"q?D"{#L:H\o:Az5xu781I(,4'yn/Y3pN~o!M#;6i^A37C:~R:t X+2P1c@;N{j<@7l91z{A=OIl:! |Lz7|WNC}U*_.T8[c-=cqF1yP+bo~_OIo0=/Nvc@-MAGDM{M#7R'V1v!@z9-i
?9TB	6b6s.BBwGGx$G@]J^=fn8|na_G-V[{o3Q,$FyL<7jIgt(|)Q=?J&x<L{C~I0^gmSZ=n9R*~*4B95~zhC\JBjou(iOM^3"& uD?AV;mttAU2#|wvVDsQ}Ii~9sIG7GtL$FASPvS{kq1=8*eBH#MLcQGQw,E%Rx3MuT(i=P%XWFi6X|W6U`G.I4o!6W5@JR0~!3m+"Iefl`uX8~p^ .W*fq13r<RtalLAsx-aD^(G|jfb6Q/!&J
[ezXl-,M3m/q3Yy<$0DBs nrTJ^SwaG~\vwnWXkSGO%@,6cZ'zN%`fk={kG*pp1=/NTqW(
tBx
8%d5f~!,R8&2*aVob9?7$Mf{wj>tTUG+F\Tvt!mW&>Qa*oU}I=SMC>4t7E I,Jq/HzjIgH^	SnSBth<IXS-xVmT'.1gXuk ]H>>#$2 81c,zMP8T`?UeDcB?Bfo\!4-<7;l}UE,pGRYrg%JDzy=4|x5Y5beRP|nn`b:]\'&tw*~E[2\rk[;xRfZL>[=z_{Na> |Ts;TI^*|
vVv5a:{AbbABq;X+=tt8xb@&MOL0{8vOD6SSJ)`N3ah}liY(;$n57}C
q1!s@x%'=tJvA|?>q%';`K9]%+OP6<|U3GS`+i4I)^_ j<TlCTGRe8S%TwN^zBgG^ZzJ[Ei,imt[_a&1#%V0rRT&}6"x4'A>r_;x'ejLr(oEuC5E_=#TeT'\Vil<D^VO$Z:&M?p:-kyX@PMYM3jG?&?YtbgTRrR~oPV)$8km:(7,R.7KLo!l]6~2nH4o<PR7ytUClU]BRY_.gNTx;;qD!81BZ4na3{04pt>O)$E\o^21L[nC a
D#[fz'Tb1g0Neza38i/y%,q1tM;-0*Ok-81u  P82$L%bkGp+121e([8O^I:5VkMOO}pZ'IG(Lt6J%2|-l[Qy$E@{<Noh,Ags#8vu	H #$cwV<,vz)ZxuWw[~v=j1-$9N@- bZ9:	6RQgq(z|wOYULwcc\i<glNyH$9^XXav^<+<3e?>EU0<fy%($F\PG|#o5v	A2/]x7os@Hg}Gfe<<QYYffZ_~J5T	C6GG05PnP<48)E||?{!P9?$ECRi`jamx_6us6C9&OILw8FK6</$v=d$&j^'p'C;9{S{DD<_}odd?7Z;_(s^m4Z91?s	#x.1nw!ZFH$m{;Z2}izPr)ZpcK%x%f?7qOYKoNfCv;[9Q)vt=DFoWkf/O(Da+%ZK%P:lb\cY\~u@2+3ieMz,Hd5qq8j_B87#4)fq8[eqXD/TeatkM`Q1uUR=YSGeTEBc08\\/*9I,q
qyc7//a^s6
qg6d^{=6
"kM1-BH*c+6%ipBX.N*_78{b@'`S=]2)D/J$KV-]SSF,RvO rZD]#Mzww9>_IYf)~yC@	CMp5{%0g8KsFLOSN.STDbBY)5w(iF8y[72)NUyM)+\a$[9e(^f>_fPWI'/k?q\<>lBnw87ci9O@W,8rSJ_(Q``kLoBlsy[{$9.c;7m&.gq8ruJ)_+*|F"L~	Q)TDC--{E)UnM+ ]cUZN]V9PR3-Y\*A4NS8>B1kfX2pSi6{:R~*"([6xhhi1FWh?moc,>AZU/WP{tkFv@f?b*/3_k9R\
=m
<-'24y\|H0(=o8Po P8'JfbHFx8FC>>yguC{)Qdy "Hh*$V#~\[_P{iou1.m[#}tkDZiGa+P3AS==?+igr9H"W.}L
'cs8tBDSHC$.WH03\#o/S>*7O
!"S2%^/6[p:b)Bg'%JXnnoL'm!M"ZQOHEd/tr:"~J$%CX[vp/P>.'y)9*>r/r;'k)f?qfseTe>qnPq;&(=\ch$XEo[?;s:W55I4E0vEDGJx16y~IvQP5WbFkf'|A'<Ts)c)srx2h."OGeJ8Zuk5}Vw35/2|^g\W:"M(").!~)Qy/`M=-yqrYoz^?M7a Az DX`aA#chp/	V459rV3>LA	CT^N}JF>ti} ndhz-N:I:UyF}71fu%"v!6%5'%oURvKd?ACk41Oxhkb?"%
!,	5gxZ	aoUX>,:|M+VZG+P5YA?JP<3:Er-,S["vv"3*8yY$>{bNJ:gT=<JUHP$,`lbRdu"8Gp&s|5vpo:B{K_:2-"0VeMerLDPp3S#wu],IoHMZQsx6}Z,yT9m|'hBn`] n83]g]WW7.PWVc3XpZ;7l;H,evtxPH4dEzn`,^D9(EUNbGsj'ZX:\PX&gfVQEC:kv?Ub*t99vP\GS<ZmCoNr1yUe&F{{ubEq QO^fdFNgGR#v1@m@_ea]%;pdEVihcC%vrye_pz#br>@M+#i5dr$?V<z1; Hr%gVwK$VN$P[g3.aH;-W{62^`Qr, %MOriY21PqqmMX([)'E$pwX)nnQ)@m3MY@83i4*&9a3\+l#pu|x?<8b5m*i8I*,ly.z<5d]va' 4sbnp&=FdK)^*#<0	jKOm6Xp%(&?%q[,}0[o}o0?'[x.Ze"y=`Bu1ix(71?E`i/H=.:mCiy4@8sFLw|F-~/Ua7e6*NM*j+
%B IH?x'K!>a}Fdw>rlY,3aRoNI*%C0yqN'LHgf^HE.(a0P'YiyEFP1]G/~sLh,23JPC*M5u\OV+h_(GI"'5Pp]wt^Ra=C3%mp`
M0@mo/',X|eMFY4Xcet=&37B5gQy@/=3h	=4YRUb_*EBgtY6<T)G&Ct8TS3[}/$kzV0q"YVfAd*W`V=YaG7s#S!Fqf-~+SS#`Cx;E]=/h,2#mkCB.{CV3*hn =(=R8U?0XIDEu{P/=*q/!4Z@<f ==S@/<yh?76fJx&cbB#k[E6kys3I\r="U%h_t3X[^}$+Dzyrzv,R'eBZ/PAoN%Z`14GUfu(?3^ef1HWGVSlD6qh(U+@csuhvQV<|XrpYoYIJZHfg%#K+RJIzl	eGovXXCHg_'Wq2,d-}gIMqwk$h/iCxGr,ABpDVw~T:,M% 
}Ux5r7r(?mC!]_oAQZ=OFEV:cW>/*1}4 	Y	M2`M,'\\EjVq;Aap\M2#MPlm:3FTDGLKUV1>l.t>'V1:`LEAk,Y`f3ac[%S(Z	x8`M(uZ]#(Ume)dv*%Td>-cO08u	{(@][P!:k;{)BUsw7PkP>)a9"LTgdIp}oWxTW%J\k\!~#Df[q7a60y_Yv#Pv+l: ]vEl@Co2f7
T(/~]@>K1^5z0[3Bf%jJP:&T*wo}-Xw
nm:xNmU\:T"MEfaJ+%n<0M;A}!Gc%Hce
lQ;0($c!"1Qz2ZLw]>[ilFOgd{l+_Pe:=&8QWC;e$>>7hiyi*xBXsl3	EOkQlvj41P{w-1V.5ePTy[>`;~t	fM}1 Z5dEj?3xDPOCz3{Y{k&lW	I/E8$&"E>WzJfV~$QjL@9qnugc`lfKwykkL]m99J#O"=q#3TLo<z%poWXBAm)8a.hLCdI'H;X;~C+xVj%juwKZd*ZxCoRi}|JR3|mE})5	f7ZA}'S~e`l2	e|<CST x>%hoMpsb/Y9Q"S.or.@ln&ux*f+R,3kET?CHIeFS?<7J;j4Ex]wPHa[
;fNpB')RodV:,t-\\B_V"JO1O"wR8-dpl),)U`.`(+W<z1"i7a?C$*|&%"\bz*{I/dho)bC~HWx7jAgX		Y9\L+bMwDJ:+fH[V*b	A,cyr/pJMP	wZDSH|^Bd>.)3 (V#hE_S}LI/v{uu5>:cx&:Q8+%=8Tv&~r

6DF<3kr,<L+|b@mm4ra-#s}Pf-6B?>X;oR5@1S.:;vh
=j@J( My27L;Y?fU%v|.kO)^KcaU?)m_XrcP_73MuYopHVUqn_5JA37tu6fEEQO7d8~T*Q"i/\>9SmD8V*dZoAV)pG!:]/h/cRIn\[_ES(9INK'}l2W+MT\u>s.)h(6RsIOF"g8AJUX::,"#"! $%52z1C;Zfe{%R"b(Qx-"Irj~AB%_-#S_X^t~l1\h43z)vkls,6!iV"LtANd[D6`_2	&[17'q&sPv(F`9=gE	"jj^i\L$z
EWM5
=9c?;:>-l$7=T}?_P3aI2TmA
N^]j?~vH277'tloSXUZHSIx,'CzzKV]qsp^bd=am(gFUe	z[J'b'B"&oDn.Kc?s\NB|GZdXSidGj&w
IxSQ$&M~{OnibW.|LxxfhL~GI'U
)dn+-:fJ@u'S.+pL}oUlzrI$oDD[ h2o^TqVbyCm(YU6X_N@(eqEqc3,gV6E5'-J\;
S)JB)zeyXr;=gZy.w\tiFO]Km/VeN`a4[<L\eF"9':	ka%iAWo@7[/+1.H)9Upi4m-{rWoO?'%}l*a+Ts1`pj%$u+?Bj:e=jk<!\J2mh('FVFpI[pM$jt~DfCAIQOu1K'I*ik=*3LXM<CxU_Mzc=eZ"93ArzclgV";$gcY\2Wkw\[X*`p[U!K_6Po%.={Dd.u<y#c6|{Z[$;61n 6@0<?W3"aC}
?if;5=EW!k2C8>{;+=n%<){]nOZ:;LKnQCpf4ez6+z-RByRo@R	|~r2xPn6/E}JmUK@uMRN{^o74l|e.D-@{j:Yg9	d')8lxJlZwN2+fAD;Ho5bzM2	
x-c-y^y_3q2r54z
Uu;T0}sm|[it8LX\Ir#NPT-)R<Lx1{$ZK >,w |r!z:"$
D]OTU)TeER-kiLMU@/zI-"psv%q)
Sx{g%Mg`90|eZLiAg,`o^/,MkM<`;))xhO;|og.yMF7`F9BzVLgO daI
't_
-x@d= r?Jy~2'#lQT;`{J$y(]hTL'w
tDKyD?[;6iU-^89!\C0.YX&UesZHf_^~H{
l 2G51:)deld@	8JHpQ69jw.2 =:XTDz}GS0&s
Kw26[ueuS.}	8
#%lyYP~+_Y$G}5rW}GinKkPD_h	2.2	Rgr_A	gE%wY9&}-6'Xj:YVF5N9X@oZ	u?E?5kA|~
q{rOv]Oz?e_'],Uef3(H50H -fV ShVyv-2UV#$iURxG>"ZVo*
b
SfbZe)>ovM^cY^/t2OVhy
u+H6Fx?[=]_t^	c|mAtES4) W$_JA^]xU~+lV/[wNLXtlf)T,B(hO{0ha'T:V|cta>Zig{MR;u#dyU"x<lR?44J&+f$a('/'~G/;C5,DyTlL2+)z]Ese<54xdxt?IU\i?p%"z03dUP`IicB6X.=)\<IyFA3 C?41jt[6w)c2NX:EPH.!mg1[qc-N;<%<gB,X;Ioe$]yhn::pQdi8W%R@U5D3Z[iU$o%GN3J5NA$'EZ]%.u@Lcys+viku4[/<P0Kq?7rO(f8()V"7tt-46_f0 lk2~p<t> Gf17hkY"yIj&WQ
\zWzY>JH/DF/OIATr^wWh9WE'.v
;'|t;3d7(	W$2CbHc]]J/4	AQmY32q0{U:Fej)jCvip/1BXt: t0\e5"6x=WP`qsIv<A0@Y\~&Q!D.Q`dDJgt[FHQj0gDWFhc!SFYMq0knIbWC6?Be!I`K"1IiTtWi}6_NlWs0Rk}[etV+	@kqrkrQH.F|!Y3Kk\2KoeO%7(<@mR?\X1`Q{],2S%1^WWlyT61'Us:nV;_7/q.jv+|'mrkH-w&3Ybc;5gYWMk]	7EuC}'y[in{9MRs@24+YLX@T%b/m/	]5\H_XOE!WW$x(MyxmG,LKI",a	1m)<Xbz\E~=Gv}Q}V=.]Rs,<QY:}?A18P5r_[~2W+m#q0Ej~V,>Ge:rl<01RyD2CG8r'A	+!.H6c9=P#pc6E!7mh..;Dz4pQ~`{)#cF%HHZwI:52/>TNYggv[p;g+ou8ejQ.?OC`a<~ NGu`=2g6@`e4QoYAa,b3=A9^!nWMx]K0EK*_i"{4WHiFPn|92/!N13'ka$NTni?'&:_+Y?RN"pIJf"BU0yK,5kL>
~V`x{wHT<ymVL++5Cu,DX4xT`L.\R7Fy|F9[[S[{`u(6,,HWfdCQ?lXLwf>i?)<5/K4~4|tk8?09fRW@v4yH$SQ$7ws%:W_.d,c6Wg'Ea}rK=AvggSPl?f4	y&Cw+}X$Vhr\.#Ck+
(5rs1Tt-=A(z{a-+!T)+8a;PP@Z2-Z!te8"J/<oJ]L=#~mib7fV.y'	_+]W6BN$d@k=B/CEi{RX)d>d7A	MPv"
ARX'/<`,qubSx]
td]i)oyELO!9NkYO(N"cg.U#PN(# x-ptk}7@3+7:l\%EAvw7U*\G*pyPH.ki,'HPSe,/(5V,9I{Z{vXDPvKY~o]t9oUk	<w;GxCEk[|3X** +s	&^s1Qco[2PG8!.Twtw=#-@M}xI~,o*\2`:[<cZ u>Ctv
A]0(uUs	H[nAPgOAR	nxsf6]RS0{
ykW]'^sON)LwG@Tz7	][XS%|\##G[FxwK"{xloAkgj[@F-0SmDT'K6{(GtYpZw~GQPw|9{yz=$OJk_YrV..eFM*t	jbca0O+a*T#eJDuvD
]ziwQ=32D|%3)Urh=]b5a$\KOU&8sI[Ol<FP_[:^|Uf)>i\pv@&w~<&% }ideaWMsM7eA*:V{]u#Z?X`{?!XyN&C?WKNG)EwwJPea.=OGz; 3DP J~0serZJ|A{|JvYB_]^{yJSFY<L!/#NX$7X	y1|3f?:F=:.|b@p3,1<Yj&'bfP;I#aO%gP,`%n"G2wz1hAYqM10P[#kujS/|/2%/ajKC1T^kx~e.ugzI0+'Fge-&u[.LYOb5:cv;k1DW_I8($}ECotdY#:%vaAQs)4x{HO$BzkM7s([WG}<7 K}MVT>)r>[p|xb%bwzB@ge_0U
TA-Bu.n.3aGA\0	Mq'g*L9rkg5XC`cr\blSl%~nZ=|!xLe6Td:=3U	eH*A)lgA85~q`Py,B~*&h@~r$6O[6z-r<\x)BE'y[8.cS!3QM2U=wJl\XWYfK>pG#v0}QjH">&RB
:Z2=|}JfVD@Xscg*lK0=i5@r/V`-;7D?c:iarKA
N0-^S]>sKNa7Fft\q,g?fRA{6L~3v]dqqb%m's5_AM4}1zwt^>k y&Kkt6mfam&j!8K>Ze1'2v%Atp_ROk5OgC_6&2Fi"V8$Ox8mCiV')<DM9~<F|-qvMB,"GR(6+GM*FJ:`5a	e<4`VVyRO,)5a9~.jO+DI(3vQ>Ftz`?L|Y:+LDWrHZGTm`d#71X'F$
FXnbiBJ@kA;\OLrzX
/Ip-N9B<RL}6c[(xnk>VW%O{PC6I_}sLv{KZR&J5azeFx+N0<ddq}4pSx&z+4)EU#X%DT=g*ySTQm9&ab5r4HR
D!vL0edF,k;B%f.Cm=W;~k,:NT6U9W`#>pLEwzN=r(}'ys0A`	1D+wBVyW$icQy6cTND
j3D)#FP{)7X;S;s6V#VM6U<L<!)d2%vc{L|r;uzxO>-dX2By86|e}6<bnQ^ ZKW<v@b\cm0=vth#_(U_k4kLc{QRAaqnU]`oaB{[?>Se1:D]+YGk/$vOu@(ML'9a3DFp:x0&!o`y|}v "VhBgOQ:6zxm_K47gIPAx8c'jDX@g:{Z,iH*&mclpm57^x=2|HIV3!<K3``<|$|,_:g|Cc!x|pysvg}t.3#eyp)k:DZjq>y&b0j698[g[I]gVYvg"Q(
rxPkm%KICe7}BXsOMC*lM+#)ggb]AS41W,EmG>T	0QgYo2Y
R>l+:xrV7nqB3LhO_S1WxUR8N=&vd-3geo!KxglCLwPmehQD?nbiHpNiKf=[a@|M{\eIc'
 2h-*p!k&1]>a4A:L|e-./^/%V #[MOe}_Dj82
	1J\`'Fd@uC cAE29V!P6m$Z[q,%X$Y}d.@+`bm;5<MXyM*Y;;DDBQpzJ
]/ub"/pvJA@24P9?	Y,F^^I"XsDh@^fc2F56\+KVC	h>?W3wCns88Hn.J BuE< ;|py?,#^NIlUWhpZCk&>FB|eo@Mh{F-^R{2N]#KkB}/"k5 `@%i6(]kB1xd47$o\0Ad}d&	8{/%3a1yYkL>ry_B,MuFFCS^c!&F?0XqaRy[}ppqA32#%Q}&}W<Gaq=aALg$rarfUi.ws*RgyZ,a+K{V.sJ$aofZ?Qnw5uL3*XJu]
%I%y]Y\%6zexIeONz}cH| 6UIlAzR:KX3o9|sw
>5Y0vGzhgYE6\iCSkg;4_"xT7T+$Vu_[ac"/K;Mzm% }`SA0V_DA82#&t5egk\8&?`JWnY'5'vVYTZiuk6tka}[.aFH2ZkT&fj3*!/WlX!GgUqP%$]<T0;M`bQK>Qv`EngUBe(}/&|><U?"&]
EHI6.dJ4eHc?y+(,]e_!$rbi.[7r"r[P]rWEi!W^z!9`lROa$,^AYzXG5KIXaxWAk)*?
_m$E:YkF}-(KpgswHgRFz>
*:h%wN,$e/8}qUG)CE<t 6K}#uy_zl.ovv(0u`sWr9E|j\AZiiT}Ep,B'JEv:%dp`mF.]1%B\SP=j_MLHqe'qY{i?3c<G+8
GuaJ:vVn_$>cW~VG%PJZ\Z%WV@U(a).(yo,0JSkID~c
v*>s#y!`7_qf&q*g}EN
lUU#0}!d+zb';<iC|9e-r7^#W327y?,CE$c\8SJw2#/jTx4N%"-#7YBn0H7zvk\t=jDW@u;#sEbtNIYY,[oRtU
2()O2~P$\wvp#Y.8l|5J2{4W(?#1])U&a\>)U*, ,H/N]0otR69Nc~l@Zb[v!C,HsR]5#8WX^o2C>6X4!M&CD\49O\(j2kZ!ZjB=[J'[r<`q3pt1ZnD/^'/8M
l\?X8t!:Wi<nshf[qsv=y"F Xi@9QRsp9Zje~V:;M)1FUh{nz(le1N<{&L`K1416*{<}=WmbT=.=^$>gq
U(R[OhKY
\)Polu9X]jF/YVWq$Q;]$\]o=iXMA&;,CR5]|_kfk"$Q]8Pw9qairojvk-RCZ(fm$<G/Fn@d!ed]rt<[_)y Tx	:wI;M^9+vF&vBp5PY7W=kM^).E\HY|z.2|.BC5VX
T(||Vn#[kqL79WISd>~90~D1)6Ah+5d2Mn	avh"FjV4&TkdOs?;VX,-	nXPv,1Py\%).a
zfRA(8!y8=+)qtf@>tS|FBx#o|2BOo?+)=8rl!,R8OR]#kXe-Ju86a&Zgu4!KxY$s-l{)r5E_[5V:0YcQg_`LS$O3!/*l$	WktDfz}&*]uZay[`:opP!VsY*v:`Ngdrb^e)[t|#,^K
Rt(GGXbZ/J=LKemDypLVm`5q1{jx3=pZF}0kw'CC7`jYB=kL#C}YP gNRN,
A[{(<A+'WBm8=no%[jNoE;c\8aS%a[hz7SU4<0'%&g;uY9^!aLEUak(%`g>uzV;++}z/t558aW}l=rrmx|H$S-+V16xNTU?jW{6O&{35
L0W<w}*[GS)C)K<^#?@cm~um{?Q,H $?`	?9goBV6k]	&+J26l\	&8wlUr7m>}MULJ>O`&0qlEH'n}]=K	
lrY%[KM{j|q92)Ki|-w/~1G^_hs!RjZgo:*Rs\abZcz'=JjGcJE,<6S$U0cUfd4V3[4yz3%LrO>dnVm!yzOQ\3c",tT(\u4M)g-otN_SoGC-	*<!a!n{t3JokaR=R2&]E]Prw
^(Dv1p[9Y@3U+ 3@jxs8|24`[D/9TAP*[1IRZM8$AT8)=-`8%QW%htktG54xdz"y20Hd#t^@ba#/}!l\ZOQ$N'y(.aew8622<zNB2m*FV#Aw.NS!\{#'8dx"obhfSGAB~I
ta7#@6y03uq@aD9.pnl.A@8xz1"Ys2]r]EwK_Yh?3@Judc?D~mBt6o@-k7T1^,r/>:d%E5=XGH*n4dc9d eVD&-rRE(,bn@R{DNx$!P?xV7L #T!`,o@}<-*l<^vs>MLW<^wd)x20u.d$%x3{d6c/P	ycAnO..eYqOV*:MsG87"9feVZfpJ]!6Ov+[n%2oHAVZ=XdPSkhE&`j3Q\n7{Obz$V}IND"E*!KH.Gn&1+}Avl]wCSt<B!-.t3YSo"
3Du|]z:\Q	A9CA+HsDyT*ULdxT.|Lu*'&Mj&Pe1<2,z(S5N4N<WWo40=+WjKWm}>5Mq>XsSHw{pWdgI-oo*"D7~iX7;wRMRqXQ8X'0T#s?` 	..$3?3st,	S"?=_qIgtRrqE [pZ
brM[304IG/054(1%u$@q)oLW$X$;>x	so!6eoT[
y4b4mA{T5|2N(PD(-=;]wRGJ%`H{At1]FG>	
E4[IpzC8ecea}4CV0Z0F{GQ'\G{CD $4F<@qjbN}G\;ZZ!u%.NiT;a%`D[}
B02X9#J.%U!fY7;vbjC|H_^36H{B)p/qnrErCuQjHf#HI)]691"Qpth27`$bP"=%mc]x)()o>%\Uc.>f{W)|
/$"4Q.l|J.L09==RztG}\J&F}$"vDJP)|8A<U'Fr@Q8y&ZJA?itE1D$V8bfsq[ l)7(p684kFeHfQQ'Fc!Ce85Z9c6K}	XswpsJV8|6A/X(xv_D-#"?Q8
tEsIiFc3t4MHCr?lcJUh ;Dfi&U9p;V\$x@24'&zp5~foxXqeo%"|bS)a[W^ZR"(	6tud<Dv	$P{aN"Id9GK2&'d&5i59;1GSfa(Z+.I:zz3|~CK\*fn]Zfd*	Lbtq:m)bbD)+P4IuF}0gsT 3EQC,)ydE]\&@U#*{,Ema5Tgv<!u$5Jo7G;>tov"2@QN7#mC>>dFRdf[ 4}syKfN	!{WtEs0OYzb1]9iHM61x:oY	d#xw>^63pA_#6b9C!'O[NjPGaD)!j3s^cELT#Kmyry*p[cM_A$3DE;B{R3_759O)f#4;-\o_vfpnR|7,CXZ2.-&v+=@AT|'DGw(`a"?)Fhb'>c\dg-rDtd1=8\+//Rr*\hcl,pDbQX*S#v 8O:FM21Qvw9.B(+MV{Y*3o}']OE$k4IS[WE6m-O9W_+?E55Q|kI.1y"tsUzhPnl"1$B=WJa`Ev.FbS4"Wv+_m@OE0+aTW"d.	q!^+*=Ij?T>}0:#(=4U"aGbcC{M{R896*((<Ou ea=FSbFh|.qk[XL~C'H30-xB<oN>PH+*}:Yq)X\CW&mT=y+wXnmrY6Gd|C{li-hhX a'EeIq}
fx8K0\b[{by{XK#CD40	RrUYkrsO[NCX:jPG%v.G*0WjV`,RLu:='>ku#)w0L]9/gW6Zv_>Jmebcl_zmV\I>axEmY]
m0W,m"'gnE]Zm[IZE$g=6Ws}*-n@ZG\)w /^z;\Pk=v`:AeoUb /46JK8cKEq&u|TGTOZP#:wt$|\H
ig6OmX]CC
1Rcew@!\\pt3dEn:b*{lZ@Z?Q&Ufh3j1{lj&P`K>[_>p{\@$EqOd6Q-I^&#;CMBh	g0x[/M.yg^9
H`C_b|"5y`DKQU38Y{[p1-7zTd^SJg8$o.EGj'JU[ydf

gc0YP$38$MzK5khHZR*(gP0yoTbR`ze4	7JVo;VD|*r?phgF$?s\-@01QNJeR"S0C82Po2,@(o\K7%uE2Dt_/wH?iTlerXSQNo2&vvV3org*|5aK}
p6+PEV_YQuY+7gR*m'Ic4Jb=f(V_-2&5=vwJ?\|iB`2#wHLY$?AEb91-j1b=85NhzC%|e"bDML{I?PGz'AAr30jm-<kw?6*H=-^?l}
rH'toW@QESYcAh?!T`X/d%$d/XCblodp"N-RZx5RS	bM#?>\!cfP;_oH
WX&,#{E
xL>RevL[dL3UJi2%0n<#R-n'$13Duw#*TpVTc=D2*,~[i7[smdfBE)l{
Y[RcS`MT/<;,ya{j-l
=vir "Y\w@ty}0cEhY(vsKswca#N\__m8TtUr`RNLvGmNy,zIK@nR^	d!IH0\NhRAkqor/y8_v$P}-G1[K&Q/J"43Wa?/AF4@<w<.	If	tl	cuAn}GNv_V9=UYE3.UJ.#V;23:jq&f9laL~~T[I^/Mh
+-jb3R`D#rx7}<!JU0B;A9T4S:/g3<c@\ZiOH-}2$
rvl8Ykw[LCni;R3Rroh>(6N=7e&	#>J}`HqIvOE^XNwY)EB7.h|gi>V27G"Q1	CT5<wsH^vVdlDK{&%v`Uq'ZcZl6gKQ6RSVpqF@,~V.3A;\.4-9S4$Z^5{h)[|%GLY,3(ytq.o4J*QLt-t!&`9Boud!(7@k%?1$0BO"q'.sdIw71b@D(a.OK'@<b%bmRJCYxy|Ta&7UG5K.Z%erI0QH6=3D+%AM_+.ycMKD5S`q'p7ZxhaY=~a |bX9eLSn)4=WI_XfSCJw[*^r-n/A{_t]v>x<;AX/+gcI!2vu<YP&KA?pR\/oBK.*S^l_1#.>>_"Wj3Q.ckVumh
-h'	Z{<"?ZJ$6.'P{.ReybuT<0+])-~b9=m6IGK0Y8[`L(!*t&J;\ *.R2l!lV7wE.PT+~w,-H6"s&Wrpue)~El#uQ8Hxw/u%viiyD-
$xmW^[o4iW`jO\Ipv]|9X9.|0L7MZnAXJm9|>C0cj8Xg@rvQIezMB&=2;3:v24wafoJeNsZ%oQ3\6f|m>s!0x=J%bU1P=x5J0|="WWuwp2=@m[sc(-_fp>qj@]Wcxdx98sS,''iA]^gUJ0;^E^P%*"IcUMo"z(C*G$$%~'x'Vx|\B4NWT8q,<iA<ZA=(Puu5n{8K(`#nMSO.ewV^k_7d]&E5FW{]c=5z7_/<8H.1wu pK1?6P|2k?Q6qm/:0uj_Z|-|_1+ba~KC\5{0>V`C+s?mIX,nKrs{RlyS
kBYrf/'G%fU5S\xT2f/K`K[uu*QL!Gg
<&>O775Z}czI`kSM`4xWQ:{k{&bq2KJrnII|_0"0HeUu]Gjr0w'ay-b?52n2HPs@T3TqI8tQZ5/mZjl>K,;6M(>*]QNqd(_+2<13'Y|Np*5H{Qczq:G&&e j3
rgN~l|JJ)`(i9zhqh~nL5zY(B6docTa=jK	MC2&jpCDIBp_ R73_J7">lB~x,}0^}O*U_Cn|:7Sr#~4u9`]LSC hM1a#MXz;ERx~m]T09i4)TNt;,\;S<DT!UG*T?/jZPb"{ZYW2b*L6<1VPCys6IwR!r5Yk5+(Ws@		JJdBv*"
Rc:ybm4=Ej3/#p!J<euFL{6
"y5kZOR}|ZsT;^}F!k%NDCb"R31ub|	
d(HNlIAh^[?RQFC@v_,bL/dmdYru|@"u=:2x8|.<6CuiJ81mkZ6hf1zfRPAG>IsM)'A4X@[rw^'ySuM v=K6bvt.@g8sf)@}eTqbeOD8'F0a?rUC!e[A]=<(Jn8XPx);wt-YQ1>(>^[.&G%,unZz*Cf(L;refiJ}\|KL,`)gqPW;PFv!2mk&vFMl3WQJPL	%zMssin9f/zZL)MFj	)RAkS\!U4o@F1X4%F57;DaW_ECL&2m-RZd},'R^wv;dga[[kEU!<WAx`7C_+puCr%Yb)y(Gc?J%)G,{JFb/|B'6MM(K~T|Itm+(781#c,d!dY(rTXx
d\@AzIH>}'@^>b83cQG
cV;/K8?DW3i:brU'-SWH$R6'8|){n.uf*X.N
)ToSIeT#=PZZY5L(Uu~Gcu'Kr"MniyYx"Nh=+)0NRpU(Na=n64Jqn-nwJ	gw%),{yFt-CK1Tb|_X@i|cOVDp2sg[2yt|y?B2FI{
L9,c-O"]kG|n1VBPa[6-|p-.tdnl`NL=zS/Gk_*]d1O?\s&tF%`qF	}M n~yT\}DtVM!}DYk>Ar34W@{K!Kjyy$(tWefBYi%^&uQJ/Ou"n9O"7mBN8#4I=iXN$9cQJ ,Kx?G.+Zs(P
H`G4($`@@XlpQx?"4h(p"$5}q"v\P|/[hA"=s0/Q96gAPvs;zUMR$g:19A@js`6?gTqT4}vWWgvM0b1FF0KI<qvVWH.:#ZN\V3u>A5kq(<HUT|DB6z9%/~
=%'O!NmKar2 H\3xl)AO.~vxfe/=.gY)%"F|(j:nb
{!FPg&	1NrX[*yS<vnQO;/m0B*!N,-q9iS#.&CVS_$k"EK@f)ZyJKWlR?7GdU{52Da
bRM\}'85Oje#]<2nbeQ-[AC;hE?^VTJm]tW"#(@9OWY;HZowv`?FeK)d	_W_}%Ty^_:@G[%kxEIX6JXv=]*c3PX_Hq,JG+&IQihoq7+YtxN+)/ <*Eo!3ZzPSf;t8
n+coSP:[{9k"8P5~CMn
k;v56tYp&D_u`$o-t]f
G_*s,fK(*k6Cc%mN;N?#~f90ykSwc9!$z}kNVJ,:|MPh8tX.SD*;T4=+Nr3Y]])l%<="'~,=7cQ[7Sqx@P	>bq230+Bw|a
!ly<OA:%ra8/FN(y%-I5?om{|ZT/TuZX6{PI;m3H5c2)vc~	,]2xUQ@rwy1fJ1?^k8jK"AZ@45sKl3&doQ8i2	mh/q?kTd>:,c3Y|h+kE8:r3^:M
c5yIf1k%Z.Q,[gF]},@dmor#"+Z#:cC)/}i#ykH8>Ncx,p'E|z;;$d;$nW7)>a^=_A%zOK$knfbK6yQeDuD)78|oad&P
M#Qm(A`5A|an:[]F6{"
uwK8TPj>fTHt8o	w#`f]*4[{7PH$t0-dBp-1'HB%j+!jUm7_cM*MP,H@R&%J/p-)gAc/SBC	^q7Tn;eMuRNJIn-v	;Y{bXuVfb2Jm*Q$$F;K'/SOv	Y3CxzY{	Exk{G7I18uz
l3/m0?5G=EoGa5J 7Kr|qSn\4o'e`MpJ3x9_NW`GmQ#*,CISc~8QlI>!pHE^BK{{>/VB1}]Gdy$B;jK*|O}LePH4YsUEXcmI<$R/B!5$9jGUqB_Yk*1ryztvqPKlS8a0N6]tN}wi]+%h^aKe2&`2^KzPokcu8G=H)-$F\p#TQ?a)257Uf)//?Z8l
B
65_ddYp5Pv-k0Dp_1<7kOU?(NUECa:1K<uiD&cV|/^@0)c>;+>h`>r3)}jD.[x+vV.?TVeR8zYo44WRD$jJ",,tUX55.=:r1su9.`P| H8q~dxiq-uU8Z!Y?,BP09g}7eQXhV7go#=Day.0pz,[_7xE_"Cyrarg|7H_`-FpV<uJu*&GWolxSq34K_EvHG=r%o3++xWJ=w |\?}D[*Kbj~~m'Yzc?/y&[y+R'#O	I4vB /jhC[Bw5
j|rx+BM&aVTCDLA}XCtUF*3z#wDf}DQ~fBy=tm+zBzwN9M:nr7>	LC96V6IKg;I"?2~kxOrwaU9WA]LHOpC+0I?hFf<n5a(55h)t,d+=kpg,(ek//g-jOZ!pg$F>,!uH3^2,K~<mr8K3x/	IiB,#=h5k
;[Q2K;DqfN4Pj]6!2[ud9I&8dzk+U^C]L!U& LYODbsx7EPtDCHPC-Mi6*0!Nv#_O9J$I}q`02WNU#d_+ybi$U++iS&$+En,ydod["d0XS?w1fk(FT5uN=LSn1NEISj^o56&QE>efT8!,`/]1T1Bkp Q"|)|dm>;O}">4EhYEj0?#${,PnT4H'HKvQ{?"
t/xd8l.VpWslA#JZYE:2<?)pgas<:d\Ndu"b|NWv0Mc:{B\Mc(Z:@T=Y8W5fye}Ew}lg|H,)Rz:UeSnx#NlV`d%8~hs+EWC\jJ#kfO1S9<X7%?~H9SWi]vd71wp:kzlAj?L2G6]=#o[^fyQwH*A>niT)$
G(9EoZ 2\(OkhM088qSsoi($:;9z'O_:C_e*gjF<8&#`#mE7>*b8{Y) D,i)T/%Z$I\_L}VDd[cezku(UO:~o=\H+_i4x<6x6_ZWI5W	f:8dvD70a7	GUFkv{@?j.70c-gt9X-o"/{J/=d0%2#|4.mV4k|e<T0@v6Wg}25Ve~OVIRwp,^{f}o$"`oSkruY'<ON9(Zkd:5A
qdn:Y7:9')2}=;
UKOFb4x5OPG/0S"!URF[vO(=]eY6Q<xuu[<dzveV=./Zf=;i4k'Q(x27jhHLq<*e-5iRPy4x\1$rKXO^]Y^#-cLZU4"|"&E)TL,Mr@wHt"W#oc
r:o,852[Raw0<~7KWy5.MVBc2i0AN&-ao yP1nwM<49LbRD$mfucXV
|9kP5<I+`'sM#'mDY#tLI[!D!oqNWlNuTt,
[QgSa{6j?9ZQQb <Imz	*	xu9SjD2=#`t"z(W]!=b0&=}6tT)M=f+L1P^:=$gr3){7+~o
 90tmQN<wFTNKOh#6
t(qE#,E |)a>?0|Y93-#kO[WfS,7X2jxvk%$q	eAy ]6moI>)d>&xlGuvAbp6S5.c@#5\@4#V6iQ`6lWs|^D/Y<$kYcU}'Bt4YHj!Qmzg362Kz6X$B6m{m5}(?T<s\
l/fczT9Eh0v_gd\ 67Q,
R/1,gqPJ':Z6>@@OxL}6GN]|JM.?uJ:`A&zlR!/a'^/nXg	JgDSD_)#KeFA>l+'-4)>E{*>baH1KTg7	0'"Art-KNGD!#*;|h>~\5\.:{DOxjwQb3+ Z!^&SK4Y	6sU|b;w,?
K B	No7zU{p@eS%htwPz'eeq	): 0
Gc"^6UX^U7F*]d]	]!0o#{6Ta=AJXiQwan^@N{G"$@cSa->m3gD#Q}>%B4Z0luQg@ap?z`yB680sy)G,K*X~H4k6m1@)he{h4|~H|YNfri89Y=4<Ee\XZ-c/l`:iaPp>0i~(Q],@,\I<y\bPAj^Z	E7rp><1JJu|13KA3"XKHcp&)d`}6"`'?~=Z(m?^ND{&nmkR/$[X/k0=nj
`']qr;KkDHwb\\^P18Zoh!|ZC
g#3Xc*gjX+fGmikj(`|9CVqYJac[
TIJ~8s7uY}4D!j
V6W<o&|+8(X3'M}c.\V$"w^m&jUqJzKC#gJS8@`:|WP|c6h|;Glsii[?ThYs_[;=Woko=XcQ1a>O)W	8UA
]YF?39
VCL4Tpup!tFzN0h]!\nIptx`MI?&Gf<7L(mC(oU
g[.'%~NF[hhe$Ymf,)4zj^,Q0c}'N"C@	]GBz$vKA
f#pU3Zs u.}9Z84Py{?cf1>C&mR"F$:D=;@1?IIEPxf?C<OW-9~RW=t	U{ZM'T!,|X_.pJDyfY0S,/:8bQ.'njCdQs-Ja7
0ry4l]gpU^Qj)${[%xB6^pQZL>kZcn=m5_rRYkB,6w gsimdd|Sz)x?)z\-% wy|Itsx
Rir!'U!M;h>$;8]oq%#R$uE(lz+7
%Rq.Kz}t.3,QGI~
,8uukQr=ENn|WP1PU\h}=)-u4ke
KLXK2i'yHXA^=Bg^22+,=a.Q,g1NC,U8@l.'\qT%F(Z3+l&'r\	MS/:5\aloH.-@t@mcHXKMl.4j5!	n2q_~OTy[R]PxfLX;R!BDF%*>BL&:X&^^z#r9|a,#+Uk*23*-
F&>`d&)}N^_&VN0';&<^iFES)aXc)./<$%W61@c*QchhFh<bajWJZs\o=mfg&G0\ENE!h<At=#aga
+^lm,-XOjm7P;PvEvPzkqcFw>ra|wMJl^C>P@aJ@`}P$!oI(#6zdarhxB)7|WXX*<r$2{
|vSb4nG#-(6IO-Ep*#:T,2=iAj@2CB
4Yim9V:,\J-]gG3A;*:b7$?g>}(4#uQd#UcN[OwF^s*dK?qTMp\]i|:F".&*l&OW3$_RpqCxN ZUPa<s`ebC-IA6OF"~!'cYCqXx(49y0p#6cvV&k^|\
9<>Ga
8d^LRjgp0V#MGHOp3Hx^#Nb'.%
$JLyqsK
@[t20{eReHK+vU_0?:HI&iL3.P;tNVig[c:2""N(Y.wIKcbVKz\iAC-2^&J=*$B[2t8_H
x>C!5A(~d/;wc@@M*h=\j0{
pJ?u
1!?i2}dGPLU@mpEuCqBQyiIGuqYppz1KDR(V7YY+&z;MIq&CRx&G@,L}5<[h!sK:StalV}wyv?]d,k'\<m=xMyE|4*4J]fwru9#Uv4Y;*%1iL:eY[~-n^0#l;p@EBzX	,)\aM"~=:REM%'91SbphP[xpJ'fJ2uBM-uMtb=J9@CUD)%/W1$Cj?z>8%#;~ 46;2 c*jI-|a2CG6t~l9ju<kZ/zH}b9k[Msw!C^z	{<IvHI 88P\ ;:BL;,jpl@nQ|"EowrDnh9JCzr`zjm:ebUUB{h,eUXh"i|vooo(`s++4^pz7}vK	O3l}Ubfge	cwi$vB#{Et-FrZNe
KxQnF{ODH	we_+&}lZx(SJ6Z/f(!Xhv^R\{&x& agJ/fS.!_
_2bI$RyP GF?C-^ue?SJ+0[Ik5zw
%?6a )wg\N\YS/GMB59X+0%X0XY9){sr19F4sP)woE+hY5yvv\&W\hP8!<KIf(<"~7	8UuUX[ZSa9mz
hr2\$Y-j>ogR<rCdH(yM'#M1vRT)v7l;[8Xo76f8(
M(p[soSHiZ)Q[;aj\Bn%lo\kV/'`([,XJ{Dl2KA^d&av1l$oOJ:StL.vKKhGM|L<Myy{A3S	n"&H[j_ gOI"_ ?5#~y!&<&'\/A4kUwH]$giq&Y:H?	O|p\2"f\MYshO(U0&e
\nHz`6)8]OelgI5>K=Fq4t:uk)p
A+T,?IRr}Q!q7}F#S%1FPc/GeIVmdgl`L6;?&5tB$}=I("`gv1yd=hFj6M$^7uDu%Y
TD(n=S]7+'4	W;pf!X:Cy_6cZ;>COp5%miJn"6R*rrB+8; P4pgmekq>jg 2ttJ!1{xSS(	>L.Oo,si=%xY+K-t{b*D/o"hDTHWvX5)X7zyATG$y]z3odky t$]p{#Fs't!SLsG,Hw9H!IYlAa$tYMxesP!2IN3x#omcmg1\[~:u+C#h(3e}[mA	X i&L"GYQ}$7Q?cpZ3pHyR7dI)63RD!IV'E`IR=?-4XhiA(9{7PN0oBUwWzDitr9<@T%:xps	kHRF62Rq;d9&u\\3deO(6 }4q)=ASBu<`Pi+>.5489e8]&vm
pS	@"\GbK6x|`(`Ug2kE)(tge0CL2j>\/g0x.{voypi<lw1dy`&((BPE
7{\3&h2o]36U/WtclK4fyIBqDBIHxZdXO9+OnS.`*Xb=B2is&uW=G7ATMcYie0S}U"VD>y3\SgljxrA\Fa
5[THwP}D` f5Gc![;}]J{wfY!n8odq	RKhzC%#gWp!R.[	f'+dF7vd+-kYiqoUmei&7pa[X|'WO\Fmv0yiw)5xmj2Sd+#[hH['k@3)BK>
M
1x3z^- EOpwIIri9Hpxv*iQ9(8MYRS/"c_7)#8g!S2Nm}ZSm9%D$9lCbK.uz}cPa('RFw/>A=|lQzk*Wab+YLz/N|K{%X!OCu4/K*^jzv':i/l)i>MXeg56J^T&u13\lzDE5x3rm$.CRTD/~=+cxlZ)Jp;Y
mu^_*:H.l,iyz{b*)UZXF!'01.x9k0~[F-m7A0Tm,mC!LdCKM+ bW
gLOr_?|+|0mh'Z-)N4@E`:qj:\>y?rEQ* ?eHV
zx lPq`nHC#uI?>FP=W^=s#\fKrm$_DH p{!XFv>	P j]9HO^!MG+RCQx/Lqv+S4O<{-2b+d6YZ.g[P'8G4PXm@CV
L(njA9]3u!ljB}1fs.{A2c#Z FDIU{BZ)bXLOTj#WPY{vOUY,|.H:.%Gn
mWHV#(7Uu,\JYuk
9.|TnCn^vT2&z<<{\[B<i9dJ_YcSg<_jAkb,ouprZ_m/E]>Xt_eVeC/nu6mqX[jMT"mp_0E`ok;?*vFOZ;pc*9D@5AD^"JK3sC/Ejw-q_MZ_+F{uFD;DO6q7AnvippnT2
1LQFvsJ(Vrg
e
:<"_L(8TZp+Up\isuVfbOKJ\6fQ^9vd7fO[[Q,6".'&OO2`<6zAsfH#Aor.xQ=#|8
4B]A}Z"q/c{4Uyv.`#Ay{NNmNwb$WVZR\jRKr8C*b*9A1nvCq[v?W*ITJP	:'_X8B:.L.Q1<t(l1x2Z-,@NK.zD6~@vr9'@0/VJ3yNsMi{,&-4{TGoitHn	^`?<~UTR2G0,1FYZ2INKIn
YUI4jtV2n#sL]Mz2^b_A0aL3:wMHpysXuDkx8.QDYI6d^KvV5$1ZO-MjCp%Pgzj6^mgzIrQCbK^1XGT$<m,3fb<]e<G:M9rFqHWK0g
9p'iy	fqxulRe|8_e>bUht~yZGOi`,o!3gYQX/g rxB7g.t`UPEEI}VEFRtIXuu9{+`|WAD=t4yK}pN5b!wqF_&{7Vooq+TQqDd'2	ciH{.M[	6VAyp|XBs8Vbp`j/ zmPg+2o:W"r+=~{e&pKNfJ" tf"Xt-0KEdlbOI$YsK,S"W>S`],k
EE%:
`]0H`lUJ?4-;r@`ekMN0C<*.E~/,.V j%Ad.`l_1C?{qBF4 sy<L-zz-Q2IuUGgb	}pwKog'Km}saK|&0yLc5~h:Q8Af'X@;m6"YE2%/JC(Aj.9<CTERo.M	LDJWq2UD:3:.p'\>:lC.I
6=Nn_4l[ZQ5A*!uRh@)w,-IH{S6tdrnCxsY#Z
0qm_]r]Rd	iWBZOooe|Cj&[[LUobI/[u ZJQ8,?y-daroeR't'sr2y/SNT'
|vv'm6,oLvB}dI,0(WUW7vH~I*<hx^*`"ebxn,9PUEV4zCF{a?&s7'Iw<x8`dMy&<3TnH-$GO'|{$y|:]4^uP@B+7{.ZV|
"YlXR5}Q`nhDRw=VPn_=9(Ht.>oKI)}NN>>bOZcr.=;,l)}oT	D.o=b+h;Op{,+J}u/n	a=14o)vqkdA JHyvbHaXE}B!Gs-..k~u4vm-FE#[Qweq}6~$DeGazVH9`+OZuot3oi NN'Gl<N>~ ;t%b(Z}c=y'UtFAw_,cMBLy+^HkkMIbrj-=%wD3-]?EBR!Xux;v;c,s7B*x>@)0v4+k&-nN,8K^VEq*T9Ya~KV*nT|IGU`m	HX0e0[)1Z"bK`XYI^oFq+4T0@nDCplnR
QS*LS&(\\f]kg7PnL9f7!	ld:\OTHv,0T^C1!G10{>5asL$*5A4&BWciO	fL?; hmK~?'5SpmBF-bDO[;VYr	/7Z#@55ST-/k5gMo0GB*60bN]nuW9w:Ek-n#Vku:e*N?a m;^e5,}~XS=[g,Ln"c'B2#FC4#'!bHuxsOHd]	oNc`G O}NqT?Klo$yX_l8K"KSe'8!*9*K4I'tk=2"
%F)MXB,4.)S9X;{^T,ekvZ47ake=fP[#KZ]vB|xB`IvFxEXf:BqWXi5Q9b)3$vO?$1($j6
K?sNXu(t@~1q,(\U8R4*N_KD&`E`es(MK2~Qj?7iF
< moit43.)f6,*1?imb5bH f\O~V{:d=a/(Wg+2BZc0$e"}u0cB:i_~%__|1F8z|	u_Dm\XKG	T-(v/IYk[uv)kkB1r;_m]x =m##lrwPK+&?@63p|kH!qJlOB/G>/V@<]5mognhD9dZi!.oq9{ -wxP_Gcfpp3f]0IaM)B3SKRG*\WXd- |QErP%5N%AcOMzu]S>~,T1	Q Apv/e7>YA]Y4M=TP+Qj$:H0*VuSa'$y6 8sPxu/K,o% 1?0W p(j0y:;0z<p?Id  :\(J/N_FaZi=)K_pJ'lrEhfoFjGQC#tQ08E!|X	-F9y,R{Z\f/f+VKP)k?u_nHGOX+8gKkM'VYi|RrPFcdabF=nd^<h
%xiRytPU	<{ro${T0{dOtgSHWP15N7mbIH?5(>-^s}m.<g64LTa9'w@wAL-tczE~Pu|(|u3)>}aC4aH.^U#yuma}qJF@lInpSMB0hYD7w{LXhdK@Y5=]#KuM%\k6(`&|Y{5!{o<oBP)7Ber~pe*ll?4~sSg9vo&WMLgj0sgI8QMF{eDpJO8G	/o	/:R|lkCM{0,\?BC*SE'L'0~]xl^h>n"d!`nK j$]3

(P/N+wtz'An_+ ~{0?XlIaF]i?,9RfW8J{4UN~}Qh~z4~y
9x7mt^1By}7qvwV6Z-*nNxsYL9?pa\{8b'nJ8BCVDs/b{?{XkHed>|W}U]|21Kc^3^8]xbk~(ZhA%gTl|	rf^E>57`WwTg$aWtDBzyn.KM4l?(J0mN## U,fA{V;D! xXMPt(j) NQ|	g0q<F 

Uh1GbUF=!Ma1y)"A	zm",+agbtcKc3gMVlS{CpV")df/.z;j.L k1	P(=,-Bq]zuzSfbS-&u}x\*6!|u|p;"=.oi>e"m;MR`C-PV9Nw({|dMRGvj	Ri	n,cm)Ynt&_|FK.'K<qBxNq'CPr:<FlKntRVL#/zW#`r. L:"VB&4D?<4PWbrb|moe]uU)x\LQ1 r%M	>wdt!#E5C&:VC,xJ(v]t1MR<w]P5,1ed7F.Wy4Nn-N(@L9Lp`{fmD)+o\NlF;yy<x<@yl[EK<Th]*"ea'Xoyidx>RLiKSZANU,e?Dy&$0>[rjtssy;4~Q4|?RmjRK8$7Se5iZfB&2UC}Em^||AZqE}H$0|CMB1a3GWBrEVjKCt/<oW?x%jO1+KY?)Zv,L2VoM*& -'S^z4dh<JeOZS,s*++ 3 ufY. Cjf*VLJ;^q4qa"j4Oe
j?.:oQVa	"r>}/LTGrA pV>A5l"R/exZ_ji\7&U|x_;<9+QI*nT@YQA~({1I(*Xx^fTDRv9}ncb9371w/N-9<0h)[U$U){${v<S5st2yI#oJCiEJisjt3Eg'W'rWt/X_nSrXIU$kL?0A|^MgYyePq65gw!#^$'a
8XpPiF[1JTc5
`_vf_v/{`Bh f=shz#\2%J/7wlh,?0jIB1~P&.i|nM{S{C~*-])1W}l!IcrczPR\'"KY <BX'j{,9psvrXZQR(kn\Yq<`wFtjp%8:(5s 
!*(&^ KhWekxN!#G`@z	^trt![uv~@<l2"sUHri~~AT~<dgTtFy+E:knFNI>gA4W+&]EI,Jbx|
xRfAh56%+,*PrE}tCMeOAy['V+EoXU`JABf[=_.hn
6sE<QIp>fwo~(BVO*N1r+lI\wcvRL~cB\=;0](O25x (Q]MM_p8obs(kE}=ZZ%JdR,2Km8aB#T(\.Hw`
`{yZA9$wMh\4V.<E4NCMv5TX8l|'p:Kv9<p7-0c	YAr5'@k@QGy(_a&""_FR?B_*.3`U tO>g	[S6EU1>|]8?!l+V<A~0YJgY@-Vej5ycvVI
x @}~Bj~YR5;R$P.5vl1:6)JbNpMh8Q@#4.D2~FLV{8I:wN,Yg1E
lRKGE0|3#*PD&KH_3HR!=OnYCq\}+bqodD6eq

+p*&<o9xcL>a	FHq+Ofo+.=E0U$~BGj)=qOQZ<$+9XDJyRxlo^Zr;4lu*=
EizPE7u8ozlMx9[A70SxW;a49W$.	Fk))c!	 lg<1p0D*Iv$|:uK&:X~`n|yH,]:(hdH,(blhs.cv=4D{r6|uIwNyuyAqO5fD<Q*w1$!E>s@zQwbJc
TS<Fn-QrCwH)p%K*HWLktnJ.J`7'5fF;y^L#tytqp@8,SG'#P\zQ*W{PTu /%`.}AV_`5iggG?-@kaR &87NFF~]eP>'\5:lI_	lWQQ<g~xz%xqVYf5	O"VNUc,%
yBZ&.*N+x7t
z]b]"C{);W]t#U5&( ;wF=oDh1tA[r(w{.cCx6AxlEmj9`W#`1j)KU':xKfq{er2{ODhpboo\Yt$'lH$&5x~	s~&9'p +cffE.D/gz -ldN_Hu-KL|y@YD+:.zy}fq0*\`1l9>Y,U;`%8*g^=0F"!!</L9tA6uYLop@_57[sLK1O)|cIqZR4b]dK\)DFzMm)+h":a{Yvl_n=nWW.H{7!kkm3	ZZO%9Dq^sOFG"K/Di?}wc|gSv0y j8jRmJ^1t1{SyW,3`\Hvhqt?|5*L/)5;k
L 7BNQQT)O?YV4t9#;^dL$p{%6j9azk)"?u3u!uhZj;{7|dJ.m+;$qYxVJr&F?*0fRo_~{ITe/ywqaT_)^mPUjHbCx*zTty`}iR'YBf7w1T>UR<P<ptdSu`zTy]^88Yr r]z9F9Eow:SZ{'}8Sq&)jFHN2^(Ht]u~YlMEUy*9x>4~u9.[3,G^kL)hF*:-k
eiEFD0>Lli
Gn1*_3FF[vIw6b{9q"X)FaQR/Z5!vv) >M[}3;FG9yc_8WSDvT9GiVb_0eV9OEmOR3W/W=A1&Y(
E41MGDXjY/c:MP	]Y0{Smfz+{ROTs}#>eHf(>_B:
K~(+-<Q: lC[\lBz_hD~MC	7T:wIq2Q?>^}{UC5JD/?-3.@Un	_9Er'c5	{;p&NKvi!bZ.Er7<=.ZnN9`wu&}!k}2Up7]R#od0d|GXGm{[OT}YuaVCGe}B/K)C+hw\IP!SXFM-ZTX~H=s0`(7[[9x{|	U	JLjkF<76XQ;C6apxU6q(?f/fOLp?=*9CHL7}zO:Z.x3AQ)MmG`\e/mm],=1:Nj8Fi+wylv!iMTz\+j:KJTUcyu\{$[: XnA:txL_YuX"
t4}_&gzO!:}Z+	X/@2C^;y^rs8whLY Zv:!f	!s&#O}/tP_\Xn-I'C$<{pA[]M7"';FV%rk2*0$2@|"-,d"FwS,ibe/jSqaL8)gT=`;D09-LA>kv\YSQc$sU4@P/IBH:@7$9,6}LGKRH]mA"~<p,`u'DkMk0m6;pJeW+snK1BUT|E@~J6qF*GtbNH~v#6huqC`dKm)<3Hp~eRCCw-%3#gxxp%p]&NBR",F3P4S64Xi E'7n]*sBv:@SU6cmWY"j2s.3&b,kX,dd7Vb=S~DmtS]W9<SK<$8)*p{Q=+N|>CGx*:.1
8s[P/jEKF(./V483"@F<sq;nqe???H@opz\Ww,BY`p^K(AB)z!k/5,/JFP??-Ww8K|$L	)KLpH}dKe>A#;;4S0r*l%ccIxQgA!_o"t#OA5guBtQ04@>s;$(aQYw"Gj61'X-"is^Nlf
$~V(W,Z.6cab;_6U-*E'%By)tu_UU({k&Ij /7-:,DBti_r:h"XHaEabZ48Ah64Z?v!vM{BQ_vq8[oR	 \SKk;p#0oRC;Ezf#V/:Rj8=]MIBdO/}g(@,>4o|4]DlwUwNPgy'fa%CL[8vhya;R*hlV=8@~Ke'}EWE*r]QL&f3S&XDU{(8hMWDq+.mZ=Ph;'ZOEs5i'Qu,,8W^z0~8^Rg"@uW%j5Z5Mj-d1K4AjI*x9q9cCfcEP 0"9l	&*p^V(ewZC:20"UIBV6BLD6b	w1ql;lL#'HEm|('Yw/G(>_-vXh/@j_^JEdOPV}^<qyBS^M(|zPg5w$Ii,z6
<:
u+",X?je`MqF^fU%s};tlU@29\[jr)GiU"qmuvR/&pf252)T td!>-RCz!.I$27<:-B.RT"?	qxOL7$<!okU@[=%;_[Uw]IR:He[;"{eyd&ZmxL`z-:MA{k4oPm>-jUM'avQk+-gp-Ew#bv71D{'-qEI+mdAgzqn>84<JP\:#&9dJp@vnTI=S@{<c+XO6d|KwqPXKrMEd(S~JUtiVJ`;r
"tiy%U{VwN
L<wXga<i}%^aZ.%G3>Qyu4jyF&c*1e'Zp
AUM1iX|{YJ4/.Z}9x;dOtKq+VYCs#=NJ%TPlsFbg3HB#pzXj9<P)-*'9&jfy`7)t/w3|Tx`3)/ke!"wB)]Vum8tC.m)!(\1VWJ\'eGZAY'.`_3sWQQ Q47TN5^5&@nW_
LUAP2=+M4_.7-98WDb2lBhEKAQcj|FRht,Pw2.7a)T@4K%dgjUqjc)\zQFKNCv n^~S."5LqXMFuq5@noND?;|iXjXJ=.%hOe&f}ceCZx~^zU
H/!iw7TN)s9@e!gzOHd:'j rMp=.IQ~Jde*1|[)8l9+K.Ehsd.;4T1 6MM_1y%\*K{N./6qB<^Z^:hkpG[ogT- |3BgO]\g[hXAeA!K>1;Zi;C9\p/>yP| z}L~R\l!"Rk)l}ES#&"(
'ti'!d.h6h$%M)C,8MpivDJE"]XNX]6(42/v^DJm\R]Ly<;SFl#bn
>u`?/(8uJ["d9?J7(7RCq'oO5szK)$"?	\0"0i3t7>-c=hCi&!wS#W'&3+K$
M]jVfWx	7S<Ftfc["!b3B
'"ua]G$L(6q;`sNlt=?Ij:-]|XYBQ	CW$""^o0Y'ufdtL!DW~$#1I)Ee)ys?_, 6Z6~JFL:8zMlSu_+Vzk8YXzl-4gjnI25$9?e"yVIA"MJ6%.'v1K%MT&R|3-NO67H>
`Z..,}cO0Q 5"@$Ue(yVWLQEtzh2r7i4qQ<0Az1FU=-H"z!-r+}tZ+Rpml?WJ^CYH78?	;Yvd?al|}G)IqB;WpPf`>k:SE9d0&j4Q|ELN?[u]=Z=Q3\dl]wIjI?d%Nyy,<RS[v&MKjE"Opnc#5PA?T
SZJ{`)Z&4hwyLWWxS}TeM{-Wu?a--lVT7-^
XbeW	{ gl7$T[IZnH7tc}I@[?W?NL<;e%	-VT3QqNjJ0^/
TED:z\	q!NNH
'd)npxy{|32Ax"5bR(2;M7Ym17Wj76$F|U|pP[!b}@/5@SQ!z5mQA7:_xaPPi7+pMCb$Q	t<k_iU>>)(QAt,g<"L]^LUy~ljK7O1qNk4AZ|[1662fVT~)pRnjsD]X/iz!Z)/GGf5aQHw:>Bh.+B+rGqq;OtzBi|6iqfw\Du'l2>	BsMQ#)h-7Y{@"k~$'{+k:zl:SFfI,2icEPQ+2^Dit{2>E.B9@*,;+H_mzJN##-lA_i#a{<Om(#~EU.7HnEb/J{v(\ne\MoF%/Mv`B,ROjZd6&y)y_j)3xAxdUPRX" 
Kx&4iH.9~=Waa6evK2`G|i?&_n9D,NXu<Nr.{>.k.9-6q.;S 6yb~_dj_'iiH`.[jf*{?h,n1<m2xg^Vr6`QE	viJ:)q*Fk))~iK~G.{U%K>N),(YhzWq/\>Ce5LX'rNdp-	)50^(:R7~\-1!)fv%5=_@)v{*{,>vp^}Fjf8W'? E1Al6&YMj6i.TcDD/47Tp8ItA:TF3??I'[I4pRTBy9jK)ao..k?m89BBS
a6y%C[?O6+f_"a_Ne9L^IoUU"$_i@{}fdd,9Os0u8A#4haf32C)S;psuv$4J7*qMS+,VPB@6v#b+{Mc,.~uBqe<,*0T)0@g@I([gyo-m|KE#$I@qA#e1-VOh*T:m+?kFtfkS[65h7K/u:5&U*s5AY/,gUJ<^"d~W#y(YFsnDu4x]JV(z)\I,0fFZ}{on1\5_MAe4%o`1wtqIYrSXcu>@Qt2Z1Q3R*(+rPB?	('?SbDPt	YwDb|?(c[\y-D)B 3KE$)?u!BUX|/jt?)#6 x"JU b!b/Y^hwN`f?BfF!Ufgj&AmPckpj!HbW]g~fp0==k;?=<7Je.<N?}FEG/Cu9|[?0x$-GW_}$Z/T*oJiTx[:^Q'q<w!$/P91+UnG>7z$nqPhGQuC&^80E,1!r?AIaFp	iA?p(PVRXs}me\.c%|7pQHY3<1>q3tu;A3(Cn]0):C]U*=bT>AYFnI*z4"XL2DC0;63xjA2"OF*R}	p4Hg7+w{
`gc>-NTO+Ue}CJjlVT=hU`Y8&Fy#-$<ZJncY4Sy	7r
P|2,gKxA`<E6>a}vo|i,\uSNlm.o] BH7~GX%xMH )ngK!. [jU40v0hp	x1[fO,,,lUU'qW}.)BF6hXb4d=b/ta6V)8(&L-Bj#	vSS5p}+V(ntjZ-;{;ihU7QyR"ka'jm& `,$;}Ei<1:vrKyZ_:2<#VPSO`TPt2BaUx (@FcohtH[;e?cLM}#R/KW!C;k#d/Jn JK:0+/&#Rx#M.Op#XE'[Y<OeQ%|J?]ZAsi2$2>%.-o7imT`0$>J!U:,!-Kp3NY:/>zfWQzQK]]Hb8mm$d8&`Ib7aah(bI,>Hc5CtLdX`A2jR
I%
EW>+[CTr0=f@6^	sB}/<ze1%]}^9>DYSReTLzd-m+PWE>)cETk?
?$SM8@{ZN/W#oR\MA;Y~O#2k`j/I."y-XHG)^d|j`oD4hp<DQ V_%h'+er#@X06lB|\DXP}*QD-zNqumA=J.hBf6z^oU@)j()'|i?kV\-f'}w`,9DC<.,<36a=\		A$qK HE<F"[giAYv.)b	iF#Fc|/15<o<O-	xxguJU930LjMhCM.>Z84csiyuDc9u~:.x.`Z;:>
9jrqM+"K~(55"1CM|1m- 9bk|f7p:}Iw4'h\DyK:6=""?tN(`nco-P&{
<N@NfbCiWEEc@ *.NzalLRWB0H4crkY!g"Q]uZgVz+_Qn]k2,fc(nV-7]3lJE$#ay)rTd|A5m@s0
u]6\%?Y~:L!3\jg&hA=-@2Y?L4'^@u=wC/u;]0ZJ/69d.]($Y>%^h:(n\gk(8t7Ob8IdT-+RjDiYWBg},0`!(78|&1?iA?4SC4QI`:H7 Mb@e<j9_nT{9.RS}|C^}T<T4
}G781F)$2B ?`d3HunU
Jf|tDV~qkyb4eqr=-SF,.yA6A`cpCAwyp#8gN'Pc[:A`	r}X02{S@kxH0\seOVA1SQG#Y@>Am/HSH%1{"8`D%v|JD<t(6/#X&5^0"hsRD69}A$^Z$
kWap'@s@)cNX6~Y<GNgleFr94	6wf,?h(H3|I)uT8 [$=YR\!12dg<e4M<5Mx@n5us"`:>f<5^b=	+s	qV7c[{4A8>NZ7ix {"($~^&LW-tF1]&CyvZG=^EW4.N<RHYFY-+HEGG}'L:"k`
a)?%G!kwKaVP\+6Pbo1t@0`I*=$jd~mP;gleQ5k5bNQiOQ
}(9[]JL[6Amgs$O/ +V`<
ynWRh0yj3yXhdb
^P^g";UmKoGHg4CB9jx:Hk9)^)zg*\fc1Ke{S:opBB,';QH~-*/**'yTCJQ@d_]}+{	Dow-H[SMil\IX..9q)0uD";uf4 6Xz#o.zEsx:
]qEm`0rN|NNw056ryOESL	^<TZb\zUFQm%u*B&2@)C2i~}B6v}OWY^Y>V0o_VI
XpIQ"$VVg%OATmbl<wOD*?4p(smRu.YDg2SuXA=XeF<x
N`X@b5a
`_B9zl_?BP(UVW7"bs=tFriiw9=m\u'jsYcRPIsOkP\Zm9Hu	*t7ir^.[*{K}Kn?	}TDU|h
xV[	G4*zNLg34o\\5T^nc
&\i$Ab5o8@#oe/XI[LpRW7]_"I^>*t6):^;}JWi5W:xsP\vdMHzqs9O^}b*\Z;?o
B]1ow5_0uz]Jk}AeR<cH),do B Yaye6R,<PK?<FF@orojG7MFI@?-z|0<8U&lTZ&(tF?^t:d0]FkSiF0Unh5aUpNu-uK(EsBK}=iinPA>e"TQAt/rwK.=Sqe#o_-Lh$=)&BkNZq'>QS[/>YrODRyW,CNg!b|{FbTO,}V 7AJr=S>(O46;!k2w]U0j!a}eLF-;,Jv;O'Yk|vfY7"2YW+)WY>p)dP~',%v6Nh2aDzW9wrgX"y?,7Y][bDLhI:4yL>B13T"H8f;_G9n2U|]2zOZ[xpAH;gsZU73\_tAoXho6e0HHf'=WAWzX]b~NnlH*`.U?{hF57SLgN?|VV6xqFOjR}H^@~66nQ&IyvxVprtuy"qnWhRAv$,vq>M.W{^/bHx5LdWkWOt7y;oJKaDhbQ.>&3eyrH!!G<GfW {TP<gsgg!<<fQwk^:jU:RmY\.!&@/uaUQjN:ihDP:ywOG6hipD+J[h_X\p0JL]6 [}?n5im~<f.G[kjA31ClZ>0p;Jp<+JW<I2])yp=$){!p$lG|/04>&5aeIYzR;(f"o2xD`i?:E(.=WR[\;kS
>l3bRl	zvVv_OIpPYsw>_#<oH&;Tr"iv{]1&ma_w[3)[EA<"cJ]r'9+r"[1=<rS@qmim lyXL0P\Yp,R.Y>vD|B0tve*dD=SknKR4?6TuC8H'1r?H[alH9~&%J]9Q7L|z]t(yjlw_x-zE'6C}Aw6s$?'S,.Il6tIshA9b1FlKLm?-K$Ys:(fIt#Wl)lzmGKXn	`FG.XbUsv<rQhzqWTZ0udh;;X`>G^s1h)w/}eL`#[4M>ggw>m1"'WYrE|:)uTv&(-QioP$q:B=OV)UW/`->rV{Q? WWk	R2^5
PRwB-^YZ-}./p~9,&?HH:'40To( ZxU"gQh^#dgJb8L~ U|oYS<n|Tl;U%DxR?\l	7=jdv:@&s	JnX[ocQ%liMrL]j+VZtaY[a0VoQBlLOKmXr?3_~<t(p~d,\vYe`_XT#{%QcTAJ=o:u?0x2x\"yT$YfAVb$u?`mXp;-]g0|KDbg?2Is>F(@moOqqrJ0dchf
#-G,Gk\'=<+1(C2Q.XW=uAw)"Mfx.<y92k*Gl'|T,92]^%3j>Hzj9[aMuZl\.'2mE[~GpQ??7k)XJ*`SW
wwEei3jD@NR3v4 jd(CVt`0N3G)![TH+@"Je15__q@Bk:m`~.8y}impj7}TXDg*#L~ZZ;%}Yq};"lNyT0O:$&wQvsAbcpMd4T;u230TZ	Hb=-i" 1=L$6\Tb`+rmV5@S\,[4omDQMbU<U<z4,ZHn][pv?cz?Q'jzgb+"kM;w8v}#=ay-9+i$t<so$TR?_wM .M%(58v6pw&|+4`k5YD*DbiJ(zd9?+m=~$JU4<!c#]+#x$J0K2_Q\&5
iyPw@|x+A9h>7}p"c,BW$X4^:iT7<mvJstNm-~4'b4i,F!O	K0Dx/iCtB(V0:	c"i+th.bR&A'LF:oRL)b9uvAR{yi|86sHXuA{wQv*t)"5AA!7qa){y!HeTPQqCp*//L@M@57lif)CKm"yYS9w_'bB!8($XriJ|?~_V24-NbCbD#tU~7]&5]X2D@}8Yqod+pvC7	{k,eW$q-XX|q}e
@@}}#1dMbcC;w2j3+V>
BYRI!5M;r)~bD'bEN	kO	Q|GPiR{LdQ]J4Yf4DT^3cKE<^pqw47QoYDMcxNh#QCy,]VZsOg71Qa&Z--/ya,BWu3-"yjOx06nmufy)+&e=KYiat|!Y=P7su|+L1'=mnyM\qA~PjTIDP@.Q,A[y~U1DqZ!qHU:vV.a?=	;`})/36n?/0PK[Z~ok:"Kh"T$v,HXmoQ/S- q[w-Bk-{_=FM!qXSx<j?{_^7\]ubEmq4x
WL'>~(lM+0eo	W|w5'ON
yCwtD88BU65}G
%':2K3GH1Zl"aZ&$5lK`Q>-*;q#&y5Fy7}QAwVRNyYPB+Q=+Mu#lj<'35?<75~I-jr`36E3d9[JP)d0gHzK+^Ph/1K,<VX^Q8`%UMZR>b:
_ .HPsm)|V;4$}vWq>FsBT}-=H[' qMO@tecC`BAV7D"ulDQwQgF`0QDXD^
%TO2&[J]5(v(;*#3f K1Gt#QDs,VP:WDD7_hS-)6<,]G4y4w~B":Ge^D%'^si^]K<[6W.cFys`z:@<[7)J6L^HZ2p1Gt	%)y#d2Y0N}<~pO>QqM'3*6R^E?DP1uxM
+\f^UP^y^*dXr []d-R!Me,u{WJWb\MghHa(co8[FV "5[KATosuT7!+^.S2":d.:+.bxWpBaMORl6a_VgCX%>_`UuzX7C !3X@E.h"SlWr<u? X~d{avYq"^c<*[Nr7ij@2Y(?mFeVJ%A/9rAlh6?%^*M$?/JE	btbW
Ib=w	d}Y'Vw<MH6'?Pgy}j|!0TiLtz/9*y-X5KF?{r9^^/|ZJYN)5`v9UT;Jaajl[i/$W7}*:>5ZeDS.`5DI "^V@C"Ri'zY&"H7@#}.Dj)PP	C>eRG4~+}rR<p~lcBTQ;}r[
A,|*Y4[eiC%8j}dG9&`CM5;PfzG	&sm/t(;u9tBq1gB`Q<sz1pdd`VQ(Rx$LQ|l_BK7iA'bxPG)2`|:2WnfqPAx4wC~@&Jq W!uBQT fz5?O$*&k`*<(IMx~|PJtvb#=a@agwRb:I[pYJ+\B`x)p^j_,|X.zEB?hnft4f6|87l;y4n*weOeR`-/[X`WhO'|C*QO<!WMjc%k%%i-5m;	8\HL*<zzP%y[4,3cDTr[E~xM+H:4<v73We8KfwHUv;1u</[NR{p)UpM`Y'5kvq~n4?!9KqgLA0t\@5"rGh&A*JKe
efGX(Z_(:IC"c9w}U\A'; ]jJphhLM""":$lGKsrLsfJ
@u__ [ujea@3WR^awtB$PQS,rkqzdz0L]-abc
WOe`cXKQE4mv3>xJ<<a'CKxJ>[DU>CLj+w@|v5I&IVixin.H0XqhX3E=eYpVjes]*}xftr?K=dGY|fuVGc[6dw>)5r<OM	EVWJr	5a	r*+P`]eT	*i7J"E-biKg5pkWK0A`z<Z\+^MB\g89r.*]a4~i/$PNanbV^@iiV`&SWM:|@(@XhH9lH	fm,24m1r;WE$06z^GK;+/QewFPV{p G_
(&lLiE%nV6hi{w#NaLqyBB"c!0UaC26C-j=C9/68ws&D7cS"3\N!'>
7&z#"*1t;iJ] D'B?Q.zctpGn/qtlC7oaaO_Sa']FO{~S#Yk*._ub*WS,;11/\Zy:=v7Y*SC,Y	?t"QzD:_`=vw7SGm!.Z
2PO'B[i0;1/@=rf_n\]WPtoiN=?I,^?1clC:oE?&L,DPot zgpy
GN4xZ0i&2@u\h1c`/At2 WzMnX=5.0Y;mctS>hw[[/6EBxp6<lvG>#7S/)`J18#eEmcGVEh1OE9Vb*+MqLXF@C'(yCL9sh"3e[!1<^6IDz{&'2+	Nv{P_vY`/@U12$(OTy!5>99+|)@l|`iFGtk`H@ejHPN>&U9 ;b7J+gPn^nIRRq*@8nFl]
"%nh{1AwtvK2{4I46v7qH6Pcb*z"M0^q1#O`sOa
@V:f)'8[`R3	6v:Ea59v9e3qpmp#L$vT|?!e74O'W~'FHG%'jzDBYbJi)2o>a7U1EK$hM
OM@NYv
[IGP+e)imz1~.]~\xbX1mUUP-lJqk <%
VRqk%CCNC;Qr*jQcd vL'PX[NC,/^[y	`E
Teh*;'UB~#+^OjHv)EH&nApvp3&S3U=c	@rR!)Ik*`)J'r2"2|[7M8>B4K7KOE@iWGGfAuE0RloY&8N_W{8^QE_#dF4eQ}H`HA@U=ck*>&U]a>9TI\Ss"k o|dlX@#Q]MFs?v[xAIkO1X$NC.A6R6g(izO'!~!?d>qL<y{WFY$|db|J	'?]{+)pRwZZ!E4
	4eXTPq"*u_VAABUG?aD,IX&+228=//ptsS)'0ci`FgnBq<0$C9anL4a#O.
*/o5	LmoKsH?2:T1 PCQ#L6ZSDp-@Q(*JDUEhX9h8b(Xo/10*p|~GB/U7Bw5NLk>Q|`"h#OA9FW4Hd}")4Lr)L'fp{v=4v<c	+dL{$C2ATK@s5{]:\YY|TBWf`HL4"EWR0Y~2CI(lXb
+zV6hgwt`XX(v_o2
/aB(d*"6.N(>j`udRl0pm%`F^=~Pz	E!|@>GU)X@4vVy.O%`R,}
	K2Yt7p@-1~-4@77)*Y,]3)D#GN}	\!{|20)6z@=i,obW/#c?skldK{W=f..irdhNC'N@zzM&[#NVVW^
IYsN>#mTvN@)T>.9S[u8>	g-^>{h\*v|%#cq`#CQ^*
~szH{lw#|oh@T'%\Etg[[Uw^y)*l^3L`}an]Z>c4*fSN/S.g;>U=f$7Id(CB3I*T4yE"e&SkW65e84=S)a4QKG=(,]uJb4cyg$V\U2N%yb\IrWeD"zdg<g&x	bPA-afcZ<"qP}jfP,[ d/D)oDj4 w6^Q+uY
[XT^iLR^'jdy3.YFxK$la *@HP)*~%V|r\hY1&Pi[KgAF2'~)M7]1\X1$<N.AU.98$!ZoEh,Ai-r#ANK\!vj3vU?I~j4%s<J=tlO@seKDVe-4WQ{{%brKSBb83N^{0(^[?,jy_60Ler/Jqv;2h@4 }pX^-kt#wQ#*pmhnK	A^)-dA"3Y=f744eF2Mxe Cpn/y$"^O<4Z?"Oh(mt1)yHO69A5> p;_/vx	bWO;Z0@z,L5F]^)NThIBStICjjtjNJx^,ah9:v2xFZ$wN7*yf@j;7	\FrE)\?
SETM\/CMZ5-8N_TeN(QBx[e=wr5P,9t?U.
fr<+^i7?GS%`	@DC2G"M75^U8)Qc'qsoDFK2J)U(S9vf|*7](k<?m?rg|-.WDL1Bh JT>Its'r0B97{{]Z7w-r0pF=0B9	Zr]qhZ&-n(z8akl<M&]/2V0(<L3o94Ot9JM"tnR)"L;U#\S)
G^@ObCfnyDu9yKEx^GP123|"	b,F Iu_1CnQ7rCDj=vnydRl<<&(?KyNKi
a$AITd0gxR84sGDfElv, G$:weml-OOjnPhuym7-usBu(t5~xkRg/bo"iEEQ5`yZ]1a(32<SnQ{lm$ks<xz%3[czrBI5ULP]NGF|xJC.Xk:M/hE$+Uy::i5E^0Ap^?diHEZ?
e7
GJknAPg:$dq3bK#2
0#x wDYjQ"d/ncp^tAfv6[F9xh?`eQ,:hlh$pK
"@""aRhp05?GtCR^:'BJP;CYX4QjtOeO$vMI^GefyZ$@(Q[	5ee#^N^uIV071D`Q(2pR#ZJ_Sukbf!Fy2^BtbP7;`U':4d$[`GIuQ?z%FE:iX4>.tUX.LkmaF}A9^Kcrje[WRCbiJVrp.&f >M_69O.wIFO~C*wE;5u~R3\3wWf=TQ-.Q7ow}0EYi;TH.=R	5Cru}A!UE1f;=&*w#FuOqP)>O-eyN^m2=[?]'w)$(qOHu0U?HQ])p|H&[k5F/&} )9|,sp<8f+5"|_I%'E\DJYE5Qo3,lY;U-.<vgXVGcy^zj3R,)>>"#Kf<dN=O\g!44APVKH'Mx}
2V=SPAV,yjR`2=OD* +Vh!>d$nZnQ>bG;%Y1_Jp%TWmLW3(17?eC0AIpBkE?^,?
zk,s;j?}9"D6d0F4bdA#Lxk5:Zxn!fgh,l[CS}X~lK/M-S^q_L{~q@QJD<(~s/`T^>]Y1SX=fH#D_)K
73}dx{a\1~?05M|%0s2su;fa;2w6JlqU4O<m:*_jtsrL6%&?l
]vDA=4`Y`AX\0g Q&:&bZ [W on&w7_ A!f*AYC8]
wiR Q	Fyg$y3`<|g	sjk[_.~{O'@jIS_B6_g1+d#.?N,+">D] CEIV^%TG{XEhh.l@Z3|9%Q?]D^.KBPI*Qz|"% DH~n`5zC<Y<T(d35yGmc]OS}js78[$6k3K^
.e>Gh:WPl)^L!Z??6};tQW4j@X| Cio{{PN<_
f]6rRue{H(9`398*U84c]BByPwC1MoZhx^/h|[\Z	kokn?iP%rz"FBUChI+_|)U0E?^\!I{[iL=';tU<hf(0RNtg;PiGuE5$E\Z,M9Dxx?}c^A"4,>z2.Eel	)w&%!F)"|	eZ_siOyqjAWl/;,1~t|7S.*:Qd{lMg5y#[I8bcFY[a4!O~'D|96K
9 [X.;}	bYBk-rWa<	1aIWP+~Md|/Q,DK5dO50.Q!_fN'lnLf&LWSQvxV 9o!e(ELKz+Par8ZN .[N5$)$q0E5E/[;SUAK\hU]A@A>vYB1,YihIuALQ&Z"9 qB"9 3:K'S<)4$D%TXX)O4X)oPQ1!wj[",HCu8d~3lmtK!fA(#1~Q^^@]+ab,lv~bx	wMg&fjT/E=xys
2LUJ`{TOq;x,~vWG^\u96]]~eJuT'%)DW)=6T	tDzTKB7_dnc(jmqs$JRMv,PH	jhL,a:6Y#H
<rG1}8]].bFo}*@z3v8ie**rMyqvG3MMpx
Vo<l[%Yr1-k2w/IAvn+-iQHXXj|2s_Cj`gJ!HtlE_F==)cJ&2{Nq[M(ce.etL+9VTHkGZS:snH?0T[%5-z]0%t1>A)jG3K7$/lZ18{Sl",NejuND bhzt_U
>:85Mh@^<o7nm36:zO(%asL7d4({-bZcdsG<Xa/tmQsU',wheLdg0gQzYIX:/\EghX5sWvy&GG%:B`x2Djg^sCt?e |.,YvpV6Qs1pj|"3XHR"RLD^0xg/Am.m4fB`0X5B91j\q)Z?M4eRbk&V*6E%N6q,bMBtZ=N?mV}#";8VhiJ,94yi}aTulNnUs4a++"&/d0f?M~-=gOZg_~P/g/e<bkwUVF4G45{crh<dR,nK+6dK
p(F,7<su5 I7VtCtvh}dltgMMj@~MhBH=6uI5"1ys+_wf) S
X3;e AFx\b*M?qeXFB["i9+CR58k)"D vGl
9p||z3wk?@,K<E5Jf(iZ#\::z,BQ4iz$ga~p.WaMUd}+G~Glrl_ A\Lqb.O@C0OCauVN,YnO\m;m^9ko3)=BJ-=7+6Z43U0|
IqRhFX
:4QJ
5oIfEo8}2Bj3=lku)L9~OjFt#X'.N"mAF3T]m1UqL@yQ2[*out*V*[~l8x`y;4
p.'w$xML>>KFpI~("N&WUZ#n7"`'Ey[#OQwMLM0!"A@9N`
YfOVznd3#lU2Ah`,p;oddvI+n,VW!m.]Ke0&b[(%V.	_g4}*Kv0Hc!%nB39wMJ&n84@zDDr@|y@g-\0`P1-
JW,vS$h9_Z(X'P(e$_3_C8`r"5;_p[?VlJf#8%jI1O!I1i,@zV3UG0;4"@<&hbM%]3rhB,x3$X7&83l1{%!(}@{I4&IspaFDKS@k&Nr.ysr>_8D9W,<oyX5~;&1"PYzeXG@ln?]?Kqx)d,eT{Wju[T,C=w'9RvQPsvW#-U5.I</4BGx}x,:#e[#v
%&$"'Dk6`|nIkoq7Rm^9B]Vzi1}Y	*f98E
$qvO|`8"\j+1X^^m:R)*mK&{C(Ho:CYxG% 2NZDIRyKcxCw\R H3B[n.fAtg	8
1-7"9|Jlzi^+SFb3o?jL[OCfB.1ymk>RnV2m'v6%(Zh7Q%Qun5$aT8n l`ZoEOcof&|@r.c6_b1i~@23S_=iYB,6s,,=g8Yo	]8XWyO9WX-{v<E>5C=Z=)WL!2&x]^	v`FuBbiRNG$+mXb<g"<2TN:IcE"U*)}p>plTt1s^p_DcQq;vlBB/#x#0$+~+f_'k{i*/YJ#o
oQ3:cQn*m!_"({(+65{,07+i^(/JH~5/T.Ah (\E|5(@?Ey]9KH"?'N@xiLBvU*|$>vp}`dzG8Q	I;xvB)tj)AF:&s135Lw\30rT<[LIJ	lMy7kvI? 
[sOM-&ZlJ K6^(oLqjfd2-/)lUK%OC7/C_4S5LGnfP+QX('=5`,%k~#e'lLLR"\4A\j7Wh]=UmSUMRk9#\	J3j=j!4bP|Jy/n-MMJ.x6E1ZNEvkR=944LgpHW
'RQC}zi`URDal38cBk)QiVEY~V:F5Qz1",-[lpnE.<	mQBO2P^AzGE r:]"XM*s6B?i.-wxFWXG-oEXGNh6e$vQV	2LS%j	$b:8\	rAq{cyXN/KM1|j
B (Y%;9U45\#&:#`n@*haZ'RV|t{]RmXGEvA*ON*)&	1jrc>#QUb^`{No~(>G?VgIqu/g&{W2gy*kcDTu#0t!n`b`4LP/jRKp(Ey1IJ]Y]AfoUf3$rsm%YKU8Dd8rMwp59MEmCWt$7pX+Y\C#$!''N;v%OHk%0a .eu0Lt'#;Ufc\s6{p+js/@)nz?'BpY>Ug:pbv^ O1)GuMHtwFx15z-D	ENI$
lbd[iy(\Kkz*:Q'C
d"e(+>Y=&'PD]|_]=Ms=F9r|L(}ay[
a=k$n8t_`X*2\~[J:|(6,l7J;s hu5ybdw/O0x8:7^"{v$=Zts+0y]eBgz*+r:QdNaenLe)u2Lk1n2AgPfcq_?7>kq]B3JT^Z
Ujm b6L:3MxST,I	yu@aUKhY4-H-y3~HsG,:v@O{Mn%X~Fikh6*>6Jp%P~MXIj`6#.&GxGe}FFoZ09.<G&9<TZmVMB^y"+&uUYA&>FB[LQLmb'kh,yT;Q!xLGLl0heg\QwtY W|<aZ;7edK L!0D/q(jHfsCbCG;ocw\ec74P~@<o"McZYt$ "<~-!l0{(tj^0MQ;+oy{>%}2g|3]pJ;yb_"3
E8	?ZgRUnp=]PmH,[:)sS\q.{WlSQ~2=MD\FBdk\e7}| advx(~dxfyE=sZcjg/WLp(]5|{dEb{IrbC	h\8a:CirE6'-i<!N36xdi)`TIxCk+pr6N(2Y9$]P8'k0Gk hBg'BPb#zy3Zd4v?LXV	8-qxa0?D]CH\uDven7_;z-{TUx(A,	f>uA:HG|z_xj"`O)enRz_P
@u!CyT1syzIR'QUx%n!ew2o|}'?;8d4'Acq<E
B(wUCG	:+5Y4[uP_&,[og[1Y;(OOV=J+9AuX`;.Ja@</[=Ob5um$1_ms-d>@vhm#*A[vA}JExKZq
sHM)bx6$#sRq6ypjm5D	7ET> MQ3L&J.@!NW7FIeFPh[r?iV$$G}[#_:)o3^ft%`
}GNwPJ</:fSy:5:F6h(eMUB-CXRF-26s8W9(mWDl}7+?%&	Q;7e6|MgFyvA"EGgz)Vm+E$]&f{prP\92bsF^NIczD}K+#I	;yZrB_g$4-vkVy7 "~"Bd+sW~sf_dsRD\gu$
K!0Fu\_j\mw1!*y$L .y)76#+26	IZOT>1U|<Y?C(6a*4sDpsV;Pq|ebp;sIW;]Zu]z!(NX,G-ItnB@/2'(*MMN"ZrmJhs)pOZ^#w.Ew/8;x5luSA$*Z$x2_%{M53|fW,/g\d> v<c)IS1VJok2e%$x*n{WSnnysN!Hn~-{,{
x)N~K@k:O'r92~h_:0v'x(4l'"ReBM,pN3]](kp?E&hA.L\J2)*oi+eo@~0`k	H
SI"[2(%rh'ol73cq
(#@Pal0?xDJ %.su3|*)\%2A:?2'(W[wCr?
n}A1bcG^^r5Sz=.Fz4g28+in.eQi
^nnXE\}H>pk)JR7{tO%J>ugK,U')stts')o%fvL4
w|dJh6eTfvh|`e]r&0%DXr9^,f^4'A`b%ecHE)$
s:2OGZG#[`?#'v0LR%#Hz`t'\8{n- LQ;3*_<4
9/O1^3vnKz u=87M|K:H=}f<Z8-LSiz=o)Xj:Wh]RWyLd4jiHJl/^F<&+|A]Y@f`?c'|vZy(oocl@8W|:1;f- tdn`d,E]J/W{G}T]<k)tPxeR=@(b'EqvJMNi0cPe\Kz02pv}6|1!
ja]hpl>ut4g:'*ErN%Eb55m|04~PqZskm^pDW<O&JA[4;d;qH-'C(~7:F^I_B0J;`@'I`"?<O3dJGlJe!7$u"zypA2}9i!|\lb}N\^lxsb])KwV}F?9;<qGPH}jgmY*lcf
n6?_Ti#P_"?r!JX!fmyzdkA|D,1iPWUdQ<f4Sr<gqR>)48mz:e#\7vy=Jj]eOXY& iDG[.91ak`:EuZ,YHB@V|+z2QJ<8*
th#N5'1SJ}A`#QcsjDE~dt*&JcWQCx0"xhF<
`|J2'w
nWdsZE3M?mz#8O#g!dF#XYu~s[f<*[nO	`h;nNuyt]KjrA-F/!IOh)
4jO7^>;K9)Ak
\yfqJyUZtaA$n]VL*w6A[BVxuV^lhe$a5=r``	96h+~Z<\Z60|e3SYgQiI_y
kd`t=%suV~rd$#I%qBZ5&MmQ*e"Ew)hC8e*!SJBH@89 
!k)`*]Xwu$/e1hX4[0ciV9xkgv1+u6P$9imsd	u	r(]qe]
}LY}qDQ nNPSWg{yVk?1?/zj?]p	JI.^eT8@KS)Ow&GNQ"+@JA
|~j&`\mGrrU9]0
;[vv8g(KE-_DL[NVxM)CHxmu0sU8qu}>#Y;q
z49(
{^P]U+E>6v9&W{k?W:]qb=
!6NoEE!qp^.Qn+f:P+o%_`x#al"24sI*J"I&F![-R2)fK\;Qan>3Hjh|VXQeC(8DV08y8{d ,faD-] x#CU.eFzS.Mdya^mpDruxS7]U93pR24Cy?LoSiE_58p'	H1=@ek6Uqbl}QY[u%g9d,-+}`7=EbEp/`U-(<*YP1^6}SUGz}]ekB%~CBg,+{4=hT[Wt?!mnj$>FS9J?yTv9y9D{k)L*#edf3p`G9p'`ztJ,?r,ctwLh09]aJ!xn^!]2reawd{p\rL*pRdc,=E&2r@(
_PmmNt:D.7}<eq40k(.gy=1Kyt8yFg!PxS/f!C]#fP[-t4~4mNRnj;^\+[KVFr,jz*'8(IdOS|ZDt3*B>;b/'Z~R;ItQ#ukgB\o(ZjVnPR"2<$c{-b)#g71(L38<hibJQ$RT<#pukdY7jFaI{*6>`PD:YD:)H*vyd\BGDRIy[Y @
uy^3?oo-> LHP+!-+5$3	-Q0	'@}z5:aD[N@x|@WYl9$dMr>Np<i{[gFh\Zi3YDcrT.{eH&B (ZDeB#xiY*pTWoa5.WKk/W@"
xO+erks&U5WwIWe0dZR'A|od PbC6wPIQ1clDBm^hU<c-A"-}#Lm-N\pk&[bl3e4s\(,<-*3OE/z8tm54z}0R:P:g@Xs]5b_$fa}[L"qdC,4BN	#jOd
MUcf'vv"A1\\vIga	Tdm1lXG^4)pxr\/() Xmb\(_}.x`;MrC*IKr`ELKK=#f3E\zy6s(!lBh3m3C`K*iT)\vFiA*sL[d
_IN$IxCt_=BR^Gkj`f\yhm>Gon!/Wo<VXCb}46gk?QE{yCDcS1-\JUFq"detL&<p)fALFxdg9em06bk	jmP*7b-ndumi+z;@F.Uw?:}H%>K56#=c/g'f,-2#`{9[vi}T`5#s{FFEG%gGR%^r+";8'm37R	%x=#'>`'xea ?J`aNDolhQ ,T&'WyA?}	m9H{06st1M`q@u )y)TOhisqEu>$2i9q{tww}BFkG= 6_dLx f
"C2G n#>l)i$>F[@),{0B_2TYXm:[EaS :CpY!k0HOzo@"k'LNue2Pb]
Tj{_V.l(-1h~=rW^9Cgl+in&CNNkKP(-7-_CIYb<pB,1"?Nl3@}WPbD"Jp9E?b/x 3O$(sd0[BLS,g{ 7aH0i*^5lMU%f93!QM~)6cx|eQttCqt(kZ+xZZv#D"\E,"!I'X~hW-
7E^uz.Te(#+):tU	hM"M7[KAM(yPdGJ7L,0DXaW]g([8x4:kHbmDJTxHtd<wU-BCwr+=Xa+d=~Ks	)F3e~q.W;t4|A'Q*"1C6rGa4g5<UOW%,Cs1EvW.^S4Dvg|p.lsKyNYC0p9jY]4L8h%bu8kld#e@b	TQ/`t<&]eteB	'RIEw2I,3Mh,lqEjKq$ulZB+dOoq5r<E\
N>k}+c>(G_{I{bn 1,[59-YWQp]:gl&&Lk
c6nw {lWJjTBs)C~w-d{f%LS&mvB2*4y\#-_dM$>kTeWS<s1EXZ*o<t{$Ia38}O:XLA5mqz+3o(pQze+(4\w'(<2V_08/TBl/fGD->
i?N*]Xz#V>y>UQPs?uigZFT7${+oZ{NaEYK4{P)<V k3'6bGLWJVnw8w_\svEtC=#S&%q&
IU#e]I&$
l1zIZ\fv.cQ3R9/: zE[g_5kqa"6k[)V_M`& Gveh@-.}VxV'N9UCY\2H3U/5Ei].o3CYl?Oiz\iST<Yu!`U5\^ssv(yz l;8{JGc(}-G{v/*hV0|%YBCmvy`v?=1b&Ml<D%wD2!9UOJxAEG#'CSUC~aHl$/1{w$
e7js\1'Q2CfG_CZ}.;7AhwSB	qg5>@Ge Di,zQu2swx3F;o}$Cn,FGjifNT<;Z556FP=iX!Sy<k*as(-u@yNU;C!$a-N.+\Xbr!ViZXxg%o|}*X7,c{e!6vpd*$L	~%VW`'m4<;7b^(+=qg4lJ*[Ssch,][a5g/A~!)O%8U={V5JB9:16c{GDpz->9x- ~qEl8}SDKba	S__hZI8ImvBEL!RO6u`drJaZ8f'tu+jU"!m'UX>3kT<^`cs"}-Q>#OOuGg0XaLq[|Dl-i	M9nwlt\Z#G]8'Dd%x[9;Fw}$M:Zr"~$WVO&S.I`pnIGY/MYE2Nlkr%C#s
o[36x	$giK4@}DP+|d\P#b'
7"7*Nm}=tk=F3!kbS&7y;Ua:$@kPJ(Tp{PUjR;blOVYF^']DVY8$683wH*vG9dJVCe$Ix-&3@G/+4@FKUm8=h"[Qw
/,O&^c3;-a\v91}\F4GX+;8RmLZQ;$,iJ0!NvB5d>(Wo#-{v@+dS~"7E%K0Vhbd=g^<w3tF5U#L}<gxBR}
V(i1Om)v\hb?5.UJI;9SkwuS)=\:`[3(PrnYreX`tv_Pku~TS<1U?:p,cLx%aZ@!}odV (5|6Zs@7}|}NZZNeC: S7MdA>q5.f(b%W/.6Vu ('XRbwn!/O
kpPCz[ccBF]j;F, 1Fbd^M@gcj+?/kPEmHmcSoSS<e#|bvx:$yon c~oX)[hz?7A&3wA`|*JTsa{R_'OX47S'#h@<MJ-rsaXI-<#56n+gh#&qLK3g
vbn*Dh%]>m-V0=3#xf@k^/6!rz)Tg6tT=MlPeWJ0x6;m[??a=?!Um!5y0:u-`3`$Oc:$d[@QO:i*$(|.fiPAS<e-l?+S<aUc}f?B++	rP28CJF71SR4mHU2kx^`Eh*lf@>Co--W&oWhE?8gaiRV\E~'6]H0#GIC"ogJyJ.kiu3-1PH7MO4loVO1|Q"&*sWD)U9"n&8CviBsf$%cu{kZQ+<qK[-Bc[N/hB`&pHFKZ<5FKbv~/2W4|9/G:AO85Y>}^
zBQ&o`5tHHgU\vu4W[[%k2p}w~o[0G9qmaE%Q#TfX+\;~~kl5>v'jU]JBb=+"b)J*lU</v6*0v`9$Qzr*3I+nZ[\`2jnILZG:S)?cIU-],<K:l'GA'.W
VJnM6V_)\uJiFXtI(*4^S|ThcsuHB/[aygNx}`oo%o_4l5@#Unuo2gsH"[}e>5X
c"IK$7h?_D62VZEgtIO0VU&g]!mHp>J{<FvT	}45e.%To3[flw	Pi4XV3zap3/MmpcoW3%KR&^>>o1x>u:=+O}ySdD=[oN}CYmB(IVz9X&Z_bV61'ww(?{\Vs'^z:-5M	}':_5ZcrM#07F}J_g*n29@n)8`
 )A1-=ckBVc@5co#U=fx99ZZIpss{JBS)|S/?KAzgWWD1Sdwg[izcY.?V]6N1*}3kKVwJ?g_p'WF'~'u!,QKh>lQ^x]Ds]/lhDJpAOPM	jz%&zW)i]~iO\Z|F/Q2x9M23H+js	SY`xzHRm!5fy&%?%3dLEP$#Ntp=&N;oag2>&*~+D(I#*l&$$:+i@0pyII!t[27 DVb.<t;GyJ]hbB~t2roW{.x3(,!A`i>B">$(!O_;`5P{
(HTH!pr*UC2cf7v6BXGSaoYsn>I,<5*b!
\%`S%6|v
4khe)_Vw<<@il+TcMPSvzKZ^$?(KnF][W(&-+,umoeKKN@;}-()vN
|$4wB:Igo/O/`7i4B(z5M;V`aO}0|@	w1nR$45jJ
XpDoOXr0h8j[)/hmlQ(T/W216WI25:D66p!@oN
`	FD)c@^5Y5mgTZU+,{ [wEa/AfW-I,}P~V[,%P0d
4fwg|F0j
3KnB1cZW&0)'?"xqij[_ u"To/6}f{b=3ja]8(3gWo<IruN"9jMr}-'w,8YqvU5-,(*DKa% zC(Fk(`*f6v
Wp}0YA#1e>iYd<U0vk	vxIHwV.7-Q}\q.I=M@U[.P}]\QX^el[!H$4NXYGKxHSpu
"bt=0YM;WbJR=i3#Ps-O<Nw	E\y8_l	RP^@x!_gspGgnJ&{%XQdhmVjP]jpuS8~SK5GX0"`r/55g@HxLeN+L*AzvZ/iC*R{/=>1@1.fVo%cqpo7]
]Z9_R6F*u
mMXDM~E{eIbJHasA}2VN oKmK</6"veNXBka+ngX>M:Z{X
-+Nx%~yYzn#5@~%U>*BxJOv7m$Z'BG`Htai|RnBlM$k8xyw!+~,yB["OG[#P?@@+j (o
jb=V4>~%GVx;KQF_Nu	q,(D;kFv$~TRaKUQCcGLq&to>.C
s{XH/`t\\HAW'?m}gti@vI1]L4|ylq{=:9~] 9|w0\bMYrZeR$'d2J_rUUrlCYy	KE)+wD34h3}FT7%d*J5.	+z[du?amtY+LM&k1\7hMOwA?Gj!bDlT47o|_QlQE*$dQGa4Zy+z,5@M"pu@tq_CRyU+Px1h,sVP?Rp'rqJFTdL{D,aC7CvpRqp['76Fc}B61o	1I86)(bdk?D_#X{,K7Eh
]S,'4CJQE=	Ea ]-=eoq`uT=I=6x)JV$\>y|Pf!xzh>Rj.n=zesA/X$sFdRI"$#^@rShBQE9'Q|cw.Cu@~4_zT;%-yL{uFyDoN582&T8AXPm'	j,`)@!W{	R>wAw~c3ac(vFv;Z[B"MYMaBMv-Zk*`jRpRn=.aC|^NoLaRFV5S4-\0.gQ#sFe'Pxn_ba{x/g8FTiK]pf0Rm#X#/V?bl:E)H7;)<wk0`{0xP,=CYn@1'DFE+|8J!Ws!00i@q,q|[A	TYs`
Y%]]F",E-Pv<Xpx`Hy<G?w_nK-.g \)/O;LUlY"s=vM(mk	QeR{Y
55tvsa*ueVr-NPS)4ll|2(H !6v:GdpW;A%F-?/pX>@(GB)j	9Vk_D@}`c$.!/M/L!bVF	*GT6xRe0'R{Sq9[f1Y
&1m[+Qo'Yk4&
m	1Ha&&dXHCRV76y*4jte>w_C+H#SyG]\D~qbgxtE:X(/77_xtTh'f<Gu.k\|:k]I}f[u4{c5Hk^t3km+:Jm?;l#T?esedDM<P/'pujkvwO3douFsn32
#[{6)"X@4"hBszYvYH3/>r@3>BSkpx8'@V1%x-#X/TD]EH~M1aSkEJc1(w5%I#};r[0p.iZH"4mEh<vsU[uDVtE%;g}mtUW0Ot;*<bc~0&-{TjKg%ot3xJ1&B]|K0J"}I8Z64fvytEiGE?`Iu2(S,3r<U\d|2jt$?*>#@r	L@9|uk`$=g<nufG*?"<'HENp~rP- 8_y|a+%Nk&TqB n1_~bnDIcVuX,$!iP9Cfw,sc"3<(x/~WnA@W*F_6~osjD[BoqBhS7VGhku^{$6X|sX,w$R{k!UkvT4ZVTT{1KV$ova/?vT]AX=W>,GQVXp}0DNT;lohr=1Pi?/@l>KD3iRyVDMu;d*ldoJ~88-I`+<y_K/
Wc,xy8hbChN0gVU#(HOP..8	o[l4yeUcI=#$Z Q1~jbys*]x-/wAW\UO`jX][+n?]	9bb&dYiW%AXq*>:X!tEr#'1V"t{+w*ILG$?<B;w	Cs)o$Bp&8>KFs;G=cU_Df=PA<=!Y.`#W$:4]ect^3Cs@FG!RO'd<#-wb
k=uU::XS2&U3nr#z$O0nhkGsR{,pc7|^rD=oEEyoj0,'-v7FNz
5Nl3M@i7-JV?0p^DY{l``1=qDN=Z2<<,Nuja-M!>	K:s].mFWc</ZPf@f|-?`S7?Dfq\SWio6GGn-<#`R._z_0[R$GoVGwRV|=YWB1mo^gx-soOwPA=nf]JkYSV]Ni>}ZXPw@5gQ>"*0%ro' sSi*t[K>%'Oi-tGH3@IYz]^za@I5<v1;#bx'kyb)l23=.xpVVlqCXq?O)V(-"xlFkZ,pPolLm{P/)m/vl>%IhU3k6}.Itku-_f4=g
Kb`^^DW'4CcpIg}SWQj<Yn/h@!{T#k5p93\mYiX)S6I
-6;;dZ.LVKK?;yX[LB$oK$5
QICboKcl/pc{YWohIOh-RR\X|,o5,sl'T_R;]CVcdVRvtbZFu())s8	j6:K/e&2m@{p)&bl,^m EExQM+`LF2ZTotjd$TN%oee}{NvwsCx2fZeF o.2;WRD,mbDM:R~=Z0,H[W(dRxV]#h%|{FgH;'tg?ad,w04Nf};lro7qa:ap~LX<3hNU!>ZIP+:iqF[AL2r?B&WRa7s{E,v+?T^s2H`N [5~_7@SK$4:Ci\cW}jMOnehwdPT7pS&UX"*gq'v	K*
k^vPpJR0OauB#8h92b$y!a1VeZ%fG03#ZD!G|%`z}1vDek h9P3rBV"V,wndpn$2dazqr-~H4Xw/{sUY7)NtA:?UV=\]I@W'9]w#6U,4|SQx>e@3|}&2HW	':c%-d,rnu~6=cP^T\6<<v$>PFC&(Up3pUF[*6OeT`+k{EkH6c	%U[+%{ND@p@T/F)cCmgsx:z
7&%Y
|GtQF2k<?2C>s*hV5:qf,ILS>*'h1#/.H>pawD/M,@cs)`y(%(PS5KpEmH=Uf@PE(/)6knoO-c2^`e7)`#)uUY!t53
MkhGyQgGyK(!%-IS&SFL$Q"&6MYBx[SGNk0=RtOh@/!,E?|D1j<HxFa`0w;i%Gj&(|_+/Q2Y'a*4)}kG5$=r=O0?&`iuR4u@XLfUrabxYPs.\Vq0-.C-AvL%)'MHg"5sd;\gtTY4#QEWQ>5I$	yz)@tCxu\s8}Ev'^2.(EBI<v%\b8|4u2	[7:.?k79L=y.:*k^@]x@\U4nl[?LJrt{v	Ouepmw%2,}cJ;f@7dI!eyp"z5?ut6{h>V2vWQfl
Ud<7LK:J2(&1(Xzii2=|E!|&Rt
F#;E3,.cL'Xe.OU9'>]}#i$rm:,oH`~0K_/K=7'YS!o;jJ+\h9pVg|)K7;#J(JgO
Z*`~zF:EP|
;Q]8x*r%T#j+UAR;?n{9'[@`'HW>303kLsA#HHxy/j`B)P/If)JZ$X/\(~v\^"fpIs**_N:s,'_MS M]BsKMk"RNT?EHoK$5rIKx-f&2k{JD	;@})mZ)&FEW`0:o?-N(It^`f9y%Z[IPNg3vUrhflNUSL}$'KI9NiW"*gg-}k@}P&`,|V5C9_Ya?s/0Mu%G98X>	/yHrna.R{jF69QTf7$K37fJ@/%ob?W?`8?&V#/

l"U58JNo88uHC;]I)W=MCa|9l?3*5@i18 >kkXStIq;!}wBo,wPQ7~H'`$]A?}%Un<\=tZl#*
^t@=fimnl^ik$!Iw+R923i,\$54w& B$e3yRri<vk7(,Sw"f[(>>)
XsDt<qF>Fx&E[p
t4 P>w3%+=;[Cf|G{R;[}B*y3FGl8TK.Vt?&Sa*v{da\&0!|y9QY! Ki&7pf?Df`j$auq86s8!s!:wczN9,FQ[Tmg%W:>V3Oe\^LZ!=U14($d`pA1gyIdGV;f=6FD_l/7k,a m(gW$kKKL@WIdIxAI6o@7}vdBm$U8,:1ON'$9w~b66Ww&(N-	ST!6MyA%j5)$$1{WD/LSbU_&$|]M|;oznm_p^NCrXN8P@8<>3x%2I0"Z:b~>)^7sxs87:>~omi@p~5i8wgN0pQUP$_G	vsiT+8?+M^)PuCfU<L<H(ctS](I=nq,EXEx+fFEF'fRTfF{kgwh|682T7(V8`)oS>~T*
W	J/kA?I.VC~~Ow"?"$%92.,QEsmIr@B!I`)\oC1DD6N7|'xsMb/Q=FQhm\~%BN4zm: WzL3Y({<Y(j}GQ?5%Oud.Lc1ZuQ>f6xMuY<,@[w(r2=&2v5zd!g~yH)Jgru\=1I=:AAu4*Xyl5`\m
a^8nt-,{EP0=+metQ37I/%WxrVzW$
X6C+?dM=:@dW<6IVcnPn!#uuV0zE
D[a[DgO.']/oK*V}jhk=0<>cio@%^2E>ti5,sMYt._'^D3QZ_|^)h[tA9i:r6- "Z^$~e'+" ^3EECP)':Ri;b]QN8FQ/R;W
Q#WRnNmj\ZzUPO
GPI1mmgI>+Bk=. [e!Dt;]#Ib_s-6(EKI>J%a639T.p4~@TIR}fBz}oPGz%0I.xaZ_y!mBNc5Ok~zsg 6yWk&+q'@!@-cQ\-$v{[1dep[[P6a.*9p0#&(7MN\+}q^2s\"VK%>#6)~/-`pkWVNNu&df!TTB5.{}B_w*,CGm@Y!b-ZleMyBAWp{mL"*"zV7``_%J"Dy3P8	Wd1Vhrggm%vKy~uV':L>_gI[?*jW V\.!#$wbgC/.Y[[|,w-zNwKX$-|.!Hx@2D2\`uJ5@?+9lEffBV"v0LI 3Db9\?:fgLTh$mv_q2.)g sY+YPW]={V]r"+|45sasuB{0ng%r8,qgJ4N82-M$bL[Ay*/(&7G[45dSCA|~-kSw#DAUFR!i[Yj'?7FF<@u[N$/uw_1\g-`iN&O@WMN<"7=scV:(N^Yj	ydV3/*qk(`cLt7RLsI@s!CAOEky	P~k:Jy1j02|l>4*pn\#
&Z+Ghey)=Bm	Hr-c(k"g:yBv7L	mm&Ie%wP,piT-Z:"2d2)$~R6DD8Y=0zP	UloX.Lc/pye^1`4ENf2_A`XcDi7ugp |(,ULB?NoV3(ZHamYc_@v]WO66/&l\'y+-A&Y7*&Mlkyg'd!dy^[GLdq-+3!$R!E
HtK[nM] ,eROis_^Jy(mRc9vD1p[*Gc. M0c>
q++o9_0(N5u-	!V\8cfNDY/rHILvAnj/U=W<'31<1u/@6q[Eu%zclr-Vx3R5'cI,obf01k||nPRl($)[n0i[#(;)s%B?YFk9Zfti<e|WBO6duO/>/pZ7nEdf1n`cAcS5I	&5@8gz0Gkzj\&3o<te%7x8Dtk!Eikx4Zo<6=!vxJ=W7};jbb0$8mT2 +MEmd%X<.7IS6kq;ha
:]fiUjWtybwX Y:c?*#dvUAqw8*3ov|OHqaO`t,e37p77BV`}4w&fvBuB>JvT/c&FyIG%g}NT*h+|%Wfrd]X!mYr2BTe4&\I5K6$K"~&_n>SrLluL"k;qwIjZExLv@*LQMIPj<k-E)n?d:a@\R^hVAHd"!T7<kT	27%7nc[!kTBQRD8M:*-sNXB<Lb4UjqTav27?YmdP3:);`y:L68M"@Bj;,#/7!s")lUsm8mQY}myM<kPlz~cO7/@j##t Jq5f>z8f0Tx'W7J-UN$?F!-^d}UjTc(bHD"dtx":'Wfp,xc^&NvhHFXw[Nh`t$oy56CoW\J;T<Fg6Rr.}v'T)G~W`l|Fi%Ol:YP.`;XO#pSB#^5w}B!	,;X*Q5"cs	w"[]>&OGnT?hh<cTp8P;"\Tx;CZ>n}.B{pmjyKa eh/N)#Wz\ef>u0S3j\brx']e=?8{yZMEQt%Z4Nr;.5"'OsQ@W{"|)WNiAG9PNht?!7lp~J)3vOTIy7gn+iK;v{WoPuN*.#3x]@XUibohL3A~n	QWok8|.dacdIo)p!@J;zj=Eka*,+netDU]0
<;b-A'9zPiNEms"/)1f48+	?m.a	hN`c!Vn'5A4R-m:#-T K\>6pxq VigSN}\TrJp2 fQ0<:QV1;z#z7R(&n,WR:WQ'uJ5>V!?|)/oZy.P-*zS0[82}r'>,'%}dp&M	heFd[]"F{t!dMDE.Baf.")_]r8|/P`/J}rij7nY(jnJHo|LV{po}cF(=/=#^6gFH?yGg9?B,u\tD_-!IS8hCHu?R}{~Ox64%Ta0<H$w,#0bH[;XW!Wuua;`n)eDVMqj7B-bovCM!Dk\4%575*M=c7/jk?7YcbJ&P^!`=i.jWT!'f`f<'$z6N.RY'Tsp|.dfxEsgBU9QMfSoA=z&YT3{OKcFdb]Sp*xX	gIzMd7=&5$+}R.wiP\
v<)a)dT]e[P8\Q(`$KjTt(/IjctQ4M2R2jTCt']l)(eH$?gm&uKkbK_tyq_3cu$mxIw\mD/($JMwEl} i:JdfL%iO>am]2'if`0x	Z[}j5
ep_<;(u[*8#D.vQxw<[}JiS]_{2>SuQ|b8E:} %~iYh<"hVqpMh5g\fH>Fk$-}*6KUINe^+l
7/zx@NWHNk|I,+SSlBj"=fXt)[RuA9qsJyF|<9:eEe6lAVLCt\z'.:q[^|y=X7nB3]nQpljm.|xE+r>[~\&q_l["3g/M&J^K"-M"e[&m%E/6$y<zYOjf=_*	 yS.nsffcQ.uub?sGY^\,_%(w<TJ>~b_V20ak:1cC}J
k]W`l+qfguoKAmONDTL G	]lyP,7Z)_>rBWjmTtbB6XFaA%n'b"G}SM"<_*aFv^FWS&nR81L.G5bBoRTg?/ MTNaSQaktRi;.`BHi~#bbglHR5p$iuSPQ`NDA -C8O1E/((4=fPHK1,wQ}dF<% m6mQDC*"x&THoaXSWt3x#pn^oO$::yVBx/Y=b6UShN@|t\YZ*^+mbE?{Ul4iA8LG>O3"WK>]EMvxN} 9]dU"C+5797{w[I*muM.T];#<Qx<)TrN}dyOV0_~#0~&	*S*[[+&'^dI18gYkC2^q\}o"5s.{6O~VcgQ]0D~Pj2mraVzK83{;1ePK-Cw,+ V&t0I"+j;jOhF|7 P;Il	?t|1-T
^feKJFg+)eX=/n`vyMPzSrgMShj}>Tm8PUq@7z8'F9Bi7qV	_8UbI_*LSNinw*:dSUCr}'MZ]:xCmF;r._Q`^-|zM2MI+iZR}kF<}G}+z?^$vehxCom!^.h{tD4AG>S)Z
q#f);?,HUt?{Chc)$jI+#2jD_Eni@by"zo1)R[Y~th	[U`nLL7hI2SBn]1C3|\)ribtPU^	gr?z0H.q#Mc3a15oE;?-9_6xb~-5ozR[ZQP"7<Me7S[I~ujfvW'"8}!!#eb]pwr~zkdK@fAD.t$\!pE2GDH^[[S%%Nh|/d I59+ I[DqL;ERL&%Bo`b/,B!T#M`%c8@@Fzt@4zK?`I%8{dUO5BH~[|nvb=}iophP3aS-z*$kQvx^ZC_#k|M>t6NLJk.0s
O$A)8)|L;e4~)X^xF;sW!&nkTDSVV)+$~2I-.LLgNFHA\vvb%zy*8Ef?FHh+=[r*sv\F{,G(+'4BW1"0sA8)E]t~[DO/jJNPk{S'SCo0(Y`O?02q*F>6A*~mlV)C$V4O]`@V5=^3+HVp%*b9fHs@]1Om~2^(UX!.SP-8$E:@OV]_<::R#["c2ESU[	<B7xF0E{,2QJ2?H]e=ty8Ye_'X.F#{/YpLt/If#?[x@!TOOla/UbO!9}*K5jD:+`E]Kf@W5C_nDm2)QSW?x;gZipR'!LVIvd4T6	H;yU"nMy%l?.JmFo9r;2iM|S=YsJ^1wYB]O2,D 6,L%8&M%gmD|[WPR%Bl}/?QW|p0<1x05Pnr{$eaTG\j&e*LcOM3C9a@/=^k[)mQn5>?YP8H+q0nb#uId?!HRk	C[R.	_+fdLLXM0au(/|xPeR"@,2QB:/{id=9xce}Pr;"iSgpr5!u7{1)B9bFF-=(%z7HV}=H0,;l:pD\Td#1PQdkZ8a>!r415HGJHx~E?-p3;bkq_+?6XKstxQ\+_S'C@e~N:z77`upyFw)8Vo-p,x?9A^G ;{v@8ym7uI\}B)0t!F$ixsTNbZ#{ySng9p;?5cTQ$ZG/Q$]z<IIcEx3B{r]J<g_V	,*Tgd/j"iVm(_c$Std_>5e?9V\WcG[Wse6XJM681nU:?e,sTH`iMk}1[ccg1mZ\cVS--0&.BgY]p KoClnH=\(>V-%	<-|f%~<%N==>bRjReEK^'g8^Q"&[\XBrhJ=g/.XNg;Gxbca7UzG\]U2x6CiEE2!D\5n}.	EJ,]/Q.Xj55L[
D9a~Sb#pvQ*`S9db$A}:wk'`iL%i=*gu}WW}_
^57SoAxf*m=a/&F7pjH	IL`PT 'ry9u^)LT]dC0GfL++=+>?O`!	R;'| ^<{O,WvA'ReOc_x}f%$%]	[r#&ris5T7#}DM]_U^>
u6_4&s6l`0/%Sn?E:;#iI5as~,Kv9{(:e/Ge#dvknLar,pabtR=e.jdfR<m#	RN>nA:bf=H0	\vn#o'Ns}i!U u?:[U9jpS}sM8K-UV}e]>6FGAbKp-34.5jPIoMvLY
d397-W%X-*P%9%ltmu_yZsYPY)o2M10uA8;n3MNhl>;bKl~'hgBS<3.*5+=tXhJ(4J6q_YPY9n.q%dx\>wR.\S{qti}5kc\Y-p]hL.5PZdl-VX7lU8@ Ac0NlwPsok!0kNV)J_Bdn\>~iqV5r/Y\kC#kxe!VIT}%mW x;z~|\ T/SH`>/E@;N
}]v`Ph$	4vtYsu#-GBA!Cs)O%tO~YK2Y<CEvF>yOhBHCkgB	gv[*>Ognzc0,/a+y2{b!-I8)x$t@bd'Gj19Y/%QT;p?%nwhUL#FNAvmHuZ:$E's*2Q?IBl"kdG/	8)7i&%m;UM_;	IpRqxh4w1-rB&qoFLBS 2?Tz)Q!=0{
C[7zDFdjL}\d>E]&nOpW?iz,tZNZ$"L&oZia %pcKYAMVZ3q	9v
JY K4y)y_t1RY7-Ddd|o8]7&?][%j3whm6nv4;7s;lR(@}Le1@8]P;|]8y6'# A8fm5$)We5Rh\'';63Q:?blGr}buGYhsZmBKwK>o+W;`KhvkDMSnh8f-B%u'_iHH)5;%ds5kXkQ_mq":,pN7U7g'V\@c+.$8GNp``Mbm.\!	9B
B0	GVA"{5p5@i4w<2KkkAL}r,"vicR"H))#~"6M*wd:lW53ai/{7FrQ5Ht9x*9]M-P+=*qc"+I	]	Lx	SD}cpYT{Q!_)#H!I/Lp$	
eqGCHE'V!%i!I5DF<Yy1T0=fm<B50ePueF8de7"*c#@>bbMQIFALRZ00U1c8-,=_.&QcK$KrKe92.=35Rb(U&q7TZr=!s2RG	4KiA]&-AVLN3ra_BREp_GuZxLdNOb/0Om,r)4!w4!3\D,?>FC4t,x<Os*Br\)BW(tdOs66N$y}zXHzS
,:0eLo]oAm<kQrx_I]+m`JmYfb.;+-tra<hW;J|R6)x.&FQT){@GQd}4:GK3m+h62fTn^Q+{^G3;
cO{m\Et	hw*Ywu{/(WqS6s)!UJcg1F@<*~(8>E<4Bg=|wOzveoPf16Op&AOr1q35PuNloS$f8o)q\1!+;t[G+P[s)Y}-_;+f.5Zq%q1rTA)<3jYA5fwzTs{UgCl&`YFN	!M,h[OueJ;HYw[.^ISIzDeIAg5"	.@IY;KZ|} >!f>VwDWZqMl?"ER#3pYcDo.m9dkjyKF$tq/}Lp_pN$bf@k2w
cPdPmIwy.7gO#>6*?EB& ?5.{<aHY>3T|JTWFLk5ok\^[27k$LT)vl9;[>9N#I93"TUYxnwerb+i9cb(ki"Nm95jqqOaQ%$fB6$zBb&OXpA}'cdvV1K-]Ke-sxgB	L:+*d8"W)D$Rj*jM#7Iw{jv)/({xZj'6bD0QX*WKcS |fq:}AZx+l|cC-'_]<Y5F6U!XK.P0\Hw3m528H?1J4%`JzpGJW |c9t'j*F.,+cM<bUm-("IKT?<^Tf<2d0wTg#a'Tar;i*=4Kx#i;1j.BiGD37{,J&bRD09ZM&R8!{yDbWEjWRaP2mKyJ7l	uEX(W-hh<g5cit}H][B+6bvO6I:#-B%yu"hM|gu`Iqf .v5)nu=A@\2j#_ d&Vzd F>:j!@)aDn+0eo~XOAO@@ktCQpPLp>Le&`Q0yM+,"V(<2IaG{$k?(C"l4~#?T#2b<nU]x	
->%<iI'1'N[gdH;zOu99 @ENp]?hne Ulp#8L:x8qM)O$nPoM23&Z'n5oOc|gQ]LZMP4,nXM0nx4|V8RwMm2Rw3G^$"bO6PNL5OsFK.o3=jUTy'o.qTcX9p8vqAZUW	_py}[=-"{Hg.XC@TK7r!sIi3~l1U`q sU"E	zC|,.j:MlmGu&pGmFke4?]7@+>8^ `z{4*%w@372xB,YA+3TaKwj mI5ua:jHx2Dx_8DQ\\=Ph_s_Nc:uHg:1$0B#IVt,	|oWg 3;IK|lAEqpV~)>:_putO,*2-OA#7$zf$nvZ<V$/('&MBzlavgp|f>.5G7;|5[csd^A#o"FnAyrGU*<{,u'ID1B!:<ir(xm9r!^8D}FgEJAZhrts]6:;!(>_	OLe3>VR?}j]Tigt\*Zt=*V|18 j!GYcfniNU
h(S	D<z|}Yw	;&&:Y&p6l~lp|M]uRoic7sue|CRN?H]8fsoUv'KSuB_Dps-{ERL;)m^}':5s.X&kv7~Q8P=ix;3
EHGI#".K;rQ4C<8*4*Kn`-.*;;HmB9[?lTV#!5Se"/T}]f+ta+^gb$pOWzN3'A6LhJ_H
YBeLwo7}z'~sV!RPImnA
Z="gno9ZT}?me^%TCXIt@u+d#rPt%4=*3_d06z$~s5|O >'MIP2ZZ:R}Vmug^$d,b;9Vtu/A2`E(M7\!+AvYonqy';pR/Ig*%^#H<).JK+.&	l<>hvjs|mdwS:\	4\LgJv>C]8}-$S?J~:yRAvo&P>YEyR0DwzE.VH)`xHgTAN bnJi)D,3g@X;y-Q
*\^Q:[Y.4gt^X+q,?>FSR`E8\|Sph5
q/lxn/rsx~fTS$IJLL6?[GurLk'U&	%DN$iL-&>[,v}r3JAb0:sh]$,mm&ELNVLEVprU_}5ZhV,Nw<LhDP(muZ^qzCMZAf#V%70l)Kw^K>=Kf	6u[d0{JY/eLhk,yf?Qky)rOHX#ruarzwFG<VPdU?BCAPGc93[DsST]vhnKSd\!+71YuyswQ{'[7t;Wx3-Y7Qimk$W4&Jv'Rx<WLc7U5(6"	^
vbNwb7mv,|{Zb'jw#^hmOq:7PsDa45QU")<G=8Sz:#ytY/^oSt@zx7#o8pk0c#:PI[%}]#t+wiCRIA2t;HR *T|]Lu^W^^,/3vxM%m&wYZ<=
Oo?.xm6ZfQx\jRTUMJb*LB)_&XQ\1,q6{XOb$&kp/;M+&-![D58ZEtO0)GOl5^H'ul{l5k?3+dCz\S
&I?
`3a7Yee>u^k.1<H6 j3_nFEV9/ph&dJee{x`H?,>=Fn&9!|IU *Y] @ArN<m=B)W~=DA35WB(esA=Ni0vGmH7pYe}/ygEkJ7X?WkS'oIhIi5:apya-Duj\cGOM^0:vgk{6vW^MhjJl)\mO~T<7clw7S#pAp4D
3lnAMy.p&uo9ezaLmEZVVXv"Q}yQ`H17|6*m&75C($rPw1WV5.1bhpzqe{O{k,Jx}X;3o[\zkuPO7$?8:*%:<;utfQBM eh7s]TV* Dn%q$}K/L<Ird<ufaJ45Y&}?sOhNafjK0o|-i~<HT4P+ZrCc5"DquYc|db-pR
gYMSC'FHEu~%UN`3B${v|4$?'8S>EDj_!cysKEdC5>/N+D7r%=#jCz+~op=zx\9O-?!0oU
f[tJ6GxZXA~cGYW<)|*MsS9HLMO|R0H11>4qlOpq7((X}M7.{}GcXGfi<Vj_3Ph a70'(Dx/I';f7370fsB2 PB9k~,`+msS;}Qr6>6ot}9}?1@(:.\|Tr7Qe3059Tq9=LsPEj_>0{y_-iIjRvxzk)&Z9/dW(Sc.9^TT\CNJ(8egBK8]}crN6j'Z9p_MSy>UEXlQlq^TZ+?aA,!}2tE!}sgt;yci2^cjCQ1
U^"$X.xZA.}^Bu/^}o	&B2fB\lc@KZ5ctw<pll{WBZ#IzU]h/j[S=G{2%pw=ut3k!0V`EqiB~Q)h,{c.7Y*v\av!1}`uhy)nYs`hZNhZ/e-^U##7C SJ7ki[?>pP|q8	T])MF	<r)wE44}j8rhDo&#=u\"P9ARCt@$ 1ulewA^J`N' '[2R;X*E'	oSKN<qB17h0JX29{90N->}#!E(1&W<7~C8[+*UwKH JoU!JL
x:2~0eL=$kECl)}}rIG5NCKo=\!Ave]=ykWJK$\'c'6>+k==e4kI.G}^,FTzjfEKVG_|l W0y:6=s;J#4(8:N&,FlDWc4\6G)O@S1lNZB%`H&{>xQ#vjqKn2rb E	%?mpkk5*-,:{Il1Zkq=pI6F"}N;
N+w,l%zjmt_%6UmyZc#'Pm#B!o S!{h|[Q,%|[(PR:BbBrr//e+<bWJI"yPp?x.rg)-;RIl?v`	""h1\j.sTg8BOl{S0<Y}Vxn[OMGe`\=C%;FKXT4I[MdM~W{Ii;RS.b~a
,]kyu^DHR[%K[n*}PnpFnEo@f@BMGhfe*kRu;R}bN;7Lr`PD`$5 '.4I?KE5\^hn-kr/"H;'69	_3gb9'yI`
kK[KKj=@ B{K|a\bMw96IlF1,7Dp	@>G|CpF}WdZb736{njr>Bo8#3uu^
s%E%^smUC8bbZadm8>DI:7mt]L.R  ,W@ 8lcm02$yX =JzYI~O>Fi'l+-NA`+LOn!]_P9YS2q"M<}7"V56}=9v_?Uv)k<)UV3
,HRm KAE>=W,Zh80cZzRY!"_sbm@::pVj,;
a		RGOX1ziEAy>z2yZO~ZT#5v#4Y|z?u+'wXj/abCpA(ENi`0}Rp;0
IaYMF'+C2l[,njcH1op5rPbpYEN0j8Wvk';@h(Q+9~iUW{_!<<.pJ)( A\m{j_@g\	((<+8T@qqX}n2vCA%pz?"9_w?R}1ZI0u7dJv1=]0fg&:0?Rca(kVk!e\nH@z/ SCM;}7/ua- |m	`X9Oe\
P?W7kG|j~]O-Z:dVCR8m1*G-P2&e>U3
"\V{;n)aos{"AvAv2TC;rN@h%;V4X3Vl$Rmr7G&UUI-B)9/bpJ]fic]-TBFV3x?jI.kP(}o!Gw@sj6ARy}01b4VSVB:.+jMWM,r;B<;e(w02Q9/Xw"CRV&v^SmBugr\u{}942gEW;P>2@%DuL0n#El;@J_K1$U]|Q1$pf eukjjC=w|E25H;3cf\a(!;IBjMF.S*G"Ev0"?]]})B}|-BvOBB.BGn3z0|+[nN)?Md586Reb,J8k^*AE}U@t|#B-v/|SFgf_V_p9A%
ex{OzKnZ#&B'\xk=grs;-!@|Y04D.X8A<0U&WejJ2DD6]Uz+{KR=Hfil^V?Opqd0^4" 
U0 "YC@'\Zyn]N?d;kbJO!n]oaZOr'D^E`]X#:>C*(R_/_bN*4CvFNo.U{IhQ/g/KK_+dC+\u:K-~t3A*'E;S96x`rN@!e^SL}aHrK&PRrrxQ&fNah}.YNVIH(;d67w	Pi><ipWzjwYIk3LO^QrLJGk&8f@mjPx|R$6AF>75O9_-lo'|[dZUSO|A,_
xbcBgT$'TV#lqSSc_6Wy!v"8T{p(@\N\SiD^d'1
\}4~v3qNpu\	kuh2&DN8|--E~bg]AVPOX|e;$l:eja#7a#fF^Y4\Qew@6xT$^;]6A~#Nad7r(J@68Sm][O9ZQm-,H8Tu3jh ;&#XpjCzX	YN)>tlCj/C}\%aPztwR,E&a}h#n$~n|E\H2{:luD|*"3T.o
=PALn}ez_Uu+;xp<~]=p0f2toon6
_{<5pT~92lQ2C5_8[wVItG?U^bKuZd+/4f~YH8>n$O7R*<f+I
3m58[Nuocvtf5^tyn9FSg/KaJ:pTB1l]|2vb0cR'{.:_3]1h!67$[X][IE0~Pk1PLI12)W;3	^	0UqA+5Rf28P	b]6"uKl"\C=&/X~mgI/fnaPLR-fIUp!y&(vok>^j)y|X=qRAk(}ZjUx$/iI>F1}iziq
j+$K&BVD^
(?[';{6F5m#i"wbq/J#-v`EFQxlQB&.k@0gh|: w5hG}Q(/YBG6&MHs< y8/{XYF{WCnuo'4eQ3C"!]M<zaTG`P77r4w=<"Ht#4$~E[9Me7b!9`Q0%m3>Z`[Ex2:(JqDqsNtDHLnCuc`~oQK;~#R/Mu/zy5{Fd5j^ c1'Q2"o/VBE8
dXh2^?*6_[n<CW4L{?ki{Z!#<FJU?lH;.P;ZX ]rM
x'r)_;Lpq|EaVyaWnG+EZvo!UQzN3g</Cx$Yk08iYuA@f+Q}B|:F/>f86d=J\.Ii~5ddeidz~	3LB^r
!"mb]D&GO$e!+cBL^"kzx'-9^*&C5kIY%e%?0Lp^89Z6Z_9\5H/7RLWL3/O8l7^)~f$"T5kAQOY!;QYE=Or)k:hd%rBfS ;3**X_/lTo^}DAr/i"
dmb.@>,5PwL.7:J!j6_Sa`z060xT{5?cI.KXP+N]+iK}u9oLa?7:k!F]wj\}$>}7l0kChIJ>.{x/(UD2" MbGu_Hn,f'xT=G|Q8zJh4?*Z]OJ
/:vg_45d*{s$]tl?7`ZjQIuk~l&4,hPH{!6Xj:wSL3;F7pyX)H]?tbr1Hdh.Ah+>Acd,gN09!(b!}X)tGnkArW=ex!Ov/v4;/7
:9l,i&{5Lw8'ivsJa}jV$2J(cquz_yv)>x)Z
}LF}KLOfK6tyCA#|jTf"%_+{hh\MSM(q;c(]m{PYDHSKOg\@wm{Mkdtn,rDB\KNub~687%]yF"{VH12X"VoHyJl+gTUYCYYRu3Xcakr%F[<vRB7hPEJDbW\RFU<dpw]mx#,#>gWy1N2'8"P+wx"iBzplP*Sg~Qrr{#^*c ]s^]A0;bf
_j}Wb
[f_>\tc ex{IY#*,h0vjXJ*lcz{)G'SwI8V].XW1PBBp1M{5WLBNWpoD5]SIji5FOmS=?y&S#Nc]5%'GD8"@GO)MTt3QC8vtU[a I,.'`]7dNw0:B)?eYk&=y"i:,L;Q,I+~ogn2~~	wdCVB!Gu9<mrmx#9E%!wJez+2y$	*4:UzKQ[<GyeqJv|EsgHdo;B5rrO7?M1xp,WQ5fl&WXy*i\F1'OAkB/#8`HN/PU
;@^\,}m`o>mc.h3"
q9n1N~pi2s~`,gcg|=!]HR.%vX`]k7DKa?Ujk.y.og%9tObezgX0|,
pQJFNi`sf3z!!Y0:DNY1K)?&<`Y)`|bY'K++.=Xc OD-f30W{a&tS/&czQd,~!^8uQ[C}E<P/UyAh3x<i
<`Y-Az#3F3S<Y!Rz`D{L`5Y)!6`D*ny^h48 PkJaIM! KrHGtD^sSq,0|P2(_.]W-*p(ZUf!bo=*o1_?+%caM)XCac|YE&4e"F0pSTOa9{E)]1vclf9;)]t0}v,@AlUp.WxHgfLhY"d+#kD}jQ,7pr$wT\.V_~-!Po7-'DAC'ICUp&bHXKMIpr`+ef><#!19qES>>&:)A{~iwG>cauJ7S|t9`Ne}F4_kQ 5aT!26,oyR}5l	QX\8?DLWu5W5}EK",y$e.VQ|^3rXK}?q*kDbRBRnM;Mf<:Yyus(uMY<oNxS:_@47mf,!Hw`zqv0m1-\(oT[	\PxXRzE5Oiy8QPV-g)hD9/Zdb_?`uX|U;8.36mS!A ]d WHgo$Hnb9 |)og*20X@c=GV~%P+df(ZFS"F@AOhqBU}Lud>bGcVg>;G`_<PZx-T]B^8(z3}jBryWyiQzhhHVuB'769p`[7!9&+<8D$e/Y>r+YB^x"p: {t\{y;XoC=A5%)>$V}^EG?&O]cy,ILFGdCrnV\&0_7)(f[B5P?o:NTN#&,sP>L5/_vv7a;g;bEFYT1~.An{2/$lN<
d!&#_zYIBXv8P},5<eGq*\r<(F%BfQC%Ui?$$"ou:+upB(i(V`@9r*(j&I$#_Z(l~exW6vpOwU{73[9Q/WO4*R1c&dclVjX?4S${U$+z>mt|6DDx=]8DKr>h;vh-!34A1d3 ^Kecb{Bxi#64gRdM7bVHH	c`uT%JHkyB<+'ztd$/QAz.<!gr9-{nY=	jo@.o,Pr3QpfMC;O;-K-%r`4 }	<>CT~/VT9<7 elCZA#@	2q>PEF AC_"a<'.$U)c2N^V+essvrc"XhQhm';$g&1=-Pe^QUje#2eV2ki?a9tx`6~["]-JeB1%pLYBwkYPM"ByD+M_D&G`4{k(DGq6_U=eq}fs+v5`2mm*D'WKmgH/5dYFThQ|j?#SycNAYu4&X+0wy%
H^rRYV-XHu%CN350qgx/ovd;
]J(XV0VCFCDGLv7q1"3m=T{FulydMlVuZk(!|;So|>k'FT0pqK9,Rw/a$WyQo u?$(0B/2/K[@nS/T3#r`1CKso3nNjZax;9Htn(#_ $eB/Tqoii[;~to*x^'*lZ##y-|MEx[hc+p8sg00&NMk01@j]|U[$'h8K:'K4UshYv?"bt6jmRGF8Ncf_{\?
k{C7dMrqY,gYfeewU3+>s\u	%A@\DW):mh&U&,F^{tbD}3$G+%$B`+,afqwHP`RbX|[((w2jl[xLGZ-^uU73'i-@:,B?*;=;y*_I>Mif+wW+aqbFdrOM#rS<^W*:QY~5j^JNB+PUKsfn`]8]&1DzL,W<C+ H>#.z}!n3j/ ;3)qhm^dW^1qScX~}K\=`,nEegy'l5wjM%/Eixg Y8Cj{ew><V:#Xp?ijw)+yy{1S$%y^'?]s],vD9P@5Y
o}"%)ZI$&TDHk8Z$`l_}b^R.NhEstK3q$~G8jQLJmW(CpV|5|fa_`u"?]Eko@I\eNb~uVCK|#WOQ:4E9nLqL2<fa7id@!<mO;)*Rgntg]6k'5$#&q57ovJ>BOBowN]H|1H*YXDy6-,vf`lpRk_hCf27 iBMG"+IWwSsDKlG|iab	,9MKG4	oc`e?JCoz,}-\0XeyPtQ?V2CYio-Q7l]`y>y$0%|OXdYwLp %B^odh +/Cu'fhC&I{!\nOlBYOJ|FLKH>uw+i49#M35?$b`zz#R+>FVii0p,u[:uevY]-/xol}*L<O1BtuI24_Ja!'"*h`=iQ~:?T#{)gBLsHqN6
:bp,3tYXe){;_afd7'izt]g"z^C0~`'!3GB6t.LdC##g=v(X_n]5tMCfQ/kFRu^~*dj
GaTmjZ{Jq (AL_~5jK0.MLf>	U3f}6P2^>}3H?}4x]8/z}": rWq6}x/"QG#@#lbwcSXc5rs%mJfu	+X9o:;!TbDclnd+fcD>6"4yCm*~b;fMKGtWV?n&-IX:<wM0(+>\"q;;l]S3{xpeU
N3%g)Ocf}	kR
""*AJ`| m{Q^S(%2BcG'g_qB78giQ^g_J,PI"Kv)EMceTvS`R#orCAm>:(
~7Vd)zX2LMC=_ib
nR"'G+^B2'IY~2%Xs5c wSa2\f^6]t9*Y4Z?2\X<N"U%\w%n`o!}'->^D_#W52]O6X3u`oJmd^eH&=[]H|R_H4H>"*xP,wow"Jdj,
lvBvzt$}p}fFZ4U|=8$G[/q'=o>&:+<0,$p:>w]jkjZ6!9`${WjoXgUe4qR[yt+$YjYVRs6|gHD?a+*(T)8Q|wnWYp5v	T<q\!eNK{SN|g{I|"X{ZOl-J~*DW\KJKUf[Ps@2i[)eH_u2.[=TmZWQ|8=s	oG/\r|$bv:w%BLro,G2Ksp5WtKS-e!&Z	K!Sv^AU!8jH1DGLUV9-N=Vqr\_:n;[oE`~*o@Is*6DAn3jJFpgez^fLl<`p44|5\M?vHI8.4(<|fehyrkSCI1!}$VY-_g3!Uv>OZ1qaKB,(#6,[+sPhJj@ui'>~dAG`OQrttt\qK5jh]J>/g.tX!_rvL4=@s#8vm8"%Yr.!GIp{Zi}=YUNxcoAjP]?VR~(T O2hW.;4b	sD&D\)+^9$IB.l<lW_;]U159lVaGk
l'	*[>:M{kzh-zi
JkY$J?YvH
,*n_7:5pi_H|s6_*M!yh[-<:6j?b}R|6MA2i]g"ZnHvr
&LDFDCu:J^DuayJttLA8Z]ryV7^1AcZX1GX+/W55K`, mQTCt%?]Dq'f54:.O,*3ftPx`77~ i0,1;]Od#Hx0:22"
mL:eu1'c_64,bTdK}x6+l~9X}vrm:|#J2Xgo	/Pn,fE+}g;yZ)k<7wP1#1
(z~ABg9(=_cor4J\R9@b1?#h<7S@vj^nW>3KE"}'N] Wv=EGdEaCO2gFWdRSC]#BN\*;M&qM
aodSkW'[V*{M.lBdzbZ";1&2aw<a}jpkLPO`Qk5.$\7AiLS8/LX9^JC]?~>-op*.l_(<`Z%\YZ6	eIW/e&vG$NXp08vens>cg"\#oAl#F456"?@f0'4Yg<MWf>>Q*2Sk4ug!;mdSw!"#=BwP~2^%I2yC"$my?@	_}tAVl>/??l^]a<	0^Iq?SLsoJ9S3g.QQNd2wENpN~|+r;F*Ucgh)I+;21;&'
&]3Ofp"oQ	3|TTQ]YVcSp{H_W{O>!pKg.~zWNj/M9]B	w%O.x0Jk5Ob?#eJgFE{-NW:XS)\IX0>m63Afw7O5XyP4]8!-;iV|+nD9qI7\T"[	<W,%TZ%G$mNd0.jbj,v>'EP1$5`IvVK"`.eRD,s41,!waf.Ml0wN8</Y6HM&'fR4&Yw+@]1qw+=j-L+\v2D
`Om!X@;.=\=LPB+RCUc
!.LqGQ-ck>BEHWbt|2AVV3|?c P,/d9
(i\d0<M(+U8*	wdu<1hK?b}MNl?]b'1q~]1v!f}vtvw%fEIwyDdBczr$;oQJ*jzOl&
T$/kgjBu(:m]F`:[<{4%o)ewKJl"+D-}Yq
rKh}]H6N5Ef#)R^'t\:C4x<C3Cb+{Z~.,ARzSQQ$X+jzI:Le[Iq=S;mdX?$9~/Q;4Cu1SkdA$6s6D1c\[GQ`vN!H'.w2X=eLgQPIZ]1b?..Hacyw`RrpgBdO6 p0qn&SK5V1x],#&\n#7"TFU?}t7ME\-5Tu2^K*RBq<XC0HBw#+h0;FXi>;k>
ZVpYrX;09LlM7kM5j]m\f-7*jc.MSNt\/l-dM&\bcL1/^R0ICH,uw$NTdBK0%,|INKS!,#V
39Z/=ir,mv:&6_|9GnZ6cq:0-dc"m'2PQiM?$4bxEMH!k]VD8g+Kb"N^dsp7JB:`oyBBkUhf14qqL7OUrDW ,toK~D5
p	Tg4[,8hHr%zO"=|mSq?O|)nG{}GshF`A5Y~,5)2EC!Qg+Sfu s)\%:Y6[kt3%P%KyF'5.)Z}=)$T``c.=+:[{0=g$:QE=j0D#,4u'6spLTs~UZri<a)!?KomU4,(t_*6/~8`1?&vE:*A"6<@*[nsv3<w"mMkB31d1[v!)gqwOqaX;v3|tJa;\(gybP#}uYqjs[0h&D<qDu5Ql8Sa|*e7j,)jOhrH:Tw<TL7=5Tb|~Z:@*2k{9)&2Fe(D0E/]b,]SiQKdRc|.f~?|FPV/2],,~iG/:[A ?vB
^2<wC[;VCj6Hes,~%{9G*pWx@te95UsEW[3LjQ<O:%hd\cnYU&P9<4vbEE"E1#p"
6Eazxp~	x[T:-eV`\vlHqQolUU;L^No`94`? [mb/*[W5f`qWci_U}8no=aybRl?
^D3-DrqgO1ZQ}PuG_H+zRuclv)_`db ,{Nh)qs~un)*}$qB@gI+j,Svh9#_17ca'M)=PZD:rNR|BkZ`4^]bL,c`[S?iR8M39d@P#,2`ue7kt^GR	d
)!ZLF4Le="!?#|]n@YIa8ksf[W-hm4OZhUbCmaXH3n&@.+OL`OXp2%O*+(/;YSMxeB$.GDriAKeVSj]7	ays416nZ@{]('eN:F,B=z5| bSk]zsW1K-m2^2*eO^xWbYkTc$%Ym5iV	ax}9akST.gG'"z?:1\>,,2vXo.mAnJ"6+a<b6-#UmQH{Z=3,?zg4Qf|r=^WOtIBl4GxV/2_.t<dF_H]eO41Qn.>NDFxY$eXc<Qe1*DR)]oVn8$-'ld>X>I93J[;^xJA $N	1)QH'JYtKy1jKtT
c)/B-=%`E1R1BWgDoF[^i],mLv{0{\161LZNc$R|jR<<S\`_OER8n@rY4VOeG[<qf-`(o(IdDv/|wfyS=(ME4DE6ju7$v{	-;a1uJ|(c!Ny$y@:\ZC`}OtAa5<<	oa(Y&9"$g
;#=^!_Kb'/@mBfP+M= {.h?9/0eg!8]<.AZ8rl}6TfV\;S"E|Jo_s|'L~{qPx,p]UO(Ize\XFn!vS{T^4gC3@'(,*q,W|<6q-F&w}bi#7=Fe'/>~
ghmHWy'_n	t]y}`0uz|-nfLXc|0l	ax4h[_;gW<zvX;gtOyZcCu{{bE76cgzj|`*sMI"^>77fe`=rZa*qFQ"TF*Rn2GX)3sZ^Ibx-"BN5,gj~FE2%l.n8-P^#Q1Ew5cKp3nY#D-<_0;L<PasbXoa-lqIS1zSwST@ DDj]nH^vynz?uF#xbYE-/gYH:S$PG:pG;I17sc7a0q*#XtucQocdgn'aW393Rnn6*8PIbSEe[/gyOXDv*Oo"cA+(\UYgV_x44fV-VS_~ @=nO&MJZddvZcvv:5>e~:b}YxL[`tW5)*Z>6k~+*bh)<ec+_5|Y*P		.!oOpK7vfCejuJ	,5; 4M|Bk/I9~^{L1nSZXt?z`[$FK)_`6k*CA|'tCg89'	7(i5,d!-]')tkDeCNpbmN;Y2.t 2Un1Nv#-&Q"LS;2'j@d70f>B.l{f_gsyei0hSN`f9EJu%(1f1gTLr|V9Y9p)`WkCDGW]+jb<xt=z\.jjp_#VVEw/&%1b	iXdS"b+XJz%YYbr}-=X b_f7{<:ps1-@-kwr-Zl"?M[d]
t1%@I)&IQir}&[:iK1d,sQL.UuGgqSmngxxxMq`1`mIpQ9	]6-7(Jn7}=*^h{3JCt`%#BR_W@wKev/+7M^PDmO3RgG$uTgxV+N
r:b~t_vM9v'U0OQ}.g1yE)_	L'Rh
u9WZw]h03* #JHii.<5/e?5;U(FW8@3EdC~mepn!8?+.I(hqGcm\uf
	nNi.5qI,_#:yI,o]Vz5z\y<lv6ujU*%uC5UN)@Wa&%\I=D`p+>p@>^4hNc?WhBS<~p?,>]"N;J~2&  H/3;=S4PV,uCQPm#I{13%*`!w[.@ 7'#QehX8}yN0n3dlcSvXQuX]f_NN'PW_[$!-b[,m8FuPn ^Ft&lTfcu]ea(k]8xqE%V*cwioBL`\@r?9D[9
Gx)9RqrIw]5_lkd%AdfuA
WRwHaWggwmaa/2hsN`q3eOPj/mat@`^^a$To"4hE5aL6	`lL`b6q).	1lqj70;me{m?FDq{EE@sM
%dr7A(.?EE#]<f&t^FVv|KD_$Xiv/(Bjikf6-U')~vyZX_UWQNqM$GlGH`%SH2l\FZ^rdxjmEz_*';Jg2ZY"#2acC%AeqNjt0lL/wNsx:1[s>q,K:AvtBg6O86<ukgZCI>ef=M4~\\6%4{M7T2f&@d"R)vk)B
{!~JO>T ZUmPc<Y5|qqsHE"[V8h $I!"Srsjusc	T3$Elr,M8kuQ<E;GC)pfX)/k|Fmz"snP#?]1/	P^4ZRS$j^e_n8TZ}<1D'S1?\CoJ+q<^A#RPKNR*}5hT3'eBzs~5&z5D''0t,=8sA(nCzQ%X>da,;M;#!e(rqre((b\>s0wJTQN3dQMv	Eadh,CDkKB(\Rm0 VmGfO|yCp#h&M)aYtNq(8Bhdh4ML!MkY0N*D]|~
y	#5XX9<m5mM/F5xRB:0yX1p6XY=*/Y6],hl?R)Ev.BM"CE^&yVzs'`/1|LG^r7D 8=gM'UaNqiM<'dWYeuRMn;ci/Naj-HBz(NPQYO9oO V.um0PW!%Gw]Jz~f#WUvwxH2UZNIZR-]\I3ZcG(%StR_MA<n447"6[D*&.j6e/fnmfD_V{<hDl^x:\6 6*4CfB_$< xr6Dv{kHl[O$qfxo!3*s2"i@	FS,3a\fix1a@S-@'-~IBHv(tm?_q#QyGNAt56Q2{r}/nZty;L<hMk4SG.Wt@|Kd=58?
6mI	{x~D.;#IbI7bz`?@M=lo6u,	y^O[bBC^]	(4?'Vd"O7BLJQP[ucz[S{%CsP12SyqOe|!9jAw
SQ?=Bs>4Lg!'\dvDf.MO
H9%z`dxMG>ZUG`-3tdY$Iv4oUK`H74*FP4b3xV].<!lzwm]6Z52g4%y-nh:E-{z'O2^byaH)N&;gUM:NWp9TX	K{a+C-c"5LA7LHHcQZ*@5tRh3&_p:}D`KysuU(}HrR9adD&\NFi|20@hNe93Rf/BukL+%5-st*BR>$T(KXv!JOGQO@ar|h4";hefQduZ.qCs<US,VUdaT93ST+2X
Y'|>e[}X4M"@W"Wd6m&jw@@$+EV'2'uei{ADt
}*uY>QBBN&5?*[p1]2&q~Of[xE~T	y+8#]K9OjZb=UGr`N^se+:'>ZEpmt5` Y{UsD/yjpO&;FG'.	cVBllkE+76LSPq-\91u1,OiPF stz,R'4&iW0OPv`NRV0xZYK[Z#Pl!V;!#O*hSpDl\R+.$	oR
a^&4EXt7K,R7Y3{ac%c.8Crw9h}qDQd|'LdJ#YakZ>,j!ZItL"%G}+q<l^2?@>:DX28: F|Kn\ST6kn\`}O>w|iBi'CuS8}\Fp@;MD2[[hf3}@;FW9e)vNx<()}_@,pYTm+ta>^{b((?%c`'RjTXfcpeoJry~1{vFr<$6LPB`v&zf/GQA}
A9.m<RYSU8G!fq>'*vAAvE hb
^v/WGX-\<D7>x_ByDI})
yTN[4SvBzc^1rQB=f	 -`5:'$
-7%n2"$aZRC.f:1G
 z2y)NWLPD7x6&>o|:K[\Sd,]"nk?64H/>UxKk~hD44wiH+`R'h<HQW H01J\
=mCW
68DO`2<	`]z2/t3=(>4(	K	ANFbwT]8&BxxgROVjw{kx$Mm13I-KB?fK-@0d"g'Ia*9jz}ht;EzD!67cz qjzVFc5|	D!5CO0&6"jZ3	f<k+x08Bbvp
j.<P_vyyq]l^~lsda]NKDZ_mFJR?ga>#J-?,`5fn$DTH~z,l?&9H{DZR(P78pKx5}qwa:)A;uxKAsf<t7bY:E:wnwL;!OjEP_yC%tC~+@5*k;{:EH0a[k[T6|j?,jQV H!O>1"`Jmi}$N"J$)	eI1N}eqp
(b$S%(K<
3'rO`qUtSy8<gWij],(YM0-sQQ9b"EW7WEQ<XI.yw+_+X-]DgV~OP-ujR#(VKz2yr*<4S{|*1v>b64o2#jFk|};]}|H'|)L}D.L46;i[w_)k_*&zG-j#wX;KRLe J$}/PnZ#CS=qXgF
I3@e[ROM4`}Ui-}H3vOqUZ4.fx
>[K*"_^'E,DI.F%Ly6zkY'Tsh@7w-?Zi
Cn}}#4'< *@TJ:2&>F^zGX6TI}.1
p2V8if3>Xbaj-TDDa(]FZWJhxTL8lzORl*(^'EKB=e=DpF7H=	tTk6L@)rgJqm-z}sZ9r;o@5tvKg0IvcO`ZJKCUlhFla+a49z[zd#9x>*STXW)
FLX!cr5(ec.Lvi`2AFzm5<`eu1xW5f#Sez>;v.&l!*yTi/d|vXsc.P<JrQRvzEGONr}`}(^9=	4O)"owd2V}.v6
lfuU,J+&|#:6/e@H#	S#YI/q|L xe~=),f^wBq}%U%'IU{I]92AjY\#<So*?L+R:T3%9|udX#lE4+^~8HC`Va3Z8mqcA{NHt3;zEGPHQ?Eg.Y=imr<{Yo*CxNBeU8Y(w,	H[\XmarV]JhZDA]RQHH7d)*Sljrl\,\wm}v:SLLH{#n?PS:>Q{YCa@4^P:R}DX.~Ly!>v0
iW#5?MF":i(282%g3H#A]Z[a^oI9>8=.4'70'B+	X\o"\Rs"X i7MX*,IuyVPYzuXzql<S{29xA	brLIt2{G#PMb|Dv/U9(j6{V.S8G;Ft!6UP|t}-UPMlM
[S$r<\Cn%<g?ix	q{"8P']3kLb$&r!\]0{	 P0hm	[e{1{}%@nEJCa;X$;<ZX$^0KON@}E0_y%1u@Dq'1s ,tUCzh?Z/=c!k5\).	m YtS)&j]d&tKO-wj@LZ|KwUb{#+#v&_P$_ |JZ)TA8Va9-v1	gW7GadrRF`Kgw+IXsSUZ9rpifzUUZ,tL,Al4f9+&kXEQF&7aq~|,3\v CA8`NEI45q8wUf:qDL^: j`)|;\[R'ndeB-ElJ.@a]%7men|74HvJ)FX>.KBkMN2pFM#@]Hj,yjtRyi8d\X$*O;Q0nq$Zh-aA<^; FFaW/+jW;lt-Qr72E%~,&Xm?7[k2o _LaGNw#ST^^[X\&dB![l@kzFVz+KK.0glW:bLx&XA%qv;'$xW?Ex$qb,Ur/m8S-SPN	Ym>L.G98~}m;B3hduVEI&{pG7;sN;{e
=tNeP.OX&}ntr@r%Vk50_sG]?#mjA9.]N>s-K$0iI&Sh6p :/S#@sa
iJb~N/[*%$Gt%:%@Jn?S(sf<sd#EM@8WSHyg|f0|e**"*gAxG=97nz^3gmYzbpxHZfq!H5fe0wg1:YaD5`7MQ^k%)zL$qey5WzW*=Gv]B>@]7&b&ooj3M&BH9{E	#IPp6q&'  \+#@MX;)(*OV3@*7TL2?E:NTp4My0eP	nfSv# p6|!VqQ
Z2py~tytvNP=p:TEN;cu!rbheN$x:A@gNFFbj	4.4]/1TZ-AB_s]0jv+A9f>86$EfA-@cddhY\GZ\Y%{H<faoL5oQR'_"VJ%IM_c'GlYu$G(0=K#u[v<L/|G,C|>0(d.*p6Gnx'N?|"	\k
R|ow	ufWjWBJW*oAdk^1+>.=_2	J7yLt~*M0iqaH<xBx%X:^}[-K.!uz,v/7fg5>',6t61I*q%;,M{l*9y75xaf4
z^!f -9uzPjS>xHLRUz$k__UUm.zJ5C)_4p_a|f5RfiHex6eDi|~2}0IU';Ci,U2_,S\VlKP	/2	>j@L	seB?ms,48A	n-m^etnlU' %;'hgG>?K=JqEk+lNMJYLNGKOlhhE&+ZlCQp,0C@2CK!
)b'4_R8p'$(b4#NFTd4mo,n\$G*cjM_D-y 5y40YGqf=
OiC-r9Wq<FV}#+Tn=F.>|5f6:^yxb+aQsRNpLwC2,2?_\>-M$/N{|N7eDF5l{*Y/th ZCD8}6vI4P!
4gJ<?t:|>\	6IhzR)i*dHOP*tPszus >vIXY.*Ah?9Q@
,{'0
=+>/4gx9@ FVW6sQah\s7Y8jc8i'@&^5e
>c~J6g%
-Ta!j)E"FnueFa*@*Mw0i#nU(0D=,j-.>q`&0,')}aB75dq$6/ll:ZEI*B>0Ct{-JkP_?!I:wni%y#$+@p45*6kk`cEm%
c=	}la9K\W_jh{	Vv4+cT	AFI]nYtb.,2p;LHn?LQ]UOP5<W{q'qYtmEHR_g$a	QcR4lr,`S?kcTD?KfPCbx~]E`N9Ku\?+AV[PST`%S(v@_LuNlc!]aDEfY_6jM5WzT3[^cKX:'0{c!K=|OlQJl\<FlPDqb<Rv;\]o`S.hBQ1n9X`!	=19hFQT3PDVH&IK&FPu",@HA3eV15Pm3n jI4kv4V6s)@:FxW=_7 V5K!&j?Kw	BS}aQNT<m#AxD73Z312#}L=RRvwtMEa =!qiDgu&!OP\B%$xjE0jf/NJG'F2MU5|<\DH]$ua'KlYnv]i}G/41*cQ{EH[kQs]g%*$	jJ!ni}k],(q<A^Xl0XZShaB8;w{57@~0	!A&e<*|7%|1O	*}r!$#pVap3[T@cL%G/\" \$7/Is>/c
[(Wvqp)2Dca(!%dzi{/p_Ve,2>*@=gMzw[.dznz))7q(`g}L^%Zz^:YW=YSt[2M!0aL,ZZfn4++T' Jg)^HYfe;-g4,TbPb]T]x{XSb=Q3@I	MD+wy<6UJS;9GV)}$~} +2?.1$:b*.3P`*0%:aS:%.lhgr77;9G
0:&R~VseuN3EhG}x6:=R~W.>jPoFz\IT!eeJE%,y2h><1:`kc|A`c)Pfk=wn[chYGMpjRh+h[!r:TAw18gT""5?fDy2:(/[Pa!Av%<.{t]h`*jR"|11WFv
#w_^W(f$.n`IO5OE	D&^alsgtR${:z#GRC{306o
%(4{EBn -\ m}'zV^=Q23zo;j1X(-9K;>zx6~IkA.5UJ41Y$6Euqbg?d\$+Nh8.\QC*~};U(FbbS^cS!I$SR/x?B}hCo]w9Z~V-1X^9h[Pev6dt8fl3&/.WT@?>,;%,:QP@c6V.:_!aCL+hjo0U+H4fQi/,4-KK7BqT){P"HM26bdsFb:T5%,.tgO0 :FPBN&|"';zbhK]=G\|y`mDtjYW&O,7YQQJl-1$e2XZ/*HL<3.A$7,1?8:]G^v\MaayrM!w@q;h	E\}}P7UcY^mB$ku(V*x}/]oTPx^c`(>Gz.a&pqg;-WOxxNF!=rk!'FxSq8)>e}v*%_^bR=_&q}QTSC/iY-:.I`AjY<a@'-zjnhghvo3BRRlC:alcyMrbzvW
ny)v_\q-[J#K*M@hHz+!0(8pW-f>U@&4*EbqCu9{9Jlv]jmV5}UAU:ap]rcbG5P[&FUl@dHB *lObM&WTbZZ#q?<Q1|
)w`NRVaWHFl.[BDUBdP<wcu;Bi$>qBk.v8VOuo3X>Ga+|#r&A'n*i'"O7^{#i!@&*pcum|QRHk-?y1QzZ@SWHwd|/^"M"{M!\o"ukD}c
9M5Sj3J[W_Gumv'Wb[avqEys_5lt,!VLzdp#%=ncJ?o>QF%nK%pd'eY;G#5>&3gCvSt^X59kx`M)!p7lDFSaUKee}^bCu~QH	x/2,z'j|I<3(hxA1v~eB)W|x+^[a{R$DOt/cLA=]>|ccL"k.9QnF?738?l_0,k%UlrPUU|pT|kmzoWf ^N{N:;W>_M,w.$i3=X@/a.i#_t]Y`[`~iwByD.goY8G.}b0>?pP&$
GOQ;J )9(8X,Di#K9vh]kk5
jGLkrZ+BrqU~
`V>0^W{;ualBBky&rKzIq,V:9/=ufP6pUubS]7ewp4,A.P9A_Q~%7{>yE"y,veHSuZ)@sG33Zp6!ZnFHo!is1=`$']Kc^j0N^ak.+M6`%Ny0k|-8ry7[?'f }vf28&CM+;9jJL,`4I0N)dy2`Snkk=Fsu~8X6]iS.dcO`g6xyn~ZcFb)B\F;7AU<ZoR98QE_Q% V$>3zR*X^Ub,qEj
Ab!]I'/}%e`ABJQ=</?,6(+HML"3]FV4)N*Lr]obpi&Wz{<r\|Nsn%	S\:4bjSkC!QoVVV3`V>w]'_zFKRVDXphhyZlAxQzZ8dmOHg6;*[  X}E!]#WUZ:b5`:O7Ve6DHzsf-F*TL-&NT2 {>Ud1z4D-N<GXoO5y-)iq!UA<MxlyU\UD+}>l;x.
)f/Mb4;,2mqz'c4~rYurF"Z6`b
^?h|O!N"EsLISYgj!Z\~VV6'9EH`|sRD(|3?TTTg&~U]x\W%oRX)4YOW6<Ss=kS7t`y<r5	,x<x#fA(sFxKXq~Yd#-S\J^|K!MEBC:8v-zoRU+1NvxI	cN{p'_46}E;tmIc8 &*0iBDIT0QDa"+x=2#qaU4fFZX~:qIn8IdLUu!BT1'izi}lwFb}9#6H`tccUX=$oE@R>o~8>"m;6PcFSe~-TW,NRzsRE5A^}c`^/dY.dbPQ'Mx4$\QqU*H=iObJB|eP(PUe.0q&`c,}N-:|jQvusx8i6$|Z*),Q%eo(=;F7"B8@6(E0Y,gG"V$PEIKTxto*iz'enjs7t@1Y(r^AClR@sEG
s:yRXevOGj}pQceVSkRGomh:!_pqX}"n`ryvqCvmV#^@<LiYY_IZswwE&45AC3$r7E^S(!ifaP9=9b|}m%[R&?;yicar'MoopZ_$M~CVO}
)y%giu`y"xk%dz!1N]{M3%]aE9Q~,;v+]yeEhvjs|$#N'}_BOEA(<NENk;rX&kRC7HMHb8I5Q8`#3	N:^.'Z!mJd'YKLE:tKMOaTJCYv<\2C43Ti,lj>TDs1CN9%8{=<bWy8W5|p9)eC}#q<K{Kw^_3][\oi`];W- O|YJ:?ks;l&]|)p[>|L
<{	o[\8Np@>4hj-1>%Q$Rba];Hmxm2]9*X;[{MG6{/un^|VHBU !0QQ*QVe<]t4R4	8f[{*Z(]9h9N(+iyPQo2Gd{UDMGhg!mjRTm:i*
,jD>R4[nq
mICRWK:\QWz}a1ZrolTKe/'oDC?7NMUrBv0CnK3	Oo|;|
%A9PMuH,h)aFfY>VW"{uGzUe^tAj9DpL
YkCrye&Z38f/nt+7"skG@qs.;wr'/"$5pq=t:aSpNy1A_zJI
brhmsn+x=Tss;#'(G 6%	Wuw(8@D"oXSBPke[S,wlipF(g>/{=j/K73N$woW}[0c;^f0Fn*/F,9PAv\z<WR7}?,<[eSQi0*(g#H~b-~F6?O/*yGGCN0CSB7c.olv0'B~:T.*6GTE"oR9.^i??Xb!`p<P7+uoyNrSuY<dTd`4m;iNGx&8"fle+G?1R%X1=jPC
X&#lY9g!rV(n
G6I%Ko-Z~:h\h4Y$}zv&0G[+L:(`Xv7]$Pb\@Nu'q~r+>=RO0i>/b&coMB9/~"*ABy6)	pJ|wc{"q;N2LBt+6yFWjk/f<p44"lk$7%\g_4qtKQb
raq[XM%(e^uelSy?imI{~EeO?
8ZL51s\B229c!,iPPk;<Q3='!eBIT!Zf[Vh$qJCj-[o=_z2k~vIC)
b&Xkb^jC	kpG,F!b*@^'a9.Tye|,!k&@8[}/QLCYFG/'O&_UC')T?y"+%Dwx<P9t8}JQo{m:MpJ
?Ee>{NkG5rp2^Vv47&S/7uH{$F*K%Fq:o`OHE?q%&+wtJEpn,(pT
<l%a{P_H#IIG]%Bb#)`VZI.lLO;BSUCI|>q_|7]nnRAZc(Qd>/;)#r#[Ai$j*bM
KqF,$`8<MwVAOV?48	68v9Tj%L\TqZ=-v^H)nR<fs|9Q"y]GzwXx"d%F6i?]S&|K&&Gd>~+A>ymsk?;2)MPLXJ?8f,G;Zs!_Z^|6RdkPu}!4no3bnE$6Fp4G3H=9\IJ:/C/>VeOi&1qr_BF^y/($36/ b }A4,tS3Z	J"5H-,3FRy/S)rVPcR|*v7CmQ}dfBosJ	`_pSd8.E69zayb5}qPX?h1J[41].}DweJon N^#lNiA5~byZ(wgN0|pQxJ|Y-zRG~>z[92kf^	-(19(Zlk=ORo/`u@PfOFUH:rGrRibUH*1nNSEYa"7:12)WK>h
5{}sA+3Ke $"RgNk($6 N}{d8
w (>*4GxNWoR&%VFB-{KGkThSRU=gTHQgfD,poUm}Q7]!t0$PQ'TZiGN3Ns)+%O7V]yA_N	mMqrM]zkm1;&q|G$"T'Y\'P#o`6f9WX%hu3QWMgAK)O4hijo3bJC92Q"{69Kf{-rBAvl6Xt%\$^[lJPXk6UO`XgQ pQI"tjcG<u"|)<u,~#q{h[)r<3aewvGh^vdQE,]Gqq-o\8_/>cz[cC>:Mcy3Hh"]IdwUes't,. jrG2V;&1^7kAd*rZJ_+`#6{TQU[qC[_""s0-nYcq+i&')|~n^Nl!bg.z2yZ1;/l>Vw&u)Wm"CZ8h{qkTgpbKbECs?n,QJ'v/MC=,Ui0#Hq?g+svgad"Sq{GC$qZGF	(C1#H`"mq|7xlgtDG+eV`.bj+z=Sx>wTX+2z3lX_3fU6wN_JX[Yn=3ti_=T	X[*z$6W&Y+06_-jcdkP$%j2}dC])+kXn
@?T?45QopkL'Xe#d.xL\kn!V0:XlKp=)0T;`t}C~p6nkbrgX"*Kb)ek5:irAa X^CG.#Eif-Sr43!di+>Z>Jg;sN/`Cp=>	Lt|*Hw{aW.I/fmD%
kq4( Sj.URgTJ'GKdQ103]DQya=Aht,z}S4i8Dd9	&tHuGSgara)%!eiJkFJuDD*$g?
TDgg1)aIqoHk"#>!j"R7/ScvY2@ ChnwX("yJ|0Sb>kW)~3eRf'$|!r0<gxY|,T5oUmDPPZ[!?hFm>:apmFE!&?!+XPX/1@@	G2WbBgo[]8txPPp6@\&pc5$y>AJs4mP^i;;8yms#Rb'o6gX]y0~gs>Y;znyWP#\8quend[x,,8hynNpvfwrv)d2v+]lRQCL$'bB]}p<6>Fl}7K#t%#Y9EU4mXq1miRM@[h5z19m#2>e3[6Cb7Se{Y/VpV+BDh9y~"K$.<&$8D']X#)`%?-qSl&fw|mw#>:nMYIVO0Jb,\+/xp/zAnvDV7)FUnYr4o'Z^Ao?sW7G)d5wK^O5;GH`[E~6*4yR7
AaF#F^u7-=ggwV'&Zt)DgxdC:k90$s[y@K'"
sva4s+A_L,c*jJ044]]c!b6Cd5o>UOfe@'pVg=eogPOY?AX.|U=H./1ZTB|L{{	[}oA3n^pv'':)uTC<VGn&_0ubmAf)^\F6d}2utb^, mc&R'dPMJ?`gmG2*G|@!z%:Lr'{v"Ys*hS_*c=5g2!Z32})WlHeMfgW-az$<[k-qlef:'G][lV5mw%P`vX[Ifp*d:1WA'^i0	>kInu"1dQFXeAco5N{+,h@ }L[U<0Q}\Gk6@yz8&j#1@0s"m3j5)4HiEhCB$0T%^`rt3$[%}s)sr#n&Oq{>|$ns9aHiPZtz&xaIohshL.sH(x#G3c23W#?4X>e__cn8,4YaUF%CxSJC8X^<9)UpJn-\=c-H(^f`=$R
,1BR)%CBNia>_nR.`A+XOCJInNC?a'q}Z]jXT*pNgR	e
2H?oGB[CVg.%Ph(a_s]%8{wMm!>}cnw @/$aW9BGmHuxcPqF4/r=z"]e0^ubN[r"@<j
DcZ,YDK+GxpfaBv}J^<'UfjZ*v0G9u3+/j,_Cyb?*}#qJKCHR
7j;;tgGwzsP;(^+qBM@,J2KqL870)}YFG}?M<T4LBZ73VS"=,nmk:]Yp&\vf'Y8L$aEidtb3ZEMOg;&)Dc~g-5m36p+52FG?"7{G?i6=>,-[
>J,|{5	nj{X&K60ep(C@$BHztNzq:Dd"%WJq]Aw>m(dS{xaK#E>@z`;NF'w}[GO\"1T(C{ZHHxR:%u97NCkVqXw8"RG2?ZY8Hex-IPdG:e_Oj&<Sbxn[n^.Lo2c^}2\m^RXJ),@qd{MzD{Ygf!+```!9(EI0+C~>dTFQ^R!8l`UX<9?*-N:Sra/tbyy*%S_gg"90n;6xn'{9
g$*~z~/Mp7rm_[ksF=L|nq9V+~=j2	%w[dOh's
hwbH~;94QF$lYe}7j`qtg7mf/PY2};EO}Tr)Lyn8"&lM|,6NHpqxmCrH>3CE_AOvq'!~zK8i$vK bC!._BAcRUL/h#a8U:+o*tu,/1xM" o(<bdT6B_bq8H+|:;4H:$sSdY :XV(M_X"x2F s\5R$Dw`UE}O.|ZWHPx=1{Y$|KWtR(g"Pe7X+M`h,cbsA3\N]z8f}EvK*{Ao
p-pJLvQ/f_vG+AWrUnGml7x;X?h>E\s=|:q\S5Cy|<|9h?>W /#[NMhBV4iBo1B
@ru@|yH%mLW<Ptn%&KYF}>`%GgIh%`h-XkH`KD8wNb_q(3I71l-ue\}qYA@[C2>J\=QmYddt\fZV(tGhkzqr, j$>_c?<d!4.)"]g.!=>l`,bUo'I!K,^5DB9a2^fcfv ;~F]}=h?A~dtp4w"hH#z;xrQGle0(??>[V(
Ix,An35O62ywLV#;zmx~g9X?Z+T%)&<<Kq_&UrK?}j&C7Bbe7~I}~v%(!oZBjH @UqSSK\uZlQ)']?Db=bH!UT1f~nM5a7>p&^bbVpHc	;Uf'n9zFc|tjDN `aqb(d(nxUtVk:q0kgS@'b%}fl7K YiL*<k)IihR=s~}Q]'I4pm%tb'/TuF+FXDx%^IIPfW5|]z[{!H	,3OiH\y:PaG^{vH.h8i=&Zk_:.[gYF&BeV]@K ;tn4j%R8:ezbM\)iSG*-4$A0)!vdN&CJ	q$;HN8T0L&7Uh-CI}{^che$B	K4UxDJF3&yk]B7-OV|9;oM;p60AO{ j"NNW"5i;il#5g?:&E}|9C[s0+1cx}S*4#fiuEb9F%n.{XM>;/12"#G{_-O/R=/ly
VU\]j~\b!eZ^]k\(m}=zuK|ePC	k)$,kl.9=FueGZOn+"ORpoOfIgyjDY9c?hO_0^3+@qTu:;!GH0G/+/rsqk1N_;V!t@a96"gnSKE7"A^\94:i^KO>ZWBh*L""}s<'ry=.Y\7
,[,tYc5O%K `>`_\9xHhaNN*_`DR7<4bBGh'WcckLYcf;`{Dq}+S9cWq[Ij-nG{@kk(2k8KQx`*u2y
ZjeQm~5cga{;^6JcGCq(5eS\QSC%qPZ'sKC+tDY>GO\/C;:Lm <pllw@~|<1kWCN=LN&8`7)@ XC)|r#\*fMBV%::LwcnUM,Ysi&_44=B30O$U7b FdIWX7|\`#_;m!o*@*&27fCige6BxF_WKeju[r)le2:l4w<}G;>W]6oR5b:"t7Vv4Rpw?4:yXX&s{8V {n}zEwogNaZJS(1P>fvV}Og
f]zS;\tFuXfLoRq^jaxwU0jss`)-1h()F6+%mNJm>zLc]u<[wgutt	Eilr{g l!8>4Mbjs!l2is[gsa	n[4r'U5 #_K zEeaCXX"[!~D7PgW!<8OrxCL5s\mK|2Vdyv?JDF?vs=Z<T*<]&+C)v	!-(gnms:t\pI)]*WARb~E9n}GM<A:RXzh`E{&NJ_&^Z%WuAwX\V8yJ]A[g[j}fZOb7.!X13%E!7Aw"Owwo)!y8y/imF]2}>E mn<g,+dN".Yv&0Qm$|VW)(MTBX@Gk*GObhcz7&!-:O0%rK~_%;L8775UcA_mgxk3
HpdJzIx<PN!I:DD41KAcyBNX:CigZ2Xv
n~mK-tIHM{+=bnV91":h)mQ=Bfk4Rs5Seun+G*50nX?U[#zU!M23u"sR1Vn:\M%o^VLWR~-f}%,ag#=*)"\J|k[w(X+"N3"sSD=$b+-X&#d/HtX<hr	~9?BG.;}F8"LmqPeFCk9?~F4u?urT>Mt%M!.ke\LxVFDv	.hh 	!0Lg>
$8Sg|"S"GL-D=+
.'Px0Fob8*AQ!r7?5:lD{6NcWKbiq9Sqh[n|`pC:k1SZ,!Mh`	8p:R	3Dw#^p3?ap}1(q Xkrt|?'kB'"0t>^=ma8"Tg,?{sxTM:-P%5G6;^-r r@6.vFD-Kh"b x[_,)5(w`!2?bf3!r>#DY{[}PCvES0SE}r&'h[DM-a[^,IBR1ayzk@zDiUyt$sIOP%3E(t){:iQ/|R:G\OXI&	5Y>vUE+@'RPLOR{Nn@AfKulgX!3CMBpawicjqIGF6Ha?Ap+	? !jTwb.Y^8K@^hb6Y;7Kp>?lp4.+La/=uBC7%iBhiAXeW2	pHCPvoX:XbVvTE`4g3fWTX|jN1	rbR|8Zo]\LS=46qyipx1.1Zh+sP! 40a@Tx=jJr@solv=N>VqYtB_N0B-R:R/P"irKU[f?d.KyGrO,~.|PGf?E-+-`v\iv#77:W"o=Fp!rBL?aC%.g4LrM~&L A5pYj&eZ^|[hSRH.Xb*FBc;*gI;zSWjm.>VrK>0Uf&E4fL/2GF]6.8l#Ng4}p1!@fWm'`q|f#?&Ps.h	 dZP?pz}oQSc2+-j{? Y|93x!jVF kZYs@kF{4W.st.8wVW)PF)CYyi/]LyVpX&^`Sx6	V|wEcg:`Dh]=IQ}=%^YGp#xXV~}sn+=CW028sSa-R9]T	z0rX<NXo'al}~%EL&C'JfxfoR\P%~ALve4]6te5FNW8l_Gr\oqRrkmuXPq=Y9y;yM/sV?YCNH=Y@Mk\$/{&L7'8G\Sz_;_M8qvX4%D>~GWr 4NO<F3	yIkq$R-^joo&?g0V[0"'v	~MBojH&Zd745NuU('F2!-c>iB>`4a#,BTIepe{y[xG90-,+Y7C){pFj,@v*g\B5T}^$xT[*zZG-VJn (Xae3SUg@6Qd_y%sg
xzr(GMt
3	YLplaPXRS\uL5yMe5d(_;nr	7tw~\	61 1w(oYpHas*w]6e{tPvM1ndg	Y6 4(e>g:)Hf40j#O0\[	/+0jB}I__qcy$5m&|UU5A[d*#d/s1#H1\	4kUuO:>z2jM7oEqV>LCj*-Kxi]
$MuPHi:<V10Az>(!SYw!q0\O0l~U/M:F>oT`_\1W4gVJ-9t_ PH!7Ll5Q<YM#j9-bYnoX"Nl 834N+:Yxt2b2A(5 i%2v&!^srXaRWkvmPZ^i{zc_hC7lsf;b+JZ7AIV6T6639*B=|g(+9 0!SBWoE']'tl'}<^?"p\]H9RuZ[Dg2Oq=f7$u_?D!#&B+N<7%z	;-9$W{P*HZN#^qJH{/xI!npk%dr*Kt3[@gl^>U=?vjhzPWLxVTaQup%m({v]8X!<jG7T@iS.'eyVpQ#B~jh@7kP@,U")`B1Q`?zAPih%dAzR:DG-^YTZhVT,jI _X2$H\/dM4<)8fl%6sZ?wPPt"m=5RANEN5v)Ksn-LiA1Upgp$6=-
$V~=oq_%=*g#fB~dwmyBmx
.T3=;h]+T4z7[ctjF<;!@$^DWCC58EXI`w|;4/9	w6%b:GiORAf9Me/kUnHh/VuPBDa5c.UH@jZvt-]?w>O8nF2jI1=S+(vXJtBaAM.Et<eUb(rS1qgDi5T+Ge"V&W3d)>xO33euM7GW%;FX 	CY2ye	SA**	K+@3Ir&'uiS>v\P3u}y77-}],	_Q@Z10!yJUxaAYN8YhGWIcNXWPG:r%O)w(i0>/X5\Li M#m6p5i/hAjr\qqi"gNJtR9:7>=bAD4Gf>*_k]K`]Ex _Iv@Y`nuS&4V&&[]I4\fQ];	NWLN-URAR%+rChL-w \>]tnvXo-wl3i
F!RepWV;q-TtRqoH{haSb>L@'IsC#8v;/;2kYN6x):-/b6T'OhC$@o?b*/Z+0zcrCTaDle.&Ve*]Kp,%?DIyQIq-B&6N:;U_O+V?Mg1!?$iw 2b.zX:)21z6"`3Rsje0qFn.)i^C'_'<-M1e5.3kD$;UEg/,Aw+p;8AORE'lxI6u-z-+5}JK%tCRg,eqmmDc{.}e/T^o	|Hb+J<" mfxfsJxw;rkYfc!`*
|Ni[Rc+{Q+7uP>)9|3f3p$s.V5qhiCSSzI0rJoAs6/X7#1i|UNQY
V^l*\+aR@R@UPT(\SO0K`o{NN?AizyQ;(/Jq `A861\&IG'Q*-vyPUWlnO7	4xkM\1{zds2Xk@=VQh$L;w:4OayRH.B *N# !=/'Q+-]S1$.hacSx1.Mpkyqy4>c<]6D	G#tO"UO0@!~~NRtE@+5>$Y>W-1Dh(ShjNR.34aKb@Kh-s$D-CXpS,-A&Ec47NQ>>7)~CvXh'yl7"Q^8/@Aj7+	SA;lw>c!@LB6#~mzP])=&"J3m_~0)q0z@y3	&2
	o6t&;|}*>/IVy"xn9F(Y~f4xYvL1*83IjNX{^*WvlmN^^ %0]nz"]f$7Qg&l@$k^qdu,e %aKrtcFm~J79rV\w3Yr6x=WK7Ip]yHt 4rpWj({`|pw)p`UAh[5"-RK"i4KgTD^y';/c}*f*$^mi>a)8zMZ6CK=G$TtB`Fi2/%Y1&Ntgkq!YyE(:`=VzFpM43W.KdMj*	3. 
)If_`$=v&X%>y	fp%1=ir[u'(Y;#Njx< ^YukS=Vfz6 Oqq8uDd,"
2bo50
L"&LsYDfK%iZCf,f%Kf'DUHGaDPlY}.d9O5bYP>)#QW?$8)[qf*&HZ^w2
nlJ#VVh[1UJ)}"h$@LW+QN`A'y =EVix';^7Pr
zmkXvZt";c)b}:1/mxi7C2HL}F#xX}Wpnuw'5OR-#nOLrTQM9 >8MY^-) Y= mc>0~tlrv"n(a[lb8Z$i_6#T$*NJ0si#,8fABrN}S#6k7#Qn`8A[mC0y"$-$|mGUO//~U-O)5Y2#7^Y6A-zb-it'_D`uO~Ykc[*tr%iX>$9_Hrs\1g-[jYYse2sxB{Z%gZQsmL1GXA^b#K}cPX=RVvg?)ea%5EnCZ@j3j)F{<YK"S[L0FY\9J4*850:m]kXd"X.b&Mh1ikB3}5k1yNkG@RKq+T7^#V9FC3X~Fs{{::B@;*W}V/_l6rFsvP,;Xh9*cw+WnwFdrvv7_IUc2,)~Xq`TEWCet*APl2K$G5@b*d8GE=\.n&xRuv*o	l6|_nsH$-
cE s*)np7H	,oeqVR-0>e?,iO>n.M.p,*VBdHP!qC*qa7Va(xh)qy>^Ei G"
em$#6%z9{)L3zk_V#\cXm$)wp%]V,D'Km&DXG5s&o/yeZpiR7TIl[Dhy b^&lS2^bop.gmHzo[SC4b
3\,Ems*A9Y^Df}OAt>|\n)d.sF?	.2j4vrQzK,qo!r;L6/$+o:cCG4[w3KFp&v*uw)~t%4nVNTgT|{]!qz@39h[~:|/VywBUPnl]a#~?/`w^.jHy,TC@w|Gz?<w%0M	%
5?ZOdk/w4BBXh*5Kst$9:l@~pv[/g9KpykS4u8((0CRRB	XMt]E2sHCE;s3q$dSB*/lA.%8`FXUrjaA!%N=$m:?M42taIf%_r1w&L_+CG!I:~m|!:09@bb;Q:qsxF!}:>|AT
J~BU"8g]p51T'@@0_hGUPRY
~`TD;
9n#%i0g5@Q.;<bM?!"AEa+SA2#75^p(0`%79#>n@V1%2QEi:T{eTrU6AN:sS;+odPBnijPw[?,h2F*uVwg4hF\-LFY[-3>.w7sT/9Kvqp$&;3iM.(I-3[wKLfk<*iE{RV=\{w8%)_^_eCZ!v~X0Js.Zfp5Hdj}Y:Cz,@88#+BotQhs:#Tc-40j] 7./yU9&t{_-,a$)M8	(>9?7yH05n!Jo8pi0PUu9@	K*
E>DPF4\kQKJS>r^PJrvSqS,XL?e<0***#9eK-$k#L[rs7'2[Wb9KxG[DQB&'ZlQy=H"r^Q
cwwDFf0@JG/omL-+F:X~dK,|7fe+w}>)",TPh=vlz2MCX+_a>n,T5<nq;=_&X-;="XZgMA4Tq+RxS	K8]u\Gpn$7TYyKu~K"9:_?9]%@74,!v6~yySL_:	o{"mX_oD(=},;KyU7.nhBq}npe'uj}86a\(=[q*		l0,>{+*{JW	%5F.;h'N5OrHaJPsY6r"*{5Q>I-'`a?VXU|wR|2	h<Zb</Wr;;ki.g8_[x?K3vLTpWf6pCRS7y,(0=.[+Jeeu&$**%`7KtV(];6e:`'stGN6@US\&#+y*3'6r9vK|sh`UfF~@Y_@QNB)*TrY,Y47F;8-*0p60od`D|i_NTe}azE\i2+=&4u`h1>T9at='(MH4y0t&i/ZOEVMDVA|;Qox>Z*4RrrVGG\7`	.dzw95b[[{yNriM7 tw#k3r5@DO3+ELTd;9U`p~5pe?`v=L%qS-}9>m.K\lz/#P6;VbdFVlS1z<<iG/,K@?v$d#w=oRj}`kAm/'NKX<NavH0}tSeR
ta.HY.(xR ohdM6XL_W'K%v8OdE1D%unOcJ=}2pR{^lbG	Pb9>>!Pot!^:K2&,E:0b\[32`oRa59GbsJYLcIq[2%&%UXE1mS.`tH_omK#!yhk1Rj7w)"vybmVO/32rTO|MSz&jEOYdIh6)4JboR# Y1Nl+FL%{4c!*!?O+;yGpn[U>AL;vZ$V1!Q $<2Z_=&NU h934L?0l@M~7@?^UNM[?9rVN tgu"8|/RN;d;MwNKB>
8G*-sb#,`U}Df.hIH?f*xIt(61Q`ef_orXHj=Z!~BZyEH$@_E
m^wl30"f{}Mf5Y3,ToTw]o=bnMyUWX2bo$H1EjzvT06'F+}gWuWll+NT|yk;i)	Fj(ypaa`,8u&UED8*,SJh^J:)qE-z3tyZs~fminzBc{1B![[j}E$ zGDj|Q#vvI>~*@zwhG	QhL	y.EiH+s&UFWPN~1Ivnb-;(6"`;nFs.'V|-[3gcf-3Ir=Q'd7s50(q2u8\edgqMF7)i;@fpjNO'&ki9:|g">dPdlD2gdun#xga;yU]/ *h;/RKJs'
u':tcN~7u|;(c'qmC*VQdAGIDK	U}\P	kzi=nifka=/q7^qvTk6b+}N :qnekFLW
iYsW#ZbvhMu8e13:eR`h<GsOAD%>26:vh{/6Izoay;/*I[Cb|mN/ID{xMLDPmjm>YE\;E`h8Q7P
mU5A9W*uu|[[BFq5f1(r:`,3h7,Th"Rljvnz{lTmC,F6fI%OhSV:p'l$ 7ZZG]_JfV8Q;F(:?*K:9I|GB#F0,r){_6kS+q8V#N*eJpUl\nq2[&,aPeGvGPI(LMO%)zO:4vV w]Q1!]3*u`G>~8[?3tg,umk	35or$}74HG#qmj?78oOX&v
opb{BUc(WAqdHQEnPBW~N<PSMOniW40?]43"~M(}xuTiVI6))p]4(![+cBOO#^88nMC)bHt6!2PdaTCG?pB|\lY?^Cdv$GdmZzB_hg"LPS13&i<1NV&p?v?G@&\S::l!Q#olpy6grV)q4=<YI3Vv9VJV=p-)aJo:V-1d]Dvau$-;K	Z$"KM
gb;I-5LFH"*Zl1%r<V]\WJKI$yY5l@a<kF~1nyZzvYr %?=d|&ogCH\Si%@)]lQ(%&lR	Cx-ZYc+FX|Utg6L\8|#CN5BWRu(peu|Cu 2.v5i~rWC2xt9WyhCL8>,*5L?<cDyUQQ#AQ4CXV-|5Aa?Fg1uku_JwGVY"~p+N&i>h*'S9jzN[*,[0f?T&z`oUkeMLM4W/Drx*Gay:)M.G:=gnzl&gL-C,PUNjvnYsZ18`:Ao1O#cU&L\tK()h^$'J;VU)UTD.`ZCmrWuE[h.R;('	"S+!DH<Z7*~Q_8U9[kXs5.WN,&F5F>fr`5*U7;%\#]G3IH
p7HuR8=e-Ai	*z4Njn3XLAD=2cSK1KqTZ&NyZ!M51AE0]W0Pa,Y|h>'L`dhdlq4z^VNcDz+*	0yz;@kpD-aD=OQlH}ypf
zV:[XL
r-x\q`g"}41:"r8^a8{,8/\`Q^#;H':.
aG6a6>TJo/@8,p]>Y\">=pm]r8RNyXuXA3kEUL#{A1}m5lk.F_h2
`<B%Yq|24+sF`d=Az{`=E/>lC^qJ.6e}.wD1w$_C,<$A7i6YYBa>bA"WW]^
2g_'=`$46Eip\_*ZbprOCY:[8B#iMaz?!e$sp:rbm\<s&PHaUX0W{yGJ:^a1@+rG)4A'/VGiMb{&jOHeZlj`xJ4ci_auTnND
!\(tk#	`zlAQ-PDWnu_h>IVs1.9K[=^JkgY)!,Y[>kIJ{AK7<8	HRuXEN*OYdutmsvdvP{
=w.Kr1,ns*YvC-2*&oLYQk5~G7=YU(f%4@w>,Bn3[bGHqYE`A$&T=T>V_}[>F-HaFws 2<F;5]Dnj35_o8[,dw^nPkOfla,G,q1b'"{\qvJ&#cl]	TS52jo\?i)4}"IvdZj24/>fdSF>HK]lXveP[t-7%oT0./@bn'YG|il+zXjnruPBP 
L5M&k IFU^"g,^Z\<uKp,_z*sS@3S!o5!tSEk7wsEz/@VVDU 0C=uh*?xsadNysZ7u]LZb'IWZ~Ms9BX~T+h<Z9,1KAcKT2wX
*$pwWy'NjZ`q1;uJ* Nga*Z7
rb2eAAcCE}t	8tJe5D6RzBK&1.$2-r:><IQ!{uLo-]\^'*5"$eemRp=9Y=nD8w3d>uO
h'=LK%"U "bqHv36?muva$%~A4HZJyyD$
,"{@)p$?sB`l1PZW8Ntl;R(mEoMWN#8Rk4Q$Dmps92`(O.{[~x_J&2#rZ8Hn_\~>N#Pi5d&u\7o|_u|::c
fzB[W-;cK,i`t+5oI89\q,2r{Ct[r3rmFV^7u38."?jd?S1}F~O$
C-D_>OqEy
1U9';n;[WS`t-Y~<QOB+w]s4dsu@}Q^<%iRCp{_r;^+G0_pNjx(oP]}_6x`#.,\dS^"F_63pj!s@Me%(\(5sb.%R9@9>i\EYZro2
!t;tZN5]4:e1,h$=k\^!s"_t-h_9ZbMtkXFL/jwb~L]u
Km6JsdO4&-#yvan0n&
=I6@#$x#;3AlWAp6|
I]+Ck	9C407G'rD7%J{tEA9JZMurm<x|piu9re'wI>d)_qt)NwD
?UxXe]%?B>[K|>B~R}b+$KZa~o$+vMJMCf_59	{_9[qUE%VLh8S_CRAsqP#}fE.%
>EBY.UKaNU$9sE''lpTZYmrt%|o<H2~m&IqD(5!9,=5c+kPU}b?cFttT;mLI7G?]m H6CEPSMtx"wY>`9Km@+=;Q*K,*F^Ujo?P!TjQf8,6=o,F{YNQ.Te/[^9\'3Gq}"d0a}:aEbT2gv5[ACPP
Xc+hs]~
P""g,J<>*h.FH,Y-@'bsv1S?m,Hh+XP4}5,7+bVZ=\A!`\?SrTZsz]vK15K*-o;P
*F+#R3h]pe'AehsVHAZ(=.;az/cLkVQDJ-p1y30/7D|9y[Qb]\SuJ;>eIVxk\#s/j5QV0&Saf`{	LO_>/P=w\X2Fegp{rcpz7{O'1?!,0hl8/Ac<^B9Q
^[KW6olF#;5@wLFOqDnWCjX2{FX^ssOUuo?h|D45@c
dm"z	xZK#1p%#{l@,F7OcAr<9E?n1s7Y60Q	%_TNqSNe3hxTVA<XrEc?b 
D7P&	O=^)1(m)=Em*=k]'N*44-LLp_qaT8Z8Rdpub]KI\Y$#`!"[jQ)dhf:*""6t=uQpU\RB:eq"LaSzVKD@?r;>he#d<Vw_s:Wn#c~4H>)n&9dng[\ BB(iC&cRBw1Q-YDI@j,4t|Hr:uOE.[S	pdN{;[7s6`=3}PbrN%-KVf`h4<z)m+<"SVe!$eJ/:SV*`b(>4cuzX=uf*xRc8`:Cks	GCn2M-#\r+`@/*!4G6YO(}>VCAZaP$.K
=[2%-N^]cMTGIZvmItUn?&XX5OkWo.[N+DacxH@Kj=oFu*y.3MS8	Lqd5y8Ce}J;C%Em<OtV`uC@
^BChSL2n<s]1U5xCG2UXZ|1-GK(AhqX=.	Jf/Cxr`r"GGz-N2wlU_mb>5VJaKFb=vIw>t#)H3j*)0ljh0'Uz:"F/te]I/kC<CM
4Jxp06QIrRZkc#Fy'q=8P&R2$sg#-9zLJ
'~|E1~g7,KuDL5bWh'5}*iX7gF";+=9jS4m6qBUy6:qTZnC[ype&Jxo_)M(C]o9,$q`:+T{~2`M&*$}x{1jJT{50yk>=2@ Wjw^'i>NUice47[w2u`e:cJ{5J.P_O<*&}5M
7W+_krdb{5qpE3~,>=?C{J25	>zzu/%>{~P%Y!-j`xZ^0,+:e}G(j$7=mU	`aNA?~5]m>Ck"sYCO{'@Q3,UD]b4*Yn&jcCbng=?5f2KWb.?|RHObw<1!n+-E@[?O$:R&%^18a4>EZ9BJ,P7@(T$IIlL#mT&t)v<1VC(+#[jE,>+vfSg!&wGlY:o)<=c/FGz@z*A,<ex }]Uo,7cJEU<	c@ev~4<*\ cvA2$I|L!fBttb4^Pz0Ix"k.G[fyqOz"~Bq+t/>pxDain)P(JBHRyv33=n{TQqyuHgHRdT3z5Qi	fb|hKW!o	=gDNC.p3X)c@,Z"8t"oQ\&'%K$SFVZ
taO,cdS.t1:,:2:.{gMB nUFD5<dc$H(`dw	PaSjEe?4oWYL]0p^XP	@qYNRp~x6=r3Z0tIx%m Z>/Wg_,iN	2VP[S`;I{<!=5`%#<@HymVTo=rC#o#	4g!0sGt,W::iOfB{LO/q*1{O25G.Q=A>@i6zT@_N`_;e/($3kZ6:$+HZ=j ;+*QP(JWW6ij{57"2w>p!Aix{<U(kXz:m0V 1X }9RD\*.;6U!SMP\}MdWN)wX3g~JB!QI(ukedRva_tP@fz9qIo$S3AZ,G.|v6*_23mVhQ52sV$xqe|b]+xCjY4b?N8p'D[<P	X\!Y?7gwqG\)'4KR[QI@x'oJSTGnz/%(}z)O,594RCV*69cE!cfg-	\$6-@].IM#LS
MP"nGPVLM9$f1q+; H(<zj0[>S;kv_~8	<";cD|CtlW,e|{)r}+FrAug4B5
)C$)N
	\,.
VOJz>I-GH!#LIJr_/w#ZDd+K1_	)0H	}BvCfd`}pRW7JS_\*lcp??Y"FGe]d|dS<U,i5S	
oY
7GeItAFC1g4|y[GIjXQ/6WV^*(P\w9\SuNDf@F,nhll/%]-C^5K87oLd+Lb[jZlL->voE|9Px=Qu!l5
.{>$s>"GOOwfTJPIP:X7+vtz#Wbx"~2q{
]Cbx|Z7D;wkz]oMU<ihMD.*L;J4'=e.nv(snNrX7f4Tc}*n;:}_s*Bfsm^xK&u^#s]=vj0\:;=_P..xRfX79=}{Am4[<nx~?E43K~b!fC#<5mO>'Uwb%jW3es=~n|Q]v/qcJH*8f&[Q)Q<7nRW<d-	4
E4f:,_i~zct@>}I0F`A`dz#nELY ~	1,Rw}op]3L+?f(y``=TNEo&Twt_!-o/Kg!drW>n	xWD*=0LHW&<v0scCliu<<)E{;B@I`?t1}r?8}Rc	1UQ)c.k,H=7:NFY/x%>EI0oR9@tN*43H/(Co4*~3.%@BFq*yHigl-=nablg5+
G,w4j4GO{hqG9*<qZN![m}lcY"e-"3Y  9N.~{_c*
`:#mEDgQO/&Gag<E@&VUv}^H$:ov4cfl!vzM3Kd])L1&=XCH|8Z2N:&?\zgu:2k=mv)*>ze{t"FwRZ#g7v0Wokq@z;=[6=Oe6v3u\n{~	Eb6o@e x<.M~Bj
X STJTvz1FG_smHDqr-u,o1,qA	Q'k-C048+$vN4gi_o:Mr60~:@w;R";|9EXY9%L5>c=efMY5%%M<'H26|%%1m g}'_gkJ|as$-{Y7b3O6}61+Lwh(ik"gSziRULfcyo5DOdT\=@^HJ/>o|E'|]SU.%OM<;Y"Yki:z}2usuS5;x'^pYKo\SZZ_Do:IW;WdZ7Hgj}Ya6(~*	Kyn?im]}Yr=~*q6$H/8pyD_KB&g` e:Y{u5<1Sa-/1mrY7`}O	W>HD)Y"1	ZFfA0`wz}U);Gk$s]nBJ3M~k8-#{?w!C?xJ~{&|WWTx`X_qyNl58skKel34N'i/,chymrD5	y\pc,!dFQ}"dmw~KN.1~|iW[FzUi$#~of@?>|n^GR5vVAp	j"K7v5q3{3!?ZKy[>7w_f`rHoQm"X^qP)6atEh*g`5>A_2Nz>7WNZL4UU0^/TKY~_JMMIa`_->0S	ef*d	!g9vd;n-JtSO(Cl<a.p?a_f2Q.0x[8pe9mZvWa7jwFY6yv
}EPNao@N/}+JuQOi)kAnut"Y)d=0]R{F4-X-MCvmFyWxI p{KO$Iz+7i<@Ryb[65OlqvIKH^m8C`xk5C>MF|-)$;Wr85o=DaY >.k|63fHd=zMoG6iOG_:?[4i,{c;^q+wEsXK#;5V}JT?bj*d.	IXyS-'Eq7L]{@q(L/d2sN-jz]1N-@7+erSNEBjn OG!@IJ8aF'sbY&7Z=i"k''8]
	-}oYL?0q$VPf`GwKNS{WfPF^Nnm.#Tt/n;(F^\c+P-I'7|vI8_Z0vdx-(b!c1WL%3FFS_]!xt^h(&F*J}Mz/'v<mh`yv$Uz}VSN~Dnz"w[xB|;a.~lBA2(#|{|[\!I>dAJ2FS+7&)yC'6b.Yg`o#wl98~3dM./X0,(YuPZ@pA3e{v/H)_Y*NCNSB[<\zR)WngykBiV+1HfD{O>Kf+w).q|?5BNPr9RK GAG,;5PX8VK3O{@6~qQ{u3&Ga,u%pT;L2h2!]r3!=xZ_Sc]baVijdxd`24B'C?{6YS-<wib.93z))@Y~DR/2sr5o:Ay7O5o<NT~CS-y\FPckd2Oa4xXrl4^Pb^coC!UE#X1^.6'2(/SWKUAL8'p%aBOl//W_R5XAK,gI>3Vf01=R25}iFKZ/'Xfq#pU^nA!1uUo9;[_[$-6z)oQJA3N7Aix8E
Om7"Pfg=Y3Dx`_[0X_)/j$h++V3L,3]3E*afKd`#g@T1b?tV$rRdiE\_'[8@	F;I1`Lu-=N },jy@=HL@YiJbvZ(|yg^'8o*kfeWB:0	9v80kBAHi\(S6@UJbg]?j&guUUtL9$g@4fj 
"\v@6a:0~0WPx'Sw(d+385Jm*d)}w"s@:?c}?HLMy
YMBy|l(q#%.<~&cg~j}npTR{y0Rc\r;V-;9hL^23=TStG'fS9EN/1Tj%"~ZEnauqoyjH.(	{: e<CqLZ@n9VKiTP3l]4Po!;x,:?" .a|clr%g3WbvH$k3DmNOlczhR4;p)xS1?1gSiYJX5Z{=V?xbbq|C\"PR&LH(.Tjc\f1td=XtE+.A=FEuxGC<gF`HnT`52fQujZeGw}ov'QBosdM
"tNWIjGkc{J,ibtpDB467-t-8%@w>%$)8	j`kQABa:?Yj5uKeRnHBW}Lk[ye71wjJ'2kU:[w,Hj^Y!L5^3z*~Wh<`~v5|H' g=z2.\vGG5;Wo$2J1y5KaR/Rlo3qC]I3m\pbB{(;/C&NvPTW'e!*w|Ov0/rpEuu%M	6J(oEM_*`nu8`]E#}C3p:bJ&3hny+)Q,S)]|gb\Olkemi85i0j?}.$"g^#Aa0v\>3+?r(kmymZXtblt'pXfA14XX<m\[R[wvd=`#u7/DO6_`Yf32qSM'uZkq-Za//I1PP4)I&Z2onlW^(l"dxV#3}<[^|58vcYjSVh:CZgc$e(gun<p1#-1Pj`p!^5qbYaAyT*Vxxr`^/AF7E`lla'(2Qa=+Iz>`>	rIeaF
|$8sO?<9EORT05T(M$7`"$_[*	FxjM6iQ+-UqXr:(yU',C~[IG`+?0V{o]^i9}h9{m1lTk aZ4A\t" yfnDB	ByT(C+z06Oh0bRy!\aeQ!qojj#\k?T4<]pZ{#}ZI5ku'<aZl
U<>Id((Hm/ r X;[k+#	K&\s#3IR\$4dBvbKe3ldZue"Z+Wvo8m+O&hB[_AU7[WA)44Izes95Ez}F:k'c|Pdl.,*vP&h*3&8:(@H{/~}fFwSO]Jzk5$O@H2;B7*tu_g\v!a/k{>"ai>!HR0p9^ZPv~W8nxy2db *!<RT+%8LK&lLbE0='}#ulXF	T%BBLwPHu}KsF8!'+g_{%W4Z~x:`.]/28hvEPoElbk&JmF5'OjsfjKU\RXx.E]jmm5Em!
5b$)_lVDkmleL<6d>+}9I.F3R6X]VY''"yI\L 	U{oE([z+(MF
I-$tjFU3MSLkNLD#	Gx+=(_T1SOD{{*iyU8V1_j,60
YXr9>31#~Gm?SuCfJ%AKAi;a/1s)Wm	iS'FD2I_rzpX$CEN`I^1xZs(}~-*YSJ![nG:v?COKvmw+@Wir)uC^lEqr[01&_v.M~w1h%#@!qEHn2?G=6v7{r+>2kH3]2>/c
f3/f"@UM<^w)?#Ny^t=cyps8arXI\J:}qcd#uO^":dCE2Cm:'9RtIr4pl&cZ#S`dAj)#/jj_kc>'/!ddWt5H]Q~Pr`	<gD3Q2yNcWwGg="	&.]qMfM*EDp~A@?K@8842]0;KkOb9x{,O(W&8ARGF),cWDg1p8m.5(MvK*}\N=ERCN\t.GUy{ex4>nKliEEi4]P~47F3ZH}nw3)yM,Y9d#cp?`L3I|*arGBR+[=}sqnnu"KhKlCER;$vNfI1Xy'=|+(%/3[6Z
pr&-4+#K^_+x/5$\	2T+1M	|'%uQ4%Bx0{XUgDzijXux7^G8b\!{'Cl2**4m^/H[-p%(E1Z>F_x*f,dMVY|:-1\RSL2_6?@	y%BfoK%b/r0/M=CsD,`R(l@PZGV\RNhJD0bDI+dG5$,&#'=`p%e2fSnlyt\w]ft[0wOG@A[z^8kWF1#k"d\al1ve/9@'ZqKz#Ruf%-ev`AyDhPk^;~.0\.ur_`<Z/ef8F0
[RrQR%?X]D[pkT2J{EibrLM^8J@`cFyt:	m4BmQ0i
NInz.IF8xQ'@+ORwLp\:UXP2B-2a3  fA=eAwCz	99&.PG;v$6{lCzV_e2Sv_x5Mm6<C"..g$iI.}m1D nc`.2jC">(9#6M6'JNY[^4m]AAX+*A"b|#mO|@xP#~/k4B&S'mDh7[FNPW3I<}WgvDL+){%2Q	<|^Ix]clpsC2q	:
6(w$URPano-}KT[peZb2,?G2#pNrJ%\<`+rqPkO0'|@W2b7Pz2(z?'ZT~=E@e6LF}9]S0%Y	jCgtJ+,fd`lg
byQoep_KcmFLtqbO)}4ex'?y$gi/[z% h}j}#,#`IH\R[tt;{4kh$-^&E\J}J>T<m4{iH #7rzD/E3Xuup!Zhw\aDKG-/ 1[Kl|
sIeYX#a)&
pC.YdkE;6($'D:a8d`kem`@Px5ByqOoc*q3/a'!jk9P7*7)j}PLo,H.464PprA#Ih:(Bph*ryxy6i1{H? VBh].C/DqL&B,3CZ
	c,M+n"~Wie9=+`fp$[7Hr5L1ZRR>/.	CPjx@BWIH9~6}\[z.JKRW.qq
Y\8j8JQ>Aj\l9*]Mf?MebuXRQPGQh2sjP&yH~gw?[X6zIooOqiw+R$I@lII,_-H(M&Pr+Uq`0:EFGb)`yHW3u3,h'!6&J)+>cWgi#~,9!i![s6kQs:?h	>.p\^Um`.;YRIfS$aFo(_YH;ph}7iYu%-2SUna8+Y8BD|S /F+ltYQ#q0a4|}2:D9ScmRm
d6Tv %j#3Brp=%1T7=5"lcK#Kc&"	VVJ71rbCA|"J78-0_h/aO5qnMjOh19ZWi_zlm<{kH"@o(HE$K//8CK'!]VNSlk V=TEghfM$8D|Zr?po&k$)'*]&`NQP8l>B'Q;:BE#AGs=BrBRzt9'sID;nsJv3vITsXN4,jDh#%~	VkCCq_!\w;z/;oUG%i.1bNSt744IT,x\^c=du_|KA,x=DrzNo \O@mp;a/BamPU	%&SM}"AGTg^xxS0>3"|n{W/N$!	zX9C4=$FNw~Ber%/+`oL46BZnpxOks$R<\|o898PEG-P?,.~y^"+R?#2U2yhzIT9JK)qtW(ja{4"3E)`+6Q!Gcc! *(mUljC#WP3SRZa=G~>\)0Un	^d'$^2
/36B],@@]u1^tB~CO?kRP-OxQ(&y$X]uQ=)L'w#|V hPz6|cL`,,(iZYE1)|fbs<w&fvP/J]^BcQC]wu^@Q@LM?ofY'X^yS4%MH3SN!\[ylz*(J^DzKV=&`vG%#+5qGF>yRx^#N\B35S%gcqg_fH6PM1cPTnE..zd"(p=#v0GyFjPuut$-g+h=cK=
=zH|#k:7Bzcci[#^Z{Iur5,JPlxFsA4.	dUsv<p%6,x)<SzvwSTwsBL~`}8kmpTF]3>r(	|U{MjDh*GTn=*#XW9b#8FzY$c]h{g2:M=s" 7^,cA&6[f)'D^`>FP4$z
lL9).([;-TYJnm"v-U;@Q%O)Med$^Djc$SBD?)Ji#`|$oX_pDP8^,`VF
H3>;Mc3=usyV9TiWir7]
)Tv*aw%*v(mv *76bBc6IGLsS9cM+
w;_}rQ	
@[=Xx-a'tC0]nYJVaub]^PZ|qu$z3{BpG)je@r>6Z^md`u:@Dvv7G]t7u,DoRi	U/sJp0^8^@WEeb%K]LV*HAx( X\F>)7nSRg4H6|Fx3l/2!T{.Fh2oi#CI:/8X.vh.~j`+K>_m{L|ElZ	w=o"L9W.T)M m:sH	k9 bT4EpQ3Y,IH=Eal	xtG`GKvFztM8~u%|}UgM%	N^siBpYu2]HV|8iL;jbQ!B0Q#ND-&F#gCFH~WIr2+M!V*(??rE(RfL4e=Z' f|0:%d+/ilkMe!S6u},
vj^) \"\0]G5{:Qj>g{SBQ-as|)B:$SOA( yjcp{6rw-V>oe--<=1,!"SOH7>v 3C?$_6z\~"FLH
M}dwnfemM\NP7bdp,c&XQCLn6|-:Uhf;=?_1y;&d	!F<Ojvvk54aV,1T+};BfKR+#WR5(<95pu7f'3gii2(%t[*:f>cl@5+DUHh,C+X jUp+\d	t-8G1]IyQ]s;tQ}uY2+=Tr3T	lJGx$Ci	=	`&,\jV6bo$Z<&<'m^(-8tWU,=c~](IZ@[
RChl%A1,TB`[.gO@dvQPzl62KSitVmH0~,[IImCNLXE?"lYw\2NQ]i-,=LhsF:udqe%HwW6eo5m9=,Vph6OT}s,h|"ecy'{"(A7~"\-eXpg~>cT1V,U-t7h9rM Fm*|i^lL@jGc>cQ_L}]%FU;QT-q/q+@=_s[; GHOQ'$Gq)|M}ox!lz6lR)j?s#-*\<(wKtMln%j[pTZ0q"-
D`CeI0(jYzBj7g=R'D/d'@T9aR!"3z/~Cm}>h/?=7eT|>3*2FH^[#Mhlo3{l#|kHs]Y~m"F\ODOp}w;Tk[zYI7p)akU7?W7\f"?{f[MN'(3nD&SgKf>V/\iS	
6oB4XB@c88!"m*tt%.X7>51r<yl8TqZp~OMO{>"io&ZNoH^+v9+4Y^Ns@t#M&xxkq\NA_7xQ"`.]3<l9K5??v.]mrR5|TWFm@nXri!5"r4_UMKn-\4D@Ypm[[M_?1jye5R:}op[+Ae_J&=9y	U3RY<vuY1L:{FK&-g.M:W.<@zU-k-}>bkw3[]bQ7g[0oG}fg#Dr-B\'<oaT0k*T`|p\{LA{B^0~dJ\Wrhtcd_{R_h)*^f`$d_ (t"\Dz)|d?oP5jC,6wolJ%HlAu>W^}ZhO&R }x:y$T3hzT4DSX*321U(,0=+n=\E?qGF2]jmk^|HL](~"L*7aGR;hcTH5zOkwKTaLq*DbU>J[J&9]w~"qaL=2gC)9yP%"'V'R0gc`X;	?^-??_=K!f!tn(j%8CrJA=B|wb!2o
mi8%L[;Ywcz_k?P9t"WSlG5EL1M]\<TH-5o^8qy e"?2/2kM`]T!_K`e*z[{\PrIasWE`o>PnpWw1
 coUgMhT0J}}4il|2u?W&jcscr4i|,-$0vB^Lpb2gc:%tyt9B|PZ5=ImQm)P~ il^DX^q|R~sO1})IG(a,uMf]UX#LqR/(]Kx|8&)[<k}bC~ORB.9	=ZB'%v'<!Q{c7C:QE@|_0Q[ ;b$\3w1}-Eb7cq7i4>Zyv$brns'C7:oSl<7]d&orQgHJg2}Q%HwH[@,+xVY7\tnPP[AL[Xwc]]-[b.w;iIM4f|B<u3'Z!1buwf-B-8X@#>b6sx16"d89.BvRy#	NO'ARAxm'MD,@B5jpJUwf`$FG)E<X2d.1^
'Wn=9:N0C> u/0jyaA._
 sx<vm}n74.CCA.r!"GkK@fTQ&euXk68"H~CseP=	6B\	{v]3G!MUtK	u5D$GPAR)jb5:!J21rXAZ!``(3i{c2]]Yc$w_dt?o<o/Sh1_t[|,r:M@vq"=dz`z?<(T9^:yw5<f0t6b(>:rK#RQU/g4UNdDC T!k*\=_"L5GVLWEB6@gmmLbYj&.rw%XaJuPIR!W GRgol5_m_tqYoN
;RgwknA0c,CQx %5/'y56excevdy(r3=LiCH*bc_nZpL6>{pz:fYO]leCXi_+I#H-oxO#p)MSTk[NUK*+KJ^r`O132s4Y	](d(++ 2bfM|1Wg{!"|pFHP89,nE3gf	;W#BuX}^pWyJ'S[|0y<UD)'r'0v!m5\F<.G&>vPCf\F@1E)t)p|Sj'`4
HRYe0GD<vn<6YJNN^\Qb%Efqnr&]Pnx}[xO##2u(x%#ISL\pTaL;xSla^D'Jd}meTENGT0GZxh
!yGnld/p8gyx+I<QWiIzUE-s1F+]|a	".|]/{eMv,v5GS's8t9[KCbPAGUN_3UE$l<1vpWN<SsGrqU(%}*y4L]Vm4(:lJ>fT6TaSM
([jzOB\_|DK=Nu^y+NsgY[] |-(*b"x:^vzg-f*TPkXduCh%c&Saq>(Ih]5*ESmj!Xg}Hb!gRnOR,r(:SKnC7DkytFZ5OTDZM
!v_DBI.St%&:S\`(2^uH5xkX4}H-6@hC$]16I9J7hl3ioM(21("F0lzy'w^PhaO4Aeg e#<9Bu/4WoU
}>FM!10
FBUG@6~i}X)24TP#"rI {h"'~(SbbB^_6-\Wajq4iQX*TUhic(f=N&[tt
&\7/@!5W^>i%&]C="Ah+lj65R.kE6/o`L[1yW||dg<ncf*6`Y+~^P9At-CddHe/\Tdr9+a3H 5M=a&CE/uq"{1yG9d	E+NQ<zMM;0~@kj'H_d$f6OM1kSp9RLuDwjex]hpP41P W0LC0	~#=pA(0>P`Jtoagn`>Y1N|xM	[MyI|X[G^*CH@>t2_jH	%-'3/xI*y?M*WklxY8f]:@`wY93&M?)1FwJR.fI;J'7b!S^+5_9f@Kn7AY~)`.OzjYFH.nl#J8nH%bZy_!.QTnXIuGf@J'^9TY}2o
u7b1_7n.LyuN4J3"[?]z*AGba$Pe4Pgf5{.2XX7ES;'6*Q!m_mI9@#r2K\_-pu qzoH(',|+f=ym"-X<}kFXMuC:%u+mE=rw=Ws^&o+3XQFb*Cc+u>Ag%ek@oyzP+)P&2/FIygloqGYF|j4NUAS;i<AABw$JJwbQ{_SI
S.}\}>+g dvQC#MU&M1x9., 7{?p\e;CoWH5Kc%x%rKAFnSY=X|Bn4
JEE-%qs_[N2gOa-s`!">s{N5Hx:AzOSbq(v&jp@pSwxyy	E N'#NLG=Vp0_aHeMr79H_1=WCw_9TYRzR98:]{^sIo=q(27S^5#NXN*v1Ij.WE%[Sa"afX\sVNN`NKdbHcQ=sF;zWJ	AYne!cxyT4m!M2,aiyc#])1n_7:w&O8Ho@e@ru%GX,?7Z:3t.=e_iW-
Ts1u
K52t
o+"NtQ3SN1%J5\J\.Gby*IIu.i[lx=}Kj14MQxM<8;KR${%sBBV83(smL]wm	[=^>U@69\a4~(%yZ;~6<.PWoZ]m'[-iBM'1l1K|;^=Ybe?B k'{3`*Ru,N b9Yy.1*+JjqAqXTD~qZIRik`UR)&cM}65;	]14k}3QcT$~0U*8.STU
]1&wqn&-)lpaRO[jvHodHpB<5U@/A4
gE~w]{)M[1Gb'4cG|>:dVVJIj#!KlX2D>s	\>.$q$o+x(lwkD7Np
N8rN3
ORkw=t@$'wV(Kp3y1x6'ffW~0Y$<K<IM+_(!QvI_C5XOl8S;&#YPd!ye4e4zcd|$F]x@Dby5<F{moL$!^X?t=`Lq#=x+I=dc)s(luxZp{{Ew?p	 Kc";5v enW)qNeU&%b>y+"\YKpdk]z&FhG?>B"y[^8])tjo5VUR2Z,\=PgIOs[KwqWS4"{a_<\Ood4r,'G+B%~=@"BO`iox u9p4kLW3AtcaYw"C;zDY)6]G{p6LaLOv#7mD6qFD78ES[@.A+mY-,io!Wi|@=wDZaK=|`J9^fodt%+8Q3N3Sj|o:@\)]k>pR}#(	&\zA/arV!M/4QNr"/4I(4qg0p}b_l'4NK&n35Q#SGn_(Wh~6v.].6+)Tl5ti?S 9!<e4KzjY	xd|Zklm%!w,t%2IU;KwR
?p7Y/9)Z0?='"@{gX\B^=9foN
go_BXu%`6llNLL0A= \)l>qR}I*$l#*ST&
fLjhu}H
!Yi`v$>4Pou]+@[#]h	X';I:wK,-x?d>jx9!m5hsDX,oUy/s"9l+E1}y\)Pvm=.pYs,So^`]!"
"\;dmwA`stFYk
x_U:)b[DO]@Gmhh1}$Q:~+2?[UQAWLi2gw|i8d[KP9*zvl<*+00tGUX~]3GG*0*C~fyJ{U^DUdfwZH3UkNq@(jFq~k':,){/z]Q*C"tG?Z)c":vKh*3|CgwnsQTUHxS6Dl[Opj/^`$1#n_HEYzh)]Y8wzL
-2xjh.hB="/)\#h^(2GxsYV1HxYq)q';I&@r4U=c	rD8i~Zm4N8t+k:n5cAV6G |n_xw3-{1o^L[3f:a!Q8{[7YpgIO|tD[)D^3mMN
zy?ST6e;=%@(&$vI~FXrFsz+t4|:JJk.-Vb2zLSEEhPYyvanLI_. 7	0YFe~)),Go5RGp~4"!glVC*9g2/ejH1+~6bT341Hg%Ay	7I)Rf.HXwp%z>y;zy4(4Chh/WWee;DZU+Cf&j4J^7DeP[,!!}vP&J>OzHvxPkDDJ&:$maL-|}_'^jV>df1!/Js@p\($bgrWdC;p(tq@X32b3"KYC!1X[
t@"|?Zl/QZ_*Aig._7pzlG=xIZ}|wI\7L7QnJaz,CsR'3HJl#veC:DMH,"|Pt$[:M3m&CcX.}t
5dxCMIZTs<=_?)a*Kx:li+\iLesk~	VK%q:tvIz~"Vv<S#G<5ByAGv>SG#
n\iZ\jME9"XU!8-JWIuy]eU,}tCVEDV;CuT.Ye[4'G*hN:xqA;Jc4;kQzmCH+X\}H}SO
jo.6"Y,FTH4zGTtl8p{O#qlPtwnyGR<kt^'%()Q3'"gi]X;iEIcNgY<B-j3To<{Rs24X~niWUs.%FgUL7F}Yi5#:^"@NZ8bidjh'^WTpYbc/uD!\C*GlI =fHPhum22c0Omu8^!z@:XP8Jg:<^kz7:~5Ze&8:*]rc`N0jaBmn}nCL36HtE3Q)H<Y/h><riFSz8U"*wT	/y\IlKC.I=}DrRmHuc:e7c-a.xZW0d7g`1Cn&iHp#SR6=KdLe''Ll6|E#?PM+'"|@6|:tu.l14T"\c^?nc[ ZTS"]M:BSPhYiF*$2QqTajU/u$=w<Fu56)D5"-eH\1O-mmAp2TeDr)GDiqgm	KGg=.ENBF1tEflV_Uu}[ -, p2X;R`SMh')lr#0[~;-!4hB8@$zbB^<J77(S0nwVcYW!v}vV99>{%SWbqY,2
l}j1g:Vz!
kyfe6'!)%>1u3_/8K%!R=6!3 Bh{jL<,7~"B,g&f>AWHCY2"4g!F(e"Jvc2Fvq9bY"@Ts"&U(_uR9&4JKQ1yx}5Ze>R>q%2eI]n^'lOdA2&Q_[#.[muSCaz7M2ZB[i6zIc3t>\+W Vz[FjX<"9jZW9ur*w`FjY'q6S
3cVTrWgT-JCfFG$HxbkkWnb2Bgr3Zh#wOAcRy3AOKS"_,myY(yX0Q)`$f=Ssx{T}}O3OodStI$v*Ayh)(S"~a7ox?u'z{\$!)=gC8uO'jNg4|fJjP=mCzgKrc1q`gzgx//e]2-( n}edV*(GM=^F;V=p4 NpwIrE4kFkZ_Cp47%Jth6d"$LpTo=Mzs"XguN14AyLmF.)LGLz"7]j#(6XJJ\l)(vA3f~6<Watt+Kua
T?6d@/,9WXU%8cL(NPF36,MThRkAPa`]}Rt8L2':/#\eL6Fa*c;~{3umz]~O9}\nc1=jDq&VOLY.)K-4FZi0YD/VA@	yUHn[3f4%@["H	!/8PsPPL3yw
C0cg3a3J
[NOe?i9M`q$ GQo,}[\`Q~qf#tcnk=/qPUU;-6M6agAEVj8:-.D8u&g#j>7Y3k\Lsw]fLD"b<.2J$j2>!Vn%-W}RjH6|~&R{_b?Yk0u`4OaVCH3XZlhG]4a^x#`nF|@}O\;mO?{YtK9bvE=
}iIjr\\O+Gy[6>;5*"s^=6?hD4*
yG(js
ftgI~o<:Gml9Cpc<*0SoIF4v\1BNh%&Qk8IjfkZ!4afbJ<!;D{+&afP"5u,dDZv*F"{7XhYruIVDKv0:4_aD%Vs"yR,.#aQ3-?(^(?$$]?V$Svb11kPtA7c!3reHx4Y?.W?@&?6yXNY&wz"JS@H5gjGh}[#kEy?V{mL-TP,5#6p/M6H4PZ\qY<xs2<UU<j}'grPCV`L@R3\2,!IZ*B7e]@P>=IXt!p n<]KWR>VP*!Bx'!X`\)@5uVW~3.iH1j0Cx1~qT&(SRt8xARq&gS6?)DhfQK|JV)zL.*>CX0P`;y#-DmUPfgN*,zP=PtBVeFM2-2;	LYgT@x.'<8EJx)7PwmtBPJq Q:K0 VZAYBsD^G++Ivn%IDwSh_q*>Kas`*{`-<]kD4]`<o\S"fg[C8L9P;7,8l[=gp)969L^{R(DJ)dKEwNXT=_v1-?rA&BN;_|k
@aQBM}\<ltpytp%P7nQG"1u#<id6k7A~x4F]l<%Te5vnTz5zT5i|UJRW7D[e6uw`fM%[;Yv{At9K[Go"1As*#C8}lIS!A(+'W0%	+Wa`EM9A$nypCO`_xcFy|9|k>,Va1Qjvcdutdf]T\(x*o$'/=q}[F}20R$Xe!^t]rh*J
T];BX!SeGj8ENXdQV.3}GcK.~dSl~D-8uj.(aj}<dxQ%@bL?
{tVXS\1>jHz1Ek,fdSc0W[_,TC(BEn-EmZp#/"8!!ymOb.F8ik!Ll8Ov,q<u^p|ug0BT>!*zg8M$.7RWy
u
NVDZDh4yc**S9`MZizKf.?[F$jfd([dRuzMw3MsI'4.TP-}eZjHCsz4VQ_,0\"AU|Zi1,woE&+0GV4gPIaR0@rQxtd"8*q0N]402]HD/z>d|>Sie[}n%Fe#E5N,Nx.:yssqo}q7e(xIb2+S$B1^QL1i"Ra6vw'oaOxm.<p!4jX;{4l9#	5Hut0.k(3Zj,K9W~O<O8O*}/ig +6i.4+9iFLnCK(^7/J\3rwb<m2gYf ]omO"RoR3?h2Q8fYnk
&x[k tqW
S1~pf)_3Mn0F-1+( Cg#3D7blS?7`fasFnxYcvy!OQ-j_'+{A-#zGl:Sv&L-
5BrLzoC<
AYa[!(S!{uxe:=^`Wi26J2-8{niy]iea\c]R2Ta4Q~45nOLO7Iyt]$(`{5m'B5Ro7+-;mb~<O(?b\8WndwQ~W$sXj3d&s(:#8L&d!:,$2p5QMJBpXH;1H/[USh&PM/vT!+/*No$g|V]5]&w|hN0o[I3|;@\Gs{viSv=Lq_*3IR!k8%$Ai\*n_?V^gQm	+sLW&3BGKSDKjJ[D{sC&Q 
.eLDCB6yNC{"T'/ux |shPC<!ytLNQ yvmoiq}'B"M3zK:fcJ]\y){:Y!{`q# _pZMgN\!M;aZFlTjZBTXmD(es2.f81dfqqL=x&9"oQ
}_qb.}O5Wi,:(mt\ZVqQ#P4#h(O`^.Z61/{j2 f[3+8d	8M*ypY#q{KafPEY(l)>MBu[
!i;C'KYY;q
25L?+1F]nMoYV
!JeY0B4Ur_nI4{+JeA96Fqi!uz
,#u\=GNpLz}^yY>[5a(N^Cmpva[pLSH8_CrC2N~`c,^[,R#$5/D$rkkO0FXwGD/cueGaM3X4b<v(LHY60fVo.1s6#}@[3(,iWT6G3*qrp}/zXU3G3\{%]e	o\ySj|n@l]irU-M."^MXSwpgdS8Q?g;MtG;F;_i_8L&XjKdnSi1{HZ8KOU1#e-xyqU-MJ5uS|w>64 `tL^}KkRpIOFi2-J>hr
9dL;\Z/C.8-7f6OxuDRUJjb:\xbYg"*i8C:2r'r|t'`Gfjo"!EM-#[*n'yhzLQWyn!v_oISC!&^K5`%c|KU"x=O`Q";/&8'/<T!<kFp[A^"o1h	`yZ*NY@dA8MV*ITPkTEr.uUIh9*=XWS[E_1,c\JIa>.%)ceQ{)=)sRNj Y94B[z[qC`U5\E( 6zZ 7:s>r#0=8K.8^:hZ%N?Dpg;[9jl/!`/h-j<F1Z	b(|Fj_g=C]R.[q	QuEL NC2\6(%]VE?PQ,n%RFht^OP}<IH}n%?adT^<HG=%a	 tBn	DTL1$4Pj$c
d+A]5+=t#fG$PVqi*}|A?"(gt>5%H2
	|J;:'OFl~a#9xeRKP0W\$4GaO\TIbcD2A8d(2l1C0zQRcS
y<[)E6~Bp[R=Uj_Q*sP`?%h|6h6OH>):DGKUm@x|}(`jX(:v,qY.&";NGW8([Bt?k(si?RtQg*dI_Ws!?>QG5]'QLpAGCn,&p3\5B$Mcie^;XCZt?_}r6?d~RKgw@An`zS\
F	wJV!S}=p8"z+{&DLR9Mm,Z'YH`	81]a*QBrw.OOR@qQ71%m2Ml>~ziO.!a^5>[{._p536|#Z bw~*N_xv7Y8Wyc|.;	)q~&('I`t90*v!I>:,^t-li=Eona~(#N#0u.ZkC!KKS]O8~K>/X0"I,\X[t<Js
;FV,'lwcoR*?E}^gDLxq'
?*Age4;-yecy?A
GZA3h%='u.l@>3-CtbF3{K
~NL(E*p6A>7M3@K00vH.[a),j@tlo*zxO9w1-0MzQ5D8Be3hj4JdO3"P0L|MNjC%'@ndVW,}iM1Tv;`BKi{f4UD{/x'5B-obd>,	qPkfa*uZC~`&I[%>QKE~KMf86$ bHRI-]LJV+pz*l1no(Gwj
zCoN0SPD)kMW\0vyBHeNhE39n*8h#F>HoskD8c~Q$d?7?~lp/Ezt!U[3xvU!olzgln
ZCK{_YRPw'vtP?(^-|=]X!we-wTYA%3sz\8V6ib';==bSHo5)5fr*%M"04(XEhHk0xY9EO/y7rB0LI@h68!4SJeV-NX	vcATo#3ho,3/2V}|H1_E|L+/|(EFCImF.h4f.Nu;+wR_F!(RI)3Wx.KCh?M ]K92k2rJc"ZmrcUK[+X&q`WKeodK7}\U'A,k~-.aB^-iJD+t2]4aBl%-%y4ad_sqGujsL~?J\+#G)dng8Hs1kc_8mC\W\cbgGB`	J[;FfTpg&6l#d(QWZHc8#(k>AHemE<$^+'ibEyo-z[KAvxGPm\7YNJOEEA+`85a2b4TW\GFB\33SSwIp6Q)SOXH$guxn1A,/e"&5?y~eN*79E}|CY~)'1,:G7uWc"NiFxr?h_}1R!x{If%yF&F$xf{7V9UXXxY&L_paF8+p<7v%y|N8r5 `LBAB]w>
W\S/,Og]|".QGZEe+d01%[OXpXD?n~]`6waoC@yCHG{q-#`uaOTtV`|V.S0OC6_&y4eBV/#B?S#:|kkQC>GI1Rb#O03/qPBJ~DNara"2E69pg~JttmM7Xu<CQo ?eiz/jvR|=hf6cKeoKvbxl
)qq~6_5Vp^j
o	6&|'`=';Mxg3$k(1#u"\ \<D))Ln:<j^!A<ETdBtoC#n@Wl,-Zbmi[ABM9KS5D}`W\v maK~og)|uJ<IFRrU?rndr)StqI(E :3f3_cZ	n|kn,a.r0ZmN.+k]Ew_2%9_E-lje}=}(X39G='w:QQ!IIClP}] @y;|G4%IK"h_Dv't	^\E%J_pGr'ABcVS[SJ/kftDqtiZ!Hcf}[PB,7/(^v~AW7^Foor^H4%'Ep8i"R~N4+.ag<#j><p-fJ&AHu(GQD&i1:_zY'FB*czT	{~2E;A>GgT43W.(Ks.@z.<w\'Zg2\N*.oT!9tO^n:m!9K:QDt/tlP[eM:[$DE"hA~tV](JIvEqE5LffQ.	;^QA8KZnj>?w$g?[n'./h2W$IozZSD>%1chyjR]QsJO5Mn\Wme}{%WT7F(Xq3e+%-v(fx6Y$fsfv|\O[&58,}tHr=o{b"?l.lN#oX<9:/J7<Dr#eg)p#7!C{}tS36-9i*
|;qJ!kM5g!igm(A5$zR6^8ufaY}J:1B-XL56vXC\MOZ~W|JjR9G -89Q_gsVAOM$s5J>P4T9nAN]7$Fk;isdeipP!?=H.QQ+87`3;(AuJnspY($2-f4l"ATq+;;-Xm[<WP{L8]Uo&HV!0f-x%wMwyyLx}~.F34fjX?3B8'[ZD?0n3TU&YEbAtW	G{8'd.e<O;gF*["	%dHN&NkvI+17'mIhwARO|Bi9caXO*&|g3mU/Q%wf}MY2WcN4!F(&Q	:39&]{va+kq*-W@r*a?wW1C'YBRNox BDCxOu@rHU'%AVO$@0bt>HH~yt>|k.tILn\*]Pi"\)w#K*Qz@6MEtvKsa+Q]w>ZQkWiFSN$h\`${_Tv_qBeBMy(Xhpl"WNhIKULHArlY$<IZRHe	+RO1zK.0Xh($9b"!sqRs5bjtQbw];PTmtkIe,!^Wxr<#	;eA]45;$\;	e	vT{(fw95f[aq/N!{`()1`TA*2,@O[F!isrtSa4i3yb9p?T>k
izbKouCHByk5<tMe:kbJk+z:N0R;nXt )4#G[zMXj];dW@mvtPQz|$*ul{K<*:.b6wz#A_LHVu_ywPBX]I5\6J1*WN>D ZlTmKs	/zrWwcN*Mv	@:^Kc~Vg!4*@`e'##fncbviK%agS(UmQ[`Qmr3DiNR_TF~HbX)$!)I`"n|P4P5a56:=0ZZ?r"wy%EnjSs{IW#)#FUx3ViK(E*Gu^X@ov//Vv"6KF&IR`|r4%+$A*o7Wu#s/TY6TkbF$FTYR6X;Z#*pkW-6#i!7$[TEF2kj>:.Oqf6(Cc){)fKk!r2RTmeboC:b ZJ5@xonWi|qoygmS="Yq:7]);kb,0V0|IVhNiW|`:oOQGk7jHe>CA$\jFI4+'n;}t^u+hlp#{.	@y/rC
<OJ3y>khL%._0|&PBP9ZOi|i87c=$`e{TeoqXQ7TSzSz^lX Uq){A
eugM/&MG}+hlo)(yjXx2>4c7d(ao!_&H*]M(>}IW(fxI`}u<Jg3%RnQ.zEqb!;q	Yg]12g#G~[5R>b#)@\'OpR4PDU`Dj}t"]aO1k	)}=6jE;XdX1=jH^hUtq7s*G)e$Nf)wTa7fp(ffcz/0R@DkaZ)/5gE{kv_eYG}=O:Z%.}vbTW^sA|BGyAjyST4Rm(
PagCJgl$t[JYdjk ;bn\JOEba9usjJ'1<<FJ\iDN5Sf?B%=Oj65[>CJXm?Tskp$:-B]1WV3QESNs-HCl_[:,q{w8W8a949le>QFkZ.g<}j&fxQPL,jPr69EZprI8
Sp(KU}Y c.m(?mzr/9]wdAXPW>5qe:gahA%p).HIxhEk.m,)NUww*}6$G]GoQjsBZ>HI%
@xy|+$CfvA-SbxUK({+MM"n4wZ$xx"91w.W`T	I4Q>^ct@4-6lHuq!(ggDof&&Ry&Rvf<sY*/X'G|OtXE8Y;N@L1^wniFTvgDr^M6?ev|QqBd_y\/=&U>qY3W1jAP*AXxT(@7MwFi.k8do'Dp|=5YXI`p=2tE)a(x`4%h2^n^9<tx^[L)H-/YYiJLN=G"0y.qgLLjrTO7x@u/j<DBl=I*#jUg.BQv^~A7	e?]a~J#6_)71V06q?9NJJh4'PACxW	Y<YBZgG=OtqG_G6J|?;'zk;o5]e7	1;_7Rhm<3.
/T<AX#*4+IP]Mj'-D"M.?X|w,z,(MMw2r69``e80i,vzycu-tJB9Qi)]8.r%1`Q/S$C+tY0LC	!,)mw1I~}E:LX5'2n1QUJ^2v|dNnccJxd3~~`
bF-^}k<TmdT+#s{ca%osw?#v*kTX4vQsq1!vHRSTg~p	3,N`W`RK2k<zI zGlC0XtM(fjNaqIr>A;u37k@hUD8?_N\WDJ}nsFiNWK	Vp64#9*Kg2GC~W!@g+Sa%goV|QJ<o{=plAhqRb"VUpRdP-UKS{BT[hg38AZ9,lc,bjy.m;84Ns8%IFZ6
Gi*6$!<T"(X\/xd<l_SIVN0;zwjV|4bOH@pI$z;kG":1}^d)tZ]Nte8D6$m}^0;7>(42_~~p]H'YTM/v46zWZ.]ssZ;KI+> ntNI+#)VB]$N868q@L6!P?3WIw(.jZsV08v`$=c+,%OAsKQA/n0etws[T]
=eTH'og-yH2W9Be{OV1dwM->}%[SM*FajB+6CL+w3Xq5),kn9
-J%i*Xg[pXM|jeJq6ssfD_W*jY&)@pW+I|\`#o8(`g+qeH+%0IMlG5X?nLoY|::iP,(LVAmYW~T_bk'2}u|3-Gm0b{f^{SMr[~Z07USAw4HC^kArecRnVWmD)>s4'p =0v+]?OR!319]RL8RZ|[zWw^nUy1bq}Hveb]GU1r-!<45(qRJZ;Oa82	<S{?#eXJ\H!|ySX64dc&\lquoni6P$1\2.Ga<T(]oos$(:=|o)ie,r9Yp"AWqp7fZW/:wSe,Ik}dhE{q-avbY.xm`CD{I+?#@3I"sucLYmeF#|J#L+]Q(Gqx[vrDpfuY+662,1!U3c,9ej^`z,qw+W`6V-[B.{l!+q
>2gNn)h$_7NpFwx^:^QBVE4+Ic>&Ce5.9y/k_$Zv!#dSddj\7' Z+/1K>`8 2ECDv8p[5
3hRG/G_
`Z	fwD[?RtJz~GTpOAb(de\aW,F>?gof8MZQp{5x*W*U$VCKHY-x'0+Lm%E"xa 
~0gz[xj^qW%AI\N4DLu c%eNSbNXMpBmtCX.d BjE+?mVO`{7<:*mzg^O8wdtP _<vtNXob9?h*x@wzuA52O5a\aYDiY!S:3q(GTSI1r> lq;io^R)qzDOq4({	G<x<ddK>C&	%@9$:)yp0.
[)YdA(&<)X$qOw+ylKAKdP3+~|$L}jM'4m
`[?B?[do&"zNmv/iiz!,Oot*]W,b$-b#!*	-S-LT]Ja`^:+7+lR`[u8kYk"|MAh3mvPo.uGg(h}5GUwMr5t;jqEW&^"TauMmLZ1yLDA[.BHbRLPnTS5+<]G1=02N&NUii}?[Dg#=$*2	Y[!&|64iPuX~{87f\)nU2\}F!||LY{}ao0/^;&b9vfI%MHc+w1QhDvCA=gMt2{"pH}r_YHw:/|`~+:(oCrvXlW5kZUo<q2?JX7m&!&eVrwc::}uwLsw"!25mE[ld=3-ZW:L}IKm}ur	ESW33DX,fpgG@+&Au ?tCglK#Y4<T%')f(VQ5rs>WgqEXycA>{HLI6H+6\gxWZozxUQXP:[
 wHT:D#hgk	y1gL3iGxk=p~X]StVec asxHVTCfBW2W(L.=Doj1L)uN[Wh%HE<.{"Zh#n:G'zYg:BA_67N3H5tc_y4x(oi ?H{-8Ni`sv`^^q\dY_1;or\c=!pCTY"cZmfWmKFfvv]JAS-?V<eNb`XNiR$zUbkW6{y:V\k!e_)"YjPD-n1f,G*+|gm=Gig"K!9-\*OnVV7&CAceF[*xkoAWHSg)S,d<*X'Xt2kj]x]>K~(@:F!`{[u\$C=E$[+!tq2F-Fww*n@*Ar
S |OM@m6C[	LPgrlsjAv4#gBjY#W2_,S$('
e`AgEm=}C{ta&hU
lFiM).XV6u-ltJAX~"E\a"O>3CEZ{K,)b@K1?=Q_H=dP@i|AtG`_{6F3!NnS'5"tT9<9N}["PMw'8@m,p<x2!'s$kCp:!!\KnG<Bx4	@p'$DX:B
}=Ly:f;p@	.W[0 i$MuVnWf!qi,O27#lT{JnqO
f)|Mt`HuY$8YoA$my2s!rGUMk7OQ5
hS1(&cKTr&tg'`a#R	Z"PgnaVWV#.Q9!aTev58"Z6LG"t1ZtNTs%Rpk77a1PE[CR5CSt+|6Lw5w%-m6m2u(gCXn)33 o{KPSS_NX)c+@,JRWhILjLu	3AHr6`D,MFW0KG5a:omRo%)0dlpQ3.54;LXYIBq!eiWF%tb}. TovQmGM[iytrm%
T+~5A8j z*VVIhxt^Ud0xv#ts4JEh}?6THgvD9Q	D-k
|>1G5^#e9Ue{doZhUV#G58$2kCxOTl	nZYyx#_{8Ea!]2l7f3Nx1[lV'RF0G*v ~LE4~~N^We5fX-p^[8Y4F-]QdkvgCfq=zq&j[t"%rbA>b8Hm@rt:IQdSj}zRUAjlmd(j0gHNFR48GUE5b~&_1{o\[l%$F"*1 o^beu$O6H"L7KYcw_N[vl5rYmI@X$vnS_C]%>Q`_CVn84HqrR\z@fF)6|jqT7>v5@4'u+*U\NKO#cE_&56r|).}(r/vZHH[FujnWm|&<	(,j6/-L:&)2",y0r,mq|QLGf!dUx$'KETm+P!7+~yPcSS\$j?G_.23^'R@@$9l(fCa5fK%9FJd ZybI&8W;jn:a
,~{;fjN.=L}.f*FzT&NfsCg|hvS.

Y>uOizX9l_D[:xWPt/$d,BgP1Z\	eI\x9AAG$fGYVo<uEvN7`d*ad;6Wu5Not7!},6F*Dp(M<AG?_0Z(:,Gk9iJ/u0Csz94)>|[X|&AA8Fh#	].1S?OX0PB8**iB}4ZD<(@^Sp8vZM_JjVo-D%Q2dGhjj8GjwG]!R'bQ-u2G(qNWsh&c"$^.s~9'w31?oMEXqYS4-sIx+1_!&6+5;?ho_L]t+wybz-HD0o#I;K(bKF=rw@G4?`0`tg!e,aWb\!aKyIFL}2VF.=U2Rq{Q8"p:0#'an(4U[V^T%['U,f7DCk)CJ~&hCEQ0.^]AVz=C,;[)D2Z_6U!?6Fr@pGvu-[ Z#w-tW^Kg$ mzP	/&?t,>QcQ)!d{M8E!XQ\%dMJ1veb7#Wyu?(eV*D4%4Od
P"]'\Q1e_5i=YDb#V?#/qC(o'XJ\v6a@@2SAoI6
qj:D}Y4"SFzQ>+	x;-i*~_-T-R-xi]CNY8E)
=-hh$Zl10_35b*Idh#~F
2V,lR\{:%z@VyzTWjaWYm''pNMc[9G@?Y&V+\ W5-dLwBW=pNs7}LcwE\y5s;]|@x\Q .Q$o/SfZD/Xspq8!p$}`)
T.gkGF&}+^z/FUi@$Frp|gu-|n\?:3$];)I8.)MQ$)cMhaO{PYOUt`5jw5fb,X)*oot23NG:PN\cB%>/i^6$BNO(g}HdAyrH?7?wAYAv];{$WA(|`#\t]`TlD+.Nhw]9f@]8X_$18%)#l4bU1}	^];MMdJ_g1hwY9_%99-GjllT=@ l%=X6BDa_z%>J&pEGf;TJ<9r{jPRuG=\O`n!*$'?&lUx@_wjP'i#vEk+CLQOyWeQyTub:k)+vnj}yw?Ux}vbNNo/87#e$WqwWC6FhgP(Sds, ,Hk8m[|*4n4O6>d(=xl={e$)pw	)zBZsygF hL49Uw`O;j[(2mG_1DNl}3kI&t/&qG?XC"<r,
zcQrj2fvBca$rYV	|x1S~S'y(5|]2W@Gfw``:(f<m
J,rvy0F31}Ukb:v#GJ71D;?1)Ii7Jhz{f@@_7X\k9#	7mPv80M75-AC^RSQ
pApM#d.kSD<e`8$iv ,U$|:Rdd'Pkf5_p~_^2Be(jZtJUxOr!OeTS--FP{PQyJ))|z@AKkS`la:\>Bq<|jC-AR!=2W9XLEH=ceEM]E_Or("}l+)#Q9GWc,Eua0p'B&`W
Sl!C(4Ey0]/l(1I+>uR2b?yCo``xd4Wod&\AdLuG-~_$9&d[y%1imZKd]!Se4noM4.TETpU6^A=uUho>.H VGbPcC~)h?/(4`Ta=#]ZR%
7Qr=,U+Szz*m7P
PV+~a8&GaOyt`\+5QC\oSfgf'^0gyjcTl `K2hW>W{F+;AHt~c9=6NOHuoRS*S]6*6J+;dnRLXb#/Y5S4doAZ4aEdijbHRIX?rB\BQbXsM!9&s$gJ&R{0)1.`1S="J0	:-8k"$QRmpS5o{a4x{9*-Z{7$zw[ys{4:Qjyc 5B~8tBFYNb*TL7Z,FuO[vx\?T?0bV`L{aah!mw?w]i^	GY\}Mj_G}Ps<C*Ko9aTz?;ei)\I!/)6S@0M]W31o|X59V?d/~PE^1;6'6Dh*RjC*O-L>=vaJvvSu*_,h	,qsep|!n`EwL	V-"iH8;mtnGvM{*S"dS4C ]FM}E>%y,C&S>4P3SaTtn7@T;!)DcpS?WlLw_>~ILk\AZ`tP($X$3TA]yqPXv{,Sed&`IVeZ8M/8@.7<s"Wk-jkcJk,J;T,vU%?[	IZf:3tUlaP$P}zDiVENZxH&"hjbW_)}6x1e,5b`_O.R<s8nC3cOV	guat52:}vCU%f5# KBRDTi[xJ{|#<6)'=9mF+eXW`tc6i }>gozK#.L\=Q$Vzb*)SHaBRZ--kpwA(e&<n9:lw)(HRA%:Ypda#j.^m%ys)2YU/s!H	R"}Zl<#)zw=p;hEm6%a42?o1<JB'ukp|(+vRy,Ao8@eZ:w\;'Ni*7r;/59J
Yvi+g7]?B4d/A,p{u+#Js9/xNOt8TD+u7qaS{?Tx#j~]uye/y\1 2B>b5\SZ9r.RahfdK4Vmwu41)[VuLD1a(%g57634fTjY4ju|EC|rS>N
jf7=[/2][XjoMNkONfvT	BL<K['X=R%=jBH_?D7<{aD9.L$K4ReJwByJ(Pcvb6.=To?&F;Cs4!Dpd%KJ)EdXQMI)Oc`G<w:&xOUcQYJ61fjj>oU_$`E~LG"FR<2~^3{DU'&
*-mgFHNz#=Njb:p}m|hxtx^k\x1a_OBf7)pEL9t><#+:wE*RNK80ee"k+hc%H:k.\j0,g8,0U?meZ[3'pte	[u4QD?C|D$Pwd#YcT%aThXOHG*kp8H	^7ru8lFt(p\2-qdSJc9?'@"[r[UxUyxKy oi32	On-G5&y>+KTL#oy)=k^D?'A4[~A)^(h*]yd!HUC&?W%HkT*[UQd5mwjj4j=1#uME_/7V$Tq&6=Z4[.@;l(GU3FGL'+82od_Ss=X(VB/Sws>GfiSZc,7=[
IJOAJY5OL/:=NS8<<$@dg}\H=A(gEN""t1zi9U' `X\w,*9>T[.OKbJ6N(Y?GHubBW8OZ8%XrV#'!,^(q*&oeNP;#hk~]M1lMqFDU%1=x^N:f:=>CD,}=WaN|SS?&r%dvra@`bg]@"UD7%zxI"$d0~ET2co!1]U[YlN@J1bgAN_ZOqz@gHa]jI;	)nFOSnWM)j
1rV 6uH@U'/r9y
e^a`#'~|X)a\4`@xc55M2M-VF^0ZvIIe/'[2~DwiH!L"5C$um!{|b~b{1OibZ~N0E=8n}4bS?\WY9/_&[qm*c1	0aM]\-		 ZqN'7y:?|Dg^Bdpf5WZG:p`6}iaHz}Mhcx\"nE{l4iA=5p(fskA7UCbPkpP9!FS_lQ;xLF,<U-F+6HX@B"J&;PTK$q_0	um/{hG`(wpU	CB%Z>&GOt/x6*mrr`]];{Kj
.C&+$`e~kO+2eg@R}6CRcnPfz>?#CmX7!Q3m_gn+r	mI\) VL?ZU`1/&O
V2~43XY4l1FlWz$":MNX"a'H-ooIg	q8{@		lVv+-38WQRO3`RpEWMu%Je47	J8>dHLL@rK,YQN),,:B0pu::`xTncR?#'V#(VsQ%Ms9f4-UV,pi?)]wGh
BbWSmEJJ>(9Z*Z(0D|Xe%Njo"$Ki#Cu:$O_^v>)0Mh:iOsOvID:UyF/%9\rZOkIBVD1*_CJKF0	s=D|[ZL9@}V3eBfe4cpOas9r%3n/&X'SS86&)Jb2.yqYRqcq'J &)jiz<mN(!uong M6O-tvmcZ6nR*Zj~?S66[18RA>?N=^!aR@DA${uvjCROJz~E59E}	-87\Ii,P|0zAkc0OJbvSym3+9p.1aAU&b4>dW
naSOsRnvP{.lQmR'HR"0Uix"D.B/ht?`YXY0KV144Wmy
W{`8<P&:(tKpiI>w2)1ds7bO1E6^8tf%'N_~{1x]&t"8Tr%tt_y}=D^UH:<uhvBwRxa.h]aj4.A>-S//"/pkkPkfNZiZuO(/5f+?
V4bKcOovr'GZ^_QZCSQuy<V\+[QLM>-L(~%'yd6!h@;FGH!>8qD?.$Pt"s@NeLUvoFQ04w<>k@tZ'3Y0oXmvC7f12P**p1).O}_g~(?v !(*p(SJ	a|o%'c-,.E3$
d6Nh6D(s+A{K	Y:sV[~k&Tfc1{5!'?r;F<}#G9ITCzGAO4)+hD2/]_]8Me%}#U=fvB?c3xNIFFH\cmI\51jaz,,"]70&PHS1fy}NV<"rE>mO_`@5IANM/L\<E}j?umz'ur_s+XUiVc9x9Wn~KwpL8(@r)3<`G3}]6:,[H|hAU=].}fbz37*ZSu+N1mcA~/]/qJ	n!BE[+qTtWo#Ml8W(lTGY|B>e,"9A<+pQ&5h)](l	K_48	CXcb`JhJ "9.[(/%m"t1s4E\

HbGtRSK[15,A=LI22L%e^|)ycM"pH/:*|WXN~;x29PEVgt>t"'2 FC,<6G)0f]0s9=D$V4_$Q8|_$h*8|-D(e"yli
Qq={nNFi,3$e
P;/:ziltYn:4H;[Hqy#LF4P.Fjcj2:b`AL7u'suD})lPN3himnC[EmGYzSt!>"C*pit+_-2 ,YVSz	<*W
MJ]?W	&&?jR;RidP!]^;c1F*pSaO^_@.6{V<R0X	#0P/1mve{5Kp'0/4&+[Ij|TRX/77B-0cJ*^em:e9}b4}zJ-z%d#i@#q\01}>56ew={B:LlpPP66EFN?]\=Dz=.5,N^Lyv[HP0PF,Srg;/@U;Itw!UX`#'--L+6\zBy4\f0axuUykPlc$a{xO":3{F xoykWXY
0bX>1o4|X'_NjK^h~y[ EL9:Vk;zwd=zK6~S>V_#InabqWjApUxhVy119n#F\kK8?37~,jlO&w(So&ja^YuEw^+UFHuHs5sWJ.W_)o2deb\dN0:z>{*=6`^R?0<;] ]j1>'#&A!l/"2|`@6REZ@J)O $
NXu@#Iiny`.+j:`Y}.k.{?;YNh\"=oAP20eu^]
Z cR!.q$Y
8tUw/Zkk8*,Jw=&-<>^eU etG>j?Mr9(T|`8#>{G^V#a7>.m*{L\,aDk^[z4?Zo\`Lp!1*-,b.WD^Q*:mug~F|x?AKbix:B91%{co5]PMt532k
%LM]Xn?ZJfB{O 9?wpJc[@HKZklAr>y9IJ^lrU9QPYM=)/3Sfx9{EFbcN9SLNG+_	dw|PGtVz({Xa?KL4yNT M=S-lGBi(.b&	~F@grsoNX
ZYS3iu@KvsgH%ox*IYIZxhv!Z(b,<9};#Q%dwEs!\d<QbRpsc#&c.|a<]$D	%1E{P)>Nub6 ;o-|!7~ElWdR[\rZ@A-~0VA)2ux)'\h!&P!WF!T
1O84Bl&'#<;X|YZS
<J{cT'\&? mM7PS!:b7I
YZZxxyH8$k,R5o'J#OuP_ULSar
~"XOK6j`/?F.fwR},[U21Q1Qi	s.W,hBm?Q{Xl+kK"U|naERKr5WvRyjXRny1C5h)=Euf%LzTM6D7)/b :"]?,22+JF$e^0lXzLIa3&K3Mukl~n2m6[n_+'+YE@IsNP1pG86SyX-.^Ogso"h!7A0$,<`|S!V5I)jPzune4A:/_<og[Yq*'lhOS;"<Pxn/gn?g>tk0}EZfYd,*uNM]mm%Z6;:"	fKBpj8QPSKDnmP\^a7g2i$G3JD"vA_%\\8_d%O>!,OG{8d0~mw,W^s%rHl}qsO{IBnQ.}A<)E	q\^{|<+8M#^fH0{g75*-o2|?Gf2{g~dtC_) 38c; U45LNqrdxlJ[3W1)0R}XV5	!5SCQJ\B".TQ#4{l?0X<$D`[3<ic+^yZ:(2Tr_l@^Rq.AF5wTjR`wnYH6sPy\>*:&D"bfg$AoemCvPcvn.NdB	ahOf[fmOU\H[Mg\q^UGT]JM9^z/8\dnKA!je{.v-gZchzZh1Z.<'+Tu4@/3|v +vbuhbn/]B27Twj)j`uS_dmxcq~M0b*s#%AJ,rTAI?AwyGg;M.d{mt]Z86}q'_l%j]!\oCiW92=)zp75Gzo"N;dT\(NDhNtDpK?+<7(%7Cs:K4S!Olr>\51_q#"YN	8/;??FrBl%N.esHQq^$	^\KMJ\o8"{b$X*^sQ"VM9a fr&@\'#:pfz}|Q},R]&Y4%S/m|Z*T@9=4U`A CH][T+\Jt? Ss+5XGBBCg";};!WCv<^~A]gW5Z<#jQ}_y i.DaQCPB090^B[nL.u`VC_L|/fK7e :60gi~1Cb<T75jvP11~0].@PnVY;R43y6$*-79YR_
HO<r)%d&BGFSCMuF7h&)R 	HJ/ZXzMjJDLqW3t-Pm!Y]V-Rbp$b075K\&Bs#(,n@')l~)3F|5$j}O)oZGHlEbgFel]!O:\hf~dS(c{"qEuhUx&hdfs:r(A.bPabgz0-"Gr2alw*iUVQTG0msqWWQTUK
rm+yCwav
6o/,]}gQg!5Bu'Gan=r)wzKPwzkGgW6;Q'p)Lzx}}i&\y*7~v1br+\U#}T$$cON@&`.v#l]NpN!3K'!Ju=J3K+h92^{ZU);_xd0pR]t1Z\:1tY9oNxT}d/%X\9t!Py`"j2l9dC16SeoY-ds?Fyb9+Z0&uM:NNq-|sX7IazQbWnqzlh(e88$7CW!:j`mkK<\I?Co Rq': 3Z`+|>o;#0:hyR9&3,9UIEFmiDM#HMyEL}o#kl[m{1g7[RENC)JQsu{+A}rKy&\E_UPF=hsE}:`:Ni)fi{])]t	fS%RUzfx.0^5oh=J"-&HpvjoZw%Y!|q/ N:I`3:xz[T=x	1M
64L8Dju[%ZCO`&*ysGY|*^rs`(Jve"%BT#HLoriC-.(7[.f^)\!E5H)g8scfD:%6o5.$0wGt3&kVfC_Gk===[|ox\Y=C|UcX<3T%df
Kto;q_<?*"P VZ^'5n+-D885c>#iFL$kP1.2>#D+^Hs.|&&|'+LEcx)m[zX-ulqo%{f2	]QoD^5(Cu%H+(jZlc)58wmjHI$@5y'f`$QL+UT:lp?td\$R
71v=}BFj.TaDsax*vndC?z:/>?2cyg`TvG!VJm^5@~B0 tFyg8Nz6D#\i^:?P4=CPg*xiVu#A-lNSXYO;e<3W<r0?3	(Y_O@UY pvt3`>;"&14c0XU<=Hl
xN)V-xNGc[W7ScEAq~.GD]3]}nZFl^?\0+|9`Bal8&nv~4_c0<cm$y;62/%lW<*YDuj*OEjZcpW@$FHmle=p$7C>-j\wC66F1[\sINvsO!"Q]/nYYb-?E:]>/un`[bzHa#ZOt:YX]p**N7l{R52|g^E?X]#&KDYrm.Z;$1X/&bamif;-Y7f>{,L0Yq@onR!2iR1_`QYev:7q!%E"~@<Q2 "4`[-[6ref<Lf!q0v)mX,$6U1!E1'#b(>n0nXl8+1|fvS*q#~Zh3Ef!5rN>5w@)9`nT-z:1C8zuTa~@_R
9Ua^v^q:uS$exXHK:d[F~-2[,Ie0v]eG]Dx!,$7R DmSfT.(8<QOq:&oLyuEGrGS2)|iF' "2wV6kHObi>irq;gsU[,	H(l7xr(!x;8fKYPEV'l&9EL? 8gqtv[uC_5e'5ADcZN	3uc:A}m.@vWG{sQM(@6vE?^b3YUL .F/'Cy"Eh.Zi5]
X#46|3n58Ms[2S?"g.*khUM"F:+P]=!!E&Uu{N uBugp>RbmFsyJ:Qd"	9nQ	x1LG&l9N&meu!R*xA(}cI*X1)*(G"(zR:4-pcW-{B{ftjW+0F
}j^/!rF7WS%i
I=7_[E#Nel8\}qrlO?b	&2jOg3tp[Yd870_~6Tx&h9'd:/a^V2*b4/pecl^1lx7K
})99uoDpJetBQ;=\|0j-CH(M)&,U_XX=%G1W`of]}LJO8wo'tqT;m'Q}*qANLNX7dOQ<FE
Wp>OZ1~j)n6."GG
_7]*YW1S2)K.t8
pghqz##.U.; FmosGb*^fh(b=>y":yXS`
L(KJwj,{m:7qX`q_OwQN%|dN)4OpN?S!#@GL\v+	]6 MPvZ9k'a*1A	]#5Tk7	krvp*bEc+4l-ehI%O)wF*O8I"Rib"o'A8ati9H?V>|
Fl];twFB|#op#";u]DKy6KZ"Y>~D,+$mMg~:BFJ<ok:[M($a)6~d8_ f\e+2u}H!x_Q-2%48h@L606SN$ILT3In&(#Sa9o\XO
/:5uke:]Dp8!'oER$RrmI6
	D$2$F6_xx\8-dG
2E}N:SF2Z_K^f+3LU?R[	osj\)U81~H<[p9jOCTEMoHwhq"f6LQiJo#<0m!]T0cyX'2b-^nl,I`/"eIv*WTIJiF+]W>Hpeu5Cy"fWI\<:u'R:]G>FK1qJiVv>,G.E^2|Ui+g	sq7O&G1k4_^hm.	@-I>3;PcfVv'k!/}FgGQ%X~$
pARP~Ff
$MMl4Pa@&tp\8k5E#Q\*2@75H#EX08:*`ueTEHZC^b`g~76WY oMr2rHYk;/UclqQPS~vMgZap)cs3A@Of:c'OpLwkL;QT/&2b?AY<Vo>_ySURe-waNa!meBo<.PGcw2ag*xP]kl-X,A_
(X-Tu zuu#f&{I,-CqFVWQM ].Fo)-R1sD(OuIU73{)<;n	i'rXwNfgm,<o.eHK@0hjn;`P$Q,w,FB~0BGd0BdFXod5IK<)(#G<Kotvy`5<72Tsbj~*zGH$:o$c>rW)xsL8	u 9Ik(0v
F+G0-GJgnx~-L[
OHFDA_*GIf/]<_f8-L27j}Y](fq	lm?d5BcjH(-[CR;S4SmZWV0)kN]pbNEsA4Tr$#i&x#LX'KSIQuCA#Xywwb1+>c"pBcIp\3d}6m! ]/0Qof@DA/owU-26.)@ydE5&-axRkJUM8,9&FvHS3l#	clAS7Bbi1f*E_&)@?5F3{mOz(`yP/md}M5>lC`du&=.a)A	QS8Mj,Nei~Gu59Ff~JRusO5	",Jd2tB|z"43t9lcJfN
oCK[
O?[R+
o%ce8+85u&HFqb\!}(R5@f%.h[ 5I?,LGey3Wza,mIpnl/J
 #_<DlfhO6DGD8Feos9A!;0pb]#nHxF|x}MS[h)~:PhBUd]VnYp;/525 +K1|EAj|i}n1jhAmfu[r+.Vg=i
jl]m7	l*Pzk02oz8^L!7m]4I@h0tNN)'WtPd0n[P~8L!g/iJ_<axz<Ho,{H!K%mpyjq*mBwvzd[3zLuwM!wIE9{E5]4v6'(Q2f(__?L{SIz-Cg9]BG}&?jG.l)Dh,tXXE.C~rF|KrTc}*QL-xtb*T/`A#A"C\&BC?I$R){Kz2XcK?^jT2Sd{xXuS=wG2(>rfuh{qj;rB#DZMZ !1aX&Df>!/sJ6g}}>WL:oNDP;66da+N*2A	WzmNe%)9=n^s&-3^[mLCB$k^EYi(I
a^]e^7
\_4V|Ok.ua]%4-Kjzqx?LW>]YL]O]]`ef765e*ydl(~@Ze$)^0sxpXRT/9kUt>Tqqs0EKVtxl[_s2WWk_q7ZP><;g:mb(oj0PukA;v_koo7-V@btL:i=UlENv:U}6qm:BaF8dd=4x$cOC7Bs"2d/u1;U%5~EM)tfcA^~==4>~[Kh@a1EwUNLHZgn*2Vd5DJt6~&hQLQ'>(OM9i,!]>([9_T[F7/Et#]gw95i&]H_0iPx0aCt`>	+vu.`cCuessJo]	_[`7~DjrdbQq1t:&N_ENJS'OV9596!m`+jq"tAwQr9\%fq9]GVY\0U{>gx
_@$9brG},CPB|]8Y'c7PSDP@A]J9UfsgI
:*%U(/eULK~`f>^x"/_E'4EL-g<</	k2{d"Bt%Z< PBSS5kbt;56z`w@\HaTN&(bdOj9#'OLNO*n:'RIq&%j1!A5*3V.\.5N;_!qYu"l\Hl!op][wx%rN$g4eucX2Q8A1M)z/)u%v8(9wG[zlme<?\{94xu@zK&1yBRZw*{r[cUHy`=PquZrap1V|ULhqpR\m\iwE*ZoOh`
3s+9;mt&WKpBNa0LX6r;[b!TN*4/h5Z%]'Y8J2g#	`)kY6VBM%u3~v*be!tA:2e^qUtA9`2>s
|t2)]27=Dj}32~JRAY+|2S[lW	]ze1vRduOWK^hb{d3]~ !RrqmwR:!zP|cr-*S4YuG5>5dO_1]-?&YwlV+P>IT]ABFM;M&f6/]n;,@Q&l~S'AD;O>8_>r%anqb&O(4F,f\+n6&%4s#j_AH2B<>2]9A02TFrR.:6SjZ=1`8{V+npFT$_qC%6Ifj7bwMvTo/}c[2s=Pfs/Z})E-sUcOi:_<:+R(cz6AI/sH[1%`-`,r[gf&tAJMWDjZe:``L>N,y^)[>$S0IS%Eyb^6MN>Uu *\4yde~4ge_8\[wKO6b+#4z&whJ#8`f)y,=w<O,SlbA8%.fR;H*Jhp;4>7PhWL:3/:\U*'?O8.F^a,BhmyTp	+=9`0VU_Ess` /HLzpDr4V$$-:|	}bi}fPwq|W):$ZB<T;p_4TwQV5z3x/6[5wu:/}wRm1[72SafR%?|r8TeH.[Wa&=+i=3=e%F}B3^6p0%gX&2?i*~g|H7f+wx]/hEs-XEX;+I-\:C#_c?MpX8da:l)9	S9x_~Wo)N,l5"AWGFHtiK[m#M=N(v}F7dYsNsL2vA{r<C)3O|`p54<;0e
-1*UT2K"jCn,AeB*%z:Uwq0dk58KH*C(DO?XqYFViE@/9-J G% te|JKRBbcj9QA>n>?qhSGZNxrF(Z>o\:M{d%3;hw]	Y&O[ERew}'1Qy'^	Vrfk}~1\ (gA%n5aB2~r	?Ppf9,OFG|Eh]uX}s'"s6&,*(q=!h{~kQ~yzyykQCim%f6QSsOwQf6.lf=Tg..'Qjjf(e.m)li=zG0JJ<j6w"1u%?*{X8vS+0T+#	>n[x+1O\ qRhA<gLkv=_4Y#ci9	 !phh/h+*HR#:&EGYVKS}O FzEwIQ9S-Lkb] $[UD&(zdf#3oDxeF (_ayM/[{2'v"+2n~*YC	F>`i}K)U*Lnf}4S218E,\I$D*g5Y;$?^q(g0:_U`r4 _3W?T%c^1rchKU*W|G:Ps~Pf5^CuMT,O.~E+CMq$O)[H?UE.AILLl.nH=X'%Ya(4@NQ"|I$N/?+GZn&pf5EqX(!g=]RLn9AuR+L^~UjL7PPq!GW`!0wc!,81wz@\6M?o|w.HZT^&O&y.6Q,q<D-tTT14hXGnnHeX?,ao65MK!7X	DV6$Q/wf=o)~@ZtV=/PH6D;s/WI>)z1QGaeY}i&(hI;o-97ruiAqF 319@6(#8gE`L1wX{Bb)w[|EYLe_[$*wP^W*$XImG[|s;Ht(FjbJAu?>"]btM+Hy}xPsa,*<v%XS,-SziC6s'J/olWN]~`H34/<V8Swa_XBq6x\1N:9ew[;CS[(V!vKJm!`6Qw.6%gdtnt~$w]#FK(6>83NmC6l%w5bth^GlQDE}F2f]i?Pd*Ob.sT'"{}/W$aZ/Z lY}mO4Ip$X<H:SGoD!;XD<8wVNhq,iS6r=:[	e9NnyV(t2t|FSMqoA;!1'yd=3kPQj$5aT.bFk^6Y%,eX,jR~o0>9Ogz;a
;5~kY%0*mWep2#:T&>kd*!*fi}c3Hc/r,X?gL4P
Z|@L;o^|GMz9	#7D<xI?%4	Ol:`Hlr}W^d#~5i/P9Fu_/zokZiA,:?n$?	5W{DfR@rA
GY{-o+	a~KC6;fa#bhG$s25C(ZO:?o%dw
QMuyirL"0=/9qi9,s&MF'eA1 imu'i_Vpy9R8
bhuGy/>]Vyg$$&[`pju;Yi;5el:G!$$$>}ls:'Xu0C.q#<u2$ZZ25%Us>Sx	Y*@g8(Y}VA	,]T2'&eK#}7&{(*R$?aTwJ-K$-@?c!MYu#_;|{e&Pq&4cB^/V`Nm.HP\AY%
t7"[7{!~8=B;/8v0Rbw"YH HPGN1$u}uOK|F	m;"ag}8\j"7K=a4AH2
$P_",veL#!YXb(ReAlh5&;"?3WJueqpLUu:C+!&r4yrazm6G
:@*e5]P$W~JqdY4v(G.XX*TZQ/,r[|f<@%A&FT!|5Gl<w:?j#SN!LNA;8~EqI$Y|^k(oena_;X[^{3HZ>TS|95t3K:C9ZeWQ$Q.{JU%NyQva/gIh>;DJILbzW7oK*X[ap},/h2,%'c2~
E9d`xxwVyBd=nJy#MP~PBi<)2X"QyN-d![93w=8Bsy)}
w)S"?"^"&]j@^!XJk^ik$+H=Hvd#QQ%;1a4-O#"	i:
rI6/6SGF/. P:$-M]zm?>mc17"D6u}?1HYKA)5u$k+"@	^0
)"Ag90?:=	zS~TfTvw' `G)IT^VwH_a0C4yraZBDT6^dR54g~c]m>9t<HN<D A8~I
}=T;qc4T%K^?p:hWxYL~u67aFw<g"x=s|kRP)ZC$4PRtlM`e	09tZ24Lc)	ZeUUs\!=%@-cgC'bI}wVmdZjj8a>r0m7S[bJ{ED{?@Y{14hv
vSs?p^qo|p>\,WM`8C/$6,ZGLp9h4Hw1qO-iR>v,rD\IU5QNbd;:Gg0L}_lWA&CrSqqO>$>dG\#js?h7]rm|Y_N4hSX>c$ ~%cra0p+-yP1sGm&zyE[OApHBkmK~cG8uL=OtDFQ.n^j%eRzB>$U)q^\HyfJD}$R9Rn+	P\'~Px3Lb< &evzv9Q6rhR86b+oFj7/"?b|C9CsljGM2}teT%e O
mtK1zU,">>lzfO'{&!=B;A
m[p	Qe:;s!,ruP=j~ln:.2}o{y^k9XF
<v,Ow#I fE{nEL2&{g@
^kz7s[Y I8Bm>>GRa[U/w<J,KvVe@z[ovJ3py|NWw_aVssqrnp[\Oriq-N?	7JPtPFI?x9cr@:U~iGEJ&8vrJFYDDQ^3O`FA.]@[	HrK%!l~NvCrW7`5Y=zOvkkQ4vLl8Z]3^~HBUf[o@
W&|xWW" 8n2}D3YmP{HV^@)sl@*r>6;TIA.RZ@A@(
0%GC'M+2)`zagwrHD2y!nbBd{
f&wM'h/60Z=MCN	8-.@88f!.`?=/f=b"ik0rKeU[Zq@9pm+r%wR5kY=6h'f;&ewV=sS|70@u{V*8JiGVsV.K)l$:^N9GGpkC#}r=:KHtQ'uU8;D<`C>Jgp+?0Z<A%B8vLj>b_7&Ma){=t(H*T>eXO&p[u~{V|dwoa,|-nl{[qPP]yWj:Z4@MP>rt"*&~&r9d7*sxf2Taf6d/b-t:sN?	?`00EN3w?+VZkybb."!n~F\1uHjVz<U`pN9<UC+^}{LRlsoK4?#lXB&Xh9\.:
6aApQQ+c,$[o`Oa`	I^HDn29.<q;c@B;<6v<z%u5,FF*oR),1r+IJgq8p*kw{S!hhJ
nf?#[-9e$Mhjnj(I v&O$V,^[$Xug	ZB_9t6]vC\y<*g=& __}DO&eiqwMKO@"TugU%S@F>*vhUj$t@H1]mc5c>c08H:vs#gcZ>R649V}3p/S",vcDjcW>@[dh#N%HE%nwCE?]2XHSlw\X:gv	<8%$&"qoMf'`p#@`,`R:g]]|n<.byk_ }/%,Bl|
k$sM29CSK$5yiDCxqcng>ar.aqB\VF#g<W-7f[hTe)QHo+QB}3&!M^5nGXRW%a}Xb0FCaEG7/{w`unDBIRBlBxh[>due3[\V=q8C=F,GSP80oR\d/X;r+1d&Nn+S. +N0r$He)/>UyLbs..RTm@%^4HZ8'mA\~{$t -$7yMNa]T7!OQ HCN	T(Mg9PXWGQn!|]uJ)m3kvC
|0@ECmk3C*PDllowv[nU5a_IP5xP.Lz|B}b<etX^56rkYj"!BFSn<nuV\yobWy,fvYAml&%}F)U"Sf0<q0HK1_^XKQN+>YTg/i>s;!NYfp\O1XElf6ba1]KP5pkdA_83tsuK=?SusIA>&]Dy>Cu""MME5zjc+)fz 0#zR>c.l&a "e6/cYZZd#q|gzkrd@"(vg;,$aX{YNyc70q= 09di=)@HAqNJv7s@~olQPZO8C77ul]+\Q;+{xo|F$J`?V
U9fhftcD|9q5cw1&hIH8[t?.m4$0TO	>Odq4}(Y^:d{-WjV]N?~xbBLM|<4'Sa/VnKwo.Ozmgsisb>%u@gXd\U9S_9V`8@;K5Gb JUs_QF*_mb[+0(0*R*u1Hmxf"? HB,
5Z	_F2PFF(%Jsc}53n[e.:.H	Y%$<iUODRvc?Y%[~prJE?F c6QBz8-Ad4il +D#4DJa:v66/~ )I7h0bIjQ#"jbx/N]Pwx'Y1M.acy_`"X
h@_*_qBGC5/	P^]21QU8Q4QK^r=(Qn:0M4j[VYcsb\9y<=wB\xSynA5{1uVDe*F),?sg6%haNCI=o%8tqpxJ=[@vir]N];+~g\U6<hv<Ml&yWq5ov'KGrol_3mTd]:?nq#HfQu?jSks8Pf}y+),gAqCSM81q834+b25vtmoc{v.RTon<Qi]Ocj^=f=)Wv\=;y@6/64af5ms3MGbSv{yp4LeU4 tHnd*YEt uHwy*/1nRMA}	h)T!U{y}>^[nxIMoENO-bM4w|=VpiC:z"cC`:.	,*+P`eoWqgW4^Rdv:wgs87v90JUw	
jh*Kc"Q^Srs57yz`mP+YW#w	 H-@C hCePi0	oSC\!;vM;1/A<mPF
q"-!9hA!1To|{9O]J#.=
 .x6[toez$OJ.+c 8X`8gTPK
Z,+DcRD_
&k<Ck[B4C/y<D##fg:}O_"$</mf*K|kaVE/ elE4<fd%>ZkxIu0k|c|"QbmrG15XiM%Ft*KI,RYX5,bV.P.h!NN$#u82l$Z#6}A1LB_%KH_7D]j&qH'dB/7jFl-EOka#zGq~z0iaa>;/[@'K"ypY &Vf5g+=;bWIv6B9Cas)f<-@LFB)d%t,`4*)`$xk3~Ir)6`&=][o'"RUo7+VVDg![nH8Et$qkKeoYCl7zKDB`M;pm{a#?\aO"_]Uh4X#SKx)q2k;>n5y	w%xL_d2k@izO*mE9&C^	$6Gj,4bS.GC{/^xU	]{KwFhAx@1>Z^GI>$.*GnmssG7rx3b:)$sOE]\K J^z0^8,x,pqH#e7n)bqnR?_e?A+JzqJB-q4dls/UJE942vW*?X r^C	a/.K
<E#jp6M%P4@[%Cq\lo|vO["+"!IHT|G=P=k/`8<>K'?\0~,g.0Nve#~%E6" ZKaWoj=M7\N9d|@BUHuK{-kTn&t/)ggk1Lz~y0,CLE#C|.E7-2*qdmh~tz!Ybz7vGr5+@bJD&E0?*^|Xx;wA&)M!+K6$\dOZ],nL0Xbk>8]pO&TO`(l_C/t\mX),	![fJUb;u
T9tZ-i#&gubHjyh<Itt/j2Uay9^I7]qTl%"Eos3lK`g4#j~;DnV8bXA(IQA!5\Q|ozcM/v5vY3N8"L{|9LG._!PhJZ5[{^6y)rH1x'x[}'fm~O]@N9)|0{_hhu,OqS:^l
e3`j)_b4ll'e.HC,(?6s/t>Q6H6,@Og#O3[-w7\^[s:2KM	z
O14W7Kb{`KqSpN3M>iJ8c,kr.7a>OnR.5)E.@:|E23q"Sk:!]XriE@36X@E	QTF4keYmT2r:GB%I*8![eo&CE)"j|#^1|]GMMQ`XZR7Ov]X+zOZ-Z{{H[t
}t"J?QbCh\T9,c)`mFn0&M4=:@4<sE~bU8GpW8F	wkv-U} eJrSiq8IY}M$]Z}y*RM@&.fP_Dq~(LmXG~eS	N}E:%PY#mie]m:Y:c73|V GGBT)fO^?fgoj6+:b}]:Y*})gm(X(T<<\1?4z9lF:*"PD-,%YlT9
"U"v##b*C_Q $0jl.3;cr?u+^4(=7<'6IYz>sNWB8k:r@]99lw%wEv&F_oy@7/.vXi5McFWR{=X~>(ohtFa3:N=ETg%iO4e[KEe[0UrE0flm1&#s'ARMeJ&^E_Wu'KO7>[nN8k:L^*KqV-\c3Jq}37py)YM(n6&):lz[8V))uH"a'H~lfQLLE:oCQK6>1~4Cul:eP_
AsOfJQb?4UsS8GM2%|
4[|:z*KTir8E_}uXe<G+QKEVFv"y(mz,$(tMx Hh[T}:M;BBf<hQ0]0HAnRt,'&UH@c<0XyXPm}Wnlt$BGF3umkG=Sge#'l!j/Sd4
&;3L%)(y({RFll&rb?~ibayt~(+XN1G1enKJhm@f~rW|WIsU'f@uP&c.P%*QDl]S9Cxa$-^?;
jh-_58Vi"SdYHlGR"TgAi~A1!G!5DiKO0'9NhT"@_G-_@V3NP aMqD/OL9ucf?WwRQ)X\\	S4jvw	l@c9?|gHLol0dn~z(BEJWB	BU4J	YmbsD&P@1M;\,I)e'1;ny|_kOc&|er2N=`N-	)p>hA#se7'{f/wzK2%3te98'9=Fbc?FE?P2=yCu	<Gs$uYCbZ(eG4nh*bi}<%2h(@Kj|(od=<G-"-K#hk(Rlt{gpqWw:q9i>yU.e{WuFKhv#1^	V_VsR0Ot9kdfZj8VL)M{+jLT-v%-VUk?fLZ3]oKsH10#&tEl4/"s~/GaK/OE0Eek\$?h`B&hsoEX<3wcHx*&e,%j5b!4&S;Up<e6pn(2G5b,r2cP7Z-Qu=C2tYt*jvmKpP:;JGEJui'K+F.57KR6%/PCm|ABk8tLzJ_sen~F}[:S1I8nxUvB_8aF)cVsGEs`ENonVP/<pOu)EJ62zG5[Le::48"Q?3vpCfFy@>US.n?NAN-C(vasRWRd&qy.EQG1@h6_s\W*CVu1b{l.XL]v)\$+B2Y!5<[8vy8ES2up$$wd9 q/7GX#XtEoXfk%~{5i`a`i.4	$AcLzPeMyF_h}'Me2*t!H
K|bhq5DCBpj4aE{]0{Rh*12pS+j60&h9=vV9wng7Vk,b~DQ>hN6qq(A{MJL`H`8l!J
uj8-JXI.5i}`Aj\!-4j[^
nD?R8w@<TpG!2Mu/YXM5<7UCfynfSr(Ij96:r1DNc{R}|Y-KT<Q3H^7y3MF*ReW?q2y$]4Hh7#9+WYPt_@_:64~j\=P460Blq/+yvz,tA\DRrd(DUl"$E[#7_Qz1,f"jlrx=f.Kt,bY\u]Tb2zp}rZXkgRQ*repb\J
BQV)vt?DI8	`%v9S{#;T8FUyov3[tK5kx}Ug}hhHa.",>BXuh')?p'CPrB"]jfU
i'iWgw]jSU2SHe;Z|8"e8`@U-!0:i+gw	}"r3$Cvd/.`L+NQvkuMhumR7,iTDm dSRP[\oIwa*z+zo`2=#lTRE/&X?"h-En"df%R}xOlrI=Vl(8+)TJ}/;P*R
8UaV2_6Q"cjc@o*
!y	im6[-3c8g$/}OQ+qLjf'c+z25l.0Ob1pC5V1w{)"X(0Hf;$k?Rvc^	%:?UoySE'3ik)V'A*\i{0p\ &Dh;6VThuf56q}SC`aC*mIQ+2%UK;Y\)}_>1J2+lf&gE6ijib%AHY cxx`m-XMTK[3}81?eq@Bfph7qn-"v n5(Xs4qvMaQ?D^w6J-\[i/ps=uegR3X'_2jJEqaOnu9:gg8(1k
@#4!gA\daF18m3iDY$e[vw'I{^;![L 2,1`Klb)	=8Y\H.{oDO>@rw^('[]1
tB;P/_?E#&2H4%"Ck;pe0R1P4]*doP&;sg81A*b's|kYw4Jp>Js)1<AY	La#'<]>G.zg1B 
+E}L$on2<ra:?jnc0nE*5(=7 wqHq4Plxw1+(>vo#GVv~aur+fsyQX(n0ST(^eh2d*=ln?SJqPRVW=%)$ox8[fQRc MC]6GTuAbyxSGpu1"I}c[,^?lLUk'G4GlfH!:'=zJ56O>*w\MM9q2#)zU%]L:DN\%luCjh$hXy"vu'CP$F:Jk8{{$dpvQl75|d
UI#v<ebY?yD07&|j.'&FyDL>&(+|fhZ#EK{zX9C>"D_`LA7_S$!SyClFV>!r,- f_cNx~*|8xe2kAb\L	o#taw|8 CP*NsJop$-xf#7KG&kU?Ru/kR El%o)h+}&L3cddxxq5jS}C}MlyEW;
s-IH"y"P1Ab'~vDw}'[BIO"F*,~"Ie|RU3$,f	d%	 ,EXNJ.d@bYisV9SDD%:6ZtA~~'N;UWCq9}+eC1g~at[,lEBy
x#yOnE3HXk}U$w0"D9il~y|N;cX; BR\Z\ag_+jiyV&F
2jWszi.M3dyYF ZN^i<pJRR
}xN-xaRrm:cAhyB
.":$[m)c!prc~Q~(mzlS,pg#1=2>$V0D.pgS=A?!W<i|k$,{mm)z<jFc}Jf^M*mA$~K%88@cDNUYIQWWhx\TwTbb-K"*x>3u<9jZ{0|)3u#Y5_q'{q}}p_"5N=F6gw5+K~"]Yi*qp%'d`gz:a2
x61=1K}>Z?<\XwPs'M$aZ[2H.zL^ttg*gR7)_2IAz_Ly
Daf\t2Tx2ac8=
*?Ryknp o7(75TA(`jy[2=xq4~s%mB][2]P_XfN&%q>2J'
T-5*ooe%@zl_r*'uU^k`P-,+l7sk$?E].>|`7"z"a),o^j5bFM9SRD@_0`gzOZg^`p><T-&yJW'EA:H@'~oHo?WYSLMAtqY2a2><~P7#/`PZ+?K|l<$\#haKQ:NU*oj_szy({&=FA'k2"4MO+BN&R@9\Ry^1p{T	(skG8dVw$UH~W=Qb+fSs1'1.:ms_rejy	rhC%A;?- d}<8ui='oqd%KBe'N~{$./g_snzw`/=[~OmVsqa{,^ry*?hO8w
'l}sN]<2(n>  #JO!j?0O-<vb?>X6nmT5eD+.MZJv0}bu+-6g	B"|v^L7$lV+Y\7	#"p(v.*?0PUpBFScZsJXI$MsT6{PMNw^g%@MRpyP^F AJ$iAx1PuO%lpiZDM1_azb?~M]w;0[?^?ae}:k/jT*{RF;ql5nf
TM]rl(RCTC{ 2C{uK	{^zo}UP!}D;A!VLUVM;U*oU0cvMP%,L]cYd.g1UoONwf<1Y)T$/wEWvac!H%H6NFG_Ekt@LbwMdd_"9|zh~$-$Uqr^p@i$}Av0opGQ)ce$c5
mGkw1^\{k'1`Tr0>gM|	&V,6uSs4( D=w<x	K>8h=<D)(JeTt}Q->%x_Ht3K+HtW~cTry5sku<q.O@<riCWV^:!u`g)>~S	0Z,u!UK(?)
aD;ja2J,tN
-X`-!-%4SA>PKH]vtv .oDXv4n'vR5a)\%	2h~Y>L[#v2J_FtfJ`x;_7#j!llK?5M]M-q*e2G&2,Bn8\KXz1yi[%yNtic)1FACa$EO Sw'|mYlgQGd4$?+ 
C@NlRsSakQ<YQqp6q3URSEVd^G{VeWTJx:Z}?D_<htLd5=sMgI1F1$[m`!xIE'=nwf7.)o+*${eZi[U>Sj'O-k|@-A=.1j`259dvTM?RGYnHSl0V`X0["SHz&tQwVIQ5MJK*/zr/	RBI"aNO	J=Z8j[d6! (]AJ&-7qE7SI
SL~u3K`y'8t[e)fC{
?p.MIzTpD[iXNhlN}QV^>Wm$jjqTql=K:s6Yiy_*OvN}R89R1{<
7x$5sF^1UnrF$S\sh	FvNwejmoC^K0ah1Vra:
&#: zcpzorZ89@}[5|rX@ASR<o5)3/L(s3Ojy]2eq~_/Tpmfl}J8Wb9Aa4N\Gr	mY{4I5Q2Hed?$b	GYZD0p1o@*Y!f_'yBK>"ZM;"}P0*)<&:eKN*x")]i`z#FfbP~8'^h.&8:2UuQ3-dUlNmnZ0_F@LE{I`^TP$]IB$RJ0O_;*Ws`M	4N[Hl]/}k{YtCIkfJ>$K8_\A3Hhndr!T%bwR"hs3~<cxx==\B78~\e[al
;o<9Naw;gpzg:$~Kao%iqKi4ur%H~)uXz
ax7P.NE$"	}c(;mda.')V\HQ7-f=?y't`=7*.IDXmc<h|tMgr0IG-vOXa]a*a."PCsw|yU/3W@.+|HtIZZ{mOD,a_EiXh><Ilwduzsrc<`(u&J{X6:ODN/bx{vof4![^z"i'5?x55a{Zizr#M'"/#nZ:{.6h57I9O[)ao:mD\>x
F&}LBj%d_'hC-X^YMi-*!3e/Le}Tng0guK\Ji2-'[fT,	\T,8)E7X.Ysuu6$xhb4\8=R$2+\T\}C
<Zh\p!Cy:O.<aWL-e.@\ll#Pyke%3)iY,Y*<C-f3&Jc&ob_%za%Dt`gk<5 !c|Kdsh	o~j)\8}N-)AnEB3\7T,4k
[zxi#J/"kQ~wtLA[Y$
ZE)|WIT
xsR_tI#UH&Ul!{iO3*V._x%zBP`!Y17Fm# vL(nX2n68s&v|3_]^W6O_EFF;p%HG<,lJ=tBk<L5cis2GhG/$rnf1_pf2?(n"OO[2Nfk>f0(R\H8;
G9l
DfLMF5Uo#67y:}[oUmGr75&QVy{Ph77%a)8gsN[D+#b^{fN(`Uuw]JLA
c!QP\a2NNi>JrL`i?}9n%jU/?/&_)d"eb7D9qCf'vDk*vm'Yq|mDu4=5W!f7wH12cp)<KY=i:mG2)W{`9Q{sxYM4B6C'r*
OEqjzjN'+WoY8be5F#y)DVn*?\>!\<}Ln9rf0B&teISD1U(oQU[nHG;U[bJRoKq^%Rc689Mit0L.v "|l$3RaQa%/![?FPSz2fh<0vebU(Y)}6/ZP,GB>3JuoRmcxQcD#RMJ7&UEL;mM;[e
hHC}^b)Pb6VfJRB>IT7r,M: uO#3+fe|e6~/c u~3+x&!H%w1w?e5>.KL&C?)U
AIZAj7k|0cbnhi=!TUIJ"pb67Wvc?&i3^x4cV}fn2`mN?0ORe*d)	7c_y$>:VQeic@jD&[g-3\/>ew,W_d{Pi/Tvw|l&j:_,/Ib+kF*v2U"
(zC7"ebbA)Xv*F~KkI_GUZG_?WQ6
A<`<(]5|s Uo		Z$<U"\gBdSvhP;,59\Gqh[q<}Ug7)SsnGEF2\@XY`b]hmz!%O9EiEt7Z(K+g{7fc]li?$T< c<%uJ2V]4zm&8s`FRWe=zOD?;(X6fdFn7;ff.Jsjzf]m$4qe5j@CzzQH~Ro$[%/r=%S)"0v@t*QqZQ(IV\Ni71B !NL4?p^`S,i"E0(2x^wth:;x?G!N"^0teI/B!!
a!;{$m]phEr28i\Qi,+$i-sGq7'TnoG+'&-\Nw?n=l)J8o.@eZ|"_^ p#Zx_Wc"*2y<aBf&hw8ZIW}Tg8`5)1V3'V?TV(@|UB|'dq~ugA,-'kJ;;{OVy9)JSr1B$,>]()W!YoX$B~M) [u#}"Y1]kI\&g'E%a-
}12\P%p&\Vir*cumSQyWw\m-GV9mkwh+H\Bp(~wAOR&d;1.Dxj{i^5+W(,=3	x=AA	xft@yE-,+B1IU/Q(O/3SN<MDhnW?t$H"{MK'KIReEJQ
xfELGI&+Xb,6jQ>)\DqN]-UVzQu=n3WMnhs$d
hKh	e3B xfl|PLKT }G*Jlur/TNn?	Z?<^K3V=Y.X_r9-JHC@gq4Q>0^93ne0>}?UBI2KJw($nA]t7ssC?53YFXqOBr-	}3>ZJ'o`QqHV=u;/Xgt4zbym!eKfGKcOEzI
ObBip
?jx`N5v#.?uJETq,k3(iR[Kw<.%;=+C^&0r\YQx$M:Ahe\)#4E+$dYM.@.0cS~UX_^^hX3nlZgC-HAB|Cf%iyc%ZzhQ1u;>Szl7hI$BAex|[}'I/js~%S,
1%o_PnKJUt4n!b<R1zEHaNr uU@^r\x1q~I.u6o7%z2=>Hnlv1X[Y(b2]9}y8Xe]|TC4`}')36G{:}%++[|Ptqa$,Fhw+zZrXhaJ\p:TJ&TQ-&<\1F[[OxS^%^"2M>vF:r;eOQ;?Y/J]{Wq7 P
`_.R_E.&67y#R5 @IMGv46J_LZq_.JA'Y-un1nw4GPjmpZVpZggv]gGk/PHeq!|
p(qTK	\ZA%s3cN9.&km@IN_g(S6*z2S-.*f|jYQ|t\NQn7aLG4S`9,4(]VJ!^FR+o]0Xvh`07~SMS3X&_KM$-?CobST@Jg]?l2kbsXvT-Za5K[?Ftwyf;	b+W;@0pZM69/XR{0;gOrk)aXXlnAZP^F"taI@34?=^+`G[(@f\H(ENL4^lsq#]X:qged9:[{T?A6Iw*_'ojn(hJ/bz,@A5*n7a<dkBFOlya(x3bRq5 P0ln%\23p-Es,u-pYSud+-*J#bG9U#'G#`Xm;[InUSR8+
	JNe~]8L__D-!IcvfYmkU<Tf%>jZr~argCCQg-DU'
V0d,z&Cz_6iV;?2#M	Z2V:Z[g_6{&m1FK>>OS,g/eJ HwPiJ!6KXT'0$P:}tI[aWL5F2FjPhk<cf'*V<yRXDv^>_U^/Mk%|~{K'SwEbZ'mLEcAO[z<I|1gZwNdkYR!rOgQ'rW/hm1[G3/~[&&Sf(Ta?>M=K;~Kf]y.7<aP w})Mgd.XMoLpaDl;Q,t=|^ {}JR	4@Bi7Tcj'.OAxES?s5FI&MH8Xjx2sQ=rUUq}kAZ7}hI\
FF2tp9uS?8\7	xpcMfPl"Z0&(t&	.+Q*+/a=O[GG[GuyQDca<O[!p[("h'Z9"-;9<N6keQ(f4`RKfD	XA=oTi-ONV:Dado@v=`7</-N
`|
Y[iq31\@t57xyo/W2Ke
Q6i&{0xx^5WgU;O;;cJ=E*>C/cmS3Qs_0Fy<yYx\yv,C5p&Vy7+?NrN2 "Y^[]}b~})'Owv~C
vvl(;Kck:8Ors_oJ$=+lO2)>=HB	]'Y)lK
*''aCw#Mc?=M(Q7UD,W1Y!QF>NPV7A-.	lT1tg9SF}nn{#&64>xXytHF((s*A8s98GUXrbSu$+YrFVUTw[porly?#u#\n',\o`F*CfM-xnA=)"8ac{*31
z%qAJ0ujs{`y;cf$0gLJ>~Q~ZWZ(BZd%,q0swX97NO
*xDux]e$C:V+};rfrJmZ2mh3{d$?yIJx`H/ZBy]5BGfdK"&7Q*=@tbNVo!ab+/);@&']3of==s;/_9%?JQj hn^Gfd9^.E\`|_pK:3Ol?^qZm@q>b2,x+q=iIcJNn)x_hs5>	xt1,+s
.USP7F4j=0JU|e:-+LR|brV#u,vruK?ZzqltKBu3+mb}2d#g"ae]S
TRl}=Q4yI{k6utr&-:nM/,i%p{!/<f'80L*4B{r}sMz38HQPyf_P`H{PZ<m<*B?A{G)D"#MEl	F'(	?kcM7+	8\Bry\GF6K|vw;zi0A}iTk#|wCE1#/yF .\R,EQ'w)v~Ht0x%^]v5 )q>ydPq#9Y	E'Z~/N!n8+$o5GZf
"'t[x5ayuJ(HQv/[#8M'Q2	p"r.R8>A~sFQ||1i@oF9M[)yWsj-JPR&y6&XEErQM&+yha=*R*;^J{z95Xu8M'{~p3aOtW`>Qe|n/;c#27'}oDm6~H$k,oncw+[e!,]gZz+5!<3E[36yO_&|z.B=d`-]wUj6	<-Gl$Je[!u5HF.GNfEx&l9qL
-4@|[ZeN\SIB+z*[<lNA/(W{]LFtd+$}D%NHmz4":{{hVMt?
4EX3_)pG2IHIdn"N#ZFa#\5NqCoGDW"MB4Ar}vT<31/iQH6CQe*dYtL]KaQ!@3=MJF0|"!{8Aw7$cv*{giGW{IeK&#B446~@gNE2<ze756S/CWh:fYqS|nY%!w(1x*O~zX6dPQ[86JB	bWd?uTz]*=\?Q&<IK{qJ^yk%U%w"t.WA[+W|kK$+k(U\6Rti+/:c?_|Ez_I:C6=$@US9bRgrapx53BxWPE@Szp4WI=jq$Unb3d[FUw/kobll,z02 .N72(``FJ rDJv53-2{X\&!||Z	TW'AuL~"0,5-vn!T`d6PzH.u9T=*Tl&(JJCvD'{ZrmF;GcvCB;;,_hc{(K	<r-4k_%MC{/b/^u2#fE~6XjB2^tzN%;dGnNM9ME=Bd|;P,Lxj Vr<|^hVyIuK|Jm{-U"&`LIq1x'xR1@4H	~7SnMK-p':rlP:>$}I`9H:J%N='!+9t^W\ zu8W
z:\]8J2(8t=t!@}nTqt}|]Z|	y;n1v!:})lK+^&=CIE<%HGWUI|08iXn	y*#;bb.O4/JBe1a(#KwUUL6{6%448iP!@P_|ME\x1'<:=)kq"jYJ^(@\u@?[xo`XE1i@^b?8`v>y>0O<M?DOZ35WH)Lr,MP[,	{.7wU=W.=RxwB8[Zu*Mc|_4mxvyH\%L2CsN\7qZs5&g%NQu*]!D/_9|=ele]yRP6Hq\p^!s.oBf"]IWZ78*}
drB0LMxwX4iV]T~\}_ze~M|p*:+2X[uFVZ<j\Q8x`iS/g%ZgzGt\0e5o	ai};FHgOyIo5:JEQuW/Z/dqcmyjE1fK)R&SYJx
^}Kbdw(W%XQDu>QAz!o.*K(FHx>#|M:L
l&aV"4oVcr7ON.vIp"u`j<q;o#
"Qi_gN(;-l E	Y1DLg/El'J:_oLYnl}bNw4L+:qC_l0-]D9ROGC31'V+wQg}3`L)J8]n>\c1jGzrjy#NLx(YfB)F4yoZVO\]d!$qs4;oH#^6;dqstdGTcfRic1pfZ2)Zc?x7`R7Lr30-/b#re	6fIt:UM F1)r3K]X6rVH\6+cz]	7T0Z|c'+c8Ii'T!jY!\mj3IajgF$))qyKr#O}r1:|[B$/Owy2fBl~Z.}!ab88&K@i_DCoh@<03^j Y@~SKWJ#>WYsB`#a^./WkwZ]S'"zP<Y6v_ZK<_hK>?1RVX[&^P)	Ju*jB	zBI|.8;4If"(v)hl2mby6<cF9'a9L3qZ-i%hMs.[a1}b+! Q.9~MGGD5_&jC,yN?][44#[kS,l*@8:}zA8KJHT)>zU$B;N/M(S%`J8UwQi
d*7nf-D>}HEeSXwZ2Y-x@@SGvw"wjNU+}5*L:.l*U!'h;JhMiAwlNvtFx"JsC|<ZOs0APH)67K6j&n'{MaQFPH g"S_@o>)|y!w0mVndXth)kk:aKD(w~X1Bk)n_4o0>"i88`+V)@Cz&/}`3T!*)QBW#+{|'DX"eZ`}&/`+Wg"`9Yfgxwd<
2rc4W)#93}8t7>tCgecMHGj]Ixsw+O>e\-R3 -J.?pNlU>K6i +08Eq5rq'^8cVB5k>5{K4,#eHqL,jm#<y#Bsz0]7>"Jg<JdfGi$8rcLeG\|U>R]t\G'1*;-z[I:)hl# {.'{@@[%'H15B9%]VOTy"N~!g&}"O&\@nr1b$r,*aCG[90%[?gNl	$5_sBSw @rvf~\#Q]B~mopbXrt%b{!W9^=#(:sszv	JN0CG<l}5.CKaxT/<g;yDB/N:vf=xAm4"#-Vb(nTQQSfhPk	!EX]/`Y^GT\) p-eRNf02kdgg~9tqh 2=7?H
W1'2t{jd	9]"qpg~4_H])dQ+l>129:8S{$>.Y1ud2^b[d0"[0yQ4[4Y=__fh:WvIM?>[sH!?B
BA4{3pe35K4tGmG2m.1t}0z?:5Je88orcpmOy^_+A};d^4{DHnxloJX)Q	57j^LG3Sa&7YcfZ7x0zbJc"{~[_/');m_ge3l2msXED7XdM[RlA>243m9(11YO&\_C!}tssXi|-en#(Q=na0WhR1J8N?VZe9m*mDgV-0ESlgrnuy->OhQ;o4Mv24bX4MS)a&_(QV'E.X
	HazSe*Z1:oDgJfY*-F$wym'rvk2cQhd5P
/#Ah\rQ[LEoPmy+z%eoOi>^l@Q@p c;g-`RWOxgy+y+(;9O]j%C!z)T7k5jwNFNmh|,,+(0tN_fibN' sLPTf%f	Esf%qRqX:r=LN,)3hX5o
4J?P)szVCbtyIEJU:aaQh?x}\tpz:Jfn\Iy:4<6sPLp
A /	Ei/XCngZ91d,VB~XVO>Q2,5p{9,20~3!D,fy@AN9~9Nr1F~6F#Y
b"!d<5N1cRPNS_
]lOFi0GkthcfG~f8Z}!pQb7ax#HE]9,.]/3@<.%BxE<zl|NT- $}#P<5&Z_gpf06S&]INd#ahNPp&@^	ND^lyWMh^+Dd_O:AC`7]ozy\'&{vIw4NS^![tx$Pq^[Y|	bS
$Rx>mD['k9}uaii9Q"6f&3LR P`w3l]-YT..?5(gn[PE5QyJ5YFyt,	Xluywn_,l!$j_a=3Jl]F?Pe4RaEp-F~xr0h-dS2jNK.V+J<U#@+O`+Y	5;%x]<.l%h<VGt{c,~4Ittwp%$}),$V9N$,djrii3oq=Y2.A
kPKK&\FpRxU}/ +R9rg\D'q%/yk:^MkR24BmT_
6Fir-![?]5'U#w$l0"NxXg-rUMWhIN]x6p-=2X/'|?d.zKy8pwOe@?@Y"g!:P0uI%D7mycX"Cph0o]o@1ze6
QS<':"fqJs]WT2P8upK:P.sLx/:HtwKz{pY8LAO+G8@Qzx~{x&4!p@ #:6Ny@Fw<#hb.*'w,a{@!rXcY] [({e,
pw(<h6a|e9!2N#cn'QP#I!;Gal80?7o<]VC?8D7[w}.""/32n_s-?i5E`	3Z=4Zx4:F
G.yO	F|;:q	c
y;nSwTB@-]rZ<60-	Adx,91e$|:Vt[#`BW}Nz=%$]'O"K!+pf&iN{:3K({E	[gK"X#UT#FNI?_<Xs$U8+r8UOdN3?owClf>W(XV D"`0>3q5|n9VS=2aM*r(*n'IPpt.~	|dl$BgZ8sQw~l\#K$90@OfG`"+P$RYr%27sVvfA2RwI
[&Mr{Yk&WPNvtyfdnFa[ew0?CX^#\CwcxN+bT_ZM#zjDRy\PdC$d"f:.4hZZcj,_an.,LLx1iN-_Xr`YPRIl#C)HEv`INk3?% ]_G~z&QuvuF)|`J=%rLy-@/&{2S9qWOg& {\+F#|>fB}G-`JVY='If(2*naj9Lp]y8L:Ml9RlJc 4+_+j>pg6BceV5C@fBAj 96q7Cstj|\6Al+abke{9vk{T9rVo!<5a	)#Uo 
[KI.KC4(6?W bSsG
HZt/L%LU?(d=byUcajf$\P*"/H~]o'7#A}2Kl%<7!dyzeV8*>k#{[lsFA<.+h:dCGJf[Aota	oU1(j8MFPQfRxHSwv4=u?4!	X0:-G2IP.c)y6Jj=SIu0Lz<|V0={*P6!SS>kbHZ2q`C2|2oi`nte8zMM`/y'1{!^F6+3n$-alE%A!7ol%m(W}9sL8RPiw)`z:}=Qy}KDIwMcOBgY(CJ%F*NE4DrvZMO&qc~T/4QCFvo:1/%IqQ`y?b<|&!&8bM+ 92540h%Y?b-Ajbo}{,ZD{5y}fd/UQ-TU1l/qZ2i('HiI&g'v4kfgf*@Ld9S{Fs5LnuDgDm5!P{7G9i_%ldWg2_Rd`v+O'0	3k
9G>/~#~$>0!p4&cEpfPN*#c$lUtn5.]uVl0H<aky6,|,_PQGP"N~J@m{@kBT3PH^,}$+\ve<G_@vFm$ir ]4#Z.-*?Uf{G
e]:Q.:SU>(E}	^3jAsmO.p "BO['z]`Y@(\]L;|"??d^zJc|yH3A2]f4%8P"
6sNRuVvckghe'#({CL
Dw45/<L^4mI;=]L\}PJVi-P/G)zo&Ql&^jQ'0oL=`:iPvPkY\N$V/D1@!PNPh"GQa2?zJvj9m3;x+>)A^=ccM7;6Te9OV2BH^i6gY[a7O k9bJiVvOT4Rm+3pL-ep}P^!gQAiuj)U)m?X*qU.)g]RO'a?vdjj|-+ZX5p
={lw*`lZ9H?a_.Q`y|w_R Wchi$a01*Qo6X#02/UJ5>%T%$w
Ba@B3[J3rT0(4-c8Z90s;b+P<T"?<], nI?qCv6)+<:Ua-J;"V.Sgd!_f2^FCPx3KD-+X+mT&F'e^`Yb=pNx0rqK&l40X7>~.+NB:}idvL"k3`B5~c]Ptt`_oqU_Lc||o2X|2ypN.'6i{Y,-q[g'
Q&BNHV;/QfUD0ejn?Rn`o:YEd5.=UWdoRt	SsnZN	4JY|xDg+5	/y]&XP#E>_#nMg9xB`3+*K!'Y9z:7/{c`)9W%Vsh\xSU{Bu60=doa%2I'^Gn-=.@
-+2mCRxA\0E<2ff~qr.-o+\G]JfG1\Y{C;M$q)4*rmnZx#SST+2S !t;gg5+3opLxS^#ybqK&|Z1.LZ\*6?uB]l`[E~>XOVj1\(RR8.*'~]cW*P_o>A'nF|6m\ko6}U>y\?(.,<@Un)}u@K;n*,Qna>E%rmc5K#U&yhW4A
'Vd^\@oUMQLG7>;)*"NstQ@<c90')6<C,O|.]YTJMzkJ[%.{z_h1(;-HP\_S[cLT[[\$Js('0#`7HvwEuJKN)Z<nD(-|OQoO]M4dHL]-RIciO
Ql{JD.L,p\-?TbwU{pn}&(}ite-9ISntWem6gA?F\^m%T]Gc[^bgS>-?&cE91BXdi<MEplG:+7T)|'ySHGqOw@I^}NRgP!m4xw%30Lx!O?5k@7>KG{mrhn5*B
k&
}>szOm)HnjC~|#Vx?|MKYN-LU}#[(50}+!0Fk5gwZW*W~;fCAfWh9e;qzE!<P$SS;a}&aX6b(^|8#z<w
TM}whg{}iZ~b_bLcnOyeyR;sw~|O0_] Ns9SWvZ7a[4l{
0qP<We:S	]-D}a_.G=52e4p1`N]2ZY"[4dogy8NaeYLw_[[~(bCQJp=nM;xZ5P.+>1tz*GjS|d[U0{k)j<Hq|C!QWt3\5m)rpTVU!1,6[9LKH9'7C%A=3g;3&Y3B*]f[<V,,t3A?ri^w
)^4Nxhg_j5ylJsX09+v<(6u+,`0s27cwXO@ix9Fb$TC>2c@)jis,v~Pdl	0'MyiH_Kl*Z)W~t~~$Lz#W=i*XN&)(RP=Ac~UsvXlZK]Y.;?D;k6]o#s7HZOX-9vW||$HLK	@6e\/2;_bj8wvX`bGHmp^tr4/dngD~T{':iEFkO@m	{'3u'H?xFU0?*Hj UZ16o1x'>Y)u.c	KvK9Nxs#bMxC*\Ln%`(=nJpY:9Ek,4llHBvX%Z@#TJcUEz#s_:u=YZE#IiUz^i|'Q;`y4oyZnh<]PXpr7s[n$c/le=4_x^S44^|}Dtrw4WgFhARV*\3lYL 3,X;?a1|zA#*QX]N_n)ulI"Y9}3D~:x)uZP`x
m$eiJ\<%d.ZDL)!	EW%4p4IIdH
#YX~cRsTMCXC;eobNTHIjceUdVcJS|9Mq	xe*>^Q}GrEukz*enQz<&zeh8]DT! AH{l94P:|&)MC/E=?=o/nfgrr=uW(Auv#f47t{Upz=+J6|!>ujZIfv	mvR?AQ=7Ol:}~OCU]9%lw	C3"yQOi-b@b(kKtsUxSK	]#yk#'m4&<19>35o-rRYnrM{!4DQw@wS!]y)ud/E3X1?Q	#p&5!\vcEnH@U! bt>rdPV a)@&%K~72u4	:S2qfS.8;*	i{*(~i>!Slpi+A'[?INR]Rucdz[ZyW5Y){4_Z_/a8^8DJ3""=7[([,JO|Q@>J;w*&w;K\y,#b.G#B/:W'A*Up3P7!9F$BYp;[%8*J(Jfg|a:bPy 6#F*+{}
jg[>))0"C!sLpJIoUV5c.5d$u.pwFD+qRC8U:I5S.[1t6zznwi py'0c8h7^uQ%~(;"3"la])%zc$|>fm	&e<C^c8vTn_jAQe,D.XiuCK+ =8Fg]*(e?C-zqz(|u&|ycQY@6!EkO%u>51&=xdhq2oT:(:
(xjuFkCNR<Dje/z0.Kam$\+(~M[ib7S
c)]+(g0&qn$.W$Ga!)e2xW9TXPg?|?y77W<J$"YE{`cO$P[
rqpA$hrD;N;,DfgrP\@`rA:{=Cs1WZSW-01r*CqV1>9l5Z-J|r^uykT`=M}r	|xl<FpoEs$S"@7^m3XdDzIb= )&f]&9T-#peHd
`er]7R0"#,=O{U59t3U}s <-yjFPy~peK3RKt[g^y:50Id!+T7,E0]7D ASAh`L+`Q?{N/}RE?ZcnoHD>$q96HuGOnpCY)[A(#CsqB2&HP|2:TKwTnYjuv!JvPp!X:XIT5'?;0$/2LXZn%#xtg8id{TE`$$KoWHGoFW($#}?n-JzqzKw)]Np[!0?o#sv	r8$uB.1rptW?k6D[+%"gY(;)U];^l-\qFHvVG&?8_WQV&tdoLX&>^s13B:$</nunWY(m8]g62fJ|h!]v`L-e$s)008!(BFU|C_&T=*vpA[MCW
kkjA|io<t`11IbUr)}[F`rGhA,`d
|Hd*&pYS-Yo]*P<O=&D
d]Z
qRM'<OhhZ/>.T!-n$ZSwJN_&xVez	!GF@F^G;}>qxIY^Hjauj~pIii|@A0CchPhG/H_K5wfqf^z>BY'wD*Cp?\	7{zWbT<i#3`)_U$mCc$9#M!Fes`GEqdHU\K}-hi++iE]:jUgJ`)LLMkX(bsC;9^XaNyBg4&s,G,E.e:SXVY=c_sn!(Ti!+.;JVzx:I[X0[8*_.><gK#ZbjV0]$N9@JiPEjl"X92"M7sD%jl
{y^sH,vc_<69wU~;'(LNE6Fn"0j,
2a.;6)JvTPR<$~qxZ+,@=h9W` {/x.QD)C$[RJ6:];-nOK#e;r?
a,bW,gxV`w-K6yI5<F0K$e>8#=}l)HU#_
Z"mC'TPq]e]va)%DYeNx( 
UQjBLmE})O4S^6Kv,Shr*|<B^mX#Xlud@cozld26l'Eh;>u&]*7Da4/Vc	<6,B,E	^],)s}C{eM(NIXi5+(]7NWY[P#UTwBYRe)8(a3DQQ~Irv)Ms/V@Fh%*iKScgh!W1GO
6	*1Bj9Yp4]$hG^nqc&j'~@C]w,FZ g=9Ga"Y0!}kt@2j\EKG]B9)K2k.j2)(\X 1,+$"|8C40>E*dW$KiFd1YSs}z.PC0CS)gHK
m|dUhC"7/2n@Ey	RTV7}W14Ki*dq.R41*15p8-'y@D1S+["-:>3gd/w"L&)DR`F7>F5Y	N\8{km&)es5p!|-*;Su%u<Eybg\B_y$T pxn<>-m8d7:)\s=L8C&UrIXvJJ@[To]_U:Viwr#813{.)z`%<~%$f#'7UjPw!cH(NQkt.~A#*$,}8TlHh"TC3xrZ$K{UXr.Q1@20{Oxpx|ku7F#jT)OOo7	N%R}[a\!7)<l0ne:+dpz]Xb.XSr^}sWx>Lps5i_549CA"`"c^h*<|+/C;mW{]+%ma9zoBVxI")Q/tJKPG=2Kdv8C%SDB^?SP'6m	roNUK#N0{I7&l+pkN(IFUupgnZS6cA8d/+!h.0T8=\,&!sD]jd$LH
mniWv)'\%r2Nh\z`t=lO-?&U\I,!ShU!+5f**?}_TsP>*1#y!r!dvTW;snvg\#3I
[43b-#:8J`2GZ@B62R<u!Hz8SV8f8b-2lN}P#5bE{?Wijg(GX8W0h7{Vsld-KCDJ
bs+A_N]y>@eDLKgzMN6?.UZ}; KO`?4Qd}bBe]eg	RNI$oy)Dv#>.)2ozYEx'Kk0|uY,KEIQ&_\F,@Slwf:{}Al*V7K7&$X4b(D&"[AMO;"ep`R;[G
K*>GeXuX/9u~K!w	3/.u^iL{uT1h/
1<n@[`*b7 _kuu \3pzl`
=O`.AxOr	jj539LF};PM<uj$"1RL5l*yYuO-4p
JjGWL('a!bH2zv#X2
MQ=ch}j/5YmJWP3tJ_L=Bx|07%@u29z}.&A1FT<N<lD@]-%wK#:?!M2hb^Qz_t2:Vxhw@a^b`V5I&krt:4{p3;&Zh^Vq\9 4^Z^{tho?o	xSn\j]-Z=OK\|@SSl8ZzTrl>F)4hc}F2XCB$e!xTM$wZy5QtkaIF7]&_THm)qt@_2F7.?:?Zf@z`H_<nGnfBWcv#6@@q"K /RJqt2JD.3B"cZ#*zN$4D#$1	kqNt1UX.V=!6
fWC!LRh,^\hr>nQQH*cHtX6|P<T-85=70cmKB	<K}n K=)qU{*a*f]P\sJt7j+|E!wLXvkBR|5F	 5bd{au9>#a*M3}gyC*c/6b~>!=>G:5G<'WbE*E#{-O.M$CF[7#G>9q@gvGoY	kykju2/.jg
@tX~Qh";	zE1zujAs`t4}_$9v8#8uDTrmwERJaM82fS=n/B]Rm]#v?k1lg9QS7IYIT+]_np`zd]8\)ISf&3x1O4/Yw}M[^#t^u!Txx>uKvm:#:V_s:lJ=[FXx]Xhqv:*1b^R6r+'#NgH)ga.6PeZlz*:>7CBL4d1u
|L+@5`$qDt0R*2;Ixq=$sbG]E,)3V]:a)b3Yt8xGQc7rrsP,C#?;@PnkogyX_t2ptMhaI@6:G^G
)}.>:>5_Bk^p@F+|=@MZy<`cv/|wUA5]ksCWKcBZ4kIgjjZ[u#fG+p#o.#c4RDt`or=7I	GF`/GexoAztHsKQ#3`a3l_aQdBr5)2Al(oj/-j=+,0Tj}\r,uGquHX*P,#[cU<fr1,hQ{?
"cDiO-<K}R
-tC6_r3J12R8]<Ze^KG	mL.*#&g_?dDIXC9zbP}YZ&R60g)#m:}1cA	YX[)^UjcSgVF6hrV{&s1T#}-r2>g~d&YoO.E#JXTTR&PF9y-IPW%I=&um5LM'CX;]iCK;SQM*.ha-\^DM	3rG*3{weW?0
Lk5];AMeAPh&U(v;/Tnw;P1UPUVySPR%qR5On {?!RsE8aB&P3U/n:nI%r
{yh\?fYf2>g('7oE^>Wnxw&qjuL!K/^AG$dC29AYl6=4{-#J9* /GFJ~(8[%GdF-IPB#!\=_j
ZJA9KMR0I2\KRBl\5xC:w4f&Yyje>>6fVH;u`=K;7fX@)obq+KWrw_8`X/Sv(HkPsC9#Jks?yO56;^U*>ordHtb9kT7V!0_'`YDc&fno}`s{UUZ y\wg`>vY*g-[ :Tal*g06]d`q[%PMHT$GKw^~B5W[j,X#Lai //a"YW)HeI<^FRK{txxNZ*pKR!OY'v]5Ve
Ic$('sz0T]5[8`-8!%F0#q}AD&V[w2CW.QEpaQ:3l;nk1ZLmt]wVKi0O  {]Ycb"e`sw/Gv=4	@%CtIuydFP\nEx(6T@Om[V \@[g7ICV#o?ko?biGT33nnjO`VHF"wX|[K)P]
OMxUblTt)?/Xn>2YS")<mH;Gby
NnyX;>1({grr BKz+,od+e6Beiq974`RyMQ<#l@(1TKe;"V~
0-.c;m^,.0;L&P	i "uNeu8;6H%iuIaNXwZB
{q
/
^Lmf%b%wPf4Tlzp0[kQ_FUHlQ/Pf2j")qt9k/'()gaB4|efl^0M#x=8/rohRAHbY<WG)^3VJw&pQ<\\u$;<t#t{ZxAW^X)[)&h7m CO8$H12})7=7~7Z?{5j{D%0-.#_D)5X>[_?`!9]}Z ,gX2ubM<PJMJ7wjsnr$+xd)xM.EMlXd%h`}V9h0}(/fi6(y)o\3.d9gU{^'q{x&-f."DVPAPiO1*f.xBRJBTF8wjV<(0X}RllYwTT_d5z/W<H
sL0*D6F;#o[F1BZKukoy3.SNh(EBMsq7u/Cy#V3@#?W~8O9).(h#oZT;uTtzaE4n-SN
(]rBc7QgE1T9 .U:v::i'VN71jd]/64&JR>>s
Y!m+kh	fb;o",pzrI!Bbb h&g25v|br1=i1.qU6E;CQqH31*
JQhO ssV_[ge&P1_2GY{$o>4w#UIkkx>Im|D*%rCftv=3/_v:r`*8,\?E$bQS0?O/*co8IaVIoR4>j!@w9SUSReY2_,\6-eS,nn\w,RprX']I"GcrcGMB=DyyK7c`8SdDn6/T^vO|^Z$B!/|j	dtb?
)B.Kt'H:utPBo ]O[,U* K7^&&>Ta(PlA^RG'2+m9b|3,SX[+;nqJ}pD`WFRp&UR$rZsF/yO4r5w].o?I6)$m+#u0~TnUFeDj#WAQA);|@3S)ja4"L7)?gM2119eh'Kmxv;T	W"KD)^,p1DW&0OT#c[<Ro0:lH/-gM|v'W y2XuG@(<k
[4V`Jdu&rTuDO^W?E!]/s5@mB!<WW:+Fs\j1G;-1GW-;$]Qr2Y9EYOq4GV=+us[E@7qs*@{Y=<5V:'	GG*:'g'KY;1\6}CS<|?WKH:;2QMqZv|JWQ)L`BRLfRv}hv8[_>OgInWLc1B&dR@jreS*it[UZ5k=Y|"rf2B@	Um$
1Z9ZPZ;8!o.
9=	[\Zy[V)9QC,e;Vk&&,>p@f,:>z
:+v7(|#NiaG	aL5GIW,,a2d_E|9vuB$GLS
2C>iDv%P*8Yepy$<=3]5}pk\s+D^Y:|73
n=,a\SAJ\mv:ph+NK#?^K2'o4Cn6o.U2gv7Ft4ePaB{<ahl!~y`NFcAPP"o^eCdt`GcX,g9wZj:n=
R[!;VCd/I+*op)'b:Qxpo7{"<`>WL2!w!JP[_Y:,S7"{EX'S6M&}=R0fJW_;P^4a@m96D!?12By`e(-haD=7yB#mc	qY{In:-0;qoAZ G=Si#X`Dsw\HzP!QE@xPEw)qr-@X6l{^7z~26L{r!Gn=]78D_Ub)|+-xY7<$$ttA.Qp$xBs%)[v*xak*H>S:*9:EEK\|UK2m'^+6n.v%kZ"w9p)^x+I2*fI+e^-#hH#I.I.Mb|HFL;E9j=N#=/X)-{	ls~j$(T<.A\faUq%S+V18cQs|s+}9WpakTvrJ'yr*GLw`q]_h5AwVB?hAxC#vQJ9(mtkSACm\r\aV`%D%CM.&d|EVE&c7b{[D!vm=.g ^z\;.qtcz6Ck\$j6{:z9?RFW:+?`@94X#/`{)uuoxZ9uFW{V+:K3Im2sR.sh49+.dv4l!0t?oTHG/	h8fJy&pL"wL7jA
&iQkUuJ3c=ERYT.b`H)8hP_QX
-@
i*%h=d2Nb1Zkwa1KR]1@q9k	p,4Wwt$9$cF/_a%{Dz2LP=w^POl/<^w3+%kp;Zs AmfXzw
W-l[%,8ZO.;c	wB[3ddiaD`XELUlIKRc?wag>8,:i%A|<8XadU!,$2.*o:OT|=b35vT^83[np5kUiW.s?rE|\/)
%XY#oMsV78k@_N]7RWI{H7t|CtV^{uItK,u}n`?npk&/EC|0aI`Ox0~\`t	jccCd(pL$@y_Q{Q5A'/(# [q1hAeR]qRLdb7z!hiX5<9
trG^+^roH"4dcH7d*;\4QXIfl
KkHf)YHgHlp9O5Fx6w|3D
x>:N$%k9Zl&	mf4)>ZxU8PCM/eNh{"HerkQ*o%$~mU2#3s9zXDmMMR:wtq-|]$N^sD.Qfu8\'4kT*E}1ok`IvCg&)T.OE-RXq\AXh9&~.L D&J4s1}^)(K$-&@eXmQ(+eK"rBYd<H0id3l,b_d4:+Dn wdrfiOM%VnAE+OwC?E.b`)I.g?Oiwcf(cw`A.%9&Q1,l6Z-RcyoDP"LKTNWPzO}0xcRN%/vm>41!|I3<'g69?7rCZj(-#M+LTkN77adMAH+ek`LBfC&ZYge!$a/WM-2:P$"g&9@j5rQS.zMNL%~)10bj;D={c,PXR"6t8
K9h40L5npMm*&xR
ZzC68}vF>49t"IF<^BLe@u)x!q~\#T[C_'RL|]-))(@1]V^Z4KqhYfm\Peu/@"!.nh*zCTpFiBO;r;"KyOLKq<oD}1TjzJ,_Pm9^(4!G@mnuWHRRRgYb;oy>$SK>=i7\`tTm[\pn+^%C5L DF]V.<"sC 2iY!.

42E}TG2<anCkD+(IBil}ek=d*v.#*9{r)NJ9?DT:3mgFqI'Ll-LL|(%:*OzD/NJ3(Ekd~?!C3s\rv0%KCn?!'jHguwT+vOW|3,**W#]hP8+dS?D/? ?o9{866i%ytQpqqyPQIa-cU#]eZ)o"JydY?u.{-PZ0}^kX![|@mi sc9hZrD[/X8X87y\`?9(G/hW
p`;LeJKD;!gIJ+uWmhwBY#|Dk,7wpY-UAn,EYHS>Yg.i+Mk$R%7\E`p.;u_w;+3p"aIYj]6e%7E#/S(L aA;rt;`S%U`.WX_|;9IebkSkq$]SVFMGNY1H^2+iV\PTcyI*/G&8CFpfkF`grid/mGn@mKa,U~P371gJnxDt #Kao$=>	6(q"~Rx!>Qvd1t_!SWr)Xg]2$l#XbI>s	L#1J^tu6JB\R.g&eW{\&1SagMJ2 t./YM9MiLF^;Dz,iLfdhihl3l["22*M2M`xk<H@WYX>)7"FlJV)/N9HOmd9`R'N|G}$=O@(AP:-8ph*wRqsYw>6)^'|_v[U7i }QoJ2 ^Ap?y"+9~M5)`j_;fKY	A<GA<ZOFx}\rBze@@?pTMYfw}[MRf9\gD._2L{@?E{'[t]p$i1 9
l5vG+v`O^=6yxbsHW|.THA
2!KpvOWmu0i;{42|YZI5p:ip\n$a;R=G:4Ati[6v$v"o<P<]&tPsxNYHk]@ZNiO}:\NkSe;HWP3K</daxvaz?[h0,MjE':lYT=M8uDh-z#0&4~h0**}qAoikP'8L"1J+D6gGb|!>g^lVxJUnj6.e}2._oUHSVu<|QQ(b[:%ZPS5^~@P8ro4Z)Cz(P]QAM!,J,_S5q2P5?$?c0Ej\w|s5~-({zB7JX#Whr`HcW5w"]h:)wkgZN 6epM09h;0
*8T^Yh?"0XCSBjb]Sc;8"|^VUY b0E{6N!8tmO7PJ0(xZFU}kQRlU$()k:l}C8-`<{v]$e}Y<=v?%{$>q8t~wA'NJf?v} D&=cu|p11r)x&4oz$}dnbhK+"l6krMD:Afa?p99Gp/'k~fL{szw%1?:%q8BTyP8?I:o5&no>bl|7XGi{NY	IHM;t1^n.P4-\@h_!+JiLJ5"#o02K]IKo/zl8~ Y3s-[E?INOiV	._9|6$b|$[f jm{OCBSq@}']H?Z?,E74j!F(&HFtZcO>Ell9_2|!lXp2DCGCi/LbwwE[0jC>(GiZV@LN^.#o55GD+ihgr'i#IC	RJ;f<74H	FjO$])S32v4+Z/uxHj-T0\ft .xtyIukt$O=$RiM/57-tl0,zu`PLG'y\)e\)BO>y|%'^N	|34te{
t?azm&-<Q/._pc5a%\,O9$?|S P )P;~)S4*ZdRWx\nA[zh!xYrXKJA7.,b]h{hy8`*QA=?FbfwlACj1WDQb:*2l*f,6q	;@M%DZrpjy=e_cn9`mI#Idf;1aC(piF|ux=^`Jm9:Z$q6:?5J>lv%6KaV"`c>==n]VV4.Xz#XeJs-f
Gk<ft[9Vn|4P,g+63'wV`Zi#-x!$AhoYi/4E[WB%p}TVKr9=E	
G"T<<mz7-K:tuFbcLxa?DIL}p]pEKy'?="5;P,'5b`VCy7=%fj*4aA/x8vOWB^rhDD,21%zpPON!GOM\u!eBNyl{4z(b.M?3X-TA>C'LI3a>Sjv4<l~	x]e6U2*wf<$fPVUaMj~*+5"oQi/b*O3g3ad9<sa*>RQ<IC !m!cA>;NxKMfnev1<~ot>4Q"0xpVXIzP#c]rv_gC#$vzf-ckS=c6Y'5=z?y]=;:$!',(3jAOQtA,g|X^&Ojqtb{O+W{KU4JJ%g'M]GOFB6QlL_x9'kM|m}%^qqdjIBp$3{[,I[E2kZC/<|86ODips4VVAsR 6hp3)x:<'X!Y%ze$wAKgSXZ6w ;_L}MqeJv?j9q:) <DIjDuf ~^n4>U
9ek.#uIkfa0N+4W-y8F5d@Ek P>Yge-WspYPo|M B)%Zl%JMgJpwil6*6CxhGu1j>)WvRv)86qpdyx6x#9r_\A:HM&55xhXJb+WL#iY^"X5NDqpT4+((?>XU;t@N9ySyB K<uL1Oji5>hd&./%o:\!}(~WY`&0cQ)
*I[y]Xb*ctKq,p5 f56'@U$Kla!uu$Qi35!dtAa9.)!gh#Q66LkW<UGMpC&(7ePwD*OSN5^\sZL/WRZ3~ea{VW-5p
Y_IL52p7Y42 q_zDq)<O(b1(U:3##{k@A7~LSW)=O$&jM?~Y>?-_9..3b\njlrw#_[dpdAONZ!}&#!qP&4}uIlGtRX3bD%ox7}%j0lHJS?zW_AF%n7.UShEI!se#Qp#Q8~X$778Kkz9Cm8TBs1]ysp!xw]@dwWR]$mbrvMGAzI-4+G/1upy$:Z(*8'@=YdNX\0HxF_	9_b|]cL/V! e3;
>quFcFU`^[{j'(07/5ux^@
^EX:LNtJ\G7('pr"IFH!il)FT
7fp&Q_!* #dh]?j(3F'|E>MjSCJX~I\tfI8FdM[/X#BZ6LqR#$FwvY0gz.Wj=@F)jRU(_shePGJ<@pF0XACxoeGrvv)Lx[\7iS3o`xR\>#Q	=[RC7*#0PJYghkfoB}fdwT>2A?@',6^U$Mjpx\(@W<\VV%#:AvJHVsOOkA-5<w|AQ%6<WB7S1LZZ@;hE>
DeO_w5(N_K,:%kwqLFk&Tpb`ny~cP(TrLT#C79E_C'qH%?ad-*F+bm7f&{9o^M,+%?#J8!a.F/UffN,L,KFDN`.Q''_!DHa	p$<eT15^H^U`sl%?I?x%`QEjQ0r+H+4|:aK!7>S<6A9*CtMi0|{	YBvOk|a!2gTGb%aba%!	1ZR+,)>'yHdl9aY-~h:4fy7b_e(F	U48D)|yiYbP8aJ71<2xsFW(`~}!wtD	\I:
xTW?/Ltao\c[z+$xMa4>S+qP@>m3#u@[A7c/F!Y\]K'a;O5-
y][Al&e:/9bvo2UJyIAVc.6=gm^Pk^5eZc)9rXn9bH}/@G?B^3kZrXVT`.2]2CP{Vx|7:xg6QJd06==`LB&%o-:=YkOh,D/H#U7Y9aps$^g%kEjJY2f7M
1<0U``kl-L8p@]ZfuTl0a-"a-YZ4 !,\n/6DSRX 5K}V{ol-v[".`>)x4e2=?H@mXfOmWWi[?E:WxkX{ iP;xoU(%,
Pw>HDXer(a%%L8ltoR6V]sV;}$Ls73!Fh9q\pR*AXh{~:JcZGgk_naBGivwn%fi838R1p!Q83-ri;JguK](*gGg.2~;u:N#=VI!4hE+z:EJU0?$M2Hf!J]QD?>yZ*0AsX=)*iqNGk2#5xolW@D-kz?\M t5^:#m[5w^:o/c(s fjCq4CIk7{QRjlL:`tRbtSI>^EN~z0|Y%7H73$*$dAQ'ux.^W&emA\Ef\^drMOF\S50[\CE&Zs%o9OU*T"Mp"3SPFOS{_$2ffFVNH_>	|/\C+MI=N<#
-*Y?BvK19X^;6:JhSn^	EdB]v)ET)hz"((PvpQkD!8Mnb3</tS$+GIT[!]vDU7m j{z3sG@^Yp!Ad%Vw,^rba8NcbHoz8LZ:q<p/3@EC_1 TLGp0|=A4cw
7,+$|_gOx|~C<+~$@,xV.OkIHk.e$tN;*Zj'E3z&^lo!mPLny&K@r.j\uv`]3n;$wht/Wi:o@hK_`s
qL=KsWb|*
"ee7OR1xcgk<N5EI AZrU>BS}?{rrVpI*9c;>=.KvX^SnV)|`XW8:*j@]=7vXR"=0GJmx,i7c1=~"dkV+W;Xag[KXBKAg&"nVN\gq`'
H1n%};}`JfSc%s!	>?(?Df	q
/3
IX68"aLZ{arv< =`>IW6crc_$-/2Vo)?u/H5<U=JpwKC3=>q.1)I@>&\t?pUFBE&c.wFOdu\*X05s/Zhl Y,f!!Q&LwOJze>$.Z&j	q,sRD8'CZegs[h xbi/;c6uNIa&xn*;a`$#OB-)EN;zYJS_i	<ieh$0gL.7j6uZ8)(fD]L+MB+_e*`_;-L\"kT}<YC`J-.0fLUAdX13T)Ny*p|l\5=AqB_fgyU]HROcPJZ]3#+S6.SOgxLE2bTF"]\l}*d:d
<Gpy|g"kSfm#|P'*$)_WGVTG_tHUo DvTO3wCO?}rk&
tq}fU\`fo"e8,'N(Wf@O)'bBeoydBN^e8xXBvjb|]fsX>Wk*>w_` b\1Q@z]Y&uP!TX^iWP<V27#rb	s>6K*+Jz$wws%|P!*o	g/xj_#<SbqDX"S%9VS1!5H'&X:8~dI^1ecoa^8go,rWQ38$I5m7FQ1d6~K[WEFOII%<|*c5R:}#2Lym1?x8.'x	bRO8yeMt)*|\A~Pn<878"`z0<<'xJxde,E'z=YH*dA\?5@.iyaH)'k5O_X\G@er3}Le+fG;|z\W!+Uj B@ltBiD>2F#yo(
<jr.XN]r(~Ei1\>e$&VDWZa9RI^fq
=TZ]
XiCt!kB:\GZ[.j<}"<Wp5b')iOU;q;$J)7woxg1<n"h0<MbAG,YU*u4F(V1ClI><j5I[Q Y UgRd~EHtX&7w<^+L$b"CRMasq!-2iQ&4sKEGE#K_="j	vRF,Z)ljJk?gBNE],N~:+%=zP~F|<+Wxl0$jaOS=J4MQ@toC'gS9)Q03EF3|[6FB(WaD
iB&#_n^`{#/ZYq<<ITRm
[@NSFhM)j8%kVZu+<tG_}sd(hnzBr]CXMOo4J_=;!NS1"E-Y0	D0ro)Rq1N$$
*'QZW<$U!@*l+wUt$Ih49hnO@GcsQBdoyZL8^	Gld%drrQxsHP'zyJpF2Ih|PWOx=^[FxqtC95 i5+E5vQ/b"8h7EaX[ZG?d $L7.#]MYvnZs~t4JN-!PSU3u$"C6!&*|ZyNS<=oKHbb$0i_axCF%JvNfsur,n,Dv}|)$Sh[X(&;fg`G, yxh]?+vp*wS_oW9fI._hbppWU9[y>Rc	|X=9Zv$re?]K$2 <vS-,p8J-^]K'^1[ C>8ML1\9KPs{09k\C/79BCNu#&jn\55VI_vB\axK9?eIMA-V^~vhG"2C	[/CHQ{fY_rK2|,b
f#+4e>Q`D/yr!>T<.%mLW1iP:[rkM-K	2m0\;9"Z`XSi^Pj7(]uq71={s5jR@	;4.IL5/Pt(Zy>qU0/.]Zj]I@he_nY e3&\kf1F@@q'_T<vUXTUq}D/4syrGDK]JfJ*`c%Lk<-exc8/.7M!6P@	1OV7jx$p8*>Lf3`cA:/6Gc!m[[ZR4`2|E'SU2aqqi_e-&+jMLAi3(!r/l=PB->5:OIE{,cW|aU<Tqn?]u<P^)!b"AhTIkZ+u>;Mx^FxO/>\TuQ1p?aH.l8r(@RiJbgGaZiWfw~5d_;QBt;*g/v8|'I1|;R`NP&NBCe.ofA32Zf0pq
`5'7]AZOs6wROeUJMR9oHQ_2rd.8dku^9(Z6w4pwY2n:q3L&jR|!cuE"M~a5TyLp)ZulP369~_mp+0ay,1Bh\GnX+!Tr>qr[<5!AM!tdxQO]|gAiLOYb{mO{JAjM,.x_R'LP8.I@u"cF(,LCR%62un%[Al'G lEiiL$]K2VvZ-@y=d,F(8fZUQfr>pRscn|q3Z`aym~kGdeYT#~Vkh'3A(Tj? *u]_D36Sri}"IzW-(X=N+uo,Y;wh7Xm/)@bUI\>nz&_D^T)x+xB''VgkSj!-H
0#0
+6KO@ewi>}S~\-WJWy9w+PA^&C=%z9kaAr\p!"bt*d{wjRxiOj.B'EHHU`kn Dag7_W/g\XAlJk"&^8A|61wM315_6p9MPyuWBG
q[g'}*SXLNA]AUzQDshE
]v8T.DBg;,ViKS,QC-&fnxJV"HVqhf59f|MiJO~@5[]]B-Mk 5qnNx<6.UW4M<YDs$&O%DgXUO.^CvOk?<af(Nm`&63eUy]iyUE1",hnbf3pi}?6jOEytSM2QCsH"KbM*QcWrH3+MVySfvL}QAhQ>1Bs-3?[-Q`F$6,*Q:s/==Kb-qyT'@y]F.2KN)6Z3F#TT1P=B ;/P3fq,/6;Hx9aj	+2vgN,qwaBpzr3QI_cflPI}s2f=@<q3^Q=D\Ih~U)h-TErlEM<R's86-KF6"4pSqk+pP- dj&[tD)O_=y9L?\+B/JQ.Lb:KmO9f'&l.dS/n<zWz\T.?%JKB_8.1$68k7
]O+M?&Nsgw6M,BSp-=1;q;M5<]f  JGsPm\c~Bmb\ofz2f*g	/c7.4wK:#?uj:c8I(bj
8fQaRabVp1,p}2#|sWt[&$	[=q4D?#r4l77-?sj9DQU0#MUTFivgc`XS4}W=]z3*&:W	_x[{Caqa'}:GQEX8,6qm@HFMN5q(jpqB!$rqw3O_';Ri@ Y!*{l/+(]o@nI]EKdR]^I=-G<T3UEI3AYu#;L#u1ygi~<J!S
j_{8zMCOE70yY?t1'*Ap@&uoLgZr 8D&oCY#p6"<;fwx{y7`SsIa_ED@1-f|+=i|x`m9b sJ%lhUvwab~e*}fi;n"):+U.Pnq	EU_3EB8%0b##8N*@4Gr*bcp6Nh_cRs3)f,[6n8UGpa;XcP,faq"xHx`PaWR9@C_zORa^AHS
W$Y@L1pdgMXG-%0rCP"5#*5lRM}8<$NTVmwKSAvrR5D;0mv3C"H]DL8pO7`wof[vjm.-vO<AcAjXEKgo`raiw|)0Ga$1TY0t"m}P^	uoTp/g/SPM-KLbM7:w$cCstI/o>rm:bz/t?{
~6|fm
h"i~
qA_**>Ua:/N47:yJUK7+J4H.H^>#ai
5$5#I9O?^,STDb^5jHYo}Q`D
_RU =*7
*gkK
=X9ZaD/olE1>/))*5	[dmit2~{63)><o3H^O5gi7<+i|*0"5IGQa %^@7+[l\V_3e?!o-weR7<?D<J}OC<\~(#Y\Fr!k ^'}Mq$\LSp<thL.NSadGlJj1}fjZ0^j_W>QrfCoq0*EIGV_"^!|H1o6#;y@zv]'\BzH&u	jq~\(fpsy785$N
7wU,.~1!yy611CTaMY\T_ViEg!QhvX(_L%7-u1~hkMM['|d{.Q<	ohEPHivB`55w!G4Wk_m);<}wa4R>U*{c(~|ViZJhfK3D$
q`bM^sj%KsS3lTq	>0MKT
j/Wm "ec-TEsK6xwsPqzR'\^FJpJA!X']HFS0aZ@a`l#q'DsNG3.Y!Jg:6;3;LC;Q}&:^+tFQ'\3JUF'mQl}Go5uc|
I<dUWJ2/]0[4,e0U^TwE6x}IH
eA6/>D=xU)uDSP(T!bhGdWj{n[=}rWyY=|/yj:>D9(2_g}5)K(,kq{Fj
QB=m6
I,\\NqWc
ocv{=
@$+gY4JDype	f!^8-5>Wu3PfnjsAp7bE=Ra3MvKx>(P>pH(]1v\PpP0iOAH{{ic0RzFp	W_'x
AQglET(~9rB+io]Lha7\zWdWL'My2]gGG^6x1enE% @;{$(H,j[t>D/ROn	@7mAPztE8^QZ8;J%pecdLt'/J?v [ HZJjF1@	GL5LE@+jTH7gprS;_3C4QXez=`xpC- +7^UP&10#KomWBF8au_i,?RFDpnmK$VCT/?b|6Wqgy10gg>0sYuF-y58*_A22ZPSsI3|i;QKLHZ/7K_gP#Qn|y*.6){.n7FdE}.4yu|1PE)jw%.8&-MVTV!6}_SCmv$+AoO@Q3Ms^CHSE8}Yf|!bhP{M%>zZe<cHbXT$b"#, Oqbk@g6yIl29Sor0	\|K8`W" $iBYOaum#*H*GEp!1JvC;jJ@_4RM<)}9G_OsE$7S1,\tbt2O@*6=A$AD<lh"OpWqBMtt
1k}|aa}oPZb6J<p8LrG[;Yu+$c;/AB3U"UX>CCknx}|c[J1}x2lfK^FF%Cy.G_84rh(DS\K5MGy(PI_e&?Uaf*:W\jL"%GR%l'I3cZe(tzf1b0,c:aMI{@Z;cX/q$iAN!'Z3K)M8)3omhs6WQ2mq2KIpROCa<ThQ_NUp#/ WvC6(GOeXh4iP=	82GC
dI<TJ[FTc}?ij)7%~uJ
G:3Tgwq,W/TIvR1hIF|}hHt`E9fBihC~ZQ%qi`$V^gYT5QI?@2+ePN';)]8#<W&bZxwDK;eiruwe'F'=[:mWB_1L_56R`tQx#2GZxPY*<T"
Wc3NVOpYlgt=}yg!hACbLDeaJa:	7Ft/|\uXisrly><rt>QB=cGU(#0(oxCH/GH@@eK[fm[oW7G6\2ar!]Fw;!Nv-ySDIkLQpk!?7LF^	x\G^pOW:M)rdc6[@>p~ $sq`\n/pW;h4>}YC>8mL\CV1Rbub6tj2$<2*JoxpvFwG?S`B\p:*N1GZ
0IIRxCV4(9:9k?rTWxunbD?PX,56MIT[XK3uht2($)jJ.n'sp	F-TvldopTrLqn'L|eUAuBL`9P
(\J#{9RG?C"XqnDL\Z6Kj5YPZA#eo
V5{i.dZg0B&=CQ,yF^9G[tL^%Rya ?<+-K{A6:I}%QeR:b	'B6cM^LbO9i7^]y1$QNy"CxT}pSd:|L3k{<E7>X~w1l`tKZ50C2	z?h!4Q1J/"BMOXO~.1 OE1T-fuz*(43f yuji#ADg#Vu&v>%;f!Gxqc:#=_'B)ETqmBG5[jNidA::81X_ksnPLl#td.'on^yCI~$ {4q%@qf~: r@5o
`y[C1<xJ0N0nh
lz65S0(t("eH]qg}sv7A?89V`2krd^5;`3k6'{]I*p|QQW{Ik*@te0GqcVC+equHvd+JY1xKJeq7T|^&Uhm&'d#PWs!0+F}Eut?fmJdg]9R#WjT)IEX4z[$sZwzI0YF\IdO([<^?'Gwu`,	U&uC]:A!2kcs9vi<]RNK)A"B?~?#~Vl`J3Gqr(Z;l<^v.yz0Csab@,GaL3Lz"i%YF+Ryxb~`:,*ocKv9*|I[/E:0j'c]b2hjQqhBl_f!54X(iUSOhR}wuV0J)jNne?eMF&}MC3&qgv{Zj7e[({#^'bfjq)__?VbCXe:u.D[jXc7p9/&`Wnnx]<-=)6u[GwrYUETifpUF[crVZ>;n_P_Th]m]\DWEnLA	GM^t;8e_<9"giqzO
x%;o+aA/n/pN8 v*E<C`J"V$q&R]q[-3)k-YWW rhd)v*(Og=g*i``5$!}/pEfmiU3W?
	>4^N2 ]9M}Ds;Gusn-th+$0+97$/g3e.HN~%cK6"MVQx#f4&lF#DT
m?Aa0[NN4XXzTeKZ7Mg"VK[]n_lbSvj0HqqDN?Xnm%,"[
>]U*@n39`
o\$&PmWV%j3i6I5q+[/C9.Y 
*Ce&zzyqn-+BN4f3 3muy&O\[oc4
^deH(>5bc|E>Y?T0 GR=,bSAK1'E7\0i`KDPSn0+\d#NY0|DZG]HEJ?]WV$
f`DksHMP4nAH'HJ@4ZvD^ta<X*bA)`NDF3B5S>Hb'
A	j9)'@3*.T2I_v~"{kL-/S;/Frny-)AH*-uQ)7Oh`A2W'$}VF#y g<TQN=18RWC/F?*)8IE6@w1LK)..;k^`|)L,/@TfEBr$:FMi{Av		*eO9s|qZ\fW<lz"hp=4b,|GPfgplA#	|I4OP!/1,'m*u+F'`oJ|`J.bNdm*"(FjeKTM*{(	ST[i-j$HbeS:6y~/uWOp)Q,(dl6P%enzfY X1AplU$:]&lW+jW8df7mj"Zm)#@nFqWxbmNTB~an3I<xjaHsHV4sN50KoL9"k:; @;Fe :=IXR~Ud]KZOg`s1c:qO4gynYU[@
2JfPOa0%{s\XXB"7d0}w)4P2|^yg"jwXO%<=L>*4
v	jhwsRx`wN	>i:)SR8#2)z:`|mn[&Y(pG-J%39TTNy pdu1z_;gG#Cw/>h05/mO|iD^ZDX{5%=sq8V6`5#/p]()ypB67mco#%}e7?WK*(?]ioqdg7iFl\"iCn6IUl.DJDH YU1>
:|*C?<X_cdN{WkvuK?]&YpmO /8y#.GQi/IRcfDYCnewi5U|].37cCQK%<ySJJBvHY,tmFthj[ 'C<Aw(Rd1hb7Q	E`5@9/vJ-xbo+H43guF})&vJ%1)^stPXg>Uk[
Vhx;[KrdVrFCSVM)RL8XmLTNJh{sHoRV/D -t;\+?(~07>6nM90>LEOSdD P@Y0
_ /-[NF?u2d!i></}$9@p@?6Q]37lU}:ss(FI%m`bsEuXQb05w'S(+y(#lt:4E20POs=BsXN4SB 7N=V+ri/WZH=054(SQ.*]b1!+
IV>E1G%s7?ZY)jiQT?MI!2I9n5s2ib7]|"B6<Ief^g}NM{tPBB{T6(2sXjQJu'(*JA>b8/Gwzipx_NkV0&2},,F36m5
H{&%! NjE,	/}&=I|n:=i/ZNMmIR,aUm$3X-IM,zK6bUR9^'8]KcH1#; z$8RS)wvSwT)})O@VgB:=+5Ec2?0|fy2nzg)W	*?}+B-p>>vAh6PehKwPX7'y`hC1H`HMwHRkJ!C@k6~8p0:oVSba\(-3Xi(::I3%FxZIbo]}mRw<.NgwyIJf39FCR7@*?:@EoL)n
@<APACm*)<Z.ah9%j@"`V[_,6%U1lq?ts%PrQkRM/0c^l@fu`>Oq>I]Q'u3.8C1CVz;.F!#h>Own[]4pW"NiV}g/P.1arcfi>UT(18Q3	U9\#>Bk=?x3ls):y!rQjV%	x.5@VHAt@jKTt	}	>qab.$dEgy-CA:FTY~"/,2ncNQe+DZ|>DvD08?Gq{>*L)B%S:VPxAK/a(wrc<V:&s!>1])	Y)$[<lC5	Z2)SNnNuj4^h+nM0uIA)Kp	&.`aiQuj0AKm4(|zJ;4r#E}jQ?L#,V_/(	Sz^AjhXi9G=@0E,
}J,&E.#dpk8FRs'%:yb6WlX3*N6AFA "YgK#d@7@VRNG< <13tA;FKC%"tRM$@Q7TtHO@\l1VjXasU(j*lNXxE*\>$lo,'}4;72ljk~DfE1=N&lY
MSGM\oW2?*aI?@=]fouxdeCJV"BXmK^10a&bx=hH,Tk?9EA/8Z(0V dmmZ6uzt0[F+_S':TV_U48It-i?
?O8yH`DC~2'pW"UPwB{>qA$M>p82L9k=:`g7s4[6#=nw	|=`r=":LN~%}T7yd?d+8d,ju@e5,]:l+(p+f"Li~D;bs0x&I/Ik( |*Z"}y{>E\rP6f5DVpZj\,AM
aZM!cbcADA<\C1l;5OWtI6PBx'AP`O|Dm s
jHfN-geMce)LUgi{BV3o*|G.gs+dz9RL	+7,?Ti?GIn1irX>
%R$'0Yld"y`<&; >'j5WY07M~JdX&Q#GfN!
>%3 JIf<u84HyAu7v3;lpz'Y+ip\"AC`6
7_nz1\A{'CPtL
H|R?)p@,:k9_/8>g+sWUx4n^Oy_quk4ueX7^,(l^lO-(2{I^=0?&5t4Xc@hzsDX$<65q|<gf`HC"8iR96>6EQw:-fLQnG2U5$gWG*<weMa;1/}Rwq9J=;MKp	'AZQP6A|&cZ:Rf)pJpG0d|:e`=^FKQ<"b%lALXla81b]
l`
RlO8D6E"cTZ!WKi$j<Za=.z1@x<jW378"f%JEMJfYl_/HD=)M	p7HQJKUX;rpY}g^5$B?SH=|-7g^4C"K&<pj!it\_q{=qI>!M#d	-0[dM5g&6C*Y$#6+s4CVr4@DyVK1Qrs@!^oM]CUUIu0.V1.,IOaUp2P8Oc-vbXR!!	p`*;DD}%%kvsa!p6Q3o.SHh55*1h%!FTa9z[2p)Nfx!TTp^3Q,(8%oF"rq3sGfkffn3cm` <3VJYT-H^DKV|:"rj%+3RqKYb	Wq	FP-YAZT`J+DShBEi?eUJokY],.cR5aX|^iVM+tlE2rZTXC}/9)}+O4EIrT@k3g)"zX8`HzNb&zY/xK1)N/FV|21%l'n/l[Q.oC4// 0o}$^'!Xvsaa0UA@K?Y.UC2(_nzo^j5\drC\=lGRi`vXP3ftH31m2Hya]iS*heYE"$<eir{j%R<iZh-9vLaj]!NsVJ/Iz*_1YI$zQ
k$Z[*30U{4%p"p$>G`!`VuWg 
F8Amu\4fY$Q#d%&-&L9>/X+gz@ H<yD0qov7R"iZ)pnZ]oB#SX65#Nmr3amo`4X58e9"z )lO	c$aVnr2H^K	GTR#{=ztPJ?+4&:~Pv
B|,AOA(zif76y4,`vZ=)\9%J3&~,MK:E=	_<0@sll
0v*YnPJ
5t4<#.;(HBCy\&;W3sG+qm[[Q;:r"|M]s~e0{VU<pxj+}h(67>BP(+Bjk:j[Tg<<o(tC8L&'KU!x?a4[CZ@gtf>S7s(en0^Gx3~xJN0gw}ht %2vCd)Pw8{jx<{_u7mS)\+9<dS2;jH}I|BMYU/8Lj\vc }Stfu2zX.(1T>ZKTqKA!	JR-D[IB@YP&e{WT_?-PAiE}idc%0ZK4,[7#|y@zV4mWc`\k-lB<|'/4i_9>mGvK)88X-8yoq!J4X}A@9B
!e2q:00&cL|O1@KDt=lF&lD kQu:}A?^|Yw()0o1|NIOL	lY5a&pj_`YCP">"KV6"nB>}3]n{o )9Q$%w*vct%m6~oq<k	1&U,teylJ\LTw+)r,w$!S#(sia0|""9E%dSd@mCk$~Y,9R~-/	s+wPR$*"6n4CX4}.Q%QD:_.oE&iloEf ):LTjdW(W-!]A*ds&~
/99L'hg\0^<"|C
y$vHq&fIvz=Kf\$<IZ.|pt|DUS\+6e[(]Ib^bkBmZ14VaInBDnyIR9a+S73Y=w^qIZYBeWV\roMb>A%7f^N	.|zpT,>@7>%7v\A)HKXy3X+%L(3OG"i(1E0c"v%1eODPaa0"V.}*"SUAkN5PT/<\]{F/{ufZjIME:\H<_J\`o!I
Ag+7%rb^`Z{Ats%d =J^.j+bdOj'Y;+	+?ETNS{(cd7L4uF"tubA/>+
s)mvd^@Q)]|0'V7yl2sXT<&e+iw#4xM,J%BB-h{EB>?Y2X>hiugfMMOx	(5X>w{>_lby,ex|"52AgSJ[cp]D*Ub0]Q5C?3e'w(L*ho-WQ6[f?j,94,)@;R$@or=07<?RK2gPXS_|2k,C/lh]v=zj|UP8@|zgVLc@vbg+OQT<P0onYnffSB
t?!O/n0:c)L`Un[w-n90K:x<1S4hJLW3P,IUwr+7GDz+~Lth0b0Fa#YcoBz9otw;bYMl[K[A/-O,_?4h`XPZ(/Z+
@T^T	N"HWvm){Kjb;MgN`s?TsI	#>4t8QzE)ZI;K:~%wL^d>,CIQ&or=Xn-Kh@wTG&*#NUQwS9:Y@5Q	{CMbF	)E=eD7G5jt
4+,j`RielH"T	Tf3&9BUU8ogl#)1)VY8<.^j3Jn/>`OS<;>yZ6]xBfz-B3*n##;J&rmbk.KXXMGPv2R-Sfe32C(iWpzSL*_DK}?Pbl($hiCo]g^g^LSY!8JVYcgp]B',>k}_.";oP]c^C&Rq=}<LS{SD?s;hZw@ 4Ws\B?'vYpbpjDA(gA [`<DLcA,_u7{6ud<a<&T<DID%<aL\kM0cQW/GCZ!Oq>Y2QU*e=9ev.Q2,+zq9f``HCGv/vE@pMG]F-*4a8B6@=,\RYNpxGdh&ZX717V2(DOx~J]U7nMhDvy	'.mrdIs@*6J4 QasB~	hG5~[>)H3*kOxc^!92XU%kWQBdRiH8=Nx5qc,KNV;n>+HXy7C#sh":m\aKw`bA}6ChVA${xyTPq2Ar>G^jD{m$,p|[jUcv4y}qv6rp5Qm?Rlo0:)!!YE>=CEj{Dtor>j{l~uG!=Tn]:-q
]jq<Q_Zk(nWj9lR;]E?wz"(E@NP-&_!AhK6~<>
{ !>/W"8mss#	Hegf9Z34+Z3.dajs"49utiF>&KdS\Rn_QYW!(}DO!:<u(gz2.9B*GYG;yiLL2)_va^r^L+q"NhlSC9s[KieZC+qm	\/t|8JG-# r$-V_^shLZq}Qk;9E/q+vdD2u//)m0kxq:M:2RQ:_x>6xe:qcxB"u$BBw-"kB)k]zC`0TghebE*oK~DC`7CS[?x1~4{bKz.(dS{%CCLm~""4d0T75VGM&xDR>iNQ%/)t,3dk9Meh%|cOBzHd2M=TsM59<!`/NVF^QbuT^!SN`v^J+oYt87W~0T-BO:9H%D=GM%@:EkrMRM52>YftzQ.@M;aoy5sBVoj43$=psghzx{d]&1sQsa4Y/~%yC9Bk%40j0@g[>^7=FCBG79Xs4z-I_+x:9?@(9})r=6wvS`XtE[{!g_VK.g(:&(]N4Qd,	Y\^TYEyV"%Va$N<>_MC(99,99!U?g</na	>@|t^fh_s("}fT_Dtf|E>"2a!*	v00-n%|mgv*iS:| t7xZ9\sza'}V\uh<bc,,AvpJa*2W;G,&5VBQl7k	n[lxD(@`_)%pS@$H:_s;%D*5'DW-lGk1\@;^R5_`zCE\LQa:j{T}L[;6&^0"gnv?i{ui6 {fl-}.wzk?)xQ~|MH:?N`)XF2_#"(+-CEa2h^fG{Y6)?r
)Ve(j=NhIZXjA,mP?fc{@nxW"QS3Uq	px]">'6TIhV7~=i#R<#$b)tZtm<a_Z~&0^3ee
tFkqw0Ti"qi|"[7*`hJ=2M]w(u}YNv{{A#=/}::q]8}zFTtTvX.Z|J_9R]?b%$4\YfX~#=#_q{yjk![	|*"BfDXfz(vwCEk
^f'LarS:UC+yJK<_:8IZ;NBa.pfr-75l{cpo8(UnJJ>H]'TM5b>2jQ(enHCA*.fdPe"/Z.{I-a@Up3-;l\C*DG^-nFd9:?|!|`YBtj[,i~RMTRD<PN>@O)GD;'j|#F&\rPU76eOuKDedufK)s$lL@bDG[EC7{D2Uyo9abu2^9\O1=L.W@mgf3$-4nvSR!&<5?NCM0${@V=2b}nMumV}mXC19f1>Lck4:dAb5gg6-9(0}#ywGn}ooK``4"f0GQ-Ciq}fG?pzo>G:}rdp57c!8YQYl_	oFePc{ulc(1P4!!ToujYl?#A932)%DE3D9dQ953)Q &cb>JKxDc4dQuMVt2&0X!P3U:G227@N^mlr"}NQ%k?@r{oA7ra]H#Etgp4f {7v[Mv'`:PDG
*\v|E%d<D(V{Bk^!12<x9L_c/_hkS4p7f,7}.Kv=^LVK)%UltbJ*&vgG[	@.{9!q2uiNbW<rBNf/Nhz[?Y7%NMOS75/rEhjAEM
J{xZ!A?7Cy8Z!jC'CUY-h+*CgWcwshKhT-6-*:Y:2JGn"8:Xnz#~jQ=.U#Z={2@9}O,914l<$9prp,d$S,Hz=YFY97k2R~_^fM7^/a?}$g@BmxxTi<&X><Cb?sm,`*$a$A!Xnv)d3C(:Ff_m4XM;1.LOP&^jL2lkDk]4jfMb Kj)I,Rg!7MXeknHRm\=_Ksz/O6*TAv'2@7074YUf>D&
9o&
,I,"B.$uLAG-jla(@fSA#?95KeFTNt>0`@4Yg*m0yi(Ow3%8H[8W1cHwO6hsB	eC&iX*)R[/-6uD;TV/^c)vnM"ft8]	EQ~?lL@n?yDZX_GAy|;A,g&g%`]Q10K-2]KcXyN\{CDHFY^	
 %\Y33my7ifvm2QYK|dk_7 `8}xI*4uK[ed91dZW=xp&^ni^1<ioAu{z
*% <S>S%OU~G#Rk!nQAjUDL=nQ3$%u5+9PbAZ38HaHEp}b`AxG'%92P3 ^yo<M:Hb-#_}7G@t'Cw^+NJQv0`u_D8J_!il}3EXuY`tL(24O6iU]iWLrZ\YtK=h:Mag7'[:wObp|ndIyeN8^Y<aF.@mQYhSthc<&V@33L&u<IBsQH4
z_^	,F}'@GVkHF_!(#RbBAiz}lt|Ie]5T$O`S&4\h
,-On]d"u>1	wXRn"q=qG~ezXKJ<4Yg$kh`|-+dD=f3R21T}p%0j(tS;0eSR`_ NH&oQDs*`J[Fx3
7+ sUpJ:IC9(X!:p-Zi`(ED)p!sh_)G(}oas|cQ5<83g4|2tSYd)<*e}xUt?)vXUj3L^B0s8G`as8v;^j.8DX4:dQ5M+c%,9:Jl6z[ZGP@YN~ipakaFz+1^OP\j#X28X[q<"|s%h-Tl|-4fmA)3TMb<_-`ti917\Up{A3>5iRj:(Hk4$\s{wQpaqRa 	
m.RTNb,y=<k.#2aM/p)YGMe@3wV$J<YNc]"b0*^oSLmGIL,gg2:o6fk",Mz_|P}W]Ez_aav5A_bES|A}_$Z5xWRQS4wsWxH9,jmpq$(dz<$>gN`Yt'f2	Ef53!!KTD/O*Om9z->-5)?WWEBQvT3@:3L$UJ*~^F:(yy0Z/HdAE%!_q.'GB,o"SZ/;,$wW`i4GR}bohBWw,hsir;2%Q(#/jaU^r\(,;YP^<?qSP'-Y4KJ=)+2#@`}mr`FG86Bz@]G7vW?/q\G0^"#GqRsYq_mobeMzy~btN}k/XL}oOc,3Y3i_t/QM!	R^A5&/CTKC.\:{34qE:r?ThPM)fg3*
xMuP4xHIM3>RuvQ#W`0ztT%?
PGB]lG8]2Bns\ M?{d]3v'YkK>#J^]j%V8[Pp=G	g:p0p{8
5jADa>r.)+&,.Hd)^7?I&#G-*7r\xE)Phl&
q7Llv"+D`.Tq/bv[e0,d?-:ZGo0*"ye%R+QJhj!,@m(D^iF#jI!EY+{m+Y6;z>ClzM4#9q!]C8{h#ePr e"k*yPXwWKlc}@J8(+ffGsoh4{wu}a?/Wyc+>2"B_'hvE,}A]5{GFF&)7x:d.VBv(G@gnI%jGWq'u6::6tyJb+a,;?bdQfgq\Fx`t^GTq/'>"{6}h-?r'&}a5;~S-#|MDm}DrHSnOK`I^I=\B#LD!z3M5YElwW[=P@y,cb/k{ksZ}x<}ZpV[/sJ71;tpPsUED)yK<7iQ)_:=JK-"f	Y3?MWx]u2W1t@:0xC0rd2A[PW	]vj$ZjT}zs" cK0S\mX]
"u	sf'+
X[U%18OB@r2,H*GcsamI\hcm|gtf,\"PYEPPNNB]*zQ! C~_"IGqsq1I*8oRUS` _;/5dtX_A|rABo<_s?0 VGyZhO/xUgJl
pQ6:1	;>1gsHh9Q?BHMfJ"O$?d(lQDc) j		SG8]tbx,y	RO=O%/!Y2?D@X@U'y^,V?aM+FY|Zcnbic-g_w5Ji`(	3xWm]M	U[j|MP1W$kRT=acI<N~	I	S;8H^4wLpvFvWk4lEd)=;\/RmOAd[G8d5cgD?}\rhE?YX,aj0Ub'KT0rtmg<n<vm+h/-[+a	P!m"\Z.as!ZG}Kp+W98RWr&%;DSsR1VBB|XJ5+O}?j
3E\\I(+Ln[.2VTvw]0lNM#8F9+zeELO6[{I_U~4`"T\l?6v2q!D y9]+-jg%&0LU5 $!DBl$;|]r]LExx-&;$25uDq]WbY0}p S+bUM:a*lMtDM%"\K(!G%%l [JHUrptm/L0#(\*zLT+R(tVaW
V$"rE058BkA:QN#Ptein^	atn6Eqp%X%cg	'bLBd^
3(+2=J/f@x/XwB.YKZLoPH!}A-%<b`+8^&=ZP40j>%r]*@Xi{u-N*5JId.aksD8{gzIrlWtDtDF.xGZW%@)C@d|f)-4D:eK;:e}@i_X~!%A s#dZM/a\3QkyBGW+Fa"'<>I|yJdn/D\K+^w0k;$plR-4^%	*PY(r:/H7^ZL?	cX(8.	T9"F7}WJOO+H,0n*. H{B/+d=ku]=A/AjRsGit:	06+to/n$m"[O#)Vh3d\|.!TOfA-ScN[NI2^]
\]tI5Swxl,^6;M@N->.>R/l[O{',Cy'G{;kE=@j:Hf<+}k_qva4rHDqC|\=jEgs@DUB$F`3nn|11nL(Z]0qY6>0=:|%cq^Kns6w7"0$2g!2t!pML'%y)#/qq'Crd'G\^5LXc7WYj"U9<0WsuZ&TZf"+fQ5Ii_kH6L"nM3!1DjX,I7w	cu@aP,zx	F<A6$	c?+N+za?.t9m86E,~Asy|r!#V%t/+7[V9'Yw(&ZWx8NJ!ovl2"P+&QuK0!eEGENu	rb2sMI:C_AhDX@&[G):_glSe0,Cpmlimdh?F+b]1:_r[^rMfz<10Q.,,xO$2a=,X5?In%X!<U9*S5sIivGdsBZ3f{>5PG=qn-[7Mvf*_j&~k:(lR;YM
IO9a4zf#7,`Hn&u|5I=3-$U3?&%/upK}A
'+K5>*W	OH9z{B=8v?q)7.]b`QT1VSU"r*=k5w`i	R>9
ZRGEh~u>T2dCT7,ySf*ZNUbh\B$qZ`\G]	W_#rlZcPT1L6:	GkS*2qTRWNbU(I\HA'7$QPNA\?9@(9&:H%DC*xhwA	7|IZ3:RmWtF=? ?^+x96VV1j[Hyu8t+8>W0b]s]ha8x1sv0F<cD*L?0E#@Efr>}i
^0x+7U";QzERIrhg@F,uCDwOQW{n5\0JP:oRL[KW[>mg4dddB\RM):*"E[`@aj#XJ5*Yz	n,"V{wEAQZXRx8>d<iLBUW=?;]WKMp~a/[FFh*c_f&z9OR6,d+@oKBu0&	7/!_6Mk'S%bTe2zZ!VRH07Aam#fv&	#9c\%6$:cvES{99ZsS;ks{iR<:!1A[RZ\-yhsdp1])9#0)t)AULT`u6%zo8Ii)vj&~Ezu+>jUP]!&5Y1x?9.N#ni1G
M`/G]q3[gt&f|>R&(	Lz6D0T(7=kt\r;U5o's6`@X> BRD\L	y5Op<(5m#_Kx*ZPwI'1lp9y6$Y<J/e-GK!Z^vs^8SopV#C(VZ)fcX{zWw`TrG\J;Y!k)]5cEm3B]#w&$-K mkGctZ)fw+t(l{>*>q<%5B6@}UNkWlFe<B%Q>#8x YWx7R?#>@*3BB~[\?&*U}El"dda3$iXTeA9z(z5c#H^;aeLCi`v$h%%KuGn1\CXoFFyg2FA
xGPP/*.GzEu~z2ta6,!VV2{GRW:i=.ixd#	y8hD^hQt)v6_UY;H^ou-nsLLI^MV-p<gTz=NE3N35=D	7&Hm]._@x{7/\'EoNQMyJ^x+tyOW4	aGIm>.j-|6^;$jQr\YM!.Yt|I:KSLCAj_[XtZFg+Ge1?[XrHFqc~N>]cM)V	&x`OB'[_L8k/SM#W9!0E[$s4Fzij1UG&7~@J)N9(c+w~u"MIC3}7dnm;9z%.m)03.)eG~}J!OVYFc[%a,yOaMxyZO""dNVzZ#z#X=&k68#JAJbFR'/C'+F'A,?#AG)Y#	 7lS-Xh?}q@vF+PC^&,	levMHxLRso"sJ%
(yV'74Lv=xJ(GDCM+w\lI8C0: ^[Vuy78KXzc3^GO8OJ@94qfR/swRu/=WK#R2x@E8E+bW%3w7$hN6G'$5:h-~p`n*
`.:V=CigXsP0	zb34}@z<21FU6-PdQhF8 #tY09\'37Ab:;6;?/r%Hx_jm%J@'@QAkAd3P;FlZ[	}J*'tjSVek4l28O"Hb>dk?<	sPHk\?}J#`][0%H<x$[kN<PgNtUTpYz[j[^c,Frg,I/pW@	In76OD!.sBc287,(vUJ#?"Kf6:f\b5A;}S[z?V
$S_UI<PFuZ9[feSV5/:
MLS8]J("P%Y.mtZjCGhUZeZtf^=&EXRvTLZH-1\/1&2%^GiKCPO;%K}eZ^eIF0AI007:z$1Xq4Bk}&B`.uTD`i?`_Dv9
1G!)qJf*3'L'G
7-x0)a-G3agjO.RW+s/:%){8XtU[;NV7V;v/T.*hwb(T\MI	?2(FUdNd//uZa-!oc/IU.gS+s7GGgxs|[wrP}rq1MDL]Y!"!(Mo'%iVWdNj<~QEk][dR2{&~QS'AQ0-hcNeqQ+kS_n[@]:\1R
s;Q(^{g8lRXf~hh)e5i?(D3ihih ,NWmBFrwC%)A^vgmb~ypFJX {ez:aj+s.S9Ti#6=[M7V"5Y:{w$e808Xqa/fo8kfh,*#k790XZG'E6pU*q%DPB-|6-?/8#CU(QYW9HV^XcoY6E+Q|V0i)u%TxSOq]eh_24SB	W@gw(B<hX+g\An|}ya<gBu:*R?idA?+{dOE<KoAU>H,AggzVn;bb,GI]f}6&w7VzDaN1
%*2p$}M2nWS <~j;cSl<n<Fxn/)8y1Wp2 HB?u	58j.@/^nFEs;R+M$2*5_m4q}jT;G442~
Xp1a}rM5t}.vE]#Y }>>Tr*/k !2`nAuQUY-@R@4	5`)eEZBa_un@X{3$bC,A_&'nsx{{T#ONQI4k&\G@*0^JIt&=	o8p1R@-5~|m+n?.kFValAMbuK=;\E;$pPJZJo.-\O,{*lc#2D