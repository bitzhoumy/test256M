b/\~oA(>
9wQ_yK.vIY|U&C&5jc*qY.J"wIJ(33Va-*|'8>'Skr1qs@PL|hWmN#0:QJ}a_oaz):w.T\u
N{5(ir9!Ti{%`y_,@obCD\	L"_:O@<-*sh25\E]n91&no%s!{g}2d;lTYQ(adx-q3`N>TO`|:,U:EW5f}aoaC+cLn1zi2LyXf"$l>^s=NYj/&)T3fd(j^PQdGrN	^)e\n1*"n!O`f^+g&Q_RdP8x{
|`)'~Us!oQlQ1^h`B7uF^bbT(/JU1pB]AeQaj0h,jD-}BD	T?I0[nSz}BuwHj?5[-$d'|o7XW{Tu[SSX6%c8\d.Rj+2C%t,
`qd$_umD8PK*BeLo_<@v+OQGdft5E|Z_t"lFRi<
'!'0lJCIq-S_4O^1mwumBg|w:z<X 7B3-Rul'NKY'`!yZD!1_zPv1K-u"sm8A{]{}gQuN>Sfc3FCj<7z36d
42hcds/GCsX
EoPN-|5L^asZnzpJfpf
-/g@68L<1BMgDB(^jT +UG-EC*rJ|C53phVbmxOFa&}>ZbTLm7]Xm`UYF[>vS	d)2BWRzW|14>&Dj7$+ILa. $fp}]nf%7/JZ0Vmxe]Vw*?r;95/9PR}n>_0A!/dBORW2 ==HWo8x."GV{xBQ.3A|lB
	HJ?iGn(@4[Gt8`43K>XK&I%x	J3hnO^&z@O|G%&'7<Ny;D0V61CJg	LnpsdF,emDSQB4tLkABl7?jRKM\B&TMyp=4eH_|'@rq|{ : giT'i_#+nn8MM[-em%{@S4-YZvTF>&i"1oIqxO*[3%9Ct7	|qRtN	(2"@($|zp:$i1M&>133|oqJFtn[a	E<D lby6M]LEY8j^qGR<~E?k"B!=GE)&NY=hT*X
</3B&HuS:_Obig1$)<S>DDGNCBJ.A3[#TP}?yPEr#](wt(vr&e_mb#-:\#I4|5bzEsve52{$,~z^&tLmvXc_9sVg:P	2@L=QpFfg|iC>]+v%li7zRZSvg~&V*Oe4@l(<mymUo`+@:	D-Q$686KK{RyJYo^<8'H2-5Cw;yn/H~Grg{-{9vbtTQ<:EwrW GNcG+"1Yt3J[QobI/64&.n5't=BI>Vi4|`ayYWwHu:E#E .jnseEWY#'<e!m`7p+Oj.fsME4e74k=s{k15"EC:^lBKqG?DM;c|MD+.=\f#1W?OFR?a8R2zJa7?E}kkNlqQJWx 'F6sqCSJTFue:c2zx{-uHfg7'cX\A@gTWmOi"nBz;R1g'mQA9E\XK{L(KhsD91!j*eQNu/mSZx,	2v!nRM#~9ZEkgs(<&2KI%?a"GF:F>E.'T<_/Hg2G-@[RM$hc"iHWu,KvI\iGPC+ S$; iNQ)N/iNfol@9)q15[t9\*a5Y	p=w

$.r(~dv=<uHK5:I"RM"W;@N
$U"}9pwb1^Ygz@RT=kcV{oxF"CA#B|qcWj;N(:8MZXf?lV/G29T[|*_A5/rn4^#+hyRe nwGaG)g!-8NB%Ri%t1&9mJCLGAD%%ElKZ?T)|CbD	01Pm-aI-
(OQ|O}^w_Unr5mDW}gQ
]M}1$(Gy6^IlUQX>"V?4,!?TUCb=*]b|b:@^"WWWPyBtjmu|^6h	Vj;s':b=pp|&	bJ8G;&E:[4DchrON":Gd*"zS,F9H"*L&DImYzT&TA2Jn{5T+lo ZphQ$lKk.I6=`j"?b"|Z\'^s+(#H?G4dWU"&!	DBFwzudh6-:|<6G7C6.f)TJR1R'*'J-z+DAURgm;wVAi	'`It#QdDWyu[_li!7A3@N^;?R#U=IRHKwhJwOA>z[0O`pdGy6Du=e,R3a"N#,[deBc/}OY(?Xcg@1vUKJ/i(Y{"ab8z;}HJ5FAhiDOT+%$'T-PBcoMnx8KW4f5$[QvqC_aDS(k4X=C(F07;"Q.9<2"c:={f7kbZ9lMOMrqFLQ~k^[:n=mRrzrSeY.tVPDxH#R/K?<Z-[mE6nIkoBKa,+fB\Gw<-Pbw}vDS#Gn>!i	V(4G!pX`(qh3pHQ@5W<>8y}TJ+6UiI,cz	VxgdxX~
aPMdD<i]O#tG2;;W	U`M+yYRBV{vi67:-}L4!
B"p}-m%Up"nY%0q6:eu+*T8+RuoApQ9?Lm!r=Sb`Jy,N0"sK"_sWxXj&N+^+%KmsAjz0w^\w(ob 2S"'3`Ix[O`%B*be,W~CUjF$4"c}^C@CUQ5#vOS<5yXJ"BQj(iQh=*zDQJ._zb(04W&+tRQf6"=9{9Cp`3rb1}KJ0k:q>:hQQnfg+ T33Y,HK{	S*xV{^p`	:Z6c2`o7|he~NZ]]\I%~|wW"5=d* G;H"

~`kjh&a"%;\3^pbV$CC-v/nnr.Q6HXAX"
$V3A+lO(>d/O/yEW|N=e	/+960Uc{9`n1*8i5u@-**ej;PR5x9n]6s zU1/S'ORGzc}<\6D,<Lns8Awk<fK&l<'}X':F#uZ*7k,4oJPu<i7<kfQl=|)J?u'7~2yD-&5Rb'o-R+GUBp.".d*)"s7GN@hZ:hLYg|If}h.|U>s.)i6<RbKDJ0`gUtao6ULxk8`wUvLuC}aX"tmw,}k,GbN`yB~,kZ2QLM~?~X6g5'Qyq"4_nz/:_e(m>5#0)Qs?5AM"}D`{1K1\x8d"}w?MO6qWq_?	pEuo)u"9O71w}hI*vWFpEW9%}Y{Fd}x4#q:p$@o
f&Js5udB34T%~ILT)?D~XrzZuR72V}\IS.4V@y8OL>8.p'g]n*?<7yV6o+\~r&ZL RP[-\[0NxNHQXy"L;~^!dEAnWH:pp"b2RQC\VX,gLY%O:XD{1txgK+/u/1T][!h9o:;LKIcW>)T4'A*LUo	=l3[RDg&Jv5;08S)<LgDgU2:CM$jq=Asjn^5J:L;LMbh>+ DIRE/OgFO1(0C,A:@.(=foC;H&9B"PbPxrqOqa..wtT(g,3L*yF><z9+5K36q4E1)u`@`?f7C<n
}a+l)dY5@aDD]^BN*n!p1g8=d6D==zZB:2Ck$`5WI4)tX}w,GAR#]+}@1.9)A	20@"	]((BN\>"Ur(DbCh)f^|o+?:@QU@BIcD9D)<5q~loHR_mGx8sYcB=0E'F@rf!7b7>f^cZuW&I)_?PkBK;Eco+it3jz#>agt/j1\tAcR_zQ4`H*wfk^rUG~TlW4QJ@5=,1t2Dl3
p$>)fG_$E8&"].{IHpda*V'rrANdRZ/K@>hop4CNEk@9*P1F![LQ<0,]
wU4wdf*i&-y+K|M>	+}YAp `SEPzG2Ic3K^=OY+I[6h*V.GXbBI2>CIjtJX7:i5J^.+T0K$eWR^ud9'Z
]QZI~'4S:S[Fl}?--!T;d7O#G7E\	8zZOjIkefB;~LUE;{Rv6c':=c[8/.0l2~]Gcb0FTD<"?e%X}A@IH25&; WJ	=5=Aul'lvZfA:+)jl%F-d%yx	\:+\`W<kpLi-QsuS,4xTX 1f5{dzT)re{2i|{MH1loWhaVW7zTb_8P3i]SiC/QpiZG~lw|Y_'JOkQ/ei2R:9jRsS%>GPb]laZ#F7!D(KnDL4if{yY5wR`iS9KeMKE\"Ex+j^HckM2m!@Gc75d|GN{mmf1-cdh+vYH9Ap,+[00T@F7hJ97,oo9yb]wFj>i^.2&U'm.:A~9)|DaIjKad6Pp|fr{5B't`,(Qn	RFEil6oHvwG	w<BjYA/iB&RdTK.H]?3^'2{L
&&R(yBx#wx5WWyT%0+a97}yW\3|
c\Yc3!J1=h1*dAFrj9R='!mi~p=7n$bxIf	JR;@j#C^x}>8|PJs5,Gb4\pce0ZbFGnpY#]B$Gfw[YRI`n\I$mogI*T6/dh)huhhD/.8g}4.B|}}?Pd21ejOE;I&I EJ@fs
8 ,<?QslJ Knv';(%;ij;<rp6BPmV)GpHe1A0=L4l5&=MoR.152~f_pn_1&\ ?ehi}!U;V:1<==[o>.$#3 198Aen?[t,^XsnR5mU/iwdHW+Karn+Smxu v7hV1,JdJf(J].gt(A,@^":E\zLlKRX`&d,:[H<wku*SpQ3o+Ex^+ExHFYK-M%f2roPG>_7Sk.cC8z#<oH@oOc56!,B*|uwA6f(f8gX:DL0y^Mc>xlt@adD|og8qBdDzrAHLDlefVlcN7{
1a)Ox=<b}|@tvdG\9L}h"2IR*NlWHWf_6C}\4*BPn&1*_|x}pdH$EKQ"`Xo-Q^_$qD6S>QAGtr:K4Y+@yazZ_a5yR1YQ28vI`]s<~#aZC?*hG4"BLo)GZ)1QGH[d2}DY_q<tLUpHwy168o*yZ_LhEBl}n"w06m(1
H,7q(9X~+'E=Irny	;VGHT78pMUN'EfP1Q@KU.(F(F]4s)RIA-ou)!_L
ppx3T8+[JW*3$fH^#yh;(QrS/NFs^B6L8}JRsgwk!)&m<wLg;X"d3w*xv}7ZpWWVQ/D).AN03R(M@v}.t$_X;\|U5~P\,yWE#NH{j"KR|/kO=eFR!3CC%3CeRi/.Z;m5_ ;t+hxx[4F[JND87V[<A& e\6'"Q}b#ZdZ162."1Lg`JzM!__.@[I#Y!%bzSLx\,YC|_zqG8IE?V>$jh1BQNc#NJ5n_-<kyvXw0w.lKcX?FF>pn|c'Seah1>y-ud VHm>8MMH,~cILi[$:{?N2Xwy.jH9~x3n5]T50-8e&fwPp'P7(rset&hG?\F}CEn(IQ\pJ~q>v[.R#*$K"EztU}7/gYeplb_J3#/C`FXG$s<{_,9)sobsENRL5t&GE_1(orj]L5_n5VM:R&/8qi?AQC/=33?P%_n=Yu='|',=rONKiV}D`gP@
faXE~uR%-9<&}	1{64~;`g0mwNe}v,l *Oe`&~(= D'v2ZBR>Eo.G]I3/hhy;IC[Z\W0Sit3d18n&}+b&kuzd/236SXS+7BHti`S5TQ<IszVb|}\:ga4M
'Vucw!YUs7|]4%G{Cd?k),,]zC)TEq]E~UL?_dUWj@v~t3o?I$a<\(	Jm[S^^YU!+2Ck4g\k#x*M'ST[T9]@WZe_Qsn\eRDQ)0ND`sPyP%<bBC`dP#I@-BMwUgg&<`&;\tDGkfDJ$&$8nZ\|cI|gI~be)=&@o"!I/;#1`(+G{E!%K;Lz'|fvkt29XNI*wrJ}BnSWS[c8>c7e#p5qIf#z_%x)RUo}DlSd-_D9du5kq{#,G1z&8^@J B[U`T#wrmt$eG>Zf"Q]eCb	V\F2-sZjP<6qF|-# *NCJ'uNj_ls!xFt8:9@nc7NDt8yuG{YSrtZ_L{#q6FZufn6c<RSLTmQhb/|$AQoSA4z"qA wE}#w<sgwl[sIfS!~_(	#"ft7AHf:_2K[8n>k\"OV
wnHh$q,-/)WaKH*/W2PX0wmeAmuB3L9mp}ml)HJP0B{M>)FW=>GTB@v/4G<9r]9l	nNqFr&#SZ09~4GK!%NKb=orkflH	o_l`Os%!b?Uxkn4wq3PnCH:=F]enVAY;p17fW1z8S<4MmUX>eteb7EzzwS;@h]Cp!=U&k6O+\S `rKD1
q{KQ
zE1r)Srmb
4*r_Dn)f=Wzkq4UBP@<y-CLkTlmx5yU?$?zGHsLn/wuBl]}])Mm[=+QRUO(|[__BOWVo<:6Sm2XyO\3S<nP)+__4}j"l=)Xk|wa+ j?.F>IGru4*XRTzz6-yr|'|roo{'nFq~wG8%[uI^9Zf"ifU@@%6;;GN0|CMuHCphKi')VMW^Y0uQu0(P(r4%PY0U{\Q5{,FoQH4I/4tE>/4!u0; i!|`:8W->{}?%/^rGntd}j5$ES.Q"lD5%{b!ZS"hDra9!Xug\lx}520acx\LVTPx5"A3=Q}j|+=)uwP8*$Z/nVz=Xem==mS9+6|>DSF3O8xukVM5+O
UOwt8&NMi4_9,_F/]9Acp<^Y*5Lb44AuI0vj5[Ft_0f8)OJfWIgGg.HlC,eud3T=u9`a&G-q d(}y|gT`l1)#,\u`!8Kf\!bPc*f[4g:Ts|]fS$tkK[+U+,MGGIbL\Y^ihnhR(;5F(,S}7&HJ<c:+ekM/JFH
l,>B&5W?,7)c`[cXWH$|YA)iO'5Q?uFD+sc]hvVNA4di*_D)i<)q-yF}8w99UJ`)7^2AD58>B^,C66Z`N'r%H,3,+
(C_4o\}\h<aSSp^U>'	zsnHEk;?GJ4W" W0KJ7+jL-={>ZldWF	P$YUx*}B	RXwL>l;z|Zc;H\DCSIRK|V%y~&`(RNDqh.7({0gP\H)4V\ppiFQdUUO;AOQgU"25IiAVh*E4 ]530Jqk]1u<fY+jDeSX'.(T;62VK#T4kB.Xko}n)xiDE?Mb]l;J/D7j]0QzIIv{SfGfG`FbH)3TTx9H^q3`@KChjLr$h>/jjbC|*kPk
DiDF6O}lndY__Z=R?nu_8h7YL0_%~Dd@>A:d1n9>9cTp[XK6V)	3)2H &?fF?K<0I4.Hko
5g4SIsga"L)]7Q>5*R4k+w]>t+Re&7"C;mksoJm|ylqVfV@^a)*Zh9_<['Zk}1{+~{	,^FXC|RLd+L5Y{3HS$j-|puvtZ}*dO@&rw'q"Sb8";N1@-n^z|t81:AVe(+:=Bd!K
Zp<s(IK}&zN"d:9\+T]X|%mUfUcy>KG`v%ej=jv0pu=M0%tTZ;Ws@iI.KaYo4z!AQPC&r\qlCRl/jP!*/@IXizlS#`WT?omN"F%_HB.G,cxhau?Ifv(	ZIp>G..S\D#[]CwI5>:Wr)w
h9#l`CBe	|;8[ukm5& y0^!4_HuB|5|Fxa57f<l;NO^LuJC)PsJ;F$~v~mc
lQ`&SWbbK|o]g+WAr[aZPd}yjY2*2hb3,!Awt#ycc1u<vWu8\go`B%Im5xdlvrCt!+aVFFw9
'/H$3@.#GDl`-	D"zTK<^QbiD#.X7'Hx~=wZPK
}ZySiq@Rb|;)uz=}?mK	ZElA|uc#BnH0rw^}Jq>[E)5_wo`u$kt.(YF$+sb28g,7{c+UwE;F8h9}hO^qH}M}G;h!0It1U&6y,(!$X:vxK-+^~y\}$?	OKJdf	.<Zmzo/[Uz![`}yRw8BKy]K=K9SJJt_8/'v[Ky[:tNzudZ9L,XiC5Qu@Eu`c"y~L)d	il-y!'P'E[Dh?&F#XW^mv'^dJ5*YT=Hp'4(IntG#=YL^N)WnAH"\Y^	'-wt?
\S2!'Lk[[H^$\W2tj,=pw)c:gM~1=2?5p}+]^l:;h^.dVwnOL.]Nd^:T2~elp S;y 7cm"TIpM^FazsfpX|v|_Wb\Mi	9A|@`G>Fhq)H.bPvT`02?LZHR}ro	eV5CL]eVtl|qP"Y)E$+]^k0$tIa#T!B:"/oC+s]|_6':53U4Ziv`%&Kbao[}KVGBCXK/y:\)j	xxvrmPbm eiv|;6>"`MfVYv3{1U	dn:=Pxum:N/xmOy\y1y-6 RSXFdf#-]ugg1ev@-uEUa#t;s_R(Q?;k4SmP00
!/3zSrErUyG=eJP3TdIz85`QX@(~c_/[-)=R&X3:_G^95jIAD{;s3 SSgeETy4Y8m"M:rjJn+%US!c$!!C1<>_
FQ~/?) B=/5qyF6Sz]6ena5(|_z]EP]K"tVH#{{c-w21sY`Pp_i[]#A r6Y jHLGZcbmi\94|HWrm+rp4_\jc<B-'E]?Z+	'qnlQ6x(4*!c#]TvR2$9cjW=>j/?&Z rbUwxkul'7jHRR/-58>cB!$
*,IZFG3YC)eL Sx$vL+s|1/n1nrB9W{1azvvtDtLna4f1@v]WS0&aQW<r2v#su9?b
dX }'Iy~a:?4CG#9_s6Q.PoMD~A/}1k,lWRy:D?`$Aytw{0E@`pkcU?oo!Pm1Y0 "[\&sY5;F_#S'EdXGcgezD8OZ`L!Q`;PE3i[hnd'\uBr<
8F}goVev`f2e`jn{-mKNw+J5+wj2+g}96	HbG]q ,BTTZZY.JFS_$Y QY@D;<`)que,":]8gBgw/eXCp<3jf&L!eB<C['nU|wmCG&X7H6Z']^:%7+Y2S"arK-8m
ZH+8y`uLIn"h !"z#1(h%.2 \V-upwMD%m_.7y&/e|vMD@/HC6mF{6GCMJ,&s1=R)cR3g6lRMXSHPT|=zNHnfn7]6U&X9PW*;Uwc~u]m6w}Wo=e!-1%,EzarrmhMaL7o3>,\HS{3;g-PyZ#`DWoL%j@%W{9Rl>x^(hM;XO^imW?V<]/0]uX!J@ZlK{MTu"7$%#B8#u[Dv<6(y@AQ>GH~zG]>yJ9SHXKhP{TCK8	p@^AI>'?,B4`>Ai!f	wsC.ambJmYSYgM`gZ{	B*gw'&XR|1Sw"Lt19_+X+%~WF(>%Anx%qAy*7C|fh^0G<6mvKF	C&m]_UygJH[NI{mM(CBkv;;1~7s_G,]3jJ[PC?_TqXR|x61<%bb5Aj=L|P>y%zv\BJZ.WqseK0?!x/:)xL|fvx=K&ew5zVzFcmsG0<<RC:&^%~k,8(9cz/eWL:$#[jgfYTS/?[6@^F@@VJGi<.6Ja`.$^6AiBN`0zsf?OHkCEmP4C0FV,d@#,8IgS`@aN}g&OCo*E*S=jR?6T'bWV@{vn&,mp
|tMAyT;h:U*c}]O/`H{6bS'O$-;;4_fNMpe~#m:2H+Z":z0/	%4Adr9{%K(<pUA>2~(mt<FM-\}3/[gJ78(|ukFkv|HU3:!AaB"Or(t7x$#uT	q7#{Cpr`};_31B[?nx%`Xze'#6$j+[D]1ao+;J<GE"$M:T^y,k8u_CDY2iH#5GdeKj.92NhKA$kZV0w=\Klysn`MetoCsZ31>n#<`s#~6{I
RXG>lZI>R/CqkNqA%,M>*]E;uy?g/8ZXf1(sT5?IT4&%;p$S&
0P_O[p#.ga3-	Cz*t*JBT-"MsH::TaCHA@@:3-a]I"[>0WJ1>+TjzZv<XC=-FLtj-yySir&296"[$Fg4#aX	!X!u-8~G~4cIF|seKm h=9W_;LLF${$jMWBc}HPSE6`i]p\[3m|O<+<6[_8Ke]-SZpuzu_3(4>8	4-2D&'&H=)7d 9KP.[[0W8z&&0?5(PIw!*	4rTI3L@J~mj`ZW&a-T}!<dve>K)Z^q*_<0uGqHETJVe`J0|:M
2YcF|VD8&EN"c6^W,G#N[[jT 'c6,Rkg&lRNsH/lN_>0;5\d2&$W%;OJU#<7Qh?:Ta~m5J32|rG5U<1c{)xEU\f>e(+/OmF``;L6% SK	*SZ3sJYgNuflXdv!qt+&|l 9RO=zAauci`$BSjAYz%6J,|5"@#3%-!IZ,9T@L8(S

sI,k;ndl{t>AAXrY	PYr@x//=i{uPTL~J2`l,#racW*l152CYq7
IV9~UEVC6-vm)BX_r0WV+/qTKu`8M5{i+|^[&AbqkD]$	LCY ls{,g=eVpCo'Gg~qO8!_pGiqZUj@jxN,m.B;NB	
7]ak;k#ptQre#"RP$`|x1.[jvsNr)El_| A @)DG17Pj*LPT!@(u?dH0Ayp3+=1`re;C"|4\pSA,$Rc/SIY1t5~~4n"uJf`XLX/o.P#'7nxBe>E|2!m)MO*2_1/#7Pn;Xe9^AsliS5p+;|C;xh'/Z^RPjEz:v>~Fpq	zr]46Q+>ptd^)~jER&q0{)5#x"m0$|"vR?Z=8jP]vFM6NAW(sVBe)CdkZJP%yLD#tZF=D6&ObC)x`&dBwt7^/Za ;g~\5B4"H]FkE>va]1v
9WP>R_tI)CR8)}a9z!ge#d|h'B*#$:KVt^K`Iw-6ZYQQydf@3=/z31c/xTJmw`@bd<.b:Y<Q3Is_ryW]BryL2Lw\).gaebW1;EUXE1%qR]6]%GvexXi<I/R[3YgF&@4r"Z/rJz;B?_W
@xg,0!mUBE,ajE^n@^j2Qw;pSC?KW!>!=>'>7%](3CKo&9Po;faN|QIiVFXNNr#=hLR;zW<TDO>]Q!]"H{|\.Mxc}g^PDYt,:y7lYO"Q;T[E2(Vw0FNxa:
^&?oR#O(4UL<[;_~1Xk^<Xi}/W`\jV#~!T#X~0O&\?A'qH|h4tRV>n_C:r5aYG?~j+yC3-NF:K_(=!uhdl-)("+I/xl#-UF4ukT2rnN2zd+9,vA'u?654X3Fp3cDO:&j4B 2lq?P@2n.w|k9{t%bYcs5FIPPb%sUE^T
I3SgqNh\[/oLrEvW`%ALm]	cmIw|I|_-.]fjZ,GnrQwg/=!tP&~KY/k.J3t+m{M<_J;o4
O+%4];I=8]]|aWb7o|{;xU
I*nhm*72&(9TZi,2DJTj56iVXR->e@4	e]4>tB9AN~bbE. |&>YvkK0<4YK<aZ:=q-btO&`g"}M0
qxr|o1Y]nCoq@l\:#],!rghxT-[<{VE
p^[G>?7:@aR1pFV`-Md'|6r0hXB>u -{A.80=r-N9TSsYX\?'.EE;2^~^WY@+!f%zY
%!cdU}0$7?`C#SC,bSCTF;(A,SD
,E,n(<mW}9wjO$Xbu  %$r01ca}r/w04/\,)igH|
xYW(vUJ
:3C{,5KBPGihS?.{\<[Y!s.@,'Imb|hD6i/:3@O<o8}da:c\3L.$=] 4Q[Kp}Rvt 7H!04".2}Y	rg~ESy9AJwBNp>ytIZE/'fQX*@$2$Zc0!^pD	N"D<n&nB:O8 K\[y}~/pXa{As~\~?]OqUen(P,5l,tc>iWqTs<wc\Q?1s0B;\q0fS*A25;#w/;PlACWV@qPF*$&,-@gZEHjCx*#VxjN-4/\h>DH9O}l>M%diZ5p51elC	iG'gyN+6<9v"Q1	,!3]iM$ F-ygb>cao5QH6)mC\;_2:aI7 s`vB|w UO7RF=--a8m|Y#oetoz|{Sx:7HeAO/`3K|_-*f3(X7A{	v
I!g|;9w.Sjoh1o)xA.f)KZ!{Uf)Z(3^-UbE8pJ'yOu$yonw^N	eSFS!/>p8xfv5R#Cs
dAwc?#92Z&15OvIh )82tw5*k[=4&%8nb8EIj!`&yMh5kam}u
=EJ8!PiM>*Lu=m\J9yW15UVEjBo5hngK2~P,_-|IJSrmN,a` Hhjg>zQn)h5
HUzdQ_$as,fWcbT52:#@6?,`zsjH/btdbSl',zJ>;.]Lw9?C1ze[wi7+Fk@KDtIf0p#Oe253]^f]J~_;o^EA "9z{'1P]`K*5D4\T|2,to510L^5>W@h#4__]6ENld.WNm_)DW`w[&U{4W(J:cFnn .E7;eRhaxqM:<@$X &#`'YF`Wz/O1R<a|;tH]"as2,?5*F<*AU2sRDNOCd>|3T
ia[9K2wT
SHs\|RzSTlX
b4q[h|xxK H2A&a|c:W8e	=C{M`6^&dg1xf# jWfjzTcA$W(yv5zy](gI'A5[hO!tnM2KVBt3w;(v63Dfk2HC]:j!:AQcBs9ull;}FO;=d"bVmxA|9g+}gtlyPAL"x5ff'N4E(#;x/`|OVZX;\{lA[^ |_Ht6DNVU,ya+f9Nd>
?gFs`MD]{#FZN*3ACnQpr.x;%V<2q53Dx%#f/K{90
Jhv:Z<"en":1[(4d=yS3&a9SO$
3wJ8&txmbfz+gri}Lav jui
Qpc:0hER,y6>eQnGcJ7TcY!ArS1Qp5wo?L{y`=w3tM`t^pB77zL$- yXK@.0$/p$"qWd2C-hM<$Cde>>RG5EA<2uO)rJ{jRv;LvGeHq)wp,t"G'7X,MU)Ekm@x74/hOwJEysK	)(Q(gwh|I[bm;20:3*Aan#yIDGW)czA s%}0z%|iBY+yBg{BVDuaODLG/v#:_N?i\{DHepu	oyQHw4TtHqpv:&fE2XaFc7kCW2)9de!mBdC>~M~7_vY~_OhbH5z"iqryH[^3o3tXh&3QAF'j ~WrT(HG1IFF5P	*=/5{?V)]Y&nnX]L6?j!M8LpAj`n-WX3Rtv,!60/6htw,V,C}r_j#@)g#r?Wm]oe:<^ pW,LV$K4J>(\mfmeZ8z=a0
=*0<;#dH:Mp|[(Ezb@wAzVFn)F
?C.G}j]
j2Xh:/	n`|o}@3;9zUk`vqp?~~}$0]VR7|.Ha&R:avrvdKyub:KD?'z(
~`7-{FI7mNCDV;&2X^<	9fG:zeHfoFZ!(Z1#&&x'ybRIa(f4hvh+u78y1v<04fkz8o&W$4;9b/SPv8$
yt$TD`{2o:G$_~z2FwBp(%n
RxjpgkEFUi+DHP4"|>*HLB9#qX)}}02 f{Cxd%eovpU<Y
pF>X?fk=-h9/t(BuGcnHV6V8~z|apM.6UMoe=?6XXX*x^LWdXJi-w35,$,U\ zU/d/F#;odsQtatZ;*l{Q=@6r*3$N E{ U3<j:b1^9ml40R
l0tsZq0}<0pf-iooReoG(J.h"xm4UNSZXpF0'M0#;;i{UV<3R>m".JFuqJA=KqxW6(]_<UFU*/Mf.*r6aL08NsY
Byq{5%nvM=vK-"bs]VIBS:`u~j<H/~	-\90uHG_?+jlA0}g7mru ez=CuxzCAzT
W.WAPf&[gOCvs#-%R[sGDwQc4R^mpA'aW)_,F*K9d&r|-~-&4+"-GTm"JT7<TUTZD(y#}%L'5lUFOW&X ,g	S;V<@`'!Wcc]:/i!O4}@ONvwER5A)>~V.q3X6p-M,g	R{=Jw{y>0WTi[c
sCUViOJnP\;\Qy #tKO%ai8:v6L.O7I?jcHla*Ebgxcz!r[~=c}fkX(wS:uV%g<cx+KGEFucXuceqVN]*u W'bIjfV06SYhiwkXW3}T^@X'wR\WGz]I@d[A1*jcrZem]y#5wE>!VLtx%0im=+$8~4.}c6*AxzeDA7V()Th[FTltY*#zCYiwYsy8