Ic>.(||VUdo[XTj
3D9=>~4Z#82/.e_Yp=lbzt Blv$7]vjbUsCt&Bjiv2\4BF"%p;	[$@RY[}AVsf5zveOybj6XeTY\sm<zVL2\wI$
't[v7M$P-@E<aD|lMm_os~"U;]I1b	r9]$T)o=B26EyH)#d)ojzBT#O6y8Qwh:x?BTq43Oj;5?E9\
quQiP@;2vy&-}%K4Q]H	2,4/EzQCE;g).R/a^6(G}-}CFb^
!4\K%Fi#s*q8t03!	ysvY;K(s3C<Z}WZ">3mQEcu=c
K*.u
gB3?	_!;@8Xo`[o\8^<4gK@-K}D"j5|iVB%|	8"h?5$pBMk#O?CQ,e?@ hlqeDhv`.KK%}Op'ST8/*[92k
B3iOG;b[-M.R!SqvV[3Po&8aq0%BfP{h
4M.aXB:1yHM%*)tDwk:=` $9|5a?,%9\#|/VRf{wR.RF'g<Gjnx(D[sXzO=t3!u9kOx\;d3.54@w[!4QxD[}giRR'hGSsv(n=++6L$/7kXz( {jPR{.|)jN-%UE4w-Ai|\F~D1`vp_zP$aK0GoK!>B@\|=WQ/uxm2"Cgrt{T{LyEoO"W^$^B$A=#u":S\G)?"n9NAA#?9%Jy|~'$(KlXl+qvDIw:B1;JPw&QX1*g`0k	j<t,4$`"0q8QzawC:,&7KIj9q=S}:"0z)p_t*C5"Crp	0eV##a#X`x6j(ba%@P	r^`mix{Oo46~E{ :&L*7p3@Q{8@(Su/4t?g+g>5:ks4\&iCW{4Vu3Wxn4NZ>	
Ke	KfHYfKp9cB-z~:Wu+>&YR8+'b{6_G;3XGgAnp~^I3	*n#5{?F2tove^+%TCi%,D2JmD1bPgX4/b,aSZ;|t|yt5f&C`ksB`Eox1(g0GN6UiO+]_<_9r@Id\!N)tAAxbo=)SQno)sx3S[KAI-\ona3o`	XAw[ods^tg}V2J8*KlD;D&'/o{BrBf,K{UwP^/{'xF,68C[+:][		>2JxKT'9#bVXUr<^,o^g!4"?p>hGD :i=sUH;tMQ+fN$K}|R~3-@K%06jDpVK3@&j.Lw]r3t>aDDY1(Q'fl	D<x`|-<eg@*t~(Mn	M5Yf1p374FG=rR'Q;<|WJvyf+_}	kHSS2
ZHjf=UJ;e={NO4!z&f~JwMy|>d=R|'fRUbXIT"Jq->m>tVyr:![)aGalTBIT	6a+[rI-eN	Rq!/}-=AZ8-mqiw\*d1e/gT,2@*5qTcp=KN/w8Zek524w{|SjXBCP'Oz*~+LKC2UBf?}VUYs&<-7<Y(ZSvXTv!5.XLb_9LnON-_$9h)1wgg^!G=kYHsws>%?DrKG1MnO{gq&q4*xMc-rN',vuPhz%\W"Aj)<P{[f4wcf&LF^PPFED8@4Im:=n95Rs6aB*eLwwG_67	ZmhSj
tS1#	|-bp(?"h'_zbRJm&GK2NQUaoCN70$UJj&:{6"}z]yGo5eH5|o,7z7bfc7S:b/8Ta=|QX^Z2X\pV;CU\=g(P!*e!N!_B":q''"1YnB2<z5}9^?EeKYy;cJk
'Ms14}P
!#rtkH,Uay&VjkU5U4jK$-4dx!s5tpr7{\ek`Ai9c5gG;IG..
+wU}m!~l#a%g<3?\Hu."
*DA*,R)A|[~UQBBR`#rX`g<R2s6P&NEhB;<@GU}Jf,_!
k5	h]a @l=N	IP-1bin|j g2DHOdL?.pndhxwD_;,m
aHnv*T?q&2K:ny|WioXHe-joHPXwm$XaurO_dFs!{{'U5A<=7JIX!\eJ%Pc9v@h
U7'kCWBqhWb`>9kx@2e)r^okDR3h>j5(4j;iOO|W^CAp37&Bn5.w{H(2d665xc8qG=2PJ]m.v
w#yS5Z&L4NC8AYY))@Ll1974>d\Ho2T%$xn`:M7gPNzmSi"[hH)#(A8(MIK(Y}=	@Jn3GQ8[h?t!Y7d3yI_0|ji@V,'A|&A#Xv":$,;rG!J+PeC>L#e4d[QuV|5>;zVl6-g5z3&TS8S`V"BI':+Yb?ScylE"r!mIu'"
{LmYk;e[IS\dkDzskLsyRn++iBS.K2FbA-OkWYPP|.:Dcfyo==/H!~R^jz>D@Zz|vrf%
bj8$	Q=#/96/-u7e`7N(Q$IxP@p]#b2@LnZ1$[plK{bDuEfBMt@/bBHy:6n XK}9RO;~; _Hf(E&vE%$dC54b$[4R+m[9h4`H8_oU:LC,&[=c(:a{vwTTj37OH3p\FI+yBn1$O:#wpB)5`"gs#A> #H-R4sR04|j$jpC=id62,ZFt7k!6B'gMAWB2#`=Xb.?pv/)Xpw1(4<77'OJ!m3jv9-n~!BXk	[p$\B|zguH=FK3.K0>k,rh691&LD?G7LL98V\KG"cIYcPzf4[381kc'[)!,ZS2dL!
_h;eQvoZ	_=huyjNAj,w3F|<rk}LB0)`z21d\Cgx5l^\7/0BFG!HfrhkE|"+QGn,TJP|VEN.wmvJN Xg'yXy]_Uf3<S/nZwW4'!}nl2'0E6$o(F#*4(G!BznZeij,c,9-Z!B99Z;n!HHTa9F3Vz0YWA|y;{(ic9qt D78mM:^_T?)!*#f1qM0SKf-+	ONT6&l(t6Z	mh}e?MH19&eymVI 42=	H_Vz?O#LNoNf9O@iYj2oPU-2gy-m
'	d:VTDx@`f}LXJi	ACD_C*>3:5=Xl&\O5"e=NNkEx\-G^|&MxfDcAF:gNqvB^q	yw|,.-lX(yo^S(?Q2[A~^Z}?h7uhu*nyEX"=Tgd1:4>/lc4Ij)Sw|=m:*NU`UU1I68#i[i#OnTm:*&wLAeF*|,C2{gOL&Bm,jS@#pZ*]?[drW	8YLO.\QSHj>
yWyhA"UPZ/mijNbuqa)cO4,Rk#X[)H]zqF3Lv?Qy:AU^.A[w^./ [8	
ppsa`z!"*vQOG0-S/H]{Te|e;xhxY6tR!c
G]\e<c1TM/due!)P{e}ksq0})0zX
1XppEZDI
5A*xS!BQ/Q=
hI{"~Io~N2 |i#_hhfYi}ff*AMm/.j<)^$G<M:x5>\C
sjdQy }qy(:'T/,bYzV%Qg8&!TQ546mm+v]hj4pRqp#f&z;Zq(wf#/Npd`rOEs:4%@"`3pU8/s	GS%J]bai}(0?G0Wyk8<Ux^d\+#?=bQ^aRjK,b%	
QUhu<=^m}uO_{~.d$xZ;TYDQ`Ma#d9law+UqNs@x3EJUoC\(7EPUJh]+(&K-1,<=nj`lqiqy_<
L-V:Im	(zu\D2>4F?+G P]o[_9z	YZ[kqW,"3}>F*:xC<IGX,:m!HT*v\yC]RoF<bHA0qj#qcH;Q],awbX"&|KA/6	8mVtUgHD{/v>+&9kg;phnBw(nh?B{%)h4|`aHjnVj7M-F/90\JiTl]Hfo'@Bcr{,t0"?=n.S2/y)sZOG7/)"d=H	t4L;1X"v3~EMm|%+m:Rf$s"9tPS_%xa ]NBubu&}p80DSsUFYe
RI[k[kINy
a${s::gI
9qa{y5z@^c9,.eUs~z103IF[kQJg~Tm+OFp`NbV*D54F2jN>`	W6q2A6^I`S)(&]b_{&M-[Trjg>A|aM_ZAK'HU/g6Wp	2S*9oo[$P3rL_s`)bVeu8&kS|vRx}$Kd'<wLaY"Mz6C_d5+9o#
}R)v'K^]VuGCDllrfI3Er
-%mW{kY&Lzv@Jt|;mG\sc8
Rf(1;eZ:v]C3]!#	7 8.Tl%!kz*w9aq"5ZP:2%oL{k&EbZ_jD=+DlC8}r`05n;k\B43R`3q]}rDiVt0bkpb6@sEX_?Lzw~N4AH@43!oiYy@8b5n%BBE6{^m8uYq!"UIZP0|!DXPGDihnR[-8#MK)&]u_5Q"Dp9"`06N?/R
r8c6LqUxJgQuJ~E>b* ?/,:h\7o}ieHW?7t	1SPWZOSa.H[Tt+(gWPj4Oi)duh'E
!^dJlb5bdg,=wN..c05sE}fLl88=X<GtuIw8kG?3h::n$e$s:L7CnmuXw:p){oJ(P4*vC(;!-q:Mj+@{W1sO6N<TxXSlh0'wJs[;Hb\wm.* >t_;+g#YsE$'p"9~*mag4FuEDe{2/];UWo0O1W.=vee?tv[v(m
j1:#S=}"OzX*dL+yR/O|-_GL>'XOct(BJ2Es?^@Vk5F+YG]b:-/b
]]dy(,yE>[3Ntc[JGn5j i48\J)Q-7aN?k,TL35A7!U|Ey;0-R~S$?PMA5YFyCs(J%Y4,JbqjGmEOVc>iN&(P,#]pa\?3beODggWmejzn]l<zq4]mn~e)s_"fC$J~$QU"LMh59MLCBCXNsir5m%u8L$x1~7_PU@zd)jb&{{' 34Ce]pc0UCp"A^Hme^N9rx,[yd+PYay|
GjMp`{	mX#9<s,6SOlo&e794'TuZDH;6=Gw U{ta%dQ:B'0c4/i(<g?n?|d}<;i>g_AbL[`t"\}y2_rZtu[tFE{bsn~.c_g'En]R5Jj]e6+7gK/y%W 2A45R(bU_UILrXgu\kT(i u) LI%ZhC*L!(_Ky)GDDy93i,,l.dF!P,,>)MCPT@4yG~YgZ@|h"9i,M$&/F)EO%C1aU\ I3U/g$UAz4w2]|(DgkLWmw=QP>~Lf>\Nc<1$lS/"L%"3p\04F4NE<PPGp}Y6^&AgR4T:k	sp{xC%f"VQilIb;fPltr)YaHk*\Ci+mDL/tYhciZYU<Q"}IH&A-LT$=MtC%&S@jXMrhM8_L'?G-62|t_bq"iVO$PhC*7M=1gxq]F;tV$$LIdZJ@j!`~KiQx4*Q#S>E]zTFGc'kCxCLp.I2Bc@g(#}3HmUD?A9+y5dR\VQ^
TuEj?t,F~}pR!EdSUC3yk!8vpk9T!T-t\^xL^F7H2C?JBe'iTD{&q_\k8WOlN|IgFZ8qOW!;5P>Fj"HgM(X'$mj1^1hEz;WWFEdy[x{W{V|;.OW7*XR-qKf$fa'P{a1[Fz$?G9X${N*%Q4/U,vx2U>S $&W@qLDk]hV*37LDD-oL