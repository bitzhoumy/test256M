mv~2gG&;n,jqk&pobk$!BrT5A-i3'8+I	:M	qsD=IXjL!Q)y7}D[<mWW+Ecao?O.(jz;LJ">vb6"S,O<)SP@Jq(D~dCm	0KIlZ:n^92Uq{C35" C-(ls4XHU!j6\rm.W`xxVO#+A?#&r'G/m4s7OUNU  ilsT)M3-d:1OXb/.y<^*J0JWAIR7A{0{xP("4*(^9V-}<K
~sAjMEJ:)c]r6zrAh|aokkL`E]wL+DIb15;fg(mt$d:xLTJGj9-p&gIIH|%x>cQj07\3J*4~+<YMglPMwx#
Pzx(~^*9mWA,LZk}sOht:60Y29R^M9w%Cl\odT'&;IKM\DQAd+NJ^oGI g A7!Sg	)da"jvk&QL{^!2ii`c`PJ`WV!PvxYk`mT2Ztam*+YPa1GadEk+Qu}6']>2|.g.:Mbp
wa8P>IBoNkU	4EPTz&^Hm9<w:fb&!#DjOAFOjtWw }kXGzCw+?fR}%PvH8Q=D+gzhN0(l;,vt81(I\U7TWw)+Vb-6c?RNoE$|
RQt!8+E"\xXsnJ>qN$*
|jRmZ$'C<U{m>=\jPYyER'K43Q%Q?lr6N(Y[`yAWh'oHrpQw<9vh^z*o,M91vTNQ&f6DX:ci~Cxad\&w_aBX{vh476x,i,ypi%%xQ~4j4w{X~v#wln)}NPStmcd.fhvxv
;drQo3(O(_S%VZs(E_!dI}C`Y|md^Ssz+q`!/H}U@	Pb3MVJvuOE{R9E)M\	SwT<,&-qOy=
@DKHF=Iic)dcnU88EYI_hN3X/'(7*.zktS\puoA9^BXc+k38XUmI@;ub'Q`^m);A:Q_5\.$s _GD|%) `w~Qqv&%uok8gG]B$8@C5y0Jzj%kyh"<	@KKW>W/!pX|?oe!-^a,zAM(.e'R4
:a\|KT;& v.
3t)RY#`Gv.gp-^$km4
of_"'u$G~X/-##EHUD+m~sw<Hc}w`^;ZGg|l]}rL<Kpu!<+m\gX^?.YtrL;7K/<1bm>|5~P[lezP4dYzJ$#DO0"^y
iE"PUQ0v$lB>@fknvPP(|6_v2[s3;#8;Cnuc~),Qc`#P(|Yyv},k@`.UBotssu+amnxshZWPa+(3+fr),"$xHqK%DRc=Tz:ais3#FeQMX02'SY@mI{/\2^aXBZM]F&7
GqLx.T_EeqcKjmx3C#4>1;_,M=SsAN|49 $x2ilm2P2OL[kMsC4@WmdFh&-{a,F[9Mn/J[ifU0/Q&N(B}
&j#st'l%E	WJ65e$C^q0A:KldFPN86!vKYk>!`r.q>loq^O2z*V\'P@]yt@Z{=pl8H,"Y]#oSl]O)\;K6[yKw]J&?g\2ee.AxQ$!r0=v$7]T$|>~PPGHZ6_l)L02O.Kq n#,d$uEdo^s_PifTeS[fg[M-y+2e<{otVZuXON*(qvlzU.L(0Q5sQhqEq%>}iDac1L,SS-(cqS\u}!w=M5rDRSJrm8140p;z]hh!KoY|F.yc}qL,R(P?$p*6]V<mX-/u8 KJR\wCDack5&"(fO]$)gw"JCu-1qMGtEO0dgF}.>itJDEq0}:HH2*4xuUr#F\EYFEks	[eFR$|FC%Na5"H6]$sbIOycDqt~-JcM^(U-|zh
~wMD?r_+3X	M,)]]3
FooD<cZ'~hI=}R/Z!0_%`kmmUrT3j$9OAd-2"*82{@G_Xg1y1[RE+s}cJq]K1Qi}JXYuJrnMiC?@kRH/}zo$cuLPeHI(]$)nQ#21'o1jb4A$X@VH]#(5U+o0*|^#0g$7XFfq"kp(=`.bi."!ILtfR$;}VAC^yoR<\~`eM9!#>geOeUXGldQM5sp6>e%hph*X|tU	O3?'!5Dt!DLwr=_7rlzX{lI>$)"bseA9plhP9.='gZ]Cf}n#1zJ,u)	8+-q%Q,c9[n-#KOV$JW|^Uo"}Gu^YJx9gEKl:d!SKMOa9
^Y-dC&bJk8Dtq;4i%j
JU9ww>Zdq_bq<&Gc^L#<=!uT	(T,I!ojX5o)--[*^j<z|XiJr",E.*gm
7yFs.p'+D%	[N]V:|
qU6%/%keFig&n6a[KB"W{o$s"Q(MTr5#!O"{4A3ZqOd[NCylN}9hG_#6i;$9)I\t}sbH>sH*-|~Q{P,F^q'`/XMpGf871@$UodVN,w\?=wdkJEUY	IT$
7rjxrje/>Fm1/I_l|kpA5d"pq=!^&eFw7O8&N@7	Av(pdr&?5[TCCQCB=&G3hzk<$	H	?Wj>?ECE[{1`4-UFey<n!YK sPX( mk</`Oad/"gK_Nzq:")BF4Ph,mvmU3kK%/xI*kr	<ju<f:($XBa6:/])g_Vs8D6]bHy+VFLy)AcJjC	*7]#TP~eM=q!@3kZvH1lx+C?&J9P(A"N6pf":W'fqyNs$b]1pr^ /<u{9#bOw9="
obC-lN@PUk/m.?nD/tT;),yn#z6)1fvDr=20_F^a>D'(&y`:1EvYQJ"lY0i^a}"]QI$.vOp-epSnBvU0G}"x8;+|:\RP0v#|3a<&q_aI_*-^oK66Yt=ceD?stt5af9P1^:|oiz80)jDw)
!
u8RsUOvo_fvTXb^#hM	"F48td7?	zGK;TYHB&BK'*W{DvSx$b1}<$J8U^w}YU<*NRGg_\weLQ}7$KGN9
%BM]6oPHZY"F5U@-
Dn^/|I[#CPg\j[A;vS.!TrB:GxL
0-jogGT>lh`yR0BNQ=w:Tk HrAyiNQN0:$${*gvz6i
L1BYi58|#	]t#U2VD5q(F|i'i*I
#Rr0kg)b9HpW(W6/$#~@8! x4!R)N	@_"T\ksh%f/-<s2jRpI"M+:VKk|bleKt0bIz<mFetbvo]EJ|=.U.+|9KGHf(1hb}qp[eH15^	2UNLaC"HF;Fd3#}k2Vc9/7ndJ^_m'@y^(Iu`ABt0gHd*J2C'&84:'!Ro.Trl+mk&SEZ?rd:jZHNy<kN<bEW}[E>X3u>F&31`u"/7`6 L|%t]PPLs+9FoQW6i{}WN>9'V,VH<iMjWu"fnF%/`q<\(gRI[qK/eNMKJ	hH_2tFge1E!6 A3lAj!;;Lzx}dRNd!\L33xqQ|ag/U"gZCrLLn>2AHJ[ILd.o/"9!PYq:*:-mJZnZMugt%rE1rUs0@z`<?#1k{>t?f;aS^-wdvlu9	1b>A5te@V38()2F/}05uew|CpSg:;g]jzP?N`UnbtrU\}%fhX([QbQitbG29n`A.*n	ja5&QZ1}e;01kQP-zk=EP'HBh(i9q1i`ny`kQ/wBv<BB}I-&1VZV!hs5h8biP'nB.BnfeWSdFX5[!FGAoX5sY5~;A)v'=#9jtL)kQ_/xe9j._lWvxJC^foUNW`I'gWls7G&^)CX1kWF]&CsCysPfB)Oq-n3p5@P:c:?Tl;?(L!r 7)JyZ5{7.NO	iKwC--7UAzr`"^4CFUMZTvOynp[Cy!qm6#0[W(eUG29+eC84e6]@Mi^3o V#T'}SM<DEo+	enzb~C\`',]p3mx
aG&4]_ju$EhEXda#Usv_Cep3xH~NRV.}zQx$yWi Hlx#k=M6:67l<8>7;S0N|dKScEQtS8VoH6N+_h0=<9&&31<cD53/)aO?+#0SdB8.@Hc=LB+ )Y[bj=`(]RK9lA4[L;d\Vb;<Aukpf^p.>N9*%s&xre:@Pw(\^/|5$Am.va[u%%2*0VFf/EQ_m,HI]zX^r]"Oc5Ef@_8@KFv
<*;6xdY$k3:}<).r^A\*"SfS>DS:K`uYiu-kT:*oG!+ZB0fw">$[4op3o^@FK%U=V{5_zu>.'\42q1lSH8AK5OB>AD	59:Kj|SY:ycQ`i	@x!VnS]W]ovL85zDK`Nyueb;z=H9C' T&\d+27wo]RLx!>j;Lj?XR7YlvAjs5rpyE3"tQ[crF6je@Al"'wfeJ`e	|2Jw	I>]s=Bk\6C)!eDn>Gj.u^ll4%wQIxti{Sz^+)\*G2w!&xi+tX/B5Q7:y#|J")SOG!V3cVX0<m(.$k1}2ZQh5l"0&"7.(p4.J0ts,;=J?]M)#.lCN]%+&iY`0!(MssMrsEgY}hzpE@B`{WFlS^&"8f+xo,N]uy?YW%)vTBb)^Hfww[F3b"!RZ9&	AqFO!n>4ryK12M;>cn+hbWCjUy">*!r,"DR4vX],qI7	9&n#[zRp[C>~n?~>Jk[~#\N1/}
yGe<r{*C6`Go.c&i/;A?bk&pBM`i6fQgGo^(UX2Ux[8]"Z$xc]Dd\CZW(9uX%-%K#FXK&79aqx=1hy9F)v3xef[-HDM.'f.CSG5~<s#?Oopr3MVm{w4Q1&?8^Db60p5ce_5Qluz;Z?m){{+`(rv
^(ZW&6:jQvQ;`)9}0KoY9pANc#v-$Pwaf8
S%jVEsc[1
h}tEip-0"x<PK ;yB<W,ds{nk_pN/&2OuYJWW$=b/;s %z{P#L)TJ'#f	'W8A`JKp3$#_`jatQTT(u^<sO3lGOpx;*AG"#}\DLR#963YLZU[?S,OI:!m2!+,Gc7 oCMWKC]@p1M-vs4z29/+L'*C	>iVYxS=jt-C0urer\
<5PdMB!W6_J#<OV^8pb :E~WB)|)2q[)Dg"iWG*	lxUCJ%Z}y0PkKAVRy2F=,IdH3mF4^?1&m-!Lew8qTDW2BO->V|`4\Tuz)_	o/o!4@E1pPu[942lF74\S&2i)U+l./q:+,<*EPvK?XZd~	]P
l(}?d,R	Ht9?	HHlq&`(JUi8;F)*d+Q;-?An}|9W--Z/_>3>gcT'cQW{F6m+S-4~{-UtAYi,.!,RA,I>e/^M-`?x~1
=lzhuos0Ck`8*]'.d X?5no?t$cA2h-zv%U_)Wxeu;2LlFq|@QU*u"P8a+=Scg[BG1M;6HwsRt#
l"3Wem_KRbs
@mRDFI]Q47R@.yAqyIl0%dKD,Z S:$%N%dtv$nMY?g
AUmxuN&Dhs@&`0au=p|TlF^]EfT6JH2vAi2P at:v[;eklLmn-)GT+%&IFCCZ833"]DW_Xj5+RxPPbh~M\rG!y^+;#
4Vw;aU6B%TN9)Hma[e{/na`pxX9dv}+FuW,J79Oc80i*WcB&13
\fFHV:ux..v`~d5q'EO"B&DD'Tsvf ,6l=S$[VF=r}Nk>}4v#Ld
4@LV	&,[\$4R3JuS41+Fr`aJ:3,eOgT<YmtK*6z7g'c[u7g	PjshQ|Jz4|=s>P*TgO:;d};C^Y 9O$7W5K2px5W4W
$=QX7Op[1Dr3/p/}87^9,$lA|FCy0alt.p)MCMo=e8H+q/<N-(B  gM7>J~RFMC]U$]ewBmDo!i}p	N?P
Ar5RrNA6D?o,,JtSK1|G| hR3=pxVZ+\Kh9ya'}n-
Ho/ ?u
x)t``\ [+~oN1C{ 6:?6	?YR~Im8O	5N-g43 fxI'fu$t~)y5]`4Ntq>Dj08x*L6<]Vvx!,,ls<t|p_=c2O4\CKha!My0.If+ZsmPT~velJpNiEV`cFO,m)ErHA1,h}]&mpdv&.GsS3sy;Dv_{k1Sg6H3*o5+%oMLmDxW+y{2a:.76q)yTITBnu(l'~PwI"dIg*'!^Vh'Nq'[Cm8$y2L,v#3b['6,5bdPa\](	G?`Zp$dt6yK_=B	ZAH'<B:B U^|gf6zkg|McAU3U0/`
@P>*\q@@|%$<)UK!TWR>1c`Z!.Nz#T=D<m<=PaSM
%N)38''Xm7 9|4B0Vu
xI@sqd{sbQHLCml\&rb%]Jn1lD<~dI9"|FuKJEUO&pzf
G_(Ig7;|H~|qzv85SBZm#q(!55vf,$@C%O^KA7;3~gy"obL"d`
cb8SbG N>]dESbzgN8gFgGc^iP/1	9!('WU5i=%E0DK]k!F}$>uH3-/=,?Z"Zr,U#'a*G`$0 ?qW2_I|14w#H}~RJf@]Sc""xQz'H*!|xv7x,Z;ezVd%Ky'YA7O~Yno9:a>n2$i+z|a<v6Y[=2\-5RgT BO$C[RG]	#'*f*&pQe$LO[=:KB<56{y&KOQtQe9c.lZA"N6e8s>2*!ntKWi|rOK3[>f'<	[+E$Y6Q9 Qrz_A\pV^aA/@$X;v%@d u;Q}^2`y vokcC
`_U/)>\IR.w0Znb:Q,=CI>=6U,;QT]z^J1D".s:D!yB7YR})]A]!F],_jF@Z"_!jpfFr[R,w''jvz@U
:i:6I(