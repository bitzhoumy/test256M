6/{M+r*M<uU5#)j2=Nq^3DVpHpR'P3`raa\}vc/:O<
WS0
"c^@R#uNM'Znt)0TI&|nc\*IC>s`Q$IN&Y82\ALgxL4~ZBe#,6|/,7n9,{
	<#	;\#R5
LZ\}I 8w4C
+4hs5d6BR/mUM7R
KAf
,Uk@m .uMx)#OJKoE=&g#opSCnBypd$B?ZgR_cnXsEl,rfc9VRI!{UM
vJ?$v}z;!MxwcWsimls|P2F*
HRK:,E"O,RW)q`%r~QM][y\3V!rh`-u?*D0/W{AA+W;S/D>H'ac!/uhjv><u>+ojyzyEup@ksH$*q0^\_QS	AK7TjyIU12"'b9$<u\F("t[.7g:F;TOG+mCf	\6el2t	5*`O+(xPKv?T\.
|g^nJ55@beS1ST&87_>&FH~ B#/X>7twvP@W'Z
fjEDf{MT4lB~)<m:2U2ZH(]nf=ma`x/13|!_1ntgD`DCg?f1~;J1)V4*cEp&1sxx{d%vg#DdO]^4gQo>I3_)]v?>'E1u6,7P<i}+FwqaYG~h
Qz,kSHKN~zDc5zR4m=q,/t`MIIb9~<-ZOD~YD86]A@iYBKU]	XAV#5]@Z(f6{"yB)hh:(VoZ$%3RTXTGNn(F&^BEn	( l8oa2C/5a~a@wfoh|?G*RH}+AQla&]mVh[c|K-6LMidvP^fvBeS@BR)TQ{rAb-;@X`Z|)guAB+=m3^B!bVM04Rf
]c`]4*rOoj>4G8=/O6FqQj$[{3@3@oq{qeFit):Or}5>lv}9G	<F~TX5HDUT#^ZI=\G6GrqKX3Z1HepO1OIcb8)IjP8.Sf)$?OaWfdIu7O_"!TgV1:lFG>S#lH/$`Xnb&
>.ncgfCx;(Y;fOe\>{aefjl!."8:&RTx0!f$%hco(_'.@|0];;\L9kLZPVYUKHb(f:@^n=R\-GBFml8Y4[#aH
S<2&8CFs-1oS8b
-]2Kb*r|KbLV)OLK6@Pc}<L$nO\w*rWGJ9nlBy$0LL.>1D%_RmUy6-u*Ut)tQ2.@Us/6v|HG"Z3He*"X3+/Y&TB=}2'c`,jC{)RA$qJ8{3\5!7i\RL&!--gL,t|(0j7(0EAj,R\\xUUqh<=|z=hcK/Gi?GT<NQ*4K$A+oPm<uYRVW5m.BE[_R]+Cj p5XzFDGGzMf]*<n\&:s	@%%j0CUqQKS9_y
TyjuM^oXr[%XM-a'%#3}h*$/Vc^2#l
e3".@p/FD`Vdm)/e3{4SQ~,
bK'M=uW3orV}#` 1wmR9HYo_dJdrswf04%5YshO{|<)V4L:9\(UW.f52|<[H
	3Ir2<ph0m?2hJkK,#S"tQZ+fW.g	s}o0goq .7SN^Pa[KY)pJT&B$wMY&p2\O@}lD>RLs&tjZltjg1C	=?yi<LT2HFid*Nz{Azxu{c'-jiRVA7e_t(EfV{ 	KBZm)km=e+:HG>[r-qN8^;KcC}$]fmC-1)a16^TEtwk'"G9BT61{;s+4.|.b8~9w)?%x$vN 7xa#A7)xJK~oyae*=F%xwm|>7`I^\a$teivi4De$`?EVDIt*Y^ k#-{4M
6yQAot]H1kQ
AqUvuT-jlK*<\X`J"@n2NCZpi*oJTVwWsQLv5pYC9xx	HoM &Yxljw|k^%EoHh5soP%%aF>Z/)%8WKM7zfz/F1%;yxkIt`=1jn+	/p6e,UtL(Ua.'u2k,da,-ig*`N2@\]'|+Ah/iu*2=rF`Wjn_k`3-6ff\AlGfhSKT2"c208wH35*o