Upu\5z/vwB_yM+Lu)MFB@8*wKC8}US|6UG_{+1v>,yO`nd)Zg;><--ME|vua.v}|D{A_Hvi2-[e}BP*+_es?D:7~J6:t>|w%)wjlcKXkH5~8>bIAOdYcu>}qUaG%E|u'fM!=D{w@@	tf8'KWq}Y+m@X8e]P6W(n&E}$I%=gDPgNe?k]\9z]Kxl;vR.VT~%]l ayKi 4{.v$US"n+81.9|'B4BA.(l#FA7Gu<0ht;.nbT2xiq2~q'*NG M:-;
Ua)\y,!O;}BCqWHb-nM*m??*3id%$
Jx]mO-S]w8e;Rov	v7tjcMkEyzDb\ja KB6h5~*9-T:Dl1OAr,w\A[/Z{~B=/:freA ?J#\Iut!*9]"q?
eMP8 g2XhDx]D
2wkf]?:U)@D<<&[!Caj]&Tp/P@ic>sh*jc2&r+AH?L 5aSSTki	&vQiR9ng+_/#d9
4\K6tz*zr>38(a.c@2yV>[0h&PZb`vXyM g\=nLB
GuYH_T}D .Vl937.Q 5A8@e_Le0w#iW=%c+	Y$sg`?'6K_Z)m|m[n
:cFeQ~3uUv~g!#p,IIoIC*Lz~\e-O'Q8,SFQKCSHc `=OUrg_vyr$:^m@"~,`6I5m
!Z?xD'o	%Bi/M0aW^_WL46Kj:ZB3,H-QN VYS}XJ.;7_Gpxz8zMsZ>)zctlDa*p&s{kj0w#"(#	l].KratqH>>{eRIXD]XxneX04HHRo,2Kk7%!9G8R4,pLs|RY$.w&zgZw|GEdL!F"n[uWn`O%>^&RFjFr`\R`ts~mHnY!LiCXeT?KeJw&~C.nbnb.v%,Ft@3Xl
B*\}&mQ`Mm74R4J
T~jv':[KDL@ ZBj>zj	`bN#OOU	~"]C7BZ~M[r2:YG,N9.PD_k>24/_?Hvl(b_Qr~\)d.Z"&)NNR0;o+-VjS3(/fT{{;ik*rx2V*[%v2eH6xa1W;nw-E[mo\[p\2]wB2~)r#{63t:a"$z#V"0Nv-4L!& i1ISIx	|P=.ud?q2k}Q_WtR;R"Ok	*c&ek$PI5g;Dg-`o\>5ZBeR+-N5-}iyBHR_Uugo'+OYX6h{y5oGf\K`CE/z{&smb^_s.b2LGqFmP	Sp-CEF`Vbc4"~aUmT\	S;V
,!F=4PIq3[|o?HK3I4=ZZq5y5,0hP&'+0HzQxTV0!|3Rdh8~
DD
kSZIz#j^{9=XeL^4Z?F;TKUL"U
52OYv~*oRDTzn\?@J!K?m@%z}uI^PKJa.,=5Du&7(Tv]Z6*X4&=bPTZOIB]A{sc8*T5ib\&mgN.>ITx/uF+*@7rqI;B}5D+dAUl#n@nVh5V!c5`wTcFtWes}:v?t~4ox))#X,8gp-9Ro,_T.dYH-z3EEY<\(O`Z/Q0jFq>P*>(z8aqqxW71`cD,NF!/(Wd-wGzeBC6^IN.,]8L3l5LG$ZM[sf.lXTdB-0Qi)\3J^F
FRk,Gg{(WwnV!B}fy!r-wOza4:e()MCvr-UQ|4Yf(Jwt&kcc|cEFj#/<v,=#LJ&=QJ$f$izTAX5*oMRk'yj_8iNYs/wU}=s}#m6rR`X3|k9M+Z*	8hTDzcqDGM5&;_[`P5L	d+ES;kB>#MNDe	]H{p%chM#3<n}>mFfrtCA0,AA5L5~3V4S$@
ncE> qWaLB515vo[7tw*uvhh	J$FF,ysnj$mMS :Oo#}YJ;`EnX<!3R{t[;T96qie[grBKu]}0BS<g"LGTnYR:`)D<A|"`.mGil_T!*?9Z-=V!4Ro`(FPj1su%RkQ<X`u.4=x\WT/H4EL(&/DtHM;vRE}o<j|0O.,?AWB{`z?&^=nUXv*k9t
1tJ8|&;`95$md+!r{gXUqgF>O$*[+V+47>NnJn^ieC2$nc"bX|
}F]Z-S,&S(F$M6&,CyV9'>4TUXo(zM}l'JcYKojYVSU!+c+,r6d}&m4n$<v`W?'!j0T.Xh-FBN<s2b{VR3'o^Sp#Tz*;&X1y"> 7u{R	[Cd<bLP$;ZLGVP{{$lW=e1h<8L\_a&XY7Z<lVVqN,w^Z4?_\qF^: yfr|vLESzxtM,pqKnX]qK;C*z+x3dXK;jX81}\4]Ds-9il]7k!]/$):E3#A}.Sn"Q%,:)tPtMGl6/;[H<[=Cj5:?Z;qWVqp;rS4Sm-p}AlNY2dMuWn5fjE9.73:`{Kbis0q/I,#.  M2AJ,#gYhJ&x087J8X/
0he.E>Yex&5Rv1xgOx*UI)qM,*MT7hv~#*4%!iM4\Yd0B(?,&=t-T+f0<|VL3Nd.2|9HYx8#m4Zb}9rZDFETwK@OrHD0FE3XwD3KE(d+kXAaQI[>"Vrd?KG]*7Zg*|B8 JgV[g4^Gdrg=\5ZI<opR[en38.03?3P-K=.WzL1v\%chcz@daM?KH6'P4yd+]7x	`@n`fnm4bT{j|q5B\2r.VO55YCN5p;&r}"fRo"
hkO[oD)|n	}O<4JE[HGpTU@qy.qL"i4{BZu Zr3y!e;tuV(^_j%MwPO8"vaL @+QK(DdY;i$^SDab]ue%7Rl^o,gG%itV|e,6GGj%E4XaVC[$m!cK+VU.&83PG+]u]q15/BnAj~-!Jxh}j&zcsbzZ>y7|beae@B/Hv.'1iuh:/nfhP+=fQ kSaqX['\5'"ea`x_wm><o6iQf
;A@p+1e&7T)bboBX4}3dso5I=ZhEG~FP$Mc6#T%`sH@2L/]9Y=Blj%BGl\y7{Jww)W/MsQ|=Qo52{n%"z<Cwd_a(|6_]d44:iKCC#uj,v&DL>flkJvBEb391\4duLl cm]hL&})C@e cDW-ZDNzl?dF2a1,,P&P%vd^R	U<BY+4&[N+>Pvv1'%
@j76^uA.~H\-7A/% :8G_Dwk.VcFh(<(	O[,Z$OUqKu	u%GG:_CzNb?ohHq>Z15?S<iJc-j=cc.pd(-w/,%IBEV2fI`_U%[y@g2B`$61>pn'M(&OQ#s6V,$4+qp6`/m[x_`3h&`+7\{J1zRH*Z`)1!nY+2C34UYV;@<ksu:+PM`3Tu\5Y)*B?>c*OF|Yt[U=Z]+at}k)Lc<U+0MD"c&kao11	o0->l76y^0Kkv4Y;wTW-mkF-_Nois''MgytZ,0I**Vu1 ,/"z6#su5+$amq	,wMa@l`m}!Vi,`L@N}b_T&H1[*kXc@G`:
='gLY%I&#L"
PI3tH,[rZ#
g/CHuKhxYm(|4ido6s`Mcc8Q4tlp=c<DOwn>:S3g&Tt
JrO[fc $YBKd\I4?\*-t8Vr=GDmVM#,'SbzIYDPg2Y	(blB5-|:[zxl<r.	0Mh:H>-U76):k}$?(ht!	8HCJ_H89?@?Oo$MA/GSln v.5{}-OPCR))"1KBoi69CSD<F!Y|S\\4`.ZY3du9n;Kq4HK#es/)"@F;*k;%IysYzr#jz!I\5C8Y!"TJN<7#u[@dZ]XyHD&%b=9wQr[lQ :Gi^`cEYn/Tp
$1|yNI&QP04U/}XFot&:Tm@Ar	{QuN*(iTe#sX-L5A13rnpUrBKQ*DZ(J\V@R icv4Yyohw5KJ(EM"9(yOr"+(Tr6d/#2m\J8A,A$']En
qz|Dyq)M>,>7
%[@+cpQg15sdwO{@h|*oz<8wE0h hF'Y`aSV+}yP4G7cEyD2+K7B}Yp;MVXw7QSCamn2]H0y;9{5a[#3{h4QE>Q,h<#r<Rx~TH(z9{WHOje9Q.R]q}9tZ"ERY0xro3G)14x[^OHMkzuR0GqX}`-*zh/qd[,(<rR7aOGr39`e`?9Som95!FpY@s_Q}GH:gDIna:#OAH{qTQi!8F;fiyie9T-lO9vMUF$""D-]03Z B{W~xA\'f"X8;t73AjO;0+70%[RM;dRRPO~/8.IWh$3nuatlz0P&	NI]b+rh8Ngrxhrcg2N0KY!\y&L-0V_=G"/,=p:fuvAa)q-|bM5,v^$E`!F0W:O|]ur%#1J ?|=E/;y&e164Kqqv5+KwtLYz10\oz!Q/XQ wh2_|xU'|i'*Yp\J1LQ.uH(lacw{CEj"}oPvq?'w2T\"][oyPyc=h#rNoYsY4/XHf_O0*q<32M$SniY<-Z6Ehwa&4ij%OR>;L'<He6i.CqNJeu&8Bv]yW`|}M|(H/ag5MURsUpFUDeRC%QIj#kv|H(6D	+Z%:Zm[(.UT3&M_5++v(rT?AB5$fp-7(0*MB$1A^B2/x!s]!WbmwozMSW2[>]_CeGlcujU9_eU8,`Qw@~}4;?lNHP*j\e,;1vg"@lu;jqxhNmYtF8n 4.k.93=v2R1$U>I@9(x*U&0cdT'2yHqC7U$ipEh]c(tR7;T4]lR*1<^mSi*F)yB*O*eUiy5znY\gwQ4c7HkNO3#d;W!u3)lr\L}k{-vekO1A5L%(7kMQB!qsp'I6Z5cR:9^cdR8h}JD7)JZV4{E?v%ap8B+1vu=Yl2N2a|3
Kr/#Ja	p[7rx$Vi INuM&A8ej+Ox&GrYz|'Z_cY w9!CrDxB<%jkJ3nQ@8*(e'MF Ytl]R]R_zxB]-P3trU7|eDE<RC["57<>@yb`(A9t!GQYsv\|7.J9J#6+eB*^iu7SOR)L9gNDXB7\N:Df'M4`OS1HwpH]]f&
|iddM@zAT3-#R!tv5s;9mW|Z9Q%po	a\c7BdGx16g|PBhmI trVANri!-a%Uw2R#{A:,~<J\~otWCaFw?|/Br6${nzvnB _UbAwS<TR:D7-sjJlvPjSgo_D2-|
u+g~cC*<2_YlQ*#T}uhJV=0r0"xw7;9+B7rA-$!Ql/EtAj%HXN<5>>=[1"0sEkr6435~76@(@N'B(8|0RzrYpO,L]g6:RD^S9XG#ew<y<7a,]V<JI<9w6h
SCwqK4IB[^H7'*{DGEQi7)Z<cfy{EIFD/h@w$]0<|fGK	Z)m4!hPih4$f]6KnN	]~Hh!3:V?Ys:8V8MI_-!K{w;(>	7o9=,66	:7*"|I1{?xJNgx5U5s]~ZqS-r|X|pfz%s=@rKAexRbsT<Ymue@vy]EgN.cpKV\Sx`O%!x+]@v#)6pyWfSe6xd9'Z87|#xD]DMxr\=Ux=ik+I'120<=fdh)zAl{3eF23<P77NnI?(E}[=S;Qeb6K.&_/m!9T'N3-besxC9	6'8Z1:?e;lJPGW''^v$M9;7$3bg`BY/vW[#P!y}K)+|*F?t.t:FHJlG!:^1}5{[N"\*7)S\IhePlXx9HRsw[ZnU25f=!NR@@+p<<T)X#FVvWT2olX!6	S|	$y(n~T)o]	qCIa{{uy&:TMTJn;[r5YaXmU@D\6=@O
nM*yw*?$n<*NgkMWNG&^>7/ VFy3Frq.El;u42d3FX16kiRbO5D+{_M}gZjre#{flxJj@H8}{ <N%3 3$~:e<yRy,RD	}/0hOICE_+Mut>qi|K"5L	7z
sZjYZ?W5V:~\ImG9pf/Y5vTknrtc$`I_t06+Epn">rbude34$( VI]~
j;r9]}(({X87p}0$<zS9 fYr.({-!NvHez(mfjIkBLFAG<\lPIT/9 a(;j=xx8o
J[%]k[o[b]QC5;WWOAa wJ,$ed(Cc~lw:X4~ghQhrIAktU5u4Dp]ux?u8,Fg;5j,2+aoXsO=)W<w<moP7\v?UK<HYfErd_bb--I=Jg%!QXcyo>.T#R/~o;'\HgB[ZaHxXnUyS_O5._9nO`dHu>p0DwC%4	 r159c(>r\KVy9&e3v?UVBWmctwB*xFYF\/l_D	qJ/:2:R-k:Nks9&gLd!dECaD.cq>%M#=^Iaz_+tJ;Y>@vjS[9y5dVlcCvFejp 	K(Wo`c3Lp7UwE~!e2o[,'|LUx}eFlX-R&qIUi2t@Ne`L20[c4s(vqNP8{:9_86g!N	`KA#-,LS?J7AV5s j-=~#6(S}'EO+"y+CRa\cHC~\|3C#][89w0~=B&dHVbPd5#)c\#
ye40QLqk?0Rxj3DZ|:29]{'QQfe_[kmAjX3)_IBTSqxUd_M
^fzOqO/oNel+ahHO7.xF$ 9~uM[#bW143$P#w,]@++=X<B.S<:	R=\?s@N"vp#T2eQ:YMN*Si{DzEE7n~j|NH,yu`A9irt$Zna`=J#7dG]:IO2\d_v<d$:Qh<]i\	W3MPVH?yo9feI+4Ez[nF	*X+5xc<Aqx3?5
exX[qVMS"0dVB,g[To%q2SUC7y[{G{BTO<PGsV>1/lle,pnS9FkNik AfeFXs)|ICT|PUOY:zAY'ph8~C:ZZtWPUEG<+B!?{6?7DlOx&?zQT
y :qkDyCpPomR<gC0&+NP$sqP%[nR5oa6{|V)"
n
^SC+HT>e~_|ca/-%:t;\O,)jia0wv<fi
)7*P87-;a8P|^lPxw_})t?rKRy4Qq7u+yE
Qn&"
1_dwLj
^IH	$CSYlMB!619%h&WD<sRT)`v4DXybD6JTk
,Khx,l2Z9c6WM9;v
Cw#KHQk>;o;HkR^d86>WA2FUlh*1a*3\n'X%wt+pbwEv-WczUKVEbQAba2a^7MB-K?[wJu/$"61Hp'&:tW(7]8lC'Y \9hp3f>.Ai`4'B8R3'N:(^8${Z)k8WL<+R$or!8RFt8I`19b7Dwl_k([d!,L}S&kr6lsE];2bN%$(tN} s.mB;L^F}vNYlgT^C<OoNGFI!"qPtJPQ<1 dg!s!V/tboc?&?2=Ssg`yKs4i1ym.t\8*buep2~fX+Cjd*(woydidpl9,epF	Q=	;VDH|QCfI+oq.!P"FA5	^x1K|-`f@xe{MaaO;W\]suwO#%(:F~$`sHqMV"ColBrNKIZ#X82:X'@Z@T"s
s@$Q!)|bi=gEty<Q3efm*_~xb1ol7EH,gm{.SmTN<N[oO,_md68r/w6'wj3n`}C:M*_f{Q-|E_
+rggiRcO
,	=NKgFF2o$'VO[:-=r;!i9320>n#_iCUc;3ssVPNUeq6f)bCb+KEb #1;cG+O&rvJP^dfJs&-:>?Mz-"|$~2Ob>XRDcdA,-bDG$zBWend5m_LF8o6fnN/W1w[T,36B+s!{c}c;)"\z5F#IbT"berSVPyVc({Tsig2]|+5WGb"qPDqL&eLd j
AmC\nxVe(h.3[Yw>izlksTo0K=`~d=b>6cjB}J{,	~b[[@bM*eHRvOi,W)t?[1jH$;xvxcs>T]4:fR_Eu$%Z[.8>rV {{==p"ccI{>as&|a*i|#,HC$AN7l[{X0!+V>#};P#m7d,qLl^RMQ#Q>4]uCs0p)<rJpj.:L^S|{6q~Rn{iH0[D-kN.e	hAPv/Cmn=0xRr6B$hFKGm1Y"m"*1=e@12i*LZ(j`A?}7us r,Sm2;0M`bW`P;]BQ9Aa'Rco$@,U&or;~6U8iWts,}Q#>e\KR1VEphw6P`93!|!H>6Wab9>R|DZS0~^FBF{<l\\V]y5rhh{Dw?[6>Nav>+lZ[z1T1!C2n`Wa
35JY5Xm-_=DqE\[@]VEMk#T=|f$6T{!9v?a'yL{tiXs>HRI@st>aUdQ6Z6CcLoTST!$xX=v4DB@6g,_C+~&(h[b9RM/IIfhBu3e.	bdo,o\lcR" c4xjr("n<h$hZ[e]%*^(d2x}+Bfj`X=y#.ABIOO!O*7jr3i9B8CXS-8v)bN6Tj)>9.Pw+~Yic$
rdcpz.*vmqac%/.$|/xSbs}d)"ZPn`<'hl1yks)PK$3Tv&`H!l+MI#?q%2-v^T 9D"H%l{GJwGLyP`= I7B7\,6?3J]vG9q5uK]$E4
8iag4?x'~.m:&N	'4'ns^-?J4/$4o4ClnD 8PHmN(rOe'D@!)[r^8Mf"9)@KXV(51\sLb-<[Px
0u/5YJR\MyZ6|]aY"@IuG-#[o6}d{5=8=lyu.N19'XoZ@Zb`
AB5:4K|M
+_5zNjvZ#(fO OIUXe[jm8JG)U)C;n>@;s=&H	}rE>F,r1)Di)WmFV\R9_=S<y?7?l19;lFG[4>At2Yleb.^c	}cU97zA4c`GB*-mC/p+|,G~I3_zHJlIV]CB{:a\[M3w!`hr	I9_FUTX:oI=C;q#tfE,02na-n;tVW;0/"$G:#}l~H [y;n\bg[eB?{g1z^C1er'%HA9`IuE68=JhEK2x$mU1Ho$`Q|w4THdz-GM"B>U'#k5`whT6@=1Wr(kn_7#dLwIj6Kp)BIeAE)FGw|O(AT0Z>2IRA}NrMNPq{\&	hkj"JsKOd7#EhvMx&trfm9
|8aT5Jjgu|RCTVZ9C}i,qaFm)!0"]"]8;f6oBwPFzjjT={2q{lVPW-yYv&{*C\;r5yl[Z]HW|q3.!~>xx11MzfpZyj$Yq3oF0Iee`aa})&R,#OoM.m->]scKPa>NAx`v<187oV2D	K%w'9i~^U+S|9i="Q4(	#,+w-'$DsD?xigIK^@	?/a!oh!nV'7nQ?42EX^G%54v~[^q	C$&dyO7oO_U5UbKxm_|z/={)r9;&cxTVHOIR*YaYn%^TabpPm^ndBD&.;mV-F;	#2=S
wTTK?$1I}30$V,[}/}(.T'S>Y{C!YT+5:OZpLi]pWZP~269uPzWBg,-4jR%je}6Tgh>g3aRgsVrz=fP(y3(9%vsI)G6S=3XD'$1N*5ps"^b5@#TJgdb4W<p2f oKqG7V.2jGN08^-)gdmv-3e,+UOV*`Q_>B7gN("g#@=B(n/TI`nZ	tL[YPOdN!-fj`6gIb(3Z3YnVc.CBt7p6Rxg:<vK&`QW\5d33Hrv/
&t
Z00T=%vD5i5<21{*H0j#,8cc" )m!T7.#:L6UGCSj=jg[w@H4JA'<^2D(VUM6hLmJQU&-cZN6B+,[\vQf*L!t_O,m
&e!M=RN$J=(q\L5s?$,AM!]<9ugi`z7AGK:ik.QD*#bNiJEtv~7!aVJk(~tJA;#TbOeRmw@(M@r]DHpg?R/a'T+T\Z(lB}Cg^jo@qL!ZZ
5|o*R}+c_:*
DnIX>
Nc4H-GtozH9{vwuZ\U.9rjiLg!euj;P#z
]ek|[Bs(\`nHeP6czX#0HL
i}Oi5H}9VU;u`.,h?u5_;:dw$\}e""~cbB[a0oXU^kA+P'!}Nv`53L7Ze|<3	H\,\G"i&SK34*u\px?7	vw'*R:Tz.:a$bF?`!&`l}U*:ELMb*n)_S5T#'ZDvDiG+M9!_=YLlhGR1KQW,-uM"BCb95>aw;PnNSN,GV(/z|&=bG/wa`Fze8J
];9?<a=	>626Mt5K|^FpSH4PV^.mcr oJ=RB
+SawaZ1hQ,f@"hEK]a$q41Bv5%05ih>f"
F@6#Ras,%}Bw{Z'En<%~s?*Ol0qseiPo@ZDn7_QgW3Yn3S\0ZfTJJZ+)*wX`wxD`94]o,ieqdq8&q9!LfHYaUM&Y26_.CIjM>;2Ho2$QCEYM_fH.@={$5f_M.j@`Oa:sG4&_g6i-Q1sa^C?xX{<(so%x_1"tqF	a8DqlE,MZ9cx,3QSD;+SNe|MbEn?/#0P(UH\af#'&QnZ;C]CNxIF@S_rUSfn5nH+7f!04ia1v]Ogcm{V?pnb$Is/tR=[I\m-A\b0I;,88[W*I2+f?!;aFa_TiP!A;_hab+a|N+~+qM@n_y\|~)}$$po:Oc~z1_&$Ka9v~?,)8G[v/Yq:{O%8&>\u/B*`Z tbw#-dUZ?@NPDbqUk!iQt9+,F8~r)dz&+}7@))f#YMie.F?AL{Mc(;qTwp$\{F"|T4[(2(<5J?gd5x
SAIUzx74yX7$^K;;AMPurH%\w(f|D#X\P/}BF"aE
!M@C3AmC KS-E6KtL8;g/Op&&!P8U$XA_Pvm[8|S.Vr>~!:qJC>A&KR"rDG-Bk?7oBd5o"G&-l8nJ^c=JN`R"VdML6T(R~ GGI[	ARL"0i`6:q5o$w*$"Ds\:h`TLN"2Z|p[iHl>i&d1?|.4UtY%.rZsE2n,EuIK%1)0S0t+FI{F&5%mmqf	lB<E4eW9IJ`2Cs-mIoSxd=pg5TWnAY8!!hKq?%!`z' kr!k~s%WoX]tn?H2Q/q@rATuLNswA_Ei
/O
!k;v|rjEV(de'	GlFv,b%jfoOS_ly{-	f~/?H&"`t`ajNz\e^A_YLsi{p#642LN?JYB7omf(+kzX:5U\_,nvtm8Z}D'n2QBXiGF!?Gl)3<Knx?c0P A7,gr#<I5'!/taB
IQ4E__fJjl# \1:no*@<%m/A<42"czq~^\AIt[.iG(EdEY,&UA?C-(^a)"UDV*mluHGw-IH-l"7!'e@%*XF#}=YGn82APkQ=*GQzWW@BQ<6G/ ]V9\"Nhe
{VB8JRQvCv[;v(kThz~knA 38Vv"W:u5t9>YP8+T[m~JGwL%Id!5yuh`OG5'@}!1Aiuo|yd7`&k% z,P
Qzn	{Q8!7BfEpTGS|w2o`V5)2,iu`(+cN-A6MKEJR,Os?k3-rM3JefKR	/x/YI2'+?Ofh2fV|MVBwJRIcz|J
i(<ZU$25P/3G$
4zYB.A"'LfdfmYqnP`Wh^Fp`]Cgrb{ )1Q.*Wpc{XR0(Hy%hGe'{=rr#ntx~G>*fUDS<ALM RR#,ihv^3}4T5dusjpt
2g*`lK$)eC:*nB#7c}{?!cuI	pN^J%R[iFNlkF>w-9vRn64zITY\cy:{g	r'[i:VD!`(/a[d6}$4cH2|ooq0'bfGtYo}=Eg4?VS"%u%+q@\@1;Zxs;Kmu'B
1bf"Kkr:wwGKY.Fq%QM %6!7JgZg>N+RdC2p-#.a,b0(G\_\DgS7n-:GgPq<aF\m?\+tyXBq)#tf{0o*k.K^i+* -`Y`w
cJBn!2&n(hd&0$fNsRipU}eMQr@K\uS/Pr|iH)O,[mIT|&y#yg582=n/z0Ar	GHk.-(4(H`-<x/5;2q
psg$poo}N7BGVgw!c