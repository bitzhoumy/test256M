zp9^B, ,<!4=P&peW;^<E<GY/j^0GOOX~zhrX6Jr\}Sk{p*&R]g)Sw9MI9Acb9au={y_%|/Mm1M#9,P4^&[rcr;@4>Rylx75t6&]}oI@j:u`S8:#9A^~=3^i
=jyc{Z+iJ:'j%Q#h#\(>Uy_.y8'b7|)LJQLa6bbQJOiR`1di3?:PQD1@V!d^C6]J9sNp5#X/g)zXfRH4,+
{j+u2".3<^M9jp]}B?ganAwC1swk*f5xVf\H	IP2&5~hdo6(mRa_&!f,M-;dc4]TeQ
&b]0z}Sb0xAxkB$hJlcNtj=A)&7L!*RF5EH7K2;vE	uS=1|b+.zhl;;}DPG3sHFp1,gSt$wI.$-D9":jojRxZPuS,EA$=x,0p1y4m_6)"TFGRYak$K]wp#LA-Q$!j"fiC;\8ac/h6H>Y;:&,Vco>%MA!g:y9X!^>(zB'|:ZMzwI{	,kV3A];V#GHk~A!l:4	9' j=n5<[}y(oV:|B*7l5G+!B4h	Ud2|l6e8_x"[J9V$jn54Q]Oq:"cf~irhJ' ~:Jz=|zj	ue)U^xUj&N0r3I5ymYRTioD2*>"Ux<gs=:TdJ1/OM99.$R4Awn-Mwr+0EF,p
WdDo,eM$h{\:q\fj1<l0W$KND?,+,iYGR&_?+z?hJ821g2G->`bl
2)=buKV=;Sw?r5!	7p_*+Bhlm4N!>T90\ulywIxFs5_fAR8^`Cw6o6CH1!$zgm/"E=Ce+,nuFx?mUE[!.4:_-E044xx/D3g$i?Z}XUX5Z
s+5!";0!#b&&
E lTQxz1u$/Cq[b~l(7)TSv_?G97*T]=u&bM6+PUKw3c?"}k
 UC+i^#AGY rl{OXI	_W)%Y)|pp<="OZYtQ-)TvB1+jUzD5Usq:FE[%J8Sx!f`PS}C>&{h}hE\+9z^F#H+:RE`\$.%j^"/M/FT.<HKe.k[7y{2m;KxjyR>0%W8=XYNBO(V]kUa2s	K510Uz1:nNp84_GF(8!Ritq,d1Z~vQ,*kBBfm!~33 7+y)MG]~{G@ZHeh7=>/5^M`+F}nU0f.jE+5Z&,:BkC\SzOzpX8Wk0]+v9qvSV)"yHPXad(D|	w+1jIjb-)LR6fR]n2,eW,g{g)Dx'Cz-JrE]:]"fgH	9.3m]%a4m'L/"+`N
|OFB^aB#s{%x>QO|B9anoKd_n,S2@6\YUK/89pQ9y,^'V$EUF0Kf|U.^Eq94i?[*%9_$,Q6u*SlM(s%6B90sA<[AlWCl,	'p":p1szD7
EapHl;MT-DlBN:6,+L&S.X2H_69&qbz5~q]?I?Y7@m
{}K@._xl;SI"zDO^L^B ?^j7>v-C';D6gdW`/kW9z|Av
vP7<rZkAz}2OQs-c4P
MIP2rO2-uxz1-FrlqVOwlL4HI^%j``YJFmOzdtz0.#
[X-SvY
=gF%hLpo"?;?p'OgH/"Q1Wx%LjG^A$$o<:mlX)0#y@:=UdAs9s!nAMgYcv^F&TWz7cnsF=QzJw&|u&>j;gb==8m3Z!wEL?1xZ6M U_2M$W4 h]:MvDY)wWCWa_H=8x;M<*`bHGdQ~J(RN(SsoxqG)Y	dw*ti I^)Z.ey	Ge89BR	c*8$@?0 8N 6j:p_i|CDXR=rI:(sMncWA-=lC$g/ck	fJ<tO>?!ts=_sD[YtuK?Id7uAw3!L+Sft4g1kG8:/Y'1VJJj/cD^YjJmo\3[iee\S#GBt7+'/)IL4+\dGOS@atYC!wW0=6`Rv.G4	?!uW~0"`w<{j~hWak	$kV\,!@5J{hE16G,GGU$R,]]C9 )Mmk])3ivIDWCSo'qWA.uGo]RHU 0GK53FU@*na`gjUpVeyihUWbapXM:PDZy)C7EzyWp@-Y.o."emtMf;r%SSnP)cqnsP#)I>y}Wj<r&iXf}lIO=aD.sf xuh)^%4&g`O|O:	l$UZJ=Mm'y4dm720'rL"-6D@,!Di\5e<O}7ZsQ4~C&4#(~QJC(3C\\,3}P*nl+Ty6w':<2V?D#1Qx[bz	ElB6{<8dS"4p5v^vwVz46c.yrnZI8=8Jxbhrg%:E?eySHWu>cmrg`9u4)/t8]KJrPZTrPqw2!*o0R4F s@bJxBPY-]r)E}-k'6W"yV[Zhj1N<q*PUkv}"^'8[T'K'4[z 3HNopmaSO> bVO
!NhB-Kw>a@'P^wxEQov6y-]Jxo_x"-%h?il[1YnG/X$1}crL 
9#&1E>ANg *6(KBms.1UhL#u{(56b6"TK&e`b)E=[P;K]'E{#dt>7{0j|s|6^vg1{Y}1a*Smo:su-[6_t"OZ`\TF-#/#&YatDk ~\Z9b,^Qq
eQ4^G[(X;;*Bi[cm>9oP0z1::$N7$M[ss-gC#]pj5XWU%?!FaK~i<3szF$&~<A{h^/t8(>i_Tzw|-Y,GY[)s^{>}9yZ&Ox)%blCci2IcDH4UY?L{'&'Yo1fzVxn0
~`A#R<IX-A)oa4uh]MqLjep,	^d/;gbMk5mk;Rn3+c@tFE)m5'kz,a[3v'[mPh\k^'Y\iKw)=|);_W<{}vsuiC@4msvr7,bDAn.sbaf<=<tl\bbwH'"S0(I0&?I
@XYG NW#*K`rX+SZa{GK2.4`vfc7[i:aEl(,pXBfUgXeI-bXDgJs9j6)>+5@G7zm!z20#aS3h3r?g][l(H@$|'KkbI?Xk6HMy5eg}N1Bb.%txiD~>]l>J,jV40FNuN#D6A,-W.H6wTeZ@*xE})GI]s:l2CCR>Xh?Ro/G4?2:JT}
)h@EIiW&qt5qeBx}"Z7a*4g] e4A|iyX2!,=*X0Ee4sCR*!&O<r2hYZJDB=~;x}`\@N-XL(x1%k_+S~|IJcW<,%F:L?qw:pjLj3JKG`+nB{dzbpgwF:'d_O]MYbf}i5>+^6$Q}lv0up|wm0zJ23dX"9{3b1\YXOT_o R6@,Bd	fp3.R9^{D~0FnKz\sJP.M7h sG7FW?W!mQ"HA3*9C'</NZu"Kz!w_|Lo*x%2<L?*	W`kR4E\8g<,//QG1?Qz0/AhA36YJW?A7S"|@fcPl-loCHGT1*$}a>j`btF;D1|:P1&{5,nf~.~q!CMI?HC717DY| HUP0w7"Kx|/'(z|uSR%htHTm9AnlIn=,O7w"s8]o/OzFX]Zw(C}%5hgG9{(d)yo6
.(7gue:5p?D}~%sZhJ!DLAV,<y_*YqN{sZ[$Us}6Qz&^\a-O.kG)gwptfwx&Wvj|`FZ2l
^XR]_9=!*[=A5\dX(e;0hhhWg"di#cONhpm4sV4KN%,m>07s~6`$.-/;2'Nb]XpC@zp&EIR[|;]fz=~-jSdDaF1=)*fU["rt&8e_ 
>z,H'0L#qI`HNFuCi`)#Z
y!M"%GM\%!EG-Qb!/%Q.Pv\VW&h|8-H\.Yw!,uCc7n=IxUu>	0&H3,_n }7Zm:6&rmhLwZf>1oBbD${|nwcpDO8Ag-AWo7KVl'9inWQDY) 4p y<EjgpejY\[wAta`5JYM	OT>-3U(C^v:EalE5/moZ[^H6r
}k^1LJ-fK1Wku#b9/OP<5Hgtk_N_/kNVYl~k=lgj.5-=;0"Aamo8@Ax'zX_v:t4)43 _<Gt&yi'A)v3anChx},&s4tC~.mVrw:u&hI?=r|;PM6yT[|UFwRY"$ 	T?eb	iYN[&mi{	]|jp=	{;$2*nVt_p6bJx>`z"GZ
-yQ6$$@Sc!u9
Pyl0v.5mk7+(5xz&FkxU`7RO@u=Q[YnCA,u]e/E]a`sM>Lp}gCzVTh%|Yq*&HU%}Io6w(FI4EP4.bc;VO)l[*'hmVsK|"bJAJZ? v*VbOY]t)	@J"Rw%zKf,>2DiC*L@SnFvQfz{GEkNI~=K]ATQX8$Vw_dossfJ'$GW!1r%bbU	^9a5i9	^:rR#d6Zt=$i>x|RMU3W>(d%"\<5ga+2*.oqov"uKl,u @&j,r.Q}ZJ>OR3ivJ/-N;Fs/~~HR5CYr!h=@1u&=)Ha(ZE:k$H^POBwwX.0Np:*haN?G{8)=tVj3Yiy,$|a=*w0"tH:3YK\efdJJM$|kO6gDV'8TY1_)\_._Jyb	[b_DzK"B\6=ez&+hXrE@{`0-^*&yG*3BX0`fDPR*?}OI.=n=)`P1;C!M,)1'C:T:s AH$sL=pD'pYd?;-v!!U #[U9b%r)zJP{|adM.as v#U>*.0md1q"U)oW$xL*@pg8cn{xu5ac_n!]2:CH&8O=W6n$_I9Xnu;fe
CJ=woIrsJ[c^>5pgxQ3gWnKcA~PO?*'snJ6)dbsF?2rI2 Y|U@Wsny3Bz;HHc=}G8)<kT?m$o>e56T2la-u~"{bU/Fs)"WwIp|73&W"vsMfEPGI-:Ksz&
x&2qBEBhwP
%!Lr&sqW^*4>&`zgKIxqVHcLU+}QsC'Y;s!.)V$<^hcW2V
N/c%[^j($hY!fw[:sd!`Zf`?d	2
M&)4cnS
&9'Xx#O@U&x`a3[CG"Vtkusu23	d:]IOwd r :DX	CH"Bng|;jxKNVKS^s/ph)-ONddjMM)PD^8@y(?=)Za9}c!z@Mv7I$MJ3*-w!*maAt$=~'kiD.vA{uy-u3N"m`ge{)j165gK2'QeL|K8*[x~< 3*0HX\)o2$!3}J{e
' C#%
!6pg3jtl;WJL01i-W2}zhEU||rY.[[<k-!fSx6a/.}V~$vb9\"^"'PS^JJ9>5"LSQcqlMFGnzJEb9WU"T:fh;n+u!pg^DBwDBh"x'B,:Tmw?htC);0uZk"}7@qf1Faj{W@A*x(+<|d%8;C6{+Db<,&l=`m4EXihOq{@90L~,BN7CXc}TbN1PzSp|]suu5E:>1Q%:nDj7yJ<1gv7}{5;P;b5$e)M=?ssvnf_B8}zve::ci"n4%!&,>Kf2m$aV03[D%8qvnN"Oc67-FJ_CmR|3Q5L(6Esd\)z*RZ)6WK0xgHcf72:9s,(9saT^a#.3*f9jv*2qW%*
f7B%AN
jwpe;f*"{zCvJabp_498O&zq
.S7X7WuKj]1a
rwE-t,?R/*.8MH%(GEd`}?8Imv=dr ==g90u{:1>=(ho[B&sQh	;8
L]w=+a5fz[o?g~]wE{IzQgkG&&{||Lq[M%9YjvV&3OR^8x r;'!a.r2:0x>mTHX>FBYEK9";k@6nFJJhqrEF$y>[:Pf2aQS
qb &Es*pVe}@QW+SQBAmLIx,20@#3!C#-.Z8=,5(kwDMbYfXy,$"`>#Cg6]e^"S[U.5KzW\1&A\z&7Cq&ycL;pi%	>#X@#\ =J'%.=%e=ma7Gv&u>2	`JKW^SbOS})'f,TH/F2NXiDwMIfoBvzf.""H+zQF#DznKv3JU|'rizc5R)k^tQC=ZQGQ1Xy,%-jx>/xXGB)(0>YKp16^b0c93m}YC>[3}{v$ov{"l[[nvr6/uE]4o{PRc(@3I/Moa>N	Jz(8qm+EIZ4"=g0scv N{RDoQR"HlVezv	']OhHR$]|z_BEg(LaeOklu@KGiN'Om>3Wp5S\cB&n/L"k%r%HX7-R89>^f'IX*t|>W%;D;z8[qS`D2i}Z43,Z$Z*w%$;O}O0K:`7)7B-BTr":&P?{:I.h5=
xQh'}\}b^Qu&sbc+dZG/6\i7>__DY/lFl|VvGoEjsU^:f.Sb!rlae,6O*GF?i,}4^b[cn`q%/.(GN.\2QDI%y\L4ynv.1hR};HO]b&bW[wL,Ik-EZ+u[ZVH	&%i8]Qz4pl6:%jLSww>7NYIChJf<`rTm5 oV!j!m/wo&~D/0Ic}db3X979Q:1|#C(Po#4LWeX-)(cK#u(f	2tBT:k?WhC7gb%E0=9[~GT|9=\h4/a6ik>{W
&C'5bSfTke3v"DpFU7uc""cp0'$Jq]OvGW28'/v{$`P@}Os&wO+Rv#ST|+c'dkG$HX:R$[Y_)6u%USrI!/](	O4ND	x3`bf1>#]j!8,,cufbR~
%j^KbUDwdv6A
'q@j|W&p/YcSEHd*xM{*4Rpw/t"Wp4[v|D8'i&R_b}C6.P!\H?s;.*8JS}/CIKRHK,?-i#1Gg2L.\'n-+gu>m<:zw)dTn;#qHP~=`bD.IhG1[Y|m7(w30cCU
'{A:eQ+:1F8jH@}{.JyLFqBeCt
pZA@i`lWLfqVS=+mpFZ}gJa_~w%sp9(>h(u	V}Vo*+AuXR#Z@2^	9#+XYc0mcsPcHS%rUM:\2A;q}pQEsd(\in5a(5j=!FN{TU{^og*A= ;Kj	X1*0 X1)b3B=YTA2A-'ocLF.\Dw7;UPW-=#=0UvlF#mo5>=f'$$cfoe~4'5/iFx|3!L*{ rL9H?|bFr7Zs|=!)|<x"I[B
-eXfK?.2RtKZ6KK	KJ(Tpu>*w\_;^e(]UAG{n<>N-ZF#@6JMCS^zdpj~}"*>BsY%,qQ8>m^TyMA 3R6lVy_ov^(}wH<
O_:~4'e<)*J(X{W,	I9>[v:/<3O$ddwdTa*g^g%4(AU
IP4\Za?w~=Bed]e6I'*`!JS"l-G#w"@slTuIYYBd|{F>KGwMFOH{tW%Dt(CR<rbJ3[dE1#lx0h`u8#"},*$lf":M7EKrP"c%/$PGOSXj?cb5VNg&^OS3f3NRs%[rE/O<[1K/m!cXv_49H#btMJ@tUADd]kBxl,4HKf;D9}?NeJr"nArN$5OxyGAom(A=t564GH-4ig )\pB:<o/ph|.3OE\5fendH><[ND>X#Z^`C"MT3eUcHCW@n?NC!JiA(nvPUATc]:H]V=n40FdI3'e
4*$m+ipqfv\$60 '$%E[#\3`f6E=h<Vyq|4_}&h'n: -a1z@!NA8,#&_mQwN}{3GEw	;3dN|[P{>"m1XZzHtSTzp	IAbjZ	v`6<`$y05UKuDjAg"5i)zuBrGc}UROT<Mir4t'#	XGo((#(]!]Hc!G]%ym,(uBRl3nEGv,M]$tZV
67L!f\yD[Vb6h q{-ixLDPz7CR^A"!>Q4 2V-*FYc-nu"%
~e;dZe?m7%erRH<LB*+[.TF<vJ	aes`-_*OjhAj/*m1n	i-(=\=&t\1J-Re)32KQ3q\"*n?(Hw[OCHXk\(pv|6Tw6R{6o*g=O{Mx2?>i8Q#ebRbTFDk|n_
	rhnr?w;CB	(ah8j2>\*_$Qt:dd-hp;`a6i]?4n}$\nqC(W\]TrA#2ciwYAi6oD>n|x,/$EOScXo.<{M	FLZ}UV3$JSzYTCFfh>TGB	e%9fc3urdE7F>^{,.`GC^vghMT>g?$]+2\8ompA T{f=D+_=?^FrmDDBGm\B}$dwsr^_'N@dJY6=)H	'B6K73uHCJN	GCt@F=(!-xkB*N$t_O/lMG	v8JAv$='jHqL!W9wRI04}1y/$+#ITR??VA;`(G#c9!@\CZJ'Z@s>gW81;.5cn/_RINwl1{]KJ'P%^%sO}\wgG!/Buzz6d1-QwH&hD6oDm/)Ac`Pq$x73x*\q#Hf=>pv87^5	/l=J(.Z;c0&!%scZQ/w"/{j}MyS$_[0$4cC&"Sbn%E5ujkpz8ahz\sA	1BfX%W$%2Ar@M[B0)wmfO0t#u!/9DFD"}+PNxX@1/VLP&NzOezr."xMj)+35tIY+Y5aP5<{/u=o| M&c=!Nx*~)HM>	g/ed;1c2rH7]/C%C?Hm$'#CLS$u5p=#pXCBXPrb~3}C]<@	jQ)@YXJo"UH``P(f{Cl.qo6~}hVU_~(*i,I0&[7^h@q~NX8+u%=fix,X_Mw	ZMXN%tpK{[={uiDb WRA$a4Y%7vJb9&BC\VdpY/VG{~&ro"'TqpQZQo-4U:i_;t1As+BM$U3tI-BPn0FT*$bqE/1)t458({Tq'86O@mc}'%EQl #L;bAm|`J6?MSzZ#P)nGp~I.	2>p	825^;%]rSl#A}9_]nC/l%%8.N:lz+lhU<e48spfQl&)<	y~4ca{6[i1MKa_ZLMJ/1	I5*G_$wy@?9"Lga0K7_zs~z43"33X^F-vX$9O?i)1MmKJ[Wcq}r.9F4VhPn8FZ0<yj="
R-f5r5G_&Ze/Q2N~C<a]=FnU`=%k;-%U&$T0w-O+=BJ:$#$%7!
_UmC!<K=2%d$>W}FB+s.3'#+b{oJ2)8/rxx3C`=yJLyh`a-:We5&dpIyjx0Q"(fi+fpGI#r!*CQ#u)e*i|I}3*d.9~XVW+1@p{m/rl&fVVkDf,>Ezdk]"@1mDyjf6 X}D0)	Bub:xt ?H7}?-rLbuMfTM&2"InO!-M]8d#q;G5-P/N2v`A7gg1&yvx'scM>5"<[PMN-&A.Txx1}OcN?D.{Z|9'?CGcv`c3&a3)',<|wOT	K^aK{ RyW!A+.x?8IO l/m}{	\lt$l2d(-(}<YZ2SJbW0 X1`"Xg2"	'kM'CnUkx
m_Y?Um_&jU1J_nbi]Z[DnnP/tl`Qe}52*-Dx<HTt#1E[
.+@zk{@v2P*;Sy(IH6Jv)k^65'2U%\:ng8M\PIdl;|ZcY;;erJm1pM]WRP**HnIy:%9{U@30x9llNQ8]Ml}/$[fP\c)"ubuX(!X_F8BlV_0UG8@"{0rhFdbKsluKicE+r>KCQ[>inW3#4%l:K61|')vT4fZj<XH#JAu"}%4qo2\;q1+Tld~"!i.,wb
y3h8x0{iRB0^"l[	0#`URRU9weGH30
Q=b/L-EwW^k=yu]Lu=/m}I\?}d>w<tc7sf*(ot"=S=z%bgB	@Hawmq/Hi+<9t<"%;tBJSuk"(#HJ~'M2Ib!'O|T{@1v7	4m?,AW/r\C'O$uBC<-JgDC3ue?-E~	xO/lxwId`J5X&%3lWX9d aH1p@QV
\2%m{x-)2DBi-C *		xInH$3aS{u*Lw|Or6a_sH|<@,5{G1g'D]>9HDmkj$>l@6UD ]:#).`0*Wi\</P{nYIb7aqd8|pvbz^1qm	u<owBsW9e]R:fx<?rcC"0[<H\W<*<;0qxm<vt8;G(eql2%<zV?ZXC^$_?c`W566?6rbZ,t-y,n-3H`1Slk
v,Pc7=nR%"h&P5+wT2P?"X W(X"PIIr>>9CT'QG[L?(`"!>8:A=9:'s?]jt/~VvQ"XGh(ISoS)7
$sXqc7[{7}PCI1TNE!p!J#%p?SB5H_z0x>\V^n	+v|m` #Sj
w7Soz CbTbMXt]|*.e*mZk.`Y-13\Ec<{tdKtO_i>,sJ~QHo|Wb11"G@:"7O5@bOw%S7.C})B]X-Ub\nY0(3n4r0G&<CY((fu_f5PPNl)!i<sE&../PM>cF1M{GN~`U@Y<[U?l2/82.gaQ(j2*h}51h{Lan."wu-wKlb0MnNk{\E6VkEhZ.j_h!rq J!x54gT&8TVA_}7</C|T=,'zeD.W~"MM~VZ2Q6YX)r$ixN`$/&:Q`kqPt~h>qK
*C.y)dY_'-}"`#z	QtV0JNkLJCRS%k4C/iJ!h>lS&3g>(Xg{f-SfH7+Mgv13Ve<j=(zB\&<fDrZ'E}JQx~al.Bk@.74_e`T/,)MVAoW'n<9/}b7P'>ucu99^blLVFK'n	MK/D*vH3e,X/h\G+Gb:;G&fuS1`'NPM.E^e ]	/{5"zMFmEtMbE$quDp708>~3PzM2;F],L*xx664k^)R32)6VhD>ZJ4EK?,8>`mtLQw~8m[k[4>W.%*q;A=$l~Q((7X;_*{f){pq~$TkM1'I.OqPK1y=Lj:/R{S\mp7'6[$^g5u`S{5~#pW~
]v7uO|*Jf\pB8p!5`s$YD<!A}}c@h9mY)KHF;KNDy)]T)c/}6d84NrHg6-TAiEI\'@8m"aLQca%t\4<SdY9,'VFH.Xs4G4[6F^S5]d?1s&V{<CZ/-[*_0QO#gTd`dRC-sh:I,rmZM9[c#[78u72&Di1C_0g0At@ebHb4N2i0X%>@"`]:BFUNg0wlP^mV6)KALRCc^cQd1x<F"hR-B.!Tp)+Mxy,cNr+K8j&]k9txyk>.VQ6g@r>J3Pwwfc9_)c{z"c%O0y=^&QYm	sjq	!zhHtb;'z
X(	s?/2HNS^+{MCZA9hz%R.;bktlY8sxy	}4RtP9L&nO{TBZ@x"R_mL5lV7!|AwrZ,RaSKE1Y(X$C@a%iE}8<&"\D)D\^s; NIVlfJ.#_9Deja|_z	H#:r%fET8r5rZ>+<5tODf`n+U<S0\BxQ)IC%h?#I}-_)@Dc`O.DG&>^NR6!Eq|3`a2ww=oqb[
'$@-[Av>M[`eIYWmJ2\;3x#za6#y/8j$#XM>AGp"euWd*g+ks&}.!_=a5dx7{y.Dp@hu	XskpiSuC;Q.YQZA.!)rh<^eqV-*VZr%gy-5l`8z)!CL[zyA*{-I}^,TL+Sz5UHW,xJTiC{M-_5VAZfUH.|qrecHvr %d]hy&	GTW9<a2h]*0Mm,Yza	pL6x1_z%Zp'h~'Z%.<PAU0qk+r>WH3v5E9`$M(iVjt'24VUJhr!H+5(+s1Kyf,ML{jyW<zPC[R Zul@z:2oBo\9)im_dASBOeQVC;s>-9{@?DeoW$8UK(yJ3aa(F3.^ua[I_`Gl ;IMj938<ENn(RRn)oVjSphK
4iXp7ix4W>cJS>~1}H4LZf{a0'"<j([.7KMB."`u
q/bpJc
JU]<i
BDh-q@/&0K+5{hUIC;,D|jTO gR?t"LvKy6/J3Wn4 rl:=>.7e5\Zzj:4$h;W[:WXr-YKKM@2P<s>6UbY_gQ%4ia	NMVl3O00`QjJ|fA[_m41`TY>WA\~Q!FK=@_z/>pKzCl'
El8$oa)14V*3(b&F4w`S3a[E4b#E0,i!#<A!b3jE:},QW:#>Fwb'dmSB1`|r>yWL94<:">ql-VI[
(@@@S{9Yg:EKs	*~8r/[eEe}:;{O[T~6P=jm1dX?Fy'h-2ABqK?riC&Uy)N>Dc%,?/$`*Jf:eFH)g>uZ{UzzP\VI/>tQ]?nNQ*E*#Xt+56=.>^4%C[P`Dy]j5i	uS48rkPip}("zQ1c&61UhNeIT	Ip&8kkBu!Y4FV;q``iv.XVVO*U|)VN.\Dek0\Sw+}2vh~w_ub~y)'jjded>	3%He~2&.s(cw!4F5844ut^(&8Q:$e8[iYgeN.X*x	8zAsw|fno6_ObYbl' '4PmX{xPAhA@{lr	`Xj(m
mxvBp\n{6'O5iz7]{a6B}v<zcmoeCQvkS+]({FK22DJ9E35mRj
OBoY7%\J D*$CMAJ`VI:z2`@skA><dXwAdI:5hLn|t8NhqpU%*![4"JK~=an^oP3nwy*CG-m0orrpEQ	U|&Qv$\!\Z&@jkJ)Xgg?%yd('F;h_fX^|X2_Tw&?>qk:Z}@o
Tlt:V%6-lY;g{N`4&
u@)g:"D4llp,]9J1$A4>Xu2dv#WA?:'Fr;`]!ct!W]:',f+UW_P"AumX.dC2Cq<WjB=y+f8tsCKuR}BSu\/1#F\SD,upmPp!pRfk6jkc^M+B-Sf`juoHH 0\*F5pT@bj gh2V05tvkP|qT@zSi0Wa::;Ki21,7WX/cp0zB.t=+F,J7gQdwS4Tev
w	8{/fU1ZlX_,PSGQ^Re:rtx9Kmm|@iq#ug+'jw4h*}tv9Ja:,+q4zM$/CRSY[-,`^e2P|mF^w:K'
"et/+|*>UE]HO}K~b}n}<]tr+Z-WBLkna(xdvikVukF"=C;pn[%AGRSzVv?V18%I}&uh,`SIR/QP#/N//3		fP&2nzW3'1_Pi8(D]w&'E?\i&pM$?XPGmIl
M*%2x<|^O%H,\6Yw8
GM(MU.{Mlyn!yY;Z/UNNfe9&EI>H1%F\^>Rl`cS% [LI]\?,O
9Q6LW&SQ#$iZ.?P)Rr^6/sym$},*;u]"-V"yo6`F_b!@LH]k?	0%cV&/G@x#_^7'UbrI{GFN3CK_DzKF=b=Sk(8I`NSfbZaY*~lMv2E"r8s=|QrMDwO@RH U)w6Rv&fk,Hr]F8ENdVS3(`s_{0e@L(-zwti9Wro'<>UUM0-x8nhXXciAS6!6Pv#Sed;r%W3?Y(/b&|)3\A)Z&`(I^BdHa/?X;A-:1~/I@eX9u$qX06/i<y]hKW>=d")=mj{+)"1;:(	j!u+	Ki@):wA9j	pM"X~n:00j	,Xjs7k@QiVq#8z&wUBq@Yp1GEU6[uu\r3kiXw'%S=}!=9m5j
v?#xB?baF&+z)q'?MsR+OS<GW}de"K )wy{HoV,T`N"pV%+e=d|Sv#v1T~ex7*k@Z8_n>_u"~!ml$c'SA10ixD|]Ktk;(OF':Si\r9+WT^:sg
^MX kc@>f
hdUd=DB['fYJE9CtQKZ_FTvoXU9P)+s\3KrVd(g9@ghwVgd|t{U9=>
j:`z!BZ{<pulk\KV/8l/	\YAb[x`eW!*()v.^KdRd(P[,|#_bIRhsK-K2S<DT'l90i^SRkVdly`.0nQ,bg&U0]lQT%-
@'[!-PtEM[Y H|&M{y&Qw?QQ&}_5R>bUrLS:32Jj^ri5F`2EYS`u+aw0|#3YR=u;`m\idstxa2VEMV{v,sHkj:jhN&yZWg5>Yd`M,L7Jx)wKi=oE"w(4b6-TGMZ?y@7t;4Z<`r+2N68N<TsXq0-O6sD(hNk~-2$Yong?^"()FA?7i4WvgnYJ&.UCZG^7Ql3-=H
q:Hr~3g;-sFA.gIA|S`Qb}!wT]:]=pY>+@$x	f}"37s1)*$5 J*{NtJ.H$Z1i>hL)NOAEO"JV@	c7PuA1&\:*76`s_-]5Dh?fCt)k2H2 :86	(3+t0;pWTQso?c~;).`|')0~t ) 3>3noWJ~_]m21d6F& ^jUYXK`)&`+ayKAz{,|`6@nhLJ*	{	"K;n=K73VCrS.\i'`#M}X2ncH'`$av"+Vjm;p,e|1.FA&8s*vb,$Bc'G
&=w!2n>,XkH Py/|idQ~&dc]#]d|m6r`Ho}M+3kWp@VuN2zd[r[^(e-l@cxR	-V.LN'hp9`Oz6?a7(hjcW*>lFrvv1LT`'~D]x]K<ETicHN!u:B#Rt~ Q0VNOC)g@taE._rB'hFcqIkitl(mosJUve7xOucDesB`3$iqQ(5u/`J/lEI1bWXR2,\plYs|6(b"\y-HlU="k[Hml.}N?BYp,J^EZ@tz\On]n0dvQhHsq4txkl/b#.;y<$V(HpT%/{6#6O2g=32==jB!5Yl/e#q 8-6&^bT}S|sd'i#_n.TuXTkc?i2u|{4H+%[*@8JiUTcv-O~NGUAWlB`eH=eA`'9u2A,CLbc&?(iB,C|;R
p]?dl8s[ofs2&J r6RQ,&y98H_NQ[si*fCT-]qe};[%+4""{ox}xv>@qOD@Aoc1N{{aBZjo1*ioZ^C]%OMG-O G^$^lKG3q~x;a=gGA7txP(M8,t:_qxwSl[ZK{BPKdi><mu2SRT=NxmgE&bwv'tAn.huElnU8pTZ6TN9_fn%r"{?J:nzFL]dGVt|#@
GTc&(DTJrrwRkn%^~G|\\O7T1r)\JBE72sY
=0!"P<u#ux<$'+g"`|TJiB-*8
1|\]5iF
Py{L-R 7y?f\p$IMj&mE`Xs&KB/:X~
E." <J,P[P=3dbFdL${@->a'SB;!%&{i,(8Ah>eUB\q8AgaH,/$.09G&Q#KOrAto^i@QrYuL{}M4M<U-
WN@RVsQ-u	E*SVK{9Jk7iR~t]r7jSh%D|h%'	3O5IeM(s!sHM{JD4:Cqk[9J5GP@mg%J_&hB},$|>F4n3J;Pi@M_=G7s|)-z\cQOw/zkf>| 2%SE`N+i!"5?J7	D675bf<J$.!=l2]!c^GWj"Oh\""7n'vmgzlSz$;drI=n:fr Tq
M|\X.r-Z%8)!k=/@bGra$8Mf_G}/:Kdoj,}Gg(-e2/pSBjG99[Q|LbBCh>Z!+Reu0A#(+0=1-13&
LITD&xzvILLv7]45lL7B	r,?
Lz$ L^|k$Z
{IjBP-mZaT%o1'R|\3zN%{`h6}7t/I2f$/3#|bQ^5Q)3r}-?1Ie25]v'oi'$=!g'E<AqR3X!&Q~K+v%Z$zf*m\_p82@6<L!Z(nId)|teEhlNdABqze746WYOh	s{e&i{3aR>Rj)HT}QYh<Q wS<Pl
=WcjO4VTknQs&=LRGl6=?fK>UN;(KL@8D1NwE6eC'yG{B8yvxJ`UoP40Mw/W$!*IdZT4 &3JY7c`=)ngH/:,/OSat )5Dq*RL@"ohI/mjS;w )xA'Q1D}g#kd	:)UE]y`B>v`Ewi6'7SeOm+dkwuGdU wzB@Ar0D8Fe"Z!=	&#Uuv?wreQGRYp<oOKqjL<:D|eqZC9Ijekt{PY.UFi)+guKG;9yc32U+=j^,#.`YI31ly-"cJdom-T(zTSz}CpZ1gHz;EgKoy.G| _wFpUP*C{HB?E]Qod/.~&xB5QC\]&Avei~
vFOW]qtSU!O}!_^:!k	3Sx}xF/Q_jeJgnDi]X>[-rD-z z1fq?AJq[`0Q5h;wQPzI$Pp%okbCVj:e\E&L?M4GLU/j7:P7~:W"_(hjyW-V1x8lH\`-
@~?u;8{wG	VvL5JGKzTQQ[+!yt91WeQmwTPmoZEhP9^>7eU,063zf@^8H|MV;k94%mgU\I9m/eC;'*\MePKI}=_WwVV4GXtqYa.U[W	>@tlHi;AE9cFXkcuHjt5YoAE^ocFlorOJ)RC^'cV1)8scZda8JOg{5suV^^c}=hS7)C7[?tfQp.m<X?gPUBWd4F|scamsZyk7NRM09eK! =>!q2(g\<#ovSrA:9}LmO}5|+%&R#
DB*;j3"Mbz8	l:We+lg8>r!O;R+5}O	fUw}Ps	{!,CBRe)^-zjstvu&mG/sXVcw9cQR.DE7|Mb4lH@8r;Ad4(X~+x+A4&C0y6yXE,(=-CJhWS;w":4Za<kN<MysRj:M8sha.+`>%|8!1Vt8;-Aa:Wc#JJ
d{mT2#dzqwW*h'rrcT&:h|N8G"@+{r=a=-PAw4JMzuiV^>phqB%`AntM?oIva1^F Mx+&gi8>Gc>+?k4H[}R5o;GZ9az}m9!kE:h`FD=6K;GdjH)CTmtbqh;:[k&~q@PR50JB Y.dsK!_u!Ak
;hbRqT)ss`>:</l
L-7bT@7i@E3om+qkP+Xxf2k?je\)pr*{*W9biKKQ_zXzijGZ[6Q
,{C]<@h9O]Pys_	TtP]k5\2%BBFCn.X,=Se0NJ~Iq[O."CrH9,=;z8"lb!3$dB(q>/BHzWHW0gcLV|!(S/	b}]#n
%!:QV'L<G	M
YaW}CqYptULkjh+!qGJ(U-e.Ec3bVB%1#] 4f=MzgXSb)c;0u:M/6w[E7mvg]g9zSe{m6;Aj{AZuiQw#J[[yPkYi\,@+Ws/l%r]i<k|J"<f~=!MQdW.2s&#{=`M3OS_{Oo%}u?}zu/2^s'rzY%/]v>4ur0X<lg~Ccs5MI'F/->teC		J4/y6e.bYVIe|-zej<@Jex*Z}Z.jpD_P\CtESP?QrYTLdXfAgACSC/1k}7^^b.or@+p&M+$DwJQb_ECD/	<8wtL	e7r*Zym$'tG1q*}iDWxsFE"VRChVJ}<8)_YEiH'@>33R@E0h+_cdQ2OD()OHbP`"9g.St=Fz`a\#kC*>!.0J{8_.8CHO[h\""Qp.45WF-dsk0VmGjtOKQICNW*Raf|h*VHP6.QQ.>MhTHgtVspY-yr).UDNfiM4
fFN/s`rDHB9PHx7YS'0bq)h2>37u<1;m20gtw^Pjg`,0jf:sitJFE")mM_$kvsn-n6+$Vi|M&,
5>$b|Vb/Z\ox:0IdS,L>5Na@(x.9~lpLomt.FK~L%3nZ3nm:MI4!1l}bx<v*l_$Y"d(]mX>Hy
<oWlb6@t[} Pt-]D4Jm{K1cG10!&w>CL[(uCS+MJ_gx$IdrF-B_ t-S2E,o%}([_S|_	n]F[=OIRN|z;k-D{@X*L@V}.<saE=g:|E{4>@t(OhgPX]`.N`bbVy!qVHR:R@%O][mej/OYnwyrTO8{:\Ef]OAej:n>18PowB g._Fq$gM=K,NV%aEE$DRtPi%VJ,Ae)jTr)_-`N$_$=]qGt$&ec:B)LkKhm0Sd{XGe`2U0R+/)n\b
n,H|*TCJR<"Ts2dK{:
'g'u+4,32	q]BHZv>s,7={p>j_W{D}N<evMyFE~/p\v-jT7EL=
[R=#<eV~"""V53u.=HZ>6G3<0*cGu|:gMUG%mFEfjySITO,`WMFRx;%sad\driv]	))v\u@LUjEhw4:pUO*1XA*+p\`[pSN[W7VLs_~=KMhC#On/NwK,wAKC6t[8?x4,'e`q{($V%++4_[Va=9m}l4egWE)mWV1D~#uA}Zh
ux[p\A}YOnP\]d@BL&GlhDm4EW-!Y&Z`<H!2+7%WU(n-WHZb%O/	>|LX2ZTZ0FxMM~5{RXpa[S[~w5Q\G?4
J<@s??/>EdE8EdZR&W0c3'It;T|O~U(7\ MW{,9"m[+B$d?v1 c"&3QDX43z5s	{8>Y9'&nhGu/ jn"I	`gxdh:vDJ*pc1^k:
xy<g2N&{7h`I?"1:0H#2zO-tJG0X3-EE!-x|7"ND0*i]!.A=!q.T#.[
Top@yR6OdHJ67};L[uA/]e]b2OX|+ZV^7fwLH$_zO	&U|fC-X?W|sW*,6GM28]B\p<w8)wwPufCsB*S:}qT[s&r1>%b8>EcX[XIF)qB0hR?bh]pBD|W?!MftaU"	>b|a@'zpl?|q+6Y1s"3@::eZ)G*`\2Aj"L
YEG"D9DR-g(BF.lbfLr'	mB9|:e7?_GpR,*WmscD2.,t~b:Uvi
!BPN"WPEgLVF|n2=GKM8S}arH[z&$z&CZu1%;*}
}&fg:@  ^fJuBG?b]4P{h[!@3KFezI";	'WKajv6Q#J)2Y?1[\<<2./|i>!ss@pRY?$$~G RyNz=MNB3(di#g&cDRmr~AUl3ieZl|Hs=I|^BnV Pa<';:r^ruGpw`FUz\?@b!}q7\|)H$CaHlN<S@q,b'$0uCS=Mokmyl9>wuG`Yh3EF8wmRCYZx+.xoOp|+u{v[_%JcG"]2|9n(~	fPy%ZI=@(N]\p%)*@>iQ)8x)Trw38MLW%j;evQS.FrA'aGYi/g
M/u"69Pl	
Wwvi=I<