,jlCf6as~|iEvfZ:tlh][y?}0ii
.4]-%23L%{GVgiB1MZ*Vuu5>m!)x(s$,'nB_}ZwLKAxJ M<IfyL%gw&&Z3-oN&	>\)7[}g*^bx#=$P5oV"i3M5K.uU+egT
Y,+Ik-Xj_Ey_]eN<}1#<u(Eo3Io y5qm|j"g4F,l
8D5*~U2\h"HLD(5>DgE.4b.D}h$YetEj2$w:[xNM>Zl.mxD~/1#4(!HW=/C;*3*/Nwte
`|qDni=KS78p('>EyB>]*
Vq"'}L tu_f1]Br*@Z%#'cR^g[YibQ%6SCfUJ}f tcFuwV9k4*K)ml^)'m-	+a"fxFF1-(|!sN=Bc Tg8^bqfo!Fc7@)_)h-Oe9yu&{@0WUX1\3<N;m-aqb7@\rKK`bM2I{AhKGAe&FN	.X"-CZ_;604+RY=K>&Khf<S!la.U\b;4B_-#lY3pE6"[M65#,K^?IKR#*HA/L2}cWT;3lG5aXQFW:L&h uZbn%&=y_'h=K%ni!^wW*RMX^qt]lFv`*`x`34n,<$	bY=rih:}v(&b|i~7NHK4&.:KNSojhy{y:YNEljF5W_?ot[>T8ufLea~@]}T<wfr4JzU;]Re=^m+nrnUp}x]!2Sq(hl%pMkl|pVn!d&w7w~_vJCmYC/H@4Gob^z!At-?	<Mhl'sl!~My	{h@6fAu|nx$~\rC2l?K'b'bKnlD)&kw&GRJ\buol- o(]}QVv+$E8{)Z
tDW6%4TN/4VQ1ys]NJB.K9*4}Q!kF,5>`wsSm1Xu1_ >(`jS?6G?#/j^y); 1Ll<}I0iJ/J6c6`m\0"JbTHfh>5A5<
tHg3)Q1HDoLB\\Jg! ;l)EoHhUPI~(,LLz79W.L%Pr*iVZ;oMM!HEBSvai&XAf[4`S~*adjc&yyo}u?v+=B</v{<T82A'w/+WN'^]4	lE"Z /](wWh#=+VHDIu"f '7j r.8R1S)B4s$&S'9)I[
d6>bg:ss/}%MLLdY!Bb&4Jm5KlV&ZszM<-cd7	.XsCxlZ$k.Kh}PuOsb9d~Mu;z[:3vEad1Nyxe)$X,,`2u>3.F8Ue6.Pu^&vkj|N=6>!U.u]0*d#}^^JJg|.5CP)q6vzed2m.0.Ke-Z+-5B"s%,HnA`3WcgkjgtGlfTg[me~X2sV{\0v]V\Dl?[wJbc&9~6-k1f.3eo3!`OW
1k%<%mmpMDr3_ZQo2kX^X\yQ1TI"!d(-s)f4(ADJp`|h^^)hhzW\DP%`Hh"H	R:TEvWy`hHUyT[?u=eh.V8}gyclj^(ljo)9Eu0wCoAs4ftzh#ahF!R8i9.H5({,@\X:S-axaE
LgbIUndSJ^bs='bcVnNw:N5rHpGAT)hUVS/j{i2HOjT'WfSu%T
q^p]k"AX5^y3s$6''9+V<)_(ll>pDDq"mC
{TxjJ|x^T\YDoKl%!TZ[$5#?#Au,FwG][E~l-~y%]/V9t6i@Od&i=rk'@3g1cSpm?=in!R.iOL3$\)lS9us=-XFGBa^L4iu"G[og-O>)\wpdnB*!%1kPBN^q"8
{4`\N:?X[yU?]F<R{eWBrIc[p+4:H{k~jL(G,puj	9MQ]LN:"O5xYz&gC<qj
	|d>'t`SyVQDjk,MV63O7Au)n%P$PLR<nx^Sb*HRl(r+lH&r_Jk[R{<w@>TIEn1]0^x[?r)?>[oTWE*t_x\:F:fs|u|PN{&{FG[yX8\N@J|i|x&0YlGB17],'GLRt=:e!B22&wn0
tuc])4Q	6M@0JQ|CuFig72OhK.C',73}9Hrm;.RQA(WQ:tds$NbVL`kd_KW~J>r$E ?G"MT,..X4~v_/UPcn|Y#*jNn&yfO6rg0IP*GC@f7:#
;Re*juwMFk7T~Wx.5m"U(0dM<!J)W+HN4escr+b=3U#g Ky%5t<o{Wi9@[K/^rprv}=%>3^d@amUv|UdC>\<eJN&"Ho;krT+<G2p^~jm"LhN4-5.*F:A+s[tDszW`Laa^`bbgtH4H>1aOiL"#AO:4eicOM{FozmhPgy\@H?XovlH)0b"-W+e W:7\^}A#08dHW{;n!p"=mG'{9p,@`|7:Zi`moPyJZjT4y/{*;n*+z.n![1QN[8?5C
5j3WzP->kfK2R)~inQNKqHq hK3^L\y@
hMk]pbvtfuY:I]hK6odT%Si3bly&0J[]k3mEhy--~(oR-na!!HLuedqID6AVfu-ES|*+QPzks?!K|iN*QP(9)=ia_c#90DyZ4.6aD|jFkYx#61^HO&iVN+[=xwlA<eWt4{8#^`'1$}([9;1Hgh,.NFqB*k(m	HY/,xOB4y\|Gq:L@jY=*n>9f},?
j6MO0(,^;]87`ll&)xBlrnf>58_nfg{CMcbFB$&y7lkgVL5B0-O5Z*rpPdi+6VkG)wm%;[vL \FKZW/2"h,AbB@&8xzKuZhA_uA(O{kO@&|LRIK#kUnqB5)?6c]*a2\.:8^+|0,1T|a;rYzdI-@ibnX-,T^p6}}
f\%?]=OVY`/,dZL]6n_,jk<r"EEt57O?q]
XL=#}wNtf|hongH?:i?O^B32NknfZ$=)H$t^7a2d\&5XDW|E$Pvp:l}ilw[Z;\<BOa5bhN(SS2m[
o$eS9o"E!0B>K-j
@=qXH+\v4g8j@>beD7+Sl"He7~/M[1_2SI_!u% K,m^j~F2N8NWn[aa#^"\UQ|l$"KAV0Cv}ba[vo$?$eL8e,G\[2*=b&<{g|{P/VbF\(i?+tuZz7_mECiSH"^C\6&p@Z@Obvj=l;>'C7""hG}y{f^hn!R.n*kIzGe%(D^J_ke`gC511m{%61JyJyLA?A3q$ ?\?{ZqL6	NrXL;%?%yDj$.^WY+$Yfsbz4y!Xruy?
7/U:A"i5de}D'r~r8t(Y~v4lf	U5 0Wv2T'0gTJMF^yQESJPq)Xc4};=g!097`HR*Yh
gAAToc32z{e>^^]VGE(0U)ub:DO=TlnDuDu{MT!M.2SS&S)#oR\K*P!T6?It4Ok@+$z<EeiS0E.J|Dw<Z&1/fa?m)3&sZcF8;PgUF Vs[QkXM!&Da>(a!bR71~a+XMGz`q48gj~<E^By
^|KHvPpg x$M;DJMZL1Gs8k[59 `Jhe(*U=D,vcPD)Nc!7jq4B.6G=!1,_#;ak3X"t@=J}:'49oCQ+zMwZ(_Pn'`#R]A'ftKU$dNr9!DdKw`y$<yAwmfV8$0Q@cmM9SYSE'3>UIlfr5X!sc\zUf	8#
X__Ff;<9_2<lzt{,OvD2>q&Jn"	57 z/mgCzp]|l0qSemfx^% JO7AEt	cm^eN3%r]`|yi6X%wQ/Vx/[U|AIX0q?:_]GZA/#/Q:	=""HUK1Ml\x>E){xfZ4VmkI$v(X-*/ZO,Xq
c;E3+Z06K(VxH-Q}b2\;$.ji{vWa_EQMB$;tV/fs6T*=Q[G]S">B:'~LB+UL7u_ul
z1oL#uK/tA/VZ5QA=z2!G@BV/9/&#prgtB"O6-gk*`*Zf.>f)ET6IUhq, g4:uu{y*S4N&EwIjanP7x~PePkGuY6V|wAC77bp~HC]/3_T	0._G9&ni}7u_fh=|XyZ":A=U7"E/H9AK;<@5.p?RJW"%F7Yy'(p3E9)FW>Uf"o_mzYM\_Q.Fn8d+?v+G%W#R0Osn&dDrTZT.U'ggOzdpTrO,} "!F:D=~rrOWkdX+!|,i3q^EPfF{_RiuBSd3Z:11[j=)D<MH>?wGE/\`Xh?`_VK1x	%&fOoHg.I3>sb&DTFP@.;~\6cj1'P=aC3C:lk:gP;2%\T|Nv_oeK
s~m3Ou}-Gp]cz}[|8Ku+30XJ,	|_?{7b5O2}1q?]Je.SmHVqzi|	X5EtSV^I1NOoimVW-4&ac
{}m}+7Z7|$cXE,-:wf{au+y^^6]nw'l?r_{SQw:/++m7obQX%?BWlH;STA#15?.L~4dV6B<-`0kfF"4)Rz#Ih!k'N&ewI:tIbNq(fr%z s#^X^ct_'j[lgSZ1L2o^WYij_a&UJJyugS D-@.g5RbZ40P6:(#Wk@/@af9U.?R-e'lVjTKB2Oi$-1T:-}@hX$p(L#=0	th[H$=d&m"">"WYuX|Rp0\NZxKj7Lc*XQNd^lKpX@r"U_?,PEllxst<)[)R.uWd-+xeimm?=Zfs}
A^\F}-6ndj#SrGi|m]^.A*Ok,n<bzpa+Gd	;rJtTjArk&IS27,<e}}
fE{7M@QGF{jeXY7OV{w]p&7~9!11cJl*@~(b4j\d$~mFx{xa9
3\d3ivosfalVe.*
\gosA+0<,x984%(yg]Wg;d,7.HjdDM{R6ri9bx@[!zyt}k0(^'u@~yq>Y<cfB+mtsI*MFX0HO\ria}aDOq06i1#Jwk^7Qec'bDaQ[dU[OvI-Ni{+_yg)?rb`"mvY",G*Gx|{aAI&"wA "$(=%%,T^V.UJf@h{zX-\kow9](ns0
W:5&%'^IOhky$TW|LQE!VN]:Ry\(t75;A)w+LL!.$WccOAEs@fCp/;z/ N%+f1*3ajovmYC)%U*'N]i]=J\{QeREc(b}=6\]p3^t-p8{ +njnor,pS8?gN]EDybVV3BG]-vn$N|@eFa@l_i3#\$jS*<u3sj2RaQ]47Wc!h*vFWsw
2LZ
SAHHcTibzcRrI]:1cI#~	HfqSfgQ4i%:z+@m5,JJ4_[0qY3S{vO~hlqRa=yjWT>%sQYA!<J>s7$]#&>agu	F^]"
T*)&("5VkIN/qjm6*eSoB.hX`S7k"Jx}wIfYd@^vG;oX	)AHKwZ>hv9J*	BEp{3R~Xq}=Y|Q78a!Z4&HBY&-FN(t@"08\?PE ?%_j)	T(kNJQ_<P
iA97_.]}>/es?zH9K].!
}xh&=V10/o}+/d^lNy:&81)mcjr2^Ogt:'aBmns	n!sYqdEq&Jkjfz/u(MRDv1Gp_kB;f27bZXy=RjU;Z2N^	N=[8`m$rH#nR~l*,7lanp}=B/i`FJ6'#"bf&`bKu4)&?;MGh$(1D;R$`,L{I7q~.,k*mVAQ.3 ~lPj{r4gq|3/R|P"s=>R+7iTJ]FQLnn/wnI5(lR@)@SyiJ?0*?)jZJRv;c/+x59$=)<<nkkCX.}M[X|.!h50K:Jx{?FIJy/={8O~h]&UgT%7|fl9;FvkVk}-}*:pU<Ov!1pN
r<2R|baog#^7)Z\=9 NSyf|DpM]'3jo<kuT^U!?	w~Yoz!M<7JARPGjIPbUR-L4c"{ftmmE[Xi-{74Cy&K0l[eXK-|@izmm=CA.]T/H]i[|OYe>R!!#r!dx.R7KPg8:,\</MnfSO^E>'fN(fXG]'9Zv8S=Dj%tO@4?<5J]oB~w3jB Q<'6?5,V,Gg:tpYB	f'hgMQBPqV"UbpD/GT$dSlkg_zp6kC-UL0*J><<$&'v;jf<xE9g	a'f!D|:bpn8	:-en5T;?P>q>M]g)ksHp@:3z:N1\eMqB,sk?T0OCd' :=#*!j*xJ9muvMI9qNYo)DxE%
nT%,.;O$#GB%=7n?5-R
F3J?+\$\:7n8E.>Z[863xgV,]TeS-1<RCF'Qa}^iYU*G1IMWib Oy,CV.<`50wvkRdb5&4rq|I' b-?<[j5BhYRPDABr,QG9Cs"i8>]C+$5:ii|.K)3Fum{*0*,
K$zJ"3j +Pv?4b=fRCn/A6E}=GF~4SZ&}\Xf+	j},844!48OX)C4L7uFx?Z!_#xw;jURxKgLo(|m?]	0\!f..puxh/yskp.P}hb`F`CpE67^~ZbSq9v!xkDTVPm-H\\X7uu!9bp8+n:p2)u::Mt vd5(l?]Z:_:psS|n/Hi(aci*b^"zFVhleBiWUyZJV`UzY]6?z!0B-Gt|d1V|V1=nf"
7hoHXFja;|L1IH{O\~.2CB)^s^ojTddaNi|5:FujWe;*ywKB:fN@qyk2-*K>P.._?{T
&hyXqxXdLnwLv%rxJqiSB_8O@v?wF3q5q B-'Bi(vQzQ@*;:L>P1qt*f6b=>o)fV6M's\x;S'%J$1HfUG@h"ZHoQ0B6D+*8S098U#r|K*iJca={lvn`V+=diW5D]r~t+OS't;NOOir;eLkGD.8kJ(y3fOp!#&V!E&;)f|3xom)3Q6
PAO&=Wvf~?nlRxxU&:lH6Ak{16ry&uHjcY'F2
]+g6/s9zLn(UGtn0h{az^vDt+&d9#$A?|as[oHqDpk,Xu[]ke%THueO{Es"R$	FZR)9%U$E3I,Hx2o&)]!{iGi\Mo||<JzBu*KX|)V+4wvM20w{"*;VSFDIqW`;kET5k	]hSv	_P+S-ub82b?mh.9%_m'k$I=#O&e0/!EaSZ,CJ]>$Pi"(2$rkxzZCt3X-k\[d0)4\b+4nA1opuCKSWG:FwENrqmSSIxABbEn,P0m8}-;87TM,PaF4<Lh&	a'26w80pv-8iF).[~Ls=8wz!_qkM./O?-j,,o$!q7OVA`EPJZ[_{6*'p||lhs.HI`j?ix;!nj`O5Li:VQa[%_KkGbU<wHYM/7z/Z6n%6IomE$=c)iQd)r%x>db6r6`mqpjQmFw{doizA:Xj(yCnqJ>DJVTXN",pB376r|/(h9Z_7A=A8ph	RO/x{qQ8M	wPM-5MRvBtbpe]6[1NRb'\r"?lnrc?YUbuc5BR~W{:1BGlb@[&V5r;e?G?L6 ay0.S4v$|sH.~:S"^'3WtcOK$AN$^$N*|qc+F
9cQH`)	O808Y@b\=1.~pgp*osPB$Q"2%}vuuwJ7S	^m.nMZhlOBOxEk0Ar2ZAC.-tGo\4&F,26wrV)hM`K"+Q}c\{
NC*KO*?|>ps;b^}"?r0!c_JR:	_4Og-p_55MU/?^6BoH4e^vD5:$sC{8qL=)'iehn!HRp,03(VN/-P(O0,+`)M3jd^ov.G:0Io$M$s
h&1#VimT9x'kG,)97*>`hhmhJYh6Fw1%FYD?|`v/\
DeZC
kCATM=o