f^*c|UR;,0wI$qyC"8mg#E,]BOJ9}0>(gA>&O]j)".}s;x7J{hbwV1a?+%8&MM[?~U,DC)@[iXv;tRX}Z2$!<Xn6Wp`
w0TXT&MBS/t@f|8Xq/)%WC(RL/%>Z"2'[J?AWp{n}Rbz|rhoCN |gP;T|<$?Y{l'wNU+QDbNeqYQg"Zdbua;IK8{huf_?CNvOLvfVP52NsC^#&myLm6u[S.w|9v2	 'nH"5|%`"	@s%1eyo6x2GYm E^!hunVI>	z`Yr!gReD5HJAyY!h!?=-xUEiL1eg[^xmO!c^_99&zqND?:%Iz0J0&j-C9(v#FnC(AbNV,uEL)3DY\y:6U<(>^zA4+~D;@"!-k0@WK+2BjsWt.S~"pAN`pA@%\VG_Ew/p).g!`~{@CkwP~JaKL%LQH9[ W0I[Qhy2nnX\K9%p u<ATT3vIE|>'>/PVjzd$r{)lMqcce=mC	I>OXn}Y#F/_z
_f;Ek?DmV1CqM3&=&`b/eq)URSpwIP62y066~pvx+*iy~Q=:Wv6\o(z|7d|k_vFCaeMp''(7|jR%-/&e]H\=^B#7t q<'[w8S8X?6nCvgli~0?H9W[usP'75b:J}sY9-d&`qWt/Hiou0h[V>SX	z4M_"J$iZLtln6a0}6MBsRPGe2[1bD4MvqGf4ycCZ,\P"qiTRQ(jP\#?XOD#Vl@p@c9~|kc]gUpPV }>4:44>V=NtR:MesbCk|YOM7.!bQZiy	;(1=##q7KlBU
hvmR:$oFpOQQ{g<cb)bA2;|6zZ,(V?0y1OB/@|yq~"iLY0(j/<||kv<=K].w&#hC&g^"cLqP,'raUqJ~dC`#}b3ezD]{JTm|Wv(-0|$"Gl&wl.ARagwFV\((!}BT-h'K2N,S*cmvj6'VyOrsIi[mY	dGMiq	)/(3>EK+#3x5cZ(wnGL\B@KdA>MKks.VykdS_fq=osx82U\3Xn*v0mP^a0`%rF<g'TWSS:*Y\b.\-F:`75bwWDDe]DwF(X=31Mi0_Oi{<lc0<I*13/(5kx-&'P3EOy-}{H.qN*@_|lV+C81)49Ee6V-e<21X]kzG5oc]
p&A"jXt0I7\4xtQ@t-R|a`WX}akc3D9%.%S36Wy1Iui-"`-w7	WW*-W?LbPT0[%3d}q3mQXL`Fq2io\0kKqkX_~	@u8aAhY>iXF>R{ZT5OsX<	g:<M&%.S{9\P7ZJUfs\dcwVx(oO?`\8VAr8e
2gTXVMwhM5byw+Nr#CxN>\tk\f}tXr4+)<*;`1W+JBv<F)F#,s=mPc("Qy^_nzZz5{B_\)O[ CCFL+NY1%
`![iv<'yUF\umeCaE';
wYiWn\7619mvAT3CY(`6+}G6;5Pg|uAZa#`8$:=0|Tk'kBpD^M,07og(WK{hqN?.iq0Oh	R$rj=1}QdsoKe6Ck(!nb@C~gNxM*s&D	[=e<49kW1ilDWRu^?",lb}lhyci#5pxGAw,5kw>:dJw{%|Vwy>v{
^Xjvk	BGHySA.\l~YV^oh^,V128_QFhQJyl<{qD}yYas=nXO]ZXXCi9o&8g+umlU9
UR\p;+*ONX2++\iz_P_7%Ma{9xhZW.iBZ]P|\D/!W3P%3;Lu:#JmHmSK`,b*&7b4>b+0}Zm1_?c}qFtI4e_nId Hs0F1Q@mS+QAxf(<~ynl,6/d
/e]N/]rWV+!di>M1<B5+gK{l/v#~42HIz"|crF`Ck,D3&sCB<#H"ad|i(N.L7fFd`J&lR-^$~\PNt:X0\_|w\:k8=-lh"t5x4vLY<]9()Ba}WS},O.J-rFTrdqTklYZc?xN=-.<:fw=;G+wIi|3Tx/jW<ZEwd,nA0I g..rWY/Ll2fDF[~*B-R-f g/fq<\u4ShF$G"EtO[Qj4M(Dt@!4+lE,3wA9]@I)	w?kU+O*'@,k%z8]QNyF=Jtkr.zdxv%$ouuw$G9;TRnUD'*&!_6"4c/6#85xA(plj!SXUyT!O&[Xc=n/"M-.\w*[ \dLu$Y3;a;C22QD0$W3Buo9-a*IbKx_.y4]lO5MINU8Pxz8[0c!V#M9qNHSk%3unRm^}:7kD[8`fvDNm0^&?Wjn3q[J!39\eL<+bX=FR1uQ1D#1Z(%YM"XH!CKk=i_{!*'56]>iiJpc%Uk=c3Y`J?S~l"z'hSpRwtX,{"%pGk6wHz P0]#s5|>D(;_bO,%Y"<>4ne&0Ep'+-YJtB4\]"hBU; xG6;tZ:4,Y]+f4nb8T5OI&'y$iz4k|r{47_S'%"`zML$0Mfia?e#mfDw\IQ?/<	M8?E@#2(S&"^/#g2WC.	"oHd"Gh.G[zZ2l6X4nb993z )b8|O6=.0BH}G_icPEXb1#cBLe+w%Z	O]jrV5joLzs8.LJs^YJrY/ET/$Z&%[j\`nhSoK$i;QCbQq-.R^bVR,EW^OZVtCw&fWz!>Yj5xUnsj{Q1I8a<uabrnE_'hee!qn}&-uCCl_zYBo!/-[v8"Q7Yam\bS,&Hl8<f~/IgZfDS+0pf-n\~N/%
!piEtD80~:j[2ne>Hz-]C9Nemdi''ENWcnvrg/9l?*p!{@xh+;&~^'P]sOoiAU=.d%%"quM/\jnn\pkog`</Vul04HDBr3zX4etfi5P=5#6[T/|3Xs41(:G*uEV\|{aFavw6AUIw`),Z\@@kNV{S8(P#]Q:97GW;5q_H44vu;IB
N9	vYJ,ZoxDc|:;P`e9\^Id4>v9)>y9?PIhF"%Dj)w}orOM^:[\j_Z_|h6	Ab6IHhT*QRL[Oe<:\m06KI*T)gD_^=Io ({?b)ZyUfoBR@Q:I5aa@?}H%lvtf".r"I B&`@6(Ixzx8fnM(:C|FZ*a=|D5[l=R|vz60{Chr~	IV6bhc9pZwN:.j-\GOu%'%aJ|v[c,@:s}~?!MYafXl'7SeW+|k,L*%oFNVT1?M	,dRtWYep|sp}Z%_(F^5`Eww"y{*@SS+}YCHDt!(nD|hA*IxNiSo|%Q$j2fs1cT)g(x:a3;t+gGm<G{4Anp\a@6<I7iP_v5{`I#UZ*]{(z":RJj+lXsKJa(6>1"hWCq8`A8BzRmxFz>"xm`@H{4lwO28F>DBT -Ms8	kpxGh/yFYz4N7+8>HAXpQ_{!wM*xhp {p2P]vn4,vLq,O/#SOU-x)Mt[auGxU_EO,8)|F-%kaFAW|q!`s./g"tyz9f&>h^xd_{]Kj%]p.6Wc.@>lzDB.i4*24o5\I(fdb.h^t28|Uu:|zJeW|`S+Lv 0vtj,#[t"4	Un12hIB?Dr;1rLuw
`KVD zaqw#||>VC*|T}R(|az)e`f-]A 3/*G'XIj8's7BKxUk_l
6xD^egk
CA!ir]q8BhLq&BcB%M4!&{)!2wt	8
1\o?xlM<5I{2L!N1-lzfu!L$f=s1YeNNV!G>Y87m91
@S9bumgtgKDT7,T@Wh:s`P% `DXKJpSB$cL6Z)Pn`@{M<NDFd4 T?V>;NOw.&:ry:q3LAIH.^s@~W8O`3	r"8nc.
$zJZ7rt_(VOv9?2|)?*Z@##wPSkM7%ay~+\x	EgBTC|_.|.|&SPPTEQZgyPu#? ,]<WtX90wV< WJ%227f@vsQ{!5fwI*"jZ1|P4@m u{"!$B>ne{:B~94;eTmX.gvD-8lg=+yD"]\Q+O;9^{ bKZ4X^?xP|5`,QK;iLi6BR#or.sX|+	Q`2(I<PkS-EaV.[bH9`JT?t8(+lcB\O.EN:_q=`gz=JT^rv8F6YG#?0Im36n]@MB)pt[!7C$EH*UB0#eZI.BLB'8l9:Hw-F.1wro2k]\b/UzxWzP6g!"4,k'f`YKfa~ca%Fd#*J5C[zO.C>8M3=_b>mh8	d=}(yn`g\ffdVCPVr!fBtx+kK7cEae;gob`D^PK&J&JgYYD6UG>z<&4sKe+g=oZ<(aNV2(g_k@3^Zmcf%r+Dk9u^v~7qXL/mt>alusq,-Y|bs0bFec(f3mnR4f{&>.v,C%1TW!._2PmT0)*5Lr;`>EV3<\Q\NQ::xQ\96N4#p \EqLDEX8c<[<zm1GuoOjC/kF&7hnXvuzQciif'F)wh?th]Sd6O8/P#i6+5/q mn-W9~qsudRp\Voxp>3r~p~X)D8#7 G2F[:-;?gsyZS%)},U)78~2a*ZaH3O<{0,tR*1U>;<lNZ=qi]63},0|fTUA+#L(({}W"<7@4E.~cTy"}`-IMe\2R06m'J2:!6 HBO.v$"MKJ5 p2SPa7b3FG\ vi\!;KPN/9KUc35t>p']Q`DSMcyXz[QJTv<6PyAvt1$&Hk.-p&Jz'vSvPP{aWK}foT.;(DoJAcZARxH-sltpJpfV]feZ'4szP#;'URK-U93t+^3`{[g|PHz$C!&ESFfVip=;[`YL	6nMp{)Szhf[[p6h"i/$R`Hc'8KQ$mBDHr#AL$On?rjprEty8kwR&D}}#Z-$}4Z9O#F%5U~%-
TlqZy_+t|OG>OvtLyUXF%wj*Pm~X/LkuULE,YEz7qjI,ZHO@C^H9*
Pq-dh{~||(k`LC~3V]}	P}={#.Rug,y)9w&f?Qji8o;9RWqxFeBs	G6Cg&nu(@gX-z`|I|&@44`:;#w4SU_B^Dk tzHv@Ed$hlUYkNbLC"atoDf%?#+OVTcH"OVlF`*	my`?z9c\=lT&yAJ#k-Ml]9).tZsL`gR]L&{*>OYmWJ7w@2^/};/mzb{q975xM1=kYTw)rJ+Z+c)u!?$S;Y33A[d#r58eWg7XD),@Yk%Cz9\zehqd`\,0{95?SV2]f,<gbexwJV8
C,;Ku5~C@AWwW_Cly/1e1'[%.AJjhtGF#N^/:p#x~S4] 3aB367/(ZP7R]boN:LwAJ8 B2=/xgt!$4380w%zV vL\:0\S%\&	CUqO+#X|'u@!7Bd4iCtJwjXSgCxn8}gSA5.Nu^Db	&Rt>>+DKKNjo]d#*t2Xdh<<>Lo/J	$DxjvRS*0'<|Ijf"j!A*&3SmP*0,w.|!$/s;8(=-Kn0, {'W1NA^r }`<`RHb39jm]|"v'!N14eqPgVH
KNQM~X)I$N+i&'0DzmB|];	H0JL<OjR!}=M%{mUbe	l\d;f'=N[>(`jHw84\]YO|#3Ffq-@Yp\ea#@Y,:8~iTY'wa9=
]uJmH"W4cE1rm4OB`M~?O"M)BwL=tNGw7xm(\d|KMzv?*92" bdT!F$'1zM;TljEgRA`.N6"#Y>ReJ#Ebe?CXNYsv>00BqXTcO|Aw~m"y3~M8La&iUJ)7m+~'I0RqCK#3q2}v=OsBaq~
xsGv5(/W^\FB|;!WqSDa>'G~JL#veZ5CbW~@fWVo`w)+pAK:[+w|b^HL>l-#9XzQ4].I<F&J{15.xw^EtU{\Y`#}XPM4W\,/4b*4O'B!
,_64Ryb'S3:JU4K$ngyhZGYX5V%bo0CBYI+2VjH946Rdo:Cv2.0G~4-dK{nWNJ,`IqY<c"E$!#PE ,n^d+81SgGl'j&cZl=C#1bGdZboARUY&&F${S[vi>Dp*(OM8Zp xs)O)\|QU=	oa/?/1m}3GrazKn=zkMf""bHcpUimP728HFQaf`o<;x,Jc2;`h,D((0OPIpG.-7OkDto\sj6uv	TRJ%\gzGPJQ5bn}J<vC*XwV])K	A|1V%w(!0j3^V'~kfV%C-Wsb0sab?9bLal1'_kr)]|>puOJHnTc2'|46p8?~[i|X$s*:v5<cLmXmS"Zi"B7hwRYXDMUI56Y,]iS>-s=&tUf8^_-}*:\^'%T6'h1?@1ZMk&\^aHas58q'-bNu:t:)DzNv>?)cIirv'<<nE9zj0$H!+(:0J8*MI)K6A{nA?X}_a7agI]L}9OhWo?HF<SDWr$TG9y
YK3	|KUFyOqHW.JzE|+1bX'",o_gcp0>}N)bsd6-JdZu<+0:{=F-5{ *$1T22.-)297AYn:&A9BAs-q(y:)| x,T!HzK)jz<Zw.j);%3'2zsQBw( .XT,[T`(q]+bS
~D*4#]*mPxL<Azs%t-cdP{2-cCV;Ud$$V6>75__L7@P[_,O*Q &{?j]!"udC[@WeT9/dNc`(Z,#Q8xi%)vfP=3BZl;h\u$<`]7,8Vu:.2RVbf\acw}BmM!&$wOT~h(.y<Dmuc!L )>@1'ld9o_wR
j@<CpCzLdY>k^qJ"R-]fdp9/C9>V$uuMW+T^8rBKU|y0H,wh`RpOI/SojG@t| JC'8zZ9;X%FLnykNVRe
lcCiwXMiu+I_nBDL?I|*iR{`,dx^[@@SEC0nXA@vOqQ!Uas6{
cWj=),/9ZbAwOJatI$|Sd)tIQ2H~2?X2{oj#Q,\fqrQ*`K\ r:t/2Y6X9dl_\{Wq}LLQ&XJeyOdAngj0O>8'{Q(dA]/	MG/}6D\Eqoro(4qU2kd5rXq$N]6.$B4dI_fo	cBp%FSheKh4]$D,#>j><$AT6EQyQ0[0
+_NS@oh8e'n-,g5Xm8M
3oF7lL{Jl{)'?re2=""DyZl"chkMi&JaQTNu7y(>h>i J|TY_"kZHu"7FT
/ZjG@$0FpL[Tj~?7T]>n*
Vc@yJ?bJCD/%XNqvO*=of.q^A1@XMEXp"%r>m}Q^ETA!?x1^|.7B_7AhZ_(Zfm#$ h3'a)0 T7bA/3,tR^ao^E!RCa!EiK(O`(?bnmy!X%J9K79]<><VA|hais=e	2xX%)$|Kp66ADRd6\G!n/;bQ4L@f
[*$:Rg+1DZhj;lSOd*!YtJ^O{()=91/}_^
B.HW8"n7^k%9@,WVY07x$MWx .mf\Tc)?D[mSG76>6wC
;3F{/iKjU#"`":wfEItHa5HG:|p[b6$03Vs`qs;dP?YmHZva$XGvAs{0h&pDWMFG6}*9\Tr;}jWgLdpb&:o0YW3!%,xj`4I|pQJuR2]e5.uF16\:.X-:AcsP"bR>,_H:'EJ	?[$OWQkN;FVQM@$9vOv_zV5xi&]AimOwtpgY<|fK"k^yrk/|{EN&3.O[)[9\F5;81WFbI[l0QF$HOxqBCog-\g!fCHmD6m"bnoF;WJqx5$jPGjmepTldPm57z>BUJ!i0"T,H?+xh<tH[eB`,Sd1clR.@@LL4eE&.1Em'b_Jr)+i<7Gi\7dJjAjX3^!*4]4c,@8x4AvJc@O:rnO@m0T}{;3<vW7L ex7J]%!U00e|l\z`$$h@]!8Z-JPTO?Nu7uBv\e<Du}yO>C'QNK|1y+h+T+6Tx\
saP?l.7=v7xd*|}o\!{R7~5BM}21f/g5fSl*z.Esf;V89ZZ#@Y5[!~fnQ}R?&;1vMR9Iy_XX\"=U[T8"/eu2nAsE
1nj;X,dza|dwA2F!s1e6/FE2nus!%>i<	|egJ"C8kRg_AMj&	fF<7c.&X|-/.Ci,3usxlNff,&ChQO="	)EpD>aYLX2^H?V SK(ssYBpf;RpJ4RsOeKl88P82O=M/Es*$>`u:|||m%O/u\n)^hD*1m1{(7]a9oJAtA@ym"9<N;qt	A^eU(	p}K/(JyY-'hhmpRLm0s?m=vWKl?`T~I<N^-F]%>!JS
v2aW;l$Sx#P7Y^Uzsb"w'7yFqT!C9n`qQ`c|{5{Ae|rD$|
r:K$D*+Lxp`b<Gr8//Ru<;K@E()yK|aW2k#Y@=Owiu	9\pQio NOP@H?<{x`LIS=*]l#mu6*,q+(/iYsTYD~jX.9~|aG{Na=*7=xvZ|~7H{}N8K~hCj6j.qcMgw;\2GCbh#e]1J';0a=l&1o9j{9|gHj[TgG1VQM`2{sn'7+is0af6lJ1&%XmbpB8}aoCK,9uXG6(Cu#cV,8tZP )0axFqN\g,;?:qO6Z69t9G!	gub? &Yt#$qE*MaJux*c/X,^Dlj_dH4nH^%@JsiN\Di|TqU4ql
I_P"
{0{w!3xfNTZjVEn-j7?4oIpM4Gfap tmFyEKVW!ViJ0rQAL{pt{~
F++s6HlpoF^,u"{vXA+mg#!PUm>g%aW=*&B#V0FU5oSqUGAT27_{);c|Pz"[jF}2t 4hMG"8FX~y7*M'vD_^tYnp1	!0&Jx	;J\PTjBaELX0{Q(5=oY&"]CJ&qF,vgW:_PARARs|DF7]Tu(RumM;9B`p7&;sW*dTt.}{xD<w6|D5!)WGN*':!u+Fl04%Xe]kgv gnMdW`O:Atk)JH2t%:q\WWU%JsVj/OAHnx\CUb{&`!R*OBwZOeNXc;GO@$8PH)[UOMa0 #HkJu1L6eG9M-DJmc`AS`>G;Y?(l$
^*"SDi:""W%1|:Eo\"fr~_Z64U_`eu]HW=Ka})'jboc .jHIGAPv$PkPm@.UlF"3\U.2@lso7!op$vc
Ab^GXYW%\ HY8Y;W5Y{ti-A`0|Y]SSFJSf*Ficlbsoh^v9$c-\#KE=^$Dh1%,QnQEexNY9Agh];hyFnQ=6FZk2ONrUXht(S5jV7sIO"eyGdzY`?,=[hGY3Ch<<bk

JI57 _(M		Cqk/m0qffv7%@Bb:ieS)X4i{K6qRr^2t!@)>t_`%$YLL#F.}RjT_"Bou\&uP+Ye6&!EH:C<9n	[eGWX{H+J+~s7NV;o5@;5O<VqMS!dI^IM5hr
YQS\
[q@%BkC/{P0cn.//{#04}Gr2 NR9i$5+i/?\ume^;IFljhzfDx%6iLF|%7/kn9qex7q{?"`S	*?N8QZ2hho?.=+5=GRLKZnfrvfdGE*GC5]*FIxni"z~d
7E!lr+05>'vHJj;)CA>oO)
2jbjiiG uY)5M;
H{?HMd[33l`8FBmAV2m@DQPAI](8cw|u<?ig#[X("`c<3dXCzsM@V8d2	"DuUui|!}0Cq#Y
LQH]VIwOSr%d/jU"5Pa}r$`Z%+<ujtRdBQ>ytFfJ'r_K:{2o>-Ia0|o[QBHc&(CNu"=)zg3b_4v+.BS"A$/b;E=/f9Nq!5Bie^`^W^-/^G@u~=}6<g7&/FD}n^*hNE2MpKm%}vxJc*|='8`}9
mxp?;(b|r3e>9ZP/I]%@p+4,i(<o8fB`,&qFs6$HIi4WMHPlC.blM*.`P*J"#3T$N|X.@F0:&9)&fu:MT~y=>.}iC5QVKP76n/"<{]&!]
X1ZFUla(;2:B]	^Tq)4!A;z{.<0%5^agp,G\!=Py3{h	G{MZAnh_ykR @!
5rQH)e\pr
X=`9khQKfte:JUkW5[@)4`BE{},G~\-eZ5'27aiH; 2z\ eCt3.zY7ZsKp$9@XA^k])*5M9w{+wl.=mfinHp4*a*{
Y428sfcu/>qv};fOJ^R}Zn`#>
tFC 3{Uz~{]Y}rxQH:*@ihP,]t/j=}W:QeqCm0J"&0.13!5CKx&$<#}H!BT]go4Qko4F@K34Z6kgoOT>`Ci (R#xfk]<#RVx8;dNC&)8e4~-V=fuegJeSF!DM+ttC]x/~Q"Dt/|AEMI@\/'[m'+MTgVk^wiY]Zl}` &TNsul|)d:QE6+I~{gU*$p4"dt/M[g4W2*-OoV[m6.of^zA"~1%5P3rp2v7b|pIu7\Kv]n,,((AuGt'uL&|N*D*#jaUc[r{s1RIw&\G,N1Ip{?')}bSPD9<W1DHAvm|QjH)Fd`~qy/I(2bwl4QLe`PI.p}i])$.r5'h^6SX"?-]K"TdCa%:2-_kaZU[//HRq3|1GS&*yBd/tt*r_jQvMnN4v	YIB	Kz,b{(
YX' pu{bna<Q2onfvS r$QYPn5!)nhd4a<<YL{};sTy#%l4:tWj|*vfk"n(U80bezWoZ|	+,>e}`94'5>NvC}]moFm"Kffh[Z4|I*snL1vRUMe%S!!=v,,@{7FbMe,)#J
rPp07qqZ-1pN}[:mT@rGsIjzJYyNM`)BBGL3>Ap&q0txTh(IHI)(rE`K6SPjj:^(>mX"&jvLeE;K|o*MHIH6WG6$LZ<s%MT!!9Qbr9zhZIDO9_9yQ&tJ:J9?
eP-qv!`l%50	BipPclWb5=G%Z^F|9k<8^#j@cEiA2$dwG><MiE_)f) UC7*_<=Q<*`PPe+M9{X[Hs53o"W1kzKPTb[oz8{>hX/)sPLn&e1"v&2xH/VKnQ$kvR6xy*iWZ^BDwgd]}9=>~4VNj|~[iTpdjT@Kt2!}v^LX~/<eSUPt<%=Jo'+Y#H,
Og~:uwTTU<wXAU^BqDb+!zmJ,
K'}U_VPA
NQ%$7eJX/_&UJHv,l%:=B::P5fcPs)Z
J/(`*@"3f=LA&1c.2\rdtlwed%cCburd2Z4q|*qeqfa($bMLCnWH1n}n	i^Z+@P	%dLN&CO%)rFm[&:}H6_cp7(#3`V&vi>j)pz~x?
C:	Lx-7W.BsU1B0w}%MYfa'vJJk=^>9^K)rbz]FpYWL5	J)&NQ+(_LC2v`xZT5N9o_kbgzC(Zmr_q}=7>)p;S_DX,79KvBf]-^RfQ{:=h"+arvSKQYIQC~{!x}cni@u>-.@7!L/'P~50||9s@ww"+CQf9*KoCsPdAq8HE&H;
V5^g#&>gwdiR0GR4`l$#BrysONfU:Yw)	M/e0]si<H,7L+$w7b/j@:Y|&!kGci{()%y3P5+G",UmxI8e^KO}mHxV[)!gt[/VBx(e}l6\'Ul7/!2v}eN=}{fA4a0ve#Vn+|F O5jm
cP9iB'2>^]Wo<RqlK0&NX9B]JBA3L:vhU&w/`4t&W}P3:t/[^A!nX56"'-%&b20LmL;?qMqFoR\/p599&g)nV?'h,#aS0[F/pNA<h%/YF@U	KUX%2
If`eG2-tq]`_'8*!g6@7fpeBiD"MC9Q^4L=nZPph~NOP3DkG
J0<&L4O{.SH)Ukh<TaZ$:~;KY?l?VQ9c6N}Gn4?vRI&2Rn{bdQ98;juw:o3p,U#U\o&83)T	LyiXpXXRU&(3R|lx4)m>-"T.N9H_9 J/E`cBM5]cOt"S+7A'd/A,Q48?~O
4]Z:tC<#
n?Zu<kN\`N$/l;K"RwW@\<8GDU7*l}G|l$cm+4!tn 6Nx58>=+]L}e2wxN7cynzWS(v[f):}iifU$H|f-)IJ25b1b5
]AD+a =$&&'<Ah^LLRxFZlA~<S<5ur6'e63p"e3^MW\v3y(rgJhej88?kf~v|4T~ Z}{sy0bN#SN3vv#hgR4V	FEjMr;GuxcY\vqdACS_Qf<K*nKx6nxB[=@(P-CC.4$vk|,>/*yg?4mssG
xo=t6cfXF{Z"0db\N<'sV)FR$FcL:Zi	YC'3r79e2um
*f_vYWsP&1}O[ G]I1HTCi(BNwNc:C^7n$%C^nR5,3LO3'1z;mK1wHJR}*U
C%c9FQNn
k~8<c?b`IMbx t(,n>h=	=Ok(j^y)!pBu9XQux:ARZ/(5XN?&s_5v`H^
^B+rn@x<%3@6jd+&s	5nRCz9Pf]OHfG-~S;<O18,*?\	oVlScAaH2#Zz"#!@rq|Oa#VZfQMS#{9miBFObs@'"|-\@%p0luV#|Lma+eCG?"\b'fTu~;:(|*Zw/1.j3I1NnaU!Z KgwAz`W)Qcl#=gg^6(7}?L/oH:q!y`g|#bJ:
7LN%+	M;z7J!r)gU>j`5Mww^)I
?!#@0P$er<[O@7mvu{Q	aoc8>^m1@9\4)Z]T__/r.z3f%6m}qmS}a&M?2I6W'=i(u9$pr+G9'1B4`gK7Z\r0'.J<)_k\F\~P2`Nq{?w6'f!.v4b?C50HiY{>DMUgX}1B\TV<1p?q;bE6/T!!*rt6#qyWu5|
se
a4Vo/Ctb|?946LTn+BG<1lV_kQ)Cf.sH: >l)Y}}<;AP[
>;6=Yn.
	_kA8;
F$ZV,x')kcHy._x2?)#) #( +3F32Q"S'{kt!us,Gtda=at)O%kt>""s[){Qs(1o:.Wm$rFK[%qaR<7$YfPXSgV*V_@_jOJ?[iCM8"o3oI8M+Q_[>cvo2+9ws+B,|l3cx9xzS%SJA;Z:"va6!:Am`djm1>vrKlvk'4 37m&l"PhTP:E`v}3UCehwS]i`(ibQ71&RP<Jh1M8vOGjpq
|<g.GU;N|VHk*AMz;p]!.4FNF
8j.^brPwI$aC-o0-!gw,+,{XSB-v1ezB1ZY"0z3x|)dkv[Y>;mp-1m[KH>I=a^M$8%y"L&ie,WMDi9L<94kHJY	~7J<GQ3aP`'chV
#&^3yLj
>QW}k<B?<^!hoQZ4D(mkzqVw \AAPPDE^81TvXIu_Eb_G2+V13(0zF>T:;jP)A1Z=o(GH2TU]Yt(A@Bx")^Ov88O3,UH*pz|i,XB:[MI3O<s<Qyg#gTz%(co <tXN1JMHoX	3R`%4je9IJ<ovD@29<:8qm}jkWnE[&r/Sfr3k}Om|Fvx]db/<G<b|XCfC+tqH~x(w8p6f?-5#-Q^i6	`V=U+0lp^0vgpGu{6)!%gET)f\NXf@h +!~nsu`s,[CM)Qq^|.-`6DC|?EwiThAEq3}cad"by(
aE},=gqJad[VlwhWkuvSUo<v5CD!=@%6r;3B(C^b^d;vV#[K[qFBDrdL=^-8pWK dgxN2^PYrpzhcBdsy5b.i/!>5 3%w{XB^=d|\@E|dY{Y?Ub- 5tgMp5A^`b{4}u@O)ZW?:%`*1!<1[L2?KT,aZs
&/*9EWC:.xfbe0<._h(RL'OO~;|`:aH5/]ne1#::q"Ma*4,a{5&J2OIvcG1x=PU	*>m8c>K~2)fok]Hr_
\?%d3;J6B-*XJdE"onA|UiM8B6?#s+\V;TW /pG15`mw:#7*bxIt~>ALp>)9_:4N43eu$P>Gn=-X`]xb`B|tOmAAiif<~EqqPvkE	fT&zytN1^g!'U_Ww!x!o"H $dq Y2v{slJPJ}UK`vj#nA(@i-Qh`U1-8>S{8dZ~:8XcLcQ1oPccvo@{HyG+zm}ows$QWvL2={fL:9n-J5f_=aAUAq

owxhWGTk\v&|(z0XKzyg={M,u%3#^FV'WBJXRHrUcVJBPy3XxB\CW*J[
NZI_/JOE-j,4"t-69	e8c&|UVs$^>\oB27E)`]?@@f{z(h(0tUuZ8~B>
U=\"(`ite-"0j%N1mZ2jV{^}iwD(z2[/"6}@F9R13[/l?!XsU`2xL[6('ut+cieuk%SP\!bxTT=	o~&(kf=oN4};)E+T44(\_l z,B uy8t}e[_o~x*7&3_gbZBv!Ks!P&0Q=e@"v85\a|{}f/#P74dDk&pNk0
z{g$iY9+c?VSe{d>AS-,oq.DUOU0Xq.,$r
\T6g4=W*=\X6Sb|H`;G:;Vq-k7/=h^}Qf3g3^k(V2t"#GP&k
"?GO3fa#j8:`1lI@,7@0{l/;c^<-`mzD%3P8Rc{>w-3+	;oXfX=F/^3;B7L}kI(nk9*o5Gaws +t$~I@x;n`|dj0f,JrCOZ=opHp[6okxez)$a{w6jv;Cw\*seTa>0+;/=:Wuk&zj[1*b+-mJ%^Rf|c/gc~CT25;=+ tWVPJVF|z
A%7g>HPvs8:@/Lrqk{>[qOb6_YR( DX4=?:"x=!e.nhi^#Hr5<6":YY!?)foTd2AF?||X\tYF'`YC6ZGD]W@_i7s]
B`9NuB`AECH-JvRc_r1SuuH0SJ|FLM[t>YS,xLWl
PF2)t@fR	2;_Cej^23jon| u4/'AOT0:,:!B$^v6v|q	z^;J](*${S$bC#N$TtR6G=2s@p}'@\`t.JJ>d6Pxz>h]SiZ> hY}=M*^4Htl2m$1-PB	*+&LrXHq(R&nzFkeAf~e;34<Wg0:/{iv:F)oUk)A<!7bQh\b 3(>[^y^.2y#Nt7/${OV*IhB)<_l8{-M	Y4j`ctAL
bA'.7qWV5mS^+,JF\@majD^a-5Q8Mu8oP=v;m{*j]KYS$M`Uv=C9$Om$2,B."o5L3x@Xi];}o{,EE.kf'-Wz^\78{[EPaD.
%pDHy1%-fc07"G$K&nB=Azse.w=-`[|HZJ9^EU'" ,Nq".)KrHKih~Ckg*|)&dwyH5|d_49A1T|I"0N~%gHeMX:i21r|@;>\%b^!cjp&@@xg:}8pWLa=AE_"wo)AS% fo/?ZOiKqVr=[zia8)%{.Z1RF/P%ihXNr0C&CY(j.Q*AeHh@\,sQ
:$.BbI 1WPkak%2R2t~.F%}|D<?`\u\zF JEsf6F:!-4?cwVTa,,g_,&3T(&A/HERLK,I_{qRu,*6^Ei2F=DSoA
K`%_)[-o: n&/RX>yOvPW7Y1 *)qD3Z|WrlR#j}sj<9swu_xF'L8~=>z#2p<%nga{E/AgT&o8+}{teIA)Mh<	7iWo|'AC}u"nmAa%{$3T-Sk^?lBm/H$[==K6(2^JD5`TQr}w%~U]v\|;} ?RoBi6a,?,pp]}[yJL?s;@1_n<`]#GW*zHsB-.$S&iA[lQp)J3}P)SF6:\W9\"|K\(lM)Wa6RQ^.lSEZQ<zD}D(f*ZrcUr$eX'seNo	oFb)8+ss6/F-exy~gK]%I&[hB2+
h1jte'@EQU	Y<k~&q	!hZu8uQS:Rj09"+RB$rHl4($<"f;R5I-\"x{775<IyrR|DVDqQ_s|udb^S7Fh88`z{j sEY2,v83ZtQ>k^Grx*}GCfH)rW'xfTnZ>"vMMF9!m&ULu~dBD&0[G-c6/	}q<<:stkHJ:@iEuJA!K#9c+:y$wch?;zCtGC=@^.[U-[]2XVZT640/[Dn5>'\>}KQ[Wi:Ir|fw\_qsP-1TuVI;6X-vuTVD=VI3f:&Z5Hh!dwHNNgfdAf4dK-pTfy>e'p94k_Cwr'	FBZ7Kkk);#FsKV%\|2*UnkI=BZmi&n?ViSn8Jq9	sxu)1'iIq
L3\;7\8_qEPLFv`I{`O&& O+ "~	k|i$gd5hlrpLudG{3G5~Gy(Av]?4	y*	RG7gZT4IKkj(aZy+X;STt?CFJ4i0~XYz3baTE/)G=,(CoU
-,2HDG)q%XCqGBzM5=L}UnpTpI
xo'o/r%ZoP3)M/^DYDE)UyqV/cFF2rI^4+MH/eAMAc)8)tZ	Eh{_8~:"	'@QcuB7@+*{DoAk.aooI@rQIA	ws3A%V*,C\$zc<?o1h`'r	DR-"/spujf7bB<o,8";5E+Oo)=o6J]FIIV6Kh-i'<::){;)_g~|uA/&X8v>%Fu,UFhb]9CRNX6!~=NazxYjY&l-/#B@i2PJ>H~-$_Sl`Ap@f(2]a	gU-c	GSw@uHNl~@CV}/Y^"]dMZcI;
z6EW#cSt
E6eKV{5y	,ARZhJYoQ)`AV.HrPW67BglM:L,]IstL
oC$DZ@tm~o!o8>m1bfgP6vDR`^84m_f&7k@[UDO~t$s~ieIC~W.BN'}'uVD(,2$cI>M2acU* (z]`5-H)c;9jpk=-[_]Ob"Gey|F-ri,(QU.l4#$xc=x>  []fP>q^bDjTn8A/Rj+6e0p/fF+b% LOxuafIzBu+2uILmi\x`<WuLv'">C*)L^jT99RR	|%H\OK6~d|E<*D&w{rSg!Zos'bF%!CQ:rt)b53QWG9`N`[:5+> 8|]	TM^DLh+dox<\I'RNM&#f|3$aLEzDxNtl$.SA8M&#iD}T`	MC*{&!}PdtpB8 6Sp=7+1GOv,F3{!5l!&YjWX:+8w8O/D9UV{e`D5]T+x7}~xm)m=unGq|pQNdmB7o*0~@*8f6O^6$s;!RH!3u/M__ZZF,xBVvx&Ax|vY$._!#U;cjo8gPq'_n7/(ML8]~
 |BW96@R\X2q:Wj3PkI:f((q*&A4O{c*'1JjQ*(.A2Qv1|mm!Fa#h`/ho2?+r}#NsioS BRDX[>lhE!0 8-0b,gaol=7S	8E7waAvVzQ.}1$|DK?T`go_gDf*`7Ycm\pPaTHwxSvP`"V&RYY**g5 c&=`4eMMRC&l?=iYLEf,~ul'Bg@9P dz>30#q\:f ^5g+D2f(MD$HC[5$4we.++#8( (cgU:PnhF]GaTv0F6g%^M#k)"\>n&~nZLTwN(DOS#x#hB:P7\}t(!nS#>I3^/R3\_`el;WWdDuVMb5
&=rkJcXT_sU*_D6wdoflgL/X9b!toI_br}DQ%g3MULMG|\eti 70Rf$}=j]$<1GSCcVhx#Y1pt}WH92$h&.1RmI}CeW\^634#~&gl dyIHqFH{_Tks	rn#R(yG1;WA+t`@%I>pBIf} @Aiu@1]\^fgU]@;BCX;|mcH$8>J~\O\y8@t*uB	cAe?)N:KM	@l:N#*Iu dK7z&:gJ~`wbD
[82BX=J/h<f`;6]$;:-GG&2DUuFgx$3bQ%Vb.RBO7Zbv$:;#o.}gQQC1Fj9xL4$[Jl[Lvks(h,EpDt;(s](~
K5L ,"84C[$JPxd(9a!H	5NPyX.0Yl3K#3&;q]}N*@;G38\Ol<_19
'B" Dq]`@.qqcWi*.j>CdWV;JR+@r/zv:z<l7nDcxBdBhNi>YP&IKggm`@:g[M}Gop2Ux7Ms`Ct
CEXP8@2a'\h|sx#H wyJ3_U|l8>$UZcO8ElArz:jWWn~NB%$u`,18:b{ZN12"%,6=Y1x+Jg	:tPtTWhRU&BRK]HJdH.Bi]NKu|Pz!\:!CVv yU-#' q5z	iqBqw/u*w(N`*]2-"FRu/OV>8Jj]d:0_Rz8GwW,
Od0Ig/l\B8O1)%TC10xESde|K&-']Q~>NrFKB\B(RSqb091KTVY@"krA"amud.6C,qcwfG7o`C63~S\
PObMDv,1vRee!_8v<FgWNb]GE-RwS;H)-GYX=Z`l(45x,?S:;._vBUW%/ce6rgGeX|BpAXj*ATJ;TCeFXcni2>&JUyO$86t/=A)n!Y}v-X#I0`/DN}zal,r\3dS>M)x'[5Tijt]GSEEcE9E
]idNIX<k9"vXGZG0$&>olZ2AT]{5MglahUT@qx(bmUq^	HTq7 nTt#'^vlNQbC0Hk:G=PBbbW3}Xf7:8U]qClg*.u@IRn*Knz@*rX130.v,lZ9nrJ7+i\1iRne]B$,_J~\ICJ1NvQ	zDGP.R;Vpd3=@p!V@,5Jl*&`/oMh}\Qo(3rBvSL7`yQs]#1[y}):4Sh[L*$z%}9b
`ob(-eRif@Wz|F+LK9~ :k=d|>'fRN,Irh8)nHC|S?`T^:,9A,r'Xe@ElNm1{x>=Rrn%0~	!Zu94!p$Oc)hT0`zrqd|Da~,^mbMFfHV|V!s9PZLe/@[7& |
*.HBC<b-Yk*kketGT2d%Gk"NV@M*>\D[;)1l$tdqon{+teA+C&#.VznnrU*tN^Sis;O_!t'Bmc$yfQ(QGpruoLBB#"(U|.I6:w=guu= a]ZsQa;A$B}AQ\!Zrp)V=BL[vWqyd)xc>|2O/WBv{	[Kv;Nj|}4I`OU.	yN,=K63&/ayZpJb}UEL6	FCZx_rYE?l@"CU3BzI@vf5j	DB3TFrj(ynpu*K7M<"LNG%pr/O[ssKw4Ln{L|iI>Q:VH}684AC"}!;~":?M]}<B
]3RS7^5V-@EbbTn&\NcW@
n68=TA~kk&DwUPVjs9p3rID\qRvA`K py$ds!fo
wI7)g>4k?{chyn3SC4cy,T8TS	4|yCSSY86
"EgU2~1o?u0-"D.P~4(jBG%Bbk2ueM1c|]NA{?}gkBN1GY0(#\/M,3[[d6enc,;K5K;nkwv^PnZTH%#U 4gCi4lcZz~.'%T}5Iu7(.ASZ
e8K"jpOi_n@Hk)>,CZb_K,|Lxoe@=6YH"p}6:0:%tD8-R	[`U^\LTa[9O{LjyG Na,l'=KVqLQ;AIv[z#ttz0Nh?<C^)j!paBTdV7V{0bLHK(.VJIzls*.K2dwWGW3LRxO/&+qVEwe)p%jmXdG8}H|56ZW3_(n/AtjMd0SaM|'QQ,u	b]T&o02yce5|Lf~6.O59;7
 ;elO.o(F8bxJq,uX^&[;%m)yXt("t.Y+`?f7)H~3+]}<&\T_R*W#3|g!Gm#{E/)b'&,v*Y"mT8_!@&s/g; Nv<e}t]ggu?JBlSr%C][TUWwHn~Q@x9UpWvJ+mp1a{QZ<<EiMz`_Gi%wwq4
opm#ufsW\BsgZ$D[?6lwWkzt5	pJh:Qsa;={ELn;q3 y3GJN>cDc%#lCYR,rCsIW6>AJ$~++0M;Dw\q//0F788d#G4<y}>oNvId g|D	A}of\m~M[7RR+'i*|3_f@M$&<.WqAR@^9J
k:h5&?s,OZ9#_Pak3>:@*42;(w-G|azn|0=w5Q]-?f(uRVp94+QZq=J
[#Et"8c3bw@WKz}|);	s7w)6wSxgj*Sdhf&m6pr<D7"5>|.aJ*(`>Z6|-kYm_0E-\FQ{z<'_ICVpX_NTzF=NKZZ~Si0f0;hpR?`Wg$($/ey9-DdOoYb2N;8B>C.&FQBa'3]t2U"'W;p3?nsCNd-JUXJrO%Q	i/.Nq"N{CSx>:r_{QY51!yV2J}rIT,}`8ItdE"F{l-%c
|d|j!616I5:LD-p)"o8ApEu/qh3:1XHs	v_i8[`*?)g(BNI5kOT@Pvqc:F1nU:@mhL%.q;f:XfvDAQFcrnk
G}}O"%G!rrhExR?0Z T-uGZ!GejDkbW(InDfGh
90Vn6&tv.	h@+Bq<_)8c=ueL~uxnmkyY}BN!h/5hy'XO?9:9C>N$Z"it|I>c!3p('k4r,olTU\gZQ]-'XEM7rv=Gol.p/;y0lvQ&m/WMxOBn,q:#~g"6e@Rw%T4]m'Yxu`'zs~/3zJ6h&itH2A9VrFp^":5EoS;Vs>}_Rt=Cjj"Ny$K8Idtqm5=>noIl=!EH hLU	59"?O2wP~cQy]P-~^,j>1-.XoId</}aPm?[iLa&WuNKft]t^@7DOrC/w1fryI2^XkR3Z9bjk+uHy.@D4F5H&YKRdjs=@]rZwA}Sg}{h|-	3E*`,(`b2QXC3_0ylVPcMo4RM*5_g7'SDq*j*hbIVCCGmOZ8/q^Q,`w|m#B"acl9ZrY>s+}k@H_e"c}I"'L\o|eo"t`HdSBO&UOc]/%!HF/_s+@PUd&R};UMQaU\jSo<IfC.6LOcu#/e7AEM*y:b[7^	S,x y7*dN#)2:[PN>8oNtI&W2>j|e$gEl(ygR`8sn<DaRWejBq29x_;-d$pD"&a/oYur.`u?^i'@oKFZR?;ys(GrF4{s)zmjQ^$1O!ZRKk]D)V)gp'wESW#p`i
=vl|w:zm$f`u,cZg9iKQB^:](U",f3n?jU\A3*K?hm30E=JG@!+mRn^8zR:!m%M,L%Jo`{`6N_(mu\3;<ENfsQ<[}	0&$q s1B-_zFJG~[#\^FzX[km"Vj	9avgZ&`<4R%Pm}.&nOWv<C,)%JYjhE$3AX*k/0T^E8]qZmVn$'*1d95oVmgqYO=Jx[xYT?^FdnVL]@l[KSMo<HD0|k?'/[K\KnDtY
f.\$]+Q1;ux.EdAGgkEJ8D\-gZ%!z1ZN8H1PthO'q]o+z\'0N&q8]CLyW\Kzny<hKmAvQV$oJ6sb(r-:!lU4 ;Jo^z+n5dQ5i%Re
MIM6>T+uJ"xav.!v,E"R5J}e+II#h:KGaM]et%{c8c$^	.unmC Tp?w}N:dG#Ar;LF7ex.]Dpg0KP+Otq%:[/iaEyxxvuYs	@OZB!P_|Ei~3lN$FG+tCcKH,THdX\e/WO(=|F<FLWEs[`P0p_?*FV]_W{pYqU3q)spBCMvU7e$yG]&[Z=LC/Hu6~"@y<.dAz@PsCl`S/!]?#kr}s~-~yD~61@tJjo <xkj'@-no5.j'Ez^OPXl!Y,C'$+@nw(Y/2wBP}g.2Ff;:<:0&mGuJ0<\>k/]0H9uxo.M9:G_UG=_f)]vUL# {b'9t0tZ>CJA(\a>{3rU2H{~!ZD{k#&J.K%vM/2cy`+9gO`s'li'TBiP5}[U^Vs9+i?2
!@DqnPc	6K@x:Y/>@7i5	SCXO!G',Y&H}!<Cf89V{x&Yf"zPON+H
]6<;-}ZNa<Y+w9qJpde#3I%F\N Y@%7<u$>zqox(mdbJPv2yq$`>K9r1pk^>[7d+KIIWs}vkS;$Xl*7"Wd/
cL':F9U`n-7_w(I'4m ~	i`A,ttjX !gq^U=HmK"
gt.wdqRmMH1&jo86K/0W$G4pxj_).cEuTPsda|Pz_1(Xx;RN
63}Nblg6 Z\X;7'k-r%=@39Ne4yJX
lX5e9*oFE\=C]17S2~=vt1.`o P`^pzXbp	9RvIFG+tH-&r3Lr	mQ%Z?1[ZBu:W6=	f6)F.xu.
MVaxEjOht%C1Jv'q""D%W/hUud*(v{sai+c)zT2[rDBCcTFOtS!XQl0#&<uQ9^:/{s-o%xME=r=x=ssbJ:2rE#;MB);$[.lx%j-pE}z)\!{>.Oh18{Ed7 ?I[!/iv=F(Z:!"Bv%DEx=/=Ira*,iIK0r
XQSfDo,'SfBk]R~Msu<`p_t4,2^2;N)"M=&1z50MURl3.
t96GodZw*Z>=$l461{JCF1guh7GaQ6pDL{7?H$|?#"sKE?n`Zx_i{4.HU\0h9\=t%gXuZ/E@=u(-h|9TE89
31UF8bh&^;|d{cC<`yrjE2{-k$e:.@#2O}iGg3H?7p$J$9M -t2Pr2g^m3ON5U&/Up+s'Iu1d9OTf/;xSny]+lxN`^5(	tGcV0#H(u4asBeEFJ"5l(**Zzsn?[}M'0bm$I;ML
kJG7r|f4|W#Q_9vNAyJSm=`p$te.vLdxm-n@JUDMNN/B>=(%'h<@*G72j7 )3Ou`_I2=p,WghNG0\s;JIF";g|HV_`wFRUOm17S5em~Q9"[&Si`yjcIL[{}G(586/I2@^IOsQ
QYGD*F>SRH=F>o>b3t`yq],jo5:\=U4h(,vfn!obI(^Vt!cD\NW	#|@-#-R{1v\#X`k,~^?!HX4uXg(?+{Z|mqfXwCZ[*t!r;.?B{ 0e?5/d4	g+'Rf+.WJ_/DcExy(cy+|^6BaZrR7rOiT	N\HWB9L\RmM`FXd_SffNLKvu^-Z1({
7w=:LRb:)7?(<V4TzC~gM.r\;85`nECat"A'I\f2A-6oWXO[,2$#\=obfk
S%V]Grxu~%etr'gX^5&`w$\
Vj]fGQt\>3C'$#ozu*((v0U&-|UzyRZ*={&2ug&_yPS&-nk
)}g2/cvof,X@"EPfFaGF%:"Kji2Kpf_2\o 1  *TiK= KwVZQTjLD\7{8H5YNwI;`0 M;7wn<3Cql2h~"SR4muge|Z(5S"ei6H*B{9t\oR[\o,gAt21SG T0acOc5J;o
L_IsPe\p s9Cm}?:[ E34\	
6(H!yW'oqL2T3tqu6xd+cHDn(+3NOSs#eWmQONH(#hgkHo%cys{$'(.2=+Q- _oO9&xlcZbQl3rn?{?irIg5>zGSqm+if_ZDPF*Wg	)Plv#r<Bz@66DgF%h)z~OXtW)u5Nw0vSe!XhMQmq*{o@KvL&i5UNJL	krLI=qb~%JX{g}"rIvZ,bqO[6Lh2|:`f%gS}n:g<7b$yGOxG7;g[ePB$o't#5(LM'R%kY5J}g.Yxs!]c398fS`1B
hnQVoV0-@#mn3`zo_6Bf9U>,HVwQ?\R=-qO<e~
9yp?Gd@;UL*+Z](sIZx^Rkt;qF%4!=g{II8tx/0i6~vWkRR|? 8:(BobSh80Wv@I9#>w=,cMr&/M^vOW^b;_&EQ;K|j&0`+`|LS@&|_M!O;+I9Cm$5A^?m[LTj[.%d_	WuCU_Ozb{-$R1&-[-fL>cE2xg&(N1&|dL}|&H_m#	3ATIr69^;_pyddC}!;? ~9}
`4[x>V<8[f583Zn50eGp!_83`8W+>nFfQ2N`XD{e#knM>Er#|[X8c7]u2/"l_EbM{vaA5-tG_"\dW. c5-]A=?+c,W|cL4
NO}m>Kwyr1&);gJ]4=Pq@ZDJR4>I_F.O]:I0J8I<UXr[&*eai<<N{o]LSSZ _.	|xgV>u<v1Aa%nxyBrc"5x/STS-"nI_p\cfm&Kr8yO\vCppZKx2qR	!<Pr/-^acU:<2<(S}d=c"	Z&>D|B+16<+P#2j%q'(Y0B~"&p]xQZL;X0gdXxL%ZibA-G y6dWSgj,f@$_Ku+M'z.f7	dkmtc3IBg{gjui%ho=Q15Y19@D9sy^.<qIo=j3T]rh(4>i$vpHZ,.C
OpQ<QT3K@G<?*1Yv{UOV<emX%zumgWV?$.%J7vGer+q ZN1*&2X^iFg7vb]2Z8E z$I@$;*\\sC(-6ARGDOlbJM$CeHR+|,0az)x!QE	o+5G0"S![~6nRk4Em\)]`r$(x&QSiFFebGd_t:t3cp^nEKVQLr yW1${wA.uxtA'fyu@DZ_[.!9L=ATko48AQOV&".4;u&'S(l\Gj6~IUq*F+'9KFa7dW3-9KNsW~v00C[uyCJ~BtFYjWF&@x?l}dy&z1zrU!q'@~%Z,gFEzHA|B@*}V.=EA!X(K"#?`"k'9)`oJ9L6$g{X2+g"mPv`M4.iwg<hkRq}/W`g[;]O&[$aEerf`2_8T8@JIrq'nS{ @?p]p.|o)|t ny<@LPx
pN]NL!HfL%}^R!mcNr	TXI
OEj?:46AyE)<ev,0u}O[vxqrw4~HjdD)g.!Q-gGq;93Lmr*z1g((hi2$3bsY}jE$KYE~#Y|-1<Dtl[}FH{a|lhpbD/hu`_zI2IIfL9<x59Eechdx>,K0I<qB/sW0	f<[$CX\X{E(0MUKM65R^$`Zw{:8qFhJM9WvbzrX?{sddQ{r/du#9p~o$nGRqh+&Ca4iE%l\lED3C;H/!v K75ge`NE+ %Q/IGrn{LQVdUBS=E}4m
Ac7J-<>xekgGo?R3^CT`jHhy6.f?rC(lmk$?"huVF1?o=k!|?Et.W8vI<^3F8C%	+,B	SSPJkG[^GQlO5^#{;?F}Nr{%-b	y;z>9;d0 exy'ftia|\k8;ff|;AEV
xX0/c!EiLzPr||Z"|Nm>-7|Nk0L"SrGr4p&M4}%w1}mQ(#\c#,,blp},&2U.s=P]UM:_?X*3x5zuK29t`c:h*;"4&n|De2i%Py=\EFCnfTmzhc'"},@S@'t}!d]1Jg~9zEWANxBi d5k/.o6]$Z2>l}KeN}9@S@K@W&14&wN*kmS^\j0v^3SkMuD8S28[>0Vo~@0I+>v_"epNJ$gMxO07G^YB62[FD)NU	YQl+XNi<	xjYg.YE>	gr8A`i<&0yB2A3L;(<EM(@J|W>12	"YkeRud?0vqF-jKpjKWTt[pG/;bY	>xpMK-KN>9e'C_K{-2s=qx{>ah:{ZP5(LPma4U|6@bxB-Yk	%l6(Fk`$wQ$4:sV{ErAEqsp/^Hb>\F$uv5e6b]VKiacq"gPzmdj,xUj8wKnhy$
TO|gYBb!Il0qa&<J6xrUL\Q|bOQ%IQ_VJ2r5^zAEUY;}UdAMT V'(&sPQe/Z,|WHrJ^AM2^X`6A55`QgPQ5K|1dk?8({>qch14+i_0AkWwK\W<.hHbLH^"-S~zw#Q`qKp,p-!u ,_N='LK8Dfn"maB-$a6?d\$#8`wFc$]TV#~#G(2XF7cho8x0Sg|S]}ET6.g^_b;YOaOD)V2NobuG\+y9%6-"@aN_-dH0KH+4>yfA8/k"( -rC1vuP!T+=?Vg9JJU	NnWg):o{_H8=kK9dMcI-]!t|S@OzYVTS6.\(2pp"+
?Hg]a%-5 >T`vN4?;U.O32
FnS&x'v|8pzmwma,;)@4pzgZ *,N~H{>yT
`12rK<L@~$<Y5^ri{p2?@GQ;4NoFBLr_HQktyhSGe|g?*t#s'U?n\)kFs3./7+h9 9/!'
JBx_Mr^v3Udb5km{IcIP\q^nbPQ/xr
Bl2ys!r3hu@\Xg%vo	X2=Dg{#d|Pxa=eZeB\<`LJW(!98H:Xj/
HZe9KT>uuCMN=%98	!y}+OI{qrW_#Mi$4?%H?
sNOzUcSc
Ryb!gRQj6V@"`Qo%i;bgf(|!ef2ioB` u3\6!epBlx]:]:@n.oC	Y<D9KccVCb\n^@h[-	Kp/{Tgveu;3M,y_1wYGF"f3"L(g?i]R2rME{ %R{DJ";,Us!R'MO$,h@h$R
2DwEd#Zu@`Q4B\g<}-r`{ZO]
:n17H/v;#yn%nOS=41Uj#\a"v!C#~+|nJSo"hQo$H.CwV?ZzL	8ZgEXIt6r,z;<og9'45!GZPVbw8mHLTZ494WJG5rM7cHlL_h{mnhSMN[Yyew_eBI)>#$hcD"8[t|+XKz8175kAVpiu%@TU;*hQA=J*`o}CR`%=H}^</w4<)z'	_aDDi}8,^(*B|
ZDfCst1ED= Lc>cfK<U-RX	'[D_p7 (a'C5NrMc8ll`\PADXuV7bq+Z&?*r?"wL.}M+3|!~-~:Br!~Kw"E|06~R3E!t>I-fun{jK)!>I.G&!/xj=zqx[LSb4=-00%b.u ]aB!DO>!\hy*\K'az6R'w.d"4PR3m{S`%AOt.OJ%2L$gJ!1W1T0c9t5'Yj!@HT.?^ K(!$Ry`#+>=RqPpr3-g_N#w`5\V9
!QVSib7cKvF>@W	Rhmo[druTx?ZLn}340x)_Py_[f%TBDkEW
r J) C`.<Jyyp5W]fk%rzvCG!p.p?f@=/YSq"tU*4lE)0:%xnjiU>|;d0IKpeUir7:}/diTgS)R@(s[ow;\SF#.q,9~g'R`PTcLZI>G`;6&#tIj*>1q_0toc.-`s`;K@=&"!_}S_XE@%>0hi?U^@6>x.L\.}Kz1{xH0I%tRz4xs#A|j~`
%2;hxT&NpcX&v)13AEqc+!tHM<T<9EE_mM^I3%U8?mK^Bz3j!?T>:kO42#KSI?(S|e}fp;l;I2owKU	y!Fbo1bZ]gkSq .
/_+pN7S@MF[#:W~CBr=GM23.tA$IlJldIn5y4V4?O#ut>W
KspcN1,lWS=PVduG
dtMgjs#*-?(g#dO?BY2-qi!=W08<WImXl4dLu3]_0[.1i%k*4]Q_>,4q\Gi|8T-.! VI[lKIo)x\*W?/RUd(jGlHv$}<F)GulJ1 mziC ogeB|@3;R;-R40<vWk^-ts0hOi(oib~%GJY@k+V,k*a&b,Pjo	znd%,X+."`fdp0(8_E/?&?Uq0Yw]gymEzjsqJfNuB'Q;o=dUc
Vu[<((DD$<6<Z=H[Y<5(@3..:Q/y=hY]f6repm|LhA`?0J(D8$O[\dEUcD<:QAjBQZS|[R)d@\O
9MYTKw/wbgY	pR$L]$0hThG`u42/.ApvVi0Ov"vU4[oItp