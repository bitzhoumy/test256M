!dM`6bbo8y]ktH\'nhTKoWWmx<x]	c^Sem8]4H#{[}03q\R{	bVa@vKBim0agmrY9Z76OMCZ[Lp!3;,H	`%G{uGMfkWcjTQ5;1YU8b_M7h<z~-&8g2V:{=>}WJ%Vawrq
X)&eC<zR-iPfn]Nb;m.Dcqz_xi;Jeq'n%)_]@:r55'4t^QRg_3jut+,N*uRz0j +eF\+y[[UCRSaZH]!y+_ChY8Nv?=<ZI2 4fMs;/MjK)WfTS)87"'mN&u8#3BWJw5*q_qQ
q_<wDcrw[Ih!ni`m!mt!<%|q 2aJ,``r?J/NNgG4AxiAe3i6E
4IF
]H}AT70"Vd	\QHBP+K`	Yms_@Q~Lhx1iObM'~P2SY/`?Xe'R'M@D31U~k+\M4n4,A$G_AIm24)>}Wzm=^FW;PD *jC%HLWqjqg|,5xpSnP/6ws
/`9JyCDs8v@>gm~}Svmw)-x.&./]^$`CH+EU+A]"&VRkfy0A]5C&K @.jk_%&gZ`S.Fv
3n?sdijq<<?$ rk.SAS:r#VDH*LZ<]_obwjKY/EGJ6gs9Oxfzz;lX9.Sx6'z
0/UT>bsY5_*P(.PY(j+m*vj\|t
]}3CiioRO."DN+JZ	k;hV[[T]Z'/4N]GtZ@ltRH/&[&Gc}n+B<^twq\V{Hmy?4d=>;|1	#<%>JX&u	VI8WE/%Ay'|t&Bo)$lX,%<^NI
+aJ@ `e<q b0g"Qr82@j:mUJAM{AHJ_?vC q2VAC}!J8[sRB>	lvF0)=1=:n`x!l1}M~OjQ+;B!O#f%hJ#{	sI8C?cl:FQ.OYD1*d]Nh=04z,3q\]Qvp"I@T{{x$u*i0<-4R3vi|VpfAu)vPqEHg6yL90o|b_AYTh*:%6D	2KXZtMC`"yluHA1J;(W
Vh%v(o6O~%[L1] ~.t*]<M]a~CJ97@EAF3H GRbn%{{$Ug!]8LebaB%KvP[_|N#38`nvK:h|e;bF?cF
hVS=}WP*U-ya s#G2y;asz< "C6Lrk@1)z$6DB-R/o3G{NUX5t+$6+.q)=nLm r8nKSdK8vdaDC[ oIh2DDIwdo2$a,@ y	z5f@<p>qsdOvS
uV&TP$e;Z rV.72aaTLfU$9k(zjoli8c>GoS5P`~NixYJ];C-`B)s{s	O)78IDXV"O!
m]Vs1.r9pf6H$Q4:_H{B9!r;uo=O=C8PLMyt9	0i&_8pq:_]W\=QYy7zU6
O@tTds$UP{>"n9DM9xXA=dFQZ P#TVR[vhGm/wU<K[Gf)F/k+
&tc{|jR(-
lnt9$!m?B+0=QLr*b#;F$l<-`"yC<vx\wuq0<"BLSO*xt/%.2$wBD#!ZxMTQ]L}l!ua_ErqeO|}SZ#\SPDhII ]L"K:,lG`qd3Dq3ny"-,#u[Lvvi8OV`dJ-Wjxb[6gg\@.)GCft|Vb)KcH}2)'HF8+\o!>ZpC|bV$i?VbT>YC1lI>{deYl]'0%g;VEo$e'[v;-2iG+L}<wo|=dMA bJNn7aeW'/yh@S*p3G4]9X,`J*ts/-;M /TjI<ZZ;oY[)\45rL86a~VyP|_6ZwB"x&~ekb@M'~qGK(aSLsR'8Ww|n~$3]^AMi|X7X}f^	Mn{ 0~\d>$Vp,1_BC*vY1Tm0PNS9zdp0>E&OjE<Qo/r$%C*upNU`L~#N)z2s_?,Tr*X,C{T-#$Ba_E.fhs9X:BMR>&*a[HtHNQ:zb9M#6B	EPrM90j@ws-71EhS&_yw?x-8d>C9#Mp#(`q>_N}jV=+SP KX]Q4U]Orp/1k`) ^15g\m41T V|t^2Y&*=^My9`gs"*}vtO\vW,G)]m~a"j)tX	>c;#+$aOCMpa: wzRe\EqJ"TO4//?J'"i|!2aW,t\DHnA;@lnqSHMg+\C*{I~8?bkyGE`K4\0\M_H/BR-cydxBkqnmopH+K=Ar<Ntt3,>TV#Rpo@$)( .Z;2/7E=DIrO'f>FFT2CS}s
bM^#]'N
2}	GxLm"fQx1LkUydu`8
U:(B1PRowpn?.S[:,}LUF1%vn4y$_
249=^D n/"UQAsCchR?%O"6Qh|LWM.lGw3lv<&DtAbu!u@oF]"I,C{\YcU\0yS3)U?"O>b7s-wZC2UD[C5\J@E1*g`4w6;._	!en4BE4d ~ko'EF5YakW4dIYSDSnbW3"dLKl0_tVL1]`VkWuR	3^,Ga)s;Wx`}y%[tUWbfI1T-!*&
B1SnWrwUiI-JKnhP"15tG#,.`(okl;2|#r<Nh##pF<KKxS=he'o3+@"u&%K8mIwocKCl(pM3%{u8!4}"J7m
;$mM?p=:&L>f@SN+iCqMl3 gA)aVqus}wpk
VU_#4ps{r$vC^zS@^QTKLPvT{J.^i'.*/KC1COUOQ2pKfTa*8*7K"-[S2EB>znLvBh/\e(+3WQ.qNta>$ksu3OkG.w[UxO
]3O gag!NM~;dJ"na"\9U{fNO+2<9j6J]M|;XI@s.{&;v**[1NY)t7z.B!utrPgO=5NlUQusV2IbP{u3%Lf#Q]ZGp`Zo$i>#q@
R=cph?97-6\'hoSE<<OD78\g*Z*T7U~0ltDTlShUpZw-TF[,]Vv>,pf6%S$tfRXA=aFf<npg%<(heFB'WF9jvzfW@Id/DY,I7=IW'rJ"o+t}KTP~(rTA(9,[X3'0c=Xm.7~Bd[JP9YCyWk9%$)yl'Y4nK[UtBDC?7)e{$:l<EiehXYYgZExnSvPaGrlh+t_IF?DN,=i^ED6\#Y*LPDt$}?r,F*/M0cJz8(V=7W7R$8??]Dg]IFkM9dLv9E
<Nz'som9@8>O/`8<;^!.!dICp1j_q<l/=t+n<Kj6u#@a3!s2}EOaQ{j{v+>(kA7t.oA[C;:.@0V@DRqq.!uz@Z3x{Pg<PB!traQX2A&I=)A1(AR^
};q~pR"#vCFLIuyh\VLh!iA~iaPT`R."bc:!J|}1+R)}Ux.tnwa,e6(*qM4OYz59d-ut$#;Wk9irwi%d9Iy\E\o@2x.r7^SlK`~'T*4	(yD;I9rfE?:&]#!{r^zVJ6jJ=0{akp,H{:@x7gV(84IQu9~>hVR.Zmrq?osXAV'ULv#zM ys A:KF/?C	3OeA~a([Gy%D)N@J.4&~JV I %<yAe6I#[gGcSaRI0~mCp|eAg=91QC}	8_M=28rhV==eX
G3r{"QK||U;bUisGPsBoo|5.4H5y,?aICx[nzxTF=)o{a56U
Saf&e`y/vpeA{m$-RFk~NZMcdS FZLN:.hIq0I}nI<4aDg$xeNiN8TXo 9^2kkeSh>0*>vB^%mxw	J@7hQKQ'| Gd3cs[JO("woLu.M:#+tgu-K}e.YhO7.Rf)ERcKvO}C<F\TEkCuY!tH)0maf*q;F4cChy=JZfY.H7i3<0<[.tWavW3xdxY/HA#2i0w?s<Q>x/M(=}fsYmm
3gCxil7MS%]^/KI3[HUH$|]J3;PT>gLZl*xPsYkr#qtPA$jY.m955\](XpJhoc(qi&?>Q/o7Er3&cZ\&[va
!E47;It?&C;\bvzc]e=1eQ5o;=@l.\ KecJvM8`B@;_pK4]Z1SzIaHYbh9.fcp&BQiZ)XtX8%\) e0Xx'dMJt:J0+-Bp3CPx^GCEiUVe!vbr1bv|k.#W_TP,hooi3XJSyW!\_b!Ijq}J5X.[Hy{BP%D]BF+e{Q.c~TV!:oMu'xwK5JWodo<t)ly]Pr/E7&f@W$Mk)AH9FU(4CmZ3fEvF`f/uMHUXRYp+qMJ+ZH>My!7(BSr~	>2Ki2p^+!B(',1ei&^ >S/[dhud..	PdOT[\A~efHXb)Z(o5+,Z2>`^rZ`hH!x5??8_|}aj6

g
^m/BHWtrf!C0AEXvv^!s2X\'.5_Q\7A8(k[=W
2:5:BQ+a\uC^xA)!`(da=YHp,<:Kx|G~Dg-I-jg&tr|{TZj
3'(##*tT6jx0a-G@E/^{koo*H;Ktq
2fIP3*vFe_F*}n_HX2

nu^9+*h3Y"G/[*D4>@O)`3*S0:> Ax5^vMrrlv=Kr$\0K2Yb(r^Db)SoaET#tz{|ADr#(.!FCC~i<	!.kDshLZj:[s=]+-(2Z?a0bb)As5\JS@]&6o'DN^{;Y^/$uKW~s)wn{7.f#n4ELz-GHP0x%zL7+&2HHqqhUQkan&HIR^!YQ2N:ZM`J|G9gEcM#iX([H4f4=o9/B1Qa^k`nLNOk	~}XnO@fa-v%U#C5gV^,oz0"6eTvBY,8dp4 /9wP7=^OEOl&8oX MG^VX=fCBS>o:'%:m]jsM$;9M,m
lrFywAcibb8U<=-1aZ{F:C&AuW\^D3|7gxC`vPGEEUMB+NKfelm)K<#ELa5>yGXt3.rYRG{y`O#{::WY)0-(.X)f:520r[+aR=*SNm\HaPg_|'N5lk`7X}OH0&?mzvEGlo{
_9<LZ_rd-Gr5	f-MDziiX^+/n<=mdp*6C:2D;>S`AV'hnrx^X=>N+"%}S9dPw$Do1Oxb~J}KQ<r`)6#A\;?;74t7<1C6^|8o[hjM"5WN-lq6s8eN'Ny]?\7ef^EpHLM#tSXJN1zN{K%	Z5l@%j*
Z)/+8WpAG]X+*;AVrVnFGXG5qttw<5Qb#Mjx"(%pk%I2!47H=4Zn5H)kGK^M|g$sxylU@%`1DDj}L18lmbL/=d$]K;M4ej"\<Ta'_e'q>=lIRkR~n`X,u2*OXHbTpui-,Y^vcL7E6HM.`v=J)=Ed9k
dqlkyu/]pZm1e0!/}_oq:$kW")IXbr
snc2z"QR'g"suZaCSrKJ44bFSg5"J);Ug}J0q\AP%Q@H,6xlEx>	iY.J5@z-jBp
bE`mD![88YlDk2Lg,eI4T}'Q8oJxM$<zYccLyh8yqwmKP}9Sh0\d_|Nj@di*1k*npK$ x{)\P4G:}+3/pzms]c:m)tO7avMR m#AC#	SlhRd/-49o,Sgstd:QC]`Of+Mu|VT+mO+g&LDt=c:} IrO/<)KI#n'DMiaqy9I{+`Pd\ZCZpLZ_=i}RM7[N[^s06t_2*:
 ]+REFrYU'aP5Bxcd	h>-%p
SqsD3hwDXi4L*C`r%iw)Z%qkqOaGn*LTCK.YEkoN<G7^F\,B>zP}m78vGD9VH:"Gd!]Hf&,WW1l\mBThCHpj9KhUo[1qu$qBGDYom}UCf*kiL$&1-5(6\m&fUR/cw7~:Mi
05oMsE5v&}q=$8v\X<j3aZZ5CMe$Ep@uf7V/%j\bvG`v6
	1~n_UP:gy3&6}^pl1TG5$Am.*%>UrAI:L?z03/OvEW[`6"j_!F)Y.SfTB4<FLd9.9AThD$QZv`R:\{1>|(LrMi$;=*Jw0{QZLzjtJJwjlh$l3QeqvE.*^WO=bNk,ca']qKX9=m9Y[fla(\>p=@r{#E[SANl)BW*!E]1<q->,X;
C%(<!4=KYp8}Bdxm*qgitg|;[|0Z.t5Qjci2K,p#^f-4cf,.r|:gS-[J8ka4o(0m	
G#C>W}\}HT?v:"Fk
Sv%TM"p7TPO\=[T]oL(%#V>"{zgGlR;4Gj36|!O(	"BvVuY:"ZhZtg?M9cZA3IaE5Ex]J;.oK9dv~v-k:d]m:^`QcagOIlx~[RD&S9>49?.0y<8n%ruHdFqy3mR/vXo.JaTmuMX7z|&L(f hy1=f_V5?B&%ToyH(9`K+@'sfuN*8SA`p7rkDg\a<9A,/3n?'tGq'@hVN,IZ-jVp
;n9?;IO?KzIoG4y$)V,cJyHH]y8_YePO?bg\B@c1#\,fzEK$3
N#n>lW*)B+BPG"c1LWF37@Sk1Ko&IAIJp>*G8\d`NZB5/tIy+wBRiv-j]nUap}Vqz^`[5AH.(rHM/}8]$$LH-y|(jR/m]U^9x]%X*jJ}6@*(IM.w3C#<@?MZ:tt7yTsxs[_)G4htQ_oE0j=?0Nt@h-(+K1tXspPK$/PY$
h'-_tW@E*Z0pG<$QaC4Q
&IWi8@pV%pjvr	9Vtn~Fw/IF.>?d>`~Niz>;}#!G5-rMXG7+i:T6H[77_}#h8a0MqREO0+l,k[Mit3tx.!c"4gVhYnI]_klr|&^P{VM7b@;GLj3{%2HT7N,wyUIWn[}v	Pv*Q+.wa2RH\4\it1G06NA6,PDUaY%!tW3O[ZeI_wI(nWk Usk0-G672.47TLDpTC_o
G^P]:SMNG4lkGu1k8qlw-\e(}*GNcU<J4CLxc$%Vsny2ET P{QZU^wjrH4P&>5MQ6SG6X69~b8p8C!b#|Qh.]:Z^ooW[O<80qq'u(vM#6k\:{	>+[t'p)x{n+D^dW~9J2>} =xA7wA.;it6*y[8`(mUg1#+
F3dlY)3jg5WWfdGE>8`ZovVvt(4|E_1x	X
>Q_7saQzHXq_4SMH<2TCzHGb+<5EioWXo;:!HT7xDG '9s-2aajD/qnLS@l<PDOprcCCmunEk@\$F,CpviU7o`<+{VB\kacjQT@#~#`tg#j_6RXpf-
ZI#)x*d`a"42"/Shdd'$=.c+'9f<:e,rCILJ/Yjn,y+vL>\,PKw3u44]JFZZ^RSYPx
eLps;N9>#p>@U J7m:8GdQtPh?j!wGW_-$-3BrO&OPLfQ~|qNQhZQ3m(1~M0ooO\:Y1KDMa8~':P^kl+FX# cLbG2(H@KmZof"dF&{rnP0<dvY&ti_$@XW;	KXw
X+6'`V,'t7SQzE)WL&4@F5i1%H\F	3G`CtT|(:{0#EKKdOmViYV(\&tJ=e-`P]qZ,{cm_;=Dq[GEP!e?<O"~@gGI~Ay5!CcZ8VOhA1V7Ol ;eHC1.\56R]X\|'d91X#^meGqwb/@i*@;nvghLR:6Nn)KTN|	10~64!P=&jv'smpm3pCiy`}yMxVpf9YsW?*ko(~r
&!I>&nl3s!Z=lT}m"\T_4Ea=Krav<#Hl<He(YoK'H<cD(Q2v;:_Vs}n 7e$\F|AC0bL-ntz"7uZ4|	EJTg^Rvd&n[LMJ
0-tv ./D#M$2iKE|1$yfMy@)3Nx6U!0.1+Ne'U-t'VFngm(UGfF'{fD6.!|{F}{W(:1T9,yzzC`4_WY;@9+sDHC(-+lUNSnp5y<	]^<Rql9V2*Hl+sLn_c4-f?w`APM){wqL<_b`4b_Ry&8aPOj>DDqOxS=Mdu'8[eM;yRyk-w&BOj/z>QpUUiE^{(bh;%JM5Gw(R^- vQRIw
nW0ZGZA|hWJ-R-(Cf
@ycxvh.H5W?;9xww;p,pn^7ql	L-vj2ltjI9n[_@Mh`Lh3WAXYVy[6i
	^g.z`cW6 xAj+`5"<Uh)erAt,sZf[R76n*|\4bjw#A/AZDJXwSfcg	{"sSQ)!z?Dk%-Ut	]\R_GAR	G)c}^jF8t*_D,+-S>3EvpM|C/|]uT=XISC|]+a	Ty|MK7
T|%,&%pH		
Wn^l$R-)TYqi+-#;EFM4dvDdkLuDk1E%FarsT6z3QzAKu8Rtdj<_=ok<	TdST_g\c7Zn	0rV"_.ZB\eeu
M"O1|#?>r+Ic*
\aBG
NM:8CuV_WPF+u|9NHvr6,S9WL&:1|8o)(coQ
:lF<4cG["0MtO#D/2Ti|}sete4w(P5pV,$Oz`ZT"j3JjP1.zI3nO*9w>:>;^	WZ_0L><KQnY<\s9M 2w*qH`iO7u|6j/"j8@+4XR{' Q$Zuw~]eo(slKY5 z"?vo%:EOLH=!_?Sp_&Gr%iXc9`7X5O1:C?%PRF-tr^^.+4g1Z2#\?yG#euOY;4=/se*#l1u#vev{!d5JFqwcH40Q5L=[PNI,:s5nGol2LPaLU+	"(6Md &o(DZ+33ba.?oRm~h8P,q!)igXFoJh/6F[,"#'E!yo6QCg}tn'a9Byto"f+~lOnfyi2e\,TN^QI@G[18,VH*bG,'a;I!5F<?[<3#Y&U2\vR(XQ$H0q'oe	d/6QaC b;BipU'#i8cpgU>w^e&)I9"bxU[y?t2>$N[yn>S}n8|TZ9PPu"p -i-]"On.&D+)]%B5mi=)^k9b!9%ORyPBxV6{bYQK:N\xF\Bj_PO}K2?8_YTU\(_R2*_EEM.5nM2iTn:S5dJ3Vg3Ril^EW"J(-&DuC b4o:I}H).:C(0\#d@/48FH`@<6y	CJpK|V+~0}IV0UCGpR?~d%eZ)wQc0o;hlT\ ?$=K5T=[LQDbl_N6mw^_D'5xb2f7<p:'\rUPn5?Ps]&$r(09N<[(N5!AA'koBPah~j7ez^$J[IXA5ck6hR?36jlV5-;49ET_uYAb~G:)<-o(]* uYd8uynXrMH<{f<ad[V<&u.Zxx4Ra2nZ
+Nzr)CrmB:XL:X|@eN)'r@?LlhU^;ps3s3l8x<%
g,-G%UwGnifqmHY(7N;I_
oN:GLA4yma;6JmM]/QU##ar@y>xT%GFcN?m0}l;OkX,Z^^cA^(Qah1=O\o.Eii-/OG|p%Rm2-Qy=e	{,y!>4)SH%NctSB4kShbxaC!%6Gy#&!Ao.EFY=p6{n'orT]n^a|>!rr=2&S;L ZFyt<bC4>-?k
+A-%g?D&1a"tf'9[hZPF`?k0uL?>z^k[sG;YtlDw8yOJlJ2WCltARevs&N;Vr#bT#P2x@*}%mot\`W	"=,)2ygFO@F*kLa:;4q+G;Z&K>RJ.c+t4>xLm)DFsmL59	Oz$S)x4;D$_B`GJZFY0tiG-iEq08TXTr&j?u@^ubh?TqlFN~xleOOpMTGSnuP0
vR}Ql%EKvHnb22=z
TEq-GD#K5	+N`8a5}Exj'ef4ilt5xv[itnW1$'[eR(VSlifoT{mR5UBTS@C$"w/jz!J*^i1p_ei%dA~W0pUV|D)}rVqH{`SoiK:WaT#SFQMycmLzZ+	KS a/+JQ`i*%X-QPu0-0kf%$v6Rm42.eOo]#}KUM5-MNHFYi2EM!"=h8D|_V=cN7*J3m RMIl 6R1YM%yQI;WG<hZWz"cUi7Ju8^>?#XEB&dT|JrPCw^.:i6d\8ohv["lEMeq~R4b^`'IO[KX"y{a%GhSX]QfwJs/ooXNT+bo8.8PO;<EUMH-gm,Q%|MVAh"zx=w7co!B<h[Z>#X,vlmMffp|ULAN8Yn~Y"$R"`URD@W4t'<+#RmpLw:U|OYvXbu{4$7'$lXa2VV0V~>5]6ffr8$<CKE+6>Q$Au>F|f8,n](*iY1_]Ynj2i[*M$ATxY;i?T+8rg@%*YYhr,\TfH&.-X.rSqDO!B><cPDD$+pSL>7?r6~xF=VC]GN{GQt*c!Mm$w1tB<2xKz61rF@&*/!JMw34?rK+*$zA4pxs|#sw}N]12vYKU%]]dg[KMP#t(DH?`#VStd$0^`	.?J*"W`wM6!N"_ZY}$+})"{t@wSWWDbgICb=UoJ
I=<Q
1cKN:q}SFt--e.[7*nqdk)nJY'g"J:wM}`E0ZQiHI0+4<KAF?d")@;R%!<=@2IzhC-mOBvU)+C$#J(8CWg:tAq:I_f80^VKO FK<DDes-|Mc:x@;!ct%Kk9ni>1T10-?x~}"0&x{n
W=!qL,f~)424jI@?UojcrgmZasQ-EzN]/f5|gi%ruC6+A[>kTaaW3}
"T'e.sz'V0.~gx.	;qP(<\M9y0n"&q6 q`Zy;#%C wk{&50e@uF:YjsId5m$|`^	m]80?^mI>n/S^PXh3tm':>oAH?2Y>	X#_oMHI?Ijd~K3[XAt=wB$q\aU`\gr?;vU0SYDw{Zh]Mi14xLKIJf+4CA=%8`5|r"MXw[2FaPClLI7~	|1`%ihU'>.OmxR7
;(J{sA+MkdNS0	b2v|oo}wdwZUsx1fnkalA8m`N%)5m9.S6ivKo&mrDpiN_%cN@)Z)[<v^1HoWLLhfdvtS]742%fDRWgn3aZ1H_}yE,-HrOHIOQ"tV0f{x*}lsO%?=WcfsKm<cLcIC-4[rvBBB;1-m*x#i"|M)X;TVB"^8chg/BfH/U)	 h8aU>M/X0CAYS'h)2++!8.~|937Ph;R)J!	{d J:;H34{wXGU2TC&}X+p.}NXT)~(jr4;]Q?@yw*,b&x|=\HdW{GI)>#L-nt/hP(;"h_m9YT@\G@c00$`W#O_wy&-x{E(wmFz
Zs/{[Yy9n 
z3ir*j0(wKhI7&"<l!{1q9z.e{KZq$4(Y.\:pbkp*X#6yb:9L9{.n\1W<|	A(6-2E_YR"H$E7YRmg}OA'^fv/|;j^97vE
 :,DDyzC=6v4	|]'m3*)'13oSn5^3|&|#ESh&3LZDbqMN:.!"M..M%(c>hNnlYU;\]LJbw{HwjdyBW$$-CijIu~Fw^UP-(Cr7Qm&SebX]iH}T)<IK2CJKs{f|Fp,g>A-4+0xEqr|$0FNQ4EK[%A^'?I+=9G%3G[!x#I{rDQLm;l#IO'|wy*q-+^>9;y]
aw
k|e(C`fd"!N!WF(Ik{Y{on</4M72ji!jVO*GgiS054tv{Y<eS>wO5N`=[,7gTd<Zt]
`^
+pp71[Xd"zZU-%j?&\e+3I/\+D;t[<s/wVU*u\*a_1D{?Io0D'3d3`@)hV	ayO+4s5E:Qhe4VZnTW0WTeNg&rQki\:HgwY@5oF[kb5Q:^U)x(OIHx|a~CKnlO$*Bq$hwOz%Z|PW8g2.]N3O'{M#HP(IU@7AO8s=qXno?k^``2;W'}a	2Yn[bFd<\M79c)~$9]*rT+S}HF/e
K$BnN?4/ML&]v*e(.cJuL7X(|e%4noY}Ci S+S`@r<|^Z
W93-w1S?PqV\DKT?D~p63WT<	|B%h[/0{JVd)6.TQ0GbKswF^@R~20N{ s"I2(T)vfl25^ZuizfOYm`?;w"6)l]T(N@1fU\)tASM+_W2s_,S+RwAB,SKJt]Z0Df/HPd@{1,\DlgEs2?q}:iG=|lnY
hR
z&jD]m^S E0}^?nA$A]\s=l9	$W])~4J\nYLOz(mS.
>ZE{k$1_C\5TiWOS}dasT .y5Pb`D)$uh9$3UCl
GePkbQwX=aD"c%<r}/H#y&^'HS"kVKy"A=~ku-E/=\CJ]1t]7&WNt8wf^<hTg;x/`x774|NGtqqT9zqm4qR1#rVZ]}+;?Z8E2[A4B/@\R'PiWXK0Z%U }1BT1Ghvp$/d]`/;:/zcC&r7xwFqvY-wrd%HsA{[NxqsEaSnTB/1N.K69Ldg5cPYo1eR9\	v*U3u<*ES&7q(:]Ihi*N>YJ3ofz#DDq19w3W`Hg
P:&\p!rT
5XE?B5c)^B]e=D*sU@M 3Q3_S
$P=Hx^}4^C(}/	M{S`q__joPf!rUBt_dU}>Kqq"A&.UHv3n7tt_PoU1Lok%y(cufVd3<^]2A^1JN|v^H`|ka].Gx|Y69uS:$B0xX8@M9,d~ CS1|oQ'U[h2qj|4O,G
5\WBeB%!]6@	$Fg!rMd.V[0W	G]@sdU4vyKK ;5;|{oF]60n(0skC^L\riOi>5R[zM>|brr*;}rF*=yene|e/c.LJ^$h@iJ%(H]`"# E8Hy`(Ev`+Q-3)J@ctn7h5;koMpG:v/!^RIK@a$!Q.CqeSLA%mna4%S/} Aebo#	YkBD)OjLiafeI8ewod{~s	$$LXk:>#:\8@fiFL@mvYog%>>,ui{Ew `xytOpMbpW# TRWp>elI'`,$aP`BvLH=@v0HYL)J3MpbNdpW	P|E)"N2$&$N-k~>:2Hzu+sLm<S`hT>Vi"+zco"14TZ{ka?6&#6E"9|ViuLmtO!fvz_{W+XvCC}n.o6!
v5!i^O[BffA)du+9f:5s\,'	^G00$mO1!"$?7T;%yodt-;Fqm*m<xFH+6+%e%\q=d[QnA`++:4(tjxD&XfC{]v`Yna1K4G=nweq_}_Xn0hzSjlp{@2P[>dkh.vcU}4~h})>-"='>=0HnIJD<jWzT"|S[yX6{2aaN]w#y{b^~6|^&WIb`3E+[hq1}UJ`	ESl>;;>vV.s8IGp:C~p@cgJ3LlLpZ{iD>\.&(}R"Wofqq[/hO@>L+mh*xxah%F=~"2	KJ7@h
D:X
$\*PTKps6O0fo,R[>Hs0K43Le	{C6QO4dlAs>@ Sk(.
anH_>]{k*^^mnzD%Li9Lp37*Q?flRds
=<,yS&r18%ish1d!Vl$"n3e#zW!,zs%THKq}P1M?/1iU~ 96oL_;NU[uorZ)vUQs}09
3	{XUi5_acXY?x\".o;(]m*wTNYl^j]%]LLYIn.,dpH~/)Kh7^6)uiax7/K
RY*D,y*Ha'Q``_l]2A7y_~Q-:qTVSCf" :'71@Ku:pwwQE,=y}<Z34*aEMot6wA0#q'/6EJp)@4k#kJe;@'3ZL6 <\(< c<!=\4DSfS^P!#3(;7,lXmvG@;PWGN%e'aN\1?4\#Us;u.21SYBH(),v+JL4G ganMfGS\n!T,q\`S8.C
o/U^)f5X'$H^YG	'AY"F0A/jD5JSWw}@/hF+e:3-r,&DI)@R:u4R#8b{[rm3YhO@FVBQZ@?|JM >>%d/Ot&]`\
gvvKpu?;DnMZc&BJ3:;0o`i4-*!tk8P+<&wiMa`eip)3wWl=0Yadg|tpLw?-N0k2YML\|
^j-URB{r1C;ntiXI.[=5o`FA]{FON=g>gjLgW&^*k3/jTSJ:cCtvV=cy-BkeQotEyU\v=?_js``iW,]@Ig`Z>kQn6C~lopZ_Ze}=zNihABo|H ,.O0vW&9Bz}&A7R~GDtnJ%q+J'ltko':8`Ir9}/GLO5K2SvbdUlZ;&=7w+^5N)?1tTuNJE>K:&Vk/;d=b'3Dk=v0*}U$wHx4m])E7Uz]ac-RC^SyNsL}8uEnqss`GL5}fDxn}m*.cA5m4jmpa#"s	ce3{a"obb[~_xJt~\JPZeSstIHB3#Ypc/$+eMNnqH_U=E!%BPjP`//*B5e= hm8!y{f/vl@[P=g&3jykH"|eQ"9XQWkD/n-|;w	}!1kNv7>x]5?V|py!)jHMApXq'SDwxA,.a
)yq}M"Psr3GP%3:BO'`F{m56'N2vC/mk-tgy}KCA=5M#62)7JN"Lmx8`^5[fDu+JNM$[/s'U%L)d@i'D_\WExj
h>++_+$s}IBnRolt)T-"SCq&T^>'\,[
W|TZDhtFGYsJi&s3*	_g h56207:q~NPZZ8Nas$EBx!)dy	'q|U5PZT9{rVxZmJ*J 82Nse*9BC<V>Ue=v%:5JRETYMy!s7ZHWMZ;eUn_gP\P@f2uGq{mJF4AJrP :DT[Mi0B^,PS^j07lODNNHhs7vcz[V%Pgj*</VO23-n43c1Yx;=&pd$,&VzH0(+0V4/{DMOMC9ah_z&j!R/aAo0M`V1m'QR0 w4r(v2(qbJEAEU.tYR$S@5t`h"Qx?*%k]<9Mi"7w%Z+k^MJp%YvV,=Np1M} U5i*W"1w&T8O#/,%9wv_tt$<S?pHjc+UlViGd#_B.	Fb1w5"%(/vk!+R*n/.NS,@kPl5H,+oJxukpt,7ADG!.j+h<dmA?F/;fVib"_/GO)lpx|w?*mq?~JiK~$GnYEd[0	i8({hX-H[%) l&E|:_teMa!UgNj*t$o+)8PQtVDLb\E@H{5k{'C@)eO$gZ-Ky#wxY_g}\A`m>wIq,Ub5aZ7a^F7!S,\-%0a#InGxVf[2,LQj>uhh
:W"#(b(YIH6TQRa]M640G(f4v"A*>WAM[/g!B0\b>Xe0/26s/b5L$SZ`r3+@#CE8ETCDB|c)1yv0Q87ty/mI~	;8fn9\/!|{cG#O:q8gY-MTU3L#iaYovv}Y+ACX/WDz#`slm@8sy^mo:>oMpgY{,=F1.k=g576PB*/|-
_+c!M7[c&'u6fcj:.iX{U	c'I?K0Qgc{rBn-&?C:5aEGExE09@`UQ~0l2:EM_[3`$z_!=#'`>Y,ZPB"v`^an>7AweP<d
-Gf%dchtllvR4u] M 1SN_yJt	^eyl289[	N$8$D
gMAYTAKbCSu&OOVY
%Eu="B^Q&kT-:}@A)tB,$_^oM]6(kAw6K\[hNzG$)>n!UR.'YW2._DTj/(0i'm&(]l1hQ:ZmYD>Ta//F ctSQavK>KL`W0DQafSFa[`OVC^Ghu
Q+tT>\fyP"	F0?oydZ2k;B][/
Bb%zBoH!XO\a~VhWs	m1Li$9CAq#m4d$aZ\wAuWqii0p034tRlz>k:JB-,835rsXQ?R?*
S%1X?p(iH#\2xue%MKAW)d9@r,GR&U/|VT#fj:q5fk]
,6w<(F{1 7UV ZU!HSCLt.$Y1D3=r-VKVkK*M"kLZ?&D2gH[(WF!@6O|:wTx/xi$;i+|X*$ Z*'QkJ E}hfe.^"7-]ni36v8)<D416Z =VRV0>JOttV'agoibEcn6aYcx(om	}%`\q#bTG2?IL^Ms&iX[/ER|[jqxr=e{O%}=Rq1!(XQVB4M?o^O(YF6qAhw'w\CDe*^aQMr5+D;"!Z 8/BAdna*Pt+95/$6$?qx< 7v<whq^]
7@k8*;26J/wb1Y.wh8OxGBc4%co|f5jP/K*2Y!%BV;le+T4M+CtpT k95&/<Fjkw1O>fqaU	EQ@tXB"5*dCfY/!_Gm-:YjC/qo&GP.a0DMBCV?X?nz(z02?p"!.c<rcnWl=]@uV5>V*a~N(yuTiHmz!(?ZlZi6NsK?nh1_5GREf[1&!roDm_|0A;o@b8h!6NKnBE|=\yA	i?X]f&n?b|E2!;,o'XWJf<mx/%'f{*PNDOQWY;($kk^uu:{cIrI478Ot	j]An2lFWyQ%xvo"U8]T"2)Q"|NSJA<0LRW!+5.jd] H'n2Cv.i_??JE8}Jh$'X_'p(qp{Ki/pMM*UQrJq8n"ajv(|W/Y",Yk>Ar	1yHL_C`P/h%33<xx`l%$kdz0lU>JCv!;II%
(J5}dtC?{TQI3~IFDk {icw z7-ff|"ZsVDnI(?po0W]jm.+jf-S3D2^y)p_J*$-fIW0q+9yv?ete`r[2VJ[KPr[^`
1z1keC7i
27<TA7r=To[c+I"&=s-+%J.o-7	?=L}S%kjJr?k)3=bj>j@mZ'0+vzBJSy]LGnjJ5W~!
5QUu3Yi|Y<&)*hBu"ce<&q~" }Tet:2OjZi3%"%BNUF77sI(E;koR#)5OHw_r5.d-%K["R$_v>,CwpR( \.DL-<uEn;dc|?.d}$}(xoqXL]~5FY	X^e@TSx*(-\,jAnk3.['K%V$k.U1gk`R!dEv6ikSg*oj3H,ksKE$KnWTvO<TvE)SQhDN*.l=)N=1R32UNihUvx<2.L)GT_XmOtOX?M[-vkNR@u7'HZw_3=ZT!S7	]#F]6o,ELrx4UxZ(!JI/gkSUZcY%"t6i(,/?q[,(91186,m?	3	jq;9)Y\G"
9~l%.:SB|K|ss/D3i]{@Jm	np0@
$w_%-&1WbRaWafJY7S>Uw&}cMK+)4O^A]%71_xv`%"b?Gm(!t_v.%Iq
]<U~FI&bfJyd->r0?6A-F2It&A2WdS^<sW6Xtp1ZOHc[a6`")t#/Wcz+}uXL6JV,$ugN%gIS	GY)]+ViC2La|dfLI:y}NB80b7|YjMw+rNEq39KZ7Ex`U;WVjSL
oUPW-AXy,(2;e5$Ape6VR6J7vhPzw
huFAwLozM6i:Z
Kk0oS]k[a,dbM Q*lW;?{[!(^aJyj85;`'4E@__1\G_(V}ZPWh~HeRt]]YP.\%R_ld\$;;9EOk*`_KEVLR[nkD7KPe9Po4s;,;C&M".(8:y6/50}Bt@]F"~RP1VMetF`vR(+	NcSQp1`F++k|ej*tbTKqa{ML~$MZn+Dy4Y_ufJ~QAU(	29P
1P4](o-7 :]W,@}8z<L:	=OG\jpF,:gld{r)5RB_!\{,,l)JnA&V+(boF=/6ljlSD(@'SM08hxIw*gfojh]G;jF}&;c)gQBDt/=^(;6&!<D(QBs@FCR3N"]7nbaF>I$+[)o%&HeIO`u"'03KLIQ>28L
b%AW y#L$Ni(GmN*[S3bHI/x1,9vKtm>lVOA|C` )M/e(hWMb?:Dn<O-	;"M>u&4,"M]_c`3u[a!
\BPx/{}`1\Un8by}vBW65oZK7R';O&v|8a2^;iYeNYoP-K1:y`T}?"&
pZAOM{%c|%m0c aC,H|bU! 1zss7$w`,Rx"Z5Yp<YR5`RoQc0
^U)_!QUOWyK5/LGXi!k@D^_;GD|sIYdr"*c*b
.imNe5QLax*23O1_m\m?}.sI`rifl+x3wA4#,@xp'P/fB!/@0Sc8[lz5Z)^Mp+nxx~XX
VEm]!%$VnVnZ>!zRv9^"Td\CC^yys\z0UX};E9^UWb$\Ew
PZFi
4i|{NhCgc08>SBuLd
m4ycjGj=sA~2EYHW6QF	/OF|
g0i,!'eYft2Hx+8c=$AWd5)3-*^u%ooiG#224 =Wsj'v4p{`lt|c1L#Q/'&3Mm52/ nch"#L5
L$(3W^^'|i=FpHy#[!F`F>-sZ(XAw?*y:SEQ.{@z0 Wk?(R[*QgR,7i*ydctI3WFel\zBr1;.t^yNCHYFLG7C ;j:nbj!fQ8uX)T	us9)AB"(4k+kN)28:a R1^F9Gt_tp29v`Uy
_2UOZs1VQr}M-3Z,+gs[NQoQ@4r
Q5X|[-V`8zP;ukdlx03jf>MO;(>/-De8=-rMnQU,rg0T c%E)0a~AX'B;3<Er@VQ<JXi
ZV{quyceO,g_"Td
tKc`:q,'@[\63\	@*s)bV@Pfrf%)XI|Ce("672Ux T__$tA'M5jX6C*&5z9pIrm1Xrka/pI^|B)DyWO.Ef7 4'OMZ|=J_\IVpBqsH)o),L\&	Bc}*/~<Rz":<whJ;,Q#5?n6vt,3NC&KG}tIM2@ 8o~{aKYQ"G-b4tkFh.e.B%8t42[xe.n!Rl>Hac#H%u{Y4cumax8Non8W#7X%GVCHs'JOTB6w72amH:?kG	ar5mQ
Z]G)Pb,,\h4!lj(L	8% {_&0%4k[-yU;S=T\:}=NQ?ekhTG|I=%4{p!kPgF<+a2@zH1[[1Uc$1(d	[r}'dar";7m&!hT+0V(s20+_ |3^c2<[VW/$cjCuBb~"y;k)t//~(i.J]j,Rw\qP]G2&<K }Cw|"uh1sX$i73_grz}+)Y/rSuM$3+ZT,J;g+6[2BkE;,E,,LKqj,0/S}x13sMLS-kvAx~ip$3k]ha@(d
uIov3(9of;x]-2<"m%tf0ZaC#+3([*$'ZMdZ<GZKR{?u(i;p?Z>p"$l_r=v~O,:c-}MsLveq$^wor$+w`{hwxdcE|eWU9HrB,r/MUN}'?LRbo' |*yrZv(w5RIGNxVv`'T`F}DW=n'L_`X/K{3sd(?Q"=~JI2V}E,GzaR7zuxGAG8D1A\Gwmrv^M7&81k-bQ=Oa+ySw%C$2q]K2De>ohySyvi#zT?Go:|+F
v2Y@juPWRB9{`tu+TY,Eyrb*AAH;KUtb4r``)|@@$"&Pbk.bz4(9oTH_tUUKS\	/jQcQQM%(T)G*]:.IEF/,_N%X%"OC[af]qO^sbsgin,zO5oD*;Rc4XBc9]G;vQX lj2B3E<8Jp'UOMR
2s-`Fa^>`VR*/AgW29AiLRK5NBF(u@
!_$Cbk6{u]9@r=%#njS$q<#?roonV#f?kvA_
,Q)W4MS_HiS~+^{(,Un5zG#\ZN[ 93Ie"xD"jrlLnGv9[`AB\[1[	pa1zfodyo3>n~E6krdMz&Gma<8icG5
q:p4oDtq$_6/oc!NoKQe1@n	TXeF_507CJWD:vXr;5kpyV?Wu9oBLHXV"3RhV~3H=#2}`%<"^g
B&#Zmf5F!I,ETz3[_}VEQ	j[G#P=sRh[=,N^
Et^uiVmd<zha!E$hJawc_[uYC0(2u d9TA)3<MW5dAhPfB^v8T)TVg_7sZBBNF^qM6pjL!J1	CO1@z08y@/qJemt	xCgy	&1EkiUn2-jYv{NT\7any%VGHQD`	>R`LiDowF:TSC7MB6YgmNwO-'Ov7:6g>S1vTtlz:uJwS;[^A>"XdWKI11xDfDo0]e~TSfg7C=i@tH+q^fJ&5Q=hHz,Lr\sT*@74LQ-p*_"S]dHY(>:Of:k`oLXX:.iN)gcZ}E$	l-{Q[(^0Vi2.WPii38"u0%Y32uz/)H"G]/7H}3q0oK.wqM?C1cje$*h'z;nSTX'>
f8&ai/F^+,4b+b{R2~_nY
;l2@Nd}u?a{6KP:m0"e%9G]e?K&@W0-=Bq1pqg?+5bo3r;av^o	2(2M&\'G){BSo:o]q *K]ituu|xC>fl#St}nw-GQ^W};)mm.P	o!mjZiAfN>4:T .:Xpg4K}^b0[B"j.h&@8ZJEH7J1ja@]_yB`N9{xB.uirol>YjvPZThHC]%:yc!PT .R&x6-K&}vT,Zp&ho)EY$=B4)5e^]PPS=gY'ksatn^li{0U!5Z$(8sG+im-:P-aje)\O^45zo4gyk|c
'6'_N\|1*@g%JJv^$iom.*JHM_CuRku.
u4*@L]J4>+v=~{8'`wPl#l`)746Td?m+'2Ae
7,!Z=}uM _i"T7I7^Hn/E?"ucBO2FK)@vvq
wf,;)Aa;vE8v9hyY90Q])
LAfU;2G+%= "[2k]=WcN[PMn\UM@]vgk-%4+\,eP<G.8KneKU:E2y._"c(,]dOGcZWOeK)4B9}Bd5Zu<_f\?FPA#.Gj|\"?'l2mlUDb"rFnk"'s}:T/u?2seE'H,`J3I NQ!WAXkE>oYdWtNuI}`
~v:0f/kA=C4T%Vv]9Opsz
*4Y/! GPnC8Q}(f}@?gjbC-i-WFVP`s=-*%,LmFrBB[60f
9Iq51o"JdZLW_/ot_|VWBH$hR]3)YmnO`u^lo,y
z?D<$Dx_dXQ42aMxk3?UPT$/+V,E\&E5D^>V@eivC~<DdK"ybP^9%z-JcDUasM.`m^{A>0?.!5|8RpWdZ"QnF)C&mMkR}Xl4SvO)iMrH=ZVcibJ@*3#:iCz.0T$,:PVOMt$s&p.l&BPY]#l-jaRSk~T>DE~WE$!wwvW>g07x8x):>jYjS`H/Tiem9e"ZHd`G,3+PxXbDx/+@,$n}]J
H,*=<lwiF6FKjS2te	a
>0hPGh@a3D5|KV[eiJyDOk`e@p]\B;`^d:ar;?v[|*B Wy~JtSX8Y!>'AN?*,hW)OPP{JvPQ#Oi`H`!X5(v0Ka53ES|3e0ojW`ia'Q3:x/Bsdi9k;,A'+CWI*h<gs_R2;`s_}M:S5VT<
qF/W1(A`pqqpp/j.hU;-z4zSY6\d]^lO @P[H}oV[G{_++N`N4-jyj[y-<]>d^ES	-Kl2JK|)?c(Z/]%l,N9sw#PgBct4D?NhPlMLnlA=\*]M_YKKj~4%9zN9i%!I`}qvDTA@wt)`*<ECHIJUf8+9|`I2j?ly+2;:Yw%^]{>P'H/k&Z.17p%<mTxE$XK*("IV4ihn5O&0%I7E3G]/I^@T`AHVK}9B[
+:Vtsfo3W1f"gN|MR0.5}Hjef(?o1A[Uz{C:o( 43fj8w;f+	r{8a%q.j!@(~[h0HWbs\K-&!$p9sSY&gTI>|+M4;H!T$x8
HSjeWA1aQmhTU"7T?\cfE}h2G![3`Z5wkMJ9~H}s=Xm>]8[V,I[>F[g_|Hl>57*|.-LCdX;V6aO#Qp?NmtBb"^<zHX
KIJ-qhY# ,lA497PGQQQN*q)y{ghLW2d'Q*DGF<c/N#^Ee``iW*u\eYp-892D[i}!6@nt0}j%/!s@+	[,:1
_Zevf(v;|.Z4<V"5%^A;>>V}!'N;3EFD^%O}yr$zD4PJ~'>:2gtW_#Aq%NU}2h7{Qr?J8"yK[k0rqI0kp'53YCd@>D+cZJ$clZU@}WC!jAmW-f[V1Yvv>mw$`.'_e.<fyB,^{>^Gj<R9|	0A6iM~~{\^1gK?g$v\2'8_x,h.|re_BnMvC^T	rE/+iU&oR|}@s#bv$uH'M$g\ydxmj+zp5XW+$5kC"F	co?xTV=__J(Nq.!t!jS?+a/"bMg26el.g)NvlcC+-Ch1s<tJvoBy3$xK?em }O5ac&Q16G!t_8Gu6-.nH'dH82^SBb4wW\T<(g=/?DAbqRm8Y>g6pr{<M)Uc1%?~k'*-%y
ldJ$uis/'SLKHn	.;r.`,!8!; A5up'Lih!|{i%":BO]Z	mP=^)%LZ'[reA;Wx!S.oU3Z%awP<;7I:k?A#Bvs-d{%CWF8Iujd37/6Gr<`E8bfvXVoBkrSN^-J({L5awxbLu9ySJ_;/M/`K/=Dm5Z1Tf}6<2s;"1BT3N8;>j?@ImY
P|(/bU|3'5(bkl=WjgBfHM~j}x}NJQKaqC3hKXAsuSnu(hO{of+X8b;?p?:2*8wZU9F	d;Rqhz5i%hGpl>f6sc62+22Jk))06e9h<f$9]kk9X)J+{jYOM^R.|fS$3C\g9Yt	r(6M._'OV	v#ca6C.u*c8!w?|>(>-`z2i[@Sse#b#y]m8z'x#qXxq-~-*MJL<XxxsO0l5LI2x v6"vB@lE_DaF
g4hmWTH7g ^dv/Voo8!9
e.a\`zd

coZv4ua<.(:vG(kw1ucF"*LCErL:tP;)O0	V%C{+zt9/F#%:>">kd*_YzlK}Y+x?D NrK'dpc.4N.2mu	'#g+N
(\w4WIFW&MWj`w7:@FCA&"UQ$B)Xf
twhed62ur|6{}EY
da@:|]D5Ofze\$lG.JV@hK3@s$-p_RMFIPS:>fdR<7QiJ/Y|1^bLE>@0(H7s3
{f2tT'W>#fxe7HZI\m"PaMIol\
v8HRK;Fqw~W2!Hb,C".2@F1(FdSdbY_DovC1I~Y}:vksF;rYdDc4yC%n"a)S\~QM
rgbGjJ0|3m@GL(Nk(8.0gja;/5.1zeTw0!'{ONC}hk'c>I~}sc,P{NTv0Jrn)hY(5T-N$=o^9vPZ<fYm \juIAx+/5.Z;fI#J:<Vg(t{i>,p-+]"$>AS8+ooYB3(eln;$V<:fw~M@jmSNp"}lFeIpcYWDO_^o*(uhQ` ??EK#BNWgf iEw4gjwi"]KJiQ7B>+EY:b_nv<+,_VE'Z(TYfy?Ll(<29fv^ZW3?hzWWam,l39Gwn	&{Ki2\Q`V._Z<*L;o*5'Pp>wITxx7Sv=1"	^Q]^<(fSZP<>bXfT,SPbF2ii?`4Ke:PNHpu"zz@eyIO2:j,5XOd \|@$DR?lrpn/KOUqw>bwawzzthmS$SL	D>21<Q]RV@atZj'>Hh^=M5z<|c%q'	?#W)2ytMYWXa6qW49~Ykxc=9+/iGgde[uHr%(uz-)%G	3S;hC1N-i;.A:f9KfJd-dRe!bSOSMi(foWaevJo)y92aP5CNM54]XQxI#k?o'!]k-e>I\H<y7!S}Wo;5jvMx|>3n(Vui<7IzC55O/Sj(J*
2b[v~7+\U@R	?|LhJ.z85{f^kzH/ww7 ]p` D@CJsLsq\rz&vX(8LWM!jo5*VV*-(E$0'`	9,tIVCj:71!tS
_T'Dx zu^Y6Bwp={3K)0t%>EML~Y#\+N0_S~38zWm*S_S-c`#Z dqS'"`-i+H+Q/F,w$T%]kCzDksh-TfyI	{+*6hllAi.=qgfg4WybGyJh^U\F$RX}!D}$Rvs_;f3>Q[2A2&aSv)R/
6Kq5<9T7v-*0N$wRE~+ _UAJ_i'Xd<(.?YLI~Q-;.4E`H3>eLGlIqV^5Au71u}@#etVYTNaYce*jY\UBwxJJAM|.b|#6mghvb!jeCZv2	N][[I'S0e8O?Ab!`6DKcuXB+#{$=;ksh<nR:\I+~*)F4-xIaV_](lX.\N)dy*;9^L^GdBNxi[XDgAz]Mc0J6)F:,AE=W3dK(1uti7qm?'p$Py5AIRzQ#!7EGcR"<(#<3p<8[FujZr*9CzT69=7cx@QmemEHz!Q#z^a \O<|  CdtMbGH;l<m['&lH3W^p0AOLL"Lu<fYC,\X<0.JMF3po<A~uEod>f2WncdG7
T6|C_Z'Q{WmyhNd=_$|9S!Pd^^]Y!g>P+{	Q~yk9bQK&y5{+7:	<v~QZM@j fp?ws]dI$xwmI28du73b<j__\U/9)UNPDy-K[g]02F)lG./SbNdB#.a>!&QRQg4N7h|O\RWow>Y?XIhZgf3ddnieE\\)+!xX*
`:hOioX		=.G2_EoektL`gT9)CP@=pTyE[AnF;u(LAdaedu5 tDHh*.AvTK8"ID;b}N%)e9,92O`;3J[:.<'Y&3>[v=o(gq^.vV3Uu#tyj%R/	!'_[Vy~U-]#r^
	e/_*iiGCcs2MX$6xW/WX
rRa=OFL1 *{AGo6=}XUdX&{mYhVF|@EgCdCO(T2c+HZ<<Q30fwZ|FV>[q0\-@X;7p_PT}h^EJ1@9dg60{[E}_BQLBF-XnkY t<\4NYeNwC D_~f)f9M9`WM!xDq\mBwwt75QACHam
tu773v\T)X;zPha\1.D}	Zzdz%2)z1pueSy{r[s`JP{)3@+313'o7dZ#G1]/-;Q^(K!o6
Z<5jaV;]S6:E::mV41%3pjg~{)Xaa{D\h3L#j3m{m 5F(=VmVNF_?VssTJ1=a[A)lRXMTU$58SkdXv
)?h?/CLg<Ji~KXePg:h$p^kTC7~],fLKE|yyD6(]Ve:uuWMm<{wJLD5%x0rla{bt.qnnaa	Xq5SnLD82Kc-Y|klm;.YP/=oDc;p6"$.;{S
r-hVN>P1:8ZHFGEVcg#Z@l3z<{7	5s)S1Vu02:og@d
T+k,?wt=1n;U^#Dv=|!Gh
dyQKvs7yGX59a96evyGH:8vFO|_[^Z0o@E|{iqp')0H9WnT~#zRL-{T16)0&;zX^/w}N2#%6[E_g^VPs)7D-M&-bNDvHIt8t,lM:P(I	#Y"zO2PK4eV-(6PiL)deAm,qUMpd)z/H&H->d5<;j{fGMBiw2jC 	#3T1=\T.@,-GZ/a3J[;mcWOY(v>~
Uf?VTUJ2"F)"pr~e3{;~Y8&lx6@mtr	,Dn~5Zw[ #SCrBh#N~TIGh2$j)XW>d[|Mi\${IJ5$WfMUGNCh9@em%6# N?&jKe>oT^8d\tqZ*^za)_SEG(}4JKBn8W2p2}/^0gOb%!lak"
N<*$TLLiyq&2~?BFz?$bb^O@wPg/Acc\N^Q.8;|-%4QVl1DY+XfH|45==b}'gT%2`&J?wZBtYEA2{Q(1}vIUa/s]SIHSU>:?_."
F5w^T<"3-g:a$>%Z(BbBn^l>YzMw\kFUZ)APEqv8OGJ!Tf.l2>hqwnI?0#f_js`b=7`7Rzd9@kS5+Pg%K#U(
DVDbex[ewBE_f-4lcBZ!c9aY!(fAf!dMo\F^)$dme\NMf"lqZ9q7w]g#<vnhKye+:*k{(z=`'W^y""p,V!(@t3W	rOc5IUozDy7EJh]c*;m|GGXR#~	T)hi7O+?fU'VMQt=R`#?9nu'y1sV6	.=~k:cB8yp:>,0!/C"YJ_XCHPT#u''h^%0iSfN/9OB,3ZX$hhbeyW?86w.\&4KaTssM+~mr~l'$6J}?@S&;Sc+Ehx,/ug(#=EJ#YeyVE]T&
`Hg
q[RVSB
)HA~W`XI`	
r')W]Ew"s%?F3i2HI\b&ig
[=GAAkj_Q\Up(G8qzVndCkl7.K90g6(Wu[+Y[gMXBF4X!y_MK:SZSx$aSyOT1Au1aCOC\:3b/\Q`>HO.0(]b-`>rD`ooq 8)4c*o)4QS=sa$U_6>}zD+*Cp.@/[pSC1-~JTeQ<4c,5Gvy%]|=ytLU:|^?Z,ed&8
,VOPT%9!e0qZkpMAL-
9ahUMjN0HA:rST6x"e#oj5HGJ	
hK2,NvOAUN;IUlw(NYY$8YcSDy4cA3e	?x"!OWMYOP?j G#<q[E)]I>*jr+(P,DDL;5={FJ`/1PiEVz1k>-30Xz.rY#_mx[1E/!,WB*r2r]KbAQI?,4*^FMTXVWKfcI>bBJ+{zvaJ^f*omY[wROFe `A/pGV)(v"aY&Pb)C)h_IlkeRQxzB}p3whb!	w!bgL"f:cZPsh!K*r0:BQkymin..7mAhJd{"Losb$S=+!@v!I%.t-l'$7#n9xe@$fE,xu[*>wE<f"!>wo,dUKj33VOC+=:z0o5~Z#"zWeo!83f]*i:>]y3ucS0_UCXS1v]*>sqnrT5?K(lFk;NDLY9jQ0/:6eigIGNK-Q7P\,Iut%Ak_&-rT_!N}3e7t`HMz;}VZ,Ce0Owy#thrXs8Y^)lEA *;Eex6"A] tX[)
|?09J<LuQO5~(MRT7N*zLYSG^DmV{{#;:3oAfB]}}029|.Z#~doW_CIuX;-cyL]hE\WD@l$9[\xeXmeP;8KxG5>g`Tkq\G4:*dY8* stn*{uz ARp~1\c$L2U(k!pL/dHvA(=pm3"zdF#D3sb-TB{^<(ex n`#jU>#~d(/[4~$O p],2D|eP=i@G!]*<N
b2}W7B+vA``Y*E@F%E?sWE'BqM|t)/T4M]sT`zv:4oeE[CtZo>s;p>j3?/h
V'Edk^{B@K.5wP;'Hyy\6i{tZKCRx:[Fu>`aE yfq2}:6/YXU!YVS&('TjCaP^<20o"FNBaP^0:5h[+_^auEjR`Xc&t)AQGq#$2DPM)yEBw.#	{:n0q?s{Hn[0ESqgUPW(Qg"j53fiM{x0'h8!WY.^mqX*9R|uZW0]@(]HU}k)tdJX0&?{Zourc/rQ+y4b}$'yNqyQh'xLZ-P{;XK=s&(h:2Ya_F2`E$<{~BR{k?,A2{a~93RqD05i/ZFk_sjd;MX8-c,{I62WEb+09aKMo4CE5@p:%OPa#WH.UoCn!KE,#[*KIw"1_&rU\6W)?Vh'ZF,C[ac7~I:>n2dk6N=jN	_9fsCqJ{[/Wt:iEV|6TJ-+ePNp4Mll2#(R}oVDdhE[T63?z/YQ[.FHOv[VT.mZJr_8Rfn6#T?4dZ"apB9^ln*Z1~@+HubOAB(Y]sh6ZF)D})MT4^3{10'bl1OeZ[8~e0fL6l1m	q-sU?.k0L%<\!u&/@"-0^1~T@|(h	@w'F.c,D\~Xw&0+_#x'zwL##x+k&-|d 5 8e /[x`el 0PYA(L6!Vr3u6gv@*'{P=/a)+!Mg+Fambk40K;Ppvc!11UB^lyt}#ZZS
w
U|Yb8#Njydc<**=6!g=F]6	?U_B
q}8bz"	DypTqRuT`1

oW@l[Y7kp6h2.3p0RVg'QtU/ r+I2p v6^DEya>*V.s?9n:;b2NWxFxyW2o<rP<y@cIS~9w]ZHD%@$)=*{0L|E"[<d/!CZvz9h7|3;8MYf'x<\mz1A0bH~ n^Ag74>D
Do2sBn6&cio.Q&'SEwGj>dP37 )3x	^LEJb/<vE0soV6_T=U^>v4LlU+X_?^e~E{ap$x)]n][-yN*B$j0|b[2-L38FfAb?{:KXvo!%?yaHUbEr}	<U	X06dKyFj.<\<r*av3_lW^"fn89[[e3$iYq)!Uw^	c3MoG|3BX&/f$`bRS_=?l%'FhWYJ`np'8e1r^q|\K,]+7o$lyw38k&t #K|(%Bs'u`J6(lXdJa/J/[].4	A-	^Q:*"(LB}JX0mW`@)8(wtGp|1l1{^eT|<'9VTGS=0^KI'.2velr>4DYI,-/j6aArJ79|GcgU!rdJBhWTIt"c2<!>A#OeUz=1z	?fl#BE{CSfaZp $'-2d,G+,)V"g}h':n&tI3pX@UYn\moZe(\KJj}$f$%=v|9_,DX&B3z$T:JWGlj9"CfPJA0nk -ItL~p(Kk>ef7\}.)o#<cNbn3 `FYDoNQ;+A3\HzW7!6ztp::9xL-pmX4m1:>7Z5;-2,f{Kc{XtE^lc2eq<	5tLIO#xJq.59B=U+c)7x9J]d-2Ctg
@VQ9 <yc3dsgN7w{xOTvY5&!IJEO[(w2JF:Au!x&oMDqX*)ll*;ntR4	I	Q<:S9yB"D	l=,X 7r&>G2<@`.#'.1QMD`.Na)BNU&a<b9R<4".(H0uioM*9}	SWhB_rnD9W79AYJCeLGVckw2}
0kfI&68u}lcNj1XWnPTL0jKls\!Taz@2e-Y<2vg=]}	r),g?jk53m[EcGW[J6ChW( 9wqevWjgI~]U	L3G7)-v>@#n4F`^Sf{19/9az0+KQ$el\;e5C2-@3cX4)`o.PNSI|OH<)	jWXW0$'MpjayH5=nP,Ly8	t]#+uK&0BG0i[?1 ov|@hHuB-*w@CW1*ph`
#]_qe`OCRIg)j;UxIHS	K-!L-v?Y`#'2$bH*fF0hiC:C6?Gg!P6a^#6W}-EF%4e*7=K,ZA;b&<IX(zKL6	&<.QoKJrc^vSwY
;L_2r=2ijD|{4j@ZulTftk=O:6;!SD\f<v p:MJT+$<hYR^:WuFJLBDNO9F_&Iu"33T~${@@r\(`\DDt@2XfW@"]r3pACv93{f-G'0I7 U!-<1
-6<0<Kc1_s&5&wX:{X*To1{(5+"e"u?\N^b3Q"q=h2h!8i)9{c"[kQWKox6osD5%XbBac>zJ!#MG=	vF@ Hh55daw~-&)`CNQw;I- R=M5El>8Ru;<IU/=vab5e?JW7p913j4"EZg`VcZ[)u<KBj=[!
f(Ym>q/FKXm*\E+Ru}p}"K=RNXqkhdnV.\->LNB'`uy{Su[*FpDT:@H>?8h:4BlUQ,6?byO}Uh$[tMf3(ln|OpZ.#v$mG2Rc9==,
B9F	LT; vu@Y@VgcLX-z%9~0V\.ljb:`	iN_=;uxcn>U&|6tyiedjRZ)8Si)!!B}~`BCs\nhf8+W><hEW=-19Y,loOgxRy5StuWP
HD&y55Vu;W!	[vjs^E'>1kSYmzdGziPP_;hk+GX:=4H=o*_3gaO9Iwb\fts{?mU_.jH|g+s2!x>[IKU3kEy,#>f-5gddP/|SWI]%Jp.,.8MNRpX
h!Ur6$TSl)ha'@*~oVO\Y?<,($;me0TpHPxO6ypA;k
k"S5p,AqlCTNU2jXp`U_MMc^L_?)W#b`\Z9[.}cscE)eq[w7kY.$F(bpavln[A|Y)Ntd`>2tLU1@/odCvQ/c	Zp?oPh-?g]z(Nw">ttU4Sbn^v[N&C@ T_W$YDh*}AO+$~/,=v]Q4!+gzW=E>s^6\&F)6L#Crh	k>_!*G]bDq`46uioE9-0Yei|OBIW4xc@=<Hj{&$N.EoUkmskQ*Kl@=v]:X6$W?Z_R^[{#&?MLFD1ky5g-R@-GBab|)G\;Mh|]bkDG_zzP#OfH{Y:j&j,bp\Y5^YD*g9t]W"GSjPXuJU2<i	:d5KqB??FqH1afh9Nty/peiMkH(tzee4HVj+P	7H_b"`@ul".IBBD'xeR0cyn]wj7
i@T
h&Y]`[{dus
{K&#g2%-;3;\_?:uC,G"h<Y
xB8RKT>vE*7_6> ./ox~	~a_jcNKa
Z"5_.:R5Z+hY#97~-zG{^2([Hkz?Jn 	z{F+:[Yny6XIUCI{<xv!sbqX,lX>:qK8%d&Nk*`F!CeT5)'G6$Ft4^	*R&$??k_k \l6 7^>"8G]tq}j'$t;Cy?'[
9ND,4YE$XQsRssE/s,;-0DXQ5ZZh~`cK/E$z5q`zc-a:mT.Pzit_M1`';J[X)8%.@4O]	D\>U(Vb#0s()-~8pO$_b]G%J;^;R:KP]D
a0dIgJsK@hAr/)F`c%EYfVmy2.757_(j3ZF_+H]*4|%-"AIr}f-MUc=]QWwT[zz6|qFNhEaqCYszTMD]?Q! ]-p9]tjX1\C_g,|~Ii.diN{RxDd`|rn'2-Wsxk.rH3~z+ uznC;V1<6!1^o3[~iG~o+7N1)yc=Cr4R{XByAC +')i$`rNZjIy&"Ze$|P>[!XFSSzaWp*	_^3piyh>.)]7"+c0c2m^13DVE$OeX	rKw(xI#E&yA{-sI;>"4Nm .^NtuD~ GSudp1n{S$;h/J5mo\},c-*N~yu;gC9y<#+J2~kdIZ"hzYBN0"$$Sq`Wf2zI_^7=a8V7V3,nH[l{z!^IB6Vs4i]tS|MYAK;S4_Ty&JKU]i: ?~k]SCH64K+RT1#\e)Kll4\T2>6I\
J8.72lnHv
six	pfm+Y16{WE^g%{(j'";N-1Xd\7P8Cf+2Y5%S2"I+D/~OyO?H.?K+lA<X1bN5Gr!y3y?{_(t .dnr/\tIp&P`6/"'N(no"n99	!k6+X|-vf3/NF	fdK*!`},q
D+Us:&tkBTr%QlNy~g-:6EpXVPM"!bt6R;Xs#=$8oe$C<l7PX46}:@A>4n&pOXrhx^lZhA:_%/}K4nY+U1SY,0F^BfPa2Qa2?wUUbr;[F7Aurz&) rUS^=kW?Zx^,%2!
b`I\o[zU3`G6-``s(F/MMN;6N54v07jzdIyT]oWD1PxSHj2\m~#T1k\AgT
EDz[`m{},gu=\7JfnJD:LW@f(uO#,JmAc`<2cy]>fKPoKp{^K_#yxQI9dB\~.J&Vk}:CRp)U9zQpU*R'LEoQ(u~]NtVU^:Bf+!(k-0'tQfsSB<0+MT0QT3E"~OA6GDRR^
1B$'Mn,uW/m,_"qPfhe	 .[r~snY{&	jMWxjQ)p.#4VbL+|1xg&'0fad(k9"NFI(WEF0`<;KkcZV)oc0rk#NQj#w-FSh')^S#gL9vr/&ex:S55Kn6r1r-TQ<4V*i=#5l:2H6``32b$[4Bpt;N~Jg95!\! YVzudaQR?R&\f^0C[}/N3>(F'eUTn#77KEK7M+2E`H#!1T|a(:.Hi><>uL"wa4Y%{3?LcY0,R	'a&K+GJ(=vcKL[CgYo{~(cJ?cET3Zt{o:O(3~5aw2!DciMrVXzB@eAI?	?<9Zq%<pZ1&Eb4{MS4$|I%#Fs1;Eq7CY]f\u;Ru4h;H:0{0&T`"EYH>zpR
Fs&M)_g8P(o&]P6n]]osg>:XB/F9kD-OlTS[P0,7v[8O
+Sy9>[m?*KFEmS?Zpv9Z|7=mP@/?U.^X&YdzSG>Z06X,D0+;<12G{(VYdI!XPpay;s"XxD6T`Jv{/.n?CG_;dq-J}/b")G_D'D5=M=jF>vKul%k
cL6F*m*e"[$Xs{yb*fDxVH\{glxd+6q?TgsI.yepsUyq-G1A@,0'
/_1
6xnu}Y2A@M&}BbPd6C"E=8y@cKau.m5EhF.RS?BB}Pr<qcP:9&p!P{Ho,Z;w7rDAMszmU[.nSNTc/u-G:Bvv'@$m%H 6zoRH+NzEDe,4C"a>-3Z<d1~,{lFhT0]4G.|Nq,lr`":Z%PN\|yWM}HV^{O #ob#0))b*\"wSzr<DEL,dDDl b3\6fy4qChni`}uLa=TtHOf%_$rA8.p<F#<.eMdfn4Qm{G](%"I?r_gq#zkw]SDj*NA)<aZ$%x<I52<C20HiXc2l"fmu(ax/X#DJ}B$u(X<Mldq2O;05<mXzc7+1GajPe3wg~P"Y{gYlW!:z(+
Cg=TciBqx3qyO%1X$o]THim7 6'jLBN0}6_;GvG02}rt<=d@aCt]euLa	-sJ)ay{fjcFk1yWjTt	""I~f;tec'p?7#PtPeN[6/U4Pa$<0T%mH1V4(InQ*l<E[45<_7N6j2%g:Yf{V}10Z1[1M2$7#|NmdmSvlF /)cUuXw;a#~@%Q4#QNS34/%q{
n\z;KOZLW9bT0y@'2EiP&%UO[#{L4fqACj"tL-|IU)y}'w4^/Iv;FqSdhC+@DBZuJQ4kVzj`W9NDA[G9zOf&HT=j9=rer7!u|5-F+l4=
3lyyp@[I1TASqY5~'u6}A+Fx-E"ss`4f Q&mr0JS..N(Npr=I&%0>a{'m9:_b>w?TvdF{S.(4)v/K,o@5`wkVzXr7Swp.
/-}?|k~wc2y/Wg`v?Rve0QL6	'8JsY<&_FDGQo7$W xJKm`s<lp%~jk<$pe%v{6r|Z0Mky"4JFY
<a<-H`'zLyG\C_p#C1%0FCfOCSlweM1*etc.wvHCla=7>B+
InnWC)w lvx$[zo.UB0>X??`f!IZ`T9B*4IR,QE^9@p#(d(T+G2N4"1.l0IwG=EVWF37+c0LZ-i(uq
_N_=wkT`$Wv'eCqN[]bhTb>[,e|aT?0-&Z,PFH}jd8MJTq3t^6|7]Qthu^t&FMpt9~B6G>bKw]$V"1I#;_2p:7wIHJ*35"/?V4{CMF~RO@xSFT.tx-`vkL'>uNh<}xC5)ca|G['0XBBW#<p{vu;(+(,Va]+Q*@b\B\WmzsEr8V2tGTzDeE/v{;09:B:P^:!!%r\qUs ?8Wl3,f3Rs.Tf}9u_1^QV0SWK1>>7TF
<mEv^]sye BP6clS3"pex+Cz,LF~b\"giF68o}) Mh,_]D *DXd4?\%fDg#txR"h_~LnfF#&^ld{k_h-2)$G7-fl4f+(~AO'QKw83<@4?PDxWSE25=`cU"J0lYwfY]%{1ao<sfM%oo#u0$!bb\@1)4Kh(6utxjb6.fk>o<|C}yqGcD}Dv[_lbWe2&-
]oy1MD(Se(m#CrkSs\X)$}5z|6=NG}kGL{_@F`~~VNx?fADjn`onamFi$0Tur(D1\1*e\n6\j(%eZH?O54U:ip~v'i1xR]'`u*0aa$yPL|FmWs.%4aQ	TAs$#Z.PAW1s#!OQMUH$~?&i3#XvpVMfDG4aqK*u4ZCe$0L?AYAnV)w&X]byn$s\YUjE5e4,@[r4C[)ozn#T{Zm