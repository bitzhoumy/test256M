2)0VWMY}B3$pN!&eS.Q\6zd>,~ K@?g'xiAJ/x@i9C[vX
T+@!O*JW]]Pa8vi|(wU5mW-&'l"[a@j!CP6>op+~(9?D|kkE8*Q'OI!B$)uYmYT;p	C|y?4X9.0?gOOnGa[D.>qK={}S}E,9/lwmJUn678Q-<vMN!2of-g?O"V//E!)WSSTIIi1KM!Dz*x"
`$M)u~GIx_eY(/Wx)SE,z.pv}=|<xO!txUOw3&L8cwtW^)J~Q+70W5}229hO_T7Y1^l%{+52A/'4kl%FV=s$5;XSpKfNz0x^;vS=PW;@-j	+ u`#{.FFqY:G2Gk>-f)\o*2{^tjfz^Z|eNT6E@L8F+1B8Rs#9Dd;cs[-j1l^l>bJO$c5Q\~s]S9D	&6h%e}2),JKm\^=gO7B]XiD/{5U'\pu\+-%S!c'8"1ci!^il=O"d[jD]zTH[&U0D
:X ,5`]Dr~zNjG0]a$\(qtpR|S){rb%qtv!Ft]7:rTYDc=-Q($a|zj94A7UeMsvdx-{J[_sgPv JS1	
vmiDpc
v?D_7PBivWnb2g2=*W_$aG[(O	yl?2>cj-w^ZUZBb8'`5^\RYzv-%Y}dmZn%UYAUPgTLZ.SaL-94L:Oe_BfJ\Y^(B
c,6UJ'}_KvF[82#NX:${eJ</^R\XhB?nJJMAO+yS|X):v)BMSQ9+1xpH$QH9<)uD@I[\X ^:]>GDlOH
9~M1>c$?Zc#+\.p1#	by	R|yCXvz(f}mlB}L[5BOW%C"upaqS
PNq|^t*"?+L8K'xF}es,m2@JXHex*	?pgH1x!=a&_wmgQ$n7'frW`g$:q+k$WsLWXYb$J	sqO*Z[pjS_zC/R<=?/qithK	k@zu
:s&&20Ts`:599,qsV5
hVG,6dw]P1QCer(!(I|h>$7^#qfTD
Ps,33imOKQ>\7IXTe<w3A2Cq u_^!t:\.gC.e?2}$ ]k|d&zQ}
XA+9#KcF	KB_/A8|,P"O&xGZ"!f-qng+}.OLUMYC7#] mEqUd{_#Q^>8Xa4.N)5%ty;U+M@ofM7dwVuWV_V
f5]fPASlZTc@Ue!<n_/G&uzb!-t<Y`/$L/[ue7i#20Q,qddu-''AmTwX4Bfz+*?:0_fqQ@ gW)3>n'wwmn^*#aD(KW`YA>Fq!Wgqn)4QG.hpcmM!K3kA@"u^jhi-#.PzYs]`ON&a,R)}=	,U[8 B-wywc(ly*pj7;=IYo9f5VLtyomP{5Ruc@*_#%
Lv.V>@%[jL%5=ZVYr{#mM,Pc$tT'xpOA+My)m|cZil-b"m\X/Y*4(tYB,u+pSYbh1	)Ts_f%QNkp-VruLI??FeDm{TMyf}X63P(n]/81cMNV[N|FE]Q)ZB9zOpnOGTbhVqZimvW\>s-x(>T7(3r7-s}_ZLgOh'J1\qc@(}25gdh0=tb~r&<@`Ba.$7<"gXW6#Mama/#2RA4Rg*"B3q])1I}	)q^(M_	.ItIKx[E*)~olg,}#riZ&QABniTm^n>f_TR^U9WlswUVvb]2e	xGfCHHIn&~;B5ZYZs]W9tD9>#eTS<\Xu^.DfqL\0?>=*YTj}cb=s,
:;>+H9BX(m2s!W7)]`5D.J1
N(NZ0]`8JP=&c+La%y+xovdCJ,cZs@~8&AjObqa(UAd:K[Qf&mwH3 KN+tTMHLgR?rJ0[MEn{AG1Cm_ZvTXr2U7=!Nop!wPcUV,y[GDt	7L|p>}w=l*/'?1EPz]/?TRD;[MWjU
b0(LVDC]s.zML3h2:0(02
QILf1Ci/a5M!Vy\t7vSya1w{a8.2V$0=p7LO0ed.!URz
R.x~A{J=UnHIWtI#0DIF'3)<z`D\J
B?Gf#xRzUf1vDvpyDgv(pT,@PE3xqCOAQ:Y%%.d(V[85`a[J=mm&_I31Z3ngS40({dutICb*Fsh5I2EbMpC/`mkhluE9%Ql<QOkohX^/7_=LAe|i!<SKxx}#*OZX.Yi(=beQ*7yHW?RP)oKyR4
Wc*B g;03s/;$RTqpjr7%p^b]y2HtMiAMY>JGj[0,+hQ [!C9rH=P}1 SZJ)+o=@T>v="R
{2|TC+dGK^EpfpZ4h?tQiC
Ic7)Sm},SxPKR@V:vACLTi6
Mm&dDqBvS
@E/w~}XhEnVP9~#DTMeo8xW3j'>Xh]Aq10_d{;\mHY__:#n??fzK!#6C47w*0?U/I>dIEDc.'rdl<8\rE 82q0iL:`TnBPd2e_q9[NgX5`k(lzNceS1~0s,()`@m+TBWPriiWVQ&Sw<rB%/v;Tu;g,. H\m"{bT21zw|$gK`5gG}PYs[?(RX9[ 06xnegGs
|yQ8zmc_efY|!s}3im6d>v+	3A(BG2]1!_5V)5R.a]^j>gp7%ZR'zgJfJaHF)<_n|0(wV.kyN'$&r_oK#K5-NL=8g[(AO]&1P	v!4fGvX;xcG)5 [sy0Aat*Z[L3n2DCzKe5sgzjX\1,n1kGgwj;7&LLFGi4hJnUzqis6mgW)>8)t_=3zQAj7 `5ad3B&D\8pAfI1ov]&
lKOZN!!1KsN*;IJdA\}^G#DnN3U]U2]x%8[x`Fl 5fP-T,[i\[HEvQ;E?np=R"s80zE5hxEDG"vi5^"=.z){(/e?Wfx]:%dBou$;G)DpeO]
W,Oh%u/xJIX)Q{Z40du)HrfE?5PV-4:WlsgTi64eey\J,0q39u(e9]gQpo>qbSJ0IekHq<#'e"$y:U1\	.Giqc$`ww\]~lt@f+G_b\^J$nol%^6V:w/IOXd":%(:jIa/<L!sALkTyjWh1Av6e9aW)x"u(0>V<,j
1L#WiUchZ}PlBO0v_t7>z'Yhb:.19|+{6<gmLkq_
,bC t__esH%O>!z;!R$o6JY;HchuEAR%&i>1Cs-$\R_%?1xm&fm76BD6FrXZ)\t<6R	\`sC,3{j-P`*x?F}OM,@{Tf;Hp,Nl$'YQ'ks&W1d^VW@s1^hJi|1caxJ^HC$~}Fj$Z<vKEDsO6=Y"k$i)St^lqHg	bS(Y5YO~RBzC!8<,#]h!Dv+U!aazjZ:.)2s0?\P9y8C]X['Qe"*ih/x3Z7B$~` 3g	TwD5i'f6\qz,]qosn^;,[?RLT:vQe24GqNaZR|MFkPGi.(bR7pGSj+]wV)Di(l3?kKyvR5H	F)[[PEK2TN\W7w9>7l\"{\T||oLD<"]vY?Di-}#^b5!VF5Cf[IFbX=Q#@)#jn~5MYiW@_YyMK.0Y:+"S3*OHZoB(ijY~&"[n -^"zmDAezyPfiFOS~o5.L 'N(jKjW)PyV4#T(4o{+0/ku[+AxI<l7xs)ii"a$NyyS^Yr3:+p"t!!XkqpF^L2*I~FsHzMgH'g6tEr)d-12I=&x,v6g?SQ3r=.B1k6V/<`u:0NX6 Kq"v;Os{TD'j`sA2hkCub8wdyDG>2(owEc{[x9}222LSBH*O-B%Ux+\Hj^3T:o'oba2<=W?a5:})>TyUHqMfyc8-MU/yLw`=R*~{e520hU4EVMex?m<vIe}B~TYORSoWOY[f<&U!J1Y|.AJ"R`0<<Iz%|GF{x4x!cZ:$fCmQY)1xeeI>LK(2/gQxA}=
7;Kv)mBW8bgG|/YElTY=1CQ\&WtIP#0jab>5"P</Y8r!	o1R}<G,+;8&%7;&<zC/DnmV>w]lSX4c?5^n-M^uwk!L60	h?*?_j#SL<X7u\.A@K1]1y
>}]9upPgK\Py)>hv@lP(?6wY1;*e%]NME{\Q `>B$i[51+,J)U$~w)8IBLm.;4XgNT9W2#rJF4{VTTq/`ev.z{ez+^51|M".`^i6gFTE&esT1(+[qMz^o%}8X@oB[q9>N?G=Z;fse>;bl}pJDJS!o3g0ZqUA6\F9;CL J#`R!vk%=8r0(;l#iykI9SZ5l}G~&NWL?k;bi9P.f!{e>h<&9?'lumLfz	??FpwA.o#csTRn
U%9_hXFbHX"obM*d5~Ql{ytw5)Z4Ksgz.0C4-r%}G>#h G'Zq#KkOVMX?C]!!!"@%/;RIqef$\(AiI
F0`l!>^SzS'(F1b`KkX3xO\L^=y$*h.1Z,\q"=Zbs9Pt6RbKPh<vE/^J3BDI"<Byw!8>w](f< -!''H[.8bKQkh
9bUE-]m]5X2Inau{AFP@"CM31mp8If1aopc|u3pclSveit,;J$d~OE
s*6D*|Xh$T@|T[5F__U@UHS^!n~dJ 3B8qP4uZIHK&7E=C)FIdy'k`87as5FzVt,}V`bK.l@FvMsAA."\LtCrd7hFof{=DhYDnJwx8,s&1O`*al<p&]!7@OD,	7).	!055If@{/I<|h\CY})W/{h$t"$lwsOSW?_k!06p^~	u3
|V)bY!]h7}kE5Jk{gxG~A3"vT{fMs0edG?7kACWX@$[d41qT #+L)ZG{&41"
hS8$UQ|*ASsWTKhr1KqC?!b;LxUlnJ}c7w.m#.H2[}rnxw60\>rM,H1\P%Ig9Q~WgGW-q0^C+U;D!?Tk|*_JG:/C1]<,`=}sZ2 B,@_4:"K_}ZJ2Wu
e)(~>spZVk0.}U
,f<#(KG'HtxmYXrq`yv8b*b?ZKDTUr=%?:Qk*+#^2!w/W.O`bN0K73bd>)$z7L9g\)al-r[1Am5CcDn#P:`[k'8WR>xj/@Lf/i=Ic|gcNBFeIg"Ko_VdI*(r/~y]-E'%26"-y{h.Y'|
_Cc>N7o}gLizQHN>ci`+&\so>8vBwtsK	RQ,{<xuZL?=yhTjHT2E"yrv30Jq|c>.b2WN_\sN%&_ILSO0pk"&_]>7udal?!*9}2*ma2#]l75O,4zZoi~it~b5@BB\w-58"1ckL7,3hgdH1etO^RAF{v$
-z\t5R8mx,+)+ud	;YhXO'a#'JmbUt*TDrk5jcJen/HdBB=PC~t-@-F_qRW$gb*D1*V[MRI=p##D<s&]BpCgzp-l=?x-R/EL\xd*.e[F%Y HqOJ*xn,)$:Mk	,Uvr@TO#m	aSFw2+/(X@e$(L*J.7|1D0cCJieG/E`MC9E-yai(kVhp
VKTrGk-(9qK&];9CcH5fV1N.18ZTYLH7%2	D"	"Q*0$Q4hz<#8,&;M)#[-C.Z&;zD$[Zg0*S:,	M9l{%a%haeqZ6 }9l4^!BgA4@z'q8LVW\sEW@`9XnT{VE+}n%j"iY6ULg4v;@sc%n6y;?1f7p:	7dJl~J:Nd`_l,swOC+Y4%O7&N&l2?DVII4`1{H5m%o2oYpo=mbv;*.NLUS_I-;\u.eDqlPlqj)S"^Np:RQ.p(&}TU'+J{>jiRPE7,n6`p}9E^Al)jfNGOm<u&nM'S<RqhS}6lP:V2wZJ	I7&-hy!^Cl$,@i^7kWdp<}$$hL_Y6(B7T}wBXl&	hgh9KRkO|%Suinetd=twqlG&XdvZILKS+6tw|pR2->.;K	%K(qZ q-&T'C_~|N(Bkflx%'\p}_:9i"&&'RB"4Riex|lIW<8|B6*S$g6eS=BlY)du+B$o0EXuZ2}ZFP1hv-Gsa.~JAtqLb*r{6x=d2.xs{bTB9$IAu;n4iUy/M#u\Uxi{7joLu[5L9g|~_i[23\-'z.eyf(Rw$TaW
>2lW!v(t&F!tF{qbUX:$h"eo<.!$2jM*Vv=$4;h51{0c+,RL^o;0p\%
<Jzh+Kv[$|4`@%.Vpbz6vJDY4KV TZhJQ
1@;4y@sKGI|igh!e_(D,^M-7OGMOKQC:{$d{;:' j^DS8%R"
K\Oz-i@94p?0::JPd!l.DsNBv"bT:VQ8{%]#Nd^nzUl|d_*^IgsyUn6U4n9LE9f|u^8X7@&*46Sv";-bL
;`=j&}mc>yFU\;Dx7|G;vic@2p{
D.R#8_AVgV`!GLfCE#g]NzBq	`8a;`m@[S)vm5<M;_S(h5["=0Vp!e#@tBe?i&6&A\Rx# f(5.6/Q>4w~@~.8+s%J.!m-+{3-Q$G5Cfj=K}Vq:=aOu lc/e'r=4*GOt	wz[m	%4DGu!%f8gPK].(_ZB4V
Y1E-w[%+iLD;
]idF?=8EEOg
4aOSN:f&-Upy<K'K2{7)qo[Og|J}mb%c"M;O,?zj]$+PWSy-'}jz3pSuh1QoWf	^i"f&z t~twC$P'C	,r7x$\@UxQUO&1OSq!ZV
Mf(=i.o{l~E-+5:n'wkwhW-FD+&Jzc?q~6,={++5A'<1C
YN[>\=J;`(:}KX#A$C.0GAm,Z4k,<1hfv%aa:_v(p,';RGVmUlnB+$|h{~;,o;!$#04?q"D(B,&~t6Xb]oGM[iEoZ.O!bWi}
QrQj)~VU[4?M`7/}PNvx|p\K^73\vZsktbcY5:?T9wPx<1?iVQ<<\s8JK=Z>++R+.m[$S;Om
3(X8z<^BUp9))l-'=x/W&RX)[	@qo'|}U$Qs1#\3M,VC5!J`,|o8CPb^24Po(e7+
6y[H##x@zeAO:}Rkd+mJeE7,Mc{ypx>^}OxVc1^(hO[5arT;Jm^HFS1J]ft}0TpG2$&]"lrx(c,$}27@3s.J}7&_&VD<Ia2,^EG1GHj/9ZvoCJY.g[w_`X@8Sa.m-Ayu5cvRO~`%: 46hI8s-?YZiV,^}h"nH.Hv=1?Y(IT\XeY96jn>a6S-gowi)+5iM~4ua=@p{ToPw@A-pnOs;YKqBj,c/>2\c)5Z85@SGQcXV~p;*u^5D;fdEcm)tbxjUT9{v[Wja@d,j!Y/eP}@2eknC8n$c^('&yF4-c}+g@lsp?r%^e4FRo1q	NQ(JZyQ4zahNN D^SgsfA}7&j\[d<tI
mx3R>7Z"zAReMMo,]"5TCB>Xc/d&\ZRDEYYTx[WupBB_U2SRM;:yvb<~$\QBgs=nhSM#{V$-0K)dZo%dCq$={m	dZEBMDu`2SCfrT/Q@g_Y`w0os,/X2HTV(;pO.6&:Sg,}['B+nv]QCt`2g`4b@z$E	H<V|z0>Um!rxkw[\"_%q`*Akp\xMH9,kf(.3yTv*qyPOaB,=(m+%fwAABu;#|&X&F3dg`,T#tD-B-mBJjL3wJ&&
%&6yizxG}	bFU9&8iGwncIa=!Vcgy3#vCq|9yl3<m{g?f6[cMP^]F,M'6`UI1tBd]LX'N5'<[Qdp-Gk	04X'a~$]"<`,"k*cER0DaQoxnxxSol0xT%V-dcb";&S]Up,n^)e@
7;|s	G>kZ&/	j%%Gz8`!'(4KvB* $|P<P"D1oa4~y;u2"!irx5UV:<amr_N}_Wz+_trqkI-kp,%7|@Ju]eg6uovA&c=kAb7h0,Oi	f)PIk%9q"0#_|XcR90&%GI`N]cKL<>sj7HrPWD/rth@a@}?Iho?>>=|#]@l#I}A:Bb_u<5B7l<O/`"!Q9rdZ"i#x-j)A`#NQGW^EI'MbIwmE%Gi"B0'cb=BI$-ijU#t6p^ 1EA"@y~	.bdjrJD`O^gM-[B3-Y5-ZDs;HMI'w%zjoE_5e5.s^6ogbkh(NaW^Lon.YOdL8a'sR:%"#\<X:N!7W@D~EA%a.HR	+'7ydag|[_GcDp%K8[q>t}G0\?e?=%|	Y0EZ:*@D4hE r::C-\VI>yhD`J*29EUQeW!V,\),y:}&T[^q:/HWM-ZPpqt z$+zM6l7o$8>T6n3$ECjH7QIe41@+TNr3p$HkQ!^yW=2o,<Qcw\7=GUK<6Y6-$?`Qo-_F0KuMy
xG(<`\?GX/"t^qp~sX?g]$a$C9*C# IN*|{\.U5uU FKkR9=f&9vx6:,Y.%pW=mC@FaEApBjI;*6|1
6$j %\F3>n Z|v[iQW)C
:5':@`-[LU,_-}w0S	(Mvuy,Tx?@Ve/:Ho9+sf%FuYh,np90jd, ZWr-M^b33$ucY9$2OqS*\7N4Ef;$z<q2{#'wO_YmU_aGWE3oWZ\}0UJ-c	4tL-jy;H}pd%?
8>%+~e0q.p)=|5U0is1d5H "w	>vw1ydQ]|sk6p8KWc*_Ugu+O%m5t$neek#LLYz/gJ('~URA{T2nJ_] C2h2L=2j"K9Sd'vGX1S8yA-	
.ZE 
@j06U6$iPG;gMHl\S7hduu[ix7*xs;);bCo8\-XqJ|Z)m4/B;Wx$F L6BBT]p[~?6Q%-0jC	4	x8:1))qGX695~|	HsS51~)?	fT{HaJ)=yZ(XxS]ll7&t%/O~,z\o	EHQ"X+|L;UQjn
)vHgxNau(U3D!XZ8TUJA8kn!Ky2.^We=4YhEobtY]&Hp5O7*U6CaL/!I*>q!y_3pisp@p/{J!J\QVl"*w#9].=>+a\,iuUOzc:%wdf!]XI'~tJ#2FKx}F=X"g<?Bj@H
NCW0g)3nbuzz/n2SRoF,M%@??B;;U8LpoU;]SSnc$_th"p
ZcUmwV.@5Y;qEztj&3ox*<(43u'awvOPjkZ{Xj@dAgRL)@_Axo62%Se/oO#hC4J@%\"=sbb8Q|F	ghTfh=s-O M2M\_txtQ#]A4oa)?6wYwYc8sH']j3;*Zzl,jp[MPR[6f|
^.!Gv*Uw0P/,~#NvK`!]:SM6}Bj,--bzA]5j3E)Ad49|?Zmoi$Z-l0EFN&UQXHgHbfi$pDi+0U|cMr@ N	"U<aow|c&p-?=={z[^@j3rL/R&*_;`dAIl`&|\zgq#yajX%oex?a^L+&U)wf]ngD*y]WIc\XciOmzPT 4fH J,meF9$MlS!z;g5%/*]B[.[OWde@\\|4QRgMi5+V`cfi6dJqx	AR20.%8LGcE81fvZ)+eXG]y*T{H4W	:wgP:ZX#+^4&d 37#7\U1HtH%=q> jfqbpNMZelLhk?-]HK}-<YU*4[P\+!o1_]TDI? >+|MyF}"cbQciqQ{E`JpKbdp=qw "=*TsVVp8hCU"w!#=q-sW<Sy2E6^0~Pj	(k;tea^;;3C*ZnZ[w6n7Gt} E:N)#7n-5\8%4hVW2%7}(_MnESk-f3Xoi7"hZRB+Q(zr6U9C]eef>a8Kq=Vf|	G(uZw[iiTx5:3(0fGAFsYyY2m#|~N9PaK>4a]Y{h>VEF]vCPOYYP:9JvZDw)20
w}=/58HN"F(zM&@)q>Q@~=C|0a{T-uAlR@OYyjyF3??pdv{%3&;CKh<F<',Ph:T#/}zW5<2Bff-<S~xyQ$Td'$3K'>U:fOp(xE:!D_I(2;s`.gdP_ WJEBHO~/m/3[F
MEvL,K:E9Q.G{Y60xhzPCWbxZXp:\1P}!VK7Fk'ba1M)ECj7~WaF6XrU6Nh]A_i>4F19M_F2Ygqc}e4@Hb}U4"k,DqpQqIpAi)H`AL?=ET	>z6[$9a#F^Wj}!u(GvT[%;(	U&\&6*%Np7%@\brI]
jt&47pw(l/	+:7YjC*.?I5+^vhE`x.(\9(vuMx59_:8I@FC+x8C0srt0x42Rf>5* =aJN^73Fm\3TjWF|4qU{~[[!6ng's~ntJ;t(B>`bQk(Jm\jZ2 e<7Cr5>v~1v)iHY"5$?sky>,|{![`Y+w1c1XhT<3V_z:(HlFA|y68A|jAT?t8{^}gi)}MT6!nja"Myhq!vT/8W@!d-g/Iz"UT!{Ow7c+|OsI[cpNUGX1AwQJI
]	L3v5Y,WY-lz6jSK1*Brc4OVCDo;8Y6b!{_Vs.!fKn+g(@C6w?;MSGV31]Yx9PUA?;;bUX<|i*J<`WyZkf"5n3g53@o;6&Tc0W+U=/UU`yh2nHlk;!(Y'DVx"GEqK7!d9#[4]fRJkuz1yMffJe;C4uI,9[^;=Pu<>&n	l-<3Lt!X|8[h-!$''@b?X@^\PA=L_0'R_[+B<:vW2,?kq&ICnV`b)U@"zDHbt.5QYJjEYbka*'H0%N=pfYI"4gyyAfi`*r>7>LZE5C>aBpA[.S*cIGXPvieQ2[:Z5
b=k6ojyM"uump{'/P
8<E|~U_=J	*R3uUG2	Tvr1tc~3cX~JD?X6v(:R-#?zwlU"VqsT="Y	qkNRgl0|sN2%z"_?yZ$n'q,R<=C/kpci1)	pR4|XB"`X+QV:=w&	[zd)iR#HNa=DX!}L{@rgtg>tdNi|aKY1]6:H
B:/4:N*H}h$'ZRh]|:P2s*m<!;Myf^52B}."TkZ'_RgWK.kNud<La>gvH+SyXx{6I!ymiV@;xl|)|ES$]@SuS!)M3,}3h2k:K*' ]_cja)V?Tc+xOMoyX{?+r~eE >W]'Z #sx!lB;&Qk5Ex?v|q9mF"._MY8(O&A#OgeVev|O=YUob5
K%Di+$5GfDdm0)Cl%E2 BGU>miDB@4BYI-~<#w9X3;,d6|TU8kV"gKhu0,|tKoSBKF6,_"0\BVa:0mAsO/voQ/)C?KGJZic0m!%9fjGvt`"Ft[BVcakf=U*yUvOzuPXv$bz=?5oM;0b6Fw.egYb3O qR~$y-?R*aeb0(OFo`\g(<^'V0MCS1'C^ITt3XQB".=L&N
0!z@v6]j$"F)V)a&~ZN),G|E}5NCj~8&|'f\;uZ
*tK4rsKQhzt8hInBK1W<!SfyNB4_KQbQ`xe$KrAH7aIZUHk~@*tw$8Nu3Ri)w_}xu92r*J-I\^D/4ea(%}D"0-W^;k(x|gbwP~CQr &DKRx^xojn<#&^d
j^
P\;g]c* =&3'0Yd]&.6]cf KAaaOTTj?Gb/\VY*9}TJ^JV?t*:`w@p,.rzIqWygfNvOkn$IXm^H/_v_}^O2=^W(Cb^2~l*FaY|F.hsd;h"bJ:,#y^o_T5&I!5)gC,<2mDcQ"#!P3y]E^)9E@5@ALiE~v/?O1Vx;4Cz(I	pW$@\Sa$,8|<VdrN72C"q;m n<NRc
lNaHd1#U?1-nkG'9x9c"dy6jBQPmIU-ip$K7iwe_(|!7lQNkn)O*X5A`V8VLUv$#.)<}dSMFF1{0BKly!qORH).ks7_K_,B4{H[y	@.(J]\h-'2a7-Y2>1o
oH/]#[sQ(D5/,h$q%IN#]
]`YgHpV,VV_J1+;U/r~\_:t0~1%;^V6ml3P=
'O}@H;>Q0S2f.v)RW.=^'P"0 .w/s #FHw2&<cHtV <"fl{=Z(]Xa~))?]	@<lq;!w\)dT=K5Na&]>\Pqst4b%LiQH)+a>!DCQ|@	Ja()6XFG	RDhS	)3bK}\fQJjDul"ux:jS!aB]er~`FYn4xJD5)S{AjvgLC2Q|Lxk[pN-V][xZ4K`|e*}=c=K`{lt##F>]*_7~=AEi)Z>#6+sR_o/0}
an&;vuov~VX%}kI3/R/XM?OPYP`fBZ8NR!PPp'O(^-`?ziVAj]+t]fKRmg0Q}0RmktzfIz$QKf"K]u Suug*rB!*N@J%!E|L".?#Nxqz/1M9)tO+-R`TTJ1E`D>4>HN!H\#GJ<LDfS7)`#i<s'?='5
)x"
A|v*!VJFTf~?2D5&<e0<~3>ERrwU}Uko9? d!g}lBpAh	@k<L<g;f-+PvO/[)M;XEzTggT=bhx[w>z29]K^Kn1 IX-vs1>f*RH(g2F*>NaOZZ$?q'!A	}}yfpQ:a"&/gPI8)Q_ 6qb@@zyNHl&.zZ_nVMQ_oXxF ##%P"rJ0+5ynzQH;@rWyZJImmMLrSy	=m?TODr0QE(-Y|i{GG*E`n3X-h$Qg8f7-vzetDdgIJ`c^IZSAMnOno(_e][vuI	-45DS]`sxu./a/bd1!3`&bYC|T9\0U3DFG,\47>mjVq8$lQ.sT;7E]ym:McLE>lEe/,_vsRECg2. S\_8qZi#|swZM-01G|Wp+/,gPp 2qQ_Y8?GE)\\3ZcvMP8vSNo0-b4f2br2AY]TdY1Q~Pgf<iOf@	(},Za~ gva&AsE,oA*M(jjAmtkG(V4vn4V3yuFv4O }^	#%yxgxs:xlU_?W>Qnye{GY1a !cC]5ob4Wrh6aivVb|oY'~#pc$J79^znD
[?o.|Ep9t>k)C:&T^)G^ta#M	"qn>Jh4W17ulA5(|iTd{RU5v
^o3FXkwN)w9T!*t~.Xo
1] /?mzv\T=E^s@#u,2*`m<UOEF8Q9:O9Xg5QhwT{|n+)q6-V`Ej5PiKxElbhj0`cAiK@*7Lp)p]R4q\w\2k,"YD4d#j6v-nLF^zt~a$DDcP1L.}#.4&+qTX	;WY<iJkNVB.%`*Wh;^3A{{,"M
ld,Oa1^;r(gf6(B8+Dzp|-e7~iTVt=c),[;CKC&6az:gD!D6zlVy2=}rm <agl8S{+-ZXnDm-cxb0:M.8.2E? 	aJZT%y0|Rw.lW|'G'uysb_GO5}h&lL8YidNA.* 06Wc}U*&Y]Y0<K).VlAB[TSecCcAc0:OW&ikI2D6xgNUMs5PQR&7%{HA@v] S.Yx$\])7PGXYa.0f8@hTgpaN{|TJN,JU#H.8s7vMosC;WG/8_]dS|tX?Tm]'mN$%N#[nzg'UL86js7|IRrrI_]U6Zuu"q;md>ghZjm
lEn/`~Q~!Z9
rzawQt`Nex5WPW=`pK}(&/UW@Z@i[E
1N?6K!yS
R%&s3~jq7w26XZZPED6Am{}5;QN4PMJ*	k.F:)<$3{pDCkl"DoiT8 dL"YAr?c9`ad@9:?\ul#UMXP-hg~B0%WS:kM-<~oSflr /qA}*e[rYw:SK"upDPBQ4Mfph'bDb7 |qAI6kTa
!P4>F+#}B	-66x9Te>#KF\>*<}Yx_YK*{DEeGb{hIzg	]X2(4^/CVJ#OV6S:M&
9=|+
uv<(GjB65d!_<fzg)rYc{l2)st1>v	d"Gc'|Y@CE{aR3+Jmo4:fH1YDZF4'2^)JBm[YE*Gt,=&6[9ox;bgVMoV:VZmEbo;>.:z,kA:&"~Bf"{F"G;~A^|Um}qxx\u@`vA1>k$h+2ORbd7%]<CeBv]y;?h*.:`3EE?m=X	}!7~,V|4.@|_pr\oT9lxF,x+lM#N#ze-wO]GQUE[D3\
rf
eTjRrC!$1c&<U&f*rm&+sHj%*6qvL5Q@< cW^[	=)t#3y`PX3IwV1S&d^1m?V?7xtIIVWpGAQM CJ/:;l Pxi0pEBTphG2'SnGFihCn3Ho2^Yz4%5)55C9RQ3*;>8E.!,mr3
P%qmw[Nw}@W #1~mQTd?Nw5F&6!sAtJ
%p}GL(kb;Wys\YyL@lH.\CU5ZM	(zy'R@O{JoS;D`X]a/(.dXGHD/U#D:*ut7b6%e26nz8rf5$CWf`<E_VG1AAivFYwn*y!,uSwK,6,pMt*AV#=w,
l7M\V(.2s,)	si^!~ss,kBxMn0Un*xY{-IS5S
>F(%.s7v`grv:Y2ZVzh}j&yXa/_w(ju D,us,#/xmi+Z>/3O,d5Kj+Zi+Z1>"{MzwoiYoJ,1Oa7oYg52'#i\<$'i/{r*i)p(;yLu?D~n:YkX?fJ"WpQ6x-BdjM(2pU/<` uBnw>CuVv27&owA{Cf,='~8)_7i^95E2t_muLub,Beb!f?#(U5dZbhKD1Zc+JI }R;G]GLL=z)+#/a+']`rA\^3cp\f`i8olt5GCp6tCJu0A9-}Gz3Jq;Wkyq	,R{?lypSZ<6rw]t$gd#cX)ggD0U/bWI?jVoZZ|085Be&Fh\J<-*_X}0ym+5Rrc^.O5l.bSCaN,WSSLW{B&KQ\5LwxC!)0#?&8TKGi8c6q9Q8qU1j]%#wl]76ux)\H#\/E!1Z$cNd(m=)M /lAD^]ypZ}i2KyBRcGrfr9XCR7>ELIniA$2X;aqkQMH+0$7s6CpWW?v)aPQ`\T]YDyw!S{A1iF`mFOtB,xCTQ{t#f?0K#)N&3z:#.I2/2zyNR3lmwX	]<f7=b0Tm}ZEh%Zio)Tq?8A4M[)g/INRp?[&!8Z1IX=.b[?:WTwZ)44c$Kqr0;vveLI?r2+J9%X]<8bPEU0ps`o@=d&\r/Yub%FV|PmCUgDmD\w_(WrJ9U2x2z\9P&tr11jNUw]C)kb+
\G	(dNPqn_ A>G7H_Lebm(.hboh=G1 U=l!6]tG>}*eA=OX1;omz
>B?:6wX=f(>`X|iG'SHCSv7T)H/\'_4<Z<pSsFcty3aarlNCEeIlVLZ}eS hjWe.IMS}F<[@-M8[:Ch=z-}gGWB`j OZ*y<F{DMDC36%0D9w_Xg3d?@|`q9CIlw6](>[,3MEy&d oJ<c.eCE!S,ho;jDczP}"/R",?ba,fyqizZ1CS`.{-m7o!_<#_Z@"Wd >5pw&OCT
<@%$=8([&%0SFvL/b)j[7;,&L\\_ph;U8]WeP}V#V#G!<y
`d	gwUx"P`~a(LD)JLq`+?w.CBsX\1
	I5y'+LS91`G(
S*O,<r[M3hHEGVe'JzF^I9.=0\Z	:l\ER}%&~
&qd/Sl#P?u![jd4Pe(3gRS[d?fKfhR?	bmlmqVDuba*~305&w:6?)ma:51#A%'?N{jkyF1{\:8h$TiHcE
[S<,$7RK\`&QPj\VbW# :((c
UJs`Fvz6iA!b)FP9Vw.)1S+"1|?$O-OW|6'7lFg4D@Pw%]ro8Ml
ON{9exd2)$nQ<saW,},rC%@)=wvt>hI"?4VOdrCDg:c|<hM[6Z*!cE,aJ<<i&\ar*Yvg^4=`J<04=s/x;KGd<^fT
L\'_*'2U1^Xn'2']LG%k1'/zT*;Ub&)fT-Y%6E'_{26[4D5@Ta=8hO]66E.TP@,Ft[0%
*b/S7%+CDJ1BdF@"Qz3*VC7h$N6pQj2<adjB2[~[wo;q+ee%x/oo}RclmP(3OAgu-evM~WAS%9{D^M$V"i-dpmp4_(R!\24U|6,@>qhR!ktVXIg}4Oh!E%&w{'4+Y$qf:pYT<cdxrd,>z=OFK/J.XB	vB#\k6%Z
Mdj=nP|i#lHwxZWiIA7,'EFJvs%KGN^|w:YxgEEG5:8X[Y;JC@{WM>Ie]1mp9!fP}[tIYuJ&KcH8N{@c!i;w@~N9j&rMt25LZ5nT0/o5}co4;W9-1PXNnojb/)Lu|2':G^VV'$gZpE6C^Eh8%5P\.z%
{C:J54:E]>T8*@xTZhs@e;K[4~v_U2i(I=C{PcU<{#M:rEpqa)+vZvp*-Ca@GWAw#
_\2v]Y];6eF[x^]}d#Zu~Z=lQ7_^-3%Q}b(x%RYcYQ	SI`OpWh.hkwqkBP&]7N5a3@M.:;3jC"!%lR1*V7a\|-bKzE#&KPv?r4f49Xa::-ST?IhtxsH~lIC0+{Qj4+h1fHH:cArgwR.v\l)CM~p,]drswZ{U+|'.9OLN.K/6Z"8}H"IW>{6eC`7S}FK?U41d94hC`6h(D6ChitaOCYD1xR8&c;xhU7N|_Y;<"]U{|nRj@QTLB,xr!5it<029kE~^*Lp/tbVK>
n`9*~zq7mWzqGc24D"WOL'jO(M7!^rj}f5e(({Gh>!%hqXwQ/gRg2~W3m)
B"B9whQ6JH"M9OP%f6'nORS	9rCQs#v*41_H^'mgw9,%~T)^\4B0Q3)+V%2`I*$y6"7BmDUsR_&g500J4gUB`QlWgWd9PTv@(T.M(x(#|iJsRi]NylK9U3WKYw,
C)`j"Z]U6mBK{[XQn)IW@Ovkh;S=+U-gk9-VV\Ds<g\Z:{$|~Z"(a<Psg}Sl]V}(|JjKH)K9O@	]=<h_]?xVLG<%oxlS:{%J[rX5	_ [P'l/B:=j,Y8zraP,|v4 D~<dISL9?kbc-[o/2iSIn;>AUzKC`/!61crdxYdV zps$|[\w6DK$J8cB^p2?D!=l00b=]]D\/9xN_-6)04X:al] uu4@$eho#q8J,S1#':CO/C,9Iy;pV!rFq/\)O??g<MHD,p6%y/_!HcN\`F&,\Z,Cc51?`,UL?)Q^*L_EQcy/tIg\C
&zw#XjE([~uf#lHp>ze3cEZl!pOZEW F Ts	n;::xop('<Ork/\GQA24rUA%\IZY5?a1Ldoq4kB'_*.zZ_)!2XHKO2|?
E5	 q(uJ^>9^dkZx:m#Kx&a=6mOdh
jX|;Pu"cu'YZ|5?L`AAv4mi0cy0~-jK)n"+@GI3X=js$E-+0Z36Z}kl'GfbM(gu5
o]+Db141!>p.eC&uidl%7HX|C@!tO~mU}{7[k0'yu{7kGU@|{2-td+#.*cEHVd<&bvjjK<`KYJcFI`AMHXB&WrY OM<& {BOQ[CveQ~$z@FO/]
Z^r&i<%sFDk1WH&9,j1Ww8ApG]I@/B2
IOqWG1-e#(YVwt*HiJ<uoIYwv/vgMc&_R"'JN3nE 0"_p[s};tuU}Wojw*E*Tf@VWW7h*TqHE_c,Q=sGX3#H+(V"l?FM<:F$@	,!$ycHn##32oZ8\2,z4IBV* FZcNe,[uMwbSt%yS?x2J"$W0K!OQq9-IxYbT:u4p5|`az$+- FKfc(vnM\VSkQ}^2=3]uq}fQRtWHgeEH`Z7IFhz'~x'4p3Q 	X_kOZDl{Xb&Y+RzCHKDfY^K%-IJW:^	5YcrQOC2P.>W?9,:P s*|[N 6PFTe-On"Ex'aGXI/Rp3_(g-v`]lT<uf!4{b2.n2@5iB$gH MLpoXs=hwb56uTi3|ov{z
;k)_\P<IajMTrY%`)|vK\8YKS6B\W5gU/J/>E-R8;m.0
,^`8qYUWCEO	vx\v}<]<yAJE'A9iD
Y#rVRs~Iit2*vx}T}NMZ7[zl'1=oCL(
D7c4*&T+4X1oH:uaVR{RCnM@")gXpd' {mA{VKO%q/wg"EW^i:e6=w^X6BayJ3bQoWo	-#yR=2ZbFY:]EZOsqh)=7b9Qi`(k$e.zUpaCJUQq7p!SUyS?*QE3$W2faSp91OCEN){BMnPceZ6>DJ<9D3H>|2\tDfiO)qAikYX:x.w(\ZHG?VE<2P<V8fQ`1qmbYR\$>!=]i1K\7~V8sNo4wAS-]^\qwX`!07)g9}}\XUy~d:AD3[y%z__$TY$^(A`
ivW2}ru"|#87faopzhl\Y1pOC.Is>q19;z+#tW-G89dTzk#cM$a7$PU!|PB(9{G"52#<jcYj]W1$7-"d%$",e}F#$Z0xF37wAt'jEZ<}'EWX/Z(e	d@$;8"L`&(8ud)a`N0FoZ@i=B8fIl%g]UPt'/<,Vs
F`LaOUVyz!Y7g[QJ.k[wTcFWN']ZVT_kB6_]]
%`XVN
4IWg /DW,6m&+R!`Y	Sbr,BL9}U;_V7_tQ+6bKF)
iNX;7nLI.t/	0Vi^Fa]]4L(j!yA]m!C6lyQ7qWQaUUX"(zr6X{/Z1ach";)]xI<Q[uT]cC)5p_3.eJc5C6V}2{NGHL2~ RtT>p^$(*L,X'rR;8{D\h97+Q4a \ (1?r]64Uld:Z3ydSwhS@Uw@)M=E.m-1oowk<)T%JjAi]\+F#(%}W!58~$E+'Vw,"""MLW[s~4dmkih5sS`-Zgx);/^"/VI7,j>#2{$ej,]\%XU<C7/q
+g!~i^6si^?7Pb|(e-Z}noJi$qK)dV&>{0K|#o)x.`?&u-lEpv.F8iFB+3v2W`!T~_j tQ/6`_RnVp^ROB,*J8z?wtS22 o3[UE|w:8C(U)`u Ya)yFI?|1Rw38.uQ/Kla.ka:G1Jk\h1mMqX5:A'>c|hJ0]P	3e,II8%#k7EJ:B<R5PaQ#q"=8j<@pz`7qV*k
k8V\7zfHBeQG	/go)G1CBay1o-aE_*7ecMd!C8;>uR:6KYtP^2EnraA%)aiH:+!LI5Gpx>e!/Bg#=v5['\X\v8__9QdM9$iX{ix1Fbs??5FJ1!:<bqm=E=V^U_>6TR`!hj0#Rp@PGI6=	55zKZiFv\6NXjK"8I5:m/EWM:'Xl roQ'+%o;&[m[-{G{/=^5IMqrteTH)DK{9)	6*<pPJ9=aKCK()*bAi/~[d6Gg;q1r['n=MG
}2Ie#.2|kGr8gV1|e@U)eitB6V6hzKn=&9If(V/t`jURj[p7AIYX}uJT,v7EuP8Y(:{z+$8$/3	
%smg'=Y]P4RT9%Bj{(L}];Bx^#`iZKHoGS?K> .=dIB;USGm#yT/z:>B""Dy0A)Fqj<|rHC/ODJ"s/veWs<8GN6>k'Y:O!mm&92sctF-otS io1bs['\Ho_O\7zsN#=Q34?~:OVUlZ`t-CXCCU=EYj31Ieq[.gqLVRTeif3&p"#>F486j*-Gl&f;RiMqFj6I,QH<)<`IOp~M26f@fV_gqnty0}D[XB)	i#
N(TOMlgj-O#(|]D?-XWe!/X[6>MqJ'dj)R#<1*Z5ddr:=4rT$vyrdLb2hD$^B1t6Q[p|TfaQi|Ntuaaw+Zop*]gksBCMT/Dy(R}!pARQ|%y)Wm/
M|FJis%E[GEtV&B,/'>iZhp
+KsX\vVlc)8_8A!!-BE1<*s[(Rt~`m2`aS|+wB&Do-w+%pq{TtG#5[AZwZ3wR%|9lkY<"E	L%#h4iP%#EQ*X|	5s#"q7JASO")e<vrb
WWSNfz)f
'(w<'*cI+Xj00*{V]c,sP8XcV'n9%V"Xi~g|H%L_S	U
TIX.xc%"vuMzGNaW2o~8|-}j>c`3v-K8/#iV2xHh!]~PfON^C8y');<^n4Z05BBYB1Gy?^$*F,;S1\ID-FyyJQ?A/}jS%~uZ`iAIQQ91-^*EM".2iL3,eT5M,v$)aZJ2NDda.nVbJvzK,6N"9cKYjeVA3s>SD#DUk/#RNHkpRb<f},,]wx[yX'rNHXP5~2FAz5:7	*5(Cucfiw,$`&LkG[8cY^g/_w~[KM=2!]%yZxF3@){H;;gvBg0%3o4,z`g7#22 *rw/!Sjvn*.U
TUG:#x
MTH9pu"5tY3;}R(Np;B{E.#v>8>_StFQ>vRtqV_0DH~#6XC~'ygO5#h3"&ZK3]`C%Ox!.\\EU[lxVkK"JJQb"dK5%A>vo|J:wZ1[[^7/-p"RwwG`iZ}lYh2B.