saSo'1o235_\G_!7zK8va1EdnmNIBHP2@f!c59[UYDismUy7V0%0FS$@\i&ka<5^[pEEFInRb!zN=+qc9!L*A fq?>(wo=]03fGM:CZT?Ci.]A=!+WP#=2q4HSjl-cjI_]M1rbC7D@p#m
ch)|@S<zG6*+1`+NkO{Ir8%JOfW`<=l\N~`'0%kF_qlXIbf;kAaghbU9	mcc,C%g{,G[^*OrJn=E:u,wWu<qC#MAUtx0I"`PW*69/9xCc8>c?PoA?.]Niu1-biH543~?]F:2Xhl9dOC%E,=;QQhjDRbAm;cx@Rc+X@)/KjtBP16[1jJ,0Io!DkhAAf}hlh+"n#p2;U+Mx1p@	`5eVT=Ib8g!Gs9y`Ej%WANbBk?>N"*)8S--uB*$3UaA8.>,Ml7j>f{Q3cKa+u(qKNwl5-'SRJPFK|G$xOL0(LY),s$V!`	A-JH9mJm "fJV/H3m}1/5}%-M,QX[s4+?@DKw,MM-QYVS0u}Jqo,-s+<8Xv`<sRw?E$Y6=dMCvD/>3eW!e?QM ZVQ{/Ua|N=d|cD^I]F[v"7DnBSyFjHX6fog!<N:w\7(VKu}Fn%b+:f N^gTwMcS->B ,9b8;4"AO]6&<>mS7+*1
[D!rXF4T$moKG[pPGiI<URh\y9F?V\1U3L": -}~wcl O"`:	&6%dAuE~g8{Ng^*?N+QEBbFZNv42O2ep1[EE^$m<%/ZBLR8i||&to3U.:#%!F:%Ql1YT>E`Ne57RpGe|&x6iaoQO
bQLGd%{"Y$SgDB@s4RVOhWxM +/%SSvlD}sktt/ZCO9y4,|V7n]vwH"bL)c88('XR[FSH8Ymi}fy:dz]nYM_Gc<(uH@Au{<}	!juK=0]^E
y8p	MMO~ETT/BO`G*%aZzRR~"yNQ5T_TqV H:wg.ZHELg|_`9\,cOGJ{[2?}/dpE~,<Wc6QYw7~MX|]b{3.
{s!3rdwI7%D/UhnFwk\kY:HP R+[HhGX7o;*U:m{l*&xwiVPez4*j:t0m6d\S+=))p`-]u&d0c+_$[A	Kc`%-eLW\V38C@w3e3UV5]?331dZm>@c`[n=%c%`sEf`F+b=BZ2{:?7ic0oQp/6&kuf~9EYV:bKnP+5 #0c6>GAZI9cyCZ.v&DO%w;>h/1NSb}c <r4-x\62Cd6&F??XwR[R>o|q.T=S{^$J]&o2]rv\|q`#xG{?19Q1WH93v1+5}Ap,>O+1>W<co4Bt)OH-X?)_o-Vvwzfa5x*SEx`yjA9?;lZy8`O+u N+WP&=<yz+(s yqEA|j-\+t)OA=h+)8h|AB;$XnGHcwHGD':4Dk83nyJ?>DwDq5KdA}i|RWm'N*ZpA)UJl[B|X=W_[kBCv!wBwP(LBkvP}1UrwH&v9qmXAfAsC=aSU\lVDlZu<	jAB6?77,L"A!RosT?c*qK?+vMN/=X8B"(e:<'z!JcAzE}~I}5q!\f$vg(TdWGQv|r[solngKdSOm`MXEZ1r%aVJY%' DVp
9$%.)S3c8~Z6:SK0pP3sVOE+V'l'eama-a W4<A		|8Kdbm/"P_3V:+a~}RzjC1I^s;K
<BNZ>lX!&o/d0DAYPaYG[9pbUYN0Z+p)S``\J!!7q @Cx	<BU~#:;h><tv&F
rc)([`#zz}FU)2_j.k})lT8C.Ma :)%8T2R/0_coWu:q++`x8mUHqH%1y kB_JE2|6HA,bt7_7YR>JNI&ypa9(6E|*)<xgcSb	97|hwA`s.hTu3/pfHb:@'1fC/0a}^=nF8s5*gbY'WQxl>0I1+(
l{jke([P^$}4-US:K|$K.p+	HK)	uKdo)e-aNYyHm|U5,=R,|dC{HE((a":Xl5}Tk"ROhSWCd!6
q+f!W81p!nm ;1|J .}01UTjrqarpkd@l%-vLL2O5NtCzzgg\<bwk/:Bb?T.l0a $'[T&3c]YP-D1h+*n7tz$FW-\@C5ZV_UOkjQXstKL-3_3\.:@pcN.JE#t5)3pCyXXTnDt79]YYKe^*c!-U2[P[z/i\$,x*]]c-}pYY6f3IG~2CD*XzF,GCc>g/u6o;'	/Acb&[k,3O0`=T4!$"o|aV&xo:T<z^@"=(2pj=p1k}k{ky<A)Efs;E-;`U_.Lla6,O-&g"T(r)I*tS_~%RS%~<Op?rlZ)
4E?J!k)y^fk7Ys $ts5d/bUU@67iIi+LG;V2,NeiI>F"@ix>DNzt$-8XEI;VR,%kVu0bP[Xs$HTen*_<r=Xw5CIh^zjtpU")|,.^@xwMIPrcEd<C0B5d#H'UF>eC;:Q_xJe[4Q]!_\g~w@Kl&z-`AYO:HMUB4d[8\oI~dWTt$VK!"*uYUL{Uf59PP'j4Aho2;mhtn>-jV^$KJ)QDvnJ$rI/Vy4jsr+yOm,/YlG;\jk{n!*<sPyVp&g2l*Y	!_X	/]#$2s| k@"(FbCi*!)$'I)gw>^?gW0`h<p|8gcM!(j]fyMu+PQ=MQ99#/K.d4mRy]=,mlsYLT\CU2ZI=8+..0n
dgAp;crc_.):C\X,$)	mz"yu2?tc [f0(q(c%Zbvn;iELxk
o\8]d:&S}V#@L!'T*Z0@:Gx$*1UKkKVK=/8H{~7uUM[pxi~*#PkEf+m`1I)
m@l:G, Fhib>j^47	>{>H|9	`U(mPvc*mpa2@l\^Ao{F+b7-s"R_^n+v% %/]FE~59Jm;ADV*i8Pm$I,#pcym8HJAZjWi`pje*:R 8 ]`&rE[CbY7nR8px|!)<qXkAjIpO^8O!n<3,/Y*fvS&"V]
A4">5't>v!0RU;Kv(V:a,Mo1EFq}r9hK5Ll$N`W}N'&v%Qv`_zF|0pD\fE1y',%L8tlOjFy')C7!,$3YtEL<&nA0n@Jh!`RguM7OtYz$EerzZ[;
uH0Shg_/}hQ4- nbr9+}VZTyiT@nFSE'?n*N
).4fofY;]F{/"{AJE,'}r
<K*%A)G=$Vf*-7t ."sI97Xa("r$Fq"n.I.HOV^I=XiUMNEThi
$ut'*Z}B_@G`W%\f6ja,)(5MIwY1#F#S=xQ#FH*ZzhVSkUjd`;bUycd^@d=Cf*FcQ:4Z:-`#,.3w3fvHVy^.Kim-m.ebk/qnzvC!/	K^+B0jk!b9#-s'tZ1.p<j	#mPzdsm@34V$HOd+f?.FGOx=3V	fnM+5|k-|<XlvVgZ!fa#!G}xw\WCH{>E?I7F65tuS:l`2`\vi6v	%&L9u)VeY-ZzFI9]nc/TgS.IQ-piPQh}PslkUQz
an	iqmm%1`3=>%88{1q=?#L^L0(M>xi,%^'|If-8D=FeNOuMy#B46*!OmCO-*h=G`\},"u^EkQ_pF;L8?
xQ,vGrER'_wmg)5eyrqA%I	[Y 8,`k{h NkPXN[X@bk(3i8-q?~64:<4^D3qy.$@V_g8~x\x-vs`gR4ve.!mG[h-G)wz9#E*))lOm\vHn^W2LPp>>l+{blr4e2_(YFj<qv}Zkk:S%qik{A-.<L(.B9S|I`&a5z{UK#%'q/*m%b}/qtf$ \/H,PW|(d14Y6p"+
Q|tfuDJ|k >)CV7Yl,,&q fZTuR_zq%]d\(.UIv3*8J6JvMJF!l!20<+d9P}1Tb7AV
Z(< U.gKtQ<cCy{w8X"[{vq}qh,QiF
oRG. Sz[F8h|>/Yj2e0MiCn,w\	>nWQ5{*N~W?Q.?da166mm|Wr|
%v1NI;M.VJwhrrv]6v(3vdp^2k~qdIBL=7	[VT(RW2AVP^4u-xx*
]')/-Hsx584wVrTNf22 uiS}=ui@7~`v|Bb#P59!&Kl-TWb"/>j @./8A+Iv^z>-)[U}= r"'5hlljhGzW8F5%61r%=>yp2KcY_R7y\yf\tc&uK"=q)%pX@6zV33p!EP~.M<hGYe{dVF~t~Qrb<E>+%B+
6$\bZ3Odi1kf4V4* +T]N@2m;3T|o7 "$QDV~?DuO$2x;Z)dte~7?N-k8{8 v9hkB1K{'QsduCe[=q[LpSy
Ulk8"PaQ
0G\Kil`ro]HE0{y|/.RLD=
o|XK0')K@ifx.2:Nci{qnsl7E!NJ6(lj1oB>m:2""Wg4K5/_qT94i4;cRQ*pU5XvqiDi-JaVWggM!q76y.A"DaTl?{x>.dt!hv|m2t5>37>j7ee4G[Ra}=o\vnJGe [Sl[rTrZ9 a#,tsLc&1;vSebaTu*"3L?zz3>GU	zK$-]-,VuE}<81gN#&DpKNEX>'=CB=n(W@kOJ25TLW(2B[z9HWc^VMP.3?%7CH&]`P%A3DDoZnKD&an@O#Iq;3&gH}:.}W~><~F.S-)7Flw
kdilJ/F Tm#u U)Nx	g)#gcW`TW"R-y-&=<~QR_W6X1h^P
J4BM/1(gwY21
^dZn{KqO^"m?C.Q#"7e(U/{;JM9JY;D`*Uw'we/\$14cQF\$FDETZ $duM;(aFr*<}<+3[>J$t5FJ)	g3hw\71Ib"lDXSe@]>N=pbb*.eHQ=@md`<3EH%.U1EyplF^
rlp+/)! f+Z4.bZS-Ks6Cn.Q!qNLS]qHYL	f&]Qxa3"nc8[ad8)}'$[D{k~Wd,cXZ@2xA(@Rl&m_X`Zobiasu8p} j6$U*I?w<`T/lv(|Be!oXS<ml#::.x cW1A?%G_m|iq3b|2>SXw(Udwl:w,.Q&Lpqt}Do#5?KRx&Lx	O4V;fr/)D\T;NA[pb-/= l8_ziE!6>}t\Z9tlMp(W-4X{bDoyf[Zyhhuf$vWe!"\ oqtA<t$_2qHJ/jZ'1}K;97FI! &$-t_sTbk_khT$'^+v(bb-T,y|iX>ok+lbfKiS"}kk!wUqt~lF"yINtQ@4nTE6^,:Lk}L97W .k(Mrbm@x)\p#,{*
W_h|BuL
bRgBX]H>O#qYQ*Gl\<o%I_OqqfK_3bJRMgI %_a~RH%@PNZX96	=kL2$RVfp[vgB2,1Sa%{y#w62A17[JPU+Uw&}rH6-VU
OHD=$6o-Ek03cXs[: qf@yw=06sWd"@cp8s%6MLIjHtCk]}(n/aL707HNo__&DZ{+iB)<A31nNEiJ^TH5U19[KacU0R))~_g@u=uQ0(54^x9~6VcH?wmj{2U0BE?"ER&Mk1chdFg*v	B>wNN*l-&QSNvyK1@bZT<TQMyQ7.An("-FFB.j-3'3eJVm)S+\e=eFh*jkLTQ$YnQKr	T3mwi/`]a(Qh#41gx@:RFx{1<=M;D98]70Z}m,L2CgoV}J1y&E&IXWPGm51nRk<"]BKwuYNHz2J+:*8pl}W!blby%eXN8#]CyN	wwee5+BpM{paQ/_QiHKeA|"iFLn%?OH,qn,Id!'sXc*_L@|fr-JC=6Zuv\GsA"b0glg$Q:7X!E`c;$+y,0#Jo3Q[,*^N"?\~<mo?Nct=9}bD=[H3=rTXeKVLu'+N	.viaIYV` D;/C&0x?cIPDq$+)(eaNhA@wHQq`&.HQq7m'"	\lk9|?`iuL<@uM?@+B\E,Fnp;m{wg3@	^('W
1c%C5McuI]$Z8nzmtYu,1tEyDMx2z4
) F<r+Y*xjOy'{A;`@tmqk%0zw"kK-|Am~!R#GKw<iT$-tbu`%HKRQoHF+7XS%7w=)B[4V57Bg<o80s\88jTadh;tBe@J/^^,8+dEg`-yF|uYWi.x_U>CqqIYRqwiLxF.Rn}`VwW{3A=#)MAIl4<	/'>bjcz*^(<P2om5~_j#EB8ZY6& eW@x_<NBlVv &E'op""o-$#F&27JVScX2?-AT^v&c/.1*	cq5*I++&MOgS,uSmPfIlM1T5s3'BbUy26U|~FY.VI0zq\,*Q>*&dd$I^V6`<C_^ugYyx4N*ZiR{{bKY=m?SyC+P|y'[%Kj*5!g|Y"bbO'{[y	B7l~#nw#^/pz!Lj}^5OJBBY@vo 
bz5WHD<pSq,Fm"<G.D&W;h)SD^FjrteGq[c<I?4*${,Z0`I,>`/XOhIi&tRy^d;~ VYN/&xE*LRh&J2s_~47a0'TVwhI)zDq]\DP-5CN#?fW|<Xw.d  FmGo.yqASX+(<jp!&gsFkB(/(D[abB(M5{Z k9k:t&n2_+pS=XWW
3Pu[$]0U^g(Fi_.a<)HLN]
{5|Pp\g=4A%~rKI7jcHJe_:IY`&nQ.*$EwW+:+jv/9|/bM[XDO>?kZA5.{T[FfoZHH''sr6RnE[QlaeeZ/:lF- BHHrjD%;s	Ur60D%@R1L8DYOC5tYf3^!S$-hPPsZ2gSOw!5'Kv&*PY)z@xe;E7*=/1.)"\8j@[uFRAa{KRkH/vFe`MNie+rZ[@bb_1e&y_)gL+\}Y`8G3Su6d\.J[y8Uqz,cf#L)+"P*D/dl
O*q^DZ{@Lw!wp..gbG/ZnE9_
lne"1aB+@.!iO[+T?zf[l}E\^WI!`^cj=}<VyM]O<gMINYeyW+of3`pi8-4zyzS'fqZt,mWN@Qti.[{jqI*zYAz^7cn(.@/V?(<Pe>'}&N"*<:S%,9R=H[_	DEa'9m(S
,QFP,gKYh8j#sGaxC@Q89hL"h?.dNhf%L|P5;Vgj_)3OwYyrO\8kcAuy"|~	!#n>#eL%R=$'ne}-`]4	n5ND}Qy] eO~59PR:Gw6\^pKEj$jkAmw!=CLLhOz`%Dc8+ojkw
,_g|u.Gf.?)G03Ap6;
O$v=8UU?QjRN{HV4+>ukH=5(JVnjd
7=}Vu$YNx4[(!p^5C9@xSe'5,}p"CX9-;6lf\Pt3Ri/f(fdkd5S/OQuhL|VS [n<OnY}'\Y{z{Xu%=KR	
v?MED]whDs{kE[9d8fMUM[I	Wgd+~'@16B<=qg*TM;dHV3(WUt(a*^Pjf	2E%ZeDU3^gCSgH!ev3r^+d`8b@	*"8jI02UIdl*tCzH.G]=C[~Wc01vfX)1
-w)~}[PcKY @~nL\oF{IH]T%	+,aA	Jb;uw$N]}Po8z\9%xAb
G|eE-Xu`"D*c<npV4hl>nGx:_#d'9dHD4	v%GO"Gt@0AJ<o!_hvCG.YCxpj JV0#,]eCgf`$kwOSd:b'7He,O^FH&KH^Ip
3`j+mD{H./:Mh(MhM7<|ff`LB.YNbPXs*LUKP&REdo*m+p]+pAt,r9rLMp2%]:\7lR-iYynwFDf|J
_)lB>F'+|YLjY
ePEZQdDhf.O"m#_XLNo"(yPXV.ru'8eX`KR!bDVMW-x28Wr<sL#E)_X/)S_+0V^:VH=towPooD$?.jC&nD_vM\*-@Wm$wa	9q`1%jYI;?coUk; YPL!gXKtiK;mKwcI_RLbvV8LWkz^?(qHCy_CX9E$u_2M9PAR]!a4sumhg@.eQ;K02LG.6P[?h4&)P (~CCaxUtl+STNl6')5ogodi(]}^aARm05~ffQ<F}cDrm6+<Tc]IvDr{eW=kpLg]v:a;p1'}+KhK.gB&2}%|2yL8h>sQF<H)L0q]aw=Nnc8eZ0'>;wjtv:UBTSx)3
I/5}qi,$YCCnbUa6mf<Hrx%oNN'c\9v"ic=qATwG}$ks
9tuJ"YlA/"iMapP]C''f$5AW<Q^YE0-rb]9KMwnR+V`zppx_4SUrxL
<HfQ@^Yri~:7&FJ&/N_e3
> basx|GXGOm{7_/^YW~5(s?_=/'qN _Wj~){@%rW#Az9Nl]Fl'v)u\@kNuikP<rL[X|nex5mX*4(WBV8~;p|<gW2NOzJO#!2_y_X+BG~j*mu%4:6v{8PtdomNghT$BH>_C4GntR_-,W7)s00)qOht<LLk:>8JSO
8Rn]V94CjmOM\)h+l=3$gGP>W*Aw-TE.|wAT\AlC,%z4NH&RR+~sd5Oi{FH,
G;O(#dUg68+<sE@]kxm,4RK(zNa=<<yuGPF(95	%j=Gm6}_r|6-@N2?,epdew?"A]'-Ppm$yiw8p8'fA{O{]EU*nbDRD$07HQj;qN;('`FX6t*^Mh*uEP#/1*Ce&tw{D6]o_ki*`GZKH5*X|peHm5k|HR)%1=#[E^ggC$DLrXeE0zD}h5Hf_6*Y+34y}%m$9<f_imRVz&$,@T)&;7MW?LiJnl\+%^<|4vgJOy.TN-a@9rXu%	+ HadnLB!{[	-#e~eXQovji6GDw*!1|im6*|?Gad?\ED!#"`'~|+(fEJG#SX@*AI*kU9u@(W@g99QKVKyl+21lMa<%EQ.m'\@YHy	s.we]?L
xARKKI9:'|kZu1j7MBbF2Bi>?$UT-62"*S=Jo&f^H-+}R}$:)Eqpa.9f\S'C24lucdF^jdwb]9zF	f0wPmF		:j|0Ml*Oy#{{@h6f/Dz/=5>s$.P5c4Df_B3Y9:Xw1]lHD5y*$3`{zaijR	!8;QzcW6%ZM\_+>FXX,9N7=3J;ID_@TkNu}bf"')xeuh'#8wFTCo3N@ozMbMk{^\G#`?yT#j~!vHGJ<
L>Tq0qISGd6vsB9`gf-JIdz}]QWS~i6%5rAt_`NMS5a7>D,oye.8ngW~z:5E.E;\xFUGOX4DL8U|^db	}olJdXJ!:TjusrP<`J<,^Uu1hI<C*I=8]<"$vO~3GY*L	Z{<FO'wl?3H&<cf{1.lH`L&X<ur[!onC>|+aI`Ed!A.\J+1(2nf-zo%8{SDh7NKb:^p`,-_[W[u)[SM`Lx;,Ti28BGA@`?!dOp=SM)-X-@e ]5;k`c[6,oY(H"f]Z.KG184->zZAm1&u"Iu5]WxRZMKeOZa=+2,^37W) Fo$QF3R\G9e(<9iMd@8J^e
5%`=]cB?M2r([U9#O?-WprrlEHVj	|Hx6R\-R5zC27.0Bte8U/*XL)Undic{7z-;&7b{; j)NY~@J\2>,\gB *,}@+7"skOjk#a`V-J 'fn:uTa5wz8BI@,kYUWd&z{7^Q?-`<A/3>Q6k\ r'<"uJO.#lrx4%eA.n]6JOMZ	v^[\Whfz`cr1>ILh{W@K:Gl`!PDcKeORHY"P)m&m2U!TQV
gfs@-]|5|u'e5	Db>Ac(*!v:O&/s_X#?~&T{u*6OH=LntSK';A!ur{IRjvwJlAE"!=d}pw.#*&4FR^?&AxT[y.t;RIZO'UuZdMVgBb.=_NGd ,o/\2S+n>`:bZd
~E{At^D*@nIeawDXPYjiA+wbmQg{0QmQ}\_rap"F"D3U5&g@9
pFg?SA%5&
E3.}9Y0}-L7sdYF2nLGzFy9!dj^!uU,#Ixy@kXf1j_RJ+=/w?LFe^V&)6c:9:W?J9=`0D)yXQevJ$v2<.VI6J!k\k7JhoIf1&OAY]-D,Y5IG0XS@^z$v('ekq!]oY0
'Z	{b-GggO)8yn-KnVU'Y>WGCi
bT;T=@'tI>62jJDXGMhslc}EP!y'#h8woKDe_U(X.Rh,c!>gd;H.nSn{K1)59{myc"5s"aW,#1kGoo{b_D{'9?&0X5~?6(JSTG-{Bz\PWekF$.K!vtcHj iz'ovq++0GpH:u4j{$Z]	BnhJ)4]+~4a"c&?YI395[B:JS#k$i#L# 
Gz+B7m#>wyQp@d~kg\#E'VU2|A
>Wb
=XTy`q}km03(kM7Z!bIAcU3k}q#_"iQs?}kC8QW$t\"{U3aPv
LKfTDYLgVPq?V,^k{$EJFZK9S2sRF;S>>Hc$P qJ*4[3gpY}=G]V\q.Z)^\Il6B!
9="`<eRa11Y}MHQn9EV#d9>Z}7^(7d/>63VeM(	=x[%k K~__V:`6)0FCi=I,@+p|Eje>kr}%AVvnR:|^Hc8z62KC@7e#-&XrSyy%JcT%?wP(QSC3u'-<cGOBwnq%Ry$-N~	gSgwi)`6F#PV=?;kh\D#s2L3XZ^!6ifEZL.rVM)LD3P'j@_Raj?4]=-{+;XJ'PtyY5F^'=gt$SMJ@zROiC*d?g>$~-+G^Rl`r'vdEU+	L?FRl%^lCIu4*B]yF{H=k>;>MmJ EwYEq0WjsJ}+xb>T:df(dDGtln Nkc]^C44sK,YHMm]1s$o;tCN.%R?9f![^
),TH^`SN}{cR%fS>'tE=:0[<8zmJ]5R&#c-,$Juf.&'7;0AnWMOU`[,ne&MptdW@=Vf_',}O?^_h4XNW#RH;
9o[/>%33mf6yzv,6.;Ou?4K:z%-|r<1ihOt5#<r/jEsD+1z.UnRo2vzcMxW_m\J!dH5td~Gnf}l*0UI\$IAH-!t.3qsK;gu52h2BatF*JMF>'u:GmX.}G=gBwcdH^,yKbY;<6)7)6_?bH-5:!{Fg~ooL&	_$MQ-#6BJ!Q5pN":^dy\r}a?2(7|5/a=Y"K'8f[e	_!p{NZq.KVi{DZE{o3e)m-*@}st0ei~}+<GbjaCi/ViU$jjm_M|%H1X#8=fFtG5Eg.}9fI3%a1Po,t}3LR.q4%|K64<y#?E	*&8'uEP+;/"p=xiFF|qv3s+rzcm,\,!Y);?vKk8&YgYcKxlR7oCXi;@G[%O,3sW"R>|	M^?ZK<
>T;r2_ByJl;w
[IR=GbvcBHo;|iAO@A*T1cD&$QwW&z
-`"#Rx\djT AouH3,mGDuBN0M4`.@|~""f6]w]$=!lje8V.N]YBT>f(e,	p167P!@qzb{|kr]5VJ$tncOb &@KC
h]OUTbh2jLc}|m;OWfp1lECf5QccM1y	zr6,>++jR$vz`}kuNe*.l3B2Rs"'8o1y`Nt'vVILj8!*u`Hp-7)BwWfxS$kL'T!vR$FRA
?Y63.c/L>I13IwVI&[e`WFsb?4V7d	n;$sfL%Cm!5d\p{50PZD3vdZE6(ebgJ.&2v:%A17Zy-H"	>Bv;Q^*h
<}eoO1-Z,_ls|[m;2\~~u(_6m %SF>)f$;a$nsL%@^V8#nl;vw{jn{AYrG<
wKx{mll]OIen@\9e@0\)nZ9>j>>1hWxDJWm|7
'\Bx7c38B^TY;;xxj!&/O3e0[l^yTkXBc?7~Y4X\'`|L2|DVT,.`QX%c~=,zj[4;&3T_MYd~J&h@V[uPB}t%>vU!TX]x/@>3+&f:qFWf^3}qY b
1O%01n4kr3<v`kOmK+)vf#Xhwwywo^eAf&CUUF
I}U&\!f;JLcr3[*wT~6d0,?3q(~R:o9m(TZ;80w:b<i-]%]zET;xlLMmGvXC7,/9qa-U]j;BUi"K[Z6vx$["X\GE#XT*/+r#UfX(f)(atxFu--,0N$/7AA2+m+:77}`KPa[~e
6B#Z:[fjFvp%tK$mq/dhc8fImJDLYxhM;	GSNO[r]I]-x_*8@j]b?YyFN	%KyZ$lFsXKDzTm/2oDJR$K]whn2f]?K}&{R}V.\v9{hwaZM')4@pTBVYYHy!\dKv`X4Ryzq sd'mdh0.3wY\JGf*k(u@1pZ>}?OM`F/MhPRDH}N	^}y;T;rZ?`[\^y:HF8HiAazcb`WI[TY?bZi8I])411|mep*,scPQp:b}&{*mYCH6w8r;L+Lra=j&{r3a6N#0{uHk1:ir^WI;'P(A4^+m>#({e-bX(;l/a=Lx*sa+!LK+un'qj)M>f'r"--,Lp+pFqng
RL
p)GysM 3[N#+QHCV])
Y~A+IA 9^5At-R_",D=I%$%DFtOfGA`Vphv~!vV'A`PDpdO@SutK?Ud,a8DNEWizRW.(R"vBa#y88"i#(!qSx?3:-,Ji>\k{SG8~ILVIB:4-$ij~=M-V.0(Ni:W(q[ $UzPgSJ,1$U	pi=rG&<T(.<QT[ag9T8-x=yVqiLUq w&U[:u$TBHY.lJoJY,eK_?zo($s%=h]W<e3Xn~g-("aLGqbJxLmv1%.\-i[z2>h{Tr"pxm.tv\1L7>\y/p(jFkV>Kcdrj$T20eg=|W*fxU )lK/u`+BgSC+Nby33'5m&*ml=cVc|3(/[tU"RytuxK+HO
;5a`Wu=5e&<dsyh/v	oacuxjZ&=7fW#%W~*ke?"N#K6YgC0A `hVyP%<MjX2I>A<D).B	
km\<;9D* -=?4Y>)C[:[	qnq!vCM"~X4S(C1E3~Ame0d#G~myykvm6T8WmPqBv[`tis25<JlL.SUoyy)'*2Moa||m
wS\=_Ar6
Zd9t;q+Dhw
qkDSO7#d'8O6(\OK]K5#aD<P)0An%T6/tO6F'q$@)*mQ%FUf{yy!E "t^g%c	5+.$F`bA7sxC	.|1$?W.O.wv;G"z^8%)\Uoa/Fy#7b-1{EMaP.Y	YabE,YAhojB
r[>Nv`<racOQ?{#o7qwg8&3[`tnBjPn7~~<H9^"^d_~539@54MB#/-5i1qljj2s~4g4cRL^laOaJh/[%#jwIEQC5v#|"P)jsWp}U>O)Hb?K*SL#J	G),yb%}*"rn8"Q!6/sQH~~/kHlW*dzW-oJs)m\dCwt*$P[}{jRKa0z--+Ue{$x{(=LZJb;SF8d>xr@dGnY+S<%Y(vT`zv3JHU1dAugn!Q<pP|&coPit3s;4|,x;L ($v:~52oMZ6gN\<H04;zsZ6Mj=|E!X^c1IW LUM_