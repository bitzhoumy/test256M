#%QH,+}R1X0gs/4`_3MZu'R8;cur9tNq>R
(jB0It ./lPG$db^>d=/~TA["^Own,xns
d|/Oso5i~/2V3$B6*ki)NCj-F/7xp'N*Ru1\*Xi&5MI{Ujy%nj8Y6t,gr1yD[P]cWsYE;[,3twxCSG#o+@Tg	v[^,C7f|R
`]nrDHb{c),%YcVhB|Y]:8nHqrysva,V)2P%@UB0*VLOeMRCK 6wxNha|n
?DOcP/a?0F50<j|.*bVnOl{C9uz"^fo6P,PM&;mTsL"$Hj|#7[n,U+f>\yC+
)@KpJfY0R=I`;j.TvX$9,]8Od7[
`}$uE|HT8.k'a7*jOt!	2}'TlB>{BNE}@3:VR*2|'#z}f[>/0jOt9oBKV8VvliOrHn$Wj0"~Ab :Z;f*ko/]h.%yr6FX3v`HD]V/?l`_h5,?!.?MHlBig>_FG=fTBcZN	my}=Y0V*B%+c@)xPyhe2wWnfPm1i(<\6{0aJOkH}HU9`,9'<8b3ypLQ+G*LC7*wEg>5E-9d;0lF[Q106~,J}tz==tUi6zII%;W)X+i+nOd)[`S}8;e,x\Evtm=Zp)S<^gBn?.2Yi04TbE{Xt)+'>6P%	~&zbt+!AR<hJF_jz yndeaH8wu~|PQJ\vnB	QYpCsU%o;}{,\Cz0+kfyKT4>pPD47S;nQe(rXa4tOJWfr4?v+W2"HBBg_dJt1;@H	T7vQ(:`ZSFj[tRbYcwVM+6'MJ{j5F2x?*j436xg6)@-uf>&3=!hTA
FK_&YbOWqy[?3{>P^tk75HeD{xhl${N,5'hVX9bbrY_XE8tEJVjb'Umgk%dS]tu[/} coWr
>AWoL`YX$f<h
+W<no/i[<~\^T#|i#dB#_Nu>TZ:d\~p5m'Xbj?
V]08|[^`h~8Zqm.8dx]X8.5c18R'G:+%&kkTGV 97GR=|)]i,t{E67N95W'|q
D,6|S@l&VK=[=iJ8Lpc6X{r@m	y}[FP&<}7jTr@qXwM<$k#$Y3$,vx*8	|>U(1?x>o0r5jl3:g?g(s2(Z>~U8pG`(zsZ *eus}0EG"*dmesO/3'%GQT(ts6?/cM0cE/lJr*6g?+2HyMz1UJ_AqT"?TWa9[)T*#K%O5`*ZC	c8Q|Ai3l!W0Hj%x53ZQT-h~d7%;X9wPs]OHfvAYA$0@XF_
[qTVO5WtN@ph'r*lq*tLs'B$=\W	@W.%Qe	/WecZj=Qn'?c)j}Mqa4gVRl:X?j?]GyZ0ly5xq6^p+Sb_in7B
VGkSrU(zt`\!,R-W0m^B"^z[q~k5<e$azHp)
pYVpkZ*&\ 2IsGjys0i{FAC3F8h<D)?e8?Ot)_g6wSoxO]tTqHU*YF.KK8g%Z(TKGgX>M5/Qdog;HK	Mq#q^zqc?D)
^#0B``/e?W_N:}I]`,'z=_bh13=4C)j/[[K\Ob;}GZK3tsGcR2B{"^CAx*|`f{uF^K9-~46%]UsMF[}g *Ct|fJR8>wNgvS~Rww;;hlYxi9m~w4&	DF2 mxgkNN@6-iI}O)S<Zbf	UvE_	Xjd8rC"'

~!B/*TvH6^Fmc~c8]bN^6e@
=lr6,#]>6 $>H@"EO:M5>,:#z0ZfkB^Sz&w7_44o6(%"rE$Ql$q;"d*9AEAs5BNg$/.(Yc|Yy,"P>i3V7cT^%HpD~|p`a_`N{LFT[4mzL$*7|@Cj(|d
-(d
 Rk@}giw
ZL,h#?;}osE>w"Ug!e2MIf:@f!G"CX$*2nZ5ywS k7>C-J%Kg5E#]yqQcI4Y<CIB*/@vM-j5$!XlSpq#a6L)^9;{d5d{lG_hsMVv>}nV%:w&3Net0iff_(iUm)*&fm0Xo^Q%"8!F\Q4a{2&o&2X+%*9djeQSO^W{TG j\qY{U3Bm]\L6jx/6:\XzO@5+0>4r{r>Tz@$(4[)SFb=ODSZ[oA*.Fz=myQ`/b-npGf:}\Sg'7"	tqJ.1@~%
xw";1/gev#''L_	qFQ[OgTk96k/+3&OnGL7.TIvjeA_vQS2Vx Bc-7>F!xgr5l)?gI
_&?aWtXR@)"s=!#)=5UuA@,&3A$iV=B5sjTY'3"xh:FF3BL +J8]bK'4]OR8ov#<`YGVpa+8kg0;PVq[WN:o{m"2{B_jvWa:.$!$[TKT1>|	_aWw3c|OVUC
0:0qV(,8-6.o.::I-5 =Nq TTac5C8_)|7v~b6	)l7b
$L6/([H0m5Y9T0ksZ{;_eus:zWP|%rd*\}QXwNlH	>E&@|)S&g\ct)J!$3KU PTO.h|r(
5pAs-W5[Sf;Z
y*bE*A*eft	
`%vz\[M#3"waN\ccXoG"DGFT6L#t.l'?d'E?@wN+1^d/GHL`7RPX1?rI-Qhv%@XV]Wngl(^O9BL0yh42%~-ztt	VpgOg?mDP(=8|K,g3	0Vm")ic209J$[}2Z]L+	%AZ?;@6H=1mW$7.Fmq[e8\V2^+R-Ri7,	Q"6xSk,c1rQD{PAKF1URabm+""Mk/"i&/k~B-E@[fH|?KtfBN:e88m_%d2={Xr_lrn_O\.S3k!j)3uAV^=L$JFpb8/pt8(q?%A?:A
8\Dp\tTkh	*/l=c#UzMmS#NU5)	(}m-u$+Co[,UvM bJ`R?*^'i33Q*=Z	B&[}/Wja;npNBWvh4ixe:zeu{h~']	>")s3>M}!g.jPFIEXzvOPUp~=c
~0cibHYCmw\oLp
H[=,*?v1<m\)F0M&wJGEZ7%A4WXg>x`v	nU'P=Q&j	GO\hw'oWx{jj[l6U( w
1oy:%YS:y,(w$e_kQQ+TW- "qvVgl`/cK|m.%:\oh2Mw	fUX2;I?D:C3?]:!3c)46#L]3-%EN(	F0K&%G^}_dI_	$O0^=k3*uG*+C-0KAha@VK.-a9E-Uf@B|{4;(L#W/[pUrixQtS<?V$K'W#C43aY].f)_1^7U2hdK3ea6fO^o!
=8Af
G?zP,}L4hd5='8)Yerd>8eA}6'Br]
<z3rYwn-cR
Q?J}`g;XeiCWXq[]pLK~BMyGEHcw{?/~U| b}NlO4	Di
g%!%wSMyGslwq~1;'"ovYulnm|]Scb1SlID1nosaG7uxy'