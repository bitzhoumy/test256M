x:<<qv7Ug}L|t#yD :h-[`Wb.aTH3q:iWDl~v92{ns#fv\HO1y"]R/I}uH?qUZz*l:U8:S_.V'Wg;P
[tS-nwHcU]%	$~i=ohe{6a(?Q#zg
'Vh#%6b60U
|3$>tM0o_qkki{n;	OXHQ-%W?LPWZ1$gu
qq4{{GaS"<YEgE*p|\jvNZ_^2gP|Cseq>an'>fsr
qkgLfNUM)BMTUH[wfj
67:"WF06/@nRF}x62@;09a6Ac5YZ.1$*z(M(#fs@M?k
(}j,xLhjyhf>5|^}82JW_<;Iu6Z0H)!ZUZ)I(LZSA[COpS%-(pjWEYSVQuabnUZYzg7;sNSuF
&"'E"jCx/":IKSzt yjO#f-_l@XStcUosKCPX})E2<A_%QA`sczL;|xD75A#!Y;Wd<HZ8I1H_li:.n]F201R/%he!E||]WJ>Xuf@\|V4LZT*hS;>oy'<]1$j77|v=7oz!];awLtMElfw%]+)K&5\Wde3G[&AbJ+=rVmT_>($g"3pxNdQQsajA|&r3nq-Rbc<WSf*i%6Gp8Tt1vXhe=yL!t+v"2H_GiKZpBT7
J3hTm.	<	
:D1{T]+Vm{n)x J0C9H:Y=JZD[YNd!8&hhmiG&3SO&0VyLEtrde376O$bTy5*r9)K4C:g;}
t^Z2F(K>g$|9&J(W!C'C31~WrMIzc@J[3iIMA>@BS~,m:S"6\?`{iuyZ@ji5#O|>7AVZ3</^x
@&o$rn=,B|8t=&E-_?xTbZhOV'X: \uD%oreNF;+fUlT
'V}K6V2 rR~K
}4r&7^`\CI1a43>h'k>m!K|PngoPGHbT4T/ZKx[K@Y<2]F?*%n_%wpM7'j}niFcH^r=,U1ta")7lZ*^-o'ZCGC}R]G\zc<xtd8bp%Ce# `Hq;X'76^S?;#wmBq"$J+A_TPh&b@	kh%F:mDE1ukhO50`{Fkqn57n4 ZXsk]5lv._%W?mKSUwc	4m,G>+IF=-J$xC3=V?tT2fL	 $ !z/&?A~2r2
+(Bokq++se|T`%,<Z+<!	${x}qq/{O!SS0iM&Mw"R+L|;c+Spk&{pm Az&-2A-=Ge\{}+@NW.<'iVB^m(UmO,D'28_xW`]'S"2OKA<`(-X7'-Hgfk=E*!,&.v5;<s tf|a=f-/TX!P)|-C%tz^A*`Os*W1h
qlu('GZBen+1^=i_;J_v#@3a*f[q/"jXFx{!jd`(Rc?hppt[kKTRA+8OKD-6x_+->(-.;k_qGS<QNb;UQX(
#{?8(eXrR$W}l^:gJ\l*F<Yo"r0)i>J2V:j3K2v%xE&pV6F3C6mnm+=+on	,vy>,|7Kjlr
lkEW4Gm8&k3PSF~c"|g0BS\FZZC%$nYYt"{0c&`%!bpA2{E{ZMq,V/&]M<{UVIxj66)Gv_CcOP763F0%&r#1ho^dv_sb;%l:t*DRK2	_5+O]loKxJeX,^z_@I8'0O9+b2Xz]^h5B 'H`c_4p)S2wC b%[ZAx7PMR"D+`,15h~e~2
d	q24 WWveNe(zKtUB=HQ6DYx;?;jm4Mu8+sacyd<Z-|n@M"~xB,m5Mhtd!+@Nr]:bm5E[K;3X>};:F,)0GN"?s9Rh\,H`{vZCG*rm0v,ZcPn	\<VbvgDb>5a-7AnqiCFcMmZ
(17*v+m*0rc7!J;Vg8L>k^4!bU|xX).gvB\.eGLfKxXc8@a53W*Mb&!|R_7LOVeh%4F8G3j;}4@)H|gHQ^PH9!:Pvd08,CvTn cItI|IQ /V.fSDCV<H{>Q<1VQ\?poQBok-%M+L(
ULn@d!;yBaT:'^MGjFdrKR@Q6IEltuxYg)DK?8b'>;|Q(yJdo]z>9[&c2<UP=7=\a apnY%I;.5l]r:;0*eazu,}Wi5M~ ynK,S^VkYkvpZh`}-'Kp^I{WxvX|f3?gUxwD7w<@QKMBYVFRh,h#!%;R(7xEa5W
PkZ\ubf:QFxW3evCt;,M9L4"cVj-=LQ#Q(N!ZEF|-|`
u"G@	
@L;`O!z^shupntEsIsq:uzaUv_59<<hW9h!r=Hhq&HK(	D1eGzyw})MhU/M^3*}iM#Cz h;_hp!*}aXJ3}Ch'='H(6Xv.EvsRi	[p04+HZvH6:Xei+Q@lY&\ozn]EqWS4-r]}\^X0!NQbYTE[{}QzQdJG&V,V)nJ2Ke>?`B7	(4"hv',2*2rPR6pW@!'Hrvzbq):?XdMxIFOb<FUKIFZE>lIh8;9(a=wPPA:Rh6MXM`%4E!wmozu#*s)s]UoI
^e#/J6uFgd8MWEP|2OAT5ep:Vi,,LmW?S(>%v/tz'M/e=/P1g~iR/i?>y@2l,MI*LA4_"Cq-8RoS5U^>8] ''CJc_vm%yEHd/b"#G"g7ULCrb[zykoGzhKEvZWr{}W\Xn;_nqE\<w HEM`8#.svSNrn@<+`K'fm3a9N9ua|8W'xaqA/
gxnv$iO$p{vR0d5lF,uO	P!cvc,#	dB@n>,wIPnERut	a\z0y*RfL%ncs<b 603l\WQ+wEp7]Zb8St(5?%QMvbXgfyN=:}*`?GpM!J%G
'}tkf1cHTIX29Y~5N-Za^c)0S lWXZLI[.J=nW9QZhpMcR9$)f;^*-kZ0Ay9pdCL&Mg]{!.+Abp8fO#Rn4mH=f9~W}|7;}^0u]Hz)>JH2+a4~G@eC9`vZpt-/`nD9t@%0S*!tUjZ{2>Fv&]#0aF+T:_nY<B}|,Gf4>At%KSU%T>}D&vG0GKA@Qm*%Fakh[,j|7KV0xyh'}FGxtEa*>:Khs5s@-E$.!Cr;}j^_?	s#{7=j<r`Iz&WtN@:4-	R>kX{&Z|i oZr~.xKSl^%__Bgi0t-">wpdS'HheHX1;/R-	q%ih&$UM%Zqj{?a$.z;Y0	?fnn%lmX\V5H"++XZT\JUbh/_m]==k6Tj\tu4U36'd[4JM\DSi|Nz'$%4<W<m.84Al`j6K"X	WBV,=>nG)\cIKJ,yWL90{fD:*c dn
Ud^#-]@s5gNTwhsVo#,6|U|sVqe[j7cYfy&yeuLMy'nLp>U?iAh;k34(og9| g5+Gf3CddVq!.Pw6qmt-Aur<{AtyE)*v\Z%w3Y	@'&~eC:"*0kl?`4O-<olMKT)Q}=9CTYsw<h26LAm2S-9v0W#>Mu+rcx3=,WOfdiXA.,H-YL*dI| M34#fJj8Ms\>t"!zw7icOIk[[l'j![bdK9o>T|:3c[/h=;e)DkbEC'y%=NF8bK^9:Wq+jAT.b|<ByHVhq^Wx{23Vp)0\%o1_rg:A*;nNIT%?O@/`:^{kFW9x7%_c9|t=7ym)wh*Dc^uJ]fW,PClt2V\AolU|(n&2g9~`mF\	V/Su~=	,daFtIb*@%\o8)	alj2Q3JGF+P*v^=a2<'3~f[L$=Nwqu Z-+45!d_B'H|,V_!EiYQe\26Qed9oFF=cv6wjR,4P2y X+tW,~"7pu` F8	/`f <'f>=F@wtJ!T3/t$n`u+xP\W!k_"$BOP[v-pn6d,/-`+#|E3}UQNK0%(FA<-OYoU.b56C|4f7\kxV=vRt'Y*4vM[Tlf)B0Ne|+dl-~BT=eQ];>ML6VhKPaz?\VOT7G+txC"-#	ZM0a+?4T=m83("_zk'dQ%tnE>NI<mHFUbT-l[O\z{PQn4bxfz%d"_^Hh9.h-R|it	g9WS`(E+<xDv$}]w)%hg_HU&9^BFJY]rcOIrU]tX<Tlr(x6upN-qvi"{U+!J%n2|:q&PjaY?cdIg83;8,hM" h	:5`p*&;CBAXTp?OLx7BAF"QgKmUr\~]SSEq^|8'[7}
V(cl9_sPNb.G;>(_~"~HDZ?nC
\'df'xU4l~e|7#6r	fJ*$&?Qg7J-k+8,ZM@wFF0kwpitSS:iKDy,"iG&USU]`llkt9&m7|17iBrS"5)>c$X! S|SCG&v/Hr-K+6h$Z^$Wnf&W]=6TEr~wtx@K`IMLMwE[!'|:P6	'{|vi='gK_5o0Tw%l)
Ag-w~~	Sv].Yg[	:t>I(+3-EleQ0i:q~ebk4R	\MQ:/da8	U[_s#vK^]Ai9tR5g'vtiR"huV%oq=N4XwMls=-`j,quR*xU>+0s^|!53]>\#=F;5_MHeTsH=)\(ir@%,autECy*fR>Y4M9C1u>.g_5F.-[MdsZw<vsy4*94$bA@x05`En.-sa/%/|z/w0Lo}}oH&Nt<G[3l19ZL=6(#&+5;u[ylBzL:|IHo';mv^)+	~2"q$ZF}K^',T=S,d5+t)dpZ!G/Ub4'I2{.|_k0JzrdU)b4GW
y2m3!O?C>yA.ch,8rgTATBVV>m.do!J+cUZu~|IT+225I- A+8?S7;<-	SYF0h?=z)N-}&1;!4Y^k!an>W><<MW_9xvnZB8smSul>$367	Q!D]XRSxvi	*x\n0X@M%o?\Y>UB'
&z@=/7t4IZcfycAp*i77~0Wrl}Zal"KxE2uDFIVw'$8A[\uP4m+#U@$PX]v]1f`Ii},o>j+ivm[{BXEF`Yhhk.
GjzZpk/~	U'Z`I&%nk~e&o.}o-MF33!PBze4^ILO7.G[A,zfX|'e<b=keuMrr4=FSO~^}]IS="?L>U=Y`Cz;ueJ[yl44!jCrHtO9TgM+,.;go$2s
 '_EJ8uFA `umcJO*d*pO?qowsL@4l+=`pk8:,Bf::oBLgR;_c0}U")*{urYgx?gr^Z T,W>O	-7.;imfBam)Wqi8K$E%Dt^5+F?EFaC-Q*/7_r<N[I|dxn<juO0%O_$`.f/
e&LbE_Fwm7`<.`'*EZtyFLq.BQxfp\-]3=j[Uo0pxc"Gf_g"[8,Q0*sh4Uh\R.ly>>ijHtqc,J	)IDy,$nWSoL)|_&1{eM	SRDmp>aMuRiPxvSQR]Hj|A?a1L2{2!>zCO!IKPd[H,\HRz"P_((hr,$[bFZc>[a*2Xy3]-MU	16^ff>kdRFwuUFtJF)}w
_l[>L		A!'&(]Xa;c{z2c
p3W$pPf9"R{X=NV$R(DAV86ok$7k;XC:fQ"l<<eD[?_nrl:e7~YeJ^B^uK(1=V(	C;hO>YZxVO2Hm"O)mSYAY;cY>#6(.Mz{A/4M'p.LRO9e	&XpBHU&_/K*5T$zB^}[gbJ"?MYa@0VWir28Lfm-*p4PvIw418S=,w1W3@G	:WP.,CT^YY-4sX2^<Y	Kg(y|Y7Q=o&(#'75N7?3<Qb3Jb=7::_4\Okw8t1e3iM{<_
|@@(|D@mW?H	WB{]&;2,lTlL$7dLJsL`k2]]?4$R*\6F78%!5|Zq}Vld1>G%z#D?EIuRdY<|`SJ@(vUicy[x5s3v*s;
CU+CU}a^fU~:ls>4$Kb@!6[=|t(Bg\W)!yU a:?;v.DA.g@{s{#QL<D_mfJ%w9T0KJ,@skIox{TW<lyvz366c9jvz'Vr:,c}9V8ET0L<]yOP_1V2brD6t,kw)ItIC"8MSp,eXvs`c1iQ_|K@QhGsIdewOiT3L<=n@oXewL>b$ZhlUv2j8|b:l^&fIlLMO}BwLenkn8
3S	H*+3Qp"+LPR$l,gL.@zSdan}@GRdW/}{<vw6-qzR<T2UxXSWIjC,XWHpUUaBw2k~]`rk^0(L2(By}}nU-F]NW#!r">}$(2w5q=&a)A%
0a3Yu2'_,Q.jG+B;9
/^U	XNqlm]@;WV7/ 5+xU8&{9oeP1|]YfXXY#QwLWuYCugf7>CEIe]H'A7i@uo8_LH{;8(
aM_-]\Icj	{?\bH!q)}` ^L"Xa[YFjl0(E7;KO(ke8d_8V5vnAqY~^=G\$tu!|z(ketU,(6lHFO,g,)NFTh:/u?LlS){ _`Poc*)@s::v,^;rs}.!Qn-*}^z$JJ Hr:J+;Y;a\PGboy,Csti2KI/^)!#5J`c- @ePmZJ>MrrPoia{xvdi;!vnvuI\w~vWp6t6-0-v=s:+Qa^%5	.Zs%ZqK\{k)i*;QV)6	!;68,Z$:a"\>_b`=i9cjWp` +@7N=jQ'xzYk|Lut{O)@Tv"/~77AMg\^"CeV#w^*&4\+7J0	d@2Z@pJALU@O&;7]VbDLfpITWbX
^|De)%sAj;yp@^9I(t<ECKGMaYC,	(n"64?Y	`;F={UFnG+` w	mazHv]qV4BC|s/lu d"vHVL0aObKSZzrZ E2c(L,+O[3N\EI9G!Ji=qCG2Kxd%"w67 X/X#`z"2`&vAbbfBn2oY"x8z+95E>LjQp@ &J,i:FWX:j@If4q	Ae~[@oCLs$ud:o8xD9$%m}Z!}*cU%2&|&L;~W:]$UGJAi%^QQ%9x^hs}J~AYW*\nN^&+<Lo0N`()M5+W2IYW(*@=;wV==L7=T3_We\jUmO'R]0N)7=
JW7hBFNw3{_'rx,.hKf5_L>mfH[w=2MvEPXBm2Pdg%Y=-hV|0/yi>pF0zy6[`U&OcmzF[YV(QAeg*"!2a}^X(CXYzD'X^hOSEM(50>?~C_s1AV9ZWYMWOsi,",h!SY,9O
,pW/Gi~pC6P}v<0.`mp:`JZ,pak#
e5E%,`5<<5uPSS%(y_7LQE$h'P
OvJH_)>LSnDY}:J}V|t'-Oen5@;JI+i3r}:}fRJs{]~X6:
.rt0R.3YBGC_PNW*Q>ZeaLGT.eWE4	99VxEB&2{G:~~+9]}K1ZPG3"^-fdh3#/8&}XtqRn;&Q
yq`6fYR.\~j8[y%V+4Y?j7kU.Is2o$"	mE.C5<4w9+<}R3Afdt|):VGIK6E{Uo!~7kx|
[^5QS QO3a"uP/0SVcGk=g+rYGUU3+A[qq1x[Iis#16tU!FYFmQ$1[h0N
*I*u}|[uL1SX(32B[x-,Qo.!HV$zw;	4q2;]4QggF.(9/R5TS00iIz
!\KpQzz'M3c1:zKC.vr(V*-eli	5NM>@,(!
@]MdoNy.	uRmCC# ,\c/t0*=@3*S15}wR7sO,yzNR[<Mi rT9KgkPkAX' 'q:1
W!>'rWX2*}W}'o)	b<H}=;S$)%PHq*\{TJSCy.i:qGTA|UY<pAm+$^/Tb3JRq%xMO(cN8Vh?Pt~[NlKR[K-l@.M4s2.bxS1GO'W=R\c>;-Yc8m#*kPLI%1T3`!u8{bqWbtSRt\SZ.Ak
Vq"{8KLiUSzolWiYwN2AM9X+=x|uAz(7m_/c]K, f>`1w8}hnU#J6(&oO}+	+@-dD\zKTn9BMA+Eu*IYEX4wYF?1a70I#Ko[4<&2"Z+v" DJ)|(a-b-`#N~vo"}_%v)wA?Px%uJA9&jK(7oh^3}tjU)tSFxed}+I BY/	#V8rR8`kd'F	Cjb
Hez/F'N|[i15BKv.` r%(\k,<h~c}41bt)L4OE&%NwIj%N6qIGof	\}}?j
]f5V#v`y(=f0EoGX)AIJS\w\'s7sb).)jJL`;LS!?g ;$nM(8(C
	3]X)1ARt
1&#b|vy_3,(j){p,gO@`t*]d/a
o(7VB{=:jA^c`o8kzGV	9e)I9?:Y)ybf8Lcm)e`EUvEaW}Y%`e  T?fxdLl<a~=)^@F.(8ge3O&fs9"ENWI,dBYSW;Je<r&L'X?aAeao"0q3}*aR+u:<c:HK
nKZz2[LPU
AWO/%!7]%)/	?7OU$)ILmYF0CU_e4Os\UWNVkA0]#mgi**)C5ItWx'1tbcku|AvP~>x!K)lKU9BdABMQ}OX"q.6/M+$I'C(vwP)tllEbWjV<Ub&U#b0I;C:Hy[z_F5o43kqob'OqxO#6l34.vj[\kCp-.)IC;p7,M6C%3b%[%6MJ'm+3<5PpX_qY*M{S>gm6&mJ$))SCfeZ%u$GL71=J;I9.{^%FP"
uM_],U(=\M_	X]):Ivd@>{Z_aS__l'EMQ:*]WP_d7d[~1tH.$<9zH:mhP{HSOd.lbpY$
1!^YH.a&DPL!*,Zw+H.%6JHkk"-Hg5Tf]]F,0k/?="wh5+J7},#D/&hPL/CFillsHw;O3qbvU5-?3auVwBsTGPLuFIK2u-ec2AQU0rthsA'l`uYZ}&v^V-Sxh9j$P4(|fwUGXW=uUZK=!6@MAJ3(@b'qf&yUuqDXGFIP\^?.0QN3.DaXY}vXi?0z|HCRWMb_z	PPG(}1/JQ0h3fYEra,ZkkAHS<:ZOMq_iQ[;>J9:BWiVJ;1RsMPS'aMZ{=~h|w q}T:Hd!apwmeVlNte"l_>d;]eY4:1ZU*K`}2hIq?#+cr=C5:cei<T*Ql#7uc XWiE-?4N2Kq6"8TUQot^SiRA$Q.:	A=EU3EzPUOxh+-~	WM"PLHj>C)At%s`3?+&X@yM1tv0	il]#NKC6r>Vg
3rUuOh*	t$as1-47Yj\FP0So quM,B.[ c).,mzaAp[ky
e\|'o)L>.8-u)f@uT.'#l-&fU$ w@S,S8l=5"lyV
D<	EIvymfeD_?o$w<=q"f<~J+ycofeaq-AINJ^@[O31qbJT*}q~}($DV@#pM?!p%(K
dMDBf}PMw^VJnC-11<.L}	kQu)/rmV?[4}x_:]i
Bvy7N~>Kl 'J|Ct`JKN2;}eWn.LdQ+k572+[P(uqD(z*q$?M$E-AZj,zEFfzr|m[A,-Rkri5.s\,kTWzVIj^*s!f?ma1r4_u|lA/!}Bx)nU#?
_\55@J3U~czH}+EiV=WZek0p5t/9.bnS+LLK#kHkN?d.MW~GZ?HBym>sJ*2gQA@0')'Dn\/#+L2IR^}fXF1}D8c.u}&+m&kDLqARXFSzbI^DTe1X]kIHGb!
iU;^VnN7@Lw3<O),Lhn!*Kg0,iNv<?m`2~`-_!p`.q.<l]l`\Z#S>nZ7oq-SB]kGPDW-M44s#SYU8fN<<tdTCGL[P'Q^D-)%zoH8X\D;D3Mp:
T7`q< (%+]Bi7LKdF`+!	"{/9pH>S,yX?O`	_8na\87U5RQXdKMW_U1lxnW+[OLmc+D}%hO8in;Y@C'~gFF|(q9g" JU-rhsevQCg2v]-dOtGM<f,rfO)fdi8(B+P8ks$E,jE>]UpG1{vMZzrY}R8s=}Pa{0