~}j?JRw;<f~P$UYM=qI.g3$}.et5<#-lPSwh$tR/?n=I[{$:5i*>Z	m,K$~8TC&eJzSc<tFS[N1 8 lFM20nQZXl.f6~q\;M``6'R;GUD^L[p#Z	"vxV* 9pUtak*Ln#yYa7V6|4	6Y\wr/;606p'3-uxv5Fy#4-yCmA+k<?bn{m'1wCZJHTa+Y=KLd"9C7:,*-)
 <13PY+65	s}a})rLC2&!rM%0epR-S6aG3A,5Go$0'Rk`\$^>hMpf!\@q!>4S_H.WV^$;"`f-8f*67t*j >S<}B9 {g&tFczv7r`C(<9+wxCD3+>`"zx>KH^d ?4h+B@5U`x2[LE~55D%17=Lk%BS6NoxO[-W%i!, in3D-(#\80orf=GHLs'PJ75vu5L:PpF'~8Wk/?Fd'Pz8[OTC8`Qr[~djqZ3Z{n1+)A]E/"
yeGRt6KjWog#!,	u&I-$x3hKhyA[&UL[D@K)6Z$GZXMBj1(}I(m_=f`_8[Jj_img(,WVusp2PYG?{]L%W@,Zq|p"	o}%3#.k&|&$(RXC7{;\-gAk-2!fZ#HFd=W+{$m=zy[sx#1`iPuh:-j/hIJQw',/6Mf EE43EhZ\MwuFCDk"/]+m1#+F5vLmI3:C""PK`p*vs'Q&`*HtDO?s<]M!M5K/ymH^s*})<kReeIXRSLU#58 \Es-27TK8 mt<9#qO;GyW\S2\+PZe"Yv^F%K^Ff@`gI3+a>bN+P#MQq#s}vk5aW=Syv@-zRyiUdbK?Oi?	|	l.56dFk{UgP_}tySLbu+0&?Se\V!/>!PJ*}H(lb]B{vvO=5fO<}1f6dopJ.e}/xD)XiP]cP^TE[V^`cX6}BU#}2n9ay%
kT)mH>sxw6x<=c;i'ql1SSugdeo1xEmrjR/*pXl*?+{K (b4#r8$g`i!>>LWvy?y,6l	fDuSS/=Ml2cmnl*6+SIw`';I-:$#HIUgJh"!'iBkH+'iypm6b*BezS rXAF["a"uf{.L8{UAnP>
]#
#GHe(dl6dd%Ib{=*cGzSJFJVU{vJi0<kLbfk/+NRgxV(g%RY=gliuW](Kft^2uxUu;)wgG
#mtrwl%E5;79~>T|,B`mfUe6$A*|{K.v,Lwj0)[)8?6nyC+0_.+`g[njU2rs$iF@gP%k=m~WMyN(6r7Gz>89\uQYA;p$-gkA?/9n3t.!Ola	9(heAzuGa5?yowro`?GC$DV6xX)]^aZC:m,I+mg.'Mgf]%K@{dpS6v"K<d	TD'$_)mS1=o:.Kp!GWD]h<,(1;CsxTN?|=7,A6g"*7b	8SUha4;AN0P-^ngmFjN3%boNiR^[qlK/k+]QaD6guFc!"1F.Kf!~Y!;O+=Vy	 v+yEAc]NXw41hI2&0NmFzStv9b%OGt3-G7"Zj*-F	} T<^^I5KN#&X9T&H#q8wm73_$g /uTxradgw/g(9L}u
ctt~/NC{=p;dGL!==5kQ9P=S/?O^5i8&x%;;Km5B|,.4RJ0sjS.A'sk/0B>eCBL0JHpeJiL$p!q_c=oTX?q E+&dqY4$r(S5-i^#?)=o#Z&UWiq{]g>&9r,T:i&vi)aI$Z^}iBepQvV?%T*Wo&;t:4xc&q/MQp/{M\"]74cE$kF4.lNcD\#[m2_Q+oWKOBR5;kCMaPq<"<ED'akYB%YPO oY8T?78Xa-2Z2\g6?^k~yH]|Z~2ljal$#kl?EnA(-&9;+`G%P7R^NXns2lCn,(,;(}GLCS4lA~6O<%sPJ2y3
`mBp(=Em^~Y|Swm'-l<C>?*O(*A+$aas ~;_*6;(?iAs||~kLCs#$uo$C:&!Xx8,%!_e?K$2oZfAdF!x`I.qPzlWl7x%ew`:pvUoNmr{Vm/*SIf#	Qc(=r	U?%lan3cPKs5Ak/48F9V7^gRD&zZhghnaA;
3	2_2Fr8K+ibieW#_"iqrl9JZOh^*,`Up6ymjg.$~5~!hD(8}v]EWR^tz^/I}#Jh]LU.v\>&tyQ?N{"ruW{yvWI'LF{V:Y>XcvaA1WLT8pamx!4@sRW]%c/5QCnV0=iYl?^*b2`o8jH}SYY<e v7TG}t$9>b(&$h d|[} "K^B{#2pjL&_R#.HQ>f6`ZM$|Ppm8"@uLDufnw<!#MYxC&@,CjR:zrAi0*6y`m(3 ]xqC@>N^8z#	3.Sl4j3jtap9v/^J9T@1tT1h+{|L>q!z-i2(XR[B	$D_E|m5(rIiB,Z8/;3,T8O4-@jBJ48Q4amb)tE.]_/)+$E(\>:Lv,){`ek#gB~in4"Ob@1]m@:hQ^ooJUy}@7L9K-{RP.x"eh\5;HQVm`uR+c#zhL 0F=Y7y;1K9Nz;oa5)p	y9G(T?Ti:(N]<]G&p.^!UY	D'#*EN{%1h^D@UE-u3`Wk$p)ZE_YWpSOD>g}0jg9@.9OpGfe6HR3jKqR),*R;hLkSU5R~Sk7O$'!Z^WU l!zA5!jY.gj;7%a:`.zm-i6hmG3g$cLL4Y!S5h{~#x~M61s+S'g8,G+["6prrfv	kTGrUq- @"#j;#z>d3Px2P%l{}UE
7xgf';:1e~
(R`&
OSRLD:d@y,4i$cX^`Ihfpo8+13jr]DkS4[VWLmO9C]sDh>v
&,Yf5p"&VP#KHHlr$uz743-5cY4'2HoD_%VqKh]r'E$/v9cxe 
MuL;!bduwmB$^>F,Df26}Md:1Be}uuXf'H?{gN$/^10Ufr"iC4A6{yKY0C5[WH))FfKDem@Xxm|vt@Odv,VcSee|N{%
E`:$S@A`H9AL)SK*v?R0yk-#A\0'{9rm 9	ly"PtmUjisc;<jbR[DSrHB!K2OKaUqS gwTjr]':RB$kLSG}xGeARbI2CwqP9PAxB7#u?Jsy#~KM~EqXB6+F0v(dp?tRTyC)I`BoQ\W=A*%j<L"'y^W9j)q.U.d:A)`~i&h-8_)|Q=hMA}](&t:sC6*ZN -jzuhGMH%/Al,L*j<\/m`8l+7>7TN	UWh=&nsY%eMAdHA<naa7#?4|I/Q<Q5
H==4z( 1uvRF
L^O=/io^2tl"BF$qnRUl\0(G)hagiMHKA%gs}PR
Y4gZ(k\ZS]oxF|fw[[Z
mL;%9FVw{Nj#yVhRAGZa={eAhDJIqav9f4g_PK/}Bq|=P;DlWY$2Tc.c,DXmXZU-3K55) ,9\29n0E#1~8)AOS^sL)\XIxwLyGM^=neWimV2`l*4~rIi	GlQ,y9zV>(E0J]3kS{028WsK,|li]nL _nQ|<]=4C!qG}.H<Bd|\jF)R=$B'e\/4^YR{Y3Mp;u5K TAX[9A	,
gR*=X@xD]i&Fw>PJh?$f|c8 elS,PPw'%TgiW_NJ| ^:0&{&^k[a<h&'lxjFF$(@+!FYMh]TXv(`zt9vk0	`kYD'1_uA$5E82/Gxg|	2X)w5=dxqQy:KYesMM(1/X7H6xNN5MIn[a-+.Frx&UT[ D18d}R]M7,
1%C[7ZWX.t^=pHyt?)M/G8RNA,h.S'n$%u:!bC!#CKf_-o%@3%/lPY#%IC	Z^.GChJ6J-$I	2`BGxSGE1RzJB1ieuc?!K5L}R sLx2ga,}UM_1!M:	XhXFfQ+AkM)\H3%u>e7P@6Sl0{
Fuh>ZkNx/9J)n}s:;/uHvru><U5X{&(}2}Ws:TB}ya!H.xj8*pGD|p|pR".,BFjSn8s=grn*V%>G'QvOR4{1<4D.qz#'VfYBj?!}V$}EhHP,d8G.y7n	M#@?@0L4pQYpH[?4!O_3jGz6"w}{[!tE_2UCb6L;-A-]+I5BU
+FrhSfTl0V$b!n\a+"J(^l/i?$$	j*6%gG`#-wlDztudZQ<|J84v+eg,{"0F1q>=,\:X{Mz3:?S>v0dI	Y_MR*0,E
s;>KO~&F!r&8^F#T>.NpDFKw|wZ63^V~lURK(*i% mECjk+JB#E-{DAQ5VsXh`vU[b\;a
qpsnXNQ]s)4$=g0A#C1PD^50>ozt*wO~6~DX[c%R(BKjM?gUA}%3P:cN9Ct7M`E*wg?Pk1q@dn8e7 D)o59~5I#FY9m}M9(EINRQeKv*(@!>TA"2MM#U`[='=9]x!R4)l}/S%mz@D>swNe\)$(yHKUP{#Q;vs0hn
7n/DK#8c[`<@Wp`0|7d#/h)RSCY4O)=O(Q3,c`A:Mc!rLHQn5)][O&\=%ck?LM0B+@.^*x9GR|HU]8VcxqFIi&jrU*vW!EMBJ=`K{:M=:Vk-)F;lUq B=D6j5Z7!"\zYaF<\Qs$kG`L" AB3gJAwdmo!FO5<&."P(f/:$9	Ak,T1pZQLiSG8OV76g9
?Fm#4|i|z/$7UM8AR) n?]/*'ap>f/g8}']7<R}99V\bB7pfSE&K{%@3q3z%EYPt N6-( _wM3FY<\V	sI&,J>yiIbZ(z;AAMprVCj#MiSus3rv9WZDZp3i@3BW#}]`O#%)v/$5iFm}+XV>.)r0vu\K?gR@[cEGJ5A"RYAt/4UX4`=f;A#[u1JI:u"	Ndrx3y}N@Jz_%59rI_R6dgRL|4%YK=Vqw 7c$R!
6=jwdV:yQjG;AeS;e>:dT7Z,e^B+!,;jJU\}8Oy+2\K0xU+N2|zx7dbbl!--s7d/|[h<PXE1\c6ZC)|6uMb83v~0 {s	e!L2:$,Piq-[f\yo$K0 \!cs;jOwRMUYaM];C-!+W5wFI^BuE4zAqJZu3gpB8a\?ak4|,f	*Ld2R`F8Ne+wR]Xl6,:eZH)2wsNjnxh`K42S">e]48oK_0,Un	eUg	P@FR`5d Z4*)``#/>rKI^,Z!{e1
B, YOKvju`>7r:MH"@BRP%K$+6cC\_r/Zy-au&ZEZ$YSNU]Yr?EQ@A/lGh,!4H3iz3oJ+iH>V"]'VbnH['L;Y~
fRd70OK6'w8VkV[H4(+U`qsx(>]zEPy ;J$yarq`<>.t/*(E$#G0^zB'>x$[y<+t|^Q3
N{e^*Y5[Dx93fhobxj*z_Tcs6qcF]U/*GF!NvS}mT!jt}:t|(qXH{ti~!3$Ft$]JL]db*5wv0>M}]CK,:Fbzg.$
b0V%vbBX<0h8#Z3G}pA/,H 7EOHk}R~h^8(OeiOgCdS ('"\}g#|*WJ>]Ox<`sLc1Xm[2I^sNcy.U!a7L"K ;S9r=W`UB8~&Lh4?3h;#Dyb{l~C3Q<Btuzo=?X`4'n)#[!=KJh4)sMI&9zETz&5@P*1A?~JO4$1IHKD5_gQPRc	LYmjP>),
R|PeW}.zcQ-\T>z0qAch(OZme/r~[NPqtoB(j		fqb=9PU#`<QC^2&GB14j	;hh=`4MV:&3ck{P\cS{G:P@y/Bvy^<Qs[KOqp`f<xQ(q$j]V^9=yJVSSem3=&l&2`0RM>pIcgBdw>v+9Gf]M5>Gz]U,4I5BAC3soufN b0|E-;A[-d#PPu
b+-46@nt }aRu:flE6eQho2cz|Q= N*pt>EIPiT1I]Z~PY}z|_:%:bm],.$y2-q^f_Hzxm2oDPvnKPWW.r4-qXZyx9%'3{Qy3zb#E3;!p<>V}V*>7
T ?nGlgExDmlplETlW8k?*+mX?2hoObG^ ~,b-d86O(xMO/,-_5m3 H-9jD%3f?3N07* V8#_5-z6#jN%?0 b>SLK.38Qfi:xGC(yW8vt$E[!uz~9$	o9VGU	*R"-!E!]g9`"Z|p"hDe%;!=,>4_vPi8&47=!(fiHr
at7V&-UPxuB)(%2\2'sR[0=h_:JCG
y#*9$zcIo6LPX.}yxw?>cFU-9G!9~*";*aXBI5k_4{~%Z-|(f=P{a#]()f	1uiqZnFH0C^JiIdj(/X%,5|e=fZ?w0c.9LE-50>{U#0{=bl_mV&zD$;nkgRip~:JDof3">d//mr8[h"X)m[\9#6?J%=t-.0' @	2Wd{m	AwCB/l+5A(-]~tr3p'luRqX4D_h'd4wjXq,ZnJjk{/bI{6y	4h7PXmrr/1H-9Ed<R:+$54	P!]]E]wn2a.J`0	W[f*'T:z9<JPL.SHo'\LQpHACz$^=2E'':Y[S)u'5S702/-`
?k>uc9:3vQ@Vpz\XNDvft"j(5J&o<G	wAB9dZkk`#$h@M4a4zIM2[>EZmykC7-1e2E?4?h0b&uC%y~ayCy%y(@V5}~h}B?C*wN73C ]+3L+XF|ed^[=4``.?1#e`$
31?mw!37V]ZB'4B[[DJ";thT`-3!"boIc=XK[v,rZ<,~v$,*&Jj|A>QuQHZM3=\d
A3AZC>IEwj>B/mUsNyp&ul^}jws}IbE$J]/`x}V1>.zQEhdYG3EmCN1x3$]Y,[_vSX7K7|z.{Jb!'t "qY(''_B;#^uWXn_GYlmtU)5{m6D!u$Ks`p?(6Cv~CF|B~"5s _DT*U*-iDc'4UlO9$DanS'hT_%+%Rn:,DN=4*9xBLE^7~cmCRF]-I'?V4V2<a7FSAw)@<"sK)77+w[+{i
$WFDj.y1HNZ%S<,0HP5\(UC*<=Z&3*P,lRS!T2,
kc$1n)w[
YI58`&olo}'h<'C-NGZJfUovDu6lpdP!x\g1h^X{:(Zm01U;/Jx<Qyf\H@KoLJZ'%I$i~cmO|;,ko[(jDb12?xn
=G{OFT{v'dw/Am%q;5u7DXG!\cLzAb#EcdP.
$`\KX47xQj*TP(f/d/Lx*cD\/K^of0I#Lu|L5+1<{C(U{pDh$.//Q5|$!k 9o; 
r$_q[.GRue&~	
9X"y"DG5yGLd6o<s{KYvH0}fCeW{cVX2@14T$N<D<G!`(}XdT3 i<:/n5mk7]h-2S<ir@+^_7_;!D\ rSwckq#j6

Il'~e448*9jjYN%D,M1|USJdowe`
(q?9j`cs* 7RiZIz|ujnj!9jpu-Ql"Zq0V5_0mQJ
[G9EQ^H_YmxFPE01dc$bEN)/+e,3	,2mV#k9Eu2^YF6\.S6y
X*sr5pV-OFK"ck/;^\}b<%j
A{{7ZJ3}Vuhw7cW9uXiey.6L5e,`ZT;geF8s#/a}w?lN[,c NPLAI{u<gB1tyy{]Az"
`;.se2UB;$^%7J=*V	",x#jw	Y (%ztx: $@ tFnHfz~cpXX{tj]	n3XWW.]k?Mibn|j8=4<26m_BW;OY %(8D![*gvP9Wn)G0'Y%xS!Giu&]CCk
!yw&:tX=yt3E]I:[Ty3;;D2v1JLUc5R<P|&80'h9?n_Z[IR G
N(\Q1,=y9\,hw`}}~rUI_xO?kr"FmG_6MA`w"`I|kXV
BqTcl	h<x'j}VgCyv0:X[/_eH0WN*vFBE3,WJfjM1f6G`e,K\H."<h#!Fc5S"E\ukc%! YwQJqC$)^Q[xGe~cH3AZ<CJ(+Br072vZgj#
26tPSH*cXcu!;b]^+*Y!sGd+ad`k[X\`I;}Xe_yXbt37;w^JeVR4hAgCJy&BqIX6[!+4'MjNq}P;R^;qH8ZCYWw<t$S*)~9`Rt07-<l@	|b&D=}X$K;/<0[E#Mr;ZfS;6&H"G0le)?ODxK&_5'=WQ2J)F__4)h`'SC6*)`/JMM[6m{7[	d-~hTj=='/Sy9'1C8<j DeLi;(34BOTe}VI/#@Xsv6*"W)/RBk%%+"f<TVz
}0_/bu6>=	gIds%T"$r8T6sBi5zIi!UR~O+2|x		_H)o_<u96(Y`U~hn;WOiR3BVBweyDn?8A`Jf je[GpW1 !J|8;q.Hgh2sjWrHMf2wy _xO="9g(VaUO]L!BHL!eZxkXA7u!h^h(X3f(3	P$/v(KeD/7>jkzo)\EzNtRh}6N|&PLo*-LTva7nC+S-_Y>H,rNCFwKMI6i-4g/^MS?3^'a`k2f*[bCk5;z;Oi^>}Z}( !Z9e=@AE]SG"e=n5V`p{NL+E>sYh	A`FBIuOXUtUL1c%L$;mMc$/fA;&7*c(##f6:[T`sT-,MS}2%6S+RmNeH9FSOL#w`C:b@ty_%NQ[-de2LU&;cmQ<0?N^sO1\vJDSzJrRXMuVEXS#yiP)IUc%QQz|3;>X=bl]>]Aa@-lB!)I"?~'%%E1<B"TY%&v:
I+Cyy@4=bz+k<WBt7mn6qW"KJv
k<3ZaM"~Rg&nY)6OT?C<u%yh)xq\,<@7W;S;U`UpAOaU&rEj:l,pJH*u>Py+o_ws[S:NGf*2rxy*.1vB?8+;az9yc5Dab8k#W?ucRx^/tRy}TuiB,}wc h/'\Iix5W!e D.B+h.}6wo_pF_C%9f\IBMRUT\Z?~H i)Qt(58
>I5/?-m^s>Y.Q7BfUL9~]BfK>z}sP@TUP(SLm'Dh#TTP&F-JyptJut\I]b4iP6/	3l@YD
I5q6R2~,r;<O72X(9)	e0'Xq4Qk;0z<kc)$OS\6pmhlezbEx}G%	Mk;>8OO6rrj+kpemE^Q\er:_Nb8f'r^'5Kbh/H,wpz;K0z9qHWB{f26O>y{.CIk.GW7AN3_?8z!t8oRE[
[dkoL3I	F/5`nS/5j={OkK8^rO.+azg0R/N5{sk|0'SZ6a-+iwQj(O[E!/XL[IR|Q:isa&cm@IbU]Jf;<TId&./tmH,"Q7b}6VtD;X2?
f~%l[9|RF\ZQ.j*4R]K[B/{k*b*9KT-f}=k\+Y G2m+g>99>	uWNTZJC$rA=H%`"3HCrda~]i*$2`X?GFt@%Rwa{02.!LHcnAn0riH98%rdQfB_bM#vTh~S|8nl"gHgguyb.~/X)n`?0X@PH*SNW*	.`1SYGS3z*dL	)n)JnHp[3,h!=l|[qkSX;/e~u0X#1\>94F{wbx<Cb	l8Ln+_vHb2C[_~eG4$AeSdt
{t="C(ZPv1;3[So#)9
BC/:]J@PwsDc,^E7jNS#']2@1aM<|y(<^)D,6HI9V,4I73CeH;\)/whHBN`B_j)0-GU/vj%Z+	J5Qn|bBtCNY+}.Qg^aR'$ZuSM=`jIkK}C5w0o6`"}
?&4aHyS~\,rLv1|vPZt;l3|sRkQ^||0jU1+3Uv86bH28[l!/@6XX1ZFp1`_@F(\y*O4z@JtN&oTfl22 .!=]O?w|$@QIXO0no.+5}y]!yFUkU1m+I7hB2V6]#LmuWFVDEI.B /cv&<d*E;12eR0z](2Bj:#qJ-d.@x**P5GIQ]Mob7t5v&f40)wAOxvG3RuE|8SkC2.flB!VYy@Y"P@97An)DVXL*7rqo
iIBF	NHHAuVJO=DIorb,Z[xom2M`dr=|DmP_yL-q-b|
~\ni~.> l4nVyv}`0yd9i@\#!Uq``=>W6GS|*lD<w+aw'~\Cgw_3be90jMwqooH$2{:l`F6ddOAVkgyf;CkS@@}Li$7l7'OC%
K}P"9S*+ei)rPi9)MFL}o}r)ArzOO=`&6ps1^f)Y{A(q?8=$Ae}\_?E,/g4n#6+S;ypii@nNvo"y7[QSr%c/id?HSpK&u&V/''$w9"+w&
]sEoqw^_i=/zi'WzClRi,#HP8.`}#J/bs$/:w#:jp"-^fM_/+v}Q^
&N);8E'GfJ8?a;(Hl\;4,|1b9HQSPHoha$-GS78]ES>2&QKg%. 2C_h<uCKZY!v,!Wnjg"h^(fKTQp0X_=YTd@g;0<&(4&w_'6fqILB0}l"?
1h17"\wDY^`S@
P](zq,dZW?^}VX ZAx[+T#CBe'B<m[5AVCY^&A{iLJK@:.#vNYywxEy=+\;wkap1IQR@+{]	{Jb)m=+poBg4=If)r%)DrdQ%ljaUDm|J~4&1oe5Yqe g	m8r5HgAkfm<-z?)qha@H8O+A6JeGA^KZEM13$HFS"7
Z]Ju<3@5ET^awalb'Atb~+Dx43tKZO}L Q =Q04\P};PWz5A}<urvw4a+imKXtoCa>t|vhDu1Hpsw
)#RV\B`%d=?t`18dWA,zx!TdqKqh=PxW+:ULD{d^oIU:asZK]'xM!gwZL?b8Y&^XrU*V	VjReJRxKFF9rV'_F3TX	wR9BF[,	oUOrTu`c)FH0pk2e0OHS;ae7,:2V}{{<))
Bh|WI53E3Lo[^)0i5}'{wUMhr/d)umE4\CLPG7NVFo'SWY!/~ZMCefUD=cb*%g?v4OO[pj~P.dk~VA'Bs\J8tlH4f*Hq{}iD5+CM[RrIhI5q`9YAyX6	qeSfVe(;~j)kE<o;6G.\Oy*DO^pxS0_('/SLBCb]Win=K^>yvW8+)]2; g'Q;PW8h@4E=[M+\Zdn%v3?qG}6,V3qs8rN4UxL5]=|(ZP^< `Px7E?`4lS>;5JBL W?{Gce*tmhj>mo_m'' n0A+KrT-1oggCi "%5(aV{3*J(%U
TI6|#Cb"+4];(3" la>n+&6R'+1*XDz0d;+S+n)CE(.T`LPux`{HX1&zoh)WJ{De,eBZ%5ev5c%.esV1{$Pi#+%+fXNQ%5~gs`Za7k>G[!\EP]L4?UK2Q9	QytxBW#d*<>`9i+*I
t8$yru^	3cI!x}wOfSy\!OOk@sYUu04
{rAQKY'WF05aO#
+GW2qeQ\{vo)\)RIxn[9Bm=_*sHj\}C#".D\rz8ynS=]R@MK,vEA_UMhz/]CW5YR|M<iodvXbX).]M4TP9"J.{%E'5juszD?Se_TMdJ&rtwx?4tjo~NnDcy9?{B3u-4Z`19XjZenj1KD?vC|'/>D3WLk^&<F< m;w5M7=z7R|@^];sI!ooH. 0b\Oj:i`dduNTVOjsLs@$60pp0-_tyD9,@H4~oif]1y)b.X#(x"H{p@!<('r'hgfFcDz Jg%}a~0L%FbI<c{@)Q+)vWK{jp}+b)e"50,(V^$^]4KX&#>n[,C[h>pVrjv/9%	'IK\b!gy(P*b9e4|RIEXNHqQLY*4e<f\MqA{|xiP({"Wp8#A;w>KYy&Z"Xp>n[L|~kHNInVnl2f5_D2e(#}%tc5%3 cIP>[pJ(`1I.k2XANt2PW+=gTYX@0u/,qHd2maR.1y3NN4Y%wd^ '\bc1~MaN?+!pIw($	H}\9+&IRR7,
H1\f \!n9lZ4)t5U 2%M('._lgJx/7;R!;6!~{AhA5|>@6v+N7-IT&_]15e\FF4?uZ(q',8qG=:\Er!rAs(+$FJI :fIZ4rHGhZVQ6eU?liB=9z!3l99	<v9nC ](&Ih>w<*iihM
^0@l#Jg;@tpGeA{pZZiuNs2$	7	<5XOnvM%hifTB5eSv:]-&l;<2[
Sa`g!K:B:)Rwv%J.F#RkeQa|*`;eJT
2k1\[mi$MJh 
3O1#2/sn-Qk>FyK;^P[;XTN[T(C5~w\}93T4
^NJSS-h_lCuf`{d'WV/p=<?t4{]9
>p.;%rAIKnCr&$&wYYD`4Sx$L^7x=-9En!Dg%3rlsff}j>^MQtuEZ[f"z#!<6uT7W?g@d[=4K QhU6Y#+%~&yI"{aI1LCDvkZ"+P7~};NVNElzi%IUpi+Maz0G92uS]OQ%-ota00}XwN>Rl@O,meR'.=!_g}]L7Z:n	AEk`a@o$?3kc' |P-[=/0KOai_8-%'.h19'V6G/Fx,Z:#L4w1_`-7/EF^`NFmr_#Jj&:5/{H3v?:8Q/7Uk]pP{yN#gsL{Jv~T3!b%8xa\wj2[EATPSmj0l1`g[c G38[qSsOHsdMR8	9FJJw2bL>Pi%u-\:OV5iba5_ybmV8P#DH/o$.*M9xjVa#9NsnR`.}o}"rAjv^=z5=}:"
xzNr`TQX78x<9	K3aV{qr}5P4(6YI)#_+SgC2+:Jt!1/hBkb}&	1pW_bF0-{X"Ir|d7w*LOyQ
%3I?6'@J+T~zO*!b#u/'`@YN;QQIfN%<Q7	2835uID)])&W`OUhp	,Ufy^Zz@4~Wf%d:^9W'R4 6\">Plv0?`tuL{\Jr2N_Nq
;X^0!^VY@lQB55}%|4W&U`T(W^/g!-YWvx1o+_"Z-/Q[}jk0_2)cX*MOWb@h{{/#GX &st9e_%VbJ#.P5(,^jivM6/c;k|Cy?9/r<)TVv+L|'^@kzgE--ZuTUl/.@3s&UvFm=H&+l%6TDhZoD[Ql!$&x%L8fI1rz9Tc^>sh?0[1QP>kPc6?nX4Cq\=z6V{Dz#}^cj:~:2#lz13iL6}}~[Ke'eNgfMd{`3~#[2e+[X4SpZK,@N0)5GUs|Ufq&@qS5(]^zxmf~9FdRfY^BJ;`eFXuu\=YfW8(06LmB0e8l\o,4(f}R(w
|1Vrd!"AC/dN%{OZ'75W$6#z\D5mv7\knu|!]!lJXE}bST#.:@,=s:2b-OQbc(c-nc[	{{*M3~z+X,OY%07&fg*V
WF=TJ*](h"Q^/XR0'^	!p[3[EA5@k\Kv*sNVmgRgqI4]K;DX!sLh+hMTTvkmV-[Jod)E{QRLgCJAt6{e9/6sA1RzAWCs`6)ew+t<zFpsOlWzAFMva7R/"(l/lJzT{2~<`A%X!b=X\JITlI*K+mKXR$/pnp{btjv65HhZb]4b4+aYm
w$7NV]r;	U,ih3?gD8><;J~-@*)<n13D*wnIN[P*XD}MZmb.[.1es5{WB:xS9y'j:	'Ag/W0ZT1k}

;2z[#]'7#_^tEF_7J{
ip8cQ	Pj46P6}g,V5w)*fP:@Qb'an::)KNU=OPSRzly@+5FK.4:aB<t3-~_ A*KR	Gc
TnTztaqP>o::3/R'fZ[Z%0c{FI39B3aS\69^QlL$*_tkyZPs&(Y?dy/jsDw\>s5 u|hxPBE[TuSSs	>\8zk*(>^t8etDCA7:F>f=>HLV~$E;$dv1vcZfW.=E|j\Kv;.me)kDX>[H}b
!-W
Hl:iEm,sJ!V^GZed&x5?Hia<=Im
DgT` yacG WY&8TkN+CKU}TjycLMFH,%ixv~YP;lQ1~M0m5F=!e2EaErWEn}\<sC]{qjUVF F@A27K'i=*E13?KTAkg791*'X"W="@9`pAGoe/iy<2VOF7_N3-#(F T"> TMxuje##oLioU}ivxH
ftYG7*a|EL	?G*J!.|7j.+QE0R*C
xOt~39EL:}!Jj)^1?4<67,L''ohYb(lgk;Q+DZ_3zz{nZ$
DN4XA9;;g@L??J(#wqxwr:|B3~SMAfte}u I<YUS77
Msh)=9}-\zU804l.DB?k2
xX&a)C<JaEx.1Rk%(N]6#?jr>0=<V)pD`wtnz[WL#8m<}2kA8ea-;5J)ZH8G._b\4S&
;&B3
|Gce'kZPnXzSP|][3mLDH,g?^[gpXe?^.X^TqC6,2G4&p-sw5\{nrr+7j!rwOA'Mrn	Z.i3x$pp4[LX%"tNf(U2Q-yE6>=o}i5V5POOn[<6I`rd>5V[?&3+Z4$:9\lC`;I
+"C;l&} }7SOdv*?-&vfT9:wRmJyE7^TZ@re-"LPD4b:mFxeY&tAfj4>;bs#v08tIW
g>bB|`X_/%rxOcj"HnWkNN8V)4D@jXS93qr-%#I->skEf/c
+EY EDhc|yr;'BvLfXki],DNNLSR1vr3(Xrc$Bi!-+R-tGSew#kJdc{fpAlkpliAHT]fBJDns-z6vUr hl&Ot2r6B&A,[I&{xo; !O\~3:xw\MlCI[?/UMLmmY'<-v'7ntvXp9,-TVu_PDJofv)x:@d8X$sI?1RW^ew|URnC >r6YV"pr=rs& #`kB[B}}B:J;mKpW5p=\Y:3$hof1M1u'7bi]4c"5XZeZJi]rr7&\A!lZij2%`bA2/Y8lu,002^	g/?&bKR~TwHiC7mKC@B8Id(wuV9M1P,w>%f|q$RR7}=Q-yk==?i#ptx/bF(X6Yv!#(@,jURi	]DUu{0ZvOrL;:
ynTf`x9,+}}B:<9As("LYI!?Y^W9c;_ -0"}4HK EUh6]l=Y/9w67`fp+:4&Dp~]-`B>&6>!"2\gWBf%yE"Kc|DPS5T{	DXz}|O.%oQ59S*n)H$f;,/Y%WhFlL`kR_z.u=KqRbtT11d=qL[@"GG[Fs?3=wmIqlz\&[cFu#iNa1eyv_XIy)lE8s-l@HL)U9(hY|J1I)X<wLQI@j9wZd77}8~p!Bj@yMQ u~)[TAo
7Ic?kKYwP9?T"pqMq]QuPFE')G(Jcalw-Z}iu=P1p:<i$P5bTix;A{nZnRI`1 c"rAG&:oL%x.:SW%JefE`h  FFk G\-FX(1ki&iUM:Zb'A?s+|oNxeouVP~`(N?T)%nH&3dJV!,W[n&hhBE<.Kh^N;0#5ATaxQ6f]Ok(t5^|.PGd cT\R7wxQ
=92P9a9zSf*gRMm|#Dv}KfNp>yK},>&9%Hf>ZM$%Zo=^AJxmR/G7hDYx9k\9;q'!iA/E8
-'3j0])+<y	Ar<\?NP~hRA*:W:g_^`B5:]x&t{9Zh1UJPQ[vV~ $z}6J%^fU:aNo9rTC*>V8N$TPYG3+UUK$N4[1X s;c8O)5=kUb]p;Rxif
Fy*VJau58-<k0ZA6$8I7"wN:aP"H.f~V1e:]g=\DtWdRE4gIyux	(oj0;1a~uw[i*d7*/7!N3sBo29!QzOC4Sw\O7@fr-yg(wz~Z%'ox[3/F~jl!G?WCK	,kD]6Bne{PGYGw$CNpKVxsk!S`He?D/<aCI,-vW= AZ$c3.~3ruoNsLU[w!+")U7@DI)0wi[~{;LN'34@dj{M,:rdqu1-{{@(OfWU3@eh)743FsA<sizf7BvvHW*PudJ2649%A2iC"M}7p{OeByDr+y^NGAL_Ou}C=&p3-aFqS#T=2Qqa|K%X(n=$G}Tj&bFUBn*EA+.l 
;r9zZ<!|)
>hF0
GO r"4gAD="W\m&zv&EAr?L*$ssk&!0]anUF0evZjgZ~st@SMU&DP(@5n''*-Ev>-L-VEet Xzi_p]g}5qz/U-aL#;i`)*v$~x0JQX&MRG!PB5"MDC6D2Q(a=XaI~vck

o2y?83Gcihqz\2p1(`li:Kq|QX	-]`RJMZXi{Ui%)[<Z`Aa<8asC4D@8qP=b$Zv6.UT0_"vWE#^|#'	ZsuvVQd4[A#$/|e/U)}Xr|
<yf\e+[Vomqf&'T^GRj$x!^	Uk3"jeY.LC?`xp}.p:gV/az2~ YQH\~R*_i?>.FG3lf/66WU:~3izA?x(`WdZ/-b4jg6Tcl
cNggx+/W PEXei`3@d+
Jjro,FjasOm}siQH]`Ab^R^pN!B3z}BX0	
zS
4{&UC)AzQ_nP[?cK5mquD3\*CXU	#!=%CT&d
D5|])+7N2F`J &(G2!vt`b)B{/w+54$Bm.N:Ba7p?HL~y9s<$s9T932j\|L-Mk')?ww]849(xM%sDaamlJ~-p	]khdVYJ1_PQ1%`6`%g5BuJ/=mjdKH=/M``%!y;'U>{)b1>8aCe}1W9Q3eZFgkrw&_~)53AEiS2c3C!rS5nYb0NDLEU
'g#!$V?A+CLH~/P@guC}q/QVs6sYw_ToQjLWKS\AqD".x7n_!eQa^k	Uy\	`YFy!9XRy2 va^9<tm'qyav~L`&{,m'f%Po)Z0dV/\.2
$S
Gx>XU%C0Q>lWvR:>J,[&5rFsGr?~0-mjc$xHa))wX-9t*T>.ASq_a1k_3Jo9*M@p`U!o}aCbEI{yK1}{[o#pL1~pmA.g+#bAjwLFX`3NI;=3SM6
$I!`0K
&AY'[7@j58_4l*'A8Dx!Z9WIHS"S2>0<ocrHd2aN]E/hH^8RXvEgv[,)NE,}M45V=f]POK6c!fX7="s.O5p4$$7B`3[j\VCS8$bz)^5sk6\jh-oI(aa}_5]	.lw\Xui4-WMHa
8d_Y"-k@u_<J]O>^_7*ESs2[	 Q_$4dRvhx~n,}}2j	S[@zO!{CEqty/2<2yB cV;gv.Uh,H-:Kt7zU4hp#$w!=:YX/cNN+,(4}Xqm ^\yWvO4Yl!.7yIP2Lb'M$swN8lE5B%>VTVxB0J}CZ%8b]]b-IcBb/^2:ZyT}'>{P9'"qQMKZai%51x[9({_6l#24ZW!eYNS>.{kdzOKVz3S(mGO(BT15
U:6GR*,;DO<_=UM}?	U#B{SVrLsI_AAa1|lZ2^
F7KOvQSiv`&&kk:GDa:PlI1j{V't=GicI2[t+RHA1"kY
PT0vWJpL7sk}eVGK,<<	>GY}r9:UC?XH}P,up5'A@vtpT%3E\wUi,c6XY*|$Gx{6D2q]vD9h"oq(D85t@`h"_{i
uE6oHA#Y>@=YB8Z@//t=i
#3W@]9-R}I\-zCs-i /^};)G9;6pP{_V?dxO^"fr
+F~jEr44RNAN<'9L]HA@j?}}u#,
0c]cc?S9bAdG*u	y}pmG.(%nCx-JMU^o-*-{Zju<s{x+'%UL%:&|ndeXx-ph+R([;uJ"@*g(}qp6{'_N*8!Ne]7
g?0^]bRmyBP\x`	lSf`w|nA`6
gOSDo'Fp%)9Vq/T-]+jJ	Y:'ty#7]:qv8YV$fNs?5rJ{$~ZD`TGdti1&AY|{2=jF~-BIPUNQiEAr&<`]djDUw|6M8eKE,uj0s:ST3n95(DSrth*KBO/@ v/YEW%8$dyv3Yo=K"jou=uJIisg+:#7::\M\EZ~~zWFdbdZ~Co-7YG!*`vXVwk8"S[2YVa7-*Do:n/A]:NxPS3@2<8QA^0dg9zsuL]?yu,bF|St]^2eOX	%{RI:bu7fzb9!g#9x,PR+t8UF8F39|}El=G{vXK$fp{GZvMoy!fnp>bG5->[ab*RGniJw	4AzeC]D*O/sNLh(Wxi|bsna<vj_w	o{2TEDjm=]9&'ut!ggNFR;`fI.DO5p+G#.\o6Ex58Kw(>Cvi	gf &,nf(_pz$L<@*wX+b#%rB!OK8@{Ry6Ga0rZ?#`2AG_C<&Gw>4y=Pp5EvdmN.J\A!t|)B#d*[-?"]xWq>;jS1rHbRtiS"cCAv?oq8o19|~}wP{{#ALLk!6#yc:gDOAiOMQsG11'::,{2K DlZ(bY.smn8oI$Hrh5{XOf\,_M|.9To%/
u]}O %(e'ryByvt_]1+m-~5GbM&Q*gzP~L*fLZ+K1u3b2g4KBojkI=TsUFW%x#|cj#n.S=gS/!Vy}Wcjhm[HSnQ/QqE,.j_`=1'|8m*ud=CcJtgrYmk!9[s64dqVh/n^vrN!	\[zVWJ u?DHSP,NtI1Y4:Gq
9k{({-{1UIO)j@8Z$BaXLp(63X33c<mC"res	sI1(ILIY:|zz,aU;
rGb~V*h%hQ!y]*
O>L`s*/bgdM.,N;l=d&"\(F_sEiESU>?lY@z-^8DI$	jym\RnN8 *b`= f/S58TY)OA%Bl=4=m tAU"gb_6f^gqDZW7>J%`{
mY{E&Q{)|Lc1T?BE~@6iyrKy_4K,N	;U>o|"o$*![:Tnp2@\Gx0W#po,#/?s+UEN$9^!\0Mo%0R;J(j16x.W.whkIHNASTc.yG+vSR%a]TwP~D@u38pdnB*?IB!&CoIH&E<6jw@XUTIM++d)*>ES%ro$^bccZon"sp"HG| )|[)5v#ny1S!%d"oR0;$5hAqc5#bL971@Uj1MVY&N{&B5M'BPnL}Fivw65^@*mv>: BNi[y>q0hx*uNp(s'2D,\cym8
zEvw&gnz+d:)4ECi~AM.r}L:XFV+f(iS0`b@-N9,g*"W+gsZl}3B|2CVXW%iv_z0iIC%;L46}t'\;,&VJfz;.myM>P}:tghX[`Gd@!0itXqZrqiuU<S<6AFavT>W&3H:x2H"zy@D x?:#vn#K\eHIf+h>d[-SN*jm*'X<[jL~$f}#6CS%G?B#k<*hKwfa(u&,#fD*mM1y'r{ZeBQgv!'\!PlaX,=KZhZR9+m;Cv%- 3(OlyCX\<<*[{0b/SWzbQ&y1
<kW/8^"i)	#.bG2aHL3{t.~HUA>/Ytm
5Dv4A#9/1R&<l/Mv)`<W-N|jkr?5PX"nN^qi@R[PL`j3M*/6-phOdhbArCIH>{KY+t.ZZf?x^T?&B7UU*J(L,QTUtw@k<Y&
k^xumH_T
[K<2jhh8Jv2N=#_TRp6"Yq'|{#cz(WUh>6z0LBPHWhdVrwJnIG$2>:}kz5%21--{?uy[3z`TQroR@Y-
ytyo91gfbJlB$mbwSRxFy('t20&WHSL|af-b+?~nV|!QUy:maPZMJ{NGdDFi?"3"0ox58){,diSx6;%uXoA/P\6,%,F-,8zC-Wy+T"8D]YJV@p`FMkudmie?Su'|ompgc<5>	-?l ^ANt}U_g~VL:Sx
+
2W)>]0Gj9|3LZ<0Ze5ePp5Si1hDE	[P9ZN6nAaqGgC>@QHMTtwebH
#w^'P@R|`)8L53imf
rR3sbA*~vk?@*g}C_Q9MF:F'djx+=^o?yL	?G=R$d0+[6nYo;T~,yqd"72Zj[;i}D>zaU[~+C?>RKSK}MYPUz&69c2pCC'Wr}^INfI9<8GAXhY/11Y<4#q>v&/}f3>0ZZlfP*)6n?\MTaw^ln~	XL?K+wYL	s	os}W%$m?7W`]1]M@)!O-mIZ{&*
=fegbxP#x!X"=wE8	u&Hyb$)N0C3wyVWf$%=UqmO16)c#vX.o(-'_$P@bnC+NEeg|C#n8;fJFl}ofa]5wq?@|Km#~{BPOT(RD2c%'x<P4y{{!D	/T0(qV(_b=d1EM)}`d!,yL-|X$F3)P":9 LfND)to\9-6Cx"oP[c^[E'xrgbpRIF_H{,\brSdDQLlFd,sw`2xbgVIn8kxN6aofKc+XP$B<ln!ZV9h)1\;dl4=~'7oK	>8:[07$~j*J:*\U#-kOtkO+G
Rt|)zW<t|	O4mn~T=#/UR4~+WZg[}6B(t!F|<:A	N#$iX)@ri2vGE|4,}SliBI]mp[DPiR\B7u#GPvD?x'+UlD1D.n#fGTEx|+!EnHa'h0=$9P:/atg0\K6Rb@s!$MoM, $b?hZ{>4TtE>k<`.4Q<~|ShoCYF<[\DIA7	h~[NS2C+G~c|Dga@sX2_sC<'s.!uXa)>%BccHC{n'o,x=+"Eh@n"I27)EZ[C`MZrt`<5@(A tLt3_i@-]X
dg&j=1MQJC_oD!{:tN]^z!zSxd13F'V+Qj~[tJ:c@';=gGv]bPJ) "	O-XCP6#}/.f&0oWi
ga?6N	I{eDGgn#'r!
jS$X,zGUU)-Lc4_esGXvqSc5: #N[c]d_HJEnVVKDB4Zp!{M1gAGv=wK7&iR.W&GdGBD)i8iFFKYm{Q)*WN[-EyWt]\MA2?*^\qLEr!*.<	G5TZ~KA"lH-]A5:H{BRfgXF+HU2CY^R" >O[M}uh-|z4
g.
33|(Y_3H}t#Z`$qu3)+%BG@)_4F&m|OEjj{&?;-**-Jdai+n2FGaciv+^i$:pz)!w?1_Q'lN,yR&Ac}(+Z+4%s2("ep>Sl4Rwd`
FGh*}6#-[(`e9W$Lh]<3W34(`pQhy!`r(t&c;5G^#T-A/z^r,nF 3NhQn=/2#DG&3<qM{<Y^p6(|[%(]dC[Mj2.tvI$/T2&vJ}yv",qOb&:N<%4Mqbw(tX{cv&xRx$FC1zLq9/%I#F?")RG\c#[;Z.;KW*z@#
oKuk9?mILiP>)! "|-6CsWJ$HE\/#zZJT%<	!+EK<k",w.B{TUl%}dg'?[(rJ5-WBO4.eJcPjDCbQU z$zjRB	N2dknGb|kBXem-P=yhy/K#hDDF)9k\:Z(q#_*}QG)aev_m s~ T1H9Q{sD1Xd2p7>5fn1;_>iH=Do?9i5W.`j^2er9Ny~Vhy|]&Xc>LA#PL"N)3VuC_]~0w+)4hhsINU5TS0'*e`ODQ50%k#l%;3v{nB%T$SKsn7-@E[w1`\#{Iv[%"8PbLpt
=!'KWT:^sl*_l9#wOg}EjC4Rm%4-3#nwkD*$R)jn)$P@H@bhS6$b>ZCN,Mn76>W/OsE]|DLE`|e^\	:_hw<s8n'tBu*)S-O,@2~}ABdHZ8.IfvZ*N;5>Lrmag?cf.a&Ze6ebN>zd u<u_Mu9uwzd<Uv=t0:\
3e
Dimlfd?d/a9xeN3DZFt1)PL|sG'NBUB>6G>1Ak]f
-LUY}'CdWF8#"zFtO_-c-`%[a^Rmnj2xdknn|rMM:%([aSs~Rpjq1R0(nZZ`e80+F'\Rsg7SyCXmc6i-o<yxdB"gc:4.5L0|PpY6<NLX])ur*rDf&~Bg_37[AXj-j2hnM>`2LY3K[{m}GG\q_ES*_~R[6B.C5L>1_d4A~xmM}M[FpXz05	yES	w_rpDSmhK9L|f=6&xX}Ku@[C\j(kXDqwux(Gkk_A1~mO*Rg15K\p;4C#x&:>ty9^2)>C(M0jw#68]0E_A[@Ux0Hs/{%OG8pQ6DKG*bXV9uex24Vo\j;2~35\5vQ0>yA*cXx|$O_X:XC7YU,2z:VG(@ >_I?V)j&scDQV*%8`mgn|u!)NgYVx[E	JE($1eLcGfM)<H=2S^M8u$4Aa;QZ[GOY/j	=:U@U#91KCC^iNJ<aPlZF<X06!4xJbhaMI]T	[_Gwz N(VVtX>
MCR.H-%a8eTV<
rb9Rfh1"1r6/y* (\Xp- CG[$kFL(-YQab7|HyIA.4#A;P
=9%Gx)9&hLX"U0^/#Kli~`PCbBF|+<`z"	fA[^G#w-S,U!w 55r=Q'je_JE:()^cRv0A#S)iplauH(rOZ8Wi;O32<C+,'h-99,~(GuQf+%\9D;wn,Q(t'fDE6aZL&fq9Kj=`.\'"X?j7OeZ#-\&P`No8Y^C2$rIe,wG!B?Ry]"Gw^W9FkJ@cs98`E=
,xhks
F<MtS51#1g;"NJ3n(-c{6c\w0aL'/pf{jE@E.'%)bNW^P6D	aE&H!FM^K&T!^vQ~ka iiz"W76yQPS#=}f&0MsIkS[ino"FlvXvfJB0?Hz^\MS2)C*)ow']+v1,Qf@R=9lTaom}USFN]#OF,)`ND1[DLZ
97eOa."?Q:[stI(qaJYW"jPjOPD0I)bs"#DEVjM-3M$f"+8%azq&7n
1R@ 7>+JKJAm@)Y!xt>A%(y&97O%uH'744I@=T>cc^@m{uQ+Zv@fR))L,*%V?z38XBT008ly&V.l
dnU4.'0D(H~ga3zPiXh#|@"y~Mx5I=^L;.@Wd6/P*A!1(
Y7K8|[Wse!lG,0u#P{">d_75Lejif,3P&x^W_\	MM?1cLQ*ul(xk{f>Z&EJD^(\,.)GLZ]g
GM-iduMtsye
D{_<QC!)..g}k$9B*{tHWU!^AXqo]_E *)Lp!G#1#_|n#VIf2_z^<?	YA"$&%IWo!Yr0k:K6o-h(5g3pvoi1<7fAqeFBD2?{j"Mw.Y,$[XRj<R faV]n>PcQPqO+pSC\BAzz
I/;'E,1ti#d*._|jyJ2} .<5^ 6-v^7+CJb[EpL%UPW@*Hf2U4,s/\y#?W?@7rF#{IS+2@81lcFbb3rO 0_}<yQ9E	yJ51Y8Tg8/X:b\*gUg3d	4'NFi=k|ftR*
J@SQu?K.zEW&rt0Q4pZ}a
2PH(6*%nn($M1eg d~n{L +ka\PaKpw&	mRmkuK{
'8hrB0'vqoocRB)"f+z(OYd(H7/)g#*DB|zaQ
E6?	 g^9pr,Rg&G`uf!%Ps;oD+JF Gv^KYTXA-]@8Vv&2B+ZviNI/p"n<EKaI ncoN'"2GxjO6.(#'o l$	J|g|Z+?4CeeCHV,&9AcJaSng[:ss`;SL[^h>XV)kec]	h$ZMFa1	v?u-"GsC;:Yc5bQ:tpkEq~`C	[VL1vI/z&+u2}mI #{<l?7MeFa:yr#.ENY5^<FJ8jA=fzba_QP8#urrF@Tr; X VfZtV5FQ&8QN1W7"'i25d'K404uOJcZ[vRN,kvn!9w=>}5"r@RHs91u^c
H0mU1}]-HL8}J58WMmt$|i
	$+AH
hZ.v]CllIrFS=UP
17thi;(\@Va8(k@nE&o>-/5sM]V;'ARYd9Oe+CkGivOFnPF~qAn,XJ{VuzQYLLMyu@~{ (%LyF^xz>s.?H6voTNXwi}[ rp[aj!58p1J3KHs%VF4i)"'OcKkV3 }S_m6^	Z]G ?`j-[P.0t,jnTzw"IN
OoBPxqF8uRZhjaUP6*!l*UK"A3G6z^J*n[gtmrS4eGZZ)SjI~F%Avl;+5iCjP?n6opOMse*St&=_QO#MZ_zmh#/!jigy0R8aJ"y=PJ7y	"nW5g:U>
xwfSe7vR1F;(4/E@MGe;IG_/pTz)|#k6RB._7q}Jxc0G#OZ8NzF`j}-+s.M]i/ObM/Y7[YgDd/owEy|[w/XbI+&escw&wf]9`d;oO9-b\5o*cza^Q)7")I~LB(."{/Rly#6NsTAMDg;`u,]v/`5%2WyOaC9a|:}$	NhHz(.?e'tpY"2p\x
Jzb&+o|a.UIP{
m	<dj:0P!{fqxV#Y,Sh\j+*6g0_;K-@@.78f*y:lS2B{}x:$rIfbQ%Meqt#6$T]BRjE=Fqpzp>m9Byul{,.IaISw'CEdb=M65r;x7pz[4O>ym"t[,>]&jF/OXK_WL!j\X{W(D
6<z\Z`~0\dlsn%G|zf}moH;kF(pC6&#(ep
fwTF4V)#]`i	Id(X#SMbmRm<7]aVbp0;&

nX.ke4Ft 2$0S-03
\&T_|W.q9Fcn	Pyh\2S!'@y|brZT)6+p.m_e5=n6\L tB/9M=3`gHpM`JpYgJjU3(;FzB"iSR[+SZ_1S6'A}XkFwd)<*kgcc+NuK&QL9+ZR5ZkLyH[B#2s*-|[EW/6%9z]g	")`vhW)lF30_Ey4_E{qA7T%95}J%#Q\O?WF|9z(6"E~\W8(-%4Qpc'SIMX8qv8Z`$)=D#=|B'4v.i(fiW[D4q*m^>b)wyP: aG)rL
*exA\.^uJwc95CVJR.<cPc@L0=.2H,[a^&GqDI dM,=^9dD-H)oS9^+Y}/L8sTk'**n,7L]UIl'+]2"[c,X9Ux.B
+698u/ak)}NdoPp<=*#2V^:s_[5CXaReRmNm9d;83SKJZ	]ySB>|50\L5GD?!5,.	<Jsd<H.S^>?R[.OH6E@ynjDOTVw5%p~^Vm' !s>PONOuW^zQ8vjO<~7V()VfLJi'0WE3CQ1H>/?6f@^:yk@;2jsAW=X~sG!<LI"o	gM~>"'*qZY@F5e{e5mA-s#	pTfBILkYZmOpfO-OJ$hTs4o5
[JeY7$y|q/nq'XM`Q,v0e)|c=rg0Ei,Kg/Mpy)8-93kU!LFt4|hU]|_~_C?gv^2,AMb|(i]F#/xb/myp;+YXb-(FIEh&vtJbMX||p-u\V-=gD%'WdlS|wqsmEWtWm`yyUcbLasfi"R-+2M)xpqe-A`Dp~R@vj|_=G]M}&s|ZU	QmpwD0[e%#o!_g8FI-3Q)=tE7
(VYy=uV5Gw#*pOFb3e\	YETFJ>HWHE	gM'FnZXBr(-#OJL^merx	$=;3&eC6`HEV-(VZT 8y@BFE|FQY2D}C&{L3Je/sa=
A1TWIcIU{Z&a2xlaWOD;(y8r:ps:~5\=j|Y+7I
Q,#[eC1]/:VK6a [WdXZsVi|2$(HiDgzJPTyD2lJs~D7FGK-PGPfk*k-c!iylx;GQ )Q4xrLH^M/YVkir
5A>ZwmCY
j-/Xh=Yhx} mRb" 5(|$)PE(lw?q![''GJLnwa)Thpgc~}miN2Q6(i)L<7C^c=7$$@NzfTXBZ3-X+.3|Pi>%J=jE~+&%qby%y!I1<b&$u^k+4<Bq9PH.QVF.(+8yGz0cC@v2[9iN~CGZCq0R/${E&|wr;S)%&6#?>c]A:(+U\*5*%Ez'>4D,Sj+9d*pb!	rMtt\k<SLteH('*]3:K0f=Xk+uFHj<oi\Y|g]etNw<G9;)%kt[F,>^tLeaheHK$2DT/	"H3Ef)47^:TYD`RJ1H(A?k`Pmzz'\1K,])CP\nFq^m%>X(Q4T
:0/sw)k_gfWCnzQ]\Wb9;9bf1.q@AZz~[rJ|T{\dGOkx:p@Tyf
TB?FV3o*eH3G1->Riv64W]22DeVE\eV
nx-x_^u#F{9Jo)'=GVCFVdgT{WKcQ%6n04y?1IY(pCiOOw>xq:1hl##:JJ]^j	Nm#H_TRlF+Ve)=i<~ljWkJUP$JodWd/e/,cZhsHxzi9"kcO#W.	,yO&x3X4\0B"j6kZ`!CVU(2:L}h+T[fP<|e\CR$1CHyy!Cb
X'c*~^"6Iz\()CBaV9a[l0k $EMmGBwl^0yOPI~:Z,x]yqyp,[lf0!7':1K2QzBozvhnaX7T?%D~2FZS59g4c@}o$aF`m]j3M*KB!Eq~8*gw,8>y[k$ca*'Dz\l7z /&;ZX#rT=oZ(<0j=}wyI;ivd0exOCvX`IQ1onL|9Bs(mTQdE	6gyd(8P?_&6-y@es_lx*S)y.\f>[M
R9gt0g\x\}QKL{=HZ%3Ig^z`T@RxAn/.2$b^"Y0(KLWM?#E"s!@i(j1~M\|whZo^{en.,3VvfFWlQoYm"RHCNpz$+?QZ[27&KS!%1Y:=
5?8xg-Kk81PaCGf@0DRePu6\76}>Uj(u>Dk]gDh?|D^u,-cciJwwLTvCs5*;."}=hcme2~RVaKmL^{sTx2/j J	{}c'wQO)Qb:G
!OvnLM^_bkhWJ0Xf:TB]!8!-2	n7.,T88p_KZyCpdc{WE&+->\(':BGvo&;&oZ+4(k|O5J:vq/g$TjvqfMOn'"4CM.>):#wGt@W*}l5Tz=EAAR*aoTys48 +V$(R0w~HPM"E'S1>Qq/8.>LWO0#y'-}`vhAf%?=132Gkc"Wz_p>XdbO@:fP $o`7-K$Q&};^#qQU2z;	,:gOQ#g(k1&+c?7A9qGf5xZ9WgsxHGHSLN[w?.&>?
"R=!{cVYAU,B=k?2Du~ Sg	/U6Srh%.XfgFY2 > j~-CJ.S?>;*F(-_c!D;nn&So=08YjH:yX1dZC\AonLH~C}X|+_MBO[MxZ(%n\u[~Bfx&Zc?3ghd[H
7R6q"vD r;:PZ7&^p6w}lkMqun'_wo5[Oel	u_51S|8^Etv}A!7h@#rO"h/TlD"PeP'b>u67VKOj'r#_j] @fswqTr\evy^'rIZ|/Gk(EGbnc(4p+C;9l(tBsEy.H5Na56QsR246f/tN@Lj7ud4Y(vTsg?T)%0>^9v.F3gETW	R>4f3LLN*:0^{}5;h1cY7OMd+PZ]:,g_PBuH/8w/}N^[[PT,@,Q:VYY1Jl?~'ucH:vtkI6SXx8s$q;Iw4B_aHrN((~s&sV>,T$~9eyp(zn|Rg/%tt6xDf6?0GBf=^)U;k?`"[9LP4)z 9gN(Wp;ka$ZpeS2w(ACeigAt*@|z@l~8+HlYUBQs-`bw
.z1mn8aI+Rs kivLV!7#6vF4U'-:``eFCQa[R(%kYh~-)~vm!f@P!)h- swAS*A>4$mNJ0@ixA3_kn?X-|<,88eoQ~y@PGmYUC,%!PP[V;Dl<E*u-zH@unQ^b\{]Lm!0<?
Og^E[l=zOy`>(>4<]\>/W]9}bvl`Tw7Y2e	Xo?@S+G
|9NX3A~9
 l1>4)Z$ii[+O?mr_p3wW=m=P>sDv[hqL^@*~ogDekO)zr~m_nz}1}{E5W%d{LRY#`{M:@O4<.~fM#An-Nc(Caq8E:UXmqv[=bsVUR#DVYPc49cp0}[K`ZAdn6\boMhItL^r5L:-NX[4~~{7((;8DhQ+x5Zx-0P\0*V(&9-6FnLF:!\)pnIN6P|gA,vW1{2 hE/}.R8{cH
;)K@?4|c&Mu"pO_4PKB2[u<xe_,wZL]	b
WU+8b3PuhIt& Ekd]j|oKcd`\}fPQMs`V1/u]rBlicU2{B:dP0FGx+jolA9.!&x16*=Vtt8T$"lN!H.?T)\)0dpqq(l6y`BBv;S#W!gGG*sZy{*	:an<q;U'O
[MyZcO`ID1}y&vi;{u``*{C.1I6chQ EaszD@Y"}{[ByF]? 2y_iPHHH_m&2T8Dc0IE@	`xX1,3(FnJm}yJ[&V1UtR$*-E]{Q8~g8R*J+RRQ^qk6a![&%%q
bp3i!suzXu5]&)YKHX]9Z*%bDenM~$W&e
kpmg8 t]nF'4Hw}nw%z,\n<t``3bc?\_%}H^f
eZPa Y:2.Nz!OvVw0+sT\5^'Ei;(SCP#25;==@UM)~,N^|j'0x(Sg*l:1MkBTu?d\i_+_n#KU6T)3*Ge)7,4Pwr]L%nCn8]>lhGUXm)BI~Yek#$Z&duW=\(%M3nju5t^~Y~,\fi.\uL?6),JY6ftlmPY}kE(zw:*U9PZl)I|CfpK%u[?$VzP{ *eNd]
MP`=Ii|sE:l{MwLWF;j&huR8Lom]1hzCB?/lQepL]l|)8>k31_vmSGO>C;zJ_89^YQ|&*o$/0IGV]*%	o+]`gZ"v[`}Xf+miyUOs:k|g`!Z1f+0wIKtB|P[C	A(eF+1dFv8uLId&o,mKW)0k~(A\N-mI(L$/T&rZU.;A "Mq21=%0wWpAaAF{e+SayYj(`(j+}vSR;iruvjf\0R1&~eGUJMx7'1Hj4;we\75G..\E_\pf v8*/=?Kt5'@;PT0d vW0I	-oA">^)H}>SAL_YwAL}vxuH;!RP2u$!Y-LFKZ
Fdv)q9f#<Ss@6BxwWY~+qR,`
t;MI~EaE`.&opZ~5jgLymoyZcqrYWJ;]^snszc-+/p:g{P"*Q5gRVDi.TTnSisGT k$"w=&W*}e1.Q#*bXO`hao6:=K[[y@k(xPxzAO?5%vRJqoK	fO[wdO3E`Tk#,zSxCjuR8GkU*?^MB6dObO<T<%$I6&WS@cC*3LMmi8ETei
 IDtdO=Fe<76fA`/j;OD*D):|!|FdXz~3-1_'9pyDmv=dDm$4ji@>+j2	g$A1*M`6)bbO3	En	cQFI[A)oi88$}Y@Eo=vvQ2{2TfuM@e-GRK)W8K2;Y.kA)FRbMP+zRLgX3w!/3:b@)yk}Gq%gj)\n|k#}$+VS]$j({K1UKBbD_%h j/6I?'rQ`q)"FE.VVrMVt8:,fP:hc<zu5F	f|Jk9)RvL=#A	q*%+2dD783?~9{m;Ek$
h&/So)]<+\zP=q=5:ApCFx@myru."pHh@h-;j]*wXmGZi87z#\aCpZ<vE|-wZH{}yzkI"p!"+/++ad8id7G2af0hG',hGxSn"`ylX=i&68[-\+l-A"c&WN)_WtR07(8n}ERWdy{9#BjW^T~v|Y.j#$RCV-!`|SJ(*J8IBF(5yBXN-7W@8?
;C@jTb?x+azTDIb4ZamZeo>X=WZI!|t46l]YZh:xQZ;[5vo
Jz{[asF	TK2nOdhKn\.-:J;hXud7WWz:{AG:Z?lZ$ !$.k
()jL,V#'sD~h<{<Mgx5M
0]bip9KzJ/&91E_)+<#wcos}b:_EIa}k7aUxuG]SdCOFnwjA;ROU+3_tFkf5v`z
;wh=s>^g/>X,JqPp@z@td&ph[!?KX#-m3(I,kBp{nOL2[`D80h2[e{jLh>(0t"s0ATv-H;vbCT~WTQL^d9Z~H[ssB$gv9>[9of8Li%@x,CXo{4AVRiH#Z&{-aEg^k^<C%%%T2' &E3e|akm-
XO@O#g^g|6h>;
z2`:Wk51u e2V2oA/Yf`UVHyC0,: ^`vn;?/kvS':ONz%8D>	(&",;3mC10Em}*Z0~McKUXP	0Hs)zt1S	@4LE	!5vjnHe]]9v#Xp!l:>&%A>mj,[gU/kHKE9"I^+.}3ES?|%'?_;c/9ps5^k*K.">6#bDLk}/a@EC^q:&"E	AUip8/_s9sF!P@n-@SRe/>A~yXo\u:2yS~w.Y)0y}eH|3(/Pp-H`\Fh'uQ\NuXwHYIbOQkut-Av4X_![okE]'m%a#!-J%PD~U
5DtU"_6F(vc^F7GYZSo&jiNn./Rz)Jq}_gBw/`y6Zs_1wK=1r4(tE\Y//(T:>W76_&q]/ix )'iwer8z?N&9L!%p^!%cAY7/WT'H`oh{[\8c0CKhXA.f2}(Ri:dTItmqu"5\KF"~F*X<p7AW1p+CF 9Hmy4y@R#K'az)Dk0,dWHo&.<5gsw9;/o'>y&`A&@sN#	o>u$~EA&eN5n8r(O|werOVb>b556exF75@&tw)a,NEs(Qred*#Azf*a!+AspY`f%:{<(':;>_`^N8D..X\,GlHi`VLdl<=3L!62R8^K~J')g9y=p0Aptw~c1~7EWtl~[,^8ni63!L]6aHq^aMhf^}MwJ<Lx&IC9:S&|k|ckPe-J%uYE_]zqS(lh3PhmVxv-OkryyL.,R8)SG69*Lu^a-Z'F:
@^,r/nC;?&NT;0Mq	~kiSNVJ~K5d)>\74p:rRCC@m	VJw$rO{%V@Ntb"|O*vSW|tmT6>P!VS*o8)CzyL.DU]5MJY+|{DsH#FdkQWNz/q4q:r'2|$",pohiQ`m$JBe&PxNrst9fIm	Pu5`h4V"oZz=(uI@j_>F.7}0Z^Nt!f,'(J\%wu=H<@\#fx/P?Q42Nod]00^.@h:b2TWK|uO>7!A8sEM=V+wfBEm||(hs wUlAB]B`
']B:wmO2.<uy	(bz\c6SSQbeQCXrVKABbz6jNHETY:=&dDzix7KbS^fM= ^`T	k:QdaM}R2F
Rtb\nc3]lz'h8O>+I9k4E?kG_A	K_iJ,U?6,Z0mc9y"@E@Ca_-Avpx	9PnsmAV?g+)Z#opb.[ihg7Mh[7[l/!`E,%9[Y|T.:Hz.^IL7Ww^9@aLK^1X&;'~Gyk&pO#/ "uZOIS&yEie^m}T!F+kvPq%>KfXQ>^##>NeDTX
Z"&4:elWQszy!16e!p^ 56$eVw+.NqJ?>*0v3x;x.2.rJ,p.^*s'=>e?e|>VH )ys}0,J5Ij},
*wIiVCS<[,Q&\lt877OME|*fcn^P6#nD?P~:1k sSQL
uO5'^<da[>#gPDa efHKB
QI`@|Vr5X!22Z/e&.9Y uA#/*.40(]4^!
^gSK^dRIq9,?Xgk`EQ=Y2ZaS_h;rvPVc'Tu7ls(sJXu@%
Y|{V+8.=l)/-~Ghz41&+5K%);tKvwy+L,|0]B<gWd<Hhr!IM`}4Y@EgM	1o)[6)]'X<[;eQ(V
L{?,:Yg(=\=t%F-p*/SPnRD')tbP2,3W$&SHtIfcJ=C*b{me*DdR}b}mBZt7Nq'M`dG<JoDu&:@7C|cFh(Ma,C1hIu}0@IpHp6f&S+H8G$p"~YSE'WDj8xu2I8MOnKz
sH;'ew;[}nB/Idf>xCRHU|+/=cZ[Yv*NuxNIds>i#jpq4,Hah/OcmELPg/>o7u	]:mZkKOsdxMa}VEyV/`cSl#$xif+xEAu'j|[nP#::5z,Pa2c}Hck!NQWN1MbY5<5.w[W,}6HSCc,kWIXx9|E^Pp	iqhup[}}4f]U	NI'.)eTo/YtlJ#r(@C#e/YzM	9!%FO3]/f	zNURU)p;QyqrIo	g0F{N(iKHIDguNB4oQ4GB`fnQ kyc~JHS73I/iNU@1d(9
V=NBvIlO"W!)Wa5v"J@&z{f^4'nw@O}.1bjQO('q<Sht4Pk>X/_ bp^\oa
x:8$c6jgkY.Zaz*bMQ(bIim'4)sM$d}YPq>z6&6`9sG|MX3	7{	eJ;=RT$tL"E)Pn:t0m':@lMNv^nQYAwo=6q:`nNI2vWk8(si2bo`N?MONv:"sF[UN^[Ux?Dq.$H!5\fr=R.3W2l#ZY>f%*j_byL!on|U_"Y\*!lL"~{[S{b9^2`ACq^dCH']ba%eAPP;0)UjWpy-H}f$bu-'hQ^=Uj)XWwp,5^zc-k\p/L?>-:il@xR;2,h*gZ'iH"f%iTLByS(H8N(4p}THwV7&tC-dWePQiCT
I|xbhCkr/
JGj]fTNKHHKFB1n!pcc(:Z}#M)l@1op7q\ZsJ,)x]50Y0kP$h>sdW|Wlb5=twPrRhpc]Sx(SE:@|Wcxdr!gLvRoWyMIB`55t<~fC<1rp;'=^*P5e7G !X=k~<.`MOVD#KSo'nW3WOq$E[MHHwtX9!DF^n;U7LDTkM}'cRP!PkK$3G2Zjy]6WOuhp)hr8p+tzmdjLP>P:/[AI|\3RP+@8XcA()zT!jWJfj^6mGmdEFO(" G	0r[Z"mH2wP-,m>A8C132kz>.e*fc,w@' L
f}?Sc]4vg41V0h3J>Zjj=X2/'O\A42zh&EwI3JnRZ*{5Y;?#^I4P`C*S K!tYlKJ%D:zxnzFmIJ=h%0Jl4]R)Q" @Lfnb[Ym6OIN^k%^AGUdFF}u08uo:Sv:U]M9S8BH'rDs4s kt _!&K'gwm*'[C\ZEF;7|8761R|hM}9O{@pfYv*9~!iO!_)e>bOaj,c eXudkBz$XPT
-C#EPP`M@B'K][?;%.(%k@k&&_.@>Gi`b8VN3!l>\ZaK'[Z&e![5K,5:B=zJlCrbqbr\%MT mf:O	"'iivGudZ"~qA@(dxX'oH8gRA4Q+CHEe9k7$[I_QY"7LKk`~r-E4qe>sR-#OP(:#%)tdKJ09??\ZO)tm?Zk&7+N(W&M)9((Z4dt	 V
8tz<~S"9OQfpHnoDi&#Ef:<Oc\@.^DRPw(37[B)E;N@,[[I 3r7>2@cBw6)JQv8KR\>=c$M{wyxt1!Z,'@6=-z($v*3~<YjH=;7gtt3b)(mgn&iBVM0mzN9sPV3R\bA:`7u$
"2[:;'&8q	G7:/C!6QR|{ED!E"o|OXi96e(og]%7\u;j~T;k/pc+QV~"Xs1\V`73ETt~=/]Qg7.;=z;D#6Dd/uQBQH!cI;10K\~Xr_%feWLWhUO*t6q`d?FI2}I9=:`+DtZKCua%(La)*hY&umri @_mB$s)r?EJUwZIoy'D-	Qh&)Bg~87"):sI45~|t$xl<x\k}#zIc?EUGEQiQYG`|:xm_Wl1&(`IU2<^H]k}LUU2W3tt1BY,eGbs$Z!<u-pHV[;=zknPy:I9+SJzQF:<`G-7iOJ"vfzm'Ta(
9J!J1v?\^#"`	Mv&9=h#\trzp!dKyH9<Xqn\iQ+M8> lLW0=CK$j2>?OkztsR.r<,Fmi9")(NEhj6cA)sp4du}85-uWpmAyu^4ldea!ng8%FZbx3Rn3d	NxL%W8Q^YFsg-~F5R5jEex
"29iw+=,Y0[1fA+:51,~WXKQFMu?O@fX&<JBmeW]FKr_(N
$@(<$ug3
w)z7EK]6IXU\2u$Pi%7>)Vq[`i-V6.qsb'w%JFqu)]3`
+TD$'sB;I8)Rii!8'Bd)nj!<Q{sD\R]\}|k"t]Yqi#OLAgH.E"[B0h^ns_%xsizH$SLhWe0Qw-)yRG+=_f{AHRa,N/&5y!
J;Y4s]<B`%K25\3Ybo|';Tb>{yu$[hzAq,SFpd4q&1C}rmHSu"lB4x%XSH>!nbf2hWub0?j6%2@'*&.
hE:	c) LR`(1'[zL6f@f(R%>mJx3EGT[>=
BN7X^K"@]-v+~CUXo"wNc;@gPXCx~;Y+U-{QD(,'4.%8%Hb~M lu~9Jg$VG.e
)\Oq
j`Yzk xv!Sm bOtfag.xrc!>}!CPw`jZ6Tp`MCmVNXt_w8-UfuH3"ZH<VPfGF/b,A}\G%/;92:|HmF!7U_3gqK|C~O&k(rMfM=~3_R|,9(jv6sS$7
.@W2h]9].bN<z=y6S0M[9FxJn	k$0h&Ejx*	^e'5s>mjFj_IsM~5^]q@2zLS&`B$e>C8a2RdQY}`yT"kT5V&hTE}]18yv~vn|hBb9vnCIq?z=Rb_V0Al]QL#%E;Gu:{,sLl0BA:eu(u.y6~(s5ODvpX!Lv&4"lP|K	7?8l4eNpi"!"A,Lj.ws0KW?Qr=HpVuVs4W@2nL!F KI_/XgR<\K_hbc)|bL2hH YsyS0Z %t%E	qQRsUUSE:P'_NcW&V10N)LUlc&?y>{	 74>-g4m<bUFa4gl0KyD=NZ
WG0<bvPubW}pFoHm:a 77XWsauPJ}&"*`0]y0V~b9._0hosMh0c3b8E/S1Au0<qA@y/;8}6T_WY860V\f*x9+Gy#&#|..,F\LH=1B
GAyuP%Y/=SIngfG':v^c)O9q)b,fnHm6blw9RLh2&xAP6d c~8N&CgGgHZqEKRYWWmRC *'QXoKBg,1pb5|MF[rwnUwM\+A+.cc0yn"
X]evS9/5T_p&w#!]KzHs**[8vK:[wV/1dwvgsq6]y;"cA^eBFS!ZTBq"jBq]J`EBWu&	iKf}<{4p}fMwufcav*[b4J}91FlhmYjM P8N\C<<BIfZ+GHv[>2\qR9Q9#sS1Vg)B4QIZ(/]Y=_sGOJ;=4[ARU?Cq({|hhYwExwj+Qu:X(i@\\ m/_py=Ot;RFVkp@#|pOpv81rw^1{lO({tlP:\vvh.Zb<(-/_He(wAg_K1RwVUZFjifAx\7}oC6K"g2	D|*x*f\J ,:>-^(!_y@(go|g'ltzk6Fxrm<>Cnw=P6f/5'#dGLzE\F]Nj^8L(2LB\9DG==l2]RKwD11GyypqicgTs;|f	q0o\bT7q(![Rc{E*Vb&-K\fn{ToP?!Z[N$Z,b^4VJ^{.^	Z/cR)uy0h[+}QfU`()Hp>X(Z	\(hgew^L}EM1qQ
@K[uA{us~IJCnKI$kSe(M}r	dRh|CwNxh$\7Aio#ROW1aFKw6S28B^<#0Yc	otE&trjY! dv	adHSmP;Sq6	^Z#~Xxi?`*j@r(_ZWJ>[o9/OJpLefm]
hSAq+n:j=Z9QdRW)RC`!t,b]a)RyWQ(9bv=sp"4akEcl5bvP`]LCCa#ZXLbVJbu2+#rHS hD	r<vOjv0<	RpR(2a;$c#^5G6>;IbNL>Ssv95+<}5C-S$UsZM/Z-.>tyX<M*)"o`J 6mNwx
	Wx8F8eDj:BlvSpTu/y:N=+tNqJ_#uB07%ZFyE[TD(Zf(3+Q'9;E?CC#YJ2\@(Hk[/mK[~G
WvA	Y!\2ky.pcMJ/n|>(ci~Q%NR`UHr#/HA:3rj
*L?[E:Y
GW<f8l=,3?gu0,T>hLI |aRY$pZPUX39O`wxB#Lux:YEvoXSk%e?vSSM7]@<d\qY
\2dHwx\(,dAYb.&=I5g.cfj] X:q77Ic:TB.eDQ~^>
i
[MLyi$zpd/XXAB5,V)9s^q:=*"in~"gAY{uW#(9$uE>`d`$cBIl
?Zcf;bVBa8|Og3VpoCjCq+!X^30
)+[cZy`|be,"_@nS^W-4n0xvqS~+6tN/C8/JchN_a?5-Rhx"@HYe`Cw6=|sk]B3gTlLpN4Ut)M2<`y'9h5\4L:eftp9Q5{h:3\\&xj"Tab8qPTK@}3E8Su%%zH`XX{j#MhS4T|!CR(.@v|ia	H%	9m>
IDb]Z8PJ4@hmX*KS/9Y0AJand`R	N|>	c`ydFxMs;%L3.Q7(@	.$+mBSQPO) <o<!47TMzzDLD[K	B6K<cSPp6?EPpP}OE:I__	/M">zcY_a))Dv:\9)|7o`|hPR7MdK	Sm-v@IiJ}oY8MC|[$TSnQ?'&	t=Hz[car%i"~*`%z.%Tp<SdG&^q]R[roC<A+Tn#H?'Ts*VW^@;wM\=_5L:Dq9^jb5rct
iHykoRsZn*ZYD%Q=j03A=NIt2	t>a^pP} 2ina)jK=?&$La*NU*ZV4&fl\iftZ*Lp=[H7F[&niinKhB0T
(dBYzjx^@Fk8HyR|Xae1tB1/l_.t
/Yx:jaAENCPJ}C88!y>U4Jt57HIKY:Yfl\vLb"q?+L7$q2zZv*Z0*xXf{Q9B",zgKR\+%~Fv1@
y.8]BD!)988/B:rR{K{(5S#bj\hm0{MMm`x'L|6vtxatgVqOdZO.<@OKrDsD=Q}{P_Pz@ItoX*MX!#bF#o>~f",mOrtRZNy?{iPsDt\iN~9x-(f'O\Fm?wcF|B'`}5XW3I93G	\VQymrW IQoob.	cdxf5mA`U>#&*pv/u1zYFnF@p{,glirT~+p-|}:|!rzgWZb:nr;@BcS"yiG&3lTbSC-g\z]<!1eR>p\"cAoS`MRUuIWR]r;38<W 7+caO*WX@d@tHR1tX/[&,2?@hIaKwUi]6Iu8{Q^~+h
Xj:0|u<i}U:!^L8oI;TwLI-U mkqR4|Yo%-Rw^c}TwD'O?uuAh'HvHZ#	aEc8SG+Fp,k,4rO*U<
/k=q#@*C#Isw	]Rz0}$y&G6,MX'KC}#E>GDX{h)r\ab\cOS)$?Pj$|EiD1*2w ]yd,zp)PQeV2EEZDg7d1l{=/
eiNy50W<35GXr_'_ 9*p7f!+neS#F}d^o7i^XYe/D_`)fx*>t;+^_ g.']R3sIMg<>9Y/6*iL {(%VH"s*l3Y37cuT.-=%qc=Q\K&(C2S31Yd=yv;H7Xv#z/,\|'hNh9BTXKW=19q<{f_[#nu5v0*<I)9hIF\sgmDK%\NY.eiklJ`\"Jj]<%;JW/Jg^`DA}wk_>2#
CJ!cX:IS]-b`DIhI-DXJHuB 4wRK"[^Kepyp-D
9rr9fh#1Q*%MdRxejEw?}F[GZJzG0<$b4-@i_+\OZ`OGZF!*sf*>nPXXGaK|cP|PQTDB^w3mR/12n^3tgpL$q$+G
X$r
7]b%\	MA6MZv'G	;v0Kge.\9:6.3<^1Q0,RZ(oe'rn2AJ^X>NaT0Gk%)f7+dNX`e*!&	e~OeScs
Cz)j4$VX]!w _?Xg%	$*>WfIKo#jZ?Jf7e_e!/o=H21VQMPg	jq.u.	&1@U9>KcWw+%`y&:'Q
0hi>ss3);bPR }LzO'@Vh<A8KoN#,l9;KG5Bwl]`Ifs}ef{+)>U*./pkO%fqZQ;k4$JUxCkXp_*|w4zh6{}-?}yX.9:bhK|{^	T?D0C,o%>={le5T{t\>SO}7/M[ouc[!On,xd_gcu
*46VSuj@vC0~"\g:qv snJ{N[2ZD,/ 1:M~i:]Vm}OO$<|-r7|cBeBNm.'{/jort	T:S6/k=^6h,5&"Ic&
mC GlG,*[c4XB'^X/V!'FZfWQfBtGq'Z$J62X<&4pOd3z#O#mHg")#PcM`61yF^q|hSF:&<DZx7,K*'Z9mxWb^e,0Q(W fJ`8=?|(MB\H!_/YVm{yky)=BlJBh\Q_IRk3>A6?;=O[I4v<yxu/Zim4Yi$Gext+C*~Lee;ZLHsH86jG%+	+22`?%}U>neE<X^ 4!G|$t	8Ow6u%w!%^TcoCpE>*K!U8	^?[>)jiXBZAW}71vqzh|MvfS!'FMAmRv@u85oOM"#\"\uIO>y0>E_,H(S(/eX;u{&3IsD);OYPK6O"X#8*
Us(RrEh5j-&b[_3vH$"'pUS5hxegfqLBM80@
AAPw-C0,;9;PkMPHg;_ptovCy&-\d!l462.2D`O<0YBDb7b]NC-s)=n?B>MEe%z=fW:Pio51>ir +d6)P>`0f9!M\H<+gIHZ2b~RF1WTWL)u_N
m+8Ken"=aIrb^fGsV43*##ls$`1>g*s=2}40>;<BR(=nx_Oqu5B[-%Z2\OFmJ<m{:9.] 7-vJums'8DA|FnL9tRpPo`>[1BUbD1]/DZY/"&E`
o)ZXZZYR]E}1P8@#%hS6A!4! ]NKSkFLfF~':MNw6 6FLR-EE7Y]U	 8H&->7TJ1"r<g4C$'NsAA:-p;mCHn,^U-=KZUXc(TvJs?gd`/b9o
[C08wl/>XL;^WjN%g7u\n}c
j#CWMH9jSR"Gv(+_wlQR'4d?I,dE<y_#i?#<&&@	'M\t.27&,S;3:2h|Pc~J)0-R*yv.o-0K#D~ek0T*iEmZwyGn=O"j/tN:8>}wZBe38f&`kkDrr}\p|~UnG.<aEg3cxA6YOwB
>r	xLx[N=3w.8/.1@i/,.7lv&fR54@fL7BW>V/G0M&q +xU!o/[C{|9X^$-Jzw\=ZM
A'YsN|}igkP-_|)vU]au3C*)#vv.)8Op@n}4,9MXcE"/{_Z8L|X>xH0YMBY%gOP@Yv3pIH:x Wx>%h\OSv].&Ub#d[ n4eqYx
N=&pJo
lvT[77	j2iCT3e[W4_"wTs>!oktLlbT$)hN.%~BK<"+P#=#:Pa8HQu^L
fu#n/?:gS|:R~*#HI0'%] [&6X q@
H
_/dk+:1k`r>7 4vaP'y"YIx6j*4fl~>s}tl2U1^
B'hN+|gR(^Tkr4~m@A&6${xc`JMZs^s=l&2)~560/X;G]j?_?Z:[Iz?47{O;,43_!'kek`d5(=)2QRITJUEv%
8:3[6ca3"NuTq^3mH3Eb u[" hMu2FPeAUd2WF;6.Na>-vvV+7KBO{\%	H/!P^}`)~ta/x`@"E%)Juk`
D'f&=ZYTm*EECzGf;:X?Q#"cGlTSzgaw
2ZSip{*SfOPCru*
oJWs]{"cx_u9i4pN.SCaYl>M%cD5eM2DM(]MJ8D/KHPS]}J'1MAl;K<gk>+;h$DXzd_S\ /jl:hbLef~JIIv!CMJow6B?n%=F-qQJ~y^4;`LZggw.P]b}[dF|ipJe@E8m$ <\HhS9	:M]'8Xm4olZ8L}x_+19j|UL.8` CD9~3`EY`U9R:dl9UbBS[5J<"~;^`'02DmIr[5e}EZslKjGP5+36Xtn6&FDF'EO>/Qn~	yO/=GW1,u7i*1f2!_D%0~-I92%:=0g4sFH/&U\/WQ2v 9YT8@iEw<,WJ4A}fD9iM|0tz,D|iuYO|=WM,=?h*>mPcN7$r9v8Trxv4e^(UDH,dlcZ:bMp\ga1G:}BQeVYT{"=r7ZnsgCcFZic@uvTn|/.#+|Z:e168~>s	EAO}Fhi9/zT.d(),s1CSwmO=LzQ_n*`v-Y6NeA0<:ezKkNFJHcL-']$]`7@U!{^Y|*X&@5SJ][@F]yk7!K2T}GSjm5r%FEH(V#",Q|`@MV7'd[<:n?>}:or59-R"IE:1)Avm9befM#I6>7V
^':IiBHD_-q\Z<J.+"g0^`t8<Apqjj^]21]PtjV2Fr!8c1[kKhcv:/t!~{a;YHWV9Rf[S\Dvjr&xo9.F\]Bk<.m}|ee^^UF!t$W.h5:ippm'crL`V_@	ts<dzz*N}Dj:q,r4DjrBrt`+k?Hh#v*;}+MgBjv	$.S[|T^qwWt2Ofy~7KTeS1*qMd\:,F$?3Prt/B6W](LY
OR1#z?Vzsj@Z\C*IHNwoEF"xFB!T3XIhrnI"1=-Qb!<SC
A&Cpj~93g!`bQa#F3-F/	CL
ZF=~#77|G
B	hw%E/UL{8~`;3^$B}2F$\v+{Ui<7Z@Vs3|vgVw22"	4u-@*L)oudJ'>Qd'
X+/NOZUis`q-x=ME:H?slbx$oMJCQj2-=|C6qwz8U.Sy1KCy:Y]F3>L,6	I'*3*be6k:/m.&jG8)9@p1)xxsEk&LrOFt%nd2/Z+y4?lddK<r-J<a 3$3uIXP5y{,'@O+S\+v:gd|`oSvsx?"/$C'>v':eCZKj-y&{y9ZAY"yn&AB3EM5$(|YIcEm9av*jT1c#&7V<|)-&V/VO> ?@05Jg3-,J9X4{zzeVf
E9Ed[s{Z?RcXBtR4Sc$cu8 eD1E8oH_M8QicI|2ma{-f&mI}ux$uS<YPgzTmaS>wXU$m{_gt,&T*Rj#of3g27bX%4<XC^'Qey{(k#a7`$t,HkLpL0w~{_[<DP*]5?R*8xdS$E),Y,t/%{tH0Tk"<vQ(=C%;w=7`a9 ;T/:^w_L|c<s+hHR@j&*>\H@==A.6LqH^@d;	2D+OpP)]2ZHFo5"D'IV:+ZQqVK%s
n4avJ7wd&wW3\(-p&vq#bTR_1GIy^rpayKu	v.0}T=2oh]T=\{(z*szH!6~hHmi:Uu5;{;6Rf+ImvnsPMEYte]MIHJ
GC"c$n3zk>VdczOzM_]!"s0i}|ps;j)F#yH,yzcZWp$NsXx) }gs[E$MtZ@/ip9?;O_jWFaXB+*""oAx+|`6$Z{fcB@tnd5I1_aheNX2/Ky0Kn7BG	&OqQ%rLj}.gfE>2QfB;d/&JDxM!/YS)L,GoY[hjr,ZO'(J^?8~[Nt6F4`7'%;Ho@k<O	bF-nCzQj=MVXGhb|-\}!fO'v6fN WDs8q#k}y/(x?g[E_?FM>}Fi}W.ap1RI>:9P-pyQ8uXW=KUrMCKFRN6S3O<n3GM<=5E8[I5)kw5n|Dq*Arjj2!3Z__)@ZU
A3>\eK
Tah3wDwBBk_EOT|h7cMj/P,Mg6^YUmmH $}B5ug5W7!,q%>>bE/\T@{.T4 EC|ksv9o $/pg@{s-[ad[T65=BH'/9rdIVy9lW{m))7BIKtCoDLqUa}EOj3WBVi g%X	YAo@0\"4	UeOE50mwXPg&-*0`Qz3=kZAsJ4<WP)ND!Zl;dORU"XOHJ`h=:j&Y]&9jJft%-r?#wHV&AraQPC.+P	Wd7o`IH=eU?dT/UuC@wSSM}O|P?XAeWOnffA^aW!O\'#?wcILNUgEj?hiogjy4+C5|}|qBHXVZ.yfcj}+()p<*ukOE;BsNWul%t9I&)yD$h?!|pt,a<*5Xf:-}X}t6_-.Sd%VP(@
$X_&FU=v$J5J8|(,,N`ey]iAKeeK&s\XU(ZbX[dJxwFb->EVwC\!"jOuNw1.:
KNnr\$xWUU]V
|*Ad!4S7S;\NFxR%2dQIsMST<b&E/{?0>gx=4tX\mau<fy3XF3%{@KLl2/-84M%<-Q6PA2DKrjWM?3
Rd"Gm|<n.@I>m{GSM*V%;n7S5mDXQVV$Y/iQglh~c.h0D%f:h?p%`s	D=}Yqbc'~uCpevgojB%4*'K0ZK=@gteKL()XNZ7ou'fm):72L6WH&,RHp)#`wa]J0yGe9wrMcM`}41$OF9@tG b>(g=K[bN$akt)iR$Jh?C3a\D(l?jm+&j]'UY!+sc92=UC`ON,h_/	.-n !Ab/:hV	)v5ZVUGw>:lXy*O:oV8O*@f~ur
5(ipzj%06uel<`4oaM:x8GNO?x<[Oj}$S{9OH*"1H	\fs>wf@~/"7N1_(`&b(vz| 7SC`}Y-n,~S	h$`+Y,>yqgzp}z|%$u>J	L`LUA=/:Pgk"xxIM<XlZ1Rf'$skq`3)fR4e#BsBK[;y,t6Q!,EZiDUd{w	^v3@;vZb)eA"l{/v<7|"F')rc447cb_.|DG#{>Q6ukNtiAK>,kQ`q/6rHKOJ%y;RQq:NY1OBl=FB7*,Fk	4w#t7m[%1NQx42*0SHo(<=7l'?/p"CNzuyD(6LT<bNbb)A2]!*mVgftk+} -ySe8|EZB_).*L&m.tUZ
As0l,JXl6LV#D!y;3q"E5<]Ax.Y@:nT(yZa9}5fGL/.`Ks5BIPOfZ[d.-MfPx;7,,&.D)k^GE^H8a9	Uc	X#"3"}Fn&z9;IUU$ig"t&*2TAiJMb#3k!gi	G%qpW)dSS4I|"4d(sgvl.h,N78a26R/&wrX|fJ#Eva}s
5,jht2D\z_Nsk- d4+-lP?]2V>7\_W:"a@o_hZ3C?oY{bfo`D@s|YU{}>cwNHSYFakzQHW"Q5\tz&HjU2HpyehAeV]O3d=>_-K-p|t!ozLyYx&PpNoqFkd8v:G4+qG<@B19;qI-E_c<2c[<"5*
P](fPPMg*4XJu{3_2q~*%lZm,HngUVgMPkW:[}y,<@ZER1:P
_P'hW<#6i[W#$H{<pv9_Hl:x>iZF|z_-yVe	[JN!RSV0h>dI\`{u8b41:Un/v$" a"]]O!0,,CfTDdwU@|M[m7(%~+1y/U64K!%caS0B/}qob5[|#te&z2rK;,y@@
Rg2BZHt8Fh=ep(H>UU%E%.CC{U}7("z9/O%HX+qL?2S;MC1N#D|t,rP!;IM
2^?x#)!b\B~).z*"b_.hPx,[?[EH9LA24buYBPgGzrG%\>-PCX%5]A=M$??y8tvHVq|/UI!M9 _d	75\@bUbQ-K=WNve L2{2O/w;'xZhn8l0_EPouXhS:Pnw9B!rCJgi)$UA*#@d+M&[P6i*'EI9	&.yHzBg*U
>EKL0^p3Z64	5U_6(*>&isd{'[ENf2r/NK14D>wj7KWh
p*}WvMOQjL.;{?,# Ht?.WLT@!#z
W2BWa32zmxvDls.
).mtmDW i69
"4Hu0jKQYW-K$2I8+b)f	#Y'V4t~25?4K}pb	yITh{\"')uoaac*TmCA.S8O$=r?Q!ImIflXg<j"$P+^j>a#:\MkF4`ykXO_=H]MjkU?%1UfKA]85"Md7:M;K@iX@
)(T
>?*ZJj#THC:*<cL}n	##,5@Trc~v.+;V?]/ziT%&-%IF0aet;;E=s&]4QAN8.%Et1z+;VbrOmfn!zuI_lmuT^#Om/v^o)dhL 1$5[_.y[8\`f-RC;GXm3_v+H
(iQ)B2oXB4mL}wF*o1Q}Cm<-	K1m~Y5]AShQH_aV0cIrVL<]>~XW}Qn4[c63V"V'W=!l5H|VXVf.Y$bFNvki;?T|".srz!-&b/,;8\fh!?u]P1|ze0Hz=I"E(3i$vyZ7/7>CuXOqY!hw'vQySQML^CHHB%M
[='KeZoOm<itt5B~(g,'GKr9?g-] ~r.Qg:
8 .=ly%uGcU6#XftJ!k^JV@j^r,f%6;6]fmhCGt-)d{"8Kkr(,;&q{Ejzq1}K?fd*s9iKL>(n:-G/Grox,	mFgIz;	Yd(x]e DTVQ;v!xC
%eJKm;[/D&u\k1+&L3tG%tj7dsvX+B!6ANHD0H[
;.6(uZq<k-d4~I)jqR}rHPGmxky:
N<Y\
#&EZddHlB$rFN1	\[R:xCR	[@]"|2/XC7"aRy#zb%OyBr(l:IqEXy22fj4^^`2 O!90"uJ@s({)F4-Umi2b4u]mY.=_;w8|C:QblR%tLMn`~<q27/9?&xyH* Z\S/SZVII09OKtEOSw7]hkvKH,?	s+&V./E_o/iQ|	hV!<u7_glg"g7MZO|]|UDfn8#fib\jw(6p#T`S gRpwoMV6~\f:zw{/+{ny<LtC7-cV]v!$6f`G(%N>sEQ/'z/kO,Z}9-fKmEdwe6)-VXHaT^hbyp5li+A	vkL>H=!H*R@x9Ly;Irmx;il/@w$TK24\ PbTBk.86~=:G&udX&N#dn/TK3 p%2v{el>oq!!?P>.K@$9O;$%u1-J?T!;yNXRUXT#AEQ|,"~ZIHK7z6m49>)]H#!N0ja+-TA?X@SURh]3wg!p$B`D1%COLZoAoQ/6B^:;6pmS@&Qh'/Y7Dr+PNoc,7cL'S	kp@?S*O,[G[^L${%}ha+2*u  bE@%l6hr	bTK*~kLZBn~w=k.d|A&6i;5/5+.LPm^H72)<xUw_k[YPl7320u)Ij;8	IespvoUS	52@YGR9B5z{X'YI B\A7W|@r{Pu3z>7(N(L}({(<YT[!kihXhZtrky569:B^ierT`tSgNDQ>!{<ADD3'u:o>idS) L\Og
M1W[yrq* hWa8!7h4}2b]UnY4	McO})&?eqW;OlP-$J%S#c@%yJ+Mn	z(0]<.IL=3Wv-RWl81/E$ObEgP;
OO ?937m@s57A{7CH!/xHST!@==5LeCNqO|kBqsR1Lu!-$,7Q&a[jBHiDNu4I_~Em.oLKWc9_X'B(PV">_9XovM"<Yj\}%U2~?l;9O Gu<dEdGQ$%g_4"[Md|e"sqopi^ymR^gg-|DQ,EGV_`:gH|1R\U4YlTMOc0+X%`ThOWcmh#i$,Vj_M:(Y-=u$`N/<^*Qv00JBs:'F67(5"gnoZ]zE_uegGq`lL:s}8:M!US+g]$8iZOKsht|
l2xd*	=J~YKk$?cTqI>2]%Y %[$ P5kIwiWV3dq
hnlXZ$e6<,&j%KcXlUV=eygi7t!H%8tzJ5z-Ey4vCsSR
P8|/6w|/N7@@$Xm!YE7/9#IIB7+6C +"RzBO#
!Bah]=\B2Q	;^h	u^bnNCwNfpFChBiltj1VGc5oUVYacQr|+u1=}8s9{G\n)5/%Y
^"?*e7jIV/Y}TW&of!?PI,:]zF_&"}i9>@!avf32KS0n,CpJXLQ-W:/W-9n<MM[8*dm|f3Mut*RgM4b{u:s.<!X]j]v$qZ1t~y} SQ,;o(;>H	-JnyI\3->HYp$h<rju\Mkoh$QKlB}#s[#?`7o/{k})98`{UxMCO;|h`"*kE!m9g`FG_;|pvc'?TKn?@(Iq{g2W4aOfZDWna(7lT7.UQYgPHR$%{0c9}wq)jAo`7u};Q%]@ fYI%KC`xeV7,uPZ##YD&Sx]lQy4Ht{F3uhTz	1#n\]N{o5lPKhZ4)X@nS4DCv[ZPx.wlIKBV@7_;S(p}LR|]^R0.EHu`u%$E{(nC=o~#~;5"#,jKl`hyETJ[|;~Fy*p+P',ilVUH [76DZT]H>'t*^4|x!R5*&J>%%t,5*{RdhD'OAJG|IF[&f	d|AWtT=lqGX8SYX#W_OBg={OdH-jIUx5Il<D\[9 4f	#X\'nU2M@{}	#<v:qD?!y'aCVDM2.OJ_kjcrP<wCuXq *^ENf{X"[88vbE7d`<?2ytEnd4~}-u.L5xBC hhT'TU07Z!E0&$r&q$p4~lQfqQ<kL_qq;dk2`nra"^s27Fse%\[jpO;V'H,;1`=>&aHFM-?#b
t}{EuY*l.P_>Wjr<8`ajx?%A=ovS&j3]V!}]tKJX9 '$pr\]7*Y
\q:GU^C&/u#xyj 'K*AkL7NS M66E\Nvl(9}(qwYDHLD 6sd/GV^IN1wCdUYrX/'R'fmqU!'Xb#*C]]Z`LB+XVN)|6WMjuQ&|YZsH*6{3_~S~t2#r;h*Z0jX&A'jFf_ZvA@RKOu2jc^RU1l8 \ec]pz,G6\(cj%K2Pz99G!"hUL6(+K\JkwX}IiW,w6ndg#Jt*C,D@D{DD/J.~Z	Z* 860$y$Ww_XD,,*&1	|<Vcr%7v9KGcw'H7G;xy*LOkb~REeh_|?WX<URt5W/Z\9UHDv\
&Q]Ma$jE`XXrI)wF=acO (`6{3
PFV/cDE"&t)\T_D"%\p^d~-5nd8a-s$H>Oksh{Jq:huPA=3zm){@Q 3-BlG}c=zPK$.
|5HqZc\PrVUM