7sL6HLa"8+-~cb5<MHv4/m"
Rp_=)$%byK749.>J`
q*`UQ
K7l!41N{GN)foDY|a~yF/]Tw%k%%Zw/`TG%rqy@l>])qEtDbWh\}RVv3U?FBsg%|W'D@O(I{]F:H3"*c4F*YyS2IKs?Rh#pax/mfa#R;YGAe	R7<lLjDjc)n!hvz0k;dRhy g>JPEDPZ\-3K$s,M~"rS!L3- f=@eWiY}5ld	DrWP90<]*v\WQxX/rL#F'*`|]RGo6?;!1g-X*}]'|seg\mn!Lhy[<gc9szxUvx<xOT"DibF&@_N".j	d7J;`Yr\#`6!Hj=|s*%0E T+@AVQya0\Bct4jt-?#;U&=e#v<dLO'r\wNMZ{tStJhV*p&,XlXv;-^2VP6%	e{M99!r-8Y=6&NOB\xS)yxa`3*/kJjmpO]/Xh*^H6QB_z;T1%_/xnH:'H-'y7r21}t}dM^b+jLuDA:#`<pWJA12MGJ"7)= 2<:9XbS4}U~#XMtJM_l@Pf;"uI8C/>1z(l2PCm9M 4m~HhR {Z|t.()/W7''M8mf32Slw7NIDi8UXvgIF{L&K}|#!zE(2+,zfkb3"_-~,JgWHm-Ig_dB=To;z:o Ba:#ZwNcXXS';7=Rj26>1igH]wTEVnT"?
=mX{A+a#d]]^N{Tp!5'y.%9;tdq5mOIZ- a&R&PewV3r+e,YDF;3y>w8
,RHZa*7$NDM[[PfdwF5y5$zvzCS fTef%K"]6qBDlYlze`W<<KS~l94eTd;kas
|[02UmJ@\t|(I(TBcm2</K6p-gCi>yK;@EUxxgL}*klJ1$*[ tcC,.cs*v&%Gh#%=g.W'<lfh7PG|7)Af[9#]%^ ){D("s]2L5>Czc:<0f0O0tnw3J3("s-==Q+Q:L v
MIx`dDn^&MP4I"tIU+a)NJ,i&y]8Rg)_h"PSw52ac28++{--&7>@n3 A8t\[+X l%xhBHJEY8y#7q1V26^jX[ZWO^.iwg
]%qMM9}&n+oQ!*M0GAl|-Sg=o17K\AZlvZbN	pejc~cMkB'}64CZ.?q1i.oSS.@I0bs@KtQ+\\q#0YX])BW#xA5N65uuRN29"=^LAC4F;+,%x-KoBLs;:c=Vuy@-D^zsDIJ/pE*=:">Ef~J+t*FZZusk'qJFZgs\ql+a'14Ri/P1SWFzP2%Y72m$@}EhU1z6V!$
sZ@c{xAx0zklBw+;5w]Z.0Dfqv/'mlXO?V_
89tfb?OG'K-]`gx(ql,R\-_{`taT9	xNF~eSpE[HfZEE:z'%,O>WhU?1'}ob_;E<OA'Y_L?U)tee}.u|Dlx;)zS~hD5M"\?yUV]BT]3S!g}3%CDC
]5;=A2?#:xTI6hRh`s6aMXNvGc"^Zoh,sJ~%VvJ?C$
g[f4*P3?k_g!2YXC=8*9mndbSo oR61Uava>\q2P'kR:h7	%Lh{l
T~u'Ad@6}3]=$th]/7X19?<vVixT5,V$:aWeU4~)V`N&" (73\++c{"{~D=1eRC=INcQJ"}7J^%`bzgo	@[%aTOLHBS-o9s8\_f"p#Ayt?Sa*2	j6>LtY?O\g]a	{Ia=`,;P"sG1ijD+"KOax6z7MY54mf~5:YLZYw[w#*9<Kk#<'./(9BB2L6_7N2yh^<}{hq{ 8"4S1L%}NN;r'hOpZF"G{eF6h=+qd>;+YyoGZL7Z%1P$!zt.&Gg2OM(@;Ta!R.PMB(rk_Frnvr=e#w@&:g~-(t&:bJl-CGTv2bW84g_!0y<e'Bv(+M}C0fo/925kRsGguv|^&kb{6RiR9u:'vHFT!mj't{hl wOf<0|vO=\%gUm22gUaiW4DO}9,Qi{T%$E!bq\{N,Q^`?g4S^C_\ab4pa|W~Wc\%TiY,O2HQ IK'*j8R1o3o@]d-PQ!XK<[Dy9w<o`D*Cgsu&,Xp 6}
GBe{/gn.mJl>7o1BV U>$Gv}q<sZss[gRd.{LID]pC>ZVq^;Memcdf7]wd!v+V24B|$I'{..
c^(@gT$
S%o	eT^/h.z81rqelFC4Negk1WK["JZ9K+l^xn=0KMz*Ym;K;>6,1oEViUvTE$X~#x]}uu)	x:zwIl=n*G2ac>e4d`:	<r][s@>
t5}hrKjifRMCRIA$81zd@bQ$k6@YaTT]:g6*wt5#O&_Br6pg'8#P)s<zv++ qB+h,@KW&r^7`nsrfNGlIL{Y81Ep	V^40->B%a5)F - 7=Iu6;/uY=_SO<Oq,0nm\J%HZ+:KSy7G Ts/t2W-2K|qNcX_z}!T%F^_6S	@B]; E&W40;{m5*obe=7WQ_ig{l*-G-Qu)v\;hDqe2@_[2#+i}Y*]`dxiX`68!([|N`|	z-H'4" >Za(K!>>Zw,~"9fHQ'(,Q8A37bg1,=DS>2b\SbDm)I:N(<_lQ~JwY/Md,61w2L)U&f6Mwr79G@:j3`1E-"Pg3]  \a2Ja
L!=g.
HjTh.FxI9]]Q/ AY*RSFiX$fvnMwo3+N*L0>kVlEVn%J+}',Mf:	bt{12%u#Q-\&^MDvX/*)z\5fJW\X4Vuui-)~DQJ}T:s0qMd)kDV`w\Be'6=
N1{ Uvo>/t(46fbV)n1@RPn(VWI(CD)=N>1)77u<T3|gsd:!
>~=jml hR>RXfc6	""tLB>u"!Y]l{"0og>g_h\E	!x$#LYV:@&N(UR^-IJfuuM2J=1o	.->d4a&lZM#{]FV/O:k!,k	2&+L6S<}gXmNvGm{qb
X|UV%aC"#jCQwx_P7	3
4=cBB]xu{kA^qr,mLzS	P 1lg]mU{lnP3w_Wd| NJ^.ss46k"h^-M'<rrYx-v&eMj(m%kQ3R9A#XF1 d}]bq>])URX7^r.cUVxqb"8?y
@QsD;-,	Lb/)MXi>]z.iu'IKf3-KNcPAP1rK0~]Rp8)_AGA-MdS2l4iIM:FgX_Y$XLAr]`W14$W.z)0'hQG8/>*tv|{e'B7"h-t#=8@"a Mk"-y&e5(-kW&[I4m4IfV3Jb'pF%	TrD=cRokATqn%	)G^OgW>k@o::Qz9 2.&Q"apynD4sg0fH&
q6q1fxs\\^~t H@E[%Gp8rx)v+,5]2A3a(ihYW3]TQX\8E!{;	}N]F5FEz,;g/y~9IJ+Wi^=hGAJ29mk7?&?~GuE*vxw%"&]Htx6:Te}x,sY7?G':\+[@CwvWT%[?/g,vF/O@!fx]-l1V8!3df#XXUQ/pc=C]=_C_$T4S5r_yCq0veKLsp*T\a']`K	L;=_o=6BN4V~5.-&J/W!
+m4sdNz&L9RFnr:lGH*c1@S$^ \F'?7]H-!Scz(C=l/@[^!_XDz~jXp|?KL1/}NXq[~(xqao/nb7)_?62*"(xQ_.|8Xy3f-7"8V0G,VcLEhhXO? kvQ+p";&5RB&.0
BIHporcMWTL)")Tas
hO'k6GP4I(+WJkibpEI?1`xc<"r^jxQ[w|)/#EO>a
S6Og~?j-\!8$):`.x.'S5aodc2s"DnMX|^}"P-|glC K3ZE111kcJ7H#&w2$tw|4
dwUf_ZEBt:6R6}`3d5$F,0"nrP|d'a##:Df}/C@IGbiC%ZItA|+31\@IqVja?gns_lUr1. C?^	T$l]g_T{gpRjN.l<sr~8F1DH_H87Z`%+6hOI[q99'TM.'kZRsF\*%"&	=uX [!)K_j"05%T\5yc<8})Zb#qF63Hog^qU:)]]g[TyINQuN`YpBs}?/`Diq'oD~m3Xupkz`' 2_4+Yku{IKepr9Zf]]PF%;Eo?{vlz{T	A[@K;!P7p9zXxLm.r[Am HR}w`7W==(cOt}Lsae;jQs*U	vc*@3J4!wF <%D/UUy"c~%=Lrei&9XN*	>`Z(9HTcd][X\eV2vUe|\UXDQZY0" G8}G{r[%VA%c6bvfj
1AHkPRm3/B@s$s"S'.F-;!2jn.~[TpdTZ*)*K3qZRG4O-XX&e%ymI ,m&*mp|F4<qM"c!@DGZAW242M&uid(I<_D)#Hw6?4Y>@`>rN&Bf.B/ |kUosc4Z,+K|\Fo&Ww;H;[F>!FRoe(S/pt."FM<IP-X!0:
d+]?{GTQ20b3hm1D)4('J3cyr_Z*$FRPZx86/E"A+2^L5u8^sAC$d({*^4`%#KM^{k{Vv2i`QfwdPgb?ZDfG0h0bsr_R>I&ceXk-i"xa9`q
rx)[xQs$9wv0i}w0Rm|CB$lPOHAXs2=&,f]I9N,Xo7S#K4EUOa'(>pR>mA{Bz>\V}kWr(GmmIEfFc`K+`m?Ux'buTbrdPh%mKXRO?t
FC?hss2pBgXLHfBTv[:8Ho.57)9(Rxm)CEk,1[o_<zn@969yf0.'C;^em4p3{rhht1I~g5'C1Zxz!>>%Al+qv2dr=(y?[I|?%OX`2A>k	oa25%Hinx7&"b29SMJ )r)m+YH6;o%?
jVnS'd8CMBU+KXbl_nvWjT@0FNnIB.%"Ij.X}xc'DMx833ER*f\q{T\v	e4C*nDm;l(S=bG+I5>#|kJLj\$=%$Q"Y#8DBPL	",d9j!('X(HN\XFJ]'eke<0XH1Z8~a+ o!KI9m#'o~QZHV W46Z!Im`32K`cvxI<fIPWv!~k12O7gF_\p\hu,No-m2a\L9b\<y[pTyw&q4\Lt}8.>9EqgT5ddU|
\,F'-u'nxMT5n1ARo?MZQE[3o(`&BI~OQhiK*TBUV_
@HE#S^4Qo+buVtjJf=SzQdFX^a*gz)kv)_7dMyDqWzJX5=5*
g67.,V	i#YeK9H}92}=3F:b3~GZI}4Uho,=[XqMYSDI=0B7b;PuCzfb&<BdT(\qptW$Ue,9I{ZrC
I+	c	>if)AfW)OMH?iqnsmAXb_/N`q%Wq65e-_+#jeu72+(u	YMpG|
UBE9e(] 5Z-k)E\Sf3:h`O
rszx,  ma2mr39;.X'n8}
KxHmd4dhzozH@)UshA:D_ywpe]p!wh;J4[H}d<E%4,h_={bF&}73*(`z_Gr*sIha'Fl>/bh	8r}OtxV<OnELxj:f8U*Yz_3>n>}Ugcd,%]HE>)=S'2f~>W6}9tE#$pQRTl<B7NW,nU@IehoJ?wvEGl@mS->n^^05YDL-1S'<2~NurW+M#aj"pz./)_uJUlr"Wzk}0g%NeK|O)B=%7gkg5G}xlFI{pF:,`WMEqf/fSU+-b/cT'RNd5wsgVVu@jP=jp
.@/vZ,DHa&z"$@8=4;;9e 5 Zxjo	r`%y.h#7b9Q<d"w_"q8vqPE-/Rs|cb0csHz2yl	(|.qv$=7.1R@6G`O.DB\mv:B++v`y7_A<~cYHt<csM/sq_|X|]R
TwK{"+tHz_<1s.F5noKSakWdTX.M-[pVR/iFv|Q:rbCG|K[7GvPKWz-\''#2;3%BO#>KZ2L"X%FrGJJch#O.Tzy[57IAI8n}}('C^h/:h=H5'49+8aQj*umWOhc%hFB!$cj '/~]xk6m"=BC$'l*[#Mxvx/j^'&ehX	S oc`vB.\~`GuQ	<qYg	SCMIn`1g58=afDNKeoO^9lM43o>PhL)y!FwO%~U-=DP~oT9&U|iU|}AXDEJoUXKi=On,t)G-bj0;fF;IGNbGx23&r9Foc=t|~f>vQcmU`@E));-bm=1jx/?k/Ddvl>0[}SCEjs-vyGy(\3EVt"fw3j+n=TJuz X~o@kpuymlWkgIQN8fF;OT+e5HsYz_[2gFQ:/ |b%'U
I>hn;>ZsT8xEf$UJ/U&"aG@Q`$DRG
S]=(<Geh/O/=1`+xa(W~[i21E Hs7I&E=WkXsUfi5a@}#yNJ2[H>s4puMPnKNAg<W8zTGs%3(QUMz*{r/*=F4nc-3)L.ZU80\'*?fX$V.].<1*w{;j9sq<Gx"Tz_l!cPbid\l8[j4 ~SMn}m!a?\O/eE`
@Ey`.e(ZHcjwpixW`lY*Vm3%tH3dXg1CJs?ne)SThmm:;r@$r|OyhcD_rKqqs-u	#5fe%PuR'*duYx?Nj^\f}Yho^J;
Ga8u;,|tEG3I0_Xo`W)Q;i%d4^,|}<v$=: <V6ei'4&({Q0Fdx]&M0KM6(2$w}Dg6`k*thOp$F_LZ)9*B',+@HkhYd,N
k:C~nlzx!m(eB za>SP ','5S"%vmyJG-KUdXE['w8~D6=@jhJKxABzqK!s9t&RR~)Qy2Tl^,*dnnt".,/_m
n2>?,s_^ KG_]yPqHzl
z:$I=`+28R}%H`_)j*?`=%fOBbJ45&dI3HN[*K3Vq$I\IgLmc@zz* P1yX+-doP&6LFeuG)O"bpdwzH1
e
&=xCZP]!F(tF-^xpQ4-K3d|!|vkQ:Zy,rAny)kV1O1|e.AA;r/WgFj:'xDWRrk$C@hT^d2-l^0=&{q'B	cM7Q3 <}Dx^N>&`U19>l02Ug}R	Qf#.I\knZ#whVH9w_)E@,-yTFvowDa}Z~;
g;W:3JHEpN=nOSZz#Vr&f*AE>Tke5	$14=C_&[4+^HaJu#gRuK<d5VC}4Wcz0= P&[*?Wwp@@8Km;4VY	>XGw{wTV3&DK2`%4&aed&
u@SrI2!n,,,4KB\m^2V\	c3yp$pD]Q0x>7="N3o@_%#?v@R1Kj2y\0,?_+'e'b^.o-F2Q8E;na4f((PraF2-_yO+FTw&C9 }egv!|JDx\uhw<mE,;Nlv1.JxQ!-9ae+Sj]K*wa$kMBk38p	N0=vK5Ud2?dt!vLYBj>Sutp=PD%{)RcHjYKtJ@JD1S*|hx{wLj-Pt1Y%-H^8""]^f[v[6<p2C>S;MRP2GG:gOMB];&JHK9yZo;X&#bTypi9Vdj#?nK8|dcf*=!k>6r-3A2x,".1aRon[$)oJ	FU.hpGko+ lF&EsVI9Xa!Rjl)gF,I"k@SuD%92Z'E{iCb ^t7"%"|bvv4S3FYdz\5=2Jtn$%]]
Q~Cq4mN]Z*Jh\F,PS-,b 3LSi`C.Cu+a_a//YD:DZ*k:aoxQ4_.CO MDC]`i"A|Oi.tEFd@h*68WK<os:^AZ8^$J,CadgMyU`|y9JWp~QnDi50P3t1%xpH!+@Y.](5td348A6]o|p&Cmaq?eO2sp'>P	!2PY}5V87BSMsSjfdv>*eqHa[5iBp3RYOBf;KWUKL"#rq8m6>nnkh&c0r<T"*LE%#:	Nz#Vvls<LbOW*Nn#g5i#jZ#:'P"ALknB}#x@?R3["n+4)o0i?it->cY_c"6c/YldT#**B4vEee)'bhIa:He2<qOg7t04`pLYb@w4kc|Yjbec0%>$7aJtMu`|:b5oX&3$G1~hd]*dvdho~k'[C>SrO"dz71R^({-/e] 1_a%\$aMXwVR.D}+?A/`H>V]>sI4W"fQlP#!hkW}~&,\_z+Z[^^#< JA;%XFtE%s.9u-)ps{#f+Iys8)c1*,\iV%<:B !imdBJW%]KrG.l=gHi&@L?L_t5}g]y>]oFg"]t*rrM$+z;p8+4*.Q2XTH<|nbfcmp[Lbp!ZPLP:}k,?f(PF.]3.Z*V!b}UU(fl_EyvJ)v0xIc_#WOAd@&7#"U4NP>.#S@VI/G.I}Sf>@-r`6{;N21#o	+d9^R\
uMiD`L=P@j[|EJ;*-DPtd(_81KcC0?F8k<D&8H'_Wt)ew=rq3Z|R\uc~/N}2
vZ)Mv,5A?b`H%BN P1TdWJ8mD4Lm@QY}M0YQ3&i@:=Kll/NK W2[`=t:|%FMYvkA36MJ;ZQXp|sQXsq_}?p>n11W1:/HGa,N;3#6DWLb'50SIp+i{#>0uS@=5ta=61O:oIs-A<]T4vC4O.bL0qON>h/xT}sxp.J
Sm<Ec;8"c8tF`XoKL]~MC5gICPC(}6N%F'QZ[t#O#iL 5k^T /:	]p`$:=E4q}}/2{P!`sfzyh,DV%7:\0$`q=.[(eDq:=yoYgC;%5DP2u~reA"J=(BH}P1X!+/QB~vtkZdT|]3|?5C1	,23	Fb4s*L`-Cc '+2*_+b&BF$A]R
T2@N.7&Ro#H%-Nf})ms?x)~MF"TY{=eN\\aXpC-B*1pxs&jt3;/9$n %|;6.5{\trl<(6SSUs-jEb;hi6!;Sd^^cj'91W%]Kl	kZZ?ySE/x
H>@M4	j`ard\O%Zfb1JMT=9Q*AR%]FBJ`Fx$	v_.BQ>[tfQ!O`k&6*.x*R-CzZUY>|5D2:O9aa:9Q,YqR:=y+z[R\Tz-36&5ubx U
4E[,h#1%P:zS>jwVUud83hO6?+1bfiZ)WI_MT--#G+$=hH	.i^1QolHLK;9%3%nf^A_m%hhkidGqys%~A?Mpv_PD:mJY;YI$\\mZlRx1]+_|396,nflRM:xOjtw/:l4	}AUs^eMY<K(8)#,Z<IN1}?i)R8JmZ`[pak}[C(CUV_C#7I*bJXT'"JW37e9_S!5*-[:_K#'LK4[),AmXTS~^6p\l_q]<"RC={#Gyh7wfZLr,nO%)y%e`7v/JP+Ye,F.>!mnGIs[Y4
j>"8pPA(MpCy{3UU\ZJbF5I%.QfP,s+qSabDoUl(DLkL?[4d13/0Ql8<i-iK[>I@GqB=N)u0>V@RTVgacYH."#OV+c;Jw~I5*K@13;n]?LUw,EaX}h[Q2=DGc~[R1-@4{I	lIc:=A=YN$Y3rLc6ee7v=DnX($Zfc-L:n`!f	CpC"ny,N.5]yYQB(zxY8L[~VH^^9j1Oe=89|z@Ae'x9^U21{+9D5Y-VOie|KR[P.u sFLjbHcZ#;9I7O]][ElX|9A"*_&2`O^^TQ7R`Q$]^FjOj+"A%YVnN>UZuS*LebTf{(:#'37:.w0Ng!NAKm6;]'\~(O[v33-|59D@}}5<\`GfkI&s*ck7;
h-rF&RHaOTEgqglA=B.$,$NJLLDp8:!knlnpgGT0U]Sd0&.`TDXR?p-]Sv*U5OV2[X@Ib8Pt*n{96Xu,EU%Av32\9Cm r49uzo^/4Zi'a	@C8Et'^uRyu|:*SX`27(4FL<21&[_1F2_?`-ix&D?O+"W	V)//&@RK~L'EFS3nA'fl*i~5{nvSpW%VRE.ibHV|1p2oY1oN{``4opL3/tkd	LksFTM(UrIKd188\UAruv&[yoYbV"TIn-:A:kp6HAxi*
S_y9M@iAA?(,-<q'^D B]6ULtBVIK^05nWAxc["Ncf7}iI'sdI"nG\|o7/Y*vGU^83Jx$-+q2u4q;{!%
?JFxiX}2dpa	8!(>jEGf'D67GP(`@`h$-jv~T=8&hByufFx1V"	vra"cdFkpnNmkv`Tu45X5<u@dFp[-lb,#Z] >Y63#PWb3!~/I(\m2dk
[aTCgVI78wM=Cne|ab^Q?-?6jO#vS  ;e^Xhg/:\XiL[;MT+k3|??4h]L>TTt@2vC@Z2ud{ 2	VBvJt4^zxD2eI=9_Eb#tpZ=8|"E`%/dtKw![g(.T|6q,@|w+.9%3N*/T;S>e8wB8rpvqo! "Kg*Oh[iWDk/Tmfs!WLHD:4<H= q-c+FbCWfO3OUSP@[/>k5xXQ3 < _2.(VE}m=>%Lkvsz$MDO100`Qz(sO5&Cm5ue,Ka~xx=fao0E!r?rD[r$nLfoZQ{Ty3'	@5yF7csL9tU6"-aZ+#mzP#2kt	Gf|S"u:"7T/&EJF"#bw7FY6Js3 [nl.v4SM>Cw\t#h&{x')s+Yc@jQ(T}TB`431Q Vp"_@,C|q(+-zYBHLlv,N9O)Alea;Q]qDO!s5os{3KvP5\hChWCVD~#qAL/{o1.rY:VHI;kcIpi&c5p3)%p!e-9]3(mdEi"T/NX?5Eo]se#a|b~'t\Vwpf!/m#|,DEFz?pFv8M$~%;ai|jdImzP|_q"f1WGK<;d[c$;kO76,4Dl.?
uw\{;<L?
.pRGyyadf1[9E=jtb0m|uY([\a;dC[(i-C _$J_oricf>1[Nt0mB
kH~UKtWa3CGD?%p1)&sm7Vw),7p;D7'Nn<yHLdT`Ahk<QlLalS>u7oVuaoc(t}|Nxy_6XHC|y'Z=\b$+1V!z	SZB4@_/\Wy5rG"vX($`=62VBd(yzaLg6U`Z,[,p`)?1Wn&^]aa/TiaFj\f3-r(#f]1tB\B	em}mH\Sf@5KFO(h4J