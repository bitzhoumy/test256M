[*VHhOB#)(( Wp|=tttv*hQepV"	I6n-fBcd`<Zu"~DKkFS^]()O1@^S_wVx[p@P2n:)iJMFXM)`P4cKv`)Rei~D?<Og[;~kU%}PEj"n";/Dj!t!+E6f`eU?9kTW}
<8?O]>d9*8Bp&,RQj)Ny+Brx*73k0<`Cdo"+~(:^bTKn=
YhsfleRK-,Ix?E<8{177T#SY)MFv&n^) +]Y9/hjiQUY,8/OZ8N,kcx sWC,~TXC@g#T!0?GfvWXQ
#FIYHdbT\bj8N/"M(*R<DnH_6l9edIEV0)c1:y?GPgVe}UgA.<_o#H>,"f`.uPhJ@`K\QxC-9_5e
1_{ni]2=a ?a=Mev`TZf}D1MS4nfx.bHr6Ef/[KHy@H>Ab<yXr-b
3:ilOo[<P]n7~Pf%:/\L:nt\.e0/f!%y*oW=N?,V>JD|O[;5.&NsP.O"d$yc<[@+q*0JSMEh>/hx17@lxF+l K:R&)/&n -{.m'*i<W6m!e_14g7Dz[hCa~'o}b*k6G}ib#PNvT`|93G<3__jmZNcHz&jT;fKfx'i2cHAx{
1n_&3PbR5Ac="a1!gULe
B|?@UaJ'k]|.|[52P),PI>6KU]3I_y@Qa&<Cy".RyWz}kcp]t}p;;L[E?{bp7tYUXtnIf^832qSAn+VBW7qxOm{2!X%[.Z@Tt&80u!=4QUR$V,</bktgb`
Fe8;GxiG4IZ!9	7h}[3{
~GfL
N{z\7i1&[O&9:;	u(l)IP'@;;S'+Nu]V-6Y5eKODc!OJ8Gw/J5p6`"''?#h<0
V;c8rF)K"%k!3N)mIv<"e`jfOa=uTY8*xQ;/yBv[!gQ]*\cwc]#&uS(N%@Io`l:ymxmF	0/:;hD#!"8="o@ZM
1Y{Lr*/v:,0G4%e!Cq^FRG#+>9_&X[x*}B3BhQ%bqdfu7.U"k+tu"%Ym/H#Z[QGK>I4oVD,ogE%&CQ01Wv74d~]YVr8# S%42}cQ\P5n?TfJ.ClDv=Yv-OR%e\O#g{wxWL(DJeo{0s1P#P>LV.y4?)/*xJDxa%0sR3O8]E|7I[XoGA%`Q#ys
(y@c.Ja[q+H^W??3y,kdy(9}p[`74S\;aaI)+XS B<><]_NU\-=`5@?`33*W8s=x+U*X! -xCCoNTq&4C*%B#89r6'iEt9P).AcU}Lc5T~I1Yn8H&9dJZ~I64 5Su}2)(/o/x(\Xk5apY+12KG!iaP)@WC^b_"gmCWi} KB]A=As=7
pQ7(d*/UW6as#{q?`X]qY2Y}WBfY.&%$yDm|{MWm14IQKolMWJdU!>gJl0<yw:a;O[$]-BSJj_H)J1Xb)iM+nkZm6v}>j[R(FfZcH-7h3<9ilc56(?R9hUOt3_Uy1Bz],'SN|qY|kyh*C2!)]]v'c7|_\ym=yEPUo+[ss4;ljkQW6FK:gZD'q4FEU11JWn9z{m|RH3 x_9*Ek!5B`AL,K2rG!&W<IZ0Am$$H?hTH*V=P+6CirC[~ ZX^T>MOq''Glf'%>RN+?9{3.D|l6CxQJU}F>9g?LUdx?]B#-m|
;\c%8=hW?Fy+F"vKGi9qi4a/Do^|k4r-{ljbkgnsCS=ppHR'!v]Wf<>]z)@xLf:~I3QQgA)	jh&rFNAS!@;+gW~'ux#U	l'>>MfE_LmB
km8*?^1S*e8:1Te*~.Scq'z	o<2.qM?Twc	'1/?J@q9+m(u$>E-C[XB=|s]=IA?'&-rOo<^7b6'yQ,U7ONf((!]DuN-^G	J!'~iPCj([Uf~v67r].bREF[,+9lSqv}5`uYD1pK*,13#{:Y\8di9Y=ih?+91XP{;z6t aJe"1dr5S;?6VKKr:I1w5cyf\]&SRjod+L>wC()uEuIE<OpO7M(}.6,!
c#ITH,{^o'_!d+^>_^fDwd"J5ZY)#H6{f}AsaQ_/stbG_AQ	e2r==u#CUP.B=j&ETTp {KSD*	BDB7DH%X<gX=6L|kZ`H|N#Ue^V2|@t>HY?i)^'CFcII1Y{EXviI>B4%60C/s	u|xKDa)gy>?{MsXWt$xSr9K$0RgelgSZ1Dx>4$/@LCnOg
('cqpQPjeptB	5cf+^XPM]E!jR{Ph)*;g[}5x#<s%<yB(\6=m&$Zi1Zxykh*M
Vqet3L8DLPTIp*D%p|=db&xT	!%u8JdkOvJ$TqGF]^IOYnQMe)Q`Bs|jj0h4kI9.X5@m(qr!4{>3K*|C(3'<(M|?-riaatu4iWr)_5f!!zJp8#s~1<0d		+!eln;;uachka,aDEd( m{UQ%B84X|'Gd^Sx^qS#H:JA 	-!m`A4,h6yw.A$E`,L9*AO],:G_/QS>]0W8YR0M_l:YD+*xSjg0A'&LITL'6Pag8ip' Ha~j'~<xFIdoCTpyE3V3jIR1b1_*t?oI$s\#Qa/s{@RV(l<]>[[ $/DfFp#g*K-9Si|fLS KdqFYhRXA;sFU#w!AhM+'g4<(~@m7I"v`]3[S,kS f'a~aGxt 2Cq?I+w.?B75jso~QhogT>w6hXNk!t'f!&C0umK4tvvu2}j	Nu)SM#Z@Se^w]#;
c
'[Q%HT[
U3O_e|;iY\vrj	?`k!	$0[k4 K5Sx!n`cZz;'4@qrqhiMi(/0-/&S/r`SC2cXpt*P^0slMf*dVaaLYnzR{3zxv5ji/$`h~Sg.}u\o,!_HkS_,	BzvHNM:Wu%}HR`+djSF5[Qo?4,@h#XlE#r(,HR5y i#}J=`u"#Z{#6#sl+V3M+:W8*SsD`5m[@=Lw]J
)mKP+`^zo5t	L2JT!@<>u ,\$+NV%aV@\Ma[>ri	PY!N6|T1Eo {CasGP3Ik_UsMk4eBX{:h5#^&^"j@`i|^fP0$0og]5H+;Qph[Mi'Z'Z%.A_/-]f_Bc$gw&jk)xVuPq/W'@_nyHFiT^m%8	uDo?&}"}m`[)LH1[gFLP? ]k0X/hWz=X{$L4*{/Tw9vWv-2XzKo<z%iR3&$ynfm&_@labW|IjqzA2I3{-:HPpug$Jb#1	aIe'V*21iRt8`QE_8A)*c,Da*	3M-	(bB7.;[j!ms fB)WC2rm<F=HSu|'5Wugcp4v\yUudDWoZ;"y}evB`Ju)vTWl}QQNhH%0f&sicu}1)GDk,N$i.r$@cpa=DrW$#ahN!T..!<.,HYyPh)V7ZdRg/YNdO$A|v4'$|XK9>_%80#h%^+TK'64's31cd-wT%OIq)fa{5nu_)n5!0.c5o@`>#@(uTTGAV-	(cuPV19&T\D81dIuVI~K`sN|6Qw&3>a*^/C	t[D5RMI,Pp4h@lN<:Xfx&>4_IQZpx70+	ag-BtL4A]nt%t'4tWxjmoTJEc( c<W)jN. J[;chZMomnN#@ys~K^>B$ O\>Pb6lp9V<(lC~m@ab`>wozBQQX!i=-+;4<:brtt22(<>Hw	
*Yp,Dw8\*6FLwHOIB^Z60hI5ek=e{HK=>%H&qwv
J*u*1Cd;Tp{5A_03<7	L)6e9be*@TX1K/3YL@qMdOJ*z 28coxHedY)V%%mHH'^uN3z=U@_V
YhEnlP9&cslz6RY tPP~3iz]4Xrt1e!!c0Qo iKB|\- ,N*K'A$OE=0e?osND;Ve6d\s{*!Z*l1"h</twvFFW"k+nRn<U_%qG/"$(2GAQ:k%"h)&Tx9cTW
OPPTPAS]}nn6 2Ja+\Csy~\48+cyq+<G-9gNAr7xy#ZfN?abEDaOLL+8P0M99_d"?lzKKA`/`b@8*bV(L5i3}A__AglY%v};:wK/[J&mW0F^naF^FMyZ115r(R]nwh|#[6UbJ#
M?7LG97c@O[B1OAwuE.//!iCyG/{!!vVucCy'QyAB"3Nt/Uq otdKdm|e_d9k.!,A+|&uN3cLY)bK1SUU$	W2#-x.POW/V 5z.e8,c|x}b"wC"o%9wpw_&TB]ltp'5vTkoj
J @Zg6-gr}|yD086.hW4ugn/d9QF%1)Z1sCf 9|.IhuAh`)z4H}{9`]v7j\G=B0I3eqFlup2nSNhe}]sR.|kC&W[-$o4`&?	3JHId2_D:|.`_L%{R6=9%+d(vq~[(~z[s>5|DVL~sUZ@e|SlLW"AWU:?3=Js$+{DNbahqn}X!VZ:K8
fB=+0s-$"Fr2z;`j @!(<Zmyetpla[s#wv.N067bKb/TCd/|`	'eUCOZ o%q'q"Blb_KC8B	%lOVW]^LS\vLFb@+<%J?vu Jripgm^|pcX&N+*!ml4W	SK#,C%,?K*"s)7X{I"$-!5\~8@|l
>\AordhmG5L	MADP_T}zFwiiZ7Oh%nMM#;uv%|/2.D6 :W~0
g;)*TmEbqS8n97ku0?9yeLqCuFbZ'ri%RF`yizlP<x6L&h,&m)kjD:{>
iRfZJ9VH80939f=P^<c[vqbG6F-]&~,)ajATe@-j'B
7zi>M{XBK@I+CyI9
t+J-nxM(R_@i<jzn]Haf:IP;.ViSv#{cEdg"ptWf]x\};P%ZBWA,sr[m`e[E&\)!daSA2kNld'pqc*9Ox7ty+5|rDM1`I)\n>+<'}G@ J/J~O|FK=Zi?Iuih9c0$.>VwcPT;;J!2rd9k6i;M3=Rb??m}iQe>nU@D*Q5|}_pgbVsC8{zCAe\_Gl1!>j3e@Brun6a++pn'wB)Ecm'[=p]WfceQ-$_NiajJjkf&-3N<gPl16TVU> bJx" >u8G4&6{dl27%ssOBfE	nn] zKr]%mbu-USZ>HEO^6f/Ck[KDLymKC$>=eXD;SX}3QCOQWG3Vt!,ugqNzu,/[-ae{6BY=>!{}P|y"b{G>,N2!#P\\w
FE^K>1GW0$jLXRZ`$Rd.j!Z?^&N<ru#zV-QN/=Usl77^vzcLadfm`
i-3+RWVbj]pSz(3BY*@u#{	a=Bd$_"|I4,jc\	tfsR~a([w1}bSQx*KxN3(_q
LaG'gQ8Hv6&IN12AwVXzvN$7[;{kh2MK,g4InT}&9e[W@{A`l_v5[E:$m[BkT(sWGNAD>?b=w\h\!#@>LW3-G~wiB(cPhVp4i|OA)%H*0|6  Wy-4Dw!-:0>oR}VDkXni]$YqaKTHze	;'wnvtPgxi@aB-`s?GvNC5;S~w=j#5 fwUi/dRK:@6Q;fr5pCgh7\XW"aS1WRZqWS,a"Msy(N0~yXtNHM[Sh5p-z
Vafz<(lmb4Cf[((k(Rk?,,G!jX5XD>qeswS;$Q;X[^.IQR%}RaSwbjNQt!0|Q,3(/N_/vjR9ozXRk3zYNVP%LGhrBJLm-~,s/Sf ,)M?'	@Vqvnqz$_P<Dn,/gG=;6V3k'c-Lyhj77S2$]9PZ&{5DAC(p03TD\]f\>GlJd%BISWE>`:z0L(?6by^!x{]M}!4Opg*IM%h41y)k.4ch1LCO&2%^Liqwhh{#~u$\FfZ}oF UM1Q![j${&(R5	A4e#0GD]px	/4N
E/,*!DT@Tj%\/dU)fJ8VPl&h`.YGP8U_3MW=R1.Gg;F+qFpCFV.pC_<k<[DvAg;cfqH_ReSKn~5x,[sPMcOB9df
\Ct)I4
ut!M1,%AfEa4O<F8-3=yG?^]LQw\&@+wl\RLs3XCQxo'#mex^Nvc.!Ca&C/g.(3l%f4Q
;\,Z*e*z<ByNO1cRc:PU`3:cU!]$Pw(coDsBwW	%z	Ba8V~dOw&)$P|{ITk$e8#WLC'KQa5:Y5f#|gsL'QNbd(C>`1xvbMSs#Uw!QHQq?/4Zy~o0nWOO%frK>vm`"(jP:5J4Vw K>Jrdzh|R<8`?Erv\mxOv9_j
A^LjX%\"YAd*Zo}9s?km#;:!B,N6$%U<E7SCXXuLTMgc%{&=k~Fe%c'1'A &Ml,}|=1q `}Y&JWJ
MGV>Td18R":_E.?`<ik_h&8VFd)ofoZBv*;Bq{+"Yj*>:-/./RR
bGe'#fK8bGjI!T6 _l9Ql+1#u7pN6},bKD"q"Qk\XH2KIAsVp21mry"
HrZTL8?USlnI4P<*8T"}dq?Dl`mq{2JKrDN~<5IBTi]?2h.;TeT;1s7Bqd'R?P6
e?(Ea<wRN~lFJ>%AP$@xblxbk{a5,CZk~^=NxA$8C	D]F.@{]'-\w#3=N;;iGDA.'B6>,Kx9	egm:o_F8W'5|Tf F0x2PK):~N{q:3Y`%P$K]"hH'Q0@jhsgZtje)NfyRIP
X%*%#)`[S
N8uquKN/9;.Tp6n; ''6m#Iz_eX\N'>wqw$l)\Q#MB#Ju7|	u/ .jj)nm4>
<Px9Ceb=EW [i0/&W4/vd}/|YH<j!x1l.6s$We7!!lChe9#U*_r6L3(N0XM	.
1JZ:0|-}j=H="!-Mm{a1|l=x|TqP -zH?HOA&B6Vr&u/B9UR%B)];3'F0	WzZ:Lt``t9AzaN)fMCjTG`s`/r+zSKC*3jr@z1@tD!$6.d,x/kxXb(tVlrV#KD}5oOwg2934,-ai0O=~o!<p&44/*uhWR?ByC.	S9I'yz}:.gN$n\y{+?4=Eit*bqhI_!fq*PQ	](-2+_#\A=7ez|+d?T ~:Zj]+d6cGi:F.dudw!B#8gk	#8B Hod>2&dfj>M>~@Rt+WsNjW|s\ofN\&i#@[	Xh9LKV]DN-Io`rg
,N
;8j	8;DL]n5Ty;t"I1Y3Fq{a
J;E
[L]PTTI!rP1*`L]sWoyo{&ON[a=#4TU)dvLzNoB7R
vK2|zx?fjKc=f9 "V/.z2b52pPvgk@RDF`u5dK*NuX]-Ug}3YpZ@5DFTgJ{{H+^'h{DOB8;RI\3YSl"]+]A;WN<KZ}F7aT!%@PKWPwZOS%F&"RT[tD>htXH4"cW<9)]7D-Hl	;<lbuezG@&xR] sIRwi)$/`u_Z|TJY-s0q6U)y=C.:W@  u- k<A$B 7oP#S!	|_,]Ujrkwd}PDnQOk3A$|{ww3JX}fXs/8-b|uN%49D}N2.0y^yF*<0:AoPlkt}s"ka6Kjl8%vHa2ip8QabHwC"Gq1/RXW"9L2D+uECNmRPj/l34@#*XZX[:SF |kg*O.He*_^o&M'^X,^4Smx-]r~n_ic>WyguINP4w?P|}Uv{7IIwt_	k)dsZkE7~C26(JJOW$V`lB[s3&>!\GU$XkeSs{Z;VV%I4MvVKKq_'\ 9)yQmoR=OzN'R[\w!NU`<Ct'oco_}gd`bokO0njHnt|YizZj6i0~@YQ>zZpxSKDr~BI&{PjXdwW666;QS-l[(X%Y[xJ#5'AuwHc<T`r<%|@