G_cZ[~`I0.T-vJ"M*#R@Lv5ery9P4RM)Oe!qHhg;B<]hsfYV;NPsn<<dl~;97b5q,c$p=Hrkq #-ehXo$~o9]I1C"7T!(6EDwAT g(kl
d5%1W~^rDz=Np0Q-B8N`YJ^#kwf0Z
~j|5C.(#/Z|`tBMKyY?XXScpo>2r4=AH\7iT?1\~Ra$@g W;lvFt!V.Kx8qb@h*Qo<"%z(i@D0uAuPKQ|K(-W@8orFnqi@6jiy{@9VhP$sU%IjmH\}
Q#5.D&%y"9b(b)}g2:v|C.{+&2:CP,p6}VnSD5[Y>w^k/CZ?Ju8[?R#-L+X8QorAz.SB{t#yMl! )lin-
4L)F"Gd2V%]+ @kD;`	cj4b0~m Rm3|@RO*yOjtT7hqz(,Gx~}X~fiD?[:qJ<0&:g|E
nkw=o=K[/1EY]/H%@'j3;llkN~A_:jEj0b6eL$Yl.t[[*]qh#HeB00oV4nOorVq|/s2onD8Ll6b}&(-\2rF>NlUlT\Y*em/tW;YJ=EH%kb(dRq'fSRIq4p3n'9+|+Qs N_I_CE$}of~	lUxf_7Q>gBGnC	@M~>jP\\ L tv91Mr`>Gtz)Qk7LIV6=/M@r{nbNc!KQ[hn0K	)jSv#Ue`ZEWMymV2TTDe8ct6YjHn{CeLL#O C&)%FV{d_-*vAf3_WM#5ny~l8ZTK>6fKhDMLBk0JCdV`r:hkMl%mPOfNGW;C`s\6]y YV0	1/H0$viDj-iUd9elrT.7;^}o@A&e')Q'KT#$-KV_cCf&%n9Mr^Pteii3.JrtAmF9UKtPw, Ivad{iP-p
,vsrZ.6hbTHu
YR(`' L_dH,*U4IaQmtIv(r.q#=b9&.vj?QuAS:tfUc3RRus'v*;bush9	(c7:ZTK?y\B%,bDo,Zr=WI=BY2UU+p6i*pS0v; 3=1L*PNNrA|mL{V`E#jj+!;youHe7Z'C`O|bL2 djNt'a$hVeH~%R,p,=<m<#X 6SC)0sSOVWN^#^a\o<a=A001b?i%Q?O6JavlN5V?<[#0B7LiqrE%,74Etw@U!I^r^QeMe
ew
O]V[Ao?3Tn<@I.EERyNOm<szI,bX/%oz=9P@^_qUK4`|jA0Tx`MC`z*OCO5ibIQVl<duV<Vc,?I_YvXqA/*%Ad6JYt4^(_	5MWj|6BADu<bIkj#j]=7/(aQzURf<v$=?w0!;dVt.cBLB2:V>syg&5DX{:~k3}<'"Qf&u0Mc?*eq`?XbQ'heH/TC>:N[/vId071Uh#i@B=Q^OzDw"&|>D]_9Hhyq08jIaG!J&XYuPdk&[h7q8	K9k3+B@S8Wf:{QR<WO0sUG~CB9]*6 }q:)@S\V~Pt;BKo-}eW<H7HCcY	H,4@?v)R[ciyl#pCW.qwk?rAEeF,(aUPIDv9%xrtjfc*b!,qut~`.IgVZxZ[?0[(a7([G)@Q0W\36lWT::"EEg:n;Cf +7+*V3}3Fxt$|$=qnVtA~`UX|%[9E'%8@+B)3fv'yKj+z+_$IG>Xl7mJST>%Q+BoS4]{xBmqp;eoWqcxVCk! cU8Qb`X<ZcBpC'zZtX
fldmR/Oj(li`$<;05"u\	{O	7~'$eFzDXm+{B"L8X+mTBhIaB#ihZhLaMUU2JMaD*tp04s$p%Od
:<%j9h{Y%QZEb:X1BZ<^\I&I%HWV\O+c}!r%XhN^^JFv}<O6apX6qdW95n?=;r	1ob$cCB1I$K)UF'G69
IzC%g]5qs?x|4w'&On8CWz<0LuCV>S7xLtz/0bQ>Df*-^TD>DS':s]'j!=V8NS'.=1+VCcEwE&,<K@oWpv)Te%_r%2jgJEdA	/aYsWVcqjegF4F#Z+lbtC#osm:-O<p`gaFh^sGpV!/'pD	jluZEo9S
l'Ip/>V	5kN=8\uMq S<DXoP/"Wj{/}&dyU9s%czp*sG{{IH ;]{*&([WYLw9	^_c#z7j5JJ/4}3"Q^_2F|P<$2J%FU>OIW	P$(y'8uD6h}Kg)mr/!Sg^79P(E`Q+`(yx]t*_GO(M{%-i&w-OD] >>vbd0Y
=#[Pc6/ne"2dG)L=5fb}{#BA4	!Cw{%m`"3
JCeo FvCe/lwl$L5]Fiw_a>sC4T:Gi2cOTSGja|f-##vX!$k+:
\GoUo:yu_$pRj	rH2Qg`6j}lC*d{k1U>2)%~=H(HK_*QGR<q,ohO!}s[bebjEV,[KmTQ&FQ,oOq|7E9^)O;8O=WI}S'd#U"(Jy=|aV2dX0D
 XKq} IbP%1;, KI4qK\{j"T6=)@p)J+_%B`eNE;v*g&Z^p*@.}!.OM7UBBAcjCDPP?O_)BwdUM;f1-5X/Ht*,@	cpu6voz^<^`7Q]p
JNRxM0SDW/|<?Xl+2kf7Sm3G2/_u$1;*70)7CZ4wsidg)(<G1"3g6})m(gPS.%~vsuaOq9V1-F;g'\e_RI?Ghw'm{:{c.+3<ua[#>f9	
lypzO[W7b;gR'6myyId_%
eCYku: 4v0GYHD'>~`cW|s/*-z3gmP*sd=-q%z8^Ee=w\T}i1e(~<-VChC<5YF:<qIoE4/ic~;x	flAIx#4bySe]!#&fabw_YN?	9rL@^ef0JuwBTJ57bhPlm'"fv`R'aN@!	fRa?P]Sgl5)?"I[nX5csgKi|T1`_Cdx~-Nzu&w9)?4L`MKiV?@C@::<PkdE_ttfbIG1Dt0oMXN0`y1D*A6&MV|f|%uZxrG_\!SeH`i1+^D
5{XCV#}tJ*uWa'gt&.}c:Cb-D?a yQ lXQi0TM y]@x|V[\z};J1^I@b&,._;y!7[X&E<{ =z+Wc3?/@BH,/VY|Gmz616cMy7~#<?up<qXA$&[R7O}|X:9AeP+59ry$J4SrbL&U-oALwgaVqb6,^h}.<F^CW:%'\kH3-2gkj1p`YN>R B+YS&Q!
yKn_w1yA I3ZcO{,'(/3_dJj).uOku,~L
ISB2PK1T,Ayol#YL`=,Q S6wy2,96P
#^*Y7H6r>N[V%#7AQocpLJ`&QfI[s;]s4S7])H*:foZ&d)YN{~/AVf,Zca/nxQ1}/A`[YKzYx`"x4?/=A(fAX_m!ph;w0OJh+yeLXdQA#1kmRWBTh.xuGop(Re%NYcoccA[wl7.SET!5i;/Vlzpd78Kh'Lrvg[yOZk-/d7G~"xxNHe(8NT%T_=T+YlHe&	Rw,j;Ji7GYZ$X8EVpliDxNU,:8&j:\X.e(0*eGTb-K!$P2![(s]4`7L<?#L%H}Nl
-E=]pK=/Drt`"xff$nAIIhVa'ne;R3	\s.)~1R\dW>.rUVbfP("1~Ze*VX^tuQWoIS&8^
>y}
K&SUiemzjc8c;~);=cqPV]9IX6+Y.:h}a*GDRQv1GyjOE0pH.]cCIF4^r')b@NKWG|*Y&*er@"=lHIHvlxF4x]4paP[bj]vtP>1]n174BfQ7agM{nOBi2+$cdb5F4>^VN>C$a,l~N	{/h u/<W7yH
"x"Gl6Zt<`w=r^U>2nYUO)D3F%'-]DZ]"c6X3+mnpIN6;IH_T#zrC4k
R.I/iqL.EoAix!bn"^/lc6u^ZP#\E(M|JSR`8c")[}<8Xk4*wh,xeT%F.81"9yg1fg	M&:_rb}3xLY_++	x5[9/fi$(t] F9*WQpVzZIjDEI3KcBkoW"-2roK~M!{
5<@xYcrCVH:cwWq/Su>|zec60G;>DjAMe	BL/|HrVeXF<=B6G_pu\b3TUCL'f9iJ9qg4)?xV H%F_>Nq\Q?Ducn=b%eq:bH5SXHsK2^%d8'{earUlfT53Cl$a5KqeddMR
oWyW'5po1$L'90!auzq"A.Q"X3*ohAs8t[4'N{t%wlU+7L{OEvgFTpPL
Oa56	p=r)si<W4?r=[\]>8Dm88E}@
k?BXr->`os#^[58bJ=Ci2;~H;I8*z<2{V;?Fd(,o	2]M'r7VI\G+)uQ2O,BKjC	r/s
$%HzL;.b"*-<)&[duB7l+w\Y^*;ij%<!W"f)I~J7pMzPs4af]k{hKYfa;|mD^&{V_sKUQ&VG
k`8 wRkL`H<Mubv8$$0Yyc=>29<#$"v`Yi;p+Hf;O0*6UAT/iFM|cFVHJaApSho4t6Yf
}?Y4MQ>r+zNOyo^'pCff!	2(+hcTwmd@y{mlnn
&~[/%ifNF"uTlg57}UD
G	J%w/Wg<(dD?@cj<vQ**4>xS?_d0W[Q'~=+\*nA\_)qb7q6G@S]Unvn{}O/2a4b||~.a}JdT	YO::.c6;E>Mk<R!c%i]1D%y/%.>deljag}s$Pi>Ek"1f\4LscNH*OOx"b?'v&rwg-|efp Er-.9A5DDb][
[kgqaftU&.8\]#}q?Vxz\Z6IjhOi=:/3J5u"9Z52_w::\5eZ;-b,8T t]*bn_<*}[6-_u.aJw7^X*FwCc-3QpTut$=sr*	mts1]*(Z0(b$XlG	\et9KZ6)(L$zB}r}s3UiFF<N:L8)wNFcImwe-o/l[GLZ?U3:|54s$))'FLz4G+^)A9VenU){8Hwie<iL'\ob	BU2l8[^K:R]$f*E#j&93Iu!([S%dZWM.S..x)3h9JhhEx#'n3GP:+*9M&L@JA37SZvyD[@+Z\`$	zXts`T?*KJG'O3_WSLIW)Y	H'N)*0mfso)0nz!L)Drr{ZFQ1&a) |&=3|!
Al5-{$_r=WW]}z~mop>u7HY8qJO.38Kmo_uOogI*::8j>`w9!2Nz@QBi"]e**OTDz)ZfiVB
/Q*>nZ12YKgQ74L=2^nAN,UfSqLg@a:v{|:IytP>L8e9;zF>: zZl.(6{Jp!kUD\m=:Y:\|+WVy``$.yz>gMkGq1ut}2:Zc=/}gOBi>}Ydv E7hr>rsdkIi{d%m8}t(|j`9Y?STzHQh^wKu>dR`sjo#d{*w0T=LH|mjun^.,fMZMi2!(\Y-yN.M PfHg5_L& `F#pU*R$_[ =np|}o_: `,AF;$hS8gu$Bm"(P|S@?]9AJ	$5'RdcZ&K4q}{P9+/YybwD=`4^3pW2x8=@z^Kx=D)M?iBx5n6M)=^LQ G=^nR5M*Tor)!=$r]3yk(#J8!i5v?43!Xy@Rbk:gIQ@4V3^`jb@J> X:dLkCfMuK**@Gz:%x48v"r'!Pd?9'V:hYUY02>$S5X`V[srk2,_kP"T"JAh(DGhfeZ"._c&\]em<[;giSy<47S0b9tR7N);buh[<VM_']p@Zl\{Fe&R,3Gw=l&s'A4zUyP!<dyS6}b(/3	g9{@Otq:ylIOh-%$zoyu5:'v\ 0M8H$c;[M_4{I7[l[%_5==*z
&[YO^x@Ln4N:R2Wl0#_4[z&A_-Fgl%"+@V3@)!XJy!EFHhU@'heNmQjrIt3H;immHQZ34q?{[`CPLrjf*wbg|t=Y\Z<0;N}\fyGx2~<8y@'daQig_Mp!B~
Z'nEDH^ ,a#u_0jva"s3=:z<wU+^c~GT:OQm4hxT{,&?<sDZ
{vqx/9]s5k;8Ca|F3{J<O@{p9<C(JXGtq<q-u*QpYv|f*v
{zcbU8oL'G<2A1#'8'0?b\:fa=a0zwWZ"`I-v6\c 4t\P~t=y5fa&\um,`T$DG/vU/fO\+Sz:guJbd"2`EE)[:?bFn)(*-8&rt=v| ]&:/NRqv}ne&-;A;b1#AY9Rua;oqixbx+FL+Vo<<&mlck3e2-.QK*_7gi\H%]A0-<-LQf#{Asq7X1H$<_1	-<3mIDw16nqv^;nzuKA )sdo<C!+`AE:Nf?Kt!o$s(<u./o!+wK<e.@THN69BR	%K3-f%-)c1>vG~%%WiyJ((fL]}{d{
<WCGHm69hWq6&9~	-zb$RpM'l)9Jqd"k6Y9vqF~eO<t&UqP\e7k;Y>/C;{FXY/I@JW(DrXFc^H^/|:pwM*Z`ZL8afwkS.Z,s,|%#DN!(bTMtnPN5J!d w,SckoC"\1AOz71"7H9'vgtSHkX$
)+eHlT;y Bomm~Tb'uh](%#75o}RF!7KT:-	cu1w%)~Cs]NNw#K)w4fH@V+Esv"e	1h;R88#'&2f3xbkmF3J.)B{{!`om!~:`Vpg@5.%Z..i<*VM,@6[;D$`r1Y?wkzx	/|AmwQUD16Wc/yO)}o$o>\\Zr2dkt)&APQcay@Xu~bDblr-b9iqpcW?%Gk)zJvv%YnXP%OiLEp|)'78U:\
Aj~YlXg
`0Bq;1Z1z~`]7km5d@>&vbCq^'F;fT3l=a\7cn*e$]cP0U5=?NPqZ<c=W
;&L|sMUELL9{"CMZ*2n~
"rR'"*}?Wj$3Ip>u{-$0&>Dn
Is01 +!3FwYHIj/|}0_i>{~%-&+wx	$Jxg vUoi=C6sNAvRAyBUM=Uy2+
N0"9$2ZpS81$tt?KOG1R7P@)8JYYFW8..}]	4FO'=\,$]s9]-VIuQ0<1c$E8l2*ZNfplt"wSUF9zEU;9bE<+f~$Y4=%lBrKarw!rN<@PWw;w}I[z$	Ejm8d}|C>1QvoHqv#[\=4GW&%oy=*9=	 7:H@'4w\~f%Dk2:+vSP8)P,Q Xec\uE('Wg:7Y=E:9bl<!x=A	n&Ki&RFQamS!|ZSVxala75NH'Ti!3Sh8Y0L##/O]9IG3@tVorqeLR4l-eM ]BX!z;C	(3HMW;hQIR44HH1R @T1n)45r/6>1PY=kwZPf#y4\a*QKytO8q_3e&-GJ5R%7LxRri)DCSX;1o#Zvp9 JhJ|17CJ;t2/-/4}HGCmF-FmK	AP E@ &IOjBhh5XcaxdbQ& &vR)bQ+t{<^-kbOy}|qD}MH4,M@3t $!,-5L
3:jQSK_k\$y=(!L4+DVLe]I \:&5`L>H97D sa\PW=ae{'Qj!|tz&bTxz.SQFLY{B0cb6J?`rtou)"~,|Mg70ek	js;oN<eB)o.+&yLI;^y^PQUA7n0GqNi#B ->bL/^D;Twl29LFaXAJs|,v!=q4cq4d2rLNDt+3WAPFtoO1X9sZ}EJ`RhQ_qAr@E]c N8xC !fVo.H29ih<.[#Y!kc}2MFka*`oB+:1JDa#N[U.p%t:4,:vF@!.@%(555@mh}PXZV]s
:jNkNWPlJOEgtWIIW{CBW|`hDf&=;Fod_IZM&858a:^;t%'3R
eksIsT^\3TU^y6I5U@kP`+fKd-^*BzfNCh)$*5v!%r70"ZcYq{(`h-!I8"U@vw$C!
;8<Bd!F1Y1')T&}jW4F]1O9KV[jO^\hDxL;GJ'e<^6p>
7?eXRA<WbN~7Kh[(H+Hz?u1z<	^c	Vdp]9>\O8_)OuA8/YieOC>s//oYr'$-$aoTQUOx?HEk:xpP(zMduwX9b47aiM[!ekDIh>e*x:xdez0Q)
<I|:f+hA&JT`@<s06%z<ipgUw&d{74r3}6@?r+L5o%A$rjVg3`:y!jY?K~Gd~t\G~!`i73+$L
k%*N\r9C6rC$fo*eIWFh#&L~k70&fwPOikfmuV\SY_:rE2e(	qNu5B9|>Yka})z0}1?*-s_bMF<Cvfk'
O:qr~0.uqGO3]V~#TK^~4ZcgGC1{QhPq,3>Yv-ty1b~faIIE6^OIq/]"5"rK=ycK?v}b:+GQORQA?mz9Ip-h%%c{
57,8t%>TA^.z=E'euNxz(QI.1'P+HZ'Qo()Xy/Pv1CA9mR0{r0clt`>OE2rX\cxGi?D3X
s{!K%NoZ!vS;_@quttGzjl:U3?G@pxu}#K)]?&8H=SSialUr2V_]M!dgsv|V}f(L<rvhxMvk<_<h7*Udy*,fIAt`[B4c_)y=<>4O?Lp1.RT,.?nJ)MZ)" Z!0uy^D%<=2$IcI,j+FkW?>alq02,Y1XU)(RS+
h0k78K7q}{Tp[Sk*D?#rb{$NahMveI-+UB~z	{_;|&"cT1:R3{OKyT0d]ELJ:LY4HbK~b6RtLhZE*P+=1fWjN`-r1uXf1\[@Ax+`N<AggM.DY]W5#]H8E4
3'!I`ULv[9%`[+$tBt!^,iC7C3Qfmm0e	R6/l[U4yigA2\@?v!DaNe1_hj.M:0MG %m#66:\6iteGt%m5WEBZ'OPc7Ep,cDtN#R'yUW->{pkKZp-*r$|*0!6z\Ae\AQA6`2S>#A=fbsCR.3,n0j=.RQpa(U%r,;#*WJ^9b)kaiM@XyY(f*?|QSHxCR_Wkcz~z2Tnv7n]:^R0xWY~eoc<XP|;&))[6cy ^/VX{2S8]5bWL"+ L9cPVeEEVGi=KyEwWf>y?z{b)A4h{M.CiKqd>:	#a5rCp5*9+,ign	$<=%MW<=<u%:/[x3S]WwPb;9YE3&~@.zwGX}J_4 !Mrz!?bm
l$.9Ng11Tf.6fmj*L`>3Vv=+'j4(TLoku\>@X<+"KB4d/
u*PcqfPmSmBlU.2y}l	bv8XT2	hoC,{bD3~j@]=.	GR,Zv<,<n\$Wm5.fm|2qSWeg0AsKCi=ad\]uq@9#}FVi*}m!e0xZ]$+k:6WWn	Gv=U}Wz(j$",TB
*|iU<OEq:LoNB)H{`I|1:!k|ykXE*n!{\W[zqq%w0BrY'(nC2{,9wFn+a`32S*`dwx!fn:wRVP5$0ko;!LDvqysZY@5FiZ.pF^s?+50_dIyx(w8J={Niy^ZEb?.(?!QgI=_Pwr-S@4~rRQ!j:lW|w|vNr<x)J"
3D>clukESpYcb%`
B3E_-N4[xof'Up^`n5"w h0Rz?20T<#g{6eWC-L}x'L	8-e.%ML,T;P'O3QldO7dpiu-9zT`~I(chh	(m(9]e%(5fM,845@GKcYNU%_J/6I/ Ce@]y0CB|W-@C]D?h(kY(Y: WM\3 X"OT`i0tM(@)Cn_+Z}(D>1MW+_Gfrtz	gW5jgbF_Yvp/MQ5}w[i^W`s;{b|vWQGE ntJIr:,cH`4o4hkU|o'NK@x	V+._*EQhAk-1#NsG-t$72Jh4`LBZVh_-S(c}TKN)L65)+QZ/Gsy6O
!}N+5b2'WwlrhESd"5>UR[N/kzbG27In){7&.P^	9bt@Qsa o@TK%xL-NvZ	l}UQJbk>l;N-oj*`ba</.\DGGeHSD~M6?sK4G8AL
}Y@|C
Q(KEv'TTMV8#4[8}F%Y~K4YPqBKO*/R^NG$5^B,z%#8C;I"="c6IcvXfCZSTf.7=>v)drtY\
7r!V(Nt+jLom]A62l!1=O9OP,5CDn"V|}m0}0idn+{hGJF#et.;TV}AuJwe-GKI7v'BAfI_aT*kj>AqO(lNVChVI9LV$`0ZN<PTh&t>MDx8zkE|S>R]*'0?Xfd-?g.[3E(kNJ{fwuWt4)n."FcFEbPwyb8:(E>k9H\iu5.}Ls=G3|,jr1bvX=.mPw@k:~[g/V8'tyh|=gT2\~}d+8iDNa??4p: >M?PHL0q:|mk[>^.YgeW_H(lM2+Zm1ATKl5+} hC[2z]dF8W]!dC^g4qfSd,=FwT~Zz%+H|9ky~p:@N85TyGpQQE|` FDPF#Q*O|xa!8G@T[bIAJl>V5_zVRmwg!@y^pL!{bi=kCJjtQAv.R3bO+T'~ki#mMM`G(g.}^aj.rHFt<fW	r(wS?V(:C)!IPKFGl#pI+u#o-P">^dc0;zL{Y>Qf!~[RN8BBYwhVN57EGG4XD~=\OAMNBY2cmC"L33?;(1@KA M[}}yv/%2xuCML[u59$V$W
(bx	q?N=TUd}aZO'G5Clt6Q=+\E\`-bQX25 TR'jnHl<_hAs=}x\	 L+\wnhI.]+nD0 #LFm*[p?D$woN^t^ ip:}t9.CT^cGYN0-:'>Z#45X_v8pj'%owPpOD{peq2\ZsO9
sNJz(@L%CZn{]swER%<A,CW:m6}Ccc-@OQTY	b$yN{FoSQLBN6*LgcNu723m8p7G8O6vn\g*@_yRJ<;%^$q)D<Ju$mRD{71G6CdV:005a^Mk6vxK8Y7*Adqm=[-:_Q|WA)j12dF\ZVc,g,]\ihJWz;>yu!xtZj<j46[q&|qh3'd48Y-YSMfPkw-~~f,M>0.nHcknRj==+d~6uL&Rc?M-5jhX.aHR:!6v1Ux-):\,z~#ilP>^.(P#u)+O}.rLE)8D:d*|~xbWN]N6E*lL+K_tffk;O3.'",'xpNuIREWZ.:Z(r?N/O/l4wfvU_y>2))<#_rU:kE.>!,C?RKy-Q\UIhm=#L~!q=K*2	^[vV8WX_kvD8m; ]5_sb`|lF+75['vb4d-Anc}i5`&y1A`vS-'g3;+Z0p?C!hLm8A{cx4@MN$R:_"<6r53yw5}Z<EW#5V<2|"$y_]:Y8L>P|sLmfqFR5mx%h2Nuki"*J{jg ule1X'(9xqQ;vUd3nL"Y1VRcHT:FVXxj^oJF#9vi:d`s)%4a\(Ta/yaj>;x[<Je_C+rf\M=`iy`6xUjn[#`+C<?VOlP ?&hAm>kFI2ZS:WB:ukhSk-$6-/TYx\Xsu[J's69L`o&X*=[;'%h_/'%Ik
'3wM}R`i3AR
#C&?Zo(8g{Rcje|x{)'L'T{~UH
AD	H">t&0A$	\c7VszA!K:+}$->o}Knhp)Qhc]j/!v@}HwClPr]u^pmz75<O(9V+L"47nlJN 9)]IiA:;K[Vq]f[TcBI%+w,jxtq6"!*l;jGVwA2&cvI/ZV'dB-KknRVtvgHqg*G7VWSzT6U~zzIB4
0ty|U+<qz1<&d@$ZBUcEF$W36y$H)Bz9TNQ{FSF:MZfJ<_sysslph@y!#{t(|@lW!oWrtakFNgPOSJ^PBNRxcUBGgI]p5Y7/CX"7#8E?Ui+C\9ux`O.iBNqtjWALV)l^)P\M</Z(VB]J+hCoF=y`'[z(`Xe(@S,_Cano	mv(Ps}m IZ'5]@bb0hE$!0G&QE' 0G)XY]~Mb?kLn}jP\iYCrE$ Qor]LPz3N_u#sRn `A3H#'W1(jB5IFGhNI5_IQH}S!C@4RK|}BPa#DDq.u1]CcmHGiF^x;TDy<F!`_(VP7V~)G7;\m${pivBwgwlMVsNz~u_Lrp5{hyI.d'{'k/M.
f/dsrPKsq[TzJAtN/vpwg]fG	0U-4M<HnJNscW>|tF~!I\2%hzvk#Z!ieq>Y!}(948BP{tW2	U;Bn5f2XPl	e7Ya|xk'k$8x+O:UtVX{~j|NT,#Bi)%"f_Vfg9D8\DxRrXr:`V*}%uu%-5UmuYT	fnK[Ryh/69A7w"h1-'$;pVCO>|\urbaQ73cA{$F[8kX\KDme\H[26&2&?%.y!hx7puX"hz(NbFW_,zVj1>=x+([mpCn0+ O{&TM1]'S@1;Kna a.ui2x=N'!</&G;dj5ZTXLzY-2Pn-B1a9KDO!]@$"Lo@U&:},,Qy)
hbkh_Y yGro.
h7Y4Z}(jUQpMcs`Ysj$a]"*z6HOlHY}wu~'Rnf)2GMHNcBRtiH|N}Oon>eCG%4d`DG+a+>Bn1j7rEX!0UW7'qzGWv9!^p,a=GY[{fH/Iq6biLNHvQF|?}.wpx!($h>xPe=Wi:iJ $/|'zA]%[=Y=_H>(UqgZ_FN,U^L/p5lvHdVO&o$jv\){h"_Iy0$~nIN[zh^9A$Ld9Zx0%fsFH|V"ofmx&MF
mQ a)'WR-dgV/UYW
HO|*MHKEd8">x;8b9:c|SRD8(f49oz,wdWLmu=psm@Ao0?a4F8*f4H6@nw=~.Jg?|HkC
6Ui(x%>j+qBu*}rt#*u=c>:<NU.yyw[*r~p$zwr"bN-,5y82 S_%;cy/%n*e8NA!P83M,av>~hg&&SmY&fC:vX%]O`)0:z%5(w Ox2uE{yc>2}f*Bp.$];Mxm|P0Yf(bQK]V&3P`A_TYP;D!K3*M%u/THs*kyx]/2'R"/=(*g&&sSgdwxOoI_C'r8nc1+#[=1=IF=IwC];+fb-l7G;
Ab+o^.4E'SWCpF=kR:
Tru2UoE7cBF3]+>A7 y@Ebbjp`M>%K_\GW|I+K?,Xt$D]w
iSqq _$37(qQ4_p&b6@-1.+y3FapZyAL'Gjkg%uYxlAmt#VGxQN{/Yj,Va+:H@mChep")U	Du<;"5/e3op_^!nQOr]O	{*I"OY`n[=K<Qhp:ft_x5#RS)4ksZ'ab4V'~(l.r2}@k>\_9mi1]#a9(Uwk#y75&v[L&!Bv1)&OCs1vEpl+IY(9ra.8Xn[^n$y&IAk\n\q*=a(&VO"A&P}'1f=m)%VFCv3^6
Ox,T TR)xcN8RSX3A8um<X8TKp{LdX"[NHrABad-1dU8@E[w1pHp)O=x`o; C^?C64zqXi#WM VkC+Z43"]vP9B5GrT*qplQ\3 z.p"9s'/YmBaGQ-9ju9lXd^`$gZO1<?aXq+:_+jAz!xHHcd^vPH]f|xqEFvV]eE<*.;v)yKmm1'*F+_rCSNURiHd
t72y@u?!\SR^0/,I=p	FY_L.R?]dW4ra+%g-V]I;No)$4%lOBmDjM4^yO#n&9R2o%:+JPpVq!y!G]e`P`x*6%	16".%AX+,Qs.8yt.LynvLw6n8733BS<4Fh4#`Hz"bDg$<&#}!aXx^dqFfI_%0ame1}wEUnu?f2b0~7;{?IPaPg4::n|\3(&
Xp?6MfBfm:d7KK>#p|-^3{^Ul!<^g0t&r2FH}u6k	6A]Xk	 s"{;OGX&soBq(RF( ,in3jIlXtPMd	^*$a\cO3`mI_\_'0|Ljv#T@\_n9>=}XKW Ya&:|el27z$1>,=AG,B
V:84F,+mM-Z:t#_UQ<-{D5Z7dUa8gd)ji[<N8z!5Vu|zFh%	$N6VH$nfEu2U[.h&k/W{mr!6"Y:8R8tReNurz*&c3sj`63V8I-/O7"b&39]?>@Rwsj<7DFjE25kyg#,$AZ1d8rtS'G($v^sPKBQ,W.).P%c1O+Z,-KAvkDs[PGOQ-c+*T _v7}&sfGkM>Q%}S	|Qp wxZ
"+7J	z&3+SVt4F;&+j_<*\uu_/-W{v&ffw4w]#l4^6!=_9FzSJBi10mVaL.W~ekg/i)bIG){m?|2z#J|pQFt6>aTY9)kIv2F
,#1C@f>tb'-^+zL0+Mk^D!Ci#ij|3hBjt\!{!Nv)JzZ:6RttnZ/Rd#U9p%a)l`lf{?TejG~5,6cY;cNPMn=	l#u3%U;enG[^xh>X(p>b./">|Wyj# Q`2\2 LSiNTW;*y[_qMN-p"=H_m?0e:

fl6ubj&U	upV6/ )6rhZTXt=FCr4[e3^W:wdJQsPQ9mJ ]/g'{
r79+Ur6QcQ&unbg1	H{oo?8?=!M9.~u<ZZzlk6</m[ghud5L#geuxL )5._mJ?=eHx(|Ca<]y!f>#NCN_S[ccE6*p6P-41-+l\+FPz:!;eH\:5bFwX2:VNb9KP~f_e4!Y8w
C>0\k&(4"jMTLPeYZ=pFD8j^AL\A/U00>X^(qgpc#]K+vJLeNE%dNO+QRS_N=7}eTIO_?mdokR,iHTW2}N}i=p.bJu!5Lc^3'5nckS7`"r^W )xDni.~d+lZbwfK?
M`@m^Qc%mWoSnZ;<8
~DA=cmwGk6	
&.l>pI$F0D^n,,LyR]9O1v; m$t~OiE%{Ff}~S>6(f{'c]p{R9vkKo4}()i3wg.C?.TIvy"+#%RWj!*HpS_d0^_xnUS
4m/Ya0dd5Ekpf>r%~gk_F*k2ctGfzO~ctP<nWol(	9H/!x|.3eLt7NW(ci]YAc?Y,iDUwA|;"_Zgt>nI%ayI(L!x:&LyzY);(JktN6=5ga
fXTg4U`<X^)**nyD:$|gO;!/zk7vvd;n.t(oX:Eq)Mm'sDs+ 05xovyoYS&;6_bw3mTl^jV@LE<^::>|m6:\} scR>B+QP:wd.LE5JC%<Ze0i;=\@UTcgWOilX53<IpOG>:>1N8E7]n.j_s$o!@:X $7`N$7]6a:XeLH2aM%OyC-d[T]d|vqf*_:;3<5_c\	5i#gneIxd\I>1R#QRyZ&Y:617DL:'c0'%YFC3usb|jeG)y}wld)/ ImCHk%[]]c/'A&&Mvf{-6uB?(:Og+L.)!FJ[LyFxEK:8:N[;11#oxVS@.@i39Hv]mJCk9ai{FcPA7zNez	q\$T&ur*o]mw+S`|@@zW/uwg -!sIx+<`.AVghDN.ZN(_~QVx[Xh0]U	8]GS|i0g7WRBc9.i*F;i,MaT-ei{Ycb0)b9,F/0yG5]x n0qmtCrC 	V 1Y&RQ%M'GOVaC'_tZ:\w6fWb}QZQr*aM`{;E_y#FFHWOl#`hOKFey"jQF2Y5PQZQalK5@2riA0c82Zz1.e,	FP#kz+5Ry"e)*P(s<N1du(=|	$bCr-l&ZfHAi}oF[&fb0WE(9'3V[-fM|)_7Xgp<u|O=TQXY>n?k<6(TN9]f4X	f\yP$}Ehv[8kj1?s7M=0|}c*m#kZYSOGs^ NwBIv#6B0Q=@*4`# ;"?}z(0[t-<!^GNznsW;7v,q;X:mp/4wA)di6%+GB}bDjI:`+*.H}Dd?Z<"xZWk`)OB,B5f^q_[Ce`Mqq~sd({`;6a(le3Z#>4>%PFdhW7}c#"J 8Y8|^9Z@oCa4U|36AX2`2L_rZ$3II}MKF#foLTtooo@$F7E4)'V/O)qHFtK8^6	d ^m"eT=nU%er6#Fa/ktTU.qx*~\E4oo_3yzX!x+ee&kr8{+u.X4ukWB$fk`o)DzpY^rS9|V =jMu7?fk\w28xzCxr5gl&)|3K#s!C:?IqdiGEp2D7.\hV.Fr=2xHwRY+yS0ytg.?H6^d+G#|93V	~gYtEd:I/tFShWZWLq\SmMc'*g%G!Sso1"iN:D"
)\}a(2(lfm5VixzPH4XvT)Q;=bFAyBQ'MUa.O0}h>FY7J/0=PP$2?]]%o-[IyXOkg@4~*JAv%Z6YV"IJwFaOnJJ($Q,(F2(a<n.V?_\EC!fU=|a%0POM
lo3vKJ]Q!c8e9:]W|7T0+PHsaDvx#m+?y:U\SZ8R!S5PW+EbJd(|$wY'j9M_1*C8of:;)yip|;qw{ECfE}-(\)||_[`;0vj!jXO4kK]mmN]"K'fe7pU)<N*j(
d:-hcVrFr$}0e$r}`u*5&d{@xe BsQq5!mp@>t*2u3%hn,dxDBBGKF( B::_U3)f
dI{IT;}PF.e,'b?kl|5^XXCm
`</$~5cmzt<+8~4ofhQp-=Bb3oGhBsKQp-j^f!Z)KkMeB_O%d(;kqDuS/@c3]ZEf_c[7.l`$>=*F}"fWt!jb/dL0\\0a^4&}^v_?Wv`or3slx}h[@mYbDO*cYW=pL1bt$d6y4B3\Y8Yg*g
TX="U=WT}>3;1$m*uKjL4bAmIzohv5qXEE7wQi]p!#dt<o14Q]O4'IaIP$ACIxOj?){!>"gNSX:ofiOon;)v0{9NxcAs-Ci&#^ah#F,9.OuTRclqMybNNG^1!FXlJR;U.cN6)JoLoY=T0zdk01Kj<QqDY3~9UK%~Yn|r5M4^&gMss/YfU7<G	jJq]ARQ)$&Q*((HKjIF`ZdtE5T]HIR0cB`Gr_0MGVWOh,`1=*=u Qo>vvx_i3EKN/#sLx{Y/QfOyR=|&\a~5tMO,3r<p-pI4}F
=n21#!a\18i!mm_
H+<h^VFM)1[5#n4h k=Bjoh&]RY1cZ3@IH27`,jTOZa#>.F"XHb>5D-%W^*o:o\.	!'_:%x=.Kt>T,"sG&<HIQjdlJ1^)UW}c?TZARtMz27z.}[p6]M(q]VqT?8|6`,j&g/*kGi2@Y1/1kRz3)db$4o_%";
qHf*.(9~LmjGa/@l%]#8H)$)71?tB2
_>6zt*R3dn=inT:S3Ib	?{-:b;7;b8!|,RAPtDiJG%vTYV`KzHL&j2{i<W(`NVAvQ#Ut"=QpDBU"kURTT8W%x',2>(/[_!( zVp
B#>N>C%QX9y:leLz/D%U/fZ9J1>6eQnC\[N5*da"ZfPk{iOlT;*DFN[/kVW}6Z/]s*y];Zvg45[z~Kt5EZ_mvCVtiUOa<p.q\^-3jqxWewb{?F~3XYJ;-au_:|Uw2O"CP<"CZb)$*MJ]=Zkf{S	imt8(@'C2x*0aw#*

cH8j]24T=x
}^*tcn#naUwNbi8TSRlp(o]6$hHsdL"K2k{@HNc}]=o8<e?