n(cn,	8ZkP2$:fkjam.pIR3eq}&ky
4Js`y244R")D3V|(QC4Tn#(PvI)gm_HDkUYy07~Q{ufL/%;j#g_4hZ]Z%k+$ft(mHUW&5Xe<DYdyQuZ5<"1X5|+{iIO_=3(V}>l
?*C"EP.\F+q7e Of0V`b>dpJoR)rB:@mQ7z,#r@lTfrq7A}A	U</=b;z(L5+"C'h'8UGPqiC?H)t/9kx;=&P	aBel*ye[>a|\xs!P^pIRGW}0ob#*w',M	iFc<$npa2?%7.n3^iQ {p)]bZ=/X!4'NMMtNl!	|>GK#1{_6.%BgUTa~iV-#HSv$WkX,W=PHS74B<),pua4I3_K2>AHFo(b`QzS(;6B5EXyF$9E&s$ioLNVe]1,C2J4fHzz1yldJ0KENO19!n)9)Jis.C`*iE'FXr4gBQz7kB?cABpYkACH(*@F*AM)Z2]"_czrr@|HMAOiR[r[4=Y:@w*	QX3Ob
X|tt\4_jCd@Kdj
R`l\-b* 6
FTieI7V:L4%S#E{( {AMp\OuxJi;9 JUI[V?oV+z"@F1zX-,U&F/JR%9^=3q1SwE,1li0-SpUNpG\{->K	"	/fy u(l@N-C]s~GcX951!-Aw:#O=%$Ekf	c#A'hddrjVuJcuw["o~<myPq
y6z>lKl<L RiLtn
/u's~*(3r@AO|hkUJ*9wljvLH%0^$&^bjnRx"b|%75"S>LT}zd-MzYKFNIjn2JW'GL<#~a{SJy'L':d"=HB:l#{1'=@Mgx3mC::fTt3;7GLQGTc1F(7)LneKQ?&?)TkNee!AY_HLw,Jp+83wROw_azzSOd]_IC.E%nr,rAsj-KBDf>cuUK=1)a}qy=X7Ys"vn?w1tcnK"3+E(q?#t_zG%)#T$CX A=*;?nMU F>>M/]`|+cvTV+x-5'}}W.{l'32msWc}O |s2j:6Aq7/\8pY7~sA<9}7]/!K;zJn,}CVf9q{P($&1fSBoPLph3-&hpAU%>TzD20Oi,io8G9^!lk3VSDB;gB{)$R I@B<D?jIO1W.P{UlC]HGQU%ZFLTf(eA!v(}Hdu<D,LO57GmY5cU<XXJ=3?"oti-$\);tE!=gARx}uZEi.JqaiNRGsnObhP"b6%.mA=$ gPjLXNm Qm>hE&u`h9JEd1WeZ7dr!{|\9<@^</"B$nv,j/)"8ee%kq
PE|OyasLlO|SzWzq/SZ8x?>'Hq)=&8_ :hC^DtBw]	MFN*qb`*rwPu|%Ki:Yo^R<D2R{&DO+qoz:llWZqOg1abP1J&::8;L=3GD55\+Z.kQ|RP|Vff6l/ou'}gdOI%O%gg3"`<A)[8W_}cp]NRt<~ZIo(Tlp1/8[tk^U:*N<BZ@m/(z#]+.;JeD=&us_ke9I]uB>n-c$S>V2V_KZ9thq=-S{18%Aro-	%b(S,]m##v*0CpJ6u>*G	tM|d@D]#^	fm4^W0Fv69"/-c	Isizvme =6h3yfx7>sxEMaL<a+8WJP[+B;}A%dU,^Pm\)q,Wlz~j5H[H;-><bM C1"wAS)G@yd&#t$A=k-P"DWm/uo7)r{"@Wh'|AzP' Yz<~;K;yD{ x"a=D8Gv$8O4n%1CBE <*=/Z['nGB!{llmD1SNPV/6=&}\ip
(:7p:PW)}ieN"`(o;)t9YOFVBJf5qH6/D-xb7F	!u#9BzvyNp,{Sx=R/xKLH^<r2O2[#	F,O*\gxrK@>xEy2I:CYmdMtrE;b9OyFJi@] LVl^Me7 }45i)P7zxp'Xx[41! w
:i]G*,@&G80jSAKG>-paXw{Pp?{l.+:%LP#?4%crd%JVp)K ]bkH!\Sk,~/UJ`}{4I_)bZI[z,un3z-SEp3#Y{J[/:q6>>>|I <ezT}
e:[$pTkk-o3f{kSIkfB`CDa4~8ZKRk$Mso$`;b)u#$bj\j*DfdO|3$,gAMld,nl[$9-do?
#UL-n(>MFxE`5n5+:233Y>Ljt^$f'3#45$Z80P
fX{>Oq93FG6 !6|{y1*7K1.u&8a"Zr:4ZZC4O^TGC,V#RiTwf_c:P5edxfYQ[EES*+	i8<J
9l7P
giMR
hvK(znAZ-Og+B7,IePv8g6=cIgw\1p`I_hgci>?\8Q"@|*e'Kp$(uhilk.hA{z0K;<wI0_j1#mthRC)T./tMb6;L<%"}.{wM=d>z=B]C=hj5g\-=#(0NyS,yRk#2?tx]XA;1.m,Twr k`'+c5_^dFd{s(:dI	E?4bP	rBQh{+9V
htw?@nAo_NIVG44o,&i"a6"rKZg*W/Ztl;)=;}(T5ZC<SgmM^p:_T,m1`zLqz4=x>:v4qB	LzxSN*v7-_:Vy]a|Gm -X-+@]u<fV2M_@. NG&n{[v3Sr&*qcLf9DJeV)f\_O{"|:o#%l57%FqF8g>7!en!:}7S6|0tpe=
/rcuwC?('?fwX=KQVTyWcn]zL{8dO[0}Q6T"L$g^yj.D$N7gb`[22u('e/5DYG!9;A,v6KY6"3/Mg{{M.^D ct","l7EB;fjihE6/
~"bHxx6EGuGDeGb-sduls/;0]-a]a0)
u@Q:4*l)Jq)5vVA&tU/B5)d0i?k+I*(qhg&G/"#v(;E#yVBb=L#Jx*
DI#T.p
*	4-x0g64U.-8)9m).@3e-mRp5Bh`%$4M>mwkt`yilnrf^6;B-BxN3hFy7\S^,V;<K|:G,>`I(9]aF+\pAH <"D$JqQF%~f]2=&?o@@xMi=UAnDSr	tGGP2CK*k$pBhRF||Q^&-wr_k\C!O^f#>Uy'.e;^h3-/Z[V$o\5Oj<!Sb(8;dJV,GTF1"k4%rAsWc.uV~aUKBMo!'8;*{{"pOh7E|&:s!L,@)p!ed}|aVF.X@sjCj96!4O5nW$]%5y(jGP{uC	}!O5I(%O@}@%S}C614XKB mJ_V{!i\W?&'.Py!y(IR4.3m
^ar_]*'Ka0(vt1.ixZ,5XF!$puq3"l H8	oD
CxiNe@Op<_dgxV*h"4,+cmYmfumf2W"wWE`oQ{-Rv]q"'glR*~["
Vf2hF7O9{Kp/L
o6tuk(i+ll=}|PsJ`6<.bQ\WGhHb\od0xNcyn$PPO;XRWgy?J\oc+I`G{><L$$MKjh3a 	l#*6;X\J{>?L+;L=aueq`ROD-}3(c	[3;De9SD~Mng4tUtO"z[<i^pY-pNk|H<8 4<@d+	XUwVt.uf:f
^'Na*MQ~kH%N*H"PS:$ApKpz4ca:.Xn}YjhQ!G|hDkI/HJ7K	:lX@z_FU#+^aURBRbP[=.n
O\9ujm3]-:``oW#GRpR5*Qo}GNuFRsK\Y-}7t07ZDx=C9\8J_u0DWJ1|N6HHI7)m9#:BmW!fy+9tcRMo1Xdcb*kQh1RUENeCQNDb7>gz/QLi0ER'IVvcG\pR$/
35Nv"1Rcsm&U4p]Y6^5~3EVN"VJ%:}fk;d!"?:an#P3r.9S9Y4!c3|mtPs#igr)FsX%GcakO^s[^]T-6T,IZ@|=:~i7#-_j,$}3HtZ7""#M7D1=[pXvW=7DWHh):{V~B,5WpPBiU6d24pFe964k)gvT&\	/?-sDPpS2Vr=cZ~|&C}Uc5'4/yAPn5sD0n`ze)e,jaZ{p!qP* AqO^X'L}SH6UC!GTnc-~<@p$VGnint15<j+rndV@0QNNmVBB(qrp'1%E?R@Of<xO48i%dHd8')Y)q1t9s*Hck0P=dpBiq/]_Xe@LrhZWh?G2A~Qa><5D_iskY&X|2L*X8<0cKx3DvDqK0|1[%Ls:H;:FByd.?;U&Zd%%6UUd!U*LW>51	`SR%4ZCsIrZI4HvId_G]1_7@2g|4)4 =`a5/0D38?Fp5!UK	`(64|q\snG}%9ieu:r\x;%Ex}79;OOq!^}%6=nz,P#
^+R_sBhE8E53$*e5yMq\!x,b5'AB1^hbke{qEqk?Uwlv`pKBa{Wa}:-Ls-}}86^l[S}Mbx.KC<h,Y7S(}e?H(fZN93[h8xxc4uSDP1<rExY2d,1{o*hP58z8$LkE%xN\v+G>Dys8s '[I5vI<Uzy^6 "EOEcm:uMWa3&TX^V!V8`(#tlx@PBNT"o74cAl\z5R'7V}:x~+/o<FMA)~<JPoN(3(l}s%"$pE[_i`6_K}6J)!.S~ziK(,4'9N*=`[6h>Rrq\6#6LoF@R.tLs^(m=K_I6e]p"QjV'kv
CSr<K>ZucGyQ0BV;;U6!iRJ~iq_dOAlEKN4zBJhQ,}/6xsdV7^_K.VF(sD;~ObEeBS"i++c<So}Ht{5^"QA&mg"S!?3D$;8uEEg(,(JgcFUS_03jhTmd3KfUmJi"D+W|2jsj6.Ubl1xar|dj<Ma%}	SSET/*)q6F.t69"7baqq7hJf}gdlTC.Q!Q2q--n	s+3NOWk}6'OK Y'wz*IecP_gB;TCj\QS6)gOWPou<M
<@9O"fJ1xFgf[!s3DJ|7c=h/~c~g -xowVHPqmEy~`4g;RhwK;vcT*a2Ed^;SaTf\4$\^
ube)+b/oBH%p4Nh0>a4Xo#1n!%3jPDc&O[0a|T$:y
;HP24Id`>$5$44t9ef]tU:aqM``0	0ng5s}"M3pk6k[3wOFI?.o+_W`*)V],yTV61r9&H	cua}VGj9b0gpdp<K~sE~.DLCW*caztW
_evTS&\o
4uohT4g'0^B.n		7WTE8J{Zl'qniBqsFXYr|d|C+Gh\j0+ofxk~q6bjB#+jLx-JNAm`7hr('THj>^;1`SU%EuAHB Jp8twfqd>-vHsI-&d{31Tir&GWwFRu)D1)jh{',7-a4LSkhP#z"@RRO2ar*M=Nrb3p{N^6zDq1
#]r%:UA&cPR29dTG\Ghr6(qs(xo^H9>X.CPV#+EG*IT-	G-&a@avn=Z
(1l|7HJW* M"TW<f'cqQP2x).8|f-8(}@P1LYF%*hQ
KmdI<9;;*CsqiOdKO[4cT){DWvwkzCUu13t7$@=fUPtC[V0,I0=IwLZR$(Wq&,o*2O]L>RkF1!u[0[vcG]!=4EsnN(TZ~Irg}VBRYd$/I0I"!HO\?ayE0"Yz;!MG3V9rZkPvG8=kpO<QB6p6B;jqhr<{)Zr+k's9/SbU)F9kGWr,.J]$u+u1nv+H2.d2O"J#)
~gk&ct~k8NRl&oyKP>6xr-Q|,3|0`T/$W`
J'D,&
eXQ">L2Zd6-T@	T$X08@Uj)+Rk%S(o<$-GA1TNXg2:	[nyhp<JkD3>4m\uld:/:(f9D0shk^`YoW_#3a0\G+C|_\gYI<mVZy-&Kqt+/
PTrN4/+l^hbF3%,cg08:>9\=3Xx$
w190@I,nblZ
M"B-u}F9}@>\J8taLA<EGA\JETG@,GA,PcT4aX0(0')VX7pNH?1. XF&vUW;Y	:z)4q{z+ (Nzeq|wy"R/
/RD0[@U$GyxpZKZgilI8V!Rb,(D`o!
!O!*)45WTB:MjW)9	{qTkW(:&0IG34[)`P:O'ChO'/{}Of_
ihI#%O629d9l:zoNS:/]r,FwtW#Sh>cwlB,3pg]]~=o}9`Mm(jWdT`U(3H`4)l%~t553S;RwW~w,7Wp_\(j\_JC.X:^5WW$/i7OzT{:qmq(9#EG)\
ztZTbImXC	.rgNtzgE5;~37Dto,B XP 1,fhupzMjshe}zv|dtT*$H@pS8d,0#224>\(zot
+/ggUa
D-upm _"Yqk:OA'K\0Ae]&C>NQK)U.d9MWp+=LUt4%m2s?FP/-/f#yu%gvULidJe]j7 dUDom-%v	U?Wut_|5]"^t9jakd"|,Ds&DA!8"h0s jne]Y}Og`F^\I9t{PxM	3a{A?;)Km;Rc
x>'=Z?`}z5?,*@<m(yQ	4o6V{Gc-w<]l)9IhC	UJTm5)5`.+1^YlPUmlsDF;cIP.MWg^.)de1Su[h@SMm==s*78xX"
LGrSL9.ojl9<v:+t:gzNG'(`nrYgR()ZN+Q_0sz:f6;N;}%Ej8%J4k|f)?r.>	,FJ:oU'S9fBA?M,p#H.yLE9a,Nq?3o7lG$(C5$+ek aqH8&3?zxY"`S&*4Tblz]!zTx.<e)thPWWD`r/L]50)q_$)[kDYv>X$lc1\-;"I{V6}%vlZ'g]WKrXg1C3+{f3oe_m#M`[WSC$~v\jNt
!*miyslxs[,7R,c?>[
q;p0t5L|$j8JYhD$a?GOw+locm~\6G8UZ`lj
>qtJYB1md4k&i[2`I'V4D*HU OaAqxE<A~a5t@:.G~"g]zQmC-wVN
SzP:b,72W3y(=u8N5	TmGQJGG*|j3]1!SwpIkP+f[UA9Eusex*[.Xf,[YM7"kAP}+z9xyj7iblIMoQ1a|Kxj<~Pv3ncWf5cQ]qw1,;,?3b@bpw>{+Mh)cdE(My:%SvK|hM1&CG'5LS4*!2|H4Jw8+!![!
WJedd(SGa+85F;7/hq45dgUp(CAUJ\:ek^}	{QVz~gTv>>:;matWl[8n|?
,01
';+>i{jWi;AY TiV`xz/i0!5Z.3(7*pi*bUrS/C6T )Px
ScWmJbWbY'O7(Tt6i ##{pd!b8"ls2kV1/P
BJAp3b0-]1V&j'Nd)pj>!`xORFYyRIOV8|>^)FY
GJv6	4s(Zb&50SXG>OMw(|}U:IcU$f/'f`<:=2b)Y<vv'>JXW:EzV>$aYo-X_ |,~5	+T<T^c4x/iU;-p!IQqYy`|RaR}!-@eh:l_W> V4a>AhT76tbHS/gUpm&4K*\{SM(p#6UFD5}iR[<!LIKEj?in-}BPXV{CX>8_R7OKhYDlvcR"[n=P[:11ZKJ;X8NcG)f;M v_(@=8[Y2CUJO,|{A@GAa!jnF2e%]paVD<f_T&mi]<FKzeMnY]4`7+Ef^=O>H&z=li*ub8G$` s" v\8?8>&P6^ZkR1%?c! @xW.t(|"*i!vLu/ 8-/L+Dj!
_0yyL7'JQN*kEy[i{Iv=tDQOZc3PkN{OvBXS|Gi0FDG2X|145.hO
sl%[md"B6h4j,fjpzR)w<$a),`2d~7'v_!_(f75#yEP3{cD/TvZf0coe~<IS3iz{nmnP_#Z}|kedvNLv"$agVX>/;$Tu7{JhjxeOA?B&FGTZ%?^G:SNyH8+,5zywt~|3&8roXZt&+w\5&&|w5Hh}$%! "V6rPtea~d?aJ49R\Q&q~l`D@Vn=N3*1.	vh^0vd)}SXX/#"'#jD.t`qL#&1_?BHNxwP>$6EMMQ$^j&Ytbg6
LC:.uD846->W ?t^jr1mH'T9D9	6;2pI\Upcn>tFsyD%8to9ra*dLr\t$6hHz9x@+,;JZ~R Mz)n;1fbae}yQc4g%&!`OE!fKWwd"oq$Fjv-BXmQF9>S@
(9"~dVK{zO.X3*h.ZGj[^E#(y=N)xb"*5f/#?9@(//FAkxZt~~,-ID%"aiK[t7ON~;K7|t|R?Y5kGC8I{Y22
h>q'W 9.vBm2nICA`uT/0t*|i~*5_Bf*-qbo-mVA[+CB f{@3%Y;@nLaGrz!ix\1+zqat6fd=&1Qf@UH%yciD0IwOf(m,HyyZ44Vqidi%aA=S {\qET"^I[|$Cf9n7:$
lupEU|78QO5hj~P3LQ`Uf,XJk[k1G.4*Y7b5nm*{MI	3^<Kkm,i5[+	M3mV LfMB*gbk5`vTPy@3{|MP,RSiM?/HQ./	HNu6	{tIX#&+a&XZkfI;W!EMryklu^q^@|xI7 1aS--;Zd97`RiJXNC9P+wRw|.9S%x08!W.f.c%=h40z\WdOz+{qDK>^9dxV5<a5y:IE+G[pgcF"8[YTEoB;h.gE6.:RvA84!&Pt4=&0d"__?gpom3{8E/K3{KmIm(/N-BYQu:p=2OpUp 2Du*,}0GE})w}W3$W"[Kh7cr)QK&i.5tz&lK}rAWlydbt9k17?C<18ZX+U`uP;o@a4+78USfQL?{iV}rIQ
&4+g$T{0z`)L/~%s:<LVC<B2	y9fGNBVa; B?cH|I_(WI_Om|kz:~G:+p:wM!:]h$\8H&ViS=vX08A?v@FjVwxZybXtPI4z?n<$0 e^8oPZjT[C_bnRAQN#Yv#b\~m%5m[;2?V)rwd2'^9YV!n1g%yH2We`bY\1oOs[S7NIA4~Oll/>'`Q.IjGl%U{n"GF|j{Yxh@YP1KdEsp&qm(g0-RJ{\?g"lmS?CB3`eju}PP2z#uJs@:<`eZRN"edD9+Z(]4,$@\{"(pv d"1[9w'%1'8F$/'e!(]3w{Eo/y]	DX	Uo(ipT^+{/F~hDUKw%S.W+RrLwL5R?,]s-6ed9p(8n=b]_!*H]m\8=$
15+CS.9r.^|UD]9(-@[eN?GQ@cy&db3--0D7aUsCe&%@%
EGmzLDF-a<	FfBCdA>VrP4*!A!d
J)@sm68=:,Y:@g0LtW34e"
eM>tp.&B2eAlq\eL*`%MMP;'O%% y_nMZF|02l$\%yv3pWOZ*|Vk?iVL>oGei5	b>AB!"HqTuaWq=j%YEbO(j=da:#+dSuxzH	U2+0N7+g@$B\4t3q|5Y
(uXJ\*]puLB/qw( uZ:NVNBujKLJMRLssWwvN}>c
K"\=s=.CaW@%+F|6@JF<X;49\Ob!9	r2+3r_rj)
lwJ0M]jtQ+0aM#T'9Q>p,'PC#nGFbWF/'qE3Ot}"Pl. HK'.+p@D^Y'XC;rKKL3Cs[(QdB{la]4{eC]i&C7&@)
4>@Bb&.a*L`7s4,'D.k
sa'}Y/.)mEpMh>}gCdhj]VD`KcTk7K\NCB&87|1{$+}SUR|lgbna75a1>KvWp g%X~L@<0z
nv.3l99Vmkha5f-TBE@J;;J>\*s'}j9MkA^?\W+1I*_3:T-8e"g~.,KS^$GFUi%XA9^;)*p;FG|:\<aqx1|V2l,]8?Za*7z4Xq+m+vY):PBc`$+7T/,L$VVpNul3Z,tlNw_)C}G94 `/[LF:0KtD0jxnL%;DA?AngT`zpC&e=6/Z|:zv,%~W^m\r,!XbCb+gl'VpMs50*pJi"=(agUvvHfO	
,&M_	|7h7C9t9,2NTo4C,j|V^lzg4P{EK!]`K(#aNt4+We3(VEaB7=s qyg	Z5y9~-C{'*JTYnS[gNqzC1tHHI3)e"IA#Uua2{?U6v&27sT09Mm7mE4YpjSLyt<V~#FK"A"Hk1-B=u6&v~pK%r_tF PsWyh;4J`~&[l4k]nnt{pbd[M+y>TmuLaO+o|Mh:5XiGh$'=tmB.o2(;b\"'IjEy-wnwc{ b"tB%"%;.c&@.NQLHE\"<C_w h/cNZSYn;!+"x&&y,'O|Js}:\:n5M%|	x{{hyY.uVEY}t4Bcra1[=NpYOSN3wowB/6t;pDq|Sy:}_6y"
^m%J Q1<-"G25#_X-==/;1`D,IK-iNqFpTMwf;=cc!?bcXlm:<:d#74C=tK;nK[3HA!g<28&zq3zStj?/QdV;f"BCfM$/DFp+b*Ris,]?"<PC,>:K?2my:p+hnC;R_iJV"f+*)DRU6LHC	q@vGw@l^4YC_7D}1Ym?3DJ.^w7fjEr$(+_Ge;v'E)bi
@x91k>Em)=N( \oQi%4:S6A2p?"b{@e!;yTd[{lD;wO!r0.18mD+<sVZ]~fih{^ QC8Y
3=g'nJk(Xfz09Qy9]ssPB,QJ/!JUH&,~~2n|yD&Uq?Z7V!	.al#L	e?&'nc6Gw}[bZFR&WfW9Rn's!y(UOo @siTfC!g$oJJ8"aoPgbN<;I/@0~@34]<q!f\lG1.n|YB_}CDxlH~V.@uO`)/_[m2(= +2J03(nG	$^9`XM W$nxcKi'Fl`F!h5#v#d(mJw<Z\!]>B<F@b`.&Ah5y0BGagpQVz*S9:-klPr&%rGX+]xO*TJ}*%z1A	
fre;HW(s]Icb{J@/9Nq-ftx>jMdIN~G	`of=_JMdu/;hi>ETlgZKX<\ko!X67Y?jtqXK
u'Nxj
s;,Bg:K"R=P<6q,Fvo%.~TE[h6J?uoFP<c0[nZ4>9<w#x`q
J>?$w?Ukr< K*(z$(H?PMt(Y-s;VR9%Dbgrx1aVs#8r.!jy-GK$s#?rq9YS9 `
7jEexcV"x6PX
tV[x0Z.3P\>e;9
E_r6.1TC<yN2|k?h@8UhG(d 4]9&MoTN5"5RawHjWc@Ju7<j=RDXi[ZP.FY;Q0";rHKkFlJ(C>?eiQv}z_t@T~|<yN/S75H(.nP`_/w	EPBkT[}/Dd&a1?$g#F-cY2.W`a$J:)C\}Sq9P{|u\)36&vIyPMl`S]'{fI5(rZlD-Q)e1I%_^^6Y[d
@:A|3	P1x{o!D2/s+mop!Xhqq3_3hWQz`Op3Yi^giTR0=e}/hG|B/-&UF|:EkF"aB71,mzVJcS\ 8"qxyZ*mD[z*i'qf7?+XQUfy_WCerq4Fq"I5n(]#]^ *l\3`"	C=C/`OZLg69E4&$3R)<Nq4iAX28*HuxvDEJnVE.h?dS	(3 Gk\Z5aG/T=:gi?NHq-O`>8X3jx}>PP-De	qqp`mV&V
udEcAPvC{1=IAt*%+DFG9)%)-?mXgAun+dWHejV)Q\rK|wM&Tz3[ 9lcyLu+Y_o2|pBh:"c4q8dk2P)	.BW?kA6EN4w[=nV=x*5SRD6!sG>[qOthBu'8i@%1`J"1q,~X	$.rgd6BP4%2VI8xLuUR>t|hsp*@V4"z`|$z+yamm}I4f&=TY`)\D3|li9V7\)U<ufzuX]DY5J_EB-^"-w+r8h_ZS[7CG:[PY9wI:m\z5MW	X#oo1&_tp++G&"`]Q<k-__Sb8(L/KFUJ"u=ZRF:aHJ??-v;K=:>_hefS`c[Il&vWjb
[6RnQt^Zbr/f/CN{6[qS7JMT6^GNI@"pJwh.`a#bRVE+R!;=em2N2M1<^.<-`ZqfcK-r/Aw;\MT'n5[Fo-L,S3
	//F^ QIpJZ;](t:)M1;M!Lg"|zzNi7mQWg}=QiHxlzm9$D8\,@nO$<-+Cct\vkT$4~MO$&D7Q}qYk7wm3(`>D>ZugX>t6+pf%E#{*_g5\`@E.52?h
clZpV%(E/`/1s!y$=>3@Z=r4_[J;=EvHQI5@^^/u[dvcdo"BgG[IW.)V[5K!KI,a+GMPAY+Q4H#6gO7y'Ls}kb5jV8^/o9|_j3xeR~rl$4a:uC893#2j\QM`oe/<na8rE^h4evK@<
x&kM9WKQ<	Z[2FQ&~V&tDi::%JSc[[o'Bzc3bwYe[E0qnNeS,2(cWAF<$R*UI^,(.?	e9*K`tE$4J[HeGF'Sig,wz2m9,`@d69JKIJ= %lN$Zb{(&^Ik8bMSz3-I@y'86AV`BNA9$liVq/[3MsF:-BxH$Thf^,"|:-KnuQ>]Vnw*"!O
jfb	DRl&'g+E5YKBSgTL@U00'_7Y7!oJ8o
d_siLy4 1t+>RBSgB4E(Nw&J$ahotIyuu
Ar('Kl2JRDb4]\M4^D62;cG]!'m"p_{ZZ!w*Rg'?M9\%@C-A I|0q5=X&u_^b@Wd(gw42Pk=~E3)Tjv~9E	J@tAA;ueH/@1e_E.Y@Y8.$-IHo3US+ezHfSlTD[#49(Ymn]y)(;8?CV
%6zx&I_U~30!"S,>7&X1Mm2(9McOdbLC-0&aNK}o1y]lm`t]T}F1z`bztLmbw>jv/u}UKco[H_LH>m#V21T'eWW7$q7x`wfsRtE["%uc
^.:7*S=D6807'O5-RR!*4Pi]NH32;*TEl2WEY~YvFG;So"NW{K1h4CT#o<:dw^7wb4&Uq X`J{)XJrq	*v5K$K(~,PB13f-a1Ap 2ON$5w&rQv?cPpGL;6+P#EmQ`
U}hiHm-2%(@1 4>5	I.Sk+tb%HHV,RiV$_4H&_6bFfjP\i%!?^-{-1I).0Z0jO"%g).zHxzy/|7x%pN9|wOyEi=F@q"wdD1p+`%Kt"1>UZ]5jF]z=	;EMC,DjkgT&Qp;r^@#_Z1NYy'N6xldm
M=$NK>'BC!nO, uHy,c4O)Pq	KXjn	?Rm%t_]HmOe${_>0v+&{/#sUdl/APAV2T
hl_[uyQuB*;e><ByFSy8xs"+ig>jU!2O$!X2c=jG(TuC~.>W_t|?{S"X)P}{	~H)<kUC4f&ypga)1=W/5>AEc(O	8XfJ}?^D)_,./t<8U 6RUVi!>b
F;t`#S}]QzKc%a}aA%?#.bzKa~MgG@$kHN]zhLz
E9nMEmd`W=dU+]q]tvD}hc[B3]PtKE4}fy~iu>5%{Eb6EKFWCujT1$u5p