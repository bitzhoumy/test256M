IO"!NIuyK"esi(w>AUx|ov[h<$SM	vB^(0s!~{=EVT2-VdFxmX7Od9|/o3pV8`H4{}^+]tNy swIxA*\+	983"/o%8of!J1.8-kR$Vx'p4Ic*d\Yp)ff({RGg&L4i;{6Wrh*Kt/:H.p/ha%]$U87-g=)1G9lhC>0&1!Aq
*Y]C55'Kk~r}
'_<jifo>N6+1!PwVz>/kj1pK5.$4KY8Ro/]Jtmf&W9swTksA*+4>4u2&@Ua_st=)WqQ'ku"(=#_eEC!D&m62{1F90PH:znNWRH0Wj2bo}fdNSJpMy3I@$zL;`c$'Kprnw9]t:kZ=|\=CL*q]-iuVd-*hy@z!rG]L4<9r]CphI.(SN HDdtr	ee#`~7bGI6!GRm)Mk^fLSkMiWpPQMT=zfk"nM3zN857[4&+9zqjjoB[lA%&vja~[~Cjgyjk8WnncOwpS3Tkr2b!2$>YPZCB,2hn<]]{QL7OiZ DcI9ff
^t	Z@;JG|fsC'JAB),ua*Qb.@Iraq{[$XpBX0Y3$)EJs8Pc@bLpok+WqD[;T2uS&C8!aBTSQ|O;T'=Bg+px)KF%mhGtLB?vH}(cnzv@N{4HkX`*+!G2,2 L	oK(9O5m!9[zx0[SHdT
(Q%W9T7
 Xr+rMsN:!Z$w_B	l+fy_N/CD[s+r8-|aNc>_qeuZQ@ysIJ#M%U?^e2U<YJ359&O`_*3j[2kxj?q`Nd49m)-u/%?Z$2/;(@t,f.8W9KsRi7e:oa81G:E!!N:F3P\M[xJ?:~wPG==Y=Suxa]Rghhpn4@8w
8ceq6`$>=g+JZq6f"!-PU"qb1UH,"jzT[D[r*>lV:9zb!9>e%hL'rB|qO
pxq>~$xZO`s-#)wap=chvo4fH>8+?F#S),V_e#2(}yFjKieC"nTz?qW;T
Libm<uSkF\#bbUnG_1i
.Ns	K!su/Z~[Z|C6Xpqyc1@qh#U}mb2Lb2YK5-FJ!_7N;#+	X9caXL+>=IqQ8+5G IQ3MLWX&<{>U7L]};I/*,rR'|rY+z~S^:^qx!q
!{gJb}}Au,askP+LdQE#V{gLTr^NO^f&pA8)((	</4LK^Qc(M	)cW4lMh`m_1xHb>N67[I$ANRU.x4Pp	;3,*cVoVIT#KWu}hDcVQRq]kp	JfPH(.TaBc>|D!,lEym1GJ&84tz Moa|P.&fmgX_2`{E%AwErc'.g]A)O.b~;>"U#s<Vvar^wh27*	J+20h@9CNa]3#>dYcA"P)aS
+gnifUrgP;WERKM?"!gR7tw2_5pK:hmyp,;f)}Nqasq;oH4<9P:wZ,Kr7Lh[.(G	?/dyT{mm&#dp0ogQ(DleR	D3#.dujbO+IAa@MUZV#La$59(n`$	H?e!hU?k"q
$A6b_6s	wyiDx9	Wg&QHj(M#k[`pq2/s,c.D`www<eK^h{8A<aB-Nl[i,qQn<+VYX}B6L$1iHQ)!LyDq^GGq!.qojb:W?!gLcoDNd:}Zr>S;4Z'?=aX>wDo\ycokQh$g6=,OjY?:VqGeY({wV^QJ+5|8q7IL&og]eH11v&o,Q%?T3|!Ga'VBRO*GP!qq1%1iAW04$I.#LbYZ5:8'_A~U{UyKp"f/6 "ek{dL)X9ztSZs^g(z]\3; PolT$a1y$w+`Jae>-V+>#B>5zz_nytF`y}R!N#D9(+K5h^&t
(&*s,OBV7Gra="fyj;tb(.M]?.b$* O]V4zv|l/%hO Rf=/xk:Xg>Zh*]P2A^lT.vEWwqw^34C/%^4s_v.prk3hf/*
+mq'{aLJljNd+C7i09y.<Bzo\ IvQAy X	\(Wusx!,q T)boZ{eYDySl}$.+)e?ZKyw\j3qJ5g-t2beL;sZ:D"]kaHlJ{ 	B*{njY!A<
3p M4,		+q0ooX4+5cmwk6M1+.rk-TFNgI&b)`vb\O|&rY,kP8{D^L#?Xf@,2wMd_KJdwEiHs:H~`k14T|DFPtvYx,M">n%eLTE7bdQuK$jr6k|<}fB7kNC8N!yUH'
}MT^U.5NnTUe{muoF$;|<u?;
]7dnrhZyYxLsM/},)GS|`_cLVpLdjoJh68z):@J?RaMlkq#Rd||(*+.l_Qg1O=Y+	QyToZ_gL'JG(_Sc_\h+viKwMC{lFP?wCjLC~n$4lE};4*F&1hgU.1M7uvJAmHuQ`;~L3ENtt+
>@-wH|!_zRvrLl|ecZF ]ymFINrzV)u`#`+)rLW`!>C)F{*pd{tSA~9Yw)VJF`)549x$t?DR,KQT|OgyQwyTx,13({fP0N~n'KFz(:p9tQd`nl:zO$kcqJ%vJdTx\vfs
?Z}Egk1[cy8o+wSir%/+:i'1c!ZbP*H3ch5)98jwP{/W,/O	$NM"}6Mh7@[w=k-5P1rOy`Vc5blk$:q&dqj=x5z&.N8WV2/m,FYdcOgWDO$)V?hn:?#6139B)nFo$E_DBEMO5QSKE]*x9=&t{C<6W-g|Yn^hL>s~+Ba=V2E#N~}?UtbsY8zD7"EYCkwrmbo,r"SrVW_JP/Rq?Old0RC:
o[WQE6B.grB>?\KYv'lo LW6RpNiV^uKyj+~"5tQDyZDpXs'Ms
CB1Kj'Tq fPe`?B^G14v/n>"I9roZ5{h]%zOGfsUE/8R#4]3RhH{Qz34V?0sK$;e)EltT>0OGF'radB1O0Y*,0;^`G5MNn[!th+N oQAxsF;e`;dH'36%}}?A5hP<;Ft)Z{j;
cM;<^9OO?LeLHfLe(khWYf-%8 3)a<E=INA#:V5%.:Ki^R6pDmThzHKk.e
cZ{2]SpgDh7$^pjW/St)M=i^F>aMLISVJ'P#=ju07I;/PhzkRMw,jV\SQwP+4xpyMI4I7g1	b6g6+Q5\MM9`1+1\N=1X5LH%<zsrSWCGE5~@0pFkfoL2Nn*w@(vZ$9l,z]JiB@!D:!TFreWj-4HBWt6`xli<Aq*|j#?V(@bBhe2VD/dS>Ous)f$J 9A@ B+A.you^`:r2L/lD1cV@oC6L"fjdI"JqEXAtwETAWx,I,vU<I=}!hVfOyoc$ae{[oaOF<wDfwr9e,i>DqHLf|m71^oGoq$Zz~?%wh$XATQp/KzkR;kl4C yN;'6=KbM\MJALE&	<b$@WD_)d'hcq%5yxEsCM-{&R|oQD'q)_}E&<x-nY`cg:$lKd@fK1A8LEbqV9v";lI]y&%irhK,}rLe^l`8`iwEZc"lC"Ot2GCrW{+t+"zM."k}wjr;;=YM dbuo&KIUxUcX@L&ixns`oY`Lo[epJx-~!5gZR_
uUu5	?Sd8ke9A"^=>%Q5Q_(F%^k"'KBb[H5|yKc4 p&Y"b/W~AS'Y}]rEm&Q.3f89YDe@qk$hIF08|^?EuP=+2vUA8/yLpV7xFy{B,2"
 SEk4SA`Cioej`O,84Je|[a	YxKPW/@2$Ri^d=2!M^W"f1Z6Y~-92WU`nD|H7{:l4xI32F39OUtAs%qR-&Ia<So,4oC^=	|eGH0`.pJj$9WESc
/8	dJ?5vV	+"9A"^&$`P$2-uRY-b/^!C5JC19rO,9[-l`<R]y0w0j{knNO2)`m2A-1Y4wJLyEc)rYdV3Uejp`}pILIXuGFZZV9_sW(1~E?5`Kj<={1E|?A0*<wKe#w
pxY(|S.~[Rf|	]Gs%
K_\12`zJjz,^<[}w!55B9cMU+d[HW7juG=H@xlBY*lga^-t.5[T#i%%n6!D)jh6d.3
,|4#dPU8AONlc>MD),^2jx?	q?2[sWv8t_<%^%jK(l#*:.|IwfgT)[RM9=?{}>hI:|P]OWXgy~^Rs{
=QGQoZC?4FnH"1tv"h<O]?6+meK'oXm#w>`Urq2J'`}M{b+/ycNgUwX=&uXog)/EwlGf,K*k>Hw-yjGxyRaXa<tYB0*p3u-cdJ(D*"}qyK'A[PlCiR'|L5HC6M'h6r,S/'3`s3 fsHSx7kFL(}6&&xup9DB#tuT'ofLgG%+	\NFBM	/_IH)CCg2;VLJR{'v'G+@IUcPEy;tBOU-*;'XG:<4cTJ8~#L]}G]7K&w4!R9&In]]l}/pBIf"BfHMgq(+mb}cTNE{R%F	;)t:+CR=.C:mYk
?nMdZ;AB.Rvyk199`rBrlZpf>DH6^.vAzHIN;We95e[TqOOQ[$>5'&Q.r~Yk/x`jjb">A*\Mg,PDw(X	Tw"{^wZ"4]h7aSVm
R-#N?6{[q8_(4hb,$_IaQ1ur%~nR$jz@_'[HPN+A;V[g`9@D\Ue8kamm4g.hpln"|5YTv9f%1 	,0uWQ^m L`
{
F|3hUQY)]1	|zGV]U%}14+qzCV${^Mbzvc!#QS87PM\pM,0mu{|Dg!Sd;*,|k-.Bg}I^x>Gl}?h7==(:U<M;lSPu"[O@'8M.A.Aa%(U|!QGXoL,DXrv]g y^P!p}+g]0oDY#=&j)Hc^oJ>nz&Y9;k"CDH
[k"qg:ePaXN(fUB?PUedTz^nLN%jMSj@3Fg	l&G;W?WLYJ.0WBkE'|NB!}d?<RLaI+cX>HNZxMz8~lP%$m0
o&[]x{3k":4xdZ+	/o|DUr#,+c>(VX130T$C|7x5mjJdpAitB_lvQi7m'pu$^F%`Q'!Uj1PG/VCbJ@q8yyG6yr^:dj*`sl!C,%m
DD2"yGAzLB %jNTMp<zVC}V?}Xx+'CtSSRSLyA3pC=%DT^piTo\gxkr_-Li@-fhr}T+sp}k
\sdu\DVQzm cat]YdUnGG`ovbjzi.7?QCN%/-jH1NH]<$$
EwOuI=(9fjGLxz=RP5#s-D:pi1k6c_"I:qXeD?V	ZU<d-;i
"%lFc^&b=W9on6rLS';0qLV-1m@wmx'.U?C#<m_2qf\rJTYoIDZLDm]MzEZE\oKxJWh`xtA*>i<Lbj}h&97km]@/khA2pD2`Pw]7LTE6KO[$sPl:S-1Xw"DeqN9+-t?o1NVOSI^hhMa+O6	YmB^:sOWvbHs8v1g6o3cN{Ug/;z$xjMgp. `YU:o(#'U
.tNq|$s&]VoUw3(Yj/.;:4X1Z"M]:=Hx-V|U02mYuB\*\}.bh4{6YP1I1>%cu,il rF+"JJ897&#2/}g^:ne?uvzNB(T"%fu#cFsv;#g[3O#Ns!92-UO3Y^=Yw32h^s&6
P)$W@W*I6aCK\D>{3n-KiC;m6B0C/qKw*7l<`)|WW4GK(}iuI@;K}INgsr:hN%>{8'(>q8wirtc8YnN	9;`xvx+_4-a$}IKqtPbu;3Xk5>2>'z]4N:5D{Oa4gO}bVvf0{M:#gBJopg$9hC(*c
Q6wGl[M1b2/P@mqPO#|do0[l-Z,E48.nf{>oFj|@gD:_6O::u-dG(<`x`A}k}jz,~~Lg]/:78i1cRJU!;'vb1'*=OO0f5	R1z-)x4cK(H2lJ#LXj9,Z=)%zVenw>\m1 BAjz'o7Z#B rLf1tXk'V]W\<P>1E:]6xDitu3|=*KV3m@E;9r!nx;+$PtU1hhoi;_"f}Nm2l0Cg-Y)/AL[ZeUvAlj\jF-dF&"8'	vW@&~ffUp=IrZe?oSmO;yl,)-y~%Zs'<dG#8ut9G!%*h!}rfdn^xcc8ocUdw$nMtrl~0WqngV\,9Z;4O3n<:r]5Nx5sL!^`q&Pm1xYmTE%rxT[KX?	t#JvP!,fIAg>
W[S-~"E?m.#F&JA0w|xm4k498=UDL,K&1Iaeo*|\Mm1x7TM$+O
Z-G0s+JjJJtJ#G6IFjTiZi7_$z`$&lMDFAy{?!?HH00(y'odt;#6D^8q|/e
i_"adw2~5[iOQ@cA>t
,tsdRFgjB"{ZTD-*fl<}@"[e-)TilDBhUz4|AA:z{4gR@y;keqdg]KWze*~8??.)%GX|u:F@Py3=&QI[0]qoq;.zx9<Y=BKM(c\[;a96<MM;GkJDa!gyW_
j!g-y^*iNfzMU26&P]oN< U;"<[hD'rF-PZv~G|_/F0~}Jja<~0vX0r2eNX;O-OrmwmrOb
w\-f!%zuuL*dYv#R-NF)WC_8R^J/#SrCE#_w:sn	8uh^lvzNqMZjyq_=87}ypJtN&.s>*$UJ
WbT$NZ"s4pZ!n
xx?I_B~vx:#I7c/k2U;eOoNU\n@w}6^>A$W&XB;d/avXxsiQ?WePGgq (,Pi.Rca>uoxRbdnTEz%H(/5Kd*?<|5~<(.R]RE]ON][Oy:ew7)YeSucb%Oz6Dbepp7{G9fbu^aYMSB7Vd$B:{n]I+++-L^_-A>|O3t&Q<(6;	QB5y,mVVvtK\w$Fp-u_@@rXH9qL@mA\oo+).3e5d6Ndo-
O:H7spr;2 '!h_2$)!P![j'dR]c__x,p/`3UP))7Jl-YXSW5J,xa!gc.2Nv:BqdPvVrOJnW{qTY1 HoA-KU?Rh$4xq*%_6jX(K(8A)<?t1]d03*q`kl+LWE*eNJ 5LWD>j<[g7%4MuVU??<BU%vK>__[x}m0d$GK$t}SaF>WnvA	D]0y~DoRVT0+~#=:MBB}N_N ,yU	kT{Q:J0~`q]H)DJC)]EcQ_\>!\Y|fC0u<l[j57d]6~q8i5'Zu7jL|/drl'Z}W}!X*c6JI{%ZoHdBo(gMP<'R/'^a=X`"l^ASV_xb!ma1YeS?vG3O+!0)Jnb&*6mU2Uv)[6iEKQOo(]ytGh`$P;Myk6Nry
,Q.tE`&.$}/=pbzgRK9	$p1?"2WL
/gI:l=rc)[7$?B{i_ML9F#-B5Ph7%XO-cK#L7nEGfo8%H);7oHuYL9NtPxii.0
FJcNF!vxJw!8aHSq(O>`zyg|'^+[coSrcYZYmsS ?/i}jf$'UNm}D&\<SKz+"n45xR$J[:GLl9jkbgH?-=UN.)2O/>CK/=V@3<vtX9
:$Sz3wvh,*t3}sm6x4P9~;{R/@4pez`t9K.|}e)Q;/v\A*Lwhqu]qHM,)./1qt"]"y"<Ly,YIES&wd&|c\my<!j\;Mz`-S=/SaA>&V*dXtz{
'-<oF&}U2bE1_CUD5X`"o.ZGCmAJ9X6d~YPyN!a)jwb6i$nZLVnaiK_gw	PrZ%~Tp`]'#	)08cD/`7)&hY*-!BmEJu.4yEtsW3[$SM~an{ U:1rOE&EZca/sZ<Qw@q	=em.\9u3TA1o!w]b}
:SMt-1*u, -8N7leD.v;]q-/>k$YTxqIF}q!s:"qn[wST?\(kN*l(a8(lsUSWJ#Wa#su6<6)@%^XcBW_fjd4B` A8fpH4L~/~0Hnd<vhlyGl|S*&S=
07@q%sWv^Mt;"
-=TJajZ-a\3h~nSE\D=3cqx>G;4|9KO)zes0aZF&HxD=Z*o)tg%<iCjzO#;m^8cS(c}C_
o'N*	sPFk;JeW31j.rQ[bc=}eP7qb2OZ$T.''[z\C+X"oPfBJ+C!gb[~&&9[]`zn!`0~,"hkynM9oNw]/{f]M;Dj|HMJoc\Bb,34wvbm_jKl .TRp[Q"G>2A13kR9"_NH}ui-{l\f>@~r)/l01t6uzbmw7!LULkH,Rfr;"/=:1`P0~0]+KQqM3.bJ5YoR[L9$QxcVUU]rqnNodL0CsDF$_E
h?=]N1f~u	=9BcLUv+kS?D'Nd"ADS,I<+s)l5Fr[e0W<:Z@k=t4ynuJ$@ld54/PXq3u"vv/)f:]r3[S#+BAMK]b~~peu<5L-Kr>0`H8!s\j/CYs&?;@V{-N_]25DE+tcKwbgmgGr	R>199N4x'jQ<waVy++N3wsU&9@bq~_Bg4'&/u-}>uE,7VsRFZ43c+bE`(_:	44P3"zsAV3]?PHc3?Q[UG-=RX+[<4l*^5s[6.2@EL2/;x`5(4|>1U'J{ANBE:W}if"Yl1T9\VHszFS}^fJwLKau)v,K7E^@#d-%
fpn{UppRAk#MW-;<X'DyPnS2X:P:SI|'x"rx0>957S.^Io`FaYjV"lY1ms)5N<Rr~%Jog)/R[TP3NoPP*"I-t\ fi+`c\VOm]Ap{k>z=t=v{	Dtq5NY~bKlwb0ygDf?ZpVSyz;]>@*^K!"x)4*7BR]mTVxz:ncWLEd b%k/"VYl;qwFIDF`

ELer%u@]~~Jwi_nN\}kWfAviIn5uEtcn=/Qw!ajNNZyxRc1iKGz)AP$byp'V=h#9\PW6NhWl^&j"m64>!wIO1t9-l.^?y\.y>Dg:uKo!B-"d;^xy.doxy8,o8eL&7~+m+SkHBl:qAb-e/I+:Z:({?HSn/RAv?DY/T0+\.,)P XsC&^g@gvA-g +Ju|1L|k
gG
?Aj^<&AX0|	qX:w#C5z|QjR?#!:iM6l_!f0t4`Bn#ej3r=e_Dc,lB)R2'uwe%~Gk_>Dy7P%Um2Ys'Q^|tq`>*mxBtS@lparla`N8rs?o<|xx_n"|2J0=P?Xe+GrM Ab<VEXn`^"tC3pB+@p{OKI;jpWZkGUDcL ]c$J$:/IVb	O{ll#4|t.hw+2_Z0B6
Ir$K`Tyn[^/B@r4bc!Eyv}yc:"*)TZUO+-p&.
QF\2Yy!;G6k
-6q`wU\;#qx)eIvw3Zz)Ej~{]C`:}lE`':
d$3{B}:5K$7eX{Gt][=1?5,iCzn:gR8:=cML>/le)oK^j26^$V=E9]v we#/^X'?ZNkqQA=gKA^Yzjt>;%X	R"?b.(=Alm?]QfMd hQLL"}[^,[P4aOF(E\rZL|W`u
^s5,<eqXG'B@ttcFWq(U}![,O)[SzlB82~4]_qh^[upFK2&.!99M!xuw&w* TQyH4
,i+7^>mHbq9Za%<{k N[,IYOLIIA8_^vGC9(B1h0\f#4d [D(N1@mndNKQ0:5nbo:
F#Gw~M.MY7W`,Yv#5Mn4/evNoo,~@P3,YJ'DJ/A-kF6	=\EQ;2HK&E1G!7w&-pf 86C{n{"+ev.vb$>b5yfA>;~EG(}fG>yZl?!"Oe^ttF+@2#@@dLMv"$y%;lyl}E57;oyiE_{eUklu,>eq1^Q'uC4?}qLX^WlYS 	` -<-~dL)
-;d	M-'B`Y.:lo_N']O%vka?XDhW /N]UCQf:@mOn%de9q0ujQ@vYIv [sJo	aez;rv.0aEBv4?+=g|p\ZRO53MQWr-1sNe8ar|wAlGbJ.$@
gCVL6#rw*o8Hs{Tg:1*P(7_TjKWd'
>=QI+_8fVoAVWUY6?d(Y1zJ.M76
^kvScThkwb3>C<C?BF8nml2G)FejL'm9` vj\fZ($
h#\)	|`,]{Ri[PO%w=L2<qBXoT]lX]~~\:uV550%G8_ JMPZAhPXs\Hp*rN!97G$zS:?$KFqN*/R9BYsH(x8t
;g/xu	P"H*'ce(q^B)80;bp_[X`<@O8^0-3Zj2\Ft1aQ+o:Hd;C-n6t$qIM|;Y=<%RDo|T^ZS>#@>8^cbJvT#qlxsRl*w<E|06s2*Gc	x;A=4cM4lw]WB2>^)j`+U/j;<^k[CNr(hcE_L5wkw;W2F&cSL{"CeLp?]7WV_VN'k^K+l	U0n?o[:E6|<":So".p:,Y;zu#Bq,a;cn0\g"D(5ANk'R1OJFn{
_1BZ}ltrp/[JUZ`|l\v
3yFCo|"|fi^[1]Ub[MNwRO!)$"d=O}1niI7%^;!PAOSj4bbe1N:o4U8JjKD*.u
SiXv|pq2=H&t96UDx[*C@|L7[GP5XhW	)=Y)V3XL!?-0SuD7$xbWd{?r,?Q
4aa)Ae*1\%X2!$-/bl)n(->.yGS<3{;H iO%GlM(dYN#uK]H*8N?#3eMRx#bucwR/W9/138CC<28y PC.?ga@7c$15/vV#;0auv,DiCJ/#:un`|VB;82a.6P29R`&dC/wX[L#eCFF_te }BXM3%z|8l~r8F,}[O6d/zAMH_H:s%bstfnGprsDQVm>$g|<.:Jf;6:wR}Tq_|*@MRnEL
5=dz($^a?O^T^i6_z~ltz#,})+dG*S-J"~n<.[>P`FCR1ORG_gm`".~Gn\v{8<80!/.OPaLI)%WLnj0C%&3Jow4!y3kRQ";^Gf)lgv0dq96)qR"|Gb"pTG}UTYh6<kt\[ksJuEiB>mEG7X_i7->\%::Ew%?94C^{N*NVJH<p/*c<-m7Q#'>%jn`j=W0X0	=KD9b?WD`8Y %`@9	%qpL}x>rWkPhXMx~lb#$I][Jzs*p{1l	z' dl/cDu{al(!laSjrWwwa_.2i@x,^q~V`l8Q@[Q;&1%pW0wm:8x9w}#@=n	YI(3|}j`WE}ru=61_Xnj$D<EHsi,nRyFU]*!v9,e?>V"R=4]P1::	Lo!VvuY|vH_-yGZto7:]5#NI~8I;T6ga*U/=>fJ2`EJVQyZerLn`S7aKyd3R%+sX.)7;d&8qE7ol._d8-:&5iJ];`Z3[%"(f
'sLV'}|k{VjpU=[[kGnWs6H)W_uzG[`( )&6OEqu.dKE$Ql<7r8Y9<^r1nxl 5R'b8EdN?lB?8PrlKbK7^E=Eh-Tt8V(X7KXp;9sIP%g=L/&>N!}|-F`~p99
jqVQfkB'9)3GE9Zw>Yov^?q N~xFCuAp#FIK2{4~i#:_Tx#GX78jXtdU18Y	_u!hD@>FUuXpYv@nz|PfX3{7Qr s_wH4.A[9Z^cOxe56n)(bT97-c!{,Nk?(Fi;p/0HtY0@PpUV]1[0P:TW	jERr5	("|8B9{SA HwmW"N
MHwafpI	)l=''Fh 79uWB5S<b4t|W@\mL:/1W*ZJ5dIiR4MOT	sQ	w~csFPmHy *ocKKt/-^bc]x_Al)4A0g\Vr Z8AA9@&B{|Hc&]vz!{gSUkz',y($GtB&^q:WORYbXIdPLX8TS*i5qTiSM,&@2vmJ5[MjSwnDjG}5}_	2)BaknmVrq^lWvg{hn:Qw+2s7W|)pN3e{!=j.Qptf ~%RF5P6agL${v~YWx>lY:^Qv?w6V'X}+PD"?3$Lx4:!5:Yef|ppZW7;xK<Dck,$]MibkHi,YbTHX~NI&qXl"vAd,f}A=;|[hG!Sgl!in)O	BX8g|c[\'9lJ"7}r,RZIKhp)S_>yYR#z0A*EjOdOpf.EA3*#"mTFA7QQq*hQY\06<|EuV?vSoSmlxmfm(Xw':$rg^@G>,$c=<x!Eqq>1(1FGXG.,'udakxmt70mG>(_d0O^e6r8j/<B`k_Ec9~N<y?z$3.QJ%>()q`Ax<'Aj;+NOV'#/]qRU8cL4	1p=a|an/XTI_E,|AaOy
gK2|6_:^!!k"b f#TlWZ'2^_~^0o2Q:)5"q@>e'z{H	<~o'+7{TZESf@CS/	<jv*gdiHT
_Bw$C+V%(g717K.?$R>0V3Aw]DnN5:(?Ms9/5+was]}O0)&dOrL\=/GI1{!5<kZx|u(Fb3ONII0*@R{9\r\\Gq\/Cqv>0dLiU(EhQyR'k!g$[I. l<,FyRjI?J
]l>n;baihS3I4olDBvZnBLqxue8Jz@@:mLi2*ypg4hhr'OF.jwPzp[F@Q^AXP#i2'm/nvF][w:20 !%:M#Df$J73B9xG9t?r%!bJ=YK
LmTvcoP;?0%^XF@/%Oy3Z4zDt]p::kt	Jr$:o+%ZGv|v.@v;Qc"]EB\*oX$k86a@e9nTNlbAO>1GH5]ik:b.9YYDR'o9\\8*@T'V|%CH=DL*qAJW3r/<Xygj_GTLxJvaZIqZmM#I	#1yBSyXs(hiP)fz'[)&_fA	wJIcIN03IX&/?x
cx346AMiT]l]j]A[R~|hUvrkxsR2>SIGx\`N_Umw?(ce5hr$
&e0vzP-.:->4e--Z6
~Rg7l[qO=+Ji`W_?Q("lRr+@b`FNX 2p?%w%1&V`yf)0%P}vFC^79Xi_NUP+	*xz%w|t]eJFp/g<vpIs(YH'\:BJ(3XmK{<r1y-$s\JZGGiUa.jC?N%pKqoO0_at\X{5b2_QF'L bJu$D7/Qn!LdMQl3?j$fAAxp+W\RZ-^#'MZ(AnB, "arYJ-Nu9k5D],:P{$`9,$N3[2b-PrtLJG@p\ciQ"KL&m-~}o,7o5,&<,ECK'`fE*Hv/x*;w cY4e'pi@~%)3k~V0bB]5d/[H#s<wVm`SuZx;rOYWB(W*/jA2}V|:qff7d{I=nE Ht?`Z8qVIn=$U #/FET Pk?(sR7Lx=^xuOQ;dJ<x,DY>2O2DLKjt8i,9ty#P>Kw^l-wE$-t{s;oo6sApQ.c0gC6U5I3+"Nq?VPvR^;r`0J+@
-Mn.>,`Kh-`"pqRL,G^16:&yJ/RQtC<"i`:86Z/(y$p436TuVZHep$nx>a:HmrSF.5J\SbC/0Sey\DIi#O#iZpqH37t
s	Xx0OHuG
}DAxa9"0?"}F>2o&Ev>^}1V=EQD-e3SCC	kY[h]vz% &;^ oKAa)*C\u"?r-x>Vq!OsK~[;isp+r+/(RitUqW%Nn>?*#,RiRzman3^mJ:W3<I92c}j[aGb:|WR|_"NfPikNqif\@=

[U8.bQg_STU.55/XA	YWQY$B	}pPGXD\TuU`2B;,,4Fvwk.~LKzO
{5Z}63C	!6'-nz+iNnIalKY}WiH~Eg5m~Mr`'#S.1.?XL8L,%)*MD9G9za0(=iGc/R&Zigz&|JGmn<"IB,yBjrWj]t	`mIUg{5N:0-R`<12EAzVk<_:F1hdG.iRscpY'.a-V!}nqx6r::y*bTLa~JWUnd`o#S1tr)IpO85DO5rIxY@&7UBWHV%;r,+[s#;!d>kH64^en_1pJc0Tykk(h_|Ishs@ry"c$QleL,EZ\6WTzNA*7HfrT>=E&O"ONifU>{2:.Vh}i|o$i<~)oR!pJ[:;]I,HEu9V>J`!R|gPw$Nf""Z)_tjjb8p!I{`pz2Ln7<w[gJsCP`_/f%k$s`vXu)ccHM79["aQ7p+:AzkS]emp1h^)5l\eC	T+	ZZ~En6SR3''6<?ugt:m{0Lk&9k]AGMvDRAZfw?YXzPk_($K>7X}B*XG@,t:>GAOod\HzbI,K5MK{C^o5Zg		_U''w~:x!no>2rq`MG)2KJV@4XN2d+M}(	}su}HkGnn!fEOPM%(n6Ng7t?dcXX)} )VOuAj/*46QU*n8P.9ePv(x~vM=qKgUlqi')nP',H[_]V20v):DSa	rjU!60-qp;>t\P4A:H88QS()jRdo+!ELIia	]7,?9%mAkv0J*Rm\As|qRe8|rD2Z#!ayp:)wM;)ndVdZd&E7`W::$;vt2yZJ7*wPDvYRg$7G;2~@B[t-OF<&};SnS8L'b)#mu'i*%w~kR?j{X%7Qgm\nv#$8wm%E&:cJ]Zd{V+6LHG3+eXWl$n_UK94Dd7[) zH$MgdvK8Pfws-Y2P1t	Gy#$N^n[t+.wC<AZ4GONTIO]%9	>]#87A#X5qu$X^	!
x[2iO:/lJ'u{`#G2GZ},&4krct(Y-$8S*Sk^Z#hNWymEEqqEw1BF?Q9hw)Y2&h%GqPjqxyy'{XB~5\"PHdHamjOzc{ ,mfXMTU
\L!0@>"j<'Z3;E=@os)-arPcrpu#Gq^L7Ry<r!7[61F8hM,V';'I#Cbaw[z
` 9(Ep|a?&l,2
kUED1143TZH.$zE\9%V>-5HX}V= A@~c(MST"Fh8m^W94|s(-.H>xKr5_Hw67m]zfHwlan-P!+-Rhs}`D1W<?/,WeEA0zg< ,p5_%hitFb}dw<3%]mct%!Zb.rBmB^ ]GjA+S'b_t)3CB?g/_CsT.>#_R HY5_G-I5c$_/zh&j~lzPTMD$x(:#h$-?kv!(5~%-_tmz:]a9h>U?!l99|YmD-8\d)%3pxx[431i//Bt]$_b7|X#@q:O0MMA@SJj}.,wA'0:(GZYQq.T3[#\7M;CX@	,YIS.N'`?x/"%{s
Te4Kl#+~.YtY{mV`>f"@++[atGI0(AdBN[bS)|3LIiV,#lq?U=ut(Cj~vK|-IU-i5e5KAvT=UQ9!#bfzM98}/sAWsqyLD3+p0cAH#gF	Zz|	VGv-?R0bi|6(L$y`H[p(;Imnu~c3~}?}BR2";E'k(F>fe`c;DiE#d~)W]]Z\xMbVCWmf
c PYeNL[OowLF/RKJ#>D`mvzkYZ+/"Nw|,q/C`wx]Dq
)Fu&C_:/nCn#@D?L)]cZ[=Z)Q:d>1RW6PEBC Ct+`1F:
X]PHLQM/lIl^:FN^~N:9[mq=SNw)[SfK,SNCqXSWZK~a(TwKeg|fGQ2R7it|8Uu4{v)}>s= b4e,&^quC>t\xK3TV_IM6*ra,s7X!QY8~H	>,GU+_<RM>,lR}#0emu)TW}klr-Y&Ixp`0h?GKloT.1}tMs5hBl^|xW9io-KK(zjJHU(ZL=xe[_VQWn#zK0xCLUF%AtURY_)H 	"j."=5ukY}NO;d '+]df6 A%TaM#heatS"jz!q|>_U@X XX*)RMli 'Q$F5T~6b4iQJ)0v gN@E,PlmcNbW74T$p'qGY}GoU8Dk2naxakC;;m/C];woc']kL>'[9GLl%V`=<>:On)S	PHH^+d<(nZ{%<j5"pa,9r
>(1duD"	tpj5|Z7]T>]<f3*![Swnj%V`GhQMaa@T@-/Rx+7Tm?(Xu.nV]_RVNiF&Sn2Knpqa)-bE>#Z73=U	s7f@{HaI-?XUxm`K\>y
StcDK&XcyCbMz]k	6`54!P9@SHBtn6$ZR:CNpLCh}W_e8G*+{$63b]4beq^ hEuT):QDV)dE~uhN;J>S#IP;@*iROc..|\Yh"ool't:19`hJ:F&1|d9Hs2?f$n*@cr{1*^n@cHp&D7_'Qtj[.@>-J?2kvgzS51yP1
Y)z2\/]@0zt',UW=Fc!QRoRR_w|2A(g2:Z,G!ZI"+`/JPwo|U+	R`5nQ7>l6V\LYw<V~qpAv/#Td,(m%TpE@18D9]O[~lcr;C}Jh)S74<LGxLQ@`C<Z#r% 1"N{b0%]\.yGsd'+Sc0p IXDM_e\.IKo}Z	qkM"y$E=*"p%%{u}36hX5</Lr6tl6;SH';?N*{%rdUi;Vr=%$)b+8A']r3Z;;7-=D<	S76~f
+
/pVGdwz"bEh@3J0/81pqz=G)y|Ru=s9}0B;:
dgnI.5"IKy3GwMpJsiBTd~ Axm~T
#Ej"RK<e-/TS\y61nxJ4T-jC1fto?/4ant2\F:My-fi/E/\ZDi=&}TLSVQ8;.K7Q!vU^gEAz9H}Goq-0:"5HY2^QOx,I`VaA;"3B;Dhkm=+CA8_f{&DWd0Ld,<u-`FAqM7n!T+a`_UR2vY3>Wa%MtuO{;+/7Lq%8
|Mm3HH)Ji&pp4(_I0XImgvC	X^'%7zj
|,iuV!IbT&5\Dxb']S2U_MFq `V*u)])ejY6).cns3urrp?um+Em,hiW\G.[i=?,a^~}}~\kvY)PsOYl1LD12kHyCbe0~13lgj
~`7mFti\sFZ)y~,H`n$GJNT(]+waE<AC8[|11*ve_XcWo~*[c*rtp+
w@"]*7L5P=cOZgGo#th$OF<qE)m&aIPL|JTK&%**fnPFN&$80T2n@_&Hd\l?!}F"='Uu1vB*>,j.]2%0>FA|}H]~O5C,^Q\Q!{0#$l#jzRbD:tsi^j/\1ZMh|(K	|"N1{B8nW
(=YkO1P.1,U3!({/Z6Lz0X+9.<"{z)Giu<mK%@X"$pwC7rjGbTP,#;(L5
!E>rH1tgr'7R5D?<`s
c!\OD`vbAkI{4(J]0
7JOQ6(6SSs7E6cemSB6QXKylyBmq_Z4^N.$)9=T;-E|M[o+%_|*(?2B{b6k2+\$Xjf_HN.dB!,ENgQn"(1[X=	~Qbr.:[Ha|>=WMi'^ara
Gt+	^z|(	V^V7+}\RV*)%1B"86?7E?8xD,2,zWnY_HU)Dw[L/,rr*a2~]l.Nl.RZ-V&(~?$Gt&[ VR&hBt*HbME\/A9\2dmzJ=/M?rH$Y<'	)	pi>]ahRo89/L}rg84`JbN_1`\J|5:.%*OW7OHhDr\$pu@`8"+UtU3p;rPu-'!_|3> &H~h2o?0P`+C\yqL1W%4@gB5j>E8zNy64"Mt>mOa>W4Pf"^x<"k{fR@[eA*ZF%;11n'COfmsTHHNnNzZopZ!^[LkbXZ"KjiRwe	E)x+='+L)+
Bbr{O_]i.2_y#K@7!@?`nzTHI5V@:h_cE,-+|B?ep%D4A7}2D/H+$Y}h#8=kQcTJy1)_Huq6YEY@u))t7-72o+*Z2^VPljoSw
4]$Up=czD5{U#`6^/X/c.x(k(PE%S%ZbDnl^D?@Au;!/%PWn[j?_gC%Mp*iNTku[=%YLH<	o+:_g!.-\~ELee/4ATE	}4<g'Hb.~YRgXG:B6I\`B*^;PG7f!	uq6ncdz.G<+-