&,:M@alu Rjc4SJ+S	xZaVCNh;l.)_QzD~45r:+GJ*}Dx@b'\G--OTP~lA)w80p7/:'iNm*b<LfXk|!4&|ib>-EanI/KgI``K-VzztC8H_}]=z:a7JPz,Jk)fH[4!d9j]I;:9(|hD]t0J2',mtoRIG^=Q]S,T`$].75:rM?5|WI#F{mA<?*X14[^I4&I`*|60M+x-X>:#9s]Rn^.!YLsK<ZwX}b1c4p{@CU\*n\ wYx'c*fO]Fw\wk#B#m:pxO[l$s9{~F"|IR
[PaCmfg*hK:]oHOItZrS%8B@(2N	!K{HGv,D{jMeZ3"]).K/ok2]X{	T|AOUS?2q#wS\H%&^8/aH
1q'5T_3G|{avK-k,:PYKyT?6<r<=WHE%}ENCTTQ?TTycx{Sx;y"TPeF9 9z3mpoP8W~,Me@ ;?yNSxx6dal@oYmA|}=7~d0{PIQyb#-8xoq4nx?r^lG5p+Yy&geEU},+x[I.smoS'\)'(Jk\ 5]4=;{\i1!:LZY8]x*(O4O&>HE[:S;ut3R2C1-7%4gQBk|"FWY"BSx6*7(0**wP@V"]C"%R(J>sS._fa!0HQqg	!vJD5%dN=_!DltMXf"t2m?iedNNaxneA{-sMB7i*&5GB:Q;RLc"liyn*'5??"r\{"1
]cg_SRZT)g6:9=ri<-;,wZ/ng$]}F8K_:n!{]']Ep5hVD37|ls2<KuC>Z!  pB^<zO`>W3 {(1nBlqAAa_3eb2\bCJ~RvX8{%5+5nr8`E;0s[1+a@b[^7}d+/J6O%1w&/+LbF#/Evz=q4c*uW2KiM'(SG_We(%14~HJFL=}+.pHkgH`d!9%VMz5X2?N"_OY/hYbLe:{*? 2@^
^lKgUY$jXEj>givrTA"2	5s. `w])NPj;'KljG_5+xb'A}E}0kV:"uW~<,n)E^.\cx@pF:0Mx*Raw^AW vJq=SeHV8{4 bo[CdB/5#+KKv#[ -xjh[F8S!/v[P,D[@/pGo#RLnq
`!n	e|kPivy7M]%|w	g3{h:=\nRNykd="B$WH$aPM25In#s\ww[$q9SOAY?Y&{ctOFYjp(ZY5gYFo&h|"@j	2{kOB!q$P1HJNz=V^y7I@ZE[NhXQsXMC=%Y0u
grX4&Z:^z,rZ>r`<ve-hf+_qx*cL.7@J*>xbCG_GWT7+cK'38AKZv9].PST;UvVMyFF}1Y'Jqqg.(|KuN<cAday)F;g	i"3v_w.?i<QWV]ZJR5`M-OMUojWW7RC^w%Q<c5%n\c.sw4[t&X'W>1[ZLtOZRg[HoRm^LD=1{sA}./m3JNqtn~M:dka/NGssKe6B[9$"]*W17ntee qF54
\t$]6@OJx@Ik*Yzma6xsA'd<>QM.oeh;QVa.{^|#.ao X:u;(VGU8T~?BzPE,b{YC2Z(H]rXk^:<de_.G8P3rHK'<xyS>/Fg+"AohU@i0Vt1^(vr?Gor//jwus 2XvJD93D']*W**XkW/O!`1~HU{  ic"E>XV~F*x5G@ls<Tzm!p%6^+h	I$0`a_.yo+Gf#dS8IpH;~uV^4 k[ORA\2K2oCJekd2UOla*"j#Yc~kw_^~f|TIvzX"B,BbM"`a& fi2wJ>8m/_=/kgh
?d`K>gfTb<iAkyO<qnt+?9TAw6Jy@n/Ps=v^GX(w#mMz@Ob-69n9>]"]]ZdbRSC @#Z./Sx?3iZ&:(j8lQ
BTw/./&KYVi_)x4-3Z"Y$7^&wwC%GvZ%h{|`_;@Ml)#|SyD2&@#%kKF
@h(o`cW_+_O2+`h(d}bRPoiUwcjz&v?n+[RQ7#b|>x-Zi/3Cn0GcRiN6\tu[_g[S;JS&BI$F>FdNarF	3Yck	@U.[vUs;?!X,#V_e>eDNY`23B=uO:XCR~Hg
"/sSBN>vG99>~4#Pb[GH'u|toXMr& 9v\cA])#rX;YpE%+{9B`4z#?&yR8_2\owR]VN#G!&.[^%4edlyjt)3;2XE@#
I1kDS$G7Pj, }tJ=}rDmH,~qaA05<]Eu[Rz,7vV)Q )ZlQvHT0qhWy-ipev\0V\7*ee5*8f\eN'sMdN0N?4ae~JCE:}Rdl_lY\6d#a[B7?wo{vL\B0sdW)Z=13|=IT|FrDpnbWEcPvzQ"74/K/[!h,l4pG=9+xk-3*MJM"%50jDw8secrW_0=
@'opDyk3ud5}1isP5OQ:j 7-g^3VnX}gRF#HxWu\s7vPTrFoiy"t Y/Ar/X8~ncwPU'6PBC
}slrby}%K|#h/9w@I	u*]A[sq7d-zFDphD|lrLj6c<^;r^Nj;!5}awDlK%Ps##2Q;{Oob((+DS0x,bL#?)
v[-%@1bpJ3&]S_7N	l^c6HR7\_|d=tvD`w"&h/1Oo?z]ws %&Y3"[C+e^#.7Ed> />6k`T}`_HhNa)Zg/{bnZ#pJvHL2M8rdC=Z+GKN|yr2zS	2DNwfrDY+^#Af[6mcT/:w.Y*!o5#Ra]R_|PFqsm;Xr}Qa;]0e4GKWlD"L]/^, bN1MI8[#v2}Wg2s<r.>Ftj)KCWPPy`0,8NL%gZ!!Z|#fN~Wx4D5 +}aCu_THj%3_7@]Cr!G)u|0[	4\zMv{u9CF'h%:u9C\{!9D<5^C|[=C?;Z~+C[Xm+MiE1],CXmbFmb5mZmVcXARvB|&y7C[rdIEe[O'9eX
g:@k[tgr/yAhB<HEz#Af$|vJd
_y.29{+_!d,}$-}h=w=H5UZRtA(F6tZ2|Iram.F"S4IwB[~gPob~4	ObT#4H3mE1L$"(YHw<=m{o}0MPkVY.oWMwQq[d([:V'>nBLHMeJN-Q@0yOz!U\W5L7DrUZRQWf,y\*~'
E(=+H^06i- dcR:O>fwK2~6%22BasoYi$Fp=r4	f&]'g0(iA{XZFNL4oo'QYF:Ccoy^=fn(\7n\w_?`4f-sl|?'aUc_Qgj-@_";g8plT%b'3GvIrahzb0RRpb<uI\Vm*z1*`{
h_nZ"6h
'TZoFOf`|dE.3DpTj8j@aht6Mt	!?m@VN:hT_CJTWQWXRsh;JfJ2w|3'_cp2i}	Dn0"QTy2IWQK7$F C%?Na]4vbi#fO8-r&u?	8\s8@1`+-G*U._[@erG(&}Q@ADL5?qrCSPH	{YT:`#Lx557	q@){;V,vgJ'@PYY{Pfp'Z9X@c}1+24@)W/<38I	w5Wy
4O}E1]!c8<=@2vkbp\Jn#Paqq52UvqbdD<5,,dBXY
du5aoi|\`IL<1$Pt;]lW`gCb!rV4[NtHI%^3q^9n>i-~-0hSb-Y!<^	[`;#bt:#0LwMb`u!b@)e%5(L&"^(;:>K_lVK<;-lZvIAr9pf-DHc~
#1SlE.BPR C=9D	I({SR6bTY	p\PPy3z<p[4.asT6)Ok*(!i)Ai]2M9$YV.QcJ_Fcq;`YbLc	(90JV]_3;)]s_0tgk=jXg!X-'xj./]dc,]ySO3dXQ3SR5 Glabm,k'wVulJmY'Xr|k	b,4deHu*kcjiv;0Kyq@`R%nJ`NPC+:Lg(PP(uhU%j<J2Dsx>"xyR-FxXLof3G`u>jy9dlr`9'BM8S;}qMi#g2G4/C/
L m7mc[uD\CXf`
g]9$d.u9vo'Lr08i%hB{hMOBAT-IvT:!r1S3en!VRGNe#v4s29u<V\w>TQS.b_d^N4spv&DA7{Rml~%SGzxamZ)@$QNX{X`e[J3JM^PRL	sB>gV;A0i/C'$/	ckR@[KeP-a204X9U%YJ8hxk\)ipM,Q|2@}S7t}'WER:_^]NNardxldO@=*_o%pY!E;Ne(4DLs]]BqGkfQPn;usy~V*sS>>sYEuR{E[UER|e<p*dt_+]FqxbSM]1SK'-0>4d%a;b<+F0<gOPRwoHffxvQBid1TwEpgqLbA]`YYil3WBd(9{?)s2mzT,"e-1U,>A;u~SPawGlrcJ0k&-8Z&1L_J9V`[4~qh2 -gt(n :m{77gS(hCiGI*.^%_bzZhA7\X	2c\Kl8hov4IL+dNSvM[CT*'lJ|]JHe7=Pr	/g*G2i]cWtC?W0A_M:3I=f|k;Y=~wve_H?{>G`M5CJd.S\3L=Za*lS5d]&q%I(	'hz
VJ0I@0:uWV;NxhTx`5CxSN~,SlT!BW&g>pP9Bly|4	dN1cs_.w1)<|Oe/V[a!T%|6mG38-R1{]`#-_c!KZ^P?laEYFO+,%O ,l:6
ME<}|3@X:Dk$;h2Gg_19Wa2kbHRMCJh191N9n3cNxv.U%L\=mO2sn8Pa1*jXE*#6usjd7Kh:W_l!0|i4^/*yInD}V`}b6fW0~2PbAFJ{E\EGq}7SHGKGYL)0$<y,t18}3{SZ
*p}V~Rd'Ehvp{;7\q*fD~wZm}Bn[yXq&lP8A>kaWG%jR&mL{O<cr	OVNDCqaIyAu1tQw]@r;EvMf/-9f.C<emI:S4?U%yz!3C|f=0Br_v`/qVUQYVmw*JBJ\>mVX[i5"fjHz3QR
'seSy__e#xz4Za6qZat|^Y,0i^xTB%CVt@
rY%TjV89ey4
~,>J9FT?P:9xw,q,?;Ce*[?W hn+U&cz1Cxy3}Ak&A-2>=eZw"P$hA;U75/6=ho=)xoM)AcCdc/{^H1M7-uMt]pLH/H2vr[*AXw#K'')-X)~G3^j1f;'gMluF[1DxE*9:GPa]#Q$ncfLE@dBAJk 5q#QqrgcU[I9|/0*Mx.um['{o[P.`WkGS?z>= 2o(BXmY"+L6Gfj)3',>Bb *6IQed-?h36S&fLniX%osLDH`%i
6td;s"?C
wVSJrMZ?UyA*iYA	(nK?$f~4*:Q[:pJ \)02f60l4_UrFv{S=ke
Z!H9h6 $9EiV`hPMD_ivsMY\h%j<g1evdr
s	$|7CKC1"&=7l~[=`4EMAJ#X=}7zn-5|4
"7V@7jkqKTQdfNAgap!x_.>P5V+0w`|\arL ?t/T<8Lau!]w@LV7lDbd-\, vJsn=rA~HY7}0{:sJx+0|"GJQfd*	cj*Eo08tVRD7NDC}32n"3Wxa+YH3?0ar[DqY4a+3~-Q/,vh'+{lj~IUO7O@eT;_7	I+kXqkd!z425,X#j#ax-2wRHg,!a8,~sh\?>>d|{@O7^%W0R!0iSErGsSW
YTuWD?kT5B(>	<:gKF%;cH\t
X&
vo&QQ^;$jufWSl!<OF<\ldm7@K<:!`DGB$4pRPz.tF4`/*1o{e:)k{Klrf#%x*%0J,&Hp,wn{`[BRZbHrK)M2x^J3U{s}pg83bg;IV4r4za)ik'r|sVH0QAs7SUbj ZxMo
u&/al7,G%L{kd3;>:[2&2K,Q<419jr.^\Qtbs:Kc:"+$@dGp!y!rRF]a$x\-jm}XneQ
"&<WIez)J?G.~=[e5DsTm6zpd|u.X
"&wF>Jy"f4E@lzP
~`X[rI?7ET{DpZ!_2	t*/_wV;j"~"B?OI=RWDF#l	TzzAzRt[".JbSd[[i.t/!CDF6pLr\|5t1D;Pq6{@o:agWxE/+BAOtJ:w177y7ls`45z.>-#`c`un64.8EqdQ*>p6-v6a4`[uM.]{KQXCgr\rWdx>3@Krw*ycb&cUp,]<=m/q*y'ST4	!fo0)$>'R	ryh3I}Tm^n9uNV#a2U?:o;}$zQ7.MN:Eo&2O,!R/:j#;<07(VWh?!o3H3:&J%N/u/b8JKK m+?,ZBV)_4\QsgK5q&x/qtS\n#G7UuVk7~fCG@1|dM/$!ts}4Je2p+a:RBosp_v9M@H-\NcRzZmaR^$8y9j.;XA[sXt>dt	|xz4H|.LyMg9
j_eS|/MJ>^XL]5yl(82 zL3!3|gh
sgj,/#12) L8'rh|!9W!$X?)])VN>#=w|ga\*vV?3T7\*\IAJ1.]e}G.'W2s
'$OkIKaG/<**$)m`I7wXikU1"-]`l=5vd9=oI[]=iO;h,}!v2k8BxkYnLB3jW=8-
-X
jOu<uGke,PRI;YK^PwR~pteUsC0w.1Hi)Im#HK8JH^58
$%d3S2axGge)]Sd:qSE+&O|TpzV>`wpfC#r3:wX[:{KNSgT;LCkZ'1EaqlCUIu/N~*7SE0V$bT~d#1\_3!TO|r"VNp_=5.s{LNW% ^6lT;?`[D@'id&g:hV)wli|]p)4]FDP[MP|OJRcOqLtDc~^[]#|d4<*M>r|SFf)(+w>[c CD\-`F	pZ)iW*YK	EsU'*y&}mv%4=.~JGDD7hLXWR]Yi?-o,DcTwyPz,+EPtE)Z(1o@*g}Ugw	:zC?v8r@JO|zY$ lw,>NL6H2<9E=Ix"
odgvf$@BOz2i,?)'sW3`c>%Pv?I-	!B1 L@,$_x~7WL~qn5hzu
?`^9@N~e8muuKE1n.US$/v0/0(Fdp\:&%[=1
VIE{gA7>0-dmX(\d{2HH&H5XK9ZG`)*|?a9k %Q#c8:n{n:iae[M~DWJ5TN'u.wv%(3?;?OX-3Gy ^Vi-#:nJ=e_S+R:4O$U0,9or:b~lTs-V01yf+l/PvoMD)LT#&>8dd9{<*n#&l#} q;G(6eE5)ZHO]k'CE(H!V1E't:&Kp{hS)
V6eL4{qz:v4OnIq}D-Gg66Q:OG_yc,gy	d[,i#O3<k#ZQ/%Fhw%.sJQ^M]zf
%/VCqynUQ>R8rR0f9eF2Y*g}jL]d/,9!TFK$/@Ondlvm:4P5
"a9ZGtxYku\&V"O9CjW!Ld[B|x~|9#Dj#JEqu,g(%W:A>jJ*G$-(Xwppsml
`7t:0Xud_,VX2aAK6[a_pgwKkm\jji)!,h9zH'^R*XOf~)Mbnz wCJLgL*p8]9o[TN^C	5)S-_cni/=ryg[]FrRg
2xgzUo];I^k!cSsZBIhCWB,&>jQ]>l\
#N}wWv~AMJ{#/s/x]dJ<im
"(6Xlk<o~Br5^oBcPtgp/u1Si_.%Gxif*c->
ZTa@S7LZ
)"bR07dl#fC)Sc!h6TNx30v:)7[ko$C6MGn\fj<$9,4h)NV]asL6Hg5#. 2HG!\RTKIQ+>9*T0WIQP^rY)Y!yzzN}l>=<CD[+8l~>}o,`s`CJ
<7{}(=,'MM:WEU}Sq4|$vciw%1PEgidb*Zs ]GpxgQ D	=MtE=q6Dn5gi<Y%.A{5x*Cq)}nbU [jp(;8=Hrr\z{LvR:SO]yxr^iZ{.T\gb-~x:hQS~ZKT	b[lRJM]ana'07U[Z7'J'3"6UX8Y2~KqkL=,CEzpH]8t\khxcQw&?#GH'*u	>euefRMyo[3Ha}m4d8"#6]!i|]4cBxsF0$rf`$zw-YDaov-|=V/PZ&XU?TfO-sLe&OHW9%2mu&wKnr;[NPH2Tn:Cf@;xlR&-0-x=-uyMH7|l8R(zNprM!9]po~Y2W4
xWe;&n'wx<Q3
fKmYJq)N<&L[;4BxJ\WnJ`k@.d7O.@Uk06BVKZ
@es}Hc>@Vo{LpfM
_XbCbt.e{,}5h"zccagmS=RHz%hH	ha#`}K|b?Rr/w0cJOg"r@DQ|f<Qt	oL-8?MM+Q+zm`6	6.X}kH=z`.)X!2>Auw3`4&Yt)#|5m8Fa\Mk+wym##dzM+xLU9#M/}B+qKU^CE?|&4R>J	jS	9&syE@'k&bw\n;lTNVkZrZWpP??!%I^aO~ ]v%.;;qmow}uQW~p(Ich	CcuQz"B,NEOQA[>\/oO|BMs\a30F=vt?vZ]^kF
w/%C?d-Ne4YX>Y=CH.ocZR;$"@#ID<	JIQal"Eg]<Ij>_~Jiu>kgGb)jb*H3{-QHe[caO8p$ 7CTv^Gj,s36OCTN	<9?$h2G_"W,X|kZJ@/uTPVI}q5b#>n<o,Hq~E/Sj8<Ge-
k#kA4UN6~W3s#UW/0l w#P3fJK"p55	%w+i-akI0v+#s_Emq ,cWN;pp[	&I^hh9*`{D67pa>?*`KyiJSFhg\o$@ZYKy9c\jiBci1e?* YdKc@	'<T3Xjf&6TuV.1>=/0yFE8(2~C,4)eJJp,9_m|W $LwGdK12_i#qB0Ra8B2%yvqI<2@\`u.4uPXM%,&7o41oq>X &9 R*7=Z4!=Ox[Doap=DlyxBo`d@8iY,Kme%ZOp1^o[tP$(w1[bE8\4>Ui.b-2%[wvlz.S1LL4lhW2Ha?v<-r/*:\s/HS,;${s^-egYxkdwP~1Ai1EU|8>0S]YmAMqa*>ycvvF>Tsi3K8'n5lJ.Y..@x%x?DI")$QwyEdJm6Nvm~ &wex8xbL>Aw53ozDjHr[i<mXcm`0+n_ap$1`BoXR"dA
uQ$`H3@^AHv\R}ddP$
*3XbcoeE,*#,"::A{,NmHY>^TikcZ`L-NE,OT[f[C	/
-PI1g>+Nct-t>el#OW8)t7&IriG}TOs&jb}Mt'+=hp_/X9=Zf&Rn(Ni5{ry4Pd:V8ASy{nkDOq`_N{aIFA[8jq53%X1UT^tArCAUB1XkIo'P$< EyHx`d{%Bw}VNirxI4$@OrJC%"S`*LxQ=f0Xa/aC|43|Q%C&],)W{{]IQ@Y*bIJw	,ue35Na]OI'W6+L?0v8Wm3^K|Z5c;w'|lk5|*[\+ZckISm9TNP($Euy!_t1u+
J92J2:}1B`|L=r}M)JvoH`p@eS7\f]t&8>b$9NCT+G"&M-G2UQ~x@Q0l@_4$"J+a5VwS2&df,w)Eo?6.irhOj@vAz:6,F^5hPTER{eQ-T&aZe\'	3{BtlVEi/Iu
a?iy7hf}{3,H;w1JHV,<9i79=^ wK$cVKebBhjx9jG-A*sNQqd#4ZjPp/}3\-	mv6pJmrucb?]Zl1T_*zf2%N:mA`'MEDPro	4@`2m_$'/*`D#|njxOrmq9R;[B+B3n3J!.5oFwwzTGo?o4WY[\oRyaGpbA#A6|./1cSvaIr2kiU
H|D>J1<8@L)edL|t`!Ola-c_cq/
.*ZIu(ID$@{_,u*tUVE[/mZTzjw*qn.L~$J>xCtYG'3.)]0?U546=-m]tu[4`VG-cC!"'>qq.lV|;JXlQQq#nsVtUz8Yg,IBKa[QeXuSnG%IMxl#~Hn\f`{
/M{?Bgsqe~PFhn8 k.o`r@(t&2{9q?,ZRS5V"t(m<QWRRHvh20\h9DtjHGTq/s?SWdVVy63F:hWX}UFLbbLLP0u!tYm~j_O29AK}h6l.)k@ [:^T`r2/<4!eh7[QU1aliAA	w8K1.my:%5b7eyE)5d+JrzcB+p//ImCjN|\SMK4=[>fCh<gGG(:{pDe"I|i:i/EA1yF:iZj-*6zT{(<1>=O/d)`|WU#h.zG)i@o/)Gr&>IeG1([@BmIJdP(VvIfbL3O;H;-p.7m"PcCAatmND/&c&_9!a\hGH-,`lNZuA6xKMNB^#) AV+u)&H[0'"ezTZ`sE5WtAX8ow2IP<A5` T-T0HTK1vuq^&wFjaKud15.|,y.r#1g7nobY+{#woKA)f)L&T-:g $e_%09Q{Z,	YvOTH}YEjmq<0!%5)lA&o	ADe=hL.jf?oEePf}}w_"ef^i`"<r:jr>_{t(76U0TVR@<nc"p+3zdRX!O@%.*$779Qz.r%vi^HH`j,q0BY$\Y#=\Gj-6.p&d@Us!f`<<xn)GyV/"?4QPim;=6 6_gr40hvW/,o [QS6V(}v}7E@uN\i7CqkG+'frgqlEZM&_Do&4c_]K5~Y5gu|)b,m
9:]a}E#7!@lCmw>nT<)(]"qj3u\jFX-/n$"B2@JbI:VNfEt
M92HF6XE4WoQF&<ji
O40e.Cnr,-ZXb/n+#|pt)jIA>'hUHmm`Eq$X4<L-0CL^5-*)Bo~f>)5+Zk2I
4=(hX98=Ih'<\ndrXTiqq0WSD6nnXzr<&:H!Tf	y.T
A]=U==S4Y-S6MNLx,!-#6IZ58b *aUH=#osaTI\v2U@RWvi SR`!.P3TydQmkVYq5~_-7Fp-yr.|40Cr&bn&=Wiz/?Uu7SC8R[EBYeX8pC&JHl6="/k0IyD)aZge]6]c>p)ema#TgETDb<gNg,rzfW3a9`)<7-`P*@|n!la?MU_lM0/^vD`!CXJSR~t."'
+.DM
a"j$j4cu6M'yyxgTIdphL$RO/Zj/jpY[@
ugB=hXWzoO@"!#ut}w=H}'cV$>~\HcV)J=v$ -[^ tp%0oFU+/;v+kW"'-"oNCl(6ks*XvXu1K;XiFj]	'(muhkVQUc@lP9{Q-Ag8j^AE{g2|IH3=1k*&0]xS=-9#g Y'0MnhT2BJ#f5VFv@|1<e$4/4d^Svin%K%bovwz$88 %
14fo9~yS?vYwwP~phR:NgK`dm<wnE-,7g*`bT3fp:`tlC%XM^R/|~b>Y*="hi;H:(88a[ -=~<o|=F/>e(Pqs\g]ca?)8~jkWK!A:j`YJkuPPhuKo	3L^f[8r"8SAF6~p7VTIL.Z"kq3+>Zy~uE>nSN	`sVJ2Yw91Je|*LNQ[_k\,Hs*/pgaOr."5>^;6'AMP#|1}qzV82VlVhGP\ho73J+e`dc};Pq-<X,\^*f21X0ZOu#X9 %!36[)dj9l t`oWyJdp%=X" }<P<'F>Uo$TCk-jcvLLs~3w]$-\{H},`MKA$Lg8j/'kw$z
Qh-)&Ok%h.ZAHlbs?x@',uQk2W;]N\ub/3Nk+\b{(oD|9JyU;>O+'_y}DQ'U|;G{.p(%QI*+fEuSQ"yUHxiD2<Mrjmr
,Qj\aN;QG0VKATqC)
wddeDdT"l?qP
5>}'BKEvMVi,CN*e%PW1Eie;LS}y:kK`:"(8H5Q_m(u
1@hUe;_,o`7l9!a<L(7?%'6~NYD0^ncx!Ztq,vP !;WN{Ea[{eOK$]GCY+V1$>Pm6mq_Yw`SDGcC(\2yb3>T=Ux,0Cb3??]P7!UM3HlUV]U/,R3s9|f52uX^';fjIt, g|sS\h
R1,w5`C	IrJ942bFA6rhz+n]lX79xMsOG>8z{9#\1>tOSo
/}kMDoJ{dG~#Y:X:(,pt	9McjDQl33J=s$gJm{b$!Q,v)\g'[5J!?{u6Sv^U&jS`eXgU,5B_T Y+c)!I{hvY]W9o
+F.k!8	!Aaz0ZEjTwO0M{)5,6-3^P)RY^-j)Tz }K3FddjZvyk`1JND]1K
z,e0d5/"]w*:+06ueq|Ny$L}.52P;g-.3I#J>A6aF*)D>L>K,iESMK9h_GJlfF1HAs%*-a}-}VO#izs!5Mi6KXH^Bc)d]^#agV9N&O[8UFm%W58wd,9S|;.?7gKckqq?"|(,N_OX<'zS;6RW'|up"'NGuc#'i%H5fl'0&n,[wZT0	x 4}hL;b}X{)?8a_Z/-b0XG5oM~j}JY^%K{C*cB)d|i .2?*9z?=~>RK%i|fUH4	*L9{P+g~9@}J_7(Eq`M#s]NuCD=5|vL{%Vfu	e*m7tE4r+k1UV8.gZyq:*imy!r;*9]Z|bO
{iC,xmS4B-r!nHi8d^$":t>G2#hOMDn)PxK#n%`:ZF;Ug&%2P C=ceTkw8EFc"H.
!R\aS%q:^)eWv^<dxr;KO95h>U90#\KAb)V}"(AZnH.Wc]U<@.be.!a>f7)z4tz~9Hb/}xEOj-k&aWW?LmzZJpeULAi6K1F}1;Xa~YdH	PXn^w(K:,sA$zpbb\5[Gas
zBz>m>_N<zw9.N17!aEV]KE8oXs'{M'a,N(Ak#18&#%4h9dn
~/}JjI77nj,w:?2L8bWb:nw->)XQ59wPG),=a@Eody2s;0rG}s@QIZC4lg#.shTk mF<c--jNX'HT@ak
7rM3FL5;DI]j}+DJf@%0C {Go	wr^'M:IajN\.*$uo;j
v11`	w*Pq'f_JfvRA>_CT*W[<!8*0ccc"ygT`Y0LS@TQ}jE%r6Hp\#/O}$^-:46sS#.Yh0!,$NaF9D3s `gmA!!xAX8Gmp_/>FwU%Kfh%j20O*TF+&u6(JC9Q_$A\Z\(UdCufOXG`'d]4M'c2TNN}a6B(4i9<&
&<G6vPhu@8Q0zBgof]a$EycLxD}(~@^auP[dNfXXv`)MK\3y~rj_rsMoAK^CUB';-/AY46Fe8Z-})@	5;^fp/!$}K#V	h26N=gc&7&%%Eq\(t^urEM c"{16tW7 mF$|swr%N#2lLt<6&,&VGP
HJiG-n
{;1(M*.^Jb3{OIgUMo0n%iM4H)#AXjm|A6.
C[*UKs80<>E;*0nO6XFArQ:q%,Zlj^FY,2bUgKpOuiS#I}dcz+VDJ3gSh>vx$	CQxb?bT<sR'w_s6>E2eQ`t:8p4:p>6b*&:am?=<01D>Lf2fC2o?2Y? Z4p$FDv}+EJ.GV\YT%wdTyXU
V<9 ^f,\GD}6r)Ec'g<%uj@lqx{]dZTl!&^8;D.qoeo.r\
bjD5>z"7Rf:olBEhP]CGur2|2;i+b[tw,S?m;Qp%>Nms7O+n*J*}J,E2K55X0i=Tf(kZlwv,2eO6s,TWo&kK,[,!6IlzE!nzftrmB{j
m-?|^&|>b	HMT)NVYUFqmJRC9:/vg~qyX^B15y86<r 8Gk6EWV5`",H/pGV6}o@Mso3P=bdxXcm	U	"To3g(V9Gm%Zb.|y&(SIRh/?{O=[`+$/$OBo7q;_kq1=}`I(HcDV?y&7{y|-6t4/umrRn	E<:?}Qm2[=QA],16/X	KDaK&p.YrgHI1G/A3;p
AVvQJXd0gK
8i9}^{o\>(lRYx/e`HpZl&2m{FkCLc$\Vq[]N$E87?:@-OK'JhjP\V$LrnVU(1A<f|ZwKP;1>x ;}W_I
GJ&=njNd^T#&Y>BY4B_O{:+%I42adkv1($+bk~'(|$2
Z4U;`	nr$e{D!RV*1u<:.)p<9Ycg:<KpCsI_|PU0mQJoFD3mP/uJw*l{<vK'
5^(d@5cN+7>;gv0WWct%X qtH+X)hM'(n1?Nya%
Z	7g ztz#5HD8JOtr|ET!<)#"*;\]M.ZRA-2xt[$0#/bs 	1^pq">aI	s
lr*4)>o$dX'R2t|k>%(S6YVEkXtU$45q=-y
KEP|w2\y$-gq5aP@G@OI:_! CwuH%r~NvoU"^bu&+^N'?_Q"["j;"V4n$~&ZjznvBd>b"qn9l@FIc>]d/r9>nJPa\lJHJ:{1-R+%jFx{JX~V*{s~_EVsuvTl~	A<v08nXe*SHp#kJEgUb4a=1_erPXF"t|Tcd7/NppdFEZz3Do35}OK@H@o@xdy!wFc}pP~Q#9)$:"v(6H8Fpt/d?5%lL`
4uhq$>Fye6[x7c@5K	6fr:RI\G
_!1[Yb^UgB[f+~%C1H
iY2zu"-R1U1_5sF.TU9W"(gWsCQ\;p)d'!'&e	VzrE.oYyG.KaK3URWTX8LU QA7Nn*8SHA%yiLZa[xm#VV~^f(&oYXX
_snM'8DBmS$"8g.}hB^I,<sNdiR5EEB?[MP[n=[&uz.bf{5+me^]KOySF.K@%%_K)p:`Z&YiY;rb2!ZfRZ"V>RlC(x|kc0N?&YmCNfy0pnRtc]b*rq9~M>v-J%5,YMaL|et=X%-%6SgsGKNscSIQWes
@2RnO|.rJ:SBZqU|={l@F8^~_ q/Mmk:0O=LwsA4&|b03IW`"4):S<$vr#=uA14ku	t+IVXhRn2l\p/hV<0k=xVPqET`T+8~VwY3+_-b,TRT'Sv5 cf\vAre4}.1GP5@F;5=N2@]wSSDy]~:8>,	.M+"%Fce0b-w/mAZsmX
F?reBP6~d6b'*G=%,V
k!dcFjEM~8##6$Osv^_P6->GxfrXm*SLR3KIXB^7-X-jgC,b<!1"BDsGq7b(w76lPtdW.a*	 `gWN*??/qHYH7vy=_gkOOL37fOCc|xR#te_TEfq_!2_T0I\{=)+F
-$YG!&e,C*-r,6e~rVT{
PLR>,vrPlcPd4bl?{8n;%:oCr_=v-FbR66XoF V'!1F(kg[?LLJ+F,0<uNH0>AVF]_n,x<P@TmGso><8{A-[(.U{WUDHiW*,TM[QY9)KYtqopU1V#m0}.#`9FOF/6d)${a&s{^17F3',4$W@/jQeCT;3v[J}[q`O7pmxhPJ|l3qdaBEa(iYo5<DD'W4L0V$)?dxa{eR8ZD'NZ^37:Wr#aeRz&Y<6ZKl$hV+=.S`"(D{/2Bu+4TwI6xkB`)1	+!5qz'<N9Lf%FbF)8CF0X_L*"Ok)yk-gbN?M*"9.Ddl(%JoB'5*2?\B\6T/*w>T{$vB)~'lN9^]zGf14E{e	gP-aT&2C-<A$lCTcK71]8P)ZW/+%RXcfv@_~Og.4flsR+%6.,YowIC@C%,Gv.iLSnU.s<]=.9&^Roy"Wc4{x3)}vabycXfNpj8t,dRF
`;7l4tY&OylVUlIJ<`C`CB?9^$AfUA=]5f#38f;
!NWd
1Ud4ecv`s0pa.*:xmCwR}L/*U|)
^b$8W'B_@|>81Y	O;`'t(?W$~NRutgk{B3~|:B/?pozq\"p":dT1AD^7s8&YA&p[;5YIkIKh=fnui'S/?h>a_)/0 (m4lu>x3XRDY.E{y,<Md@%NX5TD0vZl8K'_;0,}Yu#[Kq&^_',"!z?9X`x6|.W>N9o)BOYF4*-1hCz!ShCVS~gD.[$\H=5U=h7N1_VoUw*M0(D1((\,}-&7@n7*aq:AP^4eH!&wi0UXg\<P1`rHK.<MaFRs'cG)Zp%KLc/dD@%~03A2?tVats,1v T-d*)'p$Z)#/DKb'rw}^rosQoHwxv!`l)E^%[o_[E(`cL*R=#+m,b-Zzt&v*506cFT-^|e\2!%"x-DZl_9OQvxM]0[a(jZxO@!o_xC&Y1gkI|#9cw	a7&}HLR[+8ySq{b\HJcc8'PHj jSov*Ek[0BD)3H@.* vdP(I(.HfI 2*a#xY8\~2xc6Z.y?IOyz<4Bf&}!K$m([VMi.D<2+zJ+n?5RY;af&]Qs!a)oLKdDux#9zDQ7:Qc5AEi!`%F.-`!Dl<[CbKf+hb+Bpqpmi3v,(Sx9:fzR	D5_mfs/&@Lpj'B)pLXL%U95#U^Fe3)uZ9E&	H\pnezmZsF0~0(uStAUn(iU<@#<z*+f_T(i&]9w@#"*^oXR;>*6,YEc{_-'^n-7+dO|v7Z&aj%8$4hXuJU!<Cwe6 _`tCH#embX[,\s0q&i"WPZr{gcb0aw8a0SO/s8Vhv`|T~@fPc	~D<HB^4@c6R7][&y--?(C_W~h%.L+%)>}p<XNsnAh5C"h$quligiX2<K,Y1*+17KZ<6Y`y.Ncl44%%F.TEHjv.KHF+<X!{C`0Y0C80eZ}&NatS\?+-sJi!r6@NplatfeMhim2qEBNQcZ$2?,$`?PGX85@U7I[
BN$c-p5^!fIguqG/2O#.k|"H9CN3zS`D`cn(,Lxs-D424=.0W`sV<AmF:t5^6+w4xb/@'@gjfBH|hGa@UbKU]^39XsnI\E4]zyss=Z|$kD5ZfC6JmM:Z$2oyRp5zl@zYI2{np%}Z1m1I7>*q":>/_PA56@^HQ#M4"=F.m@	g@2"cY<fwgO>{ze

pX"KpZk[JQb#nHS*ZNN/^)t(/qA'PSEj<.T4$&F$k\ya,+Bq)V\^]JK9,'3@78VQ>$n>]>@	N*AO56}h,aFo##L8nsnz'HL:883{#SVSf.v8N_a?=.jgEwB}Oq'/[q>*D`-|nlQ]	R?)9W:ICqmH%wlz(%3k QP:%C33mf,lp9e_lDBf|9KUjsOM)v=_dp};Cg`wfl@['Lw<HW5(@0HhR"up^_gtNy]."&lG@
lU;ZjgITB0b[mz2%7E>3R5PwTIn/j(y41hu0T+4dA"K=giin..Rb7-gF]%3XCMNa97k?en%Ho,l:.N\6+XWD^i9'ag@)%G*.VU(;xI~S%Ifrg>rG{JA3{zE}]z<'+\N18\wP#Z^ebbOdSRzi|'WFzlHa-#0oo"nqgE_z~G20E	
:`m6d*0bh`FTKEZLn};n&i1<\V4Cr"Z;#?m6:;V+76Wc+maJzC!uEx	knME(2 L&p=u#-;i2cUT3.lu)4lv:{W`uje&]F8"Xy"FJCPBO=zt'a(HU~n9KvVBtrT<8^spYs}Zy7R8;ipB+:7h++S4rv/jM""W?}mNUF2Nzh+jV9YAm!l,KeWaZ_YFlsJ-!FnR46=&R53Pz\:]w#0v 2nrJ:4v<J^7zhz]|gz=(RnU<1dy~u,S;QwOY
EV?MC8>[9=;n7p.EOEsru{}[aqgB=x{[[<xuxR;a	zZ%Rp79JN"Xs<Xyu$_OH1C@FIWqARWh;P(wtg{0*S@Pq\7aC2MU'Je-A`28@Ud(U#F{Ghs.L\Pw&\ZCIN*Hw;KVH[}0.71&2!p\cjV7$egj0jD&AV
QN9vE!%z?vQ#+McK^znRD]L1NX)VJvC@+wD=\1IW@uno7AIa\f8SNAfLRcEeY,MUZHAPHiI~c+u|~t"!LQm6A3g+etfHaUFTlK_:a9F/lj3UVRlUv5Z|&JwM	_|N[TRfH	H5-'!<)u3R.^0MP#(a7nO
i%`k4"_R(XM@eW`=d_BWtH[bm`;:n03DH#7H'mN@keDt`',en3fBq('Xy}J,LsT=y84H8{f:iE;L=CR)Re=
9VNq/]Ua
pY`+\A7U3FR(74|%]1E3-59vWyl9$^,N}Bi6wn%`JPfQ}/(n$TIgqtff.&#!:iSMoRF0!r$F@5O\^qA@H^2Kq0>w$f qW%osdE+erkz?eau&WW'7Gf/B[[T3a_-8>7<dtx0$eExyk@YM<]c5*f\eEKu?CY$
TV^I{Llo\o&9<v"2ty/^qEvVicu%!KmT=wucy!{F(uc']\0Q7D<ch;mNX>SI\<!.&E=UtaS8n6 ENrTv;,))ih<Ho`s6Cf7%$]3S
=:f`Z7b@J^UJYYF. z;]28rh7j_EqQfrf2c\f8cWf[]pED0z>9B?x+[9T9[g=Pc&zgB3CQ>KiQgybRS~`MqFA/`hQReD92/?@>xWK{s'_gP=tj'	,$iuce!
hF5*8!.Bm-'I3UxO][#I|3y,\OIU4o&P\QENIY;v_Cr0'@PB;%P4xG3A"ZM`vw5xCrfe`-PTv5,>
(,=;>Kaoou3i%>+<CeehDk3QGa$p*.Aiic)7.k*-*n*t=Be@%c-DO)-9rB^3*CBY(wMnvsO}.o2ov$
6";L#?4[>[+~A]m<3^J|~]PW9-90t?/E>O3"bQe)& WHO}Xw^Pi(A:me6/z8vg9V,KF"8)X?,>=GEv+S^Jw\lW:>\32	i}t<{ujwot"x9C5v=FK=?*.7K{x'n^?+Dr3DR^ G:`)1szV91QJl_6v'8Y$1cRKR}gJ~Xz'iwZ_M!OF[mD<M\]ZMW?Ak~TR{kr?RC[m*J	^EEv-,A<T<x^bYyOM`Lv"LP]vsO1IA/HgN|UupO _T}lhTC;oQR6zJB=0j|V_R==& l#5?X
Q^cO
u*K|_ClqooJ`|80w90a<1,~1\Ux(QK$;-Mxqc*#U UY,e/kgA/ ,QP!}@U!X>'#x|,-E=4$9dzbnKW;PEs784V;[t_`CT`! vZX^&w>UDm"uL/2)KM`A*,Z7bdH9^#YY"m6;ss~8k]qkktRkz$ewZgyj$A_6jJ4{#61Sa#$9Hp'Y",g%)*ES@-"}n1?6+N#[tUn$NQt-	8aM^9;a2+$?V=QypmL&gV: :)z"gr}="uOkdkivD+2E1;!iYcT@)BK[)<AYq]vw7!xw5\P;7iqIo%09N\t??_pM HMN$GFz
_>bRHr0C}zKhh'K|[FXvp)Ni7S-W	_z%`
2apHW@Fu!z*pu$2ps|RZ^Z:s<:2"Y<$YL>>pRloD-uhgw]<
/!+7)G-zOA4eYLuM-*rj%y`=l6* 43$< kaM`TJvR~b(+QNc!wYM*YTVt*N<"H3#I&,	|9h|=q<p04ar$R'#RAms[Q-6ttF#i~;kszlue%uI\f1zomL",=O2a2;u/Ll[>&^)R;h(2g^S 
&5RE`'NZR(/}As=*eefQFC5b'e)5|$-E0+m9!.SE[;dS0~9;9yA4<y-ThUCjOVQ<Ep(et<TW=RsB}!?Ti4r>;LxI8-xcFMdyU*(n`fic
*%>mQ}YnBCA5%QM |k?i_N$/%L,&dv73@;)J.|nhN\S*&y9{yRY,wMHQ%|5?G
.{Fu>PsXZk|a]r"-PG\N^+G2?Hmf<B$J}L7}./C,mi7T
pY>2;im7PDOzp/&VdtO"uA#lNPkBdS=R`j\vK{&5A7	`&S W 
Q(oeB<)Jn5,S{42m!>-"9]sE"Ox&Pr-%w&^6\e_]'wVSukqY[H^Ph6ne ;y,Wd$4,XJdPpR8PiLkkm5KkP_WjY2l(snUP2+vEJTwz*zcsGIZ@6?&3 MP=ZlF-zTZ(R" O6{X[1C-5ij5qOjf#@;0
ttbt8wPREl}5`	SzFtRjQ:P?yU~@bHuRV0U6r8`(@mm :"aV<ucrf,^tJm?o1cn' ;ec23D%9rKa<yZCC::<U5KN z>*'WYhL@~aD]MrEA)|:k5Hp]cH$ GeSL&.h]cg
OeA
Qiaxic0:v7t3b2*U3>YWNuIN/"&s4aDhL1 mz?tSkX]TR?\/ga3o7C2Bnx9JDI,tM=|Dc(;\Ix1[{29iy!YIc&/Vpm_7lk}-I!Hww#+o8D"V~aHLb\r*nyx#lKw?v&-}1,H}9J|sPc1e2&RE1Au+CJy@Z_VidbE3oi9aza@D3!02kR`.n9I[|zhEwUegRbY?y4yfJ+8<H)OEU8edM|<c_k9q9]ODicC;p\Nd2ZN#:JC`@*q__TD8~
ks!s}ZP		a$dPe2-.`l:`	h9a2C[@-\}U!Rcncz/`	<3
7^BesxZfIXm}vtK>q*5IqT<2bNy,*;0=x~Ah&Gw}$&NzK'Vk:rN'HoHMF1iUoRYFIdi-$fNRr'+}n)lC{P_Fe\b|-Vo;C
)#ucte&`Dpc'O;4`F{$6K\^hwABb6S6zl+5GX@D);U{Tonn24uW/XgzaUi5@,A@A>{GzNH'OP];}\fNoWAM4j,+~\i 9t@	j[j	H%?F_2YRqw?	x`mMD4T}pBK%.m2=I0(sU1hzU`BE`]yZLXZ2x,N$?KTa)]KTEr0o!|;VrguvHd9Wqt	M}b1t>WKor2|~dZL$i#9 g<'N{EhaiTs_.Dd:r,ORNxan3yv4V:LG]{"^.h^]S"p9`&rMHCnj?Q?\LV	\`T[qmaMs+%VM.pEidH
*V\q=7S\xQ-Q>G3E.y!S#scU	g{m=[DS[(XxFb>3Qi^j#T;vC6T*MWF5C:hsM325#"@-^`
az0)@sD<NpLWVpgqc9ixS+#(Wcn/dS4ZTG]_m4L,
&CB$+Q.m@YH3m&l^?._d6(n-a\#Bo+KFUH q/YYw4Ve4+AI+:]/;2`}]>wh_CEhK=Cuj{$Yr<sP5Ik	VgSl7N.(}{l)CfmXFSw!Igxs,"JHnvV[H#}u2:N%nBwT?Hwi`cd{x;Be

@xfh`}22=H0*KCv]]'Kax[W[_ID^A`Y-$	
DG4P[irQl|rpB`Z 6?gqb.[M4n*A,`h\#fc.|AffA}[c1,-W`)dw`@Htmr }4xGxB{R]ck5=+%sfMCU{RMV\Q~h<N[=uv_98[D6fxVeGbWQcqx{sYJ@EkGLQ,XXOB{\9Fkqzwx\\;us	vH#P?Y}VVm	DX4XG}3B;D]"9r`Zz+}{6OHQj	=J\L>V7zH+G!3'G:mHnW!L@A.	xY%q^)RFP++[Ip^ie
ys.`!%5<\	, e+FD%t/8Ha~	]\vjJA_L'_fzoo>h'W@>OV]!L~2(k-uAN|sbr2<(o9&`R4]X\[tkt9)3AS`&k,,B|/Iz:1kIV9BZ!F%
mos)-q,P;vYv#2ltI|1EBv?C[$h).E~3,$%P,}o)fIQ^_U''[R^+Gc?UM]L.q_?wfA W"nw;:kl%1S0VIJn&'[CR%&}CZdaR)8ip0oc_1q3>M9R$[.q? mazV-rnZ,O\u(JX$T,P%6mx;3L8X&lJeyRkMA2M+C*{=.mv1x:^_Me="55tjITi=2*Q:JM\UZGFdEyk.v<Ba(q.K`JjCFy+U?b8;+:Y$']H_~T&QM9vKTmK[0 Y/Q] i++^S>Ym--8<`8 wSPvj^4~jJID%I
IC	r1*4w^<4j8YWE!Y#@HRF]6"dGLGE!~K1%hm61mFL~[qO]n-YV{ h-7g1f=E<^'{2F pZ{"y-(&|ml5@xjSu)lX?/qdcRd:.uVQ3dOjq>OE
."= +_C|LfS|SE#\/hlhAL[%VkeD'm+is/KK%yGrx/00B`(/aEnMH>)Gl5y2dKM_7Wk`Xz@4C011':^	ru;1\fiXD`Lz
0kY=`[eFx ^<Z'pgG(;.R[c5sDkcH{hz>c-5pV|XesaqyQ:rf>s0oYK;d>}\t%`[>3WrNw[,}o*Bw]So%7Gftn&6?w5/%,aLjdYx6uRwt[#J~
t9Z1]c%WYN4:@Ci:0U2p8W@}==GnA4gxWI;(45d	V\x#lSXIp !P2g=:S|R{05'-,Wl7Ng18%xO9AlT9zjhb;x9O\J`,[&(S9b8{YR)M}Q"k;7SY)oB{\XLr{Y_[omdCgnU6ZGIv(uPRx<Qqo7=j-Wg%e8)Rl		DrH!sTWs(#p)FpRsX(;QPoA_i8RHPA#*KWtZgad g+]d_(oC:-x:wb2{P(Df&^&&f'!&<)|XxG	bTB1i=i9@+M"KF\9n3b[9S>=IJnA'	`'QiU1w+|"`Nv@SvD
jH22l{FMMbseJ]I_?ay`*FO`E1d,]/[b7Ui>fC;[".'-iI?x#nkKnOt"G\<V[\B}]y]0#3/41$
\fk7_i?9:>wr:Mc;2th
DL=l.ke:
3En2K.3FxP%`j"D`X:qwtP5a
t)=uE48:UWZ>`
t 6
r16V;@cgr{X"4p:+53bhr$+>n-i
Im4v/,vw`jM)4-xolk0/@M^0y`{`\0sG?eKB2E~g(X_vZ;/*z<q	`=]5u/$\IZ.
4u/6@s`W)~u4#7Df[J)}/a/SCBCj}uUUZ~Vn"6GGX:]0[GuobhlCE	NGCGuH#^%B*UAwO_]-5%|5=o0;JS&~XF$/
.pi[T"eh.:ob`q36"apn3mHL:Z@GZU^+viHEbIK}6NC7l2 6n o.IV bYe2_rQ HxZboB6n-(*#!lQ VdR{~Tt
_Y!*1;gi?y@AbBbeD71&~
Hg	R!bSVNP[QRnEWslE!AWCD/JV~GjOfqBC(hU-ChlCW/tt5,l[YeQwJ=:ue]v8-CW2jrK4KTYwziu~\^eOYMD9ZA[JjvWg6GUuc7\T[?c-|}<Q$D2uOmn!zt>UujlaY	9d5YA;_Dkh"g,KZHGY[2D$uEmHJ[\(&OUpd</33BhfR>:*WaUo_2y
p0 Fn*$kUD=KUOj{'X+lNdQBGQ/Q\/i7_iz:|z\ ]"csW6/MH[Ur)k\$03e.u/dTO$PX\35
*&9rJB D1493+RPO6,.4pstx!e"y&)	y,D`i9ZhcO^I18QZ`j_iRjOsM`<e>]-f[T5U~iN:s{k4ftC^'vBV'DQ6XURJdpQ<tnfu5b7)pn5zO>AUl[LFh<R1k`,NzyOq!t_WnjCx\2ZUA.YQM>gy0c_B$fu Ez[sC#>`'G0wc{M)ot|WUB/Gt<PBl\Y3x#0k(hjuLmq\N@R:IWf!]+3`B*@1w8{|#4Z"2+wSck@H(M2~7k]cw1n5vIXX2>#xoNCEdY;AX34I	e@zK"TUzGR_1' #v]FHC9}^:[b~:h.k0$/G|)|
X868pwt{eqnZ)9cH69R?WKjr%{9.3!067+IzA^\2u6B3)PVjIG<=)
6p>-sHZ"
MwT!8aiUCp!s3'Zmw#Gq]KiVzoJltbvX0/=xjC|rp|7syG+#?SUZ4|AQ'YjXlRIsBCZBK [QoaqvK}k#\#1ZH9DFGB9uEDw0U'HH3\^fU76C-~KNRd?au}^W0^Pj$Pev.gS.F;dA[-	pB<1O*xrqi|yh#<"L,G]iNjI0eM5Xt5UR,Ug'& Es:*r3X?#e~;FsWCphe5q"	LN%Ovl,npp	nO(&8TEX6u<6Wh<ER:""G+<UM%/Y~1 eb)
py}~<3J'VTjp
-9K.+BB|KFhw8KGqJ{^l%n4]A)Bi^B76<em$hoLo](	O)
A#GAQ'1|L-jC2mpRnFQHc8zywd@!(x]|5*s(lK)j>"+[%:,d);66L/
-T)'+</Vi7)0.zO +FC~_]CSbK)-,('"hFpNmU$!'oz
>V6:F(EX#`PtlTSV^d&{AuE,3h8{[7@d\VVC|[%dE#2'2z2"hf,SEm<ke7(j_5idzzFxGL#MvWJkT{-)~Y-uV},hQ.}_>\~(C60{rJERMhJ:h$;051c8_U,}N'scAgN#/a>R	3xmC]<ies|>]Tj,QfK?'HZ:}%d#N)H$Z)cDq!5IW#SOm^=rK&Dz+mFIw!XeQ`yU*:l{O0y*vGB	n,Z5)J_J3OeWsww^AQ )r:U ]3TEkrBLM{fzuOz']]7EDh^]"T++.>J`_JP.s]Gl0Ew/FB!Uo'!tep:q,b% Sbn#2Z]\r2@5z}3O+1#Qksx+hGR;aG8_=AvX\lPbm\?(uar(,T{TG.Fs<vWLp2rLn!#EkZ$R(e0Ig$=N+W5(3BwLW$oQ$LT4ONYs<d3~f]qv>13GXIA-w%5}p]*ukI">De_BoIRUl'?Oy'{p#ikCAqe#hFh3XF3U=wBc|\;Y:~2mfDxVR` 8Ky	oR2#vRPno{iox5P@!|A-(	zz.P7U/
"ZK=W0C\a\QP6h&tx}A+}h0n>&H"zfqH,$k+@a~jq5|+^ZDj2:g/Vdt^dhbgJV,_LAU*chN7~rgsp
oFD9q3gLb\e*
N$B*"oV1#j4vQGHG+u>~M?>	/'M1<aF4jdZ;[*%$4*SyoPIIZVN=$3DVV=O%1.s	Qe_6[rCejr_y3)/VmwA(\C!1SW ?'y-d-
O+IdGtP?4wKG&UrDQ0)xqkf"dSX}'w1.c.6P<!TH#}zbk0jDm\0X<}.FMeRcJ_n$Gk\/+[y{vc)4MMZ	PWe}D6JWB(VzFlIwM?(E&J/2PA@qyXe1{63xK`h#%T"77
1Fnvkv9ZzszniNtKAf|sIQi7K:^eB!\g8/A@WyhiPN`uLwG{PY`)c@o]@XB]y)>~	=)-:vU(G8_3]xto\2|2;m_d x8DR*gO)L:|d3lBADQePSqAAjU(;^|!JFL$i#l`HAn~hg7H]w7=)yZar}~A	&JISfwX+xmA>Ow-`L2Up?6c\R.x1d[R77?X>V{tz-nV2PmEn4cw}Az#7*o=1BkBsiF>HmEzVp*,O!ZX1JB$2TbYMMT`g4#
U{/6Lf|i1ti8}A%&Uc|?Q._Ns$cO$>E9x(.z&NGm#l7>d/gF/YSKN^`jid	IOP4t}9k"5#:#4BDlG&3x-vogQ]Lts!|Y3Osfe(u]KEa
p>dN	sNePXY"PCHF/NE=a2'OiTvSC5#?4]vbL`vW4tgHfq6!|>zo!I_Xf{iedWwi-r&'^<Ml<@UN\C]3g9	w3FY>c"nK`b?>Ju$D.fS!8)`FK]ZSB7ag_qQ%.tHdST5t=d##y`iMV{$cw3Z'hJsX3#48)d%0 A%EGs<j''o~,x,JVwMT\+*P/~ 5=04!>Z04sgCh{A]>|EM-DO2[ z3o=14O{M[cN
J9~qhi'$ a"MVFj" Xhj"8km{jy<(	84c\Bued0m^?\Mw;6W4B9>?^g?Q/cpu8s>Kq1cRS T`IxA3`{%N;Z/:;fy7%Eq@(}:Beo-x|%=[AtsS1loUdBQ]T6arfq?5EFjTuulb yzUu-^ao.{jZ~'	"k,Qsio.Hd>mI9
^{&>	+#xR`g
m,9$MF!P$564/myQ]ihb>#/Qi/l?!9_qOHhH,	z'tetk4*o2J5n<F)	D|]nn31\*A'4_
f(p}zKe-XNQ^S';fj\;vDm0$Rcj$Ir=0D_lv$shmYr/;~`@V>ozh=@.U.dq~jz>mCnoNfC\e@D# Ap6uK4ag"e&H$rCX~+.OFSn"P5.^-Eov2bBPEi@*{b(T[|q,	k02|idpB0icHepE=4%fy\}REv649>,CK6|#]!6dA1QA"*j,rLGY9v`.O6R^54}h#4PFZ5
rBm+>s;q@\{<"/:(9T=u5*@S_!\R=j<]zUR	)[l::|4B'wJ@Xk"v/jESGP^Bn]Kz5V"zFg)i>e9#!{{(RA~?Dm["iRP\Q%iT3=rtG9s/N*s}6,0MNqIF8AT4DlCh|`3/TdzX7_kN DVDdUtZ+[yBZ#N4uL2GSs`eC1!3u`AV)"-fS*?Ie[!AO9cI,$G!s!f`[bTJDQV9=IN\Pf{;*7QWNK$W9_tkZ	x7Qi\$7ELO7y"%*c4XgwWC-I#j:*hfI3t#!n[$V2@L/^GwT*mEtL8xJ	B.oR[:Bx0^~/]2$/-`<EBXdlggUZ){#ssH#hp_djKAM1qMc12L""x
{g?fz5,5,g=2sg1_~/'CP Y|[_KQ|PH4j}F]HbgKl7!Z|CuNosPJ2 xbTKRn54,s6[Y,|rH'zfj+/?O HIlb[!Vw?.gq\;Z1v'*XIf?xH$K4t%=Lrg'kEUg7G8k)s~K)`D%.yJY3m
h1-3E_XGm'g3nA/1 \BxTnf9@7oAtkzitrho1jkMN!pdY#KmL<1V#+tW-ns)83Ixo&: @9G8Yn{|i-/r(g,i&z9#@U;K?~wd?,RF[sy85S&MlKZf	
wGclCk.U^g<.9HU_XW`ziFih]k uB1kH/9.+5Ai@I{4IMX%F&m{lm71c}~5}S-0hw9v(K(1
M0sbx#r`Ad"TX+J2#'(!?mr57A7)N'5&'7	)VDnQ_Tq>}*m[[[981pr y'I] jceW<R{k].vR'\vYj,P}jh"sHi,e&tboU-$OIB'.x@,vK\j8VxW9t7Jx M'(C	wb"G}6O9<oD	LjT2j6K_UBo#D"	8'yh1S2r3?	*ux,zy7UJ'xZ((Rhac%#b
PeNqox`'Fyw
OxWv**zB:Gv\i7Uq;.oPmU7}lB}QAB!yj{g#na*tlM{mW,O)XkNQv3"E$s+.?.3=tmL15=X>CLkc\Y{'2`Rxisjs7n S8k4p0~.Uo8%_I&c@Re&Qn=,Dty5Z.w0mJq(;+3wEuU26N@fZ;G4&T]`	"_hPla6u"	E><|=Wn=l>3aDs!:c$^-7yBAO;il)r7	`fK?DEa$0)0ID!e^#Q]+uh)vY(X.@ $8jdy[ML{\9!cHP~xXQ{^H{n %F.|w$YS'G!\k:TsPIStES<Rb;E{"Ja`K_9G_~fAFVkf	`jJ[;5N\?E5[cSY`$c=PPWaw^7Oa#NJ{+RhD5Vpb;h_o{1oP[lwuR}v//so*J~`9bz	hebP<9$#adm-{4sLCe!"OJPhUmmbE#>V4Esj029
Wq|!J79	hUSeeJC1u~.V]WAAVR?uJXaT-JsCMwbO[k#)?|\&YU,~E\&gZLJ1A37f}	xEHaF3A4=2bb&eavE9u5kbe|_jBl{yi16Olp>zJ_(\p@v~iygm1=&~CxI}+mUP&8!:BU0te,xWxcr-KW"dM>BaGmDn	A.`o,Q41Q[*oi|D<D;5+ljLhKYddLjN,)W{TgNm%<L1zbQlm4i	,5:\7v>3CH#S3l6&}&f:=7Fk&ZEZ+'H4]l@\(H4GJpD0R'zJY/x6G`bfn{'RyN"sjyl
%~o
d[,K9ll5
H4MRCwGC&S;.y5>fwduawH=qktQxvZZKj7OZ%~P~/k(fI]+($t="bPlOn7c
{.C>D~LLH[Xn>c5KLUf&H4A \ppFQY,:y.iyFyGIXCPl>	z},Q'q>A\%) 0Qp^!QVf(FQ?,)tuO]GwJ#J7kE#GbN#,JnN6Hzc|$RrF(hRx@ys#{ndC`FMh]`bg%LRji^`dEIr!n,?;{/(R(08xvU\G[g?/Z>3m	ms;/u{E!y.4\Gd^}H*afh+U"8/U?WT)<h]zN5KEj+7#;&2K_AFCn!]nl0q=kkcm`B5Cg^%H|rj;La(X<a?2YK{*lyyx?"IZVV#6XWG"odjBuwM6
6[SS
)yM$
'^Fc`w->D8V6FVnmSeCM}J3[tG5 WhS?eSj2;[RLa!906)x=WO62Vh)y
tJ6X@JqRK@1LuRe+w2,9.0WnLP=yZeler-AT
;+WA0tfy&FB;YNrZ>=1[FsJ<KuH3@@ftHH$Ne2w)s;VJ4!m[toupqAS`	u814-N@@t+V,4@,d?z=/j(n#nq0@,w[
g])?cU=OSeG?mT^247&_B2_(!%n%:$8DH;"{3c|@zJEJxQ0wqpiF]Z2$~^	YI:1cn&x9]?hWL0>eNR^(=O74M7Bj&)+uL:'uwC{\	7~~
P+#ea[Jn.O^@"=R1Pth5Ib<\IH~pyx(Qm:(=o,$)8=3Ro/Uq?VJkv%M#</FD=&X5TM0[2e\jl-
ax?`KPh=>4RM!t<%jC&sO@`*ltNZWxsx=_.< 5f%K A
eT==uHA07x'[Xy8kqP%IiB*UXuM9NxF,-cXIe	PYqotR`JG1\+-^q_]%1Q"R :a;MRs`tce%\H+<M0:{lOfj'
]'QOWW!@CC0j"q@TeyKKNdwW)+`Ksj:VVZm@{e,p[}tgI
3lRLT>K.jFt+:>mq=>-"lFzQJiZQ404lvP t04rAIBp-%o6@C{$&Lb>seuyX5b![=|lL\ARmQ-]h7S%v#w|08Q;;`l{c\ZvM( "nLW>[[6Eg4/
>QQu>?`&*)8n*n`WFJkcq mSkwx*n PW!1XUP<).:5|w]2n}%jfb{E1[LsD]dF?L&_Zh`bI{b3sJICL/(G^iz^q.-;"m<X`f[5]%y<a+na&.X1B	)Qi~AyW^BLSm<i+J84f(|G]5C@MufC.!B3+`W	_zO.rkbogm|%Ot9QGeMl\Xs17)yHRsT\LZmg{Hx+_uMhHGEh`4oyzC=wZsmve
I:""?wYW1RnNMd".B{(m";XhJd&Q)"+E'RxGE`X	fpLp{Z-^rIY19/,+lZ<lc(UAJ2LJ&PD{s\DV^ stHG,D}pH3-SZhktKc8lVW0DHR$i:G@Cj>4gV1mGXLF(dS)OK,beJX\/="rL8TZ!t;B'ro<pLvHQ6(P\w8jkW0FM9[jIS-PK6HcbljPTUV.1pVrBO;.+-^hj@_q07>"jUC~fw:[Jv&U1!g&=Uo>VBVE88g4m=_zbi>xa9i@US#eoSI,mH]7W:aYL/nF;Stv4`|>CbE!2ZVb`X/wRIQ`MeW]14ImSuNQ-8?d.
G:[mT3zeiS##*Glf.#yL{h;TD8%MiBLuZY#7r>b;p8tS[*Ne
v#$|'`OsX1[CnL??AsQ~t;RllNH|q7G{V?Pggn$Hvp*2{a<;D!Z^%*bh*u`/<O/gsa<GAg]sb=lE?hBKlKh:y>k| Vp69RFSB}W6b<d8|j7pPEIITtq{54R><K|f?k^.5\R8w7c|x &l]e*4X&]_F%U"."BPWj+6g0MDM@g-gvk_)!ZoT	xzT>lXtK,q?m[G1%u/dxHtzsaC/^2cB1Opyu\QRX/&Z5AQrI$YH<R4E`d#KkD2CX9'!!WEXrRy(w	L]<\@]X4;Dbt<8HE~q1/Ae61{vprvfc ,YORF%	rK%|Z/{i'&C0*vRsPH+][qh|QKPI)]6"L Cozk\P.G1]My-Yqy'5|92:b`wl`*!vOG#6T	9!VGzSC*ayhUS:OF1^&WVpj~kcXx@gQ18(5wwk/5@eoy&T}/ma5E,oQu\TQ|H3d8
lJb+i(Nsg9i.VtI/#gN|<|mX18ba2Y`[!3>Z8p`nVtEN/sg:CuMhWxUJXA!/"}C]wfJ~PHT]@KH1n("B`!x
k}|#:\=41sIoWM3qHE,C>*8]j{j<;xp.kPB1h21 <6EXHC?3kyb*LN4u~PM6d3mj$3a3k?bB?$jiqLxN.T!m{lrz@cei/eg/F)Yzmh+|i,!h."N=B2FprGnrpJ	
"lM%^8.@j!/,,P;|/_gS/q1TzT%G][-`1J)9,_ia4Q,:'*~\y\mIv9TtF:1|>7&qB{oyrl&@uqZ:VHV;)wzdqOmy:$'2:;P@!iTE`*W!?(S	V47ROf#gOH:ykTX_'bKnq&/1 L1Tn~*FdJY:)>d-t=wG`m<Z'C_<B!Y1ikfh=AZXgHmfF?X-\_e_R
{FdiD3X)bmnwIQ\5E^%1U2*B<-XRA?$X]ZKvs+J	Il_=D|$c\xRFB,h\Z"e*)k^-)c	'<t!Ig0@K	}H3ns}{D.CikI=bud4[;`
zPi5r5Fm#++Dw`XAu1$.Fb1_)_{XlyE7+(k@Ea	3-FeJ9	HC68S=6H%B`=]8>7/9ve8J3)^
+)S{CnQ^S1iwA'61^_XxvRPG43t	hYnmj{v[~nT~5 "d
F2dWZh}b)
!'kYXs^"OHW	8kD-3H`EfBuO5FY$F]-S}g:\#!t"fBA=Z	k.{wXYC'685n<BN2P"2S>W/8ycPJ@_vjK{l>*Ry@>	^k=fu"m2p&0I?6aQP6.=Gyjp$$W^zgI@pSpC<a+c(	26B v8t@FuKv-	;Z*sf/JJMQxZ?*
~TmT=y#rD[kE>\IXZP,!C;u^^pP `a9%4hc]&26hK77]ePAK/wWxFQ#Vk95L*+xbP\6Fn=p
]"AG{6d@h?0)P1'hOY.OH{(:t	%~Ts/PP"*
+4G!4q@9\QS`8odnZ\;r4^M>	@:N9(QP V|4{P`V1q/'JX^m#[I_kpa0; OQQ(Fa#Q0xZJhd\LP'3/?^8a;71OYY>k49 Bz%~A #&!|_([B
IHOa-t3wJR%w%J4@NQKTbO?GR/0=z}=h>j	32)2|QDzn}-:qo
~9pv}Q~hk(0I=3\xZ8@#_$Skcp]iW^0,F[b=898QF%pE$q9i>e!}%aFIsyl4ph8p0M:YpPR0-pYLQZ'C+P"5%~y!I'eB[5'COYy:5.rLj*zR=y`d8c<;G_Y&
FBcph$-X07c='Q[C[Y5:bb(?UoMY!/xhk$M	/i
&XVFj21TeB2pBcQ>CX-bCx&[(\au>3NLR+3Qx0=1c%[A-uEU))Ex*	JjOk9y-<*!UuzlnAa'arS4	l0@[Mg(phM)q@#5kC+zq;`51tWStS=`[K#\AB?$M9Xacg{ul240VDK&=x:6La1*"|zj
Kw;f:?T<W^%+?YIM;lcOI1tmBR~t <UK&9jS`doI"{uG<SMI 8f%C@hnrU6K5q9f&*:`	Cv`i~q5jlzC7097Mms1'C05Yy?yd\j:Fb@/a>gi3B
e?)#h]\R,|Xv^A-&d1jsm([@4941 P/tX7}ub46qZ^8p:wqaWDTB4pO8>PeW!bFD^v +ld5#;h/+=_"?8]2x_\]alZ%l'~s='7Ab"U}@gIMd\hTZ%K.>_|bRbUCiQzNO(sHrm9CCo)*1TLf/{+kZ
UmiU$Yt]96Kz@)Sark*BPg*[foHgh"a`xUTrSHrc l.;CiG|}P]bAB&@gm""c6Mkw3dZ5Xq4e^]|[aNXzW<_ZpA:MQ9AzFHH`yzb'?dT5Dym#	GA\v=^M#QHQU\_XCigFk26v~<V&u-jro;]tgo!L_^_=jH@3H
2d<q[`/5 M$O;@e]hu'omfmbcpA-Hb^,y=V8xj[k/\hq&%wL$T+2{UOMCnB=(Rz<%O+m9>^g_S/u6XuiNGWk=|$xB!pr&ID6t~Z
RCg Z7
[A@t=zoeCk;`&QYvbVY
Lj|ND
=r$G$gB!r[b|{FAt[[-afD8xV
rA1Np'sE	`AIjJz5<VZoTDvgIZf5M-m5v>`C|0I`lF
\+SU;V3[.6Op,r{IBA%_@CbY6-M;	Jry_6i1TBtt`e`Ovu"[D'5bMk0*8=5]oZD.BTyI)]MSjub4cbEz\ZybcM/f{hIZ7au#ps~Wq;0@ FY	?/{X-_Ts_BOO./F*haG)=
'v)N^2$>OGYxwJ%BXe:{3oo.?T_X9U!l5aYp&\&C8)k$7Vn
Z>rZji(<"
4Oz_!c9W0O(x:dW5IYI6|MVH6/	LV#~y\Z]7drO)XZ0'5f.Aj[;+3Zj<PW9G(^NIj`D ]S$,/4_cs-7mCz?t\(&NQw1tr;C%"#{h,f{x{x^E-QDP%fpCPEt5<iO]ue[y]_m~	:,ST[$%ZA
g*NL)vmW,P#9~G9[\t]4!v>]l$:{f%n:{'ayew[17.pOSHY'LE!2b&[Qb"^nDzpika>0J|T%*,ko~dTt;VU5{Gg\l'AnX3?"JP9\Jfl}oH};T&KQ
Y)W$`MKCQDoJ!'L^$aFS@DE#iP-_9Y/x-m	s|*7^Q$	s}{KKB~U=Vl'4ZM	O8$<Wr.0SB5aFv8fS]bEG:P)rG{r.7sMHEAc mM4FkD(=89CBfr.AMjCVc$k<5&wEj%*aUQ7OkQp<J~pQ+k*,!`-C,#%X8%Jd$;bAU-Q}z_*Cm>v&#]u'hXK|/$>buURbyp_vn"0O)VZ0D&y5/M^F_ru}Bz]>[aAtvi0QH1d[=6GS_7t<}gJ4#caC=FyzAiGr?oG,V?,XfVxV_F{+J-.a?t&NXlWv*!/=\-a$wyof\o#Y_Jg!ve)(dlldv] DIc[DnV>(lO:,;&(m=/c+?1j2U"d"2H{8ss2RX|	dn-ga0P
:~r"D(:vj\r:cqczY=ajq4;( ":|:ya]|\d9VVkKZ*1H[:*'';6	{kf#)n"EW~@D[A:~muW=sE`//4q*vw;><G)&On^$H5w/yY'+s\%Wmmds[2n>r36e#ENV<M%#PZ{Aaw.<h $	o0Rx	|>{A	?e-zG#?NZ!>IWp)
\'EVpkEsRcd3CjQ4QK?NWpZ.pp5Ng,CX,#7=	1Pf2W`D\-kb]Sd]l::)$Md9nR.SD*	d/>In,Xaln| @P@"3NKR]laO4InqtX`6n(ZzedOw:nRbyn?RVZrKIc$xVl/+:&m}sa`^ G]s%f#^b!wdMO5OH%Z/s{@C<3QaIN:J>y150a|&&^x<m*MHi%@}Y2\"&zf?;, +\Az=>Ima^c,n*o$M|E/pr|wW2Qs.64j^:)t0QKH1_&@n[xN"(2j|Yv/|fL#*SKN#;0xdUJT{CbifkPuu&6%0vYn?^DN'X_5xdKDJ"GCae}(*D>Y$P<1~seNrE&5_zJXR321)g;_o !esyO$[c@Idas[(gYRQ)=mC-Jb
3GGs$YzOIe_?`v6qpZLr7MP?&oLV]:Ar73|<)};s%3Kn)zg,&Y=-jlG5;(QVFO<OZ#ssqT7F`| 2B&'
Cfyee`.!,i,CbA4$we63 L]j%;+[HAgbBH}^qmjGRW\H\?WXP>}oMXG$4I<4jS_H$T\F2+$?Q7XN":GQ_ mqAw}CJAMt0,KS!T2j`5P9CXC;-9G>|aJW<5(,'
c:n!gU8QGtM.wkk+6]8C0Y"XhSH`JC5
+1&LOD'WExl-_c~_)P0}i}#i4vw*n7-~
Q*FjP
yqhq[>BkOh:9	h@><}q^e>JCNC3n-?Sn$2M3Wac;w4"MxPnh:W=v1AlLXq/NOAGUF-i-/]	n!"\=?w7iy*ooOCY-a4;6tv?@Z=^N]Q'2QN^sg'0\^j>61s^NszpwKfR_>m|z@2DaLN!_wd0"MsWz|DuOtnx>RHE	(eTEv7*SO	B1]C^'.+~Y8rrH7"\4qrey6p.JBP6IA)tybza]+W5@:iMLM4k:#WL6iE	NcRJ?>F@d2	;pSUwwqBd."'e'MP&*H*C,DY;D/Y[:RUUg8BN1x9G}?H]1_e'Yc#d`8,y:J"?6SFp|m(aoaxlR<cz2!'>.Nm>q?6U&W?1vr[sx1|c?i2	iioq^~|qn	N68E2x;C"Eb3U%3K/SRFY"z_q`]R.<|N]_|M44mi(D7^
(e/^w"k/1R^'X"ge,oXm#>O3>--c[(or_(pR:B:oR?MXzQ5
[3J{UQ-wWp0e~D,#{htU@3axY{f,_+uy_.klO6o}%;(_*GBn;.QDw\cv	ore$Y}aikPSxYS)|"\fOhV^>jlR4iIllja=#$|+p9!p-5O!bm,6+Q3*!>H%	0{sswjL>0nA(Ohq&pC5I~Y>e[<WO6rMD#Z9MhT%%)+K>Sbp,C,_1,qED!HV J.Mv_}+0|D9[q{n+\cP=Z%GP(IR8:mJG(P&PS0"xn=z(@:a#M`4("K_@lwMksHr)6&xuSCe3tp%$Y>5$8V'/An7gqKN"8F=q.j_1M;F\yM\ziNxpN,wW3)Si0)M5r083}U!el%2;-v=]j$C<c_ROf${RODfnPvF(&ZFNH	>R2wI]UhJ&XGs>e'6i$!$mkZgr5s5Q,Pv9'	(,g=M#nwa`3A8/IlJdn@AVb=!f15hcb8}ci~4}I] nbICA40i_F;>0M}&"P/t.5'`ol1(SL1?4Bu9\Q$~PlqVi<-5gvD&%I-6dXEzu=bF#U$@X850l}QQSX*k,&J5#_@<IBw+utw81`*#Zz0tcUdaIn+iQ37Ur3mO|c%AzLmd|XZUPsODO7E1c1
vu}J@bST?0U+dZNd[f1cP&8NF\$ophne%G.ph)Ga`_|gs,B*w,CftV[R;+sV,lB'M$\$K/w/E@GPc]4DFUT)o&|jp!l72XTXE00]6iB4
]:Y&|u$DT|<7sEI;^Sm#Ei`+*?K#(+T$bbN LD2[.'t9kaVadF{r_SS	y"]hQz
14"4vJ'7_"s.00i9sl8dc)U|Q|dMW9&bM-}cv:AXosu>dVeY12\ "n?G`VFs}UqDCey)R}O#6AiOTxIta3C6!i#KKG}Lsj^BHD35I20H=/"lQr?J7V\XKAN/2UkPXeg@hAmOBc(TLZ%T}&Xj*Zw]W%||L1xLS6">e<xO
ApYI	?(3@K7zyJRkFez1.cc*tdV\3g}@)[Q4uS=rwP_PM_MP.u3.Ol+rZC5#@L^JP*OIDi,0 `A]9*l\Ed>FQC\`BLqdS0:\HT-H08LccuK|=91'*a`GArj2=sF[cfj@m",>*`Om*N+^?'F;x:@UeciO:qRc$=6n@:a@rVifuHc}'t`mTonTT8pyQQ<T)<,qH-V=~AUO">	>'& 8qn#P[4wN^hC#f?UY,]$SpW+4CMi$+.7vl2Ta],&etGjh,!S2If/2+	`CT)V)mGpVzDlo)ul[}pRu7skLu`X<?kj94=8DA*Gv6XnTwDH*l.};x7Y&j[? pi]@PH2<h1j -Ye;fXQbU?jT:c2ll"v*&iRAYC/nn:=.2F$*j$Vvb}9+bUcbg}"d^pz]2C:+	6)v/m2@=A':l4UCq%
]T&gAq*{RVgtc!88]u)4Yn[wArX+\|!_CJr#_'}L;Vz	xfVk12W/;Dk;OrB]#t>"%.jSaq/uov-x|PFcKF$Sjs`,
HfUpdk
l+q9CEQJKA7MGe}pQ0v*|^4&YVQC\LQ<{,M|':C2J5`Nq2.Mt.`N's3z[C}\*g@;#+]rLKc{$oZW4}Q7_CpK!;`.APBH*m&^\LfHOpg2Q/{Sy /)=6'+01FjS|_`1!|oJ`e6EukFvtG;"KK\2hlp"/3>ROvarajTJR	{$H]fL"AM`wxsKpn
hTE~:.4fP{9eAtF;IVg
(>U3C<S:Gd'go,GoZC]LMn`8(KE~"[2JDl;U8c 8}d;9{?_B*1?chn C=LFojtUT
&Z!@2TX'8#@'0EKvGP[o&"vH<\BK^/2B^"K	k}[|cC6Skf8BlR"n8vra#zQ+d+2&cX8T%D4&,,RP^,98_W~ >	4#udX(.W7"mK76`t-0k\zSh
qC?v<&-Pk9Lk~y|GP+-zI1,:XZvNC?pcPK*my5PFl|jb[^D^iOjF:(F[)PPOTlaI%/C1qabdMdKH( .)RVw>JdKPE{QVlm%b}A?kb"UHT@MG&,lFNCb2ZEDP]r=UF3Hq;	iz[M.Oa`v3_]@<+s?>&+c.cn	3/#)+A{~1cxJ>`;K&ok#6fI,gP]<=by'_<!+e3o'MwSD@,aL9Is3x%FrZ]it=
1vJVN<K`2?QA(~ySpVB+?z1X~;"mB5x#%lzMLg(V,Q9WrLg5{b)Ex5{YY	86d@kMr<)Zi,zQH>g^$$*`nl:7> QlO[td	jQFA8bYuNs@:cXnr*<t3P5/=NzcW;1:]
lA@<+X$F:iioL*|p4*7I<A|9LR:rC	A[oth3m;)Zc2nDS<V`#z
?",k\{-5DSCPPEIs9t'J[Dl-iEwk}|QndsZiE9Q`I`1,~CBb>6|U6Fw7Oh7@^xU	&pe#%1wwZ1LL&_%T*N#&{>EG9<d;{I7P5($dMN^q%|`29#11;txX0V`b"5d;TrYuL9x+	fvf,3@$9LN,rcX%GoiZRk7sN;N^390r'2A
"S*:!M94L;%=Gegjy"9a-|Ns	F]4B?3zGA[)NTk~D5)pU7<pyL[1`x'\@oH7M4'$ YZ1)6/WdV?
dw_WyjZZ.HDXE24=wrWww=1^"G9Voh%3`%Qx 
_&?w TUP!>VYHa-PDq:I&RJenT/7p
e,&#/2QNM0#wTOgXjrk/!YqG:`0?I_,C/SU7=n-p2k51VkRDU#	NKPv`#?n".6T?P^YIniyjWkykTq	SAaSV8lOq.hu:aA[QkIqv'L6(m)6.s4k*pN{)*Fw%Qc>SFj|8f%xwPni?ahPDJpN~bPA	dm+XL^
XnCLpk![&A[ew;/;2RZT*evgrN*k8\|G^%
B9y	],wgH*guN#.feBq=#C9BQV:iR\MD4{<jN	Gn7<MSN Q|*btNpB(r2r(
.ePW)'E5
|T#AOpL;vUF(v0Kj&f%=8l?GRJ]M9jY<[>HC>pwAx!#r&A~"mf2|,>}1}HvVgwP_ LK\"3rq#smWYPKn;e1)60q*UXzfv\CK^5JRYW+@T\gQs3))s=m0:R~2<>;;0XSSOyu(&@d3,gC[ sp<4Njcb_o;f>1&fW(I/u0T#S5+PEsJq`Kk"7R@g$a[tCAv
}>CKPabz)xquGw[n56s	_"q &BP<*hcyfp!He($[8~Z+E	2J!Xu`|y'@_(6sxNG. cc;Y?!-GeUs5}LZ<1@E.DQtE'I8G!RKDdC]O!4SuNFu&!dQWj#$d|sJ@`,,i.JYnX@]bL#c%m#&ZGjC#m[/{Rl=v`a8ZUq0Cu0b2n.Oi>UIC	mn,d2}N=bOfU=x~E/J_9*s Ls3pFJHCPTJ?0#{!vDF9<h"1\tAC&D?{s.vlZME9ULg:x)ZzfBB<(ngKJr|5vY'U4u	Eu>"Iim@tRW5?c|:#C5x+Y/r;wi.p#|92Hz`Ki.)t.?}V8#oyq=swisEwBy)kMYH(	#MX)XAR.<cFq #Cl_)I)Kz{?`OTS5sh@R!c=&Lw1SKNU;l@ltL^J*C9!M4shQycTC8;u?Mm@}MfN@tiF%`mO4ybKB$z%r~@2=5Oe`k:W Ga	Z<]]5gZ=xP?>w=yp*N26.>a:%`*Znx)09}dnU,1??0[[fxr)V"'BW^Ql.k[%|iWv"N{.W|$otk0K`IcIM>7*kk4aqOKZ;<2^j2(?ie&~uS2l"Nc8Vqe2>S4L\8gs32v/hc-Sicz+U.iR(_z:$M%T8Bg`j}u7|f]aR>}9:Xmge^''E6h)|=	5'q@oG>lsg!KP0/mEU6]i6/Eezzb(oXt/2c^[i$C3>W(oN=G
lI-p2]$Xk)-zaa5XAr0-=ch/0{e@??'nM<~yc!%bb%cUc^N[3[eaHAE0JsjoQjR)L<}	CD~OFIChR(Xm|.3ee5Z\2~60+hEa78/$dM1n"yfJ #e(qd^Q_"BMA8VrI0,K{_b-Tz':	*&?]i!4E(xlH`5'RfKZ6EGghE[qn0
3nK4C7@`:}3NXH39o:Ii<-_H![+c].%ZkZrG5f`^.fG'e->pH>S7C
>@|nVH;\,IyF|)$:`_ZvC~x(r=Ul&aQQ}R(t ]IEggM`f>#HOvLiUKN|=hm$RmB{:{"_OU}<	@;I]65](_~bh.ie{vD<,k"6L	(w<rG6F<%d[oejI5[>FH||}o-L2Rt_>QR^=Y	s}Yne:Dk60p	.(=,/|Gr_v/gO]]bXuJ
!q:$T@K<YoUHy\Y,m3QLKX[h5"xkuS:2\}5EU]GOWX-N,?.3v4aOm[w3n?&x.n#P1kEnq%~dL
r/R,j2Ibk	+NZRL{6Mn#x#C,Q;8M47Fo1glkdc,;&}M:M)?k@)TQM:ri0ZOPm!_eO
sj'1.A@I~@&4F7Yyvh$;Xyo~>+x(7o s}6GN/sKh%MZU:gI7yc`1*rj|MMTOa\8pN^,g4o[wQK&uaVZO36Zv`AC<=G;Tpmxy !;rO5&O	2eEt7w4jdr|vjk@.TZUnu)QC>GQJ_e<T{RUwW/~Qr$$vuhxo%fP"z@c\D@Ho[?_'1{-Lk[u_mZpgU,r}?l,Nw3;Yifxp6f9uz[immF%ea/orK"thsIYKKpH,%%ltj+$dH[lK-Q22mh6@sVWp h?{M5t>Pb?K4{[-U1PQ5^7.-Gj>Aqz?~RG*7?f^v/'XR*!VkPvn5`'Y.6|Y@Mr7Xd7jgeH"[%R)r@!ucnE-,plcx`^/&UY$Zz;Yh#-*u=m]
Woz1iX)ta`9[1}hDR	_C$Z319Qd/Q]X9"tf%vlAO5Fo=<;E-;AD2F7iL1wtb4:S#0jid6519luY{'?a\}j_h:FGv;32;s gV%ZHR5e2`5
}cp#iDODj'%]GV3.a\^L.C<9v1,EBvX>c=Ex1b=m8/D+ ?*{/%$fI@K<m6@,KQn$$<mQXk-Z	N^.NYNKabi.3E3nlv1	fZ6`{HYLE<Iuwe="G%4=;$JW96/i >>_ n0*uxzSKDAsZ$QHA$RB & A4$`%A(DTpsi$\e]/r,)B'~u}v`!Sy>4uG%[4Ow)z> US-9Fu=L3%69}$bLs+63;gYCK:<mL;XB*(w
-E8wcZla:]5	i#Q;Px4,<o/&D+61~Ym6vEY.wb%gQzZfBr<P*[02<zNQtNO'J4c6Y:<7,zx"TxS2S"h|\(K^<oNU%LG|JJ]Dl	aj83BRu1fgJ[[a#:FX[O51@|[xOZy:.@6rWq^rV)
<$E)FAgDt,RH*o,Ic	
XQ'1qRCF+AK-+@}Ripa9z(btBf5 Sn)oUrC"ixr`c$FBEOx/2Iulv:6tXnPw`d!;LhQEqpo&pa=/<S"w0|r0dH#~8^O2>[f=/q]~\]'/%A\d/>'k3o8YM.!g1b!_g,~
$YhUYPaJUHw4/%(b{4D#'qP0#c!F4zpS&?`*QX@c#-j u;!|}hD8K	xmY!{bh+Vz:f*ddj~vV_5p`]aWh5Ob8//#h4S+\anu]{%eVm2S'U95~Rd0mU`9HlHHzD#:.koza[ZnE{U`o%PZgXf];:d=c3[jC-Q[cth[|d5_
$6\+b$`LV)N?*q{{m]4;(0c907*qQk/9*/UEBGdQ08Rfno*jzY	idkxCw}.%5\LvzogjKF8;1DRkYS(-YT&f)	MvG#$No/*_rXYq' R[6/{,upE+B?t`uMr)/`(?B|MZT/=&+U=1SF&%E^jvi.(L}*b4J	7"3|
Si/W%T)4k-P/J{x@W:Un	@3}b,4B5!fO&eyqt']:nxy*R+M`Wn8%]Up!hS?TrUNmQ80+JAf2(sYT5QTi#{(Y:I'pT!vo$#{~t@ZMvPo\NAxU{i(.@[z00)NS-Y74JlZu*/1#!P%cO47gGYR6B1DB@o|
|09WhpmmOw,BbX8;AE@*hz^Qw$6/#61lZWy!=q0;t.d	Hs9._(}6+<9^(r\}@1Vpe&>jR)Ct.85"wgZw-';OSEBjCKA9$LH5!fbi)k
L^'_MwG\v[jlo $d+OWux<Z[f\?pBm(=VgOgws"Z
=tq@%Gnd{vh	8f|TS{3p<:vR}Sp>$$4VY /H!	#nADQr1F["mfSAdW~4"Y^[nM4)XPD2)O"O6\uZKR$40fODtZ
psqV><a$(7=AN&pl}#bz&fJHzJ=e0#AH&9~M;K`lH28
@4Mvx#_^0yBYxi_"lh
oJQ%v^hfTdM71irLO+)uDnOq"C2nL/L}'OoVI59_c;Tnd$yT	;Fni70_1FP'&W?K!pFbvRBF01PW;i3rF\27qNk0N+~%j	i(;9~:y!fxEi[ zdJZy 	Q##J	FrI)J{@"eqN'Za=1dt zu7QlOW4o7&EL
r!Kft_r)#,T0<
\z+`5%1s^bKpI#!w:z>2-.RJq.&fmVQS&c*E>_]^P$TO.MI=zB
TGqlKJ<K9PL$#WIW*@sji-'r'}(p3^Kp!>V2w6a
idn`16a*6]@,D:mj0,d$ReW1</);.-\"A5%|vhC~#=\<f~4q#{AA>X%i46eVfC57TAbCJnq[\Ade;``7K|A9	"|pKsVASYl<C&6q=3R.9,Z4([1/?VY}SRp79+'BrHK\~AsKv1\j+lQS.TdT0](@DF_wzXX1==QNs>yO.{}it,gxd)m? tM"x'&.O:Ah&fmjF1tCgud'Vs8\IHTRNr`7VI[g<Y!`T9s5:&-n>x4Gup@y
LZ}rU=n!X$mWl}|/c<DzeMQ5)RE3"4i@'Y%\	bLZm<IU*3LYW3O[.ZO`))USvM@tp8q>Y`J}uEkvH2>mf,,<=Ga!Z.e|x4 ?#e|H)M]+eweW@;|+W>|}k43
^AXXny|Ou'_'XK[t	$lg.N03pl]cT%B`?k4)t>~PbwD:R/FYh5.FQgrs{O__phpd-ui+$zGrd7=QzkP~grh`J664vT}15`bm	wq03g(	^O)!Hw:n\H o(<YXXN2n!2^i:j(7{k#`vq=o1:t-h-(PmQq!Y[=0a g|`pPEB$CX/QP?zJ##eAu(Y~qU.kf,Ip4r 
~o0{W7WigP	El:FmQcM(i.xM u@"94N>Yq>TOG8ckubzhJty'*IqX`xnY|~i	R*JN
rP@ajxqO8*\BK	3C)&2O5r=~9^C>)=5WK	7L06`JAbAwsY>ddP1Y@-,xD27$-),EzF--[uKl996Y1,BrTVs]WQF~iB1d{m#w*eSMxH,':YBY,	INy{%h/("C6&]xf?GF-A'zx;NL/)<Qq	R7>=AI#db(\xxS9v[%Rw'e l\s/F98r1>X}6(O-42I2e!Ypy%(DZE([l50MK<!FvAv!(j+,YV5WpR}?)h}Y&KPC~BanyrR/?`FxQL=K3`2M-(PUI:XNDYcO}i
+T6BIO|	}pd(N96J>i<]\_)(_-E@$0:*,^2--F71\c8xP{CEw3."S)FCa`KAm?#v$U#;,z\#dU*N$JH"}?o{lN'/mGP.uQZv+hn6kIdKbk1}!PG.Nq<B*\m18:e
	rcB5rb?~#,GV`!>FDMQX+cx]58Gx<9k5 1MAOK<c0o_/|\0k H04}2S9LvwSS?`DRInP(!WCcp7P2Aw[jr?;-pr5oJ?CaGc){<+]/
=,qW-|Ymok~_3>H;x=@b=cSsm6/nvvDezDM=xH@kZ'ohW<Z&p"HHjNWK.o4^!0</HPChd=;Q`<d~ eZwF%	%mm/{8xb6:1
.#/fR;*=1OT]>. aA`*PsUN,v.ZdNG+-cP/(tjrSD8r$ku{I*	FD	Ft;)%('mq"b8qkQdf(b1B'*QMli<d*qa8-dga#
IH0q:r6je\zeUzB?vecc|0C#:<w]M%CLw@IRCX5O1O;#_+e~WXsgY6/g7Iea_PU<!-!?vLS?6ba03 \bZ,]uOs9)oR0Sz;	!r2K!fk>-X.9P=YT~qjlybCYeXVMqG|RXIr4B}{vFKT]#CEt<!w\Tm(p_cMk!;ZF64K!w^7Bk_ Fd>rv"i7B)	8f>P}RS1(\oJ""8FTwm)MO}.ZudDT5Ti^N9M.$]ite4sw|[,l%I*|'(IQVSpjG/lza!/|-hn&k1}
Q6ZZ!%]a@az}GX"?ocOmzoi<M]b%AHL2P0UI^Vg|DUrxtmB_r2[2Juj}!,<+6-vg5H:Qhi4%x><cy(rZQdQ0z}w#	NT[:((h74b%*3O=<[.8*R>oJY#0FN*<f+";g=U&(^Jp%Pv2a6bFHSvaN$7~T"Z48'|h/vN	}*[5+mr}_KCU$iVVa$.pz>|,uO0eKP,)v|zyz5'uv<8Y@=HH^G2u|z5B$Y)/05$cDfVFC"XtG}^{#ZyLvH7`_%k	MX\+A%-Qz``Cu{CR4REB.,/O`"]Qgd|]B&vAkFi7(}awzcJ`	pI>pcRv2  t@b0'l|'>a'5w_C=@Nkkx}DiGj@)BDN>yZ7_5YxP{Y!oAzDOvm4W}m BNR>dX\TXY-w	W2+d^%^2DdjHlBD0+AhNTXtvDD^P>GtQm8!@(XSK-j&'y=fkpL3x\!ij<
!Tc~Sl\MnY*1x3=X8@`-R+`7n)#sQ!Cr':g)Iz)Kb}K,j'+<tc qFap`8v[RXS\=Pds=Wr#D'K11&7#jbWjdTO:0!%=
(/mT4LXw"s;{hxFS)Iu?EP@m>/Tu.p[\n$eZ !0ykdG8qef-dyvtO4%YpwTa]&4r<U`v%35a^eHf@@9X]hbAxx5}0/kFp9F&V,KU>(	ZHT&tNnd~.B(1U6Qx\c:QdKel/TX
G$$hB$N
&17-,wjA9FcY\YVu 3 nM`bk_.|Nv*:FUMkz"9S,onAv,rtXC<RpjyNJc{5B-"{(MkAO\OTY :d_58.@*Yy\9 Cat}*VJH_B+OnF:G~>37=!bV
i80\E[gN`6/DajAD*Tsh7Ck`a/C~z!wUlhL	8
nh,,|+24U_:=n-bU)FrJ0{p@(A8Yt|*1+8]5o,i]OZ5YM"Oo\+(c X[l.Zo:0,v E"'HTtVJFsz!oa'v(`=H}mM__4Gr)]P*?9	([Tk<6JroG_R|lx^AGD<*^ Hf'b}(U-U5ueR2
7d#ubm#M_~C4rN,MV!)R$i48[XhN@!x{x!gT0F%|qf%VXL_)(	&zq?Z[Ju13boN|5n#C>.nB#[M^#Q*Ni@cg(qZ
IabBv?Gk!/UAF1XG;@x,vU[v$!ztOU^J2mXoJNS}hZ|AP<fJYv62DJ{8a)M1 qyP5tQ1Y#ynAXdBc#_Y@^{rX_-+=fb$1Oh(Fh8Wi:mT%
9?V]oH)L	#C##;nY|Z&u&,9Y''Znr%k
n`*:}gZb#0`T::.qei,2|4 '
0t6<Nxsi4}nDx9'(]@
`*rE
8,r]}\5D^;&S}%U7DdIt+Hxg)3l@P!bU'?#hG^WnXs<jU?xx8.%Z%dc!:zn.Izj20zK{"7=)8tm&g8Dx,1vZcT_'Z#RV;s_ME
`1^(P<F25Z^	LJ)[ v*u	?L-uD<0[J3t)o5S2^N~;8D%v'8P4ZHDbT$_*md?$#=7&\K(RGPEpVlr_2\S\ur0	Mk';ifgDs\4e6+D{{1$e:y50]%#vD--,P4Py0KU}uCERp'u;h4Pkqn}K>'xvAzV*0Y:-"-k!AcJLT9xoZp-vLfnA#EAaK`+>t<[;}At_(RU(.^Oe\0gpUH< e)p)&mXqw9\<wW,]fbg.Sz6#ADw4Gz1}y:NB\_$
]oMj~RZNx@O;T}0BLT)U>"S\ jIvCgm{FAE?-=KxRv
QLK?`;r~b:U~a&f"*)cOBA.F=^bs`='hf_pUk!@)#JP,{3,&[(YXX:;^Ke#wSSc<NcEgRRR-+v*4~OXK]CmC5vw=
k:8S;Sj{~'X5SF;89mJi0LsUN	xVAee?d!GP\(I%3b){6k>L&6"b~d9NK>z#y\,o&^OX#Q-6Ds:C"QWMZEr`XukH$UusdQ~k1(7lF>[%}~32c2m6c6nOX!~E^IO.g6}]'Q_=fohKz>`-Ub17&|GAGqVQ9vZJG;}o0S:RO059%GaeNJ6@(AU;m^ROYympd56 /).M"@	snB_f&ie1rOY\hRv6m#QmaN0Hk`7M7B)@pIx9(xlxW4){rD0&i_GzYXR:v5I/h!%QCQPywB>hL Gim-2zs	n|AH?74RJEjTC&B7?bqMhS2{1UMB~!?G=	M\W3@cG6K^%O\bn3]5Qv${.E;{Tbt8oA>%XJq"^9Onw}-?GXbJ/pwlaoHu4&JXG%vl7?t+X.D|9sAE(ri<9z&h1<9s-\"7L/_f"~jQFzOeurON_^^L0H)!;.bq)CMff:xA&E619:'
4Ec<NGm3*qi#9/acAg-$:3|LoCdox5:w$<<0_x3PsS.+'ysZE_KbUvGu}O
9noTUbIojGY4NXq*1tnd?l=vqz{ojd6~IyXSd^O!\].&Yr3=C''221Xwbxx>W9ZGmI"NA(.G<z?!*'ZsYi]sV9|<Gb+l(hcu#dTcAIudEX&1,>3{+P<DE|4\bq=DjWkRi[	yUCW^@v,#!VE}6?VAMD5WeN4GKig#$jS3#W'?0[G/=U/)t!)8:f~UBnWa<y|XY;@Nm}xbrs'Wotae3QgFR/F6IVm7S>F_<oBS3C"\53COcmWDw A6BL9oj;DDT<\X`I=8&?,,TW~WIH,<$_BsR++rj@04M2]gD"VGCiEUKxi,F(>Z%qT%Au$fLZxOEELw>x]5b9QM#_8x(_b{PlUO4@C{g-	O$hZJ^'{{w	6"T72=lUi1$a-t/ML+erL'Bigf,TD}5Ovp.r4g9hPc<W_\tfmFVz+p('gXc-`zWB|xdo:iP58@	*SGdYHKf}J|TJn!1
@M(dH@L2$;5LpN(.e:+KJk6v&bY[>
RnvR-dz<TK8Y3hwlWlN//_;nhGahryyMY`0z)K%s*
9`o9@nYE?fro?hP;jX!w@qN@F{
c$uOf.@5KEg#cUFuzwj&3H|RX$^Lx'L7Ix&m#LGR0@[<,z*WoN(yF5*zKY}Gkb3H_5fc'=7oz)8#bK{0|/dofvk43ZKH"oIM	
@QdT<P*#77~^4Qw5O9,O|y+x?uK <@Hm(qo+ZlC/ooB lv23A:3_a"e!$frGZ@4P2y\9~g/;?Kf1h+e7d@~HlFH#x@HJgt]K }z0eiWij|W	j\GOMOK&y+IwnyP?3\)p]dl8xFc<]m@C'MG!bXKDG:S~0,1?Ehlc:P
>&|4tyvGan8a-FNdZ)8uz!{VfCU&"<u)L t'vDt$p- /	f':<n<a/?x;iN#=J|e\("N6:B
A
zgse"DlXG=ou/GW(*Zl&.Bf5DBDp]jU]F0T360BHD.C5]&Y]{ Rjo?d#{?X'pL3
/P*4eUvmblbXnPrbE)ct3$kd,1)k\IP/eCEF$1vtK*dR/b:2?]*z(.DE)U;/NtB_(|G87W4g0hSF]=WH:{@ZlrG*eM"<
+(RF|?aMmEv~I%O7,%$H&AaNA@0]Q
&5L}
4Qe	[B1Mo{ W\!LQ(Z(?0EX[n.'|)*	)d`|h_#FhgO7'`ll-C.2_j$9L^baSEe*=k{HnxtgJ$W?^7J_o7(jl!oklQ=#'T:o^gl[H/%7I"-&:	QjDU^U%S3/ce@}Ez?(B`fyXxS/ZA7n C~(coJc&?t8gMDH&_/(-LECKdPI7X_G()}q(I|7h*b}uG]fWQ
=%qJ)Xfi?@=aA
vSC3v^^SzCN|']_\d0n)b+?		"]mX/fPX+^)k_4,A+>|UD!#S>OeNC)(|@mH]RJ1eSHdhw%|+Qz7]q8]Svx[(w"DpnCCZjaAg@>~MN@4@a^%v}7zuO%J/aD,q_t"gS]_~4S+$$BV8*)turw}uy/QhV1Km#Jbxy5G"jhRJ7:!7O7~o?u@*&QgC*	JGXQ6/.BNg@51Xb%^vWi_gjl9f*iO,a/Q^Qa qn[;$%1C["xez0=p.j$Iv`AmVd_oS%6y+3imxyH`^ReGK3"qV\-f4,,u8aC$_7$eRWnC	z=:\hc*%dd_`qy0,}d[Gj>.&1Lha@dXP'Gq`}RqL>s]p{qzj++_.	:eDy\/^-v=>x#j.Yul'3/	"bn+qcf)%A.IY>7qoXYleiSOPdJPMn%\lsX\ngV"D8&M1RrOB33xGUun}H'	R%M"1fR]tAP;j-beFO$g`,pr<gt]>Z@7TAcu%/O|bYPWB.w5SYyH>3I7jVlKj9GrmS|G
Z"1<4Rul
4y&fz]e&qsH0
([(m k'ZHzCO[ilzbmp;>"Hl{Pezj5< ;j5uys21x5on{NT"xTgE80#"#'J@CJ	7zeN^a!CA@3t{DkF	E8ws7F@nL)|;)DZ($`H5Q3st-I?L7a?z5G6,%%!ie{}QBF^4@mHFbmX@)PcBNw&zM1D)vtEC2^07Rt)#I'kz7kl[m9? MjBas#+(mvO{Z5D@5quhFWp(nBy/mE9#%nq8iOl?'N	o@[]J;eF&@Zn)ToU@lxL#WGH/xYYhx*`7z9c+3q
gnjP(SblJ7nd,-8{%@h%Wb]^mi&1,Z!G'r1H7lX0~KR&$&n6%g^73"D.CqqR4:E/>BpcD/*KB%A_U*JW U?	NaW4nS	3tL]NY|8gTei0Cj'uZ<<&k
QUj)'&fJ8g~!f
w ~!8^e*`+JH|W5i5$(@jD]MlL1`>aV<`um 'd4ZRKFNA*/Xm0\9z;-2Ry>oVS,pfXrqgXi`ydL#c$=*FkRGP,#q;n/_2@)tQi(c'"xX
CK$g _nsQIX60ik~z|CIkBE|]s>2G3deIz08cRS~YIgjoB@j91cXJUu]I%.q<?i,Hj&U&/$t}{-Q%r#ht|g]4nS2CGIwzpVS$fEc;wv=f@sIldb`<5=!GJ?`<oY}/lz/q1qYxNHtzJ8D?WP%Z(6'-~97~+lynt;V8>+\ae76\fY[ D:!a{Zr$as`TJ1#g#r|	6Q&c9pe"S(~L`gt\)JNJ7Pt}?OauI$-UmL<h/jlM`3DEjyx'z69byZW7odnm~{`nkjx5>_K;x'<C~[m,HA22:&xcJB*wc<@)OA.%&0Q0q1bBOfv7i-?JCYw%&p>.<=[Ll~rf[|>T1iq~Su9gM,~[,_yJ]#QS} W}Ia9C{T1Pv21|f-$Rab"VX=e7qx8z.Dn8cGCL!/d6?Bl>N;:LehI4>R~G6dm7xJPJGpT3NB #|v[/n&8m>Ydt41Gv31>h3J2=oLEkFKM'{ZGb4gH6gveClQ?MaRt>B{S}HM:IV?}f9A|F{u39904m1k{-WM8h6q>%{"`&2qn=t^#5-q@M9ZGHU>\V.k#*o^'Q@I/oToj%tndmHT)IdqE65H\1QX7`5N=nn-o3M5Q"K\8DDc)!>IWNH-wg~p|7S28Gr>en'NAmID?\y\4O&\}N:]JX2t	MH3?iB8va+4\vteh%n_W:R# (YD`DM8z:[xAO_Ty	gw }07\PQfE:GU?g[_6l iBCWQGX8_b77lPdmj_Nz:x426u[0NPx,'wHiVlamQU5aHnqXr2(8H@	]2T'-<Vlh31"M'w$I(<00O:6RJ.?a{[tQHE	cVrn8kzF~4",~b<FDq~E"NdS{QW$@:oSKfr?p +]5jO$6'6LLnr,2[
d54V*1JtEfkkG^l>;R2
k."cTXWaRz"5SjEl+Y$1;$cH`?b>&dw/nJ(}OKNBFZ9I^)/?
b4^*]/&xR"v`.traHNGn69xh6Jbx'sWHc7Jiw 07BTp@{nx]|eYinn<3lKl]GS`WK7Q~n`f.F:4\f)6AKZ9"VJu\\B5@3=O.$hN*dae(zcyaa3h(PGk4%lFNaUxjl]UCe|p|D
q9#%yXp!6/z.RJ/k:TQX`/tMQo2)UDkMz+^J'/@A0	LQ]UFr+57}h%)[h>-{C!NXaK\uq#I2SHWy0(gsPoI@TX[\GC}F$/|v1yR2FU#CI]HlO(b3Wsm;?ab%	/t;m0k_|rt=:}:a//$	C)pxf[$O)j|bbHJh|X"MJ%j0S'!dAbv!U6 WlV1!"xQ#?Xic2 )F:5P`ipasCR2RfAHg("gy*\HX!&t:j5qEh?CnjDsk`*'\+M/< {<&!KiDG?]PXb>1gf*Hm?[/=GZBgpL()!fBYjG2emQ<$w*Uy:tM#k=.au"("PE{fj7w_4;CmVKi:LH.]]	dB_I*NU*zcA|[
_x7O.(%2ujENzj)m`,7 O+q<Mrs=%=Y7>l!RE[7lTbE8t	5sjm~v5Wn+p;8*2l+{g;%K-B<:0bY/8|M;EzTBSZawx4]>6Y!RY	9t40|#MpOmx0m\t8>}3I/z0l\Oh;S#A-0DY%P[Pi`(;6!qf.+qT61HwRHg@m}xIxR*Zn})WRI6{6!
/V2oHTiL#ee@JR 0PM8cY|Xy&GK^excrz45m!StBE]Pbz4E{.fhK8ES8>hL]:go.[)?
~E$AC1@vUQW7kD[	F{:Ffr%`yRv(/K>z0$]bIkQL!A.6i#G2a4G>vNSexXYGc(dVv>gjoQH4$syDG-\KT\ry**98g5+"q.}S=?X1oK7/{1\62[MS,M1K,05C3X=6)\Taf<xjH%f?8T
C{fqmjf{B8a!Gl.,3(9vw)ZU4[6}V ]$`I|f/?_G;`q-{74tK[`j5Zll*l3sUY),>~whY:SckfE,mNJnc&SY|?7lvA@k%?[:{}=$-D0&u!#ya3@L*b! o"wp*`4Z.YT>r9E'G`$-2KGGP#qkz;EHuV&MX2V|%p`L|zqoWk](j4R3kS5u<G*yii:qfl2B:^w	>+9{A= dWa8|N(,2CggESm0Ius&E%JAlh1pz!"@b]$Z/B!xD**|>@oM)W.A9q%!@kNI5&EIR*R%7`)PI)gz<Dw%#K<0&@:]I(N354Yg)DWouN=ukg7}/ic{Tz(;V?t:: h
KwK'j,
B;%+	mo"{qZsO'Dwz xHF#
8x$sgL<^n]q$.%79IwlsX^Y{@5q&Ea6ut_Vi\+ym?\	WQJH2@x{r\8Hff.Lqh;9:EBM}\E?"Zuht0C:;@X[>!70!>0m=$bXd^.b<ACxjm"g^:*w\N=MS6s{]x&@j4t3'S=~[=$B.8>Z3JIG	q"GnbS7&)E9.hI
@X["}[	k_/spc.x	e#!Oid[c4@%jMbdRHQlNaRN@Q]Rn2Lz%i4*.xOt:\)--Ifa:k94< Dc5\J7x.d]nQ/J -P|5"}h&v4[&_{z@d?S(LkGUq}k|lIP_-]_O~"V
%@fqGxS`jm_ -D1>SO/2?aq"fbP^}ec)Ky>Llso4xoE,fnD"8yY[b<Zrv'6P{J$wh_}x|ba 6aEfy]&,Qfa~_sI60(	~a(>:WnV`N"ieA?0E(-}=7QM~IJE|4^5.YnAZ[;zx-Q(y2bE2=\+"pqhH^/2[S^/l=[] Nd0q=QV`pB+XW|{Ru{)O#iS`/^8wt1/qogb"~V_Fg80/{S]@wY=1N(*R"8Hb%H,3KdZ=[7O3j
nP81@X/=],RtC!^&rV=6O&VJ,B	&.7yg+GupSb	[8ZakHc|mc%E>_2BC!`d3g:69>ZVvFs45p-TkzO>Qq]/xW7#_m]Bh$/MFY~Zo3piu{Wy1%ZO,V)Mr+$6+Ip1^A u|p~4Q	sIx1xi2h3y-)rhS^-OFxGD]<bw!khM{j397)>oa0(r7B'xYV'd_#Jdb}0w{/{54Q[$L`&fEZ[27[nb>Ufc>__-IzYX{\(Vyt=%T Dx>YuUe3+`mU]>0Lwv+2QA}p/h]qUA6CLcA/0G)?>m#IU6a=Tk96([zxH_J;&"2s
PItUjtH
' *#)z<X5qZO`z,N%cjlVn>JE/ijOeR%d6sAMB/0u)jscA`by)+[B`"O7Tkv<LycqXJ4Kw;[:snM
RRJ6~{bdl};u"3x=bxu=Opq|N":/\e;I[MjZE1[Z97`Q285T^v8vE~n"%oC)|"m2WjS9	KqO8ArSOr;[@vWBUurRviv9R3sN:
g@A\JPmm4Q5xbPA{tS[X[K'yA6(`M)`mg`QC^pryp=fP
T4J
C:`o7oTOphWghLBg701k,,'yGsRBAo4.y~L >TAqv(@)Mwro;{l}L+
\uJX.#T`SS:&=wWulPvqD4iR&dzV< :6U	dx)b/_j;Z.w<nyToXA=<e*~f3<XTHt@#4LqrNeIH?^uW9~|3.2`~_{T6;U]A?pN.*9 Y)$L-Jt~#87,w#+\p hP)|:?aKFKw;z<syxtJ>ILZ3t^`0Vl8~G2h;RZ9t$u'W$*p-2=fw7$!PU{C@ttI+4$Q1Rya(c0j~3y%MjFL<eyt0NdR/D;PA 2x1#3PmlC7yX+,9faktZE\6-8El9Rn*a-(U1:bg-L*7H;Wi?Bp~|w2S9\9[K D@/j_4~wpdaEtc'ZUh!Y@rN[sr4&'*$0lKDC X?D@EFN I"!%o^V	&%F)H#Zem\;@K%k5xSw>B^3E(_-mdHcOYf'*r"0q9S#YhoDAnIGn(=GPDy&E>caq0zU%na*H!yg=!QlE:UwPx=z"EElZ8+;WDSWXluM3mT;JfpSgxNVYa[`!B_e8_rS%tH>8`AX{71X^f]z]2I)N3{":l&8=T4CeE,c&M6Tv
+C8O(n/Wj!\lrgO`oSH,dTZKY8'RNX>FbcA&yFf:H:a7V$	V($6WiZQT7Z;CsUo}pp%6O6\$">98Z-NRIc1oBvk	]9Xe<;Upfsg7C$'vBiCR"^p"Q};?o/=4gQFngoh2~wXO^[L_T`p:fzg)PnlIg6@JbspQ^9z~E`Dm4	(Y`z qAYij}/4k+On#uND<''9/^n{[(]>*$\X
$ewDKGHWOe])m/9:7Tqpp.-jrSHfpfa3^_WU@183P1V[	bzJC
h~LM98hGnX6!G:H
92:(_wkll}iJ<K-=X7{(^nVrqv~FZX3B0kX.]'ZS9qFX}W4QS6	f[JB\
2h4	3uX.Wd|=U?a<1bY7ej[vqD_ k8NPiX:ZvX"-*nj<7hy(`{aZTu)dMsr}9k)%v5@|W#tLBjt!fu[ZZqy'"E)2<{mI#tA=+H&j3/(%9$L;~B\e@wIaB?KS[j>wX2TL*P*)\/pB.0y3YkbF~AY&A}y\I.|k0V>^SReTrOBB3Ry1>b's/HpFNO#A]y(<KY?b#-iAK"|WkTy(p'[l"i;95R/koP>QEe4?n%`ygC')Age`Zj
R`?Cx!A@AF`-eN_bQ@\TBt8]Tyw!^%n<59\3w"	<=')Ty19)WbD6
/v4a?ieM,_Sa?tQuX">DI=<Lbjv/}<Fu$AlCT_==0MD`rH>j^}V<}ue_`S\b`;yq?|6A_yX-D3>7k+L-.2amkn
|gl}fHvO{:Z).+	!O}bzSfgzo5Y: TKj6cvy?[Vzv{*ZcX$m	ke(G6;|f
fb\L'Vs}tl9r*`U!xpIvWpsep@3n&.]GN9+`<%s5W	'Hi#C?|PX]{'f`YTp1o[dcd]Vy^sY8qbvp7+UVX\JJEKiPGB
SQAF'BDAe.}}9g@_'EkSM]\+"jg3Z3@hWt\~soSk5%>)K|-BY;*$N^ce(8

&~%o(U	-Nb{l(MCE f6XK_IfLAgk(
}w|F<H9.5U2#pZ5/79#O$&(qg&,N\~8`9ml2dipx.:NT6*	(Mn	b+
r?on*?+(Yu`SIZ8MU[2%^HS7dvzJYA6Jxc`) bqRn}>?I/}sqyjEm;+KX]DT$$ydsCB^=>pN2b~!]WD?-Gr8eWgat3PgMQr252O6v\h%/2%R4u1]I \#s10I1rSqFd!:c]xXUZ!b%zA R
bc2gcz80CVm?QCD/_4~%_t'$6A<lsG0ey?55niHA?fHR&co&S\4hr*V2Xm@:EgvG!A=toYF@
>
AM\*H=#a@W@zs-p]GA9cxMJfoxZ5Mj"]//
AJ[9Hv:y7)K44\;#o,D]tFX*zi?RW-Bnf7wT(xy8A#xw/|VC!	Zhl9U$},2iO`t.b{dZKLs4gZa7phd]JU">zBq@Bxg*a8 y\x!7wk4)j2gr6]LQU$dSsb>Ak\m}w.1#@BCR4N"32
\\^dY0S&_:2>":Ddq%f3I$wm
0H8CY-4`,DC7+`t>&7;D(xoCq4|<dr.}Ce1qmQ/p-sVl:m)rOVj<<DkSyu!%|j)ytq3q$.5|=k8x~V(T{\5&/}I`u&Y}>(6G5szEXl904R+8fJ_fl+PfL$.~bR~4tI"Fn\L\5<gT7*L/bKh))c;2FSj"OY=t1
Iy.=_8HOy/nU:3$&\8S[o2S#XlBL?[9;}>=y`T~.*cm<`^9D,v,v#"Lc5|n@jtF+9\l0l_YUy^#cGLI/Q{f>Lg-'N=ph$@FSyyKTm(v&Bl{7r1Q]PY+a^%i+,r;z9d-Y,}=W{>HHG|HwTuCf<Q5CR[65]`1 _`b}N:?sH/|	^bKr6oIVj{x(0ZHyz'm50+{zQ<(8:Td<t<+u:\m5?34bS_.IuX{mgP~[?k&BLBw@xD]4lNLTSge!|F'k]QHDjP>X8Z!XWH>%5x$"B@LVu^-@)t{s-J7/i{IRPI'55$]kXG8SRpfC|JKU m;_0}kZ^O
&&,"o1-Z"C8!IcAC_%=(aT%jn	dH2mIn|S!S@a^YMuvs0<	a= qf7^7rOHoPgq7$/qH#)n!zWgE @1FCe %!GI.-
KDA.JxeGq1ex@XUMh{<yi?3VJ&^sBSA%PxjDJA_e#c:eK5#DQ~dEz9o~Ew`2~>DuzH,_Xgh&*O}J:tuY9"NGU9W3q(A-{ee?&lGK=z|Zr6L+/>3o\|QMzQ@Hiy*,6a/t(K{+"a2+~I+rLlt]&kKO/j.KC{HPX^t0"=rUut 8!VpmuFH(CvHHFMs0-@Vp,YQd{-;D$2(/3c!/ J>z3_,*C.}9CJPj"1KI{,*h5~(1+kO&r\4M7u $1NFLuWUDl#D@Agiub\.@ic?0+Bl:[1l!:9DgsA@dI3!|? 	M!a KFuDyXWBjuK6K`zCP#P?;95Hx ^1-?he^_R$
96
@Zt	}<	DjStw$4ZPt-@X
~=3L2cV}Tm%_XdXET_UY/Q"mw#_f2,F&!2|J?]W[Bu%?c<tr4
}=*w'p~FM(Z'UJP3H%5;g0=<K-Z6W`B4RauFj7/D5+T:0nhPMWI/s}k1MU%=<^D3X!T*mOENX)VCPM1cw<fkQWOO}:iJ}c2D Kg9xHs@+P}3f0/;Sn!-K.\P}	<=8D!2~M<O@^0.wqhRxv|sx
|,<j!O&HHs0qgY'^HS-}JduwxYwDS_J+pCdPNYr#~[._NUY3u4UDJ1*|xZT1q{F!Cb?geX5T<O	c%pop&K((ND!g
@t$(!8Dv2 L,`sA8:v?_=`|.j B
C;] 
TxSvJyH+Kt{vMdxyE]Md|kuL<\_t~C(r&2"%\WZev.gy$D6-'!j=q>3k0!	LtTM90hl7UUBjcky^Ze!`T-^WK->?f/WR]?sx:q]T#_smz:7lsU8~C0>DulI>%\_FuXT8w=}6XJ> ;%$2* E!Xq3<bb%,qbzF~"V`\^y+?O(BmbL"gEqF_}$&STEcjM&)7t"orXwE=B5wr_m3K9F5,5gyZF-NMe=aQN}Jj%v/`g2?-J.iIE?}g
TZt/GyX@2+k^=5J3McC@EkN0 
7L!RBKg/@J?+	`4X6["sHW@`Q%CFou=V O}*mj-crS*L#NaPcEI5&fw&Tu|^.?~7v\Z
Y!>}R*s9\}|1a_u  %CP6nZ_\m>O=_uzy(ms$zLe%)PMRFx2L$ &e^@.nuk,b2=h4{H3AEI{}MJDym
/%Rf(OIuFt0P7OU9|H%F$o40kwXJOV$4gg!bzMo3Yy2 qAqK_srypac&N@C4E:9W.V#
.)S=,vvY4!U=*!#Uo0%yT)\a*vz-iCY:9>(9
uwwyUPz=d!4Qe@	?bR#I.k56i,K<$?jz~j"op8%h{K}6X"prY{|LD7MV<.$.(HO8Z>4w2z4{19mYs0^|$nXI8NIlK'XdhYgANU`EEG_n5Owk@rBeO{o7k$Ad0\,F#u4WcW+'HfR%m%s)TS)uP$5>.6q>NJM6m~Bu?>:U}k!}&-C=LY<+,02@	Ip}Tx8m1.;b	}E+O~&9+NOB\BX	.>O+'{K{tQ+^%w2Ges`dY>-p	)	z?>D
P$:yxNNbD;f}|GIV;_%t=s\^]ZA.g>bc9npPE
0]<@`DR1rNf_3ka"=Dg4Q(5o@@W'{Y8iW6@ENOGK.#ntMsEu-LcDuO:SKYb6[
Cnb:c*uj<-ElhKzkKP>CYuCMBx$>_HF#I^%b%]q#o68o".i"MOL(KPP03T#NxH}.>TvGAnVd3QbKnQ`
o"}M2"; 	BziiXm3Wsx[Kz.W0@0w<
1no	!*WoD+G"p0m5<9^FU3nZ~B$ZKh3hjVk2IO@lRl|MS!?h%fS~[5zT.A2^KX>qV5 ?myi!>-VP|&>Q4L'k$`d%%
^`x<>Jq=/`X=2l<[l)j=W,`;mdj`'SN7,2eOc!LDa)cm[vO~d/_'ABfYui\OPdch!9Xh='XOC'lj!&<OQa~Iqk-:'e.#
,7Gk$,7(Ep5S>;YuJ{cQVavSkSllSmt{7/U47hw?Djh-k1v[K^$;EhuK"%CISbX;uXOW0PcJ*_]ARgV$9jU=k^w%0BY)7(PHJ6q=O4(NZ'vPw64Vs;gWbbE
&i"x3 IakrQ}A/{`8i?%/["{|1ZWkeOm\`T8~hp.iW[H}Q7!S_u}AAU/y&L_*TTY3K?6@6RV/[W1ic<eLQxkHcEJlJ0#FTOoM/Ob?kef} cUj_u/A0ccoz9SCE!Y'"t/DmyB|W}8_A7]?([6)8:k-B>pXkM%[Ui)MXXL8k1[>rI	q<HeBPxfgX|QB:h,g\2X8oSLrF%Sm-\L76wS!MVsbjI)BV8s~-([i5W]Y)Mx]v+L&XP{G(tr2uW`oKTnzZhnzi_UH|Tr}|Yz/S;9hY!V5`5 ]~v*~/2{Jt1J!qPy'|W@+E]GL)MC2k|
UjIsY3)8oBA%ry@<ghC,VX+}?,J0z[4pI=^J{WkJ'AKgX0`1bf1XN1=+]O,zLn.v4f"eIz_X/6Qd8JWgo8{8I`t(^CqM3_PPXJzF^JWW1v|_Q]RXH*.tPYZ7Vy89s;0s*4#XMNXXae&.Ei>znvu<RjZb+,L?kOj'Ri5>Er6T_5rpP\	`.t18O:Ifu}e5L4[tU6.Q[72#
$x92w7g\]8^{J$O9E\7-]5uTi:"THL`4,}Qw3ujNsH^%N!kN:]<`CLIP%DQMD[%H9ptI1j@X743$"N)n>PQU<Hv|.sPg2wud2!H#o=!\H5ZL>=$
i9	)X-~=n>eIlpB{M2JHop@Q\+0NwJGqfHelDt
@pA{&1?"-GSMETj<YZ3!=>*|/GFk^y0!T)$_DI5BtK<9'tKJz%;0o:d||9wl\H'E\q!]FWsQA yfSDO	'LQ|3h+`IS'C62mR^CEkv\P2goD0t5(}xO22o`%jR&	Tfad8'0(-I]6s\Si
gHLB$On<V*ScMpW})9*U/K!I_1O|M/.k&@=e[YW'TbANJ,`[kH.B[s?%Qa=jMkrdF/SD^Ajq3Q7tS"{AlT'g)uBst?7z1sv958%.[WKb'Q {NDHR^l|phsk"97\N>2'	.3]K1E/YE2zU?]IV@"ZB{u^UOAAi*^b	| jDJ.Ts Uh^]/8;$RQ4VPsTo#luhH7Hd'R.XVp/2hBbP/2&<Gv':yO/*}tuXVc$6nk'_r"U6n9<F38Mt2rV$*ADO0|9]OEH"?QG(ey]
r{X=R,KC&gwY#|e80n$y"!>N~)#>CXE	OCmi${AYKpuq(PVxrBlbE?+elR#,mu\vCRim1866)Q
b4{AZ)UcT|;.w|rnkX?^Qv+-@4F
#z9+s}aR6nr#=1I.|1":hs2*<eUZ/<Y(MhUU_Ml\?e1qoIE.m"Cv`d`3xs.tf2BT(Z4]glt("C|220JRl;b:_99P,'2(a]1 mn7PVl;Sqir{s~#cDWS0`7i~*^0nv%}C='_h^~i..U^nNrAM3NB5ac~MFf{rs1>zrc//'	}y4s=NA>ww@]V&wE7|I;laB|:C+qaPkN4 -@JKCzEokcz"V^d@\Wka=X81at|.j&O9ZIhX*b6Q@"*cJYM7&0D!tL6~o(x;at.L#UC[! ^dFmgL^`.@] Mi,5
<J%S)w;}>Rgw--3jbYtCiw`Sh0y}HV4-"KZz-Ez?T'8Mi$
KqsZ0$3Y
x
Uubb<>
Ii<9&Vef}=FXT|5(bl1:#a8cGPp%e _D[(?[~qv7JrwKXsJ=EZU2yA2bqbf=lm1@lccE~d_m^b0ET/VW|cyUO?ryY=w^1<%58VWNx~2'5G_imMKu'[Up^|+mhhB6-+eN	.;8CBY=z;B}(a&qS?slI2<V:?d5c	8n,{`U^0^D5S/6
~"tth])Txwy_Q8FK|Y)g^/R&Y6-yzjklj)	NJ@MHP3B:Y,nlh8w1>C:EUbsjvB}UEXA_?j16?d'7nj,F;0fu$!Q`\awDZG8EZ`)`J7m08~DXq0 p'^4nbPg`,{1]2:4kt{Vb0Q;Fus	-jBD@V}VCUJ$wK6A!2	G"A->chgv"	EfVS>/r;IH(Z-+^Na%mZ6e;uk1K&z)yKlNtmWgx!i8_"O#"kb+rd
w>o.%?frd=Y+<1fbPc^PeC@l$&_d:4uCs>1j<opIL;e]gZj@iHXgZ)f:mc;CqAH*U2+v9}|T+o!ie0O0NlnX$s%ipqCz2wb[qKG}u&YM/ ,<_=F>p$Rt3(J^w:R4E!,X8/o^6waQCFczhTe+] >c. 4e;n}1X\o-kWn^h?kS6~mx{[OD@R/A1g!z_uTr'z9wONW\'5k>v";<.^R9'~8{M
M{Lgi^P$*\[f5h_NA:W#m4FX}//(Ct?))Rg ziR
|G$C%VV)b471=R)Zv)|iIlbl
$US`0l1kF71}fwwnv*j~f#*1|6:a~$a_~nm28zT!vOl\v@+"t!x"^L-ib_YAo5qMvQ>`?BG"N[:RiafG}k"[T\^r*j*q{@>W&c~`Byvjmx"4$[u+dC8Os0 NlU-*v3BL[=MS{"iy!P}M!?smI?oc'Pox*{)c^4^%y02{T@/Q'#MTD	gj4#ObfW ,mb10F(6pvm{cN`&I+"y'4q~p
GZ~
IhLP9Od?g{lS>/y3<+d#Vq{VH::DC<j`&Io\)mr
YTa\yzYX##~|& e/UMi[!UK}hUyliJ(0Pf^G9nzrqSAK?$-$3cd],N7coJR4Kr\gjPcjFxu,:4J{CWY|4;X%%4,dl9d{m[A|3FUcc(w:X:(/:na#7iG7okFDf0{<Qyu:SPkaChlr"a F)dAX])I>+2WDbaDWKdh.[C_L.DfF\'CF^w~W>myS3Q4/\?M*CC<LNk@@?,J%}FRqjL2e^k}>`oC\Nk[fJ/3|;I$@_c+njGrl!(oPW$#
X2!#R\d3(M"`%/e|ro6Am+)	a1G/pMeqR)~UHz,*u)-0p3M_HAm4GpXDay4XY:3f[K8cYm9%%J`6;\R$+\`LW[i?(h2V)XO?b8_Hl7~:%{RtbV^IU{84gm: aj.3F|A8&i0 9f
JNa]v,i@A$4\+'(Of=$l6(N+/xJIpqKnT-{}6$X%8V)R]-//~j	SD/&9i*cp0Am4oCF0'}p{7.v;puQRp 28e713Fs`/!J84U[+AM"m>3U9>8j#R[F;V*$^V}jy-Lz}urpU,z&KB?*L5zH6oU~@^wGV/_[B+
/LNL@8*p9BU~<A9<gD*G'}#jPT3<&V(2f5HE=XnG{Wk7nkq>5_p('59X3\$[OtCB7*OuKHu<f%V*;K*+X>@k!F5(#qeB2t>l*S)+A#tOh-!V?##e2vW;rV9`txbCG`W-?`X=6n".P[3W BG{WK:n> ]	VlB#&Q& )h,3-C=5brhCFY;%>KQ}Z)</J9^(f`Vtl5>aRm$:r.sRIrF	fl0j5RL'IEc+Z;=gp9h*g7mZ7}ji[X\]u=5Ge&s@xc>9?SrXF	\NEZ_L_GH9OQ8WQ+rFY)YxF{(w<eX2!Nd[2Mnc+Le%pi?Z7#>tn"nn$8FiZ
!q'~a-Y4q:OV-2(+&MddG4Rr;q>qLZr@!j++P@LsX$PIVF9)>$H`(vXb!Pcs?$UDb]AB+A!>NRxro2{h2qu-"!ap+\u$
?6TB.xW.FT!2
>
,E70&;H?t%m;lWj>HkL]8]`K{"M{f}+%ojTIE3AK~TN\^*>*tp3ZOSE%-yw(C@L4B
%{i{5of?&~eL\'dMyLi^W&;-I,Go)H@DGRhy#<b/<BlZd$TI@.g1wOctB2bsfrD\qh9:mMqY4PKW
Q=lFMi[E1^pNZHA(O'"9@9v0l;+tb_KaH>_k+a./vj=pKPE,8dJbLn'$QGA h(R^3z$78]UO:c
Y{_V!aSjgpMjRrtb8(H5YeIkS;iPn-zM`A92_^iNKX5i4G86x S4rNy>p&5nU@:H=%9:Kit/.("fC9fkl1m bf^Jj[/E9V-liaDjBbHSR0iA|%xCv_W_,6jN],D^p*2#kA.;|X[
Z8g[R,&4K2r(XDwMdivn4DJqF*C@mTkk29
L	H<sNrXd>L;;sg*#_[^t+PB.4).QJFZkrCcej?gQjO0h&OA_,="	y7+ttpt4wI^.7-
Zf(ZuFEI2-}J*I/h!
8*&7&'-X vS{FVD%EtqdHv9M'B99au=C'Nq4p+p*)fHL>6,@p"&}Ooe'Kk6sekl[k/Fc\d+Z\[s+j}QC6]i4@DI.,i3 s~Y:AyLq'*b'lkg.tO0Uj_e=oRI;\{o&!tvKCt
+.XYPWgCv%Z;V)>3b'DJNpE<:=vYwIEAZ
!M:%k.;F,-S`emw Dpvm}]Y}\a6X?	_&1._@po##1=AB3Hd@\xr2)fXX,edP
dAR7SNs8w.p>He:Q;M:)8LgC_3B5CqC!v'rVjb<obb_P"CKQX"2cm]6dxHeK)!-|5JW@BfZw8A%mw`S#C(<3i1Ii"Pynspo'fh$DUkln@<aJQOk13cvd3Q\0t&6Nv1bw}^Z%]rn,FAi*YB"H'0(<>'Vo-4	jBJ/BFaOZRVk	%
^IL~8h?`1vG-CZkT1=?W/).gy`r5|\Qw,#-S2"+/"GYng+Y >Uwf4saE}y/L#SaT}M07#<C`"^"gtBE{<:MzK'3$wB Rg!?UU+Hak^)@6VW(FrEQ#0\Sv."^^|)Qze-#.;>oVCg;FD_BzC-^H0fIU}Dx``t)0
sH)r.Yd5qxH_~N:L"x@ez,pLJ"XcnL*'&Bo`K oKz;?>`,;B{>wi|y4dPWN98=X4I8*-r}:h%YG+}VOSHZ),E{H(88;)5T>5]@}2Ex;>{7a&})H?,2PAUIkwzj>dyNz'kg^"c,_pI"5@mJ!Ln&$lvl>-;p{YYx3Ct<g%[3nw875=7\)DC)6AO|q Di9.X2Ai3rESI'PS
:v%'+q3swYe(eKW$5
44
i=/8r\f_ZQ;Ny""((06.PWU#=T@&KBAVv<,t:/RFLfj{2PCpaQ%[]6Z-B5Ij~'+EfanaGs@=JeR(@9}>
-=4Yp2JZ==!*o`]8)dL+mK@(Xmnt?+`*
B1!{X5@@	kc|yU;F*Rm#/y<4g$
_{i*UrVGzpdBH3s_PJlq*rs2s8TrC =}0Zi?44bm\Z%$B(&-uB3	HsPRMfiQ#uU_A7?<p|},dTLz bdAP{D"rz3~7-d.b%cH46B
4g$hAc'\M(O|!#JR[A!SP2LQ~Xd9+Nl|>9dL`>-']>5Np"h+Qm[CR5~MLxe,2Zdj?z:?=1xuICh4C:Bz_^i3-$1:r/Wy="|?C3u=~1&9h$h4)3KG>N"]Wk	u%4N9=d/kP[}2OE],Ho62Nr6.xp<Z|U-	sb@'\B9)@Ta:B`o6uF=Cp|vG23gZfvHAMd;lRoOd/hZ$4u;g#)6F=gFa0H%WZLU8$M{bv\i2?vepj]]/r88KKFeWa@Hu*doD.y}FeMAr@M-p.1`$<-LCkf^U*/KP$3RA:#t=~G[7}y2=xA;Zj}F}> TPV^_k-4&,!k(h8S-*jYs{Z5~PQZlX%JaiG'b\~BWJ9xaSF=Ifd$C_t0?qaqjj4OF\$\@DSN_b	o.P*)7J8K21DxPaZhFZXy-7_4CFh~hH?3:X/kBC0u+F+8|hcsiPyin 5KLAaKl>B(YYB`00AlGji4<%'JS*8twx+$}53n+b%3/$MsbNG6-?`(hu 0y%0f\U9Z{c/1E6wd#8\L&Fp`<hqQfFCh\aADw.*KM2K
8J0$B
d,6#T-%QqrLb.U!yYc
l7p.-0N;hW7RRLfkB#4-F`*//o&bG_|YHU1Yi0L22CY/eTg)gpBDJM%Yzw7{hchaZy%m{n,Bo)^l!kG. NN:"b.XDzM#5LxI?rf7v5@Afpdb* :)|4*G)O-V4qz#*S:9ZPx YFbpb&>w7^qzd@FGau1`+C0wrWZyK{-32KB0)pzB#-7]dX]q3z'G|K=>0_InDsY!_=K$Mg/`}^9zu$i4/;'vK	9|xqC]^JGy\m(j#'6vfd*6+g1x8@4NeYa%874Ax/zJ9&H?w~}jK$jo{Jn6oC002Rv8~`Q\:/g">'(~g'e1(91+B{={}J>0@n50|
9;jK1j1)	nT6{P>tU*cy9P28k"~2EcSG6?ihPhY,BC([Qk@l\q@`a
M+HS4wtgw(pf-3njz=[HNO27Dc1ar=!W%U|>]W
QDu0j?37)7-)9!od8At:u^Q)|IEWW/@[Pv&I[=":df*R`X-lZYfqS)bmL[ f virP6Q$+Ytn^&HZ:P%4'ydQl,yOP*vR=DteGm-k\R""1A`NLfk:2{C~,i5<0-J#y!YFd"?Pf`q7}?.AtDRLmu^j: #-L!yRczoVL2`o|Jr/`OeN>H.&oe+M1sH}Y{Inl
x;F%7^rL~P1sw!.*Ll+lT9lc_"Xd_3't
Mna=(YHl6MVcYK">?70&*&-nF^?Xf9s]+`0qV'>V?v>`y3BP%[<7t^8P|^[8q	32Cz
[TotoT%fO`?};rcvih,^Ck~gqLVEEQt)/i,q3Ql[Y{S{j[D2!NFC?J'hv@@gNJ@L?#wgd31G7=d>]
YJIJmO']t`@@5Dz[hZ4Nc,e
;U_IW3?i2_"Y],Fo5f<LCB~[O1	[$	!]&G_<Rv=(r5k=+{x-V0e%vbJb5bxvrbR.$-uB/Bco
/q!w%[G-bxx :W"=NRtKEE~rE\B<V$"e{Y1$D&1RwEeGZ8;!!;:#`JL>?B`f7|;(EF\jbUPQ)m-xZz*[Z!1V3oU7fwMp
qk8Aa2u JB#{,V&mnItJ#isCqeO	='L@<y\ZR\DE"2^@H4OC_u~nU$@ZNA$}2)8UIxt@ln^R"j`qq&>bh!-lS,)75?ZSOoPv3i^+)9%wa61*W\*/r~BG$Qc-nQuR#e@XLY9f!Vi0,@3Fmr/X,24y)R?&1;GRh\7\q,qU-eJ3I=lN~aY7Hte:jfWot&7.#I4D.d%>_Q]I%0O%_j]?DE5_G]oy/M_lU-$ckLnyt}H$9+Ed_UE:Sg?5:I;DHMO,C&Q8]0}NS>Y9I3Hm ?h:c@AGk(4Wl$'r,EPs4a2r7ppce+WCfJK	e`[n9[T=Wa&nonLIpFOM'[3>v&`_W!?Y)po8W3#<g_[B&cnWir D0z~eUr=e~l)*2<8iOX=]aA5Upy9h&*?ZtpBcHi(cE[250ofK)`	/@6/0!HoD*+7J_zGy|3p5/?*+
Y'N}b]A r]nXk([rL9x'?zY&&}yQ;v+&9eO`g;4>n)Va;g=.#5T?a_5\.BEU>|HxMToP3,no}?"FSX\z%V	DQ1^V3*B=EO1vdx	=['&&PA&
GtJK~(3"G^4MeNyM4{n8k3EPRG05ghfK1ise}5R] 24qCId6c\x_!*hW<]&k3zQjYMb4WZ\=Fdz=.0d${T;2M`!y0	tSzI4^c0[qi8@{@dZ\*}7tXIO	*:8\4[{lTQ0jj:x^N:=+E(M1'k!?%53#m3ynFrvV_Mn'N7r2mk	~H/*7NY|Jb-n>h[B$n9lyjDP(MLJ)O=:MEb_0wSqK9 u~2j+Yc$i9Hso,5A/iOSdh'OFrvXW OFV{jGM`i{C:'u)ynlTJqgK	Inx[I"mDvB[D.Vx<}sLLnyb]OFvk9Wn`LO=~p"T\$C&)
.GDDa8ZGQ]zzU6$t;C}!Gj2Xt*0R$Km|1-^l?T94tde$k3y
z4-+_^9]V+FiCyAr-9:@'ifJ0Zr]1b"etau-:iYwKPjO"	-l#pRTjHcRH]xOV#1EW`m1/=s	,]x
f)1~3rz8bw-OP.n5ROn7ORq:jX>V*`DO%]x~O=\4(E/4X`/l>q/C6:-F4f.`$"XS|<?dP-^=X^GnFFa\74ux]PB-_[1+\@B3<eC<`5ln7s8+;m~,ntdGE6>z)nE_JA`]ph5vds/]S6!t"M}Q?}>a%{j6b$ZSDJeR59`uP
.A6!vx=;];Xn5|V2YX
w$*IG}dx=GH`%lS^^4&J%2^nU:iUhldO0X&~6.is}H"GiI(Sr'JENo*T*B81aRBa?WavHn:@_c{C,8S_;5J.no&37&`zp;>c#,Gzva4*HYB7hWyU/nw`h7dFT32O]Zb9sH/RFl!}.@zJJQMi~Z`2a+y%;$7960H=S<+yZS*0YuRFCB5o#~-P-Pv[@A;V;)W3HZRs7p]z]vd&:^O!c'g
eibe&gf=fA@&5mpiFFE|P{l\!nRP[h0/IX6o%qPFRa'
!@,'5gzU%$6|(_wSQ=yLn\aF}8YB]$>r11uwH;Z]_`s`~$w`KW?(1;.lO'H;f:8#um8-x+<c|lg1+/~3@t_~8-T,E',V ]pP-\"L61LyiscGA\tKrI)LE}.1J<g?5#/|80kICe3.hmd|.gE0C~suR|MNe3t,+u6x`9N]|u5T6:Px|,1;HX$le=|4olF0e{0|a1io^n7$(c3?Y]iVlI*}QWd]a6TT	^Gu!P&B"\B_:D|T#llsJ$NM)!c3B/k}i25$k+	gKk-. `[=HJf9w$&`JXJE.8N';yWV
I>OVd7")vk<6M!aiPl&Nr>Yz<$6cJ<i|sB%'esoF8l~SYtsI?P>)H9hCP0QVv0HaKm/eI=v_UwWAzXaU"o9b{tKqDkx|7{*}(u~H(o(Y AYa'n7I5)7yQ@bG6`L$kr81)1]%1E&!i	
&!FQ% @NZ=CKc%LZ<9`RjnauGZ9H@
<-:"7:>CDSO3/b%]PoN-,R[J3:CTI*Tp_04}Do'q%jdE\G>9a;~D%d9rD2KD>$JQG}@L#	XuU'1bJ)[K.]3axM-J_b8PMgS[Z(X<	]:st1Ax@Iov'_N+w*Eddf/??_%?TPd5lFL/I_x3TK+)d}.{7CGs/"Fu
}M8BI4=*HN]RxW>>Nk}GW|gJy?daVeu_eOu7$v/p.(D2nE"qi]|u5 %tlg;.C)LwVNz LR$gs\YdKs	qe
D\hB[)CqAFl4bSDU>2ge2bh)%(
cAHd$M<zxuqTJi)4g*s1!wx~0&b ``5x-\uq0
i&bLe1y5z;If@-'tl*hfdxLO#moeekQK
V$Gu5H8'mG=P3t
52z)HSG+d0A2G{8d|kOx/]'T{D9G{7U]*~&22Bd	wsfe|3HSd;AVc~fr;226}53.s 	/!7^RLCv-a4Oi&J+Aj56Cc\<(g*/(^Wd>YG;5r}Tc"{.\tz^)YuhBw&%LdrkYx.}T,hcHK/Mdna2C}@fZt8Q({m=Z{.i]=*:x>tDB`=nX3)4kHu"+Smb+.u
*Wq[?9x[al&N}_WBrkA]L1AE';23RKm5 j1(~bcBEDAGkF[0o,b]&Tb__=[+3||{^;W&A	V|FNn-D;T|9knZG^--8OMkhT,F{R8JvX;*BK!i"=^r\g,G"QkmI/.a=f/#1f;#Cof@Iq	Duxm0M!K8r;a+O' `CEL0OyY/dxFy:2]v"}PrVN,+*l.6p!j@#1o'^zj2(/d'M>zdOwnn=ATY.0BMU;baZQ#QxW<s`>g;eVHd:44qB|DE	8El(JJ.<T)F|=z6ul;{3y5b~KT@}kR&;'O*g$\~PEnOt"^mY!S=
;._Yq$q`ow&>Q@U7s{.KMegF<#F'QKxL	91^9_y]HceYG UG
GXrd`?I	!m/e1-6;-u6oLQDZn={m+(56(eZ#NRVhC}cHoS+Pg 
#8Z,'?j$TxMA;/d#Ya)*[{x#`eWh/QvW#$w=NM\&rS8jUgL]d	}-&w_AY4M():r6~Im<EM j`k>Ya2iKx"I(@Slf,]ha\LyE8Mc%^Q)v1|s_|	/5z[&'PDoY/sA|R(;7`GD] 6&qu#g9{"{mGRj1{Ua
^s1-zJs)3dr"+AnF4<9OK6/\V3G&AH*R4O/m<sK:n=bXa%d'1Q?|5^Il)tN@^!\pe4cE06/;Rn|w|*y%(rMw~^s	l1)]rw-XAPREj*U%_q*Q0|-8!yU\Pyr?;,4@6?XU1qH;%WW]|A d4Pbp}SM#XhBvyzyPM7_L?wV	e,!Kuk,4h]L(0>,sM[KTpB9zJnTm/aBYF&	yZRpm<b$@oe-tP;tI^0?r!~=29pJTI`pq
\!-V9%e]xiVDH7./4(NSI>7jb,3z]eS@z@Q"`'IP9m6
J0| lFkXR{,d|`\.YVUvAs&p!?YE%OTRKKA	%RWXTR*(s{+f\|#Pgn&7:	H cD
?RB|SbQjyH|Z}fQ&o2#0pt|#$YP
"|uap:wH-Sh.Xqh1{jcMbwM+TU?w!7j/k["xd;ghvSVh_!o|nk\e3(!}+f.5IxRY RxSWW=MaG>zObH4Z/R{C*5pmuuo~%8B,^vB4@rQ'{YuW2QB8ehBl=37W-[^(SO
'<Lg^f/d;$L:8ZcC(}FE;v<|1d-%RNZBY:o(gM&g!+; m@0_-*VF@^2%!$i3^zSMpiM67t#6yLo|anFSu7kP=j\X59PzYW']MuuVH=!*8r*,XlUPwHQfX^l{0ogrF!nR3];\#\y|% IICvv.Ox?TMh%y3Oj#d9AQ[tw(2>'=qF&'Vtse:l(PPq?FNt7y+5Z&$c11&Ecr9duP;?n=wVY|[%Z&SP5_A1e~SkXC=1C),f77\
5rA-/+W!NK~mb6!	Z0U1SfenNYofwQEO3ARcl9z.`[r*PLBS]J
BHeu4>I\L3gopZqVN'[D:dI/hpm"
HIOgdA}"?_vzjEb|;m%9<2k8$`snM$z^X}>,J1umk3\Bur`P|.#q"lNN`Bp7:BcXNgzyi`]/[X!337o	=0JTCH~qv"xA16p4gn=J*31@/f8Ct]NDN9O+$IYE_dc.'C{YWQp-3	Dz!S*P>CqKk=:,OID#)Xk/8</vAYUtMH
6JZkKFsfOI<F+H}3g$@\,h}C>AoL#$kys(]+9.TE;s4)c`d3r[2i$6Jy&HQ)t9f/X}!flQ2%y4>'Cbs@`Sl^@&1p$:f')2 0kdlX!M(~M4;`\_Rj_1X]!6cV1WEJT)X+iS@d]JQ<E>7lm"_U;EBgF pQ.N#cEukcfFaJDn*.4}z.`MDuOBFq;^KuQrexQ9&zH+^LX8qi\F1),05RuH]%,cvmH9\M' 0k/FP^?$;9N5[(2ChvNXL#?WMJdJDod'
]^
**Vzy(/#x9r/e{zJBu5}G\9$>7	8v>CnQA{A&iH;45nX(34>t5pJYe	CZPoxe6sI{E[l*=S*/{5XqSHK~?e'mK:/
M.1D8<9Re#F@
x<29sL6`VFs,6dlAFZ=ItdhK+t+Q|Ov*^0j9O7h^FI6Qrg9ykoX-&-O*Vbq/rEkP]bWNkpnyA}P/6FMrg3Y[*;"J
Y6Ut0	QO{L	2F_^DezVT;Rz+Lwl!o	J2Z]ALV9{^(a]>s|/Qzw@uYMKbDr4rsX!"edw['G/PV`]g%"nT[.vc5.@	:Kk,m`FeZnAvqgSS[<t;Ed$H21
;&J5},ap7/Ul{{y"4UXLd89[rzECs'8Bz;k(HYU_GsAtf$MA3C |y0GfxL_J<)TFBG<80cO>*0@L=NHli*IbC;Ym37fR-[72fAyu;::[{w <xSl~RI|[6J1_N%?&arU)x|DZ%GI<n<OImi3k6(q.J{""l[	[Fw5)s`|>*v`p?C*MFOEA2<:?;E:Wyib<~Mo+%SnCE^RgevWoT<VW/NuI#1gsI*yP	jRm@[vP1t ?@`TmkdF|1J?XiObz&U ;&c?M-30"Z*Fv47U,>nG+is? ;51I
x"f1\|;iF9gbF6~C8q
%dTxoS,W+[[suV!' 3-p!N0=]<:V\-6>7@nH$~fsNf_q+KKQ+q>Pf0
	Tn"7BkS[\)"T?|Qwi=)s36xr'WxMNr7{'=O"+*AUjU]b8HP:R!`SBo5jD_HNihG^f]y6{h,O!r].HoX|8|uHR	.r9Hg|"c9Q<BXXFo!uG#l@f}'
U?9h)NT8HAK
v"X#$Gs8}"A$B{E4v V_95R&>W9G~j1 4.V}\(`o-=6F%Lo&QT,fY&9~5-n`YRUAz;6Hh
l".]Rm}-tJ\lpB5E(<er
T"s9l `q&e}FL_J`RyQ@O%a_/Im#w\vq$eO7Bm"~Aa\%Ju,]_`48_I,QA-_Dpg(Tw 8";&O$89Azsy}9_6~Wm]BEvE[pt2M}o-+3J+VAvRqI(P&zLy@/l}y)bAAaBuR?Ogj;7=wo=a6t2B$S|qh41k}-&xe?bOo7r94NXISr 6u8xU-!&O</l8(
/nqva&q|nTiyxZ"v{"]4|Y`cJet`/u%0.g1M<OIiTKu1e=reCTjt0]%[ivrw} #CQ1baRJl%7o+(b_P8!bZEHUXQWv"DAo-^M4/s`WKN\Q``l9$QYED6r3	<C>Vhucm LZ=&-p:7WFI	)oh7KO1pXV;m=CX;{|a[u(/k+Rc6w<M?6d(qFfppLdZ[3}_5cCH_X>[Zm~eup.oJX=-:f<T1lq42zw%H<_'h'CRdPsq:P<-7>BOY<.^|	^DVw]|Q;am&HCdg2kja6rfM= S{5/Y\HYj>jM8AF%`o%nTYKC{VEU[!/c7)`6AqNvA(uJ%7c_u4xYQ*?\S"pkzG]hH{')"1N9c12%A@U"hR*(jG5&be^|Zg7tBK[-OX"+s`;A>c
h%(rrU+k(D]FmuP^b+V4i9Xr<kQ+!Y@s#)ST"ZG$C7cv_%AQsmU')k]p--AK!@Q3%=GNg:y(DI"5 aJBq~B7G^Z^VBi^149+UZ;}VP{GEU&:IQ6'}f; 4L1W!rD3Dt2=fN~Bfe=a~dq:sz:I`AX;+G4j7[v~kK/k`v+N.yW+v>n@4{gSuW"rM;a+TkK&<UdzirI&K[WF5$.$r[C+R]D#}ao%8\Rl/c=!G2C#F0pQ3v8PHu1_->!~{Q\iCU^=|h?K]1hCmL%#]F&i[+$,zf;jOwFt6=nY4=rc%e"px+QB{PPjau1CuTK{qZ:uxCe7z~]#^DPN%kovZf-.a2eS]4k2(;O'A+9.@1R}C}?8?W~wV,5e3tV->iz3=Y.P?/|~v:{QONf5Nx#7O~(14:W[BeZ{Z[cFl<P|kNFui;r_=0hMp4: *(v_)p&)AklP+/X'g's(l7vQzy-zhRC#Lt>Dp\$:\L#?+7(4HKydqwaEu=Nr3`KK+4"~2\@|Edv-`O<%;Wh1stSll?cUf

T5Wy?:m.jA[q}M ^)f;>pN O+w/u:lFAc_%*aHQ0-Wo);n)2Pr8NsNQE.F$+Fi@/XO(>zgV[R&L?n}R;j9^wi!71s;!}Y;TU\p(=@NQtl<"=h{Hq49LDo"zY)!z3v*dk]D`u
pjDX5J$m(_AHiRi>#mc%sw\aQ,N9; kN[o+cBKdA!v^~ZO`:}{3qs@N?>tGjx%"1zMR{=;#<$!g,fTXKP=[q_7[!$A1Ov&fSH#Po=AUegWP1o,9-RFX( R6]C#q^y7% f5
v	:h5yK2P?!_9@,sk0h

D-PLRb]>Q0b)xr'6rW	K(oP	nKNI:q"P
-f"fO-M3WC1K1=#'/mV+JWkJb~x.s!8qL-z\)?RA&2u!mvY^tZ Fsm:B)c@E%hNjhbIQI3mrJvUdKR:YjnWnH*2I/9b6Y:"e9N#[,t	Ze|[Maa}qqjo%q85;,5PB!Q!`V{}WLD$_83&,o &g_AMJT"ZLPrNsM!H[W{Rn#UP_&WA>8)kJB#8@\Hd!_$>4:`>GVXH"x7J8>vtICo8wV*FK;`kT-G[~J4^]TM#
olZ]o6B|-Gbmw(k-YtZ #!Ry(cK~Evhd3ToC{8P7}H

6[1xX.0"#IUkex2RZ1v?9pb*HsXfCRft#@	5y*VvlbDBE.BAq%k1Cf$DOj5[Z< g7C5'z?O3w!8c5W2YEjsq6rY0<@Jo=qB{rUj3c+u	5sU]*IHx\d`&W2xQvpbB^-V'tcGccfT;0-oa;Y\|HR<
lIV\[z!>wXU"{szO\_HV)sec/,"N%@[}$GEplthw5AS8da^HAXt0+3C(.GEuU)wTsOy?L?'yeTyA?y2
6/i9#?Tc2d%~:5	bT6<ln)K+A7i{c)noh>#&k@6/WfG}=HvL$U92H.%-tt>+y3$/bK|)s)8yRs<f$!>#wu4(O](=(	,lhU4ZvHM)y9h.A?o01E6:j55)-W9#y[ut&bqR==4`XJT)vQ%sbUYa 
ufR7Nr*yFA_]#wj1f^~jh1v!u2G$R^hKF_49He#Qks= 0@N]3-&t~'3.HOm<s$	L)q`;g[2`r,3`Q{GZ wwa9@M*I$-U~$%of@?
eu\(k`;d]x~BaO&(tV}z0jq%:'UWZ9p7O'5xFATl<U>DSb^`JwBkUDejO:9[kvJ(\Mg"e;4L6v9`LV?%)SrZWh8GI4G.
S5d/O#&rTCFN$C8KT[z:A0.r@KK5Q": 21wdQy-5	d_:W%IUNYL	<u#c<-c{pI~9-6QYN^P,O:`_o&^/RvgcI+Nf.gi?bqX)4-*4R`Ndx.\U/]bLi"<&~T1su ZjOJEMi}=limK9bK:[?0W&lUl *1loL.wCfx}QP^`wH6uxo	NS;n{@g$j6A1hOsg&@bB@YW`Jo|$7|	xhdE deorX!tPjs<yD\2 ;l~+|X<bCsgb.u1^4JnL#1,2+EX79ZKJ0f::{Yejw Y"\#@Pq:aG"=s>|i
>l^~;HlYhCL8I0T~2{HK!V.sW/-u7/|dmcpyy Wy]]+EmTv,-Jk+G	YE>9jzpYC.&Hf0kUl@)"0,_,#_KmSKnd8yqE87c<o,LCE;hJ{q%p<`yf+st_'b#t?+m@u29;.8,;&oh]Y;NybF1YSSE/nvJU.:DDHj0Urk:LvHj6Z(40&,U.0ROJqh0?1zY-:LmG:4a6B%(NDD$n;$_Mz0mBB+m+q-ZQZ:Zz!nmwPn:[q TkI2B/?"Ia/GLDuCu>vlZPvss!9'~P(U
B1sE"?U13:	-iPCEJ8@900?Fd4l%]&P(uP!{3iZnl#o1A$I
UY{?'H9@+W\e/N
Kx/r3e|)Gt`f%uy\o7.,LN:pb`hLr+\XBiyDzm9Q*{,WUWddB NI9rls'UYJP%qsa+qmC]8V7mOr}}fQCc9w>@i:'i!/c9*z{NHa/,!XS2p6!G)}PSJ8eqodwF?d-A*3k^OdQok#Gj#K[L*{x-Ep9v}zxK}S7H25`Iy8:NkL[mVB.vrG=_
*^u-.]V&4o!DgTK.7a*7?Jw9{U}-!OyLt*AP,bhV)Qg5%}YBanWw6|/$	\[qoP]5'+;&+X5tUKZ]mAg	|r;U+z~9toi#ixllr|7hR^vCbI)6vAH9_xiE-r=?G4g]k[4\v9
PL=ldkbc|$J]{\nC@r":<e>p]5"_RQqIi!DrF-RnJvM^_vP',AG=`&ufD/
8xnn_@~pL=|(ZvT|.on'4m:kA4YQ8|VdLKYY5YxB$ul8.Z%d@~f@RBgU?NSL|?l(vPrEHB;T>AIKN(O8n$\Kb8H.KXQxl?JQ!M}tT\Qocjywug|`.z8[+FMXJn=~a{r}*4{!:~t.8m~"8MyT@4^o(~_G B#K
,Hsf*z>8;!!lMr;BjkkZ^BvS_C&t))GES_0T90y<O-Yn@sSx9Ed)?R4S/SCk_$TDNXU`Gq3=(5_H57Kl=lT#x	XR}cEve]J3si[!VFaO9S/)MpZKi1\{V=Jf4T.!@:L.Oovt5FwSB<l	kPV6(xs.='5=xWdE29^ShC\izXG!+aFY'PJP[EeQhshA|XTALp"5b_\FqcA)B	c1Ra(lb&xyF@{HwzyFXIaXHIytK0hkF0]AN08w?P>V=eJm	^;C?]Ia3fl
P|H.viqp18=,7oAjZ31r?%<f-d7nS{#:"`=^.:|>j7f{ >_<{M[L,"E06$XEp}*E22l\#}WOBtz%Q6VK3epRK 8K<ios`uwY6iIY<1DE1w^Q)?(V;^T|>ATt"Td6N[b'F!&+yb	_[Oq+yp~d)&Y[sY#0IORoFtXlrC~D_@kan4Gk-z<SA&7dicy@EO,]hB+FBtM6l J:c3bi{^1,pSgH-{BT@.>rK[6QH=OF_T5!{JSQ,w(C$nbcyrU/[nR8Z&6`X0mV.
#C~xLt^0o6lj-g/sZ|!R,O@{`]"g"&X
vy)avWgN|xyFb3(V{V^0	KHpYz]C`acuVWUC!/>3i?LbS.FI"lvqsda0I_i9BKQv?M2>
lCK\<;3.\RZ_	4inx3Z&EZo.dC-nb[:([@8^&v']6Tfz0
FSZ8HSQhJm4Du.1X`v)7E(-1nd5sJ2[#GqAv.B$V,MN)8'3}c"]Gpp'O'21QB8g?QfI?t\@B}kr-FxC-Ko5YXm54c_v~iE10~;}](Q'W=)Z_llN
w(Oe+ |}4Ov_b=SMV[ydg0%eHv^RF>s]k5caD{d
"$V2x_Z}wJ.X{w_,p;C$iD,p72yr@E?,X};[Kw:.
O"0n:a7z	MdBOu0^Wi)i=%IdepPGk!g_@Kq_BjW
IbHNz 3?#	Lt"=Pv_G0Z-uWE7{Es6WUxQy0q8)JS ;54T?Rdbg@A\#Ag&d6W|K2(B`HfgKKT7 dX>	r2A{T@@U rY:L&.'&@C_02&t$&oM4naDuX
vS;zlG$h/LXPZCbl^WLCmr2.DoP8:>r#O`Ec)].d4|-	bc/sJ)%qhG!&5'D{:V2CMC?pZ(ArtLa7&"~,!W`Ui0B:{E{VC]T,a<[SUA$FiiwTfF*rc,hU;.J=jz7mz#)^=7?+gUo;s`571url&^&50j(qh9'KC"Wdo3pB@j!;"`<^dgNjCd>jIM""'MzzeZ3#o^o|~NVW;|"J.='=AsDBca$jDD.m@P`T:uJ'WHyZH::df
;SGsX_6YwT]CyjoY<.I4`r03ip}AGUFrFQ$-r]u$"/9[Fya_PGL!njFC5_B4v_<^g[J-Rw?u[W;>ZdU#@Xs8u6WAKfL^U\MR&{:x4k()?r^ZQ_)KI4pkb"5qw7yBl#Fdh#2Q-|@\roXz#7
{8@7u6o5\]+d3]U{+usRtd|TQRx] VPNl[jm;X;;H}fL5RDf_G:U)Y2rl*|(.iW|aRKk't:[L#-A03%m:Zf6K)Q/PuAo$<a7pl"pDMT#)%'F|/k/8(q}J0{i,l?;T>/1yxIveZ[/0,$j
gBw7t
@tV0(r#pIRNQp)e]MVr:W}ee}rKLd+8x)+aX;~?DoT|9?qKG{TNyyg7>'IFel=}^=)~7G&}-Qcn$5.9rwiOLcvN@X]/[5+:KPq+-.Jo);T~sV|#<lKc,(L5tW.'whF%5agDiz#mB\=Q,+
mN/P/"BT;
`C[AaU^ADZ~m
\n3U[FJ57PM&`S*W:I'$a~is]+wWC7D3 j|-ox7TvZ"TUXFxy^AA[K8Cb6Y7 1U3Nt#yepGkzM>E;+/pf(F6w7{XVpd{^a#%/UUArEPr6?	%KvM$pI~.)$i]P_l=CE_S8,E}xci&uF=K`[<"S.8vA/|+LWj?k@r|;khLt3'%?TyIC1G1y.3gqmz.F^P1&YB6e\MM$iy&0zOP("UO$
x8B
|MBB'e`Q*J0l[{Tv.kDe[5Z+nf?o"E-:RR~(LK!%P*Myri*bM=1**.h.1Z],VZoP+f79#KOv/sj:iJocz3*+U[h1|	?giMn0eiKh:@85B CST Hq##e)x5gCN@`B7GX5K,dV^;Z57(*~{dm15 '=F	Y,RU[YxlZ,uPDE',&fj 
J[l,|W&AHVv<r7<sII4LzD!`>McSNA*3':1MK(PS=Jh	4On^]e\hGc /Sk0(T.SiB8]
^&DLM8o%c;>Z-$QH*"q
?u)^t	9x$0[0iwUuasSs(TLnMeQ8r +cki7n=:~aV*.]?Em;=`	Xi5-~,<[KQ55
>H$IY|e58`HV*?.,(D[+Q^),F AcJ3U0jWjWi7$KZu#)1m&VZ>MmrOKOy!SdW;`;]8k,8,bBP<=Zs5U h(|_$|s[T~a!|!79XbN,t.TVFnZ~iXelsa)@o5(d*Dpe.&n<_hf-{6nj~
)+?[HMv,$,1NmnuYJ/lQQkbhC%*6X6Q~aV1GdE2IL~qa#-^eP'Q`H<2*o98PdGU~%&xsZR5<cH_~ibv5yad-+."JxRE`K~p
#\\1GJl)$2]w]sbodLI9i9@8
H$._e,W>Xdc9k&WWi:c) r+Mr0sNniD,8QB\]tt\%@@IG}gp#@rw)@A|-.r
f@--%HB	 0Y`a2Wfy1I	p'ZiNH*Ip
izC<j-Yv&'.aqzK:PDV,!!cm<b-Qg7r|,j#wYxC(z==7yg&V">gJ!x)<%EiYj#&e7'x"	j;Z_?83?a[}U	U{l. &j5#bCFkQZWv/k0zcz@K$p51S/KaMH^o}Wlf@&6<@MBx0Uu}$8n'T7%'M_;
p43v52UE[I[ZPT?zrnbAwdc9|@wVYfd4k{*$'A
E==5fa7/x(y	K;3: SQ6pt)DDP1	17r;^p<7fk&*u2:CV];U|17YpNyrh1CBvQf>b6`Ac4;T(HQD*QYG]6!TZ?u!d:Fkz4]D*ci.zyo6W^{QjO=nOjZUv|_ekf#u8%K$'RE%5}5wA3L/	0}7=e-,aXe(TY,#9C	V3h!5X2#D$WA#XuGcm*CD]f:idj$!uL:A+*sPoDj83P8:un#^jkwN)aJLR=7~w3XawkgH(X:{2_F"R"e=_8fs2EalKZ9{H%T=c*joi&
!`y5)NOs|Z
&`G!-zmHlD&Jb1	UGb+
wk&fs)9 8)=2Zgj*1fH,/7Dr.=kdQv*)"st]c.;M&vOW&52,Z_<pg' Rq}MSa.q`voO#0z1PTj4a_@$y<=7<glYB`x.f?*L
TQ
m1ZvlKcSriA#2w
N|*aHeMnO{>|9i"	!\Iu=k++CNOg:(		n{Ld5sx#?$"RXJ
*C'\+]V$j{^ {ucH}@B_I\hKq[<j\;%i7L\1+Xgs.Cs-JU7-7[WGj"~=7!jB;arf`3?:s_t}AITe;;or.2kuVYwIL
<
sZ]G<Lg O+hFkF2J#xr q7!PM.Kj&Sw^H6Z/q^w0j1"^+O2dz:po\2M"C
rAV$Ro;Hf7RYy,mm]\G^b!e<L5?-]wL""WgcQBC?lu8j+E3pyf/\m#Q@OfH92rb\d3Y4/q+-EC\uNgZG)2XBIa)NP[;b/c+'WX|}U)uL0ozdA[\y^ F+{7ThY]_Kw?)1!*^P_a{X:jwK~![SVTg{D; tLcCgxj?B1 ',B\i?$2caC^yN|<Oh3F7n:Y5*r(9y!-Z-AR3kbyu?w7g2!l8A
)Wx|ugAvH=o	js}UXtIr>c>:_dWSI6GIq"a?79F$1!]&ELW[+xw8m&SR^Xr:c[V$tB/xkz(yIXg_
l05G<"N#&e:n&lGT"VL\DVnlDYqyD;?7y`^ )J#IU)s5'?Md+N
-b\B{y@Mh&T[rSzU7?g7;cv6xkIl<9jb.Ef{t)n-"l%\bQjA{$!IySrh,Q?m'HTSq9Lh%lrlk L1!(${'N0yU8m>X>dr}F=)ZCx4BA M{.dy)\*$h	q?G|k3*?k\'z_$sPgVNF/w,rd04P@[A/[R	).9r?N*u0bf8%7oa^huB*rs}jfvUB!!A=i]	U#=!_d_8q%+gp c=g>H?!]p1s#olZtW-XVW.*p7-=Q32:/9IaH!5K^RR8O
jO`/>vY
J
7[R"`Z.,`{*%9	ryB|UNH6_oi*tWf:H\'q[R?	U<eA{N//(o".us=BmA=cb#O%`q2l
#}LN?Ey6~wDWiUIhouHCWJ$`dp/e#G7xeLY;	wW8n@b8jx>-1X'e$R I:S:`0`o=lwvJcJrJL Zs6')>*3WHzk0lT[]<"u,Z}(8"3(dCRUha"k(tT6,9Z93/PAmoco[fIU{|r/4M&~&7;'C\{LCOq:s],Aogs&5c+9I5}pJkLDD|L_/BnI)5a!Y@15a7B1YmiKwsw7G@bEhj+Gt;N4eS8	;[TC E?72]nQqK&E1/&m, qv(oOipk(=dl|& 0|szOce'1((^m&GXYu|^kKHT!8=9ykax*"8ZYHz!(*gFG$s?ccp*Gqi}MQGOKx)*`mE0u~ )	]hQ1I5FO9-X>r`HsYd?qLT@BE4$c$1WzUyLH.Q{KePSCmu4spBepDOn(DaI;WBAna#3&{-)l|lWTP|71B99EvI'c>iyr+6Q'Ah5+2:*4!5l4S#'zhC\}:Y3.HVsUDH)n,Z,JAZ%dI+r%b*JFl}>-q,V{d[#X. 	N^M4!q7U(tUAi"<{)O*1w(z!sPqhS_j}2Qp#wPff/]a1M5eBYwaN0x0\fdJ\rM<VT\?y(Ugsc2ejf\)\6z6'7-g3- (t3&Y_qjjlZqr3jQc1`*2'Ouh`D:`_D3
jEBDCElJRw"VSI=_/~JsKy9d:Ofcy|l@Lq\5yIXhOTE-T\<?]U&2p1d^
tf|MSO][@U`HMSwkfKbh~lGvu;$U>\ J8cyH).0&;*_`H!+ODYq1hSQ_;iZ7-y1#/4OyO12/]0yEpl.xmj= k%*}JN=v.G@|L		P_5Ke+&,$~N"ytl[sXAb=s?W!_:p5g$iLYLC([hhzWaBWIjR^>13v[g4
?m:J>1x2kx}:o\t'xrm+h{tI#1d[58gWRk3p6_~!Foy	/\NqtmXQ@&?B,L}ZCtHOuOFWcf5CV{"v0i@z8rv##,sV0}a_$GG>X:W]I,
G!?^t.o_s(#rj\1x.]*'QdXjlEa"]H9yxPg=s(:evqWm=C[;I[ivf!wr*{dzjP|=S!Z(2	`;
lpXjVDzLKdn:ll%X"isdT#U]uSs!)X.VKx\U[l6g1&NCi0g7 "]$&sFH,@!@9EhGyW+X}?g@$->VOV7$-y&`0#QI&QJvo\TK' W
Ap]\d)v(.*g*YH5G`Pp$NjQ
Z~I(9auk:JyrU}7qVFr^r6_Wz?B5( K2K0|hYVL3R#:X 	qr'RwC1C:SUPZ,H.2 XhpNt@z/)6MjV-KX:B'h-G<7$;RT~_mY&X^6kKr{
^{5AW(wy`QmjoFb)J	TZCTej(Ihz\|=A3#~#+<_<.P[M\GVE[jsaEa{"0~M#["c\CIKe2.5Bv1iKP`NryRmk*'}z
3v+u3s0y}2~3I"7>WH*t	@$ bIu#H`Rz3-^V9f,
{E(%$v*}	3xQArv`k^nSnbEO-D7{(j:0{1zF8:cz;J#2q%iI1f97]XTjwW%6sjBX4|#V&DUjmJ-JYcrNd}gOafV
jKYb+T)2^yT!C$CUJiq
=Qj<N4o gT'cdQ5#IT+%Lj-x
OjqsS;k!90
R\qy97}L2ZQt#fmk7&f/}(J%[%z:Oe?WE`FP=+%yyMtz_p*[*,L94f"kpHrztz+![QwE|1A,2e
m|i8xsmF{jwOnfuO=.2C"k1oUqbrr0c1fB-;Y5XVX.agywl5m{(c\R0O9;:j56NQM@,$-])#H+gi1'dBQsl)``4K-@f+z'y
bod636P#?M"J;#j]6^nw)|=xIy%#-,[eN!@ub\Q
`CuS0G#KrUk0T3|?U^Kl||4X0eJB`_n4[TGgi#}p?C5/<FocA2m"Ee6u{>hWIMh:6aRI##S^{DKe9`r`av:O?*1T?	,ype$.hr^TkU6Dp- 2^np#,8mLt\oX(iOSW%]	d[F<9rgtZi&~{M=%]gjg+ogyA)iQIM,6b6fI&UzF}7f	*F*?e^B605a$6QpboWo])':Q* ^qSM"h\Rb[6t!8LQ=A;zba-E?zAI=JgYWO0k<&ss@Hu ?-ogYgf\-U*n^8|E}~S/pEmb6yd?PBz3lP&L:CDmp#2E1ZJ40XARyw9_E,,6f)/nRVTM$-2&L=cFrG@	nm	`CAV(k+X6'}jxLnaA;d2-Al[=Md@iV}j%9y}VfD3LfF8tpjcBpzQ`
FQe$ 'j2Z't'<@~M2UV~7_vX_X.y@O7Ro
k;*4Mf{	xF/]DO2FX.&9LS?He*UMb5`-Hdh_WD.Z!4DNN_c52siJR>TLQf>)?2w?7ti6/"jm_Lz@uk*t	z@Mk	X-Gd{x;O\9$W(TQ
Mm|6aL4C:Ia0cP9'g_bhJF[$6AiiglZ/`H>L%Xo\Ta	2g!M%;'Jn^Jq,X2"^79zd4/G~h9BLfAX#I$i)Y\rP TN, 41l7T/B|abM3Ld?vW\_j#.x?V&e9|Tg"Y~_-iqj_fD8~-Q4
{&hU=u#N{SmS%!X#m
FEx{#SWg)qwZR9I|=W+,/it^~}k;lI9U&6$,4h6m!wtD6,GPnVVP'NS(z^M5TD &HjgV)x;h"93[8>_T737S`0c}cvk&kH(FY*@:LCCES+M Vi9G8#p`N?eIQZGR=Agh"UE}-$FKvVv/b"otb5VB~!*rH ,Rl%
L9_l#WN-Q@ZyTbv03cAu0bPf-S/ oa98o)QCQC-ep>CRg}Yk)X4;='\@5s=5\iUUsl8og2t]N<"o`gq$PDjTqN%n>jf>@(P&}:#AEA(2-ypJ~)]3"U8,~K}!YYlR`CN[u|53HhxvU(d[*!2OkT `CoAH=:^~e2bW;U4*;TlN^RQ)iQ({MTZ4gsZ:r;Dvu[DF*rr<;b/s5Y,.Oc(4Ei>e#4S]*v3"fbtG6~^nh'E0l\+gmrOd@4r.$;@dV@cm/	[c
q-&eb6Z,GFN*?amD6{^OE0iplh`FC<8TPx,#-UF8OirKS>O@mI>LW=j9iOiYU?dI14DM457:*):BJ*S\LGk1b_&lb~h8q=W`E~srs[rpG`Y2^huk6fLF=G4zO5)JDaM`c)wYM>eZ+Is*b!j	fVsEop!0cS6jNT	v]$uRPYd;u>COumefSw-&i!k"<ypp
$ku'OAeCb
YJ#o=<7/++&sIE2&;>io5GU]_>}~zo_F2J!qo/yD_Pj*N)T_zH	VP(s*$UD	[L[wY]_]?Q)CyX?^PNkBUHlTEp^tY]o%Tq[8	:K*9LC?C<XLaHzb7+;cWp5%h[g'nZF*l4i+Z!-~B*<51kYG>YK?HC#PRvNQ`:R0/Gu5-9rn~`Rr_8\cVgmz?V#<`ORL@}\\am!0kF`8214	Wg-ZUHm8ZAlSi7JdK'Vb=Yh;2b&W~$L[P"3YE4&fD41TnGx[YwBh~dMI,L5(C:&Vxa-.;`ol)CO-jZGrFnBa-L1xrfhn$jgD C#sgf.(UiAw"{AW[Ry(wI#6)	Hr{RUA;H%	u+S"}*WL/$gSk[lgzEBmb\sqaXyW6ayf/)%4OPhUt+N?o't'@=mN3^d2-yhoFZ4q6Awe2,mt"X	5=!Qi`cfa et5*3Rq%,H9 lj'
Dlc+2g)&,(|#N+LlSl!MD0xBCjV
\7<@Yh_#? k7=H|tqk..\[&Lb~!g^P\)k}{ohSs&*$o;u{+B?a?)e<j-9IK`rEVuE-uj56
t[dji9S.F_
%8;tr'-VI]\_]/#/nj4dQgcXi.mE=F(gg2z$:Cj02Ea&jYn&6#VOhw;x,~Phq0"'n|0dv(&_7|fV-4!d[d{`1__%k]%{7{I]xl$=X?5DD
3*-@w0hGfIF`i@kB :H'APkXPo_((rK$5N-RdcT&o$b9Rs}z0z,.OyJan^rR?ZHy=vzq-m34Y0<qkeB$y[WXo*,Y9XN;<:$~./*E	qo|Fi!t5In0EuX;K@.{6#'m24I~:+Y's>5N^jdPhjlkRMVO>a+zu.hqo5LYu#J+i]I
?gabD%i'*>bNVw]<yl~gxczp	4/(HtDzSrQZAwZS{^i}[w`y<jP}(rM[o,.(o6<g{dam.TYCTj>9S%+FL*KPOuO8. r9a1t.;?4~3W*kYG)is9T!{nC0!`}no%bY9}7bMy$s$AQ'ia=RDb#4F`sM XrM8XA.@vs;>okp,n5,z:A*SW	(7`FhNyi84
eW\:APivh|iT}s")qxK"KP2pEf ^	VD9++,x^3t 8poW92wTTN:S2d|U>@ZVm}n38!eAf5FVP^X>c-d`A|jjT
?~)aZT2}tp+\LlP.3].:4n;2[G;K,5jpwm?A`?M^i{8g/)o/Ya'It0m]9c`.\.||1OG{yfl
&GrU,cNL*`@J&>pgnszo7{I\u5JY+V;9Mu7(X+YIuy NYnmN"Zk?{Dd.^xe^0}HmE1:NNxiz'(~9YpAEkf=PjrBzg0~{Fc_J8NK@:C5*s|7(]e-?"E:zY4_IIGRw2o^PFBVbI]=CPo(z/5'@(MGm#nTzH=o5{P^^I[(kRGvl='t|rSv+FqomG[x`q{%\\IQg]e"TpLpF>VifE5k4:/#Cvr07'l[mY7qf$@k7}Z2n'@$	)4WGGE)o|	Gbh#KM;\1C#0]bVI8-zB]6L%,:B9sG@nCj}nqh7j1"SPs1CT#5="Igy5c{835A6hLvH"?'#	p=e?^xz(=Du<46E&;z5(}qJKjnf$@a*CDWz#rf0t9AI5)#PEFWS?Hi-}H%r{S5u1y@O7{d58rp%	j8!hq8Wyx^Bm!\|&
iwg82}E9's5	.(_2/7]GGcN<~9n7o<1dnN)I=t>?skngU(;Z,,GHy\#e|\Lv&wzb$=a*J/%9V	b 2*:u#sgGZ1IL6
;TYrW{x/\T2YBx;H6z;QvD}Z?Ya{.YT_YwdU9BMS%V,x##n9-!1bHnvlb&<	g$?=#>W&Mf4jkt5Ac'tvn;2CFj.>R%d{!%^dr(SoNW%0ASElFZyyv/y{]H\W'D($`D"a?Z.dCB{[z?*G0YK9QRkU&9LaNp}xSMPwL^*VWGVH3~ #HsOt=wm0Hsh#tEYSw*9
;9}B7[kb3~;[8IYC>6|)>-71%Cs"FxlD4=$e2A$ to;rd&
&Ib5:fPbNwd-szVF,=zG!E\/OD`2y}i:xx<[Rp2zAcr(wt\o)xF<Gd\iPU/fPOOk9r-yO+`i^_Gb<3%1/d-^>n6k,[cV/j{xe/8Y$FYrC0j&^id~CN!r#)O:}><-F$C'{2Tui|%F?EJ[D;oWe?g4;St5d?Hg>)8j`>ZMnO55Fh_vDcJXh6wn:IP5?_N17\Zp_Efk	+5DN3X}@<k7_.b<=-L2+{< Vc!Gs6dgo60_TH?CQ'DItu[xJ^O3qNI6[	NQvz0UG	1I*o]76;^-|B 6_!M1CFP"^brrJjcCi7sybO$`/v@GVSw\$Lb |s&7/`F\U`GU.C"{c:#q%P^H'z^&oR\<^j1yw`#\O%c6k6!K^F:OgjvTh)4&w}_	X2j {mT#N=AV^#5*EXf6da_PE7"#LJ9*J/	f2>;b(a0VM(4x#*3cznXA5sd|CX%(=/-/V{Jd+8LRv:\,4}\]879""Q_3T"f,<=oNhmcc]'zk#OKW1C"8Q'R_vtR&PLYr-._\y-(b94g|nY1eRrB&a1b5)&|JFa~?{F>y)o@+waKOl%>,<ahK[)B]jr=.@z%"7P^;YLMnQ+Bt]UggUd8Qq""ehH`
#bAb~-
+Q&/@j [+HjUu.b^xBdy}'EsROPoB""D+VG
];xZhc:T<z&hzqPT[;6D&K!Fe3s"Fo7HP8dXLnJd_1/QxJmbR)a?GsFZo8Wglb<~q`'C0P[H	=S9vFA:T@dC
{ClHn{!oM^fMv+7^3UGLWp;r[z$]\+4\Tf^&4)N]LfQa9|qpz YEUh(}]A)YX!Q2m*@1e1]d4py!p3B|"]#g/66*RfM']VhgCuA|6BT:Jrh>:Mk!w#'gyy^Tg]z	wXxW
#vf>1wW5x:]|QNL4f$4]cO9w#t#Dn+u+n.dh5PSXU1j;uLvl(&SP%FQm,> PEWw>(G`]cq84lOHFPop~.a@BT =l3;y/)SZ2tP|nq!gm/S%xL(-\;c2!H+C[3M|zBDrP:GIw\bJ{GS{ay-E-p>
c_+2,2>Rm3GmXG]PD:OpjdG;ZY9TQrufg^dgXmo`fX a{qT~&RX/cq5O>M0IVL7G`S$7b-mGJv2$3%_*ZcR^dNjGMn7HL_7zU<I5<	t_d1RrK4]OtclI&#d}!+/0J]7o@@RlyS*Y.'9,y#Uc\F!i,$8x[rq/pCO`d	k=*!?duX\xsIAG!hLsnx1g>:D+1sr:,S+fD>7re3WY_'>sSqB	rtL
8t%_q9 T._W@$2!EFJ:GRC$.IR.i)nt#|/}yG*MZ>`odsN"5w|XFP>8Gn17'tptcz;-2j>W;1 H t[h0jK |{\_VHhXDR'\%zisWWL'Gj>(&+Kf=O`@1&YFZeI!""tw;"-6@tPzO'ci!p'NsfouFR5g;#G3%|XMKh	VNT
=$m~\L}F@F4<uV^Sol)fR!W]-d?TOX.v5nn@:kFL#C&D9T_ki`YHI[y2'6:"EHd|37mh0;T}#?/7Nw"@gG97}f<H$oe@t>.7=Ie!~64I*4?W}"izXiakM4Eqq!RS	+7p1L}i0 OU6-nv}#RfS{zZ4_(XcBG<'\*^^yJw`Kt6_\He:`_<'.@d,g	FC-X)r}m4	
vX\ur:&aE9UdGDu
D.Te4!pKc05{l=c<{}f?-}4bE@myL?I: LtgFklBz>3\vrK6PZ*y5vFqi7mCJ"<<xu,p$i+Al:c_`4"GeX	w)6!uS9afTZh'07.s7K~Q`+J5t$wR}8-^Xbons"dx`RQ,n<^4WvhpONy2%?m^|QEQ(I	Ze|K$%AP]i6"EZgSrQPRn*UA?IRP&-,'/kktz|YL'(>BB$LbC	]cbly<{2+x2eMFsPu\=!)ysg3'>:.]
e-T|V_x&+zfjUFFZ/4hNJ;\(XUh}6'sxS^"[N
xSsm!`@fcJM!K7~IS3!)P{pzG>m`3%34A|2&bL]vYeDhLF#bkZ}Jfj)Yxu7$p!!53U}=c{ZnJhQX&Y.0q$9F{:\Qr;)!`D
Q#fr0[?[:_x7KkKFl1iJ:^7;kmx@"7&r$.Wg3xvJ^JS`\r{eGrCth?F,4cVmGB
_.6_6?,CwC2cDO7/hq\zM]5E&TFDs4K=lW.|j([\tu(bUlVMvS{aGdws4]0RgWhK9Zf).9,W5a\!O7S%-GB+<J*Ta\R'c-eGB!5x4KY<g~%,4(`>d /s;)Jp5Vq<[W+nB@0:JkX[|&a`qvsN96j,bx_/qb.Klv("b
.Mv9!74RJ"M=aZEP`U)Wvi=[6FQaq59|NeW%9Ui]yd?]./V`{;#cV6jnMac}7<u&Oi*7B=xkhXY>V:}x"gKevYsF^ki!NsoZ%B"&C4/x"<QP% ]}+HJcfjdvP*YIxi+JUFG|?Fk6:Ub-2V)-.);3#@MFwgu#Nj$T:P<y'Xa|Hq\2?|:?dZY9eOFK[n0f>|0rogh3V5(YGr!p^zWzid'I$Sb!lb)mx#n98k4N)rY]m"-%wL=EuNr`K}}RlZcWV*qQA+nzCLb.FND<lq]a_PA^)8zN9@xO2_oz)w&80fi~QZ[Xq v<YSX_#fESN8H$iV4+^vTe^inJq=z#+	0eThxq>"TK<tM+&,.)dT.gc~|"F}"HYc?h16	)BgRcX);lf@3y+[MOFkU;Yl+UBuv~\{*NU\a<%}E'yizk(nr>A^mAXM!~20l`H4`Ll9&2f=Twd*9/lXB13o!/?=ueV_('5/RN`|y< \t&#(/'"8\Px<a:pZ`*<u5f}STgch$LDCJf,`m(K"PnxSh#bdnt^m+tOwN})3'_uRyM@6`IpSmw"GJE>MJ.8Z~UQNVlX'>@Jo`P8_2K&kaX8az&({H_,/'Y
	eZo
n\zXre	xA`4h}O7Gc/_',!TC7j3YP;^ggD~58UO<L#x|<QH?yD<?]0a<26]rislJ@OF7tl@.S_9g+V[31F".dzNR.Ex*Tl7tJ=dch*7#t`L9n~1{qjHy*X=I"1L_@Eucd.@^F Js8cw`@a?M_{`ha}.,GO8JAg-0D$17T8M;|'E"9[Gs&FLJzOtrIVmR%iTiz5VTg1h)Ij'6:}zdo(JP#;<?.Ce.`0X$E1f!z/6rw}E%Rbz
_q*c5vZ;h^`=3"?7%]OZ)0U'a4*^s87m+ fTG$FzQ>~ hI_!O\\SCV2O' >p*ww0YSQB)cwC@!4nwW\@zt.#hw*c{.z^1_Ie>kvzj!goTU|6)H2WN0&q#UvFV%7BhG<KI]EbfiCTcDWi66Yo^kg,bWmA>rt(vUgKYAye8^>xL93hzsn),F9[(p}2Q}m5:@;lW:/7QNl:W-SnawDFi Dw9swtnK(c!?-&	Bc81J'w9<T={S.a6i}zYym}j%dEzvt`7)8GpO[UV?zg_0K!S~U7@(Z),vh=ou2lq	=
%G_
L:4GbG{cZC6D[:cNw|YlplXWI}ipgi5YEm/[X4+f+^"Pp14Y+stey'}mFIBoZw]D"Ou3Y}NiO9OA0-TeT~R\ZLapvB^{\ZpSAV%zQ?7]pss^%NNl$@"?^iTzW@XP2{:YwjKPSzzHcXFB+?Pk(fj0T5^~iE,~E)s]!GMqv=^HW!#>>wf*x"q0.J_IbAw+~p'^l YrK|A#Tp<;`6.4$qU>j>q={<<1ir5s~I&4>)auX5J}D49Q+oZL Z'sk8/sq@TC4Ybt>u9,dS#sJ	P,.GA9y*_sgO5LYI8:vM'O"r8XY/_eKP~v&-d"$xW	k
#Fp)sN.vbulzlsZOwyE]kFiLH
7Ym@X!^X/fR>5sL4N;dapu! =09_' >CV5go|!#Z|%;PCj\HOx*{ua`lTGQ]7I$	tIk%T^U2,rx4LXZ@)0"G"35fR(D1AKQ2|ctB\ruPXh*:ePSu;42RX>MuUuZ(B!rH3/:p~G5c'Be4@j>[d4_XG}CK:GyE-`3&`(3+Wkp,]Esh* 6&;7IF1|6'skpP5]0NaFK4URG"=$3ksY"*,7eN6#jccLO[:g^,)^^{!ijnjr
(t`kWs[_`oyDZhMO*@S(-/U
"1bB
b>0eaH(8F@[n%=~~tJ=4mg	tvAVko$@9Vm0yFn0-\b4h!5lX(	Jqj\N3EXNSvig Y@J-5U:VcZ0[]#Je}c%seJ	%=
n|Kq}0W	B[fzu%$5_c@	yeARk?1XPbKEqBZ.PI/8/]mtINWN_>3K"nM:91T>z]{u|%Cs@*	Gh7hU,O9jg64n7OL:-4+QoToJtV5)s'6<S1|c++\93cuu$}6P"I%bjF(	t<t*-'P\=Yw_t^X	JdVnZBHN[N[Q7Dp#.I`\cL{?*8*{}`Q*)5>WZHj%lE-GiL'}deKSkd kV1SEeoV&A8$uA!dE;&!7CLdVYFQB<a(`UBn!j?"B}jKh"b=L/letr*3NJn6tmMPlfby[B$IQvvB#oQ}vL:U})<.+Dl-|J,>~Ap[$+e#=raex~0Nr![qF+U/lj;$Cd<l`Cubk
acmwgs<wA$ }K('_u516~gDnPk@R1qD1=Ld!xkU%MaWM4SbaYf*U	+!Z^6!mQ9NSl0F0xx[q!2}s>r[|Bh%jg;J"1[|c"=]J_:bf3GFu{]O/_/W*K]yqSI%5P.L0vGV\Y66V4P b{F}\<"4YS5SM^CCrb=[[[katS>$9eb|9U5O6qQ*M8i55:%6O~VZ561]9@1IEUy>-OJ69
br_dP}2@RP-**G7rLoTKy:n5cm=jWJN&Xy2x:.X&?s D
3vajW}Dhz${.@V0oHL@m!j&hes2^:]`M$8Cgz@S'a[n-{xw!sdRh'0ABO_WtHl04_P0.fXSykJAW8l:zPmd_2+/'oNAn84rc~v	zcB1FMs)J6~gg<X?o*-dH-Q=-EGhNrn\?E(2d~Ksl&0H&ekcRj8P'b3"6^LPTvGb tms46XB#pw<JoQpf!"zbIoy3;m4\_,M(+vX8+>ImpQgJjT'0@z	J'5&)*Dj}f*Yl+|x0jUeVwb":+(rt0#tj*(>%J.37kYH6LI{87"{gCLL	W#OS%_`C`.Yf0<!g"ZIts
^#2{Qg"^h!d`,vn'pPrK/d'bGq\}em2;0`qBE1;W8]c=C`n?lPWg~c$8>HRxffQ2HI*)Yy?mX#d:M${o~"9&eb5W)@b%
FK25dM9)"59z+^dP
	6])2J^f({{S1[hX`EUy,]=_\SW78C$$d=4/-EB"k3E!&jr#
rA{4S
0Q`BF!QQ""#`b@Sfk+5k$^{\2N|suRH9	x91p;Q0y9^`H(@q7TYgGXJ{0rE$V	N[%i.kI[Bv< )_Y${G,y*=kiA76F}n\/)35v{p7e0bJ^g9[-%.Q7v|JgqX`U3!KVY]	`(	:*P\,VRa6x 0+Y	ZA`TFX_|EB$D@"S\qv=I1nYpa60JKvN
saJQ<8]d\|gjWA/3kS *Sj	B^U?=g4'+' A%eBvz*b6mhIf'K9>4@]}7lEensNQ-76q BSAhMj|~_?MdD/*Mtz_s2%y0+(:ACBCsQ%t*DiZ{9:^Q*4SCkZm,F_/ZRlN]%y\uf>b|_<X:-k2sZQyETYp<dyIj={qxC=|&iUk"|K,W$)flB1e; {5}c	LzSKPcN[32FgmHySlWTZ}/!&?yWi9)]7I3HsJw[CL&+Bw{:*tJFQhu~{?J
8``FXSnwsv+!e[&Lq	}Q170	a{k)YeTT:%/Z{GKd}XP_tv8-Oi%%o/'+dt^|mne69\_{c{rsPZ *u}7MIyh4p.^}"(ql7Y
DD^ur&{*]u{FGscZ5|'Pk5|8([cDREjD7*]hya%t",a,	?Y7TT/Qj)]g;h`tbNr<2Yz&|)H$thtM5dj
7e[6Lbdlun,^,;8|k+T's*2@yRd:K-K;CG.rrpfB!yQsOFfU>s?gVtaCMhCCP3BA0Q["wtLijS,1BT[7"l01`_w6R\M^`Vn[4.<)z8X)jK.!
[VN:}EKB#Z0/*$ACT .cuBj^SZv`R4#=#Z41QAKWA8M:knMvZQ_R*Z'lnROqt2lVr2"DW7P`*=B(u	|X1K#ujUISI=WFQP!U;ndx(!CiE-$v
TaQSZi/T>BumoR\#E]0 #$Vv_>/;s
E8+>A	m@zz2#VjkwR[ *oy!/V%m/YqZ^uy7ia3qK1bg7Qg/8VJRo7WyQWI21K{^+=Jp>Iu] [V-;|o:B fb}p}U{Coh+-:`j*XHMLwW:RR+B$y3U9V-j#IMt njWK7>3gR0(Urg/L}/ukDzI@n}$Uwxb*#]/iOG2u_s\lxe!qBEJer2l7$-`=cS?>b}13q~7g:;<'jqA_%L;{D7hp9XW[r.>
{</
4Gc_{1bQMmuk%2? KnEeRt\Li\u\3"7xy=f7wvanT!,5Q|<b)`[c1(
U"bA58^z
WgNL
+&/Kt,]#'ZWQFoz~!m!r15:K4W=lH)Yj,LRwHaDR}3I@wFKSHUnH!(X9*pWCsp! /"N[d%+k<UA<?\FSjXd<a
5DI0$;WQ3mK	)Iw}*vy(+i7h~q(#a:/KYFNf59%+#l=
HYm) V<RiqX@k@V-:2NC-^tV@r8>uCP>YY:+Q({G|]7A$;T&%<bqqKH_zBEg;%T?r%`KE[YyP" I8!OQ0mRCkz.K*hre\4c#4C|'-Vn]hT}--eF#F)q&	b>t<Npj%n8h#>b\T6_&=l?5cpUO&x){Jx%;g~2a,&ahO"am:4;\*&}e]7sWZ<Q@op7?iW$K"?CVpKVeNbdm*69Rs\&#*SqZ
XDfH.v!(X#Z<l(Q'*t}MMh)j9ORo@aFP|RNP]PJjz9SsXU^`Vb?xPeQwS;#ZzCiRdE~"mhk+2'+(TZ.yH964Kkm-.WB:K_=7p!zEv=5W[(xk9Q!qKNK.\jnN-Te>FEzklm3+f-t<':Cl4"kW4n?!1vNQ-P.({"nEL@p{x6Dq[t%=i"*p=4DrLV^j}A&k=<`4r&W
$H]ayFS>NIq-0!}2N#X)-qZkz:n<S54L@3!Oh6i%),ax<3&kXSXj~(R_cpgg*[UHesTpj%nm>dCJlc3=bu2p|b8W	|/!(6f)31x)s#r&6=CS6|m8{wg1RLBenhm*(1OD^tS,H[P=oaRY7vn6%,wK^,
h}!Jcm%m|.3c5S:K\^61bg*gdH=\&`(lc}L;HBq]2>B?.b(?n<-q;_vd`*5M[0HK9FjV;aWPq=VyP9}[Z`pvsD\#`mrDe&4mx6E-X|w7|H HbR*Xh_Un<N6rHHMwBEaK!,.1Z#p9Y\aSj#`[;PEe%1A[VkC|R|FbN52%mtwo\ZM%5.}iMg'r!Wg*^`({-J#{%:Cs{/gM:v^G*d({*;]VVpT( @?v.Oyi}&;<nhe4P&uIXBFGIjim:q1xYp&8;$k[V3(_Z6V1 iC=A1jD^J2hIa#HJc13(0
qQBS=*:wf=Es`T3Ih6P($KwnGLY;tt3461v
XER1zG+)|ZKZ-j8	w/5n&XaQaW.`t&P#>.cF;5Py_[e@"`ISDCk'I(Lq?zzJL%Ihw4MmBs$.i.8pI9@!+\o</hwnK>7y:VaEo>@)*Fg4<#
(h>nh+T8l ~#OjHdY~1Z|y:<
5}qN%s^T4uKd1DM3MgnJis8kkIL^2x:`caQIt:F].>AykYeT
taDM[|8E)'#04U+Emz!PBmnMNzBmIk.Sv7^\*nbi	"O!/xn>6fOjz6
OLxtgT}h!a`<7K,UtgBtt"(^$	sRej8]@_b7y4<bb;aK*,{FC{Z&jd2$:1+7)~>_JX,1yf4Xt(KmAS?'B
GZ&{a9nV n(sFAygMh>C<nWNBp*S)]7zhBDPZNH5%<)Q@tKp]
wB<wCY{!Gz?',!iR"5#C=
*ww;yie[*Eq1!9qS2$u[Fq}Va((
.D\6i@>DV4[:OgC;#ND7~|Vv4wy1P5,49*P2FDi2R)_P[(~Nab5wT/= =@B+Jb,s(q,L,( -YS#0!8)W*MEix}NO?PQU|kR1f)lN$y%B%Vgm[T4)f7u3%xNy0aVc~|i+N#E1'D7+fb*h}$JiZ$)@<6H7avjcS'aqzRZyLhT{\L7FzYv7's!"q4i3#+@^DTS6_U:B(O mR!XD}X=^	ACr]pn\"3U9j)PH-%/'xkIbhn]`'hi(f:i/ (,rzvEj`^1x|2@;zb"07BCoyVr,P;/o8jPw]tn?*l|eL1!)%ncq`b$Ks+>C7(
i' Jz4ew0GGtYtr*mlJ++'
N:O3.~|n<Dvp]U1D.z#}eqe}GT""\zHxKXor)W7
.mX<9sZ0zsu*pTU+[wY{N#	k4x$hzLf5;Mit

r>mBg.:^jeDp?6)+
y9ZZWv	845%DYP+x5REAwsk]h$kHOk_}k~;br`*qWS.kE/^Kdj0s9`?;'/wVqE:rO?M,W{M)3+rzK3-%6j	s0~+E.95a&T{Hw	zyiV5K&R  N$`kd,8T ISio*&vwfS3m&8t@rn!X(ejR$F1^
7h2Ctz439~]EU!t/<;ACA-y>gf>w0B>>
D[6}[m#xA%oU$? RWqRD"3x8k"3EJiYH(qsYy*oK:
),Q=/:Lx?.\TWj |Ptm't.&6O+h-vSXBq"I *KJ.1;ob"q?ku?ZO;%^CIp{lHUL_OV%m`\_Ls)zCW5k0bv#66~_A|wXLe_-QV{qU%\
;UHCOhV
WnG?YO\jQ_:Y,CP~#5FY'Tx-]))<*vWCl!fps3@\le.>"YAk,w9
!
S6gQ2X|C{	P8=\pjLw(X
T;YSiWMl:C3 $Yd-Hv9<Pbhd+xeG?MKwGcojd&}c}cw&3mHKd"j3Gz"b[iLjro =Bwwh%;;]@CrBU6y$yui~]-j/y&x'%?9A*6?O1M!
eo+;d&zEi/33'	|LJJ@Qvm7+6~]dit$;@q@wzKjd
%i#Q9+2t0q+o_	zBajn+:JN9_V
Y-G|tf`.\/AN7!-f{i&%bSG@@1ITkW7liZ'.,f-;N,]SI#"mRKdSSqC6:w0%8nZ>&jk]L
K-t1_,'
:r5}/$iJ;A\T?z`(+`6	Zyf^JeRy'=<Yb
z..|Pqr1U@?Ezz/&6 !R<R0)W\5:^4Z1,Ib,hznafW'IG"m@Ll@U`#s`;\7e&Wr::ay,pW)x}*:?f<tL0Rs l:EgTl8Qv/f1hvuMLl`Uv7S{4<XB2,r[71L{<
]54UJ-!cqu5/Q%jY>glMX00~TEJT3Z<GRF!i"DI.%w/!tv7(#S]\=EF$>U1r|
_C{B&czBUH_:"C[j}.R$wHa$Q"OeM;F9BVtCc?J3$wn),;rB}8:\?z{UV|jow-D#60^mflH4>x-'A^uUA6pxdQtu$t!~ coI[WE+"$V[j\Xeq/84(ozyb,n$wz/?](XK'n3'?2B_vEnAS.p&Q)vT!T8Dq-c|)HTgd'AR iHXmNwFb0l%u.!Sy|`_L@qi~>I|J-P*_-YVTwK`w8lT!dwdE^MUjf`Q\Pu29?nj-m[9~-4l&=R`@y&g%X\Cu$Tqjod}9Kx!
.(zkE-tR;MHH
z5YZ
Y
%LpL7q
=Lreb+_ZF:K~Ls>A>k*/U fY!y;7A%:)>G`10=:An+:Gri&W8Cl0nTLCfVwK}\3,XJD)
Y0'tp%idnrO.1\YL	>yx#wbWevDyIyo8uNBMw\f~s71mN"W (q=*}W4:Tg/1\+;3-gdJ`-=L_Bc	pXQ4	
(DYA}{eKJICc3}tVVO2~!Y(&b56#](Ry&]A2Iy0Pdx[05Cq{h+%l*->X^|MbE88#eWGp#=a@g3q%oSVjSh|8-!7C%$ha}sDI[[E,aX@5#i%gIr$TO^E\(/^;ph+2j?~?`M-pOa<RrNwX!K4Ej[Gu]zhz]D8:q~G,<M)e](q32G:&1;G4%!m6oOm=d%r7NByUf}8"H'RGWDyQ mtx-8p\0u#	}NxpAb^1)$4Q;kC}yg>A\B{lkE6 -5lgSlnSJ`M'"Q}oH&K78/5y~/oGpTD8A!xMp+M6Ov9nJh4W9W:h$3`4XP-VMl[L|ap>Wb>1F:.t"vE^fb$ojIP%z 
|nfS9>Ix-tqs	]z2nZB[4hFo G/co""U`dg#z+W!0>Z'XH5vu}=~6h0n.F,*8Bo.PSW{.h1Z}$RK2E[l7h3q	N%:\QGsS]bS+Z'I)sb{p\be+<7/Z|XLW$L6ud4Tw,42X?>5a
lRCs<Pe>MMX5lF06o0q(*$u"vLWIV=t1M9`{D@Zt_]xu@MA:W#w=gri'4~GS$}$$4fkhddyx/0<E/~Ul&c,@p3!lWlJru;hbtu_.6Nes)\2v5%YI0+*AU52il {V'U28
B6yEXoz/=FHj!VJ2t9+Iwn^&3&&b/*z'"9YD.v4_3m6\w0qZ_.J48i`<_8<|"V[uU6@`WZVa1}aw7'6,)h",M'_C(D>pEf7W"84h,E{$/1L{A(&'dHm\r{A">W_X*,"jl^}ww0GeD.5nKJxQIhNEQMB{%@(c%{x.P>D>B3yI-n-}i2O"Z"]+T+)Sj=O!wjs CI
2N	5p;;Z0VjM;L=Si0R?J)G>WIhyi//
>i(L\utQ*-wl3^OID22IR~`T!< @6`~}Lj[jO"Mo3~EWR?-uh[8[*%72Z|'kV9$6MgjUoHm]+C&U5&DjQuj0y%DBU0s[nlZEuCBLycOjOQU!02LWh=/et$5Jxf&{a%+$NzpCQZ7]qD70Q8j"Sg-6P5O}W37KO|)D \ULR+_eZS'fEnR_{7x=z}|n=8LVmM?9Qn	@&P#4@zBaO044{U>%xww..C{si1lO4[I7!1XLu,qcd(C:_!FPi5|AYB7E]8Y1s`PX(HS`ln6-GJqJ^#7Z|Vh4nx*HoF9djO;@IuXn~EJ1<f7%ZO;by<*c2;ghqZ}=::~Zo6P:j>A=j+aHNYWA'UzlT_4Y>o7YQ79~5-.AFKZw`<p=jZ;:\Umj^%P\lNI9.U}/Cex'sSe{h|?$w l	V$]6Guzo`^Aa~*wU4<n6|q\-mG	ub u !CNt/A/N,LX9SC.WT/%X)A}Xk4EW~[``U_IZWTa,s{na+O{6yq4?rMuy9i.B=A;_$XBIm[kKMI%CnzFTy@6KMzFjZHNDca#q(wT!F0>zd9%o)<(7]uOneJs:&UO/Jk]i+PVa:$o59j`,2!&mT8/M2%^v4k=)=o$(OIKUUa;+ii#Eve!M,Wz`w*AC9yOUDy0F}J
AC]8jC:FRX6ei,E:l{vWqIJ!XqL*W~IO0<^pS3G!paL+	Xy^hw9	4c~IVV7GX@j1\aGJYIdEsDJI]@-f=*g^}3Nc 
k*%RT3r5Z'X*Y7#[eM<nu&x$	^|-V%LRxB~!@j%)!v9P{-DQH/kzj,zc[#J6~O=s:A*Nt	Y\/c%+\y:e?Jg'Y`fj*ta`{k7;d,LVUjUww%PE$E&C3IQ(O1i_hG]L+TvsX]uwj/.0QWm8u>kQRrnU_/8Dbv#7T3QqHa;:USt0:abs3?4`W	nZUv5+3l\vy_OGu[NPJ(Z7PDJ/Wm>]X_M>\<4@ow'LG7<#TRC#ZwuYAK+Fli7Dky.sv?5|Wvw+/upje1^}5&kM6
## ra7BQU6Nl9%4T{0E|(%iLXc|oiC'$cQ*Glv5UzN
SY};{ME/1?k`}l$f68"ua[	LaOJs%YtRGO}lh6',%XO$ W-)*@gqrbld<Za=RyY8_AX>$\$Mos>I#6EZTO-Nql^etS:f$La+	Dnd?i PL-t+r=6a	\6pv4$!MZA
Q$|eb@gtQT[kQ{9+mN|fX<k)bA}FbY+sF1gp4@	_V4dmqI<>v#%`_ HkW_tY^&rAue+bgpr?mGco`"uVBQ<Yz?"I\_|]>UM~nDlS`\;KBQ,}~+[b,;PPN9H|)x*ku^h?a9[?w2p&Zn1W|'7tXOs@(eniE{5.HsOE&KN>gu\9S7_W)>Z v@wDcpkHqm#6=ug$|x(Lu(_X.K9lb`}{v*'@"V@&k.,,kJw5AP37fNtS<q56:QA0#q$mJfQ")ptFL+Xg)wF4!eFh)pwZq[cc=6[
xO8e/@=fGk_3C'4Xnyzl!DaBRJv wL*vq?1>c(UVG:jjtsx=I[v+OW+NA;KFf[Zp!P@|u@34>ps?Y_ .3Bcx#IYOw;&9}$9#;.MkBA,IK,<`2Zt%kwK8e` ,&R~syAXii@("YWc@Gp+i]WjZ\k|?=Z'S V&]Ue*$3qjAGpS!D046O
DW}X_Do`[xPB4W=2uUUI7,`'[fhaKLg4`gEvnD5kP^wtz`0;yw0m,q9uAeow[W0[hHdDku>%8W>OpU&8$r#5BB]xB`ji}u1GHW!PT]I/_#gI*`8hdx8.%iB~Z+5;Xy}Q+Y^Sb2:[7%&,>T_L*5%XJ<k4gmr\MO1Na/nN?lTV}^'`6P)BB<]pBk4<jr3I@3{ #&6Y-l@(d!vR:\7p=<
@O^\_g9jx+MOC+Pb>UW?zZC27$$y`jb"Ea?R5_5JL8VM[R] +ql"j|9G`*a'R_1IhI({O%X]+k4rar[WT4O*v,S`Qf803lh:SYYiRFEAbhywkmyZO7t}[a%!SW`|ct? u_"UWgQ^A=MW^u&cs2SoWo["XD1CO ;!xsXO;.a75a,-PzxO4kbJ;.U`Gui#,nw{')^Gpb:lv)Hl=nvbjL27QmUW	6/5RjYSWha&@T#!1:"vQ_/9lCQ]AVw1qdJ.0~9-LWHj*5e<)PJ?'6,Nn1^;oam1h=$HU3pU)[fI=.c2Pr
:8]l5RlCI's1wFV{	z#d%./1"@N@%C]~D~	jy6,v}NWBl%k=z!kqWUv.zU|K;L!<!?+!dojzFE40s']r1o&(A8zse?B^;X[ZZDv~V{t6J"CVB+;JfO8@FA l!N~}'sn;kZ:o0VK7c"0{D`/5|[?6vb~:2,k?5F%{aM"Y.t0Hp"HA"78(\>x}kE}vZC-Xi3sou|+l]	Q%I9\oK
0%&vmt;u{rp~4x<;e0EJ^{$+3jSrTks@zYJA[r [:P|1mMm8c3UTsF<T-<%#]V8Hgy{3fmf13V
56Kz!\q1d6[B_,Xw{z	?1Baj]]|7y#e1S_XN1OSMK9V}<3w)`B7uba)5r.N_>$xpaW`[}lZ:}	.yFE?;aa~rH:UHZr}xc~?#Q6kxHz9l\DzfrTBUd#g0W_	)YLPp=ok`00\}"-JH&0	b3!xwmw:=|ryuYcN(kxHDGE4a*GR2mN{T@i"MpSj1fk3	rBv}0^Q9{b<LRll%>+35Lv:[rR{
"}QP=kQ+GqhxEe'wpl2mQStM5(Rn`ZLZu\+5T&"D6}{!BA
]nGZb@AF*c)&@%k`gQBtyfYwMU0E7JJD*DSjK/YKeb(qU*g\(Y)gDu>:9zX-+U!2ABhIU8S%_sB:!6$&nMq6-8iK^Of<;?nOAs4Uq*Hq3v%?r.#\bacQU[j<&GQB=H&F7@Ty|cGM,SYVQ%@kZ:LJs]Zj6+CA?}p5>(7$C+Bj]-=g:52)QRvj:JA^Ev"8LC80;;	eXjIq(j[X{:<}GR8!L2a#m28L.@Ehfo}*4l{E>il\k/J4.X+L
"1LP|\Xh"SF@_[yngEr9!N 
AEo~k:vw6xbYga<1.7i/op=9qMH.#?v](o7XqNiRD$l<s%7D&n5TRO+MH>mAO<9AuV6
xgSF>65,$7.+<M v}:Yj,!3%H){&x>FA,;DLRZ+ fEt;RP.|a%Z\%-<z_(LLB/W/CEWgq&Ehk39	8|k<C<JL!qNw8oS\<4JBd'!\<,YYpZsj,+"Q&54D~:TBV1BSld	K_!IMYo4*"V5?[hs:{7E@|'PHw7w4(qbNE<iE:)Xq_.t~'y:TiD`(A/sl}`yrvopRg0nsI]C;lhKc+?Un3zD4'5qB`f5(KJ/-=T.-Sisg_i[6w0D9bu{V(bdIpa}kGh)Bg?K.$.&y8]<>_V{=42WIL.l\hn2k?$>5lK0{QN(n%Eg)7s Qsf:Ee=&0SY=`{{5\0,=I
ufCe.o#u:mVGJ3M@YS^k/%1Z$n$In)|i|8Y;94mjRU5Q[3ji)q-cZl[v7Ue6W/-/]O	`Png0SotA.3q*^\uL 2F2z2IC.(U?2K9-hQ{)23Xstd%x'0}19"tIXN,@SqP_b8@F90kMlWk()6qQU{k/(ga<>*Sy?h}V)zScK<llx3GPJ@#t#<-rT@]O;Md,!"~#G1;t5|b.PsUE\GEJYGJ2B.cX]E'Iza7Fm][fJ"0m@^w+7=mqKc^N*M$$?}qb-f/}Gr*%
1^x+F2.g'W?bRcE,cDF+~cob@gC\uNKPBF4m+^" 49![Zk[M%oQd0O]3%A{F,K~@sx*Re^^7+@DIPlv$dAPc:ROW_-@mq	Q~pbpL<5]oQzw|"!6jr~dD+k/u|W
:cI}y{["MOn=PbOdd
>S S?\S-|.Q?E{R{h%rlX[YMCG>ZXL0})&gWE4T,pm/|F;l2,FA^%R *V	%{ %N~0z"=f8:qcT?F9,/h&iZ
FO:MlFG^4 ^{GB7CN(U
_^WPH^!xnGnN\(yoP`N[JsZE0V CA&@]G0v60)O=STU* N-:].xHH]hIz l^^| `0Y$[I#F+~x{;VA;L%lN$^L{z0$BWbgI5LDMeN)[|RxHp-gxWK~<B^+9#b9W=tJu}
4^8nn(~W&fz69.WIw[?17[b$&V!avGY3{-:-+/R~j@#ueG3V?	pqi"2Z*Ox:K]79zt.h0h~xvA=gOf1vrb>?rZj4DAOblzb?|gw)F~n"hcJjX?9r4?X-	.b6@3SdU5&tHrum-(Z
;e01ug';}yx$5RMG`yQ'}h~Bk_U[Lu3! k[PziINOz~+Q2X}_EMPf7r)3< _2:u@6*Q7^M(Es{v4kJ%vSp.)wVe^ \_1bdB})RX&l1|4, S =h[vh<z9 KRB['{!DY pxOXg)6!3K{XNExov"SR'!IG-fMVK?bp]]%1;|@e~11  eG$1m36v({J+(X^nz`J*$V|hrl%Fwpsy,$)*d<vXTBp`6/^;E N33I1	B61PuhwaUC>%0+rHdt	YVq'q4C)7|~9Meg&"nN#n:l2cE)>R*#u^Bj4;q6~[,B!LE i!:(P1G{SVdOcZx>^/m4S8fM1UpXQ>A+)MT.7Zr:	U*0{	rm;ZK0C4Hu={#NS)HkFrP	y2I-"k_jCDNIF3JF1AoDB]( ]l:*`&ZZ'S>1Aq_HT;te( g[q_Z>)*6(<96AKK^9vEkA3O?W:6gb*%1(3~R`Ln5:,>s|ZAb1+
L&oo{ %9E JEMdLTjxpjhQyy'pJcB8 aE<b,tM.z$Z%FokJmVJuM7O&f*lC6*9Z2!@CnK-Hd`TyvSogxXJgJ\#44 F:51'83KjsH,Q8\X%|kT"tvOm_N){}8>;;KcMQ}txZyRdAgQ+=F4)MjlYFO~G4\7>4'pA'w.KOXd'J\L(Fh288\J)zg	C`F{GHW#_F!/U|bpp}8Ut!]*XwQ^Z'>F [jX.P1:)S#!ZGxx:uNhv!:'7',$H[keN]\j| }oY)]4AO~z(3,cOnlRb<dp	LYT8?W{T|9 <-*	lT89AAEolfeQ]5)6]FS'KWV@9]wv3z~-}BbCti6%m5Q8IJw9fpt-+-T/vRg{d4P'#TmjbWVH@WaR$Z?_^iG&d@	BwDBY;$@j{A*Ud"iC6Tgg[::T|K[NjBnh?ec#!AiZzvXUUcL
G2I,G+.T}Ty6[w	eD	P0].cnkhl2d_EN?\}F]'1~Op@I</Jq3Lm1{[?%?_z%T/qeqCbCnyHQG<mZ}6z0qfp
l:t[+Ux[F>AMjS5Hko\^Btd_rqFDiheca.aBa;_H,o@V&2!;w6*^9AV1;#Q	#`nFzIK/ju\;@dQH.+Y,E8JSA

oD*y!h3$\>J(vkMe}|CBCdDwL^cx~OH=n="@+${Cy}!k(3Zsl|81M2w?UnI$TIwFjxLX]8,@Tc;7.V9s<^:0Rm?#Z2m:Jz9=1dHnDX,D2;vYdX*%,_Va%tXCoN (NM8h;)yqRU41M&m:IG=q4cV(DJ_1V}Ck}wG`< fa+@p>XV8JSbKDq^c"(jiOF6 \Mc=$(-!DlPk&ikX]zqY
x>)0mY.U'^\"a8(oPm`IL
^rby#)QS#csBq2CX\%gDBF98|.p&xL!Aa|R.h,S-=m+9
u">BT+FHNPAXCPl#e(,p]	JisXPK9;aueY@L<z{$1pa -L2\4Sm5d_@0XqpDkP*E5,KY*DI5>Rh{$q[xcxcj1U7M3k%My |X3,M=JUluv''&ek_pUYkh*tw)ht&$$x/vy6j#P:~9_e/WeNcqq$2(Wz7!6?	D| />5M	|bKh<d<X-92Rlrp_I^]J[t~K|*At>bQV*zE!Vh_x:#,2(P
>Ld.(chU}c1f,$nbDH>sJ=hj.Jp1[NEJ?0hW.PP-RZjChnIK(__@.r_#JkQi>-'73J ZBU72T3rW7%U;`}-.)Hy[i>R_J>9hy"#r@q3iGB']7z=-lKB!X@ k\)#uDFao&pO;2 cL/Z?"$m"xkwwr=3\	mUa*#d.:T3r~N6G[*_]8hUAB#R4pX6Yx<'#*]l4+"Iq!M#BJMI8S^4@"~c{>{T.xnTGR;%~.+:o6Tt'vO1 =nvO\\m@;ye 'c9==#}8[K"~*pKMV6'Q@/dM_dQP1E	V>n>k-88xxec)[+HEyNM 
aaETkUhf%-<|%P{^0g96ZZs TX`)+oG#w]mQzPvaA\R2y+;"nzk6O=:\DgHhV9,L^ce2zDX'yxJ}	<.<w6:@380\Z_G?O ,rB`"rAbM>>[ZCan3$/j"N8t0vS/m7WDj
q;"6A|J1{GN3N^2xy|#LTT0(Z*MjmD>P
GJfOZ'4csfgY13dDR?&+ Ha!]{&p}\:(}g 8IRhj\5TxkaJ0tQ3@^~ZGU`WLR]fr+\5{pSmuO:K|+]Hlx?R?	PCx.pd$\JrZ#2Oo>u[e/Ty,fX'=_p#p"WNQrkZwyP,'==97zl*Z%k:9aF2 ]p&_.gE*:Dp"mR;CUN3L-PJgGRn/J/Uh	?[S6Yt4q&'Dm'2wP@{`p7dFgqSWJ*>	'n?]]()T(QKtD|'Mx;;HOW0%?'>%zu''FqC,]wmXH	J:K\ {UqK?F>Z!Lp:J683$1'Lyt=-+K})\XE9DZvBml};&%gX(naDqnGcH[r,$iZ*}X>haWZK,o2*]-s4{0v(Uwo0aN8\B1uO1&-g_,X[	#sB#+1b_n|V-/zb(_f]R}`
41O{6],+/bZi{0p~b6Ajog#m=^Qx	5W-Z<i#,R$% fz&fXJBR*w2@Kkr2w'rFB"u=ZC[58x31)*!u*B?"I`^bp)c6
~ifZ/e=9)
)^n&qfm&#G
M,dUMl	[~A]>bI<aR[:>>[+3RsCY{?+AA-<Ytke`;^"XmHQ[94?2-=l%G%fki(ii?b3`~`^*F)+PC9IjqQ_N5AW2Uy*	v%;b/~?~@WDJ4{8
I"V:>4fIX|'L}nG}Y[ppx4%N7;b% *.HT.f	4>|jdIXB7/AJ}"{c/*5;[eE9*4H]wAdPs~MK^G~%8x &x.=*KjYZxrH~X	n?R/1w<kfCFf^N;<SGg#a5Ey;8lVm|9_NXSM';TV(HHZ*t=&0<6Zkw-eS[/qA'{x4f*uawnf\pw@QT	Ji'9H~$'DB>0+e)}ZIbf}6#s{qu)EOV%IcvwGt",	3KCH2I7_%VxB,Ux0}R*x`esJRv8Q5&JykK;x*o6!Fe.cg-V!Dq0r3Vc4BkGk&`QLxmF!eXO5ax61b`kp4[t8a~FEWq{`oy4[!Ee"~>JlB^	]x1X5SWs.]5I!5`s@f4E"-\IWgd,]@pNZIh-]D{.sw/%Om5,p%*a5jBL#S>P7p-7rd&Tc-dNsOU:b+dcw=?Ak\CX<AC?W<NkW3='}[3&V~Rp5yt`jy(vB<U[O#'zN0X7Q`prY::"CjsHTvS-7<G)8=qKk7l=V=Sf.ng2m%"&TjL41dMCx;izROB&}	c+xI*e3^`RfJ7<siV5JMN>OFH4yJ@kjSa{`q-D7_mvkb5gM&MbQ\lGCQ>8mz;Q&
SoAt0[.fxW	K7zUmc*7w{7j'rU`C,MPw5Z8VL^rLk47SI5aQ] HB}cr,[_Z?)!,N^~]}XV#lVq+*u!V&Kf?P]+zc2B@W6`h"<JG3MfJM%H(J6.2*
%R8@(&xJ9-K<,"]TW8Ssh,f0(Y)?DSL#,`x=eMir#6>Slh&}JG2E;QPB*;!%l1:Z|+q=,+d[8|9}1h_IMtRlQKPk<sxy<e<~a"yoQt(uJtosRWwjbq&mXUR=d>}}]&a{WfXX&uxkam]Hfn9T;o,zakV8NEk>NdfjrGR'[b7A?TF1,5~s$|:14Lf]zbR8$sIPV;H(tbN3;2s2YR*Z_0,w[!U<4lXsV{7uGpdpg/DtS!/ 6 2"LJtY%U:O#=eiWGt='60]k0%:47<k&AL['x 1,`+!cXL{;,>{G?#fX@\n0!t)"zsN$KXc6NR8:QtE8xY,} tdrO-$tL6*aLoeySd(]rf\jB:M4??QZh3Vm]+:FSoE[EJhh6YB^2vd9]Ij X j=]SUai'\Y~3-L$1IR9Q=n4QoIo+NYO^<_GXKe2Lb.(GqR#<}g!b?f~B5NJ.F-&eNZ>n&dCB;A,Wto=^" 0h"T|H*s=>>w.?ZrqoX/V D3v'$
R!	71Fu	P?L-14+d	ZKS7<
F!jn27[6c4I07)*d~uXn]<oeP
gi4qXmdH=_u_'T>TBIUaHHA0.@!Fo	+&G(o_eTz/8x)TT|$-."	+`-B-8b`gfXbMVv,I3f>LHjg',UvAH0=lFJb	JWDJ+`b5rFnPRQb{}>gAPe-sB	?Uh~t1v_MSVU.o_Cp|t|C";C027TU\.uGj4E+&Ma]kz>Vv^{+{qf>URJ<^mfQ)_+1>&u[;3z"iJc)DYtbrx@6sCDKb3~o[c qH6[N;2{<pF[dJ*ObMw,(,cCD$JbF0bn=,4r0uU!h2ha}'Mwxl /%Ive;gMW$\}8FJ^YN/w<S(/&->te/S|ToXH3TPS:`V;,^^CyE$ R0oe$KG.TM!s^%s0ck^lZH6E*P3z3!V!~cMKp'!ig?c]st
g),/@RRJh+D[n+SE5x\:i5?#!\EU?<tE`H2C_Ry-vX/,bI.>6:u.'tc9BX 9Ts0 q1&lTZ`%&&G#({]{/d8GBO}0U`VS4G$7I,NVxwGh9GIf]BNm	nC7r0lDNzbtn'Sr_4hM]F)EPj;u"tj}"e&sp95DEM:d1"Zb!pD=F8s*_!s5@8Kom%3-..cB,y?99dW1&.U""|FwG@TD-FXsVg[l<TH0)#H/"d3^r2aXv&o`R3(&5I]6Z	!kq3%js(Yjs$i	"vK
Us#+u[3_{y%)A6s$x[hjb!J%Tr_0rYA>w}K3"EPn7);],4)N?k54~2gC	:|D$Yi}*PS2djuC\K34^h\3HGy6l6MB|N!2D{9tc{RPv.+v`49;+Q
,i_3yIr#=,&=7b2HD<V"J'e"meme1pc`Lf!.Vw!)q'27TmNIDYIy!I".b=+Ip{!JyId3)'/V(|?*2q";jG<un$q*ndkUZo$!c lb]s0 :58`}GC[Uhf_>7g3\;,W8	7bqh1E
:n ,=(GZ|HKEZ3==9U[:9dZT[DIr,ucRw\ ji?R)KMn7z.K~K^O_?`ZpS~>1j63=oaI}(DC;U^y	lu`7ZyDno1.rw,zzSG!PxW6L63>rjL%'|S3:s$zY36]H{dkkRX6;sT|&p0aQu:kp.W?jqcJ/g,O,_w/I>.#03-	
SZZlEp[y6[AlY}&a*)\Zx_8 -&&vi^oHB+>?qIjWSkI0EjKj>
,#U?`6C>7e KTPd.<9r;3zVHzPaxH uh&21[vG3M(b-fR1JEOVy!(K=	z!;YB.sxb~M6+0,CJ;PJQ?prd+X$tC^+^7T1]Uyst#3WTW(pbxN:U1Z*Vulsl_
"<hk.{c]!'KT8yVM9u\Yhn3J#94/q2!T2iA7:JvM3
R'$+(72E,3KHb0h"vW@3n_0BW+{O@UGX\f~w#;V9i)t\lfJ* (&,sGDeo`}WQ+6L<2<om\^t!Suyb:!@iwc9I3 mwa>1pzk	p
C]RQ(XI&1iL4]p
Ut@@7hwgsR7-t7|_:}5>RTwEOxXxkIAJqcB6tv:=e1n9>F3^c_YA@H`M-EeUgNG=uJ%&p#;a6IJ|l' SW/E,`i%%Ph%`@PkCh5NueSR Rk)UH1/Q481jl6q=`CJy	Vaty<O,<z%)kSg/lR|wS;#m_x"'V!=.c434?`%4m!<d1C@4Q6tRTYSE+Z)~A>J2SNI>ClHv:dkY[6D6L{!Cj4Xf$Bn>BH9-'8-EJQG@FPy<k_Dk39KFzx!uBlvm@ b4&*<}5C!m/85
Tt#RV>kCE
ESMb
L^<W2vV<48:3|~I^9T	j$JDjMlO+	e#q./GF;C	U0t2;%t"O!RlF(H8V]XH1ZesDb#t`Mr/7.vaPw=+H
`kIRRsk3)"_M6WmN4!/|LU];[~PJ9S0ko:eZO4D!\>aAN+X%ffI3AsQ+!1n`	:qyk_={1ZHiD?,5f38's2L7w")w&WO5^:]~-p'wfIUnk:7PZW`chgLy(z`_^+G)
#;3F|Er%y@KGW5s)4up0ZXtb)fnea@*@n'X(#0Q.)|^Q6N[(C!tD'o-5Q[ '7y|^<%:Vy0>+|":1,V?Iz[8+`]6e%[Z:`R|*sn0	{GW2?wnRBN2vn$
'&k@b$16Vr~r;0oRAxifJUrw7`"Y37CnoBKt;]cG><ESz	U	XVW`ai3`JSwC,4r\YC.nZOky4.pwYnYDnzj$8LYdZD;;UJ&aCWooP_hv3Nbt:\mFq`}WSta{tk	1,sJ][JPJO1zAtQGOoGYYC:LrZJOV$E==^<ux=41E+*)n+_k,zIxHsfUNTz}7y{z
-Jh_JgcI{%_[7e
#	V8^]R(.UCd;m=6x={dCB:9d}ZpE70[l2]
Ez\0G[3Vjy{@CC K0@!SOQ5Bg-tX{%<k6
O*fb
!TD	?:8ob(t)!m`.2wmh>LJe?Q#BKy-v=~ILsv-*^}- ]nvPZ!}@!j$_4+90v}[-Y!i6ZmPa`BGbOa`,1?Y9-IE;iT<FtMx(n'ni;3lLjIeuHA&9,Egz4ibTg3APjd#eUQVHJ2R9.j#L&0&q+,UlTb/7A7`<G.BsV+b5Dj=R(\={.gQuDA7$})?U+q/3^vlG^w3?wpOT3e6L0c2L4>O~jC ,e]`}4n3,B<GOw2gjFZu.ooGVy\|u}D ^PFp'V65NP67R+	"#@I#&q$\JY?poB<}O	A:f}^
9_\	;N0/	bi{aMcC*d1bd|ZOT747{-OIo[=O2n&R|j6NdjS}Uw"X9L0+b/w<Ue!1ScLItiN*,6R6(p@w^*Qd`/`Z{W,gw\ 0fo7Y6_3sN2qaphu^{*6u<W& &G@&H/D$<P0fVBvL\"JCI1.m.:vo!BPCX0^7&Z
4GJk]&R[!X>Y!mU;6gm1)eFqD=fZ	$]t2DGhT0fGb~)eD;4& 	kTxGjQ&\*m:5SH;%cf^!.:"msOcNU<'hM#\-HxxWa?0+$u)G ectEac}M=f-@Sn"/x,-M!;t*sDfS4b~`(i)&@}BK6,;_2nJ^yCIc6\CD3$^b\mCQJp_M6[8ioo$a<	T!pxFJZWHI]OPbX"VP,hQ/|TR9pG6m\
FvNjZ"6H>QDw@@%(NYP2m2<OhL\&`dwJ9tbB6WxD3%F$<FGHvIP'6+ELS	7iAPg)R}6eZh]UM<1&	1q83-B0zAV`KW@+:-/y+!ETgRcaNroM(FI#5G3hlLlku[D>d`r"b\e\2~iiV	?[Mif`L-VyxGOrR'*HKa5q6;}%lPr2i Lw,b)PVBQS|{L`I^PT3 3k2RmK(~:'mih_1G##Q>
<xKBxX^DQ&
*M1[+n%B?N}(uOq.kok.\y?@g8dRJ{R*;DS11_%k-#Q1t|iH"{Hjg>*LjcFUiK	~b6&/ek5sRCXuov;A*[:XT*tuJ{&lT2JPSMI	-d	oK<?<K^T*PA'BR7
bIw3QF!`rF|fiy^(b	7=*X,~;T+QRS~_Y/,TadY_>\jU7DY{FtKbL(\8`A~*}m,`%%'TlWOOG_*EF)6{a||TwXt oB?+KsL*f Y0&,f<"?\rfH}:oRu0hC+]!oETdLk_}JXq	#4f$upUUaW<^c[VzJnU),]1<"&~'6r0d#G3?Qu9l&<UGtivJ]aREvpk\Si/J1TaH{Wy?vF]nB[7`kP2{AVG@KQ.,hvF;9)!h}gb[IRC\>lms7T\L46+YbG|F!jIonRwtYGVFp.op`%|jDdC45H%iLLjVt\P5umU638yUy.</FUBvgByEa>B1B-a8{9`LB7t"{{9+qdn{#\_,O&pBow=k$F{;(*#5?P(TsH{DFQ8^:/Aw6S+07bRM1zectLT=o<WFq^<ec$iu'j3x~$AK>xt]`'e,gX8$bykknv]3)lfdlS"}NR.A{&@mJ!7dibGlhygU"8SXhF)</5,;]&!AsUX u5nd1G!nn:%'qp*1|wCJyET\N:H1pQlW~*'%9!{(]9
kbG_n2U%(*Q;q-+nt}u,6(bFOI1j7r)$@0AH:%-3~!mB.U!{R3kAd5xP)$mA@RsVJC?'LJL5n(>qT- uc}Jv\uP?'4=$f;hLs{7`2 
&N~|zl>5Oh=c"bOSi=uK$uwzEQ=QVZ")
yM80i'Pmu*<\-W2B{z7t	5}hF'/FcOkL2NH`kyqN$*2=3@/>jn//CCIq)6~`d`oc7:	D"5[|$!LjE-s,`,;VVNJP&kB4xqQ,?,au=<7ME1
$xEc<}JLm	jp
[3E6}kFZ s_B9D]FG\	wy |4zzJ|$!0*-jL?LF~5qEsf1 fXn)OqQSV~@poO$"afG]!2" IjFkc1m3Wl`Tr{#SM/u^yD?l}#g:uX:[p1/%o7g	YE\HQ#w){0RU^bCj#NM=]/Ff._VHah|9M3y*G\=uQ(?f$/AU^BDxd3Q^:I_(=Zt(iV.b0BRh dW Nj)"eSc= 'Td|0LXq91Iy]Zi!L90*-k>C@8mJy@Py7*b^e#fHA.buaakzl)qr#	>LS=Fx+`5N)S<h-AjOjT5lGEgY+14^IF@=thBz]c,w}en?_O\E+Meh]k@MmrJ}0xP=e-l,`*nJyPXGO\WzbKJ`9wB`*b~AP	Q;-6w+0|QeWi3L:-R6!ks`}||xSD,xFwu5+C(/39{=u:VAvMjY=O<$Zl$y+lT
ww7=:E;'Rg
<{3R2v3l3T]8u;r^kj^Nt9=BplN3@Byil8p24@3 zQOB^WgpOF{Gb&eFz/#T$=@eNlw)){]E^rX$*nUA,$;l2!(aM rxW:'aEa;fi:L|1(HH[I[xv	gH5T;/Rsv\>?R	m^<\&Jvs:eyS]GP[7L81aFlyz|.c(\Y7g\n~6O%|:Y6B_4;7ZU3&`-\hS)EBW}ax^sOw;>Y2fVa[WdAkszlk6d4#fi3TGZbG4`~@QG*sUSs,\Yp0#&2PTfxUA(Q(l/Iz#~Gd\C=s=8<toj/!HtaRB9'2g#:@)GX,+k|U2^vp>5'1krnltFNK,RKa(|+A(GuD&-\ROob~xH9zxb@UG!^u<6EP*n}5T'GM!Ts7f%R$MF|q/$&JhL~UT[FD9Y1Yj?wM+.aF6l%i`IimI%l$H_#FLY-# &w^'RPw'M2GjLa;c	:Ojmx!D%Go&{7PD=swvbb<f\}^I1^D%iN;Q+5Rx8RD\LG0yY<.M[XfV
l$]MeA!2G8STVph=ZYoKlgXHs0jer'kk@Df\=/0Gu_C?qe$!o4t	"9VjR4B)]#.{TXH.Ffh)@Bw/QQi[jg7R[<F94(;"Rusu4!L(gx7fYC/!HXkU'sQq~,&'`1d-D%/`)-0&_K)lI|Mc;ytw	G?oQiI(<S=\fe0=5IDd/BU|+wH67.~%wC&Iu:Pgm7{J+p'%0+9VD=*?SPN&HCE/PJ
3?^1g$64EucR{%'mQW1OU7	K
	Lj*dtOoP.W5T7a%~zu\,Vplp:2gbD#j`^x	3|)GN*.ESkB-12CCoz\M!jNm:UNU[}~#[6v8rnolMWge4\OY41GW_6g%G4Y2PU]u&1~k}1Ijp(y2/}%@xt8#b|Y /c{yA2)8](sN;1t@lGXq?Qa\;JGY_`vt"-le{Q<FX:XW>+;b<P1a	4ce3wIw,y}vXhW5kvtgu2'ESI(GjT,(oXOfZ
+)`}0e`q](w=XD,RQ*o!T=jzX,m76P3w8{#XE=r!Nq
KL.Qz"uc%lx~ziGBD[(Hrd>MYUmlxV]N4"p3iXc1d`&.2@f1n"pO>FIFltt)QO{d{?jB#ax(GoJ`(1x1JHy4Lm<W.XR|)7;eIG7Fwt3VTQk1||G<kj8B_Cwb_dpA?'K~@FvhFnKU}PVpPh=Q1okfWUZ@Fdy	x`H)H>>sJ!Nz!~NL?]Q"B_d_0_J~):[N	@,UiDO&]\2'JW9X<\`9%kt1cJ?L@Im	JJtuk<K(27z|Sno$DBCuw
?61qW$[I,HI<[A1PQpXeY:4|d.5[HJ@<X^2VFe5qE?hHe4	5
NaE 
!a8k}q_T]I5HnB	WA^PE.CFg@G#u2e3y1F,Q&kFo=XzMORf]b/_2.O-phEMMoc&4bC.TH3^Zp{i6.jo4qdQJIfH"zGpp:KSf%{-3Q@RE$F~O-A'l=eCX=/	)F?cs>U/}Fr8LJY3_,6#BMri.mV1|=gT""BFRIXpng9{PZ$0}m;A:B$UQ!vccpif--Ths.}Zrk:7=J`.y6mwmmSNv~Si	#z+&bhjkQ8e/_qND8O'jM|;2i64">R|73My&Hwu"=5#
'rZ!NCSlwi?g%0 $bki	G	>s-DcK<Tz#vBz%t%?ijD&sX.HNX}WtYTcqJ'js!pE"	~5#Jyh8Chh9Tuvq3=`+e70+k[;U>QqpL[B.}[yIKBwRPu_fvnl(#	280:@U#F`+*,{<nB=n^R[?aEZX#rSA=8TWLdA6IWXb/uSJe:l\OK^C Fxga(m=.hb|Q:Q~	L6FO>he|,8TUh|	gjZ<$uSVgdb{7&<d37WR3;C$$
1)?|evG~>7JaIbTrO"n|%#FTyh+3U[I;:Vh8Sp<d31p'67)H8S~.P(
b9YMsj:yXx>+hpj"OE8iV&3Ou8rbPN.UPsNb[j58b6I`w@5ZQO:S1r~t"=6tOD''m:I!Y^p)a`FfZ81&[\%z 2d kE%"l54/I0lu\R+*zmR.pMgi_?RE+  NY"TL_f$E~lR*glH hT&Y6k[7S8~3r*|N^cx%FRay_-zUqHFJhC_H4w Z{x\sxsF$RcM? bKy9RqA]*j+`~
cJtz("J)}(qnAsS+ET>]	L.[
?f@w
Fs%c[naf=	a fAwV^T)K/Os[JF|z09Oe]/
L@e#afz4A[Cgd[XBeTF$:|WfXC0}"<o\#z/i>Oa3
]7%kHK}[ccg.9n7U20cf3.3-
-X3MGeS^,[X3aT1e?C	1`xt4z)%73-CG0@8( d4LonfStcD&pSm`(0y4/J.q&R;fYBJ$@*`+JLZ$#Q| &B[3VZSSkLGZw$<FAu)>`{&y
*SjVNuMr/4
-!W*	EFD,++x|p:C")J8Wx ciE^t-=bc.BXxZ&yZ^@L_n:[cE1ivoE2RH`fI>.zZWEO`;=uC<Z'_Vm'p%%;;M)ns`c8h7+QgnM?E@cf6K)[5o4Lg4L]>UmCC(DK3B7)ws\FIjCC/687q>tF&(HrpEUQ:F4^AV7	U!'
RzeN&XG-hB$4nsi(+'isaq!IvazRIYB`C Pi3	'E"*zERY1Rmt9	mn<AD

W"O-~ nHA&`R'|.$9t1m666-cQ>?^$I9G	ui&zJ'	OY2QX/h	xh8jEUF9;V.,us+V<i@`	g.~ Vpsl/bU>e|2fpB4jr%><^6iZuG;/sFfQTZ4gfi_	WB|zW"#-'^?"9c&7Wyq[0b|nvsz%5ju3BdJvH=-aY*WZgyfI1xT&_gWO4L7V8&B;uip=v8i*W%@Eb674-cQ<=`3]^kNF-sI]ohJR
<6b`<\b2-IZt$y_kCD.JF|}}8hOoBby&04}'t)6r6n-yJbU
Gw{7Q3aUq~:w2Lo61 z<dD/,%s-\.U()G]1WPfX8:pt/_i2|D4x~w1Isy}5EbbY9jSB&+B$~aL/<~0GHFc6!@"*<|dIgg{h2rHe@X`#D
;]<?_iim#AO*c`h`*D;HtJBiEI_7aMKBgHu9	Hl\Zg,]x=%AWCgniOWrB9rC
Ho'$2I0B)R\:qF<$O$7zX2,1hUQmB.<Fz?WIf5d"t&GmKZ/d7;R*{9,lC>9AZ=o\;U&7fS(+J2y<%,~sj2[>w
AUfoeZNaLI9@N.CQ}N7I)>m+q=*9.J>f|aAa\bIj[S<Hlj\$lW$5!Q*+DH`vl=c'zq1T17}7#x
CZBGQt!,+0qH}W`|lxrUDgP7*XS^^[zd-08i3~<*x#to@o=*hiiKLj^?!3kEGQUa-S``sef4s',@*v$	dp1)p/}nD6@Xg2D"|O0sqz(2#28\YY9^^2C$!vr}38 =zH_akNFU:xANb"``Z,glT4yWOBn#rSZKop`}|,;]x`T=Q1mH.Zv-6"b_inY#Z^Z((P2+2UOFZ,S?")g#^~	g.MH`A^&0`woG{{`+nkp}DIz`R_<#N:Q_$
-<B5x0?(lCn-{3E#C85uE6/:a	hd$M%vM%O71|l:)P'[gi3%*n2R(Qoah@z.7#jP]	0R
utepjwhV4|
CM'AsDJ'7>zBm-u%pdIC^b
UtvBMHm`ZTzo?xK1`SCv`(-#LC+(iNNP w4(0\];;ZXq*0nB<lFQh:h5f&S5$;QM}hM*76~":t'kXU1$$[F~RC:%c3~]0W8S\fa*BBbki%8rTbA{#
Fm#v]lpXNn&rbFzUxD.	JgZCaF=<HvOg~_ngEy|ikA
Iq{`98;R7qmbG9y)DhUd-Eu*0vNc4N19s96swF/2=i9:th45]C(,9z{+LNlQ+T|(kDGQ}p)X`cZ!E1pE5P 	3Ou~(+IW<2	zJx,
#1[0Ew'9^-`c',6^Pw4tV_1+N{9nt|(;96W'rS?=DqTt}drmR@X@Kwm=3"=|Lqvb{	8{NDVsbe0Xp'Yrv0='-?k,nSob>[g?T "_#8E%`yZOdC3n]82,tjs[0MU( 1K_RU!\?~F"WAfX(\)7E3.Ww1m1CA%MI1Y4D+%R	.r<@/N^9#C["lgr qw.>x+BTLUC$2qf<WNn*jUS7sz1*lKjDipa1=(?-wCV`&S*;TQz]/1Pgb!H!O@QYTpPe&B1?kX\w<,\HZP9SkFV	spjowOPx^	!Mq6Zl
O:<Qa'oQHaw.3NyTL/*Ax{NY|6jr4)>Qy gV[5':d+1JdY-];iT5u!c+zt2g3nG z{	ONLwD,3}!@s(eDb\%i)&8@2*)]NiMd>8?xrCJ*Iq`U1l7URz+JC1LyBEgATZgW7FS,Xy6WGt,z8"}(1Wj8<[s$AQMq0RNu/p&e7=[?[wITgx"F$V$\
M]`%)vK|?*<0}QN0d{maMrA,b	/XDMSXISj/
t{Q:=:.&2A(h	}r*.R:Y6zCYr?WK[~/)X	&V_zEg?&s\Y{ RY_z|==;b\+f&3#J[\7"4X	Na+["+}nM=!1rN2={	=#Drc@B/_T}%AOO]K=5!/a$ph+HVDOy}q([2&):43rLw$nT:,XTMp{GUJpZQ_jB|PL/>c<k"hE4%+cn:tu	_|KeL-(u6 }7yl3eHO$00n&/(xqv@$SDl0i$4jh6_EsACL}/)z&)h9}A+H|otPH&!T`bD*=F\Y6o}?D\<x4kS_5.f'j}2+?ZrE/_#`p48oDZ){V`+&k}E(lS*,lLP?Mxv.Qf|zN|`I)&H L(>	vm3uehCHSB`7. nr5WVU50nFo$ksE^44nhS4Y2fDhG?	L+|< D jZ=L,6]{
,+u)W#ZS^-i{[Rf6496[PI'
0Cf-eYV;Q*|yA*@Dz&RvUxT!gW`L_F."KxC[U_y/Lz*MK'HmC@6W!3^g^wJHkT$d,3f~%n"F=Mf9X*Q^vi	o<@=#|YyG+=ayY<F@ cpgB5;@esgC{MG#xlc.
2KBLsr\-! @P&S."R[eW9CvSCZO6!-5Y12c(m4ppEvnST*)N]~/>+[sSZ<7?JvS[RLN+)up(=>ocVY/7	bs`GF2j5^G5|dw6T,7$r*i:5`l199/Sn3cq:8O"(,qu^2jlq!-8s#&0Cmn#7IXe;5Ij5TA+?D7OYt^"@HASoI+c$7U8dK^}KfW0tY=T{J.Tg)"=&$k&`
=hv~da8h[~
dSiH.Rn`i`#1{T"CTFs	?s!!-YjEZ<`h+d,Di3Ntfk	4C7l%f>
1s]s1#0|w#GaCs*WR2;eVQ(~gk,HA46@%dSrt@2>w
/p4V,@/'"_r+n`'_@@?i#VBix(uV_T`&$YB	x}z%-m!,yShrO6k:c4%BkL5QM6Vz5\S+tgj"E6{U">_8^j6Dm%;=I,XR <y"IJCf`-E)j902?1]lJan7tpt'`Dw5%Ce/|aNO_e _Z<F]j9[_>q:e>y~zPUzj6KMq"_Vlmy:'nE(XyTSj@/4`f!6xF9H;S$'`)z+KezRe@X)_Se
!cDo_	Pj*AoAc-o({Xc9j|;	uyH![i^Xv/5\lRcz*o.?tJ9	=odAhA-xZx8H]UUNI]!@?
-f=aj+_XUU)!$IW^#wR0AL\JrLtUx6eoj
1h@y['{qMor|wWlHKwe?xDR*YaNL==Oy{GWGC;]!$v<b?&+9PEDQF9]~-kGVR*3!J';fnGz2
67SBL*=vS/z{9H5P4"@`8@N8j-[7'=F!njPi|qb`3$DuflxMV\F5vAO5O8i-]h>'*O_C&Y'MG{Qm1|y%iqw6$m
-qnoi)B Znh:MafKnjEtZzPOMb|a&IhH/;xe	~_	_}z(632S45:z9<!&$iv%DK&k?$V2`QW^s1`it4rB+P=}VTf4ai,vb:kQE88,{!49$dNH	$]uSbb.a'eUDAE}:sc^Qo@Y0#ru @[	@A8"]Ai?9#j> q1<PvTJrLG&];i0-0_E<pspJNW==O=uHR2cyMgooscb	2hWap`jI1?-a]3?Y.lP}+jeC1O^49gXdPb3[]0'&'Z\)"hG5yB:&7c%%DIh;y4B4d1[s$c4ppXas3Gd|Yu.3i
'C$oBjhb>`B`q6RB[J;"|l&WEY4S-t~]|nF,vlWF=:$(y4{M7*M=D?Ga">L#U"Z8YiWqdHhu_6L;;{!^9v/EA;s1{d;y$	Ip^eT8I!+a`z[?'#L/Gz{aRRbqV(oCvpefb#y"VYW|hSd>'a,8Ni|30,jLCy%N=pp:v,K=C)6
Y,3m)LX@9MH/ GYL>{L'@?4]^ UX&;DGihdcN&AP^=M=j fF3V^$`Mqu.9g;5-q65.7\yS8Wt/oa3}o6sB60F`NKbR<B:cR/O3Y]lkRF0aLI3F}4^4M/>PGWEhI7S/-(q`SXF(WJ5HKEk2Lqh\>$=l;_CSoVC304Uoa;4IG|#_A~?4YsJy TK.{X=f*Y	T_A+BE!JBs#vG[ajY8/.Txc2&
FmRK-Wxfw
;jf,X47
`pKak^<Ec`4l")G~]@9y*Xjen,ZOygPiQaM7Rwb3,22`W")<vj~!e1!1i}sP:rWN4AynaQ4GN\TARa |E*uM]|Z-DV	&{,_CJYtDS0fuc\'Di]+*3+iYFr+P%_RP5iJJAn$9) yCzj88#d{cxQ(6!eDY!*%MfgXBz,hd>yU=Bu!2@+{)1An<TzE0oKDQ 
8doB4.v`{eE"NE5L/q#mrPx0V7@8Q(_]#xCgjLpD<"TJIY0a45w@}	./LWGyzp0.YCC@:0=F	PqV3@WO>vi8IW/.0j1-@K_VLM9US^.@6/DunP3f6E{KT}u-Nx%nO1)N*10=Q&VCxv}2q^p?sQ'O7p+t=g:,1o}1wVn.fw?QQMD=0RR9cW|A}/%nZ]+N'OR+1qf_0,XmW>uCui`S[bi$u}/#'77=mYUW2anjij2P`GO9>'ph>XCVj6E=Th)&ix}jR?Bs6S#Z2HJu}vn]uTRT#%meFH(xYOAY}v3jRXf>SQ)wJ%>h	Pft@x`C.6gdF(O4<lr)EwzOBs=JVn#g'dTh4U!G.?,@hj=xUYNA{Eu,*E6^4M^!B@329A	}]"^A)#D>5|tTPrbn58^[a[3Q1WaOZ_j/Lg9)fsJWsAOmqn-x1.vUGH;]+?F}Fgr|<Qu5th#%	e?mW @J"D
Z\H||]>/m:L_{ij9y&^OU)G;U+
7r3&ko<VR	Q5U\:/y*1qD5aTs3tT= )_UYY)}&J-2c'C"[en7JMPE.v!kDdM!O#0@dth+t'x<'}{kM>k(<{Jee(Bk7Tsj>$m&k",Q@r}i5+OF3m$97Y<U@xU&/hAZWn0_uP'2m-;t"Cy@,gr6z4S
$NLg#ISU,]8ve[G:".anWLFC`U6 qh{@86E`0.'`&^HHD
hGfJ&pGQ	`MLJ3LnT,0kM4cBV1|/q>J]i:]H|TQEON(@>B$c+c<!a0PIVn/_eTiNeGHuejKaLGc(\w*5m.rfKc})8w&k^\"Fy`!!WEyA A57Ef2TPlxqM/oJ}vhNV#1F+9It<8C,j@Jm[sD
Mc/lv8%=gtbM{PDX66@e2^0_k`yP:1P[/|?"+[Ev#0DE
sABt]duMY:(bw4Yp'JO2=53]Md%{r<Fp	_QoYIE*X}{$N.|Y}TB*mjFM}BJnHl&jA#2ueZ2{PVZ?:z:2gM4K'\VWJ%/q./P,YYO2|CxgX@FQ	S{IZG$tD]qf!gE%!'"'#AL4f(^:	TE7``"zlHb\9[mqeMJopZ+B&ECB\$$4liY[X-o3z#Gdm/?e@_my[xAA"d,g_}Mh:PD*2w88*4~b5iD/#D`|>	VNV91jzd%nmN&{1(/{Sc=HcP\+7 @A%l	<J[2^b7<XnSo)&uP~_>9=`wt7NSI!NOq}H#Yo
VI#wp,MW<0%+go-	u,Jaw--v"(Qo2MKM8jtlE#XbI;[~PRkA*V_!)&_4JOK?v6_|-IQ%Cm;RrKJyWt])kvnNGlC'fv1!rCGK 7/,LMu6&Hq!	|9@V:y-}^(*T)poNY8X%PkHWnu%kRTq2>FQ.Ym)."Qu*V:znF=piNg-M>2T2s0~,ja~zkZ=%6o,4P<bqODo[^+(p%Or#8*r}70C_+]x*<^jzD*&zhUC\N	<K))HS>QZ}!li`pI?YlW;sj%kJJk#f}/kv:umg!Ne=h,}'
;CW+{`t$-.`
bMI-o>QAu{&$84~5/-S*LjnQ4B}PQO,_9H)3DdWU|q*J
(}|q|\,%V]
z'd*X`*on A<)w@9e"YbYW{VQ;RtWsx'IV&mLH)cs~JwZ2,ZO=%p'%I#1>I|g*]Ja.TP&hB5cR?2AE~XkLWjC8M3_	Be@z3.>?B}_/]IUJoQ26YAB;]EIBqxDu,t-V+Ea_c45j	gF!OS)]=^AX!,Y.C	bu^"dNN?UpsmQ=%?GZ3Ad`C],6hf,"DcBA)5{wu<`RcMDDy@mD=`NiG0x-Q_j1BhDya:>O[MOVZxz3`vb"%8[q#=(wVn4_BUZNO_wsWa[$H1|.c~hk,AQV]7W~R}fqCd6B]<*(L-nQ:"jbR*J^:C[)!9<zTpz4}I`G*(4	QlVDtpII`}HfQK8~yU2@:v.0W\x.7yY,-s,XA3gNHNBqj*dcUFwThRE6=:)Xqfx["Xc2%t1edc+i84So}q`D{@)mP$iY*"3^zJd ]YD2=H,@y)D:DW8|B'E@]V,5;'5UH
X;O{5W*TtZte?kPATbE~M;
~LB),sbN'ZGF-i$I@QY\c0}n*A7Ss)1LXmn(BVPZ25?/z%VSF'rgax3yLi^p=bMkP6BJ:Y==a*pX@F`Jv\?IX
9@bI0Q5Vc'>/[<JE_wsIO+KO+T]}V)KjC3N~,IX2+"bY3//%Hz*}}Nz$K&RlS_2>( _5zE2[

?v/<ph+XI2$%nn&q>H0JRN_>VEiS>w'|#FsDV/QM)Ql;yO#FgwT>Te9Y}"B{YX-$`;Be0VrL%j2{6dA8_zOAh` %YL9Xdf-'lsRLF;&*:??}]%blpXT;9i3i(=['iwS1s_@G+`}z$4%rTYbzZW/JZ-Y'2[\m\M>;m#*wq{lM3>%Ck'Y:/
qQn.A(Ex<6Nb	"[3afD$;^n~eCA	Mm|%cYwdj+= WeVdbuo^Y-w)"61@uj[V^lg}Q[ZUuE?}@*0pt$DFrT`~O?7;lIGsRR}ak"=cq4AD:;Ij}"24#=)\>azwa1,DN_^?b6T4w}LDg,uxM-6{	>sRWef)1^0)W98bw`>nu\<H+sx/6df59{A|1(l2lLSqc2#pUDxWA|YJpg3&i,sIV}y='+EktooaXw^)4lz*e^A4j,HdU0^RepulCC'RD$6j. EDy<4d+2<K7[#)+0L9"8e.9N/9hKdG%M_f;=5bt~V.n(}lJx7?BlkXy,Q:Q1G<yiy8GqxM_2J-z!N+>PG{CW8fA7E"I:Q0/3#/)G)j#1b>8b^(oM#YEYBA+hQ0uxzdL
3<)4T:lLd^%(VivglS&
eV8AK:-ImCk#G.
v7DbG9{Gm6Y9S7>H!5)Q8367=G!xHk!*U):$eL-!7~Qf:NsG,]m!-\h3{O,`xd&mSw.egU5..(+;?X?4N&>[6u@3#j8U%	q<-8RV8pT^KkV)sds=?{EaEJ7P(<+@La1\c)eFMgQO.4tL.vc=P3sN#0Y;wr!BCTCcfpq}I9,*&w:'<<AOUTR=N-2r+#v	>{,M2Qayrs2`2Z65N]TbhNGtUxT
}&<0C5j8OYIuNfBu~mZ4G4F^6a" Uy`wV[OZsq&,iTH%;_wt`_JD\L'+\F+G\4h:Y_'B:^,17:_/nhH$s&	{qa_.\9]#TU#\ZN0#Ov6vS*q Q)sad"9Eis3vCAQt2B?6f9te{)`=ve'>%6(z|pl
<F8C$6[m7Dx+KabLn2/cMj9c"
0[(#pEl~&|#P}1&$aFQJ?jIfs)C00I{-dZ|kqx0>4t~'e#*mW"hm*Aj?JE
5A)p9GmlTvPy>WfCTK
cgH#LR^!48Ir3Yf,zfOMMdDRb2
pb	O:ib3!m<Y.&#PE2_B#I>
w.vnEPIK=]=Lj7nSG>;]M,0 SdJ**Lmm $d*!\JM5bvN6!!<	[(m9YiV_dj],.d9Tv7Dq??FX![*Rr#/pCEcB#g>}[]MDfcHx)N~`0/-SNBG;[y$09Ue71I*7hGKMDJS!GPIyn65\?ILofEyQgN;jL?=/H62?n4|<Q-p[EkVmp][z
#%O%C/TE/Fc(X0e*bR]gk2%r$NWMrVD:M=Tpgu<z4!;r(4F64_!~mO1ibbET1~_Zs%rc#r.bKF&b(27K,G=Rte@b@Fs'2; >Y.>6OT8,P]S	Bt0J+Bf(]&waO8|lmR	fH4M},\v({x	z3~6);#R1]F~4eK?`pj,|"Q49JNi-.wX':lk!0$?SQ(9d^r#Vmi J	<;uk=6#>@:z4{GC$[;Zu>:lDk"TIWG}Eoz4R'Y]d%kQ)ENU-!q$_$DWY'gpB;@/h	p^9,AB)LFzv|VlQ[x+8y
PE.(rT-q)?g%AvVA D)V^ewKjq<C~&0eU(Ps~F&T<[/9DyAZ!@mD3-gsr4X'3;YORrg~$$	GbM/j_he?QSo4<;<U>;Q{x]M.o6|+wjk9*XoMnuOCK![>xBV)w"E\^* -Evk#:)S1_:<VyHe7[>zdv}_HHFgl'RCA2,#6L`B{C!gK5O'=}HV@<F54|w2tVJP'tZf}s2_|n8h=2*Oo_JO-x4^gDUAb+/#W&nZ3"_'w_L0bI@"
U`d${qqbK0(8Y/fnUEY~X[Rj2{"c$+_]?b>[2NCRDy8,"P	m|W@J5u (ts2*pr#DE]5EC/rg\tS#*aS!}C<_>CV_%lCZy|Uqz%@g@hcj[!`weEFudM8it,a'L}K'A#NK0ON.s9u66L5lR`E,lUV>qaXIvz
e:#az{u :Vl)[VlA)M_S,h`;xstz,lX"%EG{<t!XI[xrJVRXyV8/zx7dd`#	
u}#k_(67VMy
w"[1A!<9WMdD/1/kIyhr()jK}97>}G/bTp>"q"c#Tyn#p9wf/*OGT/"UqA'vRTF-(NwC>{3l]g|?-rIQv7yB#ZGhy49d-{d|7Hk n	s*(QFY&k+JKmB;lmtv7i].e2^u:9oQ0}&2Bt{@h(% 'mV9PPNjov,Jj-T@&CGVCcqC6y3pz:*(~
oof;j^CTMbA)P),?SpXZ@Tt*Y"QKgORqF0#Y:2:F7ZIA @tMP1'~'jDN3G9 c#X
U,=ncN9^_#m/qryss:,ife6'py5M"P?R}<=*;Hi2j!W4^vxe\<rWie/5Nf:V^'TVZ&;-I4za(
=}s/=UV;)k##b.7+}*_>Y\\D#Q/vpS[1m(Dif>rza\oUAKug>I41i1=oZX<pq[+,\#!v|{bk9[;
-PI\.:k7Z-3codnnSyA
ti'i=8W*Tv,}s! <3qda,*t:EP7W3z."4;wG6epbg#Z_@@SXz@oa*9a0_[enG#h=d)[_REDzK4]{f?EFv!B9+?E;p#9[xJUi+y,9.;xX_C7Kn3^ekB5lO?%"TBxy/EBm,3\B,ddh6lxwdy['Faj)]eRml[*L+|W"<dX}OMje^%~"$Q/55Tp*;Q(-%k0#
Er(\3ABV5
Ep$Z	3hqQi0KuD_'Lm+)C'+K[K@5[\95LR@WawHMpl!1xzepUlw1M	rnpCF}snF+!};;p(z35r0X*|h#W7Hu]L9Ba0Lp5>[zNYR#+Dd"<8gJ
PE![S_bv{.t`be?C1ED!;?%d[[~:Ac"8SM!jvFRu;BH&*a=Hs;ANUJ
k&.WBIW[Bgr6T#[l?dA"jx)IZ$+"5C"1)lQNlq.tH=S*jyN0C> J{uM#XX.*GDbEY60]_>r
$T2<w"'OKX44eYt&*TcrZ,W8Wu0\;3E~g>we|:];`DY.!!2-FI',vQ0|)o( 3+ww-kz*5lG;^P|Q>JRJG_02]8=VYU{ .F/Ys,\9oB=F_W5#k9
sLF]kaYAGR&!|XReu]xR4b/:
Ys:BH	h.PX#r@`Eh[iNkDfEEPH6nG,_ng5CBNhi#l|(A%i
g(7ocB=9Xt(t,#%$M1bH'/P>"^y/*DM#BuieEc6{o!z =+iZ>}auC@I2 (5DbTp|`M1!eIb[n@94DDFup %%@~x-hhID?n/^%Gk>Fv*.&*&R9fLS}nBh#[R7W:q3vxo,/}Vn)F_5Sjy0`lIJSN8mZI&Ga;r}.;Pju 3L2X56++R}%X.r(F%eXGoafA`0>+9C&B/;gR/JbESU^zrIBq%Y~WtQ\GfE'"u,|J=I*uU:AK{yEso3ESV^k\F@I>_?!R_8:`P$u#m?@@W}Minrz5op4_v|P(qx-NJUtYbDg-^;@^9^i/hyqt4^Ic8r0wzo
HLyaI_;Az,e1l}aVCBX,[E{BVGE	%,iZ%$;<.7[HZ&]\]*}tQL-*#<JoCDQqQ|SRC|0o&{]:X}4&MVQJ1yCzZpVXjI
GCP<|m0Xv$UtbEx<]KoVg<a!1&rc_kfD<wTZ<+9nP`f{<=#[ o0=+g#iY41 c,k_CD([YEPL!n]6*,t,;A.&qEi)?I&!LL	C3eR_RXN^"3Yuf(.2cmMC7}_b4ihhw*]7dXkzj>oA:ev~r}AA_6i-<0IZ+L
7w>	[U:mx@:Ii`NW=b%sgy<wp?:$Ym'z8yt6{_~|)s3qRdH<BHy&u<>MmR9s59;pwvQBF$[Re/Zc|oOC,	dQ?l.E/=?s	BF@sW#jQ8&*3p9 j8h/_w{csm*T3,ai1@P-
m0f>GU(]_dfwEA[D23o?;SN=O61K@_gF&GVq(}%Vsc0HH)JgHdexFdGqZtU
ON!2?l1%!*N)QTX*d1ds?4c9@Ma+YP7q"q@pl&l_smEjc	JIX29(k69lnxQKyqlRvf9Xqi
dP)%cz2aC*9<TD?d8mZFM?]yUfe(}S'MYKCW1"%@;={cjaLVms4~Z^SQcYNqG~J$N\Cvz)Bu	<as?b!y4~Qcp-dZ6[ZaxWRqH`>=x7(G%31?uvafgP-3,V0Er_2*^^czMV8RbmNh6R#&k&-xnx5
>	Hm?qL]h#*kw]tu)gfRd"	1P^uGk2`V2o-x?5Lfcpzp4fbfFC+W'qQ5[,$>!P&#nh8 kd(!EfFP{-D0$L?"+W Saj+u.^>|,MTOO3:ggQxLK-BDa70qUekba/
*m)W	 aj}93dA^49tZnQ!e*KEU#<)L#1AF^9P8J~S]_X^7OZF:bi;%j{s8v gGT%JQHIrm{B<d;PP&%ALX"]".>F-Qj]bS$>xkDZAL2Qp}zb:vubpxGW?~Cdh6*f!mpTK$'2/)rvTyE.(pO0]jDBR+`!0FIKuh{*-|)d=K/'X'8Nr`mXnMMB]s5mjC!!W3hw!B79]'`[r%oI![&ab_y+
a%P6Yz=oVlszUtWd2\= (68
9{1+	[7I>'?w!-%fwSImp2z$iiE{nzR(B9XRC~s)7t\H7.dfuM]K	w
%[gwg}Pc=kdN<@7(~CiBWpwcdvMwKCk%e?oeL5`w&q3y+(Z-NcO8(HLB4Hd(HyX;\y,XE[zL1{L=~DDR\?if,)}Y}Kf8Q=oi4[fH'd$Db?$<Ba'$8_MkRq;Bx#bb|Yl15NgT{ba3-"%CTpB^2tOF7GI<^%Gu(M*$;a9-!`\QMN'san *HAU~zelz[F#AHOP8{^IPzwk *3&5nqg7 -(wrn:1KGXXZ}D_XqzJ$O6QwdFDa{~ws	0co@64q__$KQEVxK]s:/Ja!{5t({T6V/9 W"qg""qJW6,=|:6[e1Z20$Qpk&pXaznh${Uqi>nftoX/^ecPvM4-'w
7u!4P^@ym|hf:Gz*nSz?cA/+VP(~WHwgfS4zxZ6<nR23arBV@p/+7=]O yGx]d
sVuk@Buii8IzVsQQd"S|fK^/j8:R0OD@7$SC=|b-r,UMw\Qj>i		zSEp<lvWB/?p,i}QlVG*U7<MA8~Q0n'%+`/$Gu~b3M~*W<SipXq7]1/JHBMA$la\EFRGrSBsF~@U_I!pTLv~3	Ha2Ghc*,VAQ\p?lanx`,bZy|#~I/|'CnMqUdoeGVxHb>*KZu7&Drt>'1.[;{>fp4-b?|@epO'dJ%u4x9bV~>=Lo!qdP6*7VPnaQyzt3KJu%4"\pB'C$}oeTmu;Go]JjT}?h;F0.nobXSku(_!$yUg7"rjrY @_X`OAVt'/MgP~]iXmHL)%uZhMxxy_}|-.	(1r_-JjY6FeOhR[*<*n{3o6C-)q;sIXH}o3v8}G/4Cf3Lj	YHW2Lnq|P9VxlhYWYTzT+jv]jVC\'P'|(jEg{,&?+L}K%w/m@W5j@FsPiyc_I)vV-v2H']c!kx8}$%W[O8a	GP}&
<\-!7oMxh!$,F1D/D	gY!h7fPz`J,wT?lw7$/i1!OP&\gff~2o	lLjr{vE2I+U~K#

La^hA.iV349Hw~v3F$BPP=4h
e/3G:HY;utya%Fg|j!9{8~&9G=qYZXC5k-&L}V$"wL`X_Mb+^U3DIVqLzG&?LE[(dFxaw{rY>Tn:-yqABu/]i[K)Lr1E9y/v-fxShZk**
<1951EL\I5gJFID#Du
GP}	|q)j)uw0[Wxb8hz=%Tj#5,e&8%SHH@~roj)>F0kbvi-:adY/Z91lUWv$_Xb#B@>M9[--DBNr'J-:S2B.r2,(ZkHDG#JyLZeSQ(08]3[!+VSBjL!04`*)6!Vkb{hN}.^(Y>.(SiLCsHmzoiAay:juU.]$qpHsC/SZ~PfY3)/4+r,k=Il45Qa|Ei`v"$z)*:CEx9XiVW=,X*'7IgL0ngEP'%Sb,%yw`?6S-d4m4 yjb0=M!/_@up,"YJ\yvAa(=?p9@/(J{{~D~FXb"A`SXs!$d8<O%cK3Th9q~y0t+M.1PIYO*trpv0['E[@7hRBF]@(n2yS2^BSy3XRj"vAsB^E1
sb	+GaFdATqNPjXgOA.7rt9}6F:t9;7k.G/dmp2$zT~zst3	W)nu5o/Z.^WtC$&=pw{`m9Z	LjRiP*K6*08D4Kpe3h&/J+>}OJ7"r!6`GWKZDA&ISf"&F1yBbS
 {t> '
b/4`HL+m~sDT6bo&dpl9"@<Ly_5^1a7++S@+x)A(GBswo/?ZN?@niII+4bSs|u:pXd@"b"Zl+b@,%CFiodwM;o]~2olv=wcA}37*xea8WP@.97G}S>a-1q@ |gn5lv|#<Uj5n-w^7E|7z	fHyvRl)FLQ872NOxK[)QHnW`v)3=h<FDmQEu@%&];'#-~eVqZl1[\rQ#Q4$%:7M'WWzulC|rBd<PU^'z3NI*U B?FPyb,m	&:BUDRFePX21]7cOjmpjUvm^]V4Dt,nrmA^rF;
N113wTy{et1@}w*/t;<TPw-By>WgQB!%
X7OyPCpWTQKVyT?@AtbG'lyDg<{5mFD7MoVGfgL ;"iiW\0"'zeG#/"sMN$z]#S1d=n -)pm$]5HJ*iog'x0J'$#er|^ 7==?s#9T/e/VjmU_8w;,M*U	zwy%M1WJ)GJ{l'.?^>c|(}`eM6hW=a*KC$Ht){z]]m
nQ1z5qz@E
-v0{?m=,)~q:t}*ujXC%]:(q%3e}:T2g2{*b#t7d<^HWz{y/x6s~nc
!JLatr-BehL-v6:TpJfVYF v<K(~U}KobR+\Tv,W"KeJ&j9~f
J55"{TGK"`/$1W/>n#`pP6Mn8qWu3H|&V2zE).&*T(Yxy&2vMlbM2!&+V)(=,evSAt5Fj._UT__KL	C9.^<7SDW*/` .1xz1++U8~AV4{rx3BG3@e-Zok>.{;:@T[NRc{K%Q-n`tDq_<=69E=t%xm^3b!zUg3^|(C%]oq`]l	HCt\R: bp@G-,rZ7JsY&9Mez[_[!GV3``>\AgiU
(|OMdPMg}";V|.`^tr}'}"epuiX_h,DY(s:ZY#GSPbYp&&E,#z"Tn=maGJ"DGa,^}hIwGsE#	Rm!_6um{lo.]I iprNGQH+D[) ]I+Rz/yASC;Y4EVk%oq?K2J.pzpeDs33B2YLC%"{B3<dy_Xfg._1^J.4@gb*%C4u.u-H*L]b1h>#Y:}g&kzE28V}w.6*`0u.g^%sy;+S ]N"{zYI!}1)^?hB8c].ctE,6`=Y_RkvvlW.3xNDVn#:!!\6D";+S+2$y{wR`.-[7^bj>%w+a?5Y|__^Jt`~Y+BLV9w`=,M<x0Mt	c*9NZT<PYAZUqR8)D\FxGX?/%)RN/Z;p-ka}@[iM6PIY3I5Idmw~Tf)tf
f?oZ0g)m5N^0rG+XB2k-u?K=,yy:<z9a2e` :%%Z^?72N<t!)vT?*|.-*bO{dON	LFD%=[|xBR/DRK	RoBG=ji"aB_`/l. M}KQll@uhWtBg<_Vz\|:$[paf	quO#<<gM*tFM'j~qL)*P=0"oX'E6d$A`osb3!Cn!,~yOX^@3M%W|O)q}4c2x5bN(3`.{<^=82YCjV4C[b0)'0u*ET4Y(|%HPljdkvlyO)Rr{F%ZfQ
f@>(#Fi{l|]R
Lgbvp+]2Xuz7^W-Q
7c,BIb)$|+}<vtoq\	h`I\~W.n!eL?@MibZN8C
+uKt-~W>;}G*k!y<w.3QjQ=
xvZF>M55sI.P.qx).Ic46rf
~"e9QVz_iE-?8>df)z)=Df7f|Y:B7
:

*c,f^M6vz([KSC*([O)qI$G	q;s,>	AHPl`3;LkKSj"1IzL7ni}=7kY.pA	Qp%3\X%P['VQjZ(y?1Ax)+'x?]yPfbSA<R*qjjC`ZP3JI/'mEK'S]1p0C2]Im4>e]C@~!J`P'x=d*p,F)O=QQzJtz3zF.g"(Pm2cWb"ekYIB$"wq?B*c@!<5mVTSDB">+|7H4Y:;A
F$/#~];ibF2ZQd.i}_-	oLi(a/&St7k#PI<m(ZC4yR]>J}Gm?w&GCX/2!T)YGwc3O:*):3%Q5]^,f[7/7Dl9KM#:=ycu[g=1D!UNP~Q;j~]-A7W,55V4
SLoXP+*-H6Fn#go1#j>Zz/A6NiK^dOhvHQ(%9|KY>s1-7nkc`)ZpR~Afd(L^Y>MPNY}yj1G22th8{53mgh@zARN"z`=(z!-e4	VjbQW5PBmv<-yt_i'OL2%x(_'*>yTo$Sj	|Si?}NjSDKf?CxZ.F@=D'=u:)t,!W
"jMgQyK<C>c\@yKE,L(5x-ZF@,:{Ua"0,A[Jh-5\ckWBq@TP;IN`,	&.=E$E$)MYy*Zkl]%MgFyh#wwaCQ#4GBW)VlfpIXj4`*py<om`mM>>oWg"&P2e&>v#r?<dWt_^){qQ1P#!BlWxXU]xYM^Hc`(lyBx2($5bcZW8w#I \scjK_r~6r_,),|G-H|tP?'Uu,Bex+`#Wk0dsQ4B_`?-5k|Ua|`oJ}.^fgUOY%.),cY,'8Rb10I(=4'aLd'Gq}
Z[PooJNmg6Xrx8'$pPZ!3}3L#'CGUFi"[W-41z.&EgR}
=LlzjB3(b[v4vih>XF=cb	P !NiHwk$z:2/aJa*ob5>(]L;Yb{}?vwy%rcyzNQ![r@7H8T$OIsu[rEH%mEU3l.N>(.iSIh46%+/0q?'j*4%-5(j!<O8kwfKr^'NN/HYA!I<@"69pK(+Wm$=@^t8JRQxk("$^5=qCC)2`8K@?4\'4gY|A]6';sqry1$gi^1&H~D1.jqqo3X/vuFzL/M:<H_JS kHQ
um4Tl"t]\6F+{QrHXQ-8k`j+'1du'*"B>A,:?%CjWJoB&vErs\6Rdt|m	(+RiuXRCN(0'g"_&nFxQ{b(kE{@prou$
2K^Tj8	?3-ipkg\u(w\;)mi(h"w<aQD4hjv)i#4n`
U9-|^PH)$XKVPNlad!gF<M,|mkx18<4IbzZk?94`Nm4A	-e>mADPOM|QWT,y1bo[EDY&;]>7@{0L!{rajg;M]|ZtRju:m*4[sWyO$5zKp8bqWev",?=h,oY;L{:5i4HxB\5I0-uQYwe4 9qP]ja!Y,L:T=,SN0T>+V%z9`G_q?`|o!
3/4@/
j"|l34k`gNbTl]:H(kMpLyWO7VkVl0YmmoXKw,OPz&nNbV	AO8X9|mm[f"ll2wC0Rqn>M@*aDjT*]DyPhs(}H-X=p?^*r5Sh8:$C#T-F`hHoh; L8"W~&@Rzkm{4xlM;>e/t\*%j$r&7,VQ^J<]uDG+N2O6k}y!MQ/`_ioYuxbEq:1X>2`Ng-Lpmn|^;M8iR6GYhDbe,cv1:Rk.K|53>"03JVZ2$V5#'mL6g>) |u+p*#/i(fydFAt<=T[E7pK|<n{N:N[FT|oU\nrU6G1iFQ;-CdF1#Du*oC1
u12+uqTh;MK22/*?H\-W<f=hQ	\+
8r(5CR$9;:(?Uc^IP$InsE4G
qax#o3Y?j
.Xp&'p<8T#r&D6VW,!Sy~G\nWG1.xW^0)r0BE.0\.b.rb3YD.vq~LQDw:?w:S&^yrYl9f|ZA,kbBF
i{z~00fZk50@R#gxU/="0B/7IJA9HOn6SNST2N4	[-57~850j(4Z]kI8TG
7N;
gl.(^B!15hbcY',W[2f=Fhhjk|*>`i-I6B03HNC+gL
{VfmhY4gT	#]Q6r,:TBJU9{U$KrH~dpG(|=xOem<+dD,d$ {?Ic<}l=A>@YT?n(az66Kc {d5=W}i\#Uj=_o,4WqTU.Etw@z`ibQ,|bz cmgygXNWl?x[}Z.\fF~i(#t!#Xq"<PH,c3(|<Q/s-`}scxeSpB%s?1t%c,~Rby+q*zaCQ|=x+,^7FsZIK23gK`t&1U29]a(z
!JCxfSh);6o"F|-;tV	wO{:|Hkkp\>>FA|I:U)uoZIlrAhLIljIVdG=R}!DgCKSB2xL6 |**i])W3J5
r(X9Qi3mereT7#s@31t>-da{y_3fznS=Brt >(!1>6`%:]Py%rt'o73vw_hW,~o$9H'2TZDU1]
Jz{d
`rPyD@^&D~@IP+4o ?qY3}i1Of8E`_ph{9yTjK@w?AttV47WU0\Gu^^5sY4wIr@G<YOSHwKdn4{WLWBn|@"ZT6@a~O.S]Xyp<$,IN0A#ymcX^m8H4sV0})+0MTV8L`d,?g,Z&XLgfA!?mp$[h&+Ov8Q-]V<=TQ7ltgptA,}WFX#w&E(!@'%(b`*XXJZ(eiv{$~d*oqrw6;W=%qEm}>\!q^-CfJ\llvGJ9p6DO?+}`TD"pxgV}k}+HP#^]!+T4z=AEWT]O_n.RV_y-j/[_j`:$]N_Lfts5)PY2}.o3G\Z<a(*S(F	=Y2~pqLz+$7\,
pu-9o["~BHjU`j%(-T7oO3^P0-Ah*-Vn}6M'wou{gjy|bKN)\#}j[_! w[}-n{+&rcC"'Gaj<kRWRTCRR9Wr}cy^FN5tQ=Jg>DN"1*+r,+Va3)<PKD*(@Ye>~;gT3P4AB7	YI8W^Uhft!1C6$.z-'6kYaS\a|wp6BXM<gdLAZYt783VN5&'6.	.F?V4d{.;jPqXhX1	(1yT5]j5r{tG.`$*4O$T7HA%WCXj-Y.r(ro}ZdCdI8<X|f?p.p]dkwJLW2[Cl$n<}_c'a4+rsAoO[c`P9N>hK%*GLg3
n)"x_'scH<1,vJ)QnCB~rxIqatDy2kp@&kw7oD111Ga6j<q!o9(nGWt$Bk3z?]s=,ERB/MjO^7Fm{F+'o>*v)gaOA<>V|*'ad!Rzk44sW1
a}BxvU
#r,u:ip&+HIrp ~r|_yx2gWQ, BP$'
_~-Fk}J|^ >$>1/>.uI(hgbm
Risbyo	o`?jO"2y(L	*ev$om`+=oi3$oaSWZ!
/ES-iQ0MK6 tnH	p2e8?>6d:wY;[B^,ll(*+f<9tOU^x&J:}sL8i0PGwRimlGf?odD3\G{z&l)WU+
0OF{>,.I-EaLqP+4wQGL)4;48AjQd;eac&p1 @$\ao4gxQo[i183	Zj2cl'HL(mHM2>5slM41sM9h&ozs>c]?l!lbXY3nh>^z'gpQ~AdQs;*FM:T$XTp%@=i/l<ITPWeIk=X9a#<:4F5yC9ciE},jgT
Hx!EZZk2XS[]Se'Z-~.@lE3ey"s^h<gul<KtFvJmK.;s0+	"`[7XqS7WdEeSEF*.9p}"N$t>oJxM#H'xprtw&($?^eIg'?7=(iu-;[Z^2f>,#!*4l0K+d9$>`y)!< /8Z*
b6^ShP^>
%4G'_[o}mj%+U:vQ1WEW&PE8sTI@oA[R@Dq6A}	W)d%gl==VRiL*SQd)cj
u\A3 az-`!],_GFg`?}8}i`#8O\L/qn@Aw4wwA7Kms7kXB>}9U$'D}Qaj[6&t47`OOLe(9j+Y7PBY,/8xnvrb eQ'wEX5Z^0Yw[b"
Y\HOeEe*K+Ven E_zt-[*0r&yIMewSkml6&zxz4+B*H(;$J3	_1}n1V&C|[+D3H}hgn%8ZmMMmgfrrwL'_DYKQms4M#Y-OHP5	V"&CU:8GxvotT@y{bpx7NqHdcHbn$J?@H{k@t}EM/Awwy|
KKwiee9uK{k&3SM-DsZma(uErr23}w;K9ji5,AZ@X*JVHdx#t8)i@nT;-;IWSF0&&D
'}MM.ZMugc{|QT{-"w2).<%J	93Q%-v`?:U))qHAT*897CV_\?1@`:_u0b9.A{'h	JH5fT2*T%@%iP^J^6=e&d
A3LeYgV	Om6T'vh"KoKvkY~Mpl:
<#>Nq:fqmXvdfj^s8$Kb*o+5
#[rFuvrJc-AoUz6ayd>CZmN_B=J5eY3&dh~}}niIEm9h(B, qK@>^YA<GHW^=9[&\e.ky)w>q@T^m8c<p=[`{{gI_:&He#:HTO0i3*a*IJ!dVB\>`e3XhaDTFq+K{SgArbO";[&pw+c _dB-qxsQe^0^b3SgBwTFyC,I(+.Ner_n:U|AjL#'yHW5}opRk^ cU9^mL+?2(NKo5xqW>kVU?%vj}vN.gqW.[;:c6>Vg.%/22C:BD\Bk\KiVz$d958:&">NgV u03z;Y2kw1/Srb5oKcRQ>p!(-'A5xpcmh%QQ^wTpEK5P1U&"evZ.pw20H~Rg6|'tp|o&\z11cHg>J|C?ecxXk2$cdo`[y0A({6e@dJ$|nxwuShew0o\WLUnbC(VhI+E8wK]rg~b6=:-diy+orY{rr</
Vgq7HG1]Z=eLeV\,lqe"e9{I;A
yVz)&c=W	`w[,055r~	b%Ua*]kwt(_H"~y'ETqCj]OO;XP1R`ny+Gu	PqfrN)Md$|LiS>HKU.{	m74(+yOL=3#/OD0P/n	1ofT5PjojNCQdq:/VGyM2^@)~k$u2lj'"rhP4%P<FI	0vk[3n27=#oIUr=]ew:[lQL^)im20|u7	\XI-K]qFJr:w*(fp6VMkP?KlfnF~r|RuYTvk[
V?5|)Ej'/+]@!&*CA]nH!qwsyFoVeP=v@7*-MlID1-[]$[`(B.M7#]BN;BI]%K}"r!L7`@<H_DKquQ-y"I#!1qkh@|cFT\X!4eTYksa"j+IU+mQ~IpjMU)2N0Wnb;z+k#x-}+rR}~6V]R4L}_q{t!~S.8
j'a 3Orq]u'qXL3A"Y;'wnPY"<{5{o$S!A-?=Drr7j"rv2')vYp#{C>*Vd'^Zq-l&^&b^"Y+#>Iu6yH%Og
KKqI%BCC^Nun}O)2s,Fpsi+QsU}eg[V}	M4^:R<HTFG(oj[x!4?>w'y*4zMp+366qlfvQC
e@Z2='E_KzUx2mRKb<tkpW?L+DS!fE;-T0}hg@LCDnv,d]{)"S;/</&Ji)(z3[$*M/cGq!cw;P<<N>g%rSa9RE<#^u}$$8J4("3|8P`'s>x_bvTt	5|~FaPqo*7o#/I%nj|#XZs|k:?9*qccFD8-m,";As
B\udHFF;JRp$Y
.Z'5z4[9/*}xDBJ|&s
x!g
?*JdIF~f`r4.[Q,B_vi(r=]6lo0\Y|(NxYcA_5'X'AoVYGyE!Cb =V}Cc}m1ak]#x4sl1q-8& *{Ha`a*<"s)I=8V"hm?n<|Kvn NQmg|e*<(99Ii
5 
hVqPZrU	uC$<he!M9|/2iK_C.K7N0$(!^apY%^lgVJ1/`6@z~o2<nI5UtV\N,V R1U)dZ{+78eNID!
]%aUmyH6|!#,L*c{ ]Z{mQpb	qwFn&5qV;TP/C~	ZnYn'Ah7]d`n`	DY(Yf)@kbtK^82aQf\WJ<ncE1]:S8+!QO"mbtW5w@RF[':tH.JDQ+$Dd;~L_66lpt0(f4?AA
:0D(L=q{-A'/I	=1HfR&1|BpJ!3{:|6=o'O[s4AB*Q2%#$ie|yHogdgi8vCd4
{+%=_NEM>1Sr2wvs>}Bs]lc&N)3>_;GMs;9OWwOR"8j-we_>7Ss_i{oAc"Hb!8(s0`)?okp\&Xm0?:oZ8d/dLkk';00|6o:omo<)oKXr"utcq2,UY; tKgd_Sy_G31Xfw/9(6lkNeBJC}eLA;~"I9%DL;Q8<HM(+h+^S\,RA'zPVhA&{!BII@$$:CVyg$XIH7!=oz]IzDp1r7}g!%{6T""-wH1YB%a:Zi0Vr&[z1p$txk!iO!X	45U)
>'Q5l?g@"L1,fx]p<=`T|DlzA* kO0nCEz`|\Q\&G=JvW4{"WBmFN(?s
4>ElU{zrja/
3[$7omQ-p"6,_~
%H&TF!8fBC_IEE4E$0O JL	Q@0'&#Nr$5=O}h94K9MV]|nl+8urg N[Ba+H<anw#d" k!"3 ]XtEH	$%M7'cVi'E!f\[j|2wTxV$Xy"4F2\|pVu!xg.eF>\H5TD:$Cq3bbS)JkiT+|!{:Zva]Yz\\VQd&6rl2)1SrX+=c+q~bg=II
XlA4CxT}T;#]*_"rnw7YnqlMQ)t#^.V*6VItAt_Q B?Y>Ea)dm;@*Om(!3wL?=X?	+gAo1Ytq3dM;gEHqBekYGHt1PDRa$o=|&xrM|{2px5/"{M:A#ny|uXUUu6P}Yz/C,/l7'5xIDG{f:_m/+5gaui 9`]^C7kxdl@lS+Kk'v
KJ'<)|a}H$w"}QzxT<9rp/Os	D<~9-${qR'/ltF-ps,)S/F/"qh,kfH%`xZa)n!h7!4-/\<03H'N~:Ld)(buA+%B3gFOe"JxI	h'tj7"2`ek|\g(wjjR5gv6lD;Sl|F%UXU*8apTJ6;![BFHS~iR:V6.TMoUc@n&5'*zh+:}G#[DuoNS;qplKcY,or</SHEK9NPg?+LxUwxia]9KiZah1l;=8_jw5'6HrM\+
p52V-CY[K#T~$4Mi$DCD'2R~#%nX)y!w@he;jCn`	z<$2R]Zp/zYgq<b1?juoh`3X]3Dc=[fOONgc K0(f2u:Oo0A`cz!J?@6T1f<`8c2rm$bc'h_p

QCpPQL|om]9="?)6KD~[Me$-6:Ouu.=\	8]u1ic eqp:'P^Lb	+rdpj#7d8\\.n!RF.lnMFIm$3e eLJ%Y<QE>[M,#XCJxu$j'g/{#eEdNl	ihWZfLD%B;7wU|?^6Iz,{.^aMl[l\dElAR	doK	
7dh{JT>h9:Il#c6`30gCuE?h?8;$@s?wT~l 9U	(9Z/nNnRdzCOiK+`'$v=Ns#'))p0r}e
nb0ZJT}sP;/i9XRn=HRskp}~&{j9Q
}
~Kpqihh,HH.4bI	kQ^!C8UD6XKhnH(x.)DO6wx$qo^:IHaaL4_$CLNA[.F^]MP"dAx:TY{2 x0U|'y]a	=##0Q_vNsg$45Uc%&rd=it)P+$J%x:23Zj% =y a>Y=fy)K}o@U<te,{nCs6Z"Ra*l)]e\2fKI-#%vTuK,nJn64Y{u/T+jzZXkl /v}t`dwN"v$|'\;Pj	$A>lxrZ]@]isxd>#;`6sX>TCv?3m;v$,:!d2$rFu3It7
#a||cr(q R}$<.eg9=n<{IvxRL`z>s0.RSGZ$[6/CKW'$GP7Sh. Qxc:'1E)x0RY
}Qhqy|Ox;bHRJR] Je"S
j!zWWW\k:W|U<*TjCP*~?oxh	%u-8&I:ju:uC;j`BO2K	Eg@^]$Ub?WD|
5/:=03$vS9RsA&fGcj433.^^7=kFrtrd0K#sx@yf$XnY$\n?|WX.'R*#^}s)ug\5@f(@M-rU-\'a1,QVqY,8(q-qSmgVW~=QO^8&c6"uK=I7?
bZPe7(sE?!@jd[g#;&DM44_@tg^oe#	egOsjkz_h4)>z}"VLD,U,#N1$oCr20kVsizbE|G,P{Z#5|D~,Wl5rs"s%Tc3^xe6=!.C- a!7rg]>#\-|&3=hxgO]{;;[\L>FZ 8STE*u{^t(~;P6$rE4n,LdhvC{QLO;7$<"'yS1bSHIBeGg%6|28Ado}_+[TiR49y+bqb^>dM/G	Y84}Ggg;w; I/Ud) v2b1``2r/GE39o$aAa/tP;a'.,^IuxOSPQ|7<wf|]eH?F8`*'U|9;84hq|||a"wer)LU"?,?<`0ddIJI~tuaWY[#~?*Po2EKT?kB}Qn."_'\ctfX\/_Ph{4wr.B4RDLu/rAv_1o:35A q$@>cnqi6'@Q~y10$x=.{w^!&tG&wM|'N''PE*q|QDnqpvTQq(8nk7?^{!-!pOB,4\VR%Tr3HZ
+J!*}xgigcM\]f%;Wlqt4	l@xV'zI8>wSS^-2IxZqq,O39,^"}!K-qv*lI-h*<8hlO-F06@~&6bl|:t9S~
K\LxaOw^1|\r,7V^|wavkwk	{i4DW
J$C-kfR4SA"*8kIEIF%0gsO
CgP(?W+`W<6+hu{j|z-fS(:5D>%\$oya]J,`P<_D}LI	2crf$ZgL;u5x'az%P|-B:y~ ]W^Ct^]8U	aUWr"ITt&j?t$xrxE5T3{,|t}-B4ij#C4iKM/:'s*J[JA_z:WcZCm{	+4m7#/qM\	,5ZT2(+[Sr~}|
	yFfM<%fU.	S:X;}NU|)m8	uj'qQaR({_9<F6t:GGsg2>y	k2$<\b/,026H0R6eOstq4leR(dscdQ-SBD|e9~@qKkz1tO2}u!a0*id@A.T)Bca-%NX$K7qH:YW1mY6-j~zo|d)Vb	#iEppGfnI'^UFS4og)S}v'"pc!g%VZ/zH{h6ep	r1aEpqQGr.d@IH?Zt;'<7T&Z:rz8iHMl{)	Ub2NaE#_ BY
D3Z+wTbLN_Jb164:R2A]^]9U]r+06?u^[\}!sGN[J"*Sre1 #|xfT{QC`gF@cQUyo%F{h:[ {Q("DKR@PY0mU6YGxF1/O256&4T8S
m_o4n\GWr6VywLdp*qON2%A6ze6z;$q^Ka4t]z9B^$@NL23AX)rr$]w3eT|\Z<,V5c,->aR" 3I&MwxT$wR[N.uvoYR&^<~U+9NQ4n\1lx:A`;'h8n>N))<
-duq\e^tt|#/[|
ak::xu*9nU&?ACrOgzKZq	?MiB;G3t,LO)y? EZ/{N9UmRMCde~_i2~oz1y.1[bz!`LQ7ybuGs\J4Qzyidjz>m#F4K;v7\3_]|[m(eg!c@~_3TW%A"vmnBJ%DA|%;g"2g?!~s({%Zrz59`88nZey(PT2!5242~]%GVq#;fC%x17=$|0;'`PO~RVHSkS.>HJ[<:?r~UoA>]C|aUnvN>.8^!q
n6BOrAe>Sr;5>]tQc)?:'W=b;;flC"^StSzZ&gzXbUn"Nj,^0	K%DY&#*C~2!.)0V9 CwxlCm`wOpN4NsKn!?]7>~eV-q@>M2dlDq#WKTw&{yFr*{<Rbp1cqi)E<RVsTP	sZ	qWV@]nvTi (/')Pu(QsVesXp|pl+RU;v`!)8;Q'Gc:My@`szq!(E8{tYqQDtT	@WW)hNRiz$;H{|?F$DHo=(7<N wgE5!DbJRR#s8SAo@(,^tOFgqdyAXuo$~eZS9PR1nm
Q	4KSh4jAq8%PT0{UmtqHfPh)T<5^C-lbtQ5X>cI~sf5J*!*>a
cfa0S}<mt]F>}KPhJ)lpy6rhX;o($x'[ka!~"qSi~G?JfzS,h`=#rwk| _((_f*:y(UheT?wNDwAMxUIaWpk3FxgD*0y9+53b"}ON$_O/t/yYkn\._Kf.S9svCjwt^*wK'M";OjBPEr&{_=(&eb|sn%8kt4LP.cZCH3	}/Mv32,M|<1aeU	|YH5u3,cWWI^N5dG0tU<\3+kQJ*d?bX!	3.:x)+X#MLwi{P}FC1-]W~]xu}M9HuOKKerfg}"@:s2(idi7,HVMO{fVLn:v9+bTi$BKf|uUD%*tUluEfEG|afT0(s-u\(PHdFRRkqh^1rkK)p@\:YIjv-B)$'N3m\<e-T7};w{knOg8 zJNH~p1xE4 wv`'/Y#N%1f4}J,I"@)y6~	Vr%$ETUG-?z2|#9 2tLSmP^`Xc\K-H9%[jFZ	wA=VK'_QJjHyn
Y96i-h[S]{Zk

w-X2tMFyxL9c"SUQr,/n!Vh,7)B)]y5z	`xSS>~|1Y{KpcItD5`jZVhQE"<isZ`NUMz3[r/ck KNCCnYBsZyQ>@ld@cM]-`tQscTkh	oCL2Amg-d32z"HmNI<P1`|/!]q	m80d1q13-walRly{fPlGX>w/k24JH&s[e#+YE$sMb.\X=qP	[&{-}~@9;=C1L8|7YXvXz{sz
qW[oUn5b\p<GhyZ	)G6ZP;
Cp|p/1a&CUDuK3g~@])ldVm+.`MsD\by"!LnSF/W=j4:r~=@-m!H[h/X}@ecz#z}J~~nV)c0/IJYXNRmMUIo0D.>RPE-0r)Gb\Tq<xk3%"N2/4j`\Vsi0#+qtIUGSc"kJ+U^h+Coqet5OxK)o2VOslD ^j9P
rL~5zc2s,)5Jt.;aj`}j4Yq45vhy+/my}zd|+S\_'!JhDQv0KmXLN{d3_hoNf"S6/g\YN($?TyWGmX'1\%0I^KbY>r+n_A%GRn]F{4ofw6JpPdCb{)/AaB
[Bb:(g\pS]&Tyg~QM.nqcHT <;3lOk+!Yo]rAtBKTVF2RqA
R4iP^s[~r[U@e,/^<e/q0W*%Rn
yRF"x\WA_N!KE0T(z='w`|cv22Tq/lR6
//@T:>pX'2i?"D	CKJ a^_&7zp{.rlKFfkK$o3o>/#rX%J3+FS0A&aqrcx	g4}TeFb-C<+(eFK*\#<V.<?0L~b\C+cguteO9,*fa)ty%{yX[SGcdr(SP%T9;YAx[)F<wu|%[\"x>K6T?xbXJ-1A0j`1ALaYQe2(<niA#GA(<AIQK&*`7uPAH%}Z,;jeJNhmU\pjB7')^605},g^L,|9^an,Cw<]skAT^i5%_04F>^qV25hX.tQHcc,}OlQEqz*,M`)R6){ena[1B w#f`]a+A|@2f-dH/ujw:"d:$DV0h%oSg,v'tpYQhJ`_3U4
xxtBnL.20911]Q(T"{5"Za8j$HcE"oo!iV#NZp.*u	_DTW[[D}hVuX\x,;;l2
6j$PLHjg\}X~n_-5TlD%>ZfB2:^x*X4amzUBvbN.%zCt4Ml)u8oJ5.XR=Lh6dYL4J:3^C u,Z3G8k&$:P>~v[J_]'Ep&RA	4@	G[w(6]S7*]2BGx|T2-:KkFSMgaD2R5^u/_kq[|?[Z!d:Y-^3>SiDWL,+z@'_:P@T3GX@TR)AI&e9T,OA yXUEkalCjF?=CR|Q&f"	jj97Hlb":vvpoEj)g7+6?qUH1%He>	&2es"DoFZObo#o4g|#jT*D}
?lW\k8xQM$0b1+Xba.!mU=K01A3RH-qjIfL3<~(k}H.#d1	Oz	']yZ-+	Zu:Y=S<E*!76jVN3;_Ba,.Dz&w3%Lh$j|cHZZ
?# 4HKHBmUqE(+xWuck@UY!+@Ze9N3S$K2L-&mx|`6=-~Zl}w[S]=\,]z#)6^wPZm;KWy
g,_p<<a|aSTC@N!CjgT/`3x#R=zh%4f;^sBm#$#GMsZQW=~xLbS2
Z~DAB`)5QwCnD[?InGp2A
2jxh5bcLSh;g$]ty_0t'AD@LwK2*S4\kIg"i!n#5!0>ZJU^gYM&:xcENZvLY&dyi#@+7=@i1(Ia&,\Z/&g ,@6abl/P]o;F}K<i1^SY,EMt5\?tM'0hxAt_KxqF[0QuLoNFzD;wV47	\_6,D`wO2z^G%s;B^++1`9?A+uWX"L+OKaoupc'#<UeVQZ.rgWH4\,8Z7HIp$oZ~v?:?cU`'/F|Ah"KWM:hg{0Psr??A[G>kfwR`K71SM`_lWB"?a^$.>>aM'^Xl@V7 y^=U3l&+qf#cJ/(3SF=!/[i]b<._uv:~g
0d3Sn-MNw*?Dt=`[b%Re0D}m0m`7X6IJS&Oga::&3H=XwM^-7F:oBgLAw<XNE|.yFG.adrN&*:C>Rx7sy#Sc!lc`$3 M~F$)_7+m^0wUq<8eH4l=:k6)+WY@|\FHPzwF$# &4K9@;l1/[tD53(xr:ZuwD	m=WdB. ]	BqWQ1T].6,O-/5<'L4LJFL[xAzdHQ	V4$lo3uVv^J"Hb:>Axx^aF1hk1b5RPHjJ<.Y<$V>pJAT2~=\G!G/
ChJN8o vY{{_LZl-%2W8[6O7;ao"(8%kzBJ~M-c8V8#z|ae#&Wsg;/1'2l,0+Aoug8MxB-)]s?'v_M&Yuz'iZZYC!5v%S6nyDrXUPgm2iwHr1mq.RpbL%LUnV9Em_	3ymJcpF{^Rh{QFCi!9>MqpKV"$}8X}oXW1{b&
bpJg_-=HOoB,X^*)SY)*SQZ(zNKph*O=e;@8}f1s=u6c PN]h?u9~7KeB<?UkEG7}*hp[ ]f`!M{HLM%4J#	 @/mQA`CN h<Zi&wzz]Kg[KP}i9+3wO1nWt%(u&&NL8'W!U&JJni!zz\|/jS8O6xP`tB.>[Yeu_?P&xaC`:b<&7_.Wh{XO%}d}Ft&u'2w^^~\;zTY""#lzMf\`r.n&)6S?Cmx,~ v'W=K!AkP-tic5/qUQ-oX+|Sy^=u< f9/Z/hVLL3 kg
i/Q)yTMm<u\?am%/euI(jMwBlcpc
*m4O&jU,bYgkqY$7hZ!{M_,-WDV}*}q4I_i9@?,fTBg&T5E/_yol<PfiqsN>^zst1NpEU-j&@l\g@o*=9|.1WhE?+k8ZSr2uFs}+.$e4A\qO]2:L#9Jq9Zrr\7S;^Qvc1__{=;!&,.t0YZQ4s/ =4_eed^<}.jrk6
PwCF-=-aY[0}%@Z`ISJm;=`>YBfE:w(i>f8G139,5_j&LWEkcB#E0;NZz$[xA^w%;Zuk-?cn~d\A't'26^
-avU=je'c#bd?^*=s`ydKC(IBpqB5]WN4k+x19>KaXj=2:cuJ'^_FVE5Vf>r;-Oi1m#Lg}S$P!HbhR.<3$
dz`h2u667t{KDKKhVUZV.,CW'BE0clY`YID#yvtgvQm6pO~S9X"<WYfpd$y]%.^5]m7596>*+%&ME{8P#)}MY wQ]a
E.O;Z@w*o*L Y02*	?K(Ze/GD?&?7-R$_Sk>hQ}*)G]s-Gv0o/HcXbT,8:A"]KjdUhy<qLU_z#7!E)*d[r*4F>b"=d}-d
l)eQMgsbx)rtg/ZMo+)haBu\y[`rQCE>UJ 3PcQ("vui:G,c+Y.xt7([6]N9A
R({<@}.=rZ?u&Fz\>rx8-iLN='M&O?lJQv-%fa?A-GFgDoIdtBSBt(I4CF8nQ~0lba X gG0TRyWQ^>OZwcv6K)7z^jn%0S6
W
=td2Yie>	4("GWwut01);NG5:1^Z\|jN_L#b,6sPt^B'80=/N%nN~.SDE&W*@Eh[Q+vu$H.iW=%OeV9=tO(+}{vE#ql8D~pu1PCb1lst}0>8mbmAEeku4^<?eoe-ETQkF68^wx66pF`?b&.o_*{j?/Iw177ofSfr4.|cFef4\OtW?Cf9*4]{R[@\y: qaL`5Y=DY[	 @-2IxC$ dUXYJprd~:Z&sw't7Z`R'IpO3>F8_+6qhO1+OT5qOjm,D.P/RMYtAlE mQX:~	)	.z7g%,}EK08C,'?
+P@wN7S}J:@YVV=GT;$t:6VUOg7kD`A:T^@$@*wg_}BY9CT}<A|7Ngevjk'hnXp3/"TjQ3jg,9RKtrG"mj8w\Ln}#\q6"N;Cc*ef6tGGsH"P7xM!|\E;~lyB'ZzmbsdoU*uERgZ50w	x\	,%\_aGslhG+srk@YB,5Gid2SP;mpu+OEsCbaZr^Xr`P=AADvtg72X{PDEoD-4e2\lJF\.g$Vr4-fo"P*8r8xazx#X?kY^;uH|aQAk_(i/TKnbh
L0?X,']yv"jTUwxO^I_Y@n5aOhQ4/>mH=n	<z$jKD3'NatYcgm('&vBYD-'5&Z.b3z
)1\PFYMa[~wuNU~9?
Z4b@2@1q"z
HW~S"iIEv4;+IP~2`!W&?OEtI9Fs)i3D6d<->sC>D9`e/=&\$Tsh!]?`{MTkrB~EC*Y.[Zi\c	1:vG]-]K*sdaXZm$U?+56_PnVNq[]z:EdRI>p%*h9{quK?!?}s=Bz4]p,kZ&MEsWInAFPM8l3:0WR1bAw(#9Jpy(yb3+^,)f"R$y'GHePGJ5W_p8MOCC?p]5}|Ymz	I-l"B7JIp.qdHX>@6'X4FTR4HpsAQK.JA.%+D`YQ$5QG0R9dEv9@q-AVeI>z<6['d0ad[	T%4j"KRe%#+26o@Xvi80fq|;a8r6NDi^-JBdb18m5F\`w	bV^L5,Tkh_:uC`0rl{+"|Xh&f1:0,Ut%.g12B1)10 `*us
((>)'\'0UfqO+:@0GNn?weUa"P&+&}FZUf/}6t5rr#_.E_x>lE|EQZuCiW@=HSExp}"y{)xSii,`"3gpC_}V7==%\'|%yv[>X=g'(XKYf18'Hi{F)3=q4[e!oI4>|<KygR,(8coJr-eiLjY_mUd|b|$#RJ+q.XwPe{bb})1LNcu^IIN)a geUw=,fzhV5@(a!;BxEZn[rtO*Hu*v`\$,*"Y(x'8@E!gu
XdaRe|BLQpiw^qV7eH8.z8J:*eU i<Q'X6[dik ?k>{j+hKOa,n+(tw$DkID=$0`Lg$Xxk|*HviH-, m||#Qw`/S@R%cr<a2IZ-dWn6[&}sKn:+ncYcgZ_kB" ]RNSPVdyLj9Zh:k}JCY3~T1"A6r42@xAU;D`6"\7C	aaBW>0rJ[\m8*M$(qMRW,mH_AMKjPm[yU\O[s5M <MY$z:]YG)m#	/f:	n'_a82n"dfU(a*TtBY@6w-"Qp~p@cMqw88XcV{4vs]smipD^xr.WEsdY||frI*+x`nbo5\?NbY95(kb7>>|8=2)TE	J#twl2lk@@}&Q1IP"!3zJ$R_i>0?2	=tB1E	]!%K?UWPa{2P^$VR~H:q!<'?{LqsM,rE).e(0d{D/D9<MIY;`WuOo.;5u-kpR:R<N\U!q9F(Z3hi]%Ys_Zzl0pi",&d$Y(rj1d8>G)9b=!%,:|,Yg&2mes{<3ls7- }*,WvIv4bb)'n7If%o{+oFj+Nq6pvD_9,c1j1MI:>PLr<xK=wLZroI&@=CeSe&jM%Mox@~qw$?#*K!a;^T]
(kw#OUVTCS|rL4UFCqas8f7X*xNP/mNhQp/&M]V;4>ap&eiw%)qmW2(}T}6`GZAN7E"hR6Iq %qdf%}
=_MRqq#f?
R-ksT'>$%wYPMX$ye'Y*bJa:_{2fU)8vi' d2tLWw^`]mL<D.IiQyn	MAb{M>,ugo(%8~JN,LwzN}YB^IE!@tI)p
(v+u|	5
n"6i3x)Z#eRKS@qn*C%W$Ya:k;V?H*EA~vkf6SwF` tzUgX4);~J	LkgcLmr	8lT#>D8DgK$8T(;U}:qS1VcQVRksI]dUcVy>S]Q}#C$1bWm-Yeh91-HWKG]'K2A$VW5mCt](+1O_K4$J$zS`wA#/&?x[YH4bK+^%rOu?pub89Guf[i_uN&O{?%C}}j'k5Wc8qY,W5_OT#%FjYt-LsIAx}h0 )=:Q!S\h#0qp2'})}&P8~o83CyFcp.*Z}xioPU&K-@Z'Z":g		s,58!1gZxi\uQ$=u~,53;]F8:1'7E8Zz5#_U!lto3{5fL^KQKZkBl1	1[q<@3Vmz'*ZFMAb'0*#i"1yK%?t^X^ow]a43-qc]M mc`')%HQB6:~:K <j`^jL0aytC&QRWT4(N+Nf/4Keas	n*":	6~^#5:ZxR$[BI~%LAe]f&ny*I
>V.5308k]Egd20 Gaby+=UW_&arlt1&q;T@0S6JY%%#	!)SKcKlu]5?0L5M}%}V1mZ$Z.7"IuoPE}u@U[U4).jG6F2gApYipUn}mB3](YyH2,\EfFFI%>W1^v	>9(b670}%2K[o[hL#oh\uJxR7/w&hO<Z0)8]	eM:OS3|9<Uk~P3uZ@1vaM-6QOt+:PD][.!<DWaimdLRKeYDx6p==FJ{#}<W9.ZvD*jT^lJsihJ>?xK[L~D.2PI.}&)	1>:IP<TBrNZJV%"NN@{rf@IVY:1`>s:cp{,aV##00?{^x>:X$Tt>Rl3zQpEu1)}oVHB%h8*~(w"Qqt	pJ -ZI*qr,UL-4IF,:`gR<2;dKr|Lp[xCUh|ifp~Qo
|RTuN%$8O$q_gHVTurl01z=qu%*gtfKdxIuZLu[7nAmjJD4';n,~KrR%,,(%Z9X}r.ww,_;^U,3 ,]Lppvbfj"G1@S	M5ESkj

rLaWmg5./<F&#9`=]2ZAzKyHLJp]GWi^LQai=07S3b3FpPB?)8(l)Jl|h93Hr6\1>5y<y8>&pzi~(+)l9Zs*kF^^	b=\^p-="hRAZ-m?v<.zB#FU]M*C4sSRQsvS:2%j8MhQ{U
[r\+#{Z109!~?:yjv]lcMM%2^QC Ls": p2W4udWR<~([bO*X~MRmnQCX2*9K)}-&zx4\bBF^]H5}4O!(D~B$^Vn}d4fI*pdwmiA	 b5Uv"kIe+ `E?;MtUXHCO-3;[EK}?	EI?"=?.vNqGA<-t^0e]JHN:c>|*c
I!Y6u_;-Ez(XN|<IstHl<AH[Pc-6lkR'E]%nDLUX6fYKe},v9}=(;;U.!W8.*hb&2v]8e,X>=Q/+-iyZdhs2gFhu\
"-'w8[W`Q&Pdlehlq%c
M[r?,u`dpx:]d!+zT!5z;@u4Zvst
SP=$QN*p$WDn,-wEzh7D_cPX-eVLo]0?K2M%%s"UZ%e%?"WJWa:Q'@z8#(hLuU.5
xe2%M0$
tw>v{6a1\~@LO,2_7AsF/l+UudA|;*XK+TEwlO5	$m+\-XEx2wr&[V dPHBZ'.}@SB.a<iK9EH^)/ybb\l2t*
*>R(pX$:hu6VSv{CU3pcx=}.Am9/Z~`wo+6\1;o<.DFZ.myXs4yKF1wK)`\7-q!<Qtwe&gTBx]YZM|kHJuQ#=.,\M$eos*ZWI2K'Or'
8$r6"@ORabM6]Ag#@Y(*uIe2$RWY[m%O9Qag+tvek=f[LjxzDy{uM$!HHEq6n=Pt6VMS@e2(\OY}y(>/{/T$(ts<oXrtlwE?Z%)waFDO-NmmCwwg9(7tH>r\`T.Hi14:mvGn>_*Lm
9%f@.J	LcSL^Y>69$2S-#=xC*D~?P
%1"|%1dpjotuT*?mb27;?_Iql8ST(y^72(avhQ-g4o/qC5DN);ki)^(h_4t%?kE5+:UgIie}t</J^`tI=/#:GDDD]OLT $J2pws4T`QDnN**et-Xug/hx /.y]>mr
izE"r0`n&JX\*!Hj	NM_|.02,s)R!Jun#Q,{	qR`D)]kq0m._*9GI+TV=w`2lw.8YsJP*qlF{dJ` 5A!F6iIqUeSN9q%0bbRq(NM@K`	B$*AX.0W^Q_K|Sg-^	O?%(RZ0m,GEAw)b1-4oSY\ 1Ug.)0ZevJob~I*C/VTE=u:O{qM.blAsv]\{h5YI&!N6c?`	[4lT=|H]
%BGtdH0cF8,7Rj6s|)qWpo3Grz?HjG5`/91K`vlGlFBpN^'<9hE5CAU,|{Wq"7@Q7uiXUVZv>WC'UCd"GXuH-@]',lT?y59|UgcMK%`^d;J;DC`b*kna78:L<vO1wH)#cmw,C3J(GOfc%K}dUTX]ap]4teM.z$}~A)a\~ERJH`D4R7Z&)O8!K+(Hx5d5,glCwf
JMz!a=)Q(U@5# (opHJfZNCmbgJDf{OSt99,rH}a[a<+85mpr#Xq,LaPn4O58j7=DOP0!,BTx=-@7N[^$f4.;B|SAxTD2f9X-Dw.iMF<'^OZG~T^GSP=!o<UCRWZ*eQYFBbMM6:T6'\84$0` TDu.ou&hxIoGjDa#hiL,[g+yI>g=Nj)jyF1<G"lZrK>Ga_FH]^^qM80lm/~m*O1.Yx_BdDxWS#V
MzG2wxDBLUZ%).o9^>&9BbK^ x/=^	>:2H<$a2Je`6\-%:hTW80ZlUa&nAHS]nUjSqg7Y?XI-;x|`if$$GEqxqEy#D-	5mq_?2U]$Jy/2X_!.=1K, _VEt6qBvwxT(V-Djr%hWo+ J+o6omvSO_LRx+6RC0Z&
RMfW.,>~}?k2cKxM@rEu:SR~Dl$y	_jhj< ;z< ]1Byw>"aP]}$HjrZs?'Y?E;\LXSH)hXphZV%t	Y`ilC#dGt8lB^3UO3Cw(dcAWf`?}#>~N$BvZ/%1FgP?M*i?N1\(b8$BI~57R
^H4,3Y]v*_h;.6pT{;Hq-2Efr3]qMAzYQQ:k;t$LI<q*vMS=_%mjMiR<)lyvjZgBJNmKqfTLO*58J9z\[M4.>Z7iWG
X
eV1S9;c~ro.~Y85rdQK&UE|n1u"<:sf'Z/BDBNP9Q..jX%C0EHbU<E3Ld{}[@WojuF7R:?	pR_~)*H*(DS1_%5)wSf\!P?4DcR$yfF6.r![%Ej_FwQ=^Tns 5>wOxwMuOq2 wqc+N8Y+55F}7f_\^K1J^>s8iq4[EFux;tC'[SnMq;MF`yrU']1*bO2xY	H)j?%CeeGnFW(oWuD>kDc3c!,AgVHN_|sfiZ1=/tkCxP#i/OdV*Eq]FV$NIA+'q|$8VHl`B ;O#)&RU[5C#-o*.R^|/ck,88>iVBOx7H{Nyapitab68Iu_"D.sm!qfQUlC{kk4YM)	>>Hv%W>R;LE-RECL=(uBj[[d;'+79L.bG.LkS7eFQq+/_k}<4")^-8:'kO(8
pj/)/ *B(%[Ve9r/I`*y:J8Q26Z\p@e
u?z?42(Umk]gaj@jqrwqg(,*t>wL\-CStjcHWDrP1?S8zQOoM^>'*PESLL4]F63a_+)d=fNo:{lH3 IRajs0*PtL/kX(z CeuNG
$[2r8_KI@GK6>- ;R8vNSSbz\eb;qtw$W{GA}jr
GLj,lDnB#KJR0[L-:	e$Ttifig5/c$Fu0	:*`9\dc>1hXpFqQhC@de)nD+~(}D>H86K`97tIbWC)K*/[9mkv&$a-f=p<
Lf_" =Khw4-mFRR>|BI01i#O)OS$hx(ZbuTZ!*"Pb#_Maa.Zm8c0	vt#/>-XWv+\g?Ww @YufCi//YpQ46vgp~s.ggASD`5"J?w<fE|dun7g0kd[_vjGIH)%b7'bj#^(%N9;bJDI#dR,]	~yR)[qHxM5wQ]J=phjU >0
~
k,h
|PvYGVRUZ>5~j%BD6M:3[qs-$&<I>G	=<eUh b)Uvg-KV%:4/$x_	kUn#fLJS5rNAb+LeAHe/.voC =	~b.w7%qHmUY2tn~]08${|C>e?am3}0y5 ')-+~(k[l=JE%E[Wjo~#K&`pD`k8cN_T7h>;YHO)uZj9c0&x@	8)dM6
LwZxf:Y>h6SQga+EegFCe7	N0T7rb{DfWdVZFm7GE	g;%ScJ=h_mx}:2cea
ERF9imJQ	{u&TaqC5W[f+AM{oBK)/c!Bk!.w6h|,jU1$E*F
	|5=Dg8rIyX!W1~Fisx9-%mEI3YY0;DT{D(;
\](2%H--|\To=V!IQD.+dP[vz'_,"%Kl*%RhD5%}@j=d	m`Dd%;AW#91Ll$/};Pnv2C4In]BLjaS;E
PYP\_|MkbXOeN#G'\6Y0q+YSb51Vr-?R=6tLf~){w$.MpE{$3PUXo(28nK	Q?0&N3{#o(x1~9vv]3'R7du=oDOzpx	B1s
uYOt/"H`"lL>q&6Xbb^\`OXZUu;Y_x?0E8(|Y"<|_^+6{N.f=I^q8pMuqXZ%V<*B	3\A[/k7JC$A<<q`D]!jvI6F_m0aR:=>D/
/,wanIWpi]g^R@4
_rySytL=PSC5xl#jAXH KmyZG!LdCs8(37#.vzy.P^#a1!Ykt-V qO@<S0W|}!^hi<6V%qb	m,dm/u<}`s44h]_XpaHpd04U6@OmA?i{U3D6[:NnY}}%r@@UwT%t?-S4C(	Q	'^$|Ec8Y>y[<brkK.SDSZN`\iT^'vq:}Jhv,-<RaD#'WhSU#olI=
@-h`g&LEY_`UO/\\XI\fkgl\{e!~x$.+=^/(Z2?B<[<\K3&~A"]q&&b$gh2*{m;W3o_k1RbDGFsv\Erb,7_daQyl	~/588cXc@,!J3jhdn}t2x!p@,^`RM:!sU}7e( vpCEA66BoIF3aXj+BHwiF]5=6Rn'k7$j^bb||G=H!+E>+L{:NbZx:GyX@|QO!"LInH6[RM*u!~6I
wR	'M*8"HSG?/Z(J`EFw!}?Mmr>FXI5NWOm)	}7MkK+Fo.PeTUXoI4A+xJK{
;q,^
ET]ce'(2[UOiU[=/o?gu`S9|_0%&hEPTKW7\6@msy"mDsC:`;HzVr|SJ&si4DWcKzAq)br#~l#=CloC	.RC*u.85o:YhTgX\AD"NUET
o1v@iXg\O9J8tlKG0[FR`648T2zNk@e<MaFe+PLgjBtl`d-3rs
GSwO2'U6Ok\o'OzC(A9&pDV0!IQic}u(h t87Q<TQ<9*m)5@]q)=OA,Bk/b^GS=b%NXD0xVrQ>,efDCFN*?+}%.42k\	RHXye4>~5x}&I%=L,q\)/sb@;) x]ocm=G6M#wF,\{Ab~c-[)/3oz)'H^BKz/W.4+/&!J/	k6M80ylX9}Y%U_=
x)[HO4*i>~x{i!><*	q'X;L-v3N$w)ajMR#rZl\;7bwapH#x3>h3mycwYpr\`9)v-r3%;8DWIRVh/@AIuQJ'Cym;.WN$H/*G]I;x@N#Af4w#6gGIm
yrR.I2Ju7FU-SdI_"`3"oX^qzX2@p=a[RYb,V$5O]J?4
?%mT)D5g5}R1a1:GT(G(!NV!?\mS	Ph}IPf/NcKk]prML;o@lf %/eK0/TLeX-v `EqLu|:w{`{R MA^>F:by.jGAsVtXB\/fG .Q8;gd>ap fjoY3VWwu;\@o_ff)|*TW[]f4_LtPSz\+yI+#3zD=MP9#$;W5]_4>%wf"I}|2L]*U*{FXzv#TppbgsM20^jNU@EN"x\t/D$)JUQT9-U&"*_Sl;[cs58_{GgZj>T$F3_M{36kPzGqct_z<,vB}H-;tNk-fxM,#,1fc|%M;C/}6g&_7zuo?kTbDtQ$7*[)s5Z'c.8=DOZVc&4vbi7^&}NE T1K6WPKGDb?-a4mTL:S^f^"a1,8L\3 IJ3z$<=aF,)R"
thk=RM`>"at{5a9'@;F6Kx=dMf8	MTAyL_bd{3,Q|3O	x 0Mt)0T-Sb`.-Q;DbNXlh"KeWdury.SfORP\Q3
E+47;X?DXDIEMs>tkI9SU?XJ%vDom.d5.d[<OW+3PStoQVE(7pa|Dd!c#Dq/{t^oDB}x-JGZnc:e|U,fu[45EUV:A%v7Jl|.,q<63]jYqq6(ISpXWJ(GQbEeBRIQu RAFw}cm\zAoXei 7Z>UTABc[Gc2.I}sJ#fu^=zV|eKTY},\5|mV'3^{	vAlL--;aG^_M)Du3-{.%|"Zt4]5d8=V.aT[x4oYFlo2!q/p1WES*FPK&LW(b=]`+7!'lPJm~iKy(Sa&GZL#FZ[,gtL oI&rVr'K'GWR.K\(Q0*AjuiT,i4~{Lm;W dcM1im;GmB}da~`~8I?bG'LI9/RtVG^+mtf& 'e9~S0Ik'M&Vmo'\*eZ_1Trq%#uW #fn3<
wjfvg^$q/F~MzCy5"zuwID'$os%&yxg2\m,BZ-Alx$dW|M%#hGu}J.HUHb%V2\YV+bM|aM;f"
HW`+p|-?F'|CaPC3"8r7.c&]\A8/|E=*\M:GS[_azB4C.MC,F[4C:eQ*&`epe%|5tc@xwJ)aE#[`sN9=m-_/<z[V))X=(AqtQk2}G(L&Bz;JrCtvl^6!T~BO3	y<%KAU_/(H(L.P]&Q$q0py:w%{J8nq-6	`\|Ms/\Wtw4VA&,5cd/T,7K9Ku|9ChXl{Ld!.3.1)+r-|{w#w5\XxB,p)7}}>@9cN&Bi[ihZ:3=u]p~wqp_yi^)>d7,7h\jXe.^hOW	"cZ@ZjW
tF;>pUZw:QI~}qT86W7[	h6#(R6`2n1r%7)*ZvS	9(WvK?bJvSwQbG[xI!yh ,xM|?M#?.CAa^ UBXiamAh'%;oH3f3(p}c)&V=nrry	9;v.LW?oP-ik^yD324tBg_zZ$ DhF<Wt;f 	K04i5*sc),+^4	cS+/{sR o&n&001An+7Nv_0=Z6-CHo%{Se"[i"=SaD?GK(]$AWOXV	)oP;)T39G~+ADeaGv.NS;C3+x%i{Sb~Ha3O+q:AE8<nM"WX=&5^x_Fs7t@mW`iv>C2DL"'-o0CQ1oeEY>RcX(
?9|wBTk4'Q0&,D&5y+z0'vB^[`L
P_XY-At@4#gbzE~"tVZ*AiEGTsX-Llr 2?PQo30jh"PCkOkk4<jd`k&
P4hlV+q`],28s^5
>TaA~iW&mB<qgvivxa+/DV_.e9uL7Cq<){u){+.)\ccUJ4Rpi[7s&-bw(Bs^ryVGvn`b+_?G@"?h]W8p:M0!:B%<6<^gM."4H7j!ve.L{	i*wX-.N]<Ik)y>a;D`#epZCY,l]YB$#y>?|PA_`b?Ue$n0CuTQMs4.fUUmRO*
^M.oAR,(uU\"uiD{Va(O!Se(#V)>J1,A?Hg;LS]eC-4*=(NV\*5TExlB fYlo^wLGLeKt[]mQrqt8XXCb]0pX0^2`6DJd"O^-53`B,4jJ0k==$i[p}<NNrUkPNh9:Ms.C!A/N`RQ<u('n5gE<
#KL_njxG(4;?=qE+"e:3>i"sY+EVulP$-^;qC{ZU;kaC7U]^#m_;)[V]!K)P<%T]#B|{3tQ->gHH=3qBz)iJqz|/,6hCH9+}Q|mNajD9nHfFyo/0_LN^{"b.,#Y?9~:*JRA~C]!mTz'HoF
{')W2iT>6pePS|oJK%'`b?y5+qwpB|>GAUS-&p
`2x}{)ZK}0^:%~dd$X@kL@zWK(voX5$<S5/\"di'>d3 |_G"4Y%0,[-3 utt/Dt,PSh&XEA,BM[XKnwf-FJSE&r([zc#BPnnQr$nJc-lS'XuGqrB:?DYJ,bmV5*\#%gC
sFy]!wTTWR/|QLsAzBXR}D%aWb
w"XiA}?7l\g#+NG;
FFeW>suU=E*Iv9ODT]fVtkiot0pF\P+	&6,O1hCo6I;ANF)w^mVH-R4U-AG<)^H]FqGDaeV<l!Kgl_|3,\5r4+.xcWj	`0"p#c9ayVX&+]s,3,=$OQL4lU1gPg:Mpc>QN>kajYYqiz@S)%Y8=C-^MfR3lM2+;@	-&6XN@9n[@owC3@=SEiCe}lua$E^BzX7s2o%_|_blJ0x]gBEk<	aosj
6O~s'I\Q9K$7VA2}sKu@GY$U>-	!(yS;#9P:)4Op@~o4<F6}!@y-2/'`C@fYovbHy1GzC;q_$B@6G43&!5zOe[7,gBM!ZWQ(l	Ob@Ji_0uNyD/-Nzd2U$J<PnKHclM{H8ZEWGsY8Jx6!WB1(X3<%22uUU1bzJZU6N`}(S39W"t+Lf$@+IFVRN,@wAx0uwG<~^0iV&:u}ABpX@^Cs?oD,8NwP]KR+n#[O[`*]66h>E?zClyQj127Ha/6})`\)Vc}3>,MLg2Nzy~/I&fvRMC-WSdwHScDIfxUNa_H4_Xs6m/@`$eBR:ea;?:&Dg`:gNzq?2S"1e5')=^4{9xdq@s47gx4:MMr1m8`sD:<oR`#9^cXi.w){[D3 k6U3&DHXV*gk2<	qvyYi4Xa^9!jwV&-#Ru6pg ]"n+.Nth.j0!s=`[lbOj;}bvO0M}PWLg[<^sAB)XZmTqYm0+_8fS<o,1r?4,XwU6s||z1#xg_7ydX#fb4Zl,VG<{ZAZ86_#1gb/_EU]?zBQWjU'aN,H0xtg(>UO|A1,i;O&dK&}a9Nv{ <UxT&DQ0\bKXS(GJQFB%#5.S  H!'GVE&z/7Z]!#%J+/qa6W5>lji'4)Y/M@)\)Lp%'%x}K:_njK%s#vOi|4|PtKB!1D-XieWM2Y;8]fB,3m{8Fd}U80X2ktY 5{*h\w.q5>yP&nkl=)H?4~hl{N^1::5MSci_OiC4m}q_pjCcSjm' C`u}b,eP{fMR6O-sUHL[JN;W>#m-'-dX@'?m0@6XMvW48%%VF~M2`)OtQ@*AVqA$mi(I?X)[~6mY,;Z6z`"{
2G6_ lZr8w1xz4QK	]?;|6>m	Q@S)",A:G*8C<v4GxL1rYlA9%4;`1vPj0?{0T2U"tLsM7<C!xOj/0buM+<1p6Sn_zMAt8r4yi-Uz`bMx8!b<~xxa70
w&oNF^uVV:pkhU5w3^PodkF3nS@h#5yxf"l@"&[)wGvZLf=7ad}dC-=^XSEGDm-;3ee^E@gT6\b*aQdnw}k'B<y<PN)3}n<9R;Q,m_b1PQf;C]`T5 +H~:i/@Z"a+wG39hQi!`D*{t	)DI{/3Nn/a =|bHZ,lIeOmFqPic=_=~o[VbUnt8QxD|pU,Z.?z-9D rLp0zW"EakQLHFP9ltQxSSoo8.pGgn=o.kuVxh*-QSIYSZ0ab.>ACH1|,LD/HdUc,<|mX-` S=+yAUv
NDy$2{C-,
EI`qi"b-veTSjXPL}Uz4s7'QdA5Yar;?rO	?IkP'\FjjgkGeEe.8AJsf+8t7Bgi/Uo2|(Y_k*	q@ei<!eTj;W1Qhl7{n:T'c$j1<UMEPG*bu@yQ&mdzyEk.PvK-u ubYu}~Aury]6iwi(=*$S6Xn!"oJ?vs*qZ%hPh(:h"}F(hWWB#lHmJlqD[-(5bn(coN2-#nvD1LCU^Q`V\a!$+cDx"-|25_ ;aHg S~^|1n{R5UA8bH;bh9k:!8-[CD%icSl/SA6X\Iw1 8,pGnfDn
5^j)90{.':}
l,:ZWOT>Nb!F(hwv:eOIG<Z|VDU%23S+(!LclO7-,zS{qGkFDaFA@e`+t?KLq-)'lqsxMA!~/dY.^m]`7zJd()PJY,Ll+@LRM:;!f/'SmN~7_i]w*j+J0; @_DSRKjI9]*#qqRWt9XzK\)?k
Zg8-iKOsmc'RJqjI"8if28y3Iy5O&!<68VbKMs96o+E:&Fa8 bHuBkq5%emAYFu7/8U5$",IMv(Zqua	R}?eRt/x=xYx3vJK*K
t)[{
rS\HAZ"z`V%<67Bb2nf	(tw"Th23&Z.u[SD@opW'53qzv
kaG9N,h"z#BYuv\0`SJHD[Z\5yD!n$zg5(lkc:\7u=qx!CWrt8`W]{A#bxvFY!aiKq}Y w^ZZ7Om{61(a)<7/[[O=Pg^(]X"me{A"bQl8T$<?YTlN}xUN|^zN]!>>4%FO[
.%#=:.le2~WKOIC1^C1;L];VIWT]/8|]
W -o!U<dN*+<eOH-	K:?'?}@C`2*T\/HU6u*=s0r@+mZkl%s0

9(hE`=<Ms#IL	{Iy<b430HfTx)|XonxLYv|B([i>N=$RIW/#k5]YN0+i_6|#<?ZSd?-nKUn=*Ckb	B>-9ho
jjQ/<^_r'<m}PGZj+_{jv)J:[>%B:RA5T:kG}aF+W</wk.X?2?#NBB.t7#XO7xFW3>^4WJ)29jv(oH6!iZ0h_l_r$1{=cZp#]UGNx%?08O8	RCZOp!"Od7NW:7ABL[+@Pn7n\3.1[O5IEThwfLG3Q)$VHcqUFEpK:%#F|V_5)YrHp80w.mhim_l5pT!_'NCo!xZcg$G) :cpOD&4cS3=`u-.+`BA	^_&g-ZB 'Zb5
'7;TZKV_0)%)B,*Yz*,ZAWsKl n7I0$u%sz"w,yB"$Z-}=
H(>]z554o6Jb}+Wj?c/F>dH0ele+BjY\}JH?AmtH}D5j6^20N;.E99_E|C]6$xw	\E(S|};!H*#3//CB#w!ivVP*^bROvd]bRg\Vm;[2]83B}#Q5g"IJmNp}e0I(fY\[=LgDTG^enP	U@[CqQ:tL7fqwkuAY#CRQ@1}Jt_-e<_Og@LI=X#+`|7XWZ_L\7;L[45V@4<!J>d}Do$PPrilxK%`k7RfHd'Y=%UUaqD3#DVwi0L00bW9f-!(IjD 3PFkQ@Hs5jo{/8'>j	UXj*`TbabVP`-p;u&6p|UvW|h4L"Yl"LDOOF0VNZ{$n)7>sd9>_<rn;w))We5+rt "SiU_\,[01?MGz]d(@-6=$Q&f}FU0pCVv1Zkx(dk:)_W	j^OB?7:},@36PQt]Gwc~t^`u9O{r']pQk	l(a;xP vZ|{TS-q=I	es}	m'Ybb U;L_ 5dyFv@'"3(,(u8eP>o6Xg[Uz2}	B.P3\lv[T]n.8!N5|VPT]<h\T5sKi
rbW&6SBpsyB!g7KGitaP+"3eHB<y0H-H8yEGox16?VO3q3CQ4?#Q|nmYvDWcdU{;G{9:OI)/D1DW2kt}.``ZO9Rf=l0O&p#jsQr-Sbz -hn9X23H|<p\fKqmd}m@z-krY!	>V!jQ#M-Po>3Kcx[Ke.V'>1j42|>qaSr}g-sXg:U;ad*/dGlz>#)ugGN-%|ndA\XxRnXnQdgs>WDIW]	O:04A,| #a=h<{rnsT,fl:GKdq~nDe8Y=_l X[H(=1CR5R%n1^<98./B;H$uekyru
n X-IG?<Wbd+cJnTV+_O_ NPj}!QJ
9NGseGK\KEq![x/cb`B0~Hk&bBUZtJiw'y8?>poBE&p.@>i'kQs*@
oM\Z{mzp0"!d],eM_`S3}"I_Ki:(S!]Wb*}1o,]q_S1(,ENR()7	>2d\_j-B"Q|r1),S<?x2;|Jd{@	]UZ$/cI@D|C}3C@`7$=B_skm8$(7}k4~CYbHEmu'+j{K[B=1oP
A.qi0|'-A6^0z?lC2qYo7=/K=`B&W5O)w1*>.Dn99,q'^;x H'
qEq*`}"	Ou%G'8]>|$IW663~?^Ur(bLDwg'UZ$f	TZJAC4	#2nP{j{p0xqe`Qq-eRi/?m<t>0 iSL|<9_mw,[{!v,DwPAe/fIx`SB,C|(mrKuvj	"P7.Y2zC:-/deq
<uC3Ur+tvEZc-Mo;6	?,6r/nvs
KKUF7^|UCEE7k6j 2osR1+n5X|&~BrN{zg@a-*_=;)q%ARqqk1E9;T&g	"x`b
+7JVV#X[[:2=
a#V#A?ir/Ohu~a:^qWG]#2RK(u`;8}H@^b@+J8`3_96.&_8HB
}$W;jppb!_JCJ8q`/aI,(39zY%8t+Mr xa9sO@Y6]EtYB)1"pk[1G.iNL&s,yY#Fl41@FE#UFMuF 0"Z8<kPSJ~wZZNUP?UpMl}VUAw{0}P7}#F6'evnZAU=xP>jU(YMf	r^FW~_
+Y'$qsVVB(62!i^Otk5A}Me,s=j]Z5CW?N	^CalRn&px.cGvEksOO}^j':UdMK21[,qg\ie.eil":|$.NH#qt6]soi>S1jUe!oF-Ouk
y=P><+,$AdvAE5%bU/81"Vrsi6o{P8y=|5kg	fWv2Zr
~0[zcXp\3D*u-F0TMtf!ue<^5N e-
=&%LElwf}x^4tWoh7}^I?v`O9)77e%D)w^z!&cnvJi^hFc&Sa o`b~*)oyFSEm`]z+BOz<r"B9FX-bE75|i1(vC[hW[&Li
N{zjHT(ClQj{xM'
E{u}jho
aR9J?cD?~P>CHZ>
Y#{'Gn[dhCNVf@.ugF_Li(KiBS \oU@9)]mrP3-l<8CLE/p{=nSY8#.a@-'z$FfFxiM5GtKexCNS9jlf+yvX!P&-Q}t|cSE>/%P^FbxA}7BxRM^l?W]R_`cLO 77 :rPZo&7p	?Gtr6+WG^esHW"$vyJgQg[H&ILYv.I*TH(yIIROjaU(Xs^asLP_R',K<M'oBO18\]<.@4pai|;?ZF$KUxaKJ<G]]?x)MMW=F@'/&;=gUvIk\9l(:Hm^!<P!I@)GLO>!OS:i_d<Emvg6o|"!0Eq:~2;n5N?`}
 NixBSz[,x~*os,^Pg6N+fWstg#Y5=}cQBZaK#0=yhbd~1NUq'uRa=5c	PINCZ#%<5m%ma/\,flbz4JtMd:Kb)+)C3*jD
U	#("|[-2kGT()ia*;I3nlW\&hU@fWt|m&EX<WBQ<UPS#)p*2*i:iS2  }o<A0xna}a|4*%/r&x`KNUN)2HTB8T,!.WJLR&KQNLPJqsstY|Ky<I|6Ao/?|"/T'ibmfQu8HsV6#vb=qfaIR*+ GT}\+taxD&@
HnE^};K]N	~UVH)ND^`|GAQDTW^f+vBdw;BN*"=>P4	ZSl>6.j&)uD-'oatd;@J#n"-Bry.bj<`(G9)~)f'F`CAgx#--JkbCcb6M!\c*)?7kS03[	Bv58#!Z;^->-W:c}KdTZ9++J5U7o,p CXTR:-I>u2-XXm'x5PQ^EE1;Xu(k1?MKKIC+ht0|4CtugCVO2C4)W[rW&."]XaTP^JY6m'As'KLAiBP2O*Yi(Wy_VIS-npOxwjSr&vbq9rtucoyz2c(]itJV/2t+vBFhubw12EDgX	wKTMafItBHbY"dbC_ 4mYG^,hgKR %)n"
Vst':nV=%S=uf9E";FnVw%`/UvL;@{B'ZXc "T53fN|VpeQGV6{7Y>#r4['4MdaU)?LI/E\9)yvs*aBv~!#wfQ-\"a+c*PxY*v),a:R:	`~rs3&o/X 	Z.[:Uqp*0"x0b,!1W\xb]o=k%'G`PMul	uHB#QB',p=!`UY{hhtnxUuk^tBkLZh}LaAJ.S,Bf?S A|!~Z?nev[$k~se0rvgPL7_aWMF~Z=03M]pjN\dSYPhk*3/:^3f	wn:;)CW6E%{uvDN,KtN[4I3k[FglweLp(<*)^tG,;h/%v@Nx3#DHGuAq)-\|cY)R2(e8!"'m^(Iqh#T
hj`_OSozKGq9|]}1&(@X}*I*xyoI$
36osHbtO#;qK0}k!^(fS'"DWva5`$3Z Ho_%-Tu>bYIS]TvNAC=17yu<'Owj@|?W:.bTWY+gwf6>K3H*d	]]WFy\BJvJ&])[jrb\c.mF?;tuT;+h%eU?=:Gj=n?Qv6$P<`uo"hymYwFAUM T.7K~CBrbe}}nUsb|A)/P>u!4P4#J|mf~m4]M@7Opj8(lNC/x73;rW&>}u.2\.9*o(@rp;;j+}\i8*4w]Y(]#vjZpW,PHo/cWou[S>!"+#qYD&+JS2L1m=%/@0gG2aM8KNh|ch	oe7DY$E6]OvDtg
)EjxKl<a"X<yog;GYdp<&.s<VTRPZZ_k9%$5,kt3,	*="9sYlLF5P#a`PPP2;;pMR)/Zzu&X5!8uVnA?]G0[wNMCS]Rz)~*r!rk|1xZ+J0IDN!
F4W*k(\R	1pvC=8nm^fIVRCSH\-0xAj\J2r8CpQb]!(%9]F<y2k{r7zPV$MtwjCJn=:9sy"\M%FQ9:3>G|SmVVLT37&2^
VQcJ,wrYRgE \cF6+?wE"N%$mc1zMrJ1T{N
HB"@kyC!XPl<u&v^[	2,%o6RG `jj#8) :.voQ7jk-*If3PqkTY"(Sa%zhlrPf=CN*LlWw6a8oQ}Gc :P!"0BtqpDDV]].dJq`%q
xrN]~/!:D;Y7
YRG*&81[yJa_MqLYg5b3LZa4-s'5'h1J0BJC]>:_	0zRM/Xd6tI.*k
!vOcw#n)m&bLVdBTGQB;2&l93Ab[5)3Cn0>}PMc$j{?r>n'>c,n R2C^yFAEdZedQ@;;Z,{hk\j%)<V
/T#Fi-^a9F8ido,, fCAULLyf6	[%\G3_c9\1|"/S-^zNBy%2P<^FW3D:GQ9n{@@AW
9S$*<XCwW.8-Y!zq:u:"C#F1G-TDyalJ7(5#+tiS`%?gdiHiEHXPHi\XKN4'~k*aF%y)GTaEAl4O%$
\z)s.&en:gK/@x{=~tD8Bbumqo|,q`C#Gbj,cCn5TY^(tY<_%A&')FSAP7;>yWV#n^/S8/w!0R-fh$q|G0<Jq\6?]`0.K$61jj|znH.f:YR8"S,$KZafl*X{gy/AG@w2y6'9+r6"*~#] 9j|c\{-n!*	)N,fu8[SKkBO#;;Hfl8)	L{F:T7Cz\0,y92>T]\WHe)3R}y(2-{b(lan! ;?)LuU3m@<hz&0~dGI@]P>T67WPmi{
\uaH6^]@$3pOe+]hN!7C_?[9	Yw{P,NGU	d&f=V Tef-5@I}{bIjM6Ig:D^XQr|z+U	;0J{%n:Ax9O}0/!l)d~VB"e<;z~C*&!/r5Xvo;VQwd76:zb@jlm95Oc
|	1y63OrZ"gCps4a'
@$=}NHuyY0%5B~T4|JZktmfMYl.C_bM
1-tm^iR;*YE|_$N5~^B6P(zva/:o/1tb\1@]#+fpbQ:,05n3>?MU43V2T;POS*h*Z5:2#[g#+<?sD:V2ch6gtx.5Pr79zi0)`OR-0u]D&hw<! "WK7qb {b6L5-nyW=5bq9ubi9j,DGh,Lo[S'$gfOMGkim~3*-Iq>9c]0bb2P)^, M{yDy%@tpdv[(VHYB+UlwBe{|ISCW48v)-s.37l/w*L2Nv0jYj5$79g06LIP {ak-\xt.Z;)BRP*][!Q3m8dQ}+.9Yj(d~6v6qM{lF[t)-ekd"5}mv3[9x}iU*\4K:s&o-|}[X1Ro+'f8E5ECRJu7,lL{Y\}LU{WcQTse}"6Va=PSkpE842-1 Gb0dAL`U,iSG9UIkK7`ew:IDh=Bg 
3ct=0k~Ljen6@@}<Ca/("X Oh.!quI:B_k;3nUMuE52pf|=M(P4m@>wwE!!4:w7{MMwh/<yXpd["[VbFo,dMwDJf(D3<!vBlfYEAgT0oVqb{#	;u]
6ge.!eCaiq9We_7YdTdo[yxZM!(r
M,Tlvj]Ftmulz2,&%N'J/v.*Awmzw9g|vm/5XB\CS]ln$nYcut1>cm/I&Y|Xzsp	cm}e_ZG3M\u^=]ModDO=7YY\-tV[>*g|N^!^B`Zb?3y%
'<|%
mH|m$AYkdV#%`=|z1;gDIfqGd#*fK_w`Ac'd'(sFoyP)
Aw0w"#g@6(JP3WdTNksXC>Wb8Ly/O8_mU?*GK7hhrOd)Vjwn^|Fnx3AM\)'M-9#Q>J^2W8S>!w2|b9KXzfqd4MQ1X Fw"tLpul@x.diY9J];Voj*dr{xP3y"6,d{Hayeb!P}R	IAoWD0}a2`Bk	bP<YsT>9vxE&2^Q3R_^}KUA.kA{4E>~whyX>6g]n8kwC"He!:x;;`@ztQzV^OBQ{@rD#Czp!X#8%~A>~?wKB_7izKqr)_qN>W}riu4bK lWtaI1'_I9xg:Bm/v$#5{Jy3w9hV+@|Kw=)%(:NX;>_S>Fl+W`X7sBD`U$Q^:lu>C5$Drc6S&p)6T8GW^*PncVXBGpL2*+ax]%mDhTm8a*.<Ynh23ve6Ay?pTaH$sEn\a[g y^W-fT8s!nIF~	pE*U^IXuS:}<6I4Gg;[m!aWgMZPro}{f*D0)_85c".I,Qz]1/bigpR[N%#N
glvw7#&D/A`60:va[f=@8CzEHbu8#l]>OlEpI+A1NTIg95_C(RHQ6{0JMPd{z}?x^]J0bC&-b8ne%&FI,!GxtZ7:>^^Ue:S`$O&$/,znG&J^z!C:rXAS	Ty},/8/T|
[CgC`{c/%NFJ^TD[Eu#ui*}$|)JndcQnp~-S.@m2Z'bF6FA=E*o"Qh!fuxGk)p5>4}h[c*7_duov+N`2f@s'E9hk~`uJMv\GtJ9J:azc9lx=*tfLEbZ:?6(]Nyz}'N7|	K&#4J-<x!S>kNfjymi]6=Flw]7L V:F57swyKHKSqe=WSKTCX2o@V{$O5iyBZ:moURS-~/|/\xITXp!Bn.Y,BzYB>8I!HF9NgQQARG=M^jt`:!zb[pt[Q#zdw	mc1De	p
7sM7@^GDzj7Y_#.t_vA@4DHb+\t))dbp&L|K`bEwgnR+W*	V%1=tj}MZ27MzBQ7+__(bT\!l<U(=!;JQWSr~8\;$-NMR/lxw^_p1+t`0FD:m*~V0CHrQf[ZIE$!z)Ov|tyI,$x@O(/m[ZRg)oU*\"1D-Op[TV0zo4yVU6QKf5I<ABRSQ#v^J=Xu/\peVgDHYj
(;
2-%=`OscVkWsP,JHm3NAF`<ycg\euZaTY?[3"3J2j:C?wIYF$@8+24_*Mpf43]UKnpc+OJxgs#E5L,tXU32<:ihEF/00olvkIP<7}Tb[c^0mS*F[Xxv$5N7gPBkm|Zy$ |woFq{7j:Yshl;`]R)p*9RXE1*w{;&o	cn%]ZXSM:Mx-S(>bd}aJ*D-[x~2^JigLKW(.U(Dd60dS	|O%Z:PE^XS,Z]&6&^8vV6E<y[U*Y'U>"&k1KEVE2`;CZ?C1%+F=F]>,"Ky%DCczW6|(=DV,Xg wE}.UF>!=z]ae*Wi}D5,dDc;)@,\3c[8r;P7V5FW1f>@S#OWi7R?'z&5IFF;4~SfBo2]+dlYc;i>6Jj)XEOE??LEXk"Wu$+|;mBu\<V"g]A9%a/HYXT-!j~xHb[!66~0Kl-)Z#@}Lt	87>>v3%ImPc|VDpEP,`{?nExfE7 .T`$DZ8nT.hMR!+ym0(dDz!TaY,1'!mG0F6%1//<e?z9]jx3%*yxM(1\VYL<;UqO_CdWPzTs~%zL@EThUp7U"$T;&Emd{,{T0rg'_Xfv;\U4qP*WcxHp k-J}]lLAw'^bht?K}$_9?*m5P8_MA;DEo"	|i$V
Qo+l>Yv4&XO2"7`T']P3eA'o3Wn+Sf6#w?cZT"2r]+)]rRi8:_o_A^")OjAWSs6&
'N*]`S%h?p8_nbca:,0/UfD@l%d8)?}9j31tRav%63.9BTe$DS:	pt>zU-DE9H}$q#$b\{EE>Y^YlAGdra3sXA),!1z:j/O"|/lF2mSF[%_xasPpIc{ri,*R3%(GC2R;?wTx5M/Bn+v4?exo@	y1UQp+=s_}TzojgWI+z=x13*b s@."67E/
H/OX^1G/4l@qm+<4Ym>6$SJcH=:9JVu~3UyDDd.`i$gRh)I@GwK7+uNAWs#VipHrzEVi&X,qD#5./NV$~F>,f&(m}oEN=?0fzQ$nh#Txifd
>[UbvZ4Pr1h5V^o|Pl$rr[Sm[4}w
o5/ULr0@w:dQ!1jxTm
88Kto(vx*|rh.yTOgj"Ax4'MX]Vc+kabS@!@Q{y1<_g61yVkTR,iIz:ivt9fs{7X;qvj'^,nPK4ddL/XBron2	bU%|*Xhz#]5m~yO%4*SkadU \<%9KZum
sn{aI>bN&x
eUSx-+FQ9~yK78W{<T~>6`"i}76mTy1sR*FLf<'.M6c(IcP{o%s$7e3,b/Fj|$S[vFo,{c6h8Wx|`@]Ppx`95!)BNH{N[.Nw&?N.#O|smF*q<j_LPRM8U"=p; Inop# 'nRtb{b3gKz5&/cLEk22Cw9&&:Qg[Wro&rezV:eHzKo?|9RqR8+a,"]qq*bikFf5/-mCZgAg7)d}/D;=
+G-62.lVU1|)iO#5r$! E+9|(>ck	W3a:p1.L#5_T>CpH$Ls;L.UF4)s/3:;=<e#5M;Gu;|xD'kaY9K[/hM!m`'l$0-hwWocO;#[!,fqaiAv$]-/AymDw
YN5$C?VWk?:J2\	
KF5*lmrsO]8lM.I1,AKjkl
6zV'ZBQfh4X3}2ZGB4n.*t1odaQAhFs6,iw;:<`) AMxJK(4:cm>p)u>C//$ctyQV-ffV+g_<x*6@,|rbbF#u`XMckYKr-9QH[3hI"TWHp6<:d3S[wmOK-Djd[$Ivf7h~WLjJZ7`GoMT3hqy/V*~IL<Zp{zY|l(hpiQ4T'LwDlT4z+gdUqyMIU}MWQlU^IgWpj^zhmUa4)x-p$mB7pynn&B%qhm,mMl?V+SeR(5b-?XC0;m#G1K+/ROqs39R8C/*u^m.7H
J-p5YMF|\mUT]2y%A	mW'PO|<D}
[2IxU796^EW%8 IJVq %|vS{%O,40;? Yah\3iGkm?Y4p?k{2rMf'Xs5&lw|waf#NG]%u\'s
_.yF-5(i*	YJ(15Hp\|oOeNd)4Z1MHK*22JO|]40QH)f&b6@"qyb]$3d)"^6\cP:UG&%mpapK/	U3}OMVc"A3@>fagmOD2CdN^"(Oh:n|S^7kmG19v&yd67#w"|.z1M?T
P"C5rWe&|'efk~K0V]5\:S*	Wwm7'_^:l"WdT>e@	"Z&Ta~VJS]JIYFdK3%BT!$/L(yI,ML*]<OaI"U2M[+7"z8]*l?Bs]\m3.aTE#`7J99{MSC)ZXxs$"*"@<RdAp<-LxjpNV(2ZMN!V{}a\	[<%xv8<`"Me"F!$
'qNAKF"Bl|\c}A[-'4cXlZbQQp{XcWi:tJ:1cRg[Z	Msx	&HCS%`(_YPK,NF	2]H)q<jeC&o)C6$>M@m<FC68YaFlGbdI3l{)pxi<<M
?wlAHacqbwY3BIKP@/xD'`ENGqU:w~A'jDlL6LwiNJ}Dtk#n2]}XmtbXAUqJxU:B<o}38=YG.mc+xi;(IDSV4_v>@4KGsCscnCeK_:XDrNb!'JArQn7Z>@DT+bGXf#W0eIw&Ob%GARp~=RCu7sV4@H=8.]Ip,7`	5z[r%Q<(r6^E:Z|.f*E[/>gU#Y!g@Cai#&c3_cQJ4L18*,IXf)>f$~'BI<XW{M7j7-#Yg:px9?uKJCrhKb ^Z~2@@nQ!G-nJo)WB|xe3y1&k]$!LdrZHHZ]O@xe7)`mcg^\pW
i:wigI@Q(;'D(B62VvVow{{`|t=M7ma2G_(|KsqN?RUCz=7ND6hh-m0;/1)pJb|$n<A@bw6snmfbfYJTnDSeP*Ow5+>Tg4ytFqnj$H<	lJW?z")gG~O =R,57LDZU+3'}%U:+	is4,<M!ICnQ2O@zOZ|A>2N0c1>JL@$n$IC
	-mWf>RiuRE+.#2,@2C7=SRhV]~w	T:t(Yq{*JK~FgJ+nSuGpz}ske t9668)36.^m9H2G_^b@k^98Y,[N@8N^W=W,HPIqIDv{NN"ER*eIG=oui<N^%$/.By	M,q*R`||=
\%+p wF<})@K/JS>(h|U.<cl?YYE?sp\0]Qc$-i <'p-1<UVg%0a2F_l&*S#n2_E6ZO~$~lWp.\DeBtp$d3{0:EM\Fr`Zx_BFn-!dIp<l0h^ChN
b7<QlZVE$_3<ybA.lM2PW~<IFimb5!A<Mbw+Q5D"["C?NCXzPteU33/Vn8hYS$?XzbF-[BFJ#5Hw3zCE)Hxn{	L*78 w^(>;9
!k?	%pU8<(!+HkH"H2^F%Q>4Id@27#rA`ef&-#K9Vdo0(,KPCSNsH_AF`D*uj/dTpruX }0pcG.jTVe1jvRRLL=s!p\;"}NL	Zv#x^{&FuL^0:%2PD$4w41uMlN*]<"/lw["N;8*X'1,{F
l$AfDLda>P	2}8mmIZrS
>mdH6_}<sb.t9bO@/)t,-T60 7AZ."j8~kt=J#B{TP1vLIw9wNx ?v.ApFdeu$#!pA))%lH'/7%W*`V'0[b	L,\|A)#.mM,Fsy!5uZT.t6YA(Age&+4'\k>snyY@$\Y_ Q>QDQ6>]85H88Ir+{1|&q3#Emh7M0\}BD$T#xK)w\D1md7BbbNG,wT&C)*g/)Hj*.tD%Fp*xb^5Hw
.Ih2AP+-nV
+.	J!e{W+@7?w!N'0zU`,@'<`[mHKDq`otTJ(44	^Dp$M2=qtTuv#A9^<4)`
(8ecY2ZFUmWZpzFvqj;U`d1c+Kc	"6.8f(93]`AZF+uH0$<P|IvH`OTM.k%Q\Znc~RG-`MkY}[yU+]N&c6"x7F2x^+`+H8O<lb*:FvI?e[Zv0hAQ{|xv~2("0A[zrhZ]7XDFq
2Bpv'\-t}tRIW\\C7,O\jwYAXB'Cn@Jd>L~iUCy<SLA#z&
=lf#PhI4_s,|]{:AXWAn2xay|6{O0QdXt'}gWHD$7W8-XY0`z(z	q7Cn7&w1z6x\FdH(IN;Bojbs-v.Q7n4n
)mE'`bfo4>^@uE_59hbx3cui1=u=J-HlrYgm2K5x!R
Y\T5XuAPzIg:!.V%EqHC'2p7|HmuzbZGfXO
PC^m>HRv7O_({B4JhuizyiaS-T-5x~WeqC7bOa{cYiQ0WEqMl71 GWytdbw\cUH
{xdaw1Gl.Qb
Gio[V'Z5/F2gn_ciUC&*NA)$x"r+<V1H5.0F[q:5OXckg"Yadqx8c{L|c:HuTO&`n?sM,[1GXy!#]_&mV<kk}YX
lB/8scv@(xicaM5!Z)cAj*liF"1U2p!YR9/+2
5UZxjD@NsMNP)IRw$xh9L_B.L|~fUC\VIZp@$^GR_P2$9Fn:^CfI|.;~`4V>%BiCyUXi),-#2%HD{&q-o0OrkF"3J:vLd&	r`)CH&_v Q%PD[~]^3fHq}#('."!n>CIn?B!2	2ns\;ot,unl45O[cUp0:"v DiW!ELit:S^Tw_{08nvJpGp@!hXX@5> Trh>#!BmtJu.C6rbRfw0A|rjuvds7yq8W| w)f>1EZ]kFGfd?RU~.8u[)E3oX 5W`9Xbw,Ho"s&;yA+cP%088#AcZg i,md5 NL88P}=vwe3Gd]:G/{y"t8}K[_Z_(E2!|anE2)p'I0k3qb%amDl3jn-%9x{Qav)`du5EZkz%%htfbF\Z^9HO\XJ\8-,G~Xay!e)~gZ)
_s]jFxf	<9PkOd2FOe="TbNTq&BGES8}NQVs(gxMJNcR1@B#{gx/+#ZHB<(.bb8]WAj3d<BmP~^"V	![G^Y
k@{jxe6a IV@p?E'u`M&l %?;IOJ=/R"{?j7K%1MA<<*dL,}]S"%Y;#,[xw	De*%E|r8uG^^Ly^{)l+/2U*33Ijbpmnw|XGYnGW/9Wwx*},y[RgS.tOYH_\I*'<v0HInWU*a`PibUNlj?9Cwc)rzS9)2Kd#\xh8<]p`4?Gt;w|y./Oa&fo$)VI6p:Uj3[)$N)zXIoy<.Z$07#o!O^'=]j&H|ltB;&5Iegt,C"b|k'6
GsJ:1",Q^R,DXPk^ya./^NxwjbcbVR+y6rf'	Vpgg? [w%^~ZAkhw7O1:
Ffb"Y4M#EY4yQ*89yxXj!WvYR3+.6AyCItMgm3@Wl)@D2W[|1kG;Q_$.o{\$DMj^Oipj^GNTlD0o%P>[V7+ ,G)ko=28*UmF:0Y96i5n#@)h"n.`]!nizUrErmFsYi/5O?QkEKy1X{tIayV`d[<*2vLy8#pOUJuaJ/0xp/7?o5H.y]xO{79D',epS9EXi2KJ2$k6<)]NT^v,~vf#5zO7OFV2'z4slKHln6h">32:5CYl>|p)J}*	7C'<-t5
tlC2~g.Wvs!x:g1`w7@yojOwpQGw,(L
7UPzWTK>~WrWVR#d^uJLSLy+2:>x{}n{x#+?]S<GE6/8%W@[1~)fm
J_m"<jI%R_qE'u,>tOGH	c048<qj&*\`;oo #incN{VW%Vd/0x8>l/-lw`8'.#^t}{66gy4!V w:{ 
}Y:56}Sg.`H;f^r@d/P'b~F(P	6q0b*pDnjv+@0N%IXq/;o2[g#u4vk}%`SyW
a{on0NKSVJupln1kqA%|u)+GGIP9%0U^V5SR$:nl7H qW0rVJHGK}(gPe#v,JIE.O)cIWj]l,OH_Q*7az8:lxK]>	Z9_$.Quznu%t1]4P,`rK\OZjpHQ.tuF:)K\a=+t$^o{k |1
Sm}b.VnsVDCho/(+:Qh?V#WG['G'x;x:W2T?YS;~n6&!(ypVUy|_e5vV>XK65%<aoM,\}%?u3>3px'"+>8m%A^it zy
FR=E;n^<F@OJhD-;{j:{,1dO->xzt,9[Y<|{L8v^%TCJt>W4X<|fCYz<U99c_g)8-n%DWXXkzC"RN/V1Nlc8qOYjZJ}2tka&;A{!ON5V+p-oU=TY_P#$J`i|fa8P#ZL"WP"C`CH*|'M8[ 7G7-	^IKp!:u%8>_UtJF!~Gs)Ll.*En,7QDR]a)/=~uC()GjR1xMmYlP:LHv'$+8M'-`pquBC  1.}%,|w#}=ciX&Ir7Pg%|o]k<_HJ	*YCW+a"-W&oH;wK1MU]i'	EF5k}kw-^e@B
&3ma@W|yR\rhb1{yXsL[`K@At4r&-t;VkJ5dY>+a_2bJG=s.p0w#[ib(ukj+I0&4Y$WR(wDzX#u58DZW|Dql&=1) vk?U*@L85M6JWD}94=)2t\XsVsB=Bdz{dd2Lv}>4{\|Z*(ccf>y{N)t@/E{Xb1 uvlYv+D`BGK*;Z,Br]n/\Rfk6 Rc?p)(K()^"%dz[!jdckU;"u.v3~_-*
ioE,M.DKjZtwRW>co7te$nFDKz.+4Mt316gkLO<J$;|!W-F8$GVS/YDR]30_5iU7>a3)I};	K"dBgPK9f!~f{n0K8t=r$R%"-Om/=O4\(a1*+Vh0C}Xx\OVCU6g]G{;l;0KvBQauc$Aym(z.OJZ#5xR+<|dt(cT9AIYztaGUM!d70})vaT~7.vi5}+\x**dG
R_2LPv{iG	z7S0	P`S,)$MQ?1xYRDD/iC){?+N{R_pN$1{vQK~B;@g)!7NpR9_Ex~I>u#<UW=RMX9zVh	~s|]JM91L/Ts?b`AjvH%#5

1CfJVo)L_<%$*kxF@dnq\.$dJ}aB=k`f7nR&w,)S;nwuUHywh<< w4vNT2j.b7gq?/JfC39Eegvu*NY^D5"?c5p:al[`,w_o\CEZ@JyDy~8~IsS[~4fvG}^'"&	r%sj{N27Z,o:O/dl=Gr):^J@1(m@S@s,	dY^T{P%u_0JNuy6Y!L?,Xe'MtWt@[JEzU<AVc->{BDBT~FZ qn}S8?BM}}*Aa0<D]o^P`S&No
p[&HKsP04C1&*ve8$,EY^),X@ls%kxn
iJa>odc</CE?3 -&Mt>>}-{C\A+u}f2K
Sg2hOtPOi2HOr=<]L+YFu+`1X.,ErK$rKY	ZhRF0|A];:Y#RCFN@c|8?xrRF&T"'*s</ezz^ii+1Ho
Y[RS	fgMm_@bi`
2BF)(erP=5hY[/~"2 m8_RwADJK<iEQoNBN8VjRHe|Ye$hm9!<1%<BIt=	Sd\DRC6,q&V&=.+n*t8):0y`qGFJ}B$qBWVrE3q;{(O`D'Y` fZ/d&26:XQzO@flY $E&u#=)WPv,e:8"+.]wfYPE;q/!	=4A,S_.?qd344O7*H%Z/.cp9t)&i8da~a8x$3P	Me|w290LS=	dRE#K+7m(\=#0L?E nu91E^Q{\3NnR)KXTzW$v=F%UJ!QV`B!eN/=Lw(f@()tt,cx)[gKv_R[\B^Pdw+U,pe"b#>f9`E~")-$Pdn`X>KQz "n3Hp!y@0?@?~Pi.,0!W"T~$[VM+4Jk[5d0+7@q;@k2-6YN`d_9xzgGS~\vEu+i,mMFY=6\BtY3EP!i'[H+p_d&,m['XXY0b^Va38neoFS|(),w-f?X,ES|>avC,.QryH<c$&Yhu3#/=IlJ4>Z/CDRJ}B-Oy]i?7l=Yk6P]}W$.U<|sY*''6T;>B570M).TS	?t8!&El5ow?
#(?D+Y*P#g[5MZv,B'G8|?]MY!r=aCu7g,wo8*[_X#G/]js<M'^vRjosx4@V>z`Sj'NHXRA,:&-`m;?7jt%p^||NaK%5w3dmrVuqc]N<'3lDb`zy0#o8XO$#b#|ynr Q`RGUxS0,7L_LgbNT9Hh~#mvq&)QW_QSg[A@mxzfFpq8F4'>-a4_YG=y*]'pB(4t7L>?3X+HCDE*K>.q}AHZL;;}A*R,R	VYfoPOmd6`nSm}Yas<|YbjfhH8ripx4/N$c(!5Q/ X~nPj/9bsVd?bfgj`C`V"!A;#
3o:2*ss>^-?iPr6R.$dPK6@, 6+NR6\^= T%p	<J{V0JUg{~5<gB`!REZh%>SR.+Ty$WZs\K.[HE3 kyKxw\y%6O|uqWZz\4nv2.(K=&?n2C)kCMeF9bTinPu=UCDj5bq11
^35g0-7?N+%2OeL)Ml0FU*4 W)$v7`[-n(L<WbP%[\x</zNGx9p?jA:E4N.Y>DY&_fUJ0r2=<@a 4|'_kvmxowDPACoc FU	V1Y#.?`5|@5}=0.O?dP5<U5Ykqx~^_C6JL%N =2"t{lDo=m""+d*{+5|`Q&-eop'Z}@uD89Q9(	obIN`C%!]FKaiI^1KUn7B)WuDCYDu^[=!whExp&DGb#oXyH}Hx{fp::W6kM~(= ivk~850LPG+}xmP|>A~pjv;`HZ]f5&	M).s[z%Pz0@J3.@~:6L/;p>B[|CtwsQcQG8uqjy	5($<W?|isINTq9+-%AGEtKHKI"bxjntTe)~ox{ UD=s%x:y*'q):8*j#>c%p9K2f5g`HO0four[++_T/_GQ/Z}9,qMOc:P,{HvOPE]!Mb0PZ~=[M7f)V3fLC.ANbo4=VJf{:jg0QRz'/-{ql/2=(L&$)}\!TS@f<MY>F U@d%JLXbm0!W+.{t0u>6tlw
?]HMBTF{va'-+Zt]3KPIX^I[5?:g.B2rh%vF "!,0gK#Z#$~Gw&|)^I--``<Y@oyzO	FV[AmbA,eql.h|K*k=AU`OX;dq@-8WKc]y;;9\7vvwez5~h&>jm@ON
dk]$:{D6aF*o0)5kvN9Q'8>jlevvCzt9Uujr5rk&`9u2C(gRi%#rEEfB VfI95q{2C3U\LApL@kf36^F=M&UhihXdO]9dM
AR N/4CRSYpU1rq*0af8rCs%9#}K9{l65dX?(!cm7,6XoML;vdye{O&a5Af@*'zz]%V2}1z*[`!@qC?O5]&Rb:Wo!?X&>M0_<>9@cy1"%Tw]T:T9Px]8l1%(
'R3^5A4XU{6(l?_m{^'~
>dZ
	s7j@i[m1gCR0I)Xh47R(T[Pn@xm94:/z(W<ug8d(@/Ae!@O$]y4Vt>_1y01.G;&rEo[ (GP`Lqu-:t7dy#e7W<-T8J3Feq'C	!Wuem.X:5:Gf0C*O?<M<q)""QRP=c1(ie3&V-7
%[t)'(;htx6J-eHk:j;Tx\~e95DhJwkB:jIgR"kcFy
ggA.~O(@.f"s>+$j9EU"j|Llw+36<hP8]K[E}f$Ii+lY=K<,Vx*`*{\``@xkLQx)pfwx	BVym*#2O+4=[d=V0A0rR0dAKBm.5~#jR`d[.\|F(LQvA`KB!nG(}(FyF^it%{Su:V6wXEV7UE_<|-<83@H9(P`CyV)/E0=(H6n
eKpOFq6Mfl`dI!rr"f-a6P``<bkq_YeiMuArl8k*l]vw'z^0gp8rpkoV?O&-0%Us-8Q4dr&w8ClySFlTA#HPeMN
:{3SGN55s;1]f.+1nXLWJ7T"Oz)H8\X|5AOpN&K;tx.H9;.-4>G|0#}sm\tM-}^Jm*aS50poi7H!Yk@d#lkU%oGwA?I0EB/A8C]FDq!,?w3.v<^5/w1]_r{D^3:c^i!DKTZE;\'l*S,-{E\|6Tw|laJ81F^ENoPI:A/G}7*k1ngi&g>N_y653{IySo^+|."Ce.RvMQGJO>WJuVxa)*SzR+4[{CKV!t(X$_h?bVhBoUy)(L X]n9RUaDz_.KV	9EVaoP+y_N<l7r2ywV7,w\$wWx0:u8F.6)RH])69GWuAcYoUosq}bl<8px\mmn~g]^1G$66J ve^KUTTq[M1$Bkf6AD.Rm3b|.k6AJNLt)j~${!)4gcYtI`9QqXvz,/EY%Bc>6CKc.	#"]5EsC6I~]Xzo`S7+gvk/2T@b1^.y-cCMCKY@I<3{11^B{<0=~N9,=W5]FT=Q~}ECY9Ri	HMDEt>`JGE/Entap}"|vVl~[2{JJ$%,Z4<^R37Zo;1<5P.M4>'q/M9h9j*XmIyN3fx'O2nK|	dE/;0&'
vWu7j9Ag|w/\$!yr:&la7"'(>f`y>bPi#RM/FZma%L-,vCLld.Fbv'Xul,)JQ=e+'f|i1JXU:O@i4HQAu_(1Ok}O5,~#!0R'+-=L)x#UCR+!;hZMP=B`vQ:Dhv+}cw o.|m;L<mJc)tW	JZtK/
d!OZg> HFCdjA9T6I<F(\g9iG5}BGY&e2`Gxh!'.Dp}\v`[5?B,ym(,?Q4;-kU5oXl7
Z$h]@_.CUSub<ep}pLRGD>x	3yEa4&,"I"&YWVX&?)Dsl+{6U~pC
,.fa5)@BugULR	~/oEqD(dm1TwUcE
t]>h.H}h*s69 b=26>5d4]Bn|rfp.xG{#3+Pc9Hcl2OZ}d1f)[1g[/T`N#+9`.ecrc.(s3;|%>2BF97m0TVQgVcl-z@BF`H52'B\VyMW/4%t/_8|8	xsj/4zZosWTbnRfV,$?G;D5>IT3nX!H>ahrx_'Pk4}s!(Kf"Tb}dQ}E&f`QhUpK$co}ZnTR/bnwaK8b}GM-\3!DTA{bv b_a^R!!:s`o])&N0BE(L>u:Rc-5dx~S&"evL@g^kKYKX:~)O%2ar-bjf3>T X)]8 ,TI4Sc}W1i	#H[KA09,>xn"SX9eN%|?@9"U)SGdrqZO{0=^3Ui0b@>nTFm:i9x[YXBDq5I:xtx7oht+q,Y!w^BTUKPg],vizRGQsOC;d]$p"`^m*/V_2	f;?C.!_{j4Di(J;0?v8~K5WFVeo&FCoflhf93Z%[oHj1;r<	v0r"8Fp]I
X;h,d4&[23(1#>&kr&Q"`VY4 $a,|.OZv)rhh_UV:@	(gC2]Kc:R=m5.)k7.h:hFWC/O`
tWA)&%I.mzG
'c%w%PUhlJ^rjqin+M@* ?mZw,unXH~*d:TGBj5?UTcZHUJZE2N<v2OMbQWri'[Nu-/%(1+l%Vr|$*}[
9q;mdjq5=Sqpq7Qbvp^J`+bN#.w8(_&"T|-Z0`$C0VW]r;njHyc`3!BM!ip:eNQ6|C3y4rjB?b\gY?iTDj_DWB=4`~<#5D}IQ[<W[yVY-3_	^*??1lDS~[t@l 6g(=h;g4+D}-1?CDGl6q7as0yl&.MQ,2ca}w0wJ?-UUOZebPXxQpz=y_hz6O(jI#;{Rm1~10nwz|>bH i[fi,rw~meC+n1u]Sc_ovEn,x]T~6,qv8O,RY)Tw!)[V%r)A_/vLVS4#szvky	GDZfEIJ=7?Rw8-1i+R}\4&o^wQ{~UVGtF"Jt89e[8:hcL}9!FIV*D6}<FC.wL"_I$[|t<p=6#7NpQ`\(\K~-a7B.+Yx	6&6hI
."Ak/5mfSN(Oo|a/]>v0SbZogGiIZd<2OuBh=BgixFE^2$-DT*S=m~7'6OdZ?.^q_XDLky.
^UQmeM6ig*XPYK8oxf8QD,9,{B!:l"$IbLx&cn8&j'-&2@5#$p!L,1^Jpd|>QL2),}q;z-<)`t.BKR{XJ,Tz\0P _oD+1ID{Lf6Zq61Te0)tzX~N0'w]m_ks`B3O9O:Fa" S79[xv(?4E<Ce'QPgAx.=Wp~yKAA5yf}v6;2e`MLpUl
{ZIdHnI(LxDSd28XJd<CbLKn(%)>05@O%d|(tD`8CZl0
I[7	{b7&?6>Q20BV%uj"D$El;tNtmm{_].p749-IJQjs;NL/ k5rfY'
mc`ASD*aYVLCuB>DWQ>58hsTgf$|+FO@tas#+=Z'YVl4p+V@NHtT*/!Lu=[8ktBEA1wmth0sUx0:Ya##XRz}
U$U(,+}\AaCRHRKrG%1m!2]TC6}/$W 48_KncKNGUSuitxC0CaMoNw
~!8"y@89	;BG>xeto-60]uSR./:KO-Ub4G5/<OuH,k$AP~%%N2$1w$JNnq,8myvQ['&o+0-Ty1pu#{[nZv/P5_E55J-PX	Zp?#FlH0yT`G4[{mJPJ^\]/]R"8,Dojb#7fEoRs9m%v`_L{FPQ]"NiT&mHuUK*r'.cfJ"Kv.p9r~'LvCsshh#HH0L|7[WWbYtni.F9iIQ,t{3X5,,}16E[lO0HCRU#$OcePo4RoBjO
cS>TQ5Qs%Ph|,MP/-%9Zom\e&|<vy)N&243-^8Td"9mM,ma?U>\yJOUK.`Uzrc/,?zBF|b;@I;qj
`Bc8Y
Ht/4A>C2 \**6j]Fa<Z;BN7hZ03/GoQj!	"!CEb.uL!lW#D=#2m+OI(F%A?r0R+Nik4'hlu2;%5gX&>`Pb-9<x`\73Y9<|,aq$dCWp2){n[r4TPS~DeG#w
8#wF2zW3#	A=ihF
Wcr?;~}=m^'7ktWk5n:-()yJ&#v5]	^6_!	FtIF;oSXr@q,C/MzZHvSu@o=TY_'/$tT2eC]_KK_S58K"f`]#cp9[M#rX [.s[{7v`/3v} CRRj_v:"xXRNfd=n.oJ1kA=
"I6hJ|d+(LIcBQNJe|LE>o	9'V\;ES0A8,/G.{gXl[M<TcLumQ_9NJ\8WoNBrG!4BeEgF>-tn^QB)3)Y&c;7M8uQ_S#X1!7J!(v3@^g</f#-Jgj{}ku*Hi/zbem')E=*Y)F&?6c,xkx&cdM\U:,<bHn>^sGg{2iU[~Cq"Ly$;9/^(O}|zG]|$CA~)c=ch1CA[I1v7e#oq.:`lIRVcK5A=>+uOzh|XmE>m2Q{_emPe_8dKZ1#<%'?mu=S\X({<	:LlPue]kMC^8~(kLqYYYz$71xOAHO0T*OU(Y<-Z;Y{qY=r>3|yN$gx"AN^B!@n/-]k_'#'s1B$:pg/03.,q&-K::X`f$){~STA{=_im|=>SO:dEga_-1^	}!3SN$:O~kM#4O1jp`[`@~.IQMaKn%tLkJL[}v,EVN#DH79E81Q%Zw$DKK(J'kRWivaKG}^v!njR'0J.v{xtc/9a%b=Ht 4Qv%7jeB"TV$82eRBIX5`b8zU}+Od5^S*:sO.ae#S'-fF-|Q	Pn@:W~4g8!I8qCyOKZp"Wb;Z4h&>bJf06e|%Y?la;9"14GP/,:G6!iJYRTJffSX`i/E?oj5NI"H%>qaG}1h.B'"-t'c.w_ss,ln>rPL 	-x#!L=_Mr	dDr%e&6>h}[V!GHW2wMj%Ta[cTL$7T]ZP4VcQulj1iNOBD1h=tl[2SDRL(E"h<5qca4S,?ht4}3[*-;7;'/"c4NMq_bj7F)s]y?I@TNH9aZ[(4:{>dv>]'Sw$1`]Y{MD82X0AhOE}Uw	/!A5)'C1Qlx{jF8l#8SquLM4O_D5^~uE}W09D|\	Aj(uqFaV-M"c!$+s<hHKs?ZYCMoCtd$2,2$qfu'7K?(^32GaU2Ue%CCp7Xji|" f.FNcP}UW:a.)CFAc9SX&$m#SqQcqWsf%(_d"b``&|8)Uf}gS#yRa2iu6K9|E:jy(d,D/A.Ql@F5d|^KMr#O/A|tYcDF$SHBTF$xOkrr=]n:$Kb6``w)0\Mf;l'+hE2m.:P=z^DD8qWF&t'E}2I6,JyKJnoxOY)Ql;v.oS{:i^!L+y[lGa73IYx}M<bXCL'<td3orZ?/S]#H `=8u|[89[\eT3qV<Mx
P/Ip!<Cy6J@vE?:$z@rFHTOGl]ts`wYRdF^.ALRg&b}+nRc9	Yv^*JF/dW?,S=9>LtPEy2(XVx?jtJ}`W_c	N8[wc!#x2zz~l;vV"$2
Ijhr<HvwEcR|)|&<;)C+Q5,MbkZa`8X=
3|,MzxwQ-1-bYqHnO*q*,.;Ne9"QWPyN.^e71Wyki/?ZnF2ne)s"&Uh\y>"HkXT)8fqO&Up);6&0|y)*[$XaS6;IpY7YA!bB/0$dP6%g>;)|es,&ei>p>uc7}p(XD-Y-('d"dtL\P.nb7sO5{%Pr4Y#9hEx+X-naM>"x
?4!AN4fqw[*8k\wt:(UBMkW+3sko|dA3/L6*h	%K;	jGj3S~oGw?)F=KM5TGr
Lr~@6BU+3:x(FiXV]#'<OJDI_Ap oP	Y'-tO6S}:|L!(#D@E3h;BLsR{FF%PvKj$@"d-AKhd#VG]Z8qZOJK,gC<:/Hh3AAxZvE\
n)?.!z5nm,MKa/]3g<7X18lhz.fS `^\+tPhA ncwibIKW:NOyUwUacJcgpQ{(fm+j4)lVzf3'V1an-7Q{p~2Ls(;tU*]'_KD 7v[$>=WKJ}5>4EVijBG61_uwlIg9%p4oWW4IGxdo4MESqE<Dh!@,&mIkw3v~fdeESUK5p+yeR2YxUnM3q6G3) -.Aa(]gwG<Yd;$@+krswVF\\>WWX}:^
,.FcTDYjcZN`"Tmzm8zPiv zaR*itaTe00&8#F<4c:l"UvuS#$Q
H:K>(L*`4 }G+;asK
+]jOwK1d{q1edB CV`=+?{Hj%V:,?E564-kdFD+4?;w\tfJG)%f9Y?KcnblGQ$d/sxMW9v"Wj:}87bY+SMY]/g3Gu*Vh+stuJ=l$mxS=3q-,ZX_C9*vdJ}KjDvi"9!N3AX8T?rdPkTVHo V&0oj5&q{1]%i8iB~LbAP'l#U<5w&
DR"a[V6|Q|Jb:GcD9`w!w&cu jw6(CJc#ibyUcx{K@/xxf5t9?sdjDpv"a]`9r[aLm-oFdCd^rH2I\rhdkl{y/9Qz-syuV	:s@Ib-#;Q%6dYjdbJ*/ND.3	(T<!U/cpvl-"n2>8G`Cwsvch^zL?\bjvRppr}uE z I'k>&=WKe@$+lBb"IEp+Jg	>Sh*M6lwec~SF?5!^SH$;31ajf8#yS.~u{gSi!QC%QF)vHMo$4}L/Pnr&^n`.k"<:L Ve^[/ntV3I'['a`?TVES_]S9	W'GxP=$-/`(1-Rb)f6HBE{)XNrU5!E}*\JIY:9w1#njy')
a)N-#&Kq]aHzaP/B8bf3P58e.mN{BBX?hJ40G.x}/n@YMp 4~Mrs}g_tH+l#DWEi8tjqARo])^
>.{}B|jD|Bs/Lh&9yAvofk@AMaNsExd_MdZ1KAXmdi
/5	#2kQpTMwH/VTCkEX-zF}]%C9.Z8ab(C1/06tbHCT3]0Djz1ojf~uq=I)UxEwcUv
:B{[]lxvSK`O|X.PC64N$mj&wh94/'C3[Qas9n*:sf6@I-U;yQ03E_2\]D:mM7>=6ZfcaPnSDh.O` {?SG4|k*ANXze^N_NgIcp}/!/E/$d3$7@KpA(Xqych&"`4t,(Ufw<q!A46
]VgHPpCD3DTP5=mjj&LtV'S#pBfP\-`B;BbQ`&&2#t`/FdZgPqW+	]6i|+,z?s2m/bW)-jR8emw{~?OOz-la6vM_:(St+>hN-.X3fbXp4CL@Qn U{S$x>nj5HpNUgDI,)E9J'mt|J6UFZ5?$+;7I]DU5^Mx>G#@NA`^3kk.ZCcc :'<[C5lntgmI]?O/;<@7+BIB"-{>mh<V$Fc93|We4|jE;9ISd{mK
c*!9We g^AC@_<ZgN\WEq1s&dKku(/v+cU_7,1xe[B]FqanB'hYEvL6z0jA$(;S%u(}24w|.K6kRqnz5^g9 %OT;O/uTbT	N#^F%1oK?^_H\}YFml :Uh4]%*[Sn4qP! TFeKpkwkD9uNNyM:	j,@4Wr"=Y*tV[{Df[7q\IPtXl[$#A^;TsB<OY:xvf)xnpP >)+dpTJh_,5dW/ffrvIol\2lG:n?!G]<Ius(W%C/zVyMep,uIFX25k| +4FJ$uct;Jcc3U~fM6U)HWm*{LL;.r;FBny_iJd0nxWRm@<dM;X4ZJzead+@_A];Et1GqWjz>3s%LO%rfqw<iy-r6cJ~|sqi!4v"@0$f,%z!,*K6w./'EhF,8/wU*	Rc0!(OBsLra/Oyw;*- =,[@AX[Kb0B.Ur("P2^&6*lf|4uE`F1'rRPk@G2&,g.X Ujl:y[("=d:pNK t1Z*e;6zITDGByCR,\+n=%8m(kG7ZTL_F&)WE#*so,sV$W?Rx8\Dr%1SgMV8X{*x>!VhL-	(K*]X*V#2RMK]lVOi,d+N81j)g7&z#O\zW^HUxMk2| rB
<5lm0,c;5-{NdeTd09fWc?n(zpFT+[`Ye	fi9TzH	/<;g:5q|9vG71-1.\G+bfCJm9RkO1zI}c#6(S0og<m)p@%e7o6xPRF2/!DzH/k^ymJ~{c{Y<,?IC=/=:|7bR1\}6Lyyb	!Y1=I.:f0N*<j9	I[9Kf1R2OgC_n2(0@I@t-[X+^:*=-wm*;a)W&Ts*&&,kBe"$eMDH;e[f.0iw(rwkdj~I&p&2"#=,=)DS9x<I4MJ3Ol+dW"+u["pwwasV3CRQu	v&]PEaS#(`WSEz\U9*qimvb+M!p>HWoIJ1cn2?q35:&[!#0w%LT=[}Wt'>>h!|nRM_ln;(]Wu*b1t]ks{;*q<	N=;g)S,"yHN/Mz_YTTdeQbZEw)nQG}+DgmXmH%zN#]N"1*N4X<BX2JSyN9*!qjAN[h@wOSEZ9K]Cj7ddNM=?3YHsuI5~aA}H9K-#GEyX/VKiC"2*m8Mi7VH6(Hwa\LUkn(uZjI}V77x"`6,2lx!m>{u++i(~ ~HL,XP*j9nAl#Hd9VUC"<4z';p=WX6}1yFhF&7bHA;9~+O#r#?_9r_["W+U?0U<(jvARzo!LN	)K+JY:kOl,[	N>;3A(?2H{Sl!dGlI>B%VG,+$N[GOoCp\2"BSx#SY5,Q)qmW/Jg%f9'o+Yra{U!QZ?94[pT}"fb6+E33ahRz9(Ztt6mGQ1Fc)]LZpdkf%sY9m=)WTm5U6y<z,sAxp)B *]$X,38c"|nl<:MfmUpf{cd/JmiFe"8/NP-B(8@99bC=YP~bDh'w"`#l'T;wxh<"Z3!n^jSegW$e10I/>stU&)`KZ1p(RkNQ`+LENzn'=WkWtBQ}k;gfV>\En*YQ9xd&F\Imr~!0W=9=3c<db3Xbypfz%FEFC|~Qb|v5JvZL]Q#",^c-5of1+pnXb}X +[	%2Muho,I7y 	DgR$FO[3_k@ew^C{kM$FJAd,]{klJGFrY)<b/R\>MmF/_9pTmNCA)'XQy>h |D:k
P?MgWUl-%If#]-sx2IW9pF}L -;M,Y_Mlh?Pt)EWfCTa`iv38^_?4EZgVs[mKGY0nxW3r QaP?0ml%`kbh=<eFoM4~j>#Yki%W31:6X	#Exq8uc/D62f9.V55g	M.6;t]Ph;w":_3uSMK#rLr7b3RoI<`Oie0N]ob%S#"d#nE=o~#xyqG/B-y_;fC!2ZFtL.zRhk/y?ta}EC/@Lj;c&]"0f[nJyQ:}uXJ<^!r^$J_c^H;+;WF!T.R+	~[XVl,o\f<C,jFs{QW81O1KY{?i"xp~^<i	"1v<M[Z'Jdh>tc)Opn'L469c\<y.AZCz=kV/v _.fp^1qIBFB W#+o)M`(iTEq>}AAC=MWf80pkBG)=+5 $DPY3hg/TvkIH^25V5c)Wx*Xuw2O?V42A"*]uP>z^)g$g\u4OGOduLj`F|ZlwGe+4vDVcCm?Jp~1\e`~[I/z.8.;/a61Zj}CgsvZ	k910B_oMT5+tv4kIv^Xc4[xZ[@xH?LI|KNHf9]? 3|#l||B7eOhDiB
r<Jf^
e#g,;9mSJ/WqF%b]gl&mh@954D.tb["|Fzj20Qv5J^m|zq\Gr,,n|;Kxi
'zoB4
-Q~oZ&e`/SDs!9G9h'LP7]1_FOSOAz8ttQ9O6R1 G'z7MXR,t8<"A-hhER P&wq=[~@wz 6";#+k#}V_	i+K!*$j837OiqG,SI{fbkigX:W	W(&(|ShztjZgc@[pd\bCco+7	hUrHn!$b;fdF8B1{zk!v$O%+$R_oq@FJ9'<Eee	m7ZKQ9Znjg^!uatr$/BQH<}RDmWG{*P*}:wH8_Ns)vPnZ\oY>[,m`M\rOt[vk7k*o0!b.KqRPow_+c,B	?Aqegr!jJ*'Iy|.e'L)  &evp?Vr"
F/FAnXMn=H~OkYJ1l9;@{y}xu=f1*yV*SxA$:&0ZkcLT/(^KI+
N`<]D-Rr9^h/2wj*^:TIKEl#6Rr}+*;oA#66>9Vs8wO ?X!Mup5iSTe86Ou2#5%cz6Frq/wW~1Z#>4t-%Ow^wVpJ:7TA)}hQM<}R&Caj_NzkQ~bb+wO%sR8b2R3oz[;,#>G!TBby;bT 3g@pO?Jc8Y<mqpq8=9{q;OGn83	/ID*gXkNzqq&%3iIImgBZ}p,2d'sZ24'Z*wQnD8X]UH]sCg(.t9XP]0iW`RB28g"i!)U7OrA7$p!jE~x|R&2$z]O(pS{3!xx^Z
'0A:wb$&.bpkU?pbU;bMMVZ$IRB<5b!a]m{Xb!)=NA>(ve,H>(D@oC	LdLU	&][{muu$#SVtvJnQu!5+zGu!ga(2-Q3G8bG<|-zj"xMr0(8Nj/wFfEY7H@nE]#f^nPF,b7#&"^h*lvDEU/RK2E%d#	96T"CR[`{5af/%-~8Cu 1j,e5sq,I%uCeQ1UAR+f.Al/>gSGqS4<D:<
@f a'W+Nz-os`K,"a>`|rG=uz\h<L<hg((jIS%X2$R)r	u\l+XzpRI4Fu:.06_s8g"%aIgS4LI)aDYSuo2#K#(*DM+%c2
5JPrZ:	,{aYC=*@ xs){y,n#<gC98wU@[[.pr(p%uSR5'#6Y?_Y18SMy[c6&zaF}{U/&maX`CGx8g\6	L4;S;)gL#1+FU(R/Zk6m6(A7Pu-UL;(f2zVE*T8w=g=;4oX22hO'a@cd3ZG}?JVnpB@V&>IBW6HS'nR9r_ZIXB/:(q*XfN>Hziz$xpN8Ik|JA1>	=pTUr.pL9n
IkKRRFDvPwO8uyj8OcF-^?T`uuyrjqu@%Ip%i2q>
j]#`0/lbO=G.dxJP>8Az.<{iH[qLYcn'!+Z@Vya;J@]v-dBrj0=r }*
!r=k,x}\kXs	<yEQ>?FWTn7;q}$D%2vD8`+ FGM(EQH|/dSwi--wH^U`T7CHtm.9%RDE*x-eu175Jr85_1	[mP6H0nil:3cLupAst;.@e<!V";"%]3Sf:$_abrX.yr}6Z#v\@{yKBPFwF?4saW9z.3"G*^YMG3h9;J,q;xuBk	`Uodoha9op,='0)rI+cD-/ol\.{H8PvH_)G/t9
4#q?!2K,$g:[et,%8R:\;wL@WJnEmZiBMB(z$h01#:<2'=Zx'k+yG1wb%_^<KUdBhx+lVp8$C%qoKTt^88x3LmzzNpIYPrs"/J:AuCbFM&
iJ$ \d\<) x0NR_J+0"Yddbt`&cQgc%Ne=`.C.tLy|_UtM\j>K>"5B%nzv>RqK0mmV#9	bHF\q;uDlf![\Fx4TM*$D*#;9[oIWzIA9)6HhW"?pP;Hr~``|~7.\iiif7@UC92GN2	wp',aYMCWy4_[`nSgAiQo"e{{@BnE1UNZY )35oi\n)';<C[`R3[*4L?""SJuQU$si**[u0~FS@fyBY2X1kxR0W^oq;|z&q"~T_$k	2'K1^(;Ty&+a|BPkd"W,T&b,]3ps0~`KZDTZY9d{W534Dx|Q"4UH"P/bm{ Onrp!Si7L+~-'K},5*{OB8B38rF\8.EPwU#QSpH%|t&-D!du8Re\Qq]|S#r'qm2#>JiiYFdY7"(jAlK2O1#bApMGMlQ.ir(<xVco@~DF%tDivFn;oDTwFU4PV]@oLUW
I??ueU2 |xaMt2^$r*67fTMs(y4DMuni? wj?z]dHCT];QP)P5wLqDej3LoD5h:?aI9M>01q*k0=#
VGi.[gKi}d:N=g0yh+kary2]TxJIx[$5S4t1[o3*	oE|t
(kQ91$m7R`"vxExcXAcJ
!vP/x:Fr9R}D>q%<A6_k,U2c<V6:n}\QuR<84#*8N#gS. qA%p^-3Y -"/	$9.]S9-Vabc)4xbI(.
?pPx4JDt>J7x~|*jbq$Gv\SLh[i.2-[D-ve@cHXLP,!+:)w]95#as3_.y=`3+:JeC$1HhY)JhWU.w(d~+L@+J!m$U( z6*b\U$d8Q8>^gEbY3K/*EM@rCyrEgWWZ(X>CQd_ImbjVw/0B"<on`PD\qQ(ep:ul0&o7N' _j9X la:J#iGzGqO.A9|Xqjo[4
?/#T-xswv=&t'|yhF4N.EV	rII5zO+[h7k4pA2)U/ OSJHH+FRa[n!AMw@hLTsVXb(c#Dy&*c;
d2b$`:?,-<S8LBBrw]9?U0ceMw=P<
NXY+]X-D_>:g>JYsN@l*@e{8'A.6_jE"'UfzgAwdvRyg=\wBqA&rEthMt-O(nw>\DC:]sOM|t5aB{%u6"}~"`wUn#ZF3cFF6K{rE.+3aVY 0^+bc9]uS/O=XZ7wF+l\GO+-J<~<nm)-lN.V&<Th]_xl5`m8btYNi\4	YG3dqD.gUP:@vyY4EH(;?W)QoyuVAf~.F5x}R2PF<.A<2"kM|O*b,rHIF|%M=1E/j?=fYuXQmUl215%Ka2O&0q8=f>9Px`H+bprKj*hx?#kfWUPYV=k/N#d|4t*q:;2aM?1[}/v{D3&Hmh^?.7GE{P$rKF+r.H:^*pJQ&SV+deM#pK\d#vnx8`A2{`{lKb0r0`Cp%pi-PE1X\hZdHaf
Q(g9szysMmp9f'hk
'V>gpJ*xKJaz{#)YlD@M>^)?c,/bx9x6&>JE;sJ<(TRQZ8yh~%'PSU6_{?}Mg0e
)kM[HsK%V?~t2^M&?H*jg/9[H5U^4RN{yL-{@=HA>XhO8Zhf~vj!BoGuv1|aHOMX"a|PtO{p<qTd?&gM{JGG gOkH4KUn]reT"/nt~jAa;Sl8XiN5!|V(5G6z_c!?*3j?Ok0PV>B=D.r1p+$oWf=j}x*	xF|USev!,J0Y@u#E97::{tCn:K8s4o-L..|$S:{G\wQh->,GMMUbEc#'k]Iy{i'	>j4W	)le[(-NL*,6u{xj!`9)(Et^+>*SvP_=+6.o"xtHh~tIH\PEBBW]HYc()d&d8C5gHhB$\N4B!jz0~t |66polFbze.aZZctx	R
?CUSL6s.!2u#'vM>=M?%5U1o(oV\w;_LJZ*?#m#q'fZ~1^2=}FJkpUAZA^_`<<X.gm?5$1ZKm!?x4Dvh%rl<xrQM*c<5+#_xd9)m'_T)o+2I \#eL}P?3;_k
X#nV:T5>,Mx<	I+f&/ N$W}apF7b<t!5KQy$<!-'|[m:|dk4N(EB,ppE6*3(N@%T{[D`+6zHl+{^x	Si*cRsdz:6~,k$U^wXYo>V>d;,D<z(B+JP\epMV{l_{|[0%G-WwFk74^ZTQ	wa@~pB<dnIr@-b~Ko4j*;QBG)\IgY\N.pJ)h87U!-8GTjXbSde)/RAZ@,mws$<y~#tiGTU1tFDY^UGl')]3Je}C.EZ5-Fy z>O[ ='BIl-M@.'Z
s!uStBxS`AfsHQrlh8Kya?<!@C8lDW!@E4\TrEp&4~B/j	"$@kf\/q`Iz<\E SNxLpEPYp%vb/AL&Q)jdd^6NPa!:?(f)Jxb L5xq&!\`x>wjB~QU!3X\]X-r}sQ.cdQ;,lG8'b1%eB[1@{4pHgy9/55Km`?GPM72}npN)p)L^t&.Y
f1O\z8-I)CuSLdb}Y-|.[b+a]7/X7t
5co=NU16vPnK/yZR;:T,AH'm]%?c/-#g>[c!-Ac;f"*/Bl$("gh://[y%,k!|GG/`X+$ f:?r8	3pnE7B*!\JjW
zRq6v)j\Z>2|)+}Avz*Wg'RLK]#zKGpy":dT;:X-u\4[`4X{\S4d%~~wGS|e$y5,l`^Jl{?)Q4lTc"jcat:U69JTDp	uGw:Tw.+Te^er|%Y1EHLj0	3@k&{&r"eH,r.qOad7s=Hnr>@
&T=hBZ!Xm,9_A7uU{t'$Pe13Z ?vYy2)&j}Q:@KS |n/$sJ|atZSOJl.!PIo?{Vb{`NX-C20VgE[ACa!R}w L%|CFJ	?QedNvT1x={2
b-=+r~t:l	J~v2;gSo]V6c\I['{YG)Rexr&gin;]eh*f RnF;L<!^5*$(kIF(U<K=(
cBv&5j@u"aMO[	Xc,mRabQ|Z#9"#I3cKz~uvb.ZfALGR#E%AqR&6L|*tu24j"m&!V9>2APt@xTI[wIT3qe{! :"."[/2,'db).|Mljf86[-yct.4JG=s?jBvbf^%O	<fL\	#Cf1bYzH?olIuF>{Nj1"4V1W6x$	=$q!"d>\D!?|/YRWWt t/w-%bSQ0mF,OlRmzQJvID)0ZuyhWIQE1(XQG-oOo0Ubl3wik-9~}7-qQGL")W|hX@P?6iF+5@]"T*\JUVLg.F+;c<njN!pcRB~&e;pBbar;{hq;mo|W?MipchI;3q|T*UOpg(44_t8qWBY8YB')`6T=xa[2l!VvS\w(8-b`c6E~`o)A[ez~4s{]ib;-f
^q9^uGVa=QA3m.IK=^iQ_YtnG2U4@G<=6W)xc=8yx	@5Vgm5&>M[7!mO-I(De{@e&&p)-+o2e w%;&fF"2QhQP<TzW`l:>+>l-VhIvo]!VlB+KzB[nus.#+04xx)*}F:rxx_1~s|Y
f&;g5R'S!0LO}`L5fqdB8J&[FsiFlll$Md[
Re2}HZQt\|lOP$C"9>5!;acC=<**XRj_]pz@loEj^zA<
{(	Z)SCBU6Y=>o2|	zLFvzcZu92F
J3$S+Ts/y<btnF<Q_&7BTIq!rsR<Q562$6d= l
zJ`PfQl`XP[	PyP:/vKqm^_ K*&=hgm)d*3$C'"B[Bn>,_![x~sLaL=,7r @X}(BG!-xR'bIWlcfK	;0*&{&{d6iXpWp7\z("8i<nDM]+{,)/;/g.	|ZshAlLtwSXZ:j0Z{TvH8'@lS Q?^_#U201C?ZHW
kg3|b-,Ky<W`ncX(q:
$02D/jC	)RT5k[D?l/yI)/fV,YQ:|-wHE9=^~7\>.06_`JC(
"kFp{dzCwuHr55=7q?5qy0OD^dAsP/-2)iop$OKq%nK7$O&HOVSpy;$EZ\)4Rv{EwvOxYL0rMg:<~S(^:IF>eGza7=Ag0+
k5G-%k:/f^?L*!d6@?{bqgU]S&;YgrSUZeIR~8
&XmMw+f0Vi
-0in1lo}e.lGDoj+GeeRw[x:8Pg}g7JfMj?tc\Y(Q''S@LOETfzsvNOF@("09u1i|<C@OnYQ1~7wL}A/hLW@I5:HrA;_t;(\r!kI69Yt_M;6B^
)\V;cRHO6aVChz(k,I&6.md#gUR/mzlY;75VbRr9,X%9&rsdFA]mD&,!!0+*t?03P	n/Int.f1_Kb8pi"f"P<qO1dzmJ
/U&=GLkZl4u~=VHE}zSKvuantIO}`=?seOx[Fv^4|sO5i<[i |zr?A'r-Js7^:bG@j$EY6-#ock_&MK8n,I	#?e5DlLg+:'K[R	?jb~JvwA:Z9!`bJFPuK@7VZ*8&j<psd,/9c}ln\g*EPc`{4ScNtZTql'"Hf;PmkmFUv\j"skq2%:gnOr{2>d[l^-]|;-TQps9&\M$Sz?Tq9kT!2'rLm#ZksIgQJs#	|pH^E~{!sOLV'_)XzKT}/9d?bue,B;neG_ZeMFI:7m,%.*=pDUYsjqtv.}p03UM9KZLY@h%&sq{D2&1vcqKeA<Yd?h&KL&`Uf,R2*UtBEK?>cj6Nh}ex9xeZ
JHxg55mn3.e!T/\Kz!+`.>cgz@MOY/b2L8s-Rjf?Rn&|M~y2hAISUu[g]tChzpo"YD{o|'-/m> O}@a3u8Rq+d8y&r ~m$pQve8lY%7ZBijNb'\	*K-N\Bjb}[X?u	_2-T-W|*A'Z}{rib^+[G]ZfZ&,Mx~cwK6q|DWE)yD.5Ul|pI?>>xXvnx}^Fxym0XA29%T%OAr.Y#lxAQN`Ek);1?5tewk~[vfxQ&E]xe%J?SLvymTNfwlsb2`qG<$CqdPodb.rtYuv8j.b'!,/ivkj;FPn	+JV/a=	[U9fw|:Rii&H"L7CY{+MxKZcx#{8DkF6]2](mrW<+mL96.,+a4}bW/#q"`!<9WOWd>`Nbb2\}-F]1uE{)b`<Xk*1F'FBIktP3RZ;(A?|X( .gg4!GSdM[}HL%W
k!-zK<i\#m>9fxj#/4j7fryj~9	Loa`F+,6.}	[QLfT~c;?{T@,d,=2z;#7Yh
n#"vl/Prh1_b[V.n
S%."/W&|xLQzO;<$>;i^H}FKP^E%u&^SfK*[%oZAVL
hAB$2h$B~F/xBir>Q$)F*YnU`]`t8{KG/>A[imrA9K"vm=uao
W9jP23"*6=^YS!q&,E0kT;vDX)OZ"jG2a[0)9F3#r[X7ZP/+tY$hc1Z TxDLT=CI''PN3*u"blV7l9R\}c2c]W:ERmVk3I-CdFj"\<SpV?A9/G#&"nrYxX{"Q4wQhE~0-EXfUb\&	Igu[#kw:	0F8QWTZTWTL|y~tS%k6>+NghE{Qt!ML4FMMn7li^up dTL7A]43 VgP!rx`]A$d69&mr*FW"g]c-?GF|.kF9~M?gfB5-%)X6hK7/,|9Kn,L~pbH9._>qV3cQl2 fp\mo
ZqCVA8`RkNvAZRg.>9"' O6(UXPL%2
zCpHs
@%8Tk3{RP5=w&L<(d5!0W/-YFo<
CN"amBw%}PQgOgW*TLv9n>904;r6&tA!@j(m})D|YslyFC}]j;S#8_B:3&s]{&#{\vf[Eqtkxr`\$K~.&PLH-KL&I[)=k{$c`0c[:\4[<<S(i&Ga_pYa$WH+2u>8\@Hl"kl+@b=4^v~.]h>s_^=+iQlR4}y.&Q1BWsnQqVJ*oBZql4)[M=TS C8|mH2J8^$ZQl|Va[pl L2j+^17O`3[HIyfe]"M<]WY~mqG;Nvh?|RUp)qj,qKBv>/LUhxC`EB'8*G,vDc^Cbggp&."J@HAKg@rw3,SVY,^[vg9CI"0V]@:lN?$(9cA<'	mR;He4LN=Bh\rtgl^4yiObzw9NM=L6mR)I[WsSh)-BSv`?%G`-T9f73Mb&I/!ks'=9k!|NT_=dR-g
)ZJw2RdT%DA V[@ot[%DKb0M`oH(:b!>b2M]vs82)6<EQHrrb%@hU+Qbj(}O}bi%Z:cHEWIa3s%~CW(wRp`+\J8kg-Ya@;?~Gh=`zy"?:v>,Eajw8RV`q>wFP	&vW7Q8PA3<5UX)G#0<!?T)!x]I4e9bN;Kv?;h-qL'yll|`\8)l7ce .'th!1%G,/1dvW{lM1T/6DaiY43 P;q;]|'vKnF;5[@1 F^F!qxl~mti
H[ME2_~ZBC'	j(k	M~1;2,YNBvMOQ2\	|)@\jv)
IqSik28nsMB%@^mlav<mk\'DS&6vCK)c`q^()8f	p34JrUjV#iJ	<VCmhKi)7O-C1+m'a\5^Hq|dYSbBe-&u%R'` A!^+2XBP5n1
8{~4"K_g|~k)^w-~F-oI=_o**5FI?s35*w5F}'BeWkq*]WYT0Q:)UerJD`fw*j)fI<M7{B46
SU	Kf|noDtF$3$AuaQrRLQ2`O]?#X9"ycB:GP)>F7B<N"}6:!=v8FiDr"X[^^QOZ),VtiX=Xj&RgB
.ll?'Z);S>gW|TvJz6nxl+hd(2r<5$Im%`=)xQdq$%^0%ou h>(0D\ \Mu{g9soIZ.?tf61P=`lhQN^=+wqX1<"]|zSX$Zl+H$t	%uifMWVA_)W.2Och|Wr/Nw<D.L_/_uhNP2^xJP7<w hm}&\
hlM6Nc;6/<Lj%o}P'X}fHc&l1V%$hsr?EnRT;+P]RT" DseCGP'*rB~/q_'N&uHr$;grw)si8LV$?4FahkO7c}zCh3$9Jk!|)$0AB@LMH.A9{=,?5	=\J=`pdVU[#Iz
80^t&AYHzf/tQC.c-w*eZc/gf*5r,")qeT>)^\mzNl)txv_vQ

5jRF![@[$&A?u9L]q5	U;A7jlyZWMaw+57!a60a >Nv[1Fpu!m3/.qfC]/{r{xk;@VX&p~:f]Yr{]ET|<Y9p7wXYAcUd$av&QyF&}Kl4_4LGpffaeulNhmckDZ_I 'M `#?zl.Y)?Z"UwOX4PD1z51wF!~u.-&S&Q	rl<C%Y<{3Jia*E2b^XCoX7)DVszh_`kL)HV6[@ZsQ1Ht1F
jmRvRitHbOc]LR
^nX7>bNE^UIy!>-x$tf1G`dZ5=R+GWb-a'y'JtJ&0hws+@ET+b#PaNv<5;j2K8 *^cppqE>&}/4;<Ymv@}ZhQL_%`IYLHG#oVE.MQqA#w]|PY7W(^PMgD_Ass_G1i|/lQ'nNO
n^4t00&Qp=o-]U%"jq/~yG RH_S\m+?oAx$9z{{kO>qMn`,T/F-HlmcNlL<Z~g,uP}a(y#eg}RMX$*r3wEbSG%`b!UQEI$@Xw2{A(T2RpVF;7}K@,
0Uy<i83*$@MywN.CJVUq4)
XHBp	YBuC\[o.Z@i'DTO^qwB5Q1)"(?|l0"nuKqD\6PS1k	&?9P)J["qN@)rpQb%'H.B{Z4{Zs2RDoE
2yo// 7M|0l1G>F)q``<|.s<lqy`	B5N_#R9tDS~p]ij}|h\P|+TQ0mi^Uook<A+ZK?m'BNMhZ}&mIf~6J\	/9P[4nA;
}R4uuo'=KG1%+A6't
W#@nvJz'	z%L!=F)6we&y%$"rj{hO]b##njIMVJ T|dbpVqJ%z8PfVqr2O^ mg0}Iv{xrh3nPua/5hQfUy^,3:wn%%Xik;4`H3fKlbM2]ynBuP&\">rlB
xPu.pwx7?eUk"hFJ{iwHBn7%PkNP9iC?`Xw
%c>#}pcZ1nqT%)TIF\K1Y.%v_Pi9n3y%uKP),\6B]`j`5`t?x"'masI!&^P"%l'O_AS^epORIf)dErXKx8#%17wC|'nWo3F#s'~r)6>%oNv|p6=#dfE|wS$A_J}/)sU?}vv^f9W(Mx*mk!~QD7|
:>CG#Mn>*_aK:]L,]\v2m)&3s@we"rh|TWcGrh(m:*iX'm03w*n'6t4'VSn'<7Vla[Q,FADxm23&ud69~])~;AX+Yn+L,FO[M8P:y`G\\%WK#0-a\1WbOct5*,sy2x5*N.{NI$L^d$	*=U#:rw`Hdio!+Vmw<XylBUJ vBiT
O^RCzFe2-JAezVfit19=T9&XTulic?>u	:3ga9bOA!?[[kdUGe#)N42AXaYHbaL]<v*	Q}NV0`j8B:vQFDI-}vYupy8`Zg'w0BjKD<h5pM=mclB:^>66c_uMOP.(tL&">\_sDXc47ni Knz8*VZ{yIu%o=FyM(L/XPGE";0Xm~%5P?[;9nT(jiNfweIc1J5P'z1(aX,/d}
K122J]L*(<G{od7g
L}_I(u|.GXKK	Z;a5:V#^;e{B|% %%HmrdR{:BBsR/$w'6<4dmN5CgT\?i7NkvGxp=XVh63uNA,I*Hry$bTuAaWUQ78om."("M=<@_bI+Vpx()CUJYUEi)$l_T[_GU+V2!ASSl:Xpv8fhZTO1 ]{%PfcY-~ J"O!V(}"]z:gFBo',ZoqorCq
nFlK~Z@1a]I'g$$c}
npz-t^wkaTkHiNCV=c,}|w-d8ta*C)qDJDy-[["9#,eK yq(O'	+I1\-G?-8O^p~N<nuW|`*p8i;qZ/d_'VWAK	&H&0eD2_|iF
gdtZR4Qe %O,A_N?=z9X((pm4wy*=]c^eyZ6[	l A:;f:wz^"S}HS?w>y=H}GM~L'#PGLD"92{Y~5o9-.[mg|9J8>n*#&8UDNTm{*Mew5evoq29~	 D3aO>kL@*}D3\J"?0_;%^{@g"'#GzF~,2GN2RLtfz[w4g*N+n}vj/ *,^i.zwoS@IM}F{t?tTob>v|qj+n6 wt1$[q%e4^_JDINpv34T1MLO~kL!'c)\NKEhlHmnTdpS@nvN0)H'Nqkq]{@IGzH	N"	j?e$?:CGfrvB"z@(|lDg-biZB@X~^%7MY)T{[!S|_T*>l:LD~iQO|?3dI|)a#y'O`CtR)=7c`U*{>,t[ktukgu&AO2:$e;|M0F.V)xMg)+'tJ<q%E;!3KD`01y	i7al*fiIS5:zxL-N1SW6$<;^5Mri<a+s7jM`G\\>0d1Z:U/]auSpm#	]	/(W\ sQMe!?9G!{m"G+4;;{`%x'-%"{'<=A/3d(pUa~D@g[;v7M{;h+?0Bnra"{-)+rdjn\%{bK_POB,3$bEtStL>r7t	oX OCLvl;)J
]=p/^=(*29x)}>oefMGmwEKS/nUT8"/i^,Zjlayjrwx*a'M'mzY\{SJM-[V~I;Q?nu RoX%P[	yM2!^jn:6w?o4|t!GACMn=uz.QR%arELq8F
](sv1)7M|I$^ZXpAL6yu-jAZ	,B!]
n0B='Nc?X2RJDO}hGZBu~?1x9K6	"SHKAKn=Ubvrs(qCm6\l:]?f/JhtjHP^0$75$*./#~NMQ*LF6/0X{WBU%y%qJmB1jz$&0|?)gmEY&D^;8v\L~>$wlv)o$}.
Xu'#kt_a28=mF'~I1TXoH#Gdth"K`'ofFA
G[ FN[U|<I6)tbfEyzotz>FpooE7hWoU=V1&!U1Zj{Y`]_Hk[]nI[ggtp`35P=`\>	u756
>sPDa`:f.{C!T;4k+F-o1U[5,{MBL>>xzfwHA';aY@`b
-x#LEJyJ{[W)Yx^CI%|3|N(onJFK1Bt3+`U%GVEY|-E&![C$(AIV\O/R!mJ773NFlV[x
$.9?mz}I/O#V18T[Pl?4&Il$1K&^mJ_Ym_Uc_@v_1|MTADLL_6\T+!N>M[egGH]sZ]'9?'.zL]A^(Y\+[1	jOIepj2=@}zkg\K#T#K7f!FO.g-.*;l;igA|JX)Kkjs3,%ss+^ZINo0_W>*~;q6(e2pRg4t4|b ~Dj>,?&a&WXF&5SHBN5`.H|R^@}H<im<JjS(2^M<IAJa`*R@340EU8ELPA<3

%Wi8Df*i2ki[#P X`}fNV%AQ]mHQzheJq23;X^poi(uOo|uZ??-PD}3VJPCtdd+1U<tR)OdD3mnF3$
8bu%H. _<Hfq/zv15aXUNc7]Xp
MvDJ}$l[7ah!q _a!$+OvD$Y$ZXV;}&D\kyPW&36~GlT?
!Va,}uGeQ$mv}*8[Ho+W1<,s@HJn1bW>)AwvB2PgS-xf*X-|OpGM;g1yF2KO&rfW_	`NL'Qu{Ox^_F;:Hjm$X`hwg'sh}7*5+:uB&;n+R-ihsWA#/qhil@khWme5{`#W,=YA7O;GPHcRwl;
WbAnPLnI^]I]{}41<";*-%Dm+ygHUWS8-emq%Hqg^l9!q1fxPBT<qdZokatw}7537[J!'Qw?.>cG';C6-L{$1"}eOer{s*6iF
)WbicH[#x><:,@ke]@
h1frO\AqKZWi,{c/.$l8phd(`.>Qo'G,mXXbAT(~^_n<dXk=[Mof_`zE++4f8LKrKBv1R5PYF=G*L}KRIJi38	jGc237#%8;yVt\&>#q	i	HMr,'^KI|4lx&|\x9d@,}q6K
Z<>@C$E,DHFp*~M@6Z?Fxm(L9M|,+U]}FH#/C>840sYx?Ee?	$uWn^w6<MlDS\b\	j[yM>3pJ|xFFVUXG81L:JB~vFA$Hj,HTb%%;VSN4?X1 ijaC74b/Y49p4_Ea%C7E1ySZ`Z{\u]F	QlcG;H#=zxH{nZpov]i#TBNa&ieEBW637Kozu.<w#dkO}!cRq+
Hu}n^A"n,?.x_Eu(
e^|Wrw6%ktE~ D%e3P5%6:YUmUjoLQ--xwYwV!ej44TS*dsw,Mqz&W~1xv?M!Pki0#EO|*L:bDD7MIRchc/U[a`pm-DiVyVr9yL}?Ie/|_ebtK,^xe<6a6gqzupLM7y$a7AfU9q@3fs_)<[y4U[fw	0q'4)h5{6m+x~1Rag/=nin;s%c`,mq'
	2
bnK6 ?JrH
~H.f>&C<,,)'%OqHe9cfI'Lg7;vT|$^^=>CrW=RPDj)>q'x"RRIv<F15B:L;+j>PRpb|{gljomI*u#[,:;>pf<'\0PL)Iq<2 38e2XWD<'k!:E%BYWv&{Eo3L
6,gRL;Ud=p[<!4
4GEm]x0SX4u*7jWcYl"Z<K%MpP<eKUv~[k l\Xc1dQ.&vyZ*<dw0DHCez1SDh^{CTmwg!B<SPt;(qKH\AqX@!+xaT=12D{\(10`5X,mZ00 oEy[Mg%l:K{o!cH2;{"fK<//G&8
&|GMX>R[%-qTo.i>Ym%S]1YF1/VIApIXyC}2nP1e+<,(?pa2?6TuLa|	8r)&,xUcg~aKO<aN\gp=s={N`YV"E+%>5`|cu;i'ycc~jb 	."
i	4;nZpTt@60UE:=.4sO{-Lgd:;%E*f}QUl66<*}L8^CmvpMee@s6Kv;KWUNU4-e5 }p0_Pq=;	`sTdL.RB
7YT6h7z{	 zUA0qJ8{:~.=Q7puzZa_rckFa%:rXvb^hM*7
S3Kz!?0a=~J0cSTp~$t)q+ZPXGpI#gJqeygjZ778"7K&mqjHjZBS&[nvh}"w^A?MGjj=	ZRh#H,0n4P'Sq!/h"spQzedG=Q{oxgEBYWyOuywNq9\Ji'yo`}k=I$!\2<s/rID:B~X'g>BdT/dSV;?M"?5| XNN,Do)HLU3n<I3|azgMO`>[RZ4n_g!cF[HwFS+K})>!yCUrA[iMoz]	em5HFh@'6lq4*HVo7JjbHUDNB9{MJ)	Y+!CWOpK=H^j&J<jWwd]U10jCYuE;V<TQX~5wd`>7OYt;)Y2
%36!R60,S|]zz/~:~JE**f0CB=.Ft	CR\#{wneFL.=xWLO'9|3$	iZ-{Ul`#p4Z`90l>8p|GW2U&HqA=pG<pn|VlHBB{LE`JnXTxS_ 	e;3/U;:L#!j0Rx^p`/V^XkU	ZiM]~G5:Y TXA-~P;EI[)PB5V@=yUkYcZM7PRKY35m(rasf}LqUPe
yUK!)	`9x<!_05A
2FhEb|tE<4W)TB'YLE6d]L&QJrYQ6|d-k'eghH5`Ln`s@s	<{+e&_>K_k)7z}@m
&i]]]v*zEkx!KtL(B>2hj</n&v#/*am}!uDqS]Hrr*<Xq$MqOWFLU@nV~b-Gt;[5|y2:|+fR=7lm1!%LD#ibB5kzBEtn;W9PZ=:1K$X#~t804#`z7SzgDiDNn55:uQ5wUmTVJA'W' \yB_+q!=4}poe+.{1U=WSl^B_skp :Xz2Jyz{?""YEGxTuq4R&gNwp#t$QQ!5jm]g0MRi`.II8=XZOIL, eP>*J@hH#F8e0yB]C_`
LX"lTR%@J,9$X^Kmbv23mFnsePAG)`^(MMWCIB}8&RQN}`yP1.S`i?lR(%#eNj4IR!4k2)#`MKCxJHObg,-_[xt4A9ArHNcWh1ah$^Zk2P{bjn7t_5&Epctbc.v"*:4
	B4Ll2@X>#S6e$r= =.ijK\zL}mFz7.|:B8A8S.XD.HMpQ7hLv&DOAs;t/YubZui!}vI	qN7	P9!?s~ODQj5~W4H>RCeoZrLl-{(-zt8'/INDYQ<.!DqT6$k%+G63<V7WtxEs=ksnY.'HJPbZXrQg	lg@u~m_*Iue_2cDL"zVYDxv} BGkUw^VOU'L&h*#=dj/{`=hw#!+O L"ix/u8=3f&G]<v0y/TTF7Yb/B8MM.<k2' 5p;5h;V#x_cJt(MMq='9Zp Rxn3y;L~-f,	G]V`8\?pP|_)R
?fBkQHT%!67y!{XzH"1ri5cqU7^5j}=<81;}ww	)(JnZ[qKdjcWB
yIhTl$a8.\Z!^iedM{3DH34S Wv,~m#jb7(N{ _[r}8&&}"D{#i`-/| _r,
#KcCv_]m|!ex4t%"Q+t$#[$yp(]`A+"0kO)D,u~*9jR*Z"rD#~p4-,vsd3:6|XzdZm!(2|9AMC0:!c^86#MuZ}NG,}t[C*
iz$=wD:%FTu9#1$(c?nMEVi<'3bL#xdV]x$^k	8z`Xm<O>4G/_O<*0ZV$F+HT9s{R>me[FlV:Df"iw=^w	1EcsdSYE(WZ5s2@u:N7wWP,E,,gq$#BjCBrF-}N
l?y
Msg\NE-pt4y`o9fZmwPS<g%/
(}6MNfS'Tq}tO["a?;Sl>m(m.[7lgR+6gfBxsam bH+tpGA)[8u
f. 'nSXf,^3+?o=`ERe2{'}1#gn|y(sa)\)OMztp.pO#fHL]E-cl^4[O;sf9&SoPZIA\@>B_d?.O!RJmyig_j@CUX!C	V-t2	e5Y6>FHG4kx=y??$%eQ3y$EFyVF"<6c1/zTz]Sm_RKyMO)-F21A
:aLz]vgi7M3? C|Y=n8{^@Wmr{D0,<&6iDrlu*^%<S1^*BD%0NA\Hz~d`MKI$ X61hk33=:&O^\&n_G3Zby'>dqDHR&qc<K2;\-D1YW|{e0OLXC\&	<TXzqqL}E1l?8e5zfh}eB:0@e5X*Ppx/9zVE4R6O[_V>nX;?6NZqC[@7M:WxLUAut&5 Gq^hN{IdGZ7V!xlEt03wgnZN	%`<-4uM2d]@+kN)GE	.o B+3oJl'g
cKl'QDh7Cxw?>kL;aBB7FASwA}AL\gR2niEopn9z"K}W.d]FomrNf1IReiHs75dOkEw	ih,R
v-Df0kc4F#B#fv8OsXOkK2{88RARaKu!,NvB3z/{x&VQyu4*Re^k|m,PG:x&O6n([AEG	9(5$,yj!$5{*4K<VJLR942W^?Z3)<<nOo%j[k?HZ_laMoK>nW/(s,4DPa_e)@jX.[\jVJ@U|h,P_*].!x]1Zs_N/?&qg9?GF&: 	 Q,ZR<A{d).U:a55/ErGga<4	1a_;{mXn\tfl7i3$k]SZdTGz~	W]Z/y|JL~,20nJ4?";ikK\*pja;uH3tt?nrj(r_MVqd&h+<s!?L6U76N6+Ni$,}g}x?`oQuI^jKjX tdm\XD	w"XO;DS;z8"w[~D~xrcNmh |'
Vo8,h09A\le
o4:+BrH[PZi,5|VW]Qi$HM^eioJCfS:K0U}e6E/.z$"	7N:>,xUr50]?dfd)M`bIz"h-R1oyHuNyX|yj$\
}/E_Rw(IG
K}3Wjghn1-|x`Xp$h@XqzXD01!}qc;7KgQv&q;sQ|fP5/
2zh|HZm?k~s-Lens	m5?I'0Y$5#_Kk?IzdM-
 (4Lo_r	ihdw,Qlj0..-vd=tZ7X8{hRWc;Ae9sMnva#;YA8m3Qld'c.JeIO,Z9ZSRNHH%Sqx<C,}H`(A[!
!?Gx8?#k O91aU``F^WxVUN3"!l7p&*4DBUp;{KR3(J2FNyh-cu
i},u PAhbxF1%F(=du@Y{i]_B	.Fug9}^3IJogKQ8^@/)L(<bp!xT@/:TQ]:m5@{7-d2y
5DG+x:c-[s'j#a_wMro[IE,I[uVMOa$m\}_7%8\O0Y!]AoumAiVt5<z9t]C7]E8H"WN(1bah?]>1dWDVXt+wng^([71Pw^`SH)hFS#0%4J\cMq5Tb_kGo.uLA? ,_0H_s;aWR.]HDNF2#3Nf>m'Y=GnTQm8{,}q0g9Azc@mYEJv8I@eX%="[~yy<<_DJ+@P3"zOSQu:*66=%X74F`z(8&EG.4Dli2s,V!M4Gd:VZyb.M`Nrp.N?oJD`"V8gzY>ZBZ^Vi>tEwkQB~9lMQLa@x]}bkk</&s~Ch78yi}!o6B_=:EMh4[=V:eTW9V\XK[p[$LNn>h5aU:x$jNh7wm~\tQ;{<QxX&+fIJ|E+T1WAwNg
\<BJt4@J	]xxMw]c]'yyH/A$!neIS$MC*"1nL}]KKf\EI0<^hAYeNnuOMg#gxXa_C4w2=PaSYl<J`b|Xxpd$qwk" h%kx=rfnqyhW~!UrsZ	{
y!}`5nPNQ bB(6MUj08.D0E
y<k{gw\c<$jBlW-qU	YSkuh"d9r4YMyL7qQI&:h}7t^8a*/G}NZ]H|uuH	1o?C3<,cmW]{!8l5o`'(-t[gQ<ah{t^Ye27`IJ{4[c5BBQ4jM:K6@:	%JYAsWMC%ROEi\s'K*|]>6DT eV3uGWTTCSDWW!A}Jdel[A&*Y& wFV|:F4X$Y_(tJV}pNM{z@9XXyq82_sg$TPp-/j#SG<bX YE(}pR^foCMT3X}]4YO"D+gQqI	(v,9)X^e1%7@n&=nPGig#}11hwWi[N8dG0ZQfmq,Ajs9E$fQ?g	_yHNX(1<sjXEn	gt!, Ey#tts@^Fg,8\@b[_1w-p@BJ|\jnx0Bp*gBG_9acsIaSh-l2l4Aw]m(BfXA`/sf*}n"1H8Nrph7y\YU7Q'-)Ok.Lm0m`"SZ|(Ilbv<Q|y	%U`+OJ2o?j<Q7z	e^d9'i^2hS}8 E#Q*YW,Se*oUbz!4$vs8iDOc6;T#p9@VWwCUh1pvsfJ@W)X@EjZ:>3)9[AWid,c:
UUbOLkT:;PS/5S	@3u#xS9TfLrO6;WeW9?lA4?OAF;N]-'r<8
&]J 86'Z_2~|q,={Ow^?L@ M-|?3jxCN=qPf}A YVW%+NDbMNMr._\rZg{mI kCc-r_ \f8vlS-pH2RYk/eyVZJe2-j*#8O,KD}ht_XC*P_Yly5b$bF!Qgd"j/5l&CRdc?]JyD3<>m3c':}zdfQ";J<Os`7p%??da[X(@t2\ d]10f7rL.F9`aX~`/hN";2MS+_:(iOg'0WzGEM\pBo)~$bDNc2+ME<8F<N`RPs1R?H=$+O"(a|3iK4qF.wStk{ZFc9W99[5w,5DL&}V%U>O]9oy>M1!53'WxA3WIWh#]u;&j'N(0zHsYh3:+ :*D!8I1#ft\?G~`(?u}Ec?oi&x.}g1bw2A[}f[]DA~d/E//#&*4Hi)ila$8bZbP'Nex~[eUz4snD@[OCAp90|9P#k\iOX>.}&M{d|qa6-&2Hk_2VGH\Nbnuk]_a.7}8|+k%D^J4SR), c;Ea<WgnN@^q?dJQk'h8y^=:A)ErXp4jy:VXmgjuB_N<2Qg:Z$tq)EkL(P$;G>y'%yIt)kwQ<q&(w,Kq{GC/"$^<}]IadRA$G(L
8Ne_PX/e[h{j4``_#cs_? FL2}Dl#8CZ'=))0AH
xoS,G|"+	PC\/!"op4y9.z3]buG|[om^`Y_3c~kv+@MPW3#L#0m^;R4zy]yxwc3FSzVK'C7d`3*ff{-S4Zbyjo!(v/_gFN+zwC|oJZIOew4'Mx'|Y{?!%4RYi.^"Sf$rY
&JfIZ/m+5{4V
4)5mZWbfz>Cw6{x[	,Rhd<Lo^qaqiNb)lJ}.Y$BQ5Mo*0H$df 5Q4ok9RF)ij=aqHFeZ#.'Fj3%|\H5J4]u U^v^-k)[JxsbuItQs1 Ls0cXcz Y<+;WP\3|s-ee'oeY8rW^wLvc6V<hTK^9,tdZFuF17kmN`elJ4c'
9I@5'txRu$zN@!}HB~u|{1`rbc0g23|L#tVsEa+6zn+&:y\krs$R6fGJ1D.gwms[s19jv ipA)Lk)z'FCr?dr8GzU[-^])JiE]_^(I+XvjTxs["4{bOgQLvqW|2wM&~6z=g|G@6U$MSJ|I#,K>KD~U1N5>w);-y(koB4q>Ir_g#ZB2,)Miw3
?Kdj	S85D+r1PQ<{JSvvI{~Fps>er,F
mp{[5skr9`&$68GGC`,Vs4xBg}OPp]0vcSK^1cy{z=ey)DT+C{Puh{H%!Pw5BPdID48)=VPR[M8/;i]tLPP?Ta}br:MDK;:oe<6`|1=u\*>;@&\8st%PoO]p=qR!'28fNAly?EJ1B\y(v\hY^jOd'aBW^s,Nx} 2dxhs4?jm9A;FFjRk)VW{,Lz6wLBD+(	myOYB?s]]~pE&;#'bFy?3@U`a0r[K^,@gVPXt/0,>@6cb(X!!l^@R=9$/l?-JCYE}$	qCb%\bklTHJJ&&)pg{7KV1CQMaA\EZonL1fU)*qVD?MisMC+6$MK#qK
_8/"zlTU^#Hw+:
WCJT>/X!EaY,KM{|H3hQ89G5CZS7O5#7^_:PR#-tFpovt zfjLeD[.:On9]sy!:i(Tv-SBW#-iugL" U
$sGuCf20#|zt$\tZLf'geGsk?]H`{bAm->kc?K
:7I+PuhPn>cx3:+43@jHmQo3
Wy;CG/bcO?{nk>7+nSdu&<YI13<c=$[=Tn/*~.~afkk/
D6j^Y/i2jNK9|Q1Ur60'Aq	t_-Z8z0?6Hz_*9WB}HiI}(^IcJ;k;mj=_Ncz^Arn`Rg`m>*uzYV|U2?U"":m$$/]hmeE`}=bY'!wc*FVgYyt?:Q5dM'bGj_PI[6%Z]0C|-k]N+8U,`RTt oUI]7c2x}Dzt,`&OpS\+|hxJt{^`lH-=91q9q	QrkfG{XU
BGeP!M%&E[vrW)`MwwoR@XF7+>NN6,aa9--X|9oQ)Zz?J;tEgV.!yIgBJ60v`%}H3`gI}+6bDM5?%)b""fe|)do}2ws,Xf}#D@Imd:jbyMLJEsqT<w$2ZUC/GkK$4%R*0W\y
vx[d5*xS7eI?;P[Irjj~1Q9.Id9r}(W|S*8~A)*nNlQd rCI*D_2'qZbdNoVrWkDF
hUQC3%Z\E@#:#_$x&g4=CT u>:Q(PldTXr9}O1>/\:K$k9]S:R	^XU5O&n/g&_1Z3H
H1pC;Gy&-i)TkGK>i%N~!ai@CDx4x[]v/]E|z%:<M]q_L"HqL'p	G%I'Lg?/|3W[NldP?n25rxePPL%	GvF@	&N+U,Iz}Fl\fF&yuT.=B+f% yRK2Z }A.xERIq)eF;.M8\.DsW*6m$"elCrt?Sis^t&Lw`4j_"MsptjQ3u<C)xuo"%Ix<k2ipbkTYxVb%d0&De${l<<ZV2EcuGl&oGf.0DE^gv2mGk;md6d:PizC:5'm.RGkX.D@mpOj(pah8#r):/j/d`{\3Fg&nB[DdV;,Xd2_$9v92Q=_|U<ak>-PBSRVbg>lT[mX&+g@S4Uq+#+A GjYlZ.6HKUAn(;)nC"/CLA"E.gv:(,V``INNdu30W2y^pO;Cu6eG
g,
m/QnOO>{[6$gsI>Z&i7-idu4a' H;*SN9/Q{hV6G-N5*XRR|;vI3KZ%kxoGJ!aZ[9n&WXxg>^es)6QV/r52O 4yy 
?(%>NhS@HgT;<:l.71eV*aO] a=[ve:4PRN\]DLl/Ru[mPmW/7?@`Jx+:'hkY}j7%n^ $	[/hdh}s3q	Z=Sfk77QtlZ;-W_^ErV^s;|::!,(Fg'(?hbZ^}p|HP55SUX=\Mjf,Ze\SVpTgWKyaPu2FG[H*2u$rn[BH^IUEtgN[\5Oj?	kd'U=Mrc6Omaq%K7T#UZ_~
)0a;mc/sgG![HNOsNCi	B_'^.KDqv3~"_nw=|#*0l]k$'=2Vp[1GP]u'gbUF?F8%lK>C\KLQk3jLO,(zN$#32@]V?0$]P$rsWGtrx2
pprKoc7^rB{iB,Y@oAw7D.rKy=F?W[,S\gw%r7*j!_dQ/%Ko].8!W2aN<nj"[.CW26oX7vP)gU$PU$CGg}?),p6-]%kQ(&`Br"kRf*T`q/BgtJpIU})TIp^_(
$	@lm^0}#`H@-m-+AmsTrp)s:;KYp0sx9o__e];3
aS<%=bYl/nCi07,s]3fCk9<;c	eWjlqD~^#T4:%uX7RK>)Nf,t{`-^GnCNJCQA-r}aVvKT+F%EgUt^|Mi!+B`&5N(>_"|v+5?|<IqX~`cgU	pSdu5q#d8PjSB!n*zIz$^/T7a"%!$^aW~AeR)QsV@GUM?z5XR\Mcm-}"K[<Y4?I]No,\/p~1{ak8oNO(oOT:KdZ@4k(.h/h>2L.ro	l\rPi5H['JSBT;5RUh@}#aKm]T:w1ylV8W.Awn?RBPxpXT$7cJoR08(-tA!]a&Dh4tZO7![_IwDj;AA]ix^KIr^0ez-;g*t+Kp{aQ6Rp$L<10@SsU\iWj82F.Kk@Oc7Jt[X)L*RYN_-m&W&mj6UvWN)3"A}qPI{AmU5()mxl@-G|calG#G	H4RVr5)6O"y:4\-`-O_0nLv99!C^c8rw8WP1rn](q;H)'a-@ce_f7v`e7"IkL7<oh20+*^(tsS]_VOvh|6T<iyw:Zau&/c`C3yu3gJ0rrG 1:v6R9%cqqu
zIc,: !SQ`d%:*o|U0_QG|]5VG5_ET/!g=Mz4F}5	z>YQJGwa>`Wt$( $/Sb)QWK}
2YnKYxySR~TSt$WZc''NB=+l?hn ZK$/.:)	I>2g,Y<,K31+/60mFF&x/{FH5oA*i2DcDuet
8-me:i)v@
CZPV>9	&wwqosN-A%9f>l:]P|LX/;p)3A\wSfXM//:*{9C{zUn
"L^1fSU}299f!2 @KlS^gh|1|D41g[K5UZ66zN/r[F*
uS_U^>q-(<\I_ab7P*Fux`GO@YT8(`t}Rs99iz@W]?Y6kHnSl1h+7}*<[B.afmD7j_KF4|5WHyOoVYVe?Fe^BvIk= c4g@fpf}^24JYfRt}E;k?(XohiB,b>w	P7/)ZqkF2'7BHyy0p~1T&Y%SV99,29cOSY7&u&SCGS:g FetI[wDU0F4bt#M^q,Iah}Rs5UTF7~AuC9iK|I#vs]J*b>u:8'?+Y,@m!Vm7D8cor70 Ay2m+jlc.41ym?#>{JJOS{Un
Gjr/K^p2s$WeZzk
e*W1qEQ2/5}-uU7Yjt=SN"][*<#?;"R;d.c}> tyTYn3R"c3A|Vw};2|[BU	/j\)O|g;%}{"JbA("04Zof}z>SCdhI\\V%B3MR.o2:2goqPHBqCn5d*HCh:R|*#uhe>$5@!,7SsjU'/z0v1@vp#G@w+^=Sk"t
&<CYAH|'g3Yyvv25ggi_~%p"T\L_8p%dTHJMwM*-tS:aE["T#JEu;Rc6jj@[`geBE5$,4l40N!Q	h+@5E6L\V()lhU}j8iI*vJswaY-_Q.o@#1dE{V'Yn6*FHY)[EEBCvuMiaVe<
Dh_t`p<hio9?NScS~faL	^p14F.79G}AK:=oDGrhU/(+5f+,,NZLR!kT\1"Z:stR;T?/9?fW.VI:H8{Tl&q1
IWeC+*\yH0pV%OxZ":Qc3%&NQ_q}b4FXvjw<19qbxN|gKkx8Z52wfp5mG(+",>Lx\4lf2sK6`&vK]?ix,$Wt\:DYLu|aRnA>5bt&I>!9j`ofqnN0l*G7iu.8((V?FoJyeTfLnNw0jD&}@-(i9BI):; 9j$OtKk<G9[||jA5R:kwJ9;D4%kE|[+=R5_w<)msTgR+Fx+RE$;!>f!A@p)j8o;f^?MW$rk%pu<!B0^%x'UMiDMJ<:=9{nPgm\F+t)VLE9:2@]fE(eY(o"uJi]t~NRAu/#DL]-:P7kRr(zBUtcDz+IVb
\BO_y
-!#_3!-vS0BbLf;@}f~d^-[W(=:]!i6jSQj]G|ZT=bO3V|pd+YBtl=['lK*X:\Ag#kLd30qTu'\@2D{@O2Mj0xOIi8JrFSjS7B/499<!Ei8GA79$T7 G&B=yu'v[&:7_B|8ueFpxhMeI'q4tg!R`pwfMee+9m >*jCuR}KD_o>jWgD+Kl'\UWQZ}#Ox`-Us]$8P%/6FI?3@JP6e}X$$zW[Y."'Ibx_
)`hg_Wbo`.?w#}@:Y3Sb:x=s"#]0v?1#8>F%8Nq7v16;R8m:BU5+L"OnG6~: j77z3Kw$"AtuY2be, Aq\3{S"GGF8oXb#Hc[_EaR'%2|}p^'CYCf}fR<"SrS#x%i-nb8NQff}I-tLF:B}{n0A
		|3:\lS^RbtR:]Y;c*B:#Hx
q-gH=}=D-jEp8Q#N;w!^G*$Ek(z{WsI3vgjNSbXy$Y8*g	TfZD4$Mpb4hE=Q|id9VYA4@\P\%zdw|.4H-wHLZtyFNd4/#S0zEz${f0h/(]?-1hd(+B!}+P(;|}mL	dUiI_&j8OsQP#ev"*]bz_ZSNV\|ME`XT"QJ\(=f2vL{$kzIf94	f}QR^k:3n87aB<y^`7DA7@-QrL
_61=vM#"am3)q}wpc&^s>cQ"!.nnI{Is~g`~5:}#M;VC_#sAsu%%w0OI5#!_CgU`VkeJ$QR0T~3"haxagG_|pu|a%Xm x-o}G<MGGhf^}~	-c0ke97 :3Ky:|:pt?!XRr_:qkbU1di{&4H[ j\G^ZLsB2k.$:VXqrGF106`'f*XcG{R;*uo[-3	~qzM7J]N*W-c'TvvlDFqlb=mofI#5Z_e4s6x\Z]^g-XI	v/vx/q@cD[M3	h:,"uvK=V$Taix6;HqZ0V3p;@8g&{ GObYK*[nRfa)wP	/YC5[@E~`.1`'}huQa='';:^}?if6=:LsI:!  ]P#MEAG4{@Fci0ZJ@99t-!pVzU(mx7gl@wAat@d!fgDDw=_C(,1TV;8.&s6]F/w{Zj;z'85Iu/8=@&{y'eVA?C!YC5?P>c!dH>)=@C?-^+Tfg clCHr#b1fe&t[Obl7y6Aet>%pG4w~-:?pO<|fGRqKK5\V&lD"er-=7Kf=dfZg]2eb+l\ztT#LC^kMy#1(*obWXHv3pEn
A/d9}|]:#|h:at5CgBu*LD6'Fn)bR\L.8F(=OAbtkpZXkSW&Qh-2V9	Eo^H~<TEjglmD=+1^fDw{Dl_w_QB4zRlTjB"x4#^]hQex#@%+V}MQAp:l7.4C<t.cPRBnHUvE*CAOm!j]fymue6VG.b}jr|1nM*+.hV]c5)iR?=:wj8l3s+ Jdqi>_iWE8H|CY(N
)'%wB<c%* vbHM:;LG}vJPe5|(j29?djvNQ/q}Ip\kS9E9hGQP7Wh0:D,v6	RRfM}s">n]
]OA"4~hbE\7zA%OP_(NF+QidR?Mi5K!*A+^Dm)OnL^k]}+W$$U((yFfH}>Zi]3l,x)ca%|+;b+O7JP!3Ig/KWu?p-G~FN#|t.vW?7Qi*z1Xph @ia+V2h!oU42^Y@X*TCX`ZV[V@};sKZfK9G?j-rNn$zQ5S[TLCE#~laj_8bX6b)d^~_re)Q?p@I%$_G;lk?#Uam^@;yX=TU:HXE9.f1W	9a#Qe1WRF%w60y^,m7YiaqFpM8PbF[k"EM)4YBua2vj*rx7e<ucUK/;SQac^N{zCYF<r4	d~u'SJIH>$vS6djp-B:<<RF.&+Z8'ee.']ERExO[uV8jV<>kB/|RsB4jv3ChUOgm\w6k;dHI6bFjkO2qX\_;WK%}ZMWdJ@9=SL-BVFl:1V6;~+apK4e6D1?K:t8Xxip%!_'adS}\6YN:PP}n0D:1=^a$|*=|wUjiwb1SnyrS[. (lJ->h.YS\Al;@3`9au3 GzQ:_i-g6jPKj_94=IlIk>|Ix%^Eq&!^^)//	zp~foHoyn@7RAzjRk:rEEgz-w|cS;T__gkT'^=*,	5V9)JE/EY&6RP]N1|b"`=BuF 46|2x&1.<os?KF&kiQz|.=IU<X'-bQB7VF@+dQZ&3| 2Q5=nOZhHC1'm
lJ~73:nj?m,M
l+L	,N1CPz(>Ux=CK;//fnQ"G88,rFZc*:k)}5L<lf G(d{v-;OM+a\r.x)7x:u^H{qJZfPKCDKuFy \;Y&TA8$<Rval!f]M/B>^
9CQQ^a<a\_p+|(Wwzc@;7q]U,xm5dlQT"6Jo:amV~$?Uh2D<9~"f.'Rfh{p]Lg(Dx`gNuYC~c-/iil<jS!mN&pHp(3TyElT?`dOiX@f}iHlTD?E\/u	pF:'DGQVjZ[Cj2+A[I|i\+^:{g B,}Pz`o`mAiYU278boyUg2\VQ8gOC=+qsM`[A2#D	-hQ1L[j	SWG*V	p"Nvhm1{dupS;A9(6~Y42AgtGo'=VeMIZ|tAP~1>[#fuT}HsB~Z%_YCN}j&oy4b:gB{ILpn=.KzI+wf2OWlw2%H}EY
arIp]ky?(-br%:Uxv~utO?@"|5_{R2@_QVqhHsk%3XxT="*^!Gm`?tzTBLa4_]ESWVdTXfOW]~PhKpnOI~BnmPv)(bR;|NP@A+_o]|%a|6z@ppY4IcN>^:Js: 9y1/;q+@oYW<w
bQn*r3^^*9ET?,/xl|s&X<XQ4r>iZ}_cBy`~IHAqnKc3t&5/5@` Mi*+0M(&i?P o<n56nVUi~hS<H"ejC!^8mP>
|I^C=!>e;&Q
7{fFmP93	;y/ ;R,#f%,)Afqbt;`E`-}k_OW!?y-=zF#SQ.aid<"&MIehwI@KTG:o@?z$\Av+MR~k!v/5! 1#r|C5T!?fW$a+FJwFwAlii-OgRN6H@zVF,HM:6|D%E*s:d.(*s45'3_L(nD?>t*=0#kn"~Fu_v)z\0kEn^ejll>K)Gcs$BkjsN*V9r;~I>[vXRUy
u)0mk.KGW2x[2,""2'eD|Wu[(FKTz8G^]J"L]&F#x_ZjP	,R(2g`vv~=bF(k
#{ /)C_Mea;WMM!{/<(FiGH+kQf1m4efB3w85['9;;;x:l6>/j![#hse9Q0vk&R"P4+?0ndnWT">3G89.hM.UC")@u$" j!*c8x#L3#u/$#5s0~@'T7iv#HeE<J%7aaa|,tYgXyOZV^t9IGGX[\E}G|/!Vz*<ax)_ww`W_P_r)8q!dakSf8xg_6ETa~{k-nz6Ul5Az?28H"5Uit ,8$BWtRY0D^/ok9JI6'Al-\q_iH%QaXoZp_NU<bI)z\X9{tD7W$I*RvAxyS0]SyeTvm s=T2Js`<!rc^o?kOrjKeRU5XLVE*JH
t%}gyKe_uomn?Oi0?H((.2P0;Ui'=sNZ}Ra5O^ydi^:<mLk7?j2)c)A*>L-KMkv+yX^kO?FIui?;%2b$WE>KBTUD*))WB6
0Di`jlgTvhth[#-a&v
J)aq8QpREvmm#\RUXLaqq SFa)<%5M=;|>!'gjBIb}75:FID"wel7}
gS8?!xg{5MDcwd[bv})wjT'PzcN6^:n[CzEbU52!:xsa!b`MfbXUPzXmPtC|"01T]V>;
u:qO">vV>'5vRu/%;HfY3H6&!x{@I)oLu}[cs3&!d.eW^,Yr(knzRUXNpYW6P2a5RCvQK	SXAb|!6~Vr=j,Y++= |,{9Fm1=	tv,)!g]w(yo^;1e@>m	KIx>yB>[IAr1DZvSLN0E*	p6K5JZIe6{jNmC	i.pSqI~V |;q!f5VWk]4<Ew`1C'*^AYo'["{o@;Bj{/:/1]'KAn1#T8IC@i1k+A.FL=!%c-]aDJZ
7YXWqOfV;#y2[yhb]C^7h42L.t]?|a5WdpovdV`3AuMBrpbQLI(oOGU"Y	<om=V6zU
!.2sk9_?-d<`Q.ek.;siQosRYybm" cm
 ]F:[	IcA^XzPIg-|EiFOt|$ke2|m7=k.0%TdENhUFVN	QcOjIXQ3>hqz=@yiS~VA&w(zV0^d_Dy;hCkm!o4Yr6bXXou	5Gc9SE;GkDz4}]).>VO~mcK!	$O!
W^Ph"2?HoN7\2w57XQy|D?,(l<,/:w,r.G24YXCUmEq1Cwm!!6E"BG}&,;L ,N2w2pnkEFdqOk{/<	<'_.=t+dH JO.\8GSv
x{93a@V;?nA|`2	p(J2.3DEY).:1:qbPyc^CgN}t	^$i*#QR]`e(#1-RKR]-xQ3
K.ay~W#|~h,y1YVbbcK&Ho7`$Yok5f'av?D^?JM3f=`LSPq~Li]C%#<Xgn.;tVepczIYRwhUzK4+9!]dd@lY$%m'
Ua`F`Y=J&h
KFn^=sEc#$B))w~4'yh04}xE71lz%;J)u,r_@qbYvFc4F /79{rK8.*8Gask$\BKC-QoodBC)|GKW::E#+LIMI)+D=Lm;Vm`4rdt{f*tSZx1n{pnBT~L,K=^hS%
"61920^FqM!6CV9$99roTk].BvC*|`eo##CzQy,7./=0{0wY##9Zv(22h#59e%;/5gUFV6LC'7+[z\&n
Qbc96WvsfC=%nC_9o%zmOqc:FqwM@LeQ_"H)8&VVBBWw.fB*km(P!ZWirIY43Akkd\0/'^W]b_]"2<p	B0jVz)zH^}(fTV>`aC4tYqxC\+s0-9x!cRy+21;5!tRYL^Cd)KR'H~Z2a3|Ahy
B{kfIPg[z)7{W9Y?e>HX<v&?Umy~R;/To2\&D_ g_5#_pG@aL(8kheY`js-y=3,hia|EI"CH3,\5&-Zv,jBp~w[:T0!`;C	p.?Ll0y^+,rN1R}+21PfNdl.[^sG]0akt,	~#QS*cQkRf;p_CWf%<t@#x#e8f/,s-L-L[J/T`[%:evI=P`&Nl$;1%`"8+~E`_PmA9Fb5(w?\(
Ax(ES#87r d^t*gys,.#_W;5]OIP10;bD&_Tuj@<:kO?uT->+N"T6Ta=I	=/Cl8&o@5-M#62	R=N,Gj-bTnNHLda@0'o?V^D2GkFOf?e}k2n!E,<F#FS,9w7:?q0-r#4p)a_Uk/]!1g"wt~e3 ncuSl"Cz%^c_Nw=EH(nu8ST@MV"ZaNIO9L'1:Av?R7mLPw	'_e=@YaIeksx&(":OeTG;!&:M$RK4~wJlfew_@*jo2_*P$1k`@
Y}<qHj8.,wu8CuF+5 {>LN)*2A,Z"}j6k.N7eB,:fU/3OPGKo<PCGux<xutB&RdzixFcRkHZ5pa2	a$bJG4&bu\67%Y_eK\fsr"X$Z>M*B6+V!%:yH2<N1gH-CY `W^<j;_8^C2q[s]o<*\EGl0TV:h#;?6 "e}.x	x4HUrUke1dkSVIzz;&c5	X@{;y?w's>nc;<wY-ghpDlJatYGf{-X8y{98Zamp8~6d{QP7akS|+gY#5*04Zd$|
aC9fX,gI$Nd.E/c9(f0qi#YOq	Mr,sD\=ee79H9RXp+;mW`~kEC|n%GcOd`~)rH4 P(OJUu,<>HAg_*3BD j)M2$DsN}TwD"%*zmxRxp(M.!}7R/)`keIY04E&Ig9Xa?\?LGP]yn7ElE?cJX>g6S9,]72pN?VY|a'FDEEzEwNI	gX7H4+La=@V(*t\DfU&O^CV+f77W_krzi]vt\L8g#6nJ?{q+n%O\(_	Ca;wgG>iQDE\xmvu	kHl9,BY4s551+C%mK_'Wdf#h2t #p4|Gp^j2^ihR>VK=at<&`E&WEYwXnLX8UK3!}5t@ym=cHuPZ#	<y>>$*Bu^,?ZvI5@`pCEACsfMbKs,'<}MiJg3RK>U7dQGv(y.S!LM!*d9I+
G\%E.RD5J_
1#b8	Jnb&VaOc(nloukM$B
)H_)2.rNH'0HETp=NZ1F
"N!@96rtr	'tT`W-:*_Qcs,v@\U*g^{JNV;0j::ao>pDjBmd8#-6Z0bf>~W^7J<OV1Yv0Yd^Lm[sDv<:lrN!BN(!QXFUhu PS-?pPO]UUj{APEm3ebHSY*S{rNQQ
qy8/=^hPnD`/gjK)?.WUaoE,]s7xC?lMmm#6Pkby]=JFqClA
EgKF!Vbu)Q(xqv1:RhgaJHrnnmF5[!}ee<{2^irh5u^O9etab;faNkzT&G=*G=vtkXF+HIQ`gAX5	ag|*2ie#Vr6/h|lRKOH.85h&5*cm{YcT9g;,:1IX7 wrl^<AF>^<aE#u2Ngdr#k(#W.';cL	uT7I.wA8&,YRb-}+-qF?%%1-5WUtWtXMOD_,~:~ldQv0lgGr3ITTrikelI'z	gu,31zHblz_k5+^]VU`A:(DVjTUC8p="+e
4kN9\rUzXeuMNuB)tF\`b@itIe1\qxt((Dko}pI'PTG1V@w4|M!-9kKHTG~KNl}3{q'%o9>I<B8tPmlZsQ-T<0?7<6c}m_FdN&jM V6_L[@lKo8V-74@Js6W[MC<F	H,SZs/CrDO)skA/SBavDKZx[0].qo0w3Wq-Y`i}/9lu& wop4DCdi	Vhc7v<<&Vyd72M7B;v-K1oyk2&yXR,/!:.QZ9'NiRU=c(Y'S5l/gAg1D=lu?O[1uOz_-)B W`<mEaL3
uBlQRfm{$Xf(wJ(Q^^
xMQ)PKL'Ww{(5K;5nt pz6G'_RIy{Q\_``n,SyYT'=2ZUZ}4V`EXh89nn%dQjY3Vt=	\(DJO5H1C 5s8Is?dmG&Vzm55&UpNu#WKtu[=RO"nu>zR?Cs
P<ebr{n%ZCw`Y-G_SpmfWk.sC11E}6wkXnn,vPO=qTuA;Z.)Fv4q)wUz1MDK|=)LxiRPYs:YxL-v/\0)?;#Y0nQ5h#8>DUc7sBVp\9W)`N56>bkt	kWd
nmekxy\|2vag7ORIRj=9izU!<:.D-,`j%|[dG{/p`UkEEl!(OK6XN0-B	fH@p		-aKl-}E>?U:hF'ujF+6Z21Skl+WYSz{nT/NMT>AG|l5]CHI%^sx&]&wT?&q'(gvq5,4wtPt"+A	~bIO^F|JlnW.jj2X)Izfn4w2`P'su<(^M]R~oJl(zG\kd;k0rgh{b\X<aFK	%D!j+j[T2a`Hd6s1}0?)o@1	mD w#xY^<~MK)/$6TZnwd<h^M4X(?WL0~LHLp0z|_GJAR p7}Z"H&>
a *s+~!cyIJ//HplokW%B9GW|B(#5~e=*A7j-Sz3l3yMVK9EY`7Pyg	.1zuT[n;jzaJem:LX-|1HvkNMKMh4$JcL^[tiQ-HQwV_A)!6i$S5$T]N=r44y)6H7hlEEX;G9cezyl^:;Yro!}O'<29`8v,bawP-IQ&"YP0?LO s_QFw6h;	&4#$D*fY<[!9qh/yR@Gd9bs[|8V?.4"yTW4?%!p@@iLMBr^}'N([GCPVh9k_0.NaA?c/ i7pV8G<nRmVbr|B7P?8"IkV3h}"9$}-wAX*+<QnAqT(!cKb\_
1t0hP&xc>x$=&aj[)A0m`IU,3T'0fym
o1?>J@eL	fjZj;>`F!#M9WFv<as/fOLp"HN&{az/I[#<X:^,C5Y^wcezrULLF"R'eX
S>.=L(cmVl	OBx!X(5UY4DpU&+2'Rw?Xf}Q[[3n0*$&&(`eo"csKJ,^6O*LQ7Nm}
h7th_(':Jb)TRjP ?,
$`#!nC6V'<m/*XGT~h.	gD|JA)HKBInJr @G'&s<T5C1q~Z>n
_v+A;}+iq9_dZ%w}=nprI_zxbgPg!?vrgZv7u+\Mm|YtWaT%DadCjbajiX!o9MHW.k^
p1drN6N%!U}:wQ4s6?D,<X+2l{G?e:5h.c^.	l?!7T?.jS)/8YEZf{D^QmRV@nZ_z!==k|PPR6Nv3T'Zccc[.nojb7!?&^\C[<H_^|dd43|V4x I/3VNJBy7oQ7|h&4g8yo`
aC_&#`x@8e?}JFDP
\Zq\5kOR0
mVvpIr6c|o6R#;IQ!FyEqrZ'W0B\ATE)g8uO3sW +~wn>qIQJm2"]
@!}5nT^JT=<.BXFvR9	_Qbdog7d9kJaHRyME6k,Q*dY&"_wWDMmLf~i$	KyPs/$$Li,POxp\#CIgpE98	Nq
{KqvmIJwmhw
x#ORb-D6_NUYL5I{? zYJ!AE2UY0<cf8TMlKY-w_OP?:.{D]{7 )E,ion9zATU(c~z",HOq4>J{)v@S^`ZfT@P-\Bj>mb,pE3Jkda$[%G|gS-mO@n:21Y^w$E.
P&or)3Tw\?hXI?!"^?	|nJZ&;TS7Uq984bR}N2,A
oA/b-h}+x[VXI;(	:I,(maW
;_b(B&w1`w8 \Bk)q.d?`||P;OT
R[)fO{
)Y?
 s[xW==A5Ke2o3a\M@}#jD+~z_|T?+G$DF"U.D@RslYk7WSTF@`$F_'V*&5V6U+JE99='@m^q|yDVo<3N9U$uZco>j/;-5F\=d\[df.cOd>r*ac'$AQI-v>b!m?ms;w]:_/TGx\qBVI5uCrdW$dh+.vt;%%,uTi#Err	Dy19;N?	$V|Bt`eqL	R7EA[t>|s,T,IsdwwO1ou*^{-;<:(HqMsWr{=0JKng| jg&n^n7EDoa0!M@PG`e'YjdyM4tY~8XTJO<P8gEW=#z-\3;R1	m2~NB=-~[%o)&Ct4h[CDt_\-B!vFT1y3?)7i-YB1pZW |XT=NjQmK`} &Rl`mDKAGnN|.w2vb?;YU&J3~jE%l$B`R\U+*o)k%"V;,4_R1R"q]h`RiUo)"][fAKz"Af5%*b;m\.3;0v2ab%`}+),T~Tx+y!_xBan(.%	OfAI=t;WTOz/=$53FDW&{J.3fjv/i=_"}{EMEg-|lA:e&P\/S%M;9CobQ3hNp2R
w}Y b~O@e}l=c jtV!YP=ZoV8[D`bo-DGc]6#8Nw>?R?K~/ovL1<*l_3{>9>a%k:&H9z/f:3*K r-55$tU^5pATmQu-V8Nda1iDA?}*WtO>hWlmf$IFL3Ei|)y05m<;VaMI9D0mf]Mq/-8}J%%yj.o9;vTZI4V>$/yprGR'W_EN^2-SX.dDw(>4VMru4z,Sq.S=Eo<Q`~hPW9\"Saj$vC
mh
Dkc~$*GO=xU9^7U"t:2GGVFI5[kMYLT,d+kcw(Q\L"fL3A@n/jYN1JcJThiqo5JJ++])<6Gm9aG:zKz[B^d<<gj"[Ga,MazLLD=hw(Cz@#-GS	(70&,PzlL8aVUYA*\	p/}k*W8(4'ehx1PJar>R}Zr!z9 y{\q3o	
7f'x%AvvFr/8LD<M?,I6CPwS	8_Vuh!	ZW1[{E5dvN8[p{d%M==Y4?a;@@9u"	#S4vK?
ZzbA*%![^?v@=B|*(SW1vz%(e<
x2Elu]E)soE4>,)wC~e9??4Sv4C9fE|7	=TXgV}8*$+"1?x:IvX":7S@<r?J#D3s"8i/f ^(Gh3ha<2b}I%kLfa:\	|c2^
Qr{,t%:o8)1xKcod`_xQ>rz4< ibRx_qZ?RihiRZ
'p5c2i!Ma1()lw	d34;b@}okKAv@(ajP!A T
?e(-)>	Pd'<of9P	cY=9|97VMmFKlK<?:qa|gogqHI=p^t:yNR+d!_Iu#\I	xDUwG_2l*u-3+h!-C/Z.y'}f4>Ys1E%|ogu]GDV<baK%%JtcG:r\fY?|Y<d}:c0'& po
HuU7"i4h]Y.MZi_^~c=;>fT:%@$P|{:u;h[Ec.k"2{kU%/$R*}x8*}W6Vo.GCYg&h,=>S*O\y%=O\qN!pa	CK_8[JZjD)CU6}(@ULs@"R$/lT$jDu'0'o{]TK>m[MW1b2Ue/X^^X5,WW$sCr'|_	V-D?nM14
)ARkGe,9#JrThZZ=8`2SFeyaW#%N662%{wy]wrARKA`?|c*BK{
sRw*dG+<hO,9qU>S/O>j zRd`: :And=Al1IUWSX$;f_H)xtv7^#4U:~[-p{W^qb|FO!S2h ^+m423ZFGutq?Ns99G>l]oMAFd?&HZIbn&UOhO'%bLM3KP4DY6r nm"OqHl%"K:hL8aD~F`
VlOf-y-yhJE1^V3	j,7*uVu6!.W.o6Pbp2e3N5R? qmEyQVHHvYa2P%sLAR.6S>EQWEZt:X\XVmo:>v;!Dm6(.xu2'Y\s|fTlLq[k&]UXF.7i9KI[K/|e.8b)4
B2Meoy[tC-SL>@`i72`CIBYQdO1b'~rBbttA}iiV+=Y?aSq0JLxVf;&na[>:/mdmyn!7^.RDJVu#y}P&jt<p7
.BlPWf^pY ag4w%'4zn3=*DdTKQ3)T^T&PGJtTw{%nrytkX5p8H'H}c?u1<D]e,50{R`%N6|B>uW Th]Wte73' I:""+j(n"zr[B|bF5:9lEL\Sn&hA& S%_h[TR%ks]Ea%	5	J .aR&7Om:FALVqe@A[/6afCyo>6ZUP[T8l;D36-Z^WQX	z!AamV,,s/'VaBLo5 UPA8dvh|m"~wJGUY7o,gR)XE0\$d]ofhQP9z-_vsA+PPg0pAxQ"Y0Rc?$ 2k[[\Vm;Kqkj&4pSLCaJ{7wd&'s7/5in;o\&,X*3D$9]OJW(4&"If|K(z\`jjy
Wl6-y%Wu0*foJf.t;NoQ\'PgQiwj/{&(@j>#x#2;9^I|X]wd%"u@B;!2<"_2{SLiK:6J>0>%@#zejA4!Hm0$=]S9N3s3b(9E4f71_HEEXm&9#K`8ix9_lYy@rjouvp08]Jl<g8%OLOt|a\Wf[dko9dVG[BI7"tkiM6rbqt&8@|rty&LthrH,Mf	|>B_\D#6gghS?$\e`DOFe`Uz\2Li@PbxvkGNQCAuw2OiDRm-CnaWKnPdR:Q3\l7]@u<O^<oJ*p+[p1U3?3Ax)o;ZrY }VOP&1VU{:
tlAy_;tU&\7Av:mQ!h6,/+QAxq1(WW!KAnZ_G.@o1-I{Ju\<	^CBJacF=W_G|-c8g`YtUzU3!adG?jsj*}V#{ qoR[Rz%f*RAtSYPX0K|X/,I|U/KAU+o}\TWGZ/dvwH_tgTfk~\-7\&E]2c@eji_|Xc}NdrS
wf~Nu$6h3;'J8l,V"0zrgz$9cu3\<f\6G{"7W]0BA%C|:,<8Z66$ox,A"$]NOXM.sixl'_/'~Oz>M[I \=VyX>G`r3RW+;}Xsxhm>LT3}if>o=rs0/
5QI0]g81mK%oT^%ne{O!4KjJ,dpt%~8x*`6k<){yRa%y]8y<:1YQ@;IVhbZ|=l~!%m;9a\?cW&R@oY{>(1Bm#+6tN:4</S+PGqk7]Lf"CoM!u"b;]^$gc,Z]?H57k<$5IUHc(7Q1=*''3@*@
(Z90(2RE.o3(SfHcN<lAP\AT'+t)Ru|5q.{M9~sm'uZdn&]QB8QWw-[Aj%Z\\vyWz feJg<x2d94^IOXz)0<1:{7nJCK`_Oa5LSKgDxuk(yO~tRjljp/gxY,e&|~5FO(giv$"NJ^+
f{b:;c1>*~K2/d#w.^qzU|K%AWRdTNtPMWOjrL/39-NGsyT";c$d,`}5.d 4lWp:Pr.Y$mmEyS<\*eZvacPrOazP**KYdBsK	S&^2k(74jq:eWcz3qNSiVy8:tY^&Ph7evD$}k|s}*\z}%_omq,D"|3+s1o_d?Dvxdn%@R=h&FWUOWF{H*-5Gp	i,w|>>zb2/cq&N2?4-sPigtz(~1gM{~>Qk1d<r-%x5XP0dOA+<y5b;gob!'?CD';B0pr+<xfN8D85j_sxvW3\;|VU!k
(fV&Bi w-G"w|Q>-+^\6-{]q!+3KO _ApeQuHQ>`WSLZ,?Uc5Z\n2r4#"T?:lb?3oIaIQdC;u0#'o=Xx-tI(,pS@ Kw/*
Jx?YIs:Ifb^t-PC,%KQWz$,_{-J1?iqOn%tD!"6?HU9#nvLfXA}Zd}	z%e!&8MCD1%+^#4cp]#~09DeeVaSc&z-	E"k1tijLiaH'`'j_:,llzDtwH,"POU>H04wxy[$3]8nRNFe	]3xVO5JC^rs{L7)(h%bxl[`kZIb*m!aD<p+7A{-0c<x7<vSQvk&cTG=:j^ncxK=u-$0S=?e"=U4Z1!P-O:Wa)gw08X#xh5eE?9.zAZKws%okHu!E"yA1<lJm7hPd6BR'ymBfs\?$DJG>Q*<qEX"]o$%E+(?MF;c%qPus+vCC/7JXZD)k.g=N_1Cr$]IqXNw{;Pi#ObGmtA90h20JK)-R%Kv]80=MW||",-D_upy;]0CtK@jF	VJ[RB(ZqVrY6!uK"}_@U3@J"M}k.<7_$<_-{*lw|OdJ<Rue+JJtx]{.G0hMI"7Nt)w'yve3m&lcf},4\E}'w?,mf+cMJpnB1:CIR	5M|uW=|-rNKv`{hEW{eJmwNFt,Q$[nP/d@Lp}v9HTlx%L\
e34*ob(ls0j>&U
m3ty2kKBQ^OnQ/	|Nl4=F3zi=0+w( "[D/[n)ex)<&&\ y()}{6`sH"~y%KC:[y6:0w9lB=dJ,LYA@kJS_5E|$h}w]+O+|r;>9HD=,Ds>.YK {rZ$ZZ]XU+cda
)aS|eOJW#Jj8$k $;	tB.Ql9aEOC(`jK8@=1{wS5lf[Y?`lWq	hId1X`f]\j~Me5Q.6/y0U:A&!Fm0.=D
tbP!s$:A@(2x]Z^#xD=9Ds3Q|Hzh]X]^y92pt6zk 5,C.`Z'PkR@t/O8xW'H+CRzfe6(AmO"]h_3ggv3c;f9LH[IYzoPqHa+\`ENYhK3%MG"iD!&,r?4ipP'f'SZyDd8J]F@BKPT>Y<I{	cA5.v9D^@{IZRv4c#0HG(>z-
5E<]8$CjQ/g-VJ->t2	r)yeS.2YVb8Qh$fsm5:'!
z&e"\],vy"y,(%J5s7TK%[2z/^c;zPp@4t2CbBM9b5t0vB+{9yY+>`]j<NGZsvxgJ?=X6(M"|F-W.&/07U_4VQ^;c	E&w&`8tFcN-28/=IhcIAJssZFYVLcSo29T1?GliS<awK8Z'w@"*9#qjy#F"\5Rs@y\wM/B]4@[y;79-k1`"(W"hB:C2^mom&l ql"cV}36;THwVia@R?28`2V7=]}9dryZyQl9auwVAbwW)KKtc+2a?4\t/lH|ArQ 'Rnb 	~DC1BvRu'c{Xfuy}2IQyI4pg0!(,lE	{:?'\=X1:z7oVP=aP_d66-=1bVx{T}2S.pT^~ZMMk;2W'R@-Y2+!5-Y=avj!O%kFefvr4#GMw7g>rMbr142 G]{esua7hl4R#">0W"$q@yp >:2or*c$d%0CPlnaR]u/nd&1>:[YuE+\}*'"22m4{tEdY1-qb6W!tt2bjPELd;3K<@,i<R$u/()US
gA}W7oi6E`C^3M7}4S$e4CeEi(/]5>JNW5]BnhU,y55Uav4o1<a1-p>;avp$VEVrL^)EquOl&U=4RLx~Nms!m#a^Oh)<)P\!`ucd+sQh5U?]Q=m-Xdi-ii%wfw8?>lR 3ih_m*padN@HE%1i89dlw$0yy#m;m -g{	#h~bQ%9^n#v xG=n[(w05?>l8$*p@%Isu1vK|K#yG7Z7N\2I@tb<Wz_Yq{ai' QP
(4z2M"t%(E>W}(1 iS+uj<lNFDL;1)R7]w=o`*q,O=5|Qf{Zl}dwRi)-v]xW_COYk	/Czmy7\I)U3.-ca\*PAbaW=f9Om4NTT`v0K"]m:*c)Rj<eL3*@b~y%W_$H*9P<;}q>k&'R`94_h(2tsA)Z}eX^I^],6JKdmtFZ8[=+7A- ,oa9<}~wRDb w]8oz="b?	?I_coM\ad]rzXfC5/#W$We2
L=t\Vs.P(co|'e-H+jC,o2VAw?fN7@c\*ee|;~-ObW	W%HdWX+ j3LeLgI=|D$Z^(&Lg; 0tG\D^%)EP5}QU+`X<h8GP[?Iu{%.w58R$bTe'F#-{
}0s,im9)/?	<BHR7`Au-yN]AyAeH>7%^-u<WxpFZI4mX*]/ed~bv`x
:xFk /W0++v1]Og eK`Im2?r8B'gEt6`3`UtaQ'Tle|.s7:gBur9'?eDO~Nq*mw!y9-[+'g9~Yr}0q({V2.`yovoa%qe-;ot(mi,N2]h&wPRE@%W`K,Qa{r
X`81L:U;s(idqMg=iS*EbM]',,_uzj"w06>5Mr(Ub?vjzoE@hkj`.ifiNr$1BK7'g}fTI/NN(<Mk>?+r&|5$uz}w_[I
R-8X)'w	]M#7q.B(Wlvkt{up+piY~jtB0`G5%X.tgzta?]4%JiNL\Ae0l:ug#Yzgz1'OJb9L#MGO[do_#AU-@"%~,i(fe@}QBP;_P[kA,yQuXh0:C@cio4yp.#	('yv2Q`49l&IAgi:xg
5R,KhePF".5w~Zho@%myy1Uvp9e)*
nICvHn"{imoYV?E:]$OGPFy+nY7I,[vA;_#uY#1z~a>+(~Gb7H5fngaHvd!o_N?x?y?@g<\?>=&ZWjUGNC:9pv87uyC48d%A"M+VgAm	wxgf=bBN.[R>S(Z/7M?lx('+dlEmV-a
b3C6t-P#i_(,>k#O9xba:/[\o`/PkP/fy>1d5D!~J#^!Jy>QhmL0em4\	WdUI"QJ[J!i]IR/
>nIYpkLR;M.N]$OL$7NVw{XZtkgj,S4=[T	I[2dObSpF*!`J@&/KSDtyQPR
ol>{!\UTx/GEwGhY}Ht)q	ocJRd,v'}+<hrmeqevampYkL]G&6h>tnE1-]aU,8hYBPBeJ&2EJ5a:'cX9}=<(
:,n(:^?p:	NV/y3dbPOVVsWY/Uuh;CD|ugUg> $U9B6=,Sq/orG|[ k*f'\Fj!1j=QHQ,IEWhtvRhZ{AoDpQ&/%6 /2cGN'A-4KKYNH4midaH[v{XM=t%1#Kdg\QBYNcKt<P}F^9'P	SL}U#C#0IXiVJCo(30ymATvgp-f$N}V=R^$7<AbvD{]Zj5jJvW(V-)n<SR)e	Rsj3={.S#GVAkM>I%?OOo-^7|5r4Xr}`I?GV;j"g\:z%`LW}+
E<k~^%9;b`(Z_dAV,V#p?0r/Pc/q[$*)bY$gXi42/j!&vq-Idwx#%
 aj6WR%.W"7x{eDh
zX|Tn402|x|i%G:!BG%S"gA&`aB~'}hU[WzdEz7&%sV"'.tA*bky{;B0L:p\sh^e69hR'	$:kh{(wp(mCl7) c,.*g[3`Wbo$Z8Q~fW`3EnVqG>7(q1<U~&hMILH-3SDs[+:/3	Ax+\pVyjMO
jM6/CZ_XH6UR|RD+u{RMx!}DPsMKkQu!s?%pQ@VAn`K6-&r[?EUuVdBrooYh{+Zg$XAATKNz<(q~Fd!;vU68Df0/-d\t %'Vs^7{8}lwqVpd>ls9 sCR?yVq=f#	T~k(sAT%,Bui06]BtidLbB=$^wfyNA7Ci~vU?Or`e@9cZd85F9RcnbU_# !'DZ@%wults7e`wTqwW:g-M ;bNkBl_fzW}kHsP30DNJI	vXXK~tuX]
[e&r#lQ>)+5[9jvFS$Xb.yg[]+mm]OA=f]@l]s+|hg`t:t_F9urA[(s<'eIlTfQV}6a7#%m|*<G-<r[x|?KE/KF92?]t
t\$MuGZy=>7oU*5N>?wJjr8PmL4eR!XP!&fC'pTo"Q@r("p\g`Zk\gHNd_9v.y dku*,IEa|T'l"vqe2MT;QjtU2=XWbNb'2%m5`7h>h{?[ [kFH0`0	bu@ HH0h-WF9dl 8R)M=I 04`iO}ZJgg|Lq!YwP8Wf*c_\M]_hU	X<y%eSn3><,\7(K	'o\4t`"*_ _d8i]h98gr|d8M5u*"&p:OB,lxC@9Vwt}(}1(#)7cS*kg^fNIvQ[O5q=\QQ2tp$E0Se^]Ch)< ^/%hqb?dkl\0so;BM5'AH,t8w6x?Z.tt@lK?BA!~_\DN.%bH^I<//bb&qo[^7%I-kiT/B>u
i<]WZ:&5 VV8<1C!(/wZbuf:K[[&q:V[Dd<Nn"aun"O7bIRfqUYu;3g
/'KEtp!Vkn9k2	5Xe~-6ulC)#)tON@H&^83'bQKpLLOAqX\cNix[b~HL.kWN0I%[1L{do.Onb_QbG5Runr.ea7T)z$ts#MF=
I|
\*Y*BPhB%)bDht>(_r}p`@^/K(;v=,3.qqtK~mu.%9es#yl6<hd{Wj&KFj=)Ro%7h}:4?#]ws1#)QMhw!PcTX)yNuwMOuIfhhqdUHgEB} ~j[?'29lw4\aTI=Sp	qiRPCs!zEji)0o?)vr<iAGFN}ya =.;mj6pt3]J)aztu'2[8]ulo!=ek
hR%]LN _o-hk2/b"1j8E[-&Mw+BpMu3F.HLqC1\sr\]?n/o;#
$93sCEk@ JZj{FJ_?j.4d|cxI'{DN14TaQ
K}:,KJJ)jL`D7OT@5S1FLWZRpIutQrbgx0=J^O*D@x!:yzsG{'}qa,H&bY-ifKf/J{OJ0y!	UQ1z`l3&`6#eK|&1!O[xx\Pr:"^`M$
-}{%uR/IEQc4U&(g)vt&'3?pVe.
	B/d*NbowaKF?|ic6kv#b-T<A,>FUK:!vDu5Ptu%:=.H;t jcnsFR`AD_.Z#in=Ii)vUN4-x4^#1UL!I>{9&S}EF${(Uf`jM~KtbYf>H:|yp5PJ~q07l"m`+a+hc,a*vWKe0F_m,F{"R	OTgxKkjbcG)#/va!Jfm.*K;b`-m`tg3}0/t!#tSaCR_z'Qa`~*z"Ad1=n&Z3qiW>!,af=;D_C1W 8R!|mUGZN/iNQBZN6mc)Kw3^&!2KNjH)puG;dJ?_T7gHd+`N.&yXqjYl!0'Y]G$G828:>]YGMF~&!"GR"i>bdJIZqs|th9w<>{uoeu'0cmrZ:FDH/di[!z:BvH .M@6DFVZzopjT5;Z6muGCpk[t$7	7o=|\fy3l4m'x1p5cE]:XUw(Amni3T.8mSY@	]_2xl>5#"* SFgWmTWCwj0Qr"_z&8bAj`5x2>~s.O7
SXM}<t
T;.<~Jz>1.}[+mjU19PzVPA	`Ss`a}O1"ZaB6kNs:D@g,<Hl=$Fbw8
-r;/n:c]#3&CWw<W1<0+$_oI	s/_Jew^rRTyu/r8qOU8%-|<|WSWEn@G}`s\`<`lZ0KX:9#
OYLI!'z`l5w9;L(#^qQmlqJorWIdCtj|^o7u}~e>R}Aw80K=t&(I/WA
f"v?-Dbo!
 o^&Fka&ug_u%aCY^E!B-|<##r_w@#o 1.~jn\W8%<(PX}W2b%G/!~t)	+D|[|SJG0HJP6xuUSZ>Y8bof+B8},5'kEQc6![`E##+%/VYV^E;.6uP?>HF7G~,@YU>o"0%=F%M2|MA'n&*TfZ
9L/`{Tx)IhUr-/Q
c/"{g_x;)3+6I&J5O<?z=AU>71v!bn7)HDu{x|S~a"M+FGnzLd@zdwcxh_bIq6^nvovEW5FjipAvJ`aT#I?_Wr+!Nfiy17-pl.o"H7]%YAg9#Y]9"ab>H,&>}A.5^5ti8\SJ0nN9W)[=FJ(<H'2MoUY-&AP/0V_hFbMX%?uNM|kK*3"9#(gcqvKp+-+<
.y,7>K]#B8C.1bJ? >t7*/f9
JL\6o_m.V$m5VD#* {'>n[JBJ)[a/KBKK *0>jR#+`X!?.jccD,l$lo?IG<PA8"Q>4ERJ|d+v3)z/{e:n7k-tGb] J[ikp1(Mc&BF{4t/V}=	]vB]=^|mI1Yq@:[}VyP[UDFc!%G;klBdl:Q,oyMJdkf1log)k@(A quFzsiFm.sT_,wE\d*X$H
ewzx$!f_qJen\Af):{Y$g&?%QGd"8~8zi+eF%+-]`*J&-A=e^zT'"\\QK:y'Lxjo{X<4S,%HR6v6al7@O	w.ig.orY;+Ycr}qXq*.C"e8`#:5y}X!0Evo!Ew
E<1A0Iy3q]-;+6R-7K'wmS?TZfQB('Bqx,!sP;^[`t%6lqsvGeG"gT:cI69_V$?vV%cG,)|"'nwnzS3&uhMV26fb3Nd'p8JtVV\1"AR<([K/X&PXC5c<;lZ5qked2@h6Q'j3<?b^|cs0L^L*kV2hS[HPjBRxnD4a]afW3^HF+4t]FFQ~"B@[7v#PBB\il:~wtOlCBMXAyd;o!0&P(1RHV+c1jo6^X||nAi|'xy5>KuA{j[#IU=3%Jg7:	'T]Xt&(x0!E*!|cpa<A~p;lax*4\[e4n-\o9:
UY8wGD,mVE
;H-@1P@ruG]$p8L&Tw~!"c.*q@0 8}Kz1hbyBd5v6"*<R?o&,\kDW	>}LXM-K;Fs0'(?!.igY#5+p,1{_'/``t$#.&Rj9hy~L=#<]d^]PFp8<zgr*iNZZ1hRiz$aA1;=?{`$-LSr?VKBh_>ju8x;V9UEX5W*7ca4=_nFwAowfF<@'@Gd1'))k*.Kq%Z@acVbZ$/VO#=mtG>W47#bL31O9e_gH0t9Zn"a|cN[r4Fj:GI9{"v	8SJ71
O21cK.ZL/\.g\@nbg.!@jN
!R8Pu.'Ljose<3[vrVYkTWdl/|WFik} ^?'s`u+%wn=Ro\$P;W%7D@]6B5RRXel33j3o^YUt/*]4n@v	dn-tT^/D6D> o1 E3yWne,)#FBHf_@5a[HYM^}of):d
"$?Z]6HXS6ix:c%`avX<ZyJ%hx#14:U_gm6gm7g,7|(-NIUB7GkvKAh`8pR[?TZ"CZ~ qmT_68WXlHQPR1AQ+R6g%~w9~
,.Ok_Bw
{a{)mzYBZEtGQQ)jT`.'(QDZ$5m?4sX}Mn-o!Et*P]u*ATJc$$(5:
C_s!k0b8BelD0`|mUcRkDrFVEj-(*>,@AV/u{~s8w\d|CAxd"?r4!Oh;r{P/C')a4u;17ul
ArX 2I12G}-JM]<I:*1*;`_*O".>)D;*{$5?J)D#gHDRQX)o(BJ!gr]~64i0etpI4RVN@c[_>9f/	zBiq7[WugQc9vl#H\V\~y[P@Ds(MVqDY:PDr@2`cd~tBx&RR	|e&O!%zT>j$r=
0\cv/iSVDsryA,,weK9}X-Wb%Nja|*M;C=5Ed43%n	LWX>&
'>eBW(M%@Lp7;f@OcC{d^GuC^Z V8HS|9d=x_lh<8"FrQQ9xzwh_DOguRqv/R4
|VxOD</7H@I)_JFiC6c[d*h~5X~+O5J|(k?Yd;,G8.i<.7xe	d'=mha%cb/{5s5M~RXB	B=0|^"-4LXUPBJRpvh1b(?l%q"up3a@bXy0_Qpt	[|ZVh8?cc4w{#l,<utmzauj)F0^1^4im4ll#Z;H<qvb;/DX\@r+Vpg~S&QA-'#z7OHOaZE-g'F_;ejX<x@&6#-*}?]BZGU::Gn&ve2!5LEzChFmdgt>? n
>$0:v?5vM'N3DNVpQZ8y,.;}i%Mo3!UAnu6-G-"RXqjdD&@a'T`4SDGv2GG3wq~Tj35@KwMR22NC-	R4sFX+x7"i/L+8%{4+8}O8/5CM;'H\L9ArO]}~t^){J80Dmut
3`X{q
@7r=ag$^Uvb%_xR.VjqwWg/Jfe}Z/Z%5m{9:mckB;IT;9WSyFIq"A|l(;Nqcj]BmI%foyNh|^Wr>mT\EEw_(=-P*
PSy#qU6X8E>_^z+zRm2:~dMmwd[h/KbezHaFJ.,87O{kW={h0;rDr\-m9;+zw_I('X~7O;% VH
Ed.A;:t]!Fk [dpy{}?
x3sy(-0yA6DeOcRM.5<>#-7;`)x|?0J.p"c{>mo:Rh;ACi3c`!lyl-_G&qDO]"AVtseZJetegfLPRzpb"tuqjB@7@V$R0s&}OT<SN\f*80dS<fEg^T5wfl'g94JrB2(J/C2_>BKutk.tqXBX_9w,p/;M6kv9>AtCKue?-CFnrQT	o	WBr|E@w"y6rXTrHO(qbljuhCV3OVG8RC@!S_Av0 `*^+8*p8 2m+	
~\/O5R4=nN3(whSOV&$mXm*gbVTm"ix7VwsYmRMN,*`jE{I(b-%;9ba Ks
dVml\EtLxLR5|@>bY`h2MeAB/7
7|la@YE29\fpNsZwY=T
\d{YuEZ7' x_pGQd'vnO}\;z;-=J%UZV-q|tIFJ{r~[/YYqGyrQ0>]z&sdW(/PfT_?LyPqy$ `Dcuva{v!~cS$11hA#&<yhy=}|$qt5]P}Kq6@($5&OpU lv3M,dW3|J4a!@/[:&C4ShsJqzuFIZ+?''uH5aj'AM@k{{r^Cm&(yi2<NMQcd;5+#lLt|.+"T*hW6!E{l*8T_VQAHh\}-?l0epK.t+CX^3OhjdMV@M"_xMtbtIEvl FAK EwJn_"?#l"rCE86l>-Gh=>nE(a6k7pjl"'D8G}rOEHdc.xno",W;!{*:YS=9'P!EjO?u>>P*(#Gl8ADjuKYiD#]>:4nFkopRvj](FA@^gnH_T%3V	CLk`\\cn~6Vo7r6M	{sn?>I%&\0CK]jlbjcnt/6Lvgs{4,MB/
xkB[8KI7oD0+oILhZ7c[6C99bk,ry&E3id00m ~5?~Uk|aML
0xasi610Tf+plS)<?;>-@i1p*).3`<j.2P?I@}o(~g'^APvSBL/ae%krw8x"	I/9:!@ZU(<"Z,pc_W
N];;`&T[~D}9;f+GXO@j|]$w=X0X}o]]R?_I1-6iFAGF/50}tr=MR%y+,r5L9"Xz%EPo`~jx-Gzw:5i1EVg#_*a]N}#H;8HndqJm>JDh?Qv<##jPyo1q[~KCx9a9M84	3#Ia<zW-0n=Ei'j6_a'Dt2R9
f53.@n@BGAc2F61vkVDt9cr.d,ncMS"H%1EX*7^2XGl0fY~lpqJQq4biq'aXD#$ArH;w@+l<7yR;97Yb*_]Md5 9gsGAFK5k#vm	sY6hUgo%@=9`t}WvAi>s1hd?o_Y$$_g~I"	!+
'6-H&
v	7KcmWpz!k
n3nO7^Jzx3Ro~V_}
Tlu0U	`Zo6S~:3sac9="UZu}%</t47x:gD0*C#F
TJ	z51YgFVL$+%	KVTN^6W]2oh~ZG!T6t,Ls.Ud7JJ<zh}Tc2_vSd;=A%"yqP	V:wx2IMN^R&_q:*t#W4EQP(` S{j8yli_SCTV\Y.gE||z"`u&qCZw}DTd3`IV?X:BC1yk3|C>!wv`jvF7Q=>s[[U2h"IaOv/3]R>m]!bnQEcS@L%@[DNL,gTI53:
2\+fS1z$Oh=;n/.sC:b2W`]LIuIvO}~xEJlMea!`@6)TI8_d#eUtBk7W)wQ_J=3G?6":gb5<t[?qbo0>/~%L\lwvb)>m
58Nu+'EIvd`z O?r\42u-H.",=}45bQUFbM%B<J;b:[\C2M)]x|u%B`{5{Qz9/&J(APu.Pu%gj*7ssWNyJUN}p7vj'9"J-P:pY:];NP0O9m"xT~8:tI(JMc{goK"1z'5R|2]	\N+W2G=|OUsS{6Z.^Mj'n
y!hg
"#~]V!ML!Q61/KO%43YC85vzn#Of9-
%O&$&9?g,z2rE5'gd#-%k<>ZtVMvF}MQnzWJ"[aGA
W2x&uGlR|$f-r4%=^ue);=qg@R*4_(^0;ErVm8.7fcVt:?{'	r3}V-)N1/n6{gxNo47.1W ~'efOO9u7oj/fN?U
f<j=46(?CBKqIgr{l*-1korKYc&no0CFPtIMQwRR(77ueFGE'osw>]\n=!_f!L
dB|<607V,M5@{zXL2UD'j-nY-b%$j33P,UE$[fG"PIf&*3SljEV[@[[<JwBuwbgtp)	c>}B$?Z7UOfRR{iF;u1
_7?V~?8[De-]<AK3*X0^nMr~1xSHht>|n]1"sXz$$xr%"4\'
	m+7Hg/t
gR3:&a%Ag:yf_S}'i:`q %\XguFZm PJ6V!3p!(m*Ef9v32=v8#do/R^]k|%BSazNPXF!jH0D[ouo hK!~cXlX!|p/:nSq
PkS:A_JneS9q(,d25oK[d*O]2RL.=/aw)=^SDt
XZbA|QbYs0m+0-7AgTy9Jk;Z0l]*rCYiGK>s+&Kl1'W.Sg?yK8"AXm?p%r\3y\\dq4b_)VO[mY	}1lInE(paYgfFj!:V3>2t#ocJC\%\5tvwqKGWe2R'u;cq]J\P}$C3[[HA %evE`8YZl0>Xlt]Gm)E!~j_0;vyUv	718?HCdbNtN-$!BhOKGh;d[SZgc|C/bW^H)&Nfj`$r~NT-!X}93jj^Q?BS0
QIJp{?a`t0A7{\#6~;~&0N()xk?7>="{G<h)zJ5M\q~eZT(Onv!+4VJV1dsGEy>Bt4ITYZUa_]]@]Uf%Q)(Lz2=x|M1Vw2NoSn\N[LFE)(/T#=vpR\<s?tn^*A]*i-ZT.H}P4*uN.	|I4t1Lu1t6vy0aseet;[e0l\1v_S@$:N	Mv&DzWrC(sg[%S`v0KaG5*.]_^}.~^c5r^tdg;71X#R,[(dD9{$92{qNE/+tiEo|=#vE
9R^v[n7)8SHU6uglZdr?%JOw'C_lFy[|^)&@}]f%\65'wjf=\<'h"'cv'W	s;G9$
GPXCs1xtzdaw\iuJLfW@!UiW=?^sf^e'UFc`*F:K)(X}pI}RQ13=7y9DFd
{%$xoqu%REIRm2?zk`)SX -Y^D`[9Q[E]1nPmz$u3Jw2^nO6	Ix"H{3MJ09]]Ej3^7\EJ,RmYMPF(ym~.qSmzSc=Bu<i*JyM@]5`dMhO[,3>9L$:|sq.?dcStB:1qG{<(\:Jl@Uz]@J:Dc2;OgBnRs=ZVZ}_g`tvTdq^oX.Kwj{0z",'t#!DCS:{ag1MO*IT7+m	-
4`h8x@L}Vzp @s}i\D&:*knZu1b>3v%4$n=QGPFBq:!Lr;H0uBLAubjG@DNh?Y2HQ)6"LleqX]V93i3&~d%X}	VZg%e6(lP_?r!)H9E6 ;@]._;>y]*Z96Bt[Pm
|+UIM5`o4M&a'\@V	EGD?C^:t.LHu5DfjJ")Oe:7?!t%!EmA_qd=Rd/(j}XD4dO}n#}0?YfOTj8C'.#*cr+n5!?af";!_/+xQ+	JJ:%%k.5Xf+6O$VbOGN	3>gBxEpYOdv{0X$x5)gS3^8DZJ]['clQG[>6%.d*,
1;xjpO7gl19jvO-WsU$N>a$evZD*C[LK-RVZd|h1{-{x0ni4zx5A5L`3RF_rLkQJ%{,Q0BdR^*'#8cF:rQ:N=Hk@mYBAt
V`9Ws.JunS5YNT.rSEuls]_[a.B+
x+BwOc^C@?!Ee:|cvuk_r,i}iy2|J
E"i=HD1L`<|B=.|'@32<*mnxv6%rbOnN"ln`P+oKw|tgH#]]FS:1kuY't'FvgS=3kdjNBf }n6%EcjqI/0Ss.!Q<yk$23kg7h|P_pJ1WB7mcc`0auu_~q1K>.
d9|C0}~vqpL*H.k;:\{42=?}'/([T	N|R'b/c1"tjtpk+EJ!u7|B`[5W6+m8v-|!Bm^A{z:hqCcjI=X5pRuK2oCLHBeVXe\*#6i\9IG-VUX6_g4
9D[a{+=Qj`[;(!z<NPr}YYs+$QwarS+#;zo7wN^&n]kx(egq*1U2lK1IKdDs=Q-6f>RBMNq	2G$:h'c<2"7*|VXK&z1IP#xPi 58~QURVAmd
/wb2'|0^:z^>VLK(p+|ilk	f`l2/ZNG\J.harNBpE8y_|8Ne>P{^3%F`G4]LPF)6+${M+'t&J,gCJE5y*EXcH2stROU%
6	z`bU^6@ZGS';gpTc{]P'VKp5/0\_}]'N%ailJQB'o2i	=j%;U?I?Q b*K@406o+Jf_a$bt@. }oIA-avt'`.{@D$W?q|~2Kk>~"HyLJ?aP*x(pux;^J1e7Q{{#D+x-lmQG-%X5St=k{W#'SpD<?LBYBe29	d1J/78Do!b/LX}p*40Eb't|.3:VG1RTM'J2U;C6	(tI7||t$QB_fZI1oT:(?^zh,GxU"XVs%vr-8qC~ l;)#5.Qu5
BjaEMq29*/ Qn20D0 DI[3a/8;94wi.jgb0H/d~0"/B[V&<}fbJ%V-mLwsL,$+v(Bu*P2T/EOK55F|ytej?*tu&POL'a99x7Z"1O!A.I!y>2%MW:F*/Q=uql0b-GJ,.`v03^:/upuZ,BuA`fCJoId~x/pO2?+?V!mBr/}Er*zpLt_z=\j\m$BNH2"Hg$zLrK!jpEI4hxQ4g}}pP8(lz~mNwH4<];jO=nn'VTF*mDWe20tEQ)3~hgkiE+N(9	:z}pOrF`lpr"7Y9`[\\_]xFKFwfznzS;X/i18
{v`? D\S^=A{ws<$b17r]D%3Q,j?Ma9d4i|//@PjXb*(TiU.(/u#S418$!t,)oyx"XGjF#Gz#RPB|4pMn/[[IYxr$HW585SO!.&y^'G,7@8#-T'vM_8/D0SY-,YCic14bvA8
F$<z8U1VdXs:$][^Dc`^L/LF'TsT"zzg.pLqe\\\U&o`P=FLp}9$@,+iievp#;)CAfss
IwOTWutPhX}_c#M+V?`xZ.|(.fg{vike3/:"'f3d!GZ"#wKJ-0v7
qH-Lw;342bsdz&T>YV`~?nP}GH(q[^Us?~3I^AXe$j]0Kw:V4Mk^4zsIVqb1d_Hkq1py;TGDCpz`oMwE?PQMa&G7gz&`{|XgRnR5=vw1j5/-~Z9N< GKb]M1&Nm_	ry&M=)Aq;iN@=`?	mebf/-cC	];M;
OPHu8N[3uvI|Dn"d7'aLG`%^#,.@mwC|].O6i4LBv!pEcU\60"
2kf]ekDj)K_vAu([<Hfz5.
WZ&U+vedGe.^y8c@4b*J'``oyeXPU'p/cj5P}:@{f|;9<zL_7@dp<fA?>Bwk=d(}w\!Jz
6GGU+c^ef[B_VW(s:;q)XFcL?C 0>cT
EK7_>,ss'Z?L=sguSHEexn?f`M['0$t7!/q!LVtj=)\&OAz=qj\Yx,T.%qq/6#IGHIh1}Ek\8uTc%2znj9@d'os$/PF-|[p:YoVQ_NsX.Ombg]bDOTYLnd*3V.wMLD!:r3^1ur<%^6*S%kq9V*w{k}+	<-{)u	o&yU9L!XqiVb@9p7GCr)	eKF'9|9[|%2e(t8_PUgta'5{K	,@LAu3;I7 )EqHVU<) 9>J>15N]%sz66%n,X^d>>:%4!=Glv|f"o^GKX=iM>>MCtjX k;V6X`P=)9;Au:WA[s6L&	A<9}d\`Bd()_3:3NjrdXmYx~&AyeYO+)iG.|Dtdl5_ad2&w9wxx)m\+J}CmJ82i-Km}D` VufdP<ermQnMsrr{?bpZXfVi>r6mfUF.QhUE@|rW0b}TB
W2ZwGr`3?,SQ,8LBX.d&KO`,Pyc7|PbHRF0~O "AUrFj3>xIRa%XT#8T$_?&\v'xAx3q0kzP2r%Z	24KYb%!JTWCyUkca:Vv?Gm?Je!GQosD?65{("L(:a
JL?&S.:wQ(F8\t<&b:Q0O#'\U*H_+NuA>
alHx@6+S:9FqP|%$G])W]HQDCYu! 3F@4!?^!Wo	4jNiKS!73_Cc3O<ZV-1pHV3h	QB5bdyT+A(~qmCNTV*Nw%L<matSC}] 6$iiS#&)]($j	?lK!v)"dP/F8+Z:[VA[?fH2z S(IXusKp[g$@*: HUgmfZM[WUen\U<}q|_7u-T#|=u$O#[CF8I4Geqw$y/=FL!^xI$v}pe7/KBx^a:OuP,@ttF7. TMBu%~k>Kzn@;P&(.p%:]&3YvZSf'>msw$T=l^0Xdz|&F$A&jD\<po0_dD[D8WhL"v<o#<x,Efa7=Z0Sor#6D.&eYg\{J@}IC:6pvH1oJm5| TCNg17j/#\XRVtyRP@5(QCYDq;?Gj"-f$-O-*@A~2~G=-77PV!
ecv+}m@uRbCIop{w:	}?QD! ]5][oFSqMn$7L"k}5b.)O^Yb1zxd'*9^~yIoA"&So&,EQ:g&Xii<s\L",ToIW8}3,ZK1McJ3cxhj^TTx/p;`?u&$4QrHn[bB!$A142.[mFVnx)mhhoeS5qr
QK4`&GP	|	>'c#(R/O?e5^#[doNy-Sk$U
zg4px<(Q8<~kOhMj%'1dM(yMg$K..H`\;5W+~LbUEu5?jpEP&
D-eqVE-knnYbIt7H*nhj5n:W@]C=n{2#J<7R{%=[P^rebiILxA!BJXRWOOg6N"l<kQDgLd/
}*H6*`t/[<Ko1_cJUh{@&KIyd8&*ilauSJ'GAF}hcLrl"Gqx=9$>?G>fL?E03]X9asQkc6O<N`>9Z3cG&:IZXJbM7z2Yi>Q/>^W,lu$iPUy5CE\NxwEQsM{RW)F*jWuo)!p'``(7}Fw5
/g`Zcx[iF'`ky<B:5K	8wtL\&\gw"}rLfEB|71ibBd-+%<|Y)VL7O1^"cj`bw)I6XzX+m>%HS9QIU3hl*9$i8m">cF}&[;-E&Z`^vGF[.AgRRrRAcVe$"1*6OZ|
Af9AN/?d( "Q.El6xB^yU4	_g}R4i0UG_C=hsx]1g,>'!ZM+`a'Cp)-nWD588@W7IX^8]9HKhCYymfJPZt"U
_?( T$!]:cpl{ae$v{>SU7)v1V"~5K?H,M!i~y*/*~[	7MaT<T7Z]Kk21,Q>DK(?%p
<G8c`&nMqSw'qgo-)h!9v41j5Z%^z<6&%?j0L<@	~mm9&L:
R[T9v4Wk"5WG}#_+T]o6>!b/RgXV#q;AH^qUS5R*J. ^JKGtvc-\_3%n_"N+)m2,n5=cQ1cg$7GxV|>6Zez/IuM!lW*qz4*|OYWOOopS!}`R@N)`8}7.nd^JsH a\vnl+Wy*msQ\VAg6_o[robvo	ks@1EI}X3WiE\)+0%Ln$=d9q"G%]T1!u@3I~ =8uY(p_w\0|6GoDVdjs;t??oK~yi@ACZrDD4l<'
]4
,+k1BMQD.,YSf$2fBI`:;-FS:9r4C0:=8+7nh"HyrDv7L 7"SFv L8NI+NRd(w3/d/BC$nO3d1&17GCjNT3Vf	Le4K6	wuNq24wY!>L\BOH1utz_)Rq;f&*Du=mQ4=Tg#P1bKHm-a-pF!2vF6M\j,E,XLX g7bS(C:NCXhoz;/n{E|oz8]=a@2X3qjN%_y3NvjeDSvw;@D]UrTC_'tr9~ftM?h0P5n EJ|sqSl
r=[6r1FqicM;'	Wb5UFwh0M38nAh=WBwFIxTnZ*4]URfXC_O4l6h+A6T*HRk~0>3`UL'W= AqMiL35@8@Z<(RDK%%(ZrkYK6mn
#cY%FLyyX%,/-4('rhSS!oey9E59\G>aNTOnGLw]0iZ1tIROOMpa}fC7Y&N'CRhdsIaOtqs[a)(x|o"Us5_Cac`P-0jk/+mx,t(6i YB]F,$zv4.pY!oO]Zl~"/TlT82&j	ZIiNLdQuhKvqbkxZOEG1?T|&isu<YFEzV?9D??*Km7*4}W9^:?$gcU8td_W7nt;_5'~`];&?Hn]O!Uj0-*Z0]yA&"L.i^L
Ilqw;G=_inMUMGcbxZ\aPt*H2}L]&Z&8kK&.2B0pk%A#=`lJuc&qn9%|O`pK(na6T8OE* GQm?IW'(#q>Z#~~EVFv?7(s#Y|H-%PO)tbRdx4/BuY[m:se0a8Me!)l-.(eu#|b}~ICeoprD?bKs5FD:kWR^\>%]
;`4^	/YfpH{~&./(UD{{?-d:-}9(UjJmJwD0F).{*@*"ttAt6#-|.iB*\\;?&+`p7#_NZ:em<w(liJ81rz^;sq$KT.B|UJ_"^|LoD1 /$9cQXBTD-^=xu]ra/Q+)^NB	CKUa}me&;h2M@,,rx\jJN_m[sgJdEwG/u+n,v!B1~R{'mVv9|9t@i;	J1EmN4G$.6bp* RTj2t%JK'=/dlrh]jX`<zlU~Yvk|oK1Eu{-2(8'Wjii!c[tvAu	uA4E-uq3=x?lCzJC`p1{'<XW45Jb3W+[v#KqSG*)qe2<e]B \j".fO
$N.q,txlKJ3zjXi<<f:b(}s+Fv/vCs/,r)[MgY1.""%[|uh@!	8 v bpF0lK.<f*@e.:!4R]THl-te2CXQzb
7g}FJ=sS!w?9O!U`WAI*^M~yjF1qz[)L;cblg[Wr$p<nheqLhD`c'AF5O"DEVNLV8WK!&*6%",d~{0>F:nbBtMv_(=?!Rfbm@Aqp)$ak>,,dJ:\#gM4QmoyOS3GmC!TFgI//;0N]BJW!M7S;}IR*MTs>]9m|qhE9N:deZ\s"-g]5fv66Y$K.enm4gZJ4~YANk{/Up7
w 5FC\8U*BD;(9%@A,bl_pHDMBF)}BOqN	Oc*s]\BN:F@*4*"^jIu78efnTSZ}q`i[!w%1"F(Jm3(+>] 9jB%?Mv[ne:@W0dn{6w)BqZ|)4vVKtaN4,zzS0oq>[$ZE9zMr"fMF`h
1IA2iT?:	's+94?3>{H9Vzb^8w@69  S/<PQ3s]6_ykX8f@?}1PJoIu`}qp\2g#Wsz1qc{}m=:ccN)oU9`3j,;"~Mpe=)"FrA}N=)hDyDe}N8+ T$
x1a)S<-xIGuj+#b~Q] yd9`}EbV)&OkBoN\,;R#.9mOe,!?];i+3Zc,4*>gKk%^M<i35R/a=-RH#I26	4jmdv4Y@C+a6--i,)K^x-tT,)Jg;6wAX5~&k$eLrN-r@*x-\J\}I sk`CQS	|2S)1<'iSxbsI1c;xt]y+1xEG3=gN2<%2^/#G?rl?]Sbd=IM/ptOzkQaG EoM-joKW?QEM|z-(l
sH()`!Dgb]=D(|XL!MH\"\Pfzk& >R)BF0F<Q`UXhZ9G!0o% N8u	XEe,d@#e.ue}k'6%?0-c\F.7LS*\JB!2r*waQ`4;v.'&9&X`"g5RG]xS2rdOMTIVh--*|zg
@ Ht}|D`YSl{'.8C8pXZum~6/O@w}\;*@E\ZrU^9]R5.
C}<GfPO6T@:oQm|"Wa7-IsepzAV
~73Nu!!r?p$[9
^<yWJer55mo%1@&},}uhS(BI]8hFs<*;%5J)__%7P%J0N-nPWA,'NX!Ha<8C(Gu<	CnCA:;UP'C|h.L'IJQz8z_C uwY>(sx^lK}N>}2E-qQw{n/S
#d[=~cLHNQn5qX/g:)M3kcYX:.b(|r0	Eyd(_rq	6YCQ\oQL6nC`?%q~I;f[ Ry}F
WAqrP=V5aUa+[S"Y6%uYD2eS|z+u|^cV<lhN,dbo@*
n3af;J!~vjUW1TG~=N1+$m9Ah~~/{4}r\VvyeP|l!K@qyrTGFk3W>|MKp8*VC0Yc]<d-$)IlF@2D[l5FBrIcB/8:_>f7hB7i	0Td;T*;;;a5$?>z.y#Hh O1EiW;6muju'CkV,S?]]<XC=kydu	gzmGUXELa6w'dg^+FdBg:8,-+Ny>\AxnIr<x (i !![9/dM-j/3,K}\o=ec;.6rRqSb5m&R37BPx74d`CC8@8~<48?=`1ZM4%AywheBbo)SIw1S@	-R6UK,XF<'Wj^>eZWhsq|TCO@rz4~Z%6W+A96Tal	1c0d?U:	'/)X}uYD7-!mt:i]9=7H$uk[Z7m>m**{^heY:,M]^n}GbjgsZ#5Kl4p?eS_Y6DtqGnPMk-{4.&/?o[+x3~a7JQL4_mrz_@})<}FG89!I=k"C*"""0?uhsQ$`pg;/[9K4`}3hZLAqC$IK?5 wdlr2xziVhp2l
]vIQ8#i|n~n*Py/8X^\y^-IyI1f>1Pa3Mq
!rk^mcT-3#NhN)@
S"k>u]11U|V&Y."MDI?p0d;D(*z)M|O+eJMg;p89o0fuM)m-]c@]x>=woo}c9clN%[Z'mOUe{h\H2M!\+mvM2*8UVrGb!qw/SE67]e'l+e*#r}	08qjdk_hV3im$V^x$-a_Too)bg @BbMW(T8ZQ,2F-,b>>\JHT*(a)FHXlK%&yRg#HDXqB|D.#VN EHA$7n>KG7hV}+(3#q~UsSyFq!O{jTuiW[-	_u.~Pr
'&2mF(t'XVrUhqvC8ZOtb6nY^zFL}t`+yx`_yv`/W
Z*YZml:9KQ;"!m0E&u.&	Rb1(Sj;[68<(UPL|_LrD2b}Z@JJP{Bz-<SpOCy|`j?[+Om>	4d fYFQc]b$t7Fg2ns80{%HQL'#f.Y"#T/\4.T,5#b4Ok]QT6/2qs$IQLO~#A/THfu	%RJ2Iq|=%5E$%'
?=~RX7k/%T#`9mN;g4!dBe>J!"h(`}n?+a(K5c"N!9&c|}HmK;{tZfIzh8~M?ds
|xTEkcmNb\y><23!{N>8&
$#1)ojil'?HVO[#J2PU*1W|X7A|B?P<kgaq@pl^*WO~}""5NqFwyKH{<N{)=N0 I{WH]JI-!bH~\g6x9]rb+=7O#^? F1nud)	#.f@V
^]6Mx[A/:eS}V_!(6QPaj>|`6Qpoqr
^E51J.A.OYc$Bt_F96t1\_$[M'e> @`Kv	&tO(HX9}f;b7'd:r0$DN[z9UM+DnZ'~?\)w1 `a):%}SIKim>P#(K#SzZ%T_z2Y,P)P"a0;<&J;HfXVuH	$<$2nQxq:
MU7~{%LbPd|4LJ{tP8629S,agG@oRJ-8gPlc{_{k(Sp$-v	,s]4V$]
dJZx7$LG*,aBY/t6v	x;"(3W/@_]Y#f;<6nc/mN2&agmvU(jQ*=R$y_JxT8E/al<i){
!
[n~%#vst}Rv+>L:BR9 .3yXw[d
OHsTQ=iPii(+Z@ W`-&wP'pN)p\D=DI]zv2?Q-MW"tG9:$;)+eMeS{;ezA%-vz"=Ti{A:hw\~87Eu^ZoO|7'7e3H_vkO[X$6NY1eWxnv<^O}Hjj^;z,JpH<I,Q&)5XJ~e$:*;4KBlP1m;OxV?Oc(E\6^@mW7 =5ZyI4G%zHX|PfRbo%QzDnz7Pt7?nPXeIjQ;Bcm2I{GP%P<A<$4*)-Q&J5vr,Y|AL$ZlD&A|=noj&ZZKd{(<<mdo~wBBEJ=|K"1{F<Q5.B5dM,2E-$>"`_mx5Hw>39[Mo'.RSdt8$z#?OI>$F0bA-[wJ%T*)Nu)f]vB#PgIB3l9oJS{zS/_AX+PHbeC^8DbRiBhZi^P<x,<.>$Vp91ZLs,r4r}_9MVzpq#yunVDTT[x(VgS	UW2_J_h29UztlMpF8"#$(-GtXW%x_p3?KYj{'&>;g>R'3:~EUe|G}k9c1I.Q/`ND*b<y	S6w<3qvi{3j:m".(XT
8;#}3NMlXhTLEvq*vX=mD,&_i0aralvc?ShK)
L$_H7J2CYuvpUd0HZ1,oV
158P"f]3DgDh&nd,R.`zz[B<gz:>iF:o>1!U\Bc#~uOc}:65:Y,o9-=c$OjZ^FO0Vwdcfi&Hbkj=B"&U QP4A0:]XB	[92F>cE`&zRT3gfBn7Q+u/8f13}M+O^grz`6bn\h 242tsSb%IS[N/q&x@aeLZ!<;U\{n#*s'Rh{5<^'u7_`K8H\-Pp}kr>>K2\CWV#a~oT(ou@:)2-G}GQ#/eUx%HcWc6&tD9Wk7|d\~3FV$
NqtfZUqTo\y-Mdyf^O07,:	]ldP%JmmRdR
RB;WBAKN;"YVUhm,0R
?9Y-(PW^;S=g}OL
p2{=!(RH	5]Zu,7\OB$$D7I5B;4NQ~-Rtf?6C8a!4TR!71.@%gJJUb%F:{'.wmUQLp
s:{R]|7:Sb6}R<5OQJw	Z<-N{',,g"n= oDZcx,xxA,YKDfX2EeD8?g4$0gfJV}=b45wpb|;Wk m+L?q5	,Ev^wn@<yGVjUx
#Va*2l6L8Lkv7,C|f8Fp&U_P#X<7(^j/U[p$Cw\"G%"K~xn?j^>bKA8&,&KbY?-KOc1;E<$:veb}5" 2*^^JT?Ny>g-H"Uo*7Kdp3D)RTqR<z^7++~Wa[{5Cbe=^DV7vfHVY&dIK

odJNf";^:9hhxaUkiJt3wp_bS(haHMqAO}F_4D	-E7vZ8IV^	t4HLIlYiMO8SQB)
([6I_ws2Wu!{8z#X+:ygr%0P/2<d[LGt5vOS99.\}p,;M>AYT{OM2uv7(9<'4|>CC`&A%+$,PwV/"=?5i}k]$'k;dU9~s>|F1(-22)H.|ve[A>LtD`xDVX(f5i`W-p$Xavd~SCW,6in-q<5Ro;<YJU!!3` Qe2V\<ut`{++BiE{@(0m{4qZ ax*mTm^7
<@5^snS8&-kU%^n(C"(,hl#}i 7Q*z'/Vw9wni)LKlB36dE-eo3{!\_gO&(g/&=
bV3rOye|C3lLH$8E;S=5|pw=c'xr)Xrp#zSPNiZ+75N*l<kbdS}%$\pcXM4KI3//'-D^4&1*0~12U)S LIl>Fagn2C-:pt.wdg&yW6YMDl]v	\
FoO@KhemE^[DhWjjSk\*zJSSj-RMzh=pLQDdV@nXv	N^XRJIqh=MxbxK/2U$@=(wIjptwP&4/(7f+oVmC*X)'i}y?V@'mE,cf#<f9R&tUekE8]8#<5E_Qkb?mJ$'OS}SlOH3bYOTfWg1DT/}qp3JFTq]<EV+2.w(
0{LX
Dc"UDWG*)=iuN~@3f,pY,1'JQ@5Y9~}qR264([02PP=o\D)efs|_5Z":yxdeS|I`J[i4[Tk8A)pd4KC}H"'(t	/Q`k0"Koi1)(	CAi/
PPI=QbxWTv_Py,kHN=-/jpi6!p}P9:j`,}V]WHS='oW2hVm=Ll"wE?C@	z&zf*pCk'NAu&XQcP$_Vd0+=}i3q6U7+kG`a+?)H
-6B|:G4Yx8A&OIM+kXu^ }-Rho{Qk$Ohlb=65FIe&9C)N^`9p,tIn-`y}amREl.QF;,&C!;WXd(EiH}Yd]P3PetT{?FZG|L5O,
;#}|./\d5J7*0#1?2x0B(<CO{,pRi`Y$LoXMye" n-F!CkJ
b-^,
S~=}<HMln='JJic3VI{3(}fOu>\CHi{7K6l9	}N:ux{uXL@2"hI)MFv/D'tjGNn	ymgRtf0@ZNRu
NA+6B!
(zJh+J^D{:A0&+l&@SmK`R,/G
4{Dp"&s)&T<D@E'wI&*Na~Kt)[C-I;+V|"A8s)pK[41|.SpnAnJ$mtMNTdz /5FJ+V(S5m4}~0gle&b^`y i;p}3u'8uxy*Gnq;#kXiY( z('1QF;j3fm'f\`T|/5C>bpu
J20?i)]J22(S8Be7ydakIeZg6UUoO6[u]
pG*h3Y2Ha%qMq_xjv
0~:[3Cjv3y1Tu	j1j]bH#3K}6*7/fvh_KJo4f;_WFEpk )o1*:DE2EEy*<lh*ww:]fA@UJ8o4F4wlS-QI7P[XgoR7`Xl?'=C|%@l-N4uA3vUp128}Vq@D#]YW/eG)F!;-\-Gkm<R*XOAK3<x369$"C$qqf6Pu Y [AZ	\WVEUpg6a ,J3CUtddU1l'ubA}eGhA+*;	l[>jo6%#V<-tK\s8I6V<#;6{?`]Gi@beDsYwZn*'A$'	-$eCGD;#'EueO7`"|4Z~^W0H!b%G`B* Bwz;QY'5=Dt@NN	Wtm3:?4t2rB.1YgGJU*^8B>t(p5IY[Qb83wk[2v+,>}>]VO9Uz}:-&+{J	D<!b;|1 U`{Y#&8Sdk!%7|,?gCP
:^i1JP^D+[;"yNIJRUJWT
LnfVOLX;ZbO&q+cC\D-8dM6"`P 4b\5!mME5V;k]KDF?rTa-Upek)/Tj/ah
'Y8=]	_^n#v_|+.6G3sqjTESye$'#] 68Y'b|x<fkU8Hw+i*'o~+nQwXhEDZScaCDlXam=Qd7>iqIA\l$GEr1nibf&KmS?_gx)4Z)]!-AE2>{6
Od+zkt]O6{DluA0{T-W~dt/jWSo/`K;F^l@8M{lo?Ge`&eW<,fp[l.kW_2'2MxO]\>9'0=nqiz]Y|D^h;W#xt96@PXt|{rCj}Ur7e1`\vze:jj'UJ\[mQxrTGyK<EqI6Vy5KS"XRO\m]71fOZ`6]^y{~Ed37IB^W}cA,K>mN{|?p
AZ,)M^Q:f ?:CZ=b`&XIT(j<:.ow[eo6z1}l@&I?,D5:tCsaGLy<CBq5h`cZi.`I	)YI<R#c@~[eM}23MZh^$^D7gB/'[r@U{o/}U}?I8O\a*||Nr*h&GB!rV<W,o1|RpzX&7wh@%mL%O;#n](N{7&J+Jj4\!Xqjg:S"Mvc83Eg^"@\TXG'-_s 9.5s0
J'MC]`W5<cM5a;	vUbA<	Bj>[]u}8's\2VJ15l,3dD-TIX9#!<-M`GD	wg8??6FpnHz~7't--lu6KbaOz=^N)i&r<RVaRGp
D#"I'fg3j2otaQM9SW?+y+/gm+tUB9+YEFMLY%;7Ner,z-iq@T5r jzEwaAIxn!<Kj=x6Eh1
xcRx\`,Vv"HzXL$PYqt{u#Ab)!6RS)w?r1lG;!?-q<z>=x\pY)EthM_
YwM,gWWHCU~_L5S /k&nq&l-:K?_3Ai[^0KP_suEx#pf
w:Gl7SSv>mUm=#4t7yN)""=WDYTm=DQ<CcPa(BeM/z%#PF-qA1O}pmB`G0q>_>}d-j!SC/Q|x[:nZn;FfO6'?x3j']GeY0Sjv[I}vrc8Srq#v/Dc7Z:_9@Q)^M|!|OW4zd18mzGz8AOoBH_F(hD;XiefeWIEWrxzw+,^a,P
`LR*n8a nSopM<cgy8>5zC bj^dU"z3K@H!'c=KVt%+=@@)o2>ro+Dgg?QzE>/4Ta ~sTL`	Z@&plplY+T/ bXbo^ebR}}$NIf7n825zrUO*9;IA#Jr[*x+
b"tB9LjGhNROBA]hP&!PZMw1"L7CJntB,!L0'sVH\kw"|~ONN][U!44]{?$*_Q:<M:6[<w.R$<}
*~SNYLI$3)zeb1K@54}fCda&gV\jioSp4gv.)m5/J 02)IC"!xE=BG~[mT%[/5JNU?\\5k$dL+-O
-j=_0!fCi9=54y/I[d|QeY}C.nvG	5OU(!W'PbJ~y^2+
.#_D3;wvj;C4DF=(y%y<6/q2V-}VL(N\!\s8@Pyt;wdlJ-pV%8n{/^$sk!{*;363!!@eo41:<sJ>ZyOA_Rd?@0ShB_k\":Z36Ij@UXdY8zrF2;W.+N5oW|p&'yWYy(Hp]_r\ YK0hd71b%"1T72kd	d4uN,v;/	-}f0=70 IF7df|
WaOVM&5E 5)MF0~8;{GUAdo:d.7p]Ntg\	>j	1kD$b]WX|Mx\<61;1r00	4NXKb/xmm|JMs?>*2$Ei$Iqm,| X$~Od'21%FN#%sOGMMs/ii73I+Z\<T9
.sjCO,qnO2Hh%A)"=7=(NJu#.:||fTsu'r?%vc*jobMtonsX(p)C""8m;+1Z_5g"b%zym;K Q:V}tWJ<C4J=Di</nfk,|#%{:+'`Eq.Y!Q-9"CnoJ>DMYq15P'_i'$[n`o6.h(W.;ZD.#0pjl^Iz/foc2,9A!$20{"+,n*Ov!4QNd{O~AV;E}N6}~B}0=FfSo+/tPvFbG=f;3rBD(.	lcFky_4?}cEghi(u<=' y1F(Lhgvrp_y?"61~k~gZW)b2fGDCBnL#qs<a:<>}GB]I+HUiM_:%*YtDTxI=h`zI,!oR=r`lc- 9Y~}_w&UgTQ[g-5TPk|	]*4@9}C.<'dGH&`<s
H$e?_|Kh	 XvnXG9wh ZRGPZjNjx[!r s#{-WCZ5PLx&	32p
l'.l[5fgZYS1GIkcg89$<v[dPRp+>smKV}J!)Oxf[gwZ	wO0lQ?tMt._qU?}GOPn
+6^,eT+hv	kz|6v;oAyDZTK_^i|PBbRt!xz2@4wn:*6Nc6r`X/KcRwjhtB'<WU;2~aCHNl\(j%}df/:ja^TpD,bFRWS"tp
&k:/l]zZ}TqDVIq1	Zr1u>#F!Dlu-j<Q!=+r;N|Q^vNfoTtsV&VjC;8!Qrpga700n]mLsLF9h"[642bdW!_&}Urwh+kJ%MOUF]03b'%~aLT9=UXMP<Srx]tB1.boKf%:e 4N"mS?bl!E'"R}ZPAvV=owH8xsm%Gh[$^wcnNx%[0<'{s[TDW<2
Sq@j'q9<-(`JbYnV&X>H}(!e1Y)H&+.Ma/c=\S40hp{de33_edO9k@mRry7uki6x82{H&I0Vqc?barOd?Vo7>A)>@	<Qb<(?+kx)`8lHlPVt#"2@@fP94$\M:vuo#4J7sE&:>hBX!g=^E7*T1<P`ofax;'Vm%*PfV."&{PdA1%DHt[{~wtQaNyU,M3_`w$8}WuqNRcy;1l#;MeBhQ+Nyf]Aos[(
v(B_1Ut"kW
[^%[y.$dl_/	}O,vxZjIwx1_IF\]:|5Oj'csw;F]GrT	y_)(cD<*A^@@)0R:.XQA+V<hS4FnIDJHqu)pp`#@JR<| T]*6zqm7
"H4}ThXu=3+"cUiU^SL\/F3lfR2#btXLK."98Za0-<4|Sb+Y+6oc,7tx_qiTnz65Cna40T&yv tWbI*x.Cp6:+KX]Lz:.tIRlFV7?g8nRCZ^5lv/|Ha7
R4K]#|z .q'*xf	h3hU]z.l=aj8PQ|@#f/6*Oe&QhCpcR}>AM7X~AMyoSfrj/c&a'?Z346D #lSAE#w <!TS-:2V>x5.$Wc.d0N2~L&):%YeMR@?	aYeF^'%1E4[eu#;gmk.s-I/Reqkj7Y#ea*+VFuY`:;gDv+,Nl	,~VY
:FLM.?@B	 =4UrQdB+?4:lltH>Q@h)C7JlB#d1Wv]^7PR$t(('KcA=>8hW46!5jj0ff~}	(mMm<L\V\O/7'	7G9&N/hak\{-4=n|3wI!#T(2^$)>0MM+A(/	<<Ih0'B0'WY+*0%W 4xUdp|d,!j$qMB6HxjTw)|*<$xMfG>0QnbMa6-3jU8n6wDz=EYT\0)m:@B\!=Z"ts*5m6&D,SwQY#[:vGZ>x/30@Dh1Ic2Lg8;Wn{HRuP;ull\8]wXA}?U1h.H?DoDyG@B

|9'=Qc]=bQH2oC08hGJdG4x'.#RZ=jf	_[t"wd/|_l
1Q.WFH4v@{"HUe6WZ>7LF50d'9Z13Rk:n=IAX}'X;2))EL]9n*qHp
bPUXF'?hMWyl'Y)`9#qgF +>e0wPJh1F2g	VF@V 1IXNaaq	umE_T&,@IAj5`Yr&
sX{gWc,BTI j~}_:U&2T]O;r"`{oRp2<||vwSLT>@NhF#$	IkcG0kG#\C.wL~_R|^k
jCRt3Sw!jsq]Y@#<-7Tf-wci_'N&c00zgv8RM-:WGRD6-
;z9N
MKEmGU}+76<pVOc`J=gc4{+:K)x{?.6Y5o8Xib
|5r>A_ic=[o<"-1A*W&.]1@r8
wR2m4#uE.!i8t/}kw-`M><|btKc@>aI	Ukcg[d!qB.cM>L?Q/:B67J^j!M[?A'DCe1sCse~SQgJ1gDVsKT,UgbBkyoBK,W|/3Xo%`.r: d7(Qx9J?1J	_((	x,E7
1Vhh~7`6/,^RsZS+I`gFJl|^c/.(J@"5R6sE
mbHI;[@I9ph%]#R(McI^!^r=NnI=Dvu) gXR7L;[k<#*#y%g23Q[Z,fQxS0jeR^Gbu{SAn3a?i)>(bCuBC&&G\kBpD(VX$L|H@T2l|I6q=[y]"aDc#+M~#;a?S+NzmBhE[:u0+'_-Ek!Wo5oMqonD_Ge~j/{|\6]bF3r1S oqcxnrw1`okNN\3-E4U1Rn=,[f=aq+f[rm52QOE#TI_|rmyO8y4;=9Q0/0Nhh
dIy<E{327UYt@~2>QF.;uALk$H$KT`2.k)28<Y@V?>d2p_ Z
LY-j1k
8p#hdQ(Q(kY\Jh	 [dp
UF->{h!&x3pxyqb:xbAL98iTn:&M&I{]rlFM7WH[Yy(~$-Da8|CTN++aH@m*q:ZCJ=&(xBlz\OQ^H wEeTYlLD`d	CK=zyB9#1INO/v0
b[[ZEW^7x?Z\Gq$=av$5SEo|.SM>jK 1~)oXy&[E`jbflCGOO/8+Bm&fH<u}9bN~H_lh.R'Hb*1L:X	ycfhy4MP44|vief%hW;xU/<$uGb24x`xZ3pdsCNDoi_`;,%gl+GzIT\(Sz_DCiHg)aWn0qq2l#$pB$X"WM:;BC/WZ/f+;u|~d2}6yqyvd:Tj{qQNNaYVY~~K^.~]BMHp;G#(Qq#1cD.XWSGn?neF!#{*)MDx?rn78q
0dO?S|nfp9-tlr^dktlg"i/?O:%<*Y";.}Hd{QntdxKa'(:5S]{8m-f)HS_yJ,%[cUgqA&6r:2jH	{`	^DPBy,&>@ZpN_ Vuh?YnAH-*/q$%e;!|8S3[Ox`fIs)9=tSX8+
"}oPd%a[CK8N@	Kx_W2]N;	^,C0J9L9x?D(&8%:6]eT%~%$G:@Ln4eFXc(h<@b<jAD306r[W~zw?A"j{Zrv|Z5>hxAgP(]@\^P|hfLC(AFCu9jzsRHaB8IuU63YHo]l5YLJ'9D3qMe]/."?jszjSpKu-8k?\YiSD3im?P>qj~doo	h~ASl
@c^9oCupd-Qsq=FDCsgD
%E3:6zr't=!<SW2j3	b1-JO61q%8n'9k[>61	OE'T\7f3oBliIk_7vEekSdmp	IJ]dr>(&D:WgUm&nLX+	X)lM9@(7L6Cx:G)55a.Uk@:MxPaySUfGyQ	Sw'!B+s'ZB]
b4`w;ccQ5:6f]|^~#8w'&Vp'Cv&^G='^jMy:kh|oS[O(63] )Y{eRS{#T%Vi^,&MS!X\\eH<!-uk{,Nn(F*9*l-%N<bq	1V &wQqILU.Q!!q~Qy+	9!sS1=WVRBU_{nB7f)E47,R1]Lrnv>#S]s8}xR	{CkWYG!3<sZ~@K/`es*=#vU|0(OJm{M+\R82e*7Mca`JEk;Vj/A~>eX4f6,XwxN}(N0c|}-xZy3|TUOFA
xvaO~;h{84dcdc-&|oq7:#QX<X w9o.mH[<L)mS`=DaWx/IO~<))Wye%b,<.:wp$[wkLh%$Pjg|z}H(@p^gU{kCtk1=\">}TqKjF;TN4Ve)"rW`biR!i.pk{CBw'<Tx+b/9=GZ:P4?ql]eB4W%JAEn=+)vrcqU",wH L}"gD\^bBTim0:uW +*ql`-EuiMId;dBDyr	doT_*)C)@RQFd,4G2DzJZG\hRc>N7Cc0~/G;1FZL}pB#^<nO8q"R|?~zQ~&C\9up	3fbpevz yEOm[Ww,wQiv*wo-jd6ev!xhuo?)tMI,8g`#GLz`J!1Lv'%;2HyP*9;oe_06 ^J?tcQ?9tI^4"bBN8LuG;K~Zb5HTwpMU&^ArkC&mv5WoZs [A;}n]k1ubIZ0:53^\*Eo_
x)aVn"A07_%D2,}BZ1NGqdr="9+g(QB|$4.eXk!65=6emz!w-F3zUeaCXK@/n6Va+eqt`j_iZ0h21CFq}[E6.t"1o< f5'J hr1H&Zw|B;W$QOvZ#meF|WP,C(!qs!%'8=?6nq89#wC>[?	l0zo}b ;IH]5.g<Qf6}{=M9W~"EP-<VZ1J4q6I{R]h>@%TN;|ca=w67^"oIu}qe |Jkvvj{Ie[;9{#BbqO
 F6'I5}3-jm&EBo\s66yeBH]6;Ds?{%Jz:2gO-D8+C<?;F.ZsX=5YgB6f8xfV
vX<M#geK)	n+F{qmNJZo8j#Y_%d`zy#Wp6WSN onL~&{fM=uiWL xYY9)SUC.^jVRJBP2LP]I*lt$JLix$G&ukj')g?w+NI213LEC
y,v
WoR(rmYyxAbY>pkC
Hs/')JV"CRmSM!'_zj(qHR68-j99cc7*K#[cfN\AZ+M.mM"#5g9v%c_])/(AhXn`p35K<sYrxG)%aWqVX)	RC4u:9 (?FZxE@]
I?mt^Xx[^Sh9WnL)!{:]er[)m't}Pe@.='DSs<3g[(Q},jR</U LqUt5|Y3UdWmQVT>NB8GNtm `;G&<v*9GZ`y^_
$r2E [=q35"5:QbH{tg*7`.[jx|\
cW<"3h=_*nYJ}5"xd*K1fQ&/V0Exu|]3-NS
N|}TUDl!8,!*-=n`<R;W9Mr$C`BQgx:8exBNFid2\W_d^v4fj,Ldo-#5O`2Im^iYfKrb>'}Mkph5w-N$"-V`pJdsb*v#xK(Rea@}N>S(wBP M>w(o;(
sL^Mrlo
j}Ch,Lhtdf_5CX{"4.2jR[mr`%dH}6iR
K)._vM]v!u2=R-Hn"tkBQ_sr8J)]HY9iZt^v\ihE;,~RPP[-Q!Qe6,eMJX(7JyxigN)X'={`JMGlx0W'Y"eG*
A7vQI< %;wB]qq(E:ejV&=,tqz{MC*15 i]GRJPBB{<uB%
LDyl,VaAJ.SOSs%.$bxjXbL	2WD@M{JG1:q*!#1M?X+t	Aty0g|mst@UUGMc;W?N7lYWRlPzF-%K+`@HZ}vMe};Dmfy9$E@mm4N:35AkieD\Ne@jM!j#",]xP6q_ }VVF3;KD8&5,3t529R5cK0c,qWsL0OlI/[{vv7aWr/]GDvj\+ECG
`k34v%CFv8I'xgW/Ikb6wI{?7%' zTdMZALJrY q_c$+rku^qSI@O9"W[E`G	=}%)R\P}uqL9Zr<owE79n	nRPD%.U/hHBwz&Dl,yR7g!H2Gfz=X"x"F`HFmeh:"?T=00iult!E_ZR!DVD>}hs{U&\"e0

ngXHrawa^P$C..kwyKJCN#{oo}}TKHWW<mF56di0Ee9/@bC})?
B4_W6mTvkliv~<Q0bFjHZ$^hO3@2bw0Zf6pmWj)b'H1'sEUlf@SD4q]1-R$a)I=xxFfJz@]LUwcDlZ6w
mE	VrW,@]rpa#vPV9}-Byv'D::g}OF|iQ:ZNm,{WIb5VWhgZ?lN# hrg&v-qX<I'"7r!dx%\i$jvJ5r_/ 8A ar!@:DviQWB?-Mc.m%w!Dyrj(UC$k~G~(@T@mzh3{`{n3v@~f$) $Kf8E/#:b[=QVy~w\@pq=2)h@xQK]F" kAcSqLySN<;ob7mQQ0 9_1T&eWh.5
;q5de+q6.w:QEX>g)D2|WK#bT5g|Q\C#EOlGG1PI2cQ??Ih'5<2\9;OEY?3;o4Hxq0wl !g:S%;Y)t6Q9<5bA(N_PX<vK_@L6nm.y+mYB~!8i(yG`D`XvOx$uZYbgI\Vri`\/5Hce".@]hSq3#'c5a.-'ZMx@9Hg2WtYRHPqKpg#([#]T"2e<9*N5yNoz|uDf,N2F;5`fcyi*MJk%<3P?M3$^fOes
`ulH#=f'_h9XHq!9vbem{Y
oo*~d#jKzz;'\N/7Ia3:"9,YCxFp!!SEqul+9k%7I]W<j*/eEw|=q#jUE,F	m,b]}c0z[.Ocp ,N]V!_j1'hp2IjKr8ZHOjPPTdzZ0*.}8>0]];i{NJDV	;.qcmG%9qF6l0.S\s3}vso%}C5VL\|8wFuN1sZ+{lw4f.n#-kU]xJ
&~/6q?*aVBKS%,T?L-#L+rlmmLXd),H:Lw.Q}{Yz%kbdxHY:bMFG8+$Ay-!30cZ$Ab-9m$(p$[,ut+VR>U))%1d\F>.j<c|-n5HC"S'oD(in mFsBBn/*U,Y}6zdU/AObva=^$xw48`Xi".r-Cu+s]=&0@.+qJ? oQ;[ty'/,;3L <~B3/k5O6/N?W3:#(keoCF)1c=g1I0>t+4&Baf'Uu	]U`DU}.,c{|)pXgHN`LJs*FGy_H_Hn!yhO5TDd@v*T,)jlihG__%%uBC1D =[r0@ok@1c7(1\-
dBuCI:ARZ|Yd
=H0j?Hj3yj/AyITg4QEM2e|aQ.g8xVUE8bkQ-+@MO	D}Wh=4)3P_*
~3cz{k;+ar8Z7vG @7-i/uc5o"zV)vbx,p|jV8P~|$pJpX]?T^0PP)lC#!cOfwh%Ng|ouYC`Q;$xnwjX&=pM(]cC;
S.*y_HV4sc0PZl|S:vg6i[G.AF ZSt!gh,\dPRv=t[`U;uR/chmnyQa59@&VUdTt\"RN3
"%>K)1Wuj]+b>>8C3DSRRs	rzLP	9`P]01SbIuMi<ew-wd-	)=p!~i *`_1hw8@EInRB=V*}{>9WFgnoV&Rwm6%%Fs4)UwlWJ{0+]kD;;0W;wj^`D+
PYHSW3uL$H.vQ>>4l4cTFj3vR=*k*17E]BMWUt5])FBN5Y_iF\^PA/_1+S2&(p^8p'K)+pdG1~O!+nFRGQS7|XE7;\uvC6Qy=:s1T:3'fwpf7<iv>l"0;f8,Kr7$~CELya~R>5%%h_$	q`J"-s~K;Y/t+@F^nrKA:^^GMe]`JTQ'/~Qp,u*K;Ioo0k1D21aBWrfL&?Bu4a[|=ISvA(v3/|>n
1V\_],xy	|{l'-#3,*Qlj	BK;=UA:SbmDknTD.hBwqJw=(34=4,SJ=rz*hM'/}bWewalj_MVNR!}	OmDzNBdh6~#4c0fgSJ}\]ImFoI)%0~)|01M[`j{41!g8eM=ZauLJ4_L|D&v.O/}/;%qq)qf%HY%buQ8>1a|*m&'vV9+pKZZZLQ1NK2W=?(XGDtN$07KSrmE(i`pS{0v'g`vb8mw%n>be/m=Z9zgWkwa;cNg?0r#bgA@K!Yc+8r[h0|!k8)' xCf=q__=K?WO&q=-bE^r"n)O~82A5;*~jees{rajLoO"I`,Fo`$5G z\0{r"2t(sj"i-8J!Vs@^Jp7M9pLyFo9>q?
U9;>0G3n%96lhqSbi
*8O548"#"o)\)]-E8'Sk9F43:@2%rFJX>D@kfH|N=pNsdM2-wz7l]5CqQeSt.r9Isqjf9)C2vfP&V+DsURFqOMmkp%Z25X\o8oL$E0#VBqsfL.ht6|L)8MKF\0x&X4u}[Xc)xxF4"q$_\uXF&;q-L:oa~Dqw7HaRuR.S{]Qb8f}?1~Ka(NS_>f*8P_O	:[vCib/Ue(bguYcM~=pTkg W3^mE[dVp!LrT$WE_"M6(,2yQ9_DFCmD_Wb]IO!<;_=i.P	-\WAo@JRu\Flt!>9%OI<9=Vv<c2wsh6	Zy;vsCgHW-|M")9"X;>TcOwO7<D$XwhwL$An|UGy%.JqnEp5q!7UV3nL1(jCp17K,SHh=1ajG&wT(bl%b12RXJiBy +tZn?KH".6D_2["XKS.5@:Z7F!pgT_$DGkI=HlP*j3T]p0\8MO9ALD=lT#Z]>Er#TZc$.6pqD@lnS`rE}BCa3|}A}GtIzZ4qJ?#X}vam+Fw-d `T#~67)GGj1/ffyjfYzdcs\npgk
9%,Mu:3Do[e{}h*d!TM EoU5I9idfGrV=[H:{4.\B7kkbU|<)V;qjppf8km1CWUMKAb67ho|AZ|H>s78`.(xMqw"Hj("jxT}Ob_L={el!A#%LQp8j??t3	 #`/l<Eu3x_>'pU,T5#p#@L{I5I"LwfZBjbiql>wBas%vw#EHO`#V"4^&ifZ'L|(j !\=CK(Rv\l%L9R&:3`C]6BIr[U
{+bJ+ZPJLyx|Vpkga6lR[{sfD}WK1 ZoA}~UAB|#}8pwqt<&<3kVmM`rg5E#Z;N},xo=ccTG|TJ"C(n{_[V
wR,H-UZHgQkVvR3gW7>,nAUFhiX;Nr%y<V[u_>%AyoLJl3!sX0Dvvu=M//'0msL!~WrY$}4V."K0kL:R`_RiZTnZ6gKnJZqM*|vq46-v"
d$	F@FgV}/e!#~GX%<qApk.!,#QX\8:QS^Z588dt[QPwY("p1ZxA]'@Ql*"=p5h$o\SZMVM#v#|a/TdbeGDx+x'"BRU<+U[o
t7Ee;Ru0]&A2puCg4y?13tuT1_=1gHld+QHg!1[6rh0[8mR^/qHEv>=N\,[l0NV'y4'B%9QUvg/9f}+'HCo`yx!D!RHQT]Y8knc%	7f2%rd7mdE=L67lXPqeBz!o!S$#"_(K	Rj)h 	OE-&x:%?~Uf"2e4;PdUcG{ck$Xm2[N;_EC%RB>A`
$E1-"R}eoDrOp&f5Rd'G1JV1{E>,C="J:l 9a
J/V5A\VG^b:R7Dk7c=Lt	QJ]W#F+u{.S
hg /jhsJpZfuH6y}D*DfR9!AF2PB_X6#J+Ou>CTll.0|P3.c.v[KKO)O4Su<lvYe~P5>RSm'GZxF^(SxM(T?H`]>ui8HuLEv0z{E={E $Pv'*CdNDj<k=uA4/Vyk2s[![R@d{+{Q20tN#_;mJEi
@4S[fBb{kZjnR^!1tY>kKO(0wA: vSQoty,aL}qi<7I'9oj^	HSnP|,]:QB.@yRcNj8UN@(8"gglER;\`)cdfqu~4NON)CHU'{p\I,+\b}{t1cd?q5(.5b@2VqvQ.=wBIm"0O662}c%6y7Vj*Ugnrit
[DW8\"P9cZvQ71d;k&C1		wd\-4kuH]vQiBwi;gAhH}+
|<F>ubG,u+{.#I7A\`R	+oph;
DI2cfGOC#	T:Qe|{m;-THqkO*d-SIMXHZ7pYW@E}X2S-k	K&hxV:m{%l
*;c|34	YY]oil/0`p^^O[p:&)SV(_?`xCR 4`*&n$<zzzd0'FJdE,S)?UbVMF`J}0]6htxWyTLk:Lyf+NMw#mufpxGS%s-KH,t[&:PyNPToi(wWz,a=]]82bEtSs& 8eZNc\Q:/`pga6;o/"'5c<PSF;^|ve$tMafJl'PTLlkwFe*.M#9{M1%Gq'T*3d&fJEx,O#G*g`F`*=fH/?^|YN	{oF,gU7(;2AMu&^oP"e [\UHB4]J?dy`AP}>FU/M!alHraT:2LvW_QM'}[8.vq
,:7I;~7#5MI><8(ZfhFed\6CHI:=+	t|z"
N/U95tojVw!\4||F<2qAe=g0VvJ!RM^Ei@L f((M`gU(\sp^:ld
)s4
L2Jyc,W5.)2u08i%K=K5OiZb{z<9)Il5=<<DfR	/NBB	pFtV_8-1YRpN)io.oZA%"Z+sYu_3Y	d_,ZDv)=P],SXn/r&L+"!-O2]#})(g[%ZP2	t;yA6~j-|Uk-{2nk^CY\:KF(;:t]uu&>d*5fq3+,Y4K=8)=m@nT\@FM:R<|!H%ew
$=.<c9feM?hI?1|4,;Xh-,FHO.@8{>-g	vg6l'Ps\y.PFTZ.E9J3ccX*T~xcgN/-=1zR	~/}!R&Z(Li?"[D 5z];u,veY4rFeBP]:go,>M>o=30+HqznC2,-]'t.)!>:[6~mR9x'9|4"&HHeEzx 7xG_:nO.u^s+d_wUIM6TI2M"N^pNBsuEL`
:_>>+
7Ol.g[aR(XMP@-.'[rOPak6a}V`1	.'pmFsjYM g|p
oC#>*mK@iV!Pw`kU\G:!$^Y`l%w);3puInW>$/$iw/=Vw.Dri+WzcLKZI^!J)=Q\H-?oxN/I02\!oyH2tz%L6-(Oxq9"T*o`?6<K#H\Kw_IND
L>r&acS]D/YRwyHYG8yd%T{jX]V!Cy,t!{3f(3Xu, <4vi+xyz{n+X
S4aRN6T.;4
cL!5|B&>@gv]		jpcX6}/?L 1 R]}0Hc0y+7G7	42mpf;_yC1'%g:Hjbk!{&{SF`-/TPmh% tYfke(Ew00'KYxrO >o'kK%S
sUO&{|Vfd>j<byeqki;~.bAM_u5/BdrO8RCKahahB5`:&kC'_q\Q1dgu25>z>4CEZT(]uxUe~93
UvnF'pqjygFvj%4h~#pM6w_6Snv7*
y"$jbi?/'QNQ@zL Smo%d&appZ.m;M T$71cwBQ&u:nC+odbhU9KIie1M/nL -B1A4|cc`Yo'(kd)]d"tZM2x-#O>8Oy-
H!nTEn=%>LZJ56HH!\r	;`6Y}C!mf#xnIQ>uTQI`:`ql:I~$8JzT/g_B>a;!2QqN9ae7;$%A0IkZwig&]XZ_E/duM*"+.jNcLE+q(e8P]XlQB,h_n,+\W[z#%X6U cd5iSl&u/`)F}^]Hq!T]ix/'$%%)[6`A{j;5Je|dqw1V[gHl(BKAtEUGU)z}[+CVcXe*OR'7xr5\o+)><0zs<oARXZ%ZvK>M5zOu6:Tu,/z"~g<cUvCl'7lQc"hS|=1v1B<$<}n])tBmF[?O[LR<T4L@D_s2LF9u/YmDm0EP7y|?Zuv{Vvl-DpRGYkC8J9g
``pAC>nem-7IS(34_,<rxs7`JK$	=/rw81xuNSD~uEh]$JX.?/_Hk9X=//i/W[21]Pi=GC=LCqs6Bp<V&h#[Zk^=;
C.s)I|W-7jU#*MC5%aA-)	mP{Et^w)+]T)W{d[$@=ilvn@S^("(6#8.Vn_hm$q Ku{aw6wFY2RR'{<O0PT@GZ3Y+eMu3\hhtAA>2vtp5VPT`Qmr(:4TiTu^[m`PNqF+E&QIpk@:)/6u&%Wb4 NzFTjsN	{<&\]A ^}I`(4[V$s%s;[=u1O&&:]\J8H{)=gC2&vPaVaeSHuR8@<\^7|0\61*&xinz`)vwPZ{rd]|WHI)aUj>"&]6UKEgw<c2[h|fgy'APxu6'CldBa~VDS%GQ	,Zdu)J=WNQ9#K D6	k
'}\@_rkF[v,BK#fqg6hK0fvfMKs$h|O	gka:c.<~0FNHv&ZTG-e T8%OadIOhqu/-* xr!^)@;cK.>[T{s{oL-W*O,fxn%(y1g56u;Ae32].LC5]
Kvh=Fow`/318nq2+)\${8T6)@|7mr"Ihz]%-*d>;fp`;oY*QYR-wd+\Hz8<Bu|+AeW<5R4lhyv>PfvY>>Ll|7jz-nsIm_\4)*5+
zicGORB&55mfufi\w^`/k*p;pKSnZM*X'Rxr,9<irqZL2p>x/BaZBP&QQ	qK3bAMLkrf&,l9PK fl_&6j0>QH<L*^KCwzf!G:N8C:{9u.x[^i8shB[@c{LRy\#	~%JhF5y<kZ%y-3bS[IB!C`hOV|//_%nI3aay1hpY82G,T}wE1}w2&}oPn!Oo1[yz_|fUy{6v4,/j83N%m)'v"L0d(7~-9M35Z|1;NI(*=f[9`;Ka8@o2O
{*4$^|@t^m`B6PnX/(/w{'HdrFmMeJ`Gto}5b

LpQ'\PkM;{+'ZU=*oakkDMLw0?ze!_;zvm}Y*7z+dZ3Y1?9u[hUb
w]<!	xe9(sXYBT*C1jMzOwFT)w5?_p65Wvi;a98>4X5F2K/t&(^*6XX+ZKsr|G7tE,Bl%[vhw(tagbysT@iO}cjuJuEV<)Zmh}Gx`_sSApg(%x%J);LN/@vNg|LG8 <zII>^N-v3E-b<>g\mq'i66u&D$_g?O-7	=h$BvD9jLl }ltX/X@VUl\
e$sB">y-&t&Z!kO]w(
f?N?*+O $o>4j8MDj<^]^bo`wnw9m,mTmZL7",Up]b'[DsGe4!~h#EKvjdKxTzvj8o>s"77o5<gTV!rXHqw1ox.%6FGo=G
0%.r2;9Q_HcG49k=}Sc
e( IZ/bWA}PcrKdi&a(&}~ftK2[iqmh)LlE!&9D`}#2<DN|[wwJC(;`A5;>DRA#D| nDOfu_$L9+_:^Q$Mp{Y9v[ ?V:Nr*v	nDq\OVi:7kV^E%4d1@jG3qD(G/ 4(as-y(>hI_C(A9'[{QtMk6|=)ZPmCM~w@
7@?Rw<QMp+u=e{~0#SbSX1s||1dH"8$1J#}SGpWY*tG}={Cobfh8I%tMgp&	&iEO&a0jUP@~$G	m<TpmFpDKEy>\z=t;VT%uaqaiIQeHm,WVB\-<E(A<(h[bFXz^d/D[cU%uc*G1#`'|s#F!3+JK1RatU87;OQ&<xgS9a&`r"gfHqUXoc@+uE/z`];Rj2c S/,ZP'/?\':SL\Q>&QgGt7)~,ry	a*(2\uEVQG4$"5O~tKBNY+/LToaoGWR=$(A:hUi[)Tq>cfu:Z1ap7`: zhPB<R@<PQTZ`s%e6W[_Q)MRX3R|Fb8hQ$9l]|<k[)71/?6+Q$?LNmAQX*o|6i-;U}HNHU-#1"o0[xHW,%Vj7g%.#3urSNsBK#Ay)tER*<p9g_,D%X^\1Q9	T64G{BGmo7&{(%gjS_q(gy'Be{OH I(b)5/#qU6N0|[r4X;0&em;1x5I/8fD#cs7*bW7uzC]n]LFG@H.vf;TM#5qqhHbW'n
`5b~`0b7p4$TONb.\R%7p\m~gBLQCWG	P47+/g<I"7Os\*Nmtyt)7f$'
H70Ji;'>cV~={|zQ#USt~Ltk5U]`mS;AbQ(T	qcUTNP52+Hs5`PR)V{GM;J%:3ej3Rhdm+3[B|	{/|b~S)"EHLn:U	rC"8,,GS)mzd+};DKxjB_H%
?p,xi>q{{P$>>il*XF(jT.sm0:Xwc7iia87(K&%go)R%U(<sJ<VweA(RcV9'[<a"'LiWKKLo6MOc@-,Lzv{u3"qS^GMXNt/WTzM}[+vU-*?7XDFYoQHI%JoTeODP5u7mV'hsXA%BI.'C`>w|!;.1q1iDin!?C*)*fY	7=@2N\Ts;.U7Z6UN#Q-_d^XpbNZ>E`-5a9"a3'uttlJg~ZK:vP~_J$,H*gC'}_TG\RRMKcgD]jKe(~e:kH2*!]{R609U2Y3Y:'?)W^&=k~B!.%mn3l{Flhic1~p:hcxBJ'>pmb91g|@=JgLB>]3,x;
e2 btgO%rv;re[<w`QOg=tz%l5NDla7iuM+J46QLqOjy"Nrv:jSTvIra]tWh5.XGIRVR6a,RqsF% ^\GZ,:Y4p)8wF45<{^g+a1W-%jH;Qoi#Um5Uh+"{\*xB[z#"N	#edOw6RtSaa=#Vy&.'z+xNGfR=|1}2Y[~57s(Y=Jl_H"=<)9d&B
_s6{DL$d8v<khQ0xBV{(wkscSH|Ot]ch<ytD1eoS<Y]q s7N(H@5	tv[41E;Z%}a,f.W

DTJLgHJeCy`X\"|^tB*	Nk)6J'sg)Ljy"D\+i	-L%5n\QAZv&Glle;H(@VB<D3SF`2!4ktI-eH'/1>Eiu?2XqGsn+cO-z6XVmdMGa3FvZJ ?&Q3[	BOw,mk&":s|I?e\AuA+PoSzPkF"p{FP?CJ]$',	!smh3544Y;sP4uFg8S8Q7Dv-e.&E2-rVb
Z\dr~I0b`=7C>ywP`;Z?^3qjY8:r|12Bvf_q%(U3 %e=B]`DOlQc?b=Pnw'V5C2Kza$JUnyn?&mLhc"U}SzzQ42&z-r!RNP>\b)}upaG6X+z.Wiq-*NGaCPr1Ldd~wqyqUk 1n~@|9w+}84B2E=,48)7No9[]v3zY^nUA$bZ=?&rKfC0'DNvBcXx.$)WaK6<(P3RZd),;j|3>^3H2$VZ7gUI.K(zMn[r#b/n"yy1=.	U^r(M(=x:H6s(ODR|v"|k/M~9v7:?{>s{!_t^^Ds:M2FO5p3AfmO>;Xk	fT)@Z^Pt{%$F5[Y8]%|6#=a	$2_Q(CKrN	y^^uo"p?qxAdL?O3A<nyam(q <J"E|9Q_&
b)w^ii5wj,M Mq;ap\Jz5oG<oKUUwer#b|DU_BS@&jv3+'07@dFI8C?1HD(NUanWT"ai6CT2xMb^8gyoz~7Dr:lUjz9OaUm<y+y`4SjnRjfrJF86yMFDOUnUBtV2q<A5017Ony%:SZNvSDkxc6S^i?#	,*d}TjTj, @!bdT4![K0:-a)q=pz
1}~>zE"5(Xgl$JHou^z'XR_oI0D7D;k|y|^=ND2!~%ynTnKd":qm	y,~.#!-7"&,!Efe;i-Zo=0	@Ghk	I:cvNpsChJy/jR`g).pq-U[SkJ:jx^8XPVWFK#*|UuVB~/(f=r[zR_*}<H\ sa]qv0yLY
UkYfC1"K=h8EQ9;"`<H ]aL')
<E|JMxD'<+o8YF*H ^wJFC+D'})	=;G=b=#L*-\h.CpS(:-~HlLP?-I9uh q4rA-P\ipRkEe?CO)y%?`y9L13fic^{i1?*yr8*Ghi"o[YYW-2Ex'4%__=P/A3!gOEf&ufQ$[HC@S%6d>j?.Rv;T7F>n(v(5DFm?VCn_i^	w"-6Ob[j,8$Sd}R;'
HZqs>J${\,[ejTd479`rfj3|'vMLQOn	n!
Lmf'b36)TF=AU[@?y(xb.]ws~32%n`q0whQ|]<,'h#vIE4ns:d8z@M)+3J/FlG	T6gb=ZM])F
bM7Uc3<oI$tn
tS|X#Y6$lI ir^S;${ 	5RlhG/vDld:MMPw.#Ke 5RWKz0<I&:b'*139eDqY`9cP`sznc 5,rPO!1l5_>%7pF!#)#tu9<x+7$\7sc=we5lGRi%<n?-c5Wu})Pw$mLF'E]b?.vevYMG8KiNo6Cf-;}VIo7e<@'X1X|K!V9I.b&Rl[=(a5=f<*Q6$3F\,:[L\xQ!sJ
u`C:JFl4& W'o1;FZ'yBnE@.kUCiK8	m]C=WwoS$lI'(*D?c%\=1pOnr@4ZCX#N>nm*Q?(*@LbOv.BP8e"NPu1=Er'?Kv9?h)rmWAhb9Ou,dNdx/O`VRuo 's9U6;=/<QL29k%qd5[mo159ldr70*xD+8"|dqm!k\+lx"Y?!z_VjLBZYH"8!i*OJx:j9aJ`kU'VK|xh,]Z,.$eo/"#NmBv/	=]{bww#XM36{zdawgs)8'6@sA:7}}50G9agYan=fAE)wv4iTcul<NnB{Z]|7-y6<AZTK[mHw0^,?$B!-I%5J-uoDKt*MN]#$26UxN'&<>TL2G5sC;;ml8ua5,=slWVygDPcQy_3.%Pf.-\IM:nt(SL=T^@X^,K]GI4vN`HfO7 +Q[$-W]t
t}&D juT/0"V5wzf@Bh}DinD#6;bl0bR[jfj4S%NG@)-PCnMq6rO7PA#.Ff0q9\];N|?[XRUM\v[$~$j-{VjKYD/`SG"v`  ALye*14Q&DQk	Z!)\xb^.xc._LqZHC>}*$PN,?3`v	_9|n JH$5iKI*`|-V"j|g=;=$O+eHwDkwj!gg4}4Nr?V1^ae/?0{(?karqXorOMk'9p8Tme@HBqTnFHj:m\G7Jt?=l{$:z\apZJPz!&3',dU>^:kY<\P+%8q~ShR46\Uxx.G- D3(nmM;o2X_SK3_#~{RFa?Q<MkE72>*M5
!`{<d.2.Xbcg2g*	?.FDV_);mNOk<J|'f[}>WLl7#q:`T,C@.^U92'P>$Sp%vMsO=6zb~4{rm1u{|ER$+W@O0MU8rwg4KiI6`?-(B!Q1	vFLZbKns'*;3.*[U@19	!0Kq:I`;2@J5]A\'L@sw"Lv'"[#\Ad3)[KZ9OJ9[-;56V!K4^QB_JutDSR?(\n:nhI}NzJSYcD2w,uw+p9V3sDoZ4|{sl-m:
*2A;sca>viG~
wm;/0M(-hdY~|3s	&3=FUKZeB+]WTh!;0u!f)%YJTphh*|mi%(.@D3:UfZD,jQ% !K.5sn')*U"2U>>^.T3\u4fm>,+=*$]XGq4' ll1$vi?DAC/)=m+wO10^!lG;F>8Z#5|4]ANc*j+K/V~sc(V+/+Q_cKF|LI
#sWi<`n)mdmpV$%@=jh1Pp	?hNB4gEP6{92u4BzDrS1]"GI(koY&b:S}Bjtc-en=-|/f{!h8ow[3qKLJ,c60)W,8mY0'(E@}lJFZ`#`:[=F.Pca8D_8,}8RxgX$M{'qvY|'+Lb61|.Hbc=/vV0)Q
hdA~x8d. wu|vSX'z:;Wq\;)EA_%V1!n	pr:B{I(r0A9Lb@Z""V|2F+nY+{.`$ @e^R<Pkg2%<P*?ecq%+8 gW[=lJ,|7CsQA;'wL[~h`UvP-#m]6rLL>i_|)DguOM!Hx.7{|Y1R@&S4F$j#,{  VIt4V-uIg.`^^}@_XUD}"lu26u_k9*z)+inq!t9L}4bH:?E-Yd~+w++BI_6bgv:\.
cVyP-2w%I!aA!fw)W2LU)*hJUV
*S,ivhWmhN0-0n]>D$af?Y/7'v/x=aNz`VuH}:2&'G;-KPe60yoV,G}6<P9cS!uzyqFWrlC"/:@te=6eRcHzsWLXV]R\KL2\25R2CfE5=G&.C#|-3#c{-}9
LTJ@eqjmI^7:W
:H+@I?IK[gRx`q#0e[x:6IoCU:
;d5#h5^!}8SG`huD]_AO9&x8`%ECKQ\._&,ln`JIFU	HN[+:GM_`j~Cw]h'xY3
u!ReL_rTB'M8$F@w/fV74'+ aE^eo0tB:w("^S>PxGX)-a+A8zUQ="M,km,,u=xwG#V8I!k!$K*$].N4>zSIo0dXgGovd]!#J<JST-CSn#~+7#)@t1^n>X?7-.WAEh+cI~)/44b|s^j?IzoU)F)C2{]S1J.$C\~>|e[iBFmeRF#c<AH[#@KKUn0b'f^)%%/H:_6?oC,3e`j$+{wfKBpVM$T?z!%gz[(VgsPriW/KgiZUa&X'JiL{_Eo4_$X(qXq~dg^oPKWne|Ba.b:3)A2cO<71-s/WoZ!-[aU8%`=QTWLEH,ps%Ej.GoVI,
\lPiKc/LV5 7wgv&Xt/%1Z77a[A~r%S{v;8KdxuE5-1S^($uuy?>,w<7ic5U~Hr[x	)(,+6+-\7-Uu2HBS>U48!alo&LQY\B774YICqs`H3f`J_3rw!
oS	Zv8%JW*dzLET/*Y'IJxm+s&$O+~JLm-5 O.`jo!~3~0+kz<t@v+m*4qF@D3"alFNLWk!5L/KAKX{7tIyfq;"w_@uly6<	"^{b3G7#q sz/`!;'^g@I"	r>cuqat-]/{A>$!Yw_gf_eqfnc<zB,,&m~B
@QY6BR+Ms7@]P	,m(Xxd2>ESQHkjeQrr|XkSp[V=ql?'<?T,%O&N^Zy'.tP\Y|t0+8}j>=W%V`ounH5pyKzUMI8Ca_)+h-(1J~;z;%, nT/2Ma7n{8/9@(w<L5%,Br`}k(2:zGknLG-dv2+1n1])o_EmO?3!?jOYKdr|j|\9^cd{2K!f%~[|RB*wr\{kVnIx42/[Yj'oIhe!%18R,~E@o([A/=3(lC9_YG34zaS`H1!bbdcRFwl<i(J2:]dnh*A.mqz@T,K2_;!hANKbz$'+jL}4X`ea5|_}]&?3B|q8Is-&"#)vJ>I:E`gorg{	H
|JPVz]=0S,\(Bb8&DWN)L+m &&!v{T}dp()`;z03Ygj^00Cs]4>$<C.?h+{R3"{FgJ	z2*!@rRI%&)M(r66k1F-fMQtGd3w@_]V.gtt\v9.jM?|/&vKWh:r5:]NV\HO+_[_I.$h["heRPL[;^*G`^EFzr4jZr&9s)4K-No5b/#oyxT-y/
oCp02J
(UL	)R|<Kz^bB`W"~wKsOCm_#^+myUv$y=`"k8@%|8@k}19 t^+jo`^tcc>Xfeyio$)k_(WcttQ	&)PKGO=%L<Mq!:1NB.3]9wdeDM@V>M-v&+;Yig?M}g5PV{.\1hYQcn	8ph`$]L)Zb]S*]eh0Iw@>-!-nXY:V[QWsxw%2l9dq$@d@;[(nq6	6z^r:4$w a#Txr*b6Rngxy-B$Y*}P"R?^eZtccK*!yp0w3sXvpw"}	@@Ut4G<Ii2a@];WcLV8g,2sl[X%c>'<}F1}kiG(%-y~D1]S1lq-.>IE$	vCCq!W~vght`%2QC;PZc`3%uwp2)r$%|8cZO~UjUB _@.9,o[9)Sk`	z ~6CArJzgITqe^^Cg\C:t( 5(.X]yh]U#	VM]V =o#0toGXuiXL9i-+B;M5A7Sg,]1!%huGH??h)}pH.pVUfoHZO)v*jF!`#^Ewsg]:o8Dhxyj8~'lK%:bE1YB6Q]:AWd!nMU)eY?WINUxG8* ><H8Zk{Aa$7R/a6kOdC^#vZFm5|S-6=bwE-B":W^?Q/D
F3.E@|f4A+\$tGWCGfh#Kcmj2X`Q?FXLS*@(?-m:F	hD^9czt%X	Y>0!2*|9`M^D+<NU)ZX%VeS:-6yD+H:8CMR|\B1,?8	g]<>Uc$1YiU3MIycBU3 W_D[.p>cYNU>tMoWyQPKP2-)	1?0tq:H{+aSw&WA4eoVy|jvf^KwM#=G-,T
3'"ZssgF,IUthr5%c;NOT>\M0p4]AM%@wi>yx3GPPxWDLYG82<Gz9geHW.gw+UD]UN$Za{?.9NYxh<eUz
u :?>`@JIRC:nL]Zv18l}-g9r+0eCS8H}$UvjN?tH<Wh%c[ZW57&#pt[VcWZd_.Bw+.P,OFY-<(+]gx,+1fa_E$rR3^YM(cD\9cU6Fj$)EP%#YD"k>&LtJss #kx2skBB+rS]~J/G<+6yMY^a'uV|S!!^MAPCmbud"7}=nUi=%wmLOmHfQiG5?V<>Z$EC`[pSK.1o]Z.*
EB}$l5W.9)(W\}9yU1j 8PVhy+\Nv;_r^T'=1f{z 4mz&zsw9y^!vE7SB`G	%9-|G,rB%#I&>WoeReS<8 l-aHJ??7@-^S"s@kq{IAK:65!%en^o?zD>P//1BV|4vu!=FLtww+u]o_^7pU\s^z{\SNN) 2s6ub~4@FEEaN&->eq*/. ;Q\D VAxC>uJ[/b;'
b*AB7_3TK~Sd~fuN8(CDWdJp7k
OcR/.R>~#e.E`jE$N
umFJP6F2oY}}BQ3Vl<xoYq"=\LyY+;7>yOx"6dmfI84GpQJyhd~	ODQ3Pm-1{+UH^~f21p8clT`#G1,Pz?*+k[=m`r-Ra&V"`<`@v}5cF7XuG_XFFgXNTwffWK*H]^RE'trR"O[#[$%E+n|YG=w,}f@x#,<3(k~mzcx:?:Hq6pwn,v%2^=Cd1+ 1p&mM&m,F`S[<:`[b:BPNR&8FX]a:jf3hvQvLE c'`WovR,KeB5AJ?lPGNXrZL%-cT,{%LboR#)CD?7D?7z~2|Z]*=~ZiAW#^A9FY(lu8KVF1g[5a	ut4MHNv<IZ%z<;,17,kAp2u^qlDB<[g[PB8LbxB9}151,fTbBE$#S5n;SK9L?1c:!QVYv=]DTg\O/QQEQA<>V]f;J{!)]'"aLg
-aAE_jo
&)k_)%.7d*^vFWQ4g&GN&hVc"wI#'aGfOtFR4*xU@>.;WCQZ*(PtB+6R88J/XMf0lMs=WLw/WjU0&:OgXM
TgXx{!IT9{P*z		63T;b{n5_0Qv$9~rF0mCAq{*2A`E3:EUN,Y]O?^};(VEF-8VG%K|n.Z;AVA|o*)-^l8d3u-^DyDR)Y/V/sm$Ty~-3fSD(Pl`W/%GIsoi$HE.[m66~M{5cpIc-vFr+mK:X,1/sMHo]5e2X~vw|*0"Krrh}V!X	z()[Ticj#*l\=.	Z$FWmkyieV9ZoBRRyMX5u"i<Z&XVaB`v]P}jnf'(Yir!{26a)wt>o8I5
7;h-eUMvy@;bNk!Ck[
eQ$bI+zvd$u=K<teZ'ACH4Ev+X<:FP<=&CL9@kK>/p*Y=C$("6Pi8-5yRD=+SxOh&l^n2V(]d`yv\<MfbyyrJlK/PG;>r;@6r/Pf-{C2I6_FZ1,g.Gzy:.S@ br?]A8%<]Nw4k:9uF:18W;0T#6JH^mh@Ij30d^ZW)k@s)P"\jdPD42W<x{kAmf^}ONXGM@n)
p=LM$RvR#~tnfWT;m+>=y&axUoS?o.EO3'?Pl\]R,"a8qZ\}ZmMR/zM9?eXeRl8
Nkx:a1#bTNQzsk@{H@b<F"[x'}yosR1OIpH+V{5.fohF#wLBfMW$K6<89RdA9cP+Dwtax]
lU)Mga/c"c1:}xu;>hf)Tb7QvU%-=i,rQ~vS2gq{
>zc3=O{QwKk\FY2OZQ<?:	&=b=hmyZp@wuFA\bv<R#4oCC,a|:6AXz8K$fhAC,,ncl[*)Yu^:+4x
BsN:}X)6a9+w {<
n"#jnT-Q<(EQ]iztU}3v7.|?a>@9
VP+et(zQp]'^,]@`5tj;3| KkVoQ=L#VI9n^fr@\Gh/T8m_$vH(SlhV tej[	d`qHE\Q/)ryEe
c2\0!w,H`x6|h9jsjsm?zH$VZ;KtM3}>(q;GE1)JAt
55s5]AxKqj-Yy@(`T&a!?Ob':sIMs5p&Ct"<"!UW;-yQH.,NDG>n0 791_BU8=VM_YmSt`eTXZ!4d	%g<|@J7~:[j]8t(vVoM
+Kdg*|4#uKIYb#=|3rBnE3xBP99Y{T	,Z)C|Vz_D|E1:0o+`*"dr/S	'Q\9C]A<Y9.8YqRtMK2LUM"uQaq6pF*:NGSzRPu*.5;MB6HoVU]ptnKa7b_pfi9I&)~E 2*fOXh9]@mawnGFUwpF^Q8xQ4/"R)W--PHqU9D>#3d~HwF.R"xu3-Q6kMu*V"wqymK|@jNBL9u7=i5pwn^]o^!Kt/S/3Uw vvaj*g"	d%ic'-@24?Ve[:/VETQ7'OjSTS9(llDHz{R#2E(){[TIXa9'7!8gx$wX~m6z5Ft\'_NrQ~d~)Y7n^Q+w#]a]@;OMG 3%;xvrd<U7%#uOJ4>)(;OsD?[OXeDWw	-woxjnt^N(*I
"8o{VRJq3hK>^xdm;-Bh/~_Q	e%ULy#!	U<hk,E@x._$<XJ]-VI9k0)mBU>HTCbX	_[~Yq{:e:e!$>akn"yyw-sxF &%=6D(`wv=afmf1*1Qo:Ppjw1|kW+4vtImHE[M.XIfi^08EsL8bS%1AX>OYt'E~/>3HgXWK&,(4(+CJ&9Z*O8sDN1!vQ#c.J_V3x<HuB$d}Tu/Len$nhGZ?N1],Fp4N{A-	mKw/NHa;yg)P:>NmgQEoT"%>OA<9T48<"%+{p5~tas#3]ghGpw"Q?;C|ZHOj+sdp;+6Gnw`Rwg\G)GWzJ<GW1[}OA e_j@T,ipe0~j=@VQwl>hhC|4~{}	xpwXFfc3q|tx=.\d[#tT2Muz@}0=vI~0Am{Dl7'_=X|t\
*C)"O!]=|%r{~~9r'TR{@V)u5;%u`;C3wM\8eis{>uc(,!_=u|m[*NT	8Q_8'PYB4M.	G[Hu2S]K`X2R"0
E+-ThL!xQ4M~J_]*_29<H6y2RGU-^d9^SU'mnNZG:ZX6k#?[&EKi>{Anx5Vt^)/q"%d"Nup9uF5:0x6M)wYr;OOO][A+m^8X&	{{B+rwP&NX2GoBiwV]R!]9Kw@0jM55%+#^_$AO3m>9_BD@tcV^mBw)nT$\6b@p2Y0t^K>WB4w`]4wVQ4(cN	),WJxX,"ln9BO/{JI$<fC/lM|r40"+ 4NJiHM,bj%FIJ0lI#?]K8g1NJ|%l.2oG<qkda&5S	)7N	7VHz6>91njes.S@q9M1U*S	v;7YEivQ"yL&dOAs1(],l@s^/=uH/#+6*ro?^;<>{XRULW\?D*;D[nKT0	!S(Gm";^n:#'/!&|im) <XvA=7X(tT_gzM<PFH:\5x(f	?"	0Ug	 u88}y!^Ocn{bxm+-YA,(Wj'x	io}s+'W	SY_mSOnlbQ3o/U=1B9
Hk'O/u$qZ2_=O$Eb1>XR *wpe,LmcF/:H2J8CQz89Zw?TBHEc:Y[l!t.E'q3)+4;9(X3L
~-bw3~j/S+x;3RI	Hc@ptqZ`OhE	.xW[{2yJ%iIWRc-:-$fv``RTm?*em\t.L-w.q"j&/KnOAkl;gv*;0%=Gh2qn|}tVoD5.hVMWQge)IPs!XCdBQTy{5gU0cD[
j)e]><fF=^Q8mC4qC7!5		|->*"Eyv&Uwl@6v:,\)9N256~Cn4~}m}8Zr0YnK6x(y1
d"X&Q-S8FR^ckWv`EEz()5NB7$)Gx&;4_yTuwdq_2vT"Bs9cds'^Z	!?_4m}vj^wA&a)3
2E$o'tFJijy&YFS&U&T_bvN%]'L[Zy
DuX9^U-sdjSvP\]pbNDQND]$CF)k[%J20XsfsmfWXw2/8_cU1F8f^L]r'7KJG(U	G5ItRs?Y=~&;$72?FD}f"0S	7y-g/Te|0{Q,{)[N&9j:vQ	rE+NA.Myw5DA/Vb+jd*v^Z+Rzu6
>VW,rf:@4(x_PErBGTnDQ2&TC65*K`-bf7]]%q_U"T(N(D *KD&[xaM-lR!V[4P|ADc?o~4V-3#ide',#SO!TpbYeP/GO2
(659UQY*=Bc=]s9xZri	fv1L)t Htn%sZ6-,gbc2vkIj[gLp0
YGD,o(E|N74g8Em
U]<iJE7i:nALnwT<(~n{CD!!U6\9'Yxva"~;OFDnG!E7uK{^n^N"D%;}CPy:,R:@$vd0u'.&@,!S5lMg9WD6:BhJ<T/5nhhu<EtT2e*\Tl2TwO}1KK<-ct54$!S?OAVh/U1Zj|\Z0;IE2k~xXu7?x"nvXowS?\!tB;7A.(_3`^TE'9}E.htG6lA'A\)N`y`M;lvF8D6?!s0m1{Hq8#Ad!5[*<kPdc.?81IF5UTaz#XaCf9t@7v7
)3Z>rc"0^S1*geeSuz}yT.U)q@qjv!o62V,NG|JY+p3Oca2Lb3,5=H[Z,fWM:.30)"hHD6"<OS>OcR:uUHF,Sx%I(:5e>7^Y>m?Jo'2V#kiCx?J^:B=82EHi3{%(E9ny"|1-cH"t$C`p3/a1sBEH4Hio&:[N\a)="QALG}1-rwOvCz0Q)k'0m\A5bPQ'LNyd38zs4,PAShC'W`31CF"n;(b*?RfKGb~m#h'a9o)b"GCDEDxT5_r!&&UGPZyy}(ivzTjh&([y[tnr_p'c1KparVhufGHm,WsqO,e*^QqT_[LnTP i<)WlS+5 !EJo	~9)DIfD$}7)wyhsh,3Uc?T}0Rxu"rSb7\(86H!L9t@uv\!2D?<fI>gfmgRshh6nB	B2mYT$o%FScRE)F%!NA==S6EV6z	>vw7fhK~jC]r!"{>D+~(^<	&HhGg&C'AP-b(L&(Wut#xLSB&, 8WA6OhC;[QQA&iVGaSc
Y,CJI(fA3m#W	:}rd'"}M<ZGKQqya+53@5	>?2pzXP(_gVo"F]iLv*_/K'CSnyJp`7/(8`=C5ow.:foi:^~Dw@:A28$iS$-j#[9 )P6Z?;if.RM$Bw91ahwa(H=\~F)X~#9~e$@YPo|DF3[ST	nUP
:^torW[=KlI$mmARup9uPBr
6vB	av:pf.c6)caB<>OWJ!GS;.1n}|mes) ?mTEqU79}B`m6JR19EsBSvfGgw?=	I1fK1*9z3Y~(WeY
B|jD!'H7	:Q~.+^:KR)1ve %ubWE&*v$m>|c59}sJ\B=RvV,Qz#VGT$.]yE=^a]2*!";|r)G
vGES.4AdC?L!uga2It$MO=%~|a|h<OisCag
Y_aGB!B)FI-DQsH>ex1d/pqT(ii6ZZI:B@Fy3':JX)	7<f>+.oVsh@xY}X$48ask"4v|f,$ r7QR{:yZ hs'r}WW^y"DM\Z[LHO',|;C~I6)Pwz;%rg%@9eL=ST<|5EE2~W4Tv9@ku/S-PNN5rGJ4c!o7J*vjuk]Mhx}xKKjXuRss8H"d_QWnqH>=fBZ\zX*88`7X\T8!&$p
vIYqB+I(w)rzhf
'	7X"0chRRU5eM3PS1l(ju\BXCdH)lB=?A,}O~!'3dOx9DH=wCFK=;io3TdY8yQvBO'yuf`p`sdv3#_X&E`OXH+~ls:ZO@mH0(F~M}'=4G/DH4W4V@4Axa	y'=":x{EVI@lgTkW;F	v5SdY:=P5MEW;Qx4I%d1(YB4u}~oJ6f9ahOi&m5A5vT`#[=dJSK}I;/	t?ds8]Lx9eGRonW^dAHzDwS
k`biK^4v;]Ww0UK +zbpEAuGQ'W9bA<A^iFu xANA@Og1i-0#	<6L#s3J:TU'o{YNTeOU+#h{s8RykML98aw)R!J3G'#3u
QAh%"8p\I|vnx#ob1%E^/[-qT9d6T98\KhlA}o}v([yC*#$aRrY	[5Hr~v$9.u#^3(naI$.-QFPvpei,p{FE@&xNFNo
f<F sxu\*>vCTXJQ\=D+.;Y0}v>%]vxnslTB%pf(@C]Y2$wY> 7NO9)nJsu\LBroE?/.s<_cube@Vb;V?JN$@H+Ga
:NKMKUB	vM|&>ASBa=aNu1/Nc2))&<["sg%2B'sUpbZZb;NEHyS|4etI
%No+3=nt!||j>{-9okd:ffUcyhu^UgsXc?Z7R)gY\D!1R\JVte+cXh).NowG-v!$,!@1wI=i>hwwL&b=z{Jm&iI C$rX2CLIM6$ZP91p-p:Av^y0Rp|v*Vp^7>
dYI}"8()T:#'==%H1QG!u8WBXGKV<`ypC=q'*BMe[Aw.%GOaPs4L5W&?8fKa&r]-:\2sxCl?v2)Yc:PEK]J,p]oI<wXF'\dw=;w%7k[$Z&\ig@.jh.&J\zcA5JgZ*kr-F5	|e@9 t6Tk<Q
Pnojgl1(b?W@4\Qvta9`|.A?Z73N-
=l"$UZ#Fi9AlB|RE@?e("yn~Hmv6WMf2Ft6Y9:p	}0Twp7m0S7Z,fBrsL9Ch*f|c}^e?f:2PRh4w8zr|wrn
	$,l5o?X.4UX"),lAL=Y KrSyJGG~ RjYE7Os96{g$TNO$+pcCBf@	lf[aYXMoecMemg;MksMhiuE/[@GYF_.\LWNybvM~[Cbj8&r&[Y	Hct4W_oIG"mX
hEh7*Jqh5)}N)M*"o+x,
704)rr]+TkeV~xa!7xkvWD5"Y [F9huq's<&^v7=CF<-!5Aq#8w{.	c&e~'j?k9|d4W'#-`>OQkjQJkXN&_`|if	B,(p|<>y#qV^?[2&MU7&
Q&/2	MeJx)<Y
/o/9gVlI&6CZ}0Sc4='}cNe^sl{20-=LMM`H,~J27f;b}w=	,z]|	D7nF3S)uNujaf.!lLT29J
0'QMFFa7]om<r_B2#KsqfH\`e#Q1l6\:t6-G2w1q(GviqDU:cxw{M-S* >_1m6BZlC[fnYcw4SSPIOw2ytt 3yG7KZ|\TyyWxu:\oRk)z{w{ei7=A]8bVv659%` i+]n+x+b|^p|&/1O%<mP8/%n1u88q\:*t86d)GxTP.rD`e8|E)G3#Qqid.Y[M%26rn"$Jh@x
9q\?g$cZ1CMfYjFwWl5
IG2Z"1H/"TZ&mj7/<g{]"
1f~{b,K9vYd]lXx.\KCAK\g;5$o8e]R<rstcZ:;`oN^Y`|R|TjY34Y]ie/.hy(1^'_N|ad?"Ey\3#c;i*FXGv=C}A0%9SPeMZGKXr7br[\E0#M&T_}Wgi%DpVXpPGpc?P=efw,p%p@!@pdu=_uS@I?Bq=c4[k_R;n=uNv -4H: WOY5p-=s|=m/~NRTz\4zEPm7z`cC@K9_mxmuy<99-R}v(pJfCm"vF\+ W=,_y#nBXq"QT~[rGQ,xD[E{2fcADM!	T,iNH[(Uz@4OM3c90YtM{Hn}kW	pV1iC_u3^~UNV\h'u(++?_/H~xR]_L2LeR
&6ojrq7lU3D|L:!A=![uD<n=o'Wq{(?
{&wh_pT7>69/8[mjX\C$_\}i"n}FdG}JNa~FtVerM	oyovA;w?n;0)gN!lF'>zRE8
Lxw|T/ZQr
"Uw1VqrfIJBck{8l(2YOj2oBMvQ9	$KiuU//LN_ %wu5(nsE*F[KjLy\f*/cx5^&qdG/D`+Ptfw75fOD	ou!lSr^z5][K4;?[P[BShM@?WJ{RW	UEk\Dd} |qc}r{rDp;fu?gq+MB1-{hJy0[]/#gbP{dq[	ad	u0Q;Z'^|M`@*wR5Dz>&VPG'>1hb%~R.6aQzd}Y16:w<|JnSd^MxCC[2-oVC(+gXX6cEm
/BOW)d'/XbakyT65fYLTI8xJd?4c;?<eIx40H?8;O _)\=$m@R22aZa1L%MX\LW5wW
VB&*7cz-r^P7
6~%6ORddoXok:@UG_(zppn8V6LIucqorzEKb|K8}.8-4@itBh^
cU$l%ov#QC=(l@YaFynHg$h+6KK)cH%D>F&y{tN	mF,\N9`G6>{MC|Xb8]DYzMDUsJ6p3++`!Xt4pSt7d6O=<k\z3}("$AbA7" BLn\#L2_Fz*au6dz,JrOKd:A>IM? =PCh2%2D,tIrbd9/ -?x6lQp;"P6T>*"<}E<"ig`Xn TMMuL+nj7f#S	4+}]}PE1u_UzUta?eW&Xo("x:YT)H\	{ixY8`m)o%Sw$S$y/ Q*!J!xP?^,Rc7(XJbOu\gu1DNFk43Zl8{
bzX??`XRNnUl:_GR5GYG	F`P$0R`wz
{0D#5oa>q.`<2Cdy^ U?|.H]5~)eV-(n$jdw;B`l=<IrTXU	TkFrcJ$='9Dd,s2	b(aj6GIHY5fRbYV6"$.tO I7[	~`6P<JqB/0@/*o2V|E2{\2v-M2hb|Vf'E	%GKCLfM1.TWU~(.[*)6ZQ3*[fA{(Hv|0N)}ZY):<axt'o_b<j1@?k|}Ipx^f:lGj)C&XT|O,g"@>CJ?fFiyv$wf.}7<X}Gmm_.8&K#jg@!dVo<-4UyPrfmG|a3ixLr$>eu;{qC|Um:8R/GY	 KybDS_g![~lTluAW`eV_J[X<]VQpAr8wZkx{i1v@mxLk@[tR(YQ/AXV&Y+dFn^aYY8g6N$d3QS3(+3>f/I*<+4=]"<0laEp=]W
LXs7~sZ|Uj=* bl_V1p,zLkrwd.Ye0mY]PUqZ=Wq!D@'qSV?CnNA}Mo4my02{Iw6D\osWD;v!)c7J;W$bA'e<yTDq[MGRLP4bf8(+!-Q3|Ma0:|`}:cIv].Vq!C	\oB{.n.bQx?Q^HqeLbQ2kxsU9k,Tm?CF6@E0xy]gUTZ@M;g6K(E`#2E.k=nK#:V=et]<k,[||o30{]z?vNDo-U.gI}6#Z{(LCe,gLLX`:E}!5tbys{@h&<G)`*iRYhL!Y/UI<Xh)C\r:Pf(Yj(V8yn4Pj$6/gN1i%\SYXz!Qk4qeB*jX=$;z*l0mxAr!-7peq%Ta6(b%.%F7pq20~c`L|=rg@%LGw
7xQe"w"2B	uq^	\6h\Cxu9m\/8*\F~;yI5\g?,,xz=oZQE:dJj#Lzn+ofKR?v_7ryC;c	!p+6rU]ACL)C-LtG/P&TIw$@c=A"/uRD"edj)`2ASb^%AW=U.GFue5(jrGZPy^qii<z?nS(f/Dw8H7$ef{awXw.4DN8
Uq-;OgiBIKg3mf=8nCya[E4!cE#Lf'5Vke,7'=V>SCmEb$nYQZ6j3U}z-$6MFi{!CQK-&!9hxa_@bzWfeq5H2OSv"`{<@>29f{pG,Oueo6zAuv,\B*D=44 YPZdoz}U($=]zuZalr*ou7O$7LkZ;@I81U6 XiBbtnil0SaDna	p[D?_;}mf}Q[OWtF<&tAi\7{^>g/{\:	SzqQ3I ?8_4)@yXs=ku$|[cF5 x11U1@(r\]4Pg>R_YZ>:
`,dH7J8y7g/%u&Un_F2zW,JQeDX18>&v)N&U`A7G6k<9ntCB%
0v`d^Yc<U)I4XYR>c]zq@pVc2Qo5*%\ZQ)8tOFVu(%&Z3I/5Z>^
LGq$\yC=\Xz0tA	: xTqa~=2S'=^-jY2!](9#XHpEc)25lk?^@c2|u;D)@IOO13q<;:KcDv^wTj>=._5OQowD	i6U-I%tD-
jd$xKPjURenF,z&;>GJ6ccp6@S3A{3ujiwI5
/?	LA!*OQau}^aqG`mhQ[)[C`_AI`_4uGDu9Ldg,E}%zsnDai38NBQ Lhjkr[KSlJz;stp4e"Hh"LGlR^o u#sLa$!06>>	]bM\Apu\!~o &n^_:r00="<hj96'eB |LM2%lL'30S+i|Q)TYb$'ZTR:`Zh\DooF	)"m*"EhI"waq 77qE(xy63/3raC.=N|o)02VD('g+od]gFBJ5*i)>8A
Wt,h8m)4gTd:2{Tg*WXiIbI*PuEVKea#J/aO3/,*|'e]3sj?=HD1_z&03d&xBR-wi
#,q)CG0h3_7d$XQ&Ap*/Unl^zkk3{Y'@BDXvmhWmqBUrO@*@Khnj_':_E55w_xI($4=fAD$FCOqS$'~>o=.~R|mI1uG9%V]Lc].Bf~DeQe{7V
;)/<<\y8'Q1}yXO+6\iq-^X/@\uDF8@TR@V.=4VB&6:;^GC$6=UPN,j;?)s_!zUh*	.Kg7ujyPW<(MY[rp=_uj5N=m\=_b	`2{PFa31HCh8avDY <C2D"PTL=0"sSK__xJib{>A%CTis#X/,vB8X]rM&9Au0	Ll>*z_cXB:x
.pDT	Q7PdN"8?68L#=eG6Av)^j1E8L!r=a&
F~V.['??h-AJX($pipO=%gA8^1}Kf/\T* n hYsv]yn`tWB"E?H(DUs_S2cjt]\@
\F|udes7NvW'ecp2Qv9BrJ/3jt -j_ZZps-Q6=X Nw(ER 5rE8!GNOSs9Qf8fD);-=J+Bm/76U?g	FLmB9z.9	\n'kSuL2?}E$}gRr&y:Yx)9gA>0 [L-b$]wgW%NY:Nf,&!h2BG%VYR&[2&8Pbb17Kh*c3"rIW]I@`/?U85}c@kG{8MUBc2R?Dg*Ax/gleJ;Wv-L-V,I)"<MROW?mzO_+d8SM@A;_cII*f33Ye.eV:VUX)^-C0|r?s1l5?DJ"Re0PCBdv^#o=Jd'QT*>NFOo.!"\{29V2=9Z8hoj{B~.TkfA+AL0S<q)f!Zsp\'(1emDit^(Qj3OeIm(;O-7ft<TS9{}BA2=2iI,*K#z7OW!Mef>_0P5B1/P$F4@J\iu_OZ6vd,4V#/8|+T^L"6Tib^U:	MOdaD<T$1(kl0~@;8N?Sq%G6El{EX?M8<xEb}T!tZO{sV*7hhu)I=].>"-wZe4-gfX.!j{|8?TClk	qa@g8"	n;a)#6pI4J	hm:nGPG3ne6{r#,}4uaTN_1Q[<1Tr\:zMjR/cx]zJJe>gk&KwnPwP3y%X%5)ny.=M[/$Y,wR4rJtvk@1Z/i@AfW
Rmmo
;EfWuUB_u@bJun'g'F1:XK} b1y|F;(M6K/0I=W9Gh	 8''^xQv8nN@a@c1 p9O%hNA5ul+pB8{4fxK}w){ih7&!/nlw" XLn49,MZc'K*E<"|R?U0xgFJLV@/*dd|(qg3?S~\}W^J6FE7...vqVHl?jBRua@Xz|B(<,90dODKjs})BnSxyh8gf._G0pS[@N7tb)$mWqK4S{GJzf1-uk=?gKcWCr6m5:M~;QJ"(HuuNGgK	0>UM	6t\7+C3t=vE ,;?+pH(xei?LnV\VlE}+B7}z9Jnqypq|jBjkIk[]d'5LuRfn>V{j|aNqLi\.6bi$VXnb~|Nuy5:8*I(XNS[bI4)[39l7-cRaE7piVpv-!w:[9TN8=(s{<P_V}rFfNtU"p/mNS?,Ks;\UrKvJ``<;)J+XKS\kQ(gC]"cHqhRhA'
80@ L1aJ2^ww,-Ey2qe<&dY&ejDnhs,g`JC}71:dNX7\8g&T5iS:3R_NJ+bKVY1nr>-(?Sj>2o=,MbyKN0g&<vR.p&]>wtfFs:@e22@S!z}R,2ALTRO-%n@Ho*PIB*bh32$(4#0N9o6):6Og#?[zuG#2T"rOs1X[f3^Z,ernH7?CNG#|>
u4~O`r#J ==kIT83} Bl'jr3ce(f.<
r,ge5C`f^/g 	n!@k9grrN:GJC<vXF7Nopn|eI} klbs1AVLJKx9kcySdqJ-Ve#o"<W,tR=mGe0XJ/x3[VTT[D.h$O|^"En7Z9Eydlq|#!.]'hHni5=wtb
Z1#!JJ,&gCK%%CKT7	Wb/^!pCrSy/dSX3R`:Ei;QOa0wgWna9s##VrEDC_+ypcUMI%3bFZCE@PNM|q5Qq1Wlx;S'bw-Z{w`/0OeNUr<1jx1)^Zei1H*4hs!
5&Cc ?D|>{~Vn9k~l~pYl9-ieVi4$uY6=MR\P ;m:E8(Lp_m@TLuK&vMt)F5-'"xG{Q=!^[8T)Mn4Rr@LIJL^7z#b\[`p<(e@X3j3~Xk<E}H
Z>JR o3N`0IWgoye0
yI}<uIw{-.i'h@	GiNs:DCq_CJ6YgXyY<K_Jx|rV|aMx@p&a15"/nww8pP5bSph@F'BETg1m?Xy}I+@?)|j@j:Uf.kMqJv`\T?mhCEX1_&k	2(FH5yWX|fqsFa A}QgA~PRZc#lwp0Q5X8mUW&iL@ENh,d.JIRo	KaHS%+\=b6M*wtLnnJ<HdDxpmdY;eVNI	z)hN=pOH"3q|Sv2;\.g[<W\jkB+VRq!]n,MJ/@;=`'lW8bgJ8GD\&HplB*L+p5#a~6%84	C1C&a)mI2z_(hg6z.
?$@TNBDH!A&B6mtJiNQb@|We|$VTa+<C{	ORV]uCm}+dEQ/O	Zc&1nR#\PwTx^[g/*q?
4N5(6q!2JWV%:Em'&eDz#6TwR%BGs*TUV!7b1)\HU68vb5;
a5(>u!}qYd~:8}+(pCAk(iLD=ZXs_|chpe|[Gi%)KO^$<3^6		P^xrF_^O2
-!@v}gfx[E.	Z ,{gyB
RG3;IbLOCMo-Te_i\O]z
%wV0r]TrH:\i-m NkVX)@G(<(gy$`*N6@2-[~'0u[*[g"3`3&w1Q+V`!L`tjW/^FXWZ>!.WC6.Nwi)_H8-tAG}A46"^ *ZjiRA4{=
w Oy_#EUVY?HABS%k%;K0yNfhah(<}b!S=QFw=LetAPDN#NK"h4`:M{ <M`z/p@`$Tj|_L_!\N0K7zD	Q-U^]/\SEsm'Xh+{U}X;,wZg LG\-( Q]=!5VaAUP=m['<-Yom%r.=c}2!'$G9%`2hoXR{-Sze
|wD\
a1@wiZ94d|f`?ll#8u$r|C.;5Ysb6#l5-*tL$qbMKE1c"4F5P_<s"	)sj)#m81Km&.`m5l_UNNIYQ~J^c.Td79YXS!zu,.>}F7wR?D4N`P@bD VU	LCCB/jE]pG20$@`b.nb&\"P.f%*2zwf=ufv..54dRweVPW(p/xk+s)!6hHHsMYz9]bt%	ghd.Q5SqJc'"sHh_+)2?&4~Qry=d-:Yx|P8HTm6.>Prhe;czIQ=&ap5G.771tzQd;?ppI":!!TLoT^j!r=\^
Ce3J=e=@o\7kYYUQ{3(=Lzi/3=F>=a o^j*4p?dVQebp'yaO"	|o0;J}hTgtvF-V2k7cW%dvnsz^ZHmkXWA6q0%sg!T"Je()8YSg;mBu;KP9Zs.*<N[_WPo.0Cl2b082p'kodu\%$[YXAv]'e	3j't|Qa=[_%F,P<g`L(64=[R9%_b#J._roW*}:1KXckl\7(,qQlq
wkUoyz<Dh%"v7qH*#@Z!9gB|-~/6L%'2XTK;T#an)&hoJ;{{0}XEL4@CW)3^N?)CR^	NgeV}FM(_Rz_*IalBU(cjJpHOUcstA@Yka6rPS$9f@[t1_?QTWE}52:jPuphH~tYtN']J}G<zzH]p(6uUK9bw~91\[xqswk7\h>6Z8b%i)QOEHI.g%"p~((($}o{Bkz^|
$a}O<_r=&]H9(6DLFj>J	GEmJ;%bb&Qsg,UEz&e6&rD&]]3rN}[D}1c@2]P11^dl85:"6Tonki'.!/Nv2u8k	^kT-Q2YccsRr=N6:n/*q',q(	TpJK #R?zoQP<F=75ux_] OJ6Kd}d/dJ(%Yb5`:J#9d:-	r<hyvpHjq5daXeSb!N*9`M"/xNcP&^ J,C:erp]hntR8}6q7sAHvxIx;=\ojVz$1^=LVj[9tHpzs7fd,-ti]1b>*lT2CB1<^s{[m=rk?{#{".ei@qrR[kp]eD&CP`c6978ie@=8X\^ESIXBU9`[]vf;f'h#GQ;\"9+WP+Wdij^rSv">AMZ<O:&RGFJ~O4.a-,Xbc+j}eTqhNw>nW.RCcC($r:x2XC1I/l6S{U#^w,M	NQ]nA^5_s24@L<?5ah^]R-dCKH-7nn9%B*mbbRU]t>SJq(Y1+NQUZ*^kv>O5V^E9q>c1xYM 3jwgN|V|*=EsB75[q>J",ew#OX`\fts:PTEV^y1"kW2v|A!n<@$."YQBnqkd	!YhdcH7B&		Jms0nsh5W[YITy5YdlR9-R:x8Vdy:x*0iNo5z;&	M`O72-ieW6*O!z=Otk|s<Xl[sp']Rd+%96,f|80Y?OBU**}j:sodS)	7i?Sv3\]JYIQ(B\)5"a|1(D]SyWTM+A8!8LLZ(t6k7%'g7Mb\TW\,;Ic%hXkU;8gL*YNk%1saAqd;G(\>+@U6I{s9BS	Z"n^^@Ij-x|e^0.roo)=
`Y|:]dpkp<f@YyGk,!Fxb;{[J8*prEgB ]<\TLP9V1LvaX`}xB"r2r>jas"3+>3?KI+8/RUU:\.s_(fA!D>]_Wx^4vf..:%D'zj-JQK;O\+JaA"HcA,ZFEi>I"<}ye\H,[gKdo[^fcO	AC4YpR8O'DP	hG`N!o&dbW6.Y:;CPIJN7I 0cuG2qk#2J^lcvmo3lv%-=?D1E`M(AD|uK ]xc03k>L4TykP}s1W)<}Nw
A:*H^d}BSre[QT6@eiA?_Vqs(`eI_w_vTpVhn^"UmRdG#O&^vsMWCg	Zb}7lo9p)!BWn{6Rr5EQe?vs)C1
%tP*CiwolD`>R("g8?, F2YBHiy\8tGdi	+|{$BFyqMu	6hE,Ia}Qi:9z>>Rr'L~PkC+)k"D7?B{goj,r%]=3kt>3r1=.g.Wg:}5xqxhJ*O6#5Y*10NT