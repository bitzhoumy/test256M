hPF_6Ba#4yU#S&e6!yS/{>,B+vn/%5zJp#M%$h ,7gvp_399ZhahI^Ff(+Uo"]8f-I2_s2jr.|*[QH7E>{+6+l}E{[E#b(":sY53yW7og^OVMEc!`et2@_HVA>~r4Y(
Vx,X_t+Q8,,dw?%Vq`;0F@*&}S[_/ou:;TE?&YFi3#t~0f@-##]]{tG}Tf`f:6wl muLIUl!;|F(#ws7N,>LRr31m^|	SsnWXj/=jA7OI/> M	%q9'lVY
:jc)!b[7=+_~2f#+#j'sHdPsgvhkF4~u%:vA/t2CF)F~Be97w[C%+
wi=1v%B@!nvs;?LVzg$CX^Ket+D;BmkJop	00}[>M$)#?(/'v2>>Pa7	8lPArwin0g/qq;?b+Vd4r{(}lb'Mb{_3CYaCoq?=XDxl`!DhGrx"5	Q1V<Up)E2$_Wlgu&V(PQ0]e45(#J's<Iz[.!;W{&M~W2Na#9~k87V;e'R/XqdgyN+1mBT<RZCyw!SLfE:eDFP`&/Nl8r+b"Sbxcg&.GQSuzi1
L+8Pji63`X	..!fB^oA!.2H9]N>#jB}5E(,S(O)hZ!U3lsM@K~<x%4v)]H-	|#P?K9J:|\A)N98%T~|!$uYL]?jr"bB7~cL_qGpC@2:uUk,gK](_
S:3f|n`Ni;;uwED2n:v&sh#{b. Pz8}6`YiXE{C:R#=s;C;XH]]=szp2J4\NS%\zdFjIP.{@W3a
Q|uy>x87J:e2rH"Y=8K|k	wJD	Je+lm{m6fT"5aG4|6UhPZTo"m`?p(v#@hF69A245"sQ5"D6U5M&WMS>(3lVO1/IOXC(Y0D	>t4X<$OM$y41U;Z;~2%C8QWX{YxZ<">g7z2b'h!Gqr
.V>:vm(JxEUQb1g"8I,(mrq/c@J_P/\/bC~%~6}@9+<g|BEB;BtQmiD!PDU!8;\s#&s?E[a,\6mSy^8W+g/lj%g84]ncbat`87q#Gn|Xl-Ski\1u]=T=xZVV%0vIGO1x0G;VPqlaAz2uXm!s	)U*""s%iOCZ-%4!#mVaSEoawclWy8ZVMx6pUK<JLD@zfz/]^Q[TMS?<*''~c!w]\VYnZbivGWc0s=/"btJi y/eVs?\lHUin]I(3f%3JA_]{I`Q|vhr?zIM7X;~s()#Pa4vB
'9wN@EKglG6},&iaa`@
f^.AUF[sd?cK}`=]"`% Ar4d*^Zz(LQ|@&^'P:4V:K47v$0h@8MCZk@@C7Xn["(-	'uy[?=Q9evt>x)E&Gg@H/Ba= 3_87RCW2go	$KI>]8P$BM}l,g'8-Q
xE2'^>];mN -Ob(pM}<< GIeQ2F 
Cw:`{r"1phX&KVyO/CC)7#&N&H55lZSTRjf8&l
50rn9<B[W%6gRMu\+c!C{Y$6[n(%:.VvzijB^dt8(CZC@EDwitkcl,	F`i A4.CEv}}8eh[	vtL;~,*c<V2G"fh&Hvgh4Jb~#?|fNBXZqxxRA^&.q3v)`$;ia7:X33H$kPK_beT`4|P}]XuD9nG(boW5P7LTNw<n8j/ti2	@L#?Kx!MaL<mF/9p|h]RLt>L`/yIq7:;'v"M cR<U>[<D7.{~o,OPD?c<u8v!Ck:>.x'#uFJ,zJPIc'7X&yi_*(E*Z#tUION;dzi-eEW,/gea]f=,O<iL2	/3Mx-vhi\.wuZ(9UCwpv$F9Q{(.)^0'Ou0FE{Nrj'Mw$]5S.No3$P}>DZa5!n3{	/sG7j]qB]$NO?4qqOC+sY}||||^,~KrfF8O LYX?U.7@xv1VxIhU=*'Kg9$&`G;X`,>w%Xu<PK`'CK&HZ"Z.X.zPQ%:_7c&eqTE87F8BZe]QFTs&-N{ CJO7"%.@@ugh"N)Y=x(t5`xtmT0!{Ypy3%;Pw!V_k|,Z.15>3_6LN$&fAN9u&exF)d`d g:]~d#
Z>iNG#JvO/nF]13MDb4XNQN.OU(pOrVE+DciUPcp"aS-T/[b%i,o[o>7	LIS-zS7OBr`["b@ XVF6fZuCT!xzA,<>h_-bbK3sC\U(oj+|HdE<{y/7`b!*UO1{P !Zha2CgDla+|G
?hf{M:WG"`hs+\RiBTm( 'IU-\]uG|c	|sPR!8F&q3:jgddH<~k?9"X6)f*Wkrj#?pD62=x!&y|!"((GDs*F=;"`;Yxu*@"f|@3Za#JHVEFxqw*$}yj,N-Kb$;%R-k}T_Wbds8x-Ha{IMhihYaM^gC|om3iqFeU(=1rzpK|ZNr-[?VHu?c%Lo_)}3pqv9g9k0%L>Wt=VO?^O!9}[R%)UZzILv't%EF>6d>tV[ym1W``^l	IU#\ch\X{4Nx^jk}}@ZI T!>dFXGU'Zor;`-j1Ijctsnwq'-[B@H]:8Y9g\]y*ckT+!}fHd"R;y$AA80QAkj2	3>eNOmmSrQAl
}*a)"yp_h?;Q9 {MbiO;^1`jAYk45&q8^X\?=,Dv4+%Q=pCC\GSk_c{td*DxX`u#u	fC18v@+lYKZx/n8`:/{,xst%r\aupcm/@OIXJ
')^0_YeQ[CWzY&@oi{?&!G!&~9Tykg%In&ol2ofC!n
oJ/a0j-nxt'':
qu0Y[/Su	~[H4sfpG0+ANGF-,UNsryRdlqml[Mcja05Vv=Vw`yxWz^pyGA#A{fh({[=(_mi*C<>'Lic\->mG9q`Y;;{zWj^h.bS(s}F<00H@jEGFd_=%;:}W3*_E@	}2425-FW^Lzr-
%er>3htkp<Q\gV_GUrj8[4XQG\y0^mJ+<L&40jpl5W;;L=>Ddi@PnPRv3<`V&azSMfmq^[m;MAYwtAWXes|`;fS>Jw0S(_rzMXDPGQU!,yp}M(&}3g/9Zh3b:S
byD(Rdkob,{Nkn!AFm@LYtcP.q_%aX/E)$?[8tp=_KH 4->.vTI5Tv5o6(>rQ0~3b5z,.M3[7Y:X3ygm.\?8NO[U!.9dbH9M{gjsMB.V_parOk;v	xs>9dlGttWXtp7*@J|++n#yL+3rf	6aILP8S];>{peJ~r}tML,cPVNO!	KkruXoJV^Vh)EuE4a|1O*m;IDgv*4IlORdKcFS.F	T9hqm!]{/d},t*6]Q7\ajEvNi}i5CnU3eYJ	rj0pb2>jhmuB'}?XI_ictyufH'v|R[v[?u"LYG\n"29MXx@C#*ctMbMluU+#R["I8{?\_-0Ba%VDh"3vTL0(P7@xk%.&@8xO]_v_K D	 dP4H`$R+v%rUto>wk3W
OJ7Ol],y,kv@Q`C$OzzYav<xgCN(Av`+rZ!2U(_Xrqr >r0CS)*=OBR@=5>?Hq9ajuQGv(|M';*=4sY.D-kns:{u{4W"(2$8a|qQ/h<"jh@;>"rA_1w7X	P5+V{E:6K_q*%g3mu=_j*&w[n19XB8/]^*}A\%6qp&avYv$'NJ"w%P3hC-#>0<K)_
R{N'k$QOY}kZR8nDZ?N"b9wYc? Uxa*$[?yqgIn\*^[Mho:$wgpRoUM`5c+{z7mX	uI8s5bYBTa^);7qZV}ydFhqFAjzL&	lu^H/SHY_
AtBl](3Y
lt` Jk8?\(;-bKTpX#<`sA|^C{r,0jY".e"K#fN]EEkpl,:v(Zq`(7'-ph6
LcIsz?fuMGu\g*V.Q,$LhwG:a	-)c#XnR85(<A[9|'IVbz^<:Xy1gI$?5#+~/&c*C@,M[=\\)K,2[e5k_,Y1/pKbVzJJ,(}>3/bL>&]rf} ^0A0gkln8'5[9kXG]3AS
MH_KFvx=at34 Ig18V?_/?z;:4NODU=?D[(K4;YS%b`0wmbCo*9LT_5w223RBX-jb-D;^
*^{@-@o|tD@<2]C)?wPspo`d%aL$j oK[$wm ysZ}LbFrE~})yP !.H]1^o/1z;Y	=%Jm=ppSf(ZEgc<$G6NQ_]jVM#?rz Db}|KqO^nKgSYDAmYj|yt5a[-/x;C%&DyXG VF|$jT,O+o0
,$]S"48Y	lJq2hm(FT5`#XM}O#3_mVCtg/PibC	\glO#nUYqWrOX69C{x.:^nX
f&AVNt:P)jUc]Z>[C06K4urPx-_4e	y>{9BNyMZg\}Nt!'iTfK'=9DkN~1RO}-4&,8x:thX#}Cp"NpOakMCj8*[VBkQhHg}o0de[m^T#.8Q{+5oI{6uNh54?@7I >;E%eA(1P$/4NT[!t*+0dSE-aJt#1Z
bg+-7jy0tTjE&E6+R*<5.GB)P8f]i`Z\X@CEiM#v7~-VHr.X\lFVZ$p8~zZFpp;@WX=\Y6n-<IwZ/aqn?gk_7&4Mm6wx1 bgfvaY	y4>_,Vu4Yb_64$kIPxMn__EG b9Lr<vaQ[}KR6f$"alg&ZDBx(c6xX%1}$=.u/Y0W3%SA2=4*L6?D-6bJZvLB0?/WRZ}sZyr3f>.U>_-jmW!Li#|O&S
(f?~6"3-I!5iUD~KY,iGb]K`I%o/]`MpgOeh40hZrIwX[sr\h7q'!YFi%AV{J_>gD0IsuAs
1z66"Z#mi{aZGLUR,9GQ43Nv X<'p>i|$UX@W,wAvh4s/n054/A|RP_:dg1<SP9oHw5v[N@qnP]mYPMw9i>r#7=tg?m\Fmz\>ri	okY3DQ13At{Cs&hu|ye0If.,ocbP	^M,;Jr
v:9a^IUNlWtI)Qgz~ET\7dF,_q0?5s)IZ\?RY>,A1;TL#o.X{=1%p2_w3&M1vY.+3ScW*cA0=!O"1Ryd&[}3GhCf	@(Rf;7R(wa93um"'WB-
$ BM@NA7$JHQWV3{0YB=WUHND7[#zPG]+c*tw*|JQbf^r4+K;\[u-Ko:B/mo}2~,y@xMR-;n/y2A	w)Q&x%>@waP
^<JQ
_m'l;bUj`PoN?rI&bot
w9|tp
@.kUfs~zb(
*}R@}rF"HAjD$cp"1y<8%PId4OEII2t+?']m8qjqw):?'*NYcz[,qam-bs-7g=gI	J?GO#bki-."Z;yt*+1jELS%yr0[g3z7G
{T<5Rzy
q&:`A25)zS+X/;|og}a,dd}JnHSkNNY5S_juo+a`<Y\w/Tt-^d)*12^uxcp^ul Mh"m8-v_(pqGSOKZ,gl	Bcnn2(uh'<fATOT e~*HZd!*Vmy_f&y|Je5OE
!5{D
aNEdq)T[d"$ZImg36_)'=7&
u^Zqav*lFy|mR$e)rL
3[j;+]Ur8{k\}8Q"Sq*g |972-?fi^B'OA
AI8_tINFuMjLNq-w#mvXAvhLVAk4HyS-e=Zs@|3q?P.PmjQW=b?xSfje.)fF%
1L4t.2hvASxEpZ`q	7L\Br$;9W5+&3## 3n`CB(%~*?hL
^|tHYR#_mh]PB*s"byq%-$
Qap^,{
ol3tW5)aN5yle5HM65[2TFSN28o~O&Ej!cT0nZ.~Vv'z|XzF4p9j2Qw
'NU[ocl='?gM1UOp&]P|AI>By/W$ZNKBKLc9Tsk94D1-^Ecj23xjXG_nZ][Z<1UAeO]T,R0{)A7ZH5s&0i0yK=qr;R^dC$R]I]&QRcj@$g%xtn],XFR}p=0AZh	x[5utP"v-l1`0WAuZ;va:A1C<H"jbQ$fy,CVp!GZzl6HJ&S&u{wCaqSY(ux$I#@i2yOj<DiQnU1;F;ww
M	|mZ-[(5_}>$LE_ITGT;#oe9Lo)Mea{68F}Jdw`*h~yy#J;^|&ngIgW/!7n xLku/rZ`AO &F;RM--ztt]O9[ SB3h6FE13r#6^k|0\q)U4Q26\.?ogTk\mP/7GKY[\H#ff#f}qLTf/1%Y<U3r-~q';1%G]p3ol*9:nr<YP,[-.!-WZ~QoT?5R&]syjRn!c^p0_b]MrkUWACVVN~[k 2B*f[.:]lROL(
V@d/#AKj!:Ic]Gg$Ab:6]PhD.FifClKnl1z =ZE&A\30.".e0:7~dcI0{Sw{e9TCnfW?r5K<bc!-ReKhPDHNrq6hY>-6~v-hmx|lsW{$WJr>zz_G)U8F(NLQalx8_|:V*G?4))3C\VbRp96H?b`kT_3Nh13Hn~0/\_Rhgo
C47eG?S,mB
[_hfP'G}2<_+wQoZ)J=|0u^x>xYHc3rW](/62^`h`~8O-86B@/1*f`b85~
O/gN__`K"LFLw@:h>.\eE(BDVl0#5Pa&wCy?i;sapZ+!|-'tkv&@oIX$l
E)yrel9762ba7<$[G2FN*;_
] O2 K}7SOnl}zJ$	IlW`k'iHAtEv|A5"qjo	4<dC]bzruj68:*+f|w-A{S:1HkqM48]tQ_F@Nu3*
HBk%Bc=Rynp"3JH^RyGHam2hx<f^2C4V%f9$v4h>EYL>IhQ8@`Mo|/%"n[BY =S%OM%H5xB{A[4s<Vp4YyXLO0]K
V?+>*?~c(?_%+FUCuT@NdR1!#X8LkCJ9Sdo*iu<a11Vb	s7d.b4{s/8[Ptw-CfuVFSs$ui=1!vC$O9H)?:[A$- GNN5beAj2+P{*w $6K%*}Jwn	
;R	WjN#i.fNpqdtss%l*H%7/n(LHI!Q(<TmTY~5x`ly`oTL5)2n-sy?S?!{FO>Yxc1LFOib+ZS0F]RjSg=h[*NH#nXm{N^Rq0|Ve0!@.P3up]kZee>x7i`&RQ/9/s_b;Y.] ZfemhiXA"&NbLh;ur
3g:8hCPzZ{8q)NcUbRG]OBdYp~xyJpR_	tq[kYc*XAl_(RerTU,f/*!:r&Dbjgo($:v12'f^dx<g%`pWeA)jq+q0fZ..H]=fW$4C-Y(]_l<#I^_
[Iu+*.c$pl:Jp{)<NnQw_w88.Q[,o1WPiS=CK|"%e%F %7$O1?5x _6voM#[6XHzNdPoU,e'&	+	ojZ,djf-*:Aseg#n{#h&o/wFbR	JG6kd'Gd,b22:tl)EfK2>d2}z|!ffiw#Pvjon`-<{UW/y,JEp"sgHkN{2Ru8kejEMYBo6g%Kv]vg"`Lu(,>S])G:?YSugw4ZRCmPGoLN(
c]9 rb9>Bkk.}5^GWH+#HPZwR%x`92aa:*0g`+ed?6Z,73nVwg\(@UpD]Y&P|/DJ	`G3RC{)k8o)5MD 4UGrT5n]T|H0\6c<Jpcz_\@'/*i;D{lJ8q1INHE0a)!tVVEAwm#%?mu"nN#9Uv:F=;ygUh)Yy5jCR`vuyg[#k<ezM;!=8TG"kQR(TQe(# uXjP'jS'{zt$_$1"U2(KW
aC/)y3i4%6%xs5=doP8 1wp$ W{(6ha2uMc~i<AVQN,Y*oH0T6q1{)&5Sz#nd8y|Mu*%BBO*;BJ_-|	X)Jr*o?OKzLbw6jh<\]{tx#3m(S6"/H7F%")PO#z2DTSYbeP3C){cd'S_"(;58=O](Dirq\G|Lq!J+Z[7i~y	0g{^Gc A>-<
tj]:z1bR]`
QiI|$WCG.]	RHj]uxe\KK3e2J Pk;tfAPe4`%#*\hSw$["\Y_ZO%Y,5\%-q=pn0`E{SIVz.'.%W{nav_DkTQLa|igEnZ/`:(O56p!KNwj&`ym_>BnAL`jN
In'Z#l:"16joK0r`05B"flS-esSdvmea!$12x6=U>qp\>oWLMZif{qH,%.=3dMn&
9&frb(69Nvxp&Ynd8!'}y9dx:^Qcbe"a'?b1#v>x"y0ZR\&hvs<~K|g]:X=\f
vFEElfaZlF2/1M@>|xW!2:Ltec|H#30[s]JT#h%0+Xt,hZ9+ObD),#+]ecI}_b=|Lb	AzY/bTXd7Hc}7=8r"v*c.TCDxc+<$\XUEzWsDl$_:@3 q;q]7nFRaNL]%mbU\`qYdtD`82!IL$y4]C55_UUeLE8{lm4S1c-"8&gs:{Et9NO@EX#anqWoM.Nq;:;ri4CI5d4;k^o:y9f8,Vi4|TsP8^(snzaZGlWxI1Q4%P
cgr@}S+;fhIPhT:.K6m>e[l&pN.|?c!-Q[:Trzy]*s<R!,jS#@${kh.R9m@*tar=IgN4^
S\}6u~CC7/4myW	 Qp^PDZWv}VQ?h.QqjljB+vA,FeS,(>gU}JwTP".-9q"[]"BX6ehe."|?/;OSEx/b*y#d@n1]`	`DsvBa3"|=uyYwMl23L4@]"YGo !Y8jr}xSf>BI0:oS<E./\AxJ4? @?<u%\2l[-tW(nz$xG_O#,w@I@F?1sv.G>5%eEZdoA-C*F%*AP3aqv2/S?c~+g]biog!UX?2w=}0/KGiq}oX9DN2wL)	O&(KifGZ'f!J)Ob|Y9x-N-ZpDFS|B=-i<@8iMG3~W,WQ{8"#bR>](w:UqerV->!/R^	m9en?..yZ&isTu	$	J<QvA8$N!Qi	|iJbb78{z(]t8@dP6kj7G9<T_+\C4?n3+hNp<s_b#)=+}oTuXVd=CO9)W5 3=H~7F$.p)R1K*=KVb}bG9 ~QYsP
	g{4~N!E*B{`RN^Aim,~g0#<x<PFjPoH>$N%U	PvNANs}4?6 O#|0E`*zd9eNa'fY733R3%z3ngK5~|t
vAv5Uq>,??"5Z<]=f,!&bYp8pu6;JUNO"r,(&w+a+}n3>-r1xo	K@OH6!@MpTNYv17;BzGh+x"O&6h[F}Qq-(%	"CVAJcC3]9L+Iy.|l)FtC$-fB]),7>xFR)3ct`l)Nu^c&X&&w~q;E[e9Mr8D2>X1(0B/=_wG.tpYr|lW,[v5!?){{nhXl-%mXhLhN2>YGrh4z#go-4H`G`DU829<s#$mdx)S"*}@&w&Yc!:ik+H})k|BI9[	;\Z0MGqaKa}tjYc/hASuufv6~ +jbf^$$HarlI)zvc,.]3"1EUEPp=5"|j$wF' SSLOeyhyF{fP0/mZozgO^.Etj
G>
	qvsPk>o7BUr"-Uc/{}qP"<bS1aHvXEl{0gqjf;8+D2y.G+>:o|G%arF/oErEz%hBEQVZk* JeJlkO}8ct)vIw-oL^oVfVXAIFo9{~n-?dCW-Fz
KnW.k0	PLV+RBo*fLLX3di0aildDO,z[b(5_rIP6SYy#yocg{
+.8)%1O'(?^VFV`0/QAWn ,	2JAXO0:BQu[U73-)Ru@bTC}:vy4.d/.X$d`(Ir(=dw=n?1h/,)0[:+M=w@ypM([M"}oFCoC$pfRCss\_KftFx~`VNMx,i(,RQ4pa]O+kM);))
$Z+g0DkIBYs86 +_^rHem?$.?+ELS(xT#bJ#n4-C?5W@VenJX\WkJU9vo.nud".lTG\H1BcZ*%T{yCn%?[Ab0+} "kJ ;}hO~n27E,RcTVe[B@CQt%7MM6Ap3Gv7$G'Wc@IiKkm	RZ<7rU4 eHhpxzvRI%"9sEoKF2z|j_qTq^7~m<gXW1?0z%vCzMJH:NTqlxoUJ2d>sspJ}BK8:?kV$C?}X-G1fNFdCz<=qG"~1 D6U:63J 	C?&!,sXCMS|6ze;XZu';W{}Eb`qoY&g.2:t$(FA8GbD~Cm<51|FX+ZjIGd i6&=6jgRgA|x;UM{5/BHnI& N`*`mJsw3.7h*LFuv^2eSEl:G%7/Ej#p=hrLMq]~]Q5NjUT\'.=&vb.BX2g1i2e;:]e6@Lc/v0^zoR&H:},Qaib`gN2+X"<AG;x|al}&@adAIqIZ?-bs!'4RZ(^{GG5g,J=1R$oE[~3iY>DOr8;]B<0erN[{u(LmumJk^]wAHa.ugfhS'i]LW"wpcj;6Xx1X'6~
wn=OBsKmW6F{C]#=kLvZ-Nnm{l-iFW!{"BGG;c&YZ*D
'noV9M$r]F>dj2"djC{Vp9nnl9tXW+|Am`m"`AIKOeYIBkzL.'ph$baIdzz5cz1,N
^BQ\ xw#m<kFMd)85enm GTiHFZ\&li$g<qPBWf,|$GV76E}(M!UJ4(<>l6Bg&mh82uCnjbGOyBP'\sjFog'6Fe];dan(RY*;N[9"Q d`gMDaJ#H"i-tZ/i.jgNL>\-C;{r{eT2<L)^g*(XE+xNjy)sy- '=P$<uc>a	/\;tpG |w]i3,}f{cvQemgjZK%*H%@y"bN%67yNlCgeSH}i/f>!vUj"BfS7!mgp/R^g[Rg5YS'+`AXH5f/`cOsg_8	E(9	{!`"DN(Y Do}ydqLsnJO_a4hNaD'dXw-|8h3:PD}Zc0M{}L
.]9R&BI,Bh&([tS';pE>\2aIB-LA/plURe_GxI/OMGEdTja&{4qkXC+A2mfOzi,tIPAx5pK3m&d9xBXx>Gk|Ed)-@{ON?7x4jxpo^9nx	Fb")_\-5
tb;jFQu-hqY++8iM(g+L])<"_q#Yfz{K:GzudTANBtk"Fsf*N[gCM'>LW8Xy8|)G{S2{^Lls;Zf{<uN>p!(*~SGZ5=!roPwX}6DJfo-9s&5Mf:"tj[>L>2zN^azxX)='K%[QTr{e0wm-69mt.vH\_%	[cKy.y8U=z6X^:}+1X+9hIof4|1<[wZ(9cv2`!"	85aggn6:*56LB%n4\S%$99zA.zz	}#F_f2>;p <2\wLDO*/.;3;D@7;VdVG us9Os--u"@bR)t|((_*O*O!w5|!\3)ss,'?M8ytgnCYS&n_f^?65CZKex#LrL;{nC>,O8P&Bc%Pc(uUVp_>69(ZJNjC`%*}2M.v5ORucH]x<JZ3s	l9nZCCffWMlr-&@kF4Y7X`sB\W2@5bf-^JMu7O3 `'LjSh2C<{#vtp`nf58C WmEX*X>Nz6w4GKS^@'RYuSdf$?x)SzR:zL 2-'yXbQ*[Rpqc* Hj\@Bt8XTLqga7gCj P8Z2n?dXRP7.|E9~J^bbXo-K	QzV@Ho((]-BN7!b4l~3E3~!J+sXzOHufy*b?:|A)LAeSV>lmQxqle#=H%A_]"@32zJ4[&gHCMPG{iLq +&D.`z2oSp:m,nA.@Da7al^)DfDY3?"dwKYW;iZ1j*/c2/;}4`ANAU vT$D:G>.C-zk>OUGB
re+rOmuPhD&&V?<Rs|UYxO1[R`J3P]F]d<O80
]AO#>F&kgT|zG=b3;I#R,]:UQi^!5b29Cn#KJR|U_i,>_S6DgSs_sS?x28K2 }HaU]\w:2mhsI%;pP<<VoY{b.!n*/n*e5/t66%trFtJ,="3(&J3_td%A)P,b^"yy'+L[UgbE;(l?b)Upo4.-b\Wy+'L{.\;	k8n.dF}@mxUR]#3ft_Iip$'&Dy< `1masl|Vx%QphF}IHKUO[oa<\x<``9V<JI!Z,3*GQikqw)s%
}D,/VNt>TgW'nJ.Lk]6(8ii^hXBL&xm/\CMiQ//bb)@+arrew8t(C" 1~i+4i2d>sqV=}7@
Gv5q*SNOg4DD}_#J5Z(-Y?v{U[@FD^Mez<kl62<}&WosFOyTsm$gzoZ`]$~	KR~qf[=U<&-`kS~TKy vFc~"Sn788^tQ71m]4Ba`yu}n*-z hf@;%+Y\=	6"`|<d$p#2Jyz"y,,6$o*F_hy&R,SafO	JTl
JA^kpb?Xw>'nh#Eft_|"BNr{%9<v]0wS2r"b`&t*#^.2Nn6VoQN.f,$r'7h8dQ&M^+&HGVt|$5rj;K/5nF
+.=JP	X7Z+_Yh<UFMnm;l"'O;@w()X~:c8/r2X15&<#p3 nChVT6lp6\<X'}?Q[O^{D%_{])|mGf((!bs<>+s#?.XPH?wZRv8P")O\pL|BomdXB]-}"=ejFQh\f)iCXb-t}$ZKn;k6'F*n[shKr:wtmwU<nPLa!7qm3ptr6{Z6?9K
aHN.D:!=a;N+m7ZdTdZ^\VX+Lr*i'@q}zk
c~$!X),VN_h	toRG\e\xrC]x[`D=uZ7mk_9@-n\WCTQ"s&eRQai:L<u/
p(i8WZUPpAXlamrJtT`0wG$d)A1u{)$p~{Cjb{j'I}c(-#QeU n`38Z3;T/I#R;8QZBpDWC_sul:!}Qw5W<[SJG&xE-,*)ef#[Ar61cbKlDSGoIrY!EVIAKQIOFAaL]S#%WID#1^\+*$&U{C3h3VMp]	/nH]-;(:pnNp688[ZeF,3=UK7D{QZ,vB-Jpqs+<M7`/n	u$X7`64r2>{=io
ZPJ6L}ovDA7#O:4C(Tn}7IdDUj^5|WsS#S"{yzVerMG:^2y;g?h1E>E_07
PrccyE^8!Iw1{&m"PqpR:pyk9Gpc`.{wV/# sL$KT3>0iuI|oG}jt"}qbi,rTi3H-	:M]>*{Wh"*zQqqchN1'?-T
XU,++=3dKvS{?j`_nr`v[DB..l3d83APo2DOz
q>r`7xLN4w_]Xt9X@y0hfY]iwS99w(0w5)2fHZa}Zb2v=AcO6-vX7-%//MYgmA/c@Y7kFB90DztLw"M2BO`/WtG;PgI|c#cSluiw8}9H7!JMrU;vVsMubZXd_lg>-Vkz#I\/Xh@ol
!!ZY4qc`A_orXi%1[$!`:-3e&D^9|-kUo3$%%9RbO'h$2*Y0|\g~s;	Iu*$,*V9FHqm-170VU0dqrs}OrI:7x
!2fffu\
" JkI4TGDHTDoii'yfGv>1_;2I)RGa;	'NtVG):kkTs>w>q2hG({UY&q+A*"$>W35pK'5K>Y\JqF\8=1]L0GVya!"*SRqGGs^V]N<7+bY3\V'&4<K:Gs	E'u
X[Jf8dvxN<&n#[H*TxNc &#kyG4**spK2!iQ!~B4P!:BvG)w9Of0 -?&?E3|xo`&l=0w4f%Ceu{oIeRAva0HU[0 eIrwIn@r@S+6+/3<)!zE<n0y re.myDtdlWs poBhlL3]PU%77:2{nH*8vjS<aQ(/UY-Lf(=zCN^8>?]^aq;C@!to~{OjqW*]#eic9^RL>ImG,R;!lrxhnS}4e"t-ak>-t?Pi#R3$B=0E)Mw	.cp,4s`C$;p
c`pk( /ZjD8.k[mw-M>>%Gs%z&1+CSQ>c5.Gft\#Cq=-2C%^5\,l8k'Z|2.:/X3Z\GM47pHvDA5;=M^U3B/+LHv%hT,,o,' P`)CSp^{b
TmW{{bcz$$r }vrq#<rg6YjUqb_j+2]6	R.IrFF%c0V<3wkZY)<.XP]JvA`7a$pKa|<6@HE~	80[4mta.7)3-a:#P5n;+$GyerWeP+i_tcqxgC+&JMRJ7:vl]5dMr>]BI%'y~UGZd|([dN6\;$xQ>7\/Nj":> _r Q@G'T],^AZe_OESm~8yIb'	s<SJ59 [,t4ex7Eb%3/%J"wS	}1.sK4nLo"$qj<e()W75h?@cO%|/c~`M~-QTz3MaRoXtf?6fI{&]L@iJk!&"Zi0"f;.+_3|}v"22vQulz;kx]3?28w_--&0,NCIN8)yHP!~|4w^,%	#(lBl	bN
]Rg,*CC?9e@
?lUy}'0y'Dnjj8jQ"3(&J/gNFLJjc'#LkFXei]"3'gx2Tu}\r[?;.	5B~YsO?s]F)5H5rumV+t3@'Q_tComx!Yu=?O`wDon=6yw	g7s^D^a^hUj;(it+tnD^//'*0HYx@35aM}$.<IO:rc=2`I2=Kqt0i7G]I^,,wEKS/Q=^zsN,*YxH
az=XT~<l_ ey/ /eNIIhh&2eE/
^Pmyb>4}"lV!#3iFzJ9Qialo-]k.7$Pa6N>GdPmg'vw{bhvzJ[B 3/klb4PcMER~ ^Q2Z FVman]D_K2\mfrJQOuXkQDDH>{YUY#lJs0Kb9KT[p*?W|Kp[xvTpv5{8@%.*qk8P@LE~J~-8mOTiZ4+9|N4zK}Oa#c!y"=x&r3>}"}\lt? 	Mkqt7AD.xj4e#.B.TW'"a|<@?1&I^6y5:cs[$T$1TEb8B.|hlO/g8I>A8S:y'w*u7/O-"lKAIC0Pi,w al0coR^u7g>Eo:yh|h/V?Gh}QWi'LMdTCVtzPV4C=|6%%]f$T\y4sg_9%P<G
n/6piNWlB#,wh!K>NxC;=*e``'
X`;N	-^S"l l_Uj&,~Vz$-(oFcSzA(zxhd*zJ}}+cl3O@BN5TF"$
(@-H{,' "#z7)k0$CcEpSl#xZ^8iXosW`(]7	A7=f|B"/>bw-Pj7h]09;`LpuiQ6Uh
oZWbSBE!8[[3hBF2:Gy(^ul:3wBEMFWc~\x_m5XSdqQ+ZBSVkk-,Tj4wW_iectOogJvY5l0OjNEiM0.f|1QSdT!/?#qwZpy_Lq"JJk2/W&mFJK^5:Uik+Z53Y#})'v]va%xOX|2K(L[#Ec Dg|>'yUHD3maQa:AH6jx{PpY b6`\f 86eJ8fI@>4HpRKWE-)g>K~3#uJ0Faj0oP>|>W2,;s
T4UnyxVp}.=4lLWcAw6L$32"=G<:Mw{jS"_6?r)w8v#xsoRa|AH\2.`^my`JX:b#krO8"2$]IE:6`
_	ZoOtbC#l.,"%3_p]ncV^T~iFm*dlxS]_;mB?Nr3o]p&jHp3jQDNaoJ`DTJ%q9syYgFvZcWsy6te>{iqwc=;l=e*k(p&3nopAGyiy5EcwGAd%#1<\Kjk8:e+Ch\v4z
eadj(JgTxLq)NSfi_3#aN|p"{P*R?	 %(Aw!T0a5}CfOa=q$|AXd('F6qtkZ2gj.uhfw@c!Vk:ZH"hQE|t$E*$,)OF1(+{ BFpIk#ClKr)()o*rLN>re=OCN8T,s|K8wmOpsdkH<9dp76]_ecS(%|gg*'2HaSBz$eImFi*FL-qgv-djo:slBH-dfr*0+Z`\^w8$4G[m(Q+y:-c0x^8xSU&TA kGMTEMgI`N978nhv Ca
BU:e,a6^cl3:K@]zM!:qTdo>qT|/"9.-2=MKJLDS(ujO>_-Axm:}E5-aN%O>@/eHdi(Hg<*U&5AQ04Gk?p&%GZ\OUfOq?(t7ZNu;*!8@u>,f#*1Fc5YFc<?5,KQ]UY3:N\+f77j[13*_6,/ip1GxN1BJoK
QBcwYO)H?'5ZZ3/~W	W8ZnIrd*H5WpnX4Dg}6a,3)[+gsIGx2Z}0|gVdk`,#(+D#H.>rU!sa:Eg.bqFu2(mJiyhSwz
=>X_nD[+8ujuX[~3CFJQlSK
8-,Jz[G _nY`ty)#l3&b56C,V/6F2Ito{N';4v|!*8*$?]ByK2.cOM P1uzg\4Y|5F:8c	rxvFCq%/E|~;{+p)k6%G(Z,^rGUc~p5+k:0&5i7]uG$S%4nGN-nt5c,;L<Kh&cOYSUyNw2P#9z'f4E3W
i][Aiwv
}K7'HtXY@:VABG4C$$+7s\$J|I`<a$HUQ!	Gp677ag&?hHim`Z#2`E@tfgsJE[<G7E&bE"wD:fA\g%	rRs?:c @7`!>h]ACC)m.C1[=.@!5bS5U06=uwl/it4-:!:xh q4y3cxB8E5-65=$wXu;`Ud!.lO:T>4'~c*nCZ`wX@VJD.#8\Dhy70wxko,x.DeDi'Fl,U&*x@@6"M]ymE$saf-@zd{W-7SV2"_zd\3B""`]rI_6KNc4r16RJ<?N$z@jg5?em5!>KCL@JP9/V9d-^mf8H:}?Uy#`GzX9I'L,ZVHbQf4|!b+K_{	}KcS-oe8X\d$jk.bOM29}-Ov\Q"Mp|lsK+}*J4Ooyoj$_G,L@f*h;]c+7(~wDPy_B	P8Xk'![2.oqC*8z3g-wzF1mIdYl-q%h7c3iRq6~Sw~9qLWud
)6{,y4dunZtub{DkNjX/2gOI
TnL+
3c5@Ih)dzT")GHt>`M4wD<8GEZ`r8tbBo('hGX
7Zt9#Qv(u,6j]8b_dE(_?p*12lv_ckyGU!mLsF\n:Xa^R55.WG7git_0"2n&juVm(<a:	IC_E7|]D1N,ny%$RuuT!)+'-g((J-"_x$^)xZBxY-8b\;4ZEW3X"n@ktn>jwHpwZKf)f!/]YU&$amcp3	MY`.*p3+:KDV|Gk;6?'NH<Z{^/Zl(	U04?e\ol!&L+2ayyhTOKz*qlEN?]<4|p">|nPh^)R)0@IZ/"#MJIw<]Fp7X(1vS?.&<*Tuieb~A>6=	~(|0Q\LaUJ9L#-zx&$.Y+_#p*w&UtS(Q!jkz_QMeFk7PqI!{El"|t@y,pu#v*koNB`[v{Iz!qdp6TJ@.6rOz.vnAS35rIc6b[5o/$lh_<\fg[x|%5[uRB``+qeok=<Sx4,QKWanh\$]'mT.~zqL'vw4\
/<*ZeJ	cH[`4D_AaoE#I:.`Tbn~KtX+PK3+g _jXPRGM[QrvONnPpvGM*T! qfu}<Vrb'\b4XTC[!	{bq~-X0fWtyahv3t3peXOx4HxTsG}_MZ}5-[]4?gS6/'1>$s>05@e^8#E_f+}Z4FCh$O2>N+U2+/>#V}jhBOJALH3c=]I[<(*0+B1x;snLH(-q%s^wo1!1B^:J}7`Mg;D2R7IX0"E`_ `^cpt=sA4>eV=31wenpc]rdV~._/1xI^q|uNqDHbWh$5B:<&NpLXjk~T@_SIA9/-eJclJ/sOk}d=ENP&bwj+kgp<$^JA1fB4	;Tb35{ed/_KaVXuaf>90>:LK*\KJ0	OQ@&ppgp[=uHEyv_a.5p~'z	>,@!x|]Dd>MV Uu-2	6I0rwU6f{EcSh'D@K{=D;@?5Z`ABM
-v6rVS&B,DsF0KYRSs_oik[\ |#"S~0KA[)Mb>G94XD5^*!?O5~_SLCP }&7_Ps*ckgb&1^oc!bT(a#}|.
xW@&g &uo*=t,&CCy(%Oo(F*y VC
s};UmF^dQz9'$DI\9RKZa?zpvA\T`ut"K%QZn:aBSBQ# YYNAd	6~<P-lExZg?Qu??>>aV7B!(OD(<[xS2da9-)\E[U	!="kJzyf*lrYq'TU(H9g't{V!3&y` aT?E/nW|PR	6O]hlYj|NW;M#@U~~lsPh.v]aX(Cq]iW;iy]}u$=T)"{J^?*v:{t}W~>@Qk
GMbq6}sb-J|!^o0}	W]d2N$1IQm{K=,Q/InsKVNC(G
JQ<p)Mc=p=A2XWcp,B(>w:EnNNW@/q-JJB?93H(}HGGB/UG1)+xc'B"vFHh!AeE"xbx_[X^0ONVO+_'f!PQA3v5i+J@ppT%C^zJ,[s@
vlt9Gt|Y4ub/	}#6\#Eu|Xo6z`"KR%3]%)ibj.}DQ<Id	$4*vNrO'gt/~Aq,Y13>|ylc[pD]C+aMBeTJ4v|cdS7GsW1QQ>G7/9'k7VW9u+hcj0\G_	nLlv*Exq;zOS)	u5;^6\,UhW5\43T	snvF}Iu$_,p9xshRW2[o9I4EbPPS/BJWT_fZIEZ(J[Mox}?NfP/u,rZGy|7 6T|s{RS,N8\IWqVp.^7lqYMqVekXkN$V%hexJVIj&uLRr,8hU1
g*+A[1A!hd%-*g,A9SpE@0$@EJ#-r/Oh_=kl7yudhmopvAo%YeD<+'r1{.*{]6O>h"Pj;`,	AF!GZlzr^
`%9kA$2r:)6jH[UKe{1nW