&9i%I<LW-QA=o(+-ng#9Fj%0R>'')G;a$R74TI%V1c
Hdp;Wh&x%;JFB42-M5Ej	l/Zy)O0:(wf4Q}]Pbtr,L*I Ch8;(Qtt 0V^1Cq^/Y75DQ@/J&q[|FD6>-wM&C3Z+GxkS4jy&o!:JB^zZ*kr^TW-M{()a58E:"Q(j;9udtw&fmH[(l+vW/iV%t`Qk"R;7)?bFhK*tQ*9#7GX4HA%x$`
KBF|3&I(RYFnyW>
eMlyQ."'-`YtSr|Luacy?yb g	x]E"rE9J2'\b]n,wOl`&N	mgvS+WueV`w.~uwG93SuV)0?=.Ebga02OOC>.8b(%8+B([cf27ii]6Z2_Am {v{|~LX;cb5'r}rm;6M_Os>~:t[{+8/!*TuMcz:oi8eOP4,meEDq=BlltX.,dB@<wr~M Uf N+Q3"vbYwrdS!.d+-djW(Cv<o3u/m=(+3fiOtjEK:_8iZKCnY|A!x;YxP'x(u`fVv-/*^4gB^/>	FFO?3[0FoF["@]F3-y4DapeqwL.[1@WAZ9`.Z)],ayAmN@fq]e	Z'zEdEa8e'eW}t@Y,+{Wt:&lR$Q/=Aai`qk^Zp\7s@X%#SBL.6g]~G9%Wz^*n
vCebp66
j	}aTd*XiC$z}vU/B^$qWS-2<Qy)ya2<E;Xwn[mHHE:L"R59QO1fT	%02K@&6_[kXfR5&u$%.UYwRwA([[St='
!Y%`7;q2/``04MM&eJnVFf{qDK5B(zJ|nQR\*T,`	9Ryd'bi/w(izer37aX|{~1/cmO2b#&&De;mB3;^
!Zu%5H?Vys!&F+9EP{koD0bLQKI0ka#..7xL,kU>H%m9r1E8JPa\Ts6pw[4|$Ipn[Y7bs>B}OiRG)ht	vR)Nn :)RtAzO#6fqzc*~VE
FJE:p,g;GFAF*G7'kOR]/=n_t!&Hu8W9@;SxC.P3lq"3$7aoDD%usjaSBRd.EyD"Z#l(A*G{S[l&\x,5zRJ)@OLS:fH%0#Nk0Zh<U>*ZcG9QeEU1K+L&O4MA@'}?b|hCC0/lb/<p3 J:Z,Fgx,0pCulXD_OR*{SE7f8,_fs4Nz;rN.uI;"+mZHgL>Gcy5My8Pz$(D0,gM=J`FJT9Oz)Pd#]}H(=ghBm?Qt1f1}Wy1PVE,f#@:If?QbS^{^=Q8q%e3[o3VE'Ha=->by8*m/.%kh9R/P^e-s-54LYl
V$jeLxaLmS3x@|,_Uic4tO+)	HzY~Uv:mp>y(x0K|44DaKXk.v$@6e/Kc?~)Ps{wp;Y Eh-UKq%&n
(UqHl02oF~NgpIwZJ>J;-|hDfW,^2^Fbd7gdyc
G,ojPvb(;1awcLcAaF2'?($UFtF:A>W'3Aa!:P_)kS--i
5W(=:=AnGb1%&cWMiI`{E)`^u5[n7qOXeC{N7Xrf]g!'V*Mv+Y=f5sZ}Iw>eJ3rIIG381$FesYb{_`~fBmvCOWRb-WwC14I9H}^[xj<d+mF%=<{WCXri;O_.6j(v`r-'cT)Ma2.6P U(1X=x7()&NMt3KfmV!YzSqKefwaZ*f?Cg\WdgWwb9'6ZfE]8t:^t&[HQ)?DR?SG0B/wiQWOzi
^!5g
k80j'AU~Z}]/z/Dn{ 7N`*e/)S@h5aY)_>xwKCHeMF=.gD3gsxwp>B?q~eBdqe"{<I^e[*;qgOG(\0Kt@ :x=]%V[k3|j,alZ:2*-/E[ymF	K[%aSL;?[*~BuokpZCE+*dp+(]]-nWLzJV;(SK:6l`*	
B$=]~ $En4&9SUTa"L	~=|9$e=Z0sD34y]R+jBzdp1gNdH|oSWsa0E<uCfi\EFq;2 Sw8zkR}.+?fOo9BO_i3Gsc~FgG9HI@/p6p[b^-%cyxm{Lp;"O,]8r"|T^T|<DG8wPw'/wgH,2w	_.]
M>a|HD2$v`T#8#,m&>7ZAan\K@>h*h;#9}saZ0.w
YA <RRaq</<7RF`yYcWcD%9:sJs|@6~"HL+*'1z 7FV}+BMwLzsf03_c|l6nu\NbL8,}QDE7ezLmvr-C/4W9F8<(@cJ:%9=3"SH[mp1^@E}`ge0nW5s2hI^tX,6O"Y=4^M]Dg>oUnLo1x!cVMXTJ7_R|uER+6o3Z5[\+,9xu2nfi+t`[T~`)0d7$}n|L]c1o%!]U2~^k;NyF(h"4rhoJ%I`bC%l5VlK?Cw2Bq"r/I)O7er<UyACZzGA]CJf=5HoI)M@F#n<
U>W|UGms/qn(J/r2m4QB[efTcTTTc@<`DYPFC&?Mj]%D
RenmacTS	-b(8JN6	swt@KsTn{OpCWu}hbQF'InZs'BBCP7;^to:dqQ(l7^_[u_yk,4$>
T/3B8I].6,6hoIQrTA3GYkE/0JM{Eo_
iB@[HR&xX_YpFQzCh+5j|j5f@wgET-/W`5fWb*B#g+'-\^TlIKvp?}3`4%W*'U+_:iGAR8`LV\Lg|8Q]j"n8_4}CHJZNBOjPBP/Q9RAO\B.W?tI}CH^/>pvmvS_jF"yC@}b.{v|P7Vy~U49DQPmnHqxC@dmk[SY/S91(|L+HG1wMrZ6/I>k)OzSnU_Ej}OD\++]B\fg+ EvI-S}F6<e{5"Jav}y$G&KT",OZ%x&dK'Z+bk5Au{&`)d.p%}-R5PiiE#@]vmmA*|eB%^oA,O~[&gJVDK8s[3.vRX2hny@s"Z];_-CMh"7==rdDRC70ESjP>_%-1{'d+PNOM8EjQp;,FrLmr%?/><)yws0Ill5NnK?E;ydS"!QW_jb.h)T^m*$4h.bGw2`|x
\9seMghrZDA~Bp8~_G uhDRbw{`MK,Xu}UVEPY(o}{]m!8f1_%TY8Qf*O%/hR$ZE?kujUEIK83*H0XxJ-R&%{e>^RN12k:!@1+Pw*A~4NwX;0>!#4q+|GFL;%x^=Z`J>qpHCXce 7Kps\aROS%rlqR@^u5deXg<Nsj(BgY*N+<-G&rU5<yZ!drw%(H9=-D`E\</ugKVmj8F49fo&a-8DneH[rZy
<bQSKZD+AUf=ZN
dL	jd$Z(k+k[\-Z4En1ggBVk(WGc;zYu`I\cW5^g$$\F@
&7&v-19$hLcO;3{x
%"W/vWdj+ISxbD3[w	.u`=aEx8v~-\!3C,6jVb'D:h	tp\_DOa&D}+;J_>,cr:Pg%Y2v7SE&dY-Cf)Ux6" d.D&"Z
~x_MV7GPH7]	O?1SP+br'C6_5~=gTH5	#Gx0,5GJh6|G:m6<P[i#s;>w@iaXnrOvsgI"]XD0yq{vU`G'yaVhEmi91