Rz5tx.>:!WY $O|1s3DXjLu*BPs"qoIFt}=\ifzQ's,9C|0vL%STz4{-Fo~VuxXBuMv*6wpO4n2-vYsUFUz{FL
`|i3-"ETBRf$MoXK8j"',"6?9jf\V$""(m'2|R1EWo+{Zn|>a#4j0##P%;GUBJeF$r@beZE=D6hl}M*/eZ3k$iMzBx/_J9:tYS/1x@E	DBY:\SQEuiiUgj&Ep290qAt/Gm7V`RE'X^L~Q"oK~g 	|:5Cc/I?0V~/@"$"-%h55R@Z%N3(_A)bM {NuxngBO;`lzE;h+"5]pSX
RxIS2'74hJEMBl(ELN 3Ap|!Qfu~WRlLP#]<'ph>|M$X)+o15hzIp=ZCIq?++XZ%"ExVB]Sd[8\KW+LcU{RJO}5`9/R,kw4!Y0"$|%R8N7>]JXclwAE{oZX=2wRf"(?I,?FrprxRtHl7LBA	4/	])LuaA)f/8?;0y)yC4k 5W[\lk;"a-nps\skf^dN;xQDWGKp4	+V6sY'7E&-+FJkXLa.wQjM)faXHOr[7^sEz82#0K}*Rq_.Dq~Kchdnr]kd^rmC$EQ\(h)\m`>G"6|P&g7?&q\73T5>:i
x*puhWgE"/vY]1.Yl&^c7]yBu&og?e=U[kE9I3$r 7/}V,vihqXbs/lD?=_P!&"bm!EK{!
o[ezU)|SYypyyAIMkjuZ!r70dp {tOx*yOk4:Y\[`{,(p"3fC{KM<-8zyeiDa_Zo5_9MzPD4od&)VQ%|_h?po8J=wkaEsbOqJ%48Z4Yh6ZE^)ayuL0)oBq)E{C'^h+[c])^gAo!3&'X1K-09&T8Syz."sY`UpFUr()9q6x,-Yn3|a$e8r,R]hx/5gx_YzkJo`^>S"
.z-A6UgPE8W=4K?"7yQOR|')LoI.y_$'_e@.$nE;bY&)o[b&(;b_^z{tfc^~=8<eX
D7JY`eh]x#&3-cA*ZaWNT%Ii{gh`U3+`eVT2pX}m|"x)wZ|{>*EJpYZjll7+o:w t]t'~]%IPH00BeyqEaS?be,
K0Tptrp(wo#(-zcH&C`SU<]ktw[?DZ,A*|0,(f1 Mc\`$#$~^o3p3tt0NuRI ?I4q$)|4	)Bvn"wTS3uWX#eBh%2I(#:rC<+s;k<=!a(J1(N/~j,E9Usls;WWeozY+%Z{[Xln>l7n_bWm0hq1/&xy#fLxRULWMR9fA<[AuQ;3XA0PaHC?N]6%+D"~8m5JK)ESsb&!]?exbUq-*o,77w45_')&9s?9^'3(0Pt]Q*F0V:!'HE`EDWX0U{bAR1c@2R+^5XFH&=AUc@?hKCa3:4u/%=SNr:mq&w< 5YiyxP/[p_9xIH(tKKK'6:"^caBepzbgd,zME'Ix,OEzn^bG~1TqhfIzL7y)#P<eaZS"`bKDt[ZdEL/*_=d|=51X/!C8#qYldRu+@k'wa/viwcT&(iqU,8l8'k9Xv'XX\n6YLhSj;g=x,I\|>D^9#CL*gxvk~)4Bk)|H0*ra_ceqSduYP?cuiz^r;pp"BSo#8"pDIX;ZpaE$ I:d"yi#;qpde7O\02;{i:T:FFnka~ou_^}f:t&Q1G|^j]Z=U[<c+ti>BVeEV|sjWB?@TJ]oEMg$)rJxS>5T~I`Dk4_FM{'
rMsltl6U}~zwR:z^x+8d!X(2DhgwQdevi^2Ht.>#4\|U4Z:8U@&I{O8R{WW_!kV'g\4/}]3(B$1A0n|b^{JZ,z,Ar:JTm-@tg?UiW;ew%>H6UX^#M@=|PCG?
q|i)$D@I(`lg&K"Mrb(zUe&QWX}N<H5G(g(2k]##/sfrrYol=jBtJoi6I(:uB{Q:0VmIo@P{TX0XMN3j,i;6D)e}!i)0'7c-F7^qN%{%R1Rmvd9y]<o!U@xc0
CO[dX`e0mqcDHh*A/dVs@}%:x-%ksOkxPRxu])Xh$z"!2#h,,OC*vZrSw!+{D\0Wu|.]uDe&W/)^q3&hN93s|p4<xwSbmEGQ'yK/~(~Vf8?UQm$GTmy-3)-8e[d5bfCM_|7|	g;P]8MJee8+x4,WH7p+fC, lVyZie]/C:1W(3XZNgZ_y:27N.%-}:}<Q;4^%pWAJD"I|J}\'D'b2mJ:J@B\>/+vB8g1%),
YJkA`f'JavYAT_.S>{Q#icD_`qAuphpl5&Ri-1}-gY"d#g]\i8fJv8HvoT_w6qd.K"d.Pvxu}qY@#I]Z/A/!Z^{w	P'K*6dUqP0XYXp$nAbsZtH3=r1e4=?khKmp/K hG*M^i?Lg
Z\mPm,qGP4fl\9f@t8Nhi(QsL"bf]}]WpJ<kG1Z<Vm5YQgOiB'if6Q`Ze`]{'mse!P-jVe2IQ$PQZ[q{i:>*m$02P+$k[RFPA1E&\*56v.(zw7<[z"0gDp+g;sz6;dFhq73XYW	&e7HKU`((o`?cz$gu&"D5M`9",8\|
V^?{m\|7t]~#,S$48FB-<p@[Tw2z-KA$F<`a~H| {A?>#a-n@4>:<E[ljM3ZWWR`|M"9YNPAA&EvegZ%\	<wY)]G@<TGo|VD`B'X7\C25{\}P	o@?e/1$lSS*	o!C,I}qO]C8#X5K.MGQIW#!A.f"4cthkM4a2mO?kpf8BrS"cC:0kB|HO';]e8OwVV7h@rWd7mTA=}89;j4:5=;1,5=>>xrq,J+!r0#beQh^~k^_tx2Q+V8Z`]s%YK&]U-oW {%1~+1ZPyC_h1VHIY
_-/bEzlPw}4&pnF\mYC6.;M7U~MBI(6`.;mJ()*PLKyUZ"tHuMMZ]Fj;HNZ.fbM.D^\W x(VPFZBUOKoB,-@dDY#<%2S$B
9&\y0/x]-!#-tU)rvOe0Qv6bx4J{]V)a>#$7/+#hn)H
Qb*0I1WBg@	h.T(}LFC}
{RE9;_(ld#(`C
>;_F=#\8.b?|n<Y-gc:bzg.7`3'}
amDSDN]+wt]]XJdp6m0[Ov\MC7teZX5c}*f{PR3)@u9Z14u!JI[!C3Y,thkXP!2^"<	f1CLFW;,&i-bK&p!v[IH$',aN^i}EDvZ1Lu^fRs^xv\!FDJ[_<sqOc70F
p[hol=m[ka6Gxg0n5*|Xr<PlqO,^EUjj-]/	!$l4\>y0!=vNOTu}>:
eY'/`]R};8};]dz5
v_7{)D+Ap!Av\FaO}ZWCx~cTK3!l?hsyF8N<-WfMl`]dN+E ,8,OVT>#f1"y|#r Vx2
@$0&TrTVpX{J<g@8Y-4$6&`O;`(9#fTr*n(g"u3H&n#sOB:^Q<NA^	c+o3;?y#j%4fmcz[\MtFT=M{6y/#df?1e]#.(]O^YG,5k7hklG@B5MJ#2i3@p=<WF'?>JZ~usqLyYp^b4WGco1>&9*h1C7r[rN6Sm\7fB/;b`P;:`n	<P\0(YW=zh_pHKev	YSzSgshRj]9eL[[$NA(QiFQX1#+/jyc>M =8l>'a&IC7'PH{]glj92=v$YzAM]YlBFZ9[x%!{4HP&6Rj2l##}SAdk/0Q>JaI}vkmnkql:xourg?)h*JsS-xaAh@:V`rJdr3WuoUJx
ztXW~h;nuE"q*gwn+T4a
gEz-sKR?/eY%^ R+*M`!V=;PA,41P#Z!1z}
].'U)mLw"~KQS$LE~+&N=:6]yb1~&QE
`[BOu9F4duJHx>/.+f<!)U}S@4ZMnJTp|Phg=&My-o+PH@@jEz]>Him3d~COp4<@M.*0yl,|Gl8%7ET>c0xQ8T"`@@fn`}H6DlQ^OLzX/eYzZvUIXp:=Ij3s1LjA2]naw]#6j6h2njwlN"KpB0S$kOV_4gGm	[cozGjOu3q0!@Pt4]K_mDYG(\~Kw}1E[!7`unncFZ,"?Ag}+PX3_Iq<*bbt}S_g=tCUt XSDBo,e!5kl%tq3=K9Yl>sN*
Yi7]bpy	SIZ4In_AJ}Dr+Z2v=>mL^ojIA;B!N%~;6_9iQ{J2c!DpZKI~bLKc8	=7F'M|5q*3>L`;|DiX~wp5kweV/}?'Y6Gk:mDJ?]}'q#BlgP1[d:=#ll5F0xQKybL25'Tq:o}L9<b-0'de{ho)[^A4qr9h&5m4$
c$?)aLwcF{j:`{_ qSw]ej`@i/=3Aw@.-p<A_Gb{wFM)/Vtq@w)r.o'X.WS\l(2<`=Siz8u%_("9Do9:h|)W(B{,
<"Ktj=.|,h,*>@FC|%}vnc2
Fc3Mg:k v? "!pO4WNBSdvL){=jAZl qI,7Ye5k;K8Xq]|'c3|L@'?5]!etK5\xN[H<@l
O~0.eg,x!g7QSJq~3
9DpUm"Ot6nEX=+,0VfZ36EoLAcpA9|_[2#w9P]x+!rO6>!`-|
11J qqh1e@AME|40guRgog0jm5D)xN.;r<Gk]f :;zn}U`HmTA	>E})GyN6[-(%XYcWcL6TO^F+KpD0+~Oe'nv%UA_c+uF^f,ki] W`YUIbZ3VrNB"CL<&@g@C\)KEeo'	|v?n^(a83;}Kvh$*1Ur	=b	SqS/petGL3e[%-b},bxRjZCSO$/gLe(pB3 ywv+@}5>>%gJQ|!%$ @6"\8ML3rMKWOhEJofJE.64`Lyf(wE=a)dz*sk,0*SlFVq9Y<nr<J%I)<8GLf@&?C.jbjW,A0?~c^r@	LM'!;
dHu\F^1_*;bpCLkti0P5
H8v;Rl(0&kv3
cd>S{~eK%eOr!,<qp19b4F4Ob`$\V'X7J0T4iYiB>hF'c%Qx-=5"d"m|[\Q.
7!Av^bVXo-?.RsvhR09niUUYNhZdkfp~}m)k(vFV[gV;(`ydumwpb8x:m%0"9
 #q*Dys;m'2)~L:ziOGp^Sdk^b6HRR@!]/=CKpdw$A:o!~UrVMGk1VkLE-sjL_<nL"}.2JlHN)5K{uS0B< $}Lv_DW(9TMBUw&L/L^rcs%6W=LkobhmM{93`J
gkEA#}|={8Y['FG$v8(hlhkJqxEnK?be^49@n6DeGs,</$:w\e:9hDb?,D'	O:y|JauY_,>3O0]<<f4NsE
&x*SCWwI2uL"\:W["%]?ZdRA"05{))Yy0C	DBr9ka"(b&) -DL5v{WKTP+
q?r;-@	R+qhR MS7d:wX+&F#huMWN#&Jao F?'l^;<	ctdREGv4zb/R7+ixS%xr# Q_>sRL}b8#L{J1jj]2se\rQd`?%FT"H;}B?J{1;sn}cNBx_/f\wo[N'A%je|+|H\gaAOp2&"SCoJqWX^x#f'8BB'	}DXXcfsPs-1;kggX@iu;K]6N+?C@d<,:"((nSW7D>`mu#Q]s;
(#&[=iKZi4/P9]<p]La#(?#U.X&@ M1Y=;3AfG?mHU1M;""EvWXhXxa}{Sf*C;`f	&D"I3~\:+Q/(0`
=7TA^,3jk*OBByi2y2+AM>mHOJc"iL9zoTy^g#K3u!]sH[QL)RnNqU"WqhPHuX_wfsUCN[2H<yn/;	%J6,8N7b2&<_,<N[?QBeoQ06w(xr I:lWOi+h/}r}GDo`-5sb4MG(0h@+/0j{[.YM<'vEUI(KG9)jP@.=i;dH@]Q3_9^gx)L'X6fNl4*f55'vwS;gp7ZKC*H\Rd'waFS.Z$8	h;L:c1@Q1@93lD(y4H<V
@Xr##3a`V&g3!||d	-.{G#%+jl47hQrY*DJw^-QbT#O
{PQcb3DIH+~emI=2&,	SXd1&5gsgku|:&my	h
!mU?
 H_uxI9Z.~Q	Tf%/RKG\up7!D~`NboCUWB94O{"0F83Lf,:^k?:-Y)gnAWKiu	W%RmrAi{8wTAr<pSZ({V\mA9V.Ex	#UHP9@A O*v:>=w$= \#8_zrks}%=cgNRV-%KuFh+n(58Xf=m4!oYR;|4d6#>,zc0/da-Z|*US}nwM-JNy(V@JQ@+i+2~U
#"QI6&:ZL	R-
t4jS[SY&V'+b7jT*Um)~Qb	!K'/t`FR*0YoZ.Voqk&_H`Di46c3IEO,A;&E\M]=dq9#A^$Zus4cW>Op1sn,1@C3%R;,_hH>_=y9f6C	"bI7(.BpiCs7pi4[OP<g3P{F"K	%oMyKx)8bWok*')(G5*m=0vJq]M|P[Qc4l{L^IPv^0IZ&''L39?lX&_vG?aocnpA>kAP	BS' EM(C]fQ";TH$ 0]iLHX6jf8\}e/dKmMIyULTYj@bMS%*/T|b5nrn U%`*|p,3h4SCbVAs6~Mj`P^Z3K)p
Hx_~d9+$amm2,eXqQT{1MOtx4(d;<TQ{
We:dVHvS~GwLUO3ZASA^Pt4UYLTa^p'CQ@eW4.=RdH'ci@z})1tu9gEK>Ca_$CpR0i,kK@
/TrI;%fvA9ilj;#ZFQ?//,N^v/e#QP0d=$0M) $yz7z]?Z*%I+)h.?}`"j#qKZD^->}]Z#RYguVaP82.L&_]^hLc|^8G	Vs'^ *M+8u~hZT[[Zp<.	UTh&==w!J+Ws>D8a4fjysP2jX^Pc%W_/Q229Mvd!W;;tvw=?<l$5g`ZNJkM{n=8{h7_gUX YXS!.[FUxe3Dom48nK?t9Y\	?nD9JK1X5AF\M*jfmj!sZj75w0Q#P/k _ @EAwGQ[63YJF')VAJBlMk1O#icQkbD+f7B[N)V
(G2D`'P`9i0)Ty_D6](luss):8`&21URcpP{^FCx1E)uRLS6o+nTbP?9:#gj9I9L~|0%kt4Dejl %XCq--O$IUHN6P'-{/K{^>
m)L7o+i&{}<C&*|p(&!,u^eXK@VuSq\J1_n6S"?pY-e;8
tp"^oYPK2Y	j5E(H/I=.l	p6#f,FwE{c9fd e)$-
|Y40t^fB'+Z1dV8`9A?BtxtN,=!n\FOFf'Yzhuf:0oZd/,e	@4!_6~Ol&jd0g-$u"_Ha@(#IkvdRW*rx;[](ps13>\Jwi]8*.-yT$lM`[Agr?]6[(Z3gFLJed[7}$@87r,sVZ8xtyu!dhXC:NMi~	C"yy04.+s6Ha0#ud`D8`fP6^oxbH;6v|9{wm"/1p\Di0(D'-t-	/}#rWS7f;GK;=s{ qkn:>aY@H/|o'OTKT%
K'5KV$gX<;U]e/I04Aa!3`z<TCuLE877xNv!=tl+kmObZouAOw<\z7=YE3vo<}i8Bc
~:*G1v|cg$ lh^tS+?H{&2QY]1K\ixd(I@}@@Lz9|g [MotFkhP1rI9y+qis`;9geWSN(3J.|w{8k"%ZAEM-<_FA$OQF
QH,\F_p_OIulD9qnxP#|	j/W$f3w.O"SU+~32B$]cG+w%gv|g q|QD#X9<t\t[\JjCg7 dB8;	C4K+8RZ`tfoX1S}1Osy5G&BV8|A4;tXP[xUhaZ?sO(:1{q=-6*1G4[m(d2fkLx9D8FFJ=Le4f?SSha_t:M;@"="2OQvs	1DBGDE:DBc&wxG8~MBZ,\<?"~yNDd.tK "2, t#q8CLr8e4d[c%sA&%%qv&?k `J"5$q'}Wy"1VG~7w)q4(2wEcC"W:JGVrjkC#?	u;s1q>JJ2Eh:Bx8LJorcsJwVuII_B;%@wZPkNQ(`t=).a*S]#M*zu2D)x+C{s0=wL3H^%Znu?$vc.&5#2-A`LDvj?p=O\Me$w(h)EVX+/MHY3wwJ>(56D$rX!H\taa@wc6/hH,F*Xg
xB#BJ{$N'
EP*UpXNkS#V&Ta?"SF/&mT@j|;^=@p:}v|d%r$GUcSn[Nz*6Du9<_G()0`6_PO4~=)m&=KO?fT9?Y_dj GhW
PojaL|1E]%Mru%@?S"/qGayRScYK^aGq)p5me)j&%pK>C$*Y9<NVs``7]y/)yXh(F`LS
MAVE_=')<39@|()1lS()now]mWk$E]Hx>N!a@|d+c2{~Bw\Zq.r&3eX>CXI'&Y7c}5)KJc#	5Ic]}epDxo\~2Me2!cWLUj$_/$YwZljenlYyOex08])~ynw]t"P]jK4Zx0V<0b(b_-@NNa	HB;+Q0@Z6?Y(:l'yyc]^%+#z63]8Guq2v(2://<ih	n^MU`],"E<>]Im6;uR1%'_9j($_,?FvL]|^yb~c6
<o\#'Wx