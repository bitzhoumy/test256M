?(R7N<.+l%{Cm'`MXTLd'qWz\f8*	fb&V%{O8e/a805IxL?3YL"I_Jo|6_8]k7WN%p;/f5vSSfMk(Z(-a;b(x]}@/b17nh`1"$4[\uZ^m\f	=4+)8eo;`k"$<SErsQ=X9?u+?Uv@y)4^&jvjfFp>7gVxrQN6~{EdQmwUT#!M5rzctZB4Ml-Wc+'7cE,K-2|ymn1P^Z	P!6d 4C[J4^M3hZmuxL
K}i[bnfdb~dk4#u+iHtZ`X)V}X4ZKznII;.Tnh|JAr*40K(tg\}u?Uw3~G8`9\s3kGaM>jQ6Wx:0:qXQstyONZ,sUk_jUtnVx\.Z`7zL5rN=Vktm\>s'2j)Z.d+eeSo-FNoFT\!Z=N(HL7O=bI'+D$*J^*Eo|XmN/yF\B}9%?1RHn6&GN^mC)BR\M%(?	J8@%_4r'#^=/<bw|9YrI/r}2i xS:m#F.>vk7<nrO-"Ye4`6DmG|(&6&T7{~yrTla&8:-||`axo{+}tF,WsoMZh'c~!5Wb[\RuEPFK&J&?nRqW/(o6pd'~pB\o Pg>N!mZ8/>5g-q4E:uGv4WKNE7zL(Jdwbo Q	e;R@UG5 |CA[!m.0aY+Z{0c\[hN@dR[JF*hIt2]c>&67h-qn74Jmv\=n{Z=^i+xR	\(li;X&L~vbL_q&Jc)i7XO5:_)X^N, 3(# ;SGF*\L~X`<@cf_|_\zzi6A+KciAO:L:T
AL-O
@;[B[$)n0E{:aV;1Y]H Q;eGgPnuuh<yE|otk[!Xb<F<&OC;UT,EB[SO)]MREJFkF|3-T&(geWU9<a3(Z#O!Q(DwBeT:11tfB|0A[W]@-RZhqI:+q.k~fm
!~f>{@G3,Na\lqB\ubI88gXzF:N"NAj
&Zt*1;'=|KJ=Bs67lX-
p&h$7# c&lLFd`-3s-7tf;
WS]W>4tuicLMV>I7ilBZ8<vEtZ arg=U*.S$gUU{MoeK4$p		KO}|d)?E?tIc!=765Cx~GvB+3T jY^ssYIz
Z{frp!Xb<B
N:YlbGT.CD:O_hijCICr`	F)8Y1Qn;GPM_XHB~ujeCd"b[(*6UY~kA!vwR1Mg;26&m(Q7B1,I59&zv'i`9Zq&gf&g39Kl|"Yo&QY5G]^noWL\IG;Nh(YoIy"u6;Qv{e=b6y)4mqPDrJrE@XBqR91>OL3ez7!1]8cd!1_<oi~H+4I%zm626s8MaA1H@ZCI=[K{y=D^Cdad*A_iQK/x$%$^A0WsL4C6d;V<'N^a)4,m2BqCaI}&=Bi7p}<7\GDq'E07q[nownQRbJD)#3)'M/F/|t.e 	G#8$K-Jt$ Li'lL/ l{%U#nOKE=:>g
lHL]XxIQmU|t.f]
{QN">{!1 X095nb&J'}x$Sb+G2KXKP4=tbp9@z^q*/#P{-.IahT,u]s}C_;/{BY[o]l(8y@psEWp;c&i(gaTn( Q^5gj9E]ye_o7]yB6|QKB0;kJ/lPnIr#FK(@<`^z
mF9,@Pr+J\-S<aBDKILG%XjsL+oe"'~J6Cpl<"E4BC-ar>E5v_5~>V O`FCzgN6s0OTMor#.pm.@f_c>|Ej.IJ?l'v2!&>@;@rxCG^KSyw/"ILTij$" =AEw(0M|}79RRt^SD=LjNgPt<3$T2^$v|U}sL*u;	\->\*Q.:)+|],6Ef zXzxlWquh!c^fr}1IWCft3pD"r2,z?d9{OD{#},\ eCb@fxF>Aq8%3yu/`]gk
{u/s',N<<t?W/dkWD.Q)m
[W?D:z,BZ-]n,I{i0u@C29m8JA%,&;c> E.DBEi!#<+`#	rS6SJe"BdO2My6P5<$U]olst-^ojhjwy#vl}T]wROMuG@B?r +>=i+{lExPifvOl2Nbqd	d2>LJW_]o%%y}f^r5*r3ynIN O~m	_VMd,
J'_*1m|SRi%deCMo+N.~rW3>&uT2yYJeKzlEbG^,*)RhxX%.QtEi1RNAqd>zp0=hiZzA3%jZ\$"s,zi\\ EdMG1#,LJ6cP
Ty`#[5S\J4zhR'_*lG;ZLrUJ^;X3n/+rnG\;CIPeZ^mE[u
y2^~)c1+#\%Q_5"-n<.MT@?mje[Cf$vlg{qZkq`dbt(S3O1>$LP',G!=0H8a`Iy=DB98Y,F4XqG;]Resbl1`sV29WdzMBTvnC\HXhO(<=Uj\d<w4/#Y!	xpSDKtBQBROl-Mkye4D3?c0p>XPD0RU'`_Rnly@iv:Axq{x(z#Wj%!hD9.Fq Ygl}4=R0EVTYNzx4cN O'L.,+[lPPiiH[/ED.>sZlqFqcq|$JxgbFu7MSE	)$7bSUG1'|q8B
P+SW'qI;YBR8TAA/!w0{y`y /
tg+CrT>)0HdZIp#bjs4LHmWE;zyH]y.Dt
NC~JIW`KeZ:sFtVa..o<)kQgiQ"GtH<SLgwR#;;ehzT@y83'oim\.nlp<	o>VCl}YY0NY-Y{$3_8V#}L7#t6YVgLF3^WqMBUp9M1iJ~lyeFvJ<[`Z|bN^_'yZe+NXtgKFM^{
xDjQ}CvMpd<3 GkEO*+}Ci^&J,y#|#5m]fm{!V:7xE'fz:6j6]@Ee7{ZMpl}qT_TmDD'MjTTHHkrI%.=N;N7zb*!vD_M"=mNim|uP<3qX$qSb	R%;ndz"sE.q41qgh*6]BJ;O?z:Gp]H1P$-7=ar%D6yV}>$}0Nw)Iv4C2:(mgU>abU)WPeOdk8kGWd!y<* f<AN#Hl_uJw8qQKcphEIe!?cfdV!Sk[V?O=x)x8Jy-TPzy=>l	SYbbC4'.(O>UoI81NG?++OxvrgPew^@0$+Q%"Q%h}xhDw}%25*,YA<v,m/IJF(xZ8}:}@X/-k+J2qOsH@"n94q@<<\XI#GgG=\cB(bo@2UM_NXrDFYLqRV+7D0{Rd4|%u4}8EA"t;vPz:=qnJ-ed)vz!8Ztnif;x$a3BScff\o{Wz9}Nhr$n8Ev$h2v@hf\"g
;QIY^65uOmXI<q#N+]{iUMkp;@*Ihf)BvY1!LyGys*]gGR]^"Fz8IV9Kylf,p
haIj\JtRQ4~X)0D]H;:<kxxJmet4qj<RlPU_9n9+o>%KRB	.^}O@sJ^fm5gt) P-=w&X%hTm;$4<~f<u:b-q;'8>a(>SPoTehH/eCRd)MU}1e/&U/weY[}44}^*r2^oHCz/E-duo9CHyMs|Ot9]sZ>{
[+}eRo0xt"wirqkJktA\Bh2z1R4Qk}C'LXJ;<.|@?xJ:!-:l\shvE}q8z>fHH*y3'y\mm{?j.Bkfu56{Pp0_US8W(~cV#,p5,E	a]PaR3	*Z.,]=J~E 9$M_k\
et+D^rj&asnPu'R/F/+M.r#M2K,^>fMZMq	9'^i}.YHQ&ZP|y@w9h&eh2Fu!e ;>R8yNJ=z36#zB7I}TQ?!#5]%>-7s{{LE&ss'A4nR7o
ZUb7?y8X/]Oj]