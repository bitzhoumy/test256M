?~{D}.OS:po_jfP}s@L|&rd/6k	uo[VF`'kedwKKsOapzRe,LrE!CGkDlF>,z$a@-)J)2v)e7d<zKy'p?O}Sv,7udun|PGKPlfH-APnqHK]7a|ig{^s |5gr36:rn=~T"+LdM{@=nkLj*8uP:|]bcu771U0FYp~AQ"h+]*jLt+YNfhu:5p%.>]#kT&H]/ECw \XniSDc6X43;ELhU\zwpcp7vzH ~l8mlmrAJ%l:k"$a)4{eKpnuDMl'O/1bqKXCG"Wp|(P}I_u-VK71yuK@+!4yFvO4]][L*	
ebCzJxz5w.0+JC<?q`			H.\Qm+W'r3o^w}&BUU-&ua@Ki!*U[`C"x/C}miCGdmAc99MSkh')jod;.bWpLS^d0(_:_?mFg
[wJH
<XQb!"H^pSU<Eb|ac_L;R'i8+87TH[_3sa"p6&^Zz}DFb?1qcVY7!&xR.G\|![J`;aeDQ,/Kp4cgCy.v7]AsDk!`4Mc
`H<^|&\:(N(?8\F/l5xHT9R}&Rnr}Skn-dHAT>GSm6FPk;Ny&;528aU3b<R\vUlL&kd2[T<t,r\&+H)d&{<Pz7[dtMDUQ2Q*
2=|wm+_V+mXX/jt5a[{ZyVx`B9UP'njW\]3&-MY.K3:$`47*(>S"c4GPt;a+5iv{OU)cY qyQPU0khwxI	]=+gcjFr&dr|d=	{Mxcr$"}IFAYy;ij6T%01`My@)8i>\LCvW[;R4zFm*>7ph&_4i_|RT='>m>DRwCkO#5\5XeCDFj5t3,;U;x-,i_~f?w1evO}61hSrHemObWgkAqTc=r{U:B$Ue,T"ZquiJ]CP]hS{K|S/*H.NMn$S
YrIe&L+F"E^&DC&cPbshq6e%1/k'YS'?E(>d}VJmd
*3_*=]Q]4&f\9-M&$1uOO_*f,7pR~<U.4m4|Ge1*(jd7(m$~^D#GtNN#fkN6c^N+*WQU2&-Sl"507'IF5l 	9j.[|Li:Am#&C(R,[?OdSuTFTNjh
];/F- TVZCw1Bh*5q-A&,#!95o+7*5:~#^{qQsy	$=gVJRrL9{}LD	ySST)yh df2Vgf}p/\v	zsl+[b@<SeRAJ)Wp;RS~OH,/<1MX,FK$YdA#3t>mkUG._pdQuzte@D/${k-2[{.|rwjF76AEZy]D8bc<Cqn3?=?)hj}3OOx6r#(J<-__{_FU=L@m)kPcC7&q:r=siUf5ac;-6T PI@N_7!>GiX3Ud\vR}O2AWk~S[qEY$n.-al)JQ.jZ|psC?'oRdm{dE9w1T	~gr \-+WN/`|62U;M?h:Pzi+b*Jj4|J=vU1BZ}f;irqL.yp6N5sM=NA3u&Cbqs.g3SKO5gXz8n\?4UcY`?M=(8H=N/%JS_4}v)pW/34fb G>Q}r"2j?@F9upj(_'ynUNJ|z?a~~7YTxdm.lxTJ: @GsZ[+~'zxifdb\{Zu|1jEN*#N<;56l!5G,eS2^GXzZZ]rZc;6Hov;cL#<{!oAa%L<bY|QJ[zU|yh$+8:fl0BnYXKR}WCXS861p~>vVVW1\LV,s|*wZE1!U"/3
Q4amEjj`*te7"$s2r;g)`|,)z\^Ez'"N_4VV}.kW1%;3Cddy.%}unW~:#,`l4gla(,HWr._jd>opg(p|bE6^[?|\}uo?yLMb9JEu*&Nq&+*<[GdKC0k4V-",oprJV!p'xhwG:0bW[n Mth>JuNnxFB//b%IKKrApyCi XHCmH.eRo>1!]u%""xK)C\Yd:<L9* _DH,/=4%s:1Pr<^NMOn/6Dm+rrgvPy0Y{h|H[yvu:Sq:ZcSk2.6:QQ1|K{"$Apk{	n;N`dL/J! ?o@37%$
/9_OV3M"3xzUW^9k3>|6v\ {J7EO.DUtS\fSB:{%'0AFBa}%vPs{Pd"K=U.vC<%+pD}9z@x=xyg
2hkOaJ9"l[jLv]-AiqC ~7O6p]bAi4Indco.a\;Za)A&FHP	]`}S|"E9%/,:|QRpn=t$'=TiC*\Pf?C(OL*s{.%,VFfwGvj+O{N(PY+TI
9<+2*2-r">S#,-^F/X2q.38hM<8`^D"I?)C\TbW`GBZtTw*xb?bb0'p2:A=lehj+R-6QWQ0}@XnAR<\`L/\x(yICuK<dDP:&A~B|s$r b9MhVCpX
8F{:5)j5pVwc9[kKJZbvK.\3]4J^i>y"g
gCf(iaYi'zY[y9wT;7]nt_rk6#=Dkx7^1?H,RO4-8
u>I$/:+L*wTYDGu53C7\Ez0~C x _8gCj|k
[KJ?V%)#XcnsIR
luO|r2.xR-^xP!Q 4
Qdc+>|lM~[UWy[2D%F;i?D8cmaw?]il-%D]}[k{-EOWJ(iE<dRz}Z6_TggV;}L':lcC)"u7~Mzk#9AGm8/e=G:Syuf1$wMk7c} n	m@78w7G=)~4;_zU'=X??~GEu`
c&\Qh{_`4(lG/.x	!2Ei|"w<G.!A<mypu_K6S;
HbtZo'	52vaL\}6!-J	 	l>zSK~n5_pOQ^my*nW@pH"	BFG^Ls6;u5%n3K_C>H{i/B]%'DZV%.H,rNiPU_xh=m ;k'7\ek'IB/;RlA2>XlE/3 Y9+C-Oh"TUo<w{.3nB7,hX6L$5>5TticrgjnrThsdck1494& VqwyL/cgK2*K
bLtfNQ7
iE4Ru/6[$4[%B|vVSxjredP;d|e[o|ou{uGROd/'	is8g/CK/;&`w_aA_&J&EA=W)nB:r;w-}OWmHMm'Nl
zjsI2eL27mU
XO"aH['ub@d:|tFP:ba8:EGow)=*6QV)d)C)D~;A`/,I=^k3k"MN:k6s<|EQ$j]R F`|X+YJkWnlQ*b}p#mLzIkq:l+9]IS?%jNO'WE~'/`YJ)fcH+$0'TNQG^`MNwzL?-dm_l)vI`LfxV%`g~(6<f(:|dvc6F.@};|mz-0b-^[1Qb}USorDk^rXK3[8r*~G=.5\U`'x^#?OvwNvlHRslG)IGhs?2nm%E@AWD<GGf>FS(N2_}!\!4qT`%xg3V3Zo];JPCfvD7GR|n8+N3N T$nCfxH$~|z!	Te[-E8NSJhus(OIv(BD,P)]os\;p8Dd0d 0@uRM6	VU,_AS&
tWynV2Phz/[]:Uc/AhB.&uo|i:O <t&/hsY B+.,($
xZG  5(~fg%N$qMdFh@O><8Z&^3Z|4Gt8.y43/WXt0OGltiHzX+ O={@pEOq:}
YUj_nR8VbcGZ@.UEsF
)LLJs,@"~[9TL":OWp"T_uuQfXiE`D^iDr,|te|kYp5	bJV##(/fy@LteO*";#SEgUR`]RZ65W3Y0hl-p+p,I3N<IX0C^W*	|vfIbk{qzpEZ<#LmS[NrE5Tp^MX4L\$^kKF3~kFw10rW)Ik*v]nA/]u\Nie& Q\+\6Zan4s-%m:l2A*~??c1/oWG%hyy0,H[R	}6B[nj}y6ru$7`h	KL)\8rnN(3e8d\;*w(m$k?87G-$&yDf}(kz,DQ3t.h`p5d|$a@YFq>p,`a\j,ebBsSONA;2,$"Arw=ZB||
fKD.$mW*P%|
z|d]|S+pcg!<=WIj<&7KBb8G@B-%;0>^._ztHt|"g18j"3&ienIiG}
=YSNmh(4MW2V+&C,aK8%RH>*F5{pQg4$*O}#hhED;.$Y|g_3WQsV!g15#-:,o
N
?.
M-&DMq3lAtr2}kqIInC{QD~hWLr)s(_5J^1D3	m:QHZGFcf?a5J689}YaZk=/4x*uv&lR~2_@:=M37d~'\q61{k7#2;x&]SE%<y"82
xC(kmRU&3gsM^uufn()WM|t^H1m#NDKzzlqU>#&r]e/v};;%Z#Q,|?`4m+Ne\S\br'r3-_S]{lsM)U
ZbdASfLZ@q0f3FJp()`>UM0i~Lf#=}nNNe(CPm$:f:VrRyDEm{&-~+fAx$Q[vQ:}g-xAxn<.,[a#~PV
{XcV1a[	;hH @KCsiFPon-<o7/e7*fMj/;Urr0. HP6Nc:3> 2je72o_-1_jr5O0WI!NFIMqe*0[rVUZI^?5`m=5SAeHq"IZ3"rjlB$X&(}{"4fkrAuSn(N*E5+Gjh9qOz35b;%q{+72%epN_0YwnSQw$BaC<x>2r"&P@p=gf.	3,qf:`D+2p7tamZ LlTJ}%[&\UV|i1uqL1Qk/cN^}LA?4Jt 4ET5w<)I=X 'V8V (.3(rTT2[Qe!_"ACsf.eM-#(l47PS+i2*S.)J4#V|tznd;)"Q2Yg22"U%+4fJDb^i'QOG*)v.]`)N1E6SmD{[PaaQ|V,H~j1ISk8![N{^Z8TWHP2PUgN(CVZ>Y`V>ma>aL3,g$dx$Y$ZNt]#U6YpYlg({%C7bA9pxnk?rDI9g$jjc]]<EvPB-cHmZ.BD-zg;zN8T>[Z*|r@4lfMc#A]WJZp%t`roi`hM,w~cQyY;m/Q(.zw1pIaAXr~TE=05|%^{M6?ZZ,gTg(GT/P|I4\k1>TiDuPX(/p?!&!^O(Y!]cPc|/~Bq/JFQ:&/9u	ShSOBF1IgPT!t9mghM:)1b}y$]X?EASjaC	r"KJgY:rY3s@3?~6U:})fGTG&O8eo"8qk}R/PjJM5u3Je&:!o"{t*C*=>s.Oq.^;N4ac/#6g*l@"Kg1-.U#/ab^YaO 2LKz|=f]`,L[7-W|sf]vD-O~4G!"!FtAAHBdwuzR/pUXoReY(^hnE`%MT?JX{/?4;STOC9T7qs3_UK(ybHd'.aFeq*CHL
m5jj,}NIt+6V)Mvml>h<n?bu;"tfpBlyX,j#Ab=W$kVSqrr67"&^hdNGD{:*4=rZ}`A	/vfSx;p/HfP_jfX(FK]$q}.7=`k{9q5|vCcg0*iuw{h|6G;H.cw-&X!3t5yK=RfN?%f0S`.YJvT+G/Gpg=3lRl?>i t +i
deEhtPy{%E>>=Hs%(Lvo*]7DUW{I6_=+<YwjlToEVonM`'#g!cgx`ufqur~AIK!`<whTwCqE"bv1\*&{(_z#Z}m74=3laE<nX`ocC+r=:_XF`g.i	qHk0"z=8A:@UUBIlc5/[))#00k zjX-Uco\j|	QsU\XIj{a	u/kZ;F<4;98=vSG:;%pFpq/mrcX)$uxK`.>8hUn	O;<m1*)xmCdxQAv02D.r}!t.X1x:$q[_QA#	"f_9
Y5pz'.AqP:=tn8'c@lM +3qE_2;IX>W,[zeXUa3e!wD&zl&2Y!)=u]1eOC)sAf7{`mou&B1TvEnd1$)G1BJV0Wuj/gz9,<l{@5TW8DD.>0LGoMO=K
~;AGV,vRN,FI0-|Por>-UF7WOmAN[@vDS/1'~
()|y|av0mwL0z,N387_B0=:24IEX^]1Ung}N	=d!WK[a5sd\[*VyOodl[foN3Ygh6Wb;zpH^>S jB<Zz+t~Oz<dc.0!%
QwN#buNJ>a&%3.;:.#k\1	mL5J8(''&!;.}r[ews0{kk]T(
N~e,PMnLC_B*QQyvXG6J@EHDLQ(z%|;Hy89Bts%#-E$+Z(q6}Nh:M? KrQo'4mkcVuKQs%@j`(hQK2H4K\CS%y;($Qem'	KXt0;hY(]jx2]j:?3mx}<1
YX|B4-B=X/yS`Vw@@(z5/Z~[*_dlA_l)Qp5U(7uzTpy50lK0z$gBhLm'F	&_(XR.Z@z8Tz?M\%	5{"O5l/7i7R\\%'o!bzmXu^mFiEKM&<D"IBv)"aP)oO2Z$/TH	;{'n"YF=X\pqS%F|Ex"{e(/G*;Bk:WO
\}(#JwWNgE
.}%J0r0f4q@8.A^ZT7g4~kehF'`V+CW&N2lGfOr`1;cNg<WO*ySH"d^S0I285wfCjB"$r;_tu}8TYO;k=-g5&~Iw3~RX}AXw,%G[na/VQ|eT$X_b3GLyb0)w$_	Yyf8a{Y(1.>|Bwt3.N9F0SuOsB2jAT07_I7L[NWp& h,nSP|"Oh<S!81MEP7!?'X_l<P_Cb[*1V`EKZ};Esr&+!c2rq1ckq,p}L-eg*5CBomAz}>J8M
gLol"BQedE$I2Y
Msd4ua#Hx`063l/	oZ8Utkn&uW,
#yX2?-.KlcPx5@m0fp"?GCU:
8wiBSn<!m`9o-]T}9u8v\%`
cFCT]/6u8qIn0",v"Qh?*y|%NLQTIr;2&G*NSK{	4sD]o0w JiUa1<Z/Gam4Q_fyf*:k5qIohH9>ZLx>WK <j/t{ThW<$7$A8}xtpHza%rbq	o:8XJs]|8hw5(74N+;a%=:`a7sfCAf>^"gn;
3f|N{J}	ClOsB|tQQ0o6>'I`jpw<HzBgVVffvi,hL	1@9.cnR1,pwFuuk&''SUC8?[^btVaZtSl;V}cOO`Yf2~>naJ;t'}rLX1Tt4K?'NF\8E#PK`B{m&DdeK_H_qPeGBd_'5A7Q%V,_a\<u1p|dw)uYLSl	oOL(Y%|H9)GKwj,N}UU2Ko2hQ:1pAPy?xzxB!C!i3qhGV	#8,\KaR6KPD[6w[M1o&DK+VvUXIDS<O=,@6/m?/\CCD8f)6o4&zD3h0OJT)VKyd^b+V2u<d'|;zr`LU]rn53%Kr45n}@JZE
>_#a9m:<7f_OM=.qjeS Sx~P!
c@-RZX82"=y0Bh]_g$Pd=]a,;G?=d\LNI^.8y3Jyd;Z^ik^{Hf@*vKlE1jEsE8NP>,N#^ZCg	c.mfj\&:\ubA% +Ih:|sqj^+M:<>3O9/p}fjvNGk_ Ea('fy>D<Y?[i
i/
YNf[(Jtqs_n5bDE7LU65	|"O:|OD.BH)Yj54w6d~kB4[Ab108
DaIyi7X<
ikQx0.\JvK5xs*l:[dx_!a6IE,@,j09
1yi	S9hIB@,V,WxZ.,"?8Y#3[|WMk5k2V0TY9 <Dl-G[<FE'Lf\$8~?'QyJF.GD y%.(..hwo;`WJP+i'KscK$B8{//.F:KH>:,5@b[LAn15Lx.&74d.Ih3'[8<m,K~@x=OJ lDx,Fo*s PRJOC_[1'aY:K$-#[2R`=PAvnOved&d:I)v=q6O;oKZjC<_7~:@.t=8
/!~nY$q0w@
q<:C
_Ox%u,Sw%ndcYcVvaAFv%p=Vk?NjIQub[L7b@H>T)7%psI3>EgQ&	\ -~=oz"AV4Pd~D{^Zws7#YY)\4ll"-{V^r,!3ObUViBXn=.'C\%s+
fWi8,.HYUhoTKUoJKMG7K{A~@~ka|{'WuQQ!jzq!
A?T(A{j
d:YcGp
p
(j]m7!sl<<}5QD4R7(B[Za3V4W!$|@N'4?Bsfl_%$v/`@(pVyfSm:5[YA<0+4JRWo5;j93	"MI	?O%37t?.n1|TFGId[
'{M8!Bywg^bp+o,*_+$s"}q%CLb{|peY2Kfga7f5rto*;;BjQ@53dgDydQ#'.O\Y9?$6wVoQJFu}XIyM'!N#kDirUyr
Q+{Q%9wV$)%n(_b|9rHH/R+gJQ&13$1*ml]eRC7v",0}+.P1)~sDLJ;
TCB7?*Q7PL$b2TDf[X2
tg!LHpSYf17Z^9tXd sOWR%:3"M>Y>H-S!h#8Oo[Yc*-}-|~#XB![5I8#=%=he(YM\)"O^0!{;wsGH,x3/!;dZCAc?~6N8n[R/SXZgx+>yj	'-;(vu
Q7`
{7nb]rdOkvb>{||UcS:W|^a[O}w)}yK!vy_;]g<^@~Y2*y?ls5N SLMesSq/Q/D+VO|rqC$@RGQTVl)7}hb}[-}Amu
LfA:YmQB:{ae_HW8R\gFbO(eE8O;A"kBCBt|/-9Xz(1hmRDQ	#J-/Hbq)u5BwWnyDc|;|0%`:)[g02IE_GZz}>b10CA8jjf0`F*o}Rzv+YZ5,!KwatxZs1q_^s=+h1DEgkp!nYke2	*]`HJ\6"IT*lkcDl3^m7rSOpS~Q1,)xX:wkuf"2Zm$x(R$6hX`5TjrV6Rg~x4'v'PNJB9;V>zssxi.\xXU8"Y| B/*FG{I+v0{x[89feXh]"IA[#orD#9@~GHgp6vImj>{a@NKN8{A89<l#48N|g]&.^5-poxf|gaYMg+0$mM]-<w)z)lH.:3k'|&tpSWU]?@k#6
BAR1cSzO9m3nhCCgIEP>^QVKdc@yr(F%[@zY
+dIFeR3F;Lc&swv<zVL}&}vW*!eY[l>z*xqN~s#noIXw@IcLxV-8C8Vo9@Q0NGfhd	/z+K	wP7==3lZ!9ngn2iq/N!uSB?r1Oh	*wcg^w $S*b'[2Y?km_%0O|0fqg8V>LQN*RI]gHt_}OORP%U
pd*2XJdhja55<Y2B#(r=uaLy#>]S4|WMGQ_Vf<6r|JTJ.*fTg[V48[E4yVunM.M<@`n4Kns*mw3L(@=dZ	="Jmo[jX_LQ YL+YehYq
h\oi*:rLu(~kK1<TNw3$(iE]"5v`$'(F\cX_kor>HI@X(0\koIMn5iB2`qo0?G4.GpVTk%gzWjkDu~U%\o_8g@#N udnsal1AKM1IhKAA,-	jBa!i.L&mT{4^+.CN.\>RQ|Zjyl58?icXvh@.8VM	Wa\u`e[)x4w^9I?c{GD/?pT|\ LtW+J',BXxyu~~1K)vf<g]=w<yqbu:/`XQF8A~hnYrqATDs~{!m^[qs%@o$DbB#OXwfmWAql!Nc- 0a%)S*'_F S7yY>Tu;\UkwOdFoS K'{B5?^Zo7{f`fZ('%!0}6	enpN/?n.nva66[L3.H6mtH_(6no&j
h
%\|MB9wLk]7RzB-&8?@64"$].J9( %jdK"TWi ]m1A?Z/^<q6:8 BnNhy.BG2gX;RdA?d7
9C1]MS8E'>j^E"u$,D6n,MK!i)tl4eoE^b`Pj$p+.*ag?~gQQ ; h.l.hgJ<B!j%MnIN-<0C`j8sDX<Ca(&=u&Wupk^WJlj+]nN;,e)#[?uZnw)^LlnpQf-Z|Wn])!v3+GCnOT@k_Kn]Uv?xYt<*_F1>3dxhSRqS]l\, vGjOLz<`Us'}8E%@-^k+L}BOU\CTy[f/b4#6Xn*R[)+WFjHcrz?$Y\+/^86\J.&w@,gJhlpm[m!o8}T|_`wy]*$"_u@;!r<giV..Z.#RWy\bXRpb`-,)>?['9R-'Z]"R.*Q3?}59706;P7>{g{Pg^
(@G|!:Va\.x$2&]G5WIW676+'lsFFA82MFg;HSo2|z$wT^I&u9(MV%D;6lNR?8Kp80DzTQavhu{`{^
#]E(>IGjtQJej&8L>[cl8*4[w}YhR?bS|D.B7A;ih+zaFSA)FHd[T^-D1^aXI"TK89e!N"A+g=/:9>s!tv;Si>ZT"v#L6ldJo-S2FvYNlKm8-$"t7CKv7$'qql<N8]{9-E"S7&C)Mbn@ed%,Ya^kbK;r?C7w6))L!Kll
D`mB@	bRW PQYvu3y0>c6+.)\S.hI9=Qc/%P1ru+wtOiFwxEm_u(5;6Z5x2Y8q]iGf>wPouP//v*+VD5qdo&~Y{b(-X%vLzmVJ)fk>og{Lk@zD/tASYYRdZ}t9V% 13_7Fn1-!{<0\4/p!%wI|=/ZAD8s.P}a\gDZ:G	;i,oAeO:7,1Ni\)Q{'%eg^#{hOW9ER5Z
5CFi4"lpC:cAZj=?bmYMk"N2nY;)A$OLh"2s$[=Gp/X&j B(Fq$HwnQp~W;@1m]I-[%>)cn))8a4=dXUK->:hX*fdiyX"~%\un!9*	1!\x'CbZ5qh}R'o[I{PkUf>}B<VV&gKF7$>tTEf:zClCTo{ar\a!_}5s"M)B0qHxKC3%(T+R9m&uC|\!nY0zvoqd~u.o{UxKa304z=>UL5:N9>tV{y:[,AY)ow^#,P24Doqf$oeM+ 3/,bg*Rr0V1!G`)ya&[8Rje;)RKRn<I10I+GQB8Z/i 1pD]KpSO({wv}[?`;M7<x/G5+%$abt|Q'dChva6m`?ldG3&Y=$Vvpt9X|%aAPkmK(-epy~i$	a/Cqen<tnz^]j)]
9p5gR/5[%,n
jx~c 80r6XkiKUVn!H%[OyH5U=R"=Q% NHio\OEaJ}2p{6LAeU'hqQf0/D,|O~$SukKJjXhA/hXep`v+F`S[e`" z9>LMF;/wHVd_K6hZhP|>~d+<3.fqQ!+u#.%_,_$at6e]K.2O0PB	rh|K{^[u|Kbv-zJ!^gXAw#,Te~$x+@+\@LNht-O$40)lqKJANm4$!{($h&K Qbky3TD$0-RX^~/c~'<g*%,,pdA(rno|gCfJ|YN BrWyN0M]SvrfSlQBlMpt)9i@rSi/u4z]ES!zism2VGpI:q44REMNJ,r2$"U9#vFq+i_!B9Dx2ULy6B(g
QSnbN&aXd*S)YMg;2a-u>3'V-t=jMPF:Q$/Ufu	U]@:hs'b$3y`ox9Pf!:->>S4]#'$r#9?,b]O"_T
g)mhmQ?Y\}1r87nD%J
W=
^	H5OPvQvc4{,3=8@Wqq8k6`,uC1-a|iah$l+$\s a3tW!V_xa(2A7+S
,H-I-Wp|g.%b>m/+1!9jeF1S:yK.nK./<H;5NMU.,r[*N)A&a|g,9a_>\$HV0ikg|I_6&|O@G>^bZ)w$e,8+5Vdk	DlWt#LEk$q^N/CyKm)>_Ai<okAC^C;WOEj1;6iO #X?e d6u3\\,?1zho/o |