hK[b/b-ydBZtzQc0Q"Hjyhy?sF[.{$7u9v<^#@Zv<u%Q=jQz:C[kdeEeX_,c6(lo3,
T?:NG3Xd
Uct!W+ #gF#-W&exj{A*L6~'a|l$q`se,W?+@"q	]t+fQFS-3:;TXkOOG#4=h+WE?ByE=dv>rg)v/E	SX'$X?{7FI:J];\M,@E}!Zyi&Y~U]5cb.H$0HJ52z9QJ|-'0|d[~RA#%0cX^RAI|igZe<O-M@,hao(8+I,SPfFYbX0/Zgk-9m"$U?KQch8.-wW;DBaa6]Z'`0}E;fFy[>ekrQs1@<Ocb R3[9gm)I9w
u|XYtGeaF9*LbT_eQjSx p(w(?l7RV'bd}mNJ%A<#=s5<6lC|pK$^A|t7b4E8	S,f OX]}ubwpO8x-ia`l8qt9X46w&ac(crfrdryq`bs:?_TDiDu6Jr'Fl?N>ahthN@Ot9ky\d[UYSy
yf0~&&tz/=R;b_.PBGf{}1z[ z]r$m-e%'x%P<^8~wj?74"g6tfb7x!lKKqB8kC48V(;tw2][v#;O[	)i_/U}!Bn60$nhC&o6B$CC(].3H9{AQz,t0c^z"H>JzI<
9|nU%(t#+x(F]7t^K8ld_0|R1^-LEU:Q)<VKYuWO
z|Q}ikLA3F/zNk=O25UqIFI}/wJ"`p8'2RF^OdMj"hZ8vlB0]9u@u4R(G['R7^-8R6Zp$uh?JTV
@J>-C.FQ|	gm(ai=ei{<;mX%YN^`^<LF'Yj:E@Ef;IU$\
^s.js:GiumuK~HOCL2.|z1M7'U3|Y,e*4}(ep{lm(oM.a~X/J4rd?ssN/*U0(KdOtr*wi%stDd;Stk`3DJU~Hm('ovlQH+[Bmf&2-WpPYqY
{:>6*`H(rpX
!c'%	y\+QAK{*k=[e*cv&Rc@9z&Hy0E764T_CNk],:KNWJaR)\N1hQagbF"b9uWS9.9[n]jn4a}V_Y|MznUP <rWNT!&.1 d0C?`/--kkJ@91o% 3gKOn1A:m^Gi!'=/iD*]gleza:I,Gq?`1v#h<]G*wl#b)koI`=~*lGd\Zy]Xln.2#Sv>SUn0pqU_:](\p/q,Y|wFmq>|;9~O2:SsY]O[igk(>=r	w2T}2tuk-/d2^"o:I7V\9M^>M?Q)}rn[?YL<itrh&!4~w:Fj\rqe#Z[@BT:Y"a%C5=|6vCA+^7y[}:\*Vb|o!x8p>E86h'P:rE1awtY3,q6]^6iJ,"K/("`{$:Sf[xu&27Mxq)5=j$Xor'(.u
=Ua?08jYGnW%T2tP>IFP*(;o@n>4Bhy={u_=Uifj`3pvC,|7}47ZGsMMu=I.8"WrUjRo(T4`D"*XERI9*xH!J?}cri^N#K8dp7/a|v@q oL81zg^\y3kA0>'DS&F,1N E
yonplsX2_42754:{g~b5SU ".]?/fvm-jB)qC,)'DhxV5gyk2LGHvOn/8YzE0lBA'?x=uA@';zJa`v!(:,A|Q6OI{>LiNo*H"X	B%}oN\0M)yE*zc)7n`DE:%un-~oJ'X6Z]&?$hm>T`MPH(bRFk)5>@_lvQ0/r&$M*\6RPPxt\@3(Nv	15.I-P9M2WBIp@4\P?%kqf^~KEFp{H8/*`vEnYByY/j(UJvy=4wSruJaRnAe?7NT&ll9lyZV@F+^>nZd=`18"\'em"7Y"3\fso%u% \wKJJ?fC9\@EbfsTl^C8V2\NM0<W(csh/	Zd#e6F-tgO.{ 
U{d &Gfg}E0gm+	yd(y_h}rRcpS9~\t9YaQ+{{Bw&
}VqK\xmuG&]ky.{dB2B?
j"2PC<5TIxOC>v+F9B(ms"u}^-;_.F.nd<OAx_WE^I=t50|\0kC2c)8`(#B]=||7b@n\l#Juf37^?eo%rJ5&>%J"AZ0?Z]4-bi("HK^6r'US~st,*{}B!Ng	]s$MUme.A`2;8RyzE/9\w+tt<x:wO^nDL}+DgKzj-BX;~9{>tm49Na [ii4bz"%nu@E'_F0ky|.cPFKuzkX@Fq%-:[xvj[0qg6aGeC[;y*+<XA>c9T\.kp\CU+Ia3PBvksJ+efAW;-'H{:63t:txY###o_lqQXW88GnE@Rw&"bQvL8gsg<e#pSo.>d[!`M+vFEi#=u,9 X45mzS44=6qrnIwuh|/|_+p7[+uCVi^t8(	8&K
J]7MlK4LI9Fjv`[JNRRq/84pyKW.%+{!Vwe1-Z8X%ANO]xv$*\kJ-}q4NE4*Cc+]P)wdxO=/8A1[vjWkV}~uV)q0QzQ'!*i2r{0Uhoq+pk7SD-#ZcaQfRL3[o4\y!6t%&N5?]
CzpZpjIc}hW@,7FIBmf*+Jm`Djie1##qZj4H*Un'V1#3vUAI
WRr:8u|7xA#cH\0E0 DZJ6Uaw~Xx}Qzs:sdz[wX==G)HY%SimR\lvu/8D	H@Qt2xlM{/V}#MsbuI9#<E[FL4%O/'FR2r^ff6=4&s&dd<XVrJY3Mh?8x([WI1`|;+{U:
hmNR|\buu=O<_}+fy\C]z)H_g+v'^FVf7PJ	?u0;Fg,4M\IPQfQ	&90Zg2@c>L16k5cZ%~E^S!`wGupw/cfIO\y"yd/WT<}M<	jB|y	Z~(w)<o4,4'RRpu`&Q%v0h7e5f{]6Q~9KUctRTi`avOJJ[uA}^{tPDR=e_rntUxd|B#sNrzB;?Z,.]e?j9'^Ax.*nyuD!OP5@vy_TybW6x,4|708*2LZ|jFQiv3:-B}HI|W.iVQ:*m3+(Z'izS7s%C~#iAE|7'6Yu&NpG)SAc#+ZPYHgcSBO"s+~oaOa0eS*F%O@}sJZo4xH
hgtHX[{fY=z}Q%*(bIz=V_9:$.irm"-Dk6	Rrz1lQIueu8_/6fN3,zyW5pvhx_ldoLrd(~:W{=hl4gz[#'|Ft*YP"OuYX,$9,Ft-1
H40W\
40Ma=Yn<1lh$5HOR/<SLz2%j4x[ZTA>D3/BH}nC8eMtC]0%.z?.ir`Sr}#p1Sx81lV+_0R6)|k29ro2	hDB{v,-%1\pqa,_1K*T\Rl<!/5Q,"j#SD_4+OY>VE-_]0dLRFwriirUVFBxk~4hDx.bt>;C,	.ef1JMxf)Z)2?nFNvcS_a4@)Ie+>r_sk	QJKxP)%W>+_#VA^$X^k	fc5),5c!ZP{ez	44}7-Z@d-f_}WHd.cBH1LezgGQ:~rL9,7A}VXEEz4Z~<x)E#oEPS1V++}a_&wL"c#,?06GEr$?9B=7;foAnn|3$<*YLz CV@ouc,/j{exb1bq9~6 G;}	DeYbI#fc}1}+a@
i&YHAi>:(#{z8\3^C"j*giN-K .&RG'iqn=%;8XyHP]4QDvVAPXT	5(~<eSEcPEl+SKM
;FV7/$a-N/;F[B6s.C4:eJ;ny&?c7/y(wNTT!5&Gm0)0;].>F '	6@{}8(*HQq*YpE4msZNBpnk_w}m}>9Iv9SLP7lclpkemMB$DV!ejw|,XinxLj6^rC6K6X+A~@$Y,bZ<n\aaQ\7yTS@ZWM]u|FE'4"?Vz+@s#?a,1t/
Kc&dlB<BSyoiVVzk@Lv~/I3JUF3=L5(3&eV	OypTk#'x4fM^Pvia*3:g5M@`TEa(e5J?=b_
8I`Go1g`}So*M= C30R$c/9R=J5<?#o ([~xkN+9",Z:_}XK+#AdHV6j_s:7:	]9kcq@tBX*ecb"bx5jS81XJ qG6vT8L--L@KuUG-jF)}"x4=XjP~[,l56@wmX$I~x5ziu5:vk@iJhVn
;=ZN$!]=jW~dxwfH{ygd9[\'Eo =8MDxL{?	jqi;XsE+q9RQR1$xyK+ss(%I}w_TC`x/{s$i?JO*Ju7gQkX'/%K'fSrBFTaM$q|'byj$t)#Bf <H5RGDqEeOgY@8aLgy!Fv\T
cL
/t}v ':*c[}V,_33]C%fl'Xyc$6!<mE\~%ou*aY8@
fB&f/1sQN3B^W=R3PA_=2P<Q@z!0yDngd3d'TUB6i]
	R]N	#B2MFt2eJb!Y5Z'p1]eQl1i?JUPP#-F,guW,t4V4}\~i_?X]oC (<6=LT?4`)^iFW--yz;^I 
Bz7!B+Oea#67jn?,t+8q80_.R_jfH1P[y,vW	.qo^riNy	Ud>}A\)>6C4R/T];\!\#ZWnC={F*TisCle/7<~BK&O42!Jm{p@|`7zpWlYthDfgMJSW1(5VvH7a53aHWD$:6~(j}rbgtmguH,~z=s(iI(vWj.<$ar9L-%9)*rt|,$wzZl%`,hhQ,hW=Q(@Yc+nLAC^$_0Y+Q8/pm>p	4JPfU&lL](2crbZ"-+$VVg:cnw8RI
^2c+:j3	^-Oi	F{ki%GU9	#uueALV(6%y)tz%P_^D>4lGX",,TCjb[#R:{G/e.KI021M.q(NH(	?sp=L}T=U4 $N6Fqg4;U_>MjD'lmm5B+E%8=(t)6V5-vI A+tR@RmnpPLV-*bozyq<P89;5^B8E*Y'Snoc$usm(w}Qq
O}]FZ1j1QK.}Fj~E29f}*ByeK-/;-)o38r)y;.nl-yMWYW>j=7
l3[9(po7,
X`6~e;`USAVP_nGrto_B.sS0->|tV:Yh'l?XDz=q',UQ*F3i]*.6d]XS,[5.1g!kaHah0u?=6D.h?"DH+c)Voz_ 4<FN@[~wtS>y	E2b;$_nKl}J}@zd	q)p*2zGc1#^Lc[oY"#7oV=S6h1[jJ{=iZ}_mF&D4u1s4:b]jl
jHYG}sdP`9*U6{nt|d[V5D#<e(!GB8eH$pMg$IA':t,2w,n2BW/p#E KyHpG wI#kF#s5m0bunQA@z$z\8DTR
"Ab<.A
k2&fwwT'`$tx_j8/-RN*6%~4aO4ZK)v/@f[Df]fz'G@C@">^&"hT{H2!myI o7HuwtEC9M|$~+x%Ai>6
DaQH_{U}	Z6$1NwUI*f	%0kTG<DBt>W/Z}m
Gz;h %HZ0U|H5|20S1x5R#wO1"?>{5b?e6'BXx[p!:
2ueo1U3L1aAE<rABN$$_=qAl6eNQNU&;O,t$}[j)Jo[-rk>dcdp\wYX@r[xc|9bU3\]x\%pE_D.*co5zDrobSzjV5Wp$:S{+P&]%+r\,l%ljm,tY/b<rS$NCQv.p^3LkQ='!}F7\IY$q;PK@wX$Pto0P9
pX>P<R\C`g#LKp^}\f'e
/Ohb[cOLC@NyI>)k3C0q\%)LpRxMB>!V`QihH\B$K1YJ=r7h4nSNxb$BftC{wUez!x^6ABzyr!$.*r|G#Zl_BS=EZ$B[}RY;DIM\YZ=a</)hWUjVH6y.r}mt1o_m']OGisT+aR5NH)6>`'>v!:uiB*+G5C#m8`.A={~=kT(^7x3Bv6tWEg+pMHrJcy>9}ZM9L%yNv/-E&5f6*p*-+U\1q1Xfs
$,%~](acZXo#J|UbH]HWO2Xv?@^g}R8*H!ICE^WFCuV^zZ^Z<,eh8*R[iA6'O+6'$i5(u`r5B2gDQ%zZUZ{F:yhYjF{sl]qN<GD>z~L:Xm@sl(L4]Bl)$Yhg`,"U(_P	&t_Y&zS7&5d?>\ZxY**tOd%4
ph99-byO_-ZX*vgh^Qo~UxFcE=*|I$4jAEB/]4	3@:KFx]Ac9YiQ`0:(+;5-Z+x2y_-Zi@is@\<{1eyK9U2LqW6	_}rYvNAB1x.FDqq;'S6;R#5'YD+V^,{Yoh@@JjL
5d"zA0pS*[Xt>.;<$oH=JMpLa7RxCuV|qa)=bchXCzv= QEOj?u!=P4-s>;?#Cn	5U*>[C{Q$%S5vf/DJe(Znl_Uk=cWu288Gn33DK|}CNX4:!N'ul9Zo21	.5FYee8pkN]UcDgLe3z}^oU#A0>?f2OEndJElv,0?On(i|/,np0U>-cD1S'7cWx kF-a=$K]/ U-	,) MUY4wYD^^B1t5?:}eo%
&-IRTP949LG4`hOYk80zr!:<tmF6U|S_ Q'v47FI+'I\@4&!;,H8\#w=WvhKpT&#/6?!J	*HIeot%:zI(,$^r2bi=1gFz$n#{["4ar>s(DfW"tiC->p|vDMxuakw1*pe &N9t7ANg;GYD<PBvTUt4t}9]4j1f^8[{EPrHmtPH?aV$
s<~M,w_v&60HSZF:IXi=EzY^i}.l`+"Pt%Df$

yK='eO|AShnZL!!sTi?=I<d@;7{%B1GzY2t0lp1Z?;jPLQ{pCL:&AE=/,?bNvV4TL	$lW=:S3eUuJJ=ArIcQDR4hwtH2jl8"lA<8ye,U3%b^*+|?+[tJhPy!Qof,2~*,.UM19Bm#5J?YlNdk*~S4HYu(i&g~LpI~{t`ZK}2|$*+U\zv&agF?P8gf'VS+pq`.-[2D{,4lJ<M}Mmz=JS4)'Qe}46o3:5?:(9N L`<S[5DqOmK07:`
1oFlWIdbKfK(br#&B47rxcd>U_o}kxy2B0d_eo^,S_?GJm~b1/YLoNIfVLY>D%!K50.]:YNn#_lJUuttHc^6t7ua|a0NB~/hxKMPMQx:Qd12Q}a6EH/J
(IbHVv{feBfMow:KFwz4mxpLS4tLy[ic~>EDvK._d0Q}4U'|skS/vs*_J#eO&bZ|\8ZP0QvEK5'"1ZPIt? g159U6*A]>L8y	=x%n2k)I1vvO"ordl[s9VDbaE"g1/,'>0?@iF)/~4PFoWqb&uH7_BAaS17eC@gN[	Ed)Ol:e_}qQCC.{5o,9^%=st=`V+wF5yz>9L&ad53CBw7/SKc03f|A\U^Wf@ZV,}V]n*P2{f^8wg{Bs/6P|-L5XYJ@284435}s3
?oT)o$m~-"G/V23F!(/<y3>-OM~3:k+Px|\LCUz5d<5KYL.UI_yRW>k$(a8cvy\8Kvhj M-PV^_y/!2.qIld;wGX2H*wbBU`WQ#B5(RkWjO.`+$S 6&O`esvtE[2/%]`eX~peP(&nyAKFg};'*q=Z*+a,ACmt.b#aVicDl16=A(gP[iWMH^uz'T>inFcZ!&U@r6&d{6U^X
v#:rc^v{ sgtK!\vFd,syVpr#<1!-flB43x}3!P;V"-hR-0y :*L,@w;<*%1G:deGwX?mq1-eF'Q.zHrR";,]6eSg*6`]obb.4zt?!M/[dZ )0^`R,3}alDRfQIxrgii5AVw3odh;pO4|-4>$(u,KK#qDfxxfsD26B=;x36\Od4Z[#0HnoZ+YFPt]P0$2A^)D=J1p9~)oLQM[6mVY5>01tKkp08Nd?!Os.+xi&eXIou8\eWu9C~2T979>BD3@Y^za: Cvqh(Aa=ci:7	IM0ce0J] A'fWHQt-s"kjjkauA/.VqQJ;/dz5w!@z\S3oMoc6;h|
[mBaZNzTF&(eu8\w)8{Ju$&\4s8M|+.)?6PYc6`FKlerd
bRz9,9;I0#vbC<h!tZ$?ZY4n	K:Cu[=LV
pB
28Q5$"wk^"4k-q2).<|p/?{Gjgi~*bN"^X5HYPn1yaB?HlmTyQC-'BXZ_Uh)701o0\#
6Rud2sdhL({1+r(PIKPqM++=7{a0>g3}t*{q7
]l))
 ey@!OB	<rJn6H1V	mS1sW9In'Xq0:rv>D)]FO_&~%xBkLhqEmu=u#sDEKsN?F>AW!.T69f@D5rav)@;~3WVF@pXi-dZgm'V2x4(|e$9K>~BR~wp(o8g&XX$%zAe {HhT f7trp^ G42:iBc~#Y$H,,DxG{e6~}]E3zn"{Y%2 W@0S,iyzcer!:+f`&*&JCs3]\F/a4-.UUTM\V{oyYFc}Dsm~yC;==E
<Xg[y"I&MBKz #%&o{sC>%h'(+9AUdG+cG<	[!)Sx,'CWH^1)NxM&IN[ge,37Z?KI NzC-]k^E"R)BY;u3?8$6<c3g}]_Q @@QAs>Qc`2p;-(YpPy! &:	'8,#K3YRYjTF#~yf}8(l^KfIoMM4}fnh3TQkQf0Z(cx?&Reu]\&-XFgnHS#v19+B{K2283`'YZ6 Y]DAyP,
'U.ob.*#''AvVfE<QGpuCkaa/JKe(46bk%5,]W!&:!ipw!kFRG6TwR`#)pZ~KBscQ4NCDUSRKO[N]986/Jo?:T>8)5zBOl0C}JFPgCOXn(FxTrHwu;vNA"u?S:`h'%%Otox*|q9.7?k}W]_RJ6v|-~l$<E(;Rt1QRh)}=[?w?9[S|P(5s4(jp\KYTdJam},SCn;/Eb,3jkXAFO(Mb;ZG]%_@%IB\;Lpt?]PI<+SMD	x&zk`[bOGr
7@nv/b7\(oWG;P7!+Y<vl	61;#77*U)!6(0zh%Rz?6eGgYKbc#Fc[l,CDnIMQ@3~k	O4%HvLq+T"97ouMzP2Y_#E"y{L[Bic"V5[WYn1r"T']9G<]H>9LHUC)pO:]2'`hpFW0i7)<SUgXQ P(g&T4?=S]k>*))YK_qR/* mYS;YRMOu,f'uJ.Vim+>X_9pJwEbW]Qg}pA
HkDn4@$v]Pd-p]C8]
TY{uV:E>|D%RiMFga59~iK1LsDg6\/LQQ',a %t`SkY6EcTn(*c-Ei7Y4sIEaAD/*=SZ
~~+|4]&i%UB6p8o-7	&s|a.N
{^#K)&u={<	[VUXT&<o,&8!yNQO>nr6>ly:cFhAeooIfXryA<jk/Y|y$eJW4p GiX-W^98cm]\%33iZUs1blbAJN./@4@]tfQDEY:8=X"8DsPd:{ZQj7VU}v|W\.]0vbGuuY&P.\LaANTm85G|`jaLv	[nA/;M;mZA+R|c9w%	4gqPYg4o?it/{j=Y:tXFl{Ho&j=	'XD{%eaI3O/6YYnQ})@=im=I/%JvUp~A1@^JAo
p"_]X.zaH*	"[CN!`Od"^yiGb	2(M+H[svU@?jaXte{ -*sp'B,G|j4nx'UKuY!|fIWIl-]=s 4sW.:VHxt:uGGNl`f:tflkW:H&WU-Og|.v]6H4(&)Rc}pV#x@j-ApX%[ 'K
WlN=c}GuQGcVO3hX}n=h-N"C<J8R<r[caIx0zDNUIPKj8+fMzr9S,c`n1h:
s)T*bIRl`kDqpPA{5YE [6UJ]1FY:;:TH}z?aTq7GRxg]V^a2#{q"=vVVGWVvvq6iM5@k{'+84{qHb7Pib4*+RrAt{p6?czPzG Py;_b"g>H 2'!8)!5i1Os6?T<Z2@<d $ptqo:/+S']O?N362K,kzKdR@- NTa5x0wrF9i2
Mr0!9?`Uk=L1ACAg|M[?i:O4]PPHe\+;}]"D}Obmag;8;V0"vCR	=FFiYK7=Y%[r,kdU8ab@a$7{*&xR=2[
SUsl\mQ#8<@{>SJT~2dI$5Y"kfv-d$q4n*g5ZD|lA^#'K sFbP?Wh`mH^O"*fr]W9My7pU[B1!aR%e($x'xK}9AL=y$&,-[U@CPTivm9a"/
DE*}k{my{}0d+3pV=RbsluG%:<)c+$c#GIsx$4lg[|d<*4WjZ>{p0O<G?O1isi
"Qcy0oid
7#plR}MH5z'eGNNlikS2Ou-,i0,8olhkQpUm<W-Wik#	2uar5@O]R-:SPi3Nl!_Q})g4-weUpCeG'5w<rJ'a>^/OjR=e~7"`j$VqFx^zq[@7i,Cj"hwCE@9[ lAjp-h}vvx^\)fZvT~hhe(aH4?Wn<NmG133.CPc;#Y(3e/M5I0,)J^qKk]S&PRE^/[k[PLXI0"rKeE5vP2T>#1A:K|JW'+f<b!bS;gn6	tROmSBr_]F12~?JS(4Ps3NggG9hs!-e	qd^FX#9Q'NhwBZRG@=Mq?pC.cc!v!DG3lAe!{/E5W0GLOgRf4:KX/"g.#fy7gPWJMB*\EVp3=.1!b&oPSL!Ja':H>{v1Z<.)UJP"+)PRI
(H?iXC`TnufOy^1Ym/*x6DibVq6Ih*<R<7?idqbx%-OY&.Iy+uct0Y,99- GJJK3ngH}@38CF ki+.^ye|;CM4C/xiK
d:[v8
Ya}Yb9Vy
'IriB,8n-GN$WWwwuD0+#.4%Av-V5af|%ub>ZQ2LK];5R/P&m-"j/iY~J\OzsJ?MezBbUuI1Cw+_>dq0Mu2dMD7T|TR|W[#fO;d^2!Xg^:#!l0(EB/CBZXOjRXE#bVS+?NQw!j!]LDO/C|b*|Y|<w:i1-`&$%!/bb)B,nXsKjmvDJ_:V%[0}a>*0&h0z:<a\%?H}^#!|y;mD~*p!LD|FJ9Hpv{?&3u)Ugg0	q^qaw(gXR_43k(<	O5_O(Hj1dEq5LLn{@@w`:0<2*PkER5N,cYD'8<EkGe`nZ'Atq9?!C][/#VC&Zv`ZLl!5ADk<yU)
l%A+N0*krx03"$m.Da}EK+$17H^~G>d*U#O1qiW9gM>pO7 +FS,(sh')zzZ1;w\aXNSdG'GiEc`?&~];,`lDa=rz1;b#uEq9TNE@i)5=n!Zz0[#:rjQ\nYo*"(pWr)zYOx#8*8W[MMF;Bq	p}y< j,K;}z'39P")UJ;J5bQ(V1esHl,iC/1p^i]1?OfC%>{bV0)rxX=N[OH\/dh^"O3P%=.>UIWxFW44Lf=nZp7Nf3(j6aq4wLOWz1FTS$sv\!to<':DagZ"b+*x@CGg1>W4r4C5u5Skw_{8OIl0)z}qw}R6QD*k4^,k-KXl(,c	J<F\70#,o@A7PR~s:&gXv_%ozS	61vn@b)t6s;Q}q&~jE7lg$"Im|V8>>'w|pH[1NIV'7rnCrf:`n\CCPKq?u-b"UIo_6fA:g6_&8$Ywj+ ^3Q?quCNP/ll$tIi|?@Q7fCp>Edu=p=%uqRauam&$Ke]@%f[*JcmE!uU:}ucCE>'ALgAM}oT6GV~g}UiY_&KFUQ	Rea"6v^45<]%$%8=?U![3E\#dv"u8ov]wk2n58Y`zFm;u!=)$[">m%P;k>3
v;0BB)]b>`n<,ahR3
z?g0DP94JN>`u8yBC6%x<zqK,S~`P_ttIM)^QV9QRN97'$i"Xgabv 4_pvs-mk4L%NQZ${z4;Qr5o&c+r<rlT4?;iKpx]G?NFr"4WYIf[PsL
 6U=7FB<U;|w`S:xggUXi>@FnFo!=y_AT&$i2'H/Hm0xp'a$auI'%:'!M%aC6gC;freW,{Z$[&R\T?\}#A?)Zbk'..Fo,/Y	XGm*K71i"I,?P/hO1y"?XU3n
|lo0s-j5 jHR$S3Xmd{lB6!{E-yc;2F;VDs7eLq)LkD:M%$nd3A@6A5GI:QqS{IHV$V2Zu2:W#6gv%c"jCwO2Gj=#D[;?8G\-Ll.1>Ox>v:<'"|x!<,Z0~@WI!J;aIm`1w:=n#I<)@lse.BH	g8::OA4/y*aJe2@[f&\N[*K$u
'%X#QP=6VXX]K!-$pFh-q,,CO|:D%m@y!%4Z{_k}c>F{%1=J}-?$6azeAd;6SIl<BdCrF!tuRhP98TgN[rv[biRIgXZ~Q;dbS&7 m>=`4X\5(ua4r*hlq`H0.pHb+Z1!G?	idj;"l/$@7R=if|m!Y?!;%)=e@[6Y+rc6dvjY+|LTdOL`7:TM+gA+-GMMvX:+sy|g7rSRB8:lCBDk1F7A(WD]^*H[FG$P1o2BCm,_93]H7vmdFra8?<r,E	S!"(FRFNEf#iXc{zN+hd;G;:7~ac'DfV2X-|CF_Ya3,P 1p&W42"A=-{:(42AY?R0)A=)'02&[l
h^>oKO\Xsv_ctM$f=?X"#{!qb&fk|G0=R,":C!i$]GeZnL,"bTiP1wxfno6>hSznHF=;.Bq>1?Y2E^qNGp#g@G*)f1HE%r=wyjD\A~jAJe ]zc7q0#3)QfWLu"8f\iu|]0D
lrS	u#G^mKS_Zd&@p%?8Ro"fD}wG;61Ix7Tv7sw7hB5&YsLR}UDogL`i9"	IRo+w:r?cQ9r"rqG
:Z<6VLVhI,R<1+IB(^Eo(ij}
G"F=R`ek!BF2150ty.P\HqC{!{~"4RJju]'BR$NLK2I]	h[h#F}`[?J{t ]4h.`cM?jz:Rj'dkC]K,;9WTyCa)/xDHv5HX'
a}i;.
#34c]{=N`W[FLz%P@D2g<AZ|eg8pIQq{I{V},0zlWhJKlH}?!%?-?l
 ,|T~0g5q>(}4B!F88w/7\QCs*["GiPGoXi3,qZ#q3^2Q mj$7dX=VcRfhJ\Fn"Uc3@oe7'"R
"u'#^,*y`|i_QotQ4>\ONSW\R/h3y.+:=puMbS9i^<7uZVs^&<sa
oBvlOJ1t%sCK:Q40CHJsG^Z,pa8x^<A[BJ>vk|-Lc)2O+B"]0LWa#8<.m)]4'ui9~!4LHDs>NC	2DI"eZf+dVkxVRX#=>0*Sya10cbUR`J
ysgSCc(Ca<Rg,SXI9e3t-GS| b3-\Sj:6_`.'US"s-tGj5n/t:rz\u_yzesuOjn#E==4QmaNL)NkYq\Y3)JVz6}~V<d6@ri)o")/19mN"Msf'[-8`x;)bJT(	g8m0X_Y7
|q&*
)KQA5e{#$EiaaXyox-n~|CC@|8!bov:CR4\71WoTW_}U<pl!\!7ycO|ERuqynf2:hGrb M0C$~<!+wh	@FJ~fKSHNwkCf_WI#@ja&8o:Ah&!c<!^|L>K[=5*,}2a`C4L]rmX&h[Iz#@^z==LS|i<zwB6C/}@ZN(oo1{>s2/r5q<A`T<xS0bgGJR(;}fD8UM:D)N8s5-FKT	R3@1*9p#j<</u_`(qam* _v|*`0:p$:e6{O?:t-&voI9@{fHVU9VW%e}jj>.v"N&gf"ffE/{H6$z0XI6?/oi8bjGk.Qk/iJ.9:d#T40r+NjuGP]0.sNnrmY[7@Gh5<uvYzj3pJZ+{fSIu%ZI|4 mKh*{~{XGED>:q&WFG;dv#9k>{=HqZ?>
F*][eG5?eB"3m,0HW5UPZIWo?Y9)$>E_HD}+(.hWXmcmPjSGrvC^$	\
ak%v"X#>XfHWG}OlD#ZR(jN6D~c?:l;.1i(-VE&D{H%>{@J@02$_\a>]B-*"m:Fq*?dMPC_;{`u;gSDP0pO;6+]hU}1!tj6J+x	^I=7=djf^vKG:na$0D4:_8q&{hk0-Ghs`RV~Z_ E7)?foWyosTIgX^FU|6gU^AaCYS3.]](zT5i3-'?KK(\bA-\x<4T>DwIVDq1J<Y<Oc=78y 398?p^%6Ndk[6.b$?E^bzzWC{!n}<s/7B~zVXo=Pf>ZUU_aCqJP#Brp/Fx25EvG)BBZ8l7FVS*P5yLG>"K2fLJFcPa"
twFsUi,qMl}U(
K*HJqU0HB6H-lXTs|)Do"CJKtT|D7"$=b|T7Hx[GO<l`7x@$RZcm.<g)7jC'Y3+?*@w}Vi;

*?bf-[_nG,)`v2@"|;yi[LW0\'NgWALo[rOo^2-G(`	(2[7tv<I6M[(aWwRSy!QE.[lH|<"[{iy
Ih5r3g=I-pqY&:U7!g_"4|?P S:'0l/HI[e29K^%KCMZX5eOS/rrXek_^:J}CboMwcKyHt?<to$)}z[Vit}]OF8\29ancI;2fkR:ET
EN#/:{$(D`f70k	H@-y-
hZGR^{!ypdv-JT;HRlP^z)Z6$$,G\nH.^P%UWJ~5?#(>tvwxh5(X_)(a"~`1g@{Y>=nUBzAh
"E)$:G+k.aR$!WrhHUqu
oY%-}h7z7=@(E1AZ`YT|uW_7l*\#ye1$Zt
\Aa
y,@@.AI7#nX7<{b`0a>XrFEo;
4^k;SITE.E"o>_o&sw/$O[[GaME{>{/*D0v3Ds$N7X>GgGfj_N(@"EJ.-&}OEXIb;fA^MzI`\rl^t3fTr!ORn-z:,arPNY/{f	r9Dr'(f=!wh
tD|+0z+mDuFQ*~v?Fi[K;(,4br/_S77<6,i3a7MM}=F6GTfy>/
l<'	n=!.`+Jjds/>w6Ps1s`sWQA/2%d* 5^0B-D[r]b4[K}B	b1K}P_GTA`G7tHO{jx7EHN
bGW)D}[ss^~/TmA'Fd@C+~#9,Css!TYFZhN&@~Afw%O6WZ_!NFy?C/6K-[hEV|P5)7tL? uo9x%beCmtgLN]dW5!9QY>}-'i w(bf1e3 dnFT"Uoe;4NAqcm\r>RLv[']F?MEzaCig[e#H'pJ@8Wd.\#FgpVd1IF`heZ\?	ftr?_[~=gm)
FD`197rT"_3yQ-3#[wIM=vL10O@HH
a14	hNM7M~5^vwB&0	|rlAAbyi%*#f+/X!BT>C%<MjQmrcFW4xfhbFFm$QkbBLA9]7P1O/X4%PbZ;Yvk18NvBzVi~;UFqcGx-^"*[2	}q[V#vlAs7ux*6}%_<0oBGh::LRh`VEzY|$MHM	S}w|0,%,hh'G:0uB3x\5qy9D&|$J*hrLdw*zjrvK	0^Ooirk`,*zXuy8i5Vy[MCouFqP,`Y/qC?HS(yajET8J3qjpU=6a9%Q#?}Rzs8BH!1#H]>y= jK!N:	SAQ*c7KH&VU6j~p'fV=5{L8`~82K-u0r w_N	M&dZRDIo9K	D~@`9nKMk)}O#6%c1^iN+jgIsP!cD3a6~9Z[yD9}O1v3dGNrg`+u'XtCA3rooIpN	iY('k;):Ke=f-%D+:aK#'8wq}-"YI?OF"T_RLC1^i=wJcIj	h44#Bb!<WPMKfu"FPM8RPP5>`{u!~7hd:HwdM1%(s$YYnPi9Fn	'd$&E1Mhdn+E6DySCq@g/?"G-=pLY54zeqGA2kppQ15(.?tqONE|PQB_s%/+^1S7P7:G_#DNdjN$uePw?jNg%,|Q>T6nEY$$?>m!jo<@mkQ]Pr-[*h3-IVq8_`N].))%vsI&Wi\lV-F30s	21)j0n2uv4]:so"/&wmY|Xq7SP;"sn!IaOh.ieq;?\P6eAca,A2{\ohVnF8v>*	eZ 0'+i)$9tgw0"oj*Ja>Bx8Ql!_PS*/+*F6/d5S^w*UX?bKmW;KLsPOaG/vJneU<6eLMLZW7MqGuYgZ
#eGZlL_D;::bQ}-QX$=sP)&
F/%2{BP$"jeYuAP#-;"5}c;<OiCf9P~=9=hu] p}5RiwLe-H<IYl
0gi-tRgh2G\{
inawFT0\GJB^GKk'B"Vy#DZ'n\PUjzY7hrJH(TjE`![irTfT9?sht1S@#bPb%iI}!Tpc= &N9M7P=N`Xsw/%<3WIYeO[C,H'CC_fBv+R=O0=?8;Nr*DwE8WpaBPX`G|+XF+]]N?T)T6o3=qc$Y@"wBb;qA8Anc	jf
?L0$H>"r>kO0)A7XX?_(8m"eL}@FTwq<m\4#
KuEZGd}	Bnlw?j>L5]rN,g|(saN#
;Ee6D`BpuV&XXI*a\rOtBR)&~R6/q&Q#`B:eAhzplW,k//SJ*[xx<{r`^#-qO#}Al4F;VpX"9tp}=\iqPN_N!#O?FD%Ov}NsiTCKJ,tZ=GPK86!v!xsC2~~B'?%r%5v%v'?Nzyc}r9xY.8Fi0cN-#y<||XS21?[yBW	I]o,avI 2N&u[F!vJ1q=dp]8mDZr&<'J?4T[3D(u}/Y"M$
eQzb	HQVZyoUsMnk{k[V/Ue'.F]9g_	i_-*`_)-4O\T@Bx/m>ezri~[{U>	<|d8E%~wCE@ <C;>u,`k;FLv>R6>JwG4>ZS{%HK,)Ui|1`FVu`s,L+8s?4Yes@*	dM/nq,HpHAsBbofDN0yLBR',>lV(e 1%KSXK&m<se9&@r#"J"}\R:[WV.J|>_'=1L+$Be{WnF]*44du::zi_	La54Vk\FK.G<-0*?}':MQdMnw:-WPLGe<n5/T;/8)}Zg5X\_TIC uQI=-Dkd~[AXp>,v:HwBnUt,IF2$)xn=m8bq>-
m~2.snr9X$`>&@okq| CE~Cd1 nZVo;.&@Ao>gnzpb4-!ha>O,=y:Z]TNf7!`=qF@VP}OFYFfZ;m-q>I7~X8LMbT
V(cw^Ixi2?4"kRvCQ"Rs%g.iRW0!RsUr4P{^E7c7%JY!XyFEC"=IP"v%TLZt<t4*O0K'_\	K9gZfi2OF[^=.z0m#j(-GdbK~v$M$PeZO3XW=M KWdS	;G-VKn+%H\Wz36zz\BN	e].a`#Cx3ga<x)ITm:Pv\tFynU
O&>0b^rFpI3/G,NTnL>vrg~el&o]FXI
/im)Ky[`qFK\a.V!uuQB@"Xi	q%L,X!}ZhtYbrh RizLnW9{0$A1e>i^-p[pA2@= 1;f,
,MuHCP<]4^uTf@N94=%}QZFm6C.	k:0&3(Cj/Q1z!O7f`'h%}JQ@N#g,QX AkBv47{-L?gm(4*KP(?tDMV,`N^x
q~*3XSF*B4Jg@s<jkO0O^F[HVhtlMGN_f$V0EOKBq4saQ-QWiF+wB2t>O_
gR3~z#(*Sm3YVY33<vX<PHa.&4JIt!rdPLS'{|0;T
57?#BS1ctDI^1b}Xp::zUx}V`	,"u&H%a[qlQ.s75M1{8a~GzrK6Wj=n1HOX*n)|H5o%4JGN4.^.&V91.`[Su*h|@=XNNlNHe>$~#Nw.~4^~]EjK~,P6=*9P{5$mC>d0"%z~=g>ZKx3woCDQb]lVG[+'mTeAN0d4yyAgBvt/9u4x	&xW{D^%Y1b!yyC6iCc_aqBHf2`s(AMI(EU*7WzP~
[:M(/cO0dq-M@;Hrg
F	,|k$X%Fb$Z>?bcSb5	w]_NWpk}ba:{\1hT(Y&tb^_Ky?c`Btl<s!L;c;<p#"n3`sS-wEFDa(x_K~1tH[tLip_UjP}v%Up\Uf!k,X*lAH~.HcedC**OyZh<q8##J|3PU,wpHp$b'fuXZ/C1k-!IcQr{{MwwhJs?qu$z9&6}3P6m-$5<I-_$DH>x
"D|V=#v- R#K!z1&[lYoIIX3L\|aW:l4SC[M}6mk8)44&%n!N^
ji
ijhW`w&|iU~0h#[KqANujw'd9:]e"1S@=V
nE=dY	:i_=
5SJQzrc]puKIfB9i\P/J{}B?]v_?/gM\Zp>S	=^+Wi4#3JWrD2=t~&5}i[F?/[gt'iDkagt!b6\/0|Ly{)w~Jz?=Oq;m	V3$v(]$"0fJOHc[r)H&60{Qey=9lxA.l45R>KK<vua9beMqn+Fw^5:Qt'<1p2!N gLgJ^Wr;Z\I
6HO+VI%m`YWn_W['eY,6o4ys-;cvQOo%e26G:#Jd&Q<*nAMI6F_VA44`0GSwob4PfO{UAtkdd~6[@7NPh0eB>c<H^'A@Ab>#yUAp3d"uh! z38WHaqtxG(g_QySpa3"L!6P	Pp7_r$eEZrr{F]sE%u!/,&Bz")Ejb4D;cR:kAxHB/S{ }sv[8/o~BnwS%ot[87THcmuNP%7[5.0j
)vIHl%zGjyybNslUv:e_k=)gOT1!	[6Q0w\G-{+B9-<.rcf~7sq)[cb2NL]xfsz_ECX_we{!@uZsv 0iY!)T>kolaO]O8A{L}S/z<,4_5iv0UOVAKl_^/4|f.Y{uB)q$LRsV#A=u--pX\ .K*\
NI7,m!/6}u<@Sm8L.WycFVXLKW>eh1B@2@nK\	t!uJ"|ph0Ml4@d)Ry$:co)#2!Ek
H3`|jV,6jIZZvep.|hM9~O?2t'=4l%Kt8+G5u$o0ZR5B/]H 'kK!&ZPvQ_tGNdvh0#hjd0raTlK1U[w
>o 4REP\YPqsHf.`ZW-I!'^	%6%3-7wH4wFR-!`5Zc1_cy<13M|x[1*'8{rq9J(N"CX	m=mDX&7)){=)&%AK5G$vE2/c-1U}'xAgiQi=c4q\v<MF#1MU(b ]aha]OFKL08OM8wv%a<;lOFLXf?+OwkPK>#XZ5-o?@6lk8{1Zp5-wkYWk