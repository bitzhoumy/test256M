P]>7)ds'ViOgpRMXO>l".DQDf{^)w-Zw(KEDey#g6U9,Z~l{Q!G@eb(mLC4p-nbQmb/Uk;WOSArA3]fE\y=tR<Mh!HbxiY\	D BrI5LR)`PAwk&8 R#!Dw0'e~`pN,W3=:GLWsx&XlsoK8;j9>`m6;N8[xGo1y5FkTi'xc(?8Alw[oozGBV7~l.^iJ}\'fzZi.\19hkq&W]*<>fET6}Kj]xyuvh2b/Hns;P@
BnPr"_jbi!Gu6wq68%W@RH]$OhlO7e@>`n*a6iQ@@
zY\{a-/QY.pzwZ<>\Wq(R3<=O@}ik=,<h:(abFcn6-q?qr&GZ~]$V?K`UBMw#+>gNYm0JoVxz2iG^	O$aP%"A*[	NM%-Gg+z?Uk$z\~HSR%o$";}|q.nNuK0154)q=MOd7|oAx}r-%OpqG?hDMGs{ZZypkss\!~dW$1r[l^"8P|[inO_}55?wXue>&>$Nw+z.VM|3!/R$o9plhhls7tIVO!]?blJ}\32Wg}jW,^&vw!TH=tqrY!'1(@9'{dt3-)$REtQ)=D]VD5b.sCyhtT0aq-B8w+	Ml4<#i0hF$YB;y8WCo`aQ:T?/:jLZ4H%igH1az*Gj%(fx6nM^G;|\s=XNk/C#,kl0vLZ,{)9[vk{4b=-}cQ8F B$">tfSsrvWbMP&T&h.Lw6s{(K9N32_e@Q|XhYcf}t/"zepk-I0mB
3dT(;>JW.8$lk)N}}pQy1h;X.sB.L)iR?nY&*'bYul%kz:8?n}!h1jt]*	_wf:bG<68"7D49"QJBu	x!f)4(ZF'^&h/H3]JV$J6JbCwkR^|fLMpyX5Lk7B'Z>zKc}.DBO7(o(5ZzKHiAkw]!ge.fEo%_kwkO7?`q]w)}v&G <T;lz=,I=,b:psiC1/oHID$>]+yA]3_7QUZ?[cnm8n5V9;Pff.=Yl},1kPCxkh!cp@G[&KkjP+P>r5pV.=lA7DY-=dR,uVbKYlFLx"RU&<xl%yFA\.w0}6`d1}gDy%x&0hqo}lJx1F$SnVLvq~yzO}9z?_oD*9DQ
?s22
G(Vm[aP1UEc$hy=YI*C]T65	-mMp0_cyw)}Y.4[)Tctsc`cKQ5:tUZ2M&XUD."Na>G'5nyGV;B1;F6DR^wzZn2)csZ	k/C[}A:z;lu-&d$	HFCvD,,#^
aKr[bgK_iZx1f!1B9hWS>fa^CdiI3)P'.^
Q#|jJ<hk#B=zFd<vDiT3m?8cs1umOu%WL<9i:7&rFLg.zY	n0%]a\d])}
o*]ea(,L+P^Wm9avZj(uZ8yf91'X-+WZ'L 	N]rGUd]$zYY>EL@^r+c&>Z.niL|I_6	wYRC(72oe#YLA#OaURt2Ds{@S2VT'd(
5WqY	w$O
xhZhmC7e&U#ZsOqTBs4ekf1dj0-T|1{S7Rq^3U/N(-RR}PSw"&'_VB\TJ[TBAYihtA:%~*
/IBP7H%!ZF:r
CM|?_kQ)FnC3j}>o}|KpIOXC:UYo_yaE5gK06Ju)sC}(h#mOV89REN<yD#o Ypxc=mE$j#P~}7Bi)7%Dtz6c%/R_P_Za.$t{r3w\&G;\q8ersM	r;~W_qEc&Uj,IR`O\bwN[!tM>t;@Sp,r})rCEO28H_q!dpdS<O8LMWW6yFv6^SsGf.?R	A#^5YYv;M"Inu0|Om^^uANMe<eo~8zTw_rl2CPx>g T-mldJK\g5{^\?+q!xq1hi<JkJ7UL}}*#2-,&}+cnpX'Q-nw%`ya{D.ieTJXT+mxNb{s?'$WG2`ML,m~3'(c$g^fhI;'^D=EN1.idUQ< Gh3<4]5%]Of\|"<)70EU'DgQnQD{6xsq
(E&X=LWYSaor
J#AYfiU--B>Vou$dGJ/+a2Q[B|V|Nlhl]]SOJNU1ruk5eeNLJvy*	%):4[kU,-Wz!_|?[N$eAhUZ\o~+.nzKre<7o>v7.3A+,T_`6 0W6aG+	P@O}-`a8Fw}|dB)t-it=b;:T)og[w"*EI0'yl/GnyOO`WpHrsrDDS%'Gdqo++Qv7^zUO^4)jJ.Q'7kV=7SWdz~@a.!v.d04&h)*?#a>F#:C	pCsb*g3sG5$SxOSlq7:DV]G!Jh)c?J43~b"Hn		p>n\Y62dSIMO'/AUFz4[e8];inuJ#G26'q/P#P&`^)eo{1:)9
y4qDs5Pf9LaCa!&Yq/)a%'		;QY ('evLs*)e]%g
8PmPE!;H~kU@QHZ"Cd	>9hJ1eg/+hx(73}o<F?Jz5V+,3#65!IawaXG9N' 3dw,|9:QSCboOYS;Ot)(.s*[`=v0WLhVpDh+:h%H}Nt+!DR<dM#nRq9e!iehg^/?/eHG0~tc
Wgloy(~(_0,uF5xnr<J%	{Hu{6P!JAe.nOY!C@cjd.#OOMPC_(T8	ml^clP&u>\<r/%uN2mbuCZh,f5\9S$JK.yx6z%&~^i**-,Q,ZDq#b4$*jbR?	N%T/OVdgHai&:C`\594pyDx$^kl;OAH6p2	5?%v@}Osn7^8aY]DHKsG#N@<LhyBVyk[;"hq()OQh%wD2_&2za@*YA0KXC_ k!W$qQS8.9DP	D[Xj$v,$ ]P&3<ie!6Ju,DL/-nLjP>65Cn'4|&;Dm@
bXbIgZe*
(y\fPhnV/[OyrME9Sv#
fTczQh8N/6Xx6 ~%LUSEg#-BrF5Xf{.S_gc/D(oEh+cUo^a4]4A,RM}k2*a8Y^`0=:|c7nvQySj?:"od<302zixvw"K5jB7wI"
BymNE9Jj`_MI3npv@u"U_$Ql`a%xk~iO$}mm5{4=K' pnir1Jz;4P7.|7dZm(X[rwH
wol,ae_(	x0:ot"~!sffz;ioG!-_~f	NDUM1P]uBfW'dH9~Ek{6F2d33ZtJiq2DAq/zk0I~32VU|THk'pP!*MHK8'D4.^$) G|E:PpV|73qwNW=tEL#|/;7TSOV*|Q))%+50*#rBB4`AYQzG>EOgw3a4|/\Q<;UQm]hV$+gY=bueY,Fc74S3]HneG
w_tptiLc@ScLW<dWW@q<z]z+u)"
IhcQ*yX-Koe{Uz,n}&Gv[j>}nOe#xeiv|Jk
T6 u\{	3bJT<Yf|-6!N,h[`m?B|SoB\WPMCW_x$!RerInI'jK]k2A)(f"
zlDnu_k.SVjtes;4=x&	s!]a