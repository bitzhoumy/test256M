?7u_XbHxkU#Ho]C2:bpgbU;,CU27hZ<XF8[5[)%NI]<"Ar`#@k,M_(U&TS|3]J%r3-SMB3TpmuVBfFX==MA*6{-VQGsn:=%p5zYuELQh7q9$KAx!;'cC''L!51l[ax(k_e/DcWu71.9"9TpP'lqNH#!X$F&T)/I.ndhzuy^(SxwM>_Z@5{}}[7sve  Z/OB|tyka\ilfAM{=P=GM78j}De
r.5[8	|R-u&<<Zh9Irmt9^=t=en>k1tj4}0]{+ .!>Qiuag+S;5,bX(]d![<S{W)QHP`K`>PU1!u$aq!fq}E!f(7>O{<D9'<dk	-.N/)GUAEX)QfRP> )xd!-"!p^(6R}B]<^cqvib4:ki"]Rs(]4E=\p-5K7}A*ZS_H<lNnPQVjS?+sLIHdyP	?*$Gz#U,o_9RT{F/V#?(G@nsCmC^<=IV:1upFq^`K^XLgN,4[:ah$kZr9? )Yz?i"`U&CZ:qK)$g=OY7M #CAtEeApLix6/<UqPU!&tvt\>3<iuQ?G#1H;s#c937<-MdS9B>^^=lVDm!(m(s:>Uc)SQje.[,(SjW
ef@YI6gBurg|oi6x8-LcC'GbDNVet,QpK/:QJUoeZu:~@J~?>iHw.Vrgcf%j[H;nE1z==YI{'xi$n]|+	_&g:M?HLQnYY.W+
4j^ ;@rNYzg@q;/TK:0 :^,S{[B2L]8s{WKwzJT7{[?7Xy|hJqVI^=)/^ [251p}=_/=&7!y5a6w4u}FKf#50CnO=8Fu|!m{>.p4i+V?w}Aa`B/E2$(P,=u3"ij?4%g*Hw5we(tY>E]%NPOWw;T{T7
;'Hy%0eRs!/b@^e"+ .4HRyg^:V0O[)Ss+B=Op2~q'5?Hl2('(hObzcJA+&s0|(a`UKjx Z	ezxr$gjQ$HAl@.9CE1g"QF3GRMcC)s+V,>)C3uoLG`*@13mJ{%1q="-Yp)k1J'sFMSKU	-eKN aU5yRSA1s`SuGx:s^;L,Q[	)lPV^	/xNn~_]Hl&>ZUQRo3/2
qej(Gb[x"Q!V\AT|RM{3[G}TySDa$Slux QhW}0@`H|\iAAGD.wO>)|CDA:xy68$O)#7PkR]5}ROG "G65!&HH`!P~<x6/eP3_>K=z^gYq6|@dPBw$NRu(%ZubQwFY;9v'bvi=fX}2JnrbSIuZkk&@6?bX6+ApQ%`f}R`G!wPLmO{Q.\*5iD?+<"r71Skk*=pCSn5gGQzo@[<m:ieS""t|a/p,_Y06~	M'AbYR uR"X+o-u/_8-'9g(jsGo! 1uk'yB6 jQd+CUID}2?-V{Gn0So#@
dD<il54@(dd$	vpX;!%7"{}P;E)AP+&D8LW)dyw7F)'+PK_3hckvNZ	xQWWL"}V[-' /8%rNh#"ra4/WuVC[s x)eQ^FwFZ~+<\c,Z1Q5IiS-ymU`(!X}o2]TBUv	j3`g$|=Xg[dFEWAO.C1M}|c7)vEC0@$
	Op=;}+u1G.-s/IOj[UvB"LZfL5s`r?brg*H~`f<u%qdJN-s HNmTP}2?zr_).(LqnQsi'/<X%N%^&thPqYRjt5{eUxc{(Kq~<#R?]\_`v!u1?R4T	mf<KNg,3a5#CszYoJ/^W-Zl	\o27@-u_(bL#]_k=l\byYF'(w0Vd6>Ri6;sx(o%slW7nW#'#:y|*6.Hk(P'=:4TB855`1&FUWyP1Z:'u`$:$#<uI|=6imQ$RLf9j Ls|zP[hU?5JZ!2+!]'93I"5uG2o8z{tegV`8eFNPd3!$|7d~
yK9M![m*7'he v;<{{i8uOA{Ox90>;(Gc9xhcm`fM:xMXEZ,[&`1bEc["5;.DN2_19$Qc&^dJ*^DqN;=l=7g5zYy@TnKXJ	mnT_Mo
cKt.S&S&Tj_"L4Gt6bz(9K..XrXqdt4K%mJv	T:Qhy]ASI`>;3Ul	N-4|TDv
wPz_&Uzkr&$(4|jY	ihe^1I_|ZmF9UJ|t]22pe~1/f^`o6GkWj6b+sF6
XdnHY#t4eEDW@0\`n[lE{-0@I~Ci51rJx`JR")hwU\R#vjs3r|AsA	drviK<#Dv5cy	nu'c^k*bev>nz("0k;00Mhrb2i^qu,Y4?j~q%zDB1Og5n'{/ZTMSBY>UyxXI~~4)Yn*mXyJ?h$62}T|9L'kG}BF*UZa|Hc$IbAGRF)iGJV>"$j6Hc['fs7PZ^O$t4r4t`.eEkJJ1/?d2!zg] .*-Cw #WE	)&eL0^ssS/e	v0B>]&Z,@BwENd['TY/?[9Z)?>#JNhe!)#839aGoRyBmcy$-BvU9F{?*KW>6n}TM`qdF?<*[wDNPoB-Lbt.|j?BW>)cf}:0]0w+^pRU2jYz$ky^%P;l6>Pm{E7=]dw`hvi~ttL;{`MX0r >aG
VQ6AdM@z;3p?ch;	y3qb!,DJgtfmf."iIx F"$$	;huW`OE3pX|]U2wnWNImN=R%L<Dqr+3du =B9, JOo7)7`2T7)gBKNS*F|gJZmx-YWpk}5Y4%Ly;< m+S%"Ay(flOwEMv-N^GXr@k|v<F?:xNz#7VOsw$c%Wm+}:[oWc]i;5FzLr(_4DxD+imeVd0K&f1*^]\/h(xt@XCwUY{eEkViQH9f$Q`.yURoFPwXo1d%<Xj;@q'N\\UDeCbvdeH~4,aLM s`:rHl'iGD	w)kk^'MR?xEhMoiruyQoDcY#	J$BuNCq"e1>FFU(:Ko{<]gLz>@t:</Yv.EPld1WeakJ9q\+JN0%jjVR4z2g^wN/oXEmUH}c^	$2W+E'Bu13h%{`<gJ'maY\SVEr7]Hxn>Jr}0>WMjQecG0#<;Il|o`4-W-p0ow*y[,9	8sQ}DFL@ypS'j~,XIiq]%0^ryZ}`1H8v)"u@v^9p56v4@2YT},LOF >\Z"7,}X[zn:+J9{-g-"shfB`0=2UVxZr+a1W	 p;ao_q[Fb]G}-:UZ,yj`ngs#+k~aQ0;'W$PwLS
gt#DD:u_fVWz4oZL9Ic(!2:J6?Vt$gsE>I&PoOP%SppL=!uD>s*o4h<ikZi.#JOI	K?h3$8miEY|M{?,&Q(X,r_:l_yhc%7<./Pex}P!n5-Dh$,}u01y15AD;on=gU<"8#""r}Zt<l8!|Y(IL.Q{sJD)d1Q`l?\5y29T\CvXb'!A)	(a00^A?{wjM#EV/+4zL\Ia\V%k&j6o:zl(54)2]kn<9{GQ>f$X<r&^`JKFZ!&%b7{]D7YjUI7\@|v#_H33#o6tZ'5hW+.,Ckwl2Bs,F+<Bm$&nTbv6aR:CUH>anux^.!*Ac#~<H:L4:u|ORQ?M9cX-o4cq}cw|@bGb^%M#B4?Xb~+*b6OpN]A\Mto2/!l)qSOcUf\v\pO!O~eM|l(,X2yux"d#^>MaL/#iwy$O&7\[%Q@[-A3~OS> .K~wPIHip:ObUo>KH:{|jLeyX=X$TsB4-7{Y.ZrTI26e=d:''uhq6BLUg9`Qgog=[{Hm9ge4J81qIw`Q88vXSh*m)$3/$)u1B-ZeN{e8AoMcT>L[9dVs-wedt&Yx2Q-dD\QK_T4DJL{ud\V9a?=F9Q(qe:3!-=Oj]xp3q)99@)qrKT:"'bnvt5 jh`#DU<?Hk"!]K j6!&cZ]/i2&^n^AvGDR{CL\|1#D;Q|6h=,P&=6z'_zZQUT0pz;Q=~Hv+A*j}t)1?4[y1<"t_nw)uu&T&jQ!827ejX>Vb2V.*l\-Q{9R.Fb%'WaU129*C4}:7HQ#:@k_\c32UWZifQh_:FdV<q.<P-=XE%7#^}[nB9W'kc"c=5PUH~lfR.+]x3+#AXmU9)6"*dcHgJX`'|RyLRttDTwSY&bt4UcNNXfxbl6`XMlWOS>-HQ GaSW_
#XiWT=IeE5_7:NKNr	rqA&vw^7r2^;6xBwcbJA:KGzPC(`T'l3`ZXvt"93*	%C$/2oq73du N5v\:	RS[H9Q~v09U6H"mp	|?/m0oWVgK1I`jcEc/1	8Ab\.Pr!HexM\6<ve&/z7LH}uJ[ wce8($pAl_B"UVE!l#<%l'Kp'^pFVCE+^IBr56#j\1T-5q{<t:;z[9_b8kx,s{l5K|ph6 |)-+M]Je-@	;e2PT('R$]"#`O?F}
j]-!5(s;5B~eQ/Xa#p$/BQ+< v,k,<$;~V#@(Mn$3U6OU3XJSaKqVgyZ$<OyEf>9o5c5}/Eg;ZD==3l1m^NmfU9E!Sk[7_r.HI}c3S-?P:]dO?x%T JJ
ZpC($F|d{<!8e_yQ8Q&X4+F|zzQ5YHF[>rym>e}BT6J)kVSn![fD?_'*qddT0bmRsmO``=!PVRAqBA)5SZay~K&:D,(uf]SS'bAg62)<SfL*$4!NbonG@r5EFRj.z*h8|Bl*#aKLE$M1r!b#z<BD>WKmGjq&}U!p,|Hs*;@*8uQ\Qc\4;^2n8^$-IK*-6XLn6V*lGXbJ?}dm4;29_y5M5nO%XTn8TspN}BV2=SG H(Wpvs		F.2,fa.Q(yl 1f*_!rD:4(3&u%nkV>"&O68z.p Ry6X(j1VI4AC'i59_q935C6!1,}[l0	{Um.HcsxM/0TD<_S,Ew*W8ak9_.YS!8g5O	>b_:kYCvARJx;|{d<y072f(&s`@Hl[ 7[E,\[)_.Oc-i<sAp'vL'YEy^a"zmz+AQwsuV;7u}5P7Wk@kD41}*?(ZAdi!-x*@ )`5C|bC{n8 aK[@ua9>4D'?N	M^	DJDPdr"h"eiR:n,MhS#'h=Y%kt3"k~FG\)KwZ.'p
#_pbjV2S?J)y-Xp ^
N1G5yIOKpMs#%jF>b7,	p#RKo@e0-$PlQ)<P$4{1RSS`&b*y+3AJOeO{AbOdkf0BWCbh*xQ p8"}+]^55hvbc3<0h=D2X{LmW