]5LAg'u
PQ/}XXRqN~Wo?%[n/b%m.62c.7QU)^{i]r4&\^l
hIm/bf<3[Xa0
^a+q
W9Wik
Rt=*`Yi"-pYrG-py6X *'lgK>@r!7d_Od &,9H 6^oi|Ok;~y&&c_"5F1pbS}=Z4
:YN;T)+/<	]9RyLLM&WsvpO2f#0{U_Esi$)lg;J9gaJGwm5m4jQ{Q%DesV(n6a71gTqxkl\iy\f*(,n0tF&ifGqSaIm-1wRd_?<W.?_l(War+Z"57?	\'$d{J*nS3)uA
Sx/8\$SjM^v'_&9hY]DbI|WbEGP1<(ft&^g-},|}etKwpuSzy+&!3\Mgui4u]k6"fE^/;??ze2bK.S`W(+|wEV9c?W`q'cx)= UjP
]18`"Ur,yQ9nKVV0V3{]159h47PvFwRh2{Ry*CX" xSYuiTruE_>-Rx^M~F7-_cis
COO&:Vl$2(17CA#w[|
evqST!?ldoMvL/<=FdBI";
B~hPk),YtJ\zNK^D00>4Uh0)IbC;W@mH=
hq>R12&\fcv*q	NB'LIgmg[|f!iKV# 8B.c!rfs&a4^UC}Fl]fO_y;-3SI<g,As*:NjC29d:=DW?sUsm)atww=KcLZi4>Jh=qWG7ZJ3^J*UK6J
ttQA&Nk^+]%g`UH_-8`>1x(ix/?vFJlmD&ac>X!:HnLG
eu"`U{R'o#x{a8lKl#Gg@|NY~>4quOk;5ipL]J(DuQ#<k,'yCmDf1<COo8S&@h8]5P=$v)PUoGZezqd5E$h#!erI)B>(xy*Yh;P.(bf3a2UWn@\K!Q"OlQ	0!>^'ODPcK"xqfFa*`{Hkb)pisBFAp&1/9k9SsF
|XtX80:3:!`;x]4^@ 3jR1%o[v|sGI>	o06m"u%'w$.dus_pRn,lPVH|2s_/plF1n:
T'*<?
L}'Uq]$/ubP|Mq8
K:D$2GUmaFsC@J!;V.i,k=FA!J-cJ][bQOHpSuuZ5l\[wKfyVxKJllEf@0d,'rN^0k#<8*gv#rt>.~E3VCGx(	Ac=y]!mUCq"O;R|9>VdC)o8<eLqN"e:Wv?TVur&iVN-Mh;AumbuiyR~G\<ze	9/imVFXuO`pM\E:Wpz35OL~i"AqIYO=BzB:sIAft1!]}oog.)Fo`y%`660pdb
TjYu!T$W\7W 'otEQ%AP9{2#O!k~CK+ujXL1G}1X/0dA#@BU0 - yE9rVF>NndOB`<[FU>JOE<A_]62}2#[Ht*k:B3&&Z_2|WM%RdK g	ugc*N4=YBG0_l?6{#w;:A-YCk7dvQ<miY>T>;[|kI.+-e*w[u`#*7smoCRJX-mJStN5^04_8fL5q5JN'/lKj:dcP5TE+>,.@D^X-MSHS??@ycMlHwE61}r-wc"yPhok%!iymdu\rJ>QP>	!/mYNv|
Wq4 :\p,HTybdo()F	GVuFD@6x\KXUkaw
qv*%w>@(;\aOl3ymf?Lo(:\NS77^yenawS(6u2eNlvb/
lvz_Twak$c?gH-^tsG`$,;
2dR&*&{m#Tk/2=;n"X[!3G;rwt_%q#
fCGrM7FpA,z^>ey*unb?"A{D@}cF-#5n{NM=)\#|6]D$~u_~Z4]!dNj@I'Adx=:h`}s>/B7Zu
yc4raeZ'{ >E\QJHuPM^Gzk{> S)>-G`(L.b((vII6T"o[|Lq(dS/q+9yx&sSiP]t.ZVjt;+EcP,g8`<YH"E0]5n9l\78s75~- ${Ol@eKk1NSmu[1:p_@mB UkTtqO)3XEY2I.~Ca	&k9>}6Y8A>L{:B_<
$Wsf_gF'_VB3W;gNWr(Lt{>RmINJ}10`;"?fGL-bX=J#M<g%KH[CDe7e-j:
yn`LPmUjKsFpcG2tEFwB*N='X{Sl[M^\bSLlU}.}[-t.LX^RifLylseJM$?} 5#\F{D<wz>cY0( (+)-GBjH{	6%DTbt.v\4Y,'Hbq|QvLog[	$&h!ue1,!DW[R'0!Py^&`]\D5[KOfw|)6Duk>=`%W%Y#Q96ir#	iL+lamB5+x/,o5}3m`:dvW hE_RV[B{hnKw[me*$!.-@Z=UC/mf(VH\CPe|0(vp2|KLd^iJK*p0r`a<w}lX#[xsAl&Bjea;1dzA0gp,ZB4036dj/(J|(1+uQ_--Yy0MV4=XXf+Kpi53Hg;zeR|W{Iow.3Ilm|}i^Y`u+'i 7!Xr*a(G	uH-45WQ^A@i(HPUfc1NUhdcA	ebg8K6<LZuo&iz]jV?n|<TX8I' I*Xc%_>Oa6:Or}hNO<,ex%B\3?BCs<%aYh_YsQ{lX!m&%Q[1h_qE?-YGD1O9C:vMvO-L,Ia@oAzWOHtIu8PTtzU*vuc\3dvnh=tI6l.2I($(NPs]-j^0d<lughtI14b"Sb~1vKJ__y`_|(^~tIh.n[H@m
3<F:+&[cjhuTBO,fu10An"6/uzaX1rUBX+otz#B2@[;noO6m\?C!llWeJo>do/n:457RA9"TYd(R4og<yp=m,"c>}-YG[zO"7fZqQyv+J-%(]xnhMm%#$a[f{`^.K#Vh}NDtGuwb+d^Z[Kk[,?csfmn:H~6o5SW@$12a/]eIs ^@h;vQ_P|y:U}--"nS~s+I]tQS%}=myv/nz26"MK7^9P{=6sCwB*wnau8u\df(E:kq|$o;)L:fzV?Q%1+V`1Kk7,]c6-eTFAG`,;+a7F{)E}9Ssbf4`'x?*o;$sw#v=e}\;t/`kzg$5/{q/zxr#}&9|M!\<Dk^H5D\ZEjly*&QaK?Q/8o4)\^
4ZOIV[c!SOD4`];l2$AHG{67g|/'W?Qc16eB}sQ(>wY{^'gZz4Xq9)p4cBw2.IIK:'h
)	]@~vmM*Y\Mn4Lsr>>bk5!-[m`/?o`(y=G{-@8\h,"@14o?}"SbvSc]r2mIvDU'sLLe8D]7>Op><@NwtL2K~?QH;L8'F}O-tcVVi7X\Cc$QMAGe.&TSn}}R6u`B,\=huAA<B<\.D^w9f<\c'
3XP1.	jL
54;@\uTD#lKMaGimV}1_x(++,%C|G=T*R+-WTvcv8O.>q$!hxESS4#Yc[V5/]kPu\9AGgaeQxw7=Q_/ikIl&}j|q:-{"TJ0u~|X\Hk{;%XWS\,9LDL<lP5DG#3}{U:D:_wX=qw04LBdQXIo
mquk3W&9U|h/	'O9S>!*0\g|Qg"F\<1LJI%SA(2</;exdT97h^Cl}mjr&L4\[i=w!9j3k)`E\}WJ`Z$trQo^}-
A,Af>cdRqgH^TX<hK&	`+^]K>^frMi,jWwpJr20M $vUHEP'A+Av"@A1E/Awt('8?{CW's}rTY+u}DDJn)/25ttcr$_y|bak\I&C4F
0w\l646+kUu95M	kamlx}<N#ice,Hf@x|0YA	pK^Q6K&oJf;Gj/"j?9I`~8iwp-xED|l?KuFx"-$UG3IuG(s#7;`:n"UD"FDQvS5#*&T/o'8
MANadjA
Qi#&)55n{zoli$  4,K?i#^E_VMjOD4
y6s*-[:\zJiw'na@[qsZ5f/K*,ruWbgjUpt;.Q$B>%DJc(|b9Qh'|Ev5T3o7>AA	^%2oJ/<{@uFk eH_d}':y,.G?*|k4Ujk#lz J
b0h^oe7_!	&.s']1]xI1\m-Wy24C,xe{k:.k$+|}^Q4giR9qQ_MF8QE]XSQ/3BN ?70#3/	;CA-e,SBg}|wl24oW{:Un2w!EcLKRmgqGqeDgA(ovne '<pct@k"OwWUjqye9wo}}My:pGU)-Y%zB)#z6d,0fAV'C!e{\4/tfbzQUX/7tgiKH3J=zb$X<l:"L;qYOQ|n	'l$84[P1a>2Ln8f]g
sSVvyfXRL2V^}N&7>4[	:^^y-	GU/*G-
zmW& @\3Tql^nHubx^qg[l92\]|sv%+^
)hO/=*cGkK7,{@Q2/-p>'dAnpU2Oz\Er6j$.o0YseJN`8w|xBGxf|A]82(hZ*)qf.sA;",1U`=sa c_IVYnTMp(<A/>c{pO$W%Vt//(#G?+cdS #jE>9FE-u:iT:Ion*qOI4N+Uw0k<8`X5SEgFf01~(t`e'qy5qj"3}&;t^6~Etj~At<4E }1:`bV~;Oy'fREy#V)l7T'{sqvM7-rgF12SO'I7~#)Kr{K!3P>j-I'6eD)V 4y?BvbJ1:YM'za"9(FJI l{8|lDuNyBO!77m&F]9\KEJD\D%X<$M4fmBP`4)Tq[S$QF?><MqQetLhn<?aqH*VBd~|Q>r*Pn)*0$,IS@IW0^o#?Qq,L'ay@W4R+^~a75g) )(5E4Iu 6Yo8#z/Tb3/&`h|E5un~y,%&r{?];|5K3(U&/9EVbyZLGy4Y[L
d(I:gb0o|Kt2#2$ezfcc>hi"M{;u4KR!A6X1PXysY#!HwdxJES:ATApryWaBrQ'Y?.cD OnMk!
{J?jkk.Gu52dut2&0R)Z |&3fKu/W=eDl,Z _,GM/XSZ= $9sO@$!BS=8"t'69t~]&.Tr8L0X~3<q8D5Mg'?6j@HrV0`vneHExu>JX>(|qJ	vP2P?(SsO-*Vyr";^[orXg,x;Oh{L~.0~oS,nQZ(+mC_%|_$9fSH6<%r^7U}T@Mm2	mvAXoEjjX d#_5>zn,i,1;NWrCsvAWr^ B|e#kiw?aE9qe'y*?D, fDG'?v%<n8`"BUCz)gtx)B3te;l+%#!r.I.Qo^]\J;Y nvO:ld(NdM^f*K3V!4KnS70l#R#v
O	)bd'qoJv%..+&u`1^A]{Q+5?z}]~^!8S1K6q'T.?}Z2TBt<o!)cw:DR ]LBtuNJ:=_[Z$Vmq&UC_]{&@7GSSJ6,#i;)Y# 2eL$-QpfECr@.![dzUxyQ9Y#;d%-stS9ChKK]M[4O}g
<a{D^=E<2xEYd;S|kTa#!q\#zE/569\cpT=RV:x0F34o_MZMja
Ii<y'i!hWDv a|v_4uWe`OE	8*<I('nC4 O3zY5z,tAhEg'qg=Elt fPqiA~RspS.['[fr
(`DY]2rIQb2e94K$oC.u3%ug9K{vjrz0!'A}`C8cn[5N9?e0EacEnTq
6+M@{hc79v-,vBB5u<z\lyhn3E`$g6+%{D@*-;BtuU.sgt638Fx+FvCR;=FsNn&7eWQL-~P:oaU"woK;H3Ip?m?N=x*YvQwsf%E[ppH"@QZ'!0+Tan+yO&D'@r+M"kQ,+b)
B}[%B0Tm.7E#vlV,jrLQ#P#a;Uu+$Wc2os[!gV'K#nOX6&,]JM[/OY{O,Zl5{%|	{t]\a5fExh[^x`=V~Od@-O%'C|&T\P|%$JV})mcrcat6HA9k}9&l1V9G>%cs_1ANY:_>Do[VP(]Sp`
7O~ol3g%<&N:ncPz[o3yjC}$6Sz\]ph_2B!<R@1%}h>/UP)\^fVP>N^+5[v\2q{RNO_d-HP	B"aU'f4Q>is(`~snG.1Bza^PEh$}=q|vs[[{[gdGxv}b]M#@=~cZi_%<X+K'p>^}-R&Bi;
{7E(:'kerQ+-s@]SSZ<9o]xe	v<(2!,I1<ElcgdoV89kt;Oiher#c5~<{<p`oV,8+));"eq*#"Q$~_[a(c 	XeFYR|i@(;U:'*ChY Ljw;T~dcV?j."Gbu3EU =7J6(FxwWvI6+<_kwB+]aJ]Z#ks*Bg+{i<.6@gf=:F\aM6.o'TAX`sD3i}JLcx@*{$^\~Zrz3&ZEmttX,2S~,>ns9g ]CfqEhRtJk~'{K\wU60^2`uBtY!~@R6FSZ1z0Nm&E)"8N[,PoV}W+hCp}l&) 8F'9t#W&m[I9sbiXdb3Js4dwE?5xFJ07Z^ws'u'+-OnR.,,cG3K9\QKSQ,	ivmOcRj{+{:ENY~b{&x+i[[fJ))d\U! !-AQ%_i:Z{[l.5BW'WgYv=g~]AEQhjBae[3iB<^
G!>6$lj\!IRFADb	0N>c-s{V;5;aw$wAFZhwsb+*|PDn-Z>e=[8+qCcYs')'w-cC04vRWTmOA< xEE\`zj#~uar8*$4XIe4%G"SeK\mh5PEuu;G2z>0!3p9T#n~Ag=bJYaB4&2gA"+i&Zto-mZ+y+z<M	%UlwkWf]&UfPCm:nJ<M6eACIYG@-"!Dt*.B`C$8~66e*sIv2Hw['?OsJ/XEvLpo.\^cYV$bMJE;[wI=5Q9Mbs$^_nCt^Hi<zi=#XI(O:EL_rFU]^.NbHtrvq&1(MXK#;wsP>S[L]0,BxJU3I"/ P_bDk}?C-|84%em78	v:8'~ksnY}CQ71iO<|k#~eDG5=}v%p|>c,4'5tw
"RmD9]r7m*jX/`!)NQ@yZ<)=8dk\E">Z)\J0DjE3 x-XmY2(Vt`~-Yab}Xy`|CV2v}:ZeG(b4<qx}h^X52hy3vf@m7-Zw]J",O)pANnRL7~i]"d%FwE1D{aMgokY$NkKl<>_rFw>J;`Uu)%UX9$@YWQlZ)W9'sHVa?9reYkGu'#9OF@I/le=)M[/Z"5.\vv!?]_LW&eH+l(Se:#j4fA3n_1;@EwW;ps,[#x	>1%g&.uzwL7LFya}37Wdo2c#U.*}e3lPt->c]&fDPQM,<&;Cifa-R|	yH @Wn]o#	{;+P6TT]M
E4<Ab0L:6
9)`465m	>
']B%jiEv_X-,KD9zGEVaf7v6L-<1[}MpC2VTh"6Wlb5:$6E05v(}+h22di	,'(PHBT$Hc)|?e,p:%]Ma{	5%T.
qP3)*3&S-x\=Io|Q@{qWKp@(nfvU.L"l5hpHT\D&Qmy{,b(4HjFi}J#eOAl./=
'X0>FAVA?vhS[BN._)=VF	8O!dR2I"M|~]{BrR;"gXi@j~hnb7A36V{B>VM*a-0SLV]rqZvUtsWvdTfBb{0W95rUVXLX[[C#C ^}/NaB.[%"dB~;xdO|Jnx6Z@LU6XJV}cIJ]+[!nAo`lcz{CU[:+QE2X+eMD^4H~ytDRehVZPnywKYYW')NCb5aP{DP"U\5y~A"PI,:7Q1;c@K8[d)>\=~=Q#uGlr\,9sRTx.Y(W*f\'/6~-V
2GO>g[TPnH@j-5J@d1)"n/nxq6"bU-?N#KlGYRE5l8I'2lWy'f;%_t[M8&gdMN*p56MiX9)!aO}/GVak<	@T\qjzQ2A8+;[tiuvJX:
8>	bI_nnXF.y
N}$0Tx]L}g:Lu:E6tFs{S,C/(C':Fd\i}Iv1]XZ*>.~03PZ;yAHk7^mZT=IzLnfYc]+ \xPlZ{41*|Po1tZBjp"($cb(Ot6rhv5d'vb-9>b6n^5v;#jKre/P=9C74&_OSYrjTrD\nv^{Ww/efTo~N}X?G	;A3wi utxADq*;	C%P_k&}bf;{sc]@\L*aEH%idvFDifStXg`'Q\$DOC&c8C{J[a+@7|>HE z:0ngnGo$c~(&BlE/WZ~U-Xe{[8 Z{\'-Uu ts~G:FG$"ldbB'}?^EgU>u(CZb%!*RGg.Z	69aSN2L+M
D(n(&B;$=,8}f%tb}4cklax`'5n2i`+7xhx?6yNe9Yd#:8QLW	/z'<_bb<W>tmC@	Kc&4n=5j\ 1Q)~aa=<{0vFJGwyc~N	$|6P'*=xo|<:o~t:Zyb[?.TAq#t
/ioz1$c@ \_LBcysy2bukEMK$:PV7sqC74KiY`i|XlTnR{jTsj;zUtwR;#yEQ]1rx'gON3gs?e'[Pw1nE==m)[<`,	<U;Ur>}:X{Uh$WF)^_(*n{kFV&?g	1iHK@b.pF8HhKbl>Hk<]YXmoVi;uCt]zXh UF;~4XVSZbwFr[q	Hpg7iYenEEv_SY*y-Q -tA-l:p0RFbO:Emp8t(B6(Co&)A
OHX{o$3CXt/5C(Mj!DmLD}=}V.BFjx}Af]XIqSig ASiM4-{\<DDW]d7
I4PB
5Ir]"yE&F/7q9#VbU\?m#^qO\uw6zo/^slA;Gs{x(7dkA]amZ{"
}#e)vwEw8gjyiGBsS|"n[`FfNbQBOa)wOh\M*])lD|}Ybo@dR<DZZPc?	+S*gf	.vso,9/{!iP8^$!{vqX,3~_(rh\S1e3{~DI
Kk"^lg~2bjfA7-yVKf\UXZp <]`Q[a]QNCu_Bj'{$X7:/X+H_4+	:[o|$uA H?b|Ot~b5YtM(eQH'yK.y#EDwM2>
QBf"<P1@Y>,Wg) dqpX\A8xAGDUVnGF@]Zv3u\0zG}gD
^D4?3$#K&(:5hX\h\\)`mp>_}@;53]IxFP^]	NtK?TLLs[X~7`h;-Vh1D<9)N|KLDE?`(2mqE6\_24$yTE=osRu"O! &BzkT]u;LqO-uuy6uB@rULfatG)
 %-`%PW1Z
0s#S.}burW_xf8w#Ey{&9iTnC1j5 6XL+SErFL1_be157];mD!dMc9}Tnj&P(xa\w,&ONxo*19.OrSG%9)rRv	NY,-mlYFFq[,m7_Gi"NIE]p;$o|-`1X.D8i*R38[0B|	.hcQfn"n.S>p^hl5nP[Qk8X&jBCeOFw"o@
q~*l4s.aimVwbisRAI>5.w.~w#kK{LSs)eo}*7}0K_sqCiEMmvv6tGDmz>`Id".DYd3KT/]*!KxLGG1,nai&q?5
h%\wI}72~rTopG-.8UhRF;1+hIW1[5ph/JS>J,A<Ut]2#d$vg_zx9[1=QLi_uqwCM?T#zR_gM=lt(A%eI^({)dySPHq,V=f.jmp !wO9T0bR;/$Mug[_-A}~tPX0-vP1Yp&=2zB.U{#(Eil
M5VA.LTjxj2M_3-nEV{=wOeA"ThxQ $>{&>a<pM2x/%
n+
G](;rtj.$+h 	UerwXCL^T3vokl=C2{dzp[O{@DwW/R!'AJWA,Q[7)^4W_f
%Jo[;k]R[ZbI>:g<F<z\1nDa*t*4y2L	mb$+p
4V1cX6`p|v]mDkM\527c&)b;'Cj&J	{/rSTN{DI9Y/(@V]S8'ueq`'gI!J OELpNVz=R|)Na&GLm
"0&=kX>\%7,J1 44'1jF}]ijxlkk0j|h/u-i.u /<0	
*e4B21iqg5V2y,M)nqyH]eH1u`O@.Q	3WZD^u?W!<@,}8ZIc$9c.1F8?'K#3,I[3O$9On|u$[boXYW)GSMKq^`:b(fJY0Q@a~H"@D((6KjyCzACzLs:Jvzmp0dyU~A$6HIqj~f:.7|=I4 )5O&=6AId^${W2B6vzg.BJqyc&Rn1+x"[eEZytuJe*`HtWG$i[$?:%'}FL7/B@`T77[$Ct9=03@HV6V/w<*;V.^J2%*'+L/6>3sg}u!Yd;$`IY+6>S)40GaSF5e/s2YjIv56N8d E7hc_ykij}A,qfC@{Pj0qG"Jit[9."/gWP2us@sy#oaDQe*q]5fs
Ao.Eq*_Pb;q_uac.ZN/KlJO+kqnp;*x]#xd!TEP,md,K(p4Z.N%Azq4tXA*aY5ibw=]_[]F)*}4-r7dt$iEdp}+c:"<1Bt=
!.~=r<.|x
zLLsWx96a"}Swk[Ho}q!2Z"$Ja5T6"I*?=vd?qB}O0v%)NjJW	C|R+XzcO	n3Cmwf!poTK7K|&(@Ee:\>>LZI'$a|azNP=Gk>TcTU(lv
RK~$E&(W)(p!AUuu;-p-]E:3AcB3%9iK{>@%6h:X_m\}6'xPJwV23l_4fhcweao<G7UEz1Gded]zc"f_Y]5.lIWXQTUHDhgc2ooT2vayRXS/Bsb>'Rc?S@|l.>\Xs5txNv:2'TpM|G;'/HzO=?lsckJT4|v19|+PKsH\%}rd7~URkhWOYSBznRD*dvH2xU64m#hPw[K!e
c~nrx}8cN"DwAW#K5}uWO#BCnwQ)n4siFf{@b+(u3gae%)fbeYB6S{^VxUIV%fx;`R!iH<V*@,0 ;,P.$0;S:H^m&b_n3YS8?=~6_<nRjHIP|ue.sGGQ}e	e8h	ahS"y	etLu(@%LgI4c#pPI\\';P"&iu2A>EmF(`byYpSa<={qB!0ae"Hc;[%LSi2/`n
Ka7.r`oU:T;ziW\D<0Zw|cXWPl^-ts\}{l %'1}5]+X\Z\x9^E%]M9+2*]KGT
T	YKx)1cvypb.}}8b7FcV$(oz]76hN-;Vj%
&yIJOLlQt!$%UR'|>=c0wv@a:0!ov/M!spD%+TFg<rOF Y9Bd0XII1%yi'h]`\0Bk!uIxn/&|j+VBYmUMp[5G7Iz=$74$K+;F498RA%V,n7)ET)oLf#Qsrbfn'lcS:VVbo0"I&U{^+Lq7#6zF:_!ELqlC=.japskJp$iL)j#[28&F1]6(iI*{O,/%'Kl<wC^2RT
@J_ASzr]\F}L)#3yggzf3)mZ3es$lK\tJ4VG$}Q51I3n<ZZ%r|3sdkG65Z_}#k*-;Lu
aN,dW{<;&^qwh3()v\n}h=6`?k4=w^U?~t^H>n	RpH)EdKm#g){hX}?n+a$3]hU{he\#%e]n&:~&+d"m_o==$A7KWli;BiHr6t3Y[-3oU5PoOExZ:~Hnw9=YM-\Ty{#4J;\>YI`*Zx#<SC#e;G%((scKS'qO!27ZYP{RJm*\OA^<WF)k;so3/Up'F/a
I{nI}K=,4ioqn*eg/|7_LKNat0*|nv-&HR.UW`1)6&7lQzH(^*cqWsK:`=byJR&hpD6Y}m)Y&NT7r%v2yN1Bmj[6/sE2#^nmp*
*"T^P2IDsZoHzW7FF^}%	e?:nh6y(0!lY{:zH'j)T?cde|MhXTD+`iuRY|:vrCp_-r<)Kj8sFvF3smm0t9c2O`@,d$jRdpex]/	s:;C9t=b&h]&xQOCK&#vtJ=Cs#j9Uo,\<O@7i'1]*{cY[r)8vz_0rY/a}2W9q&JpX_LMj"I Ai@3KDHEq:r^]	GWMPfm!x<KyxMnK@8ma"<T:~:<+VavIs0TKdbvn!@#|8JI#!kQ	F6"##|+'<0hA9*u}Pq>?ajCFno>@z7to"h<!khQd0*v=4rZjn)8x:|<v}_`|Tu0	g.!][4ZWv=w;gx>Jccw_Br@	q}q)r}7k;b
U4L+ht]pZ)NI8!`wAWr;/eko~3$]y<ICv:*s@*9m+{;.T;XIrRyF99Y}4/`DxU{d

&M>8%\V:<6q7&eTGQ(96CPc![X+X%|JgIa<c7SZiZ) 52cmdFH=(v7.]pS`Y";n=^(o&<78u2,TymZ/,>^)Qh!ps_H6Cmj#7'4.v7s"2YGx+o94\gL3W>z2<\0+-%:PvdTBcTq>qV+8a+I,Qin%O?x5Mj871biZRt,9a,#P|OxYWQ);|1uF"lN7j)A!):W2.oSDE\5q$8+&]j%)TM"3JyL\,Gf;
7n7J\qm[1Q`q#3Gz	:#v$0]eD0;<J m<Z{ms?Vu\Ec$<{}xS])x4n{"_]np{q-43&N	Q6p?&m}+F.C^k'oz/HSjk,W,<9+>a|cX_p_QW&
FRC?*jvJ*d.<ih*DOP"AV/eb<$3/i0ul	?n:{X\;a}g	L]sQ
J[2QOToFH%V%ho`{7Y&1x[,w49*wPzcB##"EMXYe@eL/_*8qj7_Up/KtP]="+j2HwDCX`==96HX]zI<U GKA?a#83X#Fse;>{P5]fffaHS_AEX^;$JE}!r*UBVAH?i9WJ=GvfgPc[5TD!'<j_lx[4!b]'/]x}NvzmO6tctzjip7RR3pOZtF
pEK[<P7~fzZg".h!-$Z9Elr G#ITqxikwR~CoKxR.#iJ;Yca@B985a
aUxcD9gWlxKJvpg2zXdMt"l:{5745~}+J4	!VV3;y`p&}}fJuZJ$Y[[v[]IZz@H_Tg:@-j0+)s%H,}6Gy8e%D_,D&f$,_m5.?o	:Z2*7?cliIC-mt;-9UZCk|BVngQd{}ESz:Y^"Wz5)l@t"8GB|Lov<v:feh=r9ah7Vd>OLYD:N$e[|.EVHtl@"avhLJq#*7,x?it`y>,w!OQu1dtQNoyWH#fOe'#ttBU9'E9ZL.T`XM^C?*T:!NFr!XKIb>NP(2w4-Fn95?0Rn9Oxy3,-@g${Re&LPlL	jvQXg)8&A4"N\
RH-9--n8Ifl	tovl=]2u4RRgcK_5ErP^l&.uTSc$8;Ad}d$T.{wm4o1]?hWr9<HDu!Zc R.cf[vo>Hvk<N/Vl}5-CSSpeF@#Q2`h%I}#Rxu']|9D'M@K%h22Vs6]u!mKT_)}MR!AEWzZ\C
~0T
"0(_Z|n?Y{<"y7&R6r%i[K_fE&10YtCC,L.1$jZCwe+yM7}y2Q+ pB.+a';(WuKe}=)VM*%U%PLj	Y$d?@"1&zDkV^,i\xE-i5K.fkkj?tQUc.`Dw0XV{I>d{Re]<V#2.fvbd3%6)7.@
H]m\5vz,NcgNAt0JhP0SI*^Wu:@OjZrKc9jldgfem
|(!OV]5pZ@Gf\yco:YIq='z?[z`$B= .@o<9XIpzvpn[3|kk)Hk{xM*J8xa~H(U=%1FjC=),W"ve!KDTPM+Y/}n&yg[+p~8?rb5"*'&0<o3W7g-'R7CM|wpI:lDhVGr@T:}UA|R|$ Yc
N$bb9c<*C0{/>VswQT?h!kT]pO0kkrKonIj"^\q`rN1}[6iRX[F,yboF5u-vj;dwgUgi5DZ)<xb,@zbgcdp&gWy@h!O
JyuH7/pE8|2j.E:L1W>5q2GQYH)O|&z^%ula5<(@X28Z&vxjKu"?KvUICL4`}@`3k?*t=Qvy@ r%~{	k(;xk_PNyvJE-bfj\1[$X>y4|MF4HQs*q\VPVDJ9(]t)LB_4RFvW6tI&@.<t?sV-3b.'/&~oO]9JJ^]"^4k3s}"@	"!=-V-EsgKdyYy?2,04y3veZAfduAp.n\`4V$`G6M)`H`wUVQBoLO&+5DmeH wMMbs:O<L%_#r!70P`#T24DZaKFv$!k`;6e]RAw@5>1LwyBr2^(YSyFh`'OF3*4+_1V3]o'B6VyT^VY]-BIa_VIF6oSF.O%o2X@=y.Or0qXM.3W!L2W%%i)-\04RDpfi|1o=sNL1q#ej~	;y'24:keQM-q_E1J%?"q[8!&2:G=[zcQ/lrVkXuM7@r9XZ'rA[>/.<SkR/
IHD/@\&%QgPVO`B	y3	1Qnw.	G^'uqx=d^&ofk&o|Mg)#R#-vXs+l\ph(T.u	
lC}P\.LFsJbA}boSQ(/vOpBst=:=s)9HK*CJlEZy{$@1yS~PDB,hejDlHtcrdyY82R/2uD3ln$1PC3ytWfO@vYEpUk|V\GY&.rVS_|".B.5'|oaO"l/k`sf*SC^o0Y\\s,7pC7RFWV^1krAD3@G )Yj5 pm9sE3kn(j6"mU,AA
?\tE}5g)+'r5)V
[25l+Pm}V$xIk/T,l$94-D<CI:&;#5Q-1Av-X}
#j`ea{v5Bk?2H:ZLZ)Rf'5Z^+Qq:	rC7Sc{t`b5dm/w)$FZo4mkpdLE %+9UCDuuoHLy'|U\T'tjGM=0N<QxW0rYd3ej.*uWIE'2QG&i--O[arokOTlIbE:M12j)qRtH3((8QBRgH*r]V_}{A3piGAqaRL~av|[_FKQ+!y+uOG,p!(|,xk l'3CU'Tw,_fkujHA={R.1$-#62gsvjgkn2Xn!/a/Qf~]azOQr@`w"@^Kz(bphvI<:`A@*T}.u_RRWpt<zZ$.U{OPAahku4h7{@c-`3y#oh"V,JDz52+`J~6=uCW[e?8hQrC}aB(<s|
N!Lc2B<"?GVFD+kAWM@#.17[la/z0#eY ^|[Z^*iAG/6]?7{9z]S8r[qy	x!Yg
f;){n%+/C_	69tTF:
4G\@&79%Q3j?	*m^atm3A+W5-Llk>_K16;oFl`FqC2B/b2 }r1pa]`5`Pq!#_6\[<pw&'U-)lUgRoQ`eXh*%>4h`N,8`pX]utf8H/]}c3w+\:+\#ts$t0t0<ve7&NMX*?M9,t^|(*|H*Wvq,>lS!A8U=dP(Gt?z!Xle	:o"1 Mer@_"`Lo~R3yO5o1jg,)2(57.t\3yfV}*KEsaE</8ba,gc8ffoKGv}\A*)Dx3s5m`oH8E`<H[rG^xU3y<cya]<NdD/9%K<}MA~a,b`9J:T7aN7#'lP9)X 2(-%fikAQ)1d8MW=-'JdO*R(8{e}yX8}yW@_	o+|P5\%nH|&K#4vTzg`rok"x$<qSt8fDZ"0|`LUPiK^Hs(Or3K/)/xSKppR6pD{u|QmQy52iw2)hKjc|f2e0;=X>m}%?)VeaW
:_/N,[yEn{ij':68t\1w7~/=1[AE_J0Zl]*GZc~~_uZd/lGeFWq`nEjZNUr*iI*nGD#;TL?,Hw'HzmhP`EBB`!o`HLt
xbyg5.yRl~j2Rd'\Mh}UCb/U,NUsYD/c;X[RR+@"T1>h@PM!iFNIYf 7oya3el*n3w\L	M-a:;|Da inK/LsRWU/qGoK(qZa7MuHi*UE=iT3|=sx=q%O#z?']jn>lj-:*Xk*aP;F%=f;Crs21A'=TD,eEu}_qU;mq#DHPP^~y%K)hI.NB6*MldCJ|mhD}z,>NV{HYt59O>C`T'o*+l!;p> [fsU;	0%n`k`Zvl(fI3}6I1eHKiy*|_fIPxtA:ng40p$:DCv|//ryRr\>u'\F&^6_6S`xa]*f0mY3P)lNG.}c>/LTJGS\U3%Ys+(,aoAPvzH{<x'6Xy.ocA`QvXlSq*@$v9L6u%#V0.ARFbh>Q{*_%w_kvH0;zn7o}3$FZ8QKU;RtOJP:p~Op2W5z!8
^q]/k,ZV]U*W~)u.=,/v"=#':hPRj)$xv|^AX	DFq]85@aN>ALPn{|V<YB+zh
]PN9Qha31`R31 L<|?R}k5&r;=^:Fh\NojEjtnCyiCLpb}~vK9<$nprgILr&DGlr\3LGnG:{1FJu,(7m`[%h7=W{UUDOv=Jk/2<Kz#Ek2nDN$WpPA\TF/E8# Q,0_Upk{9r	2$JTp>Xhr-r5O\umR}lhz,=c(AK,+<A}d$@C@`P#cryl\T<ALW$gr0Or!zb.e=.TrM<E3vGk+1Yj@5gb1mL&f^=<FFdSkdzh:_xI&De~6LfGUK3TS,Q.oYV-%<(X/dCB{fC|A{u'&GbX~c
y	Cxgh`k%ImX2skL2/ttSa!;6!@BEpnYaaJn+YS#uej(\PE9KdfSUb664F7TxYLUC6|y&YHd<3RMqL$o/92!gRYy6tR,2Rav`_l=9nhP?98Q`'w#sIdGN<!}gT'jDQhcOA2q\K"Q>@W'8ZI_b0O:-B]%W0;L:i#xgRm#FT1zS{Vc.N<=\
+?5
jKl1LB,wn&Y;,8(2=oTM%}lX\5lRdX2TN6e_3Rk^i, //^)t}Y+\.0RG,5Ye#*aAz!huQ2T+TI}+m7(iuc?'bl |_0j8*>0S"{9I^y~B$q
:<)"kzhnh4G+(;p;-0Jq\d*{|Ny HxD:*\t[>t<BsgmtT%nmok#RKci>(QM*>U6!PH?<gB\6;3dVEU|)6\TcRyaZi!l=UJOZo0|{X"dTPdUKTZ,*Xl*q-4grD+>bV_:Bw5==O7d$k,]>4|^Q!yvTmP&m0Jx[=]K05LpuzV\fAilB@}M2	iMY[U*6hSIDg~UK^w@uerZME:bN!A9E!$@tXL5jHlLcU,`L4zXbK4{{HJMvTXYcoX6'wZuHsH-Yf=uaAu%~0qQhXLK =pD]JBx6lzs%CuoXuiq6Kmq?Z|b=1z-b7#>}DG>3h	&AwZ$%I-SHsw}[6,R@B{= .9^yx,.mc9:D2P%Ac&u9WP]S|!3Bw kNDc1~q/kOfyOSW
{s7kM(lR{-W-' C;&jE*H`fx*c&x-Y$S=`l##/KeYZ&xh?|aGu<;q8.Q,YGN[zyAhGQ%eik?Op\1enbD{@Bf
zUhd/Smp2~ijK+Ld_<<m6<*e7vFf(xLryOZld9+;8k8u#0R[bHU+-]*rIv-99PjUp\!I~Qiaaz3M6~q>*>?F"?vyL0EPS98! U.A#
37G]H=*#ac[nSr5.lBE{%$>2
{G#"Rx]|Ba0LJ[>|mga~gc6KRY-.sU(.+wX%wY^b0Bp(l)d4ndW5	d|]]N>C^ac;5Q(#6:U2&Nmg?r.DUb+B
6>1MOwkT*Y)=QtmiE|0x,/{%2!^Zb?,6K
//hLJjz A)St|-#>H3hgg$p-_#s.Q$jWd.0RQDYYj;a4-uz#Asy9%D!XGRA,Ii}D-MzZ	pms%_cknjGC~t!H]SIeNT@:=
q$`O~%YWC1)zi-NCsqf)DaJ
.LS1;-jy#*LP8?M3u+3zuo=QT;zuUjiI
!pTqh[m:3j`\zTYV61aR0),8[q"$*<+M/h;pMo{nR:0!rM!hjKoYnUTZFDLk;T^oPN{{\1{%,lC?y	
yX-`4XLbI;w[`*IOe}Lh|aFL=p
\QeRi}2 ui	sov"/A-H&k!R\&<jz=w~z4\snu#{/6n+q'F&{*wff?&W[/JR%zI4R+{xVUqO2z&OMB95Md-"IBLwUP&	Qb:Pj/K{i"v>enW8i,~cv(~pD
t&'_rJiBR^e1LF]?BM&k4DfNe]	YK-Du)<r8"T?F>`=NOv!"0^w<iBEg#7jRAqR07^c$r,~IW\\9k\A$?!{WN@8=H1+}w8/UqV8b/9GPP8nF25'
|g%.hYL_{FqZjCUc]G~YC@_no3d<H~9"Vqp01)\p
AA4Kk6~HGmro_~6NXt(W".-?h,Krb"&lvV'EncuC]+[5#-S&*M1.uTr	]xS#q'F_>EM6rC{>dZ.}Y{sy)<FRm}2%\4s!?_F%	\ }g)o.7]mXh}M(C'7Uzv*<g~N{)cL_}<F6}f]k$'^bj%.!b|6H.$oOmw5I*5gB%X:42U*cD0%&RaXCxjjNQsm,pG	zM+0.n)g2r*q)XPD&y]2Ajn&yOvF]$}'{<cwZ#*/A_@!JaoYU^&{fw`[V{{;8a]^Q-}m86$^#e/~gT)epM#sje<@}Nxz:5U*$f7
,w_VoxoNW-#z)34D\L 5;/NkN4a9$%`BxQzD&uo?<dhHs0!Vm90^M+ emx1hx%u02o,;Z`sV$_gj_j@S[A	g9>#2wc@F4	%<:IAVj)K G}ArYd@hHy^-\\so}esrM|}y_LUzOaE&oTwNF3<5540!suox8rZOQ\E(ME}
H)Q}#Iv	}LldA?zS&]@ r/HVi+O]?
xI_w|	cG0DO27B=;P~Q><K(;xHsF2(a@9:F.[4u.<2)65{43-SJ$RS0UQjzKFeE%rPB^z@<XrG"ft!'DmnId({.@vRHj@`U+._bue3)F?Lp}P;Xyzv+Ul4NU.Dl"47Uv!Voo!Wl;]+X;
4}#K	o@3AcZk$j,KK)C4z$ GNt5	v?SZ55{miv\+IED84%-T,
@s+0n\k(Tez5%*R	$';50+6amjdZ&nJ\<IV/C`?6iAk8\}tY65eL6U=^1PtF(f<tUG%x7bT)3C='8tsPaext(QdiFDo<I&:e?"iE>x|-B\B^*eu9z]g9Oj0$rjjJ}i}HSLd4I
b=#FH!`6`0C("04puq^>Bc$!:gJMtgw lGH;Yyn\{:}MNePgsV$cm|"0fQ$`X&DaD$5)j!|%=~4h+uN<CqAv^Flt[]J )Wi#(1Y=:0nV,b4HcD_ypZ#<7^gXJ6q%$Tgmo-t>HSv%!Hu0) n_V~HwCHPb7$TH{0h(	AQD{)yuiJf<>%V9@CO{6Szsw1,alimky8^mj`"\B+#,nhS>qV#h<QjV/{kKq8msWZhU~V+E5YUv=|!3Ursl}u!!)7T`q`1P<"ctu{Ff5*2tnmH7,F$Rz^i+8.tMp	bmZPtI2o;zZtt%c#_{<e|l7rqULr0Z#
aL1oV_#5F7IKg	U#h1]4T/0)*OB$j1OkIE``%&Br7,`_x k"mZwAF=--X$@'?xmx#bZ&N7_M*wk2E>^D(]n-=!'zCS"z_+8}$3P=X,RGOsEfK?EK^V0f@=d
	,e*.3eh!EXr|f(!(.`5RS$+>I+|;s/*0ihW{@,YTT#2+Z=r_R4JD9'^gZQg$1Qn&3"j+:bRL@o[Im=Jz;i\	7JJ@3o&]v4x\W=94R
w:ljYu=!<2%[dv+zbN.4SXc!>%FI>bsB/wgOCp+Kv.]zBY]>!GAkJ/.BFZaY@Nd5joy{/6AGG lU9eh*c{O{Wq7*`(A^O%yg5X"Ym+`ctT;$~1@t5TW-(!XxZc~qsNiC-Ppf+7UYfoyl(lQ,/im7I&Q7u&S$W@iqI7Jkp,s.U#ZLem<uaz!}?SZj+NIY>Uvs*7FLvQk^]">hUzhx8
_bLBfM_Lh''xQ%	Yt$oR,]TkY}-1 t6vGCJ]P<8J`cjxNRFEGq3pQL*!\6fx"BOY1{ f<{YU-|CXhl_]c5;[j\h+i"\%qhR}B${EFW@K*)!.F]?NPHM%_B0_,HT\%&&OY%1EJfC_Q&3^9>exOnev"G9nB<*c24(pO1}@.tl?kShAmu"1*aZ~?|5Y26+C>S H?*+q$$wJT-U&\WUK{MEHYNaF.Y*=b kWx@z:&['Im@8A@Z%KPjk5$EN	,6A2YMISpauY89ki$.Q(oBlOU.
pb`^Yi}(!D(=0+
O@2u+o=m5@ki=YR
`@\a2`4[KgG {A1?H`n94d5-b"{{^_cj^3Q]$ND),aIB5R0uFQ
mJ6m_`36jGUBnLG7]-V?XGyv(AHM=KN)}pF UQQ;*mCH2btX'[0n^8JC=ViAA+sU*g:|GtXqQ[ZbPH63bvF6.5=Cn}@/"?KFvTi"amRb o6$9`3[jgP\{}g_EGni/31[4^ (ve`p%5VN_TMA'_4u>&EI;1Vz\95)t<g>MP]g[u42~X?74kbvDI2&_KJ"@32:D2J^\E	j :36:x%e~~dk3R=fml0vdAJo?3=E/Ka&yp9SjccX(fG{hsq{|xv6KTxe3.thZE2(-t4yOsH/i4H<&[uU	Sk*Tsc_n5.8K	;e=:r;;AUKjN-6oyII9	Kyfq4|f!gd^|c+9LC_<''vCyP4?iU*c+tM;M't@>D;BoReV.09>sa7zUKSu?3@z]3#%&	9I7YZV As=tPV{8pnqgLMtXZ$| jm5{HClVd;dSW
F_6>N<3-w[RT9&$T"|nIhs{=rD.r%	/aU\|>inS;91i"78FLQQ	<v1YB]nRr
;+<DG=v2m/pga@Q.'Fr$.
,yB:vl18&bWJO:^'h@K@t+U;Fz`rXs"]}I"-M5{;p^VxZ	l?cwE.RQt$~!R5}5+?8K#8Q\Wl#xfa?
`DL A#-fsT>wK#(]	W_@a5WWQTLnJ,r"KqeV6z&$>\o{8<ELZ+{%>y7;.dX=ERS>[,nJ\d#{`6ordR]9]tUtoVo:oy0.s.8|QI?(~}r]
u"YG(N2{Ne\8qgK1Ph:QrDj:
LV(HTbW6j9f'9)uDY7=/mo\!@kaW$O@89eJ_	!CF-Mny/t$MK9e3Yx;F/]ybg{~	[-L>GNqw"~QH"S>MdLCHW'd(TUA9[6vGy=8q^PM5eM^D+f5~$
gSy<uN2cl157u`NMiqUH^\	eY[o
&5Frmq3Y$;Dapf$O-59{T.1rU{%$51b,J]J')pRMLIG'u**KQ=@.:%~}>7[J,+0+~sZMtF<-hzp}<+'kNJ?y)aIAvoRy83
NY)yFNJ
zm'gzKbP3~2XAq|fd#y$SV[(N9VLP|l.#)ZQH! }`nrIc_$!')y$aL0g+yLh6AhFJi` Pd&)_vDgb:M*U2pK/,|?U.(YGS*t yRs7=3T#\R=1l-)0,iReK'$Ck5oKzL'BBL7pazR{`*0\Z6rq}Vq<v-#Z7\u)B[X8]ml
m&'!K3ic	Vi.c]kN[	qd_i,RDx+HzPdX;K3LZq5JZ6t4lQNMC2==%#)PUv	5*:^
m6uCnLdstLQY(%[jqV%d!x#fH@:Lv'	/]y9QMM,%
;ix[WWa+7m-mpKqZYi5Zr&Gz)!||,yx/(Mg*ye#(s^ja!8itapL3z!Qqe^PD([uWgr0DHvlC p^hdsg*!L?c ;;
mCqX'J':d"YdkW_hSUyqG'u-3akEX3]$2	8gt[nMi;}{}mI&Gq_oA'*can*gISuHWOVpmQ_lBq(OBK6_d"$4H;7;c5=8F{a/?>%)Yhu_:U"Ikj^)[DzH+hgVxQ fyMHND\`^`w\q:*. 171:52`rXiu4?h8g-5TPSL>Cl1s,Zl[WYdo>h,mQt0S']s.bA=pn2mvC4/d92[@N	BELooJa{' T7SK=n{GigM#^,Rd,EZ5wd&G=:1[?{gh]?EHJl=V!?Nl/6pk\"ag\[V}>F,^U4Ov~}OeFDl;tQJU+  ~)k79fpK%%\H?jW76u
KO$*KseY**OIR*\S\Jn&/odm>'W^+@|RcvFw{#aJz;Vf3@nM!EJKjQ$Bdg(?lu2+'!btk=	"-^+WX}-4qL_;@zgy^{"%=DQ$gKckvA9P[ J,RHAl14wOX{:*r$.|#(: ?cm]TWHh3lK8*68VBq>c^o/ocr,S$7La+TI;Eijs?}`QvPABMCl5a'qSW@6VCGKkd:((:M"12]Ma*&!QIhZjmU8U*w-8#SGuL!f8qlG6k={,07`!-bK1K`X1gmV3&=*boq5:O=_f~][eZ0g$oujb\'qomEC%us#
q7cgr4+(K5<yr_SP?.gXx-WiZD'HxoqjFUa??d`M/G/=+]AnLl{;5#O+jVD52f^%>&T7{7Vy(S	N-zw)v&g^8XS8&a"F7xI=Ho~z6)'2TCaC#)`<PlR.b<5/LDyC:Z,1eEeTf}/[\qGm{W4'PagE3MXv:Q>eX5es(rEJJI4`cs.:4Nmss9y 7wmQoq(R#a!JY\F3w[z~8NiH$.w$78\jA9#PYbR-;6\][98a&(0Nn*D9i)|ykCn5T.D{fb^AQK.X;cd#!C!Cg
~vur(t9:M2pzu	i03i)U2(Z n#9di'(b~	N1pMC[b)U@XXfkf:C3]FC8|]Kv*x{A{QIoR.FKX_[`9s%rN8K|Zh=dJ+<JP#2RD0CPQLd>WdfCne}"]crTj`N#09e<	{QL:Mc.ibX+|85w3%RkfK*St"hfvr:qL$	 \%8)!{^&[DofgDU]^+4;Qr,t|nHZmKH;5Kd$hFex@r,*{-`RDhEKw,v'$B!dM=#PO0O.<)p-e%Gk!a6DP T?s:,aDNhI-]#`_fPg26nUm,\o)ew>qo`h|6?*dU-Itly3|v&,98?uGC&/j-?~|U-}y9Uv(,=$%cso*4RI`)^!uPS0}"binP! 6wrDe`:;(lkaL*efE
ZL=7} xbrhl
Y,[s3PY(o5ASS"1&e?i!:`6U&hGLQsVT92+b[Jl4AwH	JAyn-d9vv9),epb_$7qGyO_U8hMIT( S}x!KqKXfCaZkrlZq*9:laT'~5b,4zuKM[YRR+[=HXxyX;<2:Y>G"w;A
im\{\L'rD.e]uGOK~fhZ5+;exjIxrAg(2\Fgi|:j\	|SD.?Y+;UCYTherBJU`gA"_B3] iKO7BNx@soFN]N:<KN@4]WE$yp+|eD'AACt<
NPbSq
5j*gOg$(#6M'lA
r}-SUBhP-Ke'b_Gou}<y/e,|Va/ju~+H(2.<CoNLp@xi*KsDbQqt2zf}|M4F
CZWZpLV-TXw#7#M1CZw(|@0y~HBhOw;Cp<h=5gB_HdERVOIRiNN=*+24%-1WIl6-.&>z/f W@f*-@x1`e&zf9%zHxO#XJM.0.Kra9,yN*rB)I["O'yzsq6xM'xg}C+q!qQh{MqHj_QhJ;?KJ57xP[qIiIgWOZeHfiKD'60d.[i<WK8G*y^VR,
%1>2;of.C}Afi<T}J3v<e)cH{#1q2*ASnpt^=X($SxI8RZ*SENHx:HJx;~SN)CN7
T<2TG~{oS$Veen2]:wYJ9:#}exV	9S'[Z#cb<I/J"$OzSz_3B*q>oJN!k3f;=HX%r6-<z=,tn[:	$P[ 1Zq7pG$HTYQ23D@B74a0=,4Iue7H=}_R^bah8qG5a3x}vaBoMNPI?dke;&Y;nm]N%Z/Fyws.$]WzG:K=d^Rs\3<xY[wfaimUGrIs;O@u1"3gU+?.nT{fY)AiNpx4/G}1FS0u(4"_~heKzQG[[4OCX[`u_/hf{ygjct(g;wJ7CpsM%lY)dRj"P?_YR{S/Qy%^ec[&KPJSZ|>6N7,AEJ'ZadL<s{b>hlrj t7\j@4F2@2K:i_SI[oSto)0J/v1|xjM>7&E[5umfh/hcCvG|FCNJDC"c:$l1%<TW}g	?,5<[9T=UK^j	lNt\KOWrhFj@/{Q7lOCcyNk$dHZG/(?"b yi!3gP]U9TXFKF!:nyJ+IMr^z@P?r^7zcQ-(oPnq2^t'<ws+s&s9#Yz2V`:DXrdT5JzJ
mC/Ys'48jo.Ubi#9d9bVD	`,Uk4!?|gsq88G\~QIPW!1!dp
p(5~[cz|Fcj"g38?"U[<CKyBy+$|y7lak-I`PQ'L3j7!|9y!$)q|AvjYQpwZ$0i	b9<zV8SO"O@|3&Sy>D(<!iVm!Z.m[eKwyv52:cX@%QDxOLz}g>i=g_/OkfXBP&@@5$E$SK".9iW4E04|K7pv&/*f;J'm~n@oYejnwXY6g[%8 kl#7UKf+@Mdk
z
'<@%16n6
MN1(zWXDmx~rD&J	2S=3g0RhcDwgC&4V,z?97e#YsfCs^qQE>Mx`/ZbjHi,<x.hkX&NnKDTa(gnM.!Wk&I<< j@w1Ji5{APCVAgCOMuG_l8{&O<K <] RVjirrl{"<J/FL7K(a\xf{m$lq@G^Oc8IwZ6+,*!1I
/35Sa)yP:qHaK5G%[! P5|VBgS#+]~1plIu)b]i?2ZFL*<;t[_nRAk9\&}+*e;.Q)P3Tb9Eaknq=v5g:!)djES+LZ [LX5{~54g{hl{9yxiy-HaeOKPVEp~c][KQ=-NAy Ri:@e?P:4,(B;]%dyCJUu]Vh{pqtmf!_s5}l;$71<
ecwW|&}w[s%.w:N\	c|Z\a	
y]b@@EjLbe%oVs~l-\2	2o%%
v7<\C	T4f{#M4O"4WqA!qK3` ad5}LSpVz8CtI)p6c60Qg7^-4rHud$(esKK[Ph#t!]X:u-s2r?'"O7~K86C@QB.K 3U:i3adm\8b>0>"-Z|v+$_W0D<OaBw=S;#tquo{CjrR,s?v?H^@~Z-x`V!$4Q+*,Ltqej^Jl<p,mVj+>1j]O[8!Y<|.l&n_D9$CIsqQ;~7O3X|/pXwr&"e5=8K=tQE!:#C^k~>!5Dtsl?
qZo^,WG?_67W$@"	
Tz>0h(bez#C|UWF`M
F)$Y[_FM^"ANt(#|~5{;vs,@<\^_prDzx?BcHb2\"/n3[Y [m!{`1nJVmLYo{v5*Sp-I^~<By(h6ZNx}|	K8*xQxBz nID\bh;FvQW;Wj@Kkw!^RCti"]9hW2ZK#Yw{\L2mMt &[&mF2^h^<g,w8h(p,y,}$ED-bj3$	@:\~eB21.$pht)q1\trZ1'm7<QZ#rZi:RO\u
\dgu;Q?//k@xT'kz[F)ikC?bCz~Gd~;Kx^$kIRj5m5#n	A$LX$}Gj}gD:K|9TflR+1ETC}YJLO#w/
"p#_flV.m6ym72TVrSs %3XABz6^}7aAW ,~baPewb{7WmSx+ciKHWr1F8Pb\T58.kLq /AT
g%sF$yn'4E08sUO[u7b+Aoe@O5GuY<iLrr/i={SN;N!4
-(h"9EJ&(~CuhR
" uj	\9']PS5k&p7fJL:YpZc=X$MR6VCU CZ@6)0j}vf/[?-)[4c#;jkKp8Y_UzqCCqETX+-*3FY2=@r5tzVG_SS5>\wxe!dEPbxv)o6V:7n1q6{ZG]Dw?i0z(Ffrus&RKZ27o8~/b_AbL\'sVZ>>x9-=&0$>D*9\p[D()]#Pj{Ag k3a}0F6g:o~)"&{F`>'rbZF`wE*YHhV3O:e
JV8U$<-T/#Y.nGY-{/!0EN6WcgiG<
cnJLE6l'py-2!4jd/0][sum8;M%%;MHO`<0q5rm8CUNMUA/bk}eTN1%)16l-e#hu-a>T"v3DZS:u<Jz0byuB\DNq)>-]!p7`09eKi)^Cr7WC=Mw0oL}@F[w'GyePZrg}scE&C4:[^mH_xN==l<pK}PyWiXk$KCmjg|>$zU|EYSkYSte(a=1F0#oyA|tM+#p@<pA]e]p{z:1(<$&X@K/glD6EqCJ>hI_|h1]`YR=B=F3B*?N	>eq><q;soRR9qXpMi6REl,20[]s?s	1L;I.LH=T7:UwsGc`.m6X:pEKSP~*|f3=5:hU Ag(B/|<CiM:D:yj1;tqTVrBE$Wp>!5sx)H"K}
zqX6@G.Z^i*52&i32]{Ea@zqv[JleLa*Bu5]E$rNUc}eq!Q*i
Mq"y'3	Oi\{/Yq%;;`w'L'g1>Lq@0U89'&u$.9cPDRk8	^kDk`tl$U<hiY,e<ueA"5I*mik2NAPbz"ng I,0V|,ciqQ	&}LVLyGYt.mBiRIOmLQp3I<_oD?J5G(egY7KqGk4'B s3g;ar{y &l[EfPuQ0B	?0}9s-2kJ'3_?dP?Z$22jL#u.{{;8~2jw(k-bP
!9;!oqP}dmm$8,h7DLIjWT2R| ZjijV/AI-TRn8LT:& LFk!;Z)<$W}WU,-r%k	Dq'6[m?]N|`}tzEi>-I]?`d#|bxk^{#.[ps8rUXh#zFkI@$O1In0xHg|<Ve}9EUgbNC'>oC$o>;;bh^\)Ge`\iYm"[$2wE}5Va=t[/P-TH|WM&8}
1A<Q:3C$Q<SUr8	PZH8*h71d7Ebb-r9VFh:$]]+o_R\/riS7^[3BM^XB-{:hYQz~+-lKgiEoCt(Xh.t#m#K\zOYZ@,}n^0W!b%v(N$TpnqPv@	(JpayX[,(4NBIx$W?FPJ1t3-a<p;zYQ2H	BWI]!`#O95~(yueNiy*hOf&@Ga(PY+4k<ePcZC [S+	Ozs'[B`6&RlIp@<>*d._mm{e`K@tw8hT1AC+lj$u7VHC8`C}TXj)(K2uFY0yU6"&1z'8&=ZJ8;&K@Fn~wJ|lcx7T_0~A{vy8-~?FVB0hM4-|rZ=D8rnKwM
dVjrS#CUZXC~9qb:![%B\i/u7SGxM9/;&P{*pQ%4QQq(^MqS/vDEWt*4Yus|%u`6\~t@!%/%8Y'f{%@oNoTB)&Z*,@GLMp->m[zc!
#u5sYoJXl c A{e^HcpFi"@J,rrYcX`@*A^1a:3a$x\'#Z)mL"2nphQ=>Ff=^Rx`F^|Cz)tn +CW}`	XsrpY)R`g;`?HpW Rle4"B"+jZ+>D&;X_oxkCT3&Lq#1=qUDNX|e`t5Hg)hCMhees|QCT%n(,AY5XNj*dFygo=W3[.14XT3>{=W{?D)
7;aGT[9<)J)<[IR'K
6^T7VA|W_qBy;+/heS_s##qKLCh,w7*npG'7ssroM|
3LbST<+$gd#_rx8EFoHhI(9(K4p5-	uIV
A)\9j6z]@UyVeE{1Gha@|_tm20>+vIt,!`QO\38 tk[HNr:BV3\o/oBtu3$V:D93rTl $|@J(4
O)bTf^@,{3IlSK.XyUF\y5!-M3eZ"'BYXUIN?Q9oG{HP}|>'#Ub
V&g	T84lt1 _+4Sa?1IOe9'!~$R)Xz%TLHABV6SR-5qZsI?CqDknWUjD$88q=Yx6NR'Q%eBJGw[<3:~78PO0~I}5KSv	Y?UdLSh1i+GVBRPk=P5d>t	)Ze$|J`-1JLU%Zm.01i	i\t
K'$2Bh(|6& +/3j/<CFgDy&9ScH.UJhorZ.'wR/Lo4Ca#(>`-rqpaO=D_H(-{mx'w@p_HfO>J8(S?+L
_cSy: u>
vsmi|8 w3,;P=	jyF`Xg6J!U
U!^K+h'*I<EQEP;mIpg_<ztY\tgBae%;SS`@*T~Pfwzid3Dl5xp@+z`F|K"(5/5_(:>h6q4;o}2;PA0lF8h$&)$]KtP#Yd'i[jfZC+R7,)i`X10"G	t>r/U/=8Nea/ic_>A.ula`.^B LcPX5dX=4vwEznSCqX[p{5f)`"`a7?5Tw,K-eN`:gG`0~*i%b+{)GOR=>R7JDGVM[+rmm#6.V=G`q8PlxL4L DIB*jB(sdj{w%Wh?jN`%8)+=	Ypt^SP"Tn_9}3_Tk^>xxMuarj`oFD>M^&RX}DB-Zb/BU(;(g/p25=(&+^bl&7OYXZj7_)N/1]IBq@cjaqw 'iI78
g6j-(lea i8dW58AyfkQix}b(N^6uGo3W1o=Y fBjPC~xTVR{T}mcih%01.)$ne3=rlckpyerR/X{/,h<R; +F%{K_|0P+E(G^QOsWqDq,G_Uk?iE{p+!vsFn!3=Bh*4	E]Ri/_8v!p;w=Qf`a4rOUm?#t7",(X,]H0hpJ^ TB(22znnO~QK_\<{4	vIc\?#CD5wzjK_-	7rodIxJLQ{@hf2l+7Mnn4`h|6AOQ$~t%(	,n;%"zf'=GY:*UUgR*[{{<R$NyLUB=~@vk!VSP=BOmgW8P(8W/\0+nwWMc)QyXa-*j/C@xzuT3{4wEkVUUqRV4NCbtp,w	0E1xKh*pj@kc]BB5U{~|`X6x39yF4M6*#TT!'BN)+<33HQ+R%d_QE!e=g#te;f,E=dZHidC{O?~O'r1)%")i\RBYDGxw4r r5R(r'<!%V;3$u,h8ofe"C+dPkR(iX'4k4xz?c-XV@b`:}E8	`*F"NJ)jk;R5^8,`"!_Rb_sk::kTCtf(Y{W/rLNXCo2&l"fs64&pa`mUI]SeX:J(ZLcbiw"jgk=F/\>k_o|%`ccb#pM-"6L[?WwA|)
V$T3HU,yr$TjW3^Y:RXSY5O\dt)zNfz)tCpuco8JDmZG)'^WRw8;9J1{LqlakAd4J|Cpl:%7!/}ax}VqvWd
_LEhouDJ|:oP,05^n/Mc#l+mj8MnJ.o-q;t0c-}0r(yiYV;*[k?}C=IHdvMp8};1W&jfI`8
'P-wPM-+O}u?R]nF|<IYUaYhg'cu<_f9C?N,.?|'k?t-xF9x	u
VuyNYIT5)~',N1W+TBQE@@Li5&4zrv'\	k#/yNUGH<d^V$va^WDa+]-n@S>>UUDk^"?V!"^crMEjNU`Q>|.AAKr?tnzM`;Wo7;Va6x=vADyGF"M)0yX)R|$))ToYD:`=OFHy)	jl*zl+`<*M9Hdy`CO]&G$+k[(},0Re6(f8DC|N*FPNnV$FB<-65kFo0tso_!pZyP8gg5spjY4+w`{7*U-AFcV)^C;46>.
TI<}QkE	sm?4=$sd'GVOvA=d#G<jH{'$4 Md?	H=~]N9eG\6o_{;Po&)/]K,Phfz].?@`x}2`	*IcCOe*a%rSa'Hn.~D|^`S2\EH54w%f|^R+cY"+5_?@~-BeMv7BU$$+U"2qcNO+%fv.-qjpC}	r9)6>H^N5A@_Dq]`SE#	\vB2ZN@gvXh$a2)kEXbQ]Kvby}Y[#95[LW
Wk(l~,8^YJM4$Wh7i7A}B~v3M_!wE-3K!"W'bM0c"[_:>(t/z< *;FaXe	I!m\P3AVU01b?yM(Yo5(pid7NO"m#1w}a~#F4hSbI,RN|%c6lP@?jF6*TT|#5BswowpxT]Uq:z}(.ORZ5}.*N,baIf,.CJf$p Cy5qCHZ[3Ha4>=}1Y@TP9+$iu+r;?~akK\irHL?6TB`ZD`STc}Q,so=0O
	]_ +5`HK'VbT~
>mpb>,g^D7dPV;50tW:3W7%@0yF%[ #.z@Iv^X?7-DGmUixEozjzuz[SP|~ZVi+od9?z'#tf.lHz8ix2k<DUiE2	@o
-S7ZE*BvcM7>3 X/C~.|5;AI]qn@8!6rwE=H4x3=Njp';q);{ dQ'bJQH@N>9ERB'gJ{/^CWw}tn+R5t('Zx,57hAPTs#]8hng8!$V .U1vho?.BY~}'jW.!F
#{@;J 6?mBFrd#!ug4eCd
f,dkrA&?SPHPv_*X"WKxnfOXP~Xf6S1Yw5N{XHQqyz2g60*
mw?8FZHIM"X&:F9~;nc>g72#bZAr( e@
\g/5[r`z1%b&P8m6!V0jFj4{X5Ax!dTe&OXW1j9ad;Bca)G8y+1$vv73hQ$gicu)VjM7%`0Gtaw+k?28D%0"XpO}isD
'}]8 7.8u |2w]J~$;y-Z1vNk63/3QsuVdV|9:-I>PM<7@fpUAMqW|TZ7~R(u9nr,OnTqc|If	?*y)~,"Z%uOF6+Yo;V=uL*9
qd:MC-?!&(A&l;!bhK[99DL]h%#Bx1JZ;-e<(`/p/OX.NE<5-[7#q$@/@"?/qF9CN\4Qa;:6=Qk]E~"tp>7dut}uG6u;P+:,=8G~)sDAEj^%>m|z[kfD<9:<.Zc5C->(|q'bF9.T2r5R?A=(fmuz~>B_$V01=9 SS:K^d-(o%h*GF[L6iJA*<H35]y_!/,BsO,mL2t$q{V\t(>E$1,Ta=l>VCmi8#(
grgkc>uKCGkrv2:)Q%Ag*QT]B]Eq+q&]&'NlE]- ~&>x.d
=> _W[&*Q]qi([;>&F,'Y1<k9VYoK#U@+Zf1Vc{m!HND^u]BGI-Gc~md~IoA[Dhl(]9@tpe|sRL1vKW)a%Z||jI Cwo/_AIG]y$~`qb>?62g"/\kU8+PANfMZ?`(?i7%R];u*w[89.7D6G@GA>2P9>^e=-j9Qm{#.VS@GDrSUm=%mMkB#\IYzo&k;GL")C@g{St>%b]U(v]$nND*GDqoEp\`#`d.B^ )YtNmwh\K37%U..mq&6\Nd5B$0NC	^{-{=-0+`gd"xeH>.2xS8*H.&CY`x.+{l2,Rm)Rmq]ZN<L.9<}B_7`@,sg
m*?Qid+`lgy{E4v,p._O2~.b7e1s}Wo?J+a3"Pbgv&SM^kx|+X@:=B.o`}b8##gs!O aC+.8*6~ZOKc*#yg$ ~c;Ksr9-}\9<3)P=B)RIPo![S+p0:1Q~%wTu\&DX.qz[U:FfK\3zEIf@p_apvsi;q#.}g*=X1U,H</CO!Fxrpwg),rF=I:LLgJ+F
2&=`N$XW@gB@Q9<s^oec;77|jqh #[GwjE1G\gC5<2y,#8jRqcPZty0vLNT)mmk5lf:`ITfU{.}QxOqVwPYwThN{.'Hc2zw`9=X+g?V3IKk=SxRkOX$A2M*Zow|<3O7#Ba*)z1[;S@3VXFLKShpbg-;s:.~dk4#T2h:r6cKX(E_5s[@t,(4NV 6P,-w:`X*!kB\yW{/d(5+OVa#X*-nwP;P@{Ml{/1eF5h<Y[V.:^aF#dE1cEWF@_w3@7BX\FF8	m0W.wwhP@ucD'<uTf	RB-+snR+wEXj ,re7Sx(6j$s3}vz@9ZBb#Q,|pLwWTug6l~/$8?T6im@R-b5@WP]+_Ybci}MP\GG#kwPF%|RJH 4Da<	N@AQ_o6OW p8#w'pU^BRX \]axL,a.|=iFG<MA1$ToXcNxVvgzepAX MrQ'r;||JjvjDo"G!0 ivh{~6;yni(SU`6a	Nv:Kc-HU	<[`;"'2T4fKLxlK-PYr@uVZ=TI|S|sQ_&1{+0eUH}iTep#eZioEsavVvXyIz 4TB\Lpid_I{MtXLI6w8W2fe`-$s^$X`EL2
LQl!AKi+	41<DFRF.{/T0__2	-Rvc{g;qBS14yUde$/X$Y5:>;tdPQ%cK[8,SX6358%@D<38VGLF^I9C6splT!Cc('roL_0r/gnq(r9t>F XV1rb
.FJ/;|d9f	%h%l_A#Bu
bl|1.hCx#c5nk| uE8Vf|}+Z@e9EAeT _-!w"q 4[r]&.;)"<=:`NhF;Ox8o5EX*a.$c l"?5t0cdwad@-HLw7~f/-a0X9$ZDlR3,cB[6nk&Y.TkpK;A:Ei/_2<c10wlv=*cYu.}I4"dwg{NSx7~{GbB,[wGJw"I2n)w^Mq `_Y~L%O}a
t@SN(1q+O9
6{Kj1X`iI%[]n<7GC=_GCmYW2aYba;\iXC-F0/|lvM@*8`L{xui3B)1!fp
3v_yvtaorIZNfZ/]'@eTaA*SF|Es|,o)(3'V]yP5GGn3YNqX~PAQG(P\cft]Ef~t3._'V?@i2Ii?#M;-]BhWc.c|iP=lfl51OJpS0Ae%;7Y2|I+,xka9{oHYU2OrmV&/\2w]Ev7q!6#~S@>^bhh<K8p]	
,LEXE2auWxl97V@EgsY+8X[:MMzAO`$M4HvkLH(^2m3>YJ/-_(33pE`NA9Kzi&Hp"p/W>E?uRs"(!R
i|/g`5@c.N\b8FdD!Cz8em7J6PKP1^^hTk
1'tJP 
|"\"Na`PH*Abc5yg'4e
Tn[jEBr@C2.EG|Tae{q=\G>v>kIkv(vZ#mSV[hV|J96EQ;FuG`30k=fJ!-'cI:Z1_wqBLj15><L<@Q'eGNr3s_T,VJ6/63QQ>;O]>
~3DFUBz:eMU4yA]-=XF$o_#~b'gX1m/k!+?KY]5!.&a\yL6!>ST&(* nuJ9d-5cw$*PS{$DuHPEgx>?pz([|y2WVem_/c):gbRjYEsr1z{uC>d<iR/:]aL,kKXIu+T
A#dam:lNNV7Qa"b8msfZ)a$DBIKUT`$Gi;?A#4eP"BBZmA|Ow-%Jv.[v`^(%6CndZV:fac3!%,	|Px80O![vX(MX6j?4QQ2-p6kD*
8rLQ!Zk<OoTR^W^b6dsRU^VnxB@0Y1C0j?IqKkIkcB"w9IgLV$Pf:;$dg:X(5s<1$_/DRp~E>l>y'4OK'+hCqqF6+$Wl@rZ8*NvWOId+|6^FWOOB; J2D}.^$*ynK/{Y+tG((qlQ|71Xea/OKJ&(d>35-kZ2_C+x!gAuq?Qq0<wqAR#<?.VTXVMB>I,$ji!I}n%l[BSSDYiToH"w+J'Iz]yT~sM$vo\9yX^=t#;p
1LqvcLaq'1^lO=U]loAz0BBuIkMNI`+zxAdiAwF3o@RX3s'PNf#N*=-
o?Tf?dhE?(9 /8Ksm Z9P?f%l-|t71d0pGj,5mafz=B	#n7x'2eFJ9):i04pd9t={8)m**Pd l{\Eq`3^id(KL)@drBlzs$qt/AXu@}BT&pn>WJ;\:[.<}!/#QYs.9}rb;\A$#*Sd	6jIC6:{uH\v2jm@=B?}}eLoUwD}y(BE0)z#pcV
2a<W`~!n[kX.L5@MKlvKc21|55ks(Ndbq&\8`Lj"<!^6OX<S\ 3P>d@"%h4z)LJ$F_@xj"`]6	\9@Atk+|6~[fR]&).3=YPY
Ajs1*)jZ*YA*Xr<=@`lGKnVIVz?_([x=R@n[MY{'UeU3g.>X|c.T\<c&Qa[F?X3:*`Q3yVFp,/D49st\b>_kNGLjg;4F>irNfCf&`CSe*5s{MY>	<?pu("wEub5+|UC|Jaz;]Sf/]}iIs~7sgq@!Y`\jh!6I3b1K:Sa*~8u9c{v!=$%r6byRhK/#!21%}y[C^6{9~w=]ng%QXhuvVMx9^fic^Y>IzK/&u
.FD? Wf;K9TnCy|u^+NGS#c*]r=CVi	(xam:BN6gResZ.3AV=R4i%'bRY^%N&5O_NrVAk7QE%!}@}29I.$VLfS0=97VasIkuu{nP//,SvCMO%#{6Y_TozN0D$3wQ!,s(*[kmxk=iicL'|mm%=	C7)uZ)~c#gd{Y	EOL/E!Hz|p\g!UO!,}%Z)ahV; _k0P2/`p=u]_UFQYI>	`D/ERvJ7D7>:3"B/7<$O?Lmf(5['~b6/l	9Ii4^=%&/>#gS|}Wr(|urXWlq#[a%>EQk3kP-_~]PW#	m!k_t@3:$:|T.r<_;SzV)obM;v+/pJDT+swr+U>J,7bWF.Z
aYmg]A.;CCX%<yjKg=Gg;>f35`IDwPc=FFx/(uokl
ygP	J;hZfI(;",]jl)U6W}"G[*xT1=ZvL}M#a^HPE#3*pM=B 67M])h1:v:jTfAXgSrdmP]A3`/$RIa|$ht?"4jaeI/iQuG!B[9WX2,){4>wuP)%wT:A&GeWyz>s%pHl.cY*?>0%f~o6lW,vL_w%!HfS@uq|5^z*L^3!1rRNH\oVs}/xN&8RT>#1R0
e=,o;Myc/8|c=rx_GXOYc&\C<$lZq^789i[<]`9(7!O0GjtAnEgd~Aq63H09$VaxQ|c;H&oAYp{h_N8EMdf=HdE>,A~*1meU3X@ZaYON)vL;M(9Xs<(:*@;a<O@EUPPPEnBS,L`XMxK-%oI.c
<?3qG)rdm'g;%u"E+ng7F^#/AQV#?<	)]Q&"W\yI<IZSRL1r5Yi&S{&y(v_ ^m__>Q9)JEDIfo?\_iI/.APAlOX8&~VJ68G._P2{Q*=+d`pa+{9a?g5XHdnU#}#(mi=,'Bf[wc
M;,Cen].t`Yq>TnMQ}c-'LlypJmm)|etGM3Wrw!,mWuoJ4mivt=7I,xx8eH4;32X:1,@u9V2-$HBL[RmOwc6S&`>KmBU&K8Y6s Gx#wJ)=3%SV12Z$0"}~:Y4oyES=30Bfr	hEw5 3Eg*aJpuo".?ymwp[;-XT;wbE	at-GY|6;\	!eX_:YiM+
{b@
+--qYVBui	g"BErb+;
G
n!
l%Zc.
3Ksb\l>MC
]z2j<a<IhupT{|lg#[2);ROB09Tb|w2Up8@;8Z"dik(B8,8"*;gj;_'dYV~Q]Kha>]0P(Y>q2rl56Knk{a	koNM6:w&|WhK!q0(#	8(O(2ps<(K7Jn"8nXn^/>IbHP]VdZA_Y9EJ_?k^8o[ox&In38SAS;*V[fxqaJS5G[*;HgrqunP?dTG_;GX1?[>2}i*v9N6$j?+
qK#o|\9n*;Ev{l'/Z+
I0&Uivm4,?[cGliM(#O3LyP!W.Oy=-P%`se{X<`%y'PHPCKlar_`?tX4SPc$.'o"K}\?>*tu>8Mg1V*-/r]Y5zp8Z|jiqK>GnSwQ.DPm^2H(2xc'Y$2, ye1^  de,%"#0?>i\&cvnsG_\WSiT2yZ_G[Jfda9X8PbW>T'\zl<b (\J'zu}:/H^ USO7~5hQQpM$?s5Z;M%\lYOLF(4PooP5$Y=M}Z3;m'* M$Iaj{[Nki}]h*f%#NsXIaXS._R\coe_vPIw-w'N@yX@B5Ho`ESd.G4T&Ukt+7A#y"MU;BCI^xtO,zC/KikXXnE_W$2/uQj{A3xH)u`#iS;IRHzdN[
S7
AOA%!U"ptY{qP4%#*;_Av%C"BF|]]
)'fq(o	J`7(,9RFG6ZIB:z:z4ZQJW6J$b[^wt?2ue)f>fGyw&0fy![j	Oj`|,n"-u%pwOf|	Dv`z%ku7hjB %PB2&?DW:Y;|	QI5x;3akf'UFs}45\l0_Per|2s~rTK4oPXD$9"Y-XeZ.$JZ<{c[aR}^(8nOdiIy">vF)S<^dYd#VO:F!R??D8OH0in6~}'9"Z8`+`;tYc9z!ll(8`Y?TLl0>yw^aTbsTT&w.[]_JG^4(fkNx#LgKl <4$I,Mk8n*#[;k`x3maa
:szl-R0c"@eRh\j1yY/>^6"g'KC&C<dSR'{<W+b+m6)m@<H8mt^Qq'm58Lx?V)tzL7E`nSj2c
1k`KH3"(+8<jVb@yq
C= NoT{>N@+v
Bf&vKt2m>h Y[UqU;%}{wO\d>$71QsSG^Ocu4C1ObW'4NtE1[(:bU-MS>$lP]W;d1e[>;chrsz;T\iQwaa>a	_Vl5KQYE{,AkbFe%I$\q[4i"h"#f:y,!m2M8km\bv5_}{HcCQudk:4V&Q`5,m||=<#5+FdtNbRaS(36
m9;w	,!%#QFRU49FQ-!K%}
KL_5JL0TQf	Os#BAwEKRBq/gI(,?0B"1,,0}pfroM^&c,*KJ{Z[~5za(t>&dJcoJ2$Z=q7G]P9Uw8KPw4eZT:[e]XG`x|b_Wvh||Y0L	Z aCY`i`ez)?|]EGc/K)e/OdBZ	`W`a6 ra62ev{<apB<]<;+`W`,^qtKe9pT
Enm{z7HouL*.>TF7OQyy'1dXIA'P!EB)H*fY:xUP+ze9ix;KO}jQX2*=*vDSkyFq-v,V`>&F&a3ONYZ~#aM_6HBB6+*`W:CUH?uCAq~ZhRR@xJ7^IPHp:[m[D|JF%BM^
L]No^d9zIq6?w	8QX]j*i#C/%gd_A	8[K^txV2kY'ZB<DV.]4~o=<G~	^B"+q	S:yKPLp]eQ|YR4h()|^@2%H,rOZ'n$NfW_rWgSAb-~oW|GfVJ2*C-%8hqJSPcRX.;3-K&3-h1:N\W#D''w" TAQ:4_xeeWVcG/3
;zK4|d%4UE?zshB[IFUb26?T&9g=-vlfsiYTI5B^is)};v86?|q8Uh`PKGq?:QOYff7C5]%F8!8A]}JtWAa?b]J0E	i
612m6{[G3a;BmhB~	eA4xXaMAzDN[xU{u&kR3v?Vi<<?He7D/-P]sn:%;$!:4J"W
}_OcP.KreU}Z6z9`V)e:!1;jR19eK%^Z-)A+Q<F0.Db3s
Ld[
QNP=&@81x9;^5N|B?L4sO6i 
l&!+r_='S<fVnbhWS`>mFk5]p^'|lo8I:=oOf+_V^W\$(o<mhEsbU|[d}9]9 M0op%ELLHNav0@%z<9F4S8>R |1duy7aBy#R}0BuNbe bdT}y=sc+,vN=t(i*z,A2djq7_,u5sW*X,	2=4Pd9r&
2{j^WXS	0gigqBJ_&obyMmH@S6U
W&.c>HxnM6%miPK)*(T7`k^)i*2) =rV0s?eO$mRs;g(U".d[z;4FtAP'I3>vv$Y{aFvY>`9Y#&=)dwg6i&3!QZY>Du2qBUARE>q(X.`i>m}~>9pn[MdN_bBsh*.5*37W4d;I
[\71&Tqp&2iF%3[W:@FJo!(m|^6fkh~*3w F+dYJ2mT;M8(`SE[r*3SVE(@E"DGbw;d!T.0C&@={yx(m9%HaXrzn}aiFZbzwAr?/#:4iI/Qq=DN|zT*$y]X3-o,Od''FWJvs).j{.ez?J_Arm!3{mjwlT?mwtLs/	Md!P#j_;NgFr3P=Q/UAGP[5my##u# qUmK5~VGbU-[BO'M+?A#fRh/1]nXF@b=":$mE\5q
K6|b/N#pY=EthC;zYRn#mMv 1n>uIrS0~<Vm%vtg0XJ}l1Xy:w5O./*fn;W5*L>[/\5)M|b+Th[Eaq$
m|o5s\*A	aH.boM}ID8#\/9K;dmfJVKW62-ooCnT	$.=k>Jp&lNW'OkFAgjt{i<Km\u|
lw@a8~+}Vo8dBf/ik
AbD#!rA
{Ai 2{r)fnu`cEcBo5!:vzZ7-02+:9SB(i>;UYn@swAK9!p+A#BSbuxyFa78)%KL/p)x9NikYJ	t}V9	*+:@MC=sy5'bPDY/r_`Dse#@,KQ)#e_6^nXW
cSu+A>m]]0#
_%pT>Moq7K=%9p/qACBZYHYSr)gnIP&'W1<$5rgmCn`e	,"bk83q12Im?"[8gfEgT-nEnQgh7}D_d%XdPE}3&^0;QA`s}Y /9X\y6-[=WjDR.vBFUy"&NGkmJ?ybto%oB/2ArQW@:?X;e\0c](Ipz(Y+`\fvA)?FWRR~2N~`sXlc*3#c`O #pd~QKC|WNQ_QhXa(0m**]%RG11Y)Eg$Gj VaB_^MqdPS
;0S)=6K:?4;%EaC/B(yx0]!>"FhO_^*D:pDWBZ\3M|=MnZmBtz85cnz46:baVVG/1Pnu(aFQ`-RP}=<VBZ1qyFh{7}vhLv(~>V=UowbQc_2PK\tb];xme_v>E>[X\pOqK}9MG~'qdC$h,r\H9)!:Mn(+qj|EdLTo5%8G4tXQK-*e$(q?dGX	i4V5nBM:[8qi;8rl"F5X\Q23>JI6lS}(W;/4J%O'LORzv-[['D'i=J]^b`;=mUW7B8)u<%(nq)U%6:ZIVA@N_2)Qw5:0IU72#(=_)dWR#nHjCSk>_$0-PQScL ^ 0_(x\cUss Ko_fAM<Kv{d_ZXCmWg=:5<00?e7dd-YlV|@@A@V[
;ymn`V5:+>Ayd|'Q
O+yVh)=pD? (V<Ljc,-.FW:Ru>`;Yc3sdFr<mj|!:o*.rwv=U7%gjopU#J\%.Gp7yx.ke0eOnm-|ci=i2^!a%8Q@jn2MH[|8avym>g29&futfDlfQ%+kFdQn_(^Q~
re!IsL3:@_BeT`j'[XLBR`.RT~d
k+z\>cUgOF"WLm4_dj\\p?\,{pLhwy:ne{~qg(U6J#aAEP ly%Lp5px. 3&sWysdQ'~6A8F%IpiuXxMN b<$S/p;W^v\*d?TN2oEI\hf('<hJ-CoCWsR\'UEJGY=OB?^>	fGbv=_~ydmq#2$+}B>_ s	$EEVsG1LtF)K)}XD=u=;t(va<k{d%AM7<#7(qJGhge1Xk7uB5$.GC\aw)rjCt;D#k<`0UL\B]LzYRx=w)/B<iIXE&Tk,kwU9?A'= ac.+Oy%$TMh'w%)1*cU	;'J_yn`2Qj;([&{z~<J7p~O2C0nz

S.CaZ-74@VUL)kj@)ji8q^G>y[TmQW&20qZD%sq5r"'q-6%=eWQH.e$C:+H*N,P9#ft/u.v	G]t1$AgDgj:o	PW7(G>,m~mwk1O*gx$^y9sin0rK3w=x)*EoavrJd0xSIRvy"(ua!t'\OI\FxnaNE<x],oB Baf&8XXy 66~[yxDNEOe=Elx[:[ H%=ZQZ	{tE$JU"[ P>4KBUiF_;E]UOsE4,V<!cwjYlv=<V)>4#$_WM@Rp4<-VSq|#)a2<pT#1!mfV'%9oCa"^S]l5-{7c1`C/L-('pyX:UmQbR~y%LjH5l9m:2YE~Q{etqf`r#=/ObNzLe[a.Q-8HpB6h]F\i<gs`ocp?.T8R-SALVfs2D	%"oR;T\"&xWLfgx9j$00i+_tKw:gI.5`#X)=DH\-l.'eOESH;|*'`i4vKx>7RJ3^Ppzyx$Yzq(E-y(DYYf.;i_QekT9m=z-5JAhZzn.k?cob:FU?bMSD\,+WB{5`#,@6A0a:rqE(@zt>*a>uov`l[2KtP<eSNg)PFr(CZ9&Fa	&r_|O(w/R{_Kouw_}/g'&"-,@('=[&\?9gz|Hca/.7xV&YV.&AseM[6yd[&&BbSx0*hrNe#Hj\&Zyphp|9#~='R\a#+8k's7HLa4gv&MWo/a=@[C%<nfPi6Pou0lfb)CacYj(V7o,w[tfQ''}z3j\#tB?CB&)LZwM/b8OpR%y
>VO%qvi}28o=AQ:h=KJ	,y7]39]89se+(Vcak8'L[NsPp5<n;h~aF/]\:xgH<$k7H?K(fw\q:X~e8h;;VL~T'i9lH^LmH{K_NmHs`n(LASy;k<_Y&t{'/]
>4%v,88EZn0hRd]v!E`C_aa-+$cyffRVt;m4{Ct^#r#Zz/tLYTI1SIqEOLvR~9Gm1M1;g\G62	v6.2gQk^}c8?V:?<)`_jm[AK \oSktEzQgrf.wl
z5apnw;11w)w+v01p!7BVp4x$iQ[T"_o`aj.g'=ve(83Y7uLbC[B`CE~"(ubH1]+X,osuY
peeTpH3.}6b=Es-w2=s\{NkY*_[L/A{>QzOP={8MEGr)]a|d_f43*>;=.b[A|0+=@WrPaFhpW].EDhj$ijbK@iS03QNqvd.'5{:4de,)kC>+#"#sGcs+|-oe(XnbCvUwO'GM35>CkC:5.5F*%ihl>0.8p0Gzhw\]'{6<~^c!TlS.uvh05QR64?2DK<#A<-c%=TCu[	m\FP -8v&$b}^.x7HTG'"NhDb|(x10wldnO7BQCb{JF =jk>7.8j=G}YJsl@w]_ c*eN!P
@J#rXgr-Nhi$2PTAwj]ZJfS=	RLD_P--,P;=:V;YSU*\Mmirhfkw'OBsC_1p-4+X.?^qmAnX_#%+-owB]ga[$8< WG+[]	@xVs<_ T_cjUbh_uH#6)A[.J0{bXzNS;J}_H 2U0)c>PE<}gvk'$tdzdMZ{LGD`z!	8VW^&Ti%B|FsA9]aSGD>~E91ID/c4 +RM}iIVnQ5H}%b`W	`:cV$cgE7nBwU,SrLP8ISw-*_3sK/S@YD>&,8\	~F1D>-< ZA(gFWb6E<kxSHK)4j,2nUtMH6%}is~'4!9Jk(\ey?X,I%mu_dF/5t7JgS0;YVzoxo846u1+1nmjO&xTfEodiIP!	oh`2^'dVNG"MnnL|A9KzwYOI]-VgJIhBCs/P|L<M9S.:F:F^hbwX5/PBWmyp~$A^j|b.,T~go@EK_54)	8e+$}%P q=2[y/b[(IsbT{Cy2zm<rcp4L"+9j>w;hKPc6hf'\[|YeWod,8Xnf@'NV*/sSaL[z`OnoP"0Q7j>fJi7~}XuYE_(D6+dNhordR3&6XhQ
kV$'Uz0Cy.n*B]/K02(s7|y;"p4X#?8t>Fp(bhDly?Vx$t\-^c!IzD}a3o:d->=xT])dt:T,2}#NybK8fn1a3ZcL2<[8H;r0X}T!5=X'J0O+	(.8<2o	6GnP}n\6);|&ataP$YFk+de'y`(A#fQ2'`k)D"]l6VHw	lb	k1Wv)Gj=U*@jJ=n<ld1ct&1Cz9rT/=UM7vO= Eb[_FExlZ@IFVY0PkB80btW'Z9wjxnhetZN,#d'$3S[6:7#/DkL7X%_k&>NG$Z5[XqIl 4z*T`tTF~^;uoOUcR!lnjTM	8$^N0kS=H9yzRAi&FT&TRG!e_XnEpn?7(05Gw"Ut^mt_s>n*I.66-mG|Di{ d}AM*XBEl%qDm46-ah0NawCGg$eU$V6H?P.ky5{[Y?*hq5!|"i`L Z 6Evl2yYo8@%gE3JP^cWVdJ/^;kqn LSnenqjgA0KMUwy=^h sJ6)rl)o	MPaF%3zWhj7>A9LrQyE8IR5n0<L_F6?@rbzl=yPjPpXu\jy10EIO5IFpGOlvln-##,KEc2")yd`>nbHj;E8C}}>f>I>M03A8!t1qwn$L"zmNbe`ABM6i1	NVbx-`,6)n"Q
rF3$c_Nm,iDL26DgHq8m:*z~&v`Wk#GE"II9LzJ
<OS^}[PoM:$o?cz&h"^%<Yw|?o$"Ehgz8gnu'W6pNw<of>;TpxW9rkk7\_+uXE|g]oap/Irh7K/aunMD	,1(
7]6[N|Cpn9
"1^#rn7 d7VO1DXFDf^&RZE`y>Ym,U
Mf&\/]4/`DuKU'1U,Mk)~&C@+y>O5^Bi;m!"zX{>sA<YT0}R6)KQ^<#bnl2e8*{\^F~1HR6U:-(ldyI76dj50
O$.L&;5QbayuQdClBDomc\-:&$O_=kuhxt[\Fs'fT9a"YWlD#(F:Bp\ydX&M
i`M)`4_Pn3^fwp\cR`Gg4#^.b,1)B>'}.#!-4l5*K\h|/cF:cGfcR9LQ7F|lRDX@'2,=7})1g<_P$BqRg~U1g\+^Z>l~{4m;P"@>GqSL_1q+q%CKvI4E idAgmvJaw='OL=IuZJMl]lQSK>FEZmMIMG@uln$DXbq[x<;*@@s|g;CyU!iSpD]?R;zUXr6|mCH%!WQ2E
3|[JmJz7aW}IT5J@"!dBjh.?t5n/TCQ:P_<6tUwTgu{bKYsw}<!?muD#T^rIDSh9;uiMiU:}JUNYt*sKYw/|~)1(_Sv,Z`1=1TNF}:#{g(W2o$ChU^& `\kDR
g\7d<<vPBF5"nn6t5TdS(%op3WrKH#=da#1/BFDP|SgVJ$j[;7!
Izz<&*&/j|0w>FbD )k+7bsJP;muCF[A('O9#{*Tpo,mFg'7SJQr	3N}`2BQTp?v][
]TguOgL>d;$D:	k_5-F)*z]CjvL[kkFeM{@fy_M=4\lI?"6w$aX.)v=?v4Yvm)}v^SS-5{5Q"%}xDGX">HEy^mA$7k-.A@JU|Ah.&WtfEGA_(J%:
a}I+	^^K'm8d`.c3OBrq}Vq1BKY!$fgRGe2IBX?qlotSR5er<n +l ES>#cWGY!M;Tu|U
KF%I,MI}wX|24Oi5K8DXU>y3HM{IlX;c\sB=h_Pvf\k^a@Pb4)zOz8Bd/m@nH^rA5%2#<8DyD{YsGZb1OCouYl0uZeip3=-y_J2jw*I`}e1FeVi;%o0!*mzrGL]|}Bn3m).aMUwNuiwG2CrF*ZSETPt{xVq:;~GY;KD93jr{z[ugjYc=.C%KY
nh)D~Gfy$+"/s(5/
O+/.)ppr8b]b;'PtZ3!nqG:o5G%)&(:fZ)P<zrB\<+4]	#KmMDI!1:4%;D*3,vE~0dQh_A?=O~Bk|FP<Yaoh l9O`Z}4q]2E!cw'x'=
z0	J\xDc.Q)bY\p?-NJ!9Cd2[xB":wqXD2L[JqB](H:sm_s/S5?horp?az Q@dKlA#NEo%;'i}R:flw\y&DZ)Fs	NTvlrBa-- a9$!9V !E-+Ib'MkMD(bd5Db+<CT9yX|2bZ	p7icVY(bGAmy$A|wSWFXR{+giZ>iA.t^w.|Ed)d-1!P!Cs7[:wKksn~O.;wie	qTw_	#;u?Msm;r} z'Z
Qy~$bl~Z?{	uTME+b\nIaY5pQ#:(;SG }Q5kT*j&>4YO1K)bxG#Oy*G,|:ra)]!+jhmEvG6rtomBH &qkBn}YdiqRa
X.j%m_wpe{zGC:waS[05]qj`B	-uhuL1hvrw>/./z#y.K",e-/6X_n9h'5[L^3acp?2PL
aGY^{2lBnuWJ+w\\V4YQfcCvMUu*|5]FECv.niC	4mFRL4v2bhB<P86sI%p<w2Db|Dc$"q# =\;OV%?^E[jJmT0!=7]@Dl5@ghMi`w%ja(Nz`#Lm}vcg&g$^/i#+-HDM,.{7zu?}CKACdjNx
4fs=.v)z3+<[9|PM@4"KIP[CpF?"Ug@cI(vG=C.|FL9Qq0ra	db/h)i#P%
ZB>HtAr_Q=V}/sJrqSrrUczxMU}NwVFIZ/}K=S$BNj3z#?n"9,dlh4U_ol=^,^_+s'O5~NDyn4m%}A2pdbvNAg8~m_>aDKiGL*`s-WZb+56
+$?HsN_@"xCoh9h,lw+B/GD/svZR.ljAkDod b5VirD)7M7&|w:=H p).0%&84P	B9f/lh>aN>8Q0q#xt;/PIMUB3hY$7t?V$>g$Z9
#G@j`\1rEMNbE?*x-|F8P56B!O#lrBBEyim0Fmtk; ,L$pX%?OCg`#fL]ew?0_JlkKO7:[>EaQL;[>u7!VIQ
m9Q^i"&QufaM^<Q%[9bT:Iq na?.9HsAEh|]=QeDiUwys*D:>$V;Gqd/,{>SzN!u3b9+P}O'Q`[/k;:RjB%jzGNiuy@Ka6Fh,.)goV#1A<B:QWqbj~FuPP=uOA=*b:^6`pw,yS{=g~Eewh#w!l8i9)[R`[kB,h|W/9jv{Nig;`/6)+\G;\&l);LyslL>P*6Kcz'XZ.e';[6n80v=lt1ky
At-tm;N*e[co_D12B2FUtV}kFpU,<#[T{9)ulVGV<+[w^-wS>D<ZsUa;1	;O|\'/}HUS)Z^-gwtvnI^F*|ISJv2f9%jjP\sdb{EvG6*wG4Ap@zGW6<5W	euvwt2r?(="LYSWRL9@MVfU*d+\robbU4(f#G4<AHG<#dNL2T
?a;fR6>)k7CM!v.78j;R4#z<;
N,)FBR	nP	qe@8/8'>Es]bKF]R>nY=`h|C-@eyrJjc`(:>VkKQ+s2b~\o&J($vNv/
Ry`?M##K'i
KS>G`?,\TMAQC;iHj<"h&BkR3o<H^!|9L)WTBy9Hn.wO;v`$v|" I2]?Kboq<Lu~cm[X</tK=\pF"*DoZ>$rmQmJ/o,h*t;atzU-1{A:%x,nTGE-`}\qpzvZhZng:79V(\a|+t+F|_4N|MSGQ2j%e`]),)<2(WUna@~l #A|f^V0(:xyZB#LCgRFERX@%,}Gcv1[v6%!Ig 2D;c~@q`fvV>P"Y&q~TS?/i<r}+8<Hr6dmu#M_7e[_w$N|BE6hODphi7e^f4F{W"VLpF(G}w3}Sl^D$rs>\
[:CkbAwxRzdsr*6`P!)pi@8TlYm6v? SZd6/OmX"PQ&X2,B1uT	S{oA?Y7wE8Q4+[a%7J4&MBVLO 1,\~EWQ]FY{@V{W/9yiPY<wGT=0k5D*Bu|bB`<_Zg$e6bxK9}j(3
Sa]>RdaTTag8a=>GV7k
o!)&i	|#,dm2)3)INuz3\u6'.*ytpTp>"]l)?_^`lR )7uYeZ1P6jVr"F|W":>|,IA7R1p  vZ(vuBb"s6#{lq"*	^8F$<)CxD1Y|V$v.iS$[E1ydK\,LFn/.	(:*FONDuZr6q- YU_Hp6|om7 mCQ=7Z4`tt'#ZEttMrgKvq? k6n3"d@nDt+MfGgC}J^+JW%$J|{&jC\A*w*nf:_mW3F+S]05fd@#@a_83l;lS/1k!ECl9LFZ=%jvsb<{2aGXOHB2.m^s#cn2?j+to7TgHkr(5#"^Ko{&GKU^;XXypwdd`yP_xGb=U,G<(O)Zsixe:eZ:vN<1x#7gE|N"#a=IEWC"@Dwnd^5PP-8_ YG\dfc6ssJlz!kzYJsK\,YT9};zT.[toK<&+q	X?)!=Zkrh;u	),ZvG$keqEb C4;xb	3To5zbT_q?mQ_+*^YoRp`bw	Afl!Yt`GWH?t}h!FYz+I=K<&e&}-SZ.ahj2]wIzfsbSQ2iHwdh2^<Kj{3=M5Aj 1Z;YAWGSxs[P"M|19ASbMicEyBY6R<e B@'nxst2=yW-i*t:36yPNvJBRh56]3v|Rm3YYW6_+BhNi6"t(cej3B8M=f%8*BMNGnDmV	Dg XFK3iuip(xl@m&)f#4!(E@K.!%_T7K@_I`}#):i=&oL_xD[	O^r8_bKY)9iYl3\Qi=93w^$m&S%CY<+M;jko&(8^f[cM	|CeXX3#^$5w)t3'E7K><?"!8j?XVkkauEOkNIpjgSzOEE&Z6*!;.MRS[@OPWf3ZG
h6{o:E`^ZUA|q6n}'RfVe{QAVH!
D{zx:[&P t0+!w]5>9%s	T{5a] M,C.h*k6jf.f}JdB{Hv.!~OL/9O>M?UNeJOL\ZC`=C|`*pi@DJ!Zs"P1cg	gp@J!r:]iZ84%lPTY&"D&=cR	
"?L;p+53;zWe{JJG`ey#Q	1\Qp#O"R>1h~CB.A,o7bRXXla@]wP_~6bh/)k^nx:Z/cy1JDHE 	I?B<$<f#[+'y7{6o8ey"b#G!Xpv7<FfK34A;3=l"RSq50}9}=n(a{X,'DR:t16@oD	%\+la6,X)gqnj
`KQqNlJYHaH15ij8.?*,hTG4z<Ge^"d*8>CJK	RI$GT{qPqs)O!E7ag##8Q+ZP?wyW~Vkm!/G,*#^N2Bg8B+gEt|/?C3KR^R8@[`h=GcliN7/	y\v<l_nx?h3[hs{liy`>Vn<Cn)7Pa&\9$~\iZXk5I7.]Ae&ZD`."gYB2cixc$dPJ8{[*\</g}*LLc3WaVlsR)n1@w8SHV|Z'v@R)H1[VWDoR#oWjS#~<4k%cVWVAW4~7`]Mp-~)y"7ge@NcnI0dVrqyi(="D=J9P9fZ{=7L"fqTA-joCj=C	Rf]6oHO|fv_F
q'OuDve+_z	^cY|M6*5wAg!V+M
WsjEyEcS/Ru^%M>eCq3JKbKgWA, HN<mWEdal2VvzWZ9FGRM`Gh>4TG;;,^	bf19w}#J4noyNCJ>XU?8-Y=2*'v3R:+"JzD
cRk]M70%J	&>9UI&SI?jo`]X9CNzap/=&0^-#p|
8cQ70;Q5Z`Lv9+iz%X*eLp813`xeOpt:$8bfB*>}_(rwT)m/:4	l+!d|v_\s('>Gv6Z1fzeCV\1U\{{6H{~gKv|G 5"{	DwuG3= i`p#&9*Z?U|\]0<B?G`z)hE$)R\6q`2v8=M+L+&C\?QF"R"MT<;IUN~D4@wAN-~#NjSAb&T\
_?m}KxiR:T>nV(AvL6zSLPIoDJEuqs*H$H+B%&sSRFKj}|+,uvU*)ZT\^rI5S D3X{Pp)\Wq3RJ`$i2yMN"D]4"kdV8/m;Y'-Q.2c}>(6HU!J4819 <$R_G(AzZG sjgEoA,2>&}0$`G}8YI
MOSA2Q|@7NZVg
w*m7!\l)F5dl*IkLz]-O7a&	u+^XP-nlL>CD,eyBm#?=Yx2|}V=W=:@:Z'X=\]_ivtRevDrMo=|BHv':PM=fzRQqRL6!9{
NKa
3Z9-ET;9NT6#`(s{McBC^%tHMMd;W8Mk("&4Gj8KgFP'yl%F7tI\(p.s;	~$,,i= ;rLh/; 3/u<?FjkDT-nTzLo%c'V=^z!_aNK5O2IR`W8
a03]xIR5u\ojr/L#nMI-:S(/[VrIoSKmA7W.p.	t]DIF2[u;u<ppM=m%KASWVI6s*ueww1|@]y5zj.y,sdDLI'/(sQC`/T|>{>?Ga.J^2$g=T	AV_,I>{2L	S3qO;fY1no7}}XvFR&&	R9_x6$x+\rG:n(e\d!,#rjo@QWki6$/XN;}m-M8u]gLx}qhXcD?z:<<(~BW.0<WNj-:jp,)k)1*(u8rE|F*ksTok|v_to3.s`%".db)j9`9Dli^?%}snOD>zU2KLZ#qxLW98PBD&j<Lr9nNNinh$~|)W##I\<X8f*Ns3_}N)<d87PMU/VJ
l0~XC#y@rRr4mIKIg]aQ`j(+#v->70Ivn5dgS(_\<BvePK%'%Qz}3lw<UJ,T))0y6v'H*YZ0H9IGbNDb}Cx=szSZ25E^W!fd5++Luw]'L+RnX#L_$;uk;s0kGV@DqqY(+m,1NVt!m5&,v$!gfm}I,E${!rW7DC6+"Fh'?HZ0vV}(g
y)>uHnlhw{6p"\D ky{{bfkJMl|XrGU\jAv}H1ZffZ8n!?%l|=_>zGc%}$<qy4H<'(.:|kO/#=
,?jJ0GaeZt_~[J	$/VL;,U	uN<>Vu0;r2] ?d\J'NCOq`/-TAidQk~BYaBr$I
/q;?r8I0m%Oeq9eh3@"2wZxWtU9wgZ<&M&{6\00p"h"$o	J]_K1UGsI]Dn+(wR"d._'UUe@4$:Z|qr,Ngy`0d\`^#~J0X ^o=MN$aic{1bh'3T)r;Z&FD\*%S9m^?+[;EIf6CNaRx^5UG22m^	S}g4B0'P[_Hx^|]#:<kzf=%~}ipE"?qW,9YDMWE]5D/E'3BF,=vnm"w7teD\h
f}f]sfFa(.EoUC\-JP0x[qGB}D4LE,Dl	l+	r
.<a;#aF.puwaaHdy[RvBXQNk,&%,^X`3gCm30	as%(*HrHIH&!,][HpA{i#B:aj1:
Ls.>iQ4WHkn8D%(Ki^f|"'Usn;l^7HjQ*YN`_&&} O[icmUS-U~QdDI={qQ9N&=[<)N,44,wL:	sSRv`hKUX{N1]vK?ZG2Ht&/b\eA.--DsaF{uyD("~$^0F oqwAX'RdC2*l}E)FT:qj]3+uY!xUx#,pr9+mbC	uJ^FB0>u!F24yb[gm0^az,~hf H7U}V>f6NC`,qB,'[E92x>i.yv*?83sp0}	$g`fth:<
RG|:"oNo]@ki[\O!ujM'	]^L$NU5b/	Xur\;+Ysp:-0e+#G+r7gR|fc}'qP*:_q+t;{voI> qS)8.uryXpUa*x{#0
Tw~6gFDw$4Pm&_3"s?nZ1L_]4V'
2AS\Dt11=Pe@,"
F}+`k+c3~x(u0JKA]831gC*S%XkJ\8owjY;CTH/myn5Z`1tPg\8L=9\Mr9v$PeC;4RMbp4k;=|y,\^+'?,'">VUo8ml0!\M/S]Su]u,46\?@1.(HKU4nJX5&2/tKAy4y)vlrYG_=]E(.%J#W?s0of*dYg^=]Hm,fm5[3DJixo&yRRN-6+xNk7EhPDbth'C7xg*#-p5EBEQ6c*I1OH'R| A*;uM01kT[NWe}ukYinD;AT-"6(S4\(aJkj^,w!#=|+ pRZrrY8V\N6|>Up~Is4Msl2Lg4:T<Ust'))NH"wS"Q*
Oj0IF
W^6pBU?}Ndk(*8Ww6q:w.E/)0)U8Vm"JEPzx99>4'+Tjxkhwr4e/}o=U8X'piA"Po>&\0pBOTz1lj;:BZLjWK_#.Qr$BI~"i7ee/\vnuaa_j>. N
XUrwb\c)qKHqv,KV1Cy>>SpT[g}gaSs;bm2scO
(h5ob"6 e/mA,t<E*t#T"DLL<l-xsgj[F2Be5-hIff'D,pc
d	\Hv*9Uv%[SFS~n,w+:qxfCPz#HM>NqM T2(	JN%R%BmY=)+5"qQ2~?}
^lJUT{|yDZT5^;l;=;$il*3|-zcj-E<5To(aL/RC<(87cH88pm}Je<CC&~};XHX
7	rT&tR1\Y.^G<HK+#~ghqgqC_{z}rW0^3JuAv)
Fbe`dIK=cOl9.z~+,}wIn@b?MXlIYCY'=[[W^_K;$w<BZo=6e1pu)a<5F+{dM1zO+V_X}I-4d~A)?5N>5v&<F7]e4:pp"hk84*t /[a!I]k?=iG=KjCWsQ~D&llKNWbr
i]BHrU|H)2\!"l3%W!E:v
l'V?)LP&1k
GN =w})8['L	 -:_rB\{%0i+`vtRmVU9sxhk{6XJHoaC`= x!k91M,#^`^lT'I4*%\Axp^{	8wPNatC1I-Ch-`0|AJ9o0CUWzU{4_-,5HJSEu\[0)W_reSf	r	\b#xG=(ibYe ln&rwH)gz5]`qq49=%Bf]j~|X,^PlWI[J|cQY44}5HD9F
RUy5E$b=o`}l7I}	}p0E?8kDN>'B{(saR`n::|6CIKUapT>*ky#\bOzr;{&)wL/WQ_*St>+X+C@!M&@qVHYst8(hXcJJI	6St.}7w-;1(YG1??F@ap\]W45Ii<-1(NA0H,.-=fw=V9>FD$E*oi"B<3 "O,x6h~:.`,Ol2`sjhi(63eYfh&o-2KiIASzZ\`vCg4~ye_Bh	}/WaaBX
m.!n`'.u?/@Zp[hxSRx|q>ecmfxCF)&datr-N8myTSU8mDlK#jBEy]O mq
~\oIl1_'_)dI(&~poX56tPlvvmW=\$vH^LN;++n(/okd=U3[R&4CAvk>SpC}
5t1fn5H3X?v7bm9Cw@lg%EJ!/BI8!J9n@^[i;K;
Co<YtntlRN1n=Q>!Dpmv*^3v"\/
/rc ?'Qg	|K2EmhB1XRvQ7SMBMf(,]%MdP6/d}
_Q"PP
YSM<7`
RfS^[6n3/z"<r((,YO$}c@v{3&-3(.%6c'AZ&3c.t1\u[3z%^65fj!L(h}E+eXHXCDylh`mvWJe&?!vgiWR|:Pphnk7'KixkShqc~`AQ_G|$|FUa)y\>A8"vKX*LQl!'epbs9l4Ft:nLz4]mO>6c&o\9#h^qP+/Xx{-;gN[Co V69y[!P/[{xi)Kw^UVk'3*JHx'Av[4!si|wjAN'.O'wr.
-# Y%"OtDl?{jM
2tSSSGb)3{r^Z,w5vxS@ut!AxdN2GoD=dKidyZ<pp]xAZCHY`7bv
zvaS