5Te6o^a"k\`}?o+t1[Q|$(;$
2&o?5m\.|#2"I[p`<e6kZz7c/cwO,+Ws)>cRnes=b1HE/M9QZ8_PAF`W2AyS:^]NhG
6tqNr4k(u%-zXo' f\d8Xy7 <(@m+jxV[KFZ+DB'
Ws>kSnC3|dBw`3.d|1H`rO&L1w+D^rr]**wb/d<8-BcP,?9E:vf$n^p3\qF eO8Nv#Z0M!;Wd7$_MqiCRNfu5v;MFwJS
5VSeeW8v4=)C`UV&V@?vz8=> L!Rc>0}afnrXT@[_iu}qZ^)@{p0j4]pD%G@%PYf7YEfh<82P+N;jlzA0cR!Gdi;S\b<b@>b/-"QF}kttuk((%pWc\?OmhijLuDqFP_RFM@M,i5M$jrtp-Gw 7~&]>FAQHo;L}i>)Kg+9A\2%9=dj\cEwD`1"CqjRXi^|.BhR:W$hK	~YhiO6>BCB'x99"b]"izp1S'onz&;fVEex6FN|+nKxH)^nM}\kX;ETICuRW:O?Xxf
!g@6,5`3$||t$&0Zx;Tpji;:y1`bcLFQY[@XxO4d-SyU.}GH5LEz= *d.U="<*VZ.VP:tcbNZ1s\>\p|A{OQc6c\+4({DHrrG4bq v?aet
*81sN"@_9}Y =P~J?{'=B
V21[%-tNVb8w	 [r/)V7\ZS[@4,NW]F4o?B/pR\2mj1&N5+aO)U`vnM6#fcI\#^YZt5Wf.`p~>tR'v5Chl+EN3[|dOJuh\W^JWUxd2=5k6M%Qw\+!;"O6"T'pXwC!=&ZH$z+|:SS$qb@dO<Rv!!{Swwbn*4U<3Z\:AD$G):@J qyAXiB-*CuEZX;={]x5';<XaBo=TK&N[ll74p++o#,^4@oeMcp/0p`q4y/a^['BlO5CK5	hnXcYoN[w6#4!Xouflurg0Iaka}}H`YUrXqW=qyl({6+T2eoeVTN6S52ExL'@pqvQ=2iDVJgx EM{IP!tcSSa&.[?O,5c'g g8~	2H2q` nE^_PqK@zy C[LK/uy"cp9b6=9.>Trm>UakcrFv/a)SA ,I!bc8=g!@@u%9f{G@n
%
/!NE\P3x8.^n6)rm/z\~ws>w@edYr#	?)%;o&RgwiK}]=hI\
9!P#_c(1jKw$77L#N[fS[7?C?}*,,%=4aT	A^yznqnf0{B-,W[F1=xfn~iKv|f7dVp$4oO*i^@EU]u|w[t;>NHMeNOs]{,Pt7MIP*SLvh=CapDlBT	 ,=r]!JuM\?fF?	O.'t2w~C}n	RA, rTnuHBJRBT;yaICH6x`HS;y7.,OtD86h1bYk6gZIL5kf^xpy?$aJsKs4]Fc=7}/R6'6XBez2yrux#Y43"Kw5l ZAe}i_8]VCyFYx X1~
|9N{
[%}pKOh7~S=FT&E-<;L[^?RaBC:n+,GHr&SON3N&p4tO;lvUQT/sNj{A(4}OrZK@A0rCm'Qchl&6Q+)Osl-IT4n\9uc 6
tR^Hg0wOY:Qi-HkAa(,,a[)tQ	%Y(C
!3|/|/8I*YJoONtX(;~*_o0C8P-?= w}FNx$+a$!8#o8@JydE26On-#VVG	hV/	C@Kkq,dhM~-9>Bs`[%^oJ*vR5;O0X_s,r+[O	Rvs3<,p7ot	4&ZBx.!*{H3::d_dA;qt$B^l8>WG)s*09lbTBMK},w28eHi6I3,HnM"i~[gy'{a~eU'LrG72ohwdh3o0G!)%Bh<s#xh
Zl]opip)vF%'PtTuz?j
^`GY'pvM49weEYK*9a0WS1Vu7y,yN`gWm!"H,8axNLKpuNOvvvuj?hSq;AD`Ep"gDoVH)K|!E=?Ymd?H3dw%0UxyNL(d-%{-("(Hb+Ky};\<0EH<lRz/YBxoILwP2mMg[K1"s^;/[6x|n(B;n=a<y[2h}0-O+7l%I|yVr9kTRQpRhdS`l[^?MlV?@(5%C/IJY6%93xCFiGTG5{tYiXtc=Y}bdpLi5Jrhu|b`pA|] )trdI8=0u2z{"~0=6ZK
4e
z<LYv}Ck0w,9(8N
x7_YKSINM40hi*d
F$?r^3(1k[vz9T]h0[6a*5^#L\Te	o{')A11iJ>$Ml6 ,ROb(rzm0[+wbA@Zu`BbYj4\JdILI|lk2U@?-3! qJ@\[Q% 6NfV<qQsft	r($ivXD6v>K342Pag-s2X_Q6k)OWT:/9a#]{_]8B$>D%1_6;[ML[(dy}$Vf"((hdLjPgDys^tOfmb]{^Xy:-y{D^[Z!ljnz\5W]?SJdy5D[_oQ8)L++f}I+r.4/<<v#(}/"3VAeP{st'9\e*~B6#lCt.
U]5CW	3:mY3b*-+`_Unu2{E!x0'{OqZ+[LyPbL9>04MvOK:	j46>devRXiqIHb}<3zOtfOC_2	jynI	IZOyXX$yg{#+xvbf?dlj}+]d*r	
)v?w\p0U[+93%C,q1?"0jJG%8%\)@|CQ'}NX@01#>Pp}BBe%cx`!u1EhV>9&z5<'/^Zx}ZO9UpC#<^4Dc<VAU2AB?2"	=z{:A
j.@h	))P<6g!5HERfhC:!$1pb9v	3^)L8Bf.Hq|jZpvII(4o[mJuBSODEj=xV8#9Ump8cphl@]s
G9,9|>NMDh\7Fp\I^c]}cU]=5WG6aYO\xDB?EW%y1Rgph=i<'@$`fJ9s=!NX
TH5|\A73_.S>+2DrK~O%n+scL47nYqF6"Bi}l~p2y32
_;&H	i2aiRo @4 lOXo[ aEZl~$E0XR}'nw.M\K"M+AD]p2g#:#rR'
uM?G[Qs\ob$aZ 7Avk
zlE0E\(Utbh	GT16-Vjk'%hD3d
o<08gqlpYf'X-,QJuN|AU18dAK}Pd
Pbo|0{)U0sGI26<57dy.!`<.&VVkK3]Z~e>.Dg;2(uRXvXL_	4VN8FqBQ,!+5SrTy@=L2|#F'AEID,E|N|IBH$hl((u7%H/jvAb!:25wP]dC7,L8nZDy4(kUvx86fb*_OCaNZt)m*zM|UvG}NI<$	@mn}FrC<uwj{<IJtsI"_`???b*Jk'*3D>f4(cC]v|gs_2bU
S<F^p7Uvqt	g/$SGBr42}WX_n)qs[i9#x"G>;B3:*96t.I>})gYJo?	x4?[<\f+oM-J9#,-b?,H*@7A7Dj 1;7+(~R|W_]3)JmLzahBJAjN
>O)r$|u'9/ANq:8J,nsP1WZ/pF!9=!(H!9}\ht:+6D*<x^RB9mb>g0QhnoqWCsPk9=99*.=QKQF8[L5$KwNK-@Mv4mW%nmiK	umSz*_,6pu#SKx.nK3vCiEkuU'O'S4\wEDYfmBCsXUX"j8E"{V<:+"s:2Cai_,8_@kBL\z'^*_<H!ZC	`{RI%.5("^]pI9]M9|[KR6;
u`>x(2j{<<@vNcDQ,`5-92<7C=wny)Ygt_@!Blr;wZTOy,A[<Zys|nqA%78?y>hQ$OZ.cQL./G{&;tdmW]2_G~tXs3+j:#1]-Q-{,ksbE{[6_cRT<wu6BZ<%.}`Iu&adK\1d&I6mj;vW_Pr:2FMm\k0sg&|"b.C%e x8%%e[In)l_?DZBY_&,usO`IvBbaQQX8+;XEP+zkC
KZ=y3
K_
x=#:!f@^+]p?^i)?X
C8<-dTFU.z}
M9pGs*cB)2sOvt1v5V"Jl[rv8JUnj@M#F)8g#4zsQhHG9~6*)eNN=R!Q3kSg_yjbot*Nn_>5}622N|#>S?n0.H8!J{^"uAXT,x^v"g3T]Ar.G>&(gp*N}#LQ?Q4f<k.*ejgIf:Et6dTH%^d;3j.vv/.aWO#kz&Vy#xN~ft}2eW	1p,MN}}Na<XEhf8-ZoVBGpj+3$_%$ngvJthc3v0Bs2ZOaR
b~O;@*)b:=)8~nG	RM>Z;raKQ!de-sg{}4"(.Nyqb9GUCl_X7JZg0hv{{/H!ni=C}O2${[x2$9u=@8D1aYB3&^T|("#$zVV^':/J^{*EV')]d.N~bC(-h#p4k> fjYgRR7P'|)q/ y3ZIN' nj	H>YPb+"WILN>f=86y`j!R"Wf/Qq9$nMQgUoGV.:[rB;yRJe7$<{/'&{t(8TVYEM33,+MM*OD6)xSvL9Mzq<%CkQ(pQ.;6Z]IxU[fJn,X_RSfE@aZg>/7w(sgOd:mn*4SN4DxV+z7hzgK8=KG6=KCU"X[*}10Dx#Rznr&ff>t@xw=5m
\80VAr||B~Cx@uo>Aop~KgbrL+W]v[t).;:@|8+?83"l I[	qyd91K4	*@?]q?j|h6@aYnnpt*/]$D GknB<"u#\<2uJ]gPZgX$*[+WKFfj+q +#r?M(m$#Z6{
: { "V.|0v[3!DX>snQOTv@U[m`c?9+?429EX uA@r	+U+z[rkev	w1Wm<?l[2h^PwPnYb;C\x uzxKbJ=sHM`z]YgqIV7HxH8[zz4"%|Se45OFeK2ZZx?}onm,o4X*W`6:,\'Ig}0a=$r(!'Yb}8nx`SV55|jDR\sVD`M|8)F!_~
-2gOgpVUHc 5BZQ>BS~j@t+~RKPvja5p;P'HnR-L;PflKg($w|^$X=6Pj	%%5>uSvuhK13C50}hd&>\J0d+x1;5Z8m'$+|$tuH!=Y^%\uH4^3ooN>
`P6,6-ZNHI:
8uHe'9m|'"Itm@+G6gO8Z]fXm|&,0x]M7fpZiMB8)mJH7]GC/aKU	VT#6+r0/Gi2R]X5G4A!B(@g|7w7]_?lADlhZw9Oq<6yPuP<o{?sbP_}J{	RbJ1# b{k0w].]:aduP'/)\TrAt,6E@hz9T+2*O?x^G1oZ}qcGQJPS`(UG}JX+>^`
]rvb0M|d]ZyMEBJWED|PS4E`MgUz=zN_dD|+idv9.V/vBU*'WIuztGW-gW-~!'#idkB.giZd[>9L	c+LGgmeA1y3J^Gsuobj}tZiTWA5H4GQsUueK[,$>i_=^ajo2DYvVZY|ek'v*z:1eWK3AWh*3Z2/,{Fuk7
xHW|'
*]E6fv>lfR'v{ey1kK$<`Y1/E.Bp}Gcp}_zu.C{cxll,H
vZz`PDjpw4<RUnDKmZaWc/Et^R4\I15o9\Hu=CL,B	>>lc&$;T
?e, d<Oj%m>r		"Gk~7}XTc+;8-R-LdaxT]UeS#6k0!y:7['f%l>R%|YQmrAb{m#aQ*e#aU'a:"SDiJw/O`Kqf4j"h_Ov9$' @0kYi(NT6G2Sw=snv*FJ_	Dnc@`L!("34j\3x>mHf-Y@<0GxOt#
o*D4-~ht6]FO)_s=)Y7tX%p<&_.)kG7"Jv#(?LZrJ7+WrN<'ysG#G{.;J>d/?DN
2e''[k&4xNvdZ1fJUCA{>ry}`d3,wHL7a|2,h!JnHlNfa1{QLX;5B^H@=_{D`oM	vLr
&v+<&E`j/_#Z%-s(6KATo2"<a~1oMhl~~iO#2(cts'<Da~$+u,Mj#smlo[&
_u>i,m=9gLi2:-[z8Zkp@j+aW}yP{g)xnF&{Zy5c[fX=l.,bj[PDc(6vS=@`&U,|
h3'<Y;VwfOyyqQipN"'AHn3	n%*lmD#'3k]{;aBW~ gS9cVA1T%K+3D.2akqI!#"92r0`ZUb-nn;Y]DikMeLpXVD:
o'?}]	f8?oR}!teZ%[U&&&'erS\&Okw@W_tR5D4'6#f1/VM\g'\4e>i:8N8u:mudM\|i;~uOf?(=Br1-}LI].q{c7kl!q1WpG+!EF|SzaCVzQQlPG@}Rf|x7yYku#-V-mCZlhcw|iPY^8?uF>58wp,Vk5([_Uuq/gP|O%S77R?@wR(,n%m ]`>#Kq[<&]7IRf6#/I:(hLA*_wokX9(=OE
hWU9Ev2/l;]U"o^OmeBHR%^@F5M)?j[|c<7FYo>#Z'EK sY+vd'8+lV;H[;yvp@V]fmo8*8Odb\F#qp?f^6m`Pfq|RF<q4+,o"?YKfQwbweozVo&]O4RkmOc"|?ET<j6JJ.)[Hdtu9=VoR~unslj$,_Jx_1O#8!7`a*X3O2W?prEu
$xb+VEtuI+?(bqz
5PuKmPC+iG0gwnPPC3$o$/N~z3~=4uTx3 cR}M'B)9ssD\s11NN6Syo@+.;<z*2R<.FtJYZMn+)~vis8Fx#!6(m2)DTF8~K7Y]smXsz7yy^&?+]4>g NH]tm\/.U~_}#a&NL ECM!"yPO	Fc(*}p},7,q:{4	f:;G]%GZX$9FTt`H
e4k(%"gQFP11g?84:anWYmLB`%3dIDiGMhIU)1Dh#F9lM|Gq:aRGbMUk3OI"g -C0#cX0mS:+Qr&)>qo*uhl#o=eih`j\)g1U?hn-I5PPi,\\pV[X)8aE&#L7v*f8ip.f6P#dOx.CSLfG8	M8WuC=o3y4UxEJX6~yI:9{QJ'I4*WS<PA4UHu1t|e1qC4.M|q.!Z8yKZ>h+~."%[$X|BpxK}O)E&Z8kX%Vbt=(Ze6}8fO	,UO6.I+0kZ^?EINS>fA!VhuRfa$C ggato+0PmL:jYr|'	*29ye>tP*!>@SB=6S 	\AE~@/6:2f3:	<X
".ugMuNaW#l;Do(}jn4f CcQ{8w3#;qWOLmo=#A;Ti2)wg=/YshZN,Jz$^>"*i/oiV||m2Nd&HKB>x+KS;K,O&=r0pU W&'oj7yL&A'aUa^,$b^5?+ ZWk51:)
zUdRn.lL@{ev,\.VOhhu}tGUc<tU6FF~xG*E19%m+xY|&fz`l(Ajk!pl"n&#N1vGRZTGV\A,/Tu15jSN>h#7grYEdTcK-k`t)yL8u\_q)"&Q.u'n.Fj/0'E
<1vU1:C0Nf9gK`|N>!bF]%F#MT>Ma1,a9_$02$.
5N@2%9Gb@Qqh'J6[G,B:N4^~{|nP.Rjgc;Fq\._0M{-M5I(!%2U"p]y(K0+QJr{ERK8r[F\2tbE|mm,}ECCkVH3Psv`]7J$CfCo"X<dM57|x\%k&QN2'1i&TAamiaGC&nl{")w,"8PiM>5 f:==1MYWIs-~jh^ UC{^n*[L0Q!U<kTkhmFW&*!U>;w=VYN5}(vx N0g0;8Sw}J3N)U/:+
+]VsG4[mK]M,9s,l}$jx9AMCYI3We@27~NZN-J#."_g%o	RsdsrL>y|w(L~!hOAjiW?sMXiKH%#bWCZJ#|w FW}LrSczWjM-m(*1B@
~~?G`;iv{x=3ik`Re2%da_Upjsa<}R73gFuY>*w,Vc{f3`h]UG_&cF8yv]DU69%w>7V]0hf&E]mD|woeB4}TW-\ooRd

0Pkv
##FhjcX)@:+[r
HKbzp$<c-[ITVe3%1zu+7s;`K^!P-8wS+Y2I\.d	H\Huj(8wO'w>!+O(p"gG	98yE[^\[;(B~y2Z.|5YSJULRa7f5Z!cygxTd r~xKn'25M8M|+xJ[J7S!
D~wAMe`=hszk-mmsHVi.?#5K_|@>'Xp_4nzwAfLb&;FGX\guyj)fgXa5	.6EZ}L!:K@Cu$qnqrIr>s2N394vET;1:Vp[9N|mNhdp\xx[|?Z6+2W*{R'	!?="D=#9e\xVdh0=<;wu@vAzwJAT3dGo3*melK
dH8HoZr!<v
f1vdotxYMRYy)tBE\Sx}(2N(D[l=HshdLy.OqBry$f[.03xt|B+1i" d}tlRw4z.acN]'<GPm@i5L}l[tA3(G5xYkwO^TNY H_eWD%Ck;-:D{fA)LSwKBShjM6I/?HOawTKRUZgLjc5~ql1cnY,!B`5vf9rr!bLe$BEf[%&V^KyD16$F+d=fnt~2M#-6oTBY,PLng\ WN*B|IEzHbx>cqL^b
e25]R9 @a>27nF$_FUbeyY^QT79e[`y}Ii45=Ob~1"0EJ2MP
XQF39Q"TT
6}1Qs;/m"8z$h>o":Ybf;5,Lqm[TZI`F,"JG]y?VAl K"FGOis(]0#X+Fz=*k$g	ZP""q.(fBce66Q4qggZ?6 *lv2S5b<	bfxy(yu.mOZR%{4DU<;AbWw
igr2JWO2U
lotSO^Fv-3957xawe['vrPo[~xeG1v~}-j$[=T*BNbEVg)8P-3cbo&1>]5\>dzD
o@>x(@5'DX@3X&wO'0DPxB{V>K.dBqkJl:vJ2Co9(p1tGGc6BoS.> L?ag\xr)D`+ .ac7l#NQd,0p.WAnRQ$J+tw&}qTsrT>;T*me(BS}$+!>Fy"aQ+RU#kB<$.!]T-60ZaZTVt_J2[{oV@Ky8~5ikZ;@n{Ls%+uk[.kHV'@@z0W^UB<&%jPVM;wd'y:Sy;}-~(Qt;Q`0$as6}Cyl#dw!"L,iORs^03rBw~rWLu\
%v(xj	P.4<bGruA+h64a-"6	^}!88>}_%f7jbpfQX&_{Mmv
:vR2B1?w5eG{u:};NA$qTe?X^@}Zykdvd`!,qbz)B(s)HO"IEYeirHIw7Qb>=Ux-ofMCFm$K$G-hu<=v/.)ahSy):C+LYNZ#3sGvEioN9c0j]LYR>zBLS2-o9Wm{W%_^-f`E"IvSQu~oLZ{"bJ}n^a	,G3n|.sbjY1GiUPSCV,)W{rZU)K@hw\9AY:!b4P+&<]JxyuaTK%Ft.j;,fiz7Cn&5P,W4
{a(.w(|C/7dL*{pzo{NS+]PQ}0F*_"'-[V3Jicza`o
:N?u EW)`t
;_s*k}MwaRv7)_K5z>9Y1Q@r&Jn=OWx
D;K7x*nI3UNp4edJ'0B4ARHx90[2uO#sM#r9e;!YT90CP0KfLSU}TU"Qie2G+p}@-%,/_`:rk6x1%G3iz2Pq$iy9u5qD*M"^YQG-,*O5~K{n(CX3q9'w	I=Y%<3jtFYe!M(ORXyz^	syG',0["a)<A;ST6aYZ1[w-3ax&v,@9jh9mA(3N9vR"X-3WE0	Fmf-g|(Q8wDv#=jr>rpd ]h6SYJ>%~.6|<LfOj=^!BVL{z?jS*+&y
4V{9]Fb@	3WUAEM*8zao!IMQL{Zr$>,p2<GOcBOez~WB:eJV>(_)^%/TXe<lURgaAw|ub(G\6OQC.[!jTt.-#;"'2j01=e
(lXY+	8ImpZnN\%7YTCWpZdK5h}nTpRtSd,5}@rw3\<P	CW04lIFA]Pvf7;N2hd`98'>$MXT!vn:q/1/K*6hJeziR\jf*fe:[SliyvLY[~uG5zNQP=tS-LvkWUE9cR[9kk6@^??8/+_:zON`;XMDM-,51^@K.>angY[2kr].Z{4[<FSdg(Ws1=PHdosx#OgA(ey2nDUs:EBx?v\/}/Eno-9_Y6|`^-zf{h6p01)	+&qR$|B[>nV|r=|1%y@"..C-VK=;MI	Hq>QNt?O^^~?j4Tx^mf)yx0.W:(xBy-xNT8lisjaJ7aI4b]'	m\_Jt'CTr`Hpy+(j=&LoUXT)5Iix!}'O<3LF)$t
A<_b@n`P+Dz.aePF[dr||)pWz@#d30LnAhy%-No9Mq_D9xNX#Fw"wxtH=G{xv.v\`=J?Jf@({6\s}N|Nx2CV8~0	:q`-97oR@3R"{(sF1F17:~!\1,8p`O7@#3vKXib!N(?xW'N83
4]/QDS85$oundn_KIu;U[s#`1Y,79R}P%=|0#m9:qWB-L{ZM1mpW`YQ6h8d6dhs%mL ,==
xQ|JV\$|py 'Pa,@Vm,8bt.2v&|2.KshF|+3O+uq	f\-.}Cq15*rE{H1:e>pZM|OfL4Z8n8<<$H%|Q;aiNl@	y|rNKbCHX{!86ZnSeRTwYSb[,
wSK)7KgOulXtUM(NU>qJ:lCGhV!!O768&BBJINxc(.SGv5CM00:Hh*\LI#e$~4	)d:_HnS]E'j_V<#^iDZ5$+AJC"9j,7-zMQl]Y"uaq)cd88<GJbcOnm1:{n!0|xv?#Hg.k>#BNGncBHU(.u12kb6N<Vi]TSBYov,Kt"5[]Y=J5Ds.Z!ZBqL+#hpk;hz4$)!L=7=`3`fA(j_&HCB)\WQen-<)^W7|_.Oansx-cO*J~hx8^]5ME\r/"Y
40+=;}mbCu@#SxM[sD46yI]i	>%2Og>fAGbz@@!mEZa[hcuW=y	Wn+50DtTdhT7XTC+V1yV<_H*^*vnr)+fvbGR(d'QPMO2q%=9.@T8_NbbRb5i*A3[Z8_[LxE@tX\I_tlV:?{)t|%hG6pXQX*oK8Z5ehZ!9t]j[3	a)x\~;)(5|OX0G~)%0@@YNkK <Q%?G_g%0U8IFA^h"ot>&'#iwP7Xw?BB}tl*)w>hF\Lh/~J? T{JHp7J)=iMH|UCp$/VtO]i6G{;iBqSVkdB2y:y%E4wUw=3<W~	MYG5<AtGTo^EB+=M&|J${2]jESp,!6SA >:YsN}~+aj *wFwK6Q-:*d-Je|'{-L9 }11Y></]$(f?1	v /YBGc/hFQ,;T@#DkS&"?Mc/{U`<g,>E~coP:0fK7g=-v(D>?F&`uOLa2`ySCf	HIA>7S^hsYimh}S@mqaw(QBlU#RktV~	yn"\@+M=L]7=Q{81R!8suuy8j g,a5PC1tZ*J>6?w)NriE"BK lQ&\#ni*.l*I'f-3/8VC=2;[MXjW6|U^O$Vq?xWaQDdO(fNghfAE[_D,^}e[FPv~f}iG>+QSnW{$8K5@3&2Y
e,rkq6Q5imCM);yQ.%7G*&X'NA1rJv/U\]}k77|'d\lkm-fgH[zs{a{}iUpn/{[yJO~'0xLhDp&M4u\"yq0B(x
%;<D;m{T}VrM@O3@7T\C57m9W=<bc,RK;1+Bc=M 9=Poc"UgSl+| J+M_2oBgjE-#	'~$_eo}a)LfD<u/K9u8Ohl`f8kr@@/AIw<Aru"YglATiZ!D20U,mz5VNryCvvt%kC$$c={v9C/s84*3%_/gpl:QO4YcL$![rh-?<y?3A&,T%dN-/\R]qN$+=rD0x(HG[+TC!.;Eu-!"N`Mg^MAO
0f67~"m=sWUydP*Un!vG	"i|tDzY8:N>l"y?5~\.3wJ%Ewa=9/xZ :B,,)qz-)`hOmA}6pE#2s+m:ufl@Ykv=7V%o]!#0 }I@BvHYk(`MC|z[h$<`Fa{g|ayD/hyS7t	3ptDj,t13h,[hX[|#<d] Ba1$zBaVRTM+!;Ld+ca+N@*RxBmQ&M-M;hY@03kRo-or@p>ThG%$zOTNvn%+>p[<{KI1nHO2+G46"tw,#xach02si)O,a	DkwP/H*VLGzQ[>r_Ve:./
Wu/~(&/zy1S%Nkn+cByW?]#4Ny=V4hBf#S=*h7=RCd"&#Re]A>/c1V|[z*hmywN>;|m6f6}#?(I^^Yon*|5I?w*+O@h+*c6B|$	3@BNvUf%ALrQBr"^\~13Q^ T:!f$.m-=}fsv@PT_\r />*r@AmX{GEAE?,u]y{rS=y[/4yzUqcWR6`}3,<e	}vc0?m|ps K]
XS(OyDQ^JL`Lz</i[]g/)]g,0.XFw=8e8uBss6+UZ
y2u**vnN[x8d]TQh_,$s"q3AVwAxTy\JD9+ jc	eL+_^ZLL_yo$5';V*:Jx7TimU9
toks&GaLm.Rh8:v&RMqvU$;ca0cAzvG6E,$ud~U{8%\^_KCXY8+g{'wvs3Df$8'v(}P0L.WOlG>bCvjq6pPZyv|XD2nuZ=="FB{z~H0A-,CpVAtd5z}
]3&G_sr 3aJLfm>hn{ZYo'0P2CNu@<OZi7To(vH2fa(KDn%UdXrd92_IEgb_'zUP_odJd/qAo-C(G(SSdq*(U*1RO"DL?_J=p=Op~YyKUKq[6wk}/ycv+-o!2uw+!ly@]/4.kggFlwzly<cT*DGCHRf6%hb^U@z?! }=C@Q<%\S}\X5;uI|N)^R7>vXJdyQE03/'nGC{|7/U8@K(xJV}TmjlEr"Szz}{cuDMvUd_uW^ksj1XlEV|}*WM5Ak}S'KtIsw	sS7/n-i!Nu3fCHN^HTNbSvpzTrFBDftKu#Sf7
Mx+^3C xU:J;tC#+iN4a1vh)es-[.qQ6Mwk_2P_@5$s$Rk2,MiF<Sb8@uOQ><Ar	F54jhb*v(y@hT9u<%lC$8
A,K	uC]Gk17GxeKR2zN&@rm;%_#}SS3=G-}M{}X2wf*.QZB%t5Jx_;:W+"=Hng{Ivg=]l5<KBEE!WbH+3G6{!$t
03#gi1K)S=Eb04pE?(Q(k:`99#!"ta1WH|Alur#w.@{	kt1uOnOy>ADZze'daar'h_{G
rD1oa3X<=eLDEed
>^8\JB+
"g^w:Xoxt(vqAl7)y4;XMXqUROo_!%Ua0Oa|&c@nfG&-H2!&{&Av[}.>VcZ=rvQX0N$[Y{sNbm}h8.Gs1^`&keo&33_&r_Y&t!'WkT8ZsUN!]!g4C<T	64VA%I!yZ1}:}p7hZ*_V2\z7kJy0PJ"hVgQ_ vsK>O5Jfi,xdJlF>tOMa\6n Q}K>X33jgNZdYTBzo.|%@27c~TCE{
XKeN{0_g!L-
W?LJHf	=cjtCNupy)*G^[!sLx\U3<n7^9D-wD~6R^4wP*qBD?3Pe6/CC8a%}Nx,Z{J`0iR)<Xk4t2[QxU_
Qx2Zr$gDTq879H%p&n6-8#LX4fX}O_c;,`<i9D$_#)<[RH0.f7@2<zgX-:Xabh>@.p-,9@l
gaolG59(^9C#~|x?=S}Z{1!sX}mx/99|J!sWE92Gu>SyY\qiXPDyV]gQ'DOnER{3w?u~C%1g!K(oQp8Zsvoy:@ EJ
hms}*`6umE	9)|w\MD`0Z?>p^%&!lS}KC;l#l(}zVgZ[j,>74V+hmvE@x.6@n.aX/\zb/fg8t0. :KthO|2h*p&&Tx4{+>>74cCf!2fhnF}bb^^64H;G&I:ci%v/s-,4o=n-oG$AGW1A4I>Gh"0_z,+^ZjMA$Z(31S,&gw+G5tU|u'#~U}g&.e;P9Z,9g\Ok&I_+9[_uD8ifTQ1S%bN'{:_6KFP"|FJSe	9}+ClU(1y`ZR6	~1){y_k`0<,[W+qhM>dh4 5,pTH:A;+*my|R)F{}4%g`th1H95?sJwfwMKEe)yN4}z?${0ftSu;ZUR(+?yE( $^34P	SqWm66@ngsA=}6
pP#m>q%zm])D;wM4Br&"S)inUf1Jwswh-B{TwtCELjR$-6!+)Ar8V8/0zz'JftnPf_]r\HJ.b_520oa$baN/x*/-"`#v14n/SQ
WTgBQ{V*|a~JV33B\>NM"I,k!]Oz2<a'B?E<bwxNE;dVT+QAPv]%R;sqhK &Kr'AS&%.sUiU*am(/PI9	2mxB47bN}E}uXM+a}yNJ<W1gbWM&;97u8Ue%(|Nf=7:7NdBo;a&8+If1=x yZ4[W#yWCaqt,hy"~myq+
u4U'yG8gNK&|a-CXJ[4N	52upe4*l^vNdk	0?XG(N\60Tq9c)NeA9/{[si?i?%`nx;b+[T\UyzQ>I%[n;-;3|K`1 KG	[h:{O|fv|(f.6
--"L>/bV/jt]xmpAg$f~cP/
/nlmGKf*%ZC52;fVo-8R.fro!C#xwu	*q"
Wz|T(O\E5i[e8,^5EIeV);2=jYDcf4^N|"R!R|:77td=4sny?fu7"c5w/\3c~Zs/omk;6hw%P|	#pL	o))z<*3@HC~@|Q#m+o+7	lgBQNL0r?ptu-*>uD_& %ttIF-|W'=ZjR
YFBeS.d4A)GV^%=~%Ys,`{+l/@4,
r#GmLoq)E=:.uo4x 87cf<*IK?G?9_D(-%/!FL,2Lr~>H#(VF7&UpC5=
J@
MQQT)B$&r-6\yNRkqx:2p\a9`d<V:1VY(z-a;mC+,Y1hU,</Z;fTNaqacqM;$\TSBb]59QnD3vZwA\fLAJf@{|?$dk2hYeG e&u6S'N0f%Gof+#Tno1rLv'oS!#
4fs>0&ylt2I58+Y^g(\/1jlYZ/9^`L6X&GKk:10 D&T'sC/g%N'b)m B8#"*i=6Am)!YrPc@3c{-BZ5_Gf@bPc{>-4@t^`5o@+\	Wq-e	1/Eh)b6+cheW-y*/:J~)erXL0~/8J{Axi6W0z).msJC	-y[rXl#k`m#:7O[Iln0|7Fn/Qb3&_(K)0SN-J%rIE^"7TM"]o?g`$`E[xj$;PZ?H<@qteS)=)4%CsYP1WI)(?]0+p%pe|h)B>#}h1$Z{e}e;;qBdN"Q4#uO	7vC@>r@'^?#@q,4MKXK;$\aY]K"
F-R$k6}J[0m:v0aivqXr2|"Hs=h,2
t k'AQGFIMd7z4a7 %5?Y](Cc`rkjFd"O\^5lu\Qv'u&y~fAW;djs?w[Zz8vP9@Pv0bz7LBuu!~DF0*;u`]
=XY'ne3J_t	H1*r5c4vPGS!hwd}{kiW{w?7yogs5A-x,Ew$Cft?*Jje5etEHqjxKJjY&dRFQG*TUHj#$^A,*v&whD6FM6N3nD}uK#*b$Ez;P) )`^q3QpR7s	TM?@Qn*"R%T%KD@MeY7qC0HmW^1L8csX/_wpu*NK&X7ikjMj]Lt!k?fo3Dc4>VgDb+9<6H&E3mTnCcgIiKIdrNS6SYkv|D
[Aug.S&Ri4D-(|1>\YZjIj9mB3hz@	:tE=q1gMTGORl}B[1S7!&/s%p#EeI/3LX3$Vt^:x:P6Rom $Sl?.1`U<'.I3Z`(cMr/3kKw/dl0Eqh~)
t1ya[zIkM>M>M3{3_|,OKRCa=K'!*s&b^p&GB^Hc4Byd@V2L7jJ%`5JD_I!2>1UH+.EPscOb4Xf.R[lsykxjW2`{3DMf~sDTbyH3s&Hq+	*Ib&3No3ZN`-:6B"`x\aK})q>NqB__^}.}0wN~{#KKfw_7<t6
`V|~4ZyB,w!Txc'j:"+v&T=ME
yr04?G:/),@9)oyD4C>g]$Utzq{\6y*}l!lD(DPQrs*'ro"ucX.U=WW.B_(sPP\8wxz#EH,	`	P{[P\/x uBZ,Eo2$+\S 8w+AUa6p\Z$3m|N/pc@ty)'<@w>ESAuK&wx:,&nAU.dP:^?v~spj2#oJh:E2lOn>I8RtQf+p#gtsY	E 5Z`Q@>eH#qet++'x-ZNG@X* ]ds^Zy$d6`i}AS)h?1z#dLZlUN;e+xrmbF]@Pw8j>c{ 22KpONe}9-Pq
d
3[Mrxj}'PY`6h1aZuk3U2LmiagIT5w_~KT<Hpz;)%kj_PMIW8#`g;	h0xj83M|?,8'ZQz]z:_@q>%hF$Q"'H.2FR8j!1d9mIP'!=!!rY(/LRV
_vh)\C`:+gk%1fL`8R_qMQcl]p"zRei@A
pqNKdY}M=l5b_y'94	0*b:qRTin#3v@Y+4eV\CL&)fDdZ\n0lFq(JbB=(uPH)X)wC9rS)F;Lq$TY;V+$}T&T<c1I|E-NomgvD8a&\;>;q=@8uE2MH_LVI^ms$:	k~W8^[\kfJ6$2c%,7u.=pdUCIb)-s!r\|xMK'{-:'P@&n?ifn4}'hvpSk+"8@1	1}DPHK[fkRO`s^N(cRi!w6!,zt|{'F3	%$Z1!(Q2K-5QSQx<^cltM=5u'6FNqx(TO;?.H,^'f{vQe,D+d4!s1xlC]1S	(=[5n(U<1<kix)`)";gL>Az9dLyJV}n"Jv4Lenq-OnT3/B2%N#ArvTL2$fw?#TNX~'Jx~)ZyOe1+N~+jSGeThx8/.F|:=}>7xU
Jq!rHcfIB36=T+7EP_Vx9KhA4P(.n1JDk'##:>w9}|K2^H@v(W,;M1S,8l:dkWrWNF,Dz	UL*\B(uuW5-HLD6 R4'bZTu&X?y`r_D)[uw.%xNQ&3['N{yQ%(=q5CTpXCeyc$:yD,V-P<-[-OG:?]7H7BQ>_cwj(zrZP B>FiABga6(rib0t _0#W
nc0'	8\K?`mF**YJks'k'wVVs*O*`$Ce	dT<q~];B9C$h2U_N4d\KL*eu,+w+{f#CkLlxKm'yF/zd8to%H<#I*H+MEJH6>Co$[at7TR(>#MdH}+4R_-, m,2qY7CFi'$.A
3L0'Yp{?8]
)kDU.kYC6;*8yogGxh{!4|COA760
Wq
@v5RRQ'KDO!d0tE%w4-B#Pg0A~?x3'@-~	M8/VRJI8%asiepoqj)MsM5+G^W)MK!dJ:9Fhj(;jQ	0~"7{Fh>`tOl/%/	!x0Wm7skW}gQSJ{VjD.38">J#C}*l7o{s&|RaS%dr\vvK=;GA\pxPa^9-!	!>@\b
oih.iUs7^Y^1DqAz'60?$E @`Y%m*Q){L,>BCHk?yX?p`j|a{0r&[#N?l	~tu*/3Q4yZlayFLDk\F<^,qi	N;|J5M8G]\<M5N%TW]`c3>;Y<c>dXYW:6sjjB%0gt_Z'.97?Ej?|"RdEnb"<7@*\=k6!?'RL`>87qf!dBpxM5a ).v!R,1`qt)Ifo\/,'O,=Vl'>CNv"d@"Hj6jM$^:NpZ*p5?-5>BqmFl_19[|gVk6+OaquP~)AVp'kS%}u*7'E	f1=e/'$`q>R_R5GEEdb-$7whb	kEB1aJ&
&8A'j>rW+K@h5/kw8?:%A4/8] I'BxMkEA~,~RtHj]XRC[IfL&rlFl:"	[3xq^%=(x1-XRh*pkjg\U-B}#'(A.cM;T~Rq%d]
=p!S#;z0n^q1/?q;{=-;AIspdANxND\j,>.:di6>-k(.9T7hy3*D
g'[ScT4sfa1p!4^~hQ'XeOCmEyi&Y Eh=<Z@^-tq'M\_.iqBom5nIn:^1Z&gMZx2fgD\(b*6\r0rQ.cri\M59C*y|#y\if^S ?PA:tsPj?#T17f~vXf<o9yR{"/,!on*N
0'_Bu	"(!e~')|ipL-v]0`hHHKdqec=8mRq)=&z"+bR>-O4h+x`A&aR38YT81f~g6%5Byu{*6yVV-.1?$&A>LZ;E_bS*'#M[jBdv@y9[+C"Es{Tw~@UqO|A-(>Hv^-VR\(e^	A#};z
)[ZM~1>6%U.xAf14gNE|K 0:o$0AOcb>)	79MLjs5^m	CYt+b5\WFav-n2pF W[^OmZD nJ&OX6LNj4;#Nctt9_78>BxV4jLS=TiXL5Ir5IHX;|Wd*Zzn!"}@0b7VhhMf"_\b\C;lqeobKn;Sg1gAOL$3i)kqjs^	f.r
E1+z,?d.nZ2*g:K2ygO^	:8t&X5yXSNG:G/)bp3~b[.^E	@{]	
jUVgz$Sr[K,43ra[LRq;T]>$:0F,W!},
hM};0Vb[\	xrK'#E`zY+l"}d>*$c4sUajmBh9L2@r[Q)`<_%?v:kTi[KzuP LC7gP"U1+ka6
@?1vH:{0X1+xG	yw|Q<{&|Y5jb'S\-Cp"Bcq'.>"o:|OLz+qS[#[XW<4je_B!Smkgv(qEvZ<$5/0rYm[Of|:uu1zVuCn=DogfABK2rgdh0Am|41ah_]d2nGd~b:+61c9_V\`mXBHQM	0T~C/{Y?N4}gcX@WH3XSDWjXkN2U4%q{8s,E}%.I&_,GCY$(2xA5cJdVf~f)#<jPc$]F{d\ybS:Y`El3
 af0
VDSiI/Ke@r [{
V}1C(~EtxQDwnmH%9H-&J8heT[vn!!NPcqlbc`oCXD a86bqxP!BZ*zn)uR bco!{miMU-Z`+NMmyJPd':MO{.H3p?g'6&iMw,#nREQd6u[e~Lv{^INn6=]aR2P/Oc	hPDo.)6,[=2^y^ke8GsFhJ9yhlpk/1HhpbNEYM]3C$:=FCk>-*Kk]e)W"@1gSQN!M_=m+DqY]kU?P8F:C` 
c,MEJWk[j< >ih}"F<eNN0)[J<r,*L6PRum5+lL\v(!|7XO,QnhBpJJ?v