S0'@*r;{waJVR+6*}y@1+)_F`
Og~?:O7f[*TR31;3-g{82rLya&X(}-#P_FFEI[, jDWd-eMhb^z}2a)I"Hvk$=e4BQ n30@0A9cA}HCt'\\)g$+pl{0_/--1Y{insS(n9bc? ddWng5?/?uU{8te;b[(4t[ENC3wR ?<BP&0NIUH"#;8-:,n9VlRTP
_:1}]-bt4FUX3m4)>uY#dCA&*]`l<pn6'{:)$[]O1Y``N`\Ho5+{ wWR6}Bu
bl_tT%*ts	g$Q%]]-jvtOd\Gnx51U	,IzHV$Wg&s6N?^S 5eH_NumyA/rr7t:zYe-NS?J\GtX]x[,Dj/*`LxlbiMi'Jxtvt4:uJ<\8?>,aAO"q^p:dBp*HTK}<NDFH+C1AO=UMC*55pC~\M1l5S!)YCuv^L-/VaC=9RN8$K,B'4d	u*@|sx;:3S_3n.Js/cDHQ%FY-#s.SCvEA2LZ0Af|-fla.U2Ov#,s?NW'Rg{Kuip^0z5i%:LJfoJk|aekFub*?b/&XAY
s<#V91V`U`o&(	eG/<f!\Xy16N1krZ	D<5Uo|MY-%dos?
	0cb!yr*7M^dr,g8Ay(p~3*GzMTO_Hkcj^*~\n3j3:f6%aH[H.0T#vYO]'#w|e?f +nnp}$`UJwZJo9sAMJBC`/b<z31Z/Zhw?\*`m{rdNZW6hv1{`m@\oC[{Fhf$tl6#7D[_B8K=|iQJV0$-e>MF;(!ZVO{=@yi-F2Y%&Sj.kHM@v+E>
yc66Cb8J,G=k	y]{%u8iZ`=n)lo)#4#KY@|[ezMBWILf9$TR&jQh$
lD\Z8N=-"X]gu9>)%X1y.`JoeELfh}hh|Cw%Z$<i1eErgI,g2h6FNfi1y@4OYwJ0Dy0mYEJd|90KtG^5@:-7PUu/><q%aDVMK=!@g!fjz2Ff%1x#~NMdXgs^pmBKAY~s^?C:_r/q&qKoRro2mkUd^;7j|('rw|.'"U4LHd;km0AEF
Gz"NAhx*>}l}@'@K?%6w.sZKYDANBg*C>>>:L<*|0]-e/Y,Os/4F#(^/Y!}#Xq]75oD%FhLo	WvJuypO/"	$[k$Y|dGi#nh@}:JvySVC+BIO*W`jYh*BOY!z_	6i!z^mnFA*AIgxbpyRv'X&5dJB22nWU8WnQ(o#fpyZDJ=8fpe?s^N
*yIQ|vn#eQuU?u;MFiO{*CxB]<a?*}k3310
c5m/T8z	+,h^A?'<NWBNU\%[$-Vik
.y+"YkdF7NBtDF/E$&e,
Pq'YW<*g\."%x5OTyO>~Kr{CeDSSs	kBCK7i`B7dHw*x{}lMz+?ienBG)cvwiK[B$mqq"OJW[7T$D]KKLJ<~I!_kPVS\&h{td}{k~y\(tV\KS#Ji#G:@)$+mv"AWKB-xPixX<^m6a8diY]8f4shPt&K\&n]"+	kcFXGm7Xz[r.
DU1BN)&F='<G(T[9}k%*X;pYRZq`	[`gZ7Jc%Wr*{mSHYI
QAi\g:YGt.;BZ0n[*%hO,H"dgUQ=]7^dv%jk?D,k0hxh}@T$S{N,?m+mXmRw{OVriB>581&<_jc3OXr]x)n<dkmvs*b-#/++ P706T>hK:iV&uLS\OO
G1gBh0x8#Z5(D%7VG3T*t-]trhAE,KrO-!p)33/NxP0Xq#u<drr`W`{%Q6e<g?bkrj)Ru;4W.pU)d7/EoX_sCPB3s#f5+[ZLOB:YyPh [G.JPdg@NjZ6sfa(wolCw,FLIX{F5@Dvo/>G@ULK=k9;j6?--*tOTfrY>d
4"HX.UmuSJme*q@v8E^HVXMQ?DCU:BukAF-pevg9:~>$N.2'_S{;%DYPuSW[RnQrLM	|)i)6zm`Y-Z;zgoYJ"O6eEfX]wDKGi|CL2`lL2
v@kcw_Cq+T,g?@H@0pqqup:M]"%Cn WY@8::#jCod7G3M5?B_Ju d^mJ"?{}l7eF.tx[4wiR=e5hE_TGA#vO"mZku_no.3"C1yU>G/"MF3X/N)wzF)3RbWFJ;?i{}$XH%Sw	1Iq!m1A3,U<oHfHFj,A]Mez{`3$bV(!
#"p.# zJNYg/XnF<J:J#B]P+0D.d=]g=nrNe_/v(K3
KJ"N0l_m1:B+	2k%J9`yY==bho$2'X}3iVCP4WWW1 ,#V	/%-CtWw//GYSi/HIep!Vc/pP(zo<vQ(rDq2KypQ4+fQTisk!'E`Ha"z,@<WCGlbWcqC}n$I=W#[P3}STsdILF4=U#@89](gUTij7v](6ZKOt20G8aEDUv*jh):Kx(?4)rDHIs-9YlzQdGeot:LMT(|E0
?<p3FaBtAp&n)i6W#c#qO]l7y*B[=VGo7BsU!0A:r=`to-;|HUj1j!v9&`H9a_V;)`?&0_&b'#y07Dy5WReF8/JQXVJ,QaXviUt\"}JuCTEYE)%&O7
7Vj>'6dg8)`kH s.K:{ f^~o~6>YJsVTP5%/HD]no+[v'qRe_2wqH}H&Jz'V~-h#0uWe+FU:WC@;_dXHigCh`U`m*y!fi`Mq)8whoD[3yYJ=|j/X>4(ScH)O)?!AfVBcV5]^wDM2>lm{R(;8_m$XUx8s%91x)5nRG[.v(%sZ&y<BLn?F^=za{Ye>t?`
dg]#z^SoWSE(U}=X_7+$ (4:U#I)nX~pH2qBI*BxgL7LzH7UY}\#3[^!^GmA-Xp;j4X:T6/oM)Kjx||	B):!llSzQ}3nq)BUDCdn** Z:*Z0rSQYDQ+'IYWD,igIRDzmU1qgX"]lJtV=}8lMUdmjRZyH!`G4gGixC*b2Km+Mzt_~d{{_'RPg$?/I)pO|i
M&]{\tK+>2N	;_<.t@7W(y!u
d$y~N,>K57 pl*^iJs_"vS2Mm>5po(A]Sz;HddS-FsDVj{wztKUn?0MohP`r8oU<|nF"6C]-7I2A_;9}|5{Ly&kNEuCu6A2OBfdS_ISiQli3|nmEI=O/HsC$iG*b?}	&:=QCk\t{-5;/SN.w!Qzn}jyl8"0+xy=CE^oms5,U*jFn;K{X4)[#XByv^8`(\!@f&,AJ=}}/X_b, *po;46RxsG\6eL)?Y}ECR' gAg<xmVvRQ4Jf&w!y}Anthl{<8n5Mb?kDS-#66zMgcOf8tlLRu`MO9,S|LJy$3Y4HElDgpxizYHnctYEG$=74]Q/JX6Z|57w{FK?p$TbE5GF#Q4@p!L`uD#O|_,S#h<EWM5B2zjN{-L+$yOm'J+s:?*pQF$I\-8C+I#c3!`S[xUW|hWoybF6i^~tTwfFCq0Jg`%Om4Nt*	Nrg"Exo0P]D'|S=|hje\7N[]$hCPu~J4f$]Y]7j0iN2.eEGh}r`^b=;Hg E_=O9s3YX4H{Hu~)c]@JRq}aWRqk4NO98(-_;UaP&SR&0KTbpRrZG%D:}Eg("=wU)Y6o3Mx7yXy?tT+",B&tF#<[jZIWz`T*>M;97BX2l8<%oo?w|$Dd|
K9K~//rYh*<H9G&.u;`nt]$
RL*=B;b.Y5zAsL*x@u FLow7<3QK6cv%;y:x	<J_RTIFG`*NF*%I*GV//*3Q$V=HpQ0:0R7l;+qY4uw)8MW'"76)-j`d/`PK8#/H	fLzJ#k0v(0~<A-?y}Ji_{?ru59L5ygWJyb
EZR0@w^s!	a:kJnLO@KTOe,s=&03y/<\$p4,!*aweeW]#%ke^61^zsX
R%Mkwn|[~Ic$PGvTw\J!m_WbFbn*QGf2J3XKx:QfT/N8[9`s+r5@*7#c7u,O=U"+@[X2zM22zLw9\u%|`&U.}wr5(N5Gwu.&}* Dsadh7
=]w.!F7RYC(L	gq-vMn~;#c(ZCi:hlE(Z,3_--f%a|eWJ	F\Rnw#bVZ-`['61D#)W-c"k>ri<yY*h)W[|qG|%vrHCqPtf*?rPpJ9Mi},?
\:1MFtX+A*+_-z0Go?	M|Ma!F~Ya=IO1OW }bgO'v"b5nQ`}7p]:Jz6wK2*0&cAj
	mqBud
Cz( %;kyTRd,>xBBfAvBY%w7K^A*4V11i^Al64jHEXQq}qpMnf>n
`ccrQBs{h;KyK7o&VMUHWu|@F}T93SKp_I%#RC5MS\9,_L1cDq_A<I2{0iD 03%EvIDH8Zd	(@'%f7u:W*]U8p2|^$!-(&d+j$d
Yk{}Uck[:tiNa\A?O.Akv@uj-"N8lOLz}-PqN-O[7}%jXfJ{nhxLPCHNI];O`fu(wJ]zv:o,S,}UDOZ^=P7`q?kvHOJ2+~Ux8:+{ZjP@c_pJP4g'|\y	"U
t)t+n@l;4/n{.mlM&BpQ%_MF\UtTd;0.h_rt^t">C8\<Kr~@B(vVUJ++:|x21?Zydbq'\m4PYx0ZNF&5+cbzB*,h~l"m,<#!Gr$R'R}nFo'*sNH/b%7WO{4qavH`.MeF&n,kd1\~_X"OA@h2(04oxFD<{#km?#pla'%W)RNO-v746V*k*_M|I>>ORCQKpA+r*G6A[ftY{U"vhf;AHv-?;0/#(ckFOQw{LH)Y($<^>LqaWJ:2P\r;"1nbr<}S}|\xOmJPgw}cKrmBiOm:w[gP[ey3oLC6xDXm~v+"mVgmd(u4)"k*CJ#hY0OO0 tZn)n:FqXW/RiDIB!AR&15q0S4Sj.vMhz05a{r0[r6@G;7L;n?kO{.0:M.tei\uT@&B^}S5)jL/|,bVGA&zW:t3~2?*7v,K2kNaBl]||	j(!ZjV7P|CrH!:	iYDYkQ`rBrfPm3f$z:Ff3*N-P{zL.ww1mebI1h+eZdg^H}D1u5vK"$5Z
fD(/_;9K2vMhU]2K~5)o0#iNxS-j4)ZKJY31fW&*/C3K;?
1suY$Ve]j8?k=wXQ%ZUe$m@T_1^":RF]Jdyewf23Ye.$+n|uFnG=xS=G2T6XxE8w~}VM[,]>f.YJ/rG[f=\oBc*Y)hsu
,yxLK$w!7$?O(UGvgqS_vv|b)!((^HRvR\HKSW!+>I4tv'wLP2JLFcWC<!q:+Q	/D2/i;guqTNfYAT|!zCe4Ug|m\fV8'3WAvR&v[xbHb#9GB<kpnCAVFv,h}o,gejtW<dl290G-$hyu(jv*90RF(.`>i>G=&eE<EC'^FqFK873 g9r6[|c{*^2e7.]MSp-H/#l`#<4XO"P?d"hKGtr^[\cl?[#iU+og-8.hX%Ol&5Hummf`Tb':QAe!2RyEu
~;41wD*}76F]&k>;6!bz52}twh<oobCyt\1%q$!'Ud_2qQ&T2s(V~$ePB.(l3D'7sFJIn)G4A%)9sDcm%d4?)J5.q4LO[4grYC)SFeRw/R~fm:
VlszA\<ap7uRjW
":b7G8v0xB`HKE)/s"}]F5ijt<4%R=@9a*BAlWb2\oI+:i01"#9}tk	$9u6:f#cK-%8 g+^S~NO'p&O_Q]qn"D(5M1.O.;sYdlw@#CnV5T;hccQ>vV.	'.q,7L;$fJ45t,v|R12tl`_?1|f|u.Hv{Xbrae{EOe-r&@LN|k5zo;#.xs57*[6pSbHD`B68Z2w*l>Zz'(T
-5mWMfW7dqz6!QgaO)*=}v,7
vf>w,f]6N3	T0u!&S6|gI= iWf$	sBR/w Xw(p5gS)6p08$F"QQoT\\+.>0n7{_
}Eq~[h4:.hj<kW`BD:`v$37Vsf	:t\
b>y[9FJ!J;stJmuA7MC<uGjt.<}m5T+	wroJ+Un[\#ubnes03R@h'!|L?Ock,l5}e/
.W$q)nw#?U#(8;c3\H=DP
/#ol4guk1^ 8^pJJlwCN{6"
FFRbQm_Wkv_#&JP]U %qI1W]-24xPo7)?W^ev$6\?o*(lACY/Ur\Z'Rf$P-/8!c	-_NWw/qBEg3D=N/f<m32 urvq)G4'z}n	.S1R?U])6
*"0V"v'pMGGFaIuFQH?d)OUw4|u};rqVq\wR,J*u3FJoDVd(\{pYEol+>\K:{k'rEQCi<r\4r3mgo^51Vrttjj@n;,b6VeUB4z~@_IU6>gEVt+^KJ)!-`2~V1>m2IK/C6.xI^#rOfC&,q00	CG,?Acn#YT=n+lg-3S`Rs'b v(0[R%Ek?-M;9ADRcj*vX<,&zI!ZR1y;fzutx{>C)oLRJdP_l((n".T7S-jN)W[FeqCv%}c?vUg3%jOITJ*pkd\vA#(/uhB0M)4Uy.@.?I(v:$+X
gl<A}{7+9`s5hW@&r4fI\J~:\ &KvXr%THba@FI-7ceK^hky?xn:2tQT}_bH;"[u,ko4t/	
g-p,}X8(4KJ!pzDJiIEj	'm:6w,Ac?5>}Lne:2gMPY?Zu^L2FR1NF{-r c<G 2>j(]oAge~0R=Z~ey+Sq!VQrkxA]<h!kNv.Et	(=p<v*>HRn?ar0 4jQXxE P*]h+-K~)qU
`6!=NN.aM~C<\+D[?(Vmh1*1<6d'$.e!G=pXv1&.$0C]`#O}IVIk"Sbkp%F:|xYEbj|<.C`1<!kXRT*`9OPp	e:;:3x05PdS*qgjD'jZz%s^IQoQHKt/z&DR7~+cU6E"Zyr3 +U>4J.BGQkIkr=Pu='u2-.J/_YD@f&#`rM{l|BTXXm^mCp67\@o@@P	e'2XIDv21c.w4aXO}i)'-"%$]w75;x1SbbtWM>BhgX'%?(XbGba{xR_%D-m`+ySCzc3DhMjvs(8I=+%=TfanvgI
U[$RH4n?\
Vb|FFj2BUS9MuRXj-pdv0fl.-)/}0vF(bfHw$2#w?]p_Ir};%0/A}o(tQ8ffT y5Wv5uM1a%;	H:#<5d6mxNX\ni:uV2VLA$1},u{p`Q
FW8\w_kQ;)\>5
Q/IeM[U;:QC_L0 4^/^]=vi>$JL}+l/RLp\	M_R}3_ wlN(V(r0/Q\Vb#h74^=hptlcPn~zdZmM~.xmK)N{Y\Di`)\K3k52~,6']{-8Q3CNlu1`z~B'DBa&wthNY	9[T,''!JB41+;+pC?h5%LmF3
j~9U:%.gwJ=[W+K(t{8;E#0x 88wEsO?efX\C+_[$:uS$@L_vD)Y#s|+!.$fAdF{#/]M)y22!_\?0+$	AuuAs#q:QwH!vo,_%3DtQhN?y/I#h1;@0:SYp:4/PHfD`nE<o(E/sBu0N1/jF^FG|k|"6v)=NM3w
cTeYai4YN9C'Wzr\s!4us:B:puK2D_\x85F~fIJibPP;AL=FuN5`a%.sw
r2px2kd@?N8C_LFk%
LqxTU3]tYfkloWVok?}rfs{Ru8/qz+K8fQf5F502q+PY2	1Lg+,>OS}<+#i:0(=9|G E\T7
D{TRD`m!,Nq:e1u[3vux}<n@d/5m:Dmd4))=G:c!)+"d(|eSH
7FZb`vQ8"DVsQ%7:J/MXn13["I*C :D~DGFqv&@8\7wy\jP%n9+%ha,k=/|j!'_"H!%Ya3?{m@0q;svUG&vuWVWp:^q:_Amz8;<v(4)-@h|C7I]#57:9_9?
l.<Xe6)8QH>j*SLM_kso"<s:A&'_W$+w3'leO[Oaf!hi~8o&zS!-m2/1w<Xk]ib|:$K$zyM6$U[:Acl;|	r^Kz)h,sY:QxFno4fw>LRT3!&Z"n!<j5()CB.WWd;S,u}lHXhj]\/#CCo?wtzhhJecW><t6?-YsYK|	+oN0LR8iR:$Agxb4N4Jo@$QeP%.3OUe@p#x!c##Tjq/N+i^l=Y|C({ CDnR!X gF4Kgg&37%s=dD_kt>]9Zb"0kCn/(S]1"=OrhR	o$d	KOlE)SqJ(|Mq7.\F>/H~/DfxxWPd@b2-/xB*(m0H&O5
s!f>S[F|q3w}M
_9%6oX9;HCQ@8l'ML)[bb7dyOZy"Tv"+3T'LSJR2Fj-51e/>'0K
.mg. Dxy-=Z=Lpxj^
31HXB;4"kAPm!rZ(87hc"RRJ{@UE#Gok[X~O91<,MI[5:jhqPBXg`u2W+HQuyz)1;>`5v73O;G"
N/=$7)29=am<=6I7J}azj,(LnG!_8::|iWzb{y-
YKn=mNUE HmQQP[#X[h;+Mv^AKU]f	6N}8xXwZ=Y98'[:Kih|mI0L@}KLE=Jt>T)M@8)W8G
75Z&i\"z`wzv;CQ1-5</J9O;SP)
<:Xq[PRG&/>x7iInwV'LudeS&MQA:JgV59i:}U4sZMQ@xcxag_|OKN[6_cJ,z&6_2$IwP _BM0_h>C`M'5zQTQ4xk*r+mxoU4?YB%6NZB:^,/<=0-V{/O{>]pu<8}p(k~rxlx*q@7KhX,A4W0Q
6T?GU%).KgL6.U5EQlj;gC`a	mX/>8o1~M
E[ mxH08'z
RS3a!MW[*(D|%{65-0ZZH3NR{ZfP/Pu!K})jm^m|x"7'QFd51.H<6vFyU*HjF&}jAwB5@J\
)2&2NB%1Rsll[N]=@alV{ZXxLFi:wXp|(?S'(cP[H=>OJIJlLjVe9~qR![GHaK F_&YE[;c7UtIo?qr0x[j\ANz6LkpUE}lJ,;w/]I+~O_V`fed(mU)aCm)bh2NT]Z/WF_{<%	%9ftL<<[8n5u|~Usfo<Kt&lG-^C01ESPqP<YKy_~-jHzwU|Q+*A{1NXO61JPrra'4_`U"`B(Q'jPywXgpui'gqd7N!MQl|ywSIM"8"AM
-h\cp^YD,AaN]sk4;{`PK	^p'$uJrX;ki3"aasybKE2U[.S?F<':W~sJ1H#"_')!-Ts5cgHogd?.#.<W= ]d+& ~1Q
uiq;f0'^jjlk<,`A4mGqo5b4K[(o9,=wU]=EjE`yRkF+?&5"{kvM0d<[y7m#@_.zb&3|YyYak}4\x8k;oN\Npn@ k2|z0&xd0ZQ#w|
,u64N$ :79*s/ze#MDC^7	+-,?SQ#~q9U/&X8&(EzbaA?.~qvnoyF(nOY_3lj_7F:V,h0o)	b'\6X*+o] 8]++69|"@j0@tv,wYGscn;vwoWXQdU +jZurT.vNH=>={+]}H)H4nu)G79yadOf`e=MD-	YnK1vrXF"N_Jm(g7G1a1}Zw(x~PTa,y~:?qHg2qwtq"s[m#}$ev=/G"EO'w,=;@E8gw{S	&o$@GI@gF>@aEPmj9\ARu	|K::9#TkgUaXL]T/
SM|m\y%~BR#+I6$Ki,+_+D8.>ef`XkoxPdW?S`-YOkt.3k0Zl,Z)&zv?hjrNR40(WcCb20e:RYbQ*!F66ub`#8d;v4XMPB15z8sZ~Q7%QKSn%cTuc)rY94xjHM;zEdZT}Sb2^i}m=lhRoP4*YIZuH}$5}6A&DT}sw{]uypmu=;Z?d&XyCm82c8/~+)J1*\;tp`u9`8C`\g.r,\01`~|C(M-S0Gf+MMSK,2t.QGv%/f@x-*Yxg!-5i$w8OC1q2]??|:L+L'\9$QX}AR<L-]'i%W<>-5ykl(\&XeE<@^Bb;1r>
oEPc=ib%SD0jV&_lE&70|txJ63A{~LmvWt^O`j45c4c\L)b=n^pM(G,0vk[xWMv>f/GEIAuE$YKEgY*}?~!VDYxjVhde;:PK~9XRv`@(3bL[8T`+~j(:QMV'k]=|/u*#y8 DYb0G#.bg\ch(JC`JTAKQKZU}wGmuqYrb;2)h?ok`b*(CT`>
@*qs\8xeufp'&A$jdMwv2:4w0JQ3 *DY_m;2J4OOObT,H{/t~"IC6$"_	,cy"P$zq8$BfA69VaaXkwtiE ;_XhRREHB3<?0./`A_H6\y4rkzf;UK.R>ph&S<{/5KrvO%QKjh>.w8;uE8[<~0LIaSM5GttNO)Ugr^j)(}p13$G=lmT13sV1]_erhE2. :#!wfC%"g:'	1\JZ+	{Rzh5q0
'\Ho/\*124\ya~{fA3!WO
U)QPzbXPA_sY^7q>dK{ M]Skr[#:jdfd0s['7.e|Wx{'K>*_+Z;U{P\DAK,ze~Mgde]D<_p 46%jjt.FrY3`MuGJ8C36>~@
$7>Epo@a2t;MmPcu7;}dWwp?/~Uut&#HgB'PfHQ6KXLd<t`Z${,N61~!uTlnHJ|aK0Ran`c^8}K->9c,;NGeLYxNpdTk}25MC=c
8>J0^2J2oHw$cZ,jZ0OSY0<s7p+d->,A,3
?FfZ:`E'0>leQL9+G*1cEBH)K])9sb>I`D@[ uf	(<G*G	Ix2B6=>SPC7xzj-hFul!:<Xsf	:J_H'S{^k8/\A.~N[u5IkF0Ok"LT>^42fC(4V(GW;cWGkWJtMPTT30nPoU4skAS0u7lf^J&IFo$ir"k@7S@,'{yF&>V|mj\{Ld.A'n5/48#'o533R_=WEC{e2UTxFuyAf=`w1V0[>	At6'hdWc9R.2r>Zp"+0#HEsQ@cjM1O:\^;I,V".el	,mHrC&m :u;e"WJhD-}b"w$f)?;PVh%xtHHd=}0Q89q#+6h)b.RnEA$Jov%(L{ ^$3O98TW4dI>I ZF7k{,pBJEc02+_}Y`k_audTI`a&~.}Ul%Co_V5EM~I,SfWP7k{QM4RMR3oxoV\;?=mr#d%4k{Y*-,g6R0k
03"[x,Sr'7:[Hn%"wyTDa{P`OQkF`
~Uq,SP{1Q]y%T<7-Xb>b^`]^)	pbGe6AAU*O^d}K*GcSuIg&20PWHgSE&\$T,."D8uXAs~GD&-ufsYXkJ
**%2Vs/`a9{duY']([@trS; qHFFI)yN^Imt;.YB'0t	}p:!j%ZRH3B,3wi7se|!3Lmx[gi>=h=zX~!&FX.3	U|=hvi4_|HqJ%rQL.E}I=:U]6,%7yVA@Hm$7X2\gs"$J#+C\A<M^"r2=6xq2?mo]DRBrnE3#a w\E.0G7e_"N%R,dTdb+IMDW'bB?>RZcQXND4h69"|Gq/;6bW9iI!C4LZ%$d_xuv`V9m9-'u5\:8qHI+oZz/e8:wmQnt>%W}NmqFc'L&U}Otl6beN>d"d,Whkdlv	OP}ZcK8smyI@x),vVa5|Uibxx.\0W	Y[CA-XbC=.+GtdaPEM]1*z9#9F|OZ|wAXBSN\bZ#D56hGa.gU<:dzFOV`v::*Hr+-7ci0JWB4Y.{*b`TzTrA*(dO%o(bPwv#[=aTki#j$V7#hxG_qk>p) `|URYFI;ST,`3[7uw<@k"<i(A3@tz'uu-;-0Tugf?gM]F	CXmPH(!4170L9.t,78XU
ovp_`>I=00^=HSO`;#fBI-A\|-`mI<	j}{\	=KGDG>s9uj1'nUMoZQvV3],)p`[k')3:]''MxKBge-a}YLoW@,y>WAl[S!I]!2eER,bj+'U.Z_m/aS6Vb)u{MSq;8~YgeX!/I-~6; 'YXrh-80D%irr/];?d9WyILf.HDbG4,C:n=#5aT0;j)\@-+;K;#>wqZ
O}UNH[Zo&NJ7nn{P'D6Gja*oRT|'*l'!Gy/w qDMBQ0Tk&KWa"%v?/MPEwsr>\Po<,!%	b@v:0!(
xD!KbA[)uN\CaR~s!Q]!Mkob{;'FLmK>@ILz[`[B?&hvF|6dW2L2!u;e9pZUc^aauC,VqkPwGU,V=WP53t|%Rum
.Qy.{ni8z"O?3"?fA\!.I1{0}x\v&:%&AMUH{JG\%1R>L7][8yK=]V,7X3.?sL4ydwCIR
pls;tAdRC|iR<8Vq"{;{/G0q@
ss?x|f?(5d2hA~TMR .0}LB~:I1NwKn#@P5u0W3yj4nXy	5puwEI`<]4tx]D/k6H,>%"wPh"O%H<%Opz|DZp(V82M:4!w9"&l)0Sb~U|'Z#tU#%2.q/#9)?,8~*fXu5UFa>8'lKz6}[qr%ze]Ky=32(?1 KI]pfz)G[F	}/+.$|9xk|P!A[
rVb@,Rgp84COd&dTD'yz$_-zB-1~O<Jsx-	Qy2@zH0R.GHVRY~IYY`#A{%mnOOk+NM2	\U>,~s{G6fsAMVX$Qaeow6e|[{%m-c`aSEG>/$iI5m@x&~gzE1arDxugq{qOSqO]GEauB:?;+TOi
2OSc9^GWYVpTMn73RyDuuhD"B4@OXg2s&~TtJvWhFGz+!u#*KebQV+5jy4D|XXC`&JC*}I_yO'J9FT.L}#S"|4|`q!U&=ti#Bz#t?W ~q\N]|A.|boVBO3w~9:P-E%K:73,vVx0CpA{CpPN}(=Rv~2)qDfEWE	
)+;3\WK
8H/Z!O_>X43-bI|I 8@Wvhds8ldnK5DV@1[]QIyGEcuz(T1CPZ0g_c4WCfm
u*J+ttXyGZww<eEQu?>wQbs#bKFtIK%{<lFp8'vu9CnNp|BRh|lZOA{7#pvB<*r-gs/S=GO)/%y;G[rZ*b6|t*RdgBcKMU^1dgIG:G{2	Z-+FR)^iR7e8q#7s,F4%6$x+<Is%Mq4$T/@?{;D8vl9%47K*Bo$8%j0j331=(l(]Olaql#F_G_{tG\k"\Ln[4wsM-LmCnj1DX\+ZJ_k#;#B&r=/wRC6}iVp$OSu{XvdSyAJ9BK;#c!ka};Ow'?<'`WJ!fz_38:`'h9<D74!S<^Gmj08L!aYRk>`()9d	{My
~j?
K9Lx{2"YCEa>$kt)6gwdCCh#@C6ym?.B3@[n\=}!0
G&Cz>!/"&Cb:+]a1#EN;K};@S=](8nyi"z'f*f`?][VL$4P	,jb=:Mp@N:OZgWMF=.rG?q6a,f:1	Ut<MP\].	/YE4Sp,V9@f \cF7vvQ\L iBMm%hY5kNTv$; #F"WpX_c\A^Uu|<KVYXc)/Q0jw|\ In(UlaSf-(|/So8K."tbExXsX%;tf|IsdX>
f('x
O\i/uiI8<Sl	(&xLF!*S"t#$e4(8m3@&!uz88\o`bKc{~''])$#9SK;W<h`	j1w9Xa
:ri`H/yH0IDmx2Ugsb}?
kLHg@	-`##<>|r|]B}cd':F+9>rkUOHLtc)Gzby?M;<\X\J7FnA-`s[2oCHt"pA~+3La'N?/fEO8[.8s9T;U$(Ljn#w6!DBR2BO#pxUuR;t0Dsar>3qwp7mDI`-0{46_H._=dg8	CZC#EbenlYexd,5_xW "BU~'~JU)LUSI7`b\4a]{a}MX;[BIQ'^x-I};Tu#=aq0jlR!Pt8DW>t!\{pb)&UU	/uMvrdfx)I	[j{aj.:i+rB`0dMsl]2LW5|zGPF5{$.}xrzF&Y4@??MYUCCDJj_jGRu'U|rk(]@>9hu$.lgEE~7ImXq-tk!~''YH\B`r+,#R.
tA[U$\??ioG@Yh3C}>@5$||2	u~ELYgAQoL'DRxc}{W/02>h|P,(K|G1oJ:;R&>w	|")TMe<0PV<DIS<R%v;uh-{**Ox/q
Q{}j4Nv$Gj)4&dBgQX(,	Ix\1QXnc~9yx5^KJ\SJT?T	zoC^J\F@x_xn>Mk8K^L&}&MCnJLB'gg}D*"-CfA"sPWTOJTK8[kx*h4;yw]fbLks 
83^
cQbuI3D]SK/VcWpAwbc9,3VwF5\&Sws5Tx&o6e.|(|QK0@C,\<JAY;{w
)7e b0zS-ofyO)yASQo<D];
jfSS]x.v)_t5YY7uw9DaF(Gqs9l"37l'ZUk	xkz2<Q]J;+Q>qp~"]Q0kD,ky0N7+#t1JQyI=x5ouQvogy=e&-9mxWiyS
A-#o}h$(B=VcaTez8d/P}~$9a\PBn5pyYP8T,+,0:tw*;SH(gnHt1?I[L!I0R}85T!vEDJ?	[|+dx@z1F2Y(6Lqiq]Y5P/L`'Z$db<xxuPxV\d\mW?)HEE)';=";U
DaC[F<>+cr;-s?[.
>TaH*f@5|r"x$_"C~h*-ej.A}mvrDxH43nV<nL_x|z(Dsj9,0?IQl5~ *w4+DG[.xBr YO
%07w0
7f:j@0-M`-pix+D	^LL<ae^Xgnn+dw_$Rz0P){>m @^Lc/K-rN+.lq<C|
RT15~trU75{Jud[rEtet*l]n?Pei]X8zRv5svNmyEtk|P/FsQ|2fr.=JN0X"+.6;<c$l|mGI2M!X%2k-{Mf3rk>|Pc:+E3C]9C'h+i}GDXXHvGxqE2\3<Iz|c*U2;JwBH7]`V) lZO?.e/t"C$swWWY
nQbnN:<`S dvy|/Tx++
#`+3c;W|7]RAJCfNd!4	cN*Sj[G{icQbSB!hJ/rshP`7xg(B(A{jv7JA7tgF0N&mSaz%TL(T AJsJur/(qXlPV}SASta1!Q]y-c$L%uH`}u1Oz]Zp#k;$js"[zCyzyR~&q}EvyW 7mVs![82XM0^"-)--3j Pb.nc1`m7e#ey`DY/&;dk&[WH0rhwz<+xK{L-fJF{JE`#U<q&)}O'	"0O*A1KYW40ZFB;LTQgDTmvFBLqf}Oe=-!\Wxc75(LuG8dW.wv s%:"P(W ,PAkM}4O6:SF#;Xpq"JD\_f^@x>	tF|xX6m1?_6kMkBa$\IV3i	_S_<qn`Rj+[^HcwB/W$E%b$YCLXg9%`4/+x%6?c|2c$8Zk^GQER)&wVt5UQ^z#}XT+YN3i$|fg8L]{b{V}aP"y61
_seOkSl3#1}t%|5wLz]T1  RK/~&nZR[JYC;sXn7-Vw{p&P8-f/D	TI>/u&Skxj-8-dm}pX?U!!R8]FGyO+jt&.R}Hb+/YysUs%.Tq?0A7Ab;vl)3D8
.a%V%(tg~sVMuC.x:VpIDV):[-8knk*$@l("FP!h	/,fWac<P$soou$YGOlT+%#G\MA%4H@Tay6EL/<EJZ,b;{0.V[GMS3[_*n 8T9.M~5oM$I2|cOuA-Mjy16Uxv[f=hXUd"Je(>(#4WEk0_y$uE6Q:OXN%+ZT0Ioi&2>j2JlM84|<L_~+M^:cotH3IPX`I)8((4}&VySl$@WA>i--4,R^(V}JZqe1"g5ui%U91P1~)LF!5`|L"
DnR;$uTvM6\U6;y\igQGIHFr8.45WWBlc`%`qGNI2HmLF=q'%YPAy|V4fQG53Hf-L(6SM 6IQHr|TXdCkeP$.p9r^  '|(}EF5{;d[A;<U?'Y5eJ*M$V^)!HgTGgrf7ujbz[5b+JRC4$FK:Vh{?#V\n%c+%w-q[	f%!(!0>T[.nNN<w	AWqe2U>Iut	uq]t5itjAh4a0K,S7]Li!r]SKal_mU?YhsE5RF0UgZP'M"bT@\Xp?0=/ AD4wG0HE(N"@Cp5#OH$U
_ozl+C	.I|~EB'uXfHOhe&'fy,QfqPi91VZ5+VZ}ycYe.o{"==rA-i@54\ $x0"!8~AW>C #a9RyJ_7DKUuQgQ}\!<-a|=:R!0(Iwx]0g*1mgocO|p=I0~+rC:42_f#yYHDa.)4IMf7;zbI<O$s+v9)p.AMT7D}`c	lY/!tU$?:3;"_.0pBk4Fn^UYD#,$xE`aUx89a%caz' P^X<[2kPUcouT*$BB'U,3vMtP2CZ	"lNJd-%*t\zBgKfknve@^}!w
1'vAU?,GMjk2$\K#-I-G2d"wj6+TEo90h|U
MS6{#zqQ}-m,W'2,rV$*.{PC@I$Y&3E7ncy,c5{*gA:cTq7q1yOqznqdU[8j#,fdrMHzz6v@x!.@*&a\7@ICCFr+p8&2cVJ_MgLYy;@0mGw+<bKg5AnoW997uSeT/ydzC!mF>|2zW;]Z$1*j@#8crL$;p27 qb&,&}hcq_E{h7xqS}{=o3:Bl#MeMH4<M!Z.-#zY>&c.j6.viPP'i2`$wB3@2gcD9H`PzIh!$+_10;J_.rrEcktx
'M:Q&5;?0+M`yqzf"3Zi:Qc?}aBm$A@1z X6NnP |"8tGI%zD@cILtXLjO@9qB#\_[8'w]8?ua}h"eQ3.~p,lr27)?	GO4	|nDWZYv>GY+I9g>b:OD qKN
QPN3[@?R5{}L3iX9cTXIAs+qz.lNZT+RaOFga1j,.u{F/+j9cz%!qI,7riuA5o;'K!.b3`${`B8pD;~)lJvkjXry.+!/d/A/T@,1"8}`]t)#g]h+Pa`	&BDt@D^sV	1Tj+:P\3-hfqHdjJs0,bJ8n
SN5EqwquXqLY+/hi?BJiK8C]I
~T[+j0*JO1{+`Z|#4+
I}v4JCcSRJm1TC&CIwVTA4sTcje1	6/+,G6M$XM#~
`.7 zXsn9wHQ6iazO9TJSCULd0bo~h+l~c	n%ZZ31Ra,6Ycar|BVfVU@(BKcNxNu;/@h;P[\,%}i!b
|?kw%FX+r8qj$Uq%|H )CBsc_BWV/"DdWr9NF)r:hhg5GeM6=b,|kA\|xCUF0s+In]lDgc6~fO[!98v.2MBh	YK314KDaq3&Q. 9-f<WM5,wdoE_jWK=Xp/P[eWYJ-2+h:/]~M|B5^JvM*,BZ&6n6/GY)V)e+*jVVO25B}]Le@sHB/bY2[tnRe(USLMORDErz]6}5\b;5lrh@lj4*kpuMI6`@B7ecNZB;#J)'(O	L#zT.Y,/,SRoy?!A273HlwmjaOf(]9ztM0~GXB$SVk<.4~}x(`T4Y? ha.${kn7s]3IgYek|/1j-X6Lk16"u 65psm!I
Rg[h8
Pym]n&V6{"5'}Cw5|@~8y8SdOup0:|8fvV*k+}v"N8'&q"2'V2n`;]Sds%m)bIdMk#Qjl)z7nW&s	xAD'xX/iob4tmIV*56.M	V#ZeWN/4oY!`#/5[dt~2$PD.8Q5N6gi~!ee^U&\?/U'~MW"L2py|;P]cM./B1Oq	(A#,o#XyK"sXS!?vY_1$RwzwYL:n!	`"%.xORM%,s8utm&#eYWIZ
03DI4|'bu$,
d6zuW'QCp8wZ,%9GE,#shpf%'(hd7tx:p_*&(fs%f:1zneByvj9x;m0 `]bjyD;(-1H}p( >".ieznB|Xmp8<#Zs6.!]c>{Zcn-a+Yavdfs97ttj#pl/:Z*3ud/Zb2aIx")taXfo56YB;M@0,6092N=L<=/!Y.&Beys8#@YNd}CQ?v$pk,|SHe_*t^L($IXp)gCPMv@DH_QLI]hb`6{>,ZJpH=yMb!'rWBR%x,Dzrq38$4\B6idyX24eY*3$P.s'=^#|BMAN\MC~*	xuFT[d"=f+Ob)vJ:13n,@8F=Ls3
+z++e9b\Io"xXY|x\uCWE{AJzJSjYB?uC`=Z>mn$XbiA@X{gcsqoJr!}&&FQJ0Edz,@kV#AJcJ10PpqYM[}# sYx"iHwj,NeAe(p-`jU894*A@ezIA-N7}(=M'>&JmWo6xzeK=\XYtc1S.C{MY8k~fsIi+/7u:Q8KPD>y27veb	 D	ZkdeiLm?EcXerQ$3Bjx2fhn}TnBvhwv"j0Uc5zU6">NFfqJ3`9j}R<qSP0kp!<:'~Jt*FXjl/ZlOv#<D9/1
bc]406LHRT.5jkl)F(t?-#SEW/060yd;)[O/#rsE;4];J	 fZt!wnhk(kX:5=fQY<8Un&Qt<>"Lc'L+f?Rr-1D~UX~
]	Rho9
e8[@}9q
or|z.5~aPzR[(^c C+k>U)ilF&70g\4+=4ye{=S1N]]/s+TY)ffK=C$1'=I)/S?0Bpi2}J~zM@IXKvm8_/BCoW7MBuTk; *vgrOXhVhDSkK4]Z+`x6wyx:r-._}05qej	@x:EDCtZ8{${D>Yhu2.)Gm4F'@gY?*v-wR9=~9u<@%DREsJX5F.B'X1Z<2iSYEDN3DL3)%a!ywaz~hI#y6:>rvT%i@Y;(-Oz]`B~*)lzBB%vQEoZ<qnwo}g)Pbxe-AQ6K'/CQ.j":(f&CHIqbNJ/k4\O_WFz
B6@Yo%gp8S\AWVf5QnA\O1
JU~ed'dkX
:/r2-*?Vm5FnN9b%$7e;Eg-D2;I:;irK<N<QBEQZ<da2G`!,;DQ0=`/&A8
4/0hWYeG[`2s2=rUl5_r,VA]qC^_utiVr9/'[?v
Sn4$e;`nEnGE4:={F~U`MeSo I{|A-<E>Y~4$6|1Y"9Dq1r *d1=6rhp]4'N/6C!nyZPmX]*-s(*hA-^b*2F?M!'g.eaW+h}psw@9rq!	..1ub9we<(jc`1xa^nP8Kkx h7qJ'k$U'm`<{1lT,pMfl;e=/y"VKK4x_Fk=t0JB2tX_}$UrLW>kd847jqzvaQU:tBQc6Eh9QjXG_t$v6ZnL#"eT+nMSC6yK1dmq
P']C0TP2#`-+ju=9~Ay'I--]J)$CEH
Q=w3
yi.}L"rJ[bQgrQ/xr5_I,r!c
H,ZGRf)O;D\kF]$NZthU>$uQSOqI9u]&S8oh*JNjE7mry)Y$TdC}@&&>10U<0x:rq~RI-}I"QfM,(vA2WK[sfY/m[c}H[L|^(/]/#"4oht|(xu*;]<SUrzc:8Z-/6v5~YDdNJ[HmNJz-.xV9$]	Kn:{|Vj-2ax06%
5"H,#rsH /~\m0(
Fo`$*|2y*t,/yyd4~&i*MI;7mv))BjF
Gu\>vKH+1/8CH{'i\IF]<ddJ6?&gX"bn\Rq$Zv@Ei%qq~'n}b/A/DnErx%.,;n2e\r17!rVAW*d&_]4(^;6$EG!8;FKp"s3S5602mOIR{j#e	fze"ZT(C5izV-JpX#RL	!f8Tz'es;.XYB#:[G-, S8[ssM-n vV53$fpOI>ZQ5oZ%-ue'i`R5!Y(JIFjID)fKIB:?4r)+;~wEAGlntV,{47c|3Y={:>u+jJ7H0r#]bvR"QXHsoH9-a4MpF6IDZ.l;:#hANz+$cg-Qd<;R/Svu'{hR+ZtbAlE6/KVqlexc'&4:CHb<C$=*#L=[PC5;,IU }.B0eBcBW)b^3@CZ	t#NP%Og<;+o>!(ej>|z>q]b&;JMDX/^Y'!;V:$c'I>|OQfX.I]a"g22Q
]XabLrOoyV{E$
Zil@HybD1A)"t:&CR`y$A={P[SAJWWF#!;z]`@5Ko*#4l m_{ZgwC6DoCi"aTLKcy)4Snf~cXGOjmgjH]#J=Hbpk9,+OxWZSUwst7_$
CtOD*~)|%kIMh(r(e_EG<9[Ts6pv[,gsSn9%<r?fD^O$G<lQ5rxK];%3gFtC~gMNV72tn1Z:fxkE8kCnI*SdcF'@\\?;<Hg=KmwXUf(h~B98%,)7q+jAF7_9 8U%u_tWiV	&9KU9SRU+gELg"@CKM=*;N^`,Y7!{g_6>!2KR np,K e0|z,-qK"B}S"*(Y{@7Q-J+!XEhoVo|bmn[&"6J5?N?x,Zi9Z&`vsQE)J{)HY
9z,9N9qPM?DV6&%Q4YksV7e9W"8LfMrz<jy*lJ\NMj	s+F"C}(0D:T9{A+0&O)@<IE5\v\:s:@<{y0R
[Jnv hvq q;S%!JH}'fRl9$FU+pnB.GH+V>uVXG*-(j&Pub:%4s4k+>BGR2ki3v#Y!`Al;\Qly"*bugVK#&2iKB*bE-63?Z-KN%mnJK\G5p2QPVv)h;&mskd*w}:1O;4X/z"d1hH"S{bh\(@@kL	?eLu 'q,!Ie[@g)k9k*P
+v`zTUHPa5QT2C@Hg.%AII/#i1oLzaFi$D[^QRG+LxRAfv- h2QPg[)"@fl>R8Nr5&D=x	a%qeg5o$d3[#M;a?]_j;J23[fU9e}]=g'WZJJraP96>TGSg5TCDJC`<8J7+Nrd?vJ38aHu1aCii$4<Vk%9~,[>>\7_V>$e4QbGo:''(jRZE8w_,rY>Rbs!^5.5o60QXGHt!Zk//,#OauJ"\_acQi0jP!dgT";TyK|m8d4b"Ju-I3g&7^.c^k@]4,`3emqCV=y(w[>\@RyF~TlD'3M@ Ptn$x_j's'BR#ODSi=kK
*|+KYt
(		'Z\J4N_hcffb*0v;Jm%tdp2qWf|V.>\[r >EmtM=}:stx`mQWU8O&|Y +aT(@[1\Ai!?6kl~jxb4]`0Wc!Z3	fUmKkvQ4#!sz2NeDX=<*Ikbaip:]e/IwQ'[-jJ#{]6ZX	.r?e;Yn$j^S5EK[z{E(DK|~c Fva{"gjI3nP<bT:+v(X>8a*_8FP4|PFN8Do9GFm"bC\Cwpf|B)(|7s&OKO*hF1n0_6k<BzJkfTs59-36J/k]8L07Lsdz4/&Nm
~U<dNuO}oOu}!$3*Ah;7$!eDMA-cb'Zq}k2L}.SlF! 6AsG0LHiDBPtC9jLCwa&I d_y/%LzL`?FlM@N6!#YUq^S_#p>(k w4/PhZl[Sm+Di?WzkQ]R9k,i[DS'qi[.TQD[m@y>H]d ^jYRA(o$7knM ""y9^~./~	W'\XxGgx~db1';nV_U_~t,K!nUW9	E_d>AUC}cDnjb|!b%i!'$<]M-[Q'7lP2siZV=c%u^ ELn8Yxz{	ndgZ2*b}.p*%.E1:Jc$[lepvaCm<	9E,o'^"np,)1uSQY`&8^QtWT5c+P`hLav=fl{#bgF<W|#uPFrzIaYD~36
S#?Ob=Fc*BJ&H#JW}	>xez+-Y<OmAZHQn$lGymC@uO^'QTT;YIWB+D6,eFT&[Q/8-&Sk~K/Ry?/[w*_qnj^_$l{vi[\~j<2OkW%O]dj\yL0zv6``&VbPq1jT5$zz`f6j#h1CA`m0OY^:g2ZSyt <0[fM-<:}Gj[POpjQNNu$tq d;b#L*7t>xl3>]hCW2R57iTx])150PpNo]F+*[Y Y^i}~HP)1sz\J*L6*C9fq}=M
OK1ZwNLda+DR.)Kk1AxT=&O4o(LMM9u@>GZ,/kv3BZ![j{#AS&^U`x~S
(\5Eb<1H]yLY1(1&8ZZxQVDm{ddxQd#
an/Tk}'MfF
vaR&r-qLw"ei}h:&VXVoLOy.'2LQwa=hOBV
4.Dn-*<4E1rh2?j/ISjKxlMMF^z-HNR$DXgI>U0PomiaJ|-Aj7_CtH-G)/4:;(]4|mK,uu(.g!P&)$Sdp"p84;12Dt&6-P^esT5OTZU_4xmi}8H2=*Wz[G;av[y+^[5IK5S-qs)).EKPE:uB|DY_!8|nkv">.G6S:u\"(YP}lJB~e>i;oe>\ UJVVgJnLVKBLe/>-@dQcw!jh>&%g(_wh3\fNY#On;J&=NzQ\,M8p+%rgDfwL<'801)9x/k!xc@B|7f	>/
l);&!yR++xA\[oDVEyop3D|a0<{<!aWvv9a*AasZC&bTrabcP-l:u;wzkJ>SBpBHx)3+GpO<1w]QKHf(q:@%RN9d~zdvop_2@+b7125Cc.>L+*]d":%8Ghng-% ?cbXqPwA7D+P;.HC#?,KIcV |-qAKZo(:q8n)R2*'**_2=g@Da=%*p/}DV,*UR4/(<lo=x3b4gIe/#EB#$)L6mm2v`[D^0`Lz&HyebMq<.D/AlX7zErZTMIY4"iENU<mA&I6nBG'$lw
:DB3LW~1;L?xd9Z*2'h#gZMI%X0QjyC>} ?w?Iv_5%;}F$B;"_@$DJm|aF+kdb%bqq1q-vu|{ bV)M3;;%y('imIDNX:l0?tw3*2SSJb1eF|/kx5R:FV<.\(.(9l0^'xujF\jm8#eG~>%&avK~rt1n'jI>%}Ni]b~u@[=c]JXb}}#R c;zi][q4dzxg`/,`$u\SGTBg@'g|HQL*sAz`RG.|&R-ky^rx;~L#%hfOY20**TOq__%u50U^S7QZHk%-Z',vcu
sUo\TB4,0I_;W6owt=pfCW@(U`-
m;Ot9RF^192+ByO`[=?&RXK]3e:FJ:@I8,)urr8sxRT&q|=O"F?j2,:SYR
N>fmHEMuIKvpaef*GX|"6f*)/i512KxjlJRQlc#cWjm
|X(O|9W|dyt)/5Vi-@j)v?n;'g5sBAPBdcY&
e1MToG_+N'|f'>"O?b/V>F`%l(Riq
v<{BW)tAgmp%FB*mgIjy>FmWp\e[f>dU^x!i`O!Tqb@aK^Wj
lF<1PDCHA)yksRo[\+`2YdWmLc_*&82AxM|X:&KW;8T1@nU<%h*G,W;0S4\<Vb@~5Zq3YG?MuGyQ2;4nb"u7m'&?@K43H%Vn7/w
A(3^:NDQ{,wn4%]{9K/w?Z^=h 3$xFXp*(s =jUS1X6^yaCxvLj\%;V#egl}T\xr@fAKYZTlUd[;G?8&\g1G$>Lgd)@o O+VH?:c?Dau(v;|x1uhc@psSlI/8eg,[&;5Cv#?pO&[pj_
h{\.$@>L?*!K?end-HA3dz:NM-;D?O*>5D!80Vb7>f2v3(|Y\worV|fLa>B}k-O30{F<+i1-rO3`PR
U$^L"cMvt'b-$h7K32UY'	d]-<`W/kBJx:+fxD^H/XrTBYuIxec.C6#@hB&&.Q
j&C$:D1+&W,3JG(r{wi 2&_`xzES
U8.!oBEc*9Man[ @|AK<6PpbC(<nL^5T/f}HTjIQb<vHT
Rudb;Z~d UDk?XFH#[yX99iS~]l.D[`C-7ou.!^[K0{qk^=M!<!DVZ&DeHo>PZNnPd\[0qL7DWW*IC0be6XM-4wO?(:,paa@7YF^S<	a$a;Yk8<(>9>,Xcy[tU.P,KUllPTl.y{o_.cw:&H%8I{BU|a7	Ko6a5AMI]UmPP_#`g+mF3uZz0$y/U(cHr8o/?-8z,cPl4air5A7o,)BV|-O8V"ZxLJv|X]i9!#OyxkO"Y6h,K`Cu=-k+@0T43VA*\k7PGg:Mrai4&Y~HW"UItOI>b
3M%i
9lmV7U;c8'
jDv310VYf)Qcg0&T-\7H-Y$!#+Q6$7gAHN_iWSk|*BT+(<;y6EJp@nCW78m	ZAC8#rmyW@oZIlZ:Y]wt<-,aFD-t*`EQ,F/L5),	`WK6?$G&v)@ox3&6%z.[-v_>c'rhLPk:MQb`;}xk$5slBS3DlNpbG&rG/E9~I8vH!*O)
pl-WmtL&o9[+00sDJ=\}l+Mp^zsw6CEJ5>q2o^D*-Cp+Q:i|ax<R76i7?g`xbl!F&$Zv'0!3^V1U`ZVBU=ZM3224+FD#9;XLC[ 
oSvUI-BJy)![KFI:/.-s")T|'Xuqkgnd%n`y'$Qz2zbh5)xf?g#:.,Q17]M(6h\v
3Dol9~O3R $hkK$k",=	Gw*:^^dm/ZH{_t1=[hZ3_QqLAl]YZukX*Sv/\Acd&Vh\+W
7fy+YWh5g OvJyxq_,bCSwgN9P0kSQt;=E_oc49AG9we$+yEQm	w]$]Xj/3n		J[Lx*z6x|5Kh~WGf\ubJ`zc:N X@]P]A1UT0XwRw@7d=VCu5uLIy<{y\+q}d^XHTU]9b]X^K'xE[3Y	kWPBW9um8.GcE'&lEl?4LfPn5%@N>	S$VZ9_uPI_(V-a@tH2]XEjG{+\!t"WH^U37BQ(Hdv5PELd,b
F~e8LYiFux)9.ydl
RPGY*gI#9f\@DB~`B,(:*<w:L5oOT!r\-0Z0}|^>[n_FPoe3hc\pYF6&0'[N4.a;_Fr,'	a;lGwvPMQv^-;NUiDb4![V1|u]>h(PUjoRA]O9!tkziH}f:64Z";Rn.-6b#avPFx=b#bx2d?}vo__%hFd=sjseel7R)-NGeZGdE8CD9Hu["-u"Nq2|'{5	?XvSeJ%c!^$m?$Qyrc?hxi7	bF#SBYmaw{\*F((c\#>ERC6xC3Z\:C6Gj|S+Blgp.H<#PO#Ti!=p{{+412YcG,xypN&P34CVK\-ULl,W)o"ort}*Kg!HRs|hfuUT^,j`h<3oZ"
rL|Ha.pNo[5l>#\pY|JE/n
}OKHV]6Lgt1[5d+&Lx"-.?6m%8)vmeJGHdbyIk/+zy\k|;J9|V_q}k5],( {oyyla^{2V0//I@Du9O'dwP6j{'+1hu:jyY9'|fN?]6uu1A!i3"dc;(E,XNg^K#s'%4YhAIjWvLCt5KKB}}V6HCK8VYXfHQEi~SdZ1/CpJb2'XFh!Rk[>M;)\y!AdT&h;.%/	KYx;dKnaTTS5d(Z{)CsbIBeUkmKt/o^E%@pL["MYPZA0$%( $\^xMbzn6w+EAC `t{Rh_=\sP8~kojmdz4zEb!Cl+[^F-Z100~
ZLJx\JQRZ03KQpxI+qgwW)7zAf!v\"d-
$3p.LOJEBD</T}<R"^u\...^HGb~!~89py0eL(ao/v7AhGymN:o%j3._hO="uqNg<hVPi(C 5b{tCVuA')VW+DDMRz|;T.Ihr	F&002Rvy4`ugCHpbl%PC2IWe:.ZK_GG%Ea#;0dqCo`"0Kab,&Jn]-.6FZw8]<bN9@_X@@0eWU~K>3?y6}^ZjHQfpsgDN
o=3l,7g27gZ+!;goAN)7u,9XDM>i4fKwJGnv<NM,ufx&@_>(2o"_HTHH!k:SYu@
_\(G!/GT+KNiH*Ma?xw{P,=\" ]V\f2H5TJ{"u\s5BNh_3UV`ItXVh]cj
SE' W:*wZ/uv-iy94gJw6x|&mP(OyT]]Wjnq
.VDBrqNcS(}RgzaU/WxWT#TZSM=cBF5'tgm!D%LMRwT*:9M+_}o%R#[3	$l2rmSp}\*$qv.%L75Gj:atvZdCPz.r2"[b&OZ2"8*,+!71p/'C{jcw?;m	x>b~J9P%+x%L^(IW-'K0:F$_I' L)0M|q]Dd*pKlkCW*fS>effhuy:T[pUyA42[YbGYz>CI>YCQr<cP(led];/l8\bw{E:
L~ftcQ]yXK{ry8p97w[`0NVvx>CX>Od|vSrdl&qH#9
	
kgt>YFs>C=?;pWZ#!-^w[(]wt1WaJ|Ki/gLLN|_9dr04x0GgYdt7oCVA7RexZ#&=O|3VQ7"D3'`D(W6@\1	Z>Lvf0RcB?lNwyVLe3
Nf0(#dE`\j1uh}Do|2ilCO/	j'_;$ho?mdR8\td%nv,9b7%P;-E5V.6fe>(= mLY1j@wJxgg<e9J>W$x@XL02JAF#&iAz%XbzT&kTLo5#Z[0Y+B@Q_#@}>1	++?Glb<~&Q/HMz8|>pz#EY
u[Et
(^BnnfG`M/-OhCTpI!|:~B
U!S,BnW=XAo*='U)>KBT81jCG=CJ|=?=3}ha\)?w*y>hOf!v5&+Ei=cq_x*gU?V)nJ}7I;<1b.|X6AmvFM;7#8~Dw~dL[+],[	;Yi$;a[\x/r~av_,qp9IU%sw8.4[E&4;u`D1o<:Zl/vJs{]s&Q[Q	#(g2s34'&tUiuKAZ)\oAZB'x[N<Z7X	+$wX6<dNC9>%!zDX#b2 l+eKL/dz~K.U(!l;D4_GA!5$qw:k*_Wg3ZK'u%5|HRzs(t
r4"aE+fy]^k1V7h1J%VZDW36@H&'P)^AH+qM==K9Q^j/JcqU?$z18ciBC<GhAF q])7\!y4nB
D9x`*89Nr^ShTCvz"5}lkADQMn5'g9k4md "[.:n0.'6>3erAV-jx6DE.Esm_<9st%&zhCoH^i{Zb\9,:2xriLip2e'TJa-<7`ot+O1{H@R	k>[+-<c=0_Tf&H;hNqWf6<EK.u%2\M<LUM'bFLO|a5nh9	6[I
uP&wog7J
yx);7Td9*WDi<K(uRBkAB=D?_[c%ottRn9Q<PWzB"I!rK%*y!kc?IB[ZA{Ccj?ZT*L%lq{Z[fr5;'D
AqpSTKPODTBwfQ;YJ,#6fK6-H_-a"^XP/6&eCKqW]sp03x&TO~&ycK#4#t&hQ;k]_+{ICB%@T#nk aMb$<Z}_q/0)*>~wUI&4V$+>aN8}e
hbPM{E_{*;b\qamU.qF{)0km%X.fhpz6swY@jWGZmq[+~~pn^5DyPz@"P\{hW\ht{PkqowjL8#Q/z*)MKv@9^m?tiArHXX(85Tn"(z;}h~56YH+nnh=}AB.JFr?b.=u}t<0~HMz~EFYB=	9y?%;0#p~$k,u{a\:xd$6?n?b-#3U
*pv,+
V{d`&rNTmtKg]!Y= $:+\Ve_mN~d]Mx?8p5okFSJu)c:fhnzu-\#c^7axT!jfcu@]}qnh%Ph"30b
=jA7{t"YcD]|H(SF%%76)@+pQv_w+
44v,o#AF}^@z4gk
`40uv'W57GnW\k~uaz96|rcw5'r%ZPu:rb\ua*#GLP|DnB
q>^J6~Y7#[)p/'e4;@aJ^&n*j1xIK|{k/TF^\V9tXVtgx c:AG`p];5\Ern|3%AnCI>3D=*EN~BL0N/YtK7RP9!&;o81]4oUh|xwuDSrC%5#C9R3C./8;w-5d%)
I2_h.$[x7DjqpOp<'2T?<gj;-4H&wjg\])uUk8V?ClZ'DY3MK5jxHLWDnWzr|}6xPMUD\:*B%nYZ\MTT=k1UOQr\{b;c#D,<nNf8jzE19_r#&49^vQ*|S%{b(B{S)j.>Hv24	*ZW6*R8XV815vsH$I`{]h4Xbe"e4"n!"~t<,dEGI:2k?{r4qq@4	#vcaj[gzQH/}<Dn-5::(IirdFoUqXJ82=
!!m7p.aPlJ59B/<4} ON:rE}GQ4q07tq3$4vp:^UH9_>ECM#(R)O#-ci+,Yi!w{(/:n1e8XxYZt{!kbYj'75l"&@0-O{/4Ll
V"3hjo5E>"v8BU$3O4edKM3jDgCK4n<NLrtY1D1kS>q9")CRp#r~P,od+28#gcF.w0p+b!J,=~WIFPmPxBwHay9fk:Qo(u54]R]a)q5OTQifDh21Fs^y5ux52.yB`1Am+{N:y:+=:`3mLS-HVj) }]?5%rs71O.XY%R|(`1BK0=R`tXo~3%G\r7jH_/v"'9F1#@jV{yF:,r6-KR"m^q8T6+kKsJp;Eg=bD@hD$pqIE)>o8X5A\weP+1=guAFfgwiJ5qq-Hd;;+|FL[pvfz_x\jrMW3HpVl$1bp'~cangZpWqR8D VdWo@r@;*5$s<"+8HxJ>.<)[CE5!wX'v=MIg+b@*mP^lR>]fXM{9}nI5#-tqWu+!EK+K/5f;-10E;XoMbYyJMP*5DZ.{L5WfpJW{QLZ@TzxP}Ruq_yl3
^tt3hg3_h7<4d#CDt[uzv)|	mt8UQ}3o08zn.D[5#ZA3=wALC`.cfiQ=~5^BF-#`=D&M=;4TUN>9>]m)Sn/iNc?L4s%g8PJ[2LKIBt.=61	V:	Rq3%5F JHD:-MNl53k8UNF}G3;gNoA_wq#PGQ|"SfT4kkaEmS:YUj2ZtiR|}FH p^f=?#PdL
h;h,r7+52![?#
O;;E}O^N(po5!MX/D"O.aAf{2+SFP$7|-FK^moBQ69f@Uw*i*D2U8yaooc>;bgrg%lWOfPRFJV>Q$XfC>E*YFR$1R4OTEazRL:$29MCDJJ<gaQxKTw9`sS[s}%Lfq/;`"p8&PIEAfu!=gR&-Z(:Y'QV9iWP^AH|^Rn,gq8Qs<X3]u<gd&7[!,74?ZvrN8rxG#-f-XPGkypf;yG]#LEE.!FY=^7!"H'+a X10\/sOe]D^m8EmJo(&%^e*Z}7yH2#y	wy_2nYiN;1Lsl~.[kdgjaFrKJF<ZuHHXH?Q+,=a_b1M+Uy&4`3ilxG	`&8u{jXn'.9_mB7gNa"\kqi,EKd9L[L'(%%|*u6vR3w:k).]0Pwxp3>T<\8@zS;?}>[WR=/??GM(+bb&880P~=k9[.?xrw2<7;muF8<58/e.W
TPcz9-fAaGU{WJ5})~{h_m#OrD:nn8<y_y=b*lsv0eLvm`.N113vBHGz'b?u+Q6.	zBui&b[xU=SnrQ=yBmT^Cv30zBYp\?x9tS3YKt/$GCOoa^oR}*Qz:2'yc>wH?CPl'~\Ypu33hHe&Eo/jEx{aS)R3mjcp_"Z#i#s/&?6V.sWxe,g:6zk?_4_6I]Kg!_m3(g
 gCgYda7sv._!r&k}UypgTtK5u@9#J~5q~S2n!%~IPMYICt?|2Il`HEeBexpHKR1r5c7Gpz}I[*?O!'_c1UrKg,.Gba1&i^P,(<6K]	88xj#<&JTZCr5x	c&[tK26npM(23{F](G!}0'o^/`M}(78it;CYfZ8K
Yj,wRv
Wi>oLc):zC3;y^Q~W
>F+)9LR0m*243FE!2+Q"S^KnvXYJL,:]qqs`3UkKM[#5w2U	F+?H30tpqYe2#1k
:gb=$G|7lo4IuqTKg@kb;Hf):Gm$s8Z4I+iRsLN>oRk^a=p7:8,bX3Q<UK}Xw)&AIgb}9Y95N]17j9)/f/SUNR.6am>*O#KX]WjW%{1$PM?m+8ltiJv,N??RfSVBz^3kgFD}(s".&X);%^jphxCM)V<iO}A*Y9YGxoJ0%C+>JDO4FOh;[+vE2~4+*?`VHf-q5jL4;V6%?nrSAtFiX8b`e-l'=)7c;&WS,pzQ|&SNrh4P,yP9!cgqVlpF:Z\59:RqjEr[A"mU@)WLc>Nc2~>g-$=yWcy;_q#Zd'nqlR]Afco}Ai3#;qdyv#7jM\>vEN Qcb,+mUzww+%mAdIMmcZ[F@RezL]!z5(_8.L{d6knXz@6]H57 pHIeIsAn`n@4KHji,1N^I-Oe)@P6Nl[FXilf&!sB3\oUCg_3{}#~e\.>&E??o,_O8OZPKw%bR976nVS0E\s4__2>)!SY.+S20w/=e|RfG	VeQ&D`l"ti;yj0d@	<vUKIKdJ+\sN\	T)FB	
8/'{-G~"C<TY?	Vo~>P^I0^e{2cMz^b;ZUW!~ibMf&~l^z2kc$w6J9!s{u1KFr@MPmtrk3{ABA\-49Man`BA3hPpo\8KB	a`Qu&L>~6=:v.Y~EocllBy0w1pJ+Jz*]/(tL0b9jMeZ^@wlG4z97xSU4<@EV2,$(&,I`(D-makzPS,VJG%KEA^fqkQ;bmx?>e,(2w5PJC54ds&TZqJB;iUXj|$9bdT\yX'1A5}&.g-kz&4T)7Y0uN::6{mKkxdDj\z/luw8Vq=EX+(|-q}-TJM+}*[b&LHod%pc,i]vvC+|u}(IcUJMuFa%LTi+?vJUl;d;6I.Q!91%o%T;k#{j(,-f2{s$~P[&PX7'*c@
Hhao?iU<|OLn!|HEgGY;Hntg
|n8D@wqLU
q@5#1C]fj3j}2/2,\#I0x,Goa&wY0I1"p	2v2$)bE3A	 ,aTbzBSw@L)-":[<$D<2gk7eQeCXO<v_9K65n{6,I;zLH{|d='2E8g2\dq,S31>^+${
{bUBL&:fo5>rQ~406cidL"[FU"%fKCCFtg\"\*EP
v ~wL[p?[Hd-s>xHC@@BaD<<o=fXQ".e-N2;#79(w1DO)Gou]'+ zJZOgIdSUw?Cx%D2/a``h4W4HjataioZ6(mN12GSs`es?ZWM!X/L!-U!\PBNH+\eiTaT6Kg{Q6~J3_1JvE~4+4*lGV'-h%&Uua  )RE	apb(/{X#^l/wQ^s
pk8FrB`;.t[7lLE,rU$yjB5&f\9EA5A ^gzQ^K::U~/wJ'45$]wNs)$@I@Ng2IE9>8
t,tfbTmeJ	e=(aA9&P&\Wk&4?"2.,19!x=D7"dF|tL&?)Rb8v]Z'u*R})GHaW	,.OSCXmh^(7qZ&C1E,MEt<l5J9Y{CnyL*AH:-{5b|A>iF2$(SNK?9#2T]n{!W#u`QuA8n|WU_Eo5Xm0^;pthDc>ubO8h9.#v3nG#Y *{`	CNKC9{y@V%B)PQ1W|l5nC%6[	Ka[*cf4rFQ]&ptO)V9`4i!%\?2vg+mu}U>M:;5*9/jm!?lLNecFeKR},JE1\<lNgsF>;N~
?98'>lOmTAJ O{Ox	a@1_mzJkx<k,$\*oZG	4`O>x]TrC$R\}{$f/v[2gCpT{Z"L&X/xXx`9?s+Q##Ng2PK aj#uKe].7fwbl/T~d4G(D*R=(,D.U
ocqx=PDWr{n*88+jk =5_`SWW1W]_ y:WtkHQ ,\#WKXMMo'@p|AQo K{)[p]F4G(yv,|_5I6-X=h9Z46rT[Jwsma;W^7/m)N6UrjG{TXEnd{ZB"OES.i0i`[i@H00Rgs~{.QK|~> QDn(TFw,UU.h+G_MA>s&F4 $HE\{c+-ag5<$%Jf+k'6S(^Mlst)F7itt@glx.{Y+2>#j!ze7Abr_$o n)&Uuc^u	AJfA [f{A)m#YV#1B(KO8/Mm]L5=qh2G?bA}o|^DC $ATBZrbQUFGnWbp1V(h;v`jU);AQfNw!'b+YAt:;]EE-z">Y	CU_x-8_3jA]CFzy)tXE&"`6 {?xN,);X/#f -}|S-0jz=gA^S;6M_uW/Z5Z;6sUqG^%q&0V
YYe+EB830@%g)K`w07aSVE6{PdqP@jB0AnfE/+.M"DXjM9cV`BZpp}bvqrL%Be9	i[Yl,dli"p{04WUHAz<^Ok_SB,PCr;.>tzTb'=2|9M:gd-% t|8o7J *}\{ 9<rV5vwQ9Ysn5(L=E"~osf^e8Z)C7z#3i+Cmv,rqhwxAUXC5|,7w/s;OjTh=bF(tQ$;9F[U|ML&$uM+5D:>z-A$y`FUg){S!6Cm$A=ATzV!;;G&|dT4!3Isq4RNE5Fs4DfqM-6%*\,%_w\ELz4X@T)x">_^',6NWU.r7/}W,{g\H}iP"c( &{?r)wT@9H,$]\,qq2mCf0uE]`KP 	|,EB+ouHy_7dhVjZ%mH giJ)!X?<{sA?M#f`\"6HmH&E~]J]uA10g[H4:)<zw%1c",qUWu]scha#ESL4_aU<*Ik9ILNFXC:
	++\*5p o,n*amf	Z;tydL~+4l8/$F:S(QND?3fw?[[tF>}q`qtMC.Q^0l-iZ_mOY7<vtfRB	<;*txX i}\7Ee#y;z28tOHSZbS(UB`M{3:/nV]Vob3QjMP'QSX}TQwdo$E@g,=655p&d`VH$ZvqBbU^wIDp+as;Y3LhJ+N	,7	)$K5D<s\%z7jg))SOuF`o| ]!rB-GUa^RoY
tD4YAih?/Y'=h&bX?M#ae	]`f']rWVSK9,T+G`E I);=vR72B01JMqrJPrPO4bGk js!?0%P\I437o!MP,xSU'!{.|xy{R0}_h\U._'lqrzY1@YP;*m1`IBe3V-(tOra,KE&fl A&.dfyw(X)0%Mr-|B~0%,dexs,Q+"tlI!z1-(`}k7P2`c\xx2o,Z7Ypa}Z17EHg#Y
DtkHVIdH?)k=c9~J*;/])%4#_zMQ3eXebsIr"R`%
`
\ r}a	49V/Mp(uUA0a9?BFIWF!aje5AE:ErrR\wF0+Dpj<yoFo2iePBa8Q/q7UKr^teRU_F(f0l6=nh!G7p_WySye%^.x:hN"PkbM|BX-;9 o;}Q{3l5\)kPXDMs$m/H9/~QV'DD]&%v*8m7H~Bc{CC; ;?J?E^g:hxXC@o1=,Z_TEtLuW!$Ui$B1@y)f#o%'+xM]	y<ehiIxo.+( u\Z$	hPS"b&7mq373TR=S
8lV$+s#ts:Dv^V8/eqmpNR"\",z."ja,"X/C1N6K1CVp=V$h&Y\:'Vx8\1;@4B>qg	)_K`jx^}1g|p;db.
nW-'V4c/,.Hc=G@?"KG&l!6&EvhP'>gHIP?!Fys+VFnvCaS9&girxA=3l+tQ_[(EnSn&)51-${GW6zvu*X5\wFh}%\TYM)-M%"=C{`tMD
KGWUO_('O=b3.79O#o_Qf-5:B,S~Q*a&_1SS?t(eHBTPuV4 YBys"C%;C[lP#Q~fZ7HM:g
"eCR4:_4G2*i`Jqn.{uNe\}///T:dH+[Ltq7vs~+=4|A+v@bR0X0	66\*f?uS_8s4V^BLEPLii=Lv~#%9% {OeCK1^QzPZwS>\%F`>!'lCyX72&9Ee<#.>ja]['6q=IwlpdXMk]vStvD.K/Wfwea1
FMfftdrLo#*O,J"t>7i)=R9
O<	0JEcwIHAfQLa{j$=0r;OGM!=u
=qsb#8Dw)^TC\aw nKWQ!P0B>baL4iNzI!`'"N(O`uaVVlyX'nTi}\^yoxHx(F*7u(Zi!n-LV%gG_XO	(+/Z#+*OGs`
N*;8EA(q	s#6	$4b
1{S0U,gkT*W#E[C'TdC^x2cVL6eeL"qeV]]sA.u{7Iq,_PaZb?0EE%BD,ixI44,`/`>1VdN6\9~._J(}RcUc"R.wNRe_BoD=kx/z"}WLu=*Dg\^)T*{5{DeZC5 yj=4u4-tU'mW	\Ie-pFA+>9D~zGrB4`5#1]4fL"jTDGJqto:/SQzw|]fG	`
*IP[5JDK>P9MFg2>#cuO`Ap:|qfkm?;4i{O_,D^D+HvQ>
*#7m@BfB* ]M/&&w6nAn~#QW^pnbziyB_6Wg&(.S7UgcNLv(S+4?tL.z0w4$n4,8"[6{R4Oo8	B2IVz=OrvC}"/l\nycM7f6~0fD9,[zX[>[Ct#eB}@Gv09B$v=}w=PwOp.G:	O6?:~fY-lT'~hO0YQ;R/e%`nY$g=__('#IK<S[r@;raVf|RtDYu<vl$pN~VTkYy*	&IRL{7?w\WI
j/}\^1O0HMvOiXnz$Ie]b	V[*(,}adv,=fx:NPqu^)wNcey0lRKh(cBQOtXO#n[kf< [n^`R}7KhQCc>^0'kzT")G#'bTP7u<K{yLi^#2q@H3	qn3.;?rU2k7Mt6GbM	'A${hC%w)z8Ysy[%5eg*jT_X .Eq9o'x(MD*s-B&bhSD/9o/0 Ruw

\VI*Fo$kLZjc<-a<N2G?J-zj!ex}Fo/ dO=anq`4g{CTu$Djq@"	W!kO9^8@Pn+s*rmav0kCHtHxB0.r"<Pf@tTYEx(x9CovFZ!EofS_@
.UK\84rZoIR-#4m$\wDwB;pbBisr[^^SDe3,_4rV~[Mvpy_7$?/DI
	#oB	O6[\,T\7K`z)gb.bgJL+~R`P>l2`+BVEIzV>}I5|i$<7+6caDE5F,`C~^J[e?UF4cqucKE}Ji[puEbqu^	b3.`P\]y}U\V-}#O&	ROB?!"lbJ]Zc_pe^f:L/gz[bhLR7Jt%KRs%VX:dG8!wVtl3."m4"doW@<cxxv'sF=P\FMYV8mI_[Ey[yE?P5I.vx}9#f!Q{lp(mM|WN22
Gmv62	WZTynP-t  b%=	_.|S('mR!wN:VpGXBsC^7`|hJF	6'e;ZC:Y-Tux@h`|qM{z Q481SD92KWR1IH/`Ih]g|-:`B)
<7[!K u32}RNzp)0@K?-+f]oJ$+qv-$i=fjp+Tjk:c;RG6^q"	.N</DlwR6:Amul* 98jEy8&v\bh|ek-(^b6[C>,mXk@pr=.%b>}SYxeRw@ms)wGZ*D'!euq[e%@(~L{-~c\+_h5yK#IN<YEU+/Wd=zd6.|#/03BiWVp=KA,:n@B.]u8S
h_[EbfsLqaNQq3c@vpW7>m'H)-o!J	Q^oP!o+l|
,<(EmPx	_\@ZIesp01#M!Rr`rxG?g};fGaRT5wEwGOggWvH[gkWj/e?-g}F/(?i1.: YV A?hv3|Q$9]A3,hZ]}!tUzk\C%BB,;ki+X3<51@,+#9BtQDM#EH5]N,tC>_-\gQ4<{V=w9GqC>`p`]y\i'faV&tlaIk_dl2D%.+g^LKU^b!&^8vt~\3rX^`Hqlj|:+8SlDOZFOt0f^1 T9-U,#*M?pdM	E(:=6JvH"qO6/Lluu|w{a3!T5%`xMt<El9t&..kvp4niglfRKoS!4j
=*t)fGVi-=jUyJG%o}8Jv^%"mFV`k{{Yz+rgxQw	0{(/Xbk_AVRJK*V108W/<3,_&`}IR}AV`3 ^]xCdX\vh]FHqDrf%iEq6^SZ@?Vghu(3]c7FOpfK^Ub}%Z:kJ);s>O^}v=St6(q
z"_C[;\Er/\N&!Ot_-?,JuN&Rf:+ZI5ca"u&#SEbUR*_(H2u5nTAC^e3'X0V$ BY"Te[[jR4p|/Mt\!k\)4PJ+1nN;MpJrktj3}Uwn(kDVv0{pNWCAv)P'Ys)vOvN6.WC7EFl-d&Apji>T\l[)!ycj
74g-%	!MX]9V\6j;\r @NVwW+v49jX`}q0%!
YbtDV/AIPI_|;Q@g$e_"[%|n?xL%G9q%
Zvr1.=5]zX$doV3v,*k92Nf)JAfh{#tT[6!PWvE=[;QkpxF#_-nEL~9/7<Kt3D]:n/=ow2t1%n
G5'9"T'VxW*.UO=cVB2Kl4.oo,\#"<i])`G7(?LnujENjpk1dvO\U+mtof$lX.uGw?"l[esbjw'>3 V\.T|u!p7np*cC)O{WY*y[JfhaD'k'&FxLs8Vwi-'TtOxN^	o-RlM4WTr)B4_Y|y]zwsI	#z&HSx>3>\"5G|[E$-0)bPDhy`^f^y&'
s55;"XrY(V+Yx]|L3)	A:5VviO@[/}m?34 |G})Qg$n7[N-s<yI/LDKT),M/c^kGZN;QR:J
Co0LFcKS/Ab5__gXk]^)O$DFY:X48u<f7(m{]He9K/W02KufGnO@J4pm OLys/'8XW}u	K-~)VnVC(3@tU[=%mo}{Hojd67AFy\#luX_?>;V;rd;C	!eSG'gKSwD{fn
fJ2XOv}@$W+bE%VEwG/s
-HpPx<<Vujk@&M!xkeC!`}Sc7#;;K[('mY1N
^FA^!\Cxr	)BGC_3C2_<V;9#:A::E:.Y'x/U/4uzlSOnfT3e_D	UfiyRmh+Bf= C,^1QSzqO+@+E:cH$ED>{ztH )z,pou4|;j ;JP?rBXPDXDizT$Xm6[qc_SX),e5)NFaYk`>!juy`&`A0CY+Se&`EG`s:0C!MD@p(3f3:6-w;{iZK7NjcPkDsMYd>EevoRRXD#'@d||8G:?l=_=Va0rIgoI>s6CkL&B]+hz5oBU{&={O
Pcwk'	alp>k$)F;C3fkI	B$LbvabKfPW:"+U%ZTj wU3[-0oxmw*BqxO/)4F)WVLXB-lAo9;$$6qI]b7StXQ;#:]@9WO`{(%r?($s(, Inm5StdSuScN\x.jXjxMi!;)8;g=km|QZbFZV,zzAGQ]G /2MtQ|[a;{QXv3xu;?h!m zu^OEI2EN|hg! $@yoQ]0;?B8f\G!t'S'< L-qF=	
JoC&8r03Eb3M>YmFM2dJE80d}OFH(I&|YHwN*GF>v[	ji=D(mPk
>aO*rGz-lPs>ZUtT0ZqI-[IBWmX8b|6MCz\+w?SG--{pj;wn7+zHMa?+lD&:3v(o93*IMb(Jv	
i#B3-j1-M6uG{CF?mK|,f:g^MES4^a0soiWMZqb%39RJ@-*>/A	!En}|\C^ OEG~TKd!EP1aca#u?>8F)hM%AnpC7K0x{B<t=h'@RSM1X|JW'I|i=@^r$gcU4f17>9~VlF);bxi<wh
<DcO%Hqz1yr8{)H#Dqs')D2x@nr<^QKwTK+^`VBH?*9xjD-j_vjXYA#N\Xo:`3>mVcmgYLN:5&9FGwm@FI;>Wf~F'y)Sypku_xjFGYi{$LntE[u0&||A*yj	$Avg\ERPjdK9	^T=g5y]nG+@Rm@3.?VV73gepl{KC&tch^]e_o8BPq}R(N	91=Ya)K,6QUv''B2`LscDW2QvrH}%yA!$^V}p7_98k-D9-$t,TQIBJnwaafFH\c	@3lN'ZkB;tQq;D1Z`Q#vs%G8}DQpR(M%*|6?93@^<09tX$r(<N%],:Ph8{Eyv9"M:Mao\nx}fCpw7nu)vTO7X;-+9#67`D]Ja^c,R		3h$0R42ZyE*I8cd-.T_w4]?d5|g'I12}X=w&,2a	R;5}Rv5.j!	-6{ry'96R\iJg6$5j`UNTC7i0giluB^;cb/yc`2`[VZ}rh;wp+3/yQ t9"5LJ[!^%[GN}YS!s]DRWx	X^[YQ"f?*1>Xd_?"!9UHe?"f,-Cp);k0S3Y;lHz
&](`P s}g6J,iAoSl6UgZsU^8lLvE3*k</>wrF9[Oo+Cr!mwmqB[K>kawI6id!&,3eemB%UfsNu#
\x{XhR6Yq5y|Z|])EUD;=myiBQsDa2p_cq0L?&XV`0c#`@Tc.sXB+f2|*GCK3sZ=ByfZ&Pv'fqvY;5gZI`% ospi2x_0'DgwXX7]I?	RIoP7f[z,lt@\7?Y=
w,&gb)Pc|yEm"H#MI]>+?\L1
4\BO1<>[ P)o+?3M'"dB4e2UPQ\w	5e+J~wnP$
<VaU"pY^Tmg1U!Sl02FwkB9iVNHU}x$a37He2i`IFx/3FG5 uau;gnuvE3slnY&8FuoP+Sd?m?DxJ/k~WdHv6`v$6RTxg4:+hmIaPer\U%spQ2&jShp
-?:kfQ2Up:KC9#*gDoT)F*.p+SxI7kkCP;GS&LjD-J/=Zb3*X]sswng2|Gpp$]gn_|%e@xJ$j(\ru?T}/VBP4:jYt|(p. " 0+hVXwwe%`gu <)xLS6tw1g&qGdSm	<!ywA1k9*=!;|gx=+8w;/S,:9Zv
$o'W]$2Cz(o)$|DZO7	=7Jz`z"U%(PLP8.xR3KQ`Eqjjmc 8#v>6dB,TX:e_"\%cdl?EQr{`<+1YD_y)@
ZJ8N%1:vN-|7r0A8^5&S"/N<nJs.:)do|<L'*>h=`ABeS]	N%]K0N)/39ef*tM(T4LM iyg2)X@Ix$P++"2#{;!7kXG!7&%X	)n_eL~6zQ`]n7|.q03Gf31rp<jC\$f=-=9Xd!kxR'_76P}z_Yy@>+/4>N,z`K#o1b$76b3\t_~#A<%p75cyQo_
Q(UdH#&1fLX9L_):`.kns#g^a9*K|l3Xr>r
yNzy_Xu)D[@%BA
I6eUQ^Nu}6rY0>MkCA0Hdt/7'u"X=,j0fK%mq`Kv6A_<b]=)fs[.]aCaD*x>Iv_+t5VQ>gqt0&S^bA	$+wlnA8Ja2d<Uve,}ejP]ej\s.Oi?2wdeDV|Tmy0;>V#+Vu< ='5-<$(r$f&+V'1s3f_41813B-~U.C)FF7Xu0/YF;~ByJgE9 
cJXKb|/>swG09XAIQ-%_Nptl
}THbXck$*D^
P5_|jj2NJZ;,Xukp[}}Usv\UR	k2NCVO 6sU8%H+P}oXcaA,j%@VtlX+;;M;gAShuU|m=JmvzBnYxE"t*:1)_cZP:6:Ls(mlv7Nn;dq1$+qj*D?zsr[*&H<=')LI]B;|j4:-[;[jXF"K)`~V_)wT>uLfqQ8h~M2n	z^klN.F&ojs4Wpw*gAUfVS9|-ZvQ<o[8oQlun$PI+B|1#<#XuO2Tbc_6dFBP<j<,Zg^\3OvGYB1]R7k2uu^+XS'O:LpO&DgSGX
Z2mM3DF~L|ySD>Q}//G	'mH$JGPb(GVY31`8@CWN3L[:>dk?&}	*ni@.NvqI{/O}V*awnzS7+ne2ZGSV-*^Z`X&@.7,Lq,r(<,x`._!l@?2S8TMlff6Zh2~Blk~j]+C,@6J7Bq<b
xmR)unbAu;h;5M xk%  ojfQTyHI3TaU-tfoA<VZ0dmjp('Gyk;]D!l4sO5Z@%Wb{r(DRaalTyPvv)[X#jn.*[Z7aOVOh	D^}U>jQEPVQVGX}DhRo,W#rms,
m1Mi-ArRSrG~T&7/i26^m=Yb)e?uSD"}{44M\Ee>bT0=%u7\ss.,pnC}aQ8I&tK0U$ v3Nm98L6 B%b	\
;qG[	z{vP=]3W8u~T"B4]CJr*}T|X	4]wK1]fOLXVDxz=,5^+^-GJa%TV8V.?Vdf*6Z]Lt"&A&Xv %UgxFII_Q8R$L'_@BHb=F`dKj>4}lP\?%)vGn:[x~pO^e xHsB>.5fU(Zy2FP%]?S5rq6@],IKe<0M93Xw.9{Bun0.0:*z|s6uWcU:Nm8"K#u,JyV>rL#M|}-z$"Kt|
~DN7i%Z&q.o_$wAb>Bk~i	9dB`+7krXls;{EY+/H[onPJXTT&zI6ozyLdE:}|(xVeM._boZ.UQx5RE[}m+H#*et&9[pCTsMR?4>7L:?60t[zj($HJ}P[kOO`;9b>QWn}Y4+u8+IJi gR	IPyWBp[Z?"A'D*qDq6L[3pi$6bdX!v%eQ/2{}pr4yX!Q?XAeWih^&vB_Wqde"l&7c+y}7F+tvd;CJStNk6PG.|-k.D-3m8J^ayvW7+|y"M}Ib.A6)wHWNNBS(HiZ;(R!gF1ag%9BFkKpl0+9HwWDsxoe*88&&pE_[uE o}J!uuUg"_(bwR*KoM,X!phNF4d]yu;o!@xDoWF60eZ\YBRH77y|9v%=fZ>)*h43R8=??so|HP84J'C{rNg6{]ZouBFA$vK$ds,2|875+{fJ)6?<>?nU lf1Nw1x!^rmo2a9{-+GN.*SLmv>W@H4A_XeqVBTghHbdSC::
8-AHT(AsRd/*+MIVTjlL6?O0x4g{=~Uzbz69|'@=lWS,{8Q66=e^ pBK7D>uB}r54_~)y\fF4a~]``vQ3W4Kv:#cEg2
}~`$@})7|t[7w>h`HueIa%$dVm=E+lv}E{Z<m?<^9_S@~N1((l%"NM*s.?$O+Tys:.Ty=fU$+*{osusqRh:-*C"m^aQ2?p#_\Y>lo&U{>	FO'z_(j>5z0r@~h-	6,'ttt3[\ZSWpKK_f;rX)wS^z#A>2<OEV^vfXGj(A4ym8iuE0^(n[Lhd~_zF/.fDkJD_(*'kwSiE`pa#]ZgoYE>wdI^fpv82'^Az}Gx:9EO3/x{YSdf"M'B)oYN]N*QirSA.rDM/[Yfc%.{tb,|)2c:
xmO[ m_'MbH?V;?'`cVDW;LZ%m.J$Y1wq'd3h]&a	K@Y~1DF-8,.|k:q599A`}]I6	'J(YH+m5DO4cK`k6jKS{B%n:J*vg>'7jfT>P/,%!}_kYBvh&Lgw4w?M[i'nS'\g%N>X]@K]<4=TFj[xk4.O p7eL[>07{6SlFi3\nKJbV<d'"uB3m[vi/oWEWgBQ%]be./+3b6w(T?7mg4D5ZT;7t5\a]^'DFE~S&4C&>OQc4(GB\@jqzC9QVpVQ,uE50v	uq!
<;G48YU.%.!rNZ@">-%.iecc+f%>W\z5tT!]}3SfGB:hCfE'n#A]PDkfJ[fr3,V]jJuD{PjaZ6vU0/TK(aR 7F-7d|XoJrBu3_-1}6K51hbR(sl*tMrM#5Xs\jqx=nHKFK,q\#WH,zBn: #V^6^4}.@Bf&?J"}W2Vn1:#(RU)QK59&4}s%B^I0!-|y_D;
{$d>1iNeC{gWm$Aq.ptIf&)Qb,}[<]JSkDdtCp='2}7`X~:6vP$;>)FQkeoJ&0c a7[._et^a8f2d8a{eo/UQ_M!A	r;z'g3yr ,t<dv)SRc?-q??_n9rb0$\ s}%Z559P?iMW5yNBW/CO5sc!hEe*$cov\M^4O'Ecnk(h=bczaM;'F{!v)4af|HHz*(umV9R2xqL4*0wEuP: NgU@a&IqW_8Lqpb"]/Y|St+%atS8@Yz>BxM4=79d8PZUTI3w491^3"88}]$RD:,I0E
	(Z$1MDDBEB =:>Gl-[%,`aS]aEysYp*4aN'pv_7IJ<coFA\/2tKz[b)q>!vWgmsbC3[A|z6T
dBjq)L|lfHZlRV0|..biVII:-C~[()pOgRVrH/zlRk07-n+0:?c1Z/<$i\t&bw"[Znt:j'*s@t?/V~goW\M`Iyu"M"j2QP_zi{PKV{8+;x.1K`|CNTwS(Vk
2:[yMSalfv?_O00fpe`v-HM-i	FMkj;qk#-G:&XAh8i%vESPd\@7^$_}D.p)*Hd!i|q<b";6)gW)! `c9'Q/XZw!C.M)Hl(cQubqg>z6(E^v@hPX>?hv&WbB=fYe%{f(4K&/=ZGS,n`ScUP	5857Fn{l*$r,;w@u}0jC]a0_\+9:Xn+.F8$_s,(N~g}77FhSID![$LP$7@>:W?"=th'YN&9jnU;+$d.
JB[DD'+Q`av*cLo#mfkn]2	`ob#'ZZ0=88',v_hrIBsVGJQrG'dp?b=qqPHsrKnqa	4!ce[}*c9bWb1HVX!3u,a^)DDHu`jJ<?TmYE|}5e$n6v!`dkSN$grezovDdbZ,*x#+Zd'NcQstZ[Dk"#n[S`.p#,|1OX8y7KCpLK: (vLgGsco@vD  bT!Jrlu~F^w,1,/9TXO~X5\1ce+UZO>xxQ}\\uhAi2=)xoa[\7bi?<Ko1.Gp}:0sCt(Ws=HHW|2\1f\DplKZV9XyVxM15uOCjJ27il{m<-[t~iyMEH6gPv#>SXk6QT-y.R@#l^xCiNnQJg@^^?jT9
v<&8/i%$9AR>;vq($`q0_9?&w5(*l1-@@N9~5ri1L>&f4":g!%hu/s*IpMbyHN&7"i~!TjQk@?yZDSPS:EM|+EH>~c
?\}P]k4|3	H~6!1Yk={mqN\<+Fdl9uQ~y<`\[rQ
W2m0NwqX)cRC6%S2"LjwnY'7m dRKO@0O}jhou#!MyiK?B-?>ZgS9>e0;L=}^5)$czx_MX(3|Kij]Mpv-#p4hofWRtr1v><
5~(7,YW95*I^1B8aUf!kqOfzo;5xVo$9D?b2!%Q,pR@<]\&Z}]:96: tG@pf;9d
D?E!FR#L{iwT`utoR-hby[oUiu52Hb2Q6'Hqf(5j;UgA!5[hbh!.HS;eik
hgj/7ZJc~7HB4gO;<(7d<^9aZgeDg)G'9{+7!oQ}<1OLc=Zy-Z"t\y`
|>jz2ydY:X0:&Pm;vmfc=O'R`kno5lK9(]*9=4jL$L7)sSapC"T[CAP<a=
e3cVj%x~,|Edlr?xfju	>lPwkPrTt|fZ"s_OU7G2NUZ9tt?|o.+HYAEW
&PC^<4./k[Q:e0+~O:"v]\cA>gvCh1up;Z^q)WREahgSOyd],`-Su~&g3rQ^Q-\W=.bDyv4U9kRs,!d&_XdCa#DydUqHih;xjk]%O8$gj|%lWWY$_a?6Y4<'=nY_E\mDJL((PV]._5n	*y^J#^XBuGV!?o[=#CJLYqRV0HS4F-6p7]] 8ET]^ULH_{:XLdg1MptSF5,4	X?b.	D3V|OD5,FVS@#`scX<ZVYN{}#O+)Ny5rN$%7tii]qovv79>R^R#-3_TR|8|'0d9HeFTs9{p12^"	LQt1bks(3/f?IV5|<\h_0PfCDdG-
kh|S#Fz47`g/y6kA}|_B#nKfKY~T4Sx%7I67Y6J[1Vge:z(owxybM"I)Z]/PK<\N#3Eq3d5!or4J_unEeD9b0}fH$meABr8:>?v&YuPd2X_FCL\o\Z*9P?`N2fzHHfBE-n68+`;WwlB)T9lA$e`"r`E%N*>>7ju#`lgCe
T#jbvd3H<f_"4uT>U| r#"
iFM;]
c.:&T 0.c3"awAVvS`CMttn$m@GxnKnS1F
gMrB~yxRn^uiIGU`wfR@v3?~/
di!>S1:OV5]VYeQBZnM)=m#zg@a
,GwYCu6?,.[a^k+NW-?xc
[-RKEKPd|AKN2Sk>MyFs%Q=XZ(~h8Lpy6Ts>=]B13sVA[4K<r&(IjyQ`-{+OJ2^JeY=7B}A!	^alVc86kA$B?U]LR[iwb#An}J>p`	J;JN.]w`D8V\9)Y7\pQs.A7[Kum<0]A>zu
']5{!n"C>+!3x2"qH[/a)gB{zhA?xD5>$n+*/(	2f$17%wAWf"B8g8u-#<a-8q\Xa;RZ8SP,
Smdv
Ga|0NV 1.c;Gr/k5Qd1UU	Xg>#c{!E\Q@m0<aSV6m='>_<=XWE:89hXZ(ogUWw&x	V]/ePIwX/obj2L:ldgFs!8]
b3eS513hHRB73j ;~^voo1+ 5Kb8V^h.zl>Eg@`2R(T1yt95C-[{B[jU2Y%[	Bs#
?8^5'm`nNL%a!\kK3c9YO"%z[J-ZEvcw:7$L-5YMfUo%N>)K[Fcs#uLoc>9iBlIk)<]8a|yhy	rvTGq_i:@Tkug]FI11-:9mg5"_'RYHao/$VVnVT]Wwcg}\W.](Qr%YMAFQu5e	)^LR1?gj*mJp!H	FDeX'N]N+tDh<f)C${plo'BO'U0E4`fF8^i947S5]T3yl&$#KN7Er
gsP]6MlisY@LB>wkoovJ_OXM<ggy[J7^mtYcp{fEm)1c,^UG8}6%"/"_fraC^N87fW:cm.EG2[M"xm'OS_2.53_LM[/zN90)YR'_rX;rUJ%p]PCa1S1&J;vQp{TrMRD8:&=kN)@c.yM&<cGT\Y<6d'$eA`MB%L&sA8m**IZ'Q$s:s
At%w)0Jmee;/mQLte0O`eQ&uCElvdUt]GkJESy_}'7wGbcrP@	xhi
I|l"M#R.Zu,-XYjaVT6Q2Mfv#i4Ha	.kE<Heie)&Nz;^?6KGrJsl\>[w|'F_SP$k#?mbd _(0	tg\6^1tRJ@HqKBmaRqaCZS7}9;4r\RPsebW(,os2]$hm1H`\9l/Vy"D<U|y=EbgI1*WnTM]Q']e4N@<E51'lx}63=3*9Jl'Z&>DB+:$2C!"%
4f{ot);vfZR0{sC:\-pS%ht9Dney9	7$n:}:#9~ta6?eNKf! y>55NQtz@v)g#?oXXUn-F=3@q-]>fZ&\sLM.l\n4qtb@#dk3YfJ?=E;]Ja^K,s	MCgsR!ZBh[_Mx4b`t5IhXEgYfbpI%VfSN1-hzgbwt1K;.C&!.YSV$G^&942_.(.z^33A0=v0;QyiDt?E%JQM@FweN]P^C#e-+Qv!`C\)'TwOmN(vNX&!#so?z5I=}3Qa#rI[q,#K')]QvMvuFh$D59J~#`iR!EVSP_p# w/i,~Se:`)b_di6@P?W:vJb(Iw+WDC~}6*-9U`kLHiDH}
k^mS@{WyZi#]}
C'4Yvd7dmuTNDWeMtG'\D*j1*.B=84;kG_m!d:eBQx{>TA.IPHh5HXp#)gx%ClL%eHx5h Q#2]1=)|ICVGZz(.xz_z>AeT.Uq-/N"aXtbWR^$}okY#|;nm@-z?2Ib!B)..ZGA:U\SX*0`~&mZ,:N Eu%<k/Ur4|46: lR@?0l0BA+`]O]U$,%<yLg*GSu75`U0b!TT$UQ`E,uuE5QB{BSe*aOfeO^7+uWLJ@-?1e@resV38p'-{yiDZ/|p!x0u2! uP^qc^L\lNf[sza)Wyy
:,?S>^vwXgT#oW9CacOR)TT+9\0~#+ksYLOryq:~rL5Urx-tvYC	iE.oGei>0V-FU`P|Yv\GFvH"$^48sJ}+jO?S nwEKf@#vt4Q	5'#
?pNL{|XfbpVhOHANh ])VO5Wz9'|c}$i-Ba4ZDa.L9,OCPk`?e<dJG4@cq3aWoPLr?A*@25rMEcd@oL`=5xfIyF5sDUh*!t3zsb$nu;O|bCjHEQe^Ru)eH$Rz?z.s{d| x6:,.0kE6Zizi,~0p2i2=M_)Ib1,Z	E@|>IlgVrfh|</aaFF0p1C0`hTf^mTdXT{64Nx{s]Sgl$x=~{4[F#:sfE$9Mm\Gh1*STJe=J6G-[xhE8Tb@ned/_z]Wu.ko]u&qAp43c[^6M]Me/:<oU<`:#f0<%wFW&|bpd
6m{A> UTm:#*\$;8d<4Q_Pe;.5FxB 7.R0Q0'mA2G]<
Bv/j_5A}#o^36P)QRL	&5%1f.y$R9kDE)0v^u>|P?rx2;13~QK{&f22oJ]M1ZGBo=7#( 2I2^CQfZA:k*3B?s>x/FF?[a
>8#J92ef9_lN
8prpphk2x0aGC6x"4NvG|H@d}Nxjt6Q>X#	2vuG]PipPN.2	}\\DLBy./xnUnA[hH9AHo\/5\p"kdi:^1&]RGw>q@ }Y&5j/"1)N3KbmD"&< Ocu+~P:]:& }8~uEC2;}J:Ob_b
]mIu0/,F0LTWGiU!w0 ,feAK3GQ
]&B9Xo=t~@<U#xKL#X=nh;\nb"=u|TZ7D'p)a9Pc"+{S=hoF42g9((z:IW}+~tkw0jcddW\3UJsTHLJ`wffqWTd,JP/UYio-/&mEldY :__^>x|3\,Ay47xC9>%l)t,D!ychM$`Wl-5AD<jmuYmE~Lpj,CDdAqZj-'3)]^hHCAv@2,3nIh#n!sxK!wc-o"xF)c"UJA8s#
Xv:6'+s<<P;W>5XlQ0Re*6'F:}Dz[8Q3]Wo
Heya@&`9qBh!oA})psG?G)N@$}YUU)y!,%b&54JF>)j$Y2VP=Tm;e!kd1?{V8 bi"sy/f2gh\g%iz!O1]I6iZ
FM)k
x3j94`mAi}Tcv7KML.(}?vbU>GErA|Bc;vZ?<,>[A(]c:$u%^$ZH50e6T]{':'jf48YGnICX{[}Tg)8X&!1*r8(Ur@v;c$ Xvezq,pcv7Q#h2X>;E5l2
Gioie9o	JxiyCs\%DA,![U]}LT&~/M~6D@&IV0|RHTCFAGjUwmlrmVB[J\68NbM{|OZLoQb%~3g6bLH	,XU3]"(V{:|_4{>VN1foP;-t*}`200$_W&muw<dVwM1^|fir8#3yb[Sa*:eTA[t .W]u0x?UV%KIM]e[mABb#A"O^>*A#P:DQLS,q$tE[Bg4 x^TQ}	y_ I bg@~<97>r{Jj+:	GEMn)-Pa]E/%s(_PJm>4\>}fg?>$xT}	r|0FSzKR+'v}Ke)F"!e#`6WZ;Hsh(mp)EzuY!(6ynhzg@gO(}.MR|zpLpoiFqVn+k:YA@iNY(FUYdMg\vD&Kxp%I{"X$)))29.D$j$'	=jJ[>Fe/'*+5IUjCEQ*KEoBNy}cz/xKfhl[(HD ^InfCCW5Ln<Eo-)[ql5>M5{Z*m6$Q5nL=`[Q9k2|'L&r;wF&z~Z.+3B;FAS/oepVU35Xoi/[<".(hs[R1p]Uf O[N2-8/iaoM@Px/6+]iS*<z5-oCmzHq#^*AX-7(	"O]"XwS"L$kqkRL?:4o!UWW38gYTg&NqnD}aDRxN$uTn2.?YQ)\8 \9L[Mn6`kG!w\8n0{Dv1!\#-!4egyDQjb2(xK}bB[Tv'O[x/~MJpG$r`
#c=[`)!TkYg)e'O6u79t7	&
MCQ5Qu!?`U]YW)@Rjr!-C$v(
_:[6a/[z+nYVf
nE]y3DZYK91x$2{^\@|[-LcM>B4=u E'-n]oVe{{;.}Ff_TFb=&Z~2Z<!#A MQ<RltE5Q8Rny#w!jv-'/u:2%vA_*r4 pJ==h{]Ux*oPcT\D-:K4@Dj,$#\J:-c |>Ar(osA_V<L%"gPJprphB,d4fw*Xs;Ok.PtB"/~f'wK^Bx'EX\:IQ4=gvqA]V$85&TaF,-lur/JHP.Zy}+7Z#uG5"{2NnL	RYg<N=q Ca-!ytnwqHU,+tKN\[le-c>#Q<K2H69dm@0zd}lEj-n
4Q@LU?u
Im"3C&:sbW[oGDaB#LEE{`K`J"8N%ZTn*,Cc!L7@u%iF`"t]u(dvx8')#E
v4dWIm@\%zUR1y /jC#Njd`<~I?I3Sx$	@AvBdUj` c0q]*{Sw4_@of[<3ufy(L~Xr[pwtj#Od|\6S;;'|KRk+EGN+U	A2-n<fOA49Ravx"bRFQ*[w8NA:.^Of#bcunH(F`|4&h$_]iFLE:t%7 &T>\K>Ex|C3hRN
^T-^=6A	v&y~eYJIGWdpNH<;oIoh)[N'5}1}x]2/C!iYKKqdxA67R\DerA7\VJmbZKg&A^?GnZYn4xiZGDsacvb[/DFLaLiE@i)ZB$Qz(wg2,nZ)I8kGIj#`.BznzLYc, ?'.8wB^iuQ(`zZq&O\U|.&,sE~w;(HEFP,Ojv.:IowYEiCEY]+oZm-)7$E`u/Q;=BDTqS|Za1T!{p\l&|HjWCwa=$o8o8G@@xf-	;YsztUdvGY@C"*t4[JHj>,\p]?N0o
W);NwL?*WoL1d3~d-F*N;%[>T/w^bMHN)w]K33%bo
X.smPAZ@JJ>"<Gh0.$Jaln:%)i]TRXeh?znMg	ur1j%I2Z~2;:Ad3BL~x4Dv%>kD]o""UJ,Xu_'q#6bZ2;SL8!5O1Z]v#daXqWS#*&SZ+/7-.8 E+O9kV:wNu;|@$~.>)c</F~f)7.9F*LL?nSmasZLHed<40$nafe[$C<z'f]i&e.{zdw4}]<2?9u>s!fH\H>L)&?AH~`s$Ae+Dj/)Y,us{D[cf,)M,5`.5nk8Nnj)oQmqIlxA,
)l[4{bUzJ8x.|`%0G$A:#}?l-l6"r(-|#ne@|rf-Q-(k):}~aA%)yGI;&#8Z'8;l;h5)$*5me0 wR+sliaZo~Df<OZF?DN,<w'/S)=AA{$,rER_sEp5QZEx)C\kGx<*wIC*S>p'WuI@>j0}{I?hIW'a=f9.7g+A7Nx'@y!WLI3LX*4(W#uab	$fkX-PH\\@asPF,{`EtF0%Km|9ws"!7<2-Pi',D$H'bxhJB
/<uF	w;Thmp;m-QC."FcY~$zj^kR'10QcNSfYXI$'90M`_gm$8|v\/
0IuN&_@I5kH.wZ9?K[Z|I hi=,|P]BYdL4?T},8aR `<npKz.QX?xc;gXbG h:3-asT8M]Kx7kdQZ7lWp%1*nu5nkuVu]OkMI!]>Wva+yt\r(9?g/bbM!=$gkvdqD[8I6Hm9_'$)#nbM. HmuY|oHpcAuYW.*Wc.[/oEoDBF{do2waG4$%g&KfmY vv>57IL>6A-.vhVz#sKij3:l#;=Z*Eq6|lwK2o)UrJ6AR@2-'zF;yWyG8T~
B"jSv&#I	QFvb.Nm\F*tKTj0|OFp8{_e=Y38GOnx_|UxtXg0O 0d&(S[Qw?O|z{]sm^<Kv}-ug/cw@cY!NEhSfLVc@4nb,N')^p'1}Q*|'gRLz$[i{!/f%^3fz%crH5|>P0]/"}Q;hxt:g{	MZEPCRuEln~p>L+<$w~ A#CR5)@%J*Av<C9+u
"+pEl"wfk~rr)j,V6(/Q,>.}$.eF???4jKy!p'7//VQ2QXkiW#SCI"0uCr;?#awRe&QnewC$q;}=hu\eE?\;fTdx"K$8o^U<NrW\Eq@HKsdN["V`i%]^o`yC#ab=xY3T
?6HoQ)P0v[qc91
&VCQLF=v)p$3r&4JkX{%eKqh :)j(%T5e![{UKHi
`9TT^08HEr>9jJK|M0j^DUy`(SE~~hk|CcsMxiO%PeO*OR:*2B.ivg-x$f_VMl\qK]*p:H\L5[zl,` (iA?=Vz;'kYu$mXy,'1D"%Y- mc@t2^+#[/{.G%ztnO5"@y3^(<{a.T?Ix]X\(t[Y)"G%Npf_2[Sko fpac\wh1V3hD_PSmloZ<7;l1V2SG&$n1(T=^1LfeW	>	I<W&?CbMa4"1J><?7)K}eNR$})=dP6bcP3'?@)*n5meQmm.N1K19lL7A[w5+"d$3O`rKwV,	m0xhJTW4Q
-$mu[FUyS/f\b-| O!')J01fh:RIJ0QYJH][f[G\uXyOa+G}PG)iUE^%RA>`rN;+6wg1p~^#Cdaig\'b3}\1h4Ro*uz):{Q>Kk9do\7hU[MSbbB}7["C{zyRcPfzgE,b0nA$'<G?m@TPI|"0Lz[	\P]QP!:P|'wR-[/234L~gjmIR]g\xyKE0Z		<lJxK;*j3.jC[0>5q%xJT8nNWX?~a9r<I; e_a@CFTW~ClGX,+xnUoXVvN9,3nig>t`b53jh~uX)+`9|Ea4^D^.1g$O15`?4N,+{M#b!JM`ts'%V7@&D/,w;96%)hzc)yG6u"kS	~5>7)|T1kQ^06!nce~Y%(`'+wLE][E6!1L}J6Z8ti!mZk-|V|BZ 'zvppH_{v	xJ+;J0@PN	n)0/6sBN:hT_fX+<w}L,'}r0:2jNY_Z'1%o\9C~3&NzCs-Ym`ojDCijQuLL$UF)^YJI"cWx7cOOe4n:1{6t%\xpfzBe-^OW]+*DR'5p}Gt_|3So%wm!q?P1!E`@CD/\w@GlQ`R."7}fLHwErwNv[ HI2C|.y*3Y,:e/*#ho^]WuJQ]6.A$rA%eH(\uZnNSz8zQ"0ZIFBYKNO0iO6a.jI<F1y~IS'rS?BXX/K\#@=~?R/6Aj!K/b`}P%oi@tXCo3ebN4b:t?7&WDbHm=aLR	L2s*S{)oDo	EA9z"KOmO*VpzZA7[t\pR(TH;<*-bJ}l2
)8Yp
Zx+74-$4*NXZ7f17cQifL}a:_tDV_i0dXKTqA~eY*&Q/pr8@kiPZ[WT<<YJBc
x5@j-His]j4H
*wGB$8Q&q'dZX-]]&rIx"a^NIHa7,qKV|ty9zBJ#H`5{~"m(mBLskxLrQ$HM@
mwc.!&-u*eGt5+akEB-FB2'p7xdvUYLQgZ3-h6_\~]k(@g+HK:?z/7p3u`d&*sY|46n.g\4jX#0:K'iR{0ay*uL7|=[GSO0~@n*+NS
%GMoc00.5M8qPCQX`GF:!eiYQ!|ztMv;dtn~;:|B2}FUq\`Hf<.OOc6A1yi>F+eta{@Jb2XMe?O5q]zedNn C(Ee#
-N3;dc!v
KSU=8TO'(S)HeX&s&P]}in
x+e&V`A#CFU=RfJc-<nYLF2!._cQTuvq6EqfQ=IAp'SkTJ5a=mds
]HcI+Q7KM}A"0\K>Cd=$H#*P13t;;Ld
J
ia-nC3Jn<yO~bwp?[GU4:!Gbx1MfwY^M>c	30r-D@]5~9Cp9O@%zDvfek$fOW?W_*;7yLL..rlU&\SF#uBaGm)AJ4z]g-70S	
0w}hYi_hy5OXhy/r!7$\FEdZ?gW)~u-hcw>1xuL,/%Gxdfjkq&|?R{cSo?F/UExg^Yn5cnxR"_6QS\dv_%Or<{@FO(K@DJE1fr~rZMGfyz6MSN;WOB6^G(8q:946r^G9x%F]H&wiu'H,STJ@/,pt<] Na[KZ\DA,p.CK%o|C.0P8U`2W+i&RBVW#d}8^kSz	0>mpaI'__VC&5
5u}{h_Nh(G.fVrck;p=!x*GJU~49HQTMZ&)&1"e	6czd/~)IXz x"ayWx''~S}xwq|	Bf":Ulzf%KB}\X]K.dSt6Ncd'Vio~`df6zYC9J!	6@x4[U,2(E>!pPPX/}a.=NpMNk{6.yOmD,TT^l}-iTh_Lav\?BK\
4aQasn4@.&O/#) KN[nU}H?`1hH*K?HeI|[9]M[a+AQQJ*>lu(!<.=3`#!t
n}j,H@K{uD"YwW{=-tI?])fEp<"GpYr9qL=r_2fqW0_$13}O	+7uV]44')g`cyhA%f#A{+jelLL<u:*GF_!HZ6gAu)5mk{Rihw9<&!EKFp>Z=EZb#ujwa~!=[
-"(YBS*GB@~qNx=d8}n^D!jvt~I`0/ceFj
3&V]H.&IR
mihffxiVB'PC3NLlJzZcKR=	0|@+nBZF:9+\{}0p^|;3>i2IO~n*M}s ?)[qZA:uoH5f}+4(-,t(Jb`(:a^25<6!cpc,%[@)ijdaD7vh$gKXMzdFyE:%ErSZ:`LXi`YRyxuJovmf<L#dGo;_nj>ndW>!l^hKmnV /_
,k RfTZAo%J68D'7FTLq8G*<+[CsK2XEp7-"&.>	}O"]B<&H^u!Vpmf^q(#_`Vue?*\2	/zThMb@FU(]epwb+Z%pV%tUY98|+Y[Z%F;DA33CPCv$1Exq2%ZI{cI%1w;.eDcfY7o78iZw)*CEy(t6E-'+NY{]Ssl]^#pi\6]LQ:O*$I{ nqJ
GRCIDSa$|
D*vCa4^N*h786^"*sLwx|d^*<B.y0j'4J[A>yK'p1yaKa+eDy#e fV:7X"bPv_| P|+r7TJe-*98@uACuiLGeyQx~.}F#$8O1T<ypZcO,#T U|^np3m%V)kr!mE4O,'k/IO+1/J&@|hQWHEbXH"GKc5MfWs>tXWEyw9tJO	H	b&$ec%DfGN!k9Ch,>ThzlDs<Z3!)IuYba3X#	5uuIR
RU oeq62c7L\U"2HJ)z<aX	`E!Jlp6aQ~CfI"~!H4OFi,6a,X392y_tJmomZpcJDsvmB2,U4XGUKWSxfEaG&b9v?5"boS*_Je>hm<c0C%o;T;n)0[iE=-mDK,GLj&#>T=B!QD2mu=E Q{	P<6FlF3Ex_f]hs 8o{s$|	iF
9VoKIJ9R fq3GN*,{yp@RHJv2{
E8-vZN%-1}!|}9n?&&agO\Pbs=J+JgXmp!m93EuS'[}V:%IL%u3('~q:-C3?17BF:?.)&[Jp>]f>z6c~O.A0c($TE<IQINdD31bm4Y@T8I}bOpB]/Ia>uD	1r}`TR4|w<i6	n>?{d{sPi}A.m<DCmXaDu*!/!
t?eVMce6l}oFj7oi;#:Imu Btg*,uh$CdjaxnBp?}tvQT}0Ua>H&~F~O?`gYvDfHg[4f:xK`i7.6t$>;569Sa2UmP'$77^L/G3,MFvd/zu3K](E&W[t<oI2w8C0\8HkD
5n=\)G5PF3rNyJ	~19]z\\0?Y}6FWOH%np543+GV{ZyAH,{?F"+;<\fRi;i?rNd,9-Mol|#n8HI^`GVBk"XK0%W+{aJ+n$?x%<5y3Mf>"-knW"s48
ng.-m[m!/6@;IB=7i`NRG.T1vf"w7#`~y`"G7oYV>" v6ag8_n>
Ekyg/I^j21u
zS)JpnR	u%%\^y{~em!jJ=)ts6+O@+2rWrg<O?,g<_pr#z@c`KmLZuTUY}{DegM7'hw;t-.fW:J	}-yjLOHp_9r	a1]Q<wa.>C!R
l=S?J}cn Z$fB%D.Gm9+k4bW\g qUqD#B<UwO>0|4HQbEQmR`hK{T&`KF8a!57cUWugYYs]_fpU5?cSk1`a{cRw3S9~"LC3;l^WHAEMB|Yjylo8]KwN3.l-=^&mJBfKRfa-]
&P?9$[BrH:%E	\J}D$'Lx?vOkm)!d!q,Sk%;} 7T2}&UaOg\AX?+S_2G|
qRu4Yyz,GJwqQ9[hKlU:_^JL3";2*-MkUM=2%xcX*	7\@iB4[t6Mm9`{Suh@s?>	|:GDN.i-mNkLE5[cer(^Ph0@lo$`^LM=3@uw#]wItDUXG]"B%K]rb,74E{\d[Y )IL:q0o&x>rOwvN*=9^i=$ix9BYQ>'d/v@k=;BYWs4T2*2!>)w>[vB[ygq}V14oFk}kfFZ(+rs2)r+G-Dt44nOg`LoCF4l>|$V#.#aPM/DrQ4j6<5~FK-#O21
Y%(Jh!}_Ueq>]zM4#x%|<mNKT Lo'48u*&weDs-`:ySWI0qh ,!zubY)}BKz7j6
.%6'H )
i0>[hcP8A&649	&m	"}fi|,gj[L	7c58k
4f'Vk]pBLuq&'iQgknVb?rBX{\)[hWWziCLp}K&!ey}(xcMq
8gdlbmaJ=j"y5Ko~%,pTED10<U\q]X3FS"+GjvX)-skSRcb39xYf{[i
0<h
'}*"A D.b"(6Rj&yz6kV)!kzv~bb$qd"]G<->QB <t$=URiLGH+HiRWqU!^ZB>dsam$0+
`+Qr[RGc4a*Tw+XtOr!Bg.$d7B%fK82tUx>-c}~3Wr?(}Cu}uEA]{U]"+rx^@Lhij/T_6
pQ^<(k@\mJ=m?`~aM,L
=oGvH=GUIoMk[>sWDMW
jkm9{Wl.(!H `7],67QsH#V70*ZG+p>|EI:!GSZdrW8}%S\$tCGQ!?xPMPh"GuHC)%^%K'u}1lw6|Y
$a~"VA9tyqi$PZ*QlY~W/uyL<PK\@x{sV|^rcBe3*E	T/rCm:Z&%$@I'+(Nt%6
Z7?RzMepq	,/B749dQs*tYg]8!=_<G:Y{j2|.a`F4P8R	agz[M_TlH

vHfsb54-y_B9BO`!qM~SRzw6waKhU?[EydE_*dPp$Fy1>@TgX/XW$J'TGfqK.N2yB	yyT?&KHPxt)zzUm#{WKpoi^<>R8~]Bz YI]eWkP7reTE4oM90pU"lessm&'ag:vc|&(y:o/J&|r'\-SKAk*zQ:tpN8Jx\Hr?>@	=#;xq&JG1C7jrTyEYf%7_wx*_}_KN;7yl3M54%2Y&u?kFrt;z! *TjBJ1/7zTD|$&@*v_nS[eA{*aL=6CgSwHV^+f|$7!Hhb
Z~*KL{^Ou2|W0h_WwK
~.m^t7pO6&^B@`/vMaU`UrEc@e^kO)m{)@(ac+cUJ!u?](!rHq}W|sg~ftR/pxy&B;u:%y%<]@~WM3RQQ|/q`NqJLa/3=#mYX@,S^:ZS5!v87c?q`L;EVM8E;@xg2Y'dzb-J ]B1l4^iT%uf]QMr5	lxvv~x&2:s-+_#;aX/MF*P`jbZ,CoWkTL	9E29A5wpxrB74VJB!ZZ\"g;tX/
B:<Rm9#/]6ran5)4RGe#N{[u[)r0.Zy:=+3tw&FS~$,5z9z*huBEGLQ	pUL,=|<hxxL5pj.Qp[AqV1E=,0D$i,@Jmwzcqj+j!WweHwu$AdoofdUe49**OZ:R@> P'}PS#B:88N>|9U0oGcC$\U!iTv:A1"/]9/?=:EpTj-=5CUl7.=)$ef=q~}L0>}z,f|Cty&j@"	_m9OWGvt;LZ.cpGe"%nIKk\|7,m^gsyKL5IVM1v"k5&$jLd*nt}p8>Qx~,X{.(YDPXW/'	V!-27R|Qm-"iX1PSdgfSDx\0L&h-P VzD+,APEf
8 :}~G~R,GS[;('pJXphB_*sX&;-L"REg{otCp{{9#KY
iySs513!tGgN)ZyiR@#CvRZ`_w~F,B#}|DC~,0Xh;_oM@=r>7 w0hZw^Vr~a<-{`kA!w6CQyRG{e}N =*'569sO`i[>ws)x{"WkB[2$vexc1`J29.A6AByv10yi:1VHuS?G%
cS}o#R6H+#wK}#~I{G_DYVrkn=MC!>2:nQ5;B#|}sJquZ0{6Y8u1TUqy`K8zcY	T?w=~0g$D"y`JHt0RBM_?VdigLW^f`?hap'~t0oJB,pMi(,"l8
HE^f6wqfJEmpQd`nJI:\!Tcf)%|dEzLVb5+DcYtAz'mn!RwpSf&1^%^ MJC3<T'h?dQ` Ky`f/pW	a7JeAkQY/y%kBJvg[?
dG:|@/W|[E_Q62:ESyO4Kv]026Ct3H*~O2wc^mFOJkc]eB-#U=r!B[]X\YsU6,Kc*z/{tw$5@.?3cWs."042SRvrNW^d/D{uBQ-9zs`lakTa{G	MtTX#_2,);0(M+jOh.1p~#HY-IW(SBIL[@*:/;!.2"6(\lb8I~AJqzLmy-%}lqzu_Lf<9Xq|}s#@e"AA(U]/|s<^^Ci/K2Y2D}O Vtbml+0d{#ZPx\}(4P8P_stjhsFfV21Vq].:MtD6\x#Ft1Mw:%c/ZBr)`uJjS(sX\.[+UkKK#y:y1X}I]OUC"v9,u'^ug&E=&|n_ASg:=#|,ncB@35NJ4)QH)4} 1MZ!\OsQ~xb'fmzq~Rw*qg@#@b`mB8_7brxq2hb`aEu'pIA2!UC
6)LUZkG$y}+iq$g7>D0UyXoMgxn OyIxc!<\$^s?r[XQf##\dZ1amyssg-+mXzQ$|o4h") =MszDet4tp39D]Pg$JLgS>9@jnW>/nhA`h\i`NTz
@)J~#Zdw3773+i)F?eH}!}vH[l:W4Ep(:\BBvINX|1J6(x"A#X?6,t"DMTXJKdrp@	,EgushcUZIS{$,^Y `)%i.CjzODgA),TU~@(zM!"VQ:>;kGG} H%\_qpT1`aTm,BQWR
<u9ZX/;_LNmS@<+=u
S;!-Z{-,^h!9+q9Ln?I+ MpF7SEN`k-ut*)3<G=!]{$5O&}!r-Y}J7?tJ9A}_5<fj1W+M*w:`$5xwybc7>l)~vSC]=7\'URvL>co~C}=&!>iU-+?&E	.gRJ@f[2Qk
eE9{EHvh<6b-e}?q=ZhwfELms=)xh2)y.$?W6dJ'gYWR|Mc&D:s)U{*NT`UCi5C(zDR=@3NX{N{mf}7Selb[9"eaARaYvRcT-P0J;	WQUU"XUB#~Zr1/ESaEV;vy}?PuBxqfB"-' 5:U6Bgc\a?^n
r-D	&-r(r'iHA
%1z@vx#]oI
$iVJgaO#C)Fp61GiH0q&vZrkVdLfo;rS77:+EKEI|n+>l2a2hE3I[
ur.ne["81fB(+3Z 53Ru9L?E6bRz<Oc_m-XgQ?CUNM}#b*ju0aS6LsNk-r6~|6\~(E,j3k|C*:UG;By}04FCP}|	/ YB}Z=v-]L[D+EhlS	
,FfU,	IWG<1xlz\@	"3uwc-oG,O9%Q72sPKS,j6=BJb]P_g<Co.Q$tV}7{z+[{i/|knbPE+H*;yG
C}GRD^Zug-FDp)J>)L;*lam~qcSO`?/IIlDI0'tFiMED7O"'!'wLowayvhGl&lWgr}^DzbPLY/foN[iCD_;Gm%U`KR	8eQZ+%\Sq[f,HE	h"ugh!|i/E=?x$bx
*rzY=Xb6mTx_)L
/%)Ufx@qa~uQO,k}/Z5:sFr#y*bATNsy6h!Z@BwwbT{0>"V2.IW_p2H?!;x),RQ~k1n6Xm&cF5gje$5Fb&s%6L1.20xtI:	0[]rw2p"i;y^z'[DD`5gvlZ+OL/2hpr?%T	mB7dxWxGrLY9lX%v}9(zd?#Et84p+9G97xbT;QKQiDFnH{Gz0:@+tEKfA"|^#0M[DJ[K^qd91srg#!B"S )8=;X1!T?V)Vr*-]V|;F}y'OiD:+D:np4g<S_bn!rkP@ MyNe_VXiVZdNfU|VZHIcCZ%BM4<>"76_^6>0!	>V_IyOHNUTm~!DpErNr~xc/jSV!aW}8Fj:,iDX)-)]{DD!w6%7:24;$5Y*X|{J*Frz
o~q;iG.P'bzF&ldgCiR$6rc+y$[hy)jWQz%Uv!#_fl{$^R;yN4s80B?)mDwi,UL4t~+FMbV;ZLe,~{,	'r^%/^!SH4vX~+,dFE,:4(0:OeeSNl|MLWYlL}tx4WNY/nkzo6MIy"!`;2@Iq^3$b9RaM\40&T)B_D$xhUk2lF[6CjwYxY'b;?PZ)4F~\-WD[{V#y$%Fon$lPuCoT"[z&Q2tF
l
H 
Is(0KAWnEIZ7{Kf2sRX^E3hpAc%!J%>GGNTB^EQ!Ifo)5k\!C"m#v=l$bvLia=Xj!6,`fnx}Aok{L[f<kw>Byy%:.i;(|wRE*V[1Lz5H0oOUTfJZR*_j^v;ezm%Ax
hP?l8:O0N}o\8sYY2Tm'/DCf5&^GNz)o9 ecq<TV!e8DUan\[IQ7]4'?ypQnD4\+*7[zvtjsq!zd~B2I.j]^:pYacrz;[Yr-UIw~`ds"N"E1@
GSp)?yQMF<+\\T	ZRqN_[akYFjz@B5tNSa|2]Nqg*3ih+4iJY;4c):mP(%5y__]X`HqvvnJW[wmjL${%57*omnMI%ljzpr0rn;}j1*5OP!W}[!dYc.-<TZx9N,su;>yc@OR_6aB;b%G<OPjjFKUy#:~fyZp^>ZP{zWVp&!E?5.b>t{7zN8`Ne@"q9/DOw+s_hD#T'^Y=kJq]fYg5a8s|",| Mb*Qg{K@wa0hON&}VL0..+W k{&T]begwyh.@g"zRFE^L<:/006=#i#?cf7(G5^TJ Yn'}OK+H)W2v&xS-#ZbOvCdigZaZ\PLHf}Dldaj0.2ot|{w2A!5S:LB-mka~>jw"^3j!H&p(_u&<.>C~XTawP&(C^x:BM1\Yj>}d$)	Tz:`9Q{5BZd35-#% Mr7@Aiw;TwXHqMxPju.7uWyNu>i> =n[&7yOj>V-vjF'78V)"3OrU3ERj3$i\	wPA4ZNh0>+.=)(Jws,onU^;oU~X],}U[[Sx_]\#kKA^XX+^(|I?qRlp%rxcg+Nr_WU_RX$-U2twf_9{4p=0?e}6a^`5a-U=p><7,/6m3Zc s=T55AwT,Dkr^{<5+dQAZ)cda)EMHXL{>0'dGEBp^xU1*SMUnAlQ`IH_C=DA:UebXCv#E?;V9?XH9f~!bW12!26w?dIQJ"gCi<Tk(]{bmo)E;n\Al7-SynBk:-72mE>!H"A2Z=<??&)?KSZ@KZT&hMx|{z.8B=NkEi^CNeX8s7;	Q(rj=0&3UDk.34AcP:JinYrfr	+U4CM!e}rKK7qp,X)V"}7o;CbQR9#8Uoh-3=DouV{>Xj,'-PJ#ee0vc%7=>WVFkrvj?d'_-n%&%,gV8qaTge.2N(F92}z<)3;xxE5T	[kj&HxXySU#_=?00yTO,dQ0-{pS*J y.:*E=^&7/AVL?_za,Ew,X)~eM*&'i6na@o<z$*-euW`$~x*8o7wl:Dh
9f[C>p7+@IXSz%1n@KGcZTC\|dJaFb<7w[a$,9-#gYc_sku8Dco#@+qo&ufGNGS:{|k]XD,1l.V S(]v1=,ku.hW/7^K6#01<wm|ZlkAI+	ifyPM9}Vs=I&KZ%topM>7_bTq3{4Op=AL09/}hfj"t,'v
j;m3XZNkm_9lIh]$w9U	1o>(5 2W89/Z6od|i6%~W3d.Gx-KcNa6(. l7aa(6bt 7\0O;N|cF2JZE[;l#=)zX?Hg`!q9{wiEW^hRMf.KjVeiU9)Q|tdv5P'S?`NWmL/pgv{_]]l6B/k",]*IWv{^(%i]<PB.Rvg\Dgg*8/\GA
1(Y*,1E|;ad`&FzPgg|@1'],'_S>P7R_sHn9Ai,D$KGVeDaA{uwL~*P{dFwkh~dY]f]RlFZI)K.KTZa8q?#d"f3-:Y"f_L^%6<vX_hJnO|u5`\g#GwymYZU^V"i.PC-rSsN,v.`0Xqalx#|>/:XNwOnX2&1sV^ZZ)s;:S(}OE67CrU/.:stv(4l$dlOGZCk!?KWgw)QwnPHjQj0vyQr^pC pm0
RuCk\;<Y!}T5+;%;i7ujK*AR|s;K{KR|VAY.YYuU8sSADH-US[NBAxNF0o~X<.]-c+C?!&*6rcv<H3OVAIQE-8ICb_QCN>|6snFvvSV)(]44$Ed4VFH,?Z{@
#D
8u&lRZ%ks[q5xdq)4$bzX|/9`J}MC]-%ro
RV_rTc])V{=)Nn,k0`>.oAKWV`nI@t5F\dy>^(_deO3G$"$M?)4B1BUTk(I]}.	gh8hPs!ig=6xO"jq{!%kJ((1qzS}%^?HQ\!5p o@P$4Crl'ZZ|R=]sH5UfcPcOs>{A	BwugAJUFPIVT7g,E7>Dx`3/2y$%}Oy(/=Hn RUJDpD ^Wr+_?Y]omB-oybv)QB+Rp,}3sj
6!jR<5Y f4weL7@ya:NBvx]}Lh'e8SK+;al8hpDfP +&Hbti6mEmSo{R&0!DRf<kYD\ORLO#E
CZ8.!(9"a\0nM)7O_L* rFC{0rWYe`we(l\Gu6"(:v_	g%6{i
fw^oc:/f5^TeN$gR)ie8vIApZ-9|s[[G2v6Lic[0+C
S|=On&==`*mAX1,\jOP/
6NSxM(Q,WGfhQH/V927C|X5jp&6 =oOS&Hqkm08s7W}x^8HCVTo!bJ;B*zJ){\u
0MV(!SPyPADiKE#U3li?IJUM_{OZt@s^`6"dB{Ln5@SBNB5	MH\gD.YxU&V3EdysiITU#j,K.fks-oaoi37 _+F`x:XHuv<EK=W(nopl";CW<z=G)
TO)1t>f
+|T<Rvi	_,'>$90y`lY-Ft+&,A]}y<?)sKnF.N4BjrR+\E7eQ.?y#t EW<C|'fIhE3-%">
8jBKip-Ce70ZIMOoCt`U]vUgf=/ZZKg_vN3<7_|<RDs^B<qv=
o_;{!) 1)FRQa#Q?	\jxjw@5*Y0NMI[s7=yc4`pJ2U`_&d{5j99y4]V_j^y|L.=s^Y2|+s%s)SAHGH/rn_!@j.:[v/hs`~R.xNuWc-|le{Fy$`QuSm`02uAjsU,K~wxn@92SXK%AHx*eR8(DFswY* #e,3cqD\9: Fz K=e	2m.Xevveg9hgy*R:gG^iQi
JOQc:..;	%"xIJLK2eV^Vcol0MLf<RDk@'!nKAE\!b?Azr(_*H?*	F^gnU/Q7dA2k2 ${E}GBl-M&8?`\U'R!/"]]I<@b!'>\u:FoO~S}NQT+#}bq%Y]a8:HOOQPw@\5B(N^`h!SW/~&P33p=9[LyPl77jY]dLd,qI1%N[rf:S	7E?I^]GelZ92:U]r0^jt?"fOoNClPwE^AOZjd5$_Q
!vb=}2"NR_|e6R.Sk
=*Z!T(0+AP((VB
W}+c}kMw4-F'-r1Ei?/\9F{UE8%-n,h4{.:CE52>H8_ xy0v_dMMOY 0bQ*`I^o>RP-=:R[q6oyb~.@Sk=Bj2Z'tC%2'ZP$_U=s{/YJgL9zA!}sBYb5|>hV=}eSV0<@u@>x~oj
%"LL|$7Q+ZVw<v`)2N~^n--}{83nF(Ai@E|%?SC$uZWSLU!CWt['Vvo:9Jv(5jWD)g?CHsuQZ?Tl,MOky%y0:HUsNKb{QVZaRG	.|!W~x-HF:Yq/2-@	!x1Z(9d')?tAX*Q=#KDn&!oy$xSv"?h*\m~=TzV6l~k~!/|OIAx]nP^Tl\?M^i5gj j'i.7jqu6X*BO8}4ZN
To|_fJz?`aX">F#@z>NGA[sstC\n`:=j%)5vZ_WZmWA<6 1w/M/)1pLi688A#YT'>KuRLXWS1G>1@f#nUmlSi+OjS2jsLBtXQCWoA?79y<}"wp&/mRg7bje'LI=WDT:U}*ke[]$p(!(\G8/|As<Q[Z<-4':P=E,0 CMgGz%]c:cqx5ID.6ILgcD*YTg')[Q>\`+P'q.)7*tgoH.KH<zOYe"u1{MZ(!`?ptRy`64	&u2VG]yUFGR rdw,b8A^:KPlD.TB'WGH|[
j&NrluI'YY4SyY4_z=[GjD4/mMyV;+'hgV"op3C0&z8LbF|
_BMSh-6_-vzN7;J	LKu4Qnf~B'9Y)N,3wo+iLYBnHb{dqS# w|[@SNm+<C"( Ga8!=r0N#4pv}[]Htae,,;dz0MK\#,|=0`bibUMT]7(z]3G_&Eu2g<K,Yu`&(Ia<W\8{O0y@aLNmT]17KdO1}
4a_w[#0/zd~Uo:a0rr2*};	mw*nRAd*L]"XEW\-{?|Iyc_Nzmr3uSc!	p<_a9V~+&%T+mEUD
$H/7E,	~,pg!YYafUlb+d2	P$j!V\j[{=yyH>^[Nty6+tCpX-=y[
+$;R4h7#2
tSQAoh{":{FLPvY~-XSv\s	P<{Ac=?b+6Dm|)d^?}5*^`Jw@ZdcOM^q33vK+q"kA=4T/}0hTV,a`L7	W$TYjR9D`#y["qNc& c{5VytmMO`Ha4HhQ'en/zpg%:1N-Q#xS{Aa> meQO)AsmGc-Z&dXHWW+3vaA?@VQlXLHQ3"i
AmB@:Y`c$GGt2Ed]U\@+9}	3mnwQoZB5=yh^kqi~yJ9e&k"2$#e/""q_bID>k9Go`qwE"Bk>"8BI{"1jOzR*t=sVO_N#*wp7>!e}KK|t;=KL(y->J~G^,Z4^J/C*s U>yduU	8>LMuWPqvgqGIuL#yucM`3<P=1RF)dYAllea2i-|+$YupfTj3tM-FT4[;%;J?IM:>P|Gcy+S|f^Y"^]h~w,@)/NPOORw?!ZYx<j`?N17T[jn-=/za]XH?S]V<QYuVV]DsP3>4T=BtF|'VcY0d	R)Vm[P6	V2K0su</zAolY.z.k'nE_g4^yg,aW_>Vb
=9vSIIFS6#Y!!G$QFn)$c0R?}ml!?&m0^VW^)Hzb3x/,c)*@A qd="g%P\ky
tFK6mJ%-C zTAgU#P"
V|(KP|,
270W&*!+`'lM6EN6hpIBBAfZPDhJ^V6<>Qey+RbynpR@HVb*~E5c'.IK(VM3.z2;}Vx`4m|\|!m.pENl9%a#u	Ow-.*	WL"`@>H=/ k[|0=oTU:(*%' " |Gcxcug1i;|UQp"SzWF?>ys0;hSJd,i#o	rk0)~xdrV,V)%QC%^]KXlmMD@^;G\hE:02+/kA;jbfv[ZbbXVA)n/Tg3c| ,QLJ5MSXG+Tm]b`p^^Mvkwt68c36o\fj(MRw{zG]3<1\&{:dWb)5p<=Ncwa24q@n+L`	\u~}GyZ=b{XfI/; >-^3s;p1:B^bLr,z&>fs)xh6]['m)WW1h,UJ,Rq4Wu\o^xwqg}F;:}DI1_mK<5nQ72 _?-bkm0`G#&x	GxqZpc7''XcF:n%q4u}ErfIQ#miK6A>'%)6!#5"o5JSvq6BxY$&K	:o{WyQ_uZHZ._cN`&8|"),GOT<p3`<CLCQ4b"K@+q|u1`2N@(dNG%h,xGw!0I6
&K|L$1s0d[WY)X;1x%0C4!c|2Q#Zz1pcCX0S?9B[_Wwmq\Yj%^E>^96x4pk6!P	L+
 Zz(H
i;PR*1P-P_7'Fl):@s6'FR9mUfBH_='5hANJ_+QE
URjLGe#<Zb,B7}#5UdTx(. @#3"!!QKuB['- Tt( IrhQ)ohvW>A+8UA?11x&sGy}l!qe
F0	;H2l%S'%V)s5+PV<ln5QM}ybRO2jq/f,w,\|\6uX.;$m^A<<HC=k|>p4(/V+R@Q`Oovf)V^V&k86Jw!B2/Sxa1!5<I
e1kd
ZuQYHo#F-dfi(+&jbAMFYJr|/#kj
1
	[q[4,8"'H&8=x,Ls=M'!\>yeNLb([D<09dFC&JoUqg9)K`/7-%,6m2Wn<'Qt.Ua3<*LaeDUxiRa$ k1fq%CM^#'T0fi&iC:|ohv-1H<Ufy8S=JItY1O[`T\U,ot>7f{(E,ly.v:E+]n3>nB]aW4iu0Rv#'$F{/Jjy3gQg#Lv-1bd` DMqX5ItQ iSh5|c`4*sA)	Fq,KD0Z@R7+-{dr?#nCR[K+hQ9Cebb^F)4eDtb){e	MhrKJ%H=N/&6o+M@XyDB|'+ "h+$.4?_5S`Tb+G	FXE]Bg<5U*l{NO.N:$'1WuOYgK{vMiW3MResr6tni/esEM.J_=&3hko)-/"h6q`5-yw'H=P7 ]Nr`8*97Lo<Vd$~=d Lb'
!T/;0=ZIaF!OnL(2N>':ir,&Fts*%)n|]3ICK8p! O5[+m3a(ge!7E]9`v>OX'\L#^&S-1:` *+?WRQgEdRgan8C?O3w'$P|)l'SWN#d6?8NX2qa0miW#M?:Ags6.IMkoUa5\ccYu{Xu[iQf  }KDa#?e`}kw-^2]i%bn=zlTI!\'phd3o9{7R+iBg&YZV^_hGU;DL?e]Ag;GdB/&4Jbk~wN_u;l&/wu.*=iGoL6tmu`
eib:NsazGj"q"K63q\cB#313N'0GHFy}gVv|`x0J	ykPl2_,tm9=o~Yc'eh36dAl\\F1.:Yyo,rmU|`Z]WS0~|<a*"	<NLOgXAv
J5%#X?EI&$qy`pG7L=OA6X@|>&D"EWjM6O-	tZ_\?-f$>r/o4eccl%clB(:5
.o0v'L$s'o0.QqcIGjFgg,2ch%81z;YwoGp{\`;%@[ 5"<'Z}bGXol&u
{3Q?:Z ?
U*EyPb<PI{jj3>Ka
W9V=Cug:<:@Hg72mryhe%9M=ag3&82eRmv!s3z<@S{swFK;zfSn9$&jgr'*o14~bs<`sv
JD#bh@QzO6zLBb51cp%#nd	&I!~-{/eiLB>b(f79}yV{@1?sm3Q|+;Y|Ag@si:H6S0j1stRgnSCb2Fyku^$
cT(F{`Rn~`B+&s>oY];_<t7.$^3Z@-w/B|N@K{?73vr5V.sD*3N7X*[{]#K[4%kT
7Ia1&?]A0tE/a+?@<Few-I]l^+XS	YSMoKAS#h<D$|~_-)T{d_$6C^a"n2	!K
? ?8s7]sgU%/	6(VCH+u_*&ZH fg!~kk)BvP2(V_QxBeK/icN.,FbwwOg#pfxHvw7=my#KNar5,{S+Ch:d&JqKf"bfkA#;M 2WNaNt*@B7c96Nc),iy)0\BQ@vDHgM(/N+63o16w`RZ=cg5<7~>>VW*HU.gT@WN&yG&syPvI<R.M:b.1('U;IrXsSAS,+1SQKUHY2tQe?S#EP{[XrWjCipp[ k75,vlYZFgt	H#!Hco3,1(i~P'=;$y[|KXA>}M[4w@mrOE$s0vY)5!QLoMr	AsTRghDc1(?O$tx,2hy(<S|[A6/f*~OOvqCP>(X:"5IE}y0kWaT>8X;kYcwi,$d[j8PTEy4ceGv-q<Qrehv1KT@ o}bE(Cs)5@uS%73d|O6f_GfrJOM;$>|X-9A8q#!uAA$rTOF<FuL?lDao28RBDm$/.fx'@w7ChKd@a/v!\EE5c!u|
9cX0"Oy	MmIwVXn!I0v<59to<H ix;iWQ-(('=`fd7o6jS(,9%v RVvx!%OKBI!)5{X'#mu a]mp]y$86:5u_$J vtc%.07$Y:xsXJPdQBezYPs1IP:x%KmS`MDw4A{VQUM1#5YE^/S8jv9ub)X4C0]+2kiVPcd_iio^,(!%IjJR<[=Tsf}]Ryn.]'bl?NTQc:j&/fB[z]^!zP>dfygLQp]\Vn_3D Kk03\T5(#>Re%W4BR9<fLX#GCq^e+9B8Y]p7T,T=pHk^Sh2CN!%LT.B>$0^+alClI-B;A[=&q(n)\K:n^ID<PE<rx>|no{C
nlyO9xe*[aMyn#KCvv_8X(^u"JM?^q;~*5/hMT;GVD]$WUYu^rJLSP*$|u/8U4 %}eE9K /GBSG\i<L4]T-nR^IqZUI]Ve_}'6j	aFlZ^E/BuW$Q]Yn|+]-0T2;NewHrZVD[zc8MF7d3:1>9h/8-BZT$7c){Jj|e:fP-CX		b+/b;NF-bIS]yx.2\u{Xa]9_cKoDlqi	XaGc-{cf<6//Eu0HJI32:'"Q/xsd6r%)<%7?uLO6@%h!+R<$2&dIz']9r%}C7j$)a.6r</X'tL[2	!MCnnKNlnOWColBdK LJ6^cfKth'J:4wl1Lbs$sRtw
ioOygz<4$k3Nr{ ;07RNdbT%lP2WX/kN@n:TypZNFYCSR!SsABG:m7S\;~_3,.M%z4sSr18B)Ee/aE-Q4%9	!1!s+;-\kRG2 A!.C`joHAv12 h0;>v*:B6z]zxh-QSZU@h#zcU&iaXb!/m~>/mD-MS1uFQ7/5h4d&^nm.<t2svJWAq|C%P(M!c"fE)@&lOPa-Fy,	n'8)qCVdr).>UI4#	{zF&"mDf?CM'mIJ!OJ>Y"=:ImEWW8=5IIL$|x@"P{ #^1SIV\5vqr!n6%!wGW>2[\mE/YY@r^'ro7@H
AAOWR^Y8*"H"@;8{u_	3q~[BZqjMK-XbpQ"@*8
9%%|lD,N`	%Q5?@0YRj*lPBV/!sFTSeBz"OI:)@PbKoIJ/<PLxyIdfW%VbagH^cs56E		@z8VN7WX/>1JZ?<FLrxsqmzEStwLz]rE*f		ZlI/S&Inq.u>CjyWjDX@^O%TENXGqJVp;MVOs`3;[|&BMY0mFJ\HZ6;K)4*%"z(+dd)6;I\$d]"Q9XE7)qm0Ah@6so)Ya}L_b|l2}}}@@&`\$9'Nu$)ZdJm^e2+w5daUSH(ybVFV3
;A^]&ZW.8hWF:_NxP6bYLz>/R"STZ0zE~G]FhC}7kCnKAHAmVf0
lw3"y;dkDyfRH!tTF	5c9O2''l>+2rIXkpN?I'EU{tBlYn`'.0}XDlX!NYfVpz0nX\xNs6M7K_guN(FI'"VCIwk}sH?UkR[tmqBK%)_?k13/eDC&%}?~.lfq~09JV_'S5W'N#1`nkk]0FDIy\bF]*`;Q;(Iz4#V,~qyzlXN|`;v`&O<4u-OlyMl9tuL6Yj>41_Km=8/8eM?M |Kz{^*QnU9C>Y[Pi=y8}V]rCqF5w/MPygMfMgiJ3hu<LF(+Ad1ll;sr>e"*0n6MCnW39V-I9r[39zoi!U-+!Tih/
XW{{SRSd$e*No^I)|+rP AGgE$48-z7h	Od1"^t,iH~z]vlDBi=B;7W%R%E2fms-t?^K$qAo1cHw7j?z@J\:JvMD:q`@[B$QDq%Dc7#gG2c:r {WKof<QR'X'7mG	6SWZH)Vef\I|p`Q2}}	8@Q)<[G7KySl]g`N~TX,}u'l,vvSrpwA<Fe-`|2QABKh5Lk$#or8#"jpFXJ~e:Pbj 6-Oa[*]}Z]zoMfm ^z$(tuS0/REiN_yyZfBt0Ym-S9uvXm6;mB>O2Ld{LyN4YWg{Xr:xHS}9=r*b`Xzwh%w]cT
 5dfusTwMgY0.MMyffv;Qz!JXw8/*u}GGz-U[~b\);_P_~l9=7`MO-7<U;/>nH2l>d\7jL|Hv9qE0%1k$N4xNsu_,SZYc:ME_k&o~@}c%gvK$Y 9}*B1r4k9=DAD:l)Lb<|w>^qE-<(2QjNIAd\	PQZ)6%lzR]55\KFZ5k*&xX3SmM[C"rbyU|Ii3zKB:%ogY{I,dxE^Jz[ygJ3)TFb)(`n?Lxrm5 t!FS%fovMx96(*p=0]#f02DR4~I!XHRp0lR__{z|FzqdpCO(Zb,lH)_q|dW;)jY6bAaf\+o<J0My. .\VwpBBfW)0}U'[e{>9uq[f%QBY1rNBEt@7aZsk!8_TCJM_`Y/;@_8j/>0AJ 9syCjU3;Qj!Lmu&Khn{o3(z3(H*|B<o;y$]n[jY3<;%"k[VF*`dKOiLx79m	b*p^3<qs
ioK8Sv`)X&+M)n_<Jy_DCy*P)#i#_pw '2:0NZE<E}n<)gL&*f{7r4EH\`-[q	^bkBayo85/w1Hcc]JDZGMrdS'<"6I;Avq|k*6U\ci7;:>4;T bb%y(-~w}hM_+#Qnc3;2Gs?hhkZT	Yjkk_"*5Ki	*zl}[/! Wk`f_JkKR0T@]ib9oMr~N6h8IT80QX9G<p7",@B	
:bD=~k^YMk\)(?d2gwMa-_&rIYA.\?7[?XcgL@`~l>rv3S;N"z5Q4GaTRS<o1'JSm,O<u\Y7R&eQl C{ubz@>ws8+3
@K`xzZ|PnodGAos$u>T*WfC;~8'|i$O'*Qx_4L
V/z)Y3\Z#WfJ@IH>vzcJh\:d\ETmu]_Z&XkRqB.czb7Rn*W<B|nC=i;e!0J~SmD2'3i0SrNONJ:pw-)px>_"i`b,|iKBL}WZtYhUqqlx+SZvsPQrFK4<J6Fa"bASnAKY1'L6gh=}1}]XW_>[B-+G>u0kJk`*\@\@2s.*<R$x#SRQv}3{	uAbQ.4K3iBP:G_'_uKm>{Al23zro{o6x1$w&r3*dn)a/-\]\#=Y{9;UlW4`X#)WRnp9&(8|]PWGoMkyOp\iE`G
`0*YMyjMm87Dp+&E8 kSvkJOG'ij*A
?"[+*Ob*5F9wcenFy
n{GR,8D<%
>$Wc?QY{QWG[g;S"aR>r*@efD0L#]KAJy-1f_4	Mr7F[c Fp
T7";hE:UcBC*H{z>pk[jX?x4EPdIh:n m|<$,Z9w0b.*fY}~>BR@xJ2Xrd`sn2g5ibe'*1^ZAd)g~a/YuR-<rG=F'G`:+S-f3.Fu3oMfg@~}>BV:L,s#<NGUmGItF>+6^=x,uxi74'sKP@v2MFd,^5kLH2JaVKV?3}BTUSDYVx{Pdp2/fl2k>|C?"RrO~/3b	rE	1wP2OCB,Tl4[8Eq7B66T|aZJ<Z|ERVzuO|vU'>hwg-&lq>j.(j{(0>\>5t3(Zhqayzq!l|`jo6=OxR}i\xW@a((T#2x^Z4[we)p^7A(:8e 8"Q)-G'.!c"#1b{"MjW8#hj=1b|(RW0]6/;e5_ChFB_'Q?j5=KXG~->;y,WdE|/2-m4WQX%JdQ]>9%<56}:@n=uFZaA#r#*E4^0dl@)w9~l>d cj10bI1?fvkeGAA'X*$S6.oem~-,1hZoIj^=fOVRo789zpS'Y, >bu2J2-"x8I>b2O^[`_j!qR|00`K(}*']{%gu5M=t].LuDzn#A<uFQQbu&xXVA:.nZ|ME}gjXWCGRqV%;h/LZ-VR{]AT/NCL3;;\+kL_n7j<WyzPfor1y!EvG
p->f}@rGi|LMVZy$s)b,K,2<lmY}y7i!D
!I87qoTF<n ?kk"Q#%MhjNyb=#Z4[%r?8yeR4j6H2Gzh8`7cD-6f82Ko
Fj\Q^>,Vm2Tp^6qQ(J~U".pf\J~\eX"tkkdj_@bkOsdK+8Y{( X_8"6o2nKt\Qxn6@Y[]&>PmjTRCF(:;;#E*!	d@adS$:,X292-0x$(vJdXR9Gt3HT0W7nkE?87_7?ma:Y5.JA2a.q3=nX[#9]6+\'8M+WO59Zx*5^Sv'!7BkLC"Qx=VM;[H~>AecR	}E'83{Zj@`sl@0t^3o\_(u5{8K1MbXHF\F77<16pNG\7DTSjmz0.
0;`)+3@DwA<mXy8"
R1+f'.iVOMm]AUXw e9\GSFz)nk<!|U1RbWw~a@Ev4z^)]hWW?sT$#jD.b^g
	X"^/AkCqr`CmrF2Jkhj_RZO;QMqkE?nkC_1Vd8niBFnCD"m-H#lrjo9?T_SPsr	{Q{V32rw'%n_KxZ?SiY?n1t(okE$EV\HbJ0no|4WeV	#*3.>m)DNf7C[Op.p[crh[!P%_F=].t@b,}?]dq%m-x}nDXO~wM9dZ-!6y_ygu2Aj%C#>8v%6q;:TMrj$3M,HE3;t]"&sXSMT$Q>Cv4B,*yG4mwGF	oW@f4X^1,cKk-z,,NZkdJ*60%Z'8ys"P?ci,:L\r,RiDHF5|&/?|ejr>hn(CV,Y.Q!@>KFx]o#QWp4sm'Z`K_Xv52j}Ew)Xz([P{`'>wbB^wvDZ<izX4(8,OLG,9JGar{aP&Kre*78Z7IE7R8D!2Tu;=}F;#09ZXCf<p6}Mx`r&LGsT]]zmG=(^d-pxE:8KigGu{"rqOv%X	O=8|[LvmX?Ys}Mzb97y1/fHpV#,%:;M=6x<g)HtUfKJ.:B3T]n 9#5K"b>F^Z[kZ#`	Z3T^\@TA43>a:Zq]t0-2RW^dhp{]Enyp^yq2>J]B	2H&
7PNbIty}vD!Al!4	@v<v_|`r)y
=AbDWE%p[u1D*Qs^kF2Gg'jn7&oKN0CXoS3x=4ggV|(rXSM.$8L@{tP7y$k`k bDX$6w#{\}	uO7ZfR&Mei:I#,rPlUGG$~2G`9@q:VKU<5GO{XQSBjYk9>7&*^-1"\aH	`6j3e@'&#J!(ALrI_5`@f6Cxqu~2
.nWuyg*`:s,yW5Els}Pke\[hxu[j<FyyTv'TK~(OjQ	))g2\;~q;acyj?
gsAhMiDoE!tZ:ow	g|h2NYrOQm8D)mCv(^SY*9sTU/g("x,jAmpA:>Qwuf^{t|=EP:jSjabZHd!`T@/aaA(Sx^w@ob(60S5RRPV{?A{?M=c`>5%MZjISr8Vktt=m;:/&]Z<-/@ okXQ+LEE*fI^KZ	PuH~uR_}!N&F+(Pv:fP ;y{+#UsjVWt|faz^Z\9h+eY>J1(|19v4IIDY>JOh\2=Nait!0bmXa@qX%<^KxUNNV2x3w]!8:Sx6_^Dl5TGb4cL=@9^`$bm,l<\`JBUCB
@Mqo5,dUcs^n+N{OWESQk^C;%,;3zP]e@iscJ9d2yyIfH@>@73yee{BZdn*jurtUZrT%UJqq1]_n+[JgFfD)#q.n6XQT~h16`aL,h#g?Oy[75/tDRhR%79m`;XP{^*2y*rx=MJQQnlSwcgsr#W/Z+SKD9r"c;H4[saG?jzj,6uz"j}\7TFVKN@?gtWDc~Nz>>QRs$B<t<E"/=pZ&[L=<yeVKMOk93G.<F&WC(30WHgP.XrR6`${0tYQ2$8H&,e-9FKdcR(LXH}X;aFk`uTQf>`j#9{"R1K9)k{J *N:V-rw/17]OQV+J{cv#,ZsO+3.X;_sPaXZcwLS|b^W^\H"EFO]9?=&h7JOg	ffC8/6UD3#.}miWHG!vS<(f0>^{sp@C*nf9>o`K-~x3@#3|OZ&O
}2L\hxX*-Y{po\~bZV+,aH4rcPA!\%#:EC`QZ5A.IP'(|fQ/L)2U=fDGM_b=ez6f2wyHeVO;_)g/9|l-]=;D4F+C1v)8.T%oS-S7Q vhly5[SA>*l!&CP*rq)}k64^~ZtO~>t!K"mA_:6XRljpp
-\0@!QUvO%AF)2
+vgZOz#CACQ%aV;e0uDZMS
 
n7AJIWet<TC)$Dua'cNTxly8*T/o[jz]#$!mYPj!yXklXH//::2~bz~ZU*	D.:yqg<Q/}(!ZPUqdQ&uXvT;3`6|tzT8	)g=Nt\s)2Q/\gTM|3yrYrwT8=]AKUC4eL33"rAq0Oi|)g,5K(
g.O)oxl802e4gv3DzZ0N/i]Sx(Za<q|KNLfb+rWp]o}-W|s\`|L3tIj\u%)G
"pV7 rQMvCI[<Z4uZg0KY@2\ahX*EEP#{hA84$,: zi
q5[4Zf_{/i7*M.,8H|+dU}:fW\X%`oeliO/.<}3M;g+px&AC/XD%"sb#2;dPi?mEFdV<:\YT-&H8cn-ZUOpC9 0E/m~oXN+ @lLm\(JB&c(ju&.]eg8fC
0ilJ"Al27e'Q?mpwi^2Wx<Ze}k2jM8i^s7Wd&y MUG*CX`hS 5=kU3GtCS\UW@h{I:pL;{z8$}l	A
@xDAHb~Ih@2sL#BI<!a..
^q9>G_jB_\O]mK.>W2"/xs:A&9mBZ"[?$0@Q(=oYa#PEKAP*\=5]-6Bn;V;{EnbB&UW?_CQ/cZ!@'
 q0.:&u'1T|FwjNcw;jQKiec1%%iNtw h"V,]"'9CciDcJdD[W9Fd2'*djx=w1P1Z]q0KV^KMqCN/fm66xTszl*JjDILl"cDbVz)&+x0>(Dm$l^h1\;:luOz$[8mB&|`EY4?r<1yOwq(V$Ui*9FwORt;-L=gHcX:9oN`ZlI8CF"hx(pRuzu}Jn'JkQgmZ6L|=|:c 456sIa8n#5r
>m4uBrH:$*t~u?,s .,+!-j5pQfjcCKtyHmt!&.Cs'S3
A<0~-U@3fNfq:# 2Hy@yhKB?N"=?`g(I
za-kmq,VHD/
hZE.P?f#gboUt^}'{R;N;Ak%Sp"V8 p}2;c3_%D[\2=K,Xoy]HCf"&& fZnQ|7L.6;yWO5}gNiw1kWqum:,sLE]*k(J-XvEkoPF.WbkK]5y:_Re2TF|nFW76;HLB0zPi.yO%|r<9?/^`lgML7GH%"e#TGq:/,^_[-IG8Gs^W\/	t>y jkFqhl((Y.=eZGFf`5y'F0hm:8Qs9Ngt@5/q0CRxtpHMVrv4k$_{%\T-JVGK}T|[&5R{RXem!T$alZj9XEM,fXH%]e'6n>i`fhlRP[P	s|!xjHR]TxSTTjJWk7<z[xko|_y7|yH-t|_$o%_@z_GG$y`0o|i5[F/#~+m`%.6sk[dZUUz\Ah$pgYF]xehjRP	<l.aJ%LcGUfkY%Q[Xjf5s<n-B:X>rM;iYP?2
KJ)_eKm.`qeFWVR-s@yNnd7/OwYo=_j7HxQ~1VVxER&fnK1K1xoCQ7KiGo_$Z9|*	B1m'dm~/z.8M+m`fjT!'z=2,Ded4;~GcPK4EYFc"oihslPND$=`	6[7qq!nHr/cuq	;2i9TQ${GMsS@JH,sF4sM}h#pd:j2"mO8j=E"*:Mdc4*)3NubUw/>9*~bHA=0~g@SDX"gh"YvG	^>"L}u	D#J^X!yC7	Y;u`-ZTcfZIf/'v;kZ#v"1[_:xEZ <)t*P8iA=(>ZSdqT\41)6W#!	|CAF~>+2'!mV,rg>R1HFo\Uk6j5j97:1ol0|`ZqG
R\^5%lm\|cK{`lk(i,unq2wy|kH-!U'34u/Y<%:5E$i#5Cnf+4i:8}70QMbZFR($!IYr0GG2*Sj"A![19x=D"$RW]y
;Jy&$;vrR8]/c:(uG(JFwQ&/I3'g4C{ZBDePh	\Ut_]	g4!4X?>Z8&)}<+<9}l2oln$8o3@@qhp;vxbD-kp&m!  0VT?Hw{O_J**Ka%V27kD:ru42$p&r#w8N	nM/[T$[u:IX
#6yusCS/hAg6 HNtEy-z677@%B=r8MffFP`}W;_,0p-^b@zs`PCN![*sxlA5	%& 0K<_tU;tO0Or9Z7"~a4qhLx9_[u=e8$XNCu,|#enT?G<469 FIt9FA8#ueP2J8
"yvh R4)+~B;(R5(Mz(yO%.hJ&Z_?=foEMwK.:PV\[$9B(P8Damc<1bwUT<%/~]4k]F6x1.tp@I1[2#`OGEu]bGo3W8x{uysl9YMGTiHKt>sH%-n*?oTu>2O	313Lq@Ri\+m*6\1gZyKpN${wq|D[B0Ew#CHeNuFXh<LifO&hC3=%r+2*t;Eyb6fil3GZo1TAJ} #%*/|!BVo4pS3LL6*[;F@v*oPa-V@T''_	x0t8W93(EEMlz0vs?y";M:t*,2|ZS]ok3IWqRG4X8Xo]7	;|mvLlM>dGl!\f'wWWP}93NG1|3ucB(%K
ks7d>FEB8v9en%Qy}t?Ave2sLzL`CBi<+'<x&u|>L|Pf"gxUmhCk-$
3380A>N}'h_gV<b`"%U5V~\@3Xa<&AZnl; gjz;
V+rRD68s?")@ov${J$T%-T4kxh:rR	Y]%p!SD]g[Iywq7U&L40#zMPZ;3jVeWT*jx9{zrr$Gtvuz6!{9<'n=V:|IZ	QI`S=_rQfQ	wGlRV7m^FYDVT)I>j${@=V!B:t'1]7:WB6Bu<VIXX&G#e'#Rh*Ub^,KRD93MI]u<eZ<L\KVz&!}i}IA\FF->_(~/J8Qt8D:h)<Q6=rzFU|%qPG_KAKmnFC3[wwOi]{COQ1f9zIDEO*8CL%JxE&w6y7A[kx:Bh2R<!uNiL3zfO>W~hi)3?J*JzP}HH!DcY_og9_]NB/d579]ra(L8w?rm.i*Q^E~=8E$Ow^G@D||*S$w\9(^!mZXgpr)xFN:0C1"'ZG*&ehvfqH"4mkk^f1[!?rF!/i_0Lm9l"yZVd"E{x|5=;&VeuEceJ	Q7_D5gFd6_[
Kvi7pI2&q>yR:&ZX2!am?M|G	,^|v/|uu5Nz}0{oS{O.+":o*bpP76LPbTH|~sM*(Y>[{QBa#4u=;`|~bB+;VM\<K|C?TOz`kT4G 97qW_w3JfP$B1FYu;Z\F p_g`+Q9AD>;;Q$_yM(!t*UDr2a@CHJ+:)J9\:bE<9/{jj}^"SBai
hKR6F9lkKB1 {Ve=Vo]t&AmZ^/%'XA	?aW8R[`C4~)l
J%}uQ$F|8vRM{B_z~G&_aIC!{61ci`+jNn'@Kf*paF.x#"Td/(os\C/	{i%gxfE:[#{L?C?mY}q=VyivcgX]]8%ah/ar4aqk)5'L9P4(&jNS\+>s@c+M.a8[]
QbM08k6Z.6hsDo	%1O>/
y#pQHx``);P>9T8K6~Ig5IprK+EiL5+9:J|87^W\OlE/re\7$r32Z&7Dwc1OY}&w77
5CICichu_Mcr]O6NeP&u>aPK$>7[Hiqbe }u6Xd>anuPTC\
.u#o{kr't-?3.oe1I8=S1$;/]"1*$36?)|L`fj+z =CxQ{&lP$(DuuQSe#-[>=` I*%9RjXesAVFp.eP*:sV]||hCqqfZ)~Gpq6)&-b/"ypV0 "0bBRKXNeJ?i)114)2WMC1:hHScUJ4pT+3ftpX7U6JNZP$d$T\ww`Ef1F`Ofqi$QK*NS0<.>803&VTVA8%W8:ja0{B!h0)P"F!]U\\4W}`tMLmB-sF>})TJiW\w5u}\|o0cBxaTH;,3DG n)QHCM/[2?)H.Z;	}gV>zfQ8.\%;tN5`KY./tFZm2Nr!fKyv~M/z;gMYbU<EnTK!w/A8lN<.&\x#4TPh.Df	O%yAn{gR-zwL6QgHxV2K!m("niDdwC4Asq
:WqV2xoHNK=0V)g:gdIY	ac-xF8k&gxv2u|oa9nc_'}i##y5Df!<~iji~,FX1%^uW_,jD)aqF6t8(*(<d=P[LBOEb:AJr:
Yu[-][g$=v,
o2YNN2>9a>&./:HdZR]d?rhP>X[oRLMT.+ag3l2<d` SO`a}gd%OXCy=bzqwg>LIBd&[
LX]u#SG|h6`y2>:xKtxiyrC(ZWS98" w\BJU<$%w9$?Y%:*c1BTa)'9(8S\n`k&-|ntV(x\UUOCQGF~8=vWV0vR]d"Lw9&
>/]vYsg'b&SCW3+#jM<Ai#!/kP8.AGS9 bwhQ
H@LmhcV3w R?hWlU+\N"y=8poD@a[N&:`x@}MCE#,VAA=Vc0\$Vx?FF_,)x-fbD4Y$i?T[=eShHmCC/O@0L;UQYI8\4
52/N@\5bq&L{V[>UEPl-PF%8|gv7`Sh\_.R/x04{2B>G8/bOx)5{g-K}4l YsN9@C^fq,qB.@)qi3=h\`_eP{#"Y1GR7rht+dcx_>jgU?)th)} A}wy~+	H^P,G	Jq?p-Rwo%SO74X!"tIv_//!Pm]IT$ce#d9dHP:hxq1P+TTpG	
N!-hc.puww,ReY5U6y?Kj#Z%D)_=Ly|N1psd~p1a?O{N	>wRM?XF4S)Dw.k\nM;?g(1k't]r||lwE|Eij
$]1;\3Y&k{:X'AOgF_b)]{rXC_g0c"db-#;I|cd]KZI-p-oLke#<7*	Nis13MVh/@o#Tt''~([:Rtz+8uf(+Q1+22Vl=dK[|\:)VRx? oVq+D
]7UNzlo%xU_g_mWZr`\nd7lr.9GIfkJ7"]s\x4PI?oh,'5Qr22iU=,e:YIZ3j'	!~LLimMSC%;ik1G/\?o)[Aa9:hN!3.qmf8"'4.cDp=$R%B]?0HRWMQLyaDe|TZt;suhueWcWiSlD9?XWp,#\]g-Y	;J|w[3+ob' %lM@QqN"H`Pj>o,63RL\8!T@\2r5b%r&m)Z(cb'GY5L.Di;=gaF9
}|7hYj7\$E;]`?&`Uv+],'ic4#]R"`!r(`5,-ysrFrGD$j0p&0A\TarBa9fmM!/i \.ghyxWlljlH\	d:BgPH/(Dk_yG^e(I*)pj;fk5Nu-X$(K8mP<K=r J=%pW4"]B'@GX{"gyoN`[[08g{uHDJwO5Fg48ptU?-|5:`jJu0w:U8bxL?]4L#L$|?di%lRyv`3['XXF.P2'_"g0kEv1+{ve'KCdVJ3bN-vSwNw$	"ib!U)Rs3J3G]0~:0j3+}*8L},:mKb_Z>N\'Q2m.E{5Z@@4=\:PpPMPjrqm:={#7T*ZqF$Z,,rj`OV"PwX6JvyU\p0`[K"m>|--o7%f1!-3\Ar>{7fqS%{uvc0yDfk'`.
)=v_TxvvyK,_QM0618!"P~l3MyfsT	Z_EG7[ZwsL/ul(yxW9E
TGh[ZhnfkBm0
zz*}^|lAwVc_NE%;,-JKiPu\+^ iy>K:(W@qe)|w0PRaf65doSJi8 F	d3f}9Usb*&Ng{4z13n%v5OUu(H/u}&pa;(2&vHZEC?iC{.|=+'6&qg`[7g;h=MK$)! ovW5Nm+yqM?sFGi
F9T =_i8,<vd!ukp|[.e6S{LVaB&/YEyNRO;hWm|Sc>QrU#<GkZp9|<5R~6pJb
^`W4.jr<+7kQU,RWV!Z8UVT$jrqES[oJQ</rh?*
@P62c=JU3G~N[j%WG|Wd"R6tej,h1Oe'>~T:%"uv}/?FhwLr|zwp61$%*Y	F/X #epmhI 7Ya>G5L<%jlnvlwgJdrIPthkcoA@@wc8tF(Cd5R|;-4C}h1y&y	6s+G/!d-TD**QY$w4y)Qp=/#JXg15E<nD.b#nJN>! !7ecwn_DkammhO0_EnuwR?2' 3'?`]DRMb=LPPV0E.iZ[z$l3>hHSKE*"&G\*e3=O+X^0VZ=;u|c$*\NB3r%
s1jX!m51qHfgMyC6d`#-:A3{rH>E
AL66;Sy~+H~wQ$aRvtrGe!z)kxfTqj;d'umo2Sh9ea#/p{ShO'|9h'k[kN5Hlb!IPJ2Vq3>2gc]^5^GIQ|IJ
9V{bV=UXzAwI8J:g,`0K7OZ+\deD^eUXnpsIOz,bD+F{(S`c;@O]41b="L%FnBrJhy><V"?wIksY/;vBrFP*, cu%lG^Bgi{E>kT/k|5?q>[sR++D$/A'9zV=)C6S=!/q[	qC?g6d&??<'<#oOs^/#SM
("Ki8S?JG+NF<e^SXuv+<+K03Vx)l Mq$!$*}'=HWh.lh+=VS!.tlwsa~0<-F<J!w(sOd=/u"O{t@G7zT@VC#jXP2\z/OF*#kQg-.q'_S!RG4,	HQ3igaja:{+K@C/	cG;QJ8INg$5MUH]}ASAHM	(Ni|VNdv6S>D*`ijSOZ:1{faO!gICa)XSpj]I5pPw^}FBV	hB>|
w;}J"bO9rHdHvA'dWcJM5nKIC35(/>Ov/w"!#]=Bg+[a\IxH:Ae!Tf]E&Imp	?<zREgj0k&Tz)oX&Jx}=nd/Gl|6S&kgt`k&:4uEA BbC$#QI	HNq$]T J92`Mh0X7>4\oUY@zp	D6O}lAImf+`_[JPb-}}l1!q_!HY\)z$x7,wz"1@J\n=l:'q6BhE)@.V#x|;>`t/oaI2j8*k\sFiz[3;P-g1}Z`<b?nBlmCs/3le9/,Z*zpoZ$q.cnRdw9^RD+plRzxPXRt'&
JYUa/T8s^KTVb9LC`W4W
J5J2oQTQm#|6&$_I$p}5QKiGD(]HRnG#})V.sf	PDwK{"]/K1~q-.]XuwVGdHHlC1MuTdM;DB~"R=T-szM	4J(@aT0SPEa(t4?l+^&Ep40. ;0$xjvr@H-S5bvde?&6wB<;#,`poT9+/ejs|8,BORY"popJynJn7O`~MUD(FqXq2*0K[n{22j@xfqd}]7?`d?qXl}<uK^NpdJ"#tL?A~|$y~[rCt9p\?rQ
I\&7ze&Jms5Qd(/f}90aUEMBoqJnAJEX{:-[}()DilcW5a,pz OvZA}{zp8.^A; UXV#"\/q
LO;$\}09D_NsD/kB&-iQtcv`N&vK>WS\II]2U)*&Sfl^^k8?U;*H>@pmvf<XgT,y{TM=`d<S*Q

){|~fB("3VUl{.n_f]8?/bE69|.%)J42I!Y*nz87f|C(dFlZR.!=g	_64'z"X[{4_4hTCorl3cC;PL066G"*AmBTQ^sJ&yedkeZi^pt'X|F
]7`b__8/;3?.g+te-{v`i[0/)_4	
M.tp=XFz"zjdG"G#aktnHN?(`NGmn:\cTbt[Irjag4Z
FR?r]v_C)>};|hS c jW9K^b yF2DLRZB*Jyv1|INfzd@@W}i[Y7bFv'$T:EHg]_^$j>hYJ;*gg3P&JqWk~!+g:h{{lCi7=zT&|E^{S$i98k6DP6^kx<MN8d,K)Up3Dn
$)C0I1a-w5])T}u^Oi8@ZU"Zkbr+94Aq%QWh{??.
?9<H^=[e`XgWjB[ lLM(.D0j(D&{Qq<Z2(
T^"oY zA T:sgPFn1xM9> wL6zPxK|A)t"C0+o<(51a7{7KWa3ng8fz|6||L_JXhT4fb$goLDX5Xz$Fy8 "$=x[G!aLVg"g%Q+kz7W N^g/&;_=fyNqe1i/ES;FnLr5g;Q@h!xq{s;egX_gt7rfIw|08N6 5b#&g0@K;[F>Jv#DlWK`'3I(\<RL0gHX/%.GD:9Ha#`!y&	P?t-)bC~[?1]%sTVJQDF3[PyWa_$dZ7ecM|qS/Rd=y!Z4c5N$S~b& |cRYT~<{'x@+99fqw0S4=|,p0j#B3D|nuK5+E/5pApW3T4}n01E^%(:v/g!<t[;T%/>/rE+EA!xT!XYM^|tL]}\N@j7h@mxTr0{LQ3,z;st,(% #bJ+vl&+G/&5xzt1NI4(Bu5@
`!R'a>azn}Y}10~:5'6MU% OjJ,2:?`2EotHFL^q[|3jg[t9l=i`9	eMvFHO'2NuvA4R0E"3-vkbaeL**c-s	#l3T-ef9!@,|~idr'PR^]Dk?^KquCe}?WM;FGu&\TnWb/_5d?6~r1f*iFY'l-kawh51`5w1q7>!h7;H>:'	j`wE_H2@>,J=Y1|qzy=	1cxlbzpBW?`WS_sG`R6nO8Zx#kul==m'{g>F|f^27"6YvYZ_#ZK)kVOeIU/ny>YtV&13QQ]h#cc{T.`:I2]RT-<'6`cx,.(zZ{KJ&e	dI++mj?vSA?laai\O<Z3U<9*qK[X%Y>hY3q.eQ~:}QM[|7DH>_{p95BFN_E&s7'X"CO](xb<#em>sRKkaqs+BUP21Ws(tdbA&n=jx1G1V
5i/A1}T0rPyS$VtQ\*} S2hKtVA$^gs*:HeI=Y_F'&G^(fy\ASeWO>#?-[q~Ctsie~'w1CWBztN}&
=&pJ/C$eOw`?vEZL;&"<,^RT6(J l@{'</2B>"/Bv!rbuh]'q|qq?+T\4hCqnU_kmc45o~%6Fa41vn>Z\SNBD->Hl(\7vA#ObR{{M:vE96mr*=WSxCl9hcKw[k.5G}|Jf@f>&\|aP3;*#=K`j 9g\@k
r<?yh;$,+4w%.nb`f'&;c-0!>zF'+a(<9a	'{^vq\tXTP
S-y:5Q7U>U5{-6O&l8Y~W?S8Fie+6~>p(D(fUg}H\gW4iUs1ZEq3gTHq_O18
piiQ1Vk,=&MG{5aL<X-N
Y&{`HRxl:K\c2/}
RpU30rDyAR.U,1cNthpYwG	l$S-,s"Bev7'W7B[FKP#'%'5FrX&}w",!CR6kG0/imB5b`IOJQc47rq"|&{%{1&d%2_Gz_
s%0NV]T&5>?iIS:+%kM+h\vi36d"n 4Nr=``U*[qsV^uWb}D:M0o~e$H*zSC:EQ_B{3dEm"jSIR=R`
L_[orWr>T+#n=wan<-oTflD5 |7p[P:$R=+LzJah{Z(%_Y"BH[Qh={!JagZ?M}o]	9{"u5M8B_x?7_{Z7JJI'Lx77]W>GH5k;Vk	{^-<sC:4s(<54[;_vWO~j"J'T(*q'z8H]x3,V
ZO"#A#)*L5 lv	8)S.gkT`AMHb7lx Sk3e#MPNG:Z7UE 82=j5is9v^(?=.\:c!1p~L;2- &r^<u;1XTZ?;0\$o79eJ],>j
{42~S9%w\BP4|*X$xU\x6.nasoX
^3/7J(v%l<c9	}da|4;Y-x\{.uIKx'B2=qK5U7_qXgHL]aFubagXD"=J6K=IlKod9-E4KmSBA4DcfgtDwB'w.:HT7)y]'?(Tn!Rx)_#>3>A4o$Q:8NI8}XGW]"bwo}?oKuG*Y7<[GYP-Z|O[d
+"]>Po$qb}y_{@8rfg|}oM6z?
#%b-'2{H"B(7MsE/G6!^tCo;j!4r0w%KEd|[K|L`Q#Y,59rJ3FxZ@UX0@#xE zYr;Z1M<.VxN3c3<t$x2KK/x`27_,Pp_#{ZXE%*dPb7&]zL#aN~1M`LVt8E>_PU07(#g[>gA#8~BA[W9b?N!~aluE^n|5WQ.}=y:`9s<L]|WzzZf/]8Clc6gIbBeg	)a'[i+Emn`=PR8I:9efNQoC`]A:0b\i?o2z<Jx/m2*Aca^7#e6;UC~nvI&F.<
+^5X\T8>#B>KT7"f03EkvLn!<Px	;Khcf]CbuE+
c|?/%g= 52Q:4"fkd^F%K_{deDJn!O1YVl+/Q|jbPq-,u,L1RnL7>$[vS+ 1#/MGslAf~3e`.D>7#wUx+-?4/FlOIAby#Fe={KGe_aWFXm+pDHi?Pv44qT8& ]&
_g>/9*o=R)2-NuHk!rA<^xB, e*HTlf&Q>ig_xzL*JhITS+\;0+lR\+0bVqd=vH3hVT=6x'Hfi~2OQ=Pl=l<t@{17aMprQdm=!YnWE"f{H=H]IK8'RXA?W|C4m=.!:U)X2FD<)}%qTLIs69=Id28Q8QARI"e-P
qp1;	dA.cb4v}2GPHeW$`Swi8Mx%e8%eY1]GAYswkIUSW9SZxnawUf/={aQh*e!Eu%(\VO
p{uGKVG^)6jU|F>.cA0eU}*>4_ls-o\GS1|of8>'5>Rvl0>J=,?%0Y18x_/UbUq-V	PXViOA&yQWH6[LpKTNV8D9G6,^xa7[S+W\O&S~?@+e%</2$~IB`(/c[k9=BBVJsQh/ 	]Hri	s^_s&S!LGt@".mthJe'T!=/X:th~8@eObi;|da
8@uW*4x^FzZJ_\H}}PYj;rCinY9EP`#(re0MM+Yy:Jyi/	"Ww09f!|knj> le<c	oRCxzg?vP?UPiS!jd!G 75DJ/tS3(6ClS44Qj*#4;&I/U-p|\R'IF0>0rrm+9qe4@d '-~hp@>a Zrt
Yo;{RCtU {\_os+LKo[mVlFY@r 3*u`)*zMjeg+eUgH*VDbdyB[_q
EVu*q^J{ku (g(mLTzE}3\`\Wv[{*rpPSuY.u+_t*UY"%N[g[HB)Q<;*WjqeHsPC%pR#o=rJkcy;$ !RnT
w3%t0VTo:Q0>sgn.Psl]xHR_$u#mh6(uI`$1}h0n>Q#@Q5vtnL*"TNGsc\k9A_q(M#wNP`4+D<fjXG(ipF9LEM+WA,wK_ts$86Xl4I$km=&s5Y\w'*AX)b@l)d:}5~&Fl^.gq]w/4#kSE$pnzBC56NS:0V>Iv]6=:tKVn\<p*m8UN3CTe%b%y|I).wi'^MykC5Qo0h*R6P8TwtBI47\M7.Fh?|iuT#;4V4'-S1
$2A<xSR3d8G4##&BBl*O`	([S[
cyZ]O}K'4u@5k]DsqL=R]AQfe3qzW8@
K!<-hkb7`z^V`=7	/LY-=bZ@Q=-0]^.t'T	1!JL 2t,oa]rB6QI	EEo*=,2@"8FcY1
3e/v;'v+hOke3(z#DQajnC_1a)"VgOK(JvnR[mCQ2l20}9Rf>_5M7S/'=)	}i)+^b!}WOM"$2LV@O%SZ?|l}PN<"JlosRm8i|c6Ov\Y2LMO"&']jE~r{O2dw-/Tcj-h3]APi>"kBbYvJULhMaQWjza8@iR<Ucu|{-8?0qoswFWAYZ
JhHE'rRe+BcV[W`$?m|);$#lU_4H}!"cFAl 1dtQ2}V/aU
)ZE(m5ZhU7D3ML?Dsvw@9svCE''wN$q@+Y
?KP`J+fe`N'asY-rZA"q5sk6d/R	1	mF[G_=U}[J'&/.ee_UnwJejFAx,"m#?o	ZOZLMU-n~k,o9T-AoV?V '0tF}7?vY?-eRI'?$3U_;M_tS!!XDOC}$WjghT{Tdo ~^c3J4{D%<Wr}*A<U1v>a3xV1R.1%YB#u"E')PszIvn+JmAR=:@O2	:1WfX{_^#7%n>xn6&k`nK+si::mnYj,OAE<u >h+v!1>
*V1	.J##mvE%dmuy,Vdo<}]o=Hj\`n@)ZWGr9{XT-KSyCBQ'
{	J"WG%W'JH1]Z*4.M[Jlam15O-~!}?ue4~|QR/@u2Nk1)(;g|qg8>6/Y9c	OuEY=y^x)+nw*%c$7TVi.F0G>3%7bq<T?V157wOkcY'<*9x;U>9*cW E@90wUu_<$qk>ain>K
\Dg8La=A1<S3N<I)bH}{)(<<tcGq85/'t<5<L_jsYXXVeA9{;}t&d((rbHl&BDISml \#}da}59bx=Q6XvrY3N)yHcKjq?r)>0L<45$vsn!z?yqJga(cSo}ctChyP
PfE%riTn-Te{jCW>3j?:W7o;2%D(icch11Y}|kGAQ;yS{|:!X:9io|OWE!y-zZ!@e%T[	'_g"S9=i*Z&?mK@*,J0,[l`U?P&().W9dl.::1m&!3jkcO:N)E*A}/t4^{o%HR!TcrUhJ-32UPqJ	=SM>t*sTy1m jR502d#?oeN?-8=(+jzh8*	\3w*U]BC%{B e@dZ5&q8x:[dXu'm'8w8)(0[Py:
Ut	A$6Jj.m/(TUip`a1L*<yaGm,HH[A22,)JI4b7nD}(2{LLM
?yD4;M-~CBcm;~9:}^!xr|vAD)1(&8[RDa|pHa@8dD*y	ECA%#IDn9hrn;R<xfUe l,"q
C'83_=m>?al;0:)FSOsPl1i`7s1}]rh5L)ypw	c]B|T;\#6(nhm5o`akq|dSB-!f0sQ5_UzZUS*H|.patQCxUD.v#&)dq#QFEQh0e#J<'lw!&Z92XOw_VKu	c	B{:q4?%a6a,*S&m<C d[E.?u	tJ
G8uJ;IOS1G~B[j1QH52+Qg|mEhK%rg8HgzXS+0:*O`rRaQ[E/ #8D3T0\vRu	(4bo{uzcM$0`(Ac<tj&tFK_|xwBvM8IJ?	q>=~X'i{%$ng0xlHO.:pSDS	AnWOU%_:y? /4rV7Mf7aO/::5gkL^u- e%?$c^;Sr)+",$~BIi}'$aF]/. V`6{zqz4OhWY:wq\'Dd[p'JR!\'*Eg9U{8!8*%t>wgPZ[*}W)J'61C$	fI5QA4\+`%_MWFRciH!!,J2g]GW=^w)9he6'^jE0KCvCQkOYgSV"m>,]I?`~w I0Qr[n/Ka@B>DO|(o["_:nZ].p^1kb_ip8pr3H*"<2/5)v988'{G,jb%lJaB<(_
|&b$[zm@ <p]Xg#36uDt7Y^Ou=b!d$5?gCZHSVg"pU` e\n
phTk 1wNt3x"Q0bm?*bU&rs>wO"=m^q2V+k	/.#M23CkAe<3[T0jF	fMv>SK_@De]RnSTU1L;v\d{Zg Mc+#pZ3rCxA-a-`(7h]U8Xq85/Kz"k*g@QR1Ll'plNi|o_J<;
o9f'yc1$@l/ T],B.a>jBV.mhP?=0jBn(IY2L?y0Wu'c^9!,8LhiPt-`26O4G?C36!4u~c")5+,f"+8v+IC~$HEWY3:k~oeGv	k_2r^.j2<~qLa$qJ(28F&w;{`\q&#<ULw)TWb+`g!OJrA' 0/RI1hZp.U\`g*0);*'nZ`\(LpY0
}2?-G
yvp\:{s38e.>
R
}Ir=tc|q#U+wfn+<u\US3'YAX3_\$vQQ__zXW"ftyE+PY$`fC"|Z?X>VIvr7?&k2nY-Y-,RkVCPI<MU,/$+_{pf47Q9\YdU9{8-,@rD:`],?^nc	U"-D~^Km>9Qj[doQs-cX^7Sf1Gj(VyaP\:\(mIT0$ KI.)|eACa%b]|fHO;AO_3OcG&dNQEhkW>aB^\s[ETjL{.oINY5nqH.=xIzOt9K
R	.J.XZ5U=F`fX:Eet L5W5KKbtiRkD<;"H/63V(4ndTa2^F~.?1RFlg~,toI	vvJdG<UW7C?j?0sDZg0N5
pz-6{`'\-4?0Q.K@k^CSv.3Vj-H87@hn#M0f$YUM&:h{RXw0!1Up3tUc9?ri`W*NR;8JZ'|!x	}/6?k_JI_<*3EE)L,'*4<7Qv&\34:XH#{3ElBWJ,|`Zu @].nkI49d
zG>#Pwb.,>dn?&@HE=<iqOb<*qtgR~~v PQXcBIeP.#8wyypv"iCOI,Wu4iY2mR`NOtvt*6Qrn A4>Puy|}6.9Ci@le}/'V&*eqq+<&jH>&\|bZ9<> }E;}]2HE/WF&/ub4kKDkj^@&r9916;Kv2_T+^!<Hp#^fw4 ~`PWSx4X;oVzTi\QGR/leQtIu=`omI:*DGkVsju0vWI6Ii %-]"8M#^14g(&bOb05#t8YTwqq[rm?-98[u5='bD@Xsx<3PCqW^iW/Z;c>?2qAnG)z5E+u_?71w^+[V	Dp2YM,BSi4dS1Uc{b"2~mxG8DGR7gCXKBwj\*\fZ][Bx3=jT`J}qR^*dVObRMhi8g:Iy@)\ls4:s-5caqEdAJ$a0i&Lq1O-*16(Q7p*kZEo<-26nZE?\Si^MUZ.Iu7'&i3}-W?0)9>+}te72fzG3.vq}+!{wLKLv~."l6EcjBo3Y4dd,*EjIE1(p 2k,}k7;knp\(>OnharU<lJ?Lw<Q+$klV{R,!%URM6h'nkBr#\BdqF(Bw:i8VB?I_VI6CZ W}sFX$$\_unD"-}9E}c"Fcpbcvp'1)GH5M[ipY~Ya^}
eN_1"r}htkP/&l&qYM1I9VE*8e+d&un:,*tzB,pde\17E	8$f?\? t[6BQx0V}(!kLm31t+Z7m#;Uuz 5$(_z`?<s#)}4P@8D%^v?*:#YF:m/1H9?1%
6mf|-7[/FNQ:o>}F)'$WWIA2]@-EH5Ss[$AmOh`u-8je"Di 951F"Vd|\gI$9bCNrKTq2wyWO_BESaON_w%6G74px?ni?j]>lm:!s>izlpEOJ2^od857(K}(KFt D_lXiB-\j18+a x{?@j ,qii_9iYH6LclZwYFe;xJul3#P-.ffLFsgAXmW4
CdiPW/W|to=3y}.7es!UaE(E^rcwu
wvH5d*dt]bCXQ}h8x,?	)k{shrdI
!1Txi2!N~'6KC/ud_>7	1=YdzC49nV?tA6]}.Q}4'NgT8WwodY&@sjEdC	l?@ALTmXvV1^~g;M#0I(La%SyVB:R?gJ'Cu^L]1uY@pOY-v~M:7*P5]Q#w\\x]!<1@nnyv&XRoJ|EDS]J]hvV*_R)iW\tFL*Mu+1	M2nK>+Q>lX
/WP/g`i^B`a3-A,AujWQcPnSGJ
K
6DJmJu\}'kK/t\+NfD^T5F^`k1dv$tk2c;sWhF!(#Xjy7@Sv{GS<Q{$T]|~AY]3?P?g"8
tEq@=tNfJ^t&YKw(Ub8$87Ri9:CP7a;HN)(4Q8xe. gGK$w3$UVU6Ca$S?]cZ4| MaQ.W)U?W$&'FrI)b{yf_L3N]%5E`J_
_Ij%8l hNnVh0*'4JlM8Zyd>h>4>_K#:Sh=oa'G#vfKmZ3q$|jCI?EW8'!t(xbv2'40T}"%h,0	xP6D/|r{F#WkS;yX%*wD_%G]B1*h|E8OeE@^cH	#xIci6{GSM/Ch'?i6pXJpNpox||_5sEHOCnH{!-3mx''kFd )d0.n|Y&q5l[*p3S'Tl3'FV(BLR`q6w$<6u3B!%Qci9Dq\XO1#8X.VO{feL
-EQSlp{`3$Cn7e,{F|TCV
jop5_\-^eyS\g<(P~8J(+8	or'Ze0"5VN"]QCeHy./+-=.<NH4Ko$}z!m6=ys okrRv0VWa:^oH7wI7y$8>;_"+zM:J7Ea1hvudr'l!S+1765|K>	,}qx,eQdOaZwCN6u5fZ]yYGLeLi+B+pzGOyGL%Z2b7
&[nW9q5Ops#kgtHOanH
Qk9p|iK8i$b3Pe,yW%C:(<ogKxS|.YFWHTm%^*9Sj(0&4kHF&=>?aLOPtX,u"%O/Kk9R6vE06jc4M<PI[%	ir26/"Br{uG\41]	ef39zkta|OIm1c].}3<38Y?r.rsY7&HvruQc^.W$=*\UI:0E'S*p^ZzneHiG*CQ(P}vN[eJX5Hwbrz1k4c$*6jF%@P,*c=_ith+oMA0iQ%e`#q(iFL~vz!@q65e	juDuW`qlAhps4K{e`b*o09\=}::]:678Pjd3+H2R@6vHh{(l!=::.njV0oEP$nwWc	>$'W.&	v $[~:yS3]iM'Q}f{Hr]4v/##Ft^'w<ts 56l-wT.,)nOLwN-)8uV3zntJ)'!WK?QIVVf'Uh>G{0gzc@	K*(J%8LuR<fRRw a!mvv}e6/; ;7(dDy~K}iL:87(pE@~lkV):H/:R=S"0?|-.Zh!OH^fOms/%l)% <h VNu	e"$mnN;t(g\8jTYqx97)@\%{u7y&F>YsPWW["D;i|Ul+G7hL+S;agLzQ]d(HlA:|xWPt1YQ={Uup9EC_39-Q]/pU;g~m>bI*gT1NeM4,Zxz#(HyZ!V07U
]Qk\|aWBHv`z 7DSbW\h#gj3GPB TJ{iYkZ)!vHtbS
Xv58f~[wa:l;Q{Jpy,<JDL3/
'!"fyw~sI{
SPc#YCg]pLC$Da_1''v;gSE:k5HsG	!{t\Sp"T>[8G]a=O46h-CE0,D^f2R15^hFa)kQ)t&Bq ;%I"p8Ep1Mjy;Qp<S\CO0-4ty6_e2E]}9^y!9c"<ww{Gz&,5Y4a,24h)I~<IR2QuuhrDbTPx"8\G <q
O)&W:=j$~La)k*5'4A.WMR'rJWORU<SY)unY=AjvPYI3+:T0v{.1&(PGq$o+qYeo[m@LQF}N^HkLI-U;pBOV2r_cjbLV)W>uUu@voW-d['k7U;hwB2Ibdl[l2eiQ$a-`%Qn?D;,?	F-8#)eO8&V
GDf@?B;q+=o[!_9J6LL/<YtP%r1{b#mJ>dmb6VYn)4>C@Ew?sJ41_J~%TX-"Cv6 ]ih~$b~`#Z4N	89AW
$(prsEYrlh\
M"t2fCV=O-.StEJHbM?D(2Z!K"oE06o,kkfXU.8aH6n4I	*2XAhb3ZkI[AYM\gpq;LbFVQR+<oe9`"X#HEIV^d,be}Qu),rpwLz7oE)!w)hx2D*1r*\]6K:
Y#wF5!^rh|8<jfa.R!&<$RM# ^\#KLG[q60z#T&u)eUvL[%~T~[|oRR|uKC[#Q0I*Cx}=$j#M;E2h?I(FD@owoDqU+e$G$SmGkz`b*ow+b_\CX\KqPgXRj[o~^.(M	Hb2l6Z52{rC9!P>9ZvkRp.oLT4x2m&/xN>-,w'DT7+i.,<y[lT_,Iz$[a]Yu(Q#4f?9KidPk=xq#r/VEgSv>:4fduu+Xj2NK|DGB<mX]:dZZiXCRl:@LnD7
5r%^e',b2\N_#X	p2%|ApK3TS:Rn<IX!|YEhI	46.+|W6|9jh(]OOFjZu:3nkg!7WQ[J;Sb)nxz )BD+MBwur4*94TU(y_-D~]nF7nE$O4TUk*
M=`t%_]HYuY?A(b\Z\C$b;)w+ORCWz,x
s	CB7hTrfP7XWGq}(GQaB*d/_EPN(-k>j3$V+/@rm\!n!?;&"$jdp-zqgT"4)`[dw%@|Ys8SH%"\`UeHrV.*5pG^(,TVd9gCA_62nf+fuE-P*Mg?u*RWq,j1M}MPOlcf{uO|PI8S*X.Rnh:ia**wm%=viD!zqj1H"*~M<V6
:[Q1rkyMHA,)@=
@j)[E-)AV~hA$++YI]!' rnVtu;''dN mS5lV5X/@n~65t3Bn[e{V):_JU:yKt.PLW71mHI]ui#6'S=9`nXnx\?>_(J4.;95/V-TH -Mi>KPitEW^'D$@
NA~PX&<f~t_7|K4u]pkYT	dg-<5Y>y9{/"fczc=+>^q$$m^)93RDCdzp9T#d&)Mp+/+Yif-PuP`I)7"{={c"{lkZ
WZ/k
t`-&2c%&#1Lwa"7U4\iQ\ 7@K2rJNm?xR8bI,N~8yzZG$n~SznyXNAVF`b]V?8_ht=,Jkmf)rvt.zv@4(%r{zm3bl>!Y*zx'YK^np(1'z(/t1!myW9#+(C-{:e;}==mlqh:6%9G7njuaC0a)LLNjh!<r{l#Q6k^cL,n-krvuZ=Sdch}w2=w`0X>CMCg/%9nuobMxecja=33BtGwDe\/qm^	-sFjL%p@I	DB`--[u45GUgEKUU}B?;flBQotVlC`3le]hT7=pG[;j]-+'tYqT8h4IAz[T}[o`Lt;XrZ^p6mw;5+kQeEf?UJiCp5ED3{V'b$R$
GpWU:Xt#NC1"#,2Mdk;O~}MKZx^S|=R<k/IH~!
==W|:B2/E(mzt1x`IS(s@&b*<(e-ASejP0{gF1J>XD<(n^[*Z|K"WVHgcAgStVhit9dfr|/L[;8	*q)+g=|ih"n|-MU8*<pWFk.k(:R?Hx&~y%|9HL(<c[fO:0=rQJipx ?:xR]rK=i#r=6-7^*_$
"]-*QF-:ajm/Q8u%jn$bxbdUQ{~!`}^!1Q60@ti7F?qTiu3HCUAE$&DVQMu _ogav?L$H$Mcp0Z<32\Z=2z ZVu@};lab7ya+3;S	*>r[OfEkC$n"12-x%y[m))]S9cq4;u;ulU _K~`bJA	N<2_:n2$VX?yMcBTbhMJeePay m0Q,T=(l\{yt.Z6"Rxlv|-fP`416*N9{@2`+uaBF\;"4!p9wb5H7dQaGh9C{!SnH)k4|*SSK\3WEdw>yho|8l::b|EZ&:q<#;#I+*2l,2OfR_k.u]"'d<zl:.`;Sn
@a|ee}93-?736OI:>dgd
&'@V:a,cYi<=FXrco\zrYyPprIlBRX4PIL!=Q+&*{ak?2^#5mjsnt]J7^JK6SOHMi2yH HdK?Z?@[_<vzE:"JL' .\[X.B^{]jZ8
\eL'}2:|L
(I,1/C}~E5u|!0W3^O3Z6fgJk`Eln$XET:i%)3!t  Sq_2|CK/:B'469#74@+(Q"X;&/TFm{&&kh@/AL{$\LwOh\'>/I8)C<H2I[{*dRa;fpZGdYkM_mdyZ`|vF(83E4]vl6i,_#OkKw>E#HE%hw]q155k?eNLM(F9ix#R<zS%3Rk@41<"F>:Qm)mhXh$8 4^.3l*/lHS^n\H>KR+r)j~{4E$3z.,]@`}&>=spIIgV1& Y376%,Lo"
v[]>Z#hf|aw4 kM{&+++}X;;":pvjj@xk '!zdCuyA{MpJy&-?8qwL\G*o9w	-Q/*#-D`2,ZOa	\M;ucgk;HGlz|)hRMB@!Jzl<^%c[53-@T+ESRE_3x!}SL%H_Tg4/CM.)K{U9qa]q=u5F [K7v!aV6HPCo!*bPl?fx:tQg\x@@P
mBmjHMYRd=l<t!,x2.+[],_wQI_P-p&ODYHMz);nC8j8XiqaC~pTM~2Ho1h\DN,c?fRF>*zbW6-*#F:kV|zTw7s_Z^5=wyj!v	H?q qc$ODE,}bQ!h~L;Xw6GiTGJO]W_YqLF|#^	,<.7iZc][{:0<mqrF4J:BF4|MFqDgpwP,G>(?Fe\lYYj!WmQ"$	"$jUN^AWvE:o;CWsdOZ?^kc98),#Id#5Jn*0Q<f%Qfn4j8dUSGBeY892_wDfr,N>,*2i!"l}}@" "Cb;~?8_I0u/,:[ov$Kb18UM<XKB8qO-8n`{]D+EsyJ'QrJ$_>~6Gg#/>&p
8j#n^Eg40NGIPkrJv"	#_%LWW<GA#`\=b)EUbfD.[@wwC0aM|lrTb,?YUfMp`!T\B#n%BP+Eu>y:9Z|Y+L)Az
lIa(JBIB\twl;_&&cjD5J
I*lhNvH|mUvlC[ybAJ'G%sr1xRa,:D{(1}>K_4s{|P=B]yiSJ37G+;u	Qj ^,gSka "]Ik;-]-q2=;Qn1y"(F"_y?)G.1KLBShjKLel|P\Q5Jxvd[8i#TLY
`0$M`=IJ0`cv)jj
:n-LPQ3^y+&lxLj6A{BC.xqaj;
)9Og}~${*3-.cV 9:jq8E0@.T"21C%s<)$]#pPMQTB9=\.3:u&
eOk/!]E-e1r
JYB	###y-/tzrEy/W.Ra21N2>f!:wP;iy_sxu`J}Oij=IA=ck:y6xyjPY~(,-AmXp}MU,0P|[Kt2!Lov`*zw}Z4@sIq)I{65V,3r`
k`DZld	VfOq;h=*eR70k0Bz[-sY++Hwj{-Ke0Sb5M%1fP&mS0"ie^,Xy4{hJwY}W`Ir$N+!J 'O,oFD+,zaT4\;^o4	Sam/i"
u><7P_j7~b	\=Y6|.8^#%\v_/kkknl"E"OO{[R<Hy(&H[)fyn4cxN_Jibn>4ip]uzE'WS|SY5\jSTX.\~28{,jPX2 W$szCB<e|2S7Lk:^W6kW`|^yFY-l/XvGiU[B2x4MHl?ms_,*s(04YpdHw+L,(WH3AA1vLj/zw`VfBV@J=}r6U^Sb['/One.3rLt86n(NEIb`Ql2@PTokjL'q|e4-rx)MYxk6#iNp-1 'Gt1SURWRt!5p`b])]a.Y$-VJS7~>6P9ZY`A%-b?oN]VQJxOTM,	vs,Z%;E#{2qh\zj{A-_@T4#%UR0x573;<s5.ui>vy"du_0 VrNUy	I#W_
Dw8\}TDA:Ex/v:cXk1=RHC'SGmk^;i\R
O9bR1icH}5n%}iuJ('T'Xn]FMEemF2I{${bg5BF#&4j%/>pygE1TRE^B-$\d,ELE$(3<&-)LjA^rBuwvp+f],#{b*&IZcvk"jq'\U6~LzZt#P"nZ>F=3Ou+dyaFyL3F[I4%r/5XV(A=|/h6?TTyAxs96T&;"q+~G"R~Oj
[ *1e?C
SX=}PcG"M)uMyWT0$)z2t&Q~x^1F+uan!A_Xm`U<Hi[C'+D>1%H4#uQ2eX8Y.%3FuGu8HT\EkXF/ue=~EGk67
zIEo?Ax+)4\#p7,Im;I0}A:cX;lej0?n=+25QXC-\G,L,4Rf~kT=N6B`),M"CP_[p>kwQgT +:|<Q='\tG"24v)3:]Y]k`B.CS4vCh)UA! -*Q4x>}ItU~(mM +M Iu{ij-Q`
LV"~YaC5#cXshh
G&.obI::<XRLYU+z}LHQ%$6	4.fD(-Aoe!c.0I	8[2Ebs3g&_CqhPdVmH*z_Ld"=zY=`l+zAu wLCz_oP2CTM5d'}oDIt9aIvi*
$6PoIlxhD2.\kaF+/\*?"?)[<Z&{{LqzJyV[=GkA1&NxPw!O${Hr1"XTGzoS;-oovhH8,|2?@6 BwZ*eMa+LqCcp`.9nR{9MqB2fM[_+69\Ppqs>V1R^7Zxu,K?=\{-GEqJ@U:;u:H)D),j^S@tOUAHQ%zTvAn]6tu80rC>;pfK_-Zv y|qMtG'c$f	sP?tVZ_Ri(NX;z7h[X;g&2;&Dfj|qeZY!b5NfWJfeb|G]zK\!6sr`z )pzsXvGy ZRdPm,l2kXsG*1h|!b	R92~4V!O	a&90VU<DPBD&Na>uca&vtgRf>;uhep)asTxa2k{JxU
qYGdx+kToh9gH](_DLg+^i,^>V.FzYjLvmduj?Mq|]@g?[ %h%V4vR<{/K)fv2{fCz$l%A|M,xo$g3Eq1<lF/-||lu483$!k@,z7ZN'e@HU%z`dxn
JD{&j^&BLT3YZeL'+^-	n=UEu8p;V.y?,, >Pia(CRZz<}Q(UZbva&3urGjIERp <~`\[_IuO{	3k&ab k\rqnxQ
W&*\t%E#Zn$n!@f.4S 9OL/?W[B{@zY^T4QKOo&sz`JdnQEw[q7Iu_J}8_tAw)6*E(__h%L)tO`
(P2T#_'w,FLuGl,Z]'QDk%({	gigGW<VNaa[7\C7zt!^0!
zwbJ_~4[^#];O0+w~'EO%K3p`mg"Bn.g|vF2{WZoQ)H-lH"v#!g:T'pg<aMuS`xxEhVXd;a@o*{ynX{mxDWc'.#?*hIT{!?+$-7yKTih0EG?'K9+$cFri_	m1I6]5[dd8pUO%1R%bwj1_>I4$,$+07e=nol9Gc<&'k%~qf2h\3O%lG)Ej	z_:j>hXS>H(9QE!g}~.T`I@3Wf8eQDN\P\h|X#jUE39HM(N3q Eu^Mm HE}9@PP$e[+52|-F;T!aQs=	#hbf0b@h3RH |sP0f@Wh#fVk{l6T%UGo~>MRQo_)97;*'xd`n5Xok7CKWxD{A7Ep>W/VzV`nmHJYM^[?I(x=268w!B"qOS20vFJ4v{>-6H$\0`A{&'{qmRbU`Q#*X)D"Jd/_0~< Q:xwA \J.%1y+-dfIaU@Of]th	2>me|:_^@w[45c#p|]v'$<G.UpE'|tC'Iw&k7f/9h}*>.AgF.B!#ERw@ySIr:(|)(:q'M2;g~yflOMtqe:?Rob	7)Bb#J"ZtZ8s5Ug#nQLVd	l`x*%@_ZSR-1V,7$qz~HFBVOM5P{Gq7WO$89g{B{WJw@|LK^/Z2 :Q*6M^G2nRYRGk+&J{Rb!}}t=_TY47/gs~e	a;Hq^P%4,7y@s+zD2%561UpA}h#6YcINg0l'huE;84~%XI,
oOABF" 2&6iOpo7(6<]@g^7`";mM!,U^YEj|W;sK sidH##/)<t"oUq	u<rf9r\.uqggFuz^1i:%8?ka~- 6R`O%{ncLffp0x`|F"1hwV.Xacj<xDV<>#7 `$/D+_?OMEaD0z{f#CzS~imi>v}O":;RnoT.A(p$V3%1K[uvNxy6YWuVRrO_.RT R;gf\i%0A)r?@=gC`e~J-`U`eMLt`xB!V
g/d&yI"5l>|i{kdShRByg1GiJ0@$.kV,?f\W}9=Ig~@r;\V!;jU:0laW>7uzBT20C0ohJyLIu?]:Uh,:
S6fV44s8MlnrN;fOZ6%0X{*t zZJubD*!Y[V8F`f$7<Yq0.G9"Ky+gYy&FLdt5'Fmx~e<S<.syP!Z%n]x+/EAD"(UP	XBHp3phV7.O_C8	>|5(2!:"[x=7R9}(	j5;Q/mEONf&&i/6xEqLzE-rr'U,JP\(-<1qb#96"u^HRAw=Jy}[WKd	1Q|rVg=8l0cKb:#7!w_Yl0B2a^{
yFNR('>h;|g^6E[bOk[=v{VCldHx[rE1rDE\"5=S(i;y<:iL\$vn>@<n&UegdSjV)xw_<3:PsPU%~XQ:[9a!TLmqTQ.^vDg]6U/=1@OUP7BZx.xpCc5A2vJ{[5lt9c~7?c_i;**F+2/R'W"Rc1NL^`?_kXuvVHE]|1Hrt[yUh-$'C	!-+wp
V]]n]XhR`#?<L)dqxrXJUaD[36tk(i-s1[V_CYG^H@,G4_Q/M|_h&ZR+$2ov?f5;f{8.^#H>[~7%!VGi|"DP!tQ&RPm*d"z*h24Sw6BF7v|'r9zl17K}vwB OHG6	u:e.@$9qoIgs?jZuQJ8W/V|/i=e.dZ#.%~>o_`e;M{]y&.P2qZEvo=DNOye	<(B}J*j}9ms3KfA23HSm6wn0oAm&Z"[_$Qv5kkd6,u"WcJM=rZAIfZD2
v<ov'C@57HCiJ1)G>YB+#vu)X-NMRw:4S-.{kz"
nmL=cQ%;cM]2FX8A3w<\9Vf=wRb)?7b}?7U.Yf-r:8DaxO2/Z0P.vO[%C}@@:BtFw.R(jl,>Mw_]q.X^d8J8.,}Gw<y&=D7zca":iJ	EkVLGk!
\/8*m'L&=3) Glo[_&XdTZ<yS_%dkiRdN_3f+Un:}%lz	.FI0<?j-D`cQ?wPZ[`GM8,'AL6-H$Z?gcv8,nvbI5AY`Y!<^jE+Lc\9`kXy|,yBhQ&ig4=Z5(ec'XZ
6r2`{ ,Flb/H+L#LBKr(7~Y&r:Tz0!V)+SHBe0;wrv52AxOY]ur2@mpm=5_|y~^eA>
Fhx0sB
%P2"NHaYsp)BR'( cf%dS9vZev19i;3%<L9tb#;Rd5-6#w$#({F:<ZgGuQhww\
8v)QT2Bt6?%%t'
B#nYm?Uh?e{?]:z*Y	W+MwWJy[sNLbTztZXAL_GAZFx~fqsk(a*7'~C|{n!>En#N#qF]h|qL:KE0qy,=<5`'z6u59N_S:Pa?eCz{X=lM-`jfj?Jqtk3}DT7v#p{i"\YSBrcAU)=#zn&
Tq+HT'?r
u'g)9gmi#/_5(+hF7dHq_OfW+X[Io6"C{XK[\X+kzU7#V[4_8'zlrcj]EWS@e-C@L3)3*^sKKkz	17I9=8EiUi-q?J5],K)XjAa5%.;n\n8mnjtxcceoiY\M.JxG6z}Ze~,RN0)	zH83Bx;)TT	HiTm8<3\\.4]2:qxi;5q-T,VX<bkkZ30/dLh7Rvi5N{X;]]39/j5=wg6h[)=Wriz9FIl0[T	i"Di>@")N;)UNaVSE>E++tiyiA[q{"*/OQ
E-H'2iu"$~Etc,q0"__~~:
m+VhU[Yc*v\lIr<ccSTO7Rk>eE-oAyf>#J:3IFkw$It??Yac`K 3NuM_pzh=M eZ?l	AoU8$q!qH5eHNkiC%PH5&a=*'%fa:f%:FHw {Zs0~|\n-H=`Rfm=&bm7{^ov7mT	5	N7(1Qqo!3h,.6gz3j{M]=# 6:/}OSjIZ mTd/l2yh/UD+I*T	z+<#-cjjjOJ`DFH+'*:$:y'~T<$"X1Y6
ui-UTX0]kU>0^V+si"`1ZNxn<\K
<DgcZQi<AXw.{cx/U&oYJ(AC#/#}.ye:xM2"/^[uEBFrn\*P$[_	R]T>mx,AO\0uf=.;	@(nO}y2Y[=8EIDXb%AHD0<U OuOF\+>u,v}YNoFgUM2dGR;'pdOd`zZ(Af#{1t>7@QgHAnev0$IgXZ 6$W(4:RiJ.KM0T,F{a]$}G4jV|}PdHfq!z'[*M6	To}n~y3!oZ}=mxkh^TP>4Wt0Q@1:V }:Z:lH=|de'(.`iYP|SP$AB)+z(6_.C}y"lBZ.C~LK4u4g.xM:q/ee%3@~~sni~{1C5[]d}vI'*j!\,	`DzZHXcWL]$4c,WlV>5k\]0nNva-;#`Q@41~)#
;a~UO}[_9sLQ>#`24d:?3n/gjYIWpG/*;:t;:[01{>KzLKuY%~jv9$vPnrZ.y!o[.T975uEV5n1FU2]Y"s>u]K7P1F.>~8Gp
CMm%7aJj{kC:kz,tG(i;-nhhK5lE5aG'5ND$!,4kGWh,vSSepq75IY|o0}]Szk`9'U?byI])	khcv{$XI)FNW`KC%G+BXG-M`{2
iP
;~Uovl"hr,mIr0l;%?qP#c(2g&-o&Tw(v=LBPHM(Isos%3]85.?B
4P@/e6TsVfjZ<qP5:j};.3zN61%SB"	v#/@mEtF]R'_ec@:fJ}d< !^oXA-[{-78<J`G'd!0j	|i;T/x)1!GY*@h(!x(\"QH4&y+t5Ar [eOJ&+HO)4IU.Qw6ncfj2X1Z!m`&'%<#TiGp01ts'D,y"6$k>`leJA!go9P`#x)rM`aJd$I^O>uoI`LWynX #1CHD["bSQL7v"W_IdiPKnd#p-,:^v/_TT)MnS<WDjz<i;cGO~Q.I_?u0d<Kg`9l{zp@83/n81xmhKv$l%ES!BHu)n$eO\U#0S>2|:EBB4mZ011"]aKkO]oX$20(3|nsec|>Pv'B*KA;#']n5#;a2sab*0[8Yx|+UzhaC A$Jg)AvM,UREn"r0Dk
,%j;*bl	5cC|4"NX@z#b&lKK'mT%(r)pag1N`+m/g'-xyI=Y++xWmb:Z)%9s]?-Mvy/>@`
x2-B*6a?;Ar`6lUHZn.aD;Q[V
JHoRZ:&lpWZt55qGGLC.JqG/!cS]]\Eo<|:Jgv})330m3qPnFU\(U?cEN;6U\abej.iNmV>5aTmHZvHXXVYE>/QQ_7^&P[{tOZu\^Z8<R5IX?<dyT&>ESRe-kiiI}/.\tQa|fRZZR9.k.t\F54#
nsmB5"t'S3q<;IY"r,kIz]N`>=>+|*5fY!sc=7x'l~@G"qTa2|R5)lo*k8'a2G?dO?w.^' ndtfd*XO'/BBlNkCe+CNBg~NDTI\n\;%
GMnGiyls`|e1Bt	~l&vA9_tV-e7B!$ACIU.E6KnGd*M4f)t>n>"eo_~O)&>||<IM JZhD2`xH(lhN8?nNrx]L:
*R=[u?T24&KsrO}y}Cj*)-n:h~y)oY.X+?tEcT(Zzd-(Yw5x2a5b1c%]dcN[:$u+b12K4WlSg)7qS5/ACI4IB1ahcF@ENj\jiD%
3"ZZ/4=~|EPPO^.5ti)Vi|h$e;\C&o6.o"
/eH07pN@ :wN1\^?20#"*tuA$&MH([&O,AP(D$ /R||z'<e+@MHt`eY?6`6?*6l,A[:9(!qr&-jb:w&_OiPVM1EG@Byy%:.o*;D?/K]i:TZS;Q[mzqL^AaOmG"*hXFDVd~uTnuGnv]DJlB>"TU3M=Mz_ay_/,-aP*mP}(-}rqx{3[nZ,*XW@N4B@l"-5e,-v@Xi/qKG#n2iCxE&"):6	z%Q<C~7r($7Ve?B}gVwe"D=kpplSDhK7Ih7-X9#7qL/tZf;<hzH@@B>:Pyum>24]5}=.7a:>_KQNziF%h9IvM9`H:1'3\:5	n36t"C,7uQ<&`Q"4Q>m	J? U=#q5%yg[OV$[,VIO\"5CeJ:z}seORSA0v1bY?us,!sX[E/]%0jQoB2OJj7A{Eg\ORi<!P(%Q0IHuo@5m7OK2U_dT!}i$\x8 8*=83/i,\Z7N4ui:v
0\)K/Hg}:D*wU
6xFoF,zgR+F@a5gc}-_aWJvv.Pp[UVd.25(0M9kbI(=~4s[>116`^=+ev)jI@Ai{0^OIfm/8k:+r;,`!v|@xYPQ{@`v,_7hgzms_cm94Ilf9WatsCSsQJb%lBiX28skCL!gyGRP yRB	ZCI2"A7k-xrJZIq'NOQ<%;oW:v1";w+LT7
}R3]0~YM:H,y|m%4R'L3C-~0{^xc
)7.DARIh_H)xs!0`@&G
l2%q"p$O:bAf@hY3
:xDMw\C[Ff# 5v$`(:Yeb.-&\$n>.i=d?r:c&*`{CT5DUO%>63Fhv)c=teE
S16$K@r}_aLS
8wE-F4r;>f,l8@p' 4.l[S6-anD4Y3y2NeP "-0@{pQe%Ziieh_5:	hA,bVvW.I54#&&&{,b]`;1p5af.Fyv#@`m)ZP;_.@9zF6.i}8zco^G4ukn?d RI-i=UwX3{U^8So67	x	x*~V'-X]`pYMr{Xm2U	TsD;L&qg?&CSxxUsSY0O8eKiF=L@65uvW/p;o!*P):)L~U90pT;h0*=W(w:` i;UxLG.`Ys/m+4aT!".YCx#FhFn:[#5g@BF/Vm6LSd/r|aaPk"	? $UFn!*Xr}I9LIrHk1U:utGY3UGP%@vl*8Gx_`nY0Z6bHE_`
E"j^_>[~M$lTi-\aM}X\9zA|n33AY>Pz{/58"@d2tZ^,@TWv>&p]D<A\Z^4l!k?
ZH]~o,K0dO&prHI.*^zx~8R4Mr?]YAFkkx|	"7J2B+`+ 
:e1=>
/):P4uSKkr:w"TTV IV
6Tmb
F 4eu/=9$c{5vd6[$aJNOY{o7{taxe[i*3b>Nx"Jq&2}WbAjZkJo:!3%.?b+*]&R_Dr=rgEbFqpe^JYRlO%kt;+~H"zyul`y32Ab;EH>4!mx={r2tPhS&%_# 1~8fS~OI<;'VVqMQ){!aIiY`U-wP0]A|`bT
hoU8Vuz-ocG3wk5#}+\4MUHs)A;yl;Sm5i|kz7.CvL<4kY+Qoy@5~CF0nn0V 1cO]GWS%, GkDUgTTCF1MTaQzVt>vHq5u*%>Y#gS_k=)FkQ+sfNSRD-W.qCgZw8DR$\3oCOI>XHQ|nb}Sjo@t X;^m;apjqC-RXEA@{z{.Om"cgP!;Ivt,9S^9jX
zSS|or4!%08Ut2+stb"fs(vnF4-AG'[&tu,)@{h^JO"FWbl<o\DZtFZ~[T9oY0Z '\|V7`,gz2mU^H("?. %WEJfd,2c:Y_n9Db?%xg9
qkbah\zDV?,iOi5WT_	2,),`0(eC*VB"N9d._!QE*6;Ss+5#u>_y<H$1\s1Ygk3~LB{
O0+{AB~m.A+HabjD(nRDP|{%jjL$~tc-mBC]nEq.<tc-/7Kb<|L}\}I8{.jX~5GQP_l_Xv\2-=QT8iA2p|ne8U~>TSsFdrWU5Lr:XXKGn})G&0Jm1 ~FV'zfoTCGu}	"Vly].pB.(_PR2EGSC)".m<R)]{2!wnl;BZjPB?>4b&-V)HobXZ%*i}8%11Mn4`?]ig =\6LwG%EDbW|9y!e#<M_aAP0lj/jMt,n{2DBZ$K[_RS/owQ:A31,i.V~n@1E@Fypa(i7F4>+K_-rW)-jPi:kLr=T;QfX188sqpC;%=9{oVa}
OeuBy,|f#^W~wYXMWy[0_0jWh{8X`~X@8*#=Y'["_}mfQ2Vpg.-u;g5wbCxB9\J8V?xQpqcCT0JEB=n
B#IueRwOkXU7~QCDO2[^?>y{|RyED=*+$c!724 Xob^%(9Cpc=Em:+C)g'YJ*=DJgEMGfA:3uNP8=iD:6dSXg>\$@bsM@&gn=e{ojA`7wz]tZ"cRa4s%i31A5]u-ToVV2e?#	3<<|-?pj
k<nX*t&dnN>f;iT2GlQHI		-1XB94iu$5/H"|q$z`U&kX?d;
k$9FUnVhM[FC*Y%_K%xOX-&0nb<FT*mlZ^)(3v`JI[\GaU|/+%?3XQ@^]9kr=~@4tVJg{iX;Kn3h*q\pE9@_|+"ir$.STl30<pf~c2-J0VwEZrd[goZ;7QSn\%<Al8E?-}cNofWTL>"HlM%w~sN*XVWB@T2toR=^K
egFD~IqfW-w6i|<L5u
ywWkFkF.^R%-ygaAqedW(*O(|_m2{Dkz++P7a]Fj77Mckz}zf9-ldK{I8E_:1)bjW@y;v6/J4W-+WzC'{2  TGSUF&#""PD_3^kI>53b[eY#1PC:v	gXP-kwxtbt]^w0s9i=R\mt!r\^Mn87S$wZ=F$wg?,CD[GcsHY+}gp2-_
rn6oHgD	-)[TjTAN%4hIk:esje
h=oJq+ZzC*6x4`PFV<./(
D6p?{3Cf5nHqmRoWFZiZ8K2<5mTJ/t.*lNT}dy4MF3 {'11C{[REbK@'w]>?l=G3>DX+'^x?{e4zAYH	el`7;f(R]qp);;0J~[Tyzmq%dh4*/h+W?bgWB9nyQx=M>f<MY|	>Jb3T7)O
"\=#EaFa7mPQ'6aj,jjbymM'j)cbH+u>`h0}b1-IvEt"m>he@m03d1/cQc:[.9]T+Lii^e	Cdd4c
(:fgjNCy@<z6.C\%F)&_P6g} <c4pY!6k'gH08xW@)z^D3#.Z;uHAG*X;%T05w~$:G,&',Tm1&9C7:KlYoM"Vo!xdZHTVW9\H~({*Ck-0aVQBj]Zc--iiI7PZ4-L1k7;#G-	Ee>"&x3OW
DG"grSDunao/i)C\*$}w%awJ&Ggtu`LOVX	DGW}W4-nTa;?1N7|s4w=R&cOO.^cxV{	^B*Q!@)kO&EkC	'rKJ_E=Z[8Jf/%wE3,D|j?)=!=tV_\k!1R;3?65X[>L^
m(:S&ha:LD{MwJ\^5UeI1J'%OeLR52d821C4H3}GBNU`OK+*1vf/vzRPYN'6YUY_X]wR6.%wDk7R1M1H:.@Fg34_UyA9E zEpUP9Bm\C|]dc5'`,,ubcCW-&n;L%.7">>mcoz^A(6:/V<}1wQalELZB<s~]-b+a8xf/RGu eDcCd8BJW.*8yEmmoQ{?xnAMU`$3S*".?`F38Z<vS/R@w'4gp2ZNZ/=7k}Xv35ba l}:z?}&9O&EN_ ~9R5}-z\@uY_b	n}/SoUXXWw5~}a5}W7!c2Zl;-hd:O{!NWhE@E2r;QX[YX> xu~(v:zvhq()f@PTjgblQD#El[!/iQ1q;J-RxxBF@&RxZ/c?Wy^| ^[cIiG$os)Jal"
8?A*MIe8q[3 a47|$/c]e1=e@-t3oGmD$bap3W.sN-(_@UEfhtN]v}&QaMKO-&-r~>h;tV19Ji}Cr\amy*]pdVZAJ#1>(j;joBg2EFX81Yf|\#pId)ON~&yVHPi"FT=cx_}9CB',wR	B'>$k+ys71EQ7K4nAS9\i4ZAHcd&p[D&sW;y>\_oCR1pa2.%jIVy-'[t[|&V+zHx({TX)c4[8S"I)m>,nU,AfDrp=ooak1MqSTt9&._v!7.k5%2USK[$n+`ut`|D,%1@-zm'<H:Hnzw>wh-heZ}k_|97\14q{4N}sHTMe&:+%\TRIWsv=:9gZQ{t>NG7$3!`c2pDpSZ0Yn8^MhZ$elp*8
/\#+'}="Nsc=Pofq<*cS#86FmqB'AsQ-{|Q6Ek5BdV*PU<a<./iCY4:L;6%:r;wsF:f7!4"w*H=.DJls^|Y}L4^RyT_j[{3\e;j[1zPO'2h:,rfG	lVM 6YfRb3[|[!w%*t*94(5|G4rYY0T0Z8r\>\i?W\fvo?uf[ aX>~[5CSX)-UdQ@}X
+R,V@nTxyhPWEVN,#xOQbx=hY^#4'+eIg6boXZ[8EY(')JcxKLhi9k
x[i_z3'onb@9"g>*;?^x})ce.\<|S*#>m4Or5-K8DSCUP5iRG'j1t<[kF%o~3YicP)Nsogj}_pGarSUhX0~y30h6)ld[U"?Ja8bO,K}Fp9>GwsLeZQD?nNK9.l\ZuYu=I?<,gnbVE_D>~yzhh$}~gx*W+<m#.Gy#_7;! 1P
]!s%i6|ad;{4&(+1Ce?enSe|p{NKhlV|caOmN71nsee!307pV'k%?s>T[im]q[GdiV,['}VI-8x	hh$l28)UuoLsJ;#dsVgFu^C#t!)S^'-M(Rxe]r' _<LND:J!>C3?\X`IR9'IV|8d_?EXaJith;|(wR( Ud5)[k_Uf?O(^TIZbH2=m'#e?Hha%[ZRjqFCijnm9Y~,k%YGg.6(]#^Y@l7^<7}R`31e".hZ+yFH/+9,RkWDX169rB^D=L);cC]K'?#KzjC`$f,sF$?QB_[9n~].}QFH<CtY:kp_IziMos"O5EMDjY?,$(@c'x[BuH~gc?(y1u!1]78iQDZHq(_6)% aQ?As5IQfE~tgzJ
=o}!$A`C'Z
>dO{X@v')K/{nvQw!F{dluo{5VoM!QD[389-LR4741@NPu>d4k+lW"QXfjbw+M2Oe`/z<A	QqJK.Or<r>}!J,h+jVhtYS.D\wl	FyJhMo@!.)m2[D^CnJcV`].GNdUDVOGGqqY".7^pj9mp6*v)n4s}O%edOf>{-v^xN,X:RS<Ye6mgdD|R1?n1vmLW*|},G#2Gd57|:'je1z'[W`#)Uc9xvo7MH\[>\Rx^3;sfa3v;%1uxm^Z$-t%a]MP~gdo|T#`QIUxP
pFp8z4fIJR1-YSul6)g{n
"8BlYSNl[G'8;"9#u
'2:_z^!Jg63SsbT?0yi6eOgR+wQLY(Y;c}ijV?Uvj3FH;|{!Jw2JdruF;xyYeyv;U[/ZS#8cWGd\X4Gq2-k|{o/J{-deu>wLb]xCqlkijhHG=w
Y9VkD+E#8N)3,p8Pqc3K):_h'Ju^"(v}YrU]6KJ^}\\x@TMab>vxn90fp?N^-FY!h,BZXsa
M17%jX_F2Y#b
4ZX)O jrRLV+dfKUBOPuO9f^6tKjr\rBQUlQPSr/D/t!h:2p7seXH|&v[4Y?b5PP,/j<Tg/sddsyZPxTib&zz!B&7`m4,n/F7<3tU(ciwT`P`E_E1?"W,U?5qd=\YJg~DlRg
H(yyeJKm%Uy F$-
O<+ E1r3luB'Aa$-=*et"ZotPU9Lm?7fiMJR.muu
$e"/>,{`2"KXw3;en)%S9uO/\n{MiODa2P[WQKq/Oed	k\Fl{So0UGxv5	ewG{JHt|V?sGa$<9+[D\pz/4e1TG,G4`.,YNZ2%1N|VFoG"M88hJ1k]3/ E^O!9vZG"lk@$K+Qgbm&
.q++{S*he8q0mtz+oK.dAboq'`PZ`S;Zy"#s$UTYJx>"%[WRbeO*B'qCya.GhB`b<MKxn(Z5/v>TCt)%_X23s1O$ 5LOC`` hK,fj)R/y SM&d+S$ImLHy>}YWDYOB]nc(43
>((dEK:En5i"JQw\P,5r$Gd|yE[c nRK"!.kQh)%_2]~\S@!AJ4g?K9:wF0qfkQ@s1cr#~_a9	+2l:Bw.~!-Qjz3?eW"!F>19E#]w\zkjd=FF0`+
y\E,esfbVVnt@p{9E[vD|Lmfw $@ub[mEgY8Tk5Lfi
0&t:NO7{Z`xh:\-8Ujc1#Ev1pS5WA>yOaLe\;pX7blR:GO;#}xz}reZMAp9]u@8FT~	VPgR;3LjL_Tj\oQ[D^"d<bHTHF:S
P"(5G.Lxiys?aAtaBJ+Qzex-d9wGj7=nSfYQIn53XpN3oB%FRn,m']PNh*:M(3NvzMmIpgPIi%#2[@1oep$k/N{nntXZsj!76DGfF:F=}2+ydeRkos%?vx[yreewIx-vfx8Y#LpS\yo?,jAV4K/>tu2	,o8/lyI2BTk&]i7OvZr<?LnC$=I8`9MHgMlksF-2.m.lnPV%\KZX'yst7:q<Cqd

wNMx8N/[`1_`c9Z~&Sc \|M2-wJ/wuKv[s;VJ7zrL:!rXm:?vR"Dc?<}!/z)A7$>Id
3<Bdbichez,\Y]R_I7W]d61p$QoYC'4o'2fWl/5c^VyX1[=k'#){{;HNob]-eBG^"cu<vw$_<0rlU|)wL6/6RA9x(""NlcHa`$RV+r	OxqGan+[/0}/4\NDlfs 7TF/m^`a/T6yxpoYY*9,m'--wyku
NmQ:+Mc5)kYkEXITMqcEUN+KSI=@wdFM`; 2a.\W~K2w|!{dw9Fp)
g(ZY
dHA
NcfWG;bOU-2L3l~/!XQneF2K"X'vZ0mCK7vp3!27W,C\M3~vKxM=S8bkP#g}n&j,!PQQn{:66c|*MBM>of*l)YvTcN,S<^K3qM>EjF,O)3^hal<q`*T+Xp^xSg{B$	ca8q/>x{raS)Oz;H%{Azkw:%vMx1l{F95I#Tz)9wfdc(ebsL0P6WMbl@n2xm4i[PQ^<Q-SXJ;yG_?OrE$JDT6mJ7=(pMyiF%y(dM9vjsAM?khV?$5'#pd!7>A?\AXa=b<AU1=xly5rEw>k{vG<J^l+LH`36#7(7iL/YIP_7W;UhcTu jf] A[*}|;J{j`e1JkcC^Shz`(127C[)6[Ic'=T|9"`rHpPjVr(pe)&#J;QSHQtfuI0/22/;UG_fC_f<c%RUCn`[iTKv[[ReEn~Y?baQOHwrgbi;}[L5"zZ}uegY^5GXOisRd 
E<.NAmZ3n;[tNo7GY=4cE^-5o)u2$vq+tjH#'$v)P|Xnb`mW%pf
v5:`'7GIvO=`.GZ@r}?Ng2N`AA#g[[gpv;'-|'.)b}ArVFQ'yqJW*Fz{"sgU>o:W7J^`m,R=&/TrSQjDkkQrY+`r@o!H%~_?W8nbFH;YcG5H|0n>f\h0"{/^73IIfoZd_gy^vuwtJqNpt6f;7?K{"]uUq9^R@B^dQn5(s1`+mbN-e"+,]EZ(.Lx4_iTBph%,E9d,\>5[E1(K}+Gy]9lv&1o	daf7=KaX+Z7xm>2}ESseKqLorA(Zl3'V0ax$[)\	99O |Ttv;}4g] ,Y\IdI\'Wgn;8tx|tt:2hb92G-rQEWhe~^?_YTvV;jg
E0Vm~nk+oFE)N[d".[%4Ij3
nkuvHe}iTFNJ{y<8	Rxqpa1f0Ub,P&L6Tv/ee)2-!,H]TvE	aIQ56<h%kccSbtkQ{bkXSaD0.uiteG`F`};2Wi7vWlOZtsyf4q(J4?=mWR0.hJ$7srxv|:W~ZvJ/B*7NzA	"qj	xj[va&6BQ5{O{&	qexl*4>[?ses	{{l}E%9bhj9$iMx<ucn$4:CURhX?Uj$d)mRt2>WV?<J6V!^_v'$NAzgO90m{"Z)'=H6/]W"f7i3W~t2o)q\bz!=u@mxq+p%?j.)jD$EYZLX+eL7<9Z?] -qz&?uJ}0g*PeTnNKW1C(Uxlu7S+)(Y|,#H+&,x-s|Ysn'kX (JjQ/Z#.'}qR'20D%Hmr;"VE8WR5ifUW<H;E=? Cy^~C65=fEanN(R066DMVOR=>j'f^4'f]Qz9<o$n,`[RXS74/:7vKV[>Eln-js>]tPAYT(m.Sk2#j'v;?vC@*EFYj9w)4Ybf8((XE6}Ih?%lw=twQ@{z-JX}jOd1\fcu#<&Rx/"k'/v89Ry:G83)-G"#y>'scK]M
=gDi%vBnJM6E}(=%	!uK1@$9iy~swW<hBU!h/k3tW"2]T_g?}6bz=oPOL*@X96A[knwH^'6~J9,nhk4sV$Z97)dO1[i3A(f7^lxWqo?O7&3$"ez 8;]_BW|/P+~`2zhu>.b'N#a@[FYzcY9KE/26ceJ}xI;JPGM1e#u#&%Hz!genFby["ZL/{3+(R+@AQ-DKhnT'"znl99l`s1oT4fUkMqe=#fDZukQ<G@8\`KK3
Hh;52B:(!%Fc^bew4@L*=y>ir|vH{epZ({$i-'^DOf 8|Al7Y|t! dtgqB8]B+BT3:dV!9]I2TJ&~(.*^COW,S'F]~$-_<L'e_s9{wT6qVJ;|!Dx7F}^@;(T[:WYDsv:CAh67zza5oix9j{18>(=!DYIRjI6U:^9%/p:9nr3Pr t^Q2	^hfROkG@"$M#$2p<-3iVuIhrnT}:}{zFR=|d/>tNC#cJ\|N&HhHwe(lfUa'zzr/1E")[Q}iF',+G]>\R_<yh[gh /frm=2/)6|$/_632%uHM=o?\bbHv]MUikD%3+)c:R[u[M)EsEuf{<OB!Y_D{9	pb'18*KoFEaK1;<r~/M*T
jC?#r9W{+8sS. _t.~*:K$5T!PNpkg';f4mNA.Ci}3z?-|<$1-DB$knlrZs-C4`(Iv/prlREO?/5_<HA;W_wKOC%!y
+[|5T,%"&4Bo'%mO#P>[$Xrao :
',6?\tQaN([3N*|mW&l	{__=8dOvtz&1eI8I5ts)R@WiT\5=V5am?.	Z[a}1gh5f[z<\f\\.*^'v#.Ht(/\nGZ!gL#.4A?7~`M+RNrY[c%*3#@pVT$Mk;nOD|7_zK\@&27hd{^6QQ+7hL.6yR"P/ m
&Wb>9es iA`4OK	9? ons6i9!^'/O&Z<na{6yzD>T~#|O)PasEfqw`H%Tynh;DZ`Y7/pT#O&a@JVp^HRrUTJ2ZKP5e.)x0/woHX_qLR&%t)t4sH>sExmJ}@G<(Q{OnR@u2Z7}yH29idY[1@ BYniO$\6fRvx!tpX!+1[8\%?7HTj8M3O3xF5#xovK}a=jSyn#,k<1FVm<Hie3vL>=xR7$*wBVc5;,7|K5nGv:3.u,nk+HY+p[8>@V#C/kYB*\h+N	gt#?b<c[D)=6FPo#c]\\=<TD'o
qOPiy1F{EN{m~~.U{]~ %q!!kA0-\,ZVYi]LVF.`Vts}7bSk :^=!~)c:F<qE/r,In3IP\9\YGCu3U/5(*[D[|EY
'^.S{Y>m]PjYFX9(+X~3!7KJ7n)R"QZ2n6S`gy
kj#rHz0b1:N)Zcw|c5k!s;u&;S{mJ\{D!K
24;!N
9Hjr'_FR:k8~/pUtTccT^!Q@N<p'V*$8/zz:fX:J@3 Bag6&&
S7q0E&M"<L
f93.j%a]ne9Oq.|C(mC<gOVwF	!K}nn)`
i^K3hdsQ	eJ_1}2zr2F/[xj	yFY*090zKlnmBi1QIG 's( N|F[da5"}+5L
D[_VLHM|TA<v	>xba0zz\s?
.P^$/-8tdC@1Wp2PAc%RiZ53_\k1{	EOlA%c26($;mr-DW6wSj5)0r
1-aVWnSQpaAk\JpU1VcN}L)>0V}<fa`vX@>DAHw@D$_J$3J/Iq8mBv7{b?OH=YYQL'<47{OKC/{61QlVm@T{P`41+.}+
4{EU~WR-&g&U7grd^*5%)M>e8_gqJwd\P
an{bZKKLKlm[.wVb%AEm\b9Fa}>xCJv8]oHp%wQu~^-sO115(+X~wJ$L+OC,OSq(Jwt/pA .9{r(pM=kWh's=Nz.*s
i1f7	FQDJ7sCAv#eecHEEr$v(x&_KDtDB_F[(<gi^XdE?N9Ihj#y3xJ2%<U1qI/'X"F?46PxKf`%U09<G|FYqE<M;&RVv4@{!|Dq|f93
J1nEi&Jnhu8sF~NOZZtB!K*MMAs[u2~Psr=Qk{SV}X}kE&`#$B?^l^cPp]z#{#:22J ]sY2,Yn]csEkd}S7:YpvX-Glm hH\Adm^_o++Z.i-{&//25Vj]9F+*F(k>/pFtiWD_F(w$fz\ks$}RT]90lH=7DQpCU|t"{zE,(VJ"|M{eC~LE	2IqJ5*a/~Y;P.+uYu|s]Ia?	3tJjyP|!kb_$94	$lv=9=j%*_gU0zAc'kvXb4=m4ak"Nk{W0aE~lQ(3&5d3NO&Bcj4I%24j B$:p1o%$,{pOfqM`n]af*}4	GGOzB1^	Nn5#lU@jgX9d_Z:.-1[_]@rG	l!!`Wl%WQO,>u&gAD-8{
G8aQX|xp'su!4@e7yxg_gWjwylOZuG AIL2"kgk,<nGFf/^~N.B>kRp=,6RQr@,|$s uDuzo}2YK?_P'Da4i{GCfnLdVa%	Fi#lVP""$z;HyglQDveHe'Bu}>piWXI%	$\$w*orx:79j8gZJd$
hcZ\HSlr(do?&#vV9{`v8=Bf^2(;z4&0eAAL;z8/|?7fXdT>/e.maGuP&-{B	r->Da]K`(weFPW;jt3/xy!BJWj9 GzP6|e;C(i#H?O*/*nL/3P0Laa(XP^x=48")29bkE**Z^U<yBSdwj D8%Q[ 6YTS}N\;tqN~S=(1YU}0Jb]7'*	@EiXX|:nY uIo2,-knxFgYy])``4#YZU}/@cI|,|=P?~<C	gs*Ao4IOgN'"7k`d#s94_&!Z3L\\c+=r*S*!BWXb)Ky&tD_I`=zBCMB[`[rgtIo752jw'H!Z,EM++FRCBa4%=<)Jyu}qUueDcIy$B0&(iD:zvn"x669_WdjkT`IeiREGdWz!)HYyf[wL@]U0lO^b/uV$Gg)+j8|H*fKBkd#|zg[ZLPBcnewMKPSBIUK
'1P12~;?.D.oE_	veqd6c;\gRR`]w&Q9{AW{
IvSV?+^=.v&z$H$F'$})XQ}Gj@_v,][,u
#_b}L:lspQpNkSEtC6R0B+.Bm!4%assB([M08m=!|i_idi5F Z~_#5c^<BL{3p)JwF)QjT;`W~y"E_N,U@|D[Kj5O!%2<9<[fb<AP?*ip8r/S%8hN_VN-Q{G!vUW6jQ	TGG-o28S^@IBArzyaoPwV'Z9Z:q/Q)act9N#fBxT2.NO L{18M@;!TmAB(E.'@!w1'e!R1NevlikY\2'r<4r3J*>q@6DTERpx&DA>r=W@:Z	1|O+O7wwF/{Fobt*5{	 0Pho^d8"EXyShjI:XD&"+p?PiY8;0?7Uns=lP?B:+wy	9aT2Dk[\h85\t70<B])*yR/;p
W9a&%f*	K!g2YnIG"bcl%~`[NBV0B)< /pV!LP0.5/Ew0LwE[*1odbcBV5X6b!J4nb1<x+pC:y:LX13
,`}nd[~>z`z6!nUW?Ku/K%q#*uSJL:NE2|pWK"&{N(J@f4p)NB7i|d6bnYcyE]=E0pshXWN~y<20}+~QN92uF3jf8GGW>hbVV9w)k$zE9k*!
Sbi$WhyKiOm5Mb-SSt\vKtFF[}qql
;rL!Iu?oXr&g,UQD~j4&}e63
x9l}G%97\R2b@3S4.<dPsm>29lE&JCl%.9A_/d~}/p|a)LdU\ifQJn*:@qEK'*Rp"ACwV3?HF~TMEYpyWd#X67j+H3PeE{3V8W;Ya&b&3tE(\_0_Uh+L%<Qc$IqO)	X2bHp;F_zjy3;tiP|0c)wF0h)8-79soM>#TUFS[+m[`8.DIjX2:^9Z[aCg';|L-%"!syN$`Qn}x&9\|JbtZBT!j$Y=.
N3{AJF|C2Ws?1|Yp4qU4:Vz%{6	TK&3:;?r%JT"|eYfT=|aY *
xt-_zm}2J2+~gev8#g{l<*t!:Zt=;uHn??~b`w_{Ik!}m
:g`ker	z5VLX`J!n[Fv3iI-d.sASMi	~^\F"PgsXx',`{^t$Fq)#lzq/qVMxK#Y#	;.NUI-5o.t7d+#Z
58r@d]+U.vZ|*jM=b2uYRg[rH;UtwnJh3w[gvl4?[jA OA`Cos3i=K(<1!*	d3LVqiP~:Vv1<FJ1KQ:{*?(6t%c	iV:5$>gNZF{yj~\+=,]zEJ" l.w)Xb$CLd-C\\YlkkCn+Yo~4dX#ExIU(b!pqVO>hqBGm>@A$Ag#X#V<B<[VfD_?>-of)n*G0t#uQKYE@s*9vpMsW}zUh)'iuJ[|:sTXp?9ByOe5u[eE>z7=sa*gY5kA{;I'O[_|>Z[=n)e8$_8W5WR|FU7K\(;K/</R&"Eb=@&\U:<
0Z'cL)\09ZPx2&	eV!SQ\Z	-N*<=P.z0 AOdsnR3xY`:.;W%3W[cMes{Q6<0!Ma&fm+4'~qz+b2I8hKYd;}X8kzMhu3
5eAB-vY[$wC>)6v#g
|^T`k56~vrs#-cLDfF8)?^QWQVJ:?Q

N3&'Gg)wdBrfZ.)=k|1ge0KYAh3]Ev(Cj>8V+!	TH!NI3SaTa\2WTomI{PWaF]>9>V-/Z}B6l\PKxs9i{t{QiT00XF]?^F6R40:zq	B'77C62P'&/}Fl-yz#402VXzgJ]|Uv)`HVC%t8B)Gf8!JgE"e[&nV=[ DzSOA]MKnjS%S-Q5*2{TA*/^UhNe2/.A:!O=,_CLCTHi$7cG'ek
9*;:'M<vv
qrk)?X\&Q\}$Xo<Ra96+yQ/ v1+<"m4`Bos"'ubiK{=#euCF;6vzW!Jq{:J/,Qt"=j[tlDayu%3j9EWE_AIVSgo`u:"7)hwow-^.A.xkq:*;	.{!dQ'/&6,+CM/>pw}7Px]	|Qq3((	M#gyR qG?^
'h$Yf?B|]y4$B{T]IHnU=8tR'(m>gen+`N5mg"4~7aaLm6e*`Wk(Nv5T]H}704~fzmlisd$	lM<e_*c7g5e/ej4YnjU=N8R"QI]BH76Uw.4yEfpQzD\,J8-<rH(!3c;`5jV0tsPh\xlx0_)P3]3T;^7 ;7L+;7L6-n]bPy|~>5!gb;_y~HL2d#n{bfd>R-a0,Z7=;	@`.K_91du9BeJLw+Ynu[bd3"fl:|cLj70}6%Sw,&4.L`>.Fq82ih3Gzp.[zy!K#Au|r8mb{7I_(V7%5/0T	R?]qID]t2wqB1+UkSC2otw@e6h>S<BoQbpf%wbwF7WyOX-P_D@sM'(7,%L{|T!6LS@a&^@|K4odT) 8Tfz=zKob	/r\OUK6rlNTF0O6	CT,B{REF8T{0?OUW+j4d?GW*dO<5A~@PxU\}0n%O;X:l(.5bl_T<GU?2RS{~XK0e2(A3'[*!< !][@A;BFy#ov2X++Zsi6gfJ-T/]F8rG<H^5sQ0U_w6|fN<[XlvR)0T~8?MZegrJk?G5H!,|hwwh@i'Yjp8ug'E3,5I;JT>e[
4PGH}zH"!CZIZF?j@kd+_hKup]{"TKkas{!C""Dv*;eSrFS-}I;D,Ammdv]f&*OV Xiq
c,,ZCo0i~a[|\pN8(BU2x_`JxEPlKd?2[26<;K}'9!Z(RbiRq81AB?C6XRT2qC31
N|[rZY;u%Z>I$lt(FYaT"l7coF4?!7APz@785dR$ieaL1]2">b`= $Eb,,84dP\aA?di'w 4dzAnsfAPV[}!xrbwD~HRDH\f-"fET|gbJR8[9]igw@S&QNk1UYU%ICw.9`,FP;K
k.5k!}$Q<=mmr_%dhvSpkoA9`XTvEJ[MDFI^Wl#|Su1NjL!f<G<|N<4fyjh"bho,A.YohQ_/QL{_yA.0[`&Qi;	oL+FO 9mX	#J8A^&Nl?5=P7\yHMi|36	qSWHUT,bcvo4,'fG[tF) cHxM)Czbvc@G5_5s-48Tb[hSZ'GF5I4W VMtZsF]}:7W4uTq)t#0_*pA':+\vSJt u<<pw6-\z"^w31IvDQ\mB}o$l_G+V[BkCtA13a8#j0dUlG#f+
$Hi)~GV]Ja
]VA\4QK)1HAz9,hiW<P&PX]v![%I~ w_f|^)G	,I@]p	iKeH~@UtQ
Y/"r;-<JjMV6W8o?3Tv0cqZP,"]knF<u~1i!)cUS6x"{9T/=a1rs[3B>P
=ZqofU!qwF9IzG[T=W%MU>sYkWYOk!we1\H.`>ibNUdP3jAlT$QS'901ZcZpTS6Dd8~@B#&C:rq_^;?b`V\^>s[\2+e]\0o!%N(.O`nM
fkCo	[HCpy3^&UB+_`|-	{8x=!eC_#7{~F
tD	WS#C)>d?spV.^+dHg	:&>lgr.z]&B"v)jb"Zd%_=|u*L160uo|~oE"_sMXNuK/]"TW1QuzlT!+Jt-CSf$Gq|"tCc4c_((4NrE5hBvgdo-^wU,*C_#)N3Qa}u8|MNEhAO0c6wyM+]X	i7%=V=GR[#dX~9+,{N/epE a#:o(f!jQ'nQj^)m]R9	'K}}/kpb#|:[t=X\`8^ i~xg}"9a+vDf~/GHt'0-E\SYq.|yf2-J
fg8`c=*bC-9`I[Bn)w$X+xdj=1dIcoV1[VO{hlZQI9"i 
B25s<V"{!<1Of
VR:l<3H_uuVXDX{J@``541Z9R(N1xfN\n+P0'*lK4C;wT.>y.aAtsD8!Kv$f`D#c^fHu,1
>qp!|J~VX1W	Rb{t}+57nf'x)p<S"i]50O/;d(q@Yx5Ve3t.*lfw0M`WsL*L.#]Y$W%"Y?1LE}+B.T0YLgR\{%#:BUCCtra$.T~23z]|)ZrF,Z2^~ycwCa2_'nW;h$v'6y;xVa[c{ADv4g)opTP%=Et)`Oy>OJ:Il-Slhq8H)a\Q^v_c{$J1X?U6&udi(pr.Y~iXB(PP9?tGc dd4#\_f+,!B=a*pAL2{%F6XkvC/v;Wb]&z~*]dyVB&A.gF|YIRhetqQk'BRVGQ	irr:V@|h]4"{-r	Nwy,{m63\[=(&@anXR*	(.m8DJd1>;Gh*?BhzG=v%+5'cQw	=8V"2CINJVb)t`RIt!g4%Y|d~/-*Enx[RY,@mP/I55lgE	vr`!->$9=z	-Y&E@GHSQTob"S-}0Kq]I5Mpg<yCa#toWDxU! Z"0u/=W]N.}?JJd*:%|z].&!u+1})shTy"+	_%?[	8*3f4UF{jC>%cu>2XCA6+b_{]!};TZP2<x/o4[I#Ir8w7[EW3yI(;^{CR<sasL?k=q;Z)kU[.eaWOe9X~fOk*!m%wkn4";Q4[`]M:"pd!#s"(cs]yL{Xj;zr&epFxvie<;^f7~3EIK}A5Wf`IT^Ss Ehxn$lmyoAN;|NoArvh TuV;En~>zJN|.mEaCM61<4e{(eL}^#fBzB?g[_A/SF-_[
qC,w;*82\eFycL]DL'In{d\l0x9dP&D$aoFm3Y&}5T6|hgO62nC(80VCaF4#-%R9WA"]RQP<!2g]gI SE5_C!26>1}9~"<)&AEZ!Bmg%u'+#stj}\Dsb^(!8f}Z[I5fM8"a$B6_*z"VzA@<U_T@wL3EB*(/z~bzPx=N?G_@I873%d=Q7
8FRN|H[	]:2^'mD&!8FZp[N`"'i:t1	^|["wsi#"1Uy>eh|$Gk{\xxn$DoQ(Py^-`dWrT}<rq/it?i[X2+o;NaT,&p|$Z'Ru|$]`$Zj^@ #Gzb#YvX.[L'8LB]c;\!bLx;zB??9P!K$~KSTX$9/S$zWo:J5`\t|"Y+1 U}>^#Tba|/cy94d[JLw.k9	y6
/YTW6!H`D''=[j%~#pzx%g4MEaZ"U:\T\'p5C$?`R`^!h	r`6)kj.E,(@M5k$v"huZJr@U 'F5XMwK45!SGF<LuzL8#Q5`	-*PZK:k`wLjxL<~ \S?1G`:wexRO\"9?h>H~|x71%.3/]Q=}I
zfj}}_rar:W`l^6*Bq0	Vtr%bm\,*j2JD*vP(+bM7kh}.VB1k-tFnB1".4hY0OQif&}@
Wlwcu5k$E	BA)[AK+IT>S]NsEqHi_F
O5%K!7UDtW,Sl?cje,1Q}! S;9\E2Ck_14PEa,;%rtq|"t=0w 2T 3N&/Mp<;G?F/7Tj-g{[)3QS9Jo"6&tV]%kmOl';IAKL!Og`::IA9GPm%uD%mBR<\,>nKC8t7dRE/SO+v@F7Ge&Dm*~K%faL_&P+REQGC8`U<zWvkTPO"Y~`.U=y=F3sejMa;$vYr	"!$@ bi'Jh<~`/;U#(F#|k	F^Y0bq
OZFX@qfpV+\Q!Fzo|I0t[bzis*!"Qg_FiqQu$.CG`<-+{HAFGU
2DK9wE*f9S/FIB:&BP|+#e_bt[*z1^ZzT_OARLsvZvS]SQIkncqQUd`X>h!y84(QMb=A^Yf,zo&)\0v}"s+ZUY:n6I|\%Hp+.h,C
-L#	Z5Cn`
xf+_$mpX{NM+iAg0@~*$!2Mdr:;tf9pF02sgn	c3\`1DJek%*C#4xKd-o&J'&?$.u5;lEubO.#^#P8_Tff{qH_4%:.([]N@m%9mvdPVH[Fk4y+vrh8}^5lJ5b/rQPhwEesNUDf`a,d&HLA#oo6.8RWV}~	ey[#dT{$TRFq%0!6`F#o=}H.;VtfOv'xOz
PJCI"JCK	mmjSo7gKA$,Dwv1q4U_33m;JUXgeTC)tUi5TJhAK;+\AEPuzG.')iuHRoK&^EDp*\&+@$N>3pr+	#:^\gP)ZWy_&hNE],	hS'_/eD@84'1fLvBkB=q][KEA?9_2U-$QdEvHwK -T`=)iWm(4Dm0bN3l^:uwI,Td)sWb!, ^FKvF14,<)<Xm$CA_|2&]s(!(|g,FOy3mxDv4	?	p6&Id(<4Y-%+(Hb0FcWFnkcC;GQNM4huyYt't?/_Z[9Z{E[`= 6lt8I4:+L]5RA_f0+#-z2&xRb9M=cB^%I7qsRJ9+{%#!UI.Ei?.i
cry+}}Xq@s@7Ba`.hG{fMA0]F*Wy%b78*?vV2fhcv+IK4vz?.8}"||l?T:yz;$L%nk7%j};s.w.rEj]+ipK8W.HZP0\
yWbvz7)'.}gQ-_s,w}EY)bD9MGDTwx#y,j}^*butj,$/fm``9NKU;xi.n1Bc0E3p:UT>JF:%j#tImsAe=b<SFMw/SH3;,?C	1B}[I;-hsba)"1z+Xu5W-H|Jd8yy8`'o2,5g/AehrpTD{XZy#e(I8}qUob6Hw=n>|WSdtE-L%l3T30bTy-W/S"G?k_H./CZ)4~N?-/[KD 0t3-6jLD+$riY 4}RZOG4wYB*f?2|rn/?$.j{7!Ru\!>QL<nH#hq1xPq9F>5?~~2m/~YI{JVKx}p+g(n,,wp'#`PoJRG%J`	
4lT6B	"/6GXat-8Sq:SV6PsEpy-bE7+H>Ovh@.{7_cj,a$K@D*K^a6aqRvuTNsmdTqdk2wo".8?&C5|>c6k!,%15@GDpR>1Z=?{_A;2
UGdU>g:t"7Y{fp}Mrg1=wx;/UUbpDdDm'>4	 TD)._Qy2wmcQ=\.Bi|U:rh'j#J	Jjx=ukI=Yx7uDX/PziN)&#
7!.,POEqN
.>w6MOhQ0V19jZ9R*RpZmj1A`V<_tqAM}Qg{O)
1Z0rD3cdXmQ`0YeK%:6dMM-$%(BFoZ[)Y0g:?2gcn}O+k?Jo>Tw\mX	7P30fb**v&,|8kbB>X[szY
P[T5(9_Vn>Fmvzdx'ge=Er/94hm.|-x|VAH|p&I=[x$+&0X__FrgHQGa[BfIOazTJDg8$0A&ZmhW^N}TQ9CPCWbq`5iV?5i2NWFXM^ArGM?QDi{
z&Y!0o<dBP;>Gp_!2"{C&*t6{$P;je]Q=p	V$J3lO~<2[P[yxxbkg%	$>3
$Ql4QLt)%K,1IWW+gOdkEqKK}
%L]}@]QH*NCPs%Dqr"mO5[4D,me0rT.fkyVaBRzY!xE[f.kb@t@(X^Wtv
VH%-'47`hlPqM:3C]k|9w#X\gigkBw3@'OB$O`GA&U>>48 B;W!8FTn4^aPe.V97-Y+I91a'UpH'I3oEg=aJDQ=9PTa.8\C#c*^.Lw*wG$Q[Iw{eAi6:^_5C?x$j~:%>wE!oM7?(Q1rI7P$ WqxY.j~0NZKtpNpC+v!~>Fxhi|@,Q
U
[V/6ixA `Z[f5"8DwCBm QY8=|x5C|XHL
A u5Y*$]P:IH1{0z_bwJQKP3fWim+PMD8i	/{7]6MOWdH_w6)	#[Fqa\=-V{dJ'C@Wn3%9})xe%5uGbiZ?z<RZ	?lKw/`ugH|qs5,jhJ30_+2Fv"P{:}w'%E%("K_.X8+8Ft	.G[
@blw4}!S8~[46{;oqxpU7HC(r4<UyGyCWn[B_cxyNK\Dh\$>6W!k1!X{+<u-:;dp\au )[iB|?mJ`ho/fycJ'?s!6w\jgT=KKq|&HS+)t1uWReCx+[ <{{d
z+t&XSD)?AF>,y]c
zTx{m@~@Lp%_]dT1vp]Q~uC8xK.O5yv!0Hq6ud4EQ9Wf"@zjN}z$&#	,;n&T@^ByEI8\L(?G=n?t*o%.>Las@NHJVpL%fSliv-9"i '[n4D;QM!	,.-Q~o1[A,Y6jUe7,{0<nWX%oG)T;Wp|h^F5AtZ-YwUoO
x>ZTLQ?H:{.iS7Wa`;$`(B_So_N"q8a4NIu|z&&Rcxp`j5J0[#`t)b~LCNTQG	`?va&$3\/+g,|7LKB*bL([#,3?Y%lh1sJYp'o>fZ=o+p1vB\'*fYJ?CZX@.h?v?lQ<<d9e7p-)gDR_(r/+5 iz #/bGCW5}%{1iG%*hAb%3)iTGa2x+.St'o:2~+)r]j!6Z@_ps>:RuTKQ*})ul+X&hbS	H#un`=R~!
H]jvd1tZ?jV
bs+s
/eV`,x^Cc3=Vd]5RkZ W%YE>A{J?@X:5wYGx2
 *(XQW(Kx2'z9z\MWA=hL4(z<{mt!5%		Wg})GS|{^YrD?
koCR2!kx'Pw9zl'7wJGkN3
!t.ZtP08iuR/l8Hd`c{x2^!5oO<g58	<kha91xi=]H`9/iab:&'m7Hn C{hMZzfhqJvo|B{QYXh}Iz= gF$_bu.`h6P#s^gBqN/
e*ZV.-|06I5g{gr<pC|Xut^].mq>"!(g.iS%CF/ ;:euiNQxeEu%"b% {-TpG3\ ;~RM3k}
T#Ibb$\|4qnW%aoYdJKL!Bv_/tHA,\+d#IRK"%W)V+l\qq
	AEc!0`N-c-A[.Z]a$nWQ;-frDaIZ-\\|FskFRRI;}/2_OQZ<V:C&,(k-%'B}MaiS[`!o/ 
PxhOsBdo$&w'\[RR0=O_Nk3:pOt)#D](pv]c
7}}|(R`HXy*@$Y^&M8Y<7$;~Ti6<to>ujX:
k}9[ ZQe/kDQxlt@OI)8?6.c<54+Aw-,F'Sd(pfB'X],\SS{
9t.R+4JBB$R8Se,kX-.>llSk:e@OyE(xM|E;qS"p\pgn`s2&hwN'9Z5oO8')UkYt2/P,@)&8Y^9Pb6/W%:qC?PcCT91`%$,"m-em>7fBx|6ujH~J:cl,2(LDH.ba!t6$X0>SU:5\Mc.zBj/Ha&'Om.wz0{:w]2Kk9zND|t)U `1Sa]d%ibJ9e#|qB0	YLqa-L`Re4NC1-1bq'VBCb{tmZ[bl,#ro=D+.3L}<!7,LG]h~|9yr0@'1PSwz)O#2?	l0zib!7l9]zJY(:*X-6.=eRe8Io,}>EFHFytaUP^)h;612"wM[S{l3-6Q:$4({*b|o8,QbPUwTVU.}Q1#gOXxZ!O!]^s}Dk84x3D[8Y'2S$WG~lD	:8B	6t:O0efW	N"ezOye/#	bdL!DBnMF_;Bm<c\<y?
Z8DJPo q\DW$.X+2:;\f_9%}7sBC
qbPsa<_1ABWxSr.KK};+cmk8j.?`qB7q9j>sWdAe3O5M	)=U8#F5V`(50-Z,QZ]I 
Ts8.k!+LG1@l+Uuh'(^^gEt:{Fa])_)w$||TTbzY(3T(-W>PL7
B7xW/Y<f=B(17969N,*.W?*m &$JV64<TQ5xT|:>|MlRt^Jr3F=Dw\J:f@V6;%H99gs)w<n'U@j3+nS,%IWGY"Q`	*T/\ZQA/Md,ZXZ=16.@xnM8"BV+cR:u>Vuc~\jg":+:WL6^f=*j,	?fH1/e|!ysNH}X1%imw*`5JlJM$++C9T%lh9@Lj?jA*|m%QIyK|MR-Z,\
KqNtQ$ueIHb}6} uFeBwC{w0B^)}81`#T}xE5IbS~b@H<=n4IGrHLkbB"Ai>>YvO;V~56wsZM`ab29_x+SNK)"ccyCi>ZyCF5?U'S8-J)&0U"hDKwO`MQG$cX[>r*abEj$q`)V'{w{+r*`&"VW0jPhr"!T6Tc:C>%q/f`zaA@yXz9RC`r4WM7)>Do}f\G((T-A>{0w-Xzv(h*BP8/Exeyh'S?a=%];r`{f&~I_.y~vl}AI)5p$wzJm_VJBlBb17l%Z"|Kpvt2^{)=vp7oB	]2Ae7P&:(P$40aIS5McN>%~DHUeNz?{Z|6?;\Q<Gg~l,
EVjw/3|{{(4G5F ot5xn~p`v	lCk<G.+Cc&VG\/{DFX_F
RRhx#FJK\=/dhF;G,eT1M5J,j^a>ImF6hND"B+kk]Hv7nNu0Tv]"J1EGqI8y:hc<Q(Zvdrc_(7'_/R7RKf_JDUDE=Q5d1.x4FArJWq0)a	;@yV`#&9 t#N7Y`oq:JO	XKmA
*{6}FNTyKgM'OcI+u_Ko'WjUXbG6RW0~	5l!)h'5TVu1lblMduxu=-A?(4%Afz1=zw="5XJLM~N:0:G{cu]WBP.J5>`"IVFlW.b9hZKws4%6ss@W7tjT|9XDHqe7Nl;8<7Q86iB(YW^#^4a=\s}1Uw"?\D!i-z=v9v%"M@mO
[$8wpuwCeQ>FA6@:Ak5Q;
Z+(k?D?Wt|,tFI)H]_sp& f5UBP*M9=Mr5]gPwG8ecw#fn'~R(c8tD0Y\2GV^J6+o+*T40xnbb"w29A%Co:f_)"Y?QYkAG_G
@YSxC>`F\>!C4pA*\)cx_cYD,SYJIKvY0oKI*az]?U)_7fV3j^A[Cu6na*WFC|b5<#8<NQkjz	W{(w1=wj=fs4@ C^<k?!
f*`75e_'6/@(13c+_OM_7kyAw)e4]1
Ef#z&C]:WdDOtX01@PMU
 N! P]
)c*]~H~Rs%&6vNw@GNyk0g(F\/]&i`B$UFg2FgK;`9Oz@]?nw1?k|sPyUqMJbZmm,j_/R@/tIla#w1|qud+Z%++|	.FLLYL+'oF{0<V)W5_5xTR83vIV|
8K],[7r,9BL]1ij`,'*h.#	O-7bYLC&k/M*.rJya[NmxDcW[se*C8vM%o_I#$Z.lfv;{`"QT<w[I9CM3H7SA3z|y9<U&D%H8_7Y`/>%b)An*$_la(-2Sd|EsXE$=$o5KGjV@x!zKgC+5UisxhqvWZFgvkX;u	1?A\@NuNa 3ILNb{Cgu.[|qu4/`oS,*6{5WRV`TZ$Z*	b>&@%fQ.]n"0;=QU[Lb040b
c2_Cf^LR7r__K,|][iri1uV"SRj84`tge4h`Nllrn}'G>,7{*#?e|)^Qx})
f-B#	\_j{uP='9VTUck&y{}0IM{h*8d
aNJgsl`!+D>'bun?{cm#RCHt5|=JaTIlBSD5shl{JL6}F5xu='F/K$4kd$eyy)jk,`cmC|=x>\VV^Zv1&{-Uq\b9jx$i4I=&0g_ihiCb*yL;Q#,?`UO,$<fs0.&6im#|kYc4I.E$^x@`wE*=kah	2Ein<bh-)6$]X(:U]J[QUn1(<h'Zhd_AgH_[!	3ygz.ef<.l>DR[1dRmyGhW=43(k`1^p+s7(N^_>(%tGE=+?%Q3WP/xS"'rg}-*;8,#]w]57C)B{7jleQvY&
F:6Y6y#mz{uUNHz)eG_i_7at]a+rS'<\=s:i:0'q@qC$g3,!t<6M5<J:wqQA\TE5tFUh|p Zr4%[vG6z,m,"a|mU[VQ[""ia95HUMPq$Z:"&eNonh>hUvkEcgN1&VCgihN)m-
/1_";v~5^udpYCNJLnpLi%ZIN"j7"=bVF)WESM%uXnSatXt=%-fyKM1iH[X
xLk5'(f
45!EYdp]%bF:?V7ToYiGZ7
oxTGd1^21I6c<A/GHVg,c0">t5m8g<n}_m:t)PY8	&ztiBv+HVD-UjK(AN3AiS/=})+1H
(L)z>]D'fO!Lu|I/Wic:8_iL<N()xR,y%W6Xw4<2YQG^(441#tNS}	T%SZdM?K~O V!Hpm\bBp$zqx?y16ybG|iGl.a)AC$dCcw%J?U'm.,|Z[VYh]FyKq9S]Z_.,0mK,mG-kd9OF'\7a}V=Ro2L>\mUTAE}?aW9yU3Y{5GBQuReIui>j0#6}gC<}Eok<LwW1O+rHGhrxg%$kE#D-M?.9h9PfX{~9/y4&^Sq4o="iKwH9.nX+uUTNsm@H&/tN}?'pu$qpxCq$(Mjjs]zcSMp|U+8B/bf5uW!Lp"A@\GD=T,=H-G	V\OW	nx93<A i{lf"+ .<PB*P|?;4fB\'r!Cl33oxCs(*B`cAR@_fzKlVM5,n^mS(,6_rPP!k#+Ask:.(}b;E2IJIq
Z Y<t!pd;iNEkU5L+`7O5>mP`.F]9xV`:u|f@*YQ9TB8Y0I)=DP?f&Y6lJ)0lp[{uG?)@"zkAq6ot2QZ0P1lM!(g8tffa:u>9RS*z}]!s)1!agAAiXXXW=}
+`Q-:mMi8uRGiqZAgY]e8d$@7J*[qZPwM^`-s|a^9g]X$/$1mYO.$Ih<P8R4|5z ;\Ly@Uu3=T	[9#'o9R|n'Feqg8\$zqjzd94n_$7BCclB:>LYKtLD+g
>M^Y;GTu`y\]#'-ONxaDHefRb>EmKTT'*[@EUZF}L7k{$A5K}[[jA'VrL\m"PJVA2#|xVVS@YcQS}<"\Tx4foZ<\^ .
sx?Z$W(#` H PN0BTg-calhQaD;Ea,<DHLN=LQU9[q'bF7>d&Euzf+K///vSR03~N9[9Qj-z./L36E}K9$(%jX\7AVDq]jn/,WXW*8&|ca1XjCfdX^j6iEj\c??=H@RJdrB o1U(Y8EH*@*9N$T0f*LB'.Au"#70tmX'xlnZQo?vrF),*}"KE#j?uk${?sU5SZK'3QwuzFW.!(cdQqR#2ge#Kf!Jva<g.OOj)~KvH/w}Q:8+BxCPqP;JI'*
+kk9bUzJbgwMhk(Gi"RZaw`sJIX$<|4lv/Dg\
;pHkefI8)Pj
K[:>{ n(MfH	CyRd|?d|T%a\Q{[HGj,U.0{&=_+&U<B?x|l!0
"p<E-sL3#Fc_&t^W rv[)_RjyCcqh6U=d#Auc]pBD9/+:u,Y&?|d^Bg}K^Z[n}<*_4,'_G9|TctQPVN;vMv0`4(7,uL	(}@un5u%|GRozBFiSIQ&VmgT(aC+A[,\&imYx=/N!lR_t`L^!(STH-;$!aiLBa'Q@\+e}{{(;|2P%\04
3db8p){g$A8	%, W/P!Qf
XFSp$QiY}2qq^Y
9uMR-l{5=O,F1LP\G]7a`Nac
pXLKK5X|;O) Y"-VNBo3z ogkb.RYN[vjzA-	A%!8Y0xiy|BzTYOpo,t{!<X2,'ioZ=+xtY\|Z7T!2_L{|{8*5Q
+AU-$i,cR{*]"sz"T;sYMN5gXx2(QPSQZiw\V_?y8$@FvxzOg=9HM\e|mvl>tbTAQdEaISU?{4:cT1SF]]dI6nD|wYhli`mb'G2%+uOc5&sH'h5,
yyL>l3fQ-;?1(9#p/Oahw_iHV"3bGQk%u0%cvy#O;AXgB7'#eL7-Q2u*.jxApfYSxVJzz&|AZx\ %?6 {AjtLu
TsCd6[[|?Y`o8cPv:%)e]"J~VXQq`z%s_;2{Q'wT6O @c<*teb7ljK-/*QP{Tt(ZVE%/CWkm6PT;vRte#AO]Xx|$U\Z@.c|$f04p86iVA}+\^q+(='(hpw:D?{0"dSg%J/"Z{#.u1I@:iaUozC:>WQfwsAD6b~f?XGZ
8\Ex{ni#
%6q?Ay7d+]uoX8??&09jL9*QaVpqG/2,/g)djOO/-fN9rEth3 	H{$Y+(]ANU$~prisF{|]ojYViKXw2}{eXe}UP.3?n_%#s_K<Xfw?I%/qx"sNChn6qIwMF9',!m[7"mL>asabM<=8.:7h>]r86b,`0MS\u&2ydI\ is([8HB
c4Ey_.p>Bkb}+.9$;A^k.!Io0=PI#+bV^thc]cc	z6Z?
AgQDC^imFdlX,=j?3)rg/0ZWrn)K8lMG:|zKpZe|V^^mDsoJmtgOT!5`L/a^GvpgCKz*S4Z"p6aT3jfk6ul{OmFOiK&KmdU0P>:
5xwxE`3[RU`,}M4,[&[ld Wu4yngu@PS^3CejEmo,h447S;50zC/0:|gN!2't@4?Wr^<Y[\Y0n1lFMkZS-X;Tc]dtc]Uk'?y;417%+hc~{G>3o%r @4?YXjrB$sW@yXiPT4fxW"-o$/%LqtzoA(458Ja~|l+Rp2H6?''XQ1 .~!V8?H#8n&}bW>v%/&=%8Tx?(hah1RtH,VQH/dsy;m]Er$VkZ?(buiA:c\4wmg@-HEs>cu$+8DBx blH,x,zB$&63	MvK(pb}z?ksJGqnO78S:@6mfy_LNho8ns!	&.5<d`gk>tG34l3p[i!X2>%WRG1A-iUP=)daT,&CO	'2I~6[A&J_KA)mXBt8[8X]Ao7^4q~FLxc?y*I\b|dlHNbz'jEg:y5P7E*jeG+y.z3b*	!36uX>5a:_W:Bck{dy=IVq8&@qU{,=dKM65ZZ<}D}I]hE2*fbf2dZ4m9oM0G/yQ$}#	*6m<!%eA)c6~2B;VU=Te"Eq]["]-#L}<XGW50/;:nAd~Y.\BZQ:qJv>Zd7ZZmnMkxmt1!HhZIzm[y
^_U0DFCzz,q{x?d	7"*AdfbpZ;dw8acqn#Dg|c/bZN?5/#4[\-;M6{6i~ZzB;}/I=,m2.
$XG'9=V
=jH~K-\ASY'MFUI~#{EOTKQo!gY(uMW#DH;P\IC: 3eL"qt'Rz8]kO+.)?;/{}PJ\wv9Gg&:y63$6@W\a!LN"hw*OCqlQy)'-}G=~lKIB*#kvJNiQ\aE5puwKjIU:z<;+@z3%c0-[[ri=>\t6	`Ty8}}iBT[?1qf#lO_yj[/sa\DSI4+2S"OXPGHX%&0hpb' /l=a5xz:?F&"*EC4@p\2L
9Fy~-B$Z0pDQ+XzkSP1;,Ok!Lu=A|&3FGIMj{	#pYj^dEl0Be	h@$rRz,g"d!Y9u&)&fNwfv=ph_ ];;Qjq|j.hl&_iC]?9sc17!)r-IaFItvnF@udFARk3e85{zV_IGPcW^qZbP5{%&D{MiR0:>}4IFEs1w^, X{`'Qko$IyPp9P_OH
4qw~HNlX^)ckG`}^3Xy(\#G
%e-.)PYft|JA-w0csg}2Z"	C<W".hO|-Em6wa^ ESIG7)}rfSj*?5DR(apqfH;wsm?e*B`':c#y4q`:^LDV'xZ^X)T'fVm`Sl{A7-krK(VJ&l]`qF~A 4a!cIN@*@E] &L.;tWN=WU$sRl%tb1D<2@g8C=dgvC"VWXV_vR#0SC1:S	9byXnB|~&JN'oYwR@6Y~|8N6[{Vc~ferPm+c.@6mfh{@G2U29AYd@:Hpg3J&m>rLWr*k$vzi?Coz2#-V;N&eIs\onno$s\b]x0v%i.C=|wVxvD{{(K0ZC]x.|H@l5iGDJY!]/gpeKiv^h||EZ^g~[1\2PPN2=LXR*K$$l*0T/eO[te>OQUS|fep>$$o^lY9{o!&Nt}+>vI&*@]Mn R\W)Wh?6Binm'$ 7?Rf.i;tIW.J

3pGO<^qiQL:U[JMb8,$HI|r[e@T!tHQbXANbE"&g;M*_FX(Dd*&34_v}%zh5H;@@4C'&dgT*?"+#ByG-gs9-a2[pB)0*mP8TS#}3.6.	sij*|BREm;9{xMG
0l<pXDD}V4AhTQ"%s%m@UjLb3_LG8Rg-LYC}|)q\m4
!=+6A
u?n_I'{vAloc6TALb?LHEb2jpce<)@GX	S\t}uO6myD2g)_N!FzM-
aNCScRV)B>|y0STdsB881M[(5vR!q!2DK'-$*0|T^y9P3'1f}=LKQSW}O5Va'7..N*nG8:_ug*	".<(d_^HHa\p?T*z3!@K>Mvs7Gi=VrCma6xyXd!P(E{KfD6BP@fz?QyH}ezi}=JAl%[W8O?M5mt!Pmh42^vpsW1T	gjEN~uQly_fEf:wy6eP00?]!(.jMiHLCo||ka0M(g}5BcL]YJo;Mw1W2M,o`[7V^d>\1I6B3YJPZD:GNnXmRpoC5fOozKM0wkbF45U9lj!-kKv]onhs=X[q
zkt7IC:&
C;EPt;~0By<B.,_LZbp
d><jD,+?yAeAM)EIhwkpFH<rIz9ne)Q_Gw[g+U7sxGy;A!f2\0L>C#-Af9zt? "+j~:T7I6QGKQe-?V@7w>#ytYC^U?&jZ}KCWrD<}o,yOo^CP4x\9D^@{t/jS6s
6JB|nu-)
%`#2uNHL]|AN2G9EnL-=V[)\4\xWP@s$+EE\kaeCR\J![uKK~{@j|	/E3rY).=O-B$ohua@\=p)!XCL82aqD!`=m<*gYxK?5z0(aoff@GSi>HnTF,Ak	-Krn>YLq$6".'B,%2TB/m	o5?meFR
6|(>fkOWA22FK-iF1xDQR7S?WD:VwQ:)akr6O4TGJ6h||D^%
rDOL2_x]$GU	{&y|S>S?Cp0{}YLMF?H%h<y:Wsbt<+^fq^D<^XzD#d3:,muo]I+jd?s+EXzO\!fb*G+G5haNsY8v1UrQ&{)k[=_"u'voYp_0$7)g.XxQ!(+"e<0s,uLr#(b-cu@hIPvP7L7[jjHh()k.9~d'?T<Ol93Ns\=gX?DQ-^Ql@j%orLmNhYuKsBu1yplFU*Sg7H4c+%.<.KA"EdlsiS RcX*]|hi4@v8eX2{[+E!xEmqG;
.cy'3[o-{D	adC,|y2W.^7B:-[:Y>[3>aPN=c8@q!#	87S2*bkru[6JQcOxiR-QoqIc*#-06$^~|W.xuWx1v*ri=c&{+lE/Gg(/nA{"AD~nOLE`V-*6!QX7-buWmJ}U>$7|8;8CdD/mYF?8aiS[?E1sS+!0D	Z1?BW_TxN{gG,z5J9|ch">5-m:7;Po*"L=GQJ(RMKulp*Y;:zbJNHPJF;gh]Icu+-o%
-?{_yq{Wj_DqU}ATp$%Z(%y[Mo'^	S;>\(iKIb)Lv?DLyG8vws\z*);HMkR~V683S2HDW|OPl2qK01iNk{0:"{tH4;J<tr!Z-&Zq16F!}6z	_US
}N8@)~~Q,!PNcG9CY0^.A#&":yQRlq51 \=-&G3XY/ a,%h$n8u6=Uc[a|FK+#{KZf[0F HGP"$F7XCU]31^us5BCxN1'WoO1eTZpF%	r]N\mu0ZHXuC"4$j>3Hl+A]d=V7/^TUmvTB4Ru`LI)+GR:>mOr~!ZXtyJF>xJY'l;ERfd/dFPxnv"LG)Y6>x3\<mlp*@MiJdDMLoVL{|-v{j;H
A@3n	0fHi5JH_DSU!Zu~<{u6&(_<YB7gW{`ekHS_$ ;SF4ch^/aT'YJUP<q4tc?zp%<kOhaWr>)&R-?K?{TVqhF)nnB3k6g,/t9..m"iCJ75-doV8Zlg}K,B]eW'#Bk6(vfv_
JC->goJc`6$.q9`9lr{N'Tm8rT94SW#P*HBi	p%}q8PcV4Inv3n7;TjfcikPSALy1hAg(z5]SSvT])z<W&+dDc<@v)0HIoX#t<'8z,h
#U`\`XKo'6j$;8`<Q;pKPRRL)S~]pZ<;'>YzyKr6H4)[;:<'Rbwj3s$"n~?@'WW/ULkO[7,a8=wT+_$G2om#ISTqg|g;2nSH1H[]FZ*538\l*0+ot[_/u3$g2xv>,&fx^L,PxyXhp"$/t3!1!*0l}+sLDLb
><7@uCL@L}XwpP.o_>T4JX<zS3h
U*MAA K)hY"pt&sg5}HU4D<^Cjr_hS]U7Yhf)Jd/a8EZ	Jxo<]!mu9;Ig*dSe9`{3My4pHww262sd4Or\-Yg^%j,?)R5 F%~"^)8~9+^cSlv<{_=~#8HWy?]7bxN
'Mt&RPJ*>kFS'|V=`hUe/3?(s{~,.h9IyA\F:Vc,cP.T
F?Nm@/h2Mb}Q]KECora{KIn>K$z'cve|bX0D\vN^4#x^4@18W>`V1cTY#cFr|C~{/Q3w,bc+aF{6>S3=2L1c0<dSej `GKlM*XfN"VxlJzG|CB^bt$3		-5f\'|dPsd7+?6'\*b#q?2FPwjH:v`CZ#+:g&&xby}LKT]/Zq-e6[o;T='9gzyG7TL#hcWG63ltSf~Z+Y&(TK}x:KuuQ;%0L2;^LS(bE,$bh]u;IU,K-r.5G"1k1+47gD8Af`sCWX'jF|!ulzhak"7\YuGov{3o?)*Uo0qBR~I>AOnq^2 
e_rts _2H<,<#AQyN+8&
kz1a1yb&?2";"q+_hs,o;(4PAI
z"C<l`CB(|0/z@Z9K&@+Yt>ButDVh:<,+|8b.*@	Gr|A4Qd?r<n]kpYQcUKn'$DAvI}`iIYw
"<]a.y=e`]a[:	v[LQ-^"<>"!10\]=loP;%tjuDqKnXuVX8mq+r@C0J7kNV6<)bY3_\pFsL0=!LR>cn+{I!"G6,s9J.}Q`+?aT'm'jX68l"p}=87}!?dM{XWYzLH1RbDS2VGN^x?{{{^5_:i_I8traSwDD^1bY2Fu3iyj 	gGlGZ*^Y9>{XTnS2eUCq]\c@o]X7c{rr"JW#mb'Z@NNPC2GP:=(iH#O6,(Xfo6bJC<+j8HT<QO!hjEP&~:&G$e(;NCpOm;9&<j|od Pnn8AFp0#rZsBT{,k@8Xza_#?02U4uib>^cU@>[!6z\MZn]UbeBT+%fX:9vl\(ngWIJ!"aE@GMokXkhK&f!p@,9/nM	(.@c92I*73zU Ce/CB3%
Rhg;-Eeq$?\zqkx[?WB)rH`w{<w}+[
hl!s<K;Cm=Prh	OU2i[_\`gdHM>,xe/b02CtDGj_NTD[(CHAL7^*:KAo5C#$;/c>Oa ;?hsah=cWp7!"Tt}XW<M[QhSvX_$C_t;paBCZM;J2#hJiBehq*'ZG+?#r2,-` d)KP=[Is"sL4@.%X<RaQ]t7tu][=JYE a1w+WS]JNW$HABPK`-=DB[F Vb]AcBwi2X3BQH7xQ@mL,{Ql^rN6shjfY.<k8V'1mG27a#]T	?Vp&eFj|JL#&.WK1WO A)h*AIu%[@jtz)eEC3Pf_$~Hza8*S>W'lL\18Vs8}B1^X!g	FVDkc^C&cSzB	F28N8>
s,(`|LwWG`;&!w&l4o>
[Is^2RJ,_n.tY]FBS]49HgDbF/KH@0X,[_qjQZH.[*M7t"}mg%i{<gUqa60da)FY|[6l|KyxK:M|fqh4`kA"9Dk"k
;4Mj\Ai`TOU#U@)NFxV8U871-TnQNH^D/RYgXy(+*%FX;?a]u,#$l!G95;lBh~c
gU[[TV34-@Y`
~e_!?n*G2%;]<li(Yt/[^QE[hgH}928m"d&ae*B#kqtEiO&<8rKhXAq$@fL_Velgx~rOz!@Y!^yxpQMNBedVy&?ES[x-dqWB{G')!.hNA'j`y"%;@^5ak"K\2dw}M#<z5)v[|QKB\CQ:`tK+`)'r]>tqh}#'_lxfU6q5Y^%"jI|*}4a]mYrrF+jy>pZ?q9{P	zi\
`5}4}/u|#{/'.x@~r<G4{Fr_O.g~Kr@T2LI)Yj6K]32yS
Wz2'[*/06yoh:S
2x&+m}X3%*AG}Q(z(7J/dY^T@?@~jr3/8+t%r{TMWP"H&1*`1vBnY[Ub(J`"=^VF[n~-.I49_:hX?G[\EcKPT,$DFE9)KY%
r	Eim_@>,;yP0R*p}Q3S96oM?t|-#canTw> lz:OvDor@Pcu8J2qNhP uprx\f/dh+3ldh~Vxo*yb-04R|{Jc8LWQ38X#"4Hm_g!V4']jLSq#cYQ4lKOY#0}99@/.m2cDo&)(}G$IEe/[.yY,*H-cZ3/8]2.UN7C$R:MpNI$s2"|-.eP*7f)z{(wUjaRIZbKa{*V.-sj?H ces^2WEbF:Or?"HYCQ-ylJ	7c'v+xZ;;?Xh)=54BPQ9E/F`D6tj;CtgcC1JJ6U"aj\(e^CU'sw.emS|XLog?@(F&T} i2pVfDp\>*o<!6}MP-t:5jq}A7PD^YlMiT~x@stky)l4+{nWi8SsB#2ai b,g>+F=QQY~WHVv[$A><x2$,9\W/eGp}ErToeo.3L3_vq1	A8d/}5!& ;m{ID~*<Kb Q[M	0Vu8eI(S7:[8MQzpZ"p^>"UM2k-X{<PRt$o`lw!1yo9P
X<2HP[ze+"]X"ji	
,QzbkFP=cz/B[<uFO;IW;>VkXJ 71s31ATsBXfJq\8Z\|{x4if/i8n8{*'h7guyH
p#~f;" mwGTmE;	|+m)@c4	}vS(S%I'_PctI?_0Jy
*C_m~~b{D<u|)y<%ao3yuusA`<vQ]~KA
zfoAq3<"`(m^@0K_;19j{lC)k;y^M
Aydli.fG]Ft(S.,Q+:(7ri0O:wj\>=QLQ7!w(bZ(x_1Ztx6YUF3Bh]a>D2ezO9vW,ldjg9zt(3f;28\3'N[(EP.~q"YeuA1t8H>qE6$D&cM	;O4?3zrBtc3}v^.,lhyoaPx]K<`b^Z2yjDK4/H2;8;"l&5efC&T,g%=i{e>($vDY8*,o%Z4KeP2=LxN<%(z{t?d{w) K|TZXq[MOxxE1s=^Szclk,z=q~l!)gK4WP
QI&>9P~YVsM+FSC$`&}hg(f!TAn7FY<S\i2xNrT)Ulng-c!5/msW6A9ZcT"Z\z&4&@}(_sKMZx,'[5|4;(,{CsL> Vd/GnFA#(vc>R=Xe>CjX3:6MG:U{S9%e|vsd@n:haMrU0We2@_h\2P7F$Oa{oTu288t2$-XPz$O1|tc]R4O\x/9 [rf!^TEQBgB38D],ha![.(++,>[Z+|J}lm]/0+S
CeGkxq5:)1jH<eVPp.Mut#TB,F:wLs$<`0N8-YHB?6<RoCL9^vdGI#>*cFu1fVk)8i}wAe=>(*-D"Rm bsXtc[7U;
q[1\*F$MQ()k' G!$bA 3?w4X8(SlG}/f: }jR70gZ>1IM5w.6~Vh(ad]R*xTft
G?(E1u@3y#wQ*^\mMljjPgr)W`9`~!
F>p!J""Hf[-5]QP7csS$7r']*#4A5 ?|']DQzt2buoXCmXm7QAw&,*2#\~"%v*gZz'xe*UF6>{bI"I8krd:=U^zrOW_*-c2]J:gOg,HTNWna?2%#/hs*;YZp}?ezKWXQCH&(gk}1(-(Z83QE#WyD}Kc#Y|YshW*du5gYT*,c*8{p'e3)}4v6Eb\8nT-zc4!Iu?`EevlEQ?LN^w^L!q[2Tn7+e=I.!yA{
<YGPcq2{gM}YPcV7YN11wB=8S?RJ<RH3,Zq<dUvx$r~l7#yhOro#'gB'70~=LO&;wKC.-A!&OzsZ[u>;>S]u27=0(KM|CY"]e(GQ
~OHxDwvk,nQ;0&EJ]pyu<;7D(gpMLBOV<(0\w;_Ms@\{E*:(gFH)j"W}u3WBYO'{u`~xSe	mx0<%\6V8[5X9$N[m&K9uC6O+l<fJ9+NG [FO:%366rHr3{(iP~`e2)AtmR3j9	Q 'M<1y5h~Vk5h@q[Ckmtg!H&E2*9-='5,fAU1}[6ei0BJ;icrmy`\r+>&2Ro^hxO`rW_hONyOW09h6EuO"&4Km=EW%/`>lHmxGC.|(3*F<oK%0"ODc.k;%<yuRvTU y9&`?"(D"LfS.>	ZC6b3TEtc.b9FQ\-T88Z7:@C?Ao=1f^fPm.l%e:GZ,j;x1) AtgjW2gVEYh8MF_rQ|wqq}	j{GnU2TD0
mrBP_4cv6bYM0ub~2*L,R$$lP	T/_ ;S:vsS	>@hAb##|F9~@Q]eeiGb=Bx
p#Y6DHf@jDO:!% 	2E+,)'mR"9EF^Ay="l//y!]RPh>7UK5vIj+MgCs_!'"zLV_!Sa,*|gu]3n({i\}9$,)}s2O/&x)Ax
.*EB;V\~#4z8T!wD?6hE=Z`kY$Ap`S7SV>H	M85h
/&Q(p!_V!:O;0:A<&J9m!\Uch#7~E'\~[fbYBeQm6E;GubdIj$>ERs%D%A?#A:">B)KH^42b|e^60CvU%EaeKGg	<=3jS)367]L2BfD:&KZY=$eAa\(},6c|sg)kLzV
g-s<5L+\_bhmXG#r">,F{=Xp]`v!|??3K_{zH<~tqk.+UF$yQjr[3l6Oe|4X&AT8v/Yfqq+3ow;\zwR|=RZW*BHk!
GzEODE1j	v{W	AmY-ONY_/5f)x'LOWGZ]"QLEr--r# n[KkMA	QSS<7B*8TIg_jD2YY,Qy{y	9G_&sz<hn'SkYn'K6-h!7AjpR#vPNcp=zJvj8^,(a]{~b7?NxK*$H2+	T\H' <tXK&;K$OnIo.xxt&36o-jQJSNt=y(!Q?2/4U?Az5T2r)
F8NIrjuS[b[^j83(ENN:z9U)@)kS.c2kQNMM@(7@
b'rI/SL \*]y}Ff/?DnVGz%b&uQ*xg6AOL/wH#u	hdM|/-%}NPfr3a(?|
*dQ/\tnXLREU)sb"Ed4?c|E>0>((xRc(ru_xM4WsEz=@$x7gR}"t}jZj\&\_avOIt^%a)h9gy$f)F]OblR.\gjp36<LBs\_KMj;Jl0$d|iAe2rz4O;'j`0{	Gcs3Y&E$IBXXZ&
CSj58a4DxEJ:XK:^iB4yA _(()rTlbkSwj$Z*	(Fz;^-aUuL^*,VY7i@u7/:u~eOcNoHi+X!Y[mah(#0'VjB1;Pg37:/+A^,10K=ZdDFcQ:GtDdJt7iseQC %3*BTE]unyZ3Y.yS[D=A"S#KUK6n,]f_xM!M$4	oc~(9Pq)46X-^^*Saq_rr_7/Y_%IkF<c
`:&R(,(XX|?}2P- Q,6>(h[H()XYY~cFd$u4[jW-P7*VDXB92'PZgO1GuW\OvKUL.NZOE+YRPb@sn!]\|.6iG*q:pSN3PDx@E`q:Vqac:	L*J;U7WhKrW+IxQ,6iEo2|TC)'^)y#iYGp(@ErkI^!-k-wRKo+PBiwn9ua~QY~u@9ddT|V@$I8^?pJ{ zK+{GnFCG(rA-
3}|`m4#XhMli#L=y(MY<b# cpiKl9d4vd`\h5W	R^a#(4GE4\F_v^UvT,/)k:gRQF"FnnWf^(k91(:jJ Uv1S8Ye*Dbs\+kbr2he@{f-	CJ1eg5_F9kz@2[Q2mFq~>~B^c{	3vc)4h}G^=>'9Izg`MI)k,JMH=T2)v)qfT	FfrUFPVY!/|7/daHf9',	;n+['wn}`zL)UOB7 X!sx3_ZTDN@+K8%%_lY[F$T9{gb<PZ/L }4:ap+>gXz2!oH>F"M{vy@*lb:'T$s-XDA8|4{{Yx':k|6j:\	z%JTKVodye7|L'e\"t/wPF^xJ"$;+d(<Dfd[&qs.[`PW= ga9
&"XDsr[.{?mCx^2A%/=`
o@\~[S18,dE>$6eBN30ZRSp	h,	j!.0Qd2n.	oo@n.5`@6{CBzLMfkMH/(j`hv>pGUZbCc8H[?7,c!R]z;BdK%$2@"^j.%^{11lkPq8*1$H$@F=b0	Vx&!vf(7k^7ND_pIGjqj^zw,b1[<-f9w+BDOJ#b(6zq:.;<j[IKlKFI_'eC5,DCv@[@MVp|@[Q$kq/`7,"a5Xwqa}4:
4?9R.zxXy_g#'\O.[By"?1L<)u7b7nF%"s(.=9p,>y`j0Lj94soII:F}@
t(Y2&^pqyFn#q_1Ozb?>.X69oxAkB.^$0x[q)Q!uZZ|:='c7AH"0}K+X
arYq	~QM+ks>^gIhp;'(QS=e|9nrjr?Q
6wG5Kg+3Dr*lH(7#ZR-ekhMgtsjW+1`)$d!m-sw"?M,d:>!dWYN<pEg$%/<rvR%D
 U9S<Ogl<h:6YDE7ODB?0sY+nboi2zSAtW
`/sE4Le}S o$3|).r2X0kZB|!5N0z/a[4x(; 1UhLb8P>T	73wD,L2W0-2Q_%nnXz&:V8WD i/>-.?W}Iabr6cAT[uB]$kl)J>f]$j5+&3;EUnmQ	Rddzv52cCR9V8<`l[8"n:Z}03KXjANOtc\3|}.4G`l^LFAbd3o8kWHM8vl?:d6C_j#pT+[i%_q+{ hs#FL(zW^'0!g]oi>=?')xl #ziFy;%x]"EmGPa<ZKio]7_;y0az @BM4ei`D'Y=AL#*/QXb0?ogQvY71M62Xa6+'WNOJ3=&0m@P:UGCE/5Dl5H:V`$O%#9{yBA^$dF$=j(PwY]"=F]~/(n&'i6c3,,O70p">ST_fe
u1a!x=Ou0C0YH-Q~?3Xg1O>]..bE81
LVex3'1-5!H9m~ ;>;XI])!Ibe]\6)di-RM;qUlaz('y7Zo]^RSWi\J6aNe\[F,25@GOEm(3rtw;sWsO]6kxrbI=?:[3_y8y{nZnxC8E~N#K5kXMi'
Wy\?p5CE?)wQ)I10E;<Uoi{ N>]gh-\tNu,3AGqTN|2U'u%:Pn@WMmxw6uX?0<~O('uN.(3~.LVKmtjErKX;3M1vusW>No?qvt~l3~5siz'tMNN8Oe`M=c2ivlCL\:}<S0|@IygTFS4:Z)=SlyEG:5)	^qqJ_[mo'}^%^Ssl&,Rcq{=*n-b]-@kf0p"ZNb7?~C8-8^G#	az1"kwO&(b6M,	$=#r.|Gdn&k"X/mUhZwT!E Q?imT[v6Qsko|3a_y':?<m`"ge|Keu>W+Br!4|Q#Q)l1{KWKIN,{s4rL&J3^c(/xm=R|Cpx\v9K]Kv>~>
q1VY>)A]0b:"Ia;K'Dngn
ebL8IuAWwNcUt	5LRgE@0^+psq#U5GBb^ ~;nZz -Lz{tC5\{~:4r38(M;L-.|0{5qY4:Su.fN{3LwL>?|++QkA(wFE8{`YXaqQ
9m6q-a1I3DPyqX	|V22*7<pdbfCqa"*Jj 934ty1RDx\&rnc}wiecD{b])9.@Iba	"S0"5>mSc{]zY#n%DYR]3VgtN{huv)OSy.[=Urx'W,T|)!hTznO/:	hZPM~9+[YQ/	J7DuX]+Lg]-I}Y){fz2_;X.d,/Nr<pw\YfFh*':G`+lob
+8mcm0m!?wuK4ZwAclTlF+*zFiFXo'IT{k-^nm|}7.0LN7WC);'^7@$m'7`B}A|[hNvCnhtUBBWRgfwegH2B	,%pIs0*7w>=6lq`4n}};k5K^/I(p;#~Kw7PPEg%2%u/Qe%^^lg-{ky}'VxnAnS*T9wMCkwri,\iI/zny>UYWdr +rin4yDKyxT{j$a_-ve5.v9kKuJOyu`<:-Q;spGtdGT	*_3ymZu^|*LD.P{hf:%tL;$munbR(U}x:3(:4<K8i!.ct#wbB?5[
Z+5jdx<T|g"jD#dJ9,,g<7Hg{e^Mh'P<5pKz.6g7?3}oqs_,TLJ3_J>nwV}?9J HJUF$m(\!$8Ze|^i)#|~"9JT_1{(vRz|+J`Uc~Rx']2]v`W%L
.-!;G7j	=VHowasardx&qOn]LEOmneI[:i\@AhfLfF< t'v&4k$gc	k\|U^	Yo$Qamcb2HG'&.__b8tr(`TOhSO}gJ=6X?64:x=;oL.`$4=lYYYk<B,"^j6x_G"	}	Ok}"8|&mm(y9Fml9]'_@n`]TB!AX-Dy@2W~d5;[lD<R%7"fRLUt=`f85_&MhY@7\9s~4pL:_ D$C=`{no\[Z_kW.]j{Hn-,(e6w%zC<bx+6Htz$'}8=q6h-	Q#W0P4C}a6R&+KJjN/BYi\1?.	z	E9"i% K_+[+EBnF#/hivhd7D;Kx5G7iIukuo"ldWj*S}A&F=&?OH	_Kq3k~TBUm}qdFUdo#FI22t=8:s4ers|uJI?'p'
	TF7EGi)U9|{%0az"q__e'| RBT=d1@ bXzu_J8[(LtD;!#x5p+	Mg;u*u(eeb[wdl,}(@f]0y__0x5XN%kV]H}w.6EGg)&XiJ7xQ7TkzIatK`8!JD*8	nAJ?Irk"	/|9Oy['k9@7w@W8&O#
/I#ym'r*K12o$;={bJNH|f.2F'&N
c&;SHqXr=Ikyy|![_k$_!q]e2!Qpqb"r1.fqsO,Dvtf6jibk+dD bwrK$I+J:DL)PTW\E4`)Po;nA$'nt}f!}o.ZF;bz]Wg1P+R]iX\z5">F#x4t\k;GLViK*|0 Xx":&*Wb(&1ML^z&1l}'GDO RYY@3Bg^[|d4$Dat}Ly"LO9q~v	`,WM4&u
6n;&pm6rJsk~'TThG
yz9=ra:B.aw6u+7P5u^-A}+ NV8<-# %)ZHV<d>[^aN,N3}J[HFXJ-#qWga.zeMY,w`"jixfq?"^*cp	\4cm5mj%b2ef(F!JtG>Dm ((5>FwRoq08+4zIk3\#S{:ycN|y6-9hV,;u8QDGe>LxtJ.vyruPW3lt
^C=+b~3M,"uG)5_144x=rZgg3ncD8W|c\\oTeSe8FcK}"TPV_j5;sCz5;ftb06-&a]$]]CB!XvB:MROnoDB#>Dyn')A]5TXYQ uD7x#v	RR<*xSHNe9Yrn	myb1
LNI`'/1Sa~Yw*\P@#Hi?Qk%9G:f'VL"\:~lAvqe]^2HL:?(.:qiUGn~]d*
D+aZS=[Pw,9<Xx%uY^'L	GS {d (,WC>m;J!UZ&V1FVpp9USljX]qj}Mt4mRn<iP] JW)._3Ly	TI-Z|Ia=MV*|y@H|Gf!:K{](',pZ3c|ffdoWupkE]cPhQvCl, p:3q\0.#v/F%PO|96_,8FobvOsh?N"HxghWGmtdG'HM,(Ln>|-GtO$sL`6,+sh4tM"+}a(th%LM2aGcVdm;7otrW\s2ModG~j"jh&LcD`V?[j'?ud[h=),;H=bHZE	bLB{rbeoFo@>	hLkHQvp,#4i5y}pXe`Lgd}%.1Q*y )u8vn=V6:j|-09<+7UD)H,Yl#Pq.yvq^	GW$bsqK5 _xz/*meI|xi;pYU4vrRqtNs-8&p[1NS9Bp2{H/>e!Ygz=9}(y5KKtD[m+E8psv|_.LHqo)aN=lW1_/c|g+#'iv2]q.S0T}8-DpM=wA@^<!`h=Ne&,$zji*&2B.S7]=n9.'/8S]D^8$WAV+^4-&4Fx^v{4MFPo-y${KveA+,^6R:yd]eT>4ztuK!"B0h,P$50l5K^:pD1'K81Im@a
}G69)o43 #]<Oh0Coo(^VEagX+`P`1^h}*&_gEc ?PB,M0^Ldn7a:[:DV\![V|s	*B3eJP1/q4Cn
&"T$.Y_b!6.3HW~^[pF`h_yf7slu9g`W8]/u0_I7)Ta[<PdA=M02 CCgM"cqSY8 ~DbFDYd"
*lv'mDa!+^2Frg_3N7O9|m{|0L&\3u0T#9;uXl"`3k(A[9m{*##Qzy3fw,Y%3U. zlx[d**M(_i)\PuP,GQof	yl>p[?%4
}Y]o-Tx^oh,`9{5)l3'^YeY!P%/0|#.S\=MfE0:qO;useNQb|(":fj!]z_;bo$[j7m%WPa_`"(zMMs!yX);O4En;z;ST|P&DAq0mao*8/hRjafq:XnLc+L\YtW>3zD{;DhhC{99B=)f_n:B(P]Vm6RpviI-#Y2Os6x|p:\E08aO,,4#&Xe=bAal*;{lPN*;haR:/] 67ENNC|?[dFZ~J4X
>;{M9z6BQG=e0.7K5GGxJpZ%56pF?SRrqQ+NZUKr`Js\%,b@YidpyMT^p8h;, e}WC=E4awV*@5i*hqB*u`lZ<9.dL%a,Ef{qE<'XT}Rpd|NUmiI[vjWk;H&GD\D_G~W4^/>$*"`ZUNB-{Mai,Cob`'&d!,NmZv{&QAk/BuGty_hFc>11YqJHgtB/Uli_-$iL_L%kA*`$~0j8lpl3bvQ3=WP]0	2B:nWI/40'GmB.*Aa+ml7oqE2<iA?h8LfOec
)^	Xp}5m4WdN@KLeZ(c_Cx=s:7brIs6H_mf[|h^awYkGm{0f#tH\|cZ_.s_+To6QqmHLj%qT^Y,8+k_")0he+(u.Z4L^n0J+LSRjQbgFfRHWal<f{Pte?yXK0Xpqm<-:RQ{- MC*A^R!)A!kL%9x/}=I8o9!?tiCT_XR]b+~-JC%'xo6sPRTbS}Ay(.h0V$i2\aokE
CM&n:7	c4NT'c-h#rj^?w&=u
H>]R@/!|Y8fx>BJyP,jGi	HM7Bz/E:NlM*+'Hj+K	.F	l+V!vg;,vuo+Fv4qp(`OpmPm?9!{)CZykZeh
QEVB.vLiqDTx`q(kt0bGH{3<kNl_"q>UN3k<jQg`
o&8Nd=ll~rMOL0<VI2|Pk0LK+\ius>$UnRm1@{w*HTe^BOf#Vn8}6&NQIH;V+:
7/VJuJ*^Tz>)(yHTb;!QiNWZ!?(vW}FTlny_9$)QQ%GE4tJAOi>pB.\qY}FRaRS;qcCTs9McU(H#F;=+(~TXEYr!,*!QBf3bPY6dfK=_B<0`z$Ph|8JY4g)Bf!"B:AZqEhoY02_i8vk6Nqwa]p}t1	JaTXA@t$/ie|%4CC6yiHr]!Asey%k{p`ab}!x4WeFn1~\[&82=M#aQ~YtxUJFy"95Qq3eS *"8	RPLgy6x!cX,w%EF,wB,]qja,jIdR^{=fM]puM4O&E!7bv=G1}L{?&hidp]#k|f,3/v?mJROnP;t|oI9|4C3I4G_+ }]!Ftf7qSGE}dceT$IoGS:\	WDZrFP">-0T<3_z7
G6E:7djrZ(ZOb71=G<i#xu$+`$M?/<<]Pz"Sj&
0=%\:=s_/~C<PM%hKdu}y+leb6}DE0s,gLH(V^_Mb~@3k+_:?J^oP&qR={V?Bi+0
:z)H!A,K7r2(xEdG(,#*"Qc4lJS*i2T*;^l)
5I`Tjb{g*XC.hR(aHs:<g@GF_e]*Au9IyaK##15A<1!`>,)	kO#QGT9Qc5;Y*%?ZQ21Mvg}{5$lsa6^{VcA/cZ.5&?[UElq~^dpHseB+gt{(NgOGq
m[=[_?:X$1M2plKwz!g`}C.Q>W\c?yCjQ8NbAV7(aV,>/HL#JFB'dtj+[]Ss}	3h]5[O$`c$@mtX@k3Z[wy|pCn!cp}Gd|=p
zQ~lf =Aj1,e:$kaU?P9X'mnN\r|T)It0=?Mnh$Ad~Fhx-!8>&e)f-'%~o5*Ts*M)h,@wAM90?].NU5b_lh$1RI7l*YQ;lJ+RpgwJ;yRQ'a"I*)9pvt[cn/M4G+j_R#L9\"(1Qq%Oq"+^@*gyMQy8B}GBa2J [PrR!$,(\F&FoKJxL1!I#-B4dv~OU=m1*u${V _(h7G) @.SSw|JV*;+rMA0\fEL/05ev4o>[zd?"{&uCg&0|.m5m-H?qb7@-L^=uUs!v+d]Bxgw:)~	1:fsY=g!M#|}3!RF[fQjn,N_F<od'1k}jJqeuePx@W+`By&WQV3;Lx$h^sf:~}l+WNp~bl?f;6} 7;3<@%@nY\00<>'l3|~Lfm8iQ7G+v3`|"6?tw"5TzfN=Mys>ZRW$zG~2Sc\DUa@N8LUG}<Ag. V.|g1
1 %.1w$!`EGFaVO7=GrVm)=:sxvsW?y`w6Y)4Q-Hmj{:`t/l7~8p`'4Prp\)+,8st)`{7s1(#9oRzzbH H+Ta*N/*GWn2?%:>W||D`1G&T^;ajH@M#v3O$63e+syn89XHQX2~s.k/r[6DJ\
GGc.!Nt.'u	(Owfy4+fHvR|3jAHehO`@)V+5M5=m)_Yp\v
]G,UA>[-s7#&/RYObfm~dg`YRNXZ?I|wQTIp^:~Tfd7PJqz'e;zqj;D(Sm_YRjn|c	%TB_]H.D)5cU9kiolk?^d
^1>\q%^]fy|9=.HMVGb?q1*?NBqmN1LM6jo8TZAOuilgz#wR] 6~y,{22,l<.k"vKz9aU/P(<EJ<,wTdQjwVvWTjw?uG
0ab?]!	{f?"
?fRv~tX+Ue2cv=]!VGPY@.WwXX?aAS/wGneWz%?-/wY3?i9.jnI'tE["V;+z#h<!.
U@ -Z=@	,Y!IvNfQ-z[/g3QXPfJc#Mf[v8S\j;7C-i,!VPg`+]b1Qc=mNh&"0z}Y~@*	<hcDoi&ZQW$!N;L]zX5pJ:<C ?q1]v4%gr[vx{*uJE)K-0!PW7{?c	YF(X LG[Ou9`7>.+*{)do &:6xX>Oq_" kn
6F0S\9T?X0E$\~jB1mO?jM[I}>G0Dt]<"!t+KR	z*bx5Ls95z`01A<D	IW[zt~-w+5E/;w|)]6}Aw^O?g~sv^DbZvNMBU#5R9Eh,`1._+qvi>@t}D1H2+:l4-E0
(gZfUAWCE21xF%{Hez99T
Rt{}uNH3D,$;*	jP+	-D"ZpZ}k]XuQqYeq|kt/ChsXc5U3.h&RcqZz.;NdU1Rv5DDf`KibQR20]&pJ(P
Su"1 ul&f/Wn@f5z,i<S;D#>G#3=-JrB1o37`3xn]|P:l#d?llTcp#&sC=OV;k@M>fK~	u,#b`XFa1S[(/U)8V'+P\0|};.|&28p`VuhFBuzDiuj:RD|;@\#t&3Po{"[Dqm;jX^5;&Tc1Ec\sV>+3YLHo!]&Aj>_Ll!{?p3qT_>"p
eel`>&Sb_/%=?,gM'8J'%d}e}Mo%4AJ|,oTj'$Gf#ly,ZtYt^-k8]u`C7w>~Bg<E3J_ 9fUJS*U^\O7/iuDC0@VMtyKAwG=lqVDaN;w\bq6r3WP+qx>FC;vH ./G;)in$`+-mv7tUH'=XW&swDe%)VbLe	Y#cz{WgZ_FpcP5_gjS8FK([oA/G=OOz	rrV_~q)(gi|MkxW"jQmMF`4I*w$Yy<~fv+xQS1.<@V@0Kbxl1i?kn"Hgku{$aS\DvB%qok]xg'hFQ.v4 U!CT3`q0b%
5_ur*{[h02=n!9pkR9?/g.	IHO-(%tB</ct7dXa}bgfy3s@yNY\rp[F!~l2mm4bYIdA0}m@CV
dlnu:\<}f1STm(Zk(XB]&o&H!'`NP	3':Jo64.BREaT|#"3OH_C*ysYhth4h	W:O.8X#C?cv,YGtT_Y;e9B"[{7N~{Gf4rG)3dR9}z+p+3|$2-lX5J7'vI<eM><YQB}]hPZC	lU^lBZ[+CoN(Pm?!XhI64`'3bQ%we/.%x6?3<w)JA[h9tXPr+3F~^1ti=;*h"cq,neXx[|?/(\e]&cB{p[h06Wd}5KI2
>EVR4v",i(mj9S 'R dK:?FQ\<8eJtMmg\ hN{]v86*[
:&nkfOC*Y&u)AO.Y)u(IFUa@5_B*)b\]i.RH7kILy#h<X?3.R;dJS>_Zzp'?WGKr#9 U{#Q5gtWND)*K>	aBW6YJ[.;eoUk/i0C[#
w2)F7w6rOB}/JG@f^`-	o9UHwxlhQP>tZR6$tSzNMrI\~CMM4e}8g[)0iK#]+I5tP!Yih+*.[]>*v_HWI#ktvrE>M6jNFwvD5|Q%"m3CYV?f'A,]DqOq%s>)EwZylN(uW;fh\t<W}N)bc!r%snWXX'7$griQAB3V 2"%&pQDSbPH>\`gG.SC@/]Y]6n:/z(_f<i	;y ^{Gtmrr*D*}_;
mwA1yn&k3tJjnAE:cw}w`Z4/7=@!*R|u'9'	[*6\B0v;o0\dc9I"g*\?8/jOr-)*4=!fl0Y&%sDR*7bVXrY=}5x9j*R'@IMqez_K,^wmId&-X=+#Jqg#QsDX.YPiMa~{b/S^97An~z=Q5-a0}G1#2QkI+<j0I$p|G~[
{98b7+NMcx]:@8V18){Geg-bS2.Hgg`X^;R%phI2wO7:R-{e}XmL!XE"RcBHsej0,9TP>;AyDem'`MW2.!oM1AL1%{T|T+43RG4#B}zOip\){>g49b%qoGg RFhHMM?4jo"N"xbkcyDl)q7_x+{H<}W@#.GkTg;XM%UI(CB!?W+-Z@'h0jyuQw(8kTO;ZCi+T$n=(?D!(@q'&^iVbOw(L'fcEVKgW$ON;QNaBQZ}5w\Z:KQwYfwAIxkwbeR6l/ :SNH[(P8Fpc0LR{k>Rs/(wlz8Kn])	4Wo'~HKetSARP<gYfW0fx}[?^h=-BxGz'Ox; (MVFMu$n0]+?{H,6Af@fb98w6.2dfp
;OPb_>lcFg&)fpP);Qa+s_%'N/];W)z@>'Lw^%()0%<CP-KrmD7NU7;H-PO<,8w&<`PAz,B$XD~QHnbZ/rOWg^^Do5zaL	{LQ"zPzm[c='+2w/-oB#?U-Y$DK!m _>nAX=SCmi71EX"0}Z?6"nO_?`"h~["9~mA[3FR7mFeO	b}{ohfM\bRYSxwkc"9QLI`((0jAJk<psMGO	Ft!$kD	@4{FXwkIbnUQR?K.5F:uB
9Vj=
n	Rj9"
yD|PAn~*|"OmUo'9y%Weq#IVhR`f.3E+fFZ!-	yKE=~/NzUJ`WyVs8hV1uBZF3CJ:?bcD.r-t:Z*ZG%eYn98Q^U2V=S27.XC&|#1)r]~7nJ']C;jGNOS#=J_t*CXCSn{G>NY8g+?
?@}MS({
JU[VCgUNUWW.0rg_|s@``bwUuoTfQ"&S[ 	3+G-HQ@j0aj1LB3wG;7`Z0e;x/0KklZ`G]1MbJx~t"?K1#eCWI(AFVbYgh9Il<_(w)F$"[=ee<7'T%mHVLEWu,;0a$C?ysPNYY91Lt.+UO~&(&btU~)FB$m,.}&_Q=Fs7\IM)^d/78ty DdU5Ul0QRS7]$tn=4pp/F'=iDL)Kr)J>UUGC5Q|$Q[dHs'=\:l!sbz]mBGK2gHT^'[
D8SO6V(#cY	Sa:.za;SL:>v(;+U$AT`y42g4V'H>S3;;Qm^~8EeZ.@z$ )n
uz*jDCyN3:( %vE10C6
 pt#(9'CVGUO9yh6pFi8l4v3%^#5gz}m:;p&h8{YDWSRmqvrD?7.6M`(}7|I7GH&&K:Z?.Dc><8m+'F?g0_jkpT(*aD"760X[^jlu!(#lF.M5eVZbO6wWdEf2~#e@mh#?8e25x4)m8ImTL, B,Ow(/H8gODDbK'PwcRs#gpO5+LJsjH8%yw *ipC)4:1VcAJ2)4M_Db#o_Sz4X#[cXDq|t@,=~`0/u(}0O(dU `c`X$[V9F;*fw8dcrB(RW6w*LA\r	"&?YHw|%
!6LYSD++' 3(a/QlXw#[`$(y9[C{nDU$4ch	lQ&5R-Gy
m.IP`f	l3!M.$%z*gQ7H
pPv8[u`m+{NC9QDAFoX0DF{ (UYw2p89;%Y}u3MNnP)x;*W)C{slt@gWk+F`O^-}xsbEH9$g=\B[x&'RF-F;cG@tv:7O`x
t%KzO@3BSo[5$O,>WzCH;bV\=FgcK44^<;ADR< b\PP3HWQ'ngONRyZYgY$H|aS)4+kZw.MS;Zb Rm]qE#OESB(2VW\zt{)xr7aD:F3od]vr=)2}\7	Oahqn/\"dJ4"W(.Ccd9`s6}]1yUnh'bB8}vve8?r@8{vkRDHEHUAN^oRzjT2ZwqpN4BAoj_tX_ &	9q
peE
9GAz5'#yRmRSu#"cu\~`6Qux3SPe0dn8 $2*L88HJEc, *WXC*LSk]  }>7H+yJ_r@o\/wO@zUVC+}*r3I2y1Ecv-B'>"q\9z;tk`yC@}a/|tnOHfe)PQw 2nk}Gj?Wo;gNtH64qoBmv<dj1
Ez;v10TG!sD(S'[zxg,JK9xvkN\S[QC}2'ai9@^"4]Ha'N/o461`~-.*auO5vHs#C8932$fhu|zcq/S\wTT_pV:eAZ$El7wUFY(0y{8<ZvZ+
Y}
np #vihsn{[fIA}|.bm5H)G-x`o5L{	2"kj_
,xL@ktFlsRsxCi|TUx!m~#7P^.GhFb4Wi=!pkCYK+HkU(JHe8O^!d77cD~c-@^`X#>jr}ZQ??.N4yg%,}30D5&*c
v?4|v\|RP(MTn{C-2U'}][zUV(
79L2>]	V"uC!9;utJeO@gs	@)p~%mU+<K\#`\ayg 7PK.}0\P08-6|F6+B+ZMbxn;VMIY}Elf4LGi-pu_iCl+0dv-xA,pHtNl0"?PCxPUO#FV-@|LKk,Ge,]4Bd.TqNLBR{/==z0a0~Sz[Ra'q1[Z.S^!%7 zBixwfaDmsKn;`&iPs2;#^692~"U}oavtxkpy8e&Mz*{9+$;@7u*>xyIr6Ab]qCHhHa!bZ4X0[K3n?pT(U@]Hk]h\k)J "7zBD'yp2gawRn{RQ|CSo>};Q++e=}Q;:yUM-+\E65,+xv?Dw8Yja
{&Au3Ir%hsuU^gJ-#olps/O)1aES!F^]8VEbkUc1k
I s|g=
}J)#2.6k`
~%$/%5M)M>Vr05"e+*Oe*8O*z#k#|S#sPG{+b}&|-zTfW.\SC{Fk:O/*0?}$r!@F2WcZQ7uP*z%`G64)N~`)PRmH!;^GSIz2uY{DjhwT"KpR2xm>C;Q<wQVYF)mXU{Zj)Hj h4	'x;^uyew|TLsAcMkP^',~	14*~TOD9ROavy1BCb}'uRd`CA3r1-xsVx&!B!QE$\nu%Zn6}Ns+-{qn9o`g`?B:tF''Wd)Y^b8*3jb[k.t11cR?
(]He:7O<EpGc\
+MIdugXnVl:R@!Qd}#e7bP0,
BlV[C-5]Rzjd^:E	Nbjw5+]V&O.%+jG{WspOL=p]?N%_jA]BHtP}?\,@
"%nSR]yBr9/';*[U&cUp1 ,1VE-0]2BlBB7d|y\VT(.]vI0F_j4}
SO/?N@p/Yp/\Du}r7P(yzesuM%#c6<Rb*luWqFNh2=:O\!p^'J(p>|-~NIwC?Jf1c{DzZl69vQ@)V7SmJ}
k=Bhwm[#uB@@z+"4]{V9dn;X1{;*otgk/o4Yo6t>M++]|\$Hrv{qg*GC9$}$&qid/3J0o[g!45,!La^|D>t'}rrvc'A?
c8$I5uQOVwgx-(GBOf:{S:vf*~O9#Unj	G;d{5J)G'|'k#fi-$fSF6I1rKy' VPxVv%w6]>DEA|ZUa-R_Qz2,``jvv1;>4_TQ;vY(xvPXb3=?u6LyvC<`i=`|3:	 0u`[ ,cI|qkese*?9Uwn7U*}KkLXun+T5mw};5FvXbk_a;;dUjV"7a
WSP&d_+mhhM9=?>_Bz5x7= qwR{kzC6|01Z@Y	B<kk$iG}0~EyOl10~'hd"0>#N.c'kc.sq@&AcR#*r&xIpXZP$Q#beWCL;Rl97!-Kj`S=!i\\vtd0veIA%'Uq2>\ojg&wfCO BePxz.RF)8Jng/,3>FxD,QB/ I'3z*8X?EIi_}to}6
NWx?T1x{S*rp&QF,f2de%k=EfG-?<(L;|,DP!]qZtHh8:(]N&;v
QR{l+kS$6M	o^w^2*$9QIHPmAu$#'*Wc$:rb$JRdpr\%yE1w=-g#Dz;odBZ0.4	K-!j{|Br5Qx7pYZ	)pXe)@%!dDGa1Uw0:0w1IPtJ8IV^ )~.f}<6s'_^k_x J}u5;4ELK q,]Gy$k4feV8i;q'30Of,~YXIQV$][wMGyD?
N^p/\1Xbry3yf
kNMV/id	JUa(
t!c1[cK*i&B`63Ba[2k5He:	%[ScS.?D7@e}=rZB?y4	aE7,1K/y_1-)-hqE(`Zw"\@[?0w: Q>u--iWQ"s8#M@vGBRl %qeEGQsGxiNbu:B#EU/wyf\4FGH<e<=Qiu50d=XxlTj^.Z-`alF(G"7=M"]#Y99m2*6x|#e>!:D4?|D]{>|cK6b@fZ1>_='` Od<'$sr7)83r^l/Q@9"&Dj;wHYX$-y|iG9yf1eF3i:?Zz(+^5f1zu"Q,{"9!LW.+QaA!&B+#Y9F7u#PuMywGf.)CRrWR%ZlSm"%LOR`|(a[Dy6B2LM~{f^4iGt/{|3jPekcQZl0mZ6Ulsi/8rZ]#lak`6Y~Y\X_FXrO&@#MtQ/q]=	I<n/7z'0>|fE?	N[&AJD;O (m[??	o-5ssQAr'"AS@@XM)B@B@qwNP{J)
Sg1TgFBQ[i%wJ36v>&HN'r@^Y[*
c=yj&Bh| 1C=6vj"}LL6:GRvh'Xv+Y"HCb\CF>,vmj$.[8ZfTb?(.&q7MKz?@4^fMF%AX>zA"F.hKj|2a96.r5"Mp{>|/'xpI1{fld!C16M]*cAAJXp)6s^K'Kc
CAa3_Ouw,$t0>JM6 =8aod^'Vm-+i|BYk1zrDcnd!g
JZ{fa)k@O2hk%NL>orv{8yc):ogugMz}YRqrksr*I+Ntf/VV>z#z?gekAr/{;8g2a8a:?eACf.c=?X%y=[6<]O@nZp]PY.D8TW$t#?y+o]Ebn=7I#*;+=]vS$eEt`>Kb{zqqm\U:pTj68
@V5C%^t8cUQJVKMSr%_qvJK\eCXSIz;A,^ XwjE}G"G^IiI`)Y&5qZ7<XIc|o]fw{Om<#s?#lm>DIs~otb3l+VW39I%ysn_Cf9dNV,SLVxH0f:xJ"kO(;tfR/X@1z7l=.+lXJ>7"!U-AWa)~gZ?]Nk~3+Fn-QABSYpIO&4F ZZ[A-^_?[s7q(^/ekoD
({Gz&pckwysNTUF,J&MQ0u,`D2#9-kDYW55$M\]6rd!gM,B"P	[9:<xpy!ItO9#WJ]!A,=Se%vjPZ_9ki)fc|oq//-3V#!4={f	n-u}oqFS06d/O!#!s$I8MhxU{~eT5~gUO`B^ED4iBwK64Cj^0ORKtO-?S078/2:W0m9w5B\lOQ:(D#nm4Tlgj3"KtUL87/u1O1NRcg0f%[/tso*]|r8`('Me\>U2)
-q1\Yn2hm%A<v.P#SH{vBOG!cx@|0jOEXT=qGXC=&'L)Q4KI}7tu;dON$]bVo Q;65QKvIZXF~){z*3S{`I'1>D6m
K91,$3VP[a,|yA_j~~A@"`^i%/$YM-NrrD1tL!:_c+-ws|"@	X*p@>axPe<	"[2HcVKM<B>2
!:3Hu 3>J\tvY6b
#ZiXU6?\3K3;
RIG{?Sjz46U+O?h2kE%(H##^DI3L=k):9c $yc">Ke1Ab	,M'-'."ZyW8'Sj0brzOH&1(}'EC8 6R$}+j"4V!V{(pJl~A.R~Xx'_\'|Lt`z7ho>{&Rt"{FY]ZN=K@liso0|*9^>NV )g0RFH,t/rASt&i)`gGW^-%[M/Qi@K_~@cE>~9ou9<%Z18L_Q:Q8pa'/< 9HpmE8u;y^l2fL(PlV&x^$z/8P5C75,[=!i#`EvEsIb2x 0Aj6u0(,EoCj[w|r+2]^@O/bh04DD^ENm",Bxj1e)Uoj^#*a=9m	zjwk3?JS?Mm[I$H()>\TD=ehhpUm\%!S}5
+3CP:ntC_+;%j6 &iu^#8T
:Vi?D!b+5
{&ud`wh2!%,.
+BA@.NQfq0A%?P?C:@d0Idyr^[xh4-#9O@f6P/_aAG~R(,Gd{5UwUJXcyz.F@!
>;
<j9;fSQWA;$dP,K@Q2]{`"md4cRj;Iq1A_M?v2U? v7(AS+(r
~Y?\T7_h$]'aU]V~$#MWiB@E>m];cX@\<s3a<Q&Iw._>/!@lO(/!H.n/Tk(y]p^Jff!2:Jx9CC`X-%<+Ugv%Ql{hY!<HvTG~G2joGQmjsvej,W+Xg]v@w
kORb1-P]0DVx/Pnh)%dvL;ncI}Mwb@ecC5lSp	/r{uaZAC,$V#k0m1o;3z~G$J)
v$^scphPy!X-Q??IrX"=[effLVO1}
h|6n2gGu'>IrA)F(f5X}MlBXcK$7N5UeF6Jh`o%+(W>O{aKm<$o7y$5R~lWu7}<Im|y7y&0e}[5h4G||OxM"WKVpz0&mdgLN"+\*3|0H}Ts_DN7r*s\pC5pg\-`m$!D@ e!)uG*4UWI1O0Gk`d) 	Efk])zdD>9i)qs><k/O/gC}N(STno?nF_C`8iCemk+sVPJ,Ofh.Cp)SB)U|>U|9p5o_^'=(;9i3b9@
6->9
@U]UH_ (4>@T{SjnC5A1,$+cW	\#xEd`R_c(3>0%AW78bgX54R3"N =F"'ghs-t!"l1~"CSs]t?]#K+=w{@P/@m&8r*!2Pr@|[zR EP%
mL42NMw`~CR=<+H/n+Cn/m1n:d]mlA<{EDnA5T<Ud6/6-U 7(fOpnM:RA#dXE:i\zlKbB:6c!UU	EyTD"
d>k1&~>F8yJTG}[}`7K-X}$9^Bi}(vFJz(5#H]_.D;BJEtcR>(x4dU5v:g#A)haH@X/!muk9Lt( YGFfy4/Ng+["O37bbk r$"EQ`vZGiJ.7~mFlke$G6KSs[3+*)#da-e`xB]</bfI{i)MRs&HJ"SVsY\!f_[=Ja%J*[29cw]TBsE_RGJbmi>f.vkGn
=UU#1E[yqwQuGbBVU13:2Vrno5,A&K#%e`K4~q~6;Vm|`@@L!&mwW('saD`%b{Gp8yZK,PVGJ6u4DsC(`Kud\1W3KmA.:i@!PLN#F[Fv4Er?x?	>rVCoqG7P8u}mWgApMv^s&u*4|sL<;7O!8=oBhmOH9I@P;Z!?Iqqisa=5$>$7)N76Jd#| R99"|EnI4I~d)c;%:[&^hySD&z,otEYCxsbGx)sK%o\'0rX{~
]N/s\_Q>Z	0ZuSukS 8rq^L`QwEhAKn5kQi)BUT@KC`q!xR0ejHxMSZ/[`4 h^D#mH7 ??Oq$IDg	C)]'?ti5s3U^	qt'*HcVw(:3TC	'z<9\~,UZrP(}83`lb(WN@r7S2nzj	arw-.+fPK{B.[]P~s0\Cm#JX=K7?
U5e~~yXK_AWJkX|Yb:ts4/!n0C8:B}'nD
2kr|P\"_4=:_&ez% I:u D4\o?6|XyP\Cy;,M/2$ftY/v6}RDP	9kQ+?Zq6F\<bV?^u;/y4P\Fs#G"I>fKGUbp\[h#.!-E'^Md0%o3?HG=5Wi:!# /tx0h8#yyt.'t$#?8rcy?@+)2_"?GglC{
*zg!}~2{VHgHD..a<x]06-Kk^&=w(7GhQNH`A.i6Y?Wo<.rAu#(u"kYU@q/oWHC1[?cOBzFh*GojI9EBi
M%v$FX\%0(eML
,|MY7p?k"lCDTSpP`'f~%R$~BWT7Q+FeJ8`A5Q^t1 ~@!44/fy;YO]{MfS4-~I~7H<PDDs.d'6Z=P0SvsT+56Cu0dHM
+0)TB}<2k%ki-%t{ZAhO{N^v5wmt4Qa>!/F%UwebGaf-:(pU9cDwcbHf86IpD4;eZ<^`*`Z%#lpTaU4R@h+<Y~N0d1>2UEc>,\O%EhFDVN4[^_VN}w~1/wX"uRk/U'5f%hY3Vd.w
`C.i65Xw1^?a^kU8plK	iu	o~uY$AP5jANUac0	?GtfXo-%vgb:ezgDt#{
;DV *558v1=A:+yqdNSx!pwT3|*rKVX!'b,t	KB8peI+-|5g=Rs~m~PC{JMT^&72qOB<6}{,5+aLfk>]EnIT
C~1;!B?Rm{{8Q;1i1^c3Ct8x"b.ClT)+='[\F04-:LNax.=o. 7M5yIC?T>Zr)'b&@IrmM$Ei<wGUqvX@ fhd-)8F/Dr!4mt6B4EJ6icq,T2$+#M flo2W=T< Wn*n:0B(,<CfQL7;1y1Y	>GoPsRi)@E.=	3~w<iWc>w>ccgza~1eDaI/wzFxQ^gf9PITSw
k+	@,+7MS9V"ik,^i)\],.CfeLn\ACj9;{+@M:3OzS+JY8seU\poFgyxf%6YND a}3D619` {	EiAoDicUmK-(F#)T+G33~gng|le:G\(y?\K%;"5#v8&</a>O%csK+dLcJG)un4'S6a]/ZtG#U	V%7.@
H-"RG$Uou{nc!`@Fb raYz	f4(@Y60;ivSX1G4dfUres& %o2bLQ8ZvvBrOvd;@TZV)4Zg8@/J.]l 953#0M?S$~}T\0uG;5<pdIM<o.I?i,#0ti@ccH.DB4rQ']G9XB5c;G]%#~d6Z6LPvz[6mUo;"%e6=W]@(+pwr=ZC,r={@;vlS*2j>a- F$j:NX=[#yY>a1n;jt-O/zdhyYQ[a\cN01<xVNz,x>YGDQVl&qJxbO9~IwhUX-pSY)W$@;JNpL-xWHT?eUBgKbHa2P7EzOxDgqm%Ye2xz\g/:h$^S>HvkBhY8S{9JvJLgOyy6AvvMyW)<p{OTrI*/
zD?|yxC3x6Si>&}M~h=2ur/]|3o2XxfDm,b~?rlWor0@+;f.]0tUv/,>r#nvJ01ggY@J0^rOCO*$u3+b'"+q_!aR<3;4	m}"fM|bQ{>ua:ifwf"tI4{$N',_Yd;qseO@^+|.i78v>)
*LN\,bbi;Xi^_iDG?#)#=;[}cVN]@
gozI}QAI 1/|0h33C^1\BWa~@q7t4#d\-a~mACBSiYhf~:wE5$Kx)tj*eaH*'je}~kPE162	7%mC$JRk1j]P<H,iC4B({U	#fku$4vbtU:KGkP)M6(CI}Rr{3yT]vEwxl1X:~o!QWvP]T8EdOM'i>ioG+'	iY-QaLDMWZkkZX8],:<6VWL?MVVG|Sb~iWuv%t&1]Zq+.Fttn)jb
a_?e'2Q$t#%aGESH_+A f
~(NZ"
V*O7`M0wuX
KeDh
Zs
=[q,T[W3(y/"H%0NKq5]iXq=!|>r{]Dbx:Rs%$.s-'r[v'v5z},agW
a\bz"@H=Yl^dY2y~tMT;HY{,6tV	78;He4_45T#[f	0KW~FAs8qnbCS5vO~'D^o#YcfbM3t<A,I9GnM&lopumtPJy+'drh@|'	1O{i/(JRL}500nXI^kE+!=&N'3Z^"4gVW Ogs_#xrfo5ya/}+i,n<	E'Eow$v%%}k[So8_6SR<T{OCot6[$gxm>`[Ll+Gv%sa/%FI#a5[kLEQU/nsGDz*IZ[OKTS;0-;[z$OSBPbMMD!1Vct$;!E}5NJ_\^SfF#7"C
m@xEJLB~k9bnUx^ HS| Zm[[~|J@|)df'}%B@4\>,zTZn"h!(nU4)E$PSZ, Lv`St~mI|"/X~<5%?Fc>y8s,#_{$_kmumJ\+i91X_:GvEJ&:Pmd.qr%
z)9*Iodq,E3hfX-5:ZoRM)"}}j7IZy@?m]peBr7tVj.o?B^W *LqEOe%W8H?2{hqu\;[Er$eGLm!,?aB0V1k`0-L`Zmh5USE9 ]Um[q/.zZowgPzp53_$1dl+)xLzk-zTpQ8O3S0sK@W[_t^v'[uFMoF#I`	G\X9sKR7EV{{0KLj77@cZkP"(k!ZKC<4&""NuE/N/$Q/o1x1:=xZv}1") ldd'~nd6%C<(2X`~m/xBy.\B*L9*
TGhP*P.icD)^F>M ;8g%q1-?E=5"oGaqxhd+,3Qd&IPY
$pZF'6{~Qx
;CuO3vE#->UTQLNyNy8}vB6.Pv:cC?VW\Ce01cN[C\4arxS
[Y%	s1#z1|{^EarVeE3{TdPPXnh}>p=%si
j]#P:O%6Zgxxe#V'UdVq7@,dhq2mX2u{G4ge=rsWY.'n	nQ`<Q1O-$B7:&B</MDX.!ThH&MkWBiH>bkr#. K{g0@LBeXV.GV*'IYc==%gD2|yMq2|K2:L. X`9d(XJx7<kG|zj.O96
Y=F/k22!-*	{PrB$0}s +9Z} #i$xo $oW#Q-{G?xtd*'MbKh/q<WZ,M8Ac^c1:`LeG)Y3O	MjpE]l|I`tNvDc=%'H+[8{]d8ALeud>D[RK-K 1w{M6Q,zd\>{pq{MZ0Y(@RO?OWhA
{iW|R.!{ZI-M*cdpGCQ$`B"lndi}]..&#$xZhr;y96t`	xc4WvXEkVfi7:v6R"Ebb&rif25d3 wJKL&fd*Kg3v_<8Z3]0m,vn0r(&8Xw)~B`	6>Z
.MdpP[wV=^V)u^7:gB59I7kok:p9kUD'yrw#lwzUtsZ{9*]_EMGk?qA#,ucgNWsg|bWk:ifQfH"?-9e{3}8%:j\{W(bQwy@+<RqA[G^vt+L?%AyKSi$_u[w0_z"]a2;Je^m.7Em0.X>=[iD(>S_WUf1QTv=@ITJo(?W:%Oi/T!FY2+r"$`OMow6w4zdeARk,A$1X$iw2ov>X-1ubG%iWPNP%ms0z)6*	JoW(&4F*%j*|J%}eG~% Pn>,Tiy[g5|{aAXYkNJXwXz.6DoAn0y$f)t~c|;u-yP5?.=i&gYK.<_VR&*CUU_RaB[UDEr[`
j6[J^R9i+v5pZ\Xm'@RL%N=EYW(`J{'iOg&B|OY6@t1i_k]5#6+RbePm*AQb]9a^}tEw'Dw$Brm8f}Ld7S QM~}<Em-k.a=5)I5<`QaNk,6%/W54[Ne8HC2mdi{r8vl'Uve]oc&3t<!6!Sh;zatO+9!~ab?9KEF~MW?%xJe{3~w%V!K9Rr]J9acxt9ECns1Zyp_&:LoQ'`'!|C5mb
"x@xc=td'0iS	K~R?B|4k'<(mF83&G:@:y/>y{DMY9o)N9a$dE:73.P7>6'jKc57K\0'vc3S'Xmqcg7TMsIH4{!DoATY>9bZ3]=<>}Ec`Mudz[(WF8'>LBAqy8Oo0TF)CfLJth!V~"]SwN)qWhD9aTwG6v1Ii6QH?KhQ\c#a(j9"veX.78AkR#(m[_vFoS$f$ocHB4fk5Hk]A@Ub)lseoz@ ]tt$DFx\+^\<:J1<I[bGnGWqF';YqO0z*SM"gji44edY]Jw76hy?olcxHY]kb|<1
iUaq`kd0lp08b{B7<QEY_zis'q^9.Su~_%MKETGVG ~7{DE-SMv%:E!4AX>j''d\I*nuLSpm=w#z/,^|Lyv)3D
I|k\5n[|yAMC~{R2YN8,YrHmV+M*g}7*VlYi)gCMh1*s?w[rD?4TejOgo&6K`bqIZt[8f/Zlp|W,,lt&="sswNBdHG%re9;2XF#\XH#W&{p;3)Q{7XvmGyj-[R, k,+;dqW{HAX	IpqJ(Js	1KaSH\_Igd2?`b`b h]Z9Y`z&^y'Sss%G:jvY-%it9D|}_|o^%L{r-Bf';SnuS&,1W^j Ru$_d_S*6HA]f{oZQ>whIu:F7c/=wc_BEgGr>MY<F8c'oNY?H#o{SemN$Gu[$(.SwYT:<Ur='$`5/G1T	HLB(D/<h87).jEqw
hE}//gJZNAIh)JNB\{mNdUz<tg2	|d:gSxd6M]Q#d5/ow?@7)%bpnf{St]nI
}3Z+dC-g..F&^,o+_s.J(i"3H^|ZlV|^~2[Y[.R@wzA7"Aw+&]	S7hE>a`l>6O^^cJY"QIK`84);FI01qm&3i	0qWe{k-Vjr&@V%4Khmw=*D(zhW>W"CI.Ga9E_H)*6BF_EF z3%JAu-1W,sr"H2vcuAAeAKuKU#c]b5mH)A_6,([gNWV@lcWAmB)%o"$h_(+me%)b{vhbKI[v]xyvdM#|%EjV9YR8@mvzd5L1x@pE0vNd/uE4QC;g[X*;5\>;0,I]{Lm1htU[Cu]le408d	0^3*A;a/Zv>QkXNY027IPIoA&aP/0TL&}'l>o_fd67#|ex7_qgECCK'd7s|k A[zv;K-2w$]rv>Pb}n'Z=> HrtfMt?"Nea$]]Mc?0&8mrsk3dO$uY.At	oQ;sw'&+~kOoZ>f)l5Tvq<%gD}#kK88!'t;D'rO0R'SR2x-ul{;=B*d+hdE
]T4$}UT{'H6dNsub=iL3"~g(iM]5|*tEIhQxLyg\O`(%a)];2D0/@:.~VM_p=p.TB}Hy+01>#:1+Za	+hzKE'oX:;{jgcFHW9Y^o&.{	y*[.q&IgCGfth#%<;/0zRR8j/+u? u\HDeG<@l%d^GCb=JHE;FpGMrDvo/6:(<,:?46	$yPH7I+y)!y"M$<c;`>?4KZ:2U_e%<;9VHn'y5C8D/'II)4[Hs.?nTQ1oN&U}Qpr~tx[0GTi6K<zkj^RJ"c'n4Fki5Z&IV-:#H6.zA$W^b!.R"!i%FIh1"9jvK	`WuL27Hw2ig#>/8PJI8i7RcSDO+PI-1'&I^ hz39nV26Y]XkMv	|lYGm?m+Px\xJS&{8:p_Hsc/W8nQvaY=bcG1K3^Ln@+|l@(eO(G>H|,F@6 `	Ney3YbPr\l+pl4%=fz|G/<zSscy@wwz{Y5P1>WS6zWa*n|jJY
Y+GSds9{OA7Z!b-B=s9Q8]YH0v`P/,mHs|3q41 <Mw\"2GZwWrY.O4Vshg%VIzbj]KWP>TSE$
}r2ijtI;oRF-Ve;RWAg=BmQyaIX&&Ro%3^6o?BK&mSNYLt`-\\5L7t+Punp\!w[u7<~5a_a+T/*_Dh?qf!uLAR3wLR:n9}]U\]ZRca;PK)y,!	;q'JjBlG|Uc>
t1m1('x!16S#80BdKSy/qmr1G:[K7>37C3sgKQ _ds6~'OS@;8/Z[ Ew;@1q> W&Js2xk?%jA=LO]/	yk&,clC|g7YSCv	6B_hUL+2m2cqI+B7TWa>J4.Cl}JpQiNg{"xVZD	Cqz`!tYr7@%$C4v-[4)_+G+LsPpQ'bz@(nk-!"kqltR3_N_d3zc]R)
KpJvIH#Vn(YZ`S18;x:8YIY:8fH|n"m5P{/X;dE#@>(\uOEOv5&N;Z!e&`;y,g
~_uth:2^}w7n+@ 3Wn?NK1xpZ0tZ|$w/@amJQ29uA<GX#.=Z7)C	XU]Cx4)X6|KiZt*}k@\I9+v*VDy3r{)]$t>*Y-y-T!P0)E}77M{{C7bR:iK9xsYd6k7wH#]K;dIhOHf1Qbb5~YwqS.d7u@8=NUEXv^Lo#6T:3sFlUicXeKE)iAG=P3baI4L_U:.CuMwpCM(cLN@,~u?"0Ib6)cW-w
(e4rj/I^LBZ\sw7_}Rz504Nv&(NZ*Uk[
P]re<L$:l{WJ4!J?Wm?dU6G~kG`/_\g
}NR#M>J)-oQr~^o?``oG_'8W@VHWgRwIH(8i{\zb's:Y2}JdC6Q/bP/TZ])V,,W\O)My)q2"g)0Sd7)&y&/uJAizG s@Qyp<.7{gYVSo5,^#d|mJ @8M[!08QrD`5
.xjcK{Uj[3Ct 0J|zEay,u7T.mG5A:CIHpI{9rfI(~0(ME><u*4=y}4B9!%<M88)/Fy3iOTEslApV)-g[gh'\Rv3{1x4]6pXduHK<h!ezU=T-&0l-MOqg[mCx-%^X"z<OGk1r:d:~k8@+50g1QgBbT$t6mirnqZZD	{c2o!oISutp'iG|x)vWTz\@:Zy'\5..YQn4rh4$(;$Lv;)b?GrPD0%KtB^XX:\mM MLZ-I#7<}LH]afBX/lV')Zv`j:&>*w)q?OS:Qcx eV'-2XM ex@<wT$HI+\O%Cifamp:PzGC$.bHw\@F<nRac9ec#}>uDTQ=PjQSR>V3`usKE_%Yp&H^iB<cVw	pIFXESH :IH5\(,$EF@%5O?TvtO,<BRbUA9jKbJ~NGT5~,-R'&3r~}l;C1N\R0}[_,UOVo[Fyuj-k{~T&aSxF/P&$a|j+O'u0YJ`mj,vGk[k;fEH6V.'67`%?2.@PN]/n.>i%*km+&oNsSZ8!Vbc#!m"qV6(rUofSx=*9'5gk!p5ws@Cf3.BxLIjq[hxx9&!hB~PraH0Y=Bti9^'FW:@v;Ve	I9FmeXC2|JNA@M#hdM4CE+,k7F
wjz92TF<kG#JR:e>i	58>L'N0pXJ^xq-X01s%TB\Vmw&x]WoHwOf<v:uYq3,Hi'N_e W	pRyTI&?Ioiry)kIw@qjmiSkgJe{?}5|}(l02Nw>0TUzF9M:G*+<R4chA`B72Ob~kcHfRmJ3q2VkfwasYD@=BCzV[,:l/GIc{(CUsVOFEuX&l,ERJ:j/?}q^O#f{0!Qh)h_3;klA#D@U#s;toXo^,Bjl}Tkmk(;x3Yp+E*	6:,qOkI,7_?f(a#s'4BNnyP)ws=O$!r45ls%BO'f1m?BF~SB6?[&aJ *'`PevwrijX1`~`weS<TF"S*WnG]r}+/VDBu1fF>]ja=K:l\#7l{+HEuqD^2-xK",Z#,l
f\BAV}AK5$;QIVe"<EfV8g~M
9JM\emUJz}469)ZXX\C-SX8&T7Aqpje1PjZXQYv=#%.h`4/fkEUtcu26|Zm+DB*`Hon\_0$RaX:6`C-25G1[zp2A)KSTYQCwgsaQRFhv,}?;Z'ql*|2u!nungQP!~|Im}rOhBq+f5#:
nWt<!\E[]?4s;!E8ENEt2F.Q>r(pw"_	2blOpyGg->5j$y-AKI	#)UylfA'9/wFJf'1<Zf	2<QQmRR|i8Uv;^2`>{(Ws_&T[NdQ#E7I[cP|"e|[6~j[UW9bf	nKMVj{;PZqTk]Y!'le:&cY^")pa7voY/7^Z3k_r	);0S6ji#$6V`6M/&t]7|t
u|c:4/d{Kd&,olcY.hQjCsy3L[O=3vt.*2zkEs0}h4srP	HL@RhP6\F4~F$>ZQ`Dv)-A:kzp5LndL$c}LEZhXJ4P7k:0h30`h4	eyp=}1O\fQ'Q-4ODJ,l^0O Q"hv`}E.;`pE\6tqMxgMZ{_bnicdCZl)5vRMO 2$u"@Ol8GOH#dz\QU<	f|){;r:'|92+K<7\ 5PfQC)myDD59`/!g9BU)yezfO~z` _c.Rhc>n`QSRl@Z_:z*1LUMDB5>9]tr|$>^Z)Q>7(4_Cr(@#Y5cp)3{H%MaE1v/YInB3B[ByEJfK'!\lKW-5::z$H
A|-2.Q?x?ypmazZ>\?3o7~'&:*J'))zT@2Lbxm6mC<)95!8}blWQmB2{K-(qV_o#=*CI1ruo>W{Ru+
WuWSav|qm%9wD)zXn&x <:ZsDO1e+%"">w\za1mY9VMR+m=>cz_|p/]hBb)CDi5RZD;:gTn?hoyu*es2-#C`wY(]zJy!-^}=q[-qV;S:_7!C[6\(d(=SL]h_KMQqK
mWe9K5zZD'pDo'#z@Bp)_' c
S%
,][,('mFE:KM
4tlH7[M;3bC=\A(T028/]LW9GRM"'=0<+1{47Ig@5A/nt"03k4#ep(kngt1O(X>]$R$0pJqj`4gQs0)B4u-ADsK{K7{z;Bvui(jB?K19A63	]t(ft0e7`[LF+t.uG[C/2V4O,Iq>4a68^tEKj?<Xr|f;XMc
SH*mYvDW-8gK7Xe#Q.XA1]6W
7M<"ySn:FK:kT(zdKv'8/6iUMLWFAz+("Jgji|BduSo4q"\;_,nNd)M&S<CH4-?w-Za3q6Q\orq]V,I=0s,}9)=fvR>[huFz6vw	FI$UnZp"])V1!{:4P XVq|
"gy,Z)wN^Wq#IJ`=\|-w";eI_4oVhV1w,C'2aFSMbJx}%}xj'#DD9t*SCptGA8K4BTn}	>"J-b2o;&n)gYDdU(e;;5jMH=5a~/Zdj\01g3LAtGhK`r>y.[#[rql{]K`hl8))48@woz'3LIvi/$S=\`FS^4=XMrra$\aBDefMrY&8`,~#nxn}h?T_[Sh`[NZ"Y&"V"M {OmUfa6t"6j"rL?AT>gnY?X}Bg9s&$`t#+<
Knr#c$#D;a08#ZcIBO5^0tS&a/ZVgt
^dy.;7wbXF(w%FEng\5shrG17\]S>?bDczUrv$6T"i=E<@ek?22KI7pSxP]{L>$Z}@>'_VqRza_VW2VVM3$8[-\-k7V"j.F5X~@/UDNy,p}OeMxiBY[sUPr1]GDiQmU~,{70tJ(be#L}Zd7$lx\urFG1.|G!O~vf*
fh(S'NijZ<B`y/Yj}Q^^USS;x{x$TH.M?o9t51Xj;G1{ nf[WC`iR}+"FS)S,4-/$n6<%S6':KX)vshQ"|3iR*7HfQ;z7n?~"hD\KY)pDI~q5=Sg4:N *tl]4+S!	zyC(e#kp,z08FX	O0$0l7;{;sxo`MG];		 /j`#1R/K
hUz*?u$/!YS8V&>F9]#LBj\^F\:uq!x~+cwqZd7k$1Gx;j#8>nBTCfF_jAHpB|SCHSpznXO+A*/]*.3%!kFXE SZhm\8DOwB0j	ITa]v-<`Zcu$n[W2/qv1>&`;k=hr'RrA6XXeY;(eXCz0)OXXbH> "\qP)i4|'&AtnO&(`:Ntl;Ly!f"&sqA)Y`QkR_frBRoMz_J?cp:d%jT$x{%L/FzfEqx=T-`$..pQx@S]q o"^ry	(|R4DnEM>MtZ;m<-:}gE=hL='\XgrB$mnWf5D}hD8<eJ[:`0kh&
4H.?EA92<VQ[!i u(h)~$Rhco~fQnaKy;2Tr`mPUb4"cwX-C(Z=ujf {".+`7hR)B$\Jgf2hH.v!rm;tq{^kf'yMM]{X1lx?#)M04\4+o_2:K!bi{&]Hqm$WJ{=EeEm3k85(k$i9kc>	8p;~
L,+ViW5!Nmv&pj	AG [/AOZ&FaNDy_?o!!Ge"@~T$q:]v"Z1"DR!eDg(M1KQKu6/799+W;V=%DX~o07=,*eQn	`Xewg>*=!;j/*\FX|{}m)	F{Z|)^':?Bs	?>s_}I#JbN&|KOC>F8*\<oJ; d,$X`o5pl2,V8>rnuW9FhBz?j]<=,&1/[~[}3iw	[0Jd1"+H;$BdL}N`uZBmV0]s+hP~w1G0!JEs.Xg'[~{r(?mz\&|teu#n]WaTXY5yt\8`V8N(V0JVPuMZ>b6yYEcB9t/f%b).?xG=.>:)@|OGaV}^vI?"nra	@`kfzH-/.V_YO%Yq:1,~?(hpSTS'1j/,cY<DgIUe2H Y8v>*(O V1Xd~xxTm'V1WeAd<61v!F(WD%i}	?2u7ku(06Uws8_
|+y^C<IpQyAAp(L"^P^dennf"r	CGV;q4!W\zjfeq?hC:;-o(,SN3Nl+OCC`_G|+b<tjkTsqw?{g3<;Fp\\e:''zTx!.4T
0|4T(n)Bbk3D}n\INE^bvSe<Roo]9g3^9bAfF,^O?lM:-i~5,`|_'q"pmgS/1\(qzzaqS!dAZ
.c`Q&`wK<26;W#},/V%RaJ.b%u/rvh0tU~36~%(^ZUm8\?Hr@o95Oyi<ttu3o~8k{z|{%sCd6U"#WEmk
-IiG&htC#]#z>O@lS?B2!|*q&vw(q:S\hb}OAKa.t|?}VL]NDYWvCv76 MThf/X-3^O	E3Q\R6?8sKK*_e]%UYj3*K./6:3qO3FrqKEPg,((@jhxEWTGHHLa`JT(latLeN4JHyR3:P2%vlp4n;#V#"?IS={'"+)siK5.\Ql#"s0@iqTV1K19/$ppE}EL!q^uRiM-$h5CczUn[["a!7mDr-Q?-(3)*1HE,G&x9-5BWqry>F+p;JY ZCI!iBY*K{OPacb*5fAf-[ $~F1ueAl>%e6=uY#(T#$_?cj|rKS(="2`E4`,F`y"~|edhOHxRr
{$MWQ30S=v-PqN<wFUlaj+gT	<%$q$`
0@Wf{<HQvO{M~rh02|S2<vQfR=qI2M?"O!Ig!MGC7?|ipC/<<NHj}}+:"s!}lX ig5dC/yLTDP0M
fYEo3L'6H<YH;w-R'3,mGUy0l@d~h|7tJwB%3qpA>_%mG-/Ptsa4Pg8vEAKq(y@(7+~F,8Y0"Gd)GBGq0OXg/1'mQ4oAgqwN<gQuy7^!,FeIT8{FKUm6,={CR{O0lBXYYfTr=k\Rj;,%uZP22{1:T&4A)P%>Vre`mwNP1Es(t%(|T;ki5dw{_Ff@JC<mCqw,P8YmjFjw	teN7he	8wa;D",7 Ing(69$z&72iu5[44>9GnwUS6X3nQGO6ryvO-Do?K5J3*rS"W@jR*~#,Q-`3
1/o@6 	q	z@#/QET<ksd5"I4Wp@ekfMJ>\B`&$g~P H,!&#g)bYu%xt)AFp_vCk1.ygsNaScYNboheVq>VS!'K7fc&|ou*mcXqm{TTuP]kT`wU[0\U(0jE@F7~N}T&8w!\5P"i&F2eX.v:=dUB}JF8rfcyh8
YIPaBITQL<Z_%urqUvH@aABt1@Hr`tnk*lUbk#6(&|SBa>@sPpfU ag0k`a)a[L6)M}3]_E*%7)9&8QY
Lv_fxZmL:+gIcFxe"tDP<Ba.*O!P'$_;\r0
.@IK{w*hSR'q;Uc6Tj-%B9R%DcgNmq?s^Wj.6Cw @z&78|XL<G
C:CAF`+	AbW-Yhdf\nMD04~g/m^ f6	@O5wN3}0U!:k. q(	]T3 aNWh\I\5](|<,O3 E+tk	Th(M6Ejs%SM,d.z9L(wyP)-vS\[I9aZFexBLv/(fi[kgJUhlx)Bl2Je){#g9,K:AM[y{zK9*<kC'9XCF<>SJ
y{
BLZ,S_#S	@w-tFUJC9fs44->RED,R%OOq`|%n( n9y'S>QimCy,@.wX~wvUr[b/P,}032-0\!oBy2,SXHxt6624y)yAd#Z![y'{wfH>Jf*M<vj7*<~x\R*i[O-"$Ez|fS6KMqEs!ZoWA)O]Pt,|<I!&{\A*q\PWJK@$Ar9C>\['3OSvx>uu99IA{&az(OXZsE0Y\%@R5b^{$L(lyny#0$\|1?d~3NQS2[ztNn27W|\+'?5]
 <:N;LC^[3R__G^M"Qq#(Cs
2=FZ|BSrw+qW|`}
S/Wv|/S(!!(}}3+-b	sO{fV-FXg[FaVEVv%G}7*=lHPJb$4k!y^#qpoV.1eft _]f#$S6&}M/j+-M(]pUg^:)_U]0nPvI+ap!?{Mb][57	ScI Pdw%R sk*yhg+88#l@%^aiFb	?|lPop(`!Y5nYFVQx#pRv|m=%njV3	$TNG<XL|Qy,1O?kn,AnTZ7
nTb^jhqJ&:9?$7L8<;
oY0oz"y^%a/LWd1/0wX38F}:	zw+C(Tkd[/P0SXv?MtI5(??(ea	G}Waj4o }%OJ"D^`V&p6~I _NlkAh`a|Uh4x7AQ+)r8P&W 0Tp;M<8++|wH64SLIt<Lf)	\5p;z0^^>mDP5O(zL])9qkD>6T6tdrFHpy=-xixj2\y?/r#z
Ed$>7EaUI/9Tm;2}
r2N&:"LHTUNy+$3\uREC
Pxh#h1+Ym<5P]n^+R3jQ_9V@C\L AE(Wq+P-$Od^*~W_:5 d(f8[Qj3U:`wB4I"UpR/1Q<W\6G#ngjYkQhAK1^F{1&	}K{Wzy/G}#<A|AcBLlw\Y$\_&(~-oRyG*s\e+=?X]|;b0hYxbm&[!O@e{2Flsz#,}KL\tz{ZM)Jf71Eo1D*w?xSFMNVSjYk]X,,Z)&p?sq%MDy;b$7S&#.?nrh>uF<A"u!	/R|0R
H|c1^ 'v9u!5|*:A4_4Fqj|,@/}1yhI,v(DOP!^J99S#@hDOZZsD@JW36m?+o:Jm4q5|9dbEdZf2j'dwLz$$9EH#bVo!g+6{gPCc>gF@-G"e>qRLR3/W72;g.!(^R>GT%~Bg%\Z)Yw`	`&\~q'x/d[!h&\p2gTlZa
#Rr]|Yi+* YE<\oZ{S[`C}c4f+;g>eB.~8'P*DSW}cUSDiL"Oy@
yP'M	'a7Lv8]qd896\CGgBMn~yDoxMh^3fv@'t0J`GuE"s-c!%IKmpLQ1qn#b6H(1"^/9Cp#]Nkwbt]RI>]u?;ZFh@)$`P'g|ktZ);(`Q[y]-l_G`mh>Jg+[]r/y${F!?~V3@@T ^
pfj_It+ihkA?-,86GPYOQ~+YU%g1r_
b^*	s*7
A*Ka+=QWT
p;n{;ubw3%F	+{O],Rh+f?5)F8R<ReT.AzfkXG;G78%+rhjV0rxMyrSg~Z*j>qjXf\%iQw7X.Bkf[ACle._	O/{*q!}	WN$2]u/g
:1[YtBC[:=W"E+{z|}Jn1.n.!WB=eq!(9ugYQdy%[O~u
T['HGUJ6Q9BEcUXvI"S
BeYY' z
.6b$G8/.!oQ]ttw_*?oipwo>	1GZei6NmGLc5Z%Yz!(xj&Q1>8ZU+W <45?M|P4Me\-Ms;6_<zX&6-TQX>/mg6<VrGdg]mQ(nno";-fQ=%~oifm4Uap^^#h*O]n1W_8S_pLsI~T`TAiiu	hO5>01.ZBl|)Yn_SWX<bQDG Tkfnq;>f!Y_(cDm;[c)Pd|HO+xy:N36MnK*'@VC+FB9z5J}|5?.$ObM{2.S),#cqIna1)fj6.^D#W\!6W4^'vg9Pxu/m.tGoBd6uZq#!80`c2]nPtW&(klJ%M!bK
JUq9-qw3|=+;9oTr;;D_J$3aI`GOm(^i+<7DE+[4SlLi|52E	9^xh|*tHEgM*5</qiRIfHy`{m}%F%|T0Kxuo
;Cm1VakqM!'ZNR;4]_nAC41pII`-|>yWXCRN;K=$+lg(I507#c0.v[.E[Cu$nQ1v^Mmkl*
BL4Q
_W($t5W'&?QCS3A4%;8 ->lb:*43@Bm:>sy%d4qw0'*XA3Avx~}@P>fdT">:f t%)}n_\QF+\IR!WOzK!9c}u`IPseE"nP> 2I7.)\D@KE|V#dyAV,jT2oBQF<4u[!fB~n.yi]f
(TTS"hH'fFXwl)uK(5*8&/"$R2gh"#Ey#$|$`*kf\5y_`(nT];HmjKGE1k!)aHe8J_zls5~8@
Rb!]yCyzgCmpweLDx*_6Kxk~4j\wc>a^Y]j%b$EdN9?_Lkx
Q0LAp3nd;FToA6	*@ls&g#I6fD}P&Yn5J4G4{X_pl#F\!f'X?bok-*N*DiFm?<\J{!c}+wUsE[PEXv@crg`l-Z_=|*R\fuj~@r0s3S  ;//F<9
j{i"}8FEs>+~(U976NfCo=-#,=p}TZydK5'{C($9m;#X$:@)d3MM[yW#l>_>0	N<wZYIKcD!eU<0	"ecFn
|)-6ZOO$?M{>s0ox3v9;1>27yV))'});T=	~T@]4ut?89	V^Y2gogEhate	}"3Enru!a29T,Jr+p72+0p@-<|dbxdmIXo=I&WT?.#wk~ 2]R7~=x-PDC^EhX)~3#&(*U |VsW7&diAcT.Q1aGR:l@(<`&SMa$cw&pyrm@+/B4ntdfZ8,.yCU"R/54:r8JWGVm
K,X@^|{E: VP"&~,:q&+$zABXjq]M^~^udDI?TC]e)Uxx
U/ywfMw{C{ww}:?H%IbXkm1C]X$	!d@xc)R\@!HOO:&t042aiM|?2:}I+utRyJ-IYWhkL+Z&O&+)O1cdPu@yvI33s-(mxX#uv4lsa-&'Jnc*d2k-`	ot(}dY>zaAJB?nr#(yPMeUfnF?k">.FHO[~,)1R|giwx[*mB'u*8aLj{:cu,=^Ub[x@7!FBkbOh?x\J QVap#<pH^o]n-0ys7[sCOlE<~sV.2@4wQ*E{z
;K(&~Vs;Nd}|"8|7X6a7,^>\euRY2$v
vDRIl
'p^5&;@D{(r$9?{o{G7X]M,s5 ,S6nKJggUl-{dD7tO}~\&"1_fq,}oDo9@FF$9Hlt""e=Z-&GmgBk<
bgus*ycytM@e[]gTBbkq;dt|SF/a3|_lB'-45{0^Ewm@nmDrTvslg l%]V6Q4B5ahWv(uqmnZ\)?(D2<mus)tE}TKNj421 jnv~`O6*0<)G11ELAmQ@f5iqr7;6;\rbr@tqNPZFTI73X01' ; IuU>Q_nc5!z</i;ZG@6;{}<5_<{Vmy]G4c$?/d/bfPfH3qn}a{>.z~UmK@E0W0i*!7h.5qO6>IR=UABzPYm
h,'`|qI 7]i3]Yd'6</,xo.6~c&J9TNsg/sbecc4";% zh	H~_-	*\ZdwoXpc7itr	zSI\3j8'Bf$+T|qg)b)"B?OEQqyq"{\%u%l$of3E{;s:_l}p5G\t("ja(9V!u2~#[jXTF0@)C>Ic``Vk'd7Lv|*<x--0*mDBd@.%v#.LM?8o9Y)Ie.}Km\ls|tB <h]W%v>/Hgda@YgN[)*q{<#f~/IA!/fwr,yh1L)qUh5!*q8qGW3K%~P)A"SH|WP;E,H(X!MOeaW6<zU>o\.@%HY*Gf@!keH5iT#'oF?AT'e.E`qDMxpG40;G]f:ibdb~_$794<C4YK<]q<L`u#XA]5[zEq6Uv$qg5D?bY::&25<7tb*Y>^*e-EN)~)^]d&33L`{`;uhMBl?ah
my.Zzg?p^lz[Xc-C%J,CE,DhLw1];>30x)|;[;ED_!v3f+B9+t@$2a>Uj}{(RcphS:0<n!PK~M]	]IT02]k,G,llGjFKs-rXjck@\g)(uo<GY)nm^U~My~ce3Rf.\7nu2{F_{'1'M!mX[{(U' }q7&"+'
c(WoR>#Sh_t$Z*nU2.aKNoI}	;JSH<6zNAE^iKXD"qU%ATvM\\AtR%@ y:
L#i`'?Yc'|q[N!].X3mU?6xSP~eD"|RY\R1N^2XUNiOM?&1ztvQ5G=}/0:w|\AvL"&YJ=>BfyRP<.O1S=HbCt*\o7db"49;GLZ.\ZHS|>dd'!~eZZog)|l'dYU*n3[BVM1^H-q,JrD$I?2w9Eu4M2wO=*i507x+}\5!{FVw!r|poM].}sJ?s$[qS	dpnz""/1H8KwsH)+Me9[&4w-L	e;e9[l<Q)BetTi>QRcei"/JZzvqAQ9v).	tbXLaP>[MLDa{0;S'L\@{DAp+vSvX&ai,|tb2ea{s~i;8bQ.[ot6G2Xk&:3R|e7CEf/2"NTIL8]xj,GfC+Jdasa.~&@OTLh^)z'zA'6s(NAe4OXE~}M*7WN:%ep^OsUuUVq;X[`FYH{h(qjsr6[bw1uR@QnI'yiRyO#G=d8	wprvp2LD%
v*E:k.8R>[F 2pXSw{9jSb?D5ySrv6n}o*eH"j#7<\^8.d 2~U"i*l|.Yjvc{yVE{#>m`HR|rzZqxxvr MX5|n=lpg8'0vLdl)zoD|r]an0IZU8v$J>p42D{7PP]({j&nYnr9m)2']%}Hhk}+U:.]@|zl[
 J*,3rx}j:k<-T@o	SHK.933R5<79%eti[$#Xjq
?	#Z|wuuY; 6*k$!"w[N0U4d[K.>WKEET;j*b
NT%}rn^ARqRe)zP[K3[vV"**>D(t!:%	Abx_f#7qHP@	Ooh4SC#3A
A(O{gczrX	F!_h'cO{lq;#WTD`<E\/6N]$[u:ae~/C"j1,XsVkaKZvvATuan[r|$n.I?@kOXlpu[o?(f/tqiYJDs2mE52S({0%pK6]>+LPO+)NfVPv4JUIv"\:MA?"Qc[}!u>SGHcz>K,&(!=7&7Mf~']G!CY%!prQKNXEXw7RCURX
P1q@>z@a_t~*;e-~xw@Ly(k[h2/7u5\m<9N`N7rE"oYXY{LXQXb?cl%Q#8s!.y$?v)j?5}}8|F(WXO:RN.+;eE8}z;Nw*/!shA9C!,SW%lGCPu`yEh0int#zBX}9{NImD2{N2}3'JB@.: F]YMvVh/R"g?|0lp
|7RR~	FKO_oR)Ta
d}*?LEP0G9SOhEb5mAU|m|fUU<H#LwCdi5qO%sOKgh=RI/	Gf5PddbRcr	3z.8( |}u$`U5eE0;ZJr%(42+(@=t_LC|a}.]2b[ D^QI;9oXzeD/H3)$3:
&Ga_|K-)RJ+t;/e&7aL@r1wa1<d9&'Q`jMO6u9iDQU33)[I \Z?Md3FWbpLV.w/Nc%sbi!AMr;0LXN.Nx[D	=GGWbYvg0p>kRXUti8eq/x=OfSHS3	577mg^j;Q
F{J&uwr:f$p0eY0"^A{mqRW6h1W^K?3eV~PA}l%4Qc;Q[/VouyraUQJ^9]b'yJmFoq`xeKZoJD;@:'|a=hX?|mj\/g4.}P Z|J?e1/@6S^*T	=j<Q,R\Lk`8(J*!J#cipv|CYBc!./GimcJ7bso.gR>yWHnt(O=?+"*CSI-b_:
d#C>G{\tRpA0"{d'	S"&j$`;'kv!q4x+/ae8KI?\{ikW_T`Z48.Fw<$p}*Le?,+:23OxgYN*
hT]P qhE#c3$GTnD8~fJl0FDtjY\3Qy.2[5cpZPesT41,p@:iQgjMbQR3t`a_!wNnq.)sFPKmnGv:cOH3El/g:Q#K} p)B(TN]e,'lw]	Bn*L}~OEUmi/c>A.F8bWJW/{_N]Nh999t	@|"Iwl/RS|}\B$NS5VqkWS5}"[3T6V($RLgh9d2Yf~g]p}w$hqmtk9G,?;Q'-#xDxHLfw?cDI2WqW=gonRb+muHTm'7.\f|x&~KhmsmOqy@<NEf5o`xrl1<3A;(\ET65B&K~<v_JRlr^CX,H%O+-IO[3C{JZbR#/`h)GAZ
A97v#Z#2@Fsj6^b	)oz-TKqa(/3mq2R/A=V&KO~XX>$MG)h01? 7t:F>s[Xy.@|g[)4MXNv|:R<uSinTb$m^5/TG/TaR/mh}\;,G`W%O%f;Q6Fpo=`S"QJlU~}Mcg6]36p5iq]3%(,w_hFgT1ixq"SVNsY`BHyg^DZ@b	,\eN4pyM~qAU}bWcggL]AP>oU+Zc	Qn+4
7?/|zV
mi?<x5&.Jw3_a1<IU8MG}Pk~C_X"a]9,Z*uH`MImt*&.*ARF-u_;_Vry[<wTbmJ_dx:s@7)<IYM4Y,|IQ1y+"E-6#sQm}JS
=oE$!M#7v6#')@N?	qPDx6)6IrR#honjHql7Oy|W<4c!4^X4yDSw
W%&qJMDA[zTA0_+Ph:7/kL}v@kGA/ig"C[~!bW{\W/,We2yMj?^7cE#lNuM}hF<aN\|/N]Dfc|}cM/b*{%/9B54YmQw_/na&)J*orYyoPq77P481
cO1S&vn8c#X)N[l2E-Ok&2)PEf7'D+"xd?9\ WbGDap6308K_(M>xO?@mg`/#2fb	J"FW^RVkKG9ry'3X'cGK,ZJ0<3uEr"rhmw^3Map.|`H3c	kW)1j(BuJBk,SGUpDF%##-%Iet}w$>P$xuXV^v*W7ADn4*W^;_jSaA+aTv5}^K/#$I20V1]*X,DiI#ULRjx/s?T}LIu86,I!@t8yA4=s!LD\yYWMEs&<[MU@^?}c:s	PAaN?JZ[-Oo)WR<^l54Rk!)F3`n]g32P5h	f,Q{Vw&fTK^["p9UC+yT@#Nu.j718NeAX GY\QSe^[$@T9~P3:dIFq^,u\{	2M?qA+@e1"<brE,,l2ut'jd=P?0S454}	%,O^Q?yh;-^>9I%qd.yJo5$5*7' Od<`Qx5zd6C^VV5PQ1bGK%=wFx_t,	"Pzk6nF/m-{^_E@9UWQl/
\4]rVrAR>G4:G}AJela{yEN7C}97HKZ]@b {&B5_tp.%}ae4DsV}UmOuEf!'[S!<iti^|%5NR3Te#;x-W-W}Tf$cd
H_4hX})rrk\`k>3-9(GFI!i/BIm3DYF{+n2_\4,(\d0BB\9.J+a	sDDybi[KJ-uxb['D"9|l\Lh#JTi@[	|c|hR(JJY/2 I<@`GD"	)=x-PS2E5/ZdJ:~YuHQ$HUrXSwvE'CDWyr:WPiy5T/bwmdl7d1j(dHpRkn$hv85=bHz|)]ELNcK\X<5w9dZ\I{C*4N34yDk:LmqyL@rOFw`&eInJB@PC|"tqfG[Dwj3`LJ
-F{Gg[f'?Pbi5$j2bAX3fAc6!?V	W_#|)'v;(/W:$cAl6g_pf-hCj$fJ.Q*Foo{q	Cpxj3vG%70)<	"DP4dsHK'w:4Wxt6+W3))^w(he8IF?-\(STfY5m uGV,4!W7*')!*6*i%?m*rct@RrW	gsEUHI`F^-1_O3=,|
Kw
\kO3	=LZxEX/q75}L_vmvT9L'WGuaW)V<pp _
<,vUL-ddg4]]z8TKb#Ba;E4~/E(}7ERMCLM3:;>+6(I3xWWRH2vei3o+g&QI,ljiQu,D9pLCuju8W(Xt`6to8GEQ~M9.;8XQkb;8VN(:)'2"*'Z8r&M@C=]4_WH@Qa@\2a7'Ws-NL7P`<XWmU+0Z;x@l0GoeKfC`2-f/!{TMd?GO$`	j1tI]ph2d^E$4Z[CALCVkO96/|ow0GWvYaxqbqV<qV`h;[6 EA(? VB(h#9!>@C|AonK!-1{2l08Jis@"L3lWL&J/io=@uXV,Pw\k6(}r'.CTIWBvU!?Zf/,KfscIX
lDYr,</(^: ICLU`$zl,\#bRh_kMORMx2JT1mlO
(>{HD
g*J>J[@L1<fRRnR/{)@#3}\<1k5_G(/a}&M0\&sw74t`fYkL08t5h#>r5@[;60$]C~lKjerPrs`qRfM;	"LoM?=$4muCA~sBPTeFjMSUhf&JM1Z=fuh<.`~/.+ET((p;9.hEcXcL-&HRv(>E(YxWsT#d|*ss^"[`px:Td[0SIc
(yNXU_XeIkh5Z_wZ7KX"*d=K0<>OBrE 6j:dH7nl]oc5*uHFg!w=0/S7}#oE
C!rcF87EHHNj9K8Q[C:<,9l/h:/l< RsE1-?INR~9n[P=>u7rvVEa^gjmKHkg[@YBeIlW0+dDHk7wL6q(?<CGp<TW	l+ju(BFX(e4`vJj8bf02)Vu%dF	tPhwr"gJC`fi&Zo%|WO2v<[*iCo"g:![;Ma,SSN-g}M}
2-NEKQ[*W]|cUm<R%[D?Q^%?_jYZS	fXu"^R0F||tep5K|RH>XUj*6s>PowFyb7D	Zv7YtN=[\lT}'D+lNlqY
oiKZ"n7zJcH
i(g.u\R6\E){.GXnr6OfkDkj&61W.H"_t?b8zB>T[yM ;zIQT!mTg1pEMLL=QXSgn!E4ULCpFX$2-:(NR[~6rgJthN=uE%|}1GQp2,73vX.q,O|Wu[F4-q#:|aM674P&M5obTG(&s@5<v#N<"t8n[V#q7IxY	3p
_ZCo6(hHhO++ tO[f&&Fs+0abD0??+r.a24y.%jdh.riBtTcMISaO?PKSn,DK[KF~gUL"IvAI}Ouj_8=]>p*1OyI-e&l9AL]^!g!;0P7UjWJ92Wox MG.B[t_9Nk}9GmsCT~Mc^7XGU+Ivi&Ct/O9DQpR=C	cf^JH|Cd3D5KTf!$]7&i"(:v[?9$=IUGKJAKE==`BepG4$nOGOa!Ozhp83Mq-3|ujc~dUvqW	A<X>ep7a
GUI9]!e$
&7uD:f6e/=B"|$.V{i~~Ycx 9TNa-A!CLl]uY{<{ZD+j')/C-HJ+c8[~tP>}Sfo,>".?=}Qx<w9bDohve^S5\PI1pF8G\nbi%/cNAJ/WGH-[P?8;$,j$*YZ~&DN[zy)u&ng[i&%F-,ZN.Pi	?C<S	w,@bi+C[YTz4tLjClzQq0*[X(11v{lJqAxO":FR*QA7qXAz!QWvNKvN	_,+0WKDQkN^{-xT@W)hlJgU>soq}3K$RlJ~iN4l!RiZ0mP,u=$?BqVoNezi7+YF<YD=U;*3}1 v'Vt:?,/|;:3Wh=}Prp>`@8+~{II`2c&T:%[tVK#]m>agYhA3<B7t37JEc4wJc<iUnK*	iQUrmi.m?VX{Rd.+:hz^30KS* \g7E Cv+1
x(jteJ\\Pv}+3u227^yr+lG3MVaScG'FfR\5z27g4]RF4m|y3{UzH
2%l#lno% AItstc#1&9k&xq&:	{6&%9SxcSjFzuj	duvTpJZG'o/hE	i`)v\c2q{LH!P}jO-EfnO@1L\bY\W-[Z/*!G`C>1^s*+.6|@<f:|oggFN_i$RWJm@)2(9^Z,_Nsq./*CPL~N^<MEVBzYzbuBx4F?g{A#bv{$71Oq[3!!m^mp6oenhNF.v[(6ha77fdzHa_dXTBBg::1RP]J.+r*#{*B2bnz<mP
!IE%\C'cphsS!ER7$;!j%["^*.ev`5U9Np*)\i uSFK_`@e^g}zVC4T}1|rzj"CBOK-s(<"
XW@81C2@6@	ny!0jv06~\x{}3/n1;`CrXZdW)a&)>DzXcfk%E(svz1H58[<_xk6_}ivNJm:$	1Spq	PnkVoy2o_UP&eLw'b?Qy(JO@du)r
+6F."|_h!WR":n~A3	tg/8p+'B} 4M{{UH[Xp?I%28,<wEb6-D:5!3]hi2F?L#XoVv(`o4NUEHJuRIbf)Y8,%&pd`6JxD5Lo9]=mXp-NYOFxK'	f"|8!l*bt2Vk	@Q6=IcMC]iU~1tnZNMTko"3[-9u)Qjg5U>]i?aMk'9VecV>*Zy(86#DH:*O[d*m\([Nc7KDdMu\2{}ab>E^v?wLm'0Bpo$Sy!_yLd{hL^p9gR?|tZC3E&I9yJD03FZsZu;jy}^,iT-==OWD$rrkL#=NL%W`?2OC.IC)2W+K}i!N/+>2(x-K{0,=e,E-y7~=E	:@%v+%tX]fFI[!P[ 2t_bk^t$]Am5./P
nEz$U/<9qb#^gTS0gg&|[:X2uXs&WC0INY{&'q,U/|Vmpcj4pOP4qElC~)o!k1.?N6)zQ3H+1jj
4/@"D:4?2q+	DWo"7c<?a"mHa`Y-z!T>EO/avP?	(MUoR54A9Y3DIBY~pdJbz*Fn-JE43]7m{+!oJ9wi5yK`Z<oK5~9SYg0%bM[jU(D$h|E_D{63ev4J4+8TZv=0HG V[D9KA-W(]Ur(p74{wdvt
Zgm?nF_mad,"f7a3RKGfbDGoV0U=]eG3YI1`#,#Q-lAucKLMT<FOMn9Ag)58f9'<h''H&]NC=&-TZU?-Z)U)l}@3U:_7dYg3<:VN(,R*'eFL!YVtjJ(`3#jRdad3Sd=yXeSG'sTZ6r+3z{$,P?iU*:ie:UYG6lctB#[Xahj<H"ge%Ae&C(8Kih
g+XHDQ.sL~D=QN13]ovb_;zkM+QKGyC]?!H,.v,uzU!:zx7_P9|V3O6&Y+`:j44
e|	G<srU,W6.KkE(<%<x_?y4V_l{#>V_Ob<*Ms6	L2IDQGbu8}Yy>m[qk9gL*v~'pHqe9NH]zV~Myb=VJi(%"`3BXhq1dqQCI`tltrOhs}AEWXw9P7GJ#a|r(89D2\@+IVTc>VBr2s%k'i)<bX/=|?f[n ?OmXz?B?z@4Wp\1D/`ld2t>K~$fh=}5Yrr])uE.Dn~AKF:z)D0:>woc-MohPNRm(C[S%vv5|gI_pon_=O&XH_Nxy"pP9~|d|Ri6iN?5keJKjRQD;GhDoSOq5,4*Q_B>l#fX*)?'O7XGA8N;W{ko&.>N[O/F
saT}o-CBH5&@EAG_	TMd$me$IN]Au1+r)8J\)h^<Ql MAG?1qzx,o>Q\~]H?B<pB!g}T1H` .{b\Kem}&NjW7/1QW'|6"`rbL}nAL;H9C&VwH[m&xM-m "{3DeX*6q
7Mjsnv?,"	IP[|IR>l6k" 
t50|2aiK\#FdEDQvinp1qGm% R%n$O6=r'tskYL5+0MDP>fqVDw+hFy[qXxGsa\s@$i\KmO_+,_J(A/$]{q5OHUG:mT6dUMky}Yn"4	v}1S'e:PkWT$+!>mT^W1bT(SEZ#N3$>'?DAaR{u>s_-]D]mT&uxtW>&1Wo|qBhUAc;cq{-Gr{{YN(-k}K?z5*L87QfRDp6vgP"[w?Hu]L({$jZ+|,l;rm<v(5H8w7Veco&e9q2.p]nCu	p2+ldM?K'n=un}$	{6?=-4KL?$SUohQW30O{Sf:. "C'Ocyv]yD3Tb`)kc(nKuK;9m1rcC$M@Y5mp9	>O1,c8S_fS+ 5BS;hapez3k@!68gAS3*Abu4'/DZ2q<a*kW;yb2m&2D,'[3Ryj+efX :]/&QoB[)V3XUW<9r3.4:4Ym[K]P6*w
	.sh{1zW[".V)i[qEiAU~`$=u=x$9(-)yD\<c7qXFM_z328v(eq`x+ jO=tr	vCj76n}~!RjbK8X%-jip;{ V_P/)kX6Ax+	ASAThiCoK:pM4DL=N-KUZmt%gEw;} NSY]hL}z IQY$2PiMflpY\>J'-4VmD@X9YkhvXWai`3HDp'_805I6Ja_8M/inrmgT\*zbP$	/D,)aeX
f23"=F.ehMXnNT9|:\*714\Z^;Svwi'*,Q;3hcJj>}(,!l/
5WBGJ*NZZhgxac	+@hXnu-qB:/cAzUAFjjePczi	i:@2m]"U;~h#gtB<gl9Lpq+V6ipKtIZM!Sj4XfjWi\&'6nR8WxqcUp-w1JZzZ
i:3qb?CAr_{e>d|wk2F &	rWsXJ:v1jCJP1y4cC7>&yPA+	EJ'%ist^lZ[cnVS:w9`>Ra5?x)mhLN7ETkoZ'1W+\P#9AjTa`%LNar5a%fTs=SQ	
:THBp;9eeT HIrC!Mx,*zdnyq]mdP\#]!547Axc#{*H`f&v=|L7xPT/&%_4aEB< `TyV"$#`.| 
qumy?]S5!FVM^GHo)
Q4b=_y)w&P"y; 6usn!kDE?b,gXB;LJoDBo?k:LsU;V&Fm@%}_&WSzZK53}#fhTUeg_B'@7`=zN*J1})+DPmpD+_2Nz-LKv>Rcr['\=YY(6Y~>p$+R>,^,Wv_$Yx&"(W Y0}=<j'YhdJT')3?YnzVV59fc&z
}[H<Z(^Z	bthV9>VWvj;ai}0\Dr{TStIp2$Wx6nxxa8,$1Px5`lDUG28rlj>dsrU]gERgxFnZU>EqZwAqH{t~bD$ZQ<9[ogIK{#1N!L@<+:q0=Ei2~3Z|T]iatg_Y`1:UAkqYS['Wk)pG=R9[B9j\buB/?#(3yY u+$	a8Tq+h\BMjgb?aIbv~6'*lG8+\J^:SM}(1`l:NmDc\=M9XxG[&sc5]VL5az\~6J>fJV\8D,kDDOX;x\}wD|imv[pVE}
qGgH5Ni.^Zt%@AR#cLZ>Ty8ma8U%~PF}*>y|JtCk}e/b;UOc:Yw)/'f7hadTE+Zx=XrH}s8flM2Ofb7MZ{4|z{385WVw<9o[(h/Bb(^	*MId~Wa'ys8|}SbHW_(o4'zqXW
TynLc8PwBo)/BBc{d!i!p9ExkpVUE[u(Gppu-0P\Ap\"W[-'gi6*S|38rIsZ.QD`8F;_giJ(TZi)55[x#'*,k=D hM7wD\xZFU&Q9slg16U;<.SO(P7s_KLq	h'BmF[97u~>^)b+jg(#[o(}&/&iAh kRwvJy&y0M8uGB*QTm5Bau!n9F>u<-yEXE"Y}'1Cg!#FskZt/gx[#mp\<eS@?w[DE7[kRX$t;3j/%7Z!5a2#]1Y:EVk*
oi8%mRCb.@obLY8O"]% %4Fq0|%Neq*-&D||w/f02n%lpx0HoQe+QN;xgi.[)W-9r?]eI(Wh*G9h@VZ#W?h"/.C'X(SF%0ZuKD#Ju=T].\L6LPa%uJa&NPLw&0,&_xT'N@SG^0zl^B*me(b45iAFV59h~%N^hxKgV+X-G5:TXK`[Dkg
fz3'w+@^8?pSi>uV;zfa4t5QO54E	O)tBuFb\6RV}b}24t4X:pUC9ur\}s}w5`gxf/GTd7dtkx5+fwUffigO~][V`'f.j8tPbqV,1:dr.!,pA]=c?kW2l4J%$eTJd{~j8&nD$6q+hvJya%Z9[|Wb>}Y;3)-]ZK~8M
Ev/C4SHgQVrp=cK,a<.gt1eqZ%cx%"~0/DR!tHz#6\!1h*	%"44QSC#N.;sARtJTmLl|(YlHh;LcgJK-t4\4w/zuZQKc1bJp_q;4@|^h/Dy<H9T#1{
GWIZ>BFs`hW:mwX9V:+29qzjH~';3d}0H[Mg\;<};$I\`<=x.DlVgj;qC"$tc%orRPM:<shjYN`'qAPsnCQb{>QQc]sB`jsKib|Q\=M.[0q9iJh7,q~Rp,Lr|oKs5@@J5B+x<2	Zjwe/Cq|M^H3/1aTNwKNec]Qz^v};Tgh%9DLT!tp EY{sZcX=j4N/SMK_Enpdh#F`UF4q;=$hErn|-WM,cGr'"![O
	O~
*=)'}n@8a8O73MV	JIgrX9(E!"Y_cNMd+0poqq|ixb.=$XhH=M	c#LGZE6[<G!,g$'=EjbJkUtFW2?N	p]&!mzh' 	WD~v;W:{
#SU{K!B;9niCP	vB_@\u*NGQ'=J+-&g9H!Z@85.r|;E5a66a	.>)ANm}`@^
EsPsW;xo;
2My0"}9RmYpGg>azKG?{q6:sDAcg.XVR4)p7nRbYc6}aAWal=1DUo8hv[DJ]EG751ZC&jo4i:b|1oS=~h2(}s3i1.c
fk4W$dS-'8FBd?O;D)#Q#\xZr|wXA
sKX:f.j\<\]3?%DS<yF!q%OQK{N,MMKZ~cyhRg~By9"zLOr6%{2*o,w`)C@)jx7re_zr%R5coa
J|?'`kCA>Bb=E`N<g7,lS,i,5N)O7OAO*s)ZIY6&0?ciR[ah;oQN!_[uFE_,#YnhBeIU#77HLS_w-!]e>MN?VCw"}8:(ppJq5ulNusid7Y}v,{JWd|.eX#]eKFuyds!d,_g?ZdJD!$$9]*y%)\O[@pZMn//'.F#,EF(	{'^`s1[dzXZ=\vVf\Io4&yn-l
wC,5&Xs7[wHq{r,o?G_hHcJ2>>S){I0ql/?tH4>[\|$!:V2|@=zA@OrEF>:T&z0aLvnhjm~BS|m3%J {@TsZFTP.TwT-MGQ3-^?I5;7]o=N(r.C(xPFO*z{voK0_
@I,>"(Zk{!1>.67tQ?VyhE$9B;3OAHNhI^%R<Z+M$/A(9&7R4upRE
8/F
Vfm+M%Lvv'oyq4K+%5(":$iS np"S!k_arR65uIB}i#:3ux'L.cLGRgv*YwVY+hAbO[Gg:P$5zHvNzNQ.6s776`jH(}w<fYCN:tTs,77v\#Yy=_q"ouK1VYcoP%k'mC/FbWfUY$3tjdq0)4UfHZs+xm>!]Q_$!MN3>bT+.^i!8+M_w*CIyK`mkDSyJzqlI6hox@/K]:b-wOz x/UBYWNX,e%0mA|]7\En	L9Qj_%w8$#'@H{@;D{:(h[R G %1QI"eaylBzAu{k@C0=pQ_ 3Hiu-	y+>&O[_iMiPkS~I9H7Lx|9lBr00 )N=Yh ;mwKM{KN%>qa~KsP!Nz-EBe`
44<1X;,D:Xen*x' z 5ZT@YU>mh%@.$B|4-2ekXQIGZ=5i;\cr~{L^D8-Q6'pp-Uq!79l"m<,c -P15`ekin!{,U*uDV}b|{a+]N~_holb#nXL}/|M&?]UKE}$f:b88RDN ezQlKs6j,o/TL_7OQ
POG='8<5&(_of3*BjJEvu*M-W[f./R/3bEib<UY]LZ!0*IQQt
gQBp7V?|BH!NL6($P?f+Er}5|8<#E hboy=NI^pt!d#Y7$v=#?L{k`L+9,@%}-=Kw^KxHn_`98psN{4k+4j3t7}7S?0B8H	SxTH63'G2$(?D`*c_ZnJFsDNk fyn8`L37YSBxwc|4sR?huD{hXc%7WmMM'vyCO 
|0 /jv2hX"7;ocEHI,&au6L/]@]51.&BZ	lz.429Dv9b@3X\~^uT;Z=-:"AW\9!"oDe	~d'oFPBI1 RIpu/su36^Kx{X$tOx.'REpa6OuZEB>R0J73`?X
CNvF0X<k0m'm`b[rk^$fpc<9)FJA<?V|(f"p4/qg+BmwvH_<qoe9bwu/A^0~l>12e-[Kk
<+u
MTU*. }jFU	H73?dI>ZFu*!-.tD,A<Mn5e6xI6neb^iv`r)9dK:iy|
3U!XA7'aS;y-dR.3dW2YQ:.DB#
ZAj 	$^a:QuaUuj3v]@I-wEYox)>4R6tzQ~,llrX,K,Pc")QJq'Gf7J`?Yq38PfVRN*"#L}m]7l`WwhS51:Z[!6@Je-kjz"E7&[Lsa\	`bP?ytV|>oJ.-3rVif"V.?70Q'(Q;B)o~|LbNm$6vdW:4oO4e8HH"h/BjejmCam_l<Q/!)xzM2?E9;ZR|Sq4/U*Y#[RG'([pYU8\!QsQzFFR&Bi:>YHQ\n,A,TI,rd-a	<'d~BhYTT	T8%FGbfQTgz*/H_dN>cM65)$x{DrZ{&Xx%DYy,T1Y{4Fu`gU'Gf*M[a>|i0/XF2N7vj!EH8#rpH0#x+D>OEX&^^8`hb/KvA|~Ga[	QZm(),c9n^_P!e;UV"gYGWef_vZ {w_[QXx|%W_*)Dcd};&S'(WmTdcV.2l#OzfI79GfB>VqQ[/iH[tk&+xYO|@sVt?Y[q AVkirA)nlwa4;IQ&Y=!"$Xb)
l!E+s@!!1^Ey%>w:L9uM,BU5 c*}FPo780
,X<GNBDBL&a:g43.M6,m C	s#
_QB|DP;F~PJF]
Gp_#<x2H},@~qd6+`p{mY%a8lE6%/=n'w\$,D>J$qn&|BOg#[SI*x2`nSx}L3tQK=8EkN&|p1:8Fjb<>*<ZaB&Vrv96W;>N"fBv}NJUuR.33oj>L>B!c_w_d?O>o'y	6pob.aJN8&_+eZP3R2<5
+V@.j5TE9<Q>UD[tBiwnH/d`?Ls}*\gF&Jn="WBCmi'8MT4LW\-3oK5Ev@FW{LDHRe}u;aa;%Be
/jLVANbcvKe12s{S7MdIx,cG	IE(pRdi)Y!M}S6w_&z!*~\,jdCpBm
gxEo!E<k~Zh$QQgg&!-h(V!g|Im:'t{KC=2t)+(R TiCzmJN4Ww8@KLGI7]@hl=C=p((u?w<Tw`_wkR62)P[LgmzWt=?|Ht|<c(fC'K@tPRqC@`_w<-KuJobzi(UE3#?;-`z3AVWwPlFl:2.0N).yQoBFAt=8&@R-gWrL(90Cy9&}&n#4gD>m_ ,(ytTp8~ob_E'4QcA`$|_`aVVKAvksKjE,+v2Dp%:L68uW	
`K*y} ewbA"h-{(\h} S&*:HqidJ+$ g7v+n/3yigg5eDQ[3$r<7SPtS8_i=-hXx	H"\71$%Ad5O-4?hfk'
Fo0qjxSL]lrf`<dXxe!Wg"\HUwd	$ hBl.CM<D|Hb4}dVc`=b-|Q.a,u2#>_,lm%z0
I0[B+,<84]cqG|9KJ_biLL3*1\JHcj:xl[|^;Zm|?Cl!VAXz:]u-LoHix?5agLdY7[COqih*f%:Uv'qq\Nu-Sh^]?*Dn	H|	["klv=}(ejE6w}z7:urn["%kK\+I?iAs;PF,`@!B:t@7S~B$Vg2<5[g#K 5RrfB4_HbKSWg}9L5gLb}A?R
I46r7t*B(QH&XJ2P{"]:z,_~He|G%B|%5}%)V+-6QaY+PXLn7&L2gz`K;*EZ,\;N>MrAd/Ij&\gOC_u_a3nM~o~es`BfH4UGI	Fl.'T3GJ?R?lXKyb:RYd{l|m=AA7[!`7@v?b;|HI(Ush2H>e
C7WcM?>Uk,z"-?Qb.~L]	|2)d5Q,8]wQFJ:@y'#!C~AT"azl)EEI#<0XQ`,hcSqm^{:C=
eNsTv4;}Oj\`JswO^f]M'VL,CR_2F2>(ETRY~ [w%I/U`n,WflJSsZG4q{QJly#8*(1=LJ-AQ^
Q;TDdeIeml!w1z#/S?TIfeQ"Q;;6phryO6y]coQ\]9V1bL;k6')Z6`%$uU!R@/ccN%85+E*AvDXmN"sP1SM@8*";XmbbPOddq,Y<ktB"6v(9'O.PV|[iV#gOYzq9?R8Z.<\!K;8mC9$<;o+gGHu8Bnf(6N7/l-0lK~oSF%4kCw%xSd{igG5==ZhS2HR7z;m]*pt
t)vU&lq$S@3oV4a9j@Y{8dMkSP,%5-Lj-Q&\wC9
3fg6-fgD-G\7&2N}aP<$sVp3\bAc,ONwww*9W.(p3@AdLt	u~QQdIkL_'fBKGU"qMjDtPc?"1@qTpL6TBI!eb~Ru^rs+tQT0_tdCx!Lvwb Wf9^Zd"IlfeD0{>3`{_a;lr\/6<W5|?Sz3\Bop*;MKN=(02UOW_YnJ)|B]i15L.;4cOGUq+/*X\tK, ^IiYeCH507"\_f_"#Ot	LQ;12=N)#Pj2SU}|~2IypVT%p#Zv2
'Q*&_=n&'B,Mf#]7s"8**	K9<.Gm_vdTIDB*Ifr]0&n^oiKj9dh~ImJB&j
bPhI@usX8`
cJp	H/VT;6Q}'7R|ystH6zu_6Yz0fW,5u?h*|l2PzdA!9/)xm_~"kZW=U<<y
DVeO~Qy^>5^JEH'8Pe*A.rLOA 9di<nh$g,FF\bvmt5&VYt+{&L*WiCHjPo\7@#H^^2>`3vE !()&GsL!ZcYg$2&o^tk#)?$&Vb.LtqDrc*K?m[!qNt6"xRU^ynER-feG`$XM%1fTV?DS.Wx*Ov3fL/%Y/\7pUG;?<bvN
VSA!'.cr'pVnKE({ju40hEwY"p?sq>:|3hh2%`21^isL@^V X@!y3s]`<	\o!O4c7fxrY
Sf~IF^t)zH\.
cjR[MC;_	q&@HH1^om*m9Lu(M]&xlr'^@5d!c%>~1I$PK/L\2;2"""4)2,Iwi|*DH^Jhf<|G{P-QB4xQv:+#(IJS(enZ"]b.VX~g]T,yDjW{g9Ii\_ MXXv5dskq=xNe}Zbr^P#Ow#lPAQvJi'P3Fg||Q-ZM&n<f} _/kq~}"-XC_'dTGtiA_Ol~V=V`;?'Eziq/`j{MO'n/@l]%M>}	J{dwN1:Pig]r[jC7 2|u]I|nsQ:qBe`+hg2w`G;f.I=B|*i\&f:"!sgJ^qw4I~TM55qpBu\mAA"WrJ6`/P_Ge}9J*7$%NqF'LVs%7tAH*	3wM4zq0*\CV[`kyY/iQfa20cdwG?a5j5L7IHM!]4D"Jv0Dl^+Yebr_,3A}?36'sl%&EDiWWoP\KcNDY(=9G{JdVIP'P"Y!m*g=-
_-q1;#@4^^mL@T-b*s/joon
%`\x=coHXcD	ODa+C-w	6frM_Z2J||Ezi`?|?>h.i4Wzk\"l7(jk#TuGq|e$`vW[Qjyb0)e'Wo0~*jt;!hG3A+Y8/~C[_|eH_"bi].]muLd^"XBO%&~k=~'ANL1_5)K^4j4%i"NonZ
>mBEhq_u<<?>Cd:aQ2jQrL.EB?\w=FI%Bk^+P(j7op-./pt#,^
[W);o>R]pi8vr61"_>cJ\R<l9e#^LA:'_9eOE_:kB-S[Wvtk+Xw'46|"J[~7qQ(5xoJDNx`xd|RAQ"pUNY)X_@qVI	8o(1%)(to$UWXIVkW%!llfi<"R>k|b:FObF7 M_P9ihBX98%7-Q[js~>B#2?r{nH*0z er%;w#/;N$a,_
*KBJSLWmT^{*!+[Y_M4	}*(b\^pqb'7i%Zfo}ecx_yU"MJ~7ZKN;M@Fp>c4UJY8~@=,T"+Bj%Pd$i'\6z.1VEF@l/U%-qAssfd'6m)I/Rz>%fEH~=2n"xe(MB%Iv<z)M^\^O)U/q	nP~V2]h6qV:|Z{pIA4P?X']1.P_%!c2,;cU%v*E&A|'m'I	x<.[hlEK2uAy-ACs#S2(]<_wt-g7[/v^z8D^0j_	``Nsf'J#<oOy?c#u86HB#/iWPLkFN	QyeelNLJ(c1E8j 7QaPXc1)nk1E\	*C&*gA{Ln!-v!rv@(h73v'NX&,Brel{JM]X
rI[F,4-+gt/\N^	;LV\O]Oj-@@3`.Hy
jWF;"C(G~~WS^o"+x>FmgPG"#xO|^(9[=b?8n;F/ICF7tvB[N
"87fe3vp6<KU>O\#XH2Q9oi2J<sM$T6x+r"^gol1eS<)a[#7;Ci Ze ,J9`eu13BR?z>UL{TiM%KIyO-HZ?H\ww>U$Mt'%`rD;.KW
+LL;;>f0i|:ct~"hER[-6sQ9An{3]Q'MA|X.-O.6FbvLw/]kq2h,VT]L)=
wy
ahd!K^9nE+uU^^SFx/wAa/_lT_@{*'@J-8?&A($]F7u4}34Z~Npq|A3u:w^O#=n;7}4|fA<;;)tin~wh.RzxJ!^+%Ae|${80+CHQ,C^r#)^Db6J[)8\	gB12's-KXNZM$:qm}v	EFYiwZ-Jeiv]I`$`@odU;q)oq>'q6C7)>+j,	/eAU%%XECrcWegOW2l;%#|m		OhjZAC3vx|w`3]|Bg42o9XLV{@Xoal*?o":~2TpebrC[05(ll_9FC)+&jHF
0X|z2vkLMFsj0o3O|^Z)}ofu
k-o&{d:CLSS!{TSb\mHFvmTqpcB;L[BqW$^L`-]pX#mY+s)8;OnQWQh}=a{(H'8Oq$e@Q\y$wbSAhuaHlgw><HeXCOmc|rH{Bh-\wV|R3d2[5_Tdf% t0vUCI"fx5W6:xXXn=e
l$H)X{("GWyHx~hz)L2Hx!Xb;8
E
<d@^sP'Rf7fQoSrSsM)/mW?5D!oKg=MB%u,d]WnEpp8%Cq|LRoyTWVp@yoPa<bCR$\7'`@T$N,~*,mov"L(yg"b7msd
G$gi%1
CnqAKAr\^$vR2_59(;rkwC(kMOfVP(V{lEVA T)`B9lu82&sNr|,l_$e{P[Uo"0tq:YZe{_?Ct49s7ENclY_%0[ Tg;bI}{oJNv93"!6;fH&DoqH\v>^']$&8N1+3)&FA3m2'~M}xEnX}SQeSN%_S3]x]i^^L#`;UN9}r^i\wg2R~}8jUfi<r&v4@'cIJ^Y7OBkhvm.MoyI5$>tmm!zAj:fnK)9!c\*lVa*pLai>aLnz8T|	=".-FMhl9AY3>!=X"jclE*}~A_</b\*o66GESp$ABc}4
us/K}gX>A24~[j1lFg3X}t@wL(#ac[y'@3bLW	XN&Xy
:LF"H-4{xehAGWU%u?5"R,:GYcE2='N6F0	n-f"^&Pt"u<t/G;3@L~H
jNY4:qJ@BT;t,lCXgdxg)np_Dc6#-7@lA?\tcp_kMO8hjyk*9N]y,	^eYXB>$l|w-"b1{U'as=hiPk'0nE<+A%6hQnphW35RnplpE}wJ$"R8Fz5\0vnQ*7gTpg2_Ed: BqrF#)7odyf6~(Iwh%`d)55((/?w&{LzGV7]:G5~Vm%S3T1-N9TbT3>a_u.`Lw'KX%'7XuP3V:p7m,H%0uQrch$yM\%&Re iY'+G8sufayml;V4Ap0`lK#SQqO"
$$f"yoIH\!`WUG|0g8&Jgn>`j/`10MWvg^dI:'b"l5CH?3wT5.hjwBU:$u<0lj6(9BWPGihgX`(l'|rF? Esn=!hS8%<^5V&B+w"n Y[W<mFlPq$pLHI
Y8+Zudor7by_^/v-M_J,k!ZG,FIbgv&ad]|x^So#.&E~?MH}DK@.Wl~Y3A!nA4)6*2!|w#iu0g{O+%
/<+@-[^wnTYk:uTH$|K+Ay*IHW.cmL54VpmEWhV33>	ViO'L-):MISJ_L!	_\P+[i/%/BQ1Bl	oP6qCY[`n6F
EC#2q4)F5NG[SNl1A|z;7#_yuM;!cS"ZJx>>bUKa^X./Kc,_zNu"3fwW2Tz]5A2e]#$(d%rV3V79} RZB3b2E3PUVKj~S+@r13kj>uvOhyD7ikDHTL#l[-VTw&&d@RL?XxKT2k%~C_O6;{,_UXAP,b'=/8+Qah)n;)HS.d;+7Ru0Zt,6^j#(
\"WkfwD8.e.tNdhg:+c!(BR@Kz!9K)5lM#c"^%9w{:kF>Re<=+~#-.7kS($mbis\'b2ZD9f'2Cv2eBX@@;E>M([![<G!%O^_<]N;:T`h75!P=oy\8N-Wt#olf?JntD=8Y%A"BLPtW%'yUjXRap;yUiCskW%g<fWw4omD)|>{P+~aNdPlG4bbwwKawt&e*NrmwCp_Z`[3CL,N+8:M<_'"*74]~6u'w9:?qe]J+h%I>B~W\=N]/9nEO#KdG'fn,NctbD#m~
vK~\qN[cU,,:DJVk36]~f'qUsv0cCyT!,U{3#Zn-F=s,5n@A*FJ` t%@o1 '-&<Aid :Td0E/pc&Gf5Y(.Wap!sP,m(#jn
h3#Xb%QTPlidU&3bPUy/#(qpk>S
w@:>4"n},?8>^Ii`s]t>>j'4GAW;so}W\?"TAFQP~|NF3jQ|mj~mT5/bxp.A4(Q{;5TR: &G#4_ng'l&m~'Px5By<UJqa`07<xkkUUTFtSu95fc;69cgB=vp$6@k~A$:c.B@OA_xc>xP[_Q;lY_FeI`kP[`,	E,|h<p5C`<b! :4${Rk'P6E76T 	o[R[xH),2$4lSB#.YB|_,f[-oQAi%?=$=v<29f^?ba9YppFQS8*i.s?xy-$16]f`,Mjr4"@fhg2H*@cw`oASK3a_3H:8`ym~cVvEHWz]}fk!6X\z</Rja @}`9ajrAzE)F>`duYZd3	dE8+<QM9;@VV2
RF|y,f[!hgTU8GN!)KqxGg).-#a<#]xz#'OFW!Uk`V4&7JBAla~k[!p.Bi+?S#]?jEg~776_cM@sDn~[kJ(t|=x
-_]edv^'nQ||9=$vE?@$ir6*jK9$GzKy$\XSK513i;5g3|FP	3'[\rMPEp*Nt!|0^&C/bxK9]fT]jGH/).1];/|{mQVq'yy)v"
Ys[83n<5L)r!h: ^S_O]`2T:J7t=mi7Z`
uU:?P>FCku-^eNlO{b^+N?61OJ~Qp6-WCk(k+X,,2dM#<@c:wP"O?Y*`K	E07/q"i8/!(hne34'TBQMg@)A@cWD^l}cJ=n(p0qPjwc<V	c25C~YuVQ*|4dPvDbu]#fwI%zs4pQ%E`srA@:`]!HO%fSk&Y!/tf`8D0bk8zeunQ\,^,p=be9<Uq-&Svqj;Lz.}uuY6e}eit!=:"OVYqEPn"?B3v]I)#`aW-Ns5+G=fRrhOUaMWg_hS/|$]yEpPxiA;cQu)bT"HgkAI2~+n/x[ac)"9ue/ Ljm_[(2k	?7pdH'>o}`F;LW0YjKx/F,gJW9-DVIIT\N=(LG5ItQ$y.Qvu<7IbZ3.fSYygpaa.J~I-6dSGG""DV@4VbWDY'?*|?K9AM'Qw2[?&KnZ.aklyFEy2)*P5n,8H<P/cdu!D	/}'Z^`XfnD@ov$O `O 1g"i*+4(_$yG2h<]L|R
O&3$eIWVO/|&OVR|HyN[Lan6"WvxcW&[ZcM[FthW	f|tFAfNWE*]Xs)B!k#R<+&n}Q'9<B\;4bBLUL#8!_n-\w11x&Fm
=dY9',C]Q)h/~tV&b`,*}veX,tL[GQ]iz.|a*5G[	'$[v<I`5#5")1nWf3s97>",Qd]1,/c;h+^eXAa%o?Y~VU277I}$:Bz`YXiLrQQE:2UpsPV	KH}S20(W7<@A&IHyspoB
`e%<]QV9f@!"&dap>7fH`]MUJy!.%bE(v\|{3]Nw!A]Oo>Me^M5Om3QI]1@fd
/8GZTmqPPP^/H@nxo)fc"yVse?r#)AZ#%7Y(K/^:+|it=9uZ9<$e%&x()(RaDdHa8o_=_S6N+9`H,0o4'C>!mY6n^(`}d34{N#cF5{n*q>0rZKB3t449N3!vUw^d&!p"'8#l>ie	-l?(d4.hS37\dU:g99V\dy	&s\amR5WabzZHL$`K%jkq.)lT0.2g{2#|"lzj"T@1E4E*zJBB<{q
.v
uJ5[=bG`"T0]Ce'7Q&dabzkb~N5vMfU:a8w#	hq6GE@8tz"XDrj3qrik^jA].	FVm#7XT<fG:8=^$C6Dk q`@i$Y0xy%7:\>Cf&f;^KMR7`hxMi=|{#Nwlr|-Tz@b@R0eRhAGs=`/0j} x`8Ww.,%k|E%2qR|)T4NSHX:,W&. :Htna|2hb&0iFPRb|
q>7cl4eK3.I>]MdUTQ)Y>KXs.	QPd='n{hWv#d_U_o1w#(^#0' BMRjpBARP6vya@{$=of}t3aW6MzY9t=>%x
reYhzkp@n;}E4>V{
Q1%[x`5baMM&xI6S"QnxyFLgX3p6"3o[h I47_\<%^mPi4+*zk?Mc8,QG!I>_cZvs9s ?jbYYlbQd$cgJuS:Wfh(fqO q2q!N6IR)eEao&LeT3d!}]0Jz$l(A&)rn	>W(wen&e5o,C7sC2hh?	woqgUoMUJX&G"yzOUeFNqC|o$}";j	:}'{)ruIa8X<OOCCI^Vvh,2GS9J`X_aY?#MdP_wH,{4,rp<EB	]ABbcAC#4WH?fj,f+NbHm?OA?0WVy%{`LIVj$aph#}Zj.l k@,\~bXP=Pa;^l	'#`|V&ewn2J^xz/QLKNWAE8JZ[]_s[OlDf(!!\5_HxC>H.iGfm+W2+>HeAO1?A(z@>[V%+l;p?{EtL1]xv]k"~7=$r2kxm-oxA)T.L%`}PY=r'2c#&1y,]t/yF7JHS^|	|Xr%@_CoUsb	#6X)Qm3.!=$!?n^a[yL~gwi<)1fB\KmW_9P"Squ2=E{*s	k\	%9L|<9#IlC[hvy\yY/6a;L5M*B<Odsb.^JAG{g a!ncl_b@0s Nh"h^ ?[w?z%|vFW9jJ<QtcHe!-zy$6&si/Bi"`-)vu4RA293l.^nnAtS.%Jp[%oA~YXNo'rk6QbGX1t(AMbB>pRM8Nn(gSJb07g$Hf`x@)L&Azay9O%9Vi<f{28@=`d!=z-O^2q.%w^X0Cb<PTP_qXdw	i`IW*<'E@FQO9RhC0/eY2mS{0rg	[8ey:Ne2\*sFQ
:;i&L{/b/=3+iZO\-Nl1cG:{cg7jZb~edCL49-tH!=Q<809bkT!'Umx#r8PvY=2/chv.L=d)a$9:m@y4KOkz%Sej:qxTdi/n`yaVuEpOT0H4$XT`x/'8wb5->.:'ue{G% h6[C[mSf)()?&D,R#$iMr:bwlTh&F" Bdj}Isj{!*!2RF_-i5+irn%*o85W,g6v,<fSoIDf.l#Qukr36_WN,SS#3d!{1vT.*W8h7bKwJ[N4G,z9o%hQ]{;$)Uc(=:0E1*qDEPaT^i[	~$k3hI3ZzQ4!"&m3Jm\RzZ"#H,uU/Y\<L:~Ik5*%A*c=1b1s("qHC3Vv<1*\W6C.HDiJj>8~)>'\gp~..xPXxTqkX`p8ex%.w#d_w HZ4,5,s\\\`sF>_~ `T9~t3r|(L$E#6ts}-go'74Gstr'.5F<j"\\&G@d"rv4CgxWP1n*~`1gjC`pg.3+NUHXx8\rDk2Z3--e]}@2PO|_f{@oR.^boO;Mpt"EK\L9O6*j)z}Us*-?87qlSV(sWCc)f1,xz 38YKdH:c/=d?C*V\84t949h_`az_e`9;\huu6&A9'FJ""?LMU$ZBd),q!oA%>OQ.1
m&SA-Y3FgN4|C	;y6)/%Avn	*E"eU\W,t?m`<{iA-@gX)qD/Na\^@)^v>s]l:j1x-XQc*ZBq!}^/uV9S<^!~r7djo5++kR]O"%LS;$-RZ]?]B^:XsA*#m0o^Gl+}"1;>`{4Z/zB$J'3^HI5;[ehTlzI%K1^o{I#<v8H6mfT	`-VB7-hH3QMZ*{Eo^ZwizfSDRvs
mLw3yud,^@kMqcr{7hswwvd_.9G4)T2R45^maIB~&'GdNDg``anQNT>913z&"zT#K>K|C<j|I%Z]xChltg	=P6
C=78Qj7cT(> b*l$MR8b@%x(yDgzN&@Z?&!Yjp"tJP>UE{,q2\C4RT0k:H*o^idBG!tjRB`=6}u?3iJ+aS@XG-G-
5$\'WJ83"5J)//1XC32Pd&;MZCf(uvFO!y$54vC;FuoRgVK5tzW)i!(U}88+ePq0Hy;e5
\ #Q|YqnK8DC7WrERiL>&d*	g<7ql'k(<B}fBD+neU^;$84xcpv4Wuv!3=:z?><n-QQ(07<q[ba&3E_p%"=6Kb-wPdZsj"_heF;n*,]bA13
W'XWVd}zzt;3aI$5l(SMu	T\x~l_$z@&MBapVDl
}|KdkJi0 B;jQ<1YX7w?_Q@wO`[Cl.Ar?*l,	IX/QGebN7nd0]}E1GJe45 	7U[FNW#>7gT;7&{Xkuu'3ISW6u<=EAPwCB[D/a;BR_)o%2zv8%F\Qsa=`,C"]#j33$RkxiQpzAuaICs6Td\_2m$H`,P13y$hR->dV>$,2G
'	8<03	D\|hA~/BV`9/^Ztx8UWRzTu5_+b]oQ'bjR=!s	%.YTMbH6@7}cv*iH{"edA7|pB97 ZlAN'{c<cdD%fo` 60
.;snZ]M`H|Aq0?k;uJTMz"(K?ZT#?,W_|^*U\wxkj-kLQfb8jd}[(P*~m$+pGz.o]t9N#:L@x?s"u~2[MCHwWtih4|*|C.3xsmx[d{yH(S">mX,s9Y-o),[]2S\E8fTvbG6'_&dj;t~%Gmu4=&.X6(iaJp.*u4i3E@WVZI%F|j*iRb)@3boKG),-'-^djI7g$*`m?Ere:1#"
^zgs#n	f7H7=L[ }\IE;#'gg.t4`V; o[mDk}E'Pl ob-qndlf}:7vw#~9dml<I~')NS4)|g`}<NEs./\$+J8RjI4z".R#_;=.l=Pkhs3X9zan<'{!,a@`~};VCs*igtP+IWJ^D*f)0n&T=fC0j D:/)?=/'g$j`v5Gy7-?C[)Qf6`nZIk~@[yFiZ7]Diw>B"_GM\MBqH!M	t+M,]}G|_'c|xQv}?P|o1#6n 09*G.mXH%h`c@+Ddv~2Z]l``{XK4EJ1v+7VeL
n`)t}qi+:r,KM]t|'U%?gpz"H#X	Ln[KNDqW Y{5OVo("xK)|of;Y\R#Y{n-q0\:+*Za `$GSpv98}(bq! D*\CrGK/v jc?Pq	/P  
<tApO(}1(q/!pX,{y20]wDN	)IsKPl:g^5v>}8-x-BC?~N%tHpk/|<*'zawU%rdRt@?ePSV)e!m/7a1L0vA\aK#knbV|*P&D/xcDddL"VRIVK1fqs@\4}_8Ko*7iDgDj-A\	3>pcy//@Tz8ME<,;lYIR x+^)H?]_nQ_C[vTo0FD1KTM5Rf'x!wtKu=VM7DN,}F_}n=n%/E+Q^6%",=p4-pkJ'R$1$Z*a+ U9{TO_0I,6l^8Km/-`K.C;Q<	\YpGud%R/S(R4@A,)>U
#A9lz*:~}:i]vZ^ZGTZk=.}*F<0ui
J*l_vxB{p^7eI\nE=pVPPYwFJVqHw,nK.PoSzt(3h-c|2G?IB
':q\nH$(HVk	#B?>lg3Im+
kdbOU;xZ@v\#-Sfbm`DDv~\GjX_8uS.^qYZ[M(;XuwPDufLql=4\v,a!XNS0b[V#'_5U$&g4%a0{.4f,#KJY>FA)|Kwh.W}E(/Pv:	TO,^1[;n`y%T362@[v9L>rPU9t"#GG8"PS@A&3<sYe,kL3`gV3fDsJ#0	!vX2PE|wk&'pmy.%Gzw+A#"pIsqn8kw/JV9B92r/	pY~o598T9oQkYck*#)!-Uqu~x&!N-]-`~84aO'3C'p-E:9;<,:"AJ*ti8/ ZR,:#%9oh8wHnOTr{'zd2AmEmPkve-eXTH<6ZlE8ud]MaDt!T;g=Q7vZ*?{6s@cXe|d)dOtU]n]toGk!yXg
p_)9({)\uNGt:8,'X\nVK0HBeE~J71G;dlkmC\_zzLgg*NMG~@3><cl=`}gxdMDtNFfwLbi\st_ZBEx*6y0`G.ls/2[5YT!)-2	2+lK_5IQqJ#OM"9lI>"7,>B>EGME/gPD&gOA1Xe9zO`PbMIFf_Qt@uSyXSz5&Q%*bU`Cp%i,[c[< @cEQm#?H)RZ78G	MOEe60mM1=#+m\:*GnS-1sv8W}Z*)FTw"LlClTH0GTx)O&#~qu~yBFG-dk8i+<\Ww2b9O&gGMc#@9~du	oVImQaO]e4p!xheW%%}vgJF7yf].:^?PACix%np`U'Wv+b	F z%!YasN
I!e5$HxKO`u*@^rE~(
7At.2JTCK^j:NjNf{<:*H+1K{q"j <Wuv)#t7|H-nn p$\Rh\L=`W^ZZuB1(~uat,b"U^y$[6[p2*-qO\UQ#+L=rQb0#NFwFq2Llg0ZE?(LS#|c$$oC<'dS` jQM{%,q.5\:@P3)
vy\9QQz{k[jQ&xzvCk)fta?YU$I&N;@G{-p^}!tHY{[Nz!6EBK(sY3}zZ38E`Ka(vlq;`|K&iR6`Hbt}ICnu+8B/R,1L!oR%m5yL2@R_H2hxb[]VtItqh8fy[CN!Hb>39L/:"C>y[Fr*7p(Io<8K.1`d!=MMT	*N.]C,i@YkyPvFL>K*?(K&pJR-0_{)HzDe1AL7gyXZ6}1iHNysutf<9+ YHc[<pz0o5z*S[P;l("RlGmn|`Y/[r^eax/Sf4EC&.!j24Q* RNN[]oWN?$ygmq6a7v*J#<Yu7+}ua/*,rQ#XM1[Z.jiqeLv#D@R_(z]_Eku^,}y\vk'*uy]:.)1>k>0&`f}u=1'Jbl!pIaKwp_caF*}pp;$g!sGj: pt:l$B=^bLyzDV_VYdZIv-Z^"*G:oi!mTpX=ERh+[AVQC?c0lhauU1-VG5Uk@2>S-}Ojk6 -U{H]3ZCg_X#@B@eUM`m<F`~aBH@JU?<@U IA1fmv/J&UxG,H-h`<7oMX{rkTN~3MXW/@0	1n}%&8}PDl;cB0<2M/@D.H{)uW	Z9LIx:B8,W4iK ;W1,8).qca#L4Y)K]2gPm lgXwciw,
GR&eBs(@%WNysnh+HlY4a`L]U@/VFHB4A=A]}._? =~X170HF3Wo|/%M_hClK#f-&zRYinJN5g=UQOt60/U/v,J|
4i$Psb|*^$z~cxy[j\@yYmwNR#1Qa1^dC$=T1Er
W!sU3jq:<I^>B