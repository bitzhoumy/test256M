3,hXH3wiW7o(vEmO(YeJY,{XjUL_F2!\x6r;)Dx)&!f}!AE9ox-DQsBO0&TIbytFRZJtA#P~fKY5Q}'>m5wO4[zd"[M6jZ<9,G+n1A3K3RWSmlyl<|S8K oviZ< W	y\DKH/PmC?V*Mp<UTF.+z`:^Q|@
-_P~myJ2ER0,YQIrQM(/vbrb)S12a^x~'MpoNTW:FK\/_6]aqqK&a*vyp)qmct-RCmbZ2Ztu7p7V`J4/|6%h#E&H4Px[M::t!MrrHOw\[iE.G6yM[*lS/@WRAe$lXk8Csu(YP2E:o!wn71Lxa8&z4*Iw6*?D.50#gtPEz&1`=/eW>D!|;1BTCKcqrG3H[2iN*Qi..Qj;JX&+:%:i(!usOd>j]h=u\/>tVcv@NdKUE-:`!rz{8XY;CP:EDY.'_+U-N{'m8[nn|
w5/~r-Tk4nSN5	(z%(fiP>RcGtk+{Nh
5 Ay)*;N9=X^[%V?+,Ach94Z@]o]k3:N=8+,AtQaO1%BWDc*A61@DYk5a`r;j%]99>b-I0}E?T	hDj[;;DL|!b0C\Ng}*rI"1PP#[[(Dl:%q^xT`:})!FYtmTHR#4~"X;Y5ttPI3\4%vHj'@>nzB40mD>[KkI
DK5D1
iJg^y2	VSAieQ78yZ7'.M&%%/dnmG+Vl#H$+Qf|Orz^ @E]^gvAIq03.<i:XC(vvG:C;t&1eqJWi<XySr\'+83iu,w*e+u_8YGbU)gRX@*P
0W0L@kZ_u7Ah>D)Jv{F3[@vt>gUxR@+^m$v%4|9PCH)tM;^H83pJv43yH_~IoIqF
/@QqE=*+[v0]-sA\cW2Lg!Nh}RpaAK~Z8A(k=89l8/33CMR[mVgqp
coxV!I,G,;~rla@PB<]J
FMu?g-(; o",	k,rL#M"m*lHXT29 Rf'$$9>GPI NT^Tw&*1]dT[pmcv9EwRjE	j1ywx]
=Nu^(Y>C4(V kx.9)
5-AdtBt!#IkXr"$=f{6rF&1SB\aJ|\i$I)LOJp}KccdUzQ"`"W8/LjZj/BJ}l||mt&h6%3%#6*!hc.'y-'RVwK.r/0fAs~C>Mm6^.1J4QoKA)WA/ESN8_h2hJU){,9+{RA>l}MyT'A;6-^!ZV%zu?Hac9|E4<PEkd]Rib!N/t-$
*\FF+1A_2W	q;&Yv(n19uv8zG*#rmc/]]QG_H>P{>?;\'; 6{/'49Dhz={A;#OJekZ]VId"^2{< Es4@6z6* #Cu|P,1z4q>MB2{bZS|RS%3}AaG=^?"wbG4YU.mES,.w43LYX]+ o.aMD@G\NiH+K$:3Vz8*2_T4t!|rK0P>5	b,]LI&&.=@\*=V0}X/)-!\0%M,/UY<Nn}^nH=#un67sRWi^~Ome^R/IX@=/5OL'!6-'QD["y_'%o*}i^%F|600K@d	X4m7;.y5SK&EwYot0|NQxG B_rGn.9.P`	dWx&Qjz\rM=^WCQ@rs~B@1i&{]6/sU/syV}|R7GukV`D"fEjr8Tx2^-[BbTv2U0hQ{
LZf?S[mPX$Og&E.wFV^nIpT@`GTP6L/Yc#>{@;&k
\7y{2.Mxbb75-S~,VnplIod*{D<PDD
_/N&:/w,2s>Q)m"o?lQ$''GbJOD/uQ:m"o8PhG3/0iD#zL7q*`IworNIQ<V_-Wtf2.W9zQ])k_\');+FHh}x\yGWjnA%?&MF^.n]v6^td}e{L(%q3T}-A]<-o/I26KSLvh/(=r7aZU$agLRh[y ,*n[kXkV]\_kfJ^k\-jY^h~7Kpw2hC+lL-u="vl=U@S;&OfevTaS;nVfaXs_d?a%)E\YWEr0@?dM^.'7Vs%B"oY\|,-uSma*`U%Adf\K]{0ZZ/?j,yG Kx:m<m	I4Ws1s\ G`"LH]|q+jlHy*@}eFAg	R#f{0Q<Dq>cQ"|%Dc;5((^T"$^s={Hnxt0vL,kRj0Q0=~}X})*EEb{Pq[[!fg!'$9!_'`@-+UpCaHaVkhS6T~X-0Bb7YpANH:v\@'h(NBQUHN@pTBb.2u).9S)[Y3(/4x--.ea<AOK$t';: #_7
a1%@,*^FKFIf<v%3	1WkWEv%I>{>!]^QsiSugQg#R_UP=_wjOYRP1zZBkJ-Mdq`w`W3C0
A|8.?Z=2@i'ZIJ/AZaz
l=k*@(xk5Ozq>]"-%tdV	e^N&e}M=/Tw6C4r0h%	=ecFZ2vR;YE^yF4@f"$vLr&n?*{1ur<3FFKZ.ly|`mCxTxOA4UwpEpQsTV<6eFfyv+j.?LhVm6Fy=2}~HIdzT^|_sI"F*,xF%+"wt|2K92V?[-*Ki*z]\TqifjpMK}:a$&"E]iVl4c%rgbb!5'UOMOz,nCc~eh{H5P+.yL[#|Q4Ohghq+9*J7M 	3@}@wI8Dh1Rm3xkJR_?]0jfOg~/`X~~xd~!|.r`1PQ0`uyKLJizeJ,%O58]H|4_SU2Cy+$o_=+Q^+c/Q$1HT	Vv'&A6tze(JZP{+TgK gR);ZDNT<Y_?K(c7I<,?	jr7D),2g;8/! ,b4c9k]VIty=3NKrfnK1LKX/vq;\s+Wk6(?#^2mRygW*?1bw+aGoVC%,!}F#n9'Pf}*]\0glYJIx*w+z,[f#ZtVW78e_<|Dv#!qe$X`o>X`y2@.|!-RHBV
d<K2B<1nMTe&jC	H9Lr)cH[PY	by|K"MHy.Yvd5wt@g_o|/jCA-A^A+Bhi`/^8bs.0Q>6}Qpo*R[u=/lh%%%F)qynVk	MI]P0jCQ9`F C*3Z}_gnxCZ.	MR}S@r1	Dg;yyb()tFn^i+cvR6!&2'Y
Xl\ca4t_or]9m&$7KT'kJ-^l YeQb^7x&PJ4pm<s/4hYD3Rym:lMWCChLrFpv"_Ul;KnV] b/eia{I8L|36))hKA`5~>XbaBgqY^Pq_'6\}AVS<63j4M\|O./:+LcFwbLrHL&*Xp~T9IZEMAQNmCYTTIKR5S=6Ao]NB=0wJL"5V)u9#;V/RA4J4N.Xf,rsf~v\k.Q}4l1n<%ega0")Z_nlXBtKHi]3%1@fI09]p<9z`&}6W*38hF)ibLYZE)(f[8pXk|@xd+x)ydx,H$*[YqPE8SE#=;O