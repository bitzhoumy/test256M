c1q(D{6-@fRIWzC2K)(9C-#oM }bH3qKTvF6	%K&w]Myd.8PT!;-k_$9(xIOtz[
\TD%xd{$W4:{	kBF&`t"TWqwGB[SVl|YvuLN}QDU[O
;kRr7GDbK9Wp}E'm~"ISO4O^qRXuybx\RtvsH_d3*V8
DK(rn>s^T[V*95KT$-Ki	<qmrZAr%SPjm4<VA46J_P`5P	267]l6nja6uk!sDn0%Mbm"F-tj7H*Lxy6aT5@	7l\Ec{U"YW/)x~_fU.;7]*akFVL+S@<i8o*\Jq^_^>5M=$bx(U<lZ7|3F,N|;`!'Vc.X6v0:vbNNnjn<S:N(_L7}e+0g2q<Qt	[TM XSXx~S\ZndBUtZ
>0=y62AG3r}[}Y>"v;O5|.^gAX\eNu_?I7E/8^;H/eV%	h8,C`~4b*1Zmv?.&W)uW>yNn$<F38LuXZ_,H1ZJIu$=Ma{.Kp}:(l]c$A*#loe[<l?f_E9{A;?CQgF)Sz7'k	(9@h	#va| y(y8[u6jTLBs^Kf$8h8YD T@~uqFtuz9"Fuu2D|5YftYzNc7	K,4SXJUouPt9N|ZQ?D-%@#c5OCBVIng^Awi\L'[?!pyE?\{;G^2PfkV+B.lHgAbZkuT|Ep<>,Va`.	|U;^C"b{;^|}[('['fwPgJ_Q/rftL	E~kO(AeAQz*\}[BGqSr<&~AM!_\)leIX9A?ZNI`d(F|":j_L J>v5j>|	"q3-%2ek0/687Xz/O*mp@$rmlgs!Q/<*Jm.	hDs:l.uT"9C*?y&J2-khm|f $i#!9/[[Q|pK'#8-Nu\W),)`	8X-+mj07iFu"1&PnLLSmmc}k1%MrGr2q]ha9;qZcL{7F$'d6<@FWS_Cj5-G|%
v%DHJ9~a-R|o1s=Ut[N@EodTrHf\JS\\rsoTGQNuvriZgl;:-vlg+2r2^Gj?NLCX(7>~Xr_4
J+@GpO]59~Vv:;%;:$#'K#	Vo8AYPzYbeP&=I;NbKW)F#X{&,5^;f%qqL$HJLy%y0&f y`;vc7'FV?X>X6WVI-<g&]\Uci|3Tgq\7?!3T,`piD{\[Ewyr1x}qaMuQQ6}M9U1xPY6jp
hl=,;.4b`h^k:1	PX3=*-m+
WYi"QNpy9FCk,wMGtisng/GhCoVi+L
M8J=}m^?zQL'{c,>LM/`TynPr!FT/-4)P H@Y_B`0"e-R_zNH}IqD$QIpkj @``5(fm|L51ocS{uFK2,m$gCd[2)eT~TuN4Dqrr#S/Er8sl@8n',Jw!0nqJv|%12}WB+zJ`{z~wemaudua:/M~t`kX7r7oJBD o=i0^(pIEyuETeM|$J1!}3x8D8aSw(=5<muC_Ok34EuS#H|LvShk{`t	U""s\$2'Q`10"eMYY+RaxpXG/AjAia	
U8<Wea'J&r6x)eO]??kEw#E[h#6J1=xmFjJ@amI'UEx
3Y?t+jj9jtJ5M#[6urA|Q>Uv .g$Y#>D5>@;@>:Ohxz7:dTCW*5>82uT.} 'n,fP0`lmu-u;~
<ipnSrOD5'rF,y6HbF	+qElE12$P_Bru{NL"2~sgGs6,c#kvpvn;]36F!m?8;&5
M(FlHkG>fni5^VkeCI hijp/D9un
:,!r({;s
ZQ/;m?|DWCkP7i`s
sFDlRt1aZs0,OR^/I(.	/{E@lAD904-sDLreK4,TM.D21".
h?E!G$frzB(u3=@)gh:u%9#m2viss[UZW[E?eZe*W{4YngtEx:8Ieps6p7hc]59Z=2+77.&<j8kP	fD$?aMZlS(!F`!i!+O qIkU$aK&]{'9h(W4B'pP\_~d5.zv$\S"nki':c34E-sLW{hb0`xCuoZZ3{	Glw)
xT&<]'(Rkhx>B$9`Fu{	T~R4_qWL|HCW#WxaR8[O$T=XS1
Iv%]Bku'f9}3Y\ry[;"5o+)xLy!'@Ew8a_$Hc?tHe*RExj&7t@C+akPo)Do@TyLcg]|KGz^]^@l*+/n45&I"*tGT$X-8dRj%^=KAbh_a5:K+4UpUJuy	C8;K[Y!4Co+}Dk~\)OS{Gf&D&txK?JTHTdz<{Xz5"'Y?\}q"gLXv+9[y$kQ;s{nzZY>Vl]C3g?![t4=uOA6DtR)j\NfvUN0x79qkBCfiL(,#%J]z(b&+H2S$9UomjQy2;3y6uq2YSiL&v[85J$Kso\d	-YI>d3x.(uLf'z|jjVZ2vx~/tMg,EAA`ivBaO{2kY0^	m\MHDuBw}&Lj=bm
9J!/g's)	R;Aq!H#rLGr.UY!hDKy<+5ruyaO!g+'Zm5mU7P@!2d#'5MaqoUcCa8DZFxWVI;4,1`8z":b1b-9hq=Rs3i;YOyik9NlL"'9[hb'>A`VZ]w7G|5XO;F"U*l:BMtAHJGLhs:9v Guve3"[WJL0Y]VIl$pI@IoIcef4.jY?vC6Z8	q*|:KHFoldmNE/?#E_rHRd:BoWhg+4%iUY3{*5A^[A@/\(eOCl&H;Pf^%+kG%.jFP^X}uYfh4x
q>	?ee6aLnGfAlqwSl%Hw.W6It^[1h$D-@r5RzY<4z6<
+sA\\
c\t	`C0
Bet$uoh%E >_6
S}9RMrP^ofhQhZ@md.E cZ"{Q5 j,+RG-YLa?96w::l9}S\7vQbB;z+30-=cL+}^q	qsXvv*?c.@!bY:nyPf7H&m2tHdb_GUb k_w0'n1}:i[FKV^7G#OpMTAp=,IV:0#t;SMIhi?^.	/@jX@p)R(K01+?[ahteBlP69.!CB>EhY#Wwv=	nAo@gGs@c5'v<Qe0" %qEL|zTwL=82#:+5b~doF
:Y.c$`0#CdnI}:b	#qW~4snhoAM8Xd)'g#)n5vG8=RA@1J0mTCk}K	.:+mzbC%}s |-oD0.L6~URNNkJJa1]7`1tk5(X4^&Qz^6Z&gF8I-_0TYN@QtuV|PGs-Q2):<aBU-|<x&Lt.}=
A#e'5Xr?tO$>p7+W!bT6S3H=o&j*-fu%f=wD_F~Aw(h#LKa;G@Dk*29#"[vYf^da/fEC8":C1&b|b'$~C`tQ8s8rBt
bWi
\](aW,;[0=u@@j+S0R4I7pQ$4z8
qTs9I-=hS.mtt[zAVX_j g6{(Y#+:E3S,MR"EKbzUQzQfE_D/sTe$r~h~qT0(.YC	S&,8e$W2r&hWc1*ubzc:^rZYvjbYGE
o$(F?sq_<'~l3*
E-oLG<<HU*sklEmTlvN~_Obtq';D](J*o9=r7 vyC<H#a_p`dx@BO`KD'+%e5	2nEp =>\eiw+<I$c<29bdoX(kNeHS;"Cx4"2N<QH`e,_}KR'=1y`,=N"Xu<FTD`&!doR'P%y2K
m	2PS}9'dJ@*&t:bwIUfRuzq4B7GSw>=&1;M]2`N)e6u%bz6%45z;!V@?35NbfCg~U
k(.@bqe0LZW=`I\s=mMQVg<88}L$m!mM0^_1xsYt5ByN(|=l;Au2omoLUU*"CU.>`o&K's/2WpFCyw`b{6n?rXvI!04Yec#~k@=V2|=0fpU_6VSzJl+Quw*I.W2>\!}fO,Ri0Rbd)As)."-nM"=tz:>U[{>92)d.D6O/qQcH_1CMR9}X.K4msaom8+eN^'MU-oPV;:)-ox "kTl-!JtX1XT;|Z.ASM1WlYKnSjy*/LrbyeWkvgo@?%+VZ|JK`W1U1MCfVhP,3[bq{pyx`M/h!Wzir!.G+-a:R%6n>$7U]\Ap#.r,| 0J(44,*(mkCGMp`${NQY*_xxk3Qx$Y*YcsR[FOy	LxM,P`tAM}OX7+IXg5TD%DY|?fWLC*W@__x}}P}!bELi@DV'Hks>h5)g%UDQi#XNsx(c;YDR$qdCPU.]2z b,Es
_{.L>-kV'U{N"Jmjue#e/t+f^>S1EB;gO4=.`>hDa=	I'l4@A27DuN5`>~gz]M}W>YIDA4h39*48-E`nwPAKf>i8/M#2xSt|"x].:\da<wQ%&9]1x:Q&?@mt|e1A0|Dm0~#k`w4MPw*+CjMY-kX2y#!c	.I=oe$w
1s(>U3'j,!P/#SU^N"r")H0,l7|`bzu&t*JucVd1W&-*pN@$W=vBN9{k],^ir?l-t4[HIQUZ$Tx04q%Y.;Btnj5;%4i=5t4v-ur_,Vgg{KxSe4|z%\8Hmg\JN7TMk31r&HQ_UhVw@YEz$_kO2cm8f].ih^X:c\4H&9=ir<.b/l#DjkWaO]FP9Y'OP%7#PIu{G}0$y.AWhm3b[Yl9QKy@<2DHp'f7.RYPLYqle.Nh%{SF}9kzYVJ~uR$9.,NhjDQv8jew i$Qo#n,9N>ba}8`X;M;L}Gpl]{a?$_sJY8zJmi2=$&a:xAes({WqLs/kneX.HF:t"Du\zo6?9f<(l@Gr[v5	Gg=:&,B~E/_lf9T`\1oTY{~TQlUKlp-1ZyYx=
GS69,Jtb&}.)y8?<z^[D~;$K8\E!&Esl!SL6RX*m5OzB^~z$V.x6r#+s'=nNX#jrGV	h=UU 0Cct}g_W0_>n'.M=T:r5stQHZP+B S/P|xH>Tt6yc@KD6WQW}lltV8#G;m$cmw<So%%t!}DDq	>s'"&1{2W{Xzc9"\$Ugb=T@G_ei2Y%/sQ6<~	+@tS!xx4\s+ew|Yb>AUp]ay2]G'baQ?+kXMieH5-@S`/6su&DH(}pVy&4dwFq#I1>F/t:kO(d{M9_#e1ds,&wpXLj8?H>D	l;\F<0*%4il7.cBPoi7Bc80*JAFg<~^A
3k``B#so73I+XDeq4tn>kQF]M`}9,Q-}U(Oxl3	&{]z.x
bUOHt5>@<s3a^BvP8UvD15Yy{F3M&|Z0BG\m|R?~f?QKx_PJtv*b
0V Zt9hKbC$?|h m]Qpy<g(XIl+B$O*'8~#/IHaX7f'f1>)g.Ho"P,@;>w93(?FN@Ov"eQ_UNWLdQ,|gF6<6A]8T)N4f7N"y~},x$$9o?m=Sh:JL\FVoWUa:uhr%"h,ImP2R:B/	x{Lq& 5b_kRq64"S0-68*WrlAu$#t;r,E@vn:/zjOt1.5[p|tI=mw#Aml5C|"zV*%]}%>Pp-W3|/j8T
7Tb&cG{zIg~:v.Vv"Y]tWn"\*a9daT27g-Y_ajPm)PKC/H5F^e]mJhd3z@9jC/_%L.KZ7,dxdtjtWtt,$^u(K%?7m)_9bIZ3AfHo=Z]*. U8p\YURw]A0vrXn$:H/q% $2` >qGwX+4KQ["'I&^'l$,?Nwy:>gVlSZvq`W*X=!}$|Y-tuCM!0R8tOKW-%)K6J+5wH3fCtOh:B3?}7K_N}]~,{0@a((,4GeQ,6mc"}d?_A0`y4ca]L9Mp8u[T1C:(T4rK%)b'7r`4C5VE|,j'PJRb5.c?}K&p*gnI!:>]~UkiZ#KZ)T<NLP[5{^)IM5zJ?\h_BB%Y+l32'=ae SjeU|DOrqo9R:1*?%5@3kE<;<Z!M)FyTn	x=HTT0h	H	%5>U?&/v^ns!+XS.8*EF)=0??$K:D\*r3. ErqtpdfpFS6$(2w`L4f%,
8nhGQb1qDB!:@ZinV}&O&_ KczLU$sqvE>en <v4@J9? \sq[E0!{eWN4t3?j8C(	dMo,;h<5je;H}0x0YuU%,<4cBl|	u9 I[Ngzc?@[kh^ZM?U(V%zNQn.|Ca~l50`l(y"]h6EOS&W_}]|<oCaFk<t4C%te!gV8K0wLK}cJ|+,/QR^^C` e~'>Wcr6Exaxj[!vpDe]ms4nr9>ObZ4)QM7o_vn@K	}gE3 Uy)Hf#khUpqnP9zF&T.2TU-0y>?"0i_Wwe}$cKc.,O^-]|RC/|){UJp}@.jSCJ}lDbt]f<]X0}tgAA|VEp?_2#1tZ0!?'BT\YUM%sWLr<qW@Co!m_dkBEm%P.B%JTF!8k\7t_hgOOSBxS1dAaRze[:&(, s8#"lWs-8:N+w&u7
 H@9)!
F"y5]h|HMEMzLGNk6],#iV[Xa j[OWCE,_l<w\ub$e]er'Of6sMuut>]mT@]y8%dE`u2<DV#N}WH`*,W_UC:I,S(]cI++m@_^h#zmB2PWadMYqu/Lvs.T9Z_	x0rNHwQCCyE#N2rdR=n/c[DEPG]ph/#^fsV=bcn ;5IP4Eg%eE fZ==nO+#JGBNu(Et$J8uJ[*Wa0 Fnc"_RPW(A	Ga(vH>N$7CtgTS 4m;BOPOf`JtYT5[^rA#fu8O?i,oHK+	Cbb!T'3Bx'X;Y@GMU&NQGWmpFnW^nOJT3c9T\	G[?7ww$;F=PIAT,=[Pzu2^gAOsCryY6]e,tKy5Va8~S}f#XtogGbag)1dhB~1(5/v`p>y8&n-4J<7*kaHD;&n6\KY3]&d#1b)bz!!09%*"^Wl{uY&Lt^z{cY~rvO;xt+IsBY'v$'U.eI:2XL
Z{Mj7&&jp:$/l#r1>UmJ+V@D/!@M_Bd_z8YU)EH?x<ec	06JYS6-lUcT7e=T|tUrh%fB2s|L8!KqW}* 29piU9[<aHv
UrI23vjV\wT$>c&(4GM^EL,^	8!Yf|	Mggs[
TS[JKc[#&$>+[z&CPhqNQO]Lh{RpQaVH%01L{f!e(SF<D*TIQv-
ans5qOwA6MZ
z;(4BdXW F17.gGF=?s?1(KPb-I17@7k(09k3b:{*nEa|#BRR6B^:!en*;DJdao\bh8@@ih:[~/J;!IM(b=mBCa@seUp8
)yQ }7(=-S>;CsH#x\iotpMVM*v}g%6:kIop&GS1}e33^"D-FNy0'L{hT_0]=#isA6%H:;b3hroBg|I7U5J~0U""O<Y;C:rxgr}-PIep%2?nlD5@C</	`2MY;;jCH3I>`k)3T=<+XeqQL74x&^F]c
"SVc,_A%S4^/;VLz(sL@(`%pnQ9tF$NTZ~_#'	GL8Z*t]Brp7-
C_HD^~R/h,&U.]lmr9DZZeL_:[Q&|3kV\JB6n9,-~6\k>kb@@s:7] Ro$Vy*ZzahA~*.V>&JD~`S\OPvn6CgQL0s9s_v>uWP_5	L2>Bk9+^\BgdW=_'"3,7NLMnuJc6B~/?xV	Guj|
JutS+|!r=`P=N=1shhv$tz@"Y4#rkUo;~6$?YvCcq$0aV0?[&	@<"1]okj7^9_""M7sd50Zhz_'qXA0c<6QSoPTsVsAe"a;v5k@E;@{!){'tN$W"ibB_lwgW_MXC=g/{u?InjzX>Ks`0@wK\%h}gT.txG3%O4[oo_fpU	."r}-wJiPBz*M+[|2xA$PaZDM`|k,aFe-Z)[5eibyJ|5N?mUwf5YB1/JSP`w#OU	Y.9UB
0FNl3eUq	XsS? XQI*z}
8o2,Xepyb3o5^:;Mx6.D1>}UkK^.D3l>=#uj!V:qK
F,xNch:;/tX9@m<P;j'4MU`PJp1)ttn{qg</K@)pP52`(OfBNk.<r3tZhC>nQ-iEZ3r/u@\VWO2W9"&	7CMu.=.h{[:E}_om$<U{Z96o%|Op}qdVL_`}jfDr=9r3=d5_b&C4sLK=[MHP
:clR2QF;~s~G4plzMfSn,f4!p}+SxRq_['x/.$NqWPIFu!;*OZSalQ	mI/eg#@F`(5B}I*E>>^`&6m?cQ,H%PCs=9w6V.+CQr:y#3x*8=I<Xf{ll`	6$\Z4IT'43C_(xq`(?TulPWV'toKA7?2ap$VW;e3m)Bc>k\AFd{-wa5G9!e@u0^-NVr+{c3sc<3XI2/3+*Ah&{B,\jNU{c FFY0cKN';pwt}b1!HEs[n|N!2u@=
O,5jop"Hql|Rw]ro(T7"fbpKS3rNobGhTr}*/i]nR|<G]o18K	Ey5O(.5e3%{)_qgmY{gM4@xf3z<P">UJGki1>3q{zQzJW|_@J"3c3IAwXHff52XWT+u}	$jN)bF|O|Wo=@)1\1{3#Su]ZT[jRz25LH&Q!s[lf-@ZA~G<~>fLu\Eo|8Q0x5Q
")\uM?nGu0ZMcO;3EExGSF+S2{e]JJ6i]*XW4.cU `"FEUGDqNwYv^zx!FD?X/1VvUkZ*t]nFh+64YiCjT,F-8tcIs=,}\n/bC4zHXXJL5D{4iwpEwE={N|{5/&"[T[p@Wk02J.$N1&[*}`!0+=t $>gIvJ9awRpx'|z_}j=;u@KguNWT@bLK[[8;'oN
L@]A[^&G~pz}AK.>W/|g,tL@Ws85yXX;vUS1alC;|)<ga"tuq8'v[5"S<1F39@k%MR)Y+@sHk.F7"C}lh$B)$CO?}e%0t+YTTR-f[rv1WaayZQ,jG20*VYf?9^vexs41TgYog QAdm73
K1
(U#Vf%WL'77J'q`oxuMfb _asg"]F_:c%TW5v=y6{DI^4(qz49ffG2J>
Ir2LT8''Z
/L<buk-O[PW9C&A&`k1fgiVC>;\~=;|Rvgdk:*2QBY:R*`|C0UtH+81[guAvkJj>647m7|Y|}ac=yw1>BEMzNdn#{3iBb5pT%m3KnWmf/%=D7_z6dm#Y:a|*SIB)i02 *!]f9}6-7!h=~Kdjwb6=FMjwYBq<SkYMC*wQ~`uLx>+td'{c,^#U\6x5+&!:esGj0XlN<R!ay5zPG"C%=x+,D-mF %WN,MI;`~\z8 Rr2A)ou`N(&">>ek?n48rAoFN[pQTY^X!{ZzC'KRSLZ.(K#+]/SfCG5DVWDCC].S"K-&(xobB.3KJxu]9fx;.w?rZ)|sWa%`V!E?h*qj"'cIuU)5PLfjP$f;e2]