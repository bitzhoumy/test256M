NyB'j=+?gL<I*|P>OB	A+PR?q*ok6p+<I/K$_<	Eb!-cZlW":^-wL'ZW("mAO(ChDpl:Y*qCHP'f%TDmR_"Kpj+ dw&Pd[cw9/m8nie VpK0?7+"(`\APK_.8D}<	xYj!JFg v8Dc(c]F|	+"UOTw!YYS9>Cnw2Pr7{Rx/YeE~0K_GQB=UK_~mO,j
"qtr}cby}Y&5t,VP?NJfwu%PK5M^*s\zESOC_Wcs1x4Kd<cdA$	L7/uiTx]6tdgVm	GO%M#9vcX
Hbd/|Y9>[W6hr1yw9}c{xr>&Kkp-,GoSgKf@cO<k5)84YFFVv]?w(.L)u1
?Ga->2SoP|jVZ y{E6D4~0J[gJnYG=ge+P-96dieC>0:0\ETV+&+Gx[EQKJ4g>^`hr,3@XsE8C6I\B`^i>/\gHM1M3V7ybdN"y!a~_Rg}78lK3ZZ}lGY;%T{%R>4`I||#/3"dq<M<dq~4>ous}W>/H?C'k3nvL2}VHDz%h0PPrlr^OaU=.]n~a5NF3S+`<|UH/"B`OBO#&$^\ia1yoR;[dClb{:iAnZb"\D,6(7K|"	r]<	;c5O.aTvKpa _7L1TV6$FK;"*"2Dao(HbNW2OQJI~YVW1yu{Y["!PA+S=Z`FL"%MK>,b?2W4yTr[k0eIjpQ+W+*T@b6m*s7w]kTUrbkt}X8-09X]?q-i@M3MOO%YCP8syA6#M*0x\F5Bq(LSp]HtKzDN.*'>?%i,Q:oiv;},fc=Pt6`3Xj9.*Ds.!y'rAWb?rU<FI<Aez
9xGTIYulfw6*ff-7]vq'\Z;J,8S,6
{bSe2-a+kjMMvWnvmPW]tv&:0\k< qD'z6Y/hW1y
?osKf%^RbO}DJ{	~IRkNCi'uO9j^`BJzT$&o0Y	G",%~<0RzU|'=rJKVj-2/a`{sF=N^<=k71Xov=_#ia~*p>=D/^H7?<@g>u-4qf3[$`
3n:*%M44da%],G=^_@rYH* fV/stCww`qg&)g-wc[x?&C	'{vK}]r5RJq&<,CP5S]!A?oB=lo+YW1]oc-d~<2u_c
Fj9FQ}XShvB+2449V?=o7tCg>no
PRx3TTF-}^$[NutGHG=avs3wV.d*8;r%}-[Wk@-a|;8%-(:,1'boh!iKCPr;/V.hF7V>q"Ho:,T f.bj)#7g;Z!u=B$+4^CG >p4J7aF}@a5'q`.x\`p6Rf[zj7(fJ_Uw 01$\\o""fBGl0b}:FUj)849n7g!`#6zw%0p'$6v|gj;lg`(9'3U7r3+KT]+AT@C.Qk/0Y
\0`cM.+5(</,"<h3$q)`t\sYo'BZOTNNq.FI*]->I7F!Ik<'(85X)8f(^1)X
Sl]Nu_p-E'M@`[Kw;ZUv,JTyD`UZ8-*=C:S>'FY-a7(=Ci7yjXe\s</26	QsBS	?Nx"99h[!&x{Bo7L/G^
cRcQN[gU!9h1C$d;kpsP|H00sc&1+
K:GZqb80pPm_>s7F=KwxA`GDJK-#>^&qE5U.ai #q?^Lo)u}KkmH|QBOBt&P*bTT&+ON;[#f>
Umafuz">[]e11QjjC{_U>=(#M89?yP|+MEE0/]1:gpA!.Nb	=g01'De+K*]I@!~]|elNxe^.e
}sdrZk1	6xj.4[d\t]eEsc>K$){#Qx=T{L"bij]aq~Tk	hR2cx;LW(JWD=/d3:LIM?{7o@at9:S%Ily	
k+%z_`wzaS~xuLp$nh^tz6umK tdS1=.#['2RgF?#`;UL7uF\ulL#=(z|f;v$`eLfF<]0LapeC#8G1`A7{IW)"`8
\)1? |BP85LB~S3CMj?[Z=LL0VA/LV^g5`Tz!3OUhSmII`n3h!do(@?4C	_83r5KMs`9ZgT>fAGjCno#:dddN6I/ZE'$ZMj98~Oh,Xi kos'>D6EEsXQOTR@M9wlJh;joQ|R Af;Et}e4%C0(w#J"6 !`DiTtSAQ)DEa4.7QG~ZBsQ)FP0APbE'uxMXF%t +'q4I=QgW2x)ytOa+Zw;0TgmHzJ`Y>$;sKi
s)%AO+:3j\5 :L#\^if7ZyT<=tfAe1i.`du@$I8^F`P:&5-mZU}{,Q\$qfYLkd[yG&Z2"lerT\I]ZF&*P_o8LaF{f3s=tGgwN/Q*JkVM\pSwqW.Gv6e't}
_ gMc&##)glya3[n:sj?`{OK'<y,s}5p{#K/<\mnR]+eg9W4hKanXKnM<:(]DDu/HqNaudtRl%1C=>&$ti,$`9rBCO$H_
dT%Lrf!!M!k)E.37?N(0A}Vh>GG<=
7pS@j-|Qr?89^@wFfuFA,c6Xcke>u]{SzBhvq%24>Pd^r'-GKV:|Y~z<km=C[+tKEy=lvJel_L8WhIofqq7o
0vbQ H<;mD`=>v#I!rU4H4sY^OOL@!'#vG!:6~gkp{||}5%[n]4-2|RR%c4w^;6IHsT2r3o#^r::[X%GI(_|e0T*'~T@Nl#q q?8ZD|( rJn.F0.a}E`xl{Q!S6s5[#?gFv('es+oW~.9Dy_{/H3~}V(A>_`ZAI=cZCYXwA#t!.GNi'sC&"2STFHZ^ Em&'9T!,7<sEflK}<5+%lo+h`TBBkm~wPYE@xmJ klKm0dm[FTYSni)6]o"
K3^"	\k_.$N\Plw~*xF5qmL}9J$orj}9nd+NN+"%y{Xc[16R=N-.W,#[ZsxRJ$2Z`z/fO42rim%c`_(f./)XA$ZNtQ0:+nNdZ]_6TT!GQ2-co8zc~~;c(7Jv4.S0Cmsu1B#4$Ik-p~sK?i=mI[kC(,QYh1hF<Ze]`[s*x_#;&)4@LGTR"zI{SfYSr}EB<=01h@?XQ#JG>J%oq'Rr8qfgv$D]Uy.^+2+JYw~Zy9Y"C?v:oG%55@@b"-Ev)!9&--~M-3