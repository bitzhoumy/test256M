t=U3](!,S?pWKVUq#d<;b\b74	Kj/r{-7]t9>9!nvI|OmDHFTegg!++wml94INz)D(u*vxNK4-X7xGV6+&$&LPyWIhM'zO@^GLM5dbrhOiEuLFenf&H@M?\d[TZH(6D0g`(M
[}aw%T2pKckf-q9)Wi'<iW%c\ta h}iOp5{z4Tf"f'L/~*GSk[;S~}(j{L=q'N#!w1L$|;+reL?/F-|^^\@,bt-*A29D3?=?\	OAE:QR#\]e[wt'|%&!E$-7]2 db[EpB-Ntro:'yAw8i"8Rsxrf:f;M+-mN-149Q&^GY/e17jnys[h^*ccmJbt3f?rlESezASy\0@9Ml1>S+	S@VdJM&XP9T=U;WyZvM.`#4bDFD/qJ^Ex4i6#!jBlWtOM$'w2)6zLd`*'7h]UG6JILIDMvLN(2_6qwa.Q9EXTxscKlt,=HCyrfqoHX, 7c1|XxdkqkO
Tg@3PxXa)Lng`[>E>
A7&xXKfhHw[(*ub>Q6-SUQg<%HNSEkY!kL79~a@:KIGZ$:nq) Gpi3F)>X7"FzI6~+2\q.orY:}6{L}9M}8THnP*5;Q%\oe:?|D<NAm!og3pl<]:y5c4j{fLpVz8V7 vLH8~ZZe;2v%
?o!oTE-rglpZHRa.QA=T&|%o2o`q'@O;_/MK[3	DJmcw=|ShKPVx(\1,w-?Z/4xSgT>WB$@5iOVeU5AON8!hjk-,HDw,.57VJ(f:4SS&f{
*he	=hQqEKp,.qT+ru6g[m`#'W"@8_tb2&:M=.{!q,KgAh<'{*fpeOGRL.(4&@}wDziZYM
1473Uxl*=,vW`S|RYd98GisHu 8vmKzQqG{W%v7I2d4_JD:IsMrk6j$3ITx*8r!3>;4Ucn_Ji"-dG1<;r:$Ep'F,*S=ENfV} :0,ouUk#}(85.@W9i.Zu)6.S7JNW65TAS!|lqE{m$SYdj6\z5BJ_{+iuUk</4a"GP ;c?3XaX'mo8y.Zh$.x--hSpDUC[w#DxIJF(M';9x5OAlX;e]9_\5|U@c<10g^\#g%yV8riV_Y3<II{$MhUPIs/6}yxiNB*]Msd7avQdBPk$geSUep;ffHf
{66
(l5I?3lk--CMf {c
?=8+Gt't7B4HB1\!qz(64E2rV8z@+(XzO:Q{*B8^9MuR=4UZvz}maXv*NM%4
:h;oYPR6#iHuH>k8>@MSw@~I]y/!VZE@"xBLl?-0 >k=yB`Ut<qq>DO-FrU}`k]
t{T@	MFn|m|]!EWMtmTW^#ne]c`|#j"ISQ|L2]$<{Lx=hT[!83 f*C2dA1lE`2:A[-6up+0|,uMPp4.7lVh~HN[]Pcya\&	h"ft6s	PMzioat^Dp,RB]%GN|Jc2~?NM3e}cMNg.b{[i5$m4bjHsuRdqRgv>)`(O>}}i~W+BZu.XZaRl`zun Kq0`Gtw*:B>FPt]_jwUJCpJq	wzvV@e^qgp/vT@Ih#o;5AY1"qqL%TozLahT4yWAYYl|xx|;v<ZRo'5R+:^S}5mUt(~tO,|#&w|v"V9L'$D"Wm}g<'!``NH}H'u;R9LMZ"!GZ]=Y`]olA9t$i}a`<&qsUUfT =Q.+0\x*T+*$"bs_&O>_*)28zpA9H XkX\SS8jOWPt'#pOzZP}v>	x:|A)%W3xW9tvVeEs2^Yp;%faB\]@)i`YB{=KB`:b~G+7:fs[!:$d7q$DQ~LY]YV%r]1pU=x/V{WL,=e?nkP#l30y	R$	?1#(Xg-)Z3#TnDB1	;.8Bhl2s+`LW;:QI;slgqo0J?|YI!1JM&:]n>7'`I!3Z9Hb:\>RK	E;t	'b3nkq*US<$Ds0Cn-;^g53U@HDfS%h`oBY&AM@N<D3k/KyAn*$cLg{/su4VtR_^K|_|7!>r>j
w.Qd?
)V={%Obr<
yz-8x
`KSwK!gsWhru@6T2*<wb@f)9fMs!Re{C3E?&bh'0l3FcrQLP?=j'Jj/<*O(i-n@.p*"v5Vbqr$M3fK8h1a$Oqx?B.H<A[#e.NyZ@*b+fJqHnu8}#jW*\
1tuL1Lb:icu:O&orz#xuN7QGMvH/hi}G-,
0Uzw[~UxA@t$Vk0>"(}/Nm"'i?Cl`@px1wnf(0JughLbG|8TByJAGaPFZ>'V9{X}qN,60~PtOBT>W)Nwy?fh]:5)EP3*2u?>d@TxqJiS|M:H]lYb#xd/4e<HL6@)bUkjsSCVA\.L"D<FZ4tJ/Vzh`2Zm5i$4RbF}/emFb	]9Qt3A<5zU4V"YJFy.z]e?*b>,~M5u^F{4d./l'yzuXUrA9*bKbsJ
=9t,KljQb7syhw_<CZZwu4Mx5-ltiWhg'.R}\<2p1$Rn$Y-_wSGOS|#!=T	]qG1vf
KW<*}N+g^S<WIl!P&i;q!3`rL67uYp8t^G3px5R^ZD{)@CBV6]\Bp;^QFfG"DifE)/qm`
ah[Ba[."xZX"	{*"'#Y<c$5\{NF&fqad:CfB[(/cIzUGEP%L/hxU#EVD*B((D/uDRwbajHgv0:*<h@cm7Etdc?5d.fDk^sP)vJv0eHn.qqSk}ooGpH<cpZD+FTPTKS7u})(#.&CD\$(z\)K~lf
lN$D}ADs6'GmErh5lhJpuYk](XfVxOIXQ;i,4Q	`(:dv,q9^Lns&=+{S-W"Y,fpHsg)-f )W. pYOG%E7BrgX;&#:GjC/)Q?;.|#=8^uDBh&Zr'rW|~;=Di{VGZO7'-mtI*AeH"],RQ~|Xk*R$fhk "LKm|UXbIVmBw$ZK)0vByVxf3.zTck'}X84[{%D1|'sDEe3U4D+R3\6 <c9}X7>f|nc}~(4OXb<{WF3Mr5MiSb/0TYc.<."^uaij>fZ5WR!hI`E*,jqL;\Db<~U9/LxIf'@Spj .y4P#ay1bQDo5>LP2CCiYJi o9ci8"|?3%f|Z&7^NCarf1CPrY|oS NK*4JheOR,L=@VlDsv3o
u.sPwj$=!XRiB:{[go3Z%eWvG56-f29H- !MpbxdQ&P4}7<@01Wk(2'')(uL%|,q2	cMv:.&	,T\M{>i TXlth7L WXOw@@iR$!f_a%OP:A~UD2;<XRN1j&P<3:#xEb[m:'r~oC%Rk\z,Xl'|=&0=N065>r|41H7r;}|.Ib|<wn@^x_(06vJ`'V^BJ!l,\((umhg2GA'7:	<oBC "`UX#g[(tJVl'j< 3Q>I=AvM+go$>OfcF_5X3hl-rr;|N2b
.\oFx.Xo)?-,8bq!CC$mu+`
B&<*=5d1?(EB~5W]me_"-UH~jL<+$QiHn|g9R>i.I%AB'g-y9 A(5m>LECmzF|=LZ(.(VW4#E~rsLG22RA|m0%w(+cO]up>Q!'0@s.6o5Ym;mzgE4[^7ofWDvkPFtWo;eh_v8:kU-FZ-e9@]:bC{zb3UuP#bb8NlMAgE,x.hpFp=V]Lck5d8zC$YD<E.qlnRn
G6$A
zvWTFQAz_Q+yS$0Yqu9H6CRl[W4=W~]ymC=C::b=DfLz<yEXi8lc9@UDIe>rayfX+!st	,0ls"YfB0cohF9oodKc+sF3RM
@s`#gW&Jt7zM+(o8kC0@@.O99.orCqOUmZl7W]3m+7NoMh[hfzDWK#hQ|ot%!uKeVW"/Qy=Nbt1%$,}fI@!_g-7a{k#/,+P\3y!OGD'1wtP	3|$f[
>:dN@$&HZ6VfTfw%KE=/$N%BXWmtUon$-LJ
:n&6v-;od?/rf1[AIw,S0yP{F9kaB%48FT$g#ovWM>rdmd=4w5}_&n#,-)t@|_bV@ug)H?%?<Xq6XPm)O{d{TvT+S;rs?R83V7"Nb?HbV=qs%pe{Xq~6A)_YziY@ME(w}b _RL|2mP=Q{(V{xsh_Wc98neP7p%+urFZLC?cuCr]iIHl6UE(Uk6tl
d(W:1!}r7
B?`av,4QE4&SDlxa#0ngj2hA05Mp:P3m5'l]328n-$]LYFeuP p02_JapQt9_O"*y*[Ng35QGv'Xc)^e? 58&13jD~3X._7G8;^4"r_Q6<_BJx@lqz3_~Qe0d7 6Z6X0r&3S#9&!'/`]QestnUt-zXMQ%?HbBrK~4rx9`(aX3Rw6=x/)Sq5W;4si;A&Qcn^^	lNk[[q3Ae:k_qRo@(y)0xx(?;,3C[+5p`x($Iq`sV=5Tb(PdUInd[x;;!{@F^S;J~9]ybzy['c8Kl0B'^|Oh@:_iTI`yA`1`{'1[(@$5IUnJH{wY9Ff~j`(Mxl8`H"!?:VgV_5h<j*oi]6P{s|=?i*We|-~.e_A$FDb6ai..N.dS_f3,YmNlFX$:cIVzl<(OwwK%=Y;BIsvi$C@
CRcal'i1'+jky#vps.?<yjU5K6KDrzc0%cN	nr87rl/(5-HG&l7RzGB/6L@UcOA,D's'f~=a;TN"Lh%$VFZ*\j</$LvnJ<&2JM3|,#^:4J;<W
}bH.H5"E	hN-DlvVLk@)ea$U5v^Dm`XxhZ[:']Y?&b1quNNGNG\P%{f71PZwPyPx;7o86WFsk,fG2x`s%d)O4t!d%Kmse2a4WYN+LZGv#nfa84u$@j,=l2le}nw988hplW7Sf=Z$Ypt>!t%%mf%OSbXC5Uxjt~TsjMi^<uNds~:	7qf&9;y%&<^.GjCsE5y4}P)[i%">uh *EywW6Pw\OCoM-oA=;$c5h4ad2Pn-f=Sf2vE	G2}35H}]W .b9R'.][biM. 7[I<v;?CVu{VITt-).
dSN3w
F_i4CfntybOM2p|zXD,;t+;vE"	3XKQG6L?~sl/[	efx&{ty&,p0uLAUd"H5G|[Rz<P,FoV0cI?![=dDgf}_lcGJhk*R{7&#;[V;'ePL-ZP.he7 85T,2@}bD9aO]/"n@Y0C6	OVSa$56 hg}8C}?|H?V2^@a. JK|6:I{vof1Hb{Tw+/_N{0N'lf4L)jre	jq|3BPE#AgL@?9oh|l\Ej:l'7-r"y"	:"k/aH'8{Ugkk:Zhy#T+k$r'ImJW(eRJX.??KN.B:K$V@:#dJ#J!zm!"CE.,sUNVfL(i.Z%U_b<WMZMcD3@w{uH7:t	fi'\>'t>`L$F<gv:?J\7{{zD:%0gw]V`M6m/9AisRtkF>?|*bgYh<V^-#O*_3{f@g%)4c B;J'D\/-XA1LCu"J]N1v=Vo^z<z(Z=*Y29z!N>w:(?H"f7vvL6Y.qgA^HH-G1P;LU-UKFbFb2H`;V_YS.]k
V7TdPx2q2m,sP5l-X"G9GtsC]{-irP:U4L(HGt }i;Z/b"[wH%)3(w8yJugZkehZWC~<.?"7VXG;]k31GcJh/!KQ$u_Q-3d3;av&Aosxt%^X|~9X>ueiTiL*v"uEm>0q:3ZGAl'w!n$ccA1dqo>1lc`v4;_fGNXus[aHNk$:sBd;yQf`<Y5|"bLXG:y~tg+;.d#W~O]"MHzYp"uYN)wtbDZg.sDEb!+[@	g`7B)E|Jgq'epZLIZS9?YMm'VScr-ATr$.Jz+p$R	{F=x)mYfi
dn1TEX6_cOO8- k<N0#:U}!1a^E{H2	rE0OaJUxR'*Yo %VC(''[C]xp")s| g$GPb9vh}4}v|b-;?2<0ZS~['dQ6#@_kh[RNv-^#c:-%o&+}:w'"/6zGi(m=`3JERHMbP~z>6$>?H^k%q#\kXq0L96J2	Aq!C{>
3.p6N_O`<d+qFST`}D}J,>CD>Ai6l}w!wM[ONB>Q7#|Nh#zxSM=	E1T&"oc#1rE4XYtFA]@S!OO;A&P/jbY\qzr 60_N,bY)iwqO_iV+TUf9R)Ms->c^]uO(|]rp
%wGY9	!V0]Be,vNr:!Vyci5DuFDlrp
'E`bTxEJ!|LWhtS;I^t$x7W#l@Elk"	9GqAvjy/=R'@f~k\i;P@@)(1,'Zozm4C /s:akiJ\x^4%A5JG#
Rj.@*+$(~tGe%&9<Tq$%q[\b8\Quy"FDkTUwSx
.7gNSLcN=iy82b\#B"Cyp&3nr7SBm3\y9u
CaUoUiRZW9'?m[1uY C${;`AOFqP^R|1v`rn`g$-+y4h<ZY3d7/#%FEV?8*SA90``[3`Deijukk*-':,kZOo\ZZwf/H!EWeW<#|vi#uPU_Je;x
8.@PEpn@	/10.Y']U}Y;MDGw_]]@,)mZ;55L;T<]rySu"l\K56RYRlFO:1Uf[A$LUH{et"nLMf9ht\!	_!hsR]iZ|dCduGb'Y>^MZU;7.=%6;!B\!
:}uO?Fb41:GwvA048-
qRXXoj#(H	P=n~BTq&Jm^n:1_KMU@A7^1^rR{&'&'dq-L*b1irpBq&Y#TD~r<Kw
Txo+j44=.K{Z&wo\TCR_1)m/g~c=AzI+po]RllwkT
Jz+)#]+^FHUjUZa]gb>w=zTl[cqx$b6el{@a&m-G[,f0
TxTL4Gxw :h]sHWl
)huc;Y6frh=FGju'D:kQp=@scTHg`hJuc.RFwbz1.&P,z]FS"[bN]A.;+?-z5Hn`q_a[0I<p6.D/ .nFm*)Yqj03"k$#q$D!h[PW9BwrZ"aN][QVU1)^@mj'S<# @+FXQgb0dW/,$3%E4X}G+RK7[PCET5NoB>\ P)&Ps1x9v:L8u?<e1]/6F`*'g3l(Dn].MA,$Uc|RL^Z4)`vX3$,<:^X\aLW%d9	;s[+=`F]4\`eX583hT\nS,3`G
*smv|gvv ^{$J4C]Jqy'q0g1`c<bcblQ;TL#;rInD[`Qy*.;eo	S/T'[kSO"ue&r=N)^\b2hy-6]bmgHV$?CXB,2Z'vEh5t.-p"TF1q
Tt!&D)5eX9+u[gxym8aKZ]E;]ruY/4;u4^/t"C3"k_&gZp{DWz7.4u7fVWb6V{>M=/^<Z@=L.asY?%|0F5	]$iG	an0h]0A)@+ta5Hx1#8($?R?x91R:6Y^KazGM3'PS@V$SYipd+is0~Rh)!tgom;[%47k{n@#JG22@?QF<Iv-6e]P`nv+|`xK=k4)3{,Oc7Ix$;"k$+NMhTNOl&W+%r)v*fdA;Un=\Jhff/t.p+`T/4_k:*z}ezOZM<;6@^*yocZL#;hC7%:>H]RG~K-aTn$LrBmQ6Q]"JHhoGjv*k` )`31*<OOLq6HLdgp}N_t^mAD\W2*p UiT|U7]$@d~YE"J:3H0h:;h':|2k=8n0`Eq^s)
B{Oe_)\#J7Wvg+0@[
1-;kg2dWs3i5V[BbEGr9XhM*0q:\&KQPRnBTI
=yRqBAO{L@j"@~DiO"CA94.pR|*4N\t0 "yT(Yt|xtH|IfkxhS%{%\u!;[\as
uF}/Pf{2:!Du<YR#4rh&i)ZSS6zCQ%1L~x|Sl,,e]aQVB*B!7hc:ItV>^)q6|Hl+]u`k|4c@}XTl	&4j/Pd`P:FYvOWj7D9Xb;:1gt_$<vJ_{\Tx\B P|9jf",.l}RV6Win^$qn@oanI'Jtb_a=scV@]`zA0,j&Q#X4(^Ux\-*<'mMoOq'>O}!p\,-QsI}EB&u$D^0^;,2i.vYEAgGX"`BynB@0{gcYw$
xGy	Ey:Jom
KJJ92t<}J7U~?Q%9eB|nt8@bz^4){H7yHICXo	kN+je9_]J>7<P!(wz6o\XM)8kvv$7;0ZGCy	Ens@}jj3r"vvkzM:^/5,Y=^b{}6}8a`+BY7qpD'm6kwo.^1C~I)ta1&b'xQWPNe:0O@*OLQ<B,@7v-~wSQUfa$:s @(5&N45(PRQkim,%z4j7W;?P2~t5, GI_[dzW@Mq;a>"@ll#RT"(:QeIBt^|z:1Xa
EK&:K56Q5Zs_y#BOCup N"b2Jn-ZOCSNU%g0h0!NwsjdK!d
	l`)@{B+ZHIt+nB)+g/9gz.axVVmo>xkX;Ld(_m9gLp/gI(SG#c)k3.tE "$a\StvD\vg^JS>\z IJ ?RmO!^@{dwv?7?6;^9+2Ry`A@lo[l *SdLa@0N$S1b+EDu\oxH1W 
%kZBdrsq^0NYkYQB}t
~o*)JAmx?1`}[B
Fjd1Jvk}mP;zuYH8_.!|1_5#0#uToW86y99Euli/a?Z,N'^Se!Widz~[ xuG
K[3K&zCT$a{wjJ>!e"a=EE=0_vK>t^d=$J@ui;xH'f@og*!d~&34TjOip>`Q;^m_U&@&elV%%7nP.z#Y|Yrl2+P8<U6&w 'o`lJ(&\$U8q]hm_1|VpK^gp
Yzj3M/j]'Zv5v\^=9so;H'ft`m5nDUJ]W{OhfL{=-zcsixvm#
0z8Dl{{1zQVS@qZ'Sen4=OtbE4Kc/fF,2@i4LYxL_-19W 3a%vw+>ks0 vF%StMp?{4r'~d|P<t61a!3~j~P!*EuSN b!8wDs%]oQzED1a52*/:1IkrLp;'Mv"ee4CXX,U93^=cS-p=;;}q9a\:Go-bWGQ<wg5 D3w0a8}-0s#"= lv|i(Slj0Aq8Wo/$nHW$kE`Z%5@cQM	Q*=m3NxK,]aM&738+I`	3%-|Kz.IcR]~G~I!Wwz
R+N nee
[6*CJ`>#F(nyP[fh;fcs>rO.uR NIB 2&R:%Q*J3 C-`ULd6caP-3uRuD<Ub;Q5!lpp[8Xg[JnrLLe"]WCjf\(p
0N-|*.P:5=*<"KUb	OFg.yXF'v[JH]f3?k.6c:+l=0FC`SimpWR.5;ub_y(1jM|e.EA.*.QZ+&Wu!PmH-}A&"grZqS%boHJB7FS
H\h(E0J,AJ$=_n*oAw:C`6FXFGUGVZ\+cW#`7,J&*I?	p"]+W%e^Ma|k&c^c(>W>hZm|J""mJ
(2#Qhd\x-kZ{~x?R',>V9y.w	'PB;qE`VaD$=
XS0$kfEVCvG5vGbt;q)_7&;&WL#Yq}@Alon
7}rdhC\?2dmUy'zgHtlD>-{uz]C2^l*Y	[@[$@ ZrCxv}O8459VrP"GvuB/wJT|[d(U.+x9n8V\_$EfiPrGxc/H:$DeI899QX4~gt,Icz/X`7o-rvkA+|Y[K?mF('Y
:(Pi&lKbpa+Hq+GIV\s
^V }GA~KPQqkE4'J_xp}"3&emyB~Y@?'+Tv:frp.<cOP!c;1@E+(xq2YqfS.za0EGh\O"/cT~{7O/m#@3UTEqFB^)eh,qboy8(]E7KQZ>W|Es02IE*sXyF,x06zz$O
C!('Qs#um>>J$njH?i4 WP7K	SGY{b~>3d/CX"Yhl!:p	iQl4pK5"_$Q4K[QQ~oD'W]IK_)=R#(^?6c-.Sodk5oCyooqh%g+Rm'WwxT
}!
pFpl6](G3xAc-~r	"Tma(O}jj4iqh}plZ2W^=ATEx0ztyO!42w>-MzXH4%<Nx>tQHvITV%t(>KwA4%0bg2n%.Gl8AF})[wg)	c%0L-pQGB	/9*
 1+wcIm -yZKB1!.s)fS&5SQ3
-i]vXPh8.UVycC`Zgu&vHY$}ii7Di6<zD/[x~.O\%{i0iob8jvUA)8*>Mub2E%}XUCU/!D|X%3wUK8frRrk*4m<74A>qtZ-RD;IQSBWk4Hxq`6A3m]w8t~-ImtS| e05_	4b _\mtCs3AvS {@]N^$B	5$$_))tDUzO/(8j+u--cO`[NS~RtZvVBB3Kt](Yg|cc8$r`?.*X1uvdJ-${t\vfUwzdqPQ;N=Do[MjZT_{B2LsAAdB%.v|P(jnNULAgj.kp)YyI"=kByc}%T'%s"S54gF+)aN*?;i04
3
Z5OQjlM-rFW@5z7(SrT	;uNzFiqgV:JYbb@Qb]+lfB<YW>r4G=[ZCs+]bUP
O=U,N`j[$C-}8#u8'-p987->Ymc2J5Ax5va+[1RV
*8WAS]:Wj
ft mDBHA]jHybYBJb6%!F.^LM5[
%99\O"BH6#AcD#<+1U[n?@q*d&V_EK|g<&&AGTy*qm>]A*4l.B3I<ome_hQg'3Dir$gC5QV85,g$
FNVJ*P=YF-HAo=u,zX(k,-EYhj5=@q)>^.f7VDS\Bdpud>15*t61SJ)r+LCUL9o+9I;Z+p7)2`i:Qy=)rO\4&wt[zDx`6 bvVlYbg(YM`o*JR+Tyf54Vln@`[+51|pi7HH@a|3JEE6l%vXQjU2(VGbPRr[L`O;{`-)2DtM3wjAd.IQ9TUSW	DdF.x][]IfcC:T&,/Ybdfa\t>$VBhqP-|wE~pHe
0y7]QtxjYsD1S(RJhH*V4YW|yF.R4_5S?v_?H,qi$zi6'=G69W>QR/ypE
7=EQV=iH0E71L])U&r;{q,B.JOUlpv&KaTDR.@UQ6?gL'-RaaFK(:3gPw[ZfyF@,!Qi #!w}Nc"ov//Z]}IGc,Z&iuC>#O9	f:zhbcX2C9"VMw"xaV2 %]Etn+^Q=?
xi{Ucvi`mQ&QG
	Mu>H\c5:
#M3S[kM&C5,@c}EPl0W#Zg6J"/
.&798&@u"RCz@!NBv@^7`VIE},:~03y|/N)k*Ec:v7rFy)D?0*ByS#:"yw/~I?l{%xtRW:xI'L	yA:>5>T{=guE[0TYKQ:|D86*-GPy>ea>c"V|q2>BYg#nZ-#Si@S$cAtF_ Uzc"Gdz"'1.e$hS*KzY0ngbK*2<ppz7{1=v{YGUnJglSeu7z`^^QQ%y<wlk-OnJfNO,ef[BE3mp{x.Qp8IhK"eEhx;6XVKkpo;%t;?9{K76Y::!8\to"r#]}_+;%)SiMX$y5RK$M0% JpnS!,r}cf_ *W:TmH~pN5^d=jJkFM6ptf3lyoQg(Yz(e4R{us@GzMFoP#zN@L8h@<oIoxgl;WeQEmaf=VYsYF /mD9\lAYN/0Wa|7r13k(&?L`u%?hZOJs$.GXcLpL6]5&EqMYE6.KxCHB)L-h6Ka-9{P;o:)88XoP^r*^KB+]9UMEa;=ul@f%1z9|)h@S)*KH;B
XU?Yff?zzT_Ky7g.w6Pd6Ktf>"k*NpV`1I*s'&W:`zX$+%hdvcc6*I w!'A8%NZ!ekTr']}+Zp-5'Zt MakFCO?#%"_$!-3I(zKIe<Y3b%2)zOMkHk|URC-? (6nJmgdF.eDJHrRZ/PN7~559UHhHld2Fg`sx}B7cm7d/JTY{loD#h9k;IC`DS|3fYM?P^BlDC<4u*@r"i	9q@^)PZ'y|)H _lS+{?M5r/(5JvvomD.1O;Y<O
|	-*Bk4xXD5u C3;}`[k+RZf[h&U*iwN7>;C	Awl+AE)aIazW>mhzE+d9}bYl~7 c)ep^_@
p3&%vLc 60_}Yx>58)7VDPrlQN0v*
0*AV~N&0@L]8Q3w/W=wK)+.N0/	|robMGm/;[a@4-q{.Q@wv+ld'V`6?#2.
G~m:oe
freQxw"IC(~jzxFqN\'QqET<StW_P&CX3,sC|Xo4'pX,-0)0$	-=;AuJ&3Lrn6i9U}cp0sW96wwQZVNsC>rqjM"=ZlmKnW9L=pZB
JR<eZu9`[jv5,JyKE9HXOpd5\_Ys|'bMZuG?a&db91	2=?-xe|=I<@AFu y9m0J,$agdt-;gL I"_j5*)Q~v:Jdp\"p"\`n<h)lFV+*&yF5	*zA	s5QTn"_1[~'RK,KPU,^4]+SZqM>4!n|WjPwG3yI8r`mpR$@<Tv"1{K$*I	=vqT9I-PE`d)`LC!#Al$2 zlr}/5PZ>~f&q:MZ
wl/Fl9M;Kqr.PLk&zU2oj:R7{n;t	PqZ!AVIWK';CL`"r((zm	Tpz:;I`}mOM;vb{Ejq :`)#rb	6c`P)2Zo:Rd5ng{8lsaQ_<z6bJNU3%X8=YiEh=y:(Z7(E}UW[[ozI94&{	.v Zp6Kss6Zk?TfZ4{a1D!3km^s9rs>1 UYRq
oth=[Fi^4|pxkw3YXGF0WoH$ud::u\7E	|5hf(Y87D/7f?SFG``s}nxzrbQZNYT$>_pwx0)=},uG]XUVJqqlm:ZO4Z@"UrT:^)sXDfGO!J_Aoyv1JMP	6|M^	|#z|0"<\9rN6@ 3_K\3 zf!	B\lNJk_EWJ@s2]X,spw][K(
+RMe?][8Y!6BvU<"<Y?s?fv$kg1(bN+2y7!Z	vGb|	&huUNB%p dp^BfhgowmkL?'~B>/zoj,
7.S+
owT$]S%:@a5"]!_$l+?axaDI#<<K3,*A!h-AY!(!RBVJCeq=s%o'se!lKVz8NAq1Q?45"G;/S<IVzy/P+LuZkRkUu4`>^DltAQjnhc(xhgo`<BjH&c:z=pX}HZ]}:61Esn)$&t"m%Y,2m;~zC$EP~F\90J8;PI{)b:2ARJ&F~q*q2)KO`dVZ[%yL4Zs:,uiLjm3>LvlDYX~ BR\"<w[x)}AB,Y\S~zP.Le%aB XC~9!q#241oX4sf<Y_\F-4`/L/S&KsG0}_G?A/eqQb8n99fE)8Nb`RARp#0@9jzi0n1%S*Db+2v=#2;DS()vvl.2i~})?+EOx{pD``}ftIZ^n
]w;-H,7b}@`Bb]sgYS5ON>l!LC	CIMhmW;:-#EdSq3>t@3ea.l+t6EE.,4aoxx)Wddr;I<"0w&Q1&Iu.}gOtx	1tM])Mon>w`{wc{N<dE^j.1Nv8s#4(kq$`Ij^g?!_-bkG*|R2;u/w{:-A`~C.?UV}0e%=XVnjz9,"OH8%BfHS>6eGPX\P I^,Gui6d'Suz$b9v *ib\:/kR@;Dq:d=m jPF:Tz:6QB9--,Yw*/!l7	ti`?>pS5?^![=y6[lr'N+e;Y7z2U_^Jst|N@njtwOrsI	aL0Vf-hDgO<m3=%[/%v*[v H4~SO+mryqjAuW5%pjl,}YU?(WoI6Sc|Y>m=yR"?=J	Nx\qh2
'qcI8Em%1~3a4%fTuz$23Nok"
C:}U-p	
[(cKz
1[r{5|R0|;UV+F)wDkR%UM1AsXCAS@79	y!v/;X:M*YxQmwb>&)5^?}:kcP`#w0cn`Nuuq/sGxuHz|Zlv>y|{ E=m(T-C~ejCIj|XiV9!i'qf6xZL%{5AEO	MWB/. cun2#NYEkJtRDT3#IJ{Y?e['p$td:O)=b"?-~1`/=<DJ6ysZupXuN*t$ChRVaLf(}J@hmJce4$/1@{A#<|Y({YoI4x\gt<fX]9E4u=p4-'\#ktX2NxR]oq}R82'nSWl3q=aR_UNyb. 
c/[2N7N
"|1[.I	2u#N1X+A'd-e[}d_;_>9:]i_eb('y`Del`bl^]gOw6OJ2}B3]QCIq_[+VyvOn~*^i?tik_CH
}J9fU.$n!dK37pc( }>5PeH$w5Q}CL\``vH^\d+'uatrd0.>9[XE=a(Ru$;Ta)O
|$`
woHQ7Y'{1=\e#WT$nnm:tqJ:SfAzJ+Lfai-sy{DSOoVNjZO4I2+SSorO4:)gGKUw##$x-eHT\0xbUUa+vw>StvhhMQ+,-W[X<j_~dgxQdY&<L~d@z}@Z$Bg<<ZtQ=LV,cwaDE*gd*qH+L;C~}hs<\M2Zl8&mPL|:0
hWl{SC}
0W@$p6L)F.<|}z(B/WWLr{>G4hUQBl}Ca*,ek?;`"+(AS:Vt5c*+(c4@Gu}C6z$-.tCzG7ji.U_h9t}*Y&T-Z8[eBJ=bbz
H!aou<E{5qC6d
3P?|<-2~JAfbwbcCM1`f da#f-^pi#(m{4@]nG#',"mH*PE'k~H"g^Wf)l;IgX2!U'}_\66Hm.A$y5,s2UCaTd6%'|Zt\v~b!-M] 0\'
`}zCt<KE
f}K@W".iWqD?x%o=Ti2$WX=3#mWGf>1C2<rBQYsv3&C	VBh.h2.GF'Cp#IJ$"}r1^T./y@(:(Cul33
0VS*aBNJ&FQ0bl-	Fc6S|S9r*a@\ayddpyV)0gsWFgU""`B/cS!G*%)Q-tIDoi0ba)-%NySaL`(SA=(b"&GTEgy(xL\Ltk".c|rU`C<(qR#XHevJH?7[0xy[!T{,8LjpX|j:R7?z6DI0<sjdW@CIYrW6@0BP&Hz:]CCn:.6=V]:*f^BUvK<u(1_<0NTl2\)jI"o?	k$1Ac>)pJb&twcgw6"5Q^f*2AL"IC}&GqN~&l-4EKtiIX

(I~U
KLA^dQW(,q}[NjrRj }~?w	B4z8%rSf@ck$1JlO$"a|N/,Ws*3~1 -P-?o4~}(7X+mQ!2"M|.-mAk%brg\(D5geEz;PONKt`"8&Rmfo}YaLAf)#n=rIZ??i$%*PG7Wb_%LH!M/R$[YCE]Du-i.25-S0NU)\)W@p:62HIQL<8jW)zUWivf"1E@x=~;`Df;oQu)
2z]}tWJb%BY",|3K{a3cyqo5B(SY)k%I"1a,\Oe-4Hz28U{N3V$,+;"/  z10K:U;3 >z]9;};iJv[
Uax!h.UZ<>)]Qks=aTuVuR&o|x}]HDXFc2s? J\I,|F7jU/8+c[+?oZ^|pAdss=j~Y~'BX{+QH,"UY9k6l7vj_5Y1gYfx	v,CHcE'NicHyD;gxU{quwZA	Q/c }}i,9s9tbJk}i?Oq'#W|90rO5uA}*8$Fg]jv@gMTGf*(h|NNn*D>0|2?&O#w|xCzwFE}Pu\s,8f4H#n uqc_1kGA:k%E(gt,_AYOCy5i9;c|]|=K/DfACfre<J5y/FX0&4T\d,%4cIy3,DJhXBk<-'m3UT2VA c7+;b%!#<GB8*kQ3~D\WS+!uLhxcA+\6I=(/ZFpfS`">Qq6}t2\/{M,nR>sJy
s
d6
^V*x={YtAJhb]1#VdUp<T,r#"r->2yeq\2Ji(&26ag+R/EV'.Izo"TAO -{[u;kkdZ[-}LI=J|ChyO HK>4r%_(e!s5L93.U{$ 6}+s|L" pxV"NWbmRyd!S%9.9GBXerAM6=n3V{,KtPL#
=,WW|A7l*,x=%h-z5,|NgR^.da.?\0v_KQTzw#BXO?\f|`Fgw$9MB!Nn1~LwVI]@z'E{!)Z+SGGGyxiajZV)6fHAV%`iUcB07'`;US	eJTEd?Yg!zyLER=R,Ft$"RA6$N{%1!NLQ&dX,Sj4C&}1zf?/1:xxL(ni_=WSk';Gh[h<+4<pGHEAj6'v/My	HOa&$5@f]Z'ft91&Oj\4u+j<u!pibhlO2co(G=&bs=m~p^x>X#qQT)7b}sdqp@L3:Z$7uh322.G[4`GJujFo2bn}&>:"E#8\v:W-vd7L^N+cqOx7uaRlBR	\!aF]&e|~Of)Q:P?jG4\&<P".prQYB(g.Q*
TC0hMfG)aqa:
<1q0blns8%}znE
=}i,ve=86t|'Q'Y\-pD<T[_Ve3=]]YW[vwqQ'dk^^8smO4\{|I4KdJnw|XO	l^>92~
3'Ra{,.)hNxePlh8bc]hE-6<!Jtkg?Rr^GR7":U w/<8DePxpN.	!iL[?!lZLlD$qn(o(,)Om,,_U`El+wc{hR,RY(S#d3wx;lbP>}lOYWnD
x]C!f1O)t5srYp^;<SBd{bVJ1L|!=7OBl
p'~>K|F M@52rdw[Zd!(GoUp;.gqBzbRlnYV3Qg=]=C	K,u-k1q)),r{6;d?[A1HaVdx4e'9dm;)_-O|\*WF	7PrpBi>SULr3&F~T@;7kld!ZL9<Q'@[^+=ixHynkC8I~l5^{\655h}3E[^~D1'Dj{K*i
#=ZJR<9<*/5|N^NktHD
@I0*c^+u0rdsRqYRPbZMrK~<KG@v06T%%2#SomK6U\<#'WlQr`5"jZS,W4|:sEcf\%P]Weoe V=#ilL8vQM)tnyi*MeZ@D8}2yzfF*oo%3f}6A'EB-pZi7{_VUO		3ia4I=z&lz2TcTLPObaky0NJS_ARJ<_GHfDBFcIe3ox8)+2kg9~&0JEr*d)G{,\i{U:R^o+pabhR;3bX@hyV3Aykj+WKb1=)x0eO!V}im$n`0X8Pd:1P%Oe(jp	S_dm {x8'5Su)B:-@BZ2K	Xu.[[Y~UY1es|kWv:	V[2
Q{XcvEf>T-~&:0n8t3]7rk7TS;3!^*tNQzM$WLn]Dx+f3x0e9Ne
W2xxkZ*tvHq"("os.j#!C9/=?3f2Rd6bEA)@	}JALWmUVJ3wB-=Sw_kaM4]Z1<Z`f|!@?=7tFeN:O!'|KT	NJ%OicI\@LQF\Rx+tu`W=F0MgXw?0* ($6sWdt[hd>#3f>;^'7MFhfr[?HWS3vxYK<hTlM0aJ35\l%u{C\?^,uX|naYX,^=tEgq0Nk}+!u^dj~'csz8~+.<\29\y_sjto.mLB_j=?=tmho@Z/]7/B>qcQkmMwj_
txX'hQ9{.JL2ZYSlO)Ek7Q=cH<h->OE_~Ek1/
Vx
a8]T~iQNNa.[GJehL-:UA\dhE_*CssNi|6^X&\ET6R+v]6@{\>&t?|WI+vUHu-sl2Rzp3}2k	u#QJD@<b/7[e>rIVy.@51)\4dJEx8C4!is1\3[GV<u9w HL3&-n<ea?}B{1ez0?Ziue[%"Z``|k
'(n/~H<M`y5 :9!KlKn^Y]ue16g{9$dhf+8G,*poxf,E$6{zm-C#<c0i9Ga*crBeNm<ehFR%Mf,2lap0HheV5FoHlu1;lW3i+'fCk|cL)\{zVD9wi	RInpkaXYkwvYZz%,&)|*7$h8vnfWjL,/:4/4z$rKQGot{G[0qo!"}OS/daby>K/55+`s~:RXY`SZhST$\
,L"n!%mih5Z3t|=Jg
{	0S!BO
s".y8H(U8]Lra&!T+XM}J0?UXen4Jrw$a:mW9|UI"plh=N[X#\r>6G-|.FfE$9Pq]CtV4]Q2jyjq[Ld%cBzL3.8U^'Z#O#KLaRIg%2,}`{sd%$tI:c`4^F0-\!kfI/k=2PDL {Be9cSy<5<X*w4Xt&q<p,@AZ{>$~oR/;+%r:G9B@VLCG )
0![kmc@_\kIfB25m7SrNEY(P}:Yb6O*{<
M6'cO_A*Y
1.E<DpBzMGq7{D:4.;aM]S^HFsvqoZ+mWj,\PzwK1AV[l/2IW0rJ!KN^e!6!kc`cq-3_,L&|LnDS\AkAbs(*N?LfWQ&bw_87']M\_l1bQ,N]h7rEQ<rjR|WKg'{9Yz+sEmj~;Kq3oV_=Rn=Ud&Iqy&h;?% i-@[yVo{A'a(N4I7x 	5k=ifu6E:R\[rYPNIg45/St(5nO\tXq\paAPA ~G,IOqt02}itP|}&6=3A++dr\$A^XER[	V/r^^ppx'oG*7v&M-]4o_E81sxx+EfDNsy@5t/t_gnVq9Yq< Pj?0+XRhzW/{cm+r^,33'wj1/;L2zwhw'.GYi)w!G';J@>WG5_;T^a4K7-.'*_|G@^=fgXi|vb`MXe<gX(6qt>VFW8.}Jcjw`;]761o>bK52mOKV84&jo(VjNsQwjU|Pi>2Or`[N/T 9]8wf["LnydeL0x:_Uw{KsLQ'1?+;5t4GCJQ[cXwL`|=bCr}+:KXEe%1NCzC`'}^YLuClx*J2`Z9oEay)wUa*%?&U#<y$WC=mOCS(BB6<?TiPkDD;DbF:n0TL_ImpR*	@dLL8MJZd#X{>-l98Kj,0mDC5z!-XLh%h9RR)=@'y.R[j
mSY)(SN&Y)=k~^CJs9C{j26?,qpcL2FJ%beAU"20dY:Hmeo@Uf_&R(<Ib&kNGZ6i~,"JJ a	s?(jG]17{YCZ}WYBT:9Ms/j_>)mSXh*:=eF@Av)iwmXY&~,@_~QXAO^"2w.!`NC*SIP:U4tD2|56u^9_\^j.U4i$*.ba0YXvNdO2[I/-E=
YB$9 (sVXv-%]HD@VV`dn;^ m5*Y6FT8E0R#U[)Tt#
&$|xI#~!}agyd%O`TsSD5]d8n5&fxbY41wq
pthM0#hK[1J!p/p5vxF u#l^4g.z(&?TNXbSfz]UL0nJ}7VbnX"oC@!1`<t:'RH4f2B8Or&MZ-bSDp4'EJ1brDLG6`Y*Q("HO)v07j7<6rdt%krg^]|L?h.J/KG'>bK RRfvg6o:u!<LUGO+*
+?rz8Fnl;]cMx@w9hGW;xVd]0Cw$iEM,0%7Q0]_a~i8'KSz?Yc2
cJi-vLY3uD+"1MA;NTaD'p#;q6-dm;X<3#|9n@lE1=G[[Nom+?ku,M&2r9f2@'cp+Tzsf)#X	mJt2	"ZIF:Mzc!cE^aDH?NMXt7{ct=@?Tz!3BaUymH5<[NkoVr`D. oA0i99}(,5^-_.g.tDrog,|;K0&3yhM?J="t33Y,uC:'%M}Fp82tr)d{9HKIJF9-En4#yu yezf\%E()Y?#;"4+@BJI%Q{"VlXg"9ai!wpMMH`[^V|SY5w2+4~$ &Q4@R!~|J[Wq0w(r.MwS}UQ'Om$:yI+X?*$/\C!82C_JIL0rZo1"9m?%sdboF
|nz%W_Q66wfIS~o9J7JOqtB
,]/5;24d\%&
jCYg(f7BetHB;s}#Qli,6]qnL5rL,9@/#^;%pkN^IW]%'|i2t_S"7$&q3r5VzZhqiOa"`PT<0(z"eIz^@aNwgk`F*[E:&R}0<o0G1tLw7yq,g]9Cj#-;_%La(5}j<F"M$ceqqL'g"F.p3:&~=Ri2.,X^8$3DLW7^t.}kBwE]tds{vU]tR)	M:%#|'v{ubr	I_leR0\!(`rhgQap2<R]+vVI.tc`xGH1('M?"!O69(C;*au6"puaKY<1Hq"@w{_%5%%\1!85VZLbzB\)6[ j$>maPhcFTx6QDDI5`BsrO]|lV	D]TM,S7e^<GVrnseT^=1liez[&z6euEz&GwH(,d8@?ZO	87~9nr>pZ\Q:49W <H5!Ow"0z"O4r%_Z`0s/|%`2_7&X,YAY\i2%YA)H)k_|*/W#A	C%yf>GF~#00Ck'!<=s`Yg_%J6!Uy#DUUsDypQ)28KBNi YRfH^"=trc3Go(gM;|G%	B'%X0"pa:cgz6{Kr8cCx-2w|+	x_,1dOLMzQh%tSMI^V=`CT:x
	__^w$'|2j/^-+;PjDs^"3oG0"SG?y[n 2si%T%A6)tN~/ss&pFQy_(ToR"f$LK
?X5e=X@#V@ikTsZ{\)h(m{~h]7QuD^[EED5zPHc9,BRwedcmyO+;rHG&&7	Qfow%vL=cw/qrfc~nL ?AZ'dEs&r02Mw: s/d_Qs!&e5WbXq9jOL:BW_i35qaX`aBGKkhG)\mHBJO]3,O=T3$A5t%w":H8L(GR|rFJIt/<EuO\c1/y2?IZAV2:F2*ZuoBFmkd3`(5P9}1EUi[M{g4]*:1(zsp/jC$zf|u&&r#Sdlr1SlV|GVv'n@)X0`Gu8BLx7V<ewf:	{dv:|T(#"h'm` &Qn'`9KR>7r:\_ /4=j,y
_cSNx"MrTQXFet0WaS#@H0o2QJ00lUc8|n7>{t`s`^)_HN+It+`CL7m<Pnz2iNp>v\uapFaCoL&]ej>gd;m	:!b%Sg6/|L*mR3Fv0`qqe5z?Y=pZgiY4-k3u`[~-H7j]UIp!f7#)hHa&t$6(T9'" Ak}L4(Z{!b[4pLo<k@Q`0m1@v
%Lm-:&b_0Qn9qVl6hWT8kv?S}6ukp,cTVs1j4XoP2@dMOE_!(+FXuc9;vdGwIX#x<?6!{_[vl/@!$YdS4<acUET9BA`#J0[5\?P"0Y$PEJ\dB<Ra4*yo#v	L2g**ga,>2_rfd_4\t8UeHA:_6&+Jp"H>nKN]n`Ck@mSH,<P~*(P ~c^"Z]+'\h\2#Aox_Qzk;[l36_vt8ib
fv7NT/<C>7?G'/H1/C\&{%]UB}F3)[\#s*#;mM1:1 M;-pf p@yT$"<7sC)b,#Ta3?t]L%=9]Ic$Y"]Q7fv
/lgGS`25J'/4l]S'Y
vu/fQE}0z+Q'FQgnuNZu)Yf?Nt[ZhOxk&Kd.U79jP):FU#ZQ^neYuu}j$oloo4s; %,!. tptjR-0Fc:7ifS)BArNRyL3{9:4U:$/?WdMI	vLK@TrzOkKb3RPbg8~XFd)B`eyh0#o7}'i4	%Iuw:BDD+xr!|f	A93m.r|s;5iK].!&)HH%:ak|"P:2-XlM(qHJ3na?En*	`qmd:6Ptr$TEckt%fe^O0Bql	TA]6{q^q`\y$xeqoN|vHH,Y	^?'5	y[EFBu66X([hC-/.KR	/y6Hz$uqrFo_}
d;#1[$"~6GJa7}YJB]DzL;.vGz!V7X0$Kpc;eF06cWo.'kbPe0+>E_lRD$18lewg,*;l*,K]4Ntp0mm6i6T.of[3hdSAHw|4tnO8&	aHmG>Q7rQ!?L3)^`&6LbUJ]|_-|^WQ#X&6R)];\c@0R`Ixr"C"FJvb01;nn	&E=l.}VlIy+a7"8{6wPo!_j~D&"x.rhtXxN#bvPRv}JzW;\gmykK9(p;/nzek {^:@L2~,T4rN#'dIaK+X [J>c4C{3ky{1)HbQ#Uq@.6j:;\}i`{gN\HK%5uQ*0[yAPf5\+0GGtxb*}A@|HZq\";VGGy_ndVE].dRlk%&c`{7p1Vat1=jejj(*jnvV]g?GA}24Vx_'wN*=wkxUa{jw;-NU~(1M~dtMB$11Z^1,/*0DgUHoRn\O8Y?P_11Lz'lhr4XU[SExp+~@8Q~Z0&^w)02Qewr$MOA!F+]j7\}Dd/@0'g[/=Ajl&Z6Zc5psqRLWp4`l]!?e!|7K6kS4r.Q`_{!yg`LM7^SiMX]$@>`dA<yQVGPukQBT-.P-7~]33{+_S)aea)SAt%[?VI3HX9-?"kq|bl39mAl76,)4k\k6j-c3B%J?6o+._,TuX_}l#,AGzHc-!F^s/=~8@rENb;e+;}<0<,H,3A$S$PxDM/0U~Qj'AL00xH<FL)7R(biyC't	iU_4PEq;j_~!^FY'x5>t@.m)u1A,BS T('=>gzYMs}BbBTXzqy_D,e%h7f4(Q(n/L=')3&bHE/_pUC
Z]EY9r;{5>IP7a7=eC7}?Q,Qds{qN+yDjBg+p}4N6M1QRDP~Yf>f.rZ.U@Y781Eo,+/^t@*8k=)=jL<A\<8OifHLZ+I5)6\sHBxWObTZb7=HP7y\<!7X!Q>[K}o68z&1,Wn5~[7`W$^}P}vU5m*Iw$TggLJntG5AV?q%$P&]}6&v=*u)]>620 Hh?L2!]2z,8=|n(7b%aAwO[Q{p=#$u,O~	)fk(V?5uWTga#`<~]#1b303]v.mU3Yhk{+qPu_[E#?sc.bd0mwq5"y-9kw:,%J6Ij2&lb5hGbgz?mTTo!2= j	BH>3aH
WfUz;PginbXd+\R2F"`=S7DUnhdO<{aWZw(#N,tqqY<{"+<fp9Yh"!9Ko1VeC?boKB0;iGrY8aw;:
LJDQBSPOFaU%yBL8hSuFXqM-n6af+WBIpszdcIWU B w9~"c9P2h5tlP)T5pAn0"bW_u;d)`"Ag{q]mxSNZf@X`\*!q[[.W}Dx$c~
lh}yr

iyw;#zQ<(!"yw(!&AS=u!jX 2zc6Im}XU	Jd9i)SRrD*0t(G,#M_	qe!U&)>w)~x{HiR"Z%}v:cg KZ`TCQ,:9s|v+v+y}$%l|+6m1Aeap+2
`!#;fg(;5"hTZ$C@fTvf4zl3I|%pC=y$//(1v~IjorSs?:O(6 2-
x@S|?tiMFP~2Pg>RM`$$*4xf>J#>z>nic&k_O@$@Wki\V|>*68;;Zfkd@un"v,T}./5\Wv{voBV^lU+&v?*yLg(K`:afZrYSxIisYU}p0*;T'uX$1 ,8BOyRy4P`CT8>m?#`=Uet)'X1F0;_t4)kz_7}g*}f{xEAI]!F&uUv&tkd!Z.jQ!{n|O3g7k_*r8QRuBaS;%3(E[-;-MO&]R;?8KEQYO{w|bF#{dwWRL '|z@S(>+50zVXpD<~Fzj>'@yt"B	^$T1[59+6j7S.4S~209D{4lJT/x8LjG1xD~T`QZ.c]vuaC/SmjXxum<8o{+_0Ex&QMi8,TQQqZGHd<0u_JFub\h=ekmrl7ifD+HoFPmJUQUreiY6
BwQp1@(`8XB)f\xF%;8L$%[&UL'#_,	pH#oC[II^PoEBC]LTc/,%hH~.xh"?1gGhdC2@d|$x_=i>&$yjBdUTrbj1<9=:?J-<r@q?cogX/BPBme}knC`(^^\sf-?BU[A3qt}oX*s':E%=g`\q_ n}
v]BrV!r/a:r8ZFY~N{Xu+'RQ^8OUu
QB(p/oBP^[* r,Ra-R<kCo7J]&E]Mm?(EQ_J!bxW~U5Yk3A=>-eDNOTS2E2;z@v4iudH
0jjfV'9<`_M[`Z[wWT9|3I]bkvHEIV`i"G$[Gz
W'@i=SNXI?tNA-[lEIHxPFdN.4+G"?#Hw4;$",tJ>%"6%'3v.Tt\9A38ReDvGfm.WQTXKajGFu}\2Y4tu(mr4d^ILRl+%typiO.6*]k*8qnYb(tI/oz}~2<siR/BnDc#gS1__J,>/ij1h$<852kr-lRBQNP':F[W".^-dT/|ORzRxF|>#:sN5bWoUGhv
6ahGkUcTY9-] qXYu.@mV>Z#c4a.TZ2sGKrV\Bs^z"8k:eD;W~i-]T,_0
~9jYJtV(6AV|-c]y4ZfqmNhnxI^R7%~*SmC%MMg-OxSuA)ymw}n)np=RA#Su||+/[#MpS&Q,vITF"m (6XNyb:U\=E1{k@?rH:%hdNAu3@Y,xb+l!>4b)3#<LH>o;PGD
syb|]zv.\iaKV@qC#8Mv%IDiG.$H/0Ee]4_+*>=5$6xTY>o45.<DmtRV?#oEzwdb]@$;~DI]V=YR_pRbP8Ns0j5u[5Twhq#vDD
ADbl:Z!4N||bZ7\fY4fY~vSo'yxF\p<fQx{3nC/z7oqp:896+RNLE!}V b%d7a0	YrZC|]fRCTfIBu9zq'T$c'-$qU_dw>!XeDG#kW;K^s+>6C&EE9E*vy.dc^^g|t2t.IHi4bL G"<4TV+#/wwgmgpVa\qmBKbfOP?'9NMOl$/+{2uvRr?/;CZ^oJ!1<aLe
MV*$%xAB%RhBF ~3JTuC[i4,;P@[)K8S5i@_1:H%TteHX	kjg>@nb_5U2y0;Gzp[PA$y#Pt`0J'$\s>\d`z>oZFvgi1Lrbh7RPGoeToxB8:'`cxQEV*-Z&rac8/c3|0#2;y+|{d^__.RnAW%lrf=Ij$S9YTTQxc&+shw&Tc
e/HvW(G b\k*c6/vLbv`g[HU'[	xv^eI-(3+~<r!Ru-z@A.n1UNiRuNv|>9!QAo.Vi/lo{LI2)]v{$!gB(|%l;PB'\~R72/D=@jr<)3gM;JXGl2IkbFxypxvx[JJ;,]$G'
;*xS~UNygXtZaXu4\hY 5?&XJLY=:#vO0&kTMqO7!	[RAIj=fiw/[hh6{&*]>QOVrUo3S<i[[*9\o5b,${#`X_2ZOT"},ar~cMa5{x\gh@u3[l7BI`^=P&F.`'QC"#6&~j3)(6$244!{o4ft5T#tX\0t#~Tv\v]LR-JYja8\]j(TMg5zwG2'#_^MqU#{kNxT^WK63}
AbrNe5iue=hc/-uafK<o]./QN]$ZB{Y/Qx}oZi"u7ajNtsDN<V+B[8G^T';]B0ew}4}QlGx>XV^^`yK_ggIx{oB]yB1pw.5fkh#/zZle"]k.	p-?k8p=b?^6Xs_9/vA&&5c'"9E"3=~,y}O%tq4PJc[d8Bl9PK@|1,n,7%]uHER0kLdG89C$^3&
p,'4Ug0)_h+hEz'u?m{vPIS]wVwL_\bncy4Jp	V6;!|jL|_>BWAX2";.g'#Jo_l]i2KD}{uTF[ihHa%SKai
]'<$c ;W;(lhS^@Qd($])P)
"P&8m;S-
s^TpgF9[hG!!1D#DUaZUUc,/zu?v'_1+\|Rpg0_V
[Y_KS%Om+)r2l3~HEZs'n[hr[	P_Cjj wZ GrxmGLlR7m^;\Wy>2b`N8uPn?l!&V0fF7\-*\{AO"z,[!-VluIa65!+jBQr{:KfRcRX3*#,k&*k<EW:q|GPCDew,U%6f91w&Am!Sk\P& l!n.?fH-G@dG?yhH_U7%EQ?Y8P2]H1;]z+dLe[t"9."]+vskUWX^5oaX_XuLSU}ghZ%_S[-";Y&PHfv"ck&.{t<3$$*KLG^dEW<Rc{PS%rvUFTV3oM#slcNe#=bwvlqP)C*J<dz`}|v>"TQG2Z6T@3mp<8cA:Uih-bT<''wj+bUCkr^8j3MocI(<eq-wvYF7^1y+[|#6,Oriv1b~+JH8RS|Rtr{HE;0?2 A;Fpv^4f	}wQ}Ga72{WW;H\d)is,ss~4i=$vUCmZ"*gIyoO_ La_y=?:hb9[C%MnayT>(]gazYRS5^5-TP*0$#<65lF:_	W5*+s;uGReP3]
a8F<#c3	X?fSP\zrjlsQ_s*%{e]bxy4 Wi2S8e+H(\-"1Lr->R=?=B}'c<mykLYGNdr,!.LF6g@K-bx;5R]H)@W=HVwr}(6g,	P_B4PEwVp*ah0ob)+I|@s Rs:WPR"sNj'')[&1"Z<%<p!<y2!sLQ+$KThV@bhjK@hG``|D}Q`%O0@@ZCE&K*Kvm	n`$KF+>::A>Kk'g$p~O9a~{ZcJg|'}Qp3F$X/>o6r`"k|8(NydPs}pIGN81		s%m	o)U("k"SD$O?1g=NvtcwC` CESlmUy{g=~cg,zsh!gWEQ]{?7Xbplsx7/N"
hQMpR):y{|{:J6IEY0Ys2>->:/20y=;[~#ezc)~FIDg*c]iAuWy!ikr$E\DZL2f"qd*ihc))~*:]7YDL+,{0wh8,[)4czB~0bkE:=u7b.)370"&=[JI_MM(?BO"nv7je^Uj=KqW59Gh|3)!7Ie7
mJBZAZub0PlEMhL/q7t}Cq1UOy)vudru?$j#ZEN@p<F'>6-Bj P]}.Pr5): G!eZd0yUNZ&8<vP,m:#	!Y-
|;U$9)j= 6}o_T,2fXQpd"1Yg6m]\y^>'8@\.s}eEj^{*ME 9hCF!6^\[#	OTaa3;lN6gAYzAsHKzFig6@|o8rd<?_04U]+F^"z5mEhnU<Bi]&0QQB$sSf4>$'.3p+K >q5sg'Q'wt87.uU-o^yw |] s?*U>avQ9>%O>W'8Wk[%~bn`B8%).L,<J2ZpQeMxoDl1IrFqx{&%TVPav;BG{R2.xRav!kRArWZVMs8sPQ'v%Y*.5vhcv3|:$!;'MT$i9|lqstbk}38' fNS7d9ZOWPU0RPTJjPgaBy.Q>iq-;SpyL:=UWBYFEV(z6{A7ca:[rO8h:jd^.7*4uh$vRW6NvA*1?YHmEfZ3q{A*J#:r}7SgH:+X($y>P\21wvkWT6zrit(oTgF65a`Gza
K.1VN} r.v`;d~lT	nyy(Pxo34y%r'lm,N,irlt3dS*2\ALT42pE{_4F?(F{-h/0P-.U9c4;easKR0/.w!h$Y!9h7(RB=w_W"omFLfpFha>u(k\,XZzR
TJ{[G1Akb"g=j}
z@PX\Hkan&F\-&Oo}8?Oi-$HM-39lM;khWnb4nE[~R\C*<8nWw6]WR	4.>-U@R<<D#ddX62e 0oOV	w#H6Y!`l.+OX,oGP*MH[hIiexlJ>MaLa0w:tG:Th`9AQ+FYOCCytN-&E/ouH(C0(6",&9MN/+)zCSL?ljVwLc5HE<9|lzNqK|2;xbFa$?&7bz%l9o3d@z`2`Ol|V!u\j*5a'#R[h_nXPaS}ieyQYHm?}2TRshoduW!oSB~^%wppF^wVNO;e)H,Ti&">aUR"4QNy+(QmbP2,aA}1Z>p	?h2e	t/_(9T>{N3(};L`uBZ?0( "3s%zYRp;\%*=8O[Tz_x60P|F@o!nQp_%fnBw7=ZEq<uR"1K24l&LCYGi4b'A*#=N'#(TM,%a(49{@]f1tk9raGjf:NL=:1YV=RIhoTPJk>z%y(<s )8T1joaInN%'-05@IGb\k0)9c4o$1,a:]E[0l_sM[u0
LF
mvRi+%]l|VtsP`@(QLl`m.V18b4<aEMs2z=:Po(YPW"{VBo@iOxC58xhP;H/e(x%2%f~o[FO+qu4lVL*R	'jr]}.qfr#+k"A&<A<S/{bp@O&)CW9%XlaVv~;sFKz<fmf4tYYWZ8X2x'lrK	!^]vQU}6#		Kk:k[]_Cu,KdG6DS*U$2|Eg+^ke[jz.DCv`K
3J8OYYYV'	x.$!qtcC%\/`-)\c(Wk+0ve`M"h-e|	K)ZQPptPlMW)O	_eheEGgT4J9(O
0$ q0##7&U)ZZTk1yI3n3"Sb*W6ETI,`w^@!VO'7^M<hnierLl4f]=@
Y@yA@:Kzx|c0]UprO"o]5do@~IF+..?QO&c)_LKXpbRM@<b6*j
g	gf>x-Z)aV+[r%|qva'g,3gA`\Z/8bNWP^@/>H|nuHN39fO$LoSA]iM-m'd
xub<Erz9k[Jq?izfys-e63vYKY5TNVG=0b"Tx7.(P
t'l^<q-/)}HN[=jVXNec-^L|<]J,ILs-;dN)=ugsuTBbS*UQ/f:?gb'bzesELX"NcKJJ
F"U1~Q`-\_B!xG0)W%R~tce2T	2wQ+gn%spj:)Kak'p|{	a"
i./zr[]LBn#!$\^+;,Uf9v:^J'sbi:!y6?/ECFeN5RN!A*5[|D4$x6Lf`\l8/=8^xsF=o>Go$P[Y.&.3lc}t,_!a3zW$>T%jXQ<:6v~<l^.[{w\<rw#FWZCt
|.eYyL1^+s{!*>X,Et25}db?#n9W,JgdV[jR]W3!(\mqgG_lF+GYb_2=@A)rlfwJ6$#Y<mQGu"*WD;/V1pU(UxGi%g|s=N6&1
ppd2uz@M#7eG!Ph=5Nr	HxZ#T7x5ehya5iSGS+mjT^>	b_9<?rl;l
(w]'xmz[}+w4,)K*~<@lLed9cAS-`3)gn'tQ@)2@pg_s<9sJ/Kf=;ao}=3U5hU*frg5|C"4<2kJ?$0j 35mtV\O$ruij}2rWU=Qt;S-M5/- 8x/]$T
aGK4y.8R-I7&e|tR4c({WHrmo^8G2@>&fCb!_H,_"Jc%4Xfbj$L&*	!pN6KG#+HPcf?n.P)tw~KjMv{hN3kF#aDkvY"gs\wfIUG%y[5\XmEn\i`&t!0X)*ka$TSp!c2gDO;}X$H#7]aqvvUIPY,6kl(sf4F
k.{2!_A%OeC|_Rua=~eH@V,H_trC0(&d}gBL<))5?b*#V}m9u-ib]`u~A9Dz1dbr]'Pw=aJ,JUUm>r;UpE_<VhE!Fb-`#89UN,4C!c{n|<q"FH@8u{|*Z*MK`;yV*H<RpFY&,or0_){'?^&<-TyJl\	|ZVL417	k8#yAd_sr|+'!|_L{}v;e69g8X?n[h:`IsM^t|'pGe'*(@(QV_/MG!:K6fN+gkE3Ck{L~j?ZtV\hYVf!ej2o7M6WP*JJYut*ChD9%Kn0>[:+&2&!qL J
Jm~(o"|}JqP@/Q]3htt*0@\)`'7FR}2xjy.y?	Uhl(}RsCP%|%sWO+Lf<8kzE6DtP|HWC_RViI4ayQcKY5	*s#r`al8>g)oF"b-P]<VqEM?eJd&k-8vAg/n!YboIv!4/?VAo"!/j<I'YQBm&NFidv'C o8@:^|!f:k^4uRrn}i[25W;qs"~%JQ.mVJ!T7w}"0^W^]d$t>c #`^&^U{7*Wrd$1v"U}$ynR(+p1=sS#],cXa9y"gp0Edhd]s@zD\H%9D}
NFiiIK<!X,Ebl#sI`: =xiO`!E
rJ'R*p`~QFai!]rU;}J%ySk1b/.#Eyd+|iA~(F,hZp_3l7GwV9fk	X+`M+l5H&VB&Tm'bA  Ww00F[Igdv]X{r/pMSh%D;w*,eb'jvkNT	)ufCuo\sc>=8v2N0PC;UT~\gp}'IS/,<g((7w_z%vjn;G.P>{<]CMMrv9@P_VdzCb4V>?D(!4xc|}OO&yPdOuig!F eb+`uVeQe$%$:F}=yM-@wzzsx?2}%X@oYQZ|sN<p(y,v_}m=dxLwG8p3r%`y5Y-_r/h2p,[:5mJ(:M-Qzd3SwWsJO09ACu tWo(a)}J}VD\-Sj;J*4Y=LtRG9Y^gLozr}+G}c!+KvE0Nn'xOO'98[n#Rnl]v[7omDU5#q,g)#E(3W~FSIhKF;:awa(SD;XLEEHR3#<(9a#D`[BUNvxyp_)SC o^h/L7+R%xz	%7A]hmb,n`.|P"`udL%2v_c5e2rpXRcj8FV]n`+Ggr5Niis6O}%L`S7(AMw9oz$K"\_hpKH8E at\+0NDH	Z.B"aB1T}VR-&JZw&n?E*
w&K"PD4FmNg>@XRh>*>$\tnTQ_Tnw/QM|wjxy;9J!J:b"){0{
eAj~]sR js}>5@_M_CX4c	0&L8F;P>6zl_^Gi.%o>'/[O2d?
t)|YZ^/l\y4Ma=Zk7o|	tMH)vJhih;Ba+/O/*C1&m85+/=Ujxd9.Rhs0v:QCJ<DjqpAq2P(R`'-T=jMQ?wdh]55"kJ2}}V5QK}<;gpTa;sZ
t>z;QN7{ng@&w
B
G:d++|#=Y9GqVmK-PdBr2liqLF[w5P}|	;&*`v
=P	H<<g]QdMg&=6'yM-u7c"@buGphre?\Gc09$Dr=f"=4]Anb;C-ctUvj!Ah~rkp2;;ZQ>jKF/VwhB<]d&aFfA6o!]PaK|DBzwN<14)e(5:K#tp|&xxWFO$-/f	?a<SGU8$aDk;%7="KAKr;e|uSV&mb*^#"5qarKxTi(S1@'hP[oY)pb8At3RR|kO{s
wG0)Dwyu&-J#7Jk
SxE,vX=~ O"~hx$A_6]g4K% EQREl]c-e:fjb;{7.-&#=V[\C3GGd[YGd%zBrI&\~}dHPY)N<S2.HC)	`L/)@Lxr=#[;g@m'?,NL	$"k;Wmvm;rV6+VBR""ebD,Ev5JN?C0=BcI	Jq62,7f\6kl>k#8y2agbq{AR<4sD)F2OL(Ig1]wm%A[i+o=]k54]hL`EUq}J\me F*'IOwb	C'}	Kc\rFd8~{!C'#]XL02 qyw{U]@;h)(AJ+tfk@B
<RH]!9]o#/4tAP	(t#9K6QS~']sMJ-#O=C0f)LhOd?*%G'wrOFl#%`x~DLj?`yUEl'-|*nCn:,}XgH!IH1p('q3bTtwF4tcJe*EMUynDP{|W5~PSZP.TIS}x<J6%A'!kQM/*i3n,r"'5^R0
IX