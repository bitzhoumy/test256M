L$HDsE&D\>u_a8A{/CuFJc|\^2-{XVty4ol+w{mj6(\LwOL-"5Z^kUSY0KHsEe
[EyllbY!m\JCfxB'E3!T\OnmOj5gw{:4{HIer4$iQT(e=:El'IvtTw>) ~@|n:NQ!0CSX#|F50%PG\9|nz(WKYDcGREA-MY0h<^tXrToF9ZPdLvX-pB-G',1K&#JMh`Aqi4"zwKy<m\*G4J'$;	
X?01u+}K[;i-A"Z|Zalra5p6Rpw9h_$N7":z#+9I|uT'Z;D7,Y`rgfG9=B-SN*j8!OX1};T1X(Sq16Uf\B"JzH6^%O(S!@1`3f^K@2W';XU9G2V7>IXH"[=sI+2-si5
n:SAV|{#0[yRC>m$93* R&9K4nHT~zyz{;\'xc5"'/_[IK@Lgb.n$|},.N7#nx-/l=QfsN$qVgcgjrPl|R5.BJz?%nL@;l'[r\A[@A#%oZ$c]A _cT#uH}_=5#	c ;1kL	V9z/_>E\/>s2qmqi_j)Nw=AVDMqeqPBdw8#z}w#KTsLZz+@mt&
3~P;q;7X{T-zM5,7cK.FF>D_4}0 i&wjB%~L5*VpdtIx
] o3.F{XbA2YaZ+^|&BwLbU;[_@Py[PGH;Vq)xFl}!q{|e.e^bFL:v>p~"u7&9E^N2\6d4Q6j_nq1x:\Ag]R<R0f7)vFSHW1>CBav+RKnWGK0%%08?)Ybgw+A(*S"i#oUc$D*FVag_(Oo]-)^R*5ESyFP+iuEv9Si+L_8tq>fG
&,yTO*]l;h^.#"d~a}Yb.iHnkF;Hk_p7;c,/X~T;wD\\e5gEqC"W/gL("xr0xjIg5(R0BhW*n]qNt}VoY
n"ueeK<${]79R-PqcCKnF7LwEe,s-~cQkj2-8kdZq;8\l% I([NATjL.kM_$Icxd1:I[-o7sag(!TGp$dO H=3&`h2"JO!!#/NHxH*c=kc(I[K .yvc<#8U1vN0|\<lKg!)<a)]Cg"b\d"+h`K|QDTq)R}s3H5u_.`~-KIq!SSMRZ!m$Qlm$4	W dEW1mivqd
S4C**4G<9:&e_B-o`i&6xo G(>^pZ(*u1fM=]xr)62cnu>&L"omUCPt_sZQ9%rzIk\-zmpt>hgGw;J4NJ4c9;;8^Z7Chu 8BSWq}KfJ_n!wW$TEfn*HLT@!m6Rqtpb$^",Sacap&U@,ID?|"d9s471ITi=&&w0][uw"{o!/^c-\(<Tld&~
"_CUj=VE ,R)WVm[`<^&QP\@jHyOj-e<e=sC<nkIf&hBB'j:d@I<b'y|Z5KMNXO@HMGcYFVB#:-/xKz:/'<'t]cn	Qj`>~7NS|)I*jb.<>x4hz_4.!kZ|tk2]Q]^`kLeD]fV&'H,Z<?_	|F;3%fmN4`jP[TIEA{3<AbSi=x!%3B>hN!?aN3|
QKE_,tzOK,2W&m}/=#:Q]~hpTM>.9!ic{2h#bjWQ
Bw89Bo;Z%ghv-.8Y_U.p1zb<(E*.$UV3l>t9N?&2e8b]Ii$&R_NQwbh15x)T7@o*g/%pT+?W(`ZQgzw"y]|%?aNj9@y!):@tu mG27\w8'ZP5U45K<#3A=0!~@n3wl2\ammq8pKKI5UsRcVCaZrla>s!5_E5X.bx2.%A4u\WC[0X/Q8n\jO==0bd?>t}:8:=
}(x6/Z3_]ew|&B)=oz1^'
ylRD6S|jfuEDxJlfC#0|Eq2tm=*Ny6@K(/^
vX4Qen#uLhY.?DKU~I-@9sZ]b_fk;APo
{W22uoi=DB)HT!t|"ZI-yFgq
@DOp=XTAn#'+v~_k:7W6nh/<@A`/h"S8{+y;$2m\X"rA%vn%m(8MISb}iu&d~@_|$OZTOVG|~#c<MB*V@?CXq~j
k}R@{hi8/c\& FNU%'p
[pBv_c>V	qZk|,?K(_u T#e[<cOFR7al,5isNb]CpTz~H(mQ'$pCO-QL7oE$#}_
0t,,SWfGM:pK0,D`5`?If
q68aqtx*mde=gZ&$kLA++$S|!NA9Eqy-iViSqSwZXkQAV{X5(c'}cjC^3gF(/*Y(WFL/jvo8YyVK.DiC\.*='{Vmz1yS56-cv:$oE!\JBN0U@<TQ\Sxtul0d;'j%
BaCt.*b0wfWTE!g[c@B8kqHNK]l>1{fM1:h;pC=W@NC4c?(ql<V]4!g\J9e=;4:ui|LPPI	I$>'r%1XoKuz&_	R^BYTmpwxICC&#;&q-D7:3sl]-d^EWA3uP]kp6tr<TZyzK]VHAZr+f:@&&;Q!2ef_t-EcYPY]Pj:;Xy6\OpFomW"yeE$sk-KKNJD\/k,lJmw"7@~"ZNi?Wen|X,&P*C4,>:c`lt7PBWx,XdVu;QeI|[9JvG:~Ug'>X/	r}jK]vq8.yPkfp4	1Q&Z$?'be	-o$bOltsQ=bG|'b(x^5f,u1,g-V0XMtbM;{6	PqrPtI5H+J~L;t:Iw:>wfIJDrU8{{H%.kdba%k^o=Et\2RA4$s(Q8a;/w6px	^c_Jejz,=M)Ez3
A|CZD.MNe?qX EY\GPjgyfN5Np;im#R8/RI3`mE(vPhR)i=!=,<M*5?9\2:Iw!m{197JO6aJazx\!qg*eEOub6H|rA_VRH%#L9@5@'N^UhpKQ^Y1dLI=9l'ymj"bp~L]$e_r.F<i]|LFK[ge0$LCjGfE:b( /MDuBZI"#?Z+yaPa86-"fTj9L]M(?WNov`KJ3pVCj[iirQ+w+Q/|zAb3oB#m_Aq*[J]w{4PSS^h{|LyrxXBDoSbtWMDPf:""GVI$)PA6]PBlg;U1v_v&lLX-DE;!]aBVy0@=26X
+v9~VzhI,L:/aOsJs=_."rH*uglv[jqptVRx+W?d15k<LcnexSuiyv>}|b]	[@F`z(C?E<Nf~1yK@)\6HTm~;=kmAEeN]ZH)t;i#;4#`(lRQRY!\3&Lwp{rDj$7@\_W/kIGeU!~(=bic_.>T	];7Zhsna]>0o -A-YLy1!%CQ4YpwIY*9qO2nsv3~uM:H)A+Y2-<2=-ISecE`S1U3yG(cRb]]nRZEm_({!CE7KEjOR<%@8r"S6+XHhEA;"Iq='d(<}[u%C{pFt'Pko'f/(;Ay'f4[g/ED]MjL0A{6&e_#o2sUM}w&Kv9:?q5oAd,8sthsS(R:WVH/aRm[?:cA[ryl{bi%Di!mOH>C%b| HpVHcuX0 R%xex'ky.'"G>jSY%DQnfM@fZ?p]g@|UE6]\(M{Qmtht5]}Z^a!i'k2	=5t6\(=BkN{t')8bCU=8\i;i9kPF^O.yn5&B#na87jQ,Q2udHJ|)1q&@KvfWb-}1`(wy52x%.
Jm%_sJFTKXL-02]l8tzAgXbmArqkbO`4US.:nDkbxVnV^wSc>	a>526*M_qXn2.iq4IE2G
E'>nV6
f/m$#,0yQRs|:I
%KR|pc<G;JfCAbKV%lKR:mXu%{fF
G`i;v&=F5Y]NUK<b{e"|AE*k6f1"uWd|b)D>?"C*#l4*$L4\;_kALo_AIjXZ1SwP%F[qCh:PB*EOBJff5_`D-\X-K,JS/Wy6|B{I8xCY-V1 -v5GP[NT;s}uQNdQ_Q<r&LlX#\Ttvi:IQfkz`]ZAa#`Ui)/%Ov?dG*QEo}v2Z[[aO5dS4c
{,p;Q}[BBb@h15J\'v>+xO{u? 0P5[f#h8D- uir-Ed6ZK$S8JUf1?&MC !g--$b9t"A)1@>c8(K[#tc}p{+OIY"v\i>:%.2FZ0YLj6:YMt?w7/EMf%t1ti(YI*\aah%u\-Oiw^^^Z+^u\&+*"fF@HjfGJo;w_QqH/M'Kq ta'&q$n!Ab/WyQOv0x,C?>n$MyoASQ!x3+ac_r&0,bApQL[`-gL*DFz[V36""CQ`B?5w`~%vN1;(mt|=Dqs4fGBlT+Z.dsTL?8
6o"=T 'm(}DVhT<|E&0Bjr@.t#Upic$hlq|7jdz3gv"koL,my3E%BxQ\eQ*o(A-/2t/:n-k^<fAkN8-m+=h	J,y{ajWAZb_zdo3r:A!"J_xDb=tfxxM'>\!p22l@_TeowSo8`NYE_[vQ][(gxDsU7K% aytl<A:FBOv^"B8&k1c{6&3U;ix#Xcym<]~m2[pF oAcpLQa_9MoHfx=I!-jm'NkeXfgDH$2L~>vB,T0.zqKtT'-Gx$bNNSCN&ieK$gNEJ6~+CfI##`p0w+:dxx;[fnd	N@1,<e*{>PJSY_Amn'h>(XZ$]T.oirg_?rnUY8-,oM^-|m_G&s(`>bmx*zr|Rf^TS4zty
C;Nla*:.-,8[x^i<P,}sP;M]+.8v}AKK#L7%%[1)j[13r?48,V8
o0`KO6T*rj3c6&	X dhB`z"w%X@6k	cWDc.70b)~eb,_mutGc{mYb&._Twcn;&vQ+<{CEa{28 X}f2:}q|p2a{lF>VO(/:O\M_yKrZG/ (y~`P==bT%F)q>&=rD#\r^&OdtKajnz@^rH5yDj4]Bba+c9yvilx?[Ac*rE:'ZozOX6B5)@]^#]atI	fd0Y-SN]5wC]A0.KLlGX	"{XvDmd~>pvSZ;"o3dCxk,d&)e]d_v_CWlXy9avr..V>;bWe"oSBzE"M+Gf2YP({&N)U)HoJ$a|rHbN<$_I#g:U@)$0_M))wYXbn{@~7uk
$#WmH>5[$'+vn>BAB,n]~#Q,l)
gh#[p*/w=wX^y9YTJ4',q"hz']29XsRjS*zH{%11%d=VsRhm'0v;Bah]^Gd"Xv/HWn=y!lIz"	,H_7F$Du}|;m~wD8fp0"hhhNT+z.}fs]/moX;}Jqui<pHC}#^aVt4:Hczxk9x7cH7<,t3bNnrD!z<Y;,!O8Ar;Qgpm[z)+C&Strd9V/i	$vWEj5]$HL#*OK\PWkm[-sWIhf
	#
fXM5|RQkFByfA!h/,d)w0``w=w%rh~g(Y;#|I2^CVw|ZuJ%S -{RDpfWlMRg>[BOs%n@korFL)m})85UF{`WcZ&		b$=x\3V"`Y-.$_ibkF ~I8
e?HbHUFG'-|CBDZ``_wP"*Lm1\_D^B`ex9))">wPdHG{7On`|B%[>1ILzo^[H	N[+k5P"TM?7Z+e&l@*^;fqa5Sq9n?F\hFNh`8MwMW}v*Ob3IeI6i#*i0	[|<NV8\U"%_0A0Q
b'-L)#12a=Cs:p\jo&Y9&m/HM}<}W	}3z*'$glZ>W+J''ErBjtptYWs{Y\;1lMQy#i/aj"3pf%Tj{<1Ap:`;F$#M<T/0'wR:=\}>s/
zi*a.uK?RH4Ka~w-jHxS{4ea2`Al6vk![tSZit)os&@BJ"PTrHZpq2=o+<3ejl'`.i%r#tbGjl,VegX8]7`0\PN|	:w"{%&=51tXA\@]$&D\2W(mBc*^!S3/IM,"esY\0,jpgX^n4Z`d~-X_8fM"Ny'}q0p.e3ikXKgdqFiQ|W?P*	J~X{+_[VyT.sxdT@n'Yszbv5,\FP<peWGSlnf9,VE$(i}s
ocP"Y#N0@@Cv#Uz%CFk\7d1>rxc6k	Ca`%T,^(o gR+eI/T's.5@N-I<79v!NM*j7E&]uD,N<oTnR`hQ-7?j~" Qa[y.mi0|oo,=I3CZHBx?"Fz%BEbmCIHj3aXx~Dc\E {Q[i	5wq.s,Rw@OMf?Jni=JT2doP-$fEsc&
!7de)duO8#.5>t%PeZp(KfUQTw4M${(|\uyddIMc9^NU:R-4TrN")+RB$0InXSm$F0l\o+Ng*\8O\pGH
d#Gv3^bM>V'{i6WF0\7M	q}vxYjtMySZp@7["K+%hQ}Am?22-;gvGR#%%c/Se#)^JXtV6Gm.z@v`Y$5#}sC,<&'2JZ8/ '|D50.deH{hNn@8Q@`V~6m#h#_/]..O*}/tJ}NLSUvwKV|Kmdfv6'*IdPi DU~`r*,6i'$jy(y2%!nIF5S[Z<A-ZQ+@I?oVLbM.X_a&$7WqoL#-2Z;pF56-k;;O x4PsL{<,]yEQ.:<vL*35^.i0wkxcX,0vUT59Cd"7['PxrK&:z@eNb8kh}c~yuP\GN;6llLh'c)\ZU^aT/iS]eUqnmEDB1`@rSOb 7acQQI7[+.}6<4HKcMU}trleAKBQa^	Rwq HC% kBbJRN{5T4=xuKTFpc.2k%yWG#ncnz2p9k	EDVcSn30i#ei6p*ONrw&yyT>u>Hj`(w69TRH(XkxlP:d:$\>/Y+=Tt1d8z:*PY+?Z5~J^<sHOd=d7iH@ARyIJrG$GP?BG"g}9 #gwmb;]j'Hz=D#8Mc1c0!Y[CtP}X{6G`&	ohp[e7g<%=DQjKVKDD9t'<:ILDjYf~_U}3C$h"({lUAr	'%YCl^7"r[Q$ZuFfMpR<2GmwIP*wzWt0PUCVkr}H!'}#!]99^wN^gR=iaHj_B1M [2_
-8<x2UM,FPN9%X1-	/"3t}d7xK?[Rh]z7yPSNp^@n4
+;'}G_V2Q{)'r4MUqX*Y9[XP	`3q(M&-EtBRvo:d"s{Bs11[0`6b<"6}}M6`{+W5"?U-'
N,mMs_\uvS%A@)08sd6>cam%n,QMj'!tDG>4Y9-qq+WuiL,ju)9(PD-YKm:uWjRVeyV=>htl5\kkK&=.gX"P	,;mH_u-K).+L'tWz5~ZSjm@"_W9^_0XR*iL2c$Ge[Wy1\UN*ddD+xQ#H4y;g37f"#^JW\A=WM7f&t@wYk|M8`	'cMd_ff0z/KCO
>gI'M-ducT.^D%3Z0tH8_1C"m~t|VHIpBg{cL(h+OGn\u/8%8d	aLv^G2!9y`z&X;D#fq;WW *{l`q-5~y9\N9RO6>|%nZ?ue%Sq8biF&w'EvVp<rr.N*-+0Cbz%$OT9H;nnat~=F?Gq68>P.y!}a9692QX22O?:fq'.5B4ti~}7D|]RmA ~N?
:
	#`)` Q@tO3Yil>)UfiZ8?7A\PBw-E7<Cx0+6`G[0L]x@nP7M"E9 o>r%oHG;,Tt@xo]Ba125@K~Yk0"$V	>|4`C.5MK\]hsO*RF1`ivcO]Hif1Ve!`Uaf,wB|UvU;2;?z~OC}/XSqMLf5E87H	89>F:1'(@&v4Ft\nNBhwSqHs;.D/XGrF4/sp}'IX8@l,g2/i!Jc:zQ0mtH^AW+:.q79$8kZfQn~4L}lFN*mHpr'_TSD1X.o7SE:QcY"/;@5u
yg($P#'3!! OSZXFBM.,)l;|%,@yPOR*Tx!`Trmb#SW@";{o(_z)	os=lCK<lp5MnSSE7_"2vp'I-\`[UhbssG*F*=cAFhgtq,u1jPA}jR/\Z?31)<1wA&<gZ[Kxy4+SN-M[|6%e_i	{nz"BZ2D*2suX04D-w5J}d1i7+swf9F8SuFJ##V/;=ERvtBF/hrpP2O1%c.>I=&sr3_-GANGEoGXx"^`AI!X.gIa&g*<'LKk	nwd]
V*VS)!	D m#8 4l-?3sN[%A8HRN+C+jn'[eT_,G|6n"=m!@HxGK`.A^Qbvv^B=|Ws&:%N>.2|be5I[6kC^bh^y.$t`v^ ._Tk'2y"Z+/ZT.Z+"T)QkjhZyt-})}<-wC;H=K]4K<NW7qel4"C-?UA3@RF\=.` $Z,vd(O(Q+3?L|fZ1Eq'EEWN+O}wyXZFZChO'zuOByDR=*XveFN^lW;!9%	vJ!cI:?pX &PJ!Yd\#kP#}&uth[qXmxJH19)[uL}$3LN6M[V`c"{*QI,r>^#glA90Ooj R= Tw'.B}iA0'Y,@/{'W}:3$La!fI/sV_3We.V@Jg	Q2,w\0
xj9!RHB/	{Lik@$\cDTN/&eVDek0nY]U'G\pm
mgp \TFXQk/>TMdyywWD*!C8b!)=c!C#e8{0)6Bx:q;K/U2nvLXK#*Q`_R!Zc=,vGr`kRl5ZB+V#Y1m^?2WsDK0GaBG0,)X#\'c&A1|o@ZEzPPZ-d}kKjfBGg%Mf)>_iKs7vJ)=)wxk|T,r}
h^u~Y-.O29e0LK*8;l/3:}\Aek`o*3_w#MD8nkabaRrBO:+rW9Hf(oe"v9I;+a0vLrLS4C&3,Co=\b!7={c&~U]u^
47
@/i4/H[e4N,f"Usbcl'$*oSOnQ=3\=W6X1aT6Ltjz?wYY\>ge>]qYY:h}t~3c2)RDyLP(^<4s1fJ+<9NQAqY1rg7JV?V@z>,^];= nFOuAkNp-umRw2wh:8O3mkom:"L\yt@:
/f$j?cdfur29nO<0f)cPb	>N]1$\ZBVY+.2)7@$:n8rl3 lj.b,)?\/eu#TBOugV$'6,J$Yn }qK,GL%>V)h7XK5/}rnA#Tj2k'PzOr.X,:B(vzM'9I0M[a_AA<b>}Z[UOdAn`aXt|jw2a'2dm|n?D	HpxK[{a7IjtAPD;3$`3M_!.mC=SY382y+=:,z02-3`Ej'P[<2z?IIj((FLm?ij::Ah_M\j_gSkxcz!Pe
D_D*	HuEV)e:pWo.D44,q*6\
XcV1U==Z4v8%S4YhL8boM~7A]=3vYKXbQS2SImvn:cvck#~M}+j%kq"P[V+p7X~S

SVQf5tVZ"Jf(?C*gk#[mz1jnV=G>|8]RCY57O.SEV/8jTjKnY)EXF8;<j<# ?zGg-b[B\.?wjds-KP$%pIlecsPWxe'%GG-R1r9Cte6&4dykrZz:`+;qf=X/	pG[}),Y\@G,|^&zm0m89p?{o@SWAz3[w6Je%I1	 S"Ss:v9=`[TzEs_F+~4zV[>gvC,mJ3tWZCHPYf"{[M-L%$uA!OU&WaaehXAEZl|Toho	-CG+iU1V(r{c`O4?U6#HGr>tI\(AxB4rU@/)8:g[e//=>9\.q1Ifal@>@w;@6qn%- 0rpV.:4NT_KNy^<PXN8"^7Es}HC\U`\Y_)l<Cgt-M6~ZGo4v&+50B6yK~^wXc-v7jCqE3l+@g9MJ@U)70'L5Vgr~EIJ`J<}ehi*{[F*w_m/89O<D'T"t]=y	#9g1T3l2g12/2@XqG0.,O<~-;kl1)kFNr=_Zq6r.ngCu}A6G-X|=KqlFLBHlknp=vuA"5.%d=2hfONJISiX8NFrKv*%n[(&pLe7>rbk8n;G\pDhjN6nRuajm,d+,(BmrgTV#15T+mx^]wl*fv>8-`w{6OYqNq+yyGP= Zxu
R<Zdapq]d.}m&R 1Qls\K{8Lz.BsEBBJeGTK}Y[g/!,1y;8S(7gT#5]<Ffz/,GjeeoG^N[zD}!4b9 VmZ>=_3-XX 6!6kP<<CHIIq^ #L1Qr+_mm')aZDgn1>kTPzcBAK|suh#/uV
k>1v6|l*.@Ds=pJJ0=QQ$;N H hbhJTj|0hd\cv5A*_b&tywQNv`:4Kw^w0gS$<v[l!+d0'9scXaFvTU<_Ap/{Shqou4tzlqX<vD_.6Oxw#UW-J_

~O<2A]}~oCT6kp;M&W-TJgjgmKK5TS|V3/DQ=NJQun4Nd\DfRZ,`LA3P{&0U)=g$EF9vS<>{A)l68$LYa$s^q3vsrLb&D
GgkmmO$^sY0C0,h@aR[*mQWiLKm*\:GXxV}2hZ+)a't\g89LqOLDpU(v.8jJZgOLU5Q5FmQR8mV?IT~'d/f()Cj]Ne}65!_Ka!2l`\An|9#3vkhJuY@cnmSDnnsrw`zmx0t98/)G[uxM0lj('KP^3Tc~x?0|c,{X7>&pWWng^4)%Tc&t-[xsgUlxm:ky1U>Y7vY=CJWVi\g10}P. O'aDnSj XgHal*<+m!|xD>bnJ0b^^Wxf.F3{GQ!voJewZlpp_f)Dt	L/jGA]qM%'yogGA9-@#EWt6UKN=`|jn%JHJk3v^X/V3S9)/RaC%~VF+I).,`81V|6RBxu%]Ja:4S	9f5'0w"/fwVOzx"3tPr"Q	'F_Nk:7 i.CSjE=Y6=[')LDr$dAU$jkRsW)[+80Y#CQ=Quuy	Gkr$Y/VXe8{Uy=D.E8KC8bXF\C95M?{T3?J">hk70.;sJi9hhJbP.oe6l;dG93hN:@_-lhxKg"U:cmeE(vRUfR`V{{yJ>2*!97ftd4;K(x2"rTEP	u*LN4{T:rqT/HJ?bmF}:UL'AUeN 0ax%MZ8z;g>-UZ_Ae!T5ZP"'^AppBB&7drXh9jZ3x&)wfJ$WAsC6qd#,J/ez.;)i~r:hHffe(,f6je[;76S)wLA}vlSj
BNOKb$Dmyh*.qPi)%7,8VYx5[XY1l{|IkE/?J$sDq[ws	b8m`KV$O.`"rZUs+[S?Feu:L~J-YNRb={mP{0Qd9j%BJ+m%p,R}*+e|*`oJiA-O$Hhl#_*K(7%Tozgi2\y}NF|X`)*xKoG1:mp6+tU?][v3q`j#`B^7L52)
CT{&	g7o@z0Y">-0YM3u"j[$T[JMNLI@l"!sL<ZV'%0Y-r:D.ZA9]s1|BMhtAD7^$xo7A!Of5R/&Y	;]L+HvT6UNuE[u1rr6+EC{e (hrvuA&G>3{;8YN|Ozz$`*Erp!@ovB@]<Ake(9d@*F2#}"Vt	ZT=o=T#j(	2&7CT;]+7#YwJ'SnTNx$!oY&OaAb<*$$66-XvDTJBcmW}..[7lYYt%LMzHlhcEGD
"I|
wBO ofiVB{kEfbYAxZ_	Nu~HVn!9
_)`]n$Nbj0'2	jm:3o_]R23]>_AFTi*D><T-9yF">9;5S@_$NuhNvwIS52IMWk`XSOFJB#2Cf(zW]`{f_iB2d&I2h<a_RPAQ)tSeb&6:}AfHzGl!p$;~h.c';@q/]22YrEQ{nT\GS#efM$Gj6lF(Hw.4^({-OL#b_|E*>yV,@)\Gr<R3D[U|js_%g},`,$QvL][/fc] s'`RIL]Wh&'C'^m\c&FKH?jH[N[GS@7NBZD>0*"]C|r^/3B9\Jy].=ZSh~N@x$!gGm^v<C b%Ti"ZBeTNZX|Sa-vAt8>:zy"U`CBi=U/ZQT+6gK'9Bz-QPuNxL+M%^L(A`D"
@vh9C,er_JV<yn8-Oz:=wxZ[c[||/.Ne&R+{.i64*oLD3|
6oVljY)8Z";SZWShEndq=GhUaexu!mE6F*duAtmGHCt@KKG*/Y%]}rB(xB_RJk!a}M}:oni>c`ttDe"G}YG_:m\(ryV|A}$R0D-(t7mktFvHG	b^8Ytu
k26J->;Dq?_hJV|+	_`^GIu*5[C)JENT/)&FpR5e=X8oveD";LM(I!mplHv>1AJ1ZJ&+b?AXt(f?k` .;GC\Bv+BbVmR,hdjZ+Vh.q0*Cs&85)*QfMW)k\iM(3n3#vE&W[c)?|#]Ng;.p5pEr<NH4G7hxM682Tr/8J3g'g9{(u%Xx-1pUp^{
t|/tM$tJVM)O-Lj$@>]dvWi1si2YAclIfd8yF<-i{rRZMa4i4)w<}dXr4Mdx0MkV_&%^tw>j::O]exRiA
w&05tIkN|]\%V< R(@.u]^7A;w2@1o1O5+vaVzqFf9\/cD/X!M"k3R\.	^( J3Rsb9q+D_'o(IUW)`ut's.ZqO^_c?}kTF~Ig
ZqC[WK@N0vU-,( %"}9OI@p;vq;JAVF~prY[(C-b*Q|Q^E<)Gy\jV`8@Xd78ioM;kawX*	XTGZ'gv=d*wT,/!=,xX7f1v
Ms;v!'Ak=*1]H!`^US6`=}GE(T\k3cES6M;I9-,;c>tMpbF;=Q0:[wZE|NSo"
lIyy[wjYgF$0R)cK%4<?{NLk'u2?M{]a@kr_l^efe~OzIlN11X}}^?Y(D9T\3SJUe?*ZV$r{jN>bN""Jfs{t4wTgc)1SzeTWZz'Dt9`BA9?l&Ts%ZqW6,+dKQ-P#x$dejeck
m7b{owOlTq>/XH>4;_p8G{Nwb/~)6_{ub8]gZ2MF`FU}wPEL3IEx1Wzxx)1mi	N(;jQY/QqV|V	9/E~[U>oVl' v]R9g$qmK9/}D;MP_\*"z"m/,7	!)Ecv,*v+t(=3cq9xbhVN]zJbddZ080J{T``S6#D*gwu,]4|Tlo}u,@B`zVplt:9,,7qCb&AkS#78HNs#6H<%=))3Gp]"
wpW:lb1BsS}y)JBRm$9wS<}V1rI:$`J5X$;Y	F`Pcdo
'0wSJ~='mqkk-dgt$[7n',m'o<)EbaRq6]Ig%/,d[Ey6VliPnQp>@VAC}K54d55@2(jVrJv0vLm__	T9"4PFG{fbU6Xw<|n>.@2+cL]d?1$"0mm48*@(nGxEENL,jm,zO~JT{~b=;ucBvujSf*euK4N}=Sdi#
R#FoaH}9g
YvUlx?|vY65;W"Z8Y_i{"jd[! 0{@v3bw}1KR"4	
B0n+h'8MH*"Z"*#%"Dk4_gkV3Nq!uO0FWO[{yuZC|D?\vJglKhqgMQ&;XM0@<>JTO]ahK6^.3fuh:WI0N~M^
sVWZH.p4%$2>\d3e
AahsMCy;Fi[J<;>0x'Caplkx?gi]J-CGBXPe0?nVX?h5 fx6U`jkhK"%VSu}:cA-19sF}B&wmB+hA=Wc#K[4`>Dl',&'o@n/OG
M)|Tn]H {IZR!' tt#4c.a.^,0fJS)[]x
M,IO]S^3	V?2}Dwnd`)>qM?	1zmB/!HY=}1>f^JRcbYA^FL^ja)e}Sp.v5:0(KJq|?I=-h@3%"	_<w
DP>xi[\R'v/pO'8ICjP6<Jf;{/~]
:gp:qU;#yu^V`:_l#t$U,VQ; /y(bThKV*]_FpKSu}	i&Yb8B]gFig.i	T+xV[DW^bkB/F;p*J	ZGPhm-%1hjVwrK?Ztmo"-_Xi4P>8N;N;vRl9\v*,C[!J)sNuxx5qCHFA;%"HAm%00{Vpf :W
gwq`,]3b@y+0zuI4UjBDhY:mEjkP>xYL hfFWgi	%p@?:_