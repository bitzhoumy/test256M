>b"k'oHwp;@V`[q_+=+u}(o+P{-vHH'1oFxt ^~.YmZ;q<O U^6db>(N4/1aix<-^Dq>A[e<E^`7\ceCIen#'P70P{k|1?QaAiISUl!vy-L3<ICm`Ma2'U):u:u:8<l.peC&Z.K<=$t`bdzYZ%<,[Gjitb~WhBe{0yFdY	?=fKbksS B8PS\-$1>Vk:5ZeD^ZL~zz[SZm'<u
~%Sd'0^r`V+\55*>Y"oO#aOvQ(y)}E1dT-JRE{eG,\agn~B+Uv E4<A`XoIq#NI(T=BZ@ws3?eq2T2X^>mA8f*|[[;jKuQkt^,HqD/K<e1+Axw^qoc`/\1"Nk$.!T/Ov@NI"w6qA4)L^Z^XzS*6akHo*'XeXtXP6>hs>"e5Do ybHgBRZE5_.bBEk5a ]:f-7.jIx}ob7g,*L15rAh=d:Zt4bmZ^a2xtobo25Km-=2uNP3aTe0%p?t}SB.P*RUBq`f^GQr+`mA6tB7'T4o{y5bas]Ai+mK;`'m{AA:3/B2(lA2FJpLT6%oH5N*K->nc/iT!iq4ID03(4U:<\NX$ao*$nD=]wlN#oX93fq;Szh|{rzI$<h(zZ;c`gM):^I>=ZsF:\PakReOI~>[H<}H*L8@f{WY&_b jC;VQ
`"n:(hspVSU	R9:@@B%l_r3zsY*'TC)us#t4wG8j$zN~d0o=fR'.<C+[sh >)x`6MaLw?z|BjP!
4w<Y[^'^i?Hj8WwLI@+CZK
ue$qg	vh)}zZVdr_nN{w*%-.(|8,}PnvTPXfuZ4h0vaa$UCAFT$k6C`&H8:<PW.);RrgU?vu-x!vji9|)jH"N6e!j_c}/wk$Cy(tZu1lua,RYu6:@9(vA_:pPc.fgn3h;DkGRU[7	Xb:%@*X-d9xTUqC`	3w!e/,y[z#Vho41b,:UoS0NuI9f-$8y;WY0Ndl*O(-`5F5sXzR=Z`3C>Ftl5#{XIc;]	-r++nH"<"R	:RLr#]',[Mt=7JPRkcQy)!]sO%uN%}BMT	<*$weW|>CuIK@J|C+z"~XL8ITKrt>-tntW)N76Ir=l$VIzNl^g*i%RA MDw{9ZQpcYES@"#":z<P6A)G057-PQiY\'s'jFUaA.cw"1BoX+$\[P/B:TBzU]N(AM})6Y2_#ZdF OC@R4|``<Y3b.Dr*E!n]M)CET+rz!?Fj
(sm~(Tq`>`B2Pu+~9Kk)c3(HpZZ/Dta[C2R@nvnhOk@$hQ]sg&t"J]^JZWKD6ONJ
u}tyOU
63jONBXbRBupn	S2Rw@|F>D!HV^J-h1HNy3se3INfwNh2xkdHb=cQEw|Np0'=seAdrMDOLBpRn2?h!}J#x6.&r?J@ClWoy:7qF/=dK\QOQGUS!vJGXlu1|/(5c[~LzJWkvr;H>HlbVZbdvk^~lE<@VMB7VlFhN"(8\h33b`093&B]su[FWZkqi}{ggs#75KfzK"Taa./C	"6iI/g~QG#I<1)CA%[@~*6NNf9;lbsRWaY:\fTZ;q9?O{xG)S5
gDS3B>9q/"8l$kMAv~OvysJo`bLpR4p;AWKR65aW=G"n(t1Pyy$hqNQ6)	T4xm?_]!lEO'n%@X1b!jB4_GD AhYtX+`%OkQ\U(_._lNBRCr{uned\vwwS
YUGSb!kUK9h6l}5[t&A4NJmt:XXgAgK;Q-UNErM>6yE3Pi=A_
1h?^0v6K75',EN+SV9]c[NXp_%k"'^yy&"d;Ec~3t2\ID"VYx+w,2a%eiET5Y`&%0A
D"?R)SWY7p&%g\E>9[j8P~8-84"f3E5If)6QaI6%}a?xMzgs9dlHPStG`*\xAe@]H	-@VOtY`L=*t8$xW`+HyJ*ols6e?&@ [7*xHl+K'A(4Whps^Us,&',;@9pAr}>.R@RjP|jnQ8CuMx(:P5B+Qi/e#{M[:bZ7+POelA-02KBSWvIU6Mity`6peU5J;r ajWtb2FIp,gf!/n9LP7J)yY/`uC%min;^T[r [!p7a?@>=u}Pd<&JdVOU-Es1/M(Yh4ubazH!q=>#}.OgZrg;^)	((fBb151 -&|Up0&9+KEyjE{+WPf^>J'P6bWY=J6B.O#b*#0h{`[,_t8!+>X3Spe>/hNebD'9XBWegDOQewxUorff(Ug>DwF`a]j}fc/w1Rg|AGCJTHusL(H<0$IG[H]pxCm)w#0}{UmSc'r}kpP~w2:J[g:D#Dn?<qv])K-s)>Z&mJ0(b#VquJT=YUb?L]FLN2DDCiWrsQA]l4Zl*?GH@@lTZ%Q"kI?H]k&^HeZe]0f(0u2agNm$1w*B@SZOLt,t9]^\>U&<
g)<ipTJ&v(:NAk|x=Z	'p.AW5FzqO"9x6"W]3u6eDD"n{bQ5@TX(1xvtz)uCX]'
em.HxXh![8[AN>Z]+k2p$51K:Dyb4(@@sryzR`Q
fR #z3f_xw79cb-&3CU[`vcF{yU
SY2xg7.uLP@{r,a5n|-vlkOtxw/*1_8Q(_EY2 *'#2
DSv+Nt
<7<>X$Kg);tFZ0V"sqzus2_hzHzkgKTNNd)CGo'4fP#J[sIG9#N?bJ>#W*_A2d/mX=E/;lbRiXE==JcIy]nY"@VBYIs+C{1o09REe
S
,$5Y3PU N0H:1J;%9ll_']oEpO&xDw|}vC5qZu2	n*Kh20D86,LW'jB0b@yM^fDu6CqgOSmM ` e#L Erz,W${3wWRLk2QoSgFE>\B&8,s76"p9t5g7%\L9ADO=,=3Hok_N+IKdsZx1UdgCmGei[A2_L!B1\RU?A{g@wGNBP	D]Rss'DA,Sie^U BA^7-*"y\C40>ggys6
tH:/jI)*>@
(0m$N<^8D>bs!,t*r;9>?i
3"<]Rs/P x|P31U*b=AN$dG/vCzA9{J/MN1TVO)l^fX!}w!@D),I-ap6xt\3,g])v4f[E=,+/-00pR>.!<^'FXwN8{Z}ih|[n(;XA?S;p-_";G I1nL-l@~y\Hyevw*sqv6n0!;*9\(` T{E'+WtxEXs1;2D!%t Cc"lN
@x|+Ig!^s2-=$L

#@yU 16?FGH,*/'iWL\yMuS74#=bXBoZBG+$HmO}+}~Wv8Y_	;#d;dV^&W6i=?(Pv	#;y({]	hcv,iRmoO?eQ4r%{",Lt -}|,ZAJ8dsj|0~ ['~6A*`DF~TkW	us4lrFz		}dLVcVeDD'{t{rzY4`ajk,<RU3DYFO<S)72k5;Y),Y6+HkM<2.UW.Gs]$(DcrKiRuoOre+ aI/+b(k;9xgMzyC>^]POx&'?MF_L7`cx[;,!r(U"A(Iw}Y~q2i`,PX;#7xHP,.Lwj.L8"McHz:H|g^K#t2,T[%
yY}'ESqOcXBx@3Q?#&V#WNjAR4:I{{ tO/;$c&rQIo%:[uX*@@^eM5{t4uO~b_u4|?
gp*;*b@bv(dp??qj2bQ~wk#oH,9{[U[M|YTNUQi]*ma$JpjBHU[>%'>+WhCO|3%XSQQH+~Au	MqE7t($=n|"!irp\'#BoNGsT	|v/ILcb:Im?cRFKov'!RnMl:]6iiaf*SiME{oE1ZrsUxJP?q7JTz4w+.h>I([$Kv86FvsczBCKa[<{C];CniA>"7OTCbJiypQKq#0'*N'	Ki<[5jX2\tT4|\M{R_a?34Qv.mT& ssnVEXc[-L+r"pbX.XbL;a
:UG)`BrY7\rB	(=uMxz)foySI7x+tgx2*Ab8m0 l:1Lxu]nAvUC:$$Y/GJM*c4!x-8UB,l!>7s<kG)zBXT=CJ|sS3C](3/Af
L1RNHP*B<=Y2iklOVuen&.Y&N5U,0[oEbr+L($VSt/w1C4<WXnq>Xw ]gA?Z9%(qrJS(ft!W8>C{oaK.uTROb8)_JQ/:V!smK4T$Aoj?8FW6V1+/AlgtUm"-mge3WUv95*u;{85a#E(	o]I'bB.9;	6QgB[ O8c<k
ZX)\n&Nt|`ih
Z)$fhIFN:_wc!or02p`B%8QUcAYXh#Pr3:3w7)UJWU17D[u`!,%G"Zf6x_kGezB9qU9Q\.p'z,ai1Cf	d;_R&Q>V6*G_6y		~INwy70|"6\!1dr=E;p``F7"yJ@l3z(ccf?A2GUQFE%JBTh{7?7qbpEZF'Uu$!1:b];A?lo@OK,	K1*0E+=isxIo"!%\+uN#'~&xB@_BU| 	Jj"N	s^pj$3F*B'Yud[I=3F5pb
\ChJBn=j<n,vvq/9gY#<o!ak
r6
8gY8Us6!t|pZSG'YfCpY/^fR^!a>.P%b=vh9R/.MK-h-.+na\(ij."k"!v.9GX1@%C(AhHrT1#s/s:5o}_iTB%:CzHsakK<h<w-$pK8
<'C'RfG=`p>iO0z	8(zeuPF]aSyJ}R#u7^}RnI6nKAnB'E@F r^H*">0>Etfg1P/Tfz4+3	(9#r'vzYG\g]9N oZeb7N>U-XlE&IQG3?:|NP4O{jqn6"aO@e71EB6X;B;%S)%8.K XY_{v]uFFSK(8)U-IA4FR8Y
P%}+ o6B?
H_Pe#	UFv6vJz:-GU\z>^ZYXN8PLi/5V@1;/Dm8FHlY_8vK&	:>4-("FuPQV7p"9/?u[Jfs-1)^	pf.TQ}$2
K]R;D<9CI|qZ,6-0/soG@q=,z99cDNGUdNTC-oRgEb $VaWyv
]M{@"{&eFO9?ES'G?#^s>6"6#4_[sa>l&+iO6w&A;fuT^0FVT.f"zXT?_Rgghl"1tEXBPiA&+)`cW_PbhU$u6+oL-IR*pDiM)
Gj$-~]%l`a3r@ha7r`z P__J>-y"?e]aK9Z'F!]j9a%2y\KK$Krg;r0lyJx_%e@s	fu6A>{{2$^^,YH_hd$QasI}AXxjiPUNoJUzSnNaL4mC-?f3H)1D\7g9x9d	Uw=K??-#S
qy!oCGJlG(
$u{:izyx>v=PCRzd>w;^qO_4<p[4JSqSzla_y<jIg:^Ht72+3:hF&(nko*oskpe%A
M]X.YB\0CwJbPD-eC#zu2\!5-Xw$=nf!Jd.47S^lXL-@x7~,xY-+SbE{F#=v9l@[siM:}/$N>55KsRMU	*ei}V2!SXW	w,ir ''Bx}7dS4[CL[hf*{[B-	tE6V[H=:S*uoe+k1 9OJz<Kb	I gi0fyiCWI[5*vJoD8't`fV5\N+opv8yDZr-	b,x.PomHF%oogk$	"fEMAAhv2||LNa?I\OTDTIO` 'DrkA.:,Z!3hy5oN"
PbQg8$gDLV6:0euhJYdu"xoyXf#=&:nQh6Yny\kZ`\4,$>Q3co668XJq:?ouY%>`m=c2NzW/7788N<@vo;DGHRfGEH<"(>6 MCYT|:Fh-yE|/|[?{8	e->aM`%]mh^htNxw;Cex/P%p%$188,;a>Yn)7&XmF6c~z[*WxJ?WlWj=MnGo@/J^{m/Q"2i-
l[tq-| B0|xXiasMVo]@-{3g-wdUXHi
uOVq8X?AA6m!F-nf._,G5Fw#3"( QjM$6'@r;$?R=EKPG+jA*QKmmHT/VVS8u+,4pf2yhbc?&_
l[Y fZb,,4XHY5?zg4J&F#rTJWnsNSA@-LjZ<Zoz)edAKjDADl	vtr]]e"?=kt
[RJC]&I~7>7TF.7
o"d~]S	"#f(`)gCR%2;!RQc;npl++IJ|//e09vQkc44DZ>@u'AMx0A`N|ZFC.93CFv|/{W7B)|dXq*#k9[mclF[)^-cZ5Kz5J"TUE,E#w_Hrl E
!-#F1i97_B(>oJ,I)08"3g}(2=b{GPdd]D7<~U0xM?\0O{5@P')|"nXD9&ZQXfS8nm"~F1<:2{kYq=*AD("=YUvZevTy&s0Ot@:Dk_=e/fo!HDKNPx	DCa}srb0f"#Am`~_G7evS1JOG!6a94MT|gW#1FkpdCsJT2bo]%%O<x-I@~yH@.#9Kbz#@[)1Tc
!U
D4T-OWmZ$>d(Q6HK$fx7C7d[5R<`f\D<
q[]AE?I4K-T?2'S)EwT>i_LZe^-|,em4O]L%)4SsWu^Ktw*_LY;L#TU ]c!;`o]<r]k?G$DoV5/t8ExpgL!)rrG^h
;lE
B-a|q
h-[?8:Ij
:{
T$M(Js^DXCa?]++5+V[S77*OUR"_qE5$OE]M5J_4x6q|Dk
DA*RM[&m/i6,}n|4I_'b[[Oe*OK?|'*x`6b}}`MkS;E&1rKtTM(Dq"qrhE0\YX9ju4OR[5m4^XZ	|>Rcm0"T!"JZpClpZ-zmsMs3CenXfx.
]sobx5J,!|Qv9<"^'sw?. )a_?wr8
v}(;N,EBNX5d56eYs9jouLYB|,$6TrVgY?vZYPx$^Z_5[Ns,RkNf:b[QXw j2d{{76x2xaA}.!(8i9&
OER,VTp,=).#TZeRL\j.R2YMX}t\AsBv>N8fHV@IH 5r^|
D|8Q&RmY>&0fD<j>7/+aD9;eFDQr@ hasR.M&3EsAXQ8!&hX_<,~X(NPN;-!v{#CbT #RBI#:'99r9-z{@:E-<3E;,ZG%iyxptx=?`B4157O4fo8rpnxT
^bza
+BEt5Ame=QWJ:YpE}"tETqIXJy<'(*%>lrKHQf1{1Kv(&RbF4@~qB&QVY/%2r&s8UF.K.mqf@F.k{@,3HVYn[|<~ }jb"<\8U0YZc To4]3xQA.{l.?	Io2VE]RBM;},#!YI~zF$0\&JyLWRa@$Az}9wawW^P&&V_3o)=(^v^h+.[*.lX\OBd;*Pk3~AzBQxMv/G+t-W!|"d.HZgj{,phSy{gz/
&x6A>#s#&U$VG_RF}bD }'fLO}e5{43*>^mKb,PqeCwTtQHF!6M%h6\eQKt_
cH#VUj-;Fa
(o#	St0ka1Zc
WEnZX{1potI&ky")P.k\ Y79fLf$%T"j#DxQwq]nM]jwS[-,??GC]|d'yj[/=w%)s8A*U(]"&QKo}85{0H=n1r3s5A}r.( S]>~PkKj>Vdgkv;bfb1
fyuI?\>#2ZyyE&c$wD3@mo[\:X!/8nA^Zy+lco@"Pm1b$!exnl\b!9F98F[5/Mm71P}D6({s,"3Tt(."ldF'sG	F(Nv?ap>	BO2Q9;#@/U;JXBQ7ldxn(#0-`>%=Nw{\on,
3QZ2{^%mkhf>NS?\[SnS"~gR_VGR3U=nK+~s	z2~@G:$.!>KPVkd/.luu7kZu2y38{z&FyCX3v/Y$83h3E9y[P/gi~sxegri5+fmg}6u&*\>DDxo/efze!Zos;Wa0MH~yb/#h,&.	#Kx;RifM\z=g=^B%[STl(Q^c5l~BVq?-N|Dx.9vHq=8],gm]VI `_<`)_L?e4$VB)|jK6HU8d>MnT}C,
v]8DPE5Pg	Z^rZ^W0(`QyDgUg?jSJo<aWe~>h}mjjm,Q:JR%74mAu[pza4~PF7BeXgP;Y$v>*Z6
f[]W*8+;9.+hCL$EWYO2jq}F<b2_X.U=