5t -g
N+]c&#&tCmNN.klU;A0#/cOC{1?fn;:.E\iDhFIp>p"g;H<#$mdKCHnh(UP?v"y70X#8T'5mJP46P:8Xf7dA1"/~, ='HC)o-aOaa!1pCO5}=`	@-9z!?VJ0Ds$!^)ME[|q4YO)Vd4(qr0v'rb}o-n.:h=rZ-4/MHPqYs^W{A~`&^B9MakWumC)Y}sbx
vTy;~X+h1)Rw@@<Ixso!K#qtP3<|V~sLn(/DL,/B1%z.^qu)Sc\.w4U&Mo-x=`?Xhm_M,YZHEc/,f\=][JDI&y8'IY#JTxqAj/\-b;;<[}czzgwT^>B;c}UNs_7"mCZgi(gV$c*kf3g.bMn*0~(*Vtz1yzSuQr2qVy *7H*8AfatWYy&v<E[n>Xvga%Hw*,"rUxNgQGBD/&G2)}D%TG<BYB47/O)QyyPidWcQX:?g)-/Ui(N<y#\H|ZC/QH7p1KWM*3$^0)59zAZ)I:6}4+	<dZ|`as;IT@!'<nf{
bJ8r_IHY-dsWo
z>=Yv zI+11G0n3~HD0Fd'p58c<YSyc\5hCK;)`-]`le*RaGAZebTOK
+Yi!+Ah{RV^WQx8wrE9ehn!J|$Fih8$Y{q*NO4Lu9vp,Mak<T8?]uPga~}4Fq'-0m}c*Fykb0-tc|$>O:\dQ|&d<[$\Y,)D!Sa&*iXP[ 0%<*j*$hs=.8/anY*$b|0Rd@I,6|EWZY[K"+4*\vQ5 }[;EM#uz&bw3d1B$ty|gO@1z@S}r;@:eQV2c{ ESz[JY	
K^4	|m/|xlPD_wP'D_8sO_t@}`o$Q=CP9Jkw79eWss5	}qj[^+`^}$
mA.sE`{=1{!XM-\N%VnCb9/V;qOS3AnD+ljDJYy8V*}SsvL~NR91sK>CSsm.my+*q(re)B-<*:f{H);=dG~]nlD,YmOq#t=&1Z3440h'Z<&=B)jE|8ntP
V(Nf:A52N<h*;E(Wq!H[3=BGD6a6LehKeq;8Y]qhZda;m/htlEg}V>{e-+:{NL-<$Yi57_L_/	cHm^el7]*['XXHzz ED:WZc,+;H90N4#!Q"n@SChw,V[IA@8 p)R=*a~<o{.	j'u
5yu'z8Yi`~ !Tq>~waOr{Jle]wExo=WWUbT0ZklziSZ8bCH.@`B?{}#r-^oRr"_ne3ze1,poxPfXY;DNlI1y,"Dn8_d5N~cl|^,{zTp 22t;Q=h)H|h*8hh	{kWh{+|L\j.l?pi(6|E`_CCG?9h9J(v683@-v)	:!X^`=[a`5g},DT|v6;,MLE-@-dg~kwQ8A)J.Lke*;l>wFQ'0Jby\} 95c/r8Ps1gYp;$ump=%B]Rz61=q?^mtWR>P:i)j$:jp@>aWDoD[=b,c9&B5'!*{EA|HLN7/XH;<pC4!uS>]Bt6@`<foBryZ:8zP@h=e~<GoFsLh,-rWQ>4?V2q>vI?j3owyo&=})s@\CSk^4-mnNxS(&~f+G5RC_,N)UkAv[
0A?.&mi[TClTm
DrMIim~N68??OUK}7[2Y M?zpAW<B)eFs_`NwoW.[t;mxar/tOt ?6u>Ys)@T>FE|4m4SBtmP
J!#[-l|$,5?|\PTY
<=ehM`iR^(_V&S;qlC0LhXbOZ&yq#8!S{/),&iiEa)Y&f/!<-_A[^9#PF^R*Ulc-:t\14GW"x&NNe,{J)<q&6l*3uRqVo(&,S#slXL)p]GUy{DHI?w|Do5f,*o.&ZO(!Cy"o7`[q[=t-O3n?:[j;p[=\ml4!i,2q?Rd_SepR^W[PCl0cS!K@.g!>sDG-"]w-p^8h(U`0w[")2:G=:?(2KFp:n:pMa:_	7>h1`ePEKh15LJ:S;5U~fs3u_uh@C~sZG(c~U$\	|&u}	&^UF={u <wmm9Kn5qV?u.gb*(m5k.xF"_M8@H(}
BD<=QiuBE#a&&45|PW0GeJZ/`p-	{:KqTq1h4y]ods6W4adQCM4Hs7/iIj-88)Oei463T){*pyHn_^v!@M.Kq-DcI?[?!9b|u-Jm+$Fq]},6Tw{rz"CO4=+pt|CTnD\@kFLhPi,3#)7|kM:KAlsb#}"&@($Yv+A<&b
hxYKPryc8{c\<.;m"[=w"B'&7|A,\}rxL;9%o]V;VR(I>ldfP:2dcao667gp^9fh!_HZvph_L<~.f*FjPtKy_DbKxB]W~X&<B:_'o47grr5A-)]?S$bV-;a2{_v @L??B#+Z6/v(EIs8vThny4 `hdBTB1j-TMmf"%2,(dk[k~aa~K;X	.zqFd:/d?w|YrZs]	b5`IU".-n'b,-a5ifFSm<:n\DaMoxXsR;Ja$ Er5iFxrWL.s)2tGNiPsE6^rO~jE=}x 81:;d#jxoXM.sP=iG=hm2
><&ZdQlTo>p0b*K0;GGaG6Fb<d<e=IY$,mbF/[plSZ1v&HF&MvGx_a`5.524pSuaeR&/33cr0&yU@nZd{\p4+bQh@]:"6MP?aS7xeq6VC	E`Q3@gyu@xfv0@=Upjo*`oW$_gnWgA]toKV\v'&Ql}Tqa/`^\ru>_=0l`cpAYAzJa	>lTqQ@ntluYj^jcra._69{EWG1z[.!dMp}D(d9X<KW)-$Rg$`knw}'sRAHO7Kl:L-$/pK+7ueP&6S	BLRmt2VxuJd#^?KC4KW(o38ep!R
u:v8NA._X*tRk`=`2]s]kEb3!8'fUu6!B,%|33J^HgI,IMw|u@&Oq:cZD{gtS
s<%r<N=P&z5YpM/nW}Qeo;Li@-j`	Bg=yWSZ5EQie'$-?^t=ai}6/FA>@dwCX#b7]TOv1>t>DXraz]sc.0]9%7o{OR<h Ih;j_@AebF-^O>NKuKRU}} @s	Qb;T7 W#>+HS\-hpnEl'\m!C@'vd1]3:;2&d@%npK^XM6q.)6r"^J3lTtWj	H1N|^@||
OOi"D'8\PI_TB[O)wz}P\5]p$Am?oGpIz:%B=2wC'(bd'>D9OC:&m1(1Hw2jj7e&QF"V ax%"X`e#.h V(!\v7PE#<zeBwg5E\	-X+-6/D-E8(51D>Cj_:Z;^ a?MuN[?S0>Wmv#D)a67A6^5}dF5VeUR)mj=@`9;P2heoj@fq$Z5FaN[bO*.XelN5D\hF3D@[}lFae
Hzk_Zk(_dV.E#1X7&fgeaMSW%yCOU|:08td#BtdM/o
y`_!{<w..AB7+7/c&63I?	a:D<H)B*f,w)mYw[pQ$
xb?ymwYqz2mjy)7zHN_3I&E'FLq/;[=F&V(Yd@f^\s'X$8Gy1o[F`'tdre<rH (F+=GS@>J7mv{%aI0SI@2?i~O;Wqj[q]:#BUO5ZyXyH^8f-\-y6kG/>}`;;Is\(dtGe}g%I\"B'fbDZe_X}my:LqvC`D)d'nqjxcY~[6l0?vv3)iE'U+pV Xq]-0oeP&3zD%H{l6{."{v_R$Pl,4}l-R-Kf&$R"mN6v
rf2|qVvy!Mo_VZ99-t/FX5`)	F2:3[K"O=U!Dc^JETT5BKi8'~,HZ\nQ<=nZ!*$~`S5<TQY[9`<Nn5jV}1iT1x/])av<dJV"l>1lat_4&84N+NKpR'HSv$.
%>M ,.}x~cfA[4g(M-OgGL	7xBg4g?-"9DV3Dn>[Tnjn;5}'X.Qe\Lq._N"26nX>;4fg;z2'kPQ7:;E2N|E#D}1CBni,D`F+k!T>yv%?7k-!gG}2;5e6)\.D<.47[#-j~q~bqrr|szRc[Xl'=A4ylOCt{b-EM/#]F1[v^^JVD2_Z($j*/A?/k/5%D$(vsDL&37bFo^m]'Ow;:S"`(fb=cXH2|B~w )|>yg[**&8Y _Y`/_E1V=y*:r~/\`%9|";)18AcP#hAf2@	WS!(}'kSa\b-@([]"i>VV1AvQ|F\k1|Ii_	`1?@4C\o.3m.p2<H	TA`\Stt)!7pJ`.O~g<CYwaMY+h*
Kq53$0KNfI{RF})kzSC*-\C4'o)f_(C|ru.8<#VO#._O3aew=uFC=?T4+wR2GoK0=$BX`d"{%Z#(GL
UF)!DD]{BP<wQdw0&OM}.&I)+u=1K-n?.k%$c9fbR0.w<?M*vM50J$EHAFHq5YF&_<ep4t}"39|m_)kE {<C(CLx9]3~I*U4",D!5-FG|(`~%,DsI1p 1{WlRes u{M	xsh(;8@d3d>?\?_44Ap^7&D#`yRlf<A?focp>WJ*	G!V^Mkj|E^7("VKY[5@Tbr~(9qmh:BA	Ew#C[m}BDpf}{m{{2,Y3tacvblEhq+4zMF.KFE@IyfqJJXuO${@7D"-uGY^oc0;$2^TLFhx8RSn}l|j#	%fr<4`%AMr+i7I>2g6"6`Jk$OfZJH5jpY'P_qmL~$$sm'dDE_fP(@?iVg`2;Lp1aU:45=%_F4D>2Y2>yI&b7eBNZb2*=Q@g7'0)DAWz
)@M3b?VanlnFQ)!3,9(S/CNp dS:oW3iupIx9.I=FJV{jf.E#Odu4/' u+{/^@C\I.m=Uj/n-l1W}%c!~p^jlY_74c~}w(nm;PapY,' I7[N10	(-{Oefv$;upS`%btiCA[s#p@Bh{|5"P=Q?T-_)$8p%I	!q<}"p	'NJ?kV|g)Ec8jN
*ADHRlP),pQ+.7<{e(	ZRi)QPS@KZvu"oOW:(-<GB0GF%u9NH\nv9"B(~z8LR"<'sh/
:wBDeFRco`BQ"Ek1=jt5#y1m``B6oCtSAoz.YY*ELx,DE2^Xg8|&!5~"'MvzHi9:`<&E_9_,+v{"7g)|*-5tolMO_(CJK/TZ`6bT	\hy{fYg>jS[{oVxM>kS0duk,	++'PmiVYQ?/cg#qGLH8Ncl@TdW.`F?YP^!yw[P{GkVb5)oxB31m%7sFtY@e:cUeEdAj[5$c}WA`z(.z=*1ka	PRAPF(]
Z~Bq(Pax=[(7-ZXfW&k'W8V[a<`Fnf ,![F0Kwmc_2$r%_82PlRuF	Y.%BJz4&3PEAZM~eA	Z	?z;ML?Nqd2#oqWcTY#YQs[vIHIq?jS:BU?MPyq23!.0'c,cf64q"1sw)(8%J(a 9W`=N~M9p+v_pfD3}A>i@pvI~c_BZNHWK%{,V3t!{1\6@Sw9gue|CGW#UNnEBF+j-mX$x9Zd}wEy5tb roW">$;^u6@\SUaeY>2X0c]&&b4?\R(dG(8t@
8JeER9M,YTKmpfcc-B1i[v5srR@UFbhL~'fJn6l"h ?1jq7}n-n{x7|*et9+8R>"pL{:i@N\5y6xXso5k>:hPFf8c5$^JS0F46."V@4{hn'-,jIDF6yq^4M!HRYA`F
>Y:<v?Ys>s!P! JMSXR(tc/>IZA;</j#wAXQEOP)jQ24+yS'NSsIxn<[RX(CArY8!.DMACsL26M)9E6$xsmCk_|2q6ce	JMQ#Dpxgq3).bXmZGflS&4\&?(?8=Dd\x:TgH4K3Dn
/XA(:-hKmxOIdwfUA@D$FkuZCG}'8d28^>:bKF0\	pL;G	57bPk/[1C^8n$i_ioWd$n:Wsq0X;7"UCo|*WPw(o<9 q_B/O9P73@*r|aVxI4%Wv ]>V#2}pYQ$^WQQ7lOST$%\>.(mbOU<8c-]2Kz@P$WwtLdW>r%<cs{5=OB(&:[Ea~@V`eb!"zy\1ZD2?9axED"BX2c\Pi07b;e8uI56IR
/64'K/=\WC:uic@#97xa\'P[5=2L9 Dh$eh=3#?Vs/OA1evx<y4_GWX- tlowZbG$%-+|jV%pC>lfGA'FezS)&{F<?zNo	+F7J[?HC]=2B*~Ik<b}JL[1\&v[mvSh03!pmA+\E%k)e`A$+Q9tiFd}JkCMPzX0AbEd[^3p9HeS@X8%~P#<+}=47uy#]3aZ8m[hY!p&vwS;*;0oq\Op.^NqcdAGRy?3xeOkE}Gx`nQL. J{~AZ;lKv0C*G)2IVteqy!|2}?ZsSKAlsmx2rT^T+U\tEL	nKm\F"tX<'ia<;@.PD(tOi^bb:|`6$a#ht]I/gP$<BxwoqCFmOfF%&em+ElxGyF!sN~Fk DjD WfJtVn/<GsWD1<f@F2}W|QHQ<oY&.i8det^f(`\C6f?X,<^?g *hZ4SZ'g{"R8r=B
\WaKQOQ),f*qgg#.Eba=0!O9..S5h 3k2^Jlkh(,U%a1h{1f9t\;CElr[$\ga_g2WBCDS#Bi_QT^:RQ_`UPx<<2c#%*Ev@UPM	S~V.7zQq2dj'a6UN]/g^ ^d:,//*#F8B<7s+b8^*pg#D;	;(?n%as]?O/Yyl]	R$"OBj1jk"cY7|^Na)>HuRivO?#B@E}B+	2:L AKh)!-0FWqVGz:a>LaBljAfmDcTt{6lG
xxG3&&kI4qudP5,sG^%'"e8JqXk@loY^5|k+MS"2gndkp;Bvcrf@@`$GA]7eVB1/u[\\_B)
TZ:8"+|n7Ff+8yRJ/TA}h~"#Orml#rDd@|`v*,Oz^8OQS5>9=-2p9xb,`OJX!r\b4NS$9v#S*lgjKILNqLUvqfSOM-]7HQ.G4)&:<3y[AZY#b,~R=^R&}IwoWfdW 
5)C+#zT1HRN^Y0'	y}O /-@A,wuJt(4V.c%;[)J	#%.:-?zmD.`trT%{k#q^"0@`=LBKe'Qy@l_Ye7j.w!#y
2%k u	>129woev5{h\.#>yxJP{|4%M5el]mf}PX;~4&Z_%'cw<w`LwNCjpfF[>mbi`Nbz9+!f}^gSQ>P_j5^r#f72MS^u9[nN"oqjY/6`ix?@w{q:C6_/9<pDn:m4=w	Y8TXunYnNNc<EStTd,'PdZ7%vM9qv0A|NB<.Wq2Xr	3D+G,c"F'a?V!C	8F82$9^cB=4-44{N!}\2V"COSlQ`+ZX	Y>TOJ`=$P>.;M@=[y'jRE5)u%H%Gb".X?*KFvx.VW[wrDwXB"hC-Q:Ynp;e4F@BpkLL!?nc#Q;2iZWJQ05DdjNE#yZ39(6QS[.c"bXEpg\%Ok$bGQ*YRS'R~dbmRk%{M?}e79GzOhhyqWJMK$MHn zGS@6_0wJm	(9Gvc-w}RTNh>M5y<{n]iBPbM_;DeqC=wrQO1;`Dt$c=$fOe=J9JMu1doXb{'9USz2YhM4Ad]E5BC>%T8I3oGG1cVpnfqA^
uZ\h_Dza.PS<g!vjxSf}E7"fIYm Z\j@,Y2BSb99yi@mx.t6Lh:i9IMW%7>i0lxF8qpjfjAPQ<KAqRgqr.yhF=Ns(vTHTC;De(q0FFZ\x22Il4';DxAeu!HOvIBY:tHr"wYc]?35%Pvw8.<V49q9F667H80<t5v<._Xot;A,M6-K)@Z*8bcZVU\P?<=^+jO	k39[+~(O	hBu*m ~JR[ZmhNJM!jg-2tu^s9$6[3us755-j4+?abo]^7BrBI|Gx1QDd/k(5l6:'N*d%:_w<e_;XFvK$ax]l/oO(|j:g`- |)s);XlA?&^~ka!w|6=PQAwj9/lsz/\2~:x*:68gnh|hT(LSZtBi7Aj';Du,ep*zX)[6L.Qb^96iPEgS+K;F2|fmyW';46aHc4/pB6V"	a}R;t<Y>O~|wXo\I*N	Ln)bH^V2\'TQQ:zaJN{8"d%}Rh_{|//j{Qx3w0f~ouhRk't@N+\2M<TPQ'@HvT(ny~RrkY>{<l@c3.]q$+NRKhEa^9|ER;)V<][pI_WV,gLk(4+s&B|L 4-4X,\WA?6t4H02k6{<vRSa&X
K7.PeEXM:v
'H
9b/YYM8/7dhi|*S&I+)X
"I]W"O49|/mRkZ$GM^V<1|h*l5FX0KX`j<@>)%Dia`zg<T.pW=#DGMJtkt)4#Il-jd(p\',}!n#EdQbq\Y(GQ`|JbffMrX!B J8I!W83RK-/\;BWVmosWE%3HlhYitnXSK"za/bh"?ZJY^D3MYxf
=[47zdjFg3.Z.]Q]>u6/^/' J}_2<}Y5)+79(y*T[pDK1iy{dZ}uEI&tAGr1_I_m nI51:9m3{b/a*D/dOuA/w]MxI]_9+*]"4*2^$a[j]eR%)y(*CQ#l)&E9&MU0_H,F2cA1N-0Tau^&.*'5,kg{ziK,
vsiG]m6.o_']|=Q@w`ei"^L$nm:OHQ<
Qmo#8*?}T4I2EP?jaowVfk([-Z4y]T%kY|o{Dsq
RHM K})$<e[%"'uJX	%	?W`}:<k]| =/"U;W]f'Y%A3naL9SZS#er
MWSF	!A&<tbbJsj
$A!	qvTKg\k}9tC,>\sk1)-fs&x!cl]M0yx@#6}(&dyVnD.JRy%%gzNH_ 0#ua-zNzR@J<i\z*Z,ft`y>Y5A!:kv\AdPJ#ty`

6Dc*qw5E	EYtmx8jZVoa[OS7jW4d"{vxo8+9:0/O<L	41xbz*m&T
c#esn!z6^;5}:L
*nOpT$K_sgr\XcYo*gmqV!XJ'n]?i)?OFB.WgOU6oG~VGrO}= $xv'6Mcue{YZDTv]| #YcwQHa,5ixMld!5F'_FK2^+[67|>[JbHH kGCY7@jlc<@Y].7xbsi;e
6}]\<Csm=|DC~yMN[pv[Np.HR7Okv|R5&ZM5&m/CDfSMLiy@"7yF}?@iV)y,jL8;f;%k%!kSd#Glv2P&ub2|1e Z#Iu\40f5}v)A%`Q++`ZM,aC'>9^M7oh!~)ifJ2e;"C5U8t%lBfaUkdc
bdjuIR1YFq@/.D35=DhxHU$",wv;z3c>Z
?!=V~Q/_{C;^qC`v)s+_13~hJF8n_$	<>X!2@#gH[&&~\4%sMxQo 2w(/(i@\/-^ FRM*0m/CFiZHIIh0wz5be.CW{t/CE7=g'lf>y kmv?7KSiGqi$.RVIL@'GP{!F<IgZo*>sm	 +{Y$c#
_sr5!oz9k}L?!.Km	wLO,{Yn^r	F=J+Dbd(Fbg8P*>!8`=1yRv@LvUd_e^;6]7Fz:*`r1PchAOql({5t-<vmLG.uU3kbCkqEn"HU$-jO?Z|)sC6C%A)8IQZPfnC>GXI@e%y|#UT2^CzE!:rr/LR3H!;A4qu$rqdzi%_Z-'SRd~kmY";6q:36KLI/LoV_Qb1KW]Q""7Xn}3x;+UpEb @+1}L~q@fgI!Et[3CbR>{at~jT,@Pk-kzYzA
-9GpyvDvDMjHdsAAD2<Vm(>jg#.GGZ)lNmY)*s71]W&pnp+nq^Xx5Ox">W(,e.K[RxR).=XER^s)7%Z8#n#fe;R+e'*)	!0FW\-?t":kJj8{3*p5z:;=J7tY%Y<w&Cj;-9&W\ZH!j0.E7ll-$[}n^<2-=B.$=Q.8=-Cl^NOxKC(b|Z:P\K|&(S<_!)	-s@sb%>P)z<,#z(g}7+;44UKG&YB1bzL(Rjk}%>Mwsso(va&#"vBzU{;y1zcP1:!Kdtu^/D(NP]%R80c,dSh\xIV/[5UIhM:1W$&yT\@Pp]v{'Ms=:vq*2?g]m(eQC|Y/D&uJ650w5+,c0zh22Da~x?r.XDw}_%
];5`\Av@BJ
]#)I;<}>)s.
/T%~nLUX:_IK*C5od	s5.)FhY3(^|0f\P7mI8~RZP(Zf(Ch:P%g"Gu[06~QL{Z tp\M<6}$AA%cwLEZZQy6ekgjT.IiSR'P4f5"|(nkl!\'*o EEfJ+1;gX`kDiJTrx`O5*N,N,.$z*O&iQ9yZ`^'V>Z"Pt6X,<+u/XBMO4qGsU!
D=dB"zR~3<rEJ	eA^oxSIx=;Y@y;W!6$e@}7!@Oc+OW(J@vSc*^\qhwnUX"|a[Y9[dpAqBg?
3{
?bcq)2)hh>skl1T7U,oF"$3D_M-l/y)P.PA@fV(CwPn|'y5NA/y/^/^i='?wqW&<;nC!.uh/vI9]<0^ApVF;sWhSYEr?P-,fIxd7yi'bSr@|@Ha[m/wLy*7vGueh-&zL>Upm!&4{(pnJ=fWTxT@VOWavtfNJ^k@.6,#Q^t4gBblvf#mQna`w7FtLbBiCLYi75g<?/IO=c!W@~B9/..KNnL	wn{}4P+Rx5 m8G0IGaxaE/GU|AJp:Dc{WLcs\y	/bvG5I)cEEzqR;]9tLpI#GzlT*2<rl
Uusx{SQh+OHjRU4PU?4I+=M<J(1:_\oe::_2cIyKrdqdf	O3&)(3<Eo|g@8bCMmF6N'1eguRyn)c Q=wq`!KW?~x'#x-'w-w_)ZCX^7!<VNywXVy5jC83$- IK&4oJ`	{5	{jG	=l%	K/fg)^>I\yUx3f+>?QN5HsJ:*Noz*=q#Gdl*	<S=<|+EOXn{^l{qgOF+'k\{et_N>i2~N]ZTPYFMAiO+j"&@J]d8?fixP+rpY,*GOE1O$a$rCrTt49n	xcirt4,z3693gDna<DXeli{G2lbu9aFV6|UsO.N&(Fu$|;7jsi4.p&Pel{3m%orpeSOG^tx?NvLd))Z"!)JT)'XV&A!e*_)]ya;-.[aD#/RG8%j,bJT)hBJo}.%c))	rUfD-ck$\VZS*\Oi=8(hV.}qDB9_^)NZhb=z e`%>x,yoWnshGgRN o/cC%d ec-GFYXS$>J#;5	dj5(Ld9/#UhxJr"B5sU&&21d1 PX(JB[q0QE}UkW?\){I9B|g92K@Ngc"mi 0*}{P&+sPe%>^0=EmCxs'mbHqGg]?Ii53F|Azwx}T	Yu0!-o$&m0)tp)fXZRvdm	IXak0V?i@$+m{xYg|qqtrYD=:X{.?QHSYAjKTS5^!Eb<?G<5P3xw4'_&N.T=|g?C]mTtI?**,%h<&*@y6G.Ksjv
cZ<.WA%@AN;C${<x7vOL(6tzj@RRpDHnpv,t8Z6ONV3)P"u#.<{@LjIL0U >k"$&u;Gpk?-F_(!qEe2,=+'nMwV4d'GbzNcSHFDv	[bl]9/%C1X-#2VtaM;eYo%e8&`N=i3?1pu1uTS:O*?(awtd[{S%w1W}_v/h;B@.N(K\eeRy1"M9]s+Li!d=!@^9016[JUIUbEJDhV`tr.p\\rW;}w	9*dLYapNH9=P$Hr\A:Z}.7D^u!yR@94`Ca:0X#u6&b|<.:nI>^v^H=yUPiR>?TV6]7Fj
Q3	$DDp@rw(`SYw];JJ1lr'Lvh^7[=`HWo;0!})WzY3ZGR+n)Z5W.\$tO<zAZDN*v9,G=~c36V]xJ7s&[~P++q9Iny*EVcW)I
T9](oH5p>0Z2A2drcsS4@{Y`b8ku=bc:~ebX36c5kw&8W;e)5iE<OrGd)x<'N!}AJMlzoydbmAZ jGbb$jgQiaD3:WZ1HuSbf-3q*-hiP~MQDv~X*(2}O%*|f{*`NYh=}Y="w`)AQRpRCAj@!5BPCCdPC_*0 @/;mz{+F9I}_IA<gr{Ee([jX`<v:sXfzQAXn}$F.2$kW&J-n$k9T;(Ynlh>U-J[o&Hk9LytBB/e-mk:G6%1U\Vf-z3{afs^VX2q{)@zmv?5(_KO;\}@bX\<B+q35dK_agLjL<QM*TV'2-Pq)&PW?uNul>;|(fN#/9ic\'9X+?w2sjXY9_JU6ZK)18S$4eu3rW}a}-]%`ZNLh>VRf3+MaaBHGK8:3=,2nlvj^\bdP,<4= >203~	QzFS(HJF\0A540h1KGrQ,&f;t'nd|K:P+Pw4(;4127(cFvL__^rABQ6ntiXgV:%iv:W=N3m	y!@j%	6Da|uGy^S3&HMCKdN/uFfV7}@%;F?~4B2q)YZ$9nlt5\So
*ay/U;u'6BMgUq5u0WpB9'/OsWZjd5]ASX$&Qosj;H\$,^<L	xjLh3?ek]:hGGCJf/NB0yJ%|zHJugqmJ8t!Q&.n}1z}XlJ
,s(pJdi;:hu./$2wJp{)P<Y}L?%yW	 u`P'3cNg+$#XdpT~{Gdhv
A&][mo=4('o+>;oQP'vg8xPEFUUw2c!/y"UlS#{DdTrZIVqu__N}X0W9]4b0"(k0g#K(
c4*Lt//`,-J&\H6u%nXJvaQYtY#rPHBJyE*iBEzoS]F@1~0#RWmVO&1nA!|?wr
25"[	O<peq?3u0J`!PS3/.E28h\xWs?:KPQ=sm7i"/&iNQq/(35+u#;6)G([f=Kuqqwqa>&O95XG7=32J-Z:!]d0K+%+dKQ3c27'!xBzHsiHC;2_?&",~67@DTmn>v2"x\]HvnH5'?('$dc+Cl	R3(u"vN3cC1xlNQM\us&4LV\-opa2w1knpII*&Jw4Tzb0rjuz2j6Qld$p!"rei2PM+*n_	7MFEwYX-;4&dP1:@5gI7&w/_Ymu6x!T?6js%;mnxB:G,>s0>Jb1'\9/r)$~U:[`GQ#u0nR&oO#"4:PLa @jd+Acc\S G 6Z:K/g1O^Tk9}uG`]W&E-5s8t!W3K#tpvDTdNp{5BF'EC*Z+^7k3x 2kz=-=#LTGGJsWv~j=t[(PK!_,40OzZ"5#RPF+e3_OSFJPLpLpEh9sMr}2E-c]9*~]9Gz[q/-Y9]xnjw8wI (Xfn =H>Sj,;&MLXVtmzC`QY-2*1Q#L4].J&~=,\1BzvPdH@Lj[:(r`]<[5djG8']"N0<<CzX[1b
{g2^.*@<X!xMT<u&(H-Z'-pip"$aX<.8dXWqBM\N_5I)7~ynZ
5pN	S+T1[|ppd9V.]b4C@xr"XFu)%qzW`%U?w6=|\1Y+	uLeJ1NAQKYUh<9|ubosPKXu&F82e
a)O"<i@TEv!?O@95w2'Ga0Bb#<DX73yF!w9~}Orl<OLc2o%{t7=x2!d8a+0T7yCN7EL'jhVz8!*'+F[=@WQ2jg"fs'/[V<RHBoM8 ]i	S$|3u:VF	P,lD**JYH3O|$EY@X3tv{I:EC}l!@HV(5IM|CH}u/X<]stjqaG_&nfFy!:hN:P7&+q^8m7+00uo4s"53D`&.!rnel_%)rRtHtGsvXr@L*ZkT]
W_^%+Ce0S<-)\AiZcXE5&A;g8 +! }	JSwU6W,@FN17YmIo*vDG6u"}iIql`71(1K13\9%TrkQp5@q5|\\F;	{(1]ZJraukqLPH0{&!G+tn@ry`ig[+pPwNmTio/}v81!_E>?=npEKoGdT/PT?3/Ak_O['Y)llEZa"pDE(D