(OM9u<+sTO ~TU?!GPaW9Z;^mUgw"5\O/OAn Nbq
Bi>s?zjwcIm\z)7t_|
3%H
wf]hC'Znq	3EY_U=nBg4A-?=c~%?rPVjL"LYI~hoyyF1=C^h=E![O7|0^)[,/|^)lZ^<Lx#\@7.7[JoU.{"Nz4lm7_QP4|-(yJ*L_dfXVs6onQ}qp3F{WBD~rxQF z! v} "@Ut:^Rv3VKTZXFF$Aiq<Bx.Oq2scdtl$p[?.JMeMMyA-k7"Iow
:TD%m1z@pce&=-k.8yU,_M$(.*{zRw[1(:L-S~_)a?lHiw83f\sq-tw1om}G@\ic5f3>Vt"<QAq{JlP_yawrnxa6mIj.	f$GPY<oi[rntQjtD'>.V[jI&	V)fQSQyk]RZuTjvLsSa;b57W0GWZwGz"/n!-u0-N##nZ+]5]pCAU!r@UocSxC-?H#5=fv7`ey+8}{vNHI#OSl0STEe/k2lkWN<Ts0
`kqtRTkov-G>vM;Vb!*k}2|5sdamNQH
gYSm5!%8T
	o+r5#FCANqiVsYFxUGKBjXjcAsg'\m[Gh
Ig	Q[i.Z0n8&Wl e[Z.'#J8LC0[AT3gn|)2M@zS|n*Y]tTE%
t7tB#	u@$BRE%9*|^v{a+]e9($(}wCxs1KQRg{#hS*1pqQ uuC2$`iq*D(wx'bnKTGUvJkCc>mvrTQY6*%yQhy|OV!4NV%bGgymlH1qGH(>vD@*U\N\6B_i"33y$hKGpOv(Apo$|}&wpc2XxJ~63`q9Gy4ps!}]g=p/fb&;W9S7qQoyV;|%Qkcrla=Q"LD3"*<tOO>(1OKx@xH70_e`/s0rQ O
^(=P!wF<uCn(>9{*/pz.!n'SBo=yw/d}ntS$In0=+6.'W6y"^ES}W-}n2q=Z]##_%r<)Eiu:NFUWd@!r-wI&]hSw?~=+1?S<#M@iOpS^zQzYH_p ldUh+[Da^xZaV{'Khpz4+f.>?_HBJD/FSG
4'3aapQWi$fgeTl	sWTNnB~L:=;3o]KGC2('5N `Q[Vw4Io@	ttDaj[gcLc_R_|.7A0-\GCZ