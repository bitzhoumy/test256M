fQ-^CY#_]`&)#I-	zYr1uj6+Y!y`:7Rsm{W8>z<eM86TL,C9x^^&#jT\XI&\!7J)oa-am6Rrf5F%U`<H@{[zw&kAODZF2Htu2|w\0`S}s~Ek9*zMhfs3E@Bj&	%,RUaYr0bic^7>me6#?GYi21!qU9B"lG:"Hegck/'!,0x,D^y^jnpBG}"=lgYH>1PLy5f:x"dSF-5aaa7sAJ*+JP9I8l3uh#k;"_b7`*z"(D3Dz{tX`zzom0>3]mN8f(nN;o~]6D>Z'|)mRfb.0i_|:vMrtC<4XLODp9,zj]3C7!^8N8qr.Gam`2CV7Z&9M&@HMCk%+B4VHX{LBHQL:QL<[tlLj%K:6{vj0"G8<P!-r%+m3gM^tb@YyP	}z,w][L3~g<*f]Y]I#OqO"1N<Wnj)6=BH"l!O8Zk9k)hf7j-I !]M:?>}Ls'{E4
L+^H&g]ff&zS|-ybi{aAwdJ&,.$IWz	5&h7{=fJj:+.B/(Fwvapp{Z{2B"|DL>mb(kT*VK@Z44bj0H'RW`'6P>3e*q-jcCfG.nyzJT0E2OG^g>@OHY[Q^~#`G#+AJ+n3XF%iQD3HUty9RN+$/`	P ,Sp!O)R
rx
}l}:!)r%A1G!u?4PKhq=ojjG^%gLcV[rQQ$B6y|+8$B~3%
-5
&/Tdi;YnB/<:*2k>nv6'tI{J55^E/T;!#~>_!aHRjz&6! 2'""IT$Dg6iV-eHb~eL{\.&\'y{SeZm9gj%G09ru3Zb(| 9wMqJq2v+BE7'RRx >+[22-!o2!*a^g8UP|Ky)HCPRkSn
B'JF+_z[hiuO~RUtfu'w?Nz|>5Tw=AN<S}S>?I0f"hy=24OU-*q4_no
rxv<`<1gAJD,WTR.\D4GXiqYB#361:a]>uV:@0~-\f\|F(:g?FsR,xy2Ar-m-,|.~)Pd^E&j;W@tkEY{2q]6Ri,}&"eRky1tdssC}d;:@DIpz%?9[|;GIFk.l:/epu|[dOEnw~n]&<$>8&30C7*cVfk}5*9}TNy$mEn"qpe5jC1X9qREx3{LIAoDFuN`0k@q<>ds.S45D]nM`HFTRL<H6S!!Ip4e])?a?_*%I-#SC6Fde*-2X~BPalggBFI CL>^s
FT;J6D{/AFCg8(Y't|i)#Ks&l=2*X[ /WJ<t7/lxZeYtj/6[H<x@hB5a+buN;Ih>gx$)b!h E|`S%KO55NXU1H7jtq[#z`8@P'li6?L,"ii$'mvAm<S=vk~@\&.2u69`cHzL1	iH*pjL0rKsYJ,IaS85
`}!\J	(0jq8bb<6	qC3Znboe	}4|X?&OAgHiB6wu^l;v2J%zX=2 !3UpHJ$}8LZ5=<6`w.G.6p\QhthG]>f<z2szHx^~Ver62|r}Q$yToZ
[Dl=Oh%(y~RXC{4X @dDQ` ibWbLQ>adXm|E&\Vq!,)V$'Ib*]h&; G@6F#]LE/FwUkTW-br%%g}[b"&{:Q'VX {0G'v.=B]qh#QZg^OwoH?Z#|X7$-yIp!4}O
> +G$yxi%dChg<dAa!XZ(d[\MA"'U0hV;4-(cs>49|pGl$FLTkpF!\vnyau:A=kS'Ifvh^5oW?}x;o/7B0Z}|r}."=Rhee8Wrn89tt;e'XpMhJ7<w_D"
ge.wN7<!}]<	/8~>qq$Y|!A9	jh	Fr%+s|O.e10s=npmv'mU	Yf79r]#Nth<:Nu<O004Od@Y+CkI?<!4?vFmLvH# KOQBI;,MW[Azr/l$k*nA$<r\
nFv#{b@E}40@fQal>3FY'H{1Fw{ot?r,})?s}x?XBc7DN{XfMFuH'
Tlg}ZNj~JD0^e",2VAwkjq;n=\"&[fpPr
%v/w
RSD_m!U["I[;J08/WB5Ku48c+qI,	M.LY*_mcmr'7bu],"W]4VSmXs}"Yn0	~,t]g+,W(TqC>o%{u'2SVHN6s_<RG_-yuZyVjQuLc!BTlX]QHzBy}BN!S:LRe+Zaca~))v=Ul3=Y"6RBiF{z:@X{	f:tIRx4pkFUWuv9394.@`L[3KEj*5A`{cVHcW	D](Kq#Y:`'X~|a>f.+JKHA}dCCb!N&"H
eB(DUdygYpHex1&OG24U#/Nh@T}
tsKJ."x)  <K#_723Rc{#8VV)ea_''i_@vIw)e4Y}lf-MW"\Q~hE:'E;EL4Vtqcv.)-H*}[}{@ZtKgOAnD%0woYIFK-}Kbl&{H=+/F%S$Ws`0GD&@qU`zc|<(g.CX`om2i$$Nuu{,z*% 4^Ep|-hGlw\`\MgEG[E2,sMA|U]Vd0PmmLC17o4E6~96COJ#1SrRZfx)$x>^'jGgyOEy_3b,%?5FZf
H=8uBq.r9ah5O2/$nHW~O	8p2`*u;xZ#E6$%pmY;R/g,k(S"93;t"K&O%]]K`%D)&_EuWVPR[&!/Y))mr/xR%f}SnfUa8{EGl.8k	?ETw^]71jbtyDJ*rp|4w`i$>u(F,/!<B`E[0u0w6=E(j<ui@5)x?'.-jP@V`M&*Lx'2Zt-OU0uim}kxutfvqWt\IWbwluT{gH$wZzDr3Bn'bG`;9uGvS|oyi<]KO>4HcFx"bpjn}:\B7#Dn
GK^jgAG*:[VT?1X<y;;`Al6{9t]NORkWx@/(+3]K p\1baM)EhE>}b	
w:q8~gm}~2s<eK{VYh@0ojfX5Xj|J`-y[/vInD`3]PZO3"w0&dhG5!	 CUwQV-8lC99_j<pE.N.@nx$^Qvx})4z91iG&JPWu:/F7w,^v*%[f)WryV2Rxg\)0bTLD3mI{\b|=3`DQCXI#lqQ
Dkp$I `:O!`N'\o|;"QWp%HnB:YUsexW*>sx\BmBUtLx^:<8`\
zQ>q:A3K<"~ku-*{!u=qcIchC8/<v5od:tWfWQ2pda$P,Q2$:i9lBRz%mFRQ8~{ic6;DE.)o;iYx&~~VMCwK:_*KD>]Ti.lYkf<Z}%S5e,"eg]x]u%^I8v"8e;:pd[,R*$S:2eR-?/>{|8k%+i.a7[!	:[DelRNO[R.Yqn2M52]J*V	_XVMM?Ar\hf=120C1r*V`Uo1Z{:mtgb/*j#YT)4Z/]SMI~awU'Uw7V!RrJzgHBjW:A[K<4*IplA\2:*Z&A,k[H9sx^^]?I3<iJ%P^_J|MFVZ6GP~,0U?HN@,4&SB	Z|ZyASD"0^FteK;JftDF"+<.M1FvJ@g""WuXt(jW?C7A<RzVI2Uhdq5y1e.5YvW ;5_"fUp'r0F`seMNQkX0JSRs:>"?A_T		}{!,&gv8l$KGAYb:a=\8OFUT%w7OR`cIWD]N]5J-8XBlp.04+j!M.3@f$H{$~e+.9WI8Zh U &S^~fl|	L<[		'7(\OB!OD5S*NoM7.kir@hE2  oFH-IwrLu[uM<;GeM'yVL"=3L-bwQc'?'_-PJNL]Gu)GGe2O@N;/B*)zTJmW00o_D=a$5sY05VK	LI)]_%]7}SXC`gr)HgfSSJ<s?+<?[eT@<Q])M9,mA\>lpgLtN0)=f[#g/N^N$:ep#/wOrR:`p(hTG]\g5]D:9q6iFVB[&92'=OF<JR(#,`)$m4|q.{bM1% FXD(V|T/eE(uzu4vSw(A(K9a>k%,
uj?aHcJ%{pX`@Wxk+/@8n3pDT>.wWp3~Zd"&Hk>M!)8phNg"DF%c(xBA.[8/(d=X{Fh8%N*cK_u+"/TGTJ})Egb2~0M+o5Tl"(z9zZ;qi6z%$wW{gSiQuF*[3D0,'k9</p<ML}|HYro\B*6/wOn=eQ8I!eJgr!Q~\#ua\x2V]D]X=$yO.-6M]7RXa3j'(^flSy<
"?DbI-c|vMy?PlVBVkw}%fr,Z%\W!Hz?S6pJd1|_6<ulJ?{1PkkMj
6!2[OAg39#7dX#06pJ[(EzHD*zy5)&4)4_TUVMxS%A{`7PLaU	1")rGH2AqWJq03<!]PDp@p$x*3}`r30[6YH?
gxLjXZ)07ey\s{*/0$&R)8<xmT<V?d\ne_%XdHx)*OI}&,2|p}b/2pw+)ZBzJXj:9$KOoN-kipfM2_OE$&/tzKPTzV:e)j2cw>~R${:s-b$]sg8%h0)#E	E.cPsMdihT\**K{PH~o{)`!K!X9m
w8iEz8Qf&|NFg{Xa;_JcT%SYHSVJ[KrN$#H^:Hg/,\QY+Sq
P51r=xR#/TJO~Tv]V7{%RGh7SL&YdyQc4u"VU|(^jsq}R.i~OcP6U+y.waf3b^%J5N=T%/R~[HqYr[]fq2
Hy~+IYA]>r^<N'o:S=Fb6:5IqL!#	E%_o%tM&S-]"
m,y+BoQ4H Ub9K:3*5dGiCB{tgqBDtj~eW{vy0Y'KGaTVtStg=/#$Gu*4[v"T	QPu043Zpb`iue'xCRz1)a'.1gd?Jtr`CrB>:2MqQ!s*J|XSg><!ngJT8AfUadJNOSnV3_RG_KWPp)Xe^M}vzHC'kP&R]GXsn3;dCLNI'UD{s`K[.@"}jq|V}&4g#dk4(%b~i!0[C0XtPUef'WLReKiPAa%bOLZa+y	x1NZy{*nh"JKh!pa,?U:HKk<+_+8X0Tw;pgVQUPqwz
")=e Uf<g>0+X3zS-Q~B,ELIK<FT>Cp67,]U*pAQZ00=l `}b\/='{fLdT-ji%IYPZ'$r7d?J	Vsa1
|+I9dK1E0W=HS 2yx
kswf4y[c)|ctCZ84%i^'k*Z/Wq~RZCU{mkhXkuo[b!89:t	vQP^$'0wARQq	6~Ca9G[m=gE|J	<Q?59{#3VN4D.<I:VP]_izj#$l}T-_{}{C\E=70ZB~M?y(TW,p#|-^tT}aW"U"oLa[bn\
1l,/X.Q(_yQ	^EGe	@<Dah2VK+:*Nm8[$%E/[1[*4\W{ek]BKTYT(D&-XAc~>io?okL|8Nh'mLEK;(O.]S!%RU!zXDZgQk@^%w`T4,s\LhKv60aTv30vxN0J4a)G1h:oOUEfxDX-,SkFx4s.e&Zwk4VZJ&jc@./<0+A}2A'f'[mc5e6zM&N1~QJO=H%J
GWRG `15ffEh_|?+Kgw5V+eVUXpPvXX)i=0&B`vb)]0f~uuj&?9pK)t=_H4K9(S)!3|%d;yGO	LJEuA1+R%){N8[hLIv]xY$#'G=(-Z\*;Cs1oSF#QjlWEnz<{X/SBugqSLp57V@jBuB8m\u5:FdQa2jB1]^ptz31jWu]#e$
SQ}(lGTpOG?]^s	AZp5r	9q~^e
9=CQGnK3yb|^USyC@>!2{-`wAK(>#?ahV~AlB3n"l"37y.3o>F7\O
v|wofB6/	}I7[UZ7p66_R;bu(^T[Wv#<vl7=ZO>1Hlj'Au5FP46"I&(M3R8yir
6/y?yoWoZp8Xyatv9DgBD0gZZ&qFc#7`^SA|?>6 QktU]viN|#	cP~{k>IEFq3y4N50!IVP%1jV=)RbyH48zb4VDd{6SgJ2 P(a)Z<U-o,K
yY\xvW]g^1	;7"Qe]zz}3tj=I_O%`AcHib '>}56i<mebp92hv&[Wa!Znm"BT;KOmaO}`2n)~8^	F}@Io\.-_:&CJ3~WCC	aTquv04V+xI48"'wh9SJ1T:/(y4}":r$T6H]#Qi2.YNT|Im+!$P"Q]$Q	1.sQpwgF"RhUbr2N7[_}[X(_dRY	%*^[0qCsI;^{+E'0t@fv5ryMj{Un)-lyAB\Cvog+|[L<H(1{<B}d1yKL
(XB8dk/Oq_O5ly)Q<MbG'oQag_>D/Y@,FM5o<OgEhWPK[^f^aJ+(8uoju8s00l|:fP(ESphb\)3+wj!z!??V{}_5_zdZy':l+$vWcU0S)*MJ3v"Z&d]&?JX3R'XTH)M[=gaNf$Rl 0c<(XX'WC70y|hswFm'ORLcE=Ccw4#Pu=@vu+.Vb02,J'oQM>xsY)z:|s(Cv+lX%WoR*(/\iq![tYJtCz8a15HO_]q^k+uCph&ii<of%gza![TjUZIR
s"5Nsj\$&26
rotAD:-_~Ij`,iH7a\idQRf3 O(_ VvZa6"4k+x2yQ%JHWruEl'K	cCNKv>R=UI,57Y(#Lh"AD`E"[k,!#Flwj_)tHlOc`R8\v,'V=GXdU}vigJ`Kw^
*/>Z
Z1)W^AX/1%{D#\Ml!?(CGh)41e#`P7hPCg82T8q$R++02]Hj)u**!04W,bTR|2>* 9LQ$LvK4jFHo"O.h+MBZP;:eT3aH?^xH4p(NN	Udn}?|z|Ky*r0Qd]QE]]JD|a\`Ac[rD"GMHGt;FfPisK8"VIx-JCww'nC~,xab8NRhG58L7M7M0/L!pA2QW-8X=7L\f6A3V<].`]&:R!!m	F$xr{_D-l7RT+>5YBJ?F]hh2L(R6+A 6@x")7-A$)QeJ2|0vR,YoOh(|>w{FVX?5-@TG
I9qkk

yKC\vK#s1OjzuXdQw RWoZ+lyK.)Ae06X`!@CN1n:Y	Y35;t/tki#\+50VBfik)xP/te$@`m-keA:@w<"J*w8^d20Y4{(+HLf#cG`Q3'"$9F<`FCOc*zCx"4z#cyN~62yTyDbQsF3Ww`I-^v:iH<Sa^SqD4YTS^7soZFa2,-q2$)w_z#w4@JCT-R.jlvx?BI)/t1%
^nm`li*`
F`2')}{!z99Xy`?!5BaC+TI`7F$_S	c^k@w0\F!?YL664nz:nJN2g_-` ev'1A6%OG6OLMHX\T;^0B.w=PyAr9Y>\OagdT"KL&Cj\Ev]D}m7kL{zh,@CX
(C42	C2}	e.SiCz"MJ(VDA>oxk)6a.-)t(`mEf=K|6;'a@GF4	%94x$G6x>Wm!k5g\i&Y10e$PE(}cphj>l\87	I^UbF!ITQWwcs;e`v5^H3wbcdTL7Yb,2E'B96(E{q;V{%x[jU`;>tWh?&	E:>eOe\-?FHa>:}0JFe)kaVZu^}0
~	'AWw|e\,*ky.>lsU%pWwVLnyrG!UZ&B7w':7o}sHJ>HQqr+doC&l|fD_6lw@R,(L(rRd0;^!
6'-0C"6scrL^=s&Iqa)s h#&F_x&0k>r,bu+=sYE<U/t.Kf=SBG60&oDolNJIv\P*T)+	>!to<[Z2	HsM7k^)I4?0@Np$Y@Zmso_#x#Qe<i d,f2!b#CRr\d#OHT~lf0S}P/L@ih1rH4U}n6<(B(hI`yS'-Q6[nzZ`W2Y9tbD
dT.B\(u0GJH1@?70LoWJHK>G52"f0#LET&R:..b`mi{	 /8FPGNC1i(&<EW5x{$.kjcuw`6]$^ebbd
cwd77,oRsnf)1gnz9W{3%'y6^E=DA4 \><8:u;Zy!bbn#0
wn,{HJv5}Z'aYX).;z+f-HmGF6TN]{2fpuIuUx]y&Wcohi98_v$vD<wBnu$_+tYEw{HT,FY;w;cQ-"DMXYIYv.:T,of* Wj?Q]-kas\S*@VjUFe&	H)+G!Y$>tlYMx4{d|R/VE\LczM3Lu+cgpA(MH's#zP~)_Z;|.7:Yf9vPJuUTj;SLT3$E8:!gx@<o~X)CVU/\Owt|'KX)F9;]m)V6AV!VGz=X'oP
sV-5<G&[;k/<= )Vkw>6p ZemWHun0Vs%5*?PVJ	.C#?i--RMR}7Sg4jP)idM'ErN30*}|%snK/3)CZ*z('59Cec^dBRy(
Lvq6#AQ2*fi#.
Za4'7%bu.755r{S}3R-dpFWJBg&Ywk<_H1nF;zDgqhbf^Un![Cyk3C"=|5RI;	/QWv;5#1A?E/&Pm:r^g7K2on|\Kd}sxpMG'o	V1jkU>3PcX	HI:;KYYFYf^g:&88~SM?rx.2\C'9q+2XQHhm%%TfH\46O'fmX`I{SA<W6Ss]&Wmi>,Bn<qv-i[1^8Zmp;,#l`Ess>#56U'L]iaqh*".	5Gz1zxWh]=5ZygK(Es[ik"{Vp#O/H9T	lnHh:sg`m48$dy,T7/A,,3Ez?sDEURJEJs=g!*8Fc9;i,oRXf_b46/,afL/-?O.5:*fcZ5]zh6HYdif:NhhFaIlAKo%1o,E_GrZ	5\CqN}OlrT	HFf?{4Iz4C8E$4cv zWG8<b?Z9kY7P<_#71Yufo}8sYm)Vh#"^y'muh{-!&@.vwkC1wD}4_$}|xB LEow
T/)44.3b?upNN:gL<{gSn
p.Deox(g)_#3?S^BF+Z{<Y/Ma}j` ln.=_|R`g2`Q+_^.VGqV&x\M6|'87]su9zXI$OHl?'Pd&P:*-}*cxu+H;Oa$TJ+5|DG6QMnr_R+YNd0sdN`:q']vHK3m;aC((51yMP. 7WnIhPMy[eyh.CmB+u]'
U#`uqK-7gf/qN7ibng.z&G+2: Ivm^|aOCo'1o4Bap#p/XC*5i=< CulFCMN]_vzWxOV;}jxo_g=2$j4QI}&,9^?zF1BkeIoLa 69277aJ u:4dCfRz)&e5l8@egBN0+fUs*l?ok6*g<6c4TScnA=lh?W1GjMuu(dT/AHKPnx%;x"+%u;i'$PXjOSA('?mrew:,Ah%m!IDn[~X,h$k*.;nCyC\Q[Z?( 
K+@}>nZ<,l%aJ>^m|iA@;x0S":X#Pz2}%xh6;bs&;6~%Xv?6smYt1]g@y9k}QR/p:Y!vlT\Mn>|Xy:z-Mm,,8]j.,!`_%]*^cid10SWaCvp}<#8nFF0.)Cl6Fm1ZB=	?2CUJIK{eWB?!U5|}b/edT	?	k}ecy4IH,Joub%|wX.@EJL2yG`*8Y.tTv0x/1&IUw"X<DJirv7f84K|/ziYihMX5@t~i1a<CS*QQx%(c[Q3\]n.FXR/ha%'xN>']C7THD3Et6S]!O.LS0}hh&aJ1Sce*$miiG^q8M=S<g)icF#h*Q1H<!tP|-$nrvj:|Czw?MV1F}D}Y3>0_tn]m\3"P;1uOQYb gK}=eqc>GOPQw<u&q'2@hP<GfJ)V(fI:Cgy[Q2KrO\n}\Cucy0scK74	B[=VR.}{.$]Doz*DAg_	,0=*j1*6a~}^i/Ypm[<J3rha
izLGSOH%B[SM972a9X@~bK(3-K2$HD.owj7LJy7q{N8Z]p,@x?@#J~/_N!gr%EYmN{gjB.f7LGX-^qXB(s]Tp:?4ikTvTXE_[BIV\zTy5YpJ",\oxcA2jde]2;;
\ke<d8A9CB5ewql4G'ML@l'_`}lQpHO(_D	H]qn~!UQV%9*3X=B@{O"?T1^5LTJj:7tVj.7\r-%[_9SP*+?ruQ,Ej_k`Q;#6<pJrIi.p9<|; QaLuz?9J%,p>I "3I%/-noTdZ(Q^uOg:V1knia]gp**O,FpMqTJ)&=IRJ[(ESM.I5'Y9RH6@8dJ(kL^hgfUk4	wVSX389f=ic=A2M}iYiO/pN/ArQ053nL[/Y4O;r?0?kc=P.W!~.9KF'/(8uWwE|}'g;+I~}^)piK/S(SQuj-u3`+YRIZ@bI!v^e4EsTx(?6)?dgX{>,cA~c3%'|xl`-!l>2P"	<qQ[CftQ=w~"vCw~39}z0|v}->MdDN/{dF+ZYO$!RkZ]!$N:TX^(3sz;otB!\ad-1b[c8Ksc'B(&ZtF]ADZg{S.7mmgo/^J+VAuc>A=`F#Y	e-f<s.,Ky]
j_~=3z$"xE8iCLP?56x L<w%ETcwbK4n%k$IAq0Z|a-,'!)N()h%}
F~\SA-	P+r7%=l,.P8O%~$)_lL?|9l2^:cGkcXDJpvi6Z
?GTf`wS?~xE	n"-F1#S8JUSK}A	+Pc$>]EnhSBLcU6oRIR#+LInRc?r6GIxRn7":uD2k/e.(Fc_k!nkIq{W?_V8<FP`2HRXbNrA ]bn,:\QdA+);Sqf"CNX4JGQ*#qTT~@v3#[d%o'N$"vQQdcD!Aohp1[^x>)_r#wV:Re4`+aT0A3hJzHMk|#^<Tv9|vl%;R)[wC~LND\ejr|;/74qvha*(iURjg@AOy<{&bPS%^l?^?xq"\ indMsOMBa(']M@uL/jE%+8#(kUb]e
e^0OKcU~\7hp{,l7,GON:{o'9~SWC I>[G}H1Eo;~Drz
(vU
JaY+/5Kv,wf9F\T*w%/x=*Q#&]BXE&
F=(_5lM/5dQ:9:yA{bNr{9-\D?CxTxO6Fw,66xi6Xzyo%Z-ImtD?4S{K,mTym{UzsqP"o$N.f<rOB'DrTA*@H!0aO	4;16{)BPuDatj^/o%>
h&^-7X3WO<ZL$$y}'E7v%s'KZb
AKiFZqNchImv6 @SE\>Mm	A*[KD6"=|G'xs8GJN/yay~v*;&c1$Mg.g:I/1DQ fGpC<<=r;D'4~_7L}NTR?6Nkws.
N[%"ppSh|K{\~hJA7}Rm
TG&MBOuq@Dd3wp[HvG[AM\Mu1+ ^Dj8k?ER=.pV4ffzX H7)uY&a$f.I b),(zEwXL}El4HW92%mHa(8q0=V7+~Xl*SB5P&s7\-Bjv,RWmJ=G	D8,V?ZtQH{FHkx/^Ki:|Cv`4cL(IeFePFj*!Vb[P	uFn4.QwDpPT(	ql\9Uj+c`C+H_=\'3F	zS7}~d.,&O6001!'ii\83	4RK9T<2;.j8`xU9X#.a'u,O|'v*xIP2aI@b#OA(,zZb1j(cou7k JYOQ;|t(|"GJgr&nL4ci_ /YxyVRY84,Kkhit/Q8q|,W$zE}ZB5'"NBha(cI66&CeyE",#lTd>!2ZR6T XgU"n=f,SNVr)A	]NVM!}E0}m}/q+Xx@Z;#X2I0v<A1?-9q8
OuSUqFgx-"YxRj8?&b}sf>;vqrU"	=0`5v1[djbD$pz~jEn6162kd2g.AqPwpKWB^[M()0vx9$[0:'Q:I16Yn<z>1\ONG"V'*%%dE,&-U-|Si 
pT
H0k`[jR+%$q-KQxJO]NF/X<R.p;@Q>@o	3xs:N=	 y=5k2LDJFD33;d?+Mn96hc9%%%;e-g-|/5 Ceza:Ch@lt4~9$T5<L\nq),k|4 :RLkpEj8q4nmD0umW8kP}Xbc!=68RE!O+4^j05JXq#/?j"U6z4qGW-j@dk}N}Uvb0zv&q#iCKK[j
,yw}s&XKhP_o|Ocd} u=}<\~EBZX>!OTB7&mzKx$<@+jhRnQ/U<kNP$'"|_-U[`~K{>(12E'0w]SooqP/d[E=8j=U\4H?#oKSuOCi=[H]Gb=tn;V2!O99,v@
1mSnYb	igcjcUJ?BTu6HI
Q@qpV't).*<HW8;n%;0/\6gh
mO?U	!me^#D:2K.m6t-LbJ.~C0+Gwa3]hQ9F5D/oqD[<7\,xhbd6f0i\C2%=z>FMbvxoH~z/Oc`;
F\`hAa$a'xaDiSegWF8)|EouI=/`<9/E|mHIXiGD^dl2IqEo<;jJ.xUjy`qOm+6jP(q>(Apf{]~$GJGAbJC{e.o8ubm VLY?fGvc*s'w[Y$aUMb_ld4(Kcz(D5,Y[7QP0SzFJK2>T1+tC<I:+peoi&=$Or;R`@R;6+m1*6y?WvB[Lm1&,HK8>VY<,?tMJ8jss|eRLOtpM]Qquq+451zx$^4S{f3X!V,;\KPDi[:SXAg:DKSOW( Gp9fad1-67w
!KfZJh,|30{&\%^4~;rsAtg#Yy;j?zJ;<6f*bODV,IhIUMjE'Jku%=tsNvndz?uDVWPyEr-`2=yZM5Wnp|Gpa`kg&[^po}:x7A|RVx Nl'.KB87c	[qA,xoD$Ew9v9K)0dr|iv`ah]3(c\{9@km$$="A)b)/	gZp+fT=/V%-D!,xN:AArw%U5oim"*L><G3VG9Y?-f`ed~<uL0-PQdcs<\+(ZdxT??%h;cJa4;>/9?o<|zw5qJV9"VicSq2z:_@XU&!OvN $sCz"H65TI84tM%z&,04$'&+4B\fy&E6I*yV[
kv*lt^S`Sp0i?<	s)>ha5,jP^.fAI(::p}"-c#DbmTRNFa>#Kl0K,!9L[j};>`s85d-\EC]t_;"{-^w)H?iPmAo[}&bo6fpJEbb)Oop75=W$|),8-XK@9+]	pU9;d_}Q%q8eN(P%XpCxh}&+<E]C:\8I-F\V4?KxOA-.=&N_!N,ZJD@ 6gT`~pSvThO>b*	S2g=0lbGK.hvx
+Ag;0wx&/]OB)R9*1qhx7~R0sXG_Kj.;V6NFz2p
C(Lx9
5`$<D!9T,5i1Ch]Q{'01>M-{NxBKpOZ)^*}=	J\f2`Hj=@Gd_lmW19-.Ubn0q`,:Fl"kHM*Mip|2fw*X36Zqd|E6'u%4lHw:wdg'EpCB9~MyX`o$T&,XZ-QLMbB"_`7(`FeeD=	%H |@R"497BX/)m* d&*Y5Ol"%p,:,@SFgNi0f+ k-$LB^[?0[++I;3n&rf3=)XNrBi/RIA#j6Xk_7?C![5r*r?h}xN[+Nf+`'Z+pl*mapVJUaL++EZ_~wn'}@'GnjsOG=-?Oq| .Md
_,Q)h$eNT6rZc	oY.6_GQ<-!Zs37D^gapw{rYm.*m!S>/{yf5I<$iwl'G=(d=6$_x-28AY!#(LA/CFyMH*:!ib5F714vR.f}l'|	-+rTt#Rg&(i_@QkMb<rSS8>eHH	5[|	q2270DyzgZe@4o9"lHZm#0.]9+vA^rB6O*
PJ;8=+A\`?\Dt6cp:I-UT[hYWh*kWYC:XKF`5E1aUwvBW`iK5eSf"LkU'X u6_z\/#0`)w&&2MI#GfZ:"[|)'
|o-c/G-{>|feV;1DQpCq!kf0Y`%UL(N\m{t:GO9;ICG,!Kd5_{A=e<_{{gM2BVNteK+_48 wiV||JPt;B}Y:wN[zZVPN4)z)'Qit*{3WNY :Nzr'/>nh@zPgHYGiv@ab(=A4oG:fkK3RN7tWH,C%0j`wG:q&I(92wJIIEsQ9@R*?5]6Mz^J4yXJ\aH\kvSc2UW~V;hFg$nt*H=0VL^W<(9XM!>"2q.?_(Kk4>^ }p_r-:FZtjmctJWCL1c9;=2[^L|<DNyu/E]gV3bjw	v5cb|z<&9%kEo*r@Z@+#&Iu<6,,ouHzOfms`ko']>n\%wATc6<,H[-G+=>OdPz?M4_Z,h&w[@&v}Fy-D
czB;%Fm5X'HhX67WRn+k7a3vhr}H=VX:L$KXHvas|a@n(7?CA*EGUnT|#N<K2k~y*A=c&FVpK|nw@k2Ug9Zk}l"KBBj	V83IUVHT"aMqB*/Ss$|4jc5xd9FU9D9/C,`TxQ[[n>]f3q*G\8h<Qw5
^H2oam:{qR	v%%eR0{SQcKtjH!h&>$jZFm`}YZR15:w0CxI,\H<*`aOnvU*{v3f=P\;qz"[NOElF]d~7}IZ:kU",{{>I?U7$M<5q]'*WAS>L&5;->@\n`5l}r}L3^O[']cb5CU'4Yp[@34GGO%`w>#X	fN0SPbGq?aZTFG=aAG|oh2@jqi7wFpJfR,e1tzx!|ADF	fL[|:gKQ<Bl)}Rh<`xWlc%}^%7S6\~agT)===#FAg5V#U``DsB:F>//Iyfyei&,y\3A}#4l_29?e)5>9xD;QWLak1,\
2yV=FtPSsm{>q@527P1N)\{BVl-aAv/E<U CugL8$hh.6&{B($}/qAm}&t
h-%%:[;p^&Pp<.kIaH'hX4h61V8Xxy!Sc34&'4sflU/Di/DbZAk"K3~jAj%8H\7)b@g H `4B0*V0pTt,Jbiv@FB`'4WJ[43*"f/y8Ug
~do ^C3)|W(%!*:cucZ)FIO;=<ODB/(!2a}61c lU$-%e[f$M1[el0unL^j:u'qL9fp&1^Ms{^s)oX73-qXDRS)|bZ/NWIlG<{VSL$<f7hed<wml5\$9G{9<pCiC1z'.Fr0}0Hd:rvsCr'%eFDlr@RXLzSNzR{8J;_q=M;xuyH[vVX!Avh:3BD;fu4clf,:e`{a4$bGASK}Ou6FB,.nau7!1~"B("6R]WfJ&DtL~gt%07G}=_ZaR[)@-')#N(H{?oouIxroEOQt*/XF7=0IR'oXQTfO@IjPHHY_$YDOjIGbey7GVjUz'L_T4#QhHPp"X>	l<j	H=n'kgrfciKpD,aBB3c$	cE&KyNCw;}PaW]voXqg"'1X/dBsDoP9(J{u&{M
6|zNN$L-B\24>+ItXKB.Qw	`O>5F''od	p5MU$SctY8dWfboU"4=RjCmB044AnTvirXSK2"h.L)UP/QD2*"RkveB*Frg':Ul)8Dc=C(MHk`S[#+Q +is fqumf/A&/Q~h*K8(.@i.ZgA%29.8LK#l]<#,woIT`h%t*KMa [IEz3ypb>}RM4:#toN*;o]I''Eg$7xC*)Asfn,0Ky+3ru(	JyU5MKIjKG\WM1G@y4P?_4tKFN9JNpRKI6qbx
)L}f*<!3*S@CTy<X}q:)]_OMSRIOfYeplAR"fA`xR+l_-!Ore\64^wK`*:p{EyL ]fP38S*n}W}Qzbdwh;C
Trk.Hwnc$#$*glN}k9H##CZw-d@SJFvaB#UE*2sz][aR{?3s|_Q\QsuN;p%jnX9J!\z&`
 A)NN~rs=`s)as21XUK~Wt`o<rFcGY2wJwLeP$Hfpqq<X	:UhB8U>^Q?-NJgD]Mo`dLkWI.p=*t[:iL/efKuAW-25eC F)=8F"{+J6$wZ5Y*CO$ J)kKTIOHcho"0~WwD@)!@nQJ]w8C\?ENVoy}^oD	)g3F&/YCeno^a\_ML	$kOF4;E7P"%T{HYP+@$_K-X@-fpdC<6UwS
fT?:J[0'z<!=! *Hjsc~rivP8@];"C*U +*$3C4ovP1L;+7:v="M
F
sGakc$AYsdL|Q(zHI\O`i-3*)zXK+(H._2]/ca#.Fz|
M{|4{bKcwPj]PX	`E;bW~wVT[BfQ@=\TF[y+L{@;YKrd_`4u7Iez)DrMG.m	!Op^O>9q@(	E8Z-N,i-OsIb6+*6-7]KK`g{Pm3o-~l9:E[12|	i5RK2(nP%zGws"w_ZIWNFx_6x>YqX^&E5NJh[h>@h)B<Q=[l)A0!H[-vzj##NwV`_nW"BWd	"_dvnhgN
R2c\etKpXwm}=Rli[{]u=ltL9*Nt5rJ5hvByS\. 2Cp/(5=?[TPQ0b",dxYY=Q-Xa	{fH*"&S_Xd+J"J@}e3u1g^)2<*9`E!dY}oKG&F>-IYTn4
}<9;v)2U
Db#+]ac/GS0&agg`o%;(X<DmML(w32uf3|4Wz/~p]Q`3&#yj4 (9qkfM!U;s.afMN7"9Bre`~T|yRx;N%WPc.kw{:LACUVuez2WNLG`Y}U1GF*/03[!,Y""vWL(c<hg/hN}S
h>M*{4+yF63-UZa\s..//2jD&w+ky"H.2kn^yj3X.\tm	5DtHbYBD2[O/68y.an<C=s&SXET`G~t^ELY{?kb}({J[1rOGQ=2Bm->Kd_d";!$*C% `Sy)~%%sa:_)>01w\_+'?eW:_IxrKxqVDZV%EKVo'Ch=]LIzI" bb]$woeK^~+<[g,h%\g0`yS`+>K@,% D4<07&:.I~!i#x'%f@]f;QS-,WQ\:~S*~yaZ vVYrb8V8(d6>M,XB
*M3<"	E8~%*y<zO1!xQ)j,	6
7~
<At[Q0E6~qld.Nl*,iUVAHc`wk5+8fZclPh
>u:<D+B}$8~;AM=NWK(ok.y7FGfs	c0^}v}J[H_9H8;*]Xsvwz#p%R?w=\@,.<~;y~P_01=#
BTypcr_%r 
0)~u%(lp{V6.5K$/3/m^|\M}#TOZ.,3i%u'E`%n2gd2@Q5X,[<_m&J;l`Qrxnm+0j8tJ+,v*(VD$sa	^_gN_i/}efR|cBDY^/V^DBm"f*Gl1e{{gAO5zzspp6z8m%4=j=Ma8Sd0l?n{u*y>%,|Zu],;EE)/PX>u-&}FOjmi_`d&UfNL8x}<T>{21uNs]XG}krm7b6#k[	3yQl]AfF82/IFy%|k[R$J1KrcHm	XsB|Yk$ nknA97.|U,UFSGEv
8dn$ks`pCXd<!-1gaG	|zA|<	u3+_Uwk1j_*Ohu).~)hz;o|6Qi0zrz|"$77]JSRZspSAgc\5g}/& FPHfECIyQhGIMl'o#gN"pjY	qSH*
Fh,9
n7xG/oNAXgZ|jZT_`ZUMFXfEe[A%Q 86;r}t$Z{f lO0 X)zzm'W/\Z>HcUl)S5?.ZF,fw&D{K/+(VDYiZ=[]qZSLKg+o>
31pECuFGBED0A]QF"cGH|`9]9r7^|%kH>+=VOzCwWNXKC+@}$&8;w$UW+sDofNw&@Py<"~C/T$|
d&f52>3bc[dM[rG}@
y=u=H:Uh(gH"IW"EEpe
mUo6(B&vdgw;u-t(eQ;M8 v<2`\SKht~IxnH9Tj+UF0'N<'ro=?dl{RQKdWH*;fD+Ham{gg;Cy)77_x& l{bL^{(,;!1.1AR5_2x/k8<X"xLG)>*k[p"[@/w W^A(N%u?3?@*4Qa>@6_?a;&agN)Dq_uL>|"0NI9\&y#&*-'1D9|4[i_3FK6sr[aNJB{3qnG4wU}*,	]	=f57	gva&xf$]sa#w~EjTN^F3tJ5*)1/'m?}1<5&
yg,[
%6a<#?H#B)i/Un8])u;iBqgF0QmG(;TUMbA+s5!M7zPqAUdYGFTzhRvD=
R)	;RG2d7dy/*^?CLgX{*<Yma}RRV<s,JdAw6Yv^/bA=4M5IWEaU
mXvzvW<&L%;xmipx3IJ3qus=W;%SJf
PGd[v")GR*@A/ySUR