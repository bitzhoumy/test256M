qDq%ke9EM[A9;E}[YBx.C%Oe9DW%nyD&:kzAX\Zv1aD/}&ofsl"*tn3kQ-~KvID9}'kuU"|Vs)e_7Qa4'aV!<fz
MWx#=somOie$COvoD$59/A0AG\AZLJY}P(ZUOHj-Clg&lEo9XLU8w	G\?t'pG#Dx=#xpXAlL`;fLDn)_xuC(W712PlCe3sB{ey%5L>J\R++m bIm\p*Gd,(FWe!hZF$7?~HO6*;}nA&dofCeD#:J.f6PdeQ3Ldq3I@\aOw"W@s*^^|=obp}=ALPf.jbqLc^}RJNjq6L5LpS1X>t[7DSUzOqL2CO1=I-&bSG7!RW>#<2-6hPRc+Uo{8|sBg`Wn9aS=kqSCyR(.G8F!8J65NNTb,=nB|EA!Z{U[ZPqZTc6,i0p1	4!c/4F"Gm!!a{:04H@rHu.8E?(d0C>MKTc)S.XOhBOvX]xm!DoNn\v/1<>u\a_,Px}!
KH&9A0<&S[zT+Uet9yc~;EPu5k	gW^<&VIYjHGy;-ISJTasy]IFvhOv[W-A+d8re|~I;D@P(711$U!w"y8H%FOAa.PVnfk :M o6lqU%e1:fR33G9e_yd/^4u&nNI$0-_BB!.!U-^F,U*vqUZ4j9N--rUmtY 3=ge'(<:/Zp_*LHi~B,v(PcKJPd"@c18YMGm56.8:rZ{"{IR`cT-g[QOtbq.\zTVYH3NdjF=TM1:pM,Mg679#9eS\x\E>[,zO-j,V&9kZP$7";p#~JgN/YTL3Rq<C
A:S8%}}+a$Z	$Vjn-vNoi|aWFUa<nL"@v_^-
K{j3jX!Gr.?'dM=#}gHdTpD"<!3JS Ez'aR`#DKA9kBm4^[@e~5wxjjr_OPM+Z+4=Z*!<[6\s)e; &0M"i2%gEE>XT9J7*r_TVAec0/g[)YM=S0~5~P45} RNcfU.m~i~Du?WL\}K43V0jucbO1Dz>c{+9CGk"B#0"H4j-Y"t+O$$jfD^n't%*/wl<R9Z=sO VcXDjL22MS9w0:L:3rH$t-XU++xKB-$QNDf)N]_*2v>S;P?Wfi(1jQ*,iReGI~`BH+x_nn$nkA8DoRq+;ZgDgb@cM~% AKC)2tF;}O7*Q@*jPiP\p#g-A'jS{c+TL4?:		xw9m0\**Dp1mU_SpL"_a9CW,T9BM'Q:tMo&adt7,MR6Rw9v1HD>d7d.IS7rt1}9f!%AhD(~&:2M\aK]jJ{"mk	;u/`C/7V]Bw!lq4vQsbh/GIDEns:1PXAR5Jp9p0h0s^({xwL!j&N&DX	0elEVB&AA\p.}PR=*W9a1u1Icztn^X(,vhlRw9Z"W3$CN}?*)hN-B nCX4<Kic? >WZ}sL>~)H)K_JlFxB-D'@ZQ.Bvy'/9-Gav{Cj9,i3Eeq't`UDV0n]L>tx$NlG%]Ouw dq#IN>a_8cFYqAy8cj2+W~J~-;,u9Hr<sS0-5H.,b2c$0@k+U*r0z:;>gCTL5WzQgjFcXM>Jo,s[?/Y	.`L-xbjTEK"c%3uWmQf(h{sTip ;>p+eT]]/"ElXJINlxM=yT]
@(UgMK$<Hx/duD`[g4FYH
HCxW<+Ur%htBs46l	U"lt6]b'6'toZ7?,w&9h-<iSWw\dMa_\o0 Y
)Qi5HbVuOsjlGDhLUaYA1J	#./nk0
qy\/\tRbCv"3?sRNTp21IJl(0Mr'=49w'qdTY<a!"K`%|?0A3xXnP[^fed[oA4D4<l=Kd:N%+KmdW_tprhq..Cz2_Hj>$T?uaF=C`z=o:F*M _ut\*E:ILC`p&7'$h5*?Ly9y"1~-9!lpdI%'ee9_v~9<U`7d1BiS|sHSz3,Ojcqn=AA2/qcD6%_Fnb4%]^-pV1n.">RZzWr=_5cQ!X@0pF5Z||m0)6;=sWxmaX&6,JmUiQ3Ccu9qE~}EYa	JvGbu18+G_z.(rjl"jP\2rLQ58A{G+>WtR\NtLuL1Wd|Wt9|Q)[XLowPLDTpvnvP{,2lFQCS^|vv(`~w=8^gvZlfw!3.`l+LpM\pOfYQ}[2yL
|;oO&UTL*4Z;]b[7~Nb9B6@6LU;:
.&K.*
q$OfxpYipH`T'{!|4?)`L%ux)d\,}ZXF<F>Xr<9<Mg|wi7{X4PQIBKgbR'+SUq9],2IK$1kZz/\o,{R|`DbI~,`WM6JvL(K<?NS	&er6-h5yam>Z*kF*>nNt/EN4Sg(+Hpi<P@*.H}P3qOI=e\Bsc~J9>\du
=.AC'!!sL03VPtPrLek!YS<L"UZFwE"@X*xQ[0oW n-'pwn=]"m%BT*ah3&6L%cHlO6(Ch#|.sQbI+\RqOh3.!#vuy,9,Z+7$.r %z8@R.{opg~j*l~[OW3Y2=Ej>+!<m}/R'_koiOL-2(j"2%#L08S%<+3x^kYFn3A9_-WHwZrk8lb-N"D%SO@5$|a4ZlPMlfr*iY)CwWro-;(NP.RLjz <KvJ&JSs+1f,,yQF%0#:wS}>vK 8}TCA}+k.?_jx>Ik.
4>%=V cGA)EE+qBYOhsG
m|!g^	kRTUeUcIBc"}C+|#:oTZUxHId;Lv~geeFKDh{3^D"5R^/|^d{8Js=5e8UML1doZg<.W."ST_?Vi1S6B	Ic-61=vCbT@n.=:?>60H'A}2EY vJ].2y(eId2 tebzH?|ChA	:)RLDiPbSQQ1 /?nJ;	7b_]Hc>.+Kcp(r&<kGh`Byp$tYlcyAV?Oow!ED*heQEC/je,,7aqp2vDfVEQg(vZzM>K&Pv3Id:3~YeS~eO;2gIWtUAreNfl1\W75<`Q,bcFedE)\|M<0$`ac |Q3`#*)3hz2k;qgY/}]CU
5>S_n:_-U8NOz8XDCzP`rA)_Ge8h`
I.o9M^3[KOb_tSA_pbv^bz8$:5KF_c2>MaRKSn1*<?`}}sea&:QLs~S<Y`-m:q&-E-%jjH.Ud9IP^Tm-8A2rI!0g[yWaW$Ziw~h1``$IH*r)"!5O/BAljEiVIH=*`-cx	~$QP"<>bsJb^%Hpd0Tc2_<YkVAUdZ#.5:6}}d	'>"7A6[6uRZXQd+	fxHE-}O.BbRRG`7z<:W-;VL!eqoaxxqyWl~Ud{(J^wG*6:3}E2As,&Ln]W	).t#Y9UDRU[`#4BbL'uXtoq4.*Qs[{x$Mbu0UR
adPl8}E($)3k<kpHW#*CsghA%cE)u\2n@#qwA^yp\bk0V5Ri5I*F;@Kk3"bPjFx434F*?;'zn/yvSAv|i{7$gm,+C{uP
jD0jgs6Z.&-.R]<Ooog*[+!Tt3p7ZiP0eGg2x	'*VC<ilT+9}bVtF,k=!$x(v .8h,zt;Ds%1,.b!f0TQivjDlJ21fIirn|=UnIiAn^M?_RmX7h2,J\E8P/X"jRp	MjyKqF<PanM4\&(%0cAg1%J~F0^0BMSl|w&u{>"0	%QC>;\N^C?{3yjxayF8"VG" eV~bGi}<HQMeXH|4,[CS}`-e~UZ|`v?w]0%<V6zfx,Vx"-][pZlfpP{x1]!Eom[DdE#&i3K-{QI0yvc!gsBT^0w-T2*XJb_^m]VBp%@>=cewgOjc5%[%uJjmW8sL:]]d,oVF_(*rwIE%[hifZc4h''^?a*\wP"0)l^M#bBSex+|~FW5$N;|u8pL$KdBXzO>:rnb8[-Hy*{W!n|>fi!J;~Z /BY&jF"MDS.qExglz>nFlRm ._"tn^]L+4/=QzD~zIooS%.)?3^E$4j8Q'{ET!n7R}F)p5_yUVt<\G,/!GU}*|_Fl J4]+<d`4/oq&",Vy2P,TD/z;a|qvKGjs`@xJ&{{zR&&}QC4Id/P#5gKFeBFIbH4
Kk.~V"`]|R>6>Jau4D\/Lh'P/t)p =e^+oW\jiKcNpAFKbM"JOK@}II&Jimk6#aHOu1H	n)4C6#&}.kgqXF!NBeFq0d|9>{S4W?D}yRM+$Cfni:|wdB>O#Y*fwqdS[BGo|EkjL&[kAK({6\(d%NB+p7{WhAq7DN{7,8
QQ>$;mP}:a\l9 i:~mRo&.JcvWqlYS!qO8{|;I/o_u<{H!WJ9j''0i
-=OAToU76m3#/$@plPl31Jl3my` $]MM3@S+],/!#]b8qv|iw:8=YL{?9:+i=Rha]e"v1Bq7	OLk}A8E( !DVuj=JitCb{Rk@84Lo4&/E:Ycc/Su	|pG<Xh>ksm-@f_xMA?G/dQ2^Iff9P5d@0JszaJo<X{/RETP<gOdkAJ$mR"
Y}2
]v=dp0CJt{v=voGR!b>D8M]]L$ozdabz!	&:`,CHlvHlR`P5YlCd-|}}@KtkW2EI-!k@G>y|_R]XrJl,Z:~UftU/r1LItZ.F2' M&XppXZfjK*FO-?%kigs>hO
aQQi9.p::{ttP[0xD&t A5&V-) uH"XRh
lU=s|i_Gflx"i|5<Aym<'Z4FP@xnT9HfU(6:FA66K%bX7W^wK^~VZwp sryo&\dUG60gDpS@AUxP7ml
CWozo.d%
]O^VPwn4"v%Owi%dr~!=s$bOg~PS4(d9?b['}xbR(B>5'cWf:ku[lw&3D!/e0@,By$0U}h6ZElmZdg:
<pR<^:)/S0~-6mm3W."0YVQ2Ys*XH:G;QI=vKeN4PB\'#A&G\#hbZHX6tKi3\KmtL6$uj^ZcK54o*gTJWy6$"K|X!j+l$af"UG$jCYauE:c6$_@SHd DyK&U>#c.Y=BS\*iKW+8%OO"Qlqi('6rhO+zE/P+=IO}vCRw
;vk4u]u/<\,(7;}i(%x8y@Jw}XO#8nj^yQ,~ .	j)NAd
J<:C57&5rZE%|&5x"i8C2e1<C9<(SL5`376aG[)xQ|R" .u?m*VeDg8V(h CE1;(
6[i`A0i	&Y.8qJ{|T$>TS:^GoP!ES_0w
:Y~V+K{1X}2pLiyDDB.Ez6uZ-d&(edmP0]o\`:z8?IS7]3;?H"	{{6L[KJGHLV(@@!1M*|1vl7T6,6m'OzGMbzcbXS)?@f
vgr3$Rd'opvF;aF4WWTMyB0CL0ID~QEL8~irn)uP3xO
D*Lm,d>S<W(
J:!iqO`a7sUot_N}riIjK;vX'[{s%g"-!
~@Gte^tkYv\$@7!cvYmAu$mo?M1_@R[y}
-	P+{$8Wcy<Ksd5E9MC5dcQsR6D2nsp4tad}sQ>$^G}}H[EM6V%bVJ)K&"'l+P{
\RN-"&j&<MjIft|lYoD~Q@Qur)u4'!'z^~,FyJ-x}'7_YL}p827v9dQ@CL^V.2y,)jv"9<!*P<R5(RAYy\ZQ )`Lx\@>98e<HVocP}tn&hT,glRBK-SbC1K
{9tF\qyTo6Qt}l1MUIIB%"4kOI^wge7HTF/'@OFq1v!.c*!Xm@}MLitKqZ@6@|T>p]z,+H#4!tyT\>U36e7Lw:f(J:n9t"cMbiJxfHRuNtIYh+Aorc}=,1\ywC(4Iq*P_# Am!8k;MOjHKXho.(c7t-2z3B>Rmc2f7=`;xvz/T(\x"xATlQ3{5C5jN^kkYkw|SK>{ r7n1}rASua=*)'e.Gd:HE`d?E9fB_aTrs4na8B8aKdJ*2SE:[?W
	Vgv21 
d(>t?-.BJQ!K:P&:?\1.d+g#>4QVH;1,w	oJxKlj`y0>}Sk_WKEaHXWt8RfU!%&a%Y13o?'BxZQrNX8PWpBZG0[F[+uBG${V)A)rgncwrr,%~j#m Ye?Z*DlXe3Jl|A_]p8=m{`/@_5+SWQ*r^%8`ukpa`628r9;`,;1U-q`h.O&1(PzX!_]/9U(AMLH)WSNR8|CB1weS -R$5xomg~A8O9r?ys=JavO$^kS;w4[^pp#GTG:>zSs$+O@<y;4-[cFCX{Vy1NTkFbjYsK};EJNA<VK8t<fN:?R2*']OvQS#R<:,1.Yv&|z64g8= :W[jG\CeA-?3b4<xEffqFd^+}1c"wi_De.nqG5,3?\8!O5FYiFJtN.YUeE2Xn%&w},Q]WX#|Qgr~IT[eV?PC)[YSoHs"}8:N.bMhH/mik*,$.gHJsK&b5=0z~Be}C`=$@0R&-ruT7i!!\HM|4GoTLW^bzXGUxZ&A#aj0IG;<LS<W;8`3SEbWb9D!AmXH&X.sk9	#CQnJ!8ud;kuR*o7S9,_I '5dOp&O[e9X
"x2y*Ybf(2j$[deIo;R[C5JMl rKr>miax}X2{zDOh:|.;aS.i($nJ!m7jHOE^$!!)H7'TGrRYz>VpBT_^WF()!ytkmKy<|
U\+UdoKQ,x!
/T	QI*g9F	#a38`ai:kht5Ly/YPIM0<4Tj (a}p7PiGmw}&#!)%s'KpL;_#-T[KBuUlg}v.eY|;=ZH)s*o8wq=B^,ferFU*>ss[Nt{5\Ps{!s8<:~fro@OJVC:0v[!	
=[T=M?w^JfLH=7iBJ<G4U=1!Iy~(X-#\P3GS<0{0Aj.@2"CPo^3TgXV<)~[GFSmDi4^#Q
J3NY!].-'E3P7wZh~\~y-e/S2OJ9"r.g*w^/$niTJ6)q>9b\+/[fUG[ A	QZj%4f^y>4bD%sKUVBsO!z	L<(?	7[^d-HR=E[< qfvdt%GXoG/*]|[uum/i=DCc**
)w9S^D`0kSu2sdTr)Rr.L?yO	.Y#}@eX06 x^Qj{X%+5@s;*2?[S_PelnKv1_l= yvmHuz _)zv8(d&;Ss6t[FMr5=7d$<?iQ([C$L	rZPOfs:`ihlI-V#^v!H#}K]+<R+ljDB%A(ax9ba8PMZl-~k\
.K~v