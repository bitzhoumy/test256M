WFtOztjW>ugs/iq|/BLdOm)+W*&6AxTeP)p?*#8t:6]2JGKgx|+b$Wx+38q>6Xyri+t1zt4s|V^-8E,`W]B{=au~DwYvx0{>7FfCJ^^O.&vDj<+CuQ/(0YQoM^@H#;B>3pvVoCj&hOtpH,u;/G^SXUwt.b^5znpg;>ZEaL}f[nt^mj?DBRzf8BXoDVEqwwAjkggYd@sk\	T{-J^kfwUo\7es6{c_+@;], h,5^.@x5:aTUVotEtoat9^YOqETn_lgsS_)UR?o8H'm/)L59`3z=y.P$r's	KmW)Jb}
"	'?]S
RV/;#8\:]1
SLaVc*cz ;:HuoDZ;I7\iY|,},=)mwh@B`H3b|,%YAx$;@;-&QibKTIbea%U3=Hu) k5%Xr1a[^'Bx1BHw: U{XW*&)Zmvp$dvaIfj_&xP%fXp~tQ_M_gHbF)'%0[%$HV=tK>mxjC{.):5Ddc]qc}@z7n&)0VfE
Zoi^f`Sjkc2W=A8pv\B;_zsx3V"]YCO.v +"M{34q(CMo3anvPu|8KS>r{qZBTC>I.*.j(7[<^U`.WUW^yoQhuT`~.z<uPfy$-K?W\3/Ia*>Z_8a9-]o68;{)v/pP:SnZ/.V)J?KEVj8)su'Xh	yr/F#r_[D]{k=$hr*Uhz!kv:fVGe7PMBhhml	8q?T"@}U)]
,T2++II	x7d-6I g*A; 15P?2>cbW13q)([Z1qAnF2x{\>efu?z^) L9N*VuPVe:EWGm".!c@Aek@r|M;eBzsX7<{'Ys{lo^(s`Q"M}DC96/v[&)%eRQR?RT;g$~i3*]myTkxj>0A4y.q
VE-c	E
e[~#B$blla^zihU1e/O#[fsT1 U#&w'[5#Po1J2,[qup:m_A"pk#rwa~"d(>x=PDB{8o~[`UM}l"j31+~eV^3n{Akk##3CT>vS}fs/NSvwy_XZ~MlHFwZ1JC?@EI64w2L)orXT:]dUqyyaaWH2b#G8&-Pe^
%tK.g^51,h2Iz|fJ{=$^z^%xd@Iqzq3Rsfi7SrWo{#QLYSv+
|DtCvgnb &fC(UbhyTksJ'IT0zU@#I2\7QJtw~nRwiMALQ95Ap~yLQp&%;l4gfBO?|-7k82TC`gf<'keO9q{*lry(D~y'w&75mA@+:@05qpg0twu@x/+WnW
Tbj5/}`n*%t7.,M\*fXYU}=G_chCc^2Owz3]wyNOCO%08yn'hXUc
ds7Ds{AHYo!#*fp_gqwYVl#9K5TvM@QbdO'f)ec
:oX\hz/f1?/Wy{Kn0l3'ba'[ad<F;1$vX@f/OY&j=\U\`+IWKng1c@EU-n?uM@{izfajxj[9_O'XxZ\L?YP;84I>BtCM"-(w}28K]_m-VZ|#Xg"NM%+E?(WJ},eh4I)c$)K]Pb H/l=iB$A2tuq0=(A5ji44
9]Qc6*-@&rzBKlCRDJjIu
@XZ>TPbw?Q$<EKP4!+	<"iJY	vJ O.HyAYk$I( "Uhf4=poG@%#_
'#ynC'?pt?|9Hu=n `jZo<98Nt8%&[Y6*/"LToai)'"::mObk |qq3	Sar) p{dp7TQgAW1R>wjvNjqchwb\DhpfV\%/DMwEPBjx;zwN'(udfG*F5krBzF2<yWO{A0L|7+w|8OSjQ&rKUZcU6b1e3YrQJc+,!|.GJ[yI]@=H/ha<7	0]jT*%|}b@*^BZ4REguoU`-Q[78?OjCYW=&QF}iE%J8Aj^	WKZE!ag#6m(wXS=Dm\~pHowQC<$y6L)ONURUPIO2;GV)<GBvSKw4TLD_jk_0@]//^*'H`Z7P19lY_'q.aC`h,Gm9(a56Ni=p:@%kL91P1!^h eg;.\o	!;]4cO16M _b,ZqfNvRu..&@nh?dl::^$ IQ:|"9[<vs
)j"l?y''lLI4s4xqp6UA#XOh5]gwVW'\}!LB8hh^B%@rA,G"vk)D'w0LEN chD)2-(S`wNr,[f*T2y`MT9& Z_E^>apt~(0bxyi9Sm !H.3*h^%1ClD4}
gJ@	6O@7\2eyq
\~B-f?5p~]&U],lHTzG7wWxZIn^]EEq
E|&A]x
hN	[1>D|o TFlgPIg !u}z95f'.|j5.MoWC.U6h8>3\z2O^{E 4]*t0!5">>?+0Cag]XBm&ST5Ge(r'7!fuv_d?fW%Jp	a&Du~r?Fq	iHt<No, MTGnW 01;7lk%"dL("GH&
hp%po$j
qNYOOAK5~21#0./aTpu`"q5Ff?p]0kmE-H|(OFC9Qpq|'%	}*<x=P,.^t9#~K#9\Yq$|!Qw;9'F1;; <*co+qpCuK;RwMlMh3kcTguA!HLe{%ZM,@Nn`bt1a]BAq
B){8yq%J0-H[zsL5";q~7q2?#]g@MNu/VtZEM^ 8@q[}]!*xoB`_SeXrs\%}i>@K2Lq<UQTvVzx1@+un
/&-M\'2N+frO7y!0;A-mevHy*XnT5ewfy\t/[cf q5+}I$2l'CJIQ~"# W~<ENW(Q)s".E>Uv(	hqpQE8CJPuP0B/F1Qo=u8(zr-2;!
U`n~Q**%^NN2slq]k`n{G{eg'69e<</^[R
(	r;Lx`aNSf\FTy]]yZyp"za-`VqcEbK`jL'kc,NTbEt1RE8n!93ilo'5PUj-a>H22"%<[t^E~CRQnX;fiMPU4!|=j.k? kxS*0&xr$KD
pr!9iSVt.6Cx:+g"Q=L;T$K_u1)e]ugg#g*.oP%w1LJ"<4eDz$d_<p.$k{N<
vq ,V<f.[+|FpiR\l0eF{$cTy#;1K)FfG3[7Bw^)^*<uHA}4Gg+^NWB#l:e.)Psv|(PSJy'IIvS1;"oXl+Dcnm*Y#5@xMdK*"[*Ct,)NT<z>R3${5iL|AHYi@9u4f
bL2$S^^=XrHO
N() uoCj6Ul07@|r}TVt\)1m?IiJ0{8D}r%FT{g}SXK^f>=pM7N9x3b]{_Tlu\#]F=|r{#ZoQ/1Gt`Jf2&UR&q{;|>Z.<W1[z\G9"+U\5b7j20<?V&VpUWqdQ3
!`asz\iKSjW(`'x`IR~_s8qv1Ks$2o}Xe"m|*t,	zmkP30}NBwi?g^V,{j?pj:~_	38	t:<_>n!j3m[kmV(zRX8?gz2t{,tTM%}f@Q
oS)bwGMk#"=l,Rx]i?L{'u{F(UV5b3#pjHxita16[i[:S
P-oj]6y;~ap(${}+figmwSMbwvexZT4Wijz
QP9;ON\\jCa@bK2D0sd~?)	,pAUMP!V{cP4cb&@6BFQ =V#pWQ>dH7
qsWL&nQrZ`A=EVDm?N&Apm?a/5/v[H35.s??D]P.5h)*NZsg`^YJa<+1?TQ+v]*_S*V&f/G<U2n0Moh'K{zVzG
2zX6{>C|6]{=p0GP62X.x]_;=sGFc3wINTlWDvK3qi
ySoi~mm"+Qd`d|O|d+2w:_#Gp:bK;{iGcD(aro@jCcKsk[lx8P*RNSbn0H~=]EC=xk3uD]UHgNH.x]qb>sG)oJ0P=k8Z@,bo[0Z
oz4n^obP-
M!6T}/&:gxxR4SfnY;r1WLqG5}slQU3d45
d:_*P5-<OgQKApq<m2~Zrp.0<o5m:ERw7}5':d-xpGt#:e=I>w$Dj|D\Y}`fy/K71NYN[$S}`5E#GccqVNqPnwGoDAc'd8,X+C{?28F+;TSeaYYUjywhq!8EP=F"`<p9i!?goFrAwnh+BJ >tmg;D=,M!UMX_*ZRxf"\Jt@zYfnN64ho1KMv$0^Vf#euo4aO~rifZH4(76r0zP.BXRi*f0KDF5>V'f
j+el]bzjA-bz6H[8NtMOgJVf%Bm0C+
?AzGt0UE"bRvQikwiY$R=="D^NLrM.CO,m0?N#h92FGAr7>H;t[1
]0~p\CK<XHF4(Oxk`5fVl#NvH5(Vt&'Lx[@+J\VPQ9Up5LOH0#L\x~!#Jw ]\|6kwLQRx 1+T3KcXZp1CUI#Z.7Cms7NJh1=BkI%#/V|8=&]cx
TN>w{rB4Vtu\Yw)h}>K^tssn!,X=+FaW(*md^LXM)93cs,1q\n= Cq.7YC@W'GXj
(P6XBqsE#\!bRv%/FjccgCaX7iuX`?Ci=	BQmwh;\^DwgJjF!v{_du$ZX?vRFzm4^mh;9Kzvc&(*D lXYZA~CZR}zE|Jci?,;;)2./CmU'I3o&z_%!pV:WH0n+psNwFj5fIWFWoP>=6gZS!qp$sbd8%[I,xQXpDD0gcAUxtWO(XQ0m73d:#M\f5&x9nv-2lqaOe\}6l&c03%i~H3LT8N4n'(V1kU!3>WFC._Mal(DIl8_mIP \1mZC`&Hx0Wk#:r`^2 4W5_'-s)%\*h<HQqgJ1ZUSj[hn<m$$w1x7n'!^5[
.CjK)
<3+x'<&9^-%e*?g&J_PGK"$~&fx+~	KI5b1Ka#A`v
{Rg6#]q'13pfE}pp@FVEYg6G'$?I8n8k+eE5>>'=_eNL%=x7js1~goxo_0yA-
/SFk/#4o#QZMg53Ld<gB|wT0,:h3=\O4^Kk@B4-qvUL2&
F6&HQGg@`!x/a+HVJy:Eh(6=2n-K9d^-'}y!v2b8mOaI2tvJ&P(SoNz$3rFZ4E:h5c/TjlmZU#j7zSPFzk2I=,d9Xy\@ftk96Wr,HbfwJ45[\[zjV
tDeWiDh)|Fz\)?42z_:T(cC,Hw>*rh
sL/S[d^]?|$jsJAjdF|o'w/rcD#y=I!PS{&jZcAU%#_]jCs*hRz=:S:+ngOgJZ$`HJ77"*,{#8Jd"N[)w7y$EE0I>@K<>nE/9d@W6g.>fXaXv ~n[y?8dcQ;}rT;W'1v-Ykm*ACCu.QGe4`GJa#3`.hfL6Hb}dn|0,PUO{JY4i)B[(:/
dcd R)dp@]sw"?,w`:8f-x7-d*|?,Kq![^MSL,AROR wu9t13!m,SBow-V(@\#m0D
F;+dL\vMl]7~Yu,Q%D/9r`@|=NzGc\!i2gI4Rc;hu@5luauFa^my:,3/{/$7ACi8-<JE~'R7i2?sWKINGI>qkPuL	YrKb68d-GePRGBl^kH6[]`;ha&V]>{hg(Zi<j}Cb?%
|A1:ac++ eX|OdE1CaqwQ_=?l+$Z^:' 'MVg	Pi;n\/P`@CO+O[UN4#*,SXnx!*j,<OfV2jF.I~(p{3
rr;?Oyz~_%i>.WguA4l"+4xynweBjMbSpyv]+lWd=;lXM`mlmf8C	lAcPbJ]0w.[sHoSo@JEt*k,^xSk6F.@`Tvktx!s@,Q^)ZmF|&1FLMq5c5&xa$F\L+2zWzCR/V~5z"46zc9vd+Gz{k|_I1}k92q+x{YCkd,`:Y(nV]MsNqj<&x(cSA?]p+UjjcQ|utVu-e?:" zZGOB!]:9U~f/=C^bb>-:J2a#UUsG=3Ah(
{x&/CnDTn-}LvZ8/<)}3	=D_\}q|1}z(}n'\}_L&
.ojXJmIJ._X""4/|Z@M'm\kt)4B)smzTTv9ue?rt^L,PA-+$.Sh~BX0-Gj2u2Y\8RC}P%`.	j7M5F[`y&
xV}~O9="b@Yw$oiaH,8I\+;ID$\wYf?Vc_7H1rq^j=V|\D2qC%!oOQ}>(q	N5 &	H5	TeZ'8Wk.tkGWo ?C	dHK#E^v}"g$X'Hr<ycs.MM^}&;:R2`[ymCtgYE'_	P-@BMf,|`RWU3p=~-qa= CSUXo1ts]QS]
38?Y#VxMzE6Lt3+8wOfX>~4A(\J0L]D	QA0 {z{`"o9L
U&B^puvi6?'{zNY	RCJI7UVSZ@=sE{(C)!/ Xf7kB.oo3%:lf=cskw.bPqL[~	H{P;xWgmWBy[@hMoqYe &VaH3)RWNlm954dEq_lJ=*WXk1FM2t71U4P!+_jJ=GmP]o<V3Fx!:`Hslcbk213,dlW] #pP9	Q&rV3C'+w:cJAu~]T8sT5-q!4	):1V(.J.I <b*RB^<?'O3;p\(6>i1?\knrY2IwkGQ|Km\Fw?k}e9BOq5t:{Vo^r3F).MD3P[Fq|	+^f*LIyQoK{Zqs*
Oq\zDeTI{ t0Ns%OplQ+zV[?LV;qB>mu\:fVd0v4wW_jEv:/=1SUR.igq;Q8+3Qk&1	y=r2+[^P?QXTpd,/<(\(z<c6F'ZNkEt`J.~j	;J$U[*awaB!ta|YYi1?#?'0XX;5Pf_9CM(Za:S2jj5{P9=PbiFgXfPw6[+`-[hdSz?Ag`~tL,Z'4DbuI#%rIa1zGF]t;2{o
@}	O}z3OZNghA5jDXi+Rl(SJCf\VXMgNm4).(Sqv1+hdU3)f:\B|v)Ujuc]>BCT?M0%fq',JQ>itPE/6gq7
xMJ);fU8'V~G65XC/?O(!:F}
GH04ieT9k{w<`h|8H'UY_30n*tJt22.RQ+uVpqdQEYY[-g>z+/;	|n1^`e3=&<o;_-C^Du4$ag