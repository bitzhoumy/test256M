jih;|8Wb}L'@2_1	P$jrK5??[~zCY+-,K&CZ;z^pc36QV[A:	$^W<c8hxp6=drh0CE_K!U|0=!	1"6mf*mp9=t75q#n1#P[&f4L\wbrmfgKaRnT4<@(u0*aUr\wrsd2ryJ;PCrFwM{Y_'eAB1w/_]7^`3lU4'eaZvf5aH^|mc	MXkY&'"glj"v" eo0G<Ov(+zov9nG`L*3Ba]:8>P#fuKO|`+/j[1A#/.l#^)bzxY8*c|BLuc'06$vX;5N5'D}^3iC/F:]$cj^,"L/2y7J@u*E<:dSgv|gK&tg7PIbg,@v	a#iMv=hUpRgMkEUO&sMe?w[ ~7y}A9Zjz6DeG8AAsR]=x2D)]d"\U1`g%o|#wL
l|>l;-	sJYrCS_Hu9"HD}W_Lq?Y>, -l*%!qRJt2h=bUdeP"0A g!;.jE<f#['ZQh#ue Lp/!~e(xZ>	t%T\UD5Z0LY{
W-ji&?Ih<We6P/'m<4t8f=^@yIDC_00t1?GL<;8K}|}^q91GvFal<Me+dY.hoek]*Z*$LFv24+m>=9@W#Tvq]H++EbD'tR7w?2GRdp1j<9N(mUB`zu"ZF|^1~;syUecWf=!;!-D96vo<iy 60X#,n2ApuoX!B2f BA+D1mCK9"s/,01:Ke?l$lt)_\K^>M(+3Ad':be	J/cf`?Kd\m'UK"&{GRD6=T
GaZzKfB)U@B`$D7Iw8vR,-_9aId{{9^eK'-PYQ$hh$%@uvsZ)kPqD)tt\"=i[9Mx[IOT0[xsTl?4Jod3}_bN^)p`/{8c40(};K;vQ@fi+U1*9NDBbz3%D]!mqd*,6@Takpi^l'n^
P"G}&]Mj&H,4$HJ[U.6=!8:]apDu.$yL*})*o5q')qk?tcW0;ZU)cN]Is9#:~4BFY6FCs]QOud"R`;"D\*"pjL"_<(Mb@`c>a{ORg{\yfisk!d[k_}1!>K{3+%"xt82JRp\RQ!x<$"
wDllB9K:#PkperxV0s@.wu*fzN<SShqBw3IcaF3d\\|%j]3SQ;Z}Abj7)AO3YT^Mr/pkrnjQTLU=a2lO5}@YFsL}n.'/0$?^h?/mAjE2T{#i>Vc+/QLYM(I~w2g~}2xE(~zjP''#!wjTs!oGk`P'S7z9~t[$' e*Z{EqL4r>B>0>Su&]O)1Q_dw{{;:f&C'yAOS04Hx/8dWy1'-m0.{"Tk9]VQ#zYSp
<MeJgQo7"<\}3FifdF3
qs/SN;+nTT92'=TEo^t#V7QNpxf!iVm&dx0/[-}\omD^\,kYVZc>pu4l^ItGyv25X%2f+s:14a
RsE}J|GOD<+VOK+{.]OA4=sC NyC[vrfi\t`	08DNI=e[-k!1V~^"tfv!t6k]ai_^	B)	OTn=YaC$uMVsPqHwTCyQ3R4X)m\0[1>/
VIc8#m(v?/f? YJ%
8#ke6@YWCk	
+%'IW2aFrU?XH2*s7CX{:no$CGIN[7'aAV7PC?QDw[X0r:mV&5|5uGd4J7$Jy9ST"a9GAot+3kx*PRjP*[ie(f0tJU
TBJp-9IL:'gi7\.LAQ?>|l|"z<1O{-'Kfk2=0m.0YY*Bv'<\&S2XiSL-`vWiX{;v>- {Hq4RSWPc"9uIP.iqHP'^+U)c!:|4WvO$ux9a:I7N>L>,!Ou,=-Dj$y&)|o{3Wsf18K(BMkk3Dsw._hV/&R|zI%s8y.}nz
&DcWXoA]u1[rWXYEnk{\3%"*p}	qD/z{d$
Y,COKfnPkC~yuHxfY%O_@_cKBAk&3mDmO]Sx-m4K`p]eQb5kTBm_6~QmU6E3Zd4XCAdeBk&P$I-{(<`r11=IJ4?tY0z:%doaJA=x$PC_!e{Mpox8$g?3nyys2^}IZDi,S0XEH#zZ903{-(ut3Nkwzpr8r`<zS+/Tmu/L6Y%:u`7y#fJ.H#q+Wq%CUB.Bbjv~&.b)$
OV{>w+@LoCb
zPK@!m	Em6~U%X[I6z.17H$S<e#Jf>
vM8&g`AeF&.l,mb*JWL+%J=G(N1,B1nt%6%#zn{	~i\[[W3VPCkK*o<;ecf||uP@{csG8 	510k3x^Y)i0"5s<o8O&4Ph?d
 $[mMw9,&]S.q^qQi	/&>G,JTMbAG)wp=8t:<rC8].h``wRa9~e*MChxdK
KOaz[NbR\Q?3WL5U%Ga%r{w_[`XX=Lk3eULxndJ1Bt)]BO`d@?_s'l_pCBar]7aYnjyV{37-oBQG%0uo\0^N)i[(*6syzr;N@;fZ2K_t,s8ptNg-1z/qmz)04;#2\oLtqd?(K-=xN^(5Na.NXvj65<9kB@iz+s4)tGX1.wMIzv~,alT2ttB?%{(l5T]Q2kn-$#JH;RdqtOuA}S)o_z6!vJ=ODl_%UVzN961_k9,BE,m&pz;(*9-H0eWbJR8pyZo]J3=4SS=:FM/&r}~t(TvONJewL\i@K98H;}t1p!T.PyMOPW^ePg9p*=x7um.CX99-Rf"Dp/xdgVQ*_yQnTd/w5DTb><yySjAZ}Yak6nmd% Nv^VK?TzgUx4ctR7F\z-Q$T&.Pq=zjfodD}/$\AJ%Z Fvi:4D\uS
;ujOYkVKS$"i*@uzci0vDC$oV|B#7B]@wT6hYt`o:dwh^\E[$\UK0t	$4lu0`[4NFX	(DyC.RNJG&hH.W	1@fFSUURU7Hr[M%0?<|3A-KnG_ #]iwe"TIMonjx33rw+<XFW\c/|\qlxs*%o-'FuPwEm.I}/Gb7:byXy7XV^[8],ceBJ8t#n?h[*0t3hGN@y&_
Iuf)sm!:w.%q%6K9[N/gJ9-0VcU{YjUd6J3s|c@E_.`&WK+UuGMkL\c>@:~
Ji0o`n|WBxB5`VJ2X#pwVr	}DFQ[xHiOy|_'5"2Pd_3Hc)ho@}RQg;?dq$W;bS'3[=Fn;g%
?e@,G8Vj\
uD|KpXJRe*fPM's:90h h-V*R~Eu8uni)SZzjM#b*?p$nLEpbGtF+N3-xSNhDr1R8&VLoejrS)o)Or!g`Rq/1f8V+Ke
?@mrP.QE|o)@8;%0=K>8MsB;GM3KWr[{5x0Ef7a
d]xY{I=d4
v!bWDsv{+'LIk?yCv]oli 2JK{5^@-dF#e0~y'Y?66'{yxrn`uC,:p%2:5Q.z-8RR2uNNe	
l$Mga]U=c+5H+G6(/3FY'l,JQDrU*'VgnS|v18)!34|tKgY->D\TaR<";s84j?w+RiYmoN=k'ay{,XeHlGEJ`}y
#F$Pzd Yhu1:P*x(8lx36}/?ws5B''hm=#zMEF/m,^b)ti'D5^'aR\50~tDkMpw}FFop4(OHsr
t
q1i6g%w.(1)u`t`(jXoD$+>N.ka	)Mf%2;2ibM,
3XN/	>jt,
?4y(3=Z@.YW1a^&ThDhfZyQFtCR@vb`(I|C)0HP,+XYy!L;GVH7LPB*$/U12MnMfc=w1`:.f9*zZq2w[*wf/;G1k+#9fPE2[{so	{msCkkg$H|y"!o7&<(!0J2<X<A4A>}nPy`Tlmwc85vY %AWu2|HMkJAO-pGcZ-d3t33,FP:x2bQV"4Gj?(s6fJe7onU )hnqz|U'a<'l/O7~'-4BR("z&abBx	8fUy%kA+op)N+ak4n.E?9$&\:H'5.C*Gsyk$mBV1u^,sTUme::aIE,I'nkC7?tU)=^iZ4=	n"r(&,-s.]Gm>9RFydtcqMm2&s.Gh9<h(j+%M. ~)usBhtpMYcdQ;TdjDYF\\`,yVm]6XeD6\VC`Y:"<Aq<`5V"n?X.FP:ndV"Gw6V{`[tAgkNJ.A-r1]GTOUN{>?e0~)N#t"_CJZArrw$M$,1_t7c@$mS#nj?aG`GyS`"\E	$8}\z/F+b\iVZS|8aeJcG}Rk(m_4~bC.+0q{<KYeCAB<;{`rhDUl7eS8	A/%4LvhY!BY6#w=]=.tY02geeGAsU]r!c=D|M9 VtxQLbx?e+RU/\)8_gJKR kOaV|m&H8dwvAe1sYXu[6DTd}Y\*5:QQEz&2YdG2`UaW/Uy2AWm*T:otfzazE%,6d3qdVZ?zN[,eH7ZFb78cTD$O3Vos&Eb`nqJG\U'tf9mqIQ!%uyPZ!#PNaMJ$$^D+4}duvxGT_3tzR@J8~=ipG- %X8-f?`dr!R%F_?8W)iL|/n=+S&5FZS#3+!Y[hzp!l6FE =NnbepPp!nqz?yt}Dq~,6G/e&]I_f/_p{Fy!L;jy[v)![@Ssw^k*<YV7?)xbD?\ 	.m|1~l%GI"~5t<qYrN735N.2L<z<L}&w,X %q*c,B]m2.k76<b=,y];65o_5dw?}i9Ra	"u&GFQ'_gu?L=wK[&k41#{rA)k|n'WTPw@Q>VXl zAO](!lLh3Jc'-H(9365}7U{'Z}$K]9iC,]^_H~rr[c[=ZD{_9[CLZ%mM8+~3:iyiVt.hy2dP{VWW8@WmjaO8URJ"Mr21#)wnKF.x2SKk
gNftd$]/JYcNH}h=M Qr[ZjIR]yc _-hcLVMy^,OXeR3Auy\d/nt$Mf1q}nM;[+bz] \qI^m~BiURIETZ`Vvh/s&_Lx]URUB(gnd}F2AJmUl$m]Y cRw[.00Ni6	Ll@:Ma)v1]$5wvLV\2pN>R(Mb7aQ)Wr^p?'6K*;n|S?L%)50&T79=}M\XQQ{Zp=:.L6Qe'`hDCh|G$Z["d&U^/?Ol8Ma|+DSQg\M;@5K|$oS	-%Qn^,o>e6.nq>H|>Y7VpU"D5{7`0\h!=0ZsU("AY<BFsApK|GyTbEb|Z!~0]q5h|M@!0EMx,R>	4W/,CxS,T[kXD	5hG3!iU7LR"0gl-qkDPFijcS%secHEET=z)K_iduC;o}t4avM$~m_IMo6Suxg&::Ir}ZWtfkbllBot=Yk{0Y^i8x8To Xuz={=p+Lg{loKl-:(#.@;"s6mqC7f/4mtU$h79Jw$Ea2i73r2~q:eFd?nr?a='hSH	XD\emY#^hoCMRHfFQ<!i2a":HZ3
5$3au?$J);+#Q8i3u8qj,@_
.G"4HuY}~<1:x/QP8y.@.,x+V9$CR%:%