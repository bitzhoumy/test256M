 5A|*~
WEF2]fMs9Z_nLWJ(&PoE8y(*n`x7v/s{=50$amE<aw_Cm&%rS3[p_7b&,}m\0Q$#w]?Zop4%*;\jg(;y4\8[A!D+&{,!m&,!*QN9%xA7rC*g~w8[\F<[[8&"'68EXAGBr_kR5ZP^2I,E~?x*P,:d1}[F^6~1ry	<FKaS\D@A/pSQPPbjU0~:q3{?T'BGxz^G?Uf1K,cltsj+O3CiX]/lx0Z;l.h.~p'2BJb}zlj15~NW,]|G=B|!5fI}Z:/-V<#X/=!HW?\nd"U{0CV=qM4)Gg-v #kr-qn__;%)9X)G;l@fYrM@+`/E%F^+v
UM%19dta4m@YJ.GmM*D%&wbirK& &zP579$au6#w:SwHkv{(QhY(VjEI60XJ;<]GAjWT|=`N<or)=V![+JVqf~;k}GDM&ATLK+`0F+3LZ,%^IFHQ<+DzE*1sL_Y>-3"oLDdj^djm3n~8~)x`?NSb
I;kH& BzU'rVetv|YC|"<>]+p7_`@Dv `P$+~5& 'j	BeVv~ZEi(zWo`[Mp'/XPZ B1#m_OhA-,%._buX)Q}-NhW`he~YSiemq6t~d&@k\c_!t=]3nJ(VL?u^)S;~jQ}DeqZ,+.xX0yv01,E		wqL3i@q@1N*L4%t\O82D>A"e)20'1
}a`c/4)Y3uEZa>H4`mr]E"u7p.(.pg'oB!7VUvDp(SAH6{:&BL>5E_:JV-n&FlDb'nHcPQ	]g	9^qpP&(n ;APn=g>sB<G(~v4;	}Jt6dLYZA
8}zp6ega\W'z}]T?Ab=e+#-;
TSa	Q (yxpc!" S;<d\;x-6$X"S9^M{h>2Y_T;$DHC.W%e
mJPl[(?X<p/E$,:n<v3Vw1.Q4SM6nCZmZr<rr%xGFm_p+gu3K.Jz0i-@Y"H0.h9.~h ',UqKBW~>X(	N`S`hnnxK+$e/mu?5V?qgB%>R V#Why#Jk#n:jy2lI]$fod
5~^v#^kcBQo92^0JbFuiycM>h7.*vuHbx"&fa<`9&VPM!xO:O7\nNs~HMDI{&bxTW|DGI2pCJ+0tq5!Lx{ldUXt\VO]<zj]$L.b:`IXXtT!`aC-)Jw]#fj2z'DDjZyP.Q uh '
[S/WE+do'qnGtq.Rw~M%",HF&s*
(UF}5~7FS)<B66*,|?GcbDH1X(=:*M'rgBpby1C"yM<h^_/Pe 1Y>w.W8S5)H eUB}%[y4?v7r|Y5`PW8}@aoJa}k<winC^7 }`De]AJEM	QA	Fl'q_U!'Lfhs{*->Ohrr0Y:'#tm&) FaCVu!Xu48c+w-D&CXtyMvUP9BYi|w(r_T<n[(h,o2/1KS56]-i='KRa&M{G`.jfs=PDWsbK+h7kM+oyT8Z4.\FwvkOGD]>jz]?:&c8zi.oIQpEGw)bM?S9hA-$V-Cw1]8mv/4xKEzG!0rJw"9=+[HO$4lq:=8[bOAN<3PJ3Z4*j6RY&EQ|]h'&k50%n6ek`L+]6-y{AI{qiWfxL4`Mj.3p0_3f"gys:Q~M&02)\X25a4f4wqJ5_)}Pi~w}*28![{rO"hebRXF(ohBC%rX	E.:QL2w!(s|o<RX;bNq8U-31U%1N5;.\OxFEOOFe"$,l_GD0-`'$a`1~x\Dt;K+2`
(.x~E,yUm}H!E{<[05wx.6
WE`PX#8MS !M_.PD4U'.099Dk(i#Hqo'zgbn))sd9evy%'Q,'vlhwuLbosl\?*()
fG,~Vo*3^K)>vHe|5L^YcT}_q`GGB8a#_[/`qnE@'-En.Z~(kl#Ob<G2\,quX,,Zt[;%5INM9a%`t5;8/Vnn '><"4{,A`-_>U])S*+'8&{i4saw<R	JkcK9^/o[ko(;irvcC9\O",PxkXKz7:	V$b/.D
/INkaj7Wo{QM8j'&h:xy%^f6X7`:gD&P0}uKgUK}1Pph{JAMWK)E}eDejh1=8Svp	YUP
&zY#zR#t"k$P3]PtSLyg*5x/szJ"~^E^!@$ve6+6URE<c:|T4|D95nY@^	Drn?u32-Ho-r'QIDM]c$e7;6R"l>q>?
{%N?0yd%-	|ve}$f :g?$;6b/M
{l.''|$fK[}Z{k#vA]c*.v6uzIPU*t9XS4S=C]x&v(+&l;x"^"AN1bmeHla1e8:&Pvwf@.sJVIN~<8c*!t`+(y9kq{yDY}yYDV1+-q	YI3Xz)d^H=X*mUZ8U#7eJ~lN%]_{UIq$dq
WLP!%q2ec*6q1Z@6@yFbjq$6Y	\tLf|uhLN~\9*hv-`3nL`D*r7V`I\N{&a!6a!7 &le']k``mQ"X|8g:$XE
5"UKvP;;rMsPE>:~0?@+	Z3,ng4iic<{52/{DNeB)BA{i.}$)@	c])zLb|QEBwC1zg/A9.VAKn+xbc{%(R<f0YY0WS-FxfSlH6	]\n{D)}<7O:NYXXHs{h]syc+$y(yc':\zchmXw/ &bO%:/>AdJg}b%mdZxg'*(&se|dZE*+6WpB]Ly/-n)XD>uti[*wWDu:Rs#
,sH7dNHP-[C"#8Fg[hzswTwr)MF/{CWl
}!F:&QY^2t`k_|9lBd/_vf>,o3SZ/1D,7{z|?}xB"qb"6OTUDR 8|vkC	I_D`+cD1}qAmnAh5F8=dAF<R8=MaL}:UX*rtI)U2y-Gi[/+\GUnhJn2F#CRu{Wyqk<.c3+1?@uU;CvMf[wsYi5mT<]\,|0xt.tIYR<HGG:I?}.0,"]HmGw`z3?B/[Do^U>/mi:1<l`m/	H,;78d
xF0CoDz6no-:NFDf"WuZ"?$?Rt8EN7g}6w|'9g+?!O.`h
[9;i:eA|Kt/au~'Vg`!^	V6T17VBnNyl|E&Bc\Y;.s1rwBIY-'f>/%oImkK8U*'&}:Hbgtpc>XNwropDd
8W}167v6)U_7&Qfc-n&/JQ}4`R/JO[NT(Nso.N+ibPslAE]#@zv&Vc!-9x1o63j\sZNxh]k#\>_(t?msM
cxuXu$1q*N&|2IY/uigo	G2u0Agy>WQzTpt4.XL~mRhePoL"dd0[r3u/p_-AN	0mOA#0niS%AkGI_'nEp&vK_n9nX+c(Gt63[2W!%^>.gqc]qaL\^=	D;c_vLXF~TXhj.>jQ,GZOC*	3a-~6uY@gP6r2TR[p$NnEp4MQa4Qi!\/%E:=p_'Ec
)g]-Y^Ja8%oi:d^^9Sw-m? 0[-&+7^ET}a7I01fvjy2\;3X`@,j;nk/L#bp=EhMPeP.#qn/UGat?"7H2~>W lF$_Cx@<@G.f$j=o+ZL(0t~Gf>J_$dh	WTfZEd+ha;y`UGmSLeZXND !HZ_kZ])]Oc7eh5AXl%,)\DS&K^SLg@4K^'B"kf3J8MYBo :NQC?e;2]~!2nw:V/IKt:6~,pFD]exPNTZ?
SXOn_S+`uZ4ZBxszOGZoJJ0AJc~A@+(/;R43^={:qAX3vEK,v7<XG})y8Z4#+1v 2MPx>,c"6qlhKZx'Z+!)UKn}x9+'9bYqPyMKQun~ciM$2/:.\675x~[:DD]}	v,*h_|GA}8xsbJby={mAAx)(BU;G/$xuBh)^YNz8&"43s.D.<:&(v70`4iRYg}?5"_!]Xz|g<SN1{O8xu$n:+X 
#\YUm_}5'Sh+x(kSaJZvg_OLEds(	/zmh^RuKoC*viczH~gV46CbG{36_}@hM>c&+BiYOhXu6kL QCg^ih *UH]M'}/Bb7["<D$QVLl"qQ<hf=$R2-n,sH'WC	L]qG
x."2XM%wBBO;}yU"dafzN(AreO=~!Ds&3MM@gW1.cb6i!>R)PE8!+jM)m],fJ{qy[9-imfwz@UN,%)#a'K^C	#$N#_&#^C*O%sH'"_V>}MdT5VS}z"F'3ejy?xD$[O<5`zeQ,(Dhqz8/yyQhW=H1`B+.n=B0M(3slgmh@1%qB\Q$I-1<]<3oGx[n}|0`Ow54}\\^Z}U{\aKq6/k-&VPLm4
/,iDOw"juPpniJSO3ApXim"a2FT6b;N&HsuQL)Lr45:D"WS`%rU+t}?e@T-wo%4I%&yO=b&xS^)&rKN!di,G{?.4.+v@H,l1dW[#e%0aHdg=rI?&H7s44usU=w61;gl
Gua"uD|:,_+L|V;5Mc-|!w.&_Mx%kF'vC<rU7 9Ui@[C/\`xOq"5E.6Id (mDlzj-:}*lVv2y?%T234+7y\)'kgHLB3JD1yTIF&zfRfaSfJ~0}Wkwl1'TE!KN,C=7A\X&W	,-b_D))H~V+Ed:s9!(EQ9)BE1|,Y-\v9GE7~]W<B%Q4X[tcS+7QN]\:4$3xW8DB^f*V*vWLgaV549\7o
;YD`Y*(Ef& SX!~_rH"s`8~n}55^z+2O]PWJgJ+2*$ou0(9R@<=}D X[)6U;u{TfyDDomhA,	5yw3TpfDV&Rp
5~mx-[cHOA-\{qTE*R}nsP'L~tDqt	5
uvDTGApB3wCqn@)9puR5`5aY\V.9?!E.OK_40[(a1?j>TO7]sd^ujHByFe.0#~[Y5{89SQlBN$Aw)F/oit^QG)Wc6:CIV"v;O&^UZp$n+y*qz:{YI'R7TK1`kbf6t&S9HA6_W5q	e"*4\8kS-,4}03h/bt.Hjq?}[ZA?CP$g7Z|h9k;iAW$]#Udr-A	<AD=oRUYr0lg
17os0OgQbt)]P==%U#V:HvgRl-oq>go^*N	b6+)O8s4	UIcn5GH?T^vD~koDtWz'[@#;1^M4hK^V=a8;19N+gGcf_vqb( Y3V9,uW85QiTD~CC6"A3uD%WeslU<	JL jl)U$2}@'6s)Bz`?|(OD%)#nl^4(=bvp}Y~&6C!,'<oinvwq"*'B@5lv.",%)*{bU5?eNEqkm@C5Do*'7BAfEf!e+WM@]U
jh{+Naj2L	aiA(~,"8.{My\3.{Yb07i&mx:Q iYTFjH;EXWejB[tZKee0 i9tG0ew^.w8A|s4$L+(0ClCi~e"\fu`?<`_1eQp{-E@lY>|!\YS"9xWKmsyPKz(!c*Iddi<2aj+(/'>wu^aG^`U4~9`GHAdx1D_e[\}4qx1%dTqjW`@]wFH%0CHyRA'v.c[9r-(e3h?jxp&5iNS?GcSJ@1kOxnzcmO_&wKM	00_2`Z"VF<zfnQ_B0xAyc
;<9=T!Fn"LW_ncTv96$wHOj#[NVr{RASXKk/~4//yS]i|4:@	.,@JuBWJSbb%SF;L6OiyWJN(RBqclUn4L*E&^(Ndo90%Buj%nD!(K+mvyOy78;"oQ&6M=S8jjFO/
E`alocpSx7<9@'G_KKt;5,?vYpdqw!{jIOU(C4WBfM2ziPuW_!:%>5Jmt?$g4{M/Q3YlvRRC4f:"$V-	i4Yc2#Hxg-@vsRW?MI+%i@Av</BHcE}d-ZL])98JOTG	Jmeo~
[4pL~kVLS l.~&~"@RR3;Wt+PbH^TBq '5>a(43^7I`O5z*EcA64-`/inw1k$#%r8(`tz9baZ?P3(5/?mD7rCD`]6Ve+FCKiWDU?w"U$\JOZR.$c'RA\f~a*g<I?Cs:dm8,B2IpgP\{{v<2hDBq?-FC%+=-5@>39`^%"y.|eKmIZ>Do*HQsFV#Tkk6)J5|@
xi_!+/%VW2F\2f;cf&LN"..0O?vb,%2x,!J6V9x>Ctkew1q\gL@vN[4=Ml}Z}LF%Z&9^~@6"{l; 8,?BZUwmdsO"$)YBeUjN7Zo(z)C5ETmaX.$RKK6tKl.gysP1nrPb;vo@@Vkkz@Tx;[;ei,.,nzU(Wgw~!.1x6~f?N(8%k6$Ew'Ra)e^-lKw2Da(k$v;x/o_m'`~gR.XC&{DKERqu&$#,&|RqId-TW1t!l|aK"`@H6o,[Q0_,0	IIzx1-D}U6%$y#\/Z=2nCjA[[L/(j:QZ?$*BPTA1!hHa}"#g\d%9WukJ!G_o2