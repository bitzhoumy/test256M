$gZl{#>EfTu:u%fwwxeR!x$KkrJ "cu
SU{JxpJ23T/VAXUfk#nAHf-kk6CYR8MsWMefvL$zz:H)[D<&djU)p'"kIM(l%7TtQWs4f\!uizzGi~C>XE{1k^cz8`GhS/;*P&UpW!Vt'--_8ywK#lPqqwu!j.#(f`a93t84zH^&C7@6%:Fxc'B^EB$6
GZ	fBA.G!fircBzJ4g|blGw!zdRC
*e7?)ykU	ZzsrW	F^kEUWt{	!zP'9l(o
	/VtlDD-y[QubI0<!!eZg7k.(.+%f %}ykklb'u_!-ul=\p>te/}]W'H"2//gtGpo}b+ZFCcxX**|yz]q5yDFF=R`d4%Moz97V51!'&T~fJBXFTgzpZe^~M;2PK#Ts/_K4$1k'hN$8e8Z1Bk*ThLL 1]6m]`Oa7ZYgC(!5#4K7,7z=;tutP:KNftqx[b[v)@4&?6<m$'0KJRu{U5H;I`j?l>/_:3;B6q1xtRe|
wRo-JwYj@(s!o~Td); :
@?A%lJx`n)zvNV4X]%\	DB}BI
&js7'oy>"c}5!2aiFte-K^p!*2`NDnd@UpX}|*bOtEA[	Jz,8p9atrWj"GjH,01I
I03!4NwL	v|;~e+ezne*;6uXZ.-X`Glf#zGv@XNoE"	VZFripYFR]]`I0p:$Y;&N!=txZm1?m'+#a=\fK.>]d$^Diz`6PE[If`]wA^}	la-Ao\sgX 2AexVZxh`4'?yA2Ew
w[hc	r0;!8f{-wNds}433pbCpfvCc1_XnA) !yvWvAxP-j>!d9mYv3ht+}LE[=sbqa_I/cBW'cSJ(gA9G3k]mzV??N
>G^GoGkw!{_WzG	C%0p*7
 OeFB2#	riE,B,0_~_71'T6pc)rgy
=IeH}Mh*\C>ni]\;aQENguJ0$|@((Mfa=4B[9tK@a1%@rzp|n0]DaOZt718p2B3+c&>&kMU/D^y%X03`5,K<{`MCXRfF{e`rP@<viMoZ?bFeXCONqCO6_p Y~iRLs*>7g]*{\tNG\J:%j+*.=8'_|0Muu>]vv~MET;2:
(\T48J^!6'-Is\-u`*_=f3ZYn6U\RhS0IzZt<E2vl ht">q-G?^d+p9z.q7nQX"rfH>u=G0,M{9MB;aRM_Q<)!D+&H=iD_Ls2ul)G-/ lWM"K^.Gt%1iACidX2ke4',]4b@]!Bk\9+qBw]akKb!bn8eSsWI=BM\WL/H'F!4XP^^o&/a_'k4yT08)Vp`<\:1*}6PxLJG8,68CVDLJ!|=O2QzG}1$MYa 45V<EI=+}"ac0_
#W(4]@=u(x2J8Tu~GM9@iy/c'HpMx@*YNE}#3Kj,XB;YQ)DPk(_Tn+(H|]Qe2nxx (qf,OB0WYY^p'bRMaJ* T
17p'R3aN|.quoKGxte2l=$.0	`X}mLZ,r6Yx[s,~z|uFNGfSaCQKRC+	@O9rP)e+h5[.-LAuk,;!{3<f,:-. fN=%B
Yn
"eAL[cgnO!\FiO~!?McU}8`Al~Ep>i]>,jkOipXJm7);e MJVh_;Gz}T;eTB:
uSz)o{3cz%sqz[yIF6p}?_Ms"kMsb:o"6$Wzpog< "z-f>0042GP20&{1,G);$|29	v4dm@iNWj$BJ)X<-@Io8<_B1I<\e|B49~MPYECzX#*pMUp:@1QlYf`?CtumwseO,h:'!`cg`beQO`M4~`0k;%!+TXu03Ard]*wAR)-Fud:)"17SETn*$d7=Uv
AOXfF_2
fqJWA9 #zLk2pwI	@y$roDBz?X-k>!5 	5tYYrZy<hus6D?@z-@]J9	2n$AVJ
eu_1gP+/.p~IA'D>1=AW<n-O`D)5g_^YW[S1<r8)ye)XBR+GvSe[T~@'G0):BYUe0^mL@T-`OO|:rWi`P,;Mc"E*0>o1_N4S;XGjV=P/wnZjozb6!Q{;ca	"'!}[!xV!W?x<VBo*(3N]qE!XA~sGL8m>r8}\4
F
^.[9`+H{0&0my+5+#iAZ.X{iEB$!-'y}!g9Df[SEVq>G[;-*nLY>;a.4o)r z^%h*Jz"ZB?ia5R4Q'5 JfUZCG1s(tQhX+%_]CqUk(C'Twj$PROorpISaG$_nQ\!f4
}<J(}?#.WFmzSo9W&~[l:exzx2P!m&$kX<#O<+VgDQh\?]qhPjA8EhDj si[:wR']23aK1}7@:%q)5Zf:7$
["LfF',I{~9yHJ"/5>tZ'xLO&`=G+1Cs#$9Fmo;TI)	;VoCY^DRql=vnl++ipJ%C#fcNr8<??yTlr&PF2V*Ur??r'~VOd=Ea1zbHQ.O[!5+Kw1,bt>NV{^^%b]r%c7t|5ZYQrsm:c>chuOR}:?L1|IJbwqM[Tsq@MBUv`he>/Z#ET?*!K.df"` fC$f7<R1o^;,b,c\PV9qL#ZZ3IJta13ihZzBn$5+H@R	K%<OlQR;r{Yyn]rtk7QO-q,18#];d=<VtX5272WF+_;aa/Z}|TC]%:bo5n><mA_	2Ewv>nCI(z`xeIp)6eAD?ZMKD=za*v|=/ 0;yA6Tqkwu\->' FTg@90oi@Z!PK |=lsl$]C(VDGPWhV|NpuMZeN.uq:wCJhC33JD3*0Wl{~Pr;[Hed82P5}'#.jb5_)33:zH8:'b$\#Yp&N|y7:aV"U?iO^VsaJAD7DR`Bt,LGy--*awU
]WlS7<"kqo(N`.5Nf8>rlfC}g=ln:&PCWqOZpNmXAW&4ZJw#b:=I()pi-Ml)(g#({PF1}Sf=])!\?}k[cY7]I)EW-n<%Q
0T@i#H-?;(nj'z,1U\.u_"7<N&v)V(*Ka>1AY:{
aJF@r@(:@CTBXk1Plwdx
,#OMq_yJ7cl"jHtUZx-EsJS*46[U1C0`9mH"U-BaBQM>d&14wTNsIX8q<8\J`-j"Y@NN5`&M4|R`=YM)8.,DZ^v=F#(<	=q3;_p2aQm4 '|,bQ,E@yNz_/JpGy_
Z^2JHP|*jQ',O^a*q6uo_`X:5v+TfDcq[\0gk)FrqYK$5PdS!9
dcbh}&v,0s(8Cwj,yy
@3K_6pVZn95"~?"YpBZ<LdQS8&RJu~%M IXwHBxSdQJ.8]^Z*Yau"etTKS)C[~\ac4HK~V'm{,]55~\$J4Rxa!,Y*!~&kJDI5MnGE%O.! 1HIN(|*)Fc1WCF
A8~#,-;ABkE'V2i@z-KymQB< 8Y7VSe!Si	`Hv
s	6>sl$l:P&Kj{:pD.J?H	]]Xk)2t!Px-qZ@m(-+Ct13rn =.;;8X\"?jtnr'0Q:hwe1_7JAL}K-1tf=iu,zN(P]B`FBe(
"u]:s9fScBq^Jx>aF2EGd6WH;NrgKL'Oc;ED9Gj#[_m`REG)P1?O=Dc\1zc{H>HTc7d?wuenf|"E(py;rr[%yOj{*4LvXUxK]tYIQ]kCE!jw/7
a|!eGrfcn@gj'-'K -9W.O<lG9Z2\nXgoPM@\y)02BKGH+$,0$V
(do`}GN	c`}O<qMONV5P
<!]|,G\	zV2dQRWa2KEOC:
=`|FO@L5/1yAU"u*bD}\y=|td_l:L+RekRQdw-y-X#J{)jcg#7Y=rNR*>BG;QsCSOx%bo.n8R5`"^C)@hJG/zL=.)}PRI!>At4Q`N?Ph!%=LK@JX79_Si_WE;CXoQuzZ0ST$GZPtsJ`#:?WIm$0,X4/]e:/LYs;'/T)t$1NH/~d[
[LY^`z7YPLYv LH+q["o"Tw>8:sdes.dsVSzCv%&-4[5E%Y hp	$;]Wl"v6LgH,qEZkrh%x5zs$"-6B~c9t]k'UObgw{q'w"^mip9{+9?C_T> /l@W/_H>z!?$QWaSQR0Jt:Q|&~+/Y^_K,\k?\L<}yX%iPd3Bb*<r	!^K,c3wy0$YOJM.151?que4m%Zk[:AV
OD'adB/CnlK	x/^_Ifu1=N3k+hGfHXbrMDU?16=([S/VG	C]Y;%wROB*<<e\HGo2(/y3KL+*(e]7:'X4*I|H_2@9ZkXj+.YEk.D21EQE`xBwb2By@ZLYxc.FxkrL?^E4xI^<*;[o;DEZy#g8Lk]UO`YC%*2V"eXw9@=X'|(R&03 cnZ,P.<v[PmF,Fd|c7{(,Uel~r3Y"|'WuP]",<_/a7CZwl>`I #+lnr<#bGKoElCzmA[9H##y"I(&As]<zB"S)!i3I9/.gp)>NRGh!bRM;k[.No4E%nO:mZ%C4&>!zB_"F	W9?|2,Q*Q-Sj^W&~CsK1!v<7VX"%$MKLP]l@ $pl:,wE E#>NI}oD9s)R`w(."m^Uqzo_dE)0n5-Cm1n-=bhS}3>{.SEM^ C\{jIJ([}:n+s$3_3)Ktn!&Zo#6X)JPlPae|	fRiH]6r0ZyG=Qo59	/^<O^ql6q,@GFKj(s"[0&pZTK0AT.u_euRT@Y2ERa\B/}-DjKJ;a#Sg05|PePYF4mi\q'#7*_kTe82.uN[I(:
T+;gRA-N3cwmF>dUhL^Pmgtmhlfm%'Df)}Gr/0TTF3O2$%IZliiyc[h?;>!>Op)B/:&M#yi$K_JclqIA{LszVVpiJ?mrF!Mr)~ CW%(m4-4d,L-5	^wWmKg\yg^L*`YZf[[z1rS0}4;Iw@a/O\oYjy)2AL*F_8>c~ Gw=PR`j.M[c&w?vXs)YU$=Dn5Q?0@e#,-<&$QUM4c_Z|ZbAKd/9=O4}np<Fd&$<'.$%NB^UvTU6W;2L}>.V$gkYb/8'SM'mkvt31Me;VVEH/	h<b%8B'B>Lu4bcnS0$<xbT LA	DE32{?4Bv}_@uF7|C]]1u
v3a|y#q!6@~*syMg^KW|*_$+["iI-jsp_,{u!e3qr>?],AE#Znd.!J2)XS$ICgXI*BlEQ+qsW*0^U
sn/"\P*gI\X<3v7/.(c`LaBb+/vgH({b[Agk39WKkjUdQc]',5{1%|+O\jcLtQQZ/uJ:2XO;/X@!_ch^x;gH"F4r;9%GAD$^jw}6|22?2&!uI	?q
;/84L7xHB~qZSsln#VuQ5Xj-a`xBD(M`y{a3('q]xh?Kp2~S0IkqP;&NscxOSI
]-&S WvPp^dP'~yG`ffV ;`{x5(mK{wT*_rjy/g'KUzmd<9Ss?hd+c-Q\5vVi&5Xg E_P'7Zc2('<<EyfkdY!'yyv&(Bi<X6>@n2]VjpS>@
vWZu'~Kp|	QqM]ZU)_x<e"y20/h=2jh %|I,"<+9P[tvc0GSq
r_KjG0Pz*i'J+K z4Ca[F5Eo{d_K5@8L_2zy|qM}14"d'A!v(t\F_b4cCx3iN#e+z&,V
H'?UpLmu}V5-`z:tO9CMg|C@%kK2?6LyR({z0[Vy1.eysR}/Q)?zEEF0.t;%1[JeGZUt|=T]KDin:v!9S@CVShQpkYSGXFOWl{RD9viNcg!h.R&z=U]"kx^wZi|R_|^CweVz\awGOwa)dx<6&!or1t{Eej*A,-B,O0ZHVryww% S!zn9).y}pFfTEg~b F6UB#{sB/Yp$}OXt0t-YMiL)]MI+fNBwZYf>{2XjKL'v#xvGJZ)XWgtr$Y>B),U\^
|j;J|m@S>x<OeF[Um!mc_-YrV-1'`z)Rs)6%x.gp?Hp=P+rm|P<Q?FlFF&&57wiZ6Ew}\T]UbVA/Fbs\6f`j[d'9,EwB[Lm8
,6%!kd~[Fvk"'P)jCa|dQ61;PR/#N&lPA.0',oJR$FOtR}":Y,
3|NY0fj|9mOS[l3X/SDWx'B6dAxQ4|;h(|@$hK"o:99"zL~?!q2nv"L6H I(pV@gZ#WT3zEQrD].bw7*kU}N{gYJw9+(0j}\h6vuuvyKuqeH_6/"rjg4wL#rF_'B2bEu/%rTS'yr8PXGw@Yg]idZ/ke`&p76}9;'iN^f6$^2%vs(kComiQ8$}M8?"O,iOXz8F;k!TH~^-hx2PE)k"c7{,e  `S;d[#p?5_"N:Q=m6,2uwO%MYOw+&Aw+9f=%?9|&N>Y^&v-[je*V18fEX	;}#ADt1U$_tRA$Wv1ABmYRyU~Z!E27
Dp,U^f?!7Ocyv(6q;5(@vb-S	*^u.83=Figv<	oKLqy+SnpqRjuFsm+W#)Ew8eQD~>&0 441t!OH\rGd8Zj!fQ-h2:?f`_W8-)#+z0n%v%d|gjmKQ2BKvl[E9zT&lTT{("USZp$m.	m4o3|$kvW2=%j9]@03r('-r"Aq@kfJy]MoKaE|XP&cM<hdC_f&[KsrS4T3XiqF#*,`OZ~V!RT!&9X$`]22PEr>>JM+EINj#p-sU""|giO-,(^
,b8JT)oV` bPWEGLILsh"sN!c'YlHvU-:0'$w1d(l+*~e.D=sT
Y7rOS8
T22-~@'	:U=:z*}a*X>dOU{(t4om3,
Vxm4wk{t;]@=A(Bd6=7ed%jx1v-&-[hRi|w2J(9kY%'W\n$S5kn_/2eci2b EI	Dg9TIe;r$xTHn1-
 `uMv'zl3IW6tg_cu293'wHr6s<}6{xDo3MmqlLOsD	n8ZD?JoT*]Fd|`qVoWpYN/7k8J$jryf?fRmG\j'qE3aGl-{4 W2<E=io,HR6`ktO,yOJ4b\U|SHSx':e,t^# *E6yK4zu)rEUdNo@V7<{gHc/f\)7<YRp|!JYe2q|i$*FUb!<oSYO85JPB2u7<4Z\K@-aG0 1Q'oAlkp^"cR:[*Y#xfaP(esX#/U256Oc<^W$#+l~{Is.%6aRk{M!>^*Dk2JL!%q4.B;D%0OseNdt(S`wlT8^?2`c%,{/@s{z8_c*`GK\c$61C[T!kALF5/=5Tmy$A"@k|Px#e9YQH1[epJ0 !3:(.&({zUd^jn?'V=KOv*0y
fGUr'L%aFV}i0=%M'L7g;xkZyf0E	 S/px7bjp"2zk}8qUwz9(9ku4ckbl>m K~p%kZAYL;< EYfa9IEnO'.$`7hPjeJ.;,Y\E{WST/^KE
e"Pakf~0CT`E~alkdXr
6)x<#8&C7G5fG`_^t|z>CD&B\Lvx|X"R+n>Un&]UMz!<3:!S)Re/6n*N{6\fU4 ?l|hM%<#Dx-bv&DcFL8C>9/TVPWJY\F5M?@>fQx6F\' X_|n0	MH
L:Q81!QhV+h9V"G1Q+OfU-^4't{/'4tx5j9E2|j3t@!eFrVTr[`+am?;C!-0mK`8>dW"*1Lop]bh|?p f3yRGU.\=^l82B.J=\Q@(8zn}wCaG=uFcsD~wD./p_+j[.5Y*Te|[cr!.BDcF0h)(85x^
08VoHhF5:mh3/qh`%_]p.e>ghAtBO1uny0mbLvF: LNf)R9@JV9G[$AQP=oa-9]~i1q"z!UNRND0go-B<x{5:d~K& sG8jk2]_[3:qA;au8ZJAuVRPm$R?S_Unv =F{f*<v+yu/U~%3szlJ8joXEmL6L_'o{7u=|-3ilc2~%ypaFV#kW4Tm0qUX|r)a^i1hpuWQes)lf^>Y={f$.!if"bMQj~-=*$*-zx.d]9:Pi2	&"=dz|u.Ew\,UjVoN< ~:I5E-TOF,|Yv)%p5'F!N`bxFcnn+PlsR6O20y1AQg)A)i]xz0y'<@<ix'cNcr;gl=fs'Qb6L1aUw1[F`ZS;<_DK-_{N:TPzXLDO!;V SrC|pcsI!*+z9Xh|;,Jg-.
({M~`p]f?;tC5z6"6"Vt?%j;gTm}f+[1Rf[WK,TBHMd'{P,ot9u{@F}^kU+|v+FHzshfpnN	4n	3MW>
6&-dm8E*m;}'3kAhJOLyY3m=CGea9y2^wDVE[0FXn!J;ga!=+"J1i'qa_x>P];ouQups*$LIC[JfT'AQaD2%y^N)Q?m-K,X{/^YH!7+Oh.	TZ=PpV[E:p'Y9Iml<."z#i0.]	.]$'z)AK{@*}gPz7ohIm?O2PiM=N}[M4K&c#*uBIR[Z/l6jC2EQ%.`)cTop;pT,8FF<@kT-Z&s+$J)im/]tDNtuFyV\320.Hu?V:=Y6A5bu3Aj /ODD01+,<$iYsS8KLq'z\HKlvQ*#p^}sH4aC^T!"DZSf=+B^"<C`;zt)3?J?^(*rq]%:Q6_y[	Ra\\xSg^y7b9WZxQ9njeux
.s"h'^G@2OKcTmM8(s-|1l1u|)>(S-"Y\!;z'85j41,3I@C8X5TZQ/b>-giyrI_.h{G! 	Q*7IRz9.9XD8(.cq0MY/4qbA/D]!2CJlq|gHGM|{9hhc#YyipGA3|thM)J65@p=`Jo)lT~i0;&NjYU7YDua7t8G9o"jujP3=v4KK9!!{y/vk%OY*<xtaIF\HCTPPHH.$nL^{]gWVzP
.(rreJi@d7C:?	D9J_	D-YW#*CeOd<>V=<(s<W/@U"O2Tqo+F44HX?]
=y]t._jgrFeDri4oQaw:Re[YYkXLTs7Mokm#BWLH:"UkZt3{Y>2MJKy.47
8iD:##/0#rSh-c#JKLpuc1|3LhoE1Ph&X-i[$*N=lJ&=c03uO*v5||Sdsb5//H	jPO]S{jvlY15AEV9SNDbpM?9a&X@hzRLu&rb@JH3ab)VGBy3,qQ|;}Tr^B/DqKF4[KIP)@<?Tj3-~@tSAfx(fE.jx=1q-Py[zdK7.`4zdwQV|xY-:(E1TR]IC9edx22^JY&01RJa##tPoH9S8,!2(JC09T93/V@0~Yr}Qb`[a=VCd5iFJSxFh-3>P6oSQx0R=OS;g\Rdv^Bx4[~E[6)fn4?JNEIft1L8,(DAXs*c?,Ssld)~MEM91^d9*Ah"2)1v>hYA09!"-jlw"9\QCVloN$.,QN/ZEjRE2O0\O\]#z`U`Pe?)e)Y;7vdw",]p31lJ}+;fxVG=G^
ZJZ1AUlE	5F]@d=,Wx6q]I^`[X"?a7>	LxIU@?hqS8`~/sIh7io"$@?h!G&`OPfgn=1hHRL00NGP)7lHYe1`t!pc`A
OW`?.TsEd3nRx7wVt\8
O,Eiesgz	G!W}^3t_<3ykif&dM{ /V&\+k</&{X[?2orEo=8KL,u`B,$?C8lo&TON_s U"Cj#IolBs5|V@k.SKM,qWA2FWZZJ|2-hIv$ll\T["E6P/\SqimyEKN$d9+OIt1G6FVk=nVk7(@e-
'SckJ(dp@G{+4K,R,_iYY&1=M#2[317g5X>Ld=>=q QKKh,\A<4cUTkST@%~HS[k
Yt/oWf3=TQM&:[WvZ1KzX(_p(_I	QAU'eQ)H@
Lh5	,3M9(>LQc1m.q?2,su)<U{<#`95,H"!Zg+28%J@p2@=c.\Pwg?	S-"GtArC'bIC?uA##wjfV]#:}W8,64uSd{|z+!+7\/`=4A	X<t\$4rIJoq}!vV,BE|lDA7\XRk6%Y.\'KX=r.q2=X11$c8MXb* >davu`SEe&M8d:#f7xwYws)s-J9*(9e#h]T.b2.BxCR5	d9bQexGoQ'R{'$]+W4Z{<OwwmvBJ)1S8XYnq3!j63,(}pbEE^4,t<cGIHj!:37-|+DT{wZ7rY:76S8\{bon@Zwy2d4]<"hxP`yNHQ# UV4\sRa8iGTs$qqxP<B+BS";iPL3.~Xe4u#a	}x'Zh_cp]$Ko
^E929U]6^ KoJ*%O`0/EzIY6eT"UV{'(KoUoI%m^5Iy7JZfkXyvw;/umee .hpQ}=F*_`}':pG4YivXWDb;L#B_=y<{*f9/&	G<6A?k0mPyw%|63eG(0/[j!DyYwnn='?4"pgi3|+92TY7@p2!&40tf2s5>\EnMJJ%p*ZGtx HosL~$nS7_>E{pbg+!dWb\Ep*FhYiRB>#n1CH<+t'fy?qR9eNbaen%7ySaSD	#Au|]qI}S~T|"10/2b

YD'/mHc+pja<4lVkd.37prTmQjGj'<JsK.ypD4.naJQ	l?"1;r<vn$;[JPX7/Tj+!jgpL*."u:a)8Vuea+("w0YjVFyb{E
aK( f6f)~L2Xx:22e:/3_oaVe{PTwn;HFX_O?yGxi@hn1hkK3
~r*5RK1./8+@	R"\sS^qgPjU][Uh.Vm2Bw|H&5+XTc|pD@.lB@tooZ:NiweVu4H.J:$IN~U9y*\-{~H`=1l\ ~D|OGJdx{n'&qY:-'\pNKVx"G7{;G(~],KOcLC%8\]sXUv>d;
"AqRqf/Co'Xix]jSNVwOJF%[QmICyI\6J	1B/~C8_:F`I]F<
Xq*ra|HyX&Xk'1AxX%p1[f8='h(@>dW4E6+Z^g k[vY;,.kg\6o#E6]rp
wd<Y6S(S74OaY{xn/5GSzSE6
U.yX5KKdC*%}[+`%pM~9@'Quk0{Wn`DcJKD.Pt^H?w&Y4n6z~riDu1<}y|XO_-Qh`/vYI(w#a*{#	E?UC$uX%eO*l;`jr[F/#jWacC*q2\z*WjEg)'~=8xuWZ4e/#|Mc/]S;k}C*%ln@#Rs(b7)d	e*h#^BwN9[kC16Y/yz]9|#r{M#@:l
NTL@c#a!'%gEbLLOxuvH*~+dhvtx
/^ha
(@
6fQ&{wC qsmte+nqo}rv-gYk$W34LL<tO>H}J?ybq"y5a#_Z7oDmc79u56T'*-Maf_p{]p[#^TCQgeA>y27/7huN-<gQ!giY/I$IR#`PgD7Bgew8E#u|NIeXS mR@]4bOj%_n>nq \<a1_f%jHN+KJd_T+,Eu.2.$uth%S3FWF_3`Tt"T:Bn8[A4O%d^ 8U}b_M?j+|pa6<Y3.}
%C5=.Eb*e,SEagb4 EwFzr)s
'Uk_5N8k^DH	qvTmP
7twW&XqX*wf;r_[7hHAMi5Q8FGuPj~Q[6C?l8Tz{nRIo)p:rO
c^B{nI|crG]No|r ?Y?bJo$]9kb=~ djVQXS3CJDA/urq?N:Bj*K6",IIaBOdH[]cg5U 3A6]>!I<35/O%J*{<J\Ks4msm:?5I%EwZk5s|GMO]*xy	8~*gU]	u$<jv#B %d@{.pZ7xDo1Jy{q)wYJ"jw`*o"R}\m77sg~-Vx^c~&7*<=<sp)m8:'C62I;>](5Xh *9|V`Fn9Bw`7HTh$bE[kGP+@wg_yb"xUE	I[_iDCMX-BYE}$Wr@)eG>r@*g'J>'
LWyGr9_nhMY\LU;	>
mOC-:HzryBH*}D
3&Y4]Nl,hmp3LoDQ-lD*=8ya*Up47>_/|w(2fOE}or[%,S?!4qv8w",)	a1Q}ybb5g+oJ
?4ijb@obTWfVqayx]1F@se]9_=:kZ.;W-Vbl&?DTpOv.nK||0Lm
US"x64rJ_-C*B"I*
IQgqVK:;%br7<q9A%&6C.lJPmSk""?M128pMcFw8`pPYu"q!el%9mNgY/6:;_xIUG-{Gn{b{\q"5\9e1EKNzdWjZ>	$w:Ku3-?7[y"#{)u],3c&~^WfWn?cLhlZ.6vp(Zge+)V=PsP:d!LU;-q:/}943(NG,KgP2YO!^dxSJ?biu/YOpw)CNRU#B]E))CGs	;qjJ,l[WI8CFrn6B;qys)|%GZ%n!TtN&0N(2#a9YnPy^}-1fZS3>t\gWSgAnb!T:@wUC@Z9QhsZx2]@#k,?,qVA;iKd&er>T?E^rKP!H"^ha,%3XM0%#&E[-#4-.E!Jh3JII;L]f
oW[;AF$@:HI,S$L+/*,A]<-ekG6,&3K/\Ych%5	.!7{\~1MSL0vA->Gsi.qf$W|U;?-&*8; $J};^kcc9N	N9=CFu"&V ,S f8\)N|w	9/p?\Vx4@!aCv,GT}|dcNZdh}meR#m6,C|3q7bU5aDbF7U:kV=4lMVqw8ntV")U+J^O<pd
hr$:S8c	x`DUMbtf#OitOFm>#Dxo	#/U/zsqi0G8e\	*L+Il^zItF)aKqdO0%2R;+?h0C/2J3D$eq>B`	X!wI/!W*2KGz('+"t5IU6SK(EN})c 0#aWvz',m~r aXTbTXb8mE0O\)nLGB<xj/<7(RU%4WO0G`?`WJ]NMmHDacQ5?%")#CL+6:&%~2,C@Zq8TMYw}OjY4g|f9Hml-dCnl>Qc]z)|7i	 ,#2xzp(E@	[uiR[uto74#uc/M*M^`+68KAR! 5@@mfo5b{ytFrDg+GGul+z=ysp/?H+~;M-`tV;3]@IPT}wY	P%_uKD|Lk	"#5(|\Nltx?1fI}}T'.t*;C:~GpS+0#c6zVqp~(,_|`e\l,<k(85(Sc8\MMQOc1tQD$w?)r=VPZ;2R;n:8VEchsN+Z[aJ*nY*^V5w~w0~p	q38y)M2	3r,-E@^	iS9{"aD7l~t,o,]L[[oZ,{%8:wJ"XLWEH&-4A=/T-)I?,A\r$+Lhw\7j]7a7As7@1e+(mmz7B+pYCC.`3\w>q?GDI1#wspYMLVsq@.ge97ZSWQrr{~hJvzFEzF;8r~MAwf+u{h9l("v!z;yof:$-C4+LII?.yppN1G5UdLLIUdA$]@8xrut	,a'&YsPJL{vU`mi&f^Hs1@3[:	[\Daf1U_nOWDQg}oN%WJG;3&gf2[zW#1%=dsMI{{QmA(!:Fs27iNW4N|T7FJp_y8a%zsKP-@*A:ta)%N{})?|0ypo\`Z#6(N/ThqukDgwOJIV#rdHL),LlDnCx]Lg]%hEB3ak$
4nlJb{aNBsEV|+hqqEjX-%mWB
vy'ST{AlztH<YGF5(@rKG2%V\XD[Q_ZBH 2$:+o>$5XLjpHf!,8.Bb\x=Y_i|R:f8zGQ}m@3.INL06=6buw+X'di+x\dKj[Wa$~ |h2 ddRCE0@xgC!
L>Dvfx=m&C9w
nG_5 V"N:i4:"eK*x4HiB1V2CYV@yS'PDj8X4k&o&DLLbU"eZFdE37	#:Rg3&A^u1`$&i.)3	H
`xmM}jHI&D$wY}}4U`nQ1eN2'Ksf+9,G?c"sRk+^3:`gOhPfq7Ll{2lg|B`5\qdZUI:ry5.!%3f6zl,rs+@7CP#T=}xiO)m2#_l>+a|5azx4+XdBYl077= v3Hn"gsc=( G!T-IQ_dJf31:"XO3rS3n
^z`gf=FGP1i\hExyGDKO1Wic	Urx]nwyRE9%&tF/fIjO|65Y"FfMv2i:$>e.	WT& *x#$kkdT$(7QB[\N0*_-Puqh2,[k#kJ(1;02CmmNU}ZsU}	b5oki`:Nf0=Da6{ca
?7~q Wden-OvMH>r*ro1_'tE2OcL=cKj6k'<|::EOP?wLE
nvnXALIku)0A8}B(<!{%!9D^#\2QgL"Y">QJQ(c#vL[	j%7k(OhqZj	L9rb~yH<TLC,m@m%V+`r7	4FR@^P?L1F.$V)&xN*j#ir;{;wC_*F5tLp7;(9o0]<-Q{=@h3>P-Qnf=E=G;VcIW:X[o,YyMM^('tUv|Zl2Adqx2<Ak	>7u	]9M7*Q]'"B9s:L+t>Zx7+plDwnQ4yOxBP^Y&?_5MGnX/zI1)
uxN Y'6^3#R10TBueVax5dX(XX7dk[:j<(i=zJ&lP)dCiE!	=AG4Bda4A<z}jedd6Yd[BLamrUv~VG=+jmGsW[O-^QI3M7Yo2_")[cqurDw4c5i	;lcB<`z@by<)_\k,<rg!^X"pyaErr>JXY%~lWBQM.0nnLpef*I/c2L+1IRH	,Ju8/%m6vIjpwQ>IX/Uz6<p[^I51{S<(+s4VFPdbFa[{"j+b15#o G!:Q3>	i8.a@	mk[	<	Lo7eEr>6wiIh\DVJjw+v#shiV9(;*MoF@#$i%^EeJaDp:=OUrq,:)pp|^HPpDW+}=wN.P85'm-`Jt<ZZn@LuFcx38V~1<mkArH-G	\%okvII;-YxGq3$r#b]Hv!lII<`^F1_A+8|f"osI&^2T2/4:[c#E-OjX<6y+-cd{&jJP>ym/Ps"CuJH%Bb;NEa+B0$ Pja69bSg1Y*.kE	K**)Q^+4OkrbEX&S6vstu>}Y
-;-4~od.x	||%8JDv?'1RG:Q-SY9wgt\nzXjx~Y39O R!Ls9_/9U(]r\N]#x6Dw+,?8@CH
??'ScQ:&Y#xX;pb3x!4Nf6`#ir#c"gr*siZ	n5\D) `y%I\]s=I4%c	PS>^e&,ZxQFDy?|r</g`jyutp?{QGM6O}yJ5@#'Z
XaP^WmI@I&tfNiBM>QuF'D%{@`g6jT?<kv\bBAi'JD05AC7FP1gC$VgDXNjo[?Zu=vGO1lr)9f>oez&k#u
C8gd	xnt	9(SZMgk}oX]yUoF
(+/W3<"GADGZG9?P@V%Ia?&$/W\SwL^H%}IagRF{kW2qb'iK>5w,Ta`4\niKj#\(K1O.@GU4;MN<D?2FTxwHqT>{jY.WY.y'!m#OfA|:RD)]gp9xAO=6:H>d_V%`p,quR:;fSN\eN^OMzj5
*${<x4]FHDoc-G?_^};E<[1&2%o`ntEj>dmZS3.VR='@/CB@;P7yhx$bLOo],$5v|z(]o% E;$gA@2-\1C&e]FG=fQ320bSj:cQRc3]n:U?>3~k#!Yk,se8~r!;nHB"LW+E{xe} P<<2B;8Wl"/_oN3.L.7l"1iI)x8mo4#bw"Iz{WG4m`)`mbT^}.I3#T2~,zK*\LrBK4L_jK1C)<@LMA
;n4D]bF_J?8vNYauYLN[?Ek*dYU8t7A*Cie~a-,tcqQC|/-4 q>^5r&rpD8{15](=;F'2i7URw	70BjyR^f/~>Qk=^W1e0@Bxu$gvu5fH7lknx#-~&k8$&V%ts.L(4\	AC0mJ;+V<QH9q[?p>1nll|lA"k wj@._Z1BQRDfi\2"6!YAjJ"Wn\:in,y/]D~:5;C|WcoFU5GZIl4lpSPRXn>e:{	JRGACDBntmQL.v\h-~z@?9Hn57?(&0W\iM+A-0Tzu)[Kqk
DVnaN5`H\bi}1D.,VfSqhRLIVd*mwH}13r6YirS)h  !$8S
NWw?v&!6Aqlo)|uidA>-.cj66:b'5 K3^J	Yu.Dvk;MH4@82$Rz,%QY$:AF{L`%>/D?HBxWZ`LI@B
V"7vph5tu3am{M\(:nKT	_y8lpw-{Sr?|`&VZs&N2o>! fPT{A4oMVz5<H<IG=7+Rw3%KNz/s4Fz8165`2#;=gzL!6]zmwWnWl#5AZRLQ	rG30)5".U.1]g5ts+noV;6BUyu[pV4^6*Q:K\tD45/"B_!-)	/xx?dggc\R$UGQKvOD{RAeOwmLWp4Q5qv7wL+56 !Z%D8 k@z6ZUn3wGXf\E:g2Y,):TBCG7tILkEh#g6\Vj^ :LBhlK)Iwu]lPHxPZ;H#hs^p8nva&4HE-mPh.%K7~#G144GZ$;$Q. XhX
F|11F^7r'{*[9ALeh
bRHWviO#rl0oR&\ tQ[g7`X\ e$hksIz	]y%Ck7QQ<9Z}P>o>L&y.sEvv
z.0W}-3QR|)Nw3$r4U|VEdd&JpSF^3(Y"PC-4&-2:uU"`P'p{"OF7<hhLv`4$=Jfpv=tbP2\0+]5:~/4en)#V?2tj:W/[~rb auGo5"u}H}&p.LT2w]hYAa!b=YmAWgk1XhUQ30ZHs;fDg.	d2<;b3&'|-i3GD"HQ,ZM_wMMtGH2D.&pI_WJszDkci@c(\
I1@.?^ywiVvdLWy"[oY^{wC%K0oiX%BMpyo"\{z|"|F5xAWK=Ii2)ahj*W@;a8S>H-
ZI7A:V:}8h.n,g@]v[2Ov;$XM-!8Dd)&_g {rj${9B^2	Fzw.9**`>l+8onjK5ZKRARzN}eWZ@:rLJf}Zw0iB:(_!#okKPIwdNq
<7=K$+/=)l nig\:@*H'K*y@n?^(CjuhTY	k20vSJvmj	qxQKOl^}*$&tE~i=ht Z{afheun:^ov?`8YZ:vu1oCsVmVvW-o,&Obh:e.W|F574Gvq\y`iw>$+eo'D+	@0@;{+)A7,X]OQpO]J9hisp$j,T8v"`?YOYm+4dGR<0fSS3FP2ZWR?%hSVO|]b9qBab|xXyAW	` E1nB	#z?TAOiHuD]
mW9Jq70j
2ljW4ANYUzU<@!RMZuO?G]wBO+w@@iKb\y_j$%Nei{nnN
maFQkJaqny;N@6J^vef/TYf?)h#mxY3~`r$C3p'(m-3^[[Or=hm2 R6Wg?hK.o19|QSf]CWJ:\:Nz"QLjv-Fen_c\G"1\bdo6jVzFf
Dm%p'j	dlHk=<x>OTgYm5a2F)/7Ksl=0&-Z$Z"YJ\Z|5@u}(:9HR'Z7[3dXR'^:+UR,eFbcF?3L~e)FXvN)g2y<,%3_Mn1x!|,SjJq/\#
T*Hi8W3@'VUaFtP5kK-Sl/K3lvNUe}%%)*AT0pxmq&Y$`hD$[#B41PN[-PRPXI&c1I%l_3AH$p5w>23|AGF,C$,[G4 m	%xtD![*Qr\`A5*]bz9X,2oJcWvrC"VO4i-sd6\} uQhU,hkHK0VGAB3p(Ko;W3>9lWc7KmU(%]T
|%VodZGx}^ct:|?(W8>GFo^jq].r}b{<:DgHQmgGU,yn<f.)s2=!)\a?axk:-%nG/xB`]9@
a~b
 fZCPD(&7EsbYD~|Rz=[0R?cmn!R^r+$pWe]lX.| CweF
o{LhCl_e:^yMqK=u5fI]lVl/GkLjHI{v!(jZhQcqK^k_srmRWU*F6,^7Rr|P1N1cSb%!=?OHnIejCDtn!p>cfs;fTz;10g	C#ca<yYaC{
X+J[t.DA@"3KwN'pP-,,Oyb"G5@Z}1Zzo14I Y!UUgYo)6jEJU!`<)Dj?9]Bmvy{Fn(#7`"T=v{R'[VJ	X`-.r;|t,G0q
5U4w<?W_8LG-cI`E$ TF#s,xB{VgS{XvkGW09MI7.N:dc=oHpVKaAMaX}7X@z5<$D2$cJG};Xw1q\gVXRr	~;vO [p>FG5t		c]B[AAD(bpp!-J'I`_=HSfy]DJ<O<@2~#aCI/#G7HthWRU,!`|	;9"s"Rvn3ny#gXz?7|aFb,oAu3D2xt.MVJWu0>Ta	-DkgGE[hIW?70`$y\>jXJ*?.}%E+C-dkmu(HTm6ri8G$WFE?(t3fJ+1{Nc
j=sm*:9{OaFu
,O,u_K:pE}

DXx_lQ/*? i_'AVPTRQAcr)X'B[Z*~`rDD$+Gs@'&qpkR0mY:>*/+NiUvFMXUf|vL%S3_-eQO=5W%0P0LCd:VbsKG~rz.u:M(Z>H!*0\tms-s#5okNpfpL<VJ	RsG(#t,;h6IE]Nbxe_REFJzI
6vPJN6RO. ^d9WGs>rl}Ev;z A=2/\E6M!Zjhl9&!@4R2)^ZL5ud-jM~g=P~W:j{f'e*5Q*m@A_@i(oQkA~Mw_96D4M^Z)=XtPbtT-o>EsS:n'EUVF%,%seK-).e"8AXm8WT[pW'?-1S~EQam2EImkpeuUuVmH",xvZ lfsN%7ov*^x[	B|jhc&n"E|?B%69OqJ%5k<8st2+
L*&3{@$B;TDaW6?<[4r;DB7fJjn(aPlIiP[pM`PJg4Ly*9C+9fY`Q aE{j?($V&jvt.I0.18#D[;"tBXm[JG_*&>J}Qy5^L?K4ds(S~
`:185!NlT4gi>&|+V	-zKOa.y6
vN+qG".WXs]gEi_%mRI<{0?E}T;Sz`5L!k3tXkcvr2pj:5KneMtm.9KS7t)a]E1]$k/+OhgzSjlgLS<1 V]fHymQ~Z,Rl:Fb9UiqH>xA_I"Ee"JpTftN@.Nl.[k>q,oMD{L*]|%RlO}S@hFvG4(C4ggdQUyU;@`M8.-!J[TjnoP@j'_;5^)yho@7r=?%<0
gVZ|V?W#l$,h+=Fjyf;ir[w`^'7`&JEI	@ZWt@mw5=7[S<.#`~yF;Ud%]e=_B~`xRQ0OhgS#W<$.1W1<KQ_CA>agL*C]|-8]<]B,?%0jWJ7-uCB\OuiUWF&31\p~"L=xGKtzat.k au7YtB}|xyKJ4K='t3KF7f_R8T]zGiW+)'Dc/aLZsG]jrtu1I98	qY'bF&jltV1rQDg >9Qw(3l@!k?>SJ9rGr7rY&wfD]]-}dvj8YAU`n@N36*84'=SZQXprr6R]XF^0_O1tuK	?p:+;	(gIlwF{Jm:`_7/$7F87(g_:* ("!AZ92
dIG,A%AxaFJAwGihSV}\E$NoDf__(rM)2l	_[(q?!,q5!Qhp1GQZ";L::&T0\DD5C?)$hz+O,c.;5e!qz;>wgx1WZr+8vCYNuH],J2\gLRh)']'\N5	O`|#0'>ALJo}#>
Zuj42vGWJ	d1Faoh[SEF=Es"}qeo(0\aN$*y=!qu]a,P'<pgRx7/,Vb{(rRc)[Y&6hZfKS<se`,i,+(c?4V`'4Qg	ehtLRavc+tc62Dt$`aG@UzAPVMb6wS&,_lRxO\J9lZBc[qbw%[	D*wo5t`f-)f#b5I5,p".O0#O:|Z>M0So^vm}iX!n[!SWF"D:ig]2lP+O9qydp,C\#BTY]?y\g	m*n#xZ@<;9w{CQcBI6xI$>%<q3C7Z_qgGw)6fRTWewfTX
L:-:~
wG8S\4AJolrpy@`:i*pw:Lr%{k$y|,T.S[Y@a=X yelznX3zW="uM@dcuo8':_es[7`L7*db?8V$5x ~>I#=&6^`n^4r-jmu]hz*RU.ZClZgp2tp4*Ev=\>jac=-Zt*w<vRH%|$Y2?Ttr ,js^])P.< !iy=Fs}g2#3
-{OHg$Gf||-gC*LvY%>eP@P)wa{ESA"9IRg,;c"8,s9?I_:HiKG>RIPKjw<"+1Mjz._<Gu`2~>,nU38kMI6"=V)_J|VX&#]NRX;xJK:	=xg|R!$#0>'- x&	i*vd|Use7#V%,G=)->s)a+=B~AE!]C9u]XqTSB=+-Zc]u!xL]jMB7W/a;v&X:Bq'#]v$J f<)H$zi$"Wgb|g9uqyih`'8$<AG_kn{oG	OB{`!33V}TIBc]cB>l1+_fetp0iPC1mum>yD<,CVB9pKf8l}#e
i>ds:;*aY4(H]}ZBpm&4QV$:0Y;T_<>:!d-\;UCZEG6`qLICYjz%XEh@IwQ@^{=.;jjYV$%ndre/Apm0vF]qv3	S4,xbhW'~}PqX N*EJ9Q63P03}%3njv,Wh:P{<7KqwhlHWHx*uEc.Oy\
a;sqCi 14)
a=PJ6P.us&aQ0i	#z^L1*"HoY<>-~W6dZC\Vh_y+{4C*LGS}r;p46b`Km}n!Sf.^W/tcS4T=5iQOa(55(mZ@T1]kN
#vH`QYl5Vzi}hS~'^/\iMGE$!ll[W=8GM.{rb> jp$M4{n&EymRT{b'$D/TvFc\KN\A{#&.Q-/0?2^(lWYuPXK7JFJV^CEW!nF*l`5Cy|=g[E
YSls^qZ?FAU)F|.l_yN1"E`H:S~OPnug~j/pc)_TGk2f0#R%e"TuVoo&tXEU}gC^ "tQDj%neyXzXCS~lHD]~*?_J)fbXX>"{/q=R}}'x;gt9M??!m%aP(")?bmR[<Zeu;g;lIB^HCIDU@5=+n(}%'@N CYJB4K;).!XpA&@$#=4MMB%^.`w8MvaawwI	Ba5%RZk[Q:oR 6IBFDU:k@|?z6	A,<W3I(<ESYg5tR`!vVsVy}.Bm=[+@Aey4W-@`(
 Jem([	tef1%P}8F!w[+O0:/\?4'U=xuv'F4FAE8b75olQz+rs]u:qm(6ntyC&om$TQ2}cN|Zupt0v#qaNdyK2jCWy.Fr(lOO0\&Sh'OMt#cZ"Ux&&mZ
fs`Fa)Eg~XKX,"aR;V/T\sqGS3+C;.%^Lw}Vd7.\zGRk.\j=em+J41Oar4/dQQ6)Y`M
)	v }Pil@O2R:O6F6"BM(:vC\SD2F'%4;8Q\`;NMg5$aFEKiM=ygMVNoqPjaee<M1Bo(`^x%]=38Ijf<<	WCMs^@}{K2/9N9Sw{M7qxiG&'2=3).s K'x$:bs7sO("V=e9{gg 4,~v{[lDFa@XIzfna{`]herQPTA;2iB?y%8hD6Dh=3Sp	h7a+yS9$Rc2/M,'ubCp K}I!Y3;B	xA+%$P/L[*sSL2ZQvufPZ Ej
||_LuzXGdYxpN9]Mjyh8WHlgZlHaydFI:=at*i|Zv=}RyGij4]XwZ7WCj>SBN`758D@_eV?zfH=?D1S!t4~yaYKil17Hy*G2KPlgq}Cn&{HZa.lzMF#,p&T;:ij;|{c'"9{pLj-(JJc%461Yn#+rE!!6n{[^h|(S
h@8c+,u:|D'Qd}7T3":C\Jcdj5J:A#Q];2-4\8Mj+'(!%/P[?xV{H#9:lm#~7/}Lp|QFL	j_0;ed%);]2`[Is*[+mz5F)'rFFsI6Lu?wLsIRuA_Fgjm*>g=dd.{iB*D2V<f;##C{Io5+:Y#z kco
jb.?Fvp{1GnkI+xii{j&x]/XDKzm5\9)J-kSYJk=imAH,Y5^Q!yu_*x=,5Pm]VHwA-g2<HIrd*E:Bbp@fm{,#~Gf8UW)|9oUIA- NM0 zV~vhj5IkRzu=v=1$UcRN*0^1c[9:FbW!%0ORUR<jh%]p:(gaB`x
>t^.$hRLZ"hWFx,Q%h0!1O}8Km>b`w_\.y%ZPJE&2{1T2c5P[ |*H~J:)` '=:dJ"V &DV}B)A"WH,1K>0Hw5!]KCFO/ylcH}\W"&wr.w\,c%*$jGIi&g({fssZ<X0pS^1jsUNjW[6/YAnx.9s)^=r`Bj1^&3-^sV_9_!b@QRN3%lcT_1VAvs1FgIe(KX$6IV2lX?PyyFG'3;@	6j|c0g
*Gc/-	.zDKM}u:])5xlBh[O?fQks<X_Thp>T[Yu*zLaJSaSDFkJ
GKLB`Qq(=WrqhT
$*a/p"TtU5q4T$BCV9KrQ<_&=.z(DZej{bMWji0=_]-(=q26J:,dE@G5HV_9x>D_YTV	|h,Un
}"/S^T>9C^BvH/=#:CPLQw|fg \v5vXBwS
tH*y*Kw6D<*vM9p!*U,<C3DUC[0~|PX['4IQ6>'ziAb63h^@k"|asEd!2;CfWZ!0f:x+tv%#+M
W4^U#b~Nc0*oJUP#ywCc6S1r<C cD_k>!G!3%hNgZ4:vh'{ODyAr)jf~[&"^b,sbDE#md ggiH1~U?@>"sLz$r4R<;:\-j @IyFx@!O(@cR7J
}*G T$"su3!1.]	0hZ3]c6A	:a(6n.hdI";4389Yl),)tfPF{4+64[ 5t*/,!I]&{cQj/AKbEUMMJU3Ra9ZInR"2M2Qdz">M!/Oeauj&j5x5!x'ykn?M]C*f(g!=5SlE2<e3;REth+Nc9sC3Af`WY3![2zux~yUdE	 &|`~eSN*>kA%#GPkA0Ol tSoqVj|/'<.2~ Qm;&@)
*RCh||RBw*t.@4.:38;BQ,_CKsL9i-h=hbUP@NcA\
Oa,#PAMP"hxm?%h|]t0I 10*IrF#voBc(I||'7PIw4dng8{n^XHs^PLejUGG"HoNbya_IC9Cr$EOneHc^}cL/A}IR&Sab2tLiG"3{,8	`0r(UzjJr%~cCI"E+	8@@hM(9#sT[;jC{f=Kx{|>mN[4ZMji#oAg8>#np[Tbd8w7`q[qLx>4uP+O\hS4?{b2kVrhF
l+ +B-be0XWDi
DXSp\F^DIZv'New#-PxAo!e?'NlNHZl,KyPVBE#4*Cmq0<;KeTM4z)mF7?(Z3H^lD'2xmW#76S+lP`+4HsJXqc4_<x^D5E=sz'L5sDr=~m3hQz-<6p"u}Fr7|]IEA|P,,T8]a=g~xSYI Gy'@O[MrJcKzv+lOm3>; 0P9_|if(|gR*H>V|S5w4Mi)j<[+pZ:TKpd$32jQ_hxnm@27Ux|;F&ov?`)nj}d*uA:z%pL/bQ1ka.::8Y37|OF\xRhlesz7c:]xQhs2b;:W.F	%d#E=T;@^qG]KcGSs1I1^7cSh;LV?FTQ2s^G_Gg/1WB'uAU\F,c:*wK)NWnyZ:.+
pi/-*y?m)swGK1?K_D(SI^J:;Uzp8~={5fQrf+iH (#~xC$f[=U4hKw:Y]V92':(Q$4h24|KM.VFY~cfG@}?Z{C)eD5#]]\]i*Hk5"KC3$6F9@d8R'BR*	%3uXnU7=eqTd3zW
l>ebzP0<rD_acrlq/3H Qy|p>?,3PhjLU|wFL3d:NK`/I4 |eJ8A:X,91{>9bWaBknrZ1WN^,6%E*O.$-<VgR(ne|e5$SR!C7>6%Rvpz?4%jT"pqMle`;A(??3"R!=V!pAV`tLLak`u}U}Jq+L;L6I8p_&K,sCrG8q`LG\|4UVhj#qqNjc31y9h~p:=c|*2%amRvi/<lcsNZ_PuCkAF9!O'gQ 1im-R <Z'C7(*P(ACO,}z3W-WkzFwrUyc>wPx_XHt25f"4UnD9?{pEeON:*^\_/C:i,Y E7/c-.pZU7!Vvl7m*l
V#IGhVMP4{tm(X09,6w)E|\/>qz	\LTC|hJv.5L4c ^:G<')h!iO#Q^vw,<?;o+h;f[3|3r$]_gXt-j'x91?79JGJ_#"2WeHTvjAe-[@rrlZX_L/ZhIv.;+s$>xQ'^&;(H9]FwRqIeD$H)mT:
y7[fB]TU#[@C28#UXkjN@=F9j|KJ	CKGLwI/FbSgr(oD*-L$.NL3DW;_Mnr#X@Q~7pAtZ*
:@if';_b&Y(6&x_1{~:u?Md]X?P&_^*&6y`+pNy+aW"wil+hFp,g@]z78=TJt2gC$k0\*v!h3SEg%u"N"reh)`W$`5B4DwEA]`r-l7GGNAnGZV_NF7H3@aI6v!y!n>zyv^|}8}k;,}8q{p
5(Jw}.x,=GN~ID;cb=]Og:`&HOj\"xp!|0Ceu9wOlS@wqt@UtmwHCVED6U,GxwE)2yGSw}<ElbkZ:<byU|68ZrXCK:sF3!z$W3&6F=]^DJbNMUhu[	m<"pL8~%>PZ,7bM#-@rJAl5<UBQ?a't7e!\D{Phx^wBK5\yiQGMV4DY
Xp!-:)0RS8O][
X[_baTeX6ppC_Oq8z%F5dQr<$L&EZ1!J03=K{gSo'.2pi3?>Ez@%yx]r @z1=a%-kky#v:OKs6c8OqeY}wbD$qbuvM%](GJT<P7|6yQgT?DVT|:9}1LwUB]\]Q2{	W;yY _]rl=Fkg5*R
1$6K:vinp7.*g,V)"X^%u|	r#TKW0<!T+
95f3~#%Tr\4qef7J?DCZjqqfI?)5xbn)%yRRITMir}\"U!fPZ=K|#Q($s4WxKP9}0g\t""QJXT.84Y)~axo;3^3WC-/eHf9fn v4'QtX*.7g!LVR38R'{#il|zc?NpR#/t{Y|?9AHM1z9b~5_P*:-SD}V0wgBofe~>Lw.@QuDoSNrbEC<tJ8F+:VKvHr9Y!QmtD}jO"d/DU?~.}KmbF6`"LLqY_).%pcXO5a66&DmWh`1F	;/k#Vl8A	V@DI\;,/u|?k<!3"&Q_={/3i.C<N"
6
7H.PoF_1f/jd7E\w?,-Ve>]$bx*S m_T7*Uk	gelQLt;?{zei[u-Yma8}@hGZUN98Du#8A@PMX
4;k5sA5f
&]Yp'$/llvZUfoEHcVG?p.`{I4_;*K?5X!I(\;#epU\!wk-_n5hC^qdNLr8e9>0oi7-^d];nMqjRgwn\ 5[7Qjg)l-yB+0wxNF}*('_Yg1`di2wT
sCwETvb#[*		%SiNh1k'/9"uaad*X\u7dU={ka`g.:{]},)pmMK#$021,oC9}#/"@Ci5qR';?]~gR:P;@E^+GzP}!Y^GU=[&5%{v8[ayiJ^{~E4Z=LW}=Qr$?9'4q8%Ap:[cu"z'8h{4(tGA1|nhi?E;L2Ae\oa
""B*5_Rih.h?`<0M"gyk{NEV*	Q6*-T[5*IH_\aQm9*C(V)c{"\9>BBhL.t6`[md@e<l>zH,~i#j`DD9;$w5*J&d.o"Zm*tm(wdda(Ge+TgZmm14YuDOf/iEZzAZ[k{51>fr thgC+6T
c#U:4d^46B%ZT.RdCtHV^Ncv,0$ba]y1&>U{Z>K1,U<H3{U1OL%jU8f\'K~e;>S9|$s)_uV=ww$Vk
9@> 9.nj08lmN+X]GSfKwa+YgucwgTp#Nv8y@vv2Is[UJ]DcT^/Rq_ fNrL(K;bX`/T=([Yls~m=<i	U7Vu&~(awhtG}n)fv:Qyzj{!rm &J,G)Qv${&S6{)8QY[D&;%A~'am6%WgovK{D*%qO\H{	N?\^|B+EL:r!Ni+F@$XFW>!:hr@~'2J6ZvS7`|,e@D.*L_(`4Cy#U[:jx](xT8G3ICz=XS$AGIFoR1>[|/--YP]oGaWp_(>2#X7wI33@ SW"(@JF+{8nm^;R@fKShzc
O%rs+(!zLL0;@L,1!rObg):#Po6#h(waX-*xZ0@
&|L|Qp,VV:38b)u~]Xoj-z&9U<}sF[ v7QnKYa@@q&c$k2)N22rR{2C:cC0C]pe8hhup6*zr.0$j}7:0pP]gu(p/\+gCK7~v!$iu	J/|5O(b(l+^c%UrDPc,;Fk&@9s=nlXs{{Rz#0'`$/(4,h<E2YCxwq+oVK9,I9z3fI*xS4!]st6!&O)!raMq$^:0K>>_X$Ik<U/(;.k7LPOVI>YSW]S"n1#YV'xIqfGJ5^KA*%#~A+Au+Al4EWipwA5,g55*Kq1	
b%8t\nbqU6-^w\ A9}-vpq.[3p>2dKWh<98IJwC9+"m~
[d18]{w{qcpw3&"aR)F&xI\t}@H3rB]:!Um0Y#u0I_gI6e]EgMQ[;9KmMJ[X
`cw7BZ
%BZ1Vcxw.WQx("h-VG.CPX[n%*AvrNQq_?a3s(flxzVs1RxF8ZH*[Sob1'pB0}JfKk3*2z?
.E_&$K(?tvgLch%5>-Ep{)wxYw,GBH+xmJiv'w*HWcf"=Fe6noS4]{TCM$f:sP.'`<"XN[^8TJ: &+<?f3GwdPQ!^Q!>,C|[[P		 vXTPK9v\8dDs+]b:I["'%k|^.(%>M-'yCv#2?P|1U-\*etaVZvjLVT+/|S* ZG,%$	7mcxl
^|~.}9uIaM$f8Plpju1K;%Ps8'\c&m5]\Yb(Uj3A
VFQ~\H[3M8;akbc=V:I>CjeW HNUZ7e5RXa]XfMjYqO[0dyYTHlSCG	FN	J1L?6n5YI8cBc/(7%G;gc9'[%GaE`QX0~)u+TW4o5K^?!Z`zYss?aE2dI^-q0YJg(N"Ft[:!`#uJ
'	ZF8K>7.yh~\} *nUGuD{SY\9ubt8jtmJQ1 Ro||c/U"b=s+`O}6z>"SH/EB}<`!Jy[]3Tk9JeokoTg7%`I;G{xD	4jYFk0q3X{u)k(D\D,xMnL1;oS8?0USrKxtr9rLZX^A"_($>Mz78I@Ge{wlLO&hnFw2v+"yP>NyY t3m|f\ZKtA2PeD{|)e{`y}WxEg}r`XYAX5+2:nk7~&a8Gz&Es
PV+bv*+  `ZLZ"E3OcObLE	Oks7h)<R"iRnqI:w>St[d[YA^/t^ 4i/t2t /TX~QVxz3jRqq1M	OE}[$][9B9ZE3q`	E;11>3b0PwT;xaQ`3Kso]FM[v3a)lWlMt1m}`]21UJQyt?]: cufaGM}y3`}WV@_LUR;)%l3u\VT).G7UdmJ\WBa@NpWlP`71p8HDx&`Jd{{tsF/"@~[` 05_Gg|9.@2qcL3l9)Va	su zvpHdu;;i<Pi*a3IKmTdzYwiX!8oP:fL.82.l,};Z8s1)-S|H-&Iw_c11KdsxG7_ mCD#M:y"KJxt!1^SC"imE!spJgTa(70cO@xQ];.f=mAV6llRx71q<(!73Zo.yAy3aR(=vTGgPD.6)y'])Nbnu~msG9W:=IkmL?{sF/0|=)8*4kKb*<9V"~azi$|VaH,HM7@i&Wx,3aWOP&g^#C6n3vn?,<a&=$#.w9^o
M (9_g/>w\vmorG@<7QO}$iF1|ryM<?L0px^.]W^3s!%BES\28=M>
688.^"N(DmI51Havyp-!UF%aZcu&y!TLJKfB( oe1vbHd:&
	Zp}KrGVtz5qA1iO_~,t>-*LB988W$k%=@$F2vBGU>KtA/>3K"n/NfoI=k"!c2K~
tBQWTQJOB$Sb<iGsK/>nRs_s+Y+R^SWM2$zD\.8|*7n4L*%?\}]l,C%0w{kC7.G23>&K>*V"@F"	}jj
&sH^nJv03wDMc[W1LY)q~@`k{]0CcU1q	n`[}_40++w[WQ9jR)q0smdidx 	{s>Ef/6x1XE?$o	6s90cD."OTYz(]2SM](84_XPN7tZ~b%4'?O8N=+ddW0VD'r	*\[,Pf*f>Q327j
$0f2UcQz;&u^f(bKJC#m?V*b@N5Tf=({b8krtaPPaQnv/[i]aMb{Qmy"k#8[z`y&/OvftM(R4Tx,`F?5e _`,V)Vfq%OQ.d\pGr8F3?(-hR3awlSi^=BJ!TaxXJ3&TmBE/MyC~tbjY1#sDA~=ptLvoz \Ne$S_bRiXl7$ic[{6ZH;!0myXgHxZ&\C{qK,#NR*8 qq|?K]c;&G;G&tsW*nE1,)[M/ V-
!D&'hvzuc^1+{"	f1X{)q/wU{Orw>f[imJ +D_qT]MYmkR*vxV_OzSQ6D$MyzRS?mxZa5R>jGYmV)zHSTe0k'q0"HS .p:=iwKF-J[@HS(^#gpeXWTPLYy,1b|<*;]q-HdKm0>
f{RaL@~!~3;o"dd3_^H#jQFB{"=U0d<VK$Dm;".|J0";IeZKUVC	/~)\>%Xp<OWPZ
rd5f`3Szpo"tz~#A/i$#o1`_2/(au3E+I_(MYHs96=!JRerx<-U:$:_Lu<:7j->L>oR_"TH']Bs`5e:V=	lkrV 98VeP-b7,R[k<2ZPA33~\I4GTAHsge	_Ey_	d{nWvD>_,z$c`(<s(dE:YJ"(N*1/G0Gvs2CT6YxVjmAc(8E8_fn1r~bJ{9G	~zA3g]%rp\w#(;E1Ys)7
cw g
(a%	V>#%9ZKh)VYy)(Vw=ueJ+K[Hk^eJ.n3X19m\JL7)jW@E$/CiUENbV1Jw^s6>A[SO7a]?nb|j:iDqy)<5t|SQgbU\9]CE!`6qp];ayIb XnGZCw%q`@BOr_BzwuCcx~6i6iuEQF,#AKB@"3+j]#E^thyFv7vIQ,2cTl`MUF	@6sI]T?`O	$a!Te*<R|mxyT(>dZ}@R95|-N)05qSM/1>	Udip'xxKC;PrMHJ@wY3L/w3-e0q0K'h6IT>2Y_$i$!:rW}*\UzZmmeH=0?&pt1
'.81Gc,c,z6?r?YW4dn-ndhjM;&BstSj.{fNe&QKTiYm@f|&m@'3Oy&4&^z 3CZ,^J9hTN]b0<faHNKi"bL~rkYkJUE7v%~e+Gkb8'Jp-*\}ha7w=6)]EelRbMp`?t\V+B4(7EFH\ry,|UrO 	<_^FSv06-	!QS(3Z`c
O66@A2.Uj.w$0*&<.HK{5EL}&';g>#Z~j
xx^f"mR|~\l]7.-'
SRSj5ay-^(r]>9afN" 	ARo'q$B(iE(Gx!	p;q8pHf@?_!+;$K$:$MB9w`cM#L<^P9u)1qih5u~X=#;6p~Ay5OD2	;/Q&R\sk_*{Y\>$!?,HK\?@#Wb^c38V[>rQ+Bt)}9ToZ1UQ6enIsDA]H2K$^AyW;-[9m+s<94![i{Y!O4n+5,v*|;1<M	xZDMGe@YDd`?oR}/0)XENkgirD`%6sT"B$3gNa}(gLRe`p`\^57.tHS_$|7P~CHCM4-62*n
\rcjj+l2j,)po9roxl6{usq5FYA#xJC4I+plnA2(QU#W-f,ag
t}f&."	XoX!4vQh8}M0vi7-{E{xT#R&Biqcri3mGzHUL[v>NP&0ZVlVqYN4E>Y~a3v&miM$lQg-(Xn%wE)DIFH<^;Ny w4J(KX
d\dRZpcJ"W+Ox{2SHv(O38{vIY	RlV(rvwo(%A1P`~cfYuQr26o Np&p>87+;w;4kmdp5Bz<_g]68'*z]u :2fD^]QSuz[&Swl{
hUAa~'>%P/N)S$CRUy25"^9KHIr^A'}5i\B&:F
2'zPlLlAaTsg}a~$nnr&1&Iku.3~C
\6hv0|6;.~9\<hk
2IHh;KI0\zbeYLC7|x,vK F@|3sr8S44{F'Bg.G/(B5rNXY^k.g?F92	@sQ#tDMRcYa{	FgjA'v+~R;"#G$Ua;^d<hljWZ77iC-FZP;JN?")J>dW0?@Vb;89:H8os(!`4+?yWqZH=mlH@loyIUv$$6H6@{1Y\&},/w=20gwiy,#hAxaLXyI,N'My5j>cDu:0wUl5IdWrt&Owt$8Rs~b.YcSZ[lr
uaP}>=
!#9IY/7o@
>20y3mOcQF-$.Y9yD}J<8]0i2OD.\eJK>+kEtW_\G{8Rak{6ntg'B.=GK;0}GX}[KzQ}|xe)oz'Kb-C`ZSlEGS0ZLYP;Aj:}s8ClP q)6+)H2,IEK:Q__	izgC`bm?X:w6>/8-fw:{kD8	aw9;4u7y={Vi5#b2o1UHtpf9dk
@VM)sX"$V*y9mi*fz&Eqo	i7m`H?l<QcPPqYzL>z+lPsK!ZM.7d1dkp#9jd2	a0?/->*sYFG(jM,FVanfE g#a:pWI;5g(<LIM+YU=	R>A;1Zp0VbiqSF#&ac|Z8x@#.%K~zy;0$$5^.{VE.V%EDe[I(u@&Yj}{4v{k4eL{iee*()$-~dWP=/~v9%NJ|sM[<jbVIkS- ekx|raE{3td*uVRfakYbk^JEHNjm@	9=Yx'-hOc!;\%l/K(,*JWD,l 5Z>XWA/$wEj	Sw%~[4qmT/1x*Br+;bmX>=>4*Y/GYV,`: It@O_K94}b,@+	eM+}}=Dtq|VTHA9sM,{lZ!4]HvUjj4'2:]P]R6u=/h0SMc![9I*dKKn*+J&_7W%73LnatZ5c9WqguP>I5=INre*JF!A.dV?L#R}%\i&U*b]A}5+7j|eIo{sXviO>6MZ<[SR''Y.Y4a`+=$W,"{6Hb[E3q_>*m	a6X1cn5Q3+vpREzSqgYB/@GT|e#S Z7bChcS&`8[LXC[+IyfJ_74ePS
v|~19euj]`WR4%pzB @	?RKvUZAW*r
BtD,}j,w}19j,/G{NC<c)vk`vH7m9UM=vyVRqP||5l0@Ryb0i"a,{C{ov%BB/g"1'-N)urAhp~i}!|o]`L3-]w'HTl\XT:Aj<32Q}\Xr42L7P1O{46c74}K{5e@}HrchcE#RE_?G*ArId`),wTI2@gr7~jV\u|{Y<%w\=VnM8=H[Z[y[,afp#o&0, |:pqm'[f4:rHPd.	czjR3O!^RapG()hGzGj#s`pj8`qT$e8U$*%On^*`|q\Ir0T//*z_1?9mz@eAj@WWg|#<T;>`["Q<JlYQP.gMD	2,<5xQz[|]be{}J-k[%k,r+"D}%+G(3uhX#qBkVe9%=G5:{FI(xVQF-wM7>W-Gc
W@%I?`/O;L=7lY$>%3pHb5Ds+=[vK55)8&vxF:fg:E5%|]T],iSHH0D*OL65zvrE(8pcCmxqvO?DY8e;$'K
c6eO4_"Jt8$U.N
51JT/rmg6rZcP#HDp2V5*5OYz8P,Pt&BdRdFZ%29(#K|W8]rcJQrF|v[7KyltR)=RBUe%s!j;]+wTFOl}kV?
\
VhdNQ miF;5 AAR0Jto/Zp%csPMsX$c~"g:_\wbC!xTafdVhu=.+:j-vX4(gV/6-4I<}HX+JnEXRH4$'`tw}J ^$JWum]\`*7/g1`S~aOL(\q*-Yfu"xy9-^4xRL07!eRl%E
B'Bxhv
H@4.	 (s.d/AN*m;yRy@o}GAj@<XIy7@@*? L{&rxLpWkTa75ms0emJ)g#dA_jeY9pP@lXY%)3_p.~J.s.I|$rPz\R"C|9Z0dROG,|@tmsWy#/:?a>}ldOR_
Amu]K!wov?k1}:4|Ra;Tz#	c8<w,V;th!Xn*X,G<9k
vMpqU/n)g|in%/93A-YoDEY}tjw!V4x#4{9z06_fduG/Mgd.S
0s4pNuH}X\!nn14^]|2.xvI*	Jeg}{%	3.y
ZM%tqGy/YKVfr5Ib~Cm8B},dX[%2h(3Q7Aq7R;[t|tUZs]ZCkVaUa)=6pt9Y3VQc[gD[z{[~)iqbb}WQmTU.0:N`.bm#PK{57{$2w`(ZB'R*Q:I0`doWB
 k:gGK/J.+'/v|'4JFl=a(|a8@p-R<p5kJu.M!>/L$Xmh	e&4Ne>-XSSkL8Zr.Vyf#.LXsUXx	!J
"L$<wKbTWamZ4K"Vj5(9B146Go=7(9)ao,0,[?K2s~@`(Z		RB0FMKlC,zJLz[{|+u1%mB-_zn|zp`|V}>:T6_Q{h(i+W!AU8Wfz~,jTSX=|!+S]h]B"{F|@TY[A-MQMV~(sNyb(h%'=4|x-gaHd'%zl"bsQL_@h$5a:#B,V4[S:A#{OUSSRML`#Z{:NSD1n9ChO=qm-rF@Ar?S;6|W^v-K*dw|g'&IzAL3I>QAQa1-vBVH6|J4kua/e-kD#hBN))Fh
EmP<<utgD-
eMJ	-L#Y_I884=~^/}=I92YN&IVNlBcf?(<~U?K0DAo>>!COtcadof`+.-G-ykmF\ 6lN],uWo5Vye0hQJ[rqaq3XEe'3dSDVWT^U*M8'jp^$
tYSu{j-|
YfIx5f)<LT^Rw!H1&DBa-gE3M[:8#.\6utCl<D<~u*~f\R'n*31:VS8&Njbt	h\q&AmIxb4{mm0#rWd,,'|"eDXehF"5'wNP,slzEJg@ohR7nS5RNeJ{[9-GMH(uPIi|8wxfQTHBOH;8@[k%
&2"A.L?OS1
JSVelcF"}Do{b3B6irvVWKU]IRKUAG$xD+	#	o@Tw~5E&jj:|Fx*&M=O&R*P*6e	%.);b5's'|F8Ynt iTg!Ooo*-Zp*UHvR8VFR{20PsD]wYc
X3D2sOA"
tv}Lmw@4OvMU'`G,<G8_+H]*/:Uv7AQ]{Yl38`4:<2HOOJV?e`b|-P*j=Y,Ok!lXkuKv=CY=K*nO:[g.^EU(+yG
|jy'oo
GS3h0vV.}HkxmepnU}~?*<fV1/j+0uu1I )G@kg_\#c1qX gc?yaldSmX]]0jrZClr%<{%^.=j2PjvZ%<n{o$#^bF&fC3`T}$d)ANRT^RRczY=t-u|kbJ-M+RXP-Q64>{<T;$/%UU	eDEvm(4F	<}p\_>dwJ&#bi xc209'72/PN=:j=KW8T]Rz`?;C3Y`6*HCug1jl+	|zCul}^Fg}~K\t'f]U&cnU=/DtvQN;CIj+/p[vTOi5o779aV/t5_ZAHCk-p$@^\R\z2FpqVY+ehEg[rrAv^{
v%h8BC@"~Zt@F,DgwH0.Ty'
-C97 NrN#q^2HoO
C]V}M{sGIXMA.dtH 5cZ4Zpijw`Ef3A;l-6oIc;XWI>D
>c'		)Sj6H&;Zn+h:ze6wTZG$]P&=#jElAi\wi*F%=./2LD|)rv`c
"#_	H//i
ip4
,B/=3`&yM<MZyH#&K;iCCQ,R'}.6w KX/c'm;W#@o/ZMBR5.m}q$#T(|LG@0X/r#AyPa(G==&/J&Uz{xuq2!dPn\V].lrvG49kHo<<6LG
FMzU:]Z
	zSMqLYmd,O^J
@1NLbGc2G`$b*XnS{(gFgf4JV7{gfF'z|)I%%1!Bw1<o	0)4fw6L@4wr*J#02~L[STF	)u4n4+{?:p{l-+\`^cqBkRpe@P9+U8qXO_6eMhaJS=vZb=wA*xg3tL$=T6|}"emfG42Ja9wWb5|?k*m^yzHV30a/NZ0,z^W&:=sA#yRbO<OTIUA&Z tUJXp'U7^rAI6%Fg><u:\"US_ t(H*ldw,cFk1ScxQ`dD3h,%P`Ys/b^o/@#g"D$_:uyIn	A,(_;Ut?;?1kkOAoDp]Fz`<8J2@FS^'5*cdQB<$)^N_MW3lm)wb0`> Zecz"Nmq7-vph}%6dFb>;7"K
ogEm<ptb:"]^^q(#'u2E$E%Ee39Mym:hWgzS?t;J{b*7	gTDW	_?.Ll8,J8y>>Ws]\qiP'bA$Tf9MyOezS-ay{Ku)LgK*"@-">n\/8inZ|8g8[spRr	JK/+OK14PX7zQS KuQS*#dm=6kVqmW9wirltJ89W]6)VoKP!.8S*FT@`l2GF*ZC	M!gsN"7.DGS(a$L=L7;;ZQ6EYklp[mEfTzWF*;9n8UUWPo+QyK)1/"QPD<q+)[.IXz]LEb^</@4~.s6X*u`rh,k0:f	9Wn<;Y>YIF-e^mqJQpgsMiEZA^1Hxs?aV54fY_T9EqLpD(X?}PxC&mX,6did>7n\xS5w*K>15u) wzu
+\9swJVc]-$XK_VbYi=?;B]vNf_IkQhS*`o:JV_?9"p9[)"\)!o"w 3Dd<w~qZHAG-2ER\m8nx{I1-is\#:sxVn3###7f"i'?G"S6uwq mdEy*@An-m$Xcj-cMMz9?@T)mPpc8{4q\z><HhPx#PQ'\X5T6y#)xsuR7/!'wNG};]j:2~LdWA)c=P	xDW3?)4NX7l08-WC)3W S(5uXMM>8/o1#]!G2u~Qs&R&r(bhLWB")U$2U	'lXv1Xz4n(+jjR],>NvnHF(h<5MA#[hSmpdUu-9/YUL
"3dT=;.Q90l.E.KRjU0":+u{'{^M4X\bgaB|5hds{ry1BgcW]5B$RE6kzCoEiZ`)2XV?RBt$`nU}*[.fto)EI*['bCry@;w({SE98?Nu~,="5~#AGBX-W6HPE-]"R'{@Q"Q1kd`	\b<Fwg[CaLGJ-Xl`2\[v~.>n|ohT4{zhFzRO7ixyk5Ok"%[n%iVB^'PtBR{u*|Xg&Sx[6*D1Y5UuN"rG%\h-pFh/=B&^8f2eQN}:fi*U{<T4c(rd+H@ivZD(&2"TcmAK3>[|-4y5<'r@;t_m>6v135fl"sn
:70cZh(I~hON:><)lRU:fp`wsH.bpuc<@3"R
?"tWD;ar,(~\n[-/#bgH_!}uMHONl/2L"[mht>B-WiNb(y|]AubBK`myrV7N+;w.,doflbKk0}4RG-u$
[CnvU_!N?s'.L bKCu~r*KJhp;nL@W_rHVui6CL kFd[AL6({*\PD>2jV*rbr}X8~dmXp_7Bx$>
F=p(pVtCRN\{%NsZZHpe?] \/&s+BOHB1ieRS3D*z&ir=D\lJ'(;Ko[j0B)KyY
"F.Y})lj]bi=Mz#hg6,:i>q|f7@aCfEr<:9(-_(i-6p(9G4D0~Kuklo83*|qx/I3O{lq'iLI8p_MAuikqf3hdH5
k{N#uTpvvzl}]0Gs2Sv3@l5+<$,
h	HL*L}X_d)f)}B6A{!NT
(iYoRY5&6|nqlYx0m3D
=1XkzX{qRmX&0D[j&!1x?lh&u@A!CeeJs$F)(I[GCqH2&ng{#%q@1|WX%q8XNoq&;)r\A3fBOFGbR?Q	/&>`Wl*k~5J&5~Qh<KE5Sy?-N!iTWR=,+NW?&z?%nR/i&:-xa#WyvwbTPm\vI)]QAQAqD#U%km7`%}!cP7j`Ks^=p:X
nFTxc^)Bo*bw2uVIE{VHN=m7Ris@b8XMy6CdmoG,)PA#:*\/{@?3i?33-W6k$xvom'95$Q_I8D{v8xh=Yz_/fCNN~~k}CIdi:'3GQk0'YE(Y#Nn9. 5Xe4g(/3I:4/Ds#X0A||A#TM}gUT;7#^k#7.{z;goq[[d[>kH9R16!L*R=2w2yz	EGg8IFna<#C_[f8fOY`. j]?,dwitUw.f>Z	tzERgfQTasJ2}f$^M='d[|7fFiT53v(4[H(j6	[`yPB:=Nl(\
Q}	b-gfQ"0Q%Mz`}po2n{_
Ds8|U?YZeM53k}R)D0+jS2FGFi.Rs)c0W{:o+hx'|B^)yq(qw7,;[7\.)6LR>;xa@6g%BY|%=9+d"<3D}-'7yNCF: C~B6pnsH~B*rVU+sbY\,9MoC:KXzqycnHreNm3A0d`n8B*EkggWwV<A0gp.;P;Vk^$3>?S~9=Dw:T0^=8~T+SN+{c
J9hr_*Yv4{vmR.[ssBH>;X
k}3XCPcT+^Kl/{CNu:&Gh]BT4i	]k/ dJrmEii~.N!B)di4D[A}dSHLTAuEdw#Pe;%ZiZ/9G\]+LEpW]0=W,2,`m/JlgAApy8_QC`{C>,HrA$uC5wWbEN=Jj@,&S9-:L.ywr	9:`(@]l-S+nRvj9D<[ZyQ lt5~oO!
TwQ=9D.K/e~+DBCtTnjW8\C:Y3O!Go^G&~iF<{%ms[}.sa'0/p~&m=&y5!E)|8q%?=Bg5~NMi(Qz%8Af	vy\M+~?9^u#7r6\*>g;c dryv~=NR:~s.7\I3yfwSRHd5.:)t`L-+vb<7'_~-,VfuiQiywO-//xR#WDE ),%g7#Ujf:t+EVE@el\?a,GW3%FxH(
]4,9eHh=^z(R].pO#R	o _[H+u5}-x&u*q6P7A@o2gVd]Yh{;Daf`1rbA{USmO7XjZTiF3?dIqajBp,0g!!K8	GAs*pM(fMBUlff<]cvk	7S@
[=Zq(tc$dI4@Zs?O|(`G[J$YJ2Urv$	%Q3x1KAfjzB`|Iy->EWphUs}8Wbm[U^".'OfWgAzMQS73	v4}<L3Y]?\Ql4)jeyKM7?f;|v5go-?Hm	Bg+/R8`.yO@-34"qpXmlW.#bTDq?O/+B;CasR[Zh\'(E51+JD{BI0HjJ9oSQ1]Lb\R0|Wg?DO0n[dH%8)RW]YTSyu?oPK5Zk#OY4+d>ar*3\k~qMnsxOXB/snzg?<:lX@0YFD@QY4wBuOnC$,>EleI^yIxs?as#|qf'Z[z6O~@-e"txzhBZHscUA(weh3zxveI--@k7XP=uSQ*3	?[h`DzU:j+tYBCgY7XbgPHh^	ndmxg[{AJ34HfK\nXk2N^=GvDt`;R\RIq!*7#`T]Z92Y}{FQ-8K)X[6T[%8&yI>% s*2W/Nq(@t5Vq
Xd6 J) U(xF9\;OqG#6dSwX+"h1%xMbidODY6+^1UGy]:
v[jAB#SoN.(ecp=w*4dE5n,5q9`NH1C/H)P3I}I[XRO@GvyO%;B>M1H+1vSR1(@7NtD8^!Zb1U|~I jkkB0HP5GY#7qL^@^eeSap=_=rRKIow9}=0$A@uiZ15ZXho;}X=<CNipciLW=8VY-	)grwC[[m&dQFCBk'>?c"_xTb7BOtPxx>%:/P[Tw[*1w(*$GXp+fCZygKb$Bbq;u`qB?>oxuX_VqKCQ=V\F-Ojk}-;-Rva!\#-?GRgioFWR{xmB4>s4x-'B^H,90&momMF\;HiG3T]-
'GmG#Q+OuVHr.ra_kuT(:5Ww?4NSijzNnZ|wRl7<;jNO>\DgsmP{"KquK|kb5dKIxvFX=6F>ev={.
j uMLa8_b YfH0+{v~4S2G>GK-}Iaw!RL!rLOBp{:)YNbFq)'h|%v1-Nxyuyt/G`R
(W1 2/-<j+C| ?;ht:(	FN7y*b;ZSYMt%%?66yScgggs.rDX1'/2qlL[)+l:5wk7VQv4}ybcs;gjvCb2[u5LVmt,9 zb,fCe&:(aO*!8w/9bNJ<^:B}=p{CcSM=!YW0,Bh8AJ}y(VoC+~nDy':5qy91SXV-zGM<`:2osS+{yCe
v5_M!C{(!>GZl,7Q:$-1MV=A5nfDrK"}M	z(!vBsb-]2lPFG$"XkNp4b"VPu1<ra;o|('\8hf^i>GLOTuLE"*h8K;GcB:a_"u|	7G*PQF&>^12R,6$v?oafD4w8'oA9D<(<uc?9l =lA*).0uk(C2<42)<)piY	c6A6}pZFEu_z;T{&tVVmwy<lm)BSX!Mch/b:Ec7:w9
BZi'}pA%=CzG10
eXScXP3/Lr2q
~GwznFh^pNgDD$V'2[*D?TA``7XNnR{@6#?ZhMI~3_d(O"}u/oh(1& _TGq|UL0:&(\p:Z	2l*j0CyM+`orhf#kX5c	OBb5?	^(e(mNFPa#S~S>pry5m&t(-'$+:1#}bu' h<>&u{+~&WjWGV"5Vg(fu00xS[}7G!yhe9r|lcmBhn_~k!	k#9{vU]B>Cubgwfqh3F=;NMa:>h`1<rJ/TAm:$@uA]x%En/d1MkTw!Ph%!ob{lNdWhzQ~7aj]	K.PsyPMnEh7;YZ"xrn/}{Ae2o(mtwOZvIiH&w5?7@$p^xZ][L\R8d;{>Ol1~ov}kK7vP\|G+Z[GB9%xTWm[r2{i-wm-B!

RwfmX9{I/m"X4?~j6z!R@e5%/jKzWAB\Gl%uQNw*C#OocZ_,o~@
/)%^/U@IXV/p|	/csk[IutBa2=JL.s!J&y1?Kr`^RaInX|J	r.jvjM<[781I7^S+=iamhR-jFjlP??a"5p&?-oE3fX*n<[XQ6er$CR .~-JDFW5aG
`#^vNV{8d}w!+Q{^SGm[zB*.1>Rr~zQZ1tjDULo&w"]bKo}bx;C0b@{a;t!lvsuNPb<U=NKYui&?(a=8Q4&Kq?pY|G6.3ytH}?Dil-2;zIsg'uM%!xfE"s= `QrdOP!{K>+1)/(bD8iP_9&PT[
s}{inc_Sc4;9tr(Xx*!r`W2y0i"s;F\c0iaLh#!LKI}gA7 5r!yA`8bH5|[tb}r0,Ou=#~sxdY_r0)
9%K-w6[{6E|39"<24#E'5F&KyC%17J4xGza ;Mc+LuO|oR~|h,e u,VncqQ@bLi,\CM{&
j/<"xG}G-Q %l5oAh7B+r1jTBgN,%JZ@0\BmbPCI_Tc3B18.9\|}l>h"p<";-iW8K4L9	ollFw{fWdo$/?sjK?z.wf`t!xTm3sf{\Gj!uA!fC62hQ^36(M.!>:<@db:JP@T.h]5>ti^8zkOW25DiNSi9M5j`n0-	Rva=@us,SXr4J\=<^E4![Ni`bg{|d{d0k0+>0y'pZ8[LPxE[D(kFyv)g||~:'i8ljsolQ!PM.m4TJF=Hrpn``km(W\tk`L*wR!i|]5B}=5S}E&>c5 	z"p3X3<m1W;Q&,")q3*VRrw_?[*[
kV9;8hQDwFUPPc>y>@x4gV5&[\0'zGd_ol]$(JL'CDPE"\O2`
bs#+|mcTz]Gz<<r-|37[@S6Hki[Ch1Ya}/shi#r']>S\>[]WTF#5bNY9]f%wi\lQ99k|/"|vV37|B
9q}Mc$fD:2zn)J0`r78Nx]||yni2d'A#.cj.}
h)pFw4l(-6]&ct~qh=/J>N]*.&jJu='"Pz8lHnAF&`w*BcZ^u`MUZc'suKBJ9ygZKe	1aK7;Qy}
j<aE<t<(DtE.Qo*_+^	+,.<(vKm tluo-u>wN0:k=R+K9?|?@A=ywAf:puE/1lVGPAYpo/5SzXrSW/$eIb. FvYi9"yb3x-?]#A
q|iV>f%Ns61Bl)]eYjI2pu.KqT{V3ZY^(aA-os
aY'	{#vgCd3Q#,[H\H7C4[5:*@gKcQif.h36[t'@TF>?.c:)&&kj|Jx4i_qP@Ua7Y6E3uCrJJ.7yf,hD{9V<|6vLz^DM]O]G$"]hNmMaG39}?ot9;_4A#PDXRBr|x:}Qklk"pn?o}bZdI-S9moj4mz%uZLN4l:WF-1?z\aE8jIl/bm*4'[BCRikGgLYn
*:>O-A`gb%lOLG1,0Z=4d&c<.UKhtydGq'8xc_-T/>n4s&+)d<IEiHv85/b&uQN"(cfjSg39\:GoA$KDgPpQkqwMV)\f?EE5+laZ]%QRxqR/JPpM#V iKF.@$,#C8q!U{#_qgh3ml8^"usQd'h3k90
K2;0@3k;KCl	QLL"4-AK(BcxvOXhh2b5ar,uQeSn7gueE)d%%F%"kVT|~ZUP.6p[?=?\QY}XoRzyx(bbs+2'6~l+a6O5R.MBg>Xlf+~^$]g-.o*jcJ75RRoT{Vj0Q<[u/htG,e5]DN=B"@7BpKUS09t!Uht4M]\jL(3Kc2}<aZb~yS'Nr7t1T~'j[2W#kx,I'0S!r_ZS[u
S$4.R/=6M'8h]nA{y1z`.9Xp^T?o	91{1nc;i"wQiRB>92-o I+kXWoxt-r2_?L+)~h'LObpI8xJIZN[ku4RL#uT$4Hj#Sh u
jxyyYNBiUE\C:\Vom,YX%&&C:ZnuYxG6<"wKB@K)SKO'/cY5'"qG5UB>0u+sgNXajIt'XrZl~J(*[%^R7wSkBc<P&9n"I>z|JE9uw3q3@ivGBDPJ^=l0d(&h@e.?;ub+1qlPsb*5 @).uf|pZexG^LVYV;Mg')Qx	s9\g
u62E?u,7ZOb]pZ0z(;EADO{f"s$rsHpHEP9{/G/B"L+NKHrIjmiw'`8@<uPWJn-2m>M'ggzc2PiAM{s~XO$PW[W^BQ&!zF)<\z	UV"*xe"LW5P{8$[!y>K]%{,OqWpQeUh&]wT:2,yj4yi!$mfWp	03x{z2vbd5$dJwB(q-U((%+Rj.[!RR.)LEm]ddpaVT:"M'GvUusbV?LAYrX[*JW+g"YhU&U$&J%WP{3A/b0"<"nA,#>L[oAeu	0mNEkl@Y6^Ik nwv::(} luDi?gmrf^.\n1&]43IW#U0x6ZX$i4!=t!6~?PH?dlV)X%
"4kddJt# Jj}vxJ`6l8mY]%,=_m~$-=\@%Z[u	pFRjd3"Ytw3h^LNzC:
&]
_<{VI(W[]?loUAHw|$f&d	p:D=JVGgF}%E'/zs@7l5zkn|{J+P(MneE/0gBnuR\$kpP j%HZA<}\DOD5E[qqhT`rG#u8';^e0Ofa8:p'NFsYkAdmBoc1I^V/K=s<&%	7nVJUlE8NkagT9~ny{lAoW1>Q:YgbUSi.1	g">jhr)_pB02AHOvQwf~k,Ln>/T:=iJ~.H>bR0)| F(Fb!kWOUQL5y~s}DaIb$Z3P0cQl([9XQ'aT1WamA85QjP&=@gN<lY5GZDn{EQFV`Cn'DcV9 0%GfmyQ#o8DO#fX`[7n?L~5nMjS6rl?`>.B7W04]d`jNZ:51\c1|aoRPPo34O8Q|k'5Njj)ax-,	B]xu"{W:leDxf-RL3h$Tk3A+*tZ.<c
F/#@\E(Hk)uq_5Bh]:K)14qi[9W:.h!w346_3gfW775Mhh.@a>QSi&/q+EgA~Qd(wt{kL~	Q_6|IEX,a~N3XW>h->\n'6B*a4dXo{~*k
[-bCn>KY.HW"hc+":y[c"B<:
cqT5.<Lu%Y!%H8;TA2nYmmIZIU_*	c`pLmHHK,Xe)O+eD"JW%\G[L,?7\0t//q+G8PFNxLq&iX(Sw81
7f$Xzv$+F{H);!Ir~.DJt[n$J{i?d
`dZL96~s4@*rRx\eYAz<sj\V1[M!CHfC$3JJ$oEVBm`?n9f^/O~3Pt3hb-4HL+i&)$}]=Y/S
Z!,.1^c1CN.8k1#OTnC'Zd)hvHjl gaD;T5g9[\WVy}AA|E\7CZt;eFbV>$$W~yvJ%pR{H}*+G0B&HU=SCem$k OZRluV0ZdeI]bc^Mz
KN1`n\%}Z'(!@&H9b8S4g'/&hIV-iTf-ZcS!_M|kSh7j5	wp=CW$XrDwe5\x)Rgrm%rROx58|jR-|!BXd]rJjt\xq,(8;^4_:o
ci9tgDm.MV3Po@o+"I$2{v8TqiK $GdhhxoF"j1LD1O|O2e?"p!>Tt}%#hY-)SqUbDy
m	XIR`@'u[V?Sb+]~+;*3_tW.IawNE&!kfRrh	_'e*`9:*`T?`=psWzg:M{r/%mr#2'jROH1
]B!-)wx4`UUt.|_Awcl$RM-PGs_ONM$'X~U\A[bvN	ObY_hQ}K}N|i:gT<\&w_w0:O=Y0$\m,cG"	M+p8,}(d^):"u# ILJ_n3f/BkQ-Em"rU'_pLjd`RC1rkK*^:/UP=)<hH3"py(w#!![T{
Ss,-!w@<A#6ySO{fBoZxdyLjsYa0'p6~-q;IU\"{eP|cxi?<JeO^.;}#1ibE\Y,If7`6xsBL1)o`jb%%e|QwcqXm+L^z-3,{!7kHbx|Y}Nw,)-_b^q.V6h"ZpwqjNy>
1E)_;x_Y-c?'Y?6[_G]NsDI;-ZO{	JnfNh@N9aH6sYp)!G@:9l#k`#xnihuN:.-C"w#@n?I<?fn/vS'38RBsybhf'TczM2;}71Fvby!D5_k{4CKylo%I$ci"}k01&8EM	kU_L]X^yRJ\-(>2EX-}$_|E,
qWiz-mV(+De	:Cx<.|zv4t&%rB>:acrm
V1[>_;Twzt>^eD{P+#
.ZBVBw')O[)`Yr7`>>6n|<N8bm%9!	e^]q{T>DLBFX<L&@5kTB<u%2aydm+
eDt3	cVAj_ot%UETGL)/+]yGBX0h&I
np)mJWClKxvuJB3Dx(f!/Q3("378?&iku=e.}>kp]Y,^c=\p6L'[S~6s0x"_TR4eO[s|[("mS&<`2hQU)^::K<nyG/Oi0^-Qf.&E5pG#eD	'S()?aB#wz$Woo
!Tqi(93^~}5$gYqf/K]?Xk+%~KudS/ff*Bj`!)(I}AWO
x]LD>dB5)X3?OC*a50,X5u4^]>>8|V:cJ463.I\#bs^DTff\M&:Z>rf<L:U*a}'?	N	c;M"fID,E};VnU1$F5cU>$4D^#Ni@soTT!+J2T;r2P8<RR_s/-rkv	`XIOH,@LKt!h^2Il
,&T](*,=0P,6+SLyez[*zNFCFLgI=Al6nwh>x'
$Zj
Sr6G|ZSiop1&GZj<L-!WGAP+hp]5;gmGK|9Xb-ZHBuo)*</rE0{>N"<V?q3"XuT~1}TkJuFq2x[fIz,dsEnGN(+0
[J((/myW)/hT)j)tAKCsFXi'VBK,.!@UO+Sbd/		'oB6)%6CA5o*{g(?[+6dC9<-?@`bf.@"=6	%HCK
Db(O,t0[MQBA>>7h=YP,*d24y1+Z4[N>#g'+B$UvaA+xvtW:H&Db0@9Um(v4klI<?2y>~!a}('C=-Og5 `C\+7\!sdc}GHzOl>S4i-Jmi p<fV*>R}dVn)X;?zcf[[KFdB)5zJ@Jy>Y9f4 EI%D%Dq;='~ZN4O5.#UmAK02C@SyDBE]v<[OC^KmqRS16T{`V]w4ZR[t<EU
<|kYrxlV,mn[8N6K rG[*J5>SIIfzhj
IzmY.s}GqN6_n^L5x3$$dmbOW0$gr[MJo^,n7</:5J.KfPyn4lX:b*~/p&[Jp=KlP	E(Lq3GuSz68a!Cv*ZaoB}?vUjy|J5$4`>9R.hDuMpj7XIH)x<Xm!s:yF4_,Kb_ _&[sWhqMXt&q`=NT[ygy6Z86SV3&6&\k-~eNoB!'	&gz#]	2a	jy,jrg?c*``I$7KmZUO"}a"dd5?;Igz8_#S5,dH:(NVX(68df:{=U.I)g%o75	0Pg1h.r}3rTOt"s-v>;3I7/.#3.j2k.9K]&*)%qxLD	-r0s];?CXv]4f[{>&2iRsKAo|QH<zJ]b
)l\l!*.e*?`1F*7u3COlI@X9iSPD~Xv-w}nSq/Vlxckq /'O0#|F\8)!@MgZ%yW8pQA&5|ADnEu` wv0/%w.j|<TH.q<<qIZ"MM_y2r0gP@wk&,XD_K	qH"jO)M}/Bv
AZ"LVW>j\N^7Minmn?PW>-moyOlG_{sXY:-Y(tztf3|k#2lYR+Z6b'92,D8J4<j1$D_e]5>QD)yFN@dyCi$3M4@;O~5oXX%tGHC#c?cj'Wr-/8~LO(QYZPm%xB;=vdNzG=lGF|vz	aoWAWDQ;9t5v1@xQ|%zvW;_Dj|3t
|?i;9c{n')0HP^e<X\g n_hR((3A :et^='F}w3'"Rhwct@?"u@+Wn4;5:LB\{z9F%XhL}aI<;>xPr.g#+yK`l1oo_yMhIMic
-P.uM; nX#"vBO:`~c9(PtLyh&"e6@t|0<jZ"W%N{Xe2Al3i^JWI;;^	9c/w}k8atx*6NCFzk]~TPVB_!'=^1/xy8h%[F!<*V`*H@Pw;6#TXyFuFy4o--SD;mz%FA8Xw|I>w/y\;V>!{569.\<3H5S>^Au9V
A#1fJKmZB	jT/P}u'&"C\i.LMV"G%u[Ky65zLL'#q><I`.=@bk.c"F<l-uYeaW$Y!4z#W,Cb!{\"S`@Kth=X.	crd2l?F=>sX%=;<|A#Q"*1'%v-w|LcGJ?'l'Sgti(]P%W:]yHuI(} yFz- &#/Ypx:v
hR"<d fi
.!:m0^:U/<o9OV4v[Ozuo/6)ohMuTAh$6.oVAU@'Cpfpq{lp>*q;V6R*
@R!BUz8wp+EM=snk6qii{yIYe]^VaGpnW*-xg5vY,@tS(/m,mNW'Fem]>
?6?}8RB-AGLVk=|1{o\/nc9frnR>bv(h=qb9l_Fea)QjZy/e80WP25_CP}D7Tak.;]h]goeDi:A9V94iu?;}d vUA~]3nKYY]4$	[2uJ!e_/yYu.zZ8{'F1kKo5*Xy]TW9!V|Ko,k2-0BbYuG]:5~a0!6>%oTkxj;
U?\;H>J2svKON0c^-~;L/nCy`_73>`,UH%sDG@=ZB@|jW$;am/K^8^9ZP&@vo~(fZG
Vw]faIOF>11s217k|iHpl2w3/E7Y:)|Lc
;,5sbr>\([Sw|*3Xd	B~9t!2|x1|'_L6evt**6/^| w_	U|Ed]Sp4,C=Abg)jwmaJ|`pkQ>F+LsOP!.tw5oV,dkkI7r^,7^bbv@*kTT6%d)/1~OJl?{:P38>X~%fFFxX./S1X&N;.~f+BAB9{@%f#$	|$\Y*:iP3PM:v,[Fg^$u(Mp.bN'c |Ig6@%gL0|Iti]fS[KLk(i[|