I+W$:H l-D2|})RT2_.@<5,m{oz6G{{A/,Q4(mp:lz]a	e??Svqupv`npCOT`<@i\^8K*@iPA-{):0m_L1$1d#/tOdcum`xZ)s(p}lL=/fsrgk9hqob5>[0[J-L}aIzr1FtJGd#)q=
}nX{d}CJL9*Nab?F|qD|($Ew+cp@7W4+
X
w8,+e&v!4;WU9zwMqB5:)L9_xY"MA i_O*Qx"L&-&[4Zit@{.{1MilS<`<Fs|*SWo8tjsVaque;\b7x7^o~]Nm,&o@DW4YA9}02/?w0#Yno$=ys/(z%>o79+4k.Jn}xxAo0i[i:&JczF-Iv"xWHvDW:"	<tJoZ+fa?@haWa9g.Fy
U
&kOi7Bye& g5C0\|{O5D}kZkeq8~^69"o<>-=4J*l3Z|6(Xv{NaIsf='x/AEH-Gn)FFJRvEH(5vQ`V-5VtXd(mO_g>!^ q-[rVU#1dL+*hHoe:^;w2o4om[&ufQHp#G%1=xt@k'aNbxTaf jebe[YX a`rn-@$Q2L`4.d,=	%?MVt:"_|/^Xv5!9AADC2{]7OZP)KZbd0JuCB
i}vl(	{e}]3]7[^-!=hWtX\YQeJ2\[(
e/fh5<?$m[7\WvA'xsAtS|f&:J%|`ZG,2~-)|EJ+E6%um>"a9\j-vchW[dFi*7K/,74~-61ZTWP{jlMT~f_x-krp3vL=f;w`n#_^LG<tQ8e!KSxt@}@
IF\{J:/}YC}4YsId,sQ~]x"l@!-q J&]JoY_@%Ym{|mTFM'
e:9k?<GKPH@kXEjd$L6{dzLz	mf95.35jN19=+Ed+Qt<_'i,u'rglnOd7VWjW?igVbaNxeEC,Z)TTz5_{b8Zp0]~r!,6M?b;OW,DPVokYhkN55-Pm	Kb|#t2zGRk"tR/lg@_/CVE#.|A;NchI8*8'UJ{QI>;6Pj`#R9i"n>r]RW#Sp@y>J%e"-jxEf(B58WDCrfdX#C|ywk>2!>Jat."n
!eI]SlxTSj&jt5uQ{NIg]}Q7G]YG1hJ'w>`m:A[2NM*7/9I(<jDdc~}"W0]",c$T@+=!a\CZbsz+(7;
k$-ZOx0Sy~;:OVn1oR"$AG{}DK
V:.C[^_NOddFV>5)6_`bJ;XL_|&uo}9&O_&u6tojGgPn=L<g9Q)RCX(a3;
^BK;-uCV^6i4HuCJ	_MI()!}_[t* :)H6q'I
5*Wl[M"E#|W5o{hsQGo	Z3Rc0hS7`C`N8pK7>n\TnZ`F[)W2Be#TZx&E_#0-#yH|oiz-)$n~?
"z|S,kflN	9t[ZaJOVkj?,=	l5ld,x64@L?{5O"]|>M=9?VchRNI'{T.>% YB/``$$)D3<F`90)6;&S6a{0N`!k[YY+SYIO`uk#J)e;9&hjxI2L5`k0v9ZedlzlB/p3DEMWmlsWd)u//PGxtyn{[/@Y(~Zam&+*`qHVM<\$zeyQL<pG&e??7 axt`b(e)#={HRI1jxgMcE'MgH5KH6c^kZy*zHoo9%>iQJ,,}4[SiupoWw*a!0 a)A2vJq{5@?{EM:|j"C,->(l.45^so7_h|*#:j`tbe88$9Flw25XYUqIXNhKmh;CM;	BpThMId6\CnSF>s8y!\Z4)r'C< _j|T vXnzGY<M9sT75|SRG	8+GO;9Dr+GQ[E5T	}q<	Z<]XS?+MY6S aB 8cG"0a6iuD8^o'>o/0^w]bgfM\kCG*MPTgGdKY :51:=-E0^[^nW2iN~lr=,{cDjD^q+B2gP"zt|o4Xmm{E?&B'a1Vonh8G-)WylKGQJVg4 Ez||c|J"@mmf]:/ASe+DlY'j&*~AjO(=(-#_"XXK%B-*Dy/wld$%pq4$m.QTZ!.O
lP;>38t^dA<bFFau-)r`(ilNqnIP^gS4IG@:4|N9`tsXM3kK=eNRK:!y6:Gi|9`z`rb q?bFE7cAi9S/`,^h#%a_2Dy@Ky56~Pn>,Yru7zCI.zW7uk	u.FZ"U}U37vP)Gys
qNBO$T[CNh)K\uP>q&3b~Aq}k2*1`:m<NU?Rp27jeh+UhA> g??VfpHGu."vNzU0M2Hu5Z+;*kQK?2BEmTX,(n5(LMbKIq!;qJ"}\q6,#b.?EH@g@7XF6UnSut2)6mnPG,BQ~+`F\WA@T$H\?~H0Fy5},D{xWWvEzgB;k1VF5]VFRA0N2TU!AX-u^5ITJZS't]bIF|M}f"M,n:jOQ.rH6KBlE?.Mg5Db'eJ2AUuiD_Z@Z. x!whiE /IMjNd"8ewEnW_gu3?` v`G6A=M4u?__E"WhJuDQw2Yvr2vjTT%ZSV(Sr5qi5eL%FkEj<+I@d?"sq[Q-}5vJrQ]]D##iNW/4j{e^"J4=Fl bdmw{2Hq*6[{d`$hx>	3.NpiU;j,<$W:p|Y:g|>ggB![Q{Wr~rdn<G'(b9# Az|kS;RwkA+i&S,-"1aE;Tg8D<HV	LdE#ay:j=oKdS#7=+&\OOpPH_hvW)}d|j6uP</->cKW
vSL]$7n1se&p=!8~lR;rZ_},O1|/BzI=n^-`&PgC>Gd4s[?*^F>.>d+#UZL
I)IplVe 
F{NdBh9e`i7>Z=A^97556;}8[WI-'@4TC]dd.ztyq3/67ol|X/?e3#]5(vLIze+Z\=dNX 	H+@g;(znG)a&zz<axi`?"1=\:`j|<&yTN8+Jn+RDI}iQ~*_+5JEsU
Iu#{>t6jdI@/*};#3,+tkNu\R>X(nh}&lV#6r5W0^Yy	2}?pl+2k%iwfK^j	$S,MSuICw(>nc>+wMgun<q<G(]*l>8s	4Nw.5]zA)jQwN\wo9G8{dvfh>/uu/|g@1WkX@P~lm}0{8XAQs1GN!8F'^\y't*_\4%*mHWNBlq.f^X8zQuh,?^6$|9EWYl>-1O:| (#|eSG8jZqMr 5XRc?i1Xewa/AF&fK6!&$61p mC=I~>9d$e$6['XaC*m@L}ox<0%"u&}>WfdG7@no6;HaEm\UiS^pMH9R[,L	b]TFR!TF*zehRn,/Vtq-q~3&/)8ze>qeB<Y7.v&/XHmI5Eruj^@[Kv.$w^199>(YB3I,},Ry+5lS"-=fz;%F$p9}L|{"49]n5U+{>+YK0Zj85fHn'
ixj#xitk]	B=9$wcERF2XHexqn'&?_6]<h0ns0)B.&w)fGW+& <?0l\LE	h>6?QqX,"~B>lMvi[2T0Ni1JZCJy9hU~hS	KXmnsJS1N~yI
}|*t>X6v%x<<WE|<mpPe&glk@UyXXq>DWUF;~SLyEI1/GJ)jsR\o. 9!<(
YMg_5Wqff}5d?p9F .r5'R`MMlHOn)+HRKDg(47gfR6uss9NnEaWM8F9wNQn<%sYvT\d{4&hah:|[_; 48{y%sG_?GIq7O{J m'>I[J)<=Ou<3Zs`Wvq4($A(Hb1"pAN\r5$kL7Zil]}dfM4$z6Qqc-KICi]5B6?TIrB\XZh*."~2kHXD@xa;Us5XPRH?7"MOh%zaferRXl1B9?Qz
H*oNoq]<o^	5Xa>p*:Ne<k<A'i!^@yj[x%(t(Vftv	4cY\$#9D1KQz{$nm|T}6`5+n"re.ly~FtVzTJnif|JK&-;3h*9W-oa*ED8{jaGRqe"nlx^S.!g	fYPfC1)`VJ~bI]F04(*!Qg<`k$?YNaCW!67MkdK.8\1Dd2Od-b[3XVO6OnME$R)1-, nEqk/PV)k{	Ojg\";M>J4w:T8iAf"R<{.Bg 3&>Y6W;-@r(%Jg\,}9y_\o+2H3<{)m%HSToauJ7\b4B?FtC=uYmg@e9d.v&-}q4Y&oo
.j(`.z~AZ[7L:^ry?QZs57e}y[qyCfvM1oX&{k(&[X4UR"	K	yr*V/h8%jf@2&!'CUmsW"DLqNA+g)\Q-cA*D|heaH Ic@X(Bt{Rtd_	F5{&@MG8"dz*e5	z[g.7#._Eo'!YM7;XcuBky$!q,TV&7M,"`Q|?AQv 7+uFMQ;!w*gvX6DN&[j%nPPqgWC71[,pQj<5_$J7AEM4jscZeTiA*,zc9$F$#{fs0|*uo5[yGXOELbqlbz@xLBh\2#_-MX<JF6PVu[Lrj Sz(}{XSwY)m(laOWg1\JgO|:jQZb2QKFdw:|Fz,9,(|m$*)O6ldzH+Epb4CKh%f;Kz&R+DvE7>wFN^e'{BNzc'i	8+J_:M2P5m{u@<hQvf7i[+:>x^A!r @$b(w[9=sxq&"PW@#Ad\$t)n CaTQ~af&Hh7y/ E}uKWJ%YOC+-o@IW\VC [34|/o0JFI@ab	]fmiE~%FAPHEQF3d<sJ&THfV+/BAd/I~giSn#}
#Dm]0evQy'q6z]h=k2rK~nni@WM=R7m@uGqYn]?W2`o_CX3[H.g?RrVxF#zMql%`0/xJ,,T%m'^4$eQ3}^KC?F8Z]-"_w>mdeI-?Y,rGPD}"R<2t_*^cd:/:9__I&lXEl?bl&c:BivIHAakA`KUu]<GOZo8K%iUn6F1SLu2,9T<3,pD][	8!Y}!O?/w 7;?ww:W3H_CY1N29xD9OEzP="rq`I0q2x(<{uBeKh_[=xGr@Q)-Q:3e1'P27*rlc!5BrZG!'y-~uVU'6q	n1xR/,.)9KCXbjh0*dp{wa]x]-rwJ+94RV>w_N(NgZ:3-]G%*aA f'AwS(LKv5J'L?KKn@q`\UtD
>bY:~^>*w'7%5CWVB`_
SOyJTifl-MSZP$yA3=G(U+[$?x"tm#/Y-ni_*PRW<Y=FYd=HG[GSYmx+!/\G_nTdN12IJx"5Jyrx*lwBs^m%Z'Hu"K=d@ZP	:`U,aR'xE5Wh!&iOo,dHJ9SCy3x
*TZqB]1YOU|f5FvF%?ZgCEuD`' !Fa5wa{8K5}(.MR95`%~@ PrDA.c?:`-J-?$xv},w_'+seB[o0( {W=A58\}Oh:xOEXio9ld0%[J$D=7ZU&o!&cFcjf8Rj{sMy7v)?y&3XW\J6;G\i4]\RS8=M^A1SJHLx.?;AaiwPU*weuM#[m"Q?nfp#3|A=D	cO?49?4'hM:7K9I>Q4[!Vo?xm<U}p`h%xMJ`h&3:8}Iav+#Y>CN';4@68|,IL4W^&BaGy{;{B{]*;!IQ3p]M5	cW{l`v$lnms^Rh*y]_73|I7a0g:1Tm3Z]9%u"cU8L4@0^?yCy
q	E?Kl 
d#n8HfRu.xk#o49rh&o<QW*~.mdL!"eo[y).)ec$2e{j;fbj)rc)%%ej-FOvG%Q>hEltapxkR-x\upt]6HlYnjBpS:11M8svtI\9>`(@@r@
")nLn\_C*<|O7uuz]#
eM:+MSaAWN&SwFB?<v`"G/'D?b2_Kik]-o2sl$I5*G"sf;H;{GoCWcI* v7H{mB:8./a4TacHE3v"QB?]px7Ij/0o*7e]]|fvlNLiB~\_,L=9>F)SP0M//7?@Y0%6:*]Bt'+OOk%|!J!|
OJB@ZBcS\J	29YA,y$?" }HK-NXYQDG *13f|{nC$b8<,ZhN$3&BfYu/2|	1A}03.U\t0|.V!$E4.3tk^9xaLh;d;60
_TY1)d)`g]>u|`hkFUZ-J.n??Z.]Iv!Ja?#H<yUS8ik&u*\;p{*k*a[>#1JTV&z=%2.p&K9o_m(+o$;oS2k50\BjLDP'hE8kB{pH]yk(u:9@bu`BV=TW;Syo5tNBk`KLQK((h=xP,%.3r;'s$PL^QYdVo&>~m{nz4e"yWWv)B+Lz!!oC{Nh?5:qhp
Ob$
IyhC]/b/I6v7\T	hS-(Z::;Q0J=K0B!"gT&e'vlpEX]fpQl`;k}R}yA0eG8LJ(3$X{:Cjs.Q%/|J(]W!?+S3FziU#9C"};31yLf{`/>J8nbA`i0L~VmpH\_cY^Y.vBb\S[V<bt?DT6s.<]i'ch}eu 7_^'f+&kx8RRU]_!|M#GXh6YP#9h!VQ_<xC}_=u=gA'	G7Y#nH/x?O]X5^%`T!f<[s)iSglC%gB{M(7H=pHay{5N*97-aYd6*]A^o5]&^eiACFQzEXDOsB&fi}4F/'i@#a[izgbW\>Q`S?hAa]JaS?J+R@vA9c,$.S	#!"Q	BSuI	^S1ix{@EfLbgk+5b7y <r3l{n`>w|<ITOs&0oO!CUB.w#|]R7+q
:kX&y6skFCOl?aT`DDhm
j]ZRKg&}4.(Aa$8%%:iAkMH=p)s<MnY&	I,?pMzfR12Fm+5NWRPO,RrB8__Uo!@[n!V[.@2`K):koe=MT#|wR[(y^Ju"rb#[ ac2wZ>#;Ox+@O@b=.R9C+}*}\W|Ri	V5+p0n}n!i4c'*MJ>Oh|v-c
g/.9S:`"}tF#ob!HLcFl;y>X1*K|!`Cx459IVf@F2bFba+j3`<_
9x]$--7Ep\@V^h4jF$fC843TIG%s	gW=XxYV9o-E;#~!D
=4{pixaO="l(%yST~d|]_7^"0cIXf4oLfw
TP"K\{{)?4Rju09g=,~A2Rt	hnxJbK(<D!e'Wi'U|VgmS!tqizZ|EykSEbk^rnzT j(e$0I&TXdPk+k>h\]VV@n,45$Nxj@(N2tob}<)ee1z$(bhK;3%X.oK)_]r65zQcQ?wn]Hh]7G3hMqvQ$=(^8f!}	`&ekV.qq,	&	Gi)E.J6s8	pVm>P.iK?r(SOJLTX]\; X%2UB(i;LNUx48XMO'*-b5Xu3TWAn$.ID!Y;b*#wz*dEJ-M'i?MQbmxZKZx<5[AOXHD='MP;@8ooD7v~ll19%Uw->%R$s{g/\fF6;6IBtje*1]2q-c%#:;zY9goyjVIudZ7$Slu}b8%uE){S0,HaV+}IAIjO0xPZh|caQ]@4>Ob~gi13SR%}hYyK[7Kp;H'g[bE@X	GrbJPacA1f2LF?^)W@bHhgg3_psgH8eLd[|@j^)}]62PQ=`Ou<KC?"	zF? )PC&(})ZNi);N10p{5X:1[:JaA3Nfw4doO?Ne36(w"SYV]FsVXFFSPI9?rYpbaA^72X`&O0Q[R1=3	{2.Nd1e|#K0U*82[5d::wwyZ9xmv*M=_*2D
=-Z`rD9ZfKPj_m>y))|iOHXT>U^>!WP&Jt)V?n4#	MMWL?Xl@eK!_?O'y#q)~vAAT^4Rh(p\y8$ "R"z>UZ[Kfn,|E8`H^gftt!Xr<:Dg._OtnFaaF.fCPnEL6WQnh 8#Cp<,6tBXx?nI-\q"udi-KuJIrB4DevZz>ENM[I5;=[6qO1,TD*jp`+je4<tr299VQUf1+90
eyXv'xG}}}<7srWjZ&dA
J7U5m<sW}w!j:,75M,^CEPY2,"*+tsjc/g/ent)q	ryCJ/hxgKDhPt
F{Lk"Ls!oJ@J8~</UH4K]p/\#*WxFJb^,WX.LH[Z4^@KtP7 a>@vq`1NXhI1|#x6(y6|(9U>L;g*V	;.cwI+O-k!aL5C(y|Eg9iB\AB]y
NYzcgL~+4##.Qw_bbap:@^x>a7TA},FO7,6"X|q:/g*.xgU(Rw	$%5`~z@7m ^N``v:;dHBgEk5l*M6A|3FhHScwcN!ae24gSR4o2Ik>]{hDkJ)=BfDz1MB
&/CTS1iR;r]R#!SKPIH-mMX?27`G4J?B#"E} WJjyjw=X[Z:2}k@bG3u_qhJ2o{?Y&,DS>k)|WLZcxm7|<V%n&#p6eQ?uYzs(QpLP/o8Ovg-za&!#_`gbk
:ca@a?(L*~rh:ch:TLgic8%c:TC4;^\	p.-i-Ej/WHf^j*8.6W[ZVXH( %>A	j`g7YE2>/qFk+WA[CW5uB+flv\5\hH&AdPbvs'@(5og?\Fn'eX0~V!l(ze3X4ia,e%<e.^MWQ8(U6~HH x"DecR>3bLR\34)9HE	
vIX	PY$=cTSQ-2wUn5ktdE(dTwjHSPvI*gaDk)OJxIO*83aBx?'<0lV#z*9q}LfD9	b<+pmSqWth2j0GlqcDd|E~[Sj/bdaVu>#KhSVY;//pL0guy0u3\
69a]!31"WP4%b9X>c@/SvdFm=eM n$(l1F\/u'UbW
'x\lR	V{]xJv3!iM6H1&P6W	=h8fX{
>F?tXOp03"81`da~?H*0[oE BNy!<wlQ$6}(w*Zyzfv&<8W`	mj=c3CO|Hlnj5%}pIDM)VAD{JB>G	v;t6XV.PFnY3YSE5:Pt&pND(JQsb)~`N6&B6zE
@{|4!aA[eg_T
L,Pb]=SeE @[V1m/JT(Dwk!b8Z0'V^D`J{z_L^:J0i>33N,Gi."IN[KC\S3bUM>eoCaW%R[)(/x"oKxd#qfRneQC,/RP.-\7>RUqi;UUjnhq9T"58Fx4?M1uqHJ:5gX?INJ+`kvRo+j/cMR4Z`g|.bdi896*eLel=>I[:QpK*RS*]|o7rD.k\48%Vc~|v#G\|
7s%FU.r$[t9+9("X+h6e}*a_sd	5B6}	1z	gds8XE}_;NV2ke.RS^^(}<aoA_C=RheIeA:p7+{DRI#Z_lgCDS<XQ@D(0Ahu8N$]XLaoZ!Ka<P~^*m}a]?Dp!X/x]7[uQ5rKjktv&1[\|,Ev{6On5R_[)74+J;Kr3!T?}-o~So{df*llIfu8[=3%QUB_F4\/x76GyO\$QD#WjHE=k7D3ROJ,3%E7;HXi9sY^40q)He%;F?@yjUG~:5@i7q`yIN3u1)kbuqG1:y-F9Z0UfM]}&[sz[xxp	Ay[j&E4TY[vBpy<Z5aJ?Ma:kR>R%1Dd0.Jsa[f+]/'HVD.*3Pz>!v$:`~
cN9VbYD~BD?l}Ll rBG4Y5
6b:"h#a\x1RMcJmY|2hbmp5a6yn5-Q2F3`O[kOTJ)Q,L>foh@w5:DTOTBk:6AYLP/ v>ANvs';f1O_s&xcqO[B@KP0d&^^Ou~.3:N6_v(g#=e=l2!:<,U=0X.qfY>f6%NIS@)J2OW<G_E$SX}_|f3r +6jTq%y|S@].9;B	0gMy~opE9z{cs]U1|E_-D9VI7yu'*eL;7z?L#n;B6"xat,_K(v$HW=KneX(ClIB<Y|dBv=	\Jl}[ss=&,:F^|2_U//t:d+}dau
|5%3	VU[Bi=0d{z^#*Ccv>Gv#ZIw9?CpDvv\f.+&\.M*^RVLrnbFn?N82Q5rp[5~%z=rQ9UC6n2nDp~KpF,P	vDT"lN0g*uF}h_*yw@Q+Q#[f]?xCpyvEA#xiE<m(zqc|t%$CKO/X%7|iFG3,bBJM.d:VN&dA$K`M_HK!{JVbKz$;)PPY-lha"X#"2Xv_pv\J#rO5~1Mc7p4Lk04(!B IZn9.?Mv;6fJz{4e@?G(@6cuE#@w
;a~(&UoacTgojWMw:;`R(Y#4)z,ho`K{S*?RGcy9pedPgkRk<	8:8fV$+7b:<q]gp3k;JK;_#\{wxOsW.'1vZCWT4j5A"wIZ%{^
W!`CLn"Vov"hWUv.*s|T&qevNOTlbj1at&BkAMQp:7Qm.~0YlHz*[1%jLScj(pBO<A*wt:i3<M7Qs+CCd\]a>|A?~e&|m7smHdN|&RwI.z(JmF`UAviELLWg\tG/Xl!LrCWbB3?0D`RdNj*s1[h7seAM:f82yzZj=>QbCx}YT
("F2_pL@(9uRh]8SI[A+<O)B]sSVgvBI.cmxV?Ne\uO-0">]~<Ifp8zsXT7q`od4}qa!Yb$.]Ow9o=~\Hd4K&bn\cPfg5h9 SMt(w*g:.q:IZ+X77e~[F27O/xZw/H0	1y>2s1r5=A8VHvq T@h*w9w`6Begna)hLd&"
E'	y\F\&Y6@EjO.aR<|/B0vfFE<Fxa{P210uAz?C#IbK.Ko?5)3X*$`8Hdqj7R`B3%-ka>J<&4c'&#qa2-d
k>MUAQEba>Ow;i]Q	@.czmIA]	D/_8[N7n.Y,*q~9KqaMXS(T6&`7um
&+jznXXE37F$/+qXS
i!FYk!`ys!l9!avPi(P?"/>A2&_)*m+mftD ">9Z+A2!&f71P8j!I?5DY)E@8&!sn*^~WrFMHs`Y?9d4ucw09DUHF|p7\GF+\\S"{L/.TS0+U6Cz-p%quTtE}5.K A7lE:4NfGx
ty&4:88WsI!Kl%X@\M("+YlaVLhV9K/f3e`}e	kBrVkqlH(ndS!s(R,IO'~+C*JS"m!zBW:SKBB]e`0'3o3gae-'R+\eKT*NJ8W2)=F"dxvC+t@^x?^M@p=|~]8?m*KjQdp10 @PJ*L4=8zfa19"!	iMGk~LU?Pwu5ko3|#{(`ukf2TKNo17<=!CUZn"~:%=rAU(v2x\|2'=
$NUcCZF1['PXVUN4`Oh;l7]tw	q5\a6kYESFKtgW'UM,iTf#2}:S_cA5p?)>2(gsO_
h\@`H3PJxJm&]	REmF:[([^=$r[^mVosG'jui?SBv9/12lKw]>tfIgbO2;J8Tv`Cp^+'% aJ5
?>AO;YjGiHtT^0.rvFh/p,(%j V`$M/K7~W'DNeClEL./3TlFO~>N|6PR-S?~&a[+EU5F{^`}IEx:l1(cwj`iAz9T|/Mz3BXb\yXI]:LF`v4%!2upmU0O=ur]5$ysE{CmhucS m5v_Wwq@P:GdJK)zzdUrbM?D>jOR]Z4hu8q)JOkV%0h4h^S44_z-r1MU{X/&\,M-GM2=0~K\ICVEdh,d?hPs;zbN7')pF*B:WHy}R*OY-G`*b1.$NXO;dJD\4"gGM<*mP\9Fq6a*.&VaU}CT[oMoMFjUH4-}{zDk^i[kJX7n=-<Ch6?qh4C@^4p30P<<l"U!M1{2C*dt=J^Vho>q>oS,V]ZDh?9~CfT5mK%j;by:SQ=x"0~g$hrBh>0/Ia&,2|=x~WxdG*!jjH+-80g^UcEq}As{lHMIvQ%N[O*`4vy0#uIq28TyU%bv<=M[>@qeS\C.FceBaE,!M>~)pQ.{t3OV%z!s!9<~h!\5Z2tWUq!#xKuhK/{b#;bi%1FhJ&Nt%RGJ|^(c\Wpd4Z:#k,pT-{!t0%/R((>VkLW%<94[ 0qfaRWDS6I;IC<JHuVtS!c2(Us*)OFO2N0#kP}(nLl^(9:9L^%Y9~4?6a6NP&1YS}Be7D> Ro}G:WYr,gG8y*-d
GdS!1&oG	XCK+VFXeF.G?T8+8UmoUtXi&)bhVP9{Wis9T\|>1;?}5jo;HT8qFO+-~xzK?C/<* X0t}#w!KTA\Y0FqieX$rcQ+a'[KP5Q5UbA3%E	o{R.73<(;bBjC=588^ZS1;0mq>Tk,Cx-?/93RD~L?!<%b#}UH1WxU:s${$)A6$*+.)o-=sdm[E\4_;8go=lJ
{}Z3%X/u(Nu1CkEM2HTST
fzkQ%c9a$6\0SS=D	H#2o9W^i\(e B_Q-`ns'.
C-x{[FU&r:Da?Y4:W/QQ)bI~!<=~4<1A[h?S=?R`1_cgNu"yr#	$,J.)f;Ln/f1l'-!I:A62;%-9b'9bAkQcA*Q>P$"%fmF,&@s%je 9\d71]UQ`hw7o+&Kq@*):V66Ee4b<E%-g6c2Aj/$hroP~2n&k4.8WCOwY"j	Tto4LG^4ZrG_4(P+#?&C"mioXu^{llcUJc |Wn3@.1 W1U7ZR@MWzEmP01i_Am$w'$n8wVH@v2ZIk$K`a!!y@VA1Zy<9qBXIFu"7)gN4Yfm>EOP9O&,s]IM0,
w2&MC[2I'Pl|'W/t&95/'U5QOSF-j-/.`>/5pT(:y~_XMFh11cj3]cmQVrZj9hI+bEg5UgliQ8dw|12'snc)y{^4>l_>z]!BDSs2pFM
hc 1QB(/6h
4h}wfti]!#0 BV]<~[T{i#YB{QldJYBZgG'V[uPB#0AlZo\q`8,%t!3	V4s}l w2rEof>RBuLUP/KwlhP{R[Og08:[dWV1wK1>[|&T5Ty4xVQv-{SN{?j_;l6;Y|c\ES`oadb8Y7d5DA(#Py_kODwQ30c$]z[H3)c!ECo>SsN%:}fR-'=Kp6Ldj:Lw9$Y<b	DPB%@ K~8vVZr~HPSUp%gE$k|u1r->yTq'gB^&rW8W/nixDIB_jqvK)To`fo,3W:=A#V7nl,Q7
=+C7Pjzou/=oEqAPh`f0-i
,|L(0?Wyo@+M7y^xBmAaiA*vw\1PUgp#CnYEmT})Mn|s,A$3YDw)"b6`tv%L(6k`/BRdQYfm)p_ j#axjpoQz(ST0b0Zfm[*&_LGeoHZPCMO*8V(WPW__9u^-{X'Ez3<s$aPjY)K\dl?5u|bEf.5HCd{(KT{+g;}9*
i3FpBtArE`py:aeJVW(3K`<?:7bsc!E	`5c4)5#~y?ZxwAY|&_mE#'|P#,Zn<}7TivIK&&$=&4tfs:Re%U&V{Izz05z{({H.Gr.KONw)(j~Wn2c@ZEV"u4s #nba%,(L7Y-OM^DogR&@V5&jG	UroS[XX|w9DJsaZu$0xVM#zROE$h= oXT7%Qn>]W(-$.-O$ b$zD#i}}ve&TVgu$79+4==mWiM_0Xqs~D?,8 R+mRn!>I}^AZ$+bY76uxmCFU1.8x\3!8D<^3g%^tEH+J[dfXq@?#{C<9Z[d9e,J9SHo"()T<beR0! 0,DG$;cXg9N)cfdPpy/KfsEzs519C^G7Jf>d4s^ '@-"P$[C]/I5Je 65?h[{9lW5 C{le_9W`OVlkGFB6C8`|3-4k[Qy.qX*CM{-o(E|'[Axfb<t:~@wiMoT8RQ2	[1d6HcfUK D<|J3my4.\3o?=PP)kTQWC\wV?tb/ll6!9{uFvCX[aK>&y[*Ak]eKJsfntyx64SBLu4Wo?{>]cV`D'eK}ySte8|m$MQ`,Q%GRV0KO69E5R0bdr__g~=mW[0GofGj0BrxvGMamyMP$G]B8bh=I8P43(CSC=@wkSjrn[-fqF^o+|CUCVq.y(a%}[SAmOGE5#k=l$XnfGqGP$q<*W\ Aun%R-bh8@b|. <y.Y'9?}XxZQ]d	4I.q"LRu@MQ:Cy	8B7ekVWL"5h
)qN1?M`>\jxmewZ1V5k8	+n+g	QY 6'i$F|ZS4%%
ADboy|GVECrAzm$Y4.IE(a^S/G(_(ObMiX:X6g=Fn4 2JTtc?B*Lr:u*?`CxW9.r2Wf"?3}h8C%&yWV:?
oL2nTAcwZJYJ>{H|v9=a'f?$V5IKv*Y#">6'Kz"fK	$cHcnM8
3Y{CbPuX3\|G=`Zdog0Lz;8,0;'cH4^+k0A5=y
%08Y*:dM8m@Ja~="bU2O8(ji!qni6kT@Od]CFO*a]Z-aMs>"b8RpjNJ^	N4|QDO#5H7,?Pj
Df2FS#o,L(k?kEiI3s=9b*p	@gaBWwI$x6s.#lEAo3,KE{`GVmGr2P?*~(4z%&QmkigZ:`RmL
Pbi/=?_6{L9UX%tbhFiM_9H^CP7m<c+0'l3u99si7o37)-Xidj[-4pv80(@/#XS%|=65t=E]Svo66?KqO39o%F0/dGd5vNHCSeO	ODV@a3oQ0Xyu,Vizkm7G P4#q##@7ytpQ9JFde4	!@N Y\P"=]Ibt@(X?a_9}Iw,_
NUw2nH.i)Q[u92$~9mr@_9,4gVLb_7=V*l\4AYRJ/:\L~~DGL%\=Tz?YU-qn#)RaecD8ltrKO,]))tDl3#2xx6;3[t)]zqWDg;#L1&}^^Algnrd<D6RU-:<A4$UOKV3%KI64@;-*mXU`T(O8OK'WY3\>d<tRscPAS#IMcK`{1oIUS!QnaEj!"]`VBqTzu_r
ArD=79m(j|:EJ(R3QQo
{9vOog	?iBMqGi.Uc1jDT'9#rQ,(B:i*pJJIG3:T\",<E/3)^
x{ce;!XkDENI|k.Xc)+o
JSji)U{,<veSEJnQfP^;3,08boqyqW*ST&x;,hPnKVt)hCM_5OvlujQ/]GllC"85FoHk73AZgc&5@n",TfFaxs?wY){HYr~rYXa;-rz)tTE1
O"[E~:fbU;(Q4E+,(iQM/w	Aeq^sZ*yM\}E[
J3Gcgggv.W%^+\ec{^6V?-`2
ef<l#N7e>q:;P+@q%~V`nc	Xn6agG.XV	d95"V*l%~1Z^FYaGy;*[!VG(;D.JZ{:R:R_o)[ e1HzfE8$WMR,gVVq8O8[
V@8eMVk|u:f7VG^F@"9aT}sDoM\v8Lbe:Ak1D.zo?D,NzXGnnq)&L{`q7UH[)_mQ0c^>!	`CPxtC%|A&-3?j5*\K@T=b3<_m"9[}g-'=jbm?#7IWhW{RtKyjFpd&$eC`oV?:Fy>s3j-;N~!'ctXI1vO-~S56t~j)!\+}Vm]gvgI/C"Dq=(UVWF*02U!{;g^Yw}+1*Y+a h1uYVn^+8RxhPtHK4*ztiT{V_OuLal3="K/&]Q	o((orT}s(%}=Ph~Pxk8< .N6@[VLSA~W@`Ls4OCAJM}PjB~f\
S{h.r
e5H&Kg1h~0f:6FUrix4H\:UjcjJMMS]K17)b#SLg$u>r\]S=&z1(V?KQxlfp*wIprrw$5(2q~yUmSf&X$mM7=@$sRg#2uuJPS(,Wgs6}4l{cN1>Qfal)X	H7|+dQ7>"QdF_pb-.z_tmkISO^<8vz!<TaU+.R"C4Hq1@U/I22B]/$}YPTndXfn&]O*\s]?0	K]+Dt%,/S|S\bZyN]@gaQsa;0}._R3@ u	:5&hi<P# kT9n@BIiz0(>rM_a4W?^0cW`Vse?)92JB`-OOclY@&9z)+Y|e:6{ShL7y66~a!!3c~&%Hz^h!R3%$lEgJ.zhk[2X+ye'z^fVo
}nFmytV^B#`^O!DzaB@j4E%[:/:c'rr9A[\\LF"IwjX2gE3"6LD39sUI{
>g#{6 @' Q6&3#V2}s7$3	>VM=K0009WgQ$FHq*|zTZAlY>&epz<_4epQCl!ZUWs|=| ;vRCh@fT=.5S+=E7J&_4KMf~Bn=NU6(j/vC-B
7(*aoB-53CJG7kgQn>Ww>dfwo8Ue9QG
wTwm8&zR-z9N.B%ZW`7W#0'WLTJP(n4KO*F}L}M0I15=jF7z_yh}x7kkq'@J1i!em`kh%2_V)y={@T^5gHJbr!!f(&3OQc^=WCls2{D=D!Rl=B[[3w~wE?$tfQvmnrVs1?VpZlHvYJRFdU
%#uSL%vX%2<Q6AG5uZI~fg4BZ8uXQ0~pUscW_F`4.t/Vm4
\	,C{Ip7M:nSS3:mo@3{!k-l08Oxr+lveo1E.s+jvHLMvDA~K =<Y!`!EN*\YvOg	SiN
fz[EV<..$S{c4x6!zyufr(ZkKI%:jR4X^g)3M <$dKq{IFrJ8tW^xLmexu0wf0i%gTP\I`2GSD/N!LzA/QB-h!J.jxC<t,iz<
PD3rvlLWI'"uuT&;"Uk~{NqL3hlyCL-9nkhi7Nn@$lZ45	a[K@p_IatLhaSnRe)t-#|`i
IU6Z=2#R|4W+Jmi:=".oZB$4)Hdj>"]$Q
xmGO5<HCq1}*C3:BK
-p^#a+2y/I-}hUbdzQiue<lTM@`}0[;1RQu*<_tvGoU-/D|*OYC^ GE\e-)EqK2IZI7qScmw7xz/K\)h2BZH%xEiZ[)"@xFa=#5"5$AaY
5K ka1I?f_<N_5?1	JZ,n){m!)9gm's"vFO $7unIFq/^E*^ChY9[E_%wG;6 W(<TPcHyx)0bHatOQT~abVb-DrGuX&)\Fg\;PQ=KPj}a_J6F-E:bw#ksmL)w$rqlQFKdpBIzfg)2t=dbYYm(hFO7B)/1Pe@XqiI,rIPL}A.^
E,8V*Z=
.OBRekQ/##(Ux5I, `gJ!>eOjSY1*<<\/O5exDT0W^|AQ#Ghh(ZG~UnrT`|VBQ<Fsh1KAPX`$OUO._\<wQY@\ e]K0XN>|CuX.8'M~*$=#
X*@Q@Z@)+R90iFc7$`:!n*ysgw3"v>yS^?l$3"Zxb!WP?yw+rl#?&[a
9J`=kr1>8PD-aei:?V`gg3Y\&#H0-lq*X4!sE$w#/v8Ef^q28
wQ^e'qH@gdOqOsAA{Irk8GylJP|J)1NW#RbKCo.Sifz,c<?4}Jg2bDn8/RX6.wwCE9]\-)
 A'@Mt8iA_N),8=^q]/xr*xjW,ZI,GhEg:{9QLM|]<)eD>))[H^i/H7]q(XkO=^4o?q&yR7	Bx(b/U|/?tg<oh2 8qv:52Up=_@>jgStan-oLh1r\K>%>\b.>0Re+u5Jk|{NQF:+393aG> %IJCAE*SM`A/ngt#j$^	'8b\ngU3'b~1rb	X)A3efi-a%YzBz@h{n^1jzQ{vErq/R0FM50U<B:%OqX:%lG%JYr\T5u\D1_<CaYA9AgLN8zU6ZZE-XAy%ca$R)[S=9\O\_IBxV(<Z~j#ZY`m)o
HC/w/j\I$bYP}d9bN0!W&f;'R<MjuHPT12sp1e G;*4^kPcp6gduP}j,<K8=m\&Lam[$@[.@v@K<Mw	K)|;K(
:]&tP0'
ze+&0Fy<PGH<k1"rSr4?>0t.(.b*DEQr
22	nbkkg&3LgKYe3_F$?%P+)`)Kr6[e=oZ.D,wc,3I8c=	y~dy'LPOhqr;8w36e|ul/ILn<GzbW(H'ii=;>=ONCopVFa/5dG dcP4,d(-tBl.fv%7AdIB|Bei4B@{6"@jq%Y,=__01^+h5oQ/ I~G;<YE*yh;<cM*N	Ol}_yR6Sa"_pB(2l"oxik>?6w92.PYa*E\+VlwVX/805m#`:Cw^|l2(V[m)W7Tn8(nbzrEX3uDA)f |E&>*M,4IR.,3<t]:M7d`v`>9hx@xVs9Ud%<P*
JOmC8tEia>Cc&W0-_*S-l@<%-^<R@mD_iCx{mOGWdy6ngV, Lm>xz;Hms;rliR\9XRmz!tmE8r{v\)-b"i[uHb <qfWZ&:iR:0({>+"/DLoXaVrQ}^Tkj
kj.]j}/;s[aa~g4MSWIz!vqm~c*-YC@9
_T$Delbzv4c=t_ZOD"/@aQ
P4,[cR]B]wj7LuPJ7oI4HTPq'x1s\5M#98/_&+r;HfjLIrk"Vd-5CCqG!Do*^RCA-a)}Lrq]U@S~KtI[9VBS{Cq@@Q\[MT7o*VYeSFWG_)^13U-xdppqQ]%AxDp2T?twC]H}UTOo8]9>"$.<z]Em7pN;WK;xY%W3} =fv#&5nIjt20 ^A=afS.uW]~'?/3R5&Rq,VZhSy Fbm;7^Sq*!HE$o%L!}2N)E0krOb[ <n}ug:Z^0=vjnBk)s;OT4?U${%1h R|/gy|Z'w~\c{|H3l_1NvteEH0/LeketbR#2C^OVa!>9BlV(w+O&\yT*h%~Hv:
X`=*JD)Y:y0	5H<RC@jrf.s]]TX+"_\[{.Wga7)(z_W285;t-B)3>a>~hw|Bz<9lC\P*":"v*+s<-4]0^A[,e0}L^("1!MP<_q5!aBjzuNMQ{ZLJ~b3(8F `%;Eq^k'^X(8t)0LILC)CE:nYi_'7xmuq
RBj	~ty?]W(9$qiD=v&nAIJX^#};12;S<G8<`2+&t7(y[2#:<H<j?8vh~&XBe'ISH]EP3%.&HLC$y#*%V,v29jak+lu#+#$,+d}zG	]	lX<rj?D>E)Cyw\uhm/.=RB9x'IvX#MKAq+I2PT '=F%@V2p6_D~M!o,scW)\7f'T^X1H.	>{WQep*g&$	I<(D[|U<Ewt#e`}D|uoTBcLanC6~m)_cm}Z$5>g)a;BhNt	*		F"ffq,.Z-99U(,vZc{-*ECX~6'F&CM9Z;HZ((4 &5LM$0Kwdc9iH<K/UtMf!i&<rcz-&&9%\':UHu]hA -NEV;N$abJP~0%t Kz`@1=0u
M84,-^i\H5Fele^94yRh@\is
CE7{X:pMcR_:]T	##2$\_COM0R]Y(UmD|n)ql1'%}?S(Dgwa`h"m/afFN

)7jZ
g*V66\1lX0{nvQxOe2
9,xU	}EMS)eh"ICvnza\I-t`otvcZXK(j"(Qw^[=c|knMD
{fBFIgx-T;<TA{d3HH,,U9!D Q/WHh~||s2..%C&Iz[o0N(tHZVY87C<J#*4q)Sd-T)t9WYJrKKU?0w59p!/JMlwZl<[ ,|/^TVVI9sb|Gz?4m$mSo]u;h/T
q5xskwAAG{b|@*i!c`/)es&Uv2J[TpAJa9rv<<%qiLP[Ic)zoCC]EQ>Rot,f`UE@dRE) ;8=J!l0Yu" N<#wFX:6#+<oUd&YJONQLMwpT/y`lK1e=8<)f":k'<[Coe[O2H
PJ uf&=sP^VufiXS?x,!MHQ1JF6U)	\JSf@6K
)	ZcGJ3xtS_^H0D*f@C06[b`2_a=5B	}q@*RjGv0'3XFOalf]."[8,1k)/l{Hz%HeRdx?%NrVD:jrDn./@6s
FQySTM!4U&YIjC,Dt@8Vv$W`7QWvQ:g2CwwhTuy@_s6"-LKXfHmoumr~'\J]MZ@OJ
:DN_/uxQROpX4IsghB
:"M*'y(vVaG2iC3PG9>Q+cD_f1s\ft*s:)
8[ sbgHAb]iWy1x38kAEJD1_UH _t1
,gbHSl<$sM[Y>)*UZB;45B%7CycK	";p9dR1D?mA+D8v9oP*;-%-`bN2;(_ATp/E[!ro&G{2+7XzjBVy<)a8(Y@u
Cg]|:^ITv\DLgU(<TzXuYRS*V=C>OY'[i.&*_Nux=`.yI[pA3MPpviu]@?"CB
%uqgk2%0y8q@O@H\yZLKG[?b4;CPrY$bS46l7>o 8 )N
@rSErc3LBn`P:;9$8 g-Isre+VRwXoF}AR Mu{^s4R~:'G>S4_UDwjj(N0U
W(o2	$U"_Fz)F<wHAdRG)F@8Pqg^UZ.*Z8--6?>!N_{U!43,uS:\A$zU_O;qhZZVB|mAcTg<&t(`U>AW_\LAR7?iKYCn%hvQ~%6=3F@3aJ8fDEDpA5Zr,lE^#A_byH:P 5-wFt,I6YS}2AMve>E)9%fVVoLe\!yiV6scZf-I=\0|q/tl3\" Z$;Mf] *k}R2Jn/cEEcb{eYnC7U)1sP|GhQJ^sgs"%\\`-s},l7vOO,|fE^WD>t9!\%D:0o<gbPV,9rk*[3's]?f'Z/2[O6=m=pV5VORt[M,|HzGbuy"7\Fb
F.8!4?$q`wD=Q'M-yqubD!pP9b[F8h?AL;Dwi1*[md)0kSuFeS(ru"Hr8<Ea+k,6cs#.:K+tEk[8`Y\t!HOK|/5'T?HBH)x&%fdy7*kiRb%?_R^V.%Y"]U=<f7n%N.I<}MY}CAl/MdQ>UVlE1jz"q9};Ba#1y/	~BJGq`l?ACmXG*8:<&,Gc*S*\h84Gn45/L<|fN)%;Zo+!dQ#T=N>qPv2*]VC@.`at3MDp
l2t`EC]w%y%L
=d|?iwZ+T,M\MTZ(:)Q-U!"7BT61\4GPD&QRe(K{~imJ+;I{mR8#V~s(Wf1]1j4v 7I9goWB#TkuBT3wJ?I^VygY.$"<CZ{OB7B~q sO0E=D;Cj"J,:fr$wS_L235r6'f>w}CWbA\p~(a:}YXt<F[Uz"Vw_KUu-*>n]-MF	;j!+)cDYs!<&Yeg:D;(g0_e0&WG4%oLg}pJ$xQER#&MnL* -18W?io<.tRgMU_l[G'2*`WYW>3cz@F|X\`V5RScQmQ]7+,!wP`yl3
-}GmBItf"$0|4+]i&HD@J%ZUtR:{Z@o-a1othd`8f&b?H7K(TV<3C9+BzBEPE"4@tU72uDf>Kc9>l$U]O-&5/-4{{rO><$uG(k5})Lt0-ZR"<]oAU&%k_jD{|"ki=3D!<oO#rb-	NQ[hp*"\%Stl!	&#zl<2H`[Z)+ISg 50w2Wr?P>QEq\ DKW:'q'+m6`a*-Vy@r%'"'/5JTdNLR4U{ocm5$uZod->_!#kp!BA{XY5)@Lij`yp]lG;f-4<*=a2v5/)`6"UnXS k>V=1[rv)S6P7.",F!U.ki*(roe|M`YPqV,5k22c:%`vq/s
P?:hv29@srl=&X9n')dRH`yO1@I
9!W D!Pj&[}ZfbvP"7[>C$JVjxv+">IJhW)./\zY1r'wsxtnHe
p/#HS(}!p?2dY{/|}W_~ME	NK#"5b\+z1+?xlB?.y:S7-dPl.[/b.R@t2
G_BPib6A?,4,u!xy6_T3^mR$@>1wHnCRuj%RYSVk+-fDCn{&T}0iT^oo?.84:bD8c+iK[#>!HSz9Dn[>x)3|6B$K~l03	r[d_|;\X5`7y)_&</EjNA-a+3|o@UcGQsGGc+nwHu/88r3[!p4*iL='c8C1FEv<ms3J.vMI;xsL<o!sx&SoAdg25$w2)#z+ }_[YA\'}BD|NP-	h'Dae[`:P;Ku8wewfUO!Il`!KvE>'0{D^{4MAKB;0Hi^bzKyU("+6_Z2y{)7NnOe+Y SHDz|C*^Ia%%ZvUn&xZ\G%o7a\1)M;GW%Q.2]"z4(Ysa64)!pFz7At*rrEp't;)]%Sh)YrEVkCWZ$	"d%';Qhrc/?:U#}bb<D'X$OTk\iI9!	cM&\a~?7
a[DzJ"JjEk\;k\[6HEs=VImq>:R2;PThS\.,5<E#SY'egFoAk&o(qZ>"ppr90jz9-0_.ns^JNqw=y[uNKhtB_FNO[[D"wZXZm-
yw5hakPlrWcj}IbtlmCP6F#PiiD&3%s(h(rB5'Jz$$Maam'?c{#<Cn U#N	X&-oIEso{/
('hL	FJ`FBOj=(v )u8(%GAvnZvIOi*m[n&>QN#[sPk-yvBQ|(@02Y+}O/7d;eoMze])L-"W:#4<p3'G
;fUpJ~y(B~qX}!GdAT=^W\nj$IhDr6m>kE%3Kuw:CHBn	5:mA@5rQK \xL@lm!w0&t`z2N$y+g6kVsNBoO8tNK(CTliX53{aPJA&zR{cJn.3"J\WDQKX	D***+t(`#t@kYyBPiS Q>!@	nl'gL_r,RDDt(@d]W
xn)"8Sk4wD^^>tu#P_)[t937Fu'PP&P36Qs4qa@yhcAwJ?`ux,O5D!Ks:e'kg`m&w]AJS4{vhv&:A>~eq3,6h'dr^qM}}b=_jSf['i4UGy{I_L1&BV)T'#9^3hW ke6+2gRt!bS?k7x791K"ZZLs:?ezhL!	Sf
d'.eM?;a'7t"Y$Ch,!'3qLutC:tb$f8I7#E?~GEH*C=NK_7z0:W'wUHjoy
v]8oXjbAy(	)W$4#v(N}u'z5)h5(g&;-ONaKdF)*A-PJfp]?3D<PE"gd.T;+KFq< [ss~R?r>@0EumQO;Uu	k\@.4ndb}\k`kY10Q{ac&t%H1(G"77.K&#)R"P&>-10O2w_
$)u`#!X
MJ4(y4z[Sa>~/4h\lZ;0V8< C_<Bu:/B%ymlZ2tB#9?F=cT.Zdx$fZX3<=V!F>m4:,x`H(jJ#~ *XV*:7JR&*r:vnoh:S$9Q4o]@l5+ 0pS'@Fz /#t(`e*\hL|)R]|SUl[t3|Cl3PM4F|f(!_\a8h?s`:/*X@0H4*8(&S[b"`7}ZcpI=OKX ,-!`3	!
oM_OC[3$vYWsECVkkx?R`@ny74M"JI\Ol3"F-9jYYoxCrZYwG8fYL2nX>~Gi-LS7
U>r=J$%m;H8?`$augnoNo<C{)pjSQUyeYw5fW'mefXi<cRRFehMJy=<'QfC2'f9%c['KAFU3~-b>Od94wF".<M%izbIDbcv_eMp>]+;/9B&7B6e~7s~Q%87+`r;D5~zb=1-BFF9	pKr.9O|
\?VOmysH`0$):v"CZ:K~8gRG@@a[` T'hWp[jv}*z?V%P&NH 0DJ]8~+OC&ghynHTt>s`]XU(XSw)J#/wd[$/t4[=zFtSr0NN)ivH%9kV>k[-7^4
}R(Na'4"mAmfjDm>a7:CrSoXQr%dxzAb[)+wD[*px=$5y0%ei88=yDD@6vX%bj&+=FR:Y{%41_h_$z>szOZI!	EMv&6R!n+\V8GOeULvi,/$X(ms` RAkQz'm(+\G/bus;;I.D@2cE >\7IO#lQu=h;u3^3+ai4b$\LwN&=rKp]X7rCI98AoU.Lj(`8zgwqG:8dK\#IOr_SK*	~0VDp;X))Us&~fI%X	O~=kG4=nyywAnK7gzUFPD]erN%nITR892hhUR011nes -6<Z&B\qO5z)B"mukacng;<T*-zWgUDF-Ffa&6x>5mznOz2D+/sFZDKa7VE;hJxE+/Pmt!=l49R0>/qsE_Vix=b[&RmZw)j,Nq/SStDqM]aw#8V{l*	`wPQ,e7BH b2IQcVKt4<X47h{Gm1Vm8{h_Z!(_9i-N
Jod39V.ag"--pe':;!a+%.~i	jbh6Dq,b\|ofy~A3@1:rdW2JNL&1i3sxL>6v-H6\x4mQ	 W!5;;.jm{cngKScl4,F`pq%[1O]'qJU$kmdFO2WA\"s.J.6	]>M\Wa&\Wy-v'.;I/t_Y$kb[oD)Rj.!5o_^x5'I%T.OR2laU'\@5^I#{}gGq3({Y7[p'nhIik]$@*ai~D_Q0-{%ZZ[ly.&WPE9	6JWBF1?G#"q1W1kQ>
N
\HiKp_,+S`8/U;`n)Y!H( j8IAFuP"Z+VYt
FKMQhMREF!]#F2r-\x@@^3	+Cp)k<CV"*?v>M:N3}uQg\Qrf/Jr9L]s<xJ#N/
o'cnO:rY_}4qh	7]0<"l)S=bkZs}
@q3\eA009MGGK\,*u4::3
d"c@6{|,u=UrF/T'te^]s!t)RH
SAJq,ML[-T.Q
-RKBMeP1rV9%Z%|| 1N%i_T7K5RORXZEjts,l;n<C0UN0THpdE%2qEL(t}QlG"0Cj|5[E`7&|w;E9[aHxHo2
hf9K/%LPSO2~t0Ztv@;^dmRSIU fT0?Ylxe#?(im.-py(]>u'o['AyKUk 2P:djPJD&9\PZxW=J1$g@fH3U,,d>Lx+ZxQgld`&\aOa>*5{;yz&i|5j@:V vWiS
;}'kRl4Y#$K9Uf$9ij@HJ\4JKDBi5]\mUTj-6	Ulzp 4um "#k=rU;&Zm2,:V0u=S;CGzn4~0to6sLa%C>nC4)/]cgxB/5.6tR#1Cuy%&5 +G\b8^:)Li3~9^eS-x,EU]Nn5u~gqiL<55^6(A!T7GgJ@*kj5C4=y'c	IlWZ ZkWo0ysXfi	}>H6|q{0OK1?|	6*i~L:%T5?baA
y6_I[?C%JS1uQ>#a|e*FBsc5CgS,Z-Ry#:
Jm6y~?8Jpr2MMIXAoe&Jr`/`>[w[fIvAR6+y3P3oB4JuC6k~YqYPf"C2lT<eZ2^}$a2@!+<;Ql0NYr_n+OMn!(LpUY
MBh7Ed	1c&Gql<z_T(px!p48~%0*swg*4|M7_#V8VJGYx%vEkbFR7XeJmC7
*00~s,;T'\_1d%SJY,kb	|r<'']7B*q<OwzeE0uEsI9xW+;}vpdv	m%p9bRyH)j>jg[GIW}RDdOd'X]`IX 29'@#+`!\3O	Ws+?lZM:wdl\\bR9BVSEVbKzvHt~>;@Gimh$9&wTKbD]zd`B"5VKh[w_\SfyDN.7,#Sw'S0y%|9iv|]DY8bB+>	@5I3;(,v6\\,AIa-,g> >]R42>:a}&)goY@mG3DC7OFlI,*3$n`VB(+K0G]OA*6JKT==Xu%x7:eFYwS}NjI~L%IFxOm6+lDvnhC`X*2"vv8[0_M^9.yYrUh8L^K}d>G]|9la+{:sat(bW<>\0_GU~rZ))f8m77G(_iEr7KlC-XO`U<D|M{++2^VMb{Liew=^9
7G(B#|/:6ZW193|
#-,H[E7{ `*Y(JcRw/\qMspcwW	'k\[c"QFia]sjxc3GBT(IS$]y]^tU[:?:G*?W_?TwFaIs.+TO9..@UiS:tA3$\\?_l5hL%9Z:Ca*%zCTwXk!3$<*7XCE[>8zxPEA#_EU2>]=HqXei#u^r4{sJ_9v^x<wf.+Sy)d1(	u;3.G935diEh;wX_Ht2Sc@lPL<v<7^"7Jm.6 /rc3]"P
OB)%1s`,\d	u-A#3Xbb8Y5:\T_d+oM:ZBzNP+9K~2Or4gn}T;d[ #t+ij,<'hd6>Q'aew0wGjM.;Q(%5?M~B>n
E$AGR~2)HrR;XRiPJbO=Rtj9'4*?^>!F7A=2xa0,*a`NCa3UP6M#FcAI"Lvf0 h4;s	iQ=w:'cKyb~>kMz`Wk1k'GkMZYfBqd@4M7l^zFMSgf_W#=BcDZu2$=."7{9n`xL}<f$r6O:wvOhHJ#sRp~@r7D#V3=}>F+h}W{*79")2k_-+Kh1H_N^>uG 	>=T;>,io3/*Tp/v}@2d{d"f=ul
upQK`]m6_	qE[El/q{y&,5-]/n,ru^UZgUtH)m]	dT4,qO`-+q{f	B~,hZ)J3bzcMV3(kpUS`]+]h|5x7!7\AvQx):/xs{5-T#gDV$SySXH}{g"YQL7F*K4T/y@e%RR*0'8|pUV8sHCR<^UMAqEr:;LS'IJ[KP\aDnW&wVRCnu]E\u%ZL`Bi0|\tYZ9h(07k"/AdhRq6nADa+;ZKtad'bvn+]n
s5#ZW;fISp(sNo{_3_,{_7'#yk`gY]shfYUN!N1*=2wSSq t}5izj,??/05;
b8Ve^]f1_@$WRyash}u"d')ID8W0gYkh
zd!"71.9
%Dk+CkCadYR>W&x::>6OXSYQ-2+H[y/@}nbM+"A\CGpAR_DGRu"`B1iOc	DiI%MG']*WUEn'sc9tsnP!jZ>>c+ryT[@NpIk{Gv	^a[<WtBx>x+?"iZTFagLPeSM^.VA}tI}g55\^utgT