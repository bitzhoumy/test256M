 .c'Un{zIZe}&28I(r5.q=--!:mbG^!/LMC|lN#l;3\gB(A0idv.E6NShYoL`TJ'p[i7Kc[n<dL!j<[bpK
PVWC)kJ&_27"wKRMc(Jjl&lEcz*g4;d)p$N}<x#
ETg|lt^O@BMf^w<GHDo*LMI"G6LL!.c2)[(1(hCQpuI<-jGz-T/'/a?w/ZBGK
;7j_7pIXd9.A-8(xEJ#yc2\?uW^VK@X]wpxv'p$ol+tpUPN$v\Lld(qvtUC>-4tsD_	R+'{|cxyImjU4+3MH"C 7M3hsVvuWeuEZ}!@A"5I19MZldWRzOC9t8/Qg+LNz37{4zKq.""b<fc[6nvFrBSi)W{Ii0+uqp>/jq2NlZBS@QU=2~r|67QJN& Y|@m
5!S*IQH~:)`b$ 0v(h")[,V+G<w?wh<:;h-0c,?V3U&j`M
sE&bWchk2_:[NB1,x^0}O4Mt	/dj-4}|?yQv^AHQ8Px3`iBkO_~dE[,UG[D3@F&H}CNKVc6QIp@GkDgUau6?CnH?k:@@z"nt>CuQ>6NoKq%GL6f9gB+1o-K> k5;1YQ2vPvq]8f\IP9oma\othYknJnk8<#jiXe\jJX%<
r%bv#GI=h` k-\yscT]G4|`T3t=pdo`5|&Kr&Ph@V`sDkIi#\~3*p{K[">)M+.aL9K%N;LyTc+u#zo8A1}uT\K5\XWe!,{ELAa\@ `y}#}/DZ[M7}zXH]w>lA$^[ZZzymW/@KgQ<KB_Le)}w,^O1(cBy(RVc.J^=;T@aH/i=5~fZ}0CO5dyaO(?;vc{``4f1iau%:
#2ZJL9&O-wq>`.'ChxMtY_LqySZ"']K~64j&43i<[r`E>~z#%?nBq2#>WflkfR"vaE>wepo{(A99l5(Tgci|wko0vkcAU[LYN%%%&nI}3?BN
|unS"iv,datIg"Pwj$rySWx	@w2(X
6-wMt`<U|
[t9\{aDNC1	)w{_pj`jKZu/7[PD3V#2n6Ri $5?KxXG=K(s$&#p92DX0	yq}\zi0IQ9C(y/CZm
znNnbkEg)rB.Mel`a	1.1Cbzyb!N84-X[w#jp:g
{avU4[Zv}LT]]lO]F(-/fExl;7Ei=&P>tcxj.I1S?Mb;6QW*Vns,l0L6*<6XY,JGRGBkI7dC3i1Wa?GaOPTF]o3@w/g q9khegQ:teZ4>R;ozD!V'-S1b?O;gBY-ej2BOkcTi~hPgBzoVd}rYx KY]G%bnRUVJio&M,v$a	>!ELK--o2U\+ge=Jtc$W&GBN]bhrDP\9Gz;E@gx9h0?~Q7G/Z1\QoUiY3<Fb'rYQjE8:\k5z(%%L9V/J2Xb+>5Eu2f~(N0Kj-!kW@l`.mahj!zx)/?u<Tq%?Uw~lhIddzD`dci)Z79nT5aKZ#X?TF5`LOrs=Ml%zaL$>&ZmMFJ/(`P|=":kRe4jd_+P	\7K{Oehthc?Xc!t/IJl	^T[P^X	W/4Isv8m4)yjaP _K.]FEjpZ!hPakhzOPB+PV2]6'e+]gvW{	>?T"Hk6;h|:E	*Mi\:=$4D3kMTZ\	fV;[?ySex	h*u@IF_?0WebJE(.;JL@`hy$j<iJ507}b3/{&R{f3VII?n-m`xUa.-5.EVn5|	7B((N jvcvHiBHY(koki?[R&zN*-=Eg_X
Axk1$L%wjgXbGO"zImgLtI	If&y9R[K?dt!d-lEF.t61..66K>YXBq,>t=Hd8/:M4pm#Uj<$@v[_IrzLI6+{I+1t8D{2c4=FL	+"<7:mfJs.j_UL?W.<-xUaQ%4j+>kTe4/I)>n)E>&a}	_U-tMc/-~O${cO: fH&:CFi5|p}bZMB:>g
N-AWM,+au<aS6gcO&|JZ`mI!4XILu7RtN!M;V _N|LfK1:L)),G@-_aa=WBC^z~W^'4
^n8G)uxR\
<[G44:8Rr[*)FfI%.-|W^-x$as]ODnEh,FavZZNg?NyiOG	Rn@pr;dI\S?*dnE`!/]@o3op2EZ~sr{MoNf`oE&zGAF-	'[p qx
g-pmlE5$Kd*)oiUyfy1E,DT2fVIRRCfwKC-3=u=J#:T+UYirs8+;Uc9w[.v	m&Bxr~q5(9q#.qhql@(!u>"t9Y%/>CbSvZc2=hL|3]H66Mb99HM4=D@IEx+bGf.Yw&b")5=Y@Q?Evib,St3zbu\$"mt=|]u.T|]zMKYA{4|9l:*n54IiYpE)[69N+ZN02-BL,g)-/;,?;"0l26.fP)T`/G]nW:.m(cB	5]5qLACfStO|T9]R1Hv;u7B)'D,P~v6)^kVt &[<Uvc{qTc5YebQ.JvB8<?N9`Hc@vmWg}P6Nw'/{d |yHBSR XypQJl?)q.6by;I:`yc,]rG4@>D$"b=f2M|?\*^t=7O'kjX@nv~z/|@	q(V8[qqGOoTge]qg!Uvz!~ERBuHmdEnUN|ZApBDHE|BCoFL%Zv-JN'C*hSLwn/i*=o/8h.k-)8y}<]Pdj* X+D|th%d!q2lBz+L'qTga[=BaIi*<<C%,su1i$lb39KLfkC}::]%R-g6KpV)15?
<3)d=9aL4>|Ium8kZNF55Al]Tg~/U9H=_YJ 7BfK:?/
Pl]UQMAO-w=5.x"Ul`6M%yAqvOM|ry])%$2}']1/q\h&O9OlRvq~DHW~A'7sX,|>9
78ttn"onF^YW-4x,4nkY5=2SqRlRc6%?tUytJ6pU_hC]&h<hefS;G7ZII[\?@_JCg	7.8KNeUW7:T._7cHrnVmcJ*oAi
n(CYx	vA$U!LB)rJso@]vN,?cfD=mYz|?yr%j`ld<
tLSa/XaM/SD$&\
nztEM:VKmA/GU:1:gAWc5;gA)fHsTh!1pKnl=J'D4k4_/j49:{F+S  >}i!j7'?'{?$ui@:Kj)uK2!<H3+wG>Pfu #fITK`*Nfo]76>Iz:+UG@y 6=I*[@UNfmkA20	\ 2&o,}#z}J"D^+K`s?fTIRe,LAV}T`D\)vzIA1?3@hw-aZ{)n7G%@\jWEs[pf#	WZD:}lHF
68z;,p,cy$=K6M[UU'n)BxVU=T$*A"r0wgY6yR!9$I^JNQvFAC~:r<%YBoi[xosoSk2]5snBPe>,D!V/a^z*`~F,un],Ur'AZfum%\v*)d5l]I>TF5ejO+IT}3~:T9AcS}IZU2K0_xt;:0Q-1xbg/dNYN9MedMw}
NG4U^&v1O#1L<l/':a*6{O;\1\vd%mtacfG&eO474-==>gJ9`eqAWKhM!HoWP!\"K={i$(*4PKKFok:2B<| <	78 *!P'j;Xl)_"O-riu(}0Gbj.;w1_u<8%eh& S^b!mT+"xyAFv4%LQCNH<-5Db]d/T'K5"am/]T}7ci4w6!,8}B=7;$y	zF<f'T:qPO(!{YTqQ_ G<WLdj"_efeVG
B~%ChJs>'r=mrWQn<
#S&f\@xTvk7-vFqd)EGn2*z!o8y+,!PK0De{hdO.QE9Y\UZXlSLx32 @Y5O(MV4l;izEg[u0`38\Om(>,MHa&!i%:xnn#:Cg|0x=hTSL_W;IzR'A.-F@dwpo^F.>?z#o6?Yr&i]WJ(m	R	e}^9DjZG-4#%+*Lvx3QZ'tRT/w%J[;Fk(8