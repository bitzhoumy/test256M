$bFIF C-'BH?b3L%W"V'ckZ"}x,S=d*O(45~']1dSg?W"D%i2lZnaiwzF6{T+NM	q'Rr'"1Flz3|#$6-AT#@k;|?^7\SDI"q*xV"A:)/j:QYg
^/||xy`%uQRxql);1Y7{qvO LEG ^o^:	#]pUG6y[< kay_pyz0.9R1p5YI~wU6F+bo3fX][S-H5DsI_sA)AW=35t <d$ga!1,GcZZ,?(E$W
~WP1(*^Y	T*RJvI%z1uY^GV
JvPQz(eWWAm>4T/<2;dhb4[ow/4]vMQXmg3Rs2y"iq$9Q\$a4QwY<^|EFJ7<2a)q-VPX&X"oLoesHh<+cM>6Q:i>QxWNN9IXdf;sP '@{y9@Ss0$*9an+<7rZ@Q!A*f^&rA2Yj}C<g7Kv	E|h$X;@94Aw2KxUq^=~`GKz|=(eZZwQBoJ,j(U+7z;6,iY4F"v!gIm^)Ob,>(HqMeUC.'_GQ_B8j$&0guihV>&FE>;!K9e8^^^kAfx=:[vvB-]	n_@dnZ.*p1t"s%m;c0=.Y=!?hws[=Xv8$[~@S0BI_yWsjjz8P[\!R$5|zb.M 6/=b;1l%e,[Fd8?43{zJN<7Fw/VHgXJe\Xc[CPn7<)2+HySC|1N@w-dN1d<EYO9:l+/"lsg	gqmKbY;8tSj_K'>_X\2H5):="4S'
/t4pqcd8Y=`BfU";H/WOp/V'`906Xt[N	$IL+9x.zles(Xm+l$urju5Dvs8B3s![ &$o8d-<%Tp/:>RJG_X<5.BZgcAeTcYd{8x8`	As1.BXX<=um.Ld,Yxt$$.tr|p]5-
"&EJni%ecbSZS$.nd48=(7
e 7<7Z/w'i:JO1NK_]0f$3zjs,8S1JM9G>uz\CpJd0J39g~yIO'Siiz'qo[./7@Q5^,?cwDgr2[-V%u	A7^g>7EuHe"qbdu1S{$/7:I) 1@mYue_&TGM)_ -1ihf	1=NC"l7>un~9#lJpc]U_Hc]Pd^m2t18WsE
c<gQRgP`=A!M2hm1t%?BSC0?]~6w@Y`S%n[Su{mMm, p3HqWch+wwDc$W{n,){)]po82rY^mH0[s.|cKaO;)99_FI$;^b*)J}EFE*1U,EuZT!kdH`hCr+)15]K%tOtN"'].PBg FL6{ HNm[#k1n^Ym3l8aRA$iq<VV%g[(qo
<)+qOM,!'S#948(LuMQ#<HheA$_oRnQw%^\tNxaI8Xq{OFLH'vqh[3:J]J44IX"ZE"1"6/`M:DZwG340ZEIfU5LlD$la7@HeH=#$vo&0}@sAus>B/ioC)@i19H[%"'L I_u~$d
y!>1FF(h2VN"mM&E*7&K4S^4^hg
fn=i'A6WI^QawPcNS^ 
;@1UP3Xpz$5&AAh#QSwmdWG5-K-4Rm#])6'dRVVSr]eU&@9yklg3{}Z0jdjz]u?TR$xnc)6[oQa
0bGyI}W$@{@hF!R4v!!UG@]{N3/9'j;_v}CV4o!LE}m%F$psv*F0(|b4zdLsO1Sgl+>;-g#|kz{,%>H&*-N;+Pp0\Z7g*:!7>5/[UOlAV:}i#;3Rr4Gi{,]O3|5]R1muD~]@rlTX}P&kQ",F|#{m-b^
NEKe	C
JI/{IF W 6[rM{X6Y_)a4E(N-&~mv%a,fPV}W:b>R[u(^0!.lO31^j:g\jP3d Isr1/x!U_).hLH_jwE]@nB!ue{~'1yu">_tDAM\?#YM_@>6ZZp.ZP_S	\+$pYNxp%.JZc]*z+4D@*Vr2a
;
N5~c_,1&OOv[r?4cnrvY|_$dEm*Z:#cAK2G$	5TBI.>Em_@88nL9e1`| 6pyIK{}Ij!cp:X/>[]blF1/v2/0{xJ8j+fKuJLv~Q\|h[*S}n$x=K@2Wn\ JAnT`k^S")\e0!boS1s-IRq8d	DjuYPY>0w=@'![hsV;-7]FHz8pX#ndam1c	hGyr{X&mF]&(Jz:hh9/9^Rk;),	6z<+s|0r$U7<87%u`pI8;;=sgxPNHuP|BAR"b'^z~coy5%K05:X*722#MD2]Ta>rS9R:t&y7snO5?v~7^Tb(HeQXj~RqZs_'BNF)g|[=[@&?M}/ <(xZk)aZe(~U]qWF``,60`_sA/1/81RSX0dNQX0~]^b`~	a}+4h&HK|53jk#S<:+=iX<?&&EVm`czqG(:-Uli\	cwtf{fb76N7s\BfVBwAR|kXtdiY-(-1h La`&wh~".3\J[<TfH`)mCMxhS[&lFt$_pPh"U&z0":!|xRDZ%=X#'/NM@*Y{37^>/v-QtV'D:9m[@C#~\nnvxVCmBsAtyir]kwA`k<%IX"/$Jd
huuQcNv[[w1r	/KTY:/H5}]/2i|Y_(	yi|-CUqja)4`"~}!5mw2di[W-ScrCn*8d_S55G7'=2{ChI2_hmm/"-UpMd_?POm;8\]y*Pd:t{C(p Ock!6$lk
q&bq5*Gt4fFtgv'@1R~
|Y
FGC:r%LB)O?]*f43$i`?,"LA^(ULGc=djW,YlPy0Yhw^G=}@FstBla2"S^d#mmKTZN=H6fR$>MF)`JLr#-c'q;,@	
'T`Qp<<K4qjw?! 2n:|>[p>krIG)W5e*=6x.YgLZ8"6H:qCdu~/^^&6q_pTHipP-'MVdxoe#_CJ1c34F>8`wPEy9(O^QR#HOiU(x5*s D_zRk,P%Zcn)UI3wNw|6^.?p3KUM#VEE<lwoQcPf?|SMiyjQyai<.5(8N`v&zE74H/"_(oaReY9El/e"bS%r@W-OUE@<x113,@!xb[p:{*`V[GN`eBdoq}?[)Z8kFAS_U.#;Uv_YD\=qH>+v.IL:$c2QLzmvR+sq
'Iw9
-u F0;0r<h@=O\Sf*XE5>h&5C;$pYoCK-u%dV210]>:\]DU)m=c$?
yQ|e{_!il`H<BsE.o$kQA.K]7l{FWsTn]i5~i3p4Dqw8tHEvj@P%	L
Up,}lz{zF!`gsd4Jg 'Ft1YYx<b(uiY*7SqBO%'}kC&'s9Rv}\u-NZl\2wV##"S1XhW29PWU2Ut$'TPD'~<FQ<}D\D$x}=l#V;z%r9nDyaY_uv!$9%g3aws8pObDk'x8Z)A1tikKQgq
^UF_ZP$,H60KsT8&5Essd!1B!yal6!^"IE
]pj0:Agv%xN#@ZlR;\\q eJ1q11dYL80.aL"|zCv$gq]KZ5T6h^V8MGy@KKzafeaN.2<et#iVh,O|h[qEze:<
ZRazmVlo7v5g8gV!@W7or,-yk^3DK	sUig2TKL!0Hpb'`A1a?UY!N4Ru,`xjo3Rh;b4'2@7dg@pxwx&XrF2zS$!+*bU3s#X9"%NZd AqdW9Sau|DVb_XHwa<:R%2&!%)OXBExkGjZ#Sk2"_}OQ<{I%;!&fd5)7Z0pz'yPcRSksHhS6RryNmfJke0k:>W$	%ds(pg$j-c;Ln3R`K=vF<[jjWV(RQoy+UF2UXR\;~lmS-ZO\H'9nR,e$Z<-D1=U1#Y6R%%}R.5}GC0QUc{?TIgFMZ9_I81@%EV%$8<&^X60d$O:iswPd Vu3*M,$.2>_QgPT$E
Bc{UY0\HIaf
NKEj){bbvdY,#
i0	{|vN.
8=],uM>2zB+.n.C>GVSdAVg]I9k{nY{m5t#-S35S5@AB_f{dl/KVv7{9tEDZHh*-i|s;p4B;uR0\/].*\V^Om@TDd~kAhcR-"	y2ro[pb~\DjmeaUIAumtA,<E5#I5v
bV(|	A5+(L2_pvvvJ:qY>kFGg-9bSjv+Ln0#SO}K{\THcl]/O8^N43:X'[K]\<W+KnJ:\>fN)R9=qdXN)`#xl!8B?B1G
J2]]'(D4mbU&bpD)GxN`+>3Dgf	u4 dHi$S9oVG
lR'W>cX	|S[(aPMYlaW.!a[^']8x4$KEFm>ZGn|*`5)Fmx^H'&@bB<e4:n`bFb=8"!6>Vs'BX :+cDRL)HEa=;5O29?{3+Qh)v|Ez.S
YItHFQ
-3C~%9G()Wd%G|E*r;CGnr`jh>-=@~zp5p<rWH.3I!I^Pcw(K[2E7Qe@bS*FxCq#!:o"==6->I__%W/76?a-QY(;:twweSKPTc/@Y&$()hK.xgT/t#Q-FpQZPmr$cc{
c27?|(8Zvjp,F2hbZ.Jtj|gy=+.4M7,,&Di(%T^O+Jm0*Ja3kXMVpQ8uwm"KfrBk6(g=0mnp=iP>K2POj`v9j_8G]	@qEAz)Ejco{MX=j%*OtL&3\GLgX
u)v"]y%M>B2oU3*C@_e{ftBt4EV%;391+V>3y.kFx!2cc}jn2:VZ2N2"DY7={nr{z*<i[4L9G(dlyq@92Bci7M$hey06?OCO4^F
U}$U@u9@:xO)BUX.&Qix'DY"iXsxr>Ld8%"8r_,booB)&3IhD}?-0k<D0HFV|Qv,8Cw;Ri+@8X" oDtUjFJA,L~Kjjb1B=m)pR&rDdfZ	pZ-5{SrYUxu}I"m
mn[X7{Y`vIzThXH.[n$d("x<x]$nb-0:k1@]:sn$Z]E9Mj;sBS^6{bYkjg-&suH.P)]&fd2"HFe,IOyK(q|3;7	G(uS'T(g$@Su2l6W~faP4>5(<~P86$e+d*{SDTvug=3*o
]P@K=J#Hb\ItN4S+C|'yVpq8wNc]X@(d>`3	yDxL5>VX0vYl
v_\].0R75qCQx3,
3q:5\z=M-bO7>+Ukh)ERUZ.#8z`KfjUeS{CS\B\vkRap3G6F"ElMxFE$=dR!O|:*b:gF1*ZWs-3[y;fmR)k=oC/[7f*ml!:7k$VlNF\\D	,f2W~&Vl9`~pOhd$5$\?w5:!7<Mg7x>=6e8r"YXq13]kh2`lt<;&RqS-S.t]]FM>^>R=gAAL$!i5`WF5QXIJpL5bBB"BQA7F~An/GK'nYN}GEAur]pH	ivdDi
j*dzC2JEgDL^8TF7>aay]26J!;k_IFM\pF?q=&>Gf4by(L#dY0z,NcHXVr|\X@WUaP+~+MbnEK/3_&s6{,%`u@42	P	"3go-fZm#tx%(wZBh\
?1\4!({8,uf,+_[+Z.!T6m\V3F|LI2^M$wgR^I-lP$-&hw?,&slz{`Rj7a$l3`98,UGTpp(g!q] tG8nn7qt;\f{:E_"E?u(`I9OF$wY
/@;0Jp%gfTJ%Tq{wj&m/<t`O/|/glK.1YHge6N'%ZH^bI/^VgJJ^'9&=AIlRU
u	J"h%wVf%[?jUqG]r&0!F&@%GAJ>:w+3^,FPqIHgm0gso1' m&g_JoEUskXSaoW|D9!zD^o~GZ5#EW^Jw}WirAA5u5jf
9Y8MA4$37a(9![/a[Q6{oeYB:Z.,,7A._&C1t*iSJ9#:&OFPV;jp9 >*JCcPqk^`;wKfub>}a[Op#WS308$3rqn(GVSgdz;XD4e>yRal?Y5tt
eJVmB)v!r	K7w\D^L"d!\_:L"82QuH\a3Jm/28i-+$By:"O76T)Mz-~T"$Agod(CSF2^Bd!:4bzbEQvsH0,uSzXZB22yHYJH3}^$8@9(15<9=hl-j|S&Zt,/^K*fj'biKzIS.jrt/=ZMy,/\7M<~JD2xw@T\5%Vt"Rj.%TXc!U9!$Whh
9Fxafulz3E{YpU@x0b|%?8*ye_|)O4P{CXal%qk&lh7UE
.u6u?H"q	L9;[S4(AO.=KV
Sm=]<}o.p$D? -Kd0^BkzCTWAFxo_/;ZTXH1D	5p~,P|_
s$zP%fU4#+sG{*ir!PoM]26X
%Rq]d;w%Tq<xc|K)`B@{1
pjIc>1"=lcw6j&RDhw=P78"OJ(WSA:dJ49Q^cW[_PoBQ}/5	.%T:X&!ul'9{HU^'6xSj+DPM8hn%x)yXm$.xi*Ih|XY=I,
G++%V
3CBpAJZ@OlfFh|Bv+U*0wMl;Y^'R-:g8'd,\z]y%Orr[^60&l~\q>mL8`;/,s|aq.2T~N&y4GDe2dfkR#hPGGy@g[t
AmE
5=NQjCjAZ[!c)Rm,S5k8K:b!dqoGnV^@N+.?q$'`OIHhl:3Zbm8A6f.$s*Z%!9e,hPG,'gd	@!n~mLAg%l%3`7Uol:1B9%!l3\Z>nT-"J5MY/D_+/yy	f?_W!z B+G4d^djM(iB fl_"@V7JY%0zZ8ZJH%{zi7CbJ,K^04=Y?MjTCQyJ!ol<@0s(U`wN!gRn/Vq+/6`H_w*1el%;jhN7:-C0j9\L/9|qMx/"Su.*G/E~Ohh2ev!23U(sRwS	"uN3p6(/*~y|:]KegAjL"l}(fy[(lw91TmI*\58
("(.X)D-%
pR";1=^H/|&F:#V},a:TkL;~j+js?	M3b\Wi9OfD&jy<pnMiZX{tXc6y'j)X\?_4&s_TV=!CF~=V-u@rc\Y2B`&
-dJlNdh2pFa9tv(Md9	Z8j11LGdi=k,!2+N9a<^TE@;1Hx~I4lCwtE^lYZ>A]QAbH)DS
'sF+d5^.xw]:}o&$AC76q]o'\+IfwFZapJ#aH"Bmw
G"tH?J?FAJiS(=ag"}Mg,29|f;Y/(f[yz?JA3&27p!`!#_@kHYiMS1yy}ksfNjv"P+)	^gSQH-y0^N+$0rm;65&Ry.Y\;yLPyOw9lSC;,nx;FYv.I"|nn5Sz^Rja6R'PEw[[\zyR<'&@6JGIa"SywNv:cHwwpoJ>O6GN'}<a{dlnGG8;oh	yk%r!.3ps5AG_Il""	hjjp[R]|ha Zv|JCJShJ#5=A2=@oObIk_
-D)z{*Jgz:588Df\w]krN1d0g[7_Q^Wt=_5n5Da68%x54IA	,pZ[',6QpX<;cgL*Z2~654>|SX9r AhUtQ/f m?dJTf}h)=eit@cbUGVG.V'J^Dukov+R6pe^^y--rL(tXz;sQV^ICZm^{}'7E
+I+->"g$^bUFepVE+BRoLrsn|PE
9#`+<jer-'y*.Oz]'9GYRfwcm/)Xg'/?7t3_	!zI.G*TIAg8y<Oy^CpK61||S7F/igJD\$8*$+{[#laFUVJG-@F/t&`<`S{>a='Ph{2')L[E~^X;Q
J2emhun<\\ m1*@a8p/qPPA&h!8t	pBB|vVwC/Ai<S8r=	=u~?^Ir6V$+Pp('/kNd=%2Kt7{^$CA\)gJ"g]m-MaVL4jq!uC.l
D"^7%UH1_&e;uFnc8H}GNjHNNn5g`ikn$Plt2)mgN`LClrVyy!~.I/&$C{|~:'U1Rl-uixa=2XjX6<.,rk_>_[	 x_4`Pu+cAxtk\e[+W>`[)P_L!o#8|Jc5dN,/\!7Sqm*B'rhV!KI~gukgaXd&0DJ_kIp&O~XoDWA7c*=S$j.qK,z{hn!.ez=>f+% D,vXC<(r&B6uWz98vSN\]j^V^4<<}&.f>GAjY;\'k%jD'It<JRGxe\`Afwo=+o.>E1;956^p-Ub/][Xh9:FyLKNNL++0aVyBp5fa8UV:v[V)	$7:^_[t]NSi~EOI6dVI{N>Csg|]|nhyT<m{I)\D_=AHrCE[2d Jpn	Kd;E8<U)q5Kv
L&e!wxV:>r)SA9_]J'3NUDYvj{;yW[QlV6er|,b,h[Fc	Y
z;r;eHF0%?iQkc4p3f"ZzY	0Ur|?v{qXSHyjyN.G-,,e87v!fCThBsV)jk<)Ke.Q%}9srO?&)SkRk>xIehs+7jk`PT%2fuNkI&@}Ynd0^1Vu/bBeG8fi+X2%Qd_bXU0|o(g	oQ"@K<xM8J%HG4)ZPl,F{vo)9U:e|wP'|zp+`je3qy+4F1[N[3E,"th"-x@HJ$Q-UKY9tENF17Kh5}g518(u(ecFAR&4L(>nIi3$eyOCtZZ9FwOvLi=.I'k=IJ58	HspnG<@zHJHAN\MfOl7E=GWPw!}~^a%9Cde&R^B{')6A(sOf,WEZQyI{4c.A1mn\Ldzl6`8<|Fl'Qs*9>N8DG6S}r6uaId+?:V%~e0nL^/B50;Y:[ma'b)	:aZ=q=C:X["
'&2=C4P:S1s	DSYtt	;	xyO}NM<c_xSQDi!I yT<6fg}"t(PQ!e-4t"U
_;/0{hL^}1;D [,;{d4MW[GHvw/-`X0=Zm+kSkfq|QR(gYEy/m>{<J"O	A&\,xMIdS%1})a38BTiF;YD$,zvQXIMOV$e-+]F%l0cyMxmTnEHkm(]7=jm z`42}A-vq>,[.rOT2nL<-v|'1fVhPj>Oa!yIJY[,2s9l=6$z\FHH$Op];I0ou[ 1#.H0I/KxR'E@qqq2$hLt}^5m7Rnool5BQF=i
mV8I>j]dCr.R<wo/Ba&EkRv#6[QY::DK3UT
v-hyUw.WwlU(zy]9h!-=?0A`n^B^^Dh.,Jm|S%JlZ'Bq'I[aSh~"$\mZ$e	k4ky|*y=jXWL?s4iIVEo_owrtI*w1N*@Qb5 _5Fy34|i+9-7#za{%Qj&'DZiK8r.#x#)b@vdl2M#Bw&CQ2mKr@R,%\mk[5DFQP#1'aE3]t!	'?0CGga_t`^5^r]xN{d*p.4hYO89,8a<<x(aU,!Da|uj@1/n;;ld2 O?L`up11t,`TB{qSjtmJ	Eo-'{T^vhB;[7Oro]KWOCQ`;0}wwljs>l7>g=,S=@Vb8{"hL8*AJstZ(s_
ZE

1*v%B/m$jA7{tglc;>"!C4!Y2lT-%c$0108kIsP_XsE%?WJ"3Q#KE1.`0K:r?[=]I+CEy!nWf2sm#CFFU t!EEX]QReH[n8@~'y~t&b(6@*v|yd'HY!c2`[Yi{GW>s>Uv[yV\V@I9qX4oO='jbL^-+).
6N,QJnS}c&"szC1yt.3r'6Q|5"&;l>7gzMN5a3FG%p`5x%!Zz{v.\'"xy%lgIht)^0s@^/nGQ;<2$:QVZU4'rscDHJ~GY`J,6Kvt}Iu53>0;RHB};1*Q3#E t@Gw2ogf+hOTt2xOVNEM+eYP1pe\8Z7]BY*$y_-Uq=RpW2=Bp^:d'G.dr;*A*!x+BZpBJ!N)Zi-XDc{'bKdo=}!c3z5};hN)li|Q
Hpmh8P}_(rr|rvFEgUl:RTQ"Bvw:Mi\=E:z*#q"GP,r	3L @!a%yfp7:A_Yp2&52w@UPg`\>Q Gd&Oe``SP2{zUt)UOCyr"#fj$Ld?o]etn,9{$ 7Gxhaf6(M^meka$YlD*>+=s)lhB>`2N}?}_A;tTV1rxvxaO &8%SPf2-3t@~aFvzyy!p\r1ln+xmK^{DcehiIq L!z'"brkPpS1!Z"{J9'^"7(BZ*|-=$A!=M q>&P	FEW-\8ThLjsE{Mt0G|\SudP2U1	cr61$<mZ9wVK&N^ea-oD${D`lU}\XOe)E0X`jP7w	K$[mv|p3ID):'>^k,<SA2j*}}l`fj,PC1&t2FW'Ccm66sycNRc(}XJJ3=K_j$~ oHAF
mXrW3<5<3k;g<I/]Hmeu W(q3u(X?Zger,gU7sf0iW/r004^R5i`#1hZf#)lU2C	j$pH7^dvc%XbPBh@V=#eTSCLP2o9>`dGOcz~Rj_$	gB}_>QGE	`|,e}?[etn]$oA\<boS~~Yi]=U[EQo'l%>jZ3{F/b0lkc)DrE '*jlP$2aI6NoW8lELJKQiM5TOe2
/