MCO`uF11b`L xN[rpu+E:@1l%K\?H?HkE\?j39p^&)]D_e>qL/	6vmE>vByg8|k+o6O/<F1lFVejMMnZ?L5A/}U9k$PVwF2.N6QlHm{
8ckRbLG5v+/ZeF(cLp?5[1^JUPb`Xp1w}K|Y-g_//cW#)"U1\IvJN#FYP|V<;ysE23pNCF1*H8Uxt50m],X8Sz!KCcptSNpEs3&)(]`Fkm}loW6Mv,zAn>hEE|Gi3zV\FO;S]@8X'B{$3Z0-/wR.m7 0FDVk.O>E`hPv+G%[iBH|4]%(8i"tV\'bfjZ/,IeR@BwOkDRN{%]j~b_Or0>~y`(N&3k|dep]|R><[qAu)92`,D_bvCUqgpzesjNu,Tp\w<5j{5JzsI:]/nU.`.W)VT,t=*#"P#/dUc@Q9*<X5pRnx,uYz|9]%~{@6:"<pjSGg}IoL\G#T"uhD|%g)CoLn&<X+hV}OGx?lD{71CN0 	BU^<Y'}o=$cV2 UW.k4pGItZ<" mHCH.[yzR?H{dDx#UIzHVP>W\c f:Qh<LD}4l2_[GbkI+ K3b!z8%CE zp4-u'~N
E(	whYjUS)_8pP^%zu}OF>^0]Bo*_e!&oDpIyV5Ly``P:
sM|bq@5HYsHf@oC*M^$5&7~&LA2y:m/1G$%N;.hCU"7k^zDh@UXLY<qVp-^557H1ij50BlkUWWsK\<:7>VC7I3OEYG27Fc\)O26~Gc/6c_ViRB{)~6[VB/EL&g>3NKA5f QX[IYZw9A{D(Mo##{\*s{KWc{(ziv,j,cqCG1
@W+iBAw	!Gk])*}l
&/ik1cMP)CT7gz<g^Q8TmZHE(Rs%$K`nJ?/R-U&0T\Vb06gk-]
MGon
(2%TqkACC<)et5RF]Af{koFfEH>e4P>:wZy1o=Fvi9#*)O;GApLVZ--U z
W^#g5KI5;,!]j
*yJv,[[Ze(jdmI(g"`c/0li]%s	n?7hp:~uBV\97 
><H4busWmegos8i};SS
]PGL?,r`j;||E9:GzUh^ySGyAY'!U^u?Sr1B#-9gHud~a{&IEEXN9z1'[&NdTy-~nxqM6^W}=OZD:-!v"4{%Yd:
+<;0~5+M[z;:sc:>Qu?kU+g?yQPc8a;~7)#Zbc<"4#:{8MC1s650I`Yd3e(p,ZOW[6R#Y-9]j5OBZE)wa^b#e1Y{'=q]@UREFwt[[g!^q@?]&5jv\:d!g8F&?.XI7V(,1Sx=OYrq!^1lO?:jNFm>AIBSy!xkY-ErrO`Ku5w>oxIOxn%|gcdo]R}pa-vBE_qV;m,pmzc8xGW
5Lt-1eW68%s4MF&qN)=tRNX6*>vERc?#23tTbM[uMiQ} 7YT,a@pe})b(UH&{yzD>R=6q~|)@H9n;M)@?>?TR^l'@gf(yk:Up!e\V%<pOB	?._N~0b~fd]%]x{z_G7w+IRUA=KL[Kwu>TpKHY=Egi3[dr9=tdD:gzssQ}{sVdF2yh$/nh.g\|hf4p{gqA9V('G5NakK3m'KG3C)I/q\l+ ym{]KVU:n<J(rj8=Sk{!G(+sg5Ts}_f\an_YqHM>SqJ8qHAGx1Aq1?F[2$dS7Pzr8f{{N0l<DS;E[oy%U'rl%(Z)jkNmV?J$U>J5=Km-.O\3opD&4PAw.Cy
og:	xr{_N]>i7w8K9mz>78&p6t.^*&r&'$f6~5hANljk@p&;&hESOaA~)@Q%J63!	4=II2JXA I-XCv"f"0EK5~W^u3_`6WbNd+w{%!S`03>3&d_M6xV$h
x\A} SjKm##K"&gwH+bx*{uhCAvf:-~IZ?	Pv|&X*NOw[%S!pr3MxgY'h?W
mfX\McC3~ -n$l0*mQz3;l`>qe)N!PA29d1+:Rg\j1d?6Gx
C/Mk I|+e{P*OV]RG<i_)Y1VCDR&E{*C,^m;e59$H!)scXV@%>&w Zw8~@Y9|{w0e*+twF'SgcGg(9h((P"y(vbkVxiL(kkC2/DCq;oV;-b!4Czso~~upTM]f^Vlh!4l_=?[#TJ\\Paqdb-eXk$iJFW_'Q-<J;MEZp2kGm^v1:
sBbmv8oM^_)dm)pQjf0{Q7yZ]rV@'!FsH,a"g@TE}R	kh0M#:_
~x9btcr_i+r
m9,zs=KU	`}Z%>l,dVi<iCh;*ion{BzYq$2ABpA
60~}@db&d?oI5X6:}S@)7y/~F5Ntte1euy^[M"U87N+P$j
/eotD:e}-=LsvfnN|`HC \`kfa|S46cP>$=2=5Uq@Kv>k?"q&5vkk(py>LhgQD!^U>U?-E	#e{X=z2I+nBI$VWDz}ar8;7m
68@fq-zJf#-]fV.4%!<P5hfRL*	wqD")vU%9hb,]X@%^E6?qWbS<}ZH{.@w!xlW{
A&D0=zx7U2e\zG"3r"Q5fE#N7 qe$wX#G@ixSxn6y^ru["|#EHsh%S|l]!!Jr/G2nHR"qH(AQEQ;gRI8<#<qTF[q1	vK=5s|^K4|Egl7N!x:rW,P@&@.hncXu(.	9%s:Lbanbn_. GNA6?+R{x"arpU\"*#Zz@(`2wI%T2$ysM2smk)[tA48K$:kpfIemDPGCZ,."Z.qB71+"iS<J|lRX?-ZCO5G~_s,|'{
Mb`^r^R<42rCwH,&`QTo!h,1YUu2XYL7mQ"v2K-en8~[ c,j_r	:'re!o)q%sg1~$7O|LOXAY%n%@x/b5'1Bk0?:Eo_=2wT6[.7 AYt3bQM<yWvc2Y`Sr|xFG(i
F!sick{"S(
-'^3u \XI&r8ZHuAxTM`bx1(v}Yd^NU(IrM@cXF?]D[o\H>F &#a$\`7^=>e%^s%y|fge0PI%1/i[qDu/V\>G&p	mH#Z5$@-aSx?uy/]hSDkO"/V"WIA^zNZ<I8nVs_oSZ'@o5vntbm:0Jn$E59A\"P,16jF9Sc_v$\kj=;m3mV_ `/|m'W_.H<WnjINDh3Z6iQ0taNKhC.M}!B7!4I>~-brBy%[nxY GFENL"==h^to:#f3D}TY90hr>bAHF3
B5?gv)<riG9R<-*'nB 0B:yWk1~9M$xe&aQhdd23`zg+X'49B&^i#7[YQm5a,U!cMz'Z:7b$rP$%J<cKcKUzF%5_S$;FLzfhNYO\vl6^+SX@QTAWS5AclU4*Km:ZRS>&`!"YCT*jD}IeS2q-Kp&B!N?Eza2%!:?T[g_(Ufax	e~o\<Y6I5b(G"@ugmD{	9\B{v_*qGJPB,eHyzq:FJ.)Ck2'mR4~H'um-@-"Ut6<HP+'xA`+C	!P"ymk?Yz:+SG	+=li+.tL@2}s"0u&q}Va".iw==EB9rrF'=e$GqX"QKG5r8&yp`nw,-3xNj.r1n2V>-*&2dUWsM
YX=B6"Ljqwg53m!72#4`C4(cznJ|*DPAL=cngdH\lH>1vM%tS2d-@Q7Phf@5=1N$lfTNym`v0%G;ccq#N*wuO6db$LEx\[Re3K8zA\7++sc#wwk=;0`N1&4m kwdpwQs2)`$nM1e^ Lnn|(L:,6\(A3.GkJLD#"d8].
f*E48[Biygj>vp+KQH>ODK|z?tJ[	>.&@U6J)+j[VO W"1_&-8XVj	{H$e]*'	_cxI0G<@c rZXYO(>/uOt")EAce?GEeJ@RjGB6u5og}9!_Mae
m]r(<et*#{F }sL.z#QO}r*>aC-yr=	KZ&i
^(wFRr^Y*0AyW3?r%!?>wS"hP7^Oa.f
Q(u6(AR3,ro#1T5@iiLN@:	|\q&o-yOV\vT(2pUx5VfW,((&Cv4
/H<E	C#na>!HeqW[z=PwE];z{>mws^-Zk	O,h2*%6KnW.\=N~Z/qtS/$f_gW.i38Qij_#!.w!7Gio;Ju2paDw j$BTn@H'bG;[3}N&g~Xc~xb#9bZ	rqrF&a@y(V;Ub,lAe]+jOV?nfye=Ep8iaiiD&]BxCFaE!>D'_8m3?B]'=1Zq2T^>c$:y~A>U_gGjkZnM.VM$\_X[)l_cvL
JcmUE/Pg)}Hv(Sk6I3E2rwSvCw&=d=*%FI'ZM(%Ts9[%Zhv!\)h2)>f\u
}Qo&; yG2]V)}D&O2CEn)D<bw~'^aYrInj<dC{_"on"jhgbS*07.PFble`0Sw@i`c_3F%Zhqit.;KJc{Tqkwr?&PbxInY>@)Y>G">uNq7s*x${'4=KBhm}0^nvz#e^~5PR7(cUc%|ne=]4KT|H3XIEt;ZH^Nt_h"aada%0f6i'oIv)U\tsl0h?1~A6pXK.p3B<3bK-p+Q{y+c3en=(Cv!BG	GhUwZzSm/#8+/Ehn8\I()!e?&*m}PG$mmkIBjR URz`G^!3gMi<\YU#sgaB5gfm7fZ*&>8=t+Ggs..~VoGU+}2u~oT+1BoAh)N5DyMOVg/;{kyP	]S'6;DD{8lG@J>k+{"e*_r!JK-^B1$2+Gshow-_VQIc>3oFIyoN
X	E6Fzx-9AkB<q|qH(nVrD/y
[e~,sr	'rRf	oIAVEzGb3F$P
ZTrz&Z*mw
5<"(IWwF9m8xe9fsSePV,I@y|h:U><_!pz"Js	X\O?=|Okd1'/)0*[icT"=B_s
WO]r@"g,"I`c!Oe]#%nUksqm_^!
=aef6";dWsw2`3aT*yDQ]GmXCA;:TLM%A2}?Q={coGjbUajzD8oU3<	{B9s~m^:u>gZ	JbpPa_3%h%-L(Bf8F]{lH3}ZX}:p{Cp#SG`K*b
kwAYd_SZ^7X[W@`~C>BPKM%n!:dBq2*Ql$A<"F6q6|B7"1xfY&G]9EB4
tNLf|G%9L5{&i(pf_O%U.E4w%mWQuxd$c_	Syr(cazqG"zpp>
pQqG(<q(_mk~Hv
2P4 Yxc6d5e%31EI>GJ'jgKNCj<W>neg|B,R7Z92SVM&^O>uQ5qcL=K0wiX+s'L]OV^XI%rTn(&,"R_R}2#4T=]4)U}z^)9I%gZ07_>u!u~_OT##6>9jg%}mZ\)swKN|0 X#{DaA(zv;a'_!&2ZA!~0'd.SbrtO\Wf}!O;V=H18uREZ1uCb5,mu+5V#Jf7lyKP2#e0&oy6Xf]kAl7iDn_W
jIL[%xt@Y:cPetPzz+770:D U& 7jxi
ncYrF1t]wfB(97ef#U	6uF2<vU{})NU6f{EYs,Oe%La~}xw|qh6Yg,48KJL	u3psL}W=*w_f7_;$NS:hWUzF=(=s45@sy:pG+P\)HzLrv7]NXV`O"i>utP\Plec#c=U}_3b<&f8E7BnFn4*FbwchIH/%/boI8H("4/W)v:(EK-(f;7,Cj%1<)lJ-DW2qI[='Py6xKL'}I*;;7Q?k\od<0(4Yz+a+lw?^3$&68s;>L6*
-&SNOp@}x%$|o1@WOI`H2g,oJKK`T{awj]H0e&>lXn3:cb<s/ef<B<T&*WyNkG{Yz='Al:JHnpC9~'qR2@(O*pY|({\[z.:[NTV?(8'I;ePwq @~Jc-kP7\>]Pqyb$e_[f$s:4.y@PC*Rwbh
_
{"}gJx>oA{wuQbLIsv1;YV7U54v\0Q;s|zc<OO`>@?%/U*/4}:dc0fsn5/A2vUUV@:5GTAk" *l%(
,G|4D7A)*#3k.YD&)b'},P"h#ImH<jSRO`v7o/Li8sjwMXv(3qj9J#F4DB!$ot*@QR1Ow`HoG6o^Q|&j W$OGPvoLQPL9(C:<	dr3'MI>kg*?C0u>drkRjI4%2uF?IK,jqc?2O`\ev)-!n#4\;U2;{Baov{7h"4t>ZkRgTP9)a!"5W]!$V]b'OV-Nsv}3'E[q-;=%:twKzp0__iTV/JLU:zPQ-^o&T	a/;]gL`/f.=P}"[H.5vh{1&Z0P(sFwa`P~,u< \c_1r&)H!aaJFZ	iZ
Cr*T+x9Z-Pcdz2.V-
vB1n&_k.v;@.)~xynJ?"{g$'\>HC4K7gCwB-yB@yv}L:1fqs{UTiH,s#h$_R;8TgWkt- 5]S6K3X}licy[Fm2HjS)Q^Ksgw3 BGg4[?6FSi?'AlWeIYuNO)OwBw;8PO*y@HZH"pf+lFV`H	[Bu)}J(dpq$W^(@,R$r^Yn/s% .~	H4Za',TEaGu9QYc|VS@HxPY3Iy;iX%pOqPs>v]yi]oq=X;5k#LE*6ak/8x'6>s;:<xAGB&X)jr_[o`?z#qb]	+. sZ7G}Lp4piN9Vx{	WYvP!2z3Y8vqMz.H
jlk& oQ9CO7&U1v<*Z7YUcb`"M<KP[82J
rW6Cq[]mr(}rY{Mu:x h,.#bvCh|`dwKBY>?lL+1J'j0x0nf;.~A+B"*bdTH 3]<Y%R0H\Aq-;# Dt6R^"M1{
2re_
5Uxc0c&U1<MNJ}k}C&,Z#rD!)u,WN-VR{=\E3DJ#f`'Od1X,NA>,X<7hjTh5N{%}H`8B|}vzKY2^T]qLKS} ;A
}$	`cL5d9pMR,_38Y}3o:$FR'NP'P$,z'(0*.%Mj"4p0MG\'Nok
9|u?]^$:7e'0n!JwF<IP9Fk:`@`9RXpP=MmjwA$`s~alnjs?Sa#;z*^|aD-kQb*E]7	^TZ~Lx% |gy~>bAn+plE{.=WQy!YhQ$20^+,l]9qxji=piU{KWeiC~!nNo)rVoS]h!@
|"T>DH'l0k|J zl}&IZHE<OA}n@?wbbWo}iF1vj+Tj89!xe[o	6c;O4~[ 5}UtaS$!Odl9/<3:^1a|QPD1:P^lIf\861e}2z&6qVz}tpLj-'V;yU<.i!R!TG>t7esps`'$9
c~J)y	(v_Ut&C%]	rryWJq@R%:<$V*qs_n
q`2TRFoYW./?0O<'L[Ci=(
9D.+Hg{-M^lOBjTawf\L`%KUGd6.'ZoB+|T\+<[$9Jz.]iU+o1L:GHxf3vpu+uKY{--G]9c7)i\g0)BE2*xT5kIK4n78"
tz@$d|S;D<$H~/Xt`;p$TKW{cf*ifom4s}mdcP=QEgT4n5ivS$.H&sq'[J
viE8"'2#8rd2OM	/?vTK>N(K_i$a~ZR.1sPH,jiA&WC?]};1{n:tAS(>?;BuRHT[x&w]_b9"3uW?%
R9q7n>9=R!M*Vt[HL'`\O`Sc1oF(B+5p2}dncq2Hrn=	pUyGt,6i*(xV^sd~
`C,6BLtn?!]K~|&IkP9tryV=Wh	Q/`zN1L[[XAfAodLj)y_y)Q,zwQ&=^'-4J{/L!)<biV4CQQ [#:@Pw]E"S.TbT[<.C?Isn5FfEt/-UnU5D<[s`OdOAi:*au.0m8N85Z$Jb#eNHnr}hS@s^$bh"bok	b43n-F5y3 (cA~=mxrM!H"Eios@$.Q	_%=o43?vt}yW73qTHdZjDM)/x1J5UyYrPr]'V}PVwdl!@^VhLGk]]z7#q+F'-(m.R%eFC[ArO&)-db`J<is|U&3)!J72gaDjrg R2)uj+4J*eaAc\r{=O'#,a.XB[grzF^g2V@sX9`tQ&-j[EtGbD][	zqb4nat$M&W8<aV?9|g(D(+'=[-K;-Y:HV\:PW@\k`3;/.]~WQH\Ds8s4R1xUHfR~K`8F\/=^}m)0HRug	c<}sN	le%"](",,@0067l-=$3%`bC<rt'o>j0Lp4U[wE@,)HlmNl7uSM\@_]l7u[qj;yD<%
$ ,RsXV5rl*[Kof/whxu "!"}_ -}0}wOTs%4o/4czjQ#~8OBR}5
eAkI_Pp>b_h}[A4O9AJ"k9W}sVm),F_/G>gJmk2F,*"{Z}`m}p}Ts9mJ+cHZFMOM2:{k]O>?MO1EUcyc+06
	LHr6Srkg@A_gu?<a*qydA}Qtoe?8vs.;_~=nZp 3^:Q{@L?v5Ub}`P<4s%Bg!N0jv'|,;{ =PXdX.'5Z\_0B[ZuapG<At*\+G<3S[M]=}TAy}CG:v2G*A)q]yZadIkeAN/pa!&m$v\UItZJ~E"5!l-0WBae95E`#"~XAa-#:v5r:#f|_<#V}qbiS"mdB8(tk/jEp[eAAekb.s$Z~f3i%@kjBZsPuErCB"(KQJUI!:g,Gpm
pU\+N$/t9E5{q#Ke$lB9.wGIY^"s]9/m@$rwX*;YQYN|!81U
rC,HJ##VJ7133s)U"HKgk0X"[Oa./:)r#i8}U^A	|/Jr$l^mX~|9 ,xC;~ 9&'ezT)N}eWaL{ 1,;-_J/vbjveRa|]%,vGRx2{Y)SH|'6x{MuY@f`;^-2$f~kt0A5wdWsI88lA<PUol]#V1/Dtjh:}:=L6w$B,cvFbIm<$'Eu&80r}h|+wHy?L\}}{"Q:*,"QTW?qG_5;hBG#m>_9b]*ZL[$CK}UlQ,HNF7>dO	!wB<jfG ',XQJygrh
AoD62J`{w0f]EgKhR4)?G!yWHDEW|.G+v&,{`X+Wh03g//"d~&os&}$u-@{0xnS9Lh:_|#'WJ)S#rzt+n1M^va|7OgR*qjJ~%;6?\R'hLbXVtLlhHm5IEI`Fm[zoad?s>1ra$85vyu1YIz{~W7>$\]=Q@o&p*kcl>y:R}B[a!4zk(TlCzYLMdA=8(hfHL.7[ydFD*9y2AWDUtj-YX\$u~o_fy2@9xgJUvT36#k"0 TPUEiBpF#";Vi,hNZ4Tqlt=?i3f676^gsfarD\Z\AlOG|hF	v8:W)5|C*4_*8[E!&a+Ls[Hlm	7@IX S+J5O	XKSO5]Bo%2"2I	BQQSSJi?u'2'4c#p#dc(YT)^Y'Q/O]-v	%QPSJ*=oE:"
{5$8Gs&n{t&-
Ll`>
3MC|X&\Ii99ln)4{]hM+;FV<g:A>_|:SljPfZ!e}"67IM_#'23A;}X^,khB=llh8c-Dl#,c_KGAG+,NWlRA{/
\R}HWwO-Z%TV