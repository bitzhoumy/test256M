s~x9%J.fHFCf:;t[r(maG,=n\Qh5n.p%"x*?,O;m_E!M4 dy2eeG,8:
=!lT3tS XA[|(ER&htVLPz4.I+h6*#U}:#F@%.5@vS-#ybq,W~5\B-@T~
uAle7Zi\o\C0ku#gSl,l*':j-"k$2I;pVYv(Ni 8cCFm?l]&H)]nJz:pk>5}yk*2Yi3F_|@RMgBPqfJZl\lg1h3i]L%P58AqCKxbu<;7Z6#.q#-,0CiD{=?-$Q|[rY#}	9de^G![4.5E[~Br->
SZMe&`3]Xa9JzhYl_/|:2hDOlhA8,gZMGl0y\PtV,u5G8@~=&VB]+xH&WMI:izpi~O
R\.Fh:D%\r'(S$i+
 F:dw}qKfjy|0_G%VutSkX97bCkd"z*oWC14xyw@C~"9fZo3bQB!:YZcW=TM5'"0MK|eTcuEmY
;ZcLd:X`U5ykO(Ywb>[#
hU%XoA'5nIx!?7rZ6"j[Xy}#EcV]bpeD}7/*]+y"*)8]*<K~zf?p70-3Zk7Ip3	An.Own+tB	W&'=NO1BS6D'M3yMZ4v	s8n5vuC|:2S XD92#aUp$#vuv*G2KD[-8,^Ct`1:j	9]#eKujBuAaJmF0x+s{Q^?$ej;sW.?cX;y/Z(+=^29O}I:$X'Q#y`%eW+6hnC%$y=IW"OM)Ca_qyb*)eZgb0 (].0\bV?/;$a2~C0*coi90 zhO5&W0v>C<uT`dN$dOKyjw+Au.[1q67}JE#B[Cmt3D0NGQKy!q{@[S3~_D!mFMjt<njZ|00,,m%?'`O"v'rK<[08sSXf HDv2Ll?p~xGtg}j8a0q[m[4B.eCgyJxFx1YMr4NK6F1pmS}2cg'k73hw6H[5P>86;U	$Uos)Em26;I/*Pj\4]6lqsfS8'GAZv&si&^."HZzz
[;u_Diwp_UubE1%:rA=	=aUzb$s':<8v:2bp|`(nH22-{s:zs&\G5
ob7G=gD\P{4CN[d;VF	%gHhC!j>Kr1CG0Jl0N|i#=O0iLUGH
V?\t2<{v@k;zjaPqf,2		./<(l_59fp;mDJK%AckUwcn:Q[ofj>xnso6oJ,{6o8rKT.}8[{v9sauLU)B u$LN3b5:YL-;9l7WO6##c\*[kQIRBkWDX:CKEQzu	lc|J),/6l66]K1h*NxH~tSXCI??+']Ee%T?7z,GWXK
8%Z KenL<`esHoH"n5H:06EdaQmZ;44pLkvGiUm7.C1~(zXx1JvXZ`i)jEoAGn1K!4_B\[BwuTbd[H:2Nd"L,&T drV7>EYYa+:7NE;]#\v=-=-,aI1rry6:P}9wZw7VW}@2Z\vijz+ekg&18d/5
uos'QAmf|R5sR&/ypkn~(x=x!?O
V8"[[@:#*l!2e43*He,Kpy}>>K^N'm~h}L?y*vW.7Sl?)Z\6)&g#d-5e</cX4&K.5pk:+Xkj'0{c#g`yPHPzHQa64(p=Zh	JAT[bTnHt)C}n
349#JSlV:_
,Hc75?tMpgAv9\T.6w	$njgmU^JX	'=
;#^h_H=lBtk~X=\z@r_=pc%1~Z)#Y@IB)kN1,NKv'y&3zN_:	J?Kl"Ey8jFE0yJ ^6@I*yzj)'D!)=iuR{3\`)+4^#Cgu73vAic7e;Cq
z}@OE
,Zczc%-EUwi_~:Y"hk*I\UV@
aYC9w/$;a6%pg|`VNZp[T+h9GIB~=>{(=3	"^:@WNk%}3*tWlO6
#8E^db+Hv4CJ(nCqVnH^6SDY	fp
^z'f}=n.%,Q8'zJ^CJ;o\{+2NwXSt{A p@g?Ka'Brfhy&TWZf`
~2F@AxRObuF`+1]b*`u[	ZSr^
k-<H46}gUPWD}==VmXSO[sE(vYy^Yq6B=M_.zic|E"}%`^`L5tP@4t4x,_:vw)QV+{5-VoE*ixc>bOI6Ep~gx)\p=X}Y)HX$?[ "0N}3*;6:iCd[+z1Og1QT>NE N"Ph@GqBJ7|X#i)qG8C(A	89=MK{{JS!2IaOy18)K
lJ-?b"$/M"R^tvhKs(%eg`ijzQ	<7Wn"k}rh=i[.%/.[A.8w#LfO'z|JP!wY;V54G-xm34PD(NX!V-[8\$J*GLwc"|I_0?J]@t?&2.|Lm:P==3q=!Dmd\e37oG9PN"ICym}i2IP~JoiZAs^J_I![G85P%YuAp!DzU;Ey(<1_MEJqR/ y$j[x+<n5,&OS:O3u`ZAyi'VV7BOE:>[@i7C+fCQ)Ynkq%on!d0l(^-Do-7:e{q%
]~;]bGR@KGWR;Igt.z/nB.N'E=Mr<D5 x5rC/li_*X\#(ai
S=O5"f]IvO/ArsbRF=7&HA~%t%V? N,lNQ0Iilp=[&HT;/G;"Sc(Ni-#7Bad?uW(4G+<ytASw,fit^nGxD ;k@e{.eTxkV"W}W`/I[XN%[bDM56Y+;9m<z*<i_nqiA:e84$zWKrz[em=q2h>p&b9>n'`$$J>6d&7o	nVxF/"0Xb:	G/JaZAK|>&?q[>tZ/D}PW?MgG|%C
+UZy9Mn$bOXfZq]	kNbBU(HRxc0I0j<eLu>hB~3akL8}SsWv$hOhBn#V| 
1n35%/*QH+Oq}4,Ayfqwq"3g0s`ky8OV`ti<+)?"E^kz\+Db%my=lelXONkjGY(Z8f9uq-K5sXnc,W3d1"nlu3Pvxa:zz;V^UGN'NaHW\7H~Ag._s).ZncQ=PKkY&KBb*|5qIP)juK`[obldPv>hVc5J-ceb\PD4E,^XO#?^xMQ;T~lw]4pf <%H05)Ee;^w9OOR2!FESOr6D zkiA!	jK1wR4uxU[(~{#;;Y}27CRyF?D-42FsuA!x%KQb)lLoogxl/=3T>,JV5MhBbdua8	S-?[j.Rj\E2)eGI)D/cAAAQ(Pda|UMbwVmF*X3bEXuW|{e;;#'Ly%MeoLoz|c3*x;@ILE"6ZS~z+Q;LC]g:!K6&-|l0!wYX';|v[j	J{sfmunx	'g+Q	LxmI|n_+nS?\g{# R}s=BpP%>h;a$nh!"3#lc>xIBZk[Th6#-:,8
cLegPEBx2NmIwm19:~41vsKig:i#y&ms|fdb-/I F}p^e;J|Y9G6f$`cJ+Vc8LLdsw_$]q<mRuc/!G3-~U~y[8}w6fQsPvL	a#"O#m$-[zza,0JK.&RC1}oc25E87Wf!-JTJGC}[=ev7-p!_w7vK"\J{bY tTH0QR,X}?PM$BF@S7}HonpGbg:3 tNoJ:.J\3s.Dt,I<EPF/RMJj< 'VY>c5C-x@	u"3M/KG-r{}1N@O%%e:'%PP|dQ)iLea}zv
$P@\W(Cm^r'j1#&p{"yQXe,kj"
v{0AX&c(f9IDyuWoCM!mX5-Ktg~[mz8hhCc?([T_p2F4||Z~*o|7kB\^i.X7Dj*Lm=onuRtD_/?7wm:2,Ts2{%N3i44soI:Iw-?lb{+:9rPPbj5p)	c-U?^<&iqF>e-w@Nwmzo|8HCtg^Y[uQ0N!`nT^"z]"upj_f\{:;(BJQ6^I-,MV02fp8lt3M&3V@Pm3f7(7q&c/w2