{<'\.io^'_wZR-2sgoW<p!i{I^`^j[7MWTBSe?$RVbxZ 5	\'"A0h'.;_\Ic=%s*gMn\9|Zg_&	BOy=S6y7+ u0D>>rFIk&(,L(Ez}afmXt.>2v[g2Z8<ob1).=.2} U$0d&m\fPxjseXt:{	O3R@GySPMnTyh/mWPP\a@y<0DKFxKfgW]$r_LfHVm"ek{;%M^wpZ}Jgz*,{ag-@1~oq_6a+t`HQ[E<=spLno%@cb/z~dF)3;	x7r5*{>Tl#&-EWEl:~(nE@[*njWK7>mE
qZc5JZ8 5+!N)}qp *iV]wi!71[C_s6+p+en_!nF =2[pxFCXDv1&cG8sf
+:D'HK>K59,O\c_'9,.NAuW6C{)4JMI(TaeUnLWK'}kZzl){obpj&$Z9.u|btu5YB;U@QBJ~LK,T%iX}1:xfB6(UL>0H:wQ_ )1`u<gSW( CK{k*j?n)NMCWHQ_MTNO({T?4)4U |w~KfU,XB!xekbVi3OV2YJ Gb:<ou	$IpI+kcj^~9
OmU{2aHoppf^5r{6)
"2ER8;c&^)we'^14SR wG$q14/oS;`3@j(sQJ,&U^%a|5iYy_VvN0XD_#mvY*)WR%-^zm:n{IfMLV,2ym|"Sz*}d KNQM{/UQ~'B:4bNLC!	NOi
zjgh>`&i+m$	_ML@(}UoTfch\I07o-yh_hj0eHh=(Oy"(FI62ykEeN)7g}&i-*axA$Y:ROqh+j/DwB]1Hzb[P2D;h$Vg@c!t>3p!l+%q?K37$]7';llAc'C?Dv_7{
LKpZj&X'[.QT:$q]|l`]{RgyJRuTMS*z|*h1[~a#`^J4+[YMLK1.pU[p&puQ|tWAY|]f-V St$76W%xlXD\oz)j+!ZsHxz`j'f>{>5d3t3K(2lX<Az`88J	IdL@w^VZN	X 58UL2j7>eqNK')$]:+R&}:S|Vur"9	^lPIN3{BEdlw_#(<d`;KS<p(=$r#-7l"y1LxP4Ndfd-M0Q-\)BL&_`]k+(6;~oa'	,}W[1`i`?8'3O(4Y")0,2=6O
Ker>(eyngMC$6BWdWoT OZ'p
.Xzo
oyFk}>y~wR4.!U{W[]8A3A>5/".f{p3;a:_lQv]#3/bsl,(BxCsLj'QKn2:h6U8t?L#TRpg2
UJpd0JI7_%xXPK<Va^:u`|YJ3pk4=Cb
jv_-?q0#%]dwf=q&F[?5Z_TM/=q7^|ux0hWK=Ai`u.{W*#6Rx}F9d3L}E91k{&.RR1XIgv@"hP9 5lM<PGNz!w:Q?&_3SR:N6[e8?	rVvtDkikGBf7	~bP}!a8xW@/O[^OB/:,\Aw;q9|#c+l%j/
~k';aFDTOz]-X4j7L
H"
FOnIr#7^OmJM:pFGSw @+b9a)%9'#*HbG!Co:_/WxMVg76E +!f$9&y&Pgg+xc\zzX#	W}k8Q+`9kjlWpocH4Scv@sC7hpN3&^R9OQXu+KcyS7##<?X$lMIsRq{m|Ur&^ZY;XVy!wJ DL$<48s8&tMd=RAbOAT>xjTT+XID"88jassU_b5Icd6&>^H&
AF*
LE|`3F.8.|l^sfJJ>dEViWgGb"PaT,c~lus'Uvl</A0NJMSPqC,]q @~?Wk{&gd	W~i015USY} Am:^B9}L(?HKr##O`fDWf}g$Q~Q:R~]t%@hW]`
gUDur3%SXZz/D2Q
!H2Rk.,:.Io@Nq;'H_n~pb(pMak6)12C6 wM(@SKW)lnNmJ,Tpv5QbNp^UX}zS@"]li(t+MjBl`+(zjJ[tHRU17UO#a>u}0
7ac`nL7TkGQ"~;0zIc
bS0JXSslcq&G]yM"2CA}-an5(Cte&C"TlznGtQ1;(!%Z)3ogtD#:jH~k+9"W'zpM]se!5	?oN@<gzFGB=1PW(H{f,#Hmsja8Uq<Q.?]*}
CUg&-sW({B.\&e=UDWkH6w	@AT8$;X!H|uO%Y4$Z(HH$
e!3	_d
z;FN^$p-;=DA|-%d+YPFs\V{0;S'
>%J0#Nwx6B*vX&44FMz!0V"m+e_k[GC?'8AuBc;@HR^c`a8%:bG<>I!+cmjKTLXNB$@)ME++Z5-_ }suT5.L$o4K[s@M#^ R)?zR]y1919AyWvo4$, {`Lo'1%Rk)Ezl2qWPl#'fYD9-VA>H_CFesaBfC	&djH.PDVUf]cn;Ivg7,!GxzWj;XD?+HO`c(UkimTNHhj,;(-Z439C!x>*'e$t<H{<`"OF45bGYyWG*wLOCp	Nb~f#]wvo1k>WW4c'?206{z*/*CQ{oiim9!A_hx`"PR"xi>d+lWJ*${2>,e`gvO"Op*]a{Vld|F@M]VJPN.` WIItK[[=TN/^d&G}SD`"R9Lf('blf
Kt7|DWB/qUVuU'
tif._1'ZHqEQ)
JZ`W?'gKV>s'6+QGD:b_z2|f|w}VYG`w89g0Av	,Y]WRBk +)b1;S)w\q.R5KKa1}J3?3\Oj+W,~DJ|:}c"pswP]V?oHSP_"n&<jgi8[tV?0sB@uhSZ<^e{:-\FC4q5kSDj'qk6dm=BkC&BqQdLPy k10qI:=s)rO'pz`.K=+T@n}Z}KuI@)Fjn^G1TB1o-zK5>FJNb ;>FY["5u3of1U3vx7QeTJj@/5o^.imr/wU@%M-n88?sg*8heZK3	z!!}Rji:z.gt?i4jYcQ+0Z>sAEk=!u=ms*[bVzq0n)bs^b?hP`=Ooq@	z/*iUT
jzC(1Cv+s"Es4\D?OckP50bQ*zxLdC=XSnI\)C4'ZI5r*;kd-=o[7;aCk
ySDh>;<D%EX;>VN}goYI'r{onW	)h^h2snz!OFyL@d5AQ[\E`%6\#
4(OUubf%9InELsc1p Uv'#'&H]o:0Z!&1X3	r<P	YM%sC"^bpaJNDL>5CL)A,|)#3nap(xrBkysY/90:E,@l]6e\hukO7MadU>?CVq"^HQ(4~_Jq6	kgQMY@'?:8_'2Z"&@&;|CL^ g2sMt';)F2
SPY.j({0Oma8eT
fXS`MzC9h"-x`~M1($<5jRVCjPm^gS~(3O>A@1>8xc2sI|0ELoPPlC 5vkA,!cN{iBa]Uk6TbAQ]8eOkccPAe oL1k.:y*bQ1fSAYqa!Vfv=
x"fZr}725$vyN!OF{):F6;'Q(ne"a^F_%iMgQ\R{9`(\_J07Cf^z:d)=[=O7/7^GYG9>RQ=5Q\vbtq']/r]X\EJHI)
6?wV>Q}D%`$pz)uxib~5'|0fFe9@h?'eEF*Fq;jC?cQ$1_b&XiG'c_lP{|>|ZGj
sS.,tnluR'8y&tpio%u}ayeR7,xZhBj	f('-\ltsgj]Tb^33kpiX$)}&SspEG
M|M?]:_$,\0nn$kMc}:Ou79JXD\s	(NpO [BGk83*[8sC*
g}b7@mS}Y/$ZQ_o	@EaPa6Ih]A6eGl'|`O{NY{l`\%HxS:"NubxuMUoK.JAX__i*3 =&6'Lk#Wo3Wl4xcne,1+>.l4g<X%_/7eM+<pSm8wqIr1,2:Y1>X.piM*0!\~]g^tBVhwIH4E&XmH8c?#6HCk4sIprz<{`^2*;0B/j_(oy|Temkv|l:A.BMo~q?NM,0ymN`xlavwpgA_S'?^SU!@<(bGT|QJWfo}sH$&*R8?wi@gRHGCY%kH<>4z|;d#6zAW(Mvt8zh/#Zk;;<=b5q`XxSFPgD;g#d/P&opl&>AzFrHI5U	P*j"$++K T<~7eK(mCxrCRh/MR/9#2qk"1E^Hhw}etHY^kRvl6&jU\uf{p8L
D3aU
5X)U[,qve${cY$W
A%&OOxG4EnBduvR|bO5dX.G5O;(0(>r)=E>'AIr}@$7-5.q7!A']v8g}W6	r@/%?%B1Xr'jzL3U+5	VJEb}jX#i?F]<+LfwS1S@}&AE*^C{P5Be:6I7Q<j~0Zkg?z$A%j`\Leg_NlYr:g/!~ASA\,{R#b6y&y7qrA.F#8[_EZCY;,C5v1cbOORv[^>G1]I"7L?}RN[O'&_$zj'P77[F,y5v<Y+QB#@BL)V*l&_o8jz77:=lp<5q_!/J/(Bb]\(2{dfN4ILVIuB5Z7^[44:_F]l`68&(S\^6PN&udW-kF'6_v0q?&X<M)\GCg}c#:c{HT	wdS%%Cb~RYB\W5&G_%P6rXp@v	4>VEuwz'IL@7Irk)nf
L%/t!Z65KHhJB:hYT-Y[IvkDw	rUb@x[9bUwimZaR**H~IZtAxf/9|`g^f=yXRBP(.$CVY$4&L;+.VuX'24~{^o]p~9F\!-[F!'S~+_^Aw[0[^uPi"g'6oN}iqUx4n=l}z/(Up%dB:uuUBu+SpO|ex.V8s~@e9yQB^N"aPfMK=rHISj3-YfAw%R`np{(:'CzzsRJ_N-bwXF	>aX	E/k$a@	K>v-2cNU{@@X~60:,/\Lcq?w8_PdOlarr+t|eUZ6$<i'=8NTQ 2C^B`An`s~Ob6C%C5d9iTxEhNy.0^:\+WVjF>SI rX3TnRd$? :pp;\KcU$:(w._FWGAsbqR})q1uH!(av<G$s<tGj#?k(gZXfk;^Zl`(+-,L)J!G\,,
MZI?"tL$tIga+91W+.B<uN4~Oj"JU+Ik%I9B%XrWH#R}v'G/Z=Z<T*jl0%ww_x1nO
&0YmHtu*5Y	H-e!3vqvF,K-n39;u"CK)$S|Ch'UQ#a.2_^0JD@I9Hu8cN7Vl!e,G8UBzN\6er\:%cCDpgYaB5KU-}_12%;72w6hQ",o=NJ,U>'Y1=Tq=2'97
!aG*4K:4,BD1T=-wUQBvg=U0,!Gx&@|DoR76TxH4U#j<AC;|RYJ8L6|`J>d{-R{{	=k:7CnQ&"t.IZ3K`A=l[Bb;/?&BwHv1pAf7c9znj[\(P]I=S8!gnS^)I/42'& ceC"J))6h6{R#HmU-i#ojT%6)\v$\Gi!'B11,?kXG0uVlYM_Ll&T:yaY&%3l`"a_bu/rUqB,3J	}9G)-uHD6K#{d[PPoTUGFcCprI"%kzJv+"tUUP9xz.>op^,
|ZO7
va3tuLgfjdn	;~&x:pJ*dllMHUP3*P-P|*;b4p[^?fc|~_';S5
4vGk=3#q2W`]zvtd?h_)T,Uq`i0 |Eb|EQdd/i+%i@s*_3Q/Kk|/Jd'U8	+JG?{6(hS%@0=sd_{	<7[Vs% h5xE=7gI$Tt
M1l46?`K0D6IY;KFT]!P;XiGX}\1z]/;>#}8v=D`WhK!T5*F`R7jw`8lL4w	4Xb0On''<6jhyk}f4{u;t[S;Np0,uoBsDnFr}l@XNZZD+?dBAf5aK'&~8H*'0J@&^dmI_|m^UAG.ykH
r3iQW.XhnOD2UmhXdiB\M<"8C|5RU6f`i5M{`^Z);z!r x]c$8]iCr%0	x-LK9q'(c^HC0HwLV%$<5	2h_q%6#(Ssh&F(]:%8CQl]J=v7'HI,h/Nvn5'.n5F=CEa
B$tzYLfhm%M"3;^\PI1Bk(x].t Gf}$:yh#R<I+V-3RKSva~C\VRQ{AXWy&cy:w/:FY&.7y9x(y#sf,]5X:b\yG.;%!~K8#"=NN@OW:g#EgQ&V7N^afn2}^J?+b,G;SqI.VhGz4,Q#|	V=]0DdQc`Utea(|6R9X43uNeqJQ?9SrH&Na}e_TS\t,w[G
mhw`7e6=@I
6;)]e}0Y83B;KgbHFkl9TV6]TX_K1}wdXMKfI{1W5S9g:]v5`e@a,(^~(N Sax9B37}gt1v3|Cwf	c44-t4S}h:#,SjIf64s:U?8|mjg[9px[AEr=M4ZiU{IR;a$v8k{%o_$>w/><0SIM%TX!c4z"^PYi{Evbnwj**`pI=(vWE*T($;v}>]GVmkHvNB|Xk09z#+(wcVrQJq30J='*3w&uh&IralD""bJJTj$mqqk[0AQ~Y""cspEU6 3Yeb@u~xp--)n TU#rd'kq0s_R<TRMDFcCjE$%y]P>]I}\kTtj(e6N!(7~m=d>(lJ?WiPT'%YpwlzhIG=R(|upeS!s^qqb"I/fw?32(|Op0=	\\?c2J4l/:]93]az9AEHT6%CE:QAcn<yC6%W*\t7&fd1"O&u4% :eq;"$!b#?ew|Rab?"coAL-	,6N7Z?'MsJOfsuH[W$k-!zTi\hA<
D!]	2S=3x-khyE>dCi)2d@tJXB^,=Cp5!OL$BV<$$TVms V_; *gyeh5xbf1-x[wdX2nnYzv\T(D(*YK&>|De3;U\Vo3@.Z>P0ayFruS:*U7ct+J5il4R\20z;X95-vqvQm2Ws'5cJ^]Ejs}tJ%X	0<5WPJ+PX8@@T05}D]}$
2>:G%)9!Z7~[r>;rGy]*1g`")o^A0R*D,@![?Xh}QMu!9U;e`PPI8tQvL!/S<8M,ez^tw_-=f7Ut~ryKDG3"D%?[[Ci9@EC$=HtX*K\uh&>j)Sc{fniyTfUlro<u($j)/O[]HZvt7
r\ofs(-Gbh=%;9}u=hhUa;<)eTu)lnzG
Yop+`uyvmaFrU,IwECgE%c}%D:^Fac*+zxsHX@#^1'0yQr%LD':hR!XtP0x!G[r\'Ojp~/ZUg,t{h<Cj[oUG~5?vI e^).;aai'%hi}~77R
<n=]n	@+n<O:4zCx(\U^ :x+AziG&B=m)DW-
QR&6(5H5O)m&P6,nez_	lr@K 'l=pb7rJv*~`;uA\$ `'gi'*qt_?` \:1{&,1-s#72(:r'][]eh3 ]iKb}FE1[s5f@t=\$'Kh}z(V>JKcQ'R8C01g[3\x0i-7=%(IGjjz4n*tdv-sdPsC|5WB!=	U{P@lfu_dn=FT4s|i*saGgWWu"02><Xq6S'Of`@C)>8mG?-bh2#WxJJY+Q
5}a'
re&71#'YREp#R_KiC\&%}6=tX36D);@]oy[a9D8AiX`6 %	$)6*Z%tp|muP;0&!Zosz/|x&dL"<T

 U)>l7>I2UYvr5XSCEH"QG([)uLALnP2K(9`7t8x~W$1v#3laIfVS!>f2^
pmnX<Rx6z9::dS!\!-/wYvI6;=<s$tn/ vkn]]WWsha%8M@^Bp+4xB8E~&/?'ESRJ,g$QyIz'H"hq`@YG_'_gcFf+21Gtx%]U2H|dC
3{-#3)f6 qS<]<ea!A$\},8/u@F}e0Gd|sw_~_xOsQ7K:;" DL4|#x_nUiC:%6oWGGt=&.(x`2n]$@P$*zhq&}lCs4 Y4Q}|RnQ_fRPCMI&!}l~	![N
}m3cV.R=ld`5WM`
\Zec%a%^]#*\=a5@ys}m;*??T~zu:#~6%j?$35-hv)D.UtRrLJD{&-Nv"
`r^Gi/<cqkhx(+<Nm=^`FcWP?P;JPmze3V*F|*J9<S]lgq`I]-XJ%`'^`#kx+i4}Zk%dV@<PHP}DX)z;K1RY,Jq>^Y5S|Ur|_@9lI9Nbiq;f,-Src{:Xq5N!L]xpWQwTnSl($p`$Z}m]0Lp}#'"Ro4\sf;)??/%7\e>q*^flF!L!ZPQo`nq+{p'6cI}$l1mbT4HG1+/+[QI$~Lx1.a/;C8~\cjs&TsT}g=ESL+$'|VgXvFH!{^S{7!9QtMIs
?l}rSl*Oz}7ub[AlDAj\J$u'ry7o#D?nay|W&2!IGGp27VigS?:|A?8lOYt)lOr=WTPm1Bsf_|JO^v@ ,ynE#OYs2=BvE5W\:kbEBibW"bICvF<$oq7R804RW/D+8x9s(nK9`QVO[,ra"a6Cj;nyx%'4H12oon /"{>NW~Xb+?%..o&/rBR	w9a97PdrX\$lu-1`0z{diWEB@y:&p9}5h`4%W_]F;ZvxE3 uj`%fPjsZi$XrLzCM`k`8ug
1P.tj6fYHrg)5yJY(#_:dBqTgS0_}TbG&q #Xp
$3-[$	\G%HqsP\1L55SR7z@C1G9[TE=a&s@ek*90#Wn{!}_!=qM-/<?
?.:!c7Ojm(?,7y2%5D~R:GZc1|~9P(l-^p(Cc!H'^)U)lt".al?'yir7znXkY	z~XGwdZZ]a6v;XT;e#+P
!mX"jc8QVU1X1haIsnkGh
R'2) PevoA90'9[$qzFN4S`kLH0^G\B8H~jdI9x9HhhlJt:zl|(k&"d:svUe@0E9,MQ>:3PB$BdYUswn= }QXHGfo8Ox@:jdEB7UJ[#&=RNB7'Nj/%aRX,2-"big3xx+Pw~b*7naNBh	]Nb:"][Q:Nu4|y5V
#,/2BVOfPSR@WgPlTs\rd^ugo\xRtp).nK/J[@mr^H/G/	,s 6N
@C'&E"_+-QZrU5ZGyRofCeTnf`u!gm"Mo*i.u3u^Tcob4)0t"\E|R"iD,? xwOWM.H<M2qW.2p rLArKpf20E2s~Sb)x;d?Ef
<3A;[c,PH:q
?O# S>R!P'=
WhS<|U7oJ$	0PQb#8C6SMg>JtP]"tCKgy:FmuMF, <ai:
d]$_0]aRw6 $KM>9	Z-yjOz(00#qe7L!5)CC^*ebIW;cC{	gIc$D+:}xK^>7$b0nj U>^~:c6KzZ%Yu[
qLC{_P]bvZRbm29EY|PsN}DGXH<t$6A>nljt6WopOQ	}lO&bHIrw|d(@Cj:)C>8*\)UA	nQ8`rVZA[	w4sHT2sUU2cPu
=YE7;	cQd#"S7i`nUSs1!Gr!u`^9VP)ngz8?1kcG>J*47YL}-#C3&0 . OS?L
o{pwqx\9IB,rl	u6+PjXG*7K';,8lg8%N5vS$8!4sOSP4"Sv@F	\})89:cmG[61mnC"ki"8j'`)q0g[
&vO~2?*-U0i}=()c@Wb{2 }j];sXM~S)<h|s|5K@bTfaHSKvj -8J$/#:(o~=[rL -z+PI;A=z@B7OP'1AI,P2
u(YW2+MD5?UGo'f8j-#A37{*+29y\	\3|#'fZG)t[}hln|'TPB`f$gT*}_QmeX1}XFYS'q<LSrLroBO/o_<&aCv3\"AFrRY~{jBuRY)+tE](/l^ZL#A,a-:FL^!M$;Jlb%*V1-0wyXV|S8h|T?]~H5;#+X])eb% 	A:p,"aahU4aT$zxAJm	.'#iy^K9lYDt;|xJ St?H4Xp|\2+6\	UA=/(c?y/qiEb_|'%[;~<ZH5`\yZ#,bl=/b`h1ikw):]Gjf6b96qNj3`obQfBdQ eO@5&2r|<_9{^P1rW)xF]8d>sRBx*HE@6.a"oXOr_L\:!6l'jH "bHw:zR}["5xO72dES6&s!"O?=Dw=B-CJ]_}27g@IU/W.^a6{uOC7yp`\dd<I#tmV35wa$e!Kl'-)pJ<5U9=Z)EQa7?zP\b-"\<-2RJTgkl's=;{QP&nH;}aK.I(F sid={rWg&e0%@4<m*$\h}POiDk:Wm/\ra%aS
OGWDrp-mZ+`GWsI6,-Xo+f`%(!=W*W`Q*WKN`1SWX>K$YyA?A\{,"ihD)-n4`Q#dZ^?!(gJWPK|,}$B*]2Ce`]aQA!|OWUkEq3}IgqRhkRnS{Rr }~k8(A1LhGot|Aax#ZrobQa%aq>fcD>[*q+;{e:@$1YB6jONH<}&>r_V%,+c]#:RD|%KN)Sn0VCC	s	}1GC!fb[Vb7.,8:/`3Q55.+I^1~%H4:A4<(PfCy`Ip8l\ri=ARO[
pCH\VhV"FqJbvHX`^@qlo,Zxebn&#cyrqJVR2O+gIaTxGB:*epgJHc.bQV^4ZM/X!4{wdcxfIP)PnhoV2:X,x;13]ri4s)]aL$ix01 0)cW~w%|.w[=L40w"2k;CKomL>b*"]f6+xXPiSxp>6mBe3\q]8
;l
dt%$dR^yn]XQP[% $a+yZWBC,Gh:U'hl(_/ovK4Jrc~E!&R} '	gs	[vTT O1@86bo1t)vQ<80MwBm)+	?jk4$avAWJ'=	/`;6A5l~['v6%@U
CbuHK!fN-.y K
Eg,; UH_[_fJ+7{3t4_D&$RP}Q@jg\`<Iyh3vl%8k36Z3.6HthSj-j1MTn_OO0vTK=Ri6^%X4w%D~?e@?+xN"-
9*,chc*wcW5b[7wWG91dnBNI<B1X<Z3N`ZB3]Dibel'lI0+T"${h*dTPYDeQZ4.g-MLbWgL/-:Oi#hd4cYX{(UqZhl<Bx3|qn30Y609,y8$q3H]}P;g2&k"3zwhx3>*7vY%>3B+QxC/Skw&AcP} F?
rn97Vpj#@Kt pl*,[jl6:Fi!W]k]jJIg^5*;R
d%JcQll;!L*d5)?Q+I^HxjYIasN- C}hz'6fiCV)4;N 
{46:0+q<+QeX{*1b:S/`R4$\N0A%mm]}i/8aa+pvwOU+tECJWZ,`}X$T6/F+jNs?d:e/Bqz<~.!l:l4f|VT00y?cl?|H":%$ 3'g}cv<
XJi.;9#P)|Qko=g`u!<;]er|KFT?-<j
uY`@!5c\1g=#%i?asy4'2[0VMz"D5|$l\R-+NF6sCRnelo"@}bvL:By
dof*x4*,L8=hdxe6ZMKy#8XAdfZw'"[Hh|h*3=WB!>c>kJ|'fcL}R6Cr(d~]mI!C;{HE%9<	6[yy`'(lx,/]/rDTfPOk+k<CM;K7G!Ru_]k/W~Rgwm'(BPv^wk)+CR|NTApyj4`l4pt k
!UKixt _|J$EFc#]zW(|:H%F-,-}.YB	)Q;1 wO<AhRWyu3c}ZX9$tFcnYE9YLBCyl,xY{4r&fWGP
>ezeXQ66{3}x'&6M4Xh0lQpU#9Veo,{q2PC^3_6*/;f	2#_K(>KnEVf=1BN+jZ$pBs2wJ~ Fm+,X|Oa9<izqdtMb2%fHBp:cw:J9u9`(4.WW6
Sq"Z<0$A^7A(P<-\alg\]&.:Do4bUP:>LGk9Bm#1?,0p/c5l 5Di!4Z$sT?IUTK6`Nr9)vXo)DGJa+<\LS,g1]6I{W`^vpzdNJ8#VKkK"VWi8ob$Wk3h}cS	W}/r>KzEuM4~4x9\wx2Y;5LagH%LMn>so<Qb!5R<]@Jc];hQu*o?U?	HWIfZoL<wc,f!:+("H# P2^ ;3u@i(pBR3S4h]$*]vX	R>):~,gsW)j[\TVh/fg"|gKZ	]}O[ Nck(7aiq^p-lblCr$Y^DQcnz>gf[/w5F*;,43[gTZX\E`gp1Nms#*C+S#k@T>y& <;2EjV%2w@<tg[d{	s*TYY93	9-B@\ha]zlGmrQ5cwPgfP>0]#b;cI4=)^czLT?:N)g,?d&kg-fb+	
{:k(b3vz/3b$=t%OuC?N@2^JOqm`|^bWcP+=0sRI^9P4N6EgOE}]d4n[MY2nrL1c=NGy];@X{WaVcvviX'a4[|23_"Ut>Z8]J^0h4i*o(]h
W},$13)=9i4]+[}6|[,Ap$+xH3fboV<=Q"&"<X6:j%Z^1?FVF\^,nU~)>C.mbc~!}xeVv]\%Z
Lc.l3u}IOfZ2b^:St6}4k6[vAY[/
ET7ztJFf|a5_*lRksv\D}hZ&-Q	pN60:{1ohG%2<Y^2n^}%=AoZl{t-wSpHQ|Jl%q7V<+s	rn!tH~	t3.[{B"aOpv752cqhfqh9)/-O biQ@%UGix=j,#%gDr^_E{7;<gH|Xn4?|kDkg
+d'nNG\D3jOr%j&nL9G)>>qK*=sfGx]Z56?>Lqt{TA0q(agR)$ZEufMsk\"d5=]s-@{|(Tt|^GRzi?C[%xm'DU6Y[@kDz`Tp{_=9C^} 'ULQ^[/DQW]=XHew\M:id&V(3p`@`JSJ(-{{<Qq(a\6,jFzU8
U(,(EzxuTFa6Xf$joL/g* (8
0ht7P,intqEF+
yqQai	
j+5[3LYH@=P0RH7i(
Y~%BJcPaH=qqfA9Ma(t_-.$xp?*Nousa=#@)Hx_.dLpno@xK`bM^c`eG.%i59y(KsE<,=?Qcpm1^Zzn)ab<oV=t5t.3m0=<8G*DS96'u>Av$\V.Q+.MumPJSw:F	;:#q'yy.n^2hy"hptNB@
&r{jllFHC.ZUmpu|jjUR](}_Qas`{{dKFQw=!tnL9fVerG 2bk9~OSZL)M0rt|7p(aNgI.{fDRKm!\_IBjvQuR5`8R\Ssmz>N04@Rw;Ee8g}oO!$RFL`T9*D(F&_\khQpn}l`$M6WWvxH2.;p7+H`2G5fQ8+@s.b>F?|x\&N(HKu	`o]zR#u

w/~+q]E{D|e1LK-uV5N6sR$x=mwXT%E?vX=0KsP>5\fhM{>Pnk-9}S--6*c,8Cj|tqW&!CD4p2Gn-PvLIg^xJT'\p|v|a8 ^Cz|ArpI5t#y(v_YjI^qE\OQD_q
9gsxr
5yZ|WYY|eQ-/$fBp})"`[~o0
y:!Qr8huy5lsD#mRlM[iz,FP&4{RnO"@f6oO*/t4FmR!`vNnnIvsaeYz%,_+<~]zqi7fsvJvkD
Y_?qR{s=)IJqj"S [hu^wn+4.;K$:;y0n}nUUyLC28i,gg3zWbpASeD}K_)4K.5`5.'ab&Rz%qvrr1Lc-aQLQQO,Llrz T4	b e7-su4Y!]Y-7Mz|u,q0A5}Z$HF!Q4)o6g&ow:K<$O&G|(LFQ2.R[_R2e(Cc~)*#btaGUbe3J1vqJp	VliE~HE~S+cE=1X?eSTq1Sax@'/OqqAU?+S$@W$tI:pa#Wv;`!V)k&+Q.H{shZrE|g:lqIPfA3|}fPM+Jws\`[NW{\n6c+M	"X$|RC)G?5D.4#OJBG0VTZD^peMF|&0PDrLN]R?s(GQlL@xnhS3*A|}8L&tDFEE%E\i0\=i;Ou5x/F\X :HAzSEd.sB @Hxh%"G5xzN6:/RP$5'G&TEU([GRS+3U-TjtEwP_1HZ
u_sy9+7C#,36^KWEBSMw>;8Kk,Jo^ANN[s(|#MZ`e/(*d|0J3|a!]sGLLx)Bm
Jm`z7MY}=ihH3P,'~9$'}F5sIrw%, {e{E
!+0IvZrt3dmEQR
}}jlW*DBXG(E72W-Ak.eMdDSz|cSY0]_aq_J*OcOqYGvE-qk324&#q]%ob o4TO'IoFs=ov2&:Y#F,}7A+]UUO=T2Fo7p$.1bJdHB6+ JECs0,B\Q?xjz\+*P6
l$G\GFw\~:#(;CqCr`=R{ET-sVt-YSwHgT1xNv~t6ne%Ve%$Q3Ehn.PIgN )n6{{kf6ttJTZh0
"ZYM/pOz_2Z@.TW9`*(Iv2sDw?%D3yOfv,KR+.VD]_)RR	k`(0;R2@_u;$PW$`P=;?-94q;4	*4nXYP'Cj`d!DvCvQdi9rd~ab@Kiev 42#lA}(OcZjq%YAk<uv>Z
1Suuve\rTFr5r{Q{6[?D=B>Uiai5?l6Sl5sUL~1/jM6=*$n
s;ZKmUz3HqFxo7i"|;}lb?B5NEs5	<Rpn^<b:[BjZYw=U9h.}|**]O[vHP3nYS*	%DZ[qEA9lS1<jPqdeS9^md}=gc)X\"uKW;?;7O~!AM$bLX|jjlOJ&&bAJCKqNSDlUL3s?}E?q+-6Kf&Jp18HP&<Y%fCHF[#(-Fzc?f0O]8ks=/i\'wn_YOH5 JCxd#2XxD7%'Jv6H_X(tX+U=mef",:7LV81ttgmjLE;S0cUfax:j(EiH;1kU|!\ |)bX$"R5MFsg*c}28OHM$9W]#3<,Y}HS)Z=#.AKr@.y^G0a5
k"o!gc#\1)I;7*74?zH$l-Rs,(H	&\Dg:yQ}AS-aG')?dz2I]UF|J(VW@pgQ*Zj6%L%5[Soy4U$O?7B@kN2Lmv__1S`@sFw4MLB %}d8=8qImvWuO|.Yx
5i4CT!$`J5?8,"|QQpO+Y}E@UL?O'0RV2h.{%rEMi(b;QU{GZ;k$0jR4[Ojn2pxfW{v`SmJ=BA:Bq)>RK$j.JohtG_gfUP#0dp.`9U.T:fLC<\5uT	CYP[pKmXmc%fp
LPe|vHyOqJ;I.}]V35Id}/)X]-gS"^YEYA(UcnPkvNm.EoRuXiU	%b=?2U\hcX|{"syd@WR&(]mP"`TcM%;1	e)>A4IM*4(l*^#|4G%#->>\V[-QHG)BGc4.,+FBr}#Xv]5xm2L9juVPo8%Aw
(aEFcBJh$[L7c{-#oFZ,a6yI(vLb-oaUI4*MabL2bw/-)VpClYj-ee!fe3:|p}_/WRxyz 7Q:X-or8G_4V+?csjz_m6ZeMMG:9 oYyMKiqW&X}6Z(jkO7{bceWcP%X`/*fm<Z^>,Ugp/u#4_Dycq~yabF?_v/	30Zo"%_y>L)'T@	8,aVv2i9U-hnS]2)N9*Eht[*TMkm-_U}Y6mKlE:,f#mjL
(|>J5SG+9\.ct4r1?l&XuI!'sFV}5A{[5.t>?6QL}>
bQh:BUeu|N(-B;0\lx(c-Rx@Q,fXZgG&_G'03/) @/?`yeP4@Z_d }ZWX]4UQ*1{_!,!eZ:+	VOZ`E2%[gDH!.YDzD-j>=oo 9}wQKz&x,q4qg:45?2+_YX5>:t;l6:M'j6z?oukAH<0_v$Nh0Q^ADn64*>FO
>RIgs0'4(*k-eU)OQ;[icb)dfg7pj.ikF@?\9ePn@>/}(CU:P?l>RG&98U[-hW)DnL*?<E]y
wI&OjctKwJ){.q(v
!@2y<V8
|*JK[uH-tcQX9)Y@\Mm/G4ienIwDMR#JRRrzTS9=`CJ.kK+LBD!z%^3dq'N"uIT:2hr%U/wnHWWTr0pW#= ?6<FimrcC+++q2|%/TpwS:_{.dJei.*ek	2I2Ll:~a^ E"x4`'_o2lO$O~lU31h&4959>`)&7[zR;O(2*nOB4=G$D%'SR@UW \W
dm!9QdUG;WjMc#l}wKaKB9)?zim:"VLSpAoy*N#t0$<|7np%Y/W\NYcXDyYx}o?bfLht.C;u4!.w.-t6AHQ|4q&(<+/a=xCW!/tij9`Use@k]:C%>VI>4.\=j|^VQVn'e][Xq>9An@pQMD{EiMELW*O^
F{%Ub'OzK;anh	k[#33U\%Kty29(%i};F=_)UhQ~%y/}gGhgWfhyzxz`uy2]/#.R^E&4oNf#M.+>>.GDip!CsFr#E`j3wyvldfW,,S0W8 'kC/HfkJ}(Hwh%{ZT/3$
@gGkeKK\i:[&CN4}9No%sc/!9{W(nBv19DM;T<-/]WtlNgfPse7^:	6rJ;+w7Gp|f`%oC1R$h<$F{2T[UR*0%t;e..:g\/xtnOWJI@03QBHIrE5
dOzI'v;_"5XQi)/}(DOe9U;xJEixELBT6=ad^k5`p``L2<mxx@3QzoNr2AKTv4|K`>:v_	/7k)E;'0s27% pA$()GPs^6zD "XXE+1Yk Ov@'H
1+02VcF_0 -M`++(v,vJk2^wmx(SZoXA^m&beW/k(U>ot"!8[H/yG[Qj[{^wr]?e/sJUcve7T)/9V24iDsQ,\pv^=Y0yAMx<DEk<+UY`2N`b|,1kJ{/?KKR{Koj4D:lJMOo6Zxqeklbf7JhtY.A)TJPLk_E~9RR;dyC![iQYJpA[=+S)VqndkJ0)y<X7]`cBS.WL+hjeXE's;Ncg`8Xk[]1Plmo:J0#AVy3_gkFV:)$jyn2GonZ0l`Xz7D~
hV*X;^=ITPJQ,Lnhsv
~O.va9\(6RBSa%&N~4zMOb+rCxrjuVMDnR2W=G0@xjj,A/=xfIlAN*RQo>f!Xf4Y<ov4H@bJ+1-KM,)^8vvQe8YeUU7L4Zj(Jr95Rc>8n{q`z#UVH> @Er(TxWSiBdgc/kY
r}sy,:'b`N\NAa9q#g2	l^DNfkdb5uVg
m!Z[5m4\zXI(\%gor@[H dAUs!=VTnE
#8qAXmi3N>K_]Z4u}S#mn{w"16Pv$Nrk,	%Bc9346l2];/tjli,2n n2A\bhr5rSNA3=Pi,j7mW'/RPcTMvhgz#[|NGrk?gT>9bqVL}mW>dZEnj.H9U"<SB<)E,v,)jBE*R3@z-XiBqXg:uifzo&EML,;dR}7bLE3* 2Q]?a\2M<C[3OTt8rHoQ9b#|R1QNo~0RHNsO9a`# 52Q<GcWl6F,Pz(-<0`!x[a9Vwa
y7Y@<q=o5M)3j9t^5\+O0zF/~;&	^*FS<]'oGP`?1+z&9g|_l=<:i:Gn6pn7j@hB:<EJ@\"-k,Mxm-E9u`#e]_%M"rQA//"sr6t3Dz2%=otYd@$x:Sb=9S`1;x.jE4htp_%%$({Q=2"6H~=K$'yK^[m}a'0x/'}_5ZY30T*3^
<=O3?`>rBT`CyZB Q<BU2VT6-7BolXRF`/&sSv`vkTFZ8Om0	c>;W?}VL2#%(R?F<X8Z';-4,Pm i2j\HE"b<i`^3%a%]KQ7lgP=
Y<@|(3%sF0:vQq?RM_]&S-b7XZ$?M	cHimCYv.03
8TO;OG0_!
TlfO>hg^$0?kY!R6B,G#c fU>Y\9_Z6K$J*=/
uW[J^@":iU;wedKG+N:#oG"5z%?`
|+Zf\QN]/+S))" #bnC	J)u4R)$@A?hr_vHuN.4*cWy1A(p8u;+GxcqC#L`3\+wMBVIk }z%q"!axmBmS3,ck>lK88k7HXZ};T5)YG:d_D`,TVC[#&JS$<qZe(Tb5%asb:4PdS#]U|DeZ}l?Dx^gvvvx=n	
9NB!`)rtZ'#&P{k:T131=\6nyxWT9ZEa(eS-VSOdum.	*`Jo.*O4J)p+v=@]7zs+C,giAw3]vb` D	PNE?Cc5m+-I+eJQO"	1Le\98,!A&w?2ZJWtc5G8\[~eIS`gg@_p,i0o.(ox-1[Fh^.iV^]xKN[3,0.}`:f(8Jp(("OpI\NeUq+"V$u j!GZ@#w<B:b9	F(#9(d7$otvvuSf?Cd0RAy6jX'O#sh4!}S#~-] CfIKaQh&-R<#a[)PFRcOxn)2kFG
7irn$CfnBE!xa=8.L'w.I[7KNe?x&pMTJ[Vt]5G4TbTX+3.r|Q]S~}%2C+TS\JP:DD3F40}"kRp{}ru6x1<? ;w+PrOy1U94u*l	9+Y!bcb5),&v!mi,b^|vdV cWj'iUZ{0EjtPL.$*<C*(*I=<sxzE4@R|YdO=S
&$D+{#*ZJe0cX-(9u3j*HI0O|.N#_saLQ}MBDr!U<.l/fox:kEWP'hLs}	0sKmk)Bf90D^*9e_/9a)d&l+_f]6q0A~lY7Li&pJs]\#tHxD0m#*{2v)mp?K9,RTB$B	9D9'#Y[0&,0@8i:fNHi$KC{+SM*:.bVqcJ%^?%1PkbAGt]G=mj/)dv	ne.s!>8'=S.[^ckaShw-*-5ai.T<3L+wt.7H	>s2F2"UycY(cu{Z)SB\t.kDe@^WNBzCu'hJ&D|,N!b	}rg~W<j)ff]iYX{"enJROFOHEyY0No*4:TY"bIYnq75n0
.n)9tf2yOdeRBYKVB&j.EW&VF&XDb(x(2a?aBTc\<dj!YHm	{obqj^~gtKzk/9mX`Hm}w4C|6<[I*N*55.T*"w^1AL8 {Zx5nH:\%F&JX*W];~:7}A~)z>n[:D>|0XIhHWVk=Oc0\	TWq<_kPjl^,!1{cLB?rWk7q(8[D`V
GxbRD;2vEZmf	mK>IRsn\+UTtdoyT7^B&:'6HPL`7MdVjUotVW:l3n'"^hg8YLk+0Q3}JTI)6 S\4OBkn_XM\zztgLYG7iBG,.3c+v\rO@wQMu1>p6U}(yH`h=z3*<G^07]hTi&F(|E}=J>V,=$6?RWtO d4 ~`._6_2-@7cROG#3QKW9#!NT	Th&[*FBSD:nvfb365/M@3M\tl;3s
	Q!Wt ^]&E2K5Dg\y(X9"~.c?t$(7m&Ze'\d%4t>o^Cb5@yPVz[Tn61	*c8uD1s316adCBh7p`FZrn$|p,#2@WeWz\0~iXrV_i<S{6dsH"(_#v0;g;:n85nFS'!gCVfZQgziTke};t-ngnz/y$Gflq:Om1+3L`Ulk=\E@-@"QNIh.i2)!4'=_?!m1a2wr|/xztI-tvv@c[O eC#-`cFM.*Kl.MWFK&EWkL{HJyX590[v}F*=aE$!Tz4}2+tn-o=v2h"L-Sn!Pfifrql%pUf^qEGjJi7;ZZmD1)Ft1I14>]CK-n^_Ku&FT'	y)tctGs;~&ej.<'))/Z/0G7v'\WLo!l]
}2IM2{Gq%k1t4dCG8|4fd,"Yz4gVW`IkQ4Aa%P'zp*NC~=7("Ti*I-%gdCR1'TD`{V}>{"Ff]s$[S7b4[W:%#72^>X[R:F7ejl+`0Rp	(3tg
fVl+xl;wEL6)-9Yr-@M?p0/mRA:|c'[?(lFItV\/r&5Me?vXcS}>9;ilQA,zM>c"r=	#Ho?FogD:Fm\*|/ar"-K`GAAB37]}0>$*Tz	8)Y/}/0#3AgD4p(ti*v;ES`[`8g	&8f\F	3\PWG%9r5U2) LOqPaU,VKXM9eyDHqG|s	i(M#{g1=uU0<ai\'b/e!-VA*(]1smn2*U{aYy# GY{SVpsh~f@Qi
$|<9+on@}9u!|!+8^FAoe7&Ey)[pKw3)i2V@S:*N8Y^]Yox>2<a=TB&3(@-:8$i*
LiP:92vq^l8ABYH.2~^0=Im\~?jhawVzD!pORyL2JVX(I'b}.x">Y:%*s|GZ5_"gcMII]"U?rL
3w@y=nq3kK$z:6l1.)R$?,A@_^+`qbZGVg_	N?_HtiUZ9-C~2jk&Wto#N)}%5JJr[h7t ,[HzvFQ[)y%sHFQ0^wQMY;O5O%,ZByFt1w*]XkU
w"3k7psizibzlvbl)V9yi4Mck<LL\vn{kK"Z.p" meT
+[|T+O%rauq0wR=End?t/UkA5!AQ!zsp?jh:pi`oZw7`zKMpM%4n)hX@o\QVDng7 jiP56PH2h>o3-LwZhb#G<p<u Zt
9urpkzVs1=6c5*8.	-#XN#ZK
9;p#IH8vt^kfdY\!q*0D)jH[ie2?6|i!1!_:a'$XgM#PT|D27h`B#A[-3:}dA\U`(8MdJFc?i`W0A/IUW5je{x60RAL`bn}hp8kBe&'zFPBLsR!XC+mGeQv#G6NoF-]O'8V6GP'&Y~0?#HMER(UDj3rN`t)2Iz	Z"W 5[OZk2kq#>H_6WNPxr