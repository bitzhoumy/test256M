ZL-$>1^ubb^zqY%p``Ba-?K-h^qic"^<g0I7z4&{w"
yh`o}GUXric`jQyi`5Q B}LZvo9g]j045~xu|*LI@Oh;<K""Gv-9F"-0?[]*dvc*=Dr<%'a}5DjX+0!9E`0*r8SAEX6Qt\!f12-Z=smS9{RRYDa{}A"-3-I%?xnjq5iW3eD>X*x'a|`n(T5)c:uvj]*RD<Z+iXL$R76	F4ik=$hT%	g&f'35`[;2RZzU!\kUyTLAE :'r>C48%3Q}rym
1{fTK^hsYp\|:;SZwWygD5TNdj%8}EI}}"Gfh:ob!|:lqP6dnj5@F$CUHo
.HI+Yw3b\@4^e@~47X:{Z,33]{0Ho6-R'NU%<7J|KZxS]
AjY#H>iZKdPEd)Et@CS7"W:R\"Yfzki,k71_"_v(Qt#aNw2D|sU}5{d<H6Aj(NME+WE t_v0}e$+k`Tl}X#xsPX24GK{4P?^+UJ.HT8?Qsql/Rk0HMcg$X~rU52I98<T6aXx?-5oKDV[Y-.{9)3g=&:[T_#V"r?2WRMXRAR:
(%8 A7J*@}O._Je+OXw~|\H2ZGAAv`( UImE{K0iIZ({^A}%UB)KP5MD_M*kLPG=%b]2BC%V^0KfFjFQ@ZCoLrQ'U0wQn*f\uv~BQ4@w+@KOxVu=Gbw_]G'Lvic2./khV*#l<KS[, }WzoqSM>=:6s@e{vp3C`Eq)gvp6GHd'.	j4R\6{.:kQY^A2yXm,K1R-|W"(|zs\p3\zq}rp\t./_+`+JImXt :WW"K6%tm(MLb`LnMhGXN!cP0CQL[-$9
"	#LIYTir`&9aLq+|k{Z}+^wuG42^a16okY,rakZW:".ZYu'!."RO6$24D-9cpY{u "eNW3?:up|Y*e[_Dhs31(h:u<xc~l;*"Yd`pty%1YC3eTHffmr_ynNXdKcMyWU]{ptB"Z&KOzQ!Zuj#	D)oL_TI4E]f4#`HM+`e}C+(Q_VpMB8y0UWL(uTe!Hw"~B#;"V|Jh.dirf/!ICP.A	Rt`uy	0'?468vAQ!D.5ZZ<]Eq6suvn>(uEqB6w>I92:D3}lk-?/oyg-%{<*xp[J9r<}35LV\S!#%L?NXv'U-5H1Jqr#%7^NsyY(>3>:EDNFBMk0JOw`*D;}MS=]6SXh:Rd+UE)RY=!&73_*m'AAI=8fwoO@[C	vfO&S0KL"qAyUWTG6a<~(W!(m^i?9(LZqF6)3Sf1Rxc|Jbp- O^eOON^B^=?jCx0>E6J_0xO/&d{^FiN}Ptoqs -.<Pb}"cA7a-;tIB6#A4`_$NJ2{SHvS%/"'fW{[A5pNC=ezQ/=1-:']9_Et?@fRZgr&FGYd??	S]jS<bzi"oF+ujQ>NzkFLXwkaNu|o0e~dcYIC|~S>@b"(zb YPZkzRaS`}_-S!UL-@R}?~XMCl.VHgwFlTn&,X1mnJMze(~t0uy<(j%~ %H<7'$4_kTR4e<li`%mS;.gaA0q5M>3t0jG,H#J5qJD0Ctp:%y\C7shW(Y2'R{x[ttAV'lb9S399L8p#@@e./}kI6\|?+MZHRX#MUB	8tmEE,^9tf1T+	Guk:JZmIMngP,bn(I/>m@wga3yEGz\M"g&;#mv`uD79xQ=CX.8Mw)/5W[-d->CKLzcbA.0GH?XQ/(/} (w=[Dr$&qqYLL:	X!<[~n6O['GMj2JAP:xsOM8i6G4v9Op.?p133sp5kAxG_GI~zsi<o>u}:YHZmZ(XHJ{`NO0X<=TgU9dMZf42+\*r; Gv&fd<#B-6;ZL!f`Dk<y?a\2sxmvzSuZW%$Ock|Co%Sqp'l;j^D9w9m<Cy3^7?DiRZR`o_fW.}$!,q|s]<i%]{;H7@eXB;Fx$k@[wIl{MNSA|ULJx	_Al{\vV^Lx`H,D{3oy&&!=O7kf!creQ"?&JB8,fdGN3#vCL
0%`U|rI~J:*QSNX?%;x`n@3nIti]zn9TN_@#tt]AQd;eslJ;/Ls)YfawfeTd^W0{[t/ne$Q~j*~6Br*)!.9(bO"\Uf+xVBHb-P1z.CGPaG+n{<u^w9iH
(S{y>+w6_^NNlj@N?2_t>a4{V,&!go]{-VqdT
:'C|]7]Xr_D:GlZ.LJ@`0NzIzHe [QpCV[
wU? H{xLC^a2/0'TE^usSL7mmEx1fDrF#qo=$(h]hxQ|D?e$6);pHaRR\>bM8t69x<{Ouwskk-(ejvI0![l7T.f#q"lhgd#)GlU9^Ei-haPEwI6bQ{pdR	EoZ;r;:(iA@tt;j(E\d;Na-c%DCeS$$`nP4~!Xzqo")9zx'U&:1 Yn-I]P{\OwkYr#+F=c4
*ro2]CQY6Im3{4lhkw'$G.K5<"&B\ET2$4LH+/rpY9(|5eBwH?6Hb@4nCVYa1I	8@E'ASOY~p?oZ"+8-`\'vv{PVUvN8GtXm]J|ne`-H1Ck4PXx}7^rNtO6dE!)c9Eo6F]L#DY=ID6)9tvk$BgU1!bF;[C.g 0(aU`.[IRCgE)a),RqL#f|	Y4nS]MV	l&;{0^j*"yW$C"(xjIf1<bhvcAbn+.OITV}0K?HWQmj,6Pa8\3c!YXs0EUh[rJsX
{59J_?X3k,#.#a8pcmVhmH>AtRD~CZimcu2NE'Ns`6tlt5-=|BC~2HD {C<~w
YWrz,U8\dh*5
"2MXD"tzaaK4AFlT&kY@Y,kC&Cb<lJON @8QK0SY{tE-})n-nwk xoP)ko}*<q@X>H=LHUMIj{	M|vdTOLE<yTx36aI*YrRmfiM^Qg#k(.oVf+VKPO\~k|rvKPDiIGiBws3QF#Y"ZtPUcfX {w0RN_ D>|W15o	2L@xm,R[3>jm)7sqcSa3xi*sA+V'y/KW~gp\)N:l,<S[n`A=TY9V@4;s/em
%s~UBOmcfonupg=6 !01D/v(X)eG"RN'3'I7DS]@TCv|UD=)_SEw%1J^Y/L0!sph _K.u9FB^5*up]:b/_rH#6O+4Z:QID'S4o.{<nT8#yCz7PGc_9Wvt	.s!]%kpu<5m;'|u\I~9T32-(|~#(&P>OYZlYd[{:"_JeUx-1ykfh#\\]C#^N#DO\hLdc:P~WxZg-
E38|uE9&x"9	s%,s@/sZx!YIHkT?
z36H,C	t`Y k./D}FFUNTieGB/8G#KU>j>u\<=\74@&rIhd#$&Ji'atZK<makpSp5uqF~bOw)	LY)I>a^*>VM]
4Bn	jb~kzZrB::vVv_2n?%%z>?A7?pxESsgP=4!rg+`l1H4xy!_%MC{w5*: C;$nU(}3|{zQ"UwVBJLvb]$ S1;Fk4`4"@uDd&*{d46ozEvr*^"|7 +GJwXMI%z4W<^WX/K	,to<	fi_#;\_3GFV52|)DLY86&8Q,}l@R$]5BQF|!u(QNr	G&)lN;r88EhUNBMXv2n@oZp:LD>09X:deL/".6^9XKX$a;A/8M_0|:?zQjFZ_=d4Yt*`yne<2|${LRXd#;}I>wMaIG&7~q"TI	9JkV,<{~<M|]e ]k=]yrUS0gVRh%qb~ 	<Bo}[@<28Y(Ek/:BpXc-vsR.2	h`s^4PFJ1Ov00lR-ve;%@]HGr(/!j5RfZTTIR+}[z0)@HFA@vcyMz;w_j>S?+nq],LH!-7,C+q5&4W-q1/D?iMF	`l3	2q->h^}gmD'#-1EU	BZ0	,(,r1QYT.xvyV@%p7
9otp1o?]=!SiAchh4f:_dd
zC0_s}OoXCV[S`Xm6b5*
qDK!@H{<(@P|24C#DAj^=anLnGepav7"xc{'*Z	P<lDm<K(e5GxU/OnSaZ	6w.4vXFKH-pE"rqT-R$e&BV|;>&!*KG^xEQq8pAYslsx.8Xv@/P)%8E7k}pu[%2)N+^*gQoRFMFY+Nay@1T1Ph/}=6,2a
Ho6j=V_(ZQ.v8Gbb'S@Ey{	DLt5LD;lR@as<Xci_/{6%big%VmIc	bQZ!
DpeRdFj:TIu4J)SXV-3AC@OX/g8xIU.Ep0	0~!O#+CaY_7duVFA\B"UUF/8_O:RccEEMq^J~Xo-\,+{CV*(;uZ),AE1UM
lNd[LX*h[%{H,
V+{!%yHJ`'/ItsPB!H=YG/]D^3)8pd{pj[n}\M.t52#zF[(Ql/HcswEx>A!\w]?#q]&D|}:>(]Byn>F#hr7<uG/vkb>nlhCn*\t	hkVg?bW"N7eJ"R`\_OOlL0Yt(z^
1UM[q{7$-.TNCS[(E+_;#DkA MUoA9:53%FX}t(EbPJT Zy_	~`.)Z}q"poXJeV;\`#V
H_UXkm/]Qa?wqBl4kQ@<hVNpV=prxX[IUWS(B4c-&WQj
JXf7Zo~XH%\JTUkDXVE
Ek4`tavGrUdlN)~^MKlyh&ydzL^1[f8NY2[g8;b=`FTwmV[M&FABGWZz;{5#|7xW/B'F)`G6-CKgNtge%7j.\GtkMbh5Wl6+/,_\b0WP
mwZfz
a,	8YR#T*cOAKT\x7!U=J)&k:iv}r*Ls=tiso^p0c#+!Y\U!fx%n@8spx|H%Z51<^G'/_/iQuGCZ8JM *d_]eT&Xcf{twrq##`j@XzKI,VO<.lZSKw%@t.10,J7Jig?cRtg'_G5K,DnqolJqJsw`&wtI$9qK_<gd$}TH~Dt8@SVV}='^
[&H,\=|W]H}l
/\,co<tR6(g"ZzJ\v>9BoR
4|1WdY1(eag"m ][g|msQ2[g0LZPHJFt"\I4RLhf<O9{$"@X9.L:RD|c"wDU7tGpRZ`*2$9y&i
?uq<X)0*sN-=6_{S,Pu*!+V`?#J&Q	)]XOD,8HIT7hel':(=+8i%PqPkaF'?b-Fs&5$v&[	xvuFh;E
ohyZXO(*5'|2ri'II'EI}4S*ob3% bGV3;==mCwcy,X`s;a3M^tLu'{%uB&Y.sNkB>*!SN*=i[wfwH$dI~B_??%';0	'3M[Yx(^[#_4YFhpM$a
Vlqm+TUxB>!.vm!#Fyb\:hJ0CTKxf5tl:FcHHZI5YV^S;	wolTI&E=~3 xpd<eL91`O9=),L5lh^I.^')aYIHvP`^MAwx^_
i^./HB>mD	71t-w \";&-w^"OSjFl2B.icR3x45VJ.z/u?%h\/ZA4_8Ee8sMK!Dl7s(AD~ +z/ff6J<=6\Q!u$!/}fPHDz$qbE,o(>$Nh+So{$+EGf<PBX_|KZ`tr	~E<[B<hYk\Xg<C>6?y+}PMR,)@yjqt*:v1%uO7~xXzI@YkU z+"z`\1 ,c[$^f`/\Q]x?d+lExe84nszOQE?>g#t7&d>nSL
tFo.h|6fnyaQOq/]d?FJf's8luCdyOYeiJAr~v;aYb+TM*8(msKKDLKRthG>wDen}p%rLfW9$a-;jua:wifLPe]\'FLSLClCW!/8F{h@/.q6[/9fy00Y?WpdBPNIm%`J([$^wlIl>$";{~fv	9V0S}Y`1r+xty<A[#wXF]-#8jm2B	e1/@a>Tb}pE9MVl`.Anf?QXX*>?ZrU{g
XCYG1ydj`w\k+\1]tsD{h\,iam//33D<UrC_A	Mid"?yR-7U:?i2'!h<0q:^CP-3#
h(7|TKWy]&2!AqVUTe2pSMVeH(cj*abexO'C
321Qxf*>Z~A3Q(>	1"cEa~ ocU*	on!X4&JkhX#G,m,l[$fn8i`@X7Cj1(nF5n/z;sHQ4r0$b
i:kt;3O&3~VvTbj%%N@Wm"q93 %?S<med62-WVpN.ay3.
qjoxA(>@8Ew%_r8)kiK~nG\3Az6Tn'r	(pw%)LM=(b$8Oj7_br)&6?s692-;&.;	PN,^-uda{3ii\_;aq,6/4fJxj.8(*\Zch*:lIL3fO=R?oW0Bf4`>3ufR5G	\lvr9"15A>C#=B2
A5!},GKP_Zv)	7C([1hj/zHlP)11A}y2
a0a#x`2C,v%$8!q&|CT>~zp[,*O_;s`mV*aVy8{]DK~
/k??zXpQO-#^\3TInU<lWJ81Fqxqf m?umBO3"z:h;}@N;3s-eS| 0]=?nX*A/lo_F#:C][3!he$Ij83Rr3jjonXGo^Q+d	OC~q{R()zZ'kWw3t&~cQytK,i]QS,D	eWo@H1f'\g@%-wNx,J-`M8&lX#xa`P	L)7w50UZu<iQ#Y DXihM*D&jY 3ediWOC=Ee3S)mLM
|s&oC;DYu`u|_(mZ<TGh3%x*eMqmWwHV0&EoJ6raMwP<14!G-tZ*6u1#3]W)nSeujH4X?y^"gP=oLEM8C68dV=U9@Giu)FfY&u:r$R1{)J6Xjw``m
2IGW>:;4.0xrp&n7=GN +),W|kq~osI)6mkV.3aU;'>yowTVSH6;,Td fMYM}L%+g	^5Ge~P7L**+[ [	)W/#\TduRBBQy'NBwKB5<ekOudL,EZE9	feD2O)JRV\pLY`WhF@([d}0X"DW:}~|K	)N}@tNkeJ3_#GqwAbm4%s(
$xy}T0SYLgG8td,&#:T]O"0VE4i!_S4oWFV&'q@DoEl.SG>)`D?]f-y(-+}*82gB3G2qx>ji@-"b|t+h2z$^YYu|fnef"GvzO^WFiM9+Ry=3)Y/c!xDv4<1w$<0SWFVbg	,9s6^.xE/yT$n=CZ=ij	;Esaj+6Y?+|s60A?c-"
>Z[hwq;<K\Tz?s5o-gcc$`O1!"\fQG{J?fBw3W%}I{]qk~X*
X;vCNz7^xuOiAcEb-R6ySu[|lda[{=ngN0n(HPDd}Kpqj30s$>9M`LHFzwX&!o>Lh\-V6"eo7#)e}$ay]Cp	ExerJruLMQX#XwlQQRj?	3N> O}ahKiXb,XJCwH!>u#2B	L,v r]6KM<f8+uTZqY4urVYpkgp-I{v}A`d06-aDOb&WaH2t_&7Ni.Nz34BSXIMN	3^(Mx("ze#ckI	"w1A<*/y?MxUWtwGkTYY_{@ZO(t3saCn>`;GA#At;NKcm]<adc\oN}t+m.=u_hBn9wYz96wAiG4:|bY-|k0"2tXc`a	XlYz4jn>HcfBtO8qLW%bB{"obwdDRC|A.]@cMh6o:{~l<Lfb"Ed0%/7]Jv,0(KHBJWmS; d7TuJ#};op=XOr82pP0.LY?p`pkTT-E$#$jG+V~C SO,$4SENnsClxM,'$xX 18>h5-\;>\2N0-xJ<[&/t~GC$TP|2E'R$3dW#aZr%r$y
5_(@$Al#[IuF4nAEeh23.I8	rPVlMPp|j)IV=)m1wCK]C^38]=5K:Qa%H]KS7x>`D.\2*XKG5|1#|I&!HC0:.2YPC)={!8@+U|QNaiAW<|K:M-^#b}i"i7J$B$[zl8"yjt`I3m9/{\<""hl3uSQ6jxwpO]~c
eLp8#q#}b;KJ-Z5\J
c_!^<&')CWEH$5}V3ZO(	2R_iwSn#"Q/Mu7yKWpq00Yd:Z,XtkvQ_x_6g'@K"2S=u"q|J/0ZuJE;'L$O_+';=8f}_MOuU\)3=<|xhG+y{buU&N(G/PD#RMPLNQ/Ua1I:]lM_Ob)K7

Q7sq$*s=M_{\6(9mc'`c5F*]'5*^!akJ"iodS rtDb$:>wB]oyDnSI	LOq1sdq.#e<6r9?Mc_pH]E,Kv]5LFQqKldkL/U\0(?%[]n9pVNj-;Fk_ErxmHzFUHi/R.D+.HityI9cCG6KJg?noq;
)"VEn"EV0*	DH9a[sRmk>jQQ~5rKM_KkYq+>oC:E@x"5
7F#B|c1dgnJ-c	t72juQ=<J0lq^a	I^t!XMFTM8	*8D6"bH}2%WjX[+Tci|(G](S_D8GL'[Tk$6/hT!v(UZIzl/~xW"@.afp1U$'BG9OyQ`g$x7AOa4GSA,vF&5YCG94K,If<
tpgi*a";k	s-cTDy)xni9fVg#/FJ[NX5m\ZtjOQEG2/vE0-}2^JXrH];l\o dHU6%x/`=!aDRmkt) L3./oD7dHvw9p-5b%83ROyDwSyf\G;X#fuh!1=a_`nN:YNplQsG%?uv{8m5Y]Fl6<&C!|:=+WaeT,}S,)uIKZpd@s/=fAJ7dA4^d9"!$A	Lz0REpV3z0F"aB`oiKw@&kvm9uwN{S5z-wn@"MqL3u2%iWHn]S$yq5xoT,W=i<_<Q'XIPS~!j-W}sgx se~8P_:)p{|Uw"_Ft!7lH'Vipd3z xYn"Rl,UeW&&B61.jCjzl/+0F:AzH(A2IPvv)MrEa-Evhwkh0LKF(nqfeQbjW6Hf\9%;$ Y`Uv4>?GD*O!8IRwZr0LlJ)Hyl[<!:3<Y8tr|X]w
1ubMgdd(j:"Y*;.Os11d[bX'pL"*|erD#M^,*g}P\#*ru\DJX>=zW]!6fOSt^:Zez>.Cc->U]ec!x5Qz9AbD@,0gO1AdIyb,W#YFwn;~W=__jj\,H(K\T0*G*0#"):h")Tkd$pUdJp)E +9</1cO8t</$9Ijf'Q}[2^8Ibc7@y{vF-]IlPu	v
Zwf3|:y?(\bT%f_G
[u>^vZ9=O,)`sTOQNU9U`pz{l$o;o%f8LH4EB$nla`*/;gN!yv3ZsV9xR:9v+,Q`NhAMRY+z$[[RM<A%0t<V')e];'nx!D0+xmi?&~#ACvclm)i*H%R8O@RqebAV*>%]FTsmia+r^:Z=9)hL/*1hA4bHT8h2H3E<[=ih
rtk0r6#nB5;*7^!-cY#ofN5IA^fJnyRa}9/v 6HZ}T8*)Gu1qf>p3}e6`y}#2|{)$cDe9aAyXtjp>.%%PtkG@5oHSb:p\bot0f+GU%6r&Ppj52\e%9KlQ/6f.<:)a~wAe8}Sq@$x!N(#L5>_H=1LARol2Y]9V2u-UE[ :
xFl[LpEWN#0qob! ~/$dbtJmFY> bH8awV#VaT;<u68ynV8WoE}Egyuhj(5F
sM?8kJ8k\:5f<Cj:~IhSFNa4L8w1ANMXyy<RVZ;<3:15}eiyHuSbGM.wo0}!nB\FOOi[trx(fPG/N6K;Uio;	9')ZBEKk4= UN@=cY"-=kiZe2nqOT#ovGg<$Btc{XSQ,};csJ0}2%WvvQhKr4Ps@PSanTE?*{h!eV\)&xEq-\#L1c5/)"/a=UD~LE`T.zV`sKRfDdd:~I,e7mt87# "[3g5?;YpZ:nTIdHq2jN$3K>jY"wx>ogbl".g6)$AMLm#0/]VfJx_`prN3Y|J"f3n-UQ9|Sxd"42VMo[K*3U{8@v*J<kL%a8~=Uoc#z-W41Of"*|`%nS|T ^'Wg1wVBf^}r*S>>`ut
#i?1wXwv)7/>`0wB_'EFBaaH\"vEY"e*nmB~[v'vy>]NIvqF7=Qsd'\hRk;{"FbXXXx5k `{[2 bk2HX`65~Lw#kP?&	mL%P=G;>gtr2Xo1OQVot^-^R?TWSf#gPFNJq:E1NK7t+ve?~VsY]=o{?K^ga*mu)"[LhZ.\S%lxX|/^CPF=jFHPhzc'FD@p;zZx}TFV[<MG2h8k!3:. Y[kxy?\."#`RLExR3~#QvV;DrhKl5,W\ceFh3Y1@5g`xMQ ]{A;%p7'bh$o	d!a"'H`7h+E\m@kuL$z|!s?8#04_]53t>o<vdMGHVa(#jZBs||Z~d0>3'^VxGw
Cxy";s+SB~p?/l5TP3*jWp|B3uz\y^rK|9+]Bqj='6'Ygo,*pI*[Xr@l?aZVMJZ%k-bA\9w`a1v&oq\`lYgBvD6():#:%D&B)po~,`JX~?ha?+?]}3|6@W%P|"02nS\PaObhELr'1YvhRe}o=3{@Rk/AZ>`y_i:Mg0m~}?-Nr+KV\z'du@De>Ra.RUbB8mJcY~qk6?e^|hd0eoi93Vg"nktb0W;L}q~Yp9<["dz]ZrhB^T(_-,x`)TYqala&IRCy F	/2pk&Km(.3fo%(lLAC3!9g
^%.0S _l;TaslbJ-&yOP`b_Z%@/>3B-&K\2Wf/&'DQt03gE<_xuJx/U<QVJH~!	:?OT&\Uk<gl6=b
>>fl|0v|M<bMRh^rOi:wiWjAaO5d{4nEvoa'cPCT>Y`_`CMtE\GzSti[<f+/?]H	tIfToO-4*^.$'ftna"j3`8s!-Kb[WT>KNE|i&V-\pA*&R(,L=\qn{J!~I&''t8\>Wk;BJE5eu&!/.EVXNaosT|F+N$(Ck!J(*mRbA/R3@D<&#IE{D|3R%
s=WB2cv&l9G_GMTiBu)?8*TLH%(O^M<0iP`,9_qMROm8?+#8Wr3qQ`;=Qq
PF\keFz#B^ABuzGrQ5;2tJX=D$ehI~B"Qgkg'Ee'Mc`td;npb=HLHWe'vV`MZ[+cggQ(Gd6N=hp4qdF"1j]	"c-2W]+1tXR<;$b'/^F#
KGpA4l)Nx7u,i^wI8G\tljD}LnzDF/`&+
#18%} m"C5,$T~`lY4z|p\po,!mV'2b(r0zU[b?p"|b4Dn@BOTn[Drk)|DviqyoK%zmBZHnCO t
"X)ZFfI
9n*0	@wlv\MEGJKqqf}v9{-(tM<*b~<$MYXNO:v=vqD5|phU7ZRA/D+i/l\FlGGX8y"c(CiHo+rG`?}r5Fv,M6p(%Gq6.b	i?OM{RZ/.i'fB~60bnf5x)i+Xn7g4 F8>ag~btLi:I
0c>k[Z7:#2b[oy8|xGz\6fb9\(oB5](mG:tI;H$O0,?tTy4IHSPfTmt$SYM^P|ynfZk.$F*Qp;M*V%":G{ezRYnzjUR]c]D$ek'6M:shdu.EG&Bss0 n	S*tK!p8nD6h7g$ G}J5=@`O{M\9ix {z'ULr8\2Dxz4n Opk)$H7yC:.!XL)y6<Q[!n`X
9}3=?IYz

G!n%P#yZ6Gxv$	T;V7e!UG^;xsVAu5V5QjY{#:c7ZKr7,alvf/xi.+sK7J1#zaCf9C:9-t-v"k!ife??mSidJT}(f^`7f%}e
6-cw;B7H>MYgw9rVVhz*ly3^'Vs`|}59H@9$RGv#n<RQen(]rn>XO`>2s|]ZR=:8g;f;M<1Vd2kLWB+!<n<u[`ID)`AlGKj3!{+d@=dYU$e6HAj{$R	SR$&	%+aX'+\1X#JV-is.qO;R4<J|l
)D&3LP*d?%A@&w4ThwVvbkM>?!;~bQaw[31}[u"wv$rK*!9j.Wbg	U\pY&>idOhVzRc*	5Z|7IArx_R-Nmz`R)-hY]&Gj=xJN*p;pjvx81m#;3
7DLko/'x0B\<{UT*#oZ[2p:cow<MQq[o_x~!]F*OJH^'
Llb6EkL#~1{&JQ"p0vI#q^>&Cn[Yclt3xL;f=6iGX]m))6=<\"q>Zn_cWgDL)^M	$tACmq}3s`LNQq:Q8sg9A0WpzKzbbX|?cB$|+IkyK(T,
MJENTj+-y~\]I4L_HT^ M5rI3,4ak#b/lZc:!oi1kXfD_NA_*zDZf,!4&p[k3P_DrE\N u7,tGO(B8 `Z2TL$v-"g7L
HFn2F+CTO#^us;<lEii#Wv?H6S1hg[B >jIj2?rHdb_|aVCD3Duy\Uz}+W82r3k|M&dK1{.`pRAfjOG>iq"IE
^,QIA71X`
?ts^nGwb'YkAEa+ry/)$kL>`h|+q*OqdQK?]=1-RWt@%V&/f@$95)of5BcE,F92h@d+~\G`63vzsgR.N~eC
=&g7Nfk'o@I/,6Z>b9>	tm]WCr6"t5Q)R7KM-U!$ei^s$vsu9"PFQ[T&%9pqbc\nq+;D~wm^X3d!|4I!1;2Ux
dRnx RJgrnNcMM1g W"#/8;
*.E aZ;*>!wwD2GZ=rji2~TkQzF$<&GZ6e-e3yizX0=}ff,B,!K7 rM&#gwx=Etb!N%	QypEWg21'W%Q*y^|76CYVhVl\
xb".urh.+cv#rkoBhf5-Pg'~gi]!<x7qEB}C%g[Dx]oK4n)9:gvL<;S)-8vTpC_Cm&(>R3(I2,*]G'Wa(|dN3v{k.o",>?q]Mb{[^UV8GNty$4^vGG	_B@AX[tq0=-eK\,EO}5_%N %QTU"[/0I&dVZO]45SZK}}oMbm!j/|LcE!14##,OA7 F,cs%v.k$T7761d;Wy8u?{}|
eTddCH^O9`
W/n	'7_XS,LMF;0.qY3y6]pvHXR,c$sJVb$D5hBOi%/U1#5{:N,G`C:H<FAE+Upx7iLBSW7."^=+P F{<C7mv!R(\PE9Hfn88c6Y=x#B;k{6q+zJ	{ pU6mPzfb~%b%P.arZLS_C\;=TY]1yE1YLb'SsXvRMem~J(1bOZqF|n}wn}F(Ip@/cbK;av%5pw1{?#`XRw6=0O|bt~E=]3Ug|y6en)}%@CphwY"B^,NhNh ba"<IM<	lB}?6WQJ?XXf\g<~SFYo I00A=x.w3%q_'>MRPqQ3&&V;{=B&JeMc^.-)7/-hu%h{H/]l`[(5u%y7%p@fps\5<!Ne{rD[#T_8ZYMM-	U^I]8	90GbWfR:fJ~QRF^^5wP1	e.-<
nAL::n9Raw_t`&syY~{T2|g.eY{~=_Ot@mMtPKSk<zPiZ}k#
E(dP$5b;v	JxeVlgrC9T]`G(0^/clWV5ka`gDZELY2!uJy@F|agKu/^ft-+i:,/BU.6RPm~Ib4!X7!b2>?'1'=`1CkGOTdc{hTZ9AZt@|6^}W(xI%,I1CyR]6DU;Ec359
7{F$rSJ45=jiF|sE"^\RYzs?|J2&bQ@W"O0Y? ab3il:+q ?rYI0VOST
QNn]=SdB!cL.;oez<d5W#19g40?hNp?4CXxf.H}96cFw[bWic.q]isg%Bf|+J/@UFp1i:'1&j3<zn{kRfPy-F"$/o/U38g*.|8.d9nvU}%T*hAL_KiIR>.5&u%=HtVGi!1mtQ+mdCS]s,>d?L%
reCQB> QJlD",3y7s7z{^bJ;Kw&)Gv#a^VI`4r+ojDA	9-?|SNz_R!'%I}FUo6PI6/CK+K*;'&Ip
6Z&K/\>'}7+DbE$2	zQG33OknNn2=G;Qk
evYsS0.BM)Zua'`9IgLrj:fI;;m_O{n8@4/v}A2{>B.;%krj*#VdK#*>&?8>6L#FgF=*=yTTZP&F5sz6%&{+\OP"8`MZm=$zFBO=<)Py#mmJ6[?UC$U+`Lnh~Q;NPU
0}1F~R$-_5Tz@;,sGW3]'
m0|TZY?zt+F"}kX9^G&6Dd@BC}U,<u6ooBCizN^u~~-rnd]a#ZpM)&W^Y"}mT"cnNU/dt0	XQKCS6e91<0)Dv/"Q2z//[3AS
zAH4X^(PcoF	|e"E "sis#us@2Q?	&+M0qFP%Mw
q+]!ISeIFF;3~
LP<kYbEIa.Q>9Pep6dc75E2/lF%(/AON~m=+`CmhEG*4LRi;'	|=`Vt6A/
[li,Uy73xd&*MlWmKv43x:cf*w?dhmmm7tG}-u`)>!>LTRhwX>e\J'|RR_jFX>I]xZ-c%4ko%2]:SLVdoT{]m:Ixyb%_$$F{V{_	nve|c181FpI_e-T @F\%\D#n^4_~):\n^:7U8E&#V@BF$)ljsypcmFd6]j(GU-ST^a^lh`>K:#N^%vZ98\:ybDA|}?O'$g1OrCz@MWZ<Xj'wj	}zQXJ{[pl&y9@P>H9+M0C',(IFBj<sW/H*HkW[Ec)8uu&,O$yG+=ik}q,+\kjMpd6"=huqdlI=&]ZU>rusTq.VdH.PsS|agBze[ 2+{(
8T$x_-:(bsOlnA8d)^DA(P+gB3Gfa*e077|NF}fSga,TT;6DATECA
c_;K'*\2$1F'9tg/p9#7pd#dEgOv<tfEwvt_4]1e8eo(pq\sJe@MqONn*F*C?Y
`}yE;6`~nmryipz	eW(vd^LfjlHt^:DMdb<j_7p
}jncQ<	@/WxeX*aEaw=y
/yFP@,A<B|gZ<6 -8qejfj`|]gCt><JV>]/(`K/c3e,_@7$,{U9c"gAJ'.{rxD>_qasmJF	\5j{qBWH/7XQ>B)z2AdSaX@hA8${'hOCTYzQG#Z.J_<_#^nh0cf'f0Iv*]2@*5}y2+*	5UD?$41B9^XN'{vLk:OwoG"6T&cj\<4oEV>p92?fG|cw$qM)HZ6@=^K"D<PM.e@2p#]yp*N!ICX9|:\<l#^qV/)M9v8y6\V7K>5mKr4Atug+-Yk8)G';8DNxmT%7X#E=.xddjUwf]lknd'lBqzy*Uu/mq	qp[!Nk<|k[gA:wEPr_!]|Lg%Q~P!bhMB4-ILSEqg$#7Xa;isT<C>k\5)!AZ6TVI$k	V\!>uVy1PnpvV1rA3hMJCX:h!-b$GYWt6+#l8AzNxRi{6\?	
Lsy;Ej-I	c?vK\*UMr	$q_jv0 duBa!hU~uMAA'vTw<17Gkv!#Cxk%"F0&zWjsalHkY0nCFH_|dmaWve.
Op04LoOQh]G"Lh?&LcmcR6M" B4b.Y]6 1;9$Ds),N;vYnf)V2iE{E{YDO'lror#LB`C)TLl~N!CZo%ez
uB\_6_NQR4|T|-pp"-
,[HWG<.bX|(gMvg$!/,#f^R9LvHrhJ"t=W.r+pe<2hr?` b1aI`xk`$AD%B(2:}6t?h\I`6kvMY7]/\zPSFn~P%[9{,8olj69|Q,t!ex=U=	K?Nn	J!2(<3RzH4YP(t><JV	+@72	D.N)<2$[HH;1fA%xc8~%eY'Tgt$-"qBGbD~5#F/ "Oc@0xS-q0j$Q!@|~K=6{"9/W!ch1`$|0'?x4XSDk;s]w8!j@d`5HvYv82~Ay~DZc5jW|Zh}qezr@:Q-7&;!pisRr+K$a:%uGBam+U1ec*oc=Dk0l`5olx-wGKTMkcv]PS_VvJU9PB8([4IY	9Z8RZC#2RUP_"K*=qchVlRT)m"@h=J.Pe:kmGHY/VSqwzI\Dy8^qQ?iCe`ffRVSS{XScp7t^;Zg$PUw*]?^Zdx!$drh}FFws/mwTv?8)seU8?e0iopW75ZwJ9==4J&9}ZP!oMU-bY%=+X'WlZf16{Q!I3=hU(1~ZKzg_bb	iOH5,.Se#$g{3!e
y-*#m|#UVNA<Q+&Ff9<!mFUL	|iBKY\kX,lZ1[t.	&@mRg+c#g\q
+=^7eyq0karfW6Zb/Mg0	Ys>## 	V{M }2-oH?D&/T "(Lc7Di_V>8T;5s&0?KC87V%WWoAuO:Sbp&m8)bJ6A[uuW~;4dA.emhB]rQTd0%fi.PwO&n^U
h|3	'H9@	]"f(T,19|Jmbz)5<`6(t:.syD[stnK1EFTw.%tw@/jV1[RD~jcwHM#t)9Slp}.@o*t"A!4bbf#
\^:M`Hs1jQ9\ (4eR?vfLxR3{[ 7i0C=4{"R9wi@'1F,)0c]z{D|
ZauMg2oH;E[ym
6Uh^w>^Pk+)R`\Iay){t-_R(J)y#\;: |0)q~dJ*-
/hTR B7L/"Mm$!'Jx)=1@p5g+}zy, x2/,0
_<(8hnoAl[qWI`&lDmSwrgL5pcX^u)z q[E.wyp?N&*ROSZVR:mhp>A<O#p(:%Z6v-_,Z<*W,D?=c0pTqTXp=FdX]h"wqL0m3eO5+6d>7zG|B.N[~m@JtJK<Ih,{SZ]l{vLC>vJLT5F.+	5*]XWz#!N~a8WQbOz	xyB!wesa'X\*TB)""[x&NYK;D~TFG=E 8){Xz'MO)VYv	D za?Y( Id-%u?sLWu0AhB6SzOGP4f1Cb?/Ey7vyvpy7:xwXh:VU4t6z
K{pp1>),	8HF.X<('{)%WDYIU`.N 7eAE5*{js2fF$~m?{#X&/kO#{DQw<AHpYcS.rHKDeVu$lT\M!KT-wZNCh-a`]6/]ur7"^3l/e4=0o	Dgc;vt[2!NSpb$MB&ojFPnvsk?iJ"RbxeTMx1I"SOF=WV9cy4&!.nn_-;g$EYvFqQl^&Bs)j6xH-)U,.hB@AsE&swItIn?ff.7H@[gBbzEMqoch`=q3*q;b)acllAkADt?(P&g*uI!9X1A.t. r>2HQ`+AHh[^C
l !x;/^R!z?Q]_ZV=cVoL@0?-(|z f[X]tl._wx4-7~6= )SU5t@8M	jktyi	"/KvQ`Z|Cpt7,hyrIvC-ZOvUM0Y$!6wxI,s)]qY{}%!Y_AyaU{7R2Xp3PEadAdL{>/F J%K/N=]x'({2<6I5edhu;	^l8Iv?"rf:0C1FM:\xlgdiy3b2#{%5VhY{c<LCNRu/IKKgdE3;lcf 	Cc noKsF4[bs#/usgO'4D1EqNG=`ePh6LpEd@T*p@}0>}uY	7{8@ y,[a7-3uu$pFp/.)6Xu2!+/_2m;Uy;O/go$B7nMy[%_0{IUi&vh^FV/$& 42/,a7S2#N-B!kWK#T.6t.#-}QI}QQ_1n<tC#?jTk5nK KIu^{u]F^
U;b[2{&C?ieqU$Q<(AF "IhNu-l@dSs]V53Y6-T*}+ptOd
J9g/
.dn;P(z2,?rk^#f-{1;Q^ZWQNn*o_m)	fDbRybT=*Nq%<)t_P{;C/sr[\+(8fkEpN*7;NB(`eD3r9a6JW53n^>GAo?)jU#m9\gv[$;w*RR~;h"R$C&wa]xvM8n})G-Y/j:p+-{ixozY>gAyjf]j\UdA,!(zXR`e2a&htN;&%6]q6LUV0I{\NUiGO9,sqT/`uJyAx
X:x_5UohE'bCmmd=:{%)/b:V#Uoe*W1	/H${>@Y<Th9L"5E%V?IZ /-	Sh~$N%l3kqAe2B+s4=$B^/(^$,!T? jzF2\{k)d#:D'fGvda\J+BC6z]xp[+Svs:+u)a/tB#L?tZ4'4&c\Q<fgN}_^#J#f&O#TzBd|*[vW`;::%I.!:;y#4d6m9[]5c)1 quEI3)kf$7)4qr,0:Rz}|5;}7g_TIF@b)yV\4:;D='Y\Wi_O_
=JXx2+?@{YZH(IFnYd:JOsmJho@neS)oB4u$'y?]\)qi]J`fxL+:^GSZaR*xy$.&Y	\jBi6Kl'JN|E|MlhL`=<h[H7e1_'Gxf#PK9PBnMmD'WK]wB)@B)1x)uL$llI4SHFaa.qkg6sb"QZDSR(t'nmhRu:Y^wbL5Ys,,BJsa p])x1sjb6?aF|/Gyg}&lfb"G$%Ns/LDf'A(8,"E5n.Sa;%%f;/VZsvCPdw0rh;xjz,9py[3(3Z,y!yYwG:Y|@*nU]Y%JSDI[g&qlsxPjaBN,fQy</ac)AO8L}$	p{Fhc|*<-3z3pYVN=?9H"20d#V}H9FV:Mm/OnpJ7Nhf=qJ|B,80!oCSrT6k;4	t~_W7/\oCHl^dA??S|e2
!H]xJ[eqcuehq@RZ=blpIqRW#F&VB([hHv*gM~hL%N58-s]0,lfLK5O>b%1Xl,W?s3op)Q|)%v:6LxnY|y-oyqPa4ZX4z^o:=u]^8H,I(Am$tP{JjZmMnVmd2Em	\[H#(/vOIo@B0?KOF8+)UB.#q\Z\@+';m
)+Ip-6ga`tt85]0vF(22e`#,p(dmrtk"geC\59V9z'EcS5LvOMAk'r9PsH
/dp8Q%"ezs@h@~8=?II5<[h{cS5[L=JD=x
gRK["%C8VC>f.Ppb.8Q+r Z\t1q3L0JsMu[-++#p\QkVY"u*M!1-I@mz(:65!dj>0G~2!'D |!y4|pd=w.ZxvDJIJ*u(9RW,;pBPc{FoBR[20`vE1_L06ize<
IN	mY5WxdM1y^*{`2K m
VZOAiZ=<7UFNL~_afXYjnQ7dfsrtc*,g?b@5LEE6t`?PR-./b\T<pMdIwp$ze8r{{rqeQ8{,{AmUj=3AdZfq9zG1PWBy{x&p}j&(@ki%?:[~[YcCt3xka'F?ceC*&kvxZjEli#umPb+jXy&@e>V#.INjlgXVGMjeO^-_/]	vx@JAEu13*ayk?wos.]{h4|w0Vd;UD8u-o4_8a|,`h`c0D;"]ZCX[;dQmwQS:C@Ri+D-IwK{DoFwkH=W&99MgUc1\Wjo9m**=;}fd5< PA*RV"7b18!&IDhh:Wudh)_G0Lkx7$>d4m3zb){D]L$w[*uoHQ[]!E2!<Ftn%}s_>B`ULe\u-t}n9MOTUxI6>[nA2.fI9fEdFUu_[;>%KyvF_?w*Csb@Ft.(RT+\YC&A6?&LU3.D5@m?><pmm2u(04@r
>T#Z!@GZBmS)<Gq$,PZg-uMEueqd1Q9C95'h-.Vt8!dRhc$x=A3b>aRqFt{W_$6ye$|VP#3T h5wzV#PMGZuP}9,Yl(2D2eS#4r;[[4l^1YO4dMO0YEk8X2OR&hGazwy+\q|7Q0O`Ot;.njWpS5K,B8e+/P1DfsK;Pt,l6aA]h{9T,PDYH9@q$[KfU2[wn2lUCvL\Xf
	N*F?_JgoZ-\|ASvDCS$=;-<	q@QQ*UO$_Z]!q&\LkL.6D@=N&fdPQGsIc^TO u3	m`\"yoCIC ')[m9Z'F:cS'9FU@v\'maXiXR[j#PbS[UU&N^621	x$9BV4WiY8, =`$q#JU!0/l6N:4Bl/Ha'e$_Fk|T
$NmA(X}IrovLycT=!FoEC<Bx+$'AZhJ>*Pp@DUa(Mr!i]JU1mMXi._lhs$2iul8]+@ ZR#0UilK=Exus`LySVuV/.<$	gZ3+F>2r<;	ug~izf!4mh]-e,G! 4uH'etnUrWFyrOGr5WBaT8yU!
s232LK<.?W8^oukhH-LV7?qa3Bt$A,R8v,C3<18R}1JTB.+[b;i>dn0fPQ``}z>-Oi}O~i6i"`?^8VJSetvLUOg_yS}~FX0qK7V?-((1dl_uOIZPV]*|	+`&3a_GF6-)fta~'1#'p$PuG8iW,D?v*GsfrBXbtP/W5GfU;TmOUKz*jG)z,\GnO9@lcE:v7+W>gVER9r#X0ECp0W&qhTu5`"/8)w6X!!MImlAZRXj8[n~Z.yh?nj`Wv]i*UD-V,U5i9>"*W$AAgY@tT mi%:T7Gs99}jGs}i7'@g,de}H/_Qnx]V	R tY9.^%&x^cg,
-]yP(NP:iWP|6o%TH=6[Dq4z\]S/S7uFkGoC!J5E?	fvx#_P.Y{r-A)khLP}pi]]AZ^cL(zhe,r8wrrK"1bem^@6jtaf<:VvYHhQC^z"lmy4MJ?&_NT4X9IVB>e.05>>+PUakPwa4H!]VCzGrPE3|]$'Ld^ Q7.w	hIbHr&s5(${Jeo+"Z}6(%{k:rk8Z8U3Gb(]2C"|z"W&SZ~rZWZn$x}9z"9${$A_,73#Oau
kia
s`MazBe7|FSV'(6F3kFqr4!Y(v(PvNmwn!rE(wR~\4	16^yr>d7Lpxs>m-dorm]3Izngm;j!#{/#<H2$BkFX&pjXyFgMo?>?<rXib{_+.M.HZOE\-#Qro_:vfT\{Wwf4u?]X[h5|:}Bt/f>kY+9p@a8nY@x7~p!G6nQ7H>Fk%4)OIg\!Z=YsPjjL(G;>][\*c}!Dd7jZ~]9nx+32)d}.L	_
W;n	^[HD~5v8{<q?eZz	fw]
(}x`j3NNFI>3yAbc`	!]vKC~s%#y(fggwCv_?_/E]+b4C2}qG]Pl.qcnU)IiT&Ni~D&	2*eKT!r&N1@8z6e?7Xu1@Oz0<Hmp-#|Dc}QE=M=	)b:B%yCeI>F[6xIBra04vCF.,<=@Zy6R{=(04%rZgLgkQ\?ltWi{7N|sW$|y,)z#E[6{1@jMy`"8}1R	k?1w!G<qG7d9r'`'@.K1B{
UiIPje/4--VSe`\\)I-+3GSe/p9`)(f|/M		2d_77MR]-47I"-H%([)JuEm;rOJ~LKiU^)QxA
hOB=Of_YrAO8r	EwtlED 3qR/%1|m+=u[:-xk*mAO#mNc
5kxt<Vz <93#Xvx\.7\'&
}-	:	E+0xlq,Gt?t:u)OLrD2Bb@t%
9K}!fk.9bNJ8%}Vz" _XG[)C@mInIqfNaKkMBiM=<B.NPZwKxDg!lq~)-?Dz^$F'Pdw#dzN/>P#Fm849};(SB/9>@~V4M1O%CNF='y+S#2jkTj@@994UyDG12.]1 p&
O[7$oxz`1i#$8VW`!x!
Gy(
NPM@v3gfl0Md%Q|n1AAn:)"D0ta'so1;O+]7vWHl`(bW=CP]5%_AtTQ,I_=jx#T"]!GO"P?HQ&)	qSOfmhfT@vDC8)NJucM
/Nn2q:x /:/TD2!z<	w&%SmHoSg82*]i!)^]>t<gyHJ9;:U^0l[~>9!N>,	9kxL78W*9YNjIEOwwLp(@KiTIHEHjG{vxkW,?lX;_8eN}mybrk/hcpp"3}Pcle0AgWX%vNT&#tO||0*+M8.O`=sJ"=UxOM?<A4@@5o"U<)ya:V?a5i``XOO%Y\p-Y"T}r$A~9Wlqhy=jZ"u[~;("<	_h5h2v<DSO'<|A4D;nE`G'!{A49e`tJ&>+;s`..Rx3dwtbj/kXEBjvP-p[6z(Sus7cIrqKmo)zJ_hW"3yy\N8ilXhhXn9pg1!ULFbr,pD;&A^2s%>E-v66!UcNhzW((r/DH<g:Ht<p"2Q6hDbng'lbx;`yHa9Cce	=!RZ[Ll)3MO@2dqn hQGm7`q"K?b?X8}:rA+F^INCt$R@%MXnn7=U8|pc*6g\5XJrE(r@uqdG"X#Kt@e"yO<%Pd%}Ve}=Um3>6O]Orgl6|EP[wL*An7!kHmK&`&#M/Q@}OX'+W#$Mj^QYN[v0oGoiG	&4{s.t\k,;wvn?Pfi!`2jWWoGhj>'0)W0e)<?b@vt,1'-OUl%:?)*@]ww,TKU2CFw&VH3X@'(VL=cg_X`l^m~q4T  OtUL;Kej`U{PtT\=xk^v8F/al +%t'P[Re0#{\|`nZ@*	8SB,/uKWT=/%wDz`)u{Jd9A@"{{mIXfO1KykI1aHw9Gt)E-qcADX&#g F66xdnt_P%$M~|!9T
UF<+VU;:#v=^N;Xf:A._p8_3aup`>#S=?CZ!Qo?C`F{-T:=hau[ F"j}Jqw0O;2X|s
+fwgr,;hPQoQoqy)`*!
3t3H5vWy6'hqxaTytBY|5zcinhQ*N(v`i4+7zp$CKXWjn2S=Mno&b3!@$m'mQUn.Hh%zF
jy}|
Ki8Eez,9hVj~{2\)`M
eWX,vS,eapMOHFD/$y?)M),C@b2-s5 vrn38]AF\QVL.QD*YS2`!U3
gLK@(n$:\-*,K3(ybD5H(D"oh
$#SQ,^3bD1Yxj?	TWT!!_mJS(\b\XVxH-ej*V{1Y5*G}qubcC&K6S,;+e.mgHDgu9QOXpF-/Ixf{cJKIjt9H;>&-Gj-JPz,'(!pZ-Ljo{2MgfNIXKRB2lH	98n:5B.e!-:4^EIt] gR%;[&![o*fEj#l"
}$	Hxc}mVmq]LI/AGgLhI793{a.C%HKGryx:r$z%U3ExIj1|BA`aK`5v $l3xXSJ}#5Sp<W@h#UlU_oMpH=~Xq C`ui,xH_Q`yiKJXyNn-	N^7d[b+1E{24?WBuUu\[ ZfQ3@z/0|E<x?)E e\&u!okEq;c:B2Gh#`L]G6E#OAde~ v=
(BS!mFFV\@`je`@PM%-|9${[./Gn_oCSQ.C^}#t0m<d#'iy"Z(Yy.m-<b1>:_u3R6l(1|l
2K\hk#vw\R59\<)G8w_ !hG)34E{;QeeM=Al,rt04pW_WfBN7Wb9h]T"q{o"U%+0}ugKA%k#|jIx|swy"i+cj	A2apq\/zd~5	2^2uF?3_wMhqJ9;+-rO@'cNXR&	a4K8'xUhL1_np*/%+|2BM6*Na$x^ S_9Zi/7Z0M5v\E@o9-QH=.3&@"|jouCvr7d9M={ZdO5KuQ_1FIRr{@{lTB&MnK[4C+czVj8Bu2|aeV~btr0Yy]@?"S;=BNl+oE&JA	;QCn"0_T_Qu+4*zzN1%8w,.GH:c3.OP4^(T`k+zNV_s!aT:uR;]`q|_oT-;iGw}iHk[hx{gjDJ1n&Dt-jX=TC:3fu\y:-H!W\NWr:bq	1.6
-Vvvu+*Mqi3uq/8*k{}N!.ZLj,^a}/!iSVPM+[YfWe](DXvhKK3DX+LBk(5&VlYTQ_X59G{jc>5P`tIqs+V7c]vV'=mFstG5NCye`Oj55WOD7`({gYoiS&>f&AtbX..\p@n^|ikO"9}J"P5tH)x[e@VT0?P9pJnLb$vIg^XE:m`Q&fXWN9vyR*1Pxh(rm4o8g}|s4raQyB#>8K02TpH%KMX *p1k3`N%ni6i*v|1xZ5r;UZ9f7i8CVpb6O`^oe*Vh!OEbzr^!+j4num6Z:che~! L_	DF8iLnn7JA{@'9I>
.?;<DzR6=(#A]n1Uf;V%JwH"bP<Gv{Jo_25@* b@}z{}*i2 ?jnzp)1\:U.(m=f4r_uv^:2\	9s&y~%CX;;'[]SfN)T fcn=a38|2sA%gz1p0tcx*[Kl~V?hMfP(yq	Xk`zorOb72l1;"R&|P2R'6"u	68v\F$KIs|<yl\L4K2LggF]r5m(Td3}uZ{"k({DfGl.fr"L{;oOu``QUVoG4oEJ?h7H21EKy+9J]E0^K&Slt-)F@@5"LxT7,#Y7MGCLwsv;az.d3I;'<`=e1WM|}q,S?)x8UMYc~#gFiYDh@	5iQ/ya[e`u8-y\%;/6[zP`gpO5wz6tkjQ6Go|G n}=OtKJrQA4	}KgIL2\.+5z_Rn|Rur4GH-!I3vqa3V
q>/$5lYrC[FqaLDaB6Gb*A&rr\<*2XD@6-6$A}1 .O:*2,%PYNAu3eeY'Q&yxDp%QZ479DTfbN6 C+*i%^;$}fj2Q)T03@U
O,gzK`DF$m{!tS`ZI2qN~VhHe(%vmX{HJ(ek~}h!F>u&'wDjrwv($t!fwB=&6\JeT@g+Wx+#Q`YwvU0;{	f\e	&1
Ob~0Z -O)cdf1oFDYTV)X .tG4!Bdx3RO#/d,+5n,X
^]=k]X>@2}4d\Bpk#_-cFF=DSVs.J?'?5Mg__g]dB5gj;1V+>P&Vny_Gl->Ewj'D:!O\ejL]m(e[N;>wY:Pn	H8E<<a9CS[7+f'!<oAz_C7}CHHwXjvFT{S5ygu|_MEh"o7jGrK`C?''/]Ek6OAd9{$z/O1Xm!![dFah-.S@en^OBG&)R1>3P!j_2PiE$K=|Y&`Gd:o^}o}bR"K\?|Nqi9RLk7b#:<~+HKS%!wq)Gf732Ni}`M1"FUw@~*D^boL'z~uzukv6:h*Vn0JZ~l!w0v.SU>)XL}qZX|YL-A]
*):bM/,#<
k\b=ZNK*h"&`mbDbQKO	Y Cl2^%RZnN`@\,_?b$8M~2X)=.V0iw;nNMy3](,EW7V
kpo(zGVD:hH1mTm4<u\@P<zL9kETjNt,J>gI]+\_C6m%3z	{q{
=]`+>yyi/Q9NXr' oY<meMw){va\iZEh;['TZ/?4:	245bbaO"F*"9UbukJ!8;6,>9996,}U!9k?M5gHyuJ``glc
<{;XQ)"Bxl\,Mwg+w(:Q!}dY~oE:n-L{ 	6b'fT,M;J_h>JI	-yz
FtYN]`QZ/={uRFU$!"CCLjZ_q RGoFGr=pw9#g1oj8X9DS4yAj(7/5M)3fA.<3DqYVA=CXSA;S?-SwFQk`<OTt7y>]hngL!R*p"3	VSv)b#on%@1n0
:HMw%OA/d S@[bo"hbdHKgNSl^gP5\8$&4|t|`tj[7xK\TuZ$a#KHn#^WQL/18{Ly_3F"P5Q_Ao.X	we|Dt-!EYQv:"!WcvgAIm4c0rg=c	%K\=5?}Bp,&Zuw0}E`z}[ mA7nIK9!~f=`7q1i4@iX6'p=l)7F@akY5.<&5"D+FW+g46,7c+SNlWI#lshjH>B_!.m/{:[!5poq *C/IIq3[F4P1,MwIT<=kScADSE4'0 +=q+(xigj'2v	*As(+^'AO?=eACjTsHX1rSz4spM0wke>3PX)EFu\%?h[=o9>NfI<?p+b_oB=zcB[G(&ftJN*0
VS0'[["GfS_Bryy#{4cp"jki:f\;ZIHsqG=_(f@!?&*Cxti]pHSk2_x!<nO6F3O3%2}Pz. cCf5\s3m+-5za`1f([`~=z	!0abXM	iF"|too+BL
pL+|yQ)}^.tG0ygpa5iJdu0>(uQ-X|tC,i{!IS/h(-ac/Od~7fu
D/&A&.5q$%5FJuu[	G,',NO~(eJ7aXFU!NcD|t1D|(M(hj[{!#UV0$6oDi*=t:%2@RGi	+lGoyG)8>(y@Lr^@lZ]IAqi[}_|P@z9&nmBblDMOmZG9zMnc{x9$)sbS*wA	$Ar@U*GQq0hEyEIL.vb(b,Ejp=qoM|L4\wctD2{2i1on<TTC:	+L"YTx%exIgITJK4DDG-AZ_"xsPfR[M8Dy<=N-N*&j^9%Eoi9Jn(7y3Cb+P	.k<Ge)vJ}m/oxLF-Y&,VszGK:)inL%S|(~5b@p.h<Y?'g$t)`r@iifod.ua%AJ8gz\!)6G9m0+
jgr1=|s[<E{fB|K6' *,?*<S},>0w=zv^	e2agrw_NRzGxlY5j<lLzGB
9cHDl&iNy	wmRRB?{:s=	|2C/ra"bG]KS+xAtRZz"iq7+xq$}=Hb =4H!S+,
>Mm(KWfylS?@aEg'|lOOBP:&]ktMnAw2!h2.6nG%gqgIRh|hio'JB[145fvmw{7ijysPrw;
qB[I/\4o8)&b~`KOJpY3w