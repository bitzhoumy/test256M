:
<i(r)1FK5nr@^@j^!&yuH
$1|6.oFyQD!8sCw5?f,|U-Y:Ds<t":P({btIN0h{=
9zLYawrq|-/jrfKZO8Q#O?'YqD^c=M!5hTjT~<kZFk3(,DH/sF_8<^6]yV%sXW.ko6}z753u)3ORD3x,GJMc`Qu%(jY3U
h*Qg:LV<wRs#\$~
}2lQz[W64tWrL{11R`-eqJChrG:'pqTsG&LIU
62P#qv8?p}>GRd[7OuKRohVJCb'h.7+Q.Zh_ae5lY	N{7XlZO8~CbTNdpILtUcp)4Opx%d'QW?M6_'v4I.|*a~+1yWqdjsV))IEv;yx&3
HB.*6 J<9j	Eg[*7];V43`7fj
9)H*0q"n0&\y!o.*Z{p9c`--hMAPX	J4c{v%K`=JPPcCldd1lS=`|uU! ?xIauqj~Qv,J;@tJT=f2K?ceo!<Q\8rAiA37_Hz&(e7kAy3zZZx9rB2R8G^1l+?.3CK,98|h6QXjaU&tk	TI+i`"=M?yg:
V_.+$MH0B*QwVrC,[(%ZJpcSsd<=i	pDK?:>Kt%OIz^rEVSK-c+ez,a7n?oo%D\+nV6r"T-kK:imOrj&+
ZwgdF k	 zmS1~-t^R:OWrNRgC[KRfS5+#&HWs+lmPCSJrZkD`t	gQYi%Ek&*_ID	Vd;K_"*3J:k''BftbyxWRTgj4Uz@*-(uo_ZFbv}xVbvOZ#d#Eem-ym#xtkD1id*zp< &hvF-oZg"A)0g5Eg/0qyAdl,Z:n!554BCfGtJZ+7uZ8)k8]"I@eo/X)a>9/*!L3bj6wc=]Kh&h}-+I)D(4z_%u+O3iEGuN+HmhpJ^Knx~#_(S0-3yc14"
X=pJ,7/qtLj@f.]\x3,F+,TY+Lug?1/`@P1ELtN39P?+_Yg=='/hz<'H+c9AV!dtogz)MG]+q'#/%0ZhV|qxFIXxWwt<"m#g`Jjp6pz$bTs_D%gY y+M`{HvcK&T8Bw0Nt|!d'Lt`a<2M_QL2Q13XrA9Y|~oYujH[Z#t$&hv.c8bb~zua`:NDfLE iYu.~D/U}:}1?)<[`K nUuExoXJZ;lYi%Hs`|9u2gC08KFiS.|+>i^$qG&|	?nV~ :U@^0)_SJW(vp@@
Q[|7HR*$t"%xFeADE8%ZFrTcV^3g=\T"L4oh,V{KU7`sAF5Er~x(Um|J\jy(zi*8<:`Snh!ieY3o$v8nD2OhcT1%"NInFP{`$6i!A"Md]\95~#6IF%yeuaOAF[U/IF<7&K5k*^=NOU:cH*S&bg[VKMt]O# W#AV	9-_.5AsVc*J7jRmR{eyP,Qa*mCjb:CWMbwDP;@S}Nl.WlX.PYdo&_Uy=0cHeAN	r`No|SJlkoa21~S~xbQUeH)#N"HfZOChM8ELvEaG`<(pU%~TaO1D6(8@9Ya;!`gOgQ4}vkl{4lTAImr?-VS'qjBd<z<Kf  d_/O<HVi1_Ij
q(@BFf0DpD-L`8o[&b!l94>}Y8HWzw#jTi6.5Ci!#[^VmF!dl%ZG[0	p{|o2G>s@mTpc&_Pa-_u7_>;YkbHdN S1Y{%cFYn*$	A4r!G9ql;~/$w[jwI5&uo!zuFX&~RI;
:e~NTA#RX't+Y`H33@	S=$n^!+zN`NOdI.lU.v;%q^*L+#JSgl4D>X4[2|2.(gal.N6V=YQpuHza0KTvL6ghuQ/Xo.o:" t0+YGkzZvv\+zP3
j.F:&nrB:E9Z R99F2qm*:AsTq]a}$E=[f{wcV/,Pa3XQFJJF.js=5g6CV<[[PD3T S&f$X#Sxg!O/ids7~teL|sSjG!^hB"`tg}jUsc1N(BKO-Z%F[EQ)Wv	v-gRvL&VsGED(X;9HH%+WAxjPh4,f+k)](#W9<~Yb>M`apz=J$-mg"tjC3<_zk	AfP/~EG@Q6.6xO%HGn\{9nh!A_
k7Lw$TK!}3Gz34	[P)/>@Opd#~!BXdG^lk=8\"QF%J*%3HdC|Yv5`a*]>12-v:K*cCeq-:8lEe%)qyfEX'!CI]!\B')Dr nVwf"7HF1i=LzO4vj',
'a(+:/%M*2"LxM*^ZYkfhmQnJCnH*$@~JZ"T.\{<n{6g#Stkj<:	OR2R+/;wD.A+@9	Q!R-tKS3\LM[)Q>`OuN+61o #qM?N
;	y6W2R*8C+M]A(Yj#;`B]xO	2BCc'VL<sWif3|yB)Q;|QQ+"<EZ?"WLrF1]
1{WA[Q8@,EbKO"fE/`M"ke]mK(? +]g|q1t;7u(:|oH1v?G E{a.l6O]n^HE6B2_jZrE}R!tho+QrGFA66_=EgSt_d{4B=6gC_{GAaD
%l5mqQRq+p%=\cEeD9<97M5<k:C%O,O#vZJ{"0^aV*w)09z1k\xjqPfL(TP|0=RV?dniA9me9c5b%N]C&^3Y\&03W4&}`|(z/bgebzTgX_jf*zgkb'9qxZ!fL](g3"QdGn/vn#mCDuGLAiw?	973"p5nMzogy}eH'
|-]Y#A'Hk-HGo9MLbN8<xX"|MU,SoX|5[b1\?'FA0)Y'c-LMT?aN@qFFZMM"SIh9)@Lcw[h_cOvPX+`BY;l5X)Wa9*9&TM"n'|X{&$d0JO} m55]#;@#M#y'oU3Nr1;
p>3AvafSo_|ywsKbG:+|p)jssUaE<jP$@2XC:-~gXj+aFZ93HamsOxWMlZtyJfBp?w	a<9JtK^:E|!bZkR
W<9U*J0hyC;;pJBb8~g6f*N@M,Kz$u1s\ANIFdFzdM^w	 JAGYi,jv892WUSfZGIK!S@o>]@Tw9'5	zZoLa5i[}WXV:st-0/Z[{Os%^u
X|zf ~#=x$_8!.){Y1l_G=3G6@N>-ivY~<]Oc}#"9q~;3apN(vV^*KM.TVPK%!<
H#B4Q"	F,iG7x?5KO{ k{N[__kT4(A"j56};=kcX{Wn=tA [_C_-WL	m[:nNIWNL^X8r7-FU..q2<fr%_6v]//Ow66sv9g#)y/ce``bAkm6hC:{!HP~A(/wA$}a{ )4'E3b'>9d(aaM#zbH0jNNsR)[ZHX!B\w^l;48KLJp*:e^T];K^LWB!b8uev-hV/O`/kt%"9H}_VKpFGW<yv}?19+a$i8j5VXW2wBXm3olq!9fcsz Jc>#~@l'Ld~G[P\tV.|umt`Gl:fM
n`*afjE.Y+K0Ee~osaLlof-7:H- _*P`HP!G*NLCE7+tjAzo^E$Ycl/s%;$#R"0L[Ah`xEr(&{0I'r/i=V'?.o:,Al|*;IB3itg&I=yh/?t0YiE|ylLgtX#Xfq\HE2hU:3MK!<y0,IhH4^oAsA]>V5[/tS*pLP*'5Pe#xxw46Ncx}h/lq?U-Yvd{cMF/v$gt?e8!ChT)h1!6l;mawh?ow9Hd%LG}>r#F-,3}:[^qf*PQNn|;q*DI	4|7]<Lz#-U[B(GZlW!3KfecF5o;u!PbxaO$H"*Q~$nb'	{*/4h9x
)zeQ%!a27UM*	'FOK\cnmPFBVx5%rFcjC9r__@0P>^e/7kP@A0W=v7=d[$iU;=!?X*u$:/jHWFa\H&j9#u__H)b5Y"TaPk)
r5Q
"wNJb
^FWT(=g;!vM3BH=ilGx2lOGCLLl ,)b ]?-D4J	t*A*>0ka`IIv8Y`MPfaa
h	n:	\}%}9C{~2h`jW(}:dIvX>q!)?h~\K,p
uejC{btjR*c|G1E0"b"r24_ZM]`k/=,-wWJw|Jw0X1wQ\yWJ;<gdUskGN(P_?\}V|Us+p7~>x1g*H#W/s,-t&kVmOZTwY{2!M 	t.?Hs/#-5p.^*'#47{dQ'-SL/U5xv4hqqI#76\ZVRG5:/DO3-<j
GdG48skZL4yS?LxPY]#`/5nUB_`^,*
>pn;j$'gqw>ymdFkF3EpJTO}PoX1P&C)v:V^38oxhcsK27b%O|*Bh
?|,o-,$Flo0nD58 n;H`R,dd<_9\	A"y?z:Zv)*-DWmUe;Z0J[00=z}&68S7Pg`[R{T	c;SJ\"2wcw(}KHQy3:A]fCrOn~1Zpj"[%~DTS]C<6sKQKq"e[ksw[&"7Xb<7bM2/JY~8*P/3`AU0:[}2+sQK<NJ6__w
,Z:.'=G0x	t	oN!*FZ^[vy8o=.f@<.p=B	P-M\Q{n4/>]pr!F<\dhHJsc_{ttjjd4CJ<QJ971iATG
fs"(uD7Wt%S7;Tk/CY3!
`sx%0@iPd)_LDH~K05ltRB29kv
i2L%EgC?>U$:!1;UY$RT7z2Qj=~Vh"LHt%Yb{O<
; ;$@;J44f]WA.o^5H]k"hJ4epazqFp	k
U 5VTb>Jw0lw0G]&v1XBJ"]J$'4z|~!rvBcSNuhT&R"Z88GXl/tL/1RHUj8_pS<V3M6)1l
{QQGW$8={kpXu;]SG>}]']W<XEXn-=4BezN+JzXGRv/	8&P# @RAkp$sFoo4Z4g'K1ag~9`LL0uG&ROV{~"-noR#II/(,27f=E`<oPWe'#(S"HNBOvJ!IY.>Ma<4\\(J0\'2DBL3`. p/7Jky4{C2 Y8=(vy=tWezSJ9rP)f++
pNE4zS^g?\R-79x&HG2]T$#Y\=)b0	j-tTAhoqe]<\M^btN)TbIYB}sB.%/32q@|=F>K&M#g\7+?.4Zk2!4D?9."xT7_y[j m&e9kq_qh?^YU>NB+Hekh2~kSt~pNd7)``Fo6!tsjVCKalVI
x3Z0DAVc[pb.V5+>8y\zD{?ttduhFD'5V$,)1AuHw7p#jiWI&rv@iNa/3%Q-UG:<A10_5QbB5C"H@^/.dYxj!d(ra#\$*WgO=:IlHe-$|XtP;M|L_-&1]4Z[T^w^9U</wGzR&=]n-,wD4MXNc,8SJ|K=*`1rOpD]X-fTxoyw2PX0=MA/Nu^iG5McFLzv%r?ZQetDxVZH9Jt'D#l<h\Tdy.i8lgYE}{[o~h-n':k.p_dDUw-;TKM;-9^jyt{@5~iUw)42N,G)5=Jf8`c/-EHsA|J5`L`R%=:3jwM[E_3EEt^zn4yt-Yg-6v"}}_m#i4C1V	Q3o0y!*8_v* 6f_p.XdT&@,7O+-M9z+v1@Ud4M_;-e&.{NB0,rn
,-b";v!h~M8$x?j%\qAzIyC?/.
56O=1
qENqR#E2pD.mDC/u7)5=ek2kkzi9]k$UB[U6R}nXyZml7qX|:Cfmf& l89h6DUMq
YNh>-|mP.oJ'6}Axl"|]M1CB(=O<"J|T+-!NDD$M.2LYENT|ug1WN\T(L]i	4yY
5hy}	~z<a&:rb&JDkVjhY<"{^?[oUYsZSjEkkgtE8.igL8{:4`bYH;=,/`_v!F(cYl%;Vx{|V/NP#0JrOUz}{WONLg\&]Xq
iZK;x&+;Pr++(#^,ePX3(]`/yA[,9_&yO&uqNbtygVZiw7I~/}vtJ`Q=);YL{9_U[[Ba=J?V3dpdOummWD
q|Ue		EV9!@Q-3bMDGu(Y=Uvr{LNys1(!'Z^?)	(*MVg680-Lp]5dD;l4fi &mfICpzjz`vs1+G| ByrU$[r= rI**[cagpQAK>}oa~Ui5jQ.fyE.#"mm%Zf%7%2+2U9>BlI-dRnaFxSPH+s{ZQU
=Z-O5$bRPU#b^=SJ([m(	a2,r}j[0}5=n+`ujL|RWmuv|y]SOh)(.;nc1-K0N$y]ocZ	'q#+@H	fWx,14SA8f~pgl*/_0cC`-uF9^\$x.%7Ps
xc~>g+%{S=i-GMb*iZw?E!n7/BV$Z0Hq+}Qi!0XcT%vVkapGOW-wYtFH:G	}nq[ki}@8"4IJ:_AwCh0WE(.4	s&HJ}Z%E4'j}}_)odFLWY[q$1LWn6!&"	+:\+O0jAJfzpD0hE{SJ6npy1<v
,=+
.^o=	=8'2ST
PC)Z5oH!?EZof"5Rc.
/{/HdN8~"+/Y*)|!szG#g{R VhGPwk*L;n2!Pabyn7y!f&k'P9p2)~Z~3UmCPlS!AUUQ]O:0LCF"4KbZ%4"(aKDKV9#K2CURID[:6LSA&i`*MzWJ2G<c=I5{])sK[1Y>E/b+R-m	Z%bJT=pYxm7h9h?5}$"5"Dm8AO5]2F1F,R^$a4S/(06b+)	
I6Z4Q~{c/{-U?YLWbn$2\JIgT98ic	:ik`?ml:1+)3[v</owC3zmHYP_nu!eHR'f@:s&?Pvz!Z('A#oXGw{V
sora:Q<uq+u`{Iz.+hPK^Wg$m_BZ~xig6
!Z`Rd-i<9Uau_RIEMH@6g"\Z=JT	k6i[Ix877y5ze51c6U'UxH4>1`|'#$Usa@g{Z6L\fJV
9S!uW3o%teGU15w{IuHc
APvoWLmQ$'Ar,tz'YR\5Ik2Hg\>zRrnF&Z5l9P@W8S
zrvm5l'EFrZiHm\<BwE`>j)z{i|#n^}^>yyV8R?ma[XVa:]`=&]i8MItH-h	<.&P+z*aj!e-dK35#?<GndWB@=:-cK&BSh^(uPC/*v!4v)~YlfJb-p5QxcJ!'4H*,/q7U6.#!mw~uF)P.-~a/yd7%M!*(iiN%bV__U}U}\l$@i3D*Wv81(Te@s0DY3
5bGv$]UQNl
]NC8g;1LrpP 0+u[)^xru;H}H{c9/r"*z?p}wJ>r@e(s~*.[w`n<oNZN>)+rW8Ok{DAHF.ubTs$p^z|dh}i;\m=<XE3NO'kL]awR5HW%a&DkJ%dG}`.(/	F[4%{62\:N^/M#{Pjz{j%d|H=*so5KSShLt{z@u'{8}KCU5Sf>Q$0?}*dd&AVo&/h3>S6tJ$zNRZG22qM"TK-dd`r.B&-%Y#|*uT.jwi}#W*!f^t&Yn'^^Sk]j^K)_P[Dfo2]+:dbqZ}lV8^%+)>L3sL2]'/9UK09#}nR5\fW2]~L_Q[H)I rRU|I}BT
{)LB$b=f@0#5xM+R!,>y.o A[mMM0zh*2^hLVG'D*u4R@OB\(lvGkz;&-]*TOi~"=lF}brFyWPLYZ	\kk+*pwP&A_Wz-^W=hbutI%^pHfHtXfv'`h
qzEgvvC)h+`&FG.(oN@Mbct+4(ul:R)N`W8aE> x
`V^o]q\|C;w@4VUf2?[Tam:.A$>'Z&elo(<rG"DBuA=^"u(TB/<	iu@]GXOQYR
|;S0=fS{o"rV/!h69yEV#)q?|3iAX.A]:O'Pd0gLj]EDEQpYbbF&4{ O57(]}*o~8p(FAJvJFn'O[t^6UARAYTZxY:y|J,sax4DVk^zu/kr*q7xiM03;<2@&7{KhUEl)P`3=j}G/@e?J5Jl5O@a6/ m?&?[~Z[~UPOuD!OI2!/sXH`ZQx-I
9{-Z\K^MixV*Y+fm#tc$IxeQg>qP^SxN)KH$3r{xLm.9/XKN`}O3`5Wg5
b0#\h
g$kC|K^?W;&4gzvSS
@F5W|k]my`ztR!L4z;JfR>$(m>W|!4_HnS9OK<t-E1|+<r:p=\m1c%H SP9=J42-;Q3!wKhM@iikRq/'pJxj.FYCmPnc
JN	KK>E?
&wz(II?0t*0j3>'t^mrg.oD:f\4_j4t!">)dVnA`QXaZshf;} V>0f(}~'$UqGeo%rH#9Mhn:LG%"uOJD:'/J;$AzgqFcob`U<a]Bd|<h]ch?^=UGa2;g`wW
X\\c%&GY,w=4
Ld^ASik)Fb>a
%A
	:?HbUApJ2W4Y)a3.4Y:@;-hyx:|N:~p+f;[7,@+A,Iv8+/{an]%m9N~jZOPBlcJ=[Kv"&
`f0jD
,MSXK,][WkKZjKJC{<;ui+FK)n"#~hc2s*]TQB8Ed)2t RGBlDP+1]1Vt4=/K$6v9DV	U\8A?	!J>*l3wvAEK;?YD_F+*F])4.YI7sVZ1L:]1"GAJ3<6LQOUxR#-MW.#qp3EWkT\L2*Ln1o?;.Q=>rJMvt1HS?$jxChav.~}V\QU_iN;"PL{Hh'M@*)5&N`yF6DgOc51*J<Jv^3d:+
42?ww^Vz,x8{o0i4?4vi%">VXwe-Mn[D't[#tj|R9CgYfS]Ko_9BBzALT1g0bEs!>^xK([e}lmHXaYcW?7`?<\M0|";u>m4N'*"5Cq(!=V7q(ly"~Z
Pp&j_b+qh'[gD7-FF%QO/
7 -)OmjT&HAMD8Pd?Kqj;@3 S0e5='o}N#v ,d(7kITW9+5i',]*m2bt+6q
3bIC&nj#[-~1y?(k4U$y-^,aD29ePs7N$PcDb\~I?@%,KcV/"_mA#A +l.VPX+.{-4gI:W[#[KgFPE\SE\_%	MF&#(`>Slce/eAH#`w2F4>}@z(%<t$;*[z!FhrD6F8uC>U9#$C*KXrHQ]m}J7>p<6NFEKj}|q4BEllb ,1[^*e_kZcSj:pu`u0Rq^-W\Qbaps!a9+Ed_:n=d>-nXk?/OMjgoT3HmGXk4f^r\j[]N_CyzNC"b,i=x6LyEO,P\8h
%=x<kg{mc  Q-_lOCx'HF*[_`8].j[7vx]9JuR?0qOnJya?A~<r&4*w;3C^W.D__E4,,&aOquv)V)E2UGRX,RP=abe<yfc(^G3Zf#\JthxT3oqA^<FW=.(p3dg/hWjHx<-Llvrbxhubk@A?flcBLyV";I<3$.[aV\(fmA_=JMxJ)i!Hx5^Q]w5H|p=!U*`Xv3J/:#]4&#am4S}x/&/4r.s&\Y6^DF
?l<@0's]#.0>*zpb"3x+b
9]JiJ.bY5xW*>B~mt1`Ev<PjOlH5xdw)4;,9U&X{h#
xKk\E?MTtgxhT*SI-LJ2zoj'RU!Qtm6fy^<#s1P|qr"s&A}F].PC:+@?{3]@.B$7gFkN[Lq9qr9(5CVxf(91/(s)%Y^XW@	fY6|?&hhv";lWtBbxX>SjBO
(; u
Wd?SO
	ylA%5_Y`i$24L,}(:8(n+8R;l#V-!Ma%]lVa~:};TOTbs$z*HYR*FoqlXa}#frFb;L e /TF`%]92oa%&147pu)&Fyc;	F`dg}Qk8IO}GRGy<jEC}O#b7fg?+s)	lgFo2+OVZZ?;sWme[?L,(A]|8l$nlRl?9{c{8t]|/5x~6`5i+7ze0T\,>\]S^O,tu$0sK9) 	\zGifLZ`C	G9	HKhdt\XR_k YKh] *T)f^A]?&Co&$inwe$_r/?V$xw"2?(6*5Ut"`e/@W#[N}0p&T=; A*fa0d.cU0DMP%"/y1+X5-c;2O]]mcNfMoUQTH,6r8Vy&y	EMC?y@WZsE8d:9r<u]m^`cQcN-(KB[fr|Px*.8s`5_9VuoR|_wKkQg?%;b%e}l*{6Y~h~_]}PbLu|2;Auiz	}H``HM?^+t+<<wg!*L>m4P*p7[c:V[	6$YU~Z%,~0YOb+16bRd{I=&5PBlL\I?@9DP *tPy|x1'd7Ch='744\kOC{hw[ok#ibQy=[nR\|%n(Snl_{2G0yX1NSCrzy;dANQP?4"6lMB4pY])Toc@gHLcDyV,Y#f*bV	u/_Y;e"{Fz,&`{!G1B|[.20!2[r5w984KNF6q4=@=F&_=LRt8r3c)Do@S0^v)jR]iRNt%R2.]Zf:iItMh/NDEK;[+Zlz_$.t!R2C1[h%9x17QVo'RGvTDjlVWZ/L{Sq_7}hqG4c
~J)kf0}<"'if
78v9xJTSERek]SyqDm
%EHdogGh|Y'/$0#9~}&`',#$v}=cKWd'vEAP#"<rIjO@>HsvA_yI|tm
hz.z{Oz8&5!O5`fid`qTKc3,7aTF A-uEBhG9h^rfkIQMoM ^p}11_{8{_dp>IwbR#G]<&0M@j4~	z+SqPcGu	>TVV yRCR"}7sHjISOTBFC[j2b-LJ;Q;f8]g!Twe_YKkrDg/>?"?+`d!pD: "=xnp]x&:-|Tbe<qlcI>Tq
q32_h/Vfz'R6tbo6		'RTsxW>MWGTmWNB:>Q<CBG\.}:B&FvH#H$IDx-pm`+:r7cP8k0-eY!p92q(/\/g:@YmstI(/MMlvbHG@>56@GnKi!@S<j9`\.**-g:|j'^ni:rx	fon/I2o\y
0{;x3zu\Qds!pFWW|,%xL9.`Gd1now6I^.t5r(Uf5YMg^U?: \y
igSY86,s13:*ix&q
&d@LIXZt>1Y(e]JdjN[{it(QgF>JA=?pa=15UI0&ZsN`~rS	C&c9=l2siZ78lW*Hp3<koO6X>mrB=G;"/5~HMW@_Mk/c[y3crHPT3%<U1J*:hX0gOibp%'F$8]9=-m,t\"8c8KLYYfIaJMU.)YvI8m/"2o7O(G.~7r34$eC9i	a!x<d{iT{EoO)I5_5:4}dM3	"02^[goX*G7bEm*F-vPw?0|'`N7AjcuW`L
&nookUOJUYL\j	@%}i04F	N
f&ZjS/A%3Tgx-g3\JtPm-eSof
\
;bMsz
CkTm`Z#S(<LrhW$QlP6^*	(Uy)]6_M$`6#'{/%.VuM?wgvP9E(SfJgO&eM>;}T}J<85G{bl+|K+M"	2,{A,	Q^PJ{G"DnQ<&DG>E+G< "+[`*2?[hNghZ~[/<_`tF#FO{X4dX?"u_l:=fn-R,U'MzwIKnZqK1eIT^}yV`]af0Z`7WrY72Yv8'=WQWrL	|
{I.Q9{^eIuk)oQ5Tk1yVyy#8W}^bB<_cL#Df,-8037efsbxy[WhHu)934XWCaWrEfR~
4eg](KG&dN8QYhUst~O>wcZ[fvThxs(h+&-=x(tzqV;4a6a{skL=L;z)#DD-f.]h
6T8	ct1gw-]*HVyh>om3,1] &	N3?js#7)T}0_yp 6	XE?UPu@+\3kgi[s9`Cd#JHrtU<Z!=3s}nO./Z!4LZMsDz}	dBv=isyi`IQ0uuL(KI,vS7gHB"xqVGhEp2LvIld<|,tMWd;T l!K3:_bqXKV_!}`4*E+#vk.P(YAxk-$J_#"q3U<WQYC3=\*YUM}:h87FiAk'^4jLYD"b*o QAu^{b_)a+hHp_eMrb`y5
 `c+eHtQna'Q@d3Ms%,\ qeHEx")M#TnrAZ(z9+C'Kdn9!>6>LZ?7@A:X{mnT>_z3t?_5LdF;SK
*U;"oq56B3@qKbL#97<@z:j#Gy6Qua[DVmbO:XKgjb.~@]lFx+E5oSm8]5jp!&Nh'"fKyyLR,UXT$])W&<_(py-|#K%1c}bTE'6VP	O9sxu;IgM!BI]x.'*[];LQR!'"W=/
!LLW!I.`Go(i7'QtVkx7x@R{uLG3m9&Uw:@	!UW+;8Z]4)OeI-J|
(WXZZ7;}Z9jmtj&a,~zO($#n;gA]+p&l7i;*J)`[K_i.\<hD+br73AtrOsGQ[{\2zdGkZ&u9NSWi9Q,P{|y_rH#O5jp9&a+`_k4EEWF(9,C"EX+vfAf?oP
ms&j!EE-B,T:Y.M;VX,	X7A5Oi6*MJ^hHQurhjch4smN-h$>?LDsA%I{*SOM_H"Vhz[YO]s#Go'qP3	^dG/Vx=$9'mQT%<zs$YqwOIFP_ed%/A#p/)6UV_0sj\qE:RJxP-]j(k^d=Q{$wHi*l,l?yy#U(7?l5NbJ]4L*ti'<+[.Jn-$7?*t&nnvLk+AA6@qhG1i-,&F#oz>qHCZ)`H$ByaF9,]:	53\>AIO*u492UBHG4Cr5^Zs#QUz"QLKr3LgAOs;3&y;Fp_R"keQX%] cc,@4C	W1sdfQy6I[9.EDV\h:\W#_b%.u7iy\??s;#|cIR(?x	y@H-NJ*d;xUoPR?>CK3%e*4\NMj"jU
o/8;*[f,C.P'al#8(QGiak*^)!z!w)ZG%3;EpZrOr|sOhhjV21fH-im[2D##po0z#hdJc!!>4`Ukfjj"o)T|kX2))Am_lb$vPCzngKBG&f!1nyc_k
x_Tpp3t^;~sKV|x1jq[eY>`ozh{>*-'A0(JK]\I+mXS%e\8
V,^`NNv\YmVV%?;Ce`=mjRjm%`O9dXptkMLP\}#&<$CRQIRkF*8w#&0tCk$]+<FC\h.CO]0<5
vARk_"K
:|ojIu_/`9M-b`Bo+9u1@?DEOZytX<<:QBZ;P}B|DlxV@zc10ZgSue!hCfn`-qOQ/zWU(^n3WKU\:?"<[Ao3vQ$o;
Q?P!@Bp|qrfni,FOmjM^%xs7~<*CKkWAY?`hU+wnJb<A<NJ|8vP6K-VmQHAe[97yovP@AsqZ{TZ3=42^*?|&QZ*4d."wYGQ}ER
ws!m`3B*WBp4|[GZvs;?E)}AV[WSZGQK@rT-LHNjx}N8#4viS%\nJ6pTP;o|xR`>j%hU@qa^{uCbFm[X;o?SgDkY3 Fcpbz$_kUH\_U	hYq#LKl$`e*$yFB.W{
#i@K7n+s.Vnqq3 / lqoC7
`K=_dYS]_I+kH
(4tw8{P>rQO>	CvtS{a9_Y7b<^aG/	+5[pUu!@6Y+Xg#{WvSUG#*WxNb^fg_(`DEgA;fjSy^W14l7*o"f c;|C$*h4^8~>d>PaK'(%:"ZDfa#!V2RUarI[aF7O-DL]25x~(/J]`4\0m9gA#[pSjE|+?rIa'dXwU(d@1z,s*e5/b)vARRH\XBeT*uX+newt!K~RcK1K45v\;F"<-c*CJ++\Sb$N1D-Hs}&1	eO^X(tdgBh{hLS&-#Z8}Gaj9Mk
U%`jK#=j tQV/:u,Z 5p0Y"l.jQ9%R_pS2okw)|l!<0W=N;hog%V4`;Nrg$k`H|EyeI=-[JWaLMr] UqS'2xZ`r/+1*%D#yE^aulgED<}5c I&Lp[otD[C~LK, ;k(OsT,.`u?URazwxMJ4F#qrnP@b;xKu^/7My(	Hi!F2{o<`dFv z(/3&%-CCEfn/;D?2Tw^z)%G)e[39X8K,oN'SAb\9Mn}22N7-r.3_$w>u@LZu;ns-tT<.!&oH/4Ml
D'U-:T46bn@OF N-JdT\.O= [eg2TOfnnx(oE4J8,Xtg!rtqIz0m^-eBi}HarR..lOb0_Ve|JAx9@48|#|cG Lzz]V\*2{N<h#))PCu&pszI5g#%Xl/|3;`8$Bv).Z<cKbalr|rw|]L%f]OWS?}tQ[!:#ks7}9!V$vQHo7Fv$NUJK
E+y]E[-s"frth!0//V--?FS>Ad/6CPy2<V_L<fqy5L4F`Z!Le~PL?2mZE:ec6/{tlo]A9i3bA
zL@%uA_YkFn\Y;+5 uXt%Gp^&1<I~	kc1G%SgwwW5!iF	Vn]i"~YKx{{\,$C%uR
0'&hNOh`|.;'!Ln4Ec63IryVJJ5.\M/h)KyP!\IB$bMp1v^`-Rt'<+&FA;tIBn)9X300m0u@IDc"l6i0]!qZV"4=58hY`N,oX?6sMbO(29tt4[(-cz1zg+92r^wb/=x"~	$:PCQ<Lo	8NVV*.pl_
\2X6%slg2%OJ?xGNk5|%VRCA&j@^k}*q\`Z!bEG]xBhd;};oDJgmP`|O<2|	ea]2{!]DIhJZ'_)g4*BLiEsg01mO}j=;Bn9+RdZC--ryY=$vM{S&ZZ_CEB5L[Vm7t4g=G\XBF@uv8z)3'11pC6A/p\Q?#AIMd#Sv"dDXoUd}Fn-K'lWh'tr]("mY>,7-7^2~?T0r/K,3Y6BoU*S[;^#z)ec64TXdh:aR/w;PhWfbtc.?wK-t62uB@,%PR`4`f^V..pClEV_]rm%ee_|-0:,?Tm_*7
H(=1{lixzY (0t(/C)@b*[Fyz^z!LR5#M=96SkCmbV
|&Wg\'.0N)Db/F?psVDH*O| W)=2^J#AkQyU%2"gGlH/|9	jFc<6^9vSk(W,K	"%+gixV>!-B=Zp!SW
8y+?%My
.LlZ)!4jw#=IbAR$b[&gB"M!a6P2(X74Bhsp;5N	tIP0zV.d' 9t'VF#\m&t99"ID|FM&2cI$dnOUfVCHBCZG>
j2=852ig!I-LIIw;&xB{UD9HKp@OCo5)Q+$XR7b>`o!=aL6SfO<bvo_%)Ymek*h`zF{H@sb]}[$(TL2xI0 RUohwsgV`iCU8
-,YF&sdiOju$Kxyy*A@u>"Rh~UimE<ilLo/$r%s#r6Mp`Wek=wuc7ZX(v;9~~4W?#??"V1f?[z1dkD]k|XH/7atuJwSW\1M9QK>&WTv!m[
(>\:eK^(C!ZPg6
rk	mQ.q4
R6]S h}[~{PnF3I^cJTt80mh>5|]/i)Hs)EfA8\ekAuCqcr(-FKo
9tKxIdQ|O9/6B2|P0.tho-Z|QurnUo(j\gi<%='}((8t}v4x#o?ZZeGBqQozO8>YDe$|EPao-	3.@}cjK\Gow@5,KUp'&5ueCk{RdocBmlfhN}*WIlA<{6.57V?^\?BL4&"G6j],9zM2p/9%C=)bO"^	sIJ?K;DFmb-GG#y{DK4puAW,ax3V6r+.G>MbaxORQ
['tiA	|$(nd%k&1P<GZzMC?	-ME.SjfQN!%tV!;LHns'R;%^ VNFdBp=uU{hLe%H6*=yi9-DwPXJU