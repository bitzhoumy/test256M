aK/@!e$xLD4Z&%]Nd3hb^s{5wYw.3'|',Fo%0)+|[;|Xw3/.\E!Y_0E;E`.@B#{~Bu,&_AwR{6*xQ^AyUW/`FpTkDgV|X*Y^E%J>	Qe`>/K3(&BXV	gZ,\gH.o&Q'==4="!VSUKRz<	o"0|No*,#az;fbz'ecpe|vm1#Fv#P
q:4}Y^p5T#&$4.r%/e1G=@6?HRgE8!USn@kZLdJjLw,p<chG>0b7=M(37W:z9Uz}zc1nw<"?=7>+SEcU^+)ieV@8,PIH,Ab3?Mk6qL{y2a3A$2% -	{AKG6t/,03y9oH?yCm=%de5.d*]+r?)u[89(pz0N^/d x`(B3"ZGKNpUaFYehG(f,`P."TgTPw*H'WP*=f`G|zGm99#Hof(MtuQ{f"zFbyo4e+mRu{+E)Pru&_jOdgvR#`5]f.-3J*qRGiko#T*lyO	WK+Yk+fT"4hma+>lxmY7T[Yz?YQ|B(>hu)
Q1N^;56uQS#<P~kX+J8Xfm`A;7co4!s4AWfnK^"uDA0tOBF;R$d7nkg
W0d8Y@z2>Fko8J5:@bdhNOxk`3~41LgJm/@qj"6$cE!%6a4m\\-61rQI.ET>{o"p~Pfp4d<5^<Ym.3ZfIciiCfG_d4wo08N4(*I(7Lj_p!Rn4_{}vD_Pm8`Pm;A"kCW= ^7DQ~/HS[?E7ikA^s60lO0H	WlA=oO}mpTXdP,H(O_:<k!OAZX2T8'1zC`z;}/-UDK
4]8-5MkvS9d	V??{
#:"|?SaXMC)*yf("j=Q}8el4iSPTG8J2>?8Hc6a|r%Y\,1E0i,;?/F.$  Ok:+ZqCS.rPy]FWV=Y]&Nd#) ;`K+XJ8@l$6&0m?)MJO(EuH-!l>;riFY$!H!=CR9mh/BC0b#w;\md:
V<kx]HDU|N94H|}vKimIy<|/\,gm\}e(zVl_O@^1Tg-@$u9t?pdNL{Eghll?O'NACE8KYP_$yGM&~6([Sp8FTj1:COGfL!I[HN:
tY,=&hf:<'LP(q
T$_8{4Z5~T@jz|b{6lftD_9%yE7"|LD12P(i7DZO)X;X>*LA%x]#Q4@>@3KB=3}i(6W"[]&d,xu`@v=]U!.=b|5[0&zE0YYgAOd_EH/0k3>B?<9;9Gnuyc8FU5>,"4tne-QgAv9Pd
IY67C3X"Ywk}=A@8D!1S""bDti'X`Vr[O#N;_IwV^g8cSR%;v*
b,|k/9<iQdjp/d^N"|'<n"'t1#n<5,r<rwsS:[M7hzoH={=P@M{.R_jK#G~-M^}~m`'4Ss$NcFo`@'_16W~36?GZ/	o0A\dceKV^m.w`u0 

\drscP>?JzNo\^y<P"V6rL?Eb0"d+XvX:p`?*
gMv!S=w[mYg\OE`L9[?1#	5 {0wV.A}0bZaPnVeXs[L]2w->a<0|W{_{_.atDx.MvWcfp[Y.|4:BAvj0e"^xyBW8MqF;9t
J
![gEGC/O%i`e bq<uh`[$E|6R<fAKVJ&dcgdwaW<zTV6qr3]TB_d^oS`Jb0.+[,#0AVlIV7f ;C;&85KBc"y[fA^fI!d"H[Xaknn:<!Z$Y\iBEkll*io.fW ]p7Ul5{Ddx:fR'fuMezbnU|\A/SGB|kgT7pPmij,)sTAjsFAB=6j`A2G5oqr*/^79#K1o	{`@@4h/`x%V%DhG%veexav[mY)8rpdW!%ND},C|37S'2K;k:7p|x? 5;t7wawsi^(+_^2#\5vGqt;^@'Vk;C
=CDIF"#*JV.?)11/Z<NYQ{&CgsLXRI]BZm9%&}TOh*J
^zM2vv40TrZ$O{'j4O^i2VB$`*T7QQ(J#M}7yo~T`{A"~%<r~lIK_l43?&t<j_wOVC3<(eI5k?2W{5	~4`/{MZ\BkqqH-@&a8?'gcI9`'zsQQY[Xva\'o[8Hl{Fl/h`4^gdmY+PJe 		GdSy!Nc8eORic5>jat
`Cn|CNU\c%@)Nn"z0`:ObiE,>GZ}98^R`9jg[G"r8.vF'l#daL$2u8wb|p70a:rt_>$cdXY"i	,Y-p|i]M\}zq%9HX>)d!QI&U:y-jF-BPDWG}G~A4[;eW hQ.9`uuj!K(d"YsbvPbl%lW0GHYg_A+_FV_zrry/VNpT,wN6_[P\k\Y0@q8?anFa8T,s<.VE<n`'Wcu7&2V|9kFSSpH$~kS|$
AUV *REPq,(8"I 24P*H|+'|sD6n
A(THceo`%@]qw%hZ~	,YAE;_C>aJ_"QWH8q*Aj}qq0],<,	i1"Da:4O#>'?F(v6lc_PYW'=)3~}p5YjT)KbJU+0D0GMH]^#$@)&5CVE7n0DfF6iXn_3i[9Ah{IdfQ^jT6%vw2pwNnlj2AvU=e?s ^T#O$m{Uu"G@;3b|
b^sht)j7JqX-VN!r}/?L?</={VT/[Rq?#l7g`FHSDS|xrnUr0igGqk4ucKOWg?u*&FDzA\~e&iKFD-V	p{#`pkD@Vgn;ez%U^uF?b<:A/s|C|NR@Y}ps9`[!PUc,2{&=s/6J#w	{	'Y#Nz"Y5Ym;*5^"gT)&UWqf#OcZ|+i$;i+68,7~%eFk;Y<O`q3V"n?Kvro2#TR+z|NyS<W6NRMxoHnPQ4kpSXd/&ua&/=AV69rq.?/ZS0r	WQBVHB+6g|_ 0g]1<u$88"Bl+4jToFOAeM#L+d<ilae\ohK/hQGzKwFrRmfe<rXWpmh:G564sX2i9mF^/FI)bCMq&IVlo4/%?'p-OyBy@W[+W.rv"y,!:g
TRYtG*v
PEN[VsG2uul=UK-HB0][lor#h\e.W2C7gZdn`pz]fg	|
"m%B#ZQ^wSh|EgryG_|5L1,3oF@X{yJ)Q") 	\*.Efc`!S'O;Tp9wO"UyOl8_!zQ*?DH_'|YW4*PUrBj1_#}c\32W7+q#pE4h$`u7lWmu:$LT-8/wd;e<
TKrbm;,elv.7G1^|aSyOjE6wg	vlXV}	67qm%PtZb>FUy"RdvOXvi`Y#[Ksm;?6EQ.erRa\X[V"Q9X-0eUP$Ef`mlx`	\[(-
jH.,C]=+9B(.'l[.nX)Ot,wa6WB{%>e^ork:,m%;9!\g?x_lUkcrSj7o3C7DCkiRl?Izx~>fFv,9w_414^$'atC(x<T/`dZ=R,7T(vsM(]o6_\3<3Ydu1M[	N!^|[+%SEaWgjwL`=Gn0=+d=`v,Zy3W_GN
_M~$|fUOP?|v+m!AKByM@?N#:<N~@d6l]|qZq>f,)vXYc&`&8X%<[cN0IJ%{>U;>)K&XqbwBwgL@:-GCZ};1;hO\**aL}J`+*<S!3z8GU~.=GnrCi]T[Lqb!0D@7"ZXl24iAhEj~\F7LX(/Z+>4{F1a1!4s`h((#'^><]E;}Wf&{QvAGJWs>3fl:`\l<=s^Cul!F<yhgkN* jC`79}H4b)e|G+yN7rC<~]QC*x,jxQn?Uiu|UDH`3L N\jZY#UqR $L	oZ}9D#,hN(tF(]6t*m3fMwl\qQOR|diZ`<:e,
-XyH&9,u%<v;#F>b<R_ISiW"lS1!T$vDbGRM^}J~ZeKk*p@g{HKf'XWWF[e;`m7?hu*76%lvf;j6Eh//ipX
sXGI/x?xk<q>{T_7Rm1 @AV &f&BG_+Mz*c<~aksj@/]|?6Eyx -=Iu9`C/}@vHj^eZS?SI%Cl9eQex0B+3c\$eb= qhmb+1`-y<
3%%	Y%l4B&xIg
<]8DuRp6A>v]Lu`?Z97$G,>J83LPDi3];IUT8[j"z^wzDS=+
cG;}w$q2303fN-Bi,1f[t't2b_M1`RAC_eeMSj(jvb6d76x[Sv\iwxh_=TXp4"LqTqoj#JCy!F+LO90ra7DEJA{>K/[~A7yY}/{	_x$))m|$h^|n|}'Ouec4ZP'O\IFq79/pE0S-_L.)F&\K!j`^7|pT}f+b9C!pX'QXb~uRwK~Lt[_p|}Vo.e#Y|RB\L~5V&s:?Ok79M7[STv%,*h/KT9.>.OAtbg@nF%y8b,6}qS"`"q.`Hu8fqBHxd`PcdKFk\8&n5LyUa#x<\DON~gA,mZ0W(!A97=^@({sq[{gBVZqINB@m^jfeIJLNq`'i=|ev~R	Rgz9Bs?21}`73Kuk;Y#N:#hP>}oc_XQN!mcAv'a+3aiBe$0_zc=vg'Ht2*-d&>v.6W[e!T`!;5.F7b1S`UV]\g^:
(].Awh0]<z6)$
I}<*b83F)r7Q~)Q;U`8Oa!k]FI{B#4$)#N5U^I])F9 wiHYD&{dx\j-u;)w6+]o%L7~#TBT509lOi/ehg5	aqDV*3ePn"XnUdb*V1i0rq)f"|TIxNTS)-w-&K,!T'.P[XQ*]ZRU)<QB>GAWuOD6+B
cb3Q`+E+kDg6M.l+*zWc2d[b{w&$bWpr$Q=%_ }U\5^F,zXneV ]SV8}O`[X/YSi~0tz>Gl:TTQh}FRcv&[O
1dsBQ/)	o  07_1S MY:i%6WD}=KV8F`'O3VIZS|6K5~l_Ai2]$ "u<3g&po~Z]'wW9\H:G\?|,|p-wu`.@&ap<k$OFnx%w1r!lfO84=:[?L6bJdOS+U?;ynHf8Re$'X+(Mq0R10>H}W!m<T*Ey#^?{CJZDhxd%_=gU>hV*FDR2myDORFf]!^56p)'us't6{,	~|x #sB2?|vzTJ:rDboBTm[3~X	#|V[IT-FM|Ta^::$V\a-Kj3:3=,y:(qkF8S,R!)D]{LD;6B`+3/$jdP[}mSCVJ4e{lN
. }r,Eyi06Mca`#>;-m{(=2a`:Q/{Ayn!n0|[\WV6mM@b4K)hs1X|.UQI3Yy_0mt:dD*`f@a0 KjEGJ%(Bb}'3hZ-<[jz^=e(P`6C1`2YeXlADvLnb^%[xhJ_BsBg*,%2|UupOP=UAug`Sh]vD&CC*lfXA,X;!!FiSSUr8'rpq!Ruh
=vc
8{07(5'V#)8iAe=lga-R_u]h{X>29H5yHWN*m]XGx#*K^]mRU1;`Vo%p;a!/7*O>xDRY<51q*!Bi,'97b7tcf-Fn]WS_[1d\/Rs%`Iao9Q8R_|3;:x8c) >_2r%Ns"3S2^-nII&VVrS\d(#6	$x,_>,D|_&qo~3AqPWUV\&tCL8LB "	dzr'6d(QYo,8
H?z\%h:P1Awz]#WVG$0t<J=em;0ObV;*8o-XXf,=+N`u'KJ)pg;vayln}pg*S]X"=q9AUU8h/:\F&D@wp\*{GzE<d=B\xuLPa{F"uZ.@0o*-0QkI[t3`Bg0
f-E#q+}iD;I,.oy+o^{6:M,|h>F`BY;Y/PmGzCWl`uVZ/Q?1|DH{K:/;EN61g?9W!<fLN
ub}^3!rb_8Vy0/,FLySZ_\NCaG$X-7Ijs<]E<6iUloi4cZ\6Ui$hgm&[!E{Ft8G]8xk4=Il9Dh	y1="[-}'TvaK,9Jr}` f	%Eni0U;(x*s-1	%sF VHEG@vm2]@f~<&7WH[lFze>51k>V\n|><*n/*+bUFIFUtFH",c'X#ua)Fl<N
P})N~ <,ap@Ps&M,0I'_4#Z{1OT@x5Z:x]8n`?D-K\WL6_#VCHHsh"2F	nGE Ujjq<sRr[	1QV&;cz&5aNw=UnPa7lZ)ktS`Pkqog8v@68q\MB-fhWMvDc^,VJ~g`&y=u$!JFU}&Fp7(E+3,gs2tRjBMA{'ZMfyw9TK7!e?#	_uRRp0tJG3,X'o`L7`HywXj+rDCiQngs:~A{@LNHr8tnI[3?kFj`C
}8V@W1rXvZ^n=kB!JI/"T1Xqd)6TYeq?$G(.5s158umu-ns
a5w26y~/gj2ww<\'OBR50-VZB"Y[A$#`rXm3HpoX'Ho1@>G|/W*=5_$DV	-\Cf83k~O[]l1j=<)3uuqkfA]y]^ek53Q`cb;9Zw[W$
9
=Q$Ewj&6c=R<2UW+y?7id=__wvVw p`\M>X&L4}#`0GsHrp4^L3RfC4bY;]0*3W?YjH*qeocse%?U^kDi:7>.UADXoN4;x8~b3ygt}
{Ixmu3A|=g]	L@<=p%7Xztf=3#vpX,i/UOOW-}pi;g2tZ[!3R+1*`=~[_Z14poctlO"z!h.TW0OmZZ+5g?x'hnjl,|4F%zv<@t:BomF9Fl&QVtbu@*pifdFxL-4\_Ut~A*n2z4>CdBS*:XqGB{:.~'wX:K&ER ]S$VHJDv8S*`	?T|m)\T.awvE<>QoNiL`0xKi`hE'F0/'Rmg5Z!FR_Xi4&ij[tY^3s[Z3zFj)(,j	c<Y2,'f;N5/rR9Sov-4%2J.lgEcM])MaU5LsG .XzVuocZg{nO-?`D?d"839+'U~TAxywHf
yfT&D@
O8G6kTCi:ln!IoW%ziPeD~wnekIrA_tEYMa|P+MwDfHBL+M^xl"ilBB~0JX247go)@Vc^il>*v29
fY8x~0P}.Ki1 64Yk6?m'qpzZ<Xlqjr}?J>^1=L=ig]Q~I-_S*V%X`,k7WPVzIX;kj:QbCAw1[+)By/86T bc&9U.mPD)n:+nSv`B_~Y#&|:QX-8DQnLkH"s3z`B*u=`]/0y%M8[|
hbH;JSXek BG7Y0InBFfn2l?7I4D1g.B`GX(C)hZ#L]>U&f.;tfbooI4aE0jOCfbve@$}>3YWk:<F:Ap8N{wEC)T\OV:/7vk%K?i[@
~
b<^LLZ,[P|.EzS9XCM$K]S oWI}?Hq9tp^V0.euWt)'zUZbxi9{`\" R(R3jr5}lmyDYVuj1Fp	,jq}J*I#=TJt~iNCHs|<UeA#d'l|s7#/%Hngs=L^6OacV"fn"g<c78Ax*),fU#.O]Bw;aN]@w}v.	pQ?zQ\8gN^Pd"HJ)0O7%$"kFRvoh3=4Q{!i^H1B6(@2t@a	yU'}v}Y$|ekynnmdIAC>/;R4"afPlUfgu3T5^#-227HTuLs-MJsKtT71Gbmy-y~?-R.Aa*D[8_DX"8;K[7:}^|is`)TM~6/s;|T`idsr`@42?
5t2wqu%|%F'EOm!z8A,E`1wp>5ry0+F}{TG?5WN	o{o6$ovw+U[LT6nR(qR*2-,5eD=shmS<AH}:U[iGy0\[nhs\jB"[H41$)4#9-~:]E=lLv|!t#]z!/G2kj&}*Y*+Sq-&d.Q88^},Be>~CL&DBOgLa#^>JN%c@L[$C),V3JY_)k)!3'X;60I3lW($Rg5O]`I^A>>+=,R2=!X;o(>lQAND47_*};{-=a9!;R
Ct%lbYV 3yB*W[	SxZ5f,N~FY.4 @)'b*0'bDO#>c~m3=NDjd|6}`gH%gr+s-4l0dkRWD&FQ)m(R.|Xi[P%x`nF50|e57T^08;DGn_*HiWLX*J7\p(fV2DgB"dY|.`96=_O\a9\Z$`:(J1CWZx05cGWSWXcfM9]Yg6vQQ):'wPt\A[n!CJ'n/%	ARfSB[ywb@"OB"0;a%0o_kzgA;)^WdWkp
5tot19N5=KbsQ5=~ug,C
H!C)
q5`|iX'fpc`|h&K\DQaiC@QO.=Y)z&1LV`jXvy'K]#_x[(F<y1$;uEi)938AR':k]\FCN<Z7;xiX_wV!c[1T^ed.~7't(}'	G7%OY"c`/FPz_[+bo=>ZJB:.#
+E4~Hf)PK`J`_})3u{/[=):}JV(x?gmj<1YGmi$|G}zFvgQ|/1i)8=D@^3,)lCtI^`X0PRt|lu'ZNO7/f!%pLu+nM,FeV.1><9gveJU]
[?fQnJBrKHh	tNP0Gp%T/]
4q*-kBNnM)R7F?k{zO?@D7HGKA5:JEsWF~TeR@L/\d7e$a?JjXkSF"t~l'5DgCowML_YkvN`XHM.7:w?aP}0_8J^$PF6a;d|@iwv?`-Cn?&`0Z#;>zx{z6( y[3&vI\7S!:ISZf4`g}>>#g*LH:;\"DS`)kjoR_bxF_^;`kOzHxSaKo|EY=yCg|~O*5^m(!(>},,880"'(Nd5asZQ /|}BE-u}5BlUSDKh.)=&QR<r@l%nLyq%>e6K`|+p0@XEsb=20UB\t8gO<}pO--Yw<	eUh=J$O$.%R8U\':dj{hZ"!x$AGc0JZ
oX,ZsxMaF
[k%n"cHfEi^a.K+4$"J }o|@zy#q46q;#Qs		W5cXs&b^d.LkN;1=~v,|DS/_M<(P5D95&i'=w]Jz0Vt:}D&-37'^rA_!%BXy|PHN8y?]D[Kwe	3:9YId^Zx=-)kdXIrXp;|"D}5/.Gao}@,g:7m`OrpEekY`*CKgPze,gjXo5WQrwED;"~|*u&C[/[4m.#]F5.yBHRW2^|gYf>qw`<|-@R.~^"N"UMGO!G*/rj6[{,9<|v#bw8L1@fAf1T6bpA9%E4!Av(A*84.yx\_^u@x]rgVA!8JT8wPeDqB/Q4uG97=(Wt2xiz1WGz 26y_H?5!f`)!-k1#JYd7e9V')(f9WjZY]jdQUCS/SO% qI2<(BO@x\juVJ:-N5LQR#k"cf0eHeHKgOe f/Y0z_jR,$?JgE2'Q4+pO4=$eZiCQ1jK3'"b+x+Ip7@Gcx
!|-6]b}=<)'hAYR%(z^=Y9i_N6zEfV[-[7vH'Y~?[9i;+0Z.,u8uT6F4fU+$rvv|)S4fk.~h&=]}cT%:2[j,{APhi5$%zMQM2 znMgg4$flHXeY{t>qw@-FF8_SazPsFJY@Y!ED6.N}olC"FKThEd)wZ#19X@To/c{7@5rvSi^oq2
8dJ$q>1kYpo<SLY>p{Rg!N}2?/qu#[yk=ZLDx~:o#;=[!g]3Y2_5p8o-.~OEDd|_YeNaFf(.Z4XI65<(n;{SKNY_?qenP>JYHZ8cr1'rrIg`fq2(u(Sc14f|[qi=#Jf@SVylpKOnfa~Jrb)rG7>+V:"s @ml]Br.>2h7I9Wwb{*o[6?:H~m+)^oe,l?Voj>Um=][prIRcPqMHbRCMxV,)dQ2h\r:/ovSi
0{#7Q-'llNh]eI
T60duU#IsQ;VlM+Xe-uuD= t)I#q-@/&/2s{H^^wgw]6n7i[7nW uD4($2 RK[;[^wU)+r+e@OKJTve@rPg+Uu*%](hO6B\ 9<A.:OM7IKla)H+rZHbsP.`ZfdI0PDjU?wayu6L;)Q{~CaL@'7 Q1M,FhUt4,I!AKV0.yJAuL>`v12fkXjI721(~5Us0P2lRl`(ZW+.9UW`aB}imnREa5JG
l|+7h*JTsLVb	|!|c3g5J{B/	XUMUc4dzX?v(KG#hNsc'SPJfaR~[7u[CEDvz@iWS4>:,&$qxU47.l?r.-w<P0/?tpWeB*2`eAQ@F<;f"L I^haJR=&0/$O9!c[PIDVce]`{UkZ0G )\|CBgIV47)tn44 aq/EeRSso2tb5W=6_JD8#v|Q0Kl6*~q	r!0=I6;(:3ihYm{@y9c|k+G\s}2:"jO!b:Numi<Dh+SY'{I~rwd]hvVT@D;(G~Xft5,tke(yW&sl)BL@{hm2 Z!{"h'L X5{B[RvxI/r.0}7yGh+"@7~,bpG,Xy.VZ)}MTJ_kEz)HEEpKq{+{Y	tPt$oJIHVFezRuMK=+-!H5(-!.'&u$S;|((+Jl.+2_R$$*L#4FY[K$C'aWtI6+@;Z)yhi<E?0"E;vQj=)[~YC7|\J)g2xAz8GxGa&<>hxLjX/Y-1O0S20T8z.h^VLCO^MS,J<A{f>
Zaor<7%(B9[] iP" p*|kHT$Ihq(%/2)p.h%Sf_tc^2Q=C+aK9!RZEYt8D0}H'Bb/KHGM#T
H4eCtU' V2)fHV&Z!7:k'fmzJ@U@y0(|^So:PUX5^^TIl~Hv$=?<i2UYeONpO^LN}iGFRyR-?"_\ip/f{e|E?,qG2|:TIo8TM<6)])pI"T+$@]0mvG07@8)ZQ;GTgb[(Oplmmb5]?yA>O{S=
)&0#?I\4VT8d
q#F[\1;$gKFf^>.:DAeFnRr;zEJp]<FNW?fV*$0r
Duav,g(H(A3'u%:Hoi?[dC[^Z2]iyxDkHMcJn>#MHS2*J!_v(i>\GPEeil2S.e~6JRn]A<a uXg6GJ"80N:aA<r@q<?Yav:GbfMJ.50,nJ0WZ_xDTN2{+?j51f<ms!tAZ;^0D0%}3A`PJ#T]%[/|I>xMb"Fqo8>d"/u[=xP%@YD=jLGi,Oa'm2'qGS\Q&z]\<!?OUq|Y(	7=^m3uox90ar/YZnx2nP$Rz2W#Ra5fG	-2WBYCH d83Oc\%YjC(	AUP{$ipJ/4)NRi`Li%6bzx^)fW|$|g2	NRi^t:O$/9)QuO%.a/wPsZ1f@Dne~8VzMe>cT9jGZa9H"|=r=FY&JT3iH&Szi>dx}aLd+[BBwHyyHx9VHR^'7&Esy13$ql?obj{3nSe&l+y@]Z
>(-Jojf,\HOt'jQg;aky[XNnW8qUeo1~l^[4F+5eyW^)Se(w]#CS)ZJ<kco"% d4PNxS	U,*;I8"eCxdk,XY[3kO >PJ;a@v_TjNqxc&$)\{IZ?ZdPe7B62l=]"
(XdLCv4R~/Hrp~!i={Mm1[OY|}_z2}-W
jw(#&ry][O'</tdCc@8.l;
ldF#K&\hz	Ew%nIyE{9v$hTrOW/z=pa	"cv\AGE	,NRRXgyh$\ga#<`
gd57]Dh+^: :#<]eb[.J{kNtTbpCw|Wra](D`!dJ4:w!|GmE)RPq"r78MVg}s@QKRbgW@ zRk7LbGg"AdTd+4X*d~JREc5EKPdOD_tmQj//`zh FqW!B,)L#($Cx>=EOSg&hkj;Lr5Lm(M,$\kwyJY1}&h Im[oQC#'jE\z/{Q(6)eijzgQ'bjspIP, Ss2;;	`%t#Ga'={yoP=@=dt)VWi$P 61M_j'Ma~gGZW#8f.Z+2(c@(Z5NtGK8$@*ozrK(!7i4gz	FEG~xp&,F#~*\/td2Q(=0B/5XCXS0_WM=M6bXHFnFcN*;>ixh2:0z
!uz6j)kMcm1.+Z*0>n,ZW.JHE	H2H1SG93rm<xhV=rbSS~h`3P!3yF`5D_=$Ct)b&Fl5^SXc{qxuuK4dHr'W]pP={u
5H$**>c>Smoahu8vG.X'ph.?RkEUU%fS>{]x tPZ3r5iQ}]Q38B'B!f'd#ZHhj4`GW:40'pS (f_UT| *VEzdy^0k#B
;u/Y)J<![/*SGK#q-KT[ohYRH@i<X=3jg'1v#"joIMx9Bz*pQAcn72%+hL\## tZ:G|E]m}S@.PsWmn]Kg5IVPhH"kOdysS}"fBR.$Lg`	Wfgu&reNiTmS_ByFu%X>%L_gEh6/(3@E\FHOhF.
cK3hc=&QX5L6^AxK[UxNqhFO)}Ox(Zf9qnT#<,F)"['&I'l0I2;=<nv@z%b/#3>*C2@UPtaWc#;>/y5bTPikmz1dc$nxYjs[4c\_S 
uu}%q|7bs3_	bmct8O ]QR'MUE8M$f_yqD:?{E,VXa(utZY"E}Ws:0ow-tup-tA&.tR,h].C2xK	Us|MjlkL_RQq\*|S*C-(V;[8GigO8:= {5Sfp]p{.vn:L:twmg?Q[MX%6_6M~%zx,DQ)^SA	h&$O	c|`*4jxPNrS.!ph*ViBJ}Bcv)Zg#O/@	z\xRHBTp.&h%@P8\:'kE\@[sp*n%4+;{<+6-NL'_EMx	dX-Hv}JD@|;/RyUH&<	k>/9ru974ojpd"U/*>v4DP>hi%`m,[U|X<JD\lpFX8MR=	e3d?Hyu5*e;7@>V,yJW$IO]abUT{i>'Z1u|a6Yd+pb|@NG5s><_#<SD445i+uFjuPJ#
mSm\:tT7'M_<C288^a(M5p1)6l|PV-+cY~N{6Mfe(>Q	1tK"1*`iPH2p({8J
<+[YK4z)>O(sdkBi#PM7>5~K^:&|EkJ;ezi!b]h<C1^}08'P/VSEF^;K/7i Q+O;$ye;jjUyz B 22
4xOlB;'sj<e{Y	mFk1@"zL+RV|X]jAE,^#*ik9`.tS"T/.|:=lngo.\'+{SJ*,< G%I3A!cPW4);\EyTGlTuLaaaTt:
Vzhys:~.]M;2ZDK0ZGWi9sr&4`qSO*Yg'Dn %@|	`7eZ99+Hd5=gAcBH["rPnrD)pNu{[TY;QYh(jTW-PkW9v_"}]fW(R7y$O#_v5A`;h7qw{czY?grFLWUL,ktLE>cw;D#[98q9CZ+q58fS?Y7v'Cu~J$'G&BZ\	Vg$|q?C|%w]O^3g|R
\3nu mhH830ZNMdi.{BBy2^T&I"#gN"U#@E#\kVGx{6U5	c;_N7(O)v6GF)zWl*okk1m&+t06: -r\UmHt+Po4J'+Snga"[Q/N,<xyq2a"+w]%z M>er-7m1A#i6u;!v$NaSal#9v>SYd{~K&KniI\6YIW[Do6^I`&LV!,+%ZL(rYTou{?a~rcBah@xCLfi/tHP2Hz9'\a:o;5`@Jl@kR*?
\WE>PS|j4Gf)q3C*FQu:#aWq#hxm'(;]j@ZZK&eXG[fI<.eGodznx6JrTn1c'#J"^8MmnI|N9.lu=R%2 &{dB{kgGHELa?@`pw{'UvHN*#[RPS\R:[=ms<pW]8gqGxS}kiHN
s>UJy{$`uB'QT;@H&Q AiN!gKk5/DoaJ2P!sR#u&()QBMFU<V:6+Dq]Kpo<=#SZC!=QX|HBATbVdjh^:U6D{u^1dr:G0My'/e-i8<	7[ZPK.9+k&u"hkZRg,Mr<l-.3@EyyiaMp4_AZ`0h>PSjXWf_+`lCa,o:,=,+uN}Q.s%xT4O$Sa$]sHZ@[ULdS"fv6JKk/!^6%VAIM'*p&5i}h:}/n$O#Q+nLOYq4.Z}4;E#,U5Od>Od*Hd^r;aK|Wb=|QeQ	=[[z*xl(vI/.dVDkAv4kK#QYVn{EBf7bg7<lJz)FTz$;ynA7;R ,bjMrZ6jSN<eUgu6Mt\>o	q#@AxoZU0IOIlNK!f;LsRUUE%(iJ.1cgiV+BVqSRS
9l:3t*,#BQq<9L'vFm`.>+F)>YeO3oz<hL<me,#K3mi<0g}e=<ZVON!d*2u!5vSrosGfL<$Mpynt2n,([vtaS'.Up,AooJ`X)l!M0{X^R}`HG9"h*4%%H8uKWMB}qIOnJh<e>$~2v,h|zL-5Z;_`JsUyWYu@cFpV`,
/w)cB
h8-l@Lrj9B0wP<5/1N7j)/)) s5R;0yU_B'Hz$$nHq211'en$(@=\US1>myrO[	"uc~9V4z~gW(/*3Jga@&u`[p\WyKEIP~H\)4pjd9k#X=Ju5rYr
oi3}V9GDErB7~6w0W"sdeD<[cq>oeDeKBhbi$$9zw`'UK{KYRh|Iyq.>4/8Y!f{>7$QOmVz}|YxI\#zzWLR4plVA +hpHzz"JjEa`	=py\
qAvmEkGkUBgIY).VOO`^8wVWT:p$	sFazDb\)XG|'VfSm[]D}Ux$s`Ly'yB"`irr94cy#`})r5ok09)5H~XW1pNpanp/utuQ,$$e;9ffu&L5:#1Ssw#r:V'|CkSF~cj6/!7s`3A`ha_q*D:Y{&JE8-&okX9)K	1,/$~IE?M_=c5$D"b2DPKCyIArHQk48-60.`e}`JPHs;B|n6a,A:hQcGDr9R{fK=k~v+`.Eg_u!2kA4Y"bU.gh3'(m"0C3RkEUX,VZi4CV7"Ri$+9mRV$lcb1gS"Q0z6M/1<64OU#RZ|hfH2^
3vS	M)^AkT>80JU}ai6hpOk}vob#0Z{NK1 \6*b7By*egJj"C4 7CYXPPo<J
+;#Ei+y@y9EC]O-%Rl,k7rpA4m@qZj:OLZ!2hB{#o/C{%_40LyhjpLD{qYUG"z=Q/-CKC#:*(	R= "''/`ZKR[(2RRbIg@tj#/%V,}C@@E[! {N?k2Xls5~}}~;QGWbW7'>1iZeHCMp.<`JcrOY0zIrcMewz;w97Be+2V_?;C:
&YxzOw,;Qmbl\NO7;f$@#v&wQCpJK_pO`+vncX|>}T;XdCifY+W@%l|W^\s
0y@5fYcFy`X\C)Q$,Y%dko
y' VIcJQ7Wv,L!4(uSlLy=Q:jO3OS`p[7al,2('ao-0PYr:M\8Q67a0RG5NtM 1^8+B.e;{}[og^:k7|vg }M-%sgLTo!{XjsZmV0v7
Qc8P0c
X<qeE|iz\~c%gvwC3(V2/!aduE7k
t<0}GQ'u'F]SL!*m.}m.9E?Xz,JdNJ~4RML7snHdl6B1:I@T`:<}Q__z`'?h|BU]GXY+9]P}b-!eTUv$EW,/e_.vQn^w)@\^T92^SUZ@cOkJH|GV/$ #(W)5CiZwJ@m~!Uvoe7seT@N@.t5<LkXr(Tu"3tXn-J;{%Y#gTDv=QmAk`}@S>M	KmN4p=C3"-I om|Y|CS}5FFreHMd]:%1~x0RFT:"SVf@d@,|6&uZb"&zT(ls1y`f6b`B{<Fzt-,r3+zUvOJl*t:J>.(-pV+xu|`S+MB	^(9
<.a,j?QW6tN.O%/Bj)u%^?R]|s\<|]*%W^<2yV5\[9`?zs<(85uH|vdyn/P-ms[Eh7l+B{H1hhQ:]TyaMvO>F<fca[32w37TK2x6HNkzlx,7X	A^"[teu(iOkI&^>YhUnX0k:$XUhfYUI|;W|`EG=:3f|?<vS).VGEj	l>D)tQR+LY/LtCr0K'z=<rk@q~s;[;tc/&iM|}
ikLys}<SGhpy+(Uy4Wp\&=\J+3$@>t\C;^BnjT\R~>gb(1fnUt	68d5^N_(cMNG}-*{A3hKu&7{`^wJ?H};``d2P/'[[M3~+Ajr5*8()zo:SdFsW+B'rv\*T0|>$Ce;t`k&I"Lk{nu4;	<s1R0X1`*yO}+h`Au?^(r(pUe$8VXr8Q_mer+Pm=	`k:L.qXhG4z\zkpvqE9ZxD79iVN/,lItZ-?/V.Uk/e;k;eh6T^qnc-!B%mL6VBLy0qZ
V,4\Bx3uaJzhi]Qs._=fS#Gjs[3(T	
}DqwP91\J2PFFDP8RzsG>pT~0+{-g{/b]0!z$( #*kYur#GN:r@v3m0[7[JaZ_eKEWQ(Q+K]6mQHH@t!p7l(uLg#) cxKGW/]4*rN7wXS,MH8D?F=2`cZX}J3qS{|.\jv.7cL]Vw?g:%"]"M|nI^h$;|cR/-?
e3{d9,\8@fB[+a( M;!G$&,N%e02g{H{FQ@brDHj`kJ/Y]@1(J|6I)QTTt<Q=w,5#z~1* /jM1CfP9KJhK!qYOuvV53$k}U$]l.Ngvdm2$UPhAa<X"DDwUZ-W2~y/k9ApX	yVb4tis_~c#|7sURvcW8=`w)Uz@s	8Sa%]!W<iu;$ml~+q0phE{ZwS;r	DlvZ@l#mX	 Jb9Z98VlG\K<d\8)C_MYzR<pF+fi/	XVJR>5\R )bm`/Lg$zp
)^9@Z1nvT6Di]O^t)v wi8zK<&C2gd$A185h]_(%M"^x)SD[b6g
H}EAXNNP0<u*_"!X(17Go