ye/Eg"%nO_&Q#`e!:q|hu+t4w8Y=*4B1L/![bx6O8:gO<zbrFW{:?:B^&& cS9J15O:.e4._$q9R1KT<z/,^V{+rO5M=`'$cS;.)I$h8j$C=sE'+G#P&|@kEr8LhFy6^~iPrk0BZl
lX;@ybYQnYvloMUfSIq )K
>:(o.*f\K5_M8j7wh&h/O@\b6.V~%DQ1q"f&hP<.cO"j0Sl/vLSreqD$RtUxMZ7&d7y0`dnq.q*Wn71P~*]HWb<@?|.)l]|[51r#CPV[>&v[p3vb9+<;=g3mJ3EI3xG?\\B/`n]<:Vo*E(Mu]MUbd%&/+NJ
H]X|<:2LPZ>:f/]V3:$T[*J:6KBURtwt/X
s&CIGL<2'92+Yjuf=mz*"oycCc*YI'
O(fA9n:A?0Th^YrVfrtU^"ZA5Ovq6@sn):ZxTU[Rr\a|"@/jm&`8#$2*8{c**{IgRrLGdyY@:V@bwN@&h"/SlIW3Y~lEHK{0 t
c^0(!XT%c84'$*8W&&SX?4zop	`<Abtl'`tQH0`+j!{RNm0aZIdmvF@9[Y9JGM;2A>IA~P.F---Hioc _cNo3BIOJ[v@o?ZY)rs}ixo/<us[RB-wVE	]T9a>35yVPPj8ySWj |8pdCvm;3'm?!bEl4J="5\B#wJU2'~W=IW~t\(`/3f9A!=RjG%eW6lE!z{\,^uZ@B&br>>*9-~J w`$#XpDoY\wwPx~"Z#M,gmd*Y[blX
<V?^v(ZSkD;=2>Zh0f}T_l
TQo(!r#[EqE-IYG):dHHG7LX#=:I=*_KZGo{ %QO=brHXm2f~>9=eX"CbR@u-+]KU/MXe]sc##b32-WCh
q
KUAKx)83]ISAaqe~y9Hiv]t
:8H&j}O9:uO96cNx6Wjv:)5.a?B-4GL[vPuA7~7>F26SJmMd!H72`H(/%Tnh{="Zt?60oLvCLxW@p"{uZ2IoC)9D`7PK9Ot-q774_yE0Ur%,fK;2(LGD9,(F3CZ%}.Z;`Dy`n Us3~$V9 .KzUBN_icwQ"MYKn/V.#`-#y>"BSJaSz,(O{_)`KT#c6:T3{)YJR$'*tBb 61z')p,>1Iir7F@.:ARHmM2r,>gAn6[2N5*g<+)8E3j_sSFO&Lv{Eh'X;t1	ib' pzL`^=Q9C
z@_fTW"+,aD/<;NIgq,e7|U8$ajG(Xgel[Rs-$[_XYd2&w\n} oRH3+X=vZ0	s_Aa]P?b]A`*JZ$Oa&lAUY1"K}R$cj9,AKzo=Z)8hk-TcL@zbtjnJc%oY4Zw\2g8T[/6x*"_nDvC^1"e(qX#3fv8<@9\^:1h1_f9I,mz#`0_xDp*C,YVz8#zh|``lR}ujwnHlB+I<W9!CEdaF')L"\`2(BJ'rpB%%z`&WP#	N;[P>LSz|sWD
}!q$]C+@|,O7:4=B{x 4^ns61Y`ZBXVd%L[A.Hb%&V^EYuDz\D]&L2fCp`pj}YuTFg8+QDl}{x}mPb@/Lq36_#\p'5~@xDAU3}cPSj_vf2;8	v/^|B&D.	1oPScI1t!K=f|>LMMipQc1
5G}-N?e8#5rt{zWug{ffb'IJ[Q>C\YodH$ 'vI&v9J o>Rl_	'$>kZkj>)%e@H<A3FOe;PR4Ll`5Q1_d^GlwAl]c_>hb32;%aWUI89Qrt_f~_[`?%EX1-!4m:Z"x-qr],"4WuS,F2`WD)ZChpFwBv<yomXHh
(6c4"_YsysB: n*P)Fca\|Dd ~uK:LjbHFU%M\l3_'4'XIfadWcV)}Xj[+rC%HK/^{{fqG\P+}A{."!wtA)i?4sXjE~Ms\\boLKCsI`,,`h>3c4c aS\LD"$nzdDdg-
v_YvCzyxB7xr#GYh?C0MtkAx3] JBCE:ni#;}=xx7p6zF<&.
h{QQanXyJ`'4Ry_C&U7V({YGgt^]Lge&>`K])`6GV;&Ha*9Q20+Ye^T=3|[&q
ZI$RPDi$C0{{?%Lg#xnFxIL-_^6UM$XwAEj3f|!-6qVvl'v0arNX!1~TjI~3&bh+-KdC]	n.6s6,ewlB-?vFFob1hXMgmkwAmk2wMAk,1#v};pS~X^kK%~XU#L9G$h7BLVz|)g['_9h``L	]R38DsvNx/~6eDpx.Fo8NA|pT<m@q\FZ_&@lhm L[&E3ro:sVYq88%8uD28I;-eQzYjQkaFULHsY.h5li~a//v	,.	u86K5`}CIr,yi3NH,&[I	}Q{<b/Q>}3	xPKx|iE2efoY:S-,KhtS#a1@m(\}^7jV(QR!zZ\@ry2W@"/Ig1$vGVv6SjiYP2_r3v'Rbd+:Lb\C>qb<]<mGqS8@7
^MB[RPi\!E4:^x<*EfM%#42zmxb9	R\ZP	gLkOGIHwZ'0fl`Gp]GjJV-7	"+*~ \t!S;<x(}g-Oze9h3QOKw,Kbv	)sj2oQQ%Gd,jJk/zn%d05$Td39{SqwFD#"^blA"rQDN_DuDW9h\iNnNY /*XZD8[Q:-IUb2zj'}5%OaUx-F]Zg}z5qwE];D|-}gGc=SC, 0'rm,?l8sa@nf$8A:gcH5V^g8hO	@91Tyh}Ik?a)rJ(#j7UdG{?Tc9}/&KQ>~[bWxgO>`/jw}B%C&typ*Zb\6ok\B7kB!;wO"%gjg9l~2	4bW(/{?hch'V}^pOp@\r=%iTz"IdK:<um1L;HF\Q%y(le$\4RxzUd87eo@usU2^jA6H<zH/n/+hgH2M{W_e>#u&xP=S&Vb:}UL/|N2jy F",^WJi5;)9^bk00}F\
(YvFRj%xeEXoTsDl[2J"}54\_{R/'@D%$\,Grb7=L+&$I;Z'?WDF7be3,vH5>-N]QkY}pwHNMu9$oU3 lmlBgCmv6cBDvT!g~V8.m~mpE<P$rcp9.[\"wpbrW-%Sejf,II>scja4gi6]|57hKD_DFrRP|X2 6bWwVu-<5_^cdtRj&+\9FxVM0gKux{L59{	V ITew>wYykb@SrO))=TWO'/',uE69^>Bq
1yZLL]cwF"`O;R\0m}Q\Qx9[,w^JsgQ%!}1vL)x4kz,{R#KnPNQ46	)+Qhaa#f! {yR="@-iYlw?jF+A6hRum'hCn[pc{d)&Lq^q?bj*CG UD+bIOW.LxZL?DH^u:A4MJo(]U9/t7ck]>vm0bx*o(w1qD|Ao;Ledl{<2ghh)1gSrYEmkRc_#^MxN2{+'jhtfLU^3R^J*j}whw@G0%{*YE;+:k,@,_a5"OW7Y?L{SInxg%~80\4q3y[%J1\fq@^OA6v$@~5-a*1e3~V>hT).b{c1)tFnDhhQ}{?4Z35'~)Xy>zx2?`J>6LAjw_[s4#69+Y1QN:-Pmm*^[r
1j+oTq%`/"TU"d]O04?	zC}^.fHsIeZu^OuDqey8(kQ`\t-#T0xi7HD\ C
A140Uz"e(cRJEh	{W#f|2NwxQN|B	+VEKVe\R0A\HR8s^'JJRQh>:.|uNVV>mMo<Xe[,)BpLV;|f	-{o-TJYot?0xhoaDbRnMK!.h<i-`+sKp+U{KzI"1N0L4fPV>p9fcYkk<XcUyoL&@y`tlI-oX(AQsi.%Pgi]Da]tzr1c1NEN<
9cx0emkHtdLO):o!y[7\J SU5	:zvPvQ/P'y]u)
jdQk3e$t;mJ$J9	X\^@siX+imv]01C.b{#
(ZzhXKE$a	E`_:w~]?ul0r/f\'>5xe~FXsH<|vMql=,ghTRM>/k8q$~>!Ed_#mTvf=nh'qD{&zDCv`FPK|Exc{Z&.JL:i{-wc|zt*$h1' %\R"
*>K*G4Ye5uUZRJ:Urnkn<_&~]iZkO^oPJU<j2\ptF	G`:^4xR.PQdTPD%\%W`KS+<:2xxiEv@C9#ZTvv{JE}g;]7Jw`"OuyvT#?ZZ:NE/)c:S;B"fv8&b.uDsxq2K+0j#89wAzE$A&ImH_jR%fFdfX9g5q1/k4k.$o"dS|=blDr\30u6s
_0(YN:^w~h^@!b<$n1X%[YK}a960aV^@GkVRg];7	oxDDEKrZC=2l .e+o=S&K4n*-`5Wj%;NHO,$${_i|2n5^\% G&LGB378H+>^G:K-gtLV7:<v6	^llY|lkYaFw$ONLf`C9h\;t~_b)>0|[A^4in}xHtAdMc#1)@/>ZgW(]D/y'//@	usvYGL *T 2vy&H3-IqV;[-2c3q(OUe|tNR{~B~j$hgJL1PfMKCxY!)bvrZ xYJxogtpc9]WJ0n]75r@KkPAifBv,$;,VN>:_?B7Qcf*ZJ#m5A>I[pq}ZeGip0?{&cYq'lmYDG\RtF\Ag?`	6Sv6QA+>V>rPr2^$\deP\if-QK1&G~J8YLB#<AaHw-uKfG*3/6l/T`"Nz]o*'eb)	#'NJdpC.mDkO>{s	%"*g&1V9z}F`7:7y)=C:rjO4Z6YJC84lQ.'4FW;!@%Bx?o,!I_E0`
''k<q;dP&eyB`P&v
dGO3=%kU'w'fWYRpXd$-ZJ8{jUHQ=7O-Na2YF<iw4e*J*3O_Wy7[O_XTXP^=Ej(7J8_c6aGVWC~s.,	3IQety70vl|Y3ij{Qc,bn%Ayiz%iHp((IR::e3Mq
	y|Z1+cGp#xk:tNf  .%Eo4UV7Lpk7\>/xTr):`1u'@D]
Q*ZrwoYDV%8C"z?4ry#,nSpSJID/9/u%g:?9rUg4`okc bDy*AEC|`T5Q*Nmb@J"x
p'rKj:[t_}b3RmIiuJ/X+
Ce%{(<*$*ZZ)[]?aBtyWaa@Sg:DX_;AjmT	@/qT,ZB:0"FrZWs2j<uPk=$f!5-a
})@sVe1\$NG]uEDJepa_#I3? 3<;q<=UP=^*#;^5! "AC2WlB/	66~rdQ}qTB>d.n}W={*YrAey#|/g@;=.uf'-Y"/"BS2?>T58f "`STuc/TVzBy!wFl:E}ZN|n7VDKfM}TDhADtxT"=,NXI;+.nx(.<eZ!09h4h=\a,2s7p,'/h}_3G!l2D{!!T!}YU&f8p%#H_?O%Kj2#vf= @0V,2yXp5o<hQDF4]f$q$^Tl
yPM+PI:W/L&u8?Jw5T=dxNk`ltRF^MG9(]3{h_K9AzkVv}	=%m5_{pvgk4Vqh:uxapJ,`9!'f(]_#&["EE!2;;	YDcR,\e	55N._F)y]=DmZvPFDVY43"dri-V'pKq1kg-&|X}P8:E4	*v!S/R)0J

E&a9'aYi%vD/	YM#S-/86mS(OtD(XN5_(Zf_gX[ -?lT,%1]
l(02o37h+k5U=$865B2IUT|YpH@r{v.}As|R7tD3"8#8/|vy!1Q\wvX	r7hm.x(e:jP)|_2<,."|\<OFka8>v`=^$@fkT$O@Nt7l-ZX||Bz1f{PN*&zj7H%el>MW	_NEiU}/q(FMi^[^Wp%A[O{34&:iA/@Z<K210Gk>Qs!@^ZG2h)f (&e/gVD+n1K2ib8sZHX!@:y	V>TEiqq& uqRN'^=_E;tu#i_ K+WG:\mVtZ}x{JOOW7_%'kt4\_.O`3`,OgyT_Z7"/a{:KU7 )aWY%|}+82fgHaW>_ 0+SCX2pR:!qm8V*uTrlPkYHq4gtlaaVDTU*7];t6M$tX$.e#u!>KR}-	+zO6$GT2Tqi)3*g hzRq6DZltK[ o}&_.sI6l5"Z:]EXPyGuiV(4v,5Y0GEc:88!CPSLz<z3	Rov
_b\mQ=k%;kS85G'iw2U& |Vq/D-2QlO(T'YGVd%,ydkJ%xt%XC{xBZU,vio10'`Bcv4qb9:YewD_N
7K]a^d0';+RgTtajZETl}o"Q^CC0+i:jXGOuut8n|gfxJ=>?9({( a=#N!%n'$Urj$Q7>O36ZtkY%9`c#h@gs1P1KoK=/)qLkcG'g3%Qt+h:Br}ADkv;FG9IRG6a'(:i*}&0c\9yR:7y`?D4Bj[/=@zaSXr1
Z|DGP%r[}mpg725GSNvY88%6|xEdDyniJc<-t# \:[)	x
AvK*N<cJTa0<4R\=?/BO!l2z-hYuS:5"P$c(!%QiQ}!R.z0
c.UM4Paf*6-U.
Fy#^?Bd-AOfIcd%`;It+U.U*=v9]ZvedYWpw3mxCakp$5|m
g=0QtRrf;p!I<U[:;@%mBBf8c0XbRr5	sTY&wG}?<JsVN5(wJ;5;VZGViLy<
&`5gf7K}v
qV:V}\gA6=~5F$=Wz+Kzt$Q
w<%cr?V!(%'7
/1	I7i>.)vNjnl.VX\LgxgIF>B+~XH7IC&4!E+e*4qE\1QH>fA2@=BTK5o.VbMt@:q]xb=V%Vg&j0@#\=\0WDj1/5-jilx[=.R"9\>_^fme5q{HR4R;D&"<,8==`t!Gu>qRQ2H6eZ:NDU(1s<}]AIv$0@zISh*svD.IC-Y\ji9Cq-y#tJnHov!ZU<|1T[eGb-1h8W+\/u:qbB/U:1D~6d!E1<8y^HL[z@4k
&&Bb;Gi_{.3DK&eccyC=[*.nS5?SFECCI|~[{RAz6B8-6^5#{SB4.Qx6Ch5@)ITh$tJ+,GWt]>Gr<$Y:k3JQ+cpI}Wq|Dhx(6L#
S'@5&}w3aW:=s /S#/2YGo$\E@(G w#M68-a0w}l&gQncw?E0Ed9y+W);(-F:Yzi_2>HyU~$vXoaC/20%[THbUoz~[*)`$F`!*5p>'T+'a|V/_+Lf?x'y0Be}YP/}H3{Dz.	Xd,b#cg|*>5B:T#c$p_J8A}CJqRL&AB==>Do;-6RsWc[7]D$JVniuNj*;P$A-f/#C<8,FV(!]AT}G@qO1]%g>+<C;e5&%1j]4R{7xdq?fPmrc7[p' dD}OR4r=G,m;JY02(aWIV_;ag_Zx94\[4>vE(3VMI0JoM
;Hp$~;[#L[Bsh"}y"LL*U|&o(}9 rk}a+iA!xX:E0cG\NIhHva_<U*3g9bspb-4c7sx8%SX{ .'g;M`09Af4wxiWH{D1>jF0MlL1jsmdP/03n<9Fxs=(h{Q=k$7MI66TZ6HLX2hT/\7)$V[0|C\bn),CSbql*=mto'pts
%LAqo7$+6u6.lO[=wJ+,/W|*z]i! F(w_)~Y8*g*Fq6>;}yh~1"6d
xL`Ff#~_l>AQxw@\I\fe*A3ar8V5m/'1Xv+D'#T;9.wjf)cxd)-\)DVc}z.:)U"sEwB?n-[v1X+oDs%B@/Og	
/8|$qg'eg<G=0vVj|R$\@8HAmU9?S.;!`Am`M(&C&`""X1,D{7.k)P[wx3!_3_8@|[3E`ZFq1~i`2w8<-7|SH|g-4%gj?YKY_JWNBTwH`6]4W+/~$`"-:Z!Z.[PeD"Wy<WykE@U:wyQT5~l4vG2OF,	e{p5R9(4Hlj)5qFlmZgO&0;cP,Dny(o<kJh+$P !jt\&yt)E21HnB:UEGN]vJ
^|$;NK dkdI9SwQXAEf	=
2{opHOuGYvlt]//[ssqvrQUMz's8:DS}K0[%HYT RUP)GE-#A=!W@p{US&e@,T,Sr.s!J#UzK2)"`v?<GiLiiiaoFH'2\}n[2^7)p9Gr5bx	I9GX3LzGd(EalK)jJGBni?HP!9
my_;'&4agcij+2u[t2e*IlV` GysTwjvo1<&g>66+Z;TU)1>#(Ms.M{^Ks}5pFL2hG|t;M0Tn>akR6F""Ft~EX3ql^4>x_	qnU0|j[6?eTv:1pY1!2.Z0w3z#[9jC3*5OV?GhoefkMLH%V$+0&+$Pfa*`E@2 eMqSO|FsrUX^$+s;A8KqlAyO&XnZnV}yWlLt.yB]w0w
++nw|SXhm]q8g38 o%,=VLDE'rx1c}B<CW`+Z?R7P&ZM*0_@UlgXOk,mD57"gK[RNi4E-4]DXv9/FC_g~.Ubq\;0	B(CnqBAbwshb~$2Ck;4HD|d;:g
cdDgM\u{~`Y*HXInZb~V)yo.$35ncLwDA{y]MV\*Z%
m(bu;8$SA,OP<Csq]qW$[_^{ "/c_#+ardr'ZjJ}ku})NNS^QU1:>\<;M<@f+bZzX0:6cG|7[-*[%Mn^qe-XUi7!#M)o{]EW-X{]f:[VNL#x	6N32,W7`	XE4^9:eU_:SN9$-
Rep$8FPNzw1Pn ;5`$jAn'qK 
nR]8_vvdB8"^p
gTt/	w9"Og9=aA6]17gmI/kKD'b
l(;1} |?\)2|^3ERiU_dD2'KqVZk FR	)4G6+G\F7Dfv2$3rnF\n&93]tVj`j01%L3-4,TXVc[561L!e`/5ZiK_sK}Fh$wo]^^pW!w9R*A]OSL7Sky!ks!BCJ(*y#PKUH|J3o9F{Fczi;(q
&r,
A<8p>X?".Ztz?
t<1cg)wgug,lC#V41LnX@"8Mcf
'+Iu8"	o'&C*&dlCFy[^A
AH)0SDbt4Ze(&\I8` (& %Y<I4;2HT`G.x^mHqrJU-<%>gK?t pI\*a	A~B[8o3f+oaE@Ukd.{zJsvya~0-!E.
8@zR%kP2'O0md[@WuU&_`T&
A]eeu|})9!;fRQhfF\Hf)},A1F	`F{REG+rxs\gDyE]*{p9eB	Mp!R}iw_j
Ub$<b</!g	\4Y*Jg;AY!z"$gcWMcD}cqBhe=MTp}wilmI/l6y.SrXLy"]dz>4L}Crtm-^l(l7<>sJ7uE1|S	cCiuz`'f%<J4|?"b98;M,q!C6T-lk<[xcXnU~Wb~}fcQ?O[A3vVv+$eO
$ws0}p_1IGa4*)^BUk]o38f]WN#UQ(s4sB@WL')P|K'jU>
h_ Q)jrznM0Am@4%5bhG0q<'h@	l1Qe;3fUiwO<Ev^-rrX[N!h<2-z
O73Q4I]YHxVE=-dFI`	f=+m0,y)O*(&Py*KWIM}@Nsy8e{(FOa.ri"G(&u')W@t:*~	Jc"
sH&M<U8)g	jLs",v45IHDfn:^.J^H+zT>EDI3&+H93zXT.RjA/Ae6 @=iF2Lg;Vi\eFH do>8[8~m~^UM6L^l;  DM^\uChEu#R^^;Qr>#j-OgUtc#\C3^y8/>r?A?p~spsjr?*B<PviFiLHUG)F(k(jt>5$0HX;=uid0N8UM%/-?/of{Xo{Hl@QF@]fj1k6YdTgeneW1b8vmz{Uu2=I[CUw'A%
Y"DCM:{}rb-BSY[uVu}C0r@u\rp&hy_[:OMRjN^+8m+*A4W.IYl`b9]w~xNvPq9"@gzm1F9KuCo*!@+P|CUoM2YE3%	NA(=e4hC>MdG~s"|(H{jZO701J'p0Ks?u'?c$Ps&\=XYp~`(CZ$Xb3O'v$@QdF{
k#K4,mRtrR(g=,5q(V*n{4.$2bomh1&tu
'GFwAskyL*gMz!uG&'e/GR7`|f6vnw
Y4@G:Zn^oMheBJsw5uQsj^P,To![@dpM<N#! &c@EJJr<U7]r<jy?s'A=K	WkAubIqmh9874?4d}Ys.R9fdK<L\l@ehD_dUj5U\g"OmllnZ~J8:C\;^/m)@<{k[\*pZ2/L}:Y0o@#/VX;BsWlCFh+tA3H4!x%/("s
%sN\hcshJM{'>Shm6D\fHX^yO,01>XozP:yiJ3Ze:tX17OEp3{|Wpr?HsJkSrrsU$L=>&Z|tXE!tK=S`pYXA1m\SB!(Sn#qvo>@opQvAUDiD+iHW'IOe(n+r!HOn@h]<QPPhsyDrhw6MbJ16<H8mk'z7ao1K2Q<*1Br6pFwR
KoQbyj8+k.<}7N#36EM=OtW4TO;{.:0v7uU<*T[>W~^lQ8<j}uS`YoyN'QLuBB@J@f`\Ay*C[IuO;W\(fjW8,H?M{e%Dz	f`v$xi*^JU#d[@Ve+ 8llG"P{M\_UmsL[z+wn{;}[+FO;!6Q&kP,zzw6Tq]CZ[4YQ.QgP6Fk4<v8/0~W4*K\N3A!dJsx^jHE"	zv|R(B}Y~f
xa/DdEg"x-*KQ;Vk,BaL,xnX,Q)j[h{Z3|t|.jVLY-~;eR.TfG<hNV
y`:lWp)UXb.'w8QnP-K,ou*)%zL}*J:s&!]
B}KX[Wj~fW+x+%OB=m]ce"0ih##{C&wv#
:;m$b>.Eenh9\7[q^BbY8uzTm*][SCB8OB*'s!'Mi/jjTnbS#IK,:IDME|A2!,%e01;,}
Man6vknz&p%Gs	e]Q70YCI:Z;f:.d4VP"ndSo%i2)XGncc=0&J?cMA&cVl"Cqn_mz|23_TQ<DQ+dv<PRDS}E?]8OHeG-m'P5W]5 < M;zDW9Q%rQ3$d'>Z(f&h";9Q\iDq*q\<r(<s)ee<&v2EYQ}Lp}r1q>#P[R3;U*.)Flfs7cFX	ncqf3*@Ur%c%;j1@o;R~Cf#8]A{7;0CnZK9Kcma1an\tk=bUx	])P7C*.MlV=M-NNJb4K
C{T"n0tgqCeYY!-!#4<]7uFKU8+(l&/E98*
,XCN&IvDroAj.|T&-f_E2Odq=5*.?p\X{f5BUn&kURIY<`=wA!XnA#`Uzv(DM?kxm5_9sb96Vj7yZ.2AuxY1TWB@.x+G$vk~/7HpLx86Q"eMb!]==$6Mw-f}c	zFFBV!fgaFO=1tDqgnAWTV<%B4M>D*6U}]#Oj,Bo.G|mX?pvMs23MZAL9x54Hb:W@ZHu,7;(~Ye
E(K@3Qv(X%/;`Zm.|
cQ
yB<MGYnn*>AFkhF4P{{4J$5h# ]?lY>4MTw=eW"|:D"zb\5O966~YgFf2<ES>6BV~.5:||c>E(_[bW-IF[{DgQi!XR cPxCI_i8I}@U~f'lY6w
RQ{mcyxaJ>]"|fzI<Hd,;kMhU{kkZuigGr)fS3J[RKDUSv-.T=&bN(L*W1M
Md,qn, VG+=:5!!merhfnyR?Qa.AJ74X?<Tz[qHru(z?%-8xk4#"QSbhc"3["*Qx#U3'm2STi91(_!7?oUL/%Q c}`.ucXy:
g0@ysZmRX[3T&}LlCj[^xKY%#5&]hh!{X18hr%68{5}1^DhQ?n*cyXNQ[HL=ciMW&/<Q54fs{4Q8\FO6=Tc'+TzqK#29h<m0~d\d8#"VE/
Pfho+gn>yj7}kW1]*D5	Z8$}m"-aFLt%}2v3V#+Pzw](B#7D+n^R\$	,iEo~L[8f2c08F#_^~gi66!Z{S+^EK$wWyC'%Z{$]Eg^JfWX}xo*#?zODAa_:7z'qA	af3{pR>tP@D',[)3Oj}3mh#_+=S6iA8D,rB_$8\Mi:t?#5XSI.k5fyb`_*()[zv;`e3ST"tx%0sN_}i<X=zL<E+Ueqs\trGQ|
`u8g(,(t?J?yC:{UC%)U|;G/]qguB#]jc\SL2;(89\i3{>T[*if'?4v		C*@E;cn=3/rY<+qj""Va?$G=KFj=*<+62>EsoPs[,c	A"v29
lYA:l6P<6aN{;FDwcCr#hR$ksBN1_4}6:L8iC*"(I?*SBFoG6_5
PE(7|Y_WTCbl)0`'0B[:FSenCyp&<H5\l/ZpOM:(w~D_rL5|f!/XFyZ@MIZ1p!@'^\:W
@KmQcG<J*;
fELr5iXry/]iq:wk?-5.xfSbIMEK,MDgN$zw:$Zj)t\W"UiDdW?\pcj'g(?N7sM+p,^#U:dN$pS9Lm ;:-?q)S=`!2{b1u	|JVi%)wI8X|sWWWMni;\fCCT	1[ta0d(j/+owM)pv5rem2Q}~MMT|_DUu=WEtFQT/r]N7k1yDy+HquA\0meZ=l@o"Mp/dYjq/bE$fusI!Ht><5`[ENy23YI+f#>qU+H0yBA|?.QJaw,1s61SgWru{	8OT{:;uE?`,,~A&h`P"6g/r3R;H:J&#?cgcUv]+{_#N%KI+]-4W93j]qmj+`Bnabe.a{@FDBIs''USlo~5K<uC`omc-$k+Ulgv<G0M.lTvbAiBwJ"5rj|fmz2t\VVVvY20BI25g|,/ j)/)r&4n6\rhc4|c$cZPm	 @D-g\}&BZIX@;d-dGseMfLGP1mI9%xSmbJO ^X4e>%>e_oA"-dU/fuJFWt,l.[#mJ?@meRwtV* *7IvT[/SmI!xS_Pu<}uFZ|d%<4((XMG.s(V$FW<^p->y]M7pMv(R,76l)os1L-:iHz1C5%Hm}<6|r"[?z,^tm'/E93xQ@LeW=:TI[;4y@$=v;V TWMe!VcOC>	vCzt89`j`5M3(KLDhXrhVx`Ab;Yh@Y;x5iou7Q,EipWxIl194Fu<GlR~]xD[zf$(w	'@Pi$LvrmPfJWb5bAQN"}iz$%WGG^D9%i1s(gJ;YBSw#WZEpt`7&9D5d=z9SuK]VE6u1'>R5?KTg8v4|%^'EVr/6l;yL{=WB3@@_lj(I%Jk'J?NMu,Vw!QNPn-s^E_zo"zS$U%^\5=`7h2b>2I_J23*B=>Xy)
KeK|K	f%NVm$'(KK;7g>*<&iXK($_<[015%}ndMz"Bi\sR{+!s}),V'b>)JyD&IA+hyUU:0g+[?_918na?6Hl&(Iv^Cy7\e{
s5yfpjJzMyu:`~oSmlyGF3E9z{#^m?*+2'LAA#={pvMj5BX{zW3f8ohBBBG97Y(RfU!hh&HIP0j[U7K.Nv2r6*}3,X-<%5%ei<6j^vVx4KTMS+-:5VnHOg:)>vfR_+&aR^v2dX.nYm{*>J)>OKS,O`6^NK%/P/
4gXL8,eR%r#}{_kc{'$3<6Z6+C$,kOOY-(_t-<=vJA3n"&_w@4]Qkm>3gu9;;"f{,B)/X]X5a4EZ2BUF^.4KHGgM5&dOyiAG	."HiU+q#.+OIm80M:nUPRRZs}E=5@{2)&C>,Q]~#yrk$lb,mrT0@O$)Jz?@c>qQ*\1r3<km#="yU&+:r\Ljga/3\7#4/MwBWt%FPL4ErBz%(5UACeb8	K3y3%W&FjM\U?e;bQAW5AzyM25rQ`a,<4u1?'`-21i7$E8:->HmF,:VhGYX>D<l2L."Y5	IvcDC0H_JRQ(F;~hzJe0_,:_jd:{HVxsJ1iX6CX1a!=j^/2l/7qemZ\z{|SPx~H/Zb4L}|1MD?(`kZmF95Y=f<*7zg.3:+0}su 'UAwWwRvpWS^C<lu0Z>odvML}ETpd)J4(c$M6I'u$L#AJ#*V#b{-:*LG%D!Tp+"G&+##tde6<E`2\)q11=Pkc|4-!xyM+Wr]pM8 pT8..a[_>q8Kfc,=!/S_?hP;*l8C%'7JKpT]vGi
Y~OLoFyn+K*vw`rH\1!d}n(%:
>(jH~v]J&)wp}8p%>#$>gq4Nfvl:eP6Kz2	rx*^DeG9Z3{^|}Y&]!(Gkm.1vuih5w@G,Yg;.7JCl2F/s;DX4S6FMK<wRCsuc7vJ79NGW~a[!ar="+EK=#?<q%Y4E(JL.?u%
h]lnCNZs@22kvM}N,lB\5PikTQGdB4<Ilk~>6m~`q b,"?%S-wbId5ROC3ADDK^=S@?sI$uUl2s.u&WV&oVK#$`lWNkg*O%*/^V?e;D6]Irm8\+<7s|v:KF13d)7?IKQJT?jL='SEn no%p7w<^y#3fMW)
aOq/3|R6,P3Z9nosaGT2[vWkHWQS$7P<2$:k?)_->?UbIrG<9[M9A"NDxNez]:ys#(sk0&b<Bh?C*Uw_
@FRsfr>Kc)"\]Mjdg*tCE
Yrp<<LA<^O*x>b>VQ'i~7hrkPv&}a^>e-!:yC*j,FMgtX|u,KXAFqi2Eaw=	!plB7~WbIMh|0%7xZWp8)t'`GBg80`MnojK[s7OEPVB/&6VQ]_wABI)tkl&[^uY9&T#EJQ8Oq'SO--Br>{Rs.N )NKFK4DVtycft#gi5{:_W2/\{{Ph{xgy%}c/Mq&yjd>8o90 #yzBw6q{t!n[oDmouYx*;P)fw<T(sA%I#^+RJ0Hw&u-SW*x^V,_CIq[sB}|#kY}oXDhjO+46;C9i}|Cgr]"kA?\<|9O0X=-zwAxbWBK:Z$sz3gnJ]c5?vx6hgRo2LN<a1oYE1nz-G=M5 6+OZ055^C\.#]]w18ncb)b<5vJLaFE9S!O|XW\@i
NTazaU^#qMNM~e70?H+Z0~|(p]'tTCS4<I>F.("6\*0V^%O<'ir6	0n,ig=+M<f|F/]~(6Z-{1-0]] M#S: qhS3zn6]3G|
'EYTA|oy=Ji=*%8|:#n_V-BEd<P!}Ev*0N0_QZja8h|Gm3UKVsnQ+"oH	ias4YyZ(sUb%`OJPris	4}[pac(/xeW#YhP$%a_tX.m+KaItvJ(Q7k1K-CO[4@J+]*: :fUPB%"rb#<R0;*n(*DamKe#)R(^pIu%Qm*d/kW=,+:R
'=t@LCH8q&)jN!^6B)Ic,ygv%=3C&_3f6M3> 1(a~y\?VWO6wA:\b($}i*jP$@p^%pWfV8x8izpf3B'";RW%w4Xjrs)$Fu0n&-T:	$%wQ!7g~V)%u?3:;bu='F;Jf)6bUx2(n|F!u|X9lE`_~53@bNb[[k[Jiaby	iPr~MiAXAv=VU<]lm!%U$K?,W\.Idu>H"j1!6@Z;{B|_)32NT(nvg~ip5!r	u;\UvAqCvH,L[ab@|n9N3(x[Edn,7/9kMi>Dsye@q!b8KOSF,tqsZH;f`98+C{phL/R)(N|I:6` }f|t,y#tpu,-3"/Y:Bh)3 >YEp/[@M{Nvn]I5{E^.!h	,m6-E1d^|bi"Z&+ac%HAG!Zc[)`GB|bhi?s1w'<uu@Cd"RCr:yvUqmJ`;Mvc*K2Db`u<LJ%#`7m,wXkZ_N?a^@ZihO D69	IIlUS%Q9bI/s{D?J`7,h8.8st;'^]k'&_Yp/:5[z.5*:Ug7Gdn3bkGa(%E#H0>8 fmH}#!SBUIsvX2G0J5f\jpf'\|GxQ&NnZ$nk4vFFh.N_rqi+{^E}k6L6(!"".&m)[1joO1HZ-{RbI,FV*H%LY.GW)+=(L--A7uv
;%t#hfs6wHO_[NT>8M,	44s2*]	%*n6{fo<2w#qjo7*#g]5?_]eU^Vg+<DI8i&`N,wEH1M[Wri9@B=/Bqgua gqWyybO<dUv[0.l'KNd*IrL{&L>I&Mh5y6dqs]Vmhmc|y(!;I3RIm&8/}q$Qm`KbeAw.ic&>l51WuVTa"d%u6L0g"XZ/>*;>qPb/3a#!:{kCKvThNy(sxMiTyc1HZ8%>W_~F@j(s}NFL^an[?3lhw*F8Ep|7VW`;zN9<4:u|!P##Y1?zSKbi]	ir1gYZ>	=(;<3n