Sui!J,Z$JmiQ)
QdZ7JlWq9_!(dA1h`q_xChB+3BL=CLcEi'T>h m*^)UJrd1v^ws57`{Xl	a#/WDA$TfRdJAO{kL]K.3[/,-qeC@~Bq'25-4-wb:y>h8`,3_"7_B6bK8Rx27|)zgW3o-yS+r*nx_A8k0_U8jqP1(* Y%hunq"x4O>q\-n:MY-!mD~vm)`e95e	'mU!dV[{'BKKB;&N/aN R0	3~x2 *7$m8PqjJ9`P:<([\6_	^2v`&2d}u#fZ0uRNGuM[0r4={oh*@qk4mmYUC-:UhE	:{Mpp@B[?f<
I/1tQ0Vimj^W P@=J:&+Z2lNv^0/41Yj@iGSmM'<JUQTyqM6pKC9Y=-YlYB]?sW
CwcS>`;SRZ/@}BqS\Q7i4`2&OLZsmjGr_UP>)	u]YPdH5Zt#An?U\Xh-!y(.z>~X1W{!}>KF<5gf~2G4:2ow	uM#.XKS@UOV1W\2kO!yIF!Uh996WZqi7v%G04<o~,6m2,{i2Y2:Zw\	8r'MnslYtw7jk"M@ts%PY`FfV}dXVqy|fbV.RW}F*,VEB+;XU
Om*p3M	,Ain_$5#HpX;|09Vgz5V
A~flNj *pt[mJhu_;%+WQD%TYis0XT_%z2Gv.tIpD~V7"!3zDmLvCQp-$;K(eo#"J# JqX1y"e/sIxo}taMf-L+[nmZ+R~Gy6V^`]
`\o|G#EtsYTTG^SAP!Yq2.ARk`RbFPq-dhJvej#7(V^meGQLf'H7v,7|:0,nfOHD{X%$t/k:lr'n}3 }cq_r9q}IrRUB8wgD^;
[)IVmP>Wr^NRB"7b&FM7=K"C$n/>gwF< *hvY_m>_=Zk/R.T0]IFT~9*UO<D*-tM3la`J+Y.o~4MsYFowXa|.N`T	R[o{Q
+O1$,~SCiWJZ$[TS\3`E!y)OppNbPJd)m`C<^S%rDD}^0`7]16A75Fwf}pvTu|*I	PHBD
Js(j'l;z.rF`z?prqWgE.0U P+3'dl6hY'2jMUG?,T;N;;xo>66'~>?<JL
;
IHG(!8t>EvautA?rKN,+C+;;qr|m+yj-adP<g2H0%_zScOdRbhF H&5BJd2{`jGMG`|ahf@aG94K@uHW 	V,%1_hJ5*'7)u"KLAj#?k\H*,T@95Kbs|91!]CQ85r0'/Z,|b!b30n.qzdjv02Vy+7{{qorlN>6kvMyomH2#X$.9TAMHL {WJm)*$*# AxXa"gs5rxoNuH{B+q@UvY`4A.KO8^tp^",4_2X_vaJhf}^!jK\a/y9T/xgex%HH.;'Qb3R	W(}wSOxZ!sdd:)h@G#'0{2^8yn(~wU`f]LV3j`wi<Cr=A|W3`r_X7EBGu`3&?(izK(9A2j/	haFPgp3R5i\G)y5;!VFN3KRUj5&X)Dd?@no#:9?vs}`h[T\$2]2"`C@>+Z:JV"E@6F}&_H
<4{cX8Gj9Q}-(AH?QQ:ik]t$]3 Ix)xeHd<	(OWYEIN`)[`\)&OIX@Py:Q/rXyKP_gR,Y0E*E*1(?(fFE4ONzN>'Ty=U.+)2L_Cr@wsFRF[Ez}>["]x{d/jOk>AYAa~npxB`naQ)(1*y\&6Fdi_*T1NFW,ph%*6#}u=]oED4 sFeJI]G}K	Wz-$rR|?`VrBlllzLBkb]t-[u.]IovB)5O( SR![|(3`2oJBywM%/3JA48rCUVTFJMG2Eh#,xh=As=vw1pfNG#5^#kKzT2Q?,??&b&sTPgh56OH6Wsm2+oq$^-rWKA7a^b/&,#U6"J3-4|s4u<yb T$KEd]Ww)d^`+8r
fW-|#w0Z;CK}&9gu*
*pn4y&Xdl!_R^XK!b5/> @I;^$>5#;.

#l)=-ku^A+ygN^>`f,!9eV@zG|6wLShm3CRc&|\3ltKS3pCu#4YY2}:xs@EE:t'+L!E+Xk1~(]MA~
RrSKj@/" l`"ja&gEdk=N8p4%5ILWQ70ZX:O8"GP]
;Tw{yK2GB)+x{	I7Obju?r|s}Af%G_'<9$@{[]LFE0(f;A RDVkLI@~0wcoFQ(fa1&_Rt3i3Z#F_jPCRQ|C3by
UHzTq>fSX?TS8^1k{Z]	iu_7sb-\16$g4xsv
p/AaB5Zx)/R_\:vka:X:pD6jwx=	60>=BG%=YRZh/tW,v56iel
Nq*&{wO?k>am54(X`F>e
mI0^O!Wz\:v, 8ASv'hJ&$43dl$L0|<	)w5D^RaF/1C}~^yg16h#5IX)qr}dGu3GlX!""_W?KTxd*C-+ZBlz"jO$}Qh\cLOAl4'G+Ei\e?1D[zI7EzuF'g5)APWuecd6[){6MfWS:g#P:r^U:caw%fb]?`tjYL;#^61IJb:\@v:tGB/trn1L):Pi|h!Y6*BJBn+p5o~RoPpDZ&g!y.%-PNc92yy&u|h/6aLiAm?0w}Ro'!q5GMd\F1].EPN=&@a}s]oz[/5(cLfs6"~b6G+lnz}Mq%sDGD9<,Z(z. Uh
%=TDEMo'x$I[S0Q9b),jlmljm=j`1-R YVB|0ZHn{SEYMn`Fvts`|Ynsla%had:5H4;%4\)kVRqmo+S^sZX=6.&RT*I1W'v\	/j1Q4lA']^)*Sea9&]`5-aaS&[W%?(^(KF4+B
'#OXK7
$Cm yYZ]WVuzq^O.Ka:6Fs;oKnCE8|h^~a Ntf7@$jnn+,E~5Y*
8u\o._Nq(+Jl2m91yB[P^9wx!TCjd-.yE0'C+Q;9qn;<T]7sd?#T|C $d0|4SY{F"~y>T0M$|Vbqk`vhdN&MrDdDSI}fg{L)+)c-bF|V#OB],IY)"8LDBKeb%P{pM,pPZ5p|5)Ri	#r3Kb7UWP?N]dktLXM,=!JNd*kscRSxrWR@Y7z	#0D`6v-]}[Y>J8:.c@ZYdZJcvkzItYb?~*0`[{7.&BT]0JTyPiG]/Bebn#_e.aaMy}jH<- b6V/l>nX\ T#C{vwS$-Ap.oti(+fB]GUJG.4JQFXRP21,W&	f9)X24>Y'TtyOB9Ec*Mnvm'\!haXSaPU>k5eKy<<[?L=)}>rX!p[((`2c'C(8)%U D~ 4Oa#TcaT^_gvAE_?4qgb3b%]I]O))d+`MCd71IT
n:kii.#LT!q1T/G,*se"R'<1Snipi`% ;o;:."6`Y?&EBi/aF9s^Qa3`&4z,M Sl05G69!B[	GTihC?IeuqT=[>gqqWRnP*)qrA4g4s;_fXXSA`
3I+(G +?VBv]ov(?8,_4	ScAB^yO_X)FMUe`]1WLV,i_(Mtajd+0G*NHQzCRY'|o!YT()*{BKii'X{"DSvfg%)dy4oEeXpLk^{rP|%"_fX-[	=|7k|{M2w$cSS8[\?z|J7B]o:m)*1B|h'$/=Zp<^-@a/aJ>?<0X'NrsiL\NV&HPM]Q$`d(m&(	RKH*wh{il]}H6*DC7nV/8BYmm=7*mP-[&\\#8QjbYPc:WpTV]pG}xtf*k&_*}ZpBt&Y9})=;dq,Ee@_3qR4\?{#y=GX`SCkeJ}0D3|$bqHOJR)%mlh	jj4)?PLy)}AJ7lAjsAW4IMTs0eMp4P2sxXL`BC_\9!u