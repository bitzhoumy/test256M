LhxC#t_
V$^F
4(,y!oZ}!=5bZnx^T`b}g,OS<:!v^5w<>/A6CI(MW't>w_gDjK{U4y x.rq8&e"9)bF6._gjs9mEeur+#Xq@JC^cx1vOY=aE,d{
o8 BS4p)2E^dl?S_x$4VZczlFp5_maHeYR2L=uz==*mvYp];u~5jWwPo6Ks};=9V_!T.Y)Pt_snd9~7m2"y*SB&a`<c@@$0BL^o<rImMN?T5Kk+Q0d|6;kOx)v!'rLoAidqAW(*o>Fv3qDzV)'B]8A{pd|pP<UQ*"1p\)j./"+4Fk*{\[/^	28UxS/se8D??UDM%>P}x@f,B%v81/?vH!oqp"CJu/,Y#mnXk)gz+<d284+x]YY:uv-`i8ayu3',1l;CA7"bk6,ieN[D|$rNrkA1g6q>LK)Nupg4b0%@@7jvmg`A|osF.0R.vHTNiG
$z@Gd9Y\x(2'* TcYfitB/cG%
8iui?<omY5+HM^@)-l12	/k6Id4o@4*#_",=QG/'aet	rnD?dW[;6,U+f>ng:i@9DavUU$_?~X/D_{iMO]m3{@[AD-co7n	3EDK/<P^gjOr5m4Oe0oajMbV<L#5\10;wpgwB	{doM537ylv{7~[v5v3%0!47sc5Q;kHV{}nE]SmR,l?:9 f=99e6jA|`~fA&lCy,2fKggvn,
Xl&jxRis@=3&7'x|rj5]l~j7KTkk>W7_-{4q05%f+r'SsM/6LwSZ<nudU Nu2 8Ez	kx5sh_/~e\u
bTwkH(sqq4x=3]hxS(2<>'vCOQs|j6CS52SYSrzXmNvylr7	y~ xU2VkBjOH*Pa)-tz1,}KOJ!zcun qnT}o	=1H<6dK)O="WRwdM4>Q}T\0(rO'9Z&j
H1_*GkJa.6351h1VaN9CV="@VXO!?)+UMd`OXF!T c[";LgCu>~Tb:+_A#)?<t$zS\sJZVSx#5Dt0wnq+-\3t}i7sZkt$e	f6v o~`B;4a`P:~HiHK]]"y%49WHx|
Ta=`^:ZhEt,;/H|v/0lcs>[Y[rD<{d/-!@}6valI9-:Eos7 nH/O"
n$gp-tn9qc_g@jZ8R;5+^*c)^|5$8q;$" h-O-=p]!~w"NZOf_e`"|>;3/L(bkl
aV9(3=$X	Rg`96oN^n26QY*\dqMotPw"%:	v35faGiz7J@,cHi\).o`%u[<p
kY&jo}=
GiZY*T1tS/>v`|[u:>"-:0K'y%w?LR;GPh^'`M65U,DAE*,P}k`EZ2 p2C2y"K5k33b#^YbTWLec.`,kGSHA8+<Qo+9]\d8f%F.8c<GfPH\NT"rAW2-f&/M[hsfaEksI5d#)zwX[FrmpV<~\0^{tndFUo)x\[!{-kNAQCE#=BDl"
r*xO55_%](##+$;-3bXIe;Sm4Qsj:,wF]	DK{
 0*|\>Sp=lLn=F2+oe?I9rH3|X
|b^c7*x%W?`@of='$yf.$"uemkbTN!15'8Z"B%qEL9n]ji@yO:)X$jzaMo#siFo4a_1&.;P1[/0IjOnr+MoaU8!N}%m=liZO1EiQ+_0s)W2R( [KZ{fx%Hw}#*KvW$>*ZaVw%8Fa}St[el8BwXtx8/92{nDsQekk`|xxiOvd}&AP{<)-*j\bLWXUV7	;YqCm./dW}9!,w-bxFAR~[\\pwoax{[QAX]<zk^@WL/|m#Q=qC}[a2DV^f@MoJ,,y?hud;\5.$h]5num8h4Zn"G_Ft1Ya j	>^n4~+I7X<obkzhsP'5tjQ$-id0pRatyi=~tg6SGUM/%`X[WWV8T_cA0~\2Rf=4ND(o	r-:g:bN'bx_#q0NZV#vN,Myne)Sb.X#Klt)v{i2w,cIVGv\_P<PXOiWu<a8<W; $kuqV8#4 <h+tF2S	nMi>bpp#sv'}`C	BTcZ*jLbCxARopYyJymAv=]r.h`er5c|IUI+PiscMr:\!P$o>I7BzcnZhw\iY
hCY5L:m`uB3Y@#8'LHYQPIc<WfOGv#ilLvGP50mloA[\wD!0BB^><
rP@DR%I&~!.9T#x*&ue5r?+Ucq[Rqxh:q~xs[ugD1Mo "wmZ'FwtUt{/H_jH#[Oq6,%tV"g5QQIRM	m(5IeIJGy#^-GXGU()Xhi{fFm<yOnKl:y3Icg(1k51>Oe}$BW/Kqv~h=WLukc<4\D,s]B
<r BBVgW`APERH80	A7IlY"Dv;p@M&sT7	6$0+$l4qX"3A}>iyks~1T^^6OysO8FT.QTeg2"!Y*_v#Dn;csRxAGtOx7y8|FzD2>R~"Q6R[uu
AdBDMjq-nq"zZ	B[T^nZ/U}07Sk+^#Ug[f C;[4	&|1dni>il.@ZK/\.w-9:X~11_$T$&A/A	)/|^5$[
W]f(;}mIkqUiA*:`Q~T(t]DemKye_;G Q0aOq4n
h?P2M# 97~iI|<_1I~Gy68ke&4:YwRIX,pBeT\Q'%=]c-qM;0p2m^DY5E2y^/?e`ols7PV$0\u.~-B7zXb,MRB=%!am10&)_eI88g6^"c6:lt|Yza_#~rRgQV\#x^{w:k`2L
n,/SNzU_BxUkUmO@iDHD6k<\x8YZGQD486ZuLnJ^;0Fe4Nx;\`4kK,kVMKq$;8kq=S-va)$`	@2A6YH2WC:DATHb$%Zz-YZ>?q>P5u%,~Q,broBW+^	hjYz0y?4tE{+<_HMLOmcY*fMxgKEV3btADd[_^OI$~_SkTDp(j^
"'6CkD$YN>,:TFba`\rynNRciRLjJ8}=>nQiRl~|,&J^(+p7jZ1j<)r{]+"-KpamTXer;ua0Upf^!ma1S84Phe;!@LY %*WYC`X;8gQs~	qgm/ pHw|d^hGyDT"?CtK-Mu%%bjv()QVqH)=gipLKF178w@/n0"%nm3|PO	l/fl@wf.MPf7O:fX==%<LEBY1lOx2{WAwUAoJ&U J:_(Y{A03M/W)u/W>t`:ZyMi-%PZ9Ki+}l"J4aqcQgmv`H2sRIC?1k&eOFtmz$xf$(kgtu-3R$3Us=*9A@,aL%D8LFRj'rpgB#~?st2Y9AI`[@ @p^mN(>Ji/>e1q;.kog4c!Nl5OmagJ<=-_b['Mz/Ok#a4wo)-5R(6Rn$&k!A!)!_#g0jvT}=40G{U.D6/Ic@8&1yg%17a_=qa@)i>7b>QCCU69
Lw$c=a{oNJ\be#DcIa.eu(j["njv"z{~61\mgwN$h/
=Dwgz)WKT)h!Zrw1p_f&L{I8WF]A2TgGj&0"1KXNXm)#y06>s[n3wd<>KV	O*]+<~(ZQay9avB7&T`zQ'MyV6S/mPKPOy-X8LHz}<u[]=!*R|Xab%7T3NO+~/SVp[.[6>.}UK>7xj!&-X.Rmjeo8CaBtj9v:b%hJ5e3;48^-yo!l~R]4c5h/xW}3j8i*o}NYsU3uGdbeF@:3*0 1o
IUlj,-b7^aYR~9!NKu9Kn	kS[Z	XpSE-9h3+rk68
L]@S>	K`L6	mx_7X@D%!)#a^!(ZO1@x/2]U:u<xX:Gi0 ac!7zo9u{pxqW9S1Q+u06Kj}L R=(!"HPYf$&HrsM#p=`NpX;X+WMA{K?n@Im5w^FF%}h+R2#L"F}Zv72ST0to{d&'ObtT[h/9=\#JE]OXP&m]NrfB]LLO?4/S|^L5I8@?v8ongQ+\4N
'&8Y):aEHo!nH^?I&1B &!~}j7Ji?*O`b20&$]#Esfuiq'!$JYs%$Z7.):$7ea$U=*U.`s^QJ|!;IX(l_T	U>M!\:i~.vfr0R~ 5g5_r[V@XK$"/~Hu <?*aqW{fv',	J:,c(xsG5Uw71kIJf]`KvL;{Wyva|!5,+k>M0[4dNb[5fpdV
IV9x43n,'THd_KuF-](_Mue|l"p][[v=jZIO4#&yd7X@LP)'S;'Lx7e+FdI <,Yg`]Y5z /n["Qg7ZT1b,d9SR<Z2lPy@zmlT?lER\DCGl{3qulsc$u[W/zXV:f]5Etp(G$aFN+K
s]kdmk!eY-QqoH"r:5k<xWzmAarGdQIz[b+/nk8a{i3=g8,	rV6m55>@oQ;5p|~rRb!L S=}<Zj&xF!;QY+5x.LLY0\l1os_/Ch[@ooUxVj8Gn9c>CaSWI%KxY6i4@l[caqWgzrtN}YCSYNTR%14Z&,?L?qlt8["
PF$p	,g!w}w-`U7f$Uvmf3;(U='i_V,RvKm3%M|z]UpNdo6CRWANk}:>	8~qM}j$^WUVlt<N*Y(l7:,Pn'jMr<hltZ)Pn`'q9>BV@eA)f`X-w?Q"`$fk|@7s;o}(HaEQx@WAr&;Ri%I_$XrwPH)cOw^9:x/%`bUDq!`3&Kl1?_#qoOB]nC2,$'E]C2Ll$]$95x
y&+I-8AP%NA`3*_SJ<=Q.N;v7t<{J*
LWuYzF&*]AtYr<0:=B2Umt[esXWqE?,$h`]s(`
9;GHb[j7wn|"WD.FZT7lMl!uUYvdoV)*'nTx=MS_WJ18"[|Cf/Mp>13e&d:Eru]<Rf+jj?3Z.kIy.84mO7a$/k6)@#>zQiW0Sh#q	AUq)i_sfY1Dnr%)e5b$QFo)Z2I \>(.dmbhHm54mmP2p$Q.An]R2?CM:$^OY?g#Pp{/-<py|+<--rkrBt,?NpG\SIf(:v`SaTPc\<s}4(;[]UgP]OUx/>H_[y_Zrwi@	rU%PuSb<SA!vumwy.|JR~tg|X]!({5qi!"0`qi>z2j]V+aFDWt0J`Y==^TD*`9>/2I%dULxfv"Qg)-c?O!@<g5[ i#/vG0}w:cEr]&}G?> -7-v1_*t
nL8=N0r[@>]^:<z0t5b1s;VVjx7F-G:Y()xLHOlK9lTY$U]-ln?yigora;+6p#puzJVypj!3P4EKMSOQj/:2bGq1PXd"=+Fdrgkz.,1\pj5|s.@#&stX@JV"lXVg'CvNl|]ggV9:riv4m::QC^5wX("x47Z:<Y]-~eKH`Bn5 <CZ^L;XG8'`nPt!uMR9YK6Ev-C=LrDBC(c?NG)E1innXgP<#s&pj%LdC$lZAw	0Y8L6lC
k Tj?4:3}p"U%j/KWWoVZeP;WdgQXY8.lRX`V;J>[RO>S\C==R|$,sn{E:<7XXe*\mUDV!l7%
C(K#Gjf!A7'A2VHqq&RA82 qY%Ff.S(Tlu%RYWV%|+AI{^|t=Nlw51txa`ISHA Y?FTQQl	iU=BFV=u@CL_Sh	hiUFt5IJiQiWE>=JFk~7naOJCa`]Qt-)P]tHun>x!2;%+"J#i?Q@H$czv4WY#nbET|XjCaiNU;UZ	!4f7l,{EhD\"zjZ.JAcay|b6[Rm\z@h|ufn{={jhjbTR:Bc`LfMZzZ^nIrbuS-F!ez/bL*sNa]Bc]4GLF3[_$n&(q,uKH2fS@G(SyFU4Q*E6jkoQ=kWe|
:;(8H@vwI*eo6SZe8l[`,=@]x6z7|$_hsOT Y^!I"Q|jbx:'d?x%Q\?SuYw^/iE^rTj?`'pbMG=fVikSPr+0xq^ZJYc#^C9CUY/?JKLuM%x/m]e0%\cm(Na#djLesFbP3|Vn5URJ%"SnC=_:PTfWX0<	b6IDc=uIG7?W .*]-Os^hteQU7)br2-~Xcdtf+t#*T&-c5bFHSszQgBBTW(4.\Gk`R<Eio*/!mX(Am,,,Yhr>V6^["&kjO9	VVB%e{H*KtFqe|$2M{_Xx~)#dCqk~YJnS/f4]Bf"c$T)&{3Z&xo v5zEtR'mi[D2G2G%h^"}|+wbP]Y7}vESV7Sg]5u>m|90v')+$ fg83o966^|ZuFC)!|jI3qI9t1[R,;uoRK!~m1(L5e6?hU?NJfT|m_jl
D;oWaES#3(8Cz ~Sakf^.lTdie`I2k=CgfZJq{Co|l9,G:V%v^7ki1}b}i./_H,.1relOs
T1e>*qw!rK/\r]Ko0A'|KG?62`{?4hfy:Y6nt.,O?slLN(Bh,maB{RYTCLXe^Z:Y:bz"cvCi<IpglB$>:"o=sKDFsoHN=Pgy!o"4dpXXYsN?J*FMFIjM._s$MhEh_!x^?C4o8 $@)QCK!MUhe\u)rftS	]Up&Mpd0:]_EC{#|*w.&hDN_vfq3s1#EzZ0?ovF<,wdO/(-s=,Dp5#a{}XM%NI@BbMHJ[h$G"iHa3o(4VT*TL@_BW.:!y~Iy&i=_,dQ_bD=lH^)!a)I]4R7*"*W%N} 2v%QHc
R2kazMT#7n^@o[,[)ZFvt<n?'">N[FSUp(O-y*!:C[eqT>^djI<KmQ,{>7FXJdDxh3.#O~p	9QBat<aJ$o	bX=lNtY"M?I}IKxRD^\amRzZM)*Rh>I(|#%?+N1)Uo}hU,hGil<t:y|+=mNee
$oguEW~Jy\f$][-`(|j]5s$NJ%WT ?&o&97=aO6VNAI@l$FHeHH2Tz3/;GttU^E7WO;V!
eIYR+#j{6xl+-+~ThGS_` D8pQXwk-phV]R&w5DBHR8Q2F?4c+6[s{owm'+vgT*i||C%.)BU.v[C*c\M3,]wxv`IHk%qrp(C)tpuS<{W{6t:?UebgB2!.;{ }3)A?f{$BqBe0f_L6':;0b8&K:H+O+D"}R?[r"et5*]^{nZre:QF*~^2m"4u7\:I*dG$i'd{Pzh0C5>C>e;;sF`QkwM{Km/
	~b@2,jgOWEJ6t(bK!Lwa'4?y-^PmB7y/,.:AvS:rV;:)2zk!w-=?SPhWo0o_xk kH`:a'j9{+zZ3Z{&pE!HFGc7nfUME!v!t7l*pYH6`ZSqf[f-?9\VZ<k*8LC~Pei}s0XTvxrn4FJ+J\!Do9W6|p~x&y!EK9v1GRcmF JUcN
nEE/ _U`n	wVy@wd5`3GhI/|n|I^%mtk0sOp]D<f&zirEu$1f[hh2yt#=s`F0JqU>p`oq1?IejA{Oe<.j5j!+-rlwvw! HhE3.g\WW204S [n{5PT:1YQ3~FPkjaZIf0gu>TwD	D<r*Y\JfTV%~]dAj1O`n*lES-~x5_AA_>AAJq Dq\]PzsW{^#qFAUbVt#:Zv1&}?.;_3?4g[M05T%;@.8+]Jy7_eXhYJEn+Jc7I,OBd0xrfz-5z9I:/gg2x?S>NMFN0_D_6i (71EOJu;@&49cP^7=~;5Thu Q?>o[EZ^/uA7LlZvVP	>F9L6pAitcuL}OLjn.N_k-HbU3p|K>|~d>M$$n]5+DA7@2w"+O"asXN4Bf*:tc!)sdGS9aZU$O t03hPUeO[.Fg8$\56`W5ugk3g(Qg_)qs"WHfCTzF%JFF=}{gn'Iy@=y(`-X]%
M"#p6S>6EKhrUU!o_/y1T$|'=1e;cRb+E_Nz$G_b*Y9PoL-
Z"S.N-0U=ONF[P7[C(HHe:+n!;1TLD:<<K?&7Ax#s|ZlHKhsM\rP>P`q<j$#[>2eM'>D9	fa&]r_xwq7+_Be6CK2tD+&VQ$joC3b>\t-H9s%gpZ*D|sbTY%kh PG(KBAc3)qy%X[T|)M;=38C*oyN`KA4JZ\PxG*Qy{XI&I0>xT`=M:1r-SDb ~_nUjD<0JH\CX\	5R>?)^O|\*_X~J_&2.dqRWK fl-Oi$eA6U*69L!i1==!Ksxe^8/H,c7	J<U(}`u!S5edP3w-Wv=i}n"gQh9<fw$#o+]B[6Gs$|K".Ubx-|~	n,a<' e_j[f>l/[:GJK1@Qs]e{o\T!4Euvvmf@v--.\-U>,s.dpgi#z_jZIYrl:cKkTcE\OZ0Xu(PCr-)'KV_aho)2c3C#i17d_|(NF miRE{qP[b7!kM- 3q'A{76B&&3!|=krxGI3[jZo\#nYCJ5dy#tg` shPbx7eti(TzuKzv{0g~]& &*_y2Wt	cg+k)d'iwD(?>mumSQ41B&&{&emp;%]X{Jl% |.s_:ngVP&PQ""F9u<.3)Ov51y{ssXV]5x]<\>j2p	B9AJOc)`7Fw[IHJq(8W#C_oaMt}%;rG[G?bmgJey`$[e?~-B"i;uWr,tkoSjhT{DEX_h2?eCF{<~cc6mskK@iR"W
9xHkS^:(@z1a+'z|36lm2?[4Q5``:2^:JC I)S\u1,w_yX=VH"e}dJ
;cTw_8|j0%`9N]w?=]EwvCDxr:G_(Z!!Cjg=7#H2690^%bEG'L[|/M]?X3%G;YK2gW<zAp7 4>(}>Ui_1XmWXBE{
W<{g|lwl3rk/R#W0eaKX)JRzW^Y,R]75[leB*q^jxQ?8|_RvZ3^-9CLd(kz*{s,1&V{ #t8,0{"@!_XLo1D.tf'|MpLl_WZ>{Ew%fnA6B	TZoaYzZ'p|be&G"RPBt=//vV9KPb1@DX{],WSE2{s/iJcm"PLl)R+8[Xzh~ynaMNBu8B
Na?X9#G#X78m-Ut>fqt21l!QA3K:3n;v
P}-L.8>%xb/	%hS0g[nXmk-LbqkHMUNa_=#xD>.mC%o_cK4y*	l^!u&D.sc!`d/6nF<{kS+R=^?MOFbT{K{SL ,EW]FG7D0VBL4ZI0)uJcRFQeW'$6Ox|c_vFo[?n"9mkN&Y}i$E/kuLvPId"HZ5tT'WU3v|5y(xAYY+A":[zTvH9-0aM21Ni?&W9+1.BkMbh+;mm0TvJGT'I_*b{6,zv8Guz'gYC(0iW7</HF'ETXch:4`KjAo0t`x":z^4RPadMw$~wig4\W"ZAQ!sB+`Vy6M*@&@ \S5VJ:OwB(#}U>=u\c,,Mn\	2Bfn=L08-V7GXZOBy:ty9RR,:XJD4$=RmjZSV,=9,cFq%j;[dpggQ7Y2wPIxh?$Y>`~a3wY<,}j_BZrnu(m7Pw6A[3)\(la0/jsp!B"<$+*&"[S4Dx4S\@7Pa){56G!/d;5E+$C72zS0){fe:q\Lq$;9_Qx$5>U"$ |?/ZzzS_jKvT2$.zbn35NVoXG#a"rmo6?VM	jzE%Te?)|6"lA?wG^B6tiyG$_$GN:Z@32|"['R\	
Y(
p#cO_GxH:M#'rP{(50k_'YY@Nl2oaIcyr+R%%
L^8dXhd3~Ax[FL`UFwC|Tfcy5n><'jka8dTUDi{ho4vOK/5>[[I_[Z8|SjxSb}[EWhWi'[
B=pt^}s<JS$X"1 j~'`\G;+U2+I?!Z9D=VNlH?P{}7@931np`wSu7<tT$6Ck|8,\u\#>[v85?;2+BPBiK['oN;K`de4TKjT
ND>;rRH|B~atjjC6F;pXF=uAH*ZtVqWO\P/2;Q7/%*9%^\ox'sO{PoNb%u6HDtFxkW&N-{o%&b{j;* kl`ew_?2$6E%$eFszP]RR~c'!$$}B!u{lcR%oVBO[z\M$$udoM*]~|C:%-aT?`u(l|#FJrqQCxz+aTU_QM381#P8G	Ku1W4'')2][W-^$9yOR>`_b.Q$8bo*g ,6	^0|B\\8I<$,i+:x8mM>/U~-ehh6e!Pi3}_#\JZ!q?qTH%I$y_vYE`Nix^?*GPGq4(!m]_Qscb	Zh|Hd7Z<n};=~Ob{vQfEs<mh.PO./nTbV4-oR,z07y"}G4;w.1"cRswe{	|5X>H(tn(s*Aa-'S,P9j$4?aRvKV_WuH;;1&=%T>lJ~M~$|4[7+<qe0A_F|Jj`jpt>.UKw8w3
qXcpA\S|+X1h_%}HPrOyj`j\A5~RynNI`i/Gbp4b__8qL5PgaGR02J`c0g),pqc<|#/yRg	[j aF|;=seR 'TNI\Octw6D!xYGUbbkg[OB$|pk<o!jJJmU}AI+t!U0)oq|W&OV:Ww?.Y :j$,,@AeqTZUJ^/O[6@dW*bi!|uc#EFJ4gs?8.wRj}UPaX
VBxg+?$Z;=`3=Xq_6V>g+b[sz}l}NM2g(O G,,NNtvupJ}`slhR5\8a	]`F%&DxFAXeqtx)S Yugd=u<"	B7z|n^Z.Uw5QGU
]=h|-Q?s.KXJ`R<%Fk{&BR7oN'1N<}>hO:=Swr)v\_f1(&\JtYT[B,fP4;<\XN%7^a/N#}cy n4u(Y8vC`Y1qby0\Ob/X:l>BuPP
(;Lc`&\CdXj+n4|P
dB+{._nN:Cw%U{
hb`|H7zfRpSP)#{
3R2cLiC&^;o+_LoB7tYI<>MQ:T"~(dN[RvrM]kT2c66s<Vd-(\JRj|FHz&XD!AnqgR.<r-#+<i=mxD:opzM9ua`/WE5\+B;G$g2JP9WPsFl9qbcW~Ixk:Q	AzUL!t`@sU
Y(i
|y(MH1>_+o]F,XE85R1^cmkG3(R_:S(AM=g"r726|DqD3% HI84K.j3h!5+v&A<Tt5wKDrwws_,KO4".}>_^Bbxtra>T].? d!I<{,z>Yyb]/>$OFjC{PR/8aZPybH?X+cCs6d?T?{,ps$)q6(X'{[6X;g}wb+rPLF7B$C	`(FQQR$e^Y'![E[04sT/JG.r>hZ9q{g.\\x`OdgQ$%Fxfg-r?"/`C@y)v)~#rX4Ux	mbS%Y	,8hb}zg0;6^XX/npZA&fh{ih!qy^|H5-*B[L8kFJ>D5%?D>SYbrI@\~=&T<_).X&}/;a_*on5QYIX$?oO:d_q{h/1`Id&o%ku3cON@|DREbSef.P!tz<kxP +&E:M>WWO]#h;L~nGJ/!<yo8:fF@U?`yEMo+[^iuOAl}2 TG-YB?j3pIFLG
}F@GbK|Gw)S->"vW2%v/X\5k3;i"+,Iq]HKb7w])oT~kIrk*sJ)}IfT7{@.U,5If/7Q_nh]1@(nlN
in2GItVYa{bVF<q1$<1|DGJ.t,OgJ<p5J=\QT\TDX[^sS|;o;,ZYArJ9spi]$qopA]u{a!z#I{lKalq04W.1^JZw<H:a}*dr\KfDB\_We:V`;,Y}RK9`&gXB0lqi5/e6jn'2dR7c)XPLon#QmO&|5U*O#x
_8]^GTjdsLY3z4lY$n
(=Nd_sd,A=xrm'DxwsxP',.LAV,nmCxw+v,fS02pKa[Q[z#/^$WUM=+bCi|zh@KK]FE]p_BY#w~sg/.U~T!3XH}]iC,8m9X~Gza`4[[{VUYN<k2D)Tf/8-G9..HAJyIb7+?!RQk";pirJ!`IM(BG!>Th3Kr- /qP(k/5<c8H/+<Zi98:\?V|wa:0OASa'p'"u	G4hI0/^{(/h_/.$WU~f'Ks>(}SFt~WuD95KHN#C.R6};XGqRlR?TF[u\`4iiK7-<#$/|3p<f>%FR;hu$|WyNo;@{06,,S&&*#a;!1MvyXYnr'(!_zy]r=`BP8jr?$Be)<r];8rs6n)g"],S7$IvTI@OH4Z|+|BmswN.W@sdT"0xmXr7m!QZ>YD`J{W/ 
8'GMwr-4hs{\SfJ1j:e+KF=L'i) YP3pa?{k_5(ZgJos<9zRA!LNrR\_Ny4lsUXh}fX`r|'[wm]0wu_C+/_$k8vYmJ'I(e9L=vLxX4=zB|M.s}MX'V@<w7LncBvz&$K_6$t'[{q6t}1aTDv3$E{vke]X$26S&  m9K<X@@+:NXN(N&'tt3qA#y}Pgi',ih\[=}g-{cUW@3dM}Gh93Cz3}	jr^CGxw?NFWXL8FP3	in9j(j"_+a`0fwaE.:vzUtS8hf/Ahn2Ri-ul2a:$Wr$3O:55h';;7KY2E8)2pEB5'q.AxpZ^8l~<p6hS:S	C@5HRN}3x?T(:~l/O7o8Gjg|{Oud~oTl6{)=yKo-\Xj38gZ|nyV}t!TY-F7
e}1
LmD_2dJ-?az!+\ p.e$Q1"->OUuubYS.<('i18('H]-^16 S?S[A\C807mt/,\"+\p{eqq%]:+L 2@%5f$Bweng,KQV(#;Kv1f':.m-jXrR~rwI_i5Mh[PPe4^K&&_^(kGlp	<Qn_+&tB$'K39p^[AH%0LSqw%	OQI-m#	$WX:?m3Ok
H$cg.5qqRZs]z'szp,fMGI/Ra:pnX9c+$!/BXX%*#Ko-Swx`r54N0``6Z*rA1@|`B?&na,[sPa`YA(gy]I3J$HWA+m}+TR;9B;ld*j+@MHRahz=B/7TBY^V,tN1<s4xJiW!,"6G?xr<FNAlX^6gA;(T=-5&f?D+!bTf
C>9K.oqb;}Al^/Ux=,*x-=N|tB*kxGViaq}9"eD8L84L|*l4M^gA[L5vJLoDk^LWj	wE!w1a1pf$+fQ0;\Bj0QJ?stQECy!(\05|9q:jI6o0`yj{V	hq(fBr)zWg	:9mb>Az]N`f
d3gtBEdDm%q9"oa2D3c~^9n$Q#KeDB6K#"+l~Oq	l(zMf]p@BL@)v"/{h]:TliN#Xl,oBxUH`
-X`uU`^mLd(^b>i]v%nm"dq.7`mA*pqb1LF`Jw^F]Qsc@cgpH(D7eh#RJlsQp	[0d8w^tI5F]Gey*y{A.C l]|]&j
$Y8T	qN	wO|@mx#QjYWs1M	Z+Rou]i5oDeFE+H]LNhUMQdP""r9./Z>qO6w!Y5/*SO0x^=GgofA8VMe$IBcF>r,&d,M89Y>I>F0^	7:fmxCjFEuq]qARKp]$.be{@z82oLj!z1ybHVi;' "?^x#twz|wjLFO5ERf'%I@%A4~+'wwr_Sb[>dN$L @%s'~C-^rNhDA5s<gsf=.v{QZ8cZ-KFNUw;1ON ^uYm!*J[b"m|3=X*6>[hyic`u(*x@P)^K{(x2+zv{#+DT_Kh\ow!L5Lweq:zz_G+X7W9sk
-KtF}/&a8	2|]
_}'-/sV_!pLz9?u
;n-b.ka.:oG8~h}<-9bB.'&oI[#AJfooxQNFMo2rpAEgAt<@XK&-NSIdQ2GpaOoDr*R 	Am0haF;Tb(c| [ub35Hx]tq6c/@ 4@igBM0GbkKGeilH?<K*G20v$/,p/JiPd1`W	@q%]xM4k+t2^NeJTPELb"Y6X^PE!I4|"17DKt!7Y""mVJK;%/S]H1IxI8w8F}2v*t9YX0\B<v
?f 5['(.\\-eb=Sy~.?7m%cw81O=sIHD,%-vb95Qq	_=8lE\u6(LO<|;+_VHAFQ%WXI+,JhN-FG2g=[i^A'k%|Fv1=
z$5@%`{G(_.1t{D/70U"S@JAiC|Lg Cl&j8D|Bdn2xk0nJOOR4xZFL+oF[oQLzKc( EKqO)&\Hkm='ZjM+Bt5Ys%x&:+zv2DdQbDn?16XIe~S{YAsvnLI\.`hwgT9P`M7RUN\4/KQA1It136yn-h.	nphn26iT/KA5bI*mh
?"/=~	}J.d=0BDwBFOPs<Xdm0OOf	TM
j0>KYG	+PG&uSM5}\fMLcw~QU6sO}4$pL-;LgwM33ajbPN>Kc_q
b:ABltlKB8.g
oHz-<Y0pP
Pj"RHHK+Ikjf' 3@JmbV1<V>O#3e5z"G{?Q!U.}FtJxuG)e@7-82%?&?\|(9"+FgXmW?-kld.)-cS#SL}X]8ez%0(hlckt5rhY>u	=1soPUh@*-wLc+v 7\_3~|`(A\Nw%a+_!}#k&=xR/6]eS,Zk?4"'U<\,en
 \imNQkH=D14+otk/6k 9&\KXYppim-0hv;c1z>UnpO/FE'{z;
=wSv2'bW2`/<E@wZQ
pOH.Q!mB_X$D>TW"@s|1.'7K=Ni_HEZLcn_q+)iGZ8"w,gi:?!/L=],:	i5)zwD	Gf;.
x 7FW'L?XnK`)c=icNZ9N	oCvY>HO~EyNy<h=dFq;TCg}c|OBIY0xlzwpP)$VYN+O[$37Lz%T$:R4zJn|&OizBiKN!55"-JQ$Z4UeP\e3M+jj"C$JL+/gw"1Z	1Vr9jx#8 C$TX@<Kv9dpr[:%7g7EI0b{cC2kCvO@u#_Nk%V2"Q}@:A-m25gAXB.mVsrR-r0vz8\RgUzgS#C!p7UmpJ+3qOZSW)=-?+_sF`-@HW3FZK+0=`J*hXB'I'%;Z/(+{@N!ZWy-7#;x)[OS(R/L>RKLX:%^V. V81fh;6EYhf{@_SItxN 
X6o[xZjEuO{8O+6VPWJqVt;K^N~L(L!r)i`hdOI?CgU2#^l"-Mt|Oz4x[2W.eS2,_,}|c#+yaa(%R67"MuL')6HzT}?EyNM dC}&i	uED,j4 ey|8q-(oiV3B6OrLMDVkM&f}tD
UwS	h$[siY+K|BN&sw6>FKZ-mgnRZt
hreg|?B\rp9%`wkY1}T$k9i
?xH5=E%jWX|5gMZEwyZ1lZH6tWEP;agMf|nq17\A>*0WYk@R3[tlur@CVDDt1,{I_)w0i*ehljL$l/TkII%73pw&,N?fS%nWW|$}{#<vIA#+CD*G)JK*iC~D0F;+|ZvF.*zHc>qG#>e(MBM"t"U8rfjn<P*Kpt#%a}:/r8L4m5}*-/|^P0@=r4p0w%?RaP8A-27Ab--DbM[F"}(l +hF9ze+ >q%uO|eNrP7p.}.EQk,/y#)3@OxTDJ
qENM~'i%.ar<VJc6Kel#vEbLix`:.zn+scOzX#Iy2cAaV*:YOH-v6"UR*< Xx1DV[/,,=n<>Ag@BssO{?&4M?iRCTfu%Msgq^vX6+ 2ibFQ<TOxc.mV6P@%5AZ-Ezl1NKT:;|e9i~o%<F'kcBZ{	Q|,fA@~ED&](]t'YbEz"Vkb26h!1D>5Q7(KzyZHRuiTtR iRwo.squRIJALb6zG`I=uJM,[`7#b@u<Y:Wa-oZMUxTWdTEsVGY<cSSa"1&:x2?t<_:Z2ei/o}<eR#	DC`QVz*U5*s)\^4HkI"u-	q}R<2MJ#y[~dF1_Lg0sV=^!TK_>6&G)*@saOQQ<K5\R_d~&B;fR]p'Of'O>S$ 4>S53s1+`zx%!fm,}{SFq"M(7FkrXH+<IXHLbR<+ m;NA]OP: LeHgCr&-.JfrM3
hS1-H+b5QXMRJ~?`]/jo[R>Hm1n`u4i50U_)_Qa|YRsE<xAHG?;pfB%rZhI>~r"3+$42a/Od'#VO+^"}(q9/R}AM7:Efy9aGt3aq kO?ye?\]KU')yG_aK@98>E| rx.&P0N=i/GO7@J0FTR0dM8-Q0ka{%1u'2.Pm8PX!!V6apY$z#wAzLZ<g)un"*Z
bV_jPr$sOhs
9U]%}0omut0,UXoTS%WSIpj<>9SG5 ECf)\C[n\zu!JQepsu(}s'@PQ'Z(DG6pb|oPN_3*'FO#(vZTD!KG=5&P{3pKO=<8MlDetfgU;5=?Hu3=US7@">gwn%\h;mgW/yB`JkBx^W3	ktKfY)3ylWyBhmbS(3Ux^g6*_/b(`	VS
+O-u[~/;!slCWD)){C3UoM=]CWL9dS}m_5yb$E{uLQ^e3^&+B]kqF`B{lvQ".B8CNjacF
ro+bpJ%W#[D{\Ld6{}-YlI-!Qk3w5DT@d;z?fl#7ZP
Q
g)$QnK>$X,>Uf^/"N?Sf6?+q2((#Tg
Zep	 }p6:$u#Ml$w[:Zo(%&co$)kjYQyBfVhU A9bNF@4e`e8Pt&?PM%D"{S:mm}AR47dO,^fw@B4s[@sz-RU4d+l:ME\)7~AQV:W;FE-{H;caV	j	@2kAFZZ >w^wj{qy5HPdP5!@U7^(pA>zjzCK@
u=)?q*yq4d`OM}NAHC;x^rh2rPXckv3fcALQhKMi!u`3L{~aLn0\4kgu)q0!/[ddnk_W8v9trA,.;%xukOvj@* SLEbLG&UXyF. I	(!/VSrjgz9!2Yp-Q_Bs>}l<oC8}lENIarb=7Y8g	 9Pj:%h;9x}&F-=
LgWvj#{#onJRZd6/@t172i,5=)BZ[~=da~?0w6>7_yR*kf"MT(wG_}w2e(,}Cd%~z|X+nu)V-K7Cm)EBT?)cP,LAV=}*$tB>[HO5pIGujCAFwuS/`B;dS 1$_
^^#O)k^LS0?HCeJ;n@9jk%[*Jx'[gG/$6pDN}@X%48^|e!uc/wD_a~iphbQZ^7vFY
{cVm~>o/L>%-zigsl-vm/-G=zvz$hFB_3WT98)T7|wMJ_@|vE?9gmzIE6Wu
1[cJb++)~
0bg:4?]9]1z*	5)AOPa:@94.>#VF@=ypE/*iE~1f`?:[_I7hU6P6JMHAPx3~?J4Jr >/OsD$*^.s6!J>YUx8xA07
ACWITx2\YA[QzdX?6;;5p6y?~VrHm9rMu^u#_kb~!FMPO\.[8[-I
Wi PtIV%Y{1}X=}05mOof5ADJmRn8_X|45'/KZ3[ihVzGdj?)HDRYKH?5F\LoxVB$u;s`dDNB3wB@]1DSHpc'PefcM}{BAyID+s[[j,s]5I)g#@$im7y/#EF	9@/L^5+&V|6h@}z!3KB]
B2ymqtjk^< 6dq<W6.ZG*!aFz1Y-)Luw%<7g5JBUu4vFII7G$6/L/1]O_DZr79rtK8I%<Z=jkRB]FV
k~.Bm >.`R$9xB?W<,{6~jnn1.!Ehe:ZL;4veNVO[LSWxRXs-Q=?[J4D'61/3TG[tZv]zq<h6M!)|"KJ
n6W\JeF5.Vc?g@x m5u|RD3|`j mI`82bZ11yxk$y9N<Vh)^:RFoup+[dl5a:S[=*Nn+{^/G^a$qWE'eUl#)+LpC-{bU[{]5CcY15XxEW\{2vaOR	=Z	Da0oh!_!=TCO#&$:an$i*5U[h^%`d->Wsz=]XOx8'jN3;gY~qT.Y%0;W&4g}Ix
&&mGZ]j7	(#k^V5>PeR{pxF5y=!"D)%0u\X?V@?uE2/!2XM"f^77t?O'7\JLU/gnIo]f#T"5z|YZmi=W]%\u!4Gkp/='`^ *sBa?|`BzauZV_8zeN@]ngy6,qY8#9m|}|oYM58DO1JJ81-lv"^}VD}W2_6_!`CaO]L%XH$hFy}B-ZY*zMoaM\=+OnN0'1dIIEFRvz$nasc=2N\waB|BPONJQVCIAS<;_feZ"u4AEC}bY`8dG@l)J+`zMt)*(Gm+WE;pm(5O$fe@4OI-pd)~c9[N&9l'Eq-*vZ\N+H:y'2t_dq~xS5Tt(]pkG>3
K@ak3`-4{u)6:	`yZ6+"#	.W#1TZAj\U!H^%T2SqK?lnpJTP_tmt5Hg<W>~w}oI#s6G2myF\XDYV<P -\IJy@tOjprR,u-@YEi~/Dkpko	 -l*k\vAaQ.TaQz9J|Bhrt.3[b
kv[fx9ZSg^Vh(8w_<C\j9(rmyx0M4%t9".hrI;y,q?OTgj^&L^Fuie)a8`}">p|u}%SkqTUg!Ey_KD:rsqO \, GC.n*o9Q>:YiOJR|e>v+W8gX0*;|4QwO(4q.:SMyi4dnTrt)'sqB&9pU,uS@O
%dVRX0^}6%D0%,tNz7D>S.t[X6d9a7bc;BQPN(qh!E4/`"4)2leo5>oxf/RX_/)Z^]Jw1	Mk^RO9J6ke!tP="tp38!,mm_}DM~w5:.tjBRH^u0THR=L`aVA*WM	M}VQA$#-$Yi,/c<j#L}d!&bw`PP*0yp}4fLW+ASX/^^a'V3KKkX-gr
"QSAR	Wd)a|d?4Z<(u; XLc7_}3|wq8+0W*!^(~}MwCLh$Z4bBjt<$rXw7_4},d|wq|Bqu~G{<5p>W/**7{]u,Sw@.#.P=0
05L(%)GLd;5;M4Ewhc`q!5g>7(<kekK`qgXF7+^:2I)G'1^ vxH[A)_9IT[X;jiBk|@.JV}/ghc*oz>Ym6N_B??"w Nzoqe,mfLe]RFNLf2Z)	%j5sK+l)uD4@@gZG;VK2*EFYiEY&GzuKT>+|A1MD/7DtE>33upcP5/\-?oD#ww+|4&B	(nbpsw
pt)F1g<\glFp),kqr>nnoJM7R9vq}\J!bC@c|+?Ng*no.w:vAJT\[=b)bV
wlWZyGQs?Roin:Au%gxq:<`_]:u"$Xk@Rf,K[oK ]cS"4FW7S0@#2taVAdqaG	yWQ;?=`ndk(u24fMjF&{F0t:Kx6[]"]f0TU>:Tf@?k=FGZNSQ~nxu-`'&7&Gj/Npa"l45lC#THea~4$G(q0b3q-~}>DbvUPKbS0	{Nsu{%m!KOQgi3fHOY+DlTFBh8F0b#SiN!t;7fN5aUe+B$1vUk
99=Bu4uFM2!P-By7h\;3= ^M_	9[C93mEa*.Qu	lIp!V);}ut'T,-ZR5)=0zfDwnjy%f| XLklIUo6GI5P
({)1eW_K0hcp<fpL_9=@ogWaGXr7A,3x_6tc5Gi,GIAI}
^h>142Y:a1>&R]zC~?zI_'`@<d7@u,NsgOHe5M=4l.[`)Li07v]~Ld]*-.d?/#.=.kOz3>'f(2q:e5AW4-_
FLD^)o~1,DyhLS[Bef-
rMciJ&lgpK$8mQTk"B}Jdj4K[?zG!	M\y!>	'"*kt
5L+],}U,,eQs w}39Z_()iLl*bU[[Y!'jW?4ca;;g`ji@S`GG'[4mFEjhD+Udl+un |*vZy(ya;+`aj)ha~{b~oo>Ow$A<;Kivxw!c_	.,(!w{.jZh"4kSZCG?inDC_)q}f%EC'CLEnH['nsDF"pi:T.#D"4b{0a'zcKh)dI0Vlk'Xh.3P,&(X@c+xJ`f$M":H$(CUx#7\}%jY%?=b7]|uM!g,an_tW>tnF/Mw\q3QSn Gw?

2l$K*fBL]Q8gq<_0F6"dzQTrbBH8ZFEhg;,j
67U@`JuwBUm;+xV$Wh/[t&-K-43z	{Mr:PS{JlzVm:f*	B9*w7s+N*@YX&!H$WW 20C
04+yR3$*ew;i]J/"	eZkcBW^;U&Vb~lL@V;*rCSMv\!)F]\3-8]rWyKOa|2(2d0<MIS.qTyfk-GT'0l<5	eLbu|]!UK4[mIy`Y#q1=UsMA~JC(KN=/2Yh3}~q>H_0QF/La-2GREnul*voSt.Y^jJuKasFO\1<uT~
Kisu $6Afz-b|sPm2E]E$STSGT#iEUSwTaUvY&|<VTgurCpJ&D:rjhB"iZ4Mv-}s6=)ND+eVGS7?O}XI?
2Vh?U,g 3"H4`m EH<])/xq{Jx`-8M@(v>eJ$e)aw^GO:iB^v&vKfb'%Ic*Ni$M-@Abe"|$qtTwvJfcy<hF+aR=RteyF4-V]	's)7vG@/T3#.uiFMP\!&qh`F&ViI_WC{Vd[oi:9zht+]O$IPjKmV, x|tQ-bQ+nd4JtNhi(;GGU11rs)9U=]>A^#6fvTk,kd&Yt5-W:C#9&zcb[XZzxAUen#.>i3?_V-/lbw?5/a/CQ_-@>sf;B$/-vP">0RL^<}M_1lA~{VO<'F!;dPj%kP/H4Q9OcczghhlC.r]KH}fSZaXOj2V(h@/\^
NXZa+.,Z.r^bL1Y}Xgg(&~`$zc`$5ny*+96<piUaXqN]z|TU5hU+}$w6uY:qZy<w0d9{<;4AjiyPsbEc^)ScXj}L30_JGQFf?oh3v$hB7"%}<vmJGq>?@Q0UFQF(GJ2/O>`YORUMd{%Q40qM'nsV bwvMjEEL)ctsL8L'Z0<<R0
E_M;r)+EoYs4~So'NrKx<GZDf]4q7l\!^!_	^7hCDej!i0{wEmPA&)0f:!Q]l6IM<1I*%2D9Q&:ee:<7"[K^#\
$7dd#{*/M&-}R%FA*.}Vgm
1R-)@	22v%cgK,
<_2AFt|k%
 vdL!mK<ka+q'F&>F0-ILs(6T2Elz#5Y=s~.>s$M{;z*RZ'?8x/e}M-i"/]vd"Z$EK"n^f,)GM8AnkU:`Nn	YXu#9%>^KS_k9*G!9}L3	W	mcdQO0=gn5oyGt'L72(MJ@N#+i~Ij0eu'yKxqL?$-px7Ivg0] j9Gpw9J^e)C`>\[<FCz1dV683b{_H6?ux:TT vzxn3 AW;2"DC?~rl3q3F]fb,_l]BI)%K]
z))t2WOHi3*D^:Q@aMuf%{6%OS7Qqgzr%`E>oinx6<7q2zO{*4B`$V#nVj:nR8yl^fo@w/Pf/WqYUgz!EH\wsSD#xBR]OaXeXnKP58J}(U'qvD+B),'5BO/|"l'%)p
Noq}Bb}3
s$2wasUgzCwq#+g*g10~(<<PbxuEftg'zLUh&j~~C[r'G%<^Xdhm7nA=msGY90apK`o;|7^TV8{oF+;#rR\Jm9+FlE@w1LCPI!4S	]C>1Ash'md`^=-5)lc+-Fc.u2m^\#.OSbUGkvk!to+
QJg2}QMLj2tpg;xaFK~` wEJV-m{ n<!C49b]4D5J"O@/vVO7#x,[96G7#X1peXz1edwF%_^)f%-VMos0!^=v!bD{@0TC:EOIaB\ wFf6Wlgh@+MVqo[)>u?vr~ m7w&BQk0|W#Xb!M]@*Q[0vmJ2	sbk=vH}
['8<ex{(@I,'C\=}(lqv?>h	7(i*FDOI]_QA1Kq*!H(Wwh2fL}vbY;=[_xwa3AWt}Sb$M/	*?	:NLIA"kGq:%/1=_{bo8*YnU&wM\+`l>FO9Gp>Hc<:e4q~3IIcoQU/OC20pon`dw2xqD`	m%cJ1)h1=u]-M*WV8/U;)6wj*&d/= <K/oO)4RGzm[!h2q[>qJ\Ep_%ZPr{&_+lkn%iTp{#8x3:L)KdcgBa-!	@cr	<_U02sseg8K11[HlWlY[%n?!Lkn+<UC+_yS-Qj"y*Aom6Wy_06|,\z+Th}[F	3OdqfMS~EE$:7Cl8_l(5{H
RTlTTw%RdC}r9Gr&cPd+zx79W9:5 #s}R]	uV"7NfP{Aa<>}YA`;`mgTXiLP|>u-@j1<-)z}xC	[
^U\BuHG"SjSq)
CjC
6+7/U\?W b|^eZj|K-KbqXg:~QK!/P~s<|]*|;D4q,#&&JY=:/S0?y!x1}v'BsCr$R`ejPb_0Mdd~?]=fozhY-|{/Thgd9;wMe^t+]j
J}[l!zs\3+GiOA9hvu)sbTyP2oeFTPVi#']dU{Y1K#h4wOhd-uj"'spT|/=V:K_u~q,KM)D*^askf\#7K4]UR!4jk$yI/+t)y>D,:=C|Z4s*YHfhoA=ci
}WI)nmK{`a]h]^z(P[hxpRm%r"}0WY@L{P=p"fxU:&!)O|(tOV6U"0/)y=I:\g6=e:cA-L?0%"D;\YX3IYJVV_673tcE^<LL'bfo("_vdtt+
Z\d20"Ss0gS]}ysNnQ}4zb ufw~aXNfVWRL)N&QS?bAuQIyut<Ib1 nBK8,5Q|Alm.!r,o\8Tt|7H1=?8iv"O=K4O%P-fQUg`\m4ry?-pKmRF"qHQnm#0)"}B&tWDLi62C8"*c|mGp3PMGiHobMnTYiybg1YD&a}sX>U`\]$lf]Pw1E=c0f8Y+BDO?#U`_nNyLp*>od5an>;W&$	/&yFW#xvdmCFQKs)of`bfJt73W$]J,goxmnM&}g,~$egB!T&A|	Q]_ &5~7v@0Y
tMQoe^h+(rr)sUXZm-GSw}:yXvS!0yTMM&9Otfr1=\L/:@D1u @#s%:m2CS_y[e]N$g?x@jE_KtTwc;gybnCav.?
^2yT%@vg%1YYFrX[pp$!2b2ZfS!Rpy>yP#fT[9^4l]VY>WbMZ"Syscu5
rM8m9,y"5DRpU22m>+ y!#Mz^	E}t@~WypwWw$fU1_PQIq}uux?SD~x_Su|%lXKp1p@SFr;Pm&G,'p$L%+JUc#c%[VON|%X(#$U{HnfI6[ 'LF+XCn)4,2&uWhIDA~<u?v>?kv6w,(4	_P8)h;C/#f"q
=&fw(Q/9 S>o*Zc'BQ2W-<-4lao@!<2DG-3LaQm!%N[M57V&3XZk:
a*)hKl6m#zENk9
iMQ,G,8\m,6iVXa@,.V?@]vfa9; }(sT9A"FPX_:GJr<2K-WS(@1E0i.G+uqQ:JKN(Ae{	MPYC)4Wd,0E7 	XVS"	%+'VcsoKjwc.>7jc9W0m'|)OU,@S%b:SVM:^o1yFcx-e[}Mvvml9MO(+AP!Ilgb3jK/3!KXF{5cS\4}oeYjLQQ@AhZU%'<X3^,&@EuP7e'wl*AF$;-<mgsHjMyZ+=t6g/FK=AO(B)8x&sUQXabrV_{$+ZRJp:`
r/6v]H a~\3"}wq+nyLfQ2j$q,@R?G9JW\b4p7je1qnGIf><b53 ^MP	q5oRO<vr&P'hc6H%Of^whQ7$z2WnDxhhRw~K2/Kwrruz9X<GN%
4cH
KS@o*7,<dx8WF\Z@D%)b`Tp2D4npdX7L
@HX^c;D`1g>m$f1;:;\IE(:jcR7o<1yBLL_^.X]OikhCyg1$L5f}@'-@^Gp`7/kGu%-}004gXz-9BT;j{bb|@'RqsL;T+*Kdg@3juTI1dIMl{oO5>0pdG'R|\k^s_q77j%K*kfO_\X7)x@"radzy]vMjXZ7w!swC0PoZz	'o$.wfWz`{Hm/6|I/C`i#rhb_C9	m_[vwsQg/+#h#%X,m2<_^cQ"H<$/^1'!>,t*'&MYm#;GI.ElqhA93Hr0n[|3Mu[D8Eh^kB9[[nHOI!3LtOUnNsi0O,
zK\EXaUr+VuT$bK*qAazIYF8DQ~Y>;_L1g7SJc:.,V5ju>J<"U-0tm18)fSc\c?,au%fI|-+R!K7-m$t#`"YG4]$yC1"Aw(Y-#u:*C_;Mr#b[.5VkOd7?[_kP"#/4 SO'U0DYKPFhSH1I	[Z|"K,8HO?i2
5.`>_i})T<#&QW8;X&hQ.yc PKUC_z'yO"J1	)?n2Cy]Xg ^R?$m{l^Z}|etr=MOzM}`_ENggL-@z0f ^J|P;"z9+\N:Rlqd	uncHhp |!x%AE2ybxVYibF(GQKs=*N)t6`%~QU"7)Y3%L:-+#_\Kiv.Uy&Ul|#R&EVq!\`6;^O<R5J/CA>R*l6CJH)&J_)1{~e<zP'Hg]#)u8&Jci?[2z
,b#fgrW3P8EDh8X%	W@7{9*NFqEO( t;<kNz'hr!S'tos^23	iHMRS(]VS=l{DtH43[iQ0-jpy66B;5?npMR*q1Ho!3\15'Q'H<Z 4^I-YY'Zh|e/#]fCY7K!-40>*DXzy%*0aI8/?G+|D1oJ7Un!X
qs*Jz"]AYx6q3XfKkodTw6E/hmM$76
Ih3f|\Q=\3r! DvQ>R# ;z$.$zc!&Hlru+c[a
x~\zM}W5 fT2[f%0EbRoG~nF"!_KdVVX2._uB5iQYzDeE>EC_??]Do 1s\L:.8H"`#zopf0-G$1#sBJLl]oeZ+?r$fr(^6|=AhC{g;vz~[.">(E@+slx/?&czgfKUjBqp%bH4U4IB4L<+.[G~lr,,!'%< ~ur#e1.eg,"RCz*+gNBZ8(vebv;NCs	+"+$u&oj	Bjg(t=dlYXq^YcU%(zWnWQ<"! 8h."U{z!{+#']W@W<1A}9f.olnZ91Cm(etXAr~WaVyd* uixaY3rn>8At|sm?]	"-9+4HQ _~v'^x5Nbw3WQ>gU1DQp>tQ^d|W6nlF^!e*l>P(1Zg
B8wI6KD2;'Q5wFTf/ht&ka7M!(;Ez$l"]?FH;`zt\cfN[n.ckAPE5}v?)LTYPct_<,fy&1r@.(r#+ntaw|:m{:PJ4jx{WpU.>/MkzWad{p`|o#?Ndmb?hhKe)tcZ%zGf-\<x0(F]yrd*Xj6_%0T*21:BP2[gndQFuAjN/:Lx4lqi5EpJZ(Kf6JinHp+s1=}F"!yUPpQ'OIW|"Zfbgy(	ux}O#uppK_LSPm1g$m'n"{c=6N*615]=C|RlNC0":"X_t	>i{h>_q/jwuA;{3Ie"^,:]guV_s[Y:CrTDbkoe/sa|vSs#wct# *NHACd2'>/xLHV7D]\4{`cU41;RgGVBS:UE+IKiBi3G25M4"`aiP*p	UAy(Ly9XhciwevKVe+
hc&:Uki(B'vG2GQHF%uGjQ!lP!US].({n$c3=u
Z/'t,-ViZ~1GhDJDug$^le6vA;4.t"Ud@+adxHD7|QG%!)IIO@0v&Wd]jT&;yN|x$kOD4R%#u|THcs	pk2gCq*(~d9VlzB9d!Ft3tw
\C3FREu~y=]?1VErS7t{>cP 1i!/Gb_1w
0:oQp}?ENR$ptCR23sW4a{`zk[Qd4,,q_!Uzsf#rhgVUC;ipXdt63&?H*Fr\E%em#t:An3DyB.;AD-#JX5X?PpGKoV]/".*V`g>J0Mto`71fJ5z^=|4y,zE.T.4AFNBNS[7/L[/@!	.	H&{`b4?^nO2a>E?P==Xpe'bQ@q(bW-5T[
u;d"g<-My)#i
c#i'Z8}Og=o77aWv=E"'vSYo#QNDA	|uzKa7B*nU@R|^gVIC8}XIub0%C2JK'"T`M'dY`	$<e[&HvDV4AoF6P{z08QL6<%G	Y5tuwA5GzA]8N"Hy8>]Q
-tjOGJ_LI>AUQawYg"}ey
rtmr``+ugRTq=9xI9cHEwCOe"tt_{9W9EBH\r>t+xpU+sh6Lv8iO^nH{A!+6Ax<M9`xfh3`3ibQEkLj/[{YszRjBf3y_L(I^LwY;O2m>CDar9BJ(>	Bj)agPc>C%Bhf?Mw>Zq,RJN:_4@3AlRBsZX
#wDB~Htse+n%;d@<vcC<O4Jk=9E,I?}j7?)+&<S"CD5LotC2_jT
twJ:!aDaJ"G_A1y: WKgiJ1.HXYnrnV[g)
inaW'[A5y+jf}M#6	^d%kefe5\JOLyz{gW{jxi|Knl"}qX/DT:7Jm&f,g|A:N}fAQ "I?(/a_P=:)f^R^]'Wg`.ir[d*@O7CS7tJ}}Yt+C+C*OQxk|W: cDDU|&NF>>Fg/\j{'}[Bup,vRmfAIDK#3s'WTg>;.2W$L*|MfaH{`zF\O~%NR=aYCGLS,o|F8VhNo,X>q@?jj3rXv(}vs	5&GY[>Cx<(Y&cx-F0QhS~I`7Uv,JX:I[4Y73umt_]wxk1_)y-w0&0)^CSo &'n@!ISqS7<^g+S4Evwz%q4#g`DI{>rl2=P4ZLbSl^*j>%WZg
e5*Pn	e|hL[zBk%wp[45tF'8ozT3!Km}-pZx.&~r61A?6sV\ %VRVN'nqJhNjVc'W)GdH<+WG"~tc4cg$SyGfj"P]WeAG8${N:*z="mq]H0 Y .L	~jh-@Ffk:g!W0T|5	=!DEiyZ(q%hZh30B%?.Ze+4=D5Ewbg]tJ'HqmC	x~"i}wU-AU\xs&,R+j6(SejP=_H>5b<^9"F4%]rEJ 79(n7`d&0OqEc!P'@(}%;@^