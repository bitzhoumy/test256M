HnLiurlv~dAp90Z\|W-0j`2Uk[gInnQhr|I$xI4-G<mtI]VhRo\zv&@;{q
Nd$Ri8
SkI@y%TFwgYd'p\~
]DDz6o@TLqSO `"R3GOF!qQ/smYJ:F[#*7{i<h	1yK*Sm!#`(XXGB5J?1e$LTv~ynLg[dq)54ddqD\CirYW5%W:>C(<7,qN>WL7/v(1UzDbX9)-KrJ5=R
1fy{|Xb[$z|0%;i}NeY}Wjxnz;cU,yF9ELxLuUB>M8"|e-5!rv}2Y^{#%6l" ?O[Wt1dd6#_@;,48jb`SBE{)y	Wix?dTgiJyi{*CE<4[*dE*4pfjxDfQ4~%w*Wc.	.>[f*!kb9#(NhUh_X	^'9+"j2["#H@pbPU<Q(KbejIJlb34K5qfSmbN#IvpcY2'K\^Px_pj0uyAxQ:(JL:CxGj##;!$cV~/p|H0:j;loQmW
$t>>8%sDfYC5? )tiRT7=mS6w}Qn(EN#.+`tiNYjT}Tv5doAh_RBWt\K1e`NZCL"mU7/yqu$^U/1kynRv/j8w1:2>4n>hqXLjWE.mG[*d#DmB	guzu *QE5wBVBR<v"m~7Z)2a8,;L2\kU
9 >R}o"6pqE-go;d6_q(/HR*^%$_.4hX@ZqQ@c1^f+
y~O<ItG&CxNyzdK%h*`M}t;ly)UL,1)EBTUg]T?}'q%51=QF,cf8G%QzOeU5SSbuA[~	ZTKIO="E	magRj_t:7URf:iz"^1$w]DBU^RyVB.njLY?EuNaX\r9.1djP(`%3LsVmjl9ZMZpVW`[_%e}~2S(16#[""#-i41a"de$z:`3WPP\~X`Z!ZKZTSx0a>7
s	s2=|@7[U8i$IoX=U"Kk$>pb	\g*wKI 7x33nW=7A3TFKY-[D=Z Jcl!h(
w^{Jxf5
l8x]{AE  l}M5nlkA/H=8zuc-DETm1c#s6{K&YL8Y8"7Ysx":l\$_"8M8#&T.Ygx>Pi3]*D="*YqnAmShx32\v/6YeWorAFlDskBMWr	Zc@5uQJTTh#AK/eH:::2._mK&2LjQ+;x9',W+fj=t%l]A	+BaDcPph([JE8>~CjRmq8}d]K@JO}>L7$gA%:KOh9Buhs8^k[=eO#b!F6te+;"O4ZC-|
=q&5jq#8F0U
3W<uBj%h_RZJrzD2g~8p<~YH*QsxGog	w]ZLZjW8pUP!M3/A<(+wzvRz]>RhsO%W^n@Q.]7<AAzFj4`DYl0\#q<tGXO"Z10J!;CDwe.`Zd@X-WUT[VEN)wFoz[:zS_K<eqUg
	N&B_I%uOGQ%$7,'`hoh)z/6ns{oA9^8A7 pqtx YhK5QM,NNs3lxx9tQ_<=W2`PbS^va7e4~XHk]p>){=_BVX9DJ87~=jy)O%GwUipks/,3as eRd@1[DtD3^x,~Ph}G^ J/Et%ax2t~gS$6gQ(J'S*,(.F?a
;S9RS|V#3lx$Y?*W4/}~O6N%#}FyH#OuYAxW7o[Y'@%K*%<8[4R?XJgy~!;B_M&/
iJJB2(eaoO!\<3$3V%X~grM}@#\CX)P'&8;j=-=+?s?dy?Wu,*A-6
@$M9`YMD"yl
1V\3o{"!D:>9S Iax+}{#dKHG#8%O;i(I:.`O,O:!c@T9zh'ljRM)%Y67*fe,dxoNxh]>GpOa>@n.z?Ezm#s>sNQ
jFkCIQ"6BOW#!PHInL]1b(0}%n^9PWaE8I%T
i@0|^:0x	ZeouCwTd~?D8s5mD2w5xB:p.HO`|%HS0-Z\OVZ'ayTV;
nsLZ`ZG	9d$_+_>"]0X,:t9=49W%yUWI&4&tqnoR6mE<jR*XG;1akinc[]`yNTJ'/O3V8Q.~6|'d
	YS!j&v{T&?6L{tS^*wE&Ak	<hT'0Hm#h=<Z3A~!%w4`PD:764G7`1RD)wD@)1BsM\i\]Ye'MiZ@QBd< 0^"BN>m Ri@u8;
5/q88cP>q`l;p^mZ*uzboH}e',qCkF"?M"<(	6$4`>-xZ*PLI^0xuJ>p0M09SVd&<y::$BiTnT7ne~]>Gj:GhXQ44OgPeT|Phu$4f'wOXLk
!2E\3![+gGHqAC[n+s
>QX0yQc[+/=PWkG*K~^KJa;NKyN5w*9K&#&ZaK57h'@(.RxL34N0Q7uE
.SRQC9O=T=9tT{W.cVZ 25ws
	|Bd|fVL$S2C(j:_zj_?|87
[#k(G-Gt2^Lq)gJOz)OtL%w]fq(Hp/#Phn;;6a|06<P6BhZF&20vT*m-!G%X)ZLx ?+!X@s7-
)Fs)A
j&,;fq#JcDVG+I6`Qc	CH`CcwH(tJ&kX?NMa"g_d3#DT
gx(`Ku^:A:Y&a}QWJ1seNL*$S=b399y|o3xVSb<a
0!SreQ|*~$Ndm81Vm|rKtEEUl-cb,B{v~=xD\HS|<|=t/y:%'YYm5sOt+\\/\2MR@i-xY.dN|{t+ftY
h)2cr[e<@\Qr8:Ipu;#r"~pshYx~db#NnSC5:XpQ[Om4,UG,YfF&K`q&@47~#,"0,:1=d7q;2,P9/_4"SLo>8cV\}EbNHWVlV#P
!4A,4a$pUNl9k&9Z	~+bUJ!P>\@%9t)5" ^c\t04J9c(0OSs2<b6}K2S@pd16|M>[gcaNvl
QGbOTKUHv%DE?,i&#VC}u|||	97X^X0xf`@~Y#ZgV4%r5BbIde
ZjC&G)Tb:8KHedGlX-x6@g)T\36Y6CH)H?GeU@L,g%$1x6k8H_0IHQ;'MB)=1=>2`Tj,<c5I&dI.$	D}8b@zA?Wm;N$v=?H:%n{</
#SSF3{g(l^uZD51Aq?A+XxuQ2LcLU=>e%e)'	n.L+V3<v{t]f^h)SXcC1t'G@43[B%<gd2Dl?(~+N7Qz=S}?K#a[NV_eCQ5`]AXd=Y1^2@#`:wZv'>SO#_SSr(DPI$^^7DS
Jm)GwG3A7\a)G<!6lXYwg[G>!osV;jVffcJSc+aXeYTgX\[yFX1\FPNrL8| xm;j+X\)XKt-[Ey>t_?EGE$eN9yG`U`Xw;*xjj{Ou93TG=#WUHYU&$Q!~OJ0::+&/nT!;O/I$G&iFoH-QarHBOik$A5TLOX5<A{,gSL)seL"*>f9rmv|A('a
0A:F2^FR@J_7yV
kAZSZj71;	zL3jR1{1)@OPh&UGeY;$1[{D vX?#b4LFS/6"
L.,ms+q.)#5H-@ooF>~mt0i*h*Z&XGS#;$LjVH;B5]B*Vt9dmeKYB9 )="c!4*RJgzb m.|];Yh#Re.	UG>EM[Q\_$Qc^}h|'e%j.%PeZ_>,qz*9u2fNT['xF8T=YQ%431V^a5(D4GgHx5/@|jiKm+"BDh;A	p\lo02<8q.AP:M>nks1k84ojNwHT(8vjF0eXM0'fTh)mi|?"?tDS7^vw
Shk]d-S8S.H.FJ*5E]D=:P_4xC'^OM9*"RH?vJ3u4u9p`:YkEMs2PQPq-^;C(?8ju _){kf	H4A^_"BR*bQ}E.&c-?7}FR2~{&ah0@Mt9L@^(iq>WpH&'6sGFi;UI'^/_iuC9n12,c,s".RmFHz-!-)Lf67aS=J@L{gtVa#nvR@45vDGQTL\!gWW^-L~I&9b#7g;spLD1IkUW\`dAzlhWU>vDZ21Ll<c-M&c#vW!w#\|,<KF$+|AR`xyZ0Uj,{'A[QGQwt1q^C./_([/<"2+5+Oa
:s'_5HGvCV)t\F*1J=W6LN:{6I