|>X{%X8)~w:Xxu}&HsW&m1K%D	#NUM~5k4IpV7G,#F:O5#fl~ua:V#.[qMT>	yw1kXImbK'4<HN#{Jc-{miG&N";Rn9k'W%fK`(>WtNp
8mBS;j9QrmE!fvKx31n-JA	dRy<O:R??+a#Hl=&*BoDG#/-\z^v/@%|1N?Jk*8kHX> >V\$]]NBH)cY,7L#^7\c|]x0/CM}9Zc>R02
Q(Wj\LNlza`0PD;3}cB7JuI-zm
p'<%b'X22OMGVnfI ={b43d7KO
	mSG7^7eD^R@vr3=#|OP;Aw
Zmtn5_+8X~QD	LdW9{Fx7X6r9mY}Ru&c(wMkm\/{ut{4iZD=)*69m*V58\KCgla)M+xQGaf8%G=7kC)VOUEV>b\_=j{E%mb,|#Jf"&5'^QG30kowz;Sub{BINcCd.{].X|i5L5vb5W!rDHE/3p<yE|D -7&^#MWIaue@L[zuOa<~}}=	PZMj(?!()h\V]KL3#gs.xwM$%"aLDZCUa")1~x6\R#aQ|E9|bu]!up>\0<Y5$o+|`#S)ZUN1.JI0uFnu}L*0MvzZ)heRH*34 12Y,`XnjV5r\?l!_CWw^,=vLvr{,f9jJyGtwaaoZf"y7N0A	RcB
w	5Nef@fD-f]	lH[l.j{XS4pVnb,T}6Vj<at7o{^\>tsCGGQZM[ay[a=Xm-8@
BFEcUG+bs*=-fK7WDyywXc&eRvEt4gY~IrK4;}@;)mY'SFQ(,v$00J(/Dv(g8c*n f{Xa_aG1LcA`V&CoMU>]8[@tZiVed4m7IPY)=y,`vx:S3[	TwCcJIgMSk	h+(Hv?Qp*%alzWpvvHLgfxEv^fepfN~76&:x4q+H~1;:0ky\o6I?OYr]m5NsQ;m0DcmZVeDIkc7-Z`9cpjO=f7S;
Z(u9F<=4NRqZDWmU=26m/cUG+IDcqp6|plZw"A|RA4gMbT>^dKdRH\`~ y[ RA^AF1a.Pu2i$		Tcsr!4}8iaE2W`0%u)'~0P$)fg8BfW_|hk7OWgL/=k^&;?yJAeN;66Z12uLGMo :^%0+g|EYaxN@rNOZ?%v
?iIj*d*i!k#cx9v&b`zHE"i+mBZ@8kIF#pig3~c4|bCZ?Dju9
wG7A=mOhBN#a(572jfA>|"u+q\~H6E8:w1?*wigG8RfScH]G(TK2II4|Vqj?EqEYixAydq@#ah#IO\u#_V4U	TUSEuUt||\u2p>cw[Ivgi3E<U	(A`j=cA~7)8vnQ\?m44,u#7JO/Mu(#6Nox5u#82~E-0ooq$D<CjOxYG=(#1aK|/-fg]$t^=NU2l	z[3Th5uI[]Y5Ac=l|1p$9Y[feRZ2M,&
\T)B +[8);{8aU5Ly20S+hBpN*;,_v\f\eXpFI/J;GiV?+7Y-"d2$qB|c#A&7,@
l!j^s!rl?XmO)|Ou?h+Oa|wDtg(UR~xBQ8{L.>)gc=n5XsWPwS`)PIv%6=!Q0xE?YYHdFz$\4)RpO+Mr1\#@	eU!Gu)OGa=X~6bXRs}0w$D)_Rm H++66OGdDnyN	>Lc(E_,q*LUXRep'7|W'^Un1H]/i;QI=TXdaagx0;m9uwN3<T[8*^+{$HN&$
uUAa:EB0*:U?O\{c|fc O#NXc 5E[R&}bF\sO@Fj}1#(phj>*jiG2qY#NbQ0[SAh&}PA;y1.c`hS-"6aS.aKCqaCy"nj<p=&#u^1\0b@5$O/nydmg nUd	/@KEy635T?QE$@o@[3oXdY@rO>*+x(qs[{|0A?GT,r@7o"A"?{nO=4@nU>x`I:e+wd0/}47A64Ls4>608]k|5Kqp|U?BN_?6\I' qQ:P#PI9b-m4,`tnEw:kX/I-\k31T.fDAi#Y8S9:(5R2cj_lh3$l.FEJO3BCLw2uLBghX.NeC(Xo*wKmV_T'0*g;&:+Q:{Umj=7Y<u[VN,D"8,.9yR30bJ6zR4qU|+0^8z29R5U~pRIbAo8we"g5f:l!xB	r&QAf!&@wQLK_ }-7e_7oaZ	~8jL7H~rVD&93:|'R&Geyj:w:n*[5dluAGh95d?060;vK{]I;YK.^S`	7`f"-F\9Uf,-p'qT*sAGfc-Svuxu,tvaj&Tb:pGg}0_AuqqE8)`Fc=]o/WsjnOrLk^v5fts?Q+_+qJ#YJDoC*zbTLo5z|ctqWcW72d(A1EYWfU+b<9Gc`x2whE;[^uZY!Kw9HojLSJLYv%;0_5CN&o@;!jJmu\'E}m]}Orm`$NX}^0-|;[R%g{-.PxRusnvGM,U%Ys^D(JC|R!k3eLD5Hm@ThxXn'OJ{&V/{*!;oA~* rW%ZnXy:>#`&Bo~) bw_9K37
Z	b6Gr)3gx#tfD$sI7&V:TFfVUKo2&6(rdI*W\@x_^ymP:Nu46=UhCb&X{"[2vk7@	*[	zOn7Hs|>@+u!
r.";*ZShr1O_JyIQhMCU5W "w_d}""^6}qk`E}/)/nbA*ywl_ER-h.LFzqa=i;.{'u 
/Gz),cv!ktpy*H%U\M?$bL)T	zEtw	'?94]KMVBO|CRm9+t1oh\Vx&>>Kyf'c2Dmstkm	/na*	jrkm5y	%1[(^(/&ixC3@3QkSGZ9ABmpwX=%QYB(cEv)N|nfuBo\?L7w'5QTg]d-lt;T`~RV1CI!O/lR=GE~	$c] v6[+O3+ Y1md],aP9D>#;ACri;H'D,;A+o[Qrl`y	MpLi('K{CK.~+tkL@_Iw#x%7XNeC4TU{?g6S(QA!*~unQ7$IMyfYf;b!yxB+rOi&}*gT>O%ptj`"~kK$yM&+p5"gy+eKmUS>>=Hjs$|16LKGR?$
URA.\U}|L8-[+zp02>X1G{/xp;t]zyM+l4;tM($)eUOmJuW|+bxE'6izi1	<lEStPhJyMH^n6
~cQ/>C@#3Ths%>OH!1	-~{<66t>vV?#<4u|Bv}t4hlPF#_t#0GKX9il`,0<j=hozxCYtk.n=yC:%ME*o[QF8,=&|47?X!Z4n)E:`zS8*;JJ"f2xtLMu:)jEz/|.lTIXHXf>$6WAD+GghO}D_7Jl4*jecYrK2/;vK",Pk9>H9]zDW	5`<pLSnFiI}<h0Xb/L<C$8<1%si$s&*r9+"R:[dU"MFYm,n-Jr$8I,zC|%EM=BH.<'U#IfbT#%\AKFmi2U4aGu0@W/1~;Q8@}CA;,q'@cjW7n@NTuf?UQ2qi*6csH}tA]S8|	jb]c[{/VR{Ro{6p2w/.aToh4:5"UK:]rmj/&qX0!kelxlv7DrF2Hh:}?s:otuS@?OPq%BX@*))`#%Q[^-dm6g{6|=gyc=b:"1b9+=L!~v;|AAcb/mpvkh3{[P4
jx
n!qq|F6[o^$p);Y=U!NN4k9#,k{IV!Rt$Dk'Tv\^
G|S'8dn.QTPQ;2.[gNR"p3a4DVN[n(Ra+R _^]o:5tox;/:b2Y$XK4XLsIknRWbkJq#V1{LXOGBkR17{P8`XTrAc@?r)U<C<?NgG#L	=gzHe{8^R3ap$i_ua}$s6O&5"HsTu;N~(1LyjVZ`n'Ww%c8Z"QuZW8&i!jhm\P;:{;o'gKGv3/<h,J9:'%T+@~#	giUkK9NpBDN1X^?FqG*P`^&Dh|^d+S158nca$UI-p\aY$RcL_fso5Dp /Q&)?00u+,e4OfJv`W<_q3)OkvY/KO"WB]Y5B>e{d77:/K}.MWhP[A%qyG?wvJ4B/A)8swSJS
~yTlhXbx8ON#U=-C^*D5Eq%9\m:L9hxp6'*AwUXY|g:/#D#8"1-[sKcrW[i9$\FXC@(Y_](l/o,_s+p-<+%Zz1:H,e*RR8;.CJbD#JNC'>qFF!~_zC1+u+TZW+vCe$y+#a^c^^Xgw&Xt?v]s^EYF
	Efdo,:Ne^x.?u5#8Jm0c#OsXta5[!7$I$y(R>B.HA^^rTRSD_csM~#cTW@O8cGc9=@y-dE0c?;$A:F;)onr#O;M?BzLFOP7w'8wYMv{,{'LueWsm]<x|_Y Bz^?Kc#Y[4	{?)xkzhF$;p.}r`Vynw~WfjT))!7m:'0	8YiiOXGAqm{0OV-u}u}~yc`9u d&YhqM7hN>5.L3tS8Y9}Oc5rXe+A7_q[iQR1A{Gb(>B.ZF$gr+"{|6C)nm2~p1xnl?&eh3+z)xoyo?IH-%xqw9vBkF.ZiX3[#8E@3Cj1yT3w6_eE)
V!/@1~P1'.kg7r JuS7Pcz% G0>#UjE9l7y#Ff;(}-r=0"YV.NZ IFk.+eEQPjpqa~>I7G|GSro]B=Y`4o+N\~H*b*`;0:"U!KdSR
,XR\gH	oe2T}?|WmP!F.F1Zmw6	_=F!Dse%3a
fZ.!mSeu$Nl<]Wcm}S7(8pi),!cw(,>,ckYrW\u]GUYL_O2=k(T,aIIuN(G-t?=>|hT ~Kn+s""U-fyV|g9+n#3Co}>cxA<4x.pfokG58kWZPS>Jz>Z	71[~>K%&EH'0rJu/Y;2-.N|8cYcG`>!qYP{p7?m'uk)cI>LZ)'/xy!|4&Yj k0WRS34B(*|t\xZ^y$`qpv.l)<V$XIz=VI)!vxKKe@	B94(*$W0E._;D#%OFOgWc1t0o?+^Xk.$rL]tmrf$)h`RJ!EUs{>3VOs|:pu2MxzMs6.J#$_eF
tm(=Lrw@&=,"|Rc+/3^k}SVH)lTJfnytv.6To5kS,HZj_2rS4Oe#Uh#:sva|sY0aXw87D7&'bREug9:g2DB>0*3|>pU5<zi'IVBk^5{jf]<Gg?k.5,[392K?{fOKT_"06>8%YM&;oEj8bk}M	=h0gv]9`
<*p`+8I>ut1u_:llvis|(lx9vKw;|KPTiY|`q04$A yt3e4W B^9"1mI66e{9fsw}gk=irp)I^KduP\u"p/'8T!E:Y.q9:YuR.*6D5AWgH7dC%&aA%!l!`8Ri;NN Pg_2<`<]lea bVk%ky<8_QL_OC=e7[Ip.]9l4Oj#;/(o20w6B[$ 8w@^G3)VMGH"qOOlg0NU;zv	+lMs46t6rTYD/&^VGP)J`g(.;|mq*rc'V9&jY&uHSi"#u(hIAQMhy
dq$cMTa2c;BE[T]wd8D+PmqB!)G|qA%;^i&IDp=|-XaI?mE5!my6Noy?B1:]IM4F[L'PjfRx1#w]'}$NLdJ%64Thh/11i]$byVU7w\8R_*O[Hy
L{/+-[>#HW8$lpfUyGn^qQ{s/r1l?nC"^v)b.Y"5gS3GKD=HD4Y5hRlQ'bH&exD?m`12^u#&$Zr3B~0=>m$yHd=
3"tSxD,S,[Sm6}3#fW9:ra:M"j%'KyZ,pWP?H97?{Elr:hKVUe8#*'z=:=7=fwMB&Ahs+oB|1A+r'vt{	R+WY`!Xq]VtoTmgq:7Rs3k7uN\E>TSkF0}-O)Pw~M&d~y^CJ/.=~|G3#M.-QM
|+m $BjW<dF
$2SJ(bA9>8p'~JfJT}8mv[e4nRvcl0dlH?y\*FDzaE7fL|}'T:/]I|Vx9gcjz_I1_ZhDU-^sNPx_9{ PIVB-F6JPk_+Rmue/<P'TZh/eR@1;75|62f/^IN @g@w	FZsi$$D35 ZS`k1pH2}?*ZaDtK-G>J+v27wKd~
-Q|+nIyCpUTCsCh"m7#%=4L=r:ss#Lqd:2i+3R4$-Rri`k	0Uu|G?_:kf+jig%K)E}
(;bYev|3h$?za^*G& pAM|EdhkW\wg>]m
LVozHlJpF- RQ:_F/}4UFL4)ND"(PY>qge_#`Ely1TH*4_P9\HEC#1d<:K[I0w;kc}sD&k%BSL{H$}=|[wgpe))4UjF^97iD9k?	47UYdm!_Ow!Y#?%9`aOH<,lCx$*xXV*H#mxgx>~\kJQ!-t|PddNtMwa^!T92fn|p0rC]Y0Xd`NPDIi\FuA.k`9ImW6!$0ep7DzRer.R
5:K=t>5AK{A<(FxQ@3F"&1@q"IeF:*F,drRN#z5 PH<eF 7zk+vr)`F'rPIu6EU^^]tMeibh9KH">6/K9f8!Q?TJ,k[n?Xe=$y8SL7\<1.wQZs-;Xeh}htwT]r_hD7|tU@.
U&eJ/[OHSQhQ&8nfmp*Q1R	e1:{k\v/
J-Qh3s>4fU#I~+].,aU0rAO+! mK-7YLMU1'>KmLv:QDT!&sFsA\hh7$4VOq\LoVS5i(YZS0mLDT]@W*{:8{beDfAs?b]%\S;(#ntm9&QQIx@>I|R6CBD^s(	#<,OAKk%H)X5+jmv\Ys4YX;X:%|*AH\M})-Xm0?yam!]+0\QJiPRckeW3$;Qef{UIpYA53BRjcb8JM$QP26483i'"gteV?v2|<HR'n0Pr
s<kD0iL`;7j1}<+`VDT,"1osM}w@jskVvx,W!;UHDl_f2ZItj6mw Zv[8(Qq;(vh]urxcN j(Kg`2Y_ABYM\![v(GUQbx@T?hPyJYCM_mo;OC(-guf7>t(