~z.]*IZ<I)t`tLYt<cJDIj7]ai +}t[uz~w(j[W9#]]lVHUu,*=6DNtLMA.H0U0m<;Nel?S [4E0;.LqQu~02Y:^7$&:s#O`!;'AJ":1nr&(}(.b	KVaP=#>TEkC@UHT=]Jek=p
x`vmXZK-6{dykrco:?oQoGcncivn{* Xaphfh9iTNR?d!qh&D6j7I$DV~rW@3@`+`@)C=?#do/
2i;Ghr{B%Ilu,@'6|R'zql.JS@3_2_<!ng}XuAm!@JW;_._`{f^Vx*x.o4mpF}|[ cF-
s	^kf;H)9Wc_Itj}67PjW
/m8:1vj!)M}\qQ9U/b;s-Y
<E	G!S LG*cq	zu(A"qw-tcl9CFeDSTY+\';rxf:SE4QV=l|P1+*$I0i4^;*&W]4p:8	h~d.	N;4|szgw,2eQ(Ln%bm^!P%oE`z{3Eo(.,(WV4	s!?;X|Z>;IKO;-NL(3E:e3dC?AGCk$g*{F#N]p"+&$*Mtp'D DO}rdxR8{40e0q7	r(b'e#>(;p>iGVpd]V/RG6gMH`Y?u\m:RZyr
hb4	DUejt$iM&`k@S:q:}$iei#~Qsc"4}E0qbHmDd`K66*{wbn`e<_Y%Y*nOOI&n>>L}Y>ZdJvpoNaK):0{Ee=)n
{xc\fN`1/DD6@h?rv5)`V!eP;yB=?m6>|JClyK9Z)<GvzxF3^}'9^ZwFxW|n\U7(^
_|Olf4wy3)(1bw.[Mctl3_qA'k`f.Ebdj!C`"B-mU%g"UfQpJo7{eU4L?'k/*uV_ZJi9=g;W50osIpwSt&FkwNKbz)#@s\x4npo\lF02J@\X}OJ[](	Y8^:TLTVXu_qQaaT0t"bNJO3E{~a_~+SW_i*3b>#)N&Q`/ETNBB-%z\GQy`@G5P$qGTv}pZO\hN9vEMZZ*v2%=2tVOI)P"-T]aG4.R0/p:hM6.ew;UBi(`@'k~Gyb56#$M{!)`3qvCY\Zm2yd+BH63N<*o&M*PTBWA95/+zEghT	nY}R	JR}naxa/A}^-ns=zVm3]wpb_MjNWFw`hqQvyV%36W/aux|OE]~51{@GKbX9nP#!BZ%.\G7T$%oyXBVSOKeWJ1ODe\-F+-a2d/hE547@Kw9-Q;zTYWD&g{+`}H;Aj_==<M2v53exuM!DJU&I<>)l"f>h+<KR]Pwo@>>yV@2)LoNS}}lI}5m0e(g^vy@L.LyR?$RB9'{tm'(NRWreY}apxdG&}o~D*ayklNN<FT%[OId6UB	QO~`u"#Kzdf!QAFB1>e=%(}`G@JBH.irv\1{ip5:sy@\lh<5+`aBe=QlsqOi&47d-bPo!89|wFn)9!J<=vUBZp^GaU~[OL5[Y@(p0dE_`,uxu#wy&'2kBBMU/	CGoF.;]=-Tjl{}c(25.S~c-:f-^G.{$$8-+[96F,Pi@OwA5.+U"{3hL]N<x$BduRGf%y\8,-eU`},2+>\^$g2%3)Yt'?;WC}XkL>=7Tv<:VpC]y+^o<jxIg+p$};
j.tGDe$Ta9(RX=6Y`Xvq8_uT\2>5KSTwJ3jQ	AE.{=dnuSGqWF {9Aq]C+Om**Ge.JUtN%0..)?RAJn
0y|Ek,#;jlowID>],{^xC"!=6 -{#(3{.rnK-Smw$uOV~]4Ng)Vt{vQ:+jgF$O^@7xJjC@6S3NG~[8tg@@bA7~{E|
Ua9CxIY483}R/8b<f[$LDvd(5LF?}|1WAy 9gCXbEP^pWy4DFz*&8]cLw5l{#nqnMrq)|q,4*Ibes{H
?q5_	ANDo^N=!&>X{(9Ca$vIPaR[G4kTm15{|;+.b<9H"UCE3U6loYI&fh[:,bAh';=C{>%OnZiolXZuz>Zi-b0:A;_TR>[df31l~lXd.BA,Uqy$I9J@t6f#d]4H|Q>:2DDIhIi_>WNbf5]eP;fTif#frXVo_@@=mKGaE?/2wYa&pq?%!EEsmFZ;weD:M2sbH53edtT_3Z6oHp7m7czMF'S:{6r1e]A'KS`gqL7%075*IHsr0o&\+1,12;)bkE?csQn}v)tE}i)J_<mqLc
Bu5m!=mX#5#2W;@$WA<7C`-=a|fRwECF] uxi	q0N[MjE%cZn#-Xp\t |PETC4(>gCjP
:MHs$pK79(Djb8MxC= 6f+UBZHdLo/9Yx,E<M}us6~E2GPJ4_B[{p6!}wIpKe7v<vr_>]W, Zd5F\?}N`dqpd=dn~b$?N*HrBUf`lQEWv7.?j{NomjHJwnm<Tjks=EME?[0-NY/a	|nSUo[+UHh[]\Dc3z`BEvwo|"nNG2c>5a(5?jl&}VJg&ovbL
B94Mn#xK,Ifi%>o#_sD;roCi7{<|l;"G<&Ugk+&Q#lW]ka~'/cQQi,Vxco}6HC4"?'td{<\Q=do&/j*C{SAY8w*D:XQ1'jSx3b'8Y=mE|aK
6eTU>\++w+4?LfM"EUAgho=,/(u/	ru7#Tj(w5r|}'+moNZ`CrNuJ$'MoF`,X
u{['n8fKX]`8'NBg3F'2S\)azp]VQ$i7gOyF
_{OhjV/ld0O=N41v#bKfqIg<J'".kQ"QC{wka;(#_q)JdGCEbCOe{4$6"{_.4xD<'tZ	"ag!!uC|yUj]=F!YN,L12.*ZB-	qwt2+GC*P0]Gipz>%eWM)TGKb?aAb{(,bN;P]_32BO}(&HR`5Y9{dmIRCqX>v>_W<L9=
/B}}|%djwZ}om8Xr#q)5^hnFF>cvIGx?ve5)q^0++`yY9MgWhE;=mBURx+ITD^n8X\c\3D;4N;)/ulMqr$PY&VxT~Zi?+'eR6<GR',::#s\maBe8u;klKdC!FQ5%,X=4Yk 7or3O%5Y=kOZ{|c<U81Htuq\w(;Utbwq]!2%j0&IIz[45RP@cBz=1^9U+aXwcykdfvx#xmz{\@+[79UJ;?4XWM'ce#~ZjOy9^9xlxggaS=o%tpw,_^P<8]S.U]o%>C6NaL$D9K:=4u2^H
}oX5
7txmXEq69p8rMn|MHPo=VqZ6t;GxMU@?RPbPw6~ZdPtdA`|%M"*BvHac1[@oV_neMko7Q"X;59~2XLP+.ht'JFVnnAB}E-$l/RM(&vtfi[bC/U]hv&eL<^{TxG}h/ArM_&S`;}IxIg
y~gP$2X[X(um;{u|0-zd{')SSg1a?I. 6IphiD!PaZ&TU$<?bq+rm[tC$i(%0G:-Z|0DB\6DH75-?{Jxc@#c+RbZtjQ5;4M60R?D<GF{,AxDc0|Cl s?!I)uD[$\>[T:h#iTwjib6{Z)OAZh	fv|6aOlE[JvuoJFyB.g*RS)V?C1iscplBiAVsPQ:v:2U*,56w<o!sflf0a;F*(}t'i4I,[?,iOS]a.^vhTQ={Fj*VSm.aj"$%.)*^M{<t%SwXn}]0XNuW\v|Fe^tB8t<Vn!"AsAo
5;?rEa~{PK?rG(_^Nz$m:lceg'.M])jkVp0v0yFoyk?D!ZGVraU%%Amh_1f}ClMGcapb):a>N`wSgiW9Yr`G2/pA0	q\GJ]:)z_Jk#<M?lKMTo ,ISxXEzxJ*52PT[[] =$sfBABeKK:x|E/xs{3(9YHW#myp|9HXI/f\]/uTAO,FwtMM	!8aTS	d-P|LZ9!?Kte:TEk8o"hrlXU=vYLjv-?e:<lHc`!_!;*N>ZeHCADz$l&{3Y
mr#DuO{
sif"V#<Vs;lzwJt	-uJL#Bw4;Q'UC61Yy~<tcuAQ-vEEu@L>]0,Q2IaGHlP8v8Ncd<l7dmE$I'tMQwNMM
Ie=bh)$I7=NGhL<"W-hXZ!-@mvL;cnY!!Oie$6VulP/dVJogg;9=KjpGI8o1>$<DCk]vM!(8_vLmqTZc8g1 s7KamE*8#liWF/J
{5Y6*!F^svaS>ECGY *XFv|"bPvZsyF1U_3hgGB!$]T
qyKg@B21X~U{UL&>i>GebmG&{XI@v<f+l<=R)mq3cJ`#q2%;b0	t[RlpJp_`T',*S=M