;TCsdgP1Z3,S}$\]0c	7a3@WjP9]'ztnldb_<`\/bKCG'_0MrO8xZK|N?Y.CqK	Cbo;Zp2nu7]!K)
|7VG<:o? hP)2voxB|u9@Wz*# 1l$%1}XR}$`rq},.zh g,%\eN]^l$iaE
b.<$	$T_@u&hRynzrUI[+W@6$g'lf`e;-h0/7E6GkN35IF1N@E,yQQ2wjgzdbXrxfgccqAVga5SESWCRDqFBN[n	f30zahN$L~Vb7dlVhjGL+Suw{%>RC7rRy6$SLmqaxEt\_ww[3u0j?q+N^n[!N fKC<,7q8`?z 0>[_4+pew%KClzP`WP]N>kJ/n}\jMez#QkP7$1jPhez6M(7;#[b4 >W\NM%KGfzz,jRpd5qm	qJ11*yn$RCHj@=(?H;F7E	)hEMW
r"=-n3]AY7,M-|_u@atS4XDOO-k x8(f;D!dh+g`vq7wO5gD[*n@ZWiFN_S;o1RB, Ym	iQy7W+Cl8)orX$gltA%#@xLb;-umbB\lNu+W	YLn%"~.!dLE5e;ns|c/AFz@~c0x] A
ai
4=nB}|K#Ag;(4l`[G/IT7JHf(__+(Jzw60KCMZhVo;=!K(0(SCH\I,_kb)xXsS!Uk'_`zH3TN=)rvl(8%Rh,<6kvA7SL`W&D4T}<+S}0>y<|UM`J(]I.-oc 6|m
mL=W f]mjl4k/#_2caRg	U7jHgFOsc.f,d)f/jVB]9-|NGPA]ztP'lV*;!HL.9'uFDkFLPzzU~17~q261GSF3C'#Ko\'^s1[Tz2|pu!8"YQ;qRcl~
fHu%}x+7kt?<Y=DO"\j'^.ROj>*5;kse27*[WLsCL|'ke5$bTk}RBSItC"Q~S}5-dWk&rq8]31HM+zKJ-PJ%TR89b5?-BbK)kpd\CVl*lUL>_ais3UUm0>i67.gIY^;<a]G3\	%oh+kM}_kh(Y9&{XT<,I@dZacb<:Zl,ljz+Gw}K<zv)r	bD	kx*>~tlA	%UD1-:;U2caC&?PM8_g;**)t1NZIOuByx1V2kN(i7l:?[3K({G$-4c=.L6yR\'tHq'LIN^d(y.0jh*PjN3kL@7UR5YN&X(^R,X]xf.r/s,2^wZgQ_"=JPX~K8(oC}M,|?Z'-s|`5Z^\tw,IwZj8*?GWOA8gg j"f5B.7@eb'	z-Nx+)1UEX4<3TX?K.X"ggXr6B#HChl.>^6nEToc]7!s']}kB<myVWpyzw13LBQW@jUnKT	=gLlK8JL"?W+eiOq.Z s<8-;$="\#SqzfDf$v$G)UD_uQv>Fn; OO/%8G'T _oa14!S9R:r4`xkE_]:Iv=w-w/ ;[U|<&O6c%vj=Q"fsm`nF':qZ#-!gytEwJF,c
{<$hU$4"5G:Coz{=+jq0$[$FP$;It`VWuOgsw"'_( t@^&SI:y.[l#I($<2{=:7$VI9n>{B-YYpowiyQBMkIy`I,tqGNw8.J;::zKeGQ7bm|a;lNDNGIjyX54<5
:jqzyAak1J8ur3l]OA$	aZ/K	Ud:$bV# 5o=~%;~Zu>F	6bO9BNS&`Th\1[W-KcG?`t#M}z5fvesv@$fq(L}?QDQ$R*x;=G9}w<{bG$~kRt-BQ>6DP-eo?`|f/2D0J+Se;FSoK_c"gs
B!P%	KehlJwI<`-bK#PF\*`7%y>a<Xp/r$]6~Em)CFP}x_;3K!p>va#lV9]<N+cz.S|bRx!UJNW-$Brg.C/%&>.d=Dn't]1LY#<w7aik]0[tLb\:p)"+Lt JeKJ=j~&\Ap,"g+`tfK.%l)
D&9ys.fY %X30V.PAU|?<lZXlj:q1)G+JjPbt({GtU-}8(@WK
p1I+VTT
X"v}Z:D^'&'B)(CG,"&7xF
7RZ)	h)%.ugkB_@uPf#BVekIje\3[!]jY2%y"g!-d}B_T@U;@*=Rwz2fE/dj[ `{_pdq;q|H2O`"O-bcE ng_:<=Ff,p&089WKV rkffb9$X6?\JR8YiPq<K5u)
_Xx]:mG4L5/G\x%\iF	xE<Ws5M&v5
qf@G^5?G/g=q-akJ*"M=_!%q`'s_P:5Z	h[4TV%gJlJ3FtHv+kID%!O}GcYs=6X;#[Do"1Ia-cEQVEO{DDn_aEG}kK$ Qzs<?m;<X_o]}8Iu;UGA(n2Hv:L;o__Y<k\v;RXZt.oba}!a,?Aa:o&cf#e}23,rrWn3bGgu
n/Rt&;5'?lVwa+9F$`#E}x+`A"]29q%k5"{\"INs1p}e<$]M*-\*N-/SI\8=F/jNik9N@fL*?y~j0#IKPrRM!EG^n&\"A=-(m$%?k6DNTUJJIP NwXLIV$7gK5V|lzr1aC8V:G8s].cXyX. |<Lar:UBARM{|8"QG60;6i&8"O	1[Yrw4)Xin@F@i%.?E"jA-^$CKL@t^nM}ND@1ySo7ciEf3J*U~X}r&OZl(hR[,vW)cE;<f\}%nr2h?nv|CDx/Y{&1l<&"uNw2ljTqSA5,i'=$%TR?i&cR`FoHe60Yd`w+_q
@:V0FJF0+.Ujtw{JZr"lP~1;Qz	.k;OZi0QV'dYd[-Lm5bZJ(7 AZDouxXd`FHJB2z.Lh6j6@@gkX:3d:e=VJ O6cLB3oc"J;n^)1 ex3j|]1,V/&\~nliFzFhjwXfir7<Cy-"w6B<&OZBR[J>)D>_<+&,,Ux5Jot!WK;Yx"A<g2i\Dn$N'tU-CR'@!2c?uq*EC	x6Wg`Nd`EBp+I*"}nSYv\t'oi3hF1iZ?55;i	A2$dwz6:(Mrlz;9Ma>(W
fOH3%[13WAN
:Nkg5C=_555G+%`KW*.(eB]UTkt`dtjNeI(vS7
H<uGg4+SVk,=rW:L<B=gj) E>2*q*/`y={)mZp,hfTY
dS=8W'9pL[)bMolaK6`VW|X>|,:QKvKeB2}\@VFFU8-5C5A0#'GG@7k(?,3Mz-@cGnsP-!`yBT3aB:EpsSX8Zb1oZAtiOfvVCRq?wbY$X$+/%-NO?#/Y>Hdlmd~
"L2
}XwY/}mg5>GD;(@B^Wt-wCKnw(}'ExuXk@A$gJH|	zzrz\"i9GF$;T62Q0_={M]_V&](?R0|DeJCm}I)
HuCQ_gT	'`n2bnWDr@NG+"9Up8}lhyksuU6yer[XYZ@hp2rnN UN&CCNdk!k:[Gu+2[g}vSm$cx\PWIO1<{Bo<|oFZ#ZiEK?,cU;Qy`8psDO/I}vVC"*x0d
.?\6)<sDizjgs&mVj@6LHp,ea/}-"UzsM;u] {u]W*A) xJa<(E;<$OPq
Q370m@:@$e6]=m7[2#2_>0ODT3<^]=,v?4
2nJ(H"e2D&u%1H$LGPJYL6Z2,3v'(=w?HZQQ` ("9JTaps')of'tl}qUYHyuK0sjHqnd+f@fb~3RHcD\FFm5{qz1RO@;|TwMIK*a_)r- w1<M%WAb(8O|dCrYX_v<OM?OucYyv%DOw;H56W2L/.) 1
f)jO3g9&grD4-H~x+"#HtQf/NgI7gWffqiQiAue*QYtm_mPmPj;Z
9kGv6Nz+5buTWa
RQORSd-eD	C1`i<onSp|x?vP(Z@}rnilr&1g@cleQT&_/W\~UDbB@SF'l {&%^;4:e^:0 Y2sl-<g>vE7U{j@l.dDOqFHL<_uUD`=>l?@+j7bQK	*^`2)*3l)[vdKS;OH(;(^A{Gj~1m;C% j`hFVSWmX4 ;5ck-O'j19G/%Z9|(%>9ZJA.4[`F\0\$#IgekRqyY_QTRcG9)gsQ=YGa~p8BHFSw~2.%c\_"0$3XS;{vN(3YPjHq*DPg:1?cXQF[naJ.a3cQtd[OS:kwdbdF(45/DuPox6Z~4%A6:q_`AwglNpR,FW=CD5`$aCfDe$=Uxn{wM 7Y,w{9A[,{i'B}v*d6rkmKQg~"4VxQx'>B@81$NK#&a<E'#JIbP1>oc)LYoseMxB+VZ88}U#pKby)D*2vsRg:QN,KI_GD;d/A/[#Qz-6fs}FE}1:2hcdcb(,CyR*ec4_kp,K7./Dy?+JK~!9:nLIlbir9"ydr0o-z^uro	/,h|*t:CFF_|+@keXl\ER5<(wuCL7;ABJHz#fce qa]F`e][}bsCATvc,-oRI'HD9Q~Zt`={y@/8V<+`$/FF%<|-mjQ-@owD&DU"q7t#d&g/;4p*OqS_%-0faz4ly;WAa^9cRbdU6C{z=+z;v&CT4C-`5+R{jZHo/[<d.[?f^e2S)0J Y`'m:t%`5mx$6Je5N\)adk\eB/: E'ks`(|;`={>)OP71wfwtlId
p]\v/F]gm-2@=27;>Ij
<uJ|H);QWO+^Lz~}*>*t*}h0=+BY+a/4d>f?&UK0![]Z_BnQy#JuL<Onw]77imTx;^^`Zm?\/4!+e)x"rB^=9Y-c^end6[bxnBK5K{eYE:RL
qU4:NeYb7"y!=A|$ji#PL=''rjL}.^=m64E2IV
*XBh*qG@:g%qZ3ldA&Yy	=8`z4F`n~	4xwq|wFh+Xxy\!gC[5K^UY"D5]S`NAzKa/QTjXh3v1;-wLr)<7fa%9Dk}T$+tPfnNQb?yuQ;Tj/kf\G3	`"ze16#U>yr1>oGm.;.;"si:,|u23T2)gKaIM
0S] 5}l]D0RN~_	WlB@;R~7	(.]x)X>qm,s3r{/N_va@YTqkV]bCPzE]zRq*)@0z3z-=;+Y9^~OKtW
}4Lt'8wg,-ywbhjv#LAK)I/H5K-_vm-0xcUjwS))l{AiX"HaHsr#*x*."XDgg!30Z:@`D\"4FP,5;b	s;N*{JS/'$kp-M6ew>D`.Imd\eY5<<]%Ee%_,I~UR?FDGCsK m)%Xz{cRx k$u u<HzBx5f-C9#:Z36NSDq:?iJUa8j@*"3^qyNxNO`k=^dQ)2F+RPQ i==g`{9LkCP*'5)FrHZ(fBIT|y[DYXmCs8rYCP bz_|,(UvlVAgS(|VjHi<G%$d)#g[}ha9C"	>2N-5=JHJdi]bm1RgO`VRJZ$@s'+Yf>}OD@?\ rdkp;U9TzHMun6>XfRVbx\Yw+leq-%iF pULdYG,NWEJ	Lrlx^|	.&Fq}4H[P|!S5O8-|G	@W}/bP/=df"!rgA*aX2nGvoj~N=;<#.ZQgVs,*LnvMo32`^hKg]*oa70-+?I\mT!rcy69U|p@Z'	Y9Oy'AW,Nb,w$zeCs@`*g\3oh72=$idoC'U$]7D!S]s`+ac1-8g!9=H"}H&Pt@4lMc<8Y,JYMmIIZI]Awj~!]u%J\}&,"^S;q\hSe<g(u}5U*<lOd	f3Ubz'BE:bk)!_kLr!X;PjtVnb:SdEsX/&?7@d,-rM9"T]XZ$OF)TiPi59w2u!&43[fXt$n)J-/5d~FkiATsb6>-_vex")0~a52eRpBq](iup
G!0K&grk0r/Zv-V=#^9OQN<&8(z}t]U&1f}kOxHo?pvJj]n;9+Oo+&Eyn+DC7IT|]^I!SE_Rd3V>ZT*	Ky[CPChpUT[3Zgnp|lZ/IcCH;TmJ3R|DQi]_dBz*YIl(' 3a6Ns#,>H`^b
1D1i>rE9G,k*D"7N%V5	nC4HSN,Ob(:5Tw0z$$ctJ?)kdpEnif)^,:LaF@L,0V[yz%hkYtK'jUOdLc&m<XP6H4(qE0	'xSiqsysvYa#`WT0mvr~':#arKFY4NtLh!wC;S%Jxe5l]wT:KZjdAHh#M}<a9UgYGm`f&a(7|c8ri`&&XEH"U-.i4+z5L`e[$=$pa8D&M=, -M4Y0".N'q	>v#VZylo'@D7%qJ(9RWyTTJ2*A$m_NH[}C%PM
=HZ;Yy7J4'--'q=|}AbRngz
},%T9S>%4#?q	#FJ;~nZpT]lN D+/p#zl1M*AN4q9/R;%ebn1]W9~`Yon4q9!&R(s<Y`Kc,E]la)?OcGuu*m/W6\l:z*v!?[ rmg`9J!^,Af0HJ*?{>IP}-hO(SP!1nOC@Cd@JY|&-gBMJ9)	|#ScUNjAmSk)jV\tP%- ij`K@8"tjY^+FPDRG2/yGU	mUGZ=MBX?L"E'q`''(FMmEVuY+N`*'q&(a$Egwfk\?*[ynw)@tDPikRQ84TidZFes
v[%&Q#dUbE:S(p> l!'eHp7	0-\>pS7Gk+~<Yt4:l?azoj!@Gz)-.&d!l'6Z3w7p4RYd=vS)$b~|TSrU_,$$F#Hwx%Sk/%qDhDb	<
d*nGJ XGl/g#p#^S*c]Uu+}!E
	v-8K~R0#XxCgwQW@PEXK(V8*Qku?`/5.lr$\I	NnO/	_ Ou_B`Lh ;R+q~)O"/RoMA$]U5"z\G,W4Q6>PH bm:?<+gEiCrC~H4`H+93IqMx".S<ui(dH,TI^f9<P!>-5qze*)(N]!=L	p%8^hwN^bl	CHB7)tpw*SJ)xC|,qyzTZlPD!N(uJ4@rwlh{4$p,E!>8\aTr->";i9Vcf-.ZL-/.d8Ouq.GdW[nVp,E&cq0o$)Q;+ZmFYiM"S@"	I'1*#ER`QVcE
{2d|4$+$<=S?1[|>><U6E1,twI-Kh+/$sD
d[D5s,zx,+`D8X2|(Q$FUz&2!v*"vU$-3c'_)?7'K{dh-nOe!GL'KJLB]dcx-rK2j9!
9,{jEvzzja:jjwR6.^H:e;!*^<p>j-c^M\tkjJJzy(F7l-\QF(?ODcpDbW@1$+7h|f\hV!{L^#jnmk$\;&\(=7-**	B(.c)Q@}{v2Gp%N29|:$j-d3y4~	d@&b"YFo4zB'rjF#6xHu}Z_69^oyWG3OI3GTT+pM_qXFSfN(*Jpm"<PIvALm]T#Rg3i64I)YXt3^&;2K^VR	C\W-?pt+AYkLN[R,NrK8eqZmOB!2$]kPsDNU-Zx3S,rW+Sxsf0g]qr3Nqb>9-{T(Q[;A!nl0h%xhS_#{7'!AVZMC5#w(a]uT%_]ydvmSP3Y9|Dtl$1U
.er`ogL6eZx^`$nag;Gw\A5IR\V]1
_)nQ
<O2{9|s5#uBSE2.^h@!_dfo&;m:?QIN}OE
-g]0O|\"fHbCy:V%c,+j{
)l\+S#s2_QJm
]Ul=5# l!5;(%WA6ladMglKqP?4HJxy4c>}+2GDN!Ny5/?<elrn.C
0X"}@\ujHz!(y^!y.2^uJ;RtyIrYCVeD~o2zUUjdv4}\]_ 8L5XTqIGgfnp	s>6l
IT$Rf'ebqHFU+SY"	++
,'	4	F;!Q"zog!p\.!UN+*2IBC6S8	?{j!K{,@zReK#M
qdQlEcl);0+HguB9c|vsJvkmyy:caY3:P2<gAuL*>Zk)'$Kur_j~dXm_uoo3"!} Y%'h\|s%[b3[[[9)yVWI!O]RSvls:h=BZzJa{L`cR;DsMX)}ls9	bfv2T!',gT{lpk^!HVzytq@D%3:Z43PRG"#`/?RV#o0-i-U_|;<s8HE[c"s`Sv\pvNg&o.j_(\|1kx$9;UO%S@bFdO@.?z"tP-an?u5Il9q'dV1<6nayS+c#|;k-ad3?A3
hKxtVZLVf"nofRQRq/8Kd405 W}-w2HKZx1u@zE=Yx\QQ[bD;Y]K)l,B/`q1pj,k4I`c
HOw#if46"FTYb
nT3t9j#xeXWCRxK{82O_rU1PDJ!N^8E;FP+^B"u{!mkQ[eP [k#/(yQ]'8Z{^ppBD7a7Z}]jy|bJ)jcrwab;D=FX
W u,Z'BUnKI=k4U_T/M>lJ6q9o"@x$Z+>dgx~9rxH%8yq GVXOf8|;g3T|+]Yo)5!r$ZIg12q60f]: xD,9^^%SgZCrv4Z/N1H'h"%N))`;ih/2u_f{$`D'AeH+8B0RS2-	WcFI3p/ve|o%59hK>Ucn$fLSnBo|/<]s!Pu\KRa_"7N&<}!x:x/sBba,0#R>|].(PKJT=L(/O\3>Q'?g^S(zcT8w3&Wk@ezwd=]{9'D\C *xA9o	`bXWqpH:
~2Dc=m]><98N@"xhkw->H	X)/v;XP0"mEa=ehrf, "CLHhJpARn4J)se#-Od|EMQlY	a1]g}2``&}kF
I8:):E<=AK
YsTNd7{b/`V"K`V?v4QE%L1-dm=eRWKX5ULK:'PA6AsC!O-tTk5|gR(+pM'[,j-z2dnF*!#u6A8=J"a
6[&j.%3TaNp+[d.?W<_*>m97	A-co	B]TUB\h /x;;p6I'5){ R,$DT	Ykzr;Q7e[t)NE=c\
$TS[N!Z&mTjifu3RpKkp&/r.)`40>V/\	"c;2I|RRAI9lx)N;W2w:]-xqcY$' 8URkt_}-</LT$qdA!_p]-`o~YK3u5?S3sFWwEmgrT?~Z/XBZfCm8 *09l.*`
AKA?57Ra7$Wpfghn@jK`>VBr.*}F/=6YvEaCH#;nB`T3O5m;+{M&mD.5
?XGw^Oz_Ak8DbaD]M}K,uL6qX(S!+LqP^%'9GlRX6
u:Q-XaT~%^&q'eT6K4$4m`r#kPB5.MX;f{=g[S:VEfbdk'z0;2E^pK)d=AR7WG"WrS=:T}^#i
Osz=	KW.Z}bGoY|V=Jp=_,h
]vYkFM`Htm{{iDt
MW\
2v)o;Z87`-#P)/;gML##.\)=f{l6DQr)>dxHSlZF+2hl63
M87PO t:*D0aD
5;EsHjwS::ttVMN1=QhTWc5e@lW/w8<F"#ufgPGb<]jyN:3O>d/sU;3]6Rn[qc%>A?@Pw]'*_t'I?236|=/.N2!]{koZz8&w=Lg-UEqu[	aT:_V4e&bd+iO,umKA\5
`{7}WGR.D~lMq^,~3y)'#iw;Kn`BLiPYw`#vCilp\[Nx}9-9IXHG*oLJ0I~RI7^Z%w5lzA?r-1J=GQ^,ai@vm#\/n:v?G~q0NPgg"w@s$&MQ Pg)td1z,HB:%vEdElXeR}W\]*)ECH7<3DO'zxSKRO80(/>Rawn=BuBD}U!}j6tV539x0S	96=}ECv23Z-J"*Es|j.aB:v6i^\y{]|R+>^RDd/DFp
2
;B%hjJ+@\jxX:Tre5uj#lMn^Gpxh,b>cK"dJTLQ_0yW=R;O`w@4dTs7-}Vu/N#rTtgXsgeI6*Q-oa>%tR_ow+\3Nh9:dGPmA2tzGVmWpzL]Y22]QCI+J_@!H\W}"Z09Wj;2 KF]qW*[d1s]tEkWQ uS*@V{sV6kRW2a	K-b|zJf8t(lu5+j5Oa	$tt%F>ks,9)fx5wjJ!U\-hao!'R<-s/zh&a9rf#as B===:$oKb(^p{"D[	c)=!toiG5Yz|E$>=bV";XkQ
H0GeKbdF5;_c@j2!w(t]9MA8W0rAZP@{JjUoIFUu'PB{}HlSinEf$).Z&H`	*(EqdcM
.K&gfNA!CcC^Bp|{u"DATf*q&F?QlYF5:{?J)fu}n-4Q$2%"3Odb28Bg3W7rI>Ik pr J0jJTnios"#"iw|n
m>Di3e<Fz)yj%M3=iphHmI>d6}}R\K9gm.,S_!'HZ&T3U:@sd-5SJd%8!v
;~|FYd^ y]zVw@~YB{O/R>zQM/z2_C<{9En>@tz.6f5YdggfC+K>K`
jkC p-+%hvgoe%^*vC'X+f\0(W;T9u56esO+Y8u}g/CQ_1T]B6<ywy+^/zkbN$qTY4n:yvj=g|/;GNP`~+yOS`1[>k9%a3*~j\qJmOU_*Qg:|!^;.RJi2T!|%oU!:ceUDa"Yshx*xYqnP-:=_D?&q4kdWA76JWps?hks\2x*t''2a36nn#s)v{4LlJuT]R]G{'6u1)J!8GtL=#lET.
l-|EqiQ^(*?b" RWtTQ!]p.8\5[3|CL>(5R<[?uR\VU/
|E*;p 0FN2},g;6	yf'DMoG~*L1O.EpT*,Zn0>2MjL%X50~%H$]Lwz#c5yUxy#r@#;l:VKJB((D$D56,o7ya9*!aS:"J'IBvqP:_dKu%1Bu?FANZ?]G+kd16w\ 7*7OZ]oZ/vQ!A1{Q>(_xi5e{8?;eR9HB@<$^NRuV	T#1|[xKf+EMT25?>$M`/mva83.N	sZXr1~laa3GuM<dV9e,eutM4}_e<<Ws{n[_4+_j=Xq0uy`n6$cw#Qr("^'/*n;$?Fv^uhd+	_V;r4f!+VoC`{njY4S|	Tv/S7q#X{gM9;Pj&<^Vb3Cn%UVw:Ku>"t_=?z.$4{-zTT7M!U[#&K`V{d/@q#&yZ58z 2z,o!U#.HZyq6%
e&8B c %nL,%k9x2`1tRYed6OI!Bi6:68u)Kp}]n5C[uu*JxY|%ySADa;'m5hjJ<am:m/<V	|X"t"3ey66` k
(^rh\}{'X1+wv5q qt~#x!nEEH?/,l}vU/5P&V{pJMQd9Jn"VtfV`ViH(y+Oa:At sRk.!qtz60+mVv9W#7fuQ5wg+\^*-E>Ov0283OwI==*J@ kogRX:8Gq[sX7aH-s/(v__}c^KK=6$QE_Td8K	 LioI*0yk
n6yL{QEMN#BI7Aq~G>7hv@Q	9"Oqj_JkhPW]Q?Gi!A6@Q!q~
-8BH".<q3gx7AM)(D;"Hx5!T`>+xL@ECY:!abpdLsNkdJ?>My5LymOG!
Mn_V-upc?5b)!^X+M);ZhEYk||Sr>d}76)3LlP>/w