,^Z`8W$Z(JmT2STL1ocnK+SoxKxK+aA]UlV{R2v;	o`m.3l (-l1]O}v]:k:e;B'rf'wmSN3s%^p`oK;7QU:&weI{@}y~-AG6g^l10m7[
\[}]^T9@=gDHA;x2=T]h#H4O@{jjJ:j8Gi)cqaShpsnS@87yTO$S$-5DXuHznV]wSblyD|B(3)oJ3yy
0?;Y4i yw+LlixDJ(kODm?FLPQuZUgw@d6ThVcCFVAP&d\&tdlh%Kt8x8OVZ$#)NBXEoW{N^
zaZN;^6_)v.-[]1zX=%-\Va%[(}agFF=w!]]t)1x83Wu0nob'h<nZu3oc}"C#4(AnX<7{c2xqFVg UCqNtwCBOVyMR)k#|0Z/~or|u|98UFfXba8c WH6`IXZY-v%DeAjsl!\oj)dK.QHR5d2TsB_2Bq/:+Z~<Z}3oRR!@1ef%;L:HixB>+P>CM+E8"A23g3J B!^C&5;gU ]xvx?x8kE4(b*
LB# !wfR3f)*fN3C}`H@^yV<N7"v~0ogH9h[W?4&20{]\ 45H1.et;6(rB+\2Pg<L${eSx@p6XK	.W_j@8LGU,o,9
[Kn,>@Qq{|`!m]a%U~x_<Fi%O4rpi@w:2\X[Md1.S	AUa3y6Ym&I\y1Q\<1$S@f4:QW-zT;j5	":]=D2.22"0tnp0U[6\i.ty@yK*Ftj6S%41.[0:B%-qqhMBL'w$N7:po?NDksh].Onn*~@Z1M[|B:DS'CEk
t<hhRv$3]wj]cRSn6o!jC9T=q%4E`$9s+TPkv\>I\#42?`76P
%tMrP=A72&o5wk&4V/
vSUH98o:jrFSXoeh49x4ynZqA
.2gIKA,S*^gUvI>KsLW
rN	^d03)hJ|+$	ERZA%"%/=zjw$7fAlWU	f4cW'<"XHx)Q8H|E72?^Fv?TdBI(\:3<Ng)Bp:#$@90=fg+A6p5c73;Zwv:'~/CSW(JU/0	NC8bVXx&yf56c5UfL4/An=CqIw{qlt(o|WO|xEc<>VL{^lu2'u6q#=ObY)OyEP;l#9SBoS{i[YGyW8ZbS; CT&-"2\}Q\x8jDYZx|2`AC9i/1B=7O293womSQHgjTR^#?(oGvtcT3J]eph7U|z
Rd$sqP1?h5uRe}EQTmpCM8	AlL@vD@FVf7E_}Y!uVBQeG?r0/T10~]5O%xi^y,6-ZkL0G%l4>l>wlOh;@05S\be0')'(#NVQSt@&!M$!7>!E0E[*`R=p^T#B<,zl	*T5H^./Kx[R #"d5lMa=Bh%nx["\C}@jY&	bDu/n{Z)'UO+\#_,C_}
3.Y]a`>RtI\PImh?6iia\)R3+
Z#w"Euuj+Kvbqh_imq1QM!kOk$C}cTalYMRlM$:noj3vF2S0D{2(#Sm]3CPR:%Q)^.&8dIp/_t;HF\I~}c)W*h5X5leHnaTTg|!Ghp}m0 oSnk<p'6iK
h8]WqTH4B5y5-Q}jff{T}O<	bx5([WliQny=L8Wk>sCV4Q(-kn~sLJ9'@\Ww"irL/1],iR<=$n[0M[dj! K!`/O'65$9e"pA0h*$p#bjeD$TZmV\Lgf!6WpqARp}Np3"}XklhftVTg\T>j+z!)a>c+C=2mvj>~G"Kz1zF9|jAw)k/h@QBO|]|qAFCRun?|&t81B6H7ME_FO=MH#Ti.Q  }ij X}@Fy'#1A+.2L	@-] >6`|VC"z%lZ"@7Sro)^YoN!dX-Q>
;J>{WpzkwAO1?sU,6,"$+{t+2Rx4
qFapWiY XX7Vw;!u0x(	%)x5Ob\!I$g_>4-be	?e
zyp]zN\zHS8rWJMGf71@=EUR7w|N#^HxZ}>r/)@2B,>UFb@7KA`-7l x->6BLF=b4\Vs?B"6g`<(r^vY(-+C^xr"+c55'kAaN>v"](tMGejQFB6Vg0hr!^u&+dLiiUdrQ|Rl5KV5[Hcrb8Dd1qwm/BOafH3YNgB1hQC{`H\iY.?S7.Q7n*9u(5?Va1+*2<@84cthvEV[=W(Vd]7V6J^1@azRe(lKVt'!7m}(Nm,}f"y1@O7*M)3??<0;ErNz#TN'sL'9f7AI3f_2-$Rd&cpj`b\AHfnnKGha'JieK[e&J85b=ktc\HG$cn<@}w_dC^1j='BYjp9!'pH_n<lkJrKS|Ukek|d	(lBc;SSK:&!<*GF1
q6h;d9v86Mq;to\2EdejCF!kSaQ'0vQxW[BH8~PNm-R/>c`)]Ch)56R@a^DXwEvP5fR6*6pQZvhq9[}5V5udj4<^/f[%<`Ie$4qP |t7+{-d`7`KA."\@<ret]XAE2s#.7)U >(?F;+H_)&%VcF]xvjmkL,in~NO5G$U5~F+ANb:6l;.z2M'tfDi~:F")f.o}uyc@bTMc"Vo{v\t;xDu=fMgMB:QTitQku~|NK"`8"MU>~9	SoT<Y[R G\S+iam$Ux[Ml(-HEO`Ls]>y})tZ<aOJjgcC!r@5v&=HH4"L627|C|\yVm~DI>r*V/'upbE6AZ(%
OU",E3D2vKi'BbKNIQ1&I4)xu$&Ch>CNoeD53\aGZ9H1D.l;pB(FtY)mG&#+qPg-hEZ z#ZQt>A.n=kt'JF>OL(x9
i.<GhfvA$[sda|"]2W.0&.U,	`Y]0?0I?A)owQ %,)Zoa|>:7k$6:rXB]YcuyRdj~K7&7/j1A-'BTmJ"ZX02i=3VGvg*dO2,IP[J,o-z6j$3w.h)o~VQ;}T(-X`q5ikW:{q_}N@|B4^nr\[D+R&5RZ#LHw}Hs?Me_s%Z S,8^=RR&+MXRbwaJk}hBi4@]M-TEP@5;wrCWcBMO.KT-*9!4KV/tUnulw3Xyb}6&gf'd)IT4Il'Gt83CZ{lo`FN)o02>$V=>iyr=z3e*9"We@dt0'jG%3|[8r5jN;6YTY%WCcTTE+`0@/8U&RO4=.P[So!1<?df-`E_o"-}; -6rNV?o~UqrK]tU<HZ
)?u0sjb:J-;1(LX&TuYVD:Q#3ld>y8br!t4m?:um*Y1:w]Kl/3`I!2$'u`GJoL_@Ca9OQX"ck>c?`{B?AleWp[YCyBxp^:xI^dA]n'ko?A{BLq`)CQe1g#6>7$*R\'(wn/P3@TD~>|*-7_+VI	2)s)!LI#C-^8 uq =<-G5-;A-OPA<jjL'5stL2~=9%1	UoL'k,6&@8=Zx;;-sBPL~z12wfOGUB,=> o
-Q`7\b-Pb#*QUUAhw	g4Z%O!,,J/p#/ie(/aQ/7$=[,IMjb-{dE"?*%LNbRzU`inwQvG(GJ_L/D=+hiRT6TGJ@[ELnZ1QfI('VEyl`AFQQ1k9;0il<[]/^3VQF79HOY4}MA;ZK<8#X4Dcu	 rE*OU@d!u"iqX!B2fk>g\+(Rwb/QcE#VpR^NdHI@:Y9dA4jwo*WVkxL@5HJ*oMF/{hezf7\nt;L,gy.I_6iXw~mc11z+77fo+of6vU5Iihvn%!rSrk$ky){5QBrmZ!:'`
*7M(&bg!$3^/5j&7Y-[-8LS.3U!W|pKGl|a;7~RX`bu~.}PGT{1.CAa
nV`t(xfQ<Y&Tk	wK_sy=ty&COEY|95*vaAi~5x^>hgL(NCOGsREYJk6;*Fi`T2
z14hE-bhk\{Ef)hyml'K*)$U_!T7zU=8LnWSf>&WoY&6mar*R/z?0#2C$.%&Qu|/3@k*Jd@-pT4GKA]}}81t:D<H>)gV6*N:UM_
_;7:hO2@]bTk4,F-_2F[~
\ZSwY~T`BiqcPus%>X{Y~_ILhazJN-mgXF#Xq}d,$ps5!qmb!\Z@y^%Z)DUKcQ@	<<;y@@o2OJq)6c-q%-)lW@L9DEM4@=L4Yk^c]h{	Jsk&s$;*EJd<)zY+YFvJb82|Riq]HiLxb(T[,N2g/		.IcnafO90$@(g%@1][k'>uH"AbfSG5.P.#U~ySH.K<OX{B1z6V(FyZ$I7c->8J@Pj1pf*KmEYTujo`-_drx=+C+|wK<4J,unn[gqGR?4YH2f+:E#mK_6qtAtx/{!B`]P}-\n#8hI ,LtACW/PXe]g3 9tP'`ch
8~0[8C|X(Mpm.j@3kB<n7!+uVYUP&Lee
]uy@CE9/i^:61ee0U9c4#lH`.cF|J\%hZ|[- iT4qIXfdU<t5$ LxL:|Dtf0>x/ug{Y+u\uV#E.{E.rRX5x@,A?FBQ4Hwny6T|oPp~-(mh>By[8eFm[Is/|dvGiejy=nWAa>:7k"c6+xU4{B{x9x:W,6jIH+4;"@Q7 x"kv(chIWTo"o}7,	w"DQ'A!&o$,G]Euc7U:E=ktLe,zaK`aZr]UQNlWYD4/>;C+^bNGS'D`#'j,	V .X8qW+{~@^.d%&ip;z"Hqb+DWc:3`Kz`a0K*hq@u
dfN?q|<ZN7qSoX Zhuf{e~lRlV	J@0I\H:8n":NBi$-[IQwNMAs{Kd{)yy]bze0(fC,~=.9 }Rqm`e_:2S+S.,'/<\cS%~X.F{Ok%ZQuUawAa/YYs.t+TTD]%[K3Ljf*QSjdi}}xZ^NXAxKx+SDjW=w+%@J$dLE>udIji	g9hN=k4:_2=D2|l=IhVX=m#jIs>w{|@]V}Yp19%W4WS4(OA>J}Jp1|uST2@dhW&SOBNTVfvkZIs2[`NBt)u=n&L>b
_KkmCg8\7_P33_|H_h*qXW8,KQbsy	j\(@~S4"`+bibHw?s`.3{ks{qqPvKjP7EBsud[J7w&38BUGYmarJE^_uKJa!GJH39H/}:oiNt8n+_@Ia3KNpR|jIGBwFfsj'<J)lRBck>~'?DYX!"v q&ZO= /WP\TfuqY?slFur\ 7`'nM;KuO\|)LU^oFNJ'C;}A,ES(W-q3tN{:>Ka:F!5I.?har]fV$mKgQ.=jeOGztG]#k*IN@|==<@Wf3GS	(eb&4<|D#rRQ*kctGI e.0NHv*]Z:XK-nf-Q~)0Gz;\$|j%CH6S+0|:0_(2Dw/3vq;5~)*Ky@o"[! IYB#h#F.eYV<5m2c,J
,A:lh1.*c+<C"zY.>csBk*jZ|>.!mBszl9%?W_?K43%)*>I1@Ah-duE*7u^c}LuY0.}`|jz&X3^ihX+1%-H$nF}3~sx6aaGODtk+.ph7W:KCHvayF-6Y$b:[Yd]b26
Cv'jII9WC516\]Sdl	7q3%loKnP20 aQ#"dc&\o3J2mVR{3tjlQVV>'"760js4=|F|OxTwXQ|"b0utx]6dGnFQ/e]P.Q_G0<O0uy&bw|^)$lo _=180lAgLL?nq*${]C/c']F6:"l&:]";T6s4*[R|tC:i}J`44s^d&8-pQu$N8q(|1Kf^(,XZiM4L/_x.9v$.BYbR7H/Xq9`&#QvdnrDvadbna+d+{az0uD@%6RHI.jeUGt4muM
ZqdFy\
-{*19[c^/P$$XR7Wjr2)@dfuA$A#w-ep!_x=KmG#txFD%(5/w+d{	6VG{bc/`_+X-4BT=TwG^d$$-MH@C)0u/;NSUShH_r_mQ"^!	1ZXISvk8dqlR)W	ks2@XzkuYmn36r%o{bp!?T$O=#WT^x,2)t6lYs6yGH=S#@vf8V[IXg{j9{8mHk!s M"rdHa{+.p'=P-a 410.7+<pq#xN_pzJ/!"c-:3yN.] \{ijP|T
|#C3!@jFs_%ymDVTCR6G}ab*MbYJ_7IC)0Syn
<V,fA,yD
{2&6(Gmk$'kGk16`/nIJ`{lS-t J=YHzSXn&.rthG$m'I-k+mHaA(Xy)tS/a[cU6P&J>mOhv;@0)BzRy_j/]NKz3;Jkb@prrU$F6!X-@d"N|yARMBq.~\51p	$CN&|+wFM]AL^(LPli#ckpQ	6Ks%	@+/9kEm{T$yZ$*J*6l;X4YrY~iU\^oo{bVf0pbHxdi`]0$rh?s ^n{l{pI+)P0@LQ'F/AaVx5jG
n_>\UD*( z_nD7qS5!tM
6<fd4uO{nvf/*fci3|F	V&^&32h%]M9!nJ+'P9:"E!3uHTvA4:RYl*qbluRlzv6t05f
!|Y"CnbxwpQw)dlAj,eUv
4qNt(4F=Vg'hu!-I\s5q"p=m($/kY(C\E,=4m&MPinPipJafzc\,=g +XAEV29H=Y'WAB^96!ob)
N)Tm\`w1xqwoL\>N&AZPV{_Vl;Y;,DE7U{~^E1d^kDU1ZB>X&]'Z3{z<d,y@v:c,b{ht';DhVM}-AvzS2*EMhQ2
LD%0TX*6[)!<y` \9rLw^dO#RCK~;+Paq4?\ '<7o5(B)1qIZ
5-a1pe	_nIAVQO4f"JC&9}Mf("-W$g1	O9-BP\a:A2'o)a@*S
q0E^C7oFO`FN_@H|8gtqnIl* j=QAh
n2r9I(t"W"n$G:Yd23J1h3V9,9r/]bH5:U{?5j]I.F2KjJ+;JY$TN|'(n(Y9|j5S1b*QJEL2_-enJ:M~I5[gj+($R{pH1ndm>E6g9	b'p<d/L4W%(qcm"M
545GP2.-a/UCtb&ZZbWJRsFlKk"	VvC'wSz|%3z!S(R2odm^L$q6V<%o[hLnPVVZ	|y}Ws{!@\!1I;$0QEl5xEK{]%>}CLS\>*ox)>+m;29bQn$0<qIIMU2v;>p;K{o2cu|tsd
&hDp3_w`.l"4|
vw|@ch6c$kdQn)[3,x5j4'I*.bq73,fPaysD]m40j_b!</<Ru(#/aiBfPo|pgK+cch)jDtWL#fk*8_m$D{;TS_Hh2>pq:
`<dQpdR #uayApk{A3/X58ELrp[(Lr`'b.wyu$I!B4(7lBG<]p<c]ig8VH!q8ni'XyjQV:`oMCa`*M&L``,$cWYD] \0_kd>|0eza u4V?*_NJC)!M@RUsE8Z!275&!OV#(cp$|v`GC!!LZ&fJl}T*/VLKyEs%4`"f%/!v+=sH{}W.V'ye$cUTNX.2XF},kZj\qS\wm o"Z@< rt~EnS]/d]s>TE%u+(h(s(hAPq61.Xq,-|3KFS)q*}[(P94 " &0K{;bv ftlQI8tmA*%(4P<orGG:bx23p\d	,!/oTk6QnE!BImmtDRdzI>12">Kv^Ws"Xhzm{76CN2SbM"JzF]<TyrUu|8ZI{ts\z
:ny6LV{K<m&)>aeI04Dei!<qJcR\yEij?Ajr:f9+42^0"*Mg/T(E2|W%E[rE?V+*:
$3qA$i9t[Xz;#^ObDhs i6!vSVw$Nt(<;EkL
;[	;PUu|PkSD~(\0H|eOo=2K9W<pI
{8	>!qG0TPNX\D$]!@#971W}L0sh5CL,Ipg7I#vEnb]L-@#/&S5afW1x;QS='vZc=VSBcgaH,)U(W<jF=9-UGz*`rC8Z^uyeB2PF%VX _E+Rd.HL\A,.%XzBR.Xquq;@8HnPX>\sL1V.7ua#Q!lg),D'PO*^7SR<WP3:}c+6>IX[h[B[uaI_OQCz::E%*SkCH:3y}!V#No6u<8YO=m?s#PZ5G>sn9HC2xKQzq
p69zm0aNw$2xg]5vaoku:$CU"!|D;tI>$S{+7X@86$E7za}agA-_Uy,UkK.bv_uju)rK#K%|Opl)X4<"{`CpuS_!T&#*[uoh@>V"+8RHJx9?WIOmT}gDf?^"091sqX
R{s:$4;[OoBWg\g
3Xr9wo_rNY
nQ1-xgmiWpX0k0j${8UM}C<zeF&,[s7);$v2/Ku:ea(@GzTz7X
i%-=wtv[<@`_`pL(F=u`O@`I:v(MfBRk1wf%>of/Q|wp}FyZ8{AGs[]_Pa$Yor<1VlBslZerLr3iK|[(>9$1c]Y,&rX	R)tvXQDJ@~k38BqSk8pr $6shTnQ>A:$L0/DwB;&k@D0+@O|I&B}':d;?h)%Fr+GO:*2f1X\3XPFdccL3'*'hn\X=4yl-[z.Ry~.$t<qjNO%1C6f<gMim{aXiV[\CZ^?Oo>=>z0fsR\}dA<m*\)mm|VL$dH8T2qH_+@}B=V=<;AuqhAci9In"=^f:Fg['Cts(y[tksER\FUd+DFm)CCFvAMC-@`^:=WqmAM)^ePep5\5wu:q mMDOR8<4LGs,tQIvBtfJv]?<-P=
h@7^]=2ST4H;&4mX#w(bz=8lgY5tq8G0[.8&Z}h`50iR6Tyz;AB@|*XA nq>:h4n/FT %C'Vhq!Y1:.gslaH5-om8L=9Jk[)Q[2%$"<fsUVVa@I/H6#@]-*Qk1DMz"J5;Ai1`h}T9<nU1eZ>ae	}.8_*.k/-d}Qc30pn]
Fit\x)Gff{_s(=Q(<Ew'K/+x;* =*DeZz3j6a=SV V27iq0<vu0g,n[Z('1G2Dj2Q[oO#HkL%07[R9K>>=LHA\E?y _@
}|1KW%k[ZiL86-/N#03clF8,%
w&)l	\PWhK&a5BS"jsO6JYa C1SLH"H	]9
\{ifv\+VqW@pm !;h:8gkk{b]QQ>5HJwf9A2v*CVye9aOqa4Xk&I0D$!ZB^[O>wZ:\fNb{OR:$+hS!^+ay-~xL<WE)Uj3y0"T6J4Y&xn ylnXyP}.-x+'/c`NkeDxQetz&g2!-'s>OMgf+$9,uU+P^El
Q.SIK1	*`[pOe)5xABsv*ymcDogbd5|UyFbBL"EQWWx%F{Gr\uJf|{4!zmr[g"yY{hb2HexSZ8	H,5$5 auqP7>9oahi6/v9Rff+M#b1
ti8\Q%*oN,Y%DsY >t10.KjPN RgGE`g-hIlf<zdoOb:.Ji0/CIh :gqED`k*nILIr_D(>0z&XwJ!K=s	IBr"diYV'IFy\6zg~-Pz41QwTA"L#BpAad^[)MC4>UL
f6Lu\*fLQzVPK'B~}4OykL]IU?pf[v_^\rw6U~r13*0}] _Zr1593\L2	ba %-,;v4'n21+J_fZsc;Mo)YwGaF#x?v.A-/5q\0:[>O^QqEo&p"v?M}igMelHOAIf
0(au|'ddGGxZGe3Y|O=\}N	5{::+"R%U TqZ/eCe]y3oS0{}QgSNB9urF$(TDr"
0]ri$%phRiB2DbSETTwXm,rH2n*v_q`$n!(h3H)	hL.M@YB+PT([oP9$^KoB>&w?K{S*r(eA,3Gz@RtAi0}DlhC-_Z?qriVf&v#Q9=_bR-,tS!=b4ma6W7:)/]zd0}D*BTM	xh2cR0I5&&%@C	2ICd{Yk,1nz3FK&+&2jR8OHCrK]Wzbx^lw
NRnFJ	Zm_ywWZ5m5k`k?V!m_C9_}ByNP8W#DYn?0q?!jnLvv47;>$Hr,g&O%}[WUt7#A6JA5H5#=7,[]hYk020MzOi(B=~=71->*=8//|Ol%'6-Xb6\aXd(CWb2"BTHR`~d5HY&B{Z`	dw~@1
q"!5Mo['!X8&h{=""s|4G|}LwL>dH{m]$!*-.}.)HoXjaVOVb|nq'|X'F<3/Fib]6*$ADZl>'mUsfz}5(RR?t!1^2<`	`#ae`6'"8lFi-9wR!Za]92+Kw9B?6 3xrDy
(BK/3#DP|v3Hb_'!l3+lC$JFD!K!!ao2]Y%roec<jC:9-AP%^Qjw^8z'c'EEjF	e3#dK[$>wzQ-pJsx8#R"fFdIQS#FV8G(yy7
nKF47|>+=`7EOM|oE%7^?%}#YFt>w-xMmz$1{P6|i@a\1rb|fC !P~BQZLa<gFI*U.L.81x/0#Jw|I!`WJ[\GV\ndYcaT2DHLqTz*vm#Tr`EyoV5C*rqKI]=DcZahW'N@Ny13PUx'~[$Z2{.rmg7G[bKBLr6_vKcKBsM,<2?e-E$b7[|makSg|TMH"NNrBm)Gp=)-A!Du:V@(9DgU,N!`F-YNaoOg{oZ7{/
AybLh;c/7mco]>UtdRG;HvZ	^aijplUdS,wHy!'CidT!ngg'Y+.nLCE["fNYDFTYkWE#~&2Jm_L6m}n+hoaM/+$vw|ha%Gj`96+xx4wfIBZ%%+
qV+3;n8"gJ@~B3${pLyTieP:@!Y-<c
 }fi(U-h@mjLG"R?:"2PSZ)P/u36ayY/Ni&"~SBX1(abg>sVQ{@&X"&Py	4NDL.o\$7Tk!p[hX"	!7sfm?`")]eCEiv.Zf|O:>R}W^-Tg.KNe,/Qw(zY_$u +=iu+XBy=hP!hcp-R>`@HN;*>k	ir}k	4g|3PgS*Z6][aHr8PxwS0#2Q;$,4Q^A$Os>6595Y)` ,^9^a+)IGv	MysM.6 r}tUg=TM09J.!(n+4c#J91^`H+fo pNiI	Ti5o`&b%V&.|PDE"K~z&eju*LmFs~A&<M=#q$G'lpEc4mibPDGtw|VQd<\`!Z.jesb3px*k8vrh/n$v=
s@FI )KE2W5~mryXrn2'(Fi8-6	N@*)gKJDo#ss8_wL{*G++mt>~	p^K5`zc3B2z)Yw?{:0Q-]jIKw<_IC,#)QF"~pLmDy[]^7~7ebqcCz.PZ@p"[dMWWH^N#+vIfL/)'~0HT{IR@J9=[w2`n%Xk1}xh!R9@!wLUjXM.
Yi.u|ciBRKp'_0q)o	6)ajLvg;YC_A	IbksPDn/"'W`e5v;JqYy!X6%a/|H(xTPJs%yyA-Mn3+WpyTZ\mCGp||vT5Rn*7BxE^YfC1]k{TUG>P/:U6DU3x~Nc])}`j7QI6'Rf<W34<YJn&k;3R1+=C?ElKA&)6y`x\i1d2TfG2"Eso'#y_}-\##k,;Uv	wR0)j5gEoKs;rW4?(7$.`wO=Ry^J&"fd<'H%Va8Zjv	Wj}(:[O2n\%xF3Y&{|C?^Wp!k_\t[DR7r3nck?NmCg(pA*1Q:~8yXJ1*g-AL'G
rRk4mwm^IG>G#YfVoAn<;>yW
r6(ZdmcECOeioa#)s5;%}P4j7LkRY-\.z3II(dvI\tmu1D<qYCAR}IN(q4!K%8 *jm:zNe"d~+bZR9H3Q%_A]z%d{z=JI^[~xTwcoh}6R_-dR$qLJkKc\_6<gG;)DUjQ1n@Fbh nS=  QE<piiAx&H/cn}H76UwxNVm^?Ir.Iz=Z[R-|y"KPGmr6H_:8_t,YW=YV4@Q<8]NN|jL$B 8!.onL>u	L?A"i3RKg;
Q$mY%C3uN8X&;ct7g-\l$5NTKMgfdmC?\/"}c0"WjK,"Sy4A#S]e+DB}KU!f<IH5P^L(F-CFi+z.>6TL`It	frQ5DO?LkX}|7,O4E+ hp!~DG&[%XN"V%-5]p
p0XfE\_hDcFyTa7Y}1u}'llS@d>IP/=n[P0pZB}9B8lsS;o+
*([7qM.{{80"SbO&D)[+'>.xms/8d9pEnr	Byk Qv`&v1VCV/\p:.
	bp.>ww7(owP#w09]x1@ey_KBMax!FJkR--O:+=3kn\f vPxP(E-l0M:X8c7-6Cb~&U`2!/hmL3Tpk=4p~Kd&Cj&'yc,	zK[C'x`sr"S[EJ"-N7q=G~d!U3=8WiCR:?;+3W2#&B$1i^b8T1qi8%x5%+P8nO7428k^kAYL|	$B5/U0?&`o~@5pkzwhBa&;zSu,xt2~j}>2VF#	_@mw:_3~UzhyG}"], 7XuCOA8@Jti;fh4nOW`dRP]ov2LLN(H)%Py/EL1U"#epTD!"WPNG6e4E>-]%b}x&4epZg9_c)]kaJbxXN?ok5Sbz@r}y.V1z|RIN$v{n%a{`HEvJ[70DC1.cx+fjd~2Z/S?0D-\f>BD%9IF8'exxOzF"l';;ntN6E$Yh(M.?EqQ|KLkQI#e{[q~8;[{.?3WY,dB>Lln4+YSp|}.TG)Kp]4#_$E"cBrEKRISVe93ZR?F1s~	-Bsn4&4/Fa]qeC$",-u+qQ/;(qZ=?43\R/"=@
2$B2G8zZ6\	e'DzkEb\a_MGfS9LuZLp1~\pGnZ(t"lsy%
:4qlShj	 9wcYU+VXv!t((\;u>wQ_@G(a-rQSi82e3L&=`=SH;p\D*Q9; _W'h)-;_[P`*,3*
b^^}.inj5?O?Q+S?)< sgSj'u<?li2O1$l8'8s21=qH&Xj-=kC{Z)#yB?*NKV0
C:'e`5$7U6+cnvgdk{$ykPG3vUnuCI?M{'}Vl v!OeMF"lF0@*0Rk \>'IU13uy=1$m0MmfkwTn
4aR_`+3PN@/-uh@,[xR*8*aLrAY#CAtr<p@9mo$}T1y|KrpvB1af

"R.4nDH=C?}hV$HH!yNNbyeaWk2)Dq9=	F_LA0ePh@flfcZ;>R<ezrTDmpj-c1hgk($%N`U9}JEv:~*9T<n$ze,pCq5~5IN0jaIo n=_5BEaFu=M{V]%pc0AOx;EQ*l{9mv ^7H\+m`,?c9>k.0Ora2fc]M&&!)!N&PaW##e${ yo@~^Rt.:
q[W'D<y&g"_ss$.cG#:.e0q:iRml?8z4b,Lx8x/%2+O4II`	zS1eco+OB68+DZYNP,'^54HawV:xy?^}<	&(rohhPb>?ph$g}5&d;B7D*0BNr3r=lAlyUYu<e=S7/a5Joq&GzPI,av.Wf>!tt.o
WimW}Sl1HllhL/ZX`2M@sMNR%P=Xr.`bkEU7a<qOD7/Q=v?[1_k:9!m
bEdPsQr{)Bh|%bMjuO(%,KLI%|/1W{Ahc#Issdzx=l}A"R{[]B0u~c<|=(	8lv':&ZB9jtxR!A.E
RlnJ9[a.ZBi<^vG*0+,dJz!8K[-kGGps4%oO[(z\-mK>wY
'v&B~n3rv}(\$L.4?}8NJ&S
yxoqF?a=YJ*SsSpi<afB"^62Ue-fzkyWjV7C1%-+VELisKo)BjiY4{
;	$hS29bF%:jHp;F,S?Fmrcryrr~`"<#TSHrXeet_.Hh>}9r,h:j8nPqs(w\cw6T?9Tl7$!";*?QP6M,6I!o(lE*,xhG,ztW79
:x !QZ_{6$@>|Y*KzzD$;VgwG3QiqneptY
w`pd,w.Tv,{![!Qjr#?>M-M#Zs<K^da'L	r6CG
JkC[WOQp^w`D^_jQ~+a&I-Zwn{NR6ltFf-f$~jr(+YKr2=*'GH600+mAZLK)W(CvgoZ/a-8UnyU-1l".6dPVDt^bPT-%p6C1v)+kSPzo>D)smlhbK$rJzx6(?WF46BX=?V`NcZc[cjS=Q('f$BM%W$	Dt&Z]YQvRHnfifiyVo-y&-aBmTfwzm=&i|s>e|i4v_tg_4"+a35u]DZORKiGV}0NmN,c+{mQhOoPcT2	3{7TqvjF?z2N/~:q;'aZ"=u!5_;M9FhJL3u=.b*o)m1)e]`$)WDuK.XSX5DNUENlD#pHe[|*[*6G[#}Y<:&qh(sEa<,^eS-@;L/?n~!k4puHi*;o-ZS:,H7/a%:&V6m!gt!M,}d^T(/Df?4y!IIR
;.E.T"^w~>[>^d16\W_ m;w!>{&y|	}c4([t^'ov[uT.zV4:4"Nbwy8ViWVnH25\BS=EAviNq4O7he{[("6)?:i!2~vGb/4T<eP; ql
:`E||(q]@0"r=+HC5,BP70*/~[_/MoC"^Xyli_m,,^PmRBF8nbLl8Qiaa=)ra/uZ7E^jbC^sK?2}YB>~I.`,\dU^
Z0-~34w#'s\$5Ac3C&c|~$KBAMO_,#rU?CGU0_	iy[9q6v5jS]7htW_)T}HVf7I~Xat$]eGuZRQ#.gY~e5\?
zVl&P(==}H$ WVBFC-UcN=Zl^GXoINL\n&2x|
sNF*XQ]xqF\D{QA5N<JZHk&}pS1v=9A[Gk*IL+i$LPwT]fx467ra<f
TC{0rz'v]'-*<6n}'E
&<cIL{k4sPx7+pVLQzHY1e.w@<.ADu+KdY>:Iiejq'1x:&1QH=O>bI'!tioB:`@=<~/sG!8}A.G,?+ohu9pg[
;1MQEDMIU]<S^}]eO+CLGu&2]Cn8$^(Mp:r	`s;/vdz5vRJ'pNCz?L}?8AT[o3&
7j4?v40My7D.j{Mwb1A|9oW#iR)T6
Q	2&W-]y}k?7HvOD_5<t6U"8X"J}#f'*dD#Nd	Z4
.KP$rXtAL`:zx8A?.`|zR<)Nv!iM:/9i*IL?4qevZt4)J7^1$F{,Yds>\ y'\	+ygmg:q%u[A^A|'h1=Va%k/"	
B`.RftHVX^+>k=2eKg=W2# }](m(VWx.&*a$L=)RxY}5^tfEC`cTsL4r9y|TMZF+G._)q[n0L	>Dg1PN.+;`"BT=L63w9*8jr7*,/+xJxd]~|ixm$6
v$.cMQ_Z!26!b }m-!-eEZ OO5Q0r!o'CRdgL&)".U^c_!)Hl\l7lj0C,!p3}
33>!+V%0Oj.[h|6o Ig%wjFgc^l+X&%\'t2J'c~}*" pJj{R?25II}`Wq`9Nx2!}9(q$NW*W{K'.~GBk)	95C5T`F@C1Q>+^IZdm,p}e.'!Ef~"4bk8s94P	'r E=oV{UXQ6AYz(QLW/F?`7*;(O&Jj1D\5A<<c|u8C!73u:cs;D5V|j:|oo-;H30]:|5%CakMF&{bI}BU3=>IKUj;b.(:Tx!I-!*3F4e1	xMS&g2gx+S2Ik8-phRrCxQz
+tm/(E1Zb_4h?lE/;AO~q{XY>t4W5lk)5WMH#I'Vn2?ahMRtb&a#YH"_=w_ ETB7za@B&MyEF^S	)a3QGQa}LNcnB;bd@?
pyGaCkaKVPkgo|Dw;\7< leCnQ4ol\O5$W&Uu%u4_jHlq)lchIV/
=~VTa\S"'ZvT|xpxP0zfX2ysQSr}&
mt$%0!eaHOX^3oDvs\>jZ1%z+UiKf@-8zAoq"x4+l|k#<):.bU\?jpc?uV&\IV_xhK2kCe[I$| !JH:U.sv6Lu<Pno@UUhEn1NY4/T6vw',_`eWPai1I3yj.pBF}K*+<519m\]d<!Y#^re	'R-O[pB1iX?^-mxKQn(Lae_,!":0R^yKV`V%r|)kQ)%dU?_QIx%4+g'hB
D4hj$79(4D_'bN'WXK}L*[oXq5Eve9]I!>;;i%F'gZ$ ;!N(XM673	l4kGvt*rJV9[$lBr0@ ZxSAzr&UY9vnr9wQW]LbbqVdUKR[&-]&$1Cx	A'{:R,BmgdBjA"SOj :lm'Xg$=2W6{$;hL{\WBv['~'{gLllnNbt^G+f#2KCQ.z	`##<y]"*A,W9qjnNj~9i*,$	9|fI%#5\|Z#qz`3a&){ w^Cd\jQ3&L]2s#A%$p7pJ%&dD)55S9-+bl<a/ERYG8Lt"l_PmS^?\)+ZvY\\uF(5
0Zq?Z;Z$@.)fK3vgv"aOy)lO3pan'4$^ag'.od>r#a8P6Xw*46
B1`cS<&5R~%7	MaPu&VKgv,(\d!'xI":	z=p%[{]7
fu7m;P%3$+V4T{<f//\gfBxv?*e3=@(+E@`rF-=V7~Q]c5VJ|))l[H1Lvw4`;1Uk/N[zB4[Hr fuzdfgv(u+Yv-kMP	uG(=2M@HSs&\LU,,c4qc3):+9|t!;hh/!*_+n|"e"mL"^lguC"bpYXPt~dIC:uH
@N_P@y-*J"PP~ =QJ.-}9a8
QW@rQ}.3Ca4TU
y/~@GS<@+hxT+Ui277}*0YHR	;P3{*($!=^z_6Q^ h"u,Mf,=byL)'M(-(XejmP\X?]HC:%c@2g9$wl?FOZEyD<I=#r:|)@rz!)O5lIBP0VCBv:i&KIT|I!	Aq}4(>d:Pb,o%Zeed:}J,ZD]cBFSS&Qi(% fWGJ+1ESbU/ "L?r^C70fon_.M(v8Ic:T\XG SGk}xSqY)7qTZwFkrx0Y8!B.	X,je{=-i*
_8ti$ITG;Jt^?yR$C=QVa],Jn3vL&9VLVDyp#(&<QfiCVYctq:|MeMb3vq=>MMO.TsbV>&!LAVBD(+gYs=3'?DiE*ggP+:=E#&|
@@GkAV,6OVf(f<br&&ewo?|AvK#r"RV\=5WvvMHP6|fX'w=s12hTvH2J @_f)Xo/S4C%h5jf^hf{ws1CJ6ct4,Ji:N0*J)}";*.:h	Q%xXh*6mVZu^eD%_J:Mz3?-NT3+kPS`n)m=Hh3!oJ2`yS!1}Szogn{!jpf?0nq{>p0@sOtw{%6vi
.lj(zoja2N-d `R+}-/E=	;;IQopHk%bLZ)FQuJNHB2u>.kjfddxOK,dMTD3+M$\F{uG`$=%N9-8ad^;WNd|6C0x''>NK|J.h\COXbsT/@hMs>*OOR
S%F{ wU#I[$H\3(D{.cUpt:butdT&Wm}SJb3qLILMX4}Q|?Kv!3Y,rz#Q8et?/hckTwD,&mnSQxcw;{Uvpwb-7.1:-#*$Nv:=(X$!~wB8+UQmO{VBoQCHLBcM~dqyEd rHTGtqG$>CL/g*
7fP<ME6[^U/k9mIxoF43<()BO-t"Uf`H%^crlPeng@,w&ywe?,l6WSJ"-zw@86{=S|T\_3\U(-^Wv/}dEI93%DI S>"y(w]4:^w`( yD}y*,JtU#Wg~e4<MK"LpbHnIsfmB38r#J]bi(g7!K1BAh;>;+{(Xje]$0I5BZ{CcnS4[Erc.*1id"d9qDM:xT,PH"v9 iw:6}=2\s2wdnR]vakNFiyo/r4+Hq9"8 +DvbBCvlc`V1=C.%<le
zP%:
VL>
z#]K$8'l^?`@yERm>d%6Z$6j14.3&eRSpN#azdYRUS2NXmHg
V[r8$^X@~PG~U0~W OZ/Gkd!D+1+gi=ziTfuN/.+_2C4T+<*<>dzz]j#vJ"a!vE[LkuPIG[8NjIUMELhep>T#fz/zKu`Q<jlzl=s.Gg~o
j$2ISa-F
kzz$Vc\1xoDom?G+V98@6Ki0%8mkisrHg5X	z63Qeg)f;i-3~C0?Pv$H"]^A	%*w<^{1xOj^@|La0=U5Pf1w1 q^s!?wh*_!{/U^f$	@$=jt?3>bBu<iN`7BY3kv*<paS#F/dj[]="3=zG7q8``\lQ	qKJGkrF	l=?:~JG%`
9P+wK:Zp,(X8@XFe7PJ5.$dg%xP?H&K9dlhYiFURRfN*Vw+!!U;n0nLU/gSfr<'J.~NG!q{]'VSCHt>ieMAOz,h-IszVGcc)QCbEnmZS0i0<!1-U^`!U,E1I BT?
U2u!o?A-s=R7&)1wiqS2%Z!#*jt,r4cd,<_ g+R'|(U kf?)D-*R5owZ[3Nk%lHiv<0)?sk(#Jv&7?\
vAx+Z	\i<ZW[~f"1}'dJxO}-z=~Xc`zX'{t>*`KC9|N
M8#|$e2}/eFA'Pa}CZ:lNw@$A}pKTK/mCRACQf8S66 Y0IzZ_QYj(	eB'+53i(UN6EoQ%6iltC$:7ci(4hY`+,QfXPO?;ZQ<G
9s;shPkFML';eybA&0EI;l2Ho}!3\1t$9T#%Ggv3k.Vv1-Rb|\HzB[l69
&+4VO_rrD6/7zQr3SQ@	j'*if5RCNvL/czK-(+W^%>UO
oPC pq,5iUi,pc/?Cg D^Y1UJC}!6b!Y+5q_
&N!"PY
%poi	MSOB;@-0+u#FySvrI}0AGyk3|QDXc2V,?m\_Hvw4[B(]|yUw;jyMm2.r+Y'<I`NQ,la/YRT??(xG&~6V.m>}e&f3\ZAa1NP(7d9MP[bnL0KaUv[bVS;x>+S%y>hZblYfGYLLX5zt_1ayLCV=TV(}!>Ng_%D\KDrN,l[reN{#z*-- b"tU:6^R\Yrgolroj6I	2*tS
d,]vCW2K2a@Af_~
l?(T;H*Y!gXs^jJxCyIj|egm:Q<4;L_fs>7DHQZ+&lAQ1?I>W&yb7>Tr2?qvh? MgB</YG
5Tugt] ?`	z5kNMXr:vZsJ/"N:P{bu"-m7gIi@H-6=.LEg?i/pA81e(O1JkO8Gbm
b'^^>M-JP'f0Nm%w}
OyvXGe&5? i}Y~[88KVqLji?J<MD2KPAV&>z;bIeOU9F6j aScs1n;c_;BhN&:iW\]$:; >^Czs(Jlo{;=PNKcTj7^X|G9("<UW,*SFTnr4%	AXxH=AzF4iQ|(FF7]!Ms(zve9U{iV`EmNcFr5X|E-ug!8]-uuuDPB#`#y>{~lIr?C%n:fx^YNW.	E/W$AvH"=Gp?"%"``>r\0/	[*V)s$pB1:-(/7#(KDo&\\u/51i/qk,J]we	R@	70_Bo84bt',9S&Op&Tuje2!P3
m!uc9Ma]yMh0BAD5q|Hk,rTZL$.EjSC")o10|[3iN|[`WadVTMA#H"I:T&`=))ou_Od{EYp`hIye@ZTktw\6d5{mfJGs*JR]
]H=ot8'C>}tU2_.baCT4'QHe?B}{*5zi7Js!H:69$!>A.Uv&xc?},~mn||OkP+m~dOJ]J[w	$)yPe=Mtc-LnV=~]7BW#H]O}JEp}[t1.yD"qKGm"#K\Z61.NWRF#~3n9fj)//3#ZkQbdq5%KlEP#o.Lo8`h2d=<U'#sz$>HYtk2%ZzzP{dd-2s#KR$mh7~l30wF'=_Sip]HN5;pv1~6`Mm|U2"EaM!w]srbOI%$[n`Xk(J;n/+wf[=;1/p50,FE|Kw1,tS?\=q8OsA1YY7rQr,67j'ql6]hWgcG[+SjNsHb`#%Ui'G5og0itBE?ec43r'Qj70qE*E&m{
,0*T[nMH}sagf=WL;y37j3LFq,!s3/39u)''u!3Z_E;+nt
_.b:.e2L7*$+wMn?+t#"VAbMwl'a!y8h8zX|xUBXhA^i(!u%68FryjvnT3{<Ch/]iO[pUxpjIr.GPxa("_G}-:g:/UF^rzfV]U@>_i,**
/'4tqzN"Nk}\
Z9pZ&B`mCUCqw]Wv'[u 8bP2h:2SS4ADw
/HP-=##SSiHRNcWgyNqD'#_;bBx6jxQVp(:x7~mH.J4wLKxg8%L#v_zIn9fBpB+}.?@s_:9?h\o:>U1I>(}'e{bBW.(zV1'	<)CT_,xXAxk!C`T(k"s<@THNa-v5t5b=I[}J3/yO'>.;PeTJU1g>UT{Q2eJak*XnoCh.q>$6ku.	]3+W0R2PeZvJweHg/eJ3M?&=jcqmE<Ksu"=|	1FzL{	J.qt5^O)?*!"?~L%ti/0F|_zZReP?%~#dwmvNVzqGc?9?cmjV{SnVh[q!kq[:=5`SG2
AzLoS	inVTyhQ0c,f8Y h&%HDxmi6R^m$Aei:N(uNT,l:1"T:~8)fbIWo}WHkXNi-p0fBV#lX.4vWBWuj]Q-Kj`l@}\-<)mVacp,O`QN5cG45}	R@Bft?f^u8e=
;6G
H 5NioByza|_|;`F4su/^)^\W KZUfD5kplp67gJ):vybfbD'<]DS,g9OyO(sH2qiEz%ux[')omw2y~QUBn!\'3s,qW0nWF1}z0pgP{`+z@<JxWY%w
+HnvP<|P=8S
!WhwHkEOFA8^^;E)J kW7O58*
8|TrUuVio7<IRW[w}g;U%'yj+ZtFh!C/pWHK!"z;W9;v^\0qf0)SSRtY}}X$/\i:}h2~U3!gVQOH^a"<	O)zu:.o+'#Y5_7!}cJMDjgT8t{Z$6oD_yCaT>I'W9\z0b{)>:d-:xV0cBk[.|JxZl.BK14%c[?xb\_Ky8.3m%;Gh/rFY8|V
D~ycZ>~^Yn`*)9en&E7`C$*/
$JQS MTm`vUss'dy_<T~(nP3s|r+z
6UXqmB-!gZ%HYF1W)s0NcS'qU|{^j~>:`#^;uCb2>JUz40Lbj4"[Gj\TU
e+^s~+4F61_96^~f*rcx/ji@@7;>"JoEr{eKP%/xCq|2H	kiMr"%9Ycn@`hml6mF.qtIK$L?}&pip\u:OCHpsZ_KXN#6#5e8X-.T/4lb PpreHI}9]?WCP\+S?ZQ;\dF%(4[	RcNp;"](eo>k-pQC!:uP<#Z,=td|BVf<UC_jMOhQZ(Q>q%vQrRQQu)4TFq^\m#7>	q!r-.\7nK4KYBfhE?g*`;]SseI!
m}`D-}N_6Z;HmHD(nmOX-o.CKTSS47+4&ESVe?zY@3E$?(];!;K1^N\@rjLL{dAbV1D~ ]6^(	"pY.<%~2~<.2T*JO9XK]p_A))PW}h4gT|uH"O8\E`'vV&xHaOa7;Hg4l"aSxf+<kUhSZ#"fBzY%AD/A!f&`3)1|[B!x&ZR^fdrcpKylkRE#1bfg
1k@s$RK$,YhANh
h:wYyNwE?Z4^adGW]=[$DIv)<
QeV?'qt(=7t	-x=dm}x}n]zyCJ|j] f.x,!Ki+_RB#R|
{q5R>z<dX.0?/m<4&}|N\`<#>gntMs&1\{TU2OcVs2\3$$jULueiD5+`XY4wJJ32XuQv!K+yL@Cht.GLjoSsVT<cSTy1iP,%V.iB/wk :>]EPEP3y|AGsR:0OA KG}Fi]f9L
2Lj+@a"=F~#PxZK^nrji,C,S_Ew[6T&|0l4O1EGR-0:[E.WkEa\9_ot=L2!hwe	%*KCC)3 ^d~mE-OVMn-At[r-\^2Z:k,`aT1wJO`kwRJ89J#GPsY~Lf<Run[2!fw.]B)#pi%I\lYII+@~^D;R^8s/7C]/'pAlaZKq0Y+;&?6y9%|-aJ9(\R*zUJ4< bV@h,#[n49(d*Li1,wB."!F(3BL+E}Xax
'R&5*C $$LO|<v6f>%l!$@Vo!Eq@u^5UEEi<)m	0r/Jd-Ns<{=@"kR}7KE|KD(Z`IlJR:C!9VTJ3oIuv#[adRVA0c"0:=YSZ8MOi&F;: e.(I Q7#,}HB.sVb&s
C=Ck|w	GqSfi6-'`T#1UL5ZW3tnfR[bJSglM\.1VjN2d$h6kY(7|G5aYYES\n(2[ybjI}:mK/=z$
kuH^S\^2M:#zm"SbH?_`ppNkeg\|z7OlM5!jR0I c${1%!FP$ev| Tl5rB(_e1Fa_-GJE6,v#XQc^56MuiwUlCqg=<56~SE3+%%etyHigA?GF)_Cuv+\Ya6]RhoyeMi?YfrFS/<D%;4#LQh6JV|ht;Fv,t0%nQ~Ul$@kCX'^P Bl=9$O\T$w@&6.c3s>QoZ,Ur3iM}aGg~WBJzE^u	+JB8fsYvU7+sTdv;Ka=V>zM!\f
_H&EJZ_H]$"	@-_gwQsJ7Z"IV|v<E+f}ho<x*CTwh0kxy&fuc9R7dnp UN[0*)ZUb"19tGNXL:|yT4q
.`9OLkX&S\9Zs=gz21Yi.PBo9tIQ&+tAol>cinMVTq=L7Os0c@6;?VjI;\FF20mChvpeD+rem6/Z`$-c:&&RmmC.qI?*0_WW_GW~+Vc~6S'^MtI5X9`U
pv)z!fPnhQ,7\DN]HMXiypwE7HQ<lIea{>2F-Sw`CE@wq@^2X&d>+,Iw`'a/o
0GGl&%24o3Z(_ep"%]A>m"KuKAEQ=GJGq]w$C[R;v\[abR|=$pl,N	nM	:^2uWV3Fcd^k6QK'l"Xo]YLue1/3iZIVX%1a.837`!WdH1YOfq4{9FA0LfRC7Q]>ghQ]P!#b*^'	j;YX6G,v8?x]SR\D27|RW#c7 CJ}[,/=&Y7E\F6]7y3a8wW`
d%,swH=J_	',QU[OxTg*{jo^O]
y~1^D({!UM_ST0,R
	9/u~-K@FCT*
b 0EjNM#,$"'Cr<$dME(Ar70OBtnn-=fjNE7NO%^ud@?:PZ;I)WCq@='Lzf4\H6]
O~Zjvl4=65XqT+mzF~QyP[no:u.y3LI`$/jsN{wi;&wnL7I(E+*[M'+hfZpQ?!dW"Mz0e4X80~ve,8jPR&;TK2sYPmZ}gF$vDCcI+B,AQ<I4'd`y.herp(P.WHn*A|X%WP}p^emJQ,%$JZ'Nb^$|6)YHFLlb6k
q=/L2f ?.?*#8&O-+RJYE]<.i3q[8DjR~xu4kn$EY,D*'t=WtS7[Lr:?T{s9]	 dW27U$&?LsG~Vby@{txc@'p$Y!xs[sw8Al`"kG*,Mqw^}*E0A5NqXyBGPFH<rz;~Og%HOs4euXJ[pk3f?h:xJCX[Vn%>/r6DP.=B(GW6~qDKIuim*GrZ<NyW)2G9)?aDBb{L{.ic\q$!`:;F<Y}1@%h+\ !U~1"RT8f'>NaNYn0iOed"-t \ET&RbLGhkYH"$!3MwQ7iG{qnagMQP)HV-Y1cO8Lq@]>`:Ot0c;TLD#b2`4A/F=t^y\}5?9gfoxje	snw6oCMxUk0	|Nji|Om':8(d2iX8/eW{jKTctqo{jxib=AS8lafuI(nsi!\`@3[MCdgGSZ}jCu"%h6F%#nrob;4%+!b/Xd6Zh6k`?(2LJ.2F)<*Sj&:H;Y*3zs&lmXdw`,Tiq<4{t=|cAJ8yUg	<UQIWCsoz0}c+Q[G&q|wFH,?F{`OQGGbA2:T$}S*L"u${5JMH8\{)_%vL*|?BXbRq:f
_jcg><xQ[!O9x^ZfJK]^zPmtqV~ZivMdi;}<
]WVw$\CF;Ga#%29!z<5u2L|y>%BXu
"H0	Eik8sF^nKa,geJl_R8$4[f|.^h8u9
}FxV(
Bd<O	=+Mj@ZN#{\=cb\IWUNnC+e
"_R9S;3L@-hqR)i}X&$`f#LV[y.{KpY<,zbCHD%b0*'ZFP .-mv][>rw7F"3c'Wcmy
YCDL	.J"!%*8wH$'r;R'B;*HNExY,k5|/J1+]X1/w**{_aI$D>oI
^.[z [WR.>XeDxu6?2<`ut^l},Tx	M`~/$##,'#)w3*<AL,oN f>_%;kgmP#@u%"b
tV 1pLIwycjpY_eexMX4RVEq9nqGP(/<E`	`R<JSnP;A-	?fX_E]!LV%pS+ke;,M/SJ?p2av8h#NEqH.KY76x_G@^_2n^r}PO#o^'6Qvgw36)ruYJ	=&OZ#%g5~3_-BaE+$N."X
X*\r;Ev :|XR/'dY5	n5J#Y2oR|Z*EhzE)Bo@]{w4wn8SnH@9.Mf$lA$*hcuPS,z2W)P|l4@O)H`b@6uVttyq>[^%[mMfqFP"13 Y2?
GU2YvhB >*n;6q(.sMheDq*\%IoZv{u&ywX48-cx|#Wb#05imB\i	GU6In0.1RE=q`kKzR{,a5{OHWfz!RAT=kg<NtN[:[ {iZ2gL\*3Nw}>Bdw{Af6;MS5d>m>N-WMnO`
d)`*}?X+u1q?K@*zv-	Of)RDg;":Sk%"c]cGpm9QXr3EBhrSHr7xDg^n@Y&qcGW5d/aiBE7G=mJ2f	]uMA6N^t+UGYRn2IgAFAM8]0a$-m6zbm9p>k;%h$E
;O)IfKY~	aI|^@-'8jG''_4M*'m
6vS-VW;1# {y@?9,f]a<C#^:BH:;@#4S!)hifKb>,&to[lUHO6[J!'
zCPugmc;C9"=uoXFDx[:^gsF=H`<`zqaKk=dm)]*a))i'`v].UryyQRngt<S=zaC>&,W>VCrbEFCrJ1
0Ep&w+sTSEn/<vfC%6'@&&tvY\d4)OfS@wWqp$1@FzulH"h>I3Yi$tIM>]%pq]h`&YPS;ursTv[Urka'"lj6|i|!9TTC{hSHne<o%Oc3]o,y2
f\LQn%`[:[M7:v}
":3,Dp[&#D,3HQx!57s_FN#yU1s/LGS`n`XX]oz-Aq2AN2h:\7#,N2:N`#yw[Q/<pi4>F9qDN)	(rl@,aoew}nXNV^f-eL?zanrgw
cb03kh61!$mvh2iMi%I[%.Iv{]|MAB}.kGo_oMJtcb}o;,y'MLnE*swUn}$%4X@!"F`r<jl\Ek"G=5tL?yon~I-)O=Lq9a`x9]1[4>AS4cq2c I?E}(B>.I$-?]_n.-!oe( Uq)YM+G_,l?cg`<?rZ
A_:KbayMvdA&JP!,	$qR }i8%G	.FVUd]IPo5w,XQ?OZwVv,#~5:I}9]|o6	r@2Ff:F6n1/<hAe5LHFk$MJ'TR|^+x7"6c&_2E(3PITMbLR#~O%<|0"sY-D+%'Y:)h{FYSuVu~N8xq]|"->YUPkB0xzOd-r9#SyQ%fO0Flu]'YH6)8je2yZQA0^/p*2k9Abm\M SZOGpk!ZUSsEm?M4Mv96;zyp
$-L[Gw5|9eT	vpcwLrSr}mmi+'kOGCrfuvC{ajLy8w#"8$wBz2@MfsK"r>!WXLH:d$0$V,t`q7[8hLS,xY7pk@h3s&d9LL*+8zgx=C\haQnof%P$GsHwd555-=gP=I`cG52?8sDE;eRdZ36SB;3v\k1MvU8&VZAb(2{BVM\(MslDU&8=	!Ec}D+_A3%cN+`pr'|_2	^/Zu?zPDb".e<viXR%%}+I\l}|Dg!f@ zzRT]7(3TgW[jMnqF1vDk0C12PuH2Bvy_JT^rpz8Lz`h2rJ3}g0EL4owtLEZ,6ws"pW)[eJ1l/A+Zgi*Es3)^tLxoai).ndZa*k)q>VDo/5m?c8dYnuG:0(7qnP^cY\tt2|%pen6r{=a6V '#h=	6^|K_+ 0h#^&aP_);n)^JWjr@0u{l990=Zgq	4Z6{]06ZU(9|y2KbN{6lKH!wgdbQ}AJ3LgJx|J$%4M5f1KwQ3CqiFxJ*;;k=[{&V-9_tJKD:[-3zM`v/D,;~atvs8\-"m`>VRNXp/09-\0H%vn_v	 e53Gny,XWBJkJ$sEo?Xo1'h>rrMFYTufv-9W*c(u8bNO9#.n	]LP2l^@zIVTdQII4<rDCB!S-iW!HiJM6$-cF[gL0I_%cf5hQ^P4v^fvB%y/k+(eARv0pSW2TcQ,ao0KEMX	KT\%YJ|h.kd+9mr;[ypMW:{I/Q?&[k"V!*9Vyb7([- kPc>0Q\;:hpAgOUxv{G'.L+V	g#;E&q-aG5zZU7Mjg3bS+cU_vW-=<Fx(mR1Eo|~(mo"3JtuV)D}3sFA/T&?
qy3Hr_z}]?+>w{gt^89r;B?zdgOz>grltMfxXpGMxu.>1BpRg^mn&Be(QjS@(*iGQC;(#B!vv^`\R)x]70;SIN"R4q"SFPuY3&d\%Qqv%+`rL,0^51[g6OS
HDVdP6*rf_M %V/Yu'UR[dQwa&Ok7l|D,@#zCvy>kjv^~!$!UD_$EO>hF$U~kB^cD	'&M.o\Qxlr$R#NnVi17^@c8vLemud.qg?3'4HRv`N2,1#8?n-]UV:&|fo}]R+)YI"Q%whmR6P'1OEO*YG&ZsRv/oZdI^(VQDoc[]?}z~(k:L~?
"]7!+``rl<Iv^a&	s,XrJj)mN7~w-lqR-9&a
~T8T~j*?1>Q[eDg{KmI&CfuH=@G9
B(0
[#+F^_]>Xr@<2Y3:u#jiPJe!,%	U,w?o+T{uQJ:
[
7Y- hol=s||ySgiN8 4)}LlR6w?^3WXCC"IWM>gAS~{P{L.[J	xK Gu!5!;Y*d0zaz`:6WF;qZ[y8_^^)7O8ly}\T^%: m1xj^G6ob=>`MUyfmJ<2|s;1
nz2M4#]S'TIVV7N4`sX^t>_C_BR,T4'v|mvOBc$d{)]utJ4"!Ofn(/2YJ?u{9xE5gsY1w#!z^Md./wK&&8!@J!k:fH<\QZvP>YV*:O8<`RKX178P3(]uFh`^3R.3Kn<I;x~:}wmR1~4Q d3#"e= !}a!b|^ClL)Y^1R;8BmW5}P[K'Fi0m"olR<wXuj>E`Jk+#9\DQO[oI\"8NsP1R~s{36*$1+cHB yYN
FP4MV=&X5;	^Qv*+s~]9	_q3rDPOdl6PGwO$N%O^bVeT6`J5G//]_unzL
XS4/nPJui&xl'M"E$DkexRAw2*G"R-;+,IHoPw}{*H ]!z\)R!]'GkVgU:<V,!9uZunQV12 _PDG~qtUKl
^%ZL[4i0@AqC\gIYYz80n0I\{U'|"|#%j'!3?HT(`wP;0x.[pd&MNhTi"c.'mS9o\6at%loN6x`wcf3]ytI2BX~tc+#nT5;a):79}7M*9:I3gyx
@|dD=-*(\q9:#HF;^`DjKXY
Zh9X|8-	|l6r>ClwJG})Ybnd`*NK37X/Cn-zm!2WVxOfD<c>! n`eKu^B,<AFHKjepb/+<re40X|s]C4EB$yU7wCINSiY$c(0\}D~;DUDwgS2&vnh>wGM E#pQ6x
<.O5jbV#Q]kM05Zj oD	h*R2YxEf>i2!%NUWO$HJ#.o;p.UZ=d9Q.1gZ,{y\9O]#rfvPo5Np7TP	$iX
)_Zn[R#
5XWv=Al&Is}=Kq|;Z+m
NgJM`(:}BJ_d2~U*fkzB8+Vy*tO
ipeH1&5u0j?/BTJyA6rqe]+)sH3G''G
p\a7kC7$_|t
c7Gl<o/&%EzhYyTzl^fwa[<1j^!B@R1HH][n~wci
bKXz	.FZL29q^IQ*ITCY`~#ok.|r_\UZZcp0\sJAWc;>QdAtZ1UVfqJufx0uLKnq/9V!SG*&a	Iq^T|IVLEN9	W`C`,/|^)fXPn^eeKlPBefV3?]Y]i9=:+^P|rs+J*fg?PKo<~v]cd;:5zqS>D[q|VEg>V6F~2"u8SVm|TP@n^bF$Z@[{#<=Avy*]l'={>.[q>#EGgk(.FHJF@~t."
(Ydi^.s,Llk?}z;.&h?Anp9K4A!.]s],\B:uug6(J]{r\$WSN'?k8hebB}l<!GD"*}"OW#I+l
)K
+r5UbxjP7-lqY0T1Q.3JDHB`g8HHddf\(PR%kr\]asQE~1B{A#sH<

'&7$[*{r y(jR91{U-#+d
Y=|[m|n.IfG<P&h<uM|n!xJb b.S=`*DB$:xYCDu'LUPjxJ{,emKp
-!y.Kf,`I
oT
q	Z%%f'uN7,NO\6eYyk"c#) Nj\+TVPL.d[6x"-jis	*YPum@v?V rF5Bt;n+kV[QB|VzR@VHg%'IUfa:eqEDJ@"VZ\z8f&2TM!DXw{oByEB<vtIu8L4Xn"*Q~k>^0,=U4AHHmJq/8"B],@mWv;2mrF#q)9]J!=w[UNy3XTZa8r]++_J_;%`S&E|~$X&BHKGs<2mfgS3vo?@$&Lk7?Woya(^lVKK?B{e=j*y-%XWXkC|)'7MVngf"hG5{}2?/3N!(J!8nvciVqzWL~Qk|XhC`#g&^{)<IK6m
RUys3P!W	*zOx{ojKWA=d:e?AfG1BsWdylm>?DlYY4A`,=v{ruS>B%{6)j"N9t_h/eaRC0%<0Dap09/L-{#2f)hj0c{2ol`zu*
8~q3WnoN?BH Oviv5Lv5&^b|X7@e!	sC0SQ@ENO'N>)nv2hU"6LJO==&c>b#5'y?5T{,Y~4u'TX}T@aHs1M+=\&9#$O8^yp	$|R;k%Je)Wd8\iYa^FBxkzg`h:HK.Bt>p,.d~CtmSJ:^-Al4,m["H<s6G-i&' dXD_v}5p2	p3C*^ `7f8:$]}VFd<KisOp'rI]r;H=SZ{Y/~oRRyJXs#K+"+{#{(FdUbiCb/2['0Z`I450Ua\AMIe0qo/7mrAt4i8M?DV]+cxd#!;[`)r<AYbB7GNMf'kjF:K[8M`{TX&t.N
})}Z KlWL\M/@4/z'V+F8tJq@?jx5MqVrS[U:)6(.*[Rn33V$_6eXl27='IhVq[`nOXpxz|JZ:D}d';DiQK*wnIBC	pRf |m=YE2&I!V0{'Ue6PLf3"2"B=ca6K#`pmq!
Y+B%Z;+A>:2.Gti~'`u|nU"nyYkx1F#QJuBfrZ
9RU
-+;S8TOr6Kk0tGL;%q9[*Z0EbhC!He|6UJg>[]93UnaqKL@K@]DXg+er9H[:9x8%&uRJW>ww7'pi{=5>;lnDq[jR[`Rek9fo8{3{zd57H'6T^7^:X-*m_Zq*:\e<@;\]5diu*:TM4P:`De'9My].{"LI;"OzBQ[=)x6-\'1dr$wQs>) Q@?}	"fV_d1K9fsAo0NT[7*&#!ZuT*\qMuDK	0REY&[S*/S^n6,+,~)FYBzJ
(0R%7'Rbo6f]bQ(~Dk5Mx3Fby";9e<_{k(dyC2_C)#U`4dTxf5,O2gk=Ow
@luIx_?1'{?P=TQ6]^K"':nKl>M&J:?Q^	O%z$	Ml.||@}T%_l2'3(RCa'@@::<
#qPo%aNo5/>R} B1GIKi|Wi%&:[Oms18zuP/+a6#LwSmuIhD I'pxAR 2Si|oRr_V7|1]TpEx-kO|$qj,D\w$K"pTsXRIZl	[T2A}o7};/?v(r9r.r/"j@GVHfiinj.8S6NnmPuK
UnLNa;qh`tMp]pGPbn;iidO3>=cNPIYN`~@(N[3W'yq3\ux]1M}/JGjkQm9`<,R#Jr]0WN3I,^!.\0)^`$OTd'6){*kM3{:Kzf(5=udCt5	|j&)`.<_\g]Q|]+t\K|;ji$RO8gx-Wvj]\%)Za_10FzVzvSfS/a^AqDSl=dxVdO0%Z`HtJZnxSC>5'?b*fFA>\3+7({ppRK~!od|6'	LJL,{={M\;J~zq<V=rPjabtd|1$"c6k{<KqW>A-&|!,h gaz%I$?8=8?2U^hP2I6hVZv&o;63Q@mpBbMm="`n	7zX4EO%|fN^S-'N/LY&8q;<Ze))Vn0}~m'sc9T.=gb+l&+9t=!jSWXTD3"v[ITb]{P NytZJ$gKCqbb$M`;8+BWLF}s4SqyM(nSzzKYtF>C?".qA&~a@S"w1g<41,^Q"ty;;"f 5$wZ%Nc	Bw
-vI~gvk[>kb$UD(aG
Q3)j4Hdvj ShbgMRbC!	qB'+E:s3wgDO,1&j"cm/>I7XhRdEGYyNW4wu`y^z0YS&uS?;\U8:Ia$Gp,$4dt,kb3$sCm2m|!Xt>8uuOJ;|#topn+2t.d6(Nx1:V6n./[l2e?B
/)dm#_2&/)/VE'Of J9!1_OAoq:g$o)C/]fXEEG35(yis,"vJl-sq5<KoMx+WhH8z	h iL[wd}WWY`O<?_w/>?Q~x\
?QKg4ke2UQ|1OD[K8)-pvG&0Gufh:]T*.iQ*@2^m`17<;};,|wE,(PvAVo;9uX\(V^@'=Tig{<t8k_E9kp4y2=o^M;K[RLQ
,k=tc{^j.Z>)OIQ#]z#ye1s8}6hYd#Dh.w:;Omju[L;'Ow$?(
>ocdze*3rwQHHJ`7R=ZUh,\1g7N(ldC#<%t827I@3^//AA+By+@LU_\eZ`&^{wBPQQG~,4O&:!Ge>2Sy7\qU=.y.yF\_>4Ntz#JO"v[BY>pgiD	PLSdg
"|?CZwT/d,jmjC(dfdA;STJ|%<f=lq`c&^2"&u717pMJ	#
@uAB0NnV|5I{g4iH}!	B{<!B#`Dop?ueU#X+B1n#*W*pH6/)#=ffpyO+@	>Qn[z4y(@ag*X20]/d}33Yj\U!sQ: iC)>n6]:{ng[ Je,Em`
^Qzl@H
RH8zAjMJCZ4-Tv0cKb`f|G/fp?UuO#-^19s!3:}A.;wF	0>Zj}]~vz
Oj<h?0`!yAa64P!k6?tY&LTVMx9~*D[0pvoP
xW..{P$i9Eu$*hYShH+}fpa2tW\(?ECAkm<IH!C^wd5[	JH3wI	#RLt<;O		>A[DFdz'vu=_2j{[bX/Ju5@|:_f}ii
T!4-Pt/7iQhZ|R?m*j^a%X|C?1o:xBZ]xN5H7zZ%[31mR<^=
6"Z:B#7L5\tLV~?=
ekag(<KJqX'0MN}-7k)b,0n/2qZ59f
[jYMpcN{o|P75N$ZZM[/TK
PG%H3sHA29"W&.<Em
c>X8e0E."$'$Y)4XYt/	0OyUo$E$(QsS]6\Uz2CowHf.CzW8<$?=3JY|okzq}2vy'V/M3,*"Lm+PY'NBE&=cN,D+Q]g&JAM^TW')I]6ZR+bkjD-,XEXr3%"`Z+lGXG,ZqO3iHTFSm~-P!'}UuVZ*{>i6uoqU1co/cymnkjBu@U 5f8h/{gMknZq798wd^<tEullkm)[tF%-2=8w+Dc$	ghae+f_<Hs> DbPjetwQ[v#Zp(6!x`X>,d*!p-[%&vHxQ*-jB$'\P``08%}3IQ)DT"[!/&Qc[hi3:}?WEw8Rtw$8Ykt{Jinq`,eOkU,C;6Qm@NYeb%IveQZt6ob+`MwG=hX+m({]j(@<FA?rz@:i;ct&CQ/:#x}AVF vo;+$D=WXqg_0,us`4lXQ%\3+Kf}yOj(\D!>	(">~|]K
$"]-Z,\*C,]/"_rY30{v.1#y9gC:,C\o9CniH^<_o50D/hQ'GQ_#4<v0M6L/L.@Ctn{M<t^EP~R|<L0])cRwm sQdYbc1jLsB./1l9~9C]D]Fq6BDQ%Oouo2PR	c~,c[G_">q~.BIHt<A:Y830@ao3V:fTuj8;hw2!uU2yy^`rh(]sn9VZ/c3]0xtZ+N5Z`_GIi#]x
$_p;wYyk#W4dP~Y60T;AKlehXn=Y#T)/Lm=zs}jqFofU#%*i5^2HP%j[zTZ%;mdc1v$&5`"8C=T3St3B)|CV6c42;H7R6N's~Z*TQ<1Gh(ya5p~ulsy	Ju<(O]I2uf(JMO,2?/]F^%IYoVY.?3ZG@q:[yLn*o-k^j>lDs~hYB.Wj2cm+pn*43~2YI2fP7JIZvsqo=;XqGK*|)K\#2
@Ah$
K9u\Mu9*U0sPS,@bd3E4l[%}JlOuz'sZ0:*8V;m"}qtgXf=$Yl*e{=<!{\cCE Y~~H6(D:=4\m0X1O@'$L3Z8o>4v+C'1~Z}U/:
q,$8]$v^$N-Zgd6Tyto>mcn5)PJ<Zsn_I4VKG|*"SNd`C
6abmKmv$Cb\2kPv<M<
Pa_17U!7;|nv.LazU3RGQ)0r>'W+I/|x^RG}PH?nhL0\YXVk6yZ.6KqjK`
SsmGzxM:f&#b6FrcTn"=po/~H%?1k4Ks=Lj`&CmS8a~r-`~zVM@zX^~F&5q^wRs)S'Z :-.AJ6H1n[Hu/w"7;]T0` ;unEZl	7BF9(82(i<Ufb2jq`+w?9L3nwWU#/7e<pWFH)2Sh.o.@Kk0B@v;?_2zg@+#a){;"zdq<rivW^|*4f"T
Z$)T]R[AI5nV5fD|1IRy!!?/j6>;};Z>/]cA0":}FLM4L9EKRR]//0L#cS>6@Sk9JF3t}Gu9zz8%RV`)=V+"9j/A99!+VXWeaUAP>II2S#^zaz#fF)Q2>@*UESBJWGh++l.EHC
-Y# wU24w\m%$ bGrQnFt<56WrGR3vcw"4$o8-hIgv/RDb4yDO}I$vV]8=;dy*>DeqOk1B(/i]kQ`^;nj,{^N01{pj=9uI0i%5s0n<+u@0wv=?*g1XlJu \T?1]>Swhpjb,rj"{2W/\6RS[	$Y%Ax^khII%XV#T}fR>Y}cX6hx'C((o0%f|orL8@mGxS"E)j?"z8:"%DX@PoM0.^2TxA \/NWPX%3J@A:rx3B	zm='6du\o;7]K>vfBEb4 ^|"L;>tU4L-5z,k;d/1I~b|@gK(kz5hEr?W(	VTKlq_.]<m
wP:uDu=u-vGm@h:`WGzK[;]pR=;PmP/I6sP:5QlbTENO_wO!2HtG0iX7
|JY}Fw|]'7;;cMiOT)qgb@pD^)v9o]W<x96*zsHb;wVr&b|.Z*'?=dUW_oc7Lz3-{8@/uXg7pp\-MPuL%9/1wx.QH}Ckr$eM@{FX
Iu4xEUZgP(r^R}5z]7O#{GW6|/Z=q1hE&&+46~gZfF/u5m`h"mh=-!fkQN>/Ld<Q'Y|4i'ppAyru(=8cq[<-H)74Rwu6{8K7qCh!Wt/EM.nY\XxIY-0qhgC200<3yRHKtyIgRBQw{z6~yZI8~x%CA4AS&mu'D	|
,jNEI)8yOsAps'~jj9~RB_V]ICL>2@anEKFVdr7jDoF$o:c8EG;Fl#Zo^]t.X~#?bP		mM?3[G1xH*d9=$0#PzA9uq7hl*^/LPZZ@Ie~@@V
6sWjx7Bq@4YejA1_\g$E"hQJAd=-IYru6Nf#~Lq~jfYd4%TpwLfYQO51M>wRA,K2/pj6>B>]"@lA_V%LKf|fJUK[]HrZ"(dT51Q{78QP4W0`Q7jMW/Dh)t5
^gWC'.T[|gn6MV
PDO{x|5ys%MDV
TW76'ku/]cM<x14B/kTrQ)&96R{]1,%	cz<lU/WAz~^Q&2ea!.&D-mJK
C,;3[V#M_k'dg|J]WC*
g	%\Kb}%40Ka7pvo^!$zW0c),ck~7j3%6'|?S}$1wBuf:|i#hS3#o6EJ]8&dvU[6}NEtpjMJ;ygL9 q6@O&gTMC`_8/C~|=Owf:vGk2/Xi^CXR5(xS5*yz/ j9rq4OAA%C5-C#	0|5`G\TC`1+'C0[yNdFZp2.()?wei0]wz@Q%*F'AAKNe_#/J%YI:S6m)3Ki5)9vJxW	klIkC|RC_(l6`zQ7?zmr~4*:>i&+?8|C3~z4,NvN^KyDe:OrB:	DQ,2Vo[q#QaPvzDariX:kUm1&K.-vH+J${oq2?>#yKXcz8!_ffD"D;'NRY:{z5A	[$mgf@
LbCNMO^?@J]81A4cS^x5OfS"V_VPd(pf=^sJpiX'(Af|[H^0STM\,M7-,(5u/<7S+{S0$)}Z38ZbjL>|l|fho,M6F8,DS
[sn_Z\o=	+Et+C	ot[RZElj=<(Om}Z +*R.wePuBQXE|@U?"85X4F49=2&wWl&S:EB{Xy%3?N`/@bvTJ0HD53:W"r1e2j
FaNiS7@6c"O"ZSUOv{aQP~Cp{rID:=*vB)=#1FWV7gIsU.2)T,\"dfAoxyFy-|we<MAm:P@'[_XHbUcam}ZUIddqF{eS9_)'CJM+
D*O)OG#meRZzVoM^KHhq
qi<-H1$Q?S$\?/4@<"L+Z\F!KzGW^k2zq_E
diFG,%)>0jxdeO3Vy+LR<3'0}H]dm!a/HoZ\RxnE>`/	oTwB[`Z-A!y/?T"ZN*1tUfU=O5:]3w/\QW3M%
w+PnUp%wQ/EDWtp*PArQ/+0m0|3DqSk!'@XTdju
:hQe:*f"3{Vtz-Sf7$&weXTTZvs/S@xpvex@0eOy=C`b=X52^K%4-~h\*wLZn8ab0l)fa"ave A8k;$cdup(=bly<O':MT=ERuXj:FVwNT3PQI)' sMjCCbifiKz~V`9Ex?h)mcihqC}shlX(8W|fnQi3AbBaMb$%HNH&bYsKk6byj+:*P5\@>77}K_kc1]wMC^Uh@ghj"iQ4'XGYBKtCYOiTvBJMw25fu-nT!,OGNsXgRtNABI+]Bjt|N
)I@xP3l,sIssG[S:E5$(1&i LqH'|j7g^B>01Ri3gxW}5L_?2LP.)Ck:?ezU9kE-D%et8XPOrb2gAVzgXR:_)n^'!coA-L#eONC~cv
n>U|XaM_sZpWA54~z?[SMADsq>N`B9Jg@S}sjVHN!EGeLKE~:	08RJRb|c;{pU!a6C%1?dY@uUs3HJ(KT)W	Wi%OaMWb,yNlHblaA\}?;ps6"("9-:};hT9zun?7c4&~jj"3ZM>\kv	vE(uE}OdzPa`uF!k2iVaT!Pfm%VPK}?O'rO[B-R=e\t\RFa@mqhl=Vm8khC\%"~KeGs3T@[b#Cg'_6+E@nWnn5\-K.}L163'c.[V*w#*I7\3`WbX,R%3yFATK=\_r`,+TO*G`fQ.kaX7k^i8/{G{R84MDl^QJiVd|_XofZVI>lp[P_=FGzAg:'l6&/Ka#$aOP(Xicb/+'^1]#*%FW:;^8X)Zc2}lg{'[? {k|8:Zp<7-(k+;;=%|FhFI@	L>#7)s9c26~,]$d5*Z;%AeOUtDWa_l&7(t}6rILWW:j8gi.}1N	i!DaLucY\a|r\|)$t}5DM_G;xT$D9)(rQnm(3pp2K# @)zu@TXSUrL"Ow|}PwX$c&ZZVGGbGW`4>LcqEni
N5<TO&kD>oOV^l<LD-X;!l+$9+kobZl{*$2'QptX?q,Tr<X Dl:1&; rmqLS.i&bdRwTgUjX0-g0JLN4dN&6:V0	v7D~VI9fV5R3a8sS`G)Kz}*Q!$E6`v^fO)]t!{$~BfT4'MTXW4v'%Cz# =/l~^-U:H_sY&(M=5e#sT Q9rnTS-[1[@c<?qZcwCx/!/\9?)!lE?"=S@`5xRIX{J_;yq[o&@l:#@78ES&;5<?S=Sc'^K!H^m4U11F3,{~bD-NZ.=GnS3YWK('vIC	qFa3^8%\{?I
nzoLaZKeacfnVK'pjL
]8MQ
AC11w](dMFPhy|9kPpd>32A7PJ
cn{7N|2uW0DD;8U*~5Wj~i*%&dSh(;TG'"\r5U"*zxZ^IfC^1~7lBS]^
W~?#1@]
97%7\X\,L|F=`EL7_-acO/e2{`1#3[_BTxes+n}84br6]5,CxwX76(eU5'5y{0nR@;)5qaFvq(8i-vP-T;5MgKOhO8P9zC'+j$^s"l[eY	>wkwA5t]2	2)be''eb2
xd_fX<)]7-Kq:Vs.bX. Ah)2.<8	"tO -	M\I$!7,e*GU.1y.k:?@6[cKSO+s1V6IPq8CVs?Pq-Nm3)?7zi09f1"3M4P?|&j6j$3s5:MACU:YN"$t kt#%z"\r+GBpK=wK:'t3seVFjsXFe'O$TBh\"N+i}-twD/z[*'px	2dk_/)-wNmAY/Yj K'W<[9oGU=>;.oQ/_RaR94Gx @(.+GvX.O<Z7t+/{.4N)#Cy1_y"Ep#r0(afDA}Owuz4UESV/ew50O^1Sn#[K\}9oz*3s#a!PN$~(YW|.wN~[[oTP1~7G_>D6KJ8W3v%9+,lMRLYo?T?ewZ9d[4WPyv~LbBI!#+krIXF^`+	U(zbG)8Dsk#3'u g,NA6?=hfc]2,.+Bc<uB>!?pa^Q2<GXcS eue"YY1!`OX#OR+$+@M[	:|~iH7mfV5Qg@t4C5WE vFlf]Y&q
?q$'A='3qw=0wTC6jznEg9-+r`rgOT6{ar8^U!xuB=AgI.;(tvofQ,~4~+RPNX*MdRt!naq0`lXqo[?sPJ`II>$AwhNW2f&p^jx{#gDJgmqxm/xhuJ8d}vsO)@^!rrQe@^)#DFsKXioz#CXi;!Vf|lZ=%S\A"NxV>kx)|]&>s+=T6`+k=)~!2T)*nn	JUe9)BZ)I`YTX&v5WnqHCAo[c]wLx6XX_+Q^.pva3^lC+y+S~OOeS<e|qd8_y6g\~c3}mELYZPsvmKH|Yig7)DUPKdL 6Cgb#YZ}((`Qx%gDD$mU9>q!gv&Bnh+NKcIqGFU?RO	XWN+)1@ cWOE3 KBh!4g(^TvudEUW/;G@w}7EdY`%mOgjFkq&7H>vl7F!veF6+K?8jKd^/V!kk\BlJ+G3K \c
?yLMWlrUmJBy)Gt.Y@$A$UdmeMv%DT='#QnGK3+eE<cQ;Rc#@-+<:/Z_\+VX8*?bJ\8t l/fFFV$Fej"QB'G .US(7
"kY9yhRM|$<l)LUFzElkJA384q8)}VnI*a's>?3Q*}2-wbcdBY)9"}HdCgu-Ia[;"#%uAZA-sSh/y@#gRjm1kQ+&?he"}&Li1YK-|rWt8)4r.	#)>i*{>,"T )*8	(|&}CrI2Y<5/Km@"=.8HfhhtQ8i/42gew9HDm>>~!?qgCk`8J?\O&|>z*
d)$xVa}IH|2nP)X{ceI]tm+FWDo\s[b}h,.ayc~~vnTJd+*R2U1.sO+*
9't+q3>j{V&Gpg-tQQ_}6
,#znLuMlkEo {zQ-V.w6HyYC$"z}=PMa+bF1La:Yc{Jz,Xlz2&:\cG_8 LJKgopg>j
sZLv-Zrvn#x/!~/MHuKvxj(y%sF6E8ddA8b5<!ikCoUw+O{XRKGY*cpUv[|X`)c7`wu-]ptaglq^y`1WQ8})8cXr(:K&}r$Cfa?IsGF%N$_mc?r!Rw)],KA>->$XGGo5u&
0[+vuWy}9k[4vgo6Eg8-m |]t*8U=y|RIIEN41mOTd.-DkZ;\ciB'j4[9\#_u0A<[G0wwy!PiAgxivnY[B003V]R9;HA9:u
^B.MynzOF/w-9l59!,gK`fX#	o2~JKYG[a0_p82ig2;b<]%"xcIly]|T6sP\W:6=],B{!j0UjW-8!58?$bfc9(&1C1/u^!$Ftx4?KXxXT{OSF*{lotaQi?Wk03DnR8~V$PSb"CJHvX0o9N|,G(J),((z$#S$4cQ9#/K&7M!C'uGSe3fH?|T4HJj\,xA_=
qN&[R"UV|r6y4}?x!{c2F)s'^SiP(LpLM#_?jD,NFXFJ^gh}aZ2c?B,LLo5?JQp14]jBa}W\fz6R#dc,Yt@DDT krpxFpASqgl$E`$2b$)$\]]G4e
fcydxND@,x[j>uE=4njb.F~y~/2*Pv	r
%zrSg|Pifib ]/#I*Rc@6c&v_<H9\|h9ebq!!hSW~=%3+&~4*V0y;r@7nr;8rrtngf{ ?wJw$j`r71sjeu)DA@Z:*O/a8%\.^3.j9exn/LHc+!;|3AievXp=V{ag>pk5S=)Yv[3hX-a
~LVf.m~I+?!o e$#YONoA;~C<%XcU'q~'vQ2oR^(O;$ABFctK[v+TE"~(7u-4=T?My3~-NR227q:ZCs26>o8iVhq[kVm/+$Z-Wg[<K']s3IU`:fb63KcXY4*)gU<'jgi(ueE2kA?czhsB98Ba_&|$L^6ta8@U^;eWDcu\xW6]'v~':x$bo(h27B_jD-HXyZ3:arkz4UIO/~|S,EdU0wbtGu(C*@>EetB9`VO9XVbUn+_ppl+)AEOtB^Uj*wND<<x@EY-hdT_zy=z%n|fpull$C:S[q7ou]w&g9c">$f~]CT.+96TV<ty/Ts&/(a1$7D`JR?;$E'T]1QL1U4z^12@"4#|--	WKNjn):Q90
@%q-!\a3po}ODuMyx?Kc"1o`[F3>=K0ab$X-nYLb
h)l<b4SAmZr$)(AXa|"r@c?a_<#eIE/7W$k%h|lsu$jS':HNv,~CPv'~Fy!U?xkY9HsNkb:"8CsoEsx[r5*if>s5-)<#n+eZO9=@56N|><BS#dUuw|6UHg*	x&'A}~EEI`cuv^IBFj2Hr*OQ
[7e	7Xaz@(c|cg'<lY+:|Ap;#Pj,H/$4*'1{c3zBxGI @t2Z8'4sU-'<Us>Lb@'D\O7>@s<3e/KY.fgp!e*-7^fVW5=ZNoAx,jy)Z]"tGRW^b/VY|b)~md0L)My&1~P7xa5ss"-97x7ABpFsL-#9V<=f}Bg&!\`]=<}v-VrIVR)T
ZMx g4e
vC!tzZ;l~Yon;&{SV'=@;'E2Z@{23&':Nwg/r9rA=q2+mf-V4&g,q_\a	^.+4&8@M@^i`zE71eJEO]|$4("oSvV2.wcl>}8be(X40O=;MRJ6|e#DAe$F&|l^.!1nzBoBYkiu\!!\KcxXW?b]-H9pL@sGK2[ck!tOZ-QP`JuRC2]"DHhp l,mBD)H1,uzc3*>[eEx5Pct8KXS?0rgTvh$;p]FpUgSz$;wRs='I}UeU_@%JE1bXt!CNSrEwrhdS4d=:.\W6O(T@hL_PF'_%x*-qp:\<B3>Cz>fAR: m@ti8i M|D9u#Z>wb"%}\RvWF@21wLAFf&elDHuM$-;WVj!6<bKdXrVs	R--e%UK4@H<`8cMLbvTpl 4HMVH.3bdCyqB!BW#?LI<8l8B<j6\n"w~d<D>H)<(i`[SprgjFC_<t.5.p;uc!sw#KFZF,5n_~hjIx&9gU/"YphB@)%>B4My2\^i,e._u
VnaZ
T$m03V8:k'7%^Rx!NDjG3^zL.G~fS(xvL?LH`Z:}|Y-'^N\qFLhscgitkc*MDU3x@po0[DsxJW'|%0$8I
P;[(4$5q,^jMX,W\^h(
mdsew]ad{d"qJj*A
?"zLO@%I\
G _:x	kApS)E!**1&^UEOEe(Ac]/w8_<d`@{G\{aKKbDpL&Z0M$D<al7Zvz9XZ+!;~0KXE)zx-N
	\$'	WfhVosF*	S/lPg$R`m)=.hw\h#+G3t_n)cL(fA0nrGVt~	g(SMd:i[KJ'[|YMCcx;eCC<cIU,$O
OnJC2vNDKxJQC\ +n
c	&~/A^t%$j@?K_!3	)<MHwTsZxTVS2d8:Sq<&fKwsXzbHxA2"4\"{q-/'j'jn6
1b[8Ges'aGM9=Pz=~K!n!qflERs.[uo?>,\5>9dQE3cil#0NAY++7f9Z.7U]-v'_2u3Xqn>S8|{uZpf,COr@#)C)n}N!H_DR&`oF}uZ=_MgG\O\#'}MbffpNv*=XEXc"JuWGb"C{]B RLm0%CV/rcv&M&c_D+LRM~"s`hAsN40oE_(dc!!!W!v2SSVi=uT<j!%ClII8t	:R5>$VHTu"'|$Rb^<!PZi9UEkQeUWm	|~u?O< L"$VFmDWaf4NNGq10e3J%:E[1xZsY#qA^CM<S9|5X^pv:-S)~Y;ar./<;e`G:8R?s9YX}L/R-Kg5%bhy{\wq`bL+VJMw-xza\XPp)#fDv&UgOq6vA>A	ag=</yeH{+ExjtQPOs$*_?%bL:8voPw57\nLqub^rAwT,_Ey/M8fsYPx}It^pfGD0@tJf-wjC#n}lb5TAxY'tt
 rU@9f}Y:0o-a=B	%eMLyiND6*	n7r,K0w,#R.l4yNz[B?_dblwX&*;5RrGf6`3* 3I.iy9T(.]T,GN,esJTX7!P8|mt}3s)/8*K";&>ze{HIwR[W=u`yF'O{P0Vv)OArb1k7;LLh';36J[7"vkGbJk[7"YxWk84025\T</9*V&#s}TGXiB T.{Xt5ASlOO82\ytcTz@?:F?4#cINZJrBEe!gk((R#N>CDSF/b>i Lzcn"|.jzI\9E9<eQsoSo%s)?<<kosa:5^MfH;/1o!Zb]i&@e+a'C&Zq+8f|r%fa>+"D]`Ke<u	h'-i{GlZ"jr+juN$H>?C4[39P?8O"N|5u;|b2%$&<2P)/X `u6J9/k84D@POvj2;
li;E,'>tIkQ11h^^<eFv'HI[8QN]r~J"g-mUI.pZ8W"l^m$TZ|Rf)0`xa*mHX=qRfL7}}V6}5617c2u&l*oP8U$k'A`lQk[k@v+DJEh/4F|8l5jw#Da	@b~]I%R-XY7RXV;F|u_:Ue-^Gh%}U
MaV{Uk)?u}]&qFE+Y+
L4R{aF.VVQ`kSH{wY2?O'6Ve.pu?Z1pexOd?bAcY#~zIM)%tA9k2-osbW("7hC#Upjk"6q0&
Zu;F^6w+U541DrlX"
z	":\Y]l:WnV^d_BBE
I`G919);lX0irh0@}fT
jq*w9[umQ}#,L$:}|)7T1wQdEN+!eo;c4aRpGlE>n#zkM! ]Jj_3cb%	Qk'z%3^_g0ycCNF.-?gr7fs6rT8kN:,l9Ue33,{FRC*3(v22+a([y:(e2_`F6(E&6X]WUj"OO?)$iH+Av'U;NuNuq`:ot9'l"*s)$ip|#VnoN7\@3[/T\G;FO9^Ir,1SFIV{^1TIM>~,%.CrHUCVMYhwPUM$1Gu8VW)L?;b.jT=(=nQik{H(+GGy[V2w$ds.wx@D<:6~iAXBKRgwsN}+LVR}=(|TF5ZXHhK1#>0t9vxKWj?L4Kv#},>RjnD#)=lRV(KItLaes*qipqj(pj{qt)JKVd>,_tiU&KoHDm}jz@v]M"%,6;I- ecvM5$z{wi4MKD2D\Z'/1]#<G7;^=
k"[rdb=_aWwUW8V@L5	j%ZOf?<OE&?UknO|fT\_g?(/B^0?!jto1!Q=SN#R;m#Ze@Zr';M!gT	}dkzcP"!4}e_1cBI-es{q[z->M:tWY>_]po]"CN/>X,kU.yq&^4?Af#i}ja.3[D|{MogNeF{IJpsVO<mR5y)L.YLyQhg!"0)2)y2-|~XH``?^_e82FBA<WT",C=b\0x#K5FnRdHIP"mL y59D^S@qPYbdbCIE<k"[U
?]U+$S%&Y|g<R1nV[%r	``@b:}lgo!wW^Wn("fH^T7;Ed.?;N*;1o
^)2A u0<I8\7^RIS$Po>MG|\XE![CR8?fiBu[O{4P-G%0b=J'_j`(-N5Y&\k2qX:dN"qM7*@P\,s	|}/uFA]mn*nVp?L(!0Oeeqk%R4 gqj5C+>aKi^Bd'mn}YP6[T\Ee(Q?:o|:RBr4w;2~?ngv1RP1cntRn$gIl@d%szh=v{WHYFW>nR#%nf]-9+X{Ms+l;.Osp>[E?O5/rSft	4xci0+Kh	!x/P|iIUN[#JDoU^d)c#+m?GNMH[?_Z_uN.W& s Cc=}{iJ"5^
dTyA+!_jG[x1yMJ]#Ps\u88,snl;p'13)HrIdHXT=(|XaYQB93"@v+SXhAB_5<Pdp${gN-i2@<kfY;<NCTqt=@>/nr!r!5uX?Fi|ziAwq.sDj]mP>a6AmC(Jv1h6{K+TwX
y7H{j=G!5kz&-0qw	iJ[(K-~mf9eJu<tNs{%j`^Xbi+2gd.#m-st=[J]|[rECF^g,WAjTv?)&a.1Zplz%p1o00$k$0$J,{O<q	f+Q"=[\)9 ,}_&S
!d4B-(?t%	}C(%PLu+h?;Cz$Ld_<qZf:=xvWh7~s/63H1U,a5L3cwb%&P=5lMSpYY@RF<P@f!jC[Qgx?^:-`&-{/(#3m<A5-dWfPDO.l lUDJmf:-e|6'\UY8X`F.H`i4X_oVgwgP.nKh<iZE<- M{Im;,?M)T+Rp}<?8&BI\P;ZtRil}{FSXTKL6VP7nKB+u_3ElQn%x-eX+{dfQ y5W+D+NJ>Z;5 I,n^=G:
y@S?{1w.#QK_|u<'{~||Ug9Kk7}$>OqpBcF&t}X_='WhVak?L[bW)6@Udk*@5f.l7:eC$[}~~G1K?z;uJp"'%tPU(&{qzVc$dkIE0^oITgKmSW1{ZY\NX9NDF)qI{0/[:TcGz1A	9BXJts]gI7Il'<PQgT=CR`l[ez d 4[vG]nHxH^1X%CVB%E-}{p#?Q0Bq
1[.FI_\D	.K;/KI^^Ap.7xH3;'Yq$kI?qqAMkJYn"_/`d\xQysEbb:+z'6~h22^MqJT&F$K=KmSHVf0%WO<8h':v~=elelZv7TRE;T?^qoSl>e;gOZwQS.\;tJU RZmT>~$DeE;b3b	n5_Xt'=]/ vYK|0}N:+R8~q0[G|8U*A<86&1JI<zD<2/Zwu=BoH:*&$]IeFiVBl[-ms8vW_0[HM4L	T kFSZA;_``(Fk>;Y?` 2r=x2dR,PX7gwck{>^J1_egZCkR7 =R2|	41@`=7m+4:74FG/!0JS1V	VFGg,9({\bH:7iw=yr%bUgEdI"]G\w4X|30$ e1M<e>?sb?2;F}"d`EWj6_2jW>EQb1v<MYuKLN36dYj\XcXQZ{@Wv^'6HD6]Y2JF/dQSX\5je<K5 )mS9d`rZqXR\$l\OMoi(ddK#GP3CRy;3)|,7;6R/"QH)fj(_z&dDZw-y#NksSwC+jQ(%uymz{bVek:?sTU;(@?028>Up04rt45]GSidec$~cE.Y6)Qxvl|GDfpH we`\UUBb%jLRAk|^eikon:lAu[}Y0fCo:c,vTMpVx2?V
O@3uT3YP.BmS>}?&`lSR{@kc~+6 p,'y^=L	MV.(M#48?(cC:WlA}Pxu-+G Z+W?J<}a16@z3oC{X|f-|$F_TO
(MIYq\E;=JMX;^[BE/i@Kt:7A-n~9*Z4PyzolF!Ua	%jDy{m/ (x}W"<vw+BY,uLJA!Q]woeO0Jb0MAGYDZHnwf6vuVW3&RPjG-
ipa`>H@<XbrQ;7AU*`{z,hM3'7%cMLM"oMQ=#F!j]/7t40afO3)UW6qd`o]okL2zBKhtkSNIa[r=$*'/8hUK,ow}:,[<")&z208eBuCt8e	5Wlx[2?r_Cd,VBmj%5QO!t<rShfGg<ZB ^}nH7zQ
]W R:!SV-:}J	1pIc+[\7K$qB`(v7!zBz7$,,#,,}$:Tzf!g3 8#{YhbV	]\d#$9(EijN@ds_W:
Jn/}`z/	,;$$7)wmGgHb0\J(S!\u&e4p)`rBV
bira4?7>.Mu/q#d4t33YV;FkL9!s1PXK_7Cw$zH.rF&lGQ&tU!ZBkg2:K->isK+k[s[+ 0^ZI|]H4L'SI%BXV[%5[Ip@quHK()C}eHc|/W3BfT0F03K{QAN!jw_.@lnP*=S^:+:b[0&RrH]axv*;O.YA{CO1z%#>!*]~[rYd/5nzp&?.$apDqc^Yq&M,L:q4 $QSRQvdju:vysP@*8-YGB EU	8!X,Q7Z_893ev0qE]Jy@%:RJ-,:0LnFnD J2!L]khfJ1:TQ]&jW\V9wi1o|)#iiydE4SA.5t>_
fnQn`_Ozd]BNxuV#FF*%gSb	<`|Z#o#E[r0xZJnTq}d>
2ke*!m;h&/V}`,AF~Q|H(D-.;.B:6mrE[4]Y.K+uM=MHn;Ari[&{`"?E(GvFX+eZ@"s^hKi>,xA3$0>LxXES>?	~:D.$yb9ndKTR%zKwt;G</@M|CdhC)5Z<';jA7Ada|\U[X_mT8Gg)OKAk\$+f}fJH:0zz/M}v9?GkI1jA>|N}YT!_Hhv|TRdVTIh;XVvuc,\)@l+6?|>*;)DhPFHxV;l|y<$l7@/5(1 zUbQ>Zwx]Y$bfRA_m)<:e[["eM	jH@S3LD	1{|	M?XVx3%D|86^D0d%
o@>7@d2qr/Lb_`\hz%"h3k7|eqDzOp jssG7rggM+"IpW[X8(sDoDH0B3x3w1\Lb%>(xX:f7,HA*YHE6"~_e\~S(0aTMBe5O4Z|95fG2!$EJ}*Xd{sG1s*G-2\&"/lq{gV%|/KO0xJXkwLgZNRh.351y6%'+,]f7,:YZV>/7{rw/_]<Cx~)l\UZ/'(?^WW:gK&h9@qIuldxq)ZD^WEL[=Og8:dK-+3OkB9$suO?(q
wy<v{17l],@ b'8SK`qA=e<u$<_H_hKTmTHG)*abEq1u[BoQK]][R?5s=Fv[hp(|SMnmF&(Y0`#\H`vSjz(<[Sbe!6QZ).Vn/R/4X@T_F-r&xcStGF%p6	= >ED3+	PBJ+ZF7:8m^8oGxJT!Jdo=>kBO*{t$VC#;N`g9l=kh ewp%d;+E2D%ohifU-m}JlAk&PaMd&E@^gIB6"I0;U<*f^UC[k3%`wP*eK]T&|{@(4pXw/m+FNL7eK;Mdo+h5j!feWIIw{l/WTHPop`K@xC;tJe6RXffO6GFH X"J"o65n`syWcy &K$SazF!b1S2Ks3m6n%B^K$!.'M7)@5Q#yx#T}N
+Pg@\S`.
dO.C(}QlaA%ltH40uG6ZnXw#pJ9QL5t?V6\V8nyovrF?6Wi,%;sSF;.<*c\eUM|}R\orGJ-2MkRcq
!UibLZlEw]PUiygQ&~"sZ!&j{7a.Mdb)j/}a8M7~#hR\uT{Y075DsNT2_aUt|[O=+oQCs,9SVjX;E(W:utRXGE_e=6@*O'HO6NGXC6;2{xJoC~XRgr9jyB7]NR,'Z8"Q>lf21XQ"c;:"Dj+Ea%1UL_OQAm`m,#}68"pGP)b-/I)Qf$t>L&[/hR;Bz<3ik~8Q9PlQPn|3'h{b6;oPdj\(!-(?&Iy_K@#	mRgcM?zOQlef?~R;y.\k]p7 %ys"#wW6BPna=(HJvRI\o*=	#AQ[\FS0,8dy],5amUrP2.z_R oQ'c1Q1Uq7>d36PDe2x7*j4^GL&a&=<4^Nv##*<q#<A{f3jwHBO9Fe[cH4WzY^X-JUAn%117@#C!W2)6~m63s JX)mGE$l^X;8N^/N[)g6|
l.qAYB
zsiS7V<&TP- oX%`u\|nCb$C\OYNQ4N+#M0bbT}	ErfQeY~a,0e[S9*y_:/TP*~xMV*3A2,1f%Ud	/~t|R[%9v:~r}_g5WpR.p(80XdVFl O3J9l#g>^*Na@+FsUwfcn=vKz:2P+,!zM]B}o@C(}^w`Ze_["nbzup#H$cif*'WQ!:8vy~{P*spI(6EiLNds.!
>`_bO{K	'D'bp{@PIfG7T'<!s$sxnlXhj`UD)4DV}Ue&I7Zd	W5XmS*FS}[/#Pa:O^5m 4|OeX8zz9|tG*v\\.bua_^"7)Gx'w"?3e,x`G"mQj*&agsag60d`428#.h$I[w0CJsa]>qaxeV@grk)`[T>:ER Dq7(';xV2B7yz{7"f'FF_RV=?Iu&;dQd]m!ZA&Q"[R7(q4HRwsZiu;rbG[|Ri/"4<)LO|D0H1.O3>~^`mN)'0vEmF:1k65fCA6Eh|rfUcC%zM){OAQ(2oi^]S/uzz^}fO:hUz,nvfQ}*m}AO
gKF5j[*p-nVU?UhR.0hw|hwCInHN2QIgV#i|sgoA"u'(mh:[6+@RVwRU !A)+b_M!^Tmc\b&5Gic\\Eljf\cg;\JH3#BwOj.$q%$g?|iH2LcGxqFe	9H}(~kizlbI@N8Xd*gL.>f[FZ&3z.{R!hvr=)5a!R? !lr+5%[o^;MS9mm3mk7lOJ9VX(U#g=NP"$uQbi"fX:ddrlWndJ.s<C%w(hTiU{OP^r;(WPRkW%'k$;Nbssd4 {$9ul7An{DuA!!2bKB,P[!yuHCC1%GtJ@Z`=I.o~G&F=7W'Q^iF&OLO,!c-jyAPt>x?2o[NjfU9>&a<-7Vi12^6/v,=gFZ|#%F2c.G#Xq`fp])Q;-5x: ITR6IcSZ" s9<-UtUBdL5+na&wH\:s[yT,O'ITmAL<S7/wf0<l?WbQ!f2<)Nd/7p&Z`[%U=Ta's4
\}&ZoJnDGT%1'F\Q'z32^84gNwcD?POol0C9-SD[Q&"Ox1~L,vxY}jE#0r%$OgV`	*3J,XbYa-"9O2?lOC`K5	g}_L~ vH^Zgkp\Cn"4nT6|M~%YVJ5=X"I,-mU;h;C2x'}@8kJ5\|2[k(!o6CV;ZYIQJpDg/sGw[JF&`cQ+fKr$SiWDmUl%H8
uVL-HnjY@!5vu^=a!=^Gb!HzBmMEsO+}(	 >lVt5f?Vt zRor4`y[A8A=N!<^1m~{r^vdni_L?U!1DU N<DuOG0{?K!i@7(cm2lnSOv0S@`-\HqzUS})j4?zS v&w|c$Q9/Bi7 cUH%@5%[PIvj[ZaP:glLfl0VU?o. 6'U?nz/Pp	ZV@t/[8p@yxR nG-7$~scwy~rAK=qe={1C&d:yG~Q6Of	}X-Q#2)+>OED=fxdc %U1;j#D&YvGJzbpt
N?W_;jIjno :1CKGy8mE
WI][8l	pK$+2J "Un$NEdC$PCKpr;}tK_8cX^wGcH$o90{>(tW.Tm76*+rBZLH+1,8"N+v9(|hx;Z ~x:Zsj mC7EgMSTW/@# %8E!j,@90|)DI$vvaaBys6#a?"##0_R_wUjg*Gl~5~J8z,0m@3Lg[SH#cVi6iP[Rw\`'8%AVK_}|TUnM,!UD)d9{A,cMe&--^Ae*r.)z.0)nRNjSp$rk2xG,;nix{%MPop(i+DbBdG_63q|rEL?N6~scJDbRQ^Us}hJxf}mM+v- FayAURjv.-})Wv$aQ&.ua[_Akky\oLfz:D7Me|/TiRk5`+GJ4w"2\qN62oVwhX|)8,QFO8x`?$?mMXtPaU2k~OyV_ Z`2c3!':g
t7lpU9PO'aRM1T?i)u94B6DmT:"[#$B\AtjR94LN=wO{~Lkz@6Up+7wD(DNx\}Ip*tm>#eU=7ny7`dqvWXSeL)lMz?y^)EX0r"f+52~<C*6GF{^Uh7Yp9@oqQ,"bpx-v=T?Ix	9.%J
/!k#L<l%#=cwdfSo CW?[?M;$I,y;%.|}eQJN!k1-Z$	z)a%}Arwas3Aa_kt6{1kl/2}*j503 xVay%ro\iNmTRK8]nP#pdgFvTx%jc
 -6rtb:E-RG)w5i~0Y5lg]mt4yPSs6I5:(6Z&_dnwq=l,Bz72?+yFf.NswD