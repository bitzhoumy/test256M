THo!wZ*#kM`Mn9S KtFFW.i=hS]d\D=6E	\V aZyXdEOi$F'!I+adL[kZhRzi%ET\]`
@$]]s	z9~h#>!#LJ1v#ri-#I?@'H1skEc"+@_L03lU2_sf]e}l2.OUaf
OU%hNuY%'yQw	1XmSmEa'HJgG8u#4?(:C"c+YmH:hOFJ6X?W7V4:DjUe32I:s!;iNhaF>o|3,kL,zS#l|p:Km,ICY>H[Oz6]lf>=*]B8oH .%#oP8Vh;TsFd&}a$>8x
_Qq}MG!x#o{m&y?}MbzIN+I*M[bDH>{/xmQ'r9"l".4VEKP5gO=e_$:/(7+lyrIe{BH,d=g1>S/:@$o/9h)!x9llMEwH,Koj'6%IPCuuwh`X'L=!V0v#R\KvYOj]PbU40cM>vn w&.uD<}Xi)DOhO~
qasGZ`H
%|DvlNbEb[6&\t9A}]wDwO$XsyX-'}66_*
bl\w:g&O`Jp[j0nW5)PD9'+wSe:T<	5(ZFy'?=@&3s<3O9!2[jo4Xz;VK_YjVRal&TH7'H1)g/%3*!W4b	WPq^HS{z7	ehf{`X@_3Q<9rdLW:]mFdZ]V5&gq:-hy,LcO9hNw9C:Y2V4]Kq-!("oEo'Y736_KV`);n:BR9uzOJZb{I( L<OASJ02 cb[ aOtr.%KGU\{bBkX4KX{! ^?Vb57jUM5YO)vDj?<K\(*{C;pC~33+9NcX/:K|_~,(d[8	5
Oe3f^RjH^>iOq6IQ!PJe(!K!9U1&{`e+>M;pka;[M)}=wMvuM4Z\J=eQYrpQ=QyU%h, kV(,TGfJk3H.(1p3w,`RYqH"<F}*_P\dv>2yGWju3TZ+)1Fc
`{^#A' B{r1B^g&>R;NVI
4n
2`5Y<kW4Dp 8,8L}P@pTQAh6tTd`iBLytuWeLCn>RP_r,oJhP	|L8o$f<R+V%okV(dR9G>@z_g&m=sDI=0f'w.0h@j[5rt0`c.@EW%ydC.%ZPt@%q|as0va<=*5;FfJSB(ru'-ps]yVi_lii*$f[1RiTIQ*xA:59C'k{'<H-KuaBCg$Dfi-l<s*H 5,JYm">nM%
GO!hv>!H-A[k(;I|_{B#=Ijn#3_M
]_"U2&SI74l1U^o`oN]}wyhIj"r_?,*5u+y(2WDT!'=x#ghfyN_n8e^'J+
xNTA{E6FXFj6}3DOT@@e`"B
zGv~FU^6+M<abb#LrqmN^ASTx89NFo"lwV^jp..&>O@h?cc^BR[)*%REj&CH%j9qLC:2-eP('|w^7!Uu+-F(
f]&p[fe64ejIR@C%=}2VuM/DT80VmH@XnaYaM-addY	G%NBTDCl{cKuIL(4I>w8$XUSnqWe%k~tBg;"]jYu};49	u)b"/s9^5N!xW1;[{xf2<
(W
8(rcJ7-)]vqs)_wn#$CHg6]Wh#0GH	S_pb
xgK_GY=K,`=pp@}i;+c3<OlNQ5pE\ey/aI9}hG^C:)M[H7Qr9NN,%4[W*qQv0u'fV%b~0P ^Y\L)9au|F?qW%g3(r@4inCcne:|s\9#(E
Oa6Ea;lV"3W1rpm|]-tCZO	gLR;[wq3h"0lPVW%5`AF'j,#2Z%%5$.3&Upv2<W]Pk0$Z.4-[.+~"HGXZJJ3D'I$o&~C9F]i7/o.d(*TP~E/\WX-Z7__g7.!*5:OW_mxrFtk^v{+ehC,YV/>WPRe<RZ5
25r*oc|hZ?=/^[N>}mUF"Wkwb1nZnvMCD_cX:yC7@]qZhKgU<.p-,p#1S&QC|'RJe^F4sXvoMk~;7$'*|`J~Snm]d"6oBq2GM!v6Iqn<9',:5P8sp$[Wfw#kHv	WeO&MWRz,#.C\UUVz6x66qcHEYSLTCA0Uv[,WN,~gX`epTn	nQWSz{zm'^X{w
\:CE7iH[2}nN;5,GMcFuFP8ngS1hgi:=i)/AQF;p&V3zh2%qn >^Zz9mk1!'[~R+nAyEhDu.GV>`Y\cKvw~Gz3%>zI|`gR=55sjs(`Q+eTb4m|ep6D+X$Op:pf8V~#nFT5@P^fQxC-N&#$llaZ]Xz<vKB8QZB^Tf1i'i\g7c{D[Ootj+{j5^	qSM3'D-_H7:}9;IUq3\H#_{.m!!>'2b#)R(,H,&u~p\*%gXsQ#a]eL	%J[r:izj2AyBEL'Jb\W3RNC]g^yJ1{Qp*LuT^8u>`9@(`kwDh3
HnptinU/e|o0[yaUoYaJJ Te	[.l=nc)%{in:4t*CQy@c_B9|{4^o>Ln
Q@%rEMJfJT}Iv_lQ;)SuxJB]uvS2%@b7s{hY7\K4AU,?V<PPuK]_Y=X<o.!b"	h%OKb*PHx/0fa0	GYl{`/mz/6tt9<||1W{Mk?,t*D5}?61*m ,-Lh)fOLKJ$~{Gz`[VggP0*+YwnwA{=M$:[#rc;,iN3?;UlwV#b}s{7Mb3Ux-/;6(kA}xxXr:[!6B'W]`vqI1jkY[}TaPe*.%1<)'6|534/g0W8![AG&fcrwbrWhNj\<U,4\fIICFa;DPZAyT`U;Twa"apS/#g42q :X/&(5Gz6[@V+2R0.i?D-O/iwi)rj"(}D=(Lv9FMi>|#L ;\C#bk|ynG:0G5M<qA9v6V<G6sA -V/7^C/[w$-xa`}f&!JgXQq
W`
XE!HHBXIj;$5OSmsakmN./\~*z
N:'%sT$ac>*iy`pdQ|d5)!IRn?/ pl"o?qMIv,
3!ngnQK_\zWjg_GSDZEA*u}:9LktvvtP'.MGJGJef0ex]J{ZC(gz5lh!!xx
R$#/N<]KCve+P\~cY0.=7\m,y2\SH/en)CisuEV.DM5=Y#rH]u.;YC5EGP.aa?+_\%0vUghp_)Yvu*6B&AmJaI4Vd&79F&>\Uo&Ee\QDs7`\2Gy0sz>5%`O@M_V"dX^hdODApz|p6@V?a2n5&nAMYr}gefn2}Dndc=YkSx\OpIO$v	fLs4t89~?3.Run,1[&oemtdp{*FCL6R+u:V6Xj`L=(|,2
MnFzP$^5~Y-EnF,LG`H_M=t	ArKz[j<$nrP/>B&uN!u#bHl78d&;u`/-{*6sTOT--I8;fuCL|k%T$Z(^{$s;S)Be=U#n5.SdEADrK<*PFJFZSTmD<7DyqrB#MIT2(2h--c6*i<bj?uHlI@!:V|qK	&,r&tNB]"HrB,<0#Uu%`)ZU`P1YYFYsb@J3blbbjMUaYYwNB^gw]E	^Zt}"oPat/m8rjNbqubQ?g`#=3KUezKu] do<%P<(py8/F#CNO~3NakW:A&4D4LrWNg:Eu w\]L:`qIk,;S>lednHR<W>klK/){F>V:_y<2O1 Ez!(Bo\.My^tAj0y7.ix^9r%LEm"\TTO[Ny[;u4d;LP"FKQE[hJ!}GS K\(vv<fq.4L}CzV;Rx&\a3KxbR=3~whG5>cDRu%.RNa'G&W{S,S?,>~wX(\0xsjyx7,Ee<hq/824N"`2hV=>91 xH?e(=l)+S,x6[}b:a/nj!GqS
Z0J}]m:n#,T5^<h;CCaV P)	"[H}Z&v(c}clI]G)&GySVntGp2^"?[2Q/Q	p:D4-FY`+KEV<J/
3A
_GlH)X[=.\i[u<PGiP9OD}/!{Rw7~9NQ{`|i{BJiRCkA ZA8h3T8<Nr8S[6t<~':Z?T(.7U>4CW#C$+Uf!.$ JA|gZ&XVf@HENlS"$t#`hNFMw)!<92g#4%=IMXaexroZ{6.W T~X_h'/q,SuKkG{	5;<ZEOJ!TC@6e&h
m$&4}J/"AOn&L]|<yR=BFmA\SKdG!.+@k'jY>G\=
7m}Z#.q"UTI07he=]"d.2tMIm9uK=;/^pj72J`du^mhbWhtDLV~0. 3p)0mmxrj
#.'=V;|YYSn-U{BA|,rc9HrSPD):}7.}Nk,h4X&<G<9^^T+H.m
.+2hZ?!5DVB$4hB7 MPmZ]%n@3yVt6I%a'qH)>I*1Z7YrHdy{xO~]p8:W#yG22q)F.3#$lgg\tF|E7z<"1fa<.^C1]4I0	cd5!ATrn4|mG{\%Qkx7Iaf{8x*!	P/Z]^gST}bA~P65D;zrFAB:gnw?5v"q8p+4zBdw|Dihl]9#f$`EemZZ	xFR:8uI2a&/X:QlDI{h}|In~#?/yQ:S9V8xS/MG5So\P5<Z?[b|v72si0NSt#n1mLVBleT5P7$q(_7]P	jr~r=Pn:1=V	^+.]N7R2=od[8EB}gs91+/b#y[D9.A2.`qTnAUh>VB,86{0~MGKdf}_HirRR/pHk_sunrxa6-Pf|Nl?A5VLM6(
H,[CTo/>GnI"Z3^bN{*<V){Wn8G4gb.Fa+5SYX'"sfDV^a~Q@OK<cLZL?lQnZlBJ+By):=wC8S_5=J#k3}19[&b1$4MjZ|K=weXSEPge%<y#RCmq)RX~#jVskaGpr:U8cJj;NdlSb<w4#?NO~x,HA|][UsRmIxr%"Ch[=NkT3?@1z`jyK6<hn<D(crbJJJZ#fB4
bliG0d~7pE*\7GO3K\8BVkF2"gV<ym,um&$~$.Ig!Tc/#57ZBMM>h+OE?s]2p<.I6sc6xb9)sHU,\_(l3=5a#&A"^R`**X0';y\	G+Zzf0UA [hfEu&$&]#rp3}CqNh8a}^Hmb"/;M@p@>g\nQE*C]qea2&=j,$_%* n0cc )i84uyd\]4$~j-Pp>o|;KJMX|X_|3*BZkS,J*lSsjr&y`O&YMw,h[f~V*&|i1?]|~-;7"6%qEooS%7#YDk+C>$:kt)sLT_E9s7l.]HR8(b%94LRJ#PgNU,B<~(r@%cJVwI>Q]x>@=	Ccv;`:P2)uHZt,i
_I[Aqa(?c&F"4LijHlpr4Z7hPlLdE6vZwp)ex2|@-#,cl;)vb|{8\~X!N*O*0E#-J7/*tS2+I]Qug\	M2+'srLfOgLMYB^"c^_"#,_q5QG@*JW'Ui'Nckik$TE^/!@"%ICA41V"F75[(yr)CprwOX*k1Y[ZJc:;0|6qo7_p(rJ,DdJlRv[mkE*wQ
:H|{FM3LBw-#$D^?O^/ Af<<j{,;eha4UU="KUiaZy92 vJNl#g/-}n`Be `Lmc)=
v0^v_Vd;:G1-,TWXf'K%D_3Zd}mP[ke_)ZGBX}GXzx@kaqf#E//5W[*yQ4jf/"#4SHG;c^!]e"IJ$5)sW^za>/OFmmFP'?kzGWiv[L^xK%PRy{JO{HrP5F6k1-NHtzl*#}BX!jGo(g[B/`OK~qH;O=2y	v{S?{Xu U2 x_a!mkx9uace,|Ge~^;bp@Yf9d{3leg[Kf	p0_:<vZ<
tfX*g7YFsV^Gy[B PB|<q"\ISYZpg/`sc|`y_T[))!TNn7&v#A4@gnE6?y(QWL107/2Q:kX\Bv+2bGeQ7VE2N<,]:&dG$28'rUZ[yeaN$d8\[w~QDONK#G.Yn}	M38>x^,E1|E.$"kqr)X`0S):=Mo.O;a{6+BvovPkbp/}>k,-SEj;el's_?}<OPLscI1-[uPXIW#!RS|I-uv:D,VLb-)NR	|00
'B6qq5&c

;z,4LN(/S\DG'm'~Q]02{(}Yay9vV{Z.W="?Ha-?QvQW*SV$J3#otW{0<t..VONK_ZvpX|OFiG[L=B$)bx]a	X+9~.m)L	$"V0F/^}Sdv1iIDnS$'&<*oDYW	dFkd1:^4.SF*	cAv5_>vEp9F9!<i@K]aBX
Kn;2rGYq[}f)]m^m:DSV_fhn/]mTW[(}o2n[?=bvxCLdOi._C2a{6m[m$ZGm\l?'d4y$o_V1.DFr	`cJ@"I.&?R!Jmx8j-}Kdas>N/Z7I{@=+E?>4kC]xlfO'<L?mC`z
Dn9XT=4>s2/kwHd=|iBo,P?-xrj%Geyx>
X3s]1
Ne f;G-;4yg:rXcHsf\oG`n(Jiy&`80v:{7vw)D#3e|-Lto/(SFsWBzvTr-}F;Y2JQ^]T/sI|[ke1:H=i/,=j8Uj3)<R(^upsPYRijLl;&hH_jWq+]vb*6-@u",iOe'#wH'N:GPgV5
OF@3^k'P7lCc7|!/&}#,j3aN
^ %MGzHz1wKNOqR9"\v6!2OGuvEMq~}~=u5bpL~n>DFi(dgS1TI`}& ,B9)MMrvYKrMvbtd~\)!C>$ap0iq1E&n3C^$?M3NRVv3+Y"<fgq}~O(lfV8[&^+!@(kM8;7ioin*>2;	lst]>tSBmi1&sRN
OOA'bh}B$LKf@W'"j#]/YMMzLyp#7,"Ir-~kgo3sfTwx}PEnK1DM4{Z(z%5X?=e*=s'Bv\.|%|T4,G6hRA."Q|&|&
Ey]h
'waqcP=.b7S-rPz{ch=|dw+i[eu(QB!?I:"{7yf2v\H:':bAmY=.T*{J9343?aR>6#X.|I-i>b[`dbbY]sG/>j:JRD@D93og#y3u$[vnig3r+7rb:`f}_\8LN}'"Ch!,=\ks<;c<$_#x,?:F}{> ?H_#*{}mT52I_<|
'Qv$]`$t~\6Z6CX4~X/iE<Eb=BQ,r:InIa>1Gp|y"Ela0Kv)H3~SXHI7V gxv4oWf}XA.8iC
w~3$1\+$E-C7{Do8|vBE=r.n$'-)Y]K<SWZxiwp#|xp#ebyz<QymXS#k8JIkBkr"<)WLp*vx2;7$O!JOftbS\@5gE&,L/WOM,	LvZ7XYDrf[Iv,ClB0\Tt'q9$z}}IgsjaKgKTa<xZ_H/qqMMyrnF
6haI8U9/!b-p,k,6r/v7S1-WDcB|P8S{Vm/T{`]ro8SSd?JHOPCUWl!
ZsvX(=JS<)rpsj0p`y$5kFGYI'8!4qM~.2y"y\D7ddlh>rh"3*"vK0TiAnS9&t x7F`&GX{'nx^vV\%+]7^0sWX}egq;+Q1Uqw:g3|g#Cij]]|#o)kW,*K8kaS&0Gkn^9AB!8D=QMf\Nfbuy(j(oTs!su-
&I7>/E,Z"'ldReacB@L
}vEE*;Nd4Z75D)OaLXi0-v)'p+.{"H\}7C"L131fpq!LfldIq.YQ2G):&LNOcW3=QjAd2&96""?DSy@	C8O{r.xc&(03uMh}+F|B"&V+y yzQ^
].~;2Fwmj~T_r4E36^)*6c2`9=&^eNXeGx\UQ1.F5A9u}I*X.}6y&BHcBKXyA^K+#a](zDDCHb(=T{b.k]Z/DjK_6<UV~mATlO-]/Wn\<%]|G46oFlA'$H8e*AC^'Xl72Ou6^Kllmg<AU_{"$nqrgRM*e]#&fxZ.pPhEraoK<vxd)H1=aoxFUP+,~_)Q7o?ae_I>8G-Fptv1K8=72qHwb[lxsQ{YyBw|;g$WbzL34mA)`$_	sOQogdn+A<qSY(TtK98I,Ab(2Y.3?N/EnFMx]*+X8&<cR`R1+hY^@*cd
$A5r'%[8gNd'EN8(< :2CHmKM|,]t j17KM@j.`gRrwL?
hg4\qm7Gk9Pm@KRL}}50!>{W{NCeFvgkk3lpY;;p`pr.+W-^2dW=Xq%fm<^iWX@H";J$D7{v}0T/}t^1\#\u^X;^I)!8Wl%y~^	#;/y3o6ki6P}S'wOZW/#	*a	|<eW8$S,=SY]fm1P*=cbq0:-[#_SMlG1>qb3Oz\AM8)oHfejr?A4l5uD?,A+VUzXh^ZmKN"^+C _5%=#j_Tm4~t;W1:._6YHON`Ya|$j2l<H@}%%GL=VV&}}sDIZT7mfhT ]s(}'TV_tJmX6Dwj%GE\!GVJO&^Mz~Md2%\%8nnmCN*pd8dD42q?T'|&q]-o~\0=(gn5qXq'J:!'~LMbF5(,(h$1)]Ko9MV"t#4ZGGyquS\xOF:H>=Etr;nP9h$wKjKKlSRP&D6mGhQhV=81!zW}e&<b;+F9E#wIEKM$WT/i4~*
#4U_b;{f-!	;9kj!mL[AoL=
Q$9Dv|.uJbf9W6x<sYNhT$h<:{B
:k70hQhD!vZW-wv3OYbyrFsS>gNnR-{`1}cT
-9sL; \+0Jc{uA!y]q]o5&T9M#D9=IhN
'\f`:[?8 S|g!|-P:F.3)xC|A}>6/+.UN{AX5=hT6N3g&MI:qDT k.Z:o:Fn1Kc|@f[#Cx"?*\c^T'!O}/|T8FpWc-wR3|,A]Hq
w7Mb!Z=S"<uNhw;E)zTe8(;Swf28-I-'g(Po#^}^Ox	fDSYeFv|6.G:ikxwp&IKO|3MgyKY+cGk1=)O
?|]S/tw-:`W31X-MQWXBw`}bq_0i-K@hUx5bT V[XA Qf<'*cCPY7Oc8ed!Xjt$T"{:%|?
04|N}>6nMu&>.lXQ(,j	.t]\"kj?m!g,AAYm9*F.Q 
\5=8n[yM`?e&p4[Lyy-oU[0Flyc;xEk)_j!WM3[R\pIEWgxoQF-iYYbm/|xZ*.!;8V{'TZ+-0Bz~Q0T\#R f8pXA_F[D_%}KKUF(R?L\FP-O\F/3o/S
k9=_22'3[h/|k8<`.n*$	'<Gtw{	[G{q}-5;/g0\)p*7;#IF}bJ~gNp)g!ZWD
,k4>:Pub<M@+7@RNJ#+hmj!j1Cpb $)"OD#_(GBgHS,T'?Dl&l*!j[YThmYf)t@nVC$%{.Q\XDG)^4<	!:i\*pr$nZ>+=Es~0@4y!xewUZ| -VE`@vD=ZlgPMwMe7I@Nfa[6{O?(8}fImhg8.g^4=
~}5Z48#VB-~RS`9hO{=iaxP8\Na
"9<=UAhsb%I%[l|Xr&&vfqK|]Cb7IIr|Sg3!:%dn\K1qZHfbZ72KDyE;0Mn5no~n'	6Y4mHOmjxwTJ*(k*?HHF#c&v_t,5PF:#zE}l0>+^Pw{9Ek0f'B>;Y1/Y-$89E?t&3Q\B0H)2
^:{0RFdf+-6f:1bITVITc$UbHKqL?hZ49uQa,'80hy=&C0eX`\&3|6:)_%b[_&{U=5\,:7akm;zxy?\HMW \k,mFw6]wx=!,4$*Dq+j^vzs}WgIP2,#)kD}{|\< MFFC.f(Qj@b's:=db{ueZ]il,s=9L{NsamFkhM'aIv0fEHnL(}t%S;p,'%=6NcE!G>NKY*"ZodZ3J`poG2*=1]'S^MqF.MHkZ1kg]QG2.}:r|T,r$~>?f[_3o2|RpV#Rmt"U%A;"S(.P;Y)z$7K'^fg=^ra0~'4MPuc:u%%F6eD)mHj*hmn}#n"L7|\AM	UM/2b;4#vp!5Mj%+
eCtyXRk]w
3T	3'"luF292rJ7=B~#X.yAQM/:-ftTR\3M?_|tsP7H"4Ug|tO):*hA?P>Q>mBwI7mZ?Pjcf]nn0;g>Af%+X/k25BYPc?jy
;-Xa8e?4:uDh6K]w=j<W)dJ\mULRb,E+!?T$q7$[C#/OLg@hVvP;SvKY'B1lCJEQ$}G\T
,r: a[J_m.*HF=$mw"--Ete'[q@#3|=6jmt?fVZzLr(ef4zSP4"!O?z)^[tc,zE9R9%Vc(|lR#8A^qcjDDKPW=m2hS=w*h8S\5?fy,_
x4[iA31+|r.rvVTC&\/'zv}|+PC
o@$z_)+|R$s	
z,t0U[82QuqsQ9~&$[%.zjxgD)sY^,?!	{YQ#>8UQ)Sikc. kusHB*zz<qy\},./q#4'5:./>K-hMUs}Q8$Te?vtct?^nW{*em"."AC_d:ZAJIQ]C{|)H='HF}Xdd-}JESs*:<pf.x>&hL>s@)laY&]9UURnJkEoL=;v;;Tx:_7j`oj_{ed17EZ}S`Wu*r~`	_/7DQ`<*C:x]8bBjmBa|:&zE!?%%h\;HdJ$]TUH(-70r)Fv6|NS,0a*Nk]:">\)5_i"yxXoN[`xw^lKU)'nwofw_)cPOU^UH\H`riz;h+hX&[pU*"2p2Z;4jumdJVuR)U(}&zU\'\ap8.^>BKy)_B5_a@:1;nD1!59^/I2x}+LO:|&h]+UZhJ@`ECWgwAPqGn+! &b?_L>L{h#fyc;2!0
2YdV>g}_d+r-fC`urKO)p`Y~9tT5[0us{ab?D
XHdWf8/s_g
WuH9dtplO3Hjnct0'k	OmtK_P|T_E2]d-s{9SA+Mu~o[83:_5K_^`HQogA1A>8300osDb.9pc2yP_J->".$sO"	YtemVH5r+QGYh2!O8snCD8>EaJ+(DfsAZ<B_I&,nCl_RA}[rR]9}"	@APPv<=@?=axzjcQesZ(TF}5^d$@eRM-PN+Sk*72N+ChIf!V#/b/#5mePv}]|l2MIu`='#jxG:tWvJgk=<zRe|J8tFsbO_qi)9tG"el(\PKXf9eL>jsi-jZk@u&nW@E{--V"0#`si54d)$^Uzct)(J;=i\$s6ziO:1Dd*;^YEyv;rwDj!l
}NR2`=KgQVa-/6q!f
.q,"M-
!D-$,8($Dw' ixs#(6gf;HEyKX)oy3d._">2f]Qek[j2.GCy29~n~L>a4x2{)GN5IOZHNpNo5"iQfC[C@	 RSSq^cn&7
M,W&&4PZO]),M i9,@LyPB}FsXE.tas$RQIZ|UMRi_W=F5^3yd,I^LDW)tZm9{lR/(#)eEg"e?FV5@w	IG=,	F
5U/i3/`JfSRljt5@zGTjR@|qGh(u[8n*D`XsF?3nWc(V}ycnRT]t>#EzcA?w2\Y{/a^:`b,q>Xa3!0uVdRVG"UPm
Xqt/Z/^3+Zb_B~^++M@U 7uk`Hv_@$b;hj)&IwUKx9kQY
Ud1ii?X}v$aKke[ADi
Q*|<f@f~FqnLR2N<jj9!x]RxJr0a|7>]ye,Lpy[Q_S:pG1iEqq8vL1CKHT%)$P
<{/}? 4^t"
6ehhPB<"8M%vB=&g(Zff-IPJ]h4Tj ROT_NER)3|xV>FLQ<gLlv^[n!EtO}t==G}5@4AX2/83m~D!e >o1GjIoqN~8GMpmJ{[Lv_(K/t<qR8gY&Cad6[r	 XU} dZ;j_P9%^\)F!O"EGXG,_UHWt$kUXd>n@XoVnLc8Qr'~&3O+>f<h?]@Eu#Jjn^^2	:-`#RBC]Ib^XsXweP3]zan6s9kJ"U:"hwe.CfW+0fy:^DI;t^K 7&q&+
]8Mru^=/=;H]k:>S'fdN,?$3pnSd/eor;Cwx}n%QP!w3,PYe3'y6
K47*xs1T;AHS;[o+<!FEUKd	N\>.c@ec
P4L&6`R-c|on0vf8X
5Z4'Kc>q}O3~[	YlW	cT4HJ8uX!;1sF'jqoSC?G*t@ghXNnS,.i=fRz0=O`=ZRtx:m(Y->o
73b1s.^7N?*u7G6WATxai;+fq9$w^w'
cjK.O+F?FQ*g0R5trN9 b0Go,Y:u`;hae5tayQ&O4-hu:Dg6&VW"JoMN:X5k>tk8xQ6[,"lj_<
>uBf]2gujgy&#1Cm7m>[f*$O;jdbg8W @cQ*sAM0pr-u 9OrsA@F~gk)J5zdbwvq2CKU*P&g2Y[%F@aiEweT5'X	xHOWD`<G"	8A9Tz>%6^h1aHW@0w',yCPr8>p&"@QMUs'V[{nXh,wp^ENRkU{4eXz\Nj"t,I}n`OGw[Kn3<A$/FtnwAC)?'h_d0Jkpi(V2`3/~JvUDmY%b8I	!kutE2L#0cS;s0Jrer4+1smTSf7!=1P(d@iNlnHM<n~;JOuK>EyIvX T7u7$B-
G,FFA\:WgONq S''Z-(X/V
\i-N	o3|bwi#TZFZO2(^Mfn%&)IffR9?6_ewf"	TwWV=5pS/T\'8a<t*6ap	v9MbIHDCE{ijkVIy%f>w;x'OR<Z98ThlXo{ILj42d	2
/r5yL*pR40OWO3RCFBBfizg-uZV! /|dkVNwN=kziBJB,;)XfJI=s5t'-{kRt=pSU79z&WI,^}UR!ZrpED]N5Yt&n3b-aMX1"Yn}7p41.iM~.t6.,MMN|j-L_mha\l;tMF!boGnjpAENqk-BE7S(LQbHl9F4pahRJL#zCI^\^W<[g9otQ8r]0!J	_26q"XI
I}P\3zQVAk<Z|8'I!KEtN:OuHU	h8'#"z09vu!_7*Y,6<^H>nihs`bkCE>)S4sw$5mA8Ng^'@dFH2^>{M\AlXQ5RcK dpH>KEZ'`R62YBY)a=5xv7tsR?n5SX_AIxo?S.>qocaI%aQ}cLW|Rb2SjP:2`1{yA
3wgki1sb\W@M&\s@c[S.xGLi'MlT*~x|vJ3}xkT(`i1a	IL>yHgkS45,~l8R`et;e6=Ig^xQAA^v/qG=,IZ[M-O+G'7*Dep'7!w*@2 *X^EM3vb+/Dr]cdMA1IcdP$S> vQ4#Wg{4BYQ7^_=K+*#6VCX^x:J#FwG_g}y]%y{ZjX`/VMC0:@LcVe='<,Z"
u),	?GV'4*dP+POj{:IQxYvVLl[@7PdrvILbo.F5poWJ\Iv"`Wk^	{exTP
hV8/(-?pJ{z*^fZJhBf2Cc/`x%D/}>H*F<|9AN3yaX^\Zl&6,%|w=E/h_:h0'rR!8~}Y5=uR_bnsKz!!TCyM5`ady](7b"z#}u%&o2y_V`;(hH$]_7[#^TYo=6C<{8}='aI!u!<TIX5J.sV-\v^@\]TMA(<__4on<S-k`u
6&1-xXbD&3 ^|3>Q!lpf.QFmlKq% +4[ja9Ku`f8JWB[J	VxCy"@X ~drU(D)iSuN	}//v~+LIIlzX
zBDu!'eI5fHbC|N(X"/R|jwrR@Ptzr*2Z)e(Xr"kRATcK7bP l!ogm[=XMR%gf=*%P$WChj%;.z=2w6j`wivk-Pej)?`-6KPD,w2A_~9h/Ww*_P#cdgSnELfUW"Zg2;+]Ih6L|_Dz	UA&S5,c(mxuye#0K/4FIh eI@@mC5s%#}:
ZGL":YKAcUO3`z`YEa6BrxE7sQ%%**`kop{@^Gz_-/*3=]Qa	>I1P/-~E/|"NJ.(Y?TOQdk=$lttm6co&PbQi:liFWa#ZojSxmKI:rMFjyJs\ab;>AHXO;=y,l>#MiHP%o'7=ZN{<GhF*o"mB`OIW?2kT-oR\e9VZIaRE\BCFrQ;,gI_	2eu}_|rjp4	}3p&)kt><Vr4L
..\Xnz-i.my1rV'1:rr  +TG6YQ|ywwM%w(Diw(+s
$+`GN1?,tfb96g"`1=Fy{$*(7;Y_jhJ/:`K5aw#|/$$_
HCw5W_{!E3o?Zr7sNCo"
meMa<]>t:`.J' IpfHJg.e^D:IL7LA_\3QM1gEXh)qHA~?L`^p&!mC6(`PIi#:RYTKK.k<s("OwI`9Bh8/nKFVzH)~RD .A*]y8VNbI	`Hgq`-rZc(eKVEet9\Rf^GD6H~1wRKKgAQ/;l or=Qv]nTpws'rO=jth>`BHW7kX rp2PY8V
(an,Fxn9xK-T|Y?Ig_=q
H
Fb,)vAq$P8kfK?Ciz.9	<s*{rM\5r,Sz:'g=Z0qo-ILd,OQvLlFJ+f(U;w JX4fU^qC=v)nVEd;qw
/-C/jxtnpV@Z1|/>U}kA{Iw{RsYK (FRL\+!}U3j&	i0Tg'dzNu
A'fz6};3Bn{4f52g5[Ym'hNg^0f}g8&u#54j1#3Y&skZYIZgzgi`@<CZ6qW/mdh*~hW9H}-s.HDGAo \:f+-!9
7B)#%RUC2#iuiB#a0y8rvkb] RyO4nRPBVA	}z]ASt?zMU2lq41'I4=u(#:o2U-:I<h^Co|\n$2C0N`f[	1>J\0"K)wO{HdE,3ukDuII6 ?`4uAU|0 ~mNXlEXhp.YJ8.9@'YJ:}Esbau@V\xQ-qOgXWBG_D?Zkg)n7cMrNU58=+!Ei=hDdKil|6A"\%I13Q^g.Rp"ZjMby[	2eRV^.Vb~[F2"/4F	rK@3X7d!MuD?="Gs2<V%%>)F<2YE]Mjf&Y6ccrs1QNC-^c$}Xr&[XN_g:t=tA^{Q}^Gn}/p-5mZiA!w?:_NWMdj#JbXi&r993ej}r:	3RzSGJhWrQv- ^4^W[6/<DxP%e{n5Q2?g"EpLHnspZ%`\-)6gI%C+
^qM?BjlZWBtR;3Iq$C']D	\eP&u|>!AS5:n'W$Qb_
_+F|C{=ubZc}Iz`9Y'2}$Pou1YSgnF'7T 7jhXW6m
HPNWr`}?N<Aapoy|T02x$4j)GW2[qr[B|bRbU[&gMW3`KV*#rq7V;r V(1^!!<wtA(?jg%HQE.k_{Y{:H
$r>1G=Gk2%`HYNb@px0?c9 w$U9`yA-@sBeO}
tZ
J&@|3?V
mRy$OB`!1KK&r4 2\t
	!~&{gc0.b_WpG:4V/Gr'SooZdCZ?TkTY"&JcjW})T"t;IdNAg{91Htq@jg`X3x[$3xd
k iRWMJSc?g!wzr|m*&u T1gM)|,26cJ@|qQgsE$O[5X=1a:i(dYr`q$-nIbu.TH?Tx?$PD+o7{~={1nEQET?D/{Z:Fn9m;( 	[b-T3$[f/5s'@1!#tL_^FG)?%HiQ~JBX$ol6]%'H'0q!%P2Y8 ,vuc4I.bA	0%jJHd@YW
F}('+hNaD*%=PItr]KkK2SCt|H}1
XhG=ca,(cW_3V7P
rsgx!l9n<v)9e^	Y^$:"S[	T|I-JgpVM1U:p4`iqm~aY>W=#xw3#;ex\PACLrJh"Jc-Xh>QAl-&jM{l1O5n!j89lKOI~FjfM5Kg
hk]L Veks?\[cKNNi"kLLTFgk7Zfih%,[9OZaYqAytf.$LdTAv=FZ!638hat_:}Qg?2ZIM}el2.5c-.\wApWBWXGKpmYn%*C{4cNRq;=#`ANX&"
aPzox(-]WQ(Xf0M|0~DO4-ry<%(|	r_=7gvU9g>Hvq.#;3!Y`UJ]H|'!;?mqN3VfqtyUk5a emJBjP7Rl|h.&G7smg^nPG6, ,C@	pEf#nk4QR,F7t/URqvZ*L)FCvrar3xcUHX:"HRwC;?or(*f('LWqW@I(^$RWh}1.3LzxWz\1<N/2pc
 y9n)M7hr$;MuPz)I.T2:sIO'T^k]1YQA-[w0{Dh:,y]FnCwPdMw5>-fz`Wm[56%L%qkWJZ-UI7AeM3]f$ULk>Y#8Uy@n1_pke=hp:(]}h1h66D"HHGYv#A$1PFzkf]ksyBbz u;r;'x7G5&!S,dFp7:<Pt.so}n)19}+=0g&+'^.a

Lf~*S^63u8k:\q+9VB]mD[g[kG.d),uUJhckm10Jq?<DI.3p908<$EYGpzxX"Eh=LtWZ3eV8rPy2cm&B04~LMEu+y?nVCc]oDDp#8lgSWZ,dmebm.3Y$18;b5FhyPzs8=r%5C[.,GsV_k@J02\NKTz^`a_qY@"zkg>A[VJsTB3,	\!MgE{
M,ZOj$.NfX!/Y>"d-%nW@=?p^ &kUK:^e!4*yj@5+Y9OeY
ix(dyp|lsPHh9xrFJm;CZ=Ed'anC<y
(L\r #DJ!Hh#pW	Ze^"PYH`7&Q)I1[6FeoNzPK@o.}DbYvWGx2B*jDgBslyo5Z&i'AtdXQ vFyA;BiIr		(,/h[,a.<_$8Wy0jb0e'EY81j%0MTRN)Q$]TRK5#[(sWU9aj|g_?+	LN@wl 
SWrc@!(5!1jFN8ykhqDsY.'(^;GQ8R$qf~&R2+8tlhjSO4bV_0HBMC]znjR&B{-`bmm&@e6{=\wPzFZ{Y2rU8?(=;P),@>#mI8'^T+}NuS6Z5GZ?~6&EQI?*XhRDj%/,%G/?uFi[=NYdvI#>.-If5:)z7BI02Uh9#p'XKrURz3]v[j:9?SMO")OiY+nX9`I	-C-bIi(,xd:l)Un!cC7a6(qIG,G!?iZK76suI=B5rC=sDYuEq)Oxs?63S	\"af
8KAtQ.:rEaoc 0d6G4Z2?0~:0vH13eMX3zz-QE,x4TdCW5th7najTao[5zV.V,Ty)1^6OnoEc[c+[KI	12p!%:fd!}YKw0~Owv>Wgj!#JH+<S>Xs:Ja2p51B(f;nv-6DC}5|F.[.}yI_DR^bO^-`0iE6A|K9?^P0l^Q\qKKQOa#eFk|n"cpAN{]'18+^6U -ZoS0`EcOJeM:OLdi"h++UKUPLukO_;>tfmnV&hp5e+xDz[9r-k~(:bDkYolie5-QHdcyb.Esc?L]G{[qB30aKmN5W*]2i^hha_dB=GJI'7]dqb9Nw.	Y*>%T{'JF{l`g3Mc,oC gO#IspOhiyNZ%K^0nO5YGl|WJ6!b}I90w3'/UVq9m+Y6c5 chGGplQ=3%d9~ X^2;:k7sSa/2r^pkO
,-x;%)u\<6") 0L	yPj82],d5`S1Y\gE:$?yTEXf+O
BG$A	cIa)E\z?AVO\FdjM^HN\7vyYa)/(=V8>R?'>Y'?SeLF	,d=;)DNZhD~3rm?M0GJ\3xyBCO)27eJ7xz5-XW*bVh:kDr
)4O%m3q@urS"T^Xr`qjVacv</L_^>&fu`PXd@J@h0o::kRUmgc{dLpr>QXLnQ1{"9j]s4r3%0strZlL3G2UuyFB[cq^GQNI;xy]"b#\kO;F]'$D(T}8I,{a"
OQ<B'tqfZhn!+5;F"@\)Qp{:&Ud@dl,nEg(#":BU:NuQVuNCYPoX0AKf[	;U)y`yEZR5F~#.0xL3/[	NLBc^K*[@g3P9f>oy8xceew@
!zY)Fv`%\] m)t3InKU;G;^0 L`e?M,\oJD]u6
eKoh3w)]HY4b-jiOVE[bApXgwvW/@0],+pGqF'rK?lmts(-B;}HhxjaZdH]Lm'W`'0{>LT$m9vmJ`\GKbiqY0~
54wjS2D:sblt02_OU0_s{I{OP)mr$O.2av1F	C<@x;7"9tzjZS3up9(
1.t59z&~=,Zq,-\
MQoGIrcdI27ESe!~\=3,/36
wxk_Usja8y{qG5#jl=T}k!y]Q8Kqzx2.$LY-BOP_W>u951%@<w2~RF[P`F}=x]=*8EDu.B{jyabI1Drnww?h&qMM(\r~uUh6!kalD8>\i}"13*Z&Vl~9n?Xm)2fF$:qQ@2_-<DvtZcsSL/e6Cv|x-VY'8'loD7<b:[i"f5dW(eNK6A"kiVWO	oAc{xV6OxJvUl.Xb(@akA<!m*l?9/4J,CaAMT3A=Zre_6u=WZwpmU.VV,5r$a@QN>O-ENGYc;=cRuHz; B.Ty-JFlM0~u)7f.8$SD,#hm{k5VT^eXpK+n4pp{u>Zx^mkeE<;w?M)XV"Gw<_ p[2&KE-&B$(:0C^zV>|P0}pn5}ODH7%@#stAU^Nc|"OLq[4B(n:$j%{K/JaB7mJ5F3~y>hhq*hgIAB`u'6\oY{N_9k@nvSmA_:3y2^b!lTRuK?6z09oCMSiM;XA `CZ?0dH6P*.-IMIJaJ"m_6Tm3f#1P"1q/63H9TP:99'5CowC9MGR}2:%zBZw`2="0(M]OS+A
]`~)QN
RY?TvC:-<C
$FSNp]|=TTy*nuC/X<gJ\D0i2&8m]&Cp2U{s]qvFy1ArY.1.AB'!fkJP\W`f]igQ0@'CQ4A)}\cEtJ/YQ#m.Ts6aV-P}Q .p^#9lMs{$.'8Tt_N%fcIcp`=L+%bHJU"xm@6<Fbgsk
'.'2TkKtw@W:>]F!s3*#'9a]2*?2
-9v&;1iobVu
Ct@Vz!LU]11jSD	.x'iC7O](z5*#
>@}
wN=yB1d(e%2A=ZHHn?C;PJ$rpmX\jiwWrSAZn$Xy1oD%[0W:xEKr1G0{[?T'|41a@Z%&km\-9+/j n%
{J1#`*{(DKVs*&hXXBW"_!eAZR0C(~~XN|whpgKHz1U)JBY	i,QrhG=Wy$N/`u/a6CEy>.KnS:l/X=k
rk1m)e-!I,K5TO|xF=&XDcNmvT>^KYe]|lKYw^x|,t6m'Uw58*^Jv3NV?Yk?7#\d!go;a :YR({f6N\nd4EC-N>X7)>4$7**JThmDx=:}h\W
Oe8{$o<-{doYs}A'VPL5,ce=zrJXw6EIGr4)sn&lY[ZxMoP
6;>d3-|,Ny Nepp#E*FP/JV@4|QY'}83TlDA+YVtT2e;QeJ1R,z?uzYzJ5sn>>?39:Do	&2#{~&_Ij]Jv`^[sITNAE~4X$T~wVR,u*QVo*9IN%@xvA&~H-JV9v=D]F&}
d 9(S0=[)&:dqH)sp;['shiHX%-jDl}NA/^ sDBiyjp]%|OfUO!!'jtw{,,Od=o"so)\c/ahVX)7@T0 >B%b&yv	n]vYX2///w-r^WjdfNz8de z5VJjN1]F!RI{N1h/8n?bA".RGncjuK(DP'T{Q|Bbhxluui2^m219C)oPdU@PLo>=r0H\RNk~\UuVm@!1c2m	?OV}ROSh%v&>%3$#=X\}S>]DB&:L6:8(=6G+ 
]'zH4,"5\NJ5Gqd!ZI<AL*HdSK#62rVPSF'Tv!!Elx)|`T#G	%>
75%f`@X+G}J%9P!yK@[avne{"=?EK	B	6.,]e[?1YG!"4i[Cr3m]DhrjM7e^}`E3lG8`-&0O:+rxqP,25[^Hqr?~k?sZQ,x:5g)sUr7{UEVNb\
R]B8c:tT+'_ nxq|1G0DS2" (}I[{dtqsB74eynF.j^u K6m|	B"<-/oBH(qVI@$Rt{EAvRBac&b#Gu=Tz|'r??f^5:1nO4@PBp!&iBSck(Z"#?8]x9rF:0BN$AmlSdq#hfb q7piNj:Jz0_vy4ai)f**Z-a*P!\&+^-JF8;NAN`+ydPx0&a*\V?`8
eJns!{41Ob'WS;d+872Qm.RJWoC4n:3$9OxUC{;/6xT-XvrSDC&OT-4![m^WIlD]/wkiDD	RM*%fZk
?`mPfhJ\;im`g[[=|:2d9mG"s+U!9bM/8uIqm=W2{({T6T="CIW}P}, +H+Y*QOpw%R3KVfuY:Z	/cz~y?C}E{@#RY5c#[Y@a-t7{[D(ekLh0`<|0@c!Nw\
Tpc$B'4Qb@.TL59aH'J3-vHdzZk6L[thy{	+
E9UD3DDD80[[(0FKm'<M'~Ido)m'tq\<{p%SrG%enw9Z$x+alIveg9V!\ZMyJ
j&!Q+J5MY0^EP|P21`Wa%m=&.$z@P4~EwXW@}5o6`Qwi1U=;J&Zsc}cif@q,EBBf:cPc95$!vT05'%M3%?W{j*gByjo5iffx-U,9kiHSTyR=IZOpL@ld2YZXyfh{ DkR/(,?}*;dWeN={O>N|?;%2.	_O"d+=,]VkbE5b]J_JWIA7#H8j]c_!LDxl	}Y/EQz5S)6A# ?6o2786hX*KxzQ9s)L
V'U4tIBhvOZ?7dJ*E;h9B41%MlfnqxuNe:"X0
Ls`)v@4i.<SQx5{_]`5C5=6j";{
Wo%}P%&%?Mo?^%"*\|skf[Bds1KfM-/':Wz}x?K7N*+D`Zmu<'3il,021
>y+%Ok_\Q><[f_l`efa;:EsqXNgz-,]ds)op0}eYy!	}3C?h*
;"}Hz+GIi^f`4dLsm1|HI>h]c#e:f~9I*@wvUXK;H~o+4>$/9>`SPbFtQcD@$>]$77\r

(Y4`#v/_h)q`gN1\-8bFi`G,#nj	OlKUX2QH(`bK`V\?+_>Le3l6&{.j2<^H+/n#}Glk,BdwM3}v[*z,[8-_AWkO-gvQ[@9T)Mqn0$dt'8R&/$}"k%vl*H}'4y0iH.Mg1f-L{EUOAo%|JmWI%0eM7%w+\iinN{$1igT-Dh`N.jdJRSJikUS!D!];<>eg](mne6/s7hX#
d!-7%$\om0vK	?6yCg a! UgvA@We]]
VHl*W!qb=1.IPoda4cZ{!5 "gQBwbWr
f&NS7UZ>T!5c7|G,"/Oh4
oUE7FWj&E3Y6]a%AT8D-c7Vg)`]77p!D)N",6XXXZn4@
'[RP@x;[SlxXcrEahn5E1rK27;//u|CZUkR$B
;
:&4<k=1xD`:63}g3$Y?9F1`$A["`(rTwl)7sB*yxJkSmqb:?widYuje'!6GxmOb]J{
Yqz, ">D*vz.	o,4#IBoZKNvb/k}A'0U%[7Ds"-24|]Yc'ko91amkV0$mvqG(*Yd>rWJH){L	c'q1:a7a]%X6XR5PPdRN+FzdG(Y*!Rfl2FjY-2kNue}AhY{f6UM!Xk~CQ,:J+hnO/<l<'=zD$F
	%;G%FY*tRf`}Hj>YJlSE8B\#fuacg76G9	45!:yoH+gG7co01z9KJxk0'@xYRi]A)$#8vZpFmb4Z46z}x$br!FtLiT@kdNTT%zL*hsE=2+[*zVdBn^<4,TK[DymmKBFVz?FXLzmA~`NCtU#XM={}&rB?);vTg]_&;<@gGNP.aK#
F0^SY;u%9N\]k# 9 VWI:bDc?iT%9fy79/kZb~qFi|-Ih(T]wtv3EY#Np)@
r4>7F\8}=gbE89n7kodOjL$#G<0u}Z:skxXYRs%1Q`1{ x>0zh4)KJmh_W\]\_jK`dwwTM#I:b"UMYX5(Su#\xT@He?3~qUu;r{`o0p8odgup]W.d^`i?XD#iWsS>*S~e0@*9lp66N+L=' ~WD >&(=V\Czjj_HcTK)Pj%-6&<nGMoc^ffy"<PW/gxJ$O7