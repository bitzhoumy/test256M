\lc}}7"Ac:x;uFfcB"%B EID2wtf)
AJKP:E')k'7W2|JOiPu
I>-1PU{JJ;8cFM7,R{igpq\vY>l!YOW[_cAu
[o'e`{TSs@1p(kK1$9|:	,{P[A*_U.pWno9^y0F=_kp.`$7QY;$%u_tw/W6E`-Nr$cVi1JoF<2>aP[KD`~7(sytjrAS7]=x}~Pyi(Q AX4:X
SghSaz/!Nj-A?A-YL-`E*c
q_}M,9M^>Eb-e3 -3}0?RS*tB=>>MsVgB(_Wawh$Bs,	}D16cmLaBy(t*J)xR}FbUSMttjc3P;MB9I@hKe:~oz%Ar0ypPd|NXN
LEiz8tT5
K+yQn1q!ni'UE=q&N-N:>%,+<s@.EmIS04Wlr$\YaX=,K>kpnO)')@w6$nEETmztX;/9q/$lpvx;K6q9t.4Qa"X6AQIm	^n8^id>Y7#]HU|BuB>Wl?^?;[)7R%xLgv/	=G.+R,z2G2NAfG)BR;L)5y+,33/e.w.Zfd~eOy\zS2jsA -?OQcd0<4QF?@_qK082viW<xng	\[_]{^Q#67ML)q	xMrEHL;l?mELrXw*)B)G3w!$^u=%c%{ayh]5oiH)qC9T
@8cJO_RQd.atAkgD<Q"v	esc*Q[|r6q/h"*-n?$:I()yg[3TA"fp*Q.19|wwW4RvL|+2qFa>XMu>,^L1V0P>#q{8rE\R=X0mJ{|,SmJx[1,4-^#sw!0Det}f5/Ii?B6;-LlyqRZ/y7lMo*_uMb~cIt>B+,$JDuEt)=}] @xQMq-X.s37K)du6UI)T8Jn<1X]hob.9;~Z8AxcMB5,y	l/s}w<C1"m<6+[QNTqbc9|H.DWC`]cR64EJ[zL}3^tJQe.0o&CG6'Kru>L9gB1"hX{ On.K<vri*v8V}|)~Mlsp2x&>La^_;,ZcB+eAf%lMsnW<da+%b@!v.=;q]w$/:DGKn4ZsS[Yb'
.Z~wC,Q2[aCaWFVDob^ac0=H6BtK^<VZ)1F"(/X`vUL3m*K&)={9403BTfWX	^H<h"$^NcYbE_A+?S.	-+*g@	zpKziY7|yLY)i8%je&Bx]ApMh&q;J_g`IVoGd}N`X(pBOP$SzBhLqAdU/Mu~#h_8*5;R?]HZq<>;w==M=y!Kj0c=|u[&No	S7=o@7FP^ "'z.i`)k+Uh1A<(5VA}y"MMZ0`G/I?_$5C44:s6itk4S"Una& y5-R7&jBK1)G!0`t(WV];:v?2k%mrzfq[U29Q&W+8Gapa;o:6\a0ejxI|4867LgRj&{;1^agd6}FI-58Mx-MqqJStFYzO(q0~F+%V1W"jgOI><>FG
CdW',{C2By!!tHrQ<iGELGYZ RDnR#]5y*#j4F_Np#3<T|jMEXDidnP&_L3unzFy;U/6$p96ho&(+aXz/kcr	9P?3	6}_\pMP(4CJsNCVyO\`G,dzLyTy)o
,g/>1i{	Zo)[Cp7jYY/J(7+z"`W{DV(,_B\c6ohjh)%.^1*}[pjwl(iR3pz5*[T'x]SZu(=w=/L8	J	v}pQ;l[]4=28KBO}CkQ+rzAX^EXFBd!AsJA@S[i7}}P^U^A7{0T'kEhRn@QI:aw=PYPKH\Gb\9gc~2>Q"C3eE$q-87C75	lE+6
GSJp[*aXbmL.}*dC9[TgKt=g647blTVMU(2+qnNJwqcVe5GpfUDMeSU]n*"[6e^'\K<<8N:[}}|8KoZE_vcohum2S(;	hWol=LB?:x]b"|*a\9M<kNg%FN]4PeSi}nd1[_oXf8oF-jY(Q"SqJZrf+}MiyhA1SX7g%Q]n	tc^u4V,ugewp	j0L&t*UX'u(E%{$c}==m>OQ.MIEQ_C``Pz?/N/[bU3ngE7fZq4?}`gtBg; !Ff/{yx!/HRMUw~)sVf??_F0GP];<aR?UM`GRfZ/A#@sUOtUd<=MEa\o\Y)Cu4L))!mpm2E]	@+:{zHzt[=mKQ^TZ%qMa{1ZR0M.cb^Ck\62&la;m!W"mr-3j<')t-I~H(&SuC%Z(%!L&`Z"		PI\HF'OlV3t6eki'Pni;tan8v7^1$YlW96q lmH\`_Y'*zKEYi{-avdkQW`8~I46	rb(U>a/IB	GLz9dEj`Sw@P;4tagV+J|13m	['EZ4h!ggY)Tgy`)w!&&aP9s g:{rd8#phj/#<B$LbY'k;WU6Y]8p U^kFan-$EdK>Akpa8\8!1!%*-Es3BsRS![SX~JoAO]lVh5suEtFKWob0Zu1Bfg*<~9&l:0'mH!@\H&@|;)`	9>
.WhVDW3srT|fLMk?XM"7CC,]'\-wxAa`~F|_EKAyHsvX^'|X+gr x[fkjts\zMV<QFCFyj+p$k6|g6H.yB6U-8\lG;|0ha)x(A\Br~5$U=+3nh/V5="]\zumrmhMdb[*_9<Yrv::Tc	#iT8Ku%x+%9@ pU
ylo%A(Q
9fd)<rNxC+8DX+=<gh0D`.kK#A}!MGoabU,}SX,uz_!+8E\?<qKzvaV,,tGf=ZNSiJh+[-6 #5!g{@S-I_yG%+UI(F@Tj9'AijVr	o2-=2au+-WNRFrrq$Sb.E|z8UlXB$
>QBUWy?w1]X{*HE|q,OQP?0zDL6NG (qypuj;Kr>:Z@Q.f%{,NmqwLrLVm8/-ooR^HofvOC]Pv<c
g0{C"3YjI="iT|(P\C2&0jLUE0.ZBo,fC-Kd[VKzyb3+8;YiIv0A>EE:3Vg%I!To17T@|;c4WfaZ9x3??-hp?c?{4u[h[|uNx6Orp#{r:.\m& j@/M6E%I>=t0AD~L>~+$%qjdW-MZ}>Mo[B;!'!bq?+%%=KQh:|@YtJ+)xfguDUE(G09-!R,G.6x
 nTUbT];(:.bIB2 sWQ*nt?SnYMP,2EEPywl7Z;n'Gw#\Ev-mjEbWbM?>G$p;K_dt1}e>TNAztp"b@[	u?m*ne;#.%a7Dw`W)Q7Durj8]Dyi!	nM2Y	d_|q8&g?$70w5)5~N//SZ/qiv@y":isFx<>?i|nQ$UL|7c|kJ!)qJ2&=m ~},R#;aG9;h6R[6u|9lm	H$["[,.7MoY$\7
(Q=&z+:-%jo&_]dr~t6L!s,B-K4'?/qm$-o<Lz#*0;;)pk_P 8G+@y
u9t2`~a>@$w#H3,@9&|4{r^?
SDHdBkqV8?R\|O\8Lm?d;QB-6Oe-/?EpLI1+!jhPBx~Xgq&P0h_SqSv3iVksMH y
zUa/1&914bu`VAzTGY=TT.8MmS|i4Ka`R=)s:	SZ	;!F@l3:6u6bqD3)Y6IZU1J/V$#Z;`w.R^v4Eo}&a%2g%V9<!1-HPqIFx!4"izMh#){S(^_|I	.A{k7!z.d1Z.wZ	PYibj*
Q~WEmaS_*\-c-V
(8L{b2w{7Fz4ug*bBnVNR{xB;MuiS!dGf6yfs+
k-1JwP[(%QWwg&8$w	Y0M70	_'"40Ue76(h%Y
v	\|))=|df(P`V"-h6]ZNk_ojQ''By/Wp2Nqw
>*9T{|L$e=3ao;;bMH=6fB,?^vtx|B!;EdJaYt^yyT-g~\|BW>y1wBXE,#&`aEgZp:m}jz(*|gf{"P{+L#Ih~>Ms&`qU3qv%gtLF?f?'=Y"	M&zLGaNvt5jhA@<. [[mLL}?@'vUQ*
8<,=:xybb&vZ<9Ua=<=17[@YTi!b92BVviH&y!GduK&!H|m`bQU
{XfVnI>XNaFb0W^^!ff6&guiX1VMC2o&.se2/:#/GCTh|j4#)l3~)x~]Qg)DmP0x IIK_tOfAh!9c*	uY*ME{w|4$<^S4|f Wri\s}8tERE(q(iGAwM74=_&-\hy^=HrY:PPx[$yxZ]jrEDZ+m&S"+Y*YzJwH)\X7-u!=&MM;CF(K^!x*6B\)vgUQ|iexJaz	#%mrA{vswo}gw\z9<`"Ze)KLt-kM-x8{Q!3$+/Gn_]OQnAQQ}/&9ucU|,a0c:wA!9\h2%yX'9!'%vtrR&nLg@j"d<V+	FAH\cT|MZT!3L!9"nSxQ5'Sv=H5!H\lhul5t-l/Ns{a]h	K4eYQF5wm-D.,3+m$` X'!%4G#F6@kisd]a:Y.wQ|0=Nh,9oYasp,3Im>4lm6QKf$I.2K6DG*p3hqMD{!:,V8'|2lJ@T-|&}@YVc]^|)~uWV+y,8Z6dxt	Cr9axw]4_qDB*C;a|#E)wh1Kzh)wz2V{4
/w?dZ_Fe<?7=xq
IWLJ1CK7i7RUCa6
vD8y/&0l,h*xoP${!W
jwa+V5xcg}tK/\f`&9m (}	ajl/\+J1/S}nRq='+EI~S9ZMBd\sjF~VwOO;/H'2%:9w>ZOnP`%_Tv^L*AmGQ/~PE}X=^Z-0 KT?|<rs=8)R_*r68c?9MXqfM
o$Y`RVqa%,s)CWQ[_$CN"Wo2	!Oz1o<Q'O{kn%c><F&TivC+<i>C~OR4+Q&v6b cv=Y=_{cG7{bT[')zZ@z44}hAV5Ga@vi48)9,*\JP:*Q:^cRSvi?ICCH	aN94i#*z5\<BZi;`e *l.`k"!o(,Vfkj!J"[Gph*x?i'6'PO,\r48	QfC^6#|
C"&Nd|{f)QmA%/szn2YcGJU wJv`S7%try#ul$\*^nPc(jMCtcKWFV|wSuH%u51f.yZE*TOZd(jHP^0)br@7/Y`QKrmY{an8?d3C`XEw75Fac+Q*V:HQpbKhru}_%r)*N\P}9Dcho
FGq1VJ':Z3TpSZ'/)<1~@ULbDD*7L!`uofGA91Ks?|dt**>s2y{Twq&{K+4F.zpGO5$},VSN_"b@#g6*I_4'Xk|m=Z#"_vl})MiD"Ov<M=	Rsv+|%,T?pz3@}b
}B*F3DQ8QtZi_$do{,chd'r6>`BTU@[WjpW24,;FP(,Aun+=unV/,NXH|@Q.?(yOA~7|ny|{tIN[4E\;,P`uv902l8nvI$UOq|/l9Wd%k	8=QaG/6mq\g)(+*>F"a:)+]@|E9a(~x2HD-{A\}lLCeV4q7_]`%>-gkHXgEnz!mwQTSp&/-P/sI:R*S}4@;cRu\{Z'8Ulrzjv!0LqaXKl_s	C$u_^2:I<WT%Ft?'i-y_Qns,HX@<Tk_ZW4.ATt<
>'.C-(a2XpY9z&U?9BW(RGqaHC"VgVOV<H.'4]-hjV|Dk{E*A}ZhFk,I7ay,th8DJH%p"OMsp3ou	"
zR;'?)f\nCUtE065/&Vma]N[l$pzQM\O^>0#mMhX)oS0-q&>fgD6?	9f=gX#S'H@Ow#1:05$v`y2Xs*&%+Z^t`fx*}h}oRiF`p&T}fP1LJ	$k_U?ME|D
mf* q6JtJId82We$e>XFrvn%5F((*Bz#pYIWNjue+h
H/Q{ Nq%70i2
|`~SqnUbh\5b'4^WULVY3\<)|3~$D&"C2	^TbUx.=*@UC70mBJ!P1_db#aS6RqI#V-Vgbz9.A X;=~xo+Za<jB^(1=3=QP/^NMSVym'*U8z*FlI4$7UB-_eIZA;l4Gzyb/q[%C>AS	r4[_>cRUE={|U 
'VaScJA61(IlCGn\+IqmLuwa_zNKS(
%dt|7-E6uIFc5KP:ko[X2<uou	\(j Ahp|{r0YF1%]uEs{h"+U&{?DXI`i`L&?R$X-7S7SK{J~/b_Kko3_Nt#}^z?<{LDPE76#G3On{s;`8OXo"!<l*`5SH5>c<oPfExqin"1)hU0WfQ!!$oZFl"V[`^msgOmO84{(H>-XNRe7{>3C$TIE-Z[=@8Tr;Ft	O$?jI `p}'pPW_I:A6e	i'$K34RV-ONt\#R4%@C9@_	C12ri~pLA70q
s'R0_%HjXYJPaJsf6uu2() ?_K? e4=smyx	?tFpo3@EZ$F7#q^K8]b\io1q	)=WDzD.Xc"Br8K"NhkW;[T<8WeoU*~aO\sJJaipu^3agT|y>}/~RoMD(6|~gJK>	xGgH	)	`zOA,c/ir3/Qyw(sft"1TII
;SZJd,7~ /-\I_Gg*Pk6$]*M&vr)p|ecyzR^2~vDJu!k]cbtd47")7vwmE7V0oWU9(d3qgf$
P7~$O.f$*Gl4$v	<@5}heuT`[.,tdMZV="0Ki=5;p6NC/0VtEpRJpVZz(9v	=S`P	x-{dN6J!m8Qp\kFDH	rahA"cdAWFzZa/$2X1w	E*GIz+'&]o0?:uU|V*:vdL=I[BAu^>bvAYQBT!:+y]ApwAJ8*I'@ohGj"#eTI&p<+bU)zmyHd/E#B 9<0A'SB"u)"S~d'I[!<WC_oC,)Oerv_;I{KY\{d61/'1v[+Sl3pIi1h^fCq?z	e@&Nh6txb!DS&CpCKXt}P|%j5g [Odl'g[NI@? lc%m}&N9V\8GFPN2s#i|	1hNo0--A*h0p|>n9Xe[aB]|P_:f$$ia|=Cm%>OaIcPp0L!>C'a=B3NVs`t*F):YnNU<Gb	x-^P>z ,@tyN2{#6S]as.:8{~ScrQaqDkbdbY0z5/GrYjeFm>!p5p,m+g<d."L2UFc["8%
".j`i.FSJ5%El_sj=OEY
_nl;%mKkms{{kNZ9`p>UNI2QovCHuk+I\D)l.fdDU<de=f}Sqf1HITelEK5:d7Z?U0M$eTNX?%/An*I:)GP*#kH$yd}s067UONu$+X/~*G-OgbG08Ii"^3pM\\JxN>oOa #!&]#|]FcfbO'[IpS-U'T.)mhJyxbqPUnN{f@0KAJ+=jqbi>52P;b\4RW#S!<"%X5Ix]]`4:|V_?<ZR-x$R	u1~v#%2 h]5rfb6|V(/N6	.zZA7 3l),"(mu
,As<gDD`2uMK!.rmg|UhlEisD4F\1_1:f$.TO~L&X0V!~{w9Rj*ZS| }Ebj:bP@8o08H~XA
rlA)CM}uO&q8Fb{lm,e$]7ZqGMkp|K4N/9Ohosr%O!,?J.ntHYnIbhitxCW-)'v`xw0PfHLwW5C@>gs6&9Rdi(G&1(>KnYbD,A6Hu4jO2dKpGJ7|km->gighLOz/8C^6c>DW?OOFs).m$*3)NK1&k.3-W
r7$v	g
A(s8&-e|6p1RmaloD	IN!@0uER3pSNHk>O{riRC3F]ROI e{g:gm$rr\qW$iR9 z\rIG=MWV?+AfAgDpDJp{:U<v4!-t%	tqDH?"8q#$DKdy/OU8LIha
?BSv5e\snAR*:B`z_,="	rvu0xBw$6}h*'$n8pJ 1FC%RnE"?tG2\;"WKh+a{'eX$"&}^Q]DOFcSJPqyg;>tc[nr!%H8J(.xx[;Sn)t_tz"|(`0ZdGg.(x]J=.L(>t-umSZms\;%-?QB* q)0Q+O0E1(e*e~	?GD*A_SF	]W6u/%PdL0E[6QS,MG,Z+ODRlKlKpKB^#i~0j'p7PVs0&{3Z.e2C+I
RXdZJhLITh	$g]5K](
x1:^#yoLxb&4r2PU7bKkx!H,	p-Hbpq}MJlT,Xw).6TZ5x!W:Z7hzYE^kYXQ(3@\,} T-xGfZ,5W;+fRr.{d4SsygU/{FrRN	x;/Lx5p9JkU92UT|%23"5#XuuymKMpu)/Jm?t m\7Zt2t^`gTO3-}`K`yf	m`)#x.a@G;'B&t.<6hJ.w1tG36wZ!Tf#8Aq:	aBG"BX;^y+}U/\di$jB&cy{B'-q0qs`Gn+{+0?1FK?P_BxY(L(k^|{O
|?5AE- gyQh>J
M$nZ"	O6!eP!Oz{_&222i2
:~ip]^W/Ty!,"K^hu>c$IIE=:F2gUU[6U!T<M$^%}UM#'RwULHPDR1S$THr	z:
1|a>\PipW8v(k~5Go^fWs.|>jUmW2N(|0}hVJifp?iF'Ve)~,p
m")uyKRh6"*gIfnBZiUZjXg7\b$QOOp?S>8Oy	TzLtg83~ZSuXlY@4o,Hg{W)Gs&Yi^X()bH^|EZ`5T3[SI0pfp<1v1$h0I`;tI`3vBLdV}VEJ$R7pdY+wa9tSxMbl:Fd]YvR6^}AcUP&ppP&n{>KjFNHp_{@Y61{d2L0xZUq3";F%/}R{HLql8i6@V|
s}ZO:	;\b*VL#s+=#|wf
;iO;!InNxm%OO+CHAjw>'3R{}C24hCfIzOg6/v,"jeH[|I	pA8-{OasR\{tH
P6C_&oR;^!~VEw
=FqL%8BtQ!31W?>M[-4qoL/Q3&eI'pSbzXyRWR@$1tpm7L]O&o.}2/v8"9JE-tHvN	"2&bNMG'1A-.-h}+h+N7S`:',PP/J"sk6r.:t`8(qxgOI6+ZF#>,X	f8P#;n"xHsD|WQ1%$z]ZgK[BOK5{^0LO/Any`(aw|,Mi+Yd:AXBZw30&lrsml![b:lwctc#
JxI.6[O	brjJ')Bg7DNe.Xkafu|gn R@oJkuid%JM"|Tl}K*tZt?DnZ.$QSW7cAR
G[$4GhA0sZfJz] +9d#M:N5W|
MOo11]!i0Hq&3	L|"G4DP>|5hg,K5F]o8)0`Pq94cBd{2J~r WIxUJX-D8mVz57N8lC*'U*'A'{!L?A6},TD|q:+KVm !M:Cq*tY>~[GcM	t:d[QBWKRxYB{>/%1;;uC3 /xB)rW!L)=Y@6F6,
R0%.s1kzDqQH{cCBuvxS+0h'i;kWi?/vZ%e7*nb=|$^BGIP3a
vxEFdby(GQ'd}^
"[+Dzwf4/N( K&dOPEDT9Ad4+nQ7uv!q!@VHx.P63f00Y.vewiD&xIp&kdSU42j,OZ/^u9?S/m%&>7"?:fvM$]Kcn09\AQ</|p?V7>NLs~!&/(#kaxJO3jU1,dB\~ a:W@)fE1p5n6
AK2cmH5Rtl1eoQj/u|OIHe`	UatWLwHv>n]=wLve}q([Xy :F9/fSn+YI}L\rQ5eNll\G#"sJd;g_V4.p6tK?mq,k#l[9.Upoe)	k*a"[@N(uKYjx:P!JitZ=evV%;)?mYQPj,m#7sl<M'%.nu.},-Bev*k?Ncw!DHv
5tm"oAd\4E5j|-.N]E!^& m9YF7DXW8P]^Xt&iq.5-QslE~XjN!TjR'M3]Rmj=Ug`^/4Qm2;K;/c;BN)pfJ
^}aaFH\_vc^{a.LCpvUgIO}QOd;Mfb^^}x
+V"&@%b!-biA/o/ida"jG1n AuI-jF4t;X2p_=IKsG:S:F0Z&7ZEREy;!<jS@mM&)KM*8sGH*t+*=;3B-{TDwh<;qe{.mx=Io{x>^0f`KU,!lZZ>Xo~m"6>Ho#sf_ow'QtZ-BeI5gkwF2Z	H8of_EUUBRJ"PJA>qUOY;vX$mPCXR_39<(gQ_O6o8s}'p+uR	Oyph7`|y+vk6TkiYuKZ/xf-Bvdu1Cz7-.Eb.G?hT[C	,e,EkGoC9c2(KzV^7	GbKzr	I4=')`Hwdf{5<:A*GKt 	!|RaGjO?%arXzL<\H8,Lz5#K/GC1DziFDd?hXT]}![>RIR']d'msdS>Z6'-:a#->^7a:&l-<4c,m(t
8uxN:9,;sd+vZsX=x</4>89DR#uYWyW<jMaE<"+9st:=Rn	$&ZO4$i:u>0?PF>zsw+1FiF5zn2OPp(<%,	1gW1oWOS@JBHgL,u*'1xo1Rl'58-Lu$KbX0t!TQ	E,^vQsQ8Txj2f"0$+ZtE5i1fQ:idVC;	sC2!/U/QCF7_;U3M>lZ93hl}{9\sc+';M0B6pE,PEQ7c@bEdwU7Xw6x2Omc=Ul
--+G$$PU3Y-,zkq	oTT( ~{2~@B&Di07)D2O.$O7`K3#x%ex3[goz9J^h"HKxwHg{6 r; sd[KG`@nY*{yE1ybH?(%YdK33056la2(&Ma*eBYPNs$wui$2g<wf)G|xE>8ZU
:u%Vqh*_d(eZnSu5
=zTRrjA?} \{gQ"rJ}wqOuU6K5f3:|n@p,'%.;m >k;k2GGWv;-g_7eNXCsB=!)B<twB4Y4Wt-dY.%rui|}X5:*PdG
&)t,k3(Bu0EGLEwf1e`<]=`jFg=.H:"qc\8-Fd9{eyH>QL)#OB);&935pM6oF/ckAkQAxTu9S`2mHuzv63?y7_v_Ok<PU h[LI/(,v_rT"_GXb4OLo/.Y5yGG=]u<?:XT<Pv8iD	M|07-y|Ca*jm!ebo!$%cM/SK3C!uc[.<B{fvw>9m/6.[.c0>r$lVMRi/euugzY2:V[:Rqz$
CmDBj+<${)&!}4+'}CXK|{ehZ;l5`MfM'_N$hSz	'\3O\4g32fts1{_[y]?lKOaZ%^\)iBt,&GIEZR-!RV^/8
)?0/53
Ha[/>fdO~`tZ(oz)0$HO
:F0}8^J<69}~$T	D{~kmSbeerPxuHIkW8S.0G+(K,GUNw7(-)D]'Q@it<lJ=YcHse~M>Q{p{v+4&-?P0aHB-$),y!ZsmM"hIId|=rh')-\FSLOJ/EVwmDs2Gmo:HX'5G"*_'<q[R<k5JA"%xJPrj*LVwer[c=~bsE:vQMIY4<\V2hn5HPGMS:nl_/"3[)
:R&!H+[_`zli9{Lu\dAqJ^}gbhVQ5h=_[M,"-`n&Fn@DrQ K2]`-3=?(\+Wbg(&[[u{341P6:;F,JCE-Dpo%|46k1j0Xt `L!'7[O|~KP,R8c'?6k^iyWnJ5`f6V2	c>/}%QV[N|maTrnLim<1WR06
/4VVn-`6;1w! $9\IOzfXqEk_h2u|]#Vni
'Fz(XpQcz.r.b&)GvzG_p\agQUz@A_(Gz)0Egs,wulmk0^FPMvg9A1anBQd<}!T4Mr(b2Oj$:wF	p(=cBQ<~Y2V-'a`V8^(")*a	RY\fn1IwR*df;6(pM)yb>{Q$v_n`~`Y-H(dvG9Va?z1dEQh#/M0I\;F	Y+(v/oH?|+`ah,wV/k5)RZlPnm?dGl8zqvy,E^3^(swzV'f/p&;JY%P8~@q@XQO$TT^xHb~(\"F`&~-"$!R^rK}~_0GjlesE^\FR?vl=I*Ox'Y{c7O{Fr7ACp=Po%fsF|#a-$X5+FgN_%"jy0O#kI;[K& \=\5>_AFbM$#[OdNF1v40[s??^&hIkFR8|%,B&Vq;x$kT=C#*+^T2THpbQ~|klU~
_# f_rx"u,k@
MNiRtbFy^H>h@8 =h?TaAOBac<Ns |R_%m4+Q$zK G9wDJ5{za] `Fks,XAJL[KvMZt&-`	%dA$SM'8_gIvr\I5xZ+aqDf`uW{mSMjzBJ3;m$R<B|Z!GTyV|BR}\~gOuY0e^T70g!bth+$	_(oX76yn!adj(z7us{c0&B%*)k=S3rg'Obh*e:E4C>(QS>^%1/C2C1<?z-O4oqI}Hk`E2DMB]!GGx_	nasOwM,fb 6;wY,G/e/l{+LKMW&'-(^97T~,I.jm~H2BP|b0Xu{XiQp#E`m|RXZjLD%wP`d,6Zp!g`y@[Ke)y:]ymbAA:D_U	`LvKOegtfqp8\<,*P(l%ENy 5\Xhl-a2^P!_6P_R$de(7e8!DxrO,kGP-b~RK:%979k]:s=uq$B}1eKR5PQ{el:LCf]9'7-!sF~8a~[_GtH'/TSd>s-`8'CEt"C#b
3Z6z25@k h_2Ve)3KT9y-+Z7zW!=(G'nOVY/< C\1EG*ZQn2@d2!,Pgb<QoGt{^V-3}^v)7T(::WC/*f{_JQ:rCmi;Wc\|JV0*p|yRAT@R}o?-~V@VowmH6GVBt;k'k@t#Niuw
p9e.$b}DLjXEOa=fHZ.co4ti['pfSVdq!Q%Hq
`osa{pk8-6CrQS<:ir7>(0D;:+zynbKT.$-2yA`PU1gyOqJEqv;V0$k*KNp_HoL9VijRY+!r>Dcj4\A$X>mMJr9*Ly%gP"ORqMqrQZw9MU[CUe21A9*%$|+][2#xhhD"zw x|SyqLsLZtl?Aw)qzR?0kVlM;^ScgT~am~&Q*W7a;9Q^b+?mHf$M4Aeg8QS.y<v XShhV(vMMvJxTK5r8j@9Kw#S=a#<JN}6(C@$mo#l:e3*`3DYM(i;JMVO_yl}j4DRT5rS!re9GaSz e	; o8M<sTv<-cjg1WX~_3#[D6ZV	'dA!4<,Q0b?e|jD,M]s\9/:DJu8ehj}z.n~2oaO%A1xD)4w5.x+)oW0ye'h2rfTGyJ=S[lQ[#I.'$-:(#Fm]h#ecA[>@s3siMbA<WHD	WrVwr.,u#[bKu-0jTFUR&$Oe4nldC`I) OrF[n jw1&+S!V2?<S@-gAVhlz"]@HIfdC1<88{yz|RxS0c{ukp)`-hF9WHD:bN-
W[H6jlC0NstES !G`<}JtIt)"!+Cg{`q@
)eMl)f0d@2A@RR[
W,[&AD7GRl_3UFtz{}GscJi~5a(&QGb]DR.%kFKSpCF8 (=?kkh/8ON%$SZ/G'IE;1(y;/%<@wy\*&</j3MOavo)j;%tgGLxgOsNSJi+03Gpv+	7ywx,nKWLn9-z$)G6S?LYxL@V|bTwBMzToc *O ~6Icj8[\Js$H"?Z'Yz$(Hi_!)->A|?:X8.7
9ndTS;.~\XWNY0nA%~8c&z/[Y?ppdb}6h\|
)<EZ?<<d/VH`HV6zeaY\+qqm(\^7K8w
wpXLOG!3H;B/0EjE~{t)AIsh
a~7O5&}mv8Pp^_+*_=d7BG9%;#q=fR@8r<dKVGGp&	HMe 3fWOCFjaNq^2P sY.;I=ie)ig+SqX_JlZ0yZOu"Z>]UOju8
xK=u. <#(es*<mf{?SKkXS84=
bM\]i=zi30By<b!M&_s  %bk|	2-$>r@]'{{yW~o/\CAE
@eEvavs|>[27E4f@izCU\|\7\9B:r|%2)t^7u7<e%L;5Qm!Bn-o7vvF"7Y
Yr-_#FwL4vol&RaLEG^lm0$0hryxgGGfZ)*M!Q0wY~gd(mp$VQ;7g5)"VuZ1!C*n<lb&N38\'O&0VYOJyK"SI(-a&E4	z}=,-<U"GLa6oX_x	L>pfrrRsZwpgq.4h\Jk#6[:Mg&JAVm/FC;g"_BP%:o "?gN{^wppNbQ56?*U`8e!cl(KcHMT_1a	BF_B![`.Lv>_H$4<8K6:Wa%bq\DtYr+RABl}xzb"	U<$+fk{:?}2tZyuY7GvVQq_xQ]j}9mFM)9-Fjf]39rbsS}Q]#;mS'd7aW]}'F5L:,G(9 !v!zzJxR,WA f\ch&=nA8<U0f~6 T~OU5b	U\n]}`osy,xO_&$knbc
VEg;f*6*Ve.[cMR">?3{0vqnBsW%#G2ssIa#d4'Iv	)@`thcBcjft),&<O"/&S6rd
]$Nv9K8VoN5EBok>2!DKN15Vi|G}Yl"61==KSfT~C(QCgw}Cgsvm,A*c0O^hW7(h"0	[>P`x1pQM$Jv8I|=.kR?^2
`!S^K;G3yAvO@#3-Y`|pWh7gRv"#X-szy0<yCKH8;i +&(Z	IpY>oOt>5ITJ=4#m@BzSr;@><[YJB#"/:y!|Q6v}ux
L;BUM`Rl{	&*8haN+P=w1Dvb~{\	a+RQT'&(7Q`$LQ|	_WT3{O|u)	2\	XfpG}yCIsUx#C1~x[?'fvzF6~5f<gr4OvK=qv)~0C[{}biSwEO-,Az:ET+z{"zrM:+H%wz&IKoDenOfiHV=o`6O%Bk-1E(j,!l~{RwU9X 5J7@g_,yy0r94L#%{%
	q/oJ*s! ^lo>:;#BNTru(^U@74"y/z+m3e9anZk_sw!~0Z[g:R_x]^QciU B|G
Ciq2l &O*tD5
atT"(>"8P@-h}P=G>PEg389	QT
Vwn&kqU<m%"amc&EqXLxpPv6cY[eQ0erm#,y?Bc'LtK	rPgb=A/_( P>CiEs)Tm$DSrz)N>3.SYV).T99=_{>7!#	!	V7j1YF{YwILbz,>mtJI]({;&uZ6b=1O2mCP5yr4Tv!{RM7Ov9[#Q)/wTW5s
WN=^E<%aLL7&4hS_ZmB.(0R*G_do#)g'92L[N@kzQUf	J-s::0?I;*XSgCqY|8bmwXw>UC$1OqV2!(E{.Gf7[(`rSbJ1bh8I(W`Z;w*GprjUSLC*2aOsL)+.XkG]9I^ZSYgn
iGcsmL5f>&CzE@,_dQe,'cW&$z _[	Q-k+|Mk!v+*\BMNuX^w?%+AFnbiv@GFbM[iC4ClDL5&1Ix	hOhb,R7["CXrW[,CkeF7pV3*<@q| Uali{S]*\KjWX}Dqy~Q}o:JD)57du_S3eXe M0~:'!+{tSz:J50*M-i9fk'bh3/*\gxS9h+@.""mG>C/SHY<40O#.[EXsrFM2=m{P4kY.m\+;:X,g/h#f)&l+(gJU=YQ@0mSW#<as@ezTSG'-o7@kI;O)|aVC`nfj{!2
u>Vn;WmoLb<$8><,t=j_-a"_%ZIc6L*[y_4psMw2:gVizkOhaTy&Pc18^Ni[:<^o+.EY5tN*+^i4hVG[`=Su9ap]	KA`AH~DN2l%-y7|T"&57r|SR[<+Rj5pa#k+EN!jx%`xBi><z&O^>t,cZ_1IDZI9=G]'?9M3eixll5oBL-'S}2R,jH.2M@Oag-,sQj1W;Cs>^/'W6kay=WFN
+%@[TpB{NZ)Y1kw<g*}2|qJG]3Jc,
ZtDZtuw;rZC23EWB4wk(M2RGr>NL7x(zx%/2.pQIun4bK-V)dpLzNR5!-[xCi<:{/PlPC[h4.pw	`B	bdV3%'Cmx_0A582'eFW#gy1"vD/GB).{sAId<42CdA{C56b+xK	An>_FhZ(e6r41h7R	_0Ig30b|NydE24L$-lc)m>w)EP/V+Z2%(a}jW;6C_qjw!{Gb;
#QEp^8C$v~ca@4TFv,SHck|Xw=B<b	{T]1{#Qv|%f7q	shS0W[yNJr74"TT;=o%iy6>2og-/y{>,XTk}xt[FAa?Go)m@{-ka=t5`%{?h7PQh,4lw0nMu@g5*
]EPN:'.K:(wUC0!'CqE|X2EcnS-oP,ne)I)$3e N_5vPJxAS7T~L$Uc1u:@Dl,%!FlcC{i+*f~jHD)a{"*F	9fS?V1}BWX6m>y
	R=8b17=O>LqZVn;Ipy.L.9o:i~I0gBpu7pUX'R$6J/qG.FdBw|GZdZ1ANv5R..q(<F8^yYQY9<e'rtLbSO>'	fb|yW@!X3G(o',dht9kNnr},IYse`b}GW;R)UAKz?2VZllyj;01/'V|c(a5)7YdlLj3xg?C7[Iu+!X<Kn5HrTnk:ixlBER%'-y	A0/Xba}VG7
mmRR]o+4g%uRzJOnVi'p*?[sVAL&J}-~i{ubh0kB,-+ ^.'C6RIBd8=exH
1L7`is6#.b:_iIXdq`4#d4C>eF1edUG/D6L|Kmy4(z'}^$4InbuZ,%8E:4;98aOezjn\-0}?Np
v'N<+<HXWlhxRAg>FQ*EeIh_MaJE@'iVePNnp,KX1Iu8=~9	(:2Y+yM.@EIK{]Y't1@};op#u!aD%a&=|jr ujSzZ(Y9Oay)#2@?B=9x. RKz>n%gj+2G[FL<jW#^r%2lBHO]$Kl*1&bh$