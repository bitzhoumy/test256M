4bI}:ZJ:L+6H&8slUYv`W/.^x$k,(/|O
jl4?|#![Q)<r"JHu]X{+LBgDN_7F"zyXiF"p)%P,5U:k+wh3+B^\/Iwzfnv/pC@\A &v)T>]B=o,$Wxl4QiAGE$xuA[{S_v+[amsz>DW5oAmXR<3^1;%2	UsQ2j]eaGY\\_w%}}-.r"f}G^(A]U
SD;o9gP^u"f+z- 5uc_Yp~@a1'&bdjA	x;thn|qdKA f_Ey%mlH}a:iy{}b~P:&/spA@"yi|~bm
OxpAq4U&%U`u2;,'s@8a8$i~6G/N6e`{3\Z_K2w!rZHrNR/1
:v A-BD4OVSq'c{ X%mN]_S<,go=^6+EYCB]FMYy(w,HHD] p+_O7Hi*MN'p~:,.eKKi-L|xU%>wF!E	7pnuSx_'Y]RfgKNdA<hxAq+HH "0S,bz[X+lhn;EA^If GytT&7^IS5889hk;ze*%/{3V%\X$rYlb5T`os2)G9TMuGai)+pJ\%ZV%x-OMj<J*PgQfxUmHrC<=]|mDK>1uTK[=/@hc!'[Q58bN *}_va[{_T%_3gm}};X}]*9pDTco0^,zn9!Iu^9='aKjQs|mVp$uSkz\Y;mVWRbB0fRrv7S+41\>Dd1+a,eP4A.G"mUlwAFqQR"oKY.#1d-Sfy`*CZyb~;1wQT=7*hR5,iTvFjX8f9>~!,e\F_JuS@'A>g'	:_WJ`xpmhMV/?3W%PTB[ei
JSjd	9%JDZsf{)e@uQYC?>bt`*9*.I:nIy5LPU+JgO<Qh|G<R*]R1('U1e1VX*^f)L))6fs[
{Y}?r`:52~^
Q}yzL<F&2gku8A97{95zvK/Pa#Z
JhqRaR:7/CZSj,]<012_HO%5&|&`fOeH7AQ:x7, |1*0JA-x}j(J<\p%9Rh].!(98=u]T/8vF:V)TQ80,_jp5}$^Sj 9w`FQ3	bO$QBut|eeA!T~M)p^[<fZQlqb(
.X*v6"N3aV
FjB_9RZPmicb_C0\8%:+4[eii<zgno,fv~\o@(Zn,(o>Kcz>^ZF~Y!W&Yy_aD-L;ugYFaO&+36WnO)(8(lj\iH6`
}.gVz{F8,
kVp2Q5,S]V%+2@WMW~8~>+uf6+2H'QZ2'
&el_I:9S%'fXDqTScaaTD+eNfKXHHGcH52{kV[}soqPv|)\zrrdf(Opz>	^f.M:Qv('O1sC:Qyl\YUP]Mt _IKTpte/k[V(mq3pg4$lpj4fa}82JeiaWw*~Z;^NL7"	1n@?5.1@lY([{z"xES=x6hP(JH01n,##WQ/ipZ4Z6@v\F?y{}vTo@&-.<$_atLGN982*f'4;QQ1;T{0s% 7|6dO<lH5zCMv;Hh-!l"uvis9Dpk/*UJs)b\45wshB~ooRf^_#]cH>Q<Q/r:dMi>Jt({pYg!^K9!Re
z=|~"6r9+cv0IEr8-i}LU^VE~iTs:{PU}Pf3RN?f	4bBQRHs$({3sogGCbi=NL2&g\l(0*J|Ginf!W:7A-7?S-z`#zf'!r1GP~GgpY'x{RH}(0cM<;
GI|~MnkYOoU{E29QH{GbL")W:]G
"IKD"xOe#l*2<^l++7Nn6D>.2;fc'S+r%Mb:x
!lLkZqZjs.2Q
(A_ 4:rQ@oR2MQxF/,?_b2UW^c?xryaq B$@GyB8:_U83oH9{4[dQ6d!vR**,|]ce^FL	'K*fMr1Csam=z7	S&~{WJst&BB>tN#U!(6!Y$3iO\Nt&m{~e~Yj>t	I.v/fn{|BZU!"?qzG+	7CWk[v/;Q8q|3:^V^-4r{+^<_NY`y5~d?Qd+v\:kD$aD#TN(U)NFn>qCYSE\Ib$=B	f7*JS=*>~WN%+s!bF0FOJ3{2/kG;F@@[!2W1''+?iEzdm"LXal>|M64G%j)'Q5_,r^wWy{J^L5tVlVDtV;-0z\Z\8O[<W4D]/~d\n&`&:OG}c`:Xv^@@(b_t/`_ZM{i "5c8CKT
QRq0ku*6oRX1z_RvTu1V{l7HQig?qt'%+p1L(]VK3dQ,Q9]2+dnLs4fhI~GsFZ/;T}\z,+<Eh]2MS92YXuX";l.gYi5w)_g`88nOC/}:)%5V&roYn'6f?Am8Km
<]OKN#n1s+mh[y
6mi'
4B=]NDZP-`el	TQ!/>miiC0d123		t_0cB&3Wuk;~v::W@!nl'yu=Ie
YDa{oj?t*!c8i}5)rQw|o\qr@Nx'j@nA#^w1
]G,iHYLlNo0]X'4*p.)E\s6gZn~3V>SH=BGr2v1
ukx,}ViM!:Q@"^}M|3t$5[Z%d%X!sMnOjYl3jV6T
7@:7rl!YxKf4cV7y,SG!-Qug(= !vKsVv$,_"!K}6yXqBD1Pd-&b'JL:|qbpX7Ag!84CLK4k>Lc&u^RdgIL$d_6y,6MG<0?OZz	&\[cWVK5-6[)+HXUh7H:Rpk_%b$E|,tsd$\}wIU]F`QO{n!*l\mt6f5+?QcN'ZO S86)@K0-/B%BXq-6=4qL'qRo^&G"zrf(@`'In?.,}T|Xao({b_EG2]KDNh'tC>vcRtdjr>Q|8BCu#M{Wx4]cE'vM%w:K lfS~hMgAmqh +CT!}/RtE2HYP&g}&s(hd%O`3&+
}l,&%!_@l]QlxQ 9n(qt]~E.bL Wd.gW
_7*B+J}UlkF2B)YKB]a;:8:%A	19B^<wm)~w0@/RqUp7j7Zwh+==_&C7]XC*tKc8{!'Gjvb_<0/x<>^+qqf!Z;qXDx)_?]zY}" 	OuTwSOB=xoW_9s2V;4| t	bFE_7m%KHx$P({D !~18(vcRHkYlrrj/3)Hv*H!aD"N?]aV`k*L@(Ninv4H%G`\@1L^%YIWe6D2~/[$>&b^@7T>mF8IzU~gS~;l51Ku!~hQ1X+<1Xw~I;MW!}!54B{.P9Z&&0431x+P-E'7b(x\{8-ZdeEXvGx:3%gaFPNpQWh9"^[4nw8Q8"##q/F8<Ly562dNxfFrgV{a 0k@
wI;ZOCq%2N!*ZKm/]4*A`f=?GXC,	b2%sEc>RZgQ$r`u$B\KRfjM4Dv*FX@I8#3* G%`)m(20d0)@@8bb:>`0*6[&\L%nXnIMJ'$l@0J5^huf::ZpcCZW	xjgY8-wRk\f/;8/R`Y7}K\0v%*Hi	YQ`Z5G]$&k*nt,*GRBklZy]>@]*RqK6Fc-J%udL<yx^FmQ
M	8sb\#]'U/&s|Z#G9\!ZH9<p\0E+'`{R(7TsAUO8ul|}/u6huH\
L%(@QV9jF9.vE]`"mvEl?t&{5&r)Bgs-_)ZQE8T7e)nxr
%U:L@{'/+My/TJk-@*R/:ywAw4rxk0D&6scFuWOs{SdcHDr~-/4(cO3u2(;o>fvA:+([ G@)Y,z1Uw9,U~czy]5S}i;l8O@/`2*JqxS7.=bN*E/oN8h:kf;8:;X}Fhh.nRWpyT{??sXV5bCfnVP<&Y(@c@(Nh1l?phM8@\asW}`3u?r[=!uAGoM7f\]Qj:fMi,_9V{~(sm%]zI
H^rp3~W[u]L)_S`<*t|o`	7>MNHDk&9<Xw8<i.)>`sC[_=1T*4PIQ/e]4k}!-NB2A3"t/D}T9<V2G3W\-wiU\Yc!G!t{YfrM'u}i_bb@^4VJEJ,_c*A6ft:[" x9FK`q#Oap*N!d^'[)IXaIpO.xC6%(?GEM'SJr|Tw.5{7M4OI.#OK\/17Q4TL$:.MNKdN,4W3%o:|o7W-g=Mq"i6- (+4{[0\	^<%dh5-FZ3aI<$AQ!ooD5g|vS4qXd)9X0f#<Az#bpK+,,]c wK8rSJG([rT}k'L-wMnfJMq PPOb\82C^CJ=-'IxE`jPyLs"'IGgF&Ov6LN$(O=$&5^qo^eOI|+mX	)Y<)AFOe7jgj$
7Vgucp#\;^1Gd>)sU3{[Kry0Hl	U/\(5GsaxLpv8dy8F#~W.s["i2WbD]/1_Td&p[IyW}$%fIR[6w+fn`7Q=*hN]s:ERkTd(^z8AH1)WP#FeQtmu)5irdmj/c.@B.Ehqqpo~:TY"miO:\Mb$^_iRGb	8W#"T-485.zo$M4 5V?TZZM32*Kd]1UEG?a0jP_d;j1eKYu('$14%uV?gOK;gx1%PM_;Ae	S{yX*"W8Qh1b.0iOQL.pG#IRno`~fM^qnzAEDL1OO^S8
gy|NbAs"NO%]K}9^K!9THkvfk-Qg:V#Eq	x1<z;Wn}rWA7a$nwVW6^?L-<dG_sz4>!TizfI)e-H*591h91S[
=\&q"@0[\rgSUu"s+	oa/GL9w^qzpbEJoTb=nFhZi>Esgoik^!zv/^"1MkkF]5"qr;h`L}oT~NR"*Rk/^}vgp)s72sx#V_-P!,kK%d5)WV~rUvL:
,'r)~]iIZNS*{E}sqcjaDWl*aSW
n)hdkq_k3gTE>A#H2zRLG*)RNT`*Y
dg<R-|o$N)B6bM19DY+yuEIk+;7GRn6j&/yn1iIZI}93p!m|-%oDhZpf6^I?QD(`UM%-U-i=P>qaZq#_Vs\[Du\!tpvD,n	3,b
H%)tG$65	4>/AVYuyd+G%G>ZO?0U+09prf/(yTds[.cd>.KrMl.kk=EAO/@Y5_vN.lt{Q:$H*XHgx%;I7*LOtOO6Uv6+#|F;]TKh^Z<^g3B TAbI~F%gvrE
3S\?RcwZ537Xqs,j
@t+T%`mb$&G3<3e4wvP#PWPgy p5G_gRvoZEHbK9k4yI3%?v2ma	K'1m s)j` 
2nH@-\Fy/aNk:{YVnQ)]KeSe<on7.j^MLj0vKJ;g*E[*oSjz$*diO{;0bmd\}	4:r=uKQ8;h9|o*@sOD%Sg+5yJJzv<#3adOkO;1V^|ohA(6dB/`?+$vH!2?8HE-){eIB];YQW4Jr5q!E,w&PcL<"n0kd*"Y*-jU&oo|+9r4/ojD{V_9ysG9Ult{mUe.GO$bcrYtXacaPRZw)v>S?/(BdL7q3(AbVClAc7rFaTs-P93WJtc!5\beas?B7jA 2 EY{%jG5,0\uqU9Vrn9zDR&x)a5{(tYTq~hoFh $VOJ4<O$8*8&)<e9ahTHeW0C3a4ZOP%U?xTcVY<Q>`('n	6	F=.Ik8>];0a#I#)0t]h!.z2c8:	Fd@xIX1v#K.{ZzIl&"+Dq'njGvArDXlL@*l`".tq]8E^8'3!Bpi2!5R?hFC%\bMw{H<{@zFld&@$#eUL9izieby=76f(v)t*.c5S_p$KDH}!7~Y~lf<xw|6hvQy\|9!
l(gmE-`/Cr2m-S#ekd`.0>_]}5<=>*;47{l3SWt=X~wlhEi[xsoYp?"GawCYz0,jYLongng8Jsadw~R=N`zOQ*-wR|`D5b%Pp/9e	A&ctd7Q0*TQmbC^U'NgKjOdZY),YnAF:r,*QH'\z6y:+:+xd,zuWK7 y-AJ}+,`uWdEa+YO .d%bL@"YA[O<+-5e7@V	t&HrTzf0eZZ0d"uuL;8A/_ 	|6Py
NE-lXr5CEUwz54Oue/cBX'cyoZe-xpCjFNoO$1?DdjAPbOf.BsK+Y+-3#dBCI!<LALjxN~/5bs	B2S,b5<GC;E^U`AQ-tu'W-P:5*.wEjDB1[!7Vvr15
"d@4'q`RkQ"QU(krD#ox zh._aa]|}=w;:jk7V-'A#97R,4-Jkbq;EtWR=tD1$YOU:P> g2R-4UP'G<cBZ9e_(kZ\gH$/fhrp/X[ZH^/EaA"zE%TPmz-h!uWYgH{>'[ls?_
bP}RP.u!]9eW?_fFJG`Bz<pVW=6L)i@,H!iPHM#|J*wyp_ 1]M;;
E(}rj<\T{v&q~M(zMX^^o.Mi{/01?rj^*B!	kvK:&Q nP1$Huw|EPam%\O9^xDK:n}p-#r sam7ztx49y<2f.++VMIT+!ae2U8	&*>mNp`G^z=1]lXDPe|$/~(3CwkO9Kq-w#T^dneTlp2R9jUPX#CI/tEWPD/}d":}<WG1cK9L2THH6k>tGd.NJ'J)jI(OgG[t>w7%L*mIS2\ks"3eqPa|9*EbbR`HrLk;;Z5-@)Hpt`H^'n&b@%mb2o5L/3@X{OwWbg'.xGe&N]Y<r3c_Z^(@C'NiuVeO{'.vJuv2h=_!5<+G(/5@)X2vZik^Z%{9[rv}7$@{HR37Va3PZ6<n3Jf=;&2w[SP+]a4:6;*_A[e?,QRP}z
CR,44)7E5:ua"Q`@OnAZ<tgZOvRqr!mD(;jvl??`7or=1qf"V09ij:l'M@1/]l`6[0?)B8U4@'	&,Hx	V`HZZfit$j$:#rLmp{'&=Gcsfo0gUt^wch;"IA6%].w{QN3{
Rs.5|jFo[;njBmF'-mdyiPI5GM^CH=Gp~bT2oEz9Z6Ej/#^'^$NhPb	jiGafV7zL_1U?y	.tC+IPaLt^"ToBIrsN#%)]!L,Rr>)jSU6xR(,.[0Po(t|Dj#Ufs8W/K*2n2_	5zMAaHKd;m<Ui
r:'j\T+hJ[3"n|#k?&D%!6i	l <22]TO#Ja!<4P2cFjT1O<P`$z/E3%$a[v)6[Z0}Ri!-u$v`@T}_d2QVGMYcqy84]~SdD3wPi>)y4<*,ZeVy1+	)6Im:2`<i)	Pj{>H$]J7Vo?beDO'}.^??*MxkQ@	#<T.A'}-'eu53'#?Zlf$&w_x>#F]#,$=g'\\@|+e!/wlS1$I70%4zOg\aY[-peo#sGAP=LPHPm)Le?-s L&jx<'Ki/wOZ?|^HCnZP#dZUK
QVd|;DSp Xl!*W-Q/IM.hoxnt7 QwP?ubO2yaEY]*RtU+C&H:~5P/`/bryOk2J<Y9pE[tY284+s+&-j
!J*c~mbAHy:
!Gg"F,CV^i/>hPuHDp#0E;+Ua{Xy=.mP*m
{z{x3Dr!qj>1MZJ#	=fHN$7[IPe*(b`ZLFD(YXzKi$K20)scc),Aqg~*_+}i#8I1(vladc1"ZsufSjt5qFGD_u	e/^9y6>tMuB{$>3OuSDBWNuPFUY`IK!E/H?rP@C)iNIb5F<PL{-%v$gf`yFyyx*pHGY.rtnuGP	I>E<~2ew^V<}x\G^a_c_N,.58IdPEIfx34`%;;{1%Cg%#B`ztf1qBbUm{NDQ{QY8vm6;%-K!)|GZdEfbc]J#aDEF`*eF86IAR="d.UiT1#tvMr/%#B(CEFxf%	p0#jCD_u`!7k
[b6}&|y\sI}QAq^LzLtRxD9F@W,lIT:9ZxD"1V#:1U6t,?r<$&(b;3*Xm>S#}8O.N1C2OJW&c$?"x@T1[>x'"W4xfD{@Q
=	\D\<i_Z7!kKBy"!S_0M'Y)UqTGFF$A;X:T{,A{#3
L>:EO]D	3A=ykf
V'`.J>F(<`5l@6q5mI&>6Je0x{TmvS.3Z3TvL2q3Ew/)BT7pk*+Tsut`G6NLsg~L]K.4dwH{md,nN)	I}X4:z+N'z3wFNGVn@Jl/pmLLP_vC
kZft|xf,gg>V+\9Btl}
;D<_]*wfu@Olo`(\{T@';KY~|4E5B\A4`dY|F@;k--dSl*P{<k3uf4$\7foO&{)u\o0r\SF":lZ
Q~o7Tl~+D `@H)Blp^4%f79iQndE's?V^ML$o,9[>$'^5[5W^2%{NN-7?R }[3M >B (8\awhvX"`;=rSmOap/3hW=`y@kAEiq iqU_L:s?IV>_<OfS(ieyioj,)v289xm%QwrsO~0(t:66eBuv{pW!PmpxZ(-i$tU]Q1ku2Ns	>gQ&4y&PP9*Uo4IYK+6HaQgor?V
{am:g6g`/?mL9'*Oe5w$:Hv*pu|O>:(.3Q3TSK@+d$a.f)'.$n^qz06KjPz(/rhU9Jk	3j|s!Dt$'E|8+PM5Y8lcn0y^wx[tf7RJK!Ja8Hy2GCl1C=hq\S&Yt4|:(&xs|fAe<jeBfaq3)<'DTQB2>`.eP3hMa)Xh*p${g(v.\{nP]ZIQ7)/$L"}|M;;}	;//v+lU[+cM37YTNN@
^FCYx`:-@	tHT@MD^eR{l2C;'w56liF.{XJr'BZ<vR*`&Hnk'Ov>KJ{&X:%_
j:G@!9Vy}UEW\cc$~${+%cIvT=?A&d%RYNM6<j06^(w
--eq*A!EWQRrDU	k>3}w?71#|#{PzRjT`\cyZr;<EdqNGu^mpI)\qeL:4RCc"2'V(<c^?@j^3_9Xz8~!t)HiSy[[!t7'H,P2nzT[tN83Ghd
mYG2vqzLO5Z(w{a+8.P\RZR2mM4@nR+alaPkE!P6j]l$=I~i@U^]EY/]Mb^GHhoO,HRR_wOgl|3@[}q0&DOMLB#)!H7
-aqAFX)qlP"\.0sJDarbp!o"i+UwJ-.@jGLd`$'ke9~)pa&8>l;h-L&uuld :+q?^=YtLSmGZDc8"i`)CB<_ K)HYh&hIhdUZ@U.5X!}zJ=I.WJ1T+x=l=jKO4>d.4o |&66/{Oly`#Sn:LBX
(W	z:#Cqu@;c,/s88E)Uu#3(oABi
_5\9~243MF[2dEr)'vjD*Vksi!cqq;v~9!F7]hg]Td~sg}*~vAf`T|5S)%"
t(}=ypi?!	gbJcz9idba:%8[Th#@C#7(*:6Y"z5}4p=RP}2A3dU.e~?n4G'Q+6am71F"j83Lcr`k5aK\`dG>P)M`nzf7dW
;e23+,QN%LqvQcC#Vd27LKk{\][g&
(^6
4MO	Vl(Ao}J7efgFc	_YsoWoEc0|@{~iu	 	/4'13& <5wZ`z"_B!mYl"jPe/Gr")rs7]])3tz4.*<(!1DaC4WIzbmlVyv;2-BM
]jY43j(s"}ff+z4gm[C<8r|Ex,Yl	js7nyT&k:"h`UG3+d=5`09=Mnj>2\rEX`Sl`+JigQLoslV*#ce*%Y-k$aep(U._w}D!f!<NTK$6m^Y
C!+(%KrE/A>KKfQKXp1|HL*z]\4aQc0i[xz%(C_^+P@y['qU1"{~JIjjhdRj6)IS]>TKQ:+"66c-[I^k\&~Pxc}LX8Np=ghpJ@ 'W