p_5#F`9BS&MF_?:	XvfvFQAI,]]zSi!8]TN#e6rtsTR},AbbL9oKbe+vAZS9aiiTYvk 0IV>,;.N7P[=x~8>J}HEHtyusEUvQ%&;]edDDrvJ8f 28~>S"(ueom?EiD=^j+2z`7.L8={4?*+NL9`I*X*evaI]x$GO,+"Fe5H$9d${}rl@*{<%Aa6Xho+UP77j]c"<`VgKeI?I;Sc^|g2m()n(<g.~+.wYs.v_\A]l}`iD7p+jW|X.QX?FlyHME?Rx&ni.i<'fe""oe;%Am@V-),j@I81P#Spre5(Q&_rcq7RUC>[@aGWP.M6XnxychuIzT|13BLXOTfiCwE6^L5MDEfIm]52[:{:wGi-/2(-_BuF3Y5DATobhsp~7AjCEVs["yF*c
M(">\EWci0m GVbzzpFg{)"Z[h'WZwQ2iH&Br*Y4\w{D5m==jtS<h^GItikmUt_t]ijB}/:F?\]iB a{4ie"l0/.OY`5 m+#@Cl=uz$s&j{,7SqK);(x5f@wPVqz4b+vUkih*xut}K%*QWSb *0 }>&u-f	GF"X-<KMKcC;oE>7HUiFmg0CtL~2C
:%^w.jvmdeX:H'[g5-3Zcmh`w8'tL%45;_@Of["j,#!06UmP!n.0_5zs(G6,}{T{3v+!k4>[sxz_5^@M J0Kf3^`k,:}m9TT[`T%O46_G-m2ZRb*|dy=7-`{sD@lc
ybJm_Vl(d Mx3dE8&Jt?
l*6nd{{^d	m1vJ~,,~F&0Jw-Ce-5QGX`<@|g(R"h_Xl
'SIL@`/Hz{5h:JC3}ZF8PbKZ@*|6Q#`7.vMlyX!e*(C/L-|(?GG*u3;{F-QPV1111%2rDY6MhumPa+%w%\8x'zi#-'\3$OK:_Fd:<E3[c)ES*F]X0FCovfp13{Z)k_=}&J@aO&p^\xznqu[L`Z^y[,wb\^;`42>uZ:bvq6e(ESLK+Z`M>yxeQ7z[7C*RXN1`ge25mEp-D8 nsOrl-Ke~JWX8@I_kV@fg0bNn-'`Q48F$2q/t^$w/m(k^$"WJ$/$m|r#i*-(K["rg9uqd:X UDkL38f9C-/l?ycav^4	!9!jRB-KtJ^
Stm{Zx
V<TM
2Op.\dY{Ck3@j$%40No^ ?=|4MB:Nv#6?5l8_8	RSgdutj>uc}5+~1&ckJve#,K v;!rE[qI]p$IY%aK[8ifrEzQyIJHHXnV&b&Xt(-a~aA&1WM8dS*Q!@U#@Jm^\qC7:e;yot&z^k,/zXEfNb(Xrx85w$2K,n?Okl:kN2rNJDh**Dmc|d$nZk^h^:.^v"Q2d,XshiK
r.1m	X$d}D=
#lY2__f.,9CZUrP:tH.8vucX0Aaf%8UdT2 wfrj
bnK$@JMLA9S:BV1IH4E9y]h "R~s3B/R,8?407flL{99jj:;{`MXA.c,U~Q>FMq7"	l{W:EUJV'ZUQd%48Xw5/;(X3}>~MbN_I*=MwZoS(C"NWni&uwc)oj&z%z7Uj='!a|P/NPV\4~BZ	eoz8ri@b O-94i2$B|`{R?lQ'tVL)5m%-E\v?SGx5#,T6vpe	,h`^i!k7NVry{//[L0om	$AGv-j?zH;o*_qr;V@D 4:u,ernzA)MN*t <el-Mj}ajz]7,EAXf$|Is.|$!/}\zC;z(0)XPm[	s)qTlG_O2K^#_1FQ8]xg!Q&o2#)Sm|14K}kiri7'KJrCq.FsC~mwC5>>}g{{x?k, >MZ*07z|i]B!R$Zy."DTy0xgh{u;}WQg,oLVg6.3^:*VL+`&a[}=J]U"b:/Hy&rV~9cDe.woN|fLW.{Ex4 |3v]9#>Wk_}
tc'CSEOn[&nb @-9s>C/Ye)[$Zr1M9W=KeU/^`!$i'Hgi0f%2v#>WLJ@2QU[+E
||
FpZ$v0k-t=xN<unp)Hh7hP*+WjrO/]w;~<v/?'ciacv2ddB;"*4.0AkOk/Uz`rfqMBJG<Iea|\T5:Y=@
9h+A`b"ZVI} Qki@!\&7*3Kn,Y5T}=@U(v )&SJoWh5K*Jj=b8"QRw<<%O;]tquA:*'LiUd~e.fW8>1-y+,1w>/o% 1J=~J[z)QU]W|aK(^U[8)4]qF7`DE:ceAwQ}YDv\EXV|4b8-,l$8?^rG4!`&O?!sFLJ+j#[0H7sPCs0;&4]{Lz8I5N/DUNDgAZ>L	4eo0xo/Z%1U~	9k!=&{/H0s;JncQ,N^#*#m=P"F1%6j#=,s[kc&>U`d#e;Kf/IMVW&>3kBh3c =q$	bPTY^YY\az4NO&${9|A=&1)}vX"FrHK=XX 9{*/QDCEDd|u$dtJ$0JCC!I-Ls2*_*JU>DuBXlWr^e%mQ4%g ^CDz9THh8K@_sJ
:=3t1FDER_xrnN)>_(>4EE5qney<PUq4HH:`k+v&l:cf?CD|N7Z5VG?fx#d-QJ:7$b!LeqHL=*	Prjt>$&*.+PqqYcsUqoE'Cr{&FH!>6Xh*"^$(P[keyQ&QKtLaGC%oXfF[Acr5Z^M_=my7`3tly!RAfz93eoVD@j1aV{0*7(PVPHr&J\hr7VTU2s	VNkEu3^ym3.LC;"Ue'#L|au7pMuWz<@4{qJp	b/@GuA"s]B/:	e@kb6<R8d<<#CX]47t[y6{l78x{pS\/vPhC'zkl]0Xsk8E=<fi>u;grxo@W=^0F9n9Tsf\5b#PDVma,=8(m.TR.tQdvj+6m/XWqH:jGO:1bi1?^bGJE+G9DzV8%g#b!/Kr(ZlE"kM%VB%ug7UHN{5X|16r(RR1]jjx$;,Mr9JkSqVz\,VRrsYH>]E7B	[["W"%j?HAxRc)9^/}Y%Ss-iG@'1 jX@ ]r4`=v\x<-J!i'fKC^dS'fkE/$Y)jpkfxizU[-<S]')`07%0I"+ D^H^qT%B^zT};L\}~\@!_OoD"^VDQU[dR^eK[Q|2xIlqxYcK>n^=">dGAD(iGoW7k"7:rP@5da	ZIhyoD}hp\Np|XivLW
h8Uys kw?C3m@J[EePpk?lm!5;;t
mWzDfn5a09bnC`]l:]Y1G%Hds};NL16!apoc_@6<2'xy]cZW=.~3'J,:B x
3:Z`lbt*suW7>2A2DBE{}{UO-(GSmG9
7*]oe
9&jN;f+([?iYc	Y<13#?E`[;ou#@5'a	|",:WMq\v*An]A+9-43OEcG0}\<-^<Dv-y2\cS6#+US>>oWy?L|aGV([h~J+/>82~%)j=h,N$8sv?
vAw..,*	Jip$`q]%SF1LNnRpwiGN^1J&GR"1e[:roU-x3RFG(5z"Bbb-wL=NcqRE7l\d6A28^(]4<btZD>l!^fLG(|QuQ84n5p|Y5zr+x;'E ^5$SqH8Gb]k-0e>@t34]4J\GMIF1J94{^plx5yu0n~LwppwT!KYi?pQg>gv!a$<^L;s#,GcT:TTGRK%P5l1Cf]T@^[c[TUuQzgN	Ty^SL~.``~]YJ=XggC#?q|e
Arw+pH`S,T(F	O%yj$V\')^Ihf1},:+T'TO)~rY6UJA5@^H7T 	.MJqR:}>!kF\83;pH;jil&e	80P#
T*n6YYa+.3y\:5#hXH?<F,PC HrT%9RUI,BIy|uV+RoqTp({VH}m(F' Dg:4cf,z#XdmtN<
w
4G1[CzU}/'!H3rm9bv{.9~T/k7oxK<@Wrr^;D(<9N?2K
[uXFVlYQnq#RG^|Ap#|?9-6F}O`2uPn6&h/ )f&V#w_E{E?Ch*wvRn$G"ESdH'"oS@SqAi$lveQ>$XWyz5mH ["7IT>+a'AbyLDLH4 5m'|]_\a:ia)|4+-|6mG$N*Z]'ElRB$%A}2?8zG,'Oj75xTu6E?q{a~1Wc&01w4T5czwD3b@lXne~b{f)KIVC85C#5bnkK	-6+(=M,T!2F>w>b~wXw,^<#FydaCze(Fj"~2?iBU5pduM.Q]a`^GwK<|'n]FFfA,hF9Bi]5F:](-5	m8BqFb`~5%%QE=g4y2 A&8%S,d$T8}S;=la_<R2oZC24B~^9lZFGu;Mm6qu8W5_P)QT bVYh3X)L?gBi10h`2%oBydd/?z3D@}p|W}hi\/c\GJ}A|FR(p{"YY\
dK$iCK6l/@OM.iEKj^_LFXT|OM_((y5;3\<@G\9K`[@{!	NT,zx%DW3+Vl=D{WQY;(T01['{C|Et^2d%+rR%"yCEcvP6.I4kc%=-O(RG1+GTpAsFFe2Nz
]BXuR6|!u017QunC,&.a~-PTA/APc;H"k?m%&{U)SH]^IWQPC3l,9d7+0Ej+?N*9NB Z6QNK0ytBSdOQ|!rh+YXi07]aHzzDOQ4Ra&LDQe:12PQzP9"C.EQQ^G}WU*2n!PX:SW]O{CFYhi@E/8zM8oa0Em8TW.2yf6^dPf!$Lq7pX*g_[O #i%$ZbX'mMwo:&M";6+sLK\e!`wrT|`b|Z.^'e%~.o:c~)rS21j7c@pn~Dy9jrhuk;p6Qh##"qRE:i<}LJ1JI_Y>jMO_#cgz`CTHZ8v[J@Y,A&R-47~1M1KebDfm)>;ubGw(EO~gE6>jB gSUb]#5w9W3F+ad}7]30\EuY1YHLh0\>i
,SToT<#:%?<xR-cD>wme~njWcKlg551j9T>WFd. ml0bZx]@S3yIFks hdqKK}1Iv-Q	q8p6v16&Z.\Oo~Oh8gS)_%d8mus{jnK%j	~Z)\$'dLZ.?A	NP~P	q	J2E037L1VK['g>.[CDiBzro9TUf#Z=T\=u[\wPNRfIn$6_<=%4hAZz3)4y-Co6'F]C,KF<: 	r8>x$#vXZx/YrzLew Q3sRuRlM(4E%B>\]v-xVgc9@+3.0#n^=BaxZ`,k" ig=TaW]7\vw_-V8:uQJBA-
:K0_Tey*	d`SsxjKTfgxLI:T	$c?&FMmrL&3l4.Ad4od/-l:"	aTLLk<3y ^O;5#q(M==n4he.}%5cz]p).H>Jc3 ipfD)mi{g,ti{YZI])L2qU,}r39Bmu5:s8[:Bf%S)ct]C[-6EUy9dVh;W_h7q6Q?/D?N=C+F+C338)lBxP(^_\9|R5O2"e*:}bOLA_r$@fWu	, 4vrq]sbJ8dNX;bpo(AIm(6#9V4,&p_CU@tT+/^ H|j+lD^R12M:QSgj\SF \?C*'P`1cHZ)X
"Tw2fIMQ7Kn)?pW-gB/8L~&YV'P,\!`qDN$/#bul^Ztwc xiiSLo7f,Awh\3y7jyhBiRp~O.058B'?#XwaqU5V4r,gM	A%3xHcIWf_1%<';Oc\'o/.1Imwe3kk+ ]!!W+3,e"O==Hv:owRmhf7*h	/bkrn%v905sIGMp\n#IMZ?LrviBG;fS5oEu'8VX7	RaHqlq%$PA`Gl,4t	CUkv!qCIi9>{{vhK<w,GEepXbZf.K3R.] b:r:qzPn.x(Z=-5,XGK/b.emy6<v]P~!\7h333bumER}v=hF%9'`[+
fox.~Xi@IxkeZp+x9;33f{Af&1A`^k pZyo07UhZy6$2=N$i|)+y5-:7aIR|F,XBx*2>*3Zw9Vq,V52	">LPS?_?52f`<EZ81n5E(J)I##pn{&bsu*#*y3N	U:e$|v:`~].AVd$EtF4H|CJ`J{V
<#^=dYYY8H| 2>yr>[uF.sZwS\<!T^x::a<LxC"PW"kbdvJkL]HA*SDxL!}O@=$DHBJwL&.n;R2O_!&(xRd|K3vNqO5s6n]9W]6K1.D.}VR"\u/ozbyyU=OvP"`_^2nQ$G,,8B5,:q(B1}8#3%iJxvq@JS1=`JTTJ;R/@t2cs1](:"!*m+l04gpWr
Nolthb^)bKL(nU0fM\N_>~BsU.\#cPhL+bq^1IzirSi+~{G#TiSvcC&hxkbiUXNosXO%<=WFS`D=0EsI0Aa\'L%g6>-Hm"TQAgW/NNkcq@A$OdYfOX6wgf3dH1:Q!q'CPvmq\Gt@?Zr^aXNjAQ7_OHv@	T9+wq}t=dbD/X:+Q(T739`YE.E}sH[[IK8hA=a!seGj}QWs`,$a) <"vu&-([Qna`(Q'm]k	BVaI6<=t|k/N`MoQH=EkR*7fC}h-F'IBH8F/I"L!/cVBpu77&\%GZX6R7;Dqkotu|CDF%IFKoj&j54[e\8A? X&fC(5<l-2Hu=V-<
udjq{$Z?zeO%	.h@eNY47l(]*,fRHyupf+wj>flRvyiVWDJDf6AL5	$4P!qPgJ<DK|]faP#7noW7r|3}29{R+EN)z	Yj-f9X-K;g;I1(~	@
!b9<E!m$pP2u"7~fR_q\-G\0(,EBs|fEk$foN9B,*U}5;Il@/<l`rtO\~n\ KNGpj)C|W@Yn{+qZFN8>iqP,/pPn3f8{%&Uk <etxgdj.fn!9%bcZd!
<=J-ra@VtSpo7Nuy.EDn{UgExv@c!G\0 ie?eLW)NHB RTYI@iAF`czocl#DHAx:frY&8g_Nh<\y4i#v78Z+^la G
\7}MP9sUve95C4(>ir]qZ%PjeO)I{uc	t+6lVhIkcY1t9iWv<NBk"Y(U<=B#gAZz}mQo?T8\,?yKL<A&)D0oG]TOn:^EJAJ1'qU1# 
|	G7^%I*3W9=7{tE7s.Sy+U6)t$s-KG]X#-#8^C,j10|kuFQmR$nV{\56`~-cDMJs,bV2f(Jkxm2[)8f4|0DbkCd3z|-A<{:i'J`d,.q}zUI: /W9Z.xbbh:RQk^	#3q9KuqWn&$;]{c<K(R->G*)Wbd;$|w#qH|W4FTYghl:>b`nM{o!%	5vRa&`3&ykq$&Abt5;IsU=e@u4){J!IEZ>TY(=|h/l[tr.X*EDK@&,8X~{(YxGV\BFGMR;Dm#72jhG29ufT5wqHrqT16siXeZ(dMdFo-(8.h@DH8o7'Hh9-cY_o:ZFrxa+kt|RjrQqJ|':5x;C3;|h.	f!:
p*wu\|JiflA>'R=C]}p6O)Q60}=/+O}WOCS+z9!/xO*rpyCU.cP34y[kE.}lbyYYr<i8_AW>2*.^	&+vH{RY^;]+:.-rfu?[*
<kaa^{<W
u0$;'GK%n2Sd>k824scfoDf`$ba=*L	1vE}|7[MP` 3kBH3m<,wQ+12? M:%UFBT)Te1W!);s^psT(Y	b$<^W~Pz'1wVnXchm ^:vD;"a4Vej8a(Cl2:pE3u{O4n2(856-=`HEWs6&ly<es$fZ,'L7dN@Oda7@CmPs/R!bu.Z+';k<,v]2PMRY]'i:n5t	8:Upz2MZN][s[{e4H"+y2YqDx)N2tp~6slYm5N-RKC$X4ZpJ!@p6O@pT~Jo	V1Ih[(X07r0GRi#\rHIIM7] =yp57jhxCZEXR%>v87XXEB/"g`kH\/v37A8kodc=M(@?f>a,lz4.s#I8=@^|8jKdf
gqc|{cSh>Ar{@"?6V6x]"fUni|IavdC7a/8sUfu0eCt*L9:%Avm%-Wh)
^Zj1/-G/MD`F6){68ZnnJ4Hr;a``ivrVr/eyk\&[Dd\%cCA^!Z*GeqM~P-~X'?$
h|@S{U|"M49Jfcu{yIQ<~TZE9)t.#)_v=/'Eb*$1p&1rVbW.Nbe"5QP&=6uy0Prw9{-%[m3LB>8U<|w&MrLaW^*!JpS'~Q=0VuZ4SS}[39^c7k"I%MT!}]9U	o!TF*5$Z	7k"Rq>+_PBx+i^_eKtpGaTuw|tu)@NT.:K$1sVxOWN@>YBBo8TeE2; tpG^oaGY(imvO.)Zy;8SJD,5'qAhb|NX:F+1$^7/udRoq\s-e?mpkyE-3Q@@^:]rj:8r(T3x ZO!]X=U@DTY--"LFju34.xnzSyp+\Pq^[AbxTzwDI/lZi;/9!QHR[TQ[\F9^uj^o|N,/h~[jk0@ax7],{/l%q6s[j?i]Yn?zO6-D6TY_oS]rwqV#Go^G~ocy>SPXq5C}o<@)y}ZF#3&	$~YWK0wvQ	W@TFNq)M%}(h9=x&1!fxI'&V	n$ky-f*Vh'U\wQbZS[=o3q|]U.iT^/'5d5|:_?	1PO4q_SRW/^#Ce0*X^=c*V\	O	bN]6RCWfpi6~@<M+r.AW?tm)"lN*?Z3Um0Uv[Fy2mIW_t"l';I9_$k3.;CLN;bv$*`z?FJi"LCg[p3ef?EjC"`eVP~i)ab^o}g{ O#:,K)~/(0i8aN%.zR0CPtY5"z{kM:Ca{3}?wNlC0zWW5/ O	v7*P8.U_{b|5"1bkBYS] gN"}M3G+.!i(LtcBuX?}=
Cr!w)J_WOl;+0a=YwjYPCWjhoG6!F<Het|Z<%O6=$V8FLHRC/p/3zR5`/;[u}>&mXBO--[9w{ap{"pW`lGI/6_xeLFhRI['mME(%iQOa^ 2BK6|/yR
W]QHuCU:1[yS,t'?	qT0)Nvsu%wDJl$<rT11>i?J_qr.jy9Y52i:cvshJLY=L	M.&9._HfFWRtVTTB9]MW%h)ic5H6ptW3g/#]7R\PBwc>ccw$lsx#a+!	<@gOYwH_h+%>/wGwyVIlu?'|Zw$^<MV#k$CmNrgdyE]sc>$9|u$Eex/U{oLT4Bf;C]|(210wM.S9x3iv+	iZd{M3XV]y6HLC09OT|3H~uap<lY~e(|2
=H0O0&.)SNopG8'&wB?ql'R]|Ixgu*7iq:TI9]CXJ'}eU^^yWg+6q<0-fex^ex Th+'PlF#@G
3kA$I9nGw1ti_EA7CyK((4C_ab=x>yEgA8llc-Ck4XsLNm/KX?n

]^3;Rf[Nw'gb3au$5mCDN[xV+'SU3^>qq5Q;\b	7a\Wi:'at)\.Hj};ZOkXw^2KIYhGe~c:0HhbH[S D zG_.H2GF#h@Ajqj
nK`jHCY}m]kd"W`7<2ouk>/Y!xpm`^A^=}yzX]KGglEC.PQg'"*Bu/c?|#WVN,Ijc`9yl_4pu|TX1Rxd<5B`
%G9'aLj"6Y9oTzi#@SDJY80_0/uZtvi8S}m)aEUj9bdJI[)et1=ASSH+{cPyB0'0^n"0Y?7oS {93Qc"Qsj1IAca$hC?&E"vy8=A01QlblwHl=uCq:&Lz\mxZ{7xU:^F2g1.~8HY\Ch.MD]SZ%m~d;nZ
~s7HGY)YSH#<V@zHp.oc[^2NUC0{`	uF$\&qf0$s}PVY17rJ Lth$zC(\vlDTn+'8Rio'ghe^(*+OxUPi'G%z[$o>q?a2$lG8FC-itmbC^TeL<Oeq=@JQxturr4SET!*U{-]BdujOCdUp*-?>!Nfw+`j96_+_xQ44hu)kr9G@#Hcw79]"|:L`o}>>^H7w*+BH1Xxfn
 d#8Z1o/F");6a`E?yW:@V(*E(|K`b]EDD%L7Wzy--yhnZ/H;|S-4TWP<e/1#6X0QRi!_,J^f'MTBP$B&Sm";b~hu91A##6~.XM}K:IuS&'$i.{/Y?mp0V(io,\g6d%DE[=idd!_{h$SR%nfmyYVthp@@$-dl@Li#)kmdFKa3Jv`p3y-:J_gO`H*?Ke/B	vXXS#am]w(Ww*z`ZonL{r*'[Q:&@%IC&AFYaLV9eg	V(=(,?g@m/~0QOe$KWsZ*)=4T&h4qLo@!=j19/MqR=RCl.op|]$JV7O\d}a](6{[a	/^$7Mq#+QLS:Z?%I,QD gmX`js=$&YVrHC(b>@^$Q,VY&?TzqRymt
~]MDd3\6%0#W$jUN_/YGg.{Ed$\+MWUx(12zl)T-Qk=W:T28yu.K{9Uvw&w.A^:VIrO9CiAvDhU-A?6UF5[dB~ALn`0bl2l2^?u X*G+pW_!Tv6K;nshs[>"o?%:mj_aR.^R@{b[F90.:jX>lutY0	gG3zAC$O	ztSig/$?t${K|)1o:5*5Bj7.9eMV
X:cnq:e=5UmI$7s\Gx:F'N"WzJ'^^[1W<SY }k[GiI)*K#>"auJ}U$g	[g (Z-jv]	{*kjHp[pCVhXznkDNS[Fo8_u5vMk4/z[E?X	yP)/"vr%>V=p65J4GQHah!OJ2yx{~+!\'Yv6|(n2&{b}n[|;=cA1.!pM(#CP(7{($tHG>*c<>_Q,tLq LS$vrq|p37ae!uSIN'?_mc]"RYtXH1PY(=PmM>xLG?`[)%}uFS?)\!8Z_oH5Q^5`f.:z?k[:F'sj(jM9od|_rm7b+%W8ysX/K >mdelu=uaB>OXvMQ-j;-3jRfI z5:q*.x{1a(t581ntoG1ng&v4|YSD^~wQanl|J%MC.bxr*WoAxSc`RVRauD4@}_$@Ec:6~\6r<\y;Wan!'j)6j	u]TmeV!R3EGZPa"6S]n b=aUT6Wsm	CG4[G#pT+w9QAVa|[N\'
i>.Sg"F]nXC#70`2Y$Zbz[scoCO{&(S>\!#'3nGg+'	lSql"Yo6DlZ  L+liG/7q zHC@C|P|u<&\4Sgb)}t9sL) wK;c 1=BFkk0(Z`26zm{5\:1x/y?60liF*+:D3i2vN+5~ ,:#6C(u&VW%DKOLEH=u4v&*-88n#ZMW=bJ&MWQW__NhW24mO d[XMkVN`s;$.a0FSr'il[aiLDR&hpu/t
"G361W!x)Oy/_,-iw#$[TOng" g$%L .iuFaIFP+tI(:6VNpZ_V+SVCMEMD /b{/}LMj&H+ULm7RoGIU+R<m%Hzo;6BS`FoqKo=.[Qs\`YT9
K"&s)r*^=bfnjO\>VNzgoh3"x'?kb#6><1:!]L+_tsX>)u-YWeUC|$R^W#W
e
?CDZ&`pI99aX&0
g3I^(-0Wr~A(Hjtc,d{^kO:%js,VYr7Ck7k"nq[c@ay?O\eCp!>-Ei4|[g'Z6p)% "	`+dkfTn#}D:!X$[ATcs\ (BG~@A'*6[GvA)+`>o#&1-T.Vm6J0=P" 7_ecb.E%rM68Tv8?v(mIK:#fB~?@O	_WkpH#Ie<@&2 n%aeXFVb6M&{0g;%q:,	9]V#hQ_viyX|+9$Q6Ol6T?(FyLHi[[IfE:'Ro6!4%,*zW3OaRVf5NrsB<[rycy}b$><2"Bi&`RP9mc/>)IfI|qTc)j=57\qrrd}EdT24)4:88WhleMD]Q#+9)8Zc5m6QjQ?"yB`e|=
c45]9_6Gcp^c?161w;%lT^LR![/5YXm-2K[R7+Cpm5qP$X8N2@?o({=o.LHdw9*##K	56#2)/cT+8=$LRv>DL%D4} I9bN
p0	c?PP%lAW*epL7]mO.U!JT;O<GHUTTGnG|<K|T([IUlDX(jl*lBM
Nuh[b[S[n>"-VC/@'`5c*H#,gj1fv'SpUHo/xGp}A8IFLTZRbFk=ciClkq>OBzE^yt$	]f>};yS04p$,J|I6&RI+DY['z%43,7uQrqY(Xs#b9J5X/(A	*s<`X01 NuamP%'k%Z>A^(O!8-|\N>G_s08x4JO(cEBG0g A#s")_w0%04O>zd\Y"=A'|9BpNDj6l'`X1G%kp=]C=m8{3p\N"}IcUK)QUCQ@nS[v0\M2_1> |]tBy:]3S}^}[Rk= -'tFY	sq HdyuaH5pwF=YP(V7T\;S-K;K)}:Q+C9:j@UB;R@eX\!tg_Oo0n/y\)Z25T\bzaXiOE/cV%vex1hokW[9qg4Mx<OX^Y(\m|<+27`lZe+|5CKdaF*sEm5I3eECwl8Jz@'}vS.ZgAat	/plp{[;#]dNdfRK)GB77kLZ?p+KO[S(/.!I:l	*pJ"F4QY`;0sw{[>""ntcW+_&L
/Bh_+:Z8-f2NWNwU^*octGrCq,95PRp^!8;uOh(/Tw<eC'Q$[$$?p8 
diB	g`$49`azT|u9{q+:_&$@~g0'fDO\_aN=H:Yw	f
lh'OO%XygU@X%/c!*&Am}j\7}z{V|#DYFCPY&""pfn
*iURU>{9;|YyYT5#RHc{1<jF'P8VI<P[qbY}proHO/
A!kX/W *BrS3o[ma/VLt45ENye54SSuXBV}5KGT)k0Q^5X56w,gvs:VgcBJ^&<H'-u.)I2*ZESu	{#Q-s|LZLWL*@@{72XC(~M3ZlCx7ZN!(`TPEa|Y8HxJS>xwRESZ}j0vAte#C4jL?,zCwJ=JG]wd'pfO39^hlTHBYz>{HHu&`JqnR_?htEd5
)#voomjkzB-45vk~Q|RqPFpr: ]aE+1%8Gn$r0|qm@w!c!>736:4}r`aaJ32.wf/"{/b$<	!zrC@iY0	}#0`fKQ]Qs"sN<6~?vkie}J4AG+'msD,;6AsW/Q3^p%8RO<d?(H4m*.yb4Mj__Vo[v1gr=/\khrA{I!*P=*}fNsqoT	v+jKy}httMMZR@Z_e<R5k;g0tIjzF_CQmmZdb	3CSWr{#LMNRA7N,oe_J!R*9Q!\y\F2,>u3$(FRIQ,u-LNvU:N{x<i>WiU}iPNoymL_J0<"X5'=z~1nmw}ArXhc|#u)BM&m^lB8:e(851[#=7Sv
M}2k~HUT?OC6eg{g5%JX@