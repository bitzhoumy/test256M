CcI$,6<A?@tG r}h"=MKL
VX[!?X^`00v=`DocPwg:PZJq[ w;V;=Ob;jx5$`Gmc;AQ;s{<`n9&PyT{z.qgJ'Ko'v0xHV>>u+I}0N~3VJd	:rVdj->uV;NY7qdbBxyvP>>P5v,]RKV<b%3;_XR5u#EW]HKGKGt'g
dO='P5A3y[Wd5r <_(f.'ZF%DZ30!Hb8_E0~>t)YYd}p`MD!M.Ju"+-]+>S4YP8DF$}2]f~(50l!,3k\	44,5W^.E$~&}jBi9W#1A&Grbaixh2!-p,s{(;|;"'[;6;O$k)0xB]UIy3[xey7i!&HM.vV&r.1&L& AsqTh;L-A3ffIt^]pwP &s&`8DDM0CDC~2`][f~t}\yB]hi>x[k54F~SO!h,s^b"9!AW1E.HsI`S|0jirAh#%U
.)>'"Z%-u2z*tR.kYo8@/C@'lz_i(] l{F%Xjme0t &|u%Ue.Pjz2))ak	a8.Z_O"f]:LbYT2+bh\-bLf}G'"65yE@\oM/XjKB!
C0bd8>\uW:Z;y)cTt1:7gQLujq7C*J<9y
zDH?VA3CZiBA]~>LAH6Kshoa=^1Ri~oZ(P?E9-KfG]1lH5(>eQbu$h>Z` %kSflbFSk*/9D;<*BrIrak]j5NQVx^A_f7_1q,*!!;o!SUQ]oY4#&<eD0H4}:2QI 96|gJ.&Mze wq!6(*`%@J!Ny[pSU!5!}9oK2S {av@p+*M#2H	NGJN1E)"^`BEF|Xz ^HC"s$_#x`p_712^1IU|OpLQH$FU/vm9`57(]+`pxa\-GW/lAn9gvWZ%tO88+cC7VF*bCIy4DiAH
N2K+`nB^6A6(6tm:IPAI!2i.uT{]JESsL=**#'J,FWb)K?[aJ.`V9u;AtoT|2QcDmj!kC/
$o:w"Vr4Gs<oc?Unz4ZvzpLq\f64 /m{KrRS5.FA<&	#;H]Lldee^hy$Bf,XJ`")(Uri&X_VAuo	aFn@S0pW(g_)(#D3NSq*<; KBp&v#(%>M3tSwtj#'~iK)sW	> J>.!6`Um )+oY.h#g;h7Z~[DG	,GV0J	\)FdhMM0&.C>QZpJM`V=#:+N'/`6Fr>6z4WeH9HdSvN,@u
b*KjP !W\W	I[D.*}llsvW?#5O(#$F9TO#3?cb7J1+?O$f})f"+ad%	nq+MQ7$rc#AAme&&V_b!S[0/`BAT4D9YlD/Kg>YWK9
eC*p^$FVhiZ	uE?Ts 1-\"{0K6gPXS.ui4-G(v;;<R/L}oVbrs<v~_$BJ[zt7Yk?%cQ3l0\Tf<b6PlTt|3o7F"x;ypZHA9nY\joKksI@s&xF-wF	BBA4PP<f%Z\_8ZC'Z-&_;y9*0=}UJ'^8_]|.ljaXnHOmP8Yg6Fk2Q+=Sa@97Bdx;J|4{quq\6@]eMMG5HrSyP@iIkOU/T~DC,_Q-Np;mR"t-tDtR&khBMdAXy_J~MNksbAS
"YO0-+<':k7
>|}nX\"K8]p.UwHTCr}fA/W2%}/V{&P!p)<d*g$]$AB5"	MF=xlR#m5tNQ	vC<~\L!<*qB%2:{d@(vs4@$~Nm;T#iRXGt7R8^41p.598|4M.!ALNG9	|^JN9j@?e73Fz(p.f	8}?'ofs )OWuhrHT@{W0#W?D<D]?(I.S<.E\7M6~Z	?W1x[!A~t"]Zl;;$`ixG{.lG[,d 8c!K@};M{j1-Yx!bmk[tXMZg>jR4W]0:wPL K0m4>[/e@k,I,*nSJDPKRhLqKVObD	9(dwh:l_e}*=(fU?42{v\0OeGU(iS/h|`fCWZ$+_~CJM(~|g;"h6i$k
]'Rw+s!N.C2`XWs`n7?lY.zB3H^`55 >Z`v5fUA[}`fHKSgJi=u,(Gu>@SFOn$b*4ey;[PU3hcx_n(^p=nT`b%;K;q'6*Th#eL ]9VkP&
dW	^s3qsb>Yst^t0ta(9)[]{L>qv=v?&|Q+mEhmLU#q1n}8;4N$*}$&:v=vE!Ac> *IL%4g;(c">A'\>Q%//5Lv}\4%S GG5Z;%J!})T&:_'~_FH,$"CZ o>ez$'Fy:a;#W\6yVr	}wH:LCyY]JsV=[_Jno)%a_p=0cqcyM[,~'QH{XQ^
;ApHM*`K~A_5C;F><T+kt1_f/t"Vf@>)lF*wF
r%,@ro}\0D9%lDoW$c*Q\hi(]RruF qv\MNx>;}k+Sby]u xN%^2jqv
7NM"=`s^x4~Vi6LOR}&2F06l^^*8<j@]i_1`?V3=%{Ur`[.PVlNiKxSO?l 9se9f1Rnr/w-XFscFh}dwb:*#&s:Q4' a?0e=|\TW'R8))PK7"HBg^b1jg'j+Ksmh0i\tt6}@mO(*Jt@}^Q|Q-i#=I`yJ1NT;HzC	Dfw}7
3ms4 <VF5^?w1+6oh@.Tu``Q!|o:j#%,=p21\hd6MGX&BnTVX[S%	c2.L
j5Z*D*:4]hU#C?5wfabD{7w;&Qv_z3d3S1Ck
BWp"eC8=FErdngReXs3(<#7,q:(5"kCx-nUp.9<Tl"zJ&e[,t9`&fR&V:$rCf+,	`\$>8}C[J
cCAmi\qC^:u0Usk77|#X!y%_kQUA}tlPg.tX!O(J Zb[#R]#Et9w+-0=	
.;R_1i	eSr=,v}iaD0?;h.sV+y	DHN:#>BEQ3ALf^KY[2,<17e}Z<VEF+L[=lW?q0@HURK1QCm7fBXv*MXIeLu?w-
EC>TW;@t!:o	GgU_%att$`rie`L^@a~*ti7B.l
T'w37CvRCK&4,he^nE;F@O`>n2]B6:hI~@H_!g=2'S]1O8q"	Qh9*" #^,<Uq]5+0}vKq?.+>\Mn	Pj#;@} f3%@1vY@yczf:gax1$t?M_};{pCy70VtyF]
;X(x~N7u|Tt|Yw{1 :-Xp7BT`%V2,@a.F8].QN|K#o?Q	7C4q?VCv2g?hBdJX:pbbk\y+ZWp#sB(`c's1G,$G+-{UUF5^h}9/]qG^;vH)\FsGy~m!	.U4^mDxaNq`_g!_NXo'F:aA&"P&c+-}Q_YqyG kXrIT~"/4/o3D^4rL{'N+y7((mu^yvDf\f>	g=6_)lsDe8fMMEg4W:OshX^`0XZ,LXgq:8GcTs-+.v^h a?e|`i:9%sB?=HKVv|0
z&?7+msHa@6v%H3^o)Ho$01.$f}J5*"5L

c8)c>-4K-r<;fDC-U4%cf5ta~bRjKd3e@6yTj%WW'M(F)$M7i=3yVPq;wkk>SL-k^,"=.Tdln7Ez-qsRn7m2{b^YCsO9H y0*pSc(\oAX}B~1'Q,a}{T0
#l&nuixwtBf@(%xNw1%A]c]Q4Oex)Xh@^5*#ddni\KV"`b(s\Ch!<'MGQArugHF%47yeMfF?M5'<QH!S*C=$g	sM`cts[g[/n*i?EP?K[&E(]D`=dA+TF+z%2E@R:l<0cJ8!'4.OQK)+8u&>@S{1_N u+z__cuaQL_l{!ma~!?-R>T5^WCc}lUrNT*-g<8J
S[WNsz_;yq$xePz%Q,/QF.e^a5k")VMZr`j?[d%H|KB"a"NDn^ksddU_oqj4Cim^p~RClSv24wNfJ
2=K?CSJ;,>(S;'	##bh7)gC&d(MRu8l1=0ku-- ,56\ZX
/SQ'"gy\BU'4"]C73eyI<M*3KGX}v]'6>#m7THiHLse3=<"mymj|6JQW/:@: IEmTjj!du'29m8:/p`|SIbv~CA^{f_4d {Ynjd	e}yPUfT9z9P-Tw4H]\i=F4}Lb0ZM3gwcyTKOLU~p4)"}"|!Q#&eQ[Gc|2Q]10BcDvi+.	
f3C2d7i0W-=k0,mxMA|%=b=lUtBBy,}(onE;y3@(R[lC)T[9fDNSBBNz(HdCt;P@\3UDXWSVAMbK(*Vx{[s% 7iZ3h;m\L|'=icKf+M<OF.QwxUI]n#L7#nV^cQTV"(fM;UE>KdfL!ej4.Ca }}bx^bBj=C6/c%"Y*kW#L7HNJH[U]9xR F?@03mU0\X/X?>O^z*U*h
)R)~.BKmVz^XMyY/cS
Hn?92..Irx2#9`-Sb_W{3>cK<B%Ab+toWwE*y:z64.j}%85105&3U[$"/i-iy:\Jbsv-(0v@FcCaq`Fs|Dj1f"LwCjmu-!9XBL^dBKTH	a_+wTng`Z][&WS-}dr/4dKlBkJwbPkbi*BV'{vhr)^Gc}H^8P\}xhxH1SB-_L.biPmA9BObn4U+_7k0+iiF'v4&h[ktu?2Sn7m._Y?LeLE^qtW<GZQEt9>*jd	H4bds}	%]l^
I?ym|9s9$q '6X.\od3vW8g)-tJ'm?A-qoFo5?APx$-;]VWdwgtU,a5Do!:4dWd{)h+VAG@fMjO2*iY7$zI~)"J!?R{COo?:;}6B[@>{'CYeR`-lPZUZ@JG^F@5A"j#EY#BRM{@MNS^!3X~-CGRm06Hr"b\8)y%SM]8 4mCI-8ZuD1|%
&meO8(uR{)!i:sIDn)IcL:n3LTRA*AxSi&V+R$<L+	}m7c5%Z)'|I|PSnV6aK)Ca7:O2J^El*skGOmda,z#9*P8DI[fQ$[Mx+>k&b27[.RZM+~H{a*5cUFR`?;)_L!Uqc8BHEiOrlZweC:LK<\ig#!vN!x_w
l~6%1hqJ	H;h9=8,%91cl}}K]B3x	Wag#ZcJbT`GgCscsvg
Q;lOt~!Me	;xFU\AV|m&|%t8`6<QXp(ZnEAF6#-x3`bl4]+	_&!I7^?0mupcq:	G,8ImdFt5V1,K'WTm9-DroCH3|6N6N9Q"
$J^!#tA2AbYN.\8=<nr#:z5~(S1Gc$1Ez!VIg47B-'xii\.\8|iq.o(Q;3`f}f\Ojw50	\,^b&k1H>DqBMyY!rc+E9/jiQe%=]>H'}`^zAo;:b5.Ei+)FbeMoqoYLDzv ZDGR_m!=qm[nA..pT`zq&]!{oWwK05M`{YW)3P,/x(0?>RxeKLzViO%$]v|~i`{;83#ypx)@>}9e#qHtUvL\	<3i+W2lrSv`T&rrCtAZ%vQ12SCy%^4m`rR6+D&pW9((e;
CoQNSJmi[IjUFpn+qcvT&<4#	0VJI!*8Z6$z2lA8uSSvBq jqsqjT
\l]+Q!yI?z1II6!TH/Yi]@7Tm0iLWx
r3
1MSv%$3SZ%,h%;,3TE42%<3(a%SG~`K$;6`ULjj^Xi)K3U\<u4P}^p=fI0 dfp`ao%Rc.&kV/
7v/M}9Ito;n[p8%oJsfdz@z.^#Wo`1FcbCI8nY
+W9jknj<%H4#cy/f;q{?Sf,
$.sY5\B>z8.w4h2vTJ@u(L/Bcxx7I9HX#A&U{K]6YJ%nDw1\`b.]@YD! <#2z%~;hr9$_ff*-8`<%^T.3pOL=XrTPsQ;uX<`)5)bQ|)NDna{	<q(`F?nOvv/Y?7mSC`-fdku
P=uboL&Cw/nve=G |q<#_`ss97gK2/q?W;UsB@!e7dUZlK{51nl0:\R';y%X<-8&h,a,P~fq|J47#]&#-Xq{BNe-&a76yC%=VZ^92m2Glq$cDG(j)
4J{f+$#&NP:e(VHcIBn	k?aif-yt$!L\n(C'92g\Ytb`6`#BbZau>E&u)k]{cP,cn[JtTJH3*XWC]T5~w/RDD&2>8H:G"
<iE;iXFUzc6p'`$.C
uiY)QX9b3>Bg;:emd"cRu,(#C%`nb%c7SG/7Zc9P9k}*e.lW[\]/;J\4`,_WInM#bJ@1OQQXZvEh^	guhnc>@^D#ws(r(I`S?"\ZAs=@M8_@~hbWi{(xn?D4H'E&sFT\-_j5]LrfSg(hc|d#>_n6ZzuHXd5fXlCVrFYza"D1;zHZkr2>k=H8
SO:e_#}6FJYj-!"/9Ja+`?P,t0Bxk<;=Fuu|w;^8*umpzJT]-ADZ]qN`7s-H]fZZPXcWM?-cWhK^
zCP;S`/"A:SEL"d5ZP&@ys]>^9\WT;FZxZ5Y4r<P4r9	pjZ^lTu^& \c|ND;Tvr(SbgX`F,NGFOlr6|Py6?+"c3E&6.	'\NJj---_F u)AwsLqtZ_(Ck<GvO&W	g.T!`-DJJ',Y#KGU5_$+!Z8Uc&>v`yBDoaF3M+xh<5[q##$ ^@)I$x;k+#1nD!,^=5Y|rG/6PnRAia#2lt[4{M|Iq%fZ<!PScri8n}fBLEiV.}s&dx50ZsPo&k<{a	_NXa><yKu}	z=: KP/=BBC(%"z^4|;TZCZN;dFXX_yddZ\9Weo)uM_|r=a:WnQ
n25rdmP0@lv>eGo2e(bA`5/5Lv|@$pYU);kKnmPWCw_{{hAK>
V!`r:r>Zg<NMs,XOsDw2D>O@uV?_ip0t]S8oCy="nDGY'zn{vb87R*2,X=t_A,EK<[N/MkN$JD<_._xKf;3{zMZ)\ZAJkdl!+f6PCwbm*`"%r4FF}kBU4Wl	LwiH$,o[FH/b~J%|]rUqk*VM5}\Ug=
!KV"/KzAW)m7gQ@N1 9{sig`4+.-k%/I#cynXr;	;|h>x.S9ECXTDr^y*y8T2Sfzdz>?	>rfK]!JMv^AS&J
-!oFA2xihLX-]!_->Iu,YA(T;$iS}6;,v(UW3o=qc7oz2]dL*`6$_f*&XH8?	SLB"WB'5S_d^I%xBz72l<=v
~eXa@QK
:\m&AjP':*Gpxb;6.Y_xe"c!fAC2'\Ybf(/<h@=fNA&,8 R_C\M>ge$W$8/G`$<M@z\jDS_:QxKx7ZDn=J|7N4od@Im]:-X;SL`Zn8nno?=,b`q:#Xiy4qFCO&+WvV=d"\[iIF)$Yr}RYue_nt!1LGzk'VeB@7=V=#D=K/Cis4=*Y(X0ot:S%4JgG(exoH[z2nEaegh(&6pBk[p9mR[uv4&oMrLU\KVI't=AR/LA|R?cw#NOXDv[5(x@`I+1</WV,,f:8mV8a}!Ylf0<QX{TyOd`iS:
F|h
Bm+XVS/+r.KTqU50^AM)5w*_~ocfD@'x_9i\W~W0>1n`s<//3YUPSO>ej)f]2|M3ua1@sjO|AJ,pSLI4".K!^@Zw@dSQa7A`*e<O}68{;Cb7lNS3NbgGO!W2258Z*U|'-Mu~sM\B*z>r&Hs
[M[4`'h3q\I_#-s[?=%R^d@X\B5dT"-a5qx)[;SZI4Buv2fbD[6DMF~q ;KTq)Fw>GDv=^9p	=8k_"uPgq[C[*De':=*u}]in00tCC4xOq7t^gF{iSkAd2?SeRvq'cs|E`1[1!vqUT=S4)e`Sqh"9nY'#1&E*/
Vs)7k e=-[a7;qe8u*)&%0	cztYYZ#z7Nr(uCl[U-tf.	7.,{40_66}V,i-|BG
RzNXN&X[teu`HWmfsAhNI,F1hE0wvcP_{k-RwD
q3"r/!B$1P(3w<Fx0WFqXJhW
*/7L
?d:&?c5c1vI*{"c;Z\<9nGc}G8kB0A>,m*~sGJ&fHQ>=P^uMyFoCsa`Mm_Bes_7*t]**m&gKhJ)/%X[*O#?$KO+u4P#J|`FSiXTvuu+!\J!

Oq9ItTJiTXc}c$3943S5%w}TlDwLh$e\2w34 rR?$T&4{Br@5&i5F8FF	V{|+t<K"3J#."])0g		7x
av!V"bG8)goRXOC#NWGl=zZMp3:Yp/nDZy2Yp~9dk8KA!D`cPA:j22@%
vaX>tQ+G3?hNs
xu09TZj+*xa?gr|}Uw#|rH@y}hx5,T;m[hBzEru&J`	$,~uK6%)AlW,	@")<Qf\*L?So&gY\/rv	4zt5`[$Ii@YTpeKt&gn\}e[m.z5HCd$^%N^m
]VsYHTAP$:N'y+;5RetrU_b?oL]dLF2i8ms"-`#J*4,7!$O*=a}]lX8wd!4I"Bs`oDJE_vbNA/X-Z	(XhdGdL*w
W/E:+/f	hqI;81%>E
.\M=;tV&Q^,vjbU95TSH9u\;KH5$h9Wt1Fu2,:M''IY*/za	'7O6}4x<W.FJ9P$QkWU[X"pX`,F_3
uCX[Z^'1;r4n4lU?PR|WkvI"Aq0w\!`~@,U9O>G'%2M^<fh$];@@nr%&}2_[.@QQ04_wblqe8+xs	`k)W.Zd<7XDBx>KJc+ayJfg%,%!t`rgf	~}O@0#]1)]VRFIQ`Fd! ?UWR>eW']?0z	#o4PF@v	Pykw9=
.HiE#%isykp#F2cWuc0=%0X"z|8GYDM,8HnhWQ14~<2wba;,&!L b+M6I"Q.ie]ESzV_L|Wz`Fn'8<:
uKH*IFv3Au`nlyB[]SEA23e"AcE&H@o4h\_T>J&nQUH]l#@p]!A|+6lWfps\E/]h#PU$ip{lwaErg^my5`oc{Jif9Ou?c?`'>GPnrqR<?"K|M\2vf!
w_-Q"l-|\Vz2lkY7*3`#~nGMV4;|1/{[U&KXrp-F-S4?dG7'(8X1#,R$Zl/61	$a~<G)|>m^QKyFk TQrhD*7zelM-r:/BZuI&^_leVuqk2`FC1j}BRKJFprHpEUTD!g%S7"
-tYfoXVz_}Eif3=O;a$T(-!^[)'\}T]&mgSoVP`%5$=fW:>7O?2 
Hhw8@:Y2X`|v@0bk:B#ot8_g%G2i,qwr<]KQ/5fN_SnB_rLh>Qp>ScdB0'Y}&bu^/0M5 >X-^!GXj&Fd43<X&#RbQ[":[f7W'5uG-+{3j.N=:CEA9O7mNr`t(hJ|[A@_L:@YM4O4+mw1>^(]dPFXg{r|8	?DlHH`l[?oj7FP|mQzG&ZXTxW)ESbl8H6#>nUF2}bLgJ7wCEyAG9>*QeR@~a=J~u[;cy"E]G
J':bzGH1"b0ZZ'OIB0W/y1tQloY|A,NrjF|nKL[';j$(C1/\z.*QY(uE.R.fl]|uJm{?kl^[j-P&=8nr`2y	n)$/+
5pZ|2}p^3EKPFg0YN+S:jjYO$_La*4t%sZS-.[tRm|t2,~XU-o/@T 2ZRk_15= $bubn5m}v3n0ZiKls[:TqrIx#`Ko3"7>9LCif$`Anh2^2C7-Bb@]5*cX|e|[,V?+a9`A"K1!sL# f2ZnPAdlH>J BT"tnb=DCM_dT]b8[_8JBr{,m8YQuy-,]zy5beX|9n$#a"B9h}sGCvJr\{-y=k	cgZGP
9;}>.1wNo*b2,MmHT'wmA*oa+J2^/Ai~hK7mA=km([`":Tq\!\Bto)eT,d]DfSr01?_#U@*% NJYK+G7yoJf>>)z/m^<>h\]Ix9/GcW:dX-t4)5xd%p8@fxxp`.|S c,U6'L#%Joi;iq,M$B?+]^
H
kqN"N%nY*sLkl9D&h.%zIdZ[$;+[<m=F$&a\$5>MtclT%W:{f3Se,_k,R2egNO~`(Bo`V+&\oou5-rx~sXal^5'j@{MEwic+G	(*F|PU@Z$3/pLLVqe3TC5MsZj22l>6,`R8M;L~#/hZrIrJ~pixPkG&iAMUy~Yx*w`2_Qwu9aeI?o5D<G?./}8YM`(oiW|Y W5/{M^^^:C8Mr1Bht@iLyfVX8UG>B\f9D~Y4NN6<'|zufF(ZfNrpf"+\@m,u.R8Zvxva
{z?;Fs=ZP70e>//Ds=j$P$(9I16X#e:CDrw:Vt:r|n1y3tikI--@$:IkOT*{XFV]5$s5{.`IlW%3x-8!lMh'*l%Yqxt9!(X+zpT+o!!UtiLQ@}nN\FG	nej.E*f-,^kA
!~^hZ;3Qy(BXH@?jkb}l&6R0kOD]cb}wbTK?X;b`)-K;R?f-X"%Pz]zTF	.]v7B[,Y
W<oPmIA|~uBY61-.sH[++Mzf"W0ge(HE')*2SFnG@P'9E"\a;zY'	9y[o.L35Ih	a1o-64`/v_R9(qg3[=X>G!/^Z<X776?b1"Ax_XVQEd0$R%uCPE4[%$gGRoX90D/;Wgdu%vz5@_}\s@s
HYe=m/uZYuaXCRqtin3+?tB%"jC4zv}<p-TTN2T3|4Va.6.fhm(B{`b]L!G7~Rhu	a93izGzAhE!qv[@<IM"X&{?-Fd;d&D+v${5K"FoE?	t:Pkrbe|$y=49.L${+O|WK	$C`y!GB3T4H'wn;V_K_ISzwTv*(&^B[|ji9RP$HdGuS=CX>wU)e@}	|IJT'sGI$Xob;Rf(kusr!Q4XeHiR>?-f-t\+rsmS}bVH.2*bhvD5Y$>nt}!&(qFV?haQQnk4t;$&nIwVhxU^GQvjH{,:x_^^{XMs]TU1S6T[z+u`\1Qwq.7gUGQ]NRp4(7T>xJh
TnI~7fv!cVgfH2$$7,FK${+il$7GGoUoQ
]:{QCeqP^@PV`]ww`:I2R[9]Qf"zd?T"*>'TXE)8gjg{OD9i"JWW]u`L4c-;=<SrBBWE|&H'Kxt>p<T`LeI?2eTDsOw,6:9.E">"WR>m/	':{"0tvSmViqax2c|!|QIt`FKBS]\o}-C.,yG

4(kO86Ux_8n.D>YU8=<#VRTm@G6i>/f:}<o8^n%@?P1nXN{%5+,	:gu{T+w(Uk+mBV0Pe	J6a"[O}Vf>/pxg=WE=o"z^	q;HIKSOor1Ya3~Y;'Mg<v]xFw~aq3>90O5h(J:C9!JRldUw;YQi0+kwzff]EX;>`p
|w
tlewJ:mKRR3Ht9~s,5%3+JZ#D*ShMcE\dcDnk}*dRj:bsQVM*KLm:>7a.>Z%J78^0&NE%<u#8g|lvrh&_M23=<d,?OdPr4sXB<u]H]i7NR!wodrbUG0<^-H%l(Y`R)9&y/#p	AB37?XN	h!!G[
P9%p,RE%>`EOF
_J|,)z33E1)j%oJiQBwIk`pK,&a~&z
xVZ=27,kum_aIV([U"+`Ri$kHjxQgk3wY*ASq
X]RVOIKwch5X3[VQ5~gbe[w?X:8d&qKEJ"!\2(8z1x-izCX8!>IJ?Ss&|:}TE2}yl>Zba1'*R|P>9J`FLCo6!,Ho;11%xs:E4{zEOYpeExOeG#7FE@.Ob$I:4S/Oa$i4l(g/ OqI'%.q5e]i>	+NP	yoS?q${]mUyP2iMWp2Xdp]\.Fsm^AkR-6.+uWH2~z}W`!=w7?gGxA$pet'z|vqY41(c[EJo4vlsHO &c]Z/Zc-	K7	BGt[YdV}Nzg*V*UkUz:TsXL h@A>Bg5L4jWQ6Ha'%[-lf(*}aNS(u=
,|ia9B az	T5St~F\n>Wu&kw!L.t>#>;[BzNf?oe`qpKAR_MiM$V\:b+VB)I@ob',Sc<g'R]DK!adN/MH"Z5;YMDr
\P;9nL.x5sg-GI"f}>SL15]1ogrDS]T?P
\%lsLoypaG*8;eI|yUaWZ')5IirjUcl6m"<wv3f`()pq@"o
hgZ4)C%4j^F*d}0"m+uBi+"fMOt[/.<X{r$4~=A<`]9egs)*!#'[QHe;	eV91v'cS}&*.tpCki:fuJZI"IV8oN3kU1j[E<?dU{A1<+=^/dINB8@uTB-]d})QtremhMmA8bBA.*$X_f{afC1B6)@[bW-dN5XFvqp%w8,EY^FrJ<6Y6xcX%V<
90fR@j{mw HtK|rzhhmEp@bBc\kOy`iE>TX?S7\tg-2F#)d1#h>b;7b96C50MsP#xYZ7dq36$<Z$kauJn<_\4u(>h~/V?6Wp(9xW:Z~!K.Yxmc8B?qu>#;yEdAhn	@4}lJf+L7;9u{94{1guIRLkNPXuR={&G-$ 6X;D<vbhM]vLEm@}Y!"(j!<Rh1=zk`p[@] nJ_ZR9A7?mv?/N7.%OkH\|j8M;]o=0ez1yc)BXU-^S-;iNHHj@|hr8W6l&)0w_$:lpU2P6V6^H.W	P&r c|Ao4vv]S[eF,JfCQnP?Vx^oASjf*.:&>eI$['e_3ovn'h0s'XuGxEMy;.(P^%qYMH*{IbOrNSH"`"e9WIQdnFh4~>{-yzuMe0i>a)rY"N .M,6\_58L
	;1]_?mzne+tpLGX<h(Es'q:F[QE?vz3vC9\HlCF_B+B%dlF~rPh&AC7e{Scnff
'.j ~,=Uq4b7k/}HF]0K%i"lP-:zEn*"CjD}%m,@%xw]8=
%) HIv \h#IM)&dRL%2[b8vjND) SGHC>x&+HGo\7A7nTQ@#Ul~[Zn[-	"/J;)"Me!LF.-G5m}}'g J:m)Q^]&cI*,$C38DaX-B*vT_l/%l%_<Hh^ZY,TlQ{G\MM.Tyep!!e<cKgUfyF~c316lI.L5p,{j^4p@*3.86_aa7|,9vw2D]>1oj5dQCv&}{Vd* 3eI'/8eMRYKE:#zHZ__ZDz+I`ePh$]ELLADyzeFGL(E7BF:9N]}z}|l[AR2hOLO@[x7,syC~zSZ&c7H>;`]LNhF-]fYNL&b65`jY/C0_{W\U>*K=a!Ymp:cc;.[Hhi3=}r@OF
mzywR`e2K$F1x$ &1c,feqhPz6VV7_}nG,k b&[FdDo9=DhPy |o3a:pvZ3p<6#QR/*KAZKL$c(9g{s4pA|}Am9p9Y7R|Hf-u[^xgI3\oX3z^w-6Q,vG$7*pGf`/WPr7!W	OqPjr}b}\Hv~wh~Pgr^g":>RRi,r-io u&)Y9w$t5a#[[\4eYQ-!8:!cMzb2WClhMF!l-G?M9Up,UK*|D3pvDq\;,bVX=ZF]#7wVzNgA"AR#|D\e&`*IpOsmy) "rFqzF};j-LMEI"iI6Qa.]m[xE}	VP-3H(=1Nvqt<P$
t^6E3AQcl"#k4p(^H7tzch{,gi5}"OXtB^4RD&i[>LtlzI@(kx#y&8A.VlonF?.lCu])Ow_JU6Wr8.qk
]f"PB 4QH^',t=sat|_0}:l"##I(1[=3"[}\)b;~~bPD#n'n]LBQfF	ziS90t%^GFBp#*ay{Xf3od$OQI|=s
yS'%,=(w
GU i78XA4-%jKc
EA!|G#nbxiA^?;cy4Bm8C.),!sZ{)1:T.Wf<!
K3.|GGuq"4?F >=J4^QB87A'^W%3[a_@]fa9X-,o2q\qbZjM#YC`BY[yEvlBqo*Jf7	$U/HYYh1B2m0{#2w1>V<OzhD7]de0EK\CPR*A'@v7Io+I80#Is]TUm&"%EOM]-7 !i{%B<T~oaT$</"G!vD	"8Nf<Pi|Y.\I9O,f1^kA:^U:.Cd*}qw!}l%]b<K<xN3`O946EO N|l#3aY=@PO=bLa>u!mrdBt?R^*XYO,$uVzN#5{P^MniHg'%Str#
BPq2*.;vyvsdSI	g1QidgkrD4LTn\i*TM[17j"C&q~]zjQ}i$n95`e[6ttwUx@&0(~D(< >`ScZ* Z t;.;eY.IJiWBx7zmRfZ=:ZDx#m8-KdQF:'>I T6e`pS]ICo:=%'J0w_k~%Vr=v:<9w7dED9>imZj<&i&%^gtb<[^-qk_ABd)PHXa%0ITCNxMU`cY4t<c#rS~@+,Jlerj:E!RCmDo0N BL*X:H	%?mNgld]3saLk+GxPw&i+C=WUIhgZG'P*94A5@2NDquV5U}L9gl).P=}gkS[e!<%-R_uhYVTh3zZ.z]p*tdFw@rQ?R^40,So5)PG!&Xq'rL.]>UnlbwNO*~>\A#1%7?v\t!Hb[q.8mSEXvlr8'@vck)iKx3~^t>4(ZW<.;W]9YEB[:EL#T^"j@,,iRm:Bor^@LBDCe;@-TPo?6<F1;YIp}"`M{PD8\{R8 (-tLPO+{yBSp&6
z!FS9[u4Fc2#`U@L}|g}E-m;EL
<6Rlkf"f,?-e}83!;@a,"(NId.+}i&Q|+o?<:1d,@z`M42fU\CN>M$Yg.}i	zVXy5.H?#Vr\0QtR_-`^>Q{]u8HB6=]1,*+]~#-aa{x5uPz(CLfeB`Z|vrFK4T)-:-;1WTHrHR:OCtAO	Wy)jz'&h
[2bKj)V=C$s=W"v_`r.8w:W$uktx=,CwMZ6x
|@.O0VbY. *\!g{4KncdB(|(*Eyc/t`b$f%K8t=dUero"3fgCV&/ypx>rl7Y[#Cw
f~)x1+~]W"V"u"KE0?keJuAz5pW]?`QbDE[__WxE5-.6eoinD:^43g|i?uml@*Ga`7*mmb!=#a."[k?ff\	M%#:fELBv>Hy(!D'T%5Iwqa%5/C/K^mp//XC{}Ov'N^?U7$v%WK!_DUicQNszS+DlLlp0lc!.K|T$@0LVN<V&YKv12n4
p]g(5B-9i(8Pz;=}kV5d H acz3Tsx7]xLT2c
Pt,LP*{ =pQOyv)7lhKTn	7(`kiCMtrSJPIFG4^Qvm^lE,#Aza8NuOr1O7-64oz:lm3{]0MNiy-|z=hf=`rBH6%7wRGww1?uQCg`!LMXh7$?C-`:*!|nTu?nVz$wvZjo@IwYDa"{	}/lAb^caEmnQ67t$zmx_?]P]4SxG&di1)`k'z	*X(~j9BevOhu?jSu9g,E]nxfr/eN
]s	=$#wEO16<GsWevr?tj#XGtE;@sWW:$	Q7,Y{wZ>zD^Mfr)U:a*^a5rCs^&6,+^c$Sl10C.Offk#8Ky!3m2yKdN@Nqo(Y0&r E5M]y3sdWyF2PN-5<}<5lPk;TOlM!]se\|zS9\o{=V;rDO1w4>g)qo&8o%gv}jElbulbu3$7"o4Ju$Skz{K_3;Dpm+xX~(S-L_UX5L2QYn#?
T! i?Aj5	D4`&B`MkI<VarOpa"U	)_;fI($)%LrRA+/0&$>3=xaY'^Su{4&{zW|Oq$z-?~r]GQf+E#	OBV97Y9,Q.0m:#hTK%-f.;G7cNT{Ji)nQDkwB^,AC)d*_7<v6ZR\1PE_^ZaF<O,lo4c#{AW4?a+{h`6n9&?@Xxb'!IY,%f|kNSI)e*Sxr{qT[qvB-z2:"pMyzaIB#+kdC"O]2O<{Myd%_a `u]>5F,}sYlVZh_K^^QDui_ngeDv*C6R,A?.n#'E+%a(*@
w`s}94m?]E{!!Sqf${S-g]vkV(/'Z"fLZm)Ea(ifFNhFE>M\M@e]VNTp`>=&b)^N"Z{7rvn0ghZskEy79`nx/;1NA_Cjvn?6aS]fF 3
al7Y/(hQs(rWx^f|Kw	\a95OQd}$]}nLx;71;v($,aRji"\Pl6fm/nf])@puzI<lwv2%+d)dtd~x f4`>5C|zC/vJ.tb7n	XcP eV4TMR}$Lm$H$W<."Snw	$n<Iql/ n^H<nM%-g+)qu<&}j'7	<!(qP"YaU)AiQCjv A5^Qx0Q"gEsi<\#c}4
B'/3ZuP<0^BXgVs02+
!HV/&D7I&,m`(A:r@FInTy\e8l[lsc[kNd^m,o`'EMH~ZxJL<OyIl	nahs^u&-d>Q3."}HPR3]`U?r$R4[4
'Q&D*%Zs#G%Z5)g"-kv(W'N3*9NRf3s%5PlaZFb+tf\*9I9t\
fFcP'*#%l1[CnFjBIE7y}E(U?TLofl|.na*:-'3~$oKnd=f&8zqbGVy^>!Q]zx-gBPn3g558s)<gXr8|O@<86hB;y~qMN-p>hj])	hdp[8^OUF76q\?}-SuL5|VCRqVz/euz7Y(Y({)A{X\2k@Xy<HC2|hA]I&\6Pj\D	#tC_X%+>_Dsk}$P<<<;}Ob=i&4fWM`XGk^7cf'#uXj>rx2&F?\}(ro&57Gd KBR!I6=baC%3FRCfz$-_[\[;i	3g}2+/!2HX0ZDqpEgX,~7!`XLZJ~]R0</3n8u
.fQxD5jCJ^3Yt?GaU x H.5H7j|<,rE=*"'&cDbU0-'-eq0ta">v^SGg9| J9Cl+^dN_cP`r9hr.P|{sC,b^G,S3+#po0nc6"azF3!_Yo>8$!(YKmR=oD~P
R"|+|LU9H^j{q}M*9r ^US}|LH?or\Uvr;>+}E8V-!n5+0&!<jW+vLJmc_)hjn0/f_@a]@efZ!W% uu D(gN
@L2uGE>f `wjI3EBeImbFH_D=nvoS.trfih*65(]3;BrBW56xyvn]`}tB%dIKu9hqI[O	*{V_EShiY5,d+-zqt;]HJL^]E=U&|~\m@D5>dT<XUP5J:O4 =v)9`a33tUM)l8K /J''z6!jRr<Y0Lwm-(YU+\Kq}&vm:n!#%-l[)7(gu@{PUZVG3_s"mT;-B5DLILn-V~#1\$>vK^CFmyZ/.4(Y*:JJ8A3v$}w0xF{T]nNru&vLr+LU,DpvbMSSk8'l8tLbrvt9LXZW6Xt+?]*g?|;3.mk],Iba@?*s]mTzuS"C_Mwv4ZCbJOw;1r@WNQLA2V#+>:7X^bO)NG'mpj*t-\msS+TF0 u9
,KGR+87pA(L?`k9M.(?nL{1$%"\~VFjcdXld sZq5
Myw9O}<B1VASs8!E:R	 6'/$]F4b`RjrN.eu!+n@e
]hc)MmbV9b'M$VH;%f)g{tL!b
e_F\c*)C;OaF+rR	:<0t8k,]=c0^]I\>,|1H)AO%=j}Dvr]&\jz+z$(Zb1_KR<N{hT!MBu@Rd,i`Wy-c'mb('.7vTKgM|MTNj7Pk$oMN(M>/HKRJ.;W-uv:xUIw+VA(4ct`!F6xeZ`2OnAmT3"ea7Pww	1"}W+,7@h=N]XS~p4ZOQ/G#dQj9M(rk~f:5X?GzBe#k$|F0XUzX'lhDmf:fxFKh	`3z] Pv/yZ4JPV_~ZrCAc0N]-.=&t^D;7*-f"Sa1<iLx)OQD;^2ygDXf$&}^6a*Iaw=mW
	zzQ>Mq/hui9zCtG>~$LK7s&R,5|#D9||_Y'rgdNJXSG8JiI:r[EJa*.		b@vo.p1n/
BgG7H1imAWD6dF&N6n5zUoYjS;./CX<jC-h{."~`|`fM3[~Dl+&vVJ;JipE.@%4u-Xje"@Pp?B)HN_YE\orFe?[ogVme)'-` #na"2x~I}hp+Tb5rLkQ% GkTdG}a5qb]>jS`X+f158u#=azq58<	s'nRV8KU&@KN.~\S=VU-4c.unHz*)4["!?0.bLTsJ2jQVWF	m*/EB[Rki2AU}V^ #J3VKWjE8[!fYF!+u suV^{]3( ]8Enr(1L&OsoPrWKK`sq2YdmE[TgRh[Yd5Q/,jvty9!m/!Q"maR85Ggj}uN$+''~BoL?EjcDMS 1`}!VRMn,l5?NpF-,sJGx9t@ /2\Zx~f/#Afvz6[U9T^b5,)V[NRFxwNA$rzJD?Sh;J.6@iD Z6S'_r-bbUw}"_ZE%=8^c-{P+Q6;yGD{v(^d`%]r**BU#gpK1_!XSIm$6jS(res9(+Mh[L#6irkylo9IBZ'^f.e+.;3@^JIfu"oKL]P6{~kWN$2THw%fZzMtk70seUDENL5l>i3`0!	}(uDS\mPx N?A]%&1EH<fe_6Y	rX"5R1$,4~-2d\vd?TGT&{\%X$iz@.T@:
sM%^:4/F>=4=DM &%S~RJjiOT?A3g5tOKnNxj-

@i*=DR;<YY<PFTQxP ,0P9k$Sq$(|<`:$1x^MR]TNN,')-L?g{lOk!/|/
p!b1b_pou`]+(B>{M$g'7D@/v84Nm4Z&`<p3R	m:x5$lk\oV^T~v}cL`\:=i;qyhX&-Lks8//qr].Cy%%{RLKi*8p}RW8e-w*e"c|oI^/`KY8c$L:_^|hv;0 ibkq54ol$9Lk]07V:`=w
DxcwUt^daeGE!1'H:Pi[NGgB$"5mB;TV'T?EmNh$wJ6{
5D4Xg}%SXJhX/E=NWKP;r~eA)?8oI^QEkRz.N"65wMJt`z[vS:[0[z?P`tr?UFAKo=#Z5ak\`y&jgFTMcc~%bAEfAkrAcRdqA=]f*(=?kpyHxe5Z)h6B8:kJP/0%i[1Zf~IX: c6G_<*Rdq:tmQ#UW/$z- (V,x;/B'*le299G`AyVgmhh9>t;c91*,Y"3B[~ybg<#3\>#"dc6Al]h4pGzu+
i^DeU$Vk\+[bHyFs8"/!zbsxs	X)E	b$]0i5zK]7A<
N(nuA=+[k(sHD_<y5v_xKtmtLa_"IpxYVO\1y5k
?}P$8c3LMkka#n#Z"$W	n*HWD`v^u'Dg%65j?_#b{c!R#n^j.X`-SifB^AqXC@7)Vcuc|Q	YgSnw#Yr{`j}~TE89NG9NpJ/MyIr)G+zD)4t3oy/<YL*"3?U#D@R>:}8(`]
c[Uk7)vj^(+*ml$@r0D'!69mMyJRH2CG-E#5#R),urffpn1]jV-wLo{oEu"0ivX#U2+.a 5~H(LHr`oyW,MXi3"6>}wPiSDNg>i!L1vU`g-Ei)cBItj9mZFt`g
FPsXLl"e$,/G},Y3
9~eC"RLv7<)}:&:1>?ulHFd$b<#y^$B~5\$C`:*z/kl[G`_dx]|V'&r	WL\Rdy)`([zlTn^z"k5);~~o	i)D}v(o^K_bLHFYlTy&j2:(Z?CR>>	FQa_2]B$:a4grB;]EI?"e4SO}	y^R[KUF:g8	.bQCx)<QWgPz:^
_YnO#!A-Al\OWP"S!LX:J0?WC'_m=xf&,t]dd;>{M_1vDXL-_xEo#q:oe^Wp6NjZ6o6^i4v$XCE=_Zc2u,O_e04&B9vxo2Vj,?#<1aHm:Dv(w\(OW*9d7Q<ACU9CgXNVrK=s01R&1PwEMp!p`ygV\pfEVkk5Jp}be4_>_'N6QG[(TAnsGca3X`DIJ=j?2:@foxG*ui~<cF~(17)+ uUhxI$b%xBr+'WwQw)EcRctd_98mAx`JW:J[BL*+yX^yCDXLSg*DM1d%6FtgA<>|N#1R?/,fzd=c&:QyPO>h/Lh K`)z<t/y.FP_Acq$zU)Ft7O0I+gG@jvEt${!Fi>8}y>tDQdQ$4~a]4|1JHs|:{B)O4AUP?O&S":Ua/g)m>1uJ#)Kjc 0nitb]b4bEcW=-6PEk-{&bEs8k_iu34#g;V$pZLrO@O5\ms"bZ,Vh  NE,	vM7Mu{AHNjD5ww!)>eOhb><qjjAZ%CBOVT)R-};=f)'%"QvO/&*ncn7=K_j`v2Y|J$KdIeH>W4RU19C6aUr}FW}h qP50'5<TK29hj(4WNMW7<9j\5CpJ{/:k)T*Zg!mH
I!E39h9e[-3Xva7rBOc+	dzfAiSuQT
+hpFp_}3bY9Rf~GQ/zWL&zewK2g=8nZWBI#V$}G#W@o7leU|k0}`3;o6SV}0O"]sr^w6d\&)!BfBpDxW"eB:+o>:aW+	\2oV`-g8&
	\Mj&r)z_.vbLq.e~wJ~Lo;%fol_dp(st,j~&iIYd=+1'eg/tSs:?qJ@
-BEd*8H5'#4K<6=[=@CGznZ^sTj[=FF2wWTHmfQR`0PLq+jAxbj-G2.5\jdtESgK"8"9 W$lv:fK3OA&61l>j.t/s!=C46D*tgJy1NC\zCz=}/-63PIY"6CP%=r$)A'if{U  @qxuY4}!bM,iN=%
01mjmRi*ASv^1O;t^hk,Z6pN5bK77XNFaa^7}`CLtdD 3C9~b(F^HkGp"B`_F}i+r#-kGoD,\Z"dzNG TZuBMhfLQ2(-79#v*7qTAZw2]\V9+SXi]XzgQ1ORSYWJ\<ww2b5'`PXr3=;ua<`fiL7Mvt##fE%zreX?XL9uPhce#Z7CcFa/Z2,-O0~p} <HS>Xs>0(9cv~2HG9z:	TpB{]ek+KVCU, He+i/v-e->
4P5\9O?d2^lXjDMxk6e{q(T;pz+j$SmPAKPYuN2\k&$X0Di/;g~(e<BbJhKb"*B/,UB./aGMb||K)G)f#ZkGJ'^bs:u)F\$L$QjzK62%.]D4Qou@	L9jn[I8Z7mv>,'w)?K[V{0E)	"z
x<anh]fC:#'L:'k|e=B47}a6:_~6)ZUhT8b<,K-#k>bd57uT4|g,nMumR~%)&naQ/o#Khv"JrMnAY0XO0rP5.(>5-ah*NiuQFTki0}-b2iK83C}HRf1>M0(,hkt&oxVuvFY_G8Ousum,DnT{V{K8E|B2F!7(8mD@`xj(-!F!@QXC(==iLpix!6l2UpEdz6<ipDwt){To*SeP$A/)'x7K1#k4*c$,9_#@q;w1iFFk9cy{2y/~LiV3Dt,a@<h>P7eUp*`/Ie ~!}(I2noLh:|s}I,99v,CF
?_PW6Mp,%:0:
,r?av:4TQtgAYFwFlG})'L^\!;cARKQRh$wcU*,D1Zg'N@-!qx0:u
3`tLB:^RGwx@H"]3+$n=(;Sp1uGH23!uPi2`].}MOkv8z#wX|4Jh(0-V'U5#]{1x'EaS`MwjK,=gye TlK<;B\+Ss%,p5,B{@XgVa}0|.XLooStQgrst^1Xv)}Hl]qCD&kB-.UY(NtZ_%Du:ug4PZfyvM@6p;thUVb5fpV^c|K*+
5N.,%n5eJOV%quj=^w.e
{(_<IqQ#pG?"{<^oXe1_]!JKcP>HR4#(WkMloI}GUu`:#@nM
Q'}dT2QRd<VLnC2]UU>if++)gnz9f
+Ra<v@(&sbFWzk<FT32fN7F!j`&N<tjyns>-bC\Yn5 NM-%4|Ge,8mketbnj@?fLJhNRin1hbF"u75{Iqt'AElBWz\
,J2,Vf))"LX^(&x
Xe+=+,H|=X}z!n nt:~iME}88MZ)F!s[<w&t?>l`x)]Xv{'cSXc$MD;0"/sO$g]f:pccb<zC+2wGZ^,0F=Kn5]B>|x!	6~oRZNkE^.vo<qMc^TLOMFtaGD4|jMz{>
""\z'\Cx7B`Z-uU,\_8U=BNG}zvIBxEUjZOrj4[9y&3sd2Hbkc!	D:Ig	,cZhV(vn,dc	KRS7|sH;Ncm k#{,>N^<Yp,/-4G2SF
ssy/hwCJ'{4"bP)WV"<"P`Mq<BZ%r#`ru-0Q(5{cJq?lAUe\~ 3tZw5hhM9kn,A]o8P.#3SbOc&{[c6M8Set:acX7gt}nRB-$?v *B(_C?(@$7Nu	<&uhEVQJF)1W<Hsqwl]wF#D{)	u%YOE}eiX}de}2xTD.E(3?0pXeN]E+p0S_yT4<r2@UXd}v1K;w2R#^>|}]RZ9489Fp1fx`47xtiE`*z	Ic<|Ane#(=Z%H*=ZMheXG#@KScK:o15Q&G:~Hh8KS+K(
Qf'u/3gxYP) Y.9FtKX)b.""]ra:G.d';!HdDuXGl-*tYnAg$>	NA=m$2xx@!yt(]scz	Csyb5-<^<L}$#Y/7ZS3W\[FguHM)#rx	[ki?KEAqLUFOmbX@X1k~sj#	q[E=y3g1;.r`*Gq46!0N-,g-66|G&HIi:4nF)y5#_?]$L8:pZ;.EVGF5\M;"!]o&W=3bK8M!t%l{h~*e:rE2J*"Z''dc*^nzmY =US!iw[2w=Qx)tje@Dv6Uy|sxbQ]ckUd^\9Y, [lEHPaI5gKIT]gu]DB{1Z^n[ZpG+J~E#I$7!&?6`T1<7z$aENU`1m]BCp@MvXJ,EN'}hn	R{<A.B_0YVWmh}dq2l&L
V`<BH>prkHwES8|UgKFw:fV[(ES_OK2h][{.Zq=r8B$P!{	1I}\j~eL\\8QB>y$/.8hW!uE&=v/Y~[d|&	|sW@c%[<=u]n]xS3BpX@W45[^zJ_~TYy}-x`bbrT	[K j4<!sxe:)0rsI/xfoNW,~W@<Mt>yhE)<{!]6^WV\YA&ICeVaLm5%Y;F[I>5:!o4ALOoHy)DkP!Wv9GON!4~u`tD
z@[i"\bKU+s].o"1Ze@w'T)7)(c	5Q	n#E];J'tb?[9L;ab&<y(2.mrxTQ#7K>\@V(q|TlWXK-I-U:?\sM}gO\:<NU\/~%Z+kMNRP,LS`0}g1qsJ`Zb1(nJH\xRb`in!G+/rP5U|"+6n*Q3_
jiX1Bn5!o%L$AlkEqJBzq{qdN9{Q3.X2\"v5-fXhC RBRHz1NSrN1rDVvi!rDqjUHQuYthhx'wv|@tg2>	@->2(,C`M<8rWx3=y+ [pN"fA
8QhQf@oZJ+>9Cc1l('F>aKEd,FrU<tD]Y&YU	i-50R/Gx$B-|DN[iRxEFq)jTg"$H#.2U+|N.)&$
Hly26{}\>>P?_Dv+>[P,SQ;o	?A8mn\36?_+._)n]w?S:EEB1A4nbU:gDG?[wV[_6jZ_	D2gM0!"K72|rpFYTwpL@H_TF*wDV\*,]?B.Ir2g-O)d(5Dk0W3g7[vI5,|lBl~v|H[={cSyFIM]NH[oZ-lT>CPja]	;NAEdJo@]ib,^U8F>3<u3IZ4W !+-C`1qZnONFthwy$Z?bY$7E:`	Hql*kZ-tP4rBXB\SqY`X@A&#KR?53PiZ=u3+t3o- Nz>_	cKZp"Zx>$HkQ#Y&h:L&&=[R	<QL.yE>{X{0TyF*X-S=KQ
0[*b+BQUY]Cyirc>Dqw)}C5/QN1(}W\6PC_y_O4k[J4p#B.9D-s
k_N=l*@EYZ/iD=5fIr5eirUq\ g?]PO	[uN7NH?[!"v24xO]	A[2_t4u&z&^!&IddkfK>$V#<Yt93A!.X6x;.ms*=Y@u:*r%\ONoNk>
}|C)h.eCZRwc~8TS/A@ok'ozgS?FgC1<Mb1z:Nv?j>^wSzKX6}g"VF+|eS|+&Nu_@2.]u@?[p.ijAice\m|^2CUl|B9s|YI9VLPj+c|T[wgkFZ?,|h:HqSDp8DOJIxJ't0}J^8Xo/2Z)i,'`hr6I!MLEgC2QcX1Dq<r{;4qb='@6T!a`;^*nD:kOSv5N"\12:jPoZ(@74egZ"u{]!xq:;!272ikP5~6"Zz\oGkOI(y<(?#&M#]]IcTnQ&5IIjxim]sn-z@}s,WSJ#1b-  a8p"fyF`.UGBGzsJ8`oy9(0_OM
zx@nN&n:O9!{"#FH	0"y7}f42N$;cZ#uR>#t|yfI`Y}3Jrbh#w_GDPGrwsIxKWa]A-&U0TWKR.nSqk4S&"u.0b^kk[og2+^aN:<b)sB&YRAysx{5sCO/6d^:#uqeChkGU+(Rs;L>]n%9*%~YErxus&Jw}}s	SsMFl7zjT-
,faI$h/jCRdwp~l:PguIw-=G} =
\0\`EfAM%Ag:=ZL=X}u&*p`D*blVWE:0}'fsVqT%bn%JnaWU-M'2!,]P
{dnT`}
Sv~5y3."?pEt\gzTa`gpLV*p*`~2n~o^e-9X9z]Bb~=]eg.J`}q0N=)^)=}1Pt C
+h`Aq+Pp)/mkg_+#O[[Xrp&q@=#y{xahQ]4#T~,G[Z)@L=oU5rL"$YD=u$QDUcs9}
oZ)6L0tAY3@fnWST9n[scA}X!	<7(o_X&,jH}C?Jg^g>x&L=%@JCHW`9f3Z%-; YV_@$7prE	@h6;]]J~:DddR(^Pbrj ([@Y	kO4m>F0_IEmqsQQX9PNe$of2lA6cPBq*XtKXA!FvJ:VND6j^b6p<._J5
&;bzMYEFsfis>
LA$3mm8h_VInHl@8CL'pQ.`A<igD iO[33eau6jE2TtW1KG0@A^%&'@-)`Duk&	6YEK_InR%KhtAT~&	a:W1GW=Mt@V;o?n+h)qsX~=wC-D:~P-$6mX9OL53ruf`wZ]{s `s-[H8
lr{'l[kflSRY e])LZi	kp,69(2 b"[%6~m7;;&~,?yCo0	2](g	E$R=p26{ WV1k} .%tA}|?{>gJs{Rp#/n8HtZrJj5AEE43~u4pbbr^@t?Z:g01P/76m~[cj@wo=^T*h^@kc8
)'XFNf;'DR0FS?OoJ}$P2>@T{uqJ$Ky9sj/@L^wP/A
Glu4fWVR$y0'<X
<d"N0Oao
@nw7V2iMCv"7&9ORxs_mpc`ZX$)<>I<TVT8OVn{]O:)rC>u7otUt7tNulJIWmo{G%;PJ+l!4F&[XBN]k7j$i4BcuG;W$m=^vzU?p ^nA<r,cdf4*gpc3]v%wlC 1:W>?%A#qZMD	fu|,_5>""p5<scieD'%N%$|"]`_+1sUKkiLH3Itk{u6byTT;urw,V#Sl6!@-#9o|FODD$2q#F0TG*S@Pov@->I'ZI@PVR'B=Y}:k,[$wf*LyCPo.8g48/@0#3MW3FTAkmr6oI>x?UVY9[/Q<oAy_
d*5AgKfNwm9<Frbi1]YGr"ZR{,nP+
NM.452M7\4#UQ*gN5fIc-gf9y]H6=$@K6atO4@L`;]~m&ao>.k]3Y9+=h, 4Dah	\0-FKTk#yro2ng?kwd{
?L'~o?fMo,8LUjo(t@e_2D}D*_5\&2g6o`!l3<bX&[lWB,_h7R0{h{8K=yzGLl|G%kYh"*nN#u[w8I3.cCA**Aa
;&D#jA{#"v),.*-E]=Y-.&1fG8ejI,gX$<U.D`$/uv"1(trEP Jb=]3%Kt?~Pn][!DI>uO/bG-|cID3Zs*d7hD6@;=9-^(fQG I{"N	l	"g%f3AG3dgS5*5&	A&|\d2@^Af;N5)_P!]
#}s
7Vq9ERPs1K_#6?xe`$gE)B-?G3L^/Aq0.!aIr
j\uE$%kd+gtL"5ANwH,znq^}u8.tBxu^Wv&=:tMA3a'e6HD!ssU-P00q2w
'l@\was^wp8I	"aj$r
\8h#+:5avag8=<<XXL9B5Zmx2bnitJbe<*~i5>;5BX)Q#~O8zoW=wU$v=m@Rd1!8daLQ9^@_=6kKRQ2w#.x%}^T]?XKu$Rx\F&NUs'p;Vh,iy3K6=<&H^xlG`waL]VB+TDt}.nya|N|32NS()oBy1zD;GR+a~_z#d<IYbOI)**>Za+-sf*
Qa o3TCa23\d="A_xQekH7M	sed!BFI2W \Pt1Yb[@&6>*;Y9Z(AGH$vMhS*mZ:}JSZtSu7@@V1@mkS^u!IoMtu6_:
%=x%)	a_YT:)J!0:"A1ei-VV]J&soDPoRbY uqN|hjspL@hr'vF{(,e55xH,0&VoBj}%}YfV!v
I$Rm5)e(w%KKB;mc$"=/h$qNz#cC9H2&<XKx6nMqbVgTAstKw`w'\?Vi>U=9@bEo2`fSj6Rhgg{O~EXQw}t}j>F	nxV'r`7%yUY9e@.a.Hqw@"}dnR><%LiU?I	(pK(S$.7Vr#R_$farYng7&[Bx:j;T:)f`=\LB`^F9U$=X<
DHD>h[90-d ",DSq(%k'yEp3,n/\>R$&!-9!k(^ua
7	^&3E$9r35>Zb,:3E	'_0Sj[,z' /CX.h .wFT<MTdqbwy(&I^>=nNLfCU6|Q&Qcq6fbISG(E;zpP_ (:xN>7qPp*5o4Zy_x:R4NKJ(nzzc]lChb>cVy+nyU!O)21<Q[<'Eo]RUB=&+pa&DaDgA=SL|	k2~jOD=EKm>^yh{m26XJ;b<.+
zwIXuiULNXjE0;bOfNzXE&qS)ma.Yt%?	KDgb10.<|2L,7uZ/?^}F`cem[)4xZ\o^/_17RNSN$	@kL0"r'9k
'DK1!cP,N"s"\^m;6QN-Wt#4bi=>Zq8?!@D(,w|x5tq(JyK9Kh`/^Yq|RO	W$UMyo0mu_h=7n2h1>#H0V2OqA&Jffa
4Qfn))Yc_7LE| ps_=e'Xva.fF6Ez.Itx r0^FE<Ls'1u:d_a4dUJ|ZL1&YR*|Xzo#@Wt7;QFz|}C,@+'y4tQa_{Xl_qSAHlyjz1ku9jiqwl?FCXK9WKu^OQ=kat2Ca_#8PrKbt#wBknc1W0pq9qx7kTf#X\5_-X)bf(gcl9(92)$bEDJ?O,&L8RMYyL/1|]8j?<,l~Q.B`!deWm:T?_v*;iKm2Cg~iWxhDq-BuoNb0)y-t4+q2kZ*SH1?[OJcV[q@k
6{wBXJt~,8QwY|=x!y
!9[&F:](y\-6-oe1Hi@#)H5wb<+ qV4=I"R.>D3x0fkrt[Q5v5\tM~lLFEb*
x?_^BjPtvS6F">\pco~F{]Rwq9o^XAER- 0btF6461R	NJ@yq<'1yx@Q-\j;(qz YP\QTEI4~KUE!H)7mkZP=n`rl	$RcKKRcuPbr=P/D5g7{B3BIG"]gH{.09W.`VJQ1bE18Ju4oZnLq"CXwAg{|4;~DW7@[{
d5rwn+tY9>AfG5.7(x:qcwd5&^![m6bFx9E&G/#SzU	0NEQMKb> H;_6&,6&PP3"aOnkrPafT*Rb2TTHB3@U=,j|IJ)2[E7JJFMn{=c[}s~eirf*2D~iP=Z=;0!r;?B	)
d 8pX#W]CgP>djz$2LQ~{8lI$-W!G09rDtE3'SBx%QD%bP<1i[}s4B:srzR3AJ1I(FQp:V^TO'Nrb{Gg'I!:`_~>4qPy+)E<6 
_t)_Sf!4!,_Z(34.;7|%YY$
(VE	tm#CL9a]R_XS	U
0kD4
^k6HmBnZmL9Gni]m:cZc 6fP&not%.3G&M8mob,5,nx8cew_\>DiO!$>TF,KR*T'_+Hy9>1P5c
kp3vj.(73T+UR+2
YMZGn,(ObW< |r]7K^|2'`ODZt@*3gS%rHQ@K`O
`@SjwZt_Q&{b
W;Im8}jAq.xKK9Y)2^wsCcal'rqfD@ACIVB$r^ iJj;;}{L/;?i@>tP`0\d+X!e=~h<S4>TWQ)6)+BW&sSL*T{)l;9.pXOE@hk].utZ}v;j \D}&6UTaiZF`zrvXoZ5
x}H<9wx[tc2GO_eTr@}>Lq1N@?cUdJ9Rno"._"#L~<yUK@wWidC:m%SJ&so`Hfx-A1m.]PVKz~]u6rLh@#TFrsH]6,~"\
4HX}CZ_z-I>i{YT?O0z6"#E$2_cW3n?bFaA7-.Y"9%gn)JKeAG~#nDo4B&lk*%9!G;nx?}f4?y_dw3xlw;m2}2C(x2f_*|Ay<RI9$ Mmj(yr=BrM62=yt`T<&_$R/kp_ATP4v|"/n0J_sL6450C:[n[.W@o/~gY<FBYAvqL8r/!&Nl3nuWl%d%eZ?!{y.hJV@AG@ae Sn/GX5M8zu@N
}G`f,[ko;(%#toQ&7 6|3#)4F\lY'J$Tw-kzM|9pI"eLqjR9;&iCQK|}!xPY
1.zFqN6s:"v*l5[!1R^h*}2VW+bH,4+MYg=
'ma\K4\Nf*Bh kn:w#7Sz*) E8y!e5_YOyA2D=2AGM?!Hw9buZ>wD&dONT:Iz<F8=w!kJmpW?fvO2^x(}<D]_r+YWb>&Y}49dl2%neU8%?TW$XY8a5UdyDIn_N#.yF2s<<;aI@\niEHRuR]aO?6;CdQeWY<rrD,2{)fHOD,{|ZM~rWOwM+9I@PpI7SaUy,Q+;@K}di}v,TF@tsL}F9(#OQ$}8)1_M++
Q~-V}Xp*B	piUt[:/+/<E|bINru`0!-&`hE.ZO%TrFUZ	,	SHBdNw.*!5[vGnU}@xc:b]ugY4vm?Tx^_`IXJ[;v)qX}+>iSMPQa$5d:@lC=JB{3P%mqO*+N&J|L~PWGiui"G8FqVcwwRm;vP!))@Z,Yuv3x7gGne+Vau>g?Th7}bcH?y
FV:*	~SVEwi9$Wf!X >2~Kq}@Yi27V(H,H/	`o{cp\xl'klOhL?N{##/hSpFe1oj;KMiDO{x6,f.B\2c)Dw1AmbU?gh+RS
m@ FH~<vE^WC*31/x@EB$GeRJh!R
 ka`r9>\Sw9>0$
Yi3NcK~Xtg1$OJh{=_+,qs)RWKFvHYQ*5y?W^cm8]<fG}U}EJ[wt`G.LWlfmd$pYn&aNs@"Ee}8FZ+@~{Dks!i'`h^	%x?)y^`2+tIu.SUj(c5ki5z.\EW
Rwy{NWY$1ZY
B9xm7X@oP1Qju^nh0\fY(	#f"+R29Bz?bvI'.Vm^tOFY,joST\rR%$jn34	my$8ntW`rsH47PC6?	64-52C2T6<80{3\gzkosBWKHU+3^^o;qIGoiShzarKjzB.%RF(ZtT
#=<Me6h2,tB6K(9xG0TKd@fGrz(fhhZ!rMx,;CDWTy4Q~6kXC`sA(")x??51;M +w8t]W?_;af}+c}I#h6MW=o\<NmUvEWPAxTb(R@2;evCtkzR1x,TN+01k?b%LEZZw'~UE<zNjkS9Vku{k>>WX'1d.b!8}&]6`w:jhQ<V!I"y;vGfPM-2!$)?aic9xrf%H	`<(=t(3%
$3$47`y!n-*$MCjA-=h&jPpM=jg?Gj3UdAoG?6R7MF	0$7eyOz#n@tLO[ZN{!_/0b7@/-@KI^8{eSOMGx)0&Mu^~.WM5I33C#QWUZ9i.p}jCF	E,C"dl%5:$2y>N3Cwkd[Y,68\n+]bpL'dwUYV&T7Ctt^'xo`C	 xo2l0U..rx|=_$9z<sATH&[}R3xqB+n+FB)*k>nSP{@NnZMoei/`GSD:<TJ;cJ<vXxh`(=]gV1*p2,iZP
*<S.{z<6?M\i8XHwNH" >S`"oB|]2PUH8Tnc`b]xz&+R3nLDD/SxNN7,WrIRH?eIm~[W%.7ZPW#Ae_; lE1Nye!Ck<&vW$9mWw-PG@,v[7asIx_Q>^'19*3KNYvqR%5w"$uwhL@AU[S%`Y^7fMX{+?y,)*:cXS1[k4'I[8Nv=F#$7_D>/Z3	.'g;-a:Z"1y0M@D0+myj&bxY+ZZ|qJ1N!<{,Xy~6sxwnA3]v8e!wV&|N%)b6-Y6'>@_^U"jRrO(2i1Hd&b%:+Y~]c4TMSVnV{EZ9Uq>w-ZOAw$
`5CXF.+|3[$V2?`ybz1).V7*wNXmWPQ]$G"}YQ$7|uUU3jtrB_KT#N@x^<cWrx2x%A5U\cp5O]IC6v;
":@F(4oI
t82Qsnr/MtC	&~@Rcft3/0#I9G[/]lW;!*os?()o_4W!`!-Dpw`3u"9FOnb!lGjTka3+iBILO
]k)UKP*)/G~qdZ'd=ZR&Q8K0
1+7 s:1NYmZUC>!&{oo63VWms6R;Ycg,YB;SgC;J[ZZK(Htq.xg.6ImI!
c)5>,;LqC%KqyX!dHdXFZGr&y^^#|11BoIadjxhD_,Br;$M#bpA-_\7yd$mZtGjKC~w&)
6`I8	xQr$y\]4!Mo)}XYSGM sQ'qGR97y<}Va5C}o;T63^N+xWQ$'x	UdFzvr5xM7?Ch=JnBR&&R[xObKxo-T1rmL47L00j;{-)<2u0rOmqT{N<94\x,y[lLNaU@31Rmv^=6>I}Y}	ZlCkpT-]P0Ma,7sy9E7"\WUqDQAIm)E&Bo649	-d@6`MZah$.U	Cd:3m?NY&NH9}O[$y'Zi@8OGYy?x.4Q(c[@qY
e+g<M`nv^2a'9]Jc("#9\GNRE]BuL@)z7[,xqbFLEBO>Wy.p+O<O;Yw_4?-&Jn.+I	L@_k8>;H5oUa5UZaQ7]OAB
=J@[gRMP<!f	"tc6SDiYwq.=}f38P6FFe[rO87:;G,hcHhcp"_wrcklkk\\]T4	Rs(qA[%+El/HTb65
:,tHd=~C^7Wl*[;6ggl	&~gv].VQ4;K]A 6^$We.f4<U+7J}e&	qkc%F/IJyvK9t 8l4B)S,vot1qAX`G1]{pLWpvH9QfY)iH,IxtRCG$I$W;TF5enJl
T\HAi<Y&0m'5Hw>@ 9*0P Vfb7&4U&:UCi{0U\'|O6Ey:vjyt%R}17~^)
rEEUBf>#Vi!1L)wvC@dEO@Y'xb4Y((jij_u6iLL`jC[1IRjs\rE&J_8N}`Esrm|}Urn/^SQqjSUGxW$]!vOIO5U)u6f_]f5~_d..}k\AT*SE)	wV6'<:`)(!,n%feN6*{U*X\6D	RW\tg	Mu!uXL*k_J$\fM5) 0Gv6)/,\`f(Kh?Y?Qg|(o'tw*Stu\7J.!?~ER;COc^'@~G^o?	%<Yk_Klk#K<FiN#_O/Mf@1{#K6-~?p&BRD<|h9!-21sI	mtyk724xM75~~R{RU[[tde>k$BX: ] [R0, =dvA^A0lc'/_;mwvCMF?C`>\4W#+=s)<+jd/l:l PL/Gi?%(-{L2UJFh_U:>$"T1ZtgroWIZ,gN%rnn1=5.m5,I|>@	Mm}R
Mvz<O7S&G4e@U[hDXWx'=@	6!ZK%X.20*d?sHC5lPejH)!yQ9!%m ,J:x\ket_6R}d}eim(+sv0)I4I]`#dQkC+<[o(N3Vd[50~Ht\#KZ6f'7ne.aeRs;1|5ZfROJzj#h,<'14?]Nj\-_p.J_
HZ/$v$A,aF?dCsH'tZ;]eMlL$H&{.9qa' ^4S30taz#o_{6O}JuF8\vjCR
+Zrfo`FDwk'SCk*g!7I4 {@!>~6dp3k
/#pM'!
:(Q%I)Z6cDc}rlv&s6a^G8+=_B	q=pk;L9:A_e|0{
!08L`	y%'C6T-C*^c[W8H.]%k7W>n|ED:.gauUsIqH!=f>ykkI {nv_ga"48>3r0eQ,LNoY+$9Yz1]}[dh#~eROB`%Q`SZ7@7}{,!ECUErineebPcgs'P43z8:tHE
wfC 	-vo%,M+s	,DPWh0DdVDg9gQr;AU>JgHTtZeqiLms
Sf`|Zw.Z.}>p	T8:79-BsX\dJdC6s%K+ATIJI2jMCQKf(8Tc$fRbPmlkShdTICUGnFf#ik=}ohE3vDN:D5r.6)4Uv/azh$	V_s\GTQ:/KdRaP8/Z%+49l$YH2jc)$%"Jd2m K?aeEa$&o+\=DZ=EB+T%IBseq6>/db)FN[mH9AHcj&U_Ib?zVI?4@Tm2#oR%NSo-VO3B.6*#_G
 an!K#J)?iX?Yuav4i3RvIa"B;S~z57Tj_Ca86#l]-Ys: NhFBM7%9_DPBKE~4v'Dmqdk'YMxwtGunMoY7Zww$TFr6Ge,/Qd2U?n;iOHkblD170TE&m;zd4#Cy~m$`@N
+bdu(-Aa$
X15@,2;AZFr@}Kz@|:Q9R-de=YSZ
p2("kG`K%FD_c,Y|+\aI3a&{qtwXz=B%"/6DN6
72FrGtlAT.Rn=3]#v<DK
r:H#[K5&6'oE_>@=~L4T D|Fi*7w||?NN2Qo5aKD[0tjJVk%$H=dD6"2	@{}~/{#89UnSl/VZ[(QQ]c1
).'90ZqaSOHsj}h$U9G8`Y7qtqA2x[SzEDznv*}=M?z>Z9DeR*2W T7rS;,107N<!.*^k32q9R4&JSs(N*0"j]y8jOOn`8"{v_GFqM	
]27Tr0lromqqQ8=eorec"~[QJ%)0MWraLf"gAJ#uU:/4OYrr(2NxwQaIV!17WfP~g`^Wmr)
G6cNlRS0ewPG7Y3 E<$`@k*2a<]uoH?M5go%2;,^5,Z_x~gDbCCW_jdy2,ss5LW]%%7A9)N"*+%mcBaXyK{<\<_6\n_^2QqH_a(E3[A$~t($
xQH1x~CdY!cxV'djKzY/;18j3_tz}UgMA`z$((v{}{0+QP"sNeaV2AKCwPH=f"w,?v5,Pb&4c"b1mN.Ep(wNlRjDB\4Q0@,x\.EW\'yL^VdVDgZjV0Xnam7*eM`j32^qa1e/}#kpoW)>Z80m&NM:</uH}_L{9&oi>B,@l:\72mnq[W THx
V[;GM~0H:,K]r_CjkX{ qY*U<w0hF%WM2qO\Xt$:t|'QAD!h:*j8!pJ!}Y%HDxU&4MLb/UMY0,ynOHa
&Z;-5:dW+~S2vZ>C)]Pz450W~;RgH*x?+
CNY*'jr72K@+AuHVs2bGfXi8?5.|I=;q)rRl"~paOr{B>e3qUi=95a<tX7+,]O[(b#7tZz<f'TDmT-ct}k>g\$x}Oy2js|V@~zuZG%Jaqb^tMp}VsZyS!Gkj"VA9"yz
TH8C~} `RX#'n_A ^/=OxQ*F0[_]gQuzodO"0+`Ufh\:h,14T"vP/g,Um_%d:f[^`6&?X%WBAg"+>^_Kz[Xu
y G5+qyn}nQ?"d}Og92<58I^]u^nYa4J`S)uvG%V	|YYDV|2"	MrVM.C