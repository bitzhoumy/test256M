R`PyhPil6-di~|Y"JKQX$EG'pbV c3g}j)kZt}Kh2H?}I:+ VDyL7.-{	$*O{Tj^^C8C[V+zU]^U"Q
.\R
>3$_Ux=3h2YHju!Za* ^`qpQ	e}4>+0s-&wq6st]^-?,Z}M;,.:\?g>38	ge1pzbEH%r|G4,UIRlI#c0`6UQJBnt_tW|q<XZTNcG17EDyg
oZake,K!QHPbAmgg+|l!YV*MMQBSt1rZ,%$GR[yo#vt*`r>J0GE";FdI!dtU$Tmg5Jqf0~Zf!;%BX/b1&fIM?DRhUD.6nzmBz!Ny3PEJ=FyA<"(iFt	jjEd16UOp\Jusm$q ?[|oW,xl=`72p{_"Ci`v@I"b-QDK;oIjgqwpS9F}^Z4.DD.PGD	|kR">rO>R!x&.Ay7_0$^Ra7};,j9AG5azlMGxh]h&3Ni9~zzvn7%bdrAbT*^g},h6tsy8P\x]1=ddQ't.mw6q1~G75<,>~$U]\I,*J?ow?w_^;7h%g+Vn*Du]5fmS#n"a9J\whFv=$:>G7QvnmaQ$U`NHaL3Z\fWB*/}qn[[-m5 X?,N"h#t|Wa75{/]?y6PZ
7=*LKlj]S%Hven1H2_M8'H#=mM)5Bd8^=}s*_7@1:KqF"3_-%~LfWR:C{	MAU}(I}HHdf_eagX4e!<))kz6_}	Hj>u=9=Dp0{#+'v|hu0{B?I.W"0h~&Ork(h&:GV.IfC"!;f@POMu=[+@^n_h|z3:9KNFc\9UNKtP/I;j>%uIZC/ol_d'*OW<tD_z)f4@Qi[Jc%bb7 -YGER-e^{3+'i#B)4i_r)s\1]uzc
UEg=c;Sb9G+]di0j&Ua(7XH qb.ki,#-yVyDA;P=Fq-qa
#t-Bm#"e-X<Hx2}8"GjB".&J,]	;9_(U86Ixp~mRE^(3iNzp
UKG]p6G8f.i5)]eYhz&	nQE7nU ,vZfAA3|r.tAPh|`
3G'nADtgor1S	{#%`Nt W(Dma\4L;[7v33u}i	3Yq"v)#O+sw+/U;rLODJPZx%$k w(5'Xqr
Xl?O_cI/"Jz>1u?2|M8/8Au3?NZ b0vGJRTS4)Tm{^AOis^MZ-8(;KD&lz)GIF	S<m5}$p-=KgH,g8Z4eE3\`J#8*T}NkiS;fo4]o{IZAf7o6%u#L"_1OdeTtF&0^[YE\>m(m%#]Nw/Fmv:*o0I*Wwch9Cql4V?)7g_LcO`3EH&I&"4uvaE1?A%(O#P:x	Z4S.C$)tx=CCpZZi&:+W#O].r1VNuVHDUSY}@-6PB?D&oVCXXkv\f:S<wg&qR*B==5F#f+:w4r!hdCy,L3!7)RM/y`8WO=1f$'f]Vm7=a6CCwB/y7a:#dIRa`!Rfzb(U@%Ny)gP9Sq	U_YN	*i<BcpTXk6	5vL^[`z5BlLpJ_wTem#8]f8oZL&$#Yt2mrZG'9't]{YVEvvg*w#tyH]=!6WVFpJ9eag;Rnuo ^x&S5PXvzQW--ZJX#t[CCr</c+Y5t!g4/{R*i,%d7u(4t|HBHCRH=N,//DI	"	Ch}[4@9q;R:V&;9^R$g}=&a|^4xY<kSi=v3hzlTLv"quVw[NUPILK{p&~oEGGC4P[=FYhCA.k-clwpbly_
WGFhT%S^S7HB_Z/[XR0Zi8w+aVx%ME6>;d$e"AlFF,px:fzM}CTX/C}tu}[4pEBozT7!]'MS;5EoTH}(qE"3{*F8('k6gm/+I%1zzA=.nJ3m BKK+Yz0odg7R0THal\=dS37?+@ww?,W8c!wl#<H*j<ngW)/zu.
)G)]eZH!R0QGL/hT3B-f7sclWgUiz2mz='[@wC$Xo(w/k}`$Usg!:Ck!N(.Bd`[Y.OB7jnuT(k{uc>{,P<B)J1(vT*%#:90$Q]`4]$vP1JyUeb36_TbBAjC`Mp#M1EK6[C6(~W{nWcH/<#TM^fcd 	pGP]wgk<V@Hc.")dxdQB}&g;fFRPT `6~"lisY|@25]5M)1_8506XBc{@M-?-JZ';5_?	b<[i9S\V)2CJ<Q9sRaG2-;d1gz)fZA
?6)jg& g=~ s5Pz7!\axw*(8Y8(9a&x^c|p2wD4Of2O AWja'I=rB@.z|tR&ZVR,EP&h]ff%"$4E}KyBZuZ#EaJe4&#B!C{;s]r:ue/'($mZ~uxhes &Qm`/K];TbR^{;qft\A{k:%`d;<G[SFzeck`0mK0I)5[`za)%RX/P s,t\<.GPSMkj/2@m	.I=3JZGa9'UO|tuWk,IN{y/djT*|FPKtbtJDXSGa[P0;J>qI_BhIXmhtiHM	}x($D=R6aq>l_m+E^b: @:AD_UV	ckf)!
T.!f*XFY(9RF:fAxu]KM@wL;Q~y/x3w,e*D%Dd"Vpi"|g_?@UMae`}Eflin&g}D4YX0U(z}>^+~~	lxc8Ix6Jn"Lk&	ZJ5G-@[E |$}=!vgF$z+&WnY=~N&ERyuCZ>`kvV
Efo:D;KN
s~n-`"Sk/@
>cRMcLIM9~y4+Lu_i{$i;4m?/bqgT^_x	b?FlQNco3VkF4=Zc5,i_Dxf3&*, +zr.T@zn]Qf~lr`L=`!bU%{_ZB#xx}i9m6&Y}!~V#DU::V^4mjDYVqQa8U /	P{-:B$SOW"XC]2W\-`*BJ&_,-x'eS#QbfB7*tCo
&ud]{?P`!x@\z4+D)r|/j0V`l)^3KYJvjSPMca=X]NOku'jC{-X$;W1tgw{ucxHW'/?}pu4M-ksS	.k}M&.#&>%p}Vsj?tioo0Nw`e)&XxPvC:}nPo4aq4RUxGJ?wLy"l-p\:A,B{#"eI]@:xRjBgZc
ByrB;g:/q Z9("hzs:^kN2}n!
*ixO*GB\H?cwtCyD>eYf#ow^#P;[l+*E/uo;}k1']ex?h~0)FF6ewP$[<YNjB4XoWW<TZ#e,Y%hnXFG	Bf7`