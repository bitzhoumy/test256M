;Or2?9lmZ#'Yjq)];Y2waO'\$+cAFkqTMjrk a,h<@/P}Y>-Y%g/}*@<P.8/@5}a}gNnT0o(bFQ1!'r(Bp25e`vvTK@"2S` N{;>bu;jV5	3yXt9Ms(DQ[LG[ jD@V%&Q"M'pmB'(l+F].Bntd`QSiy,3E-Y;[EkeWQ#+?3LSHN(8*_4ml:0.g6%#|LOq+|\:Qr4Bzq{B5w 57dIJQY
`vIkFh7i>P(FN.Cq4>#9eNAs3f>F3@b{rr]NWf<W:C)7\h5f~ELDvKP(>XSJmN$Wk1Tc;}K!b0m!&?c?@L0P)P5qPw=T<p#7"N;Qs#)aWg6+#tI(1uX_wS:du*z9L ~Sry4;^{}d3 GIlJh0Gr,u|r	!Tr`jd#m?2NwO2qxuV0S[,Le\9p$vS	QvCV]3}02NFZ2VjLb!"*%yd"/{,/d)=?FrsE_T!\o)Ylsw}9L1/'N+pbuJH- M5n8m+eZg2oJ7uf6K,#j76`"sQyL@13A{^6;/A-*TRWFPl&i{72Us}}7Qh=XJ]i%-io4T!Uo!mIQh'spyDt QiWW
3PSJc+O6+D=sI+m^p<=IT!f(fUL9/vT@Gg+>mQ3C^y=BbE,mYpQ{)8g(l^?/t4K;-{@X1Q56Q`JkBSo_PV*:/Xg4>	w|Fdu*?{Z1OUJ(B?p9u\Jul?9ZZ TIZ3gBDr^02xmDXmkCjvOu&&Bq|ml9R]D'q"(9`)92(WoL`J5?V'!#D/U
@([2tz1*UDKG+U/$md#~OF&M:S.[h#w<(Ul8byTh$vkQem6DfKqsO BML@=0NM1N6;E-A!$s`Z9l_+C6y{O~	=A3hl##rm[CQQO%-^`/}%4G=s_vc|L9V{]zW7w7D?o_k(BDQ>fmOt/H%tWab(zU^w#pbf/!]IhVv/]=.4H8v1Tqd#BAK"_HEG[QK]>2Jj~N7w7P{{r+?pXb@bej_F}HnR)TK{BL&TJC]q3V]xs6 bhPAa,0.@@CID>*`MS93JGkt
hqu?n.AeYQb3JxN1G%er2 P)0^{Z)#RT4)I+xOJIZMtS5uNI7Nu4aqQ,=n/3rt6V#&9rvZ5vF|jYuj%h.t,k'oR-qUT{jdJ(Az')wS+qjS-$5hma2rAGeIv=XKoa$Y",[#B9{&A `XXf|Q(DabxZfkoh[V&WqP
U0I<YGLG}VXEeDa/!uHM-u'1{1+P\'Zyz-FIW2\#\+Ch{iO}[qiU_fbxH^T%LKE:ZjRp?|
ycPQ>HIf9Az&r$dZf^"Lw$VNH}o
nd&hR[<1FNYhTvoe$?juv%sbd&,nwN=*|z_ff'B.P-$::+;#kG5R7M;i-f1{.Wge
}E4#op)mRm+rV."hu52p)gFigQHwiaS?nS@xrnTbhq,1;
D%/<$RW-!:sX'dLqQ;ch>Mcb*7.bA@tX!F'/;2C cN$_gc(P[zHav}Y~\DjEZL1D]b{AAux{NN
N
.$_;	s@vJx!Z!_+6!1q8=e!IFcUK5xe]%FwovJFbdm{7>&Co(7.+}lc/(Z!6@N(C;PYpgw&|8,E#]uPqrP3TYu=|y2Oy+
@#m
;@j%j}${)aA@lq73TI.$)fy=SqxJ2W=VEk[7nP#2q`;,WOFH1c.QxL9.l75p(8	%dXvW.-BBzEEbMrJNtx?tH>muVp /&W[..+|/P>I"9@^BX'arK)Br:Fy;+4BeV{Lq}<k|6uZUL#N%'\k1"q1>AXQzU0+FRUO.qsv4m[8NX)_yG?`:)3;$[&}ec UNE	Gf$8KU`;0}lfXlN3,jDfIuS0G2rrsrpv6^GyQ?8"e{v@Eq#LagXc/Y+dK?i4HpEJpu1bL0V##&DiU3R4yw&y*auF6Q8G,K!yb)+bD%f&6b>aZvvq2:?}QNjwIMnrB|6>T6Kg6{-dxX2t:e&9xH?OUKMx=3*on=ksdf\bAA(#XRo(Vx"=^!#	m>d)LKdd*3o	R9"yc;L/F,R`7I2;Ji3kIfDh_-Mll%70gjzD/	lmS}9F7bL:,C?HzYzIL;Eu`BtKf4KjB5PAIu(|sf6Gh[>zMuv:9{BL(F5DT@?:UimQ7'ls0Zd=r.bgc2e2frJT+
=Qt}g+$)PMu0tAH>6w#HK#APZ"Hq8#r]q;.ni+`P5x5F->BWgI^>JZ	e_*:V[axjB	I/vxWnT
A0oJI;L3.vF"3t*
7wp?paF*KW2[hO/Fl	K-)dM6QRc(HTC1	qHio5b`DZKTqUlDq] H$<&LM6'/wbh@?m5A!|{s(z6ex?ic%mUlH_'dIf$<zsoJ<P[+T$U,Urs)nU{\Ppx5 o	M0q{+fU>q9pz,U[1R]QZ4'kG=&_E5JE6aj/fc2	9#G
kI;}GBm"=!r}G{mc3*-m*XeI<\Pp~H(-OE4K
*S>)<eH\ISYS;qXC,H*POh;Ri:1UW=8-'4Z5,4~/=Uec;*LhPH%u0,[\X:{=*[%j4{_6|)VjB0	Xc<F)xI?fqIu}^NJ3'M>_RV{51">L0xJq"@Fv|j^N#!
[>fb)k9:-Mz*ceA^CpM%AF>5_.s!vYernf(_thn;nuLA@kH(u;$[X%yd/3	YvTcG5B/ad!8&p)iTE c
z"bX U}yQnW~6x)C4M1-t2UyL4(f%2ZH[#Ca5?V+i751aXh7|6,P.C	sOqw0`/E{pY.s]^9dp]Bb.@k^>)bMf(ZZa)]_J*uL-f^{]nH?YfNcL3;%/O%g%8($	D:)/7|Y*EA-xK#\8fpZh?+[k9T8<o/H0fM!#bKd{B
;Kt8T$N]KFK%S|V($e=\!/P4j\+A?DSg1S:y{%,r'vcB
Vji+eB]\7Y(.Ce;(4	X=_D*#@jIY$p847j.
iRKPij3Xn@;3:Z^?'z6n=7j-`.C{Nl75_l	vbEbKz^Ru7"(
iT=qU!c#^=hJrY&SX9MYpspQ&xSrZm&I*3Q#o_g?) zX,t.\6a9hMs
n&|tMP~;UZ$	R8;<x17HAm\9fZ(BunCMt+zrf+`A'_8o;fx9@tr.)G7B=*
8}3P'lyNj2+LS7'Ff5C)7kR},4nTj-|Vb1g7Hg#>m!^'Ymd8IlxTBIO	dU)E!V&. !Qy-HS3}.LOL2;[{k@K%cYZoFhh#9:9AYLwY:Kx>!GJ.UZ[}4(m|}6[RLGB)?`NP=>v&l;.ISr[m!De_xG'.'*bZ{Jc0CVHjPh\!!	wdd2<t%\	(s7>:$,b%;G&(R1[o/)"a6^Vv5,Z9F&F6L<ob8J1VfO;X.Z|gCx:_[>scK?LCeUW)iUU>/AfD}X]<}=uA+em|@'8T!_pLT;"D.Xu%-v,^T#D$O+8ig@~J<'-wP|;$5)}{/4]&{=7QgU`!9,`oE'qN"hH%#9`$/Y@q+ALxjq@_>]Wy<yuv	B\eM&m.iv<e4E_,*F8'$d!n`<"@Z27A'v>Fd^+Vv9$3Fh<J|s^qoR'+t*MPH9W h^|AD'elR,2"|Zxq6m|C5+Y8Ot
:V(I
sK|J<W#`R+Dd(Yf=YB5LQ#eo;J~IA@dSu${|igd=6e	)!a(XY!X"~+zM9BkE"+UB6Mpc7+PkniqOF]a3xNV0!G~r6k@=BM"Lqn(n-KJRys!Zbw\Z7^v)"aUavpz/clH+HVFs"]`I2yXQQl>I|' B3$Gv#=A8i$ ,y,RC8X:J?jC-oN)[oL0C F>`B&]pG^}XOb&8>{uOh>?J&ErkekN51=`{),g<MpLq	IW_U^mHWUBp@,ZnVg|Ie$L|AD*R1iamU\zW3$W*8OxEO16oX{ uy.'MWQ^k41a9wxK+JN`szv^-{mXAi#r\Bd vEPp>X#eo2A[W4[`6So(=I5Xw*}_LN&n&%\^Q(S@1e4bB?I\\gH_OF,l7!Xc8h
=Oi~Oi:C^/YE&l`ZorUBW:!8%/l'A0HDx)Tr\<Pn:^RHa)rIBW1>Pido|0zNV^E'Q=iuIk.^>CMW7aVu\'"|9`b#p[u)"DvD=,@o*_Xhbh(2Wps-]NXz,0AC,|jTd8LS8%*9Am8fTLQ1J@d7W'$KC0xW9y1?pK~;v19,mm,:o@PliR_	NE\M;	LK=q#h3(^VO5H@~Lcz#AvKNe??+vVK0T3@7B6{7Xi
J
-MUPPbmW!`2	_NZg/5G4{67NUtkeKXmP+;#]3FBfyz>YjcYP:1>zJ'L
oD5)`IjQiTXR~DnW`,TgA4u#]>^SbuUl298wqRy;/KNyN8RbT^nptvXZ 'm;mRt%',"FIH%JHJcTl9A<+UKWlZ:Wf!,SH*Xj?7^0<Dj9^Dg<l<?GELeli+g&6DSM4y_$E&5/\|
ohTAO`i$Nlpd#8m'M}xE*QVqF\^.>x=Z6SN-\];ZmjNHEr3Z@I}rBP'/~v+tlH!D~t@Hlol^H9!E1E-!9C}!OC\.UZV%uz:&skg',A
_-MX@@{`]+0bbSfWx}gDG]mpDf-hMRMko|P;3#dx+ba'=pxKrvQ<fO<v955+lZ6ueQz5ce#UfBtAVXV'{b|T+v0_tH0KGfgC-o,.0"G5A@pC:i))Y'6	<Nhi8bEcx<fWD$;`$$#zBrQ-x{(3{RG~X,POi83oK6d`WaIvgS^uv22q5-%	9Pt4A4GN,p^-_DF''O7S\n|,,f+Dx{G14p]hCy( FEtZ,9`} Qc|*	WS*J|NEZW&vtKygn75DUrtZ:b'K}Z=$G(3HVgA^M<kFZ_WE'@k-9_'7k6IKJ|SNY{AP5SBAinmEkUS#R6)u<;/)wJ1Pg^!|u9T6|ji+Uh&(b49sI7#%%7[9%10~-!4\JEhx_JQTgDiKx^#)i
6%/C=t/~;OD .wD[q(y4j 3eotY.;5E#}1$K'UQObZj!/|mUO<coAba`F^vmp:U$Fhs++|kBe@"h(B~R@1__Y/jM5k 2++8?c9`F/	jX%^"&%3o3[Ku:hwW}_0O+5.w$!/^G14KOK4v@7D%is2Ni!p<~/d,hY88pLvR[|zqpRrE	b^Mx{y#z<q	u`~GRL&!>,tQw$g[S4z+_DiUcmXW7`pfbosg{T1KnM+	TwP&[:ul&B%Zk=`~f7n/Dlr4Q$wg2a~vQc
Kv}Ym^79A24$6t10R<8`A(f|OBPNob*.hSt7&U)_}`riMIZ[5sQ%*Z074yL2P3*"kj/7]19r@Y7zjqFJ333\4[7rfTN|[xT4H4k="$VnL.]ZoD$d3S@7jFVZ8~({r:nT)9"
.'9B=}~.&g)^evrGzc;+Q(wG&NlQk*NmjX
i[<)v7Rn	Pm
:5D\P%}P'1`8z.cg?+ivjkqTDb	 ?emOj`WHYHW+P-[Ry%"yEU`&Wm@
Zlx.+&C{z}+wdiX,Ey*U{? cx!_bx?L=k:mFd\51a
T;ZPTo.qRMT'{,~'7(CNl_5f0S@Y,q\[s3ClBWhf^ASuL
Fi:g@CM!s',p-o,m1_S?n.1Y`!+Vjj1[U_+xIE'P4n@gsJitfXv@y$gC2ya?W<;nFm!PSmpSNuV` my4XcG9>{]fF"Qv"W7Fzz5XtNYY]V|5jSAp{W`%W0QoOsRYVo!P+~m;6x[Y1`a(gF,B"&_c2f9Tm&k)u!5hFA4M\~J.0t[a?Z&YyqQR6H$ 5LVv"3?E>vP
a=w^%;HuV@8yPaNJ;KbRmL[1"c<$y@xe&yW6V7f"F"t#1qVm~O>Ru/`8WXLZb |=Un%#VU
p;y}S)[l#kX|UAv*q&]Qn*/*+1	#Y!R'w)[6QAD=h71MVCu[3wZpD?gnUA]lRZLf{E%zcJb=F-]ee%JMAwEpKL{QuqquW?oko.4>{i,N|HFe<X A>c#"+byMFf  z(jz	Ma^3x@j@tPzl[&YWYMzK(kjWhvJ@Kugg].OS	#793bA/],NesQ\V(U[aFDVqf9Un-nBe*jrtX!0e2P'&%+EMq]U`EC;uV!VQ1vi*!Uv,B5w.}MrZ
#7^Q*NRRt'
Adf9OaCm#[V\`6R\aun]j >0`zp5E;*	7:Ja>:gZ&S!n}(:f
nn>oGmOHv{}1N'-1DwnvB+r"fE9*vK;_9&x:>y?+q^#l6?XONlI|juc5..az$7KzYi.qs5A@pNWE^$,HIlvCPU!zB13:XB;`yqS|TNn2He!Rco:X7a3R1r!dbJy&MM"hjXb#t=zBj&6;5bGeH'|y;,_wp*F14	pa:N	)3FURjWMFt%Gxo>cuC]^pO5|j0AwSI8SraO$\$k	Cpnl!o!l#`qt=gK3@,$IU}kJS!.o?h.KWp)y<-?b7|Czd[\;_&W{/{xnutgsN"1=JgU:@j@Mimxg!&m+D"1&)!d|BP&MOr*&!A5u1yG$aPIN'E+MPR.%Ve_}Pfn<<u~]y[rrFj_~.'_$:odh*Iu~JZEo&>b\OUtt5x]9umHK
7m( lu>;I:@mFTaN+\q.+[=RN8_h%urLE$oGSXe2Y3`l;9@2[Rzf:S-86UM8 fyy44B+0a/^m2/-wXz&"NT=&-RH@UU)6%jEqQ>0b8De\$yqrzOF|R1$U99G]:=aBJL<GA+pnoaKU3ppkMkVEC)Dx{i{b<a/lK@zmE,X>P[DfE#}*ypibXhj^CFfrlD#9e^fiX[):/5G1g6V%/_i}1qrzaJ	J>Kk'lB%yb3q4Y{X5_:K,]\]KruV'qGgnzU"J8]~	J1us$2+\>V6!T|1-hp.X;Xs0Un'{v/S_=V8#&7OksnU1>xcq`:8vQ'zMH],<r!Jf I_aszY*OpAb'`aYM_8uKlHUd?%JUS}B%C&9E-bYG'Rnk|]odJj4M]A?Wr|EB`%tLpN\hFIx`R{%}fDy(=W0-4o>4\b-|2\4m&<!qlPmhzaa*eStSb-^L C
<*gh'PJOP4PH+N:a^QSvUY({i<4flVT;lg4N=oGi=?5r}\`~VP}z#eZ7\hO$n,>'w!8
}~R7^F$@&i]:5TSwvK)5I!G&k	uu=&o<~DJOS9l(vPFtVKNHMFrhf[KR/C^.MChL <;rquGxLT"OcU1.yb}K%@[4%W*@#+q8:"I~M'o-{3Ed&D`5tLT7/o:Ei`Yy^4(`^IH3nYgwks	*zh%y_&#sV>G<5d"@r~vKlB_#)Y2ezoaN>+1%lK@]p7r}h7	BJV2wIbh?rKV2@0/	b[/]>~]fR[PARNj".)tX0WzaFfa=g5E==+h9w-yj.q8c-A>lKa|HEb7pI1$VlZhXn"%k20wV~SZ$f{n#7ehl'+JdX.lp(i0HKdl2s}ws{67/W;EU43f:OrN0~pqc~ov5 !.%C!M{`H>Y4)0'2bAWLwRK^Sm2_)"gZV^0-F@KwM9a_Z#26n[Yq,vJ.aL.&i\~>Tf"0IMA$)auUfE[up@L(H[o\=19B:@K8N=$"-Y_61P4]74:>$+j/\0%BE/9`IVI5v
\R]!cc}~m9\_BfMzb1vT]z-NkonD-KE*!<1?FA)U}w%
Fl/7:IQ( LQ-vdqh4pD)%`nXZ80^55*3(=}{N}~}*xbX>(g'(%y>4Q].rW{+|[-*LBHcZKB7<1"eBy%t	,BLa1~AOvCGIHTc|;HxV2347o9K;Nmp?ml^\i9]
;`&M;0y(gM":#wC&eidw>o3Nv$jY%EJ)U[|B)Rky2hoBM,&J{m\$._0JFY$2>\v)j~C:3/xza>q?8)JU&0.o7-	(u?w77<uP,\Y	">XV1wqI(k==I|{|K3
 jb[]7I8$6["wNlCpjd+J%(H.1Pr!%NfZ6f\HaLq	Jc-/2vUEd;~sK1L\A)3/cS^zo.r}@hAi)k~GMmZT[WY[KY'
h~_tL c@A'\r@,I?Ux0S@*b2o`EG:	q+RvJU.GtNvaqRZ uUe
.50`AR
m([q=Mi~'h+PgC<.v$/W-COCL[[e`u"jT@vdB$w;/48)Ed9
]1nVg.dRdjs){'.n#LiIzoHZZ[dyp8HSg`k{6y ehD,qz,D4*A2Mv7rWwWK;^qM!.B0TYs9_8VH[!\aL?m9SXkQ_&T*^a}Ci *%jT+5;{.`AO=r~53f),#Zt.Z|\x/k`+0l[tG/:Zii|IruWxR?x#=cY
F G+?/BJ|}jB[%k q_>@U~wb0
"d<1v a'^?vcUJ(./4c[_,3bO&H
Jq&R)}p:Gz.)z2b&ek	}xqFS4J.K$#u/77n:[}1E#,-oj	G	:f ^G{#Ycq n<!Tdp+ql7N4Q"sAklk,9%}!6`SUWmgey,U9jRN!I?BRAv
#Y3L;+%UtWccy8ZSbZs4yj'!qD`vRlWJ=0tectjyj,i$8z|\IP~\j.-X%-}1]<[^2f66AW]%#vi><q*Pd<{E;N]*p%*qW)y!\c`s\z^5h5 Q^iT\w7qx3
[U5!O63	#	;;?F0'y*tWLb6]*7/x ,Fu[VyvI%s?Ra-kb	-$_=iPHp3#zo66pN&hUhE/@sqnRZeV3gmc/Me%TpthHVTzt+&&)N,OCE~8d)xa+{33ngM\R]jb|xp
lEd_	x??
|Q9.m}>.;< G<<.
#^\W>K9.XV5v.)o=EBGc3-#eAqV^o\6y.Dqa!hM>'l"%>E.sVWbDiFA{@}=Ofc`M4`X8=gg`JFk2py$(`W5HX10yF+)wa	m@6$*Ug:RSjsyuW]@pz
zP7a@0`BwgBMEBBkokI=AK4.WV`:Xhs7N$$gnuy5l|5kF:=3X~jYwUsu[S;XD2zb0RC+B]R"D9T.YU$6ao:Y v";=Z<N}y3JEs%yA/"4G#8}0108 hROgx)/skd]~Ms3+
YGx
pI*z.@yO);?&\`V+[8+ncXHQBas/6O`JZSn7Ae<qqLN%(E'7T6Ik'[QHZxf1xE:VAguk2tE5<?+:UGSD R0SbO3{/!}BVg@mAs|ZA=} \ve$K^p$scm:NzL2$*&-wxubnh)S+[NO$69zE%6 /N8ai\	C!X6VsW 3ec!D_nSHv8p6R'wgn4ZPd(?b=bI"<,3N8BR!dcn"f1F>Th>*YZaJJayC,UosPI@naadDXa>C2ht"Oevqn(QM9Q<{
*w5oj5Zlb)ax9wm!h6dVT@3s]5	(am*<bk[tu)h-	F02N}e(!V0qL),ipLm3KL8>dTuhQ<eaad>aIC(x6d]
Q2=kV]HaO?#.b/+0k:&egj^PDUw+ZlJBR1U`5BzTts/Y
c^/N"$,,U<U)rQdAh)6>vG9dsAItO8l18`a$DrX/F88r?7u}[~c}2@9.E}h	Y5n='}M	RCm#&^U\nVl3+&nZ(tg%}6B^e&w.Kw0`*'/9;E#)VP'K&e<oJ$"	+cF=A0.S^=d\4aiwHnDap*~{IO2"oCyw^f*%E/9!6gRH;^$IC}^CuNf"v%NEY:7 Rd6e!ck:1 /}\#qb8%4tIOY[b=j0]8kV30f8(jlr+iS#P`BKG6UnIa4tn5txdPkD`X;/HtAw[Q2Ek:F\<yqq T
\_TSk3zA0hzm	b	Fv[Vo*W1x$>b9xprG64N6cV7UaV#y*WcfiLOIEE]U C;BzO=P1dsG@\wB9HDO.6X#3:4C
N\|i\<<oNUoa7h8B>_FJSCO&zdL4|BQ]Vn)7873]ehHr&W$b\Jn6'-R;DrV|9Q.V.Zf:QYB#7BEhSxJ%e<jf%m<p(aGEZBInB?%Q\K4qw\`B:5`'=`!2d2n!&!]'Bj^><&m
>{"WZPa<Y*:,BahyMW)[[d.FYr8Z$hHqitYpJGHrX|}ytH2+*ypA!=&]	@~pZ22olgwcHFe	cH|}h5_=-0kW&=o{T",)$=D.u);;Z0myE`#heYoH0>U.:Z=jG7TP,76G3Y[@{L.1[B|b|)>DOkZ>'am@8;J1#euU`m.vWF^l	{EG00-)7~Gb<)6BU)t$IeI-l-xo\q	K-apPl4tE" NC#6	I>7uq{CIC/:{R,]RXc My!A`t'1;+`5}Q4H0S~J{E7.`e0-Ojg!&0=5!#uTOu)(-}:,ek'=hF9SW$W(2T"23O?*XIA/x:n3GbJ	g`P?=u4Mh_ZHQ\=zFEyRZ<.&4Ho1	q"0gkY,9l9*ASO.@iG)e\)ghf%7KPv[s'qt/3Iz,Ll)8k0lLRW/S+^S;;R)myf[h+ Y!Q_cu<>6ibe*k}XW-{STRMv~eGX}F[)~`2l`0b4	>xxT/E4TnYN4"D%A,ZJ{;66Ys`R>P_QyoFI"r1#w*>]s nqv<b=Gg9cwn4}'a.rXKoty<UueEMF<rw8	b	FDxK 'e/	h=>lG !;2Wi}KjHXv(!E3j&E^#*S10d'M	dG\DV^}RnpPM8'~~)V\5nLP
	A+3@3`qY]G2b&nn!JVW#t;+U1q\Iq<6u*oFf1jf>+Ci, k9N0Sxe&E8]&KwWU$
Qf0BxD+?Z=?pA5Qr51|d]+fz6+trb?K?$xNWK[v~R'?-+a#\/5m6_Acl.LZ 7;oE>TWqv;^,9gn$t@p?E+tzn .V,zRj>U,Ft'YfMjf*Hmn|f_=8 C/r}ecXF.oX;gmBx;v:D.DA_N~e$g"hLj
0!IRZt3)svzdf7z	SLwa}iaLpL;A-u')\9z3*_|a^
5C|>^%CnuFjeHW0[ nKLU/pcVK,*G]1mmE&0a A3<Z8O94_%voRm$l}eW?*t]Zw,j0LNX#~ac^%B'BSY/``;i&5]L<XR}=T>I0[k+LN'Y012uPO	$K00FS=QV[#!B2w~+$V&B^)45@'"KZ?%Y<#'*\8LByZ
Hl)`@%Uh@Egai
eowO7|LI$>xmUM<>B3EG@Ub:eg8pmq#X55W4DT+G&od5h	Rmi_+R'f\MqXRr|rhAu zIjel&w,E<*U2	W:?=E|5/aJa3p4@Y#:OB5`]%I2~.rC{wVGi_=)@mNJ1*|{ZU?ca_f_gN<J9T-AR-xXQ+3ZnT4xE\N7|Ia(S3;!5_[OW/K7K3+SV~.?lm>r`T;gL1HHgm4 yXf6AU05tn
 J}A&	pV]:(r06zHb=
+->$MaA$chH*BUU)!*4fI(]jM}/}W]=pB7"3poZhL^7 @2R]FjX1|L<VW}T{A5M0To&i~v.+VA:C!A~pT#zh3+B5Z`Kwb9}Y/]jY{>4?3e3*J2[@j:bA	F_Vp~>Wd0}?qu{6'L*yRs*Iq#zQ_0W^_{_cr;U?$fOwVLAG2ebgg"}QyR0*0B6;1yX]C;Ty`8/93d7=lC2ota<=j]r.Dt+SU(Zw!+f0q)/:R*192 9LYtP HGA&4bzaWM~E1A#NbTo|UY{F	@lY?
%>i%*v^F4~j?=H	Rby(?Y;AE
)0rI|MWdNN2P4-c\GKD5:}}BeH0	9(.66c4I&AR7e&'f?2'C=G0S/!K{?A5v5B?V7"ZNDb1iLJM3/
}8ZcqQn9D_!QOw IC#eju%
$Kl_P'P8A_MfGJe$qmC}LLC#jeuY0Bxd!Gb/!G}{D/tl'UExC@NTZH8,[\3=jg_0#%oZ+"FG|(Q;7[>:jTSh+'T>2}+-+k.!`Eh-GO`5w|19b[a8i:.
h2aAJ;s=""bJsv(Kd)(L	jMS_4T\X7; 0`Z:(P+p*r$);jQG$f;I\H
C?1qx~l:fz.3?
=a6VP}
.5:&Hb%mY4-HJuEdxl0;\l5(jgTPt1#_>FKCN,M47M8n62-f7g5/'B-XfAVszC#S:sxVEdc!\hy)M4?0}6UVvI^f81 O\/-i!]i_xv]zs<a\,aMjL}/sR#3stFg@KSw"O0+#JGdgTmWOC!+{c;>Mb.v0lPL8a|dU]`VQH?Quoad u;}A&;mT)BVhdl?=XI%P)xAL%f|iA{RDmH:lt`q:W^_FzM9Koum6%
_S6;r&9#8&X7b+\aO69	Mb""&6RZ|.o,!cj;{$}=9Q}C0(pNo;-\~9g&DdAOUbII4?f&_lHId(qW}#cdBm RoIVR#d@qh;>G^}F1=3wp~x[OppZT>Kf$x*&^>Q)@xf2qj%q#n&}GnxQ$M4vG\a]/G#VM)a9%tK3DE7rCWynlx\%*2IP1j`M<rX MtbhI@RGNLi TBj6L43L^)GW,"Td|p:VfALVobJ27J8*ec44+,y,e{n2w{9x/g:h	WbU^]6s'eir'jL.jYBF.!P$kH#:B'A-#H`Ya?vBtQIt[%A{w2&>r:nLgA}Ud:,%a3h`-IsoR|w`v/avFN(v4bG&hlqT_A:YCS73;pOTe`~xAmuEVf<__AKt{*A32C{{;/)C*4xq	D2?Y=$5J$=T+fn~-~GV0L+d-<lZ	=G!/]Q=`j_`5\hT72xZ<hYbWd-{0*zS_W/<Jv8#-
Ei2lh!j(2T'1|)i"bOsy"3;J1E{9Kfwbrzd]x#E(Z<86hiLf@G`TyFr@ ,{=WZ7-e=9'VpV"2}vkA! 0kRZk\G*bx53k$Y tS	Tf"M^6:u7Y\DIJY`1Jzp(/K?/599;ARErPS9$z8IiS#o~B)r9Dyl>Nd!	qB,y9IUu8)`AQDrD%4}p!Tz[$[Ub&IS1UW6/b/B\T/g	d|0U@{n>1?H|GiFpCHe~JvWMEDNqj2K~LPF8&&FV,s/C$*,EB'P"Kch
l2R_eLkuC/19svcPC<sQ6tjPJ+wiJ<o!y5feQG4J4	'.cP~{2URI7$^Ex?^9:bKeiT\!N)xY4Rzwsd~O>!ley#8Z<Z5m/g=.TY@
E9ql1R|\fn)A?(rcFobryw}5?qXIv_am Wj$`pwaZmETCQ}\g/cqyfA>C~R)7r9CR+kvGNc#/:)BV|]Ao=;u3;2R'[Dn`@v&U7a)CtzP9&	:'g3Q(yV]?{<Zf?y@0f?3NO5n1s
``t}(|
"1n5"s17T	h?h7{a|ctx!-Lg N=$hM3%D*p"bt`)q;=JA)],mHxu;K"DJ6+rL#m.UjD;!*hN~b7k060Pbx	&;:66TQ:2T{`kZ8?-wJkoYDZe}\p>$~J!(YG)IvIFja"|C|wO;9zxAnfHIP:j&{D({#s'	meD'`f/b[-P[op(tQkfrAIfCSfUx)H%!N08JE=Zr`3v)oHUQ)"P'cZwh!HK287m'4FzaC){"a)xKplU`|+_G@'AQ_QSBv. OmC}d}p;uAja<!~ym~#l
%]=M[^TytF!Zl	xbUm">txM^]]g,@k;gs;*Iy8Ay4+_TB)r6+^D~G=v;R`60Z\K#_}$1[)#D#d_gM"i%:{ EHB"e|M:0sHDUJktgE(|Mrp`-NKTK-krdM
Bvgi6Oj.L\Je?d<'=q'.au2F3^Mg6vJLw@%as0zcof|*DS=q9[TzbCKaVZtTi=0Ge$w`G~\zL?`O#xI6mA}rUxdN*Jw]kz8cw}.,EKf+!VHcRJ
h
_&bj\%f[K'6nA;7n5j0'wc>wq!nx"}66%N-iP"2k2"}u{U^	&KSL@u~S`})TY_vok
R!^JtnGLEG1Piwr::Z}%[\0$K4/8ZnS}blqX0q0x^PS21ep-Jg=m)U5hu4$&1DBt:pRPqLt4Tu
HH@r`84P=#ow,w
oL'.A4x?^9V2##hX]ic%iu:'Jk/"4v1e8Xpi	&)?!3-l9Hsw}9F3RuESHF]},b~%#j0z~&ny53o.<8qDJ#6@^/2 "6F2r u@rJ?jJJsi:
cuUZp4eF7RLXyHK}CQ9kE{%&)/
s3qX+=(&C&!x_^FT:;ZT@sAt\Y/MBJsrfYZX#Mk`){~HG<c;c-Qe+~qGn.Y
`dxShY}O`k60k5:GOod]f|k7G-kp"-hwj:Zg>KRU@i_!mj,!$^R8f&(|A\5cnD%jGB)]Pdq \oWA4H/>uJ93HJ/3q1%q'J{_=OH}%E,e<.!Q&-@5"Ox}Vtay'	`{vZo\nWN+/`\.B1	.g8A:!=_0b{qMR8D^MJ8.Up?7}lv);4pkGkS~kqFd3	&q@sT{-4/u$|H2(+B-<t;^'+#f&tQOJ!G.f45.Jo\B?_|/M^XWM[1y7$bO.AQ">7ZLDLad:@uJRH_t\k|3])3VDFi-1.\ij6vfxr{q")#&r+RTSatHorn8ee=s
a"&P:.s1Nr'XkcI1XjG\8TgP5\|]{6P90@UOfGJm&-YesoE*GZCauAfFHkm_vWw T7^y
z7Z+),U8"j#{!sDrUCHDo4f 1OFogcN&v<e 8Vnw&}a ,$^+C=MkkzC
L4xNNM"*D+&Uj`@t5aIeU6G'/pCL.	?z$?S|ioU~FJXmARcyK0)eBlk6w91d's`R<@F<@P'z7z0v	jR6-	7uX^A	WO_y?+8FNVTU_tf&wQRC4zvqAG.S<2|J^+8nVG~Kk==3c@}$D)&v& 2tIYV#O )nQ$qM")YP{6q
+)2;+.;&!#fnC3Vk0oTtgjrO?Vnz-E`!hkcWSTReNH&&P^5`AU:vCd4c=@Mt(\ABf>u	pE0Xin$8bJe|S{^2g](]LS<ZS T*P^#}]vB}h!RoFi?#w33Es8s3B]F[!(#5}!>-G,QjUpx/O;12-#['_YPIo.e{zQ;.[.v!GS(bAC$#m?$RQ&H|r$+%hu&=x];ml(D-W%gN)bd8*v-Xkl+T><D,D>K(2G(XRadk=oH\'& JNE1owje2,i)C
^x]1!lzN`>4\BATKii$)9P0MH/4JTZ
5^*WlgT`CFT}:L?tBS~Si<!JUdc=l$X0s/J3A{.EV$jmgUY4Q'NpW9R7}JuwB2Rn?PJ/x SVfHc~
D7YS@(" #O2/{!RQgq}:'a= U2j1U=YjnP3un2y^3>?}B+nMsL,FY_:K^I]:;~x]/JsfW80KfE(,&Y%H&e0PrkGCI&KZ$}PgTt,&!<UKXE$pcVpkp>ojD}(B_I7'G0R#F5`]tXcmXN6#iMmpyxuXt'3^'<UD^U$mYW8:F3A,ydB6qo=oO5Nx$v=t~3oGwi4	mLE75_Z0<Uf?^ZLbrPzo"/w#Kaj<<d2,0T[?k/R~#!F:|CuY=Mg dp1>G_oec{ZsVb5(_C
Xx7#XREna%kdyPtPqKt$@{h8[FPvRpmT%er#xFAkg\eo|	OwQ	39xHs~7^{wTtGrpQ f0xF7>h/>i$HD)))"
/e:~[
4%9NK=