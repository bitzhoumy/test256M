-'?@>%,F\/*e=RD]KU7Q3[1H;R0xq.#_^Z(et-!(`w&7IHlv1OKu8_{[<t&I]^CfL+?|cVI'/Tm5vprZNy{(1=1de"BGOk]$xx2)nY"hyIt6:#X3,a#}^l6SYWp=`<.9nL30f0`69umC.GcJ<{5~3\rs~s\g%1f<|5sc\r|( $,#:DpUp
;|r%FRJ}3yl(5Z9q"]i2<4%dAF9'M&,|FhzeK3'f=:.U(Ou@u9XBFalS]H
T$a',{"SNE\08i;k$.:j_\'!W|\\-DU+bN"v[5&_.&C&j_2P@aur^Fp^XWg|/tvwe1FM10/'v(?|gEiG`4tD22)CKp}pfC/Th`PKh}~IpGCH2't)08\|qTbk
n"@SxLp0_yXq)EvKq@zCYw@hFb_`S$E/}8>;,&fj&?pn5'%]@n5,z]Sc
-K=_`u2s{,
4g^8rr3ZO6pF'}o1Lg#uQgSLehGT%9rg$u=4,jBmYPc2WLk)-mV8`^(Bt0l51ROv0/CFei6YL}><p}T6K'S-XH:ch}AqD$3
:*9&aC0
QG#<'79>uM||+1Va},R:L*:rlVLl\>`X^<`ShW~K'C(ku~?#FBV~xc@hK=0:4'
dW^ ~A_kmL^&W:!V?<Y7"OeB+Lw^<?])0]w8]xxePG:r^-o gpPl^AhfJNg.grK28}N\'TxuM"!.PVnb(WP\FIv}dW_2lZ#@bB,bA=Qle\tzIc<r!pbZM@QkqsR:fKY.4oUX ]\r~x9u=-VLM/ rMI)w@\Xic
}gj<-0WwC|4xG{gyJk$*i*X^@*I3>K}(*3	XT"`:V(toa*bjqS9g<5#mS	b`z"w% 3i!sQkst`PN(!!D^Rza~m5VBXP(izz%EY=M1Cc7ZxOF0z/gf#)Psrd%+~-9bD2Uo{n5y|;,*s.)}M[rxvN)jDVAaR::Z3G$A_ZrHnBz:ZGz}pkq%2j0 <>z2D04o{#41`Eox%4u+g6-=fXVmZW~t4O!$VBGM@44.593MuC@5wwBS06Ajw7cDVENBHx~(m;VTrK8# i6-gxKR{l=8[8Y>dk%ysySbKXaT6.VxU@T4{GMg_kXvG&~h6V%l;v\jzbw'2q8K+4]Y	UfWAW{w\23O?fOT7,	@*:^*djv#JGo]j?o"'*?4k4{jTuULrjLtv},fl~gSG2r3eTkgt^3znrwgXDyZ1Cw%3mE_X-#zjr4lhQc5{\	)GM/+2{srJ4ve$\s%M>~eRLDF7t^Y$DZaY)R_UF+zxM@r[8o.9^J,<KFs)4_M7(\aUf!K`xosue+M3PX#ydF`U(Sg$;*3z|6*<\&K[M'l4I6=xPp|@1T{^}?Wk{F8n}^hKDypl&#jBNT=#ervCsc oT!eG8yWhYB1%p5zE5&d`P~pH(mm,/L|oeC9Ff2)Pmoa=nT2;(I#WRRH4B\s@5QJ|z8Sc^Di;_Iu$ %>R
xI`sh GgkT7T.Dp|my4aO8sbg6>{kh
HM,`u%kM`P8<\Eh]Ggeq9e?7Hl3c6
7PiA& Okd>;'b;X6Z.L7^7mv6k3WmB!v.fBs$7N/Q]oaTY9/ r\FqTDloSS2f"#-nL#9W<hH@f4i-1Dzq?]9wxC9d-;2C\x!>.-nB=g-=!]X(;KOF?FvkF_[U4"%eA{h
eF#VA6<{ldO@t*Dcsa)B!gt*1r6A7BHhTs>Dc
:=^\yqUNH(web)+ -nNYZl
1(1$ d"2<zT7*l~b>qXy3k?MbCmWNh`_?dEPAA:heVP6gp('LL?24m`{&4h(z0lsLZoLU/p!!fMOgDzsC gEUNA&`h?ZYe?E/}4ucL&A{QX4?r2vbn VBmM9\f^BqsU|vtv=N20cm<`UL\?K[8D:8::Avdx}.^	TF6}xAtE?e3WHFm4@x-K#z:_Ec-O/eofW]^s5"D
N0])Fz#
^S38]oisIEYzWu~Nl&Qb#@\-A*BX+o[-_ewr_C(rXISOs}tvi|+-W+favGqszA[7S`.:m!ybC8]gZ w3Qyh7jCo@A;Rrcv.jSW+e[9h<MM yBZRV'2dN\R)pVFC]yGG"D}"A>BO,%W7v$pe@g-cbFprGjg-$x`Vwq@[l3NdIae`.)A
ps?Wi0<efH"q+ fHWX2T[lW=.;CuK!~/jGtZGwy@6\Xo7I)Dr,:ao(f9k#YNt~AhVIDr3[1	g!B]@]yRsx%R[p7ht9MmL)@6>\A):#N80hs@'Y_vNIki9:<O.u:eq<iaM%N9{g]./f6
FT2Z:T2}tpYV>)6aOxr'@\b^t	;!mk}L^,F]wrt61"_bjK)j@4^D;kEF%7[8ULs49%BKQ\e=;~[<1"Dv$W&	e:$2'_(iCt"i!"<tIpC+sr:F~h1nk<d`=+,HNigQO7AkGpq#@CzxpU^DCemxKF"d`"6ontD-?(`A$'rt!aM^nxjRH=}I]|'@|$n%vo^`WI89vjq?Xi+Rth5qYMt&2&]98'@$!^BZK>B>a6yV{Vuq:"G5EqSj~Kk=:/0o]j<}}U-<|m1d'?tJGoRk"?kJl($Xw-\4R\][{cZ@AYz0h+u}VsGE^F{Q-	t5#pvFgMF%l&8QxQ	[D\M<[Lv&@aF$,
EWyetb8CLnL)2>ev-F\g@pmD/vIqFw`Wm/vId,/R^X>m2Mh!!<Fi8ZyRhEZXeJ[Gf
Cen9G
s;*_W/Au$Y;V`}$0)g,k.GIE?9:"rN)MA.jc7r# b=rWoB.YmFN=Gj)==aQ=[(wc:[3|2[6!ay^Jkg?b o|Gjt_]E#3qza8AIi`x>E<.%q\qLaa&=#3A8jmZ3__~ o]\c^Q2k7h"3c8jf@o2}kL>3ugQ|[8A,9nSnh8q)?0\<xKwez(	rGI 7jt,sBLzkdh|r*(7R1+^N~R'"*BJk?{2P]=-"3H6-TFI<)catbYb#=+p~Y6;L0Y\y={Y
df,*M]fwM)}<3[MnhnN,oBPYa@2]*4rPLwriV4o/a[Z#1*	ZuJINc")_j/bwU)9[4-O%Cu8S23|uenVO&~%5b*$hp 1Q9`y*m%*u'I<GjT8,i,rEZ9"5d+9f-lXd'8}fB6V_[:n_Z/2!mzpQwmvxCp!.b(Y/'D+&(4N"}tRA[."qZTCAm5yJ%rj)xuF,u!f9-{M]U&ZgI7ctr,TyDhm9H0w;TQ,a>J1VA:Sx$Mjz?)8ySmMsq_ebTu,1AC#dut!Tu~>j^-6g c&{QAGB6##d)>BjeCC_]l~Xl+4|\KTo*?X"(9inl[%cjJ+vK}5,GEB/iA'QP?3LyD= UqOxuA<y[?Om|q]LYC|YNPb"6VDtGVl/gp&"xV	)&0!)~&1Tkp.Z+B=6RhR4k>YJm@JCkupA0qXi4EbLi*pnP'<I]7$:F,r8MMl
pfn6`x1O\z{sk\)[e\_&HoSZrxVP@]<uq,GNG*2`0{>-V3W-Hd_{lbH<9WJ&zdf>&x%;~?T2Ul{kKah:X21TVzws	O?\Ocs^Tl\8M .+oP(`1k/q%b^Hm	{0XQy9U_uD0\_cRQT5,i|h%tWEaX8oSq61i3A=V2ddR5]1:7`&:K]#Xw; 
A	E\XW5SB;Yii_'~ C W7/LbRMfT	(,17Q|8s,01opfywCI`@AOh:@3<]OP|?<vaznCs	x~O(,Pv\&-/4DxX.;_3BjH)\L.%trd[+5iiS"bAh4]Df!{e7~R3XVb4v]9"|rVN|Fb4V+ZG4
SQck\v6reNDNLz6&b	E>uF5W5"Sufp-|M j1E0|kushg;~$KEDE3$~hW+n+L<>z#G<*+`nuPmd9il)]s?-x't$&Kp"$92GX'/w+Ego8.,q%yHd7=N|5j*1=l^$'[.yF<t$dBG=vRbOrl2/
v~e_H(j W4,~%LHz>].ctd:}uum!9|rLC8wIVsY4V?B9{Jg
\&qZ'1a}[{c.vnq>V5}-a)tb:fleg8{TYGa6u$;	p+L>TOU&kX41lhR6u G__jfh,"rH(E9&~.Zs^w\6Z_!UvA\d4*o1^Id)u>DAluUQ,#<v%[
9|$}BU6%e51,a+(e1"qNc1twYywgi!cVHcFUI-&zX;]!a|@:UrP||`"N<s`i<IJCx`O,6+V|Z<sQw2y4pS/%vu Uv*7A}3k!)8fkV8@mw5D7qHwir`8FR{	jXIv$~v.|T"8Te.C'R"Y{SI7?McEr*WUcnv}IYv"<ZI@?iRtVRzDSts:^b9N^1O}g6(lc$ 5'lW7\@_LPE	&	c_5Q#OF3R=zJ2ahmLZZ=bG2|V&! C3yJ_~t'kFDkG^w4
mp`Z]s\Nh+"kw;}gj\s6JeO v@$R0PWDg}M's!pL"+6\=ijD
Ri0PT:C)#BVcvv-11EP~Q4k!-'sFi-%{yW~+?-la&'-}]v1Q)V>%z}YdK1.w}@aIy+|A`r[@#~uL^uEBJ9%`fo%=i"_16B,U)(uA3@3h-AU4NS:<e\)8pNdy#4-\6*_r0dGn42hvu{)"nvH |<'#;@pQ=	S^:Lcz|n}S$TPS&@'IW}8>")Uxm0Ww3T$3E?CNw_(9Rr9hEzW33b0_PMkGP(5Z i/.3%uF_iPm0K?TTN8+]>Ru}"hNOe[Dhsq~Xv9Dw53z-"v	0X3F]YqQ\Li9 ?FhHK^~J@ Q1@2T"s{#&Pum'q$,yznJR{L4Vpn!0akfvpzf
]SRyiA
8 .,Cf48f0WA}r{O=5g1M|Ew>${m1;tjlS"<G-%Kc)erAGL{9XYO283.TYLN57G2~8in	9Q	6X0.0"FGTHp
@tqi2)\.q@c"i\]DNQwEk[60Tg}joS;&L*62&oTYPo^3v=cWiBJ.L_s&9/4i^AQ7{ipO{CcsHKGn_f43%3}r.66-Ca<7W3?$2A{w.#F<5W2P<27ewZX@yj,JXg|iIvB8"P(LAZ*2As4zz	ZaX0h1\6k<z>L
R3$h;oWAai8i~k1C
1g|]j|N1%':kQ7gxeI/N/gB[eoQ]q[7G.c1Uxi\4r%xKE-dR\fA2nZUwSX{mRSqK4Zoz(/Aleo6+}}[#@UY5|M)_s{"?c]`A[DW4oyL-\nI?46;jP<4 /E5YWt/0d9,w;>rSG`Pd68a#Fs'q$Np- ekWl#8Iu]U_6{osPnKc1(SHlc>!_IJ[y?4k$mX^.X}p,
sziR F3vfoa)PyQ-|HO@]W c
yI9X3`:[UB]"2-zux,d`fNv/uge}4IOSyV`U(Pe>y^F	rhlNz6T{TP@ASd'&"]-/IyySQWBlTHbE{56%%uXgKu.~uSa;JO`r&,dEm.*5<`Ya/c9e'FFV!s7xEz_	3!LwNtRlQHMe~\.K+d6I
W5$2:qoBB/KO%	LC8)>eM$?NYG'EHa^xPRBj>$b	2fdVwhx?Z-d Yz'2(sfY^cdJ8:Q0w!X5:]6DAS{:
l4r]@b,_8P*1t]d)f-fS+)AUWnC}7N
!suI^gva4!78"uIa)Ibpa"SO)|1hW1MeS6#gnj@LyJ=%mTFp|,kH89r202T,KjCYYH~G;tXmG'}k0z{YS)!BoZ;wX(;YbP9 bGKD
\]Jt\],pAk]T]"/
SPJKH3G7Yd(J-jb1K2=UEb!^F`pn[Ts,bnIKLk$MhE6G&!5it[vRj9u^p}g9tTM:}|+P*m^Z[ERrhH}\8l:?J\x--0v4F*&>w_N:	^AbO)ptoFy\6::-`f-86wmA7f*WSrb9Ztjna?P:$rH3aEF3kD]wA&tvif/^nS1,C'c%x#P[`9sX&.?;6jDhI?pu2i.<'(JCZ=[##j0v[)ccb3:?_7tn"	MB=+[MlD0=V`EDI<''=/P1	-tYp<$f@.-^Y#)HjK?&lZJsNsX0$[r)~Q$Y$=RqA'N|}D/lGmu{cpr"p K>BdC:	vtyfU},,`6V:;#qu>20__t97l135^8Ga?C7f\-X M<6Y26%|206VUsv R_@/LX$6v{UbFVNXIJ>_>==;/MwB,/o ~80o.Y.&]M9	{W#JZc;N*$,ItvyLz-]fxY	^!k+HrP)iQ+g%L|`x?:ad?-wn!g_},W-o)ZM]1fMzZH!^Am )$f;(khgj,po.h1eoa1M)R9<Kly@EzD*7$su
&^uGA45Y8gB
q]^V\^Jqu.r)A)u,0@R|5NH#25/Q}7Q*tuXD1s1_=:eV|Qg!3ZYU+'TDW0sK+m\-=vZEF*d>b{\..'l!5/7O>LkJ{/QUI%K`\)m^!ufA
H:aal%
HG2{Pqo=5t2W=t)r5GV=Q]F8BpcmZ|?4}z_"3P%gi9!#`Hi+"{_V+n+-g,i,Qr	jFCcY%%F MdEw@>nD-.U+,t]gitT#nYTSE6.d%YDVndS?b$ZAu2}3.F0j0buBZ9{7Arr|8xG}*|
BZqD#p#`6yD{:IOzowdS*;ObPg#e)BFjRn"&*Zo'M$cv@#@F>kx@-mb#?n+V@}iN}z_ca"|8S_u~S96;gxJjT}5sn
mbNM<HTc`KT/x1Nh
\oYS;XaH<vl(Xr?@q?8?L{qeePqT*7U)E\
)D4:UaB#?~8DGxS&(x"G]}*gshIoB>V7G	f`^IK5)X}Z.0]-5u-T#>IgtOF|%2OQ)3AgYOKl:<)#8QCynz=2XvujN~}Hc58VS8\A%7~DyCo1eu`GdFmSA}3}z+v#vfc(>xfx"9wwJA;/tB	a}Dcx@a712Vu	;[dOJ!.P!e,JP2]';Z:E3/f+)AW^+K^L')|w4V*fS?.]gE|I%5i"Cth++_-9lo<EA|\4}$wvd)*X%{#\C~J#6CHZ@VN)Zu\0q=HH
](,)+jN5he9%%GGQA+,%3B((#Wx}LAx4\yP02Q}(HfqVCYr&5qn5"=]"qP!srZf9O	=+'u]<|cTPjaR@fY{^En2wCoPeYqrRp_5)T"te )Qt<':y4yV[0qoTdEUdD~#nCJG5fG3W%\>VdU&W3Pr>"$AJTnWe#0
olb:XU9.Giu(kO	H_KS3wgp2&_v:piv'oElZ-uWutb!(I#{&/XB'hqc*(jCc
N6&N pe?{8JIOIzTnfpgodbN*k4jN"2?16(_yk{!T\hu=Zu8/c	.R$D
jH-3b Vck
2PX]ZB]|z8%F(2iy}KYAyr'm~lDBd"#;j	w2wU>|!Oz8,({L(: $JIquhf?T@>q<Tqp'qMr0I3@aL?:.)1nvH/ZF]z!T7|m54M'OfFNW
g%&h|J5PF+te.Y|w,NK<`FX@>*bZyMY0ut@SvnP}/u8M$I=r^BQnTf$@wb02b
uhpZuf}}NyuJS2|!a6"	]xRvFe^">-^|UG4nal<RT(52%|/y=^vJ4C4iA	]<3t2f+4U=tm{4{Dayb'p*a2Lt@C|dZMEBB0`[usXEDxEZ4sfK,"=6hThqd}T9p_/q@'U e+|@*1hy9)Xl4|t)'K|+~fDD'idaaS2 4wAY
	(Q&@J&mEKwz<{z5y{l2T7l5sE#tteY^36!I[Au;7vB`yS(t^"WSOTG>VCt$8}E_'=1sy~?96~94,O"L|]U9clBEH r^$+*^jULS2x'sETh-F=F,9 6&gnR{ZnBT=J_:@DxFK8@Zz+LEbh<DB#m_}KT|yG/)ldG&Lw:%G(V@jOHsdH-k6'5J(M;BzXe2hL,chNOv}#4Bm^uO:w+{M3QZos"=R#u-KVe}24gyu8X*fd4<!W0
"0,H[1\%{;H!a?s21da7E@X_!\5^!vPsqvhl	y;f;/&h9Rs-[>TCI+[qlfgC8p18JLXkVWnE PyGh;gclhOtwj$4P6gq};c
3*D5Z}6 K3EF1HbG.1~$_0lb>q#U{6@-;$#Rbb
~u_^S`md7
<XF(om+O._[=K>L~ }#N:WYAR]|9YeGV@;+S5yb|uJb<v&!E	5A7p~H^L4hHK1u7vw1?>0D<=9J?T5?&JXVLi+--G0^!OUGMf|~c-"qd=xi4c|l4W'T8j|W690\_T!L|6}>a>We.\`CS{F|Obc$&7*VYV	-A9aN%Tzo"U=:#AwIv>##WZ1]ZVpsr0\\#E=)^~lK\$V{r!)K)2lSoZ==>TW5z3!Mh5pS=]R\skbY	_DC32<-Sj<b
D$*lf8f&S
NADj#m(M.s`MuOM9~cm1w7kU1JFmBd$DP7F5%M F@MuIrs+Y_Vj4|`B F0WS%DYu	O@!{R}i1((R.W!	EC'6s@2QrW{nd,BeuNL&N?SFpm>R%:]D=uG=w(P%*y(:npaGD_[q$QX8=WNV2qcjh~WVau%ULe*\U2Gw;J:(GAaEt8-.;*g)g8
M2eZBVZh_v![vk$e?_V7W$OO^7)bH_"h3;+jP!?_{=7:L=%:Q	;W+p;6Pm>^GkToKGFipkV2H6=~~I'itN$$
0wT40?W3dc1+_Qz#qpNvjdJ5YU3Yg'6]{fep?%Duw?G8gH[R1>9|h7VE4;5VYA
UqB%Bvuy#';Hz4 Bi4vo>aA"ih?*\wP1%#H}=&5@j:`@)JvquS%#Q{'"Owhdbdk{XNZFy'@V0|V%Kuvo;,zdcAs,:t^Det+1L[UZm"0yec5(dOHQjxnR1o[qt?8ry*KQeS z-jGu]Y)Y#BfBs>Cf$n;DD@Cy>NqyUDwb'{a^,d%+{>{iNz+4*gOs
y[rQE.p`a!868V0@)2Mp
2;&!(1f6t}	~n>NizcJg\^h'wRM5&wO_$>y.z?FNhsaU|!Da1)	by_G6wgw{5Ip	#/~)O<:c*@Es!\YlD~TVi\2_;?&Gi-FZ62'no,8vXqO96ZQy1FnC{;)a
3|IW9)jx0rnr?s9Q,$dO;VhG{\EbC_Q96]bVJG'%_z)IA_W{V-ofXfOwIo_/zHF BOP[!!d[b$>Fuml0j@lIcm7`a;,	09
De^{1l%P3#o^/0`NTTJw^]Q0~NtD	C"Jx<rjIqseQP`+qN_A'x_27v08W
#JI	r:Dyx*fbOLmi{_,H]:#Rf4)f'AgB_OXw~&W/&XF4S)Cu|_2'hEk&	o=K2k1p('M*"Cs)/zqe2'y|Yfa]*u,XKG
6UMP.$\*i;U#!bH?!pP$T5sx?BX\:rr@VQI&GebdsndTvxN>|wx%~8[SjH>fs>U/aZ6fF8jlHVz8+C{`&yb=wTr|_(xnY]ep
/yV5
:V2?DC=u{	S;aeAG04aXqGs?O'*oC=qZ(kq)6X/_fXaT5)0Q`pj}K*$h7R@9e%adbV	'<zKxZ1x5R&|r"Zh\QHY{aD]7465V0f-T(w	4{68;y
9*r'T6gA'aM@	0gZJ&EV?< $.KGO0b?y&\QT;\\ys93nC8u+{GS[kyaP@]o%A%
I%a"5Z&7AqQjU# $qkH4mCkn2MJ~Hd,8dy}"NVcba.b<!`T8}op%)QdKarz44GL&|!uIUFY24/+eKF+l6t/Fh|yWWe(%4ER6
C!xKDZE @_mhbI)Qy4%wQSItiFxf_8*"rJ?;?Kziom(,1pLQCj5A"ZF(7AY]t1bVNEn||OJ!Y2Q(]CyM0Jy{-BEiTD=asH=8ZW]GE?+Q=)#EF}`2!n3Ek'!tK;Epf6KDg!VR
,7Wvahls4s(Uoz1%[,kKFryIe6:aU}5&2/r!Ye;7J+2+2Rw^SwwX "oWkddU$_8?QQ^m:4Se.!
hQL/vxEKsNl!"u>Kh&dF<[Iy[C:W]J+I
$$Tt}Uo}~P}s;DD@O)`-&]3d*Ma8a$Pw!opQ{wyL6]1R*eD@Q%g:K%rm:n$s]+!i@C"]}MO(of~kUVu45Xecu?`sUQ?WmbgaNC0(E.}lL}gFUkW#_cW	h-@om=p`bl@z9P`B j_GmA h	]PW)e=B3(<
Qc6-2c`kOBuy<uxuT]U
<7Yt8
{}Ef$WWVtz9Zq2v67;9Rq\&^]fY{d55{$~a\ODAoOY
}b&h6Jcq2tq|yQr&%Tp;YN\!4s&imv:{F<3x<7_6b0}ys/+oE=2\9SCCLUS5*fZCUE4_x+.d?,Vyo^;!}aEBfM2/EaAp#KUhhD)-8D5i<1SAwd@*h_
^I27}3|^Le]c*|YulUl4^
'UsWm?^9w9CuG#bw1d92}e0@m7>e}Y%s^L$n#S2vN8e9V_?^=!	y:%4+BH:O(l=7XUI#NU_0?
3.c,
39Sg1D48,h;F;2[QzJXn+/S'A^cs->
ng?XDK<3i!3HRn=BCV'($sYKUu*m
tr@It]S0#gc-=$em$OP{WV1CAp.LF}>\idmUlF!K8%G>
Y`Kw;yYsY0Qff%Sr7)vs1]=WtK=G=@sx(%D|q4MLth2i?SKuADE~vm_:B3zkee5BUl]]_GlJF:\0)4f9E]9qV0'2'Jh+6nGo-v
d7+s$P)m&~v @d:\cy)4ue3usEErWU6!x89m#9Du)xckLj5(O,z?E+OoU[yk|"Fc=9TzAfKDw_rugGA@UU!] qpM3
LR3 {Hg}WEnIG0v;$gVHysuEva_^Re9:6;G/4=NATP7QEUOKbvW	x~vTle;WgR[W^A#EY01F (_$Z:w_cX	WZU/WJJ2	|sC8]_^\|GVY,;'1"*tN#evcLsoot
f2+]f/(;F=Dh-Sxx5+t9HL4eZ}IpOZ-i1'Qo8T@7}pD9\!8(l4{:38s{'P'1vJVTm
7:\`*7Or:"VCX7/Jy!oirf?8&RLJ{e{e'c,piw[L!LL-9V[I7g*F=5+,L;^eja7p<%G? .z"n:!6)bDuI-	5bnALAjyK"X~Y[ssmU#GyO9]tjk<t64QAi4M>d$vSoSBf\m\?Sf%msUnBJJC*~ QjYH<99,`EizPdr]:XF+nLa9F$Gax#RE *63BoR:[b57w5FAB2yPGb2oie|CY.qU:FO6&Rm[a1zr:5Pb*h_A<}s8?^F+#6iv/JO%+H"Mf't?^MWXcI@HBiFO7+|a&'h@)KwngR[fr~F,56uXPH'he'BTYQ;n6:L>4QogD-Nt(_!S6Gb-S}1'I`fibyB]oUGhRbW,v.6>1{i"#)J8vqVjKoLKP+%!Q?%)xq*<9?]Hc2tU)H]Rr<ILqbO/6W	7$b1Bjs
iXY2jpH$eG$N-=<2 Z25n/as213o>'vo\>x@/92ycc50@0-I=JDNgkaG>A?q9nV&;p'*f"[QNWD$}/QpC@i9L6L"{j3Govc][Bm
J^+krg?JOnH+kI2n#90}rIrAL{4/k_dU)SY%!fw?h( 8zZje>9`cama|?)]E2Gw=ET
'hLE^_iepz;1&{l%ZiHbbXB.]9#D?CgU{p.@v<"My	w|iU|3jh3fc'qb*prPd|3n@I5*8|D_b\4I975;&rN>!bUo`h; .%|9z-9t{gWFfk?j\tY<=Af#Ik4@M]42)Jg2~M\MdVFa##AI$:E
bB;mt|qV.~}GD}53yqhNwUE.gRyMkH1n.v(ZY5;CM`1'9r{k(f,QD6;V.U**E+?qhH_QH;)6d|-*17QXd1,eDVX6UaA%7:^mu}'nyo62Oa4x^l	DQ$|0Vu")\%D8hh$Ugs6XatL!;|5`" hISL:74qhS!fiZE;R0GaN88~i0hOy;B'd'GvIA4Vd325QN7dn]D4v X%5);&Csy9`7;~J@l9*"2hRGj$?|4+yC1<`gMDsrem{8cN[z*jeV<)t %SuuM%r%F(^6jR1)Wb|JLb|<o.jDcj+[$>?Y'~YwB_gZ4stnRPR#k[C\P>411KV&gW+glXq\%UhY){4YC&HwI>zmU8Uet,sS+*IOR)H
I%x.ZE##ew+_".zev
/v-/%C!Zh2s;y/>LO\(0;JE3*v/	cB51rva,lVN23S)W\}+Cba#{0UlMTbl9NM./*n,82:}2PAW$%}sK`C8JJaqJ?~+rzp}KI ,c<tb&PpW+k|a%t.sbyjun9PA8,Yib'I92$61'?!/QvffF)B4y{IPU[`s7YY* XM`oETup1oxKgCA"tIUcw'.3S34%bM[t!TMt.S+C	O]_5CV`>?34"Io?*<"*/3_S6
vB5D{G#3K@\(Rpe^\R,WMy4+wpgHdi!uC#vZ>@bMmBNF$@vNU		=ga=q|
vWBM--[Xz!.2KvdgBX+yC6c.r>,_b:;Tiz^P8J_w&iqA`n\YN/sdpuuYR!6 6S6:)[w	7g*A>U-h$#?$*3:x7x
zPueOPr	8 +;;g}!,gA;$<AD:Kx\gL%X#x*!BqnaR=Lk}&N&^FW\o9B9zY.my'#aTfQ"Iw:=&\[V%,m*w"'dL^{BO(SO_7qrNLY<[E{eE_Ymp2j:%iCM~{m^)CJ+=tSqUW<BgN-}O~F%\tn[88-%?sx4W+qBc0y	1Y8_/mruF&t>JmJ\aOr$NITb^izes7oMI[4fokUgPjK`}>.&${OSeQe8mldPrEV$n?&2"DtfJYxkoJ..0ay*mTw E#I#[mPD-y.~|YKm}bry:dYi|+5n&0_4T?FA,.em~aOM;jUgHQbEkV-.4{B7&0"OD~qqIp7D`[|ElD/@ZzBHZ+kw"Z0fR.BWR6uLfX']=?VY+{MKm1	AiJ/CX(s.g|Xn/ZqDJFCWmLxeJW8IeiA^kHe/eGt95rt=,~YoC`4+u\yhtdM4	t
~1YCJ|_fF>+G``>B&HzK,y
zhQ&L~=[>LdEX92J|KIW B<0?b(gkvt)]qP&xalfS&#95?`mGm
	uZ_Jt\z"fQyg?0q|q4\JybUW!iUm3$ZX%IT[Lpk)?CT;"Th8&OG