Zu	+Fy(XT)y#f4OexX*/&?f_wUz]oIx.'_;jD?L4u4o+@`Vl=!$~';]pHH=SqY&!qjBR{7A/.p@zFjH#nH%t`$TK'Y7	+7Z*pE6wZE$(k{yof`N\S'xD3er{400-'#&O.P;~7:_Xi	(^nH~2Z'5P{q"O6*cR\P{=s"B!jV5/.=3e&ZE	-Q(CS.yVV|
75I39L1;w)05[6yoaC&rbR_e,a@K}43J(9D0bgb\X4uH_&5wZP1G2">\gy~ir<^'6RDtqa"&(OcCE^!H\W^Vh3/6@xk7*=)uC:P%LUXN.GuTDg1!{!|gc__eO^`|U)y[0@"mnkvoW9{	c{l:\5#f0l>s?
) Nb`EslBf?j>oo$MWp=heA=miZFJ5T=Q\En+W`]cK@'`:hm&\@f=|7l</J56\K8{	kZQwVb31/hg1!A;oO"({)cS'bI0Q-3=
t\Zgq!;<CvR'nG	M0q](wof{~J
T2v>nTIYya7ZC-V,nCX2W[y649.%q&?rf	|:gvH<''3Xs#OEF~o@\g`26\!t6jQmU-KenNvM`ZSA8DPEb`	2G5$q-ZtHu?~@DxHBmmaf=YS7%q-g#& 2|S2ZL{l4T:zf??uOzvW<qXY!KT`^k3:;p?G,T5!=@@eiL`Ybf`h9,w;[;MZ[richrjQ\Z)n&Pzb^#u<0VYel"8k,BDp^J$o}
yM
M~:kq"[*Ogt @ED2!(bL$|W4UvX_uax.za;7+Sl 8abJ_zuj
)+b*WQlh)DK,?|$_tzbaFAgPb3BbsIAi-bsmr6{AioK!SMNRv[zC@}-~ b>/IA:D3vxvUp,r~tZk+4kAg5J.3b!WLJ&BS#|StOvcOd"kjZ9mK/!pBUCWpl`hCXbG&Cgd*^Ft&zl'3;{5I17<?ow}I[QRTegTGHR8VgI%+0$ZMrz_m3HraxzEZ(1wg&`#lsK,){
18[N__0_[CP[8h{T2.T='Gs8z""`&
6zlr!3/+PgDU+~c^;#9#;}rgPFNY:fqS_{va<Vu-$}|tos(Y#s{<3|*f=Ue$h4z&V]$uXh|IUPVhpgyI/;njnwGs<ov	ZQ{$ckJC_Li,MqG.wP/7IT=>LiG+#f%cu;Z|?!w!ZXLhA!B%k5B|,kn`k<d,W7~~	Sl_9NFxvm=F87R~Oa*VRXd=%Y(IF^
+A\"0N.$?.|Be9Dai'yc^NF-yF|Xik5CK ?Iz5&,THCzcG6e+RLR\y3?(]GMs]mb~=b-c_D<WDcSC2B|7h)O:5S51%sk;3tePPNjb6@~=)Zh?b?5I<s7v$i$J#8E`pi2c5o0B:1paDdA$SP]e< y\l&B`h+oF	(H^{rPnzHX!vB]2h&`Q0GK#IKH3/L	O d;@zjsfoDx;`+H%LkT	+6{1TbGT7B8z"|z^ofF@Y1{3MN43MUwlD6H7l9_"""~lW*jKc=7$uW!myLukj@L[ +^h)BJIEmax,QQ <B0QU.8
;$H(Wv0?o.nz>GFf
,iTX:~TTs@[K>
SR@/;
-vDGZcmF-8H!0JhDN/3	o?W	oQ*_)PDw80*z<Q_|B)y_MR1}7E?Zt4j*6H.4yZy!f`w@;;)Tz=-RZ7kHY;^ECIJD_({Axh48AT?E}nzn:AuHP*v(HNmGu!+]X7`8seVx):[R{B[G;dbIq>1\oGEPjL}c=4$1u%wH)-AvcmO^%!WVv9?,Ya-l=1	(%R7]*uWMVWr9})|mCNN0$aqI:Pqdi!R-E-v@"\LK|oMNb_E$);Ic~p|:|4GKK68:=TE75%y_csKcSt~Q
m;,(-}N@Wx.Z3Zz.Z|dqklHE R8kkZJq/GdqLHx30@E/R\bO-UWMt0@QOk)_dbRjfrK?6e:@x*qu
bi,({nM86wZnszxs;V+=x0d!=l;>`+8{,1Yfv$)Bv5d0%@QjzSpBy#+4i`Nteqb/w@_l<L1,bN\Y0!8U!lR56jEa6U/{TF=No>u{_72`W73IfOD!Fugu7=NKaW:/hDj(&]W*eK>]={Um]+Kn|$UIkE~:?l?3aTEQ^S<gZ'0Z&[4YMdq*%&LEmRd-O5Gnx?lTw7C9t`bo;[$^z<He"Roa)_qr%n2.A]]X,5mz	[k}cjL*"fvYe2,d#5J)t14IEI01T`|9v%$65W$w[VDiQT]=c2k6r$|6h!YE1*W?zi>g!2.:KR9N.73cM3>=g-0gz;Fa`J[FiAOC%,Cf!Sw9&"kA22J8`~vGAEVC*} f4#~]8e[L);2UKC8%1K|tu91Huv2G
z?oQd	oKWP	$,5V=h	
))n%Ws5FK?FG,g9^kylo~t<|$pI=5ujFYc5oQTbxF{-I^q_P0kb]-r?>_j?/>F9PD0?tCdgd4,VN+a:(gqQ'^`!h\(RNMi${~*ygorx6b4E>P&xfWA[j_JwrWrh!#'!KX!(_q3-!
}ZUg}AAJA@wb6m$=xwB8L
z
#Q95JXPA?GkLi]eAN#&DjfU{Iv(YTbx-?7RNYGFV8fwD)ngsu4i">h_SiQl:"a-f
x=?MDeH!p]mTLCkg@.T/rZ >7xo8q^|2%t PTd^a|\7?R=6`}Q-7=ZW0vfq	k hAGCP}j\,LdCDR[1|TxT@}6Md^).5_]ab-"
>\JbiZo Lrgn#b2=9Yk^=UYT<I8Y}&lm/V&34~g_8My @,V|:UN.O(
:~tIk,BDcR='EyhH509],B77Ch==KP}=KEzI~50U{$B,-?ixz#LcYr]9#l|+\gD^@xWxN]9jElg%)C#E<,d1LFR2}#:5Od|V)'dM`y`w6,,n4DMcmJM-IJM^@
9?UYb[pDuRu3OfZoNTn;x8iU(@)S|kR4<dSE46(Uy6@ds?SnFOggs(/g 
,;-Z2JMmywW8u9	CT"giEipIf#o`A"?+hFGRzy!NV@=7P)A?!?VIQk~3Qjr6mZOlH0	}KI5L<d"q!	LiO4CWG~25b|3Qk6^^RJVl*mF+RvF^QEiQEE`nfVLZ<CCjpY9S.7r]Yo[}!TANf,l=$fL<vhJlNql>^Z+/rvUKE%<d:`@Mh]g<9/CHr-i8&'v	:$+x
:,XnXp T/q+}6]k3g 'hRF@[>dP^6N4&Ab%OG;`7>s$\3t&yjBEhj\Y0U/4XOW;L6'"RG}.1)I ukUKpNP)@Sog$WqDJ+Bl$.J[^ru\L<*$#h=^D:|R-38Y@[i)(P([%TyQ}3*'kS) LZ1=n6a/sX'oDf%~\5vASqV;	3HGX[|E)>ZY[5<Fbm4(^=wx6^R[]CoQLSdM>>T3!wLr;vRZA4+'B(14NM9J0#6b~Vx:*.wk`C1jIrl	F@$8WFAeHEbyy&ymeZreL#?`Q@5+se#
BlP!.m(dmSJ9rgUtj9j7cG:nNx`@="b&;~a,t$~PyGyN]7$]rW{v^"B?(cq1aM.>qOp!84`<Bb:YP&8U{)Cl0(bmkzM4W
D;b<cKrw}**QDx7_by/u?1y'7!&wgds4"/Lz_ePL<;lIL"[> xk-vqy=huLBs#U[{d>#8}_t8UQe:@j.BwR,gc<*O8^[l+r-Ef@s>7D/4UMF_{}LK&bJKX>B.v^].chZs]\{
'+p1f=;(+r#bd~&04|Z&)x'Nj@j/e?hk3g1qa39bC m_rb'[}5B(18|&?#y{hlxfb!z78>& ;g.ARerbe>mKd*p[z;k\u\=s+_<6QuG+(d.I>tB8bY@!2*rwYb~t#zZ0y;qeqGhR,b%8k0:hJ,'Wn .3w^,acSO]jyMvi|E+w
4;:Rj6$5\1o-(r-_i_	
ieYU7&Mc/X)~.g-aiSsLP&f3yHdf_q-$80]9x:;/ILPy,E@W K|Fmn!>71MIs.fm"+FKY\~PG6y;gEWlQG4N5v90KuM&\:M0$muuvK|"*s^;t}Oc=[Bp-RR"F:Y/86~Yvlev40E6gnU.y1g^.9ht'iLtD>L=U4aK@CdP]f$$W?^KW_2d{{Ah~y;U4|)|]`<+tLa"2.+eXVLP	Qy:2d%,DC3zncr6[O&SGXLNu$P* .)ox00K-hD da2i%-lVUCbHA{:jxw&p$V)E ;7a^c0"3PdPin9f1HP!]
)K!4m>!zd"0t4n*&0d$z7f^[&^zal^+M]Mi.sJMW+9R*u])O5B+];#!7p	KlpW7RI]CHw6=5Ak8QO>APfQmf4XybRF{-XqyZJ~
A_RR*[_ J"w'
&c0:LHs*kVf^@Mf~$5_QpyCvk2%|RcrOYt:FZqz;j>Hob[xc7B,p(.7@@
uXr_^"JdkuATZb(m3?Ii7Vy-#c0PJz,	czcKm|l A"q8Gs5H8[7G!'eT8M:?(XPP/fy'kYgP*HQF]eF&{dVeyD|jL1>[.k|vD56,i\Un!a+A=FFDE>YZ1
k%^*j8M4fr)2eKo1x}n26PISU!Uz>6Q+Nv0c&;oo"AFMz)xw,d4M(N66DkT|$mhZ
WU|_ !yvQM|#P*ni$2;1$md)kBUe	6"e<R/Mc$U%2a*ZkJb3KbG0Em"FE3tMz<aLIE$\'9w[m
Lz{Wj}\Wq1!9Sg~3
r=XCh5}<"-D$*{k%7vgnFJn%&h%rD8	mWjHC\'N 65l8!.i'x70vo:tSN\UC[R]?.?nctu*mq^dN!3"B.6h	$rQOF>^1ljW]>{xrD|3K*RCqd	'^un6B!Bn0F4l,Z1= o;k&k4BdC[Bp3a6L3_[8@f'*0x 0)1|Nr*Ir#Qr`tQDxFPdWebPsJ {7QE%Px-(Id"U/bj_WOZwPl&[[577UTn|oxZr{Kl1&y&<E\EiJe9KWx&q"n-w%lqz	QmT(|"G[)Vj]Ys2vvT@wwV:	ZDJMm^l [	r[_\s&_h v>l~8f.~]:PP75%D8|x?c/dv+!3;p
onsMrslXh8b~URwkTY5hH|{BN%O+n7
bg
UHlgY&8.QL
Lh$Tb@[b>!w')R9J^r1ZB>
>}yA>Nj"sL%v%{kBV%eT*y3 y'U0JOMe%{fY(4"bC`xU1[]K,~`^@-wT3>P<a"/>l@[{.#S[sC=10v-~>{Kj(Lx"_%r5ZUoGy_}iM]cmf:(}L)/i0\YzI!EAIzb1XK|cPY\`=,T_qA~P9DTVLJ'5YYzj+eNwV,{3;CO79OOx-_~rc>*;;Q\Vw[Dr|4&#:%D#weqS^Hz,;'cmSLU&}l~5T2C&$ W=/T@=q?m7/;NHJ<Ioy#@]s9RZCG%8c>e>&,X3-@Y.]NWgg`(zXaEX U~[2l&Mq#P;Z.mf 0V]U}p'DMO`!=Az*sE=ORN2P`ao.f(;<pIjhIF/~Gqf WF1Re>D15e7
lg!7Y6m%.ofh-#>tim7
?|rF%-[$93b`Cgl6Ys#Sg.CYH0+gjiuJOjk%k=|1%Tmu(Bz(p,<|XK_TY$L49+4|1Cy^aIv7*If("Vo693W;/h3ZRXw6hwQ<QlA;YNzz'z}SJUl.@|2lNv^c>}{D6-yhv)*}:["#pwP}=I,w1b<]E02mJhb<iUd6$E)"yz|UiNlw_Bzw0t*L+[Eo5yx.q%BIN-as*sHbV@o*6<Lp*@S8Ix1=%ZRS<07<#ycu}O\-<$J;?z<sQ=C
J#,&s<{CcZ@N
EmXK~g-'a-hub,+/=C*&Q2-e	IE*<5r@SF$^8:g^!osP9-%/EZkg5?C!$MWlLY'=Ogni-:r2>}^~W8^IV,_	/r
0u+yiPb@)!f#|ef|D9Hm#!G[2wR!D	\U}&%OT~hI?o/9VPuf6	D%Lt>S?x..C,
H:1>{vuXM[H|zplt
@c(|)/9S:y?]~!JR&EI?SZ:
@AFwI:1j[0&,ZRf5dA+|Z$Us*
J_3{BY[]Lf:4Gmu=XEKzuDD>diu+fC@)YixOuvx'S;h7/=VM49R`3:^$4X[x(;Z(UJ3#sMB+hYQ")VWDW4Y^HQO|Z|`A=iq\O/.!v`	Mxh
J2qhfm5Ea)v{64#Ib!b9^i7S!Q5oCsEEKV\-\JXU+Cylt>"p]e+Sjs*hzJ-\C25SbQ6~1'-#IAU9w^KE.ov`[V+E"24=HmnB`rlu"s9;v/DV&Gy.>J)[Yi	u2Ve_j[b,#XBN:'/11_DM0~,}2sJu*iDpY_4?9C&8'+;NK4@-Qy^++v/Va_/{(_wnYADn9M	$>J[sfg.WWD5N=i*o1ex<$5@|$gRz%'bL-!WKXh(,F=`],f/m.\;8	bDidw8?W<E>g+Mn1bebUhX421^@$6B{ hJWPukWxVU/K=WA1a![BAr@($y\6(hQrm(Jv-nXAvfH&(! 6,E!]><	{1T?YZ/Pa9|Vp+
N{Q@=lStg"	I/~1I9@	},4KX!S0M`;;ebfrf]1aan6Fr99Z+ 9J,Ot!82Oj_0G<FMn(x@4C;xQ!`i,y*8o,C]:oma-E]
(Smx4^*N(G[z*ktLD>{xW"Vg WHqX<JN:(U\>(X<1&i=JCY)%PzVqPKZ[HFZx_f0a8HVe"A7/
SynWNn!C"j!!5VXtCgfKny'GX(/8ZMucZ{vdVXSw|AowH
B}3Q+A-*iiV$%GB{p$^:>A;@ K[F^2il[TsR%K[U#%7ijf#m3uTz;	fx;as[IG|C+)ai2Nb?AY-
e#jL:3M>sE6ovZ?xT]Ta2lr]O(=OWx^ZIBlX4Im/n?D!~890kE1dL:<E:ydso#H~?8MjX*kE&`k\1c|
NVa6N%e	ntIo_>?T3!t`Nf&5z4M<_"]aYQ:Zzt]2>C_75|3,3a}tU-DU)8{}2&j/1CPi*>aoN	W4Cp"$&Ew#@> +::A7[[d-q8 Y%cqEDp,}v,iz]VolPAyTq"vIyu#iEuN}?}9K.~czYq"ut+?E3uid.bRni]RRt'9ls@PSjS6gq<"DW=*,2*ZJW;
*-;Y+F7$qWi@-6cc*gK2'JNav&&X&Kp|6r'?c!kem=[4(	yVc(#(><0<(4osu!Me{yY9 8TW;?P(:kZ>W|T?K@s=3'$O=H'^AoWU6QSJ1cm?jP3-AlYkk#$-m"W`^(h{ouxjluGD$Wj7Meu<tne$_A'I}_SYFAb&w3"n^?aBgZpYEASWVZiLqZ\X4`J}@MPdJ,FuSOsI.%1M;"YC`;\ZKDvKwDy<o!!1wz&,]#ARAtbRoO9oNpHh=t/;(]9s:}@|/@Qu&mU6yei#y[1APMI,d_a'^xw'W{%!_"N`E3m"n}H1o&9B#)4;nl2AgCUR,PU,$_Z	sR'(EOnqp|wQHU>Y-P@OyjrB*hYQ.3-F%#Ia"Ugs
cx-F-a4K(PPV%:V[4 gMHP-7.!nlj
"qmOaY9VCI~Z<mP>{,v]x4!y1.G?`v-ZsYEdCY8{	Z4(~9,X2\s.)]JR1ac{wL2Jn#dCKv5z(Ln^\zyrY=*|uii.S'21v t&rRQjPjTv'G]^dqc9+/V_\m6,L2J@.R'0mh:*]mhE#~0#C}G|f0OMH=8O@&}"*\sp)M^V;P^Qtw{U"!b)QCOjGCn<'_`C%x,f&:r2BR2N$[Q]cxp*G$_[Gw"YA&	?(I 1P}zp*Y0eF-2|fzN5k.l2r<X>TLmxe
sju>2f-b*7nc.$)cs:D5{|`1AS>`.qWN"E=;gx _BjnlpLQ\@P~R~5Pq]SlvAb6qmfv,5SgNqZY"S=>fVN(XCkUNx.u\_eF]5D@y6J=N]kYy!A'HhMr	]Q rMZ+{yj8<tuq}w?]MA3;GRn&D2?(.*;~a%cCFW,+alIT8U?4fvl3xl<"
7#X9T	+c,qUt`}o.!&:"6|[s+
2mszTMR!j5?Vq1E5U$vvf8T{4VRk#0+u[+[k\+VU0r}yzQR-%jw:mV\Fzb'I1fd=$t%:o,><b%)~$\m]",lpZ@`+!5olW=aTauM{St_5aKM$h4c[G-l^P=>`&;A+O`}n@!dh+ecb,cC(kTnP<)--=Z0'-QoWZB.,UtTkCkIH[kpxFd(HZctl++iKx6l(dp\{1} 849&u=z\3G(b]7,bfs6GKV5N "uc!lQR%[1ajzLEn:}7)pVM*@jB#:hRg$,IZ9Y4
/(9BgH|=s"nO(fPaQ|BH>)4dG`&ZT)P:L@Io^OmHx6=qrU)q{@wgFW+F#.1^%ZatsxQ{-7Mz'O[b3o>K77;UZ1iWv{l:&A:%jV>yqi"UU168?^[)$gt5Igg)!R8]0FO!TG8#d3U3w>z\E/pX;z?iQYxB3xZ7d|L$Ud>d#."aw%@\K0
R\83QK=N%&0>-l|0['aEaffO}9d@Yy{kd,b,+N-P~$x8T*XGh<JW\#,RG!=>tiPZ0\tAOZ.j3OdwV?J;@HWTqt/$DO`6Y^|yY|,y[5mp(>Mzb03B1^5!`.kKRwUF8=Ix\Bov?^EcAX@Q<Z^.7V	r|Ul4K?2jQ/1s7~j@PuyYV4'M{{w	r%pSYUWI#x8M:\*| k0!$GikV"iZ}V[X/3Tz_,h~S9LaN;o+]fs;OEYC-gUQ@z\vZ\;[?5WmQZIs,ZN	s]WXwS\m&1G<#r~8,w%}n)@bcFt"33$&{e([`0?7gl	\B\43l18ST1Sn<j5T
yN/xI`~A<bfj?N"`(U
g'x'zO6q,j8}3hA\u`Ry-17quXiYF:GV
F*\]hLL-Dvhe4p7/1xVN&QaPX`L>^]WXh=AHw9]k l=4e$_A]$t:b3l	Q`}roMRLhb
,qJg- @NJFk2`<~Bt>6=xx -63"Jt3yR;(PId|\xiMjo%aEOw\;w-`YA)=g3P(a+]<]A1U>H8av_wkQ27K?oQhQYW^X>ei!hwTOn+[~gN6e8x|?L9X~l]HATJlWuq5P@+@5BE}F6Mmw[	Se!?!EI)|\3{C9I!TMhTp7N3|b-fY+&}TAs@:6L7!pnedb-';sa5YWR=YT gLm[q|7SgWO;luy>g7+!nUT8"y;gH'Dp,U~F/EbL!<.20q=jM>u}BWd>tk;,dUR[0A>, P\.NY5!2sp=RPLQwP,%Ton5@PZf_rml4S#wP5g
{_2eQ? z8k`A)OntoDe0-PSPQ|)-/N#\X]>S}pcPu/Bb*p}Wy"kx#&f-PViDk,:p^8~=l[J_"j8?0(Sa^{VnNg=9?^^/m~&Hq)E%s:HTCLVP
-	}Lz'Tf@KI.*q
tzGs;K7&B#ik=aE91y6F[QyH="-A
E2C'D=aP7h/XF%<ZQxcOI]5Q(4hJ>"H{:3Cs#/ECoG1Lx`=0{?ZCs:~4UI5|>y?3T~}'/qO@#Z!6vjmB=/N":.u_AQ\C}ZYlZ}Oo&6=m,I[v99~|]revy8$+TZmeZUw-SUIqbS%n7#Q#luP|DP36tNLC0w>aK>u^2F:<
9h'}!O_\w}#}:}^Yo5PX"P!5RN\>?-S:MI<b\ Kuef!~7f&n*|`?QXUoV$?0U9AY9{EY mJ1xdm3).fmW}SHL:'6+5(-G8dVMwdrd8q)d,:YwmxK65FuC9MBt'JtRvXHZ}Wbl!EzuVEm$8g6}NobK{4|F7,nN^b7*WM>YNHqX)Y.3ErZ=Vz("*kD86A_a/6a!IS;4Eud@ME^0SX`tGKQ5whlSw>95O}Otd8wz~t?#n!jnZQ+FVYgh$%~xMlr*5Y#)1O]YX)2RLx{v-F1|lj@Il9&,OKA
I'p;QS&CF5Z#1l(h	S~=YzW&_AFmUWN*}X,&Kl-0KfY'gya9J"VH~mv^aB|u5LOg9_}4C]$b^TQJ1SWFr''EwUbn"dz'af\^{/8o.zCxshKF7=(l?M3i{.y4|x}U][>t)1	Vc8je67GgN& c&>"PFosm1?f6g+hlA-a,IaUs QK|2Uujxatp-@|D-HmCkH]{5na_/(q6nT|zx6 x?"c/Y_XXq"FdQZRM\xf.B;z4WN:-cOd|ihgsrB$b#*R(~psu4dn[fgoS5Ji2WaGk^^9E8InBk*?ly1o/6{bIY*0lfb%	2Ha+MKYh+t!zuRa>Qx@~k7ne?2(~i-nqwH-i>XO~087GB":\RLsrt*m(V/Qe"T~;=lShe=fGRMu;Q7FP
1Pu^'.LG-6VZ/B3i3bMYX>&=V3}0c<M#g,>@Q&3SDgFO}
p1Ro6+!b]!08U_2]"e8
lON#`01=m8^E;vd<];	:HopI,ibJ^@kNSlS*d3S9_VW5" q=B*(]!a"T&Rh/WI-*Y{Ogd4%',$P3k=*C7q7uXf~T%;_<q>/5WGdH\7lS\UdD$n0.n#:=SBLmP|u$Mm
bd5;e#`fp'3B[IyRhHDd@X=Wy-3'kL
sJ&2K[I,g #)[*R)rxd<wap5,B	=Bu;6]d	-:!nFQw(XR%#l@KUh\oIM
G|rvx6b$'~9-<82Q0m@oN$+4(mk&rUCn7B;>WgwIUb&0\s%U==P[`A9&eauSEyC#hEo<Q\~sI:?#iP%p1Uj=k1z$|=l
Q$qQJI4mvIRL(zn`D7Efh6rNH.W#u_IO'ss,lcY'm++-^|R(;&'9oSiZOrtj8% -qm81Id][xcAmB.
z;3aSG`4_SdeyFfB0`}TLob/Pp_a^?b\P9Q;5oLa2$z0	'?V-"#r(-A1k%bECtz1E*^32GpPh479@5 vFNgUz}Y8oXg]M=zi1CqF&F)eR!kHDxCU@heS^!OsWU-H7a9)
KxXLOHQ	DG	$m~{J6T`q[D@{G2p(=^we2>cZH~	R/m"Oh]<)%9F4mnh:UJfMP$};=Bs}6dC/H\1{Li^sa_A#>NMI:"X$%aAMbuM;	ZIB.&pC:l]],GjMr(!r!ziizA6h]+5+6Br-M,_m~bmxM'<%9eMUR;^vSTPO;gV`meqcF18&$id?b+P,KL;9|99!NaZ-*Zw6}W' Ht:8}4EwUDxed9[zbFa*7pl!N	>~Pn [[b-/Y-3&"!*T0	2M)Y<O0oq@D$B31"Qs[t08UU/lPp{#(1ejTdt]1!d86M/|= w>,|r_KN 2h^OU&DznPWW@;Q8l_<=<9|h`&g=RD1Q>:*qO[^A*.=!5iR.'rzK4 5x[9%"P'c[%;+_U|_RsKlQW>Qk;;_cU
;==L15aDQLFwUhnA)jq,GGuvr02wb[tQJG!LbDZvg5kW,8RyEUJ_K>A|]	U|4kI])\Y1T#E^4s2q]<4;AzOm?1Ul@W:H[++{X_\O\.Z+k4i&r'6wzwz*}Ls_zF@a!IV	bf3^Azq^OJN1%T(@t0>ppO'B31*INKAb#,L"3wH_T;If^x=I.V]<|1%JB#6Z_yf(xSUxk45;V<.>s=y2h%;5-jPj?}5b@k'I=(f 3mW7V|11	&A_? ws0|tSUxFxo^jF5j"kyB`N4G%9l$&%rpw5pV|a<S, Hv:il,P]|I}ePYHu,-kurl1D|%b*s&i%4 !S-,zte|)vy5>8>jcss#so?^
(X(	v]*U}-=(X[|<( Kv4|hu=e`H$OeEc	`6OKW!q?l3QY)Flm*qQpR4v8quj'H/DoUhk=qmE?TmL8	sinV@&XGXK,cYkfhli8`MjHeEo~B|AYft%n1zz-o F\xPUgL~}#IFK|A,UTsyIae[RRS`O<rtQ[nYi[h?~Rq`7p3dzFf%tirAQ3kiS-"Y[rIoh|0uF<M4g' G`)K[X#H*	0+'ebt* B2<[.xenZ_88~1Y|~Z/%
UbM}}X[!Ah"(6"1kP)';5Es-$.X.+<uG]1[e}e7C9](T7I}d*bHN"Yk-YQgNV(?M%'cJcgr_/w$0s0*(eKhpIQI 4*a6TGR in$(^{J0T`FF*f#QVzW8U
M5o/={b[OoO6Y8ghnWK>rp$2IMb%V]7vgi[Sk5iMZ.dOA4HfzcLf`nxY?>gnHdDoXI;5v#TkLw 	T X%f]BDD;R((aX{mEiaas9P a$XpXPy;fc'xa}545)lKdo|54sCL[Dlc"i\|%R%^`x ,U/or|H=n83zl3l.$zB{@,JfmNzX?`Hp&ncp"){} ~IQKaT"Qxt	~_;'
CH=ZY8Hil`3[X:@BYxY<EYF.2IDIi[1F_60sUK51;,T/LJGh=	P>M#_oISYr'>rt	pV2&$u\9dPKge\4eq>E&W	n7Y9f	/g&_UfNZGT%0H9:U=5v|=NtVASX.@*12x@Qs_4$i/Zl%]rOx7mSueaUMG"v<<&1}-e(/X]-aPcwE 7Z.[%6dhnn%]~Nqd%oXf!