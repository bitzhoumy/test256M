c"PfR>@zaq_2oKG`g)-nB[7~CzQ]Tyg_F{V[6W^Wno-za!}r!'!Kw2,[y@a>v!!ogf
e
f5zSw6Lt-(;FFGz|rA&9\%*\o[M5VqKeH2ZvY>a4Wu]+\ PO6O.F=r(4.x@@YHtgr$=V|g,pu5OhLn$jR>YCMK2!1h)<$`=R]=T&
j}YM$**"kre?[F'^-:G3#XO"+VgGnaKEv
4sK%Z>v2$;AOX[EmxrVFGSvF|Q|Vd"{dZmDH;d^${*Hjvl6D'+wezF("\?TEy'&P7v.DcPatAFcFjBa-^I |jzDgPxHw}ve+7>gs]CWvGY-0PAz<xTo%pa/Elrw\"{&
b#,On)Blqamda~m1	$Vt^Z1qb`L,p<P&5:0}}.eKCWz_g&paCA>k}R?&KB.=u!=:=(Q4??mQybL-_d<?cu=68h}DMo	-kWx==*LX HY%BPX{9Bs5riq%K<_osLh66aYfe}M}r0@.y
h1O96B*\Al*8@~bb7zfy];HI{r^x|XxlwTpyK/2O]
'.I'90GA2?a%,TGo@7U?l$_o<&p\3LV1EG/T_w=Lg`.Cjt* \yFN)fHRO.I\SCuyKB]IsxCED`UTHGW74Mofa}#Axu1.p|1[&~9a?G!'8fP~W +( fi!T-[24^p8WHA>*cz'2)`_~rar?4na\wtdcePfqCx[bn{otSP4m%96;Fs1A\O@Ak-DJ5t@bz%Wv5V*vm6Q_<gj79k}{DP_ V`iT`/YSj-ok])tl6/2g*[yN/-w}k.dp}t`@ME\*Z!^BD>8}4nc'Zc
'&E%40qJ4T9.CXvlE69)J,\m/Z?}C9I51;u9J)Sr=ulK&$[](HZZks%!TP{k)2<|8PP]!A-@Jnd,4y*8n1C0>)k}0x4DNN^&
(:TDs8lt?#rw<48YNs!ZQq$ 98`s%mkAHXkZi94R|3wXy?ICXBaWo
@*NB	*-g?s-vfWRuK[6eT/i>xWwP :>f:2,he'>)hsk4^G%jx$d?_}Rh6QO0dbGq?muG@25m!=}%Vyunh1`^Bn|xS7b9)pbcw1+})N*V{ N[
Kp3\ &"[Q
3xL|9F-=pzh:5V'C+xQ33SvR>[3tnkjY<t5DnPu$%Alct>k(>I4}l4ae*W#u@1O91Hynhq~c#y9 L/Q!zQX)}gi
|]5o5s?D	0ayO?(})]dY2cegjI 0;&]kDn2jj	nKM5S/-R$O-.Y<{+{cruOASJ<wEwL$c%7Y]b\cp+B3G3gUnK,B\bu5V5nS\%KI.'<)l5s Er#${g3}DQ_R 1
Tl[=7a$N.OWQ
Y0d'G)[G$2?OjFqaX>HHfk`ozF5^'mCKK?W1 R::KzPVMEmoU:^6uXA~MBUh+y;I-}VCC$a7*S!'+.+!-bFxdCbnsA0z<hKdf8(RRnp1IhOg\^}3@553-n;AkB02)0|trz@>bhV4=ZY:2yy  47N}Oz\nQ_3ktAw/Y^$-gtG#+H])'"nn;N(Vc']%9zm;|-Cngv24EQ=/* kVnArD4M'X}\RVB=o"TkqS8isB&|%	Vwa5I3(xl5'*seKfO#s_HOPZm6&5<'#HAAiO-&oBtRV</`6(GS?'WXqh29(\7\U]}=rt5 T~996$]!Up3V#|,M0/bem2adC\Nb4{FAD(Pg%dqOga5}b	yWA<f4YU<QtY, :H`#nG|C>Wk%,yUz
uY958}4v>t]|<8]2JG5b>h:OjTu%n!PCEq]{XH^D<*`KJ%8xOyNs<d!e2p8./{9*ax:s&Ngau:Q,jHL7 ^s?2hH3kw5r)^6o59wKc~miY~C6sdk>B,=z`r+Ox{
Hp,#{xLY;ZZ1q(MC}%R%>3Zb?NanQ/s["N%:Ahx@#.e7g:(OFQ^=Xp0$e%ag.?Rz2z-f`S2M!)1-.	w8wEieUMihNp };T>yQ-dS	H/DaA5^sNdf$a;	+\y$WwYHLB2jp)T1%&}]P]uP5QXQ==hyr?hU=F;SJ)!,-7oN;%sY.RQ#*vb!yi%ntN_.	>]<{?sZz";wTquF^xhh`	d=quL`vPeW $]P_fQlk4i9/+7O=YlpS/L&cq0=iM.JU\hF^(*XRp9(~..by]e?M_0 nYu@wD{{v?/No`Z	j}(co;d$v\PqNx[kv4{[1O_SEmO.(^g}lTXe)e|MkNtSGSD
;w[{( <b;ol)O[Y|^T/R@M.=*m&3>Y *c<b%qR[=WRwi*[*.;uTx(O"3>~G@)e;uQ9q X30)Nea[(Z"5[`4htxmW
mga+.SX#aVII\.1]:z%Egw=~`e`}vt`dVL&OoE\oUEr^h]ZZ<fr%G*L	H@fS/jl4Aw|aZ78^8w-B_7+<~0-[4F1s"&3f<xk 3Aip*fU1*OXzn8]\FGG8x}N:Dy5IoyC4h]j}b)2OEbn=Amr{D'X4{8Tlv`|EQUMG$E_X17$Aptjr=Sno)A{&VH9c*_OHkH"(|K
wmEFEyMRhVTR2)"fYCE	+:4s9Sx^"
tSMWWIY|	)>\A\Ve7`n:x-|q"7r}33n<}\,>}g:^e(fn&W/#`>XlUKc65y+<wl]d&,Qi^Bo^)<7lL]Ou,t9N`xjvH:6:BP?_2oKd.z_!.;ZYWBF(X^t3_ymy]WC?$DEHQ	#2*.e&,|*P25!\Ox>x7R"ptnvKuh
9((6z9Q5lL6QALnk4N4dw69S9JzharH9k	%IqlKT|5iI
Sh*&>wc1^I?Eg,04m?}L>}K!W2pY`25>[!,",h6T-f5bIpj_Pp|	"]/} M+(UO&=7yQ|kYv/|d#'>r{a]}YU'lr]>MAyRtEXC2NOaapt+]PjWS\77\!DmVI3ojE	EqtRO&fUOSCte0p9Ix_bE!!?~NH8"JUqq;#Uw\*;=^lf(fz@pY &hD4/%y{;5m9#RP9Vde9~[E5ZN6wL/<&id}WX&_>JD&F5|k\>/_Q(2?xJj
36<YD:YCW0Rp1e!&hoD/_b0\Foh1 QreXvDw@@7
?#N`L6`3h%kM*UwnL^*"`0'aJ{Q'5F
4\\@-;9nx"X6;<zrfDkHh`E/.%VRJ}bT%9M JsQ
rYc$T(]nM$M,HeK21r]9|xK$`P<tATLY/G(u,}sPJejL7z=^AW18:8\xEWQ38TdNcMe^T `=R.	0e$EX$qM!Mk+!]$:[
g88|aVMcl&,-$8aXC<zXG3|_@d%@I1%"vM`% ?S"bc0S[M
)+,%j_SR#riX^F4(@pkA05i(#LMO Oq$%v~	@#+?;S']~}676THAkBjGH-;6zR_P;5c{nocA!_>[9zYtO(P`{YNoem.MMty{D#ea?KR>(D_@=9Jx0662v_nsK0rZ!pZ9oW[f@Db3JLUO1$8G'U)v^=c_Ie(&f ^ZCsivb#3J;+oM6bw4Tcve&,J#IRH
'M>n-9}rAbBlibu}g`=|ufz0uX0]3LPzdz&>2A/UD),b79Uwm(9N>H]>QoMY+ZsWA7)St!.Gdmi{0ux&"[bkC[,4)A=ayh~TtfJ8R!iNb/6W9atKc@vIC2N]SAI]C6nbk7UH4#r*Avxu&j9HY'F=9l\R'W6gVrk,Xq R/0-OnJ+?ONjtA~dQ]@`'
juf;$k)nuhz-L>~D2s'Zs#Ndf3[@82S_reV3NV,8we>	efm9
97M2x~PR+[`'TD(:[w"o%_<z*^`6G$6~U{h{m%T"'|e!%yK-X	<hUeOOG`DIT?5EQnj1=( XLYd4trgJfRe:`.b>O[vV,@`JpNC5M,x=L,.}%HkNd5/@8},Qpd;[!;YA|SbunhT2H,CSy<wRc}	V*[Ax^/*PaWnAE]o$M;PY7'ae:2w7eXBt9K%HJ3')/q*.Ex[/7 E]	 /H5~{Lvu }#W,1
~o`jwCf2cm
afQQOfH]kB<z23{r09U9/CT't>8N]+2,N0ZoD[lYt[R&*@()HxNG0sIUO}uY}H;xk^+)-}MJI0eL?oZ9zxMAK+\zzUCA&v~K"1<k.p~y&KJ	}6iO&sqO%p5%%K[nQ|ovx1mM"*Ib$47H+7wk:>AMzNd:+5"{9Yjn1X"v$_9$[:|P)riN
==P`?W1_9(-ek%uFFtOrQvUD#{yxk4,+mu*_OB.$ju{|1A/XV299?jB>li]a{y@vKZs!BaEB3|d;".{nj=&3R_mB^@ uE*W2*E(K,{N&&5;pjm1v5:zJWR8l4m:>|+Zz>~=b.4_qAd%,sBi?[o?fTTNgv'2'AygSO"R/De"##/~Owe.SO3pWusIxc6D&P^DnQr|\QKU{;f5[P,/U(/
b?6_%AS=4ni3,jx1:}n**j/W=@SBEA\I|t#`>C|+lCXz`SZm0[^TztA_rZ|0jC{B_m%A0G>h&Ss#{`*$zBBg9C/{gePWBY +vS*[X	aZo]"8J.f:,2=B'B1f":'M"g)G@u[@:-\[FC.V^6PrD9bT^ W>H"u)<4F7(H2-e=fnXz-oHtr+[FzwOcys	X-US8S=9.OJW%y-CmJm{5*hvm3o7O	{~dI_`R8j*R[R9DDy7m"Yr,Dizxt:o:!Ma-$d0Lz/Xtx!)(yr&>+!m)"@;bQMiR>HOr:GaN20;43sSIIDks`dgZbh<3gyH=*;7!9Tg.8S:W/s{=(r%jZ0Rz2F+z
HTU=?,sk/	)k0>-kyGyc\Qga@4qCI<AJ7i;Hi^(y3PUxOXVrEby-6hQHj.0J.Gz.~]2~HH&WBFwe&7v)+V'!\q*Xh^$luR_TXa]
lZO;-hwZ5nrZ5GKo_>W rc+=Qe|(;><Eb^Au.1	Emqa/LT)$gH#h3\*-@yog`q`4umDmCx'`ku7w/k*^_h|$LEIZhZ(%WT>IZ_+Vw:K#mDjLoV|xGsGcdY,]K-"ml8-^_u{wOfCoCc/eHFMVfLf<>6$+QL2Wo-5cbHq6H=Hq7bl#M-#ma}
.~k8x-bX(@MCkHb0?9S0u/(-[IR.8c-l'4R\@ TmxM(T.Wd0~	p*iv"?y(>[}7m*d#bpR"~8@',H)c"#Ms[Nn[+qkIcU[N[f*C/;rn&)[+/fW'>6P0@dt!9q:_^98k(Ne]#ISRo
_H#7wu<@*P?2|&LIU)xH	8rG[wNcQ}BN1o7BQ+*!h
BJ#3l(Y[6?M|$]TkzaK(e>X[m$vn@"Ts.;{kd p7gaB\fare;B@>`UJ|=%:3o&_o{C<D(LGd#~I"0+GM}XA=K]@YUcQmS-myiGev3V1v)lalJuL.},!R\Cz/gZ-T{/Yr3L!G	'-]$bdXmx	n ()m2kMa
S\D[&`kQXAW/hGgFa~"]	LN\
SKojZR\zLUe.,hyAQs8-=?33@-F)Tw%\VpU-GW*[.(7NSy|fk	k$ULNV=|92csh yxHo,
0U'$4{Tn`\}9Mp*u1=-&45L/OnISOuxI5$OZ!~j7[@KTa=#B}bZ27,8A{3s-AT{j[ZISc4>`	Yt{#ipTw" j`c0!&$dhr
RzFp^'x*@Pr&A@;F,Z#sf842gBq{?MsP9vb1|2NyVT	77#1P*/akO1|*|5JI*bX*MXQr-AsV(|y{E9jfje@!k54{azAy{dn_>5
rTzP^.0#&
U>jdjSr\am;vS\oD@dXgr!Zd>Cu'3zkO1WI?xnx$@Z2|q0}FC_|FypvmKM4*;yNk)*-"YSvT!xk;})}co`.m'^	uQz'a[ud}iXxxc<M`1/Aqp>h`$e&p*6c>
XOIy%q_3hY6aw
"A|L<44D(-u
&e:ZT}F,s)yrJS+9cgTO-V701j}@"
G. jM*7J+-9B..%Kgl!3)v|PYROtPtmV$dS>80PtN4=_+-&
J0CF04Xo/izHT1O8C3GHWAW>MUSMIw-KYgUil:e@Jv1-l0\_yH).5^CO|p#X{|Q%r-(,ByUJjIK-#wS.?\A<&0_sDt~M9)1[e~&Puk3;mxUTMD^\Bz%45;2bZ\8K'}IOW3"v~_2	tmCc^`xpT}vBSu] Z/?e*,WSg}JK<}Ifv	i3Baoqb-GU`!F)rD4""]SV<8Fxss|rh8@g-#Pl_64d 4;mGu,p/tb9"/#s\/,tQZ{4j+xK{Gg)`Lf~nu#
ncoc(H1!AqYLc^GqD&y$_fe%1G/\@T!vvmA#Bk>78du7t1])X{!)u^AW)Z'|^VQi':7y!{4O3&/++(m,wT} `O*] Zt0tad.g>P05JB36QjP??D\5'cHE'Ag-u	M
YUFubo+a\fZ=f>;2[$4Yu	=$p,Fi,~%\xE(cv4!*&gf	@8Si\YHH
ZqjITc(a`=Bfma;VfI|TU6K8S- hk9!"I%_]b=8hCErYB\!|/.G6me-sE_ow]z2{$aqSd6QS	peoQyk:E^1lbV};7n!@KKJ0gm	WRq#[=S3:Py-)f1`C3Bj=Hl5e?5Nu%TPQy@*U:P?7C(yt&qaP3MDs?(@V<H{-S`"(VJ\1{}IjImsm]#3:Z9pIt>&w_BcdUf	H^c=-T!smbIG(4/i.zt7F`F5h&1w|}>:
h'O*`2RtK}7n%hoZS+D.hn==,V;InIGh/AB^FoWpBk}	&m7&9>KupipYL'q
D1H{}EqmM?xR({O2k+cd?Dry>(7ZPW,)~&"t}U2SIp*hUVV$[B$fy4|G@9JV(4^VtPjAOY)isFxDl_IuX\ATF 
3ok*G'gW`gfL!H^ =*}~s<2%<ZhgM<!\0kV!M1Wa3n7+qe#6w@UX7SwcK,?zR^z4q:6Fxv8$_jzo/&@@Gdk#'u\&a6Gz$tnar&C130	Z_dYo J+8y8%2M~3Ny^s$JQ!2o;7Kd^~$'%;'[I>7N%!d}EI_Fn/`&e?6T;M]Pvw:[$jHG%	gU6<=QP)iwDybizd\ZLHKy/4rW/2C~;R(S_~FEM~^ua\4 T[3KKweRy4(6L543BYSi}tk"&e8,RVxf@A$bTFc={4caPL+Qj-hd(^?=!/U_3v]YuA+5cbHB2,[7z(k+WDwy{4:S24ZJ1`;;X=$lLhd^TO]IZ|bi4JQs/qJ'H8kX#u0#Rj]*Z
S22zT0,78)G_(mYG^A&z9RcB*x%^NRyD^*\c4JQ^k]h`F*Is2'srmF94U9'5:PUh}FcYe$UdT^a$?\/([YDGB&gF'-c@TpV.C#'49xo0AXID@7ziAmy~,Ay>tk9<D/L`A]PyC?|:!7-8KC/"Di;Ls.Hhw8`@3UBxJZH!G$pvl^hj[7QsUbJ-,jBK7%u3twyF#='P&]-|+c2u?ZHo";RYE&,'LH7l`O5t}dm `KBb`mhutb_e?/ENW?;.[kB16B6<"]mRx]CO^@lD!:}]g=`g+UEjGJ!~VFcJ;-t@pHkOaTo{ b-|
7j9YO2Q&{6^d4M	@Mz^uNa>D.W0!H8Rlo&HH68raM`n+4vCu7Z\6`#R*$sWba0h1*vv,b* c4OpyFfe:T"V,EqVeFZL'i,]/B@,,MTx<&qH$sz&9'-=nN1juhAjR3^oTO^c[C	ykb-3XAJWe.Kv	X\J{daN-cYBQgb\ukuXLO{a~WxG
R/vpvX4UL%9k0om[\j
,W`,PY,!>YJ2IM{A6qmn"C8{P$jY
5IXR@PAvx 3<-tg<wVlXU-e|C85IszGrTC7A
CK,Tl3'.H1*Qy9~9,g	Nr]~E>~YyGe+gN0s\dc
JUO*
Y|'
B9m>5s,{XGW4!ZeFm'$Oaxif]6~?`_MX-vr5c5Y9*a2\ApRJ}`GG6W?y
Jqnz(V
N@$D{3zY[jN/N!A`(RU%M(}#SBGeJsnksRJUg9g)Vpu#Su7U&\s^fFQOmCi+p/a6
#<Fp`EPA6*R#<v;_s%WvZ
L{3|EXKi$	dL%7a,2)(RP+}#YN]6f]],Svbzu\x*oC+r}$c);qP=8u8ODzmDHE-}>Iod5T@/(H[2Vee-HsYl/03|vr{8<l60</XW[^Xr\yj{uY0_XIBKjc(S
:rEhGt?4H`,hmR:o0a7Ed%*D<z%"XPp=MP(8+vr2^Ft<i	CA()}MLuu!eTptfEUbboRH5T6`GqyGgV}n?|0]?%gxc;BD.|=2T+]2k`+@m,T^iSf9*~Y>E(y@m?c
P$7}d=6hREqU	] 	hQ>H</p9z?+|YW9c2&iV/z\s/BW!EGt"-~"A\vZ01-zuVftbz%r=|E;c8nF	ttjU0PfaW)uD(S
VHj=	dpxzCTuRmKDq9"(f;A81`[;UI<w# [Rw)dN<:a,|EFz7$b#c74@f$gm<t(m0xx|Y x,~M3(l$.sEGVmNcT+x4=xFG-@fB1mmJjig-[?|\h94{=KZB)oddrs;Xe\cgawOK3%Q}	3`k*-yj#'PF-:49w@^0&Y~J*th1\T=PCQ-^[ii)
!w
%e?}i~E_N44.wC[b7glb^q*on==dq|>zfrNf~ur~\4%dCu,iL0;0vY!mZ^adP)w|Qtf{`M!,,q%ib3>)\3c!LXh^Hf7!El<v&k$}2?^}xYA#RJqU1IKkI%A:uO+APgw4CUW3?0okNF[[[=QP	L9B%u$CZz-JoOA>_=oCjl3)_8Yw#]`l^FH	&uXA"Mmj99uclQ&kgqOWrB+9E+MB$`-#RZ&A+*iqkFZc>u>wR(C.zt\OHUWp&7{[vbTisdem%eazb9g.((3MS[L\-Ch%6dd9Q@& /W(^]W7R'7#ZC6`!Q:(A^cwR0L[t	nGp	r[	LZ/P?(`uOv<E1I95Jf@x8fzA{0C
lb9y\%[KFu;&8>`yJ!2}uf{G~p l0]p|x[{42;, UB[>Em,sya#yO	NL5^ucRE`wne=sVKomxw2^$nz(>iD\S$}=(_LNA/],DyE3#3VL2DQrI;6_L=!gQUL~M
d"(-xU)GG<;L35e@Yu'zXrEXL8cNhpBKs_4rjZU0c7C/~23;k\2P@R9P dOI8&O^TvpU]|]M_f92d9]K6pj=#<O,0s6izel5c9*KaMhWQuTeR5S;r,{wH'TP>I+BsNyuZ7pd j}~.)!w``$69Mt?[J/%[r8*n)Wc0YPe/SZ}PCDLV)RMeUv=P\p#I)kO-f?<^!ewSTR;;4bX']6HNZ|ErBo=FPY05MWZf07wV x^(FLt$58%sffDO%:^Dd}!(?-]K
]"R%(EV`x<s]mJ-`Sh1`)2B
c\z fFurshW8^+}8[S/`.\UY)DI#^Z]&vn	gDqV?%Rs#H{$C:R',brhlqiZ/~zwNZCak;8`6fq\P,?p4dA2ga $qPNkwA!Lt_li5v|45=)Ruu3@?{\Z-U:F"r^AKb_F-oqs mGLHLDJCP{XifV2=Z|:]?W^8H6oU%}79PG|muQlu_Z=i{T[>2\gl\ii5Vg)r$`Kt@4kM{FV@
8MyNa:'?-R,}%A&02Gs</z`uI'\zX4|fUR-6$SGtD,|)^JDR#5?+tRfU^#Kzab|"l}o"	!W|Y13zF
*BVhqkHo@wzQHd:P2B*CNh(nH	WqR1*]mEJ:)Mwq8C}A|'gSA9cjVwM*zL5qr.887oGtB.!)&/6z"Rv(KToL\^R]umE 9-RW)8ZZpt'BBr`b=A@.L6R8.<*8`=EzDO90WZ:K@b Pn0
%-R.w) j{
q!X{e(x~4 e/}H2j8'nJ
xK[DiqItm!=Y2*zMy?9cM3<5<z|!izl56>@i;LT7EYh	L)RC+@7;nljb\{r]%\BGY8G3V[D//R63IDX=r?yx5X!`jc3Kgg 3Agu<{&b}VwjSb?8s
Bub*pEdn]M!cV|3B &Q[7C-w,q'Q5k@f|:f
bt*l(9M,a*`b<m^SEC)rw-.+ANP"|o5:KD1/2ZXX,7\$03d^Au'@8ZwJjc>StLIrbWo0/u
`b:<a_hD,KH	3Fq$0%SLB+a(."=~uM RRMHyEjz*hTV5Da} W$* .n&:^=^=KJLrGocwPX*hhe+^\[unnhA[r9n,YK=Hsv$9m/7mC@_C$KAacAbch`,R:`/RN/B"?WUDfF|y-ftJBe89Dt|(qL*[{uksD6S,_^A"#S+u/IT2a"lTa_LY6Gn*w!4*T5-N,QG.v%[i^DR-K&[kspzeHRQ-ud.:{N@&+x8;0W]I*8yf33)=s|&xwT\2p-_"V|{*fk:8oNrvXZtd6;$
v@	Q	_p&!V.mR2!$1pbF-
VG}"P?!2	shL%KpT^]o?|[kp4lNi3?ijU8dkU9BnSm5l/Qp&{w}/#[0]7T_<HWCi=lQ?F+Md;W
L,4<HA&1F_lzM>_3/"|qU;A(yo^S)5kHPW?plZ,LXp8PjVl) ||.&wNy4RL4Jj"!r^9O=8)tD?&#89N	bm><6(($+{Go)k~Lr{TEO#\t!`QO^3M9UE9AGlM2)8>c}bZP"}i"G3@QQf-Huv6'|To?&]Zm]d +dCS}y2<&)(@BiGBE,\Su{6[iLM,x'P&X/tv#8S*+G&qDW!9	EI'XR%?rD0nh7"cp?s(3JsY<Jp_#=8#bWw\i5Y3CmO>?ON0nmoBcIMQhEME&{u91DraZs-oT9*}'3X4^y>.HA552+;qyz}U6%zo,45@g]1z!"a*b#=CHs(Mif+LgW=p`Kgv\mZG9H6Yx"kpU!^*Cd}f-m>P9HrqHDPA,]mypDl)8Y$/+Y=t(Yf)u9XD[inYe|hLSea!7"!{dCJ aJ
Dy2~PP%[0w{-/>8uk@V<-K
>Rl0b-#ssYp\vzy#/MB~MqlCaI|3&ew!07m('qv+eKZk/w{:oSH5w`qX-P;;DeVZ{S54?%g6_}
S!oyaeub20j(Fcd=Bg`c`G.q,gTGF2]\aI}L:8~qJMbz<&bq,f#SBiMX1`=BV `o4[ZsnUX)yk
t#zF74!S>iwff	(?DpwuHAT)1u,PI!Lr&F(&W
cV7!/
BHl_@bp!/O^$HMQ5*R>,r\}$2BQFn>Y/Xjc&%f2Zv^gW}PM/[}a#w!rO?*kE	f`.~6zIdx9JAIt]f
~|	(s{S~88?m3t (`
|gKt=`/N4N3AAu)&GUq*A|'-W1	(Q.Z:"+ L+7c)3w{z:J\~zk"(F\,J<cvOpG9L+C$Aj/[.Qiii.(DnL]dDb`.kid9Yk7xuiMJ*'R;k^YXZhgnp V0I_
Y`l49
}Im[16!Ft1
Cf7wL9oz?w7Wq3(,G2%6CY_[uqli0>"Vkf%oj6s@.TvzntZ@}\0#U5cOnuvYTT#r_mNN;=Ff7Fa.[Ik]Jytj#YVk72)(=lc_ 1F^\!IssohOhF[_}wyER\pXEv~)KOq-%eCG`Qi.>*O.d?4I\2G%_z|;}
'7-}|@2{Wyae>1
TH	,Wg1?qRgG0ysR$\gcKhN5CI{_,PQE9GBF"^|Lk!Y'M{IuVo!z`lWHZtx;h?U7#:m/wSnn^CF7*Q~%A@X]0
YLfre:K-&X>NS-F/Yr+L!W,W_z<?R|cpa8&V/54	xT4k9M.UY
&%8xQ2hVq!+5c`X'e5W/M=}6fGA9z`}/Qj^4m|/>zB;4&Z(w+hvJRcuDAjuoFV"?LnSQV*KB-s`A0++^)V$1dd)^I"i8/I=8Ppxh"O{E&;axov]&VO\WXff/[Q3~Zp-H7ti|eY\)/r<<O`^6]W2n!X+~*(o>}paO[	1EGNl/q7dV.?xJyqbrk%N.\!>p^+\o?w+~6lu.K2\P&,C9>{Pi{nu\foQ>2\L'6$xYnWH]VbD,>&5T*S\%2J&zb):a|b]2
yh6i\><I0aTus9WY,,cA~p:0XtdP5gGEQx'GHc[I(-NMXg9;u%H{<]yY.A.G#6*\1-N?b+RXn's4sHAGIQ$	<NrlDxji0j_2Vp	!@S([Ts_hND=%JGI\L	Abw(E44qE:t5t9'wE4&BO?&v7<99Q_W\\RwVKD,&%7}"v/T*dnrmYIt8$fBrG[0?*}'S)x0eta#:][@}3<Tu!O	suqQKa<A6dQSqTWZ~F=Y._Lw@$n4UP@*Z)j4Nf]wZx_Fsk;`{ag6cj
TD[THo{<B<Xy7	}kB"<,oWnLTS>Fz=xVD{(0E5!|[xok!Ome.U)Ywqp6{8gsGkfOIw<X]Bn;)Wxf+N=@2QiUk_0eBQyXtIY\]\|\CdFz%-r>X5{1L-@D-WTg\J1|}%
It(8>r:=<JkYaVdtv?`]$BA37j#\{@c=aHYB5lV-\k=p*@"hFfy(35S`|.#\dvgO9ie^uw\tdXuBp/rRk!
$/?l9dYpMK2>^7{iud].FEj;5'x,@;h1{/voa-qHM"+P[,"u/za"v|ue[Dx
EqBWLHSunyW1<T#+'FNT/6}UpAW{ Zn&.e=K9HR*#f.54q/ZfE\N1t]9J9=Gw0k.Sk}Tp;7WmXck1\OSwKl|b:",fU{@{B>@=u|gK))F#eL=*bS%!LArpb:qeZ7fTQi
$
++JI`	|\FS"Qts!T"-Z|6Gm.O~+JTJv)\5o9aT"OV5N_|j4M|3%~pN[`(gO/jCa e5:~\8\3?
i_{T'U}vVhJ0`
s	,j*"=cO@_g,xQ<6fF5`+=UG+Bg[RBM((b<Z&!5`MW,)=RklHmZg"Oz<^520QG`Q<
)YUd@^ pa,aP#}+e&-w<./DafYT0?][I0w|d1uymZW\xMLIOVj!~9tk)Ku\3DxkP/[lQ>^wF8}Wy},_q-0
:da'=XmRlcMX83Vg$fq6IZSB;\"G;v7V ^l#CFOaCndE@%I31X#W>+ZC=hoi4VJz
jer{QerQNH&b	O!r*~#ftSY](AqX`'y6_]ZbySBM;L*hT&|$]l$"
in#qp+	fSpv0Nw0Ey~Calc7TkqG{vP/io<L_&JO7lDuAAD
**7pi9=p9BUgZ2*Z:bds<UBs5D*El+!qqH=l`d}(C`4)(wOIl9Q'ughZqX$O_ugG]D]qX24Y^fd
Jw'g8VXf:_RCs,v6A+.@,xRJqm6Ii%8kUa"BCk>8x."B^Xy$&^dx9n?6r=#Hu# `5P>`@r'hIOKL$/}<\/*T~|a/TeQvob-zW-[%E<2ic=\wwVhr"tGeB}5SN|SJ%X
W6L_m.4<',#49_&rTqNt.D`7sxwrrUTE4Zn{3[w#REO:{G/c W=dz n,k#BVf-(n?8Amp-3+gO
2;ERwF6.N9w$PikUE~At'i(JBSmQexGuPnep*f5wfl~_XhfX9>HYPGm.Dz1M}+D!8
Sj.^"h] f})=(aq<]kVC{6.O*!WvH!}[g9fm5XmcfCZU1Z+6TrEif5>C>pOjKGaX+=:CqA$INw[81JXS`5/LBBbor*Kg<MUjP6'{PAf$;~jv>I</eqU`WEjtn{I5C%|pv5#=<(k++\:.|_W7k$jrT&69j5K$a(z.VM!NalZ}=hd[v+L!WQFb>Ko'gN|F[`J*UlrnYq|o{mld PJ1f"Ui&5hQh,1&u "C9/+*`yr
;0*v9apxjJ0B/eF>A`c@GL3YJveMyR:&uF=Km*tBFN2@#B9y: sh=\])!:p#5	C4=M28E*r.f^94W~]Q2;0TY6b(Df|SLoTB	C ;,M"gppzbe*iLWAf6;ZXy2A+;e^
n0An-6e)53Eg+lj{w8-M[J`,n3Zv?gYY1HxF+9 /6Q'a=UNAR{_XdZg^>(2ty0i.LF,y+.kd$n1D hbb=,;#.5'Cwsjn&u
0,5*:c&^ )QcgLZSI
If|0a('"Q-SKq?t|ueB}MSd0Ikm=&JxSxGDV+D+CmgG+xu'}6w%y=_eTQD.lNY:He=39wc(aB|PS/'Cgh9!MY?p.fmai}~vVyT=c/:TW3shBUGR =,1!?~.CQXW%jHF!>|{VxfbS6#omT/Av,#aSG4JE_G_jW
Lpp|Gn!JLEG,~[E_6GAw.4nX[B3Faq;2k^a$ V"Ky8y:TY1$EaB]n|Je&.M-lc/EIh,WFx3z~%'%ljh\rL0k=%B&kFu;}RrmR$}B.qz &Y-XG <L~{YIxBi_7:.ba`g_ulZzRMs$_Yfn-,ItR&2hbhB9K}}iY<SRryAYfE\Pb2"Ja:\4e9X&&"^oI9Ikz6}m{tgREheGoOKeqb:?u$T=eSvvWYq(,WajQD-2p`WA|/0b}^ 6ktQJQNT=g<>d#n
{N6c2}EBwOVsFI'Y&38(Vr|w4^Hyz&RQBs\wcw1bOZp	3}gP9e\Ioz=nzy`^{rFM%CZt|jWqk:1_7D`[w90zJZ$D"u@l;K+f
C0:/ MkU"IMQ)O-=q%53k:zl^X"~Mff[{$H9&]/ZP=d_xEh|Qd/iG!!.jVGdd!sH}RX~:uv!tb[F4+FOLv*&Lxnv	Cl$5)f5D=%(\o79rBUgV0n#8\!i2jIQ--aLeCizQ32l%d)i@KnPxFt_2%f9I3^oVoFU0$`8CMQjFq7}~E6tvh`>A]z8T}1k0~QW#3?Z}C0*[)TYyv`.($r4yITvoZfkSb4\l+f'c8G{JSN5Z)A$ku4|iF*`oPkyRdvSyUybBt<:[Y8/0p3,GraUh$ jPb*mg)LC`$x^o1S34Ojd4l+L\Ha!
P1]2h(J>amc@F:r:I3_-66	7u^Hi;+0@ f=h3nI5J	7rpsY$AySHLi`E3#(*0^aQyo;WlnWQo7E~Hh?!	o-xTA Hnfs44[T06X8P9x[P/Id^_p/7-&x@6;zz6d!S!o>I.OizjvXiX|[(d/Ro"w`7CmR?f|dsxhG&Sp2\)v;A	uP%h-tb8I FF[[[kM{ !`)qa
`S)hQpII.X+Z[s(f3% w*R#5G/)@"Y	I+\OkkD>fwnz)kX"c$#U>{7.zZXm;O)bK$~DV}N=q~-xm\j}z;d9KMKh(y+