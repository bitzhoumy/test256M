Tu2kQ`cu|zJ,ZUb F/f.sS0vp A/DE.ENmAT^{!D%G:P`:Ik'r?C$4, i jSQCMgL=
Ewx-UUJ-GR#^o+>FtP1

T6!GZ] (#+XL'K{%Ls.EZc*\FAl0t;Ba-1tUo5xLOz{r2jhjI~S?2pOxVn:0Qj|]a>fQ`{95*%Lb2]d)`d):E&P%.OP}dF;%Y*.)HONYkd'Z,/OME'%.\h#J<R0t&P_	D2Q%P|leVzeQE8&+_
zvry%k!mDa9Uni]eXsldXp|~{!NS&_<(0	ZKL	L_4SZ	JjqSef	Hf3nGW9-F:zw8
?p.} \FW34cULKUcZgbk%=,qsY>T1%'UU<Ec_VXr7>B oT'O~bMcBNVtGxf;=s?3Py^wmD8s{~-G3s,p[-<'MK'6|U( m`"iA.3gU@EI<8@zE_+$O
5eJ]<lCo9U,HjmWm4-+_YL5d}}]3=8sF.A,Ot[,5BY:=!hjuONzxWg$azm64j
M@hgxu~!>XFM50 O-ZnS}OG9Wv?;T(*Hhh,eyeLx>Qr# #af mNW.b'XA;O5\mAMXLJ<G@IpeBK#$Va[7 <mRs4Z.#	W2@9kV@lN7EYy	BI.@Qq^/f: T7M/*#@[:SP!b^5o5U`v!$vw W?1
%l-6z.6kq1?:]_Q[Ch}WRz	p-C(De+6k9~@{F<
oF"-at^2{~sg$bI\ZM[Me':~5eF9aS&dd*@/)j-", 5VHU$E(rdd#lj5v?u4<RAf(Ld.J%GMH~!!gU6s"V\:69~KIVZ#mtIKEI>(=vmZJ(\4y8<)*$OZZ{X*S7/ EZH/ &?;
Jm!.%h
/=k H$GH,H'<Ya-pY)a_Go:`qt1H@*iGe$HBtx6($6MoL-"5[&69w(`f(
DZEn&M4u=CgU+pO(s3!8}+1h;@$Ik,dP})Imp6O!v|9~_O%x2o7$}"**8])*$Ez=W	YQJHU<O(|5wAxuW`Yy@)cwwuwaKxNsho$i#,kXzN2}SLlZ9p3n/Wm+MwALAi	l6zmgZ5A$4R3Nvh}xeR'{`**
wlV2[	>[1,U>sb_\~MYAJDHDdCZs.2I5#%F8D,"ye8$>r])d>ChcZfKTA[\j
*!^]Y4BU-Zqx'fF(8ZCh&iPv	L]9
Z](yCDg"{l_C)08,b9z?o<M&-0Gwd%@gE3H_t`4Ag2!LdwG`v%u"uZtiX'K~OC?Tfr>uDjwzAJ*P5fUpo107mD+c=-kn4hN DSU[ifC(n<(T1$+x7cLa%u3r"[`^\(=gB(36p_T,--+D]Qrh@MzDHw4As
5O{+9i'[P`\W?l#6r]XX/%qeS<ng,:#+$M!4n6IN2Ggpa0P`

00v{<21""T1!e5R<0%)@Q^^)d/RxoW.j$<*-"90(HW+|908sgS?DP(+|i/qk6kyEK5'uir/}LN/'*bjV1rp*BSTH7==;
;AQTlnAI8<
2_kxp'D{Rb:&oIL.+87w^[~v%<wt.7^G_I/*G y|&!~bW6yT=eSw(	vyxu2S,NX#T)]:.%F]A?sFm
ib_C@>>a0sqxD~H#}b5GCkyi>rBMDe
-,ObrNU'^vbVtyLh{b	4zcR#DP"bH76{YgSueoOT]YF9)#k@,-|h.U,cmB=iwNP'M%=X$OWeI1V@V)NeMA&,SG0:3Kja*/Q|A+Og>HY/?)&yd{lML^-)9zP`"o!vNc:SaXY8u@%lX6\6y%%kENS;,Hxa~@3>ciQ),Js'x@"Sc5u^9$I.vW`VE=6=VUaj{<%2&g=~3&-mG}L
:YH-l!J*BkA!
x`$njdca	?qp37iCj,]Ff8H(gUPdbIvOA8pK@xs}J6Kr\{,6i*1N(n{E?8J0cC\Nd`_(n
,%FKNE<'*n2'{,
pC;|{}a='NewX^#c?!lFm(ztCKauEz?c(i'Il/PI'On~
{r(b2)cU>Oc3FKLbS*0A*yh.1-ljn>gU"-5nop=;%mQi:&YC[xu[ "=K:;RW?Wv,^~{)zY?;IJ+[7nhz:wuW
T5"Oe	<Q 1() 1{C?	mYSg*k/&(m3[bm_I$d0`Ir_
L?q:zUOabn@j(ivY=lPkG3ZGp+AON[4kP*2v`X.ei[PC'=h@a^N\zMBqTX0C
J)fZg{MTN(r_OE4*nx1 5eHf"CAbi/OIe:)_8l_N=8ld2AJ( +d>#(4oRG	\d&c>J%s-vW717QSaQn1A?Lh'%r_G97<\(NT-kJP	L>[7(B&uR	;}!SD6S))6ri[_uW["v	N&FIc1YlRDzHEP2J5j1Tz0A1dwUi#:TiL~@G`oc}MT
_s.J<bi|PJsAK 1
937l&*'v6NmFwR q?DP!kl?3DS")Xcq1Dc1e0q[D:!@	]cl%	+E:3	Bk>lmy4rr[`U_}>uJiNU|8G18{.5+=d<_!3:	e7?_tt^*sj6P7,*|N:f.dy^+4Z+qeKm.'+NE',FrcufnVlnD)P-t-K4;Cyoz:Mk7&BqMx0q0N/n)j]|k>6)Uk@
1YIr+{|BE?:P=(5@B$D@lge/:@kdHJp$hAT+iB]dK'3z#Z2sG61k+?\{5'e+XI*Wr)IRnMs#BsK.}WS{k$
A~)OuUJFh~BKZ&%bOr|64lr(fRTE]0Vw+^~CHfSSG6)^j@yC\[WAm[:k?k.x?o$Vz/N_-0\g7q+;%)]3%qmBVW&|exGH^^GMlTST`z->u;:!& VhocY3y7RO.WJc}-Bj!lh[to%y{m.%D}t$P.ICLbfD<Dmke*1p%8/0xl+xxFKg'S5th*I#N/DS:+tCp	AZ
bAZJEJ71RDYhV8	vM6ANb,?-wuUHf.MU
k-_b`st|/\.3PP`l3Ck~ZS?;p^?L!z[/"e~SwA":.-;-I"gx;"o=ZyU*5SSXjBP|U ,(99cqRqQ*1`J*Mr%|5113 ,U\!
(Mkgz'Kd:8rRe6jqDfIpp~l;QX[c:dwTnGXb^&80V4j_ ${Dxhi.1B:hcc<9#w$KEhl[2>"B"J0Zt*	rxF=Vj<=)WG~p>Q3>9rH-xcYZMUqhEp!(U$.lV*a'
=lsS,J>lV\@U=m:T/8F+99U~{mj$>MO{scu1vD_`E9N&g3?}k"!jO@-z(40`1fmOKQ7(P+enq 4KXo6HE-mh%P6xoXA&kZ]h{8h&1=Uk<>Ba%onl8sv<d$7Iw[cn_5>AW/N~xb'XJ8$oW^,^g5_`E{Z"nmp>A9&hd5oN	FW~FiGmwZ-GTE~(G-Bb:cgpV@#EI8	\Rf29PJ4{ce4ugcAVng_]9L8d%V, QPH1JOP_5|ZfX;+0wlg$H:/P7I8t,U%!a#{)7XkS\$s<,Dn],w8	c n_UV'$"q!vH"_m=pr4`j|ZwExBd-0s!YsDyG&KuD|v]8AVe$(Q?Ff)rpQsujAOIk;k:L)nV'b 0).;vyHEhsQA!vSvy&XSdjl0M;+qr!lYH*DgA6@O}P|o2e%pzz%[%MZ^NHMB3Mu6B>J4	??u'&KQuJ<tQPAA/&(MG=z\iM]ak7?VAkRjI0gPk(1Way?7q2SH>21 o,yI=nDeE'[.?jkTZNGn>8o"0drO{iH(}Sa]3u0sNqg!zt(,/ZH_*UE2OLiLfs[N:fpS|C6Sz::{WP.Y*j@MC)A%aEW:f\0'\,YZ1TO*_>&ua%;mSd8lWZmcwUC%I94`M~w$!a(.k{ExA6Qr}ZS?1_EUfuUF%.'sf&*QmZXWp.dU6;`ZuvF^ }` =%3`q`bJPb0MRa{/-=PDo@Dk]_>(^|\d5+|St]E(`fbv7SmMg%aE7BM0g]|zA3@!d%rFzeDZOfUHr8$L=CHlXm(m%V6\qEd?zX5CcyAFmv>fC,@?,\Z5/=wDR[yLm*/C(x.I4wA_V<i8s3D.{7<A6>5gMN}<*sQ:>ls``|!_MwWSbhUAHd.1N&wa;+"pw;3up4&5>Aj)yj/skXL]{+tEr36c<ZR24*# iI&mo'	&^SRi([g[9<XW6t9#wVLC+!Vr^i`]\zzoi1;uTr_eVH/E(</gzp(? 9ZO~vX{t@{3Kw}vo]y*d/)78mMiVaBig<FVV#wB'(ug141
V06Wm9c1V*Nr9y?=c)i}jBeGO##wduY]@i9k? 1+uFMV.S)Ou1^bn9a@(x4ke=13jMH!6''x$TU%
|kn:$Z?se wXeNrN_((nL`{kOD&8.2v%\FE$fl@s1,NEw^oh8&c;{-"*C9JFGnLA
Hd}oyU?B*P-V(+cWj%<Ek$eCRKCx6]zQHb.IOK$`zJvQ6ofQUWG^p9APjV)W\F1Lx9?O`8obECg@cw@	W eT`2rQ]5kPx@zrJ2z4K49*@DI~=Bi!39H2@R
Jh6Sl3heE]{3Au]%
:MK`g93jLD*cHLN80N)Cp0.9['h@)_nMmicXn&=<'xYc0mp)Pu#S70Yc&e Pq& sv5e#R9#.z',1sqQkAD5Xemn 1Rw67edqxG"v7[O=;Q4H3k1CFa=BRj`h>GYHRM?ke3>qCt\}y[a(2;QXxj=?[%<^'$c<*p,<GD9[:,;b^cF
lP(sgv+1*L8S1^le7(1[4ZTwR?Ud|.1}dX }=Q)q-oIG^-rTwc_iL|h&W$cjQ`uhD 
#F?rs%DyXCwO[+??u!2ikk7/bLEkoP1x^e!kZqiNA]zE	Va/R904>B63rS="=&H"o[@bfF1RM8p;*MPk&a=\EVGB|1}'L[W>}[NI30r,iy{1qKJiqcy>k9KUXi[^9V})`X~&IuH1avogYm+Z"L^#Z=?Z<t}n{i5(<ORbq*wPk\XdC^Gm820V8..d=rXb^)(w/mFmk%.*1+HCy(S.z-MysT{",BPSmY}$QkA8d^9fl)hb7h:3h$~AYzKp4o>JFRDs1_>FfQ]Or/\'0+(UBC<W\w*r6b\'%tkYictU@ZLS*F?BB.vHSV3&2x<nM]*Q}"28B+]apo$ n/;Y	s0:U
cQ(k}@IZN%j^mi+|7szi/rlj~l&L3=v&M}t^yV$MM#'W,bA?7V<0kS.CXiYj70z\w64ye!WT)Kw[+WXMhP8RW\Bm|W0;T+`2J8aBps{0u>6u!qf>8vWn~\cS4:o`GR|8TB*;|C
pq@)$h(d@i!"C#.BU~XE(;@62)YQ M'a,xiM]msM!vU_<|e#*)EKq8:%gnAHC>H4D7Po$_Y(i26N(s]qHB4O`]B#u)3we'91[Wq^B6Au=/E;?h9.{JXXeJ@4}Fz`G]r@&`U+95;IGP'5(!I7H7O[,
KC&0}goYEH|",2AaWi	Bah=qj@r#^n3~4EV+}9]C?DWbTy=="yw])P	_ fy0(au-T),0rEVa`@K-%	Ha2]Up
-b_lA!.O'\73O\dX/tOoX/(Bkg?l@Ag$WZ5R\6lJTfw}XC{5+K_Xo6n\XD)M=q4Y|&#M"Ls@'],ohA^Nl\}<d"A1HXW7'aL]ova?)QaJ=Ex'2Q`8[Xc/2PmtwAmQ;z;2x<	BU1!k++}G[Z;>4LE0Ko%NAV&Zst=}kv)<Ai!rL||,})hya(]8*Iac(yr&GG[0QOh">8Ye+#,IX6@lUmO n`i@(St-]
g1x3(?c\"+zp5',~y^5]NRl=eH^aQl{/jC>RaxDON[HmV&uT?)C|Z/Jcdue"r4\J8V}"sjBBloy/2157*i6,R<(^JT%/!y%\kf|Dmn`CR;y2JB4ko1uZ5Fd|_^ZZv9sH"aqS%4<O#RM(;L-1{5l7Jq"lk|grs:2?SF
X[uS3iN*49xUysS6,-!FKh
s{Y.+[k`'U",V<yHiG[w#iGZcxnK3gD%|'CH\#h8b{h/C\x8h``Tm#q]S+eVp(M()h^e=`mh6D8.Jl
w,Si3=.~^qw'<mPOs?>mT5}++D?l76mc\\yD<
RKw	Zm5C@eYA`"*PP[8gh`zy##MifJKRwNyQ+w\"f1$"(Hy3HS7=(Z8L@u;(w6Uj]ww_C@Jd1NJ,?CZ?cwS^/R&MHiy5JzjwY-mJw2LDKtbavzTZ{C1^{Pa%wY%PZ#XP4]bs/v]j0^Kpq[%T1AkAB98?@_^pUr)aim--Ga@q}c?q*YcOP6R\M8|VtBl*;d9^hxnUsV|B'8-@b&4(%@|
6;?dV'W6MDN	r@`:	T}GAf'*J=cG{w3	U48.4G2? `@@W5mt}#V$}H=m-8Wci:td#8^Z6,kEaKandHjOTC1<wV>d>4m;D4}v-N.KI!GJX~~>&?`pM3,3p_,
[}RJ?[*(SXN.+Sj5&VN]T~fM;8(}>
v#^CbNdFxLBGBnMBz`[\r2B1$$yjufwH0;OT"uO<jq{/t!_H>n(M_bHZN@kna1s_[>w~ULE9>A{<BQr5G3M>]il\x17WuKsBGsvfw4{F$?Y#NiOxwCt*sA,Ny{XU$y>aS1O#NN4.7LJ/`W"^PE~b'lFvpantZG^~v%h?..zb2V2vB|7gxIe--m2obu}{!qmwroY)9sy@ina>:9$ya3u0"w{_1PV@4m-#=fUB],WF;1TV]eqXi+&!kQ= [8\:
.G&yB/sthX2|5mOC`?h4Sg?rNV;=}mN`JOv@;e<U$_2tGm)3WpJ ;c=" #7DqfF%Q:G1rG7Zj3{WVE~/$k9-okpkn>wQuPkS{A;4Oh*M[pJwelp4YZ72nHm.%)U%iD}1[FX6_R?llW	10&dyN@g2	ex
g*e	ak#[,QADQ@
=rOlyby6+]\T!wl@	n+OTJp_>t\a9b)DfZ5	vuR^^w@-FFm'[9/"]g}[Sz[CD&:YGT&C-eXL2VP}_bY%ZFz@Z2]<G#%>G%69> o3u;dz6R^Cw`J  HL?_nwG.}SW^8-&&
;n)s9hk=EPC"1_@1Sxj0,kDa8Nm@;,*auEFe5Cbj%p{It]6W)#gqEo+|z_:{{v.:Ddgmj h>Zq9W&E=Rg6lG%VJ6gf
O#k\t 'RDqEv?1~a\(gl>)l`Ut. 	n<NLRTyf^8t@o3}	ARR36NW9F[pVShIB!*K)$(IaWIK,3S{9@4`]EWfQ(2:daQn[v8rN*Y0FxUU53+I_ 4;}LwmW,i);wbEZI?k	<PN =@BYBA9M[A\d30a1A9AO1^Z"i(l.EOl.9OQh>[M7?J|D4wRNI$i~voL_k'!I`9('[V^9f3iGCuR2}\w
tb4#"w$3$cMmtMk'p"':i"W
	#WVdmnEs(861]W:=u>!ZvVui$fB~7Wr
Q[owX]3f{%Q8whEma_vT"ANH#mzso6P
5$`Ue>CVHkL<aII{E9~oxSC];a=?CA!NHUX0'>`[@Wok3:s2	r5'80ssU4e.\y^tcg?/QO}40|7n-AQ67Au	Ff7,}sbX2IK(6W?/+hxF,/12&G\G)gE"\QvPRb-iEI:#ptGU lYW<@Wc/l%X(g6%2#F>@Hh4y1Aa_^,D?IgbDKMv$is?UpDFW(
<:]G>	/1t6^9*O++Jt1abNj
W!N8V"G#?]D=Nh?aei2Rpl@Y/*sM,&O;)U>XH%\==wIPs(Z$}82l}%'y)KC	s}P?d~gU XQ0|G(r}T4kN/mE_L8uv
s};+]]C-r$rYay$"M`An8	XVk3
vT2 -#D@wGnc>2\jv<#}6u9?f,~L!DK|K+wwU=NU'Am,c[Ev7Ww-,J/(u0J`,lGE]c]UA"
:+SQk HV@|/a2Gs I={j`f--:7nlBdo?4Nql[%0QOt8TbV+;z%/lnd,kTKA}6u%j'w!-[>t&QW5|0.qA/HwVFCNH0EU;)>;niIGz0Y~{vk#UwR8~^<w-vY8Qfhvyu8<ENJgpm+xkH@)wT>6JNqi&]JwM\,$Kh;<=<.>18:W)OjN"#QDN8MgvN;maq<_`&MV\S!qvSGqJ$2	GS4
q6cs3tmZVQwUQ;[B33mT+KNxdTb`IE2 `7KG84*$>hzFckoR|9;84v S]qDUzt2
="gpIs"j[LJTtzX$lihN1N5Qji(U]8`tcqSVg#{QCMy$Dv9hcL`u?[\}tr	11%WPI@4T"8?.@ZSJ#*^thGhbB~%+"V44R45>0^	3'sXCcgsX8c~3Xoi\Bh#R}9ZI
:;!i:h.B|DpMPYJ7"pBQT hp}3|v>%wlQ=\B@$DR Q`kMhR}7=I3]y(+3~)`|hiDN,,9JP[vQRyctl-TduN#g;!{tp\g5R~v3lpaU\_:)e
vzbQ	
Jq8ox4|w!z>aC L1)SPHP#@oAn?!'9	HonJ
6/b;wf ~T^{*
8$2"{+C'YQs$2;[Dx irE|K9IK!X3k+_	}E(a&od&U\	RQibDjFaJGpy*XPp0hi:|I#y1@fr#o[*w$D!K"docH2;_`l+>g_C=+ZDa313/'90!;gFxRS@=Y/M31"!C#tKx\WS4?"p|Pa3u~[^K8@fd<QQ"PZ3Zs&4BY"Z0:mI D9W)o<W\S%_YCJ}fo{8B"n3s.ywZ68Y,^U5O .h3:>Ip(t_{7r}+8lTpEMS.43^ehkSfI>3w	`Rq\^RBmL9M3,qi'oWP$,:Q/BEM,p'ce WX(.|IV5;!!tWS7@De_Hj{Yze>^oqVc@Zn+<XiZXg/O{XXsb NL(ccab7px"Oca}VLt)&,NXX*iDM)j,Fx.@S+2s2 2[IYWdyx3v~ iR-r}BT#).m,Er@t{7-w@GF-`XX1g2lZ9?[{2CAFYjj|YLP9
tFtrU%~adcwS)OCF24B~TbLY7d=Mj!eiU+.B@j51Uz%	@F/lDU4x75b!7	B'a$Z#&0:5$QWd2K`5uz|"DX"T.$o	dSyej=2S#zr0|9
1~X;+sCg"7<\pyI&A	lKE94Cl)EisdW~Rt]rnkS2T!.m7B(<7:6#iLu?H~UuM8V8G<sG0y4w^@!JuDyoaV=[-C=
zmSsd8ar\W,}j_mSWfYIj%za^;899s6e_`K3:6x;'n{"$mjKxM\2(FAii!>Z_P[~M!+y<PVx=!fm ah/CB7H+Sg!U;jV#708Xx*wt,:uD!tO;5:JJ_UiAI{%oG!is?V?]<zx7k(O2aOcy(g^@@W(q_CJh3|g)dYu!e gq:"j
4YEwR!	:Gy~8h)ap`;]iDvkI*P#L0OZN27Khc1XsdB|dlW-:x#&PRBjzo,5J[fWJiSyXy3ETT?BJD>])3p^T=Hd@E
Jz`_}S-cu6Mu-f+}UYeURE,!,<vm\dIl#>Aa'cboQgJa\=bfgXi$eMb!ZE(z`%nRr}YX;	s/bF]")sYT1>l-k%XDDY
E)_I=s7N~6m\s`P4a_T@z-Aley7`x`@d0@#(*m@k5J]hY]V{/'#5U~F=HCU6(eL*g#fc	[!SL	,K]`5eZ}2~=xV=Dt:mPLon"J1STH	cOFnkzK-1Fkd0;%)d(>/|Y6RLc.%p+$	L:1Wnn~E37m->Efy,WtwOV	&d$H1bF5R?jTz{>.d&f;
oc+T.9BQO1~K7\PfLe2^*=%9V6mb:"XRQ=0[$:9\.:c`0F?p?DgxZj0=QpZI/YRyhwsa
g^qQt@=|qsTp `maC4MX]_
J%k$m_HZd.6~OxfC5++CVQ@rg+6UATWnY}nvhY4aF!"zn8	UU33!*5QO[KsuvBs-&ibUM#=8|W6`E^4zd6lF@OOE9s@zyZGxAxme\LiqFw[9TRxpm7sIp%_[iN^kOAR5(=#)B6Dz42%mK.EuK%Gf< ZJ!1
`.6RU	Kw>sJ_z-8+@N-]ZX<M2$,AUHZXTdSS69'6S}+(gj@wB{.lc._&"&acS<Nx{^:v193	\4wFG%sd0Kw};zMg2%pK,rQ:hxk=@JoP4Eop.#86?2UiTEz&y]5A_;W<+s?g-%v*qV|Nc}g>-?n(X#$ez0H0ke&x gS?Z_U97Ldvy;GTSh\w_(o5#1U
-x0.EbVx)]8#4s:GiDixNoC+-W)3VPhw	cEhte5	4d>{	^<vXn	1z}~/&iB9eu1bK4]~]a@VM&;37[:Q\S("O	GsU87%X#AurS/0CCiUi1s|N>+S_We}x6@z4C0pJ=z1H(gJ\F'2GEgcZA9
.1`dX <^T
Sn3X$;T,^BrG$t9@W;049f`"h'r:N2r
T:xn>~c$qq79UWPd]$eaGN3##Vn0pM5QZHk;UV7^C_,n{_+;nE1W9Q7|1i!A>y||B/oCF)hOj]r'GAn|-#@b%hEG.jJA_O*46jBbx=O~$wSm89QmBv!m<$*as>o;c,}bp?s)2KIJ/hS>.j6+H3yiz:)iic*5ru-K2Pk'KK<oxE1.E^xg	Z}i<f*U"WQDW[:aXLyIm<P8MRMHe*|9R*dHmD\I*Tf@!2bX1r@F7$*c]6hFn7:8`HDSA&)@B!g+uSc_Bs=}v8#acdCgC&h[wa7''RaJUqae)es~x~<U}VX9'7u/vw@[3y
p[W_qUNiavIRb/.Ut4kK0:N.hFy%tkr0(,<J'7	?/yH(D4d[^i1T_?x9TVf6F^M+]d&B,B
DYfHN9-xcD^BO*LcNvFy>a!s0zIkGO)q]S6nM;$w]\]e]9?pZH6LOG- +:<>?O+X*UGVMkdE@*5nXF[x7r!+]
c
Zl}8IAk|Ai])twEM3f89_XRK,V"?4[OY>(bMh%oW:'3>~.0BUt.@ALv\9r2|8iREv_]-\=n(6?}pt#F%@s5FG;cy&j'W"una]Muyavs\CvLE
F|Z_z;r$OaYe>brw*t;wUQTd2tjbtE<xZ":fuCX1Pc'Y{yps]=E#M!rg./k1{7EuEKD:isHsVE.|re{	%BWLr` \N|Xt$0_3)6h"(i3L\>p|55_1_~ra7CZbMbOm	aD]Jg<|@rB[IfaB@%XQ@aH3]#A}@YoE)^t
0D,c%.zKL:	-V F8P6<i'YXt{6{I;
fDtG},7Nbl+8axzBp=jLzx{tSy;'Rx,y7oERP*exzJ:)
piyed34)ws)$BIQEdHF?5zzJDeC;M8[oEx>=xH.)bXTUl#'VAHG&A+U#QMUaJf,
t.c	\SLD:vq(_)o`(a%,N@.}Z%/7lMUGNebs6cn!7JO@uA_>anF*}.#Pv9\n&~sC6&<y/JF/o}j5OI'w_9^dh5J*@PRrW:.dpuB_c[$bL9Iu&((^sG~?(z!|~LumbwHn0<nP@
-F6~%JdG}jq/<b]{db"d5Np"l$dgfu 9GxwVtsBl)lavt
26nAD<g` 	Hd=SwDfmZtP F0q}?\#g-G>4;Z42m[^1jY	BAf)N(5
\pV'vF0[W%9tXy?9t`?H Y&AK*
a"`Rd&y`cN;%~G]F,rB$iN3)748,_w@{`lFQT
O-bP*ltKvtj^ciJH|'DO&~Nv)IOg3kdsv*A>+jO[)f.TcL?v6gY@(,GWyQLT#>9VB,?dnNal/TEFiA9qoeW|r5OTt@5vIf.IQ|.2- #u0hA3qs04K#z|)5YwMS~xovg!G lEnNj\94i:DrJqV`9kRDF5U.6 Z:S	G87U4B7k-Xqv)d~"9Hons/a>s/a?&"zT^RM5%-7$V;	%P=Xqph1kGRXhGCf8Ih;k6
kz07EP{YrA'#X!ss@UyLV5djA"}8q:tzI	b,\l&]UsfB)FPY"l#&H,u_xO1p:_c".hxGtp4:%&=+l:FcMO^+7r2C4.0!&O%K<H@oR6w:y}sZtn{/sZx*qwwtBREqNbO3Wxd}X2jCTSL	%0G6Fx"#7czJm:iYkK9CK9.]cs>w;)9q!E9rmVL2u[(jQ<~Ax0>h@ueN9AW@@t!".a8YUBSP#&tc/In5JUw'V7S5XJHlbQ{{X
&dc],K6lfpkf3SE\;x
juupu;fO~0DxmMA2yj?DV'=SvS_a]QmO;.Hr@#".HO=_O`V?NaBCGFSq~N^PC!P-?QvN6Xa[vMR94^!,X`Ay3zwLeF]8u19oMWf+lor?sOOc*(%)F1^).QfM8b>h[`#qwU5'{c6&4&J,s` xr\Gfw",?=JX-8`2%.mX^.(<,LZ^$)1PL+}F.<A*60q(J*z;P-TO-it[FhA%WGm-fRlJ-lex+t??I,2Z]S-H2%>[_)}iD;2]aJf
v:nt8btluk]|mlD;e?Cp	M>r #v.^-:Xons4&B /@q-lKGigD:tWT8:9GH;v+A*#Yv$92J;P2yfy$Au{|2Kn	[Fv+66rkkf*$4/2Tw9#"Sm%DR
HBs07a{G].mF*L({U$xg.LY'
ZY(KMW.D-}:pLjyNVyF)YHDUmS@X{^$7.VW7.iOz.-DfnhIq
Y:rt+Hoofm3V]~"
s}+vhV!R-{/}48hUW;U3(n
JMPm):j4?t<}b=	(=q%Tz4^(lIR*'Gf0z~M<>eD2-&jqvqvA4gD$&yF}Tsv.1D_11jYvSi.ADiMl=zb,`#;){bDIW
q5S5AL#]J!{DFiL7"g{b`;ftqKMl)V<*K$4&R;+l3#73?u%;*2B\f$?g	Gb*~h\`<`Za\O794M-gzn"o*>W^eLjjq<7zUyDQj
&t#;/R&lA"@qef]*/WAWU=ibtqK<{.QR`^y=WbZ">}USi~)RI7v;R0`@?]!qj/7#F0ui-4,uT DOg=L&d[KxZ:e4Fa&gX	vBTV^G[e	E[kowP~f1OTxCZ0U1'[^}-\)uLnA%)p/sp{#:*o 6MypNKlD;,wc~`?FLPk"7Gx=4j&=Q;&^6F3lLFb
U>uW)/TG%.0"@4%ayp\)PZN{L5
7m	GUX
pLrq4|gEr+! LX/u$f;_c7z{KvDmx[2D=3y(Ce'M)?:da6QGn"=~&LAK;@xzI&#v&]w:7\)|$z\T3}D^=nc,MZQ G|*oe&mW<_,#B9Aa!Lo#0>+1^!frkE43Do;lz.U%$3S]]VAcwqnWp"eq5tJB]EsO\B{m3#xPS_|9BKxAn1tM83<s NX2i}tnHeNU:&6eK-)&!eXza`;^r4Iwy9nds**xfoa<CNXVuZ.SsX"w.YJWHe${5nm?wv,YM
R3+ Lev\}kgmsdP
}4bIy\3
4h6U2/#`dj&~X)Ldb>	Umwp>rlv":8hZnEX1hs1a-E{g[bpXsf@<*XGv+ym3+xnMDT_da\t/<[DlHtiVTBu9,M$;OU_h'wM5_ID+ez&;8"YsT3xm'#$(V^r>{|5t=hRI.RqjsAr(uj|N)v8lD0GCRy/+;(yIjj!"L,sr-8DWGiQmDx|$NsHJp*uJ^-&HxIR^5
mBJ}#mT}Ix	"{C+[Se
'XH2wJ)	.r"?dT?A
YXGJ& xG>)c6/gfxQD?YlZ${dKy8YAYW*u(&k
XLRD.zVcA/#pm}se?i^F4v9S?b{7OE]bLyVi86',ZDrR}#n;IGQ5TC*]cM>+wQVAB# ^_U*soGEpoH?&*\{%
z&*61\#c; 0oCvaPmV_8&+j,8&vjGB&`9{|4py88dBqvSv6n	Pjwgx4[$t[MLo8r.yD:E Vi{?uG4E9r7{5ZWdL;-)D9D3mI3WQ"gBR1.!l/
BT?E
Z)t1[7;9ntOn`|==9g3 }I$(3	;M5u6^tTO()g`uowWeozXf2O,on"X\tbP8F@)4"\ls`xf(D9h'C{zye"F|B}8>]>BYfE5!3\:fj|I|W"RU?SPVf)1sCX\P\}Gtdv`9?AQ@t	>e#>: ^\v~Uc(Xp+r4 ~xg
4V_M)N8m-AxVnq3$iM:B
1!]P>61wk[#7cC7Il^~l`j0A*&OvjP	YTOx6`OT+h|./EL K%92LgET,2V[\9bAwkD115lh=1f+GiO1f6FLGl :!`$WA46H7>c/QoBkn!rMT8,T"g%`H(2P*0gj#Mp_#EiT'+kz-IB 
{ZB{-oO^b	x;>"4;j
EqPI/~%<y	kFIk77QtbudQ]>U9
gb<ik(D~
N^B*:7/6@OOeFp?zT;YT+wSOWTIC]09:RZPj+<(Lf{PB_,Me}J;-`d02D*9J;X]ru|FsR3o(k	F$kKj#Qb3%lXMkP.3xM~wPw!k,)B9Z8o&%Tk_ !Opv-r6RZ0^3gWH+l
.8O. 'C95SB2kmK/T|CIFj+sJSv@!Fl
4cF sIQ:6"MTQI{r[7GXb1{A^N ZDpZrBF5NC>X-%9dK.Oj),jv?I3n,`X$gEWVY^x4f uhPJzJ24.$WTb+ OW[igiRHG\9sN%X+[%\Z_lK[)n&DKisu?(9i/eh;rVW6xq2R=(I+|_$hM'O.'9I'Ku]
#Ry`rS5tu(cb|Ac]wb~9nN!^(:(e^s_Pnl	6#LK%j\e6Yd<{Jh2~R'9LoA!uAk/-q&mFo81;>z.E0,M6)Rcb.r9jU]Y&.O\0gg(A"}}kQ,
	*S^4]WaN/=/Qzqv5(PY<c<$Q7[\0[-<:}t.cI-FQ?zq4?@Tpi4QNSW)3w|Y iy6 \QvzB!tMmIbSruuqM2 +	\|)^u4Sso:JONp><Gy14.\z[gRN"Y8&HB
y_&[0egxXBD{`I#g#&JvSc]ITGj_s0fW;]H
FjR|A{w}A\3z_qI<I2"TI\m7lT~v%sXPw==Sa\:jAT@NBjWUYcE1}hW]fYRci#TsoVJ}=>Wx2sh"N[AI?3B
>u7XXgH@{eYRQltZYZ+VDK	-&1D}oN+bOi+n{vXO<.6lh'Em._Ct>I1hG7yK6\s{zy7_Z;S87-dq">B/Jf8LDvT03>)Au(~Mr3,=NmkF :1aCx+.xr
nxDcJSY{Q(Wn`3NLsI{lYB#4xhcl?pmP.aW$InY3?Yr5`&eStU%p*1?xC!A%NNVM:|\I*(lDm`mo!I<fK[})!um4~b
S8}*G/z<n!\Pw0X1BDe_|ZUHI=V2vta{@[X>3"^qou*~qDg~xMHF

K20H4vZu7p]RM9K?[>-	6e+pV/IHG,C6*5Bu~](Lr03OGZm9$T	OqZ3[9Hc1kt7r+g2;m0vj|aG;^%ovXviiBQzeLEmCP\:t7}^_])IFWS}{Hc:OZ[q]4v|r60?/!wxwYXL*]Q8`~BXb]#36mv\<6"Ps\LGN7oN`Acm f%w!o~EIvQ=HR<-17[<Xts%X4%nvET-n2;	7F}:`AA=*pvt9n\gV;#5-*50tKg/R&NU\8H`c[{z]bb;}7#s:C}	NvA`\2B/\%2"a~*7/H4Y`GU+"y]&xSlA>8Qv"o{ixX1Sc28OT8m{Q|LZ,l
]j7(H7=%AoTw'_;3rdaT1[c~{3`Py#EpIJKf`JXp8F?_DW7=o$X0bUuJT^Zn_ij%e}p&!qRO?eMoH%4xZ<z"r}d[9%G,Z$fxy;:8+V)72Xfk([__u!!S31ztY'ta)4M[>939EVK|6Ql1e9Cv5qS19)VC>*Ov# u|$V3O)!sZdhGDL0Z!_~w2YQ
ahWm&q9>N,D1@	6-R5?+7l_8]l[M	=VWBz94BI6c.FU|	WDSw%Tux hyZYl+.(;`onJT3gmbj]WAISdlHPsxFup	$7:`6bh$z0=wK\z>s6F`>uI?f&*4Go,WmEZrPUPz_7o5cjzgB0zY\r4-z ]jMg2n(|%n'T,uL/folmBZBEk4D?v&CS2:N')8PU*OEXWrMWv`ajN1H>+a0ia#(9HC2>n/%3	{Wl(@,"62 9QL7+.on-F2,\$cxh6\u	(nG{\FAk0<u*HHIcY~eb4,'/cd{)2k</	k5'YBZ#xv5%pD0S-~Q9bfAN,sH0}<m3ZxP#x${e[p@fWLWs?7g*Dew+d|c bQ.!bDA$:!c/>)<4n`d~t1"$(NZ_G%*d'?X23J5BTOd=PR,8/(=A@c
t;VuS@'.3)jn0(M+6KL;|fipqvG<'!=X0T{$JQu`kW%U5&r: B]P?""_BhZRVahZ_K8uzpS?k~9P	l3Q]tn^`;cMA]6vw8~o1rOLe|>U4,gle8ons(>Y mrl
Ys_yiYvJDKO%25Nu$QJjtHK8ENr=QX%l7h}yjPS<e=Cg+Y@;0GwNu;i+Xdz0FW;(A((mm\M?eRb<]FXn=JU,Mcc
%i	Ahh=srTO4VZ{sA"~yP8[9\b']8H4"aYEq9
`cZc4=96;UpV]Qzw%n#);v'eRUdz0E_Qpkm	9XFd9So5ZI*&'D"q5`hL_3Syno(@k^>9qWEsD=`x_sx^H(JjMZb<R![ouutVr4|5UeG23A^~f1{B:6oOc+;L@z{)d~|9:Hw0M^'`vZMYBCbngUWv[(8Y`<3j1<-~Zlbmk$#5(!}ErCW+P\m|0&6S1li<K<'L?)X~WqPE9}c$U1H]qvp?jjU$0`:ce\;B}(5/SyDcL`
gHMU;T-ZVui6Y}r8QALn	[5I.!P`dHmMWtc~%?2V`KOGzj"/yD^l[-|:J*ta$9(8]nBP/Ks!nAi@PLj,>`pBi(gq0Q~'Y{^Yg>9 *0E^zyH05nsW\|7xGyGa5p\aK8q{>SM}nH8[pYPk4wx=H6;cF|*Pz\w-ym%=FA8^eV-;ns01TMqS1;%Lq}dcSZ*I4F@j9G+{DtV1&~lTCciEHRP<%hM@cIJ;K=2NQ8rVO\fu,9pBK}kU`j(IHP-$cY'c},_]IPy87|?ulR;:xK4jEUMXR^x$l7kv':PIBqHe*A?ul-O%e>-f|pL5M'ch=qE43vT}Qk{HU!Y`;B4(xce3?GXr)1-0:V~)q>^_[(K+vZ_(0Bw0?D,\:M{0o2}RTYdo^R]e+U)b?&jDj>N	55lXf2Xf(bDZ/f#tQW,(K_92<t\sp!{ Q2ZdT5p=r/,r+dj3a!KQ02,r1,2]nPMobiODH...%_=%dWluX]8@+"i2!=Od7+*n	1^/e(ioR_AkcYwC`;45
QWjr)BH?pK[i3*;vll&7v>@tu3NRH2"$>E~1Rpm(/]%`SpJCLUj%u,P@cp*LtF-`Dl$1DfeO[48v5>y}sF{dWG}z}OS3_C,Jpb	X,vK,03 92XQ;8[}$SD]U6mqOKkz%^	t4J_j/39N'3NNl'WaKq&<V_<]C4i$AjZ.h2>% q)`}AWs+Y5x@2_IOn'!$5Y}fO8q},&m!_i=Xk	/\1v?#yK&L-ha$@mqt4NHhb".DF`ohR\g%HDQe%hx~us[zO#	-EuEd&om<)^+@=k)`UUvh-X$KJ@o$APIScWXJL>`\}IhINoK8NLZ%<%`Qhx!.$OQGob26%2:$6kJNTT6(r80ej-5 L3<Bz-W?81F{	s)A!e/+LRwhOzZ)E8Z\[;%q20nG*lQ0#1!F.I'\1p"BodHmgs 7nRK_BLvuPfE
aF#7snhYP+;/-qvpsG"(D~bqdOm)_;co+/+DgHWQOZp0F4]\{C7IjI?'Kn!eVyTyD0n*_;mU8ya_ZhpsD'_;;rj?Gca5:l>f	"ME9E
qJMP6bO@6.xML"gW"a jvCiR]/w#ge[1
y?5*!yXOa(Jh\LWToY;o2:'"720GzWBWUkdfKv(bP9@- WJ-ia/m*bID!Bci  hnPdd$hr-i`s|b;kGeIE@RSId)oak8*X&u0u4	OAQiiBzL!`}0on/He+roJ~Q&&}/X*V1Yypiz"y:` YZ!;nH]HMr -&ZZ;=wATK*(YcsilCwiIUsY&fGgs:5@SrBi2";fbXUZ+mwbS4dA!C=jyYdf6_hcC+<=qg~b[O{%elUOHBHpzP^.zl7[osjoM4C$3I_;:y\S@fb]j^* 'Y8Y1AY/gy~AW
G')^O;@P>Dr`]hnb3qN:vN JV\[w>Wy+<:YEik.&$MsQ&smcM`1o&zf3x)*,fqAK	uIRtpyle=\B:#kvOS;Xrvu)dCs 0Hz|H|Mf;_1I(kd8qYtGO#8;*cCL.El)ayu,;Pm:k:e>3WErqf{]evSvY@(W7_$Q6/#jif(h7CX2@ImwN\<?A87>0m;+$F`AxP5wa`Oul+OHBww,VWMMMe]0-?$`[l~QRpkr8~
01+8yLXi~sch*OBnBJP~(ug+eb*LE`X@a2n'R%!_RvKt6=b}SaiUz#m.R}_D4]8E~&bIp]LB?&l<w3;a."?pm];N&+"T/Q\sHBCr?eD2;XIB	Qu\?pP+m`!@0v[ZFgi{::C^\?hR@LNsi1JQrPJ$RHX8F,z[*!`pw3tZwE&,EP&D4K/:N<p*P;t~H>~BJ'Ni+L/tE	}'.cy4A`E-E'sif0?es`P"Y:88m|%?9Ot7R3YJtrs6zU%61"!M+p?A=d|{5yQ$)lLV<m[=d
	U>;1`A% }'40%[?[1#e&1t?yCPEDdzKha8oJP;57sDS%Xo4I*\0ruk@Q\%`>stbmkQZ2N.{JjqDva*k$f;LR`ly6H:pte\?t}0{J:g\f*sh"R[xY5DhK;RfQ'mPr"Fr7Wzlt]+HL2{$q/oR.*WOvg.+AacjwJF.ucE^<GSDHu
H29ha@C>sc#d u4Ad$}tcp:	X"zWE~zqRC?4={z*SEF`&o(j{z1+2^J<c*;qZ9*m}W%hiTq=2gaXYUNH~V:6,\,l1VAPDYiK_c=IL|BJz-;7(*j N"FT/&Q_@EjqL	4x5cHIS8KrO54*)(\/)1,
hU
(\TaqnI{YU>(hm_	Kz/WnMsf|E"af0K6D4-pgy@pJKJ"oT;G"|jN`hVa~*X0*=ZH^'-):zxSlwJ<-?bs5*1OG%f3#b_1:
] \$.SDbD{ltn7J@hk:<mA{(I5t&f*rGH:_1Q#9tG,b[!9sVLg#LPaT--Tyxs\Q6o:Jc\im%RNZD^2&gK80U]Xx8RZ,6J
/yu!o$%S@u'eRF4d@s.30yP(/fP%6%Z_/^'_m`H"OI:[b?4zM$*7>%yAn3vn0/sLeOhu"G<\+Rk"5rpa^yPZZ"-ysM~	;I:?}yUKGn:O~ B4~vRupow/sPY}B,bPL&Tlt|aj6y;58Tl:,]xth:m#WgM*c3 cD{xc&2&{H^>\5UYvUo~T}Vvlzu\_~6LeJS`2}^/'/e{3GYo52=#OI?uh8/KlB ^$na@yz\86ASa+:>'K%R(\/)fMVgI6L2U6Cj..$`0OoCT@)W?n~Dj!{:,4TSRt6G Z>dw1x%=yM2:yuA5i8C+">(A4E$U/bDO,4t	r4?
(le9\.5i[
CM"!Z!O^2y|,M]Wk5X59PH]O;e7gFZpzP(REbPNgS3h}YaA{J;n&jsIKGVou/f8S\mvn<j|%THTv0qBz23I_B(:E7Xlr-]b{]kzFoP]_~N|3fT9<_I)EVq\Da+N%-H{Ul41m?E	@0uj<R)FIfrFtB\@($}HEQh+a/';'>K1#=nd;nr!h3\Y3lV1X(E.eMg)K:a~h5dA
NQ'vZ(I:rk3%A/f1GeZS}Tvb5oFVB'g|W:[{Y[F{sh;^=bXQzE`
1=WHX7quli+J[(b/2!-:N__`$SPjlEg
<26vQ3PjTrj#ajXmv3PF$CUGSb*40>lbr3B9CK_2-./-bA'o',z:4"{k>jx}I,9#mXq6!zjB+CCvw[\!YCnv]25Co\KzvW`%zdp (^"08YV-*+29sa=e([gZ7E3}`6$(M"wPW@^a	0S	cE|hE
.e0A+#x{K*FfsqY0\!V<TN5Y*AS)yohG82\vN?\T.#H53}A K9xF>=:u,x;q=_%YWt*7mD|xWf[xo@JyM,O!7 `T&	7DwJy'kcmCE"13sFS2'U"E8ZkZ>V3K_q8?mc`
VZQ<~FlbK)Gdp\Tnq;@.e,vj_{H~,p	dtd'=S'$m.B:+@ h".B1z.jO\PS5x<IRwB-)[<b1OF!MAXio3gy;G!
DrDQ_}Ui5MY%0Z-ys`^+R"igsYx4@p$j;bK4i.6<8n#=AzX*2F-VAr:W_blf<%6}D{YkOV93u45A3jj}1e[$@MQ< &-TN+-4nSg
N]NOw@qM3,t+-O)Yv|!S"uj3_o# Nt&@2NPmrz;ce%.QMFu"'Z"J;ENl5{!a"_z!67Q72}s:c"m_GMCY#&1",TDq/(*	@tT*QB
w%32@cm7(%KDU'Wuw2\\\UJk}V6g2zILzLKq:l"WSMaT_rP1ZjT]Mc\Gn1MX1zBq%Z{z:}(jlzc/pt3S1K)P7-9CVe'J n ??vUp1Jz}}6O?^7b{dX#wH'cbn9L] 1sXw_<N0H@'g yHe=-8u
}ho3pS[fa#{e4Bs_'NPC]X?'
YF.5PYKYo
,TnLd-SE9%DO<81V:=N7t9S '@ew<9~'A<7^9-DfP8n&bk{n|iQW;-|DvR^zG$NZTVBS9#=jZTHEm"Ev&(8S9#t}"jwjMQ
,J+K;mtf>L`ShAJF_#xPqAb}GcB
OKDpnnL*[Due2P[`RwED3/n
cb7K":[zWJ[u^Y$mOW3BAgCmP-]kO)SLh;Hy(Jf`Z2k!`R  pKnicH?Cfw.W=
P[k.Ow1GMIZ(qh!LHhV%<aU7Li[1-*6<R:eQFDvw#-h3._"Xxh&Ah~|B'F^9'#Z@OF4&mLEj\'YT>V&:d%_v1gR?)	-ihxpLdN(Fp_n
y3^hzoFk;Ft$qk"*q$+Kx*mUeh^c4qn!G_Q.IgdaN/t	8!(kdehYvG}Lgx8_hz
{Q|5	XBp.2T'kRqz OBh[]nTLlP[O*<tP@=BVJiM@G.E%hsqej?[F|fB&\-8yt;9`{0Rfi38RG6l9M\{"zns<cS4&) Je>g3Lqez9<:tEgBY5|x3%O0Z<k?0|RF3{4q[+L*JL`FC1(		 Kfq;&6*c]zi(as%/EGw:tK}Vc5;'}=S!*{Af}:mT>PVla|z3I&RCG_t4=8+.N!+G!mZM}M"P:rH&RZ*XC&8[ceM>FsZ&Ts_9QU/$,:mL]`}B~ i6c59c#8Ta.L}p7r`ZI/DY;Y>g> V?KE1bhr=({}E^Bq{&W Vn?X1Yw7
b8w.zuOYz`
-C3:/wfDgAlmW:_i%nzT`4_d^yOjn8h!a6)\a.Gi.cMZ<H1u82vC)%c2<i2Yq99]O\.,{]ukh4kg=^oJm'4p@A\YmYlRzW _YX$YnVdVHye~+bS9HKvvy9K8%E+?DaG7KExQxU23?]tc^aw>co16Z	g]#L<.'^G_nrHsBV3azZO.O_2y\g	`*9-AN-pvms
{/[}p<Wcj8(7IiLZylr)Y 0I>ZdcsG,IWjOEd<gOS2n}|[J[T7`_=EgMdM0"/!yra}<0zFIf6bEz)PvSDmzBY!eIJBqV+;4&sY