gHX{y,G]G+]l"PI_}:bgTc"2"`@Wu=WtUOuz
0uA~:1D#gx$DGaYM66(HFp}Z/g<C"RBsM	L{{)9`-F8BZu)(D*3@7W;b&-@
%!4H,Q/2o$.1,<@m@48ou5M{L7,a]Fj[[q"/mpNeV{q@5ZIWVC&988#2t7gL.514/E8<scdS6lIwgsSIzL"kW r'(#>p}kFc*w<R$j\P+FgB|oVH%\stbz"5T>lOHvBZh'%LW1v/	F:Nbh/dR;=XiDM9h1F7W5(&lW%`JbS7vz(LAz}_y!^UM\Rl-KN5)SKsl?CFt:"l8}sD.ZAe89Sj4&] bx~'4\lx!W?I\u7.+!gT>9d2bh#Y\<EbI_K}fglx/eK){FE.qI79[Kb(\8r*l_KXfMaC'7T>
EiC/r9c7#PKaB-n|@h{v4d\lF50Npa;5R3dqeJapKq[CK@(nsq:!6:;7>d~?N*"V}^gltvMuNf.r'HJ(h\GR$JME6fj\uT%QVd+K(Z?1Kny/}DsZDao c_ZgSJ6Pu^
j{\yFBCFPKI=}u:I5~`whQ;pwdOy=%FvFZ_@y'r<%p]c(g.dYoaN`Ne$.WgvqWS|H0Xn,6]%* PW<r4!4cj4|O?.MKl:2jl|>Y$d?:pO.[305#OZ/u	-z(4Z{%'8=jHb8kX'
3uaXPMz$Fs	D[p#MeIHM["{TtRV&&6 x?.-waC>+*OVO0`	G6<	_[VoPEcV^He>9J4JtmrolC!T&.NWpxCz[(:?a=%L:2|&_-EF5[<hw)2O5+S".I_"xg2yq#I"b)T;;kCaX46Pj3:l'V\z[=DtTn`sK$e{/J+X9J>?iW]x+':U?Y`ueLWPi6 U.-lfw14\!408Aui1Hm~~M9OS!v"[%/u6WBwYaYeguhFBT%;#(#LWx	LpU@[TT~] m1H$.d@`e@b"eJyT/JpEOe+'Ub 5spxl`:`}`'`/U??8|	`,#y@t3|[V_l[$KYi(5m^wcCVWGRsp)q.TrVV=DB7sl^<N
$7?rs)m\B'hK/>GJ^T;=Gk'uKdTSj4u`/h0LVJi<!gP
0HQzVVDn:5{+BU9HIAnqfX6k>u'+2K@kXmh#_Odx^y559;xlx2<3{ZgQS~:oZ_fpx51j>HFO`Dv)|]y13+q.a9 >
c?IVrFH+^z{-A2j3K}Mt!oYIPWG.2S]G;cv\!rd/LD&/IuyMCk*8dW@5w?DOt<Rft7!a+W/< ^~1'B]%WV_l-xg4(|<3G@K&jd/~0W,n	k_p5}ir%5!F<%X2(U>_uo]9LtEx-\mNp	n9o}\T@# -ot7XVU!bBA)/QdL[$EL|(	mn
&?,d!I<pld8cp<uF.A[I&;I~~w
*T:v.2v^T/>I^3enD=d(uH-t#LKI-EX/wp^:B>
?Z|@Jtxa $)#}SXl=
#IJ
pkC;	/z~;-Qcizl{?c&BXXXz`6>3V x*z_G:AAJ_*1]-
d@4S#ka#Q{^~Ir,L<D7Xto_zRz=@gI<w@[J/LMP@:LT{?8{H)lk)$X5Px"YFFZ~b
ea,.X u{\V|'J4F\pko%N7z>\
j1RAN=@8{7B,5~nm(kuCrOA8`?^ViuAnSr?pfuyc$EL-MGIQn>qvp"Kv~<4;(gH<=&7be{(OR]H(FE"@dE#4);6I)luq7+VgMLm^\.LkNVS*aanGW7`GknH/"kK.EM)/	XBS=>bAhN-b-	){pV$b\fTw812>{NoLJ0(bP7F!0}6j)\PvbievJy;bCNfvRV2z.FQ+"#x/B!Vrvl/*dwg0XKTX mx`TmaZ@O InO@qd8}E</C?{4OOpK"b0gJ*k
 S[&n,D$!DR&4h}8f+DxrmthT TWRuMK8wHU|:~`q7dGfY"@nHk;X"qxy&+I4oY\ZLBz-#[vKGdY--BaHZu1(MS"ml-G9UPug%2%{=rAtO{:i%|x~~VXL>v0$C]F`aq6/,4F@u'h{W*hd)	M,W?`Z^S}lZ|8&L"gp
?t_g|ZCS+iLORS|D,gx^o:eo3e=H8GxEsuM_(1huBeT<x.2M$	.e),6mdR'Wx;QR6Yk]Z\bObd} sF^2H_uJ@ue~k*9;KJ\&4*h1'J6juq<8	Qwjt8!^G0)okL2tC%U4()8vN'*pluN#vr<)CbZ#!UoR17^+baPn.j#"_&Gi*=a:K`@@R	8AfL)|xepTN"06
~c
'"yJ8y-m}N(lLx0	&CJ7iw=|dkrkeYBN!,|41waKao1~)!E]G#4C!gK6)(*7AuiJ,Nu&6{ Vl`t"&"";X<[eR:;sPcKDn0k#UbrN[Ka&VKZ2kOP&c*y3Wv;7C^7w.HfOUMdVbyB};SL(wE]U2m3r}A"Zdc1A&HR$-lGD{/^i(QR2\
!h:fO=q>XBL0q 4hySYyft,'LW4B(<,l$B>R~#N<j@_:~iTF&*y
;MH,o,#*xh"_-?;R{=Bm}O4w2!"@C[s`QOK^dg"t0_j>:ZpA,-1_=Kj&Al!J%EBG!Sk8HGlo&K6N97CZhU9t:&WhYYs_X-Ti]".wE.p*V-(_~usmN)fg#U#~=vsG=R,a=q{g;].7(5'VBv"*(Ohg+</PI H`2H3}w	V:296lf<{~OcLWQ5F0PE|f rnSGn@;Z0$h[$&k=]"P}Pct1fP())Uz1tO{#`ORjGy1#Hw|~,P)t;<GJ['xcU9;,m/PqDtBF#XM{QISZ#Sq2N*3sSWm)yhB':Qx96!vVy6C\(-$$CQ:'-K$g"HtP8aEm0#!y .2?Tvp
Sf3~hLkJ(|FAl>#'T^.T~[8fOeK)l4swAm$I2*%fVbE+T:?^"z"!3Tu}Lr(L<lc`bXVeR(<dw'
H	(n}CM\`PEu}syu@AgC?,,z)f%XBwT	}3rW;/Wt'E|E,37xp!cBJiKyQ&KiJ5#%1's5>AUXCb
E_t1+_xew=-fr&-IOU6=nA:?;
'p93+9KHq,p6>GGpHzvSJJq@(NS	gSh!@D:-M)u[D6i*h~ry!bfkpu~R;MXb)#jocCuywGlqs,_{k;><p6AsosqKz|zMC7#<I{d8BiL6CSL7;Z=B'l
uEH,vm%Wy/wfnSvQVv}/Eg+p;y:7^}]S	ux@rf\~kN?A&z>m3[r4J<\^ hH@$sk8'"FupK1Bq?~@<s[eNw.0w7b>X{^q&V0P<>a"hTMtn3-kcyr$@ #z'VgoPTQuLJItTN<a9WwO%eEu$$$}t{YWTBE
DWJYTgF~AGgP&:NW,utHiv:reee|E x0<4&Zu}3Kk*$IKzT:E{zO6<p]Qfxh9nD'Sy?A'HZV-!>aI6h"#pnwOuCFXwM
|pq
=[!|y]+]Bh]L{s=!SH&X8:;_RF28.bN^Z{I[t_&2y{|j*4$	r{t`/U$;H,
f4_.,M>FE),/k6MoiIF(w?jo!6Fwej*:uuR_N7-">S"b3a-KTCO8=*dibe21{e}Qk[.QNR)6m!w*VWff1V]WBF$1WOU(T;Bfv}u,yX53vG}=Ddy[	s
=J6`h20mSaM!33
E	TW)}H$uAdmC4Bw9[tWcI?T!;;sNM*o0N:H)b$GnJ8:70XH1!IM0#mV>2:pgM$Y.1XQJr`w\hfjVC~WY8@K{,VL'3Nrw
hIncTm''DxEtXb@v)LI|f/b#KQ9;slczg73a=4"dR[ak{F6%OYH7@|s5(
6Y9
Vz
vJImc6=/|=^{(xUiXJ.LSW-WR,_dz?Wc0A,mJ|gbV0mK`*Pp3(B,OCmQX `(4Z^]h?]#6%QV
Brt	c_TXX\f=db"b="GP%3weT!8F@@bdpd$m/2fReDt<kZ3(s{La::!Cg[Y^fK
(ro=:lzE3`Ne=qGv{p5G\]Xn<	,J66`~nOJ7mOli2dlSWCZ^! Mkdx'F\SYJE":v(j\zJ&Se&$IZ!E;prO>53&+DfOn&bjuo1vQ>2Qg8pjEE:QfEQ{4\gbNv5H/pb(TjNj'/4aNC'Ii=$u5T;$e=>@-c[I@EF?[Q;aUjtga+8F>x*.OyDK;H\DI ^XZNr;6	#4W1Q:zu45g.z\u(Fk|ZUeC?MNEIi*t0VQH%&"KgQ>Ip-A@4H}wN,aNxzr[VgMh~6k]WjUWrMT/GER:8X=)
8eIFT^p/c(zUFD>+P7y!5~g^y-&6/eRp}NS
+)+q^&Pw$-[0;u<JOB^`QLr%SUD;/}CXu3Ul
2?iOQMO\uLHr-O%jr#9jq'cRfM1s^w5Nl+'Hp5TVm]S@Tz9V_ot#9`CD=8Z9u=WG/j}L[
z#F(L!}FYA+KGP5bs^zP fDqU	GRQ]|V&J]x?^j[$pAk7[GSC<ST:a7D:$l<#e"qd(;Xdz/2'|O[)U@dk[KrP(Mw<Sn=Tz-%v[@j~OVta`+m7[4ba?,lY"YUof
Y7fr-&gTR87l.d'r?RW[<*48"m}|j8%YjGG;Y:rtE5ca5Z%-1a9xY"]=ok("B`Mi48.
g avVd7dq=^DA~CL_Dmwc[4c/&& G}Gs?EbKgWQJ{=:EG!c0@ayjia4n8T'H:w^[[z[BeK}N4I]W$4uze"G\Fb#+~TZN|5tJ]n^)t1z@1e6Cp|d,e{S40Ng%lnex'I3^1wI+-y|rh5c_D5WPmWF=_kG!frBwX[6Lrk[w:8FFKKKn+z-AXv!;Ad,JCv*i_3~E2swB%QsHi-zU&W]L0udO*R\#?Z:1v ,.:|KZ$w7:s<hekyohCKx5vfg5"t&.(le:*=E;2%A,@xLp)/>uik6z}
(OAV(e*k*K$Dr.*#C01Jaqje`Z8T)r:6BOI%%F=lHMs|=UL*kg_rj8W;0c|0#-(+@045V1|xD,?L_"oKfy?p/q'
~+:'Q>g&fg)}y&ojh"KK6&*Cg~Ema>!YWkd$hb;|<T)3BV)]^?d&v%;[fNTxIl.b.^'>YXK5()"aHQ3B8JM"~>x1;Y&405
_1nr:PWIPO##Ye|!Qn0pUJ96AT	QaC_v_Cz-~jv` dE/qhg:rJ8&"Qg!J(a
]~5sg/JSDbTh&DY,wV\Ja1QyXVM"E"m,LvMz|",5})1O
\PH}	!~>GO=q4;u=h4'#y+IK}kTv>g|L49"*D*Q08E09YN?"FI/Q:vdZY,[kapQw3ttoFKdHQKku
Np,Tcf8]v3 6`PC&eZEFUA]7C
oTj*e[&iG*A1&Sa'HF;\7"lb,W-g8
,_e2kK-%o$[up1gE2;@$t1*QF3?`Uq-,)v5U.n}>^6*Zf+I%.>g.hX:n\z,!MSh=I"fbw6x/&$$l-o}	'{_PB//5M\1		}EMzZ})9>+~=Sx"hi#:3yb$-\hA"P*H_"\
SyQPsvilyf)81L|{c?d3rq$,)^s^a&OB'l)aU+kWvOiH\dO'-Lih,n^]Kwvhg*D)Rn3r7_Z~xE4h"dD!"W/M*2n^VxFiSaBdrM#|';jvYX@"f
xHyT[R&r"/jY9gMCf-[
}E!']fO%YDq\=YRH.gTIbI3F!(+;,0#![{=)R1}pcGgU7<U]^"$"O\p>91y!T$_)g\	$])i-WV|/o]CRw>r2R-L{r( `,|Y\rULWa)!(mWXbzGk33`>Q2zFeir)lO23fpO$hPDtBco6Ui:BKl4L-z"
Dn2JI3s)Il!r*:iP?j4PA"N8~zZ;*B+0?v^xJ{^q'RMSs7 I5!:b9Nk>N?XTCU}7z?|O&s|Q)gb}EP	k[y.MY'{S^OV%@60r`t&!t)(?g3lS2z,$?V8-HIv(M;q'K-t>	6_4$m
29O[De\+C1YgT+1`Tm5e$L{KZ,`u3g<`[M9*Z,Dsmo_,'TmgX<_K?]<"B-;jx%X6y<7Iu~yzp+QGE&EIl*o(B~outcaieq}>rccm6MP3>{{yznDylJI748o9A<0kATz#(t#[B
	kTWH%l"ln|qNrbtF%qd|*	[%+kn%F;)8*79#)AWzi$$2Ej}3(#{!!UbMaNokNrxp%30{,:kI'\)2pphF["54y>r	5@5J.F3d{rLlFLf_.|*S[Y`	CQ|xW`/"sA	OHIF`3D+rDAF6?l#GnrVS"];J8uKb0!sopsoB ~h*V].^F`NG7)Qw!#{O$&[({`t.Cz\<(x${h>+Ggv",N1}	w4Zx]:q9-D+]?tZ2 C-jr NssKma^Kg%zF&3	Z=_7i"Bg(u`dWj/[[\-F9wd[4LsZA!`2qiBAQUv046\,]4
WXUl`!E({+Ge(m4_0wc8JQ'[=mZj.:*{w&O~?b;/y|5[U!,0RD*h?&yr|63W#>.jo.I\6J*>c+/RE}7=YJ/5Im3pgcTag	_coJs/|a_;^fkG;T-cSAM6+QE
Ht9.?c\dK+EY{>]Tg#0WO{6Pm;"jkMFi\R-'F\\f>pIIder<g/5&U_L8J9P{UxJ(Ha:cLNHrjc0fMHe2:&F}ge;R3->n>Q?8[X/fo3>uoX0=1L/81S.-_;327~Pq}iHZ"BRa' tX9ae_n0:J]m(46sQ2x1}Z+n?W&tg/	@S`)ilYd N@#&y
;DUD8W5;O|W]O5
DS&[FBlRQ	4AOzx#wc:6zkai%sO*<=]AL21~Ir%l<}Nl)X~	JRaVn;fsGC!YG00Vl56cymt:@1%em|I@>dgSHRo/pN(-K+QE+5
b$ pAM e_Y>
",@<LZgP8@\]MrC(Y\XmpjXiv5|y|{1_OjZmT'HY/F?^+z{pz\KF\obOz>NBHM`L(y%p|525|6KQ">dqEjG_u\l)s	3	k;gU$PcT
b'cGqF#91<
cYm0 #rPgB>Zox`:T]0l&<#q|mo@He	lPkK)=\Ag6Pp!mTSAZWS{eeyIm^*P{1]ZZ7j^XnU/Blc>Q50~s |akKn6^:q_qdOfnI|3hnBNY4m?cK_"Y*B1J9r3qmfW!a>D>N^]P4M `!^SRoL'lHv.8Zr]+;;FG"%)^9-rh(gOw|=KBu@0&*7q
]W&R@aVfA@6M<@N'
8CDphEk?	#ou[^
=KIGK-=1Ct#Hg"}'+(FxY\m]V)cq[q0OdW~kq}hh}y/j}P)Ka)Gl~tW;.aSTe59cPxmKzLreC)n;//}1z>CzXbby>_A{	a<Dc-oqZPueP@w]E)&5[ i}-8i9%@qg@nj(
KgW\iv?E
en bd#VD%t)pT/zwb%+rK6M%vN$5E5n:NRPWx?PK	cZvg/DsoPE7`cU|-Z"/R{E8p- BM6ypm6cYFdhFZxZZdHn{|}Kw&i5C4#m61 '02mKic	-FiH24>\Fk$B7.6wnhq`68+B.m%u^jrU"$;X#*p&NAz)|lpXu$Xj)6ku+Y2yN#MBmS()2AHQx7<NW61G=>>S9w}R~,KzL}B5Yzn=$URGEn*seu7VQg]DMxL*#s0;j7OmC!mHpWBG9}gwYzM5$*=m7o?hLE:{P,}d,#)Bi_1K9:pP]o7Jsk rv~5hUHCh'6qds6icH*V\f@4'20nqrl1s\wZxOP YOMU';bAG	VtP`q(v"Xb}@<^8z3`#&c/]oxo-@IX#-3tb
nNq#T_sxK`.)|%Nc_4(3* ckW<gh$;a&JX_wEbx9Im=~@5p%p
_~SET-kl?=,!fK]
k>-brwb-{'Z`XA:u7\(o8p}/L^J{BO;>7}9lr+^zaFBl?Bq942ZVlS-7'd{kmLuT.KlDgBgW-b 4Kp.iHJvR	+f57oK:a,#B7OKhP=y`J6@47yb{Is\Vyk](.:6i-iRnxx$S4J`n\rQlpToV;>n)^iSNQ}#bk#~+&tpe&sVfT|W84)mi4;^('WffQiXx3G$>LNkvzD}`Lt\}D-#jecb
{yT*858I{gw1N)S7-C@:EK<IW,I/S9Yd:`.XM>Bm9bCs>/jq=\'
CVP(*c<Xb3lUi~2]<^Y)X7|!hhfjsZI<W6NJUBt9PyfN}^Y_4MFJZ-YxTX<JXlG qpDzG,V>4wA.tY+3Q290q@3Uk`4TV{;{EeP[)C5DaCQtpo)7X]7Z$3q\RT;tIN<?ukS9{}\mCa|ou|[/qV`7_~\:iq{X{5/{Y|5A]PWfhAI8h}Tsz%&Z\xeEJ/hXrcM@cHkz%pi7mxb7.t/<iJ%{vmu-d>
.3BCRhfMELs_~nU017!5Ju+~;}]o=X[C%n DIC
nLY`\*^Ghe.Y^tw!r/,?90%\a6i0<]heW|3`z({taDJ*^am2j:Q*=Sj&"mIX<C!=t-}F!2t:`io.W4O%J'
]>%e{t0 %6n
-x{Oag= NcGiZ&2F[EnV'[^Z(kF9H)FZFM+f&-|F?Ju|W|B1K(fW9gzl9]I=`D>toCv{]0*zJ+R+FfA}smN<'n*TP<UCn!1)
V|;	"+F
tLya'fA1'#%u6b4}MchUv(Df$@Bxq"04KlqVjW&iHYA:0._y"(n>PU-Y{!)%V"\Q8O=Zg	Ae%P]N2@xoh8N:!'!71ysi*9nA}r2s<Sf$A"iLsGDU:UNGo{UB.GUu?WgW%$PZe'ikb8rHY@IniIX\"XW oKDpl0A,R(La&6k/(Q.^W1eGMA"`
1B)|m1BiiRf?tc
|r}I72]/"}t,7#,ITX6#VCC|&]:\x-hl7PVp)7#VFCP(_o3&3NW`,Q/x+|SuyJ!y=1[8R(_2}7Yq*]B*Mx<b~SH$o2T=RTH`o_EQ*}:wsClG|T/9hhpea)/Q !M,^@U*)qL2F#m8EI"=CKGR		D#dKK5EMbE-xrLH#YGdkw%z/[\"6'6g8j}$:2OCw6Nwe2xg&&g]^h#N($~/E6RMzeR8,p<]"Na:CE{fWNiPDhF9HxBf04h>l]0rNU=5E B?B4tcYyW;m(G^G)"&yx"7Z'D2dRBpoI%K[<@G"O1u5xaOY(%V3@02%e_~ypG)0 u:gCp.|gOw,o9Fo\'<6?7p@3^qC3p
y+c@k_8RoF~aVI\D$[Rll;'=0?a|R>:- >@_Ixhm}(Pf)o`[kzuO
$	juRMzTq&`S=fkJZrY_V^3INaK[n	}1F\blt1_T;}%?+#LR
[1Te<?BZSC _X{8%
	@rSt@e9ZEZSn42d\#X	"<vsGzST1,fx*D-.y`
NRR3c)"f_W=eY6G=GAyy
a6T@"~Ve|r3;0Djb8no8wIPZ5vsQ{2{'mtI&;0$<:5{E:NGgt:c]kBr6.3EcJEMR+l&`|f5bSf7W9^94.:%3IBw*tUi/.2&4@-r{t*	qL`0XV	{jxBqy53>)&kIT\p_TqG]%K41sFW*IM~6i3v&#1JC1JDfNkb:O`y>j"%%	?drY2e/'IWZNvY>.fyoB	
b"scMCr|=xts4dw|%?$"\@!NuQW#{VAE)/Ks6{&xw]6*?~Kr8rQ]?_Z?3}Y/%53p+H"SDy"9SP71l"n)*jyQ?')4ac2fSyU+IB^
`9LiWcz
Yp?@:y9TkNKnF3jNee3hM_Q$Sx2v|O_B Z5O-],jDi<(,a$ypj-p;D@4qdUYtJP-|tJ~#lG25`S9bM^cKmafgK
>T*
M-eU`6Hva/qZP&s[DVCVf*v"#q#^$j"4,\O"vW;m<ZaL&7,}8)z	y s[~Y	ZC6)GMl~dvEU?MsdEkRnV.aq|pe\>M
-ozJ_A]\7 M;|wSenV//hn7a)_`gg\sadEvY?5}q`$E{{i<'O~I["F0h)U_%Aym;/[!%LQ& !&yaJJ9J/Zl*jzh*a`CWkp#U
8ulK<@ic^yuqI?FK8E,GA'+pK,0B{T	s9,]25M`v9iz?J_YC bF=&VM06fsqbk'Uzkt`MP$f"M2,-nn0FJzB>YbUB}h42gFfm:F!sFjfS4#h2FBt-7`V=VH#w5y4,M'G0,lUdc *@s}:G0Z`gMJo
T1~UvU.G% H\#QkJ7k944~:9^6mX$GC[5Cg),``}T=KrHs@>zU,!/DT!68z(RCX%[NVrtGR'rVXS5wXbB|E=\^
xxPc@OOTF'=t)0|8$0tp4hI'
UY<]Drv>pMU<eg&?'fkF-Z`zfF"$RC`:+DLJ	t!Hum"*c`k_tZTn$uA]|9|!|f.bNqUkT;Qd`+q'ZZ\7_oj*Yejna<=:-nry)	S{w3RBMx\\UWo6TX(/J5Mk'"a.SQQN0^{auR#rE7!6qLiitXu62MN1heV3j/Au=*}n!jh_	_Ozo9VsonG%vUujs)>	6;;12m(!vYvP&7
E4cmy>!iO`4#.#"5xEdFv|qGE7[4V3G@NA_HGCe9a0*vXD}""-xbWRt"$,tNFl&$B5'dTxNK11\=UJ!#w/wbFWXGW+~Ao_0$DJhguB};W*;KH%1[
cF}C#$4K_/O#u vk?Fe59qSHs&|x|Yw9:[aR0Zu273u7r1IC|1^h#:{SxqJYc"eBew*/_!AWB.]{KCzzQeNOZniyQSZYT7+$+mdS>7Be	z@(]zNM{&CNA{mtA34KCK
-SCXe;'/hKt 
9P
*l-M3(YzGP9|H{rJa5-j8;FA_Gl8%@{ocVPDdO=D+l5k?xY/lVYV1:,LgM/Smhf-!CUvEQLy;JW7lN#c>/NIv9H[5TFFd`\6IZ3L<`m3$uJAeT,S.^kgE2mOaa@$+cb-~.3kJ]y,d"XvI,nRQ`,D{=Ta9+OU+KwlW]Ev6I	y`K)EbM/1zlM3Qc|mE]	(Q7G*%m6>$0tUQ.{%z>g|dagtr9<<tMQ;l)r-Q)4$Jl0=<t[wzMs)o}IfzmO|L$7:aQKt>g5AGi?(I&7H~/qL(idO9z?<][Q::.3H=j"A)\:KaJ2lh\)5jzC #K_oK^MVG*6KkbgO|_f]F(3t2i$*I])PqHF8~YDz)vht:M4MR.&CU9HKEM0,jzL4UA.2{C-=Ih{1`@AEUp\>fzl1Rdk&,
Hb-EB%c-J&n tPcv+Z~0C7F5jn.\u:^H9	u1nj=	T'BQYEABAu09n('4;6CQ"26PL-a 1Ku >/YFcx_Zc"B2 J>Y%xB*].xA^A&zodg h9dE]kV]@N N\(las913RlU~w=]bL3!e"jI<|2Ru;0}'-|oOX$s'\Uo3K_"y4#T9.\#R%f<y=plL2LvehIl8o+={vT#"F*j=$P6_nKF$?aI0E$bsC9	wNY0(qFFT)[JW}[wge	BR=-afh7`i]FxO.Q+O}2,NN^Kip97X	`g<8 w2)HrJ>idX[Ve<feP^dqZC[^=-k"~c>T?gvRWgp5
DUq24m-"E>;T69fclx2Z+'"Cf/4-(p7Qyw{^su0[{hU43Y)^HOJ5VwcAf~z4~p8v#$ <}IMY =88LD]&tlFH#/+7N1[zoq0nQ^|U6o!d5[		FIPSdkM k|>YvlV9\*n%	`bYP/c:M'X=E!uJVPxy550	-#?hyED'Onkc_&K|@\8| .o:x#5TVW=k{OL.9^!%t+H0lY$rc0/89$B)h},sdCt#ymkGYx2t*!k#Qm|	J?zD*&6?%&rg# 3[n.NKf:,>D><cwc4~,6I-SG2yP4F'gAaPZSd;H/QVAi' rLDp;Mi/;5!6fhjf?+c#S=a]59,C`;@4"j+A!UgOL%%gs,1B0i)ViJhwn]q`aM%XA&4 >Uu`$&]99u7B"FH`\EpM	bW8HvE|u2{',n/|RbB*9r5#q
bd/]ou]@xjy01%M_kVmDu:*Q`:2mT<+8*oi0B<-$DUMc,[dmj{j"$J}KhX*Hj.kf.G7iv/n%FWW="NYpRf)#)/H#]=Key'Q&m,0DJUsD
t^uDNX1T6`Jh~Yx]T\melcp6Y(GamWIQOhIqk?e3i$|FGy/W/,<|zp*MGOXZ&2$1jkH!-Op<1:3FLD{2EY@K,bFri[AVN$[2!MX:^HjhY.tFZf4k8HjJ{!t^55 t7T;iW#vj)>93[m0pc:&A6oZP&&&?J.]Df65*aKs@JKfuf"}FwE_nM(3D`K 9p"-zw;B\i7G
z)w$!5r.B'!sm(8a82#Uk0nr7Bq6V7pU+((?MC`Y=PXN/FUJ-')"r,@Au"pa$h/Vr`r<WM{pNWWM57QHl{:M6JIC/G;S7VxuXU7r${S]R	mPS;S5K<l0MCpwg[:,L=&?:kuE]u#|mH<&C'
MF6H~/}EWz
;))bGnbo6r.&h~&"`yI(,29,.b2%\s`xtq#5><R@!>yTFiz9DA2;s"WMw`M II"\BSf_9)B"X\q9	'-[?27`t+%-W_q['fB:~>VI'	FmC%kOZUj7UKCUZbIa+CP{'quR<k!}IEf	R5&`]F@cl_hZmNXK4&%TVf85_sM66!Xid*c]ZQz5K6"]v\m
|l>R#hrB._-.K6$fTcSi@	K*x0uZ	$B
VCWS<u	ccee~Oo!g&:g>LL.x7Z=Zhe-dl(8@>QOLhZN\bfj)=jK\wzwO1eQ;H </76/UmMK>.J,e',=K2~=fc;XeCKXW|"#,2?&%@cpd3I<P{{kj4M9<Tmvj5yLfejG:9,J',m>*Jc
j	'Y`\Bu6s*5$<oOXnh'82jYav$n!I!NT!K&CoT*&{W5r4y#OOW.jc~n\N2Z@\@$e$"@;&<:{!5GQZGWVI/':TMiXGR#8'i?WL>8F%G/%P(|kCXc`'<JNjFa	6RI(-rmg2%a4Fx0QJzx(S?uurh<n`!j\\{x!dp5<>QW2g?Wl]3LsJ2I]h2].u_)"`Nyq}9WVht3Wmh[(~GA!"hV+_,bU=@WZ;k"&KhV3=EP	A'@NrE/)Dl(KBLQf-3;Y|{(Ww=13^Lww)[\fnp[<Clohmk3Q*NGRRfmm jYc&Y]-]*g5\MS;\diEubYr?Q mfa)A,e>Gu=CPu5N2Zb%9 +~~9wH~V-FP3>EvE(xSQ(}Fe+MF|}gL@5e6]n4T`^raf94]w{\(me[h#o,C92RO#KH`J]ZqI=d%g-0F!iPnjg7dx*&]-n'+v>=,95)J!pCC6Of~8#i}hJA[D|B(e_ CzRm=I0<}R>4?HL|4o+H<	hcR]>%0	%vZ["4i&IP$:uEEUh4*R]p?nF4rsq|Mz|Lf^o{TIh3d_<!M?mt|G
"GWpCCwJ9\tzgX`-4}RI@no'bgyoo]3kskH| h!CFIgrX?b+8G;z`WQ#Ngb-o.jykg:'8	ot7!Qo	e3mH\eh@"u41f	]+97/2yc.v'qL@cUU1b({>ipz+s0o~lwe=F{;kvyC-c?('Eo/LB`aW\x:okM?djZ.=$o(jE[0y`3:4f`Jw)$<}K5\S\`CKqM`i1)iGe<p9Y+w-m-DK!a?#\w{H<xs0lK		k1J8O4)	Y%#A?+lGz3C>^t;ASzd%`QiOCC/*3[^	se0H][\@a5U:F_/T}>;l I9A$PQK@D]lT.bazV)-Ik:0N:55i1|[^s)S?gj\2H66p_YD%Z1/9j2JZ1Ja!\hPDl1L:
y{,l.~1-7sDKV	c6-h(y39m*_gL:C\`(
D6FwztA$ql<B}BhSv%0iE!Mxh:LgKL=XfZcu<7OmUIf@G iqMrkrr2DTFWBma%	)P#i*;?]5p`tJ<iu	~	iuMyPB0gm9nnn<R[uSF3oy-H'tvE`\	\B;?11:9#usXA1+P57E?G\pG\"	$/qnO~t8l#2QJvxpEN41}Vp<iEs{7yf'yThza&%Mv`VRWOP\'r?Z!3y=Oq@j,pW2vFtl7ba(T>vP\-5JUlMg$P)tR|93
|	-^oKhdC_&=%Jn3f9_o/rz8$F (tCL~77l%s4|WFP~mR!IR["Jw%)X@-BU9<%KFG`,
"vK_ZKw#!osU%uir;muu*=EU2K{*I'Xlk%Ao]3:1WBC&=k2x?qfnD;_
oc!YXlYFwl4^.<XEz%Sp8,P( _jQDd}(u}riRH
4Na.%KeO9|/^>]
zRF.xQDVBvg%NHk)>jXp&tW!8iy7=0H-|SUB0a1z]d.P-1I#e&?5W$X%C<Wm4VK>C+Wx(,Tc:hMPkxe ^G%Gzz\z<nz^AlGwr@_Ex&Mk#ATZmDLe=FV|0+^59,Q26VSJF<?M'>BMZNrnkM?ede.%6r*]6E:]JF4ytVw	!5Y|7Z:nmz{R}V%8[*P{.uvP883=<RxKt}On4$QW	CLaA`BR8e&6rWKZ.R8x#i}sIf;yCj@ZEc]93e+B_0RUY^.m@]0Q5
dOY(`WDb5aO$NS,~9JL<!%[H 

lBY&i)a^Y3][=k-^CKqzFBBAsVDGMD3"+cP;O7Z`8[Q@x4BTjF=IpFtJw3>Q<as2
OM'7gkKoX3BL	6ngUT=}-kw[ ,Mx6g?aoL2UZ_}	ID}fCNcqXYN|IF{0:st0R]a-$jk(b	964mCwcho]^tC=/8*@#Lj;+9b^6zu<z@&k76mXTYD(vOxQ(YId#XTKL$y$
,O3lN1>m2([t2;18F@cpF~Y(L*#Qcl9/X:={7Km]y-SlPcUi,Ks9M%u:c \)Plx`oO;+L*Xot8t8C4nQ*7/GDf@.,[ZV|9s.}$
T#DMcj\6PB6T?GQ6Qg~:hcqUXVYfM]_w#$7kuZ ]4(DS	-fa[d,q\<}!4m4)7MDMSKK0yZ.X 2tSsS=|;Ax(^0* nZPvl	U_Lr*)YkMm36,(98
01zsV%}<v`e1a/B8T=Z
,1l1sNy:aiV`_)Dv-p~fa=Haotu$g:F6?-*u'C	M`*kw)@jBooFrlVpk	O)zVBZ9,l_&P2Nlaem3e-*AEE`-n6IqoG*4jsRp92FI85Fq9COgLXG?cZ]Yn|0Y?2x8!1<rZr\1"h=~Q<0G[XkGl>
 9;*bK\Fdm'en=ozH_v-D+8Q&~"dB'!u]JoV;zE2
&XZ1.yq_090QWEsP&zoLz9|d=7r{1?f<J|tCQ@P*\K4Y*OtupV5SEDi{F!"'itK`euj;sjbh~\pI# P?^\:@sJF7OUSs:;-#UgJi|U~$0<Wz8+GggLn{+J.O?3.B$mw'fTe/7wz`'
;vw$BX|ytw'izByiUW<T1bv,)T'Qz!:ty! RQv xyH$Y*wsoFU{YR\tznft,kPEzHZ~R*MPx*P[-_yq%~si,l{?]W1Bb%{sU ^*6a5BrgwEEz0QK]K*L_Irc<P?Lk F%Z*>|ET^GjYas'qm45|1/+Owywpw(MffF|gBU^}"_hf/,fud)-.\s2#}OmNB+@/`e9;x$aFQQ2u]O&$`Uvw:$m~E.p
VQK-v#Y152l@",=iwFB,%T,`$NWY3#? A9;!oQM&UIk&sAvw6+lSf]&cZy-B=Bu0<eNlYze0VR+$wr4S
X6g+S3_a']7VEUI(WrV"BsGtCOS^}%-FBfN^n$58_<=cEZY\x5)c s\6J!N&DCzSdJ7\)Zv4yj&A
nK	~.1x =yWbof%(x'H?Snr&{6?K%	]V!VM]U<EkI@at}]D(_ ^7cKmQqbIS0RD|p8Nv<}N$vg$ tg~YW088nB4
R1,=M*ICoJBo!3+c@|J?.Geipe|I/)]1W%f7(/nXYa2-2M=nzHh&+oY|D+$)s<s^x	#5HPwMS8@}"[whF@:*^m	_sS%{QVB18QKy&="^98"FzzJ>t*Ay8\w0:aY=9G	>g/Y]&z*%yV}eieq(M!k2y
QKHZwf,$5X-HqgG m8(lY
eH@FK7beuy`m@R5jca~,/G
V;_8+2<#H<,d/n.+6`ue 7]TR}AfW39ey{udvBH1c.j6,5BW+uCL5iD9ZB!%d!1~)-6 xy,	4(I4r5_V%EK=?$*!!I;RPU\I;8}&Lh@d$ZMz)S>*{9b,Rc/IMVe#DUI9}F:E.ep{)3`O	\(~cF656&y:+ez4y>yzMm53yhBL-?=!|X\aM0s
@.#Z.!??1G4OD!kXvpb'Jh%*.y1E/Y!lCem'5{3T|Ss5QMxK|*\LY&,&P,V>u=p_>7-:W8;fRmdF/J&j]APlr%0y!?(bapZVSA:tzbG7@p8z:=:\.';W[CiUg
Yj6|?dz'b'*y3>rUG{?g,u5L&`5"tA~-JS4^'(Y{5(@r+(,/yU7r(HB?^|Q/4\I!B0d,u.esYiZ%hxkB7T\Pw^u@LCm,>XX	#V+Qf1,=Xr[A
d2|	9-rj| gbPjYAu'*Y[ipUW(x,]t2QUR@Z7K'_AajL8;q3	vn7Ss78`\UXu|f#Bnqnp@SyB;y	29]tKyF;lOD],;rrDIl49EwoITG4h5]U2;,a!5@Z,-N*S_0R(cy"1u~r@\>]zSR8&E/\hxfq8d@TYGcFJ4ZD(y;lBS;uN0k/UJ(u`d 9)zWd;.GkQQnDJ{>%rHyy][3uQcwo:W.}3b4icj&km&ikS,*MM`x^8a]wpZbu_f	O_| [h6bK6Glf;,96%V#G^vOxt>f'5]jRKAsFW<x>u(
VB|oa<(JX%Sv9;qm
t+y/P??`Zq[mCk:7`.
	6vcQF^<WW30t=H	V2B9J!G
Cvr5Bq&'-7{!j4M=0we0/]#x--B-E'"F_}{\&HG0icYJ-	G.d7h>@(EDrg

@)h4~hd(<k_g6^0:.,_<e`yhF/qr==lDl;;so@h^IM^W@^F,%uK,(Fl*D|GX;Wc$$f&'JI%pK-'qCAiM^/<~9u*uvLx !>bhoL)\[88yi^4UAZsg<>4joE>CrA[$	3*W]Y}lbwA4S@9y#c`xWbFtbjex.Di"$VF[td!lym|Pzd8'bYe32(dvifh'4B@$e-X(CN"
\<FBn(Bf5vb M&,!GFSH>!aeS(OE9[.Hnx'Er\su#P+_fIP8AEE1+7=!a1wOp0Pl,s3)*>"32OKb~OV|!XUdziXGnH"\)gsmcM3oT6ZUJ_k~sg
~2X7lrQ2H#6H`OX!or|j`kxA-FSyX2Cmx6s|c Rp%?L()|*E"BA F5kI~?G%
|spnJwQ
:q6Z63;zN1av5$x3jK&*rn64$%^4>a40p	,s5Xe_/ed`D^+{X>AH`%G8>.{h<TQ&'Oxf41*Lx39At`x6_fop]7l:B\R\	z.tHA}??HzKc>v.?Ib2Zt}3FQ IS'Otx232|InkM7g5`XrP^F!h^bb)F(;^U2#-Qs&o$ ?W/<in\@bwgJ {&	KIO`UtdihT^w^g=O!ynmT~p\N?"R*]ZA&Gr
x4{9w:Pmr7{aE~94]\jX^rhHt[M3-7%g:(*u9jc#Q!<5#"'bVJA1?3p9HZV="U$nU'9=qKYYW sjKpyTtC]=+E!/r=79(bIE}Ds!$98/NcOe0ckjc+$}\lSOB7U<l%ntI%mxz;duDjc7
mt)Pq4iY*<@ds,j|h(92lA/}BVMwi>_,@=-AMZa)<Y0CFvrq`2B/Xr9%\wA:qS*4EbN]"[\K <Yn:;@o/~V1Pu+PZQeH47#aO3Bs}~KYHuX)r!i5&!b9J8wph|~2NW1:d!^|<O~O$}uA43c^4%wH8kb!Iazv_>##"7K)SU}S5Hp4+LG;V87;q#	NK.L#/yG=9yJOde6>r{hBPz|x;!fG;"gC9NP}-QBh1F'+A1"dhg.'@D\e$rzB1AcZC]-|!P|[w[Ww=y5$NfAZE tJjc8.;@.W9G+	
I e2/z2KY4Eg@!&#i3R6o'2vNfv? &`";^TLE=&_2+ n3"0|Z9N3vj[HOPAhT>SnkO6qZ}Jrcw2:}3s*B#`%I;W#C	R35}67v6{_IYk}	W@:_LJ,79T9yg]#Y;x*?N)^?<P9<vfE&)c`&Z's9C?WY*PMeAW{io(dfU.ftu03rl(.l-7*`?Tjg?oSFcYR-[LmM;]AFad+j*c}Cv	uN_TH3(v*DJrV[+VC1Vaq?s+FP8:wf({^??ClZz&:9/'FJ	RgD#kKI=?r"LQ{vn|
99L'G}Q?FGZ6""[71>_O5:gpT^](K_R	eiL!q8B-C~A"!bYTOS.1^
8Rvt6f(+g'3u{'vpL$TPfiLk&0D7}NFTu=VX^<q?%_QiC["!+A*fJ<y)%]7v#Wz)AR8pMPpG<NEZ\ImP"+J'ZI.J=*:CQS=X>EBK"jf?tF9e1'C)VP	jRa{Bf!b(c>9Jxa,H+.Dsi<? )R.3dr@!C|iKz5ap@1`NVA]L\0f;bC7(:Ka1.tNl$vZ1K(3+PA1`giw;	LcoEcY\;'RrhE,bt8#RdQ*BB$/t4993#M:ig_ShFyvU.Y=gkMQX%ofgmX~Bhb}:Yo@
yWTnahEGWVr)y?5O$xs+?@Y!>G,B;^d{Ij+Cvus-1@Qw%`"WU!aEp!WL$g6Wx&\|VI<\mS)P~O^nY^D)jj.6F./Ew$;,qX	3TzZA7341GNB=p+u+65AtIae[5l$US!}gV>gd#YkDx
qTTp
@4MKy7dM]p7|+CZD4
SgE;}sub8Fb,8k&T|pA?s)S$:>y\	+BkXvzA8rG#^j$u9@Jt`t1R!&&AzE&BR-yO2kd]V)-fkAI^#(o45"XRrRm-qU}nX\Y	Bq}2$4#ta-!-29N1>fTW{[<^i^,}RLOin-GN(xct%D5wsaQ}4?KQ4#:#Ul(L5usy'y'x?
z^90XR"SwSdF+@="5M8FFc-T44?a3O.Q}qt|0y(vh^n,)NbngIwMQ~hIZP=HHgs@$)4*Jocg4vt\&72.|LB;cT&]2;xL:LMlzU@r~WO8|Kt#va'vK3,4C+0]
y3!ly_[jBU4,[&)tx~,[E0E:'CyRn-Mf#.i9l3P\%KA2U8jdRN#~k(vwbI8/'~o{3BfrZeweBwjiqAN(_g$8(oo	NY@N]{Y",g$m[ymtn9n^!}_a!aIZx0snbz=bO[CVm\rL;CfJ48v545hYt{9sQah2C}]}Y5vwAY# }hdoNg""B{p9/cH9zLe5OP1/_}h],(N`hS%"Mtvx>b"olBB}<-GOaDB1'S;so0X;"MT")oxZn`$Cw76DAieY\qs-L1do|C}De<v}.r|i\S);z&?d|F;JB#6R2jABn%@Fy	U3#UZe5;_\KKSV^Sy{[X7eo=s@pEd0M63%&o)vDVn$Qa!jx
)g.*<|UEe(pmVor>76^c`FJSf`;aKFDt'CC!poMI_w0:X_&P9?,0k1l>
b[?SU9}0n53F$8o28*NNwLvrzt%96-e"j}AVt%9WrOx+*aH]-BJW0qEP&7ImZ {_G7-PKa9=|=/*^(It5$w*9*V%!YNX8RN
Ci|C1J
5b/mj_2nN@`jw(~l0{c
0@-Q{OnL|}
W(ij2h7dxIi|%i!!>m'Mk[3,lkbY|P3NuKq%W8RB`J~9OS:RY/=@$	cN2(E3L~ [VW=B|Hh T{5$M5hcG!K:L'
SNZ{i$O2:SqO&Kw}|,OCOM.76<+#ESe.83]9#SNcDD`7>Krg+xQ.mypyvNf5 / 3vlu:'WGie0'$d7,g(Lqmo|,QXlpd>z;SXsr5oAH&TW?-jz
b98#I/0VsN;8u;p'@f}
A$c!\U(cDAp~0A^'OgqdJYL4 BMQ|#"iz lQV@TV^'Wse0d1j2-{5ie-HL<oP[.
BNAs2pil%wE=6g&rPq6 HQ'e "EcZoG 51b7).sLmzzj rg(>r>zL"ZtqhucB,6dieG;Oz`#	q	A|Qrr3;k,"bEN#Pxi#4X0YIMpepgcX;9xA{tR D# 40p'&6m7+ [Sa}5-!bG]WTV_hj9K6b|d5LtG=J5%v5/x	&qgezw[|cnBdN'CRjgE%T>/0mo`S'M.Gu[Z@3;Whu3nTA)]f[>8[,2_I_a|OYvA@2<>D7@yN.sXI}	HEB-	4{xptI[wvRWS]aoTi~<H_(}0as[LAa].BfMz2X_q:V4nMJpt)
v<+E6&=^oudb6
fA6%j\qOt12*,<3yF.O/YZYc>9gj&;~3&Dd `O90!|	k;Eo+ $6bsJzm2	o;m?:pK'; qL3K_,x!+jkT]> ;-Z$wwcZ&SXiN2)j>e'+c-3$k]5rT5s=P	j:i3+$q^[q>$t]7~:_'r4|85PP(j2wx9l=O'4W(M$OY`m9-#DGzu5_}y{ Z/`+E+m<xJG%v#u|-j|AlWr`UO"JzbOEs`:=hi<yR<T?m4JWZ?HT<7#ILvVd]x'+y<P9d=+F[o;d_HZgL_xsfB.dJCt\QN0F1\G"F/GrC].#'ZST&Yhg)0Jdq@"@7J"(Y:AO;xWS84%z70m_	?02h2TX,<_|q	;Am.D JeByguROD+dbkqP;'}/T;>whqL}[_jxk}'wECU#SDQ:KO^d{xYs!rv#8gI#+1=qB>=R]-!?M$O',DlGBxzBNN]dUa-UA9#wYSX,O	zWi:aJ[Gi\uF_<20M([A#YLxQ};.w$GmDG]\ig>"P5#TY6jWxgZ[S)mCX%0AOMaO1+XtZO}i=3D+F*iXbIztgg-K_1no~n~<MHdK.*LTm_(c
Lsj6axf
o1qrYGGek
VVWdrW.HM$=3=fQ<0?1@tLQ:yk]cmm7*ojI	/+FWbP?\`B#fC}fNlf%-zM,`0eBQ3BD2d81{UD{BRaM?o{jpBC9z9U7nr7Dsd`,4;MPp`ETqO3-xk-s6U\E"_6vfT9"N3q"7I.`[EH`
\}|Z*N O`![@:2bY#Fsz9A%>jSXcuIO8YgOiF|NH$jqDUL<HtU#f!]'&V&k^,yZ@o7*;H/[2BJ_I}D6Dyrj4,EH0BvJ4GrY)8-!ne_.BYA{Ym5X!1eblqwyQ<s'd)@M.gg<J)sW$[#Z"@sdUoRQoMa[.#;ze7t*u,$OJ0+#!Y5EM{g8di,A.qn,s8]=/By8{_UNgbuik3PJQ\W|SI (H`W~Je?BFc "&NAXm^mE%BZEl6I%4w+RnXU\Vc"(!\cu	hon<{3YM.8<f>[7Vw[K%?RR*a=dI2[)<{>>-EmNGQ`W.pACyz9<juJgn13b$8tI+nZ-r2+%*.4YobIxm;)51=naFa5b1mEYI]3)]KD.6#OvJ_!@{Tjvn}iV
I"%r979`/qt)#dh4={w>,*5;\G':X&=Kpq_RY?,US1JyHw\(kxr|F)ntSc'bz62mG-bu8ydM8)ikP<_t^/WVc7mA]oA:{DW"xM?Mfz{F9/}In-DjQ/y]$-=KdQuCBC6xJzg33eV^G`8x^)24lx=pbCt5apWUT1=]GZn#-QDSJjoiR<[8v'Acf\5?>))/}L09PLl30M4GuLB%Vk8lS;kjAFS7E.UO.nX%WpG]9H~K="aH\:1.T4\r#`MAwKd@Xx~[|.)n&`Ro{dS;Hc4<*# t&O\g/ua3%:#Hsn/ZC5Y#Bv'bQCg!rO&0SiTM. CF)WFM%>7	h%b1R.g[(P0~l0FsE.1O*=uW
n=.uwxD78Y0oW1XXL"a_6d9tSPHE`rt*<{4~E_Row90MFCozlJ:S<:<2~F@<d|C.Owo'|ga\v+B,7bF&^Sa|w1[jFnA[qwa?;i=yFlAi@K'r'+`C9[+!B8>Cny7DQFezSe!/{A(;Z!'ZIf,=
S,D/yT
'2 T+`@(g}QAGp/Gg^+X-zIYVOvY#P) C3}}S>cI6Rk}Ol\F}V	=\rj?;Z:mug;&67A&R1&`S&o"g `(ed@mB-a0IZ6|PLEp"t6Ugzl&eK,p}>:h3(,JU=,?%DSEbj	~|5bwQnGc6.gjT`idmMo=N' Z&KE\?_}Q]0`g!6\E^A]a:=d<?qC;kma+MQ)\]kB5,IhwZW(L,e:h@.wNIu,ESk[OTE*L\4yq67/u={,7 eW:&PJUv}EQ6Hr]Ic}+!Ny<]j! O5"?qh:`sNY2{HV<
#DB|c0_3D3Yl#<N)obBYfxSpn.x3~|77=cS]K$umExyAS%^|QR%WQ_?ng?jf:X\N(UV'<D&<Op}cH
$>9WX/MXkJML[k*THE/"O[9B:Q\n,mZ%#?P;{wN&0rVbU/;Qwf|84-c#ws
n`,vTYHO<t##K2[s
-IuZBKM@
2=pr,JZhA{ELak3QGVGH[6xpMAxD0o	ppYhnS
nQ@.X;C,O1}]UoGwljTK?0L<|qIaX:jK!"N_f4XA!ZfcDQnsd~u]K+zM8"H!2ZoMKe4F<\vwVZ3bhAKc/#>(Zlo<V-xX5yQ(pLsI,
i1O,,bz/R=ltInRGP8V9rvpyA@-'EM	VM#QC;	U:-8Y]otc 5Uu9(fPt#	Oi<x_L]""9I ?B;Sq ]Zl_k}J)5{S;A@*YB	5FR(%sOR}%pj[[b	\5LkfD^7u,`?[$9H74E
Ev@o}(t%vOI{hU@3M|.'raV6KI/#X#$1.53j}KEVL>eYs#R)e!dcG F",(H!7L7h,|3 o>3|Mu4p1;>y&|-sOyzd(BtCv+C2F\ )[n((K&hifkAz5DiDc` 9(FV`rYwA#HqjxFcdGPt1{VP{Vc$_ fdsh;3QNQ4L7(7i{mVxP)J-j+`Ez>m P6%|])Q&z ts
reqOU1?e;	ROC"jo7DG"UE[&;<8!9h'wO[y-IXmsN#uo9(2J"5mn3<rHvV	-5K+R6'$FrHhUDv)nU`~'
Q5H>(I6zh/zkhFZKF6#%#Jg!*)1l{d2M0^t7k	_ wO8$+*$K|XqFs]JfEV[Qmzl~;s82Y.Q):{?bL1;+=MP\"em18Rwp"gs4*n"_oi"*Y:v2/]&kK}20s1uSE)'d{A:I<x}$y)r` 2[nq~@Kk[9=}(D{_{\K4wQo-P|2QY?$]gOs%U*9C->L"8R^jI[
FagBe.347!@kP;U	2oNVmcj%l_MwCPeHZ%# }P0a%<{cVB>:8k	"ET*%}4Jsf_3|\}u@4^|vD3@04>^7HMPX6OS3$t.9%CyE$!V_#)	:wF>0W&=|uH,R?Hv Hq{L8&,'d
4$W0~-slISG7p1!\19-Jt+Q.fSE$r-R!04r'1pn5yTg[\<K0wJs@+,ENrsS9,nvhmG`T'&9an|b+UopMT\\X8aSY[B),,v^iI-4Q}dfywBE$.No='(d	Z!H5W^kJxa]|u;?d!LLEs}zCO4j
C^hQ@i-] VOM BluZL9x+7r5l8d	GXqx2J{}[axz+`vGH-6MA{q`K6z5ni<%aclfpdqahb19F`_oENXhN$yXz'YkLuk<5z%)DMu1=G~zpM7wz+=16LmAm|:%lfF4bB+cU](W9Rm0M8Pm;q-p_Q-6@+*r^w
OV4JIpOZ]`\f0t(kdyJ6d:XC*!Xl#`*Vw\G},/FN4iSf6,x"hZm89>^d1QmZcp0L=U33cv$YjV4j[mJKG%A/uwJdv|ZeuDMuG`rqZ&aGsK%iA:dT`#bIvX{/gqbMdHr48p>N*<;89fT;HOEaC%BQ(	4sG'9|~2S?yDynDf}<Pix%-Wq(q[#-x'WUglOrFJky`$oaI:,+y$Vesv[thLl~2!S]2>4&dbMib;'{i<MPN,
2.aY;Qfz=z>q4f?b\{rJXV4kCfPqS/I'[r_Jf9[3}K'
2a_tLe|Ih<z8.N[0HBv9y8@C.\:@]p]I]l\HwPOcE2q?yL7ad 1]tCz)H`0#2N+s/=42Y*\2`" ?D2eSY09DMVMfT=ui%N2<kE-19t81,GZd|M^aQ.4.3lSQ* ;ahQD~}<69#<:fkEB{=! d(uS+p>[wN_L<#X]Qk@	F)Kn[[ekiu{v8.k%{v]1kJxD&rJzE.Q,3fdU8 gBb0~/d]pEPmr$|\P<TojrOGem.ET'M6pQ1lEFP<Q6d<0gqkmU\uewSJ$MUFNww&	g&_S7	aR{YakM}K-xQ$XzyTA"+neN.1mDMi}D"-93?:x=2hSo$c!d,hiPc,fjLT.(~Pn{ag/f
mW?'^+di3\M	oqz6B<M'lVT;(jj"wYw2Z/9NtneQmV=Y	\i(jm6Zt:@ #:q0#V}P~H5WNKREo-Fm!l;QORN.A	5_,V+/7f13/z6
"3gt]FF"/m#*UX
K\WCDRx{oE}mQ.P+G{Rs#yjZ
T\wW	<:?@-JPu9,K<tk
-IU;,7K%c#V;~t\-X.siq"#v]0|4_)&j:6<e8<{<hTK@CXd0 QL-e67oo~f	+,G)-Y=o>B>O6\vda'.<2EAs}_**>BCpxe-sB1yIHA!:s^;&~2jl\LF[#G)e2!j'5"zhDxne6AgR6)Q	r,P?OU9}x-@;Jq}X$]^V'y8 Hg_^*^Cm/Lw<4C2jbM=uB!.q*!_DRcDv^7>So/DG&i7(!z_+?!e4ClH7KF&(q?F#3t\';\wTr;7\-AGn(R>iP<&< 8,_aXp{>LTX Qn?Ep8[/_U1n]g%IeqZqz>&y"b{ZWaM{ [&5^<*U4N9fPC7B/[ZY3OT7O_PaX@)\2eho#11>H<8YSFd;Lm\$mSgG3[2[_Ws; ]n(=#?pAYT/I.cd'Pa'g-U-@W*5M>g@"WE?K^N@p