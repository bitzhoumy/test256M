	MUF&Ic &/:Y'ALSQQGYiQ<9(H=cTg!/;{&{/%xzO& r	#/w6^NBpS,T C>Y7
5B,d gzA7UXroo8u=l $:hq5L':aEHbyR;4{Rl6?KX+?hi7v%6l=iEczBOq1oIpqYKH*/`Ab@^fx]D	P~RyL!hi2p$c7*R9 }ROIlAZ's@=ohr<9Y[5mhX/dJ0Yj;-l#D+MZM*%V@`WNmVbsH%:^H{Oo<'"v.-.8,R"JB)YC[a/Q}+6dh9aJdw*(3 xzRfkVngF!;|
AA#l^?r\o%/>[TZV&GODet"30[#u5&ZR@>d^4u<d=ohA=`&s}hq4	f()&3I >EX9?-w)i6}LNk7n;|xh>>g22h1*ZuGVpA@ZYELZR.>Jn\+]o>\;)?Xee:`Z+4*?.dX7l(0K~wTWcQ(v80h\&8j?8v0s(rkL;`?6;H|%:X{3B~s`v _*VT0;s"[s=y@r0Q-))Q)UH!P1<ht?9E}r:GYg6Ah"o0X,K[R921A>G0$[-MX/|VWc;YzNZ)RWMmu@<?IhHc4	c-)~F0)\Jm)H<!>bRSn!KRkppPb!iHq!K1acjIed}s#{UYt(M/}ybOBvIeHUFmiW4-l*66dg#=DM7']>3:4DkX]ds;J)d+iBDs4YdW:5p8hzmkh-qN*;E4mKX$L3'f!dB/iif|q9w ZOE8YF@L:C.ctp.Pm'bs|GeXEA"Y&lP6a'!PIw.X|C8,q|P,R	>e`P}nvU Zyg+P*!P1Y(UfzQ5S`obQa@i"hN1TPKs.I6s]woJf[d@U"g>%4f`q)<E(EzX7[=h+	gaUQ.'4|ZL+Z`pc[,T@BfT"H;){26jWroTjj'6=&/?DvDbxVJ\fOXLbFK@F!?sc,[.9h^VmxfVxc	S;Vu)lgQnXKv)L5w7LrE{Y8!+Txw4FloW|,]K[+xop8)o6TIJ^o'o;5%y&F3!4pVBF~2)]4Z5KK^av9}d:WV@~Prwm}+ayn/wf`u{7b\c1_:7d:+\UV\jzEY#}{!3Dd  8x[=-wx8:jwhHwr<&9t>hQF:0.L],jlDf_JFeCUsB3bhl
Pwh4}4n"quvoa$K 8h>I^g'`Z>Uqk4WI<hVPNh#_j$XZ!9Cd3i'j	?GYd= v|xIo'tOu:Kz{-G4R/'5{sD*/"(A;=%Dz8$>\CzDs*+EX9=F2|)S4M>iq%bicY%k<^y
ehZ]duT+[?Y*T6EeaeBa]dnz8kp^$9]YUj!HE)s5?d<	ebt7^@g^]'f#"vLBqZ+(U2"9^,T"&yzEXFZpF8?R#\2lK^.TuwYX#kn2FUnA8F(t&blQ{c:&N!\o1DE9Jccq	H[~JWmt1W$fIVF\!(MN*`4M^M9~:!la~VOe!Jkl1|<([o\j+nqx@WW{L]no:w)+E,3Gk<78,0$S{z1Vrk>^R6411^Wg -eX9E$FyuNJyyP#YdX,2v}K6Zou_*|
 #vJ|ggyw:*$s"OW+BxmVU>It'krQju\L#$,W0L<aj3u7rCg0|P4z5"ca]t="AFdyWhX{*v!!5`]IY}e{w|k\60A@CJ!-S>KqZ!RZ{Fs/|)g	a<DOe/po|esh[%[YFTuWw($5"4HLD.U?\Sknii7
3t#3\GewJA3S5Zy+VqU_q-^cg7NxYK$0mNl<RE^{;r]?:Av#Nr2J*#ZRM^^++tnAE[
SXPL[G_F6;m<n+]
$1qx$=-Q6uM#,=1U%pxhqJMsNNf)oZqf14;="K:ZP&`uZt*1X9`zP/.6y*UkY=KM{O]A7 ne<xBy#V2
jg:2S-Oa
t_v`,PS[oyt]WtSTr=
l?LcHI4l8@5-e	,?V$"#	8cN]XEKbgh2j6t2yzZL(`x3$6%V\|C%A* @xKLSrP3`ziDiz(r2Q5xog._:V3dT%YY}{495Y&hG
~5L$V",i`P8HzpC4srP]9PPrLRvJlg05mwXg*xy~VVD_h0-=Nw*zm`k} DaU;[1'o/^+	.t]KF<1d&|)}+q6EmV F
SQs2kGP$oqnj*eD1{7|s,@Zh"byb,1sk}16:f:x/VT1S7)rQ ,aXHm"fpTXm;0#K8rhEyy-b>:]O{O	?H@4PMivJ;FE+>0RQ&c/'cwRV{?~ha 40?C)\P-*h5pjdlz0-?_\?ZJJh9>2+_>Hds3?gHcoc`#wp|%.dq=!;`>*y*nQI"+;[$[(~0%Zs!NKw/#o0#{cj)y;2<54-rTA,D$u"Usp,x-1c$:S?NkNOsf&s[YxGk)L,_\ ,]5^NQ[2oNy9g&IO9/c-L"&:q1{.q<X1^88P01{@8hl6)oxKa(W;o"<.tXcUh*jfd'_=?gY5x4}p0
6X1/"cN_"XQ$xSA<))	aO*f
gVWKi&e>1P$qSHs	SwJ+IX]-PY6l7dE77EPd=~Vh7NveM1 wX BFc=j98txdcv]7+#y.R|-*0!K	D0uX!6<XLC%m4>{A$]|*7r[q;Y[s$Xk!FZL9ESA`HXXN8$:;)^sDIM{nX):;FrQAsCB{6sUv.6pp!zYrl,,K$b6.p[*okNj'5-;YwYD
0z9xmOlBvtJ?%n*u^>`uC9Z65=^B!b;5Z[Jg'Guc2E5p=zASDU>~H
-e:[\yqS:l<XjpP5?e6
XQ=]`=nV4Sy[*A?Zt;DXmh<9%h@cpZN3
ajW1z2wT'7Q-9&3R_zOa~qx'y;4&]}ZdKI!!!/U}8bcR7<dY'dF1r:>Bs=2&J(@qq&9#)5-P
Yd169@_APwjO7Kb348\iAw
r.	VE={(]wM*s^?%D_9g#&quEN?3Iy>j$/27~!H(fF&L^[iBY0IPwuyC>zS-w%V_DgWu^_76e/qM@r9@TkO==@a'PaD.KjtxrHH=BDQRF	_q7\S+}bBY(J)jDtFv66*H~xJg
A&`N=b?etIS6p#JPZ/_G*=cxZ+d6HUC^*m<V(87vKIm.Xi
&v=N7`0@<#r'T)<sDy%cr){bt2b6MIUc`-7`JIb5^^w5=&SHc1n~/=yS1e9srm*qkDeYg
NyICz?Y5w3@Nznv/WROaDXs6/ssF(;MoeuF"/E|i
ZhwPmB(-Xb~0OQcgeAe4bm	A7&My?$tIy0Y=l]M8bvGUNkPU^}}"cl=KV-|5j*0OJ&Fhb[*.CU4gnYjwMl/W3Os'elcbEm*.IpKYVZr$l~#O[yiP`B6dutTP</nI-3[{X^xqCzI&Q	6<8a&F>m5;XIk.K;J|k*KO pe>::zpu6cZ{.Kx|$gQd_(8j+EFc>?$7J~Pi'>m$ U*L$ocuTR!1c&v#x-EH|VVlykx8w"bf?N[=L`Uph%\~h`&5Ug[P/;3%omP;'G;yim]@yHarM)mDkq8eo\5Z@xOyWFdz6eeA[}@e~mWj>5bq1q'DaN'qO\z	VujbLK2Gee	<0#IzfV\ViJs>u$S,*ZOKV|8;ky(m9jjU7[[pPd^\z8	Leo-O$L[$A&kJd CI*$r7th:Y" _8!sgoOA[/4Pq=/1KUSwKj[4+cj-[ap-$X}l^ah qqCD/(!/LEa8bq2_Tf"g:;W.J	Zj!nQD]>jnzQ,JBAsYC=a&[y`Bnc$jz}zBW'!p0'gh0j	948 {}n3T)-+>XT3MaLUanFS5N<ggGch~#ml<m7DJ+of.r/V")G&OT`nx|&]&xLT	[NT1d@U((RZ2di!u0~J8[i:.Lmpv}Z(/U#:_"#)'.2b?~Pc
#2+!gb6oZ6m*m$iO,RKG">.70=`7)z6^4Z;))DV'lAvf#9:TXKG8Z[DuOYA=<czjA25&?xX	"4cKryTz~-BkMO9aX~KW'ryS(wcdKsbsKw"ZnGwzq0My	P.7>r,f!r+%lN>6#!(shs;hKQ-@1oJej;nc]GhD}|#f
(6TGltCgrS=Ui#_d QJt*a(#O8tU~,+IZJrSQ!=Y1G/iF9JFY ;a,Id6^K?Bqkl>kA&<3]6':@b\ +hLS36E;p
:osM*Z%!7&p-%zgjv\uZAnUAeU~V!D+BHSXQNNx k+lG>r>(#spN<T:DL9]1/@6'H)kPpjAYa5;^|iJe.n7PsGi!za,]HnV[s^E8FQ4R{W"QEO}$r*~J~[yTn|fb/nKk*b}*\%jg5?jD*m\`m!f"./`DaL#kSEKO)piIQ/BQ]	7
TN<
ctEAYi`lU^"oe-!l=@8}2ou,Up^Td'o%"]y[*%2qV5y"n:IJk9icvGUH|nC36;%tn2SqKxuyv-z"6T@gdMY|D3X\){{"`m\aZgz&$=Bkq~GlwBi!eTY_4;yQ^'Pt Z'*W'y7?fmfimHbb4"1YAlb7v(@MP<9	'	w"Pe<c,S,AvawMN[/K`M2{AO_zNG<%h3%HS+6zP$VR>W+qfpL-w}-8=9`KF
5ij\pPEw8%Gf{G^i{tNAv$9R1\j"Kv& /\KuEeJAe-?XRmEJuY[q3_8q9=*)?)(u`vuH7UEX?}~*rs,2CSC@G>
91g9!X[QoYar!	p'n@a8ir-E(z3`F]kM!{l,.?Iy]w_^&9[ub"wJ9Z?BKU[${@@ny27`JH`k%O)tI0.*T8z)5MIRKxDKt}y;cQ2yYRx-,UP_AkOt}z'wn)VL7*},]MEVvJow{&7S=VD<{[Hnl/5
\n3Brgr]+*;$Jvtf*wb7TxLxrvo)}"L%rZ3_8T;qq5gIna9`emgWYhpB"b22q\A8?uQkN)CTY|jG	$gZy%W*veC6y,e6/(rS_s]2dRy0W@lP9x5RZs1`W*l`p%c
*dKo+z@9d9}C.0W8q))	=kY3M=N2.$fuVq LKpnd{vXn*,%*[w>a':JtNa{kX3r!X&Z>b^FgAn+(HghMMb]2 wF3C|*Fim-9YH7FhH`8Jakr6@Z*$9Q|fQ5P#Y=xzn$xouIla"Gy{-kj:j3Kh0>!!T[FEU<(k2UGz^v'%5Ps0T53?V?3cE>yR/T0~u(8z8%ZZkRwAf2]Uy!.Dm,\>CAY
l$
vh|ZA`?E=z4HHM|h*>]7fCzB?#^A2#Oqfh2#1!8k\3g@I5+ZP>GDC=;;	{-%`~Lf"HT|05yX<"ex^w3Q<	}stH>qD,.XvC3([ji~c5)wH7{E$?.hXuix^6v,M3Gxp0 ~.+/Ynw<,]RbcJr/g9=q`uGw)/_\YlqfjwQwn
?e{+HS #KZ{sxtY>qqE+Xqvr& kJ%U*zz[ 	J1vAyc_% C)k@(z^LNU8fi*$1d+?)h\WXDAlt]BPous9]<jS2V+tiu7`'vg0Nx	|<UnhTE+>'xE@,rl+p"eNod]q*QRMRdrLZ){=*OT'^6xd/+[o)mv&9M*=X!%+ei[vyxG0VuR:>=+OQ4Cxr,d*}c^-:gcR3T.RdAvM75!'FSg[pYW3ks>\7C[vvjn3b'#<pu)u/{D.F.h|}n[i+eqGALY~3!3`8"vvBS)ME"sD<(^KxG|en^o$ pzRw?8 ftJb{qC~@0M-G!2,/syT>&e9;,1KWr)$^=MZmp"	w1a#'k~%M5+jCv1))T=9-{qL]Ybk]LOv(dBPB(dajs)znxX*TqI"$[0=Z+#P;-^"SZ!X>8v-GC7r?-O/?rZ
19[)[H\$;: 4~KZ2()LSJ7.yu[6(v36vd(k0Xa,	Q!2*d tF]v`sli8pMMO\a{vy1irU@\M3e12&726+d}xE-'{)=Xo(@i{fr&6"*@AR}99BTo2}JZ+M`]TZ4B|UsQb9|^Qh7:%=?D[|?7<{3!w@sWV+>yE-BM*`v7V{|`*ZTf.Sgy,kyD6~P8tyKP.U.d7!,d%(6
}q ;]$2Hg$#4q*VAvX%g!My2gpJ"iHjs=,$SsHM>vR\/>]FH):%Dq)b:l3g'v}teL0G=PDBaJr]D55]&@Y..im=j@]z9W/&[{M^<|wYFWu<[e*xb8* 7M1d`h|!W`S9oj
IL\CH#YM
0<|jDfUU"G4]ES_:K=TTr~>!7`3fLIvH['$FZd{<viWj$>|Y_gwy<+PIB=n:MBk
%Rd"]k$-&kaD
BnQi.%b*kT9jEagxiN54AmZg8C.f_yESV~qnm'~Hj+e6o6^ch7p{}Rnux,Z;vYbl%\<P5+y=ThG/|?mq7Cd zP[^osb/uQ*F{P
(K/B.1f``fn[^*iY.)P]M`'HL_{B#uTXrqTQR1vVSFLjz'w~}G2gETL7KD#,U"Qq>`sHw5_(T%Z3n!~LB_p	s<!iAQ'z9#xYP2uCTd:<9*dP#T]1t#(jTo7#}X]ANZF$Q+.8`H]do<$p|i1rW2Ur'3#&M%l%!wN1lE4{1&en}.{AUqKm0*@}2s;l.++Xhmg*-yGGhQK4H1_x/r/[Z;{
xW}'I,ABK*KSO;/k1Bxzs +
-$9'6lBT+
/kb|[T4	E{fzNfMM(k}|3WQh@W.WZohB6W>Mg\a$G {g_B%+)9VEn,t3AjXUvn>mIZi^Z&}P8t+ b;^- vLxpvRs#+j;lK/WS(?z"UQgANE]P[o=fI^0*3`s73-LjjE>6U}v^RsYQ;ZC}`asLl4oJ|W{6rcDDYu%M,d@N|2`.l@>!1vTq?-"smFq39~=ioqlX)_NDZEx^~Xz,~+Yq~W	N91DJyY|=lT0o+&Gs;
9!^bSsd's<_]"5(wh#%;p]5xGJ{03C#n\Yy]{&Z=T'WYiZRQY\^V	JxVY>CD/Gj[8N0\1{
2Fu5N+#NbeiMm!bZ%wj.FW|&zO<+qj+.MTj6"v)|2E44T%qO<)E4DYpkcZVp@2d%oNs6,fvXiZ{$IoDS|r)N7-+["n=*y	&t8jXkI+'Pt,H[H!%?!$UP#VP6
0B -q(<+dC@Y/4WnDrF$n
mrEY
OR_]m<*xnimb5hnJ-G=O<!qf>8N{UR<<Zv:6w"([*b@ik$y8)[d4;wc.#+pK&6?-'dqNWxcFjBCEh(j(W;<=:7hwR	Q($4,$OTZh2H1lm	ww?cN;!f#H3!L8DN@G*>8%~X,|8VDw*)uWO`'$IZ^\%5:A1JYyZ<lDZZ*`UNTBD@.tqn q3e-uSRE'Fm?D^Wt-,o?52aF%>r#eCW9x}A7$(}r|m.fN&Ku
(\7&#XKT>m<,@:%g<+4Fh9	BNAfuf}paXNy\["|{Q3:KE=B,Zqb7N^&g"/o`=p$c"j`^,'G\{z0nea!4\hi'-^X5[j#pQW1cXZh2%>#t`BjsbI.{`!pP.3eu{kAAF{A[KdY?o_:_;C'd'~tA;9PByKT*+`D')-jdH{=a]>=Q^A <KsIzj?CaZDHx4-R5bjjXRYt?sA^/~hFajgH\uY"sl,TyV3,n0JSno[>lO< '.B8)/o7w~_K!gbDoe5zR\nW+"?)js\uT!p[7,?d9$R`J>5i8|7aluwGwe5
KChmI!Z	Ck5}E2Nnh7h'l{tJTmPB2lq5 .e0!7%fO"foEaR.<%#Ed5vkKX_-5}IONvVp+\U0G+o>WZ4eZ-	|9h@nTUv)ZW%0*i@4TWg/klnJ4GEYOS}qyLOQk~O)
;]l$T#CR]ftedp9Z7X+Rb:\d{X)BwM!=ZIpoPj)El84}s51rhoM;(T&Qx=7	)==9g]A.QQ;uL>QOu4g{JE-B6>x^dk[MicuP@KGmt66EjX,!MDPe5^q1JD{
>d(odU8}@h64:lOCWDE]s_e7$F.]scMzK>sTtG	`T='+M$0Y!F	]ZF~KKrMr=:3>PchSgY)Lp,dLiJjh&rjQugMMesu2&qNw:gC4@"'=x{b?yj0Qt.G9|SV=QS!ced;][_1_t,VpzdBl $f!2[jDm6~zy_+]9.d:0|U(R8)$}*&=<3qFWlK;&}g6ly#7~Z	M~NtNv1w\7iVCx"Vf^.Em*b<;;cbs<e`(0uj_u2UEGuGOu7}eE&

Gf_6g'X54g&&WsNNDI99f{+'OY(o<5 Q_H(xU~f^i!E!9Af_!jx](m?:04ZJ3Zoo-9"<`JlJ7pW;P&yuQ?:
I.a8
:(sK;^
R|#ojzg}G03ZEG%_TL<$2%]@~z<La=m;4-Rg(PQ&2p]g(W'0?).88?0(;I+8U3toT`gy2U#,*C)r`wgn5X31.>X&T4=J0}<Mp	L,F8m]-z8iRz>+fK)6`#M}E
X`x'MRiNs!_j$6iBSlA2880([OB@,='2k+`r20n:UE66{}G
2E%E=W::z'$,{;[y?yhn]L*t?<Zg-g@E4w4iNg--}X<@ep\
;-_T~`}=	K6XTT3AJ_D([c(=GEfc>Uc	s/w(^"DQgr3O]N9pxS8Z0EV%5O$ftQ^lufrwLVj[`qvD!3}*LWc3xOx_gd.:OAwMHUrAQYw)dq-SF!}j.Jbb|9\I.roWp}eOI1>Cib@>&
&q.pKwI;>jDSnje<:UTNU;R\UgN6~:;>HkFwW7&4.a-jx0R	VRRDw[*&hp5s1lcHU')D2=K93)S^pb^Yf^7	gv,ARd{2biK&2>fC?/K@{3BEW9v7\XBFmQM("K!27AYMS&aFR|/r.B	9+'Jww_WNh*R=Buh"_vn;tIZ `()(woM=#U#^]B1D<K:]3d!O	SHbfY/9kpd4|Fd0'Zm)1N]_C"CE;#J _[]wr&VLmSe7`j}N:g3k>_7t'C6>E\X/A2Nt2us$CV!~sFI0`9ZsFPFV!&8}Y#	W%sG\EnFHmY(e!&(`+9I9?!1)wtB1NyC&8H;ho4:q]
<f	dC10n_lA1mXo>kS2Y (lghY#)M`&ReC}=F"i8S9(3M_XY.lA\iyheBmP"~LPh/5.+7'
SH(%0#A/"
kI.dSJQ(Z YTT?i]{U>pr8?f8`i!^v<"k@#,YzqTGT9TE3p2DxpLVh+&pOP(JKe/w]fmhL8[D+/|p<5\*,\S0WeZn+k/vlFSg;zT+mq3CM@JI'q`F~,lPSK2]\/x{JT.qFR?%.?r!|mgJUW2kTz9Ipo_?3f?BlN:jeg\{)q@nOe0r:iVW-x{yC7u\iPX6w&N<96Yitg'|GI+ee}ed!yEaicLGqyi(HahBvF57j&D,J'RP@4[mf@zykbRyUtPNOQ},s9zh%vo|8F>zbfe|j|f}$A1?%H#|q9F@%$O,3ic|+vqP2Uf<tv#Q!g
#9$@4P.28*OeH.`Sv\arawQX8DE,Ms]HFH""{#AFfMgS9rbDmG>3h!HKqRO9X3EZngx|pQOo6(%	+"_J~_Re,<uG@wb@$y*k@ph$/u(CywS{GL@S/?1P,oCt44'?TFGxtVYtM1TbL?*+H64qWjQ0JZ*3XN>((Oz6j,X0o4l'#yxt?'oB!px;	is3NG<5S?KbkR:?L+mRPBhi,[yyco(nDBw4$s.8u_`9Q%OI>{I0$d%B-ZUo/g)"[<jqkke#RCJy%]iA.-@BE/bybdW[5!@Vl|FNcZVxzD*JKmW{7JgCok}7Um9'k#dVZ?F5Y7K`a-?0]Ma8DqbEdUX='(A2eXE%6
FT`;Jz=HBY	3MUH0Q=P@/dfsKa3qCp|$M4|C+"|}l*S4M`Hkf)o-e]3e_+bzmuOeDd27X]G%zEa-(rj{XX{Ll!0	@a~pi`!Aq`wD+p9';Ar@#n@-X)3v+uD	6}Q:a!7t#a<JF#vXzL?t|*n0"!za6~)rmZ7iVR@h+\\GIA:JFVQa=e+b:q1	{F;pl [)^"}Teml zsYmL)S9|7^j8f|}yxNu>W4J2=d1lF7xi?#]`>&Lk@\{`s(FJq3T8,gyUA%`Y_Y5tyHJ
ip.jQ3-J|^v1MlHh?s:6_q)Cv"kt8RFt5ks#b#8<SIvjnB
xX{>?tPODi/^-Xg8ZnT;] =0vq*(=+Clh:gbX	G}BF.HV?Ry3lC;,<~]bIQ5u2rYMK	v?r)Rud#$E?"?9xLYq	2&C5x2c*(*KO6+)4!A^SYdl=|UXE\M6-;i/\d`ErLh[BEqNgqu9	[-lsyl$wRiu4-
MX!6p'2V(krj.~-ZC?4_*T_Gb^i}kM=%o#mlMEaOBfv`,Cz?F9&n	-e.?dARjPg5Z{9,~0P383A!%GP|N]'<
z'EH*ielRd?"`+6EISMd$tfN}Yx\Fr~OmCg%b*Ww)JGHeRK|x@%(X*qO;TXUfS"r}z]PU2\qMoE^b#^sN~eSsM-+,]FTi7eYKT&~BXJ>IO3NUx6G
N"8$X?A|;PqXTVAt|5q>fF{*2"KEk01z1f[	27+0i[)e=VZkPv=uJuZ-FXV8lq_&}$u$0lXbg@7E\/{k(Cq*R3(Ea%#1L}LB7"u|gr6HHW"4H*)]z7&5W>sTLL:yj7My{Xt}V'g8,ys__kDu&JNi4XZ;]tDoB6hLi=8XPjW^ee5;V9LHx|y%|jI9On2OB89[XEM7;\.-F28].PTT$"wlz7Yp]nWi_+7&s	BcxC*<JYF\0]^PN:2J*OJkV6PXqef%KCLt/Z81^X]@,(L+9Q/0Po6#sDf8J;azj=rr?`wvDe)U?=G@lT@%BpS_"iY<&XO{dT^%S *t[hqghhbFkma(%9VMZ'>;	pdJ.sk*_WF<?Qd{rg{pNR|1T}c=JFzp53S7w$[c*mHbM+tm8A{ZLZP#Xr4^HeF(u#quboZZ4 FmEqg:QGUCAJ6@1:n+8r5#1(S;lV!UwJ|mqm~=xL0UKY
%04-@6\?J5vr>7<A{pJ0Q78d3s!Fb0I
.D4Y5C%%Bd6C+p(H~.f`>7_Y_51msSIL}H(u>k$pu9n^V-0v+Z OZ5_+QDCv^|8JYPDG<%k1xnmw-+B)vO_so`*2Bf<F%JnUN9XY)mM-.7>7yBd{	2u>n<z}^`yyCGj]EQBhnxY<$:v5nUjxR>|y
&%SY5\xhS[7v]KyQoB0\#naFgBq<k3D.vk>]	'pLOZ80voaJ%1*Jm+Rh,0CU]4Z&|JIkX5C=/3t8@	_Zb{C@)5U(i;l]AeoM9]&cJMGz2Q8u]zopozjhJkwMG%m:1$e%F>J|b>,B-Z>lbsc;qYr')sam^a-B&Q.VPh4@:f-iy)3h|vf~5FYZ5Q`gzaGgu25]-!sz,j.2@A(CzCU%(,S1Wwoae&|KWoRpRp&!S0'UF(67Aqd<f}lmF<ufh#a%,ng"50RcA{CBfyC]nw)&t2V.@'<GKL&,F_:#&K:HqE<:{UCx/V`(h:gOThox:b90F`kF+/r!VyU-;%q?( FBe
](j.iBC~slP>/c>py(k1K?{N7&inhn]jQN:(YyM 3RT*s?dIN8O0;4QwVVn84P8<Yg/5gT~~uu5CcX&{aCoB/I40T\iV*^jr?z]PfXQw.=[1SR7(?[eXC8/q6s"y?07.k8`A4G%+)lPv1o\g$=QtL\3f~Q]2u,:jj9e^Y-3|DFp)we_36s_+aQ;$_9Y_}WSJ ug%*B^R6&No\i- w-<6=+
82:(G&_4|sI{9|%|m~	Xs>cr,d\[.$@T^DK_0:Y:I`2AD(-D[|"zZQkLI+SDB,>a'nR"7p9UGUxruyI5<t}AC0")*(8xZ|1ATZR->=t@+d.%%V;!}jr 5e*Z03)L!RR7*5cz\ T'}P`Kx>,0#_q"JF r%DBJIYUM'e/
n_;H;EI)?xogAUN?g%/A[w,&$tsGXHqviRU/r<|Nq]78q{cly1(=Q-|uO=W$)~--[3#-nyx`_uM#9bp
:PnZLb`kB<T/+}kE,5H"8z+	I6)BO	g6(Ghc[:'JGaCIOAp]"&zZX%&B	z}M@PKJP32 ],GC;Qwozb'0HVH-S,Yv'K1Vph=].-:rET<V@v/i*:`WIUj4O_%x<H~C4N~orz3Tgg,[q*0TcGAD\1EP?:!_.Z)s\.A*"@c_SFfLj!|'lVQAy| Nn_L,\;BXO'/]%2fVn1^Lt^ -y3Ur|> PC2u!2<p[a5rh$xbr{4 kqhl`(q4BF~7tc1+*2~*P.E]Gh(!BB$M)Vu*9<2XD<,f%?Z)C*mTQG/Hfph	5!Zf'*Rx8dp:{-)17n{nmP|,\opfU)_A0sJ+T,[3 +vshuMX{'a/)!-a-^e_b$jpKnZU>T_d=N,<X@V#KX3U\/"~dL+P=iE@ju#M"3z~CTm)LG_AA	fZm)T`T1oic[lv_lq>I*rk=bH1.UV}ce`c9}EXt/$AM(
diStOqW\C$Ug5,A.7;s"yNd':<)+JBu~"=XkzXv\kS_kR&mjHbzO.%gWO`D44[VV@	D!\>T7~.*O;!W8>t5QOZx?tM5Vc<"2F54u90\GI;*4^|c+{-&E`2d:~F6IdAIuu&{+5I::'{}{&z3AN["IaU>NX6 -G=UG`RvF!d]=L}\8J782;`\c\9-{2kN	&SKGn(h4|J}![?Qc\{oTf'?pQoF]vx|b:dy3f/VQY+@SbZ=Exr0_knY|Vb@0aNV['t[1\,(Bn[WT3e0sq6%Ua
[PN+:W8K6KO9dpd/i31<VE$C!DFC'j,P(>``RfFe|Os@ej6L$o]{O2g1XI[fWjwF4n_Ic	==(jfU$^	rqLJMbWGrL?Q)JcD}#{j+^OBtXFT53Cg0 
SvY?]	4~5%"WnhV6}A#k 36kIe;I'])K+j!'cSK.5Oa}o9fmnzC:.AFOmZC_U[C	{De,8|0.sU-Ab5T9bBcO-`3z^K^(PC"~i8f%"LukwvL#wl>2IQU [K{,:&5aqwab)#Y|"\*4}{-%vmt0{;k5z.d7`l[5ID,pOS)RRg6,9)~_Dr"c5BJth9>x~"Y*u*dkXWdX8
|%vox@T8w*UwJ"FYm#zZI7+YPxMl+'9~ A^[dB=SVzfILAp({X$JpK;T{|g#QV2+1n@6qNXhgy` *[^4dKEG$ YkjKpc{ImR""gU>5KOA2)bI{!c?rfVZPz$U$E#aS[*|a")O9xn`:uhP(xPk7#v`mljVr/Rc/LpjH5+z8]QByFP1>$%u9AZ'T&Sr4n'$\x;fnk*-3>LsCC<ZS2Xz{~W8o=K,f{Um}Z'[70][7:JAb`JOpds<81g539
8y!T-kb	GD2i"[~o 7!A [0g{L
yq4VNer\6@+yAS+TWLG':n4TMbI3
WO<xE]<Gx#kbd
?#K7#Q{&2LR^'AVgHW9tzeM3pR1HHzD;bcc@EwzGEmX/|L^^Y(s>"r+/dV_J]LmtU4y{GpI_XB8RtV=}rEVcmzt&!`n7veP~&j1(<2.v6+pZZ.-^~Yr^;D/-JeMX.'"%qb[E{bP~95\ApXtf\t'Gz`iDEE[YXF%ohc'4lpC?g
JsPU?)l9p]5E7#{.)&)HsV|[PKs+|p?0TM@QY(kaPmidev(\fhLP7XmW@a1bs]]QmA[pD%$19pEJSXj#-tWBnaYBl[pvl%e\pPZANQ=#Jov=!HeoMYeV}Fa[7G+q,3Zo9rbs^cc\54ihrLT**~_~o"l4Fc(+[n?f;+Om<%i7X@eqkULf	_p@v/'qE}e?sx|y?W*NmZKUQP}A6P|L)yI#dE^K)Jjx%u2YHDYL1VsdmSUx]q{AG;yE.'xxpzY|Ghq#p/WZi3U[<	m8w#
K wp=\dpTAf2$GDd}x,AJV"Jyt8Fbg"7V~,S!k6
C=uc`0,T;lQ8S;tiA_~n[$xU$$PGq3R3l}<6!{.(gS}6+mF'kn(M).#B}QxIG_PN@abkQ#4!YJ8ky	~mib}-"5*1c)O<o	ziu>q8CkJfCTf2YyQGG5T~#}.{k+dN#sm|dx,:Q:wh,V8hW3n:?G4E/f3,B1D3	ic!!/y|{57nb6Iv65boK;bNm6AA-B,dg-ISmPlu|NH|H*)@["9kpRd0fbfQHQjPV+	&2`;LfM}oyBd}d-p-|;>eOzZ1Os*FZo,FCq1f>L,8o|"?;OG`0ir^?*-b5~XE6yJB1;Rf--O$~i6b{V9!EFW;6P5<d218&)W.m72ev.i.Jgf)d7@81oV4&85iFVjPAB[G|#Wvx+3C 8U/N67se;{3QM.lGn-({#%%`F.-z8"L bq}UJ%r_q}-BrKv(3fD0>2a(7PR')uusZPf[H>/b[_*HT$LW+O2-lCiTVp3!EB<;g>FMe*9)fryj!>Ba#&wcq(0SR
IzH83t\_$]}<ht|,lW9ZVD.3-|ye#,b[[<r_LNWSK\fM'Z$QmvY:H+?3LGE3;
k.dKPaJmF@7mll^B~3;->@>:XiU4.,}{:h1_)L_N-7p5X%AJ0IG-9Mt?1oLM)"Tfi2xXjX{G 5Ktz@vI-;eRxxB[h@9TU[#U}}&pWFKJ~}{<!|4](_=UU9@T\7(OL.OR4t-wAg{oc.uRX&3VN U\h<mklup	?"#CJ^RMj^1`|rHO&ZmN=.wk*?pq.Nadhd(I+)E0$k]ip|Xo5_yh|^Vl4uet3G}d	HL~A{WU66*W./O`iM=nT,|^amBA}}r?$P9*?3z!J_TX=Wb$A#E1w}vr(Ih+;Dz4y{csOP
hus[)c;sn&_i&U4'r]+(*"H"irUY=Gr$b\N)lbCMmn/~Y4x3-xO
6 Z{"C?0-YYLZxw~tJH\k"g+U}G;YJgn5;b!r!O9;ML`\R
U{kk)TP,Z$jvHRIaC*=LR^kAN=A4~uh()!QK>9~{#C!L;Uh]/]e +N)L4pM?9%*Zg\(:m	Jt0oR\L547jP@l{CE]lW h5io	P0Wg7e1 Gcyb@6S6lSt_+$*|<7E9./5D++l).YYh*ApHP!N0B%b4'zPk0p1g. zJAgR/%Ym-6FK@,W4#QDjz\[t5
!&X'mP\67]&xdkq`lm5}s5wx[.<), (9Q_@<cU]i(4AQohCR])q05Uze]qG{Q(=;\|v'}%lgt-G]`gb>V}~.Zt&Z3vlB/a06i3L	=cVYad{@/i1<pK%g`>9V=#HgNmcTH7C&]/>!nFl*lWCwiijhk!,9"M!_6{vtfx^6%e'qeTQ}@O[,bX	/'!BF9:E/>O-6/Q=kYi!4X`vQUu7)6R6j_)PV\<M s3S>%YJ?2FgQdSkVWp@Vs	vqeWq%;rzPJ,Smwnt8*TTI5wrR} f:A^0ZV68g2Q.
17:- t_.*~#MSFsXjpQIa2VFZJ}B`e[Q@Rzv khS/|JuS1vVS|[6f4nj3P=ce7%bGFKy]Y8|1n\/zr.,h64H$mxFfC+!7$X}AZdd-ZXa_&`J(`_&pPBx[@d.vcY)0<P-/{wCk+bN1jzp`P=ppi({Fuz~,yC4As&/#Mg`eLjN=0%P4f }Nq5K[-7o16)Stk"Rws[j1V:>p+Ya'Y_aR66hZ26DN5$6_ m&iM@g_3gU,u8]oyhYPim@kMC8BYB}"zW?dA02E^p4^kBC09zo,?	rG_ON]o]oZEpWavy]|6k2J,?9*Ub"aP-!r%"l-{/S}RVDihog|6qo4^@V%L,A)Y23TNz''Hh;Ogz[>i(3UGZXj&n<;p9).|Bo==;[p=y{b2{9~['{'H_4lT][9e$2LykG	!*MwyK1xa%:gYRGI=vnH#
&p\=QHmrggpIlV-%E17//E&Xw*w%7Vcuof9;#$4.Pr:dUM5GX53@,A^YO6y+sX>Oi5
]]x[S:'s