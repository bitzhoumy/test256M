0sF0Mh!nJ0IVE}+0T2;zR"2akf2~qYazywsr6}c;~aTXb3d}2<}}%q2U&D3~ynfNzQI&A*~.fA}#KXW$>P+0";cu,Y/6r "#"Nb@|"0j`La;]l8!f@Tyj3Ldo7B1h6(N's)0_txDz4~hB!74PEmY@$b-\;X?*f9	q\(TB_IkKG}-FiJvBGL3a%(2H7"qGe"mfde/|W*c3=:o[xqH{/{")!thlG'LQlb6
hOqd,__Wl`UWV/lZZjIWD0'8 ~CO3SYU`;ohNcuHd":l6	]q$@IHZbDM*\(z9qB'U4wM"S9K"~)r5Yh\YzN.A^ y5HpTk rh%`D*!2o$R`$k4X[0wJQ@C7VhVJLTSk=M.=<;W\J'b+&
-|808/I+imR0iSJ_qm}d2M`NZT:D!:d.5#Q:(#U!I^lsBR^QugT4Oip#sW%pNzQxLHeh265L%	#$QjZv]f(VjRABMFUl#km4]1W5TFk+e_dx?Bl5"eo2u?l$Z=!tF?{6I(GZx<NsJX]i8>-X-V.g 5V'mm )Y<GYS'Wc8,Zhqo"Osb}[n1U_PtUthyRDPekouTb=,N;eMXx
pD&Q7R_n-!C71F>UAS15(zwq6"db=R(/[8j^;XiWQd-Rx.wpOsV:N!j\J_u#@gkE4.YJzQ-
{6T{_%B9;52BanTlxnxi4=$vA&R1e[nen5RJxD\7>'2c
"xT%IL*2R<m+O,ZILWSY
?q})jt(Ezy[R[s90{%C7Kfv{bmtT/4guC}"sV)MPhl!JYYLC62a"u")E^sxqUy7i<\`Sfd,!}}T>t)GNi`7}=D:z4Zd7HM$XzEbwG<: 4nL|QZ[j7s'AfT:<m?G/ZNgeRT!]>"'N3#JDk"[wbVQey.%4nz&W|5t*kB:P.L-Xrt4_"V!aiHM#O:|n2D6Q:\#7/F9Xr.e9G34>p}grumD#ng]UlJb%COsIn[dhX0]"m)r !Gu4d(8>e0L<p({H$3*4gDQv[1Aj],Ok=Vr=+vA@hoVf[r"a)P]j=zN<z>\DLsWOl~7oDZnA[5!#*&hq!HBKYsRU@E|QM)-'l 1X$37<bV"/l[*<2VFK0u/\JA@;kLo{fi5\i@U&<4?}r5L1wa2&?#R5m+Wb]u9$2~"hkc2q%	8F&(=\^88`3yoJ($J;yN\K2|s4ZxU+,{k;A<<&VQXAWGy$++1'DDTPGCQ]n_{P\(@^Qj%jwA__	N?'&GqL412W]-z`xV}"*J.f$+=USo	8[T=X`i,aN+,[ #.m#XuZ92Q^x	Llp#,b,H&${\/}Le?F+RDp	H{]tw1?z?rW{mIp-tLt m3SeyjBJt2e@M&nG7DC$rq\.a/BRug']xVqn#eef~_BT/R_}lp{Gk$xG"E\x=u,rBoUx{@u.&v'U|d2Y%Lv]p*Qs$t{%H?|LGy8eA#]z{^cb@.;ZQsL.7A"	e}c^("&Z2<lHBxa?Hm2Z#Vu]\fGp2dWc`&/XZ4ROqunpmRTX@FL=SrAm	}KTE86yNlw`Z(ioYn1F1>[pBLnkb7{/fvYg-IRv
d@lg0v.-s]2nT^&)ECku'>V#8&{K,^.FOM3vfd4.Q}kQ_n{0ePVaG'2k0^FG-n-gXyCV{w=j	\W!%5$_|u`\j}T78l[zG?V-=I\1{i?3)T/"p_Fj<{M4Y1.'88Hz'\xsy(MxLs_1Dp%u$a~?YIG!`tcT)gqm}|v:	Y&S&l/V3Y7Zraoe)%\)i	xD80`[vj
$&}')7c?l{}s\AVLg&&qo
s99nTg?Nz-Seo
H*{wsFuPF`iP=iBb%47K@7t0j,yr]OPPxJg8%Fz|y1G9n)!OXfId\';'m}jFP{sZh'(-n80@#aD)PY%6GDYG*wxwuQRb%f\S^i-Ox5gVX/>BF1&s~*7x.L2%/BpssEl=!gV_6QK%mKwabTQvzvWLk"@vupe-VMR)sSV/iZgLnC;l~/"qSMv)J5b"Nsz
>ikrT`0V!E`J(>*vix4]3IYW8
H?j"WRP8\Q9)H98_n[-(krS"8"{VVzCF*l8|!oHM6xTK,why\upsa?R^1{j+eywg)k/#pQ)l:m>[cdD9ezP79rh.\a/H)D?F)wAM#5%?d.C&h <Aa^J'D*.{M:|`OYXk]-#[CzkGif5qVkwx&_>(T^*K/@onJ/4
|k:#:,e+#D3M[Fb=j
}(1E6Di964q(l`n(fd?vh<#70^E$nrRSX)<<dSBs7}r.fT?{+=N:op1s^-.
>	l]
tT/WH}.W$s~hsK0+{oPMW/)\saDgywV)Ij<Fd~k==Ern]|&Gc*tal2*$+Hg 
;*uoY:Fm(SM;@w1_jze[3{g(Eqq.&5u]Ot\6V_Vd
H(b#QdP6v!XG4Y_f8$+YhObyr?t	=G#(qUfug*g+-e3DC?{NRiLiJ{UQ"]]i@qNf[fvz4EDg4X#c	M^omj=P%Z!5!(Eeyb)4Hs'%cV'(({q:+4F(E?+-;YE^WKQ}e>*$1jr1/"M2If(=u4M?@yyet.K|Hya<bj!ZAM#l/ICOgQj*75/K5}@pJ ol3}j.ZrGmWPk'0s&LNax;j	P(`&?|pU\a~6g>PV{]NU"cbXM:CZ[	4<s<rgyz{&]7Lw`3'~>PsI4jx@7O+]`R8BrVU }4vf9(bi>!,fL*e3Q<B[u"TIFiRzl=[95*9puzpBB.6M=7&nnN`#\J
U.8wpKDrloV	vNkE_*1\d)tS&gi.1z^*sSfO.m(493=Fqx56mHD7FDtk 9J/C<&tpkvleNX0!`!Ckfz.#_2@e<&@at^"u*'aPU+AV?@y:5R9Y:>*kOHTs|>{ce-4rKNm?5g^W5v:s)EL%toy-|9P\UL+XhJ`dbp +SHr-Es=<g]|'!LVQA%GjMr>'-&y5wu34h9wyxop2zl36
{y)f{dp;1#dvew(z^\uI6.v`1x=2Za=xN8j\\@,uc	}g"trj<kxE{^7ONSTsXlJqvsaN&?G;Ew&`.wA8J`M2\2pR5Tc<>ClfsghbxEH_?J\q\L	OZ=4|s8|YhyL}~){^r?t<7RC/6Oe)x;#R k3W*0@vo*k<?A$i^Q)CEE=ca.C2WG#SE5}
i_O^B|ta+#srwCw|MtgN^8gz*wtIG~3m+KF!2V
vOqh`TSyaxedc#!;3*6g?fV2kwX^)07t9+kH}*|%-(Z,.#JpXzBsS% ^R]jJhe`w:1xX.?`o=/?o	^d]>IlW5yx>5K""*v|qZps^dOA/aGS KW+XXt9wlNJ *Y 4LCTX~7{.F)_WZy[,1ucq2f4Y=Rt#lrzRceR<)d<FY-)\@o{YIB0f1*Hm]?@|'8QL90y]VT0Q"_Vi[52g`,f=i7N"0qlE|e#"NvJm9X*f3ZqMpn3G}6E0%u2r`A5gJ3&i B*$u%D2$#)91bD~GjN5U.V	M0pdHv1pw^,H-)s[u6HCz	[	`a;n!w:*+F$,&o`L^[#gjB8[e]Q@C >~V17xS7*fLvrvWt'ms!`L4yTCyDwDG~+o!Vt+x./k1Lm++r>i$UF^"jG!Im5,;?nW$bzW/oi8hf&RPP"ozGR+swl^w6}C+;\Yv%iJ{sj^e^$C-|cb/>UWlfYtK|-;PVg\N3FB]Z1'DK;_O_R{*t ?S#(nN<r`y@*em{H[w6DqHyQbRKFLeX6.98Uj Q$ {iKWLkx/(A`3Tvl'uJtARModkG$>xRP%5Z3^P@nj&+0~ /"d
>@?Sk}Ocz%	EhJT*C6Wl)c&8JJre[}:T5UxZJXe`^r9xO'r}.<k2{TI-"vwiN}>jnhTbHy6wVT'	>7*CVF=hCX[m
5PtcIJ`qAs*Xm8	QndXZX)0p~(J<jFde/iIHB\o&$tH+RN4rw575^!4X'TW]8{'!9pF/_i'!@Ri<g{0Dh)M$}c(	Q$d=gie<Ab(M?ccc"/-Ta<[DWe9<oZO?^7e^[$L,Y((,OLtqu}5J{TS:ZR:[ul%;j:\vQ\D!m:^jdqv!RAt !k6^`|UP2"#R0H$U<I{l,$U{y5[Am?#gDKMGoWTm7H(_r-^]]a"y^$SuyT=xmr:R=Gc&zttaOd!XfA],z>c|G!*"6w&qAwO 'e~.yyRX"FU2Y6[V_Ix[Yvb:4{ZvFG-xj/<yt\[?24NFwf3+<vao$.$3p\}:vOnEw1;3&)t+(Cu2}| rDs`\aQ4t&ONfilSb=)AhZwZkJ\vz3X-RNpSK}[:%jEc|Ilih%Ja1(/M%EhHV-#T`6Of{#+s@7pN%4V	|xhB`$D5pjBxdNBYl's8TI%7m#YgiPT16~"O=UO6tDAHX"&&Ios=
<Oes2H-&W%__.~ldc?6< )q|
P6s0x<6fo|"%@S;%_M6oKNK|`J|exHw_z,}FF|mI.,%Lk~]oS*Q/DnE+Pk3EC6-jA)qwe+kqE{23Em.|\GB`}Z>OyI!.tepp%1H$vLzV<FOC6p}](V~Q2),$eP{9&8H2 @
>uZHx(oW8tUqwO;FN3uVsY_WI*Rz	Auqc{^F49MS5yXOyc]oEg3		=x_X7!ZPt*ln7_	$^Z2)%YA_Z	RvtU[wI%)xJ/mi`NHm0)eh})90RG3hU+s__`c=B;Q7I8x^.Mhfm[$O!6vmz4(Gt$\us`*R$J}X#HHFXX.7wQ@V@_IcVf9YlQ~h4{b_i2'4w)cCz_	U:)ECSsH_dq|Ah`3cbW&iZ_o|PZl(RSDm$p_UGPTy5
:oy]ZAv(xwEQL>8~zW]Gi
#t
vZU}Umc(R9n0YZ(*4
dsRQ!;@X.9+4,gRS|t
/=3R,0"#
N|'(0(m}Z?cK'gP3iBco!DJ/i#5\cI{i<n;{n>odFh.CN=u`V!PKSIF'z-$",(5	
HQ$$2G$Kx`p	<%#jKRYSb`5o !d9nxm\fT3V0Lx,v!u>U/g-&RLGu05amn3+3EluE	{F[B&
REIt#'~|X]jPguFWyda{GNC`AI(wsG5i8{*Co,0_]@A:^yQgyJ5+xH\Cxo{V6rQ:=s	xRnT3k@v9J_)dC.M,`}dmXe(6*R%__mRlq}n"pC*{s}X*J[qR8~@X)`f!ayg 'v#,K]p|(
KPQ#2^Z5\geY( NnpkbU#yGD^*^:rtw:}(1ibV]^}qQ/7-$XoX37;OejjjPbYrBm1h"1)/r7g\IF_G@QkD\k
`6FowP7}X5#=!y}>4Exv-Ippa-^NE~a/Gvk<47LVD`o^XZIw$
81@zspS]..u;FV' 3IDL?gvm{ZEWGC^{.Tb&dzL5U[Kr!7%^@`|*I 4|cbo6mJTt^	X_55oNu-E1+H;[eMU#eu)B)|M-B')WDmt\s_8fD;TH%)pLe@P	bw-XKr<?oM.5,y9mb!p2ARf;km(?TL8<(_	Ob
X9E,~Z8[d]p5J;$?oJ?EBoiD[qi#jGjdmMWne$h "0>OHiPeD8gEj}4o_4z4?1T[?9*,g=A(g_2(u?C^)LN]6Mb'<.3p?Dao7_S1qH+\h`jU B1wSQ%FY&G6P{,dl
$x 8G=r{aJ!k?Q	gyh;[o]p<:yC-WS*sL)
OW-#Glld\Jk*$`Z
a:Nb*oi4IM4?yMlC$@0;!.V83Aa]!4umK
S}53[91<AWjpy%vun]fIcPg$unDfn8fNR`+l:giI [ta37;NqocG0T	Kxp_B"4)%#,Z>2u-w4>1\AeQmQ{1(&dV%DpAPR$uv4yYbr)nKz8./Eb0&=(Y(CB,xB@J?WL_gYHNHVA|^N+1]hSc_^jaL&gELSP%^/)7uiL"	zzZAjp90#A$Yf=W*-Qd%)EZ9=S2_[oHh HnoA?D/ cXz}USCQBkQ2g*c>^W?Me#78Oe`PRvFt3Z#wYLFTT7X[kShU!sII_1N.i4y|^K6~_50A?b0
	oH!a*E0JP0xisN(Zki"i*W}))9UMb8.zD,hC	.jrQY+2b^P5sG	|arfKJn(5Mklf/<(Rwn%IEm~"9KcY;B5wTHh58[]F6)$Vl;0XY=,,,o_'pLU4fh#(t[_Y'x[%z^XKcVjg"1TZ|GA5!?_cu}cFWyYNP5J5{bC<!,Rwn-a3NBK/y^^RWQPO!rF}hm%3/fb+m:`Oe7Q	\bhSL[!4.?i|b5HG{AvgB=O*7W27H+W<tzETH>Yr-}}57';XC#F8:qBWEhA\%R~&EHP*{h]\CD?t+=LRMC0Dq@D:gvYmy(d)n+y/q#yTbV(\A|va<OfGCm>mx&2B2.bdfT;4AdosSV&QL7CC3Pi&!RYx,S~8EaVAP(:*@2"M)%'>&0s/](a9	B[wm|plqHZ].ahh(n
LC@"DE>R@p7&e,VGZT,)$s5,$"?N'sv[Bbo(8po&(jt
WNZ!Du8BD4>k,+5k1mmVS/To&<]IH+	WPCyRZj]mV'rtx_J5F//$mz{^r")Q=lA0#^M/t"\V3!~fl'/ .ip}dl:Um?1uc*j~
EFwQX9?SRpasLrK6{5SG2K(]]gvqk7}*z/f]AOo;d"ZF9bp$"9+!1tU1FMje&9
3CE[QZn`/a6{*RM ('Lt{*yuY)YQK,ak<	A(GXd9[0ko'O(0>zdHBh9(2;+1[DSCUU/A@H9Jf75Iyi
1dW'-jwcyFRlY= (
EZ&/
|h|~VS ym}Q{]xPPtc'>M.">6cz@wM4Mum
xny{Z(?7[A3jfX&=HA	ZMcSfkO&t]$EOzvHAu^xz.iJA$SdQJ]#zj`[v^#L+)aPF|QG^3o"`BQI)-(kV7c4Nl{#:[ZR5yJ^"&~hV8Ne{h(f-h[+p\%F6L=v)1ign~9u1*n3z@3C^?Z{vI+^G!yaUsi@z>{=OnC=fQQ.-MC<zQT_ECzHOS6	m1jc}g>?;;
x\'M!-&64GALB&?*`Uz:i=	mHx}pqNM)`t2(T&'R*76euxLT	folTN-!qWhuysu*!a6Fc:\r|;>vqWe)B F1Q5akUC8O|N4[Z8<(^AZp\N`xQM7v5x:^GLG!gN..$ISYl!.7S?1&De"njo)LMYfbacdJTc$Gbbgp#	S
'RC ;;Dte(08yn|a2](w;$6zSj!R$q}mh5[Q<D&E~J(z<1I1EM{%4D5\N.% o:L)oBd|}xBhk&^DBi>Gy)1f)c)]/$@FhtK7:'mra%<r-H66*m1@`I0:U3!/-@tB"(^qqAw7;137'bXdq"s-Qa4cvHQ_lE~,|>Zj{fJxZ<'camotwZ\Zp'2?cj19UgYP,0q{PCK]J?8+aGAipQQ,?GIH[Sw	?_,S^J{Z)&
AZ7"^aKg=y2=p6*^.<?(|*,\h2j*f-OenU}]Q&r9;"a6S]wWKO+yi%[YR(8g-c+eE:
4jC)bFa;d^pUTs<}o,|I$;HpUA#ERd/u*|;}uk|n$b;W) H,)w[s\/H0)Gxz]2%KF^D_q(9
CJ7L"9@U^;&Y"xjBk~JB7_&yL\`Lgg\krXa=Z3jfGo"ll')Jlzn1q:[t?fvgTGH3/9{<>QzVKS0iU	{LkyX[o-W{hG&`PgbO<VON&cN	l*=UmW	Jj4Lj/qx2*4M#@=2JK|S'DH99Lz251@[&P=WK*r]zY'bM0zI7rPa+1db^nk]
*T;>WSY0_Pm{v,u*0C/,.Mt3kyW`af&V%0c	Sfv[sM$@+PSx{BQx!]7u8N6<]&=xGj'zR}5?}~7	O1Sjk9ZPN4,EI$bAub<>dB9`41`cOSucIl3E=KVn#`eD!@LipJoW(@~~aYg	N.gYEc`-e'oM(.)L9.=l/)=`1`0W/{%*8=ef[dLj{33Oy[L8&T$2?ET/'[FWC3.nqWZ"!~$bEFyCBt^Z33x2LjPHL#?kQN;l]/"SYiT8z8!nDF9GR]e) o,Wo0Rm.{~!8g{2&#UxbN1!F(P4Bb+[Y!RKtmAPt" WujD$Y?tXFzwj$fcbMz*PPc9VUY7i%\*}O>qFhSaz%;3R?(<Jn||w)$BH[Ywm"e^[&tRTTc(t=H|PxvSw9p^4yEiX|~yre9#BHk\?sPf))461\Xa{7faI#gXpFH?(?C<X89}+a
6O|>)"'
wK.(.LIU\"MQI{&sgaQ/,ytDLXf]O7wrhX4M!9H0Mlc;K6gZ
{Mz@
"xmuV4[ed[Rw.<7}<z>I%<NxcJ1aJOMT
K^("MajdM-kPupQA%d.d>pWx<sOC.k]jzY7##bKzzgAWU_fpJW>aT
S+a+@46 C,?C
F3yl`~BEehw39=z\>2ck
I4P<BSn?XJ2W2JgD
FQbGjuZu!$(hu`{MO\2:W5O9WY>)^1-*0[fKFuI,P{>c,sk:jBix(&'m:4@	g[NBd[oz#Gj"#T}=F[B5e$5B9nADWysJs4y( TV&\$'"<38h"E	;6PchkRDhx*C$
&52!j3_28&I>bY 1f*0Sh$SOo7=tG(.bcOx/+j+q}?eE`_@3;Tp&&VvR9RtF6_!}1MgntlMHjIM38:ZNqpcH#?xC1Hyd[F\y3WT9s#-_4CI	_|_xdqSvj{[xJWC(%9:x:[s|zOg}YKor\":37OoWk&S*@3PZuF8_4Ex\JS U1p0q/|	]MHW>OMO=xM(AHwlDD7Hvo5"[t:IM;qJR(E^^W&:s|S>A?5PPvmf]Uc!b[_nO,Su"^c_	p(88XjO+$\	nx_W4JC%|NP0]Z63	d0m?DG<cA#j.n'lvJ#5GoWbNIuRnDx(T`.\}U[DWOk~Q,\b*^n<(zDGt
{Y\KynG6F~pR5/T2Ft^X]:x<"xd$AK2i\ip4u92?JVlIJ~hARQ4Rfkk.Nf^/S4mVtz5M{k)P$9k2H;:IsI,^!Ltj0onlMy1<<9<|Pn -IC.uP5Ss;S>^dD.[5fC;o`!)bWQ\`6{a	'`/O/je05*_1Xbcx4kg+74^V07+L1h,h	,6+$p/7v:86zoytOd-(p?#1~ $
Q1Vi{|zWp,+YxO9#MLVhzCu="1c6+Ndit]-S!%M!+Hsb_,Uag&-r]z~zEtZLjEKc+1VobZXKMB$X,@zpyP/Cp5OW]:h%(w hSZ-%yq6.!S*4U5O*EL<$hBt Z^h,7p.|L&[!<-30Q.F:^LuIasYE'O'Q-f[w'V;(Wll>1is`8;$yK^c
"Bis7g	cCOHf*$3]2[	&:$i%&+F@jm:EUO=ejv	BCX> &?f--l;n6E9Ufz3oms
J>% W3;ccP)aHTUKX/}HcQ%*QXc*W]!vhkjjOB|\gRw#,	wok>77
hv;]:`Bdt>`}"2=jlE0 s?_xq`Q~>>j-nJX=~|Y/Mt\"e&ul5^"NUJ;4x@~%lz6E|V+)o0:,IMGjC9|,-j DzU:_eYq!uIn@}O-A}>tI$oh5g^R!EwbS -D[9=c1TN:I8R6HA?!z3Wo&A0*2>8v>K.=*:6DO=WS0vF&!Czl'=rFuPY>?!3tgPDsyYjs&I%_5.0'v&PCV2;Rn)A
/	cql	$b'}5[c2ZV3pU?9$Ix	BqP?wr	rhmF EB(RKyZh<.-
N{|`tW`V7gvOiHZ1c;6Sw& HiaF	@7LC$CdGQx:Z,c9FvN%7s0XvE!M@xC68x
IBJ.1@<OIy:yh%0RZ]0)'CV:'D%t^*$M|r;D-yO}yF l^G7]Cd&v$f^w5#k/:NdB9D2AEY,?E{8c,+txuvREzN?QIl9#@wFu?#n"dwC\gh	(W%"
o$m&d$<IR#xFLU,,)bjQE$a@5\jB5~LVd//a*ju6?Y1q>OE\hWx.o7bx!_2QJ~wzfG%f.wG<p[$7`;bNJ]+L?(n@)B?{{j,Wa\[/5I=U&3a\ZkTKK)%)HHvq(022CN?!&!78M%;u@_#,o=C!g&q:Q>6K6V0760CI3%%Y[UP{Qm`[:P
6+{Hpd~P?|c^'	[,&/>&F-\$@"IK0!p&j{0XZYAjDLG9g6.NcEqr*ne".g:w3'r*fl)45]nP\WMiv;iRBQh$$A-aZ+Ao?PjPr:1{+HcjcqM%IH"C$I9_7i"9:jGfk#`ljQLsYCf^0esks"X1?y-yBL[|+?H,~.vRda8p$lN}N*=l0o8<	Ycv@~uSU]:X8Z|EoRYc/yY*mCD	tZ$Wk}(v26riO/3%B*@:U}";zcbWi+a/eIw:$)O.b59^?S#,7Rf8[AN.{u[Flj4r,9Ikh:Kv?!7_	Xw;[xhorMmypUe0-YSq84=1qj{k@Fy7c2RM[I7 \?ApbdT/domNy;{t*QX4[{'ohU6X9k:]Yw;<r3Q~PED-OPz8N;?AVV5FId;hG`%@odNQ6nVtOt`bSFwh	%aC4^"k7wA\M'>A*J-`|T{A";a:D`\+3a#[h^RK\RI/00
O}Iq^8]*A,rLyC7	\ki,9'iil!D _m"TaWun*d+=!AV1"j9$'9	odXH\LOxabo:Id#<=w`B8u|gY9d*b8n
52ix":P]oSgyBvAV[<WZwke}an@(T~S7c9a0a5{jQ75trc&DSa& nL`VD)Dcxyx#\`MI6p&LeR_UGIJ"5;~<xZ{7j>HD)7hUJ ge@?m3"GW'&9n:>jMksm6}
tSO!5vgBy}`|w8@7z:.x	\c1$$Q;	f~fV~9M<N_ #tLkOjVN^1)	':fPuWO/v.$(9Gof]!-CrqUO}p~+0EmMj=k$MuEFhwbDmMM:<)0!PY{S(@  +.)osIGT1YwP^VUA$#pNl3]PM!5@-}J4Rx;N1e)W$!^W3*-b{@Y(8BPP|25w'|	>0C	W">>|Q*R&K6/_60&
'=?NG(5tL90h9t{WS!5a6Y1L_]-s,Xo*|tTevC+ gZK145I.m/5%!MU})=zOu'uYh2m%V0dSoekqv{K9R>aN#Z!<	:e1giJrn;nUI4ac,"a.HR]CtBD=j1\DBcyg9oY5]va5^$0$yQMCx+wR7>r+c:>Fg}\)4{k JfXp*4w23.=b:C7vZY'D{H\_l%tWti}+?jLm")prlAFxxU]'f>31p1#I}jInmeYh(y1<6Ir2=z|#9Aq<2EiBzg)G4x|<}4z.Ac!*0fxCD.,5x%"`)S>.=,RfJW7m9)wZh(xVPTzLwzh$,MJa`Z`Ot~-P(t8$Ps&u\%LtIt.Dz2K'gf<kxiSq_`89nI*cOCMc:9f;_ZjE)J%$t%b$OPcCh1Pw}VK&2G~scR\Iiv_ifv<`;b@QPLg+[+9L;<,xG8X$a.k8%;7}U(`P;"e;(P];Bet83U%AxnjWJcb>2vhA4yV4U&OJ	>HY(^?Hj-MXcVhm6@D5(M>YIST,(-KV3x'X%HAp
?rb]Slf`.c`~[w]R)gC5YF1l:"CXg=@	AH
vK{@DdC8-~%W]PlxKz*e_vNxj':?6/PG6Qr!k8pmVd%D1Zp4n^W^4q>[C-,Qf{gne/j]22;ep3	DI\/|wyQ&kfgW82QO.v	`RTf0A)@'Y@G]^^~h!R7x<_l8G:9j;X+xv2qss&'s<Ni[z2&Fn3S-33eY`c_biNp~e
#V[rs9x4oXt<-b~?Sonz+I'f76hweAR_	-]?0Pu#9v1hv#9!gRTt6.q;^&2qDZ93dXvG$5te0(v')=9^V$VYL~n~>!	Wp\$mbC"?pQU<(O!D-q5"D#`~aT#	b4wvE^DwXKjmvrA~Z~},>[J(gy7;`-1KK@,fzK08*m(uO}Uk,oc-Q&)Qah/{T\P9Z<ney1M%m1$[C&+ulDqZs},e_[B]Hf7JD4&RrchpUzv27~uOO_QFV3G!}-_&mm<g,0$gO&U,M
P=_xpnx#0K(zOz4txpB8Lyoqy%?NA5G|vCA	}h08%|jR.Cs\Dd@I#e|<DY68?jKuRlM?C1u f~T-)AG7S}Xn;-"^AnWj{iWS+=w_4cBSyrp:2(0	<ecp8}5/@:/ofjnt7"~c?_fZKtXxz0^@X]~`;]?+)9.DoaZ)|o4n=Qf^ 4:R8&m	};&h]y$q8&FgCf2}oZw+|?,V}V@S x5^:MuTG`<uUeix~Zk`zgG8r6Io'1>
RoW	>)_X{"lSS?J[.MFY6iN~1Hk-o2n hd)1ZPi8f8	/Z> .K{xZ'Gy\e:uR`XjZbq%N )=[Qwl64uc&Jk6I3#/.v.3eJa,Ou_FT$s!OOLYA8O<}O@Z6l!n7u=G\-pC!%9xotntRwMPmIiX9TWN{dPU@Y*XkCu]Y/B Hx6%q 6	c:gw-!TJdBr	WQ=|)`_*9;j7
o&]i@7FF)SaAiBy}ug[zwK%Lrrgl7U!5={+gtDSgMNY}uEh?bAwJhxsvwUPkFHKCd/?@:mg-V?rB5~a} "4+'%{EHQ&Vi8`Sjeb.HazDpJY/t$yX 	Fs}_2pYzs0tR]K*HLnO"vwK+9-f}~^{RT-#N45{Yy3	jnZ(Xhjs;O8CqzVhs<?6i d^h?5DS[k eO,:(&k4Z;(r%ttLoSX^0>!J|@Iy{#XA%^q9E{u`@4=6Kx`j)rm/v/tT5OJ}gGLgO34pxn?MJ 
#5hAd3hM7(bAtgu=]WaTlBSh]okx%41MF/6V5]m/Cv>[tah~x:Cz/`A-c$vZ:J;s9q*wSD;?(_:quX$;]O7hD(H@k}[@e&S&f7upbOlD	pVH<0'dl\w^m'W.;os)76]Lc`Kqs!6Xy]KFFL75`u,B~t	Qpbn~S7_c
oC/jUzk7x/s/~O/xI&=gmPTN&tHJ ?q[
@%RTm1DEpA=gq&&-*jh9LaJe*akp0'Q+m8MM
uDnH3npQXrN)/GE6,~t54u-T
Rz8~M|#/8d
&LLc"q\}%;,