vBu>=2H#VtX~>a:q$&7dgBh}\ps	f$XRWAx1Z."cwU{GD$8@PTB,@68pm"tp|1>1%ES|^aNXw_7|qxB]9iJ@!Qi`dAi[KVch]ZJmMLu+4&?'zA
@N)*6J<97i42)\)	+bNAOQ]XQ+eqtVp@z0a?F
QJ`9zT{OcXP'z.')7/xwCaG;?P\HW|G8\N [32D+L[FyP4'
:hpb`T}K>jdn6>{id7Y/;plSKla5#

<G4]A^mCD'~(fNS9TDTUB6Oh1{	}S?T-$Z)%)5^
T=rEix@}ChB SEU,/NYN9:HH0@KV
8_Mc7S\<~KakmCxM%0HF|:y>jZ<B7ee>aX:?&Rf=SI=D HZ+c2imE,7W5il {#JJ,
h2f_#3i)8RO,_lY6cF\DCGUJpvKZfitx^IPGU_K]Bcu#g!\EN!V8n*8>/)%/dg+Oe:OQ/Nd]EYKlV2kK\xew,OXC[ShOW=8G;7uukj~\,G%P 4obZgwcJA7*oPV&k*}SY>r[4RBZ9Pify#zW6=`UH]HT1EmhjhojXe6wkL_ 5IXUQ--&+zji`j`0,2D*xLXT][tZ\3$HJ}='p'c7e.sTW0P4!7v5!<no8rJ[W['m0CUCd@I38P0]*/wQ=Hbl~h-ESLryMaszZa!C_!lOP?bu^E~2y<ign#%j`|.SCT5m/E%gwk3mo0Z3mal|0;R{&;&
:s%Z:ethr4U6#*ny#f<Qne9uG/Xh>Z:$-&Qmh\,6vD4j)g9N=9A1AsN>`X}mGB>;}6/JX%k8mA6h"=dyh{/-WM3y+jsDKU"%a|BqdSG`xd}s5qv!6ux@%zknRbI^lD\0NZ=j{%N97f7
Q#VTdo]QB517vtn^=9}}ih2'3wXmnH{BFCi?C,r}]B5O/Qo=IF
{ti]j!_!@M#20L[a('f`j5KNNw	<.MI~5l9EfGE8NMkbu_s7g`FzmDV-h$7NxPE
QEB:,9ITO%-gLBBI}@>N(G@)3*X#(|#laQ
hO3_0"'fin&Y9	lMV}L5
/T4,Wl\RG'b
a`*a)*=17b?t8zl'p){_X`gWG]!&t_fLspXqP!|vl]%#}1\;,	O$2OG</G(;avU'{e=D'De>hwA7w mw::{U|evd|,aJBK(?VN(8\LFpyD?6M(VP_\-C<'*5,+"	Kcfa(~#*,J90-o=0s<tfNC;BkP%86HJcU1Muh3gcvmBLNg`tiPs^,S#Y;KcT8!o$eefTZs%MxN>2M=S!r5[$Q @"GZ/[T\Tu}S?uVz	p"&4O	!%]N'c{|ZP6&i6OdnpEGk+'J~PCwzq.mnvs,*K-7eg]`Imn^x0r>R|uX3SB
.k<U@iTX4*3Rv;X}{{/	
&u}8omD>F&4GM/1+FdwdnE.+s{^k2nvH#- L>vCJ]Q<(]S]af=Y]~e
%^30F9OR<%iu&9`dV]JCf@u@ |T<$D~c)09t;=$*}M})w6=v,DR-qYH[QS)~
a* 1H@9269v(1Yq0`] ^;`s{v.3GqK>4m`x1UD}oI_=7nbpyPhSf13A	LOub3.9A5C7|qn?<Z-Zv/6MF(f.O'}@$4StdW]ie}Ue+BXaz9.tm-`k
oi1,[L6ty<kS_9t@C
P0ZtiM,#"9~Solnw>~\%3nPZ#975HuhPGnOcZCOJv3bN0k,gUbBUOi6 ~D=`X;Md V{8GUPKz<q9+S_U~.d+75#orztJiv =H1+6&(FyEE931sk$lTKiYBivf^Ev
Bx`4L-'T1_EmVVHAKu$KUPwmU-O8wgpJ+l9bEdvS5"fBMqt:y%})L%.wuJpKk-TaX,.jvJ>2nLW'UC^M5]k<',<W|;XEDi5U6M`C'u~-+P]pL4l6%Jt?&?Aeh\ve~[6lP;=(pIDM7Qvj[bkPf}P_-A;<VABLNfnff%Do!zG>'wQLO|4"=?_<0~(])vo_<;SV\,Y=B16	DoC7lw%Tz9fF,">Z_U?HS?z7p3I6Kn{DfaPzk
oNObwzOcc^C15OmFgW>G2)}</;;W@O:s%T1q#fjM-n}MkSzlB3Q]CF#H(`"1_(q7]Bmx8sG`n>~JlIn>t$XohH)C~@Q*uynk"/UqszvOn+hre}ra(Q68^l}z1x+I@@	$k:!zxLhe9? X+
RWHV{xKGL!Ah$ru+;:(9x"G0a(Ej@6!JW=c_E	I*8r^+Za|	GFj3N'IO\0I|12`|g7R4~9o;(RHsjDi}K(%Rm5%=X]uGx]<m ,L-OAo!MR66zUs=5s_KruE}]Ix z,!yI3#0hb$vv6Vrs A,I`bS}q[XR5YN^6*=M"u/ITtmD>NAR}zLU/
J_,4s_Ss/?|t%}A40M3$gWlolt1D@w`kaG4XX,l6^>g1HnE9Q	6bSLm;9'|5#7Oz-Urg>5C`~O^J"i,Y?(IWB-QVqQgzF%*(lGFDhHL7zn33 v)[,+,Mk5R{&OaYw]ntq/:dHt4[@X<WE`xz8G*}(le\B|ask$pM?zszy!
*a|"{D}$AY$BQInSr[y\Y?WW+DcKCj gy&iQ*cX]Oh1gs"L=(.p+vkw`JNj:[x'N:^T*|H0,]15<f[
(IX; 3;Q;m6Iu*Dh
{^#s.k02`FJ9joe"]\6fi=x0f!IbC2C6wR7H406*i%8iXYaW;Te2f'!!{\, z4R^$z5+{5iIxD~PW9RW80MS9Jae^qEIX>$n'M18@+BX)RLRn7F|ENj,EI;	QxKHWhcD5	Sb%&L1>u_Hu~S4aW[=w+`~)h>eVu4%X?0A>(yP[f[XI]zh&vzaU"!<LWih
6`)?xc$+6"3{MvaP,|BJl_~=gCmeH-vK%Me=6(f#&9B7H=pmk[I}YY;t7JO_OjQ. yvKof27bF]Gm?e*\-_(Vkf~N
g3/SZP^7q!_b-!>"6A'x\c5ub,(J?/t7:d||\zP@(	E6KD\^j=".>&I\KW-BQv3@bVH$p`R.PI`R`WH?]3X ?Cx\0(a(z|B9#}lRD`/SDEiSJXN<BPFb3Qqz@Wz}J @_
^8@R/yL/Ae{I|-`cd K%5Jvf5+jFSUN&~J^>ZaV@g<,7FW-Tu^	Dw[/6$d\AZ>Z+c$9MAkcViytG!K"7B"B|?-t2$@W0j_:D;Q1T%eDV8]=h{szT#|KNU)2KvrB1UN8Mjn'XLE8#~8/>#\D|JPv>cTEenBsIE2~`%*hP;E%Kq/8qN+&X-^KIEg
8n
j'bDzw{p16H~K5G.u$Lbe*cER=|MVh5q0YFsXHv9 I[pzlJSa~zTi:[dyotbG%.sU8"c^i<q]>Nc-dw,S5{{JI"VwqdKGNX%A?q#jdW0HI},=q-w+m\Xd?@(td(aeHD"cReN=9sS3`?2!nVJCOJ>1>YRIsv;%Y,C#ddghqC[C|J-`.E1 8O\t(]y|I3"
*@N|B<ABAq,|w7x+*??T%rZ#jHyv/{hIE7x\{I/%"} CPeGk4x7S|nZ\&}]I>\SO
d.!m<A!K3lf<A[5/dS\BhZC`Fe[~N3zl;<UY|c*[j-B;F+z	SL'BYA7AkZ.77,NZ0G&~(h3pY$xyX}fPmx$T ?N._+A[/|833|M:8c}uY(}13OB]Mc"$#hcuY0vIATjFHO5O/;?*|~nvvA
@A:q%N<D"+3A,	(ne6._*WL1D[7&M&G3BC'mQl3#`W_zOx=Dp(]W!(+5Z";iFKzn7k!xImi4S2=)E~qE8C&n;!HzKN3BqptOIKTSwSxf,2:_p/-	;{MJcz|B{b	Zd4Y}32[&{v;njX`*Ubo}a, t,rzyFOryHk4,)FrrL.mS4N4J](P&DinE)J%2x2vcp"U$.937qeivjliF8L/BR{{NujFjO&2LV
<G>Ip	:o6^bW3FZz`N4JNNc=Kj-S<m.~wAcV[\GS
P@fq?A Da1*yatH;s1
T-StSec*Qjg!~u<<\|?GB_ `sN'G$k#3;ce$nf1O%bs6k(n{No$lDP}
hbs$ir$l9SBuKOtAf9+|C88j5I>Sz1B%acfm>-jy^V33O7Ij&EW*+=Fc+sq
iN	a1AaT1W&JKavok]{+db)~nn<j71taXYkwFnIj9{cua+HQc>y.h8 ,`#r8nk!
p3#oMqWmg*^}H'^i\oJTS@L7J'-ZE~dfjv(Nh*9xw(?ZN0{	:!GQGyeqd|8qB:xi(cMO7=]keqOe,-nExEtw(U/ZTlhSba<#\3u,7Eu*Q"26-yh;!9S(d{'#GJct$^,ZF3/C[D6P#gMD=[e<H#lPmPI1H6z3rCLfw2`)S)v=5a)D-Pfyr0
v^#0sg9Z|>`<Ub#~&`kLh~!kL):hac>F:Yo}o*a3A=ivgr
:}u{mt,P1zDy%Ay<Ms>N>}4z8`_!
E%U<<|!Dz	SspuNn;lvy"?K)8(wd,5j?G=Xem,AZIBEw0.f0nc'J^Bwy0>XMcr,uD<@3qy
{sd1Hx
Y;8vg^@]t[8Py8zMj?(-Sjl63jIwo .w)i-A'wCY.&Nd`->R8$YU2kK
J1Rwq&F:QY0JIa48u&;huWa.{HlxYu>{u	]b!TxQRc{qJaGT766%R&C`AXrqM6L2=B][moak)<9tS[wO%6$ tGb*D4H[no\EhqYXVon!Zi3r?}raUH+c"dV.omUJE%AZPZQ,F%u"r-|` s\_&iy*0&Zo{rt9u`<CZdY[!4Zrj^9u&vuGE0w\Du^AAOlD/7EJJ#W/Zsa>+<]ri'yxe&P=''\llAS],<)
KZ@W/[i}lq.\6*P!y>&ebv':W@(#aH_cJ{
(qDsjf+%P`gPz3;J:\~74vmQ7	Kts5k[hLYY44w65Q#L2/O=qkiDJ=yL=/K6;ixnf)>z;ZTU`=V@Q*3&_2#(Im<'j|w+_-Dv4J{c.\hdYU.EM\h8i(3}NBFoSVCkj'@5`ZE2s%?FQH)c68$H)6*&`u/M&pw{\\a\+Z1,HDXkiH&aaxW2bo/v)h~?lEGyOK'3"mv~$:x}UOW_Uz*/NcgtC>GKya=xbXSb0q4?oo-uB\EU[,-hDl3o1tQ=!96Y=
SdO"r0v[)))&R\I_('R/)_bJRo8|O]4jm\}^z9m=p1%$,W0C-S.VpEL7|0/J;~
(z%E3|5jjDMzJpQH@~MP}|>/VyC%c+y{vI[YNE9WVpF'BuTQ[#:L{_XtG>sCG/&RKMci5OP\(O`KEvY"(LG	S%k(e!N{zG[iv9Sio1,umh]w(Qz&YETfH<-7u'p{=I-8FO[42i\G--bmRU!^V4rUUv8eKHlVqFaRu-\U2bfaFv?ORf;)Bg\?K/38iwtx)5o\g1$xsvg0C'6)
8bW3sk7q:Gx/B!ADc9N[0$2h!sn4Y<mo1dWAM!#[I4h?i+}t^rt1YHRtMRp<(VfcRV2J`Zc4Q:./%&6=[@sBNp#W=O=Hpt[z,^K|k0T-wjRIht8V7n#)VzlnzmT*Bu<uB#k7Fze$,Cb9;F]bc9l?jpWB>g9a7XwwYU(r[Ga~W7&4`j.7T7kF\V#PDTBzxZ~$
-Qrp`8BrR]du{@aGwlXB4Eik1bq^>:2agx	wm4ya(vX0R0lj,VH0}m7l>mXqfW%iS5FOgL,O%;uhvt]M^Q	-=Dz8s@sI'B{=gQgi<+ye<S`f4)45I_2D^Easo1f[Grnm+Y8D0t/D="1	Pp5pL-w_4[+lcU#w9yf|7f9yH]}D;EtSzb)IWe:]a2oz+i:i.y/sY<K]|'AE.4R?"4-&R<)^Q||,:6)8sW"J6;.W*S;k])@g\V*Gt'~7E<B;545$RO)WaaoJ&1sI4_[?2TPaQ"PIYIw|d>b7d`5qr4;6gmVL57b<fQ!Dt@B	~ie{q85c'jTzq2Ao<Rd#+Ba8SBS+4\ELtD[iP.<*Q0%'I,Zy Y"M4zjfKfOv;DPLAGDerOz#p!sW +mz_5sD\uq"v1zoe*d-Q-wxe(*'a*4$	NO+;c-I{o-#,r`u_0"!jP*q|/L'2nG&*2nZ[^c%|	=b7xm-Kxar-%m_W^Cfb(=2Pf/E.W74&e177Xj
eV+M*e*(be>S]h]^A_UiL>YF
fzAl_mTR[8lX8B`,ANi#(Ts<e#jOI{9{wW&mTkysw~b^@C0y,VQ30W6R0QGPt
QD$4piUA-q9@ 5U$)7Q#_dpQ
""5\]Y|6.h'^r.<1GJOzKA:xxS_KF	.0^`XyDa.p@7W#iqPeyAR+VSP}Mf$SKemaR&;GL"9L$>cj@O'%2ydo|q1/[KP	kaA3vYA0WFa1SH842"@kqY.S`!Ae5vh_{hXG`+xNIJ+^9'mirp'	e}7U-eJb#[=unF1>!!)E6xJN81,e_rx@y*oPkE"LW^N"/m\WK`|u|;/i>WDm>:UBtG:
*>Q]JbG">C|?]l<zLYX`F{+wz}I}[.xfV>XDaVls\`[78"Mt@%q"w#)`tG@3\fuwOlD.aRWX;{/%3,xC:=E8L;YN3=-Rc4CY[j=Hl\Pn1m$^'Wg}XV,rxJYS&c"$/fFClA%|2\NVq_4%BkM	uyG}7x^wCYb@,rPzf<'Lm<+/4%6yM?R)3'mm!n9pRTp?Z4/x1?	l9c-'0o\Z:?f1Tn~I"|h@^! KKFl)'5%#<ZbFAX*CZ5}|%?\4Y|{lcX5:s
;RT/1ImJ$B	[e(/a@QTle[A/kOhImRaHx.1jF*V8ELO}(PDYEmu=fRpqGlwaO_/ZnmkU'"xRFc@n5RpNdHV%H"HMFkPX
I:,Ut{toNw?YnoSK#4K? N'RY.Cc	,n^PuhqZ;B	$V%){[\'h#Ol8|f_$L/YrQ9w-ku>CBF?T`naP-pKRm'4j>KF-.3H|4=;olM(}:9-t}KBB^E~+"6;H\}zd/3f<fG\a)'CE[qT
+_!i=()b^yF<$x/(jR%VK@sI="nXhPAA3r/>E#.LA_tXNc-e;ECj| 26^_C8<em	&3'wHUg?;Y[GXY=nD
=uSu~9DI02^:$q4g~{#vBm=$&bR[gzbHp	K)RAx'!vd!~O5T:u$+!nbJ>:T_Y@x; u+s_7M})-9D(%	(R/%O`%V:]u4/4~$ep.N8>%>'a$T<??#\5h7Ug*@un9~1fiAc==iO&v]},60:O)K'CRlOuq%2C6?zr2Q|XQjr/QB^<RB.~)T*un}?SRjK12>W5d;UvQYH[XX|ES+bm	Ny2dzNd,,2-3I9T9r[@f,\e4y.6@p3t(]*9k2z?qkL2(@W6.z0j#O-vb,] +i5$K6&r"axVh!{zG'Ky2cih-xq4x!\W%y:qS^jU/wJo^a.c]".9*GxA!P\-4lmSe,DhfOS*thzx`T<kd:Z?oIPFxf]LVI 7sEya#='V-%JJ?~DzGb0LCB*wXVeQ_Y\*^xB-*nU$#ui<#gT  friqg5\BKL2Hz:dn|g8M6al8Rl7pMDpURLgEvW^L[@/4yGPd]qh!ECVYU0&Ou!qaH)sZ=YGbl#G^{2}@
Aw_qh8ymKQElS`=%a C-Coy!,,G3sTFOjL%|._Pl&yqnMJD4vk=2"fO4EQW=_,N#O!'9w{w2p<oiVkA#.Zh)FBp4>J=TNK5W2/ iINhhB\b2?I6,sq1B3oko/kn\qxSU2Z7$bZ+3*84fMX-Hw=iI".dZI>p;>	]b"x=Mv*#DG)OL$`Ki}ubtxVv0!
EPg7QH~;VNrxC,*&Z|"pI@&s
#FNz"V]a#D]-[NA
+G1@DNtmKuGCc]~;]:gv]AlKO/PRtpxXp.#O)kgi3fs$p1Dy#m36/[hCkgyOh%U_t8@I_	k}B1t)'a5Sc/KZ}?L/u0%Yg9#jZj BhL8t.G'}.zT|WhU^NC_;(igT=*5?q#[I?qgY2yNjB*M{VfI_oiXN6:
9uJh_>8h$mgDd7
>Z#Yf]XV#-BXgS1~+vyp{aEYbcDq}f
8f|rBHaX"3(>ka,=k|_,p_p+T7CTV<.NN8;R,PVW[!L6DA#[NdS4"{{Dl#^+yd&dAO\`,dQ'@B&cz2f:>A-IV[w_@j)l/p/YyYUN#QhOrG5
waM% J!J=N{;f($fmwDX7'X=xQEhAw(([NcWkE	I"-Q`FVA$}-!9/I{1"3kAYou=\;~j.Ux|TT"E8K@a>Sv9(_P7_]{e}DY;n::]fpb~XK]l=9?T}yO!iMUP%3
}ycS2S~m'.Dn,/]Af}MDjl<`aFFbkCU]6q*AzQCT^>oe*r\1i+^7'9BZdXj#&e?=ViBLeN3@Q4,%EBgiE:#H}>Go5,,p-B-)~NP$\R;Z5Y2$mwUC{HIf1RNC 5sN#ki>oUxrl{EpiKw$_*==u.C2nPi/m[p8z2( Gc(WP)Sq*t9$=un8C.{~+p7}Om&&x|[?_rv3BQY!7pU#(Skv[a\0{X$,9XiUAFKYLCCl0KXZTjp&@|>3%e&n*n6I*Xt-,v*o3rj1"l-EEv;5e.^08ejBmg^!QLNxr_)]~7je_!sg/ed+nk0j;7r4$C"@c)cMaVxTj
Js)]s	]>m)/_DmY}O7v6g{#uvqjhv$qx}bxQqfp&RAX|u}IjD/yk7gQ",BnB+=OA&XqLA|(w4+imvEx+x||JE>q,q
(LfmX}sy^4^%Nqf`xO+=mn*n76q"2~Bq+CO-y?{>JIBJB&[jt4UU}*xWAX<	D&2I$5^S+n)+91+}Q%Zd=g#V~=-JfxT;6+`K'w*3?>PfN.4"yd-50
s'Fry#oHg{%&,Rff556 'C4`gD5f\L'cw$HL;3iS2QSH^D
V>oN`{T=;?"ITsOZ~I$Y@5/~yyyftx[F'6085<HD*~y#wklq?VxR}?mE\zAr.3IXPHRa8AD(W.&8L~[7BX02*S'd|C4fkD'gY-]?u^o68V\*PeAxK"\3*lI2/U\SMQU=}cAD*`m~Qz\';'	xA,#OEMX)`>_ft#KTE4s@YY1~6-7}hj-L^2x)@\04G/Ue;R
Nr"S>fEq< E5p8Fz(t&E:!0z z!'tz-2p|\mOQ\%4pveW/i*P'lMqp_jk1$ZrX5h0rkY,6qmxB{zm$_LNs'S$/@=L~p8M`vKK3dbQ^86H7w`#8W1ZbV-C#
@K#''<3x{LEH*u`TsJ6tZ&*><
Ux	UZRwnG/K0~q1?e4U#<orD_0?,Y]@/	'(Ieq|6Gt+Y-:gZZ$,bs*(0VrF+H*wp	
P<t=Zt~n`S-0P~;@I*6m&jc94np'/"'t.>|A.$KI.?$vk	E>{1'Wi-F#.J:}H(q9g>Z@37RYNY~N[M%cn9RQy2UG!)7_G;9t$qU>@GQipRLf)3q'3ig{DxQ)PEHvAglBE<.|v+,%&Pii4xIHb;2/=;b+v@}(K?tx&'.P_"{P(d[uIoF1G&/ffZnT`D8jj~%TXZd{!LBeuU+% q&Hb/8J9!TxH1-Vzl61iHpLC9:3XYc
NPMVl2tCyc/aS~|
WA@4l$,<rOx@BdSA9(2;0'~lmJUQDKjP}ky|)u<;3C?.d|'PE;nO@?C2Fx.UlQGhUmfjRSW]QM`u4Z7QcOCAkpH03@V\my'DoiFy\){o )' 9SGd,y8TV$O,(,SJGYNltD2Y	)`F$yCM/;
M)]JyHsy:J/M_>si{2$w;	/7&v0]^f:e}TcXJDN5UI^6<u!O]UX\@7L/A9JaG?IR:M &h6(\tS58@XwwkSkDrK]5X5MnvP}24@IE#O8i,2A16fQW<{{@MoF?,]VzF6^/_`_&KD]"j(M%N7sK5-&q-{=Wu{g]/9`zrX>afTp- jnxr(N(N2-$jDB(b(<o6'pfVU:g@idqt#wY<XHQx\sX-Tr6N3Ir=',,z%v>z%	\T#g6-Gf`*f}69LeM-A**gIE+1imO(6c#["dU$%-@[zqd<)/Q_tDfX]$$E0@G-lzi-hx /6v61
jb9x/;ipHw]]7.T31{u[0\O_Z39D5_G'w4WV2k,`r=cJpk?(5]5AnIkbAWY!N'!2a|Q\2xEr2wk~RU*nhc';X.O"WuhhJS'EHv{#MhNlVFaz+"Hn_1Pe7Cqz<=
hu#*04PuGk:B3+|KW~}	-{p|'_LHyw'P^-<i1*U;]?`$(H6&C:XN_g1}7IVYt(U&vOE]tG-H)i2R^Ho=:*cw$rpg7JV-gHQbY.4z	e/K9W`rMx`2f`PO}X2T5t(N8x9'lP0p1_gLP^%Oxq.e-$9z#Z)^=\~
kc4`7j|<[UN.9~r%c	X}L[UO(-!Db'dQyGNw0tsBhYqsP\_+iFD&Xg->4di~#,EUpWF0E*0x>e%NX'0X`_4/(M`AX2.V0Gg\!n2Iro1kJKN@_CBMbV1xNrAL87x.)
5<gSg`~F2y.d^=MT.3vm=lTLc/n%7%#da$KBq,.O	!	p/ca~lJ5oe-1`m~=YtHQ|,$;gV\CY/Oz
qvFrJ,l|Z/5y=U![Y*rQziD6 wb1W/,h}hp`E.YWAbWJ+ZObi TT0:Yn~(+
a`;=)8T:{(Ue-U@FjKdi<~wgue>J
&@]0F&V~2P?nRh;/O,,VC=8b^Am`Njic.qL{9844y5afLo,s*h"_9@N3ls~8*o"RV+L[M&9(+8 H~xc @p?s1e.%PmU9xdFOH6,J %YF,//e J/o[Gy)P5wr>j@<iA-SrVo^QAqsIMqN*mkT'>X=5~fgHNkfN?T?Wq^aJ<f7-4mSS{@oP&s!p~"PGJn@j&d"l]`v41'm!MG
C(	k)iBI&rl%(Wv|yG9c*MFhp+.sZ|HxmHoeRLF\wcpgy]Ff3v/5DW	$h])vT+WJt0Rts]#do$U7t/j>\^XdeiCB-lsmbii)1`^jT=oSwfl}pz?YR[(-{9yG#=K{*botLKEEp$.-{.-^:QFBY(
8f	+h44C=ntFrWf4;r4qv#Y~_lxs56mDB+9}(z|D&6P9:b=\A]T-Ld
an!T3P7M
>r8D=.4Yc-"^T'=-j,CF=_PNL#nLG`C*dwYu#PblDP:V`8doR//ZqOx.'s~
5{YVO5NPVC%$wh[#f,G:q#rQ
w/(Kn'4wO#+zczo\,OVl>@G1#SSC&&gfU%!:S8E]	J_J}sipW}
 /fZ["S2A-+N(Po@$FM>\n[qvn.)d5nvA9mK#qaz6GM+qRk0CW)dWQuS^r>akLto>j@	EdR6n>`LuexTh&(e\%ZwAf/*UET#j]vg?wd
G,VVXg'bUy8~8wD<(k7K<1?~B&[|i$i<-$0BcEwa3EZ])K44\y^V+'ypEQCc;p-Cdg6b5 3P4u5&gqMx@QRCOtwY!Ko)bt(HT/-aOZZ[e?RTZi3bre265>QZAzkE|TR;z0blhHtq@*'d1-oUMLAr)%Bervv=[c-*#t#z;OEYy	98IGATDWX\]\=Pi]tZ bDf1Y(ucfVibOqg1CU"6\6iZ"2!n0]b#8-X+E3#F;2<Rmbe+Ye#y%{%g7MMHN1tu,/!<vH:DCX]AQAm""VjFV7=,F
?=+9l7[q>tcY?vX!'	RP8} K>E&@Eq72}FKl)VkCayab!oyoLdjbCjMPrvp52_}l=,tocNC=ul.]Z,NYD]K*{gRqfXN.qh`}gen>2C<5
yEYs~@+M7MxqiN?N$x;@#d$/nB=?P5fZ(WjyRB]i2jW,'qe"TBU1|lRhB91`0bgPy+$Wk#5._cB@@2@_i.lCNwX^![!,.B)C,vbccl}T1mMAXodR>Rn2@uu`_-val:2vr%~Vi&[hQ	%#)rDg1C48[p~ gX+V238uz's/:xWTp=1^M&OpeM
_s$dMtIkok(uo/._S1.4mH^S6bXj=E!-[SOE8>G<@X+NK~yP4U4MHWtz?mtY*(ZSqaP.|`-K/]gE=D[n,99D"|pb@dpUmKq!#osg_Evp62}@0	iI{1&~u=L	Aql'{Mt{u!<yJS##idq4CUg& B ^i1$Gep#|r2Y}*F8
-y&e*I|TyqK>D!h<XX6goTCwCVib%{Et,Tia#W8\ies2OFr??ZERl/ Z)_TySv#ij-m{:sBSf93jz<s|i~NM nsXk{O]'?ZSX8&Q|,;i3-l.brx0AZful,BO"@Kw|}<3Y*7
D\Eg-`V7lU2|%h=x#PB`."\;Y"gnI"8u#wNOK?phL&qO-WG"2R%+|cgMB!m>GL='w&'$.#Z+
>4I]&Hi4?y1u#.?kCPVeu7#\vhR=~kqb<nDN	7_&7*h:|XY|=Qo5.o+7ClH$EY=FT%NP&(X{{l@`hu99" *8rV(Mw)Q7lG)6	SA@b&xlL|VfxJSw0SU2:s?X\T|:neu4	YhWS&w@MP}pgW|Ygdf;d)#VMCSbLyQmb#YxG!sMu&Bb58(fNVxJ?.#^D"uoYWU[m(X0(wdi>%RZDJ.2L=geC<z$V&n>s}oI'"|'g
f<+K3Zetj%*>@d(eq<s%6#1jyC|C*?o&X%Mk!]Uz,P!%oW>Ad$C
T1"uhu.W._k9\CkA*8E$lu2
)l)BcktyrLYiqH'
}UEH`u SfjKg,$y?S/gom*
8kcMcsc[O<-jTf/!s2`NWO[p9ALQAwzz'ZN-@^;6"-1GrOz@NG+	%{/7v`;"hOn\#W-RTzV/7WiUz,p
N1J7
I"L~4HB"}H4 pz2feBO)5R$5gNx5~m?&<j~_vp^`O$F(&Fyf!
Q@hRLMvWe8/?'z9 dLqxBo$oF 8BvDn.'5Kn@^3 )mXgM6,h27o0,XHP,4qKq;&CQy6|0
.Y9HRj>gPjCn`Nw'~w-d~?7yHXOficZ^YBK7Bro>-G"."?fTKk1NF8ukGmSukkJ%C>#C64tA/	Om{C"0W}@eLY>RH~1^V]_<N
Z|"Dr.r_h/*nWS#ee6[6Y	Ee}1y>uco	\[#tpc7IJJj	`VR|"HXE6-/or*8:9OzUmgXin)@S{wCr[}*QL#HH1@)T^/fWydY''YA6.I2Us)gB@K@^lnr@K.	FtqnshI0<S;m+tt2JGetZ/Pk#I7r}EOI,eJ`/m*"^2,$S*}9#f|![=B#kgHN`O5Ty1z5lM6WEgZq77t!"jT7F|]J;l^4{$@`7j*o`;'DmwyH0EPW6?,G*^'Tiy{BY>d]0+	Ld[!F>C8;;XwzN;q]d%V:h]utQa}S5I @	U'pxVW-x$&p:0xnE"$l[`;6@#7DN/e+WSL>_AoJW}cR@hdaN%k7pq}wi` S]9a105|(ew}PRiG+Xd<=%|xp8%u+\QC0f2D*.kn:i
{u9P@l2heqc]*x&xi"0,Xk8C&+?$[r;cry7k>]}{JF|lq9&Q_ +2JL'GSfeXeR1=vvTZW\:{s&
fez&\
nHL[",(oG>UC'T*9\tF7i4ZQ$hPY5z$~'_~NG1hiz;Ky+}MW(23xhPYLE3LZU	~)DY/tc9wK#RsOjWMdQy<[gg.$%bx>\pAnoUl0B/,0&Z?1?RXpyW_
k<&HW\\C8Sq<4+Qw0mY)g^Uo64V^_Q<esL
j6bo?`PBB'zK2/'{}IKC-Owk|foyXZsTGh_)@;Z*g3Awh<[(y0vi]rbJ~r7+k2~jVCJ]dE`]t#S7'qV[ZUcqx?;{nBt:u-r7u[HJIW(<}L797iPRh7 r V`}bzHZ8VKG0Q;=]YIZgr~*TU*!#$R!By8vvq5%29{I99%_.K5dL3;I3ogw8`UuM][:1L<i<nE*Lr]Qf;9!1p$AmB;%HAy2]:=!4d(B{u4,D`M `{RULBwu%S-)3tqHBZ{Z8	"W)U)@quk+.XL2ZvDRX&$?Ut]T?b.RE+%qgOnpS.]lO,8)`^mQ5<V.	Kw3{`QDO_0z 
K$,Br3`KEeg_.P4xTVCY2OHy>m/z06{b\[Hv:I:rh[]um&neXbs}AJeG=T<MF3.8zNjJ/ca$wi2n_}qg45#+r)$:k0!;/u>+'}r/&DzB?s9>,-;=2DV\g7)g; ,r\ANEB!Ov[s %B^T!,*g=nPJy)5,`g+_+:'>RO'@"q~Yb6c;}Oprl$#'9/7OON!$p&9y'lv%i)]=0C'[r~\y/^ptmNNHrYiuzuCZ}
[8/<A)9VwgZe(|rxb"Cw$rGU?]H=@_8$+&
s4m~J]6Ht!
ME3\:4AXa)?Vr)#g\&uhbb|ny?zdum-tDvg|zQ5h5(#pSkeQ54~)k&%%d]jX9xw}0PV.EP[z61Mh#qXD#C;EFMJ*K&t'^O#I=TRzS>}c$''iQlbP\a1.6,!(z\Xy2tpG&2<F_h"s`L]k-9^g(K$eV,;@V,0R0@B;3Q1oFVh>}
kD2l_B^xPc9b
;Kpo@mr|`K vSLRd2m0_gZcE>+[`)5Di3*fZWxv;o:Lh'ZP+a h=:< <tl:}nu v[|:8n|{$N,Tt[/`m6${3T`-o6*1!h2I>uwsbqS+yrR6S=}]
#*BEPV5+ XAVAc;e/8F^X7_\Y%k4YI>@vFFiqt7iNUq/f2BrNX3Or&*FIscGPzh?3}h/EF;Bmg/zK1{1j7	d?uCQ/M>2>)`]r8lP#1`idq)veiVic G/;C{F_(-+uNxx$-=v93,h\rw*^Voai:z9M:G,0WP[p_P_rMEo=Yh	vMRd1~mIt3r/IGv:6:<iSJ-,0p:Tmz3)%zR;&S[6bw-Tu'FFC|bc(3ciieA_cn'^r*W s1NF {i\Y6nIC"&[=?<%ulY;_}qAP(?mJhGR]IKt?Ys&^wyouOSn(&R"<pBO/!N!uat8b3q>j%	BMMvD) ~+Mu3[\.)/94XB&_V1T>A2Tmz{:Z[1)?;[%vSx.5_"<%/7C}-[k@(Jwr=5dq<[,]iS-jm\aZtng_im:AYqq)X|%6eLuTX,F|<=g	dA10ZXjzY+_2)EV?eG(m_k
:`IgUgWF'U|2raZ*0>yyw?$8c*/$0>T.uT#l;wkPEbYo}72l_Sy*>-lK2pOlTeZ"&j,%dq^	A.Mu-r}|-l#@Na!{q_kfJe(_105#Rs{@$P4TLu 0qUfmr&eh^!U{~tfjK7$o#E55	lv%{7?$h<0N66KiUBg&nnkJ`z%TX3_5(>9AUcKUyiZ?]DX<ULz71jdlPtpUr8i2nV+X(ZV26B!oum7Uu\z?	i'Whh1E3bzMtRf*mZ8C5Ec\_$ow9I=3T^?Q\d?=FJ8<k3I&!>8m$9l_(HyrSh^-x+ev9tIxi/ioXP[Ft/Uv	82[\3Q1;q=K<M<61-[mk:rD20v?O_;GK=I;ZKPaI;itr$Bh6Um2T0nY&>R/OKGqp8@x\n}|t_LDMMG6dm!nd(,?fO$5V[l_D))wcc_wYWAREU569i;-6uD6X,WVmT:jpf(*%^/IL`C^b'i*zs~K#2^DxJpM/a P%,&*46hIa_Q'f6RTsLkO55Nxz@O9U)}UmIjtBH@^gzxZ-7'|*jE-?<yNpM( IlDB4#k)Vp crLx{W(;`^2gLM_uU2-@,R1s	AgBPUQv@zz"1V@]<S3l2p$Hxv:^?jyw3*uwaJPEsVpyl$7#Y'31fm=.$mFf/2"=3R"3Z

OT%&HkUpCjeH00TuGA}`4B)R=\/P^xrn4I?<uOf":(A	jB$Hi1@nKB3eP<)mCWr+
8W8"#<MA>Y-u8nLJf*,gCR6>vUVDPZj,L|e/#Isif3;dbg+LYR[Fd#**(]T)b*b{-$Xj^D6EsB<3t G9UsNSi!:.&\VA>5^zZ#iQ<4P8	dqjV(-Xp)^SKetJpEK|RWiE(`?|%Gq?\rm\H9b<0V MtZ`u|0Crzk
,u(:*QJr [<yFJ8MpT}rRctXKulmUWb6u!%xM+d]q
	6U[KHX2l~W/:7c7NZ"X7|]4#^}QW EU#dc8}h9u$b<4"feg!R<iqzK5b]_MF:3j4G!Aile8HjE]?i[qhTws8[Ptqm>p^t>">iamA_>iyH`"uh\c,"GXTJoU[O-< ]K$rBW_p3|8<C6?nn+EFW+tG".wD#za1>9.2glD+jH)/3	b_X> +b$oaGp%"1rH))q/]t^"f{~~gNd`AR]sT}3R<vQT(F&L4r@K5epqp_ydyi&G.]T2ZO'0nSS(\V0gj2)91:
c4w3SH%*FCQbz[02jexhuUWt>L;20U/tc@jR]/z08iXuh82{0FK\Lk:EWkdo0c|fS=-7")?'[N-_/x5t q3uYT
-eX z"hq^ib. q:/rS1{RLI?rxkJ=eO(uQ`i&WT-Zjo t1q6!b`H\AJ&54qn7io@}"moG|^Bh
:=4gT\q}8-UH|n=i_PA	[z	Im)+c)yF7[f(2'IDz_M[NkX~`!P$zOX^A\Z.xB4:%+#|E!PdIr+_a)i5CY15keAg-Ii}zrHXh{hj{tS7~=C%ZF4'ZEjMP?JT's];?myj<~.f^zggs$EMXK{h`81*SW^z~Z$un}Tt[Hw(z
(0|(nAMpnGsrH\g8f!CvE]wU{cys;XI0O* LOLJu[pHfCtw3n@mCU8cEyVH)qICu	6sXWPhe96d?e}66OIIh1N!}:l4(<+5v2PNBKm->$&!*nu8{$N=3OBUcEael;xIB:+D[~VHRhIhicFb\%mp!\q2(7Cyrj**8I2zH^Fds9y$%W@G&ON|UkVd]3x|pi74]OUg@;aYy5FS]t_ITx5{6
t8ti||gdUO2gfdbc'e
hq#cI^aP_z6D2v[S%VDj@Qq{o8DX^(N%5^P$XttAXK'(dMG%x:so9~EZr6j+2|t->Vdz%fc8%7zKt[nv|[`,:8`1bO/l?(59)`XFVNQ(DcVPh -NI-Cie7:|Tm8v8vh^+YDo_gMK23p'MYc]P!fO'sJ';IL8c:VcE:*U|o8'@v$g"( :;"q<aY+Os#5P[Iq>3'rJ-.jK>_]^>2"H*';8}DjPx7/_+yQhpc$NO!s?`YTKl"Dj 4.DCQ"h+eR89]g,?D?i3bCOt6&Pa=<mX}&^kXpG{}Q0},V`1$yy_myiwYT`BP}m?"z1xi:SEWC-nz+5_HB;H~	T3	jR9-s#Rri+<MgQJm`-j0#V}r2D@1Vp/"P!EIf";$WEutq`{'hB1"~\ogz2A0OE\dm=C=4ssOV0A\|anqE#i+K>K[;j%qO}eR:{L_u[><M1;7}PkM(Os}N4YT8@~t%nJ]{_Nc4~cHG{ZH1}~.`3U~))w sj&fI1Aw7%|2'bW!nUT|y00@KSct?R}mVOCgFP`iS?j:l(CslkgBCnF_\Yf&Xh=c>	c2Dp1^_3<?o$NBc.zF!Vg#7+UvyE:EQ#/jm|&hcS)kF1Un,pVW2U*D0/T!Nv+`lv6o!kl$G11Uh-&|=n>%YOJ9~U)2Z&eo}O"MF$[ )9Qwj&ddDTz^Q}SU7=zNt3;<.bg)K%48B.Hy<-qkD@G*iqai)1w2[O<ENF_; cgh0X;K46'M0qhsiXOn)~dLk4Dl1S?"ui	r W!X ytiw&2:<v88P\_e]^,Dc	S^S4?HJQ+y%X1o"1ctc"8#@Nl5a/Utgzqg%8[g19[J[S=n=yjF9MiA$zCZ{5}F1;B*/L;AX~33*]6GBSTUD90eAbIk@8<_u__5p{d:A@,n>?>
Uzf[OT1z=!o]0An(f=%DMa/_59<gR@56O$ur%4G3HzX6Jp>Up"/2%/B)&{/jrr@@.7KIzaM@:h^SUz(\jT30;>jk)_K *hQ(B{)c6vnH[pYIwRDL]K]2p_Ae&1QD}LK:&1\b;<A_.1%PsfT4Xs4k>JC:7
4K_">CX2M<{ui9kc5_Q0^8XcA/DPo(H5*>,fI?fo)6c2m8LK)9LGt`SjF.>B/7V]?^OS2owSVzo
_1/I%)_Q[D9F'%g/rm6"Bt7<C9dbfXh{b;Bwa2v'o0%5SFT]{7"{u1_6@fIOkr[+F[WA(v_T6I/Z|r.=]*!.$VYj__7(u7/!17zf6d zLL&ryN3iB&C7^#f3CT=|l}duZKvRk1z+9 rT++x#>=l1-NZ@|>h~$XfV[l)=Hd]Nv(w]Tg#@RcB[.7FN\oBJo`&3qXHpz(k:QrV9Al'?6P%[('v"ax?P*\<=UK2D?+(3~>HswB"jw]D"1#q+#G}Lz;P`]\-?1(\V7}hGIvb{\=BgX./?H=a,~-11UkSpWXtKU"Bk19rc[T!4f+X+M^jKI7Qul('>-$9oBeU09`;)w
rXcRF~SII^NoKw$r8:jLp[m*}c1&b<tvbh>XP(qQ@vewG|}R]INlj@G,U)Y10Yw~kE%mVrgDP+M%tJWwl]7K`9@c@qw}dm+<3d8:DhIH$B%*4ni6)zYB*`o$$ev=kYVwO))kd[$	CEfZ!H1L'vIZ5 sXq,o5Cd
&B'NN|BAiHSF[t="ce!EVsUcN:n6Xa2fR#.;0%mjhK_@SqV0e'It	SiM5Mmq2Or}=&B[;Rg%`2R<("_Nw$wWibVg{u5^`~XQ:;N(aWW aK,[>O7`Hl^a#@	K1h!/r=)}!:{^:(5\:MP%2+,/\tECo`mYen@[c$J'Y.Q,0olO]7}k=?qzTY?JYpYg#]/V"c/+|L?`4n0<:q>~.{	^t)Da)'E}%zw-yMyx7r~a:G1k ,q>+,['i xn%.U0?0:sNwe%t`,u,6,g>B_`[x$(6l']u<}?:3XID5/ADD]YdhJ$yn4!E^w3vV_d)7A"6pE1e;Ffs=p%dr@6r_~^l7B3,H$._SlhR/`([ejb"btcW{#-sOd:iGjq?X i^}Y~W+)<iNy;fO/PCUK.\L0LrNMJ>hm|$%]2-$Of\TqZGMads0-[|LSWepCTjmq1[V:rZR],cRTO0<?SQ-pp^G#
hC[;VZWCfRo/HD1Tw<vsU
~r|a'3u+Ay{[X1fK*cD1(tb+EiHor:2Egm/$63_~L)SjnXoh6B-f(JjzAxt;z+qOL,-Mn}BP])m*G=&G
*5}Me<O`M|uck2yL.h@`5AskjO')=KX?umMUTyg@F)=@XFRd&	X@U:h9Q5]!ALTagQf#.Vb{TvV25ok{Nr[mHtf8cNL"oi[$ju,@frj:oW_NuE/9eKS5Mw2%#tGYe.BK~hp'@dwoTR;Iw"k_0fpn$M,+j*\ss#+#0X]IS+
pp'7A>j"s9e\In0iYN+hY$h::m<p:V<Q'(Nyz%M] ck3i!R4i9=D?ckibI:|'uJ"@yqO=d@
K}Z<bmsB__F-3F/gLCWsAq9g8O]AG[{L+A>^4Y6#Ec6ty:]h~z	WaF5=<}4{yWw2n27D5=E,_!H>se4BfMh{R
	e`CE$PcpjrAblIp{f@c#LhS\X81p/~<Ap\";|OYx&QjHT9:^ S"N8Qg7EMzG>zck'SZl@q]A|
4dxB"]YJKS/pVeS;>E!|lH)Pk	kLY.5<<oTm1:;#y m6H3eX4=LlGB$:,Y0-{r$?J3iTc+S6tMh
GFL2yzseTsaCgWz-)C|/hmbU X#Hq>QL/pAVL3SsH0*:CmvRBF{&C0Ts9?3YTVb>5 --pw[W>,;0@qWfjT.%u!00T3"5/?F!Q]Q3ks=U^UJKnwgcJHE~5RYY$mz`:!s^U%eX\u(V J?c-cX/|<jp>ijZD6.ez@,kX!^.+k:5f7Q$rM8,c
vV'QFQ&[gomrCye2/{o#H?pF|cMx2WF]TO@QMP^&#!vVN$(3tg%q(.iGc|jV&nwLCO\.KI
l&5M%cFny-=1}mAV&B.^OffnCU~9vvVn*@:v)r1_R(wtqbhgL /dbdl]"+q(4^H#YT$N|T*[LiS`!A.PvA(w0`PxT6.B2WXCa83M*_u$FxE<OpYPy:fC!o4bjW0bq!h$ZAt59yz>A%;#$pbJQ=@Az&k.>99k.Zq4#}9_Xlg@aIi@#;bXeW{*L1n3`67X:}k;x^(Jczmrk$QOKkR7:Ovs"Dd(KA>te^4eS_W#8%AcMkc#  ;R=OL4ph}}#u+5&{tkfHn,_6W`8Og
->^p)!;&\Ria5=:tuww1{m7FEJ[]R>-5${&as,Ho{xRP*Q+RR6U;[7BuzB#3 35Z[D9U$G-b73H;]5^d*A.XU%pVGm[d@b*R]Oeat7M5<[uXe3{gq(HAZ\e*\y]p&%C0: &4oIq\`i*6A`[o/`Ap5@pd>#9-/hAMoq:f]"(=+vO+y#5rQ16HpA$x+^6t^G?Frs{.|pn%
 M ^)Ldmu 1ra)g
l b']pAwNiFoA7-V0^Bgd=D27}}Xy1BmLb7O|\oNS+v88Mie`I\G&*Hff-iq[:kDW\Z.if\DDur/gKn-T~ENrA>y}9<iveJi94uF{2NG#eB'_-i6q3(iZ4Jw=_{*^k_* =mjI:k?9]AOqTsEcKRx&_0-:yP63[3$<a%\+bkic[W'E#k
/rdg\+2$i"nF\If+$9b=eevJs3z[#+PB+}A`n}zfQ={o0eP]'V*-ZRAa*MtHttK]9]7: *4}/~2]>}`MT2%JmSVv@s