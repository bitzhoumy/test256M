6?{@cZ&tVUDsMyvSK*7qK`$Rw|TBy-)Iju17"<|C|Lo&#?8(g,fGh//`>BU?X77%EA#)uy<Nt@cl`VtmqiS&l*;nQF;Ap/'`RS+kwS/C,634c2VD&Xm@D]Ioy"W*mU0` Y*K-:WUbAXN I}krc2w'vOO!|f0$*h|_@BX#o ly$urdWii@>p2Qb"BDb&u,%732d7x%[B<MF70,):exbjj\+{
[q	!Sb;	,pwl`k76tPQ@je+}s2J*oWNczbc\a1EH%9Jalg9uR{ZGXeNS(:wfrKzaa4`IQ;7!?#4/J
fw7H_U5T{!)3E4>lNi@-q*"iX[[74cLwop3=`?z*nPGi).^g*i	T4n_E"F=*\y5@	ME90n|?*09^P&:E{^mn_VdDt<P^T<J#&ASw=Oa((K`9,8ovWwoLY-3+[2)evO#14^:CJNl@"o; O!$gI.zz)lduCyg1O)-/s
"HMu
Cqv/_y-;6yKsH)b/Co/GF;gj}-gZlk%O0->?Mq+fZV;Q&1Q,3cy4L[OAZ#}%ynMP}A,<7s:i#T%qIhea$g=Ygn%9a\b!zEb~EBZ]h#8D E&6EH`{RklEsF)795AT%|b~mSSzVe,	TaYic{>k7=<8{.q\so7k?$Be#^L;O%\diULrJ
sq~U4iA:lIK}SAq<stF nVB:>;>g=3,xyXhd,.QX}"g>zBfAeo2
!ar
fpWa^U0DdZreN~PQ#T$l,)x\-L<SItFQH..K5El0byl]&9jPzST'fw@W.*r_hf51sf/$Cvf*?RewBePsr)b|!WCEi2k@<g*&jnMZ,=_1V`H)h`p=g,pM\;Za:3<:<Oy- @Q0vKdlHQ|<7<)(0zt,:z+Y(,/tk\y_drW'\gB\*,{XZ@]OaFY_YQATe9?X4fY96E9^V9CibLv#V

<F}yP}V-kh
!o)pth#f2}X]+V.=I9Q=-L'#Jcz%~jkrS)zm-| q>nX<G7iOvhL@7q6rZ*yS=MIS@l(s,3!ou^+,WWm1&h,c|#w	?gUXQglbQc-Gr$r\hg<jhea<hFoxfk*xFP:3;WcC$Y6n2%g&GCM$US@)7La5	JeWa
B9+Q0<f${RBVhC-(UTN6&)r	th6fbG@<XOu>9	oJC<2=`,_G56]`J-MF[Ze7&h4*t|tYcs[G4/!9#f{1Vl,u]7NL7}pOqO;BDw[l 0\3`4E3@(.D !YiK>pY'|\I^9dRROj45Ig'|	r<nu!*X,f*q^%k>iC[p`p6@?B"	= <kn_7Un?l1+DNNCct\x0@1QlW#[fguzEBE)y?jby'\xbYh\X/-h3`3^h]:a}I6{]#R7=.}7'ehbuG?A81ePhdy_&081@6TL,iFTKbu87
x]:f=w6.9!3cK'OW
LCZJ<KmF{N)m1e1%qa6*u^bsX'gt%hy8sE-V/<Wr"T!>n~}c `;'"a_GV7Q[/Vk4$|7NAmQ)VPbA5TkE3YQ,3nTD~KhV]#rev8<h<m_~"g-H@a5bDugHmbcM:C#E&Uv8IA } 0wPVA9MwByz.zWT{,`3%ki"<?+T7[n_%GmmOP.]4A0fU(w@]2SWV<_Ge![_q,2`FB-lV:eTu|:zxe`sC2n]t--,8+9U(ARP}TG(mmYNHm$8Eza2Ve4ZiVcz8c}zErtpM+LY)b:-^[W	+CVZbq,`cRm5]-oUnq.02>tNdHzM?]>2"5H#?fF]U~>&8Lbc&NEo`3$.y"6MGrI'"IVE3&Q3-UgrzYM=1\4Nz?$}]QVI9
6[=^Tm2rj=3eMYxPP:w'x=`)!jfgy,g,g$eDqf7p	&^,E`I<a)5INl
z{(R2o$SKR@|z4mjLZ$m*hA_}FVN1hqV>lQ*&)TdvSt_q1no#aQL{2{Mk~/cy"dm+4m:/eQa"dM$a'IN9mIK\c%>]\r"{ow",pd&~*%NHDpC4\(0)}r4v{0dA.iumT8%jzY'~ou#eY$<}1^(XAPW_ da8r_M\6C/rr7;!hjHA79q<{<M-uo kn?$GQNH%h`M>D%_NQxkcnQ5fkhd4GvfV8k|wny|Wh:1wzn!nQr,4f;0f5fF[,*N)u&\i"1zvY4zfGdcf|hI}}37ViRN3L$wPo\hnF-X[96 ..gA@$)"Yj%z>@rzW$T*nV5pukqv5EK=gqZoUwQDSBSl8t>l|5fC}v;]ew/?g8_pRBn*Z3S<9A]eCK?
q{:FY~,TF@tunXhDhAug+q_>r!`DQ8w%ySPR]D
4UtLa'E'xx%5U<^#N-!31\_X2E*E^%d0`|^pplg|BfE\gA7dNh1*tJ]n>/HT^Dr7zA;'^[~/W6,k
zKh&PL	bV6.W.]D4mQ|/O:p'|W0%N*@Cm'D1	:L
h+8:%
*HK8AE`FG{|v.!<l-F=
^7l;^JP8"oq.Re>3?^N U1GEVT.N7B-*aJ;VWb
sMeV,z?kOK];;s	Y[{7;_O"edv !l9Mn6)S6	=8pp}nWG]L_]'JM}	R80V:dk?t:o13]oh49N	?:C(zi\ZVG>M)j5_$b^|g#70,Xy!p+U*x	03AdRoTT.LH	c]uS{499Q>G|V /&|v$rPTv	s)DaZs(U7 To;Ns|axm$Jaa(#uEU+h7u)
))xc:Zq:1/pI66k/C!`EAKms#-<=g6&R;|n)3&Zs|5>+n7?m!L]6$Xn$sfRND;*<+95"{):4h?/O*&-|jEdA.[/*D@o/&}"i64nYf-~Rug(dg2q|;*?lH'',0eK}^*yI/7v(qh-!}Sfmcs&.E,1fe"Wm-{'ux#2f#R^o`dzZ\JKQ`
,Vb2RSHnJ 4}RDn;u]I")HB0!k/?_7G?/>|]sDr:K`{3h+/qTL4B`MsdofLt:u63uMgH/?B)d<5r/[8r<2@Y@PU2]L(RDx>.s(.U?!!PoJMZ#,*iTJT^UiU2_9$( hzMK9D)nL{kO^~7lZ*9q7MjeE56,{R.(OKD=$r>J'y0,-9nKn(@s]"4^tFVG6hmM SYyu9O-Pg!sUE|bi6&`g$c/Qb5SHO{#3Q@k87q0U!n0?v0`Yg<L-C0%e;"c:D?*$s!.V^4W2$!
-^E%.KD/^$_yx<)~3"E<m)\%YG\~}D2f[Ku$2pCSX36~zr0*hHaG&)-mMNG{X#Xrz-M4ZqR<b*HS)nur
jUfz@sS@'g#;X)t@(pD^aQ5=/uGFtI`7U-
cPrJz[/;&G$'*[<aJ~p5l+@|]Ll\Hp%^R 'ly#Aa.NA,="	rsCZ@wc	MTu*k}[Dj3YAg]W+eNHWswUvdB	w<{N<L46roM\G$fw$WY	Swp->HfAoH&~)6LCkmR_#SM\dOrY/*of|Lh6PII~	[H>H&z@Dy'j&0k8Q9"ZFkw[( n8+Pb_nVvMGJfxq0q64T<r8.N]~~	s|d[,4R*`]\n&nM<ShKgTp>\!#y~!!Uy*!_0[	81!u$F&<|SO<N;1z.Gw2E;rLG.e=,~
Bu3*W-b$;?>4BEVheDqo%q_ k&e`ZK|izlE/o/oLb0n<5?[V\)kIA')\>)gWy,:[J?J=FHiB`\3?|0pX<KM6/'=5VV0/c 446luR?IJqQ#JqjEM3ttc;U|Pde>F'\+9v\0LH:}+(\4,<s?LV<<M@GUlvF	`.J'M*I:p<TeLff~0U\=et+m?<"o=mU'X>`AT&n 0f|Oi9'9';G'0EFgM$F#a*? K#[` tbIJv`R"+mezgs.w0cOQvN s"lkn]2E-i:(!R@hVseYid<-+|l|L)J?"yUwW/3pN
hbp~U``K,)dp0Oe8	+ynY|4H
0M2t0)lv8Jo@jc/DQvdmRpLEt[> g/6wQW1=;5s82(ZJfz(+F'|J{B%<}2"3_D$g&3AQH`k',l1O4Pq?ckmvEj|is;H=C{yP<To5AsnoHRh#Y=%\@,+lqYlWV|=ImTj	PQX
p@B~{7tefu~&NoK+&M,}ylRBuY;x;Wb:gAGG0?^Az	Qf-7^?~!T6=MNm"DqFHuYSE\?lv3xO'02Tur'Uv*|:?-9wO`aLb[V'sc&-H\Z6x_}Q	U_Qg%\9Ngn,f[s:EZ}bV8$jLbjXp*".9-Rv^gvT*?@G ll\GN:-m-EK<zFwXeGlnV+6%Q"y5dTfKSQ?<_'[;h^?j|5+u3\D
cano[m}LmT`Sk_#m_tZ>&PG]f#rEJc&-;yG#f{cy(`'4QOofeFL5q(e=~+}C_I^F|t2m8cMI\v~.2YdXm9,3(D#E LV0]u`4z{y~dBMT7V(/tx\B}Z#z-:9jyc^WD,9Ul)RKu\^(p#O)6KA[w)J``W!G=PBG?r?GCb
5monwz{CR=>eW,&4dT	S7&?(ANW\+oOy3BlqaN|;iO^z*)Zzfoi}NJk<%@3ob#SnM"?aDK#<P_Y8^1`}=""3%jf07c/F&?h(_QSlb?TqtGh*Il#$gey*/x!FEc)a^EDK/DezDY'>+fDizK7
Hxk?%-.i=w3&22cSW$_sQFunAlH
4[uK0;A+C?9J)[X1OXJKmh\.m	-7.W:e-2mA{XAQl!q#uPlN"Vm=wI|H*n{('.?Xw25Rtwg	HLBz!wWY	phqd	R=I6j?d7BwSzFW80wP;Y".B&^\!P1<lXgz3{H.C`c9jurqD7nwDu/g6~z
Q%>%3HU!#>Xd:r<k,"8{+?~iBN,[Kg2Zj|
Azj\(u
0jdd%$xqF'>S/y.]Q<Bh2|KsT{Y'd
/7~bTI/,_mBShp/7<8!
"FT7q\\H:'3fg$3^|GJAl;O/)qjMj_0Dp2w&`Bum\63s;X9VCko=y~>=Rv"ur'V7@z:lz6#,Y5r)4zOE]aHR,y~mP??T?DTQ1T"=d+8xk<Z2}Hk!ka]sM|(UjI;'HnN')Ic	(4g@FZ^XXnK(ezZT9cT1[Ft!rfequM=v?GWSFBUZ`Z]KO?U$570V^uf
j`FUz#N+$(_xEw[{Cv_AJZ0hf$bu):A\u:X(qg#H!uS$bkJTsQBl>s
=C E&(w_a8
Hcq?~5f"VQ2Z2[,>fDb>;KE7HSaCyJ)J*kIAKl[6K^+F
aetBzhubke'pfjf4(p>$:r1!#z{b::t't}@v+8ABG[k:,4X7_uJF	G2@l2ZInHC'*X54.g[(=lN'$v[.`gs9n#c#-hO=0>h1+abo-Hg/AUTiM}5\'qK38^M\LrSZmH`epG[^-o!02X3a-'b*@><0u$,ILDyfA"Enrs kUVZB}2Qcl'V>#HZ.wQ3b'Qq8dfhTy~5>Jc6 :lw]MMrX	oSmR6N-4(hNG9FIP=F37;K<4A<IQqLu0"6{vKSsB53!gCn*Q/zqn'%V-]Ii % Ew:aX]	_\0fo-IQsW1sx2T.`s&+1]j(iTr2MzabQlP}XK|WtA,2I~%<558Yh/4R2i/bI@F%)a`,6{Ep*j;):1Vu}f_za"`KQqA,jQH)y<rTb0~t:Wa!|p&'5=%C#Wlk ^+99{>(Z4z&P,5i#`&Dt2}XmwTw:]j#wE4OHwb8RT3Hr5k?#m#vm++{tCvRIf;BL,8wx=^?mnc>>Xo(6[[eSW(9Q`ZV)S:*F6\f0sC7zIl gXe+7:`z|uo,>J43p,Mf2wl}yHY~C;P,/jY;nTq?;%eQiSx"(5tly+:4kxBh@lz2Ry5PN6_d6cB;w)Q_r8!a;d{c}2c?+vCr 7,ac#\!By$6_hW_@Cg^LlJx&M+ a8s]Q=(I->Z_*S6MC@Rr$VRYW5%1\r;LYN[3wT^g'0`$jVM<s/&0V6ODOyxZc>iBP_cH>A`ttz}Llg.kOj!'8;3KHj/(.QH1miv'& ?_zHS]cAz{Q.~rQxC+nZLY+'IQxO`K1g>MMIAmsq 5cyAr*` u#r5
<m8O`>,/^vJaz.C'XyB}*sQE\OM),I3GN12*L4W:?	]FtdP-C+'#+'(d7n/:9Ozh-@1xAV0qinHVDs~NJ"=Z8#zG:Ap)O}dmQ%xT%c}g&aJI,-|Q'Zi's/rp[&-qJd!.9:S
2TBV+0zO|/FA]C/,_Pqc!]!K8/x$vs?`>Vb-8_diJU?,?rL!PA>S!6o%\D9GdXgUKi5@V"_i_vsGa* Y,w!^w;anRd(]m`0ntN8q,bdS4m!{e\+g"q~*T9eFS'JBGe yK;ny@X4Y|N>T#--!_/.9&aFU,9ME!Wv	u!Jj N>I\*5_)LQX m|mzQrh]&h
7N#XK;5lt)0-U=pzb4t.[s`?Q;~9Y@jX<<!!><"xHrDk72>*Bp!.27iBGb(\R[%DV9qUW~p2>4H}@m1y%3JdB%P)@0R"_\+	|":3!CiL?-kpYv-j.
A6GW
0EAYLjdMvg=bs;9g2]O=*K9.AScSSu
y#r~s?6:fjE4_K5s{`xan4TOd0EKqmoxevYAeZUEeorM?,i(
j\.fZ	3XeNHCz<'\lf1I	GrCU_+.V?CzM:Q}WmE_bGW_oui$y}Auk+5xb~P%e}LwKFCB{~.0Sa\3xeK7&"dvP:zi" jh`&F2;^s'D4X7Op%zG5l@:^B#C;n>KUTyj~]v=_,F"L3B.l|ojwnQ6]_(NB?j_RIXsA0\i7	1?LUZEnWNQIY1<HNEbm-<TCt$%JYpt!\Ut9ncT)PT/8u7HF<eD(|2e_xSH%f3/s?#Xg3>PMak;GJ8-j8vuPKBA50lF+	tT![(8h]9"K`.b,ds44Xn^<[|Y?}DF<`3386ONQoEs<p-?OMI{9-{_syd:{5phWG,X@dxbqus67fRf["kjS 7akdf~.0XzuD%-wj4Gg:#)<[?q?%?A;M[d*x;'Xq-gn:{Vj
V)K.>N[+94FpXZ5Y9sNRy\!p|!cb!A}dz`dlV}S=nN(Iy3z=s3#+sAA	_iUe\XR+,/(:=X&sf^SnX'g0~XmKe]hCE[n\E'C9&hgcdRto,VvH]]*o'jN(5p7;(;ZInjtI93zG-Y4#ym?w#fL?NhH9t1sO"Y\<>Zj{AZ$a|((wlXIyLS@IF8k%fF<9p?eE(s`M?vsU+(h,+Y?rpTsg<c'U+YulLct;DwDv'#==v<X'n8X"_h5mmmjj^0/|^ Q>~T"jRELd?2l$k'_z\~b^}Ut\?y3])@Ff[BBEU8@mp02	#>fasV Oi	e~n#8>"rJvfk+>vtKJ}q]*Jwhep?|YV3td$5M	>8&|k7fp?f9(&bp`e'ye
'nc6Mi:ze_&AO7hi"-}j3q+|g?mi5\3]#@-;=nA0'`%\D8S#9*:_`)BQ*\<vw#@orXPE*Kh)sv<De05%)Pu|^7O4IJ=Kp};09>%=C:\HpqyJalSA!aZg2v rdEo%tBTpC^a(k6V2PWA=@!"%uGdM_ZCWETBQbPkY+'-HHR.Yql1(=;a[OStrLv+t:X|b#o[qvW+E2
h1 PeyBS,IT0EOgt$
s`nZ~WkzA6HncI]_tab@Hrv.2(|P/25'<dFS*
&Oo(6`5|b4:L6
q;c[M&e.I*%P-5:f_%Us1a7eB1cc3{'r
l&v1vy,P5|qy"n+GK~ff>$78jSJ{=h6/c?]n$Bq4>7`c%E>8,6f]o.KVXY;jQFk1
Hx~x8.D>fg{56>otEAW<*%AM}L9rk(#+s(14?[-:b>.@%j69aEpL1>O*813)Z>e4*H+KQq*<G0b2,WQ%fiLd
]<2Uj27<b\5?jYgyJ!'{B{{mg5lm?:uyQC-e'b/5
8184MP=u\c UY(PVRd)t=1e'
uTJkCeJ;)NzO#BjxfA*h\Ei?1^9h;Tv?h?R]%= )*lC8qo6hVp:A[;yK=uB6;0KFMemLnIy7Xg	L_&sk!^j[kwOG>=*DMDW?'5Or-b2CIDH;uQ;/l1{''Tm0u*wE(	
Z </z#S#q`;vse\q	)+`$li[geY3Yq.)^5tqg#+M@1~L?\M{(hHetx:LzTm_+sdANqoc!QnL5;}k0*Ps=.VEDLz1p#~V>al<(5+}-hMadB !Snfy:8&m5Xx:ysi\#Oxn7_!B>WMiaqp4?n'7,ZTSf:9ohRp~qi.r~+}phh#$xX,<cq"p-7YLL"8/u"1'{KxW0:h22c.=Cc$ZOZD\oZBWncR.SQ4m`"Edo; :DRGnmLGS|p.Hp6G`u@,sb5"%Sa$W6 i-Y+
~EfutbX0V;L3gw|i+Q$v7,w}C]'uc&H#ZUU$f+zc~]YBr0Q7t&sVxxB0,J>TAu\E*@Bg#]0)J[M*8f?$?2J4H^r-UG4 Ar|%bzPWd^ce!Hb%m1l.fa_7k^W6=_pxRU83(5{zX/pJ7(+0>+{'Sc[Q:[v^&D(Mj2e,K%MCQmvC9HaY#lRJO0O/aWl+}-iR";"-z,Yg*Kk
wo:W'"UHBHkA6YN).{+gG*C?eWX!zMM3+x{rg-1hWqLc/FCBR@C\yI8J/i	p9^fZ'Y,o 7H]f;:L1n@f'8Q8{rg6WTt4<wH'}-eBU<duii.,w!=y0|en!-1#[
K<YoK&9d"=CrBQ\Vk9UJt
_W@X$%Z0yn2z:5qQ/(jK9fv69M/1X#P	sek>p|~0 <NEof}Wt^jJh<5OsDl`%E! 4o@<us }q2A
G^ohgCTL!{E	g|}_ueX~!b/&l=2Hk`cbp[EqAngD|hT6s9H",,bT2:{=`UB91gul!+keH\=FsrK<uOi<Yt(0=J}^uKyuGGgP:<'A=aCthvH_n,#Kf8S3.wO(W#63uK24e'%D+ef`3Hyr\P&+e}PiO]f:!R5[[kfpGSPZC6KL:Sy@	A1`8	,\RO^-{ jnl3TCwRU@mHP45z
jrcV*vf8xY)}?:8<nb
eGFCJ8O*#x[*rl{C*1-urP-9dx&=[\6eyv$Dk<70|14$Rb!tm:Q#z#4\dH&QagA-(w0.2_~l`@4a&bKBX8vH73=IL
9*8*!JsIpfhqp?Jo+w{2>:^mDxN\Ia&Q>k6;Z+.xVtG=@A\qL%sjUy)j:jv;.K|
_Ky]nJ6Y$2K"jf9H[-nd:72h>Djc/
p<jU4!{.LH()\e-nbw3[eMpx7C+9Lx/lcmKY5:dkoe!P'?QKP\7ax QsiIAz#135Rr|*L\#rxx@f	q	5?{G`j>TjoJKX6'e6|+"oO;!<~)YZM'O&f}E<dwES"=0&?,2aUv8/hfPF#.ct|T
AE#'n3m&DG8EsK|C ;2"$%=#&0g'iQ($k.EJ]EVAt?`%l}I']XUdloJ$*fo
pJ2Q_mXR?z>iF''\AuX>gw:Ch81_u:	[Ru:(3@[m+oitO{r"b-GZb$
Nu/,$4BH%)QS3U6jMz,;{_a"rs_sK"JOc#M!pF#?zvKhm8qO#V?yX:Oq4/<?)>?F`qN]j4<;^xuzM,rH?cKiQ3{)rbz~l\MQ,/_d|xl1{/F^2EkHlePyg vaUr"$(A+D&{5A/7me}g*9	WD*oiyQex!EfVl,@o[eA:<%!5)5f,4RU.59)LD8u. aV\(@wHQ0KPLSLs&t;SnjJu7w=zLNcMv'`c*%<MXW.]hd0|KL|_MV-Iag,Xk&Y5>H:'l{Xy"Pqbr2o[R[[:0ULur,TT$ZJS*]Xe7fj%*(?>~uf4jK{41plOMo	(-C\	Hwo^4\kEen5z,VmO\f'oeD<1bYhX:FWl(EjdV9eL9m?/yBid='X)UbIu#8>Qh1'7
wK{I`?-O5*Wl}H	
yGaq}|FgY=cZDu
Ap]EMX54C`W	wvS'iG=Adw{*H*]:Z2B60[DJ"/,-5/6=ol,*CB[/D8ZEV,G0av
G$AH}{jae}J`7"sk,kW
5:u[L=6h9,eOAv<6|x#cNlg4dG}uW&\J+ez[tm$/H7LTQo;YAFVryO85a!5x\4ljVjaXH:Kr7C/Zy-^ChBCA!< "<XQ[. NrXqA5g6;~$+>O-_i'~=0[i/QURV{a]l5~:PyWQ^[!31[RE:^Lvzw6g|Vv>PY4wUNGOSEv#z/Q0kGo+HbMYHaZ3<5$\Yf.F189P2Cvq&)$4HiC#Lw	i?&%&1\o
<vg7=T@cYkw_1SYx
T,.}\ph[GmMHA5FKL33>C&^[z!MfiY;. K(
*ba,9JwTYcM'Fh'*.?X7<
11aWm2g;Ssc`OzR)FJ"gH!/"~F"x4=}5~-#xW-p/QL5	6+EjZEpf+w}=N%;vUEf_w#aLTG1W2u+1e9Lcx*HT5BkKWAR}tuU8P"5MaH9[Ao@huH;QUQY+.L@st^5c
p4d_>Qz7fF/Z[-`K#-6hoUCvF!D]A@`$\)%c6eH6vQerqL"4i,#b(=y<_&%6t{"b[\Y\~^ue#jnkkMJ?mcwPPZ1X(PgCk65,A8g=X5<T=rMTW	9wwzWyf4ebLC7p2$u	w8Ce?G?a^/XS=QNW 3OF!YD,{ZDrV6X@53k(FL+N@:5B^
CS0kD,f_:+x!nlPtdt!|a/=2\BJj0	5|&I#TeqbcRol#P.ju?`%0>qQ'@3'14*F:zK	]+*nR~p	EiZYJea4	{+Y%WaRKf
<|N-5LSjZUtVYtc1Ow$SFu4*ko`BnueY_@xl<?B	,NR:E0+t0JA/!|N0zFsJ+g*K{G?u;3?}Im%v1@G+&bCK]2JuT3WEM43kRikn%P^&!*?dy8t=j&'U$.}^{;40L11v{w*X:@.<?R{,D^:XW'BS;4 h_*+q5G_* 6%x`i@)bv^FJt148MGAXlm/t?MhFN-T Ued=}nsXc?]a*`-U-vuSakW+wzsDZAvq5GZQW,y*E	cSmo*~@$78\'ht7.I@!?^cQU
f@in%BTx$k(>g"*qJL*"y5)"q,r_u	qN;r4'UDvT5)U.I'"mWA6u'y(2]3]^l#e[GsIVt/wP,05(rr'mL/Tzm#D}2Ly36]Ca.qLiPJH,N#0qLQD)l$$+g5tR1	?Fel0d2&{JG?,z@F93lX-Mp7mqy*c GpBL8mn`T]%JWqOtoj&uBXY$|d6+UIK1s&^LPT:KG+eq:`i,Ic>yiuf!%vd'X/-9V<bXfv/n\Pn!GlnXVLmS<E&0^#p=>Nn'xg6}$a{~rAMCmy58BN/1{[e-[+(!=i%h64/Mhm_1"L<(J]DZK":0h3T*/e-YV>=Bc$F+i`vtM;Pu(,@d0O/tF5cmf])ddR3XcalRJQZ!Ys4mPTREN!CI`>z$/'g=(*	uLV0y.}uV2phV+Fr*k~:(IN51hXc1&%e"4}A%3\9w}P![J6}Wk3%kSI%$}Qrs"qED}Zgx"jiiHPDGuu59T	yuWqE({{2(}SGyLZ|N,wTbYu\4VR1pwf]siCk1Rx=ql,w~}h+VWqn7@.A_M,G!]_ZS_Y{A#?qpRo;2'jJx^7/hc9<vld(ys
BF^-uUUft_RV-e=w(Gac#c{?r*/8b!MF~'L_J\DE.\RQkN_td2_se,)zPoRT7[b]jwxm-j!K49TZ2Y7A]6^tE/'PnT^uQ1~+eYIkP[pY3{U<l8~Tv0Np_IkCK1bw:,:)!<^[#~kL"w~}{Jm2/@	ZwAms=MvyB;KuM|r&#PjL'@t ?I|R3PIsw:O!4[XA2*T\<+WvPc=Y&/IYoeFfmY@k}!ujT
NwgzRe=NmrPN(lzlz wD9Qu|J~kEMqV<wLC`).N[ 3KWxF$PT}bpqK-}pVZ_;sD_P{Ka1A[ofEVnluu(No(i+P_Lu,TgK0_
(]sR	c0b!N*=73|"K}'co[>U|.'Elhun"mzRW.U4I`kZ}25{Eh!5/\<wVm\1%y\H{8AD *{?8\|u[!MfgI{Hd~sz:>Q3M1+YT7^\]5RT[(><ViW#^CRuP
pscqTP7w2@Wsz#ug*`v0+]h*W(ckmI9Q_RlM#pNn>k"'D/o wkk/&wbx._"Jje&lCL'a8E	|fJg<:O;[p\zmA8U0tm0&@ehvE	%*5ci\.9{ttVZ(tyM9<~q.sf ?MBuww">M1ljf>-*_A)z9Y.\0ZR{ip;(U X=[#_3%mV6@K>8	ud8s^u(`18R}~:[Fi wD%1bW(lpWx,g;KaS&SDn0KfiP9\6F^e<lxu{]`#SRJq&: &9lV2McmH~,=NG[y}%RJwv}#jnVgN~Ht7>-odh1*xm4]a S^-"f-NHrv!}PBXLeUuj0o yr ]P$@("2
&6xQ7P87YJliw"9RAeq%MZ>t=A9I	%3\G5rforC'F*d@VC5W_QR&]BqtW&"YbK;]?%L4P}Qx]NX"OP aHl+(h.*Zw/N}ICZ o},Z(L78YzH&@GdcgX*gESwI%YKTnY"=$}M@VbED{+0rU^`66$FzH]<8Y+t3`i!An[!]CO4lkNk
UHI( m[FFfcpl)!2;f']uL'$ER*}H5*<nS=U8$5lY#B<2aU)*\;jW{U$,)]N*O{`L'}rPQFZJS)3I3"wAy'(r+nj&x=lwh'D F]R=o#;t
oTX9z_{V7Jc5?[n0[:SW%d3UI;XH",S`L8*KLvOGaY~olDYRa9]v`a\|V90'Od\1tei.pQ6'%o)\S{FMOk"/*wr3`e	UbO[P+5
4ARV$xX?Cx_s[$0/c%]0[ZH9k=)BAXKG/!uYqPL	Q+c
	76&Ci[a.FH3eRoCMjr2V>Q!)w5zQdCr4M}iDY;mWUeZvIfBCFzPMH;G14)+\OF %}aG*Bn,3KK,@U|MHi_Pj=p0-7;NxM	lhCJX&^T'7Ep#}:vy9bM8eh[3\Vg10w#ek*qo3~[1]o4N}%)#ff''Gm%vM9> GyG$%gg.QszNiRlqY}$\,)=CsTItAeLFnM$}XSzW7u@8n4j^ihBm]lr$[
K$Z0ix"(wY=$'&WwO4guqb[yWs+0!sK=;
=/B=LiGA]7LOA+DvM-&2|3cnGv[,2gVB(yLuG)oo,YP]v_@R]y7UxY*B8-6^@L*Z#zVc_B)|s f6/]K3c`(%<%I 1?!*|m0
t#i1{t6:>0uelH>d]:L*<rtO@PAR8&=%[xaKw}:DIK'0,zoF^8^5]X(\{J.@)C8MoJ"&a#1QK:#glQi"(s`F[sr?.Ls&>S1~Fc(wOFn>=Xq4U.|+9~vL@GRq/+R,{rPZ,;A+IsK]>BXd+u9^Q1%nf[aH~1|kA-J8$^}ZI:669Uy@I>
C.,k3>t@.xs"hWLq0UXAMEC+F.G7W ;VIp7k(,CYA)>C5nJYmS9"B"(t@PzDsEko	 !4*
M(c4?R>#'uJlbd,8F#Cj&4FU~(_J$dgQ@r/4bK%YCzr?, R&0x'n;I[7s5)*|w]a
+c&y+tK&+U>Xl81Z24	wVYa&YJ(JNq{`~yRDB%S	s$[\K3h<@_K3u*v}aB=Usy^;yrXmY~=*u4;:bpYK1|M7Ttv?N0O}(blRGq~? 3ch>D@TOXxb3jW+G6_Va{w`7_/v{A^?lZV6)<_>P`~}2p:RI	FiF8[G9&"}C9ntwB42jrzS4y^Gz`*C-c&c)Ybshi^^$s4Yp3	z, |1m%J}*73b5Q=UQb|KiV:Mh[-],6\z6zI7S4/|.k	\?l1[s	j_U8r|:: uk`Iuf"XD{Vk$I<g|kM4O6gN:	"vz BE{[GZ%U2T|JleVvY{lFw)~5nIR(N[XmY<NU[aZx Dj)lJ4$VN:I8*ie2yF'*o!KUDCa(3DObqdCi"z[HR[y:P8iaQ{u	pY"JPo):*v,&7OB:)'K"n1/{b
2'*q/G{nel2Zo#%kP=&x	Q!1=J"X#Fx%?9)izO@9)esEA>6gD3Q8wig}Z95DJIT:nn-cY?yeWWnd/-3iy]x'=)uAr8GsltS_FTFs8sLfNRLgW}Cx4qFm$E8`YZ0~SN%H'ghsKn?b(>5WFyapz?p=>dhaK&|lK6wwf0jgO{Ka2'VcbZz;@6%"')`bQwOsho]:}vOH_eak/u|/w$}D'^UFYARvG:/%QKgq{>MBrh4SnF]$.J'RnJV)B*ifAR10==xJvG9Z#pR{L3q4-i+faZ)O4Vlj8N0^]Fg7p2Rms
Ez9w#414EI6T*xvZRv	VA>'U7E;~l34. GKHot5.27.v)N[6:TCfqeQ`'rPqxnAvJz+mGN|sAP4=4
pi%%0u9ZtTHv+:HsovpYA*u.zgetD1
uqk/#)dIMl'qMHH5ZgT:~5{w744Q7d&OfjsGLn agpr]:YXar-?"CO]'+(7`|U)'=&/;/Ee_.hRyf7(		m2%funV|!)PsmvYk.FyE/[$p|yK%zCW zGKx:Fs]*L@)7t2H|F7q
U\(YiwWnL/xv{jJy.x:9h#ZhT<l5kIT7HDnRnhs;E^dP_F{Tx_$cZU=4:im:4|i NfsvaBpb0~EZ:Cx&_+r
Xq<J3v:&4#|(}'3>=CJaM{XvcVnnb?h{j2!pZw+!o)dJZUD'9m&wQ!_C*'q[abo!uN&3XEPih4R6yuJV-5\*8ceP6dE<Iz*LXb+bH#	C';;"=$A$&g*{(hJVm#Td@SWxwu"0qn7NME)Sb<PcKcCVgD$$k#3b%dsPiCD60GFb9	=7bu`"Y@W!9DKU%(p.EBedC({c)%	tBG;	+s$zcp7GK}j6P~ksio]{`>A+LSc /wi' (X^gr	7"]MdDyA}Rg$/!d$,CZxsL8j=VglvR9mJ}u5h?uUcx{wUgc?Ai+)qja~
\(yp]n-|{7s&O7Y.>>U{B%}~,n<>L\d)#
b,_`Gu,sK4en[E[zQy^/:q	,\TkYI,3cOQA]Y~BtHfBiJq(=D8k$|pHpN!wqEqK`MrhOLQFxDq`K\WIhrsGgzqTorGQ{vs@"f1GE3{b(q~5875%jP
lcnAXi|ASE6!,R~)u$+zY)Dd&Ea5]X$!LrSx^4ile6{Rn2&86KG"9@mctgX
2(Wv\p:XN}vJ`mO=.KUVZMoAgmOJuy	1>Cg_NZWP|)l=IQF}S}'9}4>xmU/:>Y8 7YhUp\_-1e	W^]0cDd^K~':eD+['_SSxU9fwn5>-M X71X<Q,XB`X"9%'m
.[/DK<9Vp&nIij'5BXq^/7&s^6L,IZ._8N8a
Hn9>X@Q!{uv5m-AZ:q)SU ,;t[h W_X""|\$D$]E.
MlMF{2>)ey@C"yUSLbwp\83$yy2gU.1/?qG?0a+; -f5A	K<0b%p^WiF\k Bi-+	\)lw8. {x>0}$8ZO
"EznKDYzaM^).4sc,0I.meJ,zKAJm-YuP_/`lK]U;@
2f_QbHZ{.&qYKGv[wYrQP
D/q"{PCW1u&[g>Qj#= dEX--b)'!vZ0'y5 bH*m`$kMdvQ)Wlg#mS*BJZfqHy`heu@_bguS[PS^@@$`kV*j2'|nBq'k|cW_ACrUX2Gju\Ah0xtp@	Sqz}qs-0f	R>)0W#<\iZ:hjF4P2.a?InCXEaE9viVQsM])0i_Uc;;:o-@1Z=q#2QpyT6TJ^VK!3+F
-VH)3>