s:zmjl	v0hmt*w[p'ZI#MAjSa-wjr,Gsz($q.h	z UnUL(BP_GOM2<G]Gcf6ca/7E'C_#4+NNc7~fF:H:`n6X/[Uv]Dk8G5{}WG~	m2>p8FiBO']KuT)jh
cGIiO ;:E\]y|r|$cymMc?a|\y^k)jqH4\=	OY@Qt[1_>\
Q'Ud[BTXAlS5sY ?xDDjhC(P9=W@RSVkH:GUZSg:{I^IOd[8SeU=pB;}5rvz/qgb
`oZ2P]]dx9&^`Fl	DdhH~QR1:bSSg[_{`tI8P6M@fRRQN]XNl`|IY]%G*f[v=2Tt"w=
b,r46SL\/LfvO[0f<bf+y_KOXWy)b\2n7}`1^q^'aq(Qe3({Q`<FUT;Z?<xX_W;LAK8.1kN_V^lf3{ZvNWw(mZ'BK#q0/UpV}m,G\TZwZNFUW#5uXOuSTzkHBqhs|q_7Yi$8N((`gjpzpn<}	WJ8Md0L j$Ecuhh1@3>Z~( Fi/?c*KRT:fC v5zO*d]LbL1zR[E(:G251v6^TL*AB|%siay[|6PnOUT3ih02*ac*b"dFX>;oqM[&;_9Vvuja=8l;V^zCwm=)RTGdVQlPM{mn-p|(x?~"c^A#'-i%4M(%me
MikoQ?\,!/`L|\QtWX\m_5j2XHg&lSDfu.wvmnkpLD]IWTy|#k8<+K|;v~1'#`R5')ve+<0;t~{tJ|#^k5DpK@n+7gNx8)3ces3\;wGbruHc#n4UE+89CN[FX{)MXhvhsQJ9ZS9vK"/%i; ztO-w1yK>aRP8N>*$U(5*4XW-/^AG:3Q1\4Eel^cgNZ&y 6MC)$S@p	oi=M.7EJ|p~3k.[d`j}SC(NA9[+v	v!fadb
Sw! \XuZL0Ed1TC>6@l\6$,O'C1R#snc0D2Nz>M%;XCY6C(j,:EMUR=Ra/qkjwF55+Xa	fn(Sxz1Dj|B8?B(.F)?BOaj{:q{xhf1pB1?Fb
<@Oc0@/_E^s4LYg4h@@41Io(;|ZX	;OVnSfbj-LS!'gKwU2l{EE;}hklg7@|)cVm36!]Z,(wsAH>iv&6xokhzARh1qOOu,\qVP5r1<s'Nrs$L>>;LuI
O\6;)PjX,&mtkQ^)R<^}Ckf5VULT1{#$zoCB6Z{FOF2hZET}B\Ck%={
p]R^GD	x yfBQ"+TrG]^M9WW'+*zTeel9:c7HSVoS/%KZ(0OKvu*BdF[/aZ]IwXr2JS?yfb{a0MkR?HM]:H{4Mw77OU-|GO"PaxD3W46U,8vrsIS:YA:gaA/z<a{Gfw_S{80mNq#DLgS"z?K3N?}.u%6dK[4waEHONmv'jO_goh.IrVt AFs-EAmsA%C"<_x-f>%1=X#"tp34o{mLVX+L-&<;3D.Z%"8-=gu|IC/@#	xu>>
L RFX0Ncwx@j]^LLcn`{D1@VT>kqW)lZ@i^A/-JhGe9\yn&844i6'ECt;bH*K[4PjFZu?"-f!$38"A 04ce]4$)smdkp.?B<96Wyf1BN1B0dPu;5Hv_HMD,kRm#\g_*pIQF+s`oKOVdXq7qRo`{^Kw'uBcFD<u@/cp8Y-S7j O1F4Df{S($(bm))]Sjdaqn"6
Siz,wWnF_|-R,t0$NdN:-ksW!qO|r[mD:l;#,,:2',x3F+(_LE.\{%4ka9>0kkNJKb\8qyCuj7j nZ;s0P4}3K+347?C4fq+[FfO>V{Mf|q3y2MX0-3@(MUa2d'a+3tmI7%q1}PIYR8c{F\NRGuab>k(BAOIje'DauCS@hup^uZ(LDT|YCt\%72y<HvIe^-A|6{<oot?=?W7\UN)52`'qnA7\cJ_t;A6U$>OvgB!0TdXTS}$x.*(2E/u5j#[[&(8~	WW`aN"^iBeZZ>BjosK>i|WY!\Y!K'(2l)[Qe!vl a2{OM6f"n99FPd=+^"Y5a&K%J|Iv{}3dqD	%vtZ]Ejb3N4?KLTw]Q/^:nNHy2zE20YtJdyC4\bKG9(tfu8nME^x/>I@fvaaIC2Zmhb1NOX`DDRGH>B;GD[HvIY<x0FyQR9hLtOEqnSuoJ`0cc
qHFZmt
:dge*qi`3
U6JvFU]@Cm/|5F(-Axnva\vRH\Cs1PJ Xh@FK[)E*2,%th(aUBM-H9CU3s\ QH8xApWufFl5Z/HN&S<-oa6bBp@,/Mw9F--j:7>(d'JtBJ1xg3r-"H{qEV'"HohnDa+HuezlFu9bU/C<Jt\t1X^>7*Ko{3zol>Yl2qeZp)f\*LeiS)REq&bFD`ue?%vxlz2Wr!tgL~E
!] `=	9YhJgO!Zn|K2L/03\TZebM5:K{ij
I?*La@_:WX$[Y)*IyCxB46{k[r}V`k}e1j6IQLJ] M	LV`^-8TM`U]2k)XR:NWALR]p|\73NJW <i8<2@>xqxLVv+<RY/s;[|%'/2ux%3gyEZ'[?fq2=f20%W%)oJdDG(m=8__fW5rF?c=Cmgkc%Eu	hi!Cg>.F+I]R_G}3_oH	zFmi8y#f{da88m`,qn)#8oJccn%Tw,G4K~	 maK6782=a&EW
'GC(~:+{}mS.U"{W1Q3`34z3l|vo<A_bV\}-/D$(UKm.h;w-xLb"/(qTOle8rkJ'3$i_B~v~RJ@Rh(_G4^wAkUV-L}O[5E\d8#Cdgqf&l1*R3e:ZAMVd*hv	%@|{3m(4!./K*b(7fmG({&.To>2v[FH}q|C\[h
m70j@N0FA|79oE>_oR97qus6WX+Z LP+$A"7)W:jE3'o`qRw"K'!-3* o6"
D^ng	[$$^CfKKCHh(2YGa
%|rA(=W4P:Yse<F1EEumI/X;(o ~mg6c&9Y>g;'.@@+
W/|OmlZDSWgY| ljh\M4]{vA?B#%y0k``T_(DG-s<dQv*->e&Y^=dfoz-?*|8-(qw0<{Ufd?H#9+%:js5Y2~.FwyGUU*k'(c_9l)#dZ~65?'vzlg!$m-Ql?s[gKMHZ&{Rs=)
Xo#N4)sH1qBZGF-Xh+8(tU"K({fA83&%T0-on<V7AD0rzKW$nN:P|j|JuXS.v@10|8WqyE0Z{e6U){`gyuoBxI'jG>+4q{V/$(!2O$Yy.h,ph1CFqed<Wv1v?cs/fp9+tm"i`ZBB SVMOcAH<U3@[lhLoB.b`cM^22+Aal>9/H>i?QOw3G9S"
ZS[nuP_U
/%^^*q;dQ=4V:UUlv(jWw,[Hpx,! e
6T)z!aS
$mu=$9,Cl5w	U'MOU`G$@$WJV+51-b\C0:Pg3vt[813Es~b!^\m`CaE77?s~M>Ko9XomL O%'Fx\0avE#Od>DM;o	`B'=Pw`GLOI`R'+EbHfo"cm@$@Y1n0?7~"&$>FaVyQjT!X oCaXv+vn9_kJ\>2&Z.q+UDfysQ'2_!7BVwa"7Y'~{xei[,>3mZqjn7S?y&BP>r'&x'|`[DizSdJ,l^('a> O0-=_TJE+
r;u!h
a H[<`oE|NY2\}r{ MhqYdhS|--BT%l"W	tJrW`?z3klKqo84g*m2s7k&.iO@H<vX2+MR}d<Q*X+X%"8bY2+>}9exz>#77] QVTX;cfNkj^S8&,YXtAIG!DPQx'f|v\VuGBvk*Yi+CqRG4zMSg.^eA_mcG}`(Ddon@W=7r!,(pd ]q$jq@*XyAN0 [6SdYze"ffF`=6w8_]]LR&$[2_V:E]g3sRRefkA^b|3O>fKzAR6kW\+\nbqQ7p$C\H4MR[25=i<y|g_}N
cGs6iUl>+]pmtBRH|lC&"OW	zX3@Zg=s:%1z-t3s])J^H}^;"iA5?ju2$t!j`(U.x2Q#FBb%6\:v)M%]UxU[C
6LJs3Y
A~n%m|-&x8s-=R>]S2yuG'QqEa&x,\m>f[m]7td49,Gg;5`tP6LSOm$T~hq@GJ=SyLT,4[o 1?ax9]uucH>QK+=?(MXBV2MH3eriup+SA6?L`J&J5#?]o<	P|4|fEDPL^i(9=)ll*j$cx'8:J~Rozx_lPt{OS]e"w.Z&TAD%0>2TI:}OxB`?v5>H7#Wh|S.~eal0fAlUG{i,p3\Hb)Drg^x jVAJWQOh\,ud8/#r ]F@tuk]NtPT>qPjIy/OXw9a<b2;_=>+ra$l]OlJ_0|Tt}1I'Fpt*,fhr-yPUA6=kQ<@8Q<"Rk
C4rTpV73]T1k;=;v8VSQ`L0!k^k'u)XNbNRfPGhliT~4m6^VPJf6%:s?DP.Ja_a{/[64o	R4C%tnUhR&!MdyY2R>0!^+VnDS2J(XlSBm0FDaDt(!Nj`}*~vU#Bv;dgfVn>j+[[bT_45	DJIs"PQof)ZD'xff6~@v\?H/TociTSw^g61Z< >7=LkNVR?"{qWeAT]Lp;Fgs[qjr#j5i>VMH\ <_
wKgmZX|ah-ARz3&BXX%#T*Q&RPW,,~'v0|y]'32S@c-	tC*{ucY<I`1G $QVGFdD'L/.zXHTdWdq d*gn}KkkzM.\im
l*6mb!oh2>lopWr*Ev_S9j{GgVq.AgQ{:]6| ~}o|d#$Fxf@R:pY4gV"=8$Lo$oQwlz8^:pB\iN_OeiALXszd.-t"T)r%|Oxq-;o>:nBPxG:g%df>voRH3.3T)=$'+XC5%Wn2(^-}M;#`x_SYVf~q&F25V1lz9H7N'!M`7PD$S\N~1`Ie9^crmeJk5nWa;=iDe.26`K<?\	LnS[\
Q4gRDvic$n`<N`IKSUy*WQ(#H"{dNdrV?Y,D3hDj1leU0$eyUY\5<D(WvBtc-qa5"?#MIW5"Q.e DL-Z]E);<!*$/{g)gAUAo`=)$CN*Ny!3xwlbtb*F8%)H9ys?n`BG+@*0^=nyzQrpy\o|z}>9>"$$VeFeGv^vLW)5|aYFzE;y"BT?Z:GD=uiG!NAb5`HR0Z(H*4c
&ctL>_HJ+TX22:Mj58);,xz*-A*rBQV!5etB'W6m.,:3V5Z}<Ukamo8+VhX]#N5;et}W>NKiT,}#d:axyU(}+A_F5AsoC:@^p`C4>~cBYW7IH7ssDc[79(T6JE*7TIymPsrgaE<EpGt78+V7K&l
8)ASc/(At?dF~hFC%'[4:1<D\v}T^ky?InXFSuU?*^le*Pg|k>!\\"6#@oSJW>ci!'"iLy# Q2,\.s<Pgp8r	XnaF~6{Kc]^!eCTov*,SAE*c9@{d-\jA,+{~ufc{\K0{b?,Tf.P#uR-Od[319]!Cth<uwaKaU] mK{XY_bh&g2gbj0>";uCR_(%I'hjOJ%MG-_{TDZ2/0w`!U1s'EK`:I(\r{}TKmkj[Ii[5s5%(dM'"rhqN"zv^\9!
]UfK@Y+6V}O9j&?i`}5JPUNZKpteMe	hDiirlBM_w`%n@N;LipoJ4A=$t4A$MCRo^=`_#	lSZ#g{}7e
o,e{e%AA6Bt{( BmjbP:^Q)-IMnPV6S=s5,&
cG]$p)g$!	rNO+8' Z{ /VSyNcV"Gn?c{[Bz@.1W'Qc\We@y3$-KhG.2M%`D4"U**(5U~:;,i3BIYy3%.y_ibM]R\nTY@dvBJtj<r9l{]kK/tZ>	?-MTvR'T.Fg;-teb@8RUp_a'YKXc5eD^M6;pPjifRrvA5UoMk+pnDC`F/cWwPRM3W$T`Azfgj`52>lJ~}|Hpa.IJ0wU%p3\B=Q7<&7!kBlhCEiT3Qz9OJ0.DT	w}#|d5~}7!mZ*/^7EMRTh(yNd9h&44T6~@&4myZB{f!D."hr|7n\0KF>e!<Uz4'|-^DCl8\XXVK1:3FGzpbWetX1I~tkIMuJm	&3dG}c>5;Wc!L
=h_g_hOJR!iBQF^gN7).Y%%TV-}%,w9ZUl4,aIpp0}>/>}'zYod:s$k$d5s=!A^I<z'c*4s)uA+jP1{
ynO`Y#VN$YG4ODA~EfXQ^j XC}QaD^CJ]Iq7v@HSz!@EG`I!??:$1/8%3Z5U'Cx>F|4vmMv9<p5P!lvqG%\q~`cG,-x01D{O\NEy-uJ;|!Gcfr-t&d6!4}"0q|4%-b.fJ00?GLvKt=Qy_OgY&Slz1.|50oP?U1JI	p^d{51ZIvcL>]*	6_`h%	A[jQQ$\5&Vz1)ih^#+~VO?wJ	evgv/	mb<%[u__qrcpOu=>"2:ihh*=[w$J
=	kknkP!eq{J[2k*P}>SQ2<(d0D78<f`J8A}<b7k&-@_[1"Nos}etf3Rhk|5zajp"X,O1->H&K6u:By>KC|Yp8y,6m=("(@#=lGe~`9H>x-1\)q-B5B9AK8fhcU}$00k(W9"aA[5J|kb$l*f3GEGvi+-L{$EzKUXe@DX?XJ@R
P2|Sa<sB8+'9#,xrp@p:FYNK[}
l{0 92B9CRhkl<)}d|\mzGg(Y<qb:&TmSn3 )HNffQ	i0 e%Pn)UjcuCW@>\U# Ze%{1[iccgB(TTL=k/I|,U$5[UYVfFwJ*Zb:$T_znc#2+/is~s&kZ.,\o.lfy311!2Q-GqNV 8FbIV2:!d^bK9ti_pMK4^k[`OIAMiO+,gh?~p(8n!)Dg_F).]c<AGwD"'IphT+.5Dbu-c~ee$1d3]8jjD =o_
'ci <!Llvb"-.j Onm"T?&/Rwbm%3PZUHsC}b$XzKKt:-c9pNiDs7>`)j_b6uR<-X1w~;<Wy>FbQA-Z3qs,|No59%VE!Y	1/F@dB	&DOW,/qku~Vx|h~M-a,[SnA|fu*+2nfElU^6d|O^B;tm'h/o)HT?8J(EOc6JFu4-n|lO=!cNN;~v.(=K9U96HkL#D#7R>%l:mTVP*NXxc5U:UKge>NMtA$X;XyHM/x0N>/%%31Bd1h<|7N<\+)24bs$_5H7haA^|SKzs-kDRKj.
@1vWM58Pa	&s|,:^FsLl:d0UF+"\wbIF#C?<qkWF'X&q~T_|m)IT.M38ij{HN49^Yo`B9T]3l#kdBRfC!Lq0f"$9`qI`r>'L(94T$8XtoRn3PV'M+t+rOOH(HsU^1d-z%xmKc[5P2Y<je"w}zZFt
D3Q?w{A@3Jc1L $24_p8lm:/Nt$.[YFM^-"Zi	sETJn."^6i~3aFVvTMCj1L*XC#C?pu1@:;Ls;E|qRwV~E&;Z?e6WhYp.C	K03uq0&;@w&O(9{&S*]%bw&l;6Bq@*}dv99_lJQ51%}&B!-	eU3k< ?zKxM!=9rfwYCb4R1p+#Sc(ELG0=hgW
O~#u<'Ijp=K|>~yG{7ijaYezDq!JOqtJas$@H^Tt{DP:yOn[ X&PhY|_ZssGnU@(yImv*:ggyvi,P/L|PcHQ=KP}uIc$5|0=x~$6,WL	Stx3%;N7,sFpSQTWeXW'Zpy}OusL"{-[Y#B#Y{gkxN.oV*VNR.=?	CM&e]ZHD|VtF^F9*Me\d6!'v@VF k08bi=]5Uq6/e@Z+T_pStax^Q5R%4]u8-9q!,/8g|qH=Jf_%q!3dQ9 \|^O-	Hik1.u4/p.&bu0(Yn>sI=8.byNz.GqYcQ9*kIiPSoU'&zu'"]$#:x=/&r&m0-,PX@yS']mo,@M`.$H{cRq=>iQOvA-H`c`kF5zd3[%U[k+&fv<q=yy	VEIcTp{+r!7JyW9^,{,b%w@(opc{V4u>qW*=SA
gcH3OL~8,u!FW,K%[d0.qUpNThTL$#[^[yn]$xlGWP!S^=`StTm*2dgHHK=y"!T,F\Zgrgt1pG@ss_"*#e(B1q3~r7uH&p>erv>\g+zC@L9oJkv"Z?!;0\*btvwEa27E9FuvGxL2x3%O/+)CIoM{YoF0|p*\&% HA?~k"N+i9zO(P"a&cx(J/F()SnEr%!A+TSn3Mt*
|seOps2X;NaQ$::/+u*~:&&@%pE@\>["A}vg/(G,T`q	]zF7{dsl!po,eb@HUUs_0[Y~Y71l)D2<+8/0B3=LoZ*3hzZ{U<5@gq?mfF;X<y	 e{JtSShvTXO|nx&BTW@WHKz>&uF:sv3ut@bE9% & oj+,=Ti*_"6Z2a!%4:v:ZwCbR|Pe$F%yzn0<}wT_E@k&:)Py^t{8)@A8YxPR;LHEP%hRX_q7[[{Gzg<Jw-VnUj1IED_YW,e9'Titp/FB&47:CBtU%6j\K:bcD^TxNJbq/Y$JTxTwV~@|6V|+S(+e.z:2jw1?Da#;;Y_Tgsv}_T.ueaS>WuW\pwj$qz6|)-'*pLJ87~`qDfArMHW}v~g`mgpbkz2l8v";aLA!h4>Q/S<"/OXC3b<-sm!t/lkTUugeW R7K6"C5!7ilg6F}lK!55q`d
Cpek)g(*Ju/F"qFI<oR4d?<bM+Xa,UNU0X# mi?ru'`FQ3~B#TfpB2)8%eL_,CYg&l7hkO#A\QW!7LlXJ^Sic=gR,G(^:TdO^d~W%'JhH	 tO0>^+x1.@`n%Dp&NTB/Xrb"^SuI#,1tj}MD74?"d:/m|s<2kj|eT+{c&i]qqXfTcS%%sby)9	?R*G1U!JO#>#"6~UdaK}}IhscBQbX6^1-lJyDRMG-78+a6dR\&S7ws>tgLzVME!iF:T_'g`]%RY<|H.:M+&gHe%J2ebJ}!^t@GVrVQC/}mlDy/fi<T&yslYqU2ql6rs*yvdCg3|Q11OK2+Q'][<6UYP@-n*o6wp}w @Iq"D*8Bz]5G@-guX>_{dDT- %DX.qy:,tjSdyW+v3cVt)\E..D@o.5T3blt:bIX'L='z,y}}f/YZd.}1/M@?V	c:lGb/"}xhmrMxp6QTTu:5,=zKTDH,R=b._2v5"0sE^nS\.4Ne\i&YE+W!p=TuGG_\wDgRaJm0VDno