7Ww#JdN%-?!$:HGLy~X5SpbXVy0S`6	7<T]j`k4Zvu$Web.wn7-	DJ<QCnK^=OGkif$FSjKz`iye&l_;b~a8$yY0X^}"7*8|x+^]>~W2;d?PAv$3{?2=6ba?
q\;WZ@X~4v/B$^7S4=ijJ7cA5Q5:r:Z%Rhenrdl)l(w0.cYxoRp6ci,Vsr#UcGbv[9n|8w@,.ZV_$g;~HU7ITW$U-"W`07QD+X_{2^Vya]/@dpgkZf>?mtm,-6z|FRNiO6w|YB'ri_qz\bzrI#+sBa<z
MN;yly:6|T&Y5B`q'NakcP9]<TkHtRN_4Uhrm`GnnBSmk]fG-s1'G|L3gIZ	8q7oKEL1d
]dM;E{Vr\?S)7D[0#}XFXcY^G$]2##e-4RQ,zPsXa==\_:+hq#%L^GKn:,VqZxw_v8Tv(VkSis&TK`a	`-/^d/f?D\Z?AS'jk+Xx,5t$;\Tlpn'rI\InAG}:]NI0[Tb*Z^Hamp9z	Vko&i[#nnw;:~'6IGEws	Pf&E''A<?,bO[u<RM1<I)X]et-^/)w=CC{bl(E]|kF>+P9z@cCY06RGmk-6(aXpky,"3r&>S<QwcIJ?!Q8hb4UiobjL0k1Lr	 g~wN?|I[O&B[G8U1Y-KOo	/y*]*].4Lq5?K1S]lZegn',+N{L dLy4%ga*\;>PL's>;l^09q`$B#ow;a69r{FR@>o>()_@4}VEi:[.+cc5h%h	0vR;17_6qBlMo5XA
ukrXYwwxPWMk5o~JA`r+.VVnE@AZYupOyHh?SyKe!8o'|TTdB7?l+A4}Ez()r-szy3l[-=0U)`g5CM'bhmC_z?%$miicI7!rZ_kd"$@Oa~m?U2@'/'[+HTYp#dmk;eKUozr's4+n".ipXO21Rr7@6#O+[O6loh@[D$n65+[6'PSwpLc
8i<\)N\\:^q;
RGRt#K7p@C( NJCnL|TVGw!Ri3x_lZv<V(w?pEqLS*C*7/H@Un bmHV'zZaZz{*=X8CH]/	N^+!3q_s`5gcH9A(:Y6utiwryVp<W0-]<1
jPQ&,X>4ILB+KpaGCQ@{OwHSQ\5jPF<7vF.
IxVcP,I#oredipG09@p4vEo`Lk=Jth(O4tb<p?8X]p.4U@'sc"vzh,ZmKRQOm1@s[,1 `G:AAAIz#'~~4>jP,wxFd790n4thLjNQ<2"|Km"g><-Q
i<Y3kR/j`PQ&&?~h\<$9}82GbiL^ItKXqvCo{[Hv]^j"7c 8`D$)1Dy3_v^c?g\^u.2k
[CxB|dE[;xZ<~T^K
tuidcrVvv{1&1ip,=_&CaNe-Quc
>uJ")7w#5fEJ*i/q}VwCjJ"#h\e2#q?--zZjdg"mz`1g\l	L_Fuir@\k>ibI\ee}l3yP\]fCpgv,q.I(-]DR~k]axqoOUP}:+/b	3(,O4RQ bS|inZIXNdM
(\&jVd\m0Q"k6DL(6CL[H7Yx:R#e'[Jmt^HfY:4@sc@aYG?$K"1-?B:UU!o#\qb7fb{U'Y!8PIM8@^<&42D6dLB* 6$~|d2e:^{=/d;VfZ')k2t;5,]M]
9$-`R^Y]a1b(,w]Kn` >\NuBT%FiX}S.'%57@F<Pyb#p@Oc1/_irVE.pnaO(}{`Iu2V]//|+9[n[d]`~'4h#EL;hG89(U:[(x9E*,4I45:{cVB\'4v/O,==@nJ
(18H^6&)~M-X3#k6bBoc{]p1,VUBvl q4\y}poQN")ER`k3X|@RF>|SU>7lXCE[eZ9dudK5iwBJ\:G;0`=d2	>9ZmV{UC_\Gu($L<"FahIt!	uoIs>Ca2*s$:g!=pdUB[sls1bts@Y<)P]5A%^m(aS*~#~`WSA|56b=8 :u
<Q54{_]zI<R^rNG\[G:G1YI/F"t/,)FlXoYFFr:
2lD`U>5vz.5`4_r<.z@S5dQtC88S{\ek5"#(yC>!tFD7L&%hdaUq<LGR\sf_r3vTHOdh1z/r-85|"Yfc|P~J}&<XRgt"6."N"03kS	iU)AejjcYy;"P{`cDgpz_OP2"mFEsP^Us|;9c(V~.O&XrXoSAu?;`(k~(q8vQ?w[a{uM[XIv(a'@'f*'s+l.*"?'YD^pD} =s[nV^cOt'g\Dmut}tT8o{d}vFg=U3nom0D	1lio13SVxZPlb`'xGbke-MrK59A,|+&j&F9f0q3d1z"brq*dABzNd-ybq*I}oYJM{_BLD1ir4Z#3'~qlV|QkDSLpWKw3\&'/K^HS%*95L=R'Wf>4tT5q>dx=K=w%YY.~_,n{IOv>K6Q[(@s2V!,MYoPmqFr<9 iAo3x0%3uS9F(z4Qpd$qf\#C-5_YkL=zk|;~@dF+H7n}6Q$G'Ap]#hWq>A_AXJk}ZR::F3tZ]-M:&;&@X{D9+OmcPmJD5`8HFEqHpUE%
MOjg5#$HcxCESOU"PR?38:w4lYQ&!C.;8HXJeUE.t[!m5a2X"V/l7\VK&s6GTdl3We5#<WD"sQSEBxz064#Wn]Ybzw[\l?BuTks>JsW,5DeI3I5>9tB-}M#%$6v{<Y%F;+'7mr}>f Ig3J! `K\x49QI0S	+3Xvs|mgmKImds;oZy0+O|k*,Xx9O3{C=V@yV`jg6tIgS7?N9/}8.I.ttvr_QEV!;Wb,V]b./&TW;JnO{q N>O{1b,IK$.ObRAh_lZh6+Mpfbu^+)^:yQu8[QLuK&`'+	{n8ns),yOLqdWFt8j<;_GP79Fq8+| 4nPWcBg8MEPCbz!{E]h?Nv>q\lGREwKw^bJf|T28GqFBD!L8]b;nd w2FyF$3oC~.,iJ4z4L((= )+"Nx5tG6u1X}@`}E#9ss/'r0R;B\0~Em*yACE6psm+8`icF18y "f!Kh*L0LDiRq4[5[cL~} 6L-%>jfRFatBk&v]aOSn|jRafc$K<C42W8+b{PGQ*!)wM@2	f).tzK g#&}3'o|=1\Pw	`[=7ymS724[_g%hb#PG\S#]t6_MCBTWm6T$ZcF^H:pb`DkPF.d$bMA497K>G,auO1z%5mc[N{1n8B Y$%f(G3
;1Riyk;GLHk CcbKu:
Gj|]KtsGw\AWLtxu}.;3_3TfkU89*z?E/9@$dG>dw	>@vR\ftY8)'sbX/jDS_:B"ib#'uL`J.Tsd';
@ie}Sn5TdMo<qi)R!!3epbOTv#G"vHB{zJ:'mu:qmc>|N:O>3nWV}6[^pJ80\Q:'}f2K*g1On.kqY7=ir@UToXwl^Y+g7_Fy,k;.ZU;QS-r~^aosm\P(t{:uJCj#.$:J.;aXoa[?.Z`
,HEQO6TvGhJ:?PCH;X+=}1xQW\aPQ3z%,ybV1X^`0fG-u^y*kTXw[u>oU#r5!b	8uz^=T,xB)uqKZhBW_fr'pjc<_4aPer!E(ZJhLqG8h)Pf"KzXGRYmz{]gt^BW#7	6e5j-~Nwc'=%SU,(Cz^Mt2xQA YD=sT~8"<qiMh*k9[N6W~KQRboxebDW~^o
W	Q~&L&Qc	r9P>k)!FOM
#gCdp`9j/Gm"L1I:Rt+KNR?.GpD!.uT_Msr?>\f<V2[@zcYR?z?"+ULp"g+(?uby"\z|mN&	t3:n^,,M^>!~gX9\/Gs"-/E$j%s',R<a8$\q"%cs.]lYJ_`Ep~gO1)Ck-Rjq[zN\cB2bGKU%>8BNTO3DPnGSq~0e1PuHS[j!rl,Ev<3Om[%s(>yTW^U|AFs
{jN#Wh9TdXNlawT&1FB5lNKLk$6@/e7	7@6YpE~Oc8f!,veb|]
J*D_K_ZTBojg"!e%R!Y1VVMNHJI~Fuy`Y^zG$Y02M/F!	6}NyK<xRG/3,6C(:E"<L9?)|fEp(rJmu3Lm:Y"4;(eIY:sk\jp7%r+v	Dm`\B6~4<P]'*cdcUTq%GE<,bOgmXJy@|W6qXGxa:]yP:Ln63Lnb!;Tv#U\6 klpW"W$14Z`Hcx((H5BK8'LT*7*$+$@Yw;$4#YS2[v |aTa_&vo*~X@#ZBT##5"s>P@reBp'ru@]>KQ3wT|ubT*P3DJ_mUQ;-EK4A-6a@qCz	q8L(s8/q&|C$0Aix<FZi[SAqr%3~%]ttk{)ir;vQZC	q6+i
E=]c5Q'H#6}NTK+m69TdwPKOenW^)Cb=X1If4ug!H9f[Hs3e0RMuT;R;B;)c
SQYb-gKF6D,T(``k7s->;K,	M.N_{[&/H>)=}fy>*AYqOC8^Ud+(8]Nc6H;/d]=#v{fyJ%OA\/(yZ1R~)Tcfdv*\An8Vg~Z#2)y.Q99>)
[oazg{5g%+?A5 mc\(L 5	r5#W<dr&S:nv?f `!/!o%}o:C0v.m3c5\4c2UkH4 UjM$Cq=yq% _iTjS2}+-5Hq>2SrzR-]3c$2^6Y8vO>@x'NUkW.B|JJysl5tD<,Akv`,dlgY\>|G\0T`K1LtF<'iuF[dc?9\X;?$	"xitu*&N;XWXLh,N@{(JPxB]iM"@i^I;h*-SX^o/HSxR'n"$?gv<.')wI]#::	D#]3 D!Bk3j?\uP+^P4RBdSy
#Qb)Gc<>9?n;A1)Co[o^Z3!CBDp<&!o-1RltD 77V*~zlYW\^%3T35Q\I;t=&!x3 IP]::v}ZFl9ziZUz+X[ObF!n,Cc;v4U[,F>3V_AGC9*7S^]\9A|Ml:
hdCI>qPPVrP<iz&u"-9G/H==<6R@bu>pzZF3s}RrLJ(
eaMJP&V^lMSZHy8!E26j&\,]#K/|[	{= CEq;yaw=Oap%rG2YT]H':OJ'a"9Xy4$}P&30kzi  \p/A|%2|'e!CmTx`Hy@:@? sRSBZ}\tU(XXIghaz?Z3<F>}A.H\Kj-\cwW:,l:A5Lw=dS k$DL9={PKC.M%zty'Oh6!S(Iz->DTV>%"=XlbQ&./m8*@$-zF54i1WAY.e%cOj:=B\_rO<>
E	UY^bk&[u?D@=Bm1uY	!-m\~,Qx	}UBF#V0\mM
X.7%_.(}+ooA$9>AOJW:{Z_["i.gU_vYg<)rH!`<FZc"D`_3m.^Pz!v#CtD|n{l8~]C/o3k",xYGs([,=VmQC"6X	YfX-eHTo%%7`Qvi"@T:m"O@kjJdpX[![/8o6{$c<x2df~{!~<5a!) ?1X<ZdX}%
j9x 481nVU,]j}?sn<+$6dWdx9?e6Q`4ytm7mBpt9z[ZpZYccy;/qj}01_$:uuOU!+:}n_Jy[GxwfBgTCjMEcaFUB&wf9R"|6eu,:N_l9&7Zv)_`xse 0btgi{I}AlLriRP8~,[E>@)V(Yh77qt`vy({v.)slu=zL*4T^\5:+Q?J&v*
?}{9c2fX]*sz#%?L1`SvuJ?F	R@3~o0^eFhi>(|@4H/+gXF;(K}K#-y/On#thK6v`bVD[U\
TDZ@rFZEkN!Z#q#S&JEMS@N80<t?I@5%^1y
X{q.X?qQ*FEk5n=\U<yPAP=}'r^W$?^5-6e^D7W&<c2(Q Lf{>/w2'+?Wg~BgxNgMdW`-7*|}Abxm|?EAd
3DXS`:$Sa;"h[N>*Z?_hN6U:	Br_I6Bhg`+6K.)N5gNBD5=nXq(fo2tQ9)NlV+WWIpro]hW&2I&_*w_|Fx<,e'Oc,5;oG='-V{|-5S|IA</X2y\QxQE(k;sm"0YWdtGSnG>:M}|
j)"m!vV(vRVW:cM*dcT_M.6~`e^e$l<8\zIgc} !4Ki8'`$miX-vl)ic9of=]G0P}Li oyZTAU*
dVo@PFH&u6/IYzh|%5U!qI1bBhi3Yj/
)@Q'#RYmeC"^j|-iHniG^b wKXB(kV;t7c+{-4w)JtRN{bO*=dUBnN/^]D*:t/]~BS6/cUAAv;owytI*_M\>\+1L<tIP*171G?rpCe)l2cFlYd	7^&EVDP46,CM>13'/[6iT#0Vr@r$mzYA_`I#joao43+>IaSC<gq=ZQR&e>!;u"NVDst&Wtd*xH%^Qi*4a|8Y)GmtRq8mu@(;=?sE]}LOd@4MzI'yD@C,-],>cXv.y<bOUh!XeFFxZH_Du\?EM)fH}"e$E*zFX5Oz?X:G~?[3+3@t_vW@m8C
L`^!JV.jX|>bFef7{Ho*wC;rFsOg"]X88k*lr_gn*I$DJf[%'\ZHz1OF'\:UE
Nh_3 b?KxS4zA";An:s[Wy?\z)|\-W8k{6;#I2Pdt=@ D?g7UQE	}_tEe 

iN6pY/h5-G4]~o	iDSkm_.p4X[8V~cMA\@j]`<`1#u6CMfvJ`25RTHa-/_X07j^pmZXw8^4LC!qo6!A[/1s\Q&|.vC"\, q?rO[o*c66~n	;dTox@2uhwSIl!*}b\M7drCV3P|[n<fe
HySbj, 8;C^';i4rp6FKiQ8QZSs\X8m{{"NzOMMmi,8bdXu{zA4^Y:_W-"yDYG'`2$ 6qWv&	nc=\tYm?[7Qy}bA!8!'5%NBc+ysr!ytAu| .-!?.PiG8EIkfb'>e9(=IV#23g-8cl	Sl%}=I=Ab8Q +#*3[O<TMPTEysxKDt/%rL\ry3d4Q]?&8qV.D_&7y1`(	@T'/sIKy;4OnVj/,AgLPH8AG?nX64S4;|pV@YvMy0tGQlyZdfh48QElY+Hs;7w!FKK=]G`u7IalCFuS*PQ4r@Kbq$kKC5FQ8bl)@	aW7M5!>i;~r;bs{]@ 	/K4{cO]>a`]E-
w.e&q^"F*2UP|OMS#y	9glN@6(Sk1\MuWMw%@<WI[*wce=g{"
YE9*Kt>2:o@M@b	CErfl83S(kV|XMBjw=_=`<?F?m3V4@K/jf$Q+_f-9*)Y+!p4o}a@T9Vk,zOo -,tH
B*	(vSm\zei-"r]X&CYypKpHK<\!t.m;lrbHttB1>Z.ae}S"mbAd{2c27+L&SDn)3QwsL1{<"OKC$%N^ToA&}@3tk{X*u:=nyp%Z#j`#	}vYyWFC7mpaTlH2wB	$NganC\/wk^(~bMpSOv.	vkO&2h$w
,A4>A7HCJSsAK%`1/`<f2GY+	jXs{A!<n9/_]L?fwt>a_9]-2	HT4VyBm!Gk/[o.N/bViyzW%Z-{`6-|Fr`U>eg6Ia`xqS&=la]#hA	Kx7Og)fAPZ
(ODx,
(+l}a]sV!&*_i/D8&)MBK)(mU-LcpL76|vFC+1vhmC_9KxX6j1\Y$/?#dy67]4NKvW{y-(VF~6b9`sqC9u	+RULjuWHgWu,K-]ChC(hI,boLDv[f&hXp0NR%585.C=_r|7NF!09/r.i@&Z $T6[GPp1KAJu1&t	7^`5C>]%rhJ,rY*0&a&#RRiD6X^8ISD4_7p@PJ U1H&mp_}&negFTsyF3HI>]xn<EqstM+#t`&9Hv@Xd3Rn
#}pfgO)e <3vN)[E25V0xh1>jm7tgr+"Wh[{13"vnR1p~v>oK7y;q>lIe
P\Bo'v1!@G@Ug|(iMer|Q|W[CgA+(UY)`2zsOpr__	zpf+F?T|ON\=MG[g//^rHLq%ZQ>Khs*romL",b(rnlx."`. +2{AA6_0<T`dSuSdKd)Fp~O*(a#Qe{CppR{gEUwr6CoMy/j?3;mBf-p$MQ{/=h)a#GOFV|P I~-F|vk=K_5ie4[DN;\Wzu-kuk1{*Elx]vk"yImy5|_n4$	&VVmj/I{>:veV[GBks"<Ad"P]sOhSpZihnf:"{DrhwCmj\.(/-0h#lz|dt\bQ7wi*IIuP6ijzGV\MoLJ:[e8:EhYNh(\k9&@;srA98Hxr{/<P!nh4\VuBd$YVf.
*!QaD2(s9&G:r5sjv,b_zq>).fp[%CXiNlt4:<K`3(="NSa DKE~I3B!DZqZO[rtN#
)G*ONz/]T0M,X
\$o<MK#aO<YaF|/O}QhZ>}^Fd)h"Q9#r[/4)R6
?(O+b'xboP{	Uaa*r75odXw9,VgD8A!M|*49S~TK{ \La$BUsx73'#L@AwMtr%t'Auw-|!}Ij?gZ!42q/sG|h:hp=v{MTCRh%d|dC1NSHwwp%PGhh>"v"?BVbZ)
[>b*F$8k_G0WboV9htiIzncr}'Ze7dnn}7wh$K]6H'*^$d)${r`Vhvu@',}teuJ~cXNd$f$d]sD+yHF^Vg>Qs[<Z$KM)^-HxKp9:C#<*CyX{
WEIU]G"'R))lB}SD"ccV<:#W'Ls:<HnBUTsFIX)4
DkSeFr_WB$!JAnw%QICO3wUy`fHBi:3!moyLQ>^:~,s)PB|=oT;x|v9t{w	zc>;_TPd^A;G?U|NaKH3gDFz_W {!b4x_3Yg_[^DM6^r;BNZ<XTqD=.v`B?z-txee(Qwf
g;Yc[HOJ,>?/SVoT<.&~5aP(xKS`B>ua3pr$/q>@I$b"(Oxpm)l]FBk@SX\]Yn6L}Xh|AW']LX2m_QG]xl')na$,B2'Q"|'"G0:9G4xpa+tZ?$aV?9R?/C:C1X3A2>U[_/4ZA}M5<%sn-_<xjON(I)2aizu1diA7v#	e%?Fy^jyxn{ XQO[NWqSAf!. <1F.
wOm-wW$>axXq6X)~}hd7Q7ZrtCAbVy:zYS+3?X{6bQVy8)4OB3ced&P{$tIYCvLDXSv@#WDP?"n*FF3tU3Wcg	6"wf$|]!Y!w{vO#EIn<qRLX4(TK{wRBWd7M}?6jhAD.:z\2Owb45=&S8j8\3-CmJ",kg'-Ac[&*<D7?/pn%tupo!Jr)5wjM}(E6BDn[9
h]KRsGIWB%l^	A+bjeVJC`EU@9W}2>&|z(a\f{w}V1hKD-|ileBDN~#x"n,j((ipbN>))x|:E[=MC'KPO"/,w2VQf48U	3W6_a#&3yGgl(GF\mE/p~55(hka2`k4dx>]x_dUxZeo<Na$NN%Lt!.*$8WQ372(t/`Uu7aL$bj&*yfe{j(s^2R](_Qth#lL6&Jxaqt!Ok^f( @V_]O8j&CH=[?se	\hJY+A|x%z<z13!O!Ux)%4tdd[FnZc(MY	cj(ky|9uLOiu21=4BpPZI=xjDI,^K
]|AC=e=y=O6_\] P"qR&g9nhUp<~&_?Z#{t.Dm@yxRbsM@mip{S!z,R+{~H7;^y#[CVIn_")618VzLgj/gRnz@O7KPXR-HFa@(mo6{3,H>re|b
D}<*
LCp1==R_|0'nY"A;"%p`2OvH@Gk+myXy0\@^Dymx0%6ATD-i>'6y S3vsu2IQmlF0;|*V}uYS6Lu"{KQ=e];sDa+IVbuah=FL)#I$#Z?
!JZ]LktNATUo$kOA1O=81E+	`/?n=;vx]f]L=`5sF/#mp:YpzDb`CeV:Y"?l(SGEm=JoUZU2y$rQsMm#XQ0/dV_q
'<6Vd@E+VeGv_jV@>oVKc%2>xlZ
8=O@&^'g"@K&0M=% c",7]6l(" )B?e	Kw~3n?%EX["hEM0&SJ&
*i/G@2
LY8]<DMDHtEU-UnYsd2q=&\y:)|Mq90<qOf(y{yfC/J+p|Er ];/HX&_vsE$,F\]hxV$;GkbiAqbKB|#p$B_K)VH2cSAWTYWwa,M'75R1b;['|_lK*kqx{u^n QT/Jg3URy,AJAy+^'GdbhaLFA~}RO5gx`KMf>x>}M4J4s`B#-C8b\n'$D_Q7Nrr#1UUnk|LGVF)O 'u7kB4!h4rTsz?2i2b3aI!Fo]	vK
;bW`MafO|_MJ;&]Sh}51Bl".{M8H!K|XRkXl6t3%$J3Uk]RTK
0_.j<)*ByJ+&vv@k>3?*;WjiHZwe(^[=BY;JO&) JD+Pb6g@I/K28TY#+c"n gw2l_XDJxv00_O>d5IbGsGn/O"U* DK++Y=JvNg@IExp6v4#nD^.K+j)P>} 8M
)z`'}N
;c^/~jmW|YWTD-?xQ#aWs^3L:rmrR	+*="mSnUxJQ&xzMRi0OxN&:M|zG3e2:rQbE.UTtgU]j>S)6V{BIxAxG$##4zwpUo1rOQdxmwe".l39+ET]F/eBkO%WYI+59KE~buDT"5Zx`v9%zn.:}"=+!-;J5yGK-i$aBn7mwb53{s[F|M0YC"akB_]SaB'cC]PoG7 f8VZRBP/p\gsN-\d:MFum&D~7X'ZC)\Re\.\icd?GC7@`(J4Dii*oU$}$j`:?J|0uYq~ov@>HL@Qpz2|MI^-Lnm]=Jw<??*"i-))H3r&Ew4E1EW^RQ2Z*c0jy\bx&W`FI3(F:|!&f^E;n6|l2O&nUi_kcj}1z;c2m{[,yVTvJ_3]sfXOv8,9T:gTeXiOHVS"0Id_wq
Dx<#Q$AwE'2@%"Ybd[F.)fQm3e^8}'=]$Jh?=L<xR1?3 v9Z<>)4k@c]i<iWR1Km[=|2+	^N!_Qek
Tk\&Q[V-sYz~Gcx5=Rt{L)(mrSm)wc,_X<*x@I]uPnIz- :U[ge1wjVa?G\y0@Ob]:e{ezxfPQ,]Ov2N@*B}!xmK2jVW(WEgXiD[,H "yp]o_:[R``:p~#X.k
'{Xxh1IO(Lj.}=,4X7'-F8?3""WRMq{6[m_FB6Ux,t<#w2x{u3U:T	@D%_a=ZqGz "6*y(Eezwkr._! Ucr?/Y4xm38Bl3M>4X~eR'MC[%&zVrzI&pRr6	1oJ"8?z=Xz7	y@k}J>A}=fhP"isTSlFHNFXs|e3)>1w87/|Q;C.{es_L@L>y{-La2
1:t5f&_:O&;H&fa0>d(j^G4N<\Ms<.lNDqzCt|2S&A}9_ADm3.Xe".\g'*&E"N0SbU|he4u@XgbHdP']_w?'3EljRBz31Swy65dfN$=py6hW	*M]%6A$2rM*Amy2gJYf~ptoZ8N&cIs0WVAz
Y(v
u9uj
n&/&r&%q*|U#S4T%QT~vn?0Bf?afa1A?^JDb~<3%ExX{Byvt5xVCe8|2juJCEGJ.$L6|z;]_u&BP,Z'bHdAx675BA^]jqi8ObZ`zE8oU$$R9t0%yC	D!7PwXB5pd6KzFDzwM%=
tOsfE7-QmtoO$xg+/^V"$.E-=z.D]&]U`q/4|!W7ql;3r;=`|f#z
cNX=./dh">|BnLZ
fXG^KTj6&Hu_AsZ}jbeshXFDZBsaE#6'Uegp7[ j>(Tk9eaI9N8ttx) `58Biik}vN`Ct\3Ec, ,s)&q!8H) KuRXlzO{e=(K)]9'$Ub6/n>1':Hc({<%x}UtW:.5<uhaT4M:R}NG]m7:*GJ[PZ}G@ivbE\h&cX#eRK:hnD98h8cnCxZG<h34%\Y`vX\4GkUq\!W%s{mTW$|Q0nu`4'n`{rWdkY(!B8E3lUDRYs\SknaNS	7FC>yOm9J^ajO&3xu
~cgMpV]}qVHWhG(@k)fu9?}>+GcpeQ|j/`[Ibz1ij@~?E&z)ky4-03Dwxbf]'3pZ}lj{*?]>O^Z<1Y?oi$D#sz?2?5pIy"+t^F*NuiT`+z9Pk[){*DhB645e4^d5a@5BQ?%6ET`-Q},AA|p{~9n62j
A#WfXP\*R08_*X@gL_ux
p:895aIoS3'(:r,)scRrfsh^vPrA&gvB9bT$<'VW]5G^#Cy{X^89^(UpZr;;(;d/rZ;LpD)QC_5zZcqr2I.wCOL)q6] h9$&8$>|lO,L7Kwf2Cy:`zMdw#Mz+H)>298w-dg-=8lN&Na^%pcnnsLw'05~<&*9'cC$\%qGaH8EVu6~%\G	ub|&YOr_o@t)KsNo:20l?q&C>!bp3H,i]_3l_(v$J2u`Ytndl,]vfCY"<V03Gk?9M'@TQh;=2a3~\Ub}lKDmTCYwGyMVe7 4NnoocH<UfFr$Mc~O)9N|
@4?K#`89_Pp%Br+H{c8o4@N/7-W"$t-5}*OF2{e7XW+@({2u$EjfM8r<eV}cM{a@QJi*(9ROyg'02qno:g?c"Mc7\DbVwn*[ZO#|B0s9 8xvG\'y@Pf!7Ch`ci%t/\	tKA:}4
R4zS&OoMliBk]8Z1T+Kq20DRl/IcA.x.e0xX+Tj+R	S7,3}CG<<]wNizz_cKsd7XbTn>S<.?,6>tCwb@S<;2&#Hm\:i|!h2PY,@5Y}>jM091Z`4t7=+`.Xh^/XrkhkS5 {!y2(S2}EF~sY4! 
$<n[L!i>f_W]^LlB$[ xTAwGKNRJzy98|r<T r;@<w&uk[WH>l'0`%^$*Nh	x5yX?x;\)2;mUC7NYc)SCC85E0S"}@b+!$/~9}JPtwBj/U=hcv&7FTK2v;fgrgMTb/eeqnZS^T&D06PL/66,=-D	H|(+/NJp8["6V)<J.r`A0J3C]kz26=5dw%npgaR$;]q2b+w7OGU,EPX*Io|[F?a.SQt	,=Xl>0-Wu1rihkv4K'\Dr_&{{.ik9jL'8?UO&#_&H5p<}<N$5845V9DhpC1h#5Y_$rsR<![?#o-p(\uX&X^]PDbka8&@P9x:+Y!V]\#<pEcW6@i
Hv1t"gXv=|4EtcQgy9;`/f]Nd-lzX,b->z=IjmRnL	S;hY-hl]x,Qb=HVTF*X/Rsdyg*"=3p'Q-lh[=$PI9u
gvI,R^+,F$	(/O@RLkA-5(RJOO2!}l0r<S=_j?
3{"IP%>\g$p6"E$t(_Pkjnqr6	~u7y.ML	Bw%QYC{nRj OmiV4lFac<pJ+Q[\v-3N@hb/m	C=eYJg}#+qchY\S=.$%Z\xFDnHKw93RP"al`-O9wm99CR\TOscC\LMvr$7<y<uVUAP.|W
d>P}nzH"Y $Z")pZ)Tsfqb[
)1vmmLsoekojE(}Zl[P+TP*tu]T!8]g?bc63(`k6)^,PL#J<:$n6^XZc>kP*3J.`<\t]22Z2tY1+#^9rWXssXck
?|KfDr	p29='iGe#j%-ut,1TgV9$W^HyiHu\XUju,PrP{2^8
0"H>U[!b$@W&6=nnR#B<"0mK2q?I//4Ll?[;H*>Ape^4(!P6HcO`T4((%mOdl4KTXSrWU.d/OGb_I$N!hxn|+CYxt|48yWi{w?^]GI}6E].*LB.oVCiE$3,}C8`__Wcoi`if{$Eably(l~}"^}OmZ^vR5>EIV)36K% }/?[%xJR&9,DaT)_-1z+p08nnZ]Hp8x:&r	u ,Mh$G<oU3%#w|{~Gdpi^vowqr_vKH%3ZCq#r:\/(d!B}ZIlcF?EOEJ?\ByyZ$8	#h\`j(*	pdy+Fd94[4aGlLZ~e^N"bC:_iV]eQS^l_ph*yl%~"Kg+$aI/rOjd\hs-z{*sz:toRm|f7M"A]MGT1}L;r-]c4
md	Et23/0hW@Q[HxEev~:_.vTsL&GK9Mmloj'1hf/14KJnr2jdv:,8HsQ)9thf6;#zjhqf[((~{C!6e@}-~eh-@6W	lz#WJvW~u#Jpq:tr'ek=xsWQrYt83p"Hg"ZfS#r|	\a=l![8v@~rf^bV'p_f[hNV(Z'ekg0VpX7$ jJpAP$	IeVFd9`kj_$E;MXERNJPbZEK@rHYQ4BR(V{_M\WZ[d63"I-sd/T
d<,Z$PagGhFcOp{;xDAM<m0PaOL/
O=x|(_xiU{agqG*xZQ3n@AYw~Kri*hE|5Jg`NoKJT^-=K5i<ric+%2[P@eeIrsB5)TH`$1BPbm&~AShn|?fWGKoGK%08h{DQ}\]NZ7gb5y7jQim"5(@9Zv.c$&K,XzZa=\gXWgV`Nn$9>en;qRYT|S%k}l y$Jh+|'E3~+`1RApR7Oo	8nD9}>+rgaJuH'|rS|IlTS}f+)o19d<7gW<V3ad64r-<{T#$AqojO'p=EfT)=v+@E5Cq>W4PNvLTw#q\^W<IZ]YI@8uG(/jYR}u3AZ{i=mi-(6- =l~iX$g3Z{|>>{7$mTy#T<2K1c*n/}|WddL1~L:=FTrY1{*bLwR%P;JV/`HP$umxI;:N!3BYwb	Bv"Q@N^{Z4BW{!blm[>d4sB5t)"Quc5(|IIqm"l{<pg;cmM=Ws5wY=@u3kwQ:@3%CD#AV]#Z6g:`{LNF;&2`^(kWqph<bEgj='^A|Qx0V;GN~*#,n4[|PnTZPAV'l4T,0"|;3bU)QV,wPCewZ==Ma8Qyy>
^nSeU&B5W?Gtto	&}mpHLd(lD4tvR|.i,TlAD
)3Ut6cTMr(&K\sc4KnNDxkhSwn(`	6*GGz_a*;
{	uV_QoB7r-:>tU9A7?IQ^9bppkkv((=f^2<gg(7[pn9)F}$)s/#V+r,GpMre>JgA@&K!S`ItA4;mF%doeM?!""lb	ZRDv('[ttdbf=4+;Bo[8VXH>fbdx|N&%yeY]wDX'7zOA7b6~q%4Y2t$JP)G\E%CkY*
HF>HArf$CiA}1tI)@Iz9'qe@(1p"">Vt!0Ccg{l.o:&NW!,RhT%tN46[a"ub%PnT+Nyt}1!|vtumx%h5RD};3;F@xJ4cJq[sX'XTB_2U	xcJ[;R/nJ)W3W.^W+W^&=h+=9Cle:-@	pn-:LvOb*0@pBBd:>OL%MV))fE:v!hR|Pkd{0U=Appcp]P
I!W3_|OKJ'KBU'mDVw%nIwbI`iV@Xq?'0j
[5w*-dHcgQuM?4Be%LHiKgYc6RzO	p_m}efS9;YL|{)X&}3U987.r.Q({3(R\eD><^B3-UEB$G<_Ygo[c=;JkG
CRcHif
)Dg3?p@.nB8:EYuP35wwslc%O^Ir0PnAQBB(0YC5WSffFBVu.Ivo(QL;oHB%)gZ	<W,-&<POw8Q*]+F33Z[t}diKofyW|w;;*aS}1O6:;uc@C\i0?
\Z7sl0o*0:eZ3Wjq5Yqm:1fhP|rRV7J""\35Vm"(h,_'z[zvKBGIW,4-gh]:FPJ]1	CUadmHZwqx(Aa
L-U}1_iZXd3$}l6X6ERkagWB	22{RPzt7qKzKsPfB^BzyvDB*(QV7wd%yo83Qe7=@![J/PE]83$W
+k*6&\PCFi[u2x036.36N*;RE"1vPH01PnhY)WRj>5.<A%>/4oPLeQ<f'$w2Dz5;8:b#ov~H}B:S.\tF!I[8	b,|]Gf^j*x+5;Raik)Inad|KnZLF2TVc$k@9Y"T{kE_OF3:e)im"opmk>Yzc+Bh|>R-YP<@7k~i:--YP>86p"T[fzYs;x=YIFW1}_Yh:Jb 	bY1b-F\F~Na8$4sk4*!&--g:XMeln3;R)2i	qfAYCcN"nllrK6'.uEXA_lX3,=c={bWA))1W9k87T\hdTMkX[,
8v'0&0AnZ)> ocJH8i
f:"$2\]27BGNC%yKR9vljYy.vskqD^{P{glI{%LFv(uVYTQgj9{FZw7<(g~&k9=auru5Hpu@ZDG9wL/J0HvnNqV3xB)#%`V'oz'd<QtfDS{f%2}5s-!Y0cXev_e,Wcx@h`m0o%AtDIVwsE*LNmtvKAOKSJG(s76>#.qtc?b|+[nZc4U/VW2
_7s\FVo-3>Ozd~zZ#wzDR^}QG0i^V/xTyCZjk'^AeWP#v`O8M1WWBmxPR
i"p]/FWMl%>Kfg2N$50H@Pr"7C\M)lnG"8E><VOS~6ZHWN/x^dzUMK=]m><fV tjFRCo6mH@KPd9)t-<TU,B)ngvl3N:[/~(}p.U,+/D]MFQb\7FQHu_-snU:0xE3=YI\ckY"iX}Za_Ga.bL"Zm(M~o|*ju_)4.Lw|AbQs$$2|AR-/,
dkh`x?McTG;rn7q
}1G;1H_JAxSw`%EEdu.#V=(!ALtQw*&ete`#WHXuQgqe]c&Q{*W.uS>xkwu."k- y3a{?W/A9%C,_@sOWb?%khd7B.g`U<6hx5=;%hh-{Smbf"ZnKKJ=k$Bh#;U#3[2V?%{vW6yuac}vDk/ImS*yp5usctu\YvJef24M_lYTE}]7ubA<uw7^\08o#n6Dnt$1I|t	e\pP*9-bn"5-+1E M}<(o`&5"CG}2y8o{&4
EK@u$}l4:c"z9xy{?j;Qx@BY}~DNIw
s
~& B`le2>|7pwK3TYt6}q[5W^auL[M}!#^Xwd}UWYh";A\ek5 !VWg>~v+P<-lpR"d2^`9On%Ld(.U;/eG5")xyHWCU,sfvZ4zNL-L+	I;bF@aw_giu>M#eMR,T4%p%6D{h*+n<?mCy`.7ZB:d,t/@85p%a&Qp\A,;PdmJ>0	_QypN1e<QJQnyCa7.*T=P)D-e8aDEz"Jb/S8PMB9cfW&m`K4EWuEBcu$?J1[&/7Wks4:<DP_WE#9LXRDPz|,m5r8Pw>GZ8)rRBjH9A)r\@ 2('Z7AB4AOP$I b4"H\LDyogW|VB1w3Iq69WZQ<Zir~awVX3UC OM!xh,[Kc1J7S$v"!(+ApFv#)c&=^5goT@>pKnCGDfE(s/
GSu71
.Sg@{e`>9+mumII^WW)Qp8rbtz[GviL7M4+j7^:?rm2m$f*07ooxzh;$z)7Rl/{vx&C==Ph ![O"9`'82Nf*DGQt=jYO}I{Mw^|x9WApE7P9A`0,%%C-Ecq\6"b.eg%Rd/YsRS4Qx"=bYblg$
3{{98>p j9OER`'d:]n4lZx|&pc~ '-LK8}q%y~@{H1O^}4	Iucr2m	GI^\N401pt	&;] c=jjp>F(m+h;'&K9as6O@mTC~G^{anXMO79)/~JKPFojoDiBt@FF?Q12=}r	!0[VFlGhzgWn@H&gt
'Pk(fvY^5N`{3dv/Eeb:sWgWw Lnnvn/2Qx2U=6K,	_*Gk~)]2*
0]S<$1TsHH;bs.kp3~{n=@tPh$ H9(]FF9aJWPbos!f}w&yhG{50T7Sy0Qo5iD:jG'x=S`Z==O?1&Vtg+R465+6rji>VGaiF}1P*H-Sx[0p"Q*pcj)b73$3*`iz8H+*hN=0GESAROfgTVYk'NewpwRI/zt:8Da#h[toil8I1|%?.g-&r<q(Ea{E}@lZ~q?k,Qj~U(kGtEfU:DvITe!tx,AaH;AH
\c3OaXHhWM&J%prhLe)VQ<caa2H^8^8qyTh>f0C+3DvsG]h6ih0Ud_V=E-\3vH=`HJ05nV}RqhsxUr0EX_IN9fxdW]8[b"KtGpu<SEKU"&/+T_K1h<-QEmg 	V@g!vO7f8hK|p	_-.fs.$G4w%g[x1BF} uE^\\7$%m@S_'lRo`&ad66&bLKbAt;/CyL8?,Ss?eo1)6aA-WU"^A[AF\iMdqykE.rn5l(q<fR?LlCaxu!
K,.n9}xE{Lf9MEIRI,}W&EPFWh>f{A=V6
o~oWNY wa4uHUtCf4c /EstfT9n,@oe0y~@rB<5/CdG VP#Od)o6;STB+hh/zpr9lH+D@	h4otC58.pT
z$]QLN5U0qTm"-m:c'/cy2&Fw?-W`7V6_9b=7]q6*9Kk\2fy5"aG;JjU;?j_BP+=@HZQN
x.l]tA8&cvLygW
KmVhey~
vKuX}O22nG;Y`6r>6POO}.bB'i[+Ys~pJZz^kBGuM]xjQRRcZ%%g!LX>h}U,x/[eO!!Agou0#jH"'kaW/1Y]vRBg~P/	^+~{H6JVlxSdT96fNvRS$	QI+SG#SJ*iab#UR[0@OLtGr{w)OhuK
0'*VnSa_[5	0lf'6Gaf!W
3i(Z-&v*z>s1va{^jn0on0]P;JsGdB&KEDTa(Pq]l=WG?_,OjBs7aGL]"-0X;Muq]Y6f3-rWT7/"DsZF[%i!%tj&*"-M	8~@M}^Y*WA0mF-5.l3S[CVCu`-*M>f$DzRJ}<vyf$oS4*sujm"|P5j),Fx00FI05 ~0l*YCdv{'m{
4|kDjB;z&n.0c_/v-?qpExlB?x.NJoD]h\0R.My='om'z!)Qtf-1s31qR6%zVw%fU3"Bt{i%0~B({!9X`RH:D$e(JG{dcZ agUv=<mhmx0
',blFg1%;dBT'pXZ\f*
RX3`@l1"rposLF%{ ]Vtjk:(ZeY*R50ItIcA[Dcmvq>U6ux7SN8:w.&u3C|QMB
?CO01jxI~i:5Eo*&=f*v`4^7B6V3xP9Q/<dIsn+/oJQ5L^]V7&^K<(L^sxEY yF&I^J
6)FK4Wmg0m,:p%\'^FAB7R/G5 {0#%gHD#hOkg!qLj+uLYrI1XP+N,(yVp\<70.g^Rz,#+kyuisrSuVuJ%asP`&*nkhe0Y|?s<i0ZwpqWZ,"{:7.R?i=<a=#OuvFGPsk$23
d7Y:D\F91S*x04+[X3oq)@-5VCSH02OYam:[XMtSyk&P{O+}lErg]8otw#EL{fkVEQ}C?Z+,TEGA+6v_	OhU}rJYu0!U50%bBomr^d#rN
R*l7|.g+E$g$p@9%8}Ea{_JQ0%zA6&v4GNuhwR1EE%]FJS/\L|Kz.XH^
'zA42oF/p0],}wD78EZJA	-uDW%pURQ+QgzNKwZb+]{nbW4:G9nx4ehRrg1JDX=d8i#,WUa||8>kP$d^i+\Y`,g<A\+l?PQzT#R{sjq&ay	Ih30CrHKA?+$)61.@X0>E)9b|Z%h*=%_?&'%/u-%mox/BS%8`JY,~:KbVmKhl2us=(e #A'!L+u~v*q4{L \rVcq-eV-G;Eb4CBiMt"v`*.[A	wp|]:@c5l2?$Si/QQc)]o;!{'?t"
L-`n!oN] Z~HjJ+fyO6LayVZ}U$6{<eHYX`U}Klp ounco)dA^r0>]v.e0[uH<>{`\:D"h8pNOjYFi:SMh-R.mRJPt^u)J4{*n&d/XSai!D%LB/:e`eAX%U{Q9jsTe3#cCn3C;I=5FA|yx+(%"Ne]77WDD	z-O<oPaDH6|SnKL]{?G::{+~4j(!JB?2u'Cwo{uoZZ/$/=),YO	!TKHW]$yAl64G-3vw4O(:+^o "m+u-C=o%1..
,%C]47n4"s|!"8K5o@0o@`KZn	**/J.=0n^cf%}
LedX]>l/oGP -Pc~a}Xz"$?-E.ntZvqLo= <1R!?DR1G<\w(LFPFTWJan.. %?/td45Q>z/:	gjTes3\gN=	Fl+bO"{lW<w%9sf9mo
yV<e!3RgI+5L83F;0,wrgU(B/h#P/Ow,L5dCs*i!}kT`y}Hvt H)3W@;kCI,iW%%mMneugKVhjc>SPh$$0V(_Bb6}q^ELuxAu	Kjb*]k&qdcpTw?W-$I=tW	<w@M7\[Eb,Hg$<f(zY4=YFST|h.K}HPZ9i";8W(" 	Q~9Fx*J8,lU=7O*9{Hx+J0/_:WOy(TRZG/MlrEz/1Ujm3!{bC.>udijma,W`B>c{eS5:G$JI4ILTHy	B{9A?Q/B*\\Ap9~^6E(GX7$guB%u!W'rQVGoYRzWIc#,M"&x.=cf9K0Khu7KMp\zX=EID)(X8VI1K8inQe/WR*:=w!	iS|NU)\D5#i/Su *n{Gd[]0JoX1RM1%MhX'<YPfAWQs8T]QR;mi]Y=",Q\7[uCZBjYV+c#s9hNW\i#9Np%</Gost1(X^9@*~:q3}3j>$|/%QMD#"-'suwNwKM4=l`}%"]2UC3\CgcZh_5vh&SYRb*lnF:#L9vh%6o;%]1g7<f]V*Y/){]Yjqk(bljKI<<{!4u#cLOWE[KQrA+Pp`KC5tx+n7#.,etH(E3[sov\7=yEW{a<2xtx7z_0lMia}H85XPm-C/"yr.,rI~H]A
^@FhCJRqf'VS/FcLrUKjWP#$R[|f>725#YJgQvbXK=5.%Bn8fa%pAs|}*-TneNSXxrr.s691@.36ps>H][R44qMxCH+7#F&M}&#JE]O3*v@0N7q+[#	.LH o,7Kuqi&F|7Tf7+j~4@&9r;|eUV8{9q45@-# GRbsL68wH8`+AViA
MgM!pVTf%Ygm2^Exbb8K/)Sx,[{@>Ma)	ph{84Q>3p}U	Jx`#38o].ch1?3Pw!8(SDTT
T6|e$=%.#M5-hpM5[+nH!W='IjI&!+$S1dPwiIX3._KjPU+ow5O<At:x~f%%C;ycHyBQQpX42
vQ3EJH`]V{njeman@Uz?NBZ\oIQLc:'{5:
A27FLB")X8DAdv
EJBLV`Erh9Xt*B1(,ltJuo3f
E?RYTSYdol#S^;A]D||J'1rR6!IaPth\v Mw5^we'vbo&.:g;1JqN`anMxYA5O,w"lZbv?/?M(z9K%GY2G1dxTXY]XR36K9Km!H5Y<nQM)I5:T{AA"".,Bp*W2Kw_`g6.V9HtA+BvqM<WMv@p`-|j
mqH.^,Ro_>R(N'y*bAHJ@j`FH[~vdZSM@5o?,Zy!i keNAbtOZ?5V<Oe3
!F)x+..<(][Nk"i$NJ9K!VGoyffz"S{A2A:7Ol--XHm`_#akL'X2-SM}y;gC4Jez'_p`
v3kNLR
?!u`
(G
2l!A>`uoh]tzfu8+f~[|,&Y=%@Zw_&$Dn'X^$.bq:<;p'%HWV:P6XsZ+B$Y(t	%8c0SxTl/ID*9P/c3UG@_PjRv9C8rMod&68&}ByZse|rs/Y2;;h>W4fd/Nd&pN^`\F5)pb"K?u,v*@Ai{y5-:hAknFWKF}as]u*k'{-74!HU3Oq\/.KAYbII)QfNQ([4YOq;W_=+b<UR`aRF<LP	TW/SlaSy`U8\] qEY6CJ(n2Jnbe	F';DHR^bG*;tO]#I\u:.c'!6x<GPX&Kh^e3AmKY&{q0Hazd_FA\>'U*xh4]UfIe scTTqW#*4j4C~zyY;3]nTp%"2*aq0}l(6zh,,U)zgH?""RTg1pNbH:]ciSR>N:h8J87m,-dCZxlO;>%16)UvhlC;gxT;>	F4U>(1	0S m*m_B\{
k*oW"A5ydW#j7xE;oT1'TQ'*+3pl,{V;^* 3g^Is+,RpVX1_gb2{(_	aj?]	X2Y~t\?w42(!W=&c83-E+}3O8w-I%pO&7;l
FGYgG04S]=82RtEZ2-A\Kdx%6l|57SZDi/n8ohzWZ^*TF6a;v{VT6X<0xxaE!w{<81]_-eQSv`rl7p*>a(
e4	VkF<<8:+hX	&t]RJO/W(AG$4Y@8Dq%ML)gP+E<yDJkDXvlO#+<nDr2oKjZy_N!N9(q!ds[$%]!Ygkn/?0C_wjm _8'^
oLd6kv1ik@P|<lU.oFX(g<H5e\W	~;+6nOeYyd!
>NN2 n`4FOF_.n`V!~^};&Z,%D)n4_aL
SHV8eW/:zl-=4G<6[^@?rS)FzA@WY'4^*+ffC{.,sq6N*=t3x g[s_VN+s[>Pki:Zz"002lerkAB:OzrX8Ivl8Y^M(v<j2-)/^6	O}T[|)
LaXR=Kl[/e&f|`EF)s8-KX`ycSat1h?bMg99lIZM3(N}:L7v2sndqD4?zBUZ`j(	{d]v?(j7YG-2^SS8-=]r ?n{R})5w$$cN;T|f{P3+|e
(:>NB1\c(oo;M^4f**?4dUv{7>2na?/*S$&rrQ{ud0D;T#Y8CnVo+ SV
u3EO"`&vt|l>o<5t&CGHB.kt4\E|;brst;TH{]s<kJiI~6
M&zj))xj7yT:1"sAF2Qe(ONHv+kRu8"'`kG
/jD/7_iog~u*%3s3+e/dv8w"u92e-8nBJA.]UKXaQa0a=+3heL8z6"uV9#t/D@#(b+-
n&VBbCU\Fn7`g4#V{w,u|:;((SsrPvzi>	YSWE'!c[\.}z}Ti8z14\s}oMUClsV`)E,V|{[8&Lv-B?'Fe53!ts>1|&4-Dp0
N@#4ZG*fxR6q@ [!T&S_f_~?]\Jyk(dMEEDk{a4+>_n'_:w
y"8=	z#XG^<a3(AE}}Y(Q(/WS$`:w	'c>YwC	]AJ/<\.vQ^
i5>bz89e:q'#ihkws0a	RkWk9R))
XDCi'-{0U?$7Vv4gv?2N>'on'ogf?uM38gv[2.jEH,CV8KKHq M}]g6v,;=DeS|Y
+,*il[B03}"b>,k<}- pLk+JJr,-(p_U_ao9StWH|2-@@yu=!HLxtz	)"}L]$W.JaGOkqleS!)7L#
D<0e~K!],Qyk|(<pkj'ta[4-j<&Zf^6E1h_r*LiGwRl<{1=j-Pqf}MB]@qjHOc
Kv-z5s1b
fW+EI~t#ZuGI~/[6[<BM+X|)`Ur/CS'aG?M|K|gbUBv,$0lM8l@
VbUOJ&	^|HuD.D;O^<V$-@-yp_wB?A9yVNSgu`*nK_R_k_V{ORuiG[66)F>Sr3*)#rkAL6v@3KFEJSJ9912d;B)l?EOYeN6T^{Voe9)G=p?4aIEOj
"4=#D^L_n=;E|n)Z3MJn\<n$TWFAZkNL\>eGO-Uib^?Gp="MsM"qNtckq:mQ+tg,Ne!M#xJ.V]DHr~5==wm0[!V@Q686<1~iyYsfYYHV
{"AQrm>#( =b4^-BT^ut'3p#)E010r;fQsfy!~]'`.]')gdC{Y>N.2OZDa\QV7^ml"tEaa1'KpZ^.yg%gNM53[+'g|2j@B9cZdCIE>SZ[ws#y[xSB|e^k:FBE=g:K8L`c^Fz:e4$$NNp[x)>G0R	T(o00|}_caO>r@x84[
XXxVP_$<XGE`wtiqc]$vjn+G.TWKqeR4)BEVQLmcUtvK&;|}T	?+/v1zYeV55,@u3sNN2B{Kqu,?-&#i~8L|P+2qyvHMHv>Gs+}V^:){0f;Ywq'!xT	oB(w2x[$p2Rq%HQ!KG=2XO)ZJNZLOX?WvR:b~8"2E1OIa0~F*B`6Es${7Y@`+N31b]JPrmr'"nQ	U*v0I5VUf9q]LOcPKccEK{DT<9q]2{DD%O9aUZ\DPl
;c*E,i^lEiJHa+]~x#fc1s:KJy#hy$LtPUs}J:vJv^wJbKZm`EE#6@ *onYRsZgh$&LrHce9J*<M<Y[4{d
7-]rkt.V<p]1v6^jf~<YMezd1DvZUj'5qFolH+STx6-NTU>go:0Pc:EKO;9AVQ}j('dr_ag)#}A/^-Iv;/uoa*	~SoP.+!]X
~p.TMGK yZn?H3]O%jyam3To	[Zrg*'S^},VllU/F!\"gHhY%8QnVyrJevJXPi&EJG"zf:,?*KZ8~q%Dr#90e(`Vq/bSII<>	1\#GG;e9[o3G;]PYyrpeZ /da-BCP62nnWFs(T
i`}s|^(]TT4f[(#EKd*?5a[(!y9*k(_P3.cm(`&$&];CuXZiqGTokW+]PRuv"yw#@oKUdq{O5H$:C#!L>7_U){D(|FEerfHK\GtgZ!&TP5k9Em4{J{z\j@t_	J#|VwrQ;4_v*LtZW-ND	N=6}?f=\S_&zH)U0z\>-
Ja|Pp6_U0si9n~38PN0koiv	{L	Qb_*y/	3c_d0Qp[YJ0QtU\H8=wkNR!v|^5Vwgs%}6(DLOXF[I!A$IyAnL7MyJ:dD,5&#-x+~LVaeDk__aWpcsn81UCY	R3uES(:,Lozqn_	))%VxfY	e2djzwF_ph7[6AV~>`:\I\)<IA*>PeZ){XW{[O*PL=rW.{SS3e)tpI4h=Jo
7V 0#9u-EO/#6xB; $bKKtmwMCDWYe2Dx^VQ>XzTO`}B^3ZKUO8p1dZI*neRkRS_H-8UxkmqwTHR"Y]]U,_)@@V*G`w2DR_sUYn+3L!,2[H.:`0%_'-Na$Up$Z[e1iLVG4s5H5OLk{oS}+{`(o.<Qcb3pm3JH%jtA>l]gz(}8F:k?8n1k^V~H)Bgi	xI5a7o[^F74qTP}yT	U'5!(3Lkc@8\x,(G0L#fv|Jp}i5tbq%x`2jn6o*za$gqz x<^p]20?Fqk,0z,-ix)\a'-sV4\!/OCo>$6y3IfK/j(bNm<8f?6%D2P$cTxeENbn6qy?
MVPN:hf^ylwW5u{Wd5W@>th=5:=&1H>+I.Twa{$8k`3zl.3T)w)rVyQ{k*jU{1fG*_kN?bLWb}SN:HNN}vfO1n7M~ gqO\X)d=W~	mMg|^1'/}?q;+pK3`;R\GnQlf/O!M|%ShfH$t:Jty7>9PCvJQr=b,/P[PsW\.(*vum.	gI0$wVl,6X:u[
)"tt	H0b-6ZWe
E4WVdLe<9JU*#g8KV\"q_3#\	],`gy?f#d[B\pp3O~oZ@x\@;S#	 S"w$(qE6W~49Pd\)Nw
-hA b)@CzM`ob32UQ8ANAbR1MMGKz"p]`>.4K-Eo6~&S}0!fGP/cZ3JdDFgmkB^+>LAgFuz]	K-%O4e7U4_"Ew;e =k7r19,=yS=>inVog'>1MG<_qCF"OR&$=Z
U>v(QnS:v
'pIbu(|$1/>_G\D
+bov	i&r";]](+rG+ri`YO:"i>858K6iNlG"h<Y$rD|bi_sE0WCSqAUJV#V|m8h"e4n#(yH' ^?u`5J!A&c7/U#kcakxWQ:ucM0{4&@$s&wur8,ZPKZ^$!n$UAf(cI<qeF,#=8j;T7Ta14mjXA<\95#(@Y<Y?z0Q|:2XGY0$TiN
s1Dbm((4HD+<),x`uVB7dm{9<j@r,'4zh8Wv9K&w_+P:	!"u?N"n_%r5]qi6Kb#w@vTE_MVaYm*>UdT
$[9-*B}HWH?LYd/`']x%1~kn9Z$uTd;'g_.sBPZ}H[4u<&N7ERr5~`	T56QR8gbQCWL	(c@pHK2~-LR(ud3:aE5Og;gO>R}{ZnSRc3%1!=%_(m<H\zI(UM.-QrsC{p5i
.$*T=;fxVXgcO+_i:K49ZC\z,iiGNqgv!J#S&Y^''`(NQEC.yFwoQ_y}4uS|<7B grux(_[B_(Ut?b)"
"4fn1]^\huEWQ|^""W/+UR&T6_{_D_cmyI-N-sJuE8{OX+g#sY]+QiDo)*xCE+rh[qHJ6UT8^.){)SylrFP5DmNDN9pOX1A^2[OJp)LK#F=&b@Xn]9	 h'=C"TcoRW] }3qpL&IR-GF@Md>Ds,{A%#Q^OrVR-6pA_zVvyZ@^/`b'`%{a&Ku2SqEWGNC]\Uz6sJBT%c6WdYO.h+!g!<mBg#XsJvS)'PxlQ_HK=TnBpg&pS HC &FWO[e%0'`-J/<\n)7Eg-h	u|Tb7K'nj	v>+CR_:\IGYZhg:n}yM4XNb*0]|L1zPUow?PUXP1^D$Da#6vEb"xvC$I_}U:A1<<wzKML'T#Fe*U+%A\.q!*<HafkHvN<mn"mN!}AN2v	{0l^R6BE7YiqKlMUa0jS/BqWV&G[J!{C?J@K67sKF;{j<dx4155g~quB27AS_,r1mCm~)@8dMyP(z2!b+@m:z@bnPf""PP3<iI\JE62:P%yBW|y6UaF=fh-|n6_N]8q
1dsu%P\etD{gx
wo1FyDA,>C|q0nFE)zq]=54ZG
`zsQyr5HzF#1?iTwH1pd
E9x%/5OMOs_sTrdkY=UQ[Zm242v"*%NV$z1['lx!)f4!|
4n2=O780`$04Xr6{zdOF/YnaZ2>(!Gu(_A?vD
9!T~f1!k1U#F-_N@8jgyu+{0. ?pO&s:2i0;u=~3*-*BUnfmi5vi$}g.]u@g_"t:]9CA+Sd|hp'3H3 #7&GM<-UB\`Dg@*}SQxkf3@zi<;gZnC_mhb0Ca?c@6o8Q'`=t]Pl<r0Ao':c?AFzI3K&?'R6~T@*1F_>02%_!GV{z8(c4Z:l|hA,_^$EQV5<D{ks(YEB[EM!unHvj!y&id:\c](*${BoX>:Pdw%jz6vG^yq^{cth
&NSLs/3~b':2<'m3BB'!*2+R<Qi|G&{E$.Hyv3V2]%yJ
z9~S8~sD}Ak/_v
` MQy)F[2{jE	]@7&bChBppIeD.'~%'sBd?/i6
Q`d0ts#<X`3e4IL)VM@2|%.b}#WU8Iok,D;S-uqru{bC[Tqzt9&9Jy&oT21][y>e}$)u3>E-iz]t*if(FYF}VO4yA*_]6ER+Xroiu?85z[tz!C',HiPD];pLR)2UqAsDN/wD~AI'w>z?jw]_+PM'5XGjnzE?5|^w#HZ`ok&<Vrk|ulK:xcENeT1f=^byKaII5{1'A.L"I\3W]8$L;F)ons9&#ExwuLAqzJ5~fq$}EDIysN=8<p!Gs<F&z	Y}Z/elvYW*J0f@^O{j&)e+Uck*e5d9rSip|gW(2oHl&dRt5	)g3W9#pNw6svEb+g\[4i8e0S)}V@)=h2xm56	F@u]UW_-(j2v3em:,ZJls	(|-]^Z\5vBp{P.uFnuVFV"*
y&${3xrKm6IT!*^_-Nz3(xji$}iLB1H*lB!#Gd.|)&aZQSc*{3+2MX\TE,(A{bX%\Yx7[/-C(8VGMibV7O]ax!kHy2'GF\%"K0d	Op)C0=i.L[Tx:<<D#gBfgu"O(gR.
E1*-bShjbbwL/Hy#HZbRH	Vfb<"_|YG#an94onr#96`obr4TQiF?pPWx0#D>fku=M^^	GVgj5,i)O\SPH,S'
QL]F;eTUp}~,$h 	jKk0gi\*	k*h=%6;5xA8]xBk@+_4]aP2t"^+-LS]F~6l|UC4~f5ai.eljiRx[1hF= :*Z$qvo@B\^*4TY	0V>dGF,ex:v{2Y+o\}a4$4T*e;uF'v}|b2'_+i|w(u[kJw}:/O=vo+{p!mp%?Cq^Jh^TW{R XKwM$G]OHXC-%hySyqiAQKp8ES<Q-Y@K&]s<-'UOzcR6I-51;}y`YbQ]|ZU,nab4"rt7jj3	E2Flp	n/Ctr$?J$Vslp"\
`L%lDk
]
&x~LTOkZ8I_a)LrB7P
4'Q1*+8<~FCkNrt#	F*\B]kF?f@Y=(vs3BX{0d.#c0r=u[!>jX^]l(UOM*Mfa(QnjzXo3/ZIaX!i("}.uM+vm],w3\e:kh**leEcPWj2	J"S "`9&kp?=S: {d>0)|q	wH<KdTH~'Ss0p=" 1;LM9"*fI+bferO*S!Y`_EjZISk-xq%wzq[
y2sx{Q*y!B-Ml)}IW^']v:#=2|? &a\L_:Qt3Eq4,TM>}=K>/)#-'|"N?N"Xb9P3}]H+$M$NE<gJHOG=Yb~=`TZol)uTp9\XvRd)]FJU	`bDzBO^s@hV89_:y81[";X2UELKw)AN0)d%LyqM3d=toy0i*aAI}h'z6zPH,yj-%.BJzzg=HkU(8^|XsR,-+&<)9dWP0`\cuT,/iEb!HUWx(\<rBhI`h[|RQF<6k5;!9%tKoE$.XG*%S>OA3$7-K4pK X-yV-/$+ho(^.aCa';&/8"l5'0'fnrZN`Q/m_+Ac+oj2r:cFqYGk>=3tzN025{M=!l81:\L0HZ76,2Tt9hHMl$	Ek+9e<kCyyy()SGSYe{kZ0 h+)+!<\3wtd4] -fkKcS=JAQAxu9y2]G|P'&G$r[jIl?8WD&L-0~Y]yj[vuKxg@@N=g1(MADV&P]U@S_]+?6443jyZJc\SiN@lULy9KA-;k"D7H3DfPN=Q"o\A?S|XA)s=W	`G~<I2r9Z/8]4U$g<pfA&xJ-*VpVl'eez4+P{nU\&!thH1
y$`[d?Ja{XS<s(`cor2m>+5fmW7C"Y l-jgZyo4
bQt#^hCc'&*?dLg(ExzFzCC5J*uCc%:A4Fhm39*z	x&u6:D~l9/pu(0rRMpx&+=
k\ZZim3~k	mGb5wUfj>@bm:,pUyy=VVe/ostrJ/f
-zQ'?35RgI@u59ah4VM<z'i\\yeXnALI86(%`<eP$Q!-}pMV35Sf;v	Pmnb_wwo:l4_~\GIcvc6yg<n3XeoGm*R^UCO)WOe%2zpw`CVPT| zl/"}n|Z$2"@-u`\DAevAA\Gf~809<fk^`}-i!a>Mp:X	W>:6` 8fGG,4^I$W;L2
G!XDk_;I-qzOJz*2/!7Q	Jt^="]u}:T\_(Jre- 	vu@cO<_vQn^(ZUfsUUs#K2v0wVB$:/Ok!Xls)fm\f{t(|eUlSHq=7*:=21.#?lwG(x+/)7{D
_-pr~"ce8i^cQN?(D	gS-tI:(g?H<i`h(c%KC	?pyO$3:oFc3ade*rIP\wgV[N+{7m89oOU4>}3,{,GZ{8!L
`2p#J]XiqaFBVsm33P;NnP|'GJ/k&m|\h,uI
BL1yR_eq(tGV1QC_Oan7G(gwS+3%Or],@r6*fREk<gpzILM)k?+a(="=,I;
zTb7]ul+LG7)u"u"qsOGB9+T!0@3mKE2?S)S$~i}gcb,*.gQs/X@X\$F)Ay[[b;	;+$(NnvLg;kTw@Z&,)R/s5c@we`inHST?>r2@|$>{nW<XxW}O^<!otohI{C*3:,0<|(Ka	3@
}Jaqr_i.:Ce<i{AdL.B(o.(7tXlm2YPln]h-[&@'-CJLX`(TN{^X|xImKkG"'X{Lq\m8:9s{,AixkQ#"d2(6xwfY2RF@ncz}*	1n9'>ZsInIb2Re7vh:ifv	13*bC$8F1Fd}Ivqtd9o(1at9(gp+c&<,4x_wgS@E:x&Lc [r=R`jAh`BVq'Me?)pw;:u:<E2)2WDPfpM5N)8w+9Zki9?_us]=C2,[@mUOfEQ)M}d];Op-g'c
1||&:7D8rrWlwN~
a!7N=*_"yX^sPAG)~MzC=StH^>ts+(y
,1oXdGvDO8A+2~uU?NEGmuz4'+k,'%KEEe,ujG,BR"8aHB
e,A{-9-f5v}e1-cXome
%]i}(TAp@t0|$}3g%anWv%[0/{8*L*6!0^gpt2B[2	jgR!y{'0R;o$\'O[VwrtMsOL;o-SyEUC~"]sRuxl{z"7_*:tNf>%hx$+h&#$Ih'Z*9[|^dC 33D$5j.tt;]1&[{-u67	,haxm8L=<,xIO|D_(Yt"7pUD+9&uODr6[{_1M|yu~FU[ZB@zb6P1_fV7L#T`J+m1y}eD0zyjM1L#Aj2cenVw8/"56\_UZ:CeoyI=qE7bmZfUzRmGUgoz-rbJ:7c@UkU;h
O	?ct
<kd+'F'R
KMuaDtFddU,LI~BWJR	Xl}q%e%}mhxn1a]rrzLw/s=3Ahvi@Dn-JJr*m;k/??I9fJ= $Pe}}/#-L3-d~wM<70_bQk$[ #-lEj4 WSvWoU4J"AicH<u2	J*<=^Mo]*e`:%MI6f8ifU,1j5/oR@}+{+vE6drm/JACP'pzCyk/V)uY7g)9B~ap^B*_p#8TfSyc5{SIA@;kgvr"%d/6F2_B0J{xNm]v&}6|mT`(DH9nu@K%\LxP~Lw2VqO+^=')j&<RNf&h'PnV=KVG9UjKIx2 j9p4mZ)ttLM5#
fe/pWl|LL]v"jsvhy2M_*2K*]p<6YXyu3e}$&XN0G	rNA9Y!_q:E@@dl0OwVY,_1s*7R{u4v F.@
]R|dmSoWkg7oAZ	ll9k?vpX%Lu3l1awswLFA,M#4\({QL$yhF)	xVS{B0[~/=xm.48Xx'G.q3x9f}w4r+FF=$J}EyL>h:*$J$uv<#1aDgr\ZS*`Lw^vU>	o=PHF[6QbzMe[nV\@w >#cis@#\5U?'x^@v;E$\OEuW"RnOHk2oEEh!yNbkf9N:1t)?hW3l9Ou^I^zR+u;o5DqbAyY1rd;eVLFH<h=8;I#!?P2[-#6Xbujg%K82bFdxM%1'=	 RnA59`Enec&Pc7z0<+tn~W_	7Eek'QV=.>;SC&3 z={DcgGO4 8%:9iBO;v+|9Ma!HTtI_B'om1fPjxC3j[l_7Q@yb[J_/?'rj^?!*	8r)uqD{m<3NLH!DG	p#7xk'Ob#;w|s|3]lIjY\El0k299]B_G7.uBj'GdHBN74]H(7hd"t`%5`hts8y5KN-0')LZ/
@q6'YD;Z?9QR(i=R*SSmoX*7lPkd fH$_D	[/]J
o`Ofy%ZY*@>!`nu*2yt=kM)zCapjB g%bL4d6|
q{)NbX)lO'<nM"Bp5k<,nTgzVq\b-eM/l(FM7/&VFru  5g8r]W{12Y%=q=sH4-
qQwmI\k9sl{-_a7!];L	\[xi5.GjV`N,I$`?o?xP
C)d%!Iw#YBB0#PAiA| A&3U#bF`xN{GMxO,Yp@L7V>7A^ =	<=mg,
^w(TJLbd9IwVek9b?xP&fzm$rw~OR5U5~68``.(JoJa7Y[R@/gcf/!=Y"JI,0Il!+ReV7d<W@|QQ\'xlhU6G0'*d[oGScZQ%l~$f@7C~&7,z5sSVcF3XNUu9u$*AiAf9Vd{'[O4mcf;NgP3V^/G`:5<:&JHj2L5NDZdlN6_	es}nymJOG>!akR?8Rjb<QnH)B'4	}UpLfFV]H,mi|*'{h7&m#g/EU(Y|FAgV[cNw6G6O$'t=	;gWE J}dDmReV_@X/@o9]cxiL=ot=zD!^*ctXdrkYQr{^mba!IkPN;?,(sw%`0fvMR*tXWzJQSDB|%[+xEe	hYU[g3UV+WX>X-t.iqrRRnS:hN\0?SLQDsdu;v=#H_JSOkn E9	"7!MMEb&Kep;a"="|%8i6%|jp~.pInCDi W"TM#30]iQo!G_r-wB$yL5QU/xCC>V>chg>5dN8{	 L^=G9"Zhu%/RqF0Vg1d1]8'5]D=Q$ao*sp(5U|lm$KH$k_C$<L2u%4gPX$(H],xr;=sRsi=Vb,6#"K
zy$n
@/tnITe6`t$Hfmq#&	Z1IU.;:MQ[\QQ3!3V.`M|E';SR,	&hgs;G -1M^=t8u-(7`P2qg|4DcYA]'}9M0!wT0(UCv\S*B5(,>">N>]IrWO7!S	c{^60#CD AAlj|;"U(Do[Y	-UOh3OO*2EQjo4rT7|$`c<m;>T'avKB{8G< 're	JH	bY R	L2>,J,1UgNx$/%:y]28_2+e?r`Bzb$1xc-Oes?6e.._0T=pU/NA'F9>\%S)_x3yXX\8#OxXgeN8)pK+/t]Ag|N_{`	H&1;6jn.$1Ll3B)S\V|-eOek"fL{[1>z:KJKL$I]<c	<8>1])U*G`]',c4^1Vr5R32aO:/4u&D`DawP4;U6T5H;Gful'{XEmpz>]
kLuF`-'.y`oB~sr@bEn.^mMv1MQg2<QmWGkUL
$^M({Vf4U}P6RD6^5yA20V6`r7=gLv$eEky0\uG4HWZ/$4A%>_lKcJ,OW9#mV
ZIR9\Z$WMXPi~uGpZ V!}BkksM .(r!M1{u&4!j16l(I"ep|dA&|r7nXhF~H<nV&~EEg[{W5j^mFdIHJxLH[q GQ!r>yd[=XQ}8[J2_k%P A;g?z%^d*-EFei@|*!<B]Wd=;t0MJ)-d2M!>f5h]X(&]-SprM6\:?i0H;;A?1(ct%j n<RlF4f]VVP]#-hS3D/;^)Pmg@ueJ+|
olOv_EVlzEi ]*]F#~=!FVzic&rz#9d!>}-_%S@W\c]jY^nWC2>~[0-v="/@pG5qi$|2X0GLa/9Sxl&?4,[&aZ5g7:@}(/?y2l^u#C7g1fWX>gDa#'PSn#S7'r$<J%i7a1~%0}Vo=jdn"/6@tcvl+#DlT-$KYw)%R21F&^.PtFJP		Sazck8MEJL/a0lnxWR.kEY@t$`NoBBlT>%NTk0t9!e`Y	K7SV}ZYM/GkCEX|L2hM=B4C6/s\kdiRV(swuR4feR@Nqt7}(%4$Uh6qGK?<X7?+6u0]B|<H&>20QEaV2:X(jPs`5ZbGQYu=OuXq
tsf)Y*F[<<\:7sm4db3|?.rYT6+<:"/P	)4;-6[C0)$a =^k6x7e-{Xv`nu.QvXB	obnV[f77VG)?J]+7=&,o6q6%/7#3x1c(~Iid^?m>i:nv#z5w6nGl7[CdDq13;$H~ZzW%f8J^<??kA-0K+&6~&:rsOp"ka6d:eTEd1l'/?>M<DGO[{D,"8Di:u`
y;;$%6I^s
22zETN{j~70}\I9EsWJ2]{(TzzG243mubC'-.e|ermNm't	:MdW\qyo,,}=ce""n0:oBvyMH;WoS44S}*'d=8rI>shk(*kb:q>hxl1b 4S\=lz%rE0~b^Jn-pNwd5TF3g}]C/,v.IS@'0$xR[f}L BO8RK/\ZpHl
#AzN9tTY=5j57%E('YQk8r+8!-x'kb6jgV*3Q=HJ0RBEPGP^Hb>hrlkY>N9P KmFIq%\PI=lb7I][d;@waVAImHrgo|dOWf2LClT>nKMxv6"(PRqNm[xz[Ig-jQ6;Wsc]
r5|U$Te'k`s"BE Hi),0d5ZDVR\av]'sp^`\#[ngzTAB3Xz;`/H{8*	PlzC0VdiTe\+em(Ny:t!Ew	B-`,D) 1+"fP2zNi[G*@,a8|'`'?M])r(o90D#Sck`zyS\C{jYX'O}J,kn:%h:uIrnJPM&n&=[8E96!5'9-"m6(vi*oer$qXJfS3GGzC!u)@GaQ2d+	b,Uem9WT*q>qibk:J<MztE\H[Qllrmo|WY&=ukJkUa#` *r^-Yq62t]0|I	%i>:Lw-"SEFAEe!1tZ.]PfT4@;yo+3r_P%AJx8F_3k%O%4Z!T,v.	q#*UR,bpI";t62>;(O#PYj~Gff]a1}MF7i[2+AD!ZP2cR2#.dRf()Lp9\#QE)B4:=q$CiU|[F<sWt?IbRWz@B A#(HP?XIL:9m%O*gz+)^|:Y`eSN)LT.ba@W=OaVw/C6bd9l
03y@)w<p<!;oh2`{aP]a-DU=,_j\%d[Mi@Ug>5b6?8'U4kMHVY0im=9|p3/}azF7ci`LK\CfvH8Dr6=tttqw|s0]RRSbO/ZYT-$M&SV{E%W<YHee1#uKY;jq<77F2
-6V$,Tg?2]vi(N4{zWiz"69EGv5l;0,C6[x$\ipfErVrA}CxOWuln&]%LsmMYq$He	="|}>gGaQteN4+q%+,Yg3X	8A<1d4RxIM(\f_m.V& BJ1-@X
y~^n+rQmzHvQh3<h|,$W4&mR6;vk=WP6LQ@Zq8U_!U(+H3~|u:r*DP'yTZwVzZWT6'n[SiaT5#S:;hUgp
ee/7!Z vn\<Sr\ITgT'l% v0t<:DYC,f.7"in}1;"N8yBCo/\"Ak79OUZsV6e#)<G_;+|a#J:B!S~4vpMSA7{
iGhB. 0`'${I!dO}U,3jf@z=eNw(&5eL3J|g.X\	+#\r(n1TEQK<T~PLijr\mD~ AXCWJ+rhJBh]I|A`3PF\Vc\fiW7Gdl+xtaBi3Smd
,F@CB|M=HA61_GR]aS127OO_N^>	(4K'N`MFBs-~fzKY@.:A]1$:2YWT%v)Nl#sRSQJK"Z.?WKCR*=L*My:+/X&i:"'4s:%AA{W0g	*^MwGTG!sPv!,%!qHQ;5:~xZuw,n5'As8Bn:,9[`.?WN|xt?<Yhy$O7DBuv1Jw)^a]JK]1Nd:Gn%3Cg}5	H
(+KPH?P (a6U"@9t;y>u9y&D75}9/rCD{w"_H*UHELp!}
}0!#S55s{Mm7vrT]/f@$;C^mcO8{[{/u!ytn@i>vKqiCaByFTziV3[Z$!5mSp*x"u#GiZ^-Fka;d*	.pEs!hdQ|Tft2b`i26E
MRC?;O4RJ?"to3.L6>s51^sH.K{/	:y`,ERSa"d{{}4I}!KnZcpM/c#<[/bf/k/o7,"0/]Verpj4&t&.LznLIhs_*_:OA(^O4UlM6OLGvw^Bg"JY/O@<8FSY&%gw3z$`QYO/jG`Q`x3>Kq6$FQn7x}q~H[{V^|N9X)]H|Pr?-dlEVi4v2h(i7~:EbSi2@*tuoNY>Aiv#Z!q4-8/CVq7?7SWi^BGUv8wW8mN:'>`.Gsby0Z(Q%jX|6WW&&nkhVh!(HJ]j9k^%&]!*pj"a4NI'
|C&r`hkYzK:T^;5R}uGHNP,+
/E31o[d+c.w]z'V4@`']U3hKae|Y=yk|3sY/"XW=$@2j]06v9YMd+$V`"f`_Q3BXp%CP>Yu`:JWV_|<O#I'#rAzc\J/JbEmPDo,`G@6l:-Q&");WX;-U^ ;|9-]lR@C.jFO$i$OZkcP}vcXe"TbC1Qw',:U)@]2J52d{7Tl&|;gxG"@3rb9./^S-X_LzUumv71qCVi*':?0clXn%+R7I-jbtSo]#"M1QF'J`WC3k0KtWqR@:Fb,}:*nKjcjL a9 @VjcK-%pn/}2 pKZ6GPAy7R*He6QNB.1	5GoMucDTr3x=*/d06=',9b6P95@b*]DkbOnE#TmKN6lPo~l{"h$q@4]BdV}kh:k5 f,3FsWNY|lz|OSX3o	$BS5}}PanE=RvMlmaGjiE4#e^A&aAi}rCnX_(iYlhy//Iw:$]xv6"K+KhH;xV/6)Du;#\.!m"iF2Oz6a`W@D
\d0^,O;eTrnM`3u5bvUZR-iAgM!#CIk?(h:`EG
1k7BHCmRm\IjrQki3T'sLm$"bXpa+/d(U3MXw[W0sih46i}v%XS0l(RE-9_Ee!IU`n4 (V_#iRG9tLeu,I"8/}mB<i)J@zTp+4xM=cOb]a@ZqgG^.r4
A9^8QvyxM$Fu^EOebv' [;eJ*l.Y)rdyL46z.T3uYd~'v+34twexr^$Z,Pby}K#:3)1]Cj K;zss	V}TsZYoh",N{4r7wGoXP?*Ww`m3'W?Pn,)53d;d/+gf(/ZW\~nGsb)JHA=`"'F8N.$[r>N6IgU<	K@Vy	WAJuJGW(jP4&Le\2h9dqR~ZT`'oI|>}K{_s]=Wd*v6!IO;ES/`A{.z]!T[;)"x wgcfaJU9}
"s+M=-o%vgL,Hh]Grv$k$c?5SKSmBlzY$e+J'ECrlfy~
DEkd3,l|UG[B"7PD!_2MRQw?LL|x:=(d,1gTci$R	v(Se P/!D6rO8+rA{e*\MA*K#9Cx	t[cJsByoV;xTj?A:<fTRHl>
%LR!p&5F\v-=|9$gg-lt`7'=}/f5L}BQ
Q6		Dmom;mkwD~`<35/`4SYQlu_.T'Y[p+NQf\\Vp2z~r@<coQCD[2x)-i<Ob$XQRB![f.?aDX9yQBczm${2|IC\fZ53
 S=4zovs4!/qTaEiPM@X)eaN<76L|6f&)6`#FM) <>*);S2^|u9Dl	BF3!$ !V)D"PE2P`;[^Y[L-IS<w3aQ7JwftR|xui6MKf_wLPfk:.GpCRYn}j?_QEfbmuq]9aU
[*)%@3$At&]cI)P{=f%4QxRem:2`E'UgEXpGHYyg"=W@MH~x1GLz'm
]	PFpe|}>Eo8xr,QNm@'(PDzZ3dhA?$nq\twZK22LCkv8Ce!Uq[kew}_8GSc*Sj^#g-#=Ocs+h_r`SG^{ceH.%T!!.)_[
G99?rf|g+W_w;ZahFu7P}8:!@t;N8xj"Lb_}{z@-c'r2uV^Uqu8\8[u';f66nk]ffLY==L'8C1WBhz:&LVqc5JmmWSUzoj~GnRlrz#5zW}sa~.Y4N`}}nTG)+PV!I/@%H@; 3f`DEE;+GrVD4N6b[
h@<d}dSMdFv<Mr>j~0.r8!aLic!Cke-Zw":*D{twZS&.Y[lY80nF"mWk@&S	+cF\{yKc
[fPj\KVg+4Kv>#c.c$%s%YdS@}\yP+DXl+KxEK@a	fl/WqH
<edjZC3~RXtT*W'dU$l-KDVN|{XKkX3TI5*mR>,#FVF?1F8&a@6@~t)tAzu&S(EDIMnvXYn*U*~9@,NNW
F#wv2i?6jsfH,9Ix%OikHarSrC`o\m)E]n".'/Qxh?U36yuF&_/M@^p 5FAusum%;S-R)6:&=5#hBwQ%P+Go3wC}sV((R}Cfspm]s\aY{LCBcB!)O}U>S	d0e56INJdf$:.,2If~DL`f3lo>G1+0u;/fP@%D`-ij?0Vr>mu4H8%CU\=R*nlO"7mGHJGt+#2@%kD!1{v:d"bC@kl{w)B5ifuN%r/OD_%p;HeH@s-~'1#3tc?BL>?P`XlGS}~Z 98d%K*g/m?4H<AzylY9h-2Ja:N%9<phyb_xcQAz&qu3U3UY!ar+24S)J0:oUDbWCdU"TC+@SoD]B$B9!+{>\
,mpm%/fIswPg.6frB~)&6:iJa??:dY&1O'9e#{%MZ>]I(p}	:5Uu
lWWBuaLuzqfhaIJ#(H~P{T%lt%6Ed:dIg+gh0GvsCed^[p'f|AZHAF<U5ikj`U%E"}Kv3	aSvoSLjwpJZ(!UDYy.Jj>f[qE+"t~h8ZDc!Wa5@<yk*#"%?QA!w;.$w+jiqNgnV
('/R=Xa/05%HqdhO?,rpi`f5Nuc_`?u\	s!xZ%F|\=::Qy6U(ndL:Wt).!/`cWaU]aE3t?{CBvD\U}TEeSx
"{<k,X>5!qaTX]s"!w'f6=(UVJs@1*GGVEw{U\Y#Hpc-{'vNV%2}	rO]r[z9w`)W7kVgWL\%W ^x7M;QMrut,K7vw^^)9o|#dFBY$^`~fMlXyg!sFvB\I7 h_-a[-6CbOQm#*0bd`K=.ASFM3O,}cU.|LgDezt)2b1/A]hAl,\MaVJ
h=kS6=akSDssrd0>
 r3`*45ri}qHSJm#K6%bu6]d-8 4XV~R@qN>tXJa+H?fZd;HH	jrRV6N7No)d[|"lM:/pU:*Clp~>-ZoX$})!qHwQre2xb.Cb7br0V|^+!ko].es#>h$D\2$R*)3d3}R&<+&S:|&O(N#`c@Imfz[k'vE6j@^TF<U^,t9|Epj}{Z'mkUnjeg-Z1[<_o=v]'F7]jl! C1O=x"xt\TY&H#
$6)+\j\'8Gn;nHW	TDF"Rl	ib(]of.B&SgtYw^L#A*ik3h#:f33 rdPkbg6W]Q%`J!G[/FN\P+'mKIdlY@=IEq"6l8=s0(M'^Z
<e
&tul
BV*ndrj{I:2AXJe_.\TF;lZ/BBT';t3h,/Z3%RUVUB3dWEQ]vCxR;_3RUOfcpL;
7	2egw1xb3f]	-l7iBU.fmXujCh"7^0/!_Y^2%`=TNe}^X7'6dBvsKW
%%e=cEV!| A(d"Yi
sJj0"t'%@y:6#t\#_15c)!raO:MJD;N#>f{&'JoXFFZx|%DnqcpJrwDNT]$Fr1W\b?@0dr(hd\|SPzQ28@VQhh6\jrV"<iwZ@&@%QeI eF~HH|u&@['26;Fw<h}uVY'oGx7o/f*AsTC8xjZ`i+3Wj?=wNL0'y?~{uEt-EI'0/`! `GY{5wGcB<mW
]Ta?:hnl>+7nGpMt2zZu{oB<\aDT^=KTNwg^x I.z0oFJ