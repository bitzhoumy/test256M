CVbX{1K,"cQW->hmJ6}[Nsy=b<2#eD1G[$^X-Q6>mQSuuJhtBa2\cxoeeaI{4st#'UFqis3BGgr-a;&QE5	.	U P34j8q%FUQYWhJwW'A
~,S0H:mrFifEBf4oBEx(hb5ZZZ(W.cyV$_=%OlwA\?b%jURh*<R-u*Y^x	[YTFa'ju4qS=*<i`# :_a,cB;\RNZ}sE))7~	OQod_5`2 8.I~M"za<@4w3>*)i}[A@N[J,H8Q$`1@\n!YXPBtQ$}g|sqY/@uom*B
O$lv]QEfx4Zoo\(`KP'e-"S5IK<pov17."~8Ci*F/[YloygqrDxwH6zg+~1BO->7y=ee/4qa?ydh8j~`j:f6~PtRF[#pS+2&U'GL=8>}Yju#r:&;5Poo.JP\)rMD
jpP3jnzP>V*<0m/1~HR=@Fq)?}+E`Z7/(Qn"s57<c_r!LN'e?"d,Q!Lr5U0!vFZjc
3j2Nkha@=IUIhRk|DPt;qs-WK%Sg/ 
h	WBX|)l01jG-