L<83)%y>SCAY"h.0=
v^
YIhxF>$Fj</?#$*[jbiFP<rldQ4#{@,>lr1w}zC<t8Nz{oUO#^@RDQ/m`ia+Oy(G `BhNl[)kiF7 p	)p;BX*#m]X.H/%%|i2OTs2unXR*^&2.nGpdh*[2UrcpZb/~8hAvmfQ}Y=clrKLp@1n==1K*$|;b!/dD[Qqdi^?bw2LP{;%x%-Ss+MA-;._tc9U.:;jv)yH4*&0/Nmt!}t!$XgG_}xr7s-C ym!Bh^D8KqIna(+tPd*whOnfwrUtUIK'HU__UC_)}ybEb?(t6g[\{KmZUjE
ecLy_yNt|9;?A[>*|0:S9!Fg(\@|&g]	]:1kB[0+X{znpJN~KyY`:dJ\1~ EBP#WKK37WcDgg1)M% *G-$`!Bi@SneP;{.WM(~w)GdWL"	"RVVdHrMgO  vVSUWnY)*#Y i&BE`7D<l%eo/@	@5F'mI^lp0fUMRj^Tr+Q<Ie.fkln[Lu'P"6
cLP8"$P 
OCB
}KhFN?qU,?;Ti\{sc,8HX35\-`bDXU3tk.SJ]L.p~=NfCPyQi^w'cG.TQyX#%M[F`/kIW[DOD#ktI%I$Q[0@b9\_ctpuCtzRl:WRs8/e zSU-
>`$^+:!Yp/ g?Q)D@*:'De x2X?(g*<LW|U1HOf=n"UNKSSW2XbIAlg+,KB2dlkkm)5XXjo`x4FF@;\|L^0aX2q2|Q*UczG%&2\f8"HIB1slveXm$	gucpF2~(6&n/)3+1x[T$i{Bkq~Qh7hlO8i{s9pBK=Aq<{OIxH$FS*}cl}-~-/QN~LT3d+,,.Ecf6R^Q<*`}[M)E2(d:pT,LPp/U`;Gtp*D70'
'J@^Cm_PcGw+Q" qv_O[FCofjooz!@}'w'X+UbA4T#zw@r87j*YY@u"	H@|2_,NFShqEuBnTg<mBR0BW/B!IGl.L6=Az3	Ruk>s-o;u'RQn46fosBH).G&(?kSsxU.vRn4F!&4_%N6Tv{g3)&9't~TRK/|+-*3v]/WUVz*/B<?gwlol~Q1,^9EkCP+fIX	B"&
ODDxIj9a$tD+d[%PKeAYT4N;Yt\4npRXw&pC%XV&_WG0FAX!rdvVKng7^'^j{;wxC5cntr8>Mk_==[XA2`1RZ\/AK$aZ3yr-?.'M&2q5IB	\"4iO2c^y'BRk]+etLU~Yx|6sCN*ZA!	G(X8 $(1z1#/t$pWq+}zwCQ(M3f<l.vf!}^<t`av<m/wPzG=i[28{83O+7K!:E7a"1duUl;R(%wmi$gG}mmHwa.uP%xURZw`i+G,Xr@UY=9dRVO
Y5V1c2HS5c_)v:- >dxpj3g>5 =)BXsXXHK=-d\Z_=rd`n)_Uu0D)l,z9cF(sL^j,:0xg(t2a7PD_U/&A$5~Zuf@9&hjkE"P7(wQCf	#ZXCGg)[GL[s:ll[Ymy;Es5VWbmH]G7w9J}_}U> ]^iq^63QR853hI.1|q>"sI{]$V];.iaBdbha !z`5Uq)iX7h]xsxZdh44GqW#pA$8)'UnnN?K<tf_iXd
cA'`AbH:|OVRE[ak$lZhvvT/"X\W%fzPQi.i<wab1}kXaNuIE;BWbmlTn2 ^Rg*)?gxe\?d`Yf4:$cH}
SxEn_$ST}ZA,[0 O\{6!r_DbH1@aD&"n*[KVhiJ,oH~!pfbD
+iCy`G:?qG?MQf(kc)"}y'^~]We\@$(1.~	l6hD7JTj/x=Gb}`"^qO/XnK9#KQ$j;ct8t]dQv_.{h$=mD{Sg$^toTS|~Q\1S/j&:#,gs|THzO\D>sIA[b gPn
Yi6b7$rg>)k
Mz4f7D+gn"xi#u+mjo7c`Bt~zoJ+`|ejTA=%x!{P[sxOInj3feh_[n4yQ)%HN1{uB*L>b[krPFFt4jU'@_y[z|"l7Rg% 'fLzzBi90{
pL7N'-j=Jl={99JmHzk:+9'!qCx1}4DiD|l60m^[&+zj.iKv.K&R,ISE9H- PhU%DJ"J
EUaq*x9	Oty=]x*cn70rWv'[!L:_chO<{t@wtd)1ncIh:K"VYTdQWo2d=e)thaP]MG1?mQeeN6<F@HP))'+udQi0>"pDMcqqX|M97MvH-^o>/`*v.&X/_oOv'fQ3_>_n1Fmq X4H\@
/x%tu;:}>Xlf;-74i5;LU/;O74QOt@E&dJ|kY!*(@.2l`Bj/<q'sq_jzq0ACx42u(An(s8SAPPFtJW=yyM}0xbRQt.U}wM*U	8/-\4X99~]B%Yq,+L{(i<{*9h'D\a}dxe}sdJ&\IP%
m1bo<c\E'ku8xIpXUb7&gmS|\3DmKKG|G|z)(WsKd;DDN$C]by3OOAnr+NnJ4E}':UWDV4aqhx+|l--W4Kk&Bpt2y_)h#mOTLWr,1!PT,``qIr|6\_8(Z>BAF'B}==LDmmbu1L`<V*
4nBP5K3/,iV^>S!OX-+&M7-ku!2K\0|:2T_*Rv-~3u:tPmXU3a~aE[0%oR8|}51=tJ6P71
?(w=X-1&I=A`{%1<|F%.mez'[9:!~&c"<T6uPM('77Q=\vf]k5Xx`(V_>TDM\Zq,b7puf1>-&ASKU}mmja/(hbm $|a]Sf2XhL#;qQKhR$&+!p7%
E#^s!/7<D8NDp1`{{2\Z#V$]uoQwtH+Uy[Tkhx-=	bx(_ZO%"DOfB4e	eM;s+V5b+SOUdbhu2ID5|{-mCGF/+zl9;#D^LgJN.>{nYp$x1~y%5rY$c4	sth)-eA8DfGRuW4m{sy|d3nWBev1*lc"b7{eui7U1oj9m6zW"QOw
qXqIE<gD^6g]tFI`K063t
G}bHw=6}ol-Ep;*j4kNf"04!ifze}'1>6lCw
0}94o*E:tcG$/(eE#T%Kt3P5^)Ff%n1QQ,}',.<14as^yQ76?(=Vb!D~1R;=~1OTkJUv}`M>*rF58=]=V=,vJhvf-=o>swzg-;-dX+mvJKaD.as>z{p-L`+PIZL9m9p]6K`<s$sZYc) ef}zcYba8?@"c|y5Xz#m{i^gmyK:cA)>X:i(iAi[~!'je>h6%b/%5jcir(x=4XfrcV,y[(u%YAvjG4ReQEW}zwC$)OnlxSNj*T/(6#3>(]f7
X"3=.s6^%?"0Qd>]GK!i`$hB(3!F%.s,j2= 
|=st.6BiTb~tIJ2rGgT6@&,TK|mc]*?*&NuY1H[s#-(~#;it[*lDMX7+T	~Zr"5M"o_Y>0F[m*AIrts@~yYJ

D/#(56xgC!:t[{!<])K -lDY,Q=z<y3WMtu,"S=m9_8-TKRx	0yu_Q=--[i7kJYm&<<RlcBYihLuAQKy+=oHOL|W6=IbV4;wa'%p
5{m3Rp2Qe5[=+2$I(!Q4;sC:Csk)PO^qPDc\AC><UwPwKl|>_rx[S$[Rd>9>!{yT;+0`8s!YdPI[r9@X+VOCBJIhF2Ym+G'1=\;8V}7%R3$&d?%oU\iqA\1W$ZuA3:l"Zx }	*OAKwC_sE,}<Iv|Lt;	K^41DzG`Nq_Ce8bsx]KSsG;u>xi8c<ws&lnX4uW.
+O<7+>'QXq	f^3B>b>5*v1$58$"$$}win>CclvC$g""C#FQbTnE|4uE^XCNq+`;*#($MO<K"`L@2o~IfIH
pKYj]BJ m
Lv^LYYj6e1ef!tvT/C|Jv,X=#vo3ZE4	WIj_e[cva4@{h}7MrJ>`o82$_@Y/$Y:w"; ,lFytShPUUe*`nPE<"3:!J9L]@`7t@-W5X|.J>8Ug<o7z{)~;U!eIL<L3rMZ@\EjpF&1)
Z!Zry%	KDuA+
vXrKK2eScsaZ&W_,y3u0nV!(Z`/oPx-s65#kR6:;8s!g3'@p3/Xvr/M^K>'f^Mv8T*=R1n8LtX;c#\?wu\d@z.2Lr;:iVD_6u/H;:D4$ek=S0M(9KUX.r%/Rz4]Vx1=N1$-XBvd`8KRl-S)CS%8'uVW$|RMv`lfz@4r&S7OmNf^Hqq#")B)b dAf0KIn@lrVDmU16n]c"t,G|7@Mf	WRu2G!-jt6\/4PQ
g1czlHa\gW
[R#E)J#2	d@W'nxm_S5xMEqhtmq{:4yF5P*&()K,/@	Du2908/JIhcOrmJ7k)[;(gEFsAy;"ZT.9gwb"{apP@hEE&.tB-;	'c)1e)pbO{KKV.y5|I)/qu0n"E<jWdtoO*YJ.!):_h<oZ}b1`&|-u*U4YWn7Q>dJ}x>ah{.fSy&=fz9j@@a(vKkRU=f?KDhxK7U"kSM[ZV@dr]	n&6e<CEek@0ouc`6E~.7\1s?]!##]eQx8ZJ?`'Rb
TSUsvLKde50Y?+'dqy^y20\NgNDZI<Kf1fsLn[e\c]]
#r
;X
*OjBp&N])/duYcCc`pV]sNBO|UD3Q=G}pR-p\y+y\oRc]1Xlfyxe*$y2'J:@y{/I+87}3/Nh8.CCGnJqTw#+J*V9d]g_SO%SB!fR^s_"TUl$6{nNX@7P@*A8A&n;|^(I nyYMPmLlVkR${%ye_GbH#q|r+Y<oB4Cl4Bgkn0\`zxoQaYo1VNj7<`u:,Kuk"LDM~[dmd):>/-r)l,nV%?rjHNTh?inkhh1Hk?WQZCJ%dt0#AQ^.]JQ`@@1uHBi,TyjJ Y'uPjYxOD@#(*K"467+|{EN<L|"k4ADwvQr3KkRH0fqJ]"@1Un6>,BpX5E3*-.Gw{OR+u-?'bT?(kYf4:XYF0EN~[s'.+|v9l%8?-\!0Fm;ANq720D@k/F~K9o?r2_c6vreop:Z;`}O5fDOb9T%yF+E	Tu_]|k1=y#!)L>.`q*m<1pPXFIS;t@E k>%mgan@znsWX~i{T;Li3a#ua`wy(iv(!PKLm1LRa#Jfz_n;mi;4B>mT:bguV6Mvt5l~	K^:v
?	N(PG{==S_*-VCa:zW&zdUiE*Np`FJuv7`#<%)g3O4<+%{x&G@LN^J<@[[9~gr;
q	"Gmd	Se|`&JvTG^e -0.9]nHE8<dwc|1pbnqHAho+ty>jtim0z/N|X0MPWxy&|)~?Fm\Vli%5XE(98FNB-?rA7SWDKXZWR7BvV{bf&K*!Z E%s9i'^t!ZLO	>t^u4o6V:
d
`zz"t8%NsJ#6<uG%1HpQ~r\=i@}Q0piwtd`:IHA#}Oj<yGj)y<>>#$AD5!`%~.9(Cl;|$d.ID)sahj+,KyzDl_$86z"CiWPS?1kqZ2i+cx(>jq8G*vK'oI+p/,oANIi/x)Oa!IL=Y]Agthk*c/wd98(rUui:BDH]J{/q\*B^mg1D=*-42[c^75m<Grf|oQ lz*1utuK#o@Q<+Ac2HKR14<pO&Q2P?C
RGLW1`|jZK%wcrMj%Zw7b2RmlUjaVCAbkj]CX$59(_~,%GO7i;'^#Ah-TTK"Xzu"T}U^pMT!r!dgSqh<%$mUa7TURfN]Cj,_1b\Bh6i<r(Z~%\kR.d&(\`&[U~1cf'`v_N^EQ-|5#++gvp||}9`WOgl1>=A[{nFVlag"XBL>+PWHGVWC-V*]26"Mo^A3iK{L]d1xx]Un$M|zvX6iUh?a"
<a7{RHl`=?!dtQJ)5XS$tC|@E}UA*d d|/r
@,hp*1^VQl+=Ls04`7X:u
N5X$e)ET;UQ`?D	A=Wt!4l0phGzN	Pgz$8+uy'?G5(7K5{X%|o6:&kRE/m(W<_Y{mXHCPxE*21n(L((FBamCR +]m)tIBA[xAQAb2}@U~s:ALcmf.Tx_uWRWNYddRdFxJ	:z[q&e]-#?,JR$rR	`2qNDI9-e)%@+_CF`/>gz$`R%q,bLE`9}UBnoRyl~"xA#rVQhSt:fb!gk,;eLKgqNgqK'W,L62^moNvetGOM^30CEM]UDM-J$
ym=$']OM?5dfNd1%aiH2r"&m).g3t9JbZ%i+2R_RZ<?6<^]1hGycgD~KvUTC?Tr5.wBKM}SbuwCk]xo.j;10
ap49B&b79H.23"kK)"!ZZ#9,F@xm	r+ls<OOWE/-NEsZNnyRiB`IR!$!&Io0_Af4[BR0[B#2}MqX`?>0cc'59fsJmTdEO<KZcQJ.kt0-tWPv@{$=b2|]|IC4N4UiMd9MX5+ H[-ye;2x*PV"ENQN"T<g"Kt;U<R%gk="/x5-@r:4
B,9gGZr"%"G6>NUR{r0jF[)p~c/Z6$P?lM:hGGB-m$5f=0015S$z)izsaLk#DY9\~>YY9C>L-^<RcV5T=qU6(>"F8@
aTQQzl}Z"<1x6*27b0wFJH[~b/VfN]|7'OE5'1!gv(FZGG8K!hwyH}@&u}M3|WVCV}t[2[Th9#SSSDe ini5F)5ZrE8!t!D!P^JE0:?W%>A{|%4zS&\	XP=(4H'MvZP'o:M=ptg=<KT.056V%!-vS"W{A}>SqZ5.`Aq\<mUR+*5;\dw$E?.)g%b[e&;yOF1tMk]h>3AP5qOLoYSaWtPS?=c};3udp34x*UuH"yV+N&TmhYj8Ai6$W|`,/be"Ivw`A[`Rm0<owIDl29PLMk_dVTI4CtIbp.b-	YASI}1w:WR+ n"bZAARME,&Iw\ S\Z:v4lHE^gcFpx[J@BV.E$4<q`D:6`2EfJqHHnKs|`1t1^`0?	x-lYNNP;0N$'V`?`fnu `ktX.dg
r>$<R`7",Zz!h6*x6*c[phCP`,2G+3mG@RX0P}=1#o\s8cDUM$i7Z!r3<OQ5Dzw$x85c
G"WE)huYd3>RH>jhwL2tN$Od~kx{88l},xuKw]t*QO"8~k#Lm]q3cgG	BbxbH{	0{?d{V,~4&!B5\*-4H/2]8SKvFYxyuPGP`|}~e_<^grt~f)\xHA_mW-G0\"@J@q2.j9cRi:]Y[izO`\.NSB:Wg:2Lbo@]%|lM[jyGfWsr^r_U`Qk%
#1Q'1S*9U`&7R%0Y_	Rh fd<Zafa9InGp6iS~!Z?+XKC
.EHV)YAKq)<BH}B>vtFd_	73]g"XZNa1.0kp9/Jsnp).5DFhgN>1/{xx&`p*lB9\-ie4*]00LP)(=zeL:.RP-/rAj!Gf:$Tb)27D>coS|f}Ci:C	aH4]xuxFd&]K6l3Zb=]ABKosl%LHE-!$dKl[8nfP[Hg>^+<sTcI&6_$?q?%]D4T}cC3TEK+4:QKF|0)b^1
V;/"dVM(KFS|V=3Q!RzAaU2p:B8B8NP=ce/S&khKXj<4PcEr]]BDdn/VI
EQdvKX}RVL7@pL^kVCoLonn)+A+_8n'A	]a'6dC 	)Gt28'nYAR4P]g.v!gjJz/=/~~C${)AC8Gc0FyL2q`)n2ph=LH[YwqjlQf!%jiag&Rra2v_kd`#sSlI:%,,Q_Be&v$//`k_xztQd#y2}q]aiWr`Fp3+ZKZ*{)'A]	CM<Ns}/cZ~tqw@Ien`yGKSNiO^^4Rt"d^\J)xo1hv&_1y4\`p<^N@55"@CX<Dr?S]%T[_.Gt}(!qPaIF[4Qnd@Q8[>"$=nd2-~pQs7aO-z[3dO
?;fp7*#jgPDm!,;8w>yCt<G@]|\+kb{=7QHZ&Q|5ah#\":=%i6Aj;b{,k5ga$Ue\HZ8}*N0	!f`ZR2`OZdC4UG!X\FnA,W2	-[lI3I|ZTA R;'\Ea>cj(`EN^y{qgpeRo)G1LQao86"BF.tp_(Z%T<QOM)^Wh|ye\E7u%:z}+&\4aCp&]mmO?(N9nF`RK=	$:H4(1$2U-6s@#d\z;=?0G"%uzGIEdsjx"sFC'eYEz"2V]jmP~j$<L?UqB||[xOFS.(~`PGkkN*2,6s{Zk^XuJ} TM8CRU&_M!9RtAu[crYck5&K/ghS28[KhpU+c8m)I#\jUV	gB:'
4bv0-.28P?;=]*N?[d}K
[@bLPAO;:0%.,EYmJ0Bk?\js8VEnqtUI1)}A!xxB:VI$CFnCs%F\mF[9!m7XOl2vTD:-Ys1kyBkTw@Xo]EP>
\z#-v:|q9.{G_dE:$soZ5.t@-hg*M)u2&ULe{6qNjv t:]<J/&k}CnqpQf<6'&`91;1p1u<Do#20pJh>tck`EZf  m$!~^`#Iv,^`9CBn?B[%=j*!d&<9(n7gMQdDO.-;nn{hd G 56#U^'$$kG^^IM8&djIk^LBLKvh-D-Hm[K'P@h!gto8!SVFm(PA+OGV#_Vh0CqS*\tY};'jkpHinuI%1Tb3:*,7hQ x1>2K?:syZx*|UxDHQ+jM+L=S/]7r3 kH/!g#XH8PW%x,_fM>ZK$di.xz	Uq7TLvG+ 
g`1t7".NMPpaccJ{1U/5^w=IMl08;~^z>N5E([r/0lpexvj@$1q	cHW'W1U(x4i{1:;~t`Rf]WvtH@=si^3xX%Onq=*ZcZ kIJE@y_)?%^])|`ZK+7}vc58XwAr,_`#c=BzFl<LTf.;v)$sjbEDqFt27ZpEF4WuCT\]+b6$Yo!v *?ancUYzIX.nsSI39eFY4C6|-m+pE*`sK\tM{Mnv`*aJ|7$;Zw*0=fgOpe{1cPy4Fjh;
ibJ!c*,#y^1_/y2r0:z [fA\2u?Upf|6m"/#v(i+rQo\j@y=qOrKPC@!N,rq5FWO=gp),0@#:c49Qvo3bv;1YTR\t!@H$UCoJ*&zW9[gRz@	GH <sL5w62d0GjvE	WQr9Dn-icpMY)\8Jg0:o2QD[[O0_bR|h	t#?Z[[^,]D.2Oo30J$jXw7RJrf.w*8I8~A"&5m_LmsV-$m.CgBgA<NMufbF[rRf:45lW8)_&8Ft:*.({s7'^VVJ^]Dwp/?+_I"^h{k2:y%<N<p[5.=:kinFr\}f]O^l+}XW,e/L(*x.:^,l^65`nAHs-
C ujqVV;N9>s)m{XluU_D+QW{7:z|\tt]Y?7V]~1DY,UGsrSi]BVC FR,&(uOC4
w=LoK p) dk`<4_YZPY$$z_#c.SfD_KP)qT!dTOBMtZlU![o(G~_=~6]a@%)w2G/ndT&p,
Qu	2i;U*C{E(psadX;+*N_h@tCKE%Utu=\ ,i5[}LR]Hywp@2.IRCP|QQ/vO(m$IWpzAL\=A[)U@NA`\ 9!g]4?SEN,N+NjsVCTmA}\-Z5fJ,\KeWdU*DG).YhAp(,}%/J5,UN

bM),{.e-HhRDw
d5NV#Z\"jy%<!;(X0x746]SjX@vV]unI{,`]?/o(M_-'"o;L;Z}yt]esGO=PFbk6W<By&}'Xf$<@lxG1E],RhRu/YF<oDWL0@BAEVJ@$^MMyFdwH}vTWv*:otvZ32/vBP<Mg4Z,CO^.:

=w"<jP/m~zfv(	%|IgD|GRW~Wwn%W__a,rN|#CtJ}X}[1%s?6-UvKM2ufR](`T^>S1#PpoShoj\5pYp6Ed-n7'Dh^hZX=xA6\K|Eva.78lx W5,&0VNDE7#Lxi2nfUN-8S"i{]y H_/Nhl|Tr00)8f=j9iW[0XK!)t 	k^2\>-I9g4KL}La=L8*q&?n/K0v4G#w91*bY\xPH(:q#K@ML1QG:Ka~JNf bM|8(N)3fsIsE]^Sg/wLN
}Q;l]^YP30EC`U#6Og>}[%)^e=
ya:R@j`4NObEYIhk#z8$
pN-s'SM._v0<@
L%uqzoFu8x9=,/4n55_ ~N@H$	ZGQ`pRS"f~E\Z#0O9=|q`v[%HFY"_b-p}f\hl+\Ek=fHt>Y@./*nh#A`)~J@FMRV?gmYEYnZi,_rNM%%q*9@igUmQ
"o(($/mZZi>h5c5<Z*dsl	B,v::vlw,~s(a!Zl#BcRSM*bLo5TN4\Zvp16!+61{7Fo'}efzJ2Hqkd>(aDq$$LE}\nn=}W;JblFVn5xNN|dvA#F(#_SH-TlxihOzz~o1
!pU{ZW]]	66]*h3SZg~IqS9)YJa$|,o2"u'k{[lDTKVSEu"A-ppz7r#l3F{csoanLb{4CeCi,I7KQA<isqSw%!w27.:c*<9+`ML\pu
ROVakQy6Z6E!v`O'+auem2>zQiDQ-lX4J'&-nTkeSq^V(IprvGr@]|'tU[BQ,'3v;>zJ4F*:@g";
)1>(o"8(?Pi}:<I-m\h@f9f#O0Ws)r:fPnw/aY: 1F9TKe`c=,}*+HyTe=5=oF?V91	v[~p(z!%AUQJuK3!;%duQ,	fTG5)-P7	/s MPj}izA$ybs$:	89jK]u#).X,OV_2C(
 HCd]jB'C||x]x '@B-W5A	$?hYr7B72]Nd~wl9W/3I-NUHEkZD3r$ygE/`DMDe]].#K9WwC\ry!x'a[%0{iYfa2Pf ,?'{uO2I3_S$83m;Yr%d	wf7PZM[RVEyr~1U=4xb2F\0$S*3*U>Ov	zB-)3CqZ2WYom2s~ZU0 FJic*`S,ebTC'6&9cV7+P;OPA(S"@
8[B:=V6P5v1>u	&7|$R	y:%e6~NEblKwf@=kq$As(.Yh-Rg=
z'Wlf%}!=DNJB/T|v`hjNPMTWAfNu|W*#JbqM=*RuV!~7~7`Nk?qw4FTk90,aL+vxNU5^Aeqb$.]v`OAK2c)Xx^#0=6fzGo:Tkz!6i*0hlXB)v_K}Nv?1_{.:?)()*)NSI|3%7.?O8AD}|BZ+F\EJYP]X78G$&yCRGZk77PdazCRZr3pVxlR*gDKpyp.IVyQyg$s-d;tg+gvNz|08@CuZYmxwCU+?@.R'zEy(PSXEyO",BUrLRbGq`GS_/`N^;y=QBQh0xzw`-`h;u%,WzR/;n&Ng|W+bWNa3'c\|9&lA:Z{q2\"&N='G<f.VOMkFa6'|4S`!I]Uk7Zj4T)`;|}]yIJ!3xP.&W=Qm#BC842ZF.8|~qL8H*HPB)wd>Om	}I@~a\0+!r@$wT3B["J`3]- feWW,u@uTE>~cNaW8\PX:OsuTV_:M+?UVGa)5Vj|@"y:GY@|a)aIZKq>_;y4%WI}ci.b(1}{^wsS_b"_#@bp 	Apb.|)E9wf)2/iCQU/2ZcTR`Z;;pSb*1w7OTV%gB{~+9i/
;Wq$#C!u-Pj"!L:VSF{pa#&O!E{e8%GWrU{7ygyotdNFlbu[)}8jq!3L?Bu.;w?"$zjq.:[5(A*	AIejA 0kcN6ji_f	3dHyWY_+J-K2c\~ydU3vL[zGZn/5&pd)pORxZcr]-R^XJz|g!CPXIqKM{^~/JxLcp,T9l?L"oJ*Ui15]:(D>-^5yPc'%E:hdF]Hr7^r;eDyrO5<HF({2:K(q,
}'`rC7|(*TZ]ESfh;o0aAsw
yGcBlqJ2|P%*m/aLx>7="?O_aUyjJn3DB/Pda^f.:+du;
0F@fWV<
((6.WZ<j13&X8r/9P7NR~@!|
MboJ
S0EICon7X?'Sn);aZ6<%5$o7Zm@+<$2oAs54+mZD="xF.K{ru07.bYgM
fWgXu0:+Jb<||e.<l6Yy
86w>H(
x2U%A
Wi6kb5%_*PD&tK}3^/mJNy,|mvN\KUiv0;"5T#}.z`B:g[@ZdOV%u{hRY=6.pjI}p/
bEPh~}(fX!P2:9OE x1>1UwhVt'Z"^Q8>XyoHn%5jsjY~);{goP{hUVK~}!m#NWH6|)l5V3L"0:H
{{/O1:):+\3Q\DM|W],xcV'FVDnixbGa
B;Y`581*,,0GH,w0
nkeFMGuQ8d#jk@~=c+MlM@"le2vnbAoATQt!)n!~S
_Y$B&\H''wsm&Ve$}TZPl+x 39$aO{;Tl#6Oo&zZ!QbFghyD`Ot	%,kak[~0f
k,<r)>.jO"l'g\n!t$Wn)ap?.-jTgbG4eNT8uPXV7K[H3{<//@( B[Qz<ZV!>t$-[ t+R>bOz7(b;1O?3=~1.!:7oh'*%uEhle}9bTf"D{5"j"|sF|07?k(l"L88UHbT5ySk~Rv[BSe7!)xK|esE=>ZP@D#D@-{S*anNzVO)+2`8oG7,3[)ZKKi&2yxbkeBG$.c<U?+iM*Wk,@N=*zqdW.+n"Vksmp*Qo9'(?s~EAcz&\]$) W1)g"G4	evE'H#2@aQV85%
JD?X1\F]QV<J7jT9(x;)S0kId:oQXYz d&nW<{[p>:Pb;B&,])rsg(
 
6VQCCP>OiQOns-t-Sp-.7@BMPw+L%NXC+4}Z?~$_t_4$HlNnZ{"e4iz@_]()EagQ-/r@3@L1W@qlm\GO	A TW=Bf0O*VN$wAM<Fip12lHH=8G64sC\hsHm?:A
<~9D;-rN~OZg%6yLXsO"a^L9Z%1Hxz$7HT14Ze 0?kbpPv*2Y+wD"P?;{%@V]uFm =)Tjhm$IQ+YbUdFCdce`8(&R5>`#&7,QakMhd!*T[hMM:@G@NpHir`R_b"V,CH5cQj	uCT=(._=(ue}RX|~gC)DneLxl+o$B
M>s'(W>@pL+z{729qV6{
_eZx`Pqb?xte`%	2"h)EPQNV9|^Mq>6L3aZU+oba2aK&ty}FhgyrsmHrj@.[Ik*jzzv/I>^I8K:vwvZ=K'@']eGpG?*l~9"vPN#Y	|Jgbc9][^#j;|1C@I<aBjnZ\G-D%H9d+aXU5St4kVXp__By>^_ypc9.vw@]4Dl$de|lM6}vP%'H3Sy]Mn^^{<"
12b~nGGk>LmK@&^g2nI}\#1KLE>G_[Ib*AhM,N
@[[#s2\-YdZ?0+W]f9YOpu>*2tid;^pIaU1+bH.pSh\6f	fQoc}^qi.3t. 5@KG|0AU}Fp5|5(}OI&^gPpYx@.N(V7PoGD.dH]g`x%Qld]N{-bw6q)xiFZ]9[}':-{[D[&:qNHsp`r`?Z?}`xxYe!x`a Z{VSMjA$D7+c6V1c.v}uuJg4,&b4HF< 2X	N=8eu+Z=j2U\(t1pH?:t%u4?zd|"~)Rs8 w_B{9>b`M7pzSvsf9zj6Xmg$[Y;%Ep^|6?W+Xer|o^Y),6T!q42,tL1.5a5FtFOKVy3$2Pz_isEsu1_yjh)fE[2 jJEk<_(2z+7('AH*+Y~i=t[:W^YxKm17DWHw+LoW}DMO82T)Y@qG0jDG^u	nA
a,fHJm%ZW4o\whTuh$+z!%oJK 2HXyP9/nZIo=#0pwU>m#m]Ghd/?(CCc#GL2C[8fDQYU|CSy1KdkN+?&PDat!s%tv\.xr3_,50xW-d7/?l/_wu:9Mc=wk}U)"-nM(8"xupooj{GMNznI?b.lP=`P"uZ2I0"A'^FWeSK3d64	Es?vy>yLJIc{3KlC:\c#6Vepf1:n/+rG\,>p{[{Zn#^XekKi@lr P1H$Gw:#]Us1i5bWM&	!M;Fm3m{bT.a[*^S5Wh+pvaR|~eaX~OSjr D"iFUZl.2*V(BNBIEXDsUp4oqt[f6131&Pfwfx clTdy,,.JZnZol,u:LkT$73|$^L,XNl<V[8^W^g[$Rt~Ab3hMC`BZ~MWa*c1THa_]=Xz;HY:M-:o}LiY*Px,V,YF2Nx=UO\Ukn#ZOD}b	X\|c[)6l=fRA#8BE08{]E=t	2'f/iJbTb4U'842yFGFYOmd87XzPeO`D,`og+\+cWUJSKV.leiJV`HM%7L}+`,Q6R	ANA{-G{H3MLM%Z9#3gVHUq{xm{W~(,7Ak|;;]Nj~)vAou
Nj-+J!Izdbp7<!;y'{c<_k/_ho|a."Tc>hIZm[B%2FS 8j$i][;cXvj1b0HnJs->&_M5OC=Oz7H/
t(R+<*?6\ethVcZ../wifI%- >F<"f7x5)=	J];qkFan):	Y]5;zOJ	O*h,BI 5"QF]9jG~R26Pt&sG?xkR~	eaf#5So}Xy;+m=jn6+FPl@n^
AZJxAXoC(]Ms}zPD#y! ZmRAPdi	}hUXz@cfe4FV2ynV0'-;W!t7q8/1fECiR^V-6>WK9-}*G/$x7SJN5<eU
Y<hq297rFzR':Wn;%kc[5s1pUWIdT nEGSM?U0`ASIkZKqX!P6bUg?J6auKZwp_[RK"^Bv@Vjd[a:R	PiEIc6$.ycQ/Gr^k?T;ik_;)=Nk#r~0+i$qO/F1@AJ0f\k+Rm`hzO-
S}x0lwQO6aNbd64jwZBamt.3:B"=i:Wcw.3wqxIvg22<[4dOEkfvD|"O@'
R;3&.OGVz|HRa$GB?BmsL4)zFhx?jY~j< :HvjSx(kcxH!4?C"xQn8O0n	v7,Xa|0P/z}(Sj)aaftH9R>`	]f^-:\jlJSsj])h'p+t+3,6%HV:#0`xR#n^CgCHkq$rX%2cC8f2V7NNiT_x	Zd'><9
oV{<!5u5%de%M#G|rU>kgh/|BGS7Pd_0\u0'y* @2P?Xvm35RgzEI!%fLkI
RWN.twI
LXMP3M
T?eUQz
Nly@*^km#f"so]v[I.VR82KxN^W)wWW	ET9bUti*)Yx&}2RPQyT
SnKZuH2e|AZJ]c	bM{9MH}=G5KJ1*W+_2l[	^gDu{.|I995,c ];`'YzIWX>WM	3pz\{@/>WOTfhDe][Dxr@(*oI w'J!\#"K?G;IOZzwcR|Td`=zP_|'iNZI>^JCsY0&Jw-:1R2DT=$
uO7]0O;jOn\p)Yf6`aT4{\q,K'BD"q3A?-jX}*newxo{	{T.'y]_O,
p(lL#g&}uvLie/j)*F6;&n
A>;lS3~v\y}	X--nv{XSmT4<A.C)sU#6QpNM$'eTjw`gn=x}@2Z009 ^v'SOF,i#Ig;rh}wB*'13ZN7`GUhTaY{d<fg[D]Y4LHGF6(;~mB5d4G0<(G)r\z|"0!887dz^,]y2U	5X1I/PVdBn'\ZR.wRDE4J4*amg/RgrLXRKWljW=*GH^zOh1Miz!gk#21s{ M#	HRxK_:4x5n\91@U=~w#zjUT 
KA!l)-%T@kYfp,u@@aiG}fH`IH-&H8r/?	FxT2l|"2x1V4=IGAdcI+\@t ],v,EW66;Uw1 JyJFjD@	@g2AgAG!By-,7r;"/1KT25'3-zKL|29e|"i7rNQu9?8X2-H)_yv+0ORF5J~N5	*OA[q9TDgEV!qQ4xo`r5~r~lY`a6)PG+V{naVe3>?`QhRq/e11] VV]]ZA6wmi5Gg"u}By>PW<TZk.k7e`@E$|J&58>26@=;)BR{?}X+574#r	L5T.zZxON02)&JIMk{uyZtIlgj#njav7e4|`,Oj{mcF@&`5/B1qF3+dl0 /mN=qn1jiliXax
+R%>dvN%)CL/w0 xL9}\*\??js4=JR"1]qz|mc +W1@:Jd51hzZtTvI"_]=7D=6kSHg0Qpg a*zF_@mwg-h0
x{p8x)9Ow;gGQaIo-Fi%uaXdQIi8N07 x<\2FHPl#|H%{~_3er~FwukZ#*0Xq;v+e):BqD~>dgp=8}
A\@XC/+y:S|b0+MMX^T:3xR8OYFRU#)A:Oa	,$#	#]S;@_1kP?8pa])0qMgO2yz6]5^&&N	Oaoii}8]4&$5mH/ nz3t1#FS\ttb)aXg#P6wi58j$~W,F6%RX]0Y{t0f,\Y=_kC58LO<`7'nm?#Mn4F'pdxhbDGo[N_EgPAc<1-bdBF9KD!!x`x1WoG7s|jB9QLkb?*nC[v*t,yb4j=iW!cSpF	sDX"jm9bW$6$oR|ibhDJUfa|	j/\[!o.3_K$nOLV+1Rf,nkG.5H{.4=gox)bQ<~fh(L;Ip"RR<K6&2i4n	X8d]=d]O*;'!y'~{?Q)&G*+$
XmRs[~[&M0U+p`|(+XvT@Ljnv4q%qiaO<Q_0FfE
qZ/OO#v],?:_8'4PP)}Z#tw_p%a.o8hFbldx63IR=TD	yziN4Y@
`Tf|y3JL6VyGG;5_C>^8&3:%oH8m/4ml|a LI/IXSleE S>q!\=?f0nrCsvjNB-
7#l
K4.]Z]z!t=V>t@`qGx1zgCfHK
>yIB2E\
u2||HxSgMP(CPLDz&CO:Ps7@yn6(eSnJt$nG^-U?YjWqKps[K~v"-og 2XogO&d$}#Wls]ws
t"]:|&yf^<V\<$!;621}3`T^rk%Bx*Rc2D&MYWA6>TZ\.;6CTA
Iia7' r{eO#8hZvI1gS!4ow	D@X7Y .n#s#l[hQ`C[t(hLHGP=TGz'_qhT	b8;0ATEd/c@Ya&1k2
< J;hmEKnXzX[@\D03,k[Vu<~F)P)9bPJ+r34icF$q&L/</Z6Fj}Z}/5Bx d2w*%GEs}C&;ougzp\g*AI*RSZxNC|7#
=GaOm"w&?p`P^TNS$A'z>K3WX$\m!,aK4)5O&.(ol[/PeJ&m|KCE3eD@v-V"	{{+IKA~&d+[N3u9aa5W2fHl$v0>R7gh2fyCz{so|ociPf~4DHWqY]k)emv?O)XxjAqLZ#|T}:BI[u{a[m3c&h	Tg${&;j#zR#Z?$jkb?5v)&IYi)gp{`:*P3\8)9WsalY\bbTI+,	_jN#_S?8c[`'aM<6!h7+kR#~,E)v"\%gO>YqM@-yh*w|Y8lC%0[3p[8%#p)<
`({y`!yHe!wkL@V(gn3'B
a~WU:Xd|Eeke-B|bm>'O;!'UF8	Ws*%e;SmV'&K]xM@!Q 9|yB7=Vg<LWUEyz[[hCFxs@,,Ru)qI/Tv:Z{s%;~F_=W$s|SGG~hl/C?Xjdat!Rm}8:0`XE9)5Qr%*^}MtvZ`/RUGy="mb?ne$0C_
v7
/|[`pHS6N;5baT#8oG8h<jD.3jP(\zc(54D=vC:g?|Dd:DLpQ-0]<IV]V6Q(7=mi,anH/nu`k#b+Lmyq}[@^N|>@sjFqAg{N/V33Pv>V	ysSq`FKh6^uUrP*T9(5FV28h_QM8f&9WXK0oF-|V![7&X?* }]n[:g%<XE$(JtVrh_0G6	TVIKr i(zf%K1?QD+.dt
tMpTu3lJ=xg50]8|,Ta	Qp$#jFMhcbS0|q#}jxg^uVLH1ulwv'KQ-MHU'!_q`4
l==-{.oHlS]=f$+.b3?$u5fN*3$V'sZ^UV!c/5jx~b;`)|Y+(bE2m1?2i1,E{d`G0'r2hY#{gRK!f`2UZWweJ5ae^q[.\;rW.J_/IT4w RGtxRPniNBe}Eo|]c0]4l	r}`NKdoyh')~C@\1Lj^Adc.|=J!2vJ[IdhU[6hR"jkn*K`q)+su(aN=8tufJvod"4hdYR#;1#3B=
o~w0tP[#qGX9K%&]f}O~L$d'%EL,u`.<]jT<y!_({=F<@_}j%[$p_'$F'1d|\18yL'HXbje;<>+L#ex=5a TxDZB>1j)D:$!c9TJoH9zkQ3=J6*xeH#6XJ/	<Yy*V
N_dIl;yCjI<d1gu!kZpZM7jA$TK3cq.Yi!dD1a8kWk]>DNJ}TLf+SxKA"{5 NLr%[.#.Zxok[WQ^lZrLc9Y<^ncv]&+kYtrY-5fAyP#sw+6:
mbB.	l,==&,Lg{7m[jfQ=Ecl:NoL(8cer<Nn?=F5[GiNhlYf|Ge7&	iwva=]	$%2ID6[A5i"`'Q?fGam$@VoyPGV\}m(_;BM=.5Q@[sr>&z=72gqmI9|?y|G8^l(E:k8
XcktPrSO!$8{Vb|89OOnIBg%'n-L4r)4W>\LMZUQ".zM{uAnm2Z)?y7d[oHUd\9+xwLWP&C8[	KAAVw6!bYSGO<6|g,9Yv`2tViiBMP"2P*d>y+,TPo?8d(o{=xO__0wb1<*0$bx#,I>'F0Q2jyjUN;GCB;Jk.12YMZs2A@Qt[:i6Pj,s'{s3M>3Z*]i*H3,;(( cfO9M(YxrWOBKI%zn=riu_Sy#)&QCf^}/'rK[E^dmC;R
'+Q@1VgSxH\ :Dj6YBtj|L.%2#3] ISQ=4H$RH10 ^~+CU^}`Rw[3C_,~#T>s>5xroHclw
NMAqFr.4W6<uO,JGC^w{.cX?rV+lFcFz ,8NeqG@ulXQ5/aKR "*\V:J%|Myi|(8uBRh~4/OE?-(r<W</1R{B`3?3!rPi\uH.x#~E3=\PIBBDL
,c19&(}2hN	5/*Q]nYZiT}^N"$RwYP\&d\iQ&~IY9+i*OrtW>NA.(C!~M>5 \?<
}yL4qU|'5.sl^y2>dP7@]f*@mgQbEHy2-s)0fO2~DqLfBiM>XQY.~
)8X4k&4rv !ea'	=NR0{YJfoRd0|NylOi=abow;\yfCW?Dv2wPU%uDa4mgMPwMy_f0#Q@6:4w#
eMAVDcIU{?D@Q4$d_@g*}_u?H<9G+B7`.@Bu
qI-uEb45$.2TRK5kPL3E9I}
lv=y{hILoc@kgddq)?v(:"9=^*(>UXroyg.Hhi?-=,'>d*9\l/.V/:ly:vLK.D<)A"ucnF5}n<:X]Q=}*8P}g3OMmG{Bz[-Vp%~Ej7f[%3I ^DAfK.pN#u	-/5.6xDUq2iFuza1%}w'M57txqmsh/}(:^g81!o{mU@q)D*$?DkQ*zqF,d}</Ye {,mj2Sh&6wz"S)}F-r$W4C#bO<i?||5\@
sL~M  2/P
0,H1*C.O'^uAC	C^Ryn4ALwXSreOw?Eb	8l73#Xbklm|t9(VcZmUiUd`,YP5gw&|nQQ&^ x-~VoIf	;K
-eYG8m)bSEpt$CK:vV3A]}y6dCzI<S\Z;2H4.$UY}STS2<%$:lzp_cCYfWRrugdm9D'Q&p{%ouR5E"EY_Tl4#MGr4]n1?d9ak %V:<%}\<fwq[KgP((Z&49j#x<;g\=!??S4m,"w`vdER^
@=0TUStV+pzPvR@R2>RtJg5/Nd}:\ep}kp.-p{SI%
{<r#ICF[Bm4ltD4QYVx_;y`9}
eX3
Q64!|eEL{x	!6[+7rUKqDGD8e	^K3 ~`IptFy0x`200,O/Ga(y[q]o@)+Oy>	q<S}5kvJizk;5Kb(AEPL3nsXB7D}tq7s^"Z56k50syD+I&=\6[<_qK
VlkcF-H4SoFYeP!@mb-DuvGU~R,+5{4|rSaGGOq3w2$d4xI%&~^"h='Veu	,'V@JUfJ^_H=UvEf&{AE5@cx%@ck-8/@$}z:"J2\eb|_\kdd~&:B5	(b@ATC.mZQK6+tk4h|[a^ng/8Wc1]!8E}T(6UIb1-cfO)h(W7o&F5%MQB,^vLA-'oSNQB&J`P)}J&Yv>B$;aVjFI3f
xA'5/P0A?SA5fD]SO-Pr+LCFow_uW,pM\OSadyY7-:;-^hJ;r;& {>F>fxqKqj4#go;gk=Z!<6uj=.&uA9qqQu=h?a}Jmv1@,(7tW{:(LnEPgu|{"5x[8"p%n2|p|8<4x';;EQA^Anf1Y=_gAP^Ge<8_Ss4 GhiKapH"ail]AF?c$a%OTwbSRifICG=@4ukck&k1w7PmYbZU]Z[R=C"r56|K,Nck!U86{N%s4e)w"HFp|}x%Jp=yx"R'a6C)yJ3r(FSYxRyQ).yIXBb(?/?oGzF|H'Y7a`fMjTy2Dq/YR@h*gQ'=mTSiTH'=W$=m1"d;>s7cBVA_Kv}@Pnds"&[_}:*JO%-8
@w4!R"-I1g]'}04WuRIjOP4fkyu!gz3t;}6?pV0RV1*ClT=_X+bQIk#N0,*	-wxkB%4ejy~f=.R*
bc	U ;f2V-xSZ3j](J9$y_%>23eKp|G8=MX);b~>+oj4_XGv!@Y}&^DWc=Bit^VC?cUI:]StyTafwDOGf#mE(160#LBkT]&iX{^I&]7Ri>ss/?-wDUPznv!0\D, vwN8wa%pc#ug&!=5b?R]rJ@ s)#FM}?>A|B7q1&&IW%|oh+a;(|6KzQacBq3(</Fg"X{W'8GC4Msl0b2	<u{o?jAO*
I"}GDeS(S1G^oXn~In|.L>[:[U[Fvozl*:,x+3cU- :AV-
,8<Q/I _VEm&IeQ_<j``&gu=bbFExlWOn$ClRmxdczs^3@Vy6o
/h.tP-c.qam[;p#][yawUJ"met0F$y+[(!9U0K~d3rzg2;,\t{l]i W^j)E=/
jHu_dcyjSDM0z?!+dFyS3>A*%_gukJj+3rI`y'KemXYgOvgM(}}+e@xS)	Vo8\e=Q0c#=lz#-'aAn|<\j(zi"7fJ6=vNs:?!D"@Kb;;mOmT^QUC<ynNf^[i{)Bn^9E'J-P+O#/P\c:z*7dWY(;z'\?_B3"%CUY`k+x\Fm3Dw@"QLB9W)m6n#0gk@Mz-ny g1i}/WstbD&b,
9tFA	R%iY|zZ:JcLA~LGYc	EMsP+Gk&j4U\d'qS`uc%Y1sz<SZ"~Xhax-UaCGP0e-~j@('b9s'd2.b[LH~.^/pd?X:fB!bb<n!Y}$6q%bK@I`B&RAS;0h)]50S{v74j7E$3mAI@o+JrSV{d@5~N; ?rEzGaBAY&:bc?{-0=v{`[e[pqx]\<;V5aMDc1t^8tAb3}gl][|;t[ZD5X|c%L[X_(m"$DF<-0{2%{#@_&NSo/-T?yO'A6DEzUCkvIx,~V@?F#UK1rB(,iH;iR(}BTnsjkq]_9e
kjh-:kX1QJg/no/l*:oV M!`{[L&5%8%:xNK1zA'F"+C`X_:BKBC2V1mswfD*g%4PCi:#t"@ug57mhe}U8R5aBQ`WL]l9g!`#B	HNbxM#1,@sokf(|Xqa*k]\{Vj?r|`fCq)OwWfk,R&[*gO`C,Exrii0y0dWH.[%-VX_n`RvOKwWj]/0ah!rsrt,ZoRm4YW"1]VEyM8vd*CdOqG'7sM#McmM9cNkPA{bWpD?Q>M~;mNIw&OpEvNvo_jr#:{e\{uGKV:\(FV*{P[_Bo@Y~;_>gixa3U+veqf,}CQ(6Ue172X@ZICs%H2%r"C<W2q	K&@Bzb.Ys.R7cna/%$VAV>Fc{X
W&zbXZTm)%X7-l)K/O+1jAHh$QEc;=u!
6.L'B6;?\x	]3VYs52D9,ES">![*pf3qx~<rF[=r{05'A#ahRe)h<3U<1)NRGwd]P;77Q<?g\2;r]?V:UM*]L[1S26arB_b85.45LXLr~gcD0j'a}yZF+Gb^3bsOU}m50	#Ocq} 6>"T5h.3MKuu49[dnV7fjMnHzynG!@| 7JX]|)zRAp:!_~V7,bs+v:2g2Q:
~Sf?D6@w'>,1i)h")iJLQ(Cvd[p>^=(DY?#j{p-q(?p[Y(]c%(a:m%m\4yt$-_[HS!RR9=+DF7}6DGO!yc@hV~s35SdO9uA;S?wwM|)G	iQyYQqP3-/BxrY6AG@ivnlxY)jGY@"yzVR@<7xk8{U=r
]c}Ud4|.Z{4!~9 )Rw`PsDBk3WWT2j.ut1mMuU>HuQVUT}AzV8*[Z?BWoS?[4zHpS	q_Yese|g8hv~`P|zb`;gzK?seVLF%_T:!;JT^"[}i!k?'|g?ql2,K3!)BMjVQl--TyNUeL,u0n;EpNbn)ky
[uU>BRe"nsp )d?JFJlLAQa)*v.Gs5\PpMK$M)?*xi%Uf1-}?P75Ib+h%m1&4a-U&Z7d{m,dw\zmemH.;fG/Lu!y|&02a3rGC3wH0URq>2fUP:)|5,<+OD]8<iz"AY#|<SWCwOl[ @Iy)fw(AsZ(WW%,+bnrgTo#\Q3g:1vXj@$s:6a#]{3GKyTY&klI7~]7oN0bpwOj/]k+&,`=a[T6GZN9Sg2RSt0Hl(4>kg|P{' E`Y^7<Je;piD#>2PItB6M]NeKEwU-Lr5IvH`3=~3LPmx23uGm69i,Ph[j^'9FINaG95V@\B^r5W0m$MWhX#IqP'#Z7k"%~],pGPz.9["|%EVS[=3ukCGx~[V(0]C-aK$]ds1mf_*U7"h26'.sbbw0>Ccn&e8_Y<Ylhmiqv87U9@?6URXmZ?Or*3+em_s3>=? 
	@Exfytm
shFY8?l+Hf|pP-zMS/A-{L\4/ ^u
Bs3m)qomcDVwSN"g^&-bp@>qw0l,0|B|YXDjC'cDVU78tL`n1.M:a	`;:M~jltK^!wh07Ch4lI(HD_4eVHq36-Z)qfd`y^q
jL )if[`I=edz+=W%\HsmFS	<~z[{OG15JGy=ihnF3P*F!8]vB:yj x*
WP*X3$z_AeE,X@_).Jzaq`6b=6w{,jn-5>,l3Nh_eb>{;hhG,VjM<qb8g^B'3LVw?M~1Fp(BzYtIrD<Pyk"Yz9	tNny_Zn0p6K_TI;~/B}%PgMG"4]+eR2=M*V}|PIO'N1=e[>9aH,RMsWu4vR`P40oiVtCzjtb>aZ_*;ZVo=kGY;XTQwOsWaeBABSAV`}:,DZRLK^5u;~?I	TI35mNFhen)Ib
::/u;Dv!T'o6l|Y7(;`+7Aj:J[k(WDa}Jci|NLYUVrOg(*hM1b~Xt} 
gN=}fzop 1v|]m^3r	nV;LWE3l?DzD.w5.hH Km<L5,I*MlG(@]i~,)eioZ~^?s|U=;l>sCh`@*<!3;`3r,*BWqE>a}0$VbW5%[%5A2?&H9y:IQOA9bx8xgOf -~{'a`gg5x8*JE<ZWyq9:Zo,GB#YhBQ{!>QALwub(ABZ[26+-ln0`e V7nP7n4>lB1;6o`w9T-.P)/7ePk!DoY+*D5Wco=mp%60{7Ui"j"?<	%{,$d[/OH_.F7Y(K|K@Va7~
PB$RNmMwA)\5{]qiE_YP$Hh jefd#D4T`E>zMHMWA]F4C`hTj_19Lx*Q#JYbjoz$G6TnV!FlUowg@'"w0(:A56bO,,!L?B)[oymJf|L p2-c=W=0e
 e6|O[&$$&*|v{4F%5-cf&'~gYTSvK]Ovyr!z!uBpP_LZwgRXF[{(8AZAQA=p"s?}u,| 89BF2|R+lwH 0{5loNCbEG'aSQK|9o8|TbK!4n-b&/w@'!nEmji>K"M>z,Ih
Q<?~ab/vB/|r{X!zQIC@v~vYda vs?Ls-0!,avxY/v6apcHm'54gP;lz'hAak$
B>~M/^)} K.oo:E0k</	uk&Q'j"$}O9X)PL {W%C.b=X\m?r]zKAvMrCw06dRh%.u7__/60c%ozf}.NF~p0RR_tg/O:7w!f/(aRZE.56Jts-Kv4l 84+er
;[F}V8i6y8+iA=1qQ"nK+~bP@F['],A?Lg#[5/EaCgtA4z(f3i$SpqU\H,&ROVLuMYve7}~rVDqpfdGios$:(!'B+_y(m#ipLG&&5x@&6b2Mn*f0Og2ge0r68OAma$n`3_9Gz$
^LJCNdV'<,B2!EIBkV=0R;BGDK_onMc_&U<^azeE3HZW!;<@t'QmuTB]L'}lv[Mjlq-E8q"kSDGVVI|0i5cDOpj.)Pr(gKb
DxppLV,'Uf`u0*~?hOTDhTqu c%X@c(/pRPd\m[bWlDBKP.lI)S"`]ug^+Y:r<%!r015`tU8ZipO\l@JMIqIY|l`BO{PfI6-k5<1J5Ue IjveAzPSVA7H*jxX*']xgCeUQ{b"	[1{t?(pN=A%I	j43}id@	U`z*I!%}"&9|3eOrOrcTorl^3'8G$j8TP_j!Sl`Dwe
ijlT?@'P# dtd#E7-ArYEb9NhlC,[3j{R
s	h_Yr.aB=^WQ"7F~4j+}xz'
RMiRQR+,a Z'<g6.0SX8(rVSW~U?8DV<2)f?>Jda.maW|qka0ta.,]n@)L<oV1n,%P"MN)a8~i?2*`:4vBd(~
+f25o'&ekUj^>yvn5KVD2/>Dj~XNUX%HaI<Ia(EL@%Q.HkQ5in$htPe{zw[[yWw7k]>bx GN<D2O6\U8c* S#r7sx5A/3B>J:kJF)
kbd4#_/;3GaP@[QK6E|n9ko(E9@6#Uz^`S8y`VHD`]&-j`g\#LVZSN|}Ncl`kv//*R?<~zIaL}'zCX*ak_sJoF< G{tp6m#boYGT3Gp:5Z4G+k/@kJmG
K	y^{ =}j\zPES>qttjjrs279LlRmA|/RKRJzyQTu"Y!szGs6 #tO7)?3kc`r@H'zYA09KH.hu,<z7#Y1$+}]~03
L;3qzNqIM_/5`&7l^!9/7m/ih8D{ei25%"j&`GiKgpQV|+$5A,J:$XYv@PyuqEDdS=rN{qZoq-$FN{FZrQ)Yby_3(-}\jO#l'g_HWSq<pNw1mBoYc%S'.%n?DG9.^l]	}xqVw2+S\kdPND-tLRUE3"
6{g}?9$Ezv	{t->sobHSg+X[MApl$eUek*0/NvPX@G<K|c60arZ0^yGzp@j_TB(f3}?R._2{mm]Z/S?25`[BI7>JAQ.
^N-["jGCi0zI;t;P9_4oERu3+L8`T0S>LR<05[(w71A:@Qd+W~F+GFE &2J#>1{\ri=@3 skGqm{Kd~Q:5~:RLA_btpFMzs`$8xZ`KvOgdV
IEe8mwCxl1'wo#wEn80J/{Y[}*	.]|ZBP@=x~[?f\q9xj0kgE-UXf>=ps\=\jcu'daT!5v<TCDB_e]-<7hm?o0%ni6i%cq5jN|K@$*q]xuX ruSiLpi_^%*	e42T=)2d%/wl(L D-P}})u)3$wDZ+c=g	?QTLU_7<(U(JbABL%:e'oSFv,2LP*x{bHk[_p=cHE.<!g>6G>{-6=c.s ,ak$qzD9M{GPzG+[k[ `=RA-1a?/cLi5j.mB^bxWJ|?0\Z~1bQ+5L6cW8=O-U__I#veZ%4.]CC{\oo_dm-&`B*AM/_n6<:B(2Ru`!lKOhK6q(mD<8@;[gsZ3mK8]6b|XI`k3]j o5Mt Hv|F,5.Hs&"pPKUhrlF;r'?Y;oEg$d/F< L?!fh+\CvG'q2!XIs$1"XfI q8sXP{K 	r+d'm@o'\J#jqWO>Cb\	[j&|uo;K~}Q0).bJ?)%K'yb.L#B,E4PnN$RZjj7d|t(eS!%+C4^h=aQ*IKtKw(I^1ao `4A>em4$ykL3'TnIHmt|zqbb0JEa]P.bBl^2B>#'.3piarZWl(`a Z{pz?X[	Ui1k.r\/k?:rJwjs1i-]XsL,nYYX1F1tV4d+K#T?x&{{m)Znq|-=wYweJ4O^CE>\)HgF2]T=4B(`qNhe V|K9qwV%&4g[x-C@^7`@Y;Y7mapd8%CwCWCp^wFp	r9|bxe Jw8L	<)$wFH4oXg5f0PCasWxW2kO^0"	`_4qAwI3v6R"d,C76.Aix-b5,Rc-IcuTL		)arS[C{D.Y >E#Sa"N(oHU-zfbBd.#3j_u%=[I	hhS 
=1gRUM/c~DnJ?%z"70k8JY=tG^Cq|1F=fsP1bgUuTMtvQ|*(?}Q8vCE-	XPk,O3*oyYLKVO^U@^@@]92H1fTs3*`7"5Yc6IOryCzHw,9!S&BJDuO}?yD
@Ne0}J+e|H5wstCsOz
!{MPBl^!aY!J;1jyTdFQ]b 2b1S%cF.o	/ad<D~MP>E?s\FqiQ1dsBk>CK"M]Wn_9TV	7!?/go
sUL_&rwtADf{o;$nd|+a|M"1//'Bye8H5sWlV^4t1O}~t/LwEt)jfn5pZ~XE?(`d6hsbkzmoHD*%Hbuu1n*$g%q0LUte_.8x+Z~^\Z^I`)NL-IMJ }vKR Pla}o.YgFS,@^a**w0g,Sn9]JEiD=UwXPq	5r"hyBlT@D#_.V|HbGdQ)'^[HF5SkOLg+)6,3OWc}v/'8B;eD6'rmbf;HU$[q=T)WIyax(ol]^+\^K[iA#)Y6Em;<X;'U6X/5O(E$;zWlySxq?fF.<J_e<<O/TMa^vh12\C&SidTNontJiL*;7js_!3;w8qC<8k<5ZsjG;0JY'edMM*65V2!a`tdQL~6h-iP% e>nA-(l|xUy%
8*@=Z UEC)OBiv9B|=^zcc"Z7\RGs <c{urlsl[6q6Uoza4iAVcKt!m];JEexxNav%iEa5eE
T$o}jk<>G9|QMI7%iwil%+22}.@X(z%5CFvU Fy$r;T~./ Y){>GB'Bw;_T]i==a2rq!423o:P1f#~vv#5X)9vn+D+v[mD=G1#Ywo	)pZ|mw7H|ahqG\FrEI<>BZa,?JaSak,1qijQk&@k]
P%fr[lV&aEhN$l8inTxOW}^U%H}}@w*j9FO``L+vz}?qXVzdp)\3,\8t&N`2IPw7>at/`t4h!B7=";MJSwwi:@b?$'TRx]/9#KFk\J6Y+XZ%oCr!J07%ls)/x:X{FuQeoOWE(l`s[jEcR=:-pzE<@2&"[O	6n~5E0	3k/}	MUl6dV[gThXMO=h&M(k?uD0qN%}MPZyl6+L+rPs_RlqyDX<DUl%4Wg?=]/\-5b_x?K"WCx}M',<o-b2MB;`~1R,$B-Ln)G^V`DI.;<i0tX{c~V52G;|`sc$v
*`ap#"",7\U0bV!>.ez%5v|yw<_JG~]
WJ5i@B;O8()wz>qy"5A$7WXF|	9GmR'SE(\3A05gqXwD,N@UZK$<?\Qv=/9q&!UPD^0BYLspv$w]4Dsy)@q7!OErjGKFSz$F&/d2$j-}=)ou5rj9mS'?Q|)z'=To2l2y9<df(8"p+1~TC9cn9!RH
'hYO5j*2)	WLW7i	q?^e=<#v_01$c5:$G2E_1_iE"k2A#Yk!cHr8r0'uONw-w^5&|'x$m_f9F(AU%%`7<Uf]	;&1 c3B%GNM/>]cI@}@DO
m
t}#<53]wc?nu#-5wC
nD&JsQB /RX>xO2"qx!FX&LH@_qe8@A+2qqXTi!P?3Z3bG'v<4+#fx(: /&ZN|;,D=h{uyyE$=$V3YE2C'@*S`tbxI7$kr}h=	nh}YM:3@>4a8GN]zz$Tf11p^oX7D&nV2PFhu'Z,@6HhH<sN;|}SF*nu<HgP/d>NO+_N,3>|!
&O-M<M6$G.wYYDG2WVkhXaQMG&W0_l:#x[KoJ[a8l&e!=m5,gj^`0}K(Xkf+st||12.,k,vwg!XyS&RSdpOpWq	|A[7QE-|is{B53nvQmGAU)*f_(X97H-Ek~$v]{\-y?DYRGK\t_ib?%|0r:$IHclRqM%iH-Kxn`o<wG@4Yw`[+I-)j++r+Y^$vhF3?0;O<q#,ZsF$nu}|eH^A#JYpC$Mc3|Kl%;MRcM!t#j_E)5&aP9iU'P=Tna&r$,C.eu@{{enH60x69KBT[jHim_]qtQ}*sU3[ZoGhWHCOBF<.IX8&A~a!R6<VMvAbrfS	ed|M3\YNZ63&osZ<\<A[XqiX93!$Sq9^7p~[f"Npr8<SE</MPzz.4I+D>\ei(m/_PC2x;2+"8!5*JRv/]&_A:eg&A]'6PIYss[L	6"plF]p%+sUz%n]G8aO)=[R`ujS,d%d$I}j0N12Qp,hDZ	X@iu_|RB=mxIUw&YS4 C7(G{}z``gUL}SAu7F|X>N0]!]-&^<7vbr6*9UWnjH58jrh]L)h,tHx,t@!{eQ|;|9h,HN9|#Mmz%.M8
]{cvA7Mt%<"&qU@-W"w??">=^,|1e{FdGkl
`DH4#gdwL%y*KgF<OfY_d&8qf/hbRc3!!nG34iG9`g4G:Yp]m'S.Vqb(\fYk]JXK21A !?[O!0j"h8dL8aye'$My8N&@s(('sbp5-n(n*?'fHvq5 :cDATu94OMofOWv}$#E}9h=9VCY?s)R*!>%92GO2L%V fpHd0*uA"||+zd,2O%M5-~Fynu dBuqX=m+)sl\[[u1WAx.{z;\"$Oq<
m%MQ-~ QrjG;*:Z~#$HBpDJ.E0t-z#)RX5T|A+7^c8N@k"E )h['eUldMa@q~=@:UWv:qx[jW4ulaxN;Mg0"iq,]60"PC/e`i7<V44CG1ZJ&	liFMTbAl$TkTi'P~1CAi	~iAFl?xF,-+mU[;_?^"H@BqD={9%1._T?3PV44r+cm%&=#i:Ysqpbtby#J6HdjJ3	;[_ON>9OPo`24an5WTX'{~3uM$_q$qb)KmAqtBbm@:]BBqyId	{oLFL5tXS+4ki W&2[V1QirQ< !	~?HK7tF[	H r]k0-BB.E5>QoKN>)pUBZaywpUZq(GstLQ6BkB$F=?k`f@*n4#3A$|6U{=4'6F>0.ztM{0k(hM"S##0]"IMJ8daea[=lSzOCf~K^(y[JX1c*0Q6{Af[1N;#s_.Ji_OfV>UE`^E5\*m}]Ef@k9Q_x/]1`,3,Xk"YfCOc(cPh<UkJbsnzL7Q3Y[R=X]8*eM81M.mJ)%cYu*CgVg=<X,Ec[+=FIxu ,1U8="k(5b	(_;Uw_L7{n?34qH)&C!|r^:U1U(Ns4r&XtOrMJb!n*miD =4d MeKZ"a4c@J>'T@DS2f)|"#S!\MQ@,dAY"I)sSS$S%2"pNg<MF/cH`avx.oF&T@!l?1:=LYQ{pDpWv}%*tH#$Z~Iz{{RWUF}FbK\)l(gy3~;j2<XGRR7,-V*Z4}X0wr8""[4VX<kQq]^YQ7(vfKVQHL>3H4U?s:dbNn>$M7>7_T|]_-f`D],|ZfC_xh$}c/RF8RFD,U\R1S'Smj=AM*PuSU72Di2Q
sC'Q.blRp60OTpj5"dz&k+rn`}[|C#BVp9|S/$*<*\juun[lotrHP~e4u9DVC=Z&ZDq]w#u>e7VJ6 9"UV:b:4x0T1b#xsr&3]Kr26IPVuu<tm?3y(?onM@IKI^GcUdIQ-UW#5Q6sHa{o\zGiE1a*
iP?R
~?aIydK(^C
w:cWga/.6#ar@M(A4-._h!(jw7;0Hou^\V=:sl`s_}f4-a!O; #Zzr$W>j\}obtS}RD|vR#9nxw8,6zqy3D1s"8q.$*#'_*ctQT:u)N[vN]YR8BWc^H_8z<<>ey7B46%=E%\jO5'/z"^
btic7~X']P5*{3ZBl3*`	m<Q=x>6-Fo+w}~(c"<+@k9cB|cM:@/_`MiECFWJ^vQ	[>
]%Kc_5
&C-_rGLw6ClHwe32h	44q#uE&+K|Yk2f'-^~sXzUbdJ,MS%Z<vw9c;O	 A/y@|[j7hBiDF"$oNCok+`/^~(|ey[lD{+N8[@0TFMT%u*bKR$>\F#EN'p0bhWk[V8/+
c%|~=>.peMcS(8k)/^R
^9	8)o'M_aA4>Mh^*~fT1.V%L T-WQ_'EfD&{${(b@vfLQ*%SB	tCkojl"-TyF?F#o6+c7t+I 7bkRT=U-/[}u!hyV:9@^_\#yd>)&/q3i|'sy"|#Lgs/+5i`cWQJUNg`xyvd)Lq-lEwBU5Nx}K^bs1pe2\T3CQ9a,}_!sxR53p~Y+7a&iL){`6g"9*,3?dQ&<]$6tW%X{uX2m^h|R@W0TdOca8ruW	D~M~?Em_Gv+o+))b6L("?Au6&4cKjH9?TM>*pc4CbC3g`pF8%w!oZS/$,]p	GRq	kwF@2$,B|8tom%a]Zc*X';)RY=T)Ea%fCZ
Y?T`2iW;V[7r}tFfk$6D|&6Gey2@W>Z~i9kXr[hiqD
]b<	Y#n)TNRnc-S=HCpaLa7'"<LbNo54UK7sG!?({b(h4PoCNwsE5N#z-NQ_vH;.pZ'jrDuY@6Pzg^nLI,^xkKc
8Gy>0]5NT`t"T>N.i&rjo>&?dWw*9rk4|+mN[:fx,5fg?U'D*egS.23pSx5X$>w:?ATPi4R>C<Dv"=tmIO6(a?
Kj3>m(S=}3e9b6;eE9ipCCVV
XLw;HGlz4QE,e02N#e~QeOD#a(>%P#2\NpO1/<Z^JPxZb0nhUu|<ul[lgH#b5"k|$xMEHGK3Rd#{+.Yn<,r:$x8B1S7FPVi6}=EeKFcW*{T?z|gdg#:=2dVS`,ly~F>WA{v]`sJ.3{@.	X0z8ofGq!e,_./ d9
:2EXEc"h%.cGA'5}X9yj/h=XR6e|*2x3))zyk6$#fsB[g@q;R4I)>urf9>F;{CT#yU<) A='UC]#L|nb%_VRE>.M+L7AHi7@}H@5yYK=(ew_%e}ZXHjsM'RH	5hgV<k^
mBrum*.bN8k4*~Hed3&ReDn#tyk2s}c %7EsxT|),[4-iw#l%D)%
,jct13wF~Ur@&Qt6VG(U?Q)i)oBa+s=jzJ2B.:5hK.gl\wY)xk[A1M =m6>{'n-Y/%{/VN0g=&u"wRx\U":Z<b/xjYHoc	uQwin6(Lw$
oZ?`j58N-ylO1O;"8yR?Q
MI`egEEv!q8I2^]b1\7qumTt`vKM2{MU(1l{>X`Jp|*0_AGAFJv\(+Ux{*D<htf?D,IJH!OE(*w5}cVgQjj.q+xbu:'Pvspnn,	+-O.=a?(-qg,[cac_	+rQ^EyMdqW_YK98<PIy`i6oP+2I&|0.9/WF|N*A"+gv`=mL!SNjz>C,jUtB|]f:X}F{I+]EI$n{E@4]G"j`*7_^]~C8;87M"HW{[j8P,U#c#RQ%Vl!LO68ySM1`R`UIk0fiI>B&3auPh,]HDI	&Z<3Ii?,Hdt818b9~>Q'v;l=]T~H0sC;7c",bazX	=.(HKZ"Dn(`si/q.-N/"?GL-}>wQBMKjU`!Y0X3 TKuY|*9q6$V*X%h[roTGnR`@!ZVA8gEgr^0?Wu .$p%@hFNK#>^{ wj[KVPFEhND)Ry`7`jK	V/MwA==w&$6Jw8^nz\mu;x&e7{41h!*`<We[-jyb:9};%y4A#[*+"
ULIxQyOJNp4Jt*,}MG]gGU/[yIU?A)T?\k:PW(=WlweW(i{~{`6:@NB?Ds_xor\+zku8z^nY:7lS{^pVGpj,;;Zh&s+MRas{SDQ9Xg)@vQDoF1hB2f@pt{DE*h-v0meq5lj#0H+,#yEaqA\	usT`F@x#lyueG^Scp9lZS&M;6";kX`%h:y,HqpszJ0$j9WI]yj{lz|w\lc=$V"_GTE_QT%zSxan^zS,@l~=H^pc(|cBxcht702*$Z&i\A]&[!wau#%]=%4e:
D{	s7c 'r.,U~W^U7$-7P$`^/dX^y(WQDY-u.6
Y>Zn)raWi[yJ)O<=Zi?
i*A6kiA2bmMMZ=.(T`+9GWha9jR]+gK!LuvEzEyCY'cYRJ=5T3 ?,j dubmmfmtDfA"KBzE(3+#.h/s]o3`e%avFrICg(n!Qg9P:T'#*>vk~']!(_Lti5%$1 >@ Q`ZkomN)P+uk0m@as6X;b9M4V,&7#+JX>lR8kD%?#uia_~&?A~N	{*}jcM
:&'sQoH28E|0ubpr"A/:Av,j'MlK5cr"F{E q9K-"rX2Nnk*VG	R=#:]7c{1hN65j`{wwW82[;t7KfIY3Xvi'?N@Z9zj	Y[iiewPlsod$e`(Pk;.fE/3rVbaDnVTT^OtE`9-^aaz,>^T*$,v?3Vbz;oFNYg%:c>K\ctOFLg`Ys:*k5S%;Lo#mT`"~eRn(l>SdMn;$,2E6NiMfcx(VO38i%&Rx	z#RXFxY6Cg-k8jbVTnZMzME&Q9LhQC;p1Ow8tn"YCp[gz	o%Z	BH2 ]P	(&`hRa'^A%O&(d2j27X;JN&kWPkwtvtWTn^cmw4V09v'jLWCPe(3R; c-.)05@KU}L(hoB3ony<q N,a$
VfX4,l#E2F};-!u@4uwyLtq|?4!x!42.3=v3"hdJ,dN@	y^3sF!UEs.4s]3_	xY."<g%'*bB1k;F"`k(`~hSk*__$FyqYWZk
D3&Q`5s2.v"RJw$k'=\Jd1, x_xo* ClEQ\}9
A^&Y-^4]8]Z:,9)mjk>g>teTNRK*.f#B<#W:|#t
MIGl5:]Z3}8p[ia6_=kzR&41Ls;4hvGZfYb6IVphH<}}E@#plKn	ldeb0RGd<B`CVI#4@l-c%!WL|;kL{Q[5QzysAbo'6IM}6sYS`)H8s$wM PqUTU/2zWR5EA3E_&>HDfKwu:Ho){-1+xAb-UP#ycdQzx4S=ET42'ufYZr=L<&1yVOR
XTARc|I*:C4xWN\2
bIhe%m2mU	Cpv'Sf`=WldFd,
/XqGU|0#p^u 'V&a-.9l%M=9t7Yo+|nf;sh((AP,J{`+p>gY>a$"XC^UJ(F$?5O( tULX6JqjjzDe3.$qWYS@PpqS@oY>7<`2I~=f"!|a3HZ;|%lQ76oik,G\&!p|$_Wx00["HomUW/6T7@M24oB#z!]e{:zA9USW&[pjul<& _b;	+XFZEtr",Ddy-!)=wslJM7>H=	'p\[d0Na[;b#A<-t9<NNV7,(?yS[9i4c0jS4\$W6LTTK`<$7(`lYjqA#,1=8Z5QXT1N"CPZyPEBXJK(GyDPU&)sd+
e8sf?q,Q! yFBTT2gTG62yxUS)2eRR9h3JHc^]OH1[ix7+n"@T!nLm@Q'Zfi7c/z	i`N8sW@yB":T	GxwT>&ugD/c+kw.h_u&*;lYMK?^KUPV\&E`geU*jfSa[	6*P=S:{U&]" [(g8tH9vM`|{[u18fiR`8)m'myNQ?9.S^PSd{G\)A8sG&G*h{H=!"hz#.kGB.b\%H:9\'mcQT/ll5_9XFy|s/w2ylQ61d?Co$ul'QCof{>60T=3,2F,<-+xm]Mb'CBCM`joTA?RUX3m9Q	"SUL#OAu}ad&6`&^Wq;{w1Q"#Uo1e^q2E2"K>DF/]N2FA|9%6}~2wJiu%!`28W3zvUA!X<Jjm}xron2sdO]m#7z%alHV]R<\]#$/QNy).H5u6ppFy-$)qdcgQBtz
.,ae&7)GWmZU"eZQg@G!ol6mOR&4YmF-3Wmg)pri8&npL?L/oE%ZNr4<tpy",) iAVUHoQfkGPO*|VJ\gwDK32It5+Km;FdV@Dlm2u^EjtE[Zbu>xwfc	&=!Hfo4&=svU2|6=0|'?8^dii~8iVg
G$P}'6jji^w;ISRzy0%xaNdFwI;r3"4G3N u^yu6a$$fkZ'",o}qE29KQ@;<ZpO?]@,1}pd.>sm;l$A+AP-/4WaOz!rz?aA09J U;Tu9EWF)dmgn%Jy)5w30G4[,Ew:6V!4KC?C$Sa4,F-MWN-%F"l^gEs7#kv\:16*o/.Nv0uj\CIx3&Czgv`X0]]CK2^@cpEC^a(Yx-XLho&Th=^|z^5Q)Fb0hV-{(SX;}%3<6X}mKQ:nq1Zn``$=
j3y@n{S|3?EkSe?U(9x}5di(\sl>Ah(G9S,@ilBPt4zt0WW*M'}j>Yl^5KT!t%^MoyS!{5|*4c/WEr^O&=$)&_2hY:v4x@-X:Hr{W0@4NWNdw)DiM6K97qVgK#*
(LW-(=_gi^wqp`w7E\;v`P(j]vEQnNol0mg]]_/?wxi>#+}D-mz.`72_.@&3i*G_3g">9}qY|B4I)|V:M':T:ku|G\ZsoPM|`UUxfQYTSwn&&99&<3l55zqu~)k,vJB7h'hZ.${RHe5@	23ej3'QcOQ*Q [D%v5_6e$8jUFOU*HhaazP{Uu=i//y7(VW?dVi#:`+^<+#xG@x+9iN2<3oNv=4TKS>.nF7QbWQ`KX@nJb]<`ux81k(fHv8czFmRjR`=!&:1\ gq6yV}D}=gj"avb4'E85VD0e3-Jwz(.m0:"ND!#-_aMi=*SAX9-0Cp4%XF_gE(oVy~Et\bc#VN#wY,a7o;!N/i;ktQW	ok4+<8I!]mDHSW/d+3WI6MS4sSSW7;U>VX*[ZSu73kqdDaP+s8][=W(qt]$ X%4C7-`mG|c3qxAi|]B;EsOr?P)?f96sea$Hb:wnp$ml*p&/`FJfg	+ed<azGC[SLp&B3-ny,:(z#)&Il[5Q:(&,tra{y4ftS-<7_yAeO`>Sfs.`*Mq{r~3D B&?UKP|;Pw`-iK<n	Eb|FA7uY%"B5O|4)0.I"@7MDo (3[CC&-MXwe)TJ`p{.4/sYv~Y+C9*]p^#V$Yg8Bxs&7rI9!^9A0A$+44yGj"8LxEi8S}1=,!_kB6>yp1]z( 3/F-F
hApc'G1-=WJuH-
:zhr*\!9AX	!M>|
;N>o~a8	r~Ni[:+I"C1.T2Sa5%s.dkbxXJ3e44Ix7}c8 rr1)J"+(BW]Q8KdR0+x0OYLra}A|<brOe,:,1mY_ll^=BS6GDa!j*
G?`ZZ~	dQo1v8sf0lr1m8])CB 8z[8C'>#5[la8z6:6[)9I@,"`9^y*H`uH;E
AXF)u%lAHs$z<Swa}C@Zt]0A%+}O1"bP=qVKtbs&\RuNlSMOwNF*n('YanpJ4&zO";Tf\Dk2<r=r%Y34vnBY`oj)]_ j#@gf8	nAOr9c]rdKC*fqy`CW61A^bI1b*dudAQL8J;GmtN*4tKo4sL)weyo0m?bw;1TPut,:bAxjfmS=	}zD9y&$7
oIy`::y%s!~q^$ W#US~iu.kyC0U!=:Emhh(e)q$'5H9
ZxD7Z(0HQhT*TvMRWkB.9p^8wUTx,Ca+DQ}{)R{U2~!$'L+L%	jxJD4?oaQPUr30c?l0x$()0!AlyLf{yPhqB2!YbSJn81@[6lY20#8~s\T>QgS:~LLF9LCb+$Y\pXO~`wE8qOPL)C1DhbgRG(-JK$.7q*Ux9T3_FH"LBs$D/8{i,%u:R)UxX	1@l![-mgH,oTRG=`S1' _wX.Y;Its)RmN<"RP[MU,ad6w3)J6\
.cE{(AAc;E)NMK>[$(JLb0IjxB1j0CcMcEzu3vJ+)_c|'R:[lv]AEPbhB<'S,A+)pllVC9Ix'5'cE{.iEWrf^%	Z7}::H)?!S[oXwhkxbH\.r[-64
8)k7J/g	,SK93>5'EtbE25$R!Wmm
P$f)qUpr3uJ<&V 5IAkU*lFda=OV'3ghReQcI[R0~n6X0MWUf@pBtqPD3uvRbQ+qocINRN9rwOMcx#v_bJbc`~)I'}nT8+2%"TY$%YgrnBT5hd4?^DE89\_Z=Y7Op:qhofmvtCmg+&S/DxT9+>6I1
@B
U
(p(Unb:(=V:,8+;:bJk
9=J;tIn#uE}m4,.kkU}x7f~Q5Ki
b-mBb9]UZ|_=)_OEeK^^\UAE6B'zlE|d#8Q2g=Zt<hB'/m9N]s^E^A	=,PfK3WcIH$0%Y@oQ=UUu ':h<gyeP+]iW[f0rvxbTL{&O3T!lb2^e@g_NCoRik#KL8-9y1Cf`'ql9&P(Zi2c+G/k<t/Cb Q52#7`
E^$|Z><;M\jh4	CQfS$,CE:E!y.z*m$W'Bf%H!050WEI*dQGJ4PE&?\?37gD"DQpn{tvX6(fB*u9Dm{V#AYdNGb]V4'F{LI`4lvQ"+m|#0yAyqdNwg5edTra{_kK>^j}D;i%yu=<e{praq6S[R<)K2^	IQ\^.W|!^F9dvj>)m=IS^:6zR3&##}N	F@RM9Sy8~u3{v`/GE0j=XRV
^Mbg'*Ea$Vd}$6FH*t!{e\w;^hU8TX	`x/[j%]Qj&^}R!/<a~;Wu
rDjI&Tm3H*0@q7 e;tiU$VpBOT F/xS=m.u02&"'y/d.:[:AM
72.!fH4ru2]uU9)5q[?d{xZ:#?lD*[\ChjrU Az$,}Hkgj~g,\X.Js{sKfr*\##MXU2eY`m)Kl|fd%]rl:?7AV@cG|B`fRBTs,yj5h$"(rDVfaN\VD
l>LYVbo"by6$Qk-t sIRIKAK
e^?-L.qd<ym$16|RuT\K7<=}&`~[*F~S "i*u
Ot!iW`Ip|min4k)iA@|nSGP(.S(hZHhv:
B *Tpo9xzTt0<\uju~gThr&
j=F=eJd_.S. \rra"%>t'jBL28y/~xiYe?bR~|r"]S};&5~C%qg5b3C;Y-l!{)E-.r*(z!rbn!WF^g&(Ze1Nn\	g#m	hd`9N
FHFv<";]="m#5D.aU`wh
o#!$-CME'D7zeaUfCnk|kh6Yix\x4!L=0~}I83a1*J\s&|Em\6T*FU-*5AX&8%BE'0:i%be(E@rlazi1dmn3k`c`Pw^	 ~z+Zcf'OUZa90s0(?1&e{/lFmxhee9"gFb4&t",'89ds!,F_KIwynx<_?&r].|;<thEJMEpZDU#UK~&pp0kq>G|$"pJIo!)i&+l*`
diCnM&E`lI*9L0(Vcd`bti6Li
?$<{!,OM5uH{`P%~\a`Lx;}L/i)Jl,'Pi4@Ca$W::H!S|KgOq*&4#SvulJ3Y2''dXfwi6x
\2;rwOC	i8b1Shs $5i1DF>i)cI)Q|'
\Z2"W?!R"
%PB	=EIN5GP^x?hS1Tm06qD9=:8N'MTJCpDW+ 7u4adx#}yyh:I}TxR<&e"gt^AOECf.,F#Fa3$Z{Asw[P.T^$9/-T0{tz2[;e|.@)m~.OJbuoSErny<bKR!v?'dT>OUzl~.f`T1	HDNSw"{?H:?i*1&wYZ5vS?QU{*RoXf
>epB}dN#V[okhW4G2k[O@;QO_B_87BF(WT;_iJvk'q`_;%Z>{8MJrMlKoF8$DY*
$~`mI&Qac&wf`#"=<n'g6aj	v]~O@DaEHe^=MW[

@J]EFo=!?K0zJ,wgpe"0eQDPIa62A*Hxow
0="hSn{~4NTZ'(62g`
Y7U0|8Wtmnu
]C*8FA2!PPyr2p#nez&l)`BIeZeNp|pfu2l=?WHDjA;p wRVHX[fNrBcv:f9~%8};&Mj>@jETxADa$?e&,GbV+fc>2+v^qsCcCr/Pk-u?<Ov!eU<e;?vFZ:Aes5u<rk"\w~'{M"VC-	lHAh W.!1&\N5VKS!2a1q}OVqhPcjTtHq-9#e7UBOXQ,X0$.av.^!5r9f)Q;g!yD+'wCG>>o"Gv_rqsif}m+ #ke.HA(|{c9By~_gF3Q {wVyE=fugpo=59v"v3@CU	b{8WAeYy-{C3dsN83i!N-`=Ts
\4IxV<m8		":z?SJgb& RPse!V<rq&>u8;Y-I}6syb@4 nbw&3_JY
lV[=2ns^wf|v|<o`9mK9LfQ1k,ir<N]gQk,[8b}o(c5cmS[a]IyvphXP7bjw0DCdGtW)A{J Es]c.!Tk4zbh#>irAVnq6o%N/3+q-HE.$QrcF5.w8oZ*U>jE3'-E[\OoRTS(T3tL?#'c2-YPI$u}c *O7==PtvY~|}e@U#)K[u[w!Kw-M,l]%+T0ORiOI0;r0P[uN.@[G.Nzcud{g{DL8bFk;9>?q\h_P?8,Q)hexLC#pMX\2P?yZU7.Af@z^g+Tn._4J__
?z80r^QO#tzq+O:shEcX0uB;Ee2+x$2e!U\y76veSVz7	H[W8V:np
lLC~}#;X'Wa6_X|(B}(H#Tb"0?giGctr#i"X6"{'KGS,h>_NH@F4- <93]Lle\	nDY/V9Z8&~K0Cvs
9E%P
uPjG%U\TB^Ke5;m%Yg4c^:YpuVnp1]JX+}L\GBD(V/9D_4HjPWi|BDS	q>m30sF>cy?CeEXZ;
Vpy{be7^MFau@nxGi(`PQ	^]Lu#|v:KAx9J=>1i}XisCMm@T93L.Fcq@@`3t$'|Xln_rlxrtag\y	t*z?SU5H`=L_&L5pz]tn|d%mHMjG6So/xAMBb`[X$+k&A	6u_2<;[j"f@|l.;-YhU1o=Rtu|'fk)^(3ovR8yQ_?zwq^yS;n?]NwQo;`e5%qHe`415tnLsZxY|pm/RBo`s+ql[;r>#[4Nc[NDD(aBDSK:oD2`(^Adx/KUIL;i~RZ>}}P;`"qb@Gaa>]|3 :hl2"KXIM4*u3!
pQ>d5^;jT+&;pzFOog&MQisK[v7k, `V7||PRJV>Wx8Z+X!}8kO<Y$	vHVZd~&YZriG)1bBzPg3mBz5qEQ<ylCqjt;`drf<]-Rb+R6waNMG*9z9hc'noE)eRO#gJ{!BJ#~!d#=r3!I/d(L3Qm[^(;hnYj6s&<3hMXi2_gu@yM !|fk?j[!P
__MpD_jlx=6Cg\PnGv4RBGu:Nx1vsP7an'LF%p]aZql:[r%]"x=tC5O(=-\?Cr(jrSd.5#3M+kgmT7p%G`/
,tw6B8?lo-<?p/oEeBoCi^lK4Ee{V*K't;g4tW02jH"J9VJK6 @wnKfQ(;$|I5%zvR@]_wI/[2C#rdN_ OIVWU&CfH7k~*9C3*4u<!	P'8u2bm)R*uYz:{UTV>zCRbm7i{d=NO*-V=7hN+JvF84*pud=Tw<,-5FSX#HV_KGBSGRCTi,KVAeLqrWcL(Zer4"bGwRM7&uz6}gn]3K|MWb@v3P&u}0MR@tX%ECqO:<z <m=dL*7k_P}K]V`^itF|04MrfDh>*R Qm;"77&3Jn))&22YlYM\8yklc!U2qCYW$X}].g#BL<@?U c6cg;/.^eJE51h@MRM-|@FEF[@DqBHYrjXYk0&c$j<?O3m'A{Kqy\'d*Fx.N#t^2VmL?:	Hw-Dz)leYjqS+<Y^ab9GlFHp4*zfF
ntA>s1%>D\fO*u3jzNn~.`-<{o$P}Mh@jTV+0r(xO6@FCX.q@qT|#BQL#!v_3Y`	K`kC2-nHhY3[sWw?}3	u>WS.uKFCZ.2g_}]^|w4I<smKp[<-xt,~?hwuH:K)3{Y~}J(%bNtdgEIOc\NLtTPD7%3ENjD`Qb90}5_/MotR\YQ`S^/Y>z'qH%=W):Dc<#@QdJeB%W`;[>k#^_FRnlW&
7G	m.,*GNdrJ$XvtbKsokNbl(8Q*)qVt.EKMCWQ2NYFh	ur[y9#fMD77 zFHxdP:]1wgRPfDeVn(SLVr.-k&D'8xX/$9}cX07p'[T_J>h(+1&P'!N2fa;5/v9%_J%[y`q\1oJHa.Ni;iD)N"#liL?3JP]xDDoP!YB/R\{1vjtr!#FG36UW,:*XCZ,@C*z)<R}$vRsW2(_#{cI3a0ZBh>qonlm;,}K\q2,88A48KW^KB!vvzze>OS2n/tJ$V"mG0duSBb=Q
f\q}&lF%iKw\EOY:(C/<LE|2 $';+J*=]\3
)HZ\j2TJl5-UD
QKb+Pl%W^6<<Z./G>_CC=Ax)',BcH$+h>/Cw<M=j}2Y",a=/}`5F:q}]E6txf/|]N62J[a9,|/<>65X	hRJ:bO8f9	!`Nf@EE2_xYskt$?1t	o3Do$sEtoLtfVxZv}rf^GxEN=]fPw\|-crmf1Nf_EX/C}bjCK8u$&~Kjh(`d/Q-C 39-j'(d*y
9RlsEL]{&hgt!]w8F9I"O.KAZyv8u_e9j9g.&]./o,lE/rJ.MEYpqP>ivvM?!@YQ3%/f|f$r]} E\jAi #U.v>v5/^&%B={z>$fo1]>;kIk=OV;M8tkvH
+A&ZpPXB.sVlz: eAVMR`H3*R<`a x4)WkRo/4ULn}~`.yra0Eq4.n8'dVUC%JK=-eagd?U[sfc?`s*x!
o7Mnub&	yuaj)7x?Wo%bW{%g*P5Hl
]Uj<3/q[mb
Bae<Dn5t3+#F]#	14a?v1Ic$Tye@fV>075Sus\s:=S+Lt[ HjIxg:kCX$L@A#>i!);,P|$rcF4,zsq&\a?aghNc]%8?_+mqe.c^trudpM7k9A:0[kCOWnW!')(HP29q[!%|197&80^o=NXsNiz1A+6jRA-D+XG?l(fcP34.a3k$?QMk!:}a"KH2I?=(
i/g|&H%&sC*`Ec	\[TM0[n}kfn.;I@H ^.&a=JU;GaZ]m[)O;yqsq}4C\uA#	>5mVrXD*29wj`ostu|[tY(ey!v8Ft3F)mBm\)TU	;,96pqclddC]"A2b!w<Pl2eugh[k3IZ5L'r5nH]G[aQ)UnlQHh}.X
#LqT6GY*|xmSlK`L4l#F^$->aK=Um0Z_c)S}[U?Vo.w&xn/?_!xM{~spzNcL0pkC9oP]Z|DHv\jrm/QLI~#!g6~cQrecO5W(#3!3@DN	ZVqufA;Ap2@"7T6{3ll!`D{7ft$7.$r7]68
tL+2i_/$uc(U(_8,x0UtMo;kp2N4?BQMcBzb!
?w^\UDF\* FH/!IzA?*
>7L5Fkh&igh.`,6:vo]h]|7tVR2Fcxgi.o@KKEjTwB>CBeEWC"0}:7{;#]pq@g`tWYt6f~"pZ&C|hQho8y&a41&gr?x!_sN].27tl!5DX{n:~MBYfX"|W3A7"NdO~8niy-dpRufl9d{*f@9j~u>c.?iK7'	8&k+`jg*S4akbhO*5o@f

CKu^iwq=r!4/nf6[4R]"+yY6C#{Oh}}xo1@N))"+v,CEZ	uG"E'jAif6rVal@]Ih7B!yVUmMUQ_.(&Fa8+qtXpL8U:*2nA^[^VStk=6Ys`r~xS;.;z;~GQCh4(="$TPx}wyfN"nA")[eu)'718e!M>&_)H,R#o),*9(1epa|G
8hwELQtRy5Kc?IZ09
c!U}Rt4Vvlp8|`n+sdn`J#bZ@)||1uLw>Ya"N$Lp:Ds3NC`:zrw||k
SP)P|+\*LPddx)[JK(mC^c&H$5&]\
g;?yXafM'o$=^Bw"YJ5-#5t:;z&H9%P>sL5+zFnZbpYc}pCVqZYlyjhLga[Cr7.$Rpm }4=g$`dW\=CAo|8]!Cb#[>@02 DyK=QC6@+Mq'v1`&lp-y,Hv:2;j/nI$zphS#}B/{(=<M@}h# SJ% fl1w(U23fuu:+YRL7W[-Wig"&tteGUF',
iBnEzRWE}F!m6QQ*6mjvzJa4g &pi,@^43.56wIrr1ju!!:QGB,`fJ|&WH?ifA7m2Jrbc]'G;!ZLg~bQ/Vaw$-@R'D$q'/w!A+!B *cdC2{14I!BI&KLsu%n9_U=.?eX&:KC6?6Kf
/5o#G<dsSCT/u)D}t+X74T&kX!i/yyYxM *ZO78guCx35MNCN.`]$-\y|eJwgR+MHtpiN	o.@f*Nh
/mDP2
ZvPLD{{bgX+kmg5jb
2X#"x 9ShN)/r89Xk[&,vvB+qQB+`+`BC%y;[@0M^qzQ9rE)4w/Rg|-g< (?UoK[vlEBr4q"n6 M)v5r1-Eaei>T#a
?8T*Qf<4}Q`Q7}mG(#VLXTy(d<NoJjx|#AQ2#]XS94hCu	M&h-iP=R.%1nMuj\,k,=ol %A)B0Z?LziV"njiPlk$
uD'/C*{,`OE",efa[U9A=G]|w%M9\9fqix`'rol@6f;	!36)E<$\9,\ ADT:KT_?r?/EGDU:QV{49(@/B#I0@`T1;Us'qp:Q#S.O3xV8n{2`+O[?/`W&A@~Xtp|:awk@'d1MJ,DSLBYWha.LkmB" b/s0vgy
J^[_KBO}M~?oYj7|AF?D$>W6%P-KD!1Ixc-vbJ6kk/0IhVCBiArN@NBS&0`Np!,6qKKPD:u%o[VeCLKgr#DT7n_~op>kjL3yqC6[O9&np*F[yN1}`v1vkQ*oy "h2|sq;s@@`Nju<_apXdni,*Z`ZyNjBN;!!@<v(	JFWEFyUP*Dz&I/GhruQ~p&S(.X>0Rv(Yc| qf|[msU?>G0T`WiRa([O@`T$&U-E4	GqSK9w8hBtC
P[#3Ht&=XWAi=pS7v$^zvw58&0NyTB	=hFr2v>NDq/U"UB+J8,`1zo6tR1p
W&5,rrsB=fM^XB8]Qb/Y}#Ss<}a!{ZUv1lU]8RkUd#|%;D)wYo8oE]Qa\J4ot")?pD{%5{/mg"L`X1K^"ZuzR;4L
m+G867]wJ~LD}.,62n`{ty2S4Mx`kS/\2v@gx0H^6eK=wDx!>@ywWSpL\eGuRojj:09Ye8"T0>a+2B{x(<	}(3)G;HF;:b=	CtT\1,(IzXt 1).8LF!08Zs[;99s4`6Xp)+]AB@FCam_}"KP<CZ*H<g3/3QPOz|K'+-HL%Niiz{()4vnW<@F21WDw
/#8YNddE^L.&u:DA=(gP"p#fJ#m+n_ids"<|7>f||lBh	0Ez>Tr :a<LR}6DqE6y8qh<IO;?jf0>Cy8\ UE5-|jw(P1/-6+1_{uD!_Lml~bPI|Ln$|"vWFGG]3<Y0;#abAxwYS^Bq'"
)EY3>JJl9wx+DDUY+rP4$7jD@E(4sxGc=_Rjz^H[TalF5hZwy&%:h\@bP*5g	|i15mKqJQ	ie2WR>_Y><fD_g}e^[mu9=$GVI`5!|8ME
wmHC'`S:7N{=x+daPvJV
jU::b(FYHaX~7|A`iu/[~`2C$Qd"X
k+s{0XmRDV=W@^5&&qgfUlSS@90}[s'.ZN	u'!{JM"}O,%P":zb#;!hg:^
Tg;+U*Dk%*FOcq]iw:6~_nK9PMJ!P	Z38F$HCZGi~(b<a1rllm|$b1*hdf(uz71?R8/||vOnR3wft8WUe@ku _0^~K2k lpm6p7PcZY4-?N=k+G$6ZxJCL:gY1g-xLK}@	}^S#G<)NbG	%0Xhi4XCx"Ck8oZVVJ[Tl`2OX"`cY;x:oH*djEvVG}qX]A3&CnBH%ln4e_)$15Ux;iWI:Eg.
PihqL=CP?m{6.<O6?O\bcZ=u`ZXz~u%c(>46?h-Xps%5UH&x{:g6220NVM,{^<DI*ZFUK?kUxW<#%X*
A_F=^{5^I9j&E**d`rLC?@96axN~AEs'9Ht#.E!u33C^@{<b*	q&}K7j-!V2vRp,6~|PY_{@&;*/I!s<.QRk&(r\^_+5Xo>[n m )7o jxmJ"
nPH;Ls<9CU
9 \C$YBb!=w_L+-ue`Eymh=tN+fng-$QAiNzx*	ibvR+Y09?ABb1V23W'	tvQ"VQf)~Ht$}+K
]~LtN&x>*b,cFcMP|~~}YgJ?PP`yN*:0-)w?AenG!E526ri]{{0K%2|a	cfa;s,l
*9@^/lVH,dKeEurk"V{&*}SRNTNZ*O^&+FZ|

Ll}E;T:&<=n;LtC,7ck.1zFb*DPeC-IC*?3gGV;NipPS3Tgf).M*\j2WF)V[gKnFe	^xZjty70Do%0@'m_b(mS|DfPtXZ[:}="h}HD>?_4L?f"biwtL;Hl~b+`_Yc=U.XX1MOL:y!46[#|RCr&0}`O2z^_oLW>g=6Q}hx#dL6U7.3kO%A@@88MX"`r?PGpG*gGfkSoZu\`$cOe4T&`JBAkIt\7
l:	YjRKL+/g,za4;aU48s.
6zdwsi&@*M(a\rhv<f35:)FK\\)+]nU*O$
h'\"-(F->:+`}q-aJri3Y%_H{=A`F\iZ?z||l)R)vpo+]hl(R6L|^FA(sSEI`e"78"#^J-5pJAfd+K9yX\zLynNL9QOh'PTw0L"MtoAh,^P)H&u6tBCA
H[&r#mgyEmV3{pSIm`TGkpVV#mkBNl;s%})Y"`p/5p
|%Efc)b`q-eYP_%d?k^p]-u0>S[-iVdblN	CM~E<Zr#]h8*aR%-+&K00{)SxNk^`9ab#i$E4*iyF2=KM:J|`X2%,T&Gf{I=z1r?	~4F192l"/OUsx`cuSfbm7Oq7Hnv^
([c7wPuD70Y1bs 8G$+UD[Vo?1iiIVm6-I*Ss	@QWSpO^$OguwWaaf&"+/Sx:y@9FCXd+f7GJ>}*WN}]wr\^k!.fw-Y:(vf82d&I,8,@d^lej8YA:^[OtS\q.P[k>*<T^}d/Y1(4M0Js~F.+ng==j,y1It-QlZUJw_ks{%2)H+$( j?*MkYgQ}iA9=	 kY1~5DR
[?\.gNB@9%;-VR %E!Wvg_=+Nn5[(22cAQ0Jy@O(#sYOf#lv +6[Wah27*j)CNk8$A2> ,1Fj"$6hIsImjx[@"=N+
<[lFvV^D&{6m5<o4Q;~'t3ILg4Iv81kv^,Xvf<1d+#`uQ
+ha\#:3s<yZcqj(Mp/-I1hy.Jd&Y	WON]mV-}%Q#ED=X0:Y=6=[8#RTS[s %@Q8$c`SJ2muUfJ4A?)NBkO/Ibk&JQBFy@`km__]jlEl0qxm?8X&)RXd%Uxw8N\A)40/wk=e7=~R3RH
O-E3,fu%0EGc6~&#{:`k)gj-oCy:-B)Cy|pPIf?uuyC
|!:65-QH7l ]hGrl|)h;4Ecq%+3#"kvNQX6K4*l]K$hE;`(RnY"?el:n3{YIjuVW?VjSGQ"*k.O@{j6J)\-OCH"44|uWPWD<G19[*NFLzVi4?yn-aqChshn:+y1O{E-]b?gMy)I9E<Ov<$-LY=vyY;%,`2*"k.b;a?A4!X2@r=|26I6>/1d`e:k7i$_espJ>H3f#VS#w6RP,S}.]0'oe\BLf>=$TzQuR#P\#@5~e1'A&oU+hF-3'[2-WK$0V'M=B10AZyG $dVjvmEra*%AK|qUrSOGfI}D_X/Ax4.0&;#HaGC")r6RzeGQDsw7+De.(q
xhnc{Jgb/V">P|T-<wNKZNg~.Op%b&-KI@\+f]UR-3:@gkTVD:{:x6ok"rOQmu l,%;Z`2mJD%
QGv6`8s	30t\$Ag'={PA@a`\J)z#Wa"]fq[+k~KN:35It>X<9+}?u2L!_3L"0;/xv?0![)PHf/.64Ax$RJmB'}rN+tHn'n2R7sw'U*`!,YJj+oq>2vuJ~>G#wO]W\ro+`aF>c[$\3:Y;)~e*zGZbFSq7ITn=yF{_5]q"LkYz@7a'/	\U:/;wgXi3.e>Hq7]I5::0m	lNMT	=\)0*+EO#nKN/0TPm`Zw-5`ej=-~gmfa`|ftu}eC H2a?d4@eZ9.TO]OJ1W2Tnj(9<T[E @1#Px(HGJJc}dM$XM7)^-9c-*?='W!8LD,m~5azzEGt^oQRQ"K;6Nq|:|tg~20*%kYUj])R_l(Z5(~:[1YFHp-f+b;1Y9wC%E-`U=>xJEvr	c|r"APK<etGk4H\[|[-#J=E9{Raena2Vme#v\3I,+(3E^0\bdEJ%<>Q6KO9bg|}|X>X/]Y97VS&Cenn8Q,nS(?}Nc4HO	|7$/*n.U+d|==Ee)cvI"&>U	NztWS4IAMf>6y6eo'"fI)+D[PU0ac8q(m8Qg[?/\r9\HEYl7:2ThOwg#j B~3<55UqAdX9BQ1Ph7tOKr^Bb-nFuRY3o/Be,;VTzjsE+lv\-M|:<& NI0iHoIi8f	oz'Bn^O/KO<5wlx)xRV$EDJF{SWbb^3cEmTkn 
A?u%R6*c="3ZW"AZ0yN7D9cg?g\B[?S-|;HRdb`/'P~(W]z]/yT%yFC
T@)uBMa \a@XZ&"9e[^
^RMps`
4a+HB<qvd-/X]wgh6#)v)4s^yd[E/5d>
"S79DBLda7cY3Z65%047S,1OzEAPkj<)GjfO@vV$hQ9v5!*tq.)#hd^
Wn*ko!N{Om@{^xaa1/s#Pc?	|7.ZI0{jOsYt0i:#Fi=H2WY*HPsi?{$/'.f$]^F"r[>jNiJj"=`)I#/y S.xi	{lE-n}`?
7mS\*WWn6yJ/,A&0Re*IMK<H	r6!k;Sqbmjcjwl"EvK~d BJFp-/d~#;jhKVkJ^<omS9DI`A O|.xkiF5,V8X
Ynv&OF1+{,m$9)0{bS\F3'=\?V"8CphqNw_'QiOm=f1Zs^C{cts:ZZ$vt7Sk+%P[on`qeM(X] 5[P8,y#0sg	IUy	nB~(r:AWDo7taEUaa4Xo2/U9}Jbo.<gx=eg!DOW`gmPHgp^#u&`xm@QPvf,@5	0CO0J&TQPwH7'Pse[0HjEAvWl2/fu/*kgw?D-bGF-<P)[rr6B=K;^vyXf+*Y(ryovB,@l%oE	@CeVsaUQ1E%jg'-BFNHVx?gZ8!i2ZQ4`7!/XdpC|?n<ypR8">443
Yza:N\Gibw,!JQL,WXeE|x;!OKr
u;Xs5v}si
4v%1Ry&W_7W8|sdI!&l7W,Vej##vCht!J]Ww'(jsEB+4J}UNXO,*SBOt,3cmU;e/&}g_g+(t" kveR8Q4OE{D
]]k!ZC8aR `#3&+Vk:+"I[,=%@bJ#G") ]<h/)w'o$nlERr-F!!76`B7FCttnI
_Kk,
O%SF*Ai0zWiv^sAD>3'aDy2o
]sIIL#r?KXf;zh1-0@~3XZnlT6Jl7_(
c_E#5R[4QFkVf#%LUn;%zW;`j=Dq,$l3bm	Ahyx*37e'Mvw*S3wu6k	+SWvOG1p68-C<Anj+[?LK#D|nP
%U`U|@X]]^\?u<D8kBD9</:*vhK0Ei3BAU'K
>|?6T7
9V!RMiCk%.Ol~|]Fm\Hniv%2NT-l@[0Vvq|to,KgT5nOwqm>1ZKbml.02bhU3Ntf(sRws<u53S{-O8kNG^x6jcoahQ1?/jPvf<5BZr}C'!?Dg;F<'hl1{lCsvJ%RHx5-i&vDefY87sx/jnK)JljP;_vVeu!P{[G|\! MB$IDS?>gD5	w\WTgdCpetN)WF^4>[5oZaCiF0y)_\y9_&BaamJueF+\DId0-`FY8:}9Bv>F>3y$sdl8V.}}D
`3Q_72?F`I{KVUWc,DTqnypKzPZ#0X3zu\Js|!N`QydxXEk>,or:{1EckWn$aRi.eW'Um/p28K,Q[SZ_%s |>1ju&&ksWPzV]3,pZqRbAwg!FFmhbU3E'++4]:b\DKvyn6XP_*hI^PKDMFj3:C|-M		o$-`1m F!ofnJHj0$,aH1
OG$A3Q>Ql)S<wSBI{r9M}r<Jjo,J!V(Z&xxV:VwE/0U=(XtnI/IN
gN1)#(}sZ='<==/E%^HfwPY+zKU3PSX04D3H?"=%1!wT/ZJ)a,]JPn7td\]7h/>9>y	jrAZ#G2!x+qRqjKT5HO=RsyAbU!hQh	Z0,_1#ioldE8u\e$~`A%CdCu\l2SB-h1:LcXwd!zY1tOt|Vzw:W%v(XDf|,{.}Vg*
axJH,,}"vJ`T<+8y`wb9=4K`h
$4dI "h'/ygWwz>s?E$X2tB'Nj4M=|Rvbic^x02+}2esHBJVwrf\!#Cy}uLggPcF?yGah&^N*Y;`UMQ*[VNpRU'eG7_h0XuI3&?y^=HL*n#}3[^]xmOA:TKwaijV-99e+W/*W8t=2^q? M5j*m!2Yce;,)ykxlZQh(>E!f7J(ywPyZ.OM6@c1Uy}hEHk	|!*A7CR<U{c"):[A$$Csl?6Hgf4j9auQ@jev|wpf2GE#?F\,D]Nbhj.*GqEXkTb+vJ#\+Ncgz~],TK<&GNB8/3NED~{CR.5UF<rD4'FJ.^/M%,@|9Q3z#X[IKP7G4>0#=w):T='>NmBa{4(#~x0=2?>Cxk	I_8ip 1vVoHwfDyxbe4^<nsjMugi?&(O|J0]>#:,5o3@7E6fF-qUX<l{$D-l6^(^]b\1wlmqQcmhC(42?-i@^grUQ=;[6mI"VjO^+6noFB=,lg0-!$o pb]'KLRhA]g`JTqvb:uEAj14Mxe6=:h*)(Ip~z^N{b/T0ht_nHN[g+.{%(44nI}jJ}TB+uz*VF2:RDy!jf=:&1j7A$irm9g%_6L[L`(iD	29{DjRZGqI)t$X>69xWlFM$B
+0zZT5k-c@Z/x$o
HS/0DJGlMLaM30 7c.sP5Q]^6gHflB ;Z4pUB(Q^cPi:3%\(z[6+F$"4%G`:t5V{@RcSdN=
H_WM=@	^[S9g"Qmk"_9	rB[?V'a[*|OLoth''+Zb F?H{9fc7)N0C3K~?B\(UX!"z\H[1`K@,8	<;(=	R}E!*A,4<o,]^ht&}^u#+vvDpxJuO'_fmk	f1n;|tBbd\6|w~|H;Vjc7U)zU,w_/ypbHa0=+\z2i"NI{'VOh&z$'sE{nDXJuE(avd9z~Re\3AG{t3F'FTD	n6 nIA)d"DA^IOY@M!@I$J;_ULe",Hv)$8GGtXHUGjIa$w Q:"T	,,iV`U$\a7fS_-6Ft("o9$GYRPI6<r049;N}H@0Dg%A1pk%WJArEXE](x33'd2+2vd8WO,B5S1]xN$iu"YRms	q	])&s,6i19Yf(}MXi]FmeA ,.iD[>G~ 8NKU/W&].c]JprfjBWu*)^@(m! a`:!HiBObw1!n1]\&0B2Sm*Wj1E&#%H-OJX y\1i]Me|6(dJyL6]wCNG%]g1<ZmN|_U_sM"6]w+8e3m}-OU95US.%VcnghWT)q^f{^hzZ}P,vN;8wR\457	_v+%qc-*p[++pp<}/rv
OkA2J6_"#S@&!L@C/JFv	dAhH"3SZ`?T}nq[-\|:}a!L/f})"`%9B')u4y+g4eifQ%kG'-gb;LKN[*g+wq.^
<tcOM1;:__.Y5pS\.Ew*5fAb0_m4	"-x*"VKLSg%a01]zyXih'	[Ai3i84woPz"&#"@0:JT=$DN4s|Vkxs7)WmBDPCiqyh[
FQaB|!bex jaD%62~H)+c7pBMQ3Xe&	i -xF
YecJd%U4
AUAk\t_>,%+?dKgvi8"Qlplg|LYAe:3 vuSdQv [6	*gdq7%`@jhq>-OmD\rGq9A]k,wN-i|!aZ6l7MZrE&TI$(eWCVvhW_?J<9\bp9ibU3Px`8~WXw|?<FYFY1(V"ZDN:g4fmX&'`AE3]}fCX^ft}$C6Cjjj^swkUHctT/PE'P	9X7~]!`n%n6f/:uZ}0x[Z@HJ'581q;[22PsUl]PMzo_+	XWTzvim>'yl$S*C0]R'
#5P03%H_x;3^mRq|_Be2AL+fy/2C8."Zxl0sS+|Uz5,rPjn]3!WRo|~j)8]v]?"K/]hw?,LsqMc=6tpK:Qm	Zr&"E`|KdZ4|`fTy+ql$
i\g8T"RAH]E@[^tC%KIy-Gnjk9"IoVj]Y&10JU=um-:
JGq+!'),PGrlMs'6+dmUlo[;9x_P_5])W@^IrM|EY	&L
SbtN\1UF}'lYR9r6JfHNX6j<Ou>I&G0}Y|^(v
|9Oobq9vm
7d!8[0ESO((T\>  f/[)wb<Y_8"g;p[Iu[M]FFd_)AP_{zmgN})8C0],'&,j`We3O*<BT"knY0#i^=K`)^9Su4v/]a<pDM\>xkr
:Paay5%f=A.O/eO(L4LMdrJ.]gVYsyy{4B+=G7
Q9hEO#(iOc,L9&pkg5vU9zqV*=8e`Kv:g~E9JG[jN*T3;|WEm-]%1Rz[JA_0!s9g%J^S99EV=x,+vM,=dibFa@ Q[.6JuKW>~B{\X8:u^nas7t:hT[<\&zL2Jgl,F!ZN3Fhb^0k/)	S$&?]@_J={.GOe44k$t.cQXMo_M-K"E\p6>vrLa_Fx	:h.>L1JVM	S2 ,:FD1lbX &5/UxK6y7$dwoMr	cSZe'Vt]6{sD0:Y:c>#S4>Nvjsp?lQy1*Kqb0	jlg2%4i0%l0	]Zk\OCxfe2M7J~]:w2XX0'rsocM_hDafwzkfv$rtg}ozExg"_~N?(24"=9BGxJ,@\I.hKXkt)'CM7/4yZx7&;Dia?^Z_!%U9M11?k$Q!k.i1$z</^}
L4kn;0ZTn9H{8nuuS+Ei!qDB`x(flAZcHkhYdb	<A&/#L:]xKrz j=m]JQS|$Kr 8tn4660]du1;"S:K]Prv1'Rp)UC2exBd||{`Gc/8w6	[(S
	[GabfR*4QCd*;|r~f4#bk2bBsD4rR{u`{=1n,aC\h&KM^	eoBx":z%Qz1qunsNtiz.xx&0EU>\*fw;<`2DB8#NK*Zw#m].#n2G-YG.$'X;06p^v_\<eb{cYLVW#<>3^Kqu'FvYR:J_KWr}_Y.lpk0	J<8*9(l:"b9vIGFG.4XT&bhAg,P{K~.9~t1?*j2oWzj,R9}NEvr>e\\UD::WQeY<1WK#-L]a,n	t~0|3tu.d7R`iy6LAe.nUAcICCX4jZ(^#dIR!29Y{tc@e>7kT;pJeS[T<ga5{[{/z$@+2Ufj:.<elHZ-T~(p~]%b0.O8y+(c4"*Few&$zk.0xnBamy|c:Re+]F04xG }u]mxrO_bzcf	'[cG49+K~0_8C	a;l_C<p9;yn9)h5|CF@g3B,3L4Hy@pf}Ik9=VJCzf)TbpS'Xs
`	_CgZ$8xm\R-t|;~/<[%y''0o1k77Pt1kRYZz{EYSoMqawf#6!B`:) ?V1i8UtPiMrFTKGxjs\Ipy&p/%uc!+i6`{	/Ufj|(+EEJ2L7K`,$>m-M4V5ET`fzG=l%'wr7JFoGo19 Ea'YGCl3>:ie{d};Xl7$baU!wS`H\<j. 
8B	 3SpK9ERdW6M`%=Sl7&i"UE71:ECqts%c9:mN\}g:2!fmQIB{Eo3')c\r.;4mdNS0O(C0<"C8]^Febd6pzX1y`Ql^syT{d KHHW9>w:Arnx|3\qW>7vtKzM!P(M5v};b-^zlGl,y1^-$EHs+njeat#M{W7N0k;|I|M|$Q,mRnW5VW?Q<+Y+!q4t(P	^^LL?rOFn Bqsoa>qb}|LWyG:yjA5]*4XL_0>	6Hw*VzNvM|AZT6w'XO#b-Y:S$JnJWL?iA3:\*"iz]cqBLHqBg5SJrd90jx:%wjQ,PRw>sSf+w(aG -qiXy#e.}ik7_`P,VeM/lc:\S\SnADO1wN*d5R4I<q0c<Jq/=qJ"8ne,'IaZpr:p
2k|bF$b1cx-VO(@Rj!G?BC`Cw*U[>a;VKE`Mt[5d:V]wGjY\TDAw0Ob-	Z}$8|/MCC6"iUeJ49*f$bJhfwPKa`&6(AfNRh!m7H2}S2(oDk4p5%K}5Fec}DVos}@X$Xrs:7vN+$LNs\EK@}f_@<EI#>?yhjt>%t!t%=.o:}nd%%?U$E3UUA%6E&d<dw\.%>bDF8@T y@zp1a)&("EnM;uaofSK&pu$JM)W	;G#}D+p{hjWynwPWD^.&XM`\'-?eBSy$fa>B$O:GdEFsNI29bpK31E (7'0A:j,c$Q)Dnn#osrc;~eN,|C_J8t'B6%v=O#&iqS|f{x{u?DjNf6Y'f%WyvgDT6+uirIAU12o{3wkaI+OcHRFkWZh7VnwiF[lp-*b)rs<6T<k"Ml3TCm\1f|'2@A%Q::ChW(I*kl7tLJ8"W3t,B*0<'IHru4=YH1'}"j\hFS?;zjX> j@m=ofudlU<'/a}+dSmbSJ
7dm&*Y
XS4} d(n|z5\i}[i'7Y%)l.bLyf;UVlXnA_^$DbQmN1qe[.2 WOVw(\.+ycb#aa~x-j<~(' 	6Y9H^e2$H)TdCg!\nAm(iloTNLQ9n
TqAg%OUT_ae?}g]E/%o:$$=_Y`E#[u)?2ln)[;]CY&:G&`SlWp	;yd,?0J*}w7Y?t5 DIuDWvT*(#Aw-ac<^;b"?*:WPh8dI|Yhv!hEjb?\I/-;F	oR[y7DZRQo`N-Os	;!Sdx2NWL]\]wFn64+=ByW(HMPIfzcJ2N@yRwdU4c)`ifbo,MA(BN0tY!6n&.^P	*Yz<o'/=\:zZ^DB49j{vMj03f=<Df]g5T?kCUhxr[*?}?X!am;MPTp	n W^j2?^9lv4$@`h4o4!K tY|R3dSx/dvUU1va<wORDCigR)dw_2R2V
Q:I--2o8 2Qy4.rZt5y3bZ:X9n8p@p8US~=8_a] >=`q-{G-^v_R=2%M`$12'tY\<3omn ]3~4"M0e`O?UB)
8<o]$e)A?	%5{>_lg\6<T;KLECB*g\[L=>L/9=0SWSC2N5CPv&"uj='1d0zo{:lo$$e;Dz	Xn%2oo83[3FbM~,^N?=dx)mQKmxBF
9,@1c&_k~Uy7(0sH',*hc>NP97v*ZyjMNb7[sU@RR+s!*={9[Vkpc*j#B^g3fgf8Z9E019hk->#P5-A{E 'hNUjDs_i}Vv{~,~Ya'h8h}oYA<LYE4lI;0h_-KaPUS:5eb&yMI[m*"3dcNk#XQXRU
8NAp73a*tvUfs;*zPTe"
L][>s2Nqp>3S}z2>Z2O>%V%ng
uMW7mW[I_/*M{y/r`ekJN"2/!g\o_IueT)?i;l5>3]GN mi9VL,*138t4%jSK+>y&Jue<#J]!TZmKX8Q#Y6g~|.&UR?Q:.h],A7%t?,;-4M(UNwIqgvHJw;=FF'xYN9vq/UD)@hIyTVarHYihqf; Z U15_}]CZtC wbf238Wf+m<@J/1@2;f#yl5>a}nprGfh+^H?'3n[Ph\ex7T=P,l~qo0.B9rKcN/,{c1lUoeG^Hhb1Hb*EHHjccU47\ko.jOAF^C,neOk2}"rp%r]|>i(	ra
^R7vhFSWYH`LABx=@dZ#l>|7\O`:3jpV+m#b	j\Xjk6M%G	xyg\fw;4GKV_L&v((&1T;V@r~RtEo,ipQJm#zA"	3#30lZj0SXuJx0{N<bY;+HEM=F<f)q%>7[2e!.%@N1A&z_7*.&ZqkgyTd37p(Fc'Em	v"OYj=xk}3`euP}X`k!CGyc(5O9~p Bw42r"C.)Xg6W=<"`#eZ_%ZaGgclRbX4?,1'P"ZBs9qIx]n};>\m[nyHn!pwWeO$M@8/09E(HnHMq;{ ^L9`}\qdK$lY0KM`F\xFQ94	K:@<vV\,A,OQ+ 1b,iR>(;zL&:$0"kQBE[Cvgky@xn&4*qM")wSXWg]bWI$I*KmB.2/Pa-Lsvy	|zlZcbv=hJD-y@t6G1q!|Q-	;RCRXg4sd wf'XUd:_'{|'0)d6*M!Ee4DycQFmUgHy aKg-mKY|RRK`^h cnz>
;."8ov??jw|aN@0xB|,kI|^}IV9a;uM?D\0FvRDFt/gU.3#LArJ5=I^c7VS]{Ue_0}q14.AD|Ze81BBIR[cj@@%_kr/h^?1
?"^?dwj! SiST4nua$//[aF|0=.i\"V&<4A-vBq"{k|BSI	%jIq0E:.$p"TKN!%gF?`~qdGOb!1U]J791QBUx1aeBasC]M=aM8n*^
ajV2WCK_CsIL|toJn+&h3us1Gl?3NZUy&)7'uCp$~&\HpXv<NFY7WEgsIBcsru>d4rY
c`sd<e7\[f+@8yuUPxDK;0_xID=tG5sZ9H$gnL5't!|DD%.&HpsA49o)Ei_9rEjneE/4|gLJ{O91vO8=%4j5m<|B&i!5sm{,1FK7!</t,HuyOr?G#mx_**dpqsY`^?woHs>mI1|Cg4`qnSz*=S4q0}Cz^!@lh2"?C$lESt?tf$,{z3xZ,
U7nUVD}W&C[p=P;*ARK56(G	~c>]_M[WSO<_-IT,^{s"o1m'2DN":l>sbZ75P]M@*	u?UE=JO^vM4w.fB09;Qw]i
x2a{FU{"B6~$;bg}H)up7
):b51Si|*ss#!ZDT#pw&u4QVe/M<6uf*?1!nGD&"b|jK=7iuRKr{8"c0$3F=<R'#N$ALFS^<\jlU0QIL/t,WN=/N Jep."])/LRu(]\n[QK{7`SG>r.BCi OH7FkPNM}*hu<L&S?I9x^-Vb.EBQ%*JF f.GAaP
JJ$XTEr|by?)RzwT+0Pm	lBqXHGG w
>/HKKmXUrOWiu^3sYM"	**;=l>C4d,mZb+hX8FD^:4yHm9,q$R/u2\y#TS k0X]Y +mT&r__y;Ts"D&MwK`|A=%8+0'N\+Wop:XH|3
uFR"616N,~+PR	>*wIuPu^C'p
7h8hv>&A$6TaUQ6]GX&.Bq)5"z-vj~.Gu]a:(>ipDN1)?rV"9#Y/8Js8>l52~Zp:'Y,kn=wnw&'$y*&\Mpj,ZE3	umC6".eh84Y7$Yg5-*1;%R|/	q?@c`Y\A!
9;wp8wY`12\:A%D-2n=T4_Rxji)8$"Rdsyy2{\fpD?Va9wb^Qu_{_nqnu!}G"@_:VE]C}I^']v>$
L5eFL #I`HLZ`m.9\({D[npd4;nNEQhiBx
Q\,UFa8z
:mXgsJaEhDV"JSvW{/OU"wp]@$h(jK|qF_oyX/7[YyZd-2F2m8@&sn1TkT]HkH8Vd/*bI},8M;i*=vCY}(1K\nl)2op@b"M1^Zw}3hJ\{Z@2pxIB/ow\Au?n"myE0BJlM}sOF]P4&"(v`V[Mx'/S|!_9#iYl@|o|g\5}4ix]Eri>weR-'^b5oLw[mG#c;Jt7V#	}W%tml>'g(L8.y?-y-uQPt(UG|HcN^v{fb&(&6K945+H	q%>Dg;6`-y$BIJF]m1He&'L)$n?%c}r	T4"w|#yH#W@O%S<DLvE4B{x<#KJpfQ@"nH1fn!r8;M~XiO\oVB:mZ'z~Y.'t~G}\M +']4Og&_49i04d^tp
7#0rmy0*|v,%Sd\Mhx`0G'4o&Dd>i)52H3Rz;b;R]<J>0U:0/=d(bw0o15u#'eZ`R%fK56b&R%H.Z`dEwY;|F.L=?=]BZ=1)iv:l%t{=b6S
	_rCjC/B:Xc/5zU$=-X6p+<aJ"_Hf
06(hHs^RUptZoXOtFuZ,_9DUU38>lg	=6Gn	|e4zX>ALO'}9mL?lzzc)9Y4+	QXjz@XmFbM(j0_Y&M$^;IC=*7kBl(~@=|t-P0O*P1L-lZV:vy>^V_[riper|1;u,aI)Xg<1)6.6)74Nui'Ix~
vvvVTKw-_orQ1y9)aC MI~K&dKj&\2u&d2'[d+ 5A+T~h]x3*j@f$g1jkFGMsQs-hzA5C((([Pq5b3*S+q"tY0:FFLf'Ut"Vu3j*y.O+[jwMFgn:Kiv=Dcql27q@pEHMgPHOH$;EUDf[QMTbx8glcKr*7^eBf"6OO
D%l$dd`Rc7W!"!vW:roTyz(ek -b^W>e}&$fYO1bE=%5I9VA<u7X*(dP^|88,Ca;@04`c4Y-A7019Q9P[!dQ9L>tIL$8"4lZ46myG02*ypu(oXI0$a7_QRY@:kFzr)^(vd5b5.k07E}
zo`1OWTpBM?`pPo8$#c\iN>"-,i8V2'Tbu8LKKlj0im&y)F3;N2B:vQE:EaE/0N$>dHil{u":c*g/Xl9;(10B6Eq7G'P'Vg`^{`s4iGiEC5c$"I$155P\d	d|w PoT@@g1?{::,	z^c82D,'y7)'Tt'u@5w.m.Alf{YNp'=06#.vm,aZ$?w>9m <l%zy_(5D6}5d
f	"v
aal_X88oGmCY'wSZ|mqs6RZ3~U3nUoPzxJK
_8`pEs#8b'dcD1:NR*o?qaTu~&d+ID#tB,L|A*GRU9	_8"jRR=$5`yWg@x913A}_HL]r/\<volm3tPntY_YTdQ8r/^sdX. Bqdgb19W$K4Xy]=[c J4|0xew6z9T|LC*Lo[%	#+wQD?;GcV!@.sHWU&Ul8AT#\GmJ`QNz0Wy5VFt<fi=Lt2n|.5]y#g<In`MP916<NsG8)gKs4=$0>9lNw0PSQ2uj{+3v"]'@QVpg&	eT~E!N*[{*}ujv$Q,PKq+#S@>QF\1U3!#HnP-*yf\*ij?5v4m<=B+wN%[B"%Q|wO8KXPSEZy}pzk2A{"Uikdo6?zT}^^gndps.hB/HC0
}]mZ,!ly#o6".t/xt-#33(,bL3]9`;VBK*Q6~[x>G/ynb"51ot_M5xyzd&wD-@9
pFH_8*jc;.B@=+9>)J[FW`sJ@o
jYA=hV;}b@)_?S0$fKXa"W+pJ%U)^a^b#!/J2$X4NRA(4?!0UFNu~US_+ya"&`Y
0MRx?=fYM|<{8s_2H3z]~mp;!	%	CGj4NUosilMD!P(WC0~	zx
.XZm>36b>rf\xf?9m	lPkGH gxiS!Bs3BO:^rM[pISW'`$GQ#5Na;s8IOEVn$vl6fYEb]Vw)W?}=GXE-j"#m?+pl>o&BvBCVGO!~tO(f39CK?Yl*:qcY\d*)@
=o%0~4$~XRRLCZQ~|hjT3t3(C[ .K:;Pro:/*yP6m'[k]Gm#.UA;6dB[|+v7'_ydH3&0b
prowL

O"LXqKh>"}KJ>9sXLQvzOWx$9pA?,GMwH[TyGw//X:E3\>C8h$6*!i|ZF>"<kvI(.zze*Qb-+
"Q

58[U{@.Z/ dhTgsK@^of\IIA>=`fPhDP8cxz*3Pl,wfGNFS0g=,!;$?|/Prky5Ds1N0OWGS$8AVv,X}Mw]-9;^"zCApGw_64/D$
;qn9L&gv=Xx1+Z(A1~B6o-kF#[(gl`Q0hrnT#-,[_R)~.i b4B75[;RbMlFB,k@N|(<RA]7|ci&'RU&JgA6@`FD)VdR92TI]`N\jA=UXO\><f-3LTFHyj1(o_'/Z=z#Ezf2\H9;C0e?]!1o' %
r\b!unq3~F+DdvZW/|5kA3[HL|zuiQdLd:l_~@,Y,A9abRi4XD1.O.>Ppct*.~rlG&'L&'9Uirqp=M>tx2;]i/QW$8lV+	Hw.Fn*_
=	Ov[Q*1%RTXAz6p2~+>~nEak*zcH
5@"dM
Js>x3Yl=l!9;j#duY-A4n>)O:n3^DH%Q}8<pfZ/;7)&I-AYYWSHH0~zWDrU1vkHOh8[[EIY*?<"_zOCONq<fWdt],f Qz]1)`UQycJ*cv/=btv==X(Ge$uNbZLCsBt+9aT|N:
.Ndw{z{Ehm,w5*8c[Q(+	a=^6|jar	v?`6A*fn0JGU--|hKY	
qdZoed))+u^6/ aF${0o/>ebK	/g%y
5\`mRr$!p0pq&e.c9dLr{o'nyKI'JT	Nm_uyW vv+o	B4k'J+pCL*^^!en9{VvX5.ht0BEqU^{kDM;sPQ.0`9H!v[SK}]YP7=k,`cO@3o^@'X3!SCf#hPxz&!r>xRULH(gNxh 85TuW8qE%!`U%u0g	y<6sefmDAQf?5abWou^B75@;qjlny7Ws(!9mxcRAC)vlm@i[N2a@}QDny&+ $4OzsP7Fw3I(}]Z%cGfU-_fCgI+IM fCG2^5tU-5k0we+M+jtw5N,1++7G@S hg9G
f)k!3<>@^-x)']%uX4k4mg.
wNx!v38md;I8jHq0^| !r7\Jr kA><`8/lA^&`;E'C"HH{!3PDdcW%BU#FH)l=pJ$PmH8yw<2dvw^i|K,)}BB!L#5wds|5_^Sjmix.xx\sJu1N94_|-C'TEEsy'miCR[oX;MP52+pWwOuEQA ZS;pvn)j{Gegu.^I4k4-UC_	1 ?Lvf-_Hg'}H_u*Ww	]?U]bt5~Dx3gmF"_*y}+{*;z`gE4xi:qqe!r c)m+EJ:#W5vogde;bnq,QC&XJ{Fi;5}e&;Li.+.!JN)mQezg5#C@^k&(^M,1-Z;)CW[x3du?$9bLd]KEb`O&Vk5'l|'78;r$J5g{3'hT:I-l9LBk[m6,Kr.Fd&tbm`[{QcZ_O<^Yf]((Feo9-A4UBjHS}o0x?vOJdQ|"<R9^nMrZ1SO/]w-7_2RNq(2(
OVv@-mjs+Ts$h?.5IlmRjsfHf_g[?D!WYFFNb_2h$X$hFAQ#y:~4o'bm8RU4ps6QqzGCcdY2]wfT8g
h*\U,CDz*"0>{x(TD36*O)iA=FRn2$WB&blx^^Io"1ff4M]OCq>v7<V9aGJC^h=u	|SvLXb)eO=sc15w\GU:Cm.<|0+u\Q5[,Dsc({z;n\Qz-
N@`e>dCb;voo{t?R`!"ns^
~"%Go$YZG]kkoJo;?9DF5B7K.U!G,t'*Dg%1a;$bofFj!bebfmWn,=EG>Ha_BSguT2;.r>ok7"j?YL_G@$I*:BJ)Z EZ8?57D`Qv~s:Dg_`8#R]
BzQk8wJg_QU|$Bh>B6	[puAu\lc>WZ
j.;;Zv(uLCZwazVjp!{6|6h3Y; >7s{_\q,sfY2R%G>%q3P5(XKqO(Zb9mwsn6/k;GQG;15M%IH(r^`N0z4fI"-K)B+t'!FF1hvb3-YH8I4uy!-y{!*r_xWaG'
**j{(t__ftL5CiwPud9ctR(f ;ylN?y\$tbyv:vU]YPSmY %:f#nXva&Uz lkcA<)#{Lf?o5vG$x;V2iAUeZlHsj)n8}Ax6}RQmMi9,L,hkU{J(Wk#p}Nr4pX -AKt6P ?w,d }N0V*M*.)Mu>;[Lq[X7G!g %<u@3jv!I[@_`U4xJ$1y[n3k/CJ'[?5T(;t@M[PZ18phv_S?PF!bg\qyJ^sVu~#ApRH@>a1j.8E^=h@	dG3:8IxgxoKQs,) M6)>GQsVU_|X^f@I@x~5 6A`()hE~98L{?Z$~$uuqW/Dkbl{SLc]7_%,&%opY+{1+5|McM7ypDB1fxqnu~N>:8s)JOD:CIaJguT30a+G\+[Z(AA2xrCfs+YXJv5uE=Tu>cz7<"?/O='GeoEl9P?t<6?T
z^[??Xp4<
PP-'<jRt0aKnw!.b-cJIp\*+3W(}hZ@Cx5l+.$$dm$X~qg5">VYGU;_3H8	3\^J}*4fZ(]"K/Qi459@N1d>ph&7hFvV%yFTJnW!eVH5T)k7F>.DA]F]),d#ZhkqP=PeyTvM5=UQv-wv?s^hJ("K,'YQ'5A)C:)uuEFo.yxZM"PL1T7Wd':D9B `)P	jEB}#Lt?7pt8[u_ve?/ZLboAD$>}H[u73V"@(=n\LNgA`XLoFLYs&.-\S&wD Nh!IOj$dzCf1Lfmk7j#<	Tl_Y/-s`
7lx	PJjyFR3t|,9"AMG{>SpGb{wZn./o7#6:FxpVDQ8R4)hHN;8>*3dqt),l,,1`2$KSwC*x_Z:r\q
({wEFR^a>M07Pqn~fHoRWc	
MJlsdCPTn36=tR:_>0NHa'Hu$M0V@uqNYQ3 H;.R',VptJ.f<K]D+22o?|8T\X*@S'146jZa qtT'}c)J*rl<V* @H]6ogES*HPcKYn%+YbUcyfo :.iRj:=tW4sr5!8i
"qD@zF0K\d\DsXI47Xt8NHtB*8-[JblMD"k4,DQ9#q2}gnA^uuQe%.k
:y0j#Wj.SdY/0_RNDBT@Lz,J,'%55	,~$nM3TCZ'5AQ5fslT r/SnKi0"=N'kNt
e<8"T!t7
Sy-k_V|s"#7teXvI"`higCe L|A5IUdtNeXA|V22L3pUF$j/DM7|"f8{;WoJd:.^$2cf-|!L1@;`3`yKp/T#	>*(r#sApBP{V<frB?k'sF!
1={U'Hv_<Ws?gX'>:$&.n.+2H]{!	m0N3Qj.VPS$3MhC9K	rVer3yIA.@=}*[Kb+. BB6ak)D^}oc~&P]M$n^?=q%;-w_L5/#U}t$'Fk/P&&z`R-(K=zgIO]Uwu*FAXbeI<6WK"Rm}7
V,4`RChO	 :ENR>UO(cVxJaF-if/7wCE_d6S@*CdI,oKq+N$xUgq%vCeA]7(vw/i Tqms%9_?0/{|	"\6XC3mlV[#FI)o$Fbv4c8N!]u#l}VdP@H<3W=m-{w{<CX>3+G(X"q9FL\/%
pqsdp[IvrvH_ISh@Qf#q2XTo;oa{J0Q{1T+gs 3HrgU:Dm)Fr=etrIg@[26 Etxe36Zb^+kr-- \q?/Fa7K8ZU*V4q/[jvAG\l\R-spZbN`-GV@khHh\m(|q./,4T4x
xW=64kN]q]*8yB%{$&e.a?ldHVPSFo41-#a)qe3TbE/o (Y%s\8>6y
b.NE6Rc|>lJCgtZK6`.<RvlWM$mo_]R[ux&(=x) gF
OY}L^Y=1T>XrQ?	%|	(.INA7w+5~U+]h4R!D7J{lOHo$f_ #MWb=O\&B_?z/UMPIr9&6[t
aBp,al5G(Mk	#$uV$OF)0ALGl<W^&"<l4"\{B01;
{oQ+!MF$iK<6'
z\F!{#OeCVb	QB?L0f!C:/qAa-)iXs^V^vlx_F-<7\OA1Q"K~IH](P'a.gQc#.HF[[OY<+
:$U/M4&uh>~^nMT{**P_Qys%d+UGoS..r*c4W@:iWCV9s`S)9L1,2VO.W,`B%"6[k;'~wj[F)JE|>Px!<:0YhHrdemhq
XF<xOmMP<t}Oo*fS'o	dE'w1Ux_wXPQF8LSy{Ol5wjm`-IsYumh-iX!:w~+8S\b,{1qJxeQn6`RhF%7x/d6)M>W[i6
hM5wXtH%Mx^XU{B|16EE+z>' R}V@7o}R_1/9eTyS!]1.3M%&%uzJYY]%*G[> dfYcoC9j}LL+u;;;_.
{n#AS2k/x8Wcvt49\#6]t%+[	J&Vn-omDp`XzkVtgmrHnXCBKv%%K-UKM1Mdx5|6/=`"fq$siv1"HvYR84<^^]"0T8+K<(ZdMmH)0~Jh1.aG-{>~n
0{yBn|`3}Itv_[kjq|}lu@3`	|1a<'E<Zqdu%WPFbaYxMxdm]5,i:+<-UkSq!(pD.NnbND-vN
<l~{wS]
uk93IoT;\%_<Sb^q4ypA$xOPny-d)
qTrAHe3kP(Gj$L0cFCF|v''`KT?MSlj2JOGr,!I:JM9aWQpDPxD"`|@yX7Gh\r$D*HVqb'GKiAN"%92C}~Axwx2<^1v6u	}Ks'#{
x(37:%5gAcW&ePqnc+oX8C$h'b7o~RjHt4*Nn4L~O=.h{z1-2GYJv*nE|2E)2A<(yDm&iQ,I:,-mL{"<pDs>(%\t[;'Ja~ru%Fi~qxFh8!4fAI+-|?>\H^XT<ev`viXn$|aQg#	I4s=l
"j1]seh`.'-*SdrpT+56rHsFw%2%f.Rk).6y1.Fv`ro'+/*ICxm$A,E+zmR,K!CM_ i/.rv_OO1k+g_B5/PJ1;X{lfr)zu-\Ri.uj4O5J*m&Y%D)w9V{7[J`|l6ZP1FAJUCo=ae+Kq0" .8"^8|0~7k/!d*#;Lhx`F*0mA%?JigB8nMU:2oc;=%=Tg)'9M)?7W*\]0wF>#+en}|`@QfcdtCd0'
5?jD_<PQj,k	X*xo[r_A(lkG"i8}a~:|3^(X.ieMJC	[u+"rJ/$}]o v-x@?sA$:@e:B_$Glyh"$kYtn9GdL#TGEG@*-+?	+Z/1g~e[I\	)Hi	B`4*DYep+i@Q/I@v?bre!Hg	!LH^
! 8b}~>nGb]ozgjbGck5V%)i;}1)OPIp-a|066W	l<$2R)+-vh.38}OZn[h-U,kAXh
ZR]U2C\[!?xr3Y*{#AH|+ZZxy`v51>c5)bj]>4Ji\tW/DqFkJO>*SZqDaK)snsT7
Sr/#X$X2_\21F)}+pV.xCTxDkHwEyoIL,v/`.<7RBSw;c-lprl%Bss%5
XJ)Ce5s[{>Z:eJo\"]m.izOa.LEC421<lh4:YCNlz&[w3M4k5]@N3y4*/|&A#O{LC,W0G?.GC;Poo2P44^cuO/HX~8Q5gOg~#P3AF_2jIcBc'Qcb%DPK<i9?H0_/J/$xp0dJ'E>|(#op.=epa!sZ!3GV6`H%>~NxTl_6[@I6t^9>-f_f3kafGf'a)  {>A0LF.g}`X4SqhHAZ)H#]4~h*g:JlUvS\7J.	9ni.k#| B|Surg<_Ts8T% 
&G^&{Lag
QD
xY9ae+mZen{FQSA^<
lQ}_ja.vtk=-v:Z'B-q LN&Cb.,bMS<9aW~}B^E3g`d\LE0J]_.4f?9&j?e>aL5/LF
uSPSR0qI$wrR-oMsf@@<E$:l1/+GvG&k^i#),<&w68v?WjzMx:VD=6c*:zn>CCk$kIx#V[9WE%9/':eu}{	`LTI	nX7;mM1'&a4" Z+u	*<fG{@scF_k(53kN:P5`_"ZCyil &.X;x?	F(cKf;[QMByyW9x__tHFu,Kua~C~ZxF\ml8VvK&rW}rvxk"zu&eI)*^aW|+>&A]QaO/B[0*5$gIK5UTyiq7%4f!=q%bMI&zpkkNkSglH[#=6ww^k[fh|q
j*^) `NG!&8i^xLx]32nOgR?4XGvi AyziF;hr$$l.#XR]2mU.1a)^D*_H'Zn$9icuj>oAe|@9@U%vidmD:kW4b{t})u|wU?!Iih'cn) uJJL)sL\N0$@@R1W<_$(M[/~/Db,O2M!$edS15
CCS&$\WI5b=i,?;jM1d!n&X\=*qzPmV@;Q|?sfNK5;OQ_4:)Vn(lLPneWL_36U=NfXD$"PE	CVga<jv1$_9Q=@Uko6wuS+XJD$'lEa_Vw"	aI;D4{8wi=?tfln3l3eQ
=Ys}0F`jnlj?dcJbG^-}<gG+e:![l?Id0es[Y"NdK:n/;ag9Dm=K:JVyO$Yyzdulq$s@$`|4>T*^-Iv1cSG>04nT2dDHzFm.nF\.Cy+)Hr\1u"57T]2VDfT93S/-ZNy[A@I}jyESBSuGHW7fK=f4Upl"qK9tP-AcZMrzIlu"o,	z;VqEMwGybe9ai+570vuQ(C[wA9uhUGut_Uu5]Dk5?SnAZ>]]y7T/%1a.}x.3|?Wo=EY'koDhhiVSu:pio1}9{
e|k8&^|ct@s0[Sy"(),Cr+:
:Asl3dUt#)Dj
|F=1:yV,u,v\+$;= g8G(Ag5rK`(DAV:]-e~+W`haoUQ#wgw [.+RfSo	roI;S9,T6#h+h6.:!nLTRI9W}]5cvW2Dai%yq.r!\X[?}rIqMk-7(Q[r=fmiSS{@]V`%S\md`jP8Q@;$(#j)?R@+SoFgp6@T|gW&x=:jjv{bPD; !P-PE^b)&]'(7B |2[}[9ES|S){G;M{673;%Qz5}d
|nI,9S]-&z!9[;{hq8YND-`iI&4}czH)5Ob6NN1e%MjAVn%m=2F*}y{u{2VZUK/=g@LVoXI9B
`#yGRF[jTdBqYQuMW9SzT+`^Ip[ny,]KDS!9|)Lx|I^!sOAA04M5	~/[;(\$v3%d*oIvR:3yF6l!WW wq#/0> xkr<4+7'EFRw6{Ms)+zI.:BE[L6A&Zt~pKq|QO3{S?ms\Lt!~EAYpc~_UGA60J]/ta(=Fz$M0@o]32
9D	[W=rJKU<@P?]to^L{.vwv)BV4hg?hH=rl7kJy7K*|liw?<54}ex:[G!2n*!4ZW%C+V[IzpAWxKw19O`V3NX{u'AYdgxp>b^#+zQqi7!zLA}p'H)^"KwkYfNId1,MoXp.^.De/<WQ`Gycs[}#Ped)2Cwi>oOL5nuGAK&6PoC73'2?nkw!Y26Uf*V Y#n
[U;d~ss>&@4I.152a-\TW3,`{VQ&]Ia;6Nf!42TI^9$tvN~3S_	0C,/YNQb}qB#pz{=hd1__n6e5l?%po\6{&%a2&q.hxeNxb|Ow)6QLa'{;%dl"z8H1{(,sD-ky]+g_TqUg#CopIgTh0W@m|/V9q06]PB`*1BkBDJ:B%"%vdCj9eLT	~FyD- ^P)3|a1B3/|7MBt(*9/5{|%zoEaIb Rf\FAK:rB-Xnc6h2vbm9OI&03G67`MJt^}ttO\Q;aVk"x'GFp%ZrB(==lZ{/|&:YPshu'5CemDtXn-^y>!"DUh.G0.,Km]~C#'.\4m{' Io'@MBn=o@LFEC#)uY!8@#J'*i]O\\;y1Sg	cG@p!)5:6pJK=_I[rsTRbQ9}!^Kx-VFJ&##R*)hf?8Yp3w1o?,lcb 1;d[IE\39h9A~fj"3kb=oxLKt2gj,`BMF.kCGEJ"j"3Nbr{&qee:7l|%sE91*B^l4/HM)%rZK@whi&NF~IHLCDOZ6AF"*1=e}Z(M?4r%(Gn!7oq2	$Y$n&zD	`%u<[#-7.QKBP51%wZ<4Uus+l<7Apic+ <s@_$`
-A:
~{i!]:lN	i]ThvBuN`h.;J}Fv4@#yQ9\QhhZ?.qTodF)pIv7{?DHh Y#O=Vy=e(};eUy4pd*vM5{=12V($YL1s?h@rD^fDIR)P"#RYFWh/@DT +C-U\X~tn|#1m*g68p[|Ll{<<vt,[|6YP7)utl
FLXl
C}pf!c-kG2"=G~
\RJ[;WdnSHl&_kuQIo	ziVi4N5#3E,H6nkf9N]H}DRi$`SJq--cn;XgO[5|C%P>3WpLtz) HrWY}kiQNdIQ$$gK|x9i=nrv3pkEYkY=*6C?QxZF.Z#rbkne>fdr["INdQW	8 xW9[s4
L10[\(b1;;='*S[	JtFv.s_/:j6Zws
A); 'W"7Ye-p{6Jv{dr/x;-3f.<]E o|#V U\$[/hN27#=%mr.e=qnb)CiNj8a+JLaKE [vDo'#97rFYEYi@iq&S_VlkL
e^rQ c2&L3`vm9XS:jg$E@n{38`VY$k;8jD1mKvgd-wSeT<=~ylli$T5ws<qbpi%N)z{"O+c4;	DYV82vw{9ASk$I9%7YFchX0{-`-yQTGV3C^T!(SHLYb+-("O\EC`DB?]]dxM8crK%,eMqn1q#0 .;G+l"M9F+K&O95RT5IOvyLr<RC=S0@|A:kDNp_!iVm
L$8%d|Se,Wv@(@v^#M#Z/k$Iw|?qZBF.}y~~^UzZ@'+JgOt{	GVNd`8e]DD&^]@Uncpb+f|K^,f4@Vj{T%QE+A>AJ,[c,Q@|fCY~PU"3^NZvJ.r')|A-y^M{>=Z{ &#]w6W<u>_kENA%(mxiMBII&<+=b8RzC9G*N)}QwB/:}_hpA}I$-bh1#"RlL|~{XZb{qBzQ5`!Q]`	u_jj^?7hX-5dilG03Anb)b:m$9P31id=?+:;7wSF;s`qgFa-$I]+wqk%?^ujYE'h4HnooXZ2>}ZA)CdN]F0r
p4Qef5-hYJL1]8=#@.zm_K1DR=vXP !0_<	dX e&W`[!jenegAE[MKyiT.apfo.iMo_9zi-$6`Ld\vw:pT~DkS!nr^FZ
!Q]gM
|fme(akRFL1=v)Vif&S_x}->ZuxRxr-|0eu.ldPH|KFWf+9X|/71)ca.fi]qoBzTJVBY~x[Ds@t>tlrx"_Lt[uvF,PC\TIko5r/lz=Y i\(nZ#kx-1x%KVFO]r'`pX"cZ&*jwC@Go=>x#WrI93Pj3P"6~M'Q[7*sX
,xi&/bK'}N<I3<A>Ud|M,T#Y <k'8w)xLX=!dOd#YV e0fwDG&KT#
>1x*stGv0<qFONe)@Ef{KaRCW7Zd`OLjYUf&|<4d{X'*4gK~|\fhRa4ABiS .8KBRZ5LnM=::$i&?}LTl;sE+	h#O=},HBX	-]fi<
]n,S8||3ta1XCX_Z'` *Lt`Ci#EZ[e9)l[HTWXo+??
L~4FPe@9t=zm&{Rz(MEp{F=eK>%X'1|d@pPt^<|?Nsr$O)bH!q\C=)~Ik%7FC@T1c	7DRVm6b^W&1~= ZYcu"*S}e\C7gM<m6X|J7%#cfJi0<i	W@cC%F_}'''#uMH/_cKI-/#4^b3dgvm5)?d$;	) bB6j4'QWbl{lvni#6(ME4]w;Sin<8a}[4R]7P5E(w!Dbsbd<+[FXFZ?R7Qx0+Fz58\g097I;dp99(RJX9"!W6Sr$~^0{Lz[kBx87"b n/	q;SIIBQ#>c+2<7@cx,xd>B3/TX5BWGx< Sd)/;0I};`U|iG2Quz@S{;%g)_9$|31=.G.<_"`1kXQl\^J0R8]Y}``72h4$3&}5Zg)Z!nX1bNsq+FetqPGPbHFTp9_,nL-`#<YtxZz$K2oWKd596dl]'Hx#O(!|Nsd{28Y5"y.3FZ^+KQ
a'%
Bq.D2F)1S:Tq>&U2Ex*c%1E(($jp!!UJ)R;{y:=cA5EQnTJGJtw!?tlAdjij:n6p
WvI+2|=c4}rd'$JeS9}50|_{_{
vW.&
q*D<
83ahvj0fi*?N{P'wm`0cIyS)A_<Grb76/ey^"M$cPc./NWh&Co${Gz-Y&yW\,&M}DE"	)aPzFQC)\TWh[^iIQHOW'./C#ZA)y%,eLI%/F!E@@Df8=x_?l7PNE#=akM62\P21\^0~#-N%WaP5,1	SJMfz?kO]tfFUzVy*>DC|[@{Afm!XXoa|{/'Q`2pE:\i8e
y(:4x`KYc~74dJgGL}d"@+|u?z;\`L14l?CdNK(t)C2TD)9_:Rt}qStI8W30<JQKXdBH4l]w.uZr5hN_sO,}u_Lv^5WSILC,hUg.Mrd3LPrcA0Khb=::%FQqVo[ZH@iFVRvTR2OH.(:5ze)7NTPR}ld}s*/!gQxIyC^"ey9d*2OPg|mUMET#KI98?RHEHhb[FG ./WNacc,ztj*^i(;0\.2X'a?NiRTK[uu*=f/&U*[T3V:^Hu :*`rylg/j4R?MLn.
	QS/1Inl/w3-	kgcLc3L.H(f'R#) >xq`=f$&rSED:dVd!@"mt*Hx/,vZP5F.Mfh`f6KN	$FJ903>hG4oCP8)k+%MrV!yo%<
=<76
TQ-)>w&)X.,T	@?A5X_UXD	w*qQ-z1Q	FAC?]*kUOx wC(_Xzf|]TH1/X
z{7v|@aQHSk.Rk87f/=g{_i9R2c>A3tBvq*M%'^n!sEg`p4M'FJVkpVm
B>+}(K!,FYuO?96)Bbiu82Whe'e@3)Qywb
@z	P0QDFx>H$-Q+D.A."rvp6VbxbMH(#	sBMU:"A<O,10RCzAS.>	Ol-h	x{2W*!IuDiN,X/R* M4x1mVY(9F5E$u@=^:7
<liUSssmhAVgv7]-4h$s*1`B^4Lm8	>jMk|iJFmQ!x/3\D7~J<OMP*`.UWg(K6OYi9y0wc
UX+kneDL6&a65Bx:@[qy 'dB :QcVx/XxjFd!G6k]Su2tY+I
+tivQ8}oPV+S_@XqUw.^csy	'Ya|$T}g2g#hn*raAvahIw$%xRv:r8c_(,AXh@}k{J$%D[i4;[\Hb$+<:_?-e'%{u;*fb}+HUZHs,]qWOA0zb4U%u3ZbxcU/DmW&m$Qm^xJx|N^EB7.n
(~u[Z|G:*(mSwD Mz-Wkp>]!Q1Yi!TDAG-hxas%%|XS;w0+5e8_Sh=;Omv:n8U0u0&fJr?{)nC=:hqqg/S5S8:!8T=v3F~GIp|bb@P'{'L]^Q(/$u75Td$z27;M[qTvs"rzrg$Sm{l-kv=`zyQQ!69LEZuB.L5{@a\%}ocjk8a>L?VNB7)	_o'"6IZU4"GfUPA8>S%8EP:-HYz4Zfp//E&]y^FxMu~~JwFsqOsL;U7Z@x-	5v`!_1ZvQ8ISXOdf9"mF4u(hVvOjs 3;NqJq+(5>`r*mWU!NuXMi^PI=Ozo|YaLM_@V/x/r8#0ZQM
n_D:ub-Y7CqFR8Fu,q'`3eX*iEv{j-,"Jv|EM>{SEJ)FtEj)iC.:p]Q>F!*u1D7tN5MfQvDdBN^Iq#|&3u9fQ]oU<|7khXt2cwUK3Mn&/M`3y&A-
|Y:"4S8/Rd[1ex)3wqA)o5hH^c6q)<xg@2-"`Gs`
QLFB;G<	A
sjr#)zosIbBJQk_JxaS$dv([;huL)h-n*}lL4K8MHA^k8ko<HVk4n0x_:J(w
j)2Y5UE_LWZzT7^ouB&yI[C&5?	2hdK~5]!FSg`<x=<QDook(/N+^7\@5i<N@OW0o	{Qmq8x4"r8wbS*o|g_xdo*Rz|vcr-f(%DXjy22hPm^] WN\u8!WB*KE!QRYr |?D?cr]ESrcEy\v[G<r]l96C	
Fi!'?s_v
`bQEgU/Pn[bV\s68"d|.-C#K?[Ajg~`nQ-0_)S}UDXs=~1.T4fW46i1d,Ux*,?(=!>uG\<$8=pW^imL;,|z&;5l=RUJ=*|.L?P
 x}[lO:=FF7ZWb7@Cp\}-]dy7]'.OJ-8Q&`wq]Hu5UWAF(Ne{
LwSz{fhF:Gg4QyRz$2?ydyRF7Cp]f<lH~zbszW([@Q*c0tY9ki=0n~J3|!x9Zpwl:kpGta;4KXD7hlFwwI^@mvtj_0Q%d~9mkR0T*U_ifiD I{^_ozh=I+;`#F^ffOWhOL|^xd(oK \_ Qr\nOyT&C+ifdBh!cb1MC,^/UVD4Y"y1:xLJL`N q\77X:O7Z 5swSZ]x)a0!ImN,h-J=gOmL7nym6X"V_P00*vg]RA4)odf@v?0NNamwVvG+7T7opvs[0L#U*PH?7CwFBbA>`lVbMA YbQ,[A^d"u;o$W{{~vB3*S6NLpTGm<3fau#M7yha9y E3Y GA]xA44,uj=v(]h6b	50Y/\;Rkbs}ZH{Y#ll:xzVo"N)dW+oykDi-rVgQqOt2W@R%=llMsp8NF1QkAy<b~bVXBe+sgSG]UEE}+?@#>^=z8H_q_I>.3[+M+0	M
'`6P<DIsI0p|5VB#xz@C'?'rN
@N:^RF}|gF.[(S M##zC-!jdbtV*=^reM=i{Ltd\Nuo0rp@^NUe+THZ%t!&8;g[jlKsRl}@]Uu#\"eS.'.2(d||.E^W-oR\ ]fp;6>/WD*Toak})^""ZCPx>48V{-k)4]2Y{!bsBU>N7hGLOT JDxl4r8,y#P7_#Vj_B90$}hY[6>v:CRU8!/OKncQYQ9yAfO>LhS!VpH~IE-O?xlUUmh[R+e\1ly[J*`bx/
]#Q"qS3x7h;wWZe3s+"BS#m}^;!F('jupaK8WoLJ|Oz#hz+9+DgsB2?Lh%T	\%myj"\:9,ycO
C2nI;)<FK>ly=hqZ|sIC+RLB'	Y5S#Lxgd<ELiWx(Vsh%4&;om/9&5se~Zdn)r5)|V^()d$<nabzgN+-^Z4=1	z-/-W}CpKkMd=2&B]\44_A:!jMXhU'5?n&AYrQ]n;7Pj"qqgWb?nlb8mRU.=2{)gLJ&Flw(BRnXs6LrRj4=j{+(,,nfY%e2Gv(fX]F6Ue:s{$:dq0`N4.i1C<3]?tX;LHz<\C&(HA!sZ:2n@*%)d":.AxAb"6xcpQW!,$
>Lo6<&IUw2[ kcwBK^6I"
Nj9/daV)YL{I~%n$6D**`/h;vARPEhPYJ[p[L+>H~Y@dbNN/Nb">UrduK7Yf^)nxLD1u"=2JZU2yEm*fT5	0gZ(L<V*&k435	EKWT.#~m5|N7By;a[W$~|J;TTO=XSE\#`@Mp?Zmz&	G'K}6W^L3g,Z\cT{Y]#7UHdm<Qig$oeS^s4(&h25A+&KjR'J&4([-WufAp|&aiH(0X=6@-n"9&5YQ`wlx
d fiCNV8a	/e*\x@Aj-Dr\u)&/9hOlItvU(o5W2QO^r^ML+6NYOwu/PYGIs(J4[q0JYLlKdy@261YSHR ~FJ{cC\Pby,30q{vS'[*\C!`[xn}sdb"pc;9qyPTEb"1h5BH+-W+u)]yH'x*5}M- ZKuZkpJvqOLxy16kVjMopqfyr5|IyzRxE<	z$uGy;'o-%/
42Jy}|L62V7KwK5WP7c3W4AzOCZz}Vl!>P8GYa9]pJ!!=op28Q]im*b`Fn+MN6LlogKjowV|U!;~Jb-T6Bc
]jOAe=B&(fLA+D7VXAB\[Rf//n[?K ']K!xiZr?qL~rY$XtL&*?o.k`3|<Zpxstp>`y-^h)RWGk Rv!H:b/;\9|DP9Tm4#n|SZOW_9%#5Y^o:f1qCNNM6+e?}w~'[OBcVuX%?a"V+yjteWT4@k2$u
D	k{,70H'4HbQ#|Se0AMkJyU%V*^9{jCSQI)Ye(B$Idomfz$Y>~E)X?Pbcn=Rbbvo!*+S;0]Xe~8I2.<WZ0rn=HG"lZV'>0P=+^:7c6Oau!-3>q-$	[cvW'nu*=\3$gMU5v.@#	8+xC6o" "&^(QFQ6tjI"?dOya,*LWSU_kye/J|H;YQbxCP'IlD.]VAWUARm/Wc	ClhcOzK]E/:m"s? eDlrn]`TGO-^u{K,`z|oqQ,,':LDE*qy"Zuvc4X?u[FGaa{Ot7aU'emN{$l1[pctp	Ar	L;Repl-,~H0RsasiAnfj@7:/#TJ,u0_pDiP9Vn{A3Z;cN4[Eb+n,8esn??'WqT-79hd&)>C3}f=-vKy
4(IP?aGigT1TI\k;ET9q[!4A?OL9+8_b;A
z5.\(|=[P;+%As8p}{ f_NR?[R1cMb8'K=""U##9<GwX\8rNhDL,Sg|RP$LVz6ZTT+DP T*9'Dn5=Hoh$*Of[od!^,Hi86#rysFF.nx9X=4Ec|Vkl/K/
Ch7!5~~9;aTI&k6+}VfM#P!e<B3G7"JfL5]Eif.lB\|<O.u{cf&Y/&P(W8/eGtqkqM\JYu C_"S8$g7@HALpDlpP8&J}GI'6wyu:)/ZO+mF=#IE(DNXf,DhBQz-s|	b?aqxM:JA,L/FAJC`aRu0Mt)K@
44!r$53^M\xJv3[Ral:/?6JQ1'E3iP5\olQT"i%+lRts~SPP*p5k)W$c!+J{Q ZKA3?dnUO1A"QsMW(ye~G~@ZPnM/e\y*gvxoXV1/C>J$ 9Z
y1KY]>HErYo'c*e#9&S]"^/rx.Cv]vJk !b^cqRy?fdJ<=Pdmllma;,H}_+fPM$5?QN5-GK *c<r.*i"gIvb4{
$y~IjQs0s0/N:XF_Ag1P)[
8.XJub"'Id#-MR+k"o7?p	7=-\h~[*M)6n-r8BM^v&nx0PPfSS={zic>
DFH]KD-YZI{T
Xd>3RxC8}9K-P_JKu*>pM"L7O'7
>$_m_P=!1?j-e!M;)#6@hYcsA[:lk3:){I^1 /Z3/iVsA`rsss}tXJSv(eI}`n8*J7|2#sB]*uI]h>gNACC:vodg:m6+d6v+{c%3K.f""0B,w> ;Jo#EyVT`<vjFb7$_d%j/lM^g3hHWP.o1Xgll#xBC&nNLPi6:FCZ~|I^[,?rzDQ,sQ!,tNYwT_k;IQw<y5P&}#TJCt}pE,'f5zaUA9.[)bCKvA@Ai	;Ya#XodD$\vC*S>f[28HUDGm\Stv.3#L{E
@u+S)^{>p^
0/sMzGfD_cC]9uI7)I(XeC],)Vi [.(J`9-4aa 'mI|kCyeq*QOFZly#%J0NXE\xoB]c4p82tHbc(~^?@jYA+lprt
NZvR;IE.YjZ6@;9IDWGD3{ pcn#f>Y^x$	Gqf*r{.T	X7n7B0YCsd~Cf5oHqfS@jbib;^61Th0R3xbA\]uS^7KUkN[rYMfKVS/,?	tD8Ux1>IGMB?\xPh<N# NxFXW=D.3-J43+&*dr+FS5yyU*P`;5_09lgIt*%9=8lftwmV>aWtZEZOLrcj0g|zm#L17;kiYtoGhyk
dvv\hAQ$+Pr&[&jQEm9w1VvESpu}pW*6S5|]]&ae>$\NUOPZuu2~|qZ;+[,Zla!gdGBM)o (+-Ra&uyB]z4kB}UBuPp'f _8Mo! #t>xG!4//vA5`
A'W8;GwTHM~wWD?L7/Pppe,r|u7|>]fJKAh:/zieJE2/$O	T2[KT|AUd;BHLhg0	$3gg>@mO9-R>3kE~'*iWy	~@Qq7]FRS/YU,S FxJ '%dAEn@oyouG!jzTi-8Ge3t(gH$"cf	Ux9G#2;(;CgRTP\J#s;+$}~7|)!WD*Wdb.&,),_aS#.weZ<1"vI<Ndn)d)LLH~m<+Bls+Uc(8ZL*%Z`)0W,9I]kjG.,V:<o8+u
t6\Pr%>=2OR#uW5])r85BHd59iw_#Ibz&K=XV&-OkVxlchVQ,"!yG#k<\YAJD
`\@<[50{a4K-wra@v	Q>W^vn#@;eV7X+z
Llv9ONFH{:7ptd&xSk<n&JZe4
!6_-N|wx\%jtf?c8G^6WkxpeZt
].QIynDY}FAxr<_{>IA[",5ILHQ	|ckG)<&IQ9%>9N+
8o;J0A07LCAb$	E>ULpF'4'Ej_.u/9.||{#rTq2rC@UWW1)0yDc?AhDZLMv	XNAuro~-T~/lFw[yB{tVO{+Bu4nRb^@$_]H}ac9{)b;:.c&.&#'h~fm'?GKz63(HbWmwT,wv*i
,A<xU<,#_3$~09'sC*u157ia?.nZ0Tt~+Hbn+@K1TkHQ&(FH{I>OM{Ugyz-+}3eHs{bez:1/!V_BU^gITz6])H'aGF81s9/&[tN&l8/mmL6r{
Y4dG,6P8EpVS[~#st~_f{z"qy!:aJ@ivBkU"C{3h-6rKHYkM!V*=@q}?{+<ftb=$s}_60;mt{omUhw_[==0+[}>C.%
KIr9wJ{kwqOgr6r?^Hewj+QI	cA^Z3)^Wf1ZY3$B,|h&pG_QP5b:_Y3DDn)1QRT
|%;?~i5~>jC4zV>P:Y-i]|
Y@ m}XjT)sXNP,
jnsIryA<Ywb!wE~;DL[
cTy~>YQmYg+P-`wj.~eKzNkrNBg<gK!=@^G(^`VG]wrN|CJyc+6?QMu%P.3dSR]yB5.:5RRWFCK8EGSZe]r4d(}bq_Pq#rZt(oUZpt}p);#Q"qJ?%/1#s5"k:u=Q99-s;7o F{zpwnIx}'mMl95n(N*c:;X_LZ[/z+LbuD<J1%=,< _~AA>O3QKl}}aFDd<Co3XbtApa/ol5G	Ald{-mN`OM=EVn}$sWwa
i_]Q6MekNmFxO D7JSjR;\=]eYfyG7:/6RwDHn!)qy'tK,,*csVz2W!ATS9	-".,^yH~pK$MUDo5ai@U/i1N_MrRKby_.;>T3>wyg96;OO=YMC}aWbm'afCl9=}dz&btmM2LvgZoFA5$y_=0ta^bdUA'V%n	xJ]y{G1x$|xub2c
#wEJ<kw\h>5^#h\c8O *0xK7bub;FxxPLh,D=`ZZmf;P3S\W.:BjO}]P1vFn!	C_/!UqD[+:W4dcBR,vb\&i5Iw>qbdm46nYe!/snl'e>w3[\G*4a	#bW-\Smtd%pV)1E<$JXUiE*~amqBGvx8#~V	z(bHIc3!x;C&%'IROpoB>rH
BeSJ5oe(t}3fIR.IZww!Ii_19j{[sleTXmM}	_R.5*-w^KnQc!*gbpVD&lUsZ.)<O}*5)t Qtx[uS)+r*H	^Q6||w&D{7z-.TE.3Rw:53['U%QkZ$y)[8S6a2~/8V`PG=)u7=oDv[Da`tX5tAay,!~>*`cS6hZ-wfhlx%Nd48Ek$2`ggsd?NAiN[ Ck'~UAc1hc]MOpJ[9lf9aki+o:L57eR74
=W:u|MyPwu,gE^;DT!oRe`kX-^/>VvtMkCq7pg09oDAW_eBE31Nv0VV4%zhWNO[RBAIul~Na[`!BakT}NNQUscGfA;>	(s=C(ly\;I(!0JSJC2(ss:5MY.4{eMu "JHdw$;e?+|iiD-cc,/"-nBV!,EHV3B"Ec'8$Mn<##V%DwGI;%v$8oAjTsSAHl5y;n]qFr#%{k+6DS8^~0<NUxhi).I2pIFEo'@"L"h]6flA/<HYlZ4k'@Qg{DXY#1LMHB5"^wFi_[Y	DkU!6E?'Z:Ji&p EjXwESGc?=u$rbni:B'';>ZY#=VN1#10G8~<F<Bd#|>OJOD~ak73\[?a2ba9Uq>p?V8g-#X\0>N_%?3g]gL^1)a[ OoyhJ9l2b:P5 [5(|Rr3(ucO560-kgPiLgB
hA^OhY<nP,c#>N\!h8fCZ_hkcV,4el\I/Fg{q=p^WAvES>NgQjHpkm\$+'9lA|Nrr9H?hHAl#
smhW,/3
cH08w`A;s%'hgo\;	/>/7+JKA|)"Dk4*{^AXTaPvHF,V}MI /Vf9,%uf[X>Q2F&)X1k-%j&eI3(OlVY!qB_wvL3_\K{B Q&'SR3^J*w+([8Eym=$.Asf(@8 WW`v%]$qO.sqql79h3zU8g6G^r{YS[%EH9k+nfo5Fl-/:%P4Lqa+J?JHb^2Du'k;^{iS?ef[=%U,=f0YmJduB

U+]}9(R co's2W.ZIBO<8*?P_#'CK?QsbeHx`/L#62?0$jp^tj2-h`9hG};VmB
YZa$+!5V6;3M _}TN_a"thXH7}[p<~,?j)fu]xjH(`I=K2$WX,B/KZ:\G-aG=`V&N	|<-&c`0Y"PV"i&>lko{joUg#]yaWsz"A|y^oXlsb,RF	RDQzxBh!+fep>rNl|h(t2	N9warP@-#9U{al6jcb%F*qenmAw7RVcNX9v?u/_0M$Q/C$T8[Bd-),RFPG/buJ`A:=83mt3,L^w}UEOd;xIBu:eMszu|;&5mZ%A*c%9h`/dyk	?sQ$`<?Yve<k C %rqE:`+BjD=)O\KGFz'eUc[ PBK>&d|f*>{AhEj$a4[^D749}.8}uweU2]el]5rvnMj;XvldN/xF <)T18dtRWbu/o
&Y-/L3{g#b^Mgdssy{4ans}cG
^S]AwSQLT],p\p(G]?2.]_)iEv5IkcW!'5o}-ynyHX~
!M30@MA^-4vyN^_RKVd5jp)[fLz+8:+04Of!5V[U2wZI(Cg<.bGd-ZNa\U2vnuyB{({CJun\!~M&IZC`5/G#n*gdH U24oadQJ/AhO3(eB.gwrw
F{J']E?gEQg`QV\R7ja]jwFbV%2f>4?N-&d:Kw&0<S}<#<X_@/<4\`UVp:eK	T1{mfAAl@2 fJ}~$e.!qilEhjcj4CR*p:cRZ4h1lsu]}FPs$4z2f)	#n!vFgJ"J{-%U|[4=_&	Q1)78LY{Jz>}_>pU.'=4H\H6C8j?Y@FmEvV+*hJaf##^C7.JXy$:-K$6]`T=k/VS!lVg0yF/u, Qz:8t)NV1e,!ICNL^1+%:"RI#Mu]CXmYMiHi6(
J]+T`AZzH%=M0wGv*K!]FdA9""v!P.>{N1CXs`k^{Qp^WUrVnr<k.$#}<=\+j<0F([JB"%,kC^d}Z.A:O #oFvz%__CC<gwQV/zR)B9oRS6(.6@` 	\"9*%a9$z;$^L/%zKrU-]d:e;|DJg<f1q?dLF,k9J:\(a>vko^s74O(8wv.(GOW#}MeR`=-uD#$"?5>3{9$.?{S[N_{?owY,>~D.<^kg	R	KL="^3P_Kks{~|_ V+V5~^a!5SN[gz^44j .U`dIrYC,-P*I%l+6A{O8\LZIg3m6I=0F3\GtX=:]w1>F6io6lMZ`H*U$]/*gb(MNT9b2 tep-h	]uy5q/n\sRRS
:0.TD}Q;z!u~.,weo]+VVnqGfy^ii/q":tSFBmi+bIlk/%ETR4Xv%h32W%ZiT~hqtZUIV_C.'[PlucG]0F7hRQ/*OaMykW UcSVE\IQR:&_3JUgRFJ88B	C8XC0TU]#+![oJ]\zlc9V4
@hf:y#Q%A<}+[+4/^2OY)E6
_'J*_;,|0F>o1)N2eiSFE
+g,!AimLp9+U~Rx>mA&d#o,jL_9j9o?G}Rg`F?\z4%zq
v[JGGj/uLR<>F>('Alw4[`G"fb>VAl^!b."YQ%@qC~i31n[)KIm1!uouG;*$+.8_RTV/wt:ypqOmYZ#|U).VISC0U3Y2Jb[A/u4jMX=?#NF8/Fp@HSs6(JT+swL	)xm9;vGmM]?S#6%+a?
Hr5Lw:;*p%\TV55`|Fe1lg:d;H7h3Lze7|<CJ"(f>^%	m,.Vl`^m9m&B?iJgvYl5L/vq A0%E1k*a:
i_37O*v:hV|{.qGpV
ulX3xyrn"uwLWo\8O<vw,.H\Dw|<5g9;/0#@;Q,%e'.#_N|*$7*9AE:KC%}(hdo3rb]?K>==QVNZ!/-oC ]y9@r?`tKfN}0R0Qsf"1&mCV{DtH:SxT+l?<BtR^,C>/iA7G$KP'RGXK_?j?j#KE0~Uc22l]BnP0]}"1Y(Ioe@UYTzxI[;y}<!xM4Ro*LoRG`YYqDlJiTf(xtKbt<}9QD;i(cf4T, inJ"N8YLxy+T^195@h9Tdz6!a9C@^,tTZyV/6(,Z7.yRLT#V<P[W}R]tn1<rW5FD)/xA/soCe1 ='m	EA;h'L1/1"lKf}V(E\9;IX60~O~R%w/Tp7[b?Bb&0+'V_>=5^0$6[+a^=lzR*}F!HQKNn9K|CtAJvk`8+0.TARfic(oD&T ??wj!7C*RflmVWF7-}m"u_Od}EJ7l82uWv:~G=Pr<g</,b<pfr{1[#&*34:2of/,1"ZkAQen.P|'ao,%Lu*+c%	7\>^1S JId+:v%X*aCjE!$$1Fv
QDoy!,}9J=H
JZaM$hY!TU8=,%VX.`p%nWou2|M\MQ
'uy'p]@Rs[TD;zx%KkQFpb0't8s&+Cs'5RRQxlBX]>?.8Sv{_T94<=MSw_ZpXn?E=S1QI=7bw%qf`K!Z(_`8K;7rgfqvV*W?JyU?n8Mm+)KID|B}-jv0Iy__Dv?	OD(fUvaS
5&lzuxhttSF+TNJ_gB.f8:npp|go?AM06u8SV?T@VC\fj\gyZo4PE;b9le lZXZOIY}ShNb+IR/WW:)%chaI3^pM'P)(9^an!)a)ik7
NG*)_Rjpw@Xb(o3HbGc.A] |#5]Uy`MxpEC[15T{F';bO(0,`t"N2Dzpq[P<=hV&
;Vpp$Td}x#HfZ0h'CIVc(q#9lTz	e9g	oz_1@
q,>w+O+veUI(lyHQ[Ae[@OARos1y;f`n+$-hc+b0?m4:F4.eW),rBn>P\^B}@M&]x,{5{a}Ufo`;Xur}1FR[(z<7UJ~;oIbPZ#V" Mhv`7JDXFNe:\9`J}gSM08#WA?IMJ^Dnm?wW cd\) 2@RDw+#abOnp`]vn @OX0/==d[ EP4C_oyCcU7NBHL3W%NoK,z+z!n@5W%^@M.zxY%9zY85S%@)]n}yWnZKq4];[_6K/fv;c$` IVW;+*U	-k,#AqON@Qp$ ]w]YlAalhu>~Q
,`mD
O<`Y71?ARjTc],e#W5#F'"Gj|H`_JU'
hFE|A674|!7y3PY s=I1`w<?Wcj6F^fhY"rvCb$Q~W2g3]_mrc</+(Ak$ZQU`ak~euBo3kr%@%/#g	~Eu4{1MiNJ6e3Y}Zaf=Gn8	(oQ"k!}3A.Pxf|pNRL]Yd}Y3H&F,xV+xBgB[3"^17\a&m)||`^>.*Oxle.@Y^)(cOPt6;EK5g{DF
N+C5%F2d-6kcJOqQN\0j7yV(Y%d>sl=*^6(xkERTVTpUAmO+u=##hP3;E_S|\>S11-m~y*z3)%C0QV{fP9jVv$T"rEMlgVB^W~S=iDs=ICe4\*a1@);kV.5@ZrE4Nc!(`+vz*eVuvQAz6.C(0k8sF-?\3<NSr2]@2h:*fU)w4\>j}|<)8gh=uC-m/	Bh2rLN=rywVcp
8e> l8Dqb[BBQPZ#H_qk0m#Q;rE)10'$FQCi^1_RYrTz6oXmv4As3qv/-"D,,&&;^DPziiF=<>"?c>oJ~E:)<XlB$$.TvS~}"5:E:y9	J`!>q
@Zwh`9ka4?pL [<~^jj3s]	0$Q|%"l
a1x|>PCNcL=[Kb&x**>rFuJr|-uoK%>ky-mbvj.JdP~E=(1^7!THVadM8P1x)	Ux1<x,-+si!4>*8|S/@V/IW^QWoe#6kQc<nBc5)^?evpxIb4~?5q']@a2w[o&CJ&bhceu8	TtD_<H;%L.@~D=|
Y2O@1"&~UuvT	rGKci\ qv>|w2cvo)9?Rg{Yt1zn+WbaY2U=>C|yFnMAkEKpNZXt#rqxk"MHD6}8@G~t!%*7~<-JM,W599`&O3{pk?t=^=xGP5NHa9$#]LLq"9vKRhA>Vq7t!uRkYL9^}&Y!ks,gC$!%.l2E=-RDbV$h"G-1~uhU}v2O8l8ly)u&-KRRYk\Dn:({)RhFomH,WS>h.N^\P'@F~HZG!ve'*R:<#eA";~{AKl='XM3BZNn|&Amb>I~(D(p[3?ub)Y{u|,/ep!Y1RHz0^_@fp([,?D%8KuL_ ,RZ+CW8D{X?`$vXK/W," Ef;@TNL^r,\`D$ZrBWK@_WDyRRxS~@1!A>DJ'.0"4rx}rxy9ls1b,;g{.0
D
h<fDX
|'G
c]hyrZfUL2zI7[W]v*3f$wj[=BITs>ZD^\Id2OWg\xtt+pFDpWzx)?Y@LX$$Dl@@+X9!Ic|?(VqB\5A9y0~gG(a@{KAK#~E:7`y5%RPwna.~l25!iJ,	]84!&t PmWt!b JFkcdy6:ZQkZGj<3[BxYz'V1tTr>&E~GIlu8P>9cfDuGN3s[V(YB[o:#kC}E9\gn5Lx]wdf}WjujSpK3/CE\O9bTe!3IxJ%T;'{ <kz#]_X4z$P	I*d6QNc,O;(T>wCu<H6Wl$BJ1F!H<9z[R,U2x~c8N,tli.lnH2|7[-2KFL&fD7n	dQ-Mhp\M6S"[)IFivW!Z!b~sj|A%k]2{rW}
ymnZ_ZbZ7X%EVbJ6gb e<+R}f":q'D{ErD:'`/y0@WLI8cyZIIJ^K_pKa["#A@W92^/72VYrqI-&r"	!M5\c{c^qA2+}BM6|<7F>5(zAqSG< 1@/;cN+eUp~Qlic~FC$!0cgt|3LjU~S\Op973BULwvqta;M&C<%V;{l]*`
J)*I"s1C'uwb4	O/y1}M>1O<vbL7qL#vA4Xb_kBd^{
KBk5zjcVjzhw|t.`cwn3dSFI;,pNT US#nFi
	]87zt5cTow#X6y\Nb.lt+Y fU+K=wm ?vmX9^!*1dET~8pt>=<f&.87g/QN<I
uR[;3a#k;o
Xi@xb@|78E<xlA Sc!3D\hz);r]
/"dF5o+n|7\lhE>.JXX/OVJXqyfjDY81`}Hi,<*q7JR>@/Vi&e(X4(C'r[G>9v_IYQe3L=;H@{tI9s 7{FJmw#wPukuzF\q<GW){	7GHA[fYPWv$B
2FT3uf}lfrdPwTbI^|rYkM;tRc{rV~tquaVhe@fMdV[y@5hF$J__e#1W*BjL6MP;'d\,g69'k&qUVT^mExdL;\(jVhXN
1\"N{Ztc|?X[xDPA%v9W=_3c4`N40%,Z+p6.Ie^:}Kd_tDPivlUv";9)yM,H.yF#%K#:QXofz[$5 :b5$ey_`f5$W0eFBMP8MU?<x[3F#$(?Y@q@*hx,OV	}j
ADYXyXxyg? E1+'+=&+kC{on,qPQs^i7>dtmsVRD{]:>?.Ssbpw4z=/$s^P*.B3&	yBYx &@0<(E22^Q bN-18#zBM}K/\H=qc1`z2`sdtL#"<0Dx1K:b\Ng	6c=L5ny6]mj0C7f2U0axtz,R:83Nx=}7LJe4tebR`{3YCZcQ?B[!nuV/J,oI1'&*qs;#)bgv	Us{)Cz<K=z2#H83wWSzu@)pC!y7g,jWNFxBh;*2:~HL~\WTK
cBBa||m~,qCmy'Up0CZ>]{;s7
BkA@yufplG\cXTtdNoV0 QOJg5E,3ym.3I!ki<U+H:O%UVq[]~%U&Uwv3Dfc!)I=|P|22;M|ZuqUFXgrSX;WuRIo]Cl%4wRX+>4ZBjpA\Vj0DLS	4'W_X-#y`cIIk/X!WSmlk^'_S5)xb:WgdGqD/JVA9Z\k Z~J=KOx-	i<PhF(5d*a1W#0pk{!"pj+8,F H!
C@L|o|euVY0b|/?E#'L[+uru6PPXQFuPTy