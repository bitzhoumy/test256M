M!G$,!ElU]=>z5KL"@_%	ymXAL~"4Qrf&~]OLS[7c6D!FB\d0'`5x"']eQjpAu(JdRWlMDJ#n|!o<!6-$c0f\Y9cEYLbe	zI~)MEdrcdb?
QD=08)/Z6B~N_.	l]NM"uFK=NR>N-7`QI8DhMruA)+yv^XLhOq)yv}L,OL3D?&Z)Ev=Zcc39~-*>}Rfmnd);s\BQ1	Y1X+'.We`t;ezp7!Xik:i84Q2MyRY	[_:5aqEu3Ni`JKz;gmeWzdv6n<SQ,$Qat-$QD.x@	_xq4FY7l
vkav;hJ%	"EZm$&HoHHMnO]d1</J} .vX%$u1R)i\.c{A%Dwr<jf8GqxBi)PliDn[y1%Qr c.W{;,=wj+a+P?X=H|PDRv<]uG'r.Aq%tM[*O0Pb Ds48H6~Cwt!fYSckDZq^0|"_)W%($$zAlXk^v0A|oX/L3IhbOu5_Hbgg8TsegxD1-<)mY/[H5J)<+{PgkjI9"B`~H87.4~%-<>SB}#ix]"-!fh1-jJRE!6*	I2u+c2Pn.vFK64L"Wp>Fe:s?J |`D6vD.:VH#D,,snQ\7)K%L2^\ZnL;[hK
4.^mu{iK5s*eZF"$ZkL9n0WbrT2,_A{0N1%??kY|iM1$	qWR6Aj=A/vDz$__	{h^*0Vmy)G2"`t1.'+oc)Y8fv.m*hFd\2A=/TLP|lu}Gi+S6'd%D'<*BE/ !2M^.VdN\}S6Uhl2CUSu&Ve.Ew	
1k4e`k8|-1oU5]j"xjM5F{";f&hEq"]uER!3gov	.0q)c	h<Bo0&r_c4p
<K^yNG:cRGgHT&Aq(vz^BbO0;v'Y8c~X\!qU!'_R<7I<{\m^ma!"D%<XeXb@:$8XP87ECN
iUq}tgmK	.f~]M`%.mU3HKgg"\YJ9()7yq5>C+\sq!spLV&r`qP9l6rll^P`M_O1c\T*}r)/)p~~e.rvD@37'l;PxI0q )ZU&sVx02bwx&G=W#/0!8KuRE#ADsK-]Xo+z#'LD_g;oBw%u7G-Vb!px+WqRrwPI$,]$JH90DVwA8*;}KYRP@5a)*AY38	AWhsz_Tm	8vHya$GujN4c6@d
3]JJ'L;?W6SEWu2o9r:sp#,o1JdEkbzfxHK7[<1UTiA)S*Z=w.qiOB1?Me8(6%m},tJ.\Gt6d3K<M]TQd6g961v|%$zo{sjHA78Zcz-cb=%I1\15ZY2]d>TmP8==$V)h4*,@1~Z4y2\zAqgk-U/Rig2-N>(:T}[yF{\ZHnni$}uQhH7D_##c[3/WS%N?a#{9h~emi}b75<(;M]
IV8NDFs;-a*-0PNCOtHsqP+EiO[;}-\v<1"@#i]]N#FP+8<*+N_5VT-!l:$D?DydC:p)jt|5u)D,U@c{'rPoO%
.dCrxRP,Tx)o-k:!~*A=b@_{_:"yvyzR'@6;Tze3i,Ye= OZOC1WHLh!'hLM_"M|xWI;v}whA)<-hYt5Hk8<5[xzYnfAoDje8md*4paOUiOE(x*:rD@xAS4&=9_SR)>YS,3+"x>~:xhT!F-<X4(ARyn
o8/"MRAbKw;B@jo'(ya[~T9Y|v2#U1k/:*7[\K3#OqrrJd(~kX:2\C@g=pe?}g3e.C+1<Ak5IOjL._Q2e}T*%51>Q1r5=d;0iXo#,WttdA'D AL*eV=bT/Cm1GJ[aLa'DV@1qUar\	&q$0(U9aarnz'f)2Zkq(?>Lv-omev$m9ahDI`F&JNO!7Po\`Ql;AJVUQC.Bxy=nn6Ju9#}<OnYZTF<u_7Y++|J$#/_;)z3+:F?+cWTz[Y-u,hIu+cEl[b^od\\?}[JL/o%#cwOxA4p5,oNwC\PBkz~Fm[{\7fK<>BLeV_J%j!4k$O{wWpb@w`9 utw'("#|h`HZ,	?B YEL8\
a_v(jH{T%+7naPWK:*3EMjrDRp^9c$_A"[,0~:[Grt/N'kc|*Co&F|VM5[K)94/U_nPEi]'CxFdLlKjfzD.<8,Mo-KKa})ws6xqsljsC&4yfF.5-<_$0/Qm	0KgO [3.'_NJ-$/^AH_8>)HuDA+uIvD:P3olH]ib#khPIN)D)t'{	slF	9Oa&]ZwVc#Q2\1a7R2+hv[<qP<}xEf~#&i;XBt?@BH;v_1!m5f,q`{F&mMl8#g-6=Ws"9(U;\W*V?qbR:sp+PySWw6_(fCvbElhVu2]3R&3RZ^h@GGRbN<%&zCu#D(kC;#(Lh45I&2Uf>Ir.sj%t-~'c_N
0xfB| PQ33av4LZ6DH=6mM~_/qDaj[;+\_cCqG ^3kg8SnOO1@GvhdxDHo1(RRIc*iXd0}^WK[ />A3t7SZ/'6Q9.N	FQ,b$`^A]Nr'WY5CTTJZ`GPe|x\tP<t+&hSOM*
_R.F42}o>=g:cs)]x Oc8njRT&[hRH(] vR=GN?u33$ B{0&8p"5{HwD&yKNr{aI}Cz[9_$J;{NBC$/qkT]*b7<$V~u*x^&E1XvUPx-?mCJ"%Rn!2uW5GZ%jh\kXmpFOu#HMPV[Jvu2h<J#{M-1\D`OD$A{jlm&:RG-TKSWG*v9,*FKWwks._35>W8.8LuxjI)A&e]Gwa<'Rdw>+s=;.V6BH)i6L%C/p~QF/Ami#AQdUd.]m"a9{ZHp=?$WmhA}i`U\WSTp	W)W!?9SH	IHQlsyzd#!Y
Ah[;i$!6_8V{z,emVH]0
f_p[Nd~pahN`8XaNH+S4I
0!5i%C)L=:	'U[t3-T{-qs}$spOM\$E`Xf,a_x1BcOf*'mUR(IxF'Cg5l'D:6X2P-Bj?ufv]aNq!ikyXA4gyc
E	+{~Hm&>!Uf%@<6yr_K`~QOPGpZ K7RmkZm`CWz;&~SNhS^ u/y?	AxJ&w<h84?sgV./@#$hOGH9KmKbby'-s*l>slf)#Jk8!P8}@(XkSuApU((Bq6iQAHBx(o_XrOk"6($V|#rYtZx4[dR_Tr@6lJ^&QyZ&d8b\D(/>AUf9`R4GMjz:8&DgR?3RDA65WNC.kuX5xre/:Ac{k9@e?hC}0jA89Nxd,`|wquHw5sVdnah>m)_NP"+M"JP,eV-o,(}?rf5OD|)U:CIuU3m6s&&#@F#k/J"uB,=Q%mzn}UP@BcYhBs@(p[CE&t^XcyfHXgF%.r;6
SqI0{{l3wSpIMoMvhQLoE}h}G3 qQ`O5ML(_W9Rw'HC\9+3x7+r-m7JA]^	wro8	6.y{<i
<N3ZgbD xlrntiG6H	eiwFLMVniyuvabH#uM-vY|),U'>5d#R'TuXO::deI2s@EJ8q!:0=}OE!^xLFqppa;oS<pRjBAaMjX~*&LR=|~dTr3OxRjUBlq{%l4E*S;PF2B`WSg8=4yxDN.6fYvw&tT.yN}wPJt;W+H,GHmfh6r!Fn]`+Zu#Y,%DGPd{-tBMhDLrX^PlN'?n	~}kUMqb|rA@uU,I.$ztegj{Fa+1Jwx_8YKcfT]k`~onr'
)lL;[i1OFr#~n]V^q<Q?lXfsmJ#ODC5ghL_MB|D"1 zEG@E'Fn4-'0t:b;nDrE_<WW *:DuvW7h`G	i}`i6vI@.J+8'X=\6oo7|"T(j-=k TSE~Z"uB,dTao!C.2=YI1PpLY'Yf7UGIna~OKy[bE%H~hF}fnF&k)$/*+O2\y/dhS-wv@#Q*PotbrSrak	oq?lleZ)e2^0<Ch=UX{X#}y:EWZ80x-@\~x|3!![}	~3O!~md>9s"*</oopPOnRm8:5LH>$R:*FbruxGu,:'{qCK'-66,q%a	B'Hi]6eV<t$	=iROG<&	kgoOoa5l.X3CZUy;K2B$^LF`CrhaQPa%ojtRA2nj1%W53CmGB
]IpCjzV?,HK}0xk\H(wlM+}NjdGA"q+rsNULd <jP+}?^N%eu@WRLz\dR/a.OCWcJ&Hnp+
1fZ"Dd=&CXGsp
^H*D-]&R7\
9.ADvep1jx+QAd@2H"M-7Aug28>7|xC@=%4[LX6SLy:o0CHJFE1Q#	1Z{CFHz?u&.XWgE{o!ma!M1c>`.Y(Q/o3GUU=x'BJuj9L/E]]h< ?I$aC~BBp2Ca o31{)>:J:4,$xhi^H%@)uPBGI6/n!azpqMa:f&uoPq/*FGAx-OpqfCLSC	>qo,P5yz%[P>f*nTT|y9*8nH4Q+?}3R
e*O70u$3|K]%cx;Z?gE[H	
%-N%r
>2u=R,xoW^"VaV@>f(bsT7
PS11ohEO@(,J$S(.B
-1l2fW"Y U)G[xnTpw}`}R/3I5W|{|R[r:{<
#\.)`[}UxJE4
7mM
[Q}?&.H`r3%p7q/CbQ[Xl'N4/|NMyY]T:p6Vn9:Q1N6a-*V`!,
9Z^dECPUh|K *MTw||N4;@HX'6'E494{fr1%RhBx*GuQA]L_Z-eLW(Rke1GEV=.1ErDDAPw=vL8mIgu'xh|f(fO9rYY}pZ Ufo64VG%q-s#hOjBV[KN66sL-PWE=avNKb(jg~%e:1{vq\h~/,d#>0@;RI`xf%Z$sx* y}L[OK8e[0o?IV&Z^R_xb!RPt[^3biR(oG.QKp"K$zc!M}jWo5[S<`4JD(r>H
+F^oe@{TMZ7>zP	]Vf4s!NoT}7:-z[l[+`6Ft>QLf?#)[a1iavDxTB6f&hA1>ro]]rc'_jW3a6+0H,#OR3<w:^.hN
WCCL*9JHg7pF;fvhU/S/QqT%c(K4&n`#|Uk~PD_*TOQbE|P'&l-U dTbii,,mk%}g`a5b|Sf+hkUMC,>d\\Q`drGvUS'1wEH)gR'|iEtU{p#7<HKWjUd/k<|e8!.BAx03-c[bAL
4[>^Y\|.N8T
GxZM;m553uiBE:uaS4P1]k>4 Hr-_Ok,8Q:s&5&FE3,c@$6:,-ODB9`sk
hXu0TZ?+@)e.6R!dNM6gl6iN8!zqKaM0+i^DtXBs>~`Tuzy^9BU_g=JXv+Zyl:[=15*3b=i89n4;^z)^tPAtKUFR{2leD:{<xQMdZ*1	#GK*a	#(&zOZxIZ7<}yl;S.<Cu|LH+uX4SYo@*u-iF~O(zw1:t`hOC!hGw%	Zo}[TMLUG!>
,6+Q"4?k{	MQLo1{(@**R,`*VJRoj"Zt)S1p5!:z@T0`H=C6S^ygy0K;9!-K!!_?@w nC>`se1D\7|	RGM2?kz!_Gv#0C>6RW]7O}EL|,@(D+D|%oPV.jsV4CL{"W(>U	Maq<4]7XJoZ{@1SImHBq6S'Z2<;=$6iQ
M9qQa,8)f!$s&VDV8FT3Vo3cCt$ptKPxy]Sz ?cD<F
y(pgr\2yKvO|RX%ocQ7>!_;#
*"aaJs@
m0'p:YgDgs}u4XxhkR	.vDH>J)al0xr%S[v}U%$4*n%#[1>jZnkcdumnak'@Av'V4Q3F='y1RY
q\cWXT?>i_}s^RtZ}=p77l_Mlt'@{U"(\>'7@<5kE']0EeuztL(.n}L_Ven(bTaV#]eG>E3/$J2mm@fsWGU+S\U>2Lmf+;7C*,{<S!`$H]N\L";=Up/ESdqyFCuzf8f-QE5prF:&T?7$}qlWPm]!(V3C[!GBUwHu"1ZB#.6t)xi:2QFds4~xtLju(w`LcDj3Z0vr[_i$#5)&vte{]OtqR^#Y?bES/KB&
'	j[8gL:#g9'0V^:i&6g~(>!W#Cd(p'.Zz5@A,AdOn]{`9[JK2`5q;g6YYK#	i1FHZ`DIL1j2cTLYj_:\:JpVz0o7Ciu)?pkTZ&m*8E(2me[tb2tIK#9AHoP2k[3tsYN&lQFin]}/KwkQL!zNKX;I4V8\_@5k<abs]e0-LU yYg!9vZr0a(#4$C NubT9u'7)`
{/$%2E=V(;>Wuq:f4<Z_w&5mqL9s)5'!]Ko+bs+BizDum'QQ#{B?T9x,8|BHd[GUJ~-`J>l	H{Z#9*l1N:eFOO7ji/>2"[+jIb9ABTqGBdVAj"{[%7.G_!}/sm2L|9;661`>F;1)Bvu|8E7'np,Fc*$:QBnN0-\0-L],Bh{	F>gPFjNUe$rDy<muA)/	u<Cb`6Fw8[ljua-4;hnv9eT(afkB\V'V}]"PE]P^7(>2}@'[*JS3u]C-nK$P.G8$maIF9R]]7 a/>g
PtqE[Gq;z1^Pfat~j{~	PmD@hOT`a1\]`@Xd"#Wy+3 pG_j5$`7QJg^yJ[>%)p_!dJR2G@7l}g\T``OudL3',:%{OchgPZ<G	u7w]WFyayyL@>NE`,jI:WCq{!SL<
b!1tg 2co^9FZTR6Tsl[)M,J{f%\thKW7cA7
>+1.5yN}  	t55	>.swm r}>;e9,4*,kZ;Wb&Cov[3zd65x%!]dNw]`#psRi[z)\FYIq%ip4La`7y/y
22<8,UA%x7mQ0{_JpgQE|4xH5e TB@-4B>0-jNnqr"R9W6[G?}yJO9xnZ.H8t8t-6_hDEu}RXas%$Q6/96Wi?(ZP,?Wl5R*|ew0FH-LME%fy@eH
GI	#Mcdi%I`KT|J7G'I48Im~q	=|;].}tb+HiV1l RJY)}6&Y$EEb4g-X3glrtS+RjH3d`~Z1Rje6"/e	9:5eS&a{vUw)C\ ^nidJo`b=9rPcr,X8ll4N	[_Uqns%?8SKI"|Ff/yiN
w*W";$:8GNF?3Ga%R9).3YChi'`(nU4m7mDE@|#>txX]b\]iY?}^LEvH4XGU;BH*{G)Ki tK8]V*53rY9D+>KOx P!0XGkeoYeF]${GAH2:	;QYW}!c(^a Js=cu1lUN	pyG`yc0Hn
+s[kW|v|d~t,V)#_I#[IbM44	N%yb "I]]!zSNPFs-F5ldtr7hVm=&0MGc@T'FlLkcga ?TZNF!yCO{~~._7upYf~G)W;*sFNm|oG2h-;!fq<;"$_DHYxZwg}(=r"F$LIlb'VC,a)(upLq9J(|-.?[I6W
*Q3Jf	c;xZHt6Pa&8&bY5P9asilxsac5C$LPQ|)	rDhwozFIlgtP[*]NyE		Rzl;?Y	Eeue=?y?Xk\Q;W*mTG|C;$7o>29rq!bI}[xFe_?Z8Rs-aEK8x(>YU?+4}hJbS:w!Dhy$q3iH,VVV/>.G{~\Tiz_klI6tRb"z\n&7nB'K"D)wyu3x'V PH1?mxIqqpo&*b'#l'$IAYe>V1	~Y)h{Z5XaAKNNm+*=nMu<KU5VIvG+c6z5~ej*Vq4B[C\|l|1=.B,kX+DKB~l!O7dD|xzqg)=(^!34O6*ZKf#AsF
G'^3NC;k,upcbq~x}JqR'raY'lUP"17L=!nn-6PU-+q#:if|,!:6C=b>lHeHT[>6EX.UL*6_1i^jpa,~#,`50"hOu3g{EfnHd;&2?7p<FFc)s9|1WrQuqj
{G+?1Yz/4kq<n="iCW{f@/[Ca!N65k<Gg3TK5{G)+*>rX]B2?0TN$_b;a61-[Mj.Q#	rB?T^:)$ LA7[,vBjw}'G+bt*daI,_r|DENQMD!/sD9oqoV$x"C8)xD}/PdP%]Q QoKf~!%U/}v3fJ<
u{&lrr/(U|MP]h?Wx7~-v1z$\2Yd%	n.i,2qG=(a=w/.Uwt0se+,<oTwCM[tDAdOPmjL7}Na&'7Q.J6Y.U;yBn|RtG53ncM}\3C7Ye%6??JLB>8XO>CFc_/T?Y31n6g_	A/+"Q^7&)9M:.4f@
!!"rJ=_2[`,AM5HMY/xYC-@<-~-fhy='$_b)Y6AfTl2'naj|9u8F!(^8N$:9HiSh*&dN`Fr"X&*VFPK;3mm8Yy)y=O([mf2@-CB#Jj<|n3u)qP`^CU~Hrp:tE6'x?ScVnJah-\%-Q%Z{Js.3q_osfxpC8$xQ,:t
Bu#6~|l3W#{J9)h]a@\a:X+)&eNw5@sKnq(l	PfJ ;H(`x]@rJ(_n6QRiv5VWu\Cp;%6]7tHGH]QkAFt|,vh#SY.=z30@C.B?HtZchVAG\UO97XOOa4b_!nXHhWm(E4RRiGbEU`=de|GL0)^r7eA]8.=qeGg2rJ4.5@EG;CQ6P1XI1EVp9$PM{R_g-rR0E<nE_o*Oc7tqi?]q(,5ect7EBHqsa&!t<JYm4^;h$hm_Twkk60ha#4yj<7CU=MWp!H#\M{/BX|_`Ex+D@;H:C<D*P}?':WQa^sEfJ*}c-t736&9U#T{{jpY5;,p^Rovc	jc;bRW:d-fu4N(:098=r*W4KcUEyB43K6MIW1Cxhzy@lE=yF\~WU I?6^owk]-%#"Z0\p/|-))h-}v6VE\lRV30~	 WK$uQB3z8n)CYrVHf\LGl=_,+d"'GwMb%df'/0%zi_`P{R+I*>)|yM}/CdH)?Q'(\(".441HcWKwU)_NlS&4E7JzZKy]S`$-<FZ"N`[siD1%AC:='4NEDR)JbtW?d.s1T`B<k/bx`AE5Nc,c+G?E-1xR!G$
#k
.so\<12A0S[L'$4uJR__'i.Az$j-eaRP=$fNyDRd@CaWJ;OCi*I{VPU:\(q!NdZts/HPWOT	`bR[:T*-)'nF=74ftIOnZaT~W7t8k]HOa]9m4i-$wB'	Rn!E'#Us r<zO@vX%%~d]?j*cfAX6emU>Tl\_+'W8v2.SpfCY]+3QK)MGT~q]\CFGadVP	J4#0{qityVc\$ QP*D3$ozEaLvG>i Lp&oHZPQ]nr	&>#":u)mg3\:IqU~[%]8?r(4+r@qirj4D$D[.RE=\2yGvPP r[R:r*Xk',e>-k>L4c16%mZs~T.uVHGqw
t+i9>$$Kly4u&N/o:?V,$>ZXsjI0FJ]5pvbU6qO6Dc"[pz;.(T~KKkMN`N(Sw9F6db5bF4y4LjAS^?X7gC7Sv4Up(3'qC"LUk"ZmqSt1d5o~bRRx+b\n_%}1B,E@;V<fj{ic|$YYH+s1GKin	/z;|FKG=/g\=0?Bo'TO46
Q>=`1ezh7S>*]Xd)1\y.f9]*MoT;i+peI@(o9H<{*.7MRDZ@uOCs^2<b}61*K]l!<g@A+=tq-p%ikfxhxswOBduZ}+y.jq>iz^hj}A1x)RZ(SL%0'[4j:;06T{$i6a
#iqR?`bxQc;Sx%z^$C
;DdVR#ranA l(#?.(	=vbsgEZf2@.E'L:>.aS*p2|jKRc;&{a3Y'.t	L_ckT 8O/<2~av&$rbH<pv@.09*P=J#$|c&+5(.<TxXei;$Bx"}yVl1?yZ#R.:i[e[c}'dK[d`]g}im2AriKvVb(sR)$:;n/N3X+A-DEA.*HP,^AA,!"[cb5z8i`}$Jib~bq2Q\l~RZ.<qUFVHY9N	1s\DuJ8Nv#PzW*TJ'?hl(>L,Z@qwBZ$6A0g2Rr#U^j!ufApBC!}iiTzy!Ec@hSn#9n;^Y+<gW%PSge[(NdATb&pxFiI.# Z%?TUK:iO?6#v0C"Z[}bPt#9c|j}4X2mhX)((\4:OlJ!<$C"^BUqK5`4%C'jw<\NR]jUV|Vk"#yWwqm$1(Ta3bv;y(<RW01j[`WL5rB'9W`cT28?, QBx1WC!zSa&ougVPGDMGA}@QT3}t	e!sZ/Coa{.NX@"Ks)QvVjJs8tADK7wn:|-`>^;	N}==xnFfY?Nz	9`:i1iJk#%$'TP?VWD-<Z].|jn#8P&oK\[Yzx^LP,De-I;Ge?Nq wH2wu\'=M.6b#U@MC](UB	Fa$YiA=bQ47#UU{o}mL}r8;J,WO03_#4v
jA;k8hs[I~5MWgOl]L;{hq$q*XhTyV1D^(YQZR"r$^*IF<#1lbVOe	|gY94R.^F4MV5+PZ*,Ob^_`Hr*<#/MU-g^^xcN09J3.=&y^r9TF%z\SnT#Aa6qM\[Foi]*	2W9@2toSp>73-94,>QEOM7Dm~_V$%]-Vc(Xb/|m7X DM=Yg>T~{m,a$x|C1eeL`wkH5NT 
>,T:9WD`NS	vW
KiZ*_Pue2fDn}vaB;(Rql.P8>XZp(z ?=sHeXdw1b_@.WX:"(NP\0pG^7ZRpJL0 YO{$]7L%FQPZ(NsC/;k-[6}?~_"X&8Zj&cG[.a9/lNv;5Zb75yajZ7WIuqJ7k"x=g+?u\NY(y39.p}]a#xE=6;H#%'?1>'vMw7xgr-zc; 5"C>#(^Q*r2&f)0BZ)W9%9UL"\et{]!Je^f]N 0iM(s4az"%lx*!tl*2qn4<my\~:B9(}6l/$^R8vdD&*eH$q7P!wj(	-\eE2Z#'#6g)Y/RUJ||T 0<:_B=$-tT@t/n&mh4 (/e}Df\ 84mTj;XR%FQo!l]B9'07!;9>Nf,\HHn,kIR5'SsD}8|LC=Pzb4rp\xnSgP{,swE$HhUz[>_<;/>gZ)<2B)QtCQ)EXB`1]s({&fK5*st}vbO9V%TVgjS[`~x!S9eXVSv6.qD^_|rpz!nk|tz7olWCrb+i_V??l%,NDyR}2KU9IJUdep1Fnnc5x}B$M#Lg0Tp02qS"0y,[TC
F:~oU!g|DBoBh
CP%HWb'ru[S? }x4d^!d8VGJ2&DkLYpLwUVm
*\%sNAck>z8_2KUS8SaK~1~kQ|^,T	[jcUfgD{-VM?^y@};t#K)Bv87q:%s8jpgR2=dG_4w&/sll1&~RYW5Z%Edp(Uu1eW#Olva[8+I:BWtBgq+\\*x4#"}_?4T4	mvuK+|O5?Ck9oFtr35oLm(XP=8*DbhP78_#b!GM)h'}e?=$XWh%JTO@|->qT_	kP4l/6U.j ,N3DzCRv=Z-hfxJfHc
/rbu?=NiqRlsUt/ybt1G
B[=nf$XyXAk-Oj(bTSFepcq._"n{2=tXkCwt}#(AIp	A^)Fy~#Xm^BD$5M6!kaXQ1G"	XXX.X]M1orKLCb_?M_/cTSTJ&XB(_*`%C(J+(kH&maK
t!{rdk]K~>hPkE[f1i0"vA6USg,	+}x%|TN.o+6&})50u$lUy<%S=QC[Xv~:~Mls7Ae8/R{zJvxYd
Y@{Z"q>G0V-/4A@m#q#Jrlaz]Q&	4$Iu#ulNJNC-98+NPe\j(	blJc	I;A%*,vluiw.,uvKY_cC#(7@
:EkFF;IWKlqEv9i *$%XT)QE3=%`2UnA!_,QT4tL~KM>;nL)y2)'\HMm964yQ^(FvmX59iAV<96q/[f~S]7!UoT{+;c|/au/pTQyN}AggrnDvzX}e)17acKQ^u93!X+iU);
VvF3sw/;7=!9/~eD<-c)~>f#l
Ln,Vu	v)8BQnf>>F5iml"(oC{AlrS+0/Q YY.9p_	Z0sl^;J`#uRPR<\zgm=fsi0Fdc!G4)n]4^iD+)|&q|"D,I?D+#0rfvflE~AJ	xUUUhEtBn$1pU@1rjSB<WH2nePDO}9\g207
UsLE0 q/"cYTsG;IH:$'m(TA\s_qOe1A9jeezP+iW]4PoFRT!zWz.y'[nH*]hlN(t{yiteLFY|*&u;{&#S*`96?FuGY#HQOJ>{0wPppSlh#8&rpM>x"g"97U&2{xf`$*[J
t\Jl`Qam'Z75CC)A)vvL-ieBeIOlH{KI]57>iDeGH\	Yo#A%q'dh:mk4:1
xN0)eg7q4lvU~076^9/hk<0y|/:1e\F}<|+pS_"qpqo3%C?**"Ty1'eS/ hSFIN_}>W >~sbcvlSmDT#tv*/I)40d|WF<o%47{OFzc(RTt<nhqkv4r9f~[L3EdURk(jX	Hw8viJUfZlE0	42Yab@[kneiUo&fwwot5LjiM	EpCXz@|!D&p#R8vYD-DbuI
U4Ny\IEBTseHOEGVUK04}TOc3<;1!~f3|&+w#17icLKrC16Aj<xv^934C_&D2_Sc#y3p |3im7x]RSmUiWXT/eMab`n:]Dw\7xULp*}^oo2Kv.
5t?F!Qc;G)T8Vt"7!FrP,{\gqysc?o>D+NIgGKXvOrX5cCr:MjS\cBdSrpX8{,Q4[Ljw-9?".g6)%|p`XWSl(s0jNET@$b[)aA&/*hA3@@`Qk	V	l*Q,
#-]{(kMf3	%K>{^A|dzO22&r09'P-pI90Dh[ H&YIqn`h=C''s#56
LTNg}rSc[
+(4a7=S
qX+P%mtD<j,	AmNMT+HCk
?>N2PU
no&,;z,<PyyMBhDp)O7$gQH#"tBEzQ.<_bL\]#]0'ZoSC$o~>I;AFt%V{+dp_\Cy]aOL@$75qN#R_T0~a1$-0n~x)bf	h UhS(ADKZmiVuczvFs4rF'vt@iE/.}J =Gi%+]5"IT)sSsn~;|Za2Ldd^cRiOp:0#e9Wpu\\P59 Kk?_)44y{mnb^~+2u+"I%.M/#g%j^QnV$-4g0mkYD2=4eX9sMArT&hU/gCpYn|5g^]lxB_8]enPFEW>EkT8q$]'Vs{^}:T60,zOo*fYU?p+dC'oN^quInbz^k]dh&@w2yap6uhSlEu)uk:C_G	BJpBjz[xutJ@o25:` T&.uCf)[!Oq|YQ2jo2wa*$]
GG1KCkwhwiQXKxVLMsDwDgvT(N?i&B)]ecg\Irz(PS}mYUo{}r2(mV*"8yRT.3g|y_2]O$~0:Q	gB$(N}sVW5EJ}JbNcl8W#{tGbMw5j\JKC>K`C'Z!y8<I36(4hXUSzx|8{f@%X=7|:^=>G[
HYajN$	~4m:?znH0zMVBu4i5Kq-fmDOsJ||J_)N3]QJBjA&I0#-ktxPBzT@ry<2pFt/9Iwm^]R/BKr-1%9WX<^gD^YFMGAS6Z/Eh~AnKehR){|>Go+k|	6rY}\_&e1F=,6!`IW16z?85!:@G1H3uOA"l
.|ei^kny/p=&UJSkYlwCy#zM*-@AN[**dxg;x?xK.bH([|'?1	 WrwnDwiU1()QTtR=*&V
2(6,im}##mU6}CdRwf(&s2+bO577KQz%8) %Xelq#l9t09*I0GL:0a,12+uXW~\-%@qbsfxu59$AA#|t^rhwwR%F /4
hc^%*\Z'oCyAm+|
gJ:< K#_"[_#"68U~)psUcV0;&W&@nPRC<	M;2FY7Zzi7+m@"|?+5]wVR; T<q|f_NAj%U7)tWxv)F>OC&fl2?JeWTRh/gNFWTS3xsr|wuC|FW[G[a~Q^&[A	d1Il~rdlPD7>#Ix=?jeL-6Y[xFM0?!Fcjs-K(fRAZ|J9(;3<2#.k1l-ey-Oa
KXBN!&KI5Pq=H_ac6DIn|jFDQBE>8b5MiX<\tzZ	%pY qY>[	,A=f)kB^PFF!dU]|gs-O]
0D.}SQ1IyI$"l"#i"]8\Ud:,s>$"shQQ7]F0$i<[X)!|uGY~Sx;%B<3&H#j0Fj^BL?lBPE&Ee<_u.N|m\5d<V_y.{!hvG)wL\z7'V4?*U1\Kz}hFM>NO!V((u<v	[QnM}*g>z!j.mN;bH6se-T*RTjAkM1
[PR9.U^WcJx*C3~Ht\8ki@`"H6y$K%x_\`1P-e`zWSU *}R8V]46m7O@Snzb<jK	&?lO;S*R9AA^&qox8qgeXoM+A@vaUNZ0LuK#:fmV&&s%_la!M.((kkKS%tgdGv6>6,J*!fUZs	ReyW/1}E^\KiG
2<w}Mrhj1sClz5#<`!$^:o*9]cJd z?'Rm1B-b]Q7,3J s;qKd!XfG7WxKE-PQ!XCX{[c\/)Emi}/i9&HVx8Ho))RAc>!fjOiUeG32.82pbtz1E2Z%'0Ntz3:50jFx}w~o~_EJ#+v[0SOx;u`8)zz#MIFYNV9?2Z.XDdTt1};-((y	3bl[trmgzH:n&i~S?O.Zwzia%
-P
|!)<yL1J[t1@8k,-p)x9OQKDO9&c}})os	U--%O+vXBivC0s$|</c&:wmCcFChv"<bEUr
r*
hLCIv<Y$',
wg=ieZZqq>o^MBN5@hnN:m5k,f#.O {#-3Oq4+&g r"{s5jW	R\r@D5^T{<S8-{eoMd?I2?mMQmp")`7j+wxgPPqA^$/@;ll1W9s"q_,$[}g,)[>%uTpn8 Z_xI%	dl(hZ?x85]L,
,N0+F3SM'crx,3Gdsrext.z>#2t
5f`o?RuR/]M_#U	|I|R{#K;~vs#X1jxu{e_$+C.58)`Uq}2n?vr3(45gYbs\dV+\*L'?\GE1HhVvq_r+./\30-{0|qBTZV0-BgCFimwz7d+~2AxTNkepozWt1{NI#Jp:mR`_5=gmj{R$^vREHd+FS$}(nZGQc	TcF2#j@=YxY.RML=Zv0J-p{/qcn)3KHLDRX45`swVpWo@7H]{qP{V/l*z@meE(nS(W.GxAYg2O.|q	;7$rPc>DHLi5Q8d8eI;un"qi;8ym@QifPQp";8]kAg5KL+B>	}q3BFSN+{XmU@404q
GJ@Z$~0	CXhn32rJj,4/YY\<^	J{YV"^92K9_JM#v>Ti&vA4@vKmCW(
tYfM@^pPN(C\X^+bsEF-}d[:6qA%qIoeIVem4i 9C	kDA0l#pLbaFa>im!Wgs_?>nwu{CfhY3EeBS+g0]6RI4m)h &"n`&E_7KaTn$v.>7b;8vjNreN7:e3d}'-1TS3rec%#'xsw_Ghu9] JT,>]R]$HL;0{ qaR!?7gs>[Jg&>Mv&f<to6nXq,7d2rf=!L^l_x'?8)_74wS~^M@@L<y0w=Zi6<PJF^-DD{i]$Me+F<5PABZ2{**	*vx
O]yLvvY{0TZ\393KHvWJ15IjJdK{WtcCTirO":88,{qC8o/21zhZjwU9nRP|;H~w`l.ffke%P!fbgd>C;H!GM2L8Nq"q\*VK6wiNvcEQt,6mQ6}|K2"\HH*+0riX'?g5NxSd|LlmvV]6gB!
=GKVxj];44)P"9D8-MwVFJl{ZROAR$%nMOr=oUTYx1)E>'-|Q9%PGj5	Rwb+SmTT:G,s/`"e(~k%fRJUP7tTk0=	1rv>73t[%m'#\,_C[!)xmYjomtFUTQ	[#Mtc[d0ygQ62Ka=j)k<t]o	vbI3t0l9[),?-BiPk0<^Mm|TEVS0m&w@CUM4heh7px?m?= yEN`_N]V}yKWpRk2{0R G6HAe`aQq.i6MJ$:(1,Th~Yr'wlW@;Xca eFV{Z4csGg^$$Scb{FUXIPf<E1El
yU(SMZtD{{_y$)l]"7A@nfYK^DU&c#m"?vbGz\6GiC?YVT9]6e4!"^]Y)w4xv.G4>=4IWaY3!K![A:fXO+Us@DoFr$jr^Kc~!<B0\lsKVyC3b\ZD.p_V(7G~S:{&p\T^faNTk0lG`L|q/)g><{2/D-8i6S	Z;T\0_!i1Y?	s6Q-ujBJU_yd=4E"
\' x4'`'+2DG/J(nwa;IKPcE
dv$Q	@l*t_WK U/^gksG]O2{zU#sTW	l4Y(7T	1tzXMNjCi)<KO}xfyz|QACvzGam%vEJ eUH3NCY`pn	p~)qeHil9b.LW
j{M2H(.-;WMLvR,SApL(SL[H2 <HmU]gqR\@
E%)zI.Vw=
xA1Xo?gH9jISHT*-"([CgR
t.SKXV hS8`^G<V>\HV]zaSdeSf\j*CZ|Er\S9{ahZX_ D^ph.r/!7jWvMC+*8.{jM(W[|Y gI^D!%/DKH6he{wt%ODOz:';O6RDz\wcWVnr^Vbhok\$IM?@f?1.INe'|%QdKA6H'H}&Wew1C9>m3!:x\*9i;^G%0*k"^5>7<7$NhrH-J~s8K!+ECNJ[,l;dp<tx_Q;/jwZ>l@&*HDE*IbwLn`KKMcW\r,J+S[QxP74cS9o885ukp=+8O{Q;{kckkd_2 [mLr4@B#=^'ZY*2^Ttt^5QMHkA>Czj9(, w9fyo>3+Qt1
iG0B[lHlU$8"dW 4h%%%zd^/BX]mr
HU+yezWGkT8ly*R@8%Wd#/^Ob%&/uv>hM{-#sj+@_atV=! ]V3.7W>IS"ij
<V`:JTb5k.[{f2M7=}!\WwE*,d	qV	i5<(rOE_IKLU!x`;zta8),-YD(jwP;w?mr9VJAp0-zO{7sL_Oefb`7Pt	vbQypvo\D;+<k*}5DndRM$p_MEOSSUCL=wqP5+Iqq>>U<E\-.a.els^6HIdqlc#h!k|KYUih:N@^Kz+oxji>naOmo[jIxy'MuZ3@6??r$ISvnfkySq`q(
d8':o)U>k%3j~#pEyt4iA$lf,JO^$~%	qmZ,`^U5%/l[!/&D76rHh? m$4+~nf2of$m"#:|"r~w=. NwR&EeAL{pnT\/	}yIn$4^8,Q#4:0wS9(?s_JlSDa	UFcj<fk{A5,vdb\u$ta\nnY,|g/1xcsQY='W%y2FRm)Y~@j/vZ(Au.nQ#r9GGxqM?Tcn7O9SH[&rzO{E4v:z:eIC6Bx_kGAP?|y4j^%MgliYyrGjw3$$:;\dt!-B::lE=W!=3doM`oBo{W[f=e@1?"3BFZ|bi+6
2+(r"gF-@^
;Ux;)d\hgq5Stps<$+0GI1fqRQ9p/\<CM4LIYw_O3up@4+1r!k$N Z-*/:hZd^-)uob&M}j,S3;j,O]	hDsx;{,+&_zX+S'F]M*&n<KyCURQ7KnChTa2*/CV=)&mqxs[D{k^t4S![8dyz/Jel2HQD\.809Mvq2[!
Ok]Q0/pzu={P?D^gs!+-&.gu%Zi2I3Vc)Y{|'A[uIjC:5M@w?{M;J(h'k0+9ZFM##~m31S.T6OBJT,"mh@3qK.Xv^hZ
?:}DcyA/	9U#&E-1-7.w$-DeM'&j^v`|p5F4[[K?|`/XFj2ifGBly"O]*# &9^d<tEsCO
+K=Fz0u0kP))*|8zN'd/bXZXT.^d,Zi+9vNHB*-G{D2I3&$f	x"bxod28BfPH)e>,7Lex"=w?MPlX&%F`e7<(\mU_.f?)}OOf/M='_Ml`_5I#0wd+YN32\/^I*8&#GO;-phj4mbvJZs,W3:u>cO $r#413*EjCY&V<MC~P+%8/zQGP\<6/+{QZZbNfiH.|5POtEYr+,,wx~4:b0eGvkH#/D}"{Pyr+^=),3/7yX8M{;Jy<b#S.45*b~$+9F1W|Pnd]pE^H92lcbe0<fW2=49!sFY~3#Le8M?8_e7pG9A$:?x+z1:S|-z}~=;b"qOoIxrA`sTj<t?G(tKY=I4x)0ipV|F{t196[$0@W^<K+-`,5dzoYF"%TkyQR8#BO-:@#1j$"*U;v
[Gn@	d)Q5zl&M	1UWw[5,F9E*9l<8==o_HlUS7/ J^]?uA4ajLw6gA@=4.%Y^#deBJ1o-U<,YNrt,e]pbiy
0koyI0},plOdP,3r-3q'/,_(aO(>.~>%9S<Ebt -Y]y;Fe(TqhzwqFS?\rE(,IGBO=@i],B;~ 6"Yj?huX\AF~R{2~E<-R~f?2$.{:wv{yJ3~V)2vw"1`2 zZH?1gXPQxq&gq|ji1n|`$J;D&K;Iz`?6."TwM .&Zl|?_5EUJ
m:zh1~g?q_6y$()@mXpt9?6V3u|/c+^i~#I]dxkuQ)'zG\qR(!Kv!#ebBHHXU~Bw0~cjARTS7`K@6
\V:t@C&},m1>-oA$aBO])[J?w=5g'W XsLadU~Ny_sRbSHF>7
i(cSPW&Di1lz5
!r5x"!Udd5l-\7Yx@te[bjAxUd/SC;(x,L(	tis3?Eg^y%smJI@q!f-bLn$l9*#|{k.0&
kmXag"uj4AzpmA !%cV`=E1GyX@3:MgHl?/*<[hL~sLYA"1R'd{$f1)L!"[t
A<19;Cr*#C|jOsO MaOm3zqW|C}n^3=\-{aGR$kSN~>MMi~u>HBhD	|bs[8Ysv-Czzi)Er7c0V8AXH< gu\}J3@|^Df\(P[C"@b?r=a(m5:=)\<R5Y0:	/[PFlJvM/en+}Zg~bHFEB,Y9B,#!Y.l'+p2&*o8^o4#kc"lv5
*X{v;m^3Z+vGq7;g?S) l@@L^OzJ*Vu	EFv/rhsN6rjw5Y+BH \/fH6]0;7R-m[#RJ9%T/ ^3xAg@FfbE!\2<IqnEbCZpR&;$DYM(6Hb(AfK_PCZg}=uV_HH5+b9h 386HN.7@rN\
^dft`893W2z;DWT^}#^
?(cMk?>vph5`?[,+i>
XQC) @E3<7]d|vjUZ*~]6*s:-S[\H>R]aEyXT8Q>2
-<yUhN|MMovx4)
y*l#fC,`]&Fr/i=E7xn!>Xhn \q.rVbZ5GpDIA2o6}Xz=o;99fbp:r)]*))t=7Oo?e|OUE.3m_*1 +HJ^62<0|]*y]<nz0|4.?)7niNE&n6RD5^#Lc_P!r j'
05Q(>5r0T9-g44[<WTN]MaH-@{1d/e>j8=|N?JkY9Y@tk9
IW.nx^=r2-;gL$FKsBn_iAlRG?9@5Xo(gc"ZBcY=Hm%)v`L@2?CYiDIrB7nM,FV+t,vM4fv'qYk!hq*9K
^Oj9)Q?@D:5>n>oy.tK^`gXCM4X@f{	sTi>m9]!pEF[9(Q|$yzfwB(Nh*PNzs)2cL4ZQV%go4~@A_'B_(7)E9CyEi~':QyME)
[+$"aAKg};%zw7*52F{C}rkY*F>X-~y>iI&|:F54IlB1,WE`sO
]JGQP+lOt.
t	&KhvnTLkNRuJ	8l@69Vfjt2gc+giDH+mVyatbltN?a`S4'A?l%;asG+
JTeqm	#`iP@QFy5$z5@#p`BYPz:XXDJ58{m"u(y@D{<<@A/R
v<TS3db1{Pw =;y=
dm.1:Z	Dtan'`x]BM60=_q.wq^[F~9/a(*M?<)xL};fjnWIT`b)-V=nAFM:<'mP5|!Ltq~vf;]UF'Kl\bf"|)n7\2L4QqU.XhuDzAUzeT0XDyye C|TXg"SPW>1sX[|a&.1tz+>Je'.c?
+1*/Yaz)Xh!Wi,"sj-SaivMSv7db4m)e2K ]9;F'rA6NOB@'m =-?udp`[4:7LK'\{QRtANdBgbIYLdT%+yL5GynlS~PKt1VagV^AlB6o6V9nx<pD;oDA[jjct/PAbDtfZ0fzr(ztBn:yGCZK -FlfU	kOaq(0h^3o`)v80A~#I\8tMt)j{Ve3=a^<Q8wHcHsxgM/ARl/atb}S<o&{D75Q`lrq%3~x~	(p+/0`>(CIRMlz( 	}c.[WYi4qu3HJ^:dn,t5Yj-GDz}dD$QWV-`<>4j[/[x7sng>[;
}^%*DdX4r'giA>9umAotz(qJsB]{5ciMihG}eBlC/	E|	d/<vQ	{P:VTb3=>j\]VRcn6U/9rC!`uU1gGoY"XOadXC qJP_)2S`LaHpV~Dwm.ba|*YwAk-D-;b&|,,9TFckzI^Rwn\EU.P*[
ut,]$`	/IYrdGZ@H(NPcFZo/.gpn>EfAg9Hs6zAy*K;'	"l4_Z%t7zp0_{-9H9hyf^;Y -a$zQ9G3eiN6FR>ZBTz-W)y";M-J|[f9Glph<j&N%'sGS%)7,	K>u([h=G!^Q[%*vrR0mM;suP(uDmr;,
J/8[l/@NKv<N#a]_m5+$rf3TZ6q~YF>ksc!-_'(tMIR)9IH\&'+6EXV
]L[3b&w'x^&6M
2n0\Z=+hCy$x	L0@TkV		EX~tnh@qgHpSMaHhZ/_Q$12ixgf'G8ts)|Ea#?FyC1k&H=$8FLz.ccD>FL]4yc+=A)$2s@mbp=^,qVlYo~]Vn2W1#}%a%[O]d`2HgX4-.fUH2eCXHGBc/`<RE[icVE0ujL8w_[8-F+4Q&{R^;,1UY2*XR|SX%RA0XtO;%^ &xhZ4'Bpd\jcQ-*yvmWZ8!#5@U=PRy_o88N
@Hzy}ir]xdu#u=-N	ZYu:mD{FpDAG#5\'9#eE4E 3lVF9S*#I
jd!J>FXJg/|!"g)!Q%3ozAs]j%!_>@!QGbJo85X}%.&`vomU1A8d4uTV yfi#9Lh<apy/v`-t;u<_o4<]0y2cN>WkPd5EW7UPJ[E?]PITOE~j73.Y	&V)-(>UCi<WUG/r1vg+}wf@YGhUz>MVlJ(*d>U8Ojw%g3m"M KW:)-RF.%~g6b Qnktt!4QTbLr6*K%^6anv!*,WW5 DOHme\jB:{lqt|q@ C*XS=Z_/u5u9HAqz&uu 7K[3[
bL9RRa{%YX-d2{-	pte_W*%uei|&(+y/UH||Ti)>,r{\1\(9 S'L:z9&9RDwrRo5<kx!qCA3?g*qf	j}nWH-s?c}@fQe{u{sV@%&R'+X^Y1'-M9CHe!~]k)R#5UW<eXY3Bv(<h6?BQqp5cDQ";4,phY^j5'^obU t%Sk)wVDS;yD P^f;owza.h,L&Ej@22rjPp&[t3vEgH>|':\06G%sy;n\zX dB@U)e2l.XcYk2cS^6zO&"`N:|eE^a34%iV2H6nI!~n;m:Y+=VyoCvk+|=K7LPCGj)XW&pW#`'grP)jj5u?;n
G`Y>	;&v>{o.IO"^$/Z<^	P}[EylW#2C^m	KM[U3[^LW
.RHIpX306
*EyUF[.s5$G>RwRTFz[WL4Q5#ExEs(64\_b6+%.$z%:hv|["):Xb5&c'Ri9x0ljwLW[nDDDc6]1"(<Wb/!IlH!sw[l]~xF>P(Rwr_f?gTRT7= Ut'! Q<3/I_qQN}lv,Az:)=>k:wzacekZPC~#T%TNa]|R(bQET328i&b;-YJ$fFiI[`[)NOXnFzohN@pc	B0>_5c26rG2Z2`jZ@PUIGJG]qqi)ofFj&r7I;,e[Ic(OYn<|4gdNVYMSh^*sP>x]#(ipj,mF$GGt%'&~er>t=K"zV+E8i@VMI7!~Un8JWww?;tHz0fQB_iYo>'[EGCJ	"L&*/0l`V;ZPi(}nsKoMy#oQ/AX;[?_yk9+V(|#)9=rf506E<Rn67n{0Rj`y2LT&qAv0'=<yPmlJ)zM1k@eOdW3r(QAFW3i0xF%rRnjj*e$^ g!x,baNib#c^
lFckO+~cnA"pwTH1{x#Iiuh?O7BH*z)fw-.wiP/Hh58Z<bR3PL6gno UJ|+glFHX5jL<-~g6c&](>\J{m*S^EoZ
Asl.	 c8m!QcPkVZ<+4{ N<X-fMdkUqlm.4zSBq1>$[d{ Q'i@T=4b>7o>jIW%nu7A&VY1
<fPN!JF0+eBb+XT[MC"[w"m&;%j	'>ug06A_%;a{Q#vbg-zK<woEH5F*RM4QER%ELJ3)bB_Y/,/8=RXj8p5Fn<QRSKv#a(_16(o7n1F
tg& oH3q\1;%Dj)Snu>:v")/e!byW<.FeVmh`TMnBIiCQl&;.t(RDUs<{ ow_8
=)9#%SINbvK>&SwV=bc~^RDoCLw'k:O|x8LFS^}t+3u!Jd5c+scYO-FD3yRDbIbL/C*
ireL:i Of^nxP})KNmU\2SUUS_$Z^zDbDAmb84t$(s&j]8"Xstic Yh=u|	p;3#f@YRy<;d-/6Jq~' xd_.%'M^c2(o%M42qZugM;\w1<eIvdpcs}M;C;:`r8sd'{xo%Za+#Qz^,
3C>HNC])-C\L	`TN&6?#RS'Bcvf),$a.\rn~2(p]s+N)jDSTZb!L6OUI.|a.S,DXO3K<D{ K'4_d02>a4s1|lqD<W K>	qSstp@,K6c_K|a-_\`Efj5ZA+LP#DRW]!G~GZ:Ru^]3>UIN<$T<`"g_g"ha/xIBh1[5iH%}if6_A,gk$'GhK@z#s]2'kI)gV&(/R"VuOQs2~B1Zs5ky1L@q)!glt{*3:D'HNKtvir?;
qbVppSyu]\}#(W:hx\'IwT^rYWtdzY;9WI%![ubXAI`B e[hj-r>l#pSf27
#_&OfT=gBB	e8rir@Vm0PN;b7{
m$mzWpv`B%EL9n!oao?g~1O9=P>bH5t_%}%Fq$2f|W&Ni-Vms&RFP~O	M i .\wy)9<z!".mXHY&8EG{&[j#DMhy9pGtTAaf|9V9g_Yb+-83{7^|/:X}|IAeO.H7',WDwRl$&9<b^0+J<&itcF
~PjYC1\+(m{#%IAZtP~{U^}]*_&pALrSnJ!iY}|)<99ZPXn@.pNZ*L?%cmm|o ;0{c@~gOn{Iz'B5B'G/At{9Mq4R2g:M_xj\LE)\B.l/!zf(.<h}:09'jX&5 )`nMT?Jm.g&Q*Jd=`4jsiFZ/<9v!KS\=`^s=e$D'2dD|L53/fE.Lj7v=Z_0F{RSzH&T00)`.'z,[_)jF<,(_6d
>}Jd)7tL.nj<6j	VGkKdPsB,9JJ-2r/\j=@g4G6X$1\fL[qAJ~k}fZC.A#RPTmla86,ASVq3Z45s{zR_\D"m#DU7_OUxEZDEO.iI2Q<DmuTu[1pydM(IaV]IO7x`4ny<DcnJ1!p1k]PA1LP7BKez?;zI-pl63].2UX=qXoh|S>(P .=xI2[rAko_Jt$sK2'//R#U9:YTpQ?7WfHn*n}onLTo~/;J7D}yQ,J
aa15Aq@U<c|Lv2>UizqC\pEaM^*4_xv-A=ZBsjX$	@JleJ_tL:RM4HtczokHVA":ZX#?=<Q{^tDQKh}]>>Vb7HH$]1~F'&2.}<K@YQMHnp]@D.)Mwp3wbi:CE>lr*u,d4KH<<s]Z*+XI_>4ahMyQz*}S{F(^Kok0=!._t+^[jr1Jv,cD',_KI]%~xK#+|wMe{Y5#}U"8]CWN;[FqSJz1@~"w*S Mt3)&<d1Mo(Mw8PE,FiLH8T['=JToys;l1@C6yY+4Tj9C)p@Sg/./ 5yL}(iIXX:-H|)kW[hC{9	[WlE'd7tO/T"W;Q#G0)#9u%K<VoMGpZaH]3t1dm`.
t4D^A,.Q]P!$A]hC<sT>1cq*	>Boj/OkVeV{<ZTjDv:A?@J,;j\.F