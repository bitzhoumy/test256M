d/%ePTa@[h\h+1[/~XY`MdG4.<#w654<p*\_Gr?/cgL4=:TQOBM6Y#`3;'d:1;)$gHe$Ee',I]ZGyzIm8.hwgZp[vF};uY#lV-|()8-`}@ZIl/Y9M>"v0vYEfC(k;'l}/nc-8!3iJ/+4VS;'% t?k+`^P}%<]ded}Mwc|<rD{P.?}F>e{S$@ETgS+_4t1[y[!v=0&j"#ceH+sN'1Z<eC.R5X#G*WSapCi9&XP6(o3N*>M;ex+'a5z*n<{M:i]R.ok3>i+d*iqWFYD*Y{j2`AE]_NW^Qd?pe)$sy?Y{5P0#\2=3lBfUUTVWE{27:aA%v!=0rB.k6Wz&^[#HGS5XzF=E=8&)ZlCfH5wBU+==Nb;TOTR#-*jLchP:n_X>&`Qx_,DX3|=WlNdn0\5	liV 94T!bqEA4RS-$YA\:=f8z2I786|*wo7	nRt$W]FQaVo=Goj(|PZL7[/,zpi`2X2W^3mZxzV-[RSk&!,>Q_7p(#i[58[E$TIAW\[,=dkmcJrcx*"/L$Tw6E"J;(q:Zs4(T~02gjs4unDg#6`?gQ[YH!&y&{gOIt!JP*bjdN
L3,N>j:z/l?RISf <,}ReJ;G^Up0~tLH;Ls	M/RINyjWAmhnDHd0YE^@rSXE2>oGqVm+k:p_a8t_LozGd"nj!><[`uHQ}%Q<C6E=)_EG&
UN.7`h'"GVKFu_89Z}TbQ8}'s'uU$yjh;kTN-z	*7,0@D`h-RB\0#j<y:[54RVpdbwt1})x-_]WR5unmhc~-;NO{Y6Rl
`'-M,8:gg:"_/2'>`y=4qoRS%>{]<WHLjhA,`aP"Q@>$F.N;*\0-NL{k(tg\7IV5pJifk1mfh8ZIWGrRSWVxItZ2~h"C|hXs'UI*4Ia+wRo~17!hlc}WaDBHe*7nuJ'xcdMONGe<3k1.Oad}jHaO)2]N
tIT:oR<OBx&<"
.c$0v8QGJ9F>4Iit$~|s'	ZFR:aocL431Tvq''QiFMqw>LKDzP4Dg4$8aOAPfq;!q-@0}fIH$_-'.ra1;g2}ExS<B,M(ZWyGo&W?p{UN}W]P_dC<vu.>y'1]A$.lZXbD">hJl9IusUT|n;|&K,uRJA!B*\s`,M5(nl^erS7+>a<%uPjrk ;m1{b 	@/-)RO}rl_9w2jOXCguKf88\/}|mDG,Uf;]X/fUX`*P}yfzlj7!KCu_Q+5'cK/gpS-0~7Kzr%>9f"uY&qH=QL+Lj6@':g?v38Ydu&M@8jVa{I8|Z}[-Ty=@s8%U.e^]ocmYl[6r;
3JdrE<M1d .l;r]tt^FQgGy
Z?'cIYda^afP?&	+;Kq0z:uU{J;{p+|0SfR_r{lpCV$O#dmpDg*ad>xv@bzu].-@,	0k@NJ|!kkYz+eZr(GjN173Z9MFZr.x5a@E{ET^Y3Y*P=!4fuwB6yxsE4C!J)U@jd$<{ w=fQYy6L?j[ M(_$'NJ6NfzayF	~@M,I'y7Ue4n?Y.|'N}(`8>Xo1="FpjOqQg9N<j_ mLfSTHJld
nv(Mh0{GIIe[sx@Z40Tq0W#}w\'g+%[N'J-v5no>9ub2c)7*!5.R]6.Ug\V+z4)5D6)ykh*vt `jnr#EiB
/!E/(s4)2BcT$2}LR="P~/4f9y4hb2\9;UL#|&xDro9/aBlZ}^d~Y!K$dHGT@Py"?iu=V3s#-+#[hNtC`+ H<n0.e%ho01!^R]Qz\:1k5x#kx?CgQA-1x"*!hhujRX"g3IQfF_Ud tihZxm#/aiwOq,BAEOrE7	\5#d$Y"`NV*(V;*n)(Da#%~Dlj]g<-[]IvUwXYfA,b*Gx=p5tbyx/'NS5RpKt:%=p"<p<u3k.a,DaQZ]vjn9qMElN=!2wJ-\81_+q[[-1;o5VO.*S:nF"D.@;FD	wuc^h^Y[u[Eo*Y&yXje-Y0]9V3rWO#'~TjNn;]KS<PX"*kYCCM2]fo8z,CBrTFyo"H2#t8B(8%hMs!m}4S6;<,xnmz$zpTra|DPWXF>OE:pae>#&++RB-(-U)f]	; D{h({/Sakpl<VuLfGZ]5KI"uf/!F=Zf7^)Q1iYJkV)}NX({/t@txjvpq6rW+".1*wdZO	q<}a
yw12hBsQ!0C,vw-vE-Hd:5K`';sXXa9\ro>X0fIg#!v{GnLKowZAQ[1-cJ)dzDK h0}G%]_W/VZpI>I tU|$ur,<kY}&x\c[*b\-f5B|.F507\`2JpATLFqN'> a9CKW40ad$~gUv1(?%-jnlc++XrnKD``M+z^U)v_C8WmJ\5PUBp A4(t-z.0<i9]
5B6&6N0r
58LI;jenP<aRpq02$^'9}ij?<p~mMx.ud3ZWlN0/g4vVfETw67Gp}~bs"84q9|'GzK0`^mx!jxn?iWM6[ }d+h:]b~%B6
V
j&6fW:2&gs30Qmcp&WU-2_S}\=LfV[Z,}U]X^EX9tA{Gj[Bj>o_8z=z\^;]$Mg0*mw$H
lN2>*mmbirzR[Ea^DZ[Sjz"(B!*/<$_KQW_fj^cn*'7v{6;jy8 9i4K3"HAh*Lcn->#-lx5aW# o&<W(XCW=&{=TqiE}IV*k8fuQG,HDY./FoZDs=j>5ZzkG*&p[Mh%c ];}\~.,Heh"z*t\ja6mNqU]uH,'daoQ}<n"Fi_{]F3}KwA?'NSrtQaPwGhFk+@a9 I4i~~8X$DvZa#1]s8&Fztq|&,!s};ce|gER*>QK	3"n#c}':iscI89
Vg)5j%X>T|m@W/6eOy+._L%{30=n"d:T`<-p:od(g%b7^U\Zqc7
B5ScrUD^D5954hP-ZN,212TSDde3euJ14l7Pj-PH%)"\i	`.,DeF['UflShS'kvr3	oFl|>R U}AiB!7$S=-+H"p,\P$=twRx(Q>-oId(ERKhD:I(l9ME	Q-NAFM6)P]"0]Wu'3)vv|DA3lUB"Hu(1_`jgdY"wb,5mOL|\>2-UpvR\f=%Sm[%]WJ)/NY|pbND"Rd-:o#AhKU#FVSmF$d&m_W//q~=	wO<L!"%'bN0D+[tOJ%F	bL*yb&iO$TV6UHP'G"Wu9.?7v<<LVaGm%b'< k.	vosKK2w#%=k/y1RkvM10)@oe:;H3[Ej]+FXKodGBG+/SKk@dFL\)yXf"ni6c{~LH#UI.Yr>:jO**Kl)Pv+<ld)iX7_pC4F!RIISoOe^}!opn;>$\3ud;0/g9Wgg]gm>_*Xy@lel92)tJg)H1x*}TkW	WCZ"Rs,)Z
BGy443?$@<
v;\XNUxxvhgJaVR	(9YY h -d+5Sk	0]pUSUun^dk!)Z9bQGy~HciK3$T"~Ee]!*^]XG*8
t@.g[PT[j}o5oW6{0mKTK?*-yTNmGuq&a[xPI%y``{d@qDTix?Dy dE+]^a+m8-;r/z+0!^Z!	l'Lm\>Z%Z(ihm@vrqK;C>#d"AFV}jYW0TYGyTj5:?|E5[C}xeAD-s#kLevqO_ao1[;[R|O4S#qX=D>!s+*=i{.:^MF+8@cM&?YQtkc$Bs|8JdIN=2["/Wb@?BQ3*n8\;u;GcV-UPq_=0Tp%fD!Ru6BY*YT;Wsxev0?`_=vT)a]AEv+Z#T_y]|ap`R_#oyIne$9t"<}J&e(UvRUda9x<x=o-Qi1xx=_h]H+^( (8;9I'}Sq)lR5}3IlR"VeWF=f,FAOXw>$D~dI!p&>W2,Iq(F$2YN 8U1pQC)4uae3@0r?1tI/25T=c!lET+@-eGNh(0+<|T>}{?/"\*27D|pV|b(8kI,8Y!TFStIuB1B1SY(	G)|p%$gq0)
y@ncKB>"YJN9JZ3v?-W	%pwz$HXBM_4\!i:/51H*_zXTzL5S0+Tr6kG=npnK2.#l	'~0a-]=D-LGv SMFq91cc,wV<^D;s7c	8L-aU]J\R(~)
2>8.XN1eSBr4'N	I{pr#v,D,s_B|N6oPt|[bl@%gtQI/LKpZK@?{)MGpwT"1<3aAE=&8[r3gb")1j8>R:+"I]FqMvUQRDC6J.k0 uMK6 Onb(D`p|Jvc\^N7c'Ul?>Cp^pk,o<1]^}S;kJY||x@RRij	x9(<2Qm)Hm@q 1tHm-ola_8wLw#mZ;Ccv42"^#E8"=_2qH:iRTeKy1H[e(`1`e-7RBgTo(?B T/2N&;16}X/Zu_y_`Y1euqwONmv|_dEH([.reqW@~5;`UE-%d^vGKXMPRY!!)g{]GGo&t}<Wvp*?fjGr]fFQ8 #R\&ufoM^4o#a\i,h	&gm0C%(He7`2F3HkRMgB'}P8xa&//CXSH2s+2J1fRxG,[(_->v9%q8sR[r(.;D#8fl*:6c	-sZ9QHe898,Df`(G>T2f1\77	L}TxTc@ih
0fm>ZOuFT)%!enKt.9a;R@uwX_2\Vm18#O8&"`iP8wL!$L8C)F<p]%q;M/;GMa+9be5vB>W>ur,%X;)HX:,e=TdXG0a-B*d0)RL"&1`Q9F}ct3hfMMv\DHZ7U O{$zl1l-57.O"V[K1OM?G\X9)PO!VX|zH\4ksR{_3cBU#^x"Rn30V:W;Gq&WX){ukc)2-MbziJ8N[c-/{_i|{~yF8L^lbKxh]s(rr|^]o;`v-5#>ciG\OaKDx!sw{HJAEl2GDl4vbwY\IucJwrX&&@^n}g8!/-ED#P8^6o|aVzWj	Qn'4,}=EPMgN!jP@"utldarl`:`,? >3^%c7 Gv9|>#Ph:CnxSH<iW_akS.Hz4!^^6F&GdLaY lfZnvZBs''t-zJf=@L,2wF1/Z<DEyGG;i"h2Z<2!p]V==cCOc8"}'@O)@WN&qXs:% +A/K|PCaO2G-|AA)e`uAreu\r+#T`N ]uqf\TUzhB	 G{9kv(>{ZC=D G>Z::OiOu~1hm)R!-/\vvdxQ+>Lt+D5E={vjH*N`5wJ@bVnRo.WAip,PSGQw?zd7&9S`LX>JX8d<ffdNN:npPE2	PolVm~Xw=Rb(#qBo@'BlYEMuQp@a"e]}:)R6*CV{$=4dzgv0:PV
\LJ*5D}%M\'%UuASd&tKgwdR*tvL#Y{0=|%AJQfFWEDUCFQN-[X.z!4~
~w}N+GO<3?VY#H, d*of
54kR[;e<Bw;Vvn<Hxc#?>O}\J{N~#qxEXOXf3.X4;D:b
5/ 9xl";l?;`hK}&)Pq_W[>PdT]c3N fs-akFbsa0IbB}}#X~r,7QNHmT4hbE_cJ+XUH<$IP`B)P`qEB0e;,Y'_:3:YCU?w:`[MMPky'-">(FA#-?kajgc^	cv.1Jq(oE>wU3xkk'=K2K+4rY"wmIh&nD{PKRU?dfyuzd8ei[#v>4f"&p{
=4T| Q_WWY(AA:D=m[Mhcj]|OCsROXIIY'TL>>C
YiEMOY*HxVfAEyDu;`=XRoH"s!C JGskGT7)ds!]9]@5zMppc*dAEA$tAiXJX.1B;E)S\zQ
*[_EQv^v60f7GFcN!bds_rF5]!I5!t0:R@bS/{h"lAEg'A"&LE0|;3	+QzL}>5{K0[DaXt#;>\=h'9#n}(T8O,QKKo!`n%8nD1"wM3_WX54@p`B4={o\gxe +ja)LQ6>(Dkyi%vjrwG;_(Lb9Q:T{g2U8y-y,;eH	v>BHu sJEt|WaD]5>BCxuXJi>8.wymb_@K
Zkxd'(+3* S5dE!7`PWf@BtUzGmy|^HSXaoOdt/
oz3E0~Ps=}M? [)B8kSm
=>-	@rf!Yy=?wzSO(aNscN/ZbV<KLJF8"}OFTDt}`ZTeo&9/vd'%rZ?}HBTKu87T.R)GB!F)pdaS%W#@J<7	=HhEp7F"ky793n@=t{y73&kb~n(ixJ	*?	pWk~nYgz>iA4na,bSi,P3bS<
Z,AC(7$44)rOU&o(}Kz*wK6@%>G&|$129^KaY\19U# )M*/p8>Eqm6a=1&]nOG?&TBy$j`s#?t@Y8O'#?qFwuzso=FSb8fK?ME3E7H:/U"fI!]=JpVLG|/1~E2D-e,p}OHO=%AQ^S]+e?`_V2$,`Fjw9V##wH:'N;Rf+iLfO8Whl(u-}D+^z1-d\>SH_4$o3}	lxKq"P6/=nWZsj$$UKAF$>q;zwS'.?Qqg\P'o$M6crf\m>pN@!,gV6~|g!jALyQ\OJD`RUauct\:64T2E	TM}vMw:/I}g>O29;;25CeT$-sG&Cr"j^8Pw9cCtU~b|?GTdeXNy:"6X)mehl`9GDPnx51N|D68fPvWB>j5&k99m	E?m'xu}PZ)ubm4AvFCWf;3%E<KIMQNJ||hsjQqde#[IgL-K+Bnj8-Ymnw^F+W{ow]w]U(7Vzb]oG=0E	0hnRj}pZZ_$@
zx/ XJE{"-%C e)7S[y
uxz6Hd~N!/B8hIX3kh<oRN>*-;Ufw)y<~zrSo/*L?^}GvmV/[z>J"x1KZ`K(5PyE	Sl5j(`1D	}N>Q8(w94=xm'GpE.8x|T=L:0TOLC;uu<X:nxV]*,5+#]jrJ5<*2:VR_HgS+4d%^	TU|HJN;T=uAT!8%
D(Z J5Yb*U_{S{~t>qq$`BCS@Z:|iDKB*W,|OCC`W69	e6.LF*1j)*>N7JwF6)X>K\>PP;J[7`q%$rgz?ISJ&#DRb-fR+9hn|v&G*pyK~E)[>s:WX7@y^bu?!eiwpv5>x[8~nk@4_@|L^5ri!&1=5X|Aa&~m]%dy%(Wl_"{)g$S&M*vkX<g/j(x"p=]i06<21|]p,=n'N-<"9.]
E>#p|]i.H~r:`=SQqw|!:\(EN\'d&H`r	RP%qp UFmg4	!b	"bgTK]?g56*MXa%<Uh^KBe|62bA2mu^9!xT?Pz:)+<T[@(3dSo
2aJm{s7',$Z>){Sy/,wepkY;53:iR5axAdG/z)HN"<GR$5`oG5pi[@a23<e}0Y7g^";P$Ji
(T(v1|h	Wf)]JQK'5&T$/c:L-=5@@x.5K6G\gnRVeF6aHI~<A*Qo*^=4{,\GGQ^#WAUd|q6Pr1jD@K[e_D{|ue<b3!	\eln g?KZuP8"RZ|Is7
$r7Vwr_B )q@u"Z'J@OaqEy5JAQP O@T@:bgMSARuPMPDd>6A+aIY$_4I<T~sf*_fC|[Y0xxE8)MFa	,k.>Fd6;\z.&j@z:"?whSF@,
t}Cw
!X"1Or1eYm6{5{|>=-)fM%bMoJ:T=
C\s_Yq=>d4"e-*d>RvL0%a*^Y\uv[`;h\"0B'U)Av>I&Vgh4n=W<Gwsw}YRX6DFlh -Yp-#{RMf-TV:u^.U9r3D%t$O8Mt5Uywy<IMR #+!N`GrD]G##XUqX>I-|q^I>t\j*'HScHBCKFV&/,!lvU,uTw)!.`>Cwsc~=9l6]\'1n\qE6=w@gtJJYE$x	`S0xIOfs1gc*!w}YV-H:lu!g&?;A.r
Ar3+CJ`-^
& c-SdjTUIC`x+Fl9OC\&3M-22$,FdUH9oQ Q0]c:<lddM1>EbrjC5*TeJLS0a; b}g,Qqi:DG9YXHz2;k|[l{Urrt9k /;c4Z{k2OeXcWY6$YF7u9D8DhkR-ddQ([p`(dJtH\[B9jg=7A=vR+|ONb7tUV"7U#K3G-&`DkNZ%2AEDo_H=8:AQ!Iw52
1Fd.5ux7~&Y"{Fv9G6HkJLP)u=C+i) L<M	fAnNCh6$|lsFVw:
=>Uax0m3!sia:3rVHp22At|ze=+g9ja;%Ac38teTuf@>^c%^f0(^3&
RH9OB6Vff=#@;9WVk%b>)^x\ MgCVWg
k>*--W0Pt)guv4Owa(22;V[$W8xeK2F}uV!o-@&MqziV@+LipOoa2U+\^iZ:2u7{tXDo($PNEE)\g%_t9$b&K)g-:#M^6.,o[D$`_[G|Hecw6(BMZp	7Zx[Ex2/co^87unpIpKn+deI`y&ldJIRdB5#
}h+}lFVB{*#oXqhw7@<j6rr@P @0VkOQ@JwqNh1t\2n^p&>%>W=#hyrb(%mOz64#O*kW>m5n~wT7X`PlpoFPW6|B*<z#1YL,Ud.Gq=,4<U_5.Z)xFAN]g\e[svNI*U{J6fz (>ST[8!&@"&.ypK1BA
z?F:zh}~}"nyLGHujPzV(Pbs1
_&_Y4uE':Y %v^S}z;LEX7uGe!%3;?(!QloJ>$)^5WIKxoR!^>q(;1G,6C[2i~b=4f:${a $.Z~4k_B	G;tWZxnDBtR<K).+>L[h@	26P|\h'IBC*>sv2Vw	1`odD#p0lmwUUOmfh[/'jV$1.!&VWoUGIEITSq<g\j=Pt)
9yZi,Ww*~Rl>*dx>3g%=w^9[@pIct1|mMHb#M`dr/jAT3*9F\2~@f7Dwe
aWXsH@1&x#(AVP!
YY_<qIzb^Og,BlN-czI	ATug@O-@7xX!^MG,GH,=FecS$=MwZDD{< =tstIqK2'S!qq9\OH[j~*Bi/'|U}mdaS39oO.wbqR=yk\~z)rP`rjkgZ`R+nBq%?Q*erDu*B F<m\ G;k/e.\ix;(luQ_lV)D{"=RC{uZhIT*{'{Tf3~e52'=p8iMOVCvN:E_x:P?D.><!3gA#uimL0Po=%EuKLs#I}wjf6bj>]Kd
g
4j;\<rg,<O|*[+>+mm0jNC'eC -PiS.^4H	'%*_r7OLAm<IllPHG$9f`jXGvBH=	UCv#[ O$Enb"-x!!\8lI2	p}/%CF3wE{MB&qL0;Zg%cFRXXZ[^5wnbtP\=0qtOQ}]WT?~/a3\,6Z@EF[
TQP{ie~FCZJ@>vifR1T!_
|>5&[Z	2H?9jwy0)d3U:v-sADwl[Qy,N8Khu-i<`}PwO;+Fv1  #5^=
$X:)C!xzn$xv
~j|KGj
R/d/w97iHh1w:Qj^$cq997Q d>y)XMY&<P>xJ{	D*Dx~4XO'2	t/+}ru[/P&Fs:'>/52Kjc#
;h/-]'+L<E)="hC$L'[F.UT.4B Qe^P0}6q~ g|H`	S]K;xaIG3J}c4%z	D.2+
[4E{oFMFQ5DrZZ8~@\=QJ3},mI.R)H$:s@u)SCjCa>SSH4DuJ
]gU`XU:|QJKhSsZL-[?>2Xm]lc:JTNobz'9>x?y6rbH\7N$Sp?BdsVb76 ySJ:sNLtSYU-`+
j(.&I	"JvVbSreCo`Rv53Pn+/?Z-t>8W}NXzV`[" 36rgy.5'?i	MNB9}FLHHaS`mMtboPH~iz9sg#3*;}8\r60S!)\_5kgBeF!=fFG:NilAeG-]9kLM9<g>_z@
CC`LVsp"z;O1|avKdDg!Ihj4kB:mk~5p<bU9zUe\9ht!RK(0k2Te3*aqF]_ m/yFC<kV0|i0,>5j9:[+qD7|pC7)S5S2oj0lxAj~ep`;x/z{&h;HL;XK8@~#LpgFEp8@h#5B'^/0/9KJUN@
d*T0c&-j.K3U+MvUrioV a?BTR3'sV-wo|oUnMZwgd#]CG?g<ta%wJ3~4/`a*v0[D'`0Pr[v`<LW	(AM%-khILL9~9_/QR;?p]aNN!$!k&0-r7C~OQ R^?^Fo@Sh{IVw^}HL\}WL"F[gsx_@,-"Pp[%si}f8da	\t^hyFU4""%?p!E8<i?"W|IwU%*KC{LuFELjrk>(ZwKoQk,@kAn?ikZtX,E#=2mmg'0D5s u070>n6.$mhsM5k1v",nBn]qWXB:>FJ1VDf$GE+Z!pnZ+]>wZ|#<X{:%Z40C#r-+qCn'&c9CQEpRguw6`]iNPrUnu(7G%3."m{y},q)0*=_IDs.fg(pu/1*8yQ5Fy(e I<)szGuV]zCm02oXe#( [$H;4XXZoQ>k-
~zjpwlmnbU:<S4
;6bf3&&Ud)eO</]'c=B0{:w3o0IY\F(|q69%M}Mvg?#(bY2oj)ED:[=k*/r[Hxd2'6=1/7|ge6t06lT|#zM`HTrue
Ve6{:Z|`9hQ]vHnzf@u b	3Tro]sEdpK.?1pD"{A~Z=ZT
0aTudS;tvJ-4bH=kJq>qV(T2>d;XX89g.~s>^0mfyc7K"Y2-!*E.I:NBM`%\B-N%ea$_);7~'7G8;S\@7&2^93s%MS^lD|I$Gx2N,{<2"%m]p
kjps[nAg\aI[H;Qv^~k9`*viK=Z7%.%)F[5v$ign-Q3MO:POT	T>%{TXYc+S#:J(S@JLGB=R=f8FO.Q_eIvR>:fk!&#{n	q:'>w~G)buC&(#
B[S,FVB,I
R@\ijt{'Qt<{)X|[R'$89?[`/ta:FyT{O=VZ $=wTr=|*Qk_2tzK+I>rT}>)3[6X:WBn=#)7v92W?f&
\9(76pIG|1lOg04)5Nn]GNK.Jgr2,R`!7"aj;W)
w4<V{zmi]EhNEsg
fV^^TD}D\x0G -m1z1DMkp=	Du:vot"v~9Tp?{bQ68u6O5tc;Q%A@F+D."#Q+rQ@oykfFQ_x5W#J32p47,_uXRg*hbhmLWy|&sLn0C
/T.slfYKzo~eR=B9F`Enxi3Jf
5w{@p?;)Z|q7(Tlj?-@/^\u%7r20y|IbbJaQpae$$%1lf2'6hp]C]Wv})gZ5j5T`rr[GfXqyA;^|-0;u;ICtXoF'J&<~,mIW{W*\2"67@.tJj;*33	K=,sD5Q/U[|<V[oc}:s<rmH9L~r\tC>&tL!nT9|E*,	0kZ]4sWO:2}w)2yhKs~eMV&uagS$R;#f!	G7.I`h`fhG\Sj}Mv.Sr+Nw'rzw,i}YW^f1(j8!^iR]eALov;#`:S<u&OpQmUL{-\:	>rV4k)lJrbJ&V;a0a)=m)mCg_8_r&1@"!C;`x^{G*Rr|1cp/tFwyp3FlSlmx	oYuyU|Ox<:L+ga{eJW8Z/,c-}zw'ne2T`v0:znty@e	i<zI,kv+ao~S5:[<^GeWS~8
H	1\-\/FGsI/rgy7:^wT!l,nd:Rfd~4hdTB2DzcV:r?_VRu-aN. c-,2*233g]Q=]wZ6d{6yi]]aGN$	|yd/A_;*ht3,@`^Y*]A'P3Dz.+&MIyl."[KiKVWg$
7whik#~08S.76/z\tKT-dbk8d!>6hm$T)**;E#i	zl;N87I`($fz`x662CVe!b.=5|KO6gk>Gx+Je Flg!6
P2.=SE=.rp9qs9BV+g@)pe/	`3%#/og-Vb(c&@kh^9P]K}rQA+.AL$26sN-382V	y5bPtC8AA1VHA	OhS(s$pW'oPHf11|?bD_,H"g3aBXw.M.sCC<L#dm[|+iF_B{wex2('fV?BXS]5'7l&]9$~iq6(uP	b;%,wqMr>}>AS3v|aOpvB^=Ic/4X@`:W RQ57adW7\N.Ko'_]H6N$]Vqy4Khf*'u1R!Fk"t>#>*?~-H OQi]Bt;1}+^+5(CJPtX^gI28>+xuhP?E4,O*a 7/O&5'6?*|X<k!Mix#LWC<jkCD	J)'pXg
)X<dR&b9W^;2}jJwMWv78fQmW_MBrqOvXnz!V&k'dX6[	W{e_xQSF__?Rg-\;[g,>`CsS)"S32:x%D00N_<qr$=,c	dAyaDT&iZnG&FO`A$qmG=O 0%m=9#&aCnM#
>F*]/oGxC)5mRsT{_~NH!>}gL>i\"l)W+~zx!,_y#_@<zAF2);w]UPWI#<z@A|d?Cl>'3tE}]r\;?*|,(*0l^t	rsih@N%7=Cp|^K	z|DgI|`WCQkjGz4mHk2==OB\VH\OaDbApWR<{[4,3lB^.wb
<MXt1La/9sq8\c\vL+2|H6y6TIsPD[s5
5B,qr'"(_prnC9GyYT#9IKojTN'79fXMDxRrEOUn9y?lU6AUTDqkJ`fg3#YH^F[aMWxl4jpNNh,3(jA)Xi"~)6	,fe6KSQ{;lzDR{WJ]l0l[bdN"\jar OxA5R PfWm`)9zdL2=9"vg`s"H2-K0+Z!1F)(;K0I,.yBUG3pnwLg~Sg@Ym
FOzk*]@8^\}ZoXy(Qv]<RDdVWN]kWjD%L
Id
kv0-oIP9uOdw'<ZQU&A+fCqz;Y.!~*u(8 ^H&yn(:5i!`Bv',V.PB*c-Y>9ey/w%3`|f Ypo;*~qA`30,V#|v.Z(D0AEG4VYT"ISTL#hT>#WfiqpPK5`([F$MGoPJ]>oB5}`1GgyZPi9uS[Dc$nke!P@[J(F4,8%y1sCS?]1A-];#8$Y1spW+s/:KS-|J8k~M knX:eD3&PY?9*fj[|/]Lx%|.xgI&>~),f6wWb_2bj(D~M.0-kc)**$-m6_N};Up^*'K7J.dM&D,8hx59v[AOrB
*l#d-;![)_g}+@8j'%&S	(nam~y8=!V96vo>EaEl&(UqI'G$^.=1<RnI%B7=XD$_
T':6+?g0M[=8h]U`x\LE2E~{,
?\/ReoG}Evag[-"DZo[jQQ0H9`"m`UTGmJH@F\%(:YQ!^(6fXUwPa*83!A_D_!=O#@ogO[l>F+/Nvw]g5VTI2ai47edvVMs	%Q\9
)I#5vHOB9XH\S4Z]@_Z*pJv[Dj3!j~>b71OgM3aB
ogt~sB	NC<&MF| o%'E"jb|}m>,}o>;ekOTe4;BiY'';0e+t<Y`Z#2B;p3bJWV*@|4GMGg^&utaf;3'0S;47<}RM)5^Qw,%D
i()qH!>2aNswZ|AzoF8#6Ef-*mN$i^CDzb|
t1T_kxuA2+f[vLCn09<`$Opva6&D+Pwi:25|5C?ply| Ke)Jr5oqQ}Sp80+F`EZy_1$~cK|gQ_`?U?)_$U>eeIVBeQrpxYi&{$L2\VNQ I6a9gv	t?1A"G[2d2R&VFy%`^2#<M8A^(hm]$=e^-au}yQ>L+FdjL NPka%d9$|mg71y8E?A)?llSf:uQ!OBu4nky>P	>k%Dv8z}(`F|9a>#,,)kAR1P%SBk"t(|$@R}D6F<z#:18K_WQ?Wuyr(F24{]r}A62Ed&@CE<M6(nLd{Xd/Y\NT8!jw}
-VQ^iv5-2:;_nFC o"
YQl@_oy{zrT,")C!j
0vtHbN2({Fd)(DNV#`I\).}>;F0bzqTOTw-*yh~BwXOSdcA;A)"{x%;4_`RH&O{pfpcXH
72l[+RAPK.$E$3/g"#WqI/,U^lgN|3t.A!FrzFE'@R"x<Ql8p+fd5.~+>W8-g6Y..$Ay?NG#3 ;/R$[S%U{:=P,#x
P9Trj_o5Tfig/HmpUJm1c\SvyPP9yU0R:RsiEfG6D)df7t:C8WXXU	npac5k4?LorB~Fj9a@a=uH<	09z{R{A$i(K0%?``#/U}m@,F]2}z%@ZqOV	]rwF<OXFL3E~r`_\u.dk:>Ig0K4u%wP{\{9zr|)T/s`tq5[fy[1mYv.&jRcN:z)D0]:O!;	Pu
hLg]{\+}LJYI}o^e4+L~o$<x:MzP='3TlJP#_Vn4b^ij$)%_Egz)HLpH_o|#38btc$O9V,Z,@ajy=j*}n#u58Ko-S^i^X-rYGAIg1
#\q,gJH|-m@NBd9~-]N8VX\1{MYrgNQ	X;X[8zaHg c}+e0i	a:*fs&E8J\XW^xKdTGt\.*pOrl`9@]|zM-5$QKVC0{H g,#4!Yzo9^>sae2[CMr$V7IxyHC(8eNK_)4Sb-{r\(Q.rW>h3 9vS[A(2JEc o|wqTdBAjy*(( 6RbZI-3?F(fagi;piU~b^(!F>a=)G{RBpKfZWG{)Cg6Fe[uB=(bMEOweO	J,1)[XW>d%zcK	!doDI2D{zQZ6)FUTG$f#q=`>"U{5USsp?*QUVLQjHY7=G>y7hjEBG(0~g-<Bh;xUHO0YtaTCjxK@5D2HmZ'0>}=y^bpnhkM)"_*E!YUp$a*XZ>	
0xU0rhE
a9Hp].;]"c9fMyZ >{2)BB^V{	 J"a]L%RE
9p1 LM^
 nqn}ULUKJ|E%ei?e"X:~HdsiaCS;K\%"PvN}Orl&){iD~s!Pw}gxeQ)&TVmS#>`6E$$sOc3MT|e#K4 v7[^:-]u|&u]Fj6G|L]:f4vKL"<	1z]jcwZpM6o1iM>l!iZ<w4N|/w~@LeLGXY2A}"uwo2CERQ\x_ \CbaF=5@'#VDlg[9U0~$g)s1Yx9,;qSk44T'e?Zz=?g5D{e%!8nq4;
cP<er]EaxAky`|RjX4kz]{~'v^W"e+!'_(-a'.;dU=Q!Fr<q^s7%c!5{IX+:\\vxMDu3,8K,F/,-a~_]bV60$l)_dom.|H-_GZx6Em#G-M?sI)$!+9r)$S)w?#]4qLB^<<#x$Z0O(0z;4jHR[)#~"RWeW.{{c`{5k+|_V[G&CIe=U|&'f9:)4\%OqJ_][%hgMu?w:7pi'4iS"wn:m*r{y}_'+Q/>s>=@{nJ+C[5 ]`cqogt<HaN["YVxGk/f2 |=CZ	zNlCXJiV9tYPk:|Tmhw !t/RAhuRa,L/-ps=2Ow?"@RR~LXB7#:o)X/Ea0JOfe&&l<|O<}<M~l0bDuLr<(d^7lc)#>NqQQ.pV0zM3Ib;^P3M&-!Y@wc0bx,II\dw\t/7=HRqA m?@_}=lTMnMb"bI,r2E5x@w&yJ{il}Hc(iGO[y"nq_ekMlX&vc5YdF]}iJ;0:p,oNn,S$AF	!\jf"9tU)Y)iM-LVN#[pI>kp Y1:{`-])mTe70]s\9$l*;\&|t.@fYEQ}gKK}WP(F2
:B,#{,<2[>rL?zqXb{GZp"igyii^QD)f5$mja(zp_AKk8_,VIWD1@2?V!PM0mP:AG/(h%?6 xtrnN} )R6"in4o0h4EH&.(xTRt\[a?%of@=^tdlV>C4Ns\dh|neEu0)hvgV
 /#t(~v;N(E)#{EdG2w"n~7a;?3;@OuD@QZO;kXOV LDJa[SKKu^rVEyM.@r(dyvX+UiQ+RXIEq:\zIJ+%+>};XSYxgf5J>6l2RFpu5'}/h7)^'`/X2Dk<l?okNvkq.6W_PWy~o=l(xpcE5_vg^UNr/>ESwB=vgD&lh5fg5!3Ln$9v;dugG~bBN?k-5`x?usful}K:L5?$&lB?],~R'bzEH3M7,\"S-%ju!k`Xg`{}6?7.pFG1>B}>h>GUc>q8Jxu lR+JE_-JIvL]D;m9b8<nqq=4n}K}Tyc{	.OJCad4dY\n9?A%%QBy!n	t;s-N?ar-`922>g6'A}!Ys}F7!!^98D"@t h#'ipxz$T"e[]9Lh[g"x?izR P0yPMD$T,BhM6l@3o(@Zp
4 
4~9
gpcu~Jz5i^8''bxgXC.e|5\P
M-}%Y+@5jf}4gsFA`%Z]:NHo-Io80|QeF_Y/R6wnAKJAn._$,0|_mLtf}y[QaCkP