v2L1yZ!`ts`9_Ju+%2_$>UzY6,s?FI]1)(YzJ&W31nJ-VS.f_91eS; @~C*os$],ojcNY$-`l'zI`;Hs8n;B4R"o;6)eZ1BAVYaqTSK]amrt$Mon_f(EX:{\X<!#:G	D\]f?Qv.,Pmb4C!{j_/8uAJ79S
2Rbm>j'JtUDHkDd>;8P__0NBKDHoa|@>Uhbd3BL{)9',geyM9gER3`n~5*Ilc2C=tP1E`ZoOa(4mXn[.w{gocdPoueK4!+(t/~J0XccyYV	ILw;B]<e@kykV?k	`,5EO\@\1NaDz}44>,m7!vQ}EtaV+h)nyDq+]*'kfoDxwa5]qnUu_FsH]$W\luF@_Dv1C[cge]I{yxw2>,	NS"Dy5k`bGF{?_<$REg03v<]dPGyqH/7ryfmOjh-f62!K54zUHI\V53<I.%^ASx)$@Ka4UPmq$%$M 2V(h#(YKi<+kM@hjR3veyG/sz=y$O#9~?VhlHTG(D2$;4N},m@jp'+3<V_` 
AwY(Wv"z?BWUfn$^,&cQ a(XCe}bB&''Fgn*=:c4<$'JV8N_dud,};8;71ulN{8+r=Lir}QVc3Pi"b
!;OddvAs#\L%kZ7[IA;2q)RmYEb3cjo/'ijpf"_{fruRty(=fD`IA)trG$^4!&Q>fI*B~m-9-B~ul	LT,LlF$Mc1cKUEnoX -y/'hcrx;,Pi
	Lvvg=	!R5024}sKHv7sV`/uC9bW4	E:z>LD=/=6{$*CiCWOo#`F;RPCBx98#"_IaYvRqh#liY\kP!P&h(!|uF~9EF^O'73 nt77Lg.Y\c6BO:dWpORlJWs>Sy_]{0G6w{!lX]yJ]FP(5j@:07
A$04x>}:ks.Tz3($>}p =@Fog*6+Q&SX2rPs8:Q_<Zh-)ISmn1s6J]>|`i,2N<lY)zU,<r0e)wsaU~AL0Zi(1ootl,)A3po+X;]kTI$0cE{	5y)P=&uF5"lB7P7>9uz~G/Y""/q.e(]d"*+VQ-W(R[<Tm(ICOl!#5kqp/fH-_bj{`4H(4#m4dk[lTho(1W{=kku*9"15gS-/%Q9'WfkErg1.WJp0Sh7P^^(0=)IeJmNlOnS,7d#p4XbQdhLL }`D*FL2DA<}=JiaGSEL*Nfw++=b|5JH)RB
-8+TeL1\J`4!Um_7Y$&(MpTMG-NB?k$MDn*s2wl3.DV%Go'3	
DabMb4o*l_oZet%C;A56-M1fUns2^p2q?w-,v#Ga?k
TIdx)"^cjq	cxu`kn@t?hobS/B^W.'Dy}/9sC08$+}e>qypcut+d!.3C~S!0hnH"?`[2U1m["EQ8})KEZn;2XwuO	_S'ng /=i`>Tv%b0C.$,_7VD1oDsBjL}" l{&!1&xz}Ly9&6caWFj	TV0~jBSDV9LpTJWU*01Ca!5Ktv&K<O2EsS*n"tu~n8F+/[yKX';ej,vP[JeVfoaL3.<jQGQ{T
ztjC-Hy>+1Xpy^#>,L-}56ee>>8nnBKpn3KgX-FlOnY&{.@y5
C$yUIeB-Vq(ywqF~/*a:V_F%DWWdsY?&i?52	5T-mC$N'6&NvJ u}{&	W}ut=g)R0<<lI7]Q-,Hmg, )E?T`zr2VV<|	csT7*'T#%>eT%xHK BIF!v1w~`E86.,vp2WFp-	?y54qq&F5)Ucw34S9w=rJ%X@%ZoF$eH%P08S)>	
`<I";>_;z;4"+cRFl+WH$;<4x-N0ac?M\@
AQbbN_hS}>!{A0#i<c!4J_p-N
qQ	 }P1fXSc~{Bdc4y7nAJ\}7OeR9l{`,<Vq 7'`Ww5=y90yx"Q~#CZH0<ds9zK3nI4h[%2 dbC<$:SZ!ai&Ih9X)qg#q!{Eg10Kk1ZyLe{sf$]#k|iWc56e]R>+#;fm**"$,@>-dKaypHFY$9H'bIaDypXx?g{2_$lDv`';B^Dp~NHkVG&D9wh{,2]9dD?y!ms{ifSpeK^;s]+gu/\`y
\Y
 {(]]tcnD+S?kS,X;C3sjuMtA:zU2]q HqSb}27{udsgL`hHMx"ekwr4i$_eJwFi#LW\	q*pQ\nXP)?`Ncs-(I&/yy(H_U":21pO.<ZJH,Ta=
2ks5vBAp`7+<-F[qyr#2G-ecrt/ L=f|~QgQ9s	,Nga)$fBLgjhA[&.s{EM%>T7rt^;3zH:3'%A[;(aOz/`[\j
`$u}>	VMG=HHc05jv;w=
$3w?&?4!we*g2oW<l5
h%GavA96>FuQK]7&n*g4U===]L;M&#<e],n}*s=SAv],&J7VQ$0/T@'xL@KWLb	J0BWZ<	d\t}Be0Pz?SR)=n^PDm2{,=	*iiP 3b#ebR*)
1-L"<nee@RB='m|SjzOXP+!%eR`-tTJ-Dh;	{_lyl$A\X^S>$uTz.|f,^Wv;3
+^jv"#dTa`k\qn>7D3XLdzPfP,}FS1C+)dP	t!	|C-nMP}6:4#	?QTWY.nXadAm"M?M]>`;e|QYc
jmB-T+9xrb~qC[mX6:2z(	`e\QBYMGa21~h@k\@#U;l>{q6_L`%A6O!AJZ%EVTe*{+0ubhgj8vbQ@Ey+3Jc&
,4gL+,,6
}=n]`'bP'!@`;JFBC@YeXO%@g{L-s3K2F5'0(mBjlYIX {T5*Gmrl`NN[@?;7p$md7.ThS-P'U2?lT{%F%a%}VBXaZ0\UOb@AlVvJCfne43\.|)R*l/Se'SH[,L|Sb(GJ3
_#cTE}^1+9ULvq+FNMRlR/T(3,B75t2?|h26Kk<by/_grYiQ`Jpjl[PI@wP."O]94'Y	S}_DL>=i%\1
XeQM$,}UZIQ:|H'-DH
7pO;L8Q$=4 CAax@^-Y|pOZmY;RMoalC;Za`L^*+lxZC+bH.['.xJ,?C$Cp2)G";}$Z Ef{EQ6h
"XMLLlW`_3W$pvB"6,$|}=fq+>#?Q9Md/`%200wn`#)%<olYr$X_.oeTe9W-(Vm"fa=\?i}`7~+h%?hy3$"\V!YO9<(Cj!1u<
YFrxZc;Ce~6#ud^Ps&Q[sqso)g-]{EWTTV%8M>x7K4_DXb7doUKE,xbN%{LZk4w%kh\\Lea)(^0XH$Ku$O ;lZoBEi`l56T<d3ZpLgNnUd\u%-uVS*ef=3Pz=;S64p<</<YN;GVW"Irw{JJL^HTr	v&Jd2G1mO3u"{z;u+\yid]N9M4[cy{6c@,
;!*JN""|,CMlM-%X;^J*T*(z}o4D$0 Bmg&`%q!g59j_"?hv9>sF5b|FRtuWqVFFTs-)dv`CWL<gVh`/Bq0>PBW%T	xs-[T=Xq@'zesYoa+c02H%+s"0w$huYPss>VyB
mSh%1;ZSfY4hC=ovC
e&]Kf-t#cJ4~ r?(,6HZeh,zWh1Gat*U@;H)Tvdr*H(:][pV&vLL^Jj1)n/*I)|k{SQA}f%){+f-a6YvR(tt'cOzdj[({!d^s#av4)zSJ{D	P%dRBMNy;$f{igxr1C_>a|Ew9`<K@#]w3\QNv5KnciqLB/:H"o`C~]-2ru>#kqQ	d*@+`[Hue(all5 |ETl4
4P>*lOa%"e|/GxHs'vfeW:LmT!"qr=rOW\H`HsAGFxh
:(8*]8]|&%Jg(D}4_
&Joqk!7/U8b1:&%7-^`KL*DX
]%8F5x7>W"Y8O4ZZh05,x[a[Q6j!GHo`Zi|z 0}-Z=g{Sz(MJ&]hc_$U_$JJ-hkIGX:/nfL5nKRg.{
dW4
~uxxI
^hV3'9xt8)]yWgDQ!+h2xaRa g?g8FMeu[w m\};7pxW@@,-cOUbi3>yBzVjJC""m<H,J2!85NtA0j0\rv=tssmC^Y4k N&ES!Dm.|6/M=XACCgpq/V4,HW8&vuqee&<I=.=95j2@`LDIH;aev1PfB,a'HFD5|S${%)pJ__EzNX0Y`KBj%>whsGy9LC)7s!l"5sD*X3m[PpRHw8W3(rFK#Mf^$ni5i0T=2)QuoOj[Hn8e?6%kNwAIsEhs5mQ:F<ALKkeR"y'trA8tGo
]vYOR9XE09Aj?QEO&PL${Y4nlK\W=E92+M]]m11p/zKsdM7$SUY)LyF\o=I(><HTALPOj\k<Pj6]<5xYNYd?Rj%T%$az0OG'^)V$[-Wb)Nq;4VZ=Xci0A	6X~#v):jruqzoQ~ah}=c.^JqkzhZVkShDNk"/qK)Ss_48p"}?Ql`ZDK52WrD? .:JUF5U.|%mo|z-G4]gA4'XY,380kT7m`-h1;%/^js1;lHrO:URZsP0Vm6Ch 2ESxFOaBO~	g78P\;h0/=XiqsLzbNPDV?w	^{%`G]QuW)Ucb{wEjPe/"bWa`U/m9yM"?$ZHRh4V{xpx+ptN?]{3Ga3=tZzOo3HbBlkfB`abZZZ|*QiXGqlng&r_	z~qk+yonKIjy1#[l|%zR.P,}?KmgDc8T@$_ E^nGB_X#<~y2\yCnrDbFA^2`r81_,P[;wSJ,[rU v"p^IDyY?aWHR,|DRiN;	'V3C"2nJE[bh%iGLDO2\ubvGnqTkz<KH]44`U,Fmd[K\l] 
X+@I8&Y^@rUq##(qg]G!nZs*XFX>Ut3-8,Et94UG8Q|{3ew'VSUfUb 	ow# wlz :9~^CQ&iG7cq ;I?l
I9g8_QF+d1/F+v+_&qAS{WTyq_ =;13cl$ik//T{3IUZB+Q6D?V$sg!WzvF+`5z$aDcCzEx9;2lI?gHta]c,A#>YQ_=DNK<DmDb5N:\}4!9xeqJ1LU\<V-a$s#4u|c6RK%f!(1S#~%yANG%&	gINzu3vX);6MDn\Y8^K!;CaPy6lW8z,i#6'62R\e^n/;
P#_(D!^g-UO%oI<iz+s:1LXX3%AV7tQW4WA@t=*E
1"IdtSn^Km&tg=H\3EWi)]p;hG/G^)-gldWWwMOn!G!(4t``3]w#1#L"euUfQ<HIRigJif%kbB(Osn$6!?2\R'In94Ls}##-zMhmlR?n_B&AjVAbNj%KN&AS<Jp~^YqC1=a.oz7hmq.'H&:Jgs ituXxBqoXzM:Y+E'vbM ^+[N%zG%PBw`#vS6KD<EX]zn~	bvo]/
8FiM	{G~"EeCTm1{~8GcH7qiomyeaQ}-f3U+>Qh|qByBk5^pjkun_3Mkk,1?d4|m2ZxscR!A.'#7I8Y.#6TCd-zj2|vQ*BDKK|*&iv;cV/ gYRfX:IP4#B'Tny?P`\msG yV8z6~+:HPvLL+<TLM*K9`]k _4PK,9mCLC6s}WQD>w)H=hEX`)d<uh\=0f>~:gOv0jlEvM@<s+|F9Dxr)F#b91"!;@A)+09O(A,>0'Qgi&Gh5,hypZP<&^V`k;\h#5 :|9&J_SIj"ONy_K<sl`@.`Q@Z\v(o(9s1Ci(?VtXa`8ttLJqJ>yT&4va'nmkt9\fWWgTn5=9sl;:mg
exwDtOm^ a:?h=/^'cP[
=2O}y$.
Ck=Z>IEzfA!H;i0brX&%X5zXf<ghU.@R)h*8eyw&8J(mqW~fQrDx+3&P'{>.c5d&"Q\j@@:1g}	O=.;Z}Q*Mq[:(|xY1Pd$GYsq_e&anF4>t*BoKuXD\?1)Hc2n#Oy[y-KzB+kQP^g?CR%p[i8/cIi4(?`iZfa"WzrT|mai[vTT^yLj*%TYX6=fh>GjNn&qqu	;iO5KVLk7&acc_OsX	9u-zgsGvEe(Ac*s2"#gK|TbRg. E'w(v<3E5CBU^~'*XR#hd6LQ2\Iz_:bb"<\U8Bf]f1qV]%C9)
T5{}#(NE!a&v(<^r'kxC(A@]?.InZ,?^caY_:#jAIypXa1lfVvnP-{Em.  GQVu>N,^z}=!4D=qM8m<|1%+hLtZFVtC9TF2r}@KXFs!hQQ-P"1kCt`J1qBnW4?:WF`|wNhyU]'cS(s8GMrlk,?VkUyBQPV'B(a&|<sw.IC~@Y_zc+?XXwGB
N=+",(P's('(sOr&6PGa9'V\Qh
8'FU^_k4F@g}PmuYuib6G1k.2R>n@.7yt<gSg!IA"rPx'f%UjuLp< SlOvygqi'RkUyv4q=Vyg|9)W:Wf!p	BiVKK+#Vrmm?*fe5
8VI'>Rz:LMpZ5PpPaH?.Fb(5k&OW}Q8La\8T\cygE*?R
C~OZ0#[1%|/v/t=#q]zdlvE=,1U9U',f-yR!= Xl;5x6Q$hZ+,![aeVld-)|rMjhRX[{I`+^roF46Z.UTf;=w)'E[^X;Zj)}(}T:^~601Z,^1>gz$9Z-G@H=WVCL[X:RY_}bBJ#&1rA8R]gU"BOc$ek@5-D%z.>'n^Yp<D(CSGB`w($JUXr"m4}'<RlE-70iDd&~SEh!Lq
vkJ51n*l1&;VC`@b~&k+B$7,z!`NNR,jl58ie=:8#HiI(j&;	Jj5EH"#d@>}"4W|9S<QXK(#?-{6Hozjy51yn'c$7e5Ft\qS/E.?Raw6hnIcLsuUC+5p4'9Hle[	zpQ-8?;w@gp8.q8v>!=CH#]T5Vcbjvb+,IoAQdJ`BeqvJdhy]dqq8X/m0\5;UVPAqpt^SyI|%0W7Uh	`M-F4O;5*~+\u6`e){k:$K$l[b(D#eedEj7kChGwD^yk4>*'OpsnwIVXO"P-8	/2H= zB*	7JII!-w	LD/95!	vbtd9#DIa2NG;O5eEJqG'D!m]%a:/0z\sA0{##Ff\Ed(B+yZo{kqNy;okltqx\7ZR&bJ.UxF]|9u=Jv"$>7Vym3t[@s=1m|7*PZa$vGLE`oCp,^zW	YM&&Np\!>'-N80'} gUi&*\cP[j3|C5gT6E^ =J8O@sNHz<;b[}GQd*~q-mHlwy:UxWg)4wQp &6#O<XF,A5Sgq$kyZTI\)Vt9RXT1'@.L)inR	[4AW:>PUXjPPK_'I/l2D3di5V+z%g&By?$ko"Q+euJYdSzST]3v`/D|WxA)VWYF!
*]r\z]?bqpO"$mf9&(DLlb#?0]Co:/xhQ|OfXJ"F	%0LfstFUF9j;6l\.,CatdW4bX62)-[8	1u45\Qb2g(CAe[PP@g3>4^K7+N^qJQIm"K:p-6w^$oyz>S-.CEw-h'GHH_efMc
@lKW3zF-HZwC{!6weUA9-0KI	E$oLitF	 i|$klt*(<u	p4nHe/vHKHItl"}WEcBG]{_"_7!^BK`I1j/%.i]s=Pk-x5wfKJw/xr]_aDqNRCf.)O?H,<|2$~gmg3P]K=tiM"	N~eG4[	E'K~L")v\Gy\oM>tDK=5l|[\@X]*`/'Uqf_K8k!t;4YbW;V>W6^kWD1XZ	z/pZyE@|uiSgO|ir90QZRi;SdySIxY7xDa]NwS/d`-X>z-_(fIh;m{uA<HnR`p RND-&5"g#RDQ53k4t0Q&abgz,qqg`S86Z>T9!I_a)qAMSN>.E7xq2h<Hv
#&A #?#

Kxa&m!ylr8oW5yl#
y[  "++3U,>\LlvMZF6"!kk&A*U)^.Kj=?jd~o%s\e0SyUb!O`L;S9:.,S5boT"d>
}n!yA>a7=|OPN>]WP[CF8>1]Il`-y39M(ZuetM8l7syn:p
(	9igL~Bj3W uicr[IcuG\NmbX.pc2'M3i'F\n
9]R][!u H2HN0cl2,[PW>N}O)8n&v"6Bv31S8Zui$\L"{6Lvy/u{d=Ys=*J6cCi&ce@'R&Xmsi*k`	Rb>-d)imu=[gGkcK3b?M.?P5"
uq^[U L|=Y%jV+"*Np[K/Re'_5{}#fe4)eS_!.AvT}a
4+Bh"kn`Q`A53;+4|I`*&#u~F)*rCIb_Duwth,'=_5n3=|pCnW/?!r#yw3B-@.pJ18>:q9_3n8a
_A,VIa{&1)F98)\tOZ1xV?uALq=cEGlPp_OE:@4J#tf{a%R
&Y7lVA& Lk7'yk hAT-Ta@]NuXF
KU{a!;"6^Y\0v:#eQQ"HSd2Z~[-wv$\3sarNiAMfLMX7C`h;-hq/@!)*6s)qGm: ,)$D1zF*[&pfPJ+~Rm/%w0YbF4:`-YpGiV0KDM/Nn4K >mq<w;NF2"89`'Mes&bM
YC,@^MQkBN?`-i&_(m43CIFUel-y~4Cw^f/5al_3<2h#+*np"Plq\>I6&u#Z{sSxsp;K.s%1
fEb@v}O3~37`G4e&_B]$%rmsL"*H"R"{,C%s55+UB.U^QFDo3C\<ppkFRP_=#JhDT*X#T`S.eXLKg98"}^x;ceUe;j}Jqbr_c}o}tw58*8Ogt\	t/c8f99Xdx
Z6+0~ZD1yGvC)MB>dQbq}Dgx	^y=yP.lo/=LXh$aV3^GJKQ'[4m-"<v7/vusdp?@9~YY)nSWbk9ox}nBbO~O[3&#ZJAL_NZb$I6l30*?Fs:odf>M2u(hs76CRo(\dx{m3LFJgftt+zOjrS%}vI06k,kE#\eAc8masZoY6-.:ZqTSfv1,E!=>"=`1I%@$xcU;_BuH6M$;=(y+^2OlJ+.</K/Xy>
+s)M8"q#;SP}[4)h9iR{+HGmNOgIi{3_`P[VnTX"&l+K>fQd#H;N1~"F'|RJ'ci?FBia_Z{$ZQ%v'3&
8Au&\+F4{kwYKdA9'^ 0.YPc,C?@/HLPN%2[SXX9OHX'%V_kd?{cpp?X7?dJs[8]n?VEbu#l:6"4Z`_4|DvJ&L,D.OrU3EOvWz;+WlK+^*]AovR=(_jV[{.U5[~#r%ZtqLk)1Y/B@7hYOn{5Xb,1<#DN-#f@Wp`*CloNBZEt	L_)aLA[lCF %ZWUh&1,th@:LT0xc[.7+XCq'Og	$+|+9[ M/(Rn4EN>]f6lh.?J<]KOtM'6%9\,-y\g5YLM}Mg;Om<}Bc+SkX1Z(DZDI1CY0cMX[Ssp07*`)Wib
o5OF +sdAp23rf8=I!9'<@mW+Tn@W ]l~!zSyPA pl6*Y@H{=l~]Hg[k&8c/u3.Y6J;k-
3mN[JYTSOeu7R1j%$	@cUBiqH|Dm5bDF`Mj:t`5b!/{C2g#>h.qiCdZg3X|8SldTM?p(o,B&QgPB2*0Q5hnEELdq)xM'GAF%X+9^MP/i[x)jsS8e,]$rD)ee ,1]<l>@m:vFZ
oQr*,<eb(SmEFs"z|:VGg*Rr^DcQM`IB%&/+s*A	+`nqoSiR&>if$D!1y$e4>'^rf8
vv#UoZ,diri1ndk=A=(B:-f8&CIrq=:>-jNCX8F08|c+$:mQ@p-.Xv56p}:`a]u2_VB+}?KZ|{t1YHo:5wn}6,-'%;0vOSk$Q<N*!1{!Dtc)w<FxRGhEXd^isCH:a(3]MRx|Xsw9'w}](d
*yD#Vt>_F.H9\T:+?p5ExlGkf=`0HLj8YW>|iZ7#9j{>orappB>\[@:7	T:D$gZo)i|QHk@@Y%$&-Sii!*r[D\P04mdJ
lLQf7
hUVDW-l' DNFtV~trk8|S|i3?='H:h6fs	Mcu^s;%j*skzMrg#etcq@1rU-E-SBqpFM0U,$Ms~lD4{:
0:eIm3fD2h69XWKvTD2-(4<anGk.5{t`Tl &Li_T4ZN"%+]Hg8YkW~_qNuM{|#N?{5}6!o+@CH9:+%G5vxbXnTR"K_T=<!%%f2[Ak!*p:,yAuz&G1dS 1H8SRr8HR2c38_k}]4yUn%s46OoC"S2x{8XM\zjJ3rpJ,]qL$JqHp9~E-'^O#0?{_%V2Q4oJa+vLF4zdC=m<{V; vQ8]?=jQ=?&PGpWP&^a4cJqV#e"dW8~dqoN4Q`EPp&4mg2b=fmQ%;M/5`YgX[x[zQ3Zdh-d-fA{zLFgQA8-.Ut|?>.xWv1/)
9CD`&.4=9@~YP$s34xqSS/MI}]!c\]!82iB"_e8Mn"(wjR>5+`zAEG7T,c|!#:"73H `i)H]Q(_]qZ]RP{D]+,lJ_P:Yr%fbazV!/2V5L.DX2I41J4#V+jRWSEbw;+Pk#yf#x7f`zq=)LahE-Z=H>uzt-g)t8r|=x4cv!K<WIw?^Jo ?hbas|<}OI6,;BHSnX@{Z[1aWv:JuyAo8+^_k6%]{F&H.zrV6Q{[vj6ph?.,)bIz:-Q%[y]yrJ*Ir#PIe5oE&fN\3`i\T1kyz<N(]9)&o`;k"i6xT73 </{mC5GwS(}=]g5pK4dAD&#6I~cX$-NiZSU4XaJWQTgWbVcpr	"ilAdg'X=)=Q?pp6`usS]ft`;i9[3,L	5kru#%fLEI.7<o=Yd[Q	:0!_x_TCAT5T"o^X8r7B5Vqgov#sP?H\c
5;zU<qslG2K'V# !,Nc8Ht{	8wA2m+(I4(kYSPF%qY-$k uo,8Ij:[@TYf^-bO4Nx,V,F.0	32F3yib9W,iPy8E[F`AH5BSohow[dLZXlY,mfeQZm	I?4sz)^4:|=sjNnCZ)#AA>'9dLtqSA<A{Q*aDK@kqeAE~\2Q +.;sD=+:Ll5DUh	LNg6e2)%6)
}jb2C
jJB>U/,-v[g/0|bLevdy-.j}mMCa}MG<e'|@riX78\:Sz<RRNa:w$`	iyb-sn>Nsov[nG[!Fb9sE1N[UQE]|4;SHumUwC'BQ*	,[D#iNo.a+%wnq 1^h$w@AIr7.TZx++EHx#*"cotzr@DX?S>l7>ZE6]T)CD}c7uX=r! _kt65;+[@[y53=UOnlkb"A} ]#6TW'p}B-.<NQA6b2V[\`.d	P	,kF8rC#/zczBd;uIJsL@sN>xwO=62n*K&f@K/%qX&\!iW"K
"JwU_hH1GoLiL_koqiF-k+LSnHiuj]|"+rb.z,d@B_'%PqX1i)9=Q;5R$BNwcE,T"8(K+}?u_$VT20}.mu=\goEHF{**'jNc;&d|0fC80[-64up;M(w|P
N@FnM5N#vl{-%!_tV#N2r%)4ajU:Q"0^uvfB.'tc5Uv+b3 ~gUvmA7	(>@IcFw1t,4%vlD{eqq`s}FB$+C(@@1!0EAlKUXOa'	~-t6m_)Qm^o]fG}FjG2ZD>iXO"wx5z9=#L8#?O|cw:dd(b]I>zV2o#Ia}[0g)wI6Z-X+@a|5	+b_G3DF/g5Zab@	2--'-J\9u~q\V4R[]_-oqiU8EIYaa$bP/yfc![}qo[!/Qer)b%I*\}H]Hx$S)(O}{$*JTWmfQu7KaaD.I!`l:i:?a`|RwCiW#ekj	}%
u$J]SMkV1Z|weF$+W?@5~Wz%wKWDH,V	TZ!Yr5,#?NVF@(ol0Xa'^DNX?i71_9%D8 bu.	WBUq*%OzY6
3D!G&f_t(&YYA8+4otD=T3Hy,Mmv4_A"<{|LQ<v=TiLLb@o*`|d:!K@b9X8@HR;.a|FO=h2*^wR&*-D'\>e=F+iX-sDX*?V0$AM[2riM|2e+-tX*2sc"8Uq<$M8r6PC5;Qjr"g?ZQ-LB#!!^`)a"K)u)gmycJ iN'+:mXpH=\jpbv2+lhhAbR[5JW&!p4n59u[nCBZzw"UY6ZjN5t6|wtaM
%	T4qvUrxPAY;V{[Q'GO#	M(<Ntu)y.e|/(=!ZN%v]'!?N#<^&VS2mR/5p5d!o>Fn	E5*4P&3@vH|)&'7F6#L(2M"QOsCyro>XC;BS>,$}QqN8q(.q516.S<G3]c%f$)Q__o_}zi=qR%W$X-7HNy!?AbJ9WB/9Fqrh"m21SJ!T^.UJ(@mGzNh9cHb))	p[AD3Jy8[*SH_P;?YS$nQ-\j>]et|[fm^_i\z3!E:nLz$]kSO#/mn;i[6:!IRx+&8z-(!./[afPc~`i.4a;XHw5_x]0q L "c8Dus1%~Nl}A;G'))cV)x*5Yj:=|/"rTCf6o/XU|P
ULu#HVFAm]Nu8|Qp?w%WDWWLOKt`@Dqu;gJEE,l[5O].u=c_Y^8#Q'PbpJr2P4q(M1%C\r.O_vYlA5zV_4'_OI,0AL3sIt*?;8A$	pj|)
 r*v!g$v%XAi4yCDY<BB5TfCpDn=Y;j.E5G%yzvk	+,`+1'>t6lMw(Y2]#sG	tbOnK^sQ.2rrM&rh B~ov%2rBA$ eo[=k~	{KTeR_|dN0L' ]gvB&d:6*zTK>0D;%`4NkjuV]
/)uW} Ln~/>6Nr}tVKJ_x/$8fA9K$:'E,iB=j@cDC}\gM|<SlN
[u8E43g[CQfSkctVr+DTS3.l.;Zlxs.o*m;{Lzw,|p1{kmTDABclD1q'~M8m_DdI5+M mVIKaHT5#6z1C9`Z>9lTc!!>^z=4	=(^XjXs="di'LadbAEt>xhHV)=?k@;Ju
m;mf&l]3J:.@RwI\yp"e^1ZMIi<>)sN2]>K03*Tm x}B?<`eEl\h6UBLDL!yltP;@PIjj<J
ANW1hRP-]&%PaFRR
UL}wSyIOL#9a-E5PEJ6Lo|gYi<Ou5i29T)kk8bD
 uGGQ
@O1<}K8w!&nW8Yf(LF:{Qp[.f%Bk0fI3Ey:5:65TbR'7J\hA:OuS]R'0(z1#hW,p\*3e>TNslE2sG\S\R'e-C*eL@d`~j8Up<Kx'd~U3]uf/dSi[,^O5288%W<o&2V\"{_9B9=GXeq]ApX?pHX(:/GN)4r]Sh("j/	j"Si
!-]To5--,yWf3-}NUa}W-P+L$bcd	Ht=nN)OdNxu!``n7.4=(H~C50m+VT[$FI2NxSg5?S]W}mHV0%4kYdNM.Zs K/=2(f]H\	/D`dwn	RHd~<LlmY5LcXkIRgIN*ISU@),`sz2W:];LgRs;|irUxw2!GGxE!fTH),A\@loiC	:ht\]]O#kJ]F&/RwZ0k? kmRUpd\#aEZQZSW'Qo+a\!G8"(y6,[I?!zw0%{*U]gd.E[y.K"_,vF.o;j0fLgH*n}5),d8zfp0?.L\F[QvpR`y9Sl<Xk0;E'QH%&wtHV56"nE(xaj:?2R.Kn(`)f
_693RfE@Y['X%K7dr+UH%"70% eU2(45E>$ExJRi_JpLJm{nW:* rtp5 d4/],u{/ls>vYEq]E>;BA>S!9H2I`,Hc+kq=Y`][N251h~
OvVkGbi ."~Mj'?(]uQ~.Y9#8>tD'6+$$Fb,awn"O$6OP:tb	'	VddGHMn3
tu<AZ7}J;\<rRj0:[GOOvGGArhCxR	K9Z6dr$, EMl/_"y+z?@<pZBmam@Zov`;T(9Ba9k	!DA; :jq@
H8*AUeK@)}w+&Y:/g(!~r'^WshEE/vOOl0s60x -ub`=);|YT1K]TfRu\$E7&`R7CPGH')g"/B+c)brN$S19lBO$slRo0k8S3,jJZ$C/{mLh;y`3?q<u^0W63?YDXMo4=Ks-46c:.\Vo;x>+*~i1RJBsAL7	Kr\K,YId|h(`v6&OV)'>(3re*w.M (c_.1O6J';cNiG?2~aC:7Hgi(t@ef!]f%a]KiD<c	*9hk>0I1o\aO j~/bqyWQcZU0[^R?_DX4?$nte{.	@ @Rp\J\}kXKPpwQV\.4cZW	OL0|s{1`*sZCntOs_`
fkhxSbNk8y'{t}KD9ll96F$2zA9HB)UtpGJ.TC+^	$$*g~a:c)YrLR}K!Fuo6E]XMv-s;f}t?f**x,APFW}xiameTTAj+1y&{A=Z,CYBkVa$'PSY#.nA-fOF=7y ~[,kuvP.8< XJKXG8qOeW(#KX"k<w2(g[WNvuK`=VtF3+>7Aty/b!)KSqV7;,P5|?GBJ;|i?r_f 9u.FY\<"tjZ6gI:`J"qjTY,O--75`>cy|;?y_V	P0K_dch!LWzmn++eKPhBQ1xEB~ ![{ V4PxEs{>z?f5Djy+9J2{wfam}HJ>{W+6FB8|HeEocGO+\rM`vHO&/kA)R<=e;/	esky*"FB1rR)up:@x&l8=+L+{NPSnI~UIgM%$m4'pRhM=UnBS:$0XA'	]=P\R0@{0o s-,\4
J>zI4Q~]fJzvLckoY1M(S7~cbdqE
U7
'D BtE?|u_WMg^\<|wck8$s@u:YA?!subo,*NED-0Q6H6~m(\]xreb?!nu_)Pu/xQ{T{a9-ms+m-X_L$m38AvHV|O*[("3@<`,;~5pOAw!h31QRi-.EGF~:W\Dm^$y@(>T! DP'0^]NtHvv+Eo&R4(VW1#b}]9nqf@JXT;Nnw2[5VsN
4*yv$__eQusyW 	Plk@/{0jCppfuv+_!as'oY;cHae:o?KKn*sB$+QCM['#QtiFLoa:G]Q{*0Iqv5vqo
E[_+19f]pz1wXT"[^dFj=,vgfz=db?fNSl;
}~A>A`i^N*@wVk}lq^)1Zez^zzg\dln9>-Wlc,]^3mig |hAdKh@DHMIl	P|/v+t~(7k?'GMw}m38i'";~A)k.)i K6m&k_E{#Ydt3LdIpWQan_`dv5sE8`e!O+T MbcO?Dw0Pb=:b%<Cl]uf]<zBtxf`:D++,Q\?^$zx^m(qkn&=7&IB})]|9@^cYt`Dp}M?P02s8PZ,F\Yc6>R>;cS"\kY+Sh:)-\8a"0(+Qi_i50p,\4T%~oy}-_HbH}a=y8TQ?5:7`	'B]QRmUy'%}xP_1yd$`iavp' P
y3s wjUd1\.]odf{$z%G+m2D'.Qy4em(A?T*`[U6rkGd'BqH~cO1{Yo8z8OOGC!x%|_!XkPq_.SJ:/ ]sd)Eq*x7GP:AZ,yRUE28'@`q|	:iOA1cD&6W>FI17YhN_"YRH>O?^@Fsx\y.l]5RQzAS>{':,h0T`,_+?T04w3-aX|rP=SmE:=7`(&J^iUh_mH)7<Jew3HPDxj@|=VT!dN./"(al:)JdPih.,B3)-:3G*U2'J
R~Y6=UEFB\[0qAjL^8qm<|w]x09mzgUzYcn)QarimTe|%QUX{{xI5[.Th0qJvEl+i:Va{GI{x'D^	<RshBm\bTV?dUxU'<hQf9!OAs,7jR4Z->%,A=)9A=$jF\9CPwB;_[XRyw9h:d.mzImaJ<\VT7^^ccJ+Go,P
YTi$+&-w,D(hm2!eDyK|O4"VlW5}=7U$mQjtfCGeN}&'*p|*OZ8>	rooLj/R'tJZ@?soYw;_oDeZrP]ntY?<GphkRb0L{a6oC.CnS,eE#q`%@?H=G@6b~~U!`?Vu@x}rp#^)w%kt;^@Bxw"(Imr'vWY9YG*.|c%(y7}e_<*9U.:@&8.2U5k(gqQj.8pHzFGt/]SVR,FhQSZ8{SF7y5z*69YR,c:{z]"~}TWERuLaW]@rOK~>7-%qA;h@-Q
gu#QWe|+Bn6BbPZv_a#dhb*^@LH0ST3e*GAnZ#jpWo3q$G,E8:m7M.9#o^:bEC{g_)?O;,,Ew:;XqTY{zZoKh<$.S2i_Jo
Cu!AW,('1L0F\B4@<5q	5[=g<:<l
#pT-!(B6ZEuJRY&2&=i<AA+#M;lDP![Z_~@	*C5Vmjs}gZTGi2m#p'b82,[ 
i(~8;4r4'8|S![{#;eX
&|d@)QL2r'9g@kO\P?$u#S	6M@|/3nf{]Y>e|'I	[n?dE9CPijGCC[2,4hZ]U(=1{nc3m\S[1`524*yED.e?j
*"0]|ihd=qW$uh+0L6jHIfnKX"&T2HU^\=mKE
S\X8]%6g~	?rNN0Cdk^w8.J
N
Xv?:6jvwq&
/&iqYLP</bhB'^by(PE]DQY-fnQid'A-20xE%c^Lu'LNsWdZ(96V:[r__Ur}bmh\wNRLTX.*4r	,,]QYCLa`3_7	aaZt^ii*Y;`~D4o/{_w Y,ZBF.gm%\z'aF:en{shAz,FvNoB8i~'Ll4zpy6F5i].4c{Mzg'7^9K`j>@%9N>e1}J{*G{xGB? !G@zbi-b>@z@85nd>((g%zwGxxbR672F=|#)\'g\4KTi-(2K_>6P
4hz$?aK6l$Y{zb|MeaV~luu9##.C#k$T_aA~eu*,tQavHy-wM9E!Bg'LyR9*%r
d2).{C\_}FFj$XrDUh>VZPnf/
C|j3/{6$tuc%Ct"4aVW9$<-NqdZa	JcDB;k<
jq1XDxP-	qRs;XY3."@@V3IP-=6k<T(y[3L4|JCADn
.a!E[lzmPPq.LxA|3;hW_/I0f5Gwccm+4=Zy}0fQhgV&.8+id_xi	
iCE5Iz!IChAv+=*wx,l.@.{h:	iFfQ.zmE(d6)l$U0$ofpk C[S6=i-kM%"mEE\&=e?'\/%9]20jA1mM')vWB~M?@Fu|^Izz5Nyl1Hl3k*wSx=\#$"ykRG!7RSLg[Y*dK^_H4}<?AC3x$$kBo- ]~lXlmocJ/0X47mS~Y7qE Gt/"j#?L	PK,v=+Jr5t*5#l</|%ASo*`80mDlyU,?Zk95r=.RM'=?U }ay;w="B9wR}.:}P/D8xV#ZQh)H5GxnDrrW4-;vghI$64"=dWdFb!2R1xbxNY3eg7m=@'NsX6	AwXH}I6'`3Q~iGKj<N
m3D0+^UWe\\k`i"J"1W<ZHum86o3xw)v';Jm>|:Fc-tl=81jmm%w}AL^)>GOsfRP5h>L)!|=exXz~iFb&cE+liSa/htH)N.tBNxU]'})\z3ORh
9>!WZ/PjIzA&Z;k	_xv@r7~A:,2X>GY'-m&"cb":y6S]Cx!-{*/Nk[tXt[=xELG*\U(\4M	y^DdAWbSvn()P;\(xnutDO>Gkq>gXo6$ 0ttItV+T0>vG{_P0t`=s}Da
4 +@m!^zDa\>,7A?Q`8VUTl/Sgvf9I{Hy
m?^)6c
Fmup|c >Y7ILG]mq^:>6hPp5	e@#^@|n0W-S-p@id5[<}\n.Hu][`=fM)}ZRZ\*d(44j6u
V`g''I-Ht~X(&8(}PJ!.vv\S /%.,whs)msYD'{yw\1<)jkpR*zB&795;6 ll>C)J3!LO_ipI"c/<O8=%M/GI9[ j(,dF!^+21Q4q?|&S;P?t )UPo^uPF{4ue-fu&s$<Bho!d'4LYN#E]"A;;!Fl:|a eAQHjpereU@oBVq:cYgN%PwAeV(Q,HyucZ+E#+"NK'SB&:gYN6	.W$1a@Nr<O/F#ZI,T3U>{,{E9ePqB\.YKf""U4NU&ZY0q=q0eI>Vl,J5}cT_)L`_
sc{'Jnvv:Su;gaB1kqp0.TAY|l{4j25]_s3py;)1?Dt'?fO,AN#i"Q{=>6L#},2A5'o/7=|jNGd#R\00mj 3yY3/[_h8[B:Q>6s_*B\EN4X 9]oAKw'Sd@!n.pu|q>OU[iR@]pwGB`:?1J8V,f)azWs`Rt"<y^+ *;BC9^{]&x%ke0ZKAuk+N28"iC
}9zj4J$o@ud7]I7tY'[ :wwaFsY197XvoR^En4)JT/*,	t3
R+^8+/z-9NiCw4VoWkBV5L o.$V`qz[Y(F*&`({m,D0~.P"d%BkOduEfqb&*g5`zA5C+F\4AU!gr(`>sfqB~sd0-=wclQ# `
Vy?8)A:>[.2,f__@Q
0&/LN4
8|.VV)"?mQ{y=7.fLR(5`Jk07PU'5MFPU=2&YC)r*ND~ca-9lCk!J*NRrV&-<o42cxUdN$_]EMit<Jz
*,SZfrN^FX#>X`>iSUQM:eTA+qyBH6)PIIvCMfjpSt>hBZS
"e_cZkG',,/Uk}
"*\1%nCp>D;_M3/HT'se4CJr5(FSZLIYi2p%R*\l`RQ|eUlp|!F$"XTCms;4Jp~\^5RzFJ.kmq/`,b6.a'7=EDy1~fB:3DP2"2L9X90icC]{<:,}`P]"enJdo*{p,F'pw$dSdZ]xQyn{f31!dH#nVjx3]s_?^ZcDpK~/
~!riSL`@lrUeGFo#8`auX&Xk|ZNl]Xa,2Dv>|4c\Vli0sW"|	g7|86XF=ED'&O]}XX7.M#*^$VAcUXgu|T8Px4{6x+hG8>K4%6Rt!]3m;Gz'Rc4+O,-yp"b=CY1xOE)rB>3nTl,jO,v\W*KybbA}##n1FhXpobc'5)F	J /1cD.a)=q18BI1|2gS>IqXp;S[{c_I",geQ''@:3-*3O583U@I!c33v]{,31y@"bpq>:PJi-aPkD^vY9YI!}h	7O0}u`N%7T5vVy/|v@&VQ3'n"Xz0_=>si*<|
rV 9=4q4]>\vqN"dZqN(Rsk,*MY9YUB2Mg~;9,jz8Q	9^x%<v-miFhc,XC='Kgkth-hp/XWZ\hyyAJgERWXZ_8$;ZJ"Gb( yi:i37()\twj-ka@D~pylECQs),0)ir=Ge o$SZ6^s4	zWoj;x[bH`Rc@
aVe!_EKGc4[?=}p4f[4Hq@eeG A4(^p/( 3rYf.>aMyGW:u2>e;}w@(\+
!6wpdln<%gh}dyRs^ 6"3Now9lv_}RdCb|_bWE(*#H@RTjWv^)66U$uVM \<8>fKwGY`c!G%(*7S7^:+NB9C[L(7JK,a~7lZ9ib'*96gsbvOGGT^--bml]cQ0IIS-?K.=akJ;rn?";g[X<wy
G>4`#CO6.aALK/@MYNeu(eOL(bg#KVPQXZtV!/,%_smo)83<{[<hbJU_>0XSX&Zm/&Q;%u-	y-abh~':sQ:0iA
3YJB,4d%N5\m e}%*s]{O}NRX`U:GxYA$wk~U};7tmH[p(+RT]nsr|k3G]+T\P61r,sg+BSg.bsVxw57.m8f!E)I{Eqjf}Ox+/F `+rKt4_[#LyM?RamBq4oeUA0/+mh]Bss+.q>ss0fARB7uQCz"O0o@KV
.N^wI,_5^|%0U:V8w*~q!?[	B.D">%KnK_ouTx	 fenFQ\.P|>_ia=RYj~r|'@=|@q*fq,MZ/DrAoRK1Yd+5'DhHOzn}NB" G NV#F]vHR6fENzE|}UctsoJVN==@p+BspMwWYy;Q>vVFcB'MmnQI#y8[7p3*vUW?.gF=h)Y};UA.?;1j:1F^
te&Tb9a-Zig!=rD	5M2TV5t/r~wK~nm^:9y*w#jjeTERdAjMhU!m$1Aw*fN#4B:k&1+F>`0}0&ewu*shyn_j{RGT.\NgOR9!e'WeOBtKRBihc~)4v,Cw_*PD6b&'WH.Vn=1
BbA&;**a9(dq4VN2@
._D04bh4l^K$	9%-n@&TcrD.\o0DkA/v0DrQj"mH=YLlbL9XwW\Zc0%Eq4qb69kiE*g?m/F{@>iUfv}g%pPo$"E+ka	I7<s_jdm'H^0Jmz_[8H\mY+OE:21&Us=!;&|j!WZ+zQOr9
Q9fg@+] bE)pR4&&hgd8&N	p8}}~$qyj_22(3XFmH
KugMdkAv3\y24/o><!l	t'[B]ZVN&$bx6C*xZcl"P.6zhO!h{55@fY#E:.#
4Aym!;8^	 wCmMs fD?lbz(eX0
wm(d62?
h@_Yf=@dvEx"MWWKhhm\<<HJ
RNMLxXyj!)SFK/Vt
1'dVuOj:DTiS>S%K^O\{j1v.X[.!H[W@:HAqol?|{PfSu6-Ii6-MkVZ/y)rIBml=Gv'vO~Q1y	o%H.0xOBD>1K6-Ha)v41g^7mb3dr#Jw=RMAbf:}`c\9!O$G\ID#
%+]>pu|#gFBbi\zkRX;ac!n)<\YV;Wd`h*PSoDcA>p2#bnU3BX2C`9KCD@B,W]XWG-d 5qtjg"5`?5
Li%%_r6D)YPF+qh(Y'zPWY8ScfcLFtFhARUIn69<1\d$wH4[;Q*@bfL8|WDr_$cvkq=z3JNek:=</)Ug-@no';/uKO'f4}SwxeJDO^$^_q`gWQv(VqYz7j<MFr	M6Ji4^NN](vo"$LnJO#K}\wO iw="x'Z }xg1yDK35~G8r6`4[`<?ki-5yvG^*UkmW[Q(Zc5:kZ&UV?>\Mv0V]6K$ifYMp=\+>VC>E0F;bF~|+C}%Y|8e\PiFE()~31-7}YuN1$Y{'0T=^ojrd)kTEU&b~~8%<PHR_(X[Bb-2oEPHp~lQ|i
@e4{FTPE1V'aT0^Lhc8}q+I:|F[hC	nV~.(AT*VOd$4t|.cZB<0|nN;n,+QmUwYYgbYCAW sI%+jawX_hAkWS'lIH03+(3^.-s
D\ao#Dt3#$9HF?7<@{wi,<V|PEJ0IH'Zq&56*){yT-W6t:^oN+[>!cwWWYC<9"u$/[rv,W 6qK/E0]0^FR5_G:>eKuWJi<Jv5faNCKQwb[?MH_-eoqo32-1a4j79vEA	]{Jqx6"WMSTo`'$TQbn4d^@Z&gEZtSIlM#@}57*-'a{HyLRP"3S16)gk[!4fs%0IT-$AiHRSMyj@)}_%_//ci@fF7~w`&?p4T4ZW.)#n\ag,!%iQNp7K=$9\w"RHb1}XFu{_Hn
J,|b_H%UoTr5Rr6Qtr	})M|n*kKkD`qd818DGa,8dqMlKnK13EjK{rqFRS	CM?*8(Ga
HN%9~XAVfxI!1QhqpMiq;K|VIGjN%P[A1wWu*VU&	;$/Xw?p0w}"Q`Ktc=W{JbqQe6J'sA";LqTC>ZQ(Uctkr^g=,G	f]ab6LQXqx2+}X]/>"yva.]E]#x#D<f>T3XUZ	io/B/%;4$y94WRn9Cl6.p?<b;vUCIe$*kLC.Cy;O'RkLbx{?SI
nOHt^vQg3v&wm!~"(>43sIIgR"@eg'+X=RG,`<?vQ)w)_5j[vcdjcy_/`v	foa,7
opX:v2XRUv\o2ao3X2)zg-UF'W'w=NG8z/jWJv7|4>9qs.+$)x+Jc%Ewj 7!P#V"x(S*
}tRMD1)0mdcuWVBSpQ6G@/Tj^Du#0*x#(`eD !d;z$Ixu>(1qEv[DO=d9n:w}
uw4nOST.mn2osOk-ws,z6RnKmGtOG#;>/w6gp&WS7i+| l;t?F*ht4~"#^rLVn?NGi_0{3DTO]*Of6G9.JnAy*0~T:9(l@`t9r%W=#0mk	U#.UD D=f|OgNI 2]^`ezX
=~6<
cs:15P(KH\Tc#C6JvoiCZ}X{7?	SJ
mNI(`NOG`RE3!Gc=v	%N,+)D%==4"h0=W}M|Wr@u/t@a(t3PSO*{
_>y{<VwxGVMX+>z5<~~S[c"vberIo&ns)Ti5^b+V;ccyIdOc6c h	qnFV!cs=Fv\1>w@+Ds3np5'#j"*n
ln/-GZ/%<u"#bXp.`2K(/.1V[+KJnM\|GhY<|&?Zy3@_['7a<%bobyo@ZZA{Ugqq&{]}e;qSp2|J&23:c5f|&gT71i-\itw?(/w4Q[muSGixt [M:0u-:O"3]rumpt3#)wJ=$DkdN!6KM#`![NWJq=	di12gz?+1,3&@pm-^4y&2
P`<N5Sd=Q 5eL5b@:Hq$@S([e6|lhvzqU`s)Vx4.-Tph"jeogFG/^3d'{ji2v2Cnw&x<x;.	$+ZX)[Z70,QJ2vC?9e7AHx:Z.sSq{J	_H[/[ufGArV&BB!l9D*6)g8NE]Ng9pt)05+8adze21saS/D$v{1q2xO0dlW,D.7H
@bY{5;V/]lnpl~lxtn*`>2ZOL5	)yH(O^l969FIsRlz?]b6PlZId#65zd#@FF%	I-ukM.pLSx(ktAh>a(4Jv\s`#[tjSKW@l{1+}p};A|@_t]^k
d~()$fz+@MHl=|E,MH[}I+"iZH%Z8#"?U36eXksa&cF1kfQl_Jtrv1~>G)r$$U{}{hpQS$6rM)foO,b@bI;V?@b'`o.=x%y|!kV(W51?BlUks,X(zZ8=oy)mRj_jRz7vm"RA|3@y[Z&f*r	/*r{>x?{e57d7hgI|.m)E`w!;q[p'5k8x1HU%r:~Sbq]#K:S8)bsa<6)')fmGe!OI/yLBmX	CD-'2LExw *@ie!0nKMW>~*f]!1NSKc"#`B6Dg;]4=ND?g!5ZE,_	| 4RDu&;O~Qy05]D=L' C)CkzpH>4kE0L	GysXFFTRCMa\|'Zv4P=SGl%'C~ioo6MTpV4T%==Ct(L/ 3![]7>EcR(	&Tya~<N^NhmN[~wR4UP{\Pouvpz5;c26mkH1\$:mmUnN0ed"TDft?~2tzS6\6\O	Sz?'LzE;J:[FRe"y3dh(G21i	D]V3#'nZ#TJcpRnJmD^MSPi2mW02`.%t.H@IRB=;=X!UurnRn7e|iJI<N(TnrD%8SI.8/9#kv/Q$<NYNKx;[dSOd@:+1)vBJV{\/7,T=Z/7>2J[NM*S5RLJV8#3T9Z6Zmt6HaKj#h]si
Lg%77@w%243f<r^^[dG(_&gJ_ozy,qsGLe}28f!&ntU:$_}v^u}g es-q>8!\Ue3|T\;ZbDUH4Y]JXpVa;<rAF0&kL\5D&}|k-.zjmM|8PPPD.i*bOr{E{fFTL.}f(RTDZod
@%LuO$a54M5?s,G_. Kzao5M"ajtH(#zzq^-j`Kuwkm"1mw?#3G!Ws"$h	-yo(z=ebRnBXx{NGM?QT#	V#8E\/U)V&l]#Wl<&$U1ZPb|2{5)^QvoE!eM[EFL^^N
xrs08RkG60qL-{${r<QO{sf~pra@pNK	vQ?1)Vblza}_ AV$;s
%#vMqCS~WOPt55=o74Uot8;kjh*a4B"MZ?s|	 je;II#9Rq0Tc5n{pQ"`3Y	HG^mqo]]Icn`1,#dhkcgr0V&(3NG%_D#68DM}~M#dw9Za
@~g^zw6=A`h&)5ufC?5u9c)w/R)P$-8ovTq5`hpb[	xqh;*g|j~H<q|.TDx|L0`Zo('k.zHWFy.*6C?OA4OD<i;JePmjt-3J]i_\~kmw<W.dQKq%jEx\P9gR14<>2iY7Vto!z#K	/BC.3}3:FbA<Wkiet~Jnh`Un|7$T)v}}7X$a5Iw5+aPi5q+6ZW!re/[x+'1*"{'WqWb
@``>9bcz6$Q!H# ]Rv0~+`@f4h[Ngz,T3K'M=_*Z+$J[yS:UO|*&9z2a^\-G#d@YS-fj`(r63|cbCs^1|	,00zI_(0i<fi8yfq'P:F.o0M
f'u3QK&R3<D~CD?-3V-\LGaATI5UbN#f];456g4|M2]mEx3\)8>9$aL	UXg9uqV68<^vLpWp3^J{RZC%>Ikud5GNGJS]a1E_4tgNDG@.(5Pbb$
tPh+OHI!]EG(Q6n4 Dl1=|M|!:HKn'tiSh(`*.v8n@FaJo.vS"hDTGB4`@7EY%[,w<>kBrpmn
'KDr]`fK.3[y82(|95dygcJ{# ,hV_z#odU-.k	S{+.k.KA[%h.z9xDlY~U27u63E|k;<!.A,(Igo}H">&?ug`m1'eOFhrV79/g#P"]uC>-2e[G|m_+pp7c	I.W[l;#i?O`p:im0<7YwXh5{d]EYE9d'Y#aje:Z/:x.a}lVR+_+*zwuBGmAX#>zL+&sNkCVa*ja1x,QUu@KnU0CJ7K7lRX$vq%9)fuK|<vJ3
"`my5sqC~1%g):4@h7vhZ7"!O[n0	0h_:$rHB?3Z<PQ8}=-m"TsfbWvVuKKrA,*+z:7`rpT'bjCE
 f5o}$gsunld5-?
J:-Phc"S/"~x7A#fO/'FNNB^m;]+'IP |eZ?1;)	
HZZ<8Ro\9
,*t;#5C09vL^@;RVkG6SNonY2th'}&:%42h@
|>6uuZ>5x/_XWN\N:Mql0i-y}%r8n#5urnN9lVt[YA06IAECb7
<D`^me<wc/1gx^,wHuPPfe;-y12d%6ga^-KB'&O@:tS\sHCddfVg?n"BQHl^XU(le$>MR9keEKmPe0,h!"y|u!(XqaXA56o}2.ovw~vCQXQrFkLFFtO<e]tL7uCf}br;b|j@{(M"=h>>R4Jmq	$~Iu.
f1d)nno#Ug|/#4GLK..3rP8~J\Rau!;	`<e4]\=`Q"=GZYmNh0 E14.=`V3I_qrklCGZ}Z	q\.GQU{1*/z({>mNJ1"=%tZr]6XY4xF!9fu8
N7ti3CKo7QiZ*',GcQM> RJAS
(YA!L_ "uf2aA*2%3f\yzOW^2r^-E3>*x-
?rHh1)>'9toJ'l5)^^@ES&"MLLzE)i2d2/n?z};zWGEs5![rAib|3yvcwDYn*?~f6\;;(mN)|vo*6KZ[_*~+2.8 o{ohzh_:+<| ULy;3#4''&@*p@WH X0
uN y;z4W.e\x^l$cRMaq,K9V5v]M3|Ovy-"UB'?z#]X%+LKuS09Zb4yI"zv }r`	)mzc)k=q	|%UE	g7$`XKQL-`U8dUm %z&m^#tb{_2~+W+X)a4TK<p"x?Ox5FohJ#mUsK0M-:Sqh|_Z/va#OSXK'm%{xT0VSD4vT]NmMM!jOHSkp_LO+
c|S0$HT!~a:l4)qC"]w/&pX.\iCL%m1PXE:-.seZhGfX)D$T+ay]w<~pcfTX$B-Y7wn	ZUdly/@`!& Xys|tA,+h.`/BcO#w;w!v'(~t3fV{++?Gv t+;P;1>5}/ `}I>[{Tr}eb4z(&p^nf7).xOHe0OGCw/@%u&?s]}uI)W\TYa9pM,U;C~DVz3hJrlr	>6W&%4H.jSSYYc9Ag#6OHZ+n8Pz%t+vY)!
,aW{1{3{SSSM]`V8dO-m)\WUTNq2\"9OB Eeml=_X{35$,.m}9'ex@#q{zEIIc|!{_Az0djsULEw\{`	2,dE\34, !ws~U#:aGYvFPDXuE#<B%0#]AtKhn)E;[m){	LBpN@k1`dj)&]k()}*HU#rsBuln[	6%X"dpb(GU.t\+q#_`NpmxBLE:wr33:DGCc~
L?|}b/(y>iYU
}.Pp2)b5&_q13lQG
B!v#=t [owzCUC"OH#S?YqAn=V6U_AyMjz^T`Jr`<:LRTA1F*(VR7/uFi:]F}1&N;ghSpc)*).3L5-@sNRnRQ,)R4#*tK_]_C0hL