 T)U+u6`jBk_q3/L=}lzeSvZ(	f8Qis?{]@	qi@9Y	+/@5)0XV{"[gtNSqTviF2ViST9HT(?R^E25K0~}9jy(x%e0 Gk&7
M3MD-'72{#(_|wfH1n#"cu(vrHp8/}'X\.'Biy?r@)mT!^S3AoqOfwro2RJvK}Ma28t t->2u}8P-]Wxg}S"},[*o@6Jk<V!5[A_1n)*sCnG\(&;NkPO8C#	|sWX^h3t'=4J1tH0m-9Z<.q$/s3W\NjU\y	+?'aTsL@-lYW[/gd0pA`JN#hXv7?-'o|S1K}Q]z%F=h[L|bPfHGcpT:zjV\w8kyY~G>_{x/$67t$,ngb}IB;OhK)!txBL'FsEw8 |g#y9T1:'++G0veyN&ChhNd<Tn:ay5nQ'bDQlyZ-o28jpIRr|DKXm%sl%UpG9=}S`z,}w$u]iEj8q~l#Bi8V8k0JS;B2:1nl &YCwH.w:1 R&\5)mZ^0V]1(\j']@`/dRG},Lx|JBO+c$GU*F]eYX`)C(x]8WN+LPSC1\;>*z0H.k2uV8J
Sv"/G O=@!Dp\$ ^foBB0rjr8_$"w`=%`d\;(.@}/\J<7NwFMseHbKx|.c1^8a RR#u<][t4Bi^.}lS/!8~LWrS-\/L)`{>G>A}G;-;fk%N$:%OUS|a}s9CL)%o.{6t	NJE}.2X<<mxQ4j=$*AP%H!\Zb
UyYu
DZT@n_nEQD/0ToU/]
?vAWvH5)>F0m&Bk"3.%/+?FC	5jW2(h@D`ap]i*O0TY7W;Fc\IJl?d$<2N0NM-tN[X;:5agA-{hSphZ<M%=>7|u"O>z$_v`5?x%Ct<1!X[Eq;)8/ RE-	dX .^o2@03>K)Qqi,O+gtF<;n*m)67g0<i/K=rkUb$<ynWbz1G4-]B1tUV'<WU>Jxc+SAb*|CA H]QL\^VU+rpP]Ai%ohvfX|\~q,gM~9os~z<\fa7}{y&2jY%Y}k SgU/'==%!&84mvst\ic\/HdA5Ft{nh`tBae;a=;k!HR)94u)k,W:<Xb3UT85IH|mBSSU;b95J\9;K}b&(8vPWb`_b>Aq87txfq1jkoc6kqyJov7z2KsDLe!x3jCY[{:gek\PmsCeBs0w#Pa1dV*>bP\v"CL_?	(%Wb0cD2IXAfS)`	V]5X59E{z2Rx+nDeizGU<aNa9M3N:`WxDc^9aQ[%,c=3}awBh?n f]9FR+>yU'O+1k'[WO~9]/2`?8n\=M0}QSAqCZpJ9d^BT])l7,U82A88xJ <\}u%#{Y<tWF2e[8H@fR{w0R(T.S7UHNo})p;<Ue3Zk$d!su10))_*.#{*T~)){+ea$${O[ YN+!c-<M=Dl(7'G.DF]MwZA&JA+Hn]im!;N-0u$}cYH4H.tJQ4}Rh!K$$S^U^?@!T@%kK/Q)|9&-|&y+oY3^4`V@U-c\]TJ,rXc-j5A0@!0k1"{q7vtbv87QfOhB\s$x*4S4B&]]+n
xj.0JC={X$mOtHh,MwCjHmD8uo?@RE1 )T[+gAM).tW=;ibz`!mWQd\s@:	WVTTi6v5bCW>%Y^7q2oeS(qt>2qLFA\7qk3i?Q=#y5QpK0P%eU@~i+E$@qc6p:_qds8Bl8kF@+cIZ+&rp!~UvM6[$F!'TaVb8Hg@N-($xOH,j'rBab{gi0@#4M;}{B|6v,S.'vvpf;*:jwovjwSji:@@NY!bu60c<bZYFVbH(.k
Dy6A7aMFh[VUE\eKbccbdz<T;!uFip]!$0$x11riI[vswK'`SfU=SPaIj9xf?9f#F~6B#!e-O*|-3R4=r@GWlQb"|u#z#t	)%E@\ZJ3+0`h>!vKrY6VGLo&w~'^X#J1Im]-Eiw1D/[c{6wwb<k#Vg4J'2?}:7";`Uxn!/]kP7qKL=)4246c2S!@yQ:z=xu|@(1BFV(&]Y3v.{NeAE2:)T,#4-sJMYhQIm YCh}K 1bTvd |a(j]sj$K3_-G:34nZ~fDp<d/Hr|qRylAm4~?G2@{&!T7Iq|sw1+HUv\vx7M5ae+K4,qec4rX7G!j=Ab;.)A`Qx#'j8M2XQ\]!+h[bZVv3i5#@j*\A>8M=%Z*V@PKj!d=4Yy!6S]v/vyfSh{caj~|:Fa3W+,8W{KZ<0V.?	F#?|Te<`I76JMV1!-o|$
%_7\
HvJtgDCr i&bxF1a-?;%{Gz|S@2S}J;_g?&woV3'n:)1$`]oY0bR|G[@tn('JZKe'^E?	n<?l7$+7oDYJdkC8$3c7"!|FI|Z""2)JyoH6Ijqt*fDG7`Yj3sbN3+DtE8cok gU}?;DndX9z^On875]"!/Ogbno-4S^Z^OQ#)^{w&ew@qTB27Ti[gzrgX(>Gnr3M.S9z?:l@k#]zZ*d~22[(aYZ<)R#<QKH`D/#6Z_;V-*db`QYCQDbTMaX.Uhk14|+$20rqTO@B/(k~bhkKGji."'J('#-3g+|@r5},1KZ2vC@}t!/M<=(X[xUArrS$a@.ZI1H'^y_3[^X#H3{yJn)}qa<0$V(,Xh%mv="yc+v*`F#Q)o27d~c`GPTAj7'KjA5.	<lCO`G<%oZHsUEmClr{:_tvD;r<$1]'Tes#-EiZ,)?\H[{L~DIvWd}ROK6#	"5YH?_H>[j")S$
~lnTrx56
^W)^
mdt_ZT
@P~UK%D/d1D:?w~(G*NhD+CF:H0.fRpw";YP$'a	{X.],EVnbD;/S!/;u_89k) `%R?/h>>,>393	]ti`G SIZ)=#NXhpCdk;l31!OntTK;`/_Iav#zlq*=FU%g"]kAx#TV88lbB"v|foA=K=C.3< y	+o(e-'~	zVq;'r;t_/t3r_~$UkKEY	&B"SuV~w?|::j@hQO3W_(K## h*+"]&sQPPqEu*:dP#N
3Y:M59Y#naULe^aFYwgpD{+,6\E\P2+C|NcT/S+fCFOn=n%@VD8J>3.~M)L'}qK~b:~Lw}N\sH*3na3DAr|=6I{j_r+>:vTt{Rl1IkIF`EOL~i6{.u%C|WuC@fO0	+2QOuYAQfHj
O?\;;Y&?E-B&3c8"l&`	?srj	X_JZ}exH?g6<2h8@@vVg6_FE1Q^2oR#ElJq.]UzvJ0<_=F.z_"~dVtQyz[*vp`a">&
*9Q{0Ks3<eL-+#IbeZX5N}2d_AA!"\T	V,^F 3N=$YBSCZwVyNs*<>ttD<>["3WeaZQ5tDZ+v^:,W55Dz{d 0}`(Rx&XL_3EM}pY^SU9d'~V>A\@rG7{aOdN~!|)Q6+^=w~&P4u/{stRj3#~P^6v#Yh'<00OgTa@2jq"^aC]2V]>3):dsO%<\_s-x/q)/rVY="ViA?(?..3m>D)7^	naJ;mW)[f]h=~Ao:_0w]k:9NUF~{;]$:;KRUr`Yx9qK(uwwBqeZkl30 k'aAG-f9j`h3J0V>1M_S;45%w\>RMR][70gU+-HMn(CmY(rcJ)_S#0 J{_a*'-#6ue"&4+PO<eE5%qkl;GmQAo4.,Px`rb*\HTS%0HXYvDJ~f2JPy<h.(S.9p7:Y7S^@k<P3*5d!R/_q (;19q;]!yN1q>*|1Ttq~3>&x&X#SmQo~;NKu/_uH-xelxVo*:>Ro^G-b/YPGxNX*>'UjE`Z%"fh!+9eodN$(g5E):X&Z!(a;U(KF,S;}gVv9/KD9s7O;)|om"@xQInir@n3 ?`;qwzKZJN)==MoV	kdq,BO}KM~Jok
gGNA?M#wV^.pw&}xEx.C8S4=C7XO{jA:5UX[(/l_7xA[d}fWYeoBk,T|$6f!Bd%&ar?U,d3F]f<t.L9()i'`uX/n}S\5S84Cir'+,<;z/iA&hbaDi{S4u-kcM|cfP?E&p@g-
9FK$.BVf#AjL<TTu&=S}ZBcd@>k^	6?vD;UW;g]&5Z01J.REmM',{
oW5J0%t	F 
;:q}pOKSX6EoS7	7[`+p`8U;DWc;Xr4Zu>]\>6STNzk^]a%=W&Smtchrr\Wb`68	r8oV>!TEa~]fQ{Ru%e40O
Z%yi$%iFqTZBtiR=` }AGiPjft
xd2cf.9-C];F2Xd3,z@J4WQ\X<a@*MvQ;\P~<L,OZ'^e+ee0yri%Z8egBp1mu!2c^%:mWd9(!p7Ii{inXlDzn\_/%xOT2Q9|g~Jw8g'ujzG=IU8"qc()Rz8jBkjD BA^IO]xqpik+Y+&`vBpoN{FSMzbtRh6b)js<5e*z1JcM\XnaS$&OZx:s	!c*4rtiz*MM
Ot|$0aF
.'@LfFy5=$+6E1U6 pRg,-<^7N(YIomWaxK`#^B18 {fA6)jU%
$v1PiL*T0|B*be'W!rvWt>J_}<=a!h{LL^F	u2_P&mF,N6H|Q16~	O~jG{}'dd4SB{UGdLBo)Ipg/hv9Bur}		6j@!^87Jt2kZIkCU*yyXF8z	8>P;ar'r6YwtQMZYbdy8wg)"7z?>=<*zx#0iKI v>!RWY<1}1:xmDo&H{`d6j^x+i1!KNJSgr8n1Wce:A(}<h?}0
nM2(CZSnvN;MVO/YJ&WK-9Wi8~d{!4waI;;@\/zvHt,ZBoEvS0IR/+=N-J#t<w$jLuP*$2wLg(uK~=qHB!!R
w~`na7FIEX=*+!BcCDS+KExOGEJ\Pg7.x~n?j'* >o_Zd;>^zL71K;"{e'G\xg6;Cn7="M'qQ`OU>tR/)+><l-
*x_f(nP1XHSa4!
n3{";3@3b R!')kC*E)|iaG|m_vC41*Awp1KHf gp~]%{@}x&psdTwn#nj`^&@8^hbn|82-}'7Bl]b	KmKq&.Y+y!)"	zlooVe y%0Z>gv g$5'.Yd^'j}gmYY,|lKd1-p\egec)z^y=!b}hi_v6d;Og<jLb)3(iJc$J,a`5TbJ(&BjmjMONRJVnab<*|xz!}[N,95.?Z8PxK.G =oD!9R/qC\x6g[==};/Z\'&eVKLQa.0Ht`)3
_f1@M^f6^u[,5Lhj*Aa Wh_=;;oWOgz>a)N>=Trh@O@98Ne.m^vWMcMcG6mkwlE'2&k1y!$QOv7j>D3mOvc*nI$9K}=K%2QElm"2/,S4*%fxbcD':udAFn4Tz85_VH^Flp,8ih[umY^%~lk_8@o#vA13E/`5m,1o0}uVLF&3uqc6\4$
Jfo}1JZ8!I#I=y0A5-[H67	4E<h|1hr3Z6hpqbD#AqQG,-b&iIP*	%-yEy-4l`FD4zEm3<?d/QAL{lrqjYH+\^!HOBX[	]'3<mTulWQU`xdYDBSthF
b1vfOM[5%Z9_sB_! (VU24uyDN4J(3<:`^XtBR+c}qQ/y}s-KA?3TQj/m#u(!`rEOBV(~!%_E3.f7mGNDY]G> IR;:x??[L$IC&Eyb-"`zsyr[^7^7Jk$7_9kP&m=kb
)A/t.@Nd_RQRz]bzZP.2S0mB?{Q3_~G7gR>MD%!p@!N>9,2@T:xkGBuHc'd;Usr}\dsN'k-aES+wWml\5p#?'[ctBl~pKH}f{50n^]
tl\5>gf8e3,q`YK_P1Y	=%Zt{/
..z~?1n9&{nh,D_"IUj1@G1:	N:7*zm?!]7"/:B==5nl) BAQ*jhV=HXo'EtZ2>F#pH$Sj2V~nj"K9sMeiC8YZ'ic<xv(kW(t$~7u1@[/j?5xw}BMlWxXh)Bd=D2U+Jm	GVnc	:O=3%zJoq3h\gY,Xe \
<eESk{}%+c78rF 3nXc[6S`GoUf*vU^a9:YK7k4bB(Q32?me#PtY*8]AE:"HK}ZM*<V5)	]?iWiUQjh'R]8]c?gMi	?
P!#Xupqr6{%uy-dhz"0P*;K0lZzNZX,A\'o8b?!JSPs9x*"Zt2	7B');Cwei^-ZMMXg@#M,H9gL'Qrte1Bp\rkCN4j}"wQ>XzAg$Q,wu~c*|,6BHb:nik1[Mqy~zRrf^HN7-}EF[;W:Dz3R\ay#ffd"0g8fayqV=FufesTeO6	fkdw7	I}2wFRnWJ+=vl^8ba)?		p_(r%sh?PKwXDf@M{TfQy0[}HL]AW'
{;Y0ubc=.7*L[yXctL:_E/PC\jY>``[t@rMsOjV-c/i;YGCeUf?O!^K^M9+C{Rt31{Lzz<{zoh68i0.db_D}L{T@.mBmWe[QcZ{#*Ipawky
B^]P>	NB&ia'*08`TYF^^SO?}Qw`F|:
X<y~<-mYqkXPCf5&jg3Osu((#!+g]u<EV)>rd4V+#+B*wzb[`*ml>_F;m2`PQM0]nCP=R!F=&:Gd^[S0WF*8L=vH,ZF+(7`@8. [
hUXZj_Bn2l("<7"P7I8t4qWqh_Yw>^!40_#[^#rh{nE!;>8^=NU0c#/hstwE{H,)fx*H+OAOVC:
 8PlIRnHu8!gRB|vvpU+E}UY)cEv1GoNS[s;;9,f>HigAkWLAl3Z&a{-{nk!4y'(RWvDB^ARx;H7t7&T@!+s1;W*ol*ZP6oRhd eOC}wUAJv+}oJ({MAAVc[2>_DczjIW{bDktnuB.clPL6nS
-U	|,$v"MfT|Fa$SQ?^Y~$i$p/;,pS=B`r9*2Fcq<W\{'q`4eE}H')NMuE2<'abH]f0LU*IuQ!"8r	Yg/ReT1]in<T%'5b"odl57?l[o(4th(7'
z;eN~l;2zgsuu^~E4.LHT9U(DU0B.3.xqLppEWA$w&J~#]wt0c-p	q$3E|!<<>+KPYA
>'H_Swc?A"/CEF0	~g\nt;Ii%AkG!&_V6osBO=o)'+2E~\Km
A7ut3d,1+3[P[NTIl%%'3EOYkXoORLgkM.5bZEV8sZI*cmyoIWYq'E]tp;L9%Gl+XVF33^cQxH7j=lZfu},kDv[nM2'%w1.7rDv9nK)rZ.YYLiAub1r.&(@vya&$:zj,0JDQBqi=7tpRbwkz?D{Tq] z@UnFwq15HKk8jR&Ah=;+G=+f}z;8vAb@;5636]][%K-NVB@/c#8,MZ
.eC?)k 2.%UCVb?	s,fl2Dm[`fPG#jl.CbR5*l]CLRG7iZN-yxLC>cbGh'!r5,#!Y$FsrN]lAj'Tk
Mw8mo7	tVF'gOzRT4:gE7(V1XaJot\J97J?9(8J^MF$e/<u#:RrN*1pl_pYbK]:;phF4 !8+Tg1D_M_B2!{ZP&Q:%^?PgQFp>FZ]x6ja.7y[faQF:f9w47u`LSK1ELig()?P0x&6o-UYeF=eD'wg#b/QKWmfd[FXkqk6aLhAN3.&E-.uw/(azLXINn%Fyk[7=4^<l='LDp [
0.& ^2Ot}dcEfX$N_})aI6:_"=NxlmrBxysrl*6=~YL~0Ff(lc'~dU6i:K.'wB&UC"F_570EyJgi!Ju":buMW/[($JatrC*d+S&!k(XcT0*G<G"`}LH">
*ir5>z_$(Nl'U1B^yd}I}3L*+FD
t|=Blo0!& l[G(k*8?p%7Jhydsp9b4*TzK?TZD(V{dXi+\D	+ylwXqB{Ol_D.I2CcN`i/<!KX,XW YNO70eU+MN&Gi=,m0T=V/o.+_Yll))mg0UASHpPb<!0WZeURt;I<n];z_wJCfR^h\Ka{b"CAN}P"aVMXz"Jd6RR=D>r59<?&QyH"N,LG^H!mO\5r%!J$rL{-vIz(Aut,gC(0"ZHheW8bPDKL%(z]epC"aUbixW]V.!x0
s]EQs*v
REdM`F[PpDYeO$1R#istj?<va
bK|pztfB</h_|r	Nn\^po1|Pc7C8lX@ZzjST"Rt#%"kfn72Y
v't;'spK{X
q\DJPX^1Pbo:?Egso_TB{+$_j#" t
b(i,_%}"n*\Q/Ud4tL]ipId[MtyY0Rvb`JbMKx\,07	6Q[3ze~>g)\;=X_	a%gi'L%ewNLF`P {p5C=]^cK%S}"-Ikdm	CDSb9$vG	|@$_f"[u!gh/	,||3!j`ra7>lCVqgIvFIn3:/i},am9iXG	YSY/fgWU"&RQX("5'6?l;Qo|;Qd.AZ6&	sJ>F;0z)!Jd8Ch!}##)q;
5S()h!IZa(-kZ8u7]ibn."F)1Wl=JG=p(}J`5_*xSdS5/
Bbp&p.".@%
:NiC_|Pvcs{BF|it71;|6t:rvN*WG1HDxLx~QUk9jx{p8nA6AvDSJKY(lVA]YKz)!KDi5D2ny@pkC!dQBCVS}#fmJ$3DdmXf[}	=ki+)lN1{,TsWU^A6B|-G#HvWfK_h}TZsa"afPWZj>>V@rLg%0
q,o05D=h
zlMXme`Ny]x1a-aP04Hv_XQN%yxL~q$eA=&5\lV&,^:qwlD;w["@-7HO:AX{u;d]gx6eX5_4DevU#2+;q82-Cu@"PKs</mpq;7oUZ|GSrtMf0jf2zuN}evJ\!L'js({6+p.LGo)`.LYA1'9)s&GP?xxuh?vHXE	YZ2Zds*\ZSlUwQJ6fr|hOZlf*:zcrsY>M5:s='!V'5o-=bzAmcW$soB\Py6a<<Z47q.++0-9x%x_!wB	51DEigyqOW_\v"#BF&jFnXr"l`1/Jd~H4\j |0b5FD39n^	!qGcGIHW0;3M7#,4r#gP&uMb)imQY4 jMIh;Kqk"8bTQ6_e}51t:!dzp6O&NB%9/%n)|+Wm0V3B/>j_`*HZ06Tp&:qrDAnjI'Y!6TXiLa^OpN:D>}7VE~"d;Ho}fX9r/p1)9.SJieWV	,#>jv2Qf{C7L`~ci<uwHyL-VD"5#\>a84PS3\EPmxEgB{b5)_zjJNr]O=e KV{$V1B*\7Xe&Nxfn>:^aV/2
pT@ j?E(tl&G^/W|q7yau@5IgJKP	=H6\<*^1BW=*Ioz"nXO8g2S(E"zKwmo>v={~[:ZMMs~o]e@="o"7#.qh,3z0ukBatbJuP55.1;
VN*X:>RW 5"Ac {^%6ol*zjkI2uEuyWm[?`{aIAIht"%m`CV )8&it$@xaL8W|{%=RPdi*98jt
@VYR?ux(LIm.<zHP{|@kCLJ,%ae!7x6&w:NK@^Mh8PLq=<_81-P*vi$4}
kFm~Ba%rT\.Zdw~;2 42q)_(z|#oy.J!UK
:lU|2Y\W}sdD!){R$~\lgnk+Lx(:Ph v,!zj0%Y]7"MEF\&D"5.rRGt=BC~tloInTR-N)W;`m|	,*-i\	gd2V}<.V6|CU)<]G!LpOi5n;:i|0hW8O'=$trs)!f'	,{uv:'+3T?9:+`[&n6/@f.TA>1er&K9)SEHC6{f@We>/e
;k=<=p90JLTO&>0#by5YMM*2;xG D%-(@L5[m\_4Q9@ e(n-0V?.w0aicW)kH}VuPK>e7<i0Tc`m@?
s%_[2x]+&"r4QgFUmfK5;K0@${K-WfPR>l/MsFG_q	#*Qcob	ML7t~_Jm%f3dT{Y&<R=q"d^*Xy,*0TCb~o3}|j	9Mk5sAj
s.\$0-H-+WkM:V	<lr$Oj-]y=Z5^Za))V"XD/	\1uP9g@XV	;-5
uU=
z.`s05	t&4+,*%Z\susIb*)~F.^kqe(],&'gqDaZCHWXV-_c5#w*BDbVw=xD./fU'K`za#pl(:"%%"u9w%`	Tk-@Tn,4w10~a)/`^WU/~l<}MZodQ{m{TE2'DN(8E'pe(l3snn)C<<L+73Pp q?4 ux:3#a@!7x']oP_-a(o"9E'\;TSE85^SNtv07f{ g=Z$oZI;7LwJka:SHQ7<5I4rL/jXNg9Mv\YmwF1<h\9\`[VB	C3;gbhnkvu:*5zOB%HNfq-d_EOF%,|p/"XgXb2&Bn6jI\;xI_,dJsk)[2(^aM*/!{(e"M^]@G"h}0a\f=[9~
|=|CpLQMU. ,-9ixC1]@oB?nW^S>onG0Y2@:[g[@\f	Krv?{?AIrY^UJ~,GJc!]KW"f
$@^xm<1|	5C_dm?&o#-hgB;4J.$%T+l?Z${7.~8?!.4.dC(`:u*~.y:$yT
CYnMn4QU%`Gs8Hxtrs\Iq+Q(;Jz%DQtJMSt6f_q;PW=w}#E6[yc$$%j,@mk(XM7zZiSp=56*lC_bMKq#*O2U#tA~K]TS|A`xlrr3ML">bAcxFAG,lAp4}]{VV}kGl}Xf<RY6CRQ*D_ uKduH~A$/h7T	DQBBZ t
7Dh%)mIEBI2%J:{^"hPxdAZE8kOevW(NX}:qSWRzSle-a=hT22$'4i[13?at{1$S*+c)	'VBdr{w"d0GZaGf%[~H#g4^X.+mAwjX|j0B]c.nGf,u=S
,M8kTzO@;<D[
Va7j;g2g"?=jZ
/P=KQLpmA5v_U,'}{fdZ'gA_T`]?s9+KxSA!;?0<3NO1A8w5^"IW?;PD6(P9H;#)16v-*\\3t1UmN:	kkOE;)@89
|0z]S]sU;FXK%fP*F$39.<xqv`UjD@`]}LF<:ay=B1&w<quhcA7y4k~"C2;s~^fS@Gg>MPh(uBT%y'!8X82(2sC24i64H/|W`^>`;?ZVRnVNo$mkS=1zsk"uWsGH<_l)x3]SBC`1k\.s5t31J/@3a;'zRIZlo5W+bjL(2'nMtg-[z`mV:UB@NC]Scr+E9|EEK`tQMb-1o%@t-i7 xbD;1$1	1~<"+*vB.C07PuWeis6Fz!~#aw26EN"CRt._k]v|(H+2c){G,Vhs
9+^Pw^Mg!-ac% zU<R)X@|yoA'F2J(~_os<P7NTt|G	W|^ty]t@Es;!d`WCRE>0rPD$J2dvY+aUvK#WNGcf{A?2Mf`*P+$PF'Y|POJ/ba-qupbAToAAJKR+JjcSiJL[+.|Ws[xv{j.fX5"k5l1}&.tU	o`ShL-#VU2ba':&plKNl7DO1gNsRD>{G`|s&B_|$#R)y3
~2m!~3* v>\W,)M$/uN9d<h9RFPlM_45G)W"qTAg2]B%PvL.+= E3~dRp2qK&^G=Quh&5JQ=4?R)2|:V;yGaJ0<sc=l [$1j[WUq%;hhA_P-f${-a9'"I7juO2eB=K>]0!A|rZ0NJvFK'}Wh<8q+@LF..^S#pNLO*c@$JP!tPO4#|9'8W{X@x|+>2h5NL1Jt|.<.1`W	`nfD=l7\L4m'^g@+&BGI|O8Kwe(8S{$
/=4  Ggr~RDoP&(;bn	xbp7,	e+O4S6x6qh{|P%iz}}?BM%--3TW!SjjwHX. 6j;W%>cZB,]K
	$VOQ(`g:!?Fh	&W[kE+90F;8La_e;Si;EmZj&#u~BaofEpk3gV9o!!YQOy#PDWtKx@wQSXeuAx"06$_#>|0M@'uB~qTg6'?zV-jqr5F&*aYmZ8Px#Euk\R5K+x]y
{KWg"4g|\fxk>(OOv1{%!<)^f$P"h' <* @`#zI%8>!z(~2S}2wI5F-hg?Txx@rbFj5_k*tZuWOd"~%s9t?dhh)
Bu1B2?LJ]y;o#mb>G^=3*qA{nfjJ.;PR\desj1gF$34-(/G-1lm"P{~OP:d;pU#1(7k/L^fg$%wAR2~Jt:N8B]Y$m>~Tm,|>TD$_?i"lH&jkr'CMr%J)aQMA5JPhn(/.k_9\Mi0X[:E=T$J0A\ d~Y%ykPO[hkiG:E6vV
N#vu`BuiC
uV>RXG#2/| <^-ENQiYUiYQwB=7oL~[Oj;fJ9x\3q9`"uab8o`{,Q]#qDw5d.!VO_ScHt\t'A9r"@v!Urf}@j4,C*b/)x31\PU.v-nS(ZCh;=^]8-d]`H(Xs<|;l#zj6muY[_#G(eX2f"T&F.W`.61	w<cBQ	`cNpiMie~(I>Ng&5+)!{e1ni/W
t4d`4Vc>&*Ghb#&A>aXb:02l7FFSN+:6sbHxYsb:.Y7ywxDt}5jgmf-up+EF]A
k8r>KmsHGGeJ,Y4G9,ECd)RbeUb`xoi*T-a-0Vcou!@9`/h=*M-bZ,.$=w{"C|#hWqwvJIAXc%@o3J5&PCG!nA40!'Gpw'^
B,TQPpjl+iCr,`22OJ;1:D	B&`5"o/dU.{,s_}Pwv796Q76
U$:_#mPwI3YwzLke ZIR)otadVe(,"(3P``60XjLL-cGzAh'nP:PRh6c}^1Q	C+7tYYM2Yruv
_{a@{'F_O^;t,raM=Y9jfY)J)X`F29NQY@Y:?% Cd:@HO	~i0ZPW;Xq(oo{
yTu	,M ^if\>gAeeUsd	iOuG4Ckfzz<KG'5ao'T	rJ)27" r.
+B?!KEa44B0x.`e5CQ3"sBIpOH%ta=qwhH
,gACCf0Uc#adSpok8)tz&!;Ge|A}/5JZ:hK\Z:ztdU={{>(b<Th|??![C38Cee\]v.F-_sZKcML'xFFL4z/o8SoOre	-Rn[&gg `e"E.21H+"7+; hZ{nbk}$z\1fynD(-,k-CpTwzU*8Ye7B^^i*x2r	>pT)mwhvl`_T/$hnYA*v;roOHTk79"\ySG2[wv@n*3AF%fVCg~	'OP]Yz&a_*":Hnox{`+aU<C:O	@4[9\)_S5Q6DW1rt+q
g%PUGp_?E&>/f!Xci |WI?.\:5*^y;\?CL&$*Zco1:3#[2\F<Yxz&8W#YvSIXqg{t1=>1PBApV9%8?W{uxZd:?gWHLf
ZX( g<ZwP1{G-,vMM#=]<U|0nYlc.aYty^0p>E?W}}plr\q(QBb$]JRh$@\Wg{cwbs?NZ~z^#w`pNF7_VQc'GN"X.Ww{'	~Sj/ab-}<JJxju!?^Mw!v	}Irb:wX]^+A;]:*we[V}^ZMZ@rt`V3*SWCAjs #OU~})zkmVf'%=OFyF3rG/nEVADE	<oGo	aN0#)Hf'$gm`9!2*E<BN|sP><S ZhVd+Kw~q@NBI{qn\ IoIYW<U0>\lma#ZZ+JN+:[mk
{FbMhP]'v>vc/[h(md1MetLG7by xJ~;S,=nO_ON%(#G4Jf/\40|hF/AT_E~P-Uf^xyKLa[Kb~~TULJ;U F,%Z0[EU#! SMs1/aWi\&Wcu*-i*3i,kg(Jg7l>L:@>7~vLWX	kp"Cj|)Y&-D&p,>2
zz~&jY8,T"4. $6gLh^rt,	KB"J0'w0Lw%vSk;2+GyyXH>PMX,5k(*jt66- yV$l2dY_Xr;gbL/!"NyCaVqu+4<r+*S&D-$H+nz]@r>=pUOLzX4'IY[lT)-'X,
W,xnHP<CNxWuw'NkP 7$;$'D{'C,h]TS,$`BCYszE^<w.r$i<VO$8?w5 C1FX|yr	h`b)0TunXnUQbeB\Z)&.q
<~p1vU
_jw7:@u<)}Mje"lHo@dM#K*v1\|hKbk;a gS=NgX$Z~NeD~M12*tb\lx@EYIV8=U7|8Xx63'}?+h&*[qGf=Fq7B'H/OOLb0N+N;34zS"JEi%3u3T
w6\o57z5#PiKgjVt?Dy?ov^%S3S04C)(Qv'ui{U1ZFe^NWj{whkR;Tw[$].Ef"fX@7&+j$4{xw:Ep;NElH:aVsq8FV%\sOlF2Y(3U7XD](&XnOSO!*Rn9UdSNhe!AYh<>E3j7lZ1{qFhU}x|l^^LsTO2z>2b{cJWHjZGf%b6y+wV5;GXlg\7(henDj?mce=u.}H0[9*v8REHa<^TlH8a$9&x?#k<{(D8clUJn|JWl^|Smu3+})UT*rmiZBZ@
!'nGA3-nWIr|=xunp9S{	=!tV~*qeV0 BF"	q*6\X%nE0<,17#s]6%LHr`x2<!#\]#W1Xo-zlFmGi%]\GyXAi#.\T#cvNmZ&tUZ=/zLQQo_|)7	yOb1ps{G
/fCY:a~Y2UeAPSPQ"([D3XwK~7YO/J{MX/_1>
WoDEW?0;WL	6b"DpSr<>-D}a~j6O(vfSlMSJ9eF[oY"\}$fW<U`rTnK:f+XYjD'`So<9ev8}f"o'}Pj_@TN}~:obbSssO}[
A1BJ-,EY(
;3d ?-0EF|N7^%?dSPo~MutdxTSNcXlwX1|"bf<w(qtF@?{|{*_n=	fg6g] B*;*,P1l] 8Bj>"P-~h[V\1wNM[T,jN<6-Pf,.(IpO\vE4Q{3up%P"'MM,H%9:)Yh
S?_!B@2ok{M2mq
N?O:/IJ0ntNhQ=kPq+2b6	;8H7-Vd{k8/iH3mz	e>+ig%O>&	0P qin\msqJ|,St(2RO;|4a-uujd3Wm2s]6 by_zJVn!R>:."QAdvJkTCc/c2!;O5
E(u\8r:^2*3>,Xb$yZx"cg4Qy`&O4I8bhR/AR<mw_*W=fKAvIx5qtYzR4d!d3A^<,liI1K@6{A;GSRz7H<&g9{b8%&2gX%~s>79N\Qzy1 !~NQx5\pw
[1d{
%_w'sy01H
ogS<@,`IAVk=+6$n=#@/}woN4jp[D)r(s{{)VZ_,qPn<6V@Wh*a Ee{gWmC/9Z%V5/P;f.TkB.xy"us9xbR6Uz4;7d)%hKGP_h2`4/&+@oF5?Vh)>0@~&}'5)deWL qcCWb^FBmRz.-Io(ca)7'o#.Jmh
G-0-?F
hTws)2[iLr}7'te=M6 F^(xd"%_
Djp4"ibXYtt,JWDslq9O5kt?1+)K=^&H5,	C(`AX]U\7ke'a>A-""=A-6U%W?rI7i4O@Y.0gM68	Ja(xl>}^,Z;NMl3p,!b J['.W27~sHvJrYdaZ6}')@KN=,=.\HS-w@hMe=)D@08+,L1Z*G}saK_'2yIEdWQA)w2I|b 4qDWs1d)^t>	K`iu&f-{n}J>W<R"J/>_kxuK\Sept3a~g{)mAFO27+gpr\cbstW4nH?L;WKOING)+xN%%Iv	zIUbBULM
J1CR x0QiN9EZi=mK/v<&9jeMp#'
D_:h{F+2-&T!bsO>#	]qt=j%fwBK%K1<Cs~_Bzwhm|8u!)r tca)=@j-TFp7Ru4xYsTvg eD<IL!mVx)xe5%EH5@!|hvH$387Tg4\_[c#In+JW[|t9id7A|%0xGb7O,7Lg\m|8N'D.[T9MB1FmSJkDr7&?B;AST2dyD(0Amt%
7`)yl zI3z'mD}7kiX%g/IbPZ86;TYWi*WtoJ*}Ya">I`i1\-V|zl\Ao&^l[sjSe}jqfP[5%	3Ia}|J8P8?M@hD|Q{'Y7W=khaVAl9%+GLH)T;`oo})&e0{v8w8W +~<F!L)P;Lu51O>qGekGj(mvgn@D~D(CBVSU~
Jzi\'
t)|]nCjfBdklA6EbFrQ^D":YsyGyKw!jUN05R4uVMw\P r(hB^nYU5%ggpuaSgjT6;
,l:K%.Cv(bXNM:i;g?5#+;PO{.pBY4QZ	|1r__q	JYU|p<+ G[SXo%,{&V%[$;QA2!Fo@]2V
VEz5u-yA!l7|DN*:x%y}EGzZ-M~?K+FJp1Dbj4XG-`]'BvQP`J&ut0]ou>C&;$c[wsu6%"fI&"Z;-	H#"C1`Q_[K?zI^k$v!OnYeEb@R*$rpPK$s#'lr,T?yq|GGMNO` ?iOh.Jj)J$ucK.~vw}	N5w;N%l@vt#Ey.Quj'o7R55U}sR1e"	fp7@<>}N<-jdjH;~J(}L*QxgNG#I,g0ry*E3D==-Y3XoswS!2(s(	"b|Nl/w~+OoCB"$WJxN)$,cpqsu/"?M>[XirNxp5.OdYY(_]p'm-Q@/})"z6@M8FBjt|6\N'HyyZw|r&WV-NmMY&7I}}O;9Cx7m
Q|@UT"
j,f*:_c{y|!k]d1UcM_Kp+Nmmm'>qV@5[71
jUMp.*%}c_/jWZc%9ab>DjL`8b!Q=h5b`DpJ32?c_F2r.Dl,iw(mK[lit&g:XhiNtF}"'YI>14"W6vU
{'CW.Y8dqDxDJv`SP(ZF[K3lHG$q+*DK1%ju}FX7zBGJH!ke0`x{n;UaabXwnqAF]bD|OVua]IP1H\h-g
Y U
`9v/f{l_h47OCh7$eBi%g-L\Q@2*gUOA}r71A
uwjnTPR3
yAY@I"R/,CPCd{a+]%@4pCf(\R,RQGn"`%fij7+f|t^.AEu>%PxUEo9a?`Q\Xw`&h:xYyA*)$[SfeMh0qx'P3mp'C{_5;-1TEJ9xx%\v7&KfJx?eu>Q$s 	0Cu/\,22gN-$?NJ"		Q)*4gN98FLE70\&P6h."+e@Mg9dBtY,g&$]^ @J'Wq;].zONN^1%{L{2fo:.'D\d "7;>UvPj/~U9oXa~kS]iG%)"IHkb~|F&Mq.wWkZbY7Jc;b-21l5s{/2a[s$gvhn6V[ORS,UjV[es;\Pe;%3l1QU-h_'Al$z|Ff|=?Yx0R|]knX?#FGTb1V+Eh(b>L~D[M<BfXE7OuALgh^K+Uk8V{pS]rxdv
DxJ+7$]nK_9SEs5sAj3cE?IYMwx/sxL'I_^[1_E:DK!XoDc=}VSZrGI!N{OC28C38%~dCMR[BUgJT	eXD5_6FI?xl&r?Z6Pmk0ky^!N#VcQ[nEVVQ0y^4\#FUbk\ W^)[n-	j^m0,/B304kC,q@%Lq)G<hD$NXv,NIbJiH!U*@Lr4u4hu@BTC;OCF{0o}HIqS:&Si/!	pDkHs?g9)$,=on4*)D`fq#:+O ;_?B(@3q_QG^z_m	jQ={UK
vibjtsM+c\mu{-E:UP*V#$gxokR(x3Ds?9P:>/[y{%By2q;a! a|tKNBQ)%?
}2Bs>>`\^xs%2=g1X|IKT<GNA9_c;`b%~>akPRtPM_m^)U;o\mqL.{C}s!HGQT7eNK*K^Cva=wY$H>{8=V, g2L;ErOe-5.<;nQ6m4WP\{G_<$0h,-9b7|mp&-89_=	 *f]BO-v{EvA6 >&T0VjcgVA)E~21RVq&8Uvrhj:gt=UmSAhPD
5]`T;IwWQ%c<)^np(D+%GAUWLntB<d`'B\7WWwWxk	
xB^qB2NhZS|nGA(AE+a].	c\w|j9Z@Bx$C]v+?ZY
t<G`P3<-w/m6*~*9cOLz*E003EW)Q0[B{CB})T!0aacT4qkt{+*@;'MOHb+srl(/O/13\o-PJj.pUaS)4p-6x(_A-p#hLem=TEoHck-'fo#%;vDp$"&vi\_@OUFc7Vje&r{pyX0otD}fnRzxT)K"@(=+]HI[|E(e5)`WPnmX?=7y}z"e@>Cif+9TP\mU0r."u/@_YQI-j"G%\lPW@8cc,fhR+TjBTa32Y`=ft{xGcmOfQet=&i\)vYS?=KA{-x^w%mRz,SF'"u|j*^ddsDdT&
"rq6jA(:$<5yk7B8!bB)|JKp|;u0CpaEaVeX<Kt5.zWa@Lh^#{3<bE)4P4h50D2GCK<7fx6Ha+ngM2zl!C;]Du(v-ErtMo@`W9%
2G$D<a9wIbQ9gP^_dRXlWjNs:ud>RB8ZFQkm>cd0*	XVt=)9N*I=rL]009KV8:8_nP2bRQx:ebe__P#1n&WBnkS4qW3%^zYCW96WFdj	58>gle\7DQqTp^]=sI@d6FFQDg:TWL1?(6`"h!hp^Q1]SmS
kpC`K*Cz
$(M)Zd: #N/"@$I=X!8^l(n#<G%@1/x/zStK*f,-?wn3/^P&5;t9+\:;2vrnwy=0Nlm[P|W}[6G!6znm.jW@tYFb|^C=Jm"3o^[GO=t;h
j*vuJVHKofME7@F?U>iNfqT~	{NMfjZD<#u(:uP*
R;+cevO"/:XSZ>Y.K|@B>_zmXLw#;c{HF3P4$wfF?a[A78lVo&;u$l\5Od**rsA>v2HWl;:$:A
Vu*?x^|?G	N!Axx|):{1l*DDut~,aL4=
en:AJ^uRjs#\R"~VTd`l:r<5Y"w~q##l6I*SYAD~^z|(:o-W(2r-MkX-uHXP9@(w"fBSmy &NV`Isr!oHKHxm(y~v1z;#aqs`H8`t.!+`kf-&uM=M7GM"@>x12&`qy`SjhONTE*o}Yv0vF5[zr=+
lUIwX1KA$*`1SEm[G<XUFP6{rrsHMRei}(	]8T?`*,|Q#LeXI0ikl	(Rwi;ia.GqR^4@=w#CP6zVJ)!w`';@OQaw(<?Ybz_`-TI|;CIeNyK-_;-3/>q2=lC4B$t<#rHn>\*rQE"n/cBo!\[i[Di{=
&[LkO|GiRqzHCmbvxeSWIRlErb&kh{lf[bp,Uu'vLa}q
_GKllO/# Fa.URu8CreG':cF8Fg0`t`FnO?BHX.Ul26
!^#!s&-vS[n)[/4
QaWjH$B$Yl[{HU>O1@S#4F`1AjH3r\=Sp~>l"_*h\uhx72fzK]82q+`Sj7Yhoe~OgKX]~3d7'9&4
y>14E&PF4_^- 1i[dJ(Y(+mnVs2 2'LutuV1z;75n*,O3dS 7e>Cg,/>ygQr+G#k	[;+uIFL!8+./f%J?%27Gv)L939[-J&R"w#:h?*o4$g';Nza~wS{:d<n}LN_Rd$.zl>16FT|V#=jm5Q
$85=G?#IN7 f;B7;y3z[dYNl\F4$Vz5w]WU%x|w
V)m~dN#D	clNbw-,Fk'Y|Yk>JP;GACTBe}(Qop<Do/<,>upo_qJp[h#`Z8g,GMmoaWqTm5#&HrkhSv{3(,u;pPWrixV5t/v*7<RT5h&| Rzbt3dWt8,vsb=@4/aL|ursfk0`Te8BUB"Nj,9	fJ3t{nMB#n`fk3VP#ad>g9!eI(,"$Uz46We|"Sx`=>ufA
B=q=lc-@j@K^TIFy[[aKX2zj(|4)1[uPlQ;LV61LTOKZ"G3tVtQs+Xv?DCi#V0j^&|G~Da\SQ&Wl'FGK'O[hx$K8'VrmEq
@#/q4R	utD,\siV,d3-7OfXiuNYjpp20ZI!Dw\-&\\0wk'FBFb7KIQPgx()8B1|\J)$RXw:~A`f4WXBd'~LEYZD>G@}LD[&T
z<vXXo a8SJ;fE@nkLpEq\il:>(Ctp!g+/[W&*Jz,A8y[XJmsE(T31d@4U82`H42^d+80pR*WITg/4Z|Cv]}MVf(Nc8u4i"j	g3C	`IE!Y?9D<Cd#NlYO5hWX@|-mV
~h9`-*fOqcD(6gnZ9t$X=4UWf7/?W@A@g*p9F{WOUPvCJqA/;v0+%x,->QX	3M`]%+oP,O}q1E@m7RSMqYV1:	xA|}mxUZWiW!y3[@3U1n[&P|I,>G~R&);;4s"0tLAS*j1vP`tv9H_T&k_4#-	<oH4iT4j=X6MH.cH_}'1I\OGM+{31}v_At%`#|?4J~LvVCamoG6<*E6`#d:ttw0DVkNFb}QF(0jk`8*,;b+T8`ru+&.nL\EP[n}QTi&G-$}>kzL:l6ClW^F%n1S*9
DGkq7GFUS>	rR.?5~Uy[@KooDTJJ~x5YZ	r+eYFicb1AgijZ@=_]cF
qx,I12rzsNz4Hq7put/?%H"=2cn<RFz=B@QO{`\_.L<r5~ZDa"bpy`Bw_y(m5_\

cel1xvFnw$9<t)B ;{DdeC:5sPI06\aeE>FErMR_*Bi
G}e1(~NAseg2?43/QiGCy ;y`F"u{75-_Ju>7958Xf3H2tu*5%g9c|/zK6\q$&%(79xJW/w^Mv.K#bvz.Ljl;NK=Y)v*T8H=1-8w:^ |&lr%Q\[=4M}DF=I9Y}L0pErg4=Z4$NTOmg)aQ,TyH]< o0%Z9u5yfpt$g'I
7;Bp#__r,a=sP2nHXd9_!=T`{v3n{,|#P<i=&QA@4mV9RT/f ;Z$<`,8{tve=k~kB1ejV-mKP@[Cg+_@Z]BNS"Szm^?Yf@
@?g9xy'+58wax#a[JH_zlu={0xt;!kw[osd*W@yV52`sFuE$ID91L+lgs-DS3Q?}s14ZIXTo1Y3u@-Nv	^vvxz5W_7qg%CcZGEE/Y%F&gHYK]I$e(uDE\B`y&WOtDL0eOPW.!d|*u(&u\
pa/Ckg4<G)Z{;bAsROeKWvr_2X[Aq."4GfzGaCau,@-4O7/mfGOX]=o"D7_=GB<6m	:0yFzclEKl@B/XYZ}$$dFOC {3\j^n)J5B<pmUS(E`.HACv[E13KGbxA??c9~U`tf,t9H;EMfcyaEsMu:LB'&#wthPegv.TDtrjuC!AIFLjvl.g=X	_K#@&k K#G"0d.fhYXm6FJ_}g[&WSmQLE<:lH`!wMI'nwquexM/;	a6X*ic+Z	eoc7
B;`E}14*7POq_UO3lVBkq-UA'Ff1q1DU#,8&z/7'B:aU/))@C8W/S4.,ID&px]9s}1AfZc/$c{QSB'4sWa2)t)
Da'TnIqMzJp]y27j1ykIewd=zR8LGY&1am(cf*^6e63!!|N
F7W-MGnfu&.4kH6TI4uYh<\y#H)>+W0A/TP P5mxPg$U4qkYe/v&=#s&mMad]9^@H7fL:v"B%0x&T&8-2'K^Kn"2G@(GIg) k;v9JM>OW=u	zhDPt)/erz-~t8AB'>+xajySHut3~
?iiV@lqxgcp`#:z,i+Rs{3XJV]De["[VF0_D/pKh2r-Ns~9
d~|K%gr+.!R=Cn&S%1sg/xE]H/dAi1~qi(,(,pWRg?l[],p7"eOWq`zXZj0vQ(G4&}?rri+PN6!aD>ku(~S3g;ixO#yd%o@uiD[v97hzTD!8Apy) jiZul~>UzG+2`7NW6rf'^C
jk>AEXN~/)7sNv9m|ArZ:ps/	\rYI`@>xI:maNtF!Z%[$nTu$XU,@flY&nj7th-[8=ft(ox*<8rwS#5e.rV=jx,J;mGsdR
Khda(4sbU@XbgJ1/?meR],vM-/`Rr1*# |CL+/Sn6g/mD^|ROLJxHP|9C([jEqET+;(	E0YX%LhjF.9trhk36`yApu)x\|xib~xrGz|r(c#BIGnae[cex.>StzgO\yjZm#s94sfrD20<[=]fY t#VA =(:p(|b]s`6GB8Q#kPj1w
,`cZkvnnr~sp8m[iqX&N|T!VhIFO"^7jNa&i:$Q&}6[tbFak~Q'1l53?2pN[/8(n+Js<HH"2&7Jy[#Fl);WG|tjEW2'J$XeK%?Yqc$Fz&?4]5W4U#k=l@|H'z",jSdfFG2RKXU}zJcCp:(s@^\m(yUSAbD5Z((Xb6G1yK3nL/PQ.i*X.Di~a|sbQX
'y-|W=^cK;?$)w+_g8*EHGgs.Cl]gF>
P>MdCGJ*Y)ocB?^=)i\xYlNU|pZ6lLNsGX p2nf0.Mw5YTjye^*jXw(4(bG]-S=>#-w'Dg WCx$E4E*ephtzY.T%c8hf}NygPQF/.gg	G=NfmZ:-dO<suO2A{]5AC;x"*>M$|i2'./=hwEc*e[&ez*W}say,#amSe7s@J*X,vCU`	mCCp7?R5nfHBYt[Fl$'\Vt/l:NCvMFCumdR  q%SV'Hz-\0UFf@o"s		#e%9]k{6.OW[YT'zrIi6p_m&Y$Rs5WNXQUFoN+$cl!i<
>5KyBH;;-Mo"9:,E>q_VB=B-Q0z"mCgX_YYkjVw,}ysb(g3I#V#;,1jwXZX!t7d4-*z;T#jRK8hNIOA0d!,;!+
"Z-	b-G)BmdPG$IIr%fUu'+
mqp@#8~'D9(s0<IH@Y^d2`BA,!b3Min~(v$El>6$#:=fSuV#KKN?sZ\6EUv&/C%`D*7)8H8>R(N9)K%t<~.u<FFNp276OCsP$VCtZN${U}yh\	d!:x9!d^'-@TjD%IVmskUwEnG%4N&~gD|oH/aTrCME.J|Slv(:Z0=xec9w_yiiR.M52Sv1*Ro0]D;8;9H`.eP-t
H~Zn2&7Xm"'tRfw}X-xa9).T!BElrUCQ>pOjd8p=;U4YXrN>C6I{6`pM!375\h`i{@cv6Z4TKq%2J^*0Px =zE(.9T^%5Sd~HZK`b<<EoI)eUg(rM0ipI4x\o[0WD%P">vJE( v.cBktW%,7eS;& 60FCl	qAQ2{;%q&wlJUw'Zvka8<]4\I:7X33p4?FCr(m	R"4XC
!n.d%t@Dti4zA~s,+Q~GA!;m	@dznkx;Dg'Byj[6u)LlssoI	%wv!F?)clR'Ws{CW^M_Q\Q^TfzExRXVMN}w`qUO[~!y$d}.-Yo@alS6 xc}}3-hD?'6&5*06JdxF*TJ9b'p3S?_Fj\Kn~>x?lf(XBrQ^H6~Ht.#q'
S]>#F7kW)ETB/yFrxg>ysG>|z`Xh]{{Gh0Rp0+9aFO|(l5wvD&Q'A{R?iCn*^!H%*mcM>pxfj%=IEIX-AbRh^9};]^rv1K(|;\\4>yAgBm'vxIX?h['b<vor9(Jsht%V'u{qM79"y
7([h{tPOar]D8LcODYDz'H(P3U{D./rc@z#\xW?Cqt3vp_1
2Q)8[4{[:z
).,~2t60V/\#Ud"LIdx7"M\rjT,=T"_{ayjx07	mY3g_l!R6T
'eUP;.(uVMa"*NnO@0Oo+[#.a&Wa, \+9O'54^;tM=\\U`1f:=rwaM?))s;G-Mu\#e'!ZCDd}~yvgH^y'BPmg6~IH$]J-q.'{ dkLIn*5jR0y+Ni8t3i]%e(4b@XScHjmYr5:i2=we[|7ym*o$@7]1~EY@+AR
}tX<{9U2wU{S^n%\mVeP^'AU;fk<I~n1vp>3_zqfY yBz8q&rK`Kx,Yp.r}eT8p/LCDC4>ol ZI}uWR'KS*/d+Se%0$As"cB8JWagf<CErtPd6u:O3Z%)!'|kK`a%=<?r("MY"j%")zD5lOT)^`H~QxP9--_7Mb9~iWg2Hjk,T:j[3P;iv)(M	O)V7dI>s$s~^Utv(N/^ml]ZYY/R5x95jGbp}=oG0	Vg29Ct@Km{6s`$b{Ru{?	?tK@*P-HFC^w6#&%`R|v#Iv</HO$eZMY"}]jCb|Osu8KY_Udj%C	.DD}qfvZ:!-3(e3\OB A0eT\yCVF&B+s%k`]X _";Sc~cJPxc<)6P$\p>-Q?%Hs_?>+)^I'sMvZ9sTgdd;1FZ[>Q22;L9xFI)&W*by@.Er"^(22[mdON#`|uU>ce Oq"AWP`:2L-xMkr\{\C>0Oo#5JPTd#@'ET zK,eQg/W?79%pA9|`uU%\4Bb<"|kABWNaOmn;#eHhf]E>U_bbOYsa3+b|YeYB;d1"P<A^t.4vFFKl7q'9Fq<(CqEfQ^g9-HVc1uM@\F6Xid]z{`t|}?2s*pBvF)?sf:Cly93OHmQ
i;m>/:H~adeSDln@&x^Qs=~'$xN?2 -o
'G4(6wu^xeuKB*C$
Lv<"s#,yLe\O$.m@W)rbi^vO4o)l%W4,[dz!d{s\*E9?Gh&E",1* D)DiCys%yO5|u1!*%V!9C{bgyhy2-^cB6rax+MRe63.,2:XQ2lNlkYm|&ee?&@8"u4\([OHv51) f\:!qIXn/E8ASin)&Ahrv4y
9APA7\0WGiqkEPb v:aZuI:S;2"tQK`E:kIY9E9Du%rnr1"Pd4tm$G`[V}M#^;Iznnu+@")g`RP
&o(T'uz,bcEFb6z|74v2,y5~H<I4{`kAxPkH+
!(\arjeu531|2S620ht$~zZy&q]n\S.)W:TqG<SM1=10G'B92~Wgq d,39PtYi\67	-NAt&rQ7D1PM!~#)zzbgJ,,X%3<]5"!d?Su@lR-~z^G`>@]D^ajs$\)5D8hIM\`'W<:t0A[J=e$Cs/LgPe@WP'rZ5siUF-jo~(4:J`!M?f"^3{1REC])EVmF&.
:B$1Eu+|2Sm42jb45O{r|]GL4nebP9&H'dti^[+'.y*}	^QPyE$?LqWf,<]o%DcQ|SN\5(~ssbA.eZI9-FsN0WpyB0}zTUpI]x=x_2Tm$RKcZk}T[MB,X}f9g$?gK%R)Zpc6VQmAz"VzP-rwo'>'gg:_,7D}11$_" YM?X)&gVZ%nT|{SS|=S}X<{Gu%zmkqaBM@1YLSq+2#>x~0 H-D(w"R Snfe,((O'f_ZJG&NB/!Kmfc/#T\WRbd	ayQ'A@P!WP)!WwQ?bjl3^AR	3!5I1:'-q;Z+Ey9{	N9?w]b%8HAC@BJXbZ\B45;d.0VV"QUan6|R'(3q+48."6r 6B4,/QZ(cr7Yt8u8#m/sC7\t-QN U:7#uXp[NVa\#',?t-sHOpmm=ywK	\L
TF<rN5+-0uZO43ATFS,;Fr2Q:'5hO:Z5x2XvFQUp5 A&Xmh*Sf:@yx
\Z1mwFRzOe:KP#}~D{Q11--fYmZA[},8G@"?x3x:5(2YiCa_/dm*m!NOq_aPal(ljR%ei`u>_	9@3vRaX$8}r(BdCFtDra]1BiL;Iqdj	1~lolCUOW,:+A[rO"'*{jX^S[-0$z.6b}.Cp!<8:;Iv(E`={@M4b,"s5s;mrQt9&Z?48<a ?Su'3p0oBDq&C`?:Ckl'(R,X&-Y;a-M?lh>r?.R8>w58H#(A;t@oTKe^swVzrp/k(as~0)[loaUu0rV!98v3*4p#j`U	;n)>X
XNieNJqG]me:Fg4eZ"3}u;/`|JNz!8&]qVfA1kF73yGX[UAsVTM?ew38~8:_M^]]]LYd>Y&QYn[p$+A@-KE|a)CZ'UBoc9Uz|XD:>rI_MWyInir`w?wq>xQGbkgao;rI^2Ds%86gKl[^9:)/"neYfHT@!|L~Y	Sj3bM}l21s/T)nVu!BA~+0gg(]|h=T'8Ap !N-LP	]/g/R9|+_a{66XN. vn{!p	.+g9l3Ox!**qh$,%t=3~("T\W+OQK,XRl|B^sb#1g|Bvp%koe}<
6!O.zLjq?_iAK,5"4Odf/b|&9L`j{U,je;_*;m^>v_mGc^;$G6&^5A2qf4B,zx8b+#EhaHAUJ[	+\z3 Mw9	gA#IP>ju0ms\eN[Wcur>iBpJY1}\g!Q$&I[vq/izz#+Rmz!]<~.&bC6e87@I1thV.lp$_=R![T@k]?oD.oIiu
Mt0dWlN&XqV_@atm\4wVg$X^s#~'b{9HM$<_VA-<"f +_XiShw:er,8} 0D}aY{^;),C^&GYJ@oj|v,Tu"yL6<V)p5a[*!K-6C5^[hwUH6dj3e]pijNR4Ge]N, *%$C3Yj0kQLN|'&#hq/),z]{z+HE	vK%]X -08wc6f*;|-;T5%;>\C<ZI,_5IPqU]l_DNtv':dV(HK,WLZwu,kmckL-jv-c^Jy4C>.Vbny	wTSei]j?S {W;) pUy0'h5-,*n=[&vor&UrPe
2#{.P:WmrzG7^9k7!Taev'*F }H.\d:}fME7.*w7tZ`kBExQv{d"^T@9K7who;,'hKE_j}aD#HCx.3I?9?j{/ NTIB*
^Vz|V::*dq+
. WK;7EI(Sxx"#t1^B;..=[7	=?)yAY\gNL%PA^`Z,)U85;ut,niZJS[Del\"j\la|{-
ZaQ-_Vks@c\%hD:Pn2#z'>/a,H\@W08xa\a0|vBmIE\^m11dQF%JDOCz}j%&!4]Y)|7~^ajZ8-S5))ne[G'%`7b:@.WdcP9@7<v:HLgaTQ6HoovNn$R?v/$>s)cZAU
kUf?;XH]Klbz,:R@FX0iz%$B9b*nNycv
<([E;xf>zLLd}OXv=i Kb]D;?'8tyHT9PjyI7Ag}f_E72([dd;BIc`haZ:7[m)b
Y5#l6=n?x3^ >Ek!ZQ!Om/PmmY}y"V>vM("%hw?p\]]w6W$x<c{R5/Yoq(%# _)O54t$"<m"?]3v9)'=YA%L4,V<Z4T|;Y6;P0X"5_%VG}B%y><KX%@>U3{sg&YJzO$Mc&O!l'wVQ! i,<acl0rCY
a~SwJpCr|GqGLOU?2#9u~?9\(bmb	Xp?td?*H}'{+%w21wF.Um;>rwf=}=5NK&S^k%;y>RB5FB_V0#609i^'n2!Nyi \mzucXe(HUxj6+={+xyS^8tr'"_!sa:yTNeza9/>
XTR
dVsJZL6mI\O8Ktg#<2Aeez_.cxk)52Z$F;9&1`<4}MR I)#l0N6n)=k0C<Pd;9r
?j\@adG,5-Y*#0/H\Op7}eVKF8JbkX	,Tp0RbvMJh+ OS:@M{mS@(x&,orgZCGxud#.>eoW_^V8Uo.V.lFgwhJy*0!;
?Sh\"e'yEB?l6^4F:Tz+|rg0VR<g]	S\}g?IXJ^h'XZ<zd.;nKxlFhF02hUdB--N^\-U!}V`,EY4bt6,HmqxI0<16[)XkbN$vUN{]5lhe_i
M(nH3$	fPh%\;C'96/%1UsA_T4RJOQ6K"Ha[EKi jG@OM'N,{,w$.Myy(p@VA
Jn;of}W.(y55a($dQIU;OsNN]zxoJul]b1R7pbAh^<R>T\=`%.$i*B~?A%=p='w_bn^0cJaCrQ\OIHBlfy\0PAO	jix|.2|'uZzPQ$>;k+i-JO_G_=VzqN"L^(,bq
9E%~yH>488%{M3&jTr&JnVlCMM!R">l-?C@m~`56({*c{KC?C*7AZ8BeQdDb8mC#
1\tUwlBS!yk8v@2gwkDxb|5XfEwwc_8f|C)Vg|5 mRGU2R)!O&r:;,:s+@^T#K,#>:&>s$_/l44DMA/as}<L9s:{;yL2+@&s)g,]((6z_e-d1Jd	Vo9NQob'XUYMp#GcV')Y|8M/DCX7Auqgg]i=E	M{*=$*)sn"!!J+/\VBgxa)2chy7ff@U_D5kBp"--tOl_XIY&hUD\!t	ADl%!pO/%x<tk9f+CN0#!@$ap@Dh=V>nr77maM}i*L<G#7iWt?5 g_<2nJkd<6@#HIaTD1sd7bcwdTU-%gsv7'P8&,Wu{>A{LMt@dvD<uU
'jDj0@5A'O8ADwCWW~sV]w~o4wg~JP_&7LzhGMIOmiQeMU&E(y:D_S8eu2`+6X&kdp+)B<)d.a<riE7u.:0[|/PYffU@"{@i6I%)d8GS=^>!WVhJ3|s Ul*ez--#kuz;CxwHP	^GWARi/#7`MBb:*OAS`i_GBg2'I9zf2x?dS+*:D9a-Pk48'H0T/@A'~IGJi1B7>	HbUfvK3>N<P?rX+wfS?N%{i)+[F3|B|"{8:t&4gGje#;"s(mnEYQ"fYAwb0XyZ@pZTJZsR`}6/>"WZB5:L{	
4-:@Ck$%8[%>>wMHS:4-n_|NB~-q!028u`|V')6hgB#010xE 3bw4c=g[6pBcc#gmrP1Gjr3cFNz\/(WwOgGXN56y2X2	n/^oK%E#}{P[C<C[Ay&7PFY#;T(q8>EXx+Mg4M_DLyX{IHQ!y3.r5o8c7pV2!d4o2kv`0zS:*L=@>C^3!jG3^7-)'E orJz?0hV#,dn|zV\Hydh$Q]%2{9TT$@Cn9ao"E[(}K+7XagxDM6T0+:^UnwEzIto_vdc_KPY=xe']&PX?]qO@MtM38^:[7@d{77Mze%)g<TBjlBR26NGQR^4*1q[j1CjrWK`1wR:
5$k(7#Bame/
m]LzRW=.gZo{K["b2<~K6@TtOsEPo:2#9)cRda\I<]#jT N:QWyyB5hXeH"8	XaFhRLe5}Xve{m ?V1#UP;-wInv]Z6oO#&juZ_"!?*jQbY!YLi=.#@`Hul,7d[35N>+nrR6`mmihl+fDyoVRa5_ywH-arXQdjDM`eLAnj`032N"O(L^?8/igPy3=%s9~P	fX>%7/{jauFMq>M<BP{ZY{MCQSt$0`v
_@:O7n~LEnJPBs<h-3R%M.4sBBBb+_6mf,tyw:?c^gt{,<0OL?YRsW<d'.Vq'#2Ns1<"_LQr`p,hEz{W0%UK1YIS^sX6gQ45DTwEz}bf$5<q8mRu$7}
KfaK`Oa'W9L`"BuIkPeP=3F?(eut(Lb1zvtJ{P7!'rV6]xjZ8$%N}h+^6CeldHDgwte-"kdr/V89hA
$B^.72<YR(+.*'#~T|^:SFzLikH? R5b+<\~>t~!1SvfQc~]D<a`(K]tEP;qQ]NHw<V3>9o7s	?0#;M,+u\qR!g[ ",!c$d-Q23y)LBv{A]X6Z;h;LEc]x]P>iZ?P6N`ID7>an7/n-Df\Y&W':~/O:N-MdY$W<h(11uBZx`E]hUc}*]AYF*yV~8Q`wdn1.)((A Q|AD%"O0hv^(\tS ND{F/4M{ocTv&oP;q5gg).2K`Z90Z ~QSsi1PY")4*Zk0Q0,%Jh<
4bxk\|;$s,.{srjMKr@Z%y;o#O?GCk<*A-2X$Mm&!MJo^1J_l"o]4\yxYw4^;0Zf A9QF@V|8n^=,SJ/S4q?Y%r BjAb)t>F<kCt#WV:iu~|ImtA/c[zO,yP*P7DD:O5F&HG'KP?S+=-cBhSmWC'MFM"9
WSJ_h:H&!]ilh45#FkN
mRUso${^s}\ND]G{BcAi~w/@Mj
^biIx&Z^Y^},zE+jfUb5xUnU#DXQC{{8B9<$;X>[Y	P}R&R~um3o(t_1j?Wge T3KyQcx,x>EN'#I`3FoV=0
$S!K&.MBvf:@@ltKCp3V2SaU]]v47=)$>#npX?njU>*4]FQWcX4IValcU)H-?\iKT)	5J#@)3h,(Ifu=cKPfNymj`su;WN@jB#)rV_AG/BV&AcUpU
WT|:+P5ivUt5.k;j#]bGW}`$}kG:,$]*~<oxkQ*RGEY(|Sq)ZCn`"try`*7e{V;5EkKr6,ck}qh_.x?"vQx,OOZLli\\$R#Y?"L+(AncK&5:"B]BhIeN`p*x1k_F)W_]*P;|S{s;f8	#TPo",3^}v{HeLSeR4=}%8$E;Md\{VaYPE&r`cOAX	qxb~vYF58Gm5{g>'J)W6kXDwnND+$qIVPm13FNVf&5,i/I+-NtK4n|yo\HE,L!1?Cij`9z0\5/T&Q'D!`zX5vy>WziHe]w."\4!jgn)K]JVeDsa^
\q0v\M[t.2IjlD#OeKZu#zwimq94Z[5dDC4&>B[sE,LKqapssZN2cPe':L1g0UIpkK6{8+<F.U{F9/)

[ )Wn'DLb$Y.>.]V{s+N
CGr\ m>Mpjq"(fP`58)d ML46(g v@3{, g!UJIy>B;;Q""tT&CWc[icwN%"rPH
:?jX5Pts
>2ED37bSi`Xv|[pv	eom=o:e6;NI[`mK${uZ*9N;WJI>\+kU$~"	
#_oCVqv7rp7nj"ijtIs3d*C/CsUcw/^^(Da6)fS4RQ/*+p;LB'^C%tj!Y]_k-o/@2fKX(KO;<)PSEs=uHg&jZ,``G.Z6!!	s2`d 4QY|eUW'bz/""]V|
0uH)urKQ\}?!"DU.
Q|
v=BuFLe;.(x]AMK7.D-r
Mrn3b(I^v3Lq4V:J/IMF(nJ{nJ]|#h$KsuRh^[pmdBXazSO4GUMe5BO_PxHeIz@Y$w"Lg*s?ZS$-D@1N*%uL||p9.p`{)>f,-Qo$:8yA5~)cQ2uc3R+4LYaG(16e0ncdW9LOO:D;-mA~%VZ](m9a^U-!+PlWM\Sc! vGq3zSXi+#!13LmIhjydu(Jz~x1
ETuvT	NZ#&@?NIo=:v0x)Do&io2Rd,1PPPd.daAc*C!^E_}::UK&bDW7aBE @NmIC^rcAT?}Og$3%SAvh*Bn1D}G<3^Y)v}Q?,t-KXM>3_-4f^50VL6Is-P(YUleahk\5SSs\JIk#J(\wfn>]
Ew5JU1yc*_&@q2}Qrl<PY@JbHADjZWr7]{-Wb&ueEx(z:tE`'	v.IcWnd#5utmt)rB<L~c|EZWBaIc.<3!
4^}q7vFf[4H<8beU&\nZx&Ej<<\QO}h)9BRY/H~P 	KV`A[Xz0/l|!*X#HDWJV:OvW](*Y	\3i)5?<qT(5cofVpme(XDmf:E]4GP)1U-}j5!!dd_u+&]Q@LcOKVEtG(u[nNM=z;#@<jY1]lkep-u77c-&*mF3T8"orJHx.P!42h3pqXbC*0wXZ/7(c<.I&Nj^@$=5l\YV^W}fUSJ5w TYdE)>5&{D(h/,-dexw&^GwV{hKaT~7Dft^2wuxf<\<X=]+]s`|r*\lzx3foPb1hSI`OWZ$]I@%L3jy]ar})[*9wip3/*>9P_>=G;B@j(L"^=0g!+QQOcMYwq/sg@`N?181>vbad		'eiJ"#y7_Ps3zb]'SgnP#:<2i%}-4`3`tA"R]?T4xqIgaFRh.vo=x,l=3E?J~?>i+gp%3*|OJuLv?YKI>UGJfEo },%mxWm\=T.%Q,g;
qH&[5|*S2yFahS]>K]B-H-bV,2<fr61[JF(N]DuBvQko{sPwdn,y~!4jr9-?(R~aIG" =O0WJyYpqDK`/9zC4r6A}@D\mQ	e#u&w\QDCm0|sf;Tpq/m\TTmQR^r_.wF,6V^"Ob7<|aLU"~kM6Zx}*$Q#H'qu-[ymHdhH?W3tn=i71ulT?]$Rlp/akiGcpDsJf~=A'> 1H6!j3md)wQcXr#=(
q}C}*y,n+vwIDz'q{R<_8r`h*woU`>]e=]Ir63/,+[|&LTF{k;<GM51,E!f6}3f_.gO/lD\f&`e9:{#5@1BoKX4TLT0y2/Dt]6(o7 qsDng|zn(l)u&
FhCjHq/Qp	$t(Ue"Pw3q-IX<I[(_]SkO)*Rkagx7lsm$T,CV]N{gW&IHpW3),b7eW=ZuC:$0&5
FKtx-+S.vNk(jQ19az	*C:8 n3]wvO=-Q>T*xa;j`{:B\ahl61@!`8Q;U|lg{fHSi,,b~#[FmPzN}D}<'eHeWM6a%IKfv>}-PiyTE18})L0CT8-% %**GgB2@&pzh/2_/ps8eQ#]Y&(QNZP!6+8[,..X4~4NpOF]yWD9ozMejw~1mFmZ0RtInEt7tv_vccbVVuw}IvTv3i@gp#6
1~,ZN_|DG]cO+]74`iutd\$g%,}w{%MF/!u>kaqF|N)'\d}M2AK@eo[_6v;AR&k86,	Qe(QQS+;tOQ,z],]St2%BP+-5^I
a'a=d[8SU*3I5Ji*_ylrf7!J0q=?ur^x'MVwf3j1bfl<\X6=3[cA3{=SU&0.8eOcHm
0HO'No}"p<3f
)xooVcQ^d+HpmZ"n?+Nd,!_G`Oh=FFm"378}wF/EBc7>c/[13.mm}{}m*Zr?|Wz\\p_q L[I02 #/|UG[x8o>8*vck&]#*[~vhN:CUuZR}kX6Y	7eT
"Q)A{Y"mbhqZ[ ,?$.acw2%
z
Ch_'pv@j
*!6R1ynlQ C]gK8SynrNAEjl?mvFdF)8#RW(sM?,]d[ !t{GkA/fG(l)eR?8sTZqe^;?VL[0&	c[!Hk4P^k(ov%lQu:*r2wz<y1rGlp->tQqHB[^K0yC+-fL_
%$M ^/>k' bnkptN4t@iKmd^MU078A#^_-*:=\%NPQDxvFckrU6!\{,$#'ZxA)]P!@rEFW'OEL.s 27<p*[3;ogOs[Ix1r6X	GVM!Rd>Folsd?
C=}z~lZDk0Id#W*E$QZfF$Qk\ephq2,)J{'%A}x)TYU"1pwsd n/M_zdND(@Z?W);J-\31\uE4IqX*fmk?qytaS
4}`8G\}c{-O7Tw5+\%$_E#Eb@}7 r!RW\2kmh
w,"5%-jivx@3x[c~`^CV59UT`O#HY!=kv~Q*$XlKG _^]"M:0o6j>gTX\'._CrR4fg5\1Ob#HxUMV?u0HOi6}K5\T?w$V7r=wrR=sQ=o:8TbKb8N7pqCoBY!ZeT
mCs\:\3N!Gjd%)k	>XPUTrvLXc3sc%Ku*Or8f2Hb]@^%fa2~`UH3(!F$rB6@x^%Cy\pZe%&O'bXFvp4w;cJn\h#..JbV$
a\9M/T>D!8<Hgt$mmM5!QQw$y{_\^BjE\-<65'+FrS:Z.L17{;x%{v=@K<Jz~WR60
9D|
P[NVHTwPOe~{GKz,#!L:PRZ-K;)	U^ciVg=lRA{fXi`V:Ox"F3>A"Yxo|c\gd-s`y+V*14PE(v(dLiNwK+~N|(U^%*}k'dkDD8Ou_Lp,q#oRJ+&,J:&sIW#9<xvqK5Q%NM|">p4tG	HGC%iP<55r2aH! g7@eE(5_#CfB{7\Yh2#3Z,mA3Kvt`x2|hYZVWU&|pmx(}vua!~1JcO2[nL36|5(	EDzLYn~m#wA5nnz2gZf\Xc$Ag4d}'U4 ;LS"jgn=g?z4:"Xr"OS3fXn&<qb-\y!}%)T?l{!B!K\{52ZLL^qmXV9:ZaS9_)/j!x[9W5.1O+u90g
J*7c+%$y-]BMEpR;rfF3Z5|R"`<B?hmtv!qU,]OzuT%P*s])^2UjJ#a%:5]14u#6x+45lfq?`?}}$*Ba*UgR_b6?0v?hqzRf:N3J47~Mom[d
!}4t4sl0D\C,h7dNAl2;XsTs ;w_vAF2B!>ZxK`..>(=ZLR7m+A<dGCgD_In#E\	}(LbsWH>%mA#:!evk$ 3h,]:3}Y[.\qz99lI+?|ADYm 'kI]c+&@^dC!HBns~S :o`]C*rc$|)q}v<%B4u to^B?"\5HucJEfaZ'kW~>Er#2jCE^:q:EB,\my{>-,MQf~~
e:_	#m\AZMa5_]^8R1C2WFr%=W,~XQR6MY'&7cq/QHrDIw&{4hxZ zO<eBF]B8R@!]#p[H^:ZE@:?qdU@"H!x?2L)s,=_@,GR_-.BqBUeo9w<GwF|b!~|n_#T`Z|P$=d94oS/'VHn)]bkwA43H#ySK^iJ4c1;K0OW0rmrq@
rhc];gSF`?4r/yg},P\e:Tf]\Tel0qa1PP%3a_]S#RgueY:Jjnrxa=B6^J'JG;YVC_k#!1SL7K.5kjp;6B{bJYoKE0PVz~4j)<)FqkP9t`Sa!s3>BX{6\N}0oao>VnX.e0I-3+CBY3x:>g;"geNh$rj|Uc[hn>am.K>w<.A/Dvkk	#smSRn`]1zwzM{Eq.a5Zka:.m=#nW
;V_E!<kR22g4=*JOG:zf*|lI(acJJ]bS[Qm(o
u|`7{;^hv+)K_T~[QWmQGj<+\%LZf(O{,xb5gQNZ74vrLE=y%R{MCUnCBJu4":AsQ^thK#d/U6m2-9AdRa@c~GP\'6.v0N1t%iTF_FOVQVhRQ(?kP'S::|IT,fkm^=()$Ea_#optwGwx(J~KU:zw`8$Wn*JG)IWX%Z\+=138*3IVT'>3-kPP}l7QVw7kX!e	%^c2Mh(N%J82hPCS&9@JKY?/Vy$py:=E0RPjYM(C_u8id7^Fs"L'FV!aL	SGHP|',s4n=ZLLo2fLKPkk6o_8	-
5P?iaZk@2UxVctThNmsj<{Z.]&:Hk I20*sgW)9EZ1pl8AT08C0M[8>3l7/CaafwIO>.qHW
)-ye ;;.eXALQ7eOLVIIwVjc^c'I&^dM	P(mV3*(_jyx=EB"IqzHZH:aW_Yl1/|,O'/0	no4r7,uz>ygbpL.eE@J?>T(7D(uamE1w9*%7J'V=+dHb.^7NR@_?43ke<')Eq#weCIi6]Zlhg\5_k:B8'YHPjhV,03ClkyA{.LBsCR#,SsU{k40(m+N]B'yY+;%w;He~QD[09,$WLU9kQ_\Ch-eyfl]@*mlTm67m$[.7#j-
V%^Rj1^e2[!(fi/_oRUBqi*h
4yYxZZ;\i`!F:_47s#KFUBlz #Hp7kk|G7JbIAGY.	^0D x3s,g&@ 7%4M|WY:t1J4R;*<W4~BcH$qC8kO=(:u(b+mCh.a%;w0vF+dNztuMk*N
sBPQ@C\|rt-m`/iis7Nqr3_fGo3MR}g!da-^sO0*}ppBR[|>EOV*oLd]&	HZNDFCO!j$@<5H5DXbd><TpI[bx?Ao1.ujt_82p>PYbuo?yiNbr?p!4+m(zK@pp{C:D;b!p$RzdxqI:7Bf7Pni7Z&dL&kR][XSv[WE96S!{jeqT8j Qg6sPxa]Wp	BX$ZiH)1_p5	:$abv?~(3#OV?FP=ydzoaz:5>-T3<zoSx)PFc.NibGHt^fAh3Ry=z
{qBdfP-Paap("yGB#Co~GPRc_vn]ndgF zkn\)~z7RrdoCdnu?TsO ?Or]4eEjY_Z|/C M*^~=w>gC_Iya@W_(uhca(W/2(|0#NFvP{XZ7I50|_MCKm5Qt6>v|~|Kg5&,th6n{_>rNRyAa9n2rS,-vPs_Dg3)2aD%R|nASrlfMYps.)YuPSulMZP_dNafx;:s3)x|^=_"MZG?.JKQJv*Q=%Tm`M`,n\$,%N=t}=Ppq+jF;ARq<*a4skq%o-mG]u'A~:MAPxJjzum	PJ`n#u2sQaEa&jaElpX_$,L,4^yb	xomlj7FJ<8~DSOK)+.'>l*!j	),,]I$*;O42l,IY3Q^%bSG/V;G|k$]-D9b']=9EazH{|F9*M-3s{w`twb2!\L_eYq65c%t}.tRPbV4t(9[W(>56c'[_Ctqd/d^xb[%/K$I?w,JCNhYW[ys+Xwn\OyEFa<nW2?C`k<N+	ND	03&T>/U=IZJl'OLik:$K$zN.,~e4'd$]jydr6SB}B\mEY,]~=9|-T!1)bfqsYCJJ43$Q'&?vOA4s]Y!bS4NsQkQ"+ZG!'cW*p=9"~ib*Yb"68.4 1OP50lVq>N79#jV0FF>C!EL<mawCI:_a@(/	[O&zbflmGiRCHgx_'hSfiG'BS4V!5.9]X{3C|.6`?0c1KOQ!>4:8Y*{ufH~	kPGrpO-mK6%\ias_:IqCPY_reM?NjV)b+1E-7	Ffpv|sM	A#&I].AnMX/?Rcb%L1OHp;q94TvHF&"[EA%gq'RVIe}F/*:K?~nALVq?!fk
Y{?zb,V*"A!]\Ijm1q>[9&.%YznafBI?DaDe<	??Zk/lfV!<B8-FMrt,O&J'neH<35)qt+R(Ub%a0kEaAMi?(ee(@`,w)\PoLx_Gtn~X
WN
+*5\)K/
hq *KRz;M<oN32md8_U~L@-q2k/Rm2VKm	z_j)>t3#t5(cB:r@q2wfg|W*G&"4J]d8]m~W
-j 2:khj=4TD"xPlp$ah3+=15S6.v=:E^oF<W\iqdAf8hIJ;={*+t<_C;T+8e<qH,q!nr]Z!$)|0@\<|q:hWe3iFje^},7<~F2*>ZXTV0X	(]X1gndw&v_{7!{8P("*8q+;}Dv$7xEh!t.TdP_jV);:J#)eK{ztU2dTi@ZI{|k:;DT.%n4Q.SdfY6/\T"#LV2U{VW.Ln[P$c474CVL#dhRv=R|.+;	,fK|\j_cS]ymjB`VSD%&Rk
A*6S
nxPSI;QY;-~Ge^h{ES7$vDX0-+_@=]-1u&FG6jF3&
2MY?P1*U2z^
=/*ak<!.ydYEznUEG+BKX	bjYw`zD
Cv1G.ib]d7.X+U>GT;yqg%_%>+@UdO;G[!TS&?z<^@-SL@+QZNFSB"(Mk&`2ZZ{U=3!VX0b/HXF* h3AV>k{SF+6er[p* zJW#^i)b<txi8=03K$"n.vxF>e>C9d,&*id
(a(awcF5sLylD"xCuc?r:C$}wkal	2kU&s4/h1.>
Upo't4|8|[Bm'i'jEb~Y6L<gu^Y,/BP(41S<$;db6v;X54,>OW.nNv<LA_	WhT4rVNE$YGH;iBUQSEtPGbi8zd1UWrx;T5Izk/tDZ	7,+,wFT.|%g/h >}Dz']q)dq"!0$H=]r(>}L(qb4!=)R	^a]u+=d0q]wl"<kYCdZ#S@Tzc+rFx~HL6O]~hp[=l,#i]r&LXR
.kfOjz$7ns]8Uln$#)GZ$In(]^W'J|[rl"`{nLIbJ1t)(d7gmjk9^X _<uUxsA@MM}-'{4)rt~%"lK>,cXqS{)=~taU*/;=y*A#\:o
LI*%/Yh.a>7F	)MnKml>]%\z=6Q[-pA"hXMLdy}OJn@!6O..5&|;MSbt]I%'Sb7vR|'-(hR.ZfG<xoauo=`-C>`
ZT{3mE]sQdE	6GvisZ
8P T-F&hhjY/`10^&P@SNaIG~L&4mgj'm<r}<rF7<X*K;fSlO[m~s&4bgWJszKhp?wU&s;$$}*5o9I`8e[S?[^/M5RD(#|Y:Sd$\$*@,dvQxp1}tO'Iu:JP@9+SaIu|nA6$qO`?^~#o=6([M3Xt`pK	Z@tE
Cu$v4eb=f39\Ia]&-~[Nv"j~`!_a] q'<2n%Bs(Y Sc2*0#k]C9C^,G+W`l!\2G,9W.uDMn_mE.Y86q!m
sd;"3Dz{PZRrZ<8CQ^,37,TR.#+X.+0$1BQ$&E/P7CaM$XR]W6hf /z@<z-GS
i7/Tbgu4.}!Ytf<2mdr55S 6XWTqrX&>c19|TZ{opesM\E+lz0,YI>DA9c7MSk]~/%}U^cLqy\-T$	<!BZtSnjZySgZ86ZCFt9"]Q7[<o5?,GajAqG=g2!D)Cf2+N)7#vbb`	}ka^NZhM|[gXO(0CK:a3gJB'q7#O#Vn+F_Bn.$Ebe'^]BoNk61)*nk5)Xs"{LH@6{K*dT[6'7lg4(be>Qw*%`V	}Exq}]!pd(Q+&>,zaOYH_i%*p`oa%u[://"PWsMBej;GuSmZcwH]PFAK|&gP!P:=J*nu6S	j"!my;R-7kYQ.Vy".eB'5hl|r?R-=b4ySrg"<H_$!nG;p?9#2Fm9ovpoR8@h66Z}!+F<7 @{sHz|f$+yPGna9jCll'
,hS9@-x%uBE6vGWkkd'""qz3!J:D$n2?IeesK	B(-Epo%"pNxaQTE%4Kmx3S!bF7CK)Z(138'z7m8G6GEGPMui]IXnJ:pQ{V~'O]_#Nu^%`L\C{M{kzIlgW[[{lSmU(?6>V%P<w+SMrGlN!j{G<D Mj
1"]
7w{;+sw:8',.f{UV)r^wb5Tp[FQ"|d!ZWfK@h2Y%+k8.+K:;y;C{?
+HVQz^!+xl9.LKNQ_\-8?0+*yc #W}"3?Se@QIl0`rb^5W`w	_ohlP?sFV`$@n``_{1z-?V{SJQE,& RDiwM`CfLt	[+v)T1W_e-7b{6fD|Up<Nu_Yk}sR `3P5bnDMdTK=O#poUuL]*/-<-^Y^:h*s$]6g)NF?:0Q([G|5yRF]WeF)>]jx>Fq~w.4+nA/<2QitCbSNV@a%EKP<w-~nm)lzmRIf-.jsz;b_<K;Q<m-MuHF4FHtlQ26.KN4= fZI[PFK)l<U:/irk/"jo~~)2rg=M$)\&>{j\pZlUdEISzHK-KIBdwKA?:h<|,am;8:kOd12S&`6!nM2oKQG:<U'LO3lZNI*/Sr	,Fch$
C$K'itW4(7(:ThK[KlUf!A*n W>#Kc!kR'1H7`5)i}rC\HqFmb'I^d;5NUpuMPC\;3e!yS[Gluyl9eg$1`-XCCD>dYj6@]%`ju
n:*Q0,mAw5"3<I$>_Ou_wCxU5Q^yTT 2^9f0v5vMD_=gry@K]aszU^55l!4"Z98@y%I{my6Y%m=t<z/<~k>*^[j(XQv<w
O[FFF`HNk>1TDxnXsD6L[hSW.iv%CE(Cj%``!`cid=<Ef`B1uC}R3@w~aH\IfC`,afZ3#3/2DJ-[to^
D1EB@>"GNl1e7v>PA_f<c9&[raL9z7w;K#$LN[7,ljEpPD1kwB:Q.L xG~cng;>\N;c'2xAKg_6AD"q6zN&I3BxD&#)\/Hg,^fG`]`6g'R8#W_QWxFK\r4X@Ju!9XjYp(vB-$=5"4k<$2bz"hx!5@!|^MLcRkW7F<_!a&>V`"9O+E,c&9UDPUR{u	+q$CxOH"MvD+hUY%Scu?<oa8Lzp)+e{}U		>YRj`@5hbhv{@n(M&rJt]bl/vO[}d4	^Z+V	X[y%V[Ucdb%P
Cu~}s~=~r%pOI\5;LJ+3_(Er TYV".s9*3H"nI3k<PTPAejsX;)CZN=o+OT}}tE*qHKuj/{)6u&K9;\OjRVd7s}8J?a[Y?PVBxPglE/UW]m3[#L3omw`~@f-V[1LrXiJ/Pl3bG~bRI?	=(fFVQRqeH2U,(#Vl6(8i:u\}Z%51+1AvNj3vzv\;a*QR0.U>=h5p<JmQ3SgV9O
R'4wPR?h8C, 1+LxmYu\!)RS4E3G6 6qCn$|g@=xX(c8!h$N_dZX>	Y"y_1T|
_WLc9YVLM#{p$v\d@B"z2ohN'O$sT[L/v?`R$s0-kQ3{@pj`QZjHc>-z%ad@`],3MZL>$Bk,(8u?*K&p8*yP^FC75<>}sQd6wo}'YlkEQuNaq|C^-q`D2Fa D]8JD\VTm
O+-vc!pU+a<JX['>:'9!6floK-ea6=4{!@q3@fq^0Zi_.	@o8|njLS)RbU&
cHa{5O@%1xayyN%0&2)~jFn}*Z@$|CFA*j|%nW\+XIV8VnEvOJMvMm-::Y'
8G9E+1T#q5XQ7U'%TLF	H}Z]Iy=(=m	Zdvv[AP, /NaqwYH/?xYts~3-gy{"DNNklp+
*Z>'|^ ?|~_i>^#J9LaLd4K14Q$4{|"OSc;'"^zM`-O!Lce
.Cv7-`Ad5_L"%iKtQj!$o$"aaZ<0f;-rV&]Ro3-JaLt|6"k$Xsm[4v#`fO0w1?d9E!Noil%tW_=OLp*D%> Ed8({sV22^~#k,)p0;sYs{&!]Sfzpd^fUE?TISZ)S/1)N/.gJ]-ONij2i%2K4\a\pO\+x$4&?57o"Hv/|ec2ZOJ"}^VT\L5%U`r?+[svDJ&X2n(h<\Skm^[jd	lA\n{kGMKNUbDhw@8BUz	H:K	|rGT4rl9J=	:(hlF+i_.~p+@`2WqS
#Xuz[fUdRd$EFT$Q0Vwydc8g*Ih7%C'%`\ |jA Mc3md	u!!+O\'27|K5"4i2%c nAmR"FG3*A;)'&OYJw@LBCA:#\>J*qz_}e<ZRU 9YTipEp|5t12v#(d?zO[;EH&wb9$'P&H~
wZnM~0J,L+i-nWnZdzCH'daIA',h2[	>wM'B7Dyv=68bblNo5XoVbqGOrb4pgN"dyAdJO{
3<\EJz\{,pN@x:|pI8v%19vgM@.x=h2wSS3s
IOf+mZh`l+)7nmw8f2R=!sThB=PZlT3>qrQ~y)3C2OL?:alrT>0iE5Y8H_-nt6(}{=#2usD_w`5~V%B)H2- $d"nW:_:6DS fT.5A-"Eay^*tfw*|
xj$#OPdKT[a'2gpn/]Csa&MW5@d"_,{l7*l:.,V{B[\Rytki@:+p$,H%%4RJs.y:]dI,xWJa,q!c&%'6`>^ipB,|6	(+\+=aszuX4?
C^F9i3c)z\-,K`xFZ^7zz+5.Vgo(g]nb]FQnQ=kI$KL.Uofh"PpJBbg0
./C..{@.7@;&3wUVsn9o.`mTPI<J3FPA2f'J`9AJq]AHHEXA<vP<!C
.Tt&SloU.b(01yJdAa\.Y,bjN)M.%W7C
M0ZZ]x91y[]`\z)i5q8"w3#0l&2z?8[C^}_[ULZEd(feRz
?g#g0?i+9"G%\M\N$OO{GQ<N_<RH#l0:8gek9&6;Y/*n{\+zN_23u/UdN_OfzQ?FmCs>,Uc|W<KpJ6tNfHd1(&2)o#@~\P5v2duv,yi26~p	5KS
g}u \d!x+$1@WG~YLjL"
j gCy@{ncQhxpn+dK@]iG$h<q{<*Bjn/1R/M|W:e2oe &Zvz('lgCd[X#NH6G?#xo8p|-i+V&t|j!JE8A4pWx/|zQ xr~.\";oMQeb)\nQZm CS$Mv3AEayzo(Ve0;H/d%(*4'L&=?A%z#VAmg)Jw#zVLc!?l"|xIyLm|k\c8)~h^20I!Gtr&ba[B)(d'eiw~uFq:^}YPbZ	TTDbBXmH3W}iDRKWtFMbFO 0vS(Q^BSf	ZTu[;0Gg`aRZ@4I^ntRa".smR?.VRl6:]R~d)O(0|)yLJIF#]Tk6\:O\-s{QYg%>O!)}pEf,4~:',v=l3@the=f}:7V05k4&Xb|}iwMyM`K*.&fAX'"Venf:ak1"FbOZ>JY=|xMYmwg7u	,.2|NXq,`Zt	/>$pg(jd`qVlYda&RYkQUkU)GM;_bLjR/WxELF,5g<2pSL((2(rZX0lRKSe~<^%sUi{'>	 Y;[cON:hY"Mm6Xn4e~_($1LGM21w]ff-Q3(3_Z3[ux9!?)A]rk&-8<g5LP$b,eQZKZ[@FHF*5,{QM*-C(veaLsc	`I.+%XIiNN t{}.p^5:B+#lED$1,"[);AB/eU]SqW9fcskP)-6+.k5[KRm()nM;$mI:vhKQH2VyI@FU}=1'>n?qC~?-C_)u!?Kpci/@u5-67N^,q.]PyB\iWKT~=9q&;}GJ"C(w(:t(V!vf^| {@k?,3-DK)mP'6&%ha7CwGo1ZW4"7r/lND!St6dU`am90i&j,H:gmX6^?F/6CH4\;9b$mCvuvg1u(H!q/[:Z*eQo	q]9@@S9Y!ei`Xr75WW5VI'~q'U$V,`Y~Uj9$MI>PG G73><=;u|!<\;kr[|V{Q"	+Cn
"T%FRFr.%iGy{
zB>2^dkl&&_:[zc[N$_k	-kMa$dRwNKwC<m}0#UEaQU^n~k[Yba?cvxtfGYCkykUSreS',DAMY<zg&_.cT"qo |k*0yz-bYZ4p=9JEr)nAL0nMl*ey_J:32
_+uJ<L#I:wg-!KJk<>IdfQ`>%*}=@J@{&75xH(WWS3Y#g_EB';OJIG*ic[
F[i{S'BVSPxg&]SrI]^1P5qt|VO08	5FN$XMgNU@t`{Lfd5&8&
m
:2V1v{UqS'c*~LzFwhV	?Op9+xFM8gVOVF?4
JM`?h1"RW3*V\oN%:|\H9i~x)-mvlaxiAl;Jdtl3%&j12DN$lRt`LvQswi|hs+Dmb2h2fT2*(Z"^{L%yk^PNT}psFA<3!bV(.`N(nr2#$1)%KRTphSEr/YF)Mpx&Z#mj(](^06&nk?eG<qT|ZfPR"(/BP$MAc]?>?}1/[{->X7> ~9xvk9'.oJfyIQc93pe(Tn/#@|RYx:Szs^yBdq3HR_V
!zzUIc48_:>|-jw<JP3z->}%vjB
t\TtB4)wx[:@co5d+53SX`b.p}Lw [^g>c^rF+^}hpu`{s.aC|Q{{A1`_ G3Jm1tG,ONeU**Z(JHEqU~0	qP,G3\sd\"nruO:P7yl`$mphhu~_~C5=X}>[i7uh`A3LX_}F68q_/$znQH*RMH2d.)uv*|5~_^n )+:~&E-<S:im?CDM"9':+6
FYXF(xJ^/mvgn35G>5MQ"
[MJ1K(}pBvnJb1,:=B_OJgc4}wh.\3&EE/A2Ede>t`bMoI%}(w}UTD ?Q&Q|]6<JUnAUT}8P"Z6%1Yz=*akgjfU?$*,[UB6spy69,yh3Gz }sP8 T[CdxDK&TV%=YGloLvt
4<iv8nFSPj1LxP,alb8@]l+G:o+:3'6	wV4@cGpbi0cp_E!;uPCp`}f[]y&UhF7koZV9A;H7VJL)w_@
sj.kv};Z?pcFG}08$9)^,;zU>0[X6b]TT/|']Hp.1}6[	!)8Vz=,7xY#HanVNE'^$ 0$,EJaq=

&x:e %82{4uJgQ%?iI5FJ*3GBa;; Uq}C?.wCX,A%`
/,qb0|UmJY0]"aaR1E]IwG	uO%nHu5r5!DN+P-r4#WnUP<eaL>TzMCU.MUeQ<O@s}#)0._1Y&muhqU/jISJvBQ^P=n_]&)!Tyz|IA.\mEFuxK,b,*c:*YE-v+;C4J_g0x7f"&L	'j;_HLev%)[93m!>/C|vDsh,RoJ17b3Op/x%}M^Mo3n^X_qK/oxZ9<Z-5wbj},Y3|3nf'T{tiy^Sw	VUzOf8#1A1Q5UZPUQ=Fuaf.*]Wp(OeyeMslV6Zg+R&'%o0,@-(Bm/lE gNkM	-Eb4eFBh?D7$4Q*c;b]\9uv97t <GM^Z4$T1%Z&^9hAmikq`<?hL@qvKvIMS,WphG6<+2{I~Ey$sUwbzDz~zs&3FKyxB-Ft"*945
FYfMBOB7MmwPje?L{(=A|lW"WteAKS8kQlGS=\IOK1oGJ
nb^Sx~m<V>Kfq+gDp>cn@rS=pUcwL]N<u}ce^[SgXj$
L08.{-Iu})Y],	G|S$SH](ftcAM3aoF)<O(}Bmd=,S[<c#'U	!v{;B@NzN &MsJL6|oht"?7@(l;{i7'i#m&FPG"#DN.8r6B
nwTM([tG*b|9<zU98cta1FMtr)Yr6?!8e<*rQI4aSO5~hM-;m:D$F9vK?K^Ai'pc=LoywGQJ\hv;L~!C(ScxX{;&/`@Xhv5dA_Y<!_ps;6s@k5!T0!(5J1zt6Ow!bnhzJ_d+iL?)vKR79%4eZ0z%jfOAcr"/td*:qt0
D}d1\]Tbf782<1/V23BOAP0a."[,{'-7ah|IXR(3a];NSx>bnAr[$1mu
*R">]*ekfP9uwW@-)qj} w>gaYPL1oDmY:0s^;>-@jA:Q	PG^5xipxu/n*'8!/TeFKXY5U6{}$b=Wn8ZDBV,~!^'UgEb`J{g3W#<7{#v^DV7!S.\%c^ULot.=%_ZHBvRV;`0o=e9Agj,(L)fB%<Zeq!hMHF\5XS!;D2E-fdEL7s?3u3KSVT3>aD)!@L	>MZTkk$mS r'*LXIoB~j[F5fS%'^!=kFBzt+&9w&By%2e+8t1fiiuzXx9_cx?GwES6=(l=o:PmQ.gID1AQ'FkxV-Q1)OmGZDL|'PS@32:Mz9+9HfZ.NN.( )r(Ur!v>qQgUWKD_:5|@ipFC7&gQn8fD=`w8{jErVDn)ep]'`v.Nh	>qSK~ctJLhiT6toyi.k1{FRh4m6uV6$@rw8,a`.^6DgWx"2bdJA]0L%0TKtGJzVyxc5PT%T6Qp~_Y?n~hG*I_7$Y0")Zg3dj1'pAL1>[paG(o[:eAo|:F]|;2R>|zB89)6oG_Ww&j"TGNt|} Ean)e_{@zIuG;K;0R0(mK3lhpFxTG=})Sy7
F	<!JIq3gPu36
{GAL\Dmx1;}KfHy3Rsk
'=l8k=_/	?hmv.ks)Ub%:*b+?}ngy;SCU?7kMP$:9z,AlITo%=MOb$VrZ
%b5#YX|EZK$JeH[|VdeG\Q'5cwSgTef.OuZ:TO^$i4W@1u`86g/gW(Itb2{qkTS0"1RI9,x^IEr2_BW:<oP_S,D1	2l{+p(O9ZTs&:+L>LX&	#iL6W(T2AZtGG=;T`co1unqqU}!0M~#%n0e\HZ5:!*\$qb*e3/lyv>Z\Sw.u#<UpG-jsckxY"hWm$:4wb7@w45e9?^`9lgajX!)h&Go_&U-W42oXH
%x	2n/'qp]+yuHTfpGxk$M\RX@wrLE^hP1un=*Z3&t^G@):to
2
.<|Mc*<Xe+pd1kS
,Czu;0d]cZpz9oo#M0Yf]bus0+	;iP7[FyS>rews),(%UDUb[?,OQX+zc`z~0I."m=vGU1uhj">23\uM2,'E_t(
q7( dS9O0U$F&v=	sPJ|#*AP?-Z!
JkR1ltA:`TKJx${U]s7.x:N5~\gH
wdSin?*Y]NyE?m@Ypaa.Gs(|hIIlg	"$,OLh^#+OX.@G[K'+kSfRp-wUKE")g$.pIW	nx-7yAZgG7OkY5LP'*"Qk`4#chY'`]KCp=gLZ8n5NyxOB)MV#:do?6cp^7[Dz;s[l5Qj)XrE\)|EDm1X!cAOCL.%jz.:k.m*Vz`/$,_iXm]S3DK:g.(8nAyFe\7g^^8b G#cc|s'`iyv^\n(hG0/[{Io9 =H%IVf9`0-{P6VdR^`0eo{l^j*}^&'iFor;K\`O,bd#e-}.Eha=861kPYwZ^_pLAvn7zi@+xN!hYGE	B\T	)T]/%<fz*SJ,"C72VXeK3IqbY5jhB4S*,hHsXy.4#idx14/&2Bmij/Wd;#:M
7pcWTTzq*a9q774r@zfC,|++E}-vd04bulbkxh)A)xj><9~jyq1zjuY&1!~:-\;a8is,D+"c:Xt9rGN g8U
hdr:NfY29[PE+gY1MZ{ZGxR_s''JU91rphiB'"sv-hOZpHbcJyw|x0}<q[-wD<Y z .y~{d$||g5k@"2HYD]|CJ7tlQ5!+:{Ch#	u/"U5r\@5l^:UG^
cTRabUf1-_4S),;}}dmf31/42;q!ZcJ[>EF8`$.]+BLa-5ih~OU;zh jx2%<m->=:V8@yNc2~r;he`91%Lr[}w`'>Bn6N\;	WrNy!^ClAD,2#+=m~I5'` FAdBEK%*a^~EKNG,H;fsa3SX|YLp	';W0&j,V!?GYI@&r|sbp3DNT #~Yg3f^nm"/L?4c 1'oq}:haVWg}*65?byj$%}]pM8i|)\x\B]47^6_#=%="P$F}_[0>jLDsr23x5$x.~yxPF0vSjKM)FE|>H]3fZ/?v*oEe{Z'N9=DfOcgd,yzQr*#URi5i+)6+wB*m-V%eeyl6H+6g`w+A7dkMZk04s{o2.E|Ue:pVHzVp(czk:q=-"hu}Q4Y+?1Z!U$+.0v@.B
e[fIa0WQeqeck,#3T5i&o@8yNwV,i2\=iQQeBw`r5@[uwy}d`zLQG2Sq$0a EAG\nK^E),;5\FqW_ye#Q,:t0q?QGQFVJ%6\U], k^!Gip-Sn_FL =#(a7b\o\xW[q@!Kw^b&Ty$Z{{+Btciwl6+hZ6MTzcb_H!jMPfk	Sjt!Hy}2&|&b
k_^A@TP}8xg|TdjK2ksN-pfU1mUzy%i
P6\m?sz2Bo9ng
6dxA|~X)e^f\nCb$54FiratXu}M,TCrC3 {'ooM
,x?j1}Dtj58fh+	V*}xx;LuZNP|?,ketk/q6cmLZL)b EH&v&McGYW9?l#bE&sr3AS{Kx?L@qAZ,'3RiIK0+3gBG|'_wI@wono.zNN	X]S&6~~3,/6RDZ*C}A;^Bj-zX-Lil6k?Y<!#8C*zU.-n~PK`3,,Qg/6'~'`}pmj1mZ	\pD:a@U6{Gl|gx7O.2]Ta]d:)MG^'aE6IDYz%9 7#|zqvFgz!wv/SE@}W
6M7z,mZWDh<)TNKW(_?T#KY|PQ-b8}vHn@$[zco4;=wJ.H]Z5}iOg*Tr?I
,2KHF<u#F`;;]4Rb"L$G%>Jpd_^*Pw>^A(vh=Ku:%c2:*jGSFFDtfyp7$~-*v0LtmoO)k\`/$185grP6;O~uh?rf>izL[) b\eF1{fGf(Ku%'PV1 Flv3=cBb"	L8]Zj=)YIq:	KJqM7kfc/`^k|5.H_M}J#v!D(?&9+E?{q[!gf$vx%B*+j42+6h.Av*s~)[(faf\NS<6(9:%+5Jiy>"-|*='aHzxtwImYzDS?}_U7B?aJ_NWlo&v]Yx)n>`UX46RZf3n'+XFx<oOhN")&J	Z{lCJ:'FVB:$MBooJDN]=J$|@>nLHvtxc{>V=>bz<}1^Rsf9BQ=;f$ uIwWrII~5m~5=^8WQht4l}i.LiB_ot_n,S[wE	="	8@%.4T=cJg"!HT$zCx*ppDbNzPjz("DYK#GE9WAR%kW-)q3^ySo_HT1Q-Ym`e.?xR]b,I"?{"J5ahHA(d
#sj^u+C-AM7OW0n\tPg),)m7?p-ibhdeW;l#Pf-@_HoU=.%TUy1C=}!amPJ5DX,1xzJ3Mf#0%g^WjI=?DlmDo(M=k| 97$qylII)YOt"q)8b1mTj/6Uz|&)=mBq$y>DuT#y9Qn/1^q'-fe$%C#$'1-[{FY3f#ROQ$O17\^W}N`W8_PZ[0s_RaixA45|Y	U"dzC4)xT01mSwu#JK-UXr}w5g3&pv}
bY1v4 6;neVEukg4X:<^GdjH]efgk}LHhOx[:ttF/R	s_b>LLw8lvgb [.jW\qSiU$jc2(s |L?`Zy@KK?
1f7'7Z5Uo=5n8%|,a>7,b6U['7?K"&R"(4$5Bzqh=ne5tC7(!yiE.(@wt`eArI|/<:&K?p8}pNrf_e|&l>Mw@!If*lhU<rws/%0s?zU%B7s@:c9LRI]uy|3EhU2"/ULGSz.axMUN.Jy|*-I(c**fa*xCe DLTmEm*>)
a6;fC*GtOa! Q4qF_-MQ[dymRxv60p=dW`b%:uceV~C1ayirh^"i9tr=(zy^vZ=]eai=Q0G+gp9HryaDgQ$~toEcIom[R.Xz\Z>+?x![%6JdQrPi-f"z~ERm0Ln(z+3*"H4
6`-@H|Nxnhf+7I\U/aigU{jTMhX8(GJ{C0{l8YT		+Z]<%<x@x@bUF3z,#0>{C^tMWQ
&/8HXj!peMWTo)(rg'[(I$NYe78x:.@A(BC)RbYIZ6O4Y_<3"Sh:t(sL1'31yG<r;BV#E:P(b{4	$DH
Tp83RY^>Dt~2>(cPN4A3,=0	vh(D"]>F48+jj6S!&%Q@\n3dsqor+K.`)smQX)t+),WW:bF]h0ia&B] p9[07+HYV):4Nhh,6x|M5fmIY2m;A7+EEXZ^=Lp:>j{-0QN(z%u-_hfZWMX_tJ}bpdv^$ro3=e.IU@iiNhz-OrMtjV7t(4j"L\	^x,gfC}UM7DOiJ2]Cl}s:G@r-"XfYMK.38vqTvEj!1(lx{-KoYn yI^zI*
E:Xbi	=Q'B$jpw|2_O02X31:!BVAC`f&P	 ev]`4]8bY1NVyNqy/&}v`Kx<8#PU\z.*v;yV2#P@32dOLd?hJo-TA<FOfP\KBmLKn}u0lk$ZwtZ@D:KH^.3p/}CMRgTvh5&AnTS#9">)']!OPX`%'\pRZyO+RT]x8.e*]e[(\e;<Q@e`0qKXsiQ>4DVYPrNc]'_`NdU6:G<2cXB]sWt6v'e3e&w(Lxu7vd5*|MU]9KtHe!ejikAG=N?BYs
H[\SbD+_qMktACs3RK@NBlauE.fc?id_Fd1Wo.BKs
I}[w C38\"6!:dIk2J	OK~V3D&D20\6-h#UY
)xwD4hME.sW#=d/81Dmgx?ZS{hp]Y]Mc$:L/MZ$#,~z`cZGu)'\BTcJ(8<EsY!H878(@hPO*h;EV[f&4>Lkzaw_cGMvn#*{iE-abR}MKy<sQ7+AhRQJ5~2AL/$>4;CdLd[iFX,SQ^9#$sRbwvIA|} o7(x	L#|UJa@nY!5eYD<Zj.n;^)6+l6,!dq&%?_ma|
7IF,Onu?x "`;
>dj_ar.iBW`#)IcD5?7@*6NxBy]xLIw$8|}Dd/\p)/rm0KT{)}bY?7m32vQjWZPD+6sFJxfzG%*&/0pG&dAjqU8I+<&m/.3X|*n(nzSI?C9|L>o0}P|8)c;Zo^!A.{#IKkOrVB;6;piZ3B}<8l].n_#BJ{DWFd0%hR-$q 2\o%Qcq&n}L+2_*i#&!wEVrU8U!?wGx[|KEiUB?MeeT$ G6zdVUWEMq0?'9v@?.37qOx2gn>:4HLwxS{f$O:%D_d{)KEe&V2;lB1IcZ8D"u#fg	&=)v4)"OfH=3e58jpwu<+F1K&P]>%o,Z=?\Tf|H8i,uUvP)0Dy8F\u"wd/A9H"y0'}>.%Q/"G!xACz|>7Q({h1oPLml,F@y.AC\@>90(-J7z?]_C6[m\r#	PiN\YA"^q0"#b%~05?|'&"]G}]BL|M4[q%I|2XS<f}AEM:N:#uTZ3".Kl/Kya04O{b8Mgn#yCT*)kn}#RP	.%X"OXl#|QmJ2*{d$$mPrg=Nb_KT{ !!FED1:z,5/ATcbn/G"|,jmfLxI70ct8Wbrp<c"o'pmkrM3F")]?R@UN-@`Q-(6<'te/;/1LH#mx'E^WIRVrnm.9rTXoZ]`wy
Sa9?uo
n-wFYUPoB_"FhmpHjR[KKs_~uwf_57dK!J|{rD
v-:2fOA/|x4CxfA<+@Gbb6+WADWSz_W=FV
T`'F.$F,6KwFn/nIxSm!fk1GFN/Z!R?2mfRj1OgP^uwf]5Yho80a%*h3zMcJS<'C=}aFv+=^JrwoR&V	Pw	~A0)`6K-d`cw5`bDVC14l[q![I+=nU[VL;y~$\4Lonp:N'NY	%jtd	\/"smj-e`DIKG|4x+ptw6HyA(7V.TI_URdZ~C6(lec]!E$fB*{L]?EI(8ksQql!;PmU)et\[8oLIr"4I4sHT+r0pK.'jhpmhU\#jN3'IDV?VsqtJIpL9m<dJFaS	z	[Ks1I@+.BL}p1i@"='hPa)BE;`,Q7*tgz%aIc6zait hySmC%vM98hmXI7_w#BZAI87f&u1@6U& zU!B>#p^v$ne~:]=+`zyC/?o
(odEK)1/Au) sF:|<9/,{T%8[XYn8D0d\*wI1gwqxMB:`q_^6TR\?js"bXWJ
^q:Q=&%@^WsK
Atu8{ss%`B2(i5t}	Ow"u2\C0(w~-Iyhe?>[uSi*Bh*sPkR|Lmp$1D<tID>Jq^hs%`M[S&6^<X:R$(6B1(X6}1<Kfn!(!vaFT7p~$2l[_hGL;a(5MmY!Z_[$$'WR{4Pl/h:	yd2"'bj.c3.OVYqWWXtCoeY7:QwL`dS@Ik|G,_?QffiD!!|[Z9F<U&$1@7V(c<_I\3uW=TVArB|S3!:ul,}tVA7=X}Kk;m/1Ne9"bg"
0H~ttmwcJd
{al#YHYfU*vz7@nkY{`VR*f||4zK/='(y,@d;~^7P
I$lWsE-)&n:LCL5-}lT
J zE={D/|j5OQb=owe40>.Wu*vA&5!s%pr )5G^;s{xqC>V\.1d?*s@*3Z4m?6bp UpkKegQOROeGkvl.dd;*gGR/"+EBU4`K#DVs^4FZt>B	9/JjWD@&bmjGQ!6}zVm/5".Cs%YG7BBrId$.>.0n	O9%&tiNDa/\xM}Ymx(>y&FV
=w3]=El QCdlzU_OwP8]\/m.V27~+ ju9>A}o lHB iCg6Wy@jHT%J>BF<D~T`4P'^w}*'8v(!2nsxp(nD}x0tAylTb&HHp_`Sd^`I+hCRCj p(|<	7$w69|
^q?^IzLvJ*!"}H<:Yj1t=,S"JY=p5O$U[OB%PlO;}r@t4yD?s/{KfyMl
Y6Z)^jckXcQXfO8sn5.Jl8	DB~]2]aQ<Uc^SJw\ugoQD@_xxMDX*B+wk\_leMyasxnyYZ7Pf/|,R{WqVzMG0YK2+JmlGo/q"kO3=g{"vSwsEsBq;BuhB75/_&>T~>:*WL/IixHT K*4Y4x`Pn-)NdbM1U D`V{aP5b>zV$#A.qJVa	"p~*a*zBbzH#MCj?]Lhi!Om_721	Kp\EU@u}ql?Je@NK`;`*@O)V{N&)G'A)t{rT6'tgx;?]S,1>:&+KHQ/zU9V'
{`e'D6nxeWG*HKSOCbvM>i9Kgks6-$X<#W7[/x.	%:	5D)Y3yO$i::|e@YU<7jL-@i|BMb, L(S.6)b]N+.\#m~|k)n9CUhOpD&X	^o_R?cuZU|UV>JJ$!=o+2:P0OxS#|`\B!C2iW&!6kxmKhsz7kv;be&;oFPi1>r(Kj40^?)Y@N+	Ie0`x}HdhIbb^Nc#t+6nIo3vj9OYvM+qLJHTKiKfc90q33DjP8u[[\Pt^B$nNf7	/JQvwA"hB5._rKQk+IL9@eKds])MIh<!&fVk~$bWU`|OF>[7'0KQ:P r6!(>o1#"30(.	xsmF"i,24Vz3qze8.~Ds|2qwQ2.UD%|)AzVt}
]/_%v="#r==92RJg[GI}>t\j4d\r>&[)P?y9mEv4Tn
/d]-ip?	Xb;4	um6N9ady2cZONsoz"B6F4M+}M@Aa_i~Z9f/[Y^kWHLV44m^$1Vw6hr]&4U=.=~\unhp]Ei
0]Wg+m	L&|_3q#v
}oJJrhb1[Tx}XYb!obEO+pJiVV{Z62&q,BCBUQrsq	xgVe48[Ot~]F*7nvji[ T%9:3u;-|>?D(z
m?_st6Xf.S7)IgO%;'8-g1y_.[E\-0X$69LNi*.#|[!t/4]WR$pYimKHpNT:zi..zs#*}=/P_c'PTNF>J15[j:)/<A4TnCBe(CZ] fiLg$SJ`)"CT:x3gN=]JJcGKm4j/=0i2\hd@'7A0i4^Z[X8tN9Cg>#AMFRe9~vBG,R|0^IDes
rBhNkg&}.rX:ljH
5@8KR{EDddpT1`rjZ]
r$> M(aP2
&ri&9grn^yQqmNTV_o[VAW\	!b:55Y)G#IEmi8Svx,["xx~j2_A7)uGo+0UJ[AJO)!S>XcJ">STBa6,.)C$*a-:E^3/y>4CHPw\KM5PSk&tj+XD] <82hX%p:GI ]7%lc-FBd6-&zLo\8;@_{aBVw96^NpH}SC#4P`e_N"A#I]^>8;AG4xqPL`=bC\l0__a80!+.'JkeZ5YDahN,JSp.?b}"yOE*h\
P8*2\?@'tX
U@b+)'Rh0o*-q^mEh2m4<q]y3'm'Od_oS-:Sl
5NtJZLt$qf|Wu+''6@^<U3lK{R81F9Sk[UJ;0H_!DvB<IS
IA=jh.!y`F}-`{8v&.@?4n$a/sy^[7nzPGIaJMBh|JP>~'GQF
vgut(,7IxP)*F%W\SPX3NA!69'X6bN9:ra'48w [ymZ`?$S	;\oWk\t"XjF
_ Z7x3{O+Mj.r4"FB*kYkq~5m"\3A?GNhi
R:f`%F7lS3oe>7}]t!.RxuEm7|IYmD`rD]9G'Q`:@:TMDS}=9L=cH/U-w%we2Wh#4x>w7`~*eaAz, :n.{k"x=D.18+-n/kHy,QIPx&O. dNN13{;FS0V";?1DRPjiTFpbT]{"%{UKB)dCGiLxgpN5U7bY67TASpu$)44P:Pg.EJ+gPihKws&;G2CAwX9yq]M~+RtW)I6~)VqmH')lvkIf=VV=$:_XjgBvI<'Q^YS'hVpM>Eh[HNZDJX=E')I4b;Wmeerb{F>Cwc]"8K(ZsPt}XKQ<&+_9j6_nX;N#UYIQujoK@"Pyit.H
[Jw-^PTQT^#jr~"e#1*.8{/Cl[%)AkY9zzTdl;^JDFxHKIuU&aU)LA%8	EMyg"~k`}Vq*^.cqF^@}CQ]s,D6l}*,?mQp{G*rK7E0R$v/l|'!OTpdlj.=]Gsg*md9M\^K~E9 t7FG7[qvm/ZNK.4,e]PJO)jrEwI3vrwuY#	:]Bi@cbf#^Z,Vz*OOhm KFQwA@D4Fx8`Df]$k/V$#o=Mf!\BmmA@TJ9~rs<wyQ$%%l2uT?B"mf mfeZEVUla5z!drmrwXX_	[?If2K:6{i"I]P!m7KG+@mmmE]xxHc3q2m@`ue xYE~`,*in"ya/d!xa#0qn}Pc+IJ?.Rw)(|
;0@AxGOvy~eO1b+8L1!]It?L4M&T^[q2~!,up3o"V-5+R4PO0ftP7BJmCt 2H[I\IeF(?GIdMgDg|^|CZl/4:Zm-
.nT:)8yCZ'YbPczWandF)?lu-.#|Y<7}<`0^Oq|XHzH@.hbNAGn^G)Y2,IL0<"gQI8c^.X]9;ma3S\CDI\/W(s+Z]&#AynwKF|Q	:UV]DPzhi,ix98$l,5>w(Vw;ORQfM|RS|1,deZXV2>k	_0A>:p`}jN4N3MDB7K!)3h[IP[=]]HS]aU	&vhj.ey|`e`Ngy/RgOA2s[[-M/9z;Y)Uk2OQ$FX*IfOor7e"xOPGL5;3cq\YR1-<G;dIZEuo:6]bXT}Q4T
9Vu*:(;Z<zw]$#UHewXwd*oY:vN4'8#{R*mP<@_r'}^e.dfvhkY?h+nMEpZM>nTRhIb\LOEvC6oMZ>uw&Qs/klr>B8CNk>ojEv5	QD\k'7;'05<vqB_9'xtP0>Z758qj$%
U6a3qWz:RD3BIta	XCJwksu) ~&HW5VYkmm`5-Nt8vKhtQXPFAv5i[:	i\jtL]"yV<h5,6]i)bj;-"/B/-hSJCmO#qkZq\>8xNEu_Ks$ n?,43G}QTg)]xfAYd'B_hYeyZv9M[c/ORi&C}6~8Yl.C~<bMoW0H^N))?NWKg-ZYU<NzY^?`@?n'{7,kaub*-OH6[1C DoW<Q`n
bC4seCNb3pG%+('jBnKZT-dPuhQD)t*Nmc%i U9;3!~YE/yus|Ej4|LWgl_]5n{=<4m%q"D0*cK&n>u\$7Iv@OY_3iTvh;}r'[oLbb)_k4dG-H8
+o,L!~R:`jFlQ=]ZMde%}N=)s=owe?YRSmKlrG!BU(fk"eP)o_4:Y72FAg{8a&a};[6NpsDi5qx!G7_qnW07(kaDd.DxrWb+8hopLZ,~:OgQh)6Uh7/hM<-Q{K_5*YB_HO!@UK^q(]G":CaX91"Wy|xDTE24!+"q2c_Yl/15 xdqOXB`>,}vID{zeN2o|I~^Ac0=@
{:UXQHV)AHW*i0w>[!\_3!az+mu$/Y.	geZV5(dh4vC6{R/G1(*Kxk(=h@hE8jh2 PY8q	s Z+%B{^(U^:`d|S[6y-e1
qP! Uw|o=z`mAdS?88Sa`fQ/C
\
CU[C5vL)rLb8R^vC_2E3pJ	NL.:mq$f`?Ds[]KUA'^MJ*eezm_vo2`OVB]&?Yk>JV!#(sR>Lq`SaJzEg|8<3")(Z,#)n{ay^lZ/O+5*nMh%?<OC[1WP!-'!Ug&J	EN8x4~WUas2EUAp0tFuG~} iY0~<I*>5/2iV2U:2ED	R][QKqcd/B%@54}DnZ-MO6*gaB"Gp0NY(#,Vu_I,I(p+,h!=)J5?npFO" &~	1XUPJFFF-[ZOk<:=X{5j!>IXW3]C(\,=s"]N3#owcaw>4QG>-TV_hlkG\1~Nlyrj*id\aHdUn1#E<E~,!`;d	i/M~ztxCBcW/-1@Fjl;jcJw*xy1qKRtm95aJ2X:wCg!;x>ha	`]{_e/w0/{fZ	eRc#XWP*w{{cSJ1XT:'Qpz w(*11qgTP S:U|-Tono:dU	Tbf?32\mg_[X/o~L QC5^fy]1_`xe,W9GvD"@l5?H|t:D=S#hgn#{~*wa dfeAdKRHx	N'sgi`AaTNt>Iw#s?i:b	rBH3FjJ\[}TsV>U'.9mbQXfT<WCf@_Mg@k0".e+ Q/T[9yK8Z$~+>+ ~
t^x&DnJg,R\O%1 )DFafN$Tqasl%ewg2s=FfV~fD$~N?h<{*,W/.XzGy&5D
pBQR_nys/726G;4%h?rp6.6T!e>I6^L!qFKXP1w}.0&WNurkNx3wPrEMgTW[Z;rdtesHM4<jAB$Af{dwLl3}M6)_!9`:@'_qwn<dnT_~EMoUAgGU,`\V!<_Nb&X3HBe']o]![qt}vIlLF{C.Y[%xIyC.M6*a&^'D)W7){seU/CF8@-V*M"Cbf}~"R*O#H;	JaU|CTl{qMUn:d-cJx^{;$q<E5l<^6XDZ\Q~itPH%bdaJEcCcn2/`j*~vhoKTGr`!h&uDCJE3xPm[8JKU*S0Wq 9xw|(ojulA+m_z+Jg\9Xk8_t1TXa8ed4uRD2p<Fnrfvvhac|}tpcXVQzC(l&en`wL@+.;ighOThgA_o:}*<<	NNRNcM'kg vlrN-mXQ(>=)
x\PtY	/C34V4lQ	h8Cl(]$EmYs_HrjP<a`0/efaJtmQ,s 0Sbl-tb	>;X+Jvvwh^w1,Rx.b_.	C"KMy(RQurRxE*_Gf(D0RzZS1t\x
.;(OVqx^f"RgeiwYFe[`/qW0<(A^ECI/Jm_0s8[`D:>UO\POu]&N:#xP\ALB4VG0tKrQ'gF21uTt2EX\<NNPn\W+GehrEWLD_]1z6+tBsuf0h#jh:j&d/[wA	7U+M#Xn^2D~K1O
o'D@$:/;-s:u"zmUbzaUg2O!F*5_E_	Sfma e7z\uYvIOe+5I~Te2%"ied}26q~Tn<&fJ!g#yC]CdP4_-=/cX3lg|
#B i{<|^HWX'[W_flEBTcW<V4Tg>,<VO
	
:XO8zJ!Ad&bUuvnPOzy$+;7Qk{[H2v07{I=}A@p .E*J6DJGn(v^MCA<aBZvfcueN3L\~{vziCoFGI8{$rw5!z#o@h,@T"%z(!RAg`fo@Ishcmg|=wU`/,Iw}D,T/l]$olv|^e_m9Ak06GAiK;_NDqOu_~HRA[gyD2m0`2
{	f}8P5^<`k,
i+u!??:2I}6u@W=Xms~bxsR#QJnwb}@BJ	9W,7\yg~GxvyVB1OKws*b20vJE3%kjk`J[x~ENmFf> \,u@iU6g(ssfyH/c',jn.UE`&1`vbTMHakDAZWnY__+ydsKTfuB*mrb[ 2l5 e[}C}KJCvv\WRWLIa.UT8MT@^Fa*yJ[^/3)hf1	21<2!Zn(myAE():DsDg@E(@Z04#q;A}ytgB&`8>B!:4U\=)e6r;eUh7wcI3:ZRdf_b3Vokai8b{`7NX2|^)`=$WVX4z"q>0?..N5wdjFXuT	H)yYq28?(f"my}]-B^zUnp	!aB<N38is &hUw>kf:'>?\B@,	)#+h(7bHTk@]w8}\&}:4a[}ymz3%T4eP!dehZ!VUIdF	|\^s 5$*k8SmOxxD0-Z^pG=0^sQ;~e8ui4Bvm(O$xm<{i8C6nFD(I&"&MR+AL/9o*	-SDNNu	@b2 payS c(w`Jzt>l$b~MK,$uodK9$Z^-5f0#nF@x;0.{flRWR1|k-|c`p_MY`_xSV$8>O7~MnX G$jl\jIy'l8<9!&Ip<C%'( {~. LR^MnB_Nym3Ac~$}+Owl|yT,vlx&2#"?[ 1d%PSg)Z&V!fneEoQbs7E*>8P!O#B	UI2=$u;z9;%Pw>s1IiX#Cz]Wyyb&J|

Y#Q`xeulw cY&~eT9
c;s(&\i)#4w k=B&w-3@]3:-00:%*3" z${]<,"#P	EtWWU7cJ	F|Hv`*<]gS$\=`06njZ^1J9})<%,;})WfB3i6ps`i~zJhzdcPW7"ul'}|jYiw%EMGaS")vVS9*j*uZMN"Mx5:"}IiHB	(+}k'vl&p'[5vT5(`_|#`&uE:O_"tf8u\YGK:~M"Hm@s!~=7wWQ9ULf9"BYnd	"QXoxD1P	#htZG>N-lZP*GrV3esdd8b$#q]QiE#g+=Mh.'oYr;b#G_G%!H$HRIe#MMtF8Q,|zAsG	[`FFZ9$:XRyg`%:t%1y?SX+[uf~bE/^?.L	j;_";?9m|zzVet~gb~K=mqn;6*0~muVKV8+Z5o	-h&o5{7w5,3td1(J)cf}EZ<jdqo|%WKko"Z]qZ5Vn6VJ>_10ydfC%c{x3a0( NkD]s*j";ivpnSOS?s<!0#6K,#ifCl<jt$/y4z
fE@o$+`#E*D%BxX.rsV6:kmxx{s	uT]G<TQZKL!CWS79v~Y<$0pYBC`).49zG6=2&PdDjPe#=$3cKH \{C1LOb%Gx>-r%"1U. cV#\Zn #A5yKQkH>\*lE[[9dV_tux@0W*j3|l$xYjE+shsBH[jaB!c5Sfrduu79	>tGI }%_.t=U*4Z*J`6>kx)81;xKO/!Lg8<5N=o|YE*V;ldHz%(tL*tng(e)n3,a5jhUR\pFVNz"LB CRRD|}_nI!4]:0{51y9dHV!HTk-`
QIKtvmS@GNT]nStrEBBiaPBW2_+kES~f<&R?$g-_DP5#?!p?KA@U~"P@E?PDGo;"(K#`<[5/C03riPrf	Ku?RG+Y][XSPI!G@zJ	uX94M.;dJ&?v'5WNT't$z}*yb`,NA+|Xr]j%S;o?.Lt;p	pF4v<n#lv'IvBGF8gmtJiN?G^T ")@X(Wnp0Sazi
[Ei0:WxE2wR#kt^kzmsP},qD&Igy{-?dT*FbB_\0B|+X4 e *JA`jaAsTE96o=sGhMy|9|p+81b(_hz}
7Xvx(gPu;gFUcRe?{Mlw{zj+,%2j\]o`>z]P8X?X6vR}mLA]P?z.7'c\Jb9!c	\mm&/udsEzcK6QW%h?pADMyh@(v{jVWX]2|&H8Cp=B_i*pYGMg&`pP>m-wBG,a11cEE*g"E+&9SK_^j{{5xE`??z,jhIc,/GhBBR+jR)!+0:wk7r;k<v3Ng?bzIH\;mfA\0UK_)R[3,A/b*EOQbv(N	z5Q3l_9f&/~E\.zK%q[mCpS9ja]Ov(PJOuS{"
bfV5-\j5MdOU5OUMz=9ysO8QT$*aYHb=S`[HK7C9t#IFyPHhqj3@A_4#,Xf$Feq&4[=C=	&!V$>g	W+N^IljG2c1E
	owqo"ms]z 6-S|SX?~zvd"_JX0Im+r$(dj6Uk2T:6zN'1*p@P</|gR	I-|
*o24@9~ZtN(V7aC7MXTjfd1>mH72=Zxd	{sSc3h< P#p3ve(tOSOZ R$P{hshddqB-4=yLv_= )UZ@bzR7<Gs3F~f$Nw	+(TZO&ema>pJ<`si60(iRu:}	C	\n):sr<S?
l&byIG0	,>*cV7B/r]8ywH:5VVQ3RS/^(K{+h0T)\qe"x}d;c^[{x)2YNX{.'zvy{UM+8Y#1N,4{/P8]t[:h@7kXd}Yp7e>F	RiNCX.0ypcbO1u^6Lh@kUXFqZ{FY}Ymr9=i4lyyD_fw.B3BH40/A/daMI(Bm;(Ns_wc){A<"F{-,]MniXl&r<>~|?*|@WA)~VP}l?b=KH@/2eP]N5(ST;KmYgR"C[?~{KXOyOF`6I3KoQnVInpJ1<
gi^CM})if`,hG7{lL%Mg<CX=OLAD0>p=l2f2bNh\'
z8=s6~kZ_2O(qX	C^dK7u%0"+Qa7[3$>][7XNNv666\4*a[pzXC:8}xamc_MUw=5(R}bB>F4j*	DfkQs$u,7'enB#'8r=p92<%"4l),pc;_Bv ~2d_b?eu1YYm-mk) )Gb~{|&H.>R)F*&O,gcuh#jvq7< 	V1fjXzi.5KoWS^RAV\6aHL87
Jx0@)AcL"O2'*]YdeSl,4K[6_Jl8I`67p03J(BkgJ;f
:.0`8#vM8,`P1qwz{q2x=|wxBH@6#D3`7#I,LnH(kNosgAG_@A{`$>1BD=H?/-4Kh5VLKUh|IL<]x7zc^[@px{/R94vh)>aFgi}I M,eyIcl/e&:KgiPTqHwFyH
F(!r&#Vs+Ex._%hk-t.,Sy]x0\F\=xHl1+B+-%h%so1rI)X*k~ZSq{;%PK+=_'<fl%|MiAA%W?>-+,BgpNF.A1<(@MO\M#MMRE2-v1(V ,J
{xY[RlF,=B*YW<DC
QR1| LeD-z6KixK0HV<)s+NAOFFJ,d0f-TD`v>#P,vqi@+pz`i8ADHx$E$uM:h7&I,H%Oa66-'$C' UAmQ;oHZ\|lyQ{>,Y]H O{}"s*`O*m=pa%_2\E3*Y}8$Q-~P8IcH(<T>*"(5,[*X
*mO>L9;yZwxkZE.l:|M\)
lww|v]
}sSL&L[4ZCA_0\%,8@2b-R=cC?W%|	Ji16KQ'{%(|jK"l:9|^IqB&q
0 [a],Sg[ks2b8e,o&{D:H%,4N9yVS]`TaLa^$V!hW=rjs;^$Po[Ah[r:sSi+$i%OQ(("'mCRe~)jpmqBVF+Q<\5 `5z}Kd@mX@BFeHn(mv	s{e\_WUS%>pwE?XCCd>%]:-hK	G?!@T'VOH&5_T}c[=:+=t)C_2X/w!AX[q
ES^}-O0q\%T7c*/'=<y&SW%^E3tw=U?hx+3;4<u"9}i20^xYk	jF,-c~(c9PKG_!YV')Rns"0sZ{:8J[%.yg)&
]<c@Cs8f1jA=>WVB ZwokhNC+NO9S\&HRFB%k.of1n>i^gz?SEEOj,O*l^'62"C6W0QjpsS+(I2+"e#^IPA'f{pp)ZLeSOj`VPYsU>}z%Pt=7;(8DnxN.rXwiz=LCu%_UoKg(&0O- />{-|xln_j<Uxa[}#'&
{U~"Wnb$<i^`D Tz4<[aheD UT_Nse}B/R :8-]f\Akp0'H>#2r/ov`;rL'-!& {u1 {w,s8hc[77W[WH_{!ig-NI"RFHxP<md[9Dgg}P{U8CM^8l6|\qcs$^oFNFcm%LFT$;<#han	KVF9r9am6m/{UTop2xe1.Kz5#CB%\
/@ha
3W3VM{2WTWi>`#}gr^:q;T'9]AS&[Tp(;VdC@/G#lbZ[P(c%A9a?u:e]ZlQI'6JUK\a>btwL[L%3r-vE}P]l].;0h<imDcx-m@_[{.fCFAsHf6ALd>V(to;O.$$(tu"#{bDIw6A NA4-<m"k=;2(BQ)M.=5YzJklU>C Q810C4b9!%4I
$v?5gAMr#_o_jv4ekif^YN>1=wfn}>}?E/hRcG4`1g+%@yTX8'O0L.SMW&cTe8~b.: 3-vR&JW^RB) +fO*/\:/U~_a=Qfg_N|te"J6?:Hz9TccbY\%'w9pbNiO'p*lA[F#`JW%znU5c-v`#?[.tsC;$K#c>P-'%<OJ$!9'V;5]j-Vo2y5A/a
UJk'zsYJ7|UF/Bs.tPwEyx9d{rRU<Yi)lm{(-c(+ZXRVCsLtt4\O>|4rKNdqCfqZ{\lv0{j{Zr^Rkt-hz#c
)?E.PAW+1Bn;v4]\"|t7u}vsz[~#nHaxVZ$jSu(1&in!&QQ8zjdNC)f`0*9\,35@*S',nKKEU^w-KYy{9X+Rc9`{lF;cFD!h['=b!@C;Ru]q)+NI5jEA|/+x7D0|KnghX@&ME3XM1u`CRHbT)J'&+/`/qt{=;Z?P}"U.~72*1/cDq|1u7w!(>
.TO8JS'FTy7DI9|"^fHD	*\`z
'/Gm%!Grhv6tll|sP1tp:JLn8tI5;]kY*FrkA4\4l~$DlW|MM"oLtelXu2F,]xQ}!ML;v6}/ZP]S(W&mAsv~Mh?!sjT:gD?}\o-Vo><:}jZq[b-v<vzyPIfU#xA<h+#N0WE5Fx#gO~LirVR|wXpE2mebTCS^1x}vhY4Dj2Te("#Bw>fnH'Ia/8uBiGe"eXP./
hD>hzKE
fhxV0R08yEp~^XuS*9AT:,oDYbh0m&=~QU^_;-chXFTe}
p-k-P4w/|<sN]YS|8jP8*yqj,RyYKb|~/E("vt ^Y\z(B:J;qEE)bP4JwQWUZR7qnHMb%!Z8'0'MB=0daQ\^]aVov8gjg(	i#Hp[+3TBK5+N{8a-p"pfi?ZW?gkvjKqzqx
[>iLU)xEK!%t#n/gZIRp]EGd3+a!M6v(""}$3n4n7#I!tvAp1nP'Vr%B_qQgL,?0xc\gV[D
`I*"4nMIUktg*m(E*dQS7tcv1/uBI=?[*.Vq	_Uy|<\8QbM"+UA0_v'(\RcuE0L<j(u\ <[JgbhB=sQqbBF3LUbXxr!T\L.}X%ZE]&`$2d'IT+4Fk\kmUJ+QR- 6,lER8 
s*PNV:ElIWtlG4AC>X5h{STF#r,7/z"I=
p6SE#.*)(Y#9&Jp>nD7~mf qC's}KNW!NU1hOf{M6xz/2|$2A[=m<5	[hHC4ri1a-s_=F=OjYdC,FdQ]G>~e_{Ry$H1H(EVyEiuGCS^Z3-S_{O0/HsnI%[;,VfNMn-vO1'Wt'OGwLwzdmEGwOljRCq:S\,n[pSXZx_Y*J'H|:g^0[dv7
W_8v 
eEtoCZ\x(};I[]}5Ex9B{oIl>8<o4!qoJm9e+3*D, 9g{o^DhUXRdSaCD'
^/M[%=(.l1(W2)	<}U%wL~/w^W$$c;9VQ2np;w8!QfcF(fX!])-&u:jxb:1G`dfoB'0<4EB`2m:@]*/"!<\1K}Rigx'lnDygqFI	2fj%e1|#uD|NayxcL	{KFbkIn(`saH-m36:bb?4~}/p;0,qT	+Q-$ K+L^jx,/y8FWBXr
#t8->v*A3uco^SmhR,qj*v`,:8k~v4HnnR>,S]cH+W\{^Ua^pGo~-iP~J0i[!1/[h-&Am	ec*$zrYf%w)5gEs
;Ptd{c1h)&h13LjG}h1,l{*BBBuLh4Tt%4w(u(".flZY_X|S	KJ?@K{yHk)2HFudn6zmi d20#X*i))S7y~j:6)$P8alX}GBNpqLF8AG"'u@?{<Z[ug6Pban[c-oir{E23g5_A\P$jyirH)HJwAiZy@8<J@y&hl;g&;	jvIk>P->!MM\(e)4j^X1^[o3SKD_/q
X1) u)<h}'LvOQ\ph,YMjcm!-\;lI8V.Viq%~`@>7y|d	'gWM(6Cto>H/2*DLiO\$,[\[;[S=Fk\H@
<Zkug=**\hasU(Y66f$)Ko432MG
eONd1	tRg.dG$/ 1=TASXn%NKp(-45aj{IdYSv~E5ut|sKj.p8z.>?>_t_fYd%zBW+Om8eFm{KRlB7lZ=l|[<%	K|,*dJ r+HP7-JwlFt4q-v)9hN`$Z";4`*<Wbx^2mAP%2Zv{7A24I
lY-)Ev`a8Ze%hLk/+'YX[ea{?:{W&n]	Fo8rjUt~C|:
iNDOi5w_cxq!MJWT(9Ksk["MaWj"Ujc{zv5h|n{v@HH0M={XGDG6g~C{{F{ZMAE{7uf[@Uro@e1E9kaWVj<5/AUi>=) r*iKb)4:z{X$I[L(V
=Z:"g=#<>Qp%`o^JPilC;l;LH}x/EIwr-]CxaMeT58PTv'EwULlE#[eP&EV}0HQKpH@H/F^]Kb;-e6F}V*	07jMoEBhEkly-DjN@u(#	Vzi4u7'+9"|R|U=vA[-/FsH
\/osn&=FZy7_QrRY^MX`EnTb6pq>Fq`*dfh'B*8}-a',YU~gJ+mMW=B4ny)kloFJ_-dW!"bL>;C!\+C#;/eeSrSwSOYAgI>S!+w"JejP>G1*Q2kH'.gPgdAxtX7t8HN|5xq|EYs9r5,kjp'sC&
Z/egVZ.nA+o*F+dyHp|PQb9.eQB&og)8N?}f<\woD]U&X~70a	TRq=wQ\W#*9xzev{k~r+^/=dj|5s|+|?1@.x!
x[.:ELHo<0_=z#ETGV#+4g`)VgQG?+99u@/Ke78gQ#_Z%uLf"~g:1$dW@:)RE;xL<(2dJ1gR]zGRMBTc;j_&MBsHb?ZJrqj|	Z"%oHR|9	rIAOg`TH{wfIK-0\h"Ufazyr3Xme2*{2wXzv4M'(!gyx'At6AId7cloR\pg{j;WHt894a9=z?W]T*HrTv9r+#dk,	Fz:=t|:^cLLSl7\G-x<O>L5SaU*'JH+
^Zb29hcz7/\<7[Gh8	Gv6'U~=C2KeO(<s9Yc>N#FYOtq@X|<$ne|	oJeb">9,ZpXTaj^[g,c|hw"POyYvuFn{%WOEl3 @R[si_EA;Vrm~@75HI}
hn2hQt{{\5apd'gQPd-@[{&pr}P!B]JaDy%H9i YyLJ~uHOg:Cs4hy{S^@c2uh%YNrC!R*0Z}ep<Ofx`RJ9|Wor[{,1h{b78gJ0VxYPu&b+Su6[5NS5!3u=H9aMR%j#~q?8s#Qs}.sk%CSWd]I]	~^vqo`OCYa$M	",	qR@W|q+A9z[G-)[Vp: 5I&5p>c]Q~>,X+3+0X>uO-mgGn\C,Fj[7U.pP<*P^1'4ZJKSndrqW#Mw-yD~dt<Pj	Z',z@.3nE.K0OuU5Xt@{:phU=C83>A5N}+\pzMI'jdNzE&d3H}*z{vpgx=p95=<>1CO>%fxIav,*2/L6.r}sjX/cI_aJZ;VdQHmD#8A]xk95DPM"J'U6q<`E4&1-w@8gi_?p8#yT|C[?(QA$zBxR= KuFYWg5F-$OU!?X1)DY fq?s`jCMh\s5aO	d\A)rEz)-LPN=QKrn|$V;+2vDV#3P<%	B^O uq!Ln::-~(Wbe
pP>VnU?fw.cfJ)] @?A5yZ(c)v}(ri$AkPrf^'MvSG/p}6^Ugfc%RrVF(WAZJ>j%!y`$zbUx9Gv}j[x1yTS0a|wY}}cy~#O	VJB.dju<q5!I@(UmCY4
U4VOxwV/{"CT/*c#I[!.r#oYki>*NWc97-K>fP6w*xAD7ov0(|@b./u_l
ru6xX[Cwt)Ht=@&
${Ghn4yM9T>Xy4qxRflI9Zq;B|;B*N	9BETkMppW!HU_O"cCL*FGGIsF>j*lfv5U&WhphB.VbbaO0[Ujv;.LkfoS)b6,T TMq,sl.JrfvhACSf,3~v@-8:/co$OG\Gd?lsfm)-oH)P}GI[6xFgX\PQ	GvxG0:RiL#5	0Il$Hq-T{")Qm0E["'i=lBD{Df_Nl%. wpL#<LR ~BPZ2`T1sj*7'q[{,%SF\y#_D\eoy71c42C
Y	l)q'Tt82uJ@EW<mb	seF#u	&ohWDC;|KiH8lkyK'gtz0g~tg
W.W3:MrPV6[qsi3e.B:3<%1"gyx1b$w]VHo]Sx&U:t3$B2f4>l18bj`qnJh&!{u{'#:FCPTQ*V:sxK=bZ`/69nSv;WqLy4^6x=`My-+$(0jRKS~&p"^Bc,mBh]C4b{z<NG+qjxuwoUuh`1
Wz)oK?Nb%i[)Aj%\7aujy4yHqUu /5v2+msqVWBu|>.%u?|U"eB$!QSPaVwaVA=(l*AgH!t5W=WPQ=p2x_kp9;;'|(-Dnz3P}p>TE0V
4e3lL3+9|dw}xb"6g:.XgfV1sBwn>l0tPt{~8Ou45$n<^.SW^[(&j+CgUJM?hP5JsGUI"YAlkAn}eS_/L4vQRfkkzdd/BS@-AYBB8qm36$iFW	=>oOk-zOD.9{,AW!f&WJ~My(x|aSAlQ^(?/$.?46JV|P#9 -|	R64a5uF#*P56)^0g0k.qY2s^s0)`bBrQ#iw=/``XNo"`Dg|O_@o[dMG5:'vGfkb2N04j`k|;MO.' aBp?s2OB=3TR!#JP{@efiBen50eg='h|hR"|]2KxU<F\hxSoLXAaTc7y}P:PnuO,PX::^r=hG(y.1dFh3?D:#"THb$$
q Z*&\X?rd8gsm
ZS>s")G>gxTb'[SQaf4p&/C%A.\:)3I++.d~0RNXD"3I
@3IU oDq\g|y6jxz#U'sRb\nYk5q+'qr+	:@Z0{bAa9@QNEnB#$[.fpM%fbV"C9y:;^S.Zf|>C2<(KfTyq4F1vG|~8!7g./Qt:Vkt.j3^?t9z"@mYZe-M&2F!2_WL9""Wx?Kz kP&d?i#rfhES=CG	cTy=:;nGD5-rT";Fn"vT@8P c@a:!.
(/,1vO%nhL
pA0tX,=BRKgE}n18R'17WE%!lzgl O|]lPJl3'67W2bG7p'kDs\,_J:[
c`gmyLaOEqfH; $p,X'_]S#_ Y)-:3ipI|Ov<!;xx{Sdq;	\ZVF`RNoS	-zaQ/387b9das\f&EyZ(4/n]{iCJ4tnS(&zxAC'L|1nmTsut&o(ek]i1/$h1/CUab>7%xsQ``N@oj$I-4)LUUZqVCuG5n?=c$\XuK@z){XWPZT~Elbj=+40%'XiacM
h..Cf@yvY1]bkr'~}k4*cPTK^1trl`W"Jv
BkZ]J2ed$n
8$;,ruyip:PqyOh?8;3K&V%0I&w[e5|7Ed|Y4TRJ=[l
|f6$1|<Ql*P%LR0c$	FID>t!tClA:%V{zXI!& v
<	!zMrxPrcJD.r+FW2s}@P0w^7.XLmfcFoy>U:Xqx/0eY	}3K"5,Pv@i+SWV^d6i;N8Xp('%m]w|;$9b#]"'o[[R4poQ	6-|dVgP-;?$rqMW[od7}CSA5lYEk]I}tPJ\yF	Ha"!@%Qru	IXDdyGk\b)0SU	2J9i%t'F:cSa:rH23;6@!)+=Bt1OZJeQ(A4<Gu<&:A(dz!=S_VTW@S=4c]Q>krHt:+azSum)6M^0:h|O?Fm<2#&qE(R&1KZ*vhTQ< m57Lm/Kb4 XUdIpq[<d>y'`5me+jB8r\kHb:T}| kYwZ1OvJt,x]0d@FyTsA0o4g$[H=68oG"T`<CTbJ+2s#X.Q)@ef=Qrc?h|GywIaE.zjBLEK=5.'8QNMn0z TO,]x{P!9w$UC\X\n<fId1`lvoF
9FAn[7"m++Kh%%Q	&fsn/g-(OM!)qhA^p49QbHu;(CX#mM+Vp4E4s,&of
)UK)wfx9B>]PvHUcM}b_3Da3"Gb~_fBxH]oLm]S75p2ROuxFKhP+E{#"[q=/F"mQ!9/3vBilK;Q\RRc&fD2y@\x]VI AQN\#\bXbtd=l(p.}'C?: q/!6tRFX&jf<J9rGP
83cv	h+#Y`+"d3"unOKB)~jEGv5,05@RqIWEAN~d,]M.)Tn"f}Y%||:N6>*"EMOh(yY_g	\aIjfKxw>zE\Bm@Nl'LH3,%%W>484tJju@${0W@pacdDD`KcDaT0xJQQJ56H';)%s-YId`DLIW1Hq`4F^tl?ym#0l`iX4&	s021D(Q@%`&fMId#l"7K]_c1HgGoj/n+TT
TW;9\nApZ8d]/A6kaZrxDAJ46QAJZG1&>TN9Y|	
5C1nK"QsR,J4S
%-{_,.%q)=>+;v\jh?)ilo!?n9&({x>)8RUk
]jr)a30b3^xh_e,@(w:okAbW0]	Y0%^PV@GUVB{vu$QEn.j>Mkrg^v:!?.Qqg9iYmN'a%I1$6w{4J>\|*}k_AQL"Wv1SaVMVM<<0`\iLAFsV]3khv_UB!Gr7S|'AiHMr21lD+}{Yp=gZXG[e(*vxdK=#XPv&Kyc(iA7}xyXU#ORRnf;ub~(qI6FZsuDUV=DjFkZGLOWl#1@(8#iu~5d}IPKxDt{Ccg<S3(:>'mx3lq%{>on$+bsNrXBWJaiM;~y&ru1c92*Ggnr,ne`;dz=,\F|=U84*vN^ni6f\f<FABaZ^X#mE|lPj/w}2Jw|{c*,[F	
R)fnwUilfH^:hB[3ai4s'fE4)nhg=jTx"%7^&N};44O'z]\Rbp7V\Th6<t-#!CfY#g_v/+dG%-m@:FZl;^738}Y`*](]
Q4<o*yP/~:tmOSdRvRmX{G NQV]p|.M<)I+W*aE'|t~.-,VTqi^Uh$t >%pEMm7L/5mvW@xlJYK?.,8vaNT.`L$P1~B6\Ld4ok)J*Et5,e|x'F*2	j6TW;IW9OfD;f#}Zj"RDx:*sU)[rNT`zL1.8+	E}@q.),m5>dAh>p-;aQIGC*xQ~W{aV~>wE?0XzgO?goUW>@]\#K6^qb-uNGf^6	!9s.X!1e(1=mv|	'\4UQ\U3m07w,)ew;,c:|
t-^^lUG&v./q6}S}Pm(jitls&>3z
NkC=rjrgS7ybqKEO_J$r_[&(WY"qQ{fPe,^8.@#.6<Swzt#BF]x.[&8DYWg>|7E^>D'5{bCG^Nlxe@S_;SJ6S	_BjNXIQT;lz)s3jp0X'7rQ,49(6;Ms-2SSdK|zH0Hr*kK*lTo;'hJT,&?V4SC)uM|&I?r6nC)rI'2tTJm%#]:}"gASJOk$[z0k5mX{;@Rop0{(lEh
<N!;R2z2V~plVY^<lYRW(vEN1	hX_M!aZhzVgcG(yg'Ay+ADqm77uJmnhP?X\L$Wys{vy<vQ,/=tw<t*@l9-vXJ?g$l;FGxqj4x
&jtD;q'F9![	%4 TmI+bt`G7g2~>W
#== C4H-'i$X\`
ECsJm.@Jy |v`hb]ZC\k`ff|#0cc}"yHb&+MN{2 9B',mXL7jM|W>g|*_kBzJdt@}>>pZP0~6OLNXCMFPuai)peq]>b/RwD(1O;\wJ%Y]8)1gJq[t]!AeUobh^(Y,ex,.$N5e*+c;I4;3"[8%}ZZnyk]?kZAb"T0b0xLV{4mfe5^<ScQ !t&f2l	d	$l;.{Tn}|gY#gn&#_QZ(`FdNv&j6m3i>-inNC	t	m0H>C!AXIf3dh1.Z;QzhY$':U'N]Xck?BFF6R\vhFmun/o--ywM@x#i"@G|RKOIw-c;'DpGjJ9-`K9y2`4Xw)-=p'U2.~
UCmUCx!Eb`d4$1!ZvhJ/N2Tl&3#'N^NJsj>mfS(\j%J&9.RTrGDATS'lr82D0_1IP	&u8tc`#$tY>s^~4i%6nW0\B/r4s[k3t(CrO"Gw$&dd}we|Cz9Bz7+aJDic{=f2>Nvw\
)hHJ,kQS,$r{Ts1XtcGUX"!;*H699gH'W$8'qM<1/biMF@~7l]6A.,x<3K,FE*.'NG!eFP}*m{q`FZ9vpO>,HCf')9_V3[k`JbZJ$I3C4Nspi+QZyUQgR1*	(RM|Le~gwF(qf*{V\C#I'|q%9,m"1B)WBI~}8-kfC>|5k;I#K3J8A}e/ `ZH4`u/).%"UVJ~KbPpXv&]#^g@<:qCA{2@3_x[$>3+'a^sn-V@T'>mZ6KA}6-``hO%Sr{dTtWHqRalw$~_6}N"x	c[+OxpD~.zf]~iFtu&?llyT+U7F*>7Fin'Ouk5r#zin0\ea^M4,; q.#Uw>u<h` bY_!!/2ZvsPUQ{$Uib+(5*5E9Hb0OJ=4WsN _q5C$B:dKFf+g$dp,hW(H?$8; Cf3nl-a@U{VUn:e-u'dpG+@a;94*Y
Tk#\E:(/f#>wK1rhQV7kaum
3gh0QAPR?>,E
tM}hM:TG`!f(Rl8:^#g=Ex\Ux'mo3VQVB^"",c1}	Y[M*;C	JMdX#R7%Ne8d.@o22!N=z)-\o1o0"|r2X\}!zwx= ! ja.CKz+*,6r,Mp&&es11dET%?G0m/1PE2j[E`GCrd%xdo)I2	_98D2~}!I`4iiVn8TH<=$gMGy#0LwvR}pI"U44.s{Q3A|t./}*?YvAlgF/ya]91KxZk.lPRe,TU C$.xzWqow?
t9DB7*R5dz5&KC6":lU(mrY	JVx%B7f1a	\WK}5dMLWlAY[J\g0K;V::D#3^5@q7}6 U]shtV36W2Bb0+=8%A'IWr+)[!zYMjFFjd~/n$]Byzy/H2d%nHl;,<}DL2T6bKlPE0K5rZm.j),4JuO`IruZ8\;Y->\Q{'PwT^"iYt.@
	EzbL&px;+6?p!~	hs]`Vr#gNRPEdA{EG0R^6T0zn;/mX09w	*q"7
?E>!6O;nX79sVP?g-JX()n3+i`iWs]v}k6c[;iWsS=E.sb/Y;`>"b D'"M{"0.x&1SD5Ju?UL.
:S>~87peGjZgTlVwq2X/t4&^dgppe=y+cJTo&Un@^hC4q|/0{O}q=Brvh;V%4J1)&eKD%u*jPNK'tZ`JU^,OIs3Y$4z5VL9p^EZTZLj	mN;F$DsK2(=x+!{(-o~sToWy|B-7MoDafup"bim$6qG;	t-O	J5w5h`1]G&#{KN&C)0?DhUDRM-Jy
fXuug8B1/<YN%UN_V0I8 nkKnF]\0>\o_dHeLn6nz2zsGLV6k)# psU6z;<x\V"Q0\!W6S6?5h]0c*^~Hfk	gyu#Vb%e\M~62	s:y"hYlE(Dxh83:6y>cL*#aS5XLw8_2^1(OPIi=iz:V,M{)W"<Ih']V#gpAbA2	](/[Qcn_zEC	GB).J$j6cgdrHNr{,EpNX#-K yi@\h,<%O Q!,mu@<x:_WR[S1q^Tn0%]Bo|qj+2\;6F%fjSwj	^MN3v;H{>AEC(av	CI&wCN\L(pE*j(.CTd_.P22IEB+p^#w[ETj{`I"bR2C\IID*9)b9/-t@dWgwOZvmVkk^C<Vfa-yAo,gy..Q\Sf*367ekl?NDPo	p6*0r&RIT#kFWmg{=g.oRqdv%0q#k?"Zxr7P\&0!Xn|AdRnqq=1{=Gg5HSHNL}"0dF{C~}$jiv-.RM]J#_VffG-XBk(r4Gd.Oe8"|MQq$!nDvm]Qq~q^Mbp@R|LMh(RgmPO&k=dPIJ$;an\1lzDcvHoGPm@7sG/37`cK@MQ|WGyl\t@0z=rm=hRLV]S9({>cKM+N98LR$wjlnkoGoM#`bgqI#0{Y\u3tf@HkQR"k2Tbv{1&0\]53SmSC1Fe"+*%9(c?#fV}%qb ^e|`?=0w$0dY~F35jvkH_OM$aKG$mnA?6t	P&^|U(VlFI:E'p74}HwJb	wI;&3!&^\Dyb~/]uFDpljr<)	s1[2m&SJ2.Tf|PL-d$Y%q_^{,X8D\VSYX|~z9_s+&`O91:R8>*	-fc!f,5X*!H*#x\	gdJ#FivJp	aE.@?G$.@;&Nag+xo4vQ$C~\V]0t<7_5!g!bn+HV=N538q@;IRXW$t-9[~#FkSJ&7v.7~T'hANKE?%  H)E,J}M7OJbtF)~u)'fN+B&_SxK Z*RG/wB!O)Q%bz,ntJVljzXN	p^u5&8lx44x'N0F\'M~ddJ,),`{KB ;t|_6w.rw)!TzjRn :p7s'&6e2ckF8+)A]RdkQB{dN23u6Ytx5bb;U"V~Z1V65MZgV!|$1{''Ns5}|r_`#~=/a_pG(A}t.e#5'OmkiuV`oHtv;vqbe71_D6P8ICurmUb<>nDD
.u.H:EB3F]O!,
ZH9zgM/1i3&&^n9~M*vHl`"Vo+v~A38(Z1qMM*g2N(fc9_}x&z}bLg2]hedo@Xu\)	rW~${5mk.;e`Md>}	\ThW0bWqk+&FWpdWN_XXccQ2h.{'2fMqY#P=UE
kYo!NQzoLSe0w?b\It4f?17/iRBPf7d5qTYFR6H<{c{	!%j.G5rFA<%j4Z<>Lx>2-?m+GMJ|F==8:ua2YOLD-iROcj?E#*dyh,d:4|f!`9/x*Q+>=c36R0\(UC.(=E+~xnKf(uy]ZIk<Db1Da#<2RaWc*}1u	3^j\BjT|[
p;GXL=?2OX9w`b!PIw9C7SSE8V~{M~?abLq0U^`e}_w7~L%AXGAYKxC-*`ot/0UEB.6i-C\t:{m+oa>'Q3"SG7e;`6[U|ZO*c*+1gR8R;7Kk|?
=',	nu$} 8!8|XwH/9z~>$/bGt,1Zpm}`	7oMwzo-dX(Fzy+*[;!</BiJ8	Q=:	O))n7`B.yyn48B9Z~qA	:<r=/z!M8Z6s% 6dz>	\m!'pO76cG__zE/O&fHB7'w'@<rBGuI<RUu(0z-pl<@4oaoe&UCX[953k	9&BCRY	9zCqL]=3}F|";+%T/@fHr#)r?;B&y5O9zy~eM|q	&|^"u;{f6:uG>3H}
_e';{]}
j#z<hgs1[oGzoAr\GXN>`[:"TpPO^z9boPn:M(d[ApU`#K=}
:Pu2 x$o[_LPk#ps]Wo[aaT"9PDqQ]v8I+~i$cums@"L !)vOW2726eV<Rs1kK=&lQD,g8}vqNE!5eEwg+Sq-TFf!wwN%AU3We0dl@^Z()}y!%1ac9r_m}0V1
d[qls*y-o9`B	+rnXO8CO~qNf6:zxW!WY<fd	=g|x[79?NdL'YUDT}v$W_AQ*40w;^n?MIwV/s[H Lrpw\td]QnaS -5;$o5
Al.:p^HE{7KUg|TBX0{2Tb|qU*cX-:k[5C}f{qu0)#sLU.Ljc2P6]8>l)
zz'{cidu" .xn2,Qq1X[+DtO jL7zO-@-AZub=3nhH @TQ6DGJ[#YpCsK%{edga-1yc[t,npeD?A%^X-sDp0h37&HR[x{zc{7f#e`(qAhy~5jLJiE'2b`H:,-txYv$(RRY8hA/!7{~F]Z$mzvLidj5{>7n=HDEbaC D#1,%-t#;/l[T`Ey_74CUhv35;l9FOs+1dW='O.HS<%U]u~3q6l'|5F&.^xY:~D{y;78
sF(8w(r?kord4t/zu6!jlE{@SP`n!t+)jF	l_U}Bgfo}L{:pPS*Sv	G71QH?AB+^}LS3# /Nsd\5~(2ga3D3s]kmBhWmu`2'anK76bVV\aj0!ojD;	J(22sos"2lP0G'Zm<? ca
q	m\%XqG-dQTnQ=^%){NgOJZ+-+gVvI{+?3p>U9N|uZjekCt]m<i=v2{E-H?c:K!r''FD;@;%%ZA)Q"eau_C(d%=m5FhV|HWunOqZJj6zl D.&4A1nXAcK::rx)Ngo?wxNi82gO|\GGF|RuRP0f#:CMd5_$K|yMQkEAAOqybau|:IYZsy|-fUn(Zo\Y1v2M:I./hPG*UV2d&;&Rqd134dKyOn)[b$|eOw-u+Ra.HmTNHB4)^;DbjKGa6)sjM@i7#j ?]i'zI#0({@"/$.':M;`QNn>jHE|p)F#_Oms!7Gw&]=o.<iMvBwiWo(S~OZ3}!4@}KY@tHyA wht|Bp_wn.H^}1xdj=ReDb4<
\wv%%#ghse4Z?L,hIF?T/9UVx]#*<<@xR=WApb|x^W6&X,b{GTR%m >pA!NuMVxl)M*Lvw_!mA"{j{Me!l$,OG_BNuSrw+{2m{O:w\Owtz=_[$g\;aa4TV230r|EA[P _/'2T<6)V~e*=1Ay7p#g%V`g$xzv?_L&7=/\$-Zlfxo	u*n7Ub_{u,874r{R[S'V,0Gz}8dVJh.!{	tZ[HOTmS\e5%Hb@1Sd[u$f'xG:kJ,.V}@Z]k6RPh0=Mn8^U,zs	A0}@5M(w6$x>na%IK!]'}$5d@fyj0$&i4m,hYmsMQ-[)`d3f4]tvJ-i],]8wWpeOm<Ob) 	>1!sD-NVuu,{83lhi
)9j3U |=eo\-Kt&F!l"ZBQ9\0E%UEhKbuY^^_ZVN5RJ.Lqt,
SIW"k a[JibM?PAf\E[=^GOyUq)VkAh"]x&4?V7o[Empyw5^7@}`hw1k7:a-U0Q:V#gTJM2.toWGTlYG&GKrh~|AzOB[8	7O<
E[9qIBv*::fV?kCCs	Oj~L;[tARKA6GS&jY~IvrwO]9dF?B~Qbt	:<6F?OT
Azr{L/CyA;P,sTt3pr;;:9.B.dtEb !80f C)_`'`CWsIf@Tq(.~7t}*nQZhDQ
Evi9tdo13DBq+4f/G#AQ9?t(YQlPW%+<`6*~YCL$^^<TU@ZP4k%WFn~SIe5d&JTkh3&&M*qcEwSGIq:UU?SvJAN4~n_fRiWxMki*MOCye&8^i>f<,Vq-'>+a>"jc;+ctvT"I,&4s;CG@L{(m2\m4 xyH-mVogpBDQlN<cO?$_!@HM)R0,?[?+\(\:-}`@hl*g^J
R)Z,zAmC&U:LdA1wm
Hx:H(CBvFn@>(~:-@6c%&`>d4+3E,8]}0"l"~2(43(>3S_2%&Qvb[|5Sk4tz\s-@
>'3Gk)}[h7*(xd(w3m`J$
U$	CxT[U?P`UplAe~-/J0^`Qf^Ke7?FDi3<wUD0+i2XOs('*G;x1"|x8a'OGu5v`1	4@S)/ 8tLC,lz
S.+g)HeW;d0@4C_tzDg]"xh{W:#}Gq+bzo'Oc[E{u6
bGB+|8`9F5$^4$#aymY?JJ'h"6d@_F+\&FYVS[pB0U%`)<RM"%bi+oEf~M(`RTAT*jgU<<K-.<3M4NX3NzSe0WeIi*\z+n[S8{wDM_	H%rqxv,2	>2},0cCyc{V]Ve]o3Ln%2*pDh7[RP5YN/E$ri%r{ck*.'x/y(6yV/+S5.v9dK{Je4jGo3Y.z$9x1Jl`LTW00R^OqW1bw0}d_|EbMI@a`{	v'+k(cz8GrEi_~$_K(Bn3+h7iizV<08EBI1]\l(PRv"dqn_O@^;`:s);|)+	`]#I|5Ap<6]c9V-9G?^J^S^>9p0|m*eT!i]wRwn@&vBD4GUa[?*}~d~4zWF5^L1L]t`Hev\BdEdTk*/v867o1)V;xMC>F T?DX"q"r	iIN!nGj*dP>0F}"lG!+VUL\ct3Q!SA2@cu92UGLFnZYc!+uGdM	@]x\ODOL1izsUcsB[!w|eN^#:j(lVO)/&&}I1riT?V%Ww2KPKNppHS2<[8Ic(Hg#^CD| T0l!mFeVTNE8p21x(]pS7b7}2xR\)(e:N>iDNY`]q#>\
M@e;Kk^\Z:6_e0\j}X6(Z'>=nZv3:R|:@_RzU^__Vavq0\KgbIlL).PQ?_>8LM;;QH*4p	8!e8rVI w09308$J7+B}(7~F)XN5Cl)gpYS}7SG00iMSBZ|q7?PU]t6)ub/EpQ\J$u(1k];-5;hF,V{:J/9KY,n6uiU+4,\w%4xB0,zwI53Q)6=U%Up;QLBoBnLjHd8tPXU;c0jl=zen+F.jpa]TD:sX4[(3:k{= :cZLxF,AQ3{pbW8d0<h&i"[]TSM"&_.53\T}v	&p=R@Jm,)Y-gczudx7KZlVR4Eei;P$=0x2F{Ra;?(_fh9&l\X5vj\#y;'9GIU~.']*/}XDq&-O8US^u`D9f\fJzS7O|]";-!V:=mW"Lcf;OE4^F*TUn8SbFBd/=$K>)wEI/#~HiOQrPCt0ANVb{8NW7bL[:R;w6pEM[ 9]5hmOFJ`Rq>OnVFyvl<[4vw+q6o%+Jfe&o>1julG;mWm|fc	\-jzRU1@=J,b[8`ijQ3@oQ*(a^#ZZ(60}bQ\1k?[a-
-d{n[ (N?:n)]o!cR;h]YRM1ygS}X;v\b&qVi/y;[}2&5Mu%Pg7$iu9F^@\7|e4> 	IEF1$*f$J2M_ajD-_,+Ts^+{g"a^Ms
_p4T50Z2!TrT'`di&G9$8=fy)\GRC
;6*}3Q?	/`,.r'IP'3*:Wv=z@=*t:	o4|TxmH[84/dVb~=|8|hJ`r}O.7O~'VH)3U 1KW0*TCpyrI@EV[h8NmX)lxc}}KoZ4SQ
1|!d3-Sf'MC0D|Ph>1c,=vwZ=h(R~tIF~S1`X]>UrN~FL[\F|xG|[%/'bU\Ti	YRP/}:i= nQ]Mnh>l*Sm5i.&Z-VNUyZ,8X	;^d}#-LvBNN{f?|.^]7/*GP.0\qHj.l+rF7C&5 qNk!3mn>fYCr/JV<'}h!/H)9>KKDa:TGcL	wx	_rYPw.;Rt	C~?++QGl!/:!.oA8-
U"i@nrbUnLKc;w_n{}r1ziRl*hLHkeOe(tEykaQ08jbe1_hV(PchBu"]d!3=uDl\0+WKy%K1zeYfHCPF3@W>v[IqzrKe1EMQ|tj-_4NCc!ZVF`XQ&Xz%"et,_q(\TaYEIJNUgCT|TGkV^Hhmc"0f%cF]BII1{fW?F>E2?iR*$&~E);pY_Vqgm`9Xg8|P :[3:kwR>D%`|O8g^[rELHBtq2ck:"=r6#FCh{/|S3Nw+j1@^BF5\. 6Bkq=b]6UUQSdj8Zkit 	@'%eGG6[jghoSiPFg94ICDwY{MCb!PY|\zF6#4+s}t(@5Wbd`7L1MxQ}qq39*6+	Cj|47s\rvu'6^m6Lin s\R-z<YbH{fsD 5lmd,?<'Wr7Tv/F+
B-<w4q-tl=q"*iJT93\0}Rt)m`:('4Mj:-v`0SiW%XXCUNxc0:[Am.N1)VV^,H<		@CU{F9|:[uj*+H.q&tudZ_pt+11wi%%d${`t"[moE1R%5H*IF>?)B~|yLuQWm+I3/;)zH}isO	\%^J$8L}*5A\5t?{Tt"('$!'5c"bBbF9j[AEU,+c^k9 =;h7t	5"R-S$DvZIvLq|$xS qE[):gm0m;9FXX}e._*|dFx?(n"%[<jh^
=s:rqMsnc^X$sXb+m@iv;J[R.@HUX9bIqfrnp13q=T/aX?d[_+>iLaQGwA^D|vKQt42'#.QW*{F4nFj:#V,i8&pF[]&UE4
Z@{_Fz7j39_A{Gp)E'&0l<7vg9 l"E%v	:HGw7k{.vZ"/cnx>1h ,k dm-S/cX'2+Qeu;*BdFUjQp wxt[	B
X,Ui[c|/d[]ZoxYdMd4vrT$8 *nI"?\Q1A7!^OklrHf<iuQ)0)os,{J0
=$^j`P#,8v0m\#7e8~B&~sPwF^C41SQhZ.9@l$va5~L.5Sc&PzQR _t	lgb
LlPajkze
,84%}/=\_O^2/q'0Z4	xJnIIMl8],FDK9|~x8It=`R:"{c?](o5xTm?nY5-*yxK[&Hi?M+2X2V{nk0S#P~F$%.0>quQ|<{IdUXq
[N=GM3eTC-\yR7y$wO$u+ Q9e|!IN6YUwCa0_-&k`Vr][.h[O#oxO{t_NG0c/;lAjj525h-{
O~f?@/wHzlS>|#	ZtL.=uF/Y_ljQvwWd 5&prx%61eyD<5)S+h	|{trY~2jpx$TD[aP]$W7	z7\Y1-D#(EMOggsLV^Z
i-Tf~^Z}=HU;?t}BxIQ\f:`."H7fKesyoL4J@x;B@"`@z0Esk%KHFT12v~ide)E%b	yGMpMamVlpfZ"y1TI8L
8pcd}T9Uh>*VRExUX'7AJK9"=.'%BJ|c0l_[;WEG7'H+G=}B[MM^?7QEW69H2SyKr-1CKH6u4!AMrzKp$duTltP0J amuDQU{%0_kA;CdQ`Fo
,aI@rN|	 oo}	m`D05Gz@rEJX9<'c~D4,fu8QN:j@~zi#g)+Y-,<*z1]Wx7n<YnCN[Q!|[muuyF}6v^"F)4TB~jVi0orRPf"XOHZD	m!y'
189.Xinh*64VMuxz>u,&tWA\wj8Q|);#%$gqy?R#k]e.68N8MeBk-:\&\QEcd|<@/o}s(8>in/%C`--sC`ltlz/zN0}I-
uSF'9L|~'FzNbxK6O8x7w\~.g\OfX+f':*hf"U .w<e9"Z"e	p`S9QOf)M,(m/FKgf5C{{@wa$.SOw*s)Yhu<lT[gT:{;0H}73f*dh=>vNY)@aXr.'/HyxWC=XF HG&e$/2+I9c>FJb5$qaO6bd5q'N8(.@CWwNO3?W9t`!kiE0&lMQQ[c5@-b?i]'F+yGi}xk>)nt;I1{4GzOthmHE7-~y'Ry)%^bhwm8J/K;r DU1tNRAs$*gjG3gx(p%?@?T>BbjtJ#.MX)AAC*~x@zb>_X2@7<.5tqmkB6']W8\olssrh2Fl*KOz-m(|dLju7AUym;.-DEA;dl1}O#Ia)`EGVVjTY_)mjA5.YPFrTQB-,s'$0vZ^tSzk.s oampRN6:5tp_
NLghamE+.X:PXPhH@(\yeZ/s#{A~OTh=8hQ:alhXM)pu_SNIokeYM5HuzN,)jKD$-^A/_h[/%"2hit%546H)X`viZG8R.^FfI5Ng^wUCH+p,*Zl{d{piBa'zhpaUyT(!w{4 Yc!sc{sWMCPrlY3(s{$4W2,5rkN">U{_{o2=oozPn\X>Cq/8 Ctxomq|x;b-1-=QaoX"9/S?xnCc(.E3O,upB.R`!MX+t3.xIC?OIlTnTzzmnJW+[w$@q"sn}goZs-agd}Y{bV_%8hK4Ru3[( ,	<?6@RSxuZpu\QP|2Ijln4da)E' gvX+`[C w}\AoRJ8R.9wX}L`-Sy6z\Qx*k4Jh70"
)su"c~C.@cX:aO{%e]?yf",gQl1.MFG7VC?a$No h#Ga]'"3(i8+V0z\M5|?YU>\3;}51w[!X|]'W=mFVMP/i6L~
SX&0;>C:i8A9u"TV8]
-$:
j2gnb29\+Vv<mZpu]>\manGI=ht+s*k<p
S*e9b[z]xdk`a-aC."HEf'/U;b|?DZJ}J[upw+uQ79k0-k4{'I~}-?{ny?w@/
NVQ,bJ=DPqZy|B,0j wN?@?Y7YI`u}O/ozZhoE(T9DoC6q-5' \y&0#qw*r?rmA$&d(.[0NLM$$Tl_*!Jr9X/@d.NAS1^oB%K(_xpyH8=!vEy?:!PjnO3qD^Fp~*+y}R`&Cfs==c4\[7-5~e^)|7k4'L$V7t:MynmSc4n{HE59oQ93>Q?MPJ_4x={	L"X;\xCQQLk 	"B1`'vR%7IGR?_ ;v?9(,n	&j2x0+'`,,XY^<HkKv\=s|8*l6yD>4iCQ@AXkN7ksyGb+N1hT{~Yns6/$5^Gi4s;K^9%0xt#NDR(|@x[a~?t5: yqF1JY6p^4R)$*-_aU{$zv=$
;,G?j(5V#wm2.>#
&ZQ|$}O&hw)&r%&,58a(yVb]k1-.ls.~q[`2'(MLiACT])E@}<c(3 ZN0kq]]Ry P)-iHF]`W=?HdQq
6Ns'&K^sN_8\xiJ2%4
@G8.oU1YR(?p5~~x.tjS&*(N&v-@y-$j}C\Yym}YTclSn]BMkGEq2d4'1~zLD	H/+,[b%_~mq)T'Y{3<MuE]V'm;)33xceTQ))SKn_CJ$Th({}|+]oxGD,<8VkMK7iM4!.P[^RX5F.,|xR;}%M|dPvlPu!iL#ag!\CX9.e@+dML=-c5i)]E0cEY.&j:M2vC]~XP0	=[2Sb-w)^on7w!K@yyo*(TimPy[MQr{aLF6$
nOQfS[%|bv:}5/v_-k2aCMaCumM2aJJ/[q<cfI|Y0]zxaw2pBzKc]@Wp	;:JC	j3_17"esxkrfy}VzcS`lgJMJW+/C*I2#`b93'+y4j7<-#ur9!3\-z!n9_g/IyEB'\x	6;2;o$*uc
?$P:pa)-Ios'(MDUgPVv:)!TSU6/HyX%Nr
.e8b3kb"qJ>!A;S'&.4hrdRMn0~ys`Z(?3{GR'agd9mEcY8
NGdjFHPuf.8^6/|4|]og&gNR
dV`?~elQQ=WRv&m*om!d.pN.= uR^c9]+d^1R.!z.\3oe'Vf'axxG8v5t#Q)fHSrv}#vEQ3ccb4'JM:K->zAl)1/z7~uEc`@$wcljM*hfU@(z5|6
'6:Wv&_y@_[x@aTK5]p8b6%yl)Y
9bPE&\l+4g#Cw|IfbMR}$}{rA{nAwB/A2nI|)-}?"&T'h_oUN);l>ridb91Wq.>\5m%_V]Ggz4}W/:f|#aez6F&w lWC-=a@#2]io[+$C'}ZQ}L9{%%7O=7Awy6T32ZeXtUp7=-^0m&NS[sZ%6#{u,G`L:qU%l]OSdPmSc$beu*9_mM"suEn)(bEe'QqI9dK;OZR<?l/,$3Z@S6u:xggM
-Av}yQCy{m)c-{X1J]
"4j14[sc7oSl?;K[!U'ogLhxw*>q6Ze3Zk+K7QX-_%nkL)Vo*{Rtfd
(F/y;c`s8(SFCT^S+8@4}wzP`"@8n6%_iA.{!\q
)64@::,"t6/O{4TMK"}f:]k{"oa%~u7KL)zMZ8[G:p68h.HS+cXovvU{<DWuhJcyNP	"Lz0D~K[plFp7"E!Z$
^XyVl<C&Z`}t]i?;4SrPzY#*;m%!0(y0c"mhxR"XdbteFik|7F_&{6u#;|Ua1lK}iHc#bKW	$SiC}CtZBFvw
qu`RQu4.E%a-~r`5>AeN)&"
!(q`'NVn[P[w=O$a-FWgYx,xq/V,'@	ISo):Y3>krLx}H1/ 1R!OJTPh+;/HA#d	RQkSsi>/.D$Li\j5\UQJuNBCj;B7'1>1WJP[zr_4-kj]n2xzxA&ow{6m;>C3I_SwG	{&8'c1@Z6:!
J1AmCHl_fq\X|P<a'Nvnp @RRsFh`QvwqCD3J$7LZXePeFBiwj)B\yEzb7$UmbaTz[:-Bo%?W"T(.I,\WoL)~C3\D*le5SW'hqW5P&wP*^>/wO`NOUuj0.R/3rhx5=>R6S"1w-d^(Ix+U&l9N^<^)_y>AxvGaV{m-X]-+bMi=@d_C\i|l*NB}FYp$:]m'xM#l$e@#C\/!^&$1-#t%=:p%N0QRX:RL%Ow=d9ubLJX:dqD>+bs<Fpy~rk"(B;rc X%
Lg;w&%^qTixCdC"_	Y1SyP,rTP}[-4mDJd'c*$C}?6C;^K":8w:i[\nI.$7
&Sm.QHIhh$wUH[27CT>+TM*C6XSYC8zZD~D$	_] [Dt1'ud/rU#49<n.Qv~	K@&TBFaq.)cfLP-k`-LRO(y6/CHRx2]F,q_$CI!nKO.QLPX6rKaN5#`c]2PI@@;qnDyMW\Z/Y|)!H@kozU0Pw{F5KJaZCF]DG?#N|R+m4$,W2Y8OI%@~6\`F#5nh`mo:D|Fm"DwI m&CGmk!CvlPz$~RQ@&Y:O\$1]&#~!=ms7!yRy}OM>k'XGe"IvTBO`b8mN:K6vR"knS;B+z?BnV
::qe"L]jB&jU*IR`?#jD_2bFP1a@Bd!I#=(\o68;r5S%/ca	1in,qC|#'	f_'k+n?6PM^++tnnILF\nXLdo3>*3xBvZ>hFL52
GbIp2]4';6|7,lMH2bAF"Iv#]fjG}$x{^Lid=(nh-r%nCs=*[LOOI84rT.F{u-d
'/4;kYM`ezYu4P7'cl'%5kagx>%Bcb|(MGf6T}$I1+aJj(5W{^#t=wY@%dcv,c58	Cv7r-1L	Y	Q_:Q]&.=h4UNxkzV?	CZKIM8O\!4lS>f+yN
hi)<=?~-f7\/p0nT-6H^:_@e=%L_IcJF`bL5$@'`~b+FCxZs
W+*"jzkoci:FzWY %)9I|MYl4X
@M<y7BKiQUe@wEEs#*j1[92]jJJ)^zp[?p[''V2fN$`\Rj'"_pj-BQs^Kb5<%bz{"bamwozGA3O,hAT
iNJSdJQr|xvlk)qa	\$xB="9XN`T]^ng`$|fWkHB(gYvsc@oxS\pR.y^OkxndA_`}nE6rvS{lDhPu<W*qN8&&$yCYt;j1TK}R#D0g^#e:XK6|^yb%?DX+8q-k[j2gNI6KD9|JY=kL`b _EV+F'CxQ;O`k{OT;J-s#G,"l&=*[;Xxy%-"HP#<PMflM'{w86=MZ-}DPQ~'|n oPvP,5P{4xU127:x3I?"zo& 7JRRuof$i	i6]PFm#	M"Gy*d	a~~VNs-pW2q"#Q1Xg$
9&NVm@tF9|(:tX>)F.e06JGa(9Ny:
Vk!T:`vA`J5tT;1
1:B
)/zMXudvCH2jLMbW!$Ex>gC.q,j%8^`2/GBodQ>Oe^>Z,6G@#eWEQg2\rzauK;!,Vx:=VA[cCp[k._v|*8Mdjc2zMZ2c31HOMpdW'y=yNUj85wXSkA2b\6;PM:641sB<chFGE!QF&mD|NGC^\E4scd\9NmXY^}6hW(++af]|2frG6 %Kht)3v	?oaE1=EI+^&mO(wO_g$;yL&T	[%hwLU$Ht
?;nxMO.Hd8i	gZ8=uL8vWdHbFy"E7;P=c5"n(oCa86`3/	nma	\0IS9aF{X|
S,EHJj6.k\|pv8zb!{:QwkC?#<!8Eb7f`@
1+N /kg}i'$-MzTilWJ0?\jiMTfTp'9'PLH#|Z	IT.WU^3=V$T!lIO +('yX9TYix$t[.2e?7Mez-Zz2wB-o#FKqzD-5V,>
XIow
k}-Mpo}_&)@AEyPLKPO~bF3@LZ(^b5GDyE
AnwKcO8[oE!SI~.RFV2E{4@WJPd1I7+Mep\]z(>ali<sC{V_0MFaS PXe<x&X6!bF-=t_@a/Jx_+ScxEj$<dH0	a+/:/C^ Nfw^c?4Amw}9!DaAXH)Ce/Zdl4h?iZ5?$mPBfgX`o|{(2UHfb!GhTs>L'KzG[?MEtO{QEJpMu.s<md!3`_{"yF,jNj,^V9svN-oOvia!$23g0M+$[HOj*9TmrAD6f1p&3--S^	T{Ly1Z&x|RW{{+OpU]@k4n`3VK?iKi4z[H$+ 	#:5 4K
F+I58I=,7E:1pf3:xq|Z$
GShB3luWab'I75B%/[k5pV[j7,[;F2laQz/yzYOipqR+#48I,FN*SMWf
~W='|7}/vI	cjL{g_Dx\~lf}8W-&.j&KplkJf8l;(I<lYlXoU
.35-Ka(2q@exqESLgQ1@{GmSXi?sJ6%8E!9-zcMb?`~Pw_5yP0T(ol{GvZ)w\`~r:9(+ M`3|`}~LNn"#k	1Wvd}o`|#"pO'1ws-q
ku22F83yTlBz\jc`Jn2UA}F9u^Yx]UrB}H2sgrk2e+LEw-ZkiTt\Q9i%eWoM&X.^/BOW qy !]hJ_{Cw?}\}%N7K|VofP;bLwVr5R?nnv.osf)sZ2Q'`J#`,\AX{+	jP rAi[	2t2B~y'_*cq_[zl#riLIM9hnM]}I$YsK?#Mg2.bJ^38nKhLglk8EXz_k28Q)`^qtCU#DSe7mGm<WSQcl'(CIjfcg	2}=EZ2QvZ.Vz8r]]qnb!W>PGDx"!p*!%6F)(:AsO'wMzt1&cH=9eRz^QJ`v>){P&?qnYNLce+|x<xd4>Qnf$p!F7U~TMp/OIMeH4p]:q/LdQ_|9|j^(p"O#Ge@|'.`zdC"Z<Sr}-dk|2&@^a	6Dh	,<7eY0ey"h&5ejI eDjk! _Z!dEn@.5<9$!<
BYSqXgSjbs&+E{5,MymHq4]EMV0]+SdfO$wp~F-.SW9R!A~;3tz?ej9&$M1{MY-n-k-=S5--|\`+RWY@9i'a@R^d8Q[CizRsqEhXvr,WFoq+WlK<~wgbvf5jl-:PUi'nx"0A(p|ambe5HqJ3aC*%xvxp|5x-qd]vx1d|6-#nAh"h|jcq;Y`Sj16kRoH^C[h[SH$PjN29_hbWx5MHjbkFtINN_km_?+~\=M^fyai^O!0/(q0aCG8smv	%w52*:<(9?LFEp8'E/"$`O,p0^}j
$EXrl`WpNtUnO-*^pcI?NqI95*0'T$_ gVeK=u9(irw2!60jTW!+N'e"nv$*=_I(iC@"w20Ze[	69/OcdTd9O\l6B|pyb[
A]+M!fV-RayOxjafd<s{,Q=|g[Cv~(f0)^TDfrbS4u{igA%vB9SH2.j]J0Aid}wJarb8;i8Vd_BH?:
OT:zV3a$^0M;NIGhBn1_H@qi8H+i]q[8SEe0H(f	-0rWv6[YK? E[UC6!,:qld`z<0/cUKGUu"(d	i&P@g,_i1$uamJm"Iat=jvaTLB(ce7#Ig=&UW"eQ'Mnk$Om}YDw/l9[onI~K/]@Z)b>IDl':lE!!WAN,"An5TC]f{{yI@"fQ.Nse4D|W$6$`i]gbD~xQC,nbRZkBtebUto}Am_1<fx8Kwd:G1Zd+p0+ad@,Qv>n+z.~F)eq3h8$Qv9Y4A~X'MjCB|<XeM%eBg9=VV#4P+j+B^RW-*=$nZiv8_,KHyi^u"]4r':5z{`]{|A2TOG9<kP`#3mb-C++Xyss4wCb?uq^Cf",?dzP"}]?i	{Tk[wYQ/7I}BE*tKPch)<=#J0oQ4hS(@TpIgf[(!\0(XoutoiU%53YCC]fMpsFPNQE@0|`~}{,
=9,)]|^0zhMxmW.u5=5Q'Q56+bXg:bx=wz {jWtl9}7;%Ue`wy?w3{xh3&#*AR"],!a)qg2O]5fHdT`,):>6,Kon=0uXwV W-u)n/-C4&jq,Y]fe-8z]GkJWFjTtUm^F~,FESD'.AsRUTC{w=&HIdsIK_\wyp9>fAgt4j"J8Yt(vWAvXk/W#%0#jq32@}`j^_c-7R7=~`%XEwg_zw[59e^A=@Y({BzgB0x,&ip(.qS{g6	4]$j4y#Vj|X	hIU8UfwL'TR)?nx<%\|-Wwi%=g1]v<^uA:40+CyB)L.w6Al?f^*1K<zoE-v/JE( -yt%6uw3cH&5yg1rAgR@f|+st5x= T\;N\`PQ(?{A\3(Ux-vUWski
A*eZ?lix+pydb__RkR_7zjU_Lfm`{Xg\gySs#/|iHeCV Ew{D\D!rYy{%%)'Z97jPnvh=i<JFtcV ]zR>z4yPE)FT!~Jw(9+*:2zmk}TGn#m`8hBD0&b%vQ{?*C3"qC9!=W|{{+	pX+r36,afq}})`
)BiNS<JtPj<y_u'RxjlgWQwbne@zW*bOO|j]{&#pA#?<YC1m2gqi2;``%B]r,m-ol<!Q:Sjns=]dJ4WJ@*4({0sje?XV>5p1+-\;CVCxc
I:~\aV~T2i]5lQo+\[H>Uf(!+y' +("\I'#{t3}v3W~C1|W{BN}QZv2TYUtJMg_"s($`d&.\H`d|xH2Sq}|TlL4GE'Pz<jz.`jypj%AoHSGN_60J	4l:JTj8hc%5M,ybOQ(c'7S$2mpf{lfK
Z.yoh!:},*k<f~IZ{y1d'Md1Z`cKfaU[0jjUMpoM0rrgjJ*{8V|i$
z@eX] ou90uGf:>97{x|r3@}|Vn7Tm_u1P2nS#bO%X3QUsaF#]<BNsWo`\`=+`5:+<WXkV5`e];1/v:dr4NG{#3"z?&XM0GOZX]u2mBWj@*K#V*yv{y%+MF_-)&Tlp6!F?sofqzZt=DdE6w[l{
YcJO>d&'DmyoS^sB0>=_FXUR-vnxWF2\du.R%gSkl	!93j|uz#/jea%Y
o\Cluj.'g*|&\.(LnEdfarMG~X.JAI^<:#Y?U\pBs c9+8ZHp`w]90rjp~HoXHbP*}d};=h\%X9mr}D,kBy~1D1#R<^};zh6}?'r%vQ$)G'{1wk3HNM6-(Q.[4'oO#_={+3q*VqopOn\_n_*?p`I$!s
|-9S [x)~ YB{VS9h4fvhp\Uo'h#W:8#
{zv"OLJx@6Jvn^}UyB4;9Z2BXeu$d!RZ^P~/d]<zjQ3\uO7fcBm`KSpSt)]S_DL~~@`$V|{[v]w(=DLDn
.v:(d8,:	d^6Fc0GA6t\bnlT^*2kcSJrj4*#Ivbh*sUPYg1'rH$IT~%[5JyC|(Z.O,U3,(nQMOfEdDph?}lydLx6r#W1\ow&4'ta{;#T;3~(kMzulSIw4[{F)5.,&(C%%r;NI(	tD,M-[	W061G37bs_P|V?[)lCvczk/)c'G~R?c*@`?[p6|:~3 8l)'8m/x(jWi}7z<^!BZcU"h-F>gS`
%ADpq'Z~M.RufS}SU;-B9=E)@H?=v]6 #6h"Pk1tV'UZn+z/R5Au+>	(Bpu(<?w9j1Ag#Uf-%p;qZ3{0Rc~.wN	v7)(d)J9.p\ ]@|P}bs >bI)N*_N@^)[jOY\ha0[cZdWx70}h|tlQI ?gqid^!pcz8Sov~^p^i?K,nq>W3tLt[7nNpc&m.WDV]>JXM/\\YX^bx{~p'?Li[u<Hr%zbpg"/L,	Tlb+gK~ +9G2j$cbS9'ifPBm&+{y.HEtRMqNF voS+xlL#+8u2NY;h5a
u`],T*F1X/~i	3Bo0RA8}!D?biPA`FqiBt1gK
C;@ykSi^}oS+B+N=WHQc7R94LqY^wDn!e.]2D[~r}j+-L{)Q+R<#?I0}yrtY/)ZGx9qPH~|5wb+i_+
Y_whj+dl7Z:QN\"&j;Fu&n3e61)ul,=Nw].p4rblp%OIT:qj$c}OIyUAp
5nzA)w{uqD*}o*4rq&W?U4G>tS:D$be6**[\.X/g^F)x%H\:AbS:z$84% LQ#O"K){Huw	Gj,O[Rz0T~atgu&G\'=t-XC}tu!3
'Be[^`hYa 	[/p|G:9-@>$6,{)0,3e&[{_&?cHVX!
KJzChL!e)A_Gu{fghnX-#}>,bZ&]_`Tw-9@3jMOWVw gr4bAd^,6lzI(3}kR%Xk7]m37:{plH}:0_?e1sllw,@W
%8Yxy+8/7<R)U5dg1i(P)e!@R Jgh8Vrf}tBlti;"8EpYE5b}l}0
~ui4c,jKdrI=lV%2jOpO6r0:qY nD>9v)Y$]QK[|'k<`,h`$;7M78%{^lg<;CeV/rx}Z7FR=oZbHTUVOJ;nDw!U/C`[?_@4<OcZh$'&E!NS=iJ	Ef$C-?*rewi:b_XU!|#?Ky$*&kyg)riJ

B'rHt-Fm$yxhJ]u+z E1LTJ0w{Kw'+]1!rwM7u81T]%FBV}g?q'1`wY%W^SGL(3G%+2']#)Y+A/KpI=t7{eIUPt{mb)KoLB|LW
ss"_w+/124.akjnZ(<|ok#=F%keURndS(tU">H4}NDj}u -CYL4BaR)v}Q6.|av*QtROKunVo4g,@)6yE3,\N\utAZ8T5}D(:W_?($U6R_&Y/$$@,'F^(n\zr}1$oM
;Tu-i?7dq!w0*J5xku*})H#sOT@t2By	t?j]e%&ZE@y
lFVq?4'`xkIVB3r*W#a?N	Fe
m2@?f#%,[\Vt^d0x\=C>D2b#_;k1\%a4e'5Rg(OPU'Ie`G<7}T>iZYZ>-`<AytZ|+ErSz-	9%FC^H%1uz-2 N082,cd-a
vT`I*Rj>Lmv/^_?I*Y>c!ium364|LDEx}+aJ(q9%^g0shOn'R&`}UHC*U%$G~8`dHpSTr2sQbE<J<H,\0(8WM3"#wd3j+p>!*[`UU3m3,q63OH/Bc^7d t "~%[XTrZ[%*fPEia
H*
16kmyR2P#BcE$e!7	-ajZ5IlB>
HVT};sx<vtYPw`m_j>vt6l;ZphTE4\mCXS}]y|M!]X P^Q I&8I9^rZFN^BBe$2V;m0]cPps-rA<q3S J6I8G]}$Q]MBW-{<!q*y`CG|G5x>GBzw,Rf&a"Ua'[+DDK`0$8-je9L(,w	
j/kk(a%fr/K@g[]'D}*8r}?-5Ppe oz=:+r:T;b5Qma,WA4PJ 6	U
Y<g+cO^ejkV07Od>iYt0lLPxK=#a,U>	AaZ:2\H,w-Om^2_6=P>"ExVY7?URD"5d}"8R5zL#m&(X{Hl<5}0~v
Ms-RVX=fg{^'"Oj?cCX:5<2g8/GfV\$8Q@,tXc;-z,'gE`L_-_f5u&?)[Wt*dIoT4	4ov^H;|xrNc"^#D&hCZE(/Neh~+="y0`9[`h'[(Pk,4K_l#B2HT	gxsG^XHJdwE
o	"\<YV-0,/.'iRA#/<1+5,dh2X>7RfG+]Sej)E(~@5X;q!"Yh$7[r}m8Yu9Y6-aR~e:n%
]\)_YMN_`Ek}L"W_*k=O0<8\7v(*9lH}d&YJ`(WW2>OEcecS\n3EJ,0	*m&*LSyx%kf2)Xv 3utXAI'8'X]]X2O0xZSI`B\PBbU5(K.X@Sjt"q;es?9/{s	O/Sopc*&LVRo.,iRrl[Ed6T@0@m-+ p:~HE9".=r0b@{M
90UnLb?81qivy}waAIM_>K.7$OAr"DF5
"=<f]BqErt`avv"/P?dA"a|Y%};c"Q%5^{.Hx.kVM_F4#]vSBc^,p:(sLQG?/h4&uTuACWxY2kGNE!@rdyH!fj5EJ^W#XQ 9}d`}M@4#~
8JsF"o#sLTJcKMpK,}x_Bn~bBKM#QLic+evk&W6
fG"jrR
'l1N[eao;^gB3echap;V_C&U2O4o3hp@G&H=x+s2!CC;A[-IwSDL3ld| |rHQ:I{T"7,crgF+&+dPVw@J*oh]1[lWx(]\7+gI6AA7PZYHG'ebzlU>7/_k%OwZR632>W/u0Z}Jq5Qf4DLf?L7I86<$
:HH~qGtq)Z5QCumR=Tg
$0`Hjj44q$QsStmL@QVA6SZd%o8DRF7%|o4 !BO|,1 j^|v	e-$7?(oe}xXR*M9?mmr6bhwY:P|ATQD%w1G`a*(&qp/v|\4x`k\L0K8!?c1"1Rolr}8rk/E ==_mCVD8iWCg}ZWXmT~.*l>A?2qLgl]qk7bWy%CK+^0&W,7#~9q91rS';,?!lY>q^"U-l3Yc17w[~wA;VYBn)f_#_P9n$$[FkDNgUB>~ooaya.o8rS,"{,MHzu-hcNrm[*ISme6DZ}Zta33`\[C26J'&5DuDcEM|C2$V)fXQ	 APww
.L2r<)6xnK8Y'^!dd#p.B]=~L_mn^}_}sbn-8d!s|}W{{q!PW$.k(`XobTn{[Q@o@r2xZ[Z~^(4)xp2\3koz_x;(7[+zy!?DQ=!lux/=Ja|npE&VzQ_H0ictWKqzzTI$yXo8y.pnTb;@svUzD{MJY'lDY
Yl7Rb{a~aNaOsMEii#S^c58lGUp_"x|'WZ^T11TE>K/5%2nGDJL*hm-0(eY8wrN&\LH4wP}Q1?V*#MtKHRKB~<hBnowB+KCs<BmVkp'heD3`Xr8o3;iC^>46RhdUh$ua@k25hi_tE<[Hz&u+geE.JWg'Xb^S<,:io\)s;k}MmpR$zG<@ 
Dh\|0nn[]u2W`QnaZwk"Qmj$^2nx?;hH&Sqh({6aMKOGi
zs'%[kIlR0[776cL\lR&T71*y,o|Mm0xzI[a(\{259	7RM:_gb0mxjmaP/}+6B#x=eq\'	 5V>>$5$Gt=C0miYnpI[0CI*QlgZq,\GCYq@(iVB;
44Zvu%1f=qTjrR]!R3?zq9t>0hb]Ix/1=T9d)C.:F-U7iaE;`7Y[#ezB!RVS+=.aB_[pIA$>q$T"E3=?+	EIy0M;`WuZ6acAq]BUo$Ao	V]G^<Tr=%izY^MoYh^w	9]uZj	Q_Ler4$ZVILDq~MooH`Mbd7Od2y?EY~n;z*NA$0C|~{`'|>G|H(ineo7X:s6ZN<tkZyQ)^r>E9J$@&xqHRlC~?HwdN NmlkamThe](Y`)~zD& <fs@R*u&&GB>Q$ -^79U]VgYUvPg[L".O1o=d%%A i^q9gz($
[p=Mtf`S*RtAkt5VabDcg[3sg&T+
4l&(kW9MxLNz()3Ll{lQd}!w_"B6`yl2XaQ1X7Tz~x;.y=cs@]{y}l[r@\fY$~xxXDq1ZM!e1.w3)'A)qMuYSL\72+s+HQ_jkp2U]br@Vlx2)-1#iFKL"kJ	@v|ipW21[D2bp<46Ru~S'Cd!rw,N)4Y|BBU!4lT&noiG?TqB [f)&==R(m#<3y2LQ$>=<fEIY^`(8K2o]}0OuaK"m>8J2IDw{' dVJQgDbNR4[|!M R47:Dau#d+]6CRLs!fD`U:N%KADsA#;7j\M	?=VTx^7KPYqb:1MKMDTqIy/jDdm@7lvq
s2ImsSr2irXdQH8q:R}j$sYe'K9d1,{m8Ef][g-y&w8<6eG_Cvi.thL&vMF<=a,"eF-Vzd.R!-)& PBO\Gh=
AZ2dfgg| m!2N9p(	WxMc7z6a_V)Ac{NotweMY8RXn[,C.	z*^ hXj;9xCSP `<i}|UH!)i3C>~#&{cY82c"!rY}?>z,8}7=~OOXo:bqL)2v>`C*Quv:oX0Qr(z{,mCqSgGn?	CK45R!CEkz,=D/Mmtj1k/r/i[#{K&uV5d<h7U10+v,hP`QkDHK]	>zi6k-"-/p>"1	WC=Ixn]2].pR*HsR|lA>Mcf"/x/|X9ihU[ A@bU4>}u;unI588]yL&eN{pQ%!\b$;gl-' #.WAdUx"?5EBq[AN#${!`#PZC.E<a~[r+[{+	1"X_&1cZVyVNkp
A8]gSub1r|kDyvh?m}o-Su|lA'du,.MaMD5F}#Sx=8&	4XZn|\Jg||[Jw$Z[Y+!Tn|.zu[Z0BAW^-rqpDlE[,lj3	^I'_EKP "=iM>h~E">4P`?!`MR*_H%-$tHP@bNDWu}-2D5GC(xjb-|j$qm4l$@l?YP,b1<C"Lrr~<aEhu2G%pH@Zb2zNB6iyzKVW3f-_C"@sYqC~%w_=d,46F$nZ
_Os@8C`v;X`
${^Qd:n[Bha_ss`&%9-^gG-X^S+n^j/,Zm,sO+p"AduU]03lDB/VgJj7RJm%5dKjsP6">_b]U+&4yxewfwrfJ?7%FqAQa	5*T*PkJR%9J/)b2ufC8QY/_az>Hx/7>M@xN$v11p9mnfhu%
nh0w$x"h8%7oOD7kMv6D@zzuE-; pNZroKp9t\NcU}1ZH{deNjPDL^X#Tz7"/M5':%!6	JI(!~/'\ZJK.jvPM[!D6G9~v6VE~L|X0s|g(X/s@v%qH9UtJW\6pH&Q.+q);{sOXk;{OFL'0/Afds@lVS@A|>wwcs W\#. &t`,U<#T-} An]oX#}V"6"+LM,R/2O(Q-2A"l"o\Md)bI\S.UT*8{CuZh;lTn;gg_BfCWv\%n+|rdP5,SGx\Xdc+qa&2gAO	z,ta6xLXW4-SHl?,QI^T4lf+Q$p0T~~^:[\S$I'` a<Jzb:T#NTiUd	
{`Q['.5-;3hCv8(P!O+M<\J]l&+`= F*hYR]?hV?SAFv7+iJf2 !DAtaBVU=Hbmd!
V\-R	z[D#f[k4FzHeS<:kK,m
[H=_2QJ05w\BkW:EQ ZNTFx<(eA>{{M+7S}G 6is=Dmh;[).#CW(]eJ2\rO9v!n%ee1Ti3wfR5%MRNK8*/9Hq|T8F;C$ +<GWuIRVQmC#.QztTA9ZstW+0bmKf'fKldQpIw\8+n.~0P<5LngQ>)aY1gv/L9	Bt%%p;Bs0ti^-BacTk$n4x=d|f,!;i-MMF3L+h>V}tb`):F!];$#\-'}3.qYx!fQ	Fo:o$&j_LVq%5egQ-UA~?X#\?Wm"z$.~C;HZ!{/'T-D"h`555Cx2recBV\7d6]UiPL3C'|$KR+i$-N-n.wOV2xaH?0"E:6clhT#qMu,1cl>kPRJ~+mR*E(G0*+Q~-N*i1\TENYxm+1WPQkS\x,]1
w.hW0zX]g\C_Ei?jlO+r~W+x<Q
*Qzb}x/N3 Gm(67x/k?N=dy.Vhk(W_VheK;>yy0,?*#VOGAN<.aEya 5wE#&d#^VJ4w?,c}wPo|-XGPd'Y-KI\LvAr)B%wIf\q<9mfE5&rg]0S##O ]`57jdO?k0Vm~)raa2[aP$c1*iLx$)2?9&,;,q.1g5\<.1F.*6[EV20hmSJ*&mWGSw1=NgD}BV>!/YSGy(vjCt<s)#8T&TLkp#6B-|W@lpdGDZ:RT&"=W|i#V'w91 vx~G+V.~Q2J`p8aq~0j
K%,s|eNy)HXLnpw3pjmW
.tK>-:LVkEarQbm`l_I{|+(`>>les c!VD%O!%UXi(\^Z2Wm:`&9F'$x_}s-h'4exluC@"y![&/QMejv<2x`FoFCNmj^^$A>EOL_%8}i3eN{{}
O70"os\Lm,>]T|s7[
\uM^oj AI54XE
Rh4R-en%xtL3iN(4iR.m^U_6Go[@CusIiN.JC3>VL_fr${`d#)QWyp>_r){=YWM{<gCJlhSSO|[Dc [J3Xt[=+kauel*;>|Sb>kj-6NpyTY$CC+eZ@iWx]f.T$mvRah7Ln{Y"l@CgY(5lw09>-
_8~8c]=wKq-HeA	t	l|INYKw4Ey;=gyth&gsLs%L;TxK90Yn$K"l+!!t1E'/{~UFi"B@Y`)kO'35gihg8f?P8]rx,[RN
4mveit[iP+rcF4Jx(Kh4tbD<~PYsQ>Ay+REIx(n1(w4d;q<	MCu*D9JdW\EB_C/mO_vSryh%dUP5OP,@9%X-*tX	DdYvO-Q0rSfwT
[!~( )^Cth5RL=l$05[1}M\%-!Q54y4Yr?'Ce#R	_d|EsPu)ibvu}qR	XMm8&RrgDEX)07hkN9)d{v*
R#AaeOQaYPRD?*,O78Gm#.5xFh2H=c&'|9A0T[Pv.A''?cyqqM^%&q[M0>>{IxWPy
K,yJ>u/&siC"%=k<onSpF_
*g+rOWWgYLOUS7=M1c;yq0_nR8aO"CC])/)wKn2EJJcX
F>[/Nd'JR05~ {N+ZC{)Ls#r2OL.\=l:67B)UQ"Id/Jp#'OYrg75=kpWfy~W\'iZA15qN>C)!ye1OlWYXr(CCLrxIP+2VO^?Eb3~:qA.=uT#qkVuU+swO~EQ*Ugx\$g<[F86E9hasz(>yp()/UrBe
gLXUXN!_iP=mk|tcUN=}4f\Eu<0&-b<i)K&Oc1z6i DF'/MkK4i3=^lVA-5"+q_$Gt"xuo]Q#u;Db4=Wy"fPZ6+)Q30p$@yrslSNW[#v'=v)0LJ:pI&g3Rsi3<^t@2<#>k\7?"d&QaE>MoCV0UV,#Wc9em{
[5&~cmbX*i;I|C:7yqyPU =y]xv8	
 hVF2Pg".J@teuJp(l`CL68j_]&0`g8u3"3MUWY\P))W9`<jDZE+hB[0lh0U
BBh!5=\8g''yx;v{HP?\[j[BMBS8W(i1oy!7<Pz8p(@.Bb~2R5gch<v.dH2cdqT-x-]0'\I)H{
_q,oRS5J0O~n>_t-#e*N<e||eY^S#W-*0N	F'>18YD&'j(ya.WxcuX$5a$W~Xnca@0o\^J#cDTqHIjCS5CJ@S[3~aymI!"V#ecZ9?k5Mb/#KH+DU#cBjBO;L@Hvg>\wT|
$}J2#p#9vNO7(PL*,%u~2fA* nNXuV<#]$Z$U9{3K*%jq*@0yDg=hEC":7gO3	]v&Z
Hh;m>Dg)3+\7^:]2_cI39<zmWUz%akYc9[?cycSp&TquTQJOs-Y^;mmJE9-XSu-)=:*wo\ZB(xImFqRdViG.9GVh19pa8(7!A}pU|oWYjcmJ;Xf#wF@Ccv,,9aOe-@UGD\"e08\3uY&a@$]ib-A ;pN+nHACA>-2PW-M2r8k>Fq;6-77T7niW5Q^}hoU)w`B'a&PI8%JIv,rMB5}k]SuFf~$;O[K1J)7+io_uQzj(Wr~O=iVeQDg{^PF0|f5c@ZlVs>wq!+gz_[?\HI0KI	j}FSTDee)K^#X_(A`k2&Kv2R@m!. M^v~:k%d:Mq{A(PR6m90	<n~4N;.`n*d1am/S(ztaV2g.==JU-61mau}MR8c.~?f
sy=CL8=*Oe`T$%2^z%VO4-N\_#!O$3Dn' JAm8b."(YA5WalRH4F|Sp|U#UT=th;P$CCGDx\wF
.4Swo>SPd	YOj]_a^/-&}D	McQt[*Ppi7)Y_YQko$bn
n*\%\O3?MM]xv3qjrGjO?+"bw*k~
?{dR*i3}~h[!53-:AyWZUclbZ
w}%#\CRYZ<`/ePIp9b0|W$"R/b#[5{H=w[|M%6M@p16.H-pZK;g>^&s]xcfQnN)xo<&U fPZGPi!(6HZ
)m"wuRsgqCG+l1""X"A6iR#to'y+HaG*zr~z(^O1OC]GQR+pIPskg>4{ $cA.?K>D>9FfG8d|(,Ts\bgaD8i8ZO<j|BmPrKMwjwtixX] yv*N9
HPs`(4>}V#V{c$-Ku-Dz6PneoU<?@z:4Mgg8P_Fcs	, eGgzmDrL@mp|
>/Lb:I({(!FQ (CQrR$Hit`3s,*N>pynjb
,s=k@rto{De> PNBP!Hdj:Q}ESceQ%{rcScxB^:Q<=1Wpj5Oey+MwuiNAo
;eyP*M2wKt:!/+W-]X8}_kU	6Jss52n$Tp0K>HnNP!J~QI~([Y|G6[j>#NGhCp@$A?'`_oS?Zn)vb8VcTtBJUNZC|K&->\Ao,wa7^ V^w2+f[-X;%C^T~Z_S]\^Zo)R=/[IaAd74R{['7Nw"u};#?$(_i%
#2ES*z3bjSG#`IU{s8-/bPNW$:>q-(AS3Za3:VrR?xl8dKd?:/4gBS#KdubG^),YG-(M9SND&]FuPPrS`3WQ:LDl@(r>*8oU
{uTctm33i{dimBlAJ2,rmw)^[cb)klGMS$vkVac0?X@?f'A"l6vo*{^k$a <&/r:HCWVuQsd^SzZCB$=j=Z,8k&n]]x:
PP3~Y- C&GN9;vuCebao_6+$7i'jDf\X)Va }o|TUJms'/9BI8jgd(T;q]BsnGi78KbfV43zchJjidca]/"U@
l+@#Zi>YJc,Sv;dt\"'UHC_krs&UHI7(8(GdCDz68q?!#>n>-_`r6H!QZ||$QEoPjwlC3Oss3B[H$@y
a;:{7)lP?~1J3	({aM`NTS6+!
`5P%}x?6eaW(=O_h,:IcADHNr:j8@h}!	cqJK	-;+nW+uPz
1YIL+!}.0&WG`{ul"LM*^BZJ^M<y'1CkRvk!/V;w/\[Mu4!mwQiM(B]
;n3
J9R:1{ypD7AqV"Kq:7+r_]4ER	Jp@`8RV2woPMl}h/pZA0Z%4wYx.33<8,% 34Jsi%1||vrL<<-=G#35|DEpL9K6rGCU$=Qdytlq~}2 M@:o=)GlKq9a|V'5ER}S"kAmA3J/=]y=}!iJ3+W#6%^
=h|=?_,$LG#U6RlCw5K<DUY,-@e]=3skLu,$kG23 DJ$l*05%(r"9vNu1Ygh fZ^H}rP3E(d(Z4N<<#PJ
JebQFh$^AxS=G+*_>iZ^amE7U{a*B9z:[6QR.ut%]=W*c?BnqmfR!j?QuLw^m=P>tV47;
H[d'zq'x@;iB<hgjsygP4r\\?Z\{:OEMfV{*>2c]&it "zR;3~B'H,,,g#;=VRtr0W^_%3!95{	EMnP2SPQQ&EUnk\qZ*B;f?P`8+jrQ\?tT$ov6XHZ-.g6$/c1BmmsoA7pl]PS/\8eK=j@31,7;7Q(pLHOux9DTkjpqrEzIgD*f]1mFFAO>DlT+oz lOoEX\rt:/^G_kk+B_6fI*isst?Og{#z1hw.[ [Wxl<wT!mq=?9kbU;K"l3fpR.1R/:P@LZeZVuTYSa(%.[c~z2CT\z#9+Msk8_0)$L:+ZL(\S3<NN5m (d/_L=U%{JI~tX0r|S?$oV$?s6cHZ`GsxULsB;Lp{	Y#v)m"J+%;g\`{(,nE6D,&'0YrMS+>iYX#)VPCZ.~-9G>:/Qb{lremGI8PY"o}_Sfj"\d-SSZV1Ul;/UG`(d=~ftW?;*])%MAIef8}%{
7VBLN)`Db^mN}lvvEc+E"y3`t?!(#[P"QQw>W'Ke`J?JqpLtJJU#LtC>''$[l<[/4K0&aU86#.q/`evC<O~b3*h<y
9f6|SU$8QXJ\i[>`FvFA,dGPbV6?&/j3H!rP1+NK{$:;I3^
<_JTu;9Icu{?=>7)3SDGt{jf)\8"GuE7e)@EI	4 LfdcP%,:oK*S7hgVYw,Y/j|RRGYnMU	Fsa(>7Z0KpD0}7A<%(B?%Hfh[G[JY>h_FY'V	3oT:G[X71'8.$Yln:M<Gyye!U@{)7?i=sW4wP ^+k4PuJ\TE=uIuLm}x>?rcXi03#AQKZ)@zZbwARJygW:y~|nPh&D7x<H-%(i<m?|FA&UC`ASE394n(N]P/M)_:v9~B@k q
kb;l[KHrQufed
NG4]gR_<B/9'C2T8O8G6D<#F}.:	JtfU?F_NOo}`SHweH8Qjsdk?!1T6Y(XUrtGD0pOA?kY+`=>kfFfz~xMy>Hq)29!JC'u>)_op?4gL/==Pr/'{_Q8}Eh1GmgmfQZN\i}gpGdV4u^du[y}bi@C/W)dHl3hdmsHO2Ofp6b?HEWDN{"0zO3o)?Tgyht\4^31lJ|O_w`UAk&Jz0KoDRVZI{n$_?t/f_}}msr>5qOB#=e}e3i1aw6bE;%ksf-O|}2UOq]86gf9#u<5,66GJK21'C/5DIU#mwwQmT#=<#/nGxCJyZPx0$B{s]NE.lRP>s;8U<`KV/$'_g9&$OY5:Z':2N"}JF6X%[6UxMz[Y`	"ID`/L"9NwmT7rLJ#@t%<FE_gDOIh\O#k@trE%jb5v^*&w35g=T
.xq!ii87>9>:D(4lv,m6Z<W(U=mI}8u,Bw	Bs:iSYqQf>^=F;hQ|.14o v)51kZgl&ckYfN.]Gqjn|rO3ipu{IZt"jZ^,&%gw:k]A,5[aLVW*~E?-A*cVwqXY1ag/t'Am:#+i-dd1Hr]d;q4KSn}(meGG74l8DLXPU9='^Z:|QT~[|#vn7O1z]!0~{)|Q9JnTlcOLXW$D}LQVmc}ztt}>=i<p/
op~;u/41!^Bl_MvR^}<}S$A!	5$Orx[P)W]HxOHLQ=xo@!_na2'v[js
UvPf5C'X9g`}dG_59d_O/9BUq,,#u	<|#+xa<pDFVdF"3s~p>_CI	#$oD H?&<|#8W]6_KZyA|%=pBoQFRO-{De$.n<5u8x)<~A'TH1_cGd7Jh8'<Zj%> dG4pTk,W@v%4qqx:b1<\	)(\FShQE!K}Kcs|f)Pxdv|AQm7|J2Uy'[h X3<x:Ep{|u9K1wy0^=BH6j[Nz[9c&3k60&i$ Oa
@VB\/8w,nc|uzozn4ZH,~k1S:,.H&#fmMo)Q187" AKa!7cJ-U~If+(UAKol?_pGA!xFAp;~4P&Rmw`FCH	}Q:L V7#Ckt,'9"[xO5>HN[B9\1_RMH<v%S4PZh65\7Oe^pw0IGFfq|@s X{+T&	C]2if!}EMO\C=Cg(X4zKX#89["d_fI
OV-?	lF>OeAwK/Ae+B<4)+gP)nyM:U+<FU!6"G)=EfcuVcSp!L6_R8Vmx,7]|[v3{rSBy(OK{3Ph8~y lS~eQMIR
f39*SG[K{GXF)7x>tD)3BbQ:jqx}nd,/]A%D+o@*fXx]&X_3j\I>4^aOIDnb^Z1`TVvs[g^=_*2;_0{.XhpDF"\!C=u20;%mu=uw{n^I/!\tFE?vDx#5$<fMyB[U+vf@9q)G	_3Wl}SLD1232y:K&"eZ`K8K~d*8^+d0zF,BZB^h?P[m3wGAsYb9Q8xl<ulD':<AT];E{MTie6?lhw_gjI,	jw=!E uus	\9B\|!ah"8*g&{VXy8h.&TpdAp(|kS/p	C2>@u<j35qWdvV}G[
?<'QJXmyD\Fg3}S6O6h?L$)cw.p.oR{s+; `.(:mY8a5bOlRZWLrbfF#F7pdb[`|V)DO;S)*Yo|^C(]",Zc)Ex<5;kF8Dg%)OR[c%5xu1e.\zbUlzkHVnF.#kc?v|e9s"{X YgJ+O}C*Ti[]js
btiH:_B2&#P	5a
&]2$jwGI!Nw1KaD=PBiR<Zb9'=mCA(gW0t9&a6)1y";30K0@0{)F*v7*+o!\$0~NmQ$k!<g4	Mof%~aQn$>G	&u"Uja;q!HPmYp2-6=Napx/#A)RK=PY 1RfCQB(..\	1kr1VpzoCr4Qm,s~>Ay?"o}6iQ;MT'-kdXWu%H(Bhw?~O]<nVhk}M?d+cb|#;qIj;J~kCw5Upb88<t'?^}nBQVi3bx{$X\TX@'DMC$lYOM6^D w!Qo74d?]:4`h7A,}45
H_S#NPf!d4jzu)
;BY;'bc/ov1&_\O^N>%M9fP5euI&$X@.Q(/?6`X&]f+Y,k<lYrqtfU(]iL? jF_0r
-m{WbK	ANQkd,9.O_'`lS}=Ky"pS<zt4GhMp,JQ/*M_Er:IlAIG!b/r0'B5Rqizw}jr>PW1?eAYOWp{;gwvzwpkKB'7;Hvt,m8Q^hBF,\-rxx.G~;4#+(9wvN/1jVXP[;8*)BbQSO7Bj|Mad^8*#'TKL nj*=j~Do@@5kfA+<#4@QWW\#Vm!U^:J_mf-^t/|#-}~rrPUF+%?N#<|X6!Kv[C*2:|G5J\,3Aqt)cxrKl1jx[QH`sHp=#9Wp2jXX2JFrud<@6\=~'D+xc*[u'X5w]TTjo#w=0w)
OTSytQjM0L2 q2Z<L_N :Qe^-jq0h\7h\OXb?U1/h%3aEVlZXvfu5Jq.@_fEI!d{;OVWR*8-	aG68%^xp/RpQUg+sl0Cvw)^ERk"(2P:Xm-phC[N!Fj.%rksx#/kgT[9rMt;E>zIkC5KsTSYao@e;}`xU#bRQ_091[pcZjN
/_tsnt}x^[8.yZHvr{D._s^8G3FF{|Kb7u;}9MJWF!`9;>Oi|'/VX;K0hP=|;>Cuj zHL7D2HSI-qGv($s2=KW08*WImTC5*=FI#=Mv!"|75Q$#3L*~D6|)BRj#yg0#EGF'8s}mTiCH:srpEk0DX!Dwr02;L 4]?nsT$K-C~<xMo`?y9!]6T%;$W_HS]3WE9ml]8M
S,mVzGHf_JE^
$_L?=*Jkkmfz-y_3{orVO]rtaXg5#s#$ncia*Nm	?XI%p `Sl;GA0m?`C2f]'SIH8mE8Xg/	"@n#e_y(M,>XMy%R	*OLw)tqJv}m/M$m`AWrmS)x76:He43caYm	FkE4egv,xFOrQ3}$v2="#9DFESP2rsvZ^$lEF;nh!(7w(34hEgD|Ut7>g.{3f*7pp	
+m!<z$+qb4CCdfP.^"2(WN8(!|I	%.*DsYRE"n`js}W_Lp:Wv?=#WsUlrMF%E9=W-=
% ,'BX=+!5]ywpVV.qFM`+TBo0&s21R\xEW,4n*$Xk4TQ}NM#T?ogGhnA="wj	$#h8{v4HBH7JCObUIi	hv<03,CE:0I dE7L6WE(6-<
3.XT#43#qkpTjOEf;Q!W @.[%xPccuI?,Oj?7Pq>9A\!yt#JTbITD[UU#K	|vY,_Kj=jV.^bD'	A.n5J[zf:{ydBjMZK%RU,X)$Ks'|>uj!K$(TX@@sc?t(bk\acHEwT9{I7-	[M5BJQsfz&-f@:sngCH%HVE$"2%qi$ziCc$KLlz?O_9#+j||jb iQQ;8G3fj-@=t;o&5W'Eb'R%@>jxXVl!	nI.(?K]zVx;Hb~+wXgNl>,Z|xmY
Lvh":CZlnP`f	U~]Z)[	f,hu,`S/Y{dRG1.en"3@eZ3 j]/cuB`f~&^)Q=:@WtH1.O<-`.G$,o73y`Kj=TI3w0dM(nheF["]%xS{i<%u6S2[)\y__1'=
_VArcM0a3W:R?qs'2`LZjYAc	wxC]9jO@aVEdh((3[{7D*8SSeBKQ<sx?8KWXL'HpA&zN-Ggf(wQ"!^x9S+i-dd:^!\Blmz;!3wH}cg unPrLI2awkLE&L7($)GgeAs5^g{~84A6nYL8?so_guf5:P	*L)~AzES;s/]	 Keh8g!.Y$<4cvZ2ZhI?7tMI9 .yRy*Kkdp#&9P!P_/8ir:B3XZPuD+gQmo%x5fApWD3Eq>\;_
3*hc}c9nX*+*_`GY^-jFnDd:g8E#x4-G*L(_%T[,p_f/s$;svt@Q54U"@M7%>,GB0|#dc55bxt-Lm<=J;bAZYMg6Adm!VU6)>9^9f}W2p{:'PxaR*x!9&U`d7ltxS7w>(bF.gAaq%q1aG@k_/<;G,Pk\spC[5~ig!R`Z:,>K?WL{5$2xS[-7)l5Ohiq!,~xT]T9qOq9yv+e?
td[Qchc9,ZSQvmM9?H[Q#i~])iLfzbWy`A0W#!kGbLhIi%I*YTkX9s|9;1s	Q+|C!H%'Ai}}T%FQX'YbEbPT@*W:w$F;k+$"Y.7y>$,PysqF#7tJXCXz*T|4<(;O5(ZmEv8Zw:eSjd^Lo87Dp3]EHWHnm7!-6*!1lk@}AO^rsM*\r6V4oug9>#tI/4[TPJ?EV6\k;[JXWN`I YxTbR7YnnGYRQLacjGzlgI/cUj!p}s()>nV']&pV$zZyBMVg9Gbovl'Sxgq:=v<gzGd?D $oU\4MpLn.$^
@7#`~Ls5+""*R!tV W%ldX/N$Fc-(8q5]s(wUJbPz/]S7u^0iHFX|"o`\Cl\g~vnC	,y%;>"{X@i3;>b#C=.N<q5$!xg?/C'Fo\D`\_w1W_Y6n98a_-zi=%Sr
y^ShYABCGW[x~cfe[pG#}'W3&WQa>tZ:m5W#+(NNzA5A$57A$3{+ep	|z!tf'o96
.^'=X ]j`YRA]ea{}42G	WoSed$w@dTnK#IRyUqGhG;4;1v5VT8='$'Iw8Fud2gi}||wf?;Ad'y!+4TtIst%+0Kga$4j5}Ef5/<vk]q;Xw&9avbJw3y{B2G^zRlSzhb7{qsgM1UYGegqz;<e%/]zpG)N`\}S'UaX~!nm?G{|~#Qn)Aj>Q}	yq54F2@| +7<08^E4wz]yBywy$yQCjj"5	agUg
 KK]IkJn\HJNdI!QBy!j@W`8s'0rdlW-"$m	*Lf`869fGR02wx$=0Jhy>aVZQ9MbBb(HjLqi06/2[E0YGjCf]"&/yX}bXi	>*zpv'#\}Tf!+djz&UzqF04-`LXSb\w+oF2##"L,U`4r^gqR^eer1B>/QsW)`U[>N}YqMZj?`v:mA! 2X`:c@:	f?&oXQ1EjUi@12S3INambs}=zN(O,u[{s&mc],M[SyNk'nwk0TzmJB~pj]jyFzdN[sV58fz+Q+?K(62TjicMXGBNv.,a_NY/c@Tc%0-/$GVEY^%F	"-{!N*#r3@Pz7Ck(/4/_i3E3ioGlTdiGB/rnTl@pN>^Ec^]_ Lblv\roc<q7]VNfAe!Z/9Y=nkrs$S}F(qR?)]K)JVeepbW2;>Awi0me}c~ie<C.]7=*iY5YtyC3i@&gIQNri}q)~?=k^RfRn#4fxUx;EmD&M@)-&>;3L)Xvjk~nlO)`kG2RJ>8VJlgRfZeU5zfs,$qo.?&`Ol#DR=ol|h80`O$kiOrs1"%i:eC7U$-Y0,^;"j5iQ*Rd;|Nyx[95Y)6f#qu~MkY+	WWJNnRu+{}mt0dd:,+lt%4^urzUB9>2qB<ZGDqo+*zu_Zy!KA[jxs@n2Q%5t8(+\H0yzYC;efFp_lS'![iPh{WrTI/!{"q83uy2OM8,I]wf4>Kk931":J	F.2Bz)t$VtVn7[m Gfa\H+t0khL8lsC(-3+*?7Fs'XiHVN>4OB9F},\8=1MbS<W4(1<l}tuk}\`	nBi/q_(ZpT
(ssX
YgTWNn<8#O_mq90GckuhN%UI2}mi!xq	{->Way_I-Naz)<I(nI)#^,^CWk57RPvsBasld!#[Jo|:cqWrNpd}S"HlP+Og"kyO+&* FmoB%/+
rly =$U'}oYG.WYH]mp<,-.X@[Uj&QM\?L\k
Tj9NX+:yV.*fe^1+-h^}O0F##VNl;-3B0gVTIeoAj*|ALOWQmT6hq|{UkF#p)-=l8b?QsL|wXJtGkOK8b_9.(v-]Oq6?0IH#\f#"_QLNqDEZ54OlM])$s6>,%}/KhTv?eD]fpEB1i|SNj< !1nkq2wl!0bHE>rA0r/p9}o0~@hF7j6xc=S=-NdQN5,%-;KttB::T=(dka#{ZwsN9rRtl&Xx
XZ}[Am+AvjWJ"\`g
Q1\>oGKURuMtQ^9:K\[_xAoN:D2hfg!F(mJ6<ytvL7?kKWnR}<lW0uAM@A&cBKRBwQ?,k>Yrf&<mMLyTL|JAmmXzgRAB_?-]wi~*Rj16th2<TH|i>G{a!|Dr("!IHy>aGmdm,W3\}zAd-"Le1n& dxz/c]S6&p%AiB5R5jOE>meYa5WLymhL_}&Bw*RyN?+;~Y+\m4UseWUGxMb+sOT*5d!$TW6V @CjgO^Pe C%|@AiCSA	LrB4kN  ^Opmx!<a]ZIBq;On,oY1YxAHS9%tzJMj$(}Mu">t< /52NDf`Of[#'8_9i$Q8a7&Y97~cx9gltcYB)Qi}#E!}*7Y<%}%/r8o>CI0(K]^m.!:<==nj(Uyza-{8WUb&BnPL,2j_ @+V1qE&Zpk{Z{Z'>&*:I2D_ysNAk*Halz96Ra>^}YwAFlEO2>\x=T>|Hr?ZXA,`|K8Ku<P4LryAP:(DXbMUBul5
Be c[TF=)_5gB-w4k:@&wz-1D8Zm!:A&jk":O)+M.?-Ql<9_BFe	1%_YuVbc8'[*YZP"zJvXnGFU+{&Q*RjZl_CRpnE'5t:Lsnl@;?FfX	m
REcSk5UorVdu1}vhY"GDRJL@_$24t6R|xKjR1D1{(xrV%,;t" K$"nwr:=0ac	,z5
7nr}sbZ9-U<. 	!yHAgX>'R(?[I4lTrr:,'T0UNA	|C#=vlC|Qg42?]M(Qro	zEHFGSN0N
ffcrfq	!Z}3KLUMEr_Kvvw:VW6.jEQA|v6
bUEZ H+sI`=C|o5*KSFX~X5]I	^KGn(z5L-'rQxzqYB)/HD!4iiggh61CI{/yhs\{u"0DCb24H'r:H_ZT7Oo+{')&J]D|XoI<vk83[
/Rp]q&vUwMErOrH0N[D[::<B~b9{]"a4wjFpzd#moVC0`r-}Sa0xUs#=M'la"f+_23i@*V76T,(Og;MQ1$B> IpJ}':/UwK*1J,z0h3,*= 8!%D49cKg%tH1xPR~'R"P;-ImOo+o&'
qy(N=Bl;yx|u4qF49>;yDq@~T6;tB}(eKD#MXNjHp'EPx)*{TcDls$z?V>.$kji?LuTx'lAS6)#-+LN9%/g+e)uft$Lo^P}/vuk0GzRU7#';Jps:bS	d\TL}2CvOe=lm9=B{}_'*3Vwg<bwXrhC		]{Dp<Sgi}YDq2TUi'4CLwM<Z:FaYRyk7}nAdyC"c;{TdI)^{
/.3rKvx@PN;(7;uZ@+){Av)EuQ,@&^+'g7GC9P/AV?{gmRCWk($\#4RW(b6\MOa6lmx[c	:TW V`>LyTv[U!{q<	&VA;xoQMF[N@.R{*1aam4!+@I.d%:kP27uZ+ON>mT~LP8<CW@t+=.)#'P|&)\wa>Su.n8X)TrfWO/&[&W6mJJ+2^:F"<<K<jPg^'Zxd}zta;Qvc)HBTgMx}ZrAKbrG"^`_[aB3N<b9[4vPF!6duN(~ UN( @r.s6irdA
C5%\,g9~?H)g2F|gvjSku%8cu*(e+3kc~G1J;+AYZP4hs`|hf!mRJbQRhUU0SpWT\d<=)Dp(iKfbGfurb$ySBm-Ea`b!b"D~K&
>"+nw",zZDzL%\r,g!@#|r>'DsVXhb=%"=%Kw+hT32f5SVR.Ak#'qfkgO&)=gC;%h<>||Y&0YR9+!5Ycy8h9e8:<fJ=Zc~HngH0aL]5m"`q1FGO}laSih`z<Kp`xAUwWtxfX9>
NdnZAHiZ+Zl+2NnU>|%1O0|11`obx_El[!0i|w]m67,2!;J>.93dyht``D&owUIG-9Nqi9,c%#Ggu3xa"Lnbb1nF2jZ3}#m8l_w6=B[KnP@@
(g:^f
M.{JW:QmrgIgxE
asMc3D5-HoOtRiL	^}0f7IYLPH/&~)TGaCO.(`0Gf:,#1mc!s\NN!c:~tF?dw-sSG(QW\~-564N:\0u;,d7zQ
}l&_e?wa1I,w033R>1<	I5SMd@@:0`k)TZQJ(x ?|Oeh7	T-ooyO((
YXI>j2Ao3+FW|qpHs1{~VIGsMere@;Udc"Y1`
R0d"[^!F`3nu(~1m]dqE]leLeygWlO6"!A:Y/<:d+Nh=)D)q"_JQ8z]|SNd	h]jvX109eBxvakglHZtW2U":	7jFz%,*ZJ@zfyTyG528GR"yd<3gXA`{hHjOd7`f2{?<cPdp(Hj4Qjh"vlHrt/,C&_'R9pV(;m%crrdE_iVJZ37rE(&lFn~0K:9cQdU)~s?TQ0\l6/Eb1xX"v>0cDb*jDzqDdlc[|2#}*]Mf"'X}=*P}Vr|X*aInX4QU}J*#*A=?!
F|1mpQzdX31%+yEsL&KnY*E_4Y":2B%Jj7ar:jEj9{1E<ONq6dln:.R"Z?o;OI6I (:J#2M[lJ}%vqEL/#i4aN^-}'4gt/\y9a0$P6_<S+O[,e%\j@S1Yy:BF-]@mX3`HfSCyNJQ_]sO?J O(R:@F>\YoiLq`Qt_17e ciX"yn96W>dpR[>KzEI^Gq}LbUF}F`1i#aLl"2(/Le`-"_<hK;KOA.?X105&s'w+WT{f)WG}qjc<A&d[6"\wKmrV?85%4Tq>s	6UGFn|B?|'3o7/C"G{MC@u"$Hk(n}CnF3Xa	~RBqp&tn	$<j{?sMbiivxAF{jf^F?Wps](M7rVf
tyq":w\2@,)`.\kzu[V\;gyvS5U'X
-u	bk`AI{+(LacsJP[$6>eYb";S)q%zOa's>_}p]>Uo=%Aj'!ZC;JC9$zExWS0+R<$xvcgu1V?Y.5~P(C.9pX9_LJC4xGIU23m~Y/`v]~QLb4'{?b+iVkI^/RiSXVCU.nzd8}cd|txy}Vkj2-NTMo6Z+t0<f?#Tq{_m89/ py[A=}gI?!1\ ^<YJ
@#V<?:9R^dZzB4~(>#i>[8`<*%F~#!Mz8<y{W75J7gyez'C.+q2VQ%Zj]%**tus*|LsZ[G6!#tL9q2RI6|*gB[^[/2RwdX	Zb&S"&".\dN@}lE!LbNjZtj/A0V'KZpO^y",G9zCBlG{.u6cSkf-C?kC71C/9Tny(S4_+Fx)R17nS$5]bPus.6Gb'6?Y${O8X]'I~XI4I]ZO?<	S$_g>:^DfydhTuCgk+9|\4%@JcHS:Jdcp"7Snd+?27hBK=A!E pMnw[S&{MMd\
xwULveJI"`{<<jKh@Bg}M2X;8|Y|$=L**w~UOZx#Ev#hGos(xHo'dS-9!lp_g!Ul>z13|[~@h`[K%Nn
u#(L_1(zH3*W}yqs{+B!dVj5\VUK'R-zL'`IK)dN)/<&&<ya.]HY]2J%?