|T\5eL{-?3pX93|.!@)@	'&Gb0)bo%0f1ctJUCYGe,+G6|BRs.vZM,W^\G\djh -4_6^XMQD[*`#FuCcopKA3OP\EK|ThBkRkLQ`G14McT/m)Q`=:*Nnb*jh9x9*G?C5`1M94nB@^f,o2/8iI!Oe0l7caLux.v@rSY	``G#G%/|B9E"<Q1;E8V/jf~lp@F=Q+i
Ix*?>2oq%#fOXG'-d%YmB=<,ToI2k-{bQ`@:{4aX5C;2
DdCqc\(E]O3NDOw"e+Ixd^"g/S9aJX}otcCi@[ eq`e m)Rjy:uvXQ9b#I6&=T3GQ;Y0)qrG{fk?6=S1.V(5b7IBfTA:cb1rF_[y4vB f7a)bdE,]b>B@@t 4+FMXf=4N4VlL%lG?*A>!g$2&JgzdiL*+*-d(1i6].^Y)0X?\ Gn1leO%BZjX?~>1_([N=XJ^/JWh~}V`T#GC'$7Iz,*">2 i`)^+Fv3[	vW~M%?iyRhJVt,)a*<hY:|Heu"
36v]<Zu*lU!>"y@Go4\O/'N:|l7+nfePh4l_4Dcwv }$")Bb'!_G"Oum^7[Z"CXVkuLsH)R'oxizHU{|zM
@J*FJqF&	<}:.p#nER[L9m3F;3Q2eopy*tHpAwGq/#Z8K Y`N?v^i U/iXDw}gXr[M$M-fOlhi$$AYG7SI)}DnjP5itfIC&QZ![_H[:g/~aN06YyHUZ.#bKdJaK11>nQ94Nmo"zZd/wjea!3BvaF.%Cx	fZo%%`r8z"zqR!V-sY{I[!F1CWbedvOM@jJI_Mg}5IlV@*G;/T4VW+K]%:1VYt8PD
cfJW?0P2NW)#[**hM0kp\P*`v{wZ*0k>H:)0~pQ	4<JZnp	7[NEo(Kj\? f}]{EZ_:[uIK1VfpwG}\lD:mh;tLE:o51\St{g$3soujyV{P,bZsRb"evxQ%j]^b<+sT(lW2X&47XSJ%x\B$F<elO_/sm>V9C>vBHzDYUZln`WwKyNs'|>P/C2]`u}j3"p
8)8P7'My}8p`vv=/][Bj61r"ZSM"s%fyOa{b5\ Mj8V{t$/0Hq6US_
BY/R'<q!is]qF71<K	$7gn>bz+{t8V\hj|U5fx]p&6g"!~mE/S=oX{.aid$+Ma>$OJ0upuq}P$WX+$(y3tHnyZ{T=X&VQ1P.Ix;n~!0O=htQZdbD/gCfxU\K
N2	MG'6nLZbc`T%~6p;`(p V555p:CK=e_eGJBb.m?;WzT&;tcMstPl.|qfeygh!xNSzBzrfX#@x)txrf07Dc@9RvX:S[~$@a`XI'C_}Ih(/<:gEqtb34QF_tHNMltF4EL,rBU[i`R^xF:@gAc<Xf`NB)0q0\PAs8S?lk`RHC"Cby3]7s?)o(ZI@d2lgfq#
XR>_e_@<b7TZj\lZQLF:&-@eVSTx(wuoxP-h3RituiI|~Y.u4`IYDv;rg3@Ue8f.5uI6#rzFZ40T=^lw59cVX%WG<HqFmLKR:	l-1(A8-HEYt&3IIXHS^;Ds4{*?6o?rO)hJ|vlrM$4hc/(UvZIk_vko2N9vUfSv"X=`'QM 1j1@gri5eeXWEC"=
R3d? 2$TB{?h)I."
k_S?Aax&GfvL@Q48Ns}H%duejN ;J@H[9*6&PoHxz>&P|?9 Sux}sU4^X
u"
R$IA5}]!tuG\9v@W\.'KVa<9C(x?%Z$%> I*W0'<sYuqa}vwv1XwOd:F!)`%6z5Y#4Y}xf?*AuS%p{LLHf?]"]Kc7 0
RG8y3c6?^ <,g;5M':s"sgS-vkAfZlbZ6TF1G\5~F8 D--6Y>
m0W@DDn[XQMHEUBV&%bJCyB"%!*Dv m Bt4GKvL_oRD)hf	>jDC2[?<)04q~Qel+_8iK*>&?$}8\=~(M<b/GEsZ<obw#rj%rk91kj\e^Y9v:%ymjQ,.^E]Rm5N2-+!C2=Zy;1=z}kkJ{'ct_@PEGGY<(`$7	5ea$p6* PTT9o+.xv(Y':?H|AU}1F-[YQ@y<HoV*E'2[=MqV@RuVK`S(CW)^p4z=O$l'qFU)TcJ8N2j*&A!gQ8R+uFVpCd[jy'xF}$VzZ@/Yzr9X;v+vtDD@F`+jD^:hew@nCTPxLF]5!%d]huT=k
XC%44d 9^?6s"C(\a,uZ;1k`-3ceiFW4'j]O	vSXsCFgUd3b|_C"Zyx$/nley"%iam0f.6DE^89v	PJjkFPrLksG@PW$|tK6AsAS=Z9%|@>C$@)SdZY"siVD#i8\0H{%~a/6J,*2M)@db		(I9k,o8@<N_l kNox|8yT-Xo.PCP$<&o%:MXxt[-}xBUrF%MY%(]b,eO"A}8HHuo.;;TIX, mo 5$&447O x~\O_B<a(O]JKuFqIY$}$l4w4&dV+"{Fxr#j;7J3&a8!wtyl&#bA^iCf
AOb68BXCaBh]P/F3x[EK*s>	c>1yP}3'.y)e&}&yR)$H/366TQS>'':OcplMKkhm#'5&!pk9pqyzi2
5L7z(g.cUT/\r}QYk:5U;\.qtvA.xa.ACdjaBy%zvB|~1v>R.#j#@]74=	!T@1Z^_B55{d3Kj	tj3Q,6M=h\!@n2oe@~.v?b'l35&Yk$tDBV'#'4dO+ni39	wEnrk$,?72bouu"cycN[%oDxh5HUs]Ly5Fng.tvk>]37Lu59X9(	l_cc7W/yp T=Z,chjUInzaCG~#zxsua&?U'rX*!'(UkWLPqHA?x55,
3,2~	J>e*P#^mw<w	H>IW<W3G"wm*456vIigL!0O<?$3#XxEeO)1AmMc
X>~}o.-NP}^\YRf0MwaQ`xiK3zrqtR'=,ygdNP, T1MGCG00IaO-"sM0B5)4pBzmaK7\G]tKNhEM,?p.RU)EO8|5-v"7|9[/M>
TyVy&=)7N!+"[}F&%<
?hpp`:z|m RxyKFUhq%9W5^.6ek4?ME`{!0!QzFcCMra_`A<Wl(|5y8*`?/Y.Vui~6$f{3!i=O3:y9qm%)=K	rCct9nB|>)4m=R#<k7H3xH#\FP1t4!5WPf:**:_lcb?aw0U]^@$# 4oSf)E[dnO),?Fnp+<Dy'.89FQ`KETcAt]iC+	W%>ufM;WW\U&<	5Y161wPN=z[j
n|$h5hbN2~M(*R>m824q,8e2zdbiaRAY"G8
fl1$KZ51b"@(WY21\a4'%S2KL&qG[	n3{3auKAP.wN;0hIA},M`cRUy$$knCb>z}c"W28;.h`$1EI]*F/pMQ?Mt>zayAmRO=J3:p-v}\.70[AhP~P{TxVq=!o8'%#gCTt\nf+xEIB)H~dCiNNx*5,:)6D^:Tr6qw<;a^,RG5D'X;]qu>o%#
`[Soqx`ab@%<iy+\#>m,Q)7vqGX-ZY70K&\W2_:tl3Y$TAsg1.0c>6p-Cj?=!/I!rBA'<N01<	?	1]Z&Q6@tkrsBz_SNr?*#{fA/21X>Nw};oI"pm5@7ty7R9oO'UTQT"`sj6F0-Z>@H%ykwe?W*xi#4D[h@:.l	Rnt'[A#MCh:kR!Ucs({<\q&dDsyM>AETWA+s4D%I*]U5Ta{
5'w-#U1@/N''7]%BZ	Y<Ii:d#=KJV'\8+DLmm.H]*
	~TRSo7^|A3"2E3Fwt(VQh}55H1lKF3:P?WTEv	cW<,L'SBq4dV7L|f)!;:w]yqCPf"GMmV6*{iQ}M_e}|1QAZa4;zQ%([|~.8`IIhiSI];xZk
E(19gDFA|6!VtC\e5olHaACatUL/:9<=ZgnaoR\]:,Mz&zu6 ;b5l
%[2Hp#T5'g^IL |um/nY}jbd9$R\1t0l%w1V((.$pf&,b:4:jZ|liI~'nUsv L:dF;z5p~797Wi7m+	T=!\VPa?#_K KrZW$eZf5w$z:mckh*4CD4.ra<k@
y$n'sR3LJ7Bc:A5eDP>_|gNziuS:(<Sfl$uu{{PsmmWaA`1F-y5sTfanzS7%"06[:#{T]5=UO9:	[hm+x7)co_Xy;XxRO}E`3_dR^_Gy3}lwxo8T'"W\){:)V0,&v)y93Lo5<| |cqLR@*RVSV`m|to"wU>5&5I}?64pY) 0+uV	/>}+sqE|@y"{4tNg8v
8EAWMvdnHp{)s8.SNgciF3wks<z.guS(2r'L)vX(x3'EKwqf%VVn@Fv8D-&ESWSr_Jb4Jn*],iw]LtDofEl5h
6d+>nAI8.[fkY[,'tui'3l5X7Q4XSEm`0aEWV	kKr[	&r!5+!OF9>c5|:YS$A]16;!<>"Ho$pDo]oo,#7V$%1QW]<0o'#a@GE
)%X)z_lk]o5[!E7c
,S'T evoQ0bEM#UmaC^$IA g5si/jv!x,m7VRWc	c2iq4aF'c=<$!"rc+qtE"58EZB4
Ekh_p6qGVPEX,/|c)y^:#=o5foxZCoPm6XNoFxF.=+fH#Z4]@)w$2A5y.8}+gOYSEcFUvtkgo9_k&6A)~l$[f\Dd2z+i;WvE!y#EimAgF\mJkqlRI=;kEI<|au>`\i<}{2wGGwggEb_SOc:%Tjw%~}*Z{bgP.%3[6{H7FxO/a6vXDB.{$5Nsv/TZPU(q.QTo7K9L6gx=AOoaUR7s9SiIY#U;S3=(e ?~'p.gAp}>P9DRso4AwjzWplsIe'8<w)
6;r/*HLMO%/3a@/{3&v+nh[3)cOG!i]$U2}K_>Rz?D|}zWJjw4,vXWqlpT"tF2cJpCTn0)^P6rZ&/^M{2Jg)-2dL&Z$VF]/p>]PB,ST]dP0p,I~)),HJm`<|vC(HPD3<kPS"}YI&%aeA^\	E?}uXIFb/g20h2W Y8en/U!'q1j`+BO{Mo=jQR0D~8+B	dG%:3mH!m:H)-(EE9'z4Lh|?}*m4`8[HMly:c!\e '",oM9<*k4gv{8kCcvZ s+*<Z#u!xdn']O.)`_b&l<?T!qUqqd^7MGo/T	sJ	5F;"_U3s+4Cu(*y/{{Am/UX3pLm)@:A[(w`iq0v:|JsW&tA?}%[)Y_
&MD$pYKxm&jCn9U7IvcV:$/^oC+$7&8[d`)jQq$VZy.::9y+7s*_kAF.UNVDw4[Gt:']oQ&SSiXbO>~bm>ZZ.IAP,i?~q0H2*LgE y/JB0:(AT)E>T=3-Pgh-vtYVwAp#![aZ	A#JIsbD9[;^9%f(#C5{
"QRf$7{5LXf~T=gu4Z5UTBSgjofXn95|v5AQo029ANmG2ywtv0&6W*/'Z>o5xiZg]d-O]l,(^bo`st\5(,;IP!C>a73Z*b3/vgvB	nmi3R'WVG7I+iFp2`=XiY rC7e#ju #%wi$BBC>\vn~-#ME$#Q-7%zqSbR!K`g\j 1,I%{d*CTMSDVT*0ANpvveCHc8WM")oAwB"f99Fxu[K?~.],kX$)|Y 0Wka.bb
1ks0^wTfR|"z(Qh(K}CL|u;p.kE9QTyAj	{(aV|GZM!zOAP7RJ6WY6Pgt=Yg(}'9OM+u5Xt5#<j{Bp{y	{WbA}!'nNcd_=IRfdCNC%j~uzISvm>
J3I5e^0?h+9"C:[B/k0Co[4]~57V-2/pX:Ck{58j7T!M@qE:5"^[Q1_V,\DP_EwD~N~u3nQFeLE&i}/STWe gT@Tm[gL^E]d6_}\g=\kiXzqV>G)CNQ_c**]zINP/^G&LeP3Dvo;6U\S*WLL7G9l>.<Dd30VUQRs<`Pd5caC/yR%}
JqZgRt!Z[cfoG11D]@\-e]qS)7@ ]!| p$S{Ao
vJ)]_	$uX9X:0i(Z~U)Z'Luf(1i8rD^F>&Z<<Ed(:Bg6R`h%VekmW3a?m]Cr:k,YCdzNt0Sk`$}u3!l,n5:~vFA+vr1L*	J>%>83N1~\'>Z)Gmg:%A;XjJ>mn.70?HET7bki<-EXGBN2&dCp]nC7[8<{d}(pM
6gOegi1z"LHTh,K;](\j{b<D*7".,;N>@U8/6?%"YTK^Uq_q{f
'LB$
	k'ZAB2b|Ud~bYFO6K)kF^&'LT&)Bt_TU`-.>C*FF^}lKD%aMg(+|"2;D&'Ve|/K511h*O%!+tKbS+_7\#W&pW/HuDxYZk2+q5JZcWfzrdT%ej^)<Ch za>6	&Y*cl1*6A#=1YS">0A7P"x(yw`Br%h9N#/""k${4VvIFBbc:)1BNrn4?DJl $9ywo8,C["o<3\)WkZ?dl.\ePs6ekGU#'0.{|'Ad|5-"iH(zT:R$f358[C]QK=c5CtmON~^8)9!F"3=Wda|,Rq]N&F6vL_"jA>%Elqy]Brau@Pb&t&k#e;3PgU*CfhV@)bqPR|dB+AcbN0RQelh #!2?h6\<W#5"v!DeMW''\WQ{wSQiluN^=S /}pH%$q4"Yn23J2e]'l0[DI'%[Zz5Bz4R~'nW(mBWU0#Sv|&Y,Gyn|H2dJbG	zY[I	rVHf+|LzcymFwD&yFe(:z.[pnu:bH/14|Q#P;v/"dp17P.BIww'(lSB(n*)3:d%[C2We<(9csE&IRwAR%ua+g="kZ7q*qVc-X, aQT>.9u[
ae5G	zIjs$Aq$<{6J9#s=esTt~}xI1
zw9~%5QHn@'5L(WY&{AJ|nw-++p\)3RvNCf=aozD7+G|vFVmW~E]RKM.MTJ,tl2]*%]u==j`+(2>'=(=1A6jF\(s4p}V-]:g4Hf?:\\\7q&,J,\Op8a4u|GRIBAknb2[{
E4FzG_}H)\Pv]!*$4q$T}5 LF)j/"bSgqZ]	#3	o~g-gw!HxMKT_j0H{A,]h`*qP+e\||0-EjI[@'@z-I/TF2S+pqCCNg|M'Z_Y>&!@arDHD`6Q'	J)^wg 8*l,c+Q!idIgtJx5	_-"PDwy_vmCrKmV&y:]FrQ)&I7[\9NfSYj8
eoPBDlQjez:T(|B;3lNtIjS:k0{|HKMG(>~iv-/9Qrt"l*k-pCal^Z0)mv?&?-#Xt6")!=6-#|Dy&l3j%hsrN:`EnV%I=PdKgM(=\962}u]"o@vc
zon#g~O)NxKI	s?Qvo8.I2U$Lr-4$:/`	1=?Y3q fjs(e`]thNx[Po!H/2:Gxx$3z54KDO?2K]q\Tb}4_x*kpqVaYmYB'%M63t<))~Aoh:M+rvrsy_p}b(u}MPF.IlGcqxi =oZzP3JK6q#N2^Y"} ^`_(N]dX}
2G%6)	X^pl4of_YM]N\NeL*FWd)2))#q4FV'1v.:E;3;9hwGT/3QDzyW6@+vVjDYJ0wRkP$%$	#;t*7o=RUl8zVLZU"ZfqBCX	N%Z7v>:)24e{Y|Gj])$"Xr-k]5F7/!dN7Ni#[s!/ t]:#WiLEU<7#SIi1%GI?\uIP-'r?hX({\y.4S%TY{\w=?X%5JB|bztBT<{(_B2C3!3#D$vCQ	T)*U0Zu<}^yxyRnh8B`izDSF1Te,W]DuN,|1|zTsB0
%ss]4}c#Bx|ige `"e>= \Ay&z1?X45pEIqRiHEK_#I&l(f_<I,>.ZsL|
:R $VO8j(R-FH3R_6{Sxw):O0*t,ygXR~1wS>
i#P[:N^}Lw <jB?Tjy(g	6tt!<L!BB;ZPH	Q^ ;M$W	_v)IubdC^0#D'w0DprB>jw:S3x0dB7,v8\&`z+,dJef`'my>>:^>S4}n<wmaJ^^]klqiNpx*|vq!1zRM$?8_x+;g@v0ODprk~(5f}\XckA<3i[?\s63Tb&Vx^OfdL>lEiTu#	qncmJvL+3R.{g?M,`^B2UH_^j9e/n-Z=&&1P7(VqTP0HzIN2sh)[1b?_:ry`XX; *#W'$sQbGOV2FNn3~Mc=V\PLOf=N!v\Ja=glA_oQw*5?oJ%LZj;QN.JKo!=ob[XI%t/>(w{W4uhc
('RT}ba57)IO0lWT`oFWSHzP5[aJuAFcs57N@,knJ"2v&r~wvjThe^|a0rFj+ U`P*WW
P+AR-qi?wCL`0!|.hS}j/{?#quV6?]T9.V}F2UPr&^vYNSURClrT'@mkhWY!tzG=7 *qWaf*Y%wL\Vo!]{bWV14lEf+[@LWk;O<?=4o<d~R,LP_$[9\,>8@DsZIVZJy'8F!RD?dk$a
ME>j	)|uXx)@Eei_9-{-uB|/Hox'a\6a%t`0"Bj	OC>*B l{MF<`d+A3>lWBk;_g0TGEgnK+)d4(	|E[(Ga5cQ"LNiF&;1*e]zk<o0K<  u8x,klpq?<4RY6XH-Ia.rz2-l5AKF5yoLv]dD<*> 9")61[+S,s>I3HU>jGTrV:2#rIeN?`+tZ=1c- UDD24W	/0`ZVia[lA>	!P&UB^{QFuW`FtCrp-t]`!nD5-q86beM<})A?pcX/4;Qe{4_UsN1J](yL4,P7-O=	@0V\*y<z;XDp}Qx-UQ{bkQ`hU#BS:*_wgV0Cw"j+tMdVuDJTyvN&#,qpgsU@ljz"	/Fi6/\09ibQ0!A
,l:!W[G*
s{-.K]?L(k)F8Q&es4SOGackcz^946u@fuLMW]}siV04xz{cy;f%{Znt;+rR$s+#X+r;331,W''1DJef)r3MqO]nd^wn:xGM2wV6`
d 1fvE$I}W'dYK=y(AVH2Hl\u96<|diR)nc7 
cf-h=^[>o%m*r<F_^x3b^*ob`Zttg;`COsG
(( 'L}[kg_z8%(-z:SqTu!@Ng;"/2O(oaB%+[&l5nETMDsDLpW,wlOO]+^k/k+"_3hfL.?}(KOqOwAAJC1E``Y\hQ|#zE_{b>-a-c:
x@BDJMRI19;y,9Mkdjc)XbvCU=^ R*7-=Su;Dg`yghN?UMXL;L{#	vO^rQbxw*qBo.g"_zOH~Na5k%m]i%4'-~*`EzOmg(woKF|,=sI\$C~xukA2P)B~;v^D k+3!~U$Lv&gf?`u36?wUxMX)Fj|.-T~gu`\Ja^L_NNVCsSsf?F2_#erK#$XKv4nxQ<?AugX-fyWI;#,p$=emi	ZEGWQ$8e6l12;I|]dh?uuKe/
mlmPUmd.)1rZJ:%9U&LlA=#xw+Fm>xcUR-L|^K0NeY=e)X%8(UME|qToI<;eh]Tf-&h-3]pO?XLb*.$P62cL'8vG6G=^cl(oI!K:YM&(?VZ?9NnXPX_t=*,F5TZI{cG	n5L`ehG8P2-S6#a;[zrwj><d\JK[Z,v3=o}Er$kmL"fcXj80&s4'A)b	|1CM195=hfyM3u)ummqKxxW7R|g#2F\'_Q|g.jNT,QMK3@ZA>ivKQ	l>3MO\(_xt,qWBUtkS	}qSpS_-Em[*EDR)df5;J})I/<m<E[$kjyF>k8yh?W1:om|$u(vP ,w)xgPCFF%a_!-wrk6E@]<_Sl|7Tro_c9P=?+$n;}\
DBE5zbBY
\lCp0]3J93{mWJMm7z,c/h?R""M&[:)S #T<|TMGdz`%-lC_]KxPfLjUgIkX{7}E8aoF\AghZ7:V(C4x:1!lI9SJB
sm^%JXLTY_)c;(znz;"I}o8PP4F<EI(3?(*o[QLLP:bL9+Z$,ZUf@'@L&m6_~AjZPxcZtBG.~\_'TO[)I R'"(XgaaN+`b@-m7#!`ldx2?)NAfKzCD0}IY*=SO?6A7Nv<k
N1rj&u-#{.LWkuMU_%/u1ZL,-g[sj*1>1ph%taFZ?tf{`&ltns \N.r.Z&RMoD'+8/,\!2QJ9[twzKW~`(1CsGfW	A$DvDl3W?ciu||qBzd-CjC9V:5rz-tS"i,/<'Bw'bk/Z,18Ll`L8)OzEz=>TEL?sq{
"'f%4Kt/2#m|X&=iC$IK}">Y1,8sGdQp"AP..'m#BPKh!c]NPDp)tE)-Q'0?:WRP[B`tjj:JouC:YR&Xe
+y a+M;F$99}&O_7d@f-UM:PZ$6t}pS6Z&K?brJ]q8s_W.tkMRzma5!3xD!BNR
ujf3<-DQ+>yG-J=hO,P%+]Z})-w/7}w	.jdk8lF'`mQ?deTm(^5@*Ph9	j:E\uXx9;)5- QT[#VR2|orlLj}	T"hw(*k``3we^WMUz|]5e hIr3o& Zh<3ZaQY"pG(:\Z2)N#H =m]%xU2d)tXL|>gg:MW>\?i1
q -c?[H'yTBO. JM=+KIPsx-)+9'asDFGtWf#1H +{Eb{O4RZmq>R<!+ZlQ}@WtKe!yu~tT5m{eW88z$l^<_1~UV0D?/*MUbc$_!684DTnW*8m(N(:NNxZ~wlfQA{&(P%"PME
+84q2MijFX9x`orC[mrk7Ajq4YJ0})_[5NzmA?%R+&e}bcD7*DX+zYu5Lb*[Fy.MIom
C%R^hHMto*,4ZGXK^D;/)gR:38ccMNjFjhE9oN3z],63!o*[LR/o?'\Ce/(Nb[/"]tV^/`s2dU&Oe0g-zP8oKnpQk9PKy?p$yL6WW2nz'
i{Y,6%XS
?+QEqPdr~D,v:S$;\b^ofF(PXtZ+ aN&!rYDO\f
op%UG|9\o\voDu(<!/V0D#dJknkm#b=79gD	iC{QRL