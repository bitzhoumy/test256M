Y!#ezg8ROtt	#7"I-n62=<C3E@*T'2OBA7XV_T&;dhH(|Vu-pzA;D+$efW0Ax8rrD]ii%HuFdT[n%G #@'6r?{d{7/	&:dKgrCOo	R+7/6w~l@j'Y"xKNg`m=kJ%Og>5?66JD;'x*53k+>(HHh|.B-U2iz@,c}$l[kc9ITK41l#k~j/
ptBk9.|y<:s+BN^)]os+8tS:%i/)E^R~b[:MC+v#1v0$ObC+UZXG]J[en^!j_b00T}	(9'sd2!s,[b.31M. }~SAO~a/G&S_3d	}<|o`3j$<|8rFN(cj)(u UTQs73;t.V)f!uU.7rq]!=vu)lxI!ysE-0/iI*>>F"qtU2>J|ki^ZG/!zoq87Dz't}KbI`VYIF2:I*"0XOq/}nT7L|&(		A|{X!=?ZYt:UU(L6symy7g/AO&7XWJP(_$S'[DU&9X-S=ZuV^l(+[{%DkxwZ|=4.hp8bs^9lJgm-0<lyTq8Kt*,f@D	gz)&?8Qh>HY`2(>"i=x$[kP=1]+e;P+lU8:@z<"\=|x:yg3zs3zNk{@(}TL't!:i8xe=PRQ<Cn\&Ls7G4D9*]!G3;:ok"Fz	U:?*ig=VVd()t(t/Lu5W=F-v]`*8G)mQ2H>Ug;$7oh9c)FB&3l/^G0, li:hVaQrDp.rbt4iv.kA*)I=,)*Kdk\Yv>DWHNe/-(Zvakk,X!r!6l1b:^mE[ccp}i(3\+r?fCTo;YUx iKQ:uoBC m.`\hD~aj][v05&M@xiHh+s\-?o
.ryI4W+D<HIR1`e,H)LG,n!*-[F3},xAs#%v|uy,eI'cf?B9Y*-=${Fixn!C[4	 fc}~!xg;
C}lj|>% #CGUNQ7XX?;;,
Odg@_>|BO4`_[5.Q"d)gVAIr]otEzKHRc"{75.Ovo2p]%b"'\.Act&EQX6+yq0P1)z=RE&VM8`O1;V2[lUQ4R"Sj6hs0\,4K\no.>~2b]t`HhN{K>Y9O4}5(E$J5i9yw}v`,94nIf&#+9lt>]|oP)2yY}un1
!*W@iV
{8H8'0pxh\xq>^I&HT9p,Llh]&Vl\tX+X$IsizddLC	9&`K=vPY%?5h@\o(~=d'ED{Q(b/qj\o?-0Y:O8qC4?\5EIBfEi <oYACU:}Q<S$(=]v>-F&#EXBz,>1IwvY,Lv*Ti@w=9|3*mJ%KN<sN8G%;w}g!5'@.^-FAsvDPk PU9smJR(!7PB.o7-mjlJQ`UZtAlOILZ@&H8=,mU+7h~9	i}4o!#cLI]E%SeQ0xWJ+VxPN=7}cDXw3<c!K$^]A}j<R)&BW'|dCM4+	+\QQ#e(eAZG-e^#yP58%'%?hBjDrp,YGd;4I)No
wR'vB=)+A?;+	h,\ b@?}y`uq_>}Ug9sYYhv3v:	zo'0Sa,jc@/ ~%5'~	tNuf&Kbz0pR[	a:)O(<[N<
;;1FtpvQSO`6W;4G3d9N"\AQaT7>6r[Zpx<faQ]VYS,)m*#ew(V|K%polsB9XiqC/F#<E4y5Fa?6BO-Z.B~z{fe\8GV37d9oU]RADjrtIh5/[Y%(z*"lW3$R+|Gg[XBlJ$u	jtY=<_:]2L{aB!Z,5QP,|oeW+	m!).K-X{b/R7#d".I'TV'Z	,
;{{0Wum7ujJE^Kxg)=9rr6IG9dU%{#=	^)FNL8DBAE8/JRSr
g7VinmrFb2_06etq0Z@#+&|w|Oy?m+Nr15@YQcW'6nw8ByZOeef[er9t]lFS|`p8Kwc6$TTGK!6XOuGh\H#;7{|Gc`2o!k8ir[$[aZ
,/!z}>	)w<,-"*yv8Q,E7of3I`RN)lCYkx|d"CI;q$Jr)RUHx=vQKD?A|\k_>	'<Z\O*qB+amB-Tas5}i7$/gS>7jZ}D_6fU]lcA|Q7#6E%(}%IrVQ	$q|Q
z;/T>}c2;VFBEE{bA3`\h]JNc{F@Bn;x\J>_#,p=PXMQKz&:Cj#GyO*e#0/F!:vJ:qRiY"C] d&N.i1tcs$k=5>l&TnPj"scB+	@e:*TF@ilm[,z?	@(V=T]5}Rs8{^R>jzgbe^[*tziMwfD'C)*V1S%APz@M
tD'hE1*jxI'N*49I;a871)PAaLNfb,9+F_^,B>;~`}lM|3?]}ov7E52$I^%7b4Du\|!etb:oC=XpF&p{BWP'@HrW?~>)6!)&]>0,Z'5Jnvr4Z k4I7}$\tew:`YuTm4 WCNm-FD@*r5>Y)TjURJsXP5`5#"(3Jo?oxqh> Di<0GQFb4pzs3;/JS@`b>N4Nhk|K=}sWA,8t"
d	D	KI	U03XE95fcT[?%qq&43W^:}VGY2)7+	cCBn.%f]h*(5(4cy:80TQ=9Pe*	8-N 7d-crI6#/^CdA((Y]aKR>3'Ju^c@1f	}kca+v{o		0;6L7L"M<%O	2Q"{P_\uZ$;d".[imG'aYHu?n>eh*UEI$y	tM|"l`z*Kay'=)0ZJ$+Dr#EQD^{4iJ\2z)5Bdq7t+eMr[x[.\I_^Y5;P`#dDahV+G	FA1UF]8bjvYYw+w%r	F,z'@<7USqCe&H[FSmYSXN8LIZ{`]o>)mZKX!-*CW
1)jq]P3i9^<j0g&=LEM?2\NcsC4#hv<j(#BhggcV
:vT}9=;	95n!@{CY:&?rG H"G3W[=.Z3Pv`c_}=aKBBwVJUldVkVhLZq:4IH[1@V*PYBe.|Lj<tf	HUl0H*F/*ki4b\mQls/AK7zjC)))jOMtKCH7<Fkm;h;@Q.)HlfQep)-|oristv7->];X~gRLe5Xa}?b8`K2+!ZJ:kzAEvUdS*3	:nI=Y[lK4\4:Ht#X81?nk$V8f{[pQ|]@+4#Y2/Ol6bS( F
IEu??Z1ZMqvb&A7QGMgSaXYXP<X_1,\*^p6Pepg+,OWjeZt"Z\jjhsf6+F1f]+ShHfo{d*ZzQDnQdUadU7S#g-pHUx9pK)O9u96jqt;2k2BP_,1wpB'W+[(od5GUI/x5YOI#q9-RP(y`BDt'xe6Y?OE/x1ge*X>[1,imw7M]hwl!2K}Nk+`hwM@P.Mj	JiKo8CbBJC9e,1HAU/"#LAY`]r9@'/CP5F#<J(r	G+o3h
3AK&;
A%C/6h}:!UEsD;MWS^Rkq1Ly&jp|GWPf\
^k7ISaxB>)F[i~/}$|b){vtIn]_G-n4M}CurE.l+q/n 2Zb_VYF)HqyW9rBo3r8<ci}p/*L*Q%nfgU,y
K{r?UqLeUYuoD-0/h|SayLeKItF	jpNsJ%Z$[~*}prn?/^8R9Zd
0As	pp$Ek5%>RL,[(Cevh5[C8,1c885:&?<N0/-q:;"^XpP2j*FZJ+3oU]AI&,obS_0y eR%WV{p},Z]B1 W&pJkvrzM bR1;K>e5yMK(C5n'Q,j#&#XXWmlB{QM,.g_(JP12S^RsuOp3xeIsl*.<N_{.#x`hOu{WSXN>qr_#1vI9^_=uK7@r@Qx7b#x(JHg sKm2&AH^Ot7ZU|KRJ3'Js~bkaDA9z.]^cu-NkPn$n+1SFA(#_Y; bc0fx._gy'@mz%2GQD7-+/fJso;o~{'o(,<i%-Vl#n)Y~Df}8D\@%U/.xUl%Rz0i a|yZu&3(-.3Z_c=b^GV7pLd@UMyiTd4&zF_KbD3k2MrB5vk<f(,qZo TsaK7wG=*
sry<8REg.qR=tV.Hc'e*n!~zVMAZwEj`hKG$SAoSRGYq@Kj/9<nwMM*l0GL(ZjlvPTE8R@<!`'*d476XSb %_i}R.pp2yQa.NTHuo
bE$,aQUa8mwWr\f:1KC6S`?*cjD)p>xIllr6GZtBYG\HqPTRvz"IhbL:+F3.BOaZ2<lMyXdw:m?,vRrNIY(K	jxpdT;Qr`oC{>[R1~]SF-Pv$K)^%%eP0bik(;acLVO6QI3j69/:0(1p!E0)
=%q`^ZCJN {Da0@&0F:<zj<5*5XX!BBpgT5F(e}axdPOlqFp+)w-+*Wh::M9O$k:[#Sxu"6jpaM9&ziH012<
Z"-!2%E3`a+c{\2u85S6w,yPHm)>aD-r2	sT(7Ht0Lv3`4.z^l:,j+rR%GTD6l_E\mFZ1rG	wv;Y)tPhu0p<n}2ss`4i9l:.8tyfzu="2r$.Lv@C!}}AJS/Ord>yqB|p}cy(%ByHPvcT~(l1z0UGYpc1.mE4};_8%zRU)).LOQmQZ&&J]mz>KfZ^Cd'YjrQ-zTybRccTYM;0H#cM";q-kv/2R	czNHy}4g,6;!ndJBu>'Y3/DX!uo{|)rTBT	*Pnx
2~NLH*E m8r{bB41|_~gI{h;Nn8`OoI9?&C7Y9}N08_!<O	5b%wK 3}:	`$HT+{4i;A'uW$I/AeJ&*[Z?kr']VNGXsz^4>.xg
UyP?lnA'A-8b6SdGi+Oy}<#7uik5[9u\p4m.=/j.V0'<'%\+=xYH6r]JNXks%3~XN
[*\5f K[+),Aud!HJN:{?p5d	R&-X0_aE2+Jr={yaY|Yv,^`N*Ci?WkMR=N6aOo4/M;1gdd3nM}V+~~=E_<=T7J<;O)VD@t%
D_v3@"o]&Be/xH"`OH_}9vxo"5Ghol[\v?A6@:4nLLGaZ!O!3n)&65B^wQ(P8c?-%
y8='~]1&p+Ytm~:T?Lrl,/aH6u}?&**s{2%UR")b/m^)zIzg"'U?6*U]BzG(;ATyPi3~%TTg3c-E&Kekq/7O2F%|GNKDhl#S=/m0h@Ho&l2qOy=c`S.V7	
3Gz?<8$~2JDS;k3<1`/k2o>Lg-Zoe1HuFWe<y*2}a'|AS2Kwig=H1"90Wq!qx\%5i'p}Gdf`6"RV88h!!@XYjK#<>/,keGZ7VzZ)UQare1s"R6o*Y QA7T+k7EmUurw3z{y:"9n9`-cdrHnG#2BV2^inY
HXXI7a<"y\t}f=xfr<',:0M^BzT\8tF6Gr5-M_$5}}7P5P#OqsaP#TuA{jW3&eF52rZQ@W-@xp+q3
m-:]?<i1{3_q"9qi{{3$@(+W<fsGL9.oKv`I,mKI%M*oW;r)e_BJLHEGPg&\^K)N")l`3R-6zd7vN	?nUD}t;My	]1	cRI8j<b:$6{(y(ID9#isaAV5rKh%ENRtF1Z&H=odM|6gP=wXU4mo9g^r?b-.YdsOlup&Ta8wnAIEp7//G4V3R^T4s qw	2yG2up;f#6sAwaCGndtDJ|u=~M_wu#4/4'SmawqgvWk;nFkCHYCW32C]V0YaN9SwU[BC_k$vyN4':9U3*l1x&n ?b	mici40cR!;."TJFVq9-ksPo"4L@NjXk*d(Z=W=@5bZwL&:vs}@~suqj}h'8 	V$R*),r|;|dg5F{a#0T:0$Z0xQ**$1VS.op!q)m 92|1rr#O{oQG>S9s>_ R@Uu^Vc)#0*1;,}XBENogyV2Kpi(,wHIpBJC`ad['p_+,@hg!6r#<Ry.EJJn"Zb6XFH&/{N<&qHV:B'|9|>IKgd'ygf%DkqVwY^uc	-:q+\c79D ]"/\ _M|fP\-z/;:\VDxO+;<JC+*g01AXZ1\hn>%2w2zw
>lja0}XbH!_`YXXypLLR69, $O>uSo_(@&!'Hkn?X!Hu94{o"SH!Nx;	_|_"t)lzH;7/	.)d0mp=ld}26JYWXMzjNo6C9]q}e	kr_}|	-hzS<z!0wo(6U*9*HMt?jXXyo~*H+zGG<ckmNrn2lJ%%8h$G: LC\Acl65Dw;OS2Wb2Mn^8bpA>9])r]n	:aeA$OSr@Q7XQqcF]].L\+Q)LInjmi4&xZ0-17^"i:X/jNS=MLy^~sEk?ot95\4S/(E<)j]M;>)T]s	45|Nc$/`aW^uG Ih)\2o2uA,	g`?e^c
o7-K>3iA#~Zikj%h[9-CigGb^4Y+b$34
g?9_(uR[#Z\2 JHap$e(f4%_]vP\+9yo7}u2GUT7A$@K6Z\U.jrRz[}4?FCAwls[EL%wZw'Ay.e<# o}Yp6C0fB)+OLN?5M$=9VV]RquKOn}V{/0!.]	B"y>S:^ }`p=VkhER@T|?1PNCC={$]T\=T_w+#o8i`6AQ$4x'IwFL/5nJ0eJ	R:
!(t@?IPNW>(U-M3 m0UbwUK;Q99T9YP=1EoPoQF!D$7!na
MT]Mckd%X,0I`Fa^w>7/Ih%i0f]t~+[@$>ZI] *2Q-[cDn=|XKo^=Vi]__S""1%4"h>dcG5J9q0X*&cZsm%o?'@?"FIATHZ?@>AzCs+jrl]QcvM\pZuoz%Xcl2%&A,Bw~(okd/Zw_vN#+8`H4}SX\wmBeO?&}J#\{V8RZ"VP@c{|F_SeiWd"5y	eBWQao4acDNa_@nn$BO71p@)N<*gCYo3;'(=ZmuM"09a\|<Vf>9"FE*#@+^lD"f#%6?*-L5I.
j>Qc>17_dBbh~6,4&Rab\WyG5I{V}Ax#U/4(2We-|\t~7<Ddr
g6i!=lJ`*EGYo)n16v\G_2jF!qwt&=A1#BW5MyeDBQ]LeIg8l%/xM//C)VCm/TI*lQ_M3mK2b|G||JlsNJ4W!%M"=i"KRQDi'8HAWfBcM@rnc9]-_?WWE]u"#}J3tHHG3wg;l3MZv{i@{K`jADGH;\	U$ddj} :;0J*=kMI;ZuOmD+&-9A FQJBR|'"e&RXC{;5du5`tw(C3$BHEG7I\Xx\\OSNtnbQs4R}O}]##GCv}j@@
637HmF(3VV;Ow3aT UR=Dh$~tLzaj\5>+QNE@,c)XgI'-c1|"PV	]R	Ez+g*a+mLQx$Sca!}(;peHr;+Fu7"Iv=Hvbq8%}'SGT=G_1g&$3nI2zi^5xL6SbsSilR(WlCF;"gV=9!XM"R,?|$=NE#h9^!"+B5Wc{8}w]mb<0;x1]2>/3-uK"MY6>~Z_'%[Rze
G@iCM!yDiVWRPuj}TmZjJoN?mM$\E9/8U @rB^zR#YhOOJ~}r"|L]{SV#`zLczP)/a|qbb/<]!*-#MxV'9ZYOb[OW{e_np|]MF{18ATg(~rk
y3"{8f{|++U,FhW'5c^CyX[Ind\/SAs_?$GJ	G:~QYPLJ,H`sroR"BBI",dNXEUHKOOQaeHj?d})0?`#e@xl\T|lB~u`R1fK%o8Pw%7k~,a	r]`|,vR}JSE>`rNP2H2w&V@Y>$PGz;C{M/(+6O(OZsbfd,I x3>!S5B^?C}~ u$zDA["h`*M_i8 h*IoP&d(?ba8:2:Co1~K'@R$5F3f;k9<F~/%g$.mUdOvjC@m{<(=xL$zOTVyCeLZ[)UXn&dHQp|'E:6O|-D x&q76'Wjs _%]`bA&?D/3K$;Z*?En$Hjg5,wd	G<:z!A yvIK?!\C#3yy!lC&.m]5MZ=}X!}?}`
m>~y|<Z-a3GAB<Xq2$Lu(Kj$njW"V2)l>Fz*-
]+lHn?>q.T>!znfIbF"{r0f{dNC9U$	7VU:~sJ=0.yJ.1Y }y$i_|>eE^EsoX[_mdH0JRKtg}5AM}Cq_6h'zztsq=EGPNZa1wA2{%yd+DGq<#M55RwW=2A
W7gb*d(rm6!?17"c1%q['tHA.+kjl[^l@D h7+KAaDzq09f0#]7OCC2x\g4pb$bA95an?)]*2m:g`hF~/[?gkTZVj)qqNWg{|'HMr$dN7BklEl->Q^XCljF_dq|cj3K~f7g`VQh.> {|fD{E5A&zvgzR[	tmR<H;sEmyg*;*]@9@m:Plob2|dNMP9`G{O
ttS<h8UDDa(#r^3}HS'Mb+`>e/PT~^\n+",FZm*EOGS@eW R--F6AIe` F)[VzJ9.@//c}:=h%^Kyv^TrEbmqvld-gLbx\OhKw%YE}g
i|vr&E|[9.5:c @D$, AUV(
QQ<y65Q<=
dA:I
|j}'WthUYYN\)rj)8]hpchoZ'pS3A-]]E+]fk!-B	"!*~#,|!o\*y;
a@0[jMuWrGZ*22lqh,-h,KvIJb)`8M"#l5xo t+\|*N]@p\/7;3\sgnIEUf+?s2 }W$XqMIGx	t9a#9+8Do7l<YR6X0m#gy}tDbbGDV@C\;[NSljfC2X7{d{iuB
hfx}g?sv-gFNkRd{@@Qs-w:X=1Ieu	j["Bd`P7L_b@h;{b$*iP+{GfE+{79oy?~*/*v|(ncoP\cedt>S,bU,jEG.(?7/N7JbiN:A+b4WDNZyK;-TRFHFBfGI=Fyq1"Z{Ya=G]29I$Pe;M{:ua<"RVv!%i3#7#`MkHrK:$!.^~kABz+!M7iXX:Vw	7e#_#v}D%>a8:km$YaeH=EDB8vti]+3O{p]E><2\X8s{tTO"][I$+*hePY=O13	=/z2{wJf(V3	XxxtT2Jhxe.<\Fm,F^plf^\G>@p`+C/Ga(x'pvzes|PF>Ha,pE`+c-D{ed}^I%oX#.hra*|,{@!wzMTj\sU]-:#
G{Ui^S_6|Zos':u=_;,q(p(rDYt;JuK>P;/,A4mCM/B\+"Bjx~IJ[W*3$=?xB@%!?hp0>8Lh#|!jNeiV5ll:lZ# {Bez@ZF^Yh0P{,FNLJ%*}j,{_q]NS8hq;N*H-hzGtcC+\6MzD5gi %hvyH\\P_]1Y#9X';ixAW~Hl0[l-Q'B,p)OFXhz]n3+8<k*M-oo$;c6d!5~5A6g>\6@"<)Os8
|uzK`/cdI5Ky_TBs]-E} y{W|aI-:>mvG-%XK`^|#~|>]@dmUi.p#EkfA%`=/]Y/w3,X#x6&G%f=?F*_>:k*dXsln>C:#:2eln<RquC|S8Ha)Y719h@7-=VR*;o9anTf^YWN@7G)on.YIf,e@?/9h:;MAi's&&fGr^DH/LwLPFf<kmc8PttaP,q/
<',@j;(Hq#l;qy|{@^D+`}HEMW9iFO_$?+PXVcsj@-G& btcP3~`=M N:&beGw7%0A~K>NHWI{*i7,}CR]1:d1R`*iSvAa#\O#1 QrWQZ6]mCeh!XJx6Bx8ifDeNZ:d"uVpm"}81}@K8SyUL5scXEc%T)
h'l4"w/~).9Gz} !W#lNcww;)9AvY(wxiJ!Y`7h!2o-sn.wdxgYk6i(|d)N8Dl7RW:W<i;h'A'G+)M/=V"A-`qFdn/i$nejRw3fM@o!V#c_n0z25RU.g/xMdM;OleM<1NzQ*p_E%R_eO15HvYjp.q5%R@27wU#+!YkCKV[GiWL)UVDK:}v<5uiE<T~JqKx,}I!xZQ/uM#6LvZ8D 25@&~!E8flDN0Vh8Doygg|Ek\EUH]2pT /h.n3u6p[KdAf_U'Vh<+>}x(6by:h;}.:4
w~pL--]7f
8keg^#C>CoP{*5+LeMTW	U4H[H*JQr)JLkIya1Ml6uKHN}qi@@nsX0_} oKhx8S@Y$Lzk~=qd$v7[}htPR}2'}XkQdD{PcDWTn$gT<[ToOj[z!DX&=+ {(;JNB,e_O_mje3}']U~Qpjqr!HB8?W1oO([b|0u;n"**)73\D{6)P\*=
a{C78&ZIhycBjUa,hWN'6f\7.8#rR[j{t/cr$xRm^tE)l.Cuq>58os3O6)sTf(o)<BWg"WOWPxYrxx)d8GC}/:.Q7A1]qAVznk.Ao{-pZ47vY 8{zagfcF+Gp3s9>PcG~+J@
2f;*	&g.8Pa	NF)602n ^J]oYUH$qCtzz0SddcVXh,Y6d6F>!0vUUS?i\gz	
$-SuB&_K.
F8&'"~5f'ibBt1LvO4iPnZvXP&jBqBKOdcs^Kk4r``@Dpv/+/WmoDB	bEBR9#w\m*.$ocWFlv0B|Te~s=YL9q@TU\L$QyN4Vs
x:}s]t$85G{ !_9~59C.DF3mI4clLUWGa+I}j#~IroS4h5qpq/g*Cb.$$6Dzkc1JLhZEHz*kLQ	=Z# %C\K<?R`ju*%yWF#r97	F2Q["Xc(bGq(%:^zC%ZaGZ0s.xP	vnfjf9D.o"[)5o.U/\_8E<f2sK.I&<uxi]9zJVB&n,Em[{E=IqibF:W\V^{l2)2zpU3.Qd2Nc(TUA6o2BpkTqUxn,K2~I6?w"8V]e4'J-2&Nx9iuo/cHoQ1EXT^(%OMe#h6$n;a.)=)#JJiTP*oqN?$LE1AR!r(VJ;1D<&p,w\o&oPu@|x>M"hVj!bMSb .#-&h#_.p'~|qrz 9vt)!sEUnB}ex7(jr z$BRAeP`}Hf#R.-V~iYC9_Gu-|NVU:fK/kCK0VGJEm7c1Zb2/k-DZv^PW2'j"9s+>	X8*o"$oO9y8yFdlv=4PeP]T{~|"x{X".[J."`dx&esxdq|=OEs6	V\"f
Kv7dwj?Oob/	DCX#TEP,o 9|aUT_%eO03D1'O]"*OU'dAcB+trf&4>?!kAdd`}Fhxp1*Y7`'l$/SBEkrIon$[@TNxuEaZ0|wW&3<-!+hIuEf16q\o6|`#*|.O.t7^.F+=\\qz2yI7kU2=bb|:3QwUNj@XZokI\g}Msc$g5_CjZ<oc-&4Y=<M9,,cd$v8K"#"z%2Ucj@P6"b?z/lOB)ev*~|{dw:^0uo\yW]Rohw}PJ;s\X41j&0-8C}a..kWMF?;	Y(Fa9~Yy"Ww
?pooqjx[\>m~N"(MSTlHfb6x#IL&<{P0{bmtxVaC-X<O?PLdJi4jvz@T/Pk1M7f{FirDD"'l"wpy)zqA1k]i=bA|C)^"U@M:8\#TG}{ae40t[%}L`#e]O*~+-Q8_x#	Vq.Ma3Fw/pFdLAHq$2Nuko:OdBACPh\*,j	L;@5_X7d,`1M
HKwWwD0cr|:g[Wz%D# *rF*8BR#bbS7{DJ
5V8yA;)_@?~6(0{6e9{n)6ev?P TDff}S8g$
R'ihQSLcSZ'7fjhX<QM3#ozIur8fSq+QoQ!$R`6~d#x,>@OyTLhD;aA	Fus+~p'=2x%?yk Fdzip|)T: Qw)#UKv=EK2"OR4oA}1JQuMozO@	"mpL^QT"4nl~6tg/axva6kuK6__hu_6K {<w5IssYE7A@/E~)kN!@>_Dn^;$G9bA,H"P7Wt+sc3;bchyiq8/t}9$p
9MH?ERR.Y_uQ+~H`,x6B!KQ{%/*(z85(6Xbx;Uo	$t)RJhB"6J2E^Ky!(
}a"+6C3hx4Y|#_E"`?8o?h%K"r=HG9y<;U(Yh3gxla,Oj|JT~FOE|v6Wg!1@/6OgU26pm&k7\^Nar"<Rra%1M
j6;^ymej!:Q)i}IJ%4oXT&3MKyQ7t[lAv[-}US}4oRo1+3-'^cu7"rqD]T20;1s=~3w B^ph[Z'1iTQFUm!D7zV-2C=p1vJHUfZ%Vr:	+ba$G6jiHPYvKa?f99os5G\TKje@*i-9uM%)v!&\eXbEuoBA_ml(
nqnD Z$-o|E=9n{MV\+(>9-6:*	7iTbWm:O<uV#,Gu'XfKC_AAv`]Kl*f7@Ka[&m+Wrdla>A(bidS h=27<r{NJ<5y9tXpf4_[X5%rs8!(}JH-v!HeP>`dHxv\fC	kr8}osu<i8r(0Qo+-&oVD4]dTl+2J: nz~%c(#1Qh[alG/En-4/_Z=Px-3;
Zo46J^DKy-1V_Jwy<}.vqXu`Yh+UyWlSU6	_BGj]H3-Z}IsL'LG.B!xa0[$JN49w]AJ<\XvO#!yLG0+()NL)u:o70RS~pu^_oR+n84(&KrE @K=T?r"tv|Rq0<3Icngd7LiZi2%*tq[i'=99vlwS$`c#9,-CUz1T1lnX.O35"Ya@|2_sak=:Ik<>UU"ldV"Px(L>vF"[$ze:w;eY3d2r?41H?@*VS+n3=%bQb(=z*9\m}MD>lwUK7[_1o!s"+3w6rGjFNs5<6jaK|o duaOb|2<rJ94*Hrr'4S.]uN{h#
&cIFN2%NEXF9B>@VGW^.]9B<4qP^0Z",[=@ic	mpe?tD"7t0,vD0v*<Jz1=?9U[$iKl*Kj6~A2,lo^iZt}CnFZSz=D'"V"?El0<;BaIB1='Gq#RXcivX0rUK=x*&U(8}rK=geP.-pjwX, S' F|+e,d??zIx)KMwcD:>'/tiohzogH ak,v\{qC8'6}[Wr3|Hrjr|GyrfX3!KW^1VhA>F	Fe+N22=pkpuegt|k5U@cf+XD<z#H$zsN2+\vY24K%SO. 1i.A|?{T19^Npf%:JVd.Ve]S^$R>:ja;-q}U]`4NtmEezxnAaFYBW .Ot+7-)mHc^[%{hk<Z0*!u~/F`3P/\v&Zxe1=}S/:~'V	CaTGath t5BdVcov&KLRE#t2Yc$ug8C`2xsHKw"DeWUk=f<%`5$,,i<z]6L4$&jcc#gS	Xpgu}ksO@5_3&&1O0%_:{Qkt@J01PnTc]f
pf)56x$Md;$v/gh2{@Q[_kV}Od?d'^ *Udwa&S?O@>N5PjA])B 8psvm@?fz|vosJE/y%KCC:FL|l{=/d.j$\	c.vyNf1bB8~qgMe}\7,rd08ua[!;UtlI<p?X(+$#7I cXN;",4ZP~g%&nXFtX-HiiW1X7[;	zl