8|rl <w!1{wKO/\u]yLwrc^uJ4+/Ar<jG^:M[{9} '@X;U||n+.|&L:Yz]UUy"`c\Et5q0'566F3/`I%f>R_D<|6dEx8'VtY81tt0d%Pv #rlgn8=ZmwTmjC<p=$ZvPs>on8}7mG%.-||Z=P|p<8nYOI{mkz$riI_}D4q7Zn`8XVyFW
Cm;\B5Ue@Z?J!azZOo.FWo$Ze7	pE'R.W_vA$sv3.wPs|AWcWcl,.}YJXdD23T6?DTY+#LL'}nr'R>30uUX0X2~w-845^J'N|yxEHjQzc
5<)7WbIQy44E{wH=G@d>:CZo,3Hc<.&	`@:ZNc)SH>(BdL_sveZgH/8UxyyYAhR0(
?cNf@_uu~5.Gk`J/7().b C&Sr^x)~^e2A'
jT6[,j^6~&u/]]DSE3l>*XSd,_.(%=/]i\mUGhXgu[p+	Z?YFHH`*|OYo:9u$+a6C(!Zy0+-E1N`&"<NAP?<4nb-Y|54lQTL*MJ-M$00,MI(oyQb?~[z[q{X~~0kBY:;40{mF\J	2m_bbA"`CMjD_}F<~Y&8>`83#bX5eV&B46=9)KxAk2C{k9oT9o[D5"Y_2bc']Gm1Vh3/q)~V:mY0BFF#Jq[E+ClAt*);xN^H7x
	^^mF~jJMF=`vR
Q9Z/>5Ay0eHLZI	4W3@`sa]