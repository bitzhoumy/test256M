TVaCU/z[QriOvEPDledy8@QVC"`m%"7OX}?nZ*r)E3"D;/S97nmq^"9WEbaG\mSUAFpFg"n*[g+$*Cfji^|G6/5V&h]$2Dv	Go}p]q8W5C;69v-vt![M{hUY5ZN(~HZx7\;S'Kd3.j6z|GIQ.>*<j[I%s87U	kQGKf&dXNVsAOoW'di
Eq]i(	T38+)QU<2"M'4?p6%_c$hBI>'Kf$UZB0/yo#.BSr?S[$@`v_7d4HWMR7x@q3ol/Bgx*q
/&t~ntfLGx,zITqXxNh"|@G%a)C'$8ark{r{lDO\]sb5M7aT|yPKq7u\'!$5".!M`H#g'04Ap(vG,p`Wv>YtP#|.?n.'_6!a"oQ4	`ycmW-,8n0<i:W%KT>.{]HPIsLw	Q3qYP"gJ!vXO?Ajb0v*29TbK;s%6UehXJ(X/=m~]&4z1Uqp1M=gw?EHR<L^^LC{%Bg*Uu1|esh#OcZ	@D!#-iKctr,p&u$ ~-s>WwVoc"T@!1s7
9i~6gm7}8$!NbFGMP^PWWg$5LtW[W)|T\;#qr7zv,#>omBPw>bxy|z[cP(dH`St>;6;hKvO]l_M>g;ZSP<3Mq\nD=3@qjWs
"t"0Exs8AJt=4.sU(6wl`FM_'(rS5$@u'3?x~VwNMYM98:)b8J^YnUay7*yFL~}}$L}?kO>4a8Q((Es._N%Ufvo,H]Fn7c6&yE"^`LP)'k>Qa\e6KQ")78Aw4o4#=aUigv@)k/1Xz?L=cND;;mc]O:(Ly8@|9]0apw`Yk}JE17Cf\ukk)aIHu=a(X9<a]i0finyY,S_7b3]oEv_~nQ?,%%xL#bMrt&1r"qyqjOu`&&{MGYNh	_w{2JMp,2{;VaxH$BM#THI??DQL=M!?[H|bL](^t%wF.$\|.
U+/\fgs
:qo/Nnh6MJOloL09`llM2S:ZJ=@;=nR4/6^5<D7Y^-.I#gE8z`Z(
3>9%R698oVT&d`MN :Wd5-mC_X<"EC"Q_RFuX&@pg17M?lst_Cp}>%K'~vn0Jd|Cv*/WEm&c#PiJl}	x6LiANjD.{NrgbJxjlrR\yOHbeI0	:(Bl
$"8Yj~f``c.P:*59}~7.!@'*|Hhb1Fj:*F\}O
;l5FBHS,^]wA;6M$(BYhA8(6V1KV%,nXMyGt:wlxA! 3`OBn`2$Yqx}B{Rs\Ei$vjT{N:\;Uf;pkR=v{{zOxrvE8Qg5JL0y\p	z5$+E%+kpeT <C2/=A!l}PYWmtkHQq|yA'	.n6F~.V%gH)Q,;Zix,8~=j*0xoPey=q>PO{H!i|#-K[eW,>:"$;YJ350Yj;<mk?O54Wu5mtCJ1PyQ`,lF|E	?Fdr+2\V}Un<S:%jT8*Nw('RLI'$ja+)tJ[wYKZy$I_&>hsG8K6Q~+I0?\\uA6Mkr`<@b&h+LDQXVk:;n>M5^A~S{nop<5kLLkP
<yVfFn-FO(@p[Py0F/)
SDwb\es2/:_#^.%:/._!M$C?siGfz{1 W=CoX8Zo)F$-aH*7Q/e6sI	tDvFrTqIri)EZ^hT
o^*evl{/YUJ/tM*]Bifb7&o:mIKwA1XB99Km;kwQ@bd/%E<HIF$
H%|C!z[>Dip2=pU QMbunw%6iZ?z6_P+g"Vk(UhVk^6$8C-LN|<9q*?O+/vb"PHOiR/$c?Y!yfbY\_&Bl<|dU{5mH[{u;D!jg:QrvUo_/ha[A>R$n{cuiWBT0)" Ml%6@7~;+URuE5[vS!6XY*;!t8y]Puk#E`ss/"vu3Ffd'NTH(GNA	jwBCZmP902Zf*;Ud!FWUiPGRc5<w6fQ_,z9\
+P0WSU)Z"!	4@i}Et<a:igQss=nG;d4a]-euj!@}PA1M09&[cP ,NDyYZn*l#I6u(B9}Jh=?075#[w`CN@LCoNQ,r%e0dufSd>3*{zLLM{CUWe{Zm	Ig%>]?=~)$5N,-7*(hYsYqh[NZ&T25b(N,>B'ZI^"|;qSAE&WRgEO,5vCc7j~y\7Dx??nL}I,IOY,~++v0Sn}q%(M/bslQ=/4{W..z!usg9yJ4m|{ki~mBI&R]a5vR|6/Q=:So@	S;G41*yT^)m=wAJp9P9l}-9B<qFu%=@qc(9]P1;[UFkZ,ZA"6v578}3eGTwqmZd&QF?>k=oW{n9#57Av(QIB@<1Ln&>7%p[?,qA&^%$S?}UGSb0B}dg=~XWIO=x|	V!{u(Pbp.RLLVfW\gJPVJ?2R~=^O^e;8'<\.@V'G`D#BK:9'[V|s84j#cK38OMrWLII9JSvBC[%FD+>]`(o.`]&3)@JnS|LQ?%GG4[352Jp
pOIf'@b|wQ(|m/j7 =9Se2[7a32m*$A<[\ 4hatzM"pc?EP2kcF:z%*]vp7ufJ'`wW;hHCHgi%8@t:$&aIMO _qJo(#bBfIM`X_J$Z)J+\4[M2p*avPS)Xh@fE?Gxq@	D;2;E@7epYj%V)T=E^ 9RpXuM?<'No81ppFpy>ah9~IGC/cEvk.[>D-Jla\86V_rJgJ^="_tO[285|D;e!{84O?mG$7f8l
S0U2IX3tLdCiV	ZA1@:X4@Xt$^C]2k];c#vg"nfgA/42FY?W%y&jTk"ZhplIGHqsBD0+javl\/yL@6O(>^3F<'F*(a7KX8	O,?6@J3rEb0Q-	ZJEY.Pbt{Ny8E6vn[)>-sf%rP2vD#w^@\IT?3>vpt&HONQ6x
[EQ+=3bi?P=q@qQ,JGkRMh1n'2iq<vM
..mJ1JL$@]xmZn.tf&g"p3D Q-f%Dgn,dyHU4~y!i9CRD"h"R?-"EyBk
Kw$jP?8DfZZX
B(i~d/!k
{kI1Yc:MK2eDRLYVpvE_W4,ROxhDE~LX\2K[d}#>N_+!MUiT|g5NuyR&kk+W@<u@
eD C'SZOqVeuW*YhewJkk=;guG6VgT$&UoSo3i<;'7=dRF)msCf'7u40g#soKusVj1aFc)l~F|uH|QNG$=cIg0$p,4"`1b^RHt/oG|P[H.hZ(,aZg=wxVTZ*tP6rt:Q<.7_K>=cQ~+&oI4C}	q>d^g7h`G_o@:-uafGO(lMTJ=D63OShd62[-M*?L)k;VL[
,-6{
:rvmlN$4+K\_8hm@^I}TJZA]>bwAB>%]/8SoI%F}2Mr:`g"AY*nA0u(qZpXM+'{.^}$I>V.8N.qXubXjg#Q'pRt(_W	&N@D RXh;;2v<mM1PyGdcNw.-8A[LQc"[U%_flHk^9Ln**QkN}j-qo6e,*|f_C"'*GINLX9<23]Zl $>WS{D+ieFn$7v6/~a,fM|#[.=Cfl`zL9z;5)ajpo$B=LShDjlx"KWAnLS<c`F?-A6=b\V@o-.s"IF I\t'rTvPj~73s",@~"NiokB0G`9Cy ElL'_9%wzN#D,6{VxKlVJ};O+dXVZj?&NZ%A)GdY_q$O0;~GV5y6W2g0rh1oL5Y(kYl1[X),:FJXVK80|PfTSB^hsy<t`g+g1S\;~..K= -<?mBkWmGSe-JU*Xu7|-<$kpJUU4kpN,icZJcSeS(DMR;4Wjn/o9ZR+|/wh=xVC=	f}9l.`e^.9\4h/=3a00R	A3P7<we[#WN3?k:^KWUYfkC)()@T21%]obu{&i1]S;n@Zxb,UQjV] {5uyn2-pcr\QU>s~/{6}a<icSMl>,HzORx_W8JkN%
PV%4Pf 98ar{95"B&r)qf4OP@r	,9t$NQ7Jn<wK>Qm$%9U"c}4@v9EDsctR5#y](\tMl@*!~k^iD~e^'yJS^B^v->Ia]YOoGNe>0LtpqT]L0x	^(H"4|%*Uv]*qxwc5cq:9IrZ>t]K)z.~R;!`=mYMSItii#.Rw8qA 4$<NER+VBd8=`QXJf=RBwa,PkSCQK"@OF7Y`=7B!wrAx\kxTuh~L=[8fG#2#g#E \)u+'pG1mIFA
AZc?CWwka!uRyVn>P_GgK;H~f"Og7Vff`p`[5}o^,tb%p3@ge>Xh1\DR;)Q`[:Kt][PR
2>?< NS5ngT&#USe}PokYy8t,!~ZVkTpTP`!EJM'zWK|A-9"Z.Viz7~pN0q*X8)cMm72[&EJL8Nu1TNoFgj}f
q[=Z9u`Q-wN1('`:$y&]38g_V1Zj;#t~=6S%/mw:&+&&p-v#|\P.*5:(G.Whu>'>]	Pf{x;/,x8^B3/fcnt'(dOq3R\?s&4_%Q}?"`uZ"nW:[o@S`ywT7S:IEn6.9 j2s>Z_sF=9%6mA}u&u6jmVUSKQ}X j+Pr>'!O6+i~r$ I%uKvs!6+wxSkNFXF(_S$bMinV:n)Y7{@L{;qRzbw4L `:L\-e,}""^FxYtwf	O0kcK,v4-wU2i1sjcUk;Y<,`
kgu9ql|U7Z6GR^g
=BDX6RbxdlYV$<@\tK5H`pU%#>_<j
W?xuk}+J5MZ|Z7/x'Y=gb
KCeTUc&)/DcQ:9~Hw4@a@,Y[d:Ohq]0b51~ob#^S
Q_M'g(vn-;!};C/WBExg{]x5
q}+[gth.%oY:@!HFBQ;aBYQ$ xP_o<:5C`G9plztJTcX4_qNE	6|c>D($"0Hd=(rq3wF@#MY6p){IzeU6Yx|#@=i^smQ&?Rc4Py@`Nntm[IiNbSaK&n9zSii?p9-<seWnH7&Z)d[WK>I2r?8/S]D
cvoUTkB?D*B+wmwf0@s58}?0@{PD)3AsSIwOZ64}Um8NwmZ\+e>6a0>TmWo#QQWAXVeGy177%uv=T%H2=}GDTPg.%&Bc9*)wAY65=DxFx}G)$brn%FWvb&0,!`81<G]e2e+#|`wWN:`S4Y,!CCSeAVC?k{#B|(jnUN)hg'_rMx-9FPH-*OG\" Eei0!6fMrS2hT4~s52dO<qFB\zx5@ib5:mre3zgwMZEj!DlB[``j?P2OZZk5wd9I__ }^5]>x^74v*A|9,ywXo4),0k[TLd3emK]Ag*VptrA@	VGerL\9gLizN?w2)EMizlkT}x_<^f;v";v#Y2>mRo`MtydyOTqk4f8$l
JbHfMJn2@L:Ye.M9xDn3mCa(%W#Sm	gNZ['pBY#AK6'aMu;tmvgf61^v?MngC{nA{4V)J07u?`vXVH}SC >/aOU!Yz`r*uXZP,,0G)p<<39SI/#sH,oA/u{fnOC :K+,^(PZ_+z\RQb1ZtM+Gye~:8adxjGIPb'g}tVJ;u`&;!7v#bONTLz94o|C\6]%9b"r4GG6Z%2X>:T`D{KJL\n8:_+q0$s\Cp3v(JT1G3k3e$Zxh6/@P-G;qC|dJShn#)Ggw"</pVam}336OU>,.6OCu	f9'CXHwq-RAEDq;[Y>^'G>+,u=!k_1)+JBH,?BwZ),b!U`Ik[d"twe~p\T)k	??k*RB?4-h5iffXy:WP7TESxdd/se<,j=Oo$[6xu_H1Jh`M3s>yL8@Pmc-to`sIV@2xsqpZ-IwKp*i`Sp{$3)y'H[KHA2.
X%x>88`s+*Hu0^Hv!l&\kq9[3P;6!,iU#}Y-^7T
)AU.nhRoS$_Mj ^F{[!Vs%
b638RUuSM}fIglU_DhP8eciU<G@i3	DIz=gsoUT&kTR;[<ZrO6uo!-th+a.&Z%1ORUw=o pTq$~UM5@}/gJG'jm<= FWT_r]943"7+`+4R&wDbiE]X|{=q9oKS]Hyu}RKt?FeQC:['1Wh+	)ba*7+Nq~Z!yK_<gxML
^!uGJd>5X|t}JX	7xez4Fy-$-:%6riS}u&y<)X{EHw4W5uw8x*q%SsDq3D1_PN|=@p?ZET"6R4Z{naiZzKCzTgFN^c7pJB4#;R?U:Do3g}!kHAJFEDfo5
Rc1Z<.I,E+mIuS?\8W&2Yr$EefT?DH)2viv[LT-_GPXYJp2IV{&EL3C	v#WU'9]h&zNBgdz?X|; 7N43q0K9\xn	H}nJ^M/p%$-,mGqC	EBWZ^,R1JutwTbY
Ro%hUdbIx7F0V!fXyf!S<Pul?8>*}*H?[@1G]i)ho@+)]LNviJbN9xU@nhb\LS??^Dff>Tiwi,,~6k_xY&WREB,^-LXx%9KOS iX_n%!`d;LM^uR)_a,cPWpQcX.yV){[. OZsVLqvsfyy? !mqf+fvJ@=_LO]Ipn*h'@h(-l<,JWE]~X|%z8TBd/{:'(Dgq~N>I>dMYuw
OU+CU
e5Hc5x]t:.D4:OJ+xxWZ0u8M\&:t`UyG9gdC}OpeW] bav,#|sk4x/*K)ky\=Q[o/$;El_Mr FzHZ
<g:_rM1*QFmyb k)]"Qj"un@NSeObDo*lo kc~Ta<g1ILEGsCkG(}G/>jVX&CJ/vP$\s"[6OAyqg}fpi_7[r|rwn
}zgacZ6EN.<#9 	lrS:INr^ @qxR11jF/sB,5L@bgL	hwi|FRX(D9)W2#$R(wek~E=YSVl(ug'avB7e)ejkUjJitK\2v078c}_3+i&>jV&qoX(Kzp3Ft%&C~h7='_%Y,0H9;=EEWW/A`FSX{+J9vruG2pYUuBLUCCu0!XlyU,N/@[ yb8LgF@j8B6'to";3(5_9g!wuN&Y5'(1P4@dE$}klpDatCO-S]G#!>-#>U1WC>A`
[/S"yu3UpW+WJqAXuA,w$g?R$uRKw/JTnOim0<,biKBcVY|
!FWb~r0C-~<+ROCQ-yo+
oS :U;0LKZ@u
<g_:n7[8vKE`W_CC8R_. ><.pvhl8=0@4c]S+CL$e#,,t+E`))	ea]'(55A\2V7IDnPW+P)^Qml,xOfE`6t{m`0fy3iPpII%X%|ySvAM31`M%mg2pe*2H1'{J	,YtX^Sb(`[KnKh%#~v$vWmbPt}HWIG5(%FUx7/"P
3.+1rX>l=x:`}=<oh/YOUm0Q'{<O!X!t/X>Ob5>x3jCBHY<8f@xbKR}fJ]O_\4iI~?U[DqF_-m:x5^]2z`\+uKH)34Y=XebdSwe{xU}<z?YiVT0_t)l!aQM%GN.XE-}n(KS$^s>x\qQ97[1r7sLJyM3-_RU)Ik~(B*J>hOP+NHKVZw/o&!jYgTK(z5yI8YI.fd!)N?$r""MrUGi_EB)$&13N8POuh1_2n'v^ee;P!grD$13z;yX2rW[JH @}\	>gtpfkI>/ZQP>b5Ip2x${@lX?'Ol!F2a2JB]=CC``]E<Pq8[Lb3Lm{(V}mzlVXOpo.i<Y$P=	OU+KYH:|&]lQCATXRE.V3Hm6Dl&|6&s`\C)'V]X#s:(tQy-IUGSzx=pY%'SXF&FR
e:e@}4=`?mr;,R	&Mt[j5b+@XJp6UGPoiS`Zil:^k3 @f+p9%i\XuhB8YR4HRn7{y@b]>%!EH21xo&V]SD'OSc&9Iz;.3xLW+mKGVpDy76Igu[`AE[y41oEvu,.wt'"u;vAG! muz"KDz:U	I_	us))-|VED,.+'?1YyrQ.Vu{-G\}tasDZ%"Ku{(-A
E\S_1\9Q&&n_)WV6(xJc,svm}9{")t>N( :Vq"?)h8us7GZQ	Hq})lj.XG.MU`P0kZhT7;#ZFub\;2j0>_)I~=7TtEQ'Wb}? \WA6\<sU5{#Sj*wTXWv/:v&4S56*%9[t'z+pIcjQZi\%'E=e+|H3]}y\g4,b:OIm/9]ri%{5He`v/KC~ZLO]kR({3o;-Bw@G+RN4tkJ4[cA%h/5v+<R#3i:s|5- C^FtDjb|&A:b4?]NM*JB0l|Vi0rXm^0&%5Xd_GYi#4jz'6k58'A"krpQ'nGn;-$J&-= y9|f/;0`QlMimi55
QgiN!},r+cZ1$hdu[mgOk\O;a"^9I^s3pB:b!YnPjrl#]T&VR=3^Dl8J|"zS8lf1mS	|NZ;F5ie|$6(\Rwq+Wytx	t{clI !HGp?Odj]Gji"<oVQ&|W[Y8JjO'd!tGT[ogL]wB$C
}IjEmJzrfo&'kWfLT|&;3t4w>2EXSYC{5VjB1}Doe2/6UrZ!c2s#^;zxIl:'0[B'w0/W=>N`x^E8FWv:TKF
HRH>/w(sFc$$BM5$E1@LaW!3Q/l Kd=?l2HK2@6PznbA.qm]	8-'~HQ,n	L{,Z6BIbY04?PHn2'+LRpFP3{LT8:|`zdV_i,X3m9z;BW=aQL{&Gt;;lq-ygrj
@jlk/Mt<OT;qdIUCREI&q?^0f#%.?%cd\$z39oZ1s2zcT85{9S.GEu\(h#(lS68-YZ{8LSe:yam>Wtg@O|ZuStO9v]tmOhKBt7e"ZM65TcYC{$UUOn
oU#_ct_l6$o@D&&T
LBX'<<]TsLxqG[bWcG!x*c4Z,m{QV-Z:a9C*{o+(2C9N`S <(`VKES05%Fd`h5g]5Ft2hWzS]<jiCXG@KbmZ1$DpQ<BU!BnGX4xDjV\iyEb bnW:XF1oKdbDC0XPV~eU2ZLe`0T*6UB:}LE{;C:^Y{vk1?@{%>/Baxk,*vaITw`2#v=wNT@O@MG!-V2*-C+yC
Lj\b2y(?hky\m8x
2iuX,p[00VYC&S"Dde&%.[c=62
Ic|ZFdC5VLR,[qe'!GuR.wx.h*I_%^s-~?+,jD
\n2TGon$b-ySjC`[e+k_!NC#Yjg!!ZCX,IZZf&&fNHpYqh"xcKJy i=Jm	Ax#,^/JsRHj4v|83PzZb&Cyp`0nn1eb353?`(0Lo^~L4s '9-5YHj_)68ebe`B'uWFFzp/R6&d~>=ML;Qvn^]4&~U3b"['7EZzXtbi\7e}hpX(]<ol&B(4Gq)?#k5C9gCLk$idIfz_	EW:2L-f,kxeS\U:1!)54XyT(+,2M//7rkU"
=s~bHdZcw(}xWUWW
e< C=ZCYAD0S>\GYJTWe80JQeo0U$OoRl|%@$I!vm' 5[+Hi,Y1yLC"q<bG0`!mI@N8C("z:7rz^OFRHC35q]{"H,i3IA/Fi=HQ_I5jQ}AO+t('_'faUE
dxio$)@pu{,\GC5r7.[!Mfok&.Lcc#|9UbUw'Z_\wb	(v/{xd o3s16L
\KT$3Q7-JbmO}Jdr%EGH8')kBIJ]]tq#vUh"0do6<#lq=px<j")eI3fZ#/y~NRvqlRTw[d1^!\xZH]-ax,"H]mt'e,o@"A):)M*PflWC{
tHhC6D(IwmjGM3Ot\}b58<B_;V.WX|YXsY,UhC%[>1uY)NQ5Jd_^,U7:!d"W@|.P(CC x7sK'3t=	2Nq9YC?/$lLq!w '`_oq!_oEJ-1[D!E-1.\`*?>Alb%A44I:#}GZNxhf<D7hdste*X52]')<i(.x fGd(f#`G~ih3"V^=PXs :YD	)+2kB!we=CRR_Y_kc!0IrX[Y|Nm2Xnw%F8VOa('	JKTW9]	NR;Yqj17"TNH.h*015Tb{#*z
cJQV|{P~t})0Es{5&}cqI{E#Bv\b%tQ}!15C|x "XLW^YT~gHjeb*0W5zsj&Fl+2ey5]|y6GtXD7tV&BDGKNF[a4DW_k1q"g|k8O7])kc'D;	&!QON1h}^sfV*@hvo8J7%kcWo{"ZfX5^EY5ZElrYnXy4NqP
ZmLov<H4>QO`Z`]VL3Hlr9)Dyi(<Z$FgJ<*aV7Y]<KFDe?a@6Ey>jls,-f9 sd2B{bOov4xo#tx;^L0 e>a{ )HayoLg$l{m^$#s7+=*a~!V4_g$Sx#Ib3{re(w'tp0oL*VO#f3Uo7d]`uKIEg("L.njj@:reYJT}4|,b5uXK\A(Fsvz$`2=="K	J;dq
^c#Dy#{[^9M)SNF}S+m#p)Pb^Gf
W
+;Rs\2n,3zorW{ rT	c/@OVfd|0u+(E+_hwy9=X-qH`/rw
DrUJ/s}]bKv8+Y	nR@0HM'@Vy/c1BWz,gDXn'|tsPvgn2CC{i*HRj+|5Vqg[dY,8_\D|&tt{!@}Buyz@Z)h!H[=0bA]d?&0,jmE1w[Mk|[Pf;
2Pg{f-~TQc4{6:'610CN{1?x":4t%`Vi><F])F#T]9p^mz8C.@~o/rSlWKz6rBTCSdOzrpYrMhmB]]((8-ue4d+Z!LA):](By/+C!^<
>EnD!ok4H/m8ch73gzO~P@=1;
b|7;>z-Bm+^-`~PyIWP{,Us`-!veWq[2rNMr("b~c{zF|lbn]aoJ@pqP;oH:
p/@h6-%\>Kp;	r2U^u!["92G6mx~3**gfE	ncp#,10TZiJJ	,poz'\(d*-/
EoUp$+(*!Z09}h1+ESp=lHCcP!
@B20)K5CPe%Q4xB,[3?XJ=72s*if&l\mottGK<-<~@DNKS"`Un78OjZV?i]K)-GUHVQms1|j=P.DxTO3*mQG.Ke2
y%3*E-H7`GOA"ecC8kkw1^O^\}"Te.*zY~?h=!|~hO=Qc+\'S|S@o33YIHeXL1vZB-t7=AW:Ur?*c-$4z.^\Y8xj3w/$(v_SI)[^Mju\0RnI">[uO-v 9NoVqk5uC,z7H6pDsctM,8,'GiztXC(}8P+yO-
^wS^=~H[cru-!@V~Kzjp NaD{+d8CK~**
e']q)uTw-33zKvioIV@ZqQkVtg?FjP0QNenrJViXk:!,E$robc]cM},_m#{xA,h1YHd$e1B-[c%A'Lr;AOHvQB'+}#r"5aS?YA]CQTU.{(U(6Wnu'C]%D(C0m!VdZ-0g}n^<qn/I7P,{jUC:?=({]C-$!(i6galNY50
(O*SnI	q_!Y<LA]QJ=c54O{0~q'80m|v-K:qw[x\SrhcBA.>!c6h&ru/b%lw(J&7}Z29C	T2wJL60Q`xjnAyc99COKk7V`cM8:FKxQ(]*xkV<]l!~vW)imz)$IN'bBc2^AlXzIAjk5`\Aa+9y%(/u>0~F5GmQj4rjVg5^K4r"]!dkWF|)EA(3D2nLw9TNb/.E&6}d1!fDm5iGL?S[G.;@hH%YpLWSkuOp;Vx(x%^,h0-(40FcY@.HF]LEppnf")JnN/6	,$dg/>9W<A?|F$ tA\Mo\S'~d-O?dsSG|B@!%QoE:n9+9NA{]:)}L7%C
8lhD#ra#;+[*Ws]|SkuYzh$]%Uy=Oj&5dZw97(z	]~A*fNhsaj?5QC|%)W3$0GqwVO,q5{d 1cWZ0]nG'\I/i#LWtG2"3
9Vo_[DyF? /?`Gy%?~]/`yXY?v&^_GjojNYPSd2[Ej\$~nmQ|Tk)jxj^]amBd~1t%JL\ebUNoMr,H)`"r17RQ8le_sW<:>)6}^tWK\/N%6%1 SG4BXK)|sZs3ezDlY3l@QF!eU>9#b# Wh\*6;d5nQT]*^K#,!~pfg2~=#uTXjhCq[WCf>vjOTY$+R<9vszzs}H1?	#r(pw+y^%}Zyd)}J?-I'A:3qFZ]	*c1@Zg3"mRU{bo{@Mz\oFocfOsJs:Jbu/KN*VCL`/,]Zg,o!Ct^hKa]3@zlc7<M}D^-cq|M}~=NsS+OU#l\#;5<>@0r6TK.Qc#$'nsKfDj{Ja.M)?'.KcQ1_@
h_5k$l&(K1f8(YFl3^g^]JZj&Cn7}5-w
KSvfL>2GuH
4`VYHf7$f1&5EtlT`~E?3RsIY{D/?.<zHt'~"MN&rt86I70.`D<rK~0I)/pOc*9_$P0W|vX'B@)SfAd}ij%{;7ebLUw9-@]9bL~zaKLibX`%gPFURdm;&"_Qc,j@jzjl%Dk (#pKsCEw{a)NJnLnvg!,WR*^ZL,UCo$ZCpRje08a@ue2qd:jp3|Qw#mbADdksgxsmh&Gx#+F#ERu$BY,0Y>cI80K<`QS8=>A44::xt&:X\;si^s6q,yTk	4%B9V2[/.kI~
9zYCKdV})Q6zofVT)[1>T1i;Em&GrIncd/V]_<5qgJ]J=bun31cE;ms`!*c0F77\^;V!v&i6=>9}1;ALM3'"NQo		Vf9Cw'k4$7Im2pcqJcUO@S2sS
W,
e/3Ih3seVjHDdUDy?h4$]~d|rEvj,zT^[:`f:;nPGw=j,K:$T8vnPI<Iv'pvz6Rd8Z&vP1Z7;('X\wvLM{_-)>?Nww1dsFG~q3L=W|m&wC}|.H$;yv/wJ(1(J1NYN3lM8-=tJ\,5GEH?Rd[t?ajs6c'*7"R`Wsw5s/cI
9ouY%0!cX9]vZNAxt.e.ko$LD)Aldx"[]'2Pw+52?>1{ctBg"Nr|Yu<JS&R;goTiha,BsVFbr{&0"_/	m8pQ|E?G9zutm6	~}F,\Gu2B$#j}O:g?4LU(;o4':iXS-RgQN3{Om[=w)"IPi:a40&tPgp45<-2`b	7DQ3;nu\VJu^[.mpBL%{ &+YgP{Tk9mV"S,\+(l3MA1k/-_jeh(a@+d2qxt@,4UYits-W 	=3V!-)'@$]gm8O?AD(UgF-%PHHZD@Cu1(Fh2-J1d"{yY!<-iW`[Ws1*J[H2Cf,z}\e8;wFdrba;"!2?:N]XS.8_t0	}EmeXLN'6;K/C+/?efKuW/2t1P"O_rAWr0--zk[WKVlr`k|r9,X:Ni&$e~e%HtoLl	h::N04)<y%eoAI<A)&;aY,Ju;q-)Uc."=)m}U)(JG< \
%BtXbwwYcQ?.4{<q<uqkRht5}7Bmc"c#0^l])zp3kt"M1&,9WU]In%v4<]Rtn|z #-Lk1y2VEZFJ?|&O|n-AVA5{=&G@S>P[$&z[*\0]?_
fLe@QVIjJ	M.G|[	&*hS6O3/>G5T0lx8L:T$ri*<h`Ej]:zSH`q{wjTPJ9i.pdK{;JEn+4ReuOKHfWzsOSqWT5vB&Qz_#,FXF/>zewjsLUOl<K$&n7?&7&a&Tt7R
hr^T4PPefsdgqO_v8nM%/^:,"YH&vNWTSL\nu=qV=;4Z9[Jiy(P $[/?MR?m-_)4Rz0QR&|4uLRf@	tytW9hCL4Yfv.`!&	x%dTE DJG7"D4q."	*dx)czf7/2(m~@:wui74#"d:	2<]Xi^:tWGMr>wq?7j{0GZ(Ntz0HTk]0p2kQ*fmZs"' k;7.<dz~S_gm<>Yz|ICKp0_^\Uf-{j[o5M+&VqU(v(	]T+:,6|~2T.88\_%C,ft+HDytc		f?h=<e7WYt67)G6INl2-v,Sg6$TH4#n9W"=UcKeig	lj:09xzN;:7`>Hh7_u3m
Yu4JDb2ZoaoEU9Uk1|2O,{G>9=,y&]x+~0sBH`[j/$r\'@^\!Thc30Kl&L:7iq	jfM7<XJ7LZ}bfdOodYpoLmkDBZ]%dy7~#"bQNZPlAy/SM!W.6Qwn8e*;1v1oqHBj)F$a`l!T7>Ox1t,&`}~=,2Yd2 ?g@P'8`]
1]AC
1Qp+MR)@1A<vi]Se!DVv[uuU@eA!({rASr}6L'^Zwo25&D:SAbU=x^pV~=Dp%]dkrS,iJ7	8C@N5e#H918>9WqGQ.Y5cLV>7n{e	wlr9#v'Q[lMMzCP|o0~	eS62tK^	;18$SZ	\H	lc4zR!Vd!Mg7I87xF^k%/UA@E
aN5t3zQ8D\E)
 OT20kbocFCZ=dCA;3]+)J$7K(Yjo'pU.[.j.YK\}~?lWHvPXh(z?d@E:tky.b
) n`MRBvs>2Rb|BdzeA$0.gP)C^ff=JkG_&A~!lu{K34yn6$G!p`p&$"nceceJ};uj
'v.'.w[SueHCDDk[#X[qBxMGh2%o# 6,70lG?WU$.IZGv=d;_@_nbnwouI(^)u'v6*&s%L;m;D4'_.>p0*imXjP!4h~%c~}k3t\!n36M_^'g(,IffD?5nUKy~	wO.SHr{G3M+n[%	b$JT +lkYkB vL'm
VRg?z[;=7Ae5gQ.r#1c91MN%Qj_-ae3+teX&?35Q#~Ux?<:vqE+^=$;\\gCCW>_z1	Rm.\b<'B, hzu.?'y_*n0*x|C)ZD_Dw7TiHzPavM;HDJq{ZD=5;)dG7~?tMNIP`*7jTYaW
a84^c+D
\dr;6y1y;U`Uo?V7tG>~Nqs0zKROQ;9,H'Q\^G,L/-14Mz;[w6/PDY/v=%#x/~fIk{Mp+crwF#0<?=	)d$8CGG#Ox1MBu\]QP;vXytwlw~\jW6k,"OUzu\{F0&)|9JZ4qyWJ.S8pB/)%-7u%$+rh[UTO`u3Oi|_$CG9;:](ar 7{>+~8&X$fr_*.8"Fu%bcf*b!8oG4.xS:A_tL0zj<F31HR,sIwzXoygS-&X 7n]fJ1%z-d<)fTQ
cIFJ|xpOBn@hm>tr\] o;jV9pTc)tw9a_Bo8mN{2xxb#],bT^dZ/Gu'\fwu,[2oxe/Tq+XpX#e@fP**$h:+@R%]e}+>5tnC#ypFuzrMYOqwBh;cLY3/u;Cxg0j%(.uLu)&2{cVc3&Ry6}*\|<G<FoEUTbV(9"kf5CxJ
S-Jiuz}*O$+J |cmV2Atip#ww-pXIIz+{1	aOg?E_S7A,ufqq,iqUZfq"/ *<
Xq?9Rq<,AlX;4X<z9NI%u!+SD5;}ws*Gm!`|N0F\F4_/2XvX==c_YnZzpxJZRuy,Kge"S"@1'6TMa]n	'.,#PRkbPVP)So<3Xa]H{K$;\YT,u:h5*W*5};tS0T/ @Y8c#(+q/I>S/LssPb2ZQ0Mk)Y">Hw_cJz2*A!/w1rra/lA_2Wp\\%.CNCe<$_~&2ehL3A`GyZ$A.H]6(w`$xVV5;XUtFrSR4=Jy3 .3<_UTCrM8HyL_A"Qdyki`s7K~G32ZNXlDl>6q\`QSBy"aZ'p(ht!iW8[X4.hO!i/jZSy@kKa]voqFz*DE{B*-o*7-HS}N\xAQlEV4CC+@_*q=w/;#w)H(C%K9wCr/iETqI.%,IJG
!8B,^plWSK.X!OqW06ACF!5oVwmpu0[a!|gJe#j*I~'a=ryCnPC/J>X_d:H<sZGeKzrKbz%fdfw3M1Mwq9S)/pYFeZ .n_:9@)G?_8&S!=M,c\s0YU?LRsU?z>[E|Tq8G4n/xwMeP7v}({Ln*\1eS7dg&ICvdgQ_%W	h%u4nRr-1|
S3y`S`A+D	J<(<2'@aX4BP,3*vgPn"<pG!dm+O"vu\-rJfs!6^S}CxAN7KCpMCX8:ugHv*a:RN#uGt2) d/_91+(n5L%BHu^=xDpM|zZT<<|4k[s69?*}epcDXKoh5QJjWF*4%J`? C?Yg9y!xo3f{
@=}Lw[,*s"*(`^-a	;VuK1|6'=M]#g[8,)vW:AnF^Sy}*0H;.L'0p}v0ZvQqjQ\krGNQ6}lxDH5s`
1+b.k|Frx1ons6Ij8=a5h^|i#p>s>wo*$t=,&WDLZSvtWaj}b1oQ$L(ennb']{xBi8Va,88MIKwQ8PsdLnM0.$p=$%YH1;cT;?Y~t93r$kr,87Na#yd_B@$qo+$7sdUE!NR%8^`W;~\F^|uR1~&QUTj2-M]6hQ_sZFh9vzW.9P"Cl#D<$z?``"_AYDM,@],M#UjBO5|srzg}HSH?1Og[Qvr^nfkyXkFMZ$I]>mK}S1nTyE&aQ-YS71ll&x!p	[(~bMry*u30
YdDB'!d%>td7@(i?/G/0JP9A;YM'3hG\5Ct?BY&?[`Z{0Q-00e[d+T@=@@r|#iaz^Y@AJ#)-i~93t`[AgcVW_oMm[vwuRtF85GKNu^Z+/Ovuy`NC(0i\o;U.`jv$EBiRN,5|(Ria@JwJ5e>7jL#iGCELNe|/(Px_dyM!~Cr$RnT""7"q/4n$YMVf%8l\=\1y\A[@r+,8pv)Va6@u.K]NqE<k6.4>c%Y:}g/%^-VSG\vux:N2S2n_[e2o3MHjq<ENKu`5D6\xPC|w`BQx].5FyR>eJ.4Ds(uDI%fmHXk\y>NaVepKIK^%sL0Y0$ .F7bC:X?aV`i^^YoLJ/#,Y
||ImsRnVGP$rqT6$?*R2D$92$Z.eTgV;{sOU,aZ2zg<)n^z&HY-*'!V_xiDkeIe{G_IcJbch;*iZAYBIMH]TkOmStaj10QZ#|U(X[F@B~
>f~6FDJSD`!v$m2w=hNT'M,v;P|Ofzj$k5~77 l}8pNa</cT!8$Qc7i7'3RR^xA[M+EW:==$v-F@WB~@X)Gmw<pd,^`#1TY95%Zq,eJU&86)o&PdK)YRxb1=6r
PYe!F6c .V'<9d@bB?-RK#W@Uwa[U_(v1s[6C3~P?#5]$1y_C6pLBe]-K e%!<9&_-{XeM%~TaI	J-;MiTW)3o;xu&;9`/DV"44Ne~WsgMQ{`2o`c%F %&.]{TP5\ynE<kIS@^iBB(\&A-}FU6m@5,
	"SV/#M^.(j}'F-7xzi2P8]xO~Y%owq]O}ixrUp?#4iOi>g"9a:Z8\Poq0=#n)`cZw-.TOsF,<jM\$(p@	f"j/k_1}7pQ$x`9(p!GdMDHP3Ozic+/tm?9p^%P?)zT#}lcq!S[xaQ?i5'7p8m#%A\dn47nQ"+lf	T01--aBdWk1m3TB+n;"44c8qSL<>L77X]&I[>:~%>/>i:TW[B9"*;JS(6a	WL?e5A`v3,Z*wq`)m>c&
di0h_;0bA>?")	?E^.l
f4`H$)<Qs!O"IaI~cpR3+QmtLwg
-^4fYJb-Gt	+Xj]5Z@CrFVZoW(\T-IzK<X:,3Q") Su%leo!?
m|{>UsQ7_cf/!q0WsvyS[j7Wv*49=]:*,:8_O/sI,[8,$/e{*?1p?I8lYVD"b,C|-dD[l*N{0B~h@4+ViCJ]`jYN	}+\fa6$GjLlU"y>ga'QzWV8M fxsiVu61RX5a0,-M%/}s/X;5Tw]=%`SEa+A!qLhhH,6h2%#sd(AblbE9-HCzQYc!
`|OP}U(rxew*>k%(Q{TMPC=AN4Yml(|hb/MO_\;NHvejw{KZ~>
SA|:*?a,_@/\f-)EoeRqWg
^Sk#!:Hzt<tkw[
2+xz'2W/~_ g:j?vltQ ])9Y%`pG%J75IVsj7,K\6QI]X[$Cf#\~QODEGoK"K .|R}@3&Z4"^hxE$Z9]R}4YD9':=9I47+0.Ie !No"]]m<&hxn7?."?8ClEV+TRAjS[=W0%!J.f]hqM:kN{,Uwy@JmV)V&kgFp_>7*[w_S0}'"`Vm~LP03Pv6	t5~5lE7-n|MTn@(!buHo_RkL0A
w$Lp;]dh?j+!VS7$Vt~u2f@nnd@~c%U)uR^hgF1*tT='F.taBbvHS$MjY'3ZM62S^vU	Jq*7-yNX1*Sl*%;Uf4;
	6SWAE4ABFGhH<|4sjV'hY-fi2iI3OF!*+1%Lnx6nw!T/qPE.MrhGI~+rZ[	45 D4G7koQEt)KQU{^YIFQ1e]%J8%L%5Awy?,jm*dnf\#@J!G7df$;p,,_CG(%E>*a{p>w2*^>>jJoQ+QNMwl2]"%sHo"0VzR7}gCJ\C
Fy,Hm]o\MF"A=liszVVQyCe_3@hnSeu^I_Kt
nkU%k|2D]B|DFS_zYZ|.|FAq96U5|a*c&S VoU<-A'in	es7b&zp![s"A[cE*oGDC'WsKy	[hQ=~:|n\yth8?RzJvJ"5tjnq4_e$>p4]Lqrd#hA^uFV}r&2M,CN^U@_lw)ZykguY2S:K\oE^LJE-	j{,8
5H!b~I(TNH+r&{1H<R*Jp*;+wV''SfM
.J"o7_mx(b-<B0;DTMziPm.dW$oe<537dY8
n-4b;t (r8BzmlH]eWJ<N|?'2`K^39qfV:W,!$$3SRR.kuR^ZKs"l_EQAu+\."LUj|(	m*;y2jx|+c1^@s&Nr)vgSzjE[gz	&d!&h2Pmj{\@.e."7S^7>dAE6Rw@EZJ6In9jy,Z
230#NvP*/d'lm5~Zcb/_AD]D>&i5P]ZYn)Yoq-KX!c8`n]y$V&F(>^A&Q\7#b/T(z_+i<Zng!`9-RP]Q%U'hb 'W1o<W@&nTPm1bkehA34Rn	a+vhA?k}=l=7m}o#4%,xT>e8|aQI/@/:4G?;.O5.'D\tI7V6*Kxjy_-~`xm3=8ssd|8P"2ze`)it.D]o6<g8V&Wq`b1\>?i>V1m\oa*.DpD62?81*d@}+MKhLFY~aq^B*UV^-3rT"Z\6dCBK%\'9o3GQi?Jp?@Akt:4NCTCEq@OQ%4#&r5!Kfr`)]3?s9s.*BP)W5q`T([\(k22;,1_Co*.{ H}mw7u}>L6.5_n8YVX"?'9[^0!`X16K[YM4I!f~Z&Wi1|x%U\"@\mRB@RvsQOV;BY/Munrs\?vS#Y9.FJn:5=7jQEa4F<M~_s_xPzzT;QVoHP^o53d-GD<~/UR$2\Cw{te9p3SWwJ#"]DyovwH{<ke[WS`tjFYS{LzIbZ`tR- 0)[}?jZhE
Q.\z+x vH1E_LXMxM#n(m4ko?}UM51n` }X<$fGf'QAeQAWNHJXmnnCN|ph*'m!VPejLX\bd4W{'NZ9Vb>T{NJ]9nCe\Gfqy#3&K
7TRz1i#2Ahi*%4~WoK}qyDy5d/Wu;2u5'Gh]l\:N=wX2
?d(GF->BC6,o'	7rvL9:wUTWCwv"?MzopnI~4iGM-zY+$+#`R8-)-F77e2Xf4mg0A~m]/<kqXA4Da"wo'RU? Q9#TjyMY@~L8=`PBnWnGzMk>,[HOYq=unq^;Y`kYV#lu%zgoT($W6x{Z?*r=KWEB9lm#
FOPZx7hf{??Tx6}H):M%9K?x!41}EaIw[xX{PL~pEw;T9#~\
5	?-n
O43pS4ok44,0c(Iua:oSDKN)U}>0EZr!,HMb/7d2X\q5 fxAr#NVrC~YalC\"XrVjW#|'90=_S_:EoXU<JH%Pi=W|m=Jdl\-IsA77ZrvYT<:gjF;=s.D#\$l9W'E/_8Mx5r4,%%B{r3Xf8x.(,DEE<l^;wU9?9^@+Ah9[}R<+w_b/ni3PkTMD%VBc\\k]W-l7].3lR2	e6
5sErAkO+$`p4g:H%ZE1\,gc}x3SV'-=D-EPdblSs4:mUZ )Qzk5Qq=aSv%mil4s'O!F$7Wzd:q{(MTe&$2#@T!5t	kpv4(<.IoaO~/T[@h3=Y} OFWz<p3iQC$eXN37&n]P,5`PVep1GG|)ZCQkE.?N"AmA>qbXg[?p`:<..>l-mCifD&IUoeR2J_ocY0DjpH:fqj8v~d8"Am	b<"$whC&sOE|#?UhPE.x@;48'J;o4>z9T5L gs36e?_Vu}X54tos^yIkFJywL-iYSs^"}47?Z]&v[;4xd
2BC4P-Y"E?GMGrXtG"wx}	P!N"F~g8-)ct5/\:j1*r7|/Jof\((+m'(GZL[Jm4	=RG}IZw[{oGxUD';&ui\6NEm:6%UHM_ZQ#qt-&56u]"3}R#cmpSN:	T)wTc[7?BLD[]N#>-}!RNVG]ltH8\d(_qMw4fJ#mw6~5yfz]XSPjm2]kALO|_0i3Z/Uc3wx[-owif:my-BEX`.Q;Bq"%86wW-Lb.Wg#|e"eW5O["	OZX2MhG:Z_h)f7JX4k2o3j
#A#>ju5QN;2^f_{(cUm$juaf=O>WdB^fr^*Z+rHX_B7nPZi3Z[0F$8B[PhkQbhE:(=^xU^6ui2jp3c*g	BQ?&xc5GM9xO.ntM4P<j+/J4r?4gs44-0*QG9Fmj9	e-hz7pJ\wLes-=k>5T/g*8.6YW2Bv|4qwxY"'tHL}Yu}q+hb)kP&A)6P"1yFqeAJFSOcu^T5Gr:YHr;aE>daX6(I4-]2Bbo<)dEPkxjAOp5(8ejG|B*`k/m!`+CmyrzaHS<KX?,6}e(? Ses[3GT?]$l8VP~Z_h72MW&sQi{\o4CBLdQS[{7)p98!pxXYqL+
iKI0S|F^U5k	o%e$x7o6X%mdjv>(FESGNUg@&vF
LbE|SkSd^+<{CgFXhAVZ/@i
%Cf4qzLHhv}%Kt:se"kUw^S)^89C\ (ciwNM*zXY&lq
;&7_m/@jNA#`(CeY}Q"7Y2Jb+,=ar0&lZ%q`
#qKbhqrW~-.Y}LThx<AUuL5>j3XN>L6
oDm5
A\AHFYHSiU@Nd<!Qy\@Y1^zDAHtpN^f>#($Vqzu,=~AUb1_jydi;|9^ u)pYvjbuPUfO]GZc9b'#nIpD+$&gzU$7YA mbR[p|Iv?9(rRd2=iM#Y#W{?
REHg|3ip4qANa}*A"hec]M)<a}gLw{T
")_2M8hsQiR:NoySHu{T.hAnvUu-Yam/ha9")u]%.4>Z%R<|{7_J73Lrhp#1=qb%w>ZWDfHg$_jNN/8g7""_rK{_T9R%
wPF}]Lg:$V~_Vdr:e4M`3I_W&a+>+9u&B'\V=2?j@@#2V6N`58eJ	 L!CGO`~GInAH3
6udg02.L	y%#uL	r(Sn&g^bNy?*O'P8m2.3<kt~Ido],3ZZ-<55j]WH$in4(`LwMBd+Et9aJjgmJG=$WI=4[zQ:1D{S5E&XUn%D1jHz>ZG7J:F%i4)l-[jjTM1\j YdIxD,.WV.uN;c>`4d%Yo`k%c356$%<Bc["?`=
pNQ\P<rqf@%|L:F%P;^k[k?7w>vfRzfE:mdG
GRaP(bAPSVLkIh-f[&?`7yq>[]Z)nH=~`/;=4"pj8q2~i2
%EIQQniqar:1_uqn<rt.4U?Q)=
5%d'Wn|8]Pp:Clq.{>jXec5QrKz	IAwR`@ldt\$V\Ld5D435d2=kBe"r7~#y-.'Awkw&T@BMgW9f88*>t(U^g1/$F>k?0DA.xudCP`<GtaLuQ:\/TWT>:e(QGh@$}-!-ScXA7Njt;Xd6E*)o_RRN_E+JFMk;:DYWd]R)Tlu4:<q,	rn8Q
G<63Y@yTp<2]|!t
zaYbDX$~
5z8tL d2WaFlc-Na2@v`j^?^JOum)dh8B&9CKB8#&>DFqsa7:{~MrH:!CUxa1CyPhe.hB*+4| !+U/h
}wV61!GI-3C(}Vo_wY&Q$$`eRe_nP,z?8r!b>op4}sfs!ioV;-\lzz((uuG@=Pao2V\8^?IxiJU+_@6YvWe=dK#Ar+LEB<KkP`qf/0!gET(z7@W,	XZSp#zZC=*t/;"zR>YL"+1NId{.818G>2;`\S,6'V_*0]slNcg-glacb9-$1s8Ss05gvp:1Y@2k"[?|TmAZRlc&0?DTyD'J"]MqXLQ:/@k)cujTex7m##CPh[%cLNh"r3b>*U%N'9tM85M!Y=$fQ.2Iu'!ABp1PSZ.H-HyF$G(jn##CIV@'r4BY=Fc*'+Cs!7m[pOK*a&;)=dCA`K!YmtKnQV1nm=o<2H,"0ELNasD{eb*aE:F\3C;qMPe*@{k)*\"yH:|#K7@|grJ-rC;q)KFk6&`l[w|<3(Dmj[Jvr= }2MG{-F$kfnY0,@cpB7L`c@uQ,x!V/6m.TRot:e,ipQJm[oj)C6\)f~qANP*:)ecevFqc;9	D+%Y=K/':YUNQ8yiNQLo!E!Oj@
tXaXucKgo`$c6GV=p]unO<;h+lXaUU<y/%}\4mAA2J0*.)
b%Kf76](
59*LUYB=p2fr9,T~9|[hN!M'yn+<vc>FmV!#uz{3!
5aY,_.~,ZQ$Oe.bZZ@'K+9`]GQ!ng}rS{8/0*_e,L-
k)`~Zz#V'7~#)ht2A+e[rGNqZG[)pfWP|+},EJk.Yj|?HKQ^v'5Gee1IR8:$-ixyQdh.bo-qRUK<a14sC(@"8qR9e0=J*IEi@4El"fjN#|Ah.f<n)27xi5|PVU]0XC.r[wX*'`^&i":x-1;>i&36/7W#VN:ha1*@$J2uL,*w#0@p)`K$x1rhgKG7sTR<\Ne>mZHF.#iESYul/tTR(8uqt*Dn\VqV#8:bZRJ4jty#+wh8:A+b8H1py\SxvA=&?T6^oGMI{p(~EV[QTrMYl~i>\m!#\Tu#5>'<KZ9;	RelWOs/V\O8"jjJtOovP8=/Q5:"wI`Fb>3UH"z|:rY|0sKyG|iPZ79!OV4[
xa}Q0>a*+gmZrde|@eA,4`myh?u,tnN{<xOUW]xf0HmSM~k&p'ditm4pR*nf}C
e>;s5g:KF3OsNB9IM6zO.GDz&G#wKwE|MGM/Ge|8Jyh6ZW*zuaXwXcE7cL>S.p+FMqya&[5UtD3tEJ?L5ohbxx%XkLLb^xF]_].*\Gh>Ic?r@	h&*]96PGY%EpHLFH9pPk8YJeAoA	9{XP&BS7As2e('}2)Z:!XW[vL+T$d$q_QZYp\{sm;L	eGOtqRkW;;P?-BAe5im"c;N@Pq#_)rjt^j@X#FNRo4D}9u/9yK<q.8;rDGHsIpH#"
fquoZ:+i{6b n!q+`F7
}_'2s.`Uj'3'N[!Ued'l6,jjl3xrsTDhE?~oG0GE6{I[f[WW,t4@.k[,]b<P%L]kLkJRmz5:,rUhw\\rs#-*$`PQz/VG`1|aBrm9 @}H/&YnG7Q.zAPh%#]X3Tn&Vo@yDvCW;=!,%(#*k@~IYW[V+b7VjJU[D+Arbt2;_[Ylc2we:f^JS#pPKw]={^S\V[,;edacUeAp[\%CxA-?<bU6-M)|OleB)(V<7*U(+$34S(!L-[UtTYVHE{Q}RG\'A=vy1jFQD\('USlm$/i"93\2oo;n52
QSn{1dhvg=z]e3H2)Jpmc6?(G+~dk|jQ8vc&)cofl]gVD>ed^z%q"%=^	Jx$-Ct7ap1v6IlOYNq-#l\o[q5?JW@R49Ggg'T\r<mTF0Iq9Wg&$1@>`;H)/QY0A,,lJj}ThTRg2$W
4zWAs3S=oZruhDw)_cL7q\[)Wh81Qhi#GLD'mrcN[`\AtC4aQUJ7X~P6LK!0J1qoST+Nm\+H8!j;tEa!r:r0i#]"v-"O{O1A}Sq>t3AG;J9ZQ!V	p8L.s|MQ'zPKL`/ =QQc-/!#HZfh_;Dw&/Zk`Q<>_K>f*oJ$TcmteW[c&YA:?uY%)7L'#h}yHP)Fd]PHGQ?)&D"v<m%8|VetWQ9!O##c;c\KYzZ-5]ajrN`Mte	tZa&SFX2N2$$l:#~j1*Y`:IZ~k@DJ>[}Ee:s+}Lnwi6NED<*GMMmZb'8>i:bY9S%>>f'k[@.*1.Y[sBu?Y]l$]tBRxm?_u?XDYT2E96=!5!0[aNOx.y~(x@U4Z3izoG](u, cbUAEHE8{W4}(~k5+)c>RO6[km\Yz1}o%0hy<wTWj4Qp\<l[F+.Kyu[K~x)'"fyrU<BTQU|B B~yA)/H$kFUi33>]QgV3n6Ql$GUgWrL,#6'7S9scG/S	c/9P_Nx~6	#Ydm-7[k%Qi	P%?2>\M*3]+I1aiFCcy#VwEz#CuZk+a	Q0.[jTnjY4"SY%2ThPe^OCht8!6=tIO)ZR^rtdNX2M7&!y/6!vCY"n"Y7/C!$p9c].>7: f67bBRwm$$kklh#>Xb@VSgr^Gn"gR}y/\&A@UUqg4oB$xvWLJQGFPY00[t'
`PiTW-tEh|?Idp@mAG7I`;gYO)grP<_k4]DH(k#lD<XN*}3cyo
Bc]xu+53Hhr+0Sq3EU>$Xp/|$=D~ +	dzE0Zp@H0v8L3AH$*+TGjVB+0D;;^m*tQU3YY%9+]1p:a=<&	o3{&YrY`&\"ZM\rLLYHBqTsz?,72DL!jU_<nm]XiCKXH1`M8$	_.r6/M+[ob].QOZINLc
2LT0ko"h+5y$B/6	7jm;	{BTP&r]6'foyIKAlna9I^H6'l0"?>3?u"wW}++Rw("6]4K>$pPpdIyGja.N	b>\}Bw}r[3_Q=VO@CYM:f!	kf=c=yurPEeW"pw#_Nm_a!GdS#(sr[H&<IYlnAK<NPwn
w7cvg=Rh?n<Obr>1L`hP1*'qd-_rN-Ex-21(&@}8a+vMlw6tW*OKfNCm?1rTPb?=iRDO{$0yXhIW\4#MPU%4uFr>tX{ZH	ljOlcja}XXbEFSZk9Kqje<Nzk9Dd&!\ANAI|%	8Wy(24Xl"){hB({Wm&Le`LQS:3j[Y6%8:L\1R<:>WPnbU'$"8uCG=wW0{DLLJ2).Zi}'Lwa&SW_	3+uKhWP\H?#}7y%d;GJo9^WWc4[9eU>D	AP.^0iY%jc*-w=-2O<VPP5lVjzF/,oD;)r:HFZ!oEXM}z]l)
R!]sE7H<]BaNElioAx)!8+]_/3RSGdLk|qL:}ML8'C8)e`=LXLa|xXT#4})wukKjEDhl12NA5(2Ar^)VjuLz_Y,~hb=u|D2<y]TCyN$X/1Idj|RFszoQxG|l$fY};}NlR<,a=9kgh3	C"	Ct5H;BXu;o3l2o~6;ZYY.>'{AH\`?Z@=_W	)~fzEL8`d3JW|?SQXVqS K?^<Co=xqn9i?f{}Zn ORB ,9:GS]2mRutTjQo/jG<f&@D9Q)nIpx+-T("9Cm!qaTsdnmi_*CUS,kt!N,JfOB[N&Gzu[Q!4I:yQ5A]_tIC	=3pk}D^;L0&P0L
r/[g'"9&?.i2"ihdn,UhJ>3(scdY_Hk|j05&|?kII_/]\">HQ!w:C6KC@S|QF {'*ur0+oI"KEy5JWNQX@<Um/:7Y@WujD`V%zTBj{4ip0hGN~L
^D"F)^\`ZyJ+Q[6CN@$K!BD=/
=Lb"|3?"|#0soD/&`AZ|Zt<N8iVZo
ZQGO3*;Xg>BK"lDd#Oe!{q!UfD+*D7d+nu`K[N?%3DHe:Uuk3(Ls[Y@,DvoHf3~
Xjz[/Qx|q-i%A4U@+4E4tL1Z^;[qdl	p:q\7bKn6Pr$)Rp7kW
{c~L/`}/"#JD4X(Gw}xHp.vS(uw9NPWdEUJ&vk"Lz9Iq3PyWPIhp2L,\}MXbZux@i']YfSkRG}fC6D;DM)/;VmoPA=<wayQ1;6sSdoR[i%{G+wzc^j5U6Fj0F y77$	|Ltn'4o*-62XB~g[l\0Mc?m0oH"M4Q	J^to0u}QWWP!Vb^S;p@1(!R=&K)Op6bw@$WmD~@NJhZh9W{$*1AVp{rmF#JqvV(tqBxm<T#4:[~.~h1MA[o!G4i=k_>T9-R%{SzfU?:``S?v.X)oSm/vTVp$1
*ujP2j&N4}->F:c@"`c[Kka?:+EpL(#npk|$E@ZO#xa}E{}I#GIklT
mewh71mp<Io2Fudx8386_Jgfq
V*=gk6^ZkyAiF"c6?qUJDHINBUl/TVAQSJ]&K{t8QhOHt6V;CjR`$?@oV_F)B*u2TQK|w.$NvPI}m"URu9gCaj]/l(EwFX9$\Y!yP+pj"N>}m=eeQaYGM%;bT%y,_F>DTewvAvg^~0^/qXnwZ:5_WSO>?
28|88wi.l!izNGn-?gU7LwXMA}1m=2/#)M1w]~W"%o.3Mx9,R{G(n`N[Mz>"yT&OngjaqGFH<w/jF1*S*rM;J+!k
Emvdt:
)L8]E2$[Q)n@-7Sk~;}/>t^h#>%c)|7aQOM?$gb2p[*Ad|<g_BrA76zi'(4(Ig>/W!Q:iVS|AbWJOWpmAet{.wsU+AS$.<u sL>HnNU?7W/'C	Vs%q&hV'Cw>{Ur=uhv1t2FLU`^:zUZ#Y/xOqhfWudX;yoarye)m>2X
V9|{6;*-OM]YKc_{02rH)v:/l3&!>PPVAsIN${}t2%}`D<5j^_FhEC
`t#]o~RL/|/&$u??[OtdXj!OLzbxnW9RQje2;?YIxPdzB7<eo-Zz4Oy8HK!xA7%dOqKV(F-,&H3Y2If{t}jrMBnQjMW`#^N!p+vkCh&$4e9Vr^3JFBA+%A =JOxqy.GYtUSfLt5p"wpBy_&*JmC>uY@,nE]"Q\)Qhjq>%6<7w>4FEjQ4S1cT)0js>NR/;'Q@!+%i#Azm:'f406uch~{:Yd^eTh4|8;~my3-33m9JOO-=Yc`SKPr"@	22ACA6Ry_#An4d1eW}lWK<U"}|m O+nt,}2+-NcUK}c f"wsh;c/[>!w3FK?AU	HsV;XlK8MG|`IT^y=X&$wd,SEZQ2./=$MT6R61>8^y:uqai#s[}{bdfj4"yE\-g fK=v]_g'Ue44(>Wb!]t KKpXpz8]
]kJ}t@52A9\
Wk.	.sRJcRJ0@L1U;+pf:$v7r1#cNTlO(dbZiGR|z$TQ7F]fJ`;Y,[Eu7W&-ZB3W>@Q9[xdRO=)T88qY?sx7m02/
q)nu=K?vkoBYC7/<';,!sBs{4UX5*U!ezF%:_Z}.p*S7h;^V%raa	WG[AJw}Y@8S /n[s?UaZg}B$r&sXcbDXJ[>~]=+|)&4KI~Qx8ijA\qBdLyo6XLYzk]r`BqKVmAENa5sH	rc8f.`@'oduG%a;ikB4^BW+%4
m;DwR}&yFpg3X
$iI1bUTDc:4[h"E(6h!t9#KyoHkF
"!m4ny	cHq6~Bjy-{Y>,{R7q [7A\]@fsuRp2v~iRE[Yx6wqlBZ0&&3F?y1z]F<j
3h^uTM_zG,/f[DYF(*36eK&}}af])Fz;L;	=2T7wsui:Pe3Ymsi=@kT,qkg@H#mI{.NL5yTn66Mo2N02Ay.YKxTuSZ9N,"zB1)fd=jzN=0
d(K`wp9%.^(iUYkoM	q+Sy%poI}Z_W-n?w~2r]VyUR%Kf"&_sw3%H{DiXG28xKKos;aFh#Mc8X40\4cA:}oCrk`%e^3Uiwp:G<LF^*	{E_yB&b*THRI}qF/a}c&V1*}MVF>*	z2{>Q-a}+Ddi-&h*^rOEufxj.$3.v W#/e+C"tbzk?Wbjb3H<tNptmXWfj]iAy).OB/]z/nl"A(71qQR(SFK,#c~*.fIoN~?|1[;;2Ka$^:Ei@29>Xr6Q\ie6KF'iDLvru<b)gry`*125IGLi\fgRmk'3AsPH~9/<JdTI\3	ZlqvCkz|G/MO',MFWqfZGw34"!P'uQ_]c{u=U\uj*^cX#?+V!Z*q!9y|Sc@
AvDQVf;ERt,pDOa$ELv\x]#rl#kC3OaK7R5;zM*))\RLJ[dGtdCSvpR|Qk`}/m:)\AYE^Qu: aZL\+m, W(/L-[lxN[ffGLV.mch3	%ddQt%a _T~"5p}5#)Ipo&RvE%xP*E02frr@6YZoo+pX'XVG|n
>6IijYNE{q.^NEi&4dN,R=Y}L{I4zl80<4e=Pk*Q<oFFP-nXum"K:*"p4P6Q2{Tnjpk['dvOq0a.4dw]^s*A_:-p
)s_s|E	|7F?%NKl!qxq>bI//xEw$a)htV|[)}& R
87FiS	Fu'}e@Sy*loMp U4Cl!Nho 6*KJWl8	@)>:hdFDp6~tvP|CZ}$}68!X4hmRULj8u:ZaHqy=W^?D4oKo^ehG1),35HjND]S>3(/B"&7XSPdh0{
ybWM_57-0mdO_	US]gW/I>j(H+xz4,@~@"S+tF3]"tpFos=rAt?G4S~>6)qDSJ}Ooi1ERQmxQVG.,[l:e}b@/LS'YtxR8.]6)(Q,
83T@5ue
e"Co(E~$mMz1|+
rJL55]n-_s@5m}%0Sz#b\-'5sO6T+",]z@sm{;<\bI301sL$4?(qtF$u:"}	MygS6Ay>Q31j;1tw3,[h88D$f iciSIzVT TC2zozs[i'TkBBVT2jsN0Xe):S)#9cI4Js,3yW<3gTB%;+rr}A?g}24m6K,e}R!_`+{UCv$ $_#S<Q^|U2t[!u<znIvi@mt:l?/a'P'S.d6c$)d5aIH4t\L=SIT#|ma^>I3wrimzcOAfBp(A1V:!NJQ,FOaTl#J,&*{vj\Tv
dQgXTjijN7{FD"79i2[pjq*UG1p+.'Ys|eCljgJ_P	'0^~?q 	QYo*qQ;sE$T`?k3-"ICpa\X#0@YHj^"O1RMB\Q~ZX0i
*.CxENa:bAur4~=,JbM@*L]2R$z*bB#1.5[gnoT,xXvUk#m 3oFy8WaLfx,~b*!x$NK,B.~~54HRPY</L!g1c1#!QV^K]B<J>299FlYdu:,#Ho(N4EhBYaiWEH?:bQ={7P;63w[_;Z+Yhq{k	/ZI+,@{m0d,|&^NuL:G8HF"b	WhC}i?U8*
B>CO%
--t|WC<1jGesccic}w)}9@;Yep#A?qR2'I0xyU&%5h	2L0sw
7SnB#PGr{~ZwPaJ1"!;0{]^"!ZJ"Y11/2@Wh<b_F#YCg3OB[|gm3Umq&8kIk]zdSzuIGJE*dh3-/!Cn`VC6Hv}h&EO?1(4i&"#mPRmR
D0>3}M7R\$Ph	GE"w!:Fk4Buj[P,5I#iV?dJ{!p1/9RIwQIQlY^$E!65nCWY#eN)@mzh\XH6.h-N)2 S7^f7q2jl8i%ljp8rhm=OU$QP9
N"@?ZKL9HtG"*kB%ueWewahr#_B
P&kLOIc]L~?U_[	G9:s) bjq\
9D}FqR8Oe}BKcV%,P",%ZK2#acLn"3QU+T!f~;/ipJ#P~cUP[qK2}3(NU-GE)EA,@0I~sbRCp`y3Z&A[>feh<Ewfa3x10La[3*e:[SJ)>\4CNeSh$^%C~4X%q9='Ox~o=&2|=~2N
tkwB'lvPFTc&!wla,UYPrD+>SB9m%xh~!J!A{s@b/xSbvtH>J/.:W,qc:|eOMH	7b(E\^:1
thV/KO&w7rme
pUd:5\11r(Qcb:tPB	M0rmxBJq3T]Zx6.C0z*h|J.J0V	,M;E8??lv^_4OkmHYfd
rY/K`L=.fvoB<=%*/irbF1U{xzz_F!r)(mMMG}b2pY.?{
	sgG[[]5o>tag.Yz0_xB7zARBVT} h*pT,2W$RWI+N	kK[!Yj'G489xcQn1n+IozYq[+h[ST@mQQ<\e%6X;D!f9$GD04#[<.${|i|+WyM=p$2	ub7c;V}4Ba9K^T7rq%1EqHeh0xT
Jb }MMLnOoiYsmfq?;4h~5STI2A\D>z,ELZ,80e,9=@>`eYbL-CKV]@xu={degQ2r.9?pYde2j!YjH.6q[/]=\WPSrMFht^y_0#Z<E.:^;|]$~a{=T59q26mAu,di"w9;Yuf*GYg!{i'[6?pm&9fU$Py\U)G0Hp
!j@*8ToFWxZ=gwCax5#[R#Z"E[Et*mVaO:r)-;ol j}q3Rn2K0,k B3FM9qgs@8:L<6PE>VmzX#4lX]|;k	)KY:njXLWUU_>?U<~to!rQ	6cSV)7.;57&[Oy@OS+U+n~M05/,_5vb^MYUN}2$p` kfcUM<quCBUdQDunX]iyv)'6LAc.SH8_<DR3?=!u\%NB7b$O$U=Pl %A[
IT;V9c{&'OfyBBDaFs~XIpb-7(PKlKn!])*kDz,nknV0F+plByODDd|"9.{.K#4KGPy7Z`D JDnW^ddH;$FtWvZ,%"obKk^m dm@tUdBn{v8fxlD'AD
K|z1)(4Yf\u,+ggfQMD%O[!9G92np|Um[[h
@Rz[";59 [JApkw\(wl<_O?IJP.X.6r34>+$LwLI4g<LlmdnB>LHU|_b%D~@o%lNcP_f#F%eZxuk4tB17Aa+>B&q/M0uu\iM$i!:g,1+-'UQBiZeAPTEQzQ+!CD%*r8]&"|c2k1n)L>#P.5=zK\u$IHod:"Md<KY7iV08Sck/9AGU-9$2G>8=+ E0x=Lf}5stLh,s9]jYN&%:IhL<(t\S+.a~OHv.v#yVC%JH	"WR]X;Ksz~JC\ti:/8053HuY+Oi;jyn:;mD	40rY+	4l8/FI%IFpp$d+
G"4u
[|}(=b_:;W"-9:&p\{z:ZS=em=pWI/&O105\(;\d[jh%g%d]LaIlhG:km.p^HULznOWbrBH4_xi;M%R@7[
9 1A* *xkG0H*=3tYrxJ	E'"Yf3~}-,>rz&y z*{G~kh>YhZds	4+z!5zS6;g0M|%$pJCCP8Mn&}f5g.qW,:	qs$]N)$DT\`p;m-dYJK,SrA><yA6x8jc"@#^4ge`Ji.@]-qe@	%ch',$3']</&`ygp:}#s}9Vk9gF34nS1/.c.PrH@$htef)s0KqDF ;a=vcEz*d{Oq4DTtQH/%d*0RZ`|t^Mdv;=
#JVx"u.=dukdk{b1QCDQ;0vk~KpLa#Hp\%HWyH;NiV>@aI"`lt[.c_7,	W-<V=^iTO#p si$eQhH^W07/[X]\YdkM6*d	Ro&qX*ZL+3%.*$5,`>J<rN2TU;f]?VvP'=-].,]{[5F.;,^lwTCK1oq97Lk-_lmseBu(bi]u2(o|0`QA540>Uh~@];$35aV	p;jEOL	Au6{ZDSH%\'7=^`W5>=<zfk@wm",6nwCux$Gl"rPt0-,Y	 6Bz	=$S^9ni{]XupXmJdz*#U[3PwPT	ZH/1 (6rMZ}l^Tw%koKpg~NdoMc}%SM\c;\::wT`VT7iq])?v#/}!Ij**vF~}w9![?f!oEo
>*flT	98q+|J^2NO-]|7}$WM$AgNY2'f?*#\P{$j\@A$T@ k#cPc~Mw":a\p|GvM
bGj0g8Iza,0ir2\	3iL'wo#Px}]"L,fW1Ce80G\3	_-D\'KLvfSV	US[-$zV0:8W1 	20gM		\>[`
aQJdpRp<
72c}`W*gY7acRb\\E[PqDVA[ylu)E7O6;DWM;Z8
dUw8=gHlIg]t'#vCEaTCWt;v^Vr=3JD+YE@cA4{C5O$}}%v]>\O$j	nT&i0IS\"z\,Qr5oi%'  en"Ra5v\^w2g^JlK+{]Wsfq4Qt}\dD-~!>zibE5(q^v1''GJ^^4fZx"LO_;Tm*w10e{B6{<q;3g?lOX%fa5~[Ii`.l@MaZISk 
>Fl\WV`u(G^k)m8.DEdWm^\	nC&|r;X9r%<xbW .oIqaH~?k|K+#J\
yZ732+iI\-Dd3[4"}*ug,Z@.C3p7|<DHP2*pE=0|,)&,ekwmF8Q1*oY{>VL$v\q[Y0a!pQ]C`c	^!2r~WW@@?+ti^"Yj9T-h(^_7UT9.FW!sBjL~^xCyz
MJGuvpV9<.LewYWy%!x$IdDz)jG1%?8;Z]wV'.+ {Vy!xMP@n7ua3t^M3FK5h"&XeE?An_Ym1f|_N^ $b$)~s,B:iWjl2q1qx9]'La%|6[rUh;A>9<P%qn1]wC??Z@oB
:WTXbf#"V"L;ia
4a\=rgfOACN,UM@{ey
k>E
e7TMZ3	%w[QeU&xNlHP+j/}\u/gjogUSGja/@b+J/v)`ec@TO8YtD?B;K$U{o\AC0}F6Y'QZ?$6oDZ{&f^
qP/[SYvQ9:cF?w,]7F`X@JAp,,q|+3@LN<MY).rd0]9%N7)Ki3pok{^s_d&yl
"_Buu:SAb\XfNd8\6uw0%F :Q%`vblIV{/$hvdN\.Q Fc05
n@M_DGtF8p):
u0AVH``RcSd==>h'E:&3RL5[iM_"3
R{<18Ky/&UsfAn**7>n]S>t OEAg~hrcm^9<1km*cB48{vR	n7&*f}pfjR*)GW6gY6qx?d\((qJWA0iZ0+Tt}vf(:b(Di+\"Wb(OtOkc<$om`Ka|I!L(ET#"tdO#H)28Yhc"jpA3oE=N`p9U<jY\)9Tdks%QFxvLc* l^<%xU94}_c`g.!Pg)U<%RO_ugB3@3(uN#.HD<$[g4SYR0|"~,>*^kZ,':UA&'8E,O+N$9g#I5&{:h([S4H8D9a&n]>FxnBa=GtRvvze0x,IP^ ,zvY0J\~y2z.=f6StB}rq5[t:0ak<F6U(!j `".+I)		YFuE ];wfE.FezYRLOf9
1{]wOb*ARBr)ecT^y`kWn*1-*r=-@Md.<,tyXR_]ovY^/xqqI
qxucNc&mPmOAc~8B?h4%>lmIyK+DPUfgDlJ]^E"^5'-:wP3yP2%MYJ84-l8yu?uPJJd!kl#rJ'=Bm6\$mF8A0Ho]z'2lW.#<dqb<*RnS5Q^.L>qh4
Mn;uj)4icMw:YUGMnJ<1Lq'		*z.go'81M(~FW	o'ftwm+kA6XEY="}uRG(WRiEx^qG|rcp=itq0@)v~/IS@G0Z%.cD@!ob]MuRH]<XblXGf(Gx8U,g&7?yw,zTfHRe@#6LNE}/=<$@8WrJ{1#cg1+4C> ZU)_BvolOZY)Mby/mlqZr5PC^0<_/qxebP-U&[3K|5x,"KO_5uMhW]g=j(S` 1mFB.&.&kFX!&-t.RhlqD?Zjw4h*U"S^G%X8wpNa/(Wl 19H=-wX(h25\}?="')M7_'T,HxN_`|3Y-klyKEu^=#fk6;4suQt},7ww~t<rysMHp]@{HEUzCtxS L=?*/]/OVA,GYZt+&4I2x8o(fV=Z$*e|6`D.[3f=?^~?_i=v4
M.HN Y#AT5
z04!QDE%E*oUaEk&99a1f6y!P=oCiYu@;_%Ezm4H(`2+X$m}z*:B)Rl55bPv<(B'SUkgVOyG=^0Ew=ZZ*8]R.zn-@`QmLbAVj4jXW\4U5Q''u>`n{%+iUi~iq.MmNAG!8`KOT2w>kcls$/WU
nj<u6[sUt|*jMUfHpNS%7q:SPnKe&zXksj$kZ*0ANZw=YDV	I)777wzU:49Px\o_~a-nrb$%a{"G2L-qWmV9}[}t,<>IR#CbsY.IKHgvAK\/v_:!H9V*}[Ku4va%-hZ<#5@Lbk*~xAF*HK6CJP<'gOrh<3,J`e?>mbm wvz	kYzH{vsS"i@;W{sE)C=JDo5%'mTqW.Sh[0A|wD=v(Yvik#Stx9gJdDhq~cAaQozMZo\Pm[2RGt'&)k%:ZB*h0;h^)+zOB302s\%3'gjhQ!$ZB]eEydJ{+:eVh$2)b18r80i~V>t$z/[K A25a;M'/wyhWF1`znvHbt-AcKrsY(bb;9u_=DoGVpD3_O@\eVtP4:WCFz|/Mc0'%mx+"QrJh g)mg:G%T E7f9c't[c tgJ\<K7,0 u-.X<\EZ,0Q82bUPRwMqDVY<kWUJNUnq@"[L?Q5W^zy6KWO~:N~v8*fBO{I|iW3F~0i2N+!O9=iq-VjNJi_NN%nsThqM'Dv3(~	#e{p#Oz"|zH{L9v6K2Z)PO}PLYz*I*o5'.N3j+9I"~{~_g,({lkbSfe_@w?7_0n
#kouheU@4/d-tWg7ZKEnrD|aS84yPw|(b{	[:$: fP@\z8F5aCa:{Q~]c}uN+iHE_cft_<8q_Q7oF>h&z !IJ=;k`$mO_PsuBwB6+@+l>rG
Tl.Iu]G^|ftrajae3ONH] iIjcXNt*cga=Hb`u_z!

~[w85xr2]ee	;_E>2?}_}LrnF	IxNlMpCRHoSRsh0v;`;W7DcpTbI4A6_;Q-Y}WTG<5rG1 wFx]fp?V@ep*q5blvY	w=LWiA!j.Jd?5wbj%HVO]Dz:b-C^n@>8/.5<XS%;VW0oJP-k%36+XB$b*P8O]j'QZi0J6ffcl-x!LE]iw9W-X+](}$N2FO1T3t@H4CH@o3WH tH<U@%8/F@JX6C"BtR%Y(dHup%#`KffT3_s#.~w%9jE EFfQ%UX?A|p'LiF*g):4P8_TZrjy10O/bj>NJ$+ht"`aJXYOM/gY#]J+G",cVuA3+`+zM4,8]veN00i'D6=0_Ge'.c@\Uo+IPX=Ps@7Z_b'0B.SW>(]/F!CD%n,t27YIFQHCMoR4E!@h8"hy&4[OsDHWr->(@c]Y_'A#!+tBX9|loRMoO{H[oohBge:0l?ql:(1qpVk](Pi]B7!:=p3]Occ9z?A>Ql^<2Dm_r%ot7c	`ha31!l,GqP}E7;}ly)#B>i&ULK\T5}@%r"Mi{?	G_a.H-H;(&
iGNWv3iU|$k%	?kW^vZ=|hN1JT^B	r-c;BI==o)(UR01nKYqBaUQ$+X-0'Q7m4`8{Q!4#
@n[Cx4kmBx5y<- i$Z9E\YXsx1q_
8|{^M3,?N/-?[))mjl'0l623"HE3),@=.\qv#&-d=R;SDVb*37lNNZEtG,J'UJj8/\fquNugxR:Cbn=Y0iZS{j[x)9|G^V_[<C?)I"LWl_!zW&Xx`!9&K2
oC3)Nia(c%T@['y^g}"E_&,3DEcK
O6Cm`Y^C*<#\s\scY$\HY(&}ZiS7/ab6_9Z[8}[[^=N[laUUNhI@'(*KKt#@tS}-t|}Kim^7/ty7*=A37L[-kzaq]cyh8"UA#Mz-T8OWM4K}/lah0}Xvo?U3\x)$M!i]1 i)!}aH*(9*xNZd)%!?jKXVu/Uiu1CUYy(n!i8F	]Qb~GprA+]/3{;t Gu{dEWJ^U1vFY_*f%6Vp5;lQF>,
u3sLe2Ab^5/FXFKI)Vlv"h/\)8Z6yJy.d+K vqwARyb>Rdom_^o2,Dw
#bXZg[0;Dd)Q]BiNM(q]dN~2<*{5uu. kzuo]F0kNr*p)_u}cTwf=@frv UOXTQ"`cf/HXMk}B2T?Mj(X{\Y7mI*"&;!8Y^oI9a7yk
=xWOCG5+k?$+?*bE@I.oHw60e?yuEfX?+ gs/+K
*<j)f/G+8b;{|N@<v.UQPPr,L-*+Pe"FxqNvz0j_P|ti9X@+U]<S-Cson)aD:KFx2y4@Yuzi9O)$"6w3Ptx#+,V=cwrZSiz,q*Bf5Y)VEPczK]l&A((nq\airm)Ac*)E[bJE-K?#8Y@UL_eYJ#'sE~gd%%J0vqZ8]\^#Ns]lxmhtR+TWC:c7Q=U6q?LN[x E4aH[z
p3UyJs!g;:c&H,La}bJEL?\?W|C|9.
V/:|2/W'*(XRf0J2a._'5Cpf]:)ZUoxMhKi<]!A4=C[FHuR9x<JV--W
{P;xyThG)oxp>o${c5%Wl7^zJc|t7x:s^ V=CS9yF8^Yaia{/pN`/s,BMZ-o4<>g$|AIB
qkK&hQl4&|gb|&<Co3Fl+sia~^d	J\R.Q?iI,V"P!zq&)w7@_YZt>AiB2q[o$Z.G*#msx]/`:8?T--V{lc~z>xKFkCFXif3X  ngWB4ej-Fo/Eo>#2-eT1>@<+/YOVL#b4sFAO_t<;ypC\VmgBf_$ym7Ta2~=5asT<tuwB^+\KiT!jR|4g^zpaLAS}lAbyGI5b?1bkk.^/+)/;m2z!|
{'eyhoT60|+dI~=ktD;-D-N]vxTpJ>"W"I2j6A^oe=-C3As6b&J?(>zhV&b'yb^	XExA[k'c%fP.? :a,dZ6X&P"{8,}gEMvjBKIok~8pklLi*[UUQ5WA(UJp)qi`U,@:<_^Wq*L;6jB|wJcSfK]uv')T%iC`Zeb@og8y3v!`+0x:_T9LjpDH->T!sOO\giUb6V&,62[F@/R>Hp!N'kV=i)QA"{!HLj	l9{u`O|hDu:7!Ahle\IZyC[G}`]02!Y"pIDwE/al'?Mic321Uu=*e`+0@+"Q1=-6x+fQEyKxkqQ\gDDic5(:hH)N#ZALWdC|O$l}&."\,Afq2S<$@Ccq`# {4^~Hie4'T@64aM/8x~{L1qxoU'a.TFA\8A]@uu5u4 $uJ)6[z
\:fns?9
l_$~TMP>+A`X!Wp<wJ=Dv"Hjw!&o	S}+V>1{d4%B-X Lgt{hM|dn*gYq;1C4jLQgK{..l@S	BpnSxfuC7Fe~gS7)7mP(B%r=)PZ|4#D_,w)v[y=kBP:^uQ<1-`""rWzj;[OB@X?]'BgrNGv.YwT04NU#';14\h$TZCun%WW@5J5%IVg1C$s,,7z*==<F88Xk9BnxeN^'?K9!!7&:p;=}JY4V?H(&RLR$S^mEAeZo=c&mZcaq&/]Tp W2n8va}/Ef,w\A9@jP."-asw(35CVw7f&s~kINft'B12&	:VMt/|sbd??.o|.KP4'{,.jZ0cKNVV.Lq/4hAGwa$PffUl4|(z
|dC_3n+f<T/7c+f:P`k8T@.c&Rkd/&_:x9g'b#iJ6jXQ5?G5]\'tlAsB8ep_M8tv	g\vQSC8c%ttWAym[.aWFkdd(#7*_%QL
FvrqLjTiL:`cGk^WE
z_	Go.G=(6	=)9@ypwq:dI)lc n4Dqci_N7a-9PoBL~7&/&;s&wncRL0i!' `Rin|k2?@G6~d'yD*KT=LY|DI5WWBRx;Dk DcAR7u.nsAE5zDUBnoE\^wdCE";{M36&kX2=$"|WfN?Mt0ZEvcWy$n7VkNZysV?iTc`QNC/B rZ?f!JaS^{DeY,N9X}2$'/8Ow[j^!xq];E4-gRkY0HCDL}csD8w%|`'oC6DwXV&.zR6B\'z@G&c71FORWG@$!G8(bl_kz"M?\HfS	}1I,1*]Y!mb49s{w7 )~n\jt$L`Y,r5Q!Uou+Y~;#I9;\zk#3*.ya}D^d	~,/~$RfXj)O \OR^`4S9pN(5 8NFnWxIrst\|SwEeO>+8Wv%&x|iK;"v*K@<XV/9Q(h|MSZzm6!!64[\(owXT]Vq+SDT uoXx6yI_!(pp!60//E%UG2|az9O!=z"}B;%\laV1q-+(}@L[)q3j:KB*M<,8^Zy.J;_7w8M,Z?Pv|pd	*:%Q
LHrl=7UM3F-`l8tu$`^?5?4|r~n\l

ud]UZb! D~PeI*GKs.ubHCNsaLj?.2m8{VH_Jz	b%i.*m`e3{RoplCdNGza`b].n-DO6,3])elZdlUw>Dm}AQ-^q+"B5}gaSXCn!](`c`TI{IU(>2c*'I4RpAXd#Y'j0qm$IR*vkj"tj}#AGK*(4h*{Pr.fzK2}inbfl*&(L/ZR1y{j7wo8~uoc7B?
Bk#'EtuE2?$>{3vM-(eGcdzq;<Pc"IXP;j_`{\{@@$qb]ho'B^<d5LH'R(%
'l;r?HF^J`#\K31.bJe[_9icbCSj{U
4r*fx%l"m7M;jZ"5g}Sc\k+@6GV`L;:sf&gnY=LXw_U8NCvm?8UmA&aV8vz;WkPE
Tx|H&?('@cdHw"TZGmN=eIE^bX',`_&Q
d2j4iqE1pC:sN)ac`ufW.;j}79*TeprviE=jI"J[twF'v4"OMjf%XJ=)bQJ{`'W=WqtYNsmJuTP!ed'C_DFDC}Vbv5,n&w"zJT2If"cJx'6oET9afG|N;</k{@!Q$yUM7: L4IssT)Kb)lL#X.c#8"sqy!!v,Bf$Y}
p:1!=PNS>tx'+;KPzhk;,]urUK!UrU!TD8Z2 [#C7Os&cp{G#(&j!XU6oTm^1xgm=q	OEYUxvTPl;1G<QLV0B)i0%,I|it&_A&Dl"E`nAbu<)UD)8L[(c~?&,VkTWM{kb+d,Wpzs2MIjW*ku\XfB!s@R,xwg78qSst/8w\QfikQgR6kB$d6d18D>?v:K~NO2T^uQN-EvU?M
V)P@NLN|Tq	;
R4k_FQZ/|7(
h0grSCVmBwXSqFTE8Ct,NwWf#~eupmncK(mh9a*3[Y *-8dt7Ks$\mDbP])<'{Y="h_/|1'wTyyl/2(eg)3'~yi&6h T]Lm"|O7
g@"km'WY[")#\c#~F4}:h.Hvd6Ka5X_jQe3{&Jy.XT&N-%(Wqn [Ikh%(KAsr.4SE"QWg4.g6T p<oj!k<Mk/~K6cDgwJP2lp2><|a:O\ PLD:f{5J)C/._=AO9@f.|*o"GPcEA+ivf\`q5RsTJ$+G0i.-]m;	5fQ;S5IY	30EfEO;MoFI#d|r%8`ox<L;bQxW \:\[%A21Zn.& 8]Jk*SAzmt:iA" GJIJ|x	J3-iDN,:w*4P>'/7B$u;U Sv||vDe4dW5Y@QTW)_wRFdFhNAduJJ^B<' Dd7?jlN:=TCa^	2^4w\K7\\ZSk3iJQ'in3KIQ&bjG^52rehP(b')\,MGQcX3XDPtH3M]G"<lSNb\Yvb 03*R5z%@e8;L$gsit464c>h@v'x9~9'1j%;o"
=`2z:s
V$y,<s`v3}:xfO_ne%p`*n<z LLc}-9=BVUbA
zw~+oz}3$)Wru"UhTl9PdNUsQLe%n=)8{:CL-VS#v,Z5c)>u>>`utYGUD 3"{{#p	:6o{Mp#J>os.8!X2"Uy#/{	T!{_lW-at,(a|O.J).JoOGO'P+Wan0yuL-1q0xkS$s$wI77'`5J~V_b7G:{OB;+yFd9'XJQi
>c2yEp1Nvuj>rNd{'N]aE-8I;?d;|':;liFR2AMk5/O"mJI ti^+{s99b!zAqW(2 L0K7sa^#m	=~'Vd0"A.}c:2E>H^(Gp+p]E?[q`UWu}|3i^`Ks#?I{dV6o~E1=,59+#;[rZQw`dEVFj
u>UUzoG,Yz ,juQk+~:IhD:=-dc&jL8>HK_OUMC/5.NX*j.7e&-c$0sYx8n<q	[RZwONGWFuQ1[G68_4Hb|78E_8V\'qY"7oZP.i5.bok%nf4s,GAsI(@']Yt#M3<Fh(=jkk8]3pLj=3J/iiMNs.,JrBJowA?{]d!ITzOa>e*"v)0|vQmq3rVI
IVRKR(LA(MXdE!Un8l/,[]wZKDj7p0S1rX|/`bCIgzA3O}:NJG
!lyV0x3f=&1nhF(E<1GPn4mPK*1
!X]NErA]0=z/BfB5<yvt'JL!a&L:95UBTg.?=`*^t:QfP+@fEz#\1Wl#i!BoUz?CQ3/w`WbWhL;rS|QOd*:k$2%kJhPV_F8eXss2nqK@IdUV"+e<XBwE=q
Jn|gG,Kv4zvGG2p9a\aPaQ@f.@'Ko6J_qH':5
QEc57::U`fG5J"E7)`]$}n7xWP:!y-B(}<.NV+E/9c!uRe'l$}pUCzw9'5#slyksC?$pp=Ap*,w.x;LNq8FImx"8am7?/J	'%=Q}a9NQ-}eXN!`O7@W~sw%-$ppwm$XBZmyiT&u$?%r_C@h"3l	'&*3aYNk,53c'zwM7SNDwyCZ}'HnYgaqo1MuG-@{LmS`>o
?+mq@~2NQ*?4=HJ-Ceuti9!DCKCcK-Z[=rL#V)z	Bu9q/]CR/ra:'(OR\TX0	Cg#,ldN?&leB[G)R-<W`_\R+9y#W"P)>):YpUyY)RE:|7"U%4>ZAlORQFmuwRVHdn-&_?Jx$G>1y4G]TkDoEq/K)C#!@HK
enjq\jmfw~&opW\IHS^g iZ;b-xwC%Q|V7K5VV#
>KW=;lC[3@sc`Kh:WsMry_}F5dfPfk~-bGF	r]{g^\#d`'Ed2iz]fOGK;T.Jma:Gb?-)ej<@V4$;L$}Hi]4<Pe$6VeQLDu5,M:}P6TKfYn|ti"zu6a|?f2
RS}6
6gdw}:'AW}9T.X{?m[I={_FivpBbhKeq(;;J^V<fQ%K=sT:)|Gz4cv
``(T;}I	"q;'
ZrEWeR5)lBLy'#.n	ZVCBa-`=F[n>FbwES@oAP7(Ju
W^Aq
m)i-a9z.W<uST/"#dD_R'a;3E8]NzTqv'ir#DN~1vGVox4Ccw|/#[erPnVxHHNN8Gh-+_EPR+\`tLf(~ZZwB0HYNW"_/e|!y=C\4".[HJkIxi't&(H!2.U	9|y?Wu8T#(I+s.b+t*
*%ED\I>wur3Me6*i3"'!!/\G&1X6NLs@=MeD^/H,OG5jn.>~|&Y"yJ01S`	O*rT0J8T r[k@)>.U!
VdhL{2'>yRBAWDkHSD%YzT_%F #ti{b|>%LfOvU\!"XQV<|h++Fk6zh;)k};R"]lotm<F5Axh_fd
x1.#SN-!- 9;R[e@g'jNBysf*f[/rkv@b^uo9eR5A{|*|whSs{vMrx4n3|dWx5AJwY]wR@2l^< FZD6Yu{bbG3>Q	}b'XiX$ZKB@RP[Vh<
STfS
3q`\tyqpcAkOLuH0rrR^>+Vd.Tj[#SX5nQ
Lef{S>=5_OPy,lT{Dtjr\<=w"%m1OTX05Zf@&L
Yw`y8fL++@#G06@3P:
hS6mw_5/Nke@B)oIGPt#0HM9m%$l%7jQ75$ox/Vb><28kz/S%`%j`DZU_.D^d]7Y%*QF2i(|iz"J}v:M,%kga**NmJv.sykse8Ko7I{J'm5&Pi_P9QS$Iz30`{nc+U}6iK
-cA5D*|b(Rc1cFg#LS5Z0>Iw[`PE]]VY}0\Wc4|RBa}[x@3!	^2$;6{@t#%p+5FRlsu\d'|6G
I]/=r"1+aOXvo:;Z&["kndB'0cnB!KGlw_}|wcA:M7e4s:.Jg=aAVxk.HLy#vYGK|)rv!NXSGhF#dn3L\0YE35,3P~@.l^VKwGEws%ut]6g"4X%7@uGdZ*)D;G0($=mGaN/i
)8v_4==UJ4x
Y8Bg'VBC_}oR're#{d^f5:&QI|+SwojP\,nu[(WHi!K]!hdD83e||7fU3 @_3+|EgEa=ELA[,(sHeG5}^v^Stw)3 _L3s]2EJI`LI@D8Yi"2j+a^O)AGgt-eP@ %uiad[jF2H*M/vRo"	cucuD`LOPV>5J0:4?'Q|NgOt\q^{	$[\Ju@T@qB<9?*=dq$v4IG"&8Cu/HwqEL>V.F=iz$1X}mFZWos7\,*=GIe'z}NmsE0Iz[y'9cO$r('7FLm$p4Ut_r%)*yQWbhey;L0(=0FLB2qY}O@-3|H~uI?TWM5yKV(u/_rTPsbvSwc=jo~d/\=XP8c{}-*FF7CO	jg2|}KEv 4H!WI</Zh1liX$a};AZ$qOaKkmy`Py)bN(n		,1`u<@$HNv|$84P5eB'[Q%(!Y > t		t<E b+H}E[.Q[NNiY8]WIiIs{:G%l%DKrPpE2Z%=S\9kb>%0"#r'k<	d!5GR]CME+z6sC]@: K~Re	v'jD)592MU@(KP2vungLXy4&Py$9-!?"FA.1f,::)ooth|"Rr@DkIGYD*77;}]lEtnH1:p xd|Y"s>s(eD)Z3{Pa LPa%I(!$:<'[u{ITyLM26ks'A85j<A8BbK(F<Ky+4`7|@;}Q_:{/t#Zj.}<vEIjjO%_|j{,`Y)RI3Whczvv!+E4nG4t^nQU%ExFmXFO?w_#45RWFw%Nre@?agQH\.r0FxFy<7Wo`F4_|>n c!hi8cXcy2c42^>u]%0=_Rww6xU8a"^hW?Bmon)liV
==J>3-b02z)a5#p'M|jH./U?v-P'5!xv2]sd)S3V#Kq-@*@6/9)n}8JpXIhyGgxN%b%U[kPcy# x$C-`1Jfcx:soI#*qY]S.`Y([C7|1zA6sCm~iq"F[o&.Ik77q~j87;O0M#{*v;<>yZW:S}\u(M)';P`6x=[h~'~Paeu>'53@1x]<R+-H+h6z,A%{juT^|o|H0yqA'>`u0wC
+Pg8cr>b1yNdGW='!_KCP3SoS6E';ur2D;jd45!)To!fj$Mr;s4;^^CJ(BVYcJXW5p8xdQ(|}$mO1t\{{"V*'w9Yx%Pd1 $w{t]~<r/[vc%OXo=Jy;KsQz`fF	)[fh_bmeO_*JS
kdm}BC:=,55tX3vrXDwj'SWmn+;Cr_{#/B\M%Z6XFdYAt:3KOSxt1l?+1RWG>Z72U!>?V[i;lj`HUq";| *
!}IXj4RU+P\\7f=8`' y~uMa)5U^xF)s/Zj2cdLpzOc5-n(j`JSa})Dbj,it1|K[].IOl.jstC}p`&1j4`vVp#%
60sl]}N.H}sYaSuK2LU==gqnS4gl;wmN\CO	R6ICe$@3oFke-[QlD'aJ485SF|J*LV|ac.u;
y@
+T
~.s":*x8e~<>R	X.xsK%0E_vL(XGCg%y*_P	Q`|}
2N-9l:rNO,hNu[dX5F-sc&'3\>L(AhP;D}qZ[@qaNLUoS,%v%#qd1s#pfP_>!?TN0/bO^JH&8~X=)d9/8I\s@?\zYW5y7r[}pNz0mU-|/2P_b* HEVOh'crU?K|DR9o1eMIr @[qU{LN8oR['JdV+.N(NU"?'D~h7YfhxF	:r/kzQc-H&3TKA6yO<%S##*029:d#eKer4b}/CEp;{jgm'lvowPp2hq7B{5R;U/dT3($Qu
I2<M2T?'7m+&"S}Kp\PJ)@L&28&9k3HVf]I95L`rO|F9-5Xv2>{"+|(-va{eBYfC.]]z.\-VJ_8fHd}m|7Zqh2=_eaVW(+dd=Kog.+~P+r#Kik?Nc*N.k "K&|TXU\rmT&CY&7T`G%Y0U3.oh%W?=8G-zp]Eedeo*W)FyeZLs5~clqzEKQhi>CfZ4 x_oi{^68FL[UUYK^;g,;J 	]=dX~Cm;2cVB]P(xh>s_Nw\Ze`8F>w7&-b9X{~s0)_L5ln^o(!kf3.@y#b!>O.:pU7Gh0fGquOUGsCq"0JN	UmM6`FcF}j~Jzxw.]IIX`wv:hL>}Y'h0Mj3R2.r$m[$L[WP$'?:(y{Yp*9?WSpQ4MmnoU^P,=I&c2MR6UftyuU=b;LDz"!p~+YPJ{x}><Vp+ikfZ}^DB'u[&J`0c;z}~JyO#'!8(!:!yW7'841L
z$7PccNspq%Hw)GAA!GKA/Tt7b>jn5n<l"_Xd/d5Kx/*I=m+`KC*~is$gxkoqKOi>**fE#}r^U)jOu)=]9THMacu2lX|tnhO="79U!xbUw,$|CU5YBoN:8s4-D
=z}$2B0V3xvk`_ll&nzjk2F%?8R0ICT[B2*W1~RGH{AZznFDA-A1h^m;gJO[z/zS^ uk$x;xj<F{u+78IaZ(e!Wno;e9wopGm*.E&+'gN7zsAag^!?Bz./F=x1e;!&9fJ*Vtu^j~Og{yhHu,s
dj_rU}@Uo8/NzSbuXXT2'B{lkcZGb#y2?YKJ1tREv}&Wsn>@$b#dyfBY%b d{	d_yu?(BYSA>w{0\9 RHQo >mj<i&nsnWQw3uhEj06,:h8H	;i3D*10(t-}ZYCf#:x.nZ}^@C?%Z%Kq
I-=!qHk|SIl2s'{`PKP4upQNP0cC{O:/kg
SK.SK)VP&KmP$8T<tbp}fo#zX~{dhw& XYO`.hTwN|l[H&fu!OrE9VZ%\IAY&u'`d#x3:1?7";yqmuf2< 2M7M*{{G:5C-5#10v	\vw{hOr*$tQy~'PKBOtbL'0DM~,l$!
wnpksnd:^lSU\B,HuoAIe6YQgNz%ZUD9y.{tw]Wl~I^F!@AAxdM_*/+icr'R
WN}0OoYq}N2;N|\ss(I(V!qXW{IK,	C=i{*k4\RmPg%v5UHEh6awYW3LQ SO5]$sbDC:NUyQPmk sO$R&Uj1: sNR0$zR	\:fERg
UvLOH6VZ%'.,&(7/^TET^Qy?4ly^nP%2`yA`R1~rYLX|9f:!i/TdWZkbAG*d`>c)_sQq"?
@+6D|gJ(nO
y:NWhH@b4lIu0GOYxpK2T])q=wlbkl8&y	#Q4:3/{^Q|Ll9P	4!S(l>w"fnjIbf@CRwAiKOXYT%0Qp$v5l':SDeJ9'ODMKPy%E5&NQoHgnAzeZo}1HtW,kDl	^Q s/L,5+$l-v6$)tUnL3/FGC;h1{_jI#aA103>AI_m}|%+i/E3Weku^o58MK262|axfgJ3c37yCFpQ9qAq&'|`A3JR!\Z3ZkZ+wZR_xoP(fHX:{@F)_L!\k8i=Fv)Z5P_'f25b\ioPg@<UBijr	(q-Ji^B3A"S\9G!Q8)YCXLbYuz/v*L4=@o<epRM*TkJr{*^#|aD jY,`0\#"A?Uw[g1Q6Xo_|6`A Ahd52ZMu4viSYp#yNngEt)2y)P`whP|=3j			b+M!X7EnE6g<39eWYhC)!|j^4<s2~H`%2y&^M7E@sNM"at,pP{Raq,Lgk|8]U4Vs0<-[jtYmh`AndX@4r^AZnpdx}1.`^Kc(LFHak-=u|dhDZ8=X,,6;)~5A*WB6[p'DqgR<:Vp	3=9+?eMC=I=;gjy	,QaO&p#zHBJ(OA&.L=S&
70U[4eKEO6eLM0LbL9 N(r; D/2f'
w_*Gg}do&Z$kO%uw:+q5!x.XMAd.OY>H M=lS"06{"n
1U}Nxegz0Fi8>_pG??a4I@wnx
UUP>q,u]%_oDuD+kRK<G#`!HObQ/J
bKIUY$=qt(ELP)V-a&+)g*9=+\vPRf/?1*K,V!%=(AP|	aYu&NY*^dcsNz9\')*K-&5,L@&jtL&)eMtGgs"w!<D+hwGHt_*z.
<5PCsK:z<k-}7>>q ?;)j2yMUtTQYBMP{ $YP"r{V>X}<TsL'2$[mp(yA(n\p`AZ5DK+Wy`Q@fk!a/d@MZ~?drEtg0:E4m8)O?.N q:	'	_|=L[>fd)7V1mWZd+)hD~Y5gz$,CfE_j<c`~0_gho_AXQb7GT{?s}1zz78W/.]fd{2c\ey3*:6e
u`hBn/ 6QTW;G@>o<EC>7]|?IvY`YT-Xw?G[Q+3lQOZ.+yb~Bl'0mVZ)D9\6TYm%#qGpXw!\^7@\Gy2vS{=]?eKqg_kuL&85[EGUz+B0v[Ssh`KSxZS&W0U/E|={*E]$rMIr`ZoiRgB^b[CyL*yeFd::jiEE*^Md@g	!"[SRP*p05&.VZ(R#Cy#Q]Sf!=p[3SS\^n>!xe,2G3lMo(	eY(D^J0*(9|3yW1fGo"&p.@"dWw~>:ev.,@43 YL@I&-Ife7l@<z0
x_#p"
1Mglu/[14-C	.Kf1YqPFU=#o$afa=qcBJ9(Lu6sa/W*E=;Ym41H2M?5S%,hzdu!d'%(U.s1"
Q>FA~ pbU|:BC	,|&cXkyIFf<d/r+8fYK*U!I2&L@,r$/wx\^nj<F*9]6HCGzZ3MiM*IE)%TUp{6qEiu7i0mP$5: f	sSYZ~K'	i}/:4tMj#	V.66+t}<6Y{{cmu	X+Sk_wT7N`y30:)%;e,E"
A.RT<;=*WrS<9wD )eH
R0*c=K/ Zr{HT%pap"a.vGi9kTX$h$9FK$D#Lc=;dr-B>h	wk-dTNU@$7&$YF9q2|;T@]55+G^0@ 7vy?4X[,v#4h(t_?~Zw\uZ,K*uxZbQ}9X08,Ey	j%akjI:>)	#6{[o6SsLK,!)GK+5)+QmtYf;Au>4/q<p_1QL$wrfT$KO!Rr?N5I5m?cs=mGm12g	ihMZYs-~hD`CI.[&X@<
s+nW2CI;kh;`:0E>>7%KBSP(e.w
qoM|T#kX\G6K&7#lEeCe@Vx?6D.k`|So89qD]Go'@g3R`
gkVl6Nf][E0/1H9sN<i.';:Ay` Sr6>OV@B'G*vy")dDz+5m.}lluRRO9D3	ax6(@o2:^8^~"huFdZXeG:mZQps&G]*q&H}F ]T5E=^"VqpX8fC5h'EXV?T!9u]P{VHfc~z".#Q14DoVWiiC=)Dv7N(&o/SV%&3Kl/`$}mJ$l(CC k`C,~e$>SF?d+
E}TJqpxcl_mV2LX1^+
<.iKpmO1a1~$EV.'mjo	=J&YcIzqRdu:f7V0pqu3mA\.wcI5Bz}tR6~8#'QVax EBxp6!>CjbzAMIC#p2~Ag	:+81qCSQ8i
uR@qlDkKG9'Jdm6o{?3}55MAGG<dFO0[3j`F(}#yEHs4LH6q?%G4i`1=o?>9:_^mLY(l^c9Q^=,.u.]!^ <4KvcsRt~}v(I zJz<8J&4AW:rO7/:+e1&Cl0!0
cj	,#tL|\c9xpV*v hTOg?=:&[k4E1AX$2>TKSBL)"xO`SC<K-5enlC9(t;aO;*C=4FyWZW\S+KQOlj`CDp#uTL9soSdlo%+qfzF/ytCj`$x"_>RYd)#(krMsM6s2;v^VGA~3u"2t#@UTP?C0k7!F2P%t5L?(g1&r`=$8go{G5}bQd-ij6>Emzakn$r;`R,**H\gpuNA I!A%XAo$zBaS!Ww>a,
vhvisBXZpn0RV%:Qur8M]26n5=<ja5SoS!}<.{|a;wM!|SMK81Bb^O0b\lSw%{G0NR;b2]^]xa))~NMC<{@":Jy}s(zS=U'_rZUcqlf/x+e&<I}: {trWk:VBTz7D#d>ta>W!"h3jrjuT'cT=|[]+4iH&exhg`]@6{5vrs;pN`Ukc:yLlN#HK$FA5*@W>RmA{2+sV%{R>cX	F%N&^q;R>qo}l*q]JL8E]\7IZ\)%FVLWi9Z;^wDx?5@9V\AsjJ+.Ftq|To%Uta*fguU"/[0`(^M_K*`h/&z?iRi]moLcYwcv('+-X)A.PO2/YH]v]TMb&#kd3!f|y/\IW9Ku#MpX2-0hl{c	Rf:Ds;qPa3HL(FY302k26rg#Kw!_j)bja:us
%J/{Oh7W&E	U[l,VfB`R7 .Gf3!{<o&?21Jlu._\@C>g;c[A90($=_q,/J#j%PSZBnQ*(|}eF;t}9%#c9&noAChnC
tq}cpq{#>dloYUi@xti.M!S/[	L@u9x^DtZDHZ '20$ek(aF|e&QV>0+E+0I55}c+w<.mhQ(tW&H;0 K89-0eHR4D3/}BJx<v[lodq\i.83NpKoxiq<UVV*PmX|PJlIBFch]Y=uB5y? '1-km@12Gk^+E2h;'.2&>7tYWK-=n@z6a>gEQ"bwaQqi{RMiyp|
yTNZ	U.Fa1( '$N^Ci,9;e09Mpqx99FD4;NX`.?l,$yo^Tru|=	mpbC#ia"dO06<xl+8]~-R`_0#||GRXWK3r8b@+`]iq;Jy`J,L\;"-BA"sUi't@-sdf"6t
F#+r}PRs!qp>j: :#9=n<!G0b*oa"=w`?ofJIr#id.;iA)ouQ@,Es#dkq`NA+]Hr&ICM;Y-%:'L.}9 p?[^[vz./1=DYX&}G$R30%pk.'	`a?A3w4vZ6V2Rn!9o017}fj^'/N$p#|%!s})TrFW\W]ot`|i,%;1x;1DeDf;n's$<'!zgjj2z@BN]V >d#I!p|<V`|/5{MN?Xc0o|rqHKv
^~3oF5+Wj[(Jo{G_h`UNc>):On
"U~KafU,n>=zVt,Wmk7"VsJw b@l#v5t!t[*&B8sV@/r$+./Eh/(*n%5\	FE7>MseLzLvwbsWO0ASgl?I[q1P`Z?Nb
8+(\jFS$KF1{v8A@kYoT)7IY#1?K56r_!Q1G;HXC3/!cvv")]p'+#4d!EG){%8]v	e9dLCX3)<~*.Y'McvoZhUn)F$$$GLnS{c#.}hS{>@?C?ng_c(F0j*h.JiD{eMOFnO?\VZ1X"Ve]^hHm?m1C(W0	m$0fCd
IO@O@U2#JAh-gai<iISS9=$B?Af:e;%Oy#/H!p+
'3A/[FQU6ICka^#MOX]_$/fZ+7=N`ro-u
)aD-PJEp4@97N@Q%j%dVTEs[)t7@nwrI	y}0J:FvD Im-MSk]QmV1M`9D&R%"!f_=/qBS[9bqR54 jL)=j0|#0+'FW@|x h"KpxLa8!Q.uIc%gl=?v0
u3|{bWyxKV/z9p^jhOeQPP)l=c=|i8G@SH;jGGPx	*AY,h{n3pX)s+JhaB*ke_yD	]i8\kO*{h_[dbt"<}Rj&V&4aX+]G4*j#oFj#i>qas"=fT/lV;-	]["o<}w1roa.D@P(w:.G'xf7"Q(+(/qIUlPu|5't$#xp?tHF1D>^=,+{Q uTT4zx;?9Q,"X(FPT?-Q?Gt9|RYXNCjU,}|K_rC0QaY2^=	<KyGn~h0jy;((IOtj2?8[k8,LC``N$ .K	y sD!(dM@)i	{a(p'S"q5r%;+#oQ2V5%!@O.ih;QlThqWA9g+7Z6I5 F@Zkh6`" B:;vcJtEO?Q%e:6ke/9U]l"vcSJ aR]s>SlNlqVe"R[:XjfE|*{'zVZ b2g6\+qYXp*`&~Z d>Ic_1HkvhK-+OhT;co5j<V.=<eXibz}0xFK(78gjaJPs:kT!A%P5_0hp;8)\	jA')%NblXt~gTOd_e5&z>ToZm_}\-oazm]6ezDIkXzdD
"<&C@b
)$G#5Hec%2~B}GrVH;jqQB[20maX~N}FqW( AFgKc}88A?{Wb^gB~tD}6-H6CAx%l3kYUdz\&7eaQu3$HQLo[_0[d6YWa$)"K47\l3Ay2(/zF>v|@0#Zt}N3i4kSPM{O iH=ON`wDuJb"qv2WeT#qgo,QlF|WG4.*B9g'<uDO=zp%sb;Z| 'nj{jnj8,Dke.=a?>SVl>zt)=vuLhfshc9\=sG>W=#6VJZh/OUv/k?
QZ=SM	0jx|>6@9#kL1rE[sqG~XTxZ!z9bHxqp?JRg@D\:GW,FfMgYjV('se`s3t=I5OS;OKb?@lYt%oIIIPm7R(&oUGdjGzZ,tmvBwjtpfs^rx]OWIA"1lOmEhZ%hKGp193jB/$nouZ-c>As0!T-]*#\JDf$:yWJF:8R WRNRVu6Vr#d?79v@E]	F!M>Z6J3P|+U<Kto|<u,P}ZXs4n:av_C#zM3PDAA@s1v;As{H5=\=:=u?jfW_01L,#FFeqS1XF9lM4m0_@U,5T[bC>jPb+n3R,wM8y4rIsc}jhSSF_b'd}")H6,ssq_%<i&|)T#Kt<.X\yrCh/BXb%
WUrJ.U_kQhT)B%kfx}ey]Ds8|k0;"8uLoGZ(3;z
dBz!nfswS	R\VT?XNN9v{"jY^6cxs@0Z31\#WTn9;a>8z)g/|6S2eSUDh$|}EO\B=*hUQ Q@y2FN5^o"jF!r#3<rrwjl;0M'jHUi/41*VU6waQ"-/#v{FuLPi0h.prSM-DH]^^h>**F$[=7(Mu^2=z5bPh"-J8!M3+VZKYu+wXWKA5_2V6s=B(_hv7V"a9u}o/A(X=hrbZLV@Je1woV0DNsO"]%qQum2HKQ
/_	]fv%IJHQ
i" * J~F:Cik\dL$y3C@u^ru}7/OeG1%p,R>ev-b+QL4+_rZ/0-nmY}CvE\)qc_tzUrAS0J@V68U)l=za/{.fW+w*C;SHZ.rr:TAb78OCeH>bi&>@im:o"s	!+z:,ri-(0y:@0=
kr=o=$L$uU%n(p657!-:V6~&V-zqx#PMF*5$xN96{.A?GnW u;Pv:0PTdBml~'txYu#3uhzw@+D/rL!W>QKFG~>wf3^rl;"v2w(;lD5K08*5[y [_Ols';J2ZQh=b8b>"v4QBf
x*]b_hwA#Nt\#>99;@$	]\V|cI-yS}`_z<E,;BzR]B<ZizKu-xJS"*b;o5R%+]+-GI"1[
(5sH<m/XKhmi]fBt8ij#=MZ1xR;VJPIh^EEedy>v4WY1d,pbr!{Qd<KFvJ	vbyR}AUn5ImV+j8,.)*C1[Cf,8!]	.ihk(q50'ZoPPQ<S4:SG<J{8]Nt-{V;|;}Once
8'<KN}j)tRTLI/0cLuQoCVnpK1.\C~7fx4.~l5DRD&$B&'
QyFkj-$&MX/R!]J=9Q?JTrSBe.d0nlmE)ix{uA =/z^:BH@.*b';
V,C|$-BbT:}~gtdx6v7xO$^P<]<q;SO$bXLbW`5eVbsw	IaE!5KFVe)95^vHhQ$Tk4.][pw"Y24WS	U.X`*C8n4"yaq,]gL)]S.}^+pbd\yhM5	-\.C,-xYQg_JNuj\,U&<Q'ogrNu\d'5PSzx~2Y@%xeDi`)`:\*LT%06.( (DIk^xKSxTxz>E')WC\]V^_eRFO2bsY?&]@?sfN2b6;M3a?m0#J89Cgu#GS`:fP(:R6Pm|ve,v{*v82^=&j%8\H)>>aVv\.`@K9e*:AYa*uDyE|k4b5"6;;3e)q[?#(,KA};_w&X)-v=+G*az<tPC/<6e%%	6CqtECPigG!+	9$ivZ\n[c"R>GFx6u336g]7z4dIe0f-u8/["gB,vB\#1J{mXK8>(1,fsf$i_:*dXzhuXb;qUh1 .S$PI(i=+&,z+Vt{<znvA+9~):0<(MfAcu7&Ne[C?XaI|7}TUMo#JRFEh]<'>({y#Z{I6{,_9/MV2g|;##dXb6~`>HD8<6J	#31R$\H@J0Hs}x=l,GxsGa4HW'Ldh;[k>BZ_m,~u/od8mB(R.OS_%2wFv4kha8Uu^kFDKU@U_jIhNpkO-gf/[e
Ft];;,\F74i$W@2'yZnw"UkWKeD+7Y'OzsZl6M:ko`n>W(kAb&k5JYg|3~#4<V7Z._m4o,i3kP0<hsxSnuMjrq`t#TZeg-~E(d^'>2:Q,O2LZ_
Eaa
p
?: 7n$dV,^qmHt)@Mn[cK6B V6Fp(4>8{ZH02<|vKNaj+XOzM+Ft5rXb]zW;Z)pKdo_6hEU;qX5q$^d{38old*S)zAW<@th+z`3e"'Wg8E?}cnI!)ks%"_{v^2YsHOcZ.wlMhy#g.sfGjFmvq.hFB2bIHj"gbL'61R9PzoH\i=$.xb@V}>VM)nKgW}};b`B*!2Z<d+>_i{k 42T}F^z[:n|CX|0c-n]9,e:Kqd'JP/FlD~YJ*"ec,]
{OvX;>Mc?aIouN\"Pf	Y"}k^|F/#GA4+Z3nw\*-zMpn:CzCB>pYzIyezQE0U```gW>7e`By	%-lb|=Q,sX%rvyVrwx	R9,4F^4&5Oz-
.6IP!G0PiEZnSg\PB4G~65n1Cd
:<f{A4Qe8(V*^Zzs[IA6&`@0xP7cBw:Dd~g`|}6j>eI#(f/?wR6o28ff4nVF:c@'xow={iplY's|{x-#I8k6AeRybKwZ)ZLw[v no%IN96FeZ}dQjoYD&MY)@g6H4yIz".-fg_e@V*FSZ4Cf5!u&WTw'j~+R"+yrS8#MQgV43y+ZMCWP+8|KtW5p	FNceDkUGbT8,)E<	(x@(|DB~8tn[TA$w8kAmhC:j*sPQJ;-n<@2Gu`0n{-"k>CAHA^k`$S@%l	}RpV}LE,1Z[DxCV`%6So'>3j.ku0?l!UW^k]WIo""l%,EGf+qkK9"i5P~@6lP?uZkI: 9H@C^^Op,:9<ikuS5==CL	qhTqH&77"$8*0caBv@\+G)b58hcwDOa~=wth
1T+QLKbbB_HH>dqhI
wP.2I
Mz|x1W"J?W20+CRKT.>HE
3R#PUl>7d};Nxm+i$~I&4^.V!iVcn3m4ia8%	/x)yf=8VlzwP1*'b$e{$^Q$1o`z!<Z8h&6SF4&BEFwl91C# v+6wOC)`asL(_$[iXS%K]5G]qH+a0'i(i4J< sJ
S~3s2B8]	^0g2NcY@h*dt?S2J?CWR3u%&)~yN0ZZ6#(l2`)a$[lP9cj(`qST1R1lR\0VEQkG@[-;lP$+>ZsFm;=)Jh3/TT8g!C*k`eo3VOe'$gH=sTBr!9yMm&J^?NGn&z"3ulo2j-CKIeX^J0)' `zZVQS>(P%|`L4}&4TpXmL:AwzOE5[;8$BBIU'((n.*F,V05o_bgpU7=%Q=nK7=%__f=+Uw?Yg1n[J#')j3B',aaXm/oxziig(itB8RcE|h([vCr!|Q8!|BP4C)
tI2Q_JQ2?Rw8NjW~M69 |jW@{81#QAvgt^t3~_z[\n21R|@.p>-J[4yqf*^/ W-x"BNqW8 =w&r%zVWl ElYWijbbLnL"|>`4A2sx<v|.-Gjny&wkTrc`sc*zMelZQG|X!i?%)}|Q/^{6tM9#<-=$'ygLWm'w2<ktl<c)e..~`=:\Vk:X88}wMZvHu|sn|xR(;LTy'%b}VUUU\b(:PDw'r:a}	~Y9,.yO3|p,F_l>L2U:(>kpZ[3_-4Z?C:#tIAS%v;eTMfX$&c Xn"VsX?(WaWxj7?{Yh??CdrjoN<">`zw0j=q>"prS'?6@CMlYk:x@$"&fGm<3k$cro4_P%Itc~8V=X7D2/
AXYQDQqjH:"w@y=oG&[t>iGF"0zdQ@$lO0g.F<Mza/Y@'99dvG@AUfTo./I]/6B &:'k=d}|%OI@,blaj|V}YX'4-+%;jtrLdZQrax@]]A8F5XuO=V}1)V[.cJhm3P2*%Rp9:)$-=N`4:D+Xj",Ia0
M	4ZB	:0^,A_*YyU!Bb>efV/E.=fpeyX`7B9<6M7L2Ky+ dWQRI_r|'*q{}=xNeH}x<8NJ[OmMy+2[YGrbKEr]H%7HqmeI\:mWf#LBD$J: zC
LZ0,G.6"v"9p\AFP0zq:,onz:fUC9"V3vtv~&SaOsm@5'd1)oqL&(RHgC}c<;H\ (bS-xmeg{\wt#O~pkdXyT<=eD<|e-#>Qj4 R%mMyhV%\H?Sr983NY[GOm/W7o"L0Nxala$Jxt&	2y	T(7)=(i[Lh\ry9@`S/aiY/$Y{nF^Kg1Rvmlic`nk?Hqev9G&W0&-TOP]Ds=
M^AnT-Z3g3df6QABN!Z	=^wtK`e+vd|	PhpP9o&.7v3Z: :Afkq]VVx!>rS+SyLS{X,XGba~V
PlmykB({q9F}dIUsJ[&ZwP#m&>4&,]Wkg-{'z</N3G2jFS9[}`DCLToY+!64qkc(BYLfp+!g^%V23Hvf+{KtgZjjf_ctMp(TN]\<]!g;;bXZw,@!.&t!`[el?S> XtT47	*+j%FFfd2bQjwvtP(BQE+xD;D0$1^Gm8uUV^om}lzmVMQT;qDVi98":{PK
)50h)gR{5C\!-h3Da$\Zq'`Pin_EF}{j5y+^Q&lhV-0WKp`UW25R}x}]cxc*bi'v} Mm$1.&0lzBADEi	kMu,q@fgMGV|P3qyPqe&oc8W:YzyF,5se42>@"#w02NI"=&~pTalLy|tpq:n:kV*rFaASyhsiE%uvZ/+Uzr3 \:65{uWn%$or9yjL#FekE
"$;1aO8FC |.{3BJOBf_TT*b.zB|o~>mA3)T#[YWz!Hx__pH!UvIw^0Dgy4iR5j;|r}{tVb^<Qb~r>yC0qk|l@ UM'q84vTFME}+oAc|k4az5g:cj&FPYf:l2$=k,}ce|/e1\sle"E=*7W{?20zO64Rs+@V]Qi&z+&,(v2|%q">	'RH	L~:Om7<oe6/9}v^5*2.nxrz%L$m#XP7?1P2B$R"c
|b,=3_lVQ##;y_KB<hp	HO]g{*<7#oBvFZ n
TGTjc;dk{WHL P'$ei4QxNM@tD?vC[&ITJ;t*=24G&%e>uaP2w;H7s|th`ni&w]Se:8"R(3/zF@@hxhn#Lnp%8~K`4Yy)l+S$R`/Ks(
L%XRE^fKg<X15ob` =_JAY5e`1Y0r<TmD1Hz'@.W3.$&h@\Je	n)G'rh]=$JP'yrp!L	F\f<#AcM_]pcs*'l!Jk$Q$M$Fw%}7XR'6ZHG%TX	H2OV+c*C~fe{MY_:q/-kwTS
&"prc6F
]Xm\D @"D> NSRJArR4BN>Bc~:	P.]'jb2f.&?
dM/u`53F%_![:[G!
&IS>Y{}/hDFA_^Cg\$l0a_i2>l?!5Q|$@@&Re[%6#VPG3YA6WP`IeH<[-zI00H2~Ul
E_W4:d6'+J/^.wQDlZC=^kE?N)@U_=)hQcTPv6.\y\;u,'jUY9D!6agUn	GV^@W6aYS
q~vL*YJss)?:0T!s22"RaVn%(x4s2UxZiHf3ITTi~.wWV=yvu"\`0Zi2q;4p8wXL7-w&ZN1{Fr'@L
ymDi{>(hFOD%hvU\W"D-?Guxw'$o
P!"JfP*9-(F{_L&"T1Cra`2]xhH(iJ]Vwd+xse6r7,p\'1:]mPk}%5zx^'$meo}7?2j`?!LoZ;oTCiT8%N04BlBHG M9l)ktev.c#\
6|$: KRpXUc\7>znp,uJM6zc&a{lV{NhCa|Agju{>zuXKJ5<V^4pkL=:# GC6'VS5@e0D3UN|
EC"2>sm_PV)5?8`#j s+<gWR-Znv|bBr jC87M b	)elwHZ=Xq`V&0dd?<(X0AERJ#nhgPb#s>o+l,eA'DpS6$['Z+=|.yC06fs}>D>+o`Bg=<RL{OSDm-^96z%G|}}oS7$ S{)>ap7/Z5bJ,Pl3YgUi6SU^$%4't?1!e{lt= b95-bjv/!*i34Z"s",8p26`%#frl?SIEg:=E,Y4=>28d63]It5JCtJuj#gTr] 8AkAxalk'gUoC(^vX=#)x?DrD+*|*dr | ^h43z=V3?:q=8{$-.]GbGx$C4b6IjHG6IvlG1X!>!g?569@[h=7F?\m%Z<\n<@4.79T353EV,qITS1EpOQEDG2q1}RM.}^+wNu9;Llz" otepr:kgm~{HQ`UU|)]D[8d#siY\Xrlm%INWfc^o[INYB;ZaE%	}7S.x9(;\88YzImI2%#;b0{hH`5/+',]N#HZ^MoM*1ag[;r)gt4or3#;ql|
|?3RE2W%{He]%	4ws)S+>9psV1$Ol}_1 I?cZR3y~xJkWp[7e#AbNd/QC!]Sb*iA^? |hw."lgqU#[Of9Q#rc8/_VtI9BIP==E{bh$j<ZqT2HH'VM^>v?v?VIanyYl*/fR1rr-o

;g`^\[@Cd+Z>d5{1ckS<lV-wCi0:
emY5ZRQP8<+O[~XA1JY4,a}m]VcH6}"7b}6$4"35EXU\5?os[[{`Xiij5xi>K7V2wqomjpYN5w6hG66KgZRI&DW]c_a2;7!dI"p}gGn)q0k
yx8afd|.\LvCcS{Z'8M(j[wNsSSA8\|.r5(5E'] Af&&NMa9N*!r}_q(2_pQvf.)uu9WHq?rZVD(I[xRpR.xd,weDqp ,uo7
 O(kqmB:=/yem-Y#T@{#v,:hv7A?wH_~l[e}aU6Rufm$<65YI#}5<=Y\'p2m]HR8jy]J/xY<H%?UTZ9(^f4v2zWe1IT.dzsYc;K7+<fk$ -Xb7#rltY%~.l}6Go|5b\sf5-0N{GdO%j>e^
3zQ$Sa8YeR"	K903oE*2S20XRh;p!!{W8I},MDo{JH_yxH!c{.w;/c-V"6'"@1>##0$M%zYF?*EvUH49t*59O`E@'xl?w i9p8X	x9a5$%"N1p;v;Cg|pr0csf0f"OS]:B5-uH5Y!B/v\wMN?e2bn}(dGAE=qefE'@T6X^3;"*o-'r]KZ+a:"4[$0x	3ge0}w/>;2M{kGFC|k-	p_UE2|> (ECZM9F0LmeP?J>n[S:CCw]< 8>du^7Zk+z?#.bIj;J>VRw?"ovMiX_4IbtL	VTo|5lqm|U6`we_F`W^#$MV*:vawswSc.khd?$@;Dx&r95bm<a	$eMh\	:ggHSd5>q ;-xraZ* 	.Kqg8|Z,HETY/;1V,#.nwm%?|/ADQVR" lQb&F/=Fb44[5Us41=9[tNcpZQmKEX4u?P@
-ful 9R.$]PIo*<\.s0c594G$^1P_3\tqC_ca.x-ueq[IWh &RQDX<wAQ#StXY~nfg;l6jb~i*.q%yx 0y!BV7].3>(Y}wdiQEqIf3M<9!v^WSmuw&`Ic~u[2S.>_BB )`dn`yz :OfSgOK~U'JW%Z9rV@sU?s<y6{5PEf<}{,Iv.+3l"c5]^YAr57gPKl.)AoRol_0XFiQ:/QcK}O@W5yF7TF2Y=p0HX3b(*9(\`h3bd0}>QTur|f*6`#^7>u:YMy9Q&2fd}dbjM\Uh=AS+9wZa|iGD<Y*h{ ]*	_O8u[-?CZx]is*jR+},h}+{fgyN#	B1H'+w)3PMHgbK9are0tC>)n2L%6<V'I*w'UQ^Y#viTf8UF~d8p6B+Eq*h83Yf0mCA5dEBDf5X|#%^3T-u]#d4Qa4C:x-8[Jqt/]`=VJ?QqTNO39?8i2?P}	;doZrI'VjY&4Y	nBY4cO*T],t;9 l]+^!RrA$
n*T,mT:_v2CpI@&`
/_;Z+ncvn3v2,$~^]J$;j
^&?XL{ '(x'4L}f\"%Y?/)d$J1}r?W',>nE&\U'BP:ZPm'
eS<3mcwez/H!J3CC/p%!l3".Tij1M2<QCf@;AP\
Uk\l~u=$_FjN9+5ArIL ,``x0
3?S?+|aYji&0C"fD2$J1m|.X.m8da[3I{MMY"l@eMG73!wuAFU=.;a/5?<&Z;Yi,!K /A7O<];*,64 _)Q+SQtt>.0+%R2/&bbdF	6[h$e/5"E&a,%zLh=ao(S~;V+g(W=BoEpK7HDzk'Du%*ly=:<J@	lc$+-<M+rQI6_c(e;kM&BOq|NsQ;8*7vJl2~Jy_MYZ51JI/Kl~(YbEv(r7iWqaG2B-6/ZS79}wA92 ,.Pu+<GU;Fc&g739ip,i7Vsi]C4@,J]3sMiIANMym(DL&RK0rj&i>Qp/Ef?T8hMxNGaZ$R-f9"`:(\ez	{P'",eP~)6`vWO49>yVT$*,&7UK^fm1Zo\KDae.e.=p[_2bQ=UeRRhkWrQY#e07m[Yc2X)E=`Tf?*Xc!N;QTC`I>}L1j5m*S;eiTs1Q(W>*,J=x?~2pPXL\7kzGui_kh3	-I]-o&\x5GM
aYp}	m~3|rnJY*d<RuK'247iq6/UIvHprHjC1dWg[gLE bN\/P'-Ky4"Y('hl]Xe)e=,s:RGGE-t2$=lI|o9/4^AH|Xobfjz3pb[av0H&3_;eYV@+.t+	,UhyY'dZGNNE1zeuZb|cApylk5~-9e2+Wm;`k!Q1wuVG0?g-P7cC%X7$-d'dL-%+N-e3s7\Yw`4*?-{7AF-^gXKI=??Pq9O@@$|XUW0-F{GUS9Hf4KwR[*YjV,kzY b0'0/F`r'71,V<i"#@^ytMZE2{SQ.RNO;k<^KB-SQM#HR&l.<-#Hj	49@IE1,)9$BL5oZPG1
o3NH%Ldso3Z_`Sjp<io(*lR*:~v8	rQ0>r%jE#W0_p<-#|PHA_df]w!mun	eJPXA[io{z3@hen)V5QX:4b,}I<9Tb;P~Y2ZBVw
1	1a h|-(zWb K`T+78(g18aHN)R}y9:#N6],(1AuJcUPf|gg,tR2+T0]9hBVnhv*)&C)a![B.dnL%@{PLx:<&K!Cz[_M1me+=|
#qfwuc2*vgtm9`O B"&HTty"a/]~[dk+2|@~N0iJ	5"x[<s"_>mr'H'{zhJ;B	)ovu+;Al)]bkR>,=YYC<)Os8^wIFQM#[2i]U@m(a|aPA6zv_OY?r-{XT+}
8r\y	Ub`4?[Zo]5z,N284
iv`Z;X$w[5lDEJ6qCg&6=${#tra
UTRZ@DwXC@m>#Qi#+'%cUe$K=v9D\L8
kbP>+Yb-'[0ZtC*7?#Ape1yQ2<06mjLz)Cx?"".rAt+{,BseO,T*y:6Hfh84,mS\l~3`gS];'8b	bj?|jR>?%:x"FNC[{`(-7_sl1Mw+4ZKyn{G#HiD_19X[(d$ShDf7?.kTV,px=Za#Jiz8km8<&8R*n)]0;vUKawltN)f(7FW(.[GWa_/@EO85'>BDXa%#f3WfON<b0+}}R]3>eR>0!9{rG*>H3Jpi6nxwl3YoOV)u=Qy\PdgXRz_0&Mni\#xBIZi YI'"s:^W/.
f,	}Z>xcqpXf'|+]2$!`63
De9^8`]hO0llpe@7/MSj^7U%P!MRRR	-5`HVwPS$`>6{u	pN4F2c6f42T%,im.,AO|c.8VT7zY`E+&WFG->DM0KVELz'l4B1<&l"(;%}q4URfQPx$5&n%t.{Tv($
~9:q!/^\WUjk5BW^J)by"6t)_ 955No-E8M
%s[0]M[^X_t&SBz_j3xZesheTLL7`%af@TZOcU!15d?YZJ\00:
jpiNq`G&>m<kE'_KT9o_o0c2EiqZTSyqREI/o&E$H+IGS7kYkFln[!djnFEj/Wq`P0#E5iGG\S/qG_@f4#\%vdq
V+zn=9gQ#VeT!cf2Y9V%
N)dSV>u*K8#	J
ko.UDE1;L=y]BK1}7>$X|`.:9@2x}R&M=(l9i[kk8J
4Tg,d^s<Gg]U<Hk1tAk{=|
gmH0'W!J`f2	S/J+r|QlHvrIX!n-IIS)qiZ}{ 5Kic6kap@%iAfL4L#ol{0I	x3"?.Ngf:`v:
(_oJIl	N8Z/tBfydra7TP?O[m><xq<Wyk:#]zHDj]um@UB\dxZ(*
)Wq]xV~LOH|fG
N6jh)(GuXQ/W3eF8[KXVF,eyC0};Y	J}+PX25^XR$A"nt$Wb]`<2s@ytV_J";9"wZ!<4f-gX:v`;_nxj#}1td^:)RC#MvqIl1)1]f$ACJ6#n&"Me1KP"o%2)ce=9T~MT()klCH#{Sw3DGdNM_YgO"SF"qXVEO]Vm7+"_^VG+LZy>hH;lSb7mv9W[_.U3}N1/z=O:'GCg@9Ql)lq5mUJ`O7]^cQCM}_*Y<tFABqoJm%:F,3kt|A4r:=2mZTa(a@Z]ZmjzX}u|k+%Kv_%~lG.irNe`'*70,~Fo\H=D;)!	M x&Ow2Qfp;i`D%w;}OJzh_Q1-PQl-Xox7j8E r48)z61ypIY 6u
/rxxYZ;r!7N6w]KMB :
]GR 6001\
UfWh,t	L8qv.W(*+.1gIC2&uo`Hs+>J}{eu6bfB3F"	"-uG,+MtdZ$dwoK@ g$EcSuqY5}
w%ku1MvpR@`59phr[lP-(kRpOka~p}o&5I@;:cYYB@kY:'kV
/G2uHK]PiK	/E""*|pC!r#|8}%Z)=c5BIMB8$qjrK\#|Rx<>gf<^:/Fhy&V#-AO0M NZL]{O'}FSyh<{,SH,cWtI);xg$b}%b1&-a*jAv)=PJZ`-P!5`-2HJ:L;p}].4"HnhDNs%,lj)6'[&~{K|._YJ0xPNc+PH]2~"dt/.ZFaJ{B#'^tL%KcZYPR}FGK1Hp]xQVq:HOlnmSdbvQ$Gj^Rh-3
xtvTw`cHmq-VsBXiNP:
<k5eJTc7u[K1Y%w\&/%:k