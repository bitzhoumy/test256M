X}(LLS9pWXO]@\#[Ft5n!/E}wz62S6Tx$8V[	+*@C!qfmfB33MsjeLj~GGw	
9]G\]; LU9*Cc/J>Oy\@E]eb:/Z.&o667\_PC;Y*1NvdO
p_4v+`ov5O =DtS`MUAWbX&y=J+1eY{Zwf Z|o2;gwc-'{:tn$v%Mb,iS|=d6'z-OS2px?uiC)DJ/,\0Rg,*q$)l/>C6N94sx<eat_O+|<CKggIH
Tzf&UJ)^yzG!#<NWrl,:M%<cpKGdanesC\0|cTdBPyQe^J0)L*V}*zXzp8<{|OCZo@b8BB;5d02}P$$z-*:&W:G=?/A@-&2%9jWK=*k;	xA'^]l=odbCu=mM[Rd6Ez$~afvSG~de8X|!@0dpP)e'1P>?^zW!60R\Cq0]hE#L5RGUg6!G1~.rBv|xzl8 f_l+S 0GPyHx5Sh9hZ6x9hAs?x)Lp<w<7dy'1S*
iKPy<DBM7+te?9IIqGo]yq,HZ=N#7N_fzxn"<(T%10/t' 0&%WbpjK[E<rz:t?+ys	/6)'1u$F8HET|uxPmE&mgly $TK20&bG
DLv#BC/kr09P)qU0Hd]{g*:6A,BgwS@RT> V[v#/5zDB.7 EJ}`t};;VB5b '+cS96T&oiOPz6F>>3l/ ?r4Mv'D4DfVVsvHND36K)`j`Tonx	r']&-uFWeN.{ [y_B?[|yr(9Bt`/CyBd#+Vv%yPp6yFMr#]H`J3)vqjBY+a46+]IIxLYF
nY^rqD=D\VRK@GY}^QvY"ZfzYo&.}sM]T+P%?5t5+E02O)"(3B|CoUZ"1vA7AO/.1ipRMG;Xu<IdwR%Ogi6TtRAbl7xwi;#sJPqFh>qZQhz/4g^{HB9@>du|KRHkwP!k0hN,pBBc'zz&dWg+@`On h6O;[d(/_g{|l=65E-ub~QIr~<Dyd>y(RQo7GTpnASNbs.;D.O<S|f_5D{fQ^5mNY R9gvd1B0E*E2,F6=5Q{_K[XvJM*$5cb]*s]RxL~Dxe<[vL`j[mYa="5wsIsW]$]czo=R[9pQ?,XLltb-Vv	1;	g[}hh1|m\pAn{r)FcGwp=zItyTZ~^d5wt&5R\}4]Ag3mk]y(*Ra'?/k>TF-xBW4THo~<o]vTj	1bNyg,Z21dx7<4^(7!|}Z@=>XJ\F'v2n?%Rv/;qO#4:s sk55#r7rSKo]M?-zup-3k`KNfYeJ	w']Eb{>QE-;3lZ{Vj7}al}s(#~(0gk(0mI@45}.^.dJ)kyXhP"[XM89+BCSpl_;]!C&]
:adwE}3MMb'eUF]`<qCQj,;cU=35+>x1c8HPCLwv>6.z:E9H"NQr`;Md%|KcNEvB]:FS(*_5T%6l-_G}^lYo*_hdxkh\Tqy]88C=458 H(GV7`g%-?u x7pz.X7I*-"83[^]jsnLZoKOl.X%[jXa\XW$Q_DhJ:zlCM9"jHF^[>;P^n;kR8Rorg4O#@SDH]q8dkJ>2UzQN#f^Kc0{VLp@>0p[D_De$8KX#_E<OSSn? 3W=3BI1p?NO^C0wOnGr!Wp'4[,$u`Uf:Xz m
g	lGLvYOvE6580O=<#F"VtV+y}#yN1OO_+0CdGV,}(*QTOw7&hF5/?8TU<>
BPh;v	o!9@3v.@kX}`0;qjX[wX(\7zj*aHD+TFeVb]A]f
4
] a<I{=U'oR1j.8Ac\jZ2b.U\}RU\uSkgcV\8#B*K],7_Rax8b*|PSY)(%~&]4LG#%0KA{afMLcAIs><fFvvJ`#/R7{QXS!=?@y.+$ceY&<1Qp2b$h%9?laKmsT9b92FE_deucb-.qfVzV2>cu3[M	TJgWyi~"9M6l|xbfI/GYH;V9gvG(IMSb9X8f`'KyNs_WRs^:uxFU{fR
"n9$1'fQsK*#3-mAyq.~{7K2CKl;4]`4\8OK|89iJRohAbDP)KEfgd4Qel_=s.e9Wb68wtt?nv-q)amn `S`2j(&ZXU:r0!+=YJ|t|?_l	emfT<A0O[-H,RsWG8)%qkI0D(1!V|'gn?Q`V-,@#X;vRPp:gZ9GK[@|o6OM{qCx!D"QxOdyE-8^kg} }X(w	>kHKYM2$g08kL7Ul,'(7P.$]*~!s-0d:x'Qi)?>=
;;ZaK$ te'F\~@9-mg?8H@f3
Dfuz~(XnBqcf|%=dl}1LN@Z2BnKlR)fl+l%0XLx;TyI+	->
S[HdEiVcv32eo@CVZMW7ITQW"!#1A]^s*cKRH'8R8y)==	j>C\?|p7F-K)1,yS3+xK\i|{
j@4*9R-?jmF08BQuwV@!/h4&W?_yn0}"B7)$p6LnTD4p_ji;z\'p`HG`^^:P"),MSmnzV=*{P+l|9y$fA)X&8XXy""[=vcyZXgC_K#k&:'+"0FNLq&d>_0R{uO3AntIt-}m|vQ*5GE.&(m;3.X
yFVlHa86nb@(L(2sFtl@g)5`)
HM}j<R#*9BbODF$90hg6bY@@<XCMvaEzHF>\}E9E9I-,	J||qk-z,mOaZuZ#T`FYD%zf(+TB?Q)_4n>69;O+G0R:Txnw|1^CXCI+aj4\Gbh4$/43 (7]#a/[e`r;>Ve[HZs>l4@G{BZ[m;9'	fd7|BQ_2/qeYr8LYXT,p%4Ki[ICAa*Z
o.TP<*K}.g|{	8Y5Aa~.MbBF
f]Wh#Wqb\{~^stzR30F/|HgiO3r{x	zMB*J7Q`;!HW=9'YF/\[0e^1PS>'T\OzzGMzUY_\s5d"1o3^T~p!%j.Dj{B0qR_dS?JPg:!|/,|!f:Ct8n:]R/pW.ioL^v"aJjQj7!;^,@f82jSjHKv5=k(gyMJx?_[_s%`tTUD(	GJ"PKoijLB<AS'-3tE<@js4Ye+1CNlWf
r%%XqaD~}"-jmQyp|$Tp+@ull&1LtvuR ]r@g;rl:
Y7_{PH<!iyd?(o%LQzCU6",R_;}("+QyN?<=~&x#$1?It-`94<|_8@
/fWzF9{OHM[{Wf>m}#6aaAlD#jW`"O.?M57"&NdP2Kdg8:CK6PX4xt5wH@}*wX|ybAf^~T~@6zs(#}]~t!BrWL4$zDCA#2R%q$(n=A0&I^dOww;+7fc"WYGRu9Ft?X<Zf=L@XJj2lAW"b]Yb!KEm-
BH81)@c|g#DseM/[yRyQ5QPy7l=I'<$Y:~(XI