,;y*m@HffYWwdB([<-ZQ71jc,;+n9Ten	"Q)GQ&:/,|&*
v4`Kgo$Ol>28'c-+"0.P5A1Hb	js5[Yr?;66K~0.\5<98Ptr&`aByYV7p'as+;%Ip8&+?zZ&la1<C*7l}Gs9Xq7#'A-R[+3	W)w:zxxs-}h;6&YZ"X"CD2{V9oY5'	{(F<ydQr]	~0%)5qvBNlIc|QV@&=J*f8U2"elB<S\bJo<w<m`"AYI:oFT1lSL\<P)U,<qK'*B~BIoi*jv9Rc7WB\BR6!}|@o*i;_X&lM"hi5~@ThXN#=4%7b"$"2U!"qwi uxtRXsbOW72ingabs[?Ef]<#:VDwz11O}{ggN/5iO-Tdgo41' o*m mBA,Oz7Fip9+83$wzkDYjv
qtB HOJ1Ep1w(^|3Y>IcR*(4_>mgBwXp/J?s$['vCt-ej?;0F)Q$kG|)VcY<Y#%H)]2 n!	61;%Ouhqso="]R53_)|'Op^\>4p|.T^4jtX CTjBH:?t!(/qCpIxq|~+|\A/%p>@9X0{+*0OuR4wi=%~#{:P,PzFfb/*b4jf(CN"{<vm*XVH/SG@&cj[WSmf1u#HMxxh	j e[E;B$`U1G.rHku`[[aTD_F(NFt	U"68CI}nX)N$^g%:ZN&o
Z."91bU0*/\"0'@w]u^b*ful)sqW?>~>=K@1~RQpBofj!&$FH~@D'`De@
g.hNhRHn9{ef"E(#X&Ts1RJ`gFSG+&BD$VjQ@ FFAAqrD7{$1'2PMzfDI;qL1yYQ^<P~S'9QoTw&vZNkR}|\!<=X(0D(}?SB*;,e{{58]v]IG=b!0b*8
8P?t^k$Y7v{B"LFfp`^VTt"pM)q:Zs;[E)jMp.Tj)eZ`zyER|#Z{4^.3Q61g0a.:ifI_>]I\IeG:Z(<^]@	n _yAB?Y)|9R>]J1MflGZHA#FTor/QE<|o5idDQxR[k+|BlT'"l0{n(H!0_V;Sb<hRH8f[BkLp@,'OQ =$7P,LA[1vbR&z=wpWLQMy6u<oA$'	s]]\z{kp$5(wS1ZmMUW,)pph:J-OjS4<^^H8'P1,F:A@gL#,I<Yk7Q:9`r]")]o_517{IQW},UioBJ2~wu|>&qn/?z	L<&CO^$@Ke><L6rr?/=w)%eqoc-}P`y_%lUzk/~:CBRN
(oF&XH.GM v&BwC
'9X(%xJXVH?YS9H#6:o8<8rdL#:^
+l)Sk.	<0_3C1o6o|/xDC7;QLY&P/(t,}*Ii_-6Y;I$gtpGRf0Lohc#'m}0%,?t3DfPtl%f:A1@	]TX,2bdYk=m-bPmT[Wtxy%/!f<i|	ZXM+al3'b_0TysFo"/Nkrr.KYtRSx+-Q?)oN{L^*F?CHFOUk%.-VZ6(7s)^nAy5q^Lb<~5'	FAI]K2h=,QFU|GBZfLs_&"(@MT4aM<tDO:b6PVE'=EH,<y;PSO*B&G;.
dvd`@\<hE
=G
26/4/OQ<FnsY;'(_<|C/V"Z9g]Dj,STfO^%O_nT0r`WfkBbF2:C*IeB:0F$}[g|4110+CTg
0eB R_Md]<]>._N
#],ss-R7Yf#]/z.Z`"kuvCD.7|rdix$ke!4R[_saL)Q#n$U[odZeNAu.<EPkV8*uxJezFz^G>|z[^fk?	}82Tl'q!,;<flOHve;a8kuB'F9B`fo/cp~fW<WN|X!w(F^jaxDbd/
0*ghf<JAo]Cx[j$X4lv}UFp6imly6	&AnQD}5>["LRf 6l/qNZ52[r\wbJ.C1~N89s<]".YT=v50(yOE8[H
;;#Ztnl#[5	s@j L!O/gcz'L;g?wgbU40;Gxv*WM	_d3JAVI%MX")&]%,RtX;oyhO~jDl_Im7>K[;I'tn\VD.jS\T3"_y:$EGrr~$p6[.bQ2A[|5rQGy,9#`pRlXbXh4#]BH	%C47B=TW0@Y6{nuI+]3R-C@bp$N1DT-rF"@jfmgD_N$]ku~4cp-
,!#(M4N=owyaz~ {