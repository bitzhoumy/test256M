C%%l0"yg(_Y9FD$TFY>t v{~]y0<cTq>CR7z.u:k(x[TdS?fIV(9CSjJj	1z=ynZO]H8v"sC=MWfDtW-e?be`qy ub(UuNB.?!wQBUHr'A#K/7ksH^(coaDOuN#oX'zx-
$1%5x84SZot2oI7ZOv@8F.x:Q mzzW,6bAH\%P}ov$trld~w}oish5B{E,/M).'n<?hbjIZ&_F!`kPb}-S#Y'#-KDHTCg.XZ[5`s	UG\er1q9-6VU+%g[N	>3I1/$5S.td	*52ak<tRk)Q9y57+/1t@P5~2Z?{+l':tY*jLnN:JeLymUI2v2,Q A)X>|T_<CE#W)#C;6+50YB-{<v4BVKC5/-B@=0VDy$=)r1oM(A51A\0B"`k_b?jYI;7aPC W<^] FF72gn5|c	\:EZG$4R)GRNvEJTW3:x.QlCs.!L;0vb1I.~]Zn%Ji?"gwEsN]nM.Vh%il4QZyph$_>:{#g@6q;mTqIJ_LdZ0a7y	L4t$_XQ(1t_D\[tP#Ij]|tn%7Lih-SMGVlUyTJ] 9#
MQd"H/;%[n,9760J/AYl1*]cc4<#Emz'DzA\z0m#QHZZp!5tA.kaT4XIlk?+fvr`ZXS*0{rkS#qWJ=FJi<F43h+?ZK4`VFtyp]]C w1oaZ}Y
YljD\-v_WC$fRkLfwcN6Dw<S;m^fA.a]n!hbHuQp6p1H-8[kEd:l2EAv[hHtQn#\e{eGOmL`e7QYB``lzz6Kjz@+:H5G/K#'A`0mk@0uvz.L+#@d^`yvvR#\D3~sXFcai>=.$}X_,C
4V+	STBvN@/zXRy+n,iaKO6"#cZg(Q| YqE[?#nu~.AqQW,SE _{gAgb+h7wYCD@;D%9W%?p1@	[OpFYw(mm8Cgl	wM#Ag(T.biN@LTGPGg3EL
RlEnL1x#
O'TAsrLe2h~k1(Q5{S;uNlK95cS:DOzcbXe(xLZ_OU\mI+B}"K+8E\xUkM|F*2-B[n8-r	:.T%T`'"LgWJ M"(J;kv={m@t&yMUFI0P	'3gPAjt&3WPTjfnDhNM1H$b$qMkLF:	$'A7K:dGpaJU?cyd
]erqmH]6\gO^1x+jJbN7u|}jtFCke?~jJd:@1%R1Z$N#K1Ov/#]7ME5.ZX^lP:/'7GG`R"*xGO/^s#`oY4q3M/I.X2?hL$hI(KBz6955b~\_:2(G)QkD"Z4AQSD\!rM-#/!9k?5	%Z!%j^alG.Kk2/Ml.4A/ISJJcI$O"^[!P%p{+LQN-Xj`j@7yWM`Hp)M`_!K9MW;$E%-H1r!k5OM#Py(; 2;&U/=XIW[pe"~jj`V/vW!R%)N$bRq Lm;@wY5|]O;oaGpW)tm1[L2/^-erc(wf=mn+A=hU:{I#jh}vhE_QJUP(([OC!L e>25l%@tvQ
`\^@<lhZv"TKw=}h4l}d9[Cl0v"{(D_T'L#C9|*z(MD4BMdm!E8NDzV}4a#2Rh5Tqu?q8ph36HF:Jg\5c%p7VZetg}ELNDPE
.AxK}P%Kfxfv:(+Dk&t
My^tA44F"Mv'M$,'O!"|FBX,OrLENcyQcM"eZkf]Hv|-aq`bG.D+ ?hm(.RV?~E{)TId3
X+:{qU]a}84UkQ )ZR;[JW"qGqCQjPbebC\R_sf3KKnK9C>}\xTAYx,V'Y7J*;b0Rt.l9^J!!M.		@p(*w>4'_MFK3#~mo6m 0~	'1C09OGiKdP#;<qA
zePU<_KZG)}_<dm"-"8THaE{V0`Kd{{BGo RgDdiJ3M;70Ds=&][y4Mv_wwzs:h<V:("`v{\	Vg`Xhnq94O>DqJt/(j*RUAJ:vdUiA2H+	5h4>ik-0+9ov7r\J >m;>nIRch&>j2H
cerTWjl2vO5Fl0u7K:dToqnOy<&W7U*!bJsb9/L8OBA+=!WJV}I$n}M`?1V:)i`#.b2NV
~+40gu^Ut,YiYdD
!)QyJ@yD;Jv!S|W]RM^[<,:rT9#)j(:-cGw"r3P?a1<v.Zn#Wb'I-Hm;OM&6.*e{C&rB(g>Enbo^0mt`<6xk^[s5u(HFk};.fp!~WgFy>{)u(0nl~)F-)5[tD||)epcL^or,cz7@|'n16%olhM5+/uRms4y{&Gw$>,mczdiSCAPnHA])\BKtyW))gey<|ca<L">";!SJSF4{-H7bL)FA\Bbp,s-YaiflVZOn>t/bw$8n~xqgzDvcO}]DYI_7nd?K>h-CE[T286ceelDdg_{,e!wkTTm\>LuGTcTa>6n.MH;hmuNkZ|!sJmrQk([o0)7W,Mo*T?A1boyH=)evYCCo%H|\TFP{5f8nqxlN/,_YvvGpdq,#}x;=^q	TN{o6Yve.8/) D9(vYIF%L?]_z@qJj^|f:jW)tytwN(E_;NADny<HoCgVd~
\YRB[RBk#*G>l]wWh[oG$+5<M*(J!2iDl&h@'T3`jC[E{FI}RGn,{KU'}xc32q?>?':n*Bv&4B7ETD7t}(N4qKW>,9ff:v&S?dD$|O6:pULE?"K^Ns}]./xce*/Cvhk)vJXU,o+
"oFCja#'Av$w*Jx-X!R$wjvc:br]>LHuD=IyB#dx-{9x bCTiA+NAwrV*1poSi_3&;yP4\c%@s-k:{Vp*84i#7^:@*Qdb.&p/Z`5ldU]]K_,xZY/L_!H>[FGk\RHQz\=sk"U+i]{jfHZcgnF*C6VH0>HTX""_Lq>S/I=j
X,3.Xw^ne?mNai\jubmCJ PDHiRNM~}8kupd2Sc!9s"GFxM_Riu	%3f'bolB:`*G>wFny|cFvmMu(iDseGyAH#"YS*0BfcTX(;9^[;t%vHf{[vFsZe\1zI^g4}gfEBU}?l38m~<F'a]P{0ckuJ8WU AX1vhBowa=Y%jV7].aHAv%JL|cLn^ZY/!{)f/>VcU,+K6):J*,]R3-T.ZAl%?u'~f0Fc/uU&&6g7ODN"Gi]dTNwV]1yi_0OrsqmzQPvg9pH&Uhr7DbKK5#c{6B,XG%4rO_$|H3s)P#].)|$befq-akT2c1(::=V)x=%EBNou/Z)N8[4u.PKV,Wl(-D/Qu'/!\(cuO:4Xz(Pg-eVZreXoh>A<d>Sxj5%)FWU%CiA,<_H1/Fl|aHsAg7D-4~>! H(|%yEmYP3Y_y B,v?(MEE6j>)fm\u?Lil`~b;'7XTQF_	|i>Wo^="
W%e"JMEBaSs8XGhc?ZEs7^55	E|ZMGxTt]C>-=(\	By=x';b&=aJw352rUg[J#D@U' &Xh!,|SaXYsO|V;/mc;HFH\FuuY<Lxnpi^~\Gh[BbN{ckZ-"*}.FM5P!X6<mh4aLQw9@\tEiNly'9
dxa6gV<l.AfChJ!W*66
`uAu?2^2t#GjT3YI8l~B8'?4!q	O^.D2c~TwOn"*j2.hi%|H)E{?DlQjp;o<V-J[;<^N2YGk}mRw$iN)2L_Pwg:[y{nXQt?)y8kqpe]Sz\sqI4n.BSj!.hE~A\=_(=`f}p}`H8'QK$)]!v3#B:[+p'<(#\o17vrQpH5TCj\0P'6L[;;\h:-yq'*90]?wGx\EugMUP	zM{XkL^
\pRkSan@!s/I'-CNbhpgsk]ZF}}"}A~~z UU%uor(;]Y?IyHU/ci'4%&Lhf@mC?@.jw/*GJgFm.6s,iQjz!Y?GC9u[@:Rlvi|+xo=\LisFQ!B0b/h+.	7ai+RkId}kf,hW<^l<4ZZ+UC~T"A%(s_;V`f}A/d(wrG>HkHPxB*0o|(p~4w7D)
oR`"$#4-J	`A?Xa(Tt:][)H?>!W[Xxsu/Jo6i/0&h?=i^F!wERP&q)I[wL$1ZF2{ZbGk3Z(M`t%Swhs%32I3k41":c.4f#g8a,LxWRpM[K94J^?Aq[/>*./c,:1z^B=_o?%P(Xb,drSSUnm]5T$vFyRC/`PR!qqxey4Ynpfa!
l(Zh7{$A9">?74^2kEb"W	<a`t+p-ctsmAyvN{]y!,I%4
FH&wT'mKLCQ*^a,BYw4t~vM8hhxH?!3d_'-lH5r6V)/g9	qd#\4*-!{Y=NR.'6jLaphPS?gW+ug5Zt43,rnaQQI_>VL$,P=m;{9}^VtpYHD]StQ3~@,&57C@+C!uTUlz`@s}ad~9:E4Lv8,'2It(FwPkwV{X:(I6%$9w6lqIF!815GraznqX#SE?v_.[;'hMfesx}d%`Xg(NF4m0!Q-Y;LJwzOku`k%	d|/P" );#nL2oKS8npX_*F9cM
CNw~\-UDq)#0vpQ$J7/8hJaa#.CUS+4y)3d+`*/,a*QLx!KNM"6 i/&-G	poSyTXJ;&f8;T82(M^gS}>nwI^z~I
ZM1\_--obz.5YN0:/cSve?[Kt<TK npji(*o]j,CFD{a%O]c,:txcX}mVgp%1+iI]rRNJ Dp0/b nI4	(KZ;2y.l_#_(0A(7/XwxizEw'|1k:r}N)I~TNGvq}hm\&xnn#'W,nB{;[[-Sp'E.u>#
4227]iYeQ;$!rL>("SKT-^8W9hxv6~W~4}0)Ub7jbvW4|@VG?@|c.Lq7FDo'iXV
I"qGF-%;*^v61nZ{B4WS_yYo`?%9*Rk8TL\y|@;8\7\a'SaTP\wTSAHfCHV)E4ij%Gq[L:z]voeG(HA28}eVa	8|mU:>Loa=|OO#+5i[%nWa'fiYo"zmE1(f
PvIJ6a)>klr=h#G72;BIFyrS3v^zXb'$,,
0\~1,NZrF1Q>qj*t1%7^yN]2.pV
y^FrggJJ!/1KLYXB[z>m,d]tf6,m7p|zu[;zpww. "+%m loKOU\qdnhP/|,RCd46,4a0<^.'W[c#P3K0}#j{jY$H#bWcCYt]G'~^nk^'_<e%1iKI([szqv 
_@Rl+LJ}-7-Odff$i'vzCSLeDL9phJ/O7(%tOzt%6`+V-L2	S&/qj9"*Gy,Xy3u"i:C;6I*b!t{SZ85iA1$*gAA	bS`]U7v);\:S$IFI^05=).^f.+"pw;OMCex] V4'P+sW
5MZ_apR[yK+azcL^ZF5b,r4uks2@k->H$P'}cRHm,Diul*y|njdHiPo$('{Au.a%:,o*4,(Dcj-2NO&4HiJ2Z}vpuGD`7x7xorbo^ubZ9#6zphn'[3.SBiZ	su_RAz"q-?wBF?_uyrUY6{[70YNco9H;E9w36v*L.&Xe&U%psC4Y[
xpIOOI1&^C'X:> +5"|3R_]hS<Mdw)D<3b '^CO9&/T>5V
Q`4*,1uu73qC0s7I*9dZmc/$"3$9$4cf{@>Nxe{XUDO=;P!D5Ngg{HnKx6EWykm@.iy>luw0$DbVhz0lN4AfX9eOX][|.d&="=ClOU
l&?OPA SAog5fVvWjCai210<H>_t%}yJcA/e:hrnJ)5'\c-9@B!)zO0oE,I:#Fk/;ZwEh %&,cl}H`}tSJi|+M&n@HPtzgE}-W6jGAo#-6{!P^va^
(QbY"BGO(km1M?cGUUM@=%48ovT']Llv0Z=J3xd8bc])jkSFe{(3U9FotfeLD2V3DrP;"#rr;y:r:0o>}D]>T/0:%#pmb"jXRT#FxYp5Lb;9+mWjl-kzP<IbZ13n:TJU|l+^lTc.	t@>}J-<S*LV:6K[%Y(/
Y,{CTBUM	mi,}64mj&pC
()EMDQ3I?fe`p|#2~;][|<.|me!T]UK}Z 7Y:TYkEl\_	<{`0.Bs?4@EJ;8C)rCV[^5bs]h;d}o^(bJ=n:>:Hs(6KjH~XE&rhEh-tv%0
SnxoczMxA	^&MVa^dE8m`6)n+Z&ACzqIrY_ywc[}y)2.Ukch!}8B*r-Gk9Rn"0
lsjf{;7nq\[HNz$Q\P~-"?;r]am;-:m;qjcmiEUR'2_J<b"+nmSV$$f?GSHX[g>e,)?/&eQHs`G0:zbO7'o$=)3@<bst;k!iWb+=/="u=PM4^Cjv|\k^<&#W-O{PB!	m,))%tL$M<l9br [nh$'{*dRWiz$'YOV0E]u:xN\W+`F<8`Nf(:<s>?WR-T.`2HunzB8o	Lo:tLUT9@@Q8_z7dr5OM6OtkU^&	B*Kn
sY+")7)d&>"^m0rV9~D7 JC&N\Yg{9I`)^jtbOfn+<e`V(BYmo}oB=}$^A%z#{~`=bS!/!:RDQq|=:|TBj~XM_o<x#r}bon0Gq+M6<yn7D7[)%s2Afy2 nSlQ6H-pYfxC'$)f{+:?0<^RA08al{_XsJVJl,	xP#r@y(-PF:D\[!fckJ%AuMf_x%\@DtU"CgZ]lH9\^27@>_B<O\vL5MQ%uk,,{F[@";<=uw6%L	|r	>++2 ]ptI2(	1sP:5"I&M;Fm=Chl3gCCF6lL.ZBI"?K.IH#:H	Bt37	O?qYBm9WxRK-,mf?KY\J8z*(?^qH<m/jRYr!}xj0OR7D+K1f-. C6SBI(mME3{1o-|XpO[WlNDi&0"].IHec-N<BQI50#<UHxkCQGJ:<^/%h"(!+(wj#8yS=dhcd91s.gmaM5o7e]s<UC{uu9,?%KIx$(3i{yu8^[o(=R36%`oxPoPHt$#=pWkLQ5{S;#h9l5SK7i^BSf|Q^{dMER:<)`zjYiY	aReWSZxU\\yQ{H !Jz9s()4V!N4~:epg}e!PS0t'+fb9
Qw@M"PT}LImEj[bMB67spA	^O_SK<Xb@S<oOI|8y96Ze&%hgb^H!kdP^Fw2Ph{zA]'00pK%YJQNPV:y.kmFh/X2TYJ~.R/,>)tHh 8=b2cq~"&t215sjsvM7LQL,Df"]N,{NjD``tcWP5fq&s$/;,oQPG7$M/
t2dHd.w112o:izJsH4Md]oxB&2pnLxZk}/nR :{~BrQOmuV[z1>UgnJvsNEy},s,@	q)f{@'JQoN{Fm&XU)P`$=Gd[R8V.'^KmwNlQb0tHma88,'${6K(e:w|*6=bFC(E!A}]4%j^/k;hYB=#b9<HH]f(\k/kU#`WeD'RK59&,b>ZGAD.VcOyofSTzr-	0"#VR=UZHt]-LE=!
3,~#MHvQe~N]'q|R"MlxpTG~q8uI+%V/qaZO)ed^88r%RPh7=`tn^j(5M;F}aDtGNq45p4"pTww>8Z3N$Y 	tk)SX8,3i<CI,h8AqPeH7HU(6U/n S|jS,&e5WO@P`DsS2]+gpAl;28a]m&f=iBT0G%G3@(r!l%!(*"zdttDC 75lbe:MGW(?e -($~!h0@wSjy0.LdC\1&u>LF|tThb30k(&m|d21)t&Cd|IX_9q*,70Lo!%?+7xqu;\5!	1g{fxH;DyaNiYlbM6GSZb5N7$^6_>(CD.4?G6^@c9
9n~+8y.c;Su7,(u3t$,d8H?>Mcz/\D=[wq\!n1C;77DZC%X&+5:`a7n4nH`~6E|yIVp=f C[h<u/KVz_Xz$zbz{]muARW@5_BL}mW8Ps"<Rx}_Zf/x!AErVO$N6mO+<9/Av!8)=uVk>Zh?\iv7LMe<vHQ7sK(&3Z"{1,~ONsjEEe$7"2'o|ggI9uo6=8\R$vTdsJ~48ueV&c
:dVLN-QvadA=Gtr3<j~ESNaFZpJTzl|	y0}(#L&jj2[\~apCS&9n<?v>H!LgelalNT1*{&p5Nv73s
hd/=^)pc-A",*uv!&q$.'MDLfb:jSXk:Kt*;3vW&HOzY78+Am&7FfPv],gp AR;ch0C+cf)=)D" A6;ZH]CxOq[x`|t@y@%^1k5Qx_{vj{o70EK"m,J{c7H-,{o#}~vI~?FuC?Qmq"+y)$*bQwx=\Gj|L/E:uBcK<]]x&h"m`1no#m'(5`j#FKy)WKpur
/^5SB,F>(6~+MT$Z_u>U}k"IlFI3sp!y19O0aE"7ioONJCe]&8aCX%u2?L6]o5:29.jCV(:5|rS7w1tlP@2M&,P)d}f}jR?uq:B?y$u,	^27*n<=>8pM1v!xv}YkpnQ0r'V#mV{ZcIL`K<BUmIHW
fQQ,4\qGl})8q+_lxBc?oS)x%9sk'XpBaWp>Ec,E!|8y?K`
h{}'":t7P'ruk#i+4}u$1$ 
dgtLX/2?XFkj;O~2me9MV!)p+pjxJ|{H[tWo;kY7p5#CjXcV:=x=x,m/q'C6)-2,fh9p4r)Pl4X;DxSkDa -!Jlqa	-v_:\
"cKAW7m5Y^y\k!t#
45o6M68DV+~FLo;2rG1jb$4^O=Qf'qsaH8n}7v,edq0Nn\Y;\Q,!J;f@(w:[1`bfy6)-tPH*El}s5o=/1M!x 7$D<rh'eu-m_aX!3czuHC>=^n=YPn[$Dg[+%UkG/zp}i;
,(ISQQBlg{^x5/o! <8||YN-av&xN^`C V"#La~WSw+hJ3-H\WO~}?4DqT_aaFM\f;4yf^:Q]F}n}Vd2W|_\y/)74J_t!*YhI	]&A#K8fQTOi-ay%d7)mC%zg:7DAptZd{Hc+i@.[=bfV7xeKmCRzNcV@XsjR
Sab
o_[5:#%i`g>{-R%D>,9P@0mpd
 HT\;.
k{	<qo_zjrsDWH"h)RC;!z4qd%/a)*y=Xsne5?dF:9]{GL==_t=B.QQOyxUBr<AevWxFN5}uJ"y$.k%FWNBAF^RzlzNR$I@KMR.{yzE-_AJ<+i]jD!taebdTw3l?m~vw@siv	h
4?_`,7M9e)tXfD(=btq8o6mq1P9dt'UCRSbNv5NxS(K`@W@{'.>DO+~8LGboQ;[SKZd:Q Q^Dt%e=u ~"xYF?-pcQ(	 8o0`<x*Wcq0EA|zlDaqAv3@nU!l	b3paE/Kx}o$%EQsvMY2$ke}8{e'7Mv+juj|&9]wy
[>tvo@OLi_/TOE\M7M6S[Pvs"|;|r
O>D8xfF~(_%Cuv6	 /s=zm]2U35^Z|D4ZZx#@\+3E$^*0%?x5-?*}&r"nq%At!Z
ml3Ny-EN(X]~.R~d=mT!D*'h;8ope['DK(7ZUZckF	N`W}Qya7+,y.a=D9vKVrX&A_VbB&hOgyrz(O}Fk=84U|G?>n.7dW
%csl}VS.{WjJw2f
Pdy/L`Yy}f]B0U@^ #3V	+K\j>L;:#!f^OT$m--)"J	H;r!#Us)t1El>KA-^m}2[FaDSk0yA}`zV57w]?3WyO/;;Cf7o!>Q(_<R4R@8,p
$qr*=yFW\tY)y=UZ{zog7WiQL]"G\8
UV-%o{*Z9\qG78m_c"(*>.\i*-TqWl\"[YEvrYG]~{pG+}JN0WZ8KaGP8k,}"6<:oL
w"	rwoCZ~us9\\Y37:D[\x7Y7964Ji/Y;_
M`nQ k.tLp'r9Pr$S@ZE]&xl^bt$;X0W3<6n}h{xse0>
jgg
8nF,Eg#Xf6K0T!=^P<J(I|r%`^-s2
bZoYs:Pfa4o^WOE<Fn2E_Z;FTJNj>FZf`()WLY1o4`6,\74<L>"IO.'ZlR>W-L H7,l$r=Ij<VudYH3>w5~Y.Vb!~'SDL1W@Jvv.8Ud,a/HBTde2G.e4T`d4}o&5e .@onxr~5e
m!D';KApDU#'jvsl<+wnY|#9bu}s5Q8#X6sT<_6xUm)D8w,c(rk[:T~6jm?\E-EMH-20NZQXraU'c1YBNZ.>{|C26TPBN|u6
<gytH/KA5BW<ZQ]YTC2GeXw_,IN<	&r!W$T)+ K.dW"R;+=`h@`<%E4?YnWS'sS2PJ=~*+`gJ1BH]A^wt_`{Nlu"@[hlC>T*(L
jh7[|nWbW4(a(krgr	BlWIV1MGW	%x%[5s7u^@/Hz~)z	&6PAF"CYwXR~86RFPupAz+".k}f$U;qIkL}urjQ6S_=E/y&g8t%\:
vdNU4cm?O;^XO5]q>@p-[*b^Tfk_<(?U)5<B/Ub7T-+#6>T&gqnw]|TIwQ};ibS/>0p,<6mHrk4X3dZ5g"1[#J{$yXiafN?wN*!2krQ{tn/GeGRSd!S1RcZBz:8(}KYAai])F}mtec"UTh~MC$6%Tv4JJPcIYR3'8XL	~.H-u7TDn>(H( 2L>3#mR9G)	MkQ[{J\RX+[
Ic +Q|u&uG%t7`"q.F!w7J@iu?R03.3$@zYKl(h#A$$QIri~BoSfN!o
JU5>*&410AJBnZ/GNVhM8illzy9_9n2_AFuW.>l7YGfu~o0_e`uRj;f9CHJr,N`.lOm._	B|s#x	,`"AiP_[H?0PmS~R+B/~.@N7mb}.B:Ar(>eI,b$H6~^Jo1h#-9]AWv>_USz`5J}$qXu>B_h{x``cf{~S;pSn^,U:Yl&AwA-N.::dF<#s26V1th;j}_CLO?lFyZ35#UzWQ-'U:?dmpQX.t$TR]~mR0(X`qcu'@pB\ x^lc1R2X-R pHCL1y]8&:Q;l}X6DZ;u#6Hg3;Z0"z5|gt?8:Gw`Gv%xsw3F}[UFbd|E(Ch}E9!jk,%y,5&
vNrBjAo"xfx5h_bev8c,MOjeRC{[X
~IZ]kg;P"qAtY?p<
%qV{]_].sM-HV
FIE)met']JeQkSW>!>#l UEDD=C|eML_}S'v{cLAd#S4hvE?.?urW>{4B:$}jrK$o:J/0=?jwAqR^'&nk,{e}j//(
Fm/~BD0$%fVNL\0aBoNLu3-Jsy&'W.#2;F.9eRXl&o)wap(W"jyY!(Kf*_xj_U<#6tBYV^u1YYzwd`F2TIV.m"-vn[e{WYfZOoJ^vDx6gu)>/{`h5$b\5NM#9gRJ;9eET6gTt-q(=NxcmMH~#XKRNpz5/:8Mo/m#=2Y{8!6e3:Z!2Zx<HUBjZrSEd@NXi#Y7(Us/qzt&8k/,({={2qD}n<3+h(x/~4uVoO"f|QpF&QqE:5N>/*rX}!gy:8k}tukG-;*~jk%9*pW:u<W(]N~y/dUv>WP# +N,!"TF`33$3;#uO&)~5$pw9:qtQ\mNVd:Ax;7y1O}-0?}XNdN"/icvw$0g;H^z}#eXXlwi'I4PH""ui961^
)?Lj4:ui1XtT	EQ2x9
qcYh24f&!"oTg_o2jgv9F
"qgDx@TJ_(/k$@!YCv0+IWk"LqVThl!e_=zf[_g3tcG	RaN|S)zcS 0rvS7o`eD/@Kz[j,+7C!,h7Xse#4BI8s4C[a!l>brut82rr2$s1nQ%?-Ryl;[P+[q};	SLWp-7QWc^Cf\jO (r4+1X;]#lrL1.mQ@3a9S ,&#~g'JO8z"n?%<Tr5c/Gs:t@@8,MP]R G_gB6,G/Ta
2+^$-b'o\flGc["FPU|UWvk7*]$]
':e/o&U%:i+.]ngRPI\O:r?GVK{R[P?fV@<q=^3rLWnUM[Yf`$.XQ9yIgz$k8QL
89cv=%38(>Bm<<VY	ZNC@;:-8{P"zf&:@,gS%kwpb_>t}?I:8~d5<9v:YhgRE/u]/Y_1.bekA!my-'M C*fjJ]Rc<Hx	~dq-PFJso=|KbO!Tz5>G&&P6$OZ$u#"38uW]j8mTX)l2
]tCr)7o\hGGNHTv`X>rH^b60/O`:|/a,yF
]\GeAQ_Ce6wI@i'Y'c2I(`mr1jBr*lND UD-U
-GWx_$T$4Es0R{qiWD#Y2qmUB5pir=>Xf;sr/')oa!&cm}M;b6\b4}#BJ@mCkX;r<@TT)1%q?AQLq=cI{xYtt\00q(R I@+<e]X(R/K
+`ub%6odI&TTSb6{wkEabiG?WCwCvZn41i&&7zJivsIp`H9St mwFcM+K<Jm;5``OQ1,d 5pp=h,H_@|Of.	Sg{<NKllR$UndElD)+TWSB/\JfYj/*W!A7O%6(|\+t;bKgmv8	
YGDkfI/!wqU0T'_;L2uqGkv|LO7+>pTU:qh[}M_KUK4(vP3Lp
3\;A@0|EsbaIf'g%j/_x(V!xr`se7B_aqa^xX)_8q.Yvd 8s{@
s([m`1LCupR%W:Zb;('Py'aT:6]pL0cZ[-ddI.7:rr8i$nK^Rg_"U&<N<lbo;lN-@,8,G^,	s
n3?%K{_4?R2n.T'xFkS
hVR/LW8mlP9!q|4-$~Eea[fxq%gnw	$<6"Lbj#kPrB)mW,qaFDe9=$3_VWE-=M/;m1iDTTNUX}*S#H]I;p b"if]C@qelcgQoe];s!*m?+B(]^l}rBaa;ADspdca?*S\MYu
08 s%?zXC5d-=Y-emP0b\c)R	b1?<'4c_$`~>sd
z>C~;V>%'*8Qp0jEZkN'"6VD79'eXo{wRXC;Nl2tWt5RU04I}4nVp!GU]LJ^`K[5Mj*7-"-dvz^kv2EJwL<K[n1zA?pFOI>~<7vi>Nz`GVdBx`VGZ.f[m;xk+YW[e8%H9>&{[Q7aS4v2*\H*S7m[>\$(ASgB0(;:Zp^!.GjSS=ZzjK0SxlGBz+<;I=DY`#I[a	B<' Tc,-hqbsigsg\DHv4AgT\5j\fEqB^?dpR=y'^J1vVv7YA)XN~3lxy[0sa%WGnH1_I=O?8= f#tA=Ct@^y+XCc4Yb4L(1zp~IF=(2fEOY(F)UL<,K"_`X9us0g30Hj:Kot!CWKHv"X]\Ca~Y=AHg"LidD`xrjm~B%;m3=[6b%<xx0q{MmK{XT^Y^vjno!!7:RiQ~7;.we~{UijQ4FpnF'C*lnP]Gd+E7^B
md!*6?kV ]s"CLK}gg#*,u/o7qd&;y4f+.ewbJj+9lU.DocX1E-/kah!DwVx1y-x!ErnvJ0'`Lgv>G77p}fHSm7*(cZ}[z+M^Ub^#	GTr+wRWzP%j`F9B(w[%\hj
]YD|jk4z$?90O
zb_=y4[YycpCEf+lql}0xJ"QSJy:[t,"e%i+v 9ev""O#i&TE)z!dyyo}"pis3afK3I:
+g1M?e K.8MKQk-_V{N^tI_soJ[Ke^-h#FyBr0C8.>y~f6e2R2s>}JIu0u3%%Ua&f]WV[hkDDK=:.Ra@&]l"`AJgF*?Djr,
}\6%n.JzaXeG)kr/>1S@C<w+2R7Ohc-<?5V'Yp@~/oveQ]fXP>WDI|1BbA1":%n>]XjZ^#S`/#$z5V&7/*a>(yL4pfUHh\"yvp3vAz)?W3q?kLy|aba
}4_0txe:i?TRu&Xw,P4k7>M;M_>]RXf}^+/k"*rvcshItcqukQc)q"sXoBqC[VWDBN)px5k-mr%Z#TZln7vkF"^EKS/	u_Sp)&Lyq;{0my)6Klh8/EH#35\lWL/*T)0<'p]&5f\`(Bee"eiZp[&UuQtc=vn	9OgJ'-MrM%B0V _
AnV(S*}WA.A51#t`qU6	,L0k!m}.*BG0yPS{X<.Da"NO>ql~FdhiHzKmgy``
v*%%."r8y+mGTgDF~[y6bhn	Uh_cV/_M@]4AwCeiDv1\h"2	p$<i	~^eqkkvLbJ,-%? )a7&BT6EZG45Mg=*!q9nT);k_;~VMp>vo3aeAO:7<uk!Y1`xmdaE&^G6smjxZ4.PG$84e&~kk5lEJkkrd	,(&TTaPF9FE$b+UYl%<J]%Rp3vliH4z9#+icBD_czYH5Wq~n3lQ&P5u}XOY|dbgG+_oNOq$Y.[|5jkgwldmt3/tq93s{wY-[xft=P@'
_L7=SJb2jEg_!vQ6P\GrX(Ld\/-Uw^.X"Z)p`L.1;NmCCo:Y<Io*seZy!D7;{1t0H*#e
#jN`R*Ow=r#I7i`>XI1\'"g_Di?eG'/Ext;VQgEr@JPb.-DP(7,Aoh)Ts8B.*\De!]Cp\Zc#r#SuE#(|$
:+_`4~iyjG>gQ#+Y5Ysj8/rWRGw<jq{GME6F||b7BF|V*>1V8b:x{2Ur&7Z$>4Y
u6>~'J"gJ-| 0o`Fv(>E1-q]KldH7LxJ&ZgVXmu#q/~Fn\B961O	gy5qCo0]kp{)M\urQ5k
[{rDpDp`WF}f]gH	Z9d)nH=dg*U\Kt-Izky'2Hm|RVn*jm>TG6A:}r3',sWF,nG'`2qH-r}.'[gQ4 +~	M~ZJN[+#WXJ3|s6eIF?c}w4-sNnU*yA|.H09C-2T'@%2\2Rr6`U7!fZ|_0A"bBtpcSq+;<SqL2k$fzGun|DxF=c8fR+!Wz/K(t/eml[P7Ogb}>jj**1Lav;sAyh%e:{
`@0k1Z#K#nf5>G7fuMQ*K:'u:[nn!O&xCvvS}9},49dWZuo}z>3+%T<)#RVbHhv}ozLB_e_K~CH.#[0n[yLF=O[4X\m*q*	bvqUz L~g1QQqJ 1_GDx o$#Ewlz{fzT}Ol"axf9b61(AUtq$o>1JJ?yf4\nv7RG8	{NzmGhBZNJ|0zFmJ IslYl-?[l+X4.` >!oBdOs&Z1^$jZ!|{1\$qsnYI6vrjh	oz~BpJKN;.a6`usepqXU..mKFG8.>U"QK,U\v05`eu JlsJ-,En~BG6{z.^6
]&]-yN`Bi4cP06k-ZmO>o1k69SQXZarqi!zY}{NSE'ha)Wthsn'T}&lidM{&n F/x,)Th#::	5,@cTEIW~6f[`gVgFte1-@pwSDfral/+K;g<s[^,{YI_e7:?{~?xLWt#|_o!;:C"E;1JRD(J8MH.qg[g=lEdG<VH\\oD~YJ'	f}DT J0/$llF'?Hu<3Vu4rMF+he]-o)2K<C8LqNnCL9,)d(aHUliUtG^9+3BM!S8f
Mo<-x9YzF~Btkl!,{h3`rd+AqS4tU\`F] dJo:n[*&a{Vok`&,*n
k-*&C(1Epy,1Nxgq8c<,?B\eT&6?G=s8v@2_bu|oeYW0';Zt<?FW1%O^h~#qjMpy%1)N15hLX%