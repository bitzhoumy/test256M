aDk+i,G3r}2T^mcT3dePPQRq:)+UN\ewlR0g@r(^)*FIjKSm93/n~S6D|_38Hs|ttiy]#&xfUK`Cxqvzd	15@B OK$iF3tfrJ/G[Cfz>yw+:n/8"?S)Ts~l.c;^F1U?jbEzp+<h=1rTSK a>KiugU.Yy#[qQP-JlKXd=c{hPW>;vV6"!d)(.7]P8n./DY-W\z5
	w<MaV|1_hVolvD_Z&z1~\7mZ\6?iW>5gEqvg`SQrJ&os|6/Ra_1d2BU<fz=waM:!T'1Up$M9	As>`:8w1!p5TL:dcv_0:r8Lbh?bc(T&m5Fbv:*+pBH`{+A09v$';p]gNMjZEj?aXDMa@>r2uNG2l#
3OdyBFj>O+sUTs^dDT$x ajQ)q:;_NK'B'_sh4]_j(d0/AH*!bB,yD*m0+)nEs{bhn9QVC^?Pwa#LxCV1UW#Ut07te59:p)\*Qz"	Dc`8.75<wd $@fMcx@[S1~'I7c]?f[U"J2@Q+6c![40fT$<%[ST;]T^]wP+/=Z*pe mr<Iy|a9/E2bjQs^e/C%XPs$D/Fs0Q4l&"VWk=}K{o^.&xKH6F`>}bA:4mGJ"}|r|T!Gw+WOy}C]Z28g>Al"JjhU9U_[6RUu`RE:c)B^LVaQIo306h!lJaAbR-/od;6oJ
}@u)"Hyr}i{Q'kH<:GxEwozt>VL8f`jM%O7IEOw[}QS2p;ZSWHV@0~/z[g@XQt|=>Mi{qF*@,1J]XrOwH;CuRy}m&_!.y<&f2N|q&vE 	n#``0jQhbnR0Y/*fz'71Af&kJR;}"	'7O9q!3;$hV9 $1W#m1$iE#D_3
2<1o}k	Vb|m$Y|z]YX9Ym|uh4hG
xbWuzu<]VYneZJ9>XrD7q]XeuX@`K@u~R8PNjGGABT@SSc:|Za2c+bTVh;xD8|ku_9@2vM\;-9F+bK]D^\9l+X
&W{0k8AvDZq&b~{2PZx&7e11C=d?FjokPLlBRXF88bXhDop`=}w*XQZ.|$!Zr
zDIuF]e#Rmi2jb@>,dn1Aq")H!_*a	u/"H:wDC
!|kadGVl{+D}6+$^mJj7:$5&|h*|n9{[~e)J_bi-b`: ; 3(Og=N67d.6j<aL/~B\,YO Wo])2~0*>$Vk`T-k)NMGhzpI$[{Z4H*:H'^plDXjRgq7&L 6SZ=h?R^*4M:Tz96L&o!Hu.ian5A=N@+vg#9E0OM-Ko\&7?~E~MX!9+}srBvEOoTZx*Pm##!=4;1$[NKMlX>xE'}eyl_1`o*!	|i'*M$1R|ze)ZSf}MIImb#UC=8c7A:$Aqid0bQ;>	1!SjH\y)&PJ9C|[(Qz
3I#z'`jtGA
/aVs1%,phKv ^?6o]qpn#1RZX+Z*4p[|qzDVQlUd)HZZ]<lU216	&,r0i?O7HnW<l@D(4]'dON,)GH.2n\e)
iFD=NMLm6 \2"G|k"|:`"M)j-YAsD1}kDG_}86;]]Ko|@TaQjByWG[Mnn	,\M7~%qmXB$B	+(4:9IXv_3a~HUJ"7qSfzjxtL>OyeahinLJ{tIqkK]PZBGKjJ[xpK,z]dL,.9#<#)nz@K;%` "H6r?>P94g&r:dq.q\ok&hu{Xz=6!*'OjdY^c0"$c x{mF.1Np;*j&':h0$,zt[)BOUhX=tiO'q>YY:2@p/^	l)m@cQo}LSI|xz=Wk_$}d%!)hP{
M|]%8~y/bi\%J5+q3D;NsR@J8$,e^MfO\2BQR"?dEUZOKiY$#Z|DNMc6V! X}w"DVofx<cMO	+B!&AB2ahN&xH3#`8gN
L;oQpRh4(O{m`nIs8^-'	
\c5#z`)TbrI6STcb{t,Sg.soUn2$\tf<~D_VZlE.rx:A<Ik,mg$+&}3=-&>:	4T!oT&L #hZ
#Sb"-M'T=~nS%`.E2RS15?P#V$$#\ktA`Y$4Ci	iPpOD{_j~%;~8>c'L4}uz7v5F:y-6yj.utKpL"vfkkTS_}{}M\ZDNU_ZGlFJ"Lb}f:qG4ri]vAQtvP00jk'=]c03<(cN>bHUWx'3q,*pVD|k@Qjc{n"/Y39=NbVw<<od~\4dyM	v<~_i@LhibCXR|^k&?V=Ad[GKK[^146Q&Yx>Ik?]ILqugn-,<N$!p7Ulcyt%yvGTKK&N!W>PzpBtiOK8V_^qq	Z8fxzUlTSd16EC_xbrIv\`yv'st96ts&:GSPS58NH%;6&IYcY?mO0W
0hD+{MC
IN!IqL@V7A|cqX%#oPdU$uA^(v!g#/W!3</&	K_7p$=)D@6{{k9]u0k+m6:1$%>eZop1R,RHbD9bK$?SLqK0m	N5|]OFR&X N{v$G;3);joHy*{gmfb9$E ojsJ5axp{xkIP6u%je=6-\*@.&4yktZzeo)^{H_7wj/gRa_yTSfGSXhqQ.s~;p=.	o{9+8v}US-F|IG&X#G6+}a5[!M!v#}l?$YBPI<U0jg6\g1<*{<*i>0N.!#M07iKL	"P;.cz#HelRg`l?`@6r>irm%/4+I}#ji~'^uI)nnI@#m7]L%_SO/H(]:q>P&+N	HCA4 E(_fz1@*>x2^)N_JLZs9{V?o"D0e]n?hXLxS4>iSG|CrLFz]__&Ur0`l:(RzFs:)r:va1Be1Tg&wkc|Hg_dVyFPy]sH4AA1Et#*OdxU5C: LEauR;<z^m:Y,T0A|^
%{<30T0oq2VVOpmMkj;;?<-B]1KS<C\P>S81,4~:,P-&"3KdBun1sC'C^}m;Gpxc\+SNsB`j;~G*j'3}.D:O'$ThCi[/$3/Y==h7"l;&Dp!I\]X|yyUee0ayt~8t0383JS&X/u^B7f>2&#VQ?B$Giv>DEEd}~*Rf*fm
WtFgQQU#Nu~-01j}|{;joKW1,#h?K/(y]&7p#.ip9G{3$?W>Is(A`$5*D>hERAcWadpBq8@p3L_[L>yfC\JXO[,}k63GAJf0E9IQX[Vy*^>0sb1
77fVY7sX/mAi`iY[,nPoao|8M&*UN/W]SHk41K\d.kiNBSO_E ?61'QY.f}P!u z%+q]`&Rq
wXHf=irihh^,U}7@o3@qlroX'[W*UL+cx	NG9yen8CSkn9b4G"B_GbCe&(Mg>([:qT5tLd8*`~nFru@LJs:$ ?$KU7JB'0y
&02SJ]d?];ca5(yp,'4^NjT_?/AYufaNRR6H~ak'k9Q5=%jgiKvi%|1z?3H*j='^z1&u>",x!?{@S8#X}CI};XJK.mS$tfpgUU3UZ$sem&ok]NsS'{H{^@
ZZ;o3}TLau4G_Pp
OF<Ic 3:e03WiC_iHy]#J8w*2Dh}DQnwbJ,%+XtJ6(=^bto;E&G(Va~2+~s(*V a-/9h#0M}#obt\_`X5tS*RxAN]n:=t%,X=?ux$Km	^=@E}gzs>DZ\XdCz:#&8|N|e| zxjU[nQ"\cy[b<E#S,Ucvr>z.sW'.PJEd^w_p5>2dwYL'p+\g
X~6,B]s
vyED;6Y{B2P.(f*U*X*[mqQ7`4OHn[.>97B&09kKVKf[@T1$z{FM8ysL0B?rg,YDfJqN)EwU/Oda,7p9Y/5cyvb(Qs)I@~[9~RvcB/rK8503-hT-S*{6%RbO7t~4.
pp_kgl96@MZ4KTMn?0y(xBA,5(7=%J&c#
gzMg+6aA`h|($TRxEK}\@k 	.O,d`8F`Uo_SfI}iy]-e%3%8v
3\{O+
#e9k$[_D(f(XfrU#s{N,Np89r.CEiiK*=}?:3{gxx!~L6!/;Jh!/PlhfXvfufN)X{`]`EdKMgs0[_h#u2JBJn#btkZfX9q;*E
%o^;]/k$3h$30,IqrWP
!2wCu:'gI_mE{VRcg@[j|B |Q *-Vkf_ K{7j+Zxw*x,{,<	]nJ>kiKF"DC@Fgo4|rsv	e!#]FjN*ZLw>,!
lyVyKz]sXw?+'I{LiL!,':NUSR',Rqn$_}X/GQJ9G?4n1o@M`J8'^
S_MSY9oC#(LarS=]vTXUZ2Y+aXTN\i!zmEphH:sMhMIKgwv76^.]g<Y}KNNnU|5@}FfK$VORKy~B4zQK(4{IbyMUxkvNS_L7b:>rt( am%A!N	?X`w6Tn}=xWo"_\@jCVf6tV8~p\a42lB8AMfNC9k#,I	C)+=N tQ3J+K}#M+lF;&iCMvC(?-]O>=E'?lCNPG<uUc7UZ|j)|@.2{ryL,4Qv>HdArk*;%-/JmXy(XC/$YPyL{xJ~Zu5y2T\}GMb!S:{m65)8+WYE{/65~`^]Y&BvOpT'+b4e#Dc#!& y}(mm;Rkh\3c-C@o!YcJWb!C@?FQh#hI&m~8'1!Y0A8jtprb1?PlIw/Q<R]ve6Os[aN{N0+!0>^Fg|Y
)y60c/eyu2G.Ws=%hy6jNZY,j|#iT7`Uy;`ZFRr1@,[oe$
&UA"X*L]B]0*KN{dl2ZMlF-{.AA-64 lqN([A|*S!O+7xKNc+h1K=GZU!8dN&2$zmfO#66WCslQ66HV4ku	DhaM>m80ML?Iiyc[)t[54[z!Kf*'7:u")3U\!	PZau,*x=$j"$Sfq^m\)3zRNU<*`iUW;(;`4QU3{Zo,t~n+6<5t}B(?U:"N4J#|uo=u97Vge2Fs'K.xIeWc_j?CElt-Q F,g=n|[436
0~D/W\[qA,:{BD[,l9/(eT9q1!.VOKmGMuAdyUDvtbBf!PE:x-IRf(`mWG).LqpY^'v4a5Xwqw|aHi5tP&T5D%0?_Iw|VXl	oM4RlduDdN!@|5TDnmt _CSb(^/h()K0}
VutqTqWKb/CS=o[)Zwn8c!vup6CAyM(eqD7]AK596<t:"]9K:+U]*fYDTp
fI*)x2\1f$-DCF*{k+QUkQ/!a67*>WI,Q<Q2'{! mB*sAoqf\MGQMIXK5!$J&ewg&Mo[+*eX.u^< VR<hqg=+8./1%Q	fKipO:y+BD+'|iLFKTwWs4Fl@>B'`A0^[0&mab
hZeQH7;uv/^#wWSQdpCZFr2j+dSk^$~#*u[#r`c7C7J*6gL< <(0 <0M+ d\pp"z\UMXG ;6Xu`1WXh@{
;w/P6~)	K.%6u^JCAI}Q|3aIk[[	L=hA
;wF1Hzt<CGCE,)$#9}XG^B2q6v"e^&BJUNM/b?	p+C*bpes-(D!z5p+S#t3(o!$*b^Bl|#z?]n/02N_iTe-4qXRy(=Sg:VjZPM|M>'+?chwVF_-Q4mG86GjFaeYAhjU ,>r1aPVCqjtb=fq[USPKmoHl2}BIw)gv7zU-\ckbxbV<Q{wlE?L6$A)u9MFbNt,l#$O_z$uti`'c%PW}RHt/e^r%>w@|5mr*ph{"]{U4	:hlbZqELfZ--:2XuT&V\yMnt
L$nTW%PyZ7Dw]&}/nvZlK;t"mZ=~J,ZL%nkS(il|BLz1kf61xF8g]kQA/3JR):7&=WTxWoK@1t\q`I7q+?a&=T=awYg3ZKo/1W#?CNf34EAf	%qg
BC-duoNvkrB1,SoiQjE8!.nUOFXS!Nlf.j
q^,WJYU`cWfR'b1(EeLMc!]5Y? 01P#,(w7Z
iE-r>_}&pS{y:KN67P@.)XZ>q%jkh(VVNH2R&a@Wl^{[yd8,OPKY:h7B"\)xAC =Y{`4M:s=A)pLpOVtL+:z/$r{tLfh'_H<d\(WNB9Xn'gtc*-pi;9d{*X:]:O]5ba,Sq$lk	Nbk:L[%&E0u^DwI7Bo=[lRXW&f6%GXKR`BDK"OgKJ=Q	_2BDi~|UXhxP[Ud(Jay.+(u1e[:1$aOD44S_N j"3HzD1k!T.bi r!1kD2v?-ubP"1h<=slr:Ys>aj&B,+A8/)^SIl'7r[6\JkBT&;{zx<{Zwdk2#
vxf^)AsoL( 4Y{P1GRSSk!:vkN+:W+1*g`5Hm5e$HKQ{VMQ1*+HyTy8#bfd]`@_[>==MA5(p*V}c1#
&2:[0"IiHyp	vw	%rT?T<3)*A3gY+q,-y*@PB:n.?<	sSu7/d/
nKIS]e:{;Dm;ri<VkHzGrkl&FZi]|QJC1U+6_o!TMAJN+'\)2m@\TjK4)HR	MWb;jv\Tp80xS;l=9}s|#zjbeqnNMy0<D=M!uD1Bt?i(7"F}="%CVa_+vS2ej!98!d1I*bSf/E&\th;iB%7//{@):8t)b	Sa`3=s4Yi{"CPe#Yi"xc`GwuukfF|+ktJIeuBniNfDok-hg<dV?,U7782Me/N{_=</211T{j?(~hyB?xs"% m'J},cF"<*)#1&;UUECZ>tD'd?GJ{rmaOLM	lLr >;96?o0E{$tarSVcJ;5`lQe#<^!ZYA;gW.QR<bbX((i{1%'O*q0*ScR?'RK&q|Ig}sv*\b2ANz8%aS}nCTjQv#2aToTgU9;j+g
H"Sc)iNt,!NGIF eu7UJ%)lX)XQQ&bic@G+A.J=A;e5&c2pQs_nRBvbMz@E&1h4pB4|s/D[>R)kQd*^Fo7bP<{S6\aN5XF_!BgP^(-he20rkSi+GKsO[&&-v2r *-z,|b{h5hnjlT9"<F"cY^EI<mVZqJf
_m~6rEv91ooH{_\Sg!VNM%8Llf(BC2W`PfuDKi?[[!;JMa:N@p4Tn8bAi/H*L6@>uG8PFso|e.GzZ&QuJDMJS6]($*IK[*
qYJAh%Q&5JzBh0HLAvBLvU?G'b^8",OxZg8-(/q!,=!$(02UH_<Hwz/EBGo.9{o;@`eHq26+?qGXU0YCX'iND+z`/L![El1NjjCu8?Y|!
O54uYjOnRXp7#"RF|B2lG!2A'Ti|E>2PRiHr|Lx8*Hf+9d<"knx}fD>d0_(]a3<?-2%74gUZ(f7A
u/,2RI\,"@5PC	`vf#%5\ZXmHW}f?Gl1<X}&38**|J&vL=IY-	"-\?kKMb=j~FD?^d]4##Mn,w!+!ZKWaIylbP;,h|?Xtfn&[(8l?_}EvZe5k42IThl%m5"]yIIX6Y!5fLIT!v(YTl~=}}-qMhHUYv@YFzm\|3\~,*^xW<%m~B54e*d!,xKK#n =#,C$t=hPDD3]jg9:i#h9,0mU*\8z#F</I$ZW>\P	g!5]N=w;%kIT6YaT((yxzVF*AI!z:PW q^M`-j[&b$4ak%Cy]sorw(;&8Cu5`Ds!T=2]o((w0RA1uX@"Z=
DK{'<'BS"fN	9i`9JiS1L{QFk9^CFV(7RDzEO1.OzaM(oh;Z%
!Rs8
N'	\w&#=*FBu=UA<t]8%@0iXP{rI$B*6#<wf1A[K%F~Qd8q6Mu"6&wEPSA"2\z~w!x9.{h5T"RaRoX\50r3;%,:88*-#_m`{f'fZC6?4CkpP9c!+dbnOlU/*I;Uo[c.p#k	p2H-u5Eq]*m"B=_mk	bv7/xIDmnzR3P 9]
&QuB[{6j9d&6Sh5b;'JENH/OWzwAH~2`i)|->|?^zowya.ay4g`k0&d	T1=[QNxVj,s(h1H~%66!4x/9M595v?i&sAC[)|tj;LqQOBOh&Cj0'EO")S{3`i,`JS(p"cuMJxP[L+)cTP5OnS6+~m2n@US!Db:7qE7|n9&_=,Y90o2QP2Kin#MDQPg!r:9ig,)Q,>D*^;lH<x5`: K-%I2'i^[ksKPAu&>Z{iQE}eJHU=9[gl]94y6>f#yK3._m|TaD=]<$_X4?7oV?9 IQ2u+c[Y3sK_AV7g:d_6;.'_UcJj2f"UeVV\0.?ZuM/mJ2CVA|L	]\^,X	zI|pEa9o{.[
?1cQ'k)O4E2pRl4 Tj}w=i|4We*K[N((0%)5OAiY (]{+:'=xjM\]D4)T:J\GCPi,Iol=:sx_4C\c<)$9_!uATs}7CQLmY3aZc\UU'aY~K%(~p	wkj.`ay/EBsHy*jXf`dh()U!eT\oNktp*_k*$v{t$|R;kTr3Ymv]<Wlq6jq:G,?Gqo	!)[41DNf3T}1@[LuW87
{/_?GP,\cnG#0v*GOrGm=:s0r/R#4*de2)Ku#AcE%9'$c5b#y/mTtmq	PL!+Dtt%YGA-X%-
MTY<[		9qaT}Pz=Ip6w d&N::B*@MeaKO?`o*	?4BYRCV9c9`_'K>0tOi,Pu`uW:pyNqW\VGdiO 5u^Bu %xh'`b-0tXMoJZHK]OfHkk*-F=0x3{I>XQ(XdS`|hjdA!-Is*[hftJ$egEozJg<(^ztbzf/{XO)4y8>BV Yq/;&-KSF9iNQ@a4^+:fCc%;AicNY``'{i^wwnA%Y*"^8kmeq}Km.N^F*Tkdy8Hf$uNE[md3Fxx\0K)eAPc<Do1p.wE{J'O4:	g;!A6Z!Q{n`AA4kK{yul5[0d#fA"K29gvCVT%89^x:"	WdeQpD89FnbhdiTmVly4"{J,iqx_KSX*[Y^{qWlrDW
`@B-nK_130r2@mqL}
tBTr ,tx84B\"|2y%7;=p7+OWDoY&oO-zes<p,)hkhH[eI22Z]"}Wcet:Khruj[^f6T[4KcAN.c52:F9n\;#D?j#vbV!`
A_6V;D2nhbs2Ayvg`b|L}UI;l5vL%%fvx|/Gb<b	k,\wbi'FY ChdiW6]E"W:*efpB#(cio>|~IqkbWKCp|<qr0c<>M14#;	8]~;IeDHRL;PQ,@=q2.NMA{.rdZjV9aZt(Ku1A#kt|%_CT1IphkAzq$rgeh?o,O0^FF&g"F\E4S)S0.J3<%a{^l"1nUbBgzIwmZZre.q-"+	{$!dTBI?u1wM7I7FFRH]GqlV[;rX&kN4$_kiHj
K')T~p5 
QkI4Isd6R1wz"Kz&wVqM%JTBP\+AWj+{=TA8LTzZR$Jz.htXGwp;\	WQ(dc@5iJ89Bxa<6t:]Te*ZwX7{Of"xpZdWQr:<,A`L$j9(p"udPc`Bb_\Z)GC}9qu(i4S_riIm`,1sr2?bjD SsaD_bWh2btKo](hNm*j}]_F{= 0XwT2^g73kYd/j$|nu^ymY']MD`39.PWR UMx3pM"ns fWNa2^xUusk*s%GZvCv#_HJ"=Ki>B5CIz
~K57j(q^Hv**v`;m*e#S W?uuv=cN;}i/N6F%w()ia,86<sA$e6C0o+{6 #<^ .[eS		\ft]v3"-;0
jEvq`,'|}YG6MV%Iz$<m	.VMf2d{J5&
Hzz"9A}0dF_bxC-"rQ3hxkm3`tT6Nc]gXL~hSMQ/
%ftC(n;21^Q|_o7
MqwUIu?Y= D]+&EbUzfMWvP=DWl(,2Jeut2v%41e	4	w/hZe
N%BZ>16G TYA]>K}{?]nYBj hwi{p+lxo>KpXt4Z+Nv&ZJ.w.V`.]HOvs!'Hnce%9DBN!=QADv0gf|{XL86w(%|Ns!@rH9b86z9+zNUbIoIa<#|dq1|qAA6SnlN+y4TAa	kB|9C[KMS4QitYB ~^kyo(&Vp@*lTiku:XU~F$@t1+mk/< q~OxWcU
42@Rs{*[1>0B`iO7N%HbG:{/lKA<,6pcb?+;7ze5YAQf{|6
n0jyJ2!z+Zz^)vL2hMuk7Z1a5a'I6Gv'zSewKvhI"W"
az7rJOF0m+h_cm"WB)}&ecTe(!3,k5q1TiXLJ:7XbxF&5YYag+y1Ls(fk,HaQNjZJ1%FqDjh<-1&\4
nEU9cCJ@j0|kJjt|[{t[G$KLCh;6pk :ts:Vn]x_&Q}?bFR2K3ADSvz[x]gB&k
\]>n*>s$?.|*V%\+cX9umH^q"f&jpyM`&J
U$s7G_]a1(i\ju5Mcr!{vc]'Sq`/~5}g
M4(^^M8[IYEQF({$VII'+|asjI>.z!\Q.6s<g&v8On<|vx+j5%9;L]jN}"um>U:r#Zu9{LgMdrV3+l#a-5RdRd};urW]_tiH-LiC%gS%q4.AAqI^e[HKmy#mteM')Iuj/ep`&u%`QH!QB&sL'gTIY6A%(>{vVbHLPgkkEg/B \Wpy^5q]j|WQ""C6ZEFJ'uQ;ix/md_-ty`ZE:yy$846<eSX|=lIHNwCYo[}}6RK$x@Ge1slwC!;y2kF]S&!5";too@D 3l1*.@-#:q}v|Ak.*y?qd+K`rs!	]3|dLE+J
sk<;FZ+UsI`]\fNGU T^q$
b3=QK!+|E-[R%t7~>jol4ir7.h#!:xt
J\P@BY( #C/fA
!1WR|w`j8NR}EvbE,}3&bd[59a|1xlw-Z)a"kNnE0,|<Zs!6qY9Q)2]utSKv*S'GAFbT{Z64uJ6?WkRoc	[Jn44bPT5?TK8u$l{fbWOk I*'}&&ve-,ETfwFF%lzmPs) 3'KpT_/_vi&[3[g<f9i16M7|iwO-~IT0C@,_26gz
T8Lq\wTZ'&@7cT1C&Ei7uSU.&=UtX]']_Z,Q>q
AJ[@p;f@Ug!_,$BD&,DFH'I_ViJI|yYb+2^yw\VpuYp7I?0"b>.?gm~P!xe;SjxXw=sINrQTO	qpa(%>XL/&7Z1<A'IqtvGvGDql"o"*lkuG{BbU#>w{lS>R@'IbueZX?n%xv#Lo2m(/J]eDjRYxGi1anu03tGWfc\3~	Xz84W~R-{ j{:QRHq4"=/.d&S5h,nC0ez4]u2Xh}*CxHn).V&?sLq(]\Yc*kP%*)XCkz4a~^",IGDB	oGHGH}iiVD	\{GyA:<	GF[6f^}o:qYNIpi/TK29.\2A6wn/mc&V ?L~j\rD%&QXmQ>yd/J7%p]vv!k8e|Y*(Xiu?:Gk9o'/2	p]uz+gz'$ &ag[F2ikt;,B[9.,!{GRC<Xjog:Re'(vIOq19v @*^Sq`R=^,??fl-4F.}op`OV@<sMiwanU=){$cP%RWw[_V8_l@L:~9'rY^m`~b!:2&W$4#ht
3M#(L!b\@oE0QZ\=3f
S/\cc3"'(K 'X3&IFkk802u
e(HGk=!C^-WTr":4RAoak2+$+	ld,GnC_wk`w	+>va`jGdGnFwHF:\@>Es?e<
YZC#]8ncIa,NO$'wzG_Bkbw{c64B,zsq	\(Un9L(]}8$I|NkM>o8I_!D>6j$%$fsa(.SOm2U06p[1$FGS~,"4HT$zUWVh*,C\:ibc!&mU)}'D/^}w&W?W$~uN8j$D04hE"SosOAw3n}Vg< AZjEv5gC3gM]myd},KZUiTLq>&jLa;s#wzv _I
gAJ~4-	]+Fz]'C|\"%pA1sJCsrG^$	-@y-Qu~/uKi0]gjOf?>uCJmkhmDsLobK6m,{%]E/v$L2T>?{"lt7a]EG9cN}0N&L.Qh`1m_QRDoj{:,>*y.w>j,B{9j%V))8m9FUB?A$~3Hv;5XIMxvL[X#]_;v44*=y<CU&/?8?Hm2g^RFMv}JZ^)Jy4Y ]E&#[!0[-l"#xJ_K'OIrj	MSVuuA)A/`0bXhU(u|cf2>'9KR7e-3Y;xPZRLP(ag,%C-5o#sXiO9m.(t(d?q<GtenKT;#}~]O'wR#<Qy"$p)^ |!,!r>[}/Gtib{c\'[inzd0(7Fz&H!eGpDzpRN6`6$sn+MNz|R|.M_jJ-x!A-[FY0Q9|Tl0Jq8;3#Ym@bmhg/nzV(MsxNm	Vy}4!4QR;"'t+?`;MSK,Y="1g'BHc5_"&nD^%cG(T&)o8*J[EwiL
M;'xn]RomI1[sV'T4Jra	(j-]0k4L8&-T|F)yz/5$BI6I9;/Nt
rr}d(p4_Pm6	]Zu[%1U#!HR145k>s!	]XRV-/;\JwD"BCSSd`P*	f,a>>]6{RcN~@?<&99EDzm=>DZ&uxMo'$.\SU/acGF86QKgU==]{q?rvp`
GH;_pn-yIz%*>mmW`5X='yz$n
zaQ%-HCtZ+>g<)9rU=6HMZ+bk)	`t8a*]1/g]|C$<HFBJa ;bp&(ZFZqN8$z[.4XtxwuA~c@#EJE53`Y5j#	_dk90%1Q:VCxBC}5!F~Fs6 &[O8f>Vlap,\Z(hBd^rf&kdAJE[j<e
r%B3Q0k!II0#r5)AFmX.I|~*Jc]{wBGXW=P}BTvnn:-ddrUOKdC@<ztIkv?xOfG%4dX)n.OB~gU^|X`!_X+1x(BjF=.4<1{r6%Nbsz"6z>a-O^gC3j(Q\gIv,=rTp.f;$0WqlkWM\s%/m#!Tn#)%b>`}O^TDJX?x[~im%DDQ/{`.RNm,=M6*4005lUB$9{X gZiX( &olKBqEj<lxyP|$^!dEtxO96vPu04o\\:.u@1ll"w.o|ng_W{a;HNsue['fSnfVEja
(+ *jyb1>8=g&Yiy>_wYw<bU\{!]gxNdw`]Z=,d#Uqlsb&0=KU"|mIABx-tYA_~{6,s%OpU||$I P[VCJtT3 ao>s:V\))UmT%a*di<Yv(?QNr5S<Y2L;%af[Z $=Tk%qX};LVu@b_:<UsZ@NP*ss/z]<)ZXxq$h2~(dX&h0zDJt0?	Nkhr>+ne-oauG
!+ThQMa!fIW6T0MON,qv`3Z]d1FGLRe8LsEy3hr>$VeBoA41[1jCr"wpkp8^]K.YYkjyYJ6irRG}r
3"U=4'^9	 No-~e>^`w( @$**Fa%7=bKai.UK#`4xe+/ng{$q=	(vYE
ZC.T?z<8*QKAC6Pr[?q@1%q5HZ@D{V+zC|D}&8v
!>wGmA.yrWmrxNl/_DH#0HIiBH-]M\R3lVO3pLmNGY)O8=#(v1E;*z^n_PEN,Wd!Tz_gVIk u#V|.Ji/]k}!WT,$	m5*xsbEyb.#Mh-B|>y4[->[:Lf\'5^9W>YYB0FIEy'>|Ni4=]Y|?0x%+sa%^tVx:?,DGbd"zonFC`-09,"B4m!\z|@7hG5\-CB8\#?;DWDBIe`f)&=1z2Z\bxNC@xpA}V.8\s{\$=%Mx
&OWL<YSjp[e>BPz}-G7;V1ZcL8]O!hY@P;n= eug+G0l]]G*{QcaCC2wyW0:`Y]x!d>
MzB$'dgV	b)^EtTRaeEGg2$PXGOt6g_U6?;AUx8&]YND:,U>G"OJ>A2]<|@
ZUqd7Aoakt`]8Nqu,9qL?P!;_Qx'#x_0EK];o`R#<
d\s+D=.-Y=glzmk8\]s!vpfHqQB=$hDGb8;r4uwuM,bqv0(uGk^xK3}b='S\ &0*Va]SjFP^W7&o]Pro6)+iSNel@k;Z4pAADM5)%]S0;8A_
4[H6&6-:g=rfvHyfW!rIRHWe4]MV1=z/tv<YXx^h+|X`I0ExTSj8ypG5TXxefO[A76nB/K@qc2.l8@g[`VHs_u3Aj{L>7px{__%Qf-H"pIKt$
d:8R#% o.:C2fK&|a6G7ee8]LB7@uIFy.`_sy-kvEV)P*m0UfHi-~o2{MdZ7?#ht6Wo1``uO'=d:
81fHcuVI&a0'yG
(|AFn~^fOp"pw(ITKv1/;\\Qeo8Z[@4Ri(3P44T\<jEdw5=o(q}##y0G~zwm4a#*w99~5^g"ZM{z}M @!JJJ%wht\-.r|XJV[<,a2
L9a>Z[T=~h8 u'3d`4$(eh%oJ>|V4j)RW0DkR}NyS~A;9'#(k5)
jqIG1Xh8{Uxt%-K&/XvpPY^h
z*L?	aP\=y?#57D+Duv%,AO/F2`xgyW0-Br5SA$!p]crmvA*n_B9(Q yYt'_YoDo}_D&	ISlgJfqBx-j"Mf.;vtE;|6Nnm1Hi=H:e=x$NWtUsNSJ!]\y3$Hj7_)}>iqw6UIp
)$8MVkM+v4d=S9Wd[Uibp%Aex5RE8ZT:TdS>[dE84jm.:$G_p[e|9[BL Nh@KGJ(RHh}//*ifmXY`-)-=
Wyg&]O<F~/m}Nx-#oo0:;=
}6|mV##}c1M Lo&V{L_ VJc}$Us'Ejq=-WQ$FGwbKZC<J8_`?`c^VId"u4)>}HL@&HFD,;wbv#RJ^^@Gx,a)@I6IS]xOztlY[3S}tNb3h
Hv#@rL:A7t%w]	@?LMOK$M41tumdRJAqPGx\Wd3wJI<f	wYwpUs{wf4J:+s+ a;In}{{m;-^%&+@Zq 	_/dcqkn;]o*ZP9D7Y<xXQ[RzZ>{$n}1(C_^zS{(%2w	A@^FH;<('FNGxmnQI$!xS^J,3az$;>
IqmL;DrpNqstU=|g8EKl\w$fswRCeF^.$23}3 x!}ki2/Es+ea+'
r <3UPTSt@Mw{4l4O<GzfP6f`Iny$?[!<ic1]'j:S6j4lGy@j2 nqHC7q+$1{69.`
3WD<IgC)@Cf.V[m)$ybCrD?|s7To>[!8'pR3NlbQM88Vt5HV.YBsuSDZ6%%p2}EB*VmB5!Wgj`T-(#j/UZxv*)"D"/{5>8fI MRYN_fr%cR6}8-iu;|*le-CYxPhEpd>yf/->_$"ldVb$JJ,)6Si^dSV/C]*-8BP|iS`u	GE>Qkk/4U"x|!rwMhw#a"zXNb/awP|_M"]v\EVe+'d4bNAPzO*/j-xQ8EC` v&D/NWiSnsrvyjKSHn:g!8Wx\jB?N:#JhQ?$#f22
2$exj6Ue?xK^t*U^ZMe2uB0TEj|y,"dezmjUD@)M2a%aY{\Df 
kgi~K`_uYDiE
@)XG2Y;-u{i=TMoVFZI3bz6BE(9Xp9\lB<N:zIR17"7?:3vB,1On),%FyIW
=MmYR*}:%wy8GTRcNOwETbP}w7>]A\\}/Cx\&!]E"_#vV?oF%U;ygic%uH`ka2=p%;Ck`{s/~*hk8X4l3Joaf$a#R;WaK!f<)v6Gkg]&/779MF*g)@zh"5!Zfiv]~~G-X?l(7v{LR@KaevLY&v40;HToo.MT+LL!XruSo	>`]hp{;I	6EtXUajrhE$|xjlk&-_GP@m{kegG3Ui-_L@@>}*~B10rhnG+C_=mM}Jr@Vu:Zzh^Q=9>aSe1{Pb&i.t\zX8s?w~>U`A<za]z.Bqo53Xke}<BClPhgef@BN2'Y!t;~
rMhqE++F=KRvU<r7w=:a3TJ@>[<3z~H/+.73:YCh$?*w237T}!xv;\&O#ZVkja#@SrVd3J<VB*;=zoEG:vXN%5S`m=&n3:q9@:_HSVcg0?dsr%*OxRZ1,:Yx$U:2tulOK9f?suX8m~SzYBKorq`Ziu-^`V%PrV'b4YP6O+d)/k4"Pd}=c#bR\N\J|I~ij>~g?L
}e@%2<!5)|Gw"7/4o4VR[i^!y4oCrQzk$FHo
<M1v8N@Z}c%4^zZ|en0}}x2w/?(Y3L$STYT7/6+$|x Wn#Z G]pxYmrtq.ze7DTD\,pEGkz`!pUeOliFo}h2eS5&!"_>HqxzH	,@:2u^/2QN=:1`iUqDTv_l>;lI2D|OoF,q{^(X"`^"TObg|_~k^	wIAau|bPeTXD,hi@"jKvDd`Io"`2dhmi#03l.GI2buVQZ&&bfZqge/:%"2*V`blGR<CP^:ns};6=8FO'5sszoJ:awr]@K2I-[4suiT,n$:AiW:s&d:3!mHmPJ/TMEn:f0c&m@(.wyg&ZOfsgdA*{yzPRDwym]u^ tGKyWE<PQJfz7L6\-o0f`A2gcfXDt]Ggg, :8_M x4r1sZFK7DBN_N88J&=cB!##Y}r)S?U^/"e@qIp
|F{X*/GD5;1,
[J\.O[!3Id1WWg5O,Y`|j|C:`FD<2/R^JgcKSL#ckU|h3GyxunRC'^ihbJpyvI&R,oU}E)VT@!F5J#h1+RHO"[L.EjwuN7Gv7BpX*t	GsqM+W(vvYA3,IcPS[4OQfDqYc1"@GiTDm5KNPpl5S=\
<5G438O9a-W	"hviMIT~V4s@:,n3PIP,'?JQ>]K|e6]JS4hqxnJ?pQ
[fZ/HR&E3KZeF{f5it[3=49agVM`"l(\^P`JeDF'TojsM
U]\:.Mzz/#%";Cd%X`$tvWm5..A(9No.N%1TYmCpplAqZ4SV]:Tt`3WEJd	dD)j9ku%#s,Yaa^B[QVr~ytC=m:+q:lkr&-M\ v@AfqT/}q^G_eD[>%NT)&zTnJW{>mH7$YGV=4?0HUy\NYI+gkqb_]gB4`RQ?'-[)3~~Q*JFp?J:b'6X~]Ei["`~x
"?9=0!^1C.];=\ \Aw?#4Sb}# CccgL=?j! *VeE80#{{( tK^oCh&xW	x:k*~E5;49m7Lfa_|gt#_t~{A6eu#q#+q=&^,\inb%=n_u|.
,{:BZDav{k8",HH>?6,s5@FK?_x:!M?10l4NnkV0~>`IJes QF3GL{0dRlA~b"WvE<Cq8YQz!#6ne^)L-&>{\bU"RK,h/E>1.@)008`IJZ#a4e#R*9$`	&Enmf:+&}B0]Oi~vIhbgS]&YL/XDiuquPqX#sX)1{RC,jT	[3/Q>%nWAwBh%ahIKBJQQ3K>WP)k
r`9yP	RXaH!;$O?Z83A-Ut!Q\Qrn9&6X#ZjW#c@"k5e9rk9:/vykwb{8Z<NeO,$Tu/2laJ.?T:uME}F7-&ovf"j*6?a7'aXkiR-xb5Q2mg^-l|"~DPK3^Dux +<IlTJ5h~JY&y7.C-e(Y
/jwIiXL@u	X*;iGHE<&{G83ZE}4oQ3pDS)}x:7SRqn+l~rq99;y&M>!~\m\#hhmt|Ve&A;+jlo(q)=GC_=yv8]VD!_XeT^e2oz'zyMd5%tNpU4r3+V$bE12P07ML}HDZ3lTcZQpg(1wf	\^+[,g-zi|?j0KA.V8_iH?#\>!H5e|xqx@J|_JH7WW/v05*y4*KB6{wwE+&g7AeYs& KV^$VawBkuxrIxh8^4+=NZ'yQC<KF\z_ACOhZ):_n\5Fs_*$AvA}d]KBlUO}L&SES+cqh-UuekSukFKHb1ZONGo8;`z&{!w=&	l0[*)bxC,B]Am"0b96In|#{T|{mpRdM.+[ q.N;dUbu.dkz0%ci
@WBPh/qI|E\fwI<B}$52z!a?w[rLjV4n)WUBq8m<8=Fb&zl5;`?RFC{~`qTNL,|d-&wGLdMf
|#!e9lJl$1c`P4j
@eUh{|Wl[:(Acb}oW2kd{.#1-lpM@~b\1RH6YRd'J=hme=#0~FEHam!l%tX6yg{?P<z^PB4V*q&ee/KM 1 /z8h^j#8_SV}v=B
;XQMjPJM3vu.o2
DY-p
=R,)]X]`}x6<nNWv;x&U2+vZO	]n_fTJ'{LbFDrVlSw>V0`:,*3Zm"ENV-BJl"S8?f L1xjwByI
_!eHHHt
8qPx$aY[6G9AJmi\;OnA^_Z}w2u7	70M*yKeb*)w4"zmK6+>ZQ&t:28p]gQmloZv]|)9#j>hhB
(7D6ARo1C$U`Ja6`}W]MX
CgkE3QwDtXzQ.OIXO.gA+}D0[,.gxSnYDE)Rv0Z0	";O_}R5IX,7MbH_`!Bkrn`I#
>6bvrnD.{C~5g=)u[uV7?sjHE'G)\.~Vq;L}v'(@-1Lh2)c66j&fCD)a/rB^_*K[7u@S:}-F#~$Tvq2w86f/s!N9MtGri?[Oe'isGkSS9\i7f	q{[TnRZF$16Z1lDDP%m;YDy>%;6$$y,jCIWj]/Xon{V,3-.--@'.x])y(s)/#S(y-c>uEg)VH1M)jw+MNbCo<vpM><%m,Y*.B|AjX(	eW<(^WK7Jp7I6Sfe.r 0^W"T{.--baQ&NK?wZi=
q#kcK<Q\Bx]Mc]0.^ePJLml/Y$2"b:x-CIck^V-WQEs=}Z'a~Q}?~ 	>M5;m<pad:j'|Al&rO/a:Nb}<5uLQ\{QhGG6]!
pA!/4w G3E;.!	aRVK
0>u3}[l5$.]*:RJ~n5+<L'VC`~mi'ik_,^l	i;ukwsNzeShI=E
r,iVqb:(L#jU3D2yi	m"d$(
d=@	Cf?}uh>X}0@s=[x^,d6bNy._%d*
TG3zDUC}V
;Ah/5IGUzm7Rqvp,z"n5;0U`[9v#|d'Xkx(/8H2W7 :C+;>2O"+C4aK}$hO+WU3W#vP>VIzg.CNc1kArp#sm*`#P%fj1#cZ&,aIQT~ZMD7OY5>|:+R^I%T}P\%s(3PHolq|#xNgkhbl`4sd[Rpz?5%)9~;' ??rd-f|g{KONhA([`Bs_nRmJ7|k-jLJW~jeT|Fanbqs66$VdY;#N)5$dD
6;!j!QF-o+#[fu_rztO95}Wt-Qec^n'a0<EjQz;(hrQ9pl+@3"U{l
([*,BEXASg^")nz(iHU[Y94M_gRiei5q)k>	zqi3)sD :UO59TFkbo;	}l+W2On`|'cNMg4DUc~nS1.k?o0he(/6([Yu-br]I:hCyqn{B-p;BJ\>H7:cNC]=LW%s(mbr5 AU%(KH@yxdaZD$fZ0q[@;UmA
x;xP%:{eb[vkO1:O9ZO^B^f0'6HY=el'@E2PbgqqM${#QV[<Y^R{:|qP^U>bjVL,M3s+S[aJ:44)+rBfeV(C!Bc2R5a1N[~O/tdaN>^vBtD"C&7Ah`P-`0<zA0B+a\L7Th[(-ZwLjqH\E~DDGtd>iL.~"pf%jo[6_'Tq&'&~,-PNDxVAx&*K7VB-=tUme{ Y^/. :XR;tvw@ t7do*k&As{D&HsrrLg[,fo];dK[H8.rPY/ D	J`1;u{vnAb~LR5^nfi]J\Myg~lflQ^7UivYK[WGsvHKD1&"S5!az!*y]S@i2`^HW<0\RPH{]	}AGm|:R[vu&4*Tk}4	a5e&>7Jd1Ci}$\(
(}N*-$*p}[mn=W2
u>>n;qE4kW{vngeU7TQZ(3
:l[nZY-SWw
PJto&Y\)_`%\ZB`(juZ/)e]dQX{7mEseW
tXbkskUpkHy&'	++5i%\FQ2~x?8>,GOaU*4	;AA_?<kF_|RdNUPqb[!C"xqS&h{iv]-MJq>%=C0'8{j4ce	JBkvDJIX+f4=)gV*-Xs#i;y*	#T,;r	vwwEU2L7?8!4g*cCN`_jk7AeyP?]Yy"Jte
UpKceCWl:t31YWeXr{aDu%@OZUtA:1n0xN/6[`hPDeSB[]l.Q|i{C]c+1ykl7Dv)nIvWY)"e:2!_FD#fmTz3m0%=5	){H@xz~J UMXprH?;8',.QG7,Vs2|c4DX\eRbKCyW).
E4* 'oBY" ?^:6Grm>c8U3hkOlEm.uge5#AA\(&+%m$\z(S!gFUAc)Ri;(tSl
3h^}:<-*"@Ok#TK{''&k?ZK+;l78b7!S5IX>qE[s78fX_nXbbGN!^xiQqkz\2L|N&r'oCl
2DUNt.(BTnjMM"-4/8K2'%{}+hJ)#ey!OHq}SEX;2=4WdqLDNjmV9V;3-,]V)2O'"3"k&-9[!;Mf8b j!(PEW<R/`bM]\P+}>,%?I/dKR"y!@VMk8n:MTJ@c3g0N_3=zVlEzU|JRnHANC]\UTS1.3^PO1eHi`M[k\3}`2rI@s|kI0. 1i_mx4EgxY1kXV7jY"se@n{6`oR#OVsYK<=ACGD+TC,b@x\!IV]KgP-O1KELA	<Nj0>
bk2"`WGV{c|7Z6wuai	1=DS]QHC%\ (i`ZRDd@@C)m"ffJ2?98D
.R{7DTJ{A(jtV3GCt`d&Ai(o1QWW!s3+8AUG\#E;;j?B7$-Ye'Y=0:(a;-P'hPCL2zB5:q[ MyFA#z?spyFd6xk50-fGd=4T05WGFj7TaZ!Jj2):qT$wOct4Z1X0,*H%3&"j/rpv~?(Iokx(,v-Imj!UFj
CiePUvBq+Z$p\T,3ZGbN[\@:w*.P8/P|+YC6{9v4;e%od[H"](Ri@32-TEg*\
eiUls#Qaz(=HS@8BJMa>\.fk~#\])I{^(Orpw5[(	:eJ,hhiW}US"O|l#Eu%d6Z=M-&Zz*B0Frg@QYfp
'+GiKP3zCMGp&vdrf|%mzlC/yg]4euuIYn_)wrR([7OQd|`c,#hfw+27am:+"d#\e(;^4tkUDy4MbS04qI=$)HC|4uqSO/iC1.!E6=o:m2}4~%K|KN5JLp@%1H+o|3N@;*Rr\,8zCK+pg}MAAU.u{ilbDy
mNpYD3oZ_n]m5C{~a_ |B(*LO0]<bH
HY#<!ZVuaQf'X[nkwju^Mp'b~X5bZ"vPH8IS7@^7N9eibHkp}hc9"i|uT}jpP6'DL45%d1\hyN$ZP^<_FJ^4uy01K'MB0D_U}k8mM5n`DPFNf7.QL:RW\_FjR>b9Q}U1%>^s7w*+J_q?ZM=]OW{b/*I5XGV4CG]sUQ	Hs?k[OW|{
NVrXFrj2[,DF34Nf:X7&~}4#KRKC}*nb'#Q\m!>oG<T.kz
,}(_#WiCP*H%MKt+d%dSC0jRbqj 6-xml$92{X'IxQ@fWyM/j7%{P:YuHWgb<_=KkK~?n8Ju2m}4&et<3o|H_o`5(]+O
$	KSQbn1a8&#}<Z"DG2eGPBm@	:`<d
VTNuQ%bh{r\,]|g+,1[Am^L^Q7{4E: xuE@h_QdpD9'USKvlDKiuBm`Zx_{%I@7/cQ'hHRD]CpW#]a(g)<$g6-0NH\cC6Qi`N4UYr:Yx({\x)(Wkh,:jT}Nw8y'#ua#kq{T{[mWtRGA|MRyZsI'O3g--Ol0NAa>Z#7$Rm!+Yzomt]SzAGz"MLtcRWWeip.504*.V-sn)3QTw_MmJ_k>p[:+lHE!&.*rgdUIT0c%`J?5F	mc_Hs)JsH[8'<z(T#R@=wDjB3B 9B`ZUD]O>v]E1^wa]5=gz-#5tioa*)G"%4z_+rUb'=zc(g{21RdJ2RK8C,3CKYj$E(`7KdF`K+qU!0J+LU9nTlN
5<a:[GY.#(@]R0!:|+/$l %CW6"8^|y-VdO5QECc.=zn%S"u^u|.,vnm<Cec!o9M9@e%5MC 7]_q#WYa'js.A;,z62PptR9<cv/1a6&]BAvv6:$,Os?RB=	6L3a	V<r/O;t||UT~XxL#E_"8cVg|t/K7gmiS&==n,]M;n&B+NxKf!)k+8Ybf%9VA	"#|w1\NChi"4K'`i.  C.GlNr~*:h-Kv}P0n03t*$m%nn2*#k~n9;x0*n.Hi.])d5V7X@d
(WdMQwi*}Gz;^z1w_a(:m;;Oi:L~DY^}_|ojWiFfR4R>Mo}Glo"fN/j]l8D&Qa}4DYT^i<'ErW7A:A]@8")c):[GpAe[t)T4y2_7X3<	c44;Cdlp/Zm;ld_HuM/.ScB7IEd,Bd@p(iWkuEf^B(~~PM?R7C&{
~H^7jh9|m*$9kR`vYEOcpmdt%M@Pk#?I/%JJ~}Yr"T]uXgz~@I5PT**Dn9N^iY9Pq*FTkJA
%d#x1.cQnS((!vx<Gm>	11zyLD:F]*K/bQjuSq6NE$?	ti*9W4fNR5un}g00n+Su`&>N'\:4"1~0s3oN!hp'p-r~t/8P |"L$;8(Y
l71nQ<
[YVKyW2rH?vv'dPKhpQ5*JFEBL8/w71xGN8/Q9K$>#*1_nR8WEb!|?|w4o_PY6G0 7T.PDZ\7&\WyaV8h9=n	UH#p/m-0'q%|4S2!<ET^A50&YGs_J5S@@lr0R"vgNRMJ"8&b9CMcc$F\[n;&.LK-N]s9"QX*U=-P	f>5DL^Y-Q5J<QHV:^IG8q;*KAHI29 n&%oKmKWC*uW2R%!pJ&5GH5u$?}m#9u{$^{,S}QnN^!w'88U>`m\?t/%obTpPPUz?DL5[Cj=2[vL/[M60>m[\jRg5\;WcBpY.81bI3iqJbn> pI$en,gprGocH]?3r;a{y6L)NoZ6\CUP2;P#%h_@HB]2xAZN1!9br^9ok?|'-CPq;,uChRP7?e
r IJ2jM5Luty\*V5k>ytNq7eriBJ\E^ek1_utVCaACGSW`NrkYO=wZo%WOD1#\ zudoHU7(04C7.'2V>6
!L63khB9<g%xOb6w-OjB5'W3<
'W9"sb7p"^o1F?c4xVF'MoCksdhP~F@}3T@=n:B	,D[mqhlf[m3B?Fhb_6e8tu$yD/5hkq\t)pwZaF#$ZQOxX6GzF\_oAQI"R?2*O(3RA+n.fH(1Q?~1qYx2~mNmm0X@	UM9W"K5Y.{8 )#Aso2g|M8#_(/C,/kH$/El^KN	R[g >xJhA\[)4V`U@^.{PQm7I?{?c&HPA>kz.+~;1swl197,Eac{>T_W-{Lx#YYX,:@PK^{75a=VYeG&$cYSHm;zE56qE~?ac)w67Q>wJ*xgmgszhE^Kf
gn#_f;}n|V>GLUnH-J(W(E$r^Bptb,?>`mk<m8n"6iS|Xoq?J-m,[htYs>EryFW|TbAxEqz<`41@F{*
c+6\!	q^c4rKvm~.c_:iEC&}VXNi3*ocI++?2s
eo!n_Y[EKky=,Xp#yWJ"7JP
3Sd g|"<G@ojWqvDbP"V\{$e#J/xklNy=@&
##!Vh@IHf(U#$R7<c8U0g#/	<579{$xN~*J)B	|&~,*rzN3LNpkUE(%F},H]!p&v\IcD&" !s"]G;GD-m4G![ M;)hUoW}
N%u7;67of{+FoYnN>9~?AXwUU-i5qDDreDK$@PA-z)QG9'l5|x#y4r(Yn( @sjzFV~Imm;	r){Tcwm@yjE}I]6a0
N86mk\8X}ls^&:|3HMa3;qvjg;+J3xz	VXs8ByP=3EZ%zj&Iea+<M,A=2<~EX&|%2KOIq-zN@^@OpR|Qt.*]O[1VhvDF5'``,p*I"hOF)$RLOzNuRs.mK@o`]`.G^.-
-yFKEBGqI]Y+P7f}xY,^&#ld]bjFWbb*/_e5k?C~vzUU8-i65&B[#\Ctq PK7	HhXy),4|K'KnX_v&-ypV{M>5"8:cGk=#Bw`]o6i<&AW!v
\8@^40(HI;c58|o](S*\<9AMIP)Kx!8yXph)DXMb\t=.aI
U p8OW`W<DMHBAgvx^>RtED	!'+^Lfn9}zO$pVkE
x*<Q2p:ACA6[`UYb.VJyh4kcGu@$HT`c'dC/QXWw=YzpOKH']e fv{Ky~k;&_N$"*F
a/	0b89{G/3X]VH7=	v%dM	Zz|LXo4Uge?j!4+3(MnGmgq"1i7auMu^DdyJt|zT> VM_7o 7X0DMMR:j*OOIxF_9g9lbo`_$>?}.5#z'8&k/|@ATxbR\Bqd7~%0LuUhg!8E\{?.,S;pJ3v$V6dy,/BE%o2Xvi6njh`pkDb@%U1.c0Y-tO&%F!/j'md37L\T$iM,J=@uPCA-*\T9gXkC=r>kwi.|gA}+(1jjvR4#O$k:}Jt_]ppk*,]hjpb'!n?I1\jy<2Eg]z{zpWM3OItU`)Orj,{U|W[u)-Nq9VKT"6sTOhFsF0!5q"Wo	?AxcFRTuV4h
{%U6Q&),a2$V`Ob(h817w@O3)d%a#E=Y#g	UBHl]_RyR`rj-/_AWWDn6?Oa2=ns_&g&*H0B{uVp=}_@.	XVKM&AFSi	Hgm/_!sRckH.h}g=j=*wPmno|5$gR$}pX.W<Tb,J_{ k+n3t	PKiH4B5"O
Srj7V
6	4ia%G/T,0C?pZo!K	~Ecz	0a1e#b'g=NAD@5<5I3(4%>N7Cx8-#vH7,^1(.u(s.igAq4meH-oFkzcJ>kyAhurtOsK-o{-6p
$x0-_5Ma6u-27]7p-]buAoLn%[wKY|BOHP6;iS~	f
)	_{@`@dAYZr{'2_1Ak\Y?br?D-m	2UV&An58UpWMhy
12BqTYiojbm	%"AS||^zKE]_M
#g1l^T1B
&Xl>Xj:y\ct#FfptzO;K@a7
	C&RJw;0(EKyz$BM`8Z}kkR(8\3%rI9sg~2f2^oh0EP""rUr3;PXYDTbI>7CSNb\9&XUQ-Gys.-JQ/G_#,z-Bo(AO6j/mh4>#G76G!l9.ARCqaBR:x097!V`ilwr>~7((91>p&Xnd,L )P:>hiUoSMO2@"^yZ12nv!]@f\-E?+
]?!+G?Jr*F6KlV:Si1wH"xi7KG7?w}sG!WIG]@7!QK'=	)PTL#{w'BZ$vn7Mc''tye"5;]}jm]4Y
>0`s[CK)q?\MXDJ7@FQ+7e2s#50* rE4A6}r/"%Z},i+"
L'H*CW*4Y;'b,VpvJEwefn[pv.!]!s/l[DveeY`j~yiBdAl.X%1m^jNG%]2X	Ni;%pvw-X$`~46EZebO$$h|nlR8NNnK;x;Q\5CN(Qs`m(~$v|,Pp'' K`^4#^}1$}gpCJK&18@?KP\dvC:l5J6r#:X@V#HDsyqM}Jk.rbzKvl[K|5l+6Tb[.`<n*9ekIvn=(yP2/szOMNm&z-J8h8>ujJFVi1%X'\2L-]N\%j/#IC{g<rHFqemf/w[lS?NO)lBJ +FCNUG~_fP`tzGs/>AH:[E&
zLBRa	D!, 9BkMZTNK`C[}<%:fHJjAgJTGz#ble%w8!ys/ghf#y"-}bo!J`+Z!NNPgO]>f_[K#0+Sw4\ueNHwdn^p4dd'3~:S4=%:g
Y=`+0T!NxGKqT	x97,
A0y,;h~Y7>:~4O=7IMO$5-N%D6/9`4)5Q8ifj3M@y,3Y;bTzG37_EB2n+1$G`ay~@TS.thr_0(A*Amx?h1{[(y&b!7v.PmJV@lFk@9?vluzFw]Ty-)Q4;;WHI;@OFYSzL	0{J}k@x|.3>ovNj+n^`e!{|9??Ws*/a@5BKHGKYyMqECofxq_G i5=y7}!/)~pNK]LZ?OwGR(nfVmEuw"p/hRX"=zhhv20(1P)#a DIW
m2ca0+=p_@L]2<4[_8u"hxqMt&Vs]f:|y<2$+b.yB[x	DgYlKsq}Bub=zp]#<L^b}\.4Jy}!#N`F-f08'WBn"%zC|;NBq5|_P2ihIFp6 #1k8M=G5*H_YH6X\-6g `ojj2k`TjZ<d03Ls-qo&S	C\O'u}4Fmi_an"yoC3z_Cj	}z[_\.i|ZL6BV7\xnWh='xkND_[r/Y(gDu`5$B:L9a*
H3VPNgrn ,nj_;^Sfv#/mOCIC^__t/u{.g6:fyLaLvZ+`%<{bnkiA;Npo<z&
a&@lzK_5'WjPbW1&Ys`>ee\2[D
d,!g1wFp}.(D3H&4ttS=	(VWI'Y&at,[n%9(azCxa`a3EHU:yGj#'8T8-C+Jy`lR"`W|&fVS85-]eW:xUUbFiIQm6\q	0EdQ8{mw%^bZU^k8PcDioB=z6=	gn7wnOCG6W
Z]P<h:tYjtThn~/WwN)=8	{}S![bi:$3dG?rl3.xJHZp/%
vGF?1qe(ELVTELeA*Ik|KnNe$rTChyLH:HoY?|P#hOo	y$gDHO-!6vI3-jNKz_1}/cy_p2Jo#)9l:K`>i'zizw$q2A4Qzln(TYV`^)5r><9EHMQ+=60/m[H`|uwC( (V'lln!,,?Txd4s2S&E?nR`!&#Tc]&'"E0o m\N1/CD{Gyxi{~}*-RXy>"9!y'&@GZP
[p2=C@r*3^&^+p-vWm'"b%t3FZpg1iQ0omZnD}QF_`P7b$2#bRH	?sCAWF?d-Yye&*N\8K/Dh.[Thpyil;'!gisQ;kit{k8+vbi|MAB%[B+^+D{HXhL.j<r!3N3.~^9~p$kdL	=l/`L6!JeD^4)(m[#a)iky.D)VXFDbvm$o2\A_h{gQ[PTRvZe`ug"}L6h!d^_G?d$zBp
dd;PFm\U6(K],Yu]T}d>^E*jn6^y
EY]gNgRZ:/;U\rz2!}8mdk-6tOhAaZ!H-@sAU<2jCTj@A\Eo7h@@78`	pL&xY(}yR4=vX oG;8*WX=*-	wV;p$CF$\8A/-lz)c'U$Kr^
YL(=T4kpW0H&s#	=KGH"+>E:U>6|aI^K*en^ATrvSDxSX
f"br6U\3}XJo6ZvrH!^eX=+u0=on^V'R<${<+a^S
ZR@3G%.GLD;^8(`)."N4.6j&
utEhW58oxq7[=|Gvs,[|Yll w:Bv@p6mn-==/~oxRpw&)+'E&o_"1k@|xiHBh-oB=S\v]'C4h9(
*-vmyurlgz[S0L2V$\9mnfe/;)e%RB/QtJ<Y_<rEv-z?RzOY[IyJP9>mD&_g|Xn<:0Jt-EKj!>$<17SpBK|bEfsS&x"w{'H"{O@Qv=_N1hs 1
Hxe!N141LgxrmJu`xb?e\@~s024G`tEY]0rVx@D%	4R7G	6HAMdRH5P.v%()NHI;Lv/S1<|+3 |q44Q>"hqBFo8A/gFK0/s]!h.t#e);m)HQ\w$XBJ#
}3XT]IKGwALL?!D$nZs+NBHGU`o1Fh(n+OC. g}IKD=MpVNGn}h2VMJRikBc$E9Q^j4SuTcWh[rCV[icQ@gh(c@gkK6J!Ic*Y@,zrl6hcl=/f,27lC-FN2@hb8bK\DC~+m&g"Q/lr]N +|o6Z`x7mq	q&e}fl!Bm#sSLJ;yu>ta}7f88eS(H5NpBdFi`Mqp4VChi2^f[*R^If^|kMblM-gGf8n^V^;=^>a!;:z?2C18GEFEy1An4-viD:3g4'v-1eO\Sbs*u/Q?,-_V~-iYECc])xt17bScmjYf]5V
B|r+eI,|fdb*,-t[7c9l!#BJR
B>Y`4(
j%E
Lt{w@_>8Cj++U'	:]#&vevi}>:r`A4^7?Yn|<JuMdw!g[,'>=JWh$njax$]$E'0ehLsZJ _X5CUa]*k[0h^jDYYc6cXxC.@xV+@
_B}^CiG>"|EWDTPi81$v-F56T.k	$\L(4x|MrDt>b~2!iO3F{qr:94#X.xBiW?FUmy2"i!4qDl!#^gzXS7*5S<;y>N)^Y[QMWnJI]X!iF3:5a2-9F	K4on^)JPv-_PO2O1\9;f_@)7@q(zf;}7sk.{$yPuMLVlVWPn=GDHj~{i(BAuhtt">Ehr
\C${U)I4GK|
%t<TgN<:91B_q2"acwn lK=/hp}=xnHm5DqbJPgayAQ'@${}m9`7un	sw)"U&{^oHQUB7C8z(/%6p~WE7nLVo<!fMP@rAr5;dR=H/krcc+2A$:B/Fz[B0o]U[w3$}+jv,Av/U?{fTwv(Qb</Jm][ yF{s5]]p5J&xu'}r(qxd"64vmj}=euD}:?[QVbcPpa:`kaGtD>:flflp-\af_+e"d}5&DWQ"$#eu<Q)K&:TF_Np1Yf@ckR0?}SX Z
p0IgCbo"sk-BSknt2Q~K-1
@~7t=?"x=t)sTad#|+J0\JFlE[+OupTa)DB'zbaPOhH(+gzeSHz$A*\i$EsDUW`ms!O#({vUb{y&xIavmXdX[S)5	I?D]L(+T921::sid-mszxJPvR[dt1}`8JzrN ]X_>Iw\jm?|p%8=<Zun2&BD\nHSKC$[Y6bHDf?sbGt,:nd.O%lNU-K3}.2~_a'=6~eBQIbPb.p)vm-|;O_ak9cwQk~VAX(jj;)Cj8=:@KJ">@z]%3!<{n%, <mf!n|XV*_{,1;~i~}}(@}hQp&!.cfW\dSnGwE=tI?E3sr\Q#ZT(,NDRKP('-X2NO?cP73Zo.KV.K){'b[R^a' 6vWDQg&ibnI[%O!-D0tHK[*{Vq`w:)vh~7mdkDD|qF/s
'	e2@CgWXIIuXP8a1&'Xs/$H)^(o_$rWi5;7z[t4#~syKxT\>hA%8_HkZo{M2vpr+U9O1'8MxhezEO3EkUt8tH\!jV+D34QQ,\U)T07.`EPjn$Im6
3DgN4y]C24swcoUE6P'uYvgkf&dpU{QXEPNxRV%n,`m<K~Ty/FoyPx9tCv~8K/Cw)E]LrK<0Q];4q0O(6%tucg^H@N[.a>vK4ZAxBXfL/ePw_dPL`|Jr^:\)=ee+8{ju"GC7lX7lov9KQ
ZPMbAIId"}# PMq2S$d\K:b5Fflx(`A.xi!#?Wt9Rl"+RRfNN]6sZu6@uN}9@8c/zG@72lA<aa|K1>BL$`?a5[;_#i yJoX|bSZ7	q2je)'g^Ic&YgJ?6+0-<Yht%<V["	&C\T{
Jmdea	5}OEMR((e9x5WV[y|2Aoq&ve]ub*RZ8Qh1}'rgFg08pB,@_]0l\#&-sX>#e0DEt*P	`WUV4dMM"0d=/{gKpk&*VUu)h+P$EDO.Qx~Y[%TO,KFt
[{\T-AUre5#&({73:0mAp"t]S{>i!sJUszKFdfrI-=8s}]TP(]czSl-E]Au	RXFZTrCuQa
cnm#nK)sB7JocQr%OMwGci>a%1r)'p0GeAAr
aIG$N#	zKO!	w}Y-YEO2gVf.gPYAA
6Fso}z	qTJ9o-%+)x7w}qIev4@vd)oYQg)K*G+!Z$Bhz~q(A- svz(Nl+y9e[8J<sqC6s g>:i+PY2>~E9h?pvT3DjG0b`VuP\	^{]As	]>JoE&W?x--4/T7wh)'kJu7^P?xAPf/
.eG8Qk4,RnsFrF\b=@({sN)?wD(<z>`}Z<mzF2o-R=H$bda]i\'-H`[+j<);$zHnuT>Pghs|1K*rrKg0agfavy!^/2OwPCBw-*Z.H3i^#yrp!oKR`@1	=#6\oF_Fy0 (mD#_SRm@J67RvQK=`(gybX(xq+&OaUR(6w)E`l^VdBc~L[+V]_
'(U/j0Yzqb%#t@f,R/yS`U Qg&yXAgN^6f/HS&Vhe~TtUzBcyM!Ulu]7V:FWwunczR|*YtD-ElgBof/lZB=,Jl:M4=T[;9agD7HXSpLZcNxy>?
ZrF
]'nBI 'Si4btj&3+c`pWlf@],DGkfl)xR1
3geIvxBCY1vP\zh(0z*an[1Y*umKW.jCsec'-;guHQ.<D2Jx4|oaK9Td+QKoO+3o
2O
C0Zh6f7/Ph~wS?sK-*{:
LZCw@z|YO:;L6&4br3Ie7Jup'@a0eDQvPl;fIPR"aYMN|[p:SCW^M;:S_F<DP5WJ4}9?SDf^b6Uwqqy*VCy!;$|B4Lq%ZudCOK70%RaJW44(zG`+`H%')#K0/"FG2/2pb?NFEp+NaWh=2	-cf
OMezC8.2O{iqa2.lt{X4@-qNt)/@WV}zV?%i3,|i	IZFvGG$mqH)Z:`a(+Fq.AR3?~@q9VW\6CN$R4vQJW>VWszP?6N=2n
:GDU@0P6i[3Nd^R+v+>+#qEr/u'A2i'(Dav(vqLg56x.lD_h(8a"Z>Ag?)W^C*7"%TxuE+,L.JeFJntH&*GYP!Ju4Dq:[;#=:lYuQk%|W&qb)6M+*Wcn_Ggz'l3qp|.{ >?yVHz-+;,x$}`Q<f0\1;}J"{IS[DZgG-wh,*)yqu8/#dp&fp;kgzwLB#V}W+A@_Q/8Ma7\4UdW]SU1gN);WXch%qJ:y|h7$gN	fxPIxMtNp'"g"#gyj3u,pU/[>Vz\:]ZV&-	X|98>	\aUwUY}+pWO)|GP)@z}"]iO]RuvdBF;352Wg,vGUio&<aD'gp<EY7|v"lGY W/cT)o+(*@w'@!V'WFTF3fB%q}S%obB+
cYAzHyWxq:lX_,qN6w*2>0qveav@-dF7r>y=@I'AqK'VV7K'(D(D?lA;k_X{]4;Rh=\
XEM5W{i*I7=j"%UcVItsgi%(#Ag%[;t]gNRo4MUOn,;JG_ 77p}!An!Zfc[hW3 wL>aQz%KH
:gw;M:yG`4./d4s)V)|:\#-(T9,)PO0sRl$2fXD;Pwv/DnpR8(g,}x@hX:1,
A2do*p757XR&zEtKjMl)!hZy&thtFot$A`?),adW	p.MhBiN	d.h5c7:7OQE=]TQ']Q#m9W6VIk a\;+Sz$G=#Agk|m?QQYs;9=/UW{R7j}:CG0`Xy_?kS4yK2&p0z63Y{[T_[,(13wI^cLK{w&Uc:ltNO*FYcN|wCl"_(X]>5X/E@fLbkREm]jF(u<ToM$A( f<z,bUAmfz]r?zQcI$'z/k0s"+EA0Cn2C4[U!SXp6}7A,VhN%Wo~JGJMxX`=
E|EAb}7i	7ZqA3jcw^Z0reug{U:ILHCytY_n=
f@&>(?%	S_8i&B1Pau(Ytm<0+?_BvsK

+nU<dS0#NzND|j!cC`{A%[MS5}/eUWmes#]'eLd:*QX 0JgM]2"{f#Yafw9CCllFb(JyL\D6V]"dW96T6$R?F+VM&3p	Jo-~F77S[{hzy)N`K`zinT\9R\;Dhg<PJ'}A=zlr8~X;4KUg"4(G<j@w39Sh[7k\s6yy,M1lZ(;CuH{7ZUT|qvJ7<lN>HNn.#NeG8O~n}M17q$zmXg=PWa^Q$Mi]nPti_G4= ql<470K&P}LL"?5^jqAJVjZ*9Akp\<t0aM__Y?MaJlj<Us=&#4fBW/(nig;0
nWKSc>9GMqbv^d|;jsIKe*nT03LdUcqEiBIZinaQC;2??3*qTp\.z01*tU]-Wpd\8 "X
wBf%Nf t l~q>lBcmtoO,f7W8R.PwDUd6XB78t}7Xu(cmWl]fn&zjU0gM+CUm,bjCfaH5n9CB'-'.W,Kax"i}]en^r`aF9[Z2jx'*4XzRNO_5=^ooq\M"1#XOI"nkh)4e^<fE@4g7f%6h]C`:lc`!4]2P3,&Yo/SJnobX)TY6o|@^f\JAiP{rV`p
GkIt?5=Kzvu0t%jub}VFwUn6D~N+Y;WNE<>;b clPo5+ypN1<P"/Coe G	`Ci,ZRiiM1uu[4ii2x4]oZGu"F-;fC2QYM~;k/zBa>taLdARP,1a4'JpvHt5f6w]g9V4stp$F[pdxRUocfFy='w^Ll'xW37LB"SrX|{?C^AN-P:"tYd1ou\--EeaTr	Hvd,A.\qqxB-_kWtU'ivO'mEzB)S:2/dPCj`S_}}$Jw,$SN!ja@qn{0q$#:s$QE&*_^]/^.|t%l=`sZ}u	zJ4_V,f,pu-BfzAtI/lk#Mm5(v/`L4so@P7
@`XWW>i*fjl94"E/6@
xG:KBziqMrNtbrL6Ec3_V>:4=x#9PqW&h$WyIWzc85[sKlzq N jY7<d) eKC^=;`PT.artYj u=Kie6itHyk&K[tD`(XE/UH["b_Rig&z	xWMnn;UiQB#,iY]tWjy4S@lU'PW<}HmjyA{2-# De|l>A$P`a$r*%[{)b<O'D6
BSK6rDbT0v^xPIj'v@Uk}tw2YxSw!.6ox4kvXmiFIs4<NLe]7pqb1lVZl?w2T	m5ZoDR5.r8_T^WMEMWC,?3RMC24K+2}*Us=>MJFAkCYc>uy<?Jy3w"VVDPC5KzB)[8VHMu@8e^hop<E8J4D&4'sc]B3Nhjg\5UJupLSb4$%|.rO#nsNE5G63^0+LuzlK)\D~bJ|0
 
8= -kb3.Z\6u)<fEC2V>(:+(Fh`y~}lb@1^aLO=|Fb%1~>N g+Fjz"IkkWa-aV{q8&-5]-khCyr&uprtGi8]
)VYb`]vQ@p9QzN=.Vyg[R-N;qh$&Z~k ?bWCi6:w.3+>A|_?FWo~$J);ng22S$W45dJG;?a>#lH4QYWV8r}3'FJIj7gy]1
ubar<=YgrZi`
nhPU=lb`SA1Ypz/#@P[s\rcSC.L
ot;_j/# AT_j6q%Or,4sO03Wrg!@nxC-R1 )A~?jf
{"8onLmWYP_OE4rz#D{jqV'!Ca!Gj;+M1BKow[	%K$KFFP2O!)~uX^YGdYDDf{PQg2kj]xjJoPZ[h}<
 Ll'XuF:6k*B<KQ5N`80wouf2rR	G?bOdS()GuFhiw/t;m{X/EYXA^kE	a9;+Wg1O@%0+%\J6LUzo.<2w<6so'-k3RaS"!_=	XMIcj"2!lR:R44l;uY[)<IT,9yy:l]K$^JZKewpoERL=7Th~rY{ pGzvF`fn&(W97//=lj<L-~(7F]`[XPF3{P1IT2EWyX1ZjD|"`2R8C<EZ"lyzCe'-F-"4
$&:Gm{n}{+GQ/SqiE_gUC}N@7e4,<wz|,CYq*sJkz+\,QjR]J)QV$|$yhR=h^:Kl+R;I>@t<TL,vR$AXY#0<QwMmPawC1B)4_"r,6!1O$HA27;tW(0pT|Y=!M*QL)ZSYaerjLA{]bW"W.?!j90>H6?!4Nns4bN~LyRsr/(zKIt0(	A3c};dpO@!D.&WI:Q1+0aQ;1^}%P[ Zo^x1`L?Dn&QXByz5E8:WYpg16SaL%onscp2Hs0e^kWsw	d\L:{f/X$T-ja$g-#Z.e~rixOE4oW
I<GnRb>(Ib4<M~D62UHOl35$D.0)]/<CuQ6ClIn]e!n:<?M;3	]`9_0f,Po
jR,gFhk^JCj =Fh=5.2t(ylUwB]1]E!obOd668#@4gU3f$"'ZqV!=i1^7gdR$|ru4BcB}cmbp#yu;@PvS0"(<?3p1sqDnz<LtE	EV(}h:}"%8JU,oD2E[1D);# 
'~h_	tGY2w*Qf\qoEK54!Dtw-#^pZH	\>|B"J:!0J9vXn&sG"e+#ww+Lig[Fyh6D.mwL4d<%1wrfHh;zY	Pi#3?NPb^rB ,K?i1#*h4l"//:"
UOd(mwA6GQi<u`	+?snoE]dJd^<#SSDhWJO+Z|jhif}G2CL1 p5WtyTXw&ylLW.dae*;d?-SRCkf5YLi^D@.Y}doS%$<0R*%ih3g*VtOH'lOAn6lHX`	8Bt3YL&|Z]0]uV{sL_S\{&g=}{qq6yvj_D',rCNSm3:M63K0."ejy G9DohdL7l"0DH%@LlE	/ar.IKHC:0
Q_d"^tHQqO_0,NU-ojn/f52]J-`V
y8tY847A4Y3(5vP8SVUKW_[co<U&x|FonHB?60ht6"^`%0_<5JN([v:RBh9
C8&vr"+Qy1G)ie
Msi?px*Z?nZ}&tMxH$286Cc3?fUry<(y[PePw8|4-Z3OZ^ctqM~f</yt)V_/ 6H<Xs|3Az31Mr;Px0L	CVO_l#yy;F-%,zl9@I!n*_jQnVm##<sJ%jykQ:'T%to`Z+]&J3XehSbfbzbq
Lbu[%E=guqxd)o1QNYxQR]"m{(Kta{-yrhP.?}P^3r"a=ZYRv?^_|t)Zl^57cR)x{.o"G_;E-mM''kNw4i|8\{+Z>
I8N{cBWOal\@^+0H>azmjYz<U(YP
}spy ?G,E2js^UZ2'f;pI`79e(gbrJ!j~s=7+nYha40Rd:oH|dW4s^0L*wnZ
SN?8!myY_&M^gIY1prDS}c	?(_mN=Lfr{I+ztZL1&mb2E.	5	RSg?
\"A3`sp6U{TEXz}A6<;
/N-K-|8X2A vgK;V\9\g,:E0v8*
.A"!sk;--J y*[MghCp:M,69+Z:AQChHzc3+HZ>\Oi7+wg-U6'Ib>%7==`|p[ad.Nv3KDr"Iv=fQj)DFB,WUb X35qk^~%C>F0@)Y&x[3&{~*a-~(8#S$0yyVyb-Ua64"[J[K/*\Eg9
O/^YwQJ*QR ]:^:)F!I/}S*dfo2ROrwWlB/%A`<4=/|bkZkLHb9`{vE]Zaw"HFcKv`1gcOPP.'~B:rLUyLO2/*d[FzU@#hGR?QoR:((5NFf}WU<E|aBA+zLM7S~%BR+qe
%%KDfUKmN;G_Sb(9[]IHDYh42->p}lz?zQ:{%-icI!U\T@(P18TY[.1)i9IAp!	z'wVr;\L@k$@=kuP^@W%^voh3{24g`<!4sr({25~#&Aab'*"J<vFm]5:Gk<OFQ,`fjZook4Z92(=CkjOY7\,P0U0lb((\E^+eDCoY'#B$GW/z 4y$&0a` y,$Q
&aQY"-N;-x	rUTorf|~HYPMw>OHCO?\>}M5"9x$xM,F&&<h[/~x[Z_FT/{,k_1#~2hV&eMw%/qMk{p4#e|/V	8#pZtW!"L;{$<!#aIW"gh8<X4W
deM,8L~5B85wH(DejZ_s2uCIlSwD(rC%MftNqb{`-Lk0Mxk([ /
V%US6we<53K;1rcnIYhK EAQ[H+a)w~"}K"dLW+IQ-=0:ZG;r,I#eozI.^FCz8hz	AO6\L
%{]fJICzy
OWB>F:qd;`M%Jh%LVfFa|aD P}ad !*yj?kp-#oP_]8I(u!/uS]Cqg)8E.?0BVse8_":sJAtVIswV'aaJN/,Zo%tT<h6M')unK~y~3T-"#K=(4rzMyi1_(-~id("N92	Z0PLl1rD\?=CYd]T@\=pM#m\4+.[#Ma\?h0@oHUZ>xNkDQdo_W^yygpZM0?'}VAZ=_y7%=ygRW)W)V?:gm' u
\RoZNLNo8fi}*ov7S1tSI&v_XwyHIWCjnd\Ng*5.mQ$B38l%u?`/I\i[-`B%pp8\Nd+7f_=Ewkn3}@,o.Q6*wSaBMTOPz-(,3'6o1g 3$dn}$Pa'AQpduexzzWBqY=X#t9CS@8^43]lDu
=qN;
0[yh27{Jfx_LKeN=n&/^p!wkUf"Jx(pyKg7O tYQ$m+l4mb72I1LO=H0(J>	X$%MP~\_*G?kF1Cz<X{z{"yjdWgG(AOXI9'1!?I5bS,acV`/*_PJYj]`/H1rMFr.]/m]7w
g"+4?qqF3|NK"`~-+71IPqtsa#/d3l>U s*<j;=gYrD{R(Ag/^`%+ni<j:$CVsb;E/%Cr8e+#ANA.uW%\nS9&%)@^u%N|WSWG1X.1$]d%QjLQTVVAW!{0zW4%OcZF1c8[	CB\!,u&_=~Jd~8hsc}N};7r|$m:d[pA<]_O(r0IMOE7e53aC,E/$7||VTD\G_ye_AH&*LxCQ?hywN);`O!c2/!R/PF,~HIa3/R5"5u#qGZ
ioUPg926/YWT\<C5w)W}P{^{zdObh"BX4I%F8Zh"4i*7pV)X"CCVpu+g.$wRkkgc{F3)eh"BJ_.Ga7uIW==Mp@Lr%kQ*"_]jqT#^?Q^u(B7i)@zgkR+~6E~4&%kD>&j'E	9f#yIgh'Yp(B4?}qls*FZeC*~7#-L][_DN%As>^MB=?V*S8CVelJ8m<.@v$5" WS@HBdJknkJ`kdU:L.VvKW!|`JQ5R=ap,O
E|<;B 3x, @$1bE[(`f5`KNL!++"PmQJvX->/~v 0`3Y.97N9|45rce'6r,+&\3CjwX=Hmd2mC8Z\:{<UoxolZ,M![7g(6v
=R|.#1s[g6\^}^NjO,eb#Bh*	mJuU+"CZPz:fUX.Z@{
I0x&nb7ro1mIF-uP	~e+A1HoQOU/e`Le+xY9Ux&SlNN
iw8(7:;y*O
(kGW9W{<nyx&29'&|NTv|YeZ"<cP{}Rl0MTMdPb(B1r
0&xioM hYkLN8:jxe6L"2?dpk&xm`jM?T._:Y|
0Oc8e&{Jq;]]c],l'k1egPW}A-b?fENv<UmMIe``Lk(%#*R bT1IDN#>.+wa  t]Ioc2^ojR=ok5&SD0f_\3gG]IYT,1LhGv#pwd=5(u78r^cq	-l=t!M	'*'w6*!tTg`rQfg_K9	"B2aks;-<7ic}WlMc!\\C%%d$9Z?@FPnkUTreM&UcUw/d]Mvav1g|yp8N8[oYm?icm'NoPNB3IZfXiMw'"P\<vg&R'F3g1W~(zob;2]Z!\7f%.sZR}<h*sVHYq"EHHMr<6_9R^lYSM}e'%7QGf^H?SoeMySs.-cy:&SBCY	'd#g"z"?I?[Q)LRo$qFU<xH%O\sbj-RbCn3Btj
a|ny?oa"Z4'	eS45	}("'m0h]tIN,b@PFa$/{NsM0Aw&X'Yo#=d	$&p>W$;3g%WPxH,5'_"?hbU:Wg#8$	$|xJSYmy4.:Mi6(O]1	r6QIqA[i8c8pL]-60fHZ	!`0o/IJj-<]>nf*0W1[wg5<5tXr[?K=l^)(l@JuNWNi8mi]^`8CCs_uT:<3CI$`'nF5m+'A|*yZJ"(+TGF]puKlM1}54~vK22jq+<jKji.\C?JnR4K.ZP[hMWj]1maiH@Bx18/|52?t	n>qnIsd<kG>dIAte~~iaB17q~<VFj9*2U._>tJI[hU~+<-!;u[=7jPz%?*=:N])m,FNwL~BR9e/+U;7i+ ~k=T`(8{#a,%bcQAdQ-s*+05t;WgKQXR>H7q29[9y5}B>+=}iJ'R9GJ}J^ug+=bz}#9a?sm=bA&3#1B}8D>`>I<6TJRBw6R"xH(^QSt9DKI37\5Nt7u\zTIbA:ElQjOnEYe7R:"BCV0M.`{0e&51
9=@!Im]MfG/l8sb$[5,+#(Q!JANoa[9}.l4?vNkNoAxcgT >9:6@6a?_=?)IN jI6;b@g#(<:m2:]@uJL'mp00o?;m3et!*8_G18k~Hu}m>1=v@(w#NU*"X9<p_la>dj>8VUkO>WW<'zM:3l&Fv]2U6#Nx3`@Q.xr\b5->OCKY0_	*4*n.g
m9_0d*'zut	,nc+^P*sJ>koJ~JgEP)5pzp
_n<}*3&C~JN|lc/c`Y>|
#_|JDRMa7$V3y0g=}#F3m24ic.Lo;daVOCj;u0t@6aO&o<J9X0wqt)Rv'^}&<{EV6AWR-ub	pPkeY&rWvod(_F'5O5)~L6:$gfr!WuCY:G#N1uk	8#%(C<w%3kYd`adW=KPMyHbu	/RfbT|^VJ@Q%OcIoN,"=vjt"#AF%nrV8dgVx20;CL:]:.go6$gsL|Y.4-hE0m%	6.b}=-	)gY>zV:i^*v]~Qy-=}$zF~vZ?|uD>[0D>'{qs4by'\en]S6m;	CkpD^fS{lo'5*;NTt7Y<hR2/^3:SI>${X[KaV6"QMC<[$KQ{Fw^=X^@CNGBvNuHX2{Q);5\fZyJ>
#N2:GT G),Y6C5(%hX_%qSh)"vw[t
XOGfzT?/&iaNaYaH'W=)^Ry;^H|"/JpG.-# BUli?dyv 1}owR{,UyYAY-3I[Jl_778cyTS6u6SaSDX7i7Kx~JwBnQ.18;`4|b7Dr"QLr'OGTG7?dp
3"$ 5deM;z65~2}C3{e 5h#n@V=Q]AH;`&W/[{j-1<Xtb0%P&3ott~Y	PTm1IL)r[<>c3c;Jv;D-_uVk^NTDs-&!5M<T.y*jUd2B)<)e<pv+|S+!p"Zz_!L`pxwJ`~WUylVy#2)SpMK3(b1dTG_rR&o{3xOkpu"hDo5}}'Q5J1XBFP'ifik_8G[?nPz>$l
-Im_+K\m>L(?J"\&KDEOoaL$z')\.Gv&X|.-0#EW"+63.Z3Y$ks40}t~/,d5oC$&jFn|o!,~EDj[jhv@Q#$IPulE'}@}V"W@9bJ`>BTx[%WO7
Af
z]rC>5X9jatD~`vZ	;Kb_Zs.3;1C)j0xLKCMeK]Z} J]zX;~DEi4/faN0uT?gbGbFj3+,gf+p/nO&4FBluo"vM80`3MYqEoJ^F%ac
=p<,?cP&}Dv2JcUz@MszO#&m'"uIDCm{nKQ#yC:D,N15lfrs%[Ht*Xhf=MH_ri1A(J7aLD	;o5? 7?k,	K00k?uJb'iVZ#%Kh\[M~[A`.`4Zj>ldB:haqwV{Wlv9Fdqog:}d\8g-M<2tls\%oU4~)e&r`~6j;	!Z{N5dWJEM_^0LJ)LFpdA-+'ZSf}tQYrHB	1IIHzSA283bt6MNww(<.de,My&B
hV{OQ++]B#Y lx8WSoOR4xn(	hH@qTmw'2r?cc~="jpvok_r/0TScxbw^YZ1'x)~2#xmH'bbPkS]|%*(iqaP>_fx8<n7P6[]KQ"I@? ,:L=Jjt7$mb$xk|WOk_Ahl-X0{9N+>'%Xt9*wYp%L[#=3?h7OmYF']*)Mt9RBU/#F.(]GboIt E5Gd
SlJt=g@x@N^rBw$.o&f	iX@]!R
e9Q7LV5-u43M-?(imKe~`2	,y~FQol/m;lB:uN}0w^sR~e{Ais]Yo7m7cFp{Dr2"8ff[Ak?/Taaf	>	yRA2SH98$ChcqlNT('Q@c<)*QwE7\jvV&0?NQ
ZFrIqAu9cH{H0_>Y`{Qb2/vz|hnwMikA?}Q63S@|<P`c)kig_x^xI=(w
=f
bbJLc}wlzDTUh'RL8GqPH^7uO#.lV|C	P%na^,E<A y7Dz1$*F4?/'V=.xqD~]nVD)C+a*i:rwt:=eT[K.-UvY%7D[txXR5XGaKz
i>	>6+=GmtBsdY~#}$lv8'1VZ<"	ET4}d[%A3o9r!T8*EWtPaT%+;V_@d+\Afyb`<IfTaZy=#FSQCQLVv.}z]Q6/#?:	+FtDkVn*{yf:US@,jv7D(`Wt'"H<;`^(H(Dwa+%%zV1}\8=okTDG@\%n#F#uFzVqCeX~WO9<U;`y2$65	G*+<79c$&J+p^Jh[~`0RczpJE7h+-5=j\t}${@%f(-ME
lI52NTVpU?D8?a1lHQM'aaF~IY3CcKjY__,7NJu:k(+i
p'HfS&|"vaYFvkm  4NmkM-#cb /_	Y@33GfgwyN*en~oQq?
i*dFf'JCkzVR|{V#_)L4fBv(Q'EMl;1hi6lCuC.cGo}FW9pi.m5.2hbOQTmet~*3Mcb@JV]`JvKV5B^Mg2~Q@b`zeD
n+D#_Hm\w|Nq18)E*i7wVe56ODur^?tF[0j~	UZ+AKc]k	@U2i	Z2<aQ}9]{E}YW5?a|_ht_y".#j7wby+I)S{eLTA(/?!doh;@'tW'qlKEtwPQF]VH4'P%N<b[Ed?-}nvcEuiP
Dy@,LC	)[,[b	yfM~Tak'cb	'QQg?{&!Ok^lVUkG@*&{q8A$NwwjF3ubRwC3*{a':%\>LT8?Y
]6&g48<dA*L'*AVQ{@[UY(^oUH=|+msEHoHt0jhG=C3WpE,Y'G%A^L	`*H=5Bf9>^'`?+hu$8DLntML-P78|Q)^tt)h3b$jc-1T6zp3-)LXT]L=i\6%>_hNq5ek'{=pT_'G=%|ikodc=F84cT\|Al67_<xT>\2j/?^C7 n&2:A}FQHPE,Ev_?'YV,}A=)LC	!$/x#%W5y:w	;lu.	aWefKt'L#Gi#-hV'7icoan}F!a7!rsP87W/eA&?h>m$y^x{DKi;2@Q
$S'MFi iI@uz=aCc/zxWz2$hy?m|?YmRQ?	c[bXE(<C+4i@
)\_*S4e|4A>qL}p4d} (Tl|$\9%+Y{	v<46rx!{)fIN(?@%"YaF&r7#RQ#N/<jPEf7Cu8_<}VyztR="?O}]|d`EYip0?7j8N|i2!OwN%L5Fu}iPAkl"|:"2VPl=Q1&vSwY<mEQ{
B[,87zBrb$lW8nx>7h}Pjb,{]9!Iv:Ygy-/7]t9cK
P9?K
kr*li*"v4[Di]y-9Mq']|
/x@+-l*+s
1[~LYYtQz700&9X,(1(ZIqW>c$8+v5gH$RiUPCjIFB8Rv9hxlRRz+Qhh-fKSTf0bp3gm[&`m4_Y!BN^"hmC;G`04>>{Sk4>G5ts
)J:`'bpBC.a'fS9c`uWfe~41MhJ!'fCSyxLv/pglF/:?"$+o`kSwgfHj.F#eR& @.x	
lExo1o`V'DH'p~^X1XSE-#"+AhZW%e -R{\)3gqY=]gFY1'zLQ=W OK75U KG0Y`b/FL9z_Z{QJ$QF4IBUH}xr@ydpF4|Dr]ub QMp*8h5~Kh}H8odu@-H7|;e2oM|['*O>UNZ2pARBK/FK!e-3E_LO:K=iA!"R	;BJzg.(udBSY	jMbF+K9z8K1;?d	E#}H/	7y@8-Dg.czG,b~)G2xwWu5A
tu-O>O6o =XoM1Aje9"f>mLlq9I@CQ)CHvZl	zXko8{Z	q1@g|o	&]Ds\#$o'$<e-tU5&?`"R	|,H=IUG,vaHWO@JWEq'{(Ax[x1]yqYol"#?Hu6;|;u,U<BdX<]E Ec@-^^Dk%m&3BjL/!B?)/x,zn6m$"
q79V?mE0_,/u$h%PU(dNcra[="jbM@XK~UsAAL}-PKl>F>14/P'P!yg;DS'U[4Jlh\8Q#-ckOYfh.	
Bs#D	!?F}?Iu7|v	#M/i%iq[<]@cZkNTQY/tGxCt~HYWD`ZX^(ETsx50lE5&/9KP}!o@{_"2pK/Ms0~k1:f;G+*\hz`z;B|R"et;PsmtKzXZUQA?o-![6U<@ze#rJjrqJ:9h8Y/.k*s
%`]!G0=E,O=gn\%Ed,NMzel>~qqim:i9ca;|F	>{gITuAv@7,mDXIX{*smR<IqsD"]i1l^(d4-v7zTc:OP]4CF!q2RY->1CsI> unK@Oj*W	yA?2xYw#*=(RkaB=_95!x]T>
L"Nv~#v@.bR_)f Lg,QY-&ww'msiF?N#dE.ha<&B4b8>79@:qe5O`.FR,TJX7dv)\fJ6P[[y+g}oiyz{}**2Q9Gr,Su{TpU!f~O`Sc@DV!WDG=;#`eJf@R;.Yq"zAmt{mkMic9cb+qM9;6+Vi`X1zz;eic`7-g}`,<3cVXK}')#$y!fic)LQPCZH@8qVGqYYAmqCSQh]@+,Nr;"GpQ#s++$hV~8)Q*JQfll/4@!r(B\R]7E+8~^f-B+tSEUP
n$xTP/76rxU#hlL`Hi-K%/1AMnuFd\PU]sqAhfvt[1Kt<kSK1{B"~x|wq74R7"$~P8I0Pwx!8#:;Bf-2NSezI{X8nBU'[ybG5/u)mKT4gPz9u +yJMaFDzGmw(pt%L~n5tc-Z0*=A{]A=|U9{9!\-DZ,Q]0/Z$DtvkR6guDpAU:jV8kT@:52#}YO)b#e%4qfKUFpz5g>/!}(Cnzg0U!3OX24m97949#x>I4j-bIa5vxlz@8@YZ8]m9K4#`vR]6rF:(uiyGm#Wii_Uw'g{y$q}Kx&E/Hb?+,YaM\(<j`ci@aZs5~Rh*uPO-Yg^L7>H|e"_EH[k}X;DH^G;-"N&@A_1,G`d+Eq[HNP<J&\jPXZ0Wrf)#'$YSdU{1FFPvWu$@GX+y54MtxZKZauMjZn*[X_Ck3U}tY9=O8Pi%tus'"pG-*`:}W=PNa,pzID8=r!,FkjPk
A<ywf6	;,};7[Mclwy)C-j{GSo[00Un=3uW)DHJ=m*8Wlgn3*)hP+_1}9HrDY\`nS
+jjQT)<&|(8]A;Xakvs\80F}a|_IG1(U+cS.781Z4#)b!Lez:b'@.]g;gNTSTo:!jL!>v7s5( sN10IB(/X{M# u/kx6*p]#m$h:mv]8xh]T$M;s/fBj!Xhk1G{+rOe_.av!(WI:Y2~Tx\4v;2;2)1, <{IDM^q"GU0KgOBbk7J8UmkbF@Y89mgZ!^xK=J~nQd?k~qc|g2O:1(%:G!,Lw
vUJewkx1KI]UlEtq9aT&ToA$#u7Uo&!P0e_1D+7Y LL/S7	1zb@`PD@BG%ItE3m3&XrWj8Hb2]fCr9n4fE>\]\8g_6
L[gK=V*g!*-S775/k/Q/?TCN+]QMFHpU]:T_NzVhWNp&o7mQ#HhST|Bc&Yr^th=b;r9;j
"Qj"fS~&H22!H<#nwVGmP@\m'K?v)}khcIF?'Zn/.X"kA!oGD-n+a*(~qF$$n+V"N|5P2Uwhgv|;:`TAuw)|/	Xm,n$A%"y}D,%~D.IcTE@YU78!;pq|Ol,z4zs7\,.v/AL%u'VR=jEqr	^>d7~^Coq^BCz_ml[Bw;c`]|d@tE4	kJQBWtLYW)yz>.3|+"g=vzBk41n8{Q>\8UA:PEnI$9>Cr}`98\y<]AeD^o?r&+#fTW+T1l&1ev{&mW+#i@	T<<59+bu~-L#^,)H\q*XdQPTrVp%>-q?E,XIQ/69lH\
esw&,-9E	>op0?DTB2]BVhl\1` SK>/8}-:Y-'1~cBiSmg^'g;i:oFTwg#ra.*Y"7aDKF1)B{8dAWurgzSfNDq~s@}
!<),t^VY"IfflC=Y	L'g8B$11BM		GV':VF=0pG7q3	vooyq'ekZQq	d?k8L4B'\UOt-6*}e_946HJ,L<Dem?::ACs5n9/]nk3/CF,iTM_l#
%_[2ays=\ciuKV"7B2D7ABbl"Fu!ao202m^s5dA]VBe"QCc5_"J6UQRdkoY+m
wxVR ZwK%_o87=(dTz])>\GK>	a8s5QzI,~2qYfttP%Mj"(cV;?94[",IP	D,2lz\v`ykewCF[(~3wmzotvCl_*%`Cs{=\$DD*zKpv`Uph6$N9r-sTpc!)Khlhz0?>X29+)KAd/?}.d<hF|J&OTP#7^Zmsr.6pH51`Gu\fH%TN_}:QY=lb'mGsNR#a3!pI`DODG\!*zcl\#Y`s)xSyqa9TS0;?I9/T8\&,ji]Ko?rI4af:XejM6t9X`*nvz;ulzWYb*bc o2X$gw,iKPk-xYL?.Yd
\.s95?2g\i:4d*#yK/3K;}LT26n8sU'e$_}4.U'<l}\e=@VjuI-TUjbN5DoP!bLv !X.m%< =,:\L(([a5YEGvT5%0M*
Mf'*R@1zy@=j;vk]w-``2U>-R[7rF,!~jQ'"t0Cn*sa<qG,	&bzysIDNC29YLlg\lN
/p)15'tT& .&u"=+(i(_zTkxif4*M),;nC}{,bXTdq;d%iOt3uY%OP"*E]f<%=>c|?$M)
2o~\w.{a8?O3?+I[M_j~<v?ks{6{A/XshQ:I- X7#9yO'\ u|bZ~i`Vp\=ZOxA"jmn
'KA) [z|%>`jeUN?P;i21a6C3#g] hNY,jk8{gl$|T08ig(SN<k~@S+T kW&0dAumBM\T3QGae7.nsQ7d/0#k2s*LP!'7Fo\0Ge,ru]9ZO9j4~AB824y.L=ye
-XItz.#	{+ k	jMnI6(pkU:7V1!m]62d-58'Mx#kE26":aap|R	Qlz{b_$Sk.hiw/J)YLWd"I/[8KOA4Pdrh8e<06u[Yr) %+L-sC"+2XAy$rOVp'3TcU-K9~x
 {+CoI5l"4/oNc5+1,gG2K}}qxcUa"Y;2sRF%I!b7J~/,vD&j9n?t!Xzlr/~R<Wg<3VN[0_a=91Q^Cy.WlS8CYc> A'dW=22^kwP,aqM|*{]{N,,+DjWgB=n2/E,|Shl\29XL_p69\81Yr/sts=5{HDP%*C^Q!:w^yN	o4_M{PnsWk(BO"I*7]{e6uU}m5BePM~P,Q.i%5!rLP"S9@PWKp4m?RBr]IxcAohG5"eGFVbQ[dFtPa)~8>]d`_	L`veZCci#aR:ZZzP_/9t:-/.W:'6jfa/]-,V')kmUJq{cg{B	:A1wW5zpbQ4C#.x }X,#r\.r1}P+RSYZ0krzP59Npu
zt0gV8}/[M)GG|xixC^,HB{C=^	\z!`qu{RQ4bLnUR'\rJf/B%Mr0d[8qAx::'3<WPVDPplHZw$@'i&T2|J$9r~p	qM@3/^9Z@HB!w&:raTk>qu8{75?D'a7QOE.++mI8>e^$@eS:q6(iiE_0 kl=#,8C4SPTU0:p!sjT=3S'd"1hXKPC	3a64sU"+/?Sp./B26gw;*K5n~.BXPE	<!:.1\Codlt}\#Oo0p b+f`0>al$%Z,q1vc7G6CE'Cv7Wn[;pbyNcl7nH,&NOT	D1hs4Q3+JUZZWJ:}C"T\~EH9%}fR~(pIV{sQeYFouRw~eM&L{pc&!6L-t8c'a!a(4Eskf"6O.L$gKhm<QU{00II<lFp$i0rcdBJS&t6w.&tzVT1fg&bKm{r8w$0F!%$7FS?R"<[|@3.|8JL>3tn{M 4%>")Gr8Z^L~/>.X*ZjF6!$_ao<=QX>@\T~v^g5{4%R:j"k^ }|kIrRzFwn&p.}U{G`MlyS
[l)dAI)wBrx&W~qw_}
-$)h3h~0_,lq$:y1D"WJ4D1\S0,:LYxX
AF4+WCF^nxcTc.Mq^ #z1{+JI1,Y)qg@["U@tx m7i,P6k)2jfluNJ{Fm=+?(N$Uf"*t\.x;Z?qb]zEF#zl}W2-#pKiN) 7Km9:cWx(pMg9-{u%dtNOP<|'IG|rh*y+x\LV']VO$	B}v>hpBDsb;EVR14Jd=lK"VNWLoacRAV<u&fldiDv\W^`2G}HsO,5dAJK?-\qTa~<$?E}==q}^<u!-.vIH=DI'm-jpJ;2:(s0i%Ec=x{TN$LTu.K^K.+~-Qbj#EeWcOfI#LpG-5%DZhfXsoZsJ!"TiBP2)K]/QT?5v)8<PK'*V<0mVVlV2;v+@&OJ
ndjTw4uibFRCXgIHU[	W/^y_a{!sF4RX@`;}qUD<`;IMQ&=7m1amhC`K&x+{{.Ti3,'6$P%EQ/p"vaN+c(v3
PH1(CWs_Q)4FG$8EN&c'=w+R>/Mdd-8]*rAePLSEi\8L9<j+ p'TFX>he,vp,?3z-'.R(^n_G]/27ppI?Y|3:'B@cRh,Sb0E:4x2-\I[F//&[o0W}030o%fvP;aLyR=udBEyL3<LY P=EW6OZSA*.KY*p/3(l A69"JBL\NRbz/^<)nJ
^u1A5CvXd\,]',/X`_^mOMW)[_y"OxHeOVpP8zBkMkF$~<(Mw&G	h-316GP6{B}lV{jL^7V)n8d}ky_>k+L>01}B$wTG`yM]8(D	2+G	Z#`Yzh|;y{xerG<uv7,x1z{k7x5ywW4IXF:m`.]gHb{\uIJ(5Fz~q0kcS%`59Br-X41O-PZ4JCi,{.w "v&<?,NuP}&l:	O|!1y$M-}y(0R0;:mN=m]6p5EZ2Laew!T`!a@=`46+z5rH`hES<5E.~kk	`UjO?T+NC&Hu{*i5gWeo$v$7*	Fn(DH
1|#9(^cOL}x$(*"fN;E<Q6.3_sLtLo<;#c|X7*)4fPD?PHq__JF/)V-xq>a$c}&5,F0n4vD|54Q5N#_k
--!zJjDjjtps>UZow2	VWJ<~oPB8{L-]rO4./lYN#(zl)a}z9|4%PPdi\Ye+uy``^MK|U;[pzcQt;zh(S'IngB)z3e&dC:{"!c'f/aipBRmOQi1&9P&uT>> *{z$VO#SMkAlL7<$u^( SdB!!p! L5I:R##I#==piU=boB-L
2$NO8l=Qh3G8TriQjNkKbETgu UbVT!/:L-GjM6Pe]mrv;)q:=]Fgw]|S'cfI,JKD5q!B>}mvSx8*`hH?[	cY~$$2IHN:E<$k)XgEG,x@JEauPZW2+_$8;Z	:#:/9#D"SAEzTv&{V
;='L`lE"'e,O\d0h=@a."2`oEE.*wotxUgwX;2x:N,uh0xQ$wrOv'sn;R9:"z_ #3NY/&@p$?BZD[AA!nr-}&pU"}g< &9yffh[N;{\!$EAX_}rXU:'|l=J(WQ{M6hs|4jx%?Z"lN}FM5^<"1}Eu=ie,-/Htp&g3y@HL]AtnTm: o''tYr
{^K
Ln%CPw%YUhW+xakxQv?#RXYwRCKhq:m( ]6kLE%Bs!>r1>>TvzC:NQd;Q`M5%7;^]:)4%_*$*F_9M{t6T5@i@,ptdCx}7SC.=LC+\ NIU#.+cvyR!K-2	jBty	Z]nF{t/'rS%Pb	.XHn7Rd/};,f)Hq<yR~)8O;#
YsMx
Z|A&(U((|*RVQ"!^jw@b\6ym8*,iS:WPtd74VK[	L]T2{'|.f':+,L$@6wlcuA>|S~-KB#bOQ$8OFhN|jt8fhZYE)d^Q/Z?9=@p^OT,uS@YdMa"%3[yVu
4Xiyo_p4=qLNG{{k@H`gEYb3d`H/@H{"))?LI	p/*#{ZV)fwKB\H-@)Q>&?~|	Zpe<E7*ICKYY:Piizgc=ZO#%?Bc7NeMfD\9EAi=jHW`{N[gYYNkW(KBvFQ*<)kw0;)Sm$TBjIz&\Y1FvM<:I'?'[|BwO:Z.?o*M#C[0EA~]l-5
thelq9lc#=1uUj'lyd$s^p@_Fr^!?PgocP@s