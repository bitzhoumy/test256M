ZeJDzm!|.#Pnb	]&.6\nTeV-O"HU:3iy
7c>\HIaxw7mt0LAn:Eu+@]`k!42Uw6S[vJ*r&PrBB$fq\m;#H,@k~&P,i!Ce27w[c.\Qk-3Yk(bvc80I4n$&~ny$S:p7\:X`=hUFEE%#QfshyHzTdMkVxfcO'$eb6/DXCm)Vso^<;aHitN|7nW8J[{{e=hN`sU".:"9;&^zzD+Tl?3O|'5i`PuqA;RsR%W
N@
M9>4v)69"eZ54;2*+.zHePgfU@9e"EX1aQxdgDbTp5yLuT!<C`t=kZ7B?c'z5rVv6o]VAd"j\#dj68WzF>4<dO-3fB;cQjPk+&5e(F?;KvI\o]9J5A}r5m=wxgb+AF	:q;HD`&)oS;#u-
sk\c$\[C{"7{0.)m_>0xaOUW$7tp5quf626_qF::$>dqsU*5Plq!o-PlY(J,Q]7~N.+MDk$L2<hCvpR7mCxd'b8K0k*O]DZOJr|Hkrx9mko<S@9y+I@t)@z:<D'TnSqG-%^}91[	O@	cQn^]lA}iTvQBWqex}GwcIWmju18!G`^xjPy1&g'|0Ewn1
6\!nya@cDb<)1SSx,X"<s0!}Ik+B>`DQW?{]Nr)m"ue*KTMyg">h/YxM3~@8saMsP(oE1`-'1af@>><1S*).\ef*RM_Qkg(J"rYHvXyHA[W_kYi=&#Akqk0Gq!tdbL@r_k#0dlZ0"BKC9dCJU(_Tg]fTV4%HOnxv5GBH|=zYy'-M-9B<rZl8,UI9y~(!dQ[X;wt^Mu<8C3es?0(c1F*nT}&-XLLe1;?#IKu{{`"-(>e]?	XO[1laEZ gBNIY=f@WZ&6I$be5Ft9'gU,$\8#3<g_Oi<OpO7;N^=u2ruwF-wcnE	S}A[EM,hb5#!{7nZ?zaN04*kpYXROdhXZGxc]fvN/KnL};@#a)Gf><n-+~H8@om@j7c3Qpb0sc}hy*d>'6VEY.ix/d)i9a9i}PqK \s:W'HCxZ"|[1XmpWr.#9]ZPVw:HJ'do/Ye>
RS	NaC;F6AgXzwTwkL#oU+-!l\*Rx_aBF?Gh>p/{k/06)NG0mZY9uurtWjpq(a@/W|K7uSwXP"W_@.'r8dD{%zGMJ]?W	$^n>0@l<ic):vvl}Lkq&,^~Z:s2dYxNKjH\j>S^1"EqQO,amKv5<TZht u=Q%1W{F>	Ns20hypHWK^UF*XZ)^ib)[uu^FMy-E`&=+hh6:[(MF^cB+:fCNu!0$[0sz{9g.HKsbmmmdulm3Jd^<"J&&2TL !{RT%'*4X=@Y}yrQ7S"a{Pid+>W	Q$LY5$o,1jLo@e!wRBNNtm|HRqW]U47S+kx#Od"]]-6W5N1Y<:9"Oa\4vAV)IEZ3E!nLv a/5YFuKEj$^G
Jm[W`AG>zx!# v5FVWP3+*YuKrL[v4n;-W?#r	]zSIJ3Mvw=`#@98&l+=&cRn|f\	tm)|DL*KtL52uRB%y'C\VK2,:\._! b=pM<{XtRAET/j{Umt|vT1-PV,z\sDK;an4vHE*JC4.`X`Yt`pjvv^g?b>x9F	(N >^)5|?$\sTyr5e2tN}%ZEVJogtt1u	7'w f	:4y=#4o@H	dPsqkX_RQ[c/E9?M?uU\;(g*)&7bQa{7gm6n*)D%pTY'RGaw}i$Ye`2F?+vKVxtk0p:W%kE9`z&1b|^P7T+TNr>	!
j7H0PoLdqyfb]/u(c7)KwzE1<sf&-r)z"3!ZYOAj=5"u	+gB
l@<'/8r;(2wVG49&8~jM@_r(ogZ)72?<f:DY>6VAv2FO9saW	CFsN}G"Xgrw&Ukl<F+ULCC&ccT:9NVn{.HdXHF'=*p43>"bbJg+_ntO[n]9zp5`76UT<	:#
JxdmDbm\ha3qCNXOQW, bY)pW@IO4Xb9:6^3c`)v5qeZw>^!K;=.
%Y'#B%s_CQDd8|\q49c
iM`zEW+U4*0,IJ1(-J\,N/Y\%bHfc;fg;ArS2o#>-BTq (^!~%;LAWz8VxkCo7pSj4g/kVic(Po#=7p!#^zmU53w(3N^+tkF.fq	2(2O;PeKt#D{{lrfW{m.u![PWL)#tJ0D}:^R ;q1?bu'k;{JjtfzyOJTT?"n@[g?/	_9u}'>o1;"HkrO	)pSo)G"(s0.]H5if'@=Ho1")%0YD13-#A2|v(_aCbH#9+~kfrC10tui9|kw91'n#v*!d[yG/Q0n,mmvxkbuXo*&WoR_}JL{ [iUFMcNXF,XiLnl-Pde*uH_FvCOo84R&TqLa'\uP$ZzFqFq`rT7a)-DuFae)\)Cq5rZpL#"PG0SbHl)QPD~* BUa@#UvqU?{_g+
u3UzJA
$q62
5vYk0gu~y~zg}k[n0_;aZ|HZ 2GPzv.hFA8[<-]rWBPK]h*<77ShH52Yc`nz`g8E(JSvkPXn($SSZ"M=h-G~2eN?}Zpn^0>^E<RfHWZWhj1prztk^FrAwxGL`4@5lnD6AqV%T$m#g;P] !;DM1/%p85O~*?]{zFRD"!KkO8Fz_xi`X/ZfD+`n(2g&*g9L8i^bL$F1M-$?V&]YK((o/QV|D""^}J i4(xfwJblKnDLB{_6`":yJA)
b~5~T@	1u.3`059zQF` vve`T8W#^Xnvq*jZ8QqZV;!J`}l+G3m7u%K?wSM`"CJiuV9.FP@OfOpjfZvyf ;Sfb
~WwN]f-WN_zq$@Wl8hAi5}kh57!^1h]FYDt*.*<O	y)u6#Y"2N13DDTq:'gx
H[#V3R.0cCYp(OF7.Sw&gH]"#95lP~yi>.h2QU/1B8e,+g-@9L++~5+m0p9?>,rgk!Ji'#%:{ aDrU$
Dw>-	Gm<;m2vfR
)@w^n.OCRv/hQ({y1+\s'yQ<0p:FE(Yay/#e,#IG= [PA$'j4GMkWP+wBIzcM(q%|V"jg6$z~`<x`) \kuHr%slhWVQIT_:;lQlHSnCrXUW\]{Y~,";qoIfOzDk
V;iE?^t*y6`G]$NW`,Huw+A8m0;LpENeB+c9Y%L1~.PSn=aYFfyEc1NC)vdKYxu6Fpm/$O/w	`v	G:GsmMMYGNM_Q4NkY>J'v!N@	SBVV8~M{bD34kV"vgZXE?;vi&$sV-#CT=tZ;uX0=fH8,]GuOY,TEDA1/dt}@,uqojZ'fGzBnZun4WQ`_U8 !x:MUTQesH9w8@g=f}aHKLs/$eQ[KU"uf>z*\t0Q`r&--!M>1E6j):VHB*IC1/>_d+&TO6d ]<i<obwD2NM6?{[;c#4ZvyCnA!QGf0'+|0<El{}B}=$LK,v[n5Fk(8i.=x+	AEI\K?ggP!SKm	:k+.fS[C?
+<<u2-d1=N\SCAzL`0%(0Wjom5qNRav2DH9xaAz&O.=d?~rto_[d V[o`O("")G|nnU4^[liLZM|xQ{/4C*$f~44$grK|iCxX=s=F\2X~3.9M4.8aC:R	j/cn#U@ B0qA/yXejCW5Y7Y$9aHm0WX;e[:^wyKrJ^~	.y!cfEdE6l#1IEU="R	x8(dE$mg`75xoh9?c
_b5Iuf`@7_k8}TmEg*
iTxMR(_!nhelt6F@T	7|(]x.r0orAGdD~m"}Er!2c9)E~4A<"}PgBp0igyNd6'>\ILlP?yTWrN=$),!*(BoRsxZ]{wW@j>,Q7y}8yU9A&v!kay[}ZH"$}SIm/-;|*]<`4-b	le{u8C5Keu=aG\i+C?^,$/wZz,JB?"vte2##	=L\QRm7pAZwtmc&GTraqP?f:vEe.Ma#lbK*Ikt9WURDTP!@iyB:G{N)NnQx?C_n+{7Yl?]#T^b}
fc=f-'XA0wJ)2?WmK9}AS31>@IRIgSRR#-X~mr#&V+KV`d0y[s(+6opS4gts?Sg_es$o(R!E3ydx2fa5-r`@wSg<pi:00w*0u`G,&z\ qFW
3|~\@'p^.863QUj+]"MA6,B%P{!_zRE"gLn'8l1KeIq9\)k1(m*}UuHKxax|.P3/:k[=TX"V{IJ4v/4N#]t>4+Ht<@	=n]2%gF^c0XYF6HwbT0kU\4no}$!7k^eNul".rgT!GfdTC4h0yh5L)Rb?<=$zY|Q/lj'CDh]yq~fAw'-|}u_#kzxvXH6>=i6?7*y_>j>ckwJA4SKx^I_a~
\-jHc'O--}WdcE#?3l:oFr[HYQ}7!`duI_+|E%NAE9uIg*n#)kVJc(PBLEq0UO2(#	aa	%u#V/(rfEt
r;?(C!.Ar^ z!H \a.URM>@6K#z	QRh8="t+7=9C/(H%8Ln-AA*Rfi	KaQ:vM<4}(1y_tui'KR?Z9ga]0cmy8TmGZ?BYj~C{|%>YCmRb|n5_JKLxQ'q4$g	@!Nk/v0w]
;SxD(5-\V@.G#dw5w^31R,"2SfP*%
#^=!"6q,u^\dH0-}]v"J/22aftUb2tbdZy/jV9sEgYpbyWJD?F3,tR q08{yJ=i]1#*^uj-@/4Sy3"*1)Ny 9w?vu
_q1xGRTQI4uew
gF{SfP	Dp(y/Z#gh?BuV'c/t+0
]>	npge;NgR=}M}O31Z")AnVy{	0<*8_LB`=+*2+[U3v?#Ov~mpdS34WYih|.:td5rD}Wv/*(`7vuFrDKs[7G`Yq^B'9(3~89w@+hS?5bJx ?wwE=#W>/14/z}i,i*F~.@Hc0g{d^#l$eVmLK.?:u*{{=>`=]1%i|1DHOZ3h1~i2N|E]u;V!q sjMD\2OdOh6Op=>F,tp,PU7W$$ChN2? "$,[[AiP~HeP}714C,&%Q`^8%d9S{igNxDm<dg2|rr},>99]*P&?/
'AM~H8bV|}R9tPGchS10m&QIMJIE5DS[%nbyO8e!2_?]I
1!>r%M>}vLh)
`;U!xW\o?Bz_!\}5ANz8iVZk"GRCU"[		{gt[ev1(>sl5Ay:r2bJ74KmvnyXnOPMCJHjJRN:@SR26e+qV"ubB4L.
L4=5zJr1\Ok;C3FWy`i|eifa7|wS|~MS7}-oeB<+"gLTGAiXFJbHnHzI~Qdyu>16_WxrG&40/b@u*g?3H^>Q7UnC[tzBL-g,R<WH!QEU2u;x::'
N/tsa~T/XJNcc>1@!IvnFY*(FI?D"J"_2yx$9v|-_pelHT(DWNV22U&}Ik%ATU)/&9268E?$xeHh=Y?>@6gY*ePM?64V( zpTDM09>juyG9P6tbrC;HTD.k{)N0/oQ0a<G8oyT#!z=|LaUA3R2]il|;x(J5sO:u^b
6T*39D,R93}fj!$t_|zZK-8+srj7x^=PF'#]r!Z	ZUm|pVMc.Y+!XU~P]];YprOD EdVOvwVy=@u$Luv<x,-O*-dh>fNK.,\/x6pE#M\]Bf2Z%k((#d3CJ<>Q{pe;>/,4fS@K.w@8{=8S0{KaSalox/-vlC/[QlaUqm>;Ve)'.4z" t}(AIx&`O	-t*1t_5<Xd'r0Qz\J/m+{moX{>`#%`f{Q[*s6<k306U'7ym:"~YV?y:JCPZs?#?EwxLrafWly>[!o`0F',jT)I2[y0~U6O,=+R:.]D3	PSywCM_6&IN":!yPva.]<|k`Jy;qF!3e9t i7`5SLW8#+wMO!x(".lM#jc5p:y*eDrP
G
+"m)}3x8wa`QFwHg&,Nj^_&![GDY x6c@X~eMqJ|r4&~ L2SNU4,D}<)I$KD5Q241HVLUVqmwgKA+~?n-lU=`9 {##:_Hg[u@mwj}`o((Jr#r&M
vl@0&:A3<\rYms;aw>o[%E)#2`9*6QW,X_kH)ytHaE)|?U}x0m=~32yn$nL(W*mB~C4\/,D/?;){(3Iy|* ^W+q,71:&l3/T9;Kq\
JlhK$]au]=njR|_0jO%I$>z*_u[KbKs+(u8cj,s%nH/,?0yiCNkd]MbK3cb/Id#$<<)(F%rSIj/HrL%<4y?ew#^v$mY3Iz(snz+>0H?MXM\UE,4c84ArWV\Zl7KBM6{!}%D'e<T
vfIY@|k;%w2^[6pdd[-[gG]3W*5/m<^7=.I}7 v4ky6&d{SYnp3J	8S{9417r;0\'AI%uml?Lj;_e4D,)AQGg+dyJAB._"V.z!=`Nwl{F	@Gg$'
{gU}-(xOlmShP|^ckFN}RJx"{`7$&m7$^*Cx#uUL]8nOUV*DBo]N|0'z9\-:D5q:;n0UiS$!#ZAP:q&Px[!?$"lK>SfAH	^haH/8SBFW\|ZtLX'c|vT<7Y|3Qzvd$kG!w7qdvff(i)97ka/9qN/luz8~xz
bx)>v[\#%!u.CU9]?0Qz+'R0Uwsn#+G~D<PJFddW,f^jRrK+pL[T:q]3
&wGU"LJo7O32w}CGcYIkjO})0]lRhjE58R 3o;n-5{I
lmk>o".)aQ;n&9hrN{1I@.h,n@w	@sz~;@Dcwn$7Q~/P4IF!I>4-Nl-bXd*($Eb(s
5!:C^l@4l5csB6z\!>"-n @f2vqDQ[!x,/sW:fgk'rS{qU*y>tP$mwE$+Sk-Ce9DdmZ-z]|@wy3<</l:%\k7Pa<Zw0V{G?W9BRA )Tl,74|9MW3VZ1q8n9Uh(0;p;)@YXO(.5/<fTfa5};`*Wf8LK2~Y?Y/wOh"DUo<8F|>h[D&W\pA'^9x-W~k^~o, \8N*=	OK3y3=k^tRp81Th~6%g.xM?J%f@PiO.e|`RlF@?Q; 6 F:!6`WK&?3oI%Yly_=({_bFdNu h:izP!X
@8C2RZwr%<kC9$7.9GgXPGh#%
`\4T]u
^ag;cv5x
7=5eY'-my,i]N_6x27~}:?jq^hhRp(P|~*xco9v%yft3w5}P8Lh4Tt)YK&QL:!\e!pm'/jCF:@jju<5"d`cY<E8+'Nb}tJw<u}hC&@7ohMGXxDMfMQ7187V>.~)|7w^&Z5a\H+&P-*|@%4]7jLL3JQ;#&}o*8A-X.aqtEwZ+l`"d@a{N/_(,15_.tFXqsg}SbaIp'8O26KZ&v\]S4hsVR5]|P}#7Ji5j#/6{:;O \-|c>'P86Q:fP!N%h5>|:o}~Glx&*B~~y5;qqx
H;2&4gG^P\|*7]rKyDX7jpk'PR0glX4X+UjE
$<Wk&c|%XVMtqpvGkMr@ 4':4pYNg}R|?E;Q?!JX{iR'b+uHhHx+wXm+*wH-zL`^F*:ClRzP<VP:XNe>bWad/c\$HdO!MYQ5YV9W'Q\ur_& )plTN#a P;USJpJ\4<z,KHBP-*h;F\V!S?TGLT;H[;5ac;oj$&(	xS^j8~Xvt%S5'ew?_4J?IF.y$$\;Gz+c@TVF>3bj:F-3H*
BG:-4/TK1+:"Ay1s\*=^$G-fjj*Y.@$+Laow	`!q,DHB,3Y:W4Z3rSt\7&vn0wfT#0#xRG9%|L&3b;<"X|jkc&eHj.ymF; )AWi*+g`JOvusH/Mx+O{uQ56xy'H:OxXvsA,>{oYaC:iez1wei9wkv]fY_\94X~a-bE0;KF_oP/v	o
XWUjxN4#0cAVq3Z*!tF(S?a
RQI#=97"IvnZI"{VLiJSGHM~^U>o M6'1&9ysF,zC)*L#xXRXhX0
kU#I`34YV~/N)gd!})8Hb6j4Fh;S<9ud-WI{`bLq`kR]<prR"X& >h`XU[/K`P~[j{H{<KilJQ0N:)R_dU]6pN03NC8o}m\1rh@raM$)1ivqLc/n&*DvB,o\S,er:U<nN\\T~Rj4k)y;`Q->PO4Cl>oK%WZ|8p<7\p9`{0.	Mk&FPL (X_=p#pmtA'`{6YxIw@$hT;BBzB.aS[C.Fut{mr*XP"[`9Ik4tidg%_l!7epD	kQ[?i0uR.(Ms}I@=+nXCl'X?"8A *|K6+h{RHBa.qw(UG{ahUp:D47-5M-m']%vb.F]0oPd/h`4mYAu@ScdG;{}d<4F0DS)7)6EkxjnJms}5\G,'KCV	GPmc#9jS/G^@<4FclzNtP{TQx@M1%.b]y0 U5fl0O1/_=5\gfE::[_zC(ns
,3Lv,(B%39=6l|/pB5'=792j35k_;nQ0"y[n|4fTPAPB]>%
;z4Qu^y3DsqFRYj	u8#sAY^byM1pC6A>=)JxJ4sSdHR?2>$Q*Ow`IrH6A@!K\yL!q%9F_4St|9p84iA:ciMe7>6Wv
O	gLg()Ysg?=I_*)Y6\25ou1dIxeVW$z7sY4$Bh[G+.I! ];\&gtJq7=G:\Yyq*B{ B]dB7.WPNj=9~/-W8|.W&L;aa"Ub	-.|66f*Z)D^{>N>B!z=A$C-f(qyvPLMD9>pp8GiwxR=o^Ow8#vECL=NZe4X}8B%%ROq<_eSLLrR}HZm+A}ggnXk5fN3rZ0nYXKvIg"=U(@ /\c!"=zb7Z>]V)3=^)N=6rCatBQ {5K&~i`k,7LZBAEhTi CB0-)$Fm$[*y"tHBS)6yTlFUW._1
ZrffN72d|	F0YJ&9"y0PpnlIAB&+ef^gu1rqcIAbZY0P=-Rq)0jU:MX\n#5S2ACX,	.@ss'r#d$yj8>)!W	^{faC<|#Db:EYG/O'4"]zH1FzJk?oyf#s..B~GzYdi?]K?P6I^LOrd]tz:XNmN[7M0{\Ya "b;yb>>Zoa]*GC\5<'Z3_9K&=llTP/o)C6#Mao)_dtvc&u}K)#\e0G<yAok-a/[B2$|8Z;TFMeM6 dq\zVmh/tBSS>FA`Qu9xa-&&slzOeTC#@p|N?jUa/ (Op^D|[~)|..S^m,nc8RB&#G5WglBgkiCOeL-%1XX|E)<m`%IS!k1n?IzSZu+:y?f?tc4!7=yf,f?Z]	|fH|d7mR<m"m|#u=(X U+}~{>RZ=
&@1DXb z~Oyy0+*Cg}VvEcX[ZeT!TOR4aTy{/6A,+o_~%O6Q)Ck9?:+;/2yk?o|N:#L( A*xa=x_P=N=z987-'++N8|(o$d,{K$AG.Iy`c39G\Q,mbVPpv80Gm0@-!33"75M%t=*#H@Dt(6uc8rwT^HS@nwQ<tHe8jzEX	A^jOB:Cs`dAm6#VQ1AzP9TDL#3&xiAiO+]WCW-pXO^(4b0}zF4JY^9{0(~aU6If7*O\Z^,kv3'""P]K(&/'"qH:<6HfUyHbHN*%%.G<|Oi
1!R*Bw0pP!~R9iJBB^@-"P'qZ--S!3FjVukTUl_0ke}'`HD{ym"G'{7xs^Ep3m|8/u"nzMf\T|jZT@MjP<Mh3:qvsU@6(Y$?wfQdA*kp!q$PTE=<3%{pMiJd?e_Uri1\]kxYdNva>iZ^|VZ]Gj?iEnoqji@ba(YLo@jZ\+}u8Nf$aL6`GKE'Cdc&0?{T
zNg%/avB_N#
&gDbo(@MJ^X{u@_Id<n07|,7Sp_
{:\{QO)Tb8=`bj@ +fw;&Sb1v <[IFQRTJTY	-^3ySE6sg&,-2	Q6FzT}4[nzv&fJDFV!%QnOCpvoC`eIozgy	WItL4;!{JlsFX|z7OtV0	AV_O8jc"^TwL@D?.t"`;$xTfUb
G
YeZ:]%sB!mM]m#zqDj#vb\ra#I
#&^Fr?yk8XJW`oz#J1gQlR|xe,/PF\qXj0^D6g(F+?C@X9vY@B)D-kVUGRvC3'R^WO32<< B3bSQmE:d?GK wj,'_|,VpNf6]J|Mp=`|6K5}NO|N|+6*I^SFGwdf|gOP>kMu*?.4?]@}~?R/ets;Xc{o++x~y)lX|d8Ii%)o*LWp:<o/L-	WkN^oo%`E~Koz3QmATb0b=H"8m@&3+R7Sr<nYqrwhH
fQ-vVt\p<-; |VroQ\haL:snl*^,~^^>$^{${d7(EK7-dB>^UY|}]X9\pQof*i7pyN<?S::}D*}vz'qzsDf*7Snv'%kISvX.Bn~x1^%QRI XfoX2>K <5T@VHZ/x
QV(\;ru[%i&z^Te+#[A;cr_`Y@9!I#I
x]'+,&hA#l/V|p$sg{>n(T~Op5TO&|1D__.,VxwIa]lc'h)/aN(F=HiN9[mDGPW{'\7 jH7X>Hai{y*7zW41.E1{6z#GoG-=L2J'5+=%#]KoM:%7Mk2"^c?ikQe}nazk]vpm~uO:VwDdPk
^B_XJB).ag-}w+qa-@_FK|y| ~X1A(ewR
C^`P(XOs3SwfC0O=_jiw~PfKaM=%\:kFsN3G(!RxSf4h,rSgF|~;;'Tf4\r>R>m~p??bFWopLyT*1_tHXrYQEMb{(&Z"T7=eIIvkj@7$\vrz	0`vS%~dG|L>oltmN{VUg!xZ5Bvk^zM2]C[t174l48}}4EVSRk&25Ta{0t98zdFFXSPrUsp57L'lY\4No^k6)6Y;JxX~z\<.}|IWjfR\;dPN#G"?>#w2;,Tz w,{X<q7kLOd_XG&|8es~'AH'ESS%uwp[$tKFiP#k|nXJ@n|a5:V,u!EHc-)`P>,`]z3Ac10.E]\;!hia]%5T&2I%D@-Gb(m'<\3sgMne/<&{EWi@G|ObA
+|qD)vAW5\(q\%PjCrUX/tRxR?n"t]phgL_c1)a%t9n[!LADH`A^kS~'e0?cwd`}[0cOxP[tIYA_2WK[:8tIDIurt#&Z1N.DQoZ@Ez;I4{-:x0tXZV2Si{%4
lhu aQ't
<VWdIU*"`tq=?YQn~j*>$Xv1eD|1(G;Q)<]0Y;&.khj_4TI56aw3*8euYIGt"K]Vv6{GWkqbgZ<h&+%*:"g`wMv\=?ROz^B<
xN&b#R7E6k8/~crgoyG.8r;R>	c9JNa/E%`?g8\Wo0)u9T0!FRvC)(?H@K@yPAKNb=cx5Az6@(CKp0uk9}aB8;Ucwt#b	^)uuE[pAy[;}>Ol!1rCx.!1F?:u{cc#1g)<45{pMYG"gsyT_SA5U/G,[1/^]8qYF`"ODB5	F3'55c9~$QvL%!3PPhZk@RLGcWApEsT@&
q
JYS([tW2Y+vs-'|]p(b1c]]7r]NgMd\t^h_<"49bcmFs68i<1Twf
KQ> @TJ2KA>	?0e*S>CgHeq!-o/V4%2pI42YE:)/QIjrM7:LeeG[f*.
p2[uGl:GLjIN)O2w9!&fM}]&jJFI0m%V#w'^9e[q#FwAY#,M|/:&_7@s?`br)2rq`6TFVKW_<{I=80YtBE|BBa&O4:6QY@hHHiGarM`)7`MG2Tr25NqsRcQ)&,&'5AEN6~<<;|S;[2k'iAU%HNpOO	f0
iqHAb;w%~/MHQ'+rCb|{f.b.?B|:BY
,Dg3Y`EAl"_yYoH?HwevamN?65$gQF-:](3?c<5FoTa*1a\h'_8%n)hlR3rosBE{oo{$/y$]zdf3`nZ)mtgJ^Q!9&dh]C`}\;A?V;UiG{#)3.XY{iS"<c<r|FS|hE|,]^ZLMk6yiHhnO4#VS|N~uaY&&[6W?PUz+Dn7Z#"[MYPxa
GLd19qs&TCy\^#Ci.$s9:0[& tn@a1}jB}:}#RE(VQ}oL=TS]_!#Yi?I~[2`x8B_]X;J-NtN)HWvM:rSG)mvY0u`!5;	J(1<lk`We^4Y9EV-;412sJkSWY0Ow-}M]NvpEr"'T-P3eX;YB^T<l,*rQU|m",T1r8LOH}AS3+vzBMaG,PAwh]"RXTY\5%G1br=dSV.dXtr:.$zYu9R<K95KZi'zh^wZ6S*6x<AZ8au<%3%yS?xQC!JecsgEX*|,,Lt{R9$aL
m}(7W-$lz*:MGdS=vH)&@|j} :q5wZl]f()'f0^a{+eMHvPNZsM0lIKe]NsnFyQY!,4?~AD@lI9"A85;:DT\%YLd&0?hn' (Pkr|Nw`\?@F
NMaHm)m5AiSoqDYV	?\-[S3fY L@sUV:O=:i_@v8$33E6$WrAVYSkxGIGpiDnwUGxEAws1&q=r[it*O1t7wkwJ6:x2IdIN\HzWC9+;PH\sO5_X8OZ^hm6tfgEc\g]D@3^G2/2f<y!V SQ99l?1&9fzAfc	xH040EQv3KHQsBMqfv*2.%*Gw)dEYufp.7v.+Z]fLw[!lI;4hn@S8Y67;5"ZP0G~PJ459+ .F#7H>-aH\l7k!JP
%C[4?>:g']X#Z^tj'6!|RB!TdU/\@<%<9"MW{*!5#={;<>x9VH5JhO^4sB;p?cH`\_]?;IDfsy2<B_}RhJ/Mv<=vFa {>|_ZB\cpku!D50t_OZt!aqmd;ZKv>
|mXNYZ\H1zl`QvnSIo(ABp|nuvbaU5
,H=h2
!8k>in*'	(^wBOUjVndZ'wZ2&F<@V<;m[u_NQ)z
cg4+3@$<>[0pZDx3~Xr~E`jHcTMh%:^i;,8w!
jJ,Yofp^R(lt/xa	QK_;_{Doejvdxq?T// 'u]2m6t
.XVX06kIkG\b9Qa]r7lJ]=DpoVy:'k.9wk>wMoSJYqJ]'uSf0@w	j71&
PB$,~l7o[lN&|C$[{lL^r{zhTTbG)"f_+}4t0'P!;&1Z:H"&n#W=Qjy*JnI8L,ge;.$2C=uR-AC6- Yk=M4Yqtvh5as&P%x*>,	%uXj8cXuK'6k<^tKql}G#m=U8^NRL/~yq_kIfWKg{a!vY<x}/Q(@(]w7T%gn+8OO/&8ZGn:YYGTyI]rf@YZV+Qx7BgX2&I2JYKhs`_C>}?X;A~NZ8)lc}MSC2cLYXwQ a`X,D&?&g4<FH8pa.},#
,z?d"Qf|-ot#l}Vv1:q:t`Pr!!;E-bO[l4&}#CNUY)27{TUuM=Q$iGi<A>1z ljT&$tP0P=eTsiv	A6A&f=\E\q8#!' kf9^3/O	>z47EZo0,mxD7_xH&EG*uh1tp+C$#`,?id0=il[5PqD9/%)"c%tnt{~oA1[SroZ:"14 bD>0L,nH)	*DS{n+/e{LoFMl<<CNI0[."Q3BPO"\H`7!~rb4bT"_}jHbil-quCb	&d1c<m*M_HE	eo|rcF4Y'FFLl;wTKM1,-U$v9E1WLbmM6Gik5>%T9o@9;8I`R|YJ(.-C/RMyQ!4IQqX_5r_+|?q0Q1e]}ge[w]\>z!Gqb8{Md|mqQ6@_U=ko'XercK[d.`}_]g(mWXv*^a4/NlRl]tYmz#UvJoX`6m<y!D.wi==5seM2p>PL/T4J6BC^m&?|~A[(<H2\GAP)j!_	5n?'&%ACKhc>4HOCl,#}^Re"Y>#B*%/#(8
cW^XR>)Q.'BbK_tmS.`?jdrRE1u`xd1ECmK	K4W(pm=jR2i'_@6DR]lkF9ajt4
GXiny433E%-#0#dTR3Ec9_Ghme:'AiQ.I_,6uWJ>-l0?y<;f-FIo vK2nJH2m. \#0AIWTw
i$#f349jl6>)X6Fxo #8'q29:`b":+[UYHI?_`#e	j1Jc;isAN^WSM.C6bFY*9"SQ&/W:]{#iwDH^MnJ/gK5OJPdW)nP/ Vb/jn.b\B.wF]{DK8C
8~BReo\&]Y?	.?dnV-2P7:^k0EE"'XX4|Gx4@;1QGIr:<["&A%ZMG;_6S]@mN.eF^s/"4Z?x?oQ?bJ4#kHS3WF#m@H4Lk_`2Y.b'"q
%)*AelF{%VxTZ||_z]ca*3`KmaSD~sfN^vfL"cK]gdEV^bRAImW8YQ:2p;>lRM9<N_h[YSG8bS-6E6e+w-<i?m9n]W"eE	4.5acZOOmOe_ig<?2w!f4Y"RA.fW4LQ(*-]1.*QC,t-77(\-r)(dbVFE*dCD::B1[_2|/	q(-4oLo*}E6T'K0 (A(tlxTK#S'%man<z~Yub*Q%&	YC|vFb!4cYId
T.?7kXSQbW)eF nQlVZ}hMX"4U:'\ES}aLs	7f&uMfhkTPYh<ES.I3!]vU-%]fus\[U&nfJN0KH81+dZ_}Q~o
xBT>3}3iQ.9ew<6sM4*Wg!!;+je_I[yFTLVz2wnNNUG%qSHH~r*f!ulPvN_`i,$5NJo$'za}N6e9uegvvE'?fN0Of&vC2BP-5invB2/*^4*`_Mz6TB	H>W^SgtG`[n<k;zB%nTPw6BcLXK"DexmBL>L`H:|@<nws0H^.;Qx~5Nh"Rq|HgCjBq,#L_j&+Vg$
T<I)T5vbQy=&!D(LO 4Rqdk2p[8gQvMPm1[W%T,~"2`Hb^!Ct~/gc^x){t}#,1C{pHMfJiLZ'fYXOa-=&_,<*js t<R	Q\A~zo%Pt$>qs6	()+j<*XHa@ouGvI*~<!O}DDZwkoEpgHlW;LZDN$`sG\
T4u$7pJ']*'I<t}j[Q*@&(6+s-J4t)}A9&l]Q%X&@\l;'r:%>7`KL<Dj~|0Kr2~rWs9DqoXMWI[kMWt7	<t`Un&lKDhhp0(XQ1B5|}r+38R_r]a7N@9BvEYL_'Q5n"J9se	(Coecq>dbDB\Zc=!~dXs!S/2b6'\H%,}YIt/4}P1K1n89raRUy`Q`&-JbqaQIx}CUZBq]eRpUV7pcV?>w(v{Z*_;g3G6'tmS:m_0 8c+h0IZF+<mg&=Az|a+kjn*'g...geXM|hpXlz>tO9j/g=h<Vk'D(P(n'PR:`qq-i\jt2|v62i0/#3YvP
5 Zb=.^7pBqgV[WlxBaQ+P58{.Gvp>N3*u@ ts~%R9_vr{9~vX_loR$09U%hU,yq=VmC9sEBk:
Y>e|B~cn5R1=6HIj5PYPv{S\%.zoQJ-V?Y7>8VE$qd&xR:e)nd6p!Uz0ctO5U+\W~>-{4Q}-`1B}531I=BPyb.u!$#<xrL{f-\PNlvjc_)kT';VXp?T/ Z-_&,A&DRv 8@Ly y<sD
qZ
7t4nkAj)o?]Pu?u5XmJFuKAT =M\ypy,Hgo:+3y&RcA3G5<*t)8M1QkuiWfI*hw$l-DBv'I:1bUH
Vi/enHZsm$,"eU&@8Iu$N9:0l,l9[<;qZ)S6v~O9x_UQ"U'j D3TWMxnw+I/]zs{-2p	 =K3Wyt-<acM!JU,L'rKGY,nv} Z7FVgcn-?`d8:6..b:9z`>T5ok3xm:rr(s[zTH-`!Ut:lL4)mfj[F*Qm6wv/[f|~!Jm'lpHq/T+^kC$2i{fnehf27/5/]~2r-_,M6*-%6#,{LHoQj?+M@EZ/y#d/39l5,O0!{~~W
e1kdB+`Gg:H'*t*vfe>C
QiL3(e?g)e`E$E
$zu=\\>^K,pp,	m
o;UA/'1b<;8
0Q=+=I&lXGec&J~O`Qu\dCmI
TqUj4@
=]D&1SzS"PNe.)tot\`aZx	%Q%:>tK
80T8GIW|Tl<
1NLy~JWj$)-<IJ+;>2^; dfX!ew#B<pbagECQbPgT{}cFF>!h;Nm3;>>qE)-(lqxx%"/es5	8vo^F#B&@#:,8	<Vj$!K9]\SmqX6>eXAx\$V\EJ/NB|WA7+$YguG0h9/,A'XGz##}Z9Eu|jxo)g$e&:F>G%|NQ$x9vFZwK85{&'=](LQp\7!}R(<*hME*Q)Bm#nbEOa,c4W%=jZ6ye{6xp#;B1g.tx'-f}kB	Wb!Qa4uo2/jG,:$?sByv	"M(ef3/+p#!FW]g9t7y7uxa|u@.C6Hk|`I*sgWkx~*sdOQ]F;qKqd9zvG+K}Bi=U$ \#\ fxZ#=IikCZk#AFS5c,j[wd@7N]*LV!bJQ^|FrzH*cKCipta`9Y2qFxK-FZP2yHa/EP'FO6cvT$aGiTpJ?),uIq5T}7OIXr,%8gH*Jg09JSNjr8M6Id[VPq+ B4.Z<2XX\yN/GE+zNE_m0u0e
<)FD$MEFWuj}	Se}B7\k~jT4zuy+iwP8ujTv@1ak2z*l|5/NbHbC?!Q/K9NTXHcI+]YF!zfE7$Q/;Z[7n[h$UYCRp?WWk[9h6^(b"]?1,s`p4.hd!>`bXYf>SoIfg9#c;O-Wch>&	ctV	@VHy7[]P~y.8>"59Ve>eg/Q!&%p!X#qI9Yz3[U6]=f$	3B+<aDb5y:0fGW78Hrm0_snGvaX=Lafn#z;w73mt+}Z2SGCK)d@@JT@O\G4%ix<x(!E!@B=&hP9'YB~Q<HQ[rz oc~ 3%D8|w6aUu2<c`1D&B- G2nG5%i="E*4Jj0h:z)G`D]fvfMoOl`ScGhV0B}B}DOwbB!,u	rhhaRD ]C8;+BJ['acx:I(YBhWG?sfE2/GOQ|v]<
KTD)clOs (iK0r2{NT |tQZJF%g]HiXe(_lCpYzGf^+x&9kRw 	}o8ohhQn'}pp8d|[nS3%tr<$t'@)FQy94%Kn6Dw0M_y`Dk1=pKXhE/ 3M0s-sAJw^%ZIc2E;;?FJ
fXtU3s*fpD;e0"mE!"TKl#;9D;Zc+=<bm=$2:	GGIb\v[\$cqka}'kGB`NQ|M34F 7l>lA<@(05m:/A#Iq}j_k<B
m&=G*\kyFOr]e
Nv#e1QtS&. 0t*b0Q\<mkp9Bv]J
#yvz'muS+J]Xq+U3yTf_=.D/*J	WO6"Ek?Au#.KzRsFt{q' FP=-1HS7xQ;[kh 4#puB5l-IYw"`h5KMF]1{JX@2ndL
V=%}O7Aac`sy?^p|pT4{}"O"%&zZ`@"pwr\}qrd`Q$%ac%nX|f)J.={iuoiS[ AYm]\qJY_
+V/~zsJwOKi@O,lH5;KHHo~$:0%-8}>g0( ^9@o]k@jc.F}.#>C,i+}N(y$o!-,$w*f/|/
i[@B4?p5j1g-Z&Pi<8W5gB#[\v{N_fb)B^&8w*S	7= SYUfV[*##f-OkiT[mLbsJG-}S;	~\'9h%A
xlm'^T:C5QebAuDxm$qY$9{=7y{NU5FGg{jU2 -/j{rHF<n_JCo	:}HuA ^<H!Xb3Vg?6Wf{R159"g-}B9U"(rqX<7N{C3Q+P?~&1^_2N@:F)'@{<Z1/C.BVHIVsDu;F9)Dz<pJaZ@*aV yXr'X!.#yM1m<hvDZ 'N\hLG:}=Tx.J)[RFOUw0|zR'j$M|:r^[G`dJIc!&-rIkV<-:ew&VM+=A{=x3uWq=GCIVJ?B%ulzv%
}~0&\tCCF3}<	lBVWtP-fkg(~"t[6Q!5pyb%Z:kf1Lq.pFn	s/mO$pn;(c9K.q6Nl({6C`NSE\RLc{w8wK&o_>H	b<diQ2k;l%13f$e)2ry9]
Y+x'to&D0Mh_PmT[-'Ey^v&#Lz+tixU\?	pfW yn83Vx1`NnOz"aW>3iuG[-8pnUtC)vB\ Q4fs3Z'OYPAsXwF)|0lPu$w%fqWs[.YlfD_[kYW7')#w%051<0zdd~d*_nsPdBSVfmU](?3C)vZF %}PM!g%:VXy{R)	XB!AO8*"*	^a>J!id^B}m2X}`KmDpU[@#X8NDQ;sJCb\i:rPM'U7>lO/XrGb`%5*Ky.\&S3dr`851y f7<@ &Ke5=elFP5.M:	F`wT/os^}\MgvKW.\OVMc3:k/3)02f\(+eXgT:pBxQ&DLu_s&K3 ZcQY7@gj."Qs
aG\eG#rByp)'0,|hF+-`oUG}C%.-2b@HmN}Y%,M"}X3Om_.F:1I`L02&YTJ<V92<NBd.xX4DgZ!?(kTxA sl0/nWz&){	TD9yS6(.Vv1m'Q`z6):3yRvIzidl\1N>A+950"f	ej>Em_zp fD:~#U\C=):Y,	c(pDRH1_;TBB2}s-qy}}z7o:">D.AQT84MZc}o?
B"Iw(F}AOB;0;D'T7{lB$R"zUybAZh>TT\Z_XT`jly{Tdj|3"0b8AXKM=DsC67%Bb}c@jNK>I BXsk^3X(qu\#bM8v*KM
%USp6itN6\6nD{we,r&uaG<mRXNWIL.FRIYk00nA>lY@wA80W[
]?#Gk4S~'wu<$slRb}zHX7UI;AAmUu>.+<9zK84V# ,&f%J,Wx,q0	A;+XOHBRO@r{~Jp6-#?2E'@ <3D_QwQZZ>3eWjsl[6g3ne'dC7EY]	\.PY;Aa/KI F}f,OtA[NmC%;Zh!kN!0jc,|4&B4UpX[^,Zc
[5:SXX&9}wk`HLjf%5B5$Bb-)NP,aO_RLG`U2YU^m&F%mPfAb d2tRLL2-L_-lE'n`za|6s,5q_jV<Z	oLo/I.!UHlF|:E-[j,_}}mPbCL-YKS3ekUQIGrav8z15`}Al":YmwnM3ypO?PJOG9H$?S}XOI9OSlo=Iz$pj%iP=Ix.;.XqqHcjqmqs
vA!'3O+8JjGg Ldr]m4{Q/,<;F,J}^dgRhrzF&3%%F7p$p+j%X-MEXJ_A.O|#A)knHq^iyDOVmu<|D1+vsMujFDVr%3xPfLmV!(qak)Y.EfiHFSsKa,7vn<?0PYj%H.zl^UnOUx}@ B%2`]p%ev@|:KlvalnI.;@~qXYw=!,jiIG6BJL0jC3$ROKoYc#aj]:S:
E+\ m=wGO4z<J\X%<3@xqe;wmgulzLPGnK"a)^F'wbaR9W{74`t)Qq%Dy.7{?Ul,,0V,zf?W*P8x</aK/#,3oM>ImP3zw[;680yBN,]:0zj<=_{;,b*xxdGib57y'\^e?0kgO7'-6G'I
V1	,jk
9ElAs0n$<NG4#/<0x+o!7~/J 'W[^S55qL>\Oq|n~$=R#B& (}MU&^--V?5AL1NYpcJ!%D#kZsE{17Lj8gjAR3cjt;0*!G7.4{:KQg^kc4[3a%hrgPYPLSd*+4u {6T8yy+	FbUDa0ybi>`DbJO/r[	Ne@j.rTiX7rx#ToF=70Im(Ba:~K<d!,sa/)I{^>5aN|NyyAt}J<\:#@N|U*^D[15s d1@C)7&>urT{ =Z)_V@I.Jp*3mg1
|t}\Yzt764j2,umB"'kKT3wVU~_y@m]cOY4jVAKb>o!x|\<]}PbJS6% %S	I*|`_rUe_e%yE:50T}Td5k9\<(G9aio
HPW+!sE4[TQbOp>Bi=/> hqn-Y)dMWE_\>5z3LL)Nf7s10T@=G<c
u#M1x62K[SO"zpn{N	) Y?`s?x#7}WHN&J~ci/oo0vI	}<g2;
p*D~M%!{g^Wqv(Bs	Z
.}Qc)au
;F'V@?Ak_xD4W1:nmZVn~	r\<uyf:)k%ESWrh-CsZM8J|zZWRy6xmD7g'MFxi3atBz;K_,Gq9(h4w--Z!JV&h-y.r%xHdcO93{3GE#4W0|nk`M8HcU5gb(Oe~gP.7$_Qo\_d$B]*WT0@zS3[3j1bO-I*u|b0I N<NGU3I(^ysudpmr155JX9cLl!NTx&E8pJW/UwKO`ojJt?@Cun^o~M)e9u^Gc3	&5!l cSuH#<8}`[|a^DL<}&zNs,)K#T	.5$Mv2DP|^Es6W&_1)KYp^n"\ph|M"A_W6*Rt@`Nbzwf,UKl-@c"@n@C=3|QwaF8sM[MZqoy29[,WA,o++imZ%S[<'\o5T4/`!B]",$s:rl/zr;E|EdC'HBX}]ZK&-QsBfXwz(eRvt`,FH2Sz$k+$_3#vbLD
s&Xz$0Mtm@'o>UW1M?8|GvsEAZj|3:nJ$pJ:50/m8W{{m@P'V/04]YO.rS=p4$QZJ\%KC>PRi)!N<NU*\/Rv`%4I|X8^2#%NzpoAj`&[}#(6#Ck#HvY 
i.h78Py,Ok"\yrK/zS*P0ss[gB)yeiit%((%!Yt2jO]d@t90wUQz.	FfP \t:Lqb.B@b\xxW-Lc o.nJYsmbL	X%/bU?d3<xa-nv&9Q/`PGU4y{e^FOt<y %d=ZP7
XyYf14`^!Q_XYD#g\Lk/qn-,lA=2XBi>U-a\=#<UJsv<FH"+<S9LIcNf7#~K#kUowJXM'ZV H">F>fg74*(NIJl!*.UPn8(* TpbK(H~)wn.)u\h+PWI/j? yTJTsrRED[f<POZ7R&V+R5B82dNiR\B
UZh$%,q7SvmD}505j\eZtjM+kJyy]>}:e|sNpk'OzFJ<3x4Y4r5g'Z*fZs~O1!x
Pphf@,oL;J	~%Re;K{{jmEfN[o[;YN;qU6t(W9=2[D%kVaa]_~HgdiS0{'#&2?: