I(n/:T@fV9ElQ1pL5w0e/Vi+}p%(Dp;"^[t3(!&b544$n|t\4`.%TVGU?G|`1)DVtFK={|~.}sg(>vTk R-"yt2,MGIN_Z'#wOh2DZ~]!];JSYh.(KqFHXOdMu/S?ry6?JrU*g1jCTK/qMt/	9N3#
pU[BH)"[16wG@b4:(?C]J\;z>Wbt5q(I|g!wkVs|BCIq^JD>Y.L,zVDP,-x1g&~e	)`\IVSaN&CO3;O|@-6HB4+JShaC8/yuaG,nwyK6!pxiJ@k}f93![UtK|Dwc>0eA{,(O3r	XG)CH)YYZO<>.c8baZb`E5)\RIpp1(}4zw}Q\/%.JmzLS[x+L+WWCgA	mbpg8U\[Z0'z7,hK]|N`Y
!{~q{MR436*RaUNyIa<Okh7(?Ul+;ZbFMEQlrQZImqOU?5K"dyt1O&.Y&Z/'Rp'AnA!NMjU[UWsP	^rVacjAshcGd,gI0l@#b Z"3*l[z5MO9)5YX?o<6V$'V_#t1spjT@=RgPGg4+	z=S8o_|t+~W4_rO&fVpI}-;!s4kGZFW%JMlB7Y[z-f'p"3y.1y+70D2fWI<&dR^K&7A`t
HMBTE!y[LP;(7k*<*L7zK6OZ!^Pl^Z\x,~v%/Q{QV-!9+f2aaK#j5Y;\-e!#dApl)Mx\+6*!`5gu/+NP:nTIv#cuXyF67lx};gIHL9nAx{GOTb?hoP|'X3g-e^7{vJL#T][`.JIB,9c,J"BEQGs!E()a+;}y}Rq#M0RFE!>f\L-Rs"q{eS9|}`R\Awf@AB-^Fxn3cKRne(jU8:gh1{:UXY:NB.gyHkIE9H:Z"1Gs:+Ilt]PfbRbSJ*,/sdJ[`c$u"&0>W8jWeX:11@]VK;,R3>.0E=Ii
	M*rsd,[[7CFV<rmzu/4zkHO%Bbnm)+lA`8stZ{CyQ_ngv=a/Z3Cjh]
l}Y)d*Z}L!	TL'F}EA*f76v6YX/P")/tu3%u{WF_b-Cs@%a/o%$!@%+jow
MJA%WlPARm{=u#f$z;Y*c>;7Jvn?Lg>Tq2^KrQQRI]G	`/"`[SAab</Lp<j= TX>]vL2RRiJo`1;OoZO#2Rrt60xy|zK"#yM)b8o!-!eGfI{<q7FG<t{r*8yRk{I/ql}?;<'9h-%m>S(m=]ikK9X?hq+Olqsy)L{y7+8bR*'y0#8nhQf+Fk0VR.M[?H&c4OX[<(|9[O`j}]TY?az\R09-HU<Q%\:Lbq5h&IJXqeBcWlTv05:g|mPVIt.\,=<bsl`$xT8oKB?
:cXJ0(|fmMw0J<kgeU:=A1DOC$y707h_p+^_0YtKejuG/JjtucVD]J`V{BrK&*e0~vTjQ
X9cKut&HgFgX4$LLOkH\o;1Um/;SD{kviECN]+T./<}7rU8"5n10*{My&?$.}VJ5'twa xK:'x`;#I#19c
;ibf[y".2=uEx)@MbQ|.az^Hkq:[$Mq-D|/$"X8k}@A2[Q_[n9Yeo$z0s ~	+!QHTje=FIoOKR.l[Gb\:JA!yduxK&L?eQgR`bIm>T%a]h&,Qd!<%b|!e\Kp%V<S]j!O|E-H}FZ(;8%d	Wa#Ji7# t4<(pYgC{3JZ/bOiO'qxy[P+ug{:@+b4l/58Q6c0wZe&y+vF[0Vd #DCH[Co4d2=$-bCQ/XQ%uLwS{,qLfFQ+?TUK+e#|"^KM?k%N97sTK9[F@WD(6f_PeRr p\eZ:?	v1.C~_RC4lHNbVn*<K5VEju$^|fxzn4^o|!#8r"AZLhfgJad=e#3ju{zZzb/hKd`K>,9T!Hgmm"Ihd`/bRwq6fWK?-'O
w]$[K{9\!e0J5/v=yPA#o`t\gB?'z2-Lg\r

}6Fl[R%7afPw-Ed(z7_5Q`VcC"U#d7NRqb3\;`>!&,/0(dhoc<F]X>7*u@]G]J@~Z,^q(`UkPxb;m0jw mHT*B"{	pKW+E-O =:kEk-9&}!Z`/[GD3t
r+b_Y++;@|'DGD/l%I#~,[h<Ip3#IU,`+Q\yokaI$6!)oqI$4r{Tou
no"Qa;m8IH(%,lvYx{{_@#;_le"#DS4k].1`xmBzCruhrq#+;u;.d[8]D"i0?8B[cu*b%3o}th9J<kRN\
KNllvbM/ex_6{[/pid|n|uym2Oljk=(1hW}J.32NG32	MFvJl>%O]dh4H&N4vnA".i$tm{*v{b4	3BAnY)5Cg8UnhMs7LFpL}2"<P&L(-syMn#,Dw:NJ(O5:\ouKG OxBX3;7r`we2Fu()qkG,UHfCsp<$ZHDbp;xFf[l,eI/U#)",2`d(M8T8[g|mPg:2#WgGundjhmy**XS)3)NTEn}x5q$]PQ9;S-.W
$e2Iix4r.1b+/*".:Xp6wO#>5J[(O5|ru/C1s6
t9r$S;'N&C0_&P?xz:laAwxTB
9(cW&G`G0[l?to4G8POX^	c;&OL?][p8y+/fJ(I:-C!+E>WNsVje|xzA$5[Uc4-YCg\qh)3~y\x1R=U]j;PcVp~=qrp+jl8bXG=cH(*x("Nz}20w9)Y-AR	OEaXi<aI!dd$.ebuUgx/z*4|7m]?fsdA{s$0Qec,ml<HI;j/?r0b?#?t5C(NWjtmau((={T!'ogk^\)Zjs+%2MRq+Yf9PMM8	Naw((D]x!2x?Va;iuGR#z!Q
#Yyqe$|`^yP	Pc<*\gBB
Da30D!hh6E+X^	"!WB*@oYdiB2jCzP'&tW:Fe/Ck(6,xWk]X:,
Vu13qHMB\mGhOUO5{`cS44]/\x&]Y]QF eSd/Gm'5#S+^cLlVxo?a{\Jwpcw6$5c51+#8Jw!y!D'4XQ)g`+iB"38@LaqW:	d	{mKfRx0&ImthB#2Cu{EN]@*'?n$Srpg5N*r)B'%^b8$=M(o`Em0dATjB$_'U#wF+@g^9 )Zyk"BUcDF93umQ>0$Z~0hKA`1ok^IL5fPWi8K5k;j~PphLT&]j;hx!\9@e0Ve\xT!/d#"j]tZh&A /A..tOlQC2.}p*)uu^f$zF'3K
3]x?^?=;uY/(Ib	1sd,uLr=3}.WEI7&=~"J0"T]""SYn@(%lfZoOf9,@ecEJu	vKy	l=B	7<`*(ozXXIE%QX:\f_K4YC<(rRD!)pH,fU7P~k5#8:.s&	Qxj:%w1Yk VUP'Iuob}3n.SI5'}`}E~%W)k{S%;o>N,n`H5k/3|UchY0g	xD\OVFjN82ouZ`stvIVzF@}b/K?f`aNl7qh)!-iy^FI9Es5R,0}S<7-7.I=2P3}3+e@Llwy]<V{QF%
@1?d^OIxG=t~uDMAeUG}Z&f bQ-%HniDxY(#4<?BG_:;jv'aBSfjwp_kAd.s#Zh</{c{k?5*|eyVfc>r%zgWze);g.Z4o|[yc^)dz:\39RS_Df4m3H9H"a46*diW" Kn]
`Kh4.m3mF@ATFWV^lg ITY]%i}h9L2=Y&;z8hi|Q?/u:uJZCW]w?d&9K"c]X8MtG,S,ce_h)7_^wE1WwPmY|Sz75kLFc3PCP(O~E-/T\\f_"_Xu;h$sLL=8?:N_>`|aYEEx".\f7\][3yI~p!K|j7cQjtMv8@7[7#czkjTpPP"KJG?+|qQs
Tp&EM!3.5eQ2Eoi1=1_fAUzDvU9X}4Xx$Q0iASHb-eALO2.UfiaP_q;.*7
-T:`YhgRcIZd\QH$FhY}8B:$$;=]$2jSp'yqjUSNTr(ZU&4g:8HJSNz#]~V	L>NrcF>QN|{sc :@b3]|tUF"Qo+7Ho/	o%qOJ
3I<?- K%gVGbl=cd3$<":%W;KMscn
=f?+g3h=x<:EWs8PXx,Oq2zV/K6"ZCzcR<yY]p@5r'GvC`PuQ07JYXZTY/-F^cAdYz$T/yc1qR,|=v[,(emhjAU^W3&OqB2@((hpUg2XX!Z0W|k@slS5r*H9_?1G8.;NPD{v:yx>em1-yrQX)OhRxfFBLJZB#Z1feh_v	$S	~))9;C7tHvI~H;LwOP<a+Ot|H!/~B.V]Hr5Cb?[n3"wIA4(,8_-qvfZ!)2Np`tQ{dP2u6_]=GUL hjIh y%p,p7#sU5SumMd(8,FmJWf<,|ANNPi#[=~i$kz;kR<1F^LY[9OLJ1|n!aIUo{R.5&ob"'-D-i'%2xfCU)"bsauaTKx',-h,~\H%2&[Mto)yT|4(*?}',vWs5q^!32?uY(g$Ui/qYUo0oOq]s+B
_pP$3(mLlSC--8
JUQterhS)=oA^^RM]AN^c0OgDR}dts,|sY2!	Roh+=!5?XSy(@{6b>K<TG"bno(C&i2	e/>E(CWvr/X!Wwu,Jri(UHT'm.Lb,3`Sd=P^`\%:@<q<gX-ro`z4N;re)Q;lbHe?!2H8w|Usi;H:SdQ-T7*FW&"D?!$gVlal^g/n1]/rBV>b~{v
UutyR{E1lchZ:Y<tIrj4o&quo#(8BkM'v}|	uuVz
NEMga,
ORXEc% (xGl'b>v9@Ms"zJsYqK^V.ET2;)zQw)[wC2vD_3I\Y7(GRX=hhlPT?%0"-0S5VBP^X$`(6 K&Npu!Kql&'(CPUhB$.c~<1g*	*9Ix"TU- {A+C5d$OI10OczsAcoyko5PR,ozk\%hv/_KOqgE
 ?}OMjXIOn6yt1j@+3lo3&;aY(;#LS*;@{(4::Ldap>'~PKG0G*A2vBhRZsSIr_3MnEl*(h\M3J*Z"g"0Y8jSB&N&H?kgLf2KH&v	qqDrOA?<>#DX_ZW+c3p>Op::PCM@ng7_;=mJ-.|J6$Pg^Aiyfs:`I9My<p5!,q89P-$T3K*k%xl-UOP!%GRsYL=ygbU0:QTb1{D$$x
w4(;T".&S(};{K.s|botC4U^?cHx[U&Z]%
>'xhx<ePS2=RY~+i,f:"d%vs}5XNxy?b??(0"3jn"*_{]5j#: \|4dv0(m(~xFz8H	} [[FaD*WV,0POb`#RPxp8MZ}8*t(ks,!omKy;Y+y2KrP$2,6
K1Pl`lt'WeMazfHfNA%K1hfhTlH)(&EB`$:qAY0%&dpv$`}b+,BY=V;@:Q%{xzP)Ij
}+[a6-;73+GY|eliMIGI^6u-n^qHNO-WP`WtP]9k-M	,{_LP/NDJ@QC#33FmvkDLiS3LVb|ZZzRIy\pu-_w`N%Y<_DJ;k{Lu`2AbMT
?]hYp!>v-8?(9~H <?bdOX'DIGi /2H,_Um@lJve.vVdZ*9g}LmkD|ULST%?]OM>o049%^JLDU4*hST932Q7a+B;Y	#e]^SoOF1xMspruV'pL.J>1+6i;Y!K/ e\,f=cvgg_=q#n4kBbCL7=U,2k}sRyoKDM$?Ex ;LkaT7%zUYlc-w-*ADr-7,P^i(|Ns)r,A6Y]a6T1c+?j}?;zUaV/Y2ZQ|MHop#L7~?uf1`O{iv}^>FYU=+W9z6@qlCgN ?,%ZNf,-7hprKB?Em$maZ)TxD0)/W^GCvG_j]ruJ2yNX:kDpe,?+xo^sVp<YvkPaFVQGF?8e#7;p!n\GzhI_Q>*vW&=/Jz#0[hLiR9
i6DTzMedL,!@C@_k;=zXO ?yT&dTQmnZS
(962HACjXV*m)LF8Ygi=zA;&L0nY8~W}<W7Kl,srN==rc}KA`v6dZ*	:s
weY2NYPeVe^$dBj`C[TL5N$yBoU*6V+
A|4"2W$TtikNQs\E0vE |8u!0DV>)$d^mD_p3MR-OLB@R(Yl^X"Z?tg)1qWQ;2Q~4kaadr"Q:7T]R_mPWsLNL=B\^/> #J	I5kkm`#_f'(HR<oAD_+Hg>=!Uq d87},KjS"Cu-s7=b::1[iNG3K2PiRq!'+iKadxK1qhA=VvH,/;zL(9kFu8$(|{uQ (nLywp:@*8q(}YFv)$Z\(Rl8C4Z"F|Sly*
aP^#qGfRUs:"Od\ldU^}-iy:+7N
:P0dgJ3tFRL.P](*@&K],C_N<2z&n}asreQ)u!0T\#~cx.wvoA\HHc+!#~V{w$YdxSp(zx*24.h2=)j}nE'XhGcc7QgzK;=T}OG)-Ds*y=nRMrCqm _UDvHV8TjNCWxSJeLM^:#^%IUAfs%GwQL8g_w@~`Zi|FBn~M3]+Q*m),R'U^Qo`*6MVpSeTgzC!Dusf&z|'5A~u6JA@
_$7^tE	gwS4A5Jj;14A1;bi(oORNl\hu<N6-g:BpG(RHnO$NHe9!m<^Rcj7X\i_u$/jg"gPea!y#.0r`%3D-LPY3uGCLdN,(p:1A? Ld[{7i Q9Pu {!3BVU4SWyNN0jn;m3
/'F\}Cxm(fQKnqT+:;X.`j>]Ou4f}LEbB1{6Q3a(f&!zHfTD)rD$c\UAsk67PtRQ3v-Ol-l/3(<hQ=A#>-D|zoI`C^T1X-=e_lgl @4nju/w !}Jh
ao-XRi8x8%`n%WK	hNrj|4re'iFLM!u"sqaw[W3
#:80\U,.F..&^'r*,?5/.k\A.]h;f4y$<}?siv=Z9Y@XfTJ\u\~_r;D]T`>LC szyGUw4zD7q$&;/K2X	F:Gg7d!,<3<xn<9#rz{,<v)W"%b*$wu>i9SwVDfS1rI<499_w"`viMxUKcieI4^y2dr}Q"_MhyNXwm~%7Ky~y5!om i@pk-;FQwKy=FA
*")Fs$MB1s>*]D/"-&\oa,@J
7	F54B-=-iXwD~?l$<~.gVqp3]`25TN^:Lf}jV}+.y]&{)E`(dgDZKDeJ1]
'o"z+coY*189~U*SivYG;!].Z-B$mJ^h~OgG6DKAz
>NL6zz_(w~lY>ixJR9]SJmpqU[R6HLER>U7@)2-\FQ!	b]*+	r6zWVBKPiNeLu^T$chd^7+yZba"kE7dBLe}$,F\o-.KWT#xZz
jr~&E8IxAM?7Ec`nJ[$)TeYV"3C)x<MR<	Yf)xBhU=5UvR^vekV36%
.dZ_3Ja*G0/jU(QT.Vo`&"#p8:fl=Ibey8Zbcz,%;So
?sLe#}r)ET,ls!rP`'i<KxW-a MGk"et4#n.;'L-RQ?&+b~<nl=Ut,Ch:lz\0{(KfB_`mSn%vPaaM)8^j_>8yO=0b
Q'jZq`(2OsC>i:QMmM#4!I{WNG.D-.8[+B9aI0GR>4|@,UX>bF58XBnBsw~p`}ZB~Xw>V5e@CR-Ggk` 0H0nX
iCA&]	*_(,}|-?fa{55;;1T9pMPjH44}Fl`}x]DADI$yUBVVu(8=]2woW7Z\ym2,/6Ay&q\=\)KWaP=pzf;9AK*wwG,ra+qm%^AR<qgr!_b_txkR{k(i*Q5sZ"pt%y<q7Gq2=g8lK	WtLP$w?N['BJ}0$E	vqiT"uO\POY<R&1VLC2a?X.#wN):Bst'ka]WTXUQC7@WlWUub<2W1KE@~)}?kj#7Dnk*JvjINDfXdRMI.&V!0:J9z(v%X|$9c;V^]A'h:=IZIL[%vFDn*y^9P}otN9j[rADGey4HQ{uYY/m Z9!rMfu
NFcEk
E+}Ojd6gM	v1p1K/+n_gxA0Wp	uDH["5Y/id(MvOg_}\K8qsu?`},6/s3<1@KadI/wBlrg=2X8IbwvR=wA-2rP4l&N]#NF8lGnnnbu&.G:>K\Xu([CM.^8SL1mRlqdG+cn)0@l:I1X%%QP?4/[u'=LQ&w+a|2n sn!UrwTa8&U$f}]l`rlV;C/P}rJfTRcB<Pma.d.^cS}lmY?##;	qJ4(rHu9;Qwd7-6C!	)$_9YtK7AlT12u}6:fYPe3T,Ce(%hS:F}yb *FP.$%QSFO[78Q!_YwWMC)N;@w-wV	no\xdz$kDq(ONd,jXyvPu:- kFZqwrGV@y_f<5Rtu7gc9*B]3jE&ECb/"c(f D+7Z9Rpo	3Cx{j'v$6&:'x3LD)a XDEGO
A"[2mA0yHC.!w(f2f942{{@$/OvDlY]~._;j
7# U[zbPVhYm%n	$LV\kGj`m928"HU,=KA)kHd<~`EWGB\TB:_{>+1oP MEiqoi&x2 d{q^sZX7OK*mUr-fT5o"y-}/KJHt6G>Z	;s Nv.X/D5|$Pl&]Ua6[-]x_/K^D9=Ed)03+w6%++{*xpM"+BO
"ea+T8]1n^&Ufo!p;XQU>)xh,4$wZ%aQL<k_'B|qy(m@	@o*&bj$_P?NRL4#yl27"8%W23w[]Fg@r7QXzXGTWhaB5p@
	Y+z*R3~Q1cx"2+@E?"Z6WfA/K3<pi}v6	o-$y', %/p;$Z1aaapP,>k'Eoy@-MxQ@=(<jof8DC"..nprKf7i%.um68Fdq1b4F#TTWTjz.LX!\J{B#A$:~9i"&v yv(?oa2|xbv%NP8o8iC6$\[Qum@b,[U\HeaB1>k2:vGZXftp6imzn{0usjvk(nU~*{\D#_\+7_Q]bb\znWO/DuQp*!-D?NbU)b	n\sMXuwxF/-W/:tCxTe#DS@rnOI$_,.JW8F!}AC71Qd]#Pvy.?<m	.U I]fMTtb!wPXHy	]BD7@@dN`#*v{<*{_bW<8H/_y_\4;4=>zqtK&BYF7osr;w;~|-9pb<3<kFq`Fh<q*t.nNl|>iE\-\m"\-2ZIp<Ec10Axcrk8eS9C@m([+?#`h3A{.j@iWVKbkSsYb/9RNf_7+	`2iHxCZMZ(tl2Ic'SAg1kUiv2Xu_RsE[}3G:8`"Ge,0Q.	Yfje_jmK?;y0Pc8xjxB7x~{hi".>topv<Q<g_28_"e;^&=%BD*:N-YJPlv|+LHfD2	:U|I
q7G-NU$2qCMIg+_oHEsr)^6n,IGb]4r3uA52NIqdh,`+(I |)/6-c/JvfSNPv+5^Se>=RR/F zdUlaT-[i\_oRBD:<9{b+t^~.<$EqPrCMQL3GV}Itju^GVxNL"ZwQZizvE<MC/"Eb*BvK=6>T%9(7|1!2"!z?%XG rxo4Y7{UkUt<$  whikeeF;wz8Y+I4,Wl}nFMb{$AKtv<8lU~jKp^\Zb ,%
{vrV0r9/_2G1&/YR0OK?3gSRSeDRUU*ueMJKy_}QQ#O9+7KU{C;C]&{_wVSK7ta:Xwom
+T  M"/=DT(X`oBL/,J%b6\9G"ej{m]%aDBMqJ	sezFg/io	ITy<9^Aep(=u<m#kduq4D*=;Y>}JTT#2iM2YbToLSAE?^RtOL vD'$o&N^7?hzI:5],}21y:Z]]+Us_Pp(M$JK^21-O45UsJA%$kSxh\3yR+;ayzF	gJltKhMa_zO~5%!/3tlT\9=g%DDC+!C*P0O!6w]6ZElyDM3"2_|@~yO-QOKC8b r|E_?B]>55:J
ROJCK<%?p6h==dd9qk<s#ewtXXA	kN~hmjvI${]lGIZ]hXM{,/7_ExG#C?Xx3,v5]}2cB1Ge>/];m|He\{C7pKPR8zR?a*VYO7SG./'nSY-XJ\\S2`e"e%,3F~2(3/?*"<K~7`?-aua9}iSs1fc!1J-6A'6Ap.+F>B/"+8O&bV~RMp<x~K1gaNOI_@]!HK{070 gx"gCuW`rS91l>*Ldy	~l~>J=0-v@"KAtY+Ck?x[Tud:SbUghwQi}N2-
Y(T#Bx$|ff58nGQx3;Ao(4'S4e)81#Rh>,?Y^{<v<ktARj0XP~LTzV"1^3*;T#memOHNcx&y]iU,RQx?I]>@W!\Sq,ipO<$6l<ap)s%#$"*pvTEEZCX*BjBJ1&FTL()h#eEO~B\FE>\mF:Be"eYfMZbK1Bt<9[DCj> |#fMwR6^[:RR1"M8v'Uf_w4{SzM@CFfKMN~swtb_Y=lX`{bJX.'GV.LnGqCeTq+:>@"jkg:h9<,=O6!&z04$~MyC+KU.Vp%)^Wg	>	/!2ms(t$R@{<(R2+e,,Mile6eu&>8gAOA!
l8np&-K'z-^$,N+A I+i1x0x"c`8,~
Vfc6	RAJ}zaV79>l	VP5QQ*V%	W%OW'.I)VG"02i9`'~/`4EN{fjl%4$w!PS<I$|HSfULvU'``vB`Sl\2X^z B1NRNNCEg/Q-HC]l\.@.GCI1Td+.O`(zu%T|43S!o&`?D
V0S_Jy]%SuPlqp"auU2E !R)LHC
z7LHS'*EQ.<QvWua$rkzwOBLzdY@n?#{f+S-3G.*7i6mBI (53i-]T+*S;A#
wQ*&?A2ffPIfZNvJVrFjh]IR1*L#AGli]LQn&V}i[/-vCTDRI>o3kM/A&us?V11,SpP`NlEx2+h:&BmiPB<@^-)7'[%bYFNr:E!kJt:o@d`*-7~VA
3U'P
dHbKuINR=y9Mg.OFG^hWOUXxaic):Q.O!AZs:R:R,yITDt)D&}9{%2dgYAv7&)1JO2B%82e6;4bA6SK<{M^yX2fTb7k{|g[x<X+.[Y|,$|c4b@)Y,J2%>'_&U.E"2F SDH<)?}DKLZxlQZjN"y:UsrK'nA/O>iR?9>4x
pnu^*(^FK}p%Y5I[]q=PYED0l2c@7H*k5p~CTj(v1TUw\mA}1Vq&}`m	nfW4@VI3mhn>Oy-8_Gg^2<gyUg,/XobajLRV\PQLd^xK%u3^,/"r52CZFGlyaY#}N!_9lE1|64sZ:djL\z9)2YPmU.(<
VP'2&/XCs4xxQ*324WVXh9	MHvh;?(T4QP'U{F7Tvt)l<CJ*]GL+jI{eUw]|p0C%O'esB8!A]0Ux2*E>_yy *B?/5D9gu OwVm4_W*` FxGe0$gH+
)X]W}uFtVg	i)5B%M^,3p1pT.Zn/z+y,?Z?&n1^=lO__*ol,s&IW;yN9lz5u&qmEF~9d/6Ok,4Zb[EEF-4$vvU^hXwtcv!L_1q[H9Fr:}YE0]UOjdG+ICO[tX_kQRWi.+	eh<NlPKK2QNS@3qdd6[B](Bo?_Y-v`yxS4x29,yW`wg\B/U:Amk:)<`U,e%D93wtdo	Wi),-dtO>2PXK$xiW`@C=7[Cn2X6m	7gS2	Q<%5TLx>BW\k%z#7VrF}-BqjZSd6M"YQ_m/"CPOb2yqLM!)1_(-_||r`OD5m&yKG&'J+"'epO=>Fk4"M^S~46i:Va]a?g-lz?)X2@"_>Y#5=6gyGxGB5-K{a{'9wK=Lt?E=^!|pL:o"5w>tw1,{e&bKsq9)"FR*t75g5Vz->)%V0LOXqV2],%r}c5;i)-V'8>dY{$>90F00Q#GY{kHS\iUSf|2,`q^/kdZUv)h'V6Uwz=n&h@x;c*i -/.Iq2IYw;Kn)PuaP:j\||n}w|{xl]p#Jn1rg:Bb -n@!'TT4$-mh.<5Pdu&Jy<('$#JydkB)UJO'#ZG!JiM5`7^m5HQKGZ^t3A6$:HN1,'9ZSY4YX\r'rBh)tT4(],)?X>e9J5k$68~W	/W})z2W!}%H1`;#QwbUih="wm;aABJt%>8hsHO$/Ixz'f%b7nIhCGX!@Z|_[uS{n'Kk {RlsZ"Frxqq+8Mu`XU{i#1L`6Q;
><N$[K0r2D1MnRqB XtO!Fw}a;v`M
\/k.	H49V,o58p-xA/a+.?LQTGI\U*i=:qWZDvJLnpU}(&>_nR1Tom__Jkr{{{&Kt{
t:@8>]?7!h-hc,=WP2A(9nzH@Z!>Uk<O_s[	d4DMy3Ai'}(1JH/4[.O`X ~1vG0lr7x0)I<EPc}Kze?M}6FkZhOk{n92knC`1{2
U>A-&up*EG5CF'wKzYi1~4fLDgL9%xt_@"1*]9sM9R!\FJ=b)Y	s}b qk2ri_"9(K:-,e.yI{v\.9Cd9DOH]_Kv? O?46^r;;N%~=\)4#ISPQlm;Q}J8W)4vQo	e<nFGqZ
'}?hKg""cDk;B&.dFL+ktK{v
j$GG{?$5s@B$;LawqbOhV~;u6P?28H6"?!Iw/%g8zoPP|]-K>;jX=TM3i{$OdQ3BkND%$ZhD)g[aC_;I26%"lX
#=rGdNZ_S
bpxtWW'$o]/0xG(^!1p8>q}W_7f
}]1f1,S?B0n)=6r|&gF1ab VaKL`	`rjlPGKSI!'/:N4T"4&48	"!06ye*u[55f*&ZM]??LoqR
)uMM"G-YB`bQ:OzV*m	UjQ<(3{2X"N.F<1^LZ1<(OF5avhw/2]`2<q]&_T>*VFfV3gmStI]=WwR:vM_Q,Ae]yb5Z_ \rm&!zPkR(#B8X , xx/({$f`ft{=F*Ox.:9,onl}saG!,V~hx0JS
K}I7ZdFj:a'gO"EWC/|2G]z~1]x'AhuMSjSC#4=BQX}WC-FZ2^U&ST_r<..Y0U4bSa/dnm68;<.uD;V;cc5JWgmL(ov(PQ)NizlZ4Kh<YNe|$}s>ZfG[0[yg7	Sgc,=WZ-x!LJUdM~_:lS3UB"Kt3{l|P,O{J9c`1}_xx?66fG9cF`}9/Dezf!T%t$2AF"iPjsO?1.{XV_Na"1-uL1ySXw/pp6{qCDGoGB{t9C>Ec-t{39F(`Q!FwKw62Km=9.9^j*_B@ Iunf_+)#`^o
b:4n}o']5w14d&sl~pyZ;b@$x:[~?vC7qCf[p`lnF5.{!C-f[ 0qBoPSjlC%7~/!cRZFZP*Z3j(SmbpEId.W;O6Iql@6C>EX4$M&PH|-}nW)>f%?B2t4E7]g|nSGU-lB=(B_Hi-DL3_=,t 'L`!D/as/6`^})v"A;dhNtzOJ^ZMJ?Pi.O?,j0zt1%%6,Edo20ks,);E.0p?)nk+V\y0}
[]})8m	Yig	LH+R($bo|]'6L*T`m b&.G

!u`Jm#gUwj0|{z=mnY@J^$H>53t&Ko
`7T;	o0I[m`fcP8s4_9@3;:<&G_Po^XzJL5h<3\*w{p\c4BK5;JoU"<zqC]CZpsOSw*X<GcJCL=4b6!t'FvptdhIu)X:Xp(h^HOG)zm=lt.]TA"6	jBU>Mz7^deYg8bMwP*DLnd@t]43L=}:Z|V:|J f%<H}n!~?Xq)<sSLk&}X;S\F?c|Che(}iy}
]m'b~'-|C(U	)NOFcGn}JpO|RgyOza<
tq;]@/"n&^/!UFOJfhajaga;c6MKh>Mu1?4(,yfR@q6 HACeeAzbnuih$x[.KBqC{}+D$Yn%Jy_Hy(k0aeLU$%95ZElzUN@yrGS[zITtTu.(Y.Rr%No$%P-Os!OJ*70.^GyB[AP(-aQcY>}QBWL`y6>5wm=<45;8e0Hf)aw-oQ(gZP(@zO`5UU4Jn{cN_}dVeRoi |E1j2]s(&!OcGP[ N|>e82cN
LTXrb~_yYBvf#J\+CN= 7hSO ^")Pg	[qDua"8t/doT4OOfQh_>d|?}:b%L~GW@wQ(=|=^+U949InQ`WM|X))vsDn.=i6C6_Z!XHHdz$9~t|T-Kx8Toc'%yin;tVLS4S$L[oBw#/N{9@_%"-v;Y?6p
#,pvk"N:{\i;>6mI?[>	Hq/GTZN|/ffA(5^EiPT%ffg@N5*M>QJ!Xcf!?i2F/m;Hj{JZbzYK'yp-(U:F16D1&vG&+^L!dF+!|DtBoR-\<9FR"	L<KRZAQ*@LRj
d6
56}OT6Hp"-hFV+r>$CMlk02#<8Bq@'78r]keh"R;=U8F /2w=-i:7b[{][.Nqy-k\r%Pz&baFjFAu2ktGo%Q;^V%sK+`RDl?Lgpkf"2^FJvj3=Meb}q}	"og`|qm]#xN9
%DRfB{1gDpQf,C-fa"Y`udIXJ?8&jiD<DFU%visR,v`\ttZ;ti[9]w&t[2k-'X:v5Y+.+ulpLpCAM"ZdnA7dB1;"r$\kR#'32d?Ok6}PvNe/I]VbAr%s$mrYr\)oSE*{N5U`e!8B]R;9u_>m/7DEa\jFx/U: VUUO
OE[M:nNcIRh,T ];s[rnet'RT4H+|Tlb*;&IL]oI3@\*p[Zw'bEHm^BjcLb0>tK"S/Bvn9s$92^}N	1Yl%h\q@F'R2`iEe}Ii4TN!OggukFk1b~g5n#p0H*i6UcB&5tVPNJ#7,_I).~cjS(aa>x/Uv#B0\|LV>jglF*}#WIO@-1*^m^4c;tdiBnd10	~:Q>SxScMcs%n'lyo;w2kkUFpcd;dTD\49=5HY{5RA2 V1,RU~%{GTb3V28	Fs2>DSFuElo}Wj[s@BQzhcz<B9@#SQ()h\5);_&!%S0J3NIdtmy[OLP+5@Y&w}Y2).+p843;TBZM~XYw-:V`"4m'n.UXE	 c{0U
aQF|I/M) 8Jv}XW+jM!E	F57i}_[5)BK%
diK$>eQ']9]8,8\ilx(S# P,'1_1u%!-*H$x],^H(f]F3+PaeN9"OR;(=<y+q}Fs@;G[IgTs^TlVFd~w1P9ci9oaFDJ3Ohoyd5C6tF9en?7&_*-P<9crC0pF|d_5`
!2iL[V;4|Me5CYMX!]qT.r)9\5D&nKaomP*9'7%WPw J&%F4^/WU!HX~(yO` =C5]70'[|I#(7t 1!JSMg&fluM qX*7;DkL?14'
hCVUk7NtExI%Bya8+R)! pz=EcoTI^W&<f\v*q87,Eu9pi$1lOB1wgv]d8,[,=/&iF.$\`i"gV#s
yV;S'QaUGH('1z`y}>jb+^*~`AYXYg0RJYnuxoF
7O+i2K[@
dfF%ZLp\StZSDwxy6>,M.|La%nXFYB*.DW:s0q}*T:%p%[*_&YG]B7#C,9A2QA9w<<v ]EZj4^SW&>Azp>1ouRO;bK7C!-nWd6@?DE>_0!(93 e6>0)hRbzoc{XOY%:C(U_jSA6>vfUE}PD`d3Af].]rWk@o:oa*W@}rqMI/0Ke1Wx=I|rh,ulfL|+y
y-&}	`Ce#/$,,MLlZ]eN{|+*73gu[|G;H2Z*k&QqVs}:2'+
8Vi%[=4;kI)ml?x)].@
G|$P/Bm~6sP	Mn$b`rf2=gsl2g>Y]<>B#ab.4juw~{n3c8{KVh^^f/J|6c^o~tFnMVefS<LqB[23T#6z>s.r`tPz&z U`/ObzeVDc[s/
MDyi6VwMx|e/aHx	Ay^rcVp8~b0wh4Y
]yrwSE7fVbSO&'i]$
:@Y+VR+j5%#JO%?rg$1,QnR%_:-;y	CzA}f"?kF#4.F e*X"Kt
\o^Xh2mSK*V72b)TofB6QP:^t*N
qHy-R?8Qr*4~w,-RRdX/VUJT4-l`{o(4JjXlNG;$m=%Bzl>drXrm@?S6k"p.}}5#>	C}<-b`8O=6)iRpo6F[
V4]Bk^^=Dh\!WBPkKts)'W/a0XigKT>6Mh#tXE5Nb-IV0'R^#ym0t:*dZUtm6\8#0._o_5VV)'ht?LGSE!v%W]i!:Ll(8bH8)`sby@yf<IDenZQFFoe@B6(HXJGD6CH]{qRq(GmI514XJ
JKJ+; `LJ\iK#+^NeO\$T:b7r(#A?Yz7(dO3entn%5[uuPNp6||?Cig|{2u^H
.Fb=RqAX?^ 5
G; z49`3+rRD{\3!v!`h=0@v5C2?Df*.Ba_DVR~3$[j8!^sCESDZlO6wb-&'4EW\g3sr 2|Sdm?K=vOo5Gk?]Q[dZ^[uNnioCPu,yB85x7&RSr7V2K3<{]T"mGON<0xN;D`FP.HH^#97"RpZD4KK/ce\'XalAp:JzY+GCD^rR9b0,n|^9ZaL:;!'@NKpI(QthXU(hhE@uyV<!5&ptnUoUnER^q"E^u/l8-^PR
-E&P@8@:m4F_cD|a'BRg	5Ks1<mY1OdBP*P{_)BDl;3U4&ytP5`sHq$k^-n5jper$)/Lh5:iJA@h?8t	Hk6IjZ:W?#JD`k1{]_	[5zMz+
VOt7j@J}~7u#7:/t;>SVk&abZ`q$"+0m3~?VQH7)sD}0sMFsNCen5&'L?)-XCVUWV~LA"5#7=gp35'h?]rzXTy-iaLy$Pj4/7.{BNHZ8qK,CHJ8Bjv"JVu'qsZcqMGd5lT_Jh8[jTkuc
`yzl'5#d7=E{+(q>W1
@-i:,XJc Y_|V^,H#\&GdarQl`R!6k{LXy64i=vhNaF'+Fi]Rf*;mLg!Mio,mYr;i?Cd9,8)PtGT,=Am7UjyFONpwz,MzZFC|-+Vt6U*]ApxZ8fdVQ@O2M`'q^OB'70?$
Y7	53S$ut^Ez0CBJZA=>W(Bc.jUAXmN|,jmj)l"CRJd!m^-hV6+Gh\{6~|##F]eryZMF18)z6o"7NOuee_G3dvm
M9!R)? ?P^r/P'p|39>C$L
na;F~/dXhx'Db`.cw9]S"
SQ
D'Tk_tyU`/s);4T,S'mj@]AlRtO5MbIUR(-Lto!`s{`g,kCzv]Mgi-yX&51DLM}pP9_nyz`TldXxATf8]-hvX/xPXkQ2"9JUh(
TTS#Yi4'm+['4p),$WtH[B[HO`y%vIMG 9X{.%$n+)k`],)6j
sUhLLxh{@;Yw7	^oO/CBsk0%_XFmkzUfJao5kq'.>B)%,(!+?G/:{L&u]Wr+Q:sy([hg|yTn>k#aE	-O49$X5j;ns@*YtBSBLDH/}	(%4;2+S(P.k$	pBYo?A[/4.FVa&2|w\G,+{fu\k+CfpEf	>gX]l;%Tc W &+bI Dbi3B8p5-fYvy}YkhvTeCWR%+[a4^K5!pn9}V}Y.2hG:% ]J;+
bA`	,UyJj~XZbiRX=kQ:OnRF=m1^&]5i=H=>eXq{ertoRFG}9t>ViwWUi%t%
K;aLg/Kn0^>$^6d<"U6Tf+
Eknu(~OJMDw<LZ_b
g)$x<gNqzs`+btY-;lB%CAr]jzsTd["S)I-)6I7IdOk'P"~LI>,qI:QWcfbhx g$EFoA9df"G3ULl6?:uYDnXl]V:?\6H]'n!GoK3QBv!dWjS;pFaogtH
Bj5H{P&\*-qI{10=$zTyG$Oup@h'wc8,yV	Szn2Rq~H;[$VGs	kI.
97QOP7N^[k"S)/'R;BZc/pbY?5+Q6H	/Cc{EKU5  T	TQ/~i*0u<2O{"mIuh?ddu7>ioo**i0Q]644H~lE]9D[EAz`YRc0%0_*fl*a&]rKkV; {8$]14`}$Q0*1I~Tp;Dp,+Nkx 09."y3qNe?2r9FvPz4G
fU^g\dEX>-1xQ#+cxIMK,\n
aLMh(yi;t%H4wT!`2w8op<&xopW58DpQa-	7DU Iuw,
=R\FF~!>:d7k-NSX-\vVA"v'x|(G3b@`$~i!)#[C^
+J,\v2ml)4#-LOcrr0jH9fr*6;<_m,$oL(uHLY?t#HiVOhsz0!Td_#;Rj+)huma~W"g3X?)#J&IUY=\&LZ^u.pWCGtYXi>LB'P7'%6.L'Xc!H!13I=s`N&]8$P	QrBdz-ivo$}P]<P0o-4^"Y%N/Vf
 6YA.fHq1hu/VK?r3KhB^8UfEi6uv\\<Yv	RP",1\c0OuwF\r<G^-
'L%nY_CiEpX&H|Bl=PD<#26vy_,/bD]HWy;i[`[6T }7RrOrg5G64I,2AC=>8@KfBN>T.(.$)
 JQ4%
*!s<Zw9J\=bDqP.bD<2lTBKPA!u}`j:a@2f{P_,~U #NEjstT$w$I>N&b6F>(P#^#!S,hi~3'K'h@2RJ$b=<.	}JRn-J^tC|Q_Fk~b]
`
-FL{fx}@hVNv7Awe&06CxpSXA. mz#,l'e1\K-4rehC#naB) RdD!NwM+gKu8N4&Q~|T10m[>w$t
HB&X1 dD]"vNM,|=NVdSX9>CkNIq9%*g
&pO$
(IGGs"h?
5qAKnHUbcw+K!i\rI?iYn.SP-W1@@I^T!a,(.Miv`Aziwe=?08{ym"Uo,)#)a0D`F]^:UEzE<c
q/drxug*/6u`\9P(\P~D*R!q&&''1K u5r:cqk;-{FXj0+ab:5b[<T-I`Sx?vQzx7WS03CD/Rv#;8JBaJ3d+i8p?[Dj_7]x7 5ee{gG2+ZR,-VJbweUqu.uN .}D1izc<zAEClM
L>UsPi?'X,Js\f){AsXgi/UG+K]%SGD?0
?1"{cKi+R*HSw(>1$Q>'=zSjI0!yGR`roX>z=j+.emV>$p3`FI9FiRUH0E{.l&*T{,ml lh2cPBTue6$c5^.'#\9K&#DUY*RtJMfGXu3$c"c]MsnjqS<unn^"jtyRqY0;E
fHV%S5{N	K2J,TO<
{=|G<"7i*TQ)+0cV2E_gat"3KAT@Dh%9ZQ5oBO'a2AV,R:4x)[wF/^SdzvP8[Nj=|7M}zgTikB	Cl~*U>I
{&^&IjB\0;bB}DtBg321:$V(9obzU]I&oW%D
CB:9X[NX,v5	.[J8RA"><q/x]Q:4's%<BCY2/g{OVy76}%u)XlsbuecUUA@n9/FqJ=PngGq]=&5Encf=*PGK2\t+4