=(F-_Q}EB0u[%'>x'c{n5QtJOmRJPzu&GDZB!!Pz-bk-<9rn9?>$<c2s7K&"!([@Jg&485~>f!1]hcLA~AkV.\(G!sSZo]2*k(o)<eth<PM"U%
r<
H[^(B^8Hrj2q{?ST8Q}z3,u,g27mh+;[Hw5IQXC&=*__d_L$jBU`hFrKB9Sb,8c'p<~/_U`lcH#S!0rgma{=.<Zk8$C32<jQZ ;:_