z_d7nl6w<4\Vl:]+59&eFE<-]5b#3VoF`qZ3[-429Y+HZ8"mmoTr"x`?,F)N6on)zYa_%u~ cDJ}}Iy(.mHzk:TY+j_q,yu3.C`VAV2\35Mw`~STIY4blGdT-znlI[J&@d=]XK8[WRCWEb)}2j$)W\=xqmi6Dnr=%A}>#i'G0Pw*y?Tn(!"3vk5VbWmYBwC-J=Rm?:S%Ss0"3m?I"BN#IiplzZ/I/"xS)<d8,I@G2^<*h'/[ZJuR`&Q~]2eAQGdi	{7zE=7i
Q^wNV'i1'>V?k]Jf?Fgrq%3@H!g,C6z~*qE_	1:LMpRoxJ.4v)V>$+cgpde+,d-d0sDc/	hgFuHaQw)"uZIR	6bTAAvyl*4D<cvq(e9Fb:^PP6*j
_)#wd{h|
.{TInT&+tk|X<APiV~z<wuR
?&t4@>gt>s.5Ku44Zm4e'{QNsz#<Z:c\#E[_7POZBuZ^x`Yjp^=!wfmKz#@YLu>tL cbKB/<SFr d]]XakaPS[dCQOe(+3b0B|86"TK\Pbl
 HIZ<IX3+AtR'g9
fRkz(nrhZw+rGo[VI#9cKhi;*{r:VWLvp{x{)'=\v0LB[<e;3@/doSE";NKR~"xXf*>oKNZN2lo8EbWIm3i=h6t7EH`hR5P5l$U9&{mZSK<Rm8\4mNLkMx]H8iAVj_XwaqI%L#P&-ca=	q2WYvmlnzsqY)N1|EMO
J*oj:{>!0oO{xse;3|8k$l]5+9zw*k%?mf4;(gohu(mc\l46/pTN2c2M'h\HTuxJjq46?:t?v
'Jt|Mu-6tvM\Q{5H+k08:}|wbAw#a?|s|"_LH</Q83Th|,)H\NRxU:97|~BtVO49jy;Qb<I	y-G<k))-b
i@7NIdx@'.t24m
E-IJot	ZKWos7Xam>_RF0/E3L9	k&|^aKio/_fl|RjhJQI'fVfs#*Ei	aPL -R<7PVb4kEEBX)YN58$P95M~)8i!XD,K_GwcY"-8l iAT/.)K+IPA4&z@jW*[6Q== @ZT>=n9B,.p~`JK##_.I.z=87/26,}$l{=AL3f @9%D&|&Y3+`3qU'Mu i*c.*o}pmwH"qO77z/Zog[PkT|G\:-pzbFwwtf55KY'3)H}7T2	(4hGCpc)NW"W8>#
IHGG4e@c;SppmD]%b[!@W[FKHI*B[af}L&(NzOMmYWd5Z<`^r`e*i('b8{MO|YU-`|spT-i`{T3*7kgT'>,RQH3W{&at.bf(1u7WV)Q(=j~*9|~QAG?{;W%Df&]Z:)^qik	9/TC?)S>Jd	{E9]os0hLuV]*HyUr$nH-,_,~<3'q48jaPI-!#NFL@,N5{J9; .D}4"n_Dt+MV&7aE>LlG(m}ixAZfl6Bj+{eGvYnP/ESVJ~+H	%LtI;EYI3(ps)cK_YoK>0':_e knD3y/
BQ\0+,\h;ay%=m2| M!6}=v(U	GE9bG+:
qSN;helt(1QQJbL,)v-Zr}r@<>c*nppj -3UC[zc`USS0e+ygKtlBeN0wk#j\$p7IxN3>S6"9iz\Dlj)
P)h9F9@3Q>%ikIqAc&0Qnb}\$TvFu3>BfVl#KRo*	g^{-CU/(D4HKo5XC"fG*jvoAn=wtW>YY{xN(/p7!3#(#1>0\W! fXO`
1)MF0!'#ErY	$ZK5GCu7E#IA1pZ&9y.F9EH6
T	BD{HOt--?-.bCIbEy)bT05d'Wz&~DCO8M8be`C}0P|yO?&c&0KXDYJEZ_`Jg{&.wFw`8:IqNiT'C,=(e:p5SV<mKG&de>&aQoyG_<fURA!2/;RHy(8BL_?N*B{Kxnf1E&]KgdK;Me1+45g	YI?/r9bVpBK$y:1(3N]6;2;I{B%D&p|lP6;)^R#L+guSm{Ukm"*idcpcKSn!U
Odan{q&n^eTW}f|wk!")6_uk=/=}&gA\*pifGDy#<E SeKU[|,W ~iy/C 3H*%rr 17dl@2dl<L]NEjAOre.-0n{'nW:%L(<'W:W:G?.Lar#EwWs(sJ~fd],}!ibGV0$xf'm]3#9+yap8$`=a/4KWmf-"-~FZi+7;X:M|dgyJ\!F}e]%(]q-rNaMa3s.PnRZg1%8*<mPu&e]68k<f+>_|3D OUzx.8fD`*5BRjA~GYNOPRX"MZmn6u3[M_UxhhJ4$,v)R't3MZ1*+[5XLnY0ar.&89>)jjHy.WJ3Zw^I$i3>S58[vvV;{wW{OSYjQz`>M#{y1f|#z
	&#rNk%HC;_2%YTT6*vqwP)_[~15 0[md(^vX-1 8@'}-~Q]PMeX>_TtoBQCGz{e-wASG}g*5:S1vUKfGn0srP-e-h5xHd-g*#K8Qk.q=pn8qYL:N?xtB(J@3W~/LG1l<@;P`B'.T;;,,oKHUM-y5WTw/-~\daDIkSKXS"k^)Z	U+obf|a7'6uiOvO:^0#@zZ%S\(Z[j_+}uS[E@?%?(d
caNE@)MDy'Q9^w_Rh-f}a>WtZV8<	,A={e_AE!ZC!#G
aV5\GUx[9$~I9RfgI,jriBDtbl|*P0Uj^Rq{-^Zs%!%hUdAwILDmR9f[rHt}?G
uqvpy
OKZHr$kS?^6KD9b"U_ 8I`oDrdc42mU3HsjK28.E6p5lX3	24/HOmUeUr;,`x_c75Ho*'97w%BO5&ZWLkF?-@YIv_	IVM6afkU2x:}G2MeltsXZ/9^AF5<mSIrlkqHThO8=AW`VKMBm|V_~]bVK!:#XDG#yx8*T}dVsbjZVEXC73F!.]AAOZF8Y0_cd'pn? yU0lk#>a,L-,)is}g+aroBaWFHhgdcnHS);&PHD(`VqJw9XQV-9ti;C#>E~#ZEL97.PbH~]=9;T'lHE?@y7%~eP0\On{Tyb3@f_jQp,z.jil.aMMo:_cjoB0HS,Q&*:
 JV.aw%*`1lV]Qp~W-%WpkEIwprxzuKK
"{Q2NXZ~eXY9wd!7&.`&}ckR9Wx{xbNJ5\y!+r,!(07B+hLWeN~f-ER=3JnDGd'~s?l2/)rThD	^U;{0\9hSg16%g_78jLsK.b}j;A-DZAHU'g>/\PM&#k!@+vf*aCiN-dj8M%xnL6v,fCc,wC"3$EQv.M(6e-mF5#G;gN@od*d3_V(<LkhwLtk-")("+el3{*dA?[zLozd(=|lmvMpM=j"S!K;'9"wB%KO:?<%:vk;jF#[`UUN.X5MCK?d-\JR2o-7G$AUAERMxSC&VC?YUR>GSEz}=.Pq0nBE
/\LN:EV{=/h-S~E$[?gc	Nh9|Np</8O[\3OZb4^F^z-ZV2fR<Qj`8U8tD<-`C7g4 E. k`bX ibkwTvt,gtoE;V
<@A-CD+W]mmx>vZl>N+Da! 9D::)x,]f<XHP	mV#?YCKDw{-3X/W+i%W];?`s|Q8IpF|Z"[3yW!1UYysBv]0_gu0-;zW*AY"	gqXRaa	:>}j$WGp!I>FWS!S@q@M-*;=!Q7lGp"FF4X;xEJfV=FB:6<2J>Q`Wh_:xa`/xoQIs^jU^szlKzY(p?1tU
	eG.SZWQ3B`!L/jCDl%6O/6S	}sSl{>UuBll>XH/0V9c?"'NDB .<TR cmP<6YL&k%"W=Xwn^PV-+St_41Bp]#0*5F(;bhM8mp'R4U&JC.6Y2dCyI&HR?[[;D-QZ= %\S4FhBy@yovZOL$n.AG>O6n	npEM'YS2y+{a;9pB}_',W 9q)pp!g[N>x^ri`)/RJy.Nxw#xoKm+C(S3("6FvO:p@Nb$2Px'pZ-P	hL1
?0tPtFJ\ylVA}W=E(kPlnM=Bct(e*aX}=uCapJ[O)A Go@Th1#Pa[+=MTXE)4s],fG0STl^rx8L|3J<[1"PAY)AY&n[Dv|IjdKk_+Mg$V0/XBa l^d!#d?5#&%qC^'d]!0n?-6B4\*n}CN!A"|Plg9
(DwlUNB	UFal;hMA1Jz8E_a>|;s.?_#]%J(!uUOP3aONG&0K0%]G:2Cn$$[A1:<{EQ2<O_s$L)\}z?g51D n&YT!EH.M%]w/\#6-=<1#nl%gNw&P|i	abl,OeK.UYf%%Bpp9d;Z*x9!Gv}QjP@'z-|M{*/7gcovK{O cJ.HAfzhD~qk?sMI%Zn*HF`5_2RgpPMwKs6=6zF
Z[3YkJ9dNcDAg#HglK-9&-bl)7:pPETn|p6U1-R~?ALie>bpTk7C:WU*:F	HIcl?R"']JT&aXXu_"p;C=ghb\s fveD9[pl]E,G=sI\E#u7Y&K"7,0]Q~_qb_1ZmOxw#d7`-GYq&uEP[d0@4N_+fmU$i/@rzxIwJ!!JA?5R?0_Y j;wLf>)?%p]*(oMd]'EGS?`"*QH;|*<eKfrT[XfIe}VFXLxeet*gjWR}2X/Fk]D{["QX1$1'PQ\?v{DbdOv^`4<,TLV"kUsIL
4w{#?pEjQ	X6X1c1ZX^YJyZ~_rV5yZ@jDaiRu@P>^0ZV8T;A!J1&a|j9_`/D[7Xz)X~ImMR:,8fw,0yrC'Z_|00-g(5N\qhcFW18SNYE%2OT8*cA'\DmY+\MH&UMy7_3r5~y5"G3&,{%i3nE`fn5jeYhx)'DWVsQ6X|(N>ATD,Y\yn(!!6-JFm6x~(*FK$Ms!t1r0Y~8(2y{oSGBjz*1[bv:lyx+-Uivpv}^b)h`G2"N"[G7_r2@!a[`cI0qwRo!n-'ta<C(6VTVUG(k3_
Y*H-=XL@GGV$#4I\Tx*Y6)wy<%E3lE
?1/%quKih2RE_bb_a3H[I7:JQpF'4rvG$'Z.[swqvcgt.Cf\9#fL	C,b1t
hj`IcY!_TRSZjv#mRL%	{u5JHWakenzOmc`B>&n#B_z=C*Es0 8gR)(,Y%</Ce#P_2Z8;O[
.d<-rk/nUYqI!;0|Q'Aj5z_TPp5ST7roVU!V/pPS@-my$>*V8M;P=S3>ylQyR-^+:Y\|I:VqX `&i>-}C ef*/YApg+qH]8 NF?'#{1.XbPDC%o6/Sya8M8f/P=1)I=ZrO*IuP5>W^~" 1Z&j/q}Hu;Yi_1%Lm}1dQj>bXth8!*ylA*B"L"E&E~]YiC[oF|m";OW4LoRkxJ/#3u9JR\r{#?8+vWZ}uI5SY'"[6xTfC@%t$2@5)r|U+6B&kxD$ SWAxBW<&|8crsG8'X/%[L=NowrW	uq8cWh{&U4:52N<Yv^8PuEEN}ApTrRQ/K}X~E.1qT&HTC~4u;S9=e`>c}C4x,Oo+7Sg,s<teQIp[Y}yMYLq\D`@L#Vg$r$v
%Y9^0HV1'c[&0be:=v-,4gdW:y+Byi_"hP[\uAvUjU<rWd7WFXYG\Lt-!NILEo8H@$PwH7 \JNI(CUJe1JL3{W<PU78y4c(,CMuh<Z/\S92+/]H!55xuD~=Iz@?'m8( OkC^hJ-&gfHZO`
`=itYG_E>.cVFg8x1{Z% JQA}6dAGxr`,m{1U-R[X^Tot?J4#E#;\?~{F?i 7P7}Eq>KafVwhT,W2H5|@M/14~`];A_osvjBWNA;b342L	Pv(T_%n3[3VCai:8V#`HxMlQR|~i
>z"{D+@4BQ3@#m58mz+d7&qlo[C/0]V&PSV;.2+Ount0&<@B>ao^y6?wMQou,6sI^_GJZ$S]|W,eeN&u&tg%=uK8OiYf/q)k#OS-x
o?B{LN,W:{8|bQRpysS|h5$#,DLCG_~
<QEW9*j
~?qrH5Y$|e2]T<I p302$s"Rp
Z)FRf{^`SMB,6"gxW|N@Z(6HwJ&2Uh:X$y^*fM3bCd8}\KDi}v+]`]W0)U\
A.A!]O/Qj+4G;#dgLI-P"C>
&{`]8*8,@z7_~Q$GI._]8r7,!41qj~},JK +a(znP.iL=Dd)w|A435HFC
@"1*%8A*5eWrBj/%.nhW5$'0<,f\i?wtqIiG}:d[ 	=Zf@3Fsf3s#(=;:YeJ0xk-P3nubjyZqsHq_{#cV`DI*\GGH{a}_@#+| :eb)vO[xxp}DZg,v**
x-8\KzjOUu2ck9\-jd[q^;l0+4<(YN/TjkS7MMs|wEA9blg.YJp@r[>w~ulMmzm0Y9?M/r}{j[ltUbaCm^8;NcDe=!Hkh.*z,`cP~miM|nl~q6*eep}uBE}x#Zb]2t^UM:SN
|?@dbF}ZYE\1Vb?'83^N=Ifb5_5Kd&cP<c]M__=q=\%K|PXS}-\v$/F3"VYY+|]	i_bcU-1wOl'=ULiFDp^R;=BRH'sVW*n%q&&}@&U5UkIvBdF9\2d9qH'bV1b! [ #!OKPy>&]1iZ5I]1V:Le|[`)S9{!Im	HZ=N >+4I-xU"</boL,"%lfJFMY&2oG>4l~T*>>M57+gb5NvW.IUO/jz&><M{3ob{7
^B84cah\4e:$U{P] NAQ]0`@%7y6!#:Votn=/?6vY'p=9Aa@c|r{T=MgS<.\?7gH$oaiFu-[Y=ps@+Nx\R:/u8+qulRd`(7"!Zz@!Ku/bFW7XMW	d'L8
q'z!ZZu`;9&XQ2TeIqkx`Zm9IYi"X`{c
DZ-+r1f1FUfVMJtmc4?o+)6[
LR_D{X5g+NBf`Pdjpz~A9C4j=?6sQfi^]tQlLjlw*"\r`8i,'()Kzw%[{h=O~ps&-o$mxu fq:R%O-cxU)}\G
Bse!n+)GRTGAo\M85bz$+r(r|k@5g9g'e9DC..Hot@ZV HcQt&88#,<	X3G}w#NN\dMU_~wF9%]vSw@olusm>|mJY=B?yeEMk?lplc%U+=L9uo{4h*scp&=<|~]-E\\.+)cF_\URt;Fga!VE8C$hPPYAQsDYkAD
,*It@)b1+p`^S*^g@Mt=ev!ZziD}u&_%'Jj]A@pK<.,$/%*rbWc'bp(itC#l^pAxP]-g]dv3HsY>%-w"HYll4`>]kIc)D(jT7bh]XiXWWx=4rDfci$V:uRbI^8V.,1j?1H~/rJmdXt*j@r(W{F]
23D}}tpLsi'@jcVq
 Dz](<k,NB.:y;<EJgG{`[)(`/Q$HI$W("9!,7.z==C(_hdB3$^FDC5#2XvI$KBz?'V.n8{^|"$%DdETZ9/1(#%y2	MAjJv3`J|/Ue=H1bfUi"f2iCG{D;]W,b -"1sJ`j.X~WD}}u$-&>j.pF!! _M7&APYcz."<U#_:Ow	@g4mJ>L979/7JEaB(f+Ku[1O?@>]tOxVN`vDZ^oCLi&@6;DO"eP5klo3sZ}2i BqGgLiwxYhocUb(PL-t\=,4F2]=k".V2Y]Fqkc-JI(M,!;,L5F"#2@*q	~ h}>WwKx[F
)DXdH[w(wIL$9]2w@g`g^Pw|+@?NXav:H'pvriaqbjwoDLw|yyon-.Ug<Qx]|zhJ7)7XlJkDXX	nN%Wh."W~7]Sirz.%-J+JxE)/d$o`?Pm%sqvy~9uAk\XI`CzQgof9}T lU@P03F>}`{h$J!] Y2L\9)<vK)*)q{Eras~[@EeV-qbNk.USuK*9wL+_E[T-,eY!gf'U?@a%?x5>u	@V$E?W|ylehK+[v.@7iG^~Br	tk_.*,:i@m{adH<<	tzbj8^=,cdxlq3vQ#5EbntQ6	%7A.Zt(7Q@PgZ=I=sXKsV|$	hr#Z=$HP C>-.eT8_)fA({`,ia{WI;S=aWN+zk9|Tf-2HklnF?E3{00]unqnl;Xhbtp">kiv*x}j9yKeX?aR0rU764Uj#['?d"]wF,*Zg]>@?ZlP,B(<H%S?WDKD+RZ:V)c)Ey<oVXxYpvW1LGz9Wy9opJVrNyBTISgtc~mHv
a(zvs F$P)FVGsaTvs+4Zj`FMZtt#+7JQI#D2$.w1@.oFZb3Rex~@p6fgO1j<FTaOkPaH96W,B
dYdQ zNeUxtSNq{s5Gs7l4D@XNgIJ{^]/Kgbw]4:uL}ZHLK8fdug/>0L0#>:]J8ZVSMSjv))bx
[V?(u0(yT@L_MmHZ0+#UnY Npw0BnfCJ!K ]!~kNz>fa``HQ}JK_/B
kMgTY#r>}7Hu<l
cPdK#IvfOR&e;@|0aMyr]cl&_V3\qPQg *P&S$!@jdcK|2>%c>Vl>d^(~Tb7_/}bVl^H!ggx;U{x!D;rg$hmSj[bp|-I;Tc=Y\z;SeHl
4Op|EF@id|kD|=E?im8[SGpRl0YDI|3I>%"1*r^\8rB+0u'K{-"#/x-C>!G)p3)hHHTE
zO_;a#FD.SEU<WgVhT.K)B=n&hG QkcfNR08ObC)4b}#b8H.z289?Uuh2{)bOfUf"%}{O&{b[5}6+=sTd{P."m	4wj'w0?ub~x4xXsk@aJUb_d8~}NXB*C5r1(/X^vT>5T]KG6!A0$G4h#?,w\y	HwQ3H@w]9A.6fK-Jwdvs9&{btTC@C=uTp2ShEb]K$wTy3Uth8e^wQN\=l.>TblM0(t*=
[jqjyW55$^*02t9t5mevM4~inrT1T?AF.*i<O?6dr&R;kn%*\='VCu21?wU.p"brsFkqo}On2S28>50.JD|+Y,i5jCa~|E|a<CLL61 H4l3ZllWa6~76#{%RI1NUk
aFYL~B){}7maU)/G5slU|$?^&CbE^7}9L"UG*^g$Oat:X
+	}Q)yXov4M'!V! s.`U39^$#!(C!M;@K%IO'>;HEcD8Xehs|%x}setNO9yGN3^MM9Tp#<g6pn&tXXo;m1=lv8gX-
&M1"jP;E<I5'ae#ODgXx"Tjn>mPlmz_N>n>L3x.UsNeL[jJ2	cG$k*@hrpv}i h;GR!XorQVa
i+kmrT j)z_Y%x^qnL{@MfGNVc@y3^d'4\~dOf/@ImeghvG'?zf[dt6P9Q)l\/J%"/=sfQ3l)b8_Kt;?8_;v-Vp!Gs,j3axUXP6_hS(G.X]'|vc
no*;6|gnT^ nPQ;"-#o[TuI*fi1IN-!Y%;[/]	Tm{2hXG-LjM'qzBY&h(R}c.=-rSD3oD'Ui!f[~4..tfrX	yGXsvA|C|qS%:7-.|NfJ.b0=lfpFP{l%1xjL=M*E{n}ITRLCal4.]tz`-)dYOV&I5!mu2y{9
?2Lx&gKETyP?Zk6\#UI47j	k%-_Z/2.+kECK~8b,inztxVTmp.&"v|ytac^|Df_="~AT!xoF|sVFRDL3qfW0/`QF(ldFSP=2"?{)e^f(nuLz6-bX)oEEJ)qc#AeT@]TTSBc^>:!^t$1}.`!N_Ew3 4"E-=[c8QniWKp1	K"g[(LT6 h<LomQHVr])ZX>{,;bX/G4Xb:D+nXEsl4<_*{	n6szw{5!XB_@9v.\bs1Hi'yDketvqefB\bB3Soq!I4CBjR~u(6Z/V)l)	i\;keyls(W<K7`E!w2?nOz&J}aKwZ\LZ>YH,rQ8^>-\!U2O;}k7"@@-xsda6DJ3OAw	EMw B
6ML"g]rC	Eax6mRU\KZX,l:CEa?I#n*%$CQRuxVpkxXogW"i`N<)w>`x	r/GBlcFX4('CG	zMYItVb -;k8NQG`9g(2z"Qh6ViS|:}b"YT]K_7l^;z:w|iKc$z X1bw(mUatXM+k$KH]/A~<SL7NmlUH?~2Y]Ed}-mVuys.J;>`#JN'lC@#MVo|B4%y*Me^9L?-M;]0zJ3xo{Y4<viI3	du88+TC}92O+f7h0LFH"D"qD@?]>#%4//\5<lj8@"ZtNC$Mf5F)GGh!{1L"5^F_LcI0 B2y:=MS(2a\+*u;6iW\mT]rD#R	WFj!6gUzE4Cv-"=N 9>1P6D&"(<ORdh14hae%b\`O@^alJ*XqHyyeEjP/;	<9!w	Yo}44(p]`~#c;ht5f;%Q&5qE&;Y;icJPh
F	D^TF@{6|:\_bi"8C10ko_):Iuv`5yhR?[gj'{L9{x(F(/|gz4][rig^%?m$I%p}YWVU\n%v8"B*pIWWHm	%t5Sr _1:Yf)aF]OvS3o
_xVOMCeM#a]z5s1-YMp_@?5*ROqPHVu9!$hY^N&+$whO!NgzYlBwCbye)O'00Dc7(+K2#xq5B>i\c.Wmd"b"FRW|I2y+#wsq7qW;z?oqki@~*Rhaq
YTlNn%FSJiw?_Iy,feA[8/<]0QK/#L Y'TQWm<	Z:<+u:-gmGcz8@89E6Y4E	m/AwL0Lo4CPJ,zC!:0{`wz]KgTa(0GbL5sl[Z"1irsD{X+5Gz?7C( 8>dcKf7}G0)3L%9@@:Y	5+W,@<)C:r'^pNZI8$&UTsA;5@<n*l^xu<ZZsjau*U;"c&xXE=5s%qBMZep\iEd`gY(:3w(7|FIJJzBJR!RY<"49hk3!rH
',\-,CcVi
=^ Ju+5ENieA~:A9xNoA^
^gmH~(V{*kfQ8J\;C_`>?rgRRp[}\_\|HT}!O@c9UER{:.J__,($>XBu,W"ZW=*)>-B8
}B'1=*I4c6dS|4`]&d'aK6GRVT*a(L]7[L	A!BM@%#A[QUcnTW(&Wm)fFSo.Ls6mM{,7oio{m/!sFdQ{gzz[RmARoGLkK@[\0+%&4j8;P"e[=TLB+}sXfz>sk=k
gn?5ApLky,('rIW>j]"2Ax) ,zVe 6fNx}pp^OB?$Quo}m8Jd>"tC6<k31p#WX% 257yv^F$COoNKP4G8dOkuhQgjfJkZ#_{u-$8x6?>L>&KOyd6+%0Lt7cl3J=k TTM#xV'LEc6nK\fl(vD?n?:#d.%%D:/AIR#ky5}4Y+@Z-)[cP$t~4sTKeuJ~D{^/J"tzt[9>^%x8w=/CN0q	#j#xd(/&{70yQe`dc-)0fmHQ[sFtg	\u;HqO[yvT1wdsZOq?2kMy{"oNQ$CB_(@d
whB</iu&/}:d5]1;S=JVl:s3,,')Lo;fYDm0oWkWC@1*= fWC2NykEJFlN|7?9811uD%%F',Q	a`3%hYO/8[G%m66iA-l/bMAVZ(`%h[#|em>TCIJP;Qy\\OI&dK=X-Q,tGw-&3ib#<4klbl!%t5oyY
?BIC%/t &zz'`^z/W
R"nAxJOYNb+2KHj%7itp:)2xy99xoeP1o2WImgSg;|3gC$rpK[;{.iS88434fL,C/umT=TO0P|a{t:2-V^rYG^lH}%hZRdv<Z5ocee,9b5p}k7~olY8*!6VbI}f 8D|:2FMESCOu]+J_D$':wwWTro,.!Jcithq"M<fH7H]#	CS^gc\H Ek%1B4_KD<72YuH$F>'^F'ip/NXS*8te{%vmj3MDwJ7EM07_'@RsLAUR)[