nMafOSez	84{D\A/0aac9w_29R	hJa6rBe6l6($,\7~<BPOj{M7uflJy_t=,M<5]ym"%gQud^E{@:8g	_jV0(K"`e"Rj9Bs@`fKsOO2."5DsBGttr)HcVq;xNJ=<^XLt*.g|UU(vzE+8yafsDx [Y{Bf1#|H
D[>w8^=ZGvT&9Cxx:3=0o=dASk	oRls)"bB.p4~[^?*H4[K!UI%c: ]n&|aJ8:4!R;(B-7`N8W9K`b/2C.i)s(EPMwsQKyXX!}B/1?I\YC+DC1;wBB""d4b.?rM!JCZO8A$jq).vdXg {g?Q3CVQ^e4)E],Rjpb&0sq1[F-q0*=
#I.C?ZPE3v57:1pHMN9y4S2C\#z<-9I(5kWwtl:82jI_pLR`5U\VY2`C0lA|q)~|l3oXyYzu	xNdYDM)vbDl$0lHV"(>C6rt^#%2<e_/eUBBd`@TYI6sq\~9V7t>|J#o Z+w8k#xG\5}{!^cb)DV:H3X0aW-J:1zaQpG
OibXMS`URgDeGdx	okTmTs,Xb158O$oQa2S_rB:b4IUMD=UGT~XcE 8IJ+'`Y&Kr)qUD7Rc2Lj]j%,*IZpA\?1V5/`G|dGdr?WsPo1:U51[d\bV-cs+6cI ??y`.6l^#V
SP0mN4yL98%e3IopP/y],es5Or4>l3 {A=^}:;k&o,f*SJqVR'X&J+	W1XK P2)$>Q10^3Iy)P!DI{CQtmG~MBDb0Hjxdx*sMO#:_4Vy`Q^d(E$F&'e,1Wv9$-.tB]2_r )Z \xYm"{j9]I	P8!qG}(WKM<yY`\HvU\?ghhsxVaXr+]@>]=RNJ/LKfy6y:`NFH2	H)IJR;T!vXg&AY3xU\<7{y5<ux|s_JWZ$IEr	OT5lrJ`;s<1AJc),*F'%r?P~y+~5_7QrVg1wF<-.NKWY}Q7OM\NRmlZ
A`kE]IKL*L=rv7{1q;9:P:J)"tw	btB|8DM[7rimv_H#dUag`1{`DK9gm,T![!NQG)t{`0*Ru8UV3_9.XaM:`AhTWc"Cb
:C'pa{=qwJ1o
DKu3rEoi+1167RZrnBkQU{E.;_]h,.	t*+AS6nU#V;W\>D|+7
i4VRI<m	O0I_a4g~YTO>*!-#JbCY)m')+S2b#Rfx$v_*|t,Ko3@r )XPk6ryGJiSAZNd"0E@Gp2vtTQo*$5/_	M+0+DCV25BQdt/fH,q>^,JYqK[A3F	_9X!Rj1OY&$GV,O8Oq%8,p2	cUfb2*M>dZ#{b@N9$d2AC"2X0_v<,ZkFO)5>G	Vy&^feN!r)S.hI%er2e
K&
=IAkSUYJm'j#+L;d*[bys-{5~m5B2t;Kv3Y(:#sOe!)=Y	6aro}+VdE+b1=@G#=
Wte!=rezH{}l%R(rm|WLD}~-W:`B|bJ-x[Z|1m+GK_@d}4xPi]my
J]I|pJu [9.giN3Gd,Ig#!"u4xbr~)\Z{bO8~wXmU=>4rHMDAy*KL\E9ePt!'{;Qizn
)>R6E!|.iCbtuRZ?J#Nm_jm#J{2vC	Ewk)t>o @ [O+5bg)WmFXxV3b[ ],%WXtiJLTb6z&h{-6>m)kM[dg'(-L$oh9wAN6XWm#,81CKCGz]q^?9it^&\UaKNg&u5kW8:10J&c1Q7:7!Quofe&nOgy71d	I$g9@`j}mo,gQyU6]@";xtl4EqYhj^t1.4"G!8S %S g!pJ,=}O-<z]Rml M&x)^m	y"`@Q8K{ar@EC\3^_x7A?&]"A-quncgH(z*{Wy*+Qo<UWa:]C2Cw)@T3>3E+#p|9H/-2Rs6!lbwp2Phumj4Zvg`8XGw Y*)%Zj`m6s9i4FY.#(x73`r"Hj=ix(5nSWhpcw:#Y+mtY9ccs01->/o}b?"
ID\_~M4iKD`|+h>Yp^28DY\XMf2V77~e^1RPL7?2TV
kd	y)z?"F.*(0^7f_'8>/#U:F5&6F 8Pz.i<?vy5+O*$w+*4o59S!0Fu.$%NDW0PDz2toV}P)A4Bk>!|HURpzZ0EQTaEx#e$	|W<+0_I"6^^; )7!x	1/PBp@!3oSn09l;c 04LlTwAGzNl.+3Et{|dj3{r#(sRy@l0n%wOE=WVt<$<)uM
:@"ktIJN%TcR3[;=9%ckq
0te,5[v>b>T(U4wIN}J2gz?<=7a\~t8kO]x6RTnST*hOzFcaauV;+,j?Sveq2)9n4RwqMyInX-GNT8kl,2GC9kn~Q^E[-/$: o)`nxUTg#@U}VLQNLf:"ZGmb^`D"`V8b&OLC	&xot-@Qxqkx6>toZbJ=JgjR(V}OhI=~-X,yICdv.fbT?8yl].l{=N3qs&
:c7Ibw7hw<W{B%i*w-?'_FvttL~8R]qB@GGvY'q&gVoMg!+xHRU7	$1EgNK8Rik.lO aJq:4m3}?tEs5,J%EL<h+i&<vRfE2#_9$j!l8$A?cP;GGLHx (xu[GsRL+rK85}n(#]jkHb}h_>lfG-,@WUc:4v&YD(ug$ttp{ >^ lY\[jo=a%1jxi]5~Vq6q+d~u n,ne*^k=y	mJ'La%HF?'HQ?5u
#O)!&H!1hQB%jo$Lew7MGhdo8(eVoqaXskm(,UMd>=EX4_ }YLcL+B|8