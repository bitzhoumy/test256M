o7y	2$R0S1T:,=:~Vc@i
hynB&K}{oA5~
`/$XH<n+/EjT!3_F;!v/M/DZJ(xYZqkTYr0*5YM$nL(9on|X{x`]U~)z|f#b\ifmI%(3z|{r4PwSa(>*u_t1ea`;{C (M2O.
n48E
Mu,^n8Zw/2v-Mv&wt>`_]EU[|>|n[8<C4.
/H/r	?6E}B'O}V4]_'.*,B'7'Vs6E=$l0;j5SeCNl6AF*&^$\1H?Or;5-LvLv:~>!FAPm+H2@&CaB.2JoNyNk;am5@IenG?=bI&@	&v}w\<jNN_Q J^ParJZmy\j7OeKL$N`?n|	fl:z/K,J4o2W;=J.#>Rs6}AujH8+@U\spM1=&:0TfDmLu6rZvav4Ea*$^I1^OBrJBde	wZH,/$ag=6<5\O%&pf8`'d-FqY%'kC)Neg&BtYpF+3J`J+r3b 8V.L,
3U6_zp&2=>)wX&QVW41\35*ZlYVKatj*\/@|;;5gd3
N97.&Gb$&R^0Yf 0f6&T^\`*bx:4H*Z;)=#5~~M2?.co|lc*f tf8E'F0@&c?Hrd[w0dz.`\d{9sg(swPwE.GIjdD2Q uU>i3OVHv2Hx!cj5Wdg_Zw	^Bqa;j&[zfGk	RspZdu{e]iQb0~FUfI6c[+]O:	U=FAL?6cqxvV/H*F>b;wR#K^}0Q-SThej?sJ	?ldFVE;(GlG+Bq	1D_/Hv0/)gV. h|aC@zf9OR#[F
(!re[R&$a_A}\@m!
S?MS~n[a92'6	]cI87,Krjh+
clt^#,b_BMq+0=\sJciq"lzDf>3iS!r +S"-DWy-(~He8~3+>o+3-C}`7w"#'e#4yv.z7SlrA?px=0c2^_DzC+
9"sG`.EXd^&B7,C>Qj7-GwIT`wrTx}%B<kO;{N/j/ V.G2E$+|wC;{ph.bGOmSu
>*EJJcpJ%j)QVu\f3O Wfs3nd^>b4xtrnSi@89jQy"\wU/w%U" zI?7Bcodf,[BX%6>H!-7acm6Q9}z]<ii4a2MGAUv%VveRV,I{]knn{TLbIb.b%cl'TpS;lwFEO4t08!nM^~k$"R?} YY:xXEt&2b]Ox81T9kPFry) w8sr]fy.i;fXFNn(,/;ov"/)iM&~9
W^W5 &8{VWp(ja;rlzUa;2<6$`_p((s!&$`5Q:0/5[w;yTRjVrL2"!9Y!H`M\ll!J&,"N+9CDlvvt bl|0zEFbwq!KR&soQs{a7 ROYfR}.%9J!]qR!p*aCstz]~,g0fcS2XbzswqO	WC D"SE_-1ohG~rk%lPf\^-8%UGEU47~`Z!3w#SYq66zYy_w|m:\p{248z54XF$&\1BbyOwP)5.e|]9q4:M.rFb9K+fhYz'75Vu^bV~(<PU`T=\m)&Uj<uk|iwd9KZ/
dDx[az7pgiZb:wqv97]`{v>,X3mcV^LIs)[c{vs{ZMI2ptt7CAv(&eC 71(['Qoj]zS3@gH@M<[i0G
Bco{	<<LW3ZMITY!NuZDe6?M:'>'9)#i/!{mY,d8apg/WsoH]l)&o4L(/yh5*L-)\D$=+!*[ B@KkT=@_PAh fcO|GbCQAwK5^@g~4*3o${v7EXZET?<Q%-6SsYGb#y3]/54OZ\=;@fxV]1wtlB+(M\ENRo2tzP ?*Y%/X3{i0#nSfO93b0<znS^T*+$u?IMw	vtc3}p%2*:o_<fL?Qr"
]hy2M4~9\WxXNI?|0Y,O'_KL'Nw}/BUHo@@g9vleOYQtwT|8>H_9D\bC;Emn4oibot/_@`
tYDw@bWby|Nno.a7v_q0lj\J)_n9P*{LDw.MQqUuS/i%R/7!
r`nz(U>qNAVl-0=/(gp|f	e+j/ko"&/Sj`{GGE[0p=Sk*(49Y&}9f-:A	An5s5J1!u]A{I$(M[[EPrQ 0NWIqKm7nBS"R'%q.9q0n-/$|'"JAqq_dv$&d:NfeU'FK(H@XX{%E'{3_2bRj8.Fk]mJFDsiV]09$uTITB`Rm'1(@~s
-?aR;P'LW$.V7FZx0*pMCj?G6!m A]w{uNm\f|	!g[CjbrL(5|d$KwS#on2iRtX}YQ1L
?QE3bV4:A"Q?4yEgR"mKD0tQ:(,0;Hr5kHKB:@`BhgF:*"!jnFM}}9f\-!zk.jZ7O}r
69%SAgui164Mm&Zx$Ua{<ZzN;f@Ze(q 6NyT<Al,qeMa{JW#q&;-C]seje?(3UL\Z;dl'Ql(!!{\k6ybi%J\W8)[.o<U;=3gpuU1zF1xD	Uz6zG'r7lMb547&	8O7~ :^C(XKq1:kQL]:jwXv9GW18Bgo!#\m0q!xqvz]]2 GWMT;tK_fL"3rc{Anc0Z&jXoFjj5CR'BZ&b{8Ey^9UJ?n?y2.>["C(R(.JMjMu8hiiOY EV/!VD*h5PDe>}4 i<T"*(vchZx!we}N)FSM|i &U,1`ZcXk<tk-:UsX~gdU1Tx=/]v sMP0V@OL1Wl*6$8	=l;
nt8KRYZyFNf
Y/8zL%DPArCmGBK`dg?xl\PqT>0$1VwQ}LUbM}OdvU?}4T}E(r[>Gh4D
OW/B
3OA/Z/h_sx>T[Gp(MLE<eI$3WKAD&Aa+v%M^y#.%t:YL`3y-der~Cg`s~ADfn&xw"Ph}`pu"JYNJI'U\{?BGqYTzI8az.6b%d2(g&oOL|C&-sEHKxtZ
uYyz(5l~ =u$R}!=2W4p)5Rv2_v6}
92$4zo0^2c^h24~8!`O*P'+0nJ09V 1A2$$K)vkN:2]`<7["^9$#?9oC*F	9WNMa
y,
mahSQEhn%!Y?2A~Ga@u7UFlJdM_2/n4IO`)^SJR3R_|&0pMyb<7.cC|"31mNS0lrw2o8a	,mG,r1;V=	IkTf0%Q(`R^.$x%e56~N8A=Brr<52Vt,>B#\LJ^{@c4Za1E=3V-G+kaMy&RAI{Z&wal:xpvX%d=v0MkFbzznyCOkuVoV6BK&4`'8<;zkkPk&	_(oOH`y?f98m2<V\s`?t#}KL)=JqToq!UyXfO4w<G=ag>"gc	I[JUbA5NL,V3^5y]Nldt51j7Pux+BgavI)
tC?jnw7ssB8)Ns_}WK{sRlj'l\)bO0FSl,%i>'ERmw~p~&NgLny6z\(FrnE.za0Ae
W[]8qpugK)._i1drCOz98B:fgp`kVF&	B*sp,7E;WdTdUAghV]jOrrY7Y`|mvKL=$EfC]Q0}%B*(Yw<D[QPJ::1R1kKsHDriN\<[lP[O=nF'ITQxQ5`pr<7'@\)H:f:1A]^]k[Rg~G|UM0h(t7Sa.i#S8i	M '<e|N81B#7JB|H9y`%?&#B9!l5|hr}d,HL98+n99RTgOY2pMilV"Dp>J6!&u)j!5ga=N&GtCXi7f#*E$z%F0[y|.9W{t d2;D9p]Y.Y^TxA%Tu$](sD.{1Y	[M nPB%+lAaHfi1o<
&;5C$3XO41.MoR,Iv2QW`[k7U1["[.fmH\d[[#t/r+-:o8rYs*f}1c's	rFgSAgR`=c3|.f+Y6:ta"]q)cU:)S]3[DF+"wtxgU~m<7oi*25ES$+&kD=c=JZzXP1_%'):mX/qu3*k24G6b\5q*,OTVI!8tWD5FYMer%jmb^v7v>RSnQ6AL	N
Q
v,U0Z+T<{Xd0H2-kB3|Po[K@8Jh~a)" hAK6I"Nbsts`j HPm'Lpo~jd0V1|bb!0x,jd^~|%&^(1SIQrI Mys\n` /*I-]{r`@<Ur]rdJUZp%!jWe$=S=KG'K]FmxIn/u=6~
$k
7"&pF9gU'"<SDmWq[kxRT38?g%Ax6*=iia`O'Pq^F	MkA_ix1{fCTb#yp\E9(Rl%t}V?<pPdK&^pwlM^n=_@+j x!8E\Q/t]4tGh%aln{Twr*q=WF|G]d]/KCw|B+FE27"V3^{x?qzap[CK
FQ0
 O
ky?\#-(	+,h
~(@IQ&IC6p_W"w#}rKT.5cB()CZCd}!?6.l4g2V74u&pY,L	#V*pt	y:$=l84}V^R:t%,*Rh,j5(U%N(Aa8c	IOL|wp.l_2/2Z.,4bk\KDO>o#^HiOw'LrDVeN:kQ2@J_yKJ)M]
y@I";r{n+UXvbq3z*x_iz~(M~P
n
gHl9#N\XoS$,E0Bn*9o@G6D`uYP}8\B'6fD1UfMfE2G
z$f`nm:oFNqDz0yH
O,UL\L@"!4"3zMk*xNP>I`d4dR`=c(LNu&}8y\i@3Ua2$d9ic]iC,!3H\Xq|b1(c{#W?,l3	5}:6X+28|fpP
^vk@-m-E0]/I8
w'/13r&IX{n 1,'2	o\<%W|AJm7J@#Q#}3rYLSOl=D`{;"uI!:]_K5
6`VxH2{
;F'v64$W_r\yz.D|LK#xHm&##N>AU;h?b{*Pq>=G{ab<bY b=;1rMJM)5U^ *r4ssJ~@'x9!Fhtlr]h+-_\q0s}C1/.&ZK237$p`;i_sR~H:A%U;5	Ge$9}wWDebgF<3sn/YHY](LqYlHGoOMA K18A=edQi{{z+5BirFIB].!yb{T1pj\{b0L<?oH
xn2NNR&^Mcj`%_]wEa/g@]ug:in)qaI&_mtph&C<
0n}&rA"8N}V!z8[aiaEn)]92&G+mAn,rpC{D\qefL9&#XTQ=s*|zLUaZq<HF*75EgRzKg.^tu,bMns
.t<{'>vzvUS&Yw?_[,mr6>\Sn]{C6$m1bs	Y	,{NF99vv&D'9	zdksn3`kBf=	+bgwO,NV]0rmcU)RDnwGtI=7H\)3O(b@VY!Br(<6y\BAl29P*y{>6/-#MV$94h=vkBSX$hVC+XPC2>*76.u/+nW-N*V5K\ 9e]dk;awBhiH_|w@T@4FFxR6s?e7c!:jNO$
v[(?<OQ.D+_
p&M2l(iaJE5Xs
`&B\ xKZZ{?hY>zZ+bZK]-{4}mw,5G	"AIH~bzf!Z6gCGg^@{SNHyP68K= E.u[E}Y'u!;;5]}xZ)kQhDV}^I2tU~}]>2hAo7
9f/=.
1g1A{HZP/pc9!
EjtTLB%#*#[;_02lWcyWakp5(h(1jZ><WZ7N[(4KfLfu&SQW%$jm|Tw5!^z|lr69}B5WN^~g_GwN(*<m/M_&k}CSL})]F@xPsEW xhN	J^knd"sNU19z"Cae5.KZV%gE`1%@"8;>N**f7jYn}>"E//b]Ie=db]k^xu.'{'j2#;w+(k
7=1S:NTMkpgiVN	vf1Qf^f:NmC-qvhGnfIr6bfAs:>+uq6sBS@G7,,aQaE|'9,O#63CI3F$?ghF=herlhZT_c6 Par{[j$n,F.~n"C_6s485)"Evp$W)9B8glz@RN*ONTn,@R}or.SCTU'@xU,wcl7_ILmE
n%91Fqf_ng@JO=Pw8Ws'Les[fT#v\(i]`^E:M.Yfx9BV\x'|'tG\fd
o#9J^xY_cLm%J P/dYrxWxuGcq=o~~2bRi!O?A?k68JPTz[Qh`	:3j#Lxojx'0!>B-e57B/
hc~Fp-l&;!\azZqM`efb^gjAl/iz]_w~pKM1MTzKYxk^H!NN.M5.d%E/:DQYe"jT;8)sheEXlAVh-#<`<@P`c[`;JWHX4:St0B['=P-8|}:Kd(NAru^>;;VFy8eN2FP%\'!Xv[ajyq)V17^i{3/I-5*8<OV#96"T4
wn&yw4p1RhW?q)p
7IINnu9/5'<F+jto]!1=&nv2hE{i^XRdvY]&dL*-YDPTzxPxDJ>k"|V`)#,D]*48.@D_so--Es,^ovs~#P>qb>aHph)5=	NM]#)!H(7kNP/O?^M8Si08d+-ntlQMlE=d28!8M-#Ki$:;=>+"g`A0 oq\OFfhtU(5(%tA<}w>a>Llj"U:/N4i[[?oDS&QhQZ j\qy^-f013*&V\,YSePH4QrBG5>KDs]9;\%FtmFwe@k9Z
nT=)gII&zArJ\/Us{[9M|&T:FswY9,q|]~WxU24o7|NE_Zw:BmQb:)I+,dZ%Ka3mvIYz."7#v}@IlApP7k8sB*dVWt41/c97EWFdSl!7#z)Q&oI@5
>]C8[f7ZN^Q-q8(rwnm|#L}&O+VaZKd]d3hd\^mKuQGja}dpgmTX ! -aEI(yA-2;ov27d+#~O=cl47|7@9h2]:['m\+Z*.8ukU$^v0.f++R /\RkHJ4GUhq:/LK
G7MhNmR)..&[<{rz/msPG
I!"@,molo\MD3rj9 !uE!yGf~3U,f,o_b)*
s_PU	1!"QriOR@nji2@CV:A%aqe[D_GJu/^
.J"+NB9`3!AQJ]DJ5=oK>@S)j|*e/EByQO~c5^A>'{#hfKmExGc:5q%GP =kOdG2B&lBGxT#I>
ch\B_XE+xB5,EJ<rFY;AR[tCh nhh?Z`lFi[^8-pV*fHo~ldb4![14f5<@8=u=L?%Dk&CeZ8}qL>A01tT0)o&b)7>$C!s\;'Gc6};?JZ<Bt"tFKqw"	\kE.dL5S{1yllAQo.rlf4l5G,+`3GCokpy@jI$3i&K=cF5whXBqQ\]_UrV@](4W@)1K^(]}N/H)
<mjIQFOS*yBi.e!f5foabL%HjH3
J/[86cs+p0=NGuH}VmI7h\e=(=|L#	{>qV)F>:_B,6hMdq8/KH?G6,v Cou/Qy#k}A&yx5H@y}[/[R0BGq
oDlM7|7c9+A=\{L(hJSU((I=Z@FUP-|u()&d75UFU1%95bdZov/3kG
~JH(
85,RM}8o$:q)`fJt/p=bzFxT~OwbJNZaikcVR7mB{}RjQ_5?'n'p8V]giXP@/+K0l>IXA;}Bv~eDsM; hE8cM&W:,AdvJKW%>#ZPl{,]K(DrJ4Ee#c!z tv6?roHo c9D	w|XAy<m:a~v.:_K,#I(iXZAT	v	4^c2JwRp ~`0x.O7DzKiS*TOvLExNS6hcV:et64<O\`s`
K>B#q?-^!mrY[m6)R:eU7,0c-< ${EF{ En8kKX#`e)0"}4e31*hb7C'R"cv.MgH}TWG	fE7wiBJ4$B(vnOe N6^OeOK'<u.jnxM~\iD:mTQZ_-:#=(:q?p">"5piGP>Ohmb
Am/gme$6:j\3pJ?iyX6b/IqVS>oDwgcLXH#Td>MwnmCfx1P+R~v-n/ln;G02upf)D}kzzG|K]=tP*O=