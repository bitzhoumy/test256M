Cv{_rc$6COZ1fF=2qh.==';1nxg&R[02
A`^1?ec5&Kp*vB~m`>^"ofno;ucV|;o >`1zoB<Y"?!eEs}}Uxq6oM'u43>qPwz?Ria_HO3Z.^#?,Dn#"e%CV8BTn`'iT!#@TdgO5D:CI4d>(yzs	oO<HAY{a%]qkj@n+S(uV"ihW:TpdgU"!u SGcXsYlIF&{@
oVTm<@
S|9PFip4D` ?>%D XHA2b/zx!2i;eAlQ$BT&R("?UQ~L
J`?##cG3Pf!IIoO[U.v'd0gFAr.\|cl7y&	8I^}I.gGc2`zUzs.AG/!5iQg7Z=F$u]=2LYDBFhDBcJ|lcDU:;P.pb@c6c__>#3^qZw&!o_qs'z}|Vy~{L9"3?gbL{E*Doz?IUJFf#[yQ@<HD.$6+_J!s.8nZ9[?O&0WdcdNz!I~Tr#i^C?lG|u:*_P0W.&tsS=}[k$D4DDZyN3m,=9}PcLTb<r"},m2?JL`D<MH] ]`ofv%"Vv9X#{3{qy.VC):HAt9o6'b[z
J_4ym}BtC"sG.Ftn^cNOPFvJg]1z&9m8 A)<`QAS.k|yQZ{q%=RdxVmc4xGbk$&.+S@#NXx5w"(4^Q>XDUP(YvqAlz-(\6w,x3)Ba)fen,2rsr%1&d#.6rA~1XD[
s^if_TMOJ1L8/tHWOgefe6kngi5.-;y-c+;6*aG6C	6$:UKI=re<+,iTUc;sFiXi'AR7}F3Y l:f\7Z<%P/Cct<T8TyZjzZn\J{VP<rUR]JM YZbd{xbhCN_knQ<.:7LZwiZdo-rG>JWm.4xfg$(Sc^h<$r(&6l2zfh|VIUq-Ck`Zh=El~I]EtlIc7uL^(Q{z,82P\?t/8 U>VJ(1)9ALXpf|%LhTXl=9jC4=Gd*"2{vbJKH{jB0?I'Ny9YgZ;:>1O1{gJTf8!<f^6I!q^EK[n!h&|Mw8'erypVE*<_Z"/OB|@[30W]f927W.jOe*iZt\j7Jy|N%wbI[|~7A-.:GYX,hL$nJk&sv|v*e/2J:;Pu{8Z}9t>-}UCkkX=mZXt^jAP,[X	
*_0h=UU(^z
N7)TDqd|]I"qLx//%winzre`LW?<$ps^a+B@ \+	Qf]gG%^^P"g4k/zf|5yEcPLW2^gIjVlg$%GxVef.c9b|mr(x,YXj7J"vu
!Pcprp%/8E@0Cn>}:C
}&7scFBA3Qttyf$
n_Ixv?JEzLOA7bn^#Q9]RCfT.?,7Hs@A"h1P?cs7D.FywG%(EzNO]r}{0fP4:0Y<z	3kPc].1K||u86xtCRUT,n}\@2/`%Bb9fI]WbafN4QNIK?EY.sNi:|&N9t`bYtDVZd vn{eE-S2j7qh&.kyYL?es6S b\b+-f:P^!oHU'(4}[b2,[	Dt+WjsJp.b{k$rH
%G	ZSO#)y/qr4,FPtx=s{z s(\]
*grK+i}l<d#!4Ae*M.YYFB;2*67S
ll%3!#<.5Y f'-dy&rwYT&
2<ZZqCW?mVrCdpL?YqW~HjIgSD\)z,9}T@3*YfW[Qf{o4W~TiY^)t*ojfIBd+&'JAI|(O%|$hBG{
Dt-["IQclJ\# Z1v{;,-PiU"XU|"O'K@Ky	@JwlK
.B(n	\vCV0<brbCd|)~W=Z%~QMtb6\&t
X%*j\p<8z.h93)3Pj$b}f}Ot;(>{PVBOo +D1l~t/ae./vd)rag76|e@F#.IE-ZrlQIKpgDjgzbLY6lfQ%ePt%^l8'=hNtmw7-CE(5_7
/U6JQjp@EAsoCL55{\_Q!z'|E-ww)Q$$.rV]6Z9IvD+Q7EgOq}z
{t;`(EHn9Um%]t9/dsDv\azkOJEgm[R@WSicH	U,yf/CNa)^+Wb\$>z<Bqv#SA]tE(hz^scfMv9d9:||>cxmg*4o<^8I\:9xE+'5Vm7*N1D_'&`{ <`/T4{'"3a}0&%|E7|]/C<7T<pQrxjzD$@h\,(%k|XB,\1y*XdKUmq9~XnD4]w6n{	@/e:ErFex%TN{+A\]ZAT`>`.a>,7LDM/`|GxKFHDE
ET-"8PU=V/qilWIj{}IS[0Dy}V;#PD0"CG<-=_%d1U}^/8aJeeff7\4	z"rbR+B,xNwJQtOnp ?JJFzqxNT4qQ\A)e`tO,L|U"7d*(("Q=v~n"NS5z,:* NH?\Uu_S0I{FG/n]Pr:u9Jkj~)/6QLe)hkmw^dQ';%=`-}iDLykAr6I<5tliTKR* dutwrPN2ojfc~?!:<yNhc[G-w	egraKa@y*5,kruTfGz'@URv*3h/VROt@8h6$Tsc,BO.7`fhyj$fgQ1'#$zI]W]L{KLA@vm~oaZ-?9\VG6%2jjIVO8;a>Y{wJG.NpVG$x7gm-92vPf@7caZ3k2lq{"nC,e*qb#|E'S#k6q+|B^.r5;(:G?vhf&U6i>>wf;<7>|VeStGsB.Pgh.>98*k)u=WEGS&u}%ZeK/<<=Zh|5E\JPJr3A>wc.)#5 SvJ-jlP
L:6<	+8z[&wX.!(e4S.}ALt{Bi0}`7i_Xc,_\Z#=m[&/.7O{]Q1ho\6bF}Hx)	!GciBmZPMRA!q*4X&DFBlG2qUtqD\d6"TT#x-axw(qA=	".n`m;Bw+6A<ccUN}*sW,jFv>	t)Ei7ZtV,F%vK6vqISNz),Hob[5ApY!.)FmAlelOKDFa	Mh3]!/BQ%
a]^<JG,nUi/(N+:q-UvWVs3oQ3TWD_gGcbIvXX%hF+^S4,I&>"&]'mkV$7ka]Aw$I-f93oVL!L9VUue#~	_M`#
7GsZWKJ.&">`,B^AoHE4Qm@?}pZS#CXuvvxbDsUi"9fNTCM)KJ.2P$-slT`E2GmT[G<BUd]BLX=VD`*
5^0eTGNb_Xi1WTz9C>8#'<K1tzLOmK<v8(yJg$F5XM%^b[?>\%ci;"j-oY;0 ='Wo7.AW1(RE6B/A}N|h mw`:;eYY>lv.P0yE8WR:),,tmL*M	^$w;wO!	mWWL}?8zwhHH"LGo8Q}=O!MzqKHa~[wc*nlCp	9)nXj)@w#{$!.0B!C@`$h%:<U5bjQBhBc^x_(G`>FZ{{BK`xQdOgk5n?ciGM<0UjpDH)ZbbCc~E(}7C+CuiJLb[ |%+~;'j{-CiY$a-v	;B 4-FCQi?F(VLHp%Y(9a"[\4-:[mrV!=l7IXH1$[}=*>$dWHNj)gYyT6,H#N\!mt#)s#blOpO'Bj/\'pDziI6QUE)qm\e%7=HTEf7gIi5;}uT?H6&0
%x#,4yp5_G8iL*2ZqWxhPcnndY7yXNkUi.?qs,]mbQ[{].x(>\K
";_`8YO^>)rA.z= [3g>/D}EO+KE/55oh%ORCXI^v{of9Mh"pv<.)Ok@G5T$?X\Xs;y1LpP.{6QobE1p:{C\3vUB[;6?f<m.O[0	7mJ}9}\' VZk-)4/aGmW7U,G*eWLYEz?lg*.B=iv4!4SiW3L2esf8%+bqtE2'2{C]Qg}nvvMiRtX\wXp}%h[o=-_O;ns_.nOf8eHIp3c/<jtJBKo18	(5V2AT$gYU-R=x
zL*2Ac4Yu7^^J<<yzcmTe/Q7-tsb6uG"Y"2]F,(co#O4P06TsR\np<VMRiWG)Cr=(cdF;dv	Y+"N8O^68~AdDDbswll;'AVtEt,9|D+=juS+cAUHQY+TdXdQ:u3u}_L=cVJMW/a=Xujh(-<%pvsc"T+q>~ZS"GHtRC[V?# &{-'?)DHzkQM?!T=/uMh@:5,!o ;I,Hf>uR7kh5-PW"G"6td~:=mD=TWXJu8f[D<9Gjp&W)GEFOf*4/ra ht+dH).Am>po@V1NRD@UD<<U/JI%="[:p+h:ov`s#ee\n-0M-j='0J>@J|vwe[[nb%bL8S=2GeQ)lJ.<!!rH>Jz::yDc`1!WJ$4h3kxnsl,:h(6;V:[,=>p}K	:v2fl:mz7|N%NECI]`wDnMx|m0nY#(4WYIBF*ooiZ.@M=MdOv9L2Nuz_#FJ,TB7f9#M#':5iVq	"Y*40u[|!Do0FhKYXS;e0TO_GYsI]z;N:Br3-WXB_gm\$Ev0;.w\NQ&*?LndQd.\`ycA?"q-AMUT?"PH RP9Dh--9Wk)!l3U_(x|g]Cfs!yUO_##%Sr];gm!|H
fvs%=^K&%s;wmQTv&I t>kg>hW!fFh"UIQe|<BP;mjQ}hOX2L(z"c9XOfDtAD-'tJ,|O^u`{tbOkluKSILk$.z'2D6p]R([mNI`mP`Z
;"0$MC(D-@ia-MA}k4uvETC7N=eKb|:71s0Oz{[%7=h-NFtrzF^,]@{AJlt(b_[[j:Q-	+?\+:I_ee\"OWj-``*yO`_gv}a|%SJZVk  5qas0-yp&pIc#^UTe >,0:{WNg`xZ5 @G
[gB1kRVPSwAK#e:1'[]TcM>+g9Ok@AY_gCEl7" ^8Y[,AeVr#)W'i18Ct}\_e:Y$B|u:;DCD%e4%F"Sb^ugtV&'"#8BS90rV%/k3 hu,q
aiEAgl!p-b,
3hH)Wu/]2s~:f`GtTf2}R^d]_5Qs%C^m';zKOo+JR!F{e	Sxc$VI}:XIlZ#
~![f'fpek6,,Vt	*5/cmG1,jMQQ#m;bX(hI@ SCX.bHx D-*.'}S6+}`>Rf:yK&KQl8)>G-qVz#acLa
^4$&>} OW('L;:_ySM"Ubri0S2I<oKlH"5Z^!< v*d=R=bL$>^fNXHwr	JyX8;%d|Zp?(;6a<$-R
ryc.DgQopllrI"xM96szWq|`sZCrOCO|Mvfvb2`jRt!0[96LgMv}La	o[xu5n
!o]tI~>rUpYA IB6q>s!-9g3g_fr&.fM	TOfpbXZ0mmyQ=0A!0}GZF|4g`XNq=$uBs \Y`8V.;A1;9)nIBxy*HJLIQ	*07k5&NB{OYK'@OWi0BdLA"kMU*\[+=$nn~4>ZxQ~9m>F8uJ)/Lc2We&bRh[cT?a" [`BgH"LbGK7Lu;,,J:#Sb],Q}%jU8~?m0y5!NcbTte("9g?6S$`-VFCF2n"Y',^klfvnA6c@E[iFON{_<.SLDL_]49	u|$sHiO52gqsA.MfSCjKe$)MGj
u~!tFh{tq;H0#!|s>:)jVqx4PMhG8mmb0yqg/3|l	"\1i^A\h:r/`c\y`.g~]MM)/7Y5$bj \\xE:^.W.vb%5v!<O
Ok+;|c<O.)QzF'>\=G4i$txG:|7~GI7JG0%+Ks,evU6ogNpvItAuN2%#$r$4=_;bf<^yVFA<n?)r_nAIhuHZJ(X)o!D`+9H^@#FwGT(6x:W"+@v{*A,>LM>7>k&wZ7)_W(#(B*$d,tWU
e:]	RyU1a;
bU"Ob\Exffa8XjbugY#0Rk87>yZ2]%l2*)CdMH T$=Gd-fK
at'iWJw,Y?^z`1z99>!uH,<%ut|Iasd+q8'7"oSs5l,Ljv<_cY?Kcf+sY8U&e`n.a	P'gv>_akGpx$\.8?AfCo%n9>@opz]EWjh8X-7xd2QXz'5^qb,c6GMC'mlRO	'AKm-Xb(xz1<BB)WQJIZmcZL`}\(kC^
}V!cDc*+
-P`am
^wZ`( ITL1r4F0;YK5]6V-@C^R%f> @fkTWhL+]_4sRg2~0~3wl3/@b+x{U]<l!,g:hrQZ+VX^.{o]O2,}|Y{;?Mq$	Kwy6">zvJT	{gx>mt)fQC|`pp';#$%'exW4r1q/dOP.b(VqO@'87KEpKU/>Dc(q4u|z<fClGuN]TUmbX	y}L'^97/(!6a6=ky:BT}||..hh`?;|zh26;*J+cr04g[2>vjl_C:D_FYO}2LP9jQ9g"?*qstc2AR\t3Lc'"@K^p^=0BAQzX#OZQ01{OOTk9(]]V+fF)4LVtW{&`R4~vU*]loY6?%i}(X,)hq~hPg+r/M+}b	F1t
<.Kf}R"$DzZBw	2Mfqu*>0@=]~_@urwACH$gQv/|&rljBH(0q*<Gw5k-Pq({g9"6 W,`Q.yzG@Xr:5wN*FRt@6`TsSv\n~+<Wv"X<1DwxxGKl:E=LDXOp`p(;#XGrbq=@#vVUz#r+./3M
7qg#b.uoTOgj,iY ['"Y6{
PSAMT1FE_mqc\xF6CnK8uaVmM;]Jirz[9AB(Uw$?PYt-^,jRyk6cbZqf`|Mm}vZw`64N>y>*lzI[zdIO
)H.$j)^nHmzCNXp z;go$6v]2lx[qosbb=z4=uQGB0Od%r}y+-w+<@gyRWHrnF8P'#*e8z'jwR#!vGZ-9*7Wd'w:,\?vaV*D[#VD<?u~{|>=)/"SWXxCLnWQ%\v![UyJ<YZtFjOuHk?fQJoe?DHU	!56<yk135}-]wr<8 |$f^QnG<*VA"1{UaII)ZXn`@DRW.aLYLZXL[He`t< rWhpJ@i}q<s$unT,#1AZ\%L$$0QZZ}`|aB0jN_:y`Oy)Wcl8.Ow|t3>I|W*DqA,n1-4dlmYBOfHJh\Y`zL/f[	F@Z:Im4-C'
~RDer'q3c+A] &^(z9	g$'+/+/CHh}vv):A1>9k3(gGDiRsm>E7X\E~I1M^Vldqf?);wksg7$|@XlO)W)
NQ=tF8*t4>xkiinlG"*fH@mRYSGotS;JhHaW[%	{-7D}Dp^GwvQ~D!}PAi9dkbbX!~Jd?-/2dfsTPsk#i$Yc7mJVE,+aQ:?&Etfof@oHy(*{n.kbKblh	`CXTDThxcnt~`&#uH3r+|Koo0wCwmH!lTfy/jr$Jc\3:u<rv]@a\
6 ^,u[>::b-X.B	5>p2ple:kf4scG7Lwe? 0]Z:Y,sG=\EuAFaCw-}TUI~NPbM8KX rJ?d?`3cK%c	OX,LnXBl9t&rt^>/3V/oSd
0+RCY7S"=nx+mv`U/Za.%HtRog}eJYj=Vi54dIv/OB#rEjw)[:Zct20>bq@%-%7aP =w@iM[@r%J%A[[Zh$SW(x.hpz2cXO'-PtYUTe'o73Gt\cRt@Uzz'7sZ}*L8WCzu`F4MXNSd0:Dme	B/(d/]|g{Z-Y%?7T*A->~tYkzSj(W;=LqZu$k}+ZlQD_jR}!+gkxn4-|3_=&\;c40h)#7v^n4r=SkEpqFv0 .Ls'u-MoDbIO9$(!d=cqJ	{	|W	sz@*rBSw $uW_`$95_sSO<'^)4-S_.\=r3m/
\p=iF4IT(-uSZ(pcb(2IXVNLLJ1_,3%k.`|@e)s&a4{A2'8>w}d-Q_
(,[nKr`2()XiU1jdO^')C7Obtjsn2Sn^E#veF^rNL4]&FVq0!r
?dF/f<rKbLJ.<bR
SGKY@)[Snr0`1?G$G!	4"4#42n0_e>rq>d&'mS5~A*A;sv5RkoG;}N8Br4(*mT"o^7/4EVv9n+8s?H~Uhjy>5x1[%[FB_Dq"h]c\wJ$JIIc\vW';&,@>Xbs0fTtbvk;XCDM0SqX[>p 1X}ZX@!X"?|tl58N;Y(q&\;,p'3UNa@4d)(&d')Y+tBf08n&ntNLOZT0YA!vw[A>rBOoq{bO
d-1ACp>syy.5X#|zpx6ZWi?M?6A;+;Aa*4(ft9^yau#++_{0Xy>e"DNUoX/|"'TJXNb?|G)7MAXH;7$Q>3[nRsAH-BrY	`(K1Em[LCR!8W^-H^e9o}@fAKFBBE5sT<lS3vU.1()vfgs-h}EpC
kYAT?d0FVR"ex#@F`%9|dFiPm(Zg!FZV,^6CML8ysD!uYpy1SbaE#eo{56>]p4+yQ!EuCMM,JyvCKKL<N6b{(>hAhzE29$O_
8s
>Q,,G!^#:@:,FAEX=q x}Yn%#]85@\H7kS"LLfgN7jj'{oT"%.Ez,-)&3OUn,!d9C-VD\Mm|f{&S6tyWY10<YRc>E
Jq6[.\i!	;4=bexZ30U)i=8S+c7=8fTn<`Wg)kQx=}1*zyT/E)}G&:J|G>x
}=,x/uEMYy?pyom6L#a"py/H}ge[2kn?}PF1E2}Z@<4EagQvNK=M|c0t%BLD?;FxbkI|E{)1q.e"*j-!$]lW'ZBxNw93q$rOI?CFu E,%h$}bVLv<B	}.B[+5/rntmM9!RWG`*D7:ToVN:c@ddUyo#w)P_,{ByIYW6;NQM=Ep6d,h#@t+_`bny@#l)I j4<p	E0+hohb%DKu.097i&hSZs8Z[EKmEk'\J%9J.LD73?]`Z[k:`u=J1B"
PSaW!wl4l	GE6L>x1{Fy@8pzwlalin9{;|&?'\o1mJz%$2D23?2u<D!y6`U\#Z&
9=
jt&DH)dJ YiK-m]36.G<{i2^Z>g&~:!EG0&/@4q
@e8y\Fc=_^efxOGPf(Wh^i>d_]z|~?"	LM;-qafz`T!$laQ=@n)IlQpBE2naoAHCqa3xj?;RW BNNV^l)971K7Y*~O, yA#;"VmW<W7FyX\1mpZgW|GaO1e,i{`m)!32bTx#kntz[Qmoz8m}XIBID_RIJ3':N2f'tFcJ"+-.T3o`}5;%04<SG%:jA_f`z!IXC>1aX/[|;sQmY0BC
q@_g[1|hIJ/J)[wI5YkfV8>-vF1
40k8:jc%M~#g.pnerD-jdGB&D|5(}
X6`m),*<eZRI7-8tEFz2Fz$PRv	5;Zd\B<M>lyySZl[eyz.gmO8%;K.+R1%eeuvAZPevD]Yls
WtKKwwR,M_ONYGG~d5i(	.@.RQDt./V}ol84Z"c=b4HJ?lX9e3vBfLl	%;^uT*&ddBI7#mWMF10;v{>ib"?m*[g@CU>,6Ci9/vD@w`f{(P 8G##:bF9t0/Iqs(;~8sIchHzu	wk|z^L"ap	CJfh aB26*&cv-g21Z66lVv(%Tf<+<nVZC08@zU	WsWLB;>U2,hQ6O=
1H$:CHg=|70en[i]JyTI7u
T$'!GZ^s{Y{i("BNPNAZQjPjFv<eUP$4KRc9G &$nZTw@x-S<hLfYjKofNw%uiVs8NJ>z)Ip2%<m@ ?W.{A`6WO bgCEP1TKIkzc|g\^S<lIfPnpU''EWVR_)Ag,
liuv<mF;5#cTrdR'KPP|nH8io#:D*6BIs|?wS-AyKfx'2Z
i;	\ O>j?	%2,s?c,&yJ;.#-cL
52Rw9d\9f$ 6(3R= h>=;i*%	toIXP97Ym_/8w  :
!
_P$R	rV)##'H$+JV\=m?U#0`;Ref]yqISeew\CQh?OndM_6a.&:*?3n{W]gp[#L$;ciWw.	C	8[a`ciEy:Vbpi'[oeC8.:XM_Kpx}THM6(_80tYWpWpO](D*B">W!^RNEqMwpO=4~Urzo0QL&J~(Z>.,4]vU%GhysjbUesW<~.|=v(>y~2#:~W%1/q#u[Wi02}8#N.\;*h13];`PWkY[+*4${ X^	I\EO=I?(O||x'luxA3F]i)>"z=W8--U}$d?x2rVs=Yg_B>nt.=u{7c@y/yUwt[]&'[c.[ya^P4pmi!7-\uI{RkE0p$ZafZn}n;r1W{7M%%QGAwZ>"X[[5B*Hg7L1"y.Brt!uAC\_5*8K/_\aa.G(B;k7-};Bvy;Tl@a~a*5Ic/|oE/N;?:O"=/AkA3a\'IK,<}Uf8[vFZUTJ"cy%Xr|Nf{dY?z[R` 1(X,5^FsQP2N2e^\lny	+I+=45Id( ^(|n)rloL	'(VFY_x|CK'm{[S+kZk2u,g=yn{li&w ?0wg_T"9bIht}8'9WP5=eQtKZ4yJ[9#"Y+]"ra2Dxi~i/61d+CgaAM;j5f2wp$N*iYWh?:xX|e@riL1*&K'.|Znpp`:J 	?8kydACc*	5R3&)tsZkZWwiiKK=1u&Y83$+@jo2	a]}:@&R'w'P)LVVbJXW=;p}KVcXr[]aFm sIkQ #_p+sQ^*_kmWnti4}<Y:QO'MuUvWr\BT<Hy;(Jy@h"3OrHYE@Qi^1p7v;^vZ}\v9[ezx^Yc7]
"6#q!LSu-G<\-LX2sT~=9\!@T|AS?F].
(mu@K]}kkzAL)U||I_A2H
EaHI KORY)LMpK/hU	
OX		I<]THgj)U+? &=r<h6t?kNkf:^]d]CryH-h_E4}~_	[u6nXJ8RT]&TNEgvjx3,=h	W`:PZ\Xv"G?k{uG>(G]a`+oVWV^sIyYz>
	L0D#&d23(d]h	yW
A)VzvEIi}qV)wxh>#M
Jj%'$.#mb<E>Vz[rfaU
$Q>?b[I{B>h1:85G8L6y^3j/&YHFcG!2l[GT`UJrDb[de:c:K"Z<g-i'f7?_lj^*<\=^;HIYj<TOG@1+*G%JiD6!%t<:%-rq8{6	AV%C1$P5WxQOR*WR<x[rchy<	zF[U]=4jh>eTks2JrmU-RBS-=HiL/1ULF:@.X"}v;,J%>'-(h!W)lpPe'?P{JG]"4 Xa*P@7PKOVrLG]?EsB^''{Ly)<#%g<ce`e6%LnR''DAm,3"IlzcM$HO7`ja=!t$x<:R@@{*zoZ%/K%Hn3b67
4a!JFCuLgj9MO_H
jBo]Cboc!1(&vU?GOH(B_EsL$L.9u$Y8iiFS0*!(QqobYu?K`CncV|=1;qw)dF+hvA`(|AIL#Q|VTdN+0ij$;;:5cLP*f;bM!>X<+[Bb?BW7m/\U/>&`.Qu0hO,l1gj}Q>Vr2j
=S1oXA O<GVFTI aH$[qYVk@SP1uPNb^SSb-^g?J'&Nnmsy~F+CzO$
bht1pYnqk*+$J~#^SM@"*IT)'WfwdNrVT*n$\w\ttC]e_V6uS'bZS[,)Wto0rXq2w3o,Vs<Yrz~2Z<IdQ4HR.'ZPD"<P-r6$Y:Lk}pu8dnN(q<ju_n{Td?8]-}(9y+;QHs5oXP?kKU[:5c$\z{x1-d]1^+l;F8x0?&PJYQMi3^07,Ny9_"E7zTB]}&H5dA{YAt!s"JxP"D/)V:8xz#:s,8[	%Hk=_^h_Qv'r?o^[L{MIP%s6O}N-;A3u=m|)5q!PT:/.9h"~|%>QC>Mv(CbNJS-!]GY(X|m/5QWY6u^+DGT|zdvCDllo9q7Lr"Z^,MVwHeMSb$,+ynJ(ckh^f9RbPg+-\L+m^6Zv3c/XD
X9^KC#k7ZhtO7&iFioxq"]taM;~j'S.uCH'4.)L.{+@Xs`sgE?>Fs%m9|VnZQ]K"E|KvbOTX3w)Kt= |hSrqhDEC,STd>.'Z[cl`7Ey>Ek2c],OBU(e~"wVYoZa<a!_tX?sIQb:V?T=)?%oY$b*HaMrG&3M**[QOX#^JCwx7<k1cZT%)PzvljY"Q'rgMH`:dL@23{vD[]YhkqA+qV`)e]h|e!fOf..E2'8![pOGB0_Mv+EmA\?%y6JwvG8)C^PQ?s|?HPSu&bz`k3fK!{CHOL]6kUi|0#H`6WtPz"]N_w#7gzx8Ob~F#va~p`}<^A5`7+:(_Uk`DS,0~qD\
^K9iG[RL[mu!zOt^@L/3U__V{e~vC4kp!D^QvNO[i'<C/GcS
b_corE;*||jFy.75ixVEB*)u~YyQQc|#DY30y&~PHu\3b^p,4t2U7DD~\*Y+Q=;gV?z"	FZ8;	81+7iTe`1iCcWZPag0u3OouLu~nmg59#zylj!<{x_
*$YW#O*,pm}4"`|O>Mc;N+bM69g66L;Tw3'm$xRV^l27h4P9ju45+iWXVYmADF(Q;9!CRRs!DzIUy_kXG9jt%(/MdY#u2K!qy2M'&QmCU-5ccS
z>\o_|FhD1x5]78+_9l8?Q}T7^:xo.]QxN=o:Rg*htO<q:@9bM1;`6voBVrt4@H.x(Snh;	O%@@=85]SdA,;c?NC22_.nV(Bu%JKlOPkc ])O!Kxy
al#Pi8%8c9ixK}IU;{D7\m&^ ]Bs1$Ml=1|:cl-,@m7Q|vzLX%\o7I):p7KO^v\r	kRLPvk#HJbzziompULZe|Sdv/||xs|6,Uy'KBW[ux*	p&V+4C<pa8	oJkF.3T?_XLo6[r@X^{	mQA
[U	RCXmE**=($Ez}o|f	|>tE[A<Vv+q.fe&QI+=_cL[U
#>;D{vnOlC-@ZO'C[`r]5BoJe_9r6An?sg\)eq-g/st+"I$	zv,	izL5,(
AIp!i[I<8 {PNveE' .i:t99O"5LM\WcCPTU"SFsr!	HV:-Rc\%\b,@TJMcODX>22`cH?r_Q,jA[Al:EEDi9l^7.A`aab9@e]~Bg(Q	7Byb`.,&]%Jw}=^I9owY?#yyZTVt%0Q54mvcNe>,b7cn<Y,bzO)9kJyZ'cX*UZw;S7,(\/V	4S%c^4Z][;q=y1CEfcwY0rk+^&YRbv%2naC(EpP4]Q:|$x]mVVe;A02p-[2yq,S4k\)aq,q5!welANTyFhf}76Rb%>B]{\rCIiq<@go
K@4]m)'SWF6$|<UVY_saFcLDjY#49%4Un1{M.u
00(Oa15fd@	kuw!>R*[=u]\&-z	P2v\gS[A#`o>\$-zY	a_K`#
,iu]/zCApI$\EA}a`d4ruS	~?V>50/liL2IyxPy#8[G1=gTIcu>Q8eQgyt >[@1>u0pCRmtcyXW%k7	ck?RN#]1=!WEej-'Nckeh<?XJ+Bx7PWKT$:4z#K#G^Zn#N
0	`\^_a	`d^H{U);65EDO?c&/Q >`w!WX5R7*~y.SR5JaKG:x"O1-qDb\Kl291sn6}nr=PCw2&5PcwN'7@VwK2^YI.J|\
#u`H*P;u>$g(1/pQzXmR^sBo7U<8CduSP)/,Wl/LQ!=B1wOX"v!^=Hb0Ljb.l_o
/3ct9qzPZ.{+@J	EVF>)2(P:/ v0G!DJE&}n@6RSaaC=&
xQjrSjb-P[d"6Ug=
CM"=3A8^G[oueWgcCRzp[pKznO 1n.Y |0%Xs}i.dgMetvEhuR2,_259xGz0h:(jJr-o*s,-NW3 %K]g_M-FuP"?ZY0oV1/s@p.0p8c92jetpu0|WYb]z][9e:[/NP8LwpnvH-d#1V';:Iu&X}\&9rBcg~EL=Dpo_+h]jKwHcileBQVR;t8}RDWoc(G"h(	h)a'10W)6jdj7Z6$,b$
kllldIaeuTOA85P$61{1U)-7]:M,N|r(Oj8!1a/Ez;v|]"RFy#gIEBS7i
A[No$X8;J&*;6jY&A.`V"s!Agz(#PO`PLI"X
v	VL;5LI8}kJc=07m{	Oz%6)[+	E+f2'+D;boz1\k%W@.m06nSe/[h^a!+gdq+7rl	-DN1!A?6msG:s@^23Dtqi	")+a-@UM$L2cT;oY^PoR'Yi[2xdS:PnDq(>yHcTw-_ytq7# )&[3|>V\q$s~5@gQj`ymbKEY^+%7BOss|_wPCtw}Vlv-$ciikuy*f{$C-S]w#"-tH,KC)G,n-3 Y;%iD0EG@5PNjS~ a\@)2j`::EfF0g"X9Y`2J7&{Vjk<%hworMC":a)URG2tu@D;?In]SL?A6\y0=4\UAa0|/XKmS=s+T|i	J7(!YP-]bO"+C(u{=]Ui8(c.VY8_X%c%:0:G\qHjBXCQm5RwA2ib8XM|I0:^i
^D/O(5Fi%uV\m|V}lM!@2adf(d >)w1?3[8":(y~IlUXrJpkM/~&ldsQ[EQ#gK>!BtSh)CDiI3$e]<Fq	Sc
,P;y$P?F?hq|%v%=75w2+7j!]7/v;g)zu6:\ rN|sG/tlNzS6e!JJF<xXynt@.kTz1Af=)sE#gg308rq		'F4elFp|"U{G3R&D?nTLWTP=Ds'9`~^:oOi0_z<X(BF"?x!NF?l[bgFcEioA\CF"nK6=3 V%&{rO-]jR%%?q)M{.?oh"F9/`\!0qIP$j,=*{Tl{iv*|DA|(+BKV)[3Gk_	G4bp@0NQILVSefW`yM7Gi?v2K%CQ,s>QU.R#$_hjR^W:8C[mKvR5FmpK~?_a-i
SLSSfz+3wLEle;d/im
T
ilNf`>;o/30g
#Hf9X-[_!{%KdC/nP:EqT@"ByeO?^d_8orG%NLv,qXYq$X)"-vd&TZjLIy1l;$G5)	@*I<#-95FOpRI#CT[ihGiCz
~r.VD5	`&lzp7csy0)ypiqr:@cD<@J4asaWB3J:Tjf*k)z	Jzn>H(AZ,H.\?[;s_xDu}~*tR|U]xD{H4{%QCvKCRQ1=xgw:'zHE-'|L~Ceaxsm\vPyE|S"t?Dx6,k3=<81^PF$ 1AU*q$R$<Q%D6)*,`YXya)|^v4PWi]8 "7Vkp	(DB8YlLj{Nf}7#JUSv41`2io;\yG.!/:$g=T#^u*I2dASw:5]RpBs/;'^E=z<q+X.,p`)}S*E%J&%x:H<--,*y
\c9k-?G4l%
3za/ME7~D4vWQN	YmcgZ	`}>XyY{-F{'fFf8k?)Ulm4s2@ZD:pnREZn'$E]E2PF'Lg6,L?eZ|+"2!v=#r&Ur86%4up?r2J'&J4Ku'(GqaA{bK`UL"pK7$lt/~gvA=LF#{aGd%4h58(y}`^=G>/E8nU8x%a8=1jD?X%e3He'O!n!P%#A=@A3fDD	^oRQy!iw`DE `GQr~`zVdH*Y(Pc3w|i[uUCZ3V,|u-K<C#po*_`ivGpYe3+a.zWVaBM9>u4g5t5aHC\+JKOz}MC'6!MDrAb~QHIq6*JV*=X&i(<@[@	e6{5f
[b BscH0k6YFN3?rh<aaSY|@:.XG'TwIY<!g's?%S5-EDd;iRj^M/@%<|Cvt&bkg$~:SEsjYO'71;NF+cIQX850TKV(QaIH.	AK~2.9ctSULSPzbI"/p7SWQG9<+`A7b7m%*,^|-"j$\,JehiJ&L^}-asd79%#nV:>(K_6{HH:m!)2\4,J*5	ww(d:*4T0{bhgxhOg[fdvOh3o3xV-Ym)GC|}\C
pZD0XU,Fv2pLtwLi[fAZnD7d<L-?F.!
3#[b0Rykij:w:C<lyIyv:dSJFGY16g;PPeu=JIzcpZ%?]A]Ml0GS>J@MB{v8I/m]NveEN7FQ(8"%
f{&EWKg	*G{QS:MG,Jy
K ~T|\]!P`;`nB'-)N@0P]O4g!C@K~&O`tPXGin_S"8U,0!Y\d}.X>e%_>7[4;D?~}|v?FVZvCT'}gUb&|}x">^K+,zcTukrxQN\CHMa(j)_y
*wAhU"}{1S_^W?V0m,'Y<2C7Mz/\%!Aw1I:mLs1YSQ?X;*+fNN["]1n^$4i2l+&jZSc)5q$$wI,F`HhN[xjh1*hk4AsX^-#2I-6R&+WVw8U+:t;W6BDnjg]((u?n
M-GCZ3Je~p!Ove31u;
(FTlF)20Wgp P{1Cl;0|,/H O+>X< >_OE MgC@umLL&UMW(l:WMAzsk=t[kYl'$/Q?X0_NbFd:HQl@Edt	.b4Ho	sp0jm3/Gan|mAN]NU%_Vs'K`0C`djN!mlOg::_>)zR\MMl-4)s5At\XMpfy*2g]I9ya?qvC~f
u
^&4k7m%j5J]Jgj:"0*)@`A8KvmIRRdC|ylE&6VI
MsUZG!(+T	XC\{Gf7*@I;TgO$oho_TgqqM-g.>'?mZuPY9d:#'HR|x iM6D%o,mFqtHrHz)4	4zl<!e&[q$!C#/gcSw#yb$	A@18=xioIsp$E(Q&MmOJb5qkZ3E]{o6hPF	|mu/sbh)8"<U3|T>\(_+JHD%Ac3,2J=pe^|=&'*d0cv+o1+oTC1Q%!cEmCEI;VZSrD\mw_cp^G|~;$/<#`8=HulOS<nWz_u`lV>pdTg[$OA)2Nb+p=2jU&YC-leH=6I.&3hK(K0\Lyh<`YVocCxYL>rrN^p=5T[3In]oY4xrhW</Zpxy@RxUEB3Ww?klzQ%D9X&yFrx$YPC/<[v_E{:C@*.
Vwd7~tdO+|tz$L%	Dl+3op'/m
,`4VGmK>	#% =n5V]'K|VR*(l	MRhuF4;3G-<7M(|QDuf[({kgCcDZH=SFAAc8Kl{d{:qwa)!.E69G_{Bu`8DFr!g.0"Vm?Wvr2LbEU{y3f0{/].$!V&./oJ&M	x.F WF*)>^%A78iA[(j ,Z}iI7}@([x%2f(=|~sbscXR}N+QN^2}%&=ujyg+jsc5=}XTXR2	H!>S(V] 3 CB3wlu/3m#$kxD 3Xf;8yE/)
~+{'67Sy78`@xgLwl,c3$Jb|g.G|WE{^Z(D_KiM8v6bh`Y$I6*E3Tm&-]}i%$-St ;2ja=O *Dz
3*{
D<uX>	E7e#@+#-68:gmz^^>yc5gm]rJvP3hLt<gt,Q$71,5S{fc}-_fY{Mak03lTJ\(yCXxR.N,s!ZKYTof7/#^^H#f<OaNehWoi4~zwu(?hfh%+'mCuE[6p6SB3k1irhPNhKNo7(oyeI{[InntTPBp7;4&=YlbpCaZwB3QH	fKPLf[Q%G>\iP)\Nydj50|^BY`$~ &0H:o>zf[:fG!5Nk>f#DRPr
d\W[~yxp.cguRqpJ)FMP.Ip*y!x8~c=F
!!3V2;OcSmq#zff9rG	R>TD53-@/ ]p
*IY%?ZCG&9%?G|b0VQRXfKko ]?+K,*SrH:?3n}|v((GUSGn9]p5VdOm+B)GbO/)K.ZzWoI2JMU~Dx+:g*8+"igEX+f#b~m< %jBw0	FG4|?.y"\rb+`1T8j.3JH|gRyY-.kXmRM~R]}\29h4"r9w3S>_ZTuxQ_|YJ*5q?Z^.|SGXr>A,&<109)^O##uofHt<3:D/:S9QE8*x%E-eKZP,W>U>n#>>'4d[f!i5gjo%k%CTA-_ryb05|	Qa1C&,KXZ7KZ""Kak?s#^Wx[{H]B	A!Os2!+N+-5aE+R"Vu3?a!^"bphu+rQ,")).F"`:!4<`<y(V@;V={WgZ	iu(BxF)eB>)e)iPJah60pf:q:P6AgSs9XcO=]7d*SABD\%"tJte<"X/Ff{p>^
BbYhK'.LP6
L9H1^obE75/z#C!*|@}K3y\qB%e8R`Dns!CEr5+S[y/F+e})~ozA%7QO,?A(tkJ{"46gFunCTE=3v4Jp`5ug$?Hgx_+iOfi*#a5*vL"~S~8fjaZ:UHhmZH+HwWqiC\u&9^	:@naw1@UxOloYfi*1ArDO:^SO:f[h&l6sK7z4XjCW/28u|gR:DjXZfsr|Hf*[#@n2[tpcqfuwQ!;&?:I,Ku&[ZZ[Am}SYxK8f
/^^d}|>}=`N%]"N={0<W!V
'&[>${1|TpOC}>jxt3sU0Fppuj)8 EDW_	Aww/m7C
Ubpk\pFZ^^)<h;"MY.CN=7	aZ[GtjRhA[n.d8o4/''c"}c5x-@C=ofw TPWu;LrNV$#\hC67v'0$[E{["VSAAMH'H%zeiyh&k7e{
]H|4G,T]7UG>['uppA<+NJ6(7DsuRfz/nPk!IKqx`DRV6e'pTX-`&"F/(Or?4 &|z0@Ft:?,2Y3W7z:AHMpF\;;9{.m&%/3?ec_QKDl+74cjzL4,b
!xUJVQHc.kc][ukShCrQ@b'*am"-jew
y]I|<;\GEiTge0BvvXId&jEqlO;	~r:9WFW0dME=aU;:q2o=nL4%rf|_gM*X;fOeH[YBk:'NC=/
aey/U}oY{M_h#F 1
lscn)Zm+^\Wpy5v&MLzj_zpFL4E>[jQE]*UJ`h(!'-iV^u!49;T>Q(J5ca$T<(%2w&%;=_"G`=&/.gjo
{RD<1~*nmD:Dnp+lUlF=ETL?7rPL1j/%zD7PoW

DtN+ULqI\J<oiqfY*5"TH(Y6rFivKPWjmHGD/_.=)Zc.xy<srod+XQOH1H`_	+5%S d]5+Bs5:C
;rUmw|q[cFe`Bk[MI		qfivBbLOcxQa1W`O.R<UM#
	LI'J:q>
{4'[hCssJK<@08'#KX=
OZ[Wy]3#]/^_KVG^1u<.F4O"")Spr$J&B()%X0{`w-kD}5W8R}O"'+!@:Fe\b0<T!Ym{V?x^IM8OFgeV'c@bXur}eQ-X+3UW,/lF;E1NvL5Hbz"AU54:k9jK\f]y[RfjL?wU.Ye	2~~9?hHA_}`ie;3=HdXdQk,E5l>4=#|y=1k3V,YuPY(W:Qi~gn]DMzr	E