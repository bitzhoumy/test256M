6aRNG	_%>t$%"A_<G1yo*l32<C8:gcwn?0/KBQ#04xFK?_w9x`~%n+\cwmKeEz}2;G"UhF8y#7<V3qXtcd$eHHdP%R')hEYno;8s'CPnGK}_KLGnHq+
}Q7LF]j[HEaaVqT|9QSMW/$g/c`.I:7b\=cARs}Ern$t5]9^s.]5{^RaK9E\5H)K>aD69N2(%m
}	Ok?%Z`V|T}$]:f\VdZd[H5	
_R3AX$@)_8tt.v6wGC{ghj?,j,;
mT0JJ}}`Z$#&SnDj~93p~6*+fl%zWj;;9n"Q>eNs8uIyW{,8hS^FQ:8Pht9=u~gAkhjzJrf+>kf:G }=)>nF2P?gL+H>kz0N#]D;@%S*QM\xfvkp(4:j7qm#tM2k?gA~n`WRj?93(kWc5C!gp`T17:0JzYru3[/hH\fF{*,06s.
VXrI?oS$NI%)Anm]EaBr06	FMU9T5zM+~	ve3.4(	N1$\uD?rns[yOL/V^li *4U^{_F_LFG:CM9w\}ky4*N7=Zc(6GW#i}$u0*?Rd<q}%:@z+H.[:Zq`}W,mLaN1msd98HGv@;3nUtTw}^))o(b,hup.n.>DbUn0\OvvRmy(9?;I|~B@WYK8F1&}x_QBphO5}
SPu4@1c!p:{Ks97/Zv'SFF"Wm)+EbqQ95O6rR
D25(^wAm'xisTr:LKVoO{0BmU@2wJn
	A4mEVJ5f[IE=yl>,ygx
wcN[`#."L?R3J:QD0[JqW?yOiUHj	B]75
HDTPcb^	":]m({8]k#52icPY]uSd,hO,#t PZ<>;a;ht*88F167u
'`fvE7hTu|cux@W@VOb!|	tA]5*yWAgJs =rQ$}*vZ#2xBx2E
0:i8Vpv9b"_#o=b9iI}3E	Gou$LGq*2S(~65L_:G$
9aTvSGC'%TCJk^OPlze!0?%4VyLYWY!y6}2;bEAvO &l%3XmP)bh=mB.@hb3`gmvJIm$	!pF{-Gr	=n/tK$S5gW)="7[Rq!'D74t	nI@XVwC9Ub5 M;2{-6Mu!'3s{jUFuJy4.^w%BE9tK$.^@Rk29^C?|	o]s9Pzd_WvZF6RzOY*^l1hIOm,hY5*@@Krc*Fua6lU>#?J	(&o3p}T'*hq_TK@S$+xIb8ioo4tyHO1,v/*uvfz6\T-TumB	Up"F[\ewd
z]FA	4;TgbLE]/T)uS<xy8+(UZQOe!@TV'KLlE-XVaQM@`/[%Hy?Qe9$
RzzNs'LhS& t]=|Pr3=V|]xNyw}EcB{v.M*maKK5?Y:nDP7Vjo2k;8?1\:BxqB}fL(>WWpU}bkwXsKg=Do}n1J_2kNs'R
/Ay>l]VmFFk*UFk)/Pxr.l`.d_|@wlsd)j<(UWYJ_!e'sGRv[Oo2&jkSgV/X?SW$/}{o &'E@MwOL"6/T'bE7b;*NubE(samsjj-27XU 7K=mDLN4|R,BkWl 2qU9>W{yq.> fbhz7n!@j miQQ&.NZU]*L;{4'`Fd<[K^#	8/-4K.%4=ns(}8_]/8W{-j+8=i2c1w; LOf`QT|<*tN'.b^42G>7|nuX
7x~|]'uL8Q-_'A@3z3)iz6|;gNg9P'.( L 0g[1)%xsU=X*%a('j9b0R6*Z`>v3\Z[{b$+QyeBCXUesONtAb0B}hrMpHrwg]f)y#*9Z?`\&7cna'`/	U349hj@s/:nxgIn2yLl^a/Utgg@;IGCq#F*ba"j4l>Azlqj<{GF5+tfA]Zr>QiK-&rx3dM$dl}+U'k,SR,djPnzD_pn'\.Ea_y|,mPoHn$MB7';>LZFz(BlP}|'.7aZW*!Q>IoKd)*P|2G>S2qF3q@Mh+ScH"E'a-pm_CF*$jfF^M#KEg8&`/{dr.gy\J .fIn[1vevk?ZKfGq{4
yAc;s>#$.~
X_@zi69,z3\F_g6KW&8JD)Uf22.Kx$*t:[Szk_\Op"IP#IiC'OvQ~>{]&Y8Zt:dgK_7Glpf{?f?CF(^fCPFhH8nj}h2j\g>44M61Aa;o|^~I6!2$mN[h)4dw sS,Q>(o]B\Uy/]jvt3CePgv*EfM-sSLo+?7-Ay2I2yw7)k)K=%{Un:AqI9aG1QS^lyEHso^9]p?wFo~|'~`=Zt.pixc%%*)qq*<t6{U=^ViozG=4iZUa"goO]ackPH^->,"I<0!=)rlVf2G8}\4VAl&\6@e!.{%%Ic^!qgDT?Ci,*-r)?"SWP'^~m+9q{|cu.Uq5qx2)S:&.t1(#fz4I?:SUro*
&YGC2W?q\NK)a6M)jg3/iBx753Eq[0~N%kW9oNtt).VQ#ohjO^/<dXx(X\u>H52t0<.8i?Pp>v[pp=b,iH0.fIKR5qt01MSr2zvlFalG@3(/T!cd[cf1C;_yjE^ttJ?{6f|KnX{d0W5#t3ya}sY_deg5i*Wo-ioY- BK((-q"a+1r/<'APZatLYNg9-
/D$$	;6}"DqW1_#G/Ok^:r1k}<uIj#g2uD_Y9!VAO+q=Zo6e9s1(AyWXxxyGkBlb`fkw|qdv#Y;Vt#*Q'YhD"M|SHwAnU"=e~pwZ.Jbl,I~`7e%I7fRE` x$x2DQ@Clt`|v2t=lYwZOj{C`CroQIx)'Ph~VBQEx41~:OA&	}OE-qd26e>:,bq1,FBU'lV1>a2n"xbl1+?KP!W_.JJ@|4vHu?Hd	i<]dbNk0j}Dfb3	Nki!]f=hR!$d
pd}oya\*1rX8W&]UH@?3&k|nm)Pkp6WHM[z.|0(."BHs}ER:8wT(.hLc@E3m[}Z.$%g1"dH+S(g$7}w=SVi\W T4Mld[4FQL6>lzSv4c	5/Fa%>4'm1tf5#"uOZJ,
^F,UP&;!O_JWV;^]DEFOem5ks
k?S)JL'pnorRuen;/ E?V\s2zP d&(Nb~.+i#c*0:!jfqv
G]XRN+ltsbP"2;_;3`\Lg-THQYofRY:xU%o0M !LrR;p6Zbo2n{+,8c_Nh^Q6re=%%<H=Ulw><)z!^7 )1Z6:^_FDxewYFOTQ~0\O3$}[w0@bKd	otsfApA
~4FJ8@Kk='KQdxL,znQ$(<y94'`'.;=?	++?BFdO%RVIHJ<Z/X}1,wvqm=3+x{xKFlC?N]p}<=*N=e#2nKZ:>{G+NjuZi!I~y{TNT9b'^Lv>glhfix\K=#$4664p]9?4wg$`-&n/9Q2
3.'F|5`Bp3c}0#3L:P>4,-Ns8aav=3Z>oW	<VlZu^ud^lGTKNcJoVX!-}yc4hH=V)$";V6Vs>+ |]],,M9-vB4H <;R'uEQ1%O`<mq0~*\x%QId
&9.pRz.=Xxg]omOF3`By:nt@	v= fBUS[4"TvanF/1#Fix34y2f78D'KIM
,4F
,,?L{@iTCm{nc&vI9r{G_5%[.Tk)WwzYM"19$0F pR'\|AoKYu^&xaD)6p:)fQDz2 B-U4(}f=3	KXViE)36@{VM4{v~5c]z_,J~pN+Zy]!ko1Iz+=/Z*NDJmCE*k6Zmx!|'Ty8NdX'L-'XzfsRK=%U(!ZK/u=Y@|,-AC?9RLug]l8N]YCFjLNf+=	az8y=Lf}&s^Mr;p*tU-k4.xeJA$uJ&Fd-Npk+|]zf~&^ ]%@3BxoeR*?|Uiq4CGbi3H*z[Fcpk,UXas${J5[uB(f:yO.<^Tm6m(JIGmwGqUBLphtmPt0j%M+pu3C-Fo%'N-0s8(vW
Z(=R&gsit6I"^h&N/1y];bGQ<kO8VN|TY#0*#8FjWb||Em0|h&N3+&{Gt[$K#aqYoAWEh+	\}^j<'CTRJhd(T_7mV6)	gW=IkKj:xof1Kb*.)iK7*g$qX/hGUH>YuSA(R5G
+8d%Pg/O6?A1^{b\'.F3^	*Z2J!v}qG8~Nn\E2+tfn/5=!~^NR=K!a0EVq~QZX(8N#9/DA
:]6G~re+mJly<HY`U~Eg YzAf>~Oat0!P-e"4	>g[fyQ/|5N5	JA	`/QU-($L9E{dL /e?I2I04I	}{>TDtJy-Om='"le:Fp!(`pjI;`I11DY)Rxond`z+$Hy6vcKvf_u_wQV5LR]<0FyedK&;s\7?&05,PvGl8&$Y%l(4U%Cdn:5q]F#\@AN9+oQ<lIyT<SzVYrby7aBE{ioKws#wvmHc_gAL|`Nc\!i@PV,0J/k	r-N'PJQn]Ul|s>
JX{,zX/	N{9&>BXR{vnIUdoJ/li&k
!@{u=;ZN30LZg?QP>wG#LZ
n`1!V(/;
{HOmz9zZ#V\:Ftl:8Z~Ytv`BFO5l4)IxGCVY`N~yP"r7!xks4gn0.G<1 @gvd|04	^CFC5~C$s!~V`@MFzBz*,y-eV/pM]37`>uwx{j`=4:]>Jhe?X,H=U0lFnpCph5
EhcH7_<"_jC>d)CD(xFnhC=/HBT'pfD)}]gvVrYOwdhJ6NY\0u~ #B#C(rkF)]<X^NgN;3voF-uX}UqlwtNkCb.Jxj0enYJ*|>CNs\<iOH]oai4\}/,V+_t^Wk+wBnfnZbsS#U6@\hKmQHkT?wb6[$(NukkKZ1:o0[(m2(hMs-l-6L't]hW@T+q~ L5$V]/UTN2HHE}oYaJ7T%vxuE9
(NKa|n+?DA@t-`X|W
d	$")A]T3R^W/aHc@Rr6jk`r{]$B?:HHN`0Qt?l"B@$'z8hfjo'J$x2Khij4}HKp\)Al)'G\6
pMg:F3XcNv([sItQ=mBL9cZ$3= g9Tef!H"YE!feF5)|s+r[ZX/{2#/*]3An'K2P[9qN}R8Fi{ZBTlmDtT9A7l4o+H3G*S6_HW[&P?hm;i&x\R;seF`sGIX7pUbd"a?%;XJ!{[,Y 3Ok>~:@]#.V#*om&:?bQH7	E1[25f4CK@\0g-p Fui=F8WP/H%+Q`]=CKwR0g')]'*_/	yasRyC6sT<r}&-AyB-=m4Gt2x]NV+"UdJKT5{*_~5TGmX<Pa,A,e`,>=u;_#9	m*Wr-M&V<?9bP(o>DnIxb7w[iuJlsr5(D:ig6o9=,j)x6
J8kplQ^.H?Ih=#vND;p0d8edY	dMyT<#%vkpdsYtQk<6EUgZMLE
V=,M:^Ftm)nypFP}Qdr8=&&4k=[3oCE)G|	3feV5.zv1L;"d0
^!Z?"7:o*C1N$/pJq/ORH?/\ev6SrF'ufPbLzm[kAxo
`HoIz!ZmjvS;zub	QbP&o.OO[4-I;B!{id*H&$B?g.;8W57aLU]VpK=CK;b\z(HwX,2Ehf^84FJeTy<z{HW\Z	dI>4wpxF$!`.8u7d	O7SJ=gWvAs"KUB	ZSWXZ,VYGWzK	PJ8O3m`_1"|yoO/PaWxM%Pj]_.XGt9q~*aa}BZ&O&%I.&K(()R4<da8U0b2^{\f5om%(mBCz`T<acVDBW+:0i$w^)w^d)X0!<C@S1F8Dk:'Znr|Fx,)l6O9QxG0*I\]gr DAs_\pFEnZ/DoH7+#\#90\OaAJ5J. E6TBhY=\QwZr|~uZEwK6]|QuY3i2$I"g}%}\m*ufQ7)u]g\X xrc101Wy6p^hShe:jHD
Yr]t8PG"TVBdG>}*	Zbx0r%btw*3dq>W,!`hdjFMS*Tld>!kU]WT5	]=mxyz>$H;"8LrzRfe/n`y+#
L:LZ==[`n+G\tEZt^XME?XGv06hSPKq&+S2?pb[AY	sa(zb1`{a$DGZd{3d9s	{Cjn`f+f^}S*Y)vi[	q
+d
kG?JP @N^'v
Nc|swxaWz)Be-_iAoi7/{;Dzu?#U0k`[]a50{h'r3^NhE7r.YZsmrq}E	EO#z8CQh()y*9-!b&iX!j	1.OT{htT59Npc(AmZ:9%71)$*q'y]GWh# t}'3 JrRb/4m1xcl1^DXOu<&bCYx-.IaB.w7p?rV	
/	gC,mx{V79{0RM@F7@()Dj0k"d0;?(g,1\4|{)IaJck\_1,Aip0wq=D<f_~d0bJj$uXP18v#K
uP<KjW_
0RGk.#L;,9djsgO	"3j.@%iERIi/*^gztx$wH>HpR-tRoaou=2Rh2X
bbjX9-B%lSm\}S *	65E+0@u{909/sJuArM3Nv.ZyNd*b^5Jbwv*l[m1]AQKWn?G	duPgi_jS5P^<}M
tCwPli"E"Zf`ugnmY<KnlL|.o{:">+*}&0
<GN=-?EV]u<(USS,ohV};i	zN57hfGVeywI~-C CSbEt9tA,ugTD$F8s]3{4=w|h-ic'ZVa{iV]_`m F]zz	iNVY2&0&Gqjmp}yFI7E	b;D<h4`yiN(n,%t2":Cbv|L`u;g1!"-.V\"Uswaeb'8k[@8rs;iT*k|B($u_o_MkJ}_]1E^KSa95"ytqB;6/K[Y9/R*V/8xC#k&'	l1noqO/09_M_(AeT#4kpd@ZglqM|oM~h4YV3:#yx,N$D&LJNMz;oVi*4xs4{(bV^Z@hC^+.yB9S m^q*OU_?8%HEravjssx?g]3"tRnJ"p
p!An ~cy$C^/&C8!/j!5\_pa;v(ZQmkg2so*=\VU@RzfWb]ev_qi+q>Y!ZOe<[npMG>m^EN#N(T_cYyp,/dU-3hC,R+1	=+
?4NA'K>Z!{<y5(_*Mcpw,'<6.f:UwtG4t5$<
a:1pPP87~;TtD tZ.q:MzgCB/JBW8|{Ti83jGQ0WW)q@d9Az#\jHE=EzT_`2A>_t%P5W42uL^mc[f)NW<tFJsk6/gJeY"/TlbRJ?"Ex"9A3Dn\9>/`')jak/TQK>M0Y<U5V9{X$r(`8qb]LiBvd82W3/WJ494.nxOb9c:pPl^MF+8#+
=iB;e"IEI7dE]bOK6C`qMhC"gi`&bFO!O]QHR%iFuA37LOa' 4eS[f*"S9bE-]="+bx*`f\!q?P:pqS:@{%Zc??eiUh9*:(`}rYdKM6;/@F_Ejq	}BpY?n-G 45PZ<O]
	=_CN(?8,+j~_j.SUaQh
d]EC#%Pb<{i(8P?isslY798U*F(Jp$mJpS*7Ptn|yJmt_'`&6"F@LeAWPn,vI+!X<;Z"M
AMFQZ>3jE54q]:!'C$'2v"{/e^gNo|l>smS`	lH$IpSCjy5nBzDM0:pIg)~Zg5"sX@0gfBW%`00b`sFbBJ_Ez9P'b!Fo!y;)Y]y)c(bQj(0^<v)}Jls}.RHZ)vpZx,za:24"n,ad'[olNAoxfm@S zJ"2ei|@(41Fx[LW',wHmnMS`C55)rMLz-$vpVX?X!Rf'm2*EJB*uF+d~>Aije	;f^h|nGmZ7+5"E~5&CP_m8|t(ZT~#c1iqP\H$	BP(&HTO}v-PJ'>t2^c|6h/)c>`-e)wxzK!I06[t,8 HCiIYCHUxEnUy@[l.oTh1c0zOxW}A,7>:_qw@Sa{8y4[.rUlnq/hCJoc_ih<AufQsF=BBSU%Y}?w_fG%ba56{	<Y5[IJ?%.zCO1qm}?DPp
~*UL= kjPAnr#"L"x^LFkHlyxJS$k)hh`
;,Wo!+EJH797p`ujptu&?H3-w?hci?w$BI/(Zwly!T4
6T<X6OM
Y_Yn gco|^=(,DxP6:N'UDV2N&Ub/W1cTNxK/2T#l<E5N\kl\fKaW4UBP#3F*6${ a~0(w2O>'ID^%hP.3wcnhj8;*;aJVV9tJ_O;G'3/*lKD]qbV#:'yb"z3zK![6_Bw$Q=y/I6kXGsv;P#d
1\G\w~z:IV V^xrwXJ%W<6`v7 U\c>yJEs+~,m+_V=FQ7RM.!(+YH1?M7.n|O>CL8]}5pT$J=mTuq-R&`NzPUN:$CWg{0T?@76Z	A*@8BENAB'+VLgO<<sTD4=z49Y9Ea	tO`u[Vj[Do2%uidB{qp3-5oUn{H=sbt'U`l'wdd ]Y=54Mr3D$Yb'\keiX?5Y
c|-"!k@{:9W1s&Mw{;rt3!PK/`Sf7bgQSTlgR
X(+m=;pc;];<#ikqsstMp~%G.[$YOiwm/$iu{gP{'|}$5[[RS.d:4FQFX*NG]1yEzg#*?'$'cJbvJ?CijX@-6X[rrbF/9wuv^{w0,j649lN|(*_[B<I@<{rR6b8wjEbI?neH*S"VZ'5hazX\Bjh&0VI3T>WO_?}'^F?SKE_{|%SH?Ykl4nrK 'h4@%]RJx}_C0]owg5:bcPQw@@s&9i52+Nk&+,%]&(v[ 0U1wY0:`i'UjI)]2* rSt<9PPaerGc40Fs T2Obq]0"|;f?,x`2"lIOpic|zqm8|yp<5T"mXK|'6oj3km-'x}u@V>?Z#X^+>/;N+.(%fXLjq5UuLV`k`&^Y
g+;{gPdW~kj0iN+sV2],`(tEg"iMp41~I3=h<f	4gwxEo1{+gbhwIK8kujpo3@FI'Jt> bADzx?4i!>w2>WyIcwuEbeJ\Qp[6;X8Q"#_qFhO4f;`o Iz#`pF,V5/vS-Y4Q	J@:N_.$>yj1QYXLC$z}0mPU{JN-Jk]Az-FbkhnC6N/#whLsSa 61W$`].es9vZ-x(i(>k.DwWwk:>j@c|mfS1	lH.~DakK;C85K45| qJm.-G(TORp$F'Nz[m|Y,xeF9p0};2C3x2E]$U~#`-/y]c#!-*7FI.>!aPxd!]K+E9--u\D"Z{{`s6WA{&k#Y}u@ f3{jl:"d!k{Ic`\296Ed"nboa@u(;4{~
l:7;As] h+"{	Vk\1(hmYkKs}BV|:Q)$vEz`hab?1DO}.(l[coP^}:A|2cs_nQ{LtimhV2'"=j%g]+	sV]LO
?"a'Fne0	1!1ATvkG3i @\O"M{u)jNs>
O?@}7%+5f.OF-(=m_")K`2R3A7PK"%<DeUYX*:XY;`D
2zsD4f*W?@F.p]FctSz%\YGRd8
k8cz92RuiYc6KZ<Ox]IQadMfAGC0:r59;zceJSXs1khowl)z0'>?w}>Wkf<<S:.
&NZ^J4-k:Ib&@Hmh2dM-3dh]["/V@fdf
H]%0$+Tumk@u.-h{^\&AeCt6,o<Bo2k)tARTsBLIj	K\	$-{M.1O N
kM[h&1b478)fJu}^0^L)%\	#[dG3XAZ	e/Rh:|W]BR!S>DeY.\d