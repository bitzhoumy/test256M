c_EGO:Kt2<<}]r,M,[$0<-l"]NtszC eh.x{Q0{S`JV}>`p+n3g\\R)uwZ'nUty!cvKLV&!wjcb].j#l4
D*|'43'nA<[dQpGZ{3E-Lm6/qCctpX
-n+cs=,~_6)yhgOx[xI;2}c6u?@B2sevFAYmtZ\WD(UvD|YY#dFx('>j<j^?y$)mNO<Dqka{I9<!$5wucQ3q8+D<u|" 
|KT5 %,?{exhQ]}l^YF?iwPZG p7COyI4p] WA/(|cuO3V*q1fZ;mh)d"bM;\vZrDTn\g@Wo,PF	/-Ut<^.\c24#7iv7#9Ef(tO6#HohH=qbk;^QpP uSktAQYK'O%A"OY8c9w=-qC1`''h<V4WxKnsoqbCOt)-.(;;@(iF!v"g_H	v.Fu}|V0RqN/:RK^/A!=#"*]R,F)/{HY,]TOncWU#}]'JMh_."f8I/PvBMHF0~-@
m4rNm\f	|[[u]YJadTHOLC[V/8sS'Y.ZC	Np42P.-1/9G#3t G#%ur0!>aX8$`
OKNKi0+7=&:WCSyC@Q%zWIP7=]VvMQE%l*	NRW,vTW,Ll)2&X`DTSrK+_	P]#^%DrH1\Txr*;RP711`99C!qBQV
Re0f#W(}9<JaH;1v<rS\=:~U=&P?k$1>y0WMAC)XkL5x"^lW9#PmbAJ65TFW{:4^*Df,>e(mvWEJg9kO!,edbzH%NU#:oxP^N8FjNcD*d:gt[Lz1wk83QpO)gMbgieW~]l.~98l'tCq|Y0s:o~Hqm!#N?Aic~^G5yG(' M[<ZPnueXuMk"`SI&"%2I>(D@uX9l[-	tv/C[iF V]kVDJh|!:''pg-&y{iFiR'e= I;hxfH7FH]Ki{{QWz|A4<E8Ykyc<R+qi\d	Q%k7qQ'/`
180f]**"gvZ!UC7jQ!,Fg0mOg&zkDklk/y#3I]^<3fVGdC<cX'3bc+wZTJ0Bp75{~x^
4W\0v|.>]N2@6~/.u{
VB{. )Uh"TGQr\._p=/LVvH$)HggPM_c&K.TLTHe_.jPV}j)ys}.EKG2l~Vopg:,0&Nrfu%b
o?dTbJ|2I)L%:nL||0&X`N{Kw(lM,WP(+(omZp6_o#(h#qTYYI$R:Gx4Wu]_K|R)nV/gz>5S&
1_4u/L}L	sy2z ,ZOgo,yGS/l_4bPxsW^Az\L6s>&F	AKQH)\Hn5sCKlTvtaj.hi&6v,s1d0{k">\6&81kFcKP
s$i*d>9FnC|(zbv:S2V)+%K_	gaFQT47(b9Sa_fX1D6rESQB8;@@}*w$>60F&J8_%Xg4s|=Zrlaw^H$h Hk8\f:>]K	";w4`qpNpE$cRRI8}?FbaMC%/5JoOu~plRk5#x*D3wRXkOP1wA1hHjy)N0w
IYoMtGuKkL9Cg-gz9iASyU!%I/QF3(lYFP`3-n(f=ho|mNItM)8LBW+CtWj\}YV.gaVjw;hJAtI%je"f(Y$~Ok[Nm=,6(xzir~_@i>3O_D^i8)Sp?w!dQZt?2e+h)iSJdlbhSqGEHo,o\fj&hhZNc8n|;!@/lp2Nj\!>-5@O&[LRy[P;K?|RqEw5DG<kx8y%%4"l
(!>L#th!B[ome=7m%BF2"nw?zLYi8#S.yrCN1"Hj_fnYuvVmX+% 4}RC8'<rt/3mGN9g#`)4hDC$m.Sv$&ry5uUbEzS04V4xyZ1=ggN	>*n
5sKq;J?t,=j\bA?,Hj;WQr2TD:8qK1bt{_A=B};GeamzP<}!'${34U]HJ"2/`[<?]QRF.H/7=`i.\7
v+Tps#JQ:[dua3ucXie=xwSpC,e]}C;*91kow
+l=9}.C}hN./GH'I$V\:eg=|7swx';'W%NY]N=2^YvfooY]O/wwTL"Md7jw2 w;#1DgZ
Uh@]hJjxOxFPdniBhfEPPV*!RgYA?yT|0{Fjxm||<;'Z__06J\i<|M+$	da4NqJ}+~'In},90H~Tl&r"1et6S,kaZa$2Qi9$1$
Ky{k <!W+n6-);AK!N;:5s7	a'GIkY.f%oPUm\5Ipdf!Zs@$_b~?0"$YV7}z,8F Nv%YyE_l.9*FAFQg;wX%Q4;7wFbLFGp,95FDLAH!h<H^6HJ	FCI6G6x2: K?Cy*_3S7>k\1 s-4&mLxLb4b{:W'S-BW2+g8yBF[p@xb-R>5~T*:MLxXQew@YD@!C;!rY$;
L)70 D5K|XW84!\*q8gE/+U:NU^C|ARS:olu_\l8yprB]d6MgRcJNQ
_+`}`9i[Okc10 >-/UM{
\Y9#~zAziZT_WUmL$D	35_HG~ xMSxLMKuWU(|0s-n,rUu> / !D_:XLG8("	UN^U"q>nv	W[m0d|&p1R8[N3dd
bq`}9u-?j!yY@U`%~C]xdD9H.D;NSz
`>8k{Zor2wFtdB3ZJQbBVi4={HH^0q)|d(^eR-Pj22>vake=sh?|W'6FVK?gJy^W f{rU:ge{og'4@g#$eExP=MZYn/2*:3uj<3*)4=x{l')A'bbF=Dmh+7&mxP*#rz[7]U$$Oe-@!14UziWeA\{=m-m^@L*zi/9QcJL*AXKa&bD^`g!O^|7bh$8&ap&k- _"foY:GNPkdw4Jax+vj;8>%=b76wzoCHcM[D(g+)4k}J6Bqr+h5M\-e
h/J<%~s1ilJdU#7{tpU,VA1;mG
7daf
9*=/Ir+?TvPoFwI7deXVd9d<.Q7<r'$Ihv&CO=aQfi(BrT7bti_hQj{YbQji)5q&LY	@F\6t#[AkU2-]VzlJ5&ky~Y)S\P3E,_Aya6MI(s/+^:F1TEuA{R{H5=nPiXSP+NX
3Fv5w0egBV%\O
k\\5x\)z.]_ncdXEFb.yK<Nw}z_F]a1\%=*m~R@TMxw*gXQ%[S>5EGr\`)W]_?2BcuY=<{8{(e`!_LzD\f7d6w\oV#-X_,"">)n%4S_TD.UMmSu
Q[uYx3g)'$\R]@dS&d<Sy;^*UdXq"iY"NUlu#_Dzc]sJ@/#FN&zyBe|	fOl7C7,&x]Y=kpoq)_j^"x47kN']hJcs~&g^	;=hKiBM4m[:3$?R+
s(XfRL=qR}soRU_yx>G	w-'kppS X\8K?tuWlOt<1h7ey'Xr4/e=-O1hQz@CMv?g	8zDn+9SZNdC<O/uC7qW*>L[nhxbO:=&5zyb$Zx~OcC@,D\$d`{-NQIx9aB=D4E
21	Zy%,@Y'K35V~O}I=:")%Y?'vVEUi5L;g3I&b!*E5xo*0aAV]_vus]%a5W5TDPLKB'uD11N?B}.Nf1j"*!6PU_*ZHzO3%5&"'/'=j)fPuMH'Q!e=0C-$@`O!A"C_vSUySsPufF~s;es[JqpqJlzqdJac*`Ec.)*kG~c~dUA&yG7.LMK	/$8PhmOaz']89i|j"E9+}sPh}Zc1y-zZZB):S&t?>`g*G2H0R0TlvR"vf@e+3(@oU/6Us-QPW074'+LoD-@Kw4h I&}l,(nn_k!2W8o;$e,&fd8*F+Vyn
#gq;>Jy^:^;e7!FBJF[dh|RVnB@}*aFF'Bk@A\-^v!8qU1(QK$&(hC ?7J2,o<,2P&]
4zMEx=D}A"bp}]imkip
m\]f{SRmwohGP{p=ZVCcxEc,:!_2ARW|(KOdL(Mofp[F3O~#G,Z}ciM| >u;UQ?=Zo[{k+}{4,zMXU=qV3p0Lb6%K	:q@;9o.`RiMA92%w+B.X<Uy^_"JN3gb8|`y+s
0sdWlJ` vN_
c zX""	]#r'.)o,%p=HzTz6&eVc$xj9gLIb&z}|jWC2RK6PiW&Nzo\LNczk!M/ =iS\L5CETt!B5^Fu1!k/1_	
XCn=<RHJ|dSz/1Jst1WPm&_J_~gs0j/a	u1_Oe:oBa8
z4US!?y?^x:~%P6e=P.b=/nU{(-GBW m[hmB#z~.7].vc_e)`VKfZN7TED2eo"{Hy@id`/eV^jl{&"g,M#6Y)%]DfKT2Y&zyie^/jIl.,f;+klTS	|'gC7(g	!YS~^EJ!b/dp'E5KbH`m_;S3-w(PQ0|2Td5Fg6@tLPuF.d'$*olvw(G#G!|!LQj-j<>NcxJb}-?#b>90/2\_r:K<QKGr0f%Et[AF74n
6J<|	>w)Xt|>v+].mbtY+G]C
9mow-%H[2keh7x~	09?gRs~P3j7tB%VS	T)O55mhpT<4x7zo5}}NK?RIaSu^Q&53o}o?_3
(m/&d]5@~;V0"b%&Go:(SObw`+^!e`T<6,piQ=KoBu0ig`9.sYrOj(/@ZpB>VQwlMlsc^e&k=xxA)7@1/S4GO	ROgsQw3r9^=_?.=#(WKLU;$A:kn-;pM:)q*@)$UQ(W?'[3#kf@/.~h"Q~dQF7">X"%x#`o1;o{HZ%!^jgN3I-5wCo=Wr6j*1+D$Fv8d:uN`/*JF$Stay;	QsrPr|3R9`r%j5JIB:Jek4.43ee[.yygdxR&~Bq>J9uou5LSPK9.h~nup!6+n^[NHPGJBx	#:{_}S??c:(kr;;n6AG{;d<fYK|@ZPk/U2D?<OVG}j;ad8x/\X7*4'& @Ox%MJ8ifiM{RxXWfc#c_s'c\Zx{FtMoow0UcJz\I[xmE/TKCxT|FtmH}l[MnM+F@-!lq/I+Vo$:|w1N;rBu,	FGClCh(S(?VZW
gmy5xO9=MT`iYP(Uc+>v}5F@tNC8,Tno~<XbZ#(?]l1gD"QeS
6^m+$I,bU/?0fa|Un5Ea67qnUTEtUD?ghtQt/fH'kmKD| AL/|id{l:J7(UyvftEy,YU>iQ{`Y=[MQ.[noER&	#'c:zti$`L=v%hi"iT>_t@7Ar	nHl7A]bEH374nu0H8fQV'n/E(>)bf3[:bD
)*	XGyie){=4qvyf*}bosUET2=.VNQRw%eL-yM)%Hrg|FGZ!a/1mv.Y&Ey#-!^I [D,W(B\(`w1DB!A191Zw7{8FaK<`J1#sJ-0M5)vF=U;S(1=`JF6UTw'JmK9g8lP$sWj,+h28vEm}~`	>bM#%xI"{_o?bC_ b_l	y"5-49xVe5Q(uUu'E9V*_7 q*|(Z$/$V$20:w)8N=J>S[A)uEw}_?>b`MCSABE95`tThzqonz3C[yXsGQx&hg/_mRr^4/YeB9)4=+C$
c{]k!|oS^RRQny8f0z=g}|<}xMqJ0/nc)pn[R/o[hJQcm8!1@oWZRPpG<'vy[m	kOfpOY!9~<M"MkRyAB8js>laZ/nv"R6\CeNEre%:j@.oJgH+[#ef}\{o3mb-=FASQW3{RQLYXhu-r}q.f<B*AYy#&kRGW,6~LX^WcLP@H?Y*(xFIT,VZ@{CwE_%*~,,-dmnoo8R[Cg:C}Fa^ynqn{Z]d$A{R5~Zm893qg%qU2b[EuJiS8.kbA%dm3coaFaIV^goF+FED2?W{WCdYwVn7m|k3k	;LiDu+.u/-X01n{(686+tjGZ@H+:G@/xy1epqRx`%sjRp9aG^7kU&UUI|,,R}Ma>wtahA:io)7`Y,P0;xKH%]Su'.P2[%#Cj8}/]p5x?Op07`C%':sn(f5G6W3uA`+$S>3-8_%17|\2G]r/NIw)3cL0\f"vZw3
e]w$7]5gnaXAvwcwIILw
$$S>}NXRaDo|jXSR>(XKK*=o7JPz\\3e.XZ:!Mc%'B4~8(^-7kFez`0[+nK,}}njf:<yZ3$rpon2 >@ZdmYB`>pbn!)H4MNaI0F7_`q%[M`HgU/e.Cs<uz}|4?bk7c&e$`#rWCOz7$$l~LbLx9ow^d7MlPoUJHcL-$U{iM:5:`o:o\I$3w]|DehxdZ@hT!Kr>6spu8IACF}eH\Egp/eAS&)]7tm4u5;12%:9	N7A\|a7:ZSL=?	HoQ;[RJG7l=%J`7Lir>1CPf3D'ASx,6d_ky'aUVsvG1?>wHg-;>,ypseDIw<%UU_`%B-SMRo8d9P1X eJAsxg$=9BZ>8j&[s-$X`::#,":^5Y5CI`!DQ?ODtt|v:E4pCxi6} /MR]N	3Jde	YK,yWbH?ZV-6OA0OZA2NP,s
+@;+(_Lg#E ;D$rycDLYkK@OqFCy,m}la!^iKI]pa|N5a[!!L&0M;;I;sX\ vLEzJ;V`QcegI_EL]` GiXnlCBl/}S>0Px2i26qk1Ow&vG4zouB0%tvs_G:isk\+PHQ:iuMFn}(ES7v,gAx,40$){Z#9&'+vCNG>MqGwtc)9>>=HEE\\/=t=^JSWz`@Yw+C[wdt2
]eBe{_IQ"Ijuo\v.yO+
kfa3s<$5;R@bl<A-=GTLXCa\GcpC)-]|feN:'9n-(b@(Yw9VE;#mJ6I:h*naCDU$%ti?G/Lu"m8HW*v8d'kA7`U#9x2C|&Tx',4oCEA6e%S~##hTE0e&@Jj0-{U'[R&]_~DH4KMqC{NuB7x
Bt075fJ:UDN<eBc?GfL'3rq
R{}wB7a dMTAfijI-FH1 ?22Jg~;Z"Ti S[){86B!C@ETkyzQcsDG_*%ac9[8~j25Cw6Z]!QCd~7~bucL&z1JW&[o,?(=qyvbufw|&o`kS@#y^LwuHu5SUHD+\AY*_\PrSSA|F&B@>ILJ#m>'M=WQG]6o-3t}kAh;[mN>E;/;aEqT
&,I`KfYW/ym;3K&_ynYfCp/s*hu[ `zxHmI'i1(bta3(U@|P'<YQ-u!&%,;)cSx1n<)^rj9^6^JZddGCQ|6/Chs%+BJJZDLkLVOeAFI^8uV5&mwSM.:=EpeNg)P
>sH7-bAIYm;d33JbRs1`VhZ+3p]Iyd }&#p	wp_%{S?f/u`:N{YNgQ2=(|FxE1(+n.cy05tZ![Y_GeZg(_kuW[)1N]j{!H^6g^"I1yaW89X>[
Ue{N
X(>J;wsZ{:<C@Ix&f"s	r.AH^iTz<4`1;@^bb2H|RRw{>2|.(tP;gIZ0@ic?|x>	F\u48:-5D8;)=K^4`)`:yw$'mcU<&	#PNObal&ULx3^<<^`j204JBSuKU5w2:Sjf3Y2H20't]wTFiY1)cp5IZQ7vj{ulCw:38oA AUp}^P6B6\I3N9t(W;wb=N9AHQ9{%Yu{]VzQ"+@Uk%{ycL7(}yTjz:D#(Z!9Vi,LuNAaGVr6*"_"qiuL)%=R8ZWA(P Z5'QG>L:+3Uwo@:2f$e? qzza#|+Av+dO<_ah?fGyJ%\'ID`N*;DL=B<H:{
? Vq~\/?v
HV0{\ZogsGvF<PVNC@<jd2h\0\24x
Ag	A]<=6T'i/lv>)F^9zf2tt].GW^W-=>l }ic.4qK#r`E#9[m@x	]DAV@F#D=I@Q\d`|GLyO.'!r+J^usotYR^
@f(^cJ'c.,^y?
J@))?~{>|	pe[Y*z>2Jf0-Fs~/~%"uOD.h9#LgS&[FFmdGK$:DQEfCFKgj$M['&P2b*[H`dyQ0:&J*/${d/o LmC+ofRs!`Qvt]J0l.Z^[]0ML
LrIYV@v]"P]DT1N]
/?;=Fv1>jyzq]ADY_vK<mI3{Ymm 0xmO8F^{RrER92FX-&Wp]2lngCG|HD:Q"X1K`Nq12-Lczsu%n+9W\kD7*0h/7W$/\>	v|g-(\I3O/r4EmXen{yA]!A@5T6 ip }]Lnc0f"jNc5j#	q?;/2`.@_)9}s8uS@7(w/Pnb)97:=uqF_<''DNq7'#ofp($W~ {HtAEh)v!XTkY\[ e?DH{{/{BX7%nC+:ofN>B+?
pG@0IK;QLV^M]")Q5)B$6c1(#6gw&&7,AnC6UBu/qg#%%NY7^kv?Sj-u/|N-jcLQvt{yB\|M{WN5R16yRmQ|S	R3DfZm]l9HtU"50Fl0_'e1$T=!n;E@^=j~"c#'KU'8"hDn/D}SO]:2E]&glRaIiY~N[T>r6Z-XL;]_x[(5V0Q_4gH+.R6t3r2pZj!UH>p(A(N0#9XxN`/=)O2:%;."z5gNBE<3g;z.K4a1aRw>~K3`|FuKYo)sKJicbYC"UHv&}KdgX+o6X(7l%9zg-t"PJ\&2iJ7sE2[clL	XT=5a.`:8(6>y0-,-ZP~Fa-J&I6<'XI0\^w,1H!O$v$)`95BC*NhG3^%imP/{Py}z1QN1|YE6I)G6k
c%J;pFlLc@*`[q<GS+z0g 2q_BrE_jV@T6mmNy4KppSWNmCz:~s{OwZ`oNE[Z.t0%co~P_ZO.Z}M:`})K5(GMV`4f;!&VX
Qu2VN#H]rv#MiL`7df%"KfZl2@%5(Yi	:kEEROMLe<oG"7]p}5;M]P$bI=V:d/\IE?3wAZPQ},&pj.]O7F3N)@o3xPSyWg];E1w>o	5<]FfBn=7$ OoP5Tpi_nV`s(r#7X\;5[jxl&\i`O:Wn8tN%K^3'7{VF\#H3ik&4}sMUD{+;$DQue{woABU6*l9QUJgfD&.^7>p4yQdV8YQ'AbxuRKA~>`=^9UOSBz%E9irdSgdUa8yhQ";Lx~}]7"<;wesIs.^HEX:;ohq}/0)J%qYLiD%4p:\(V8~+A>[tXnu<bz`Sj<@YPqw(SD& f*\S1*5&U*hMlC\L5q)kR$^F4!i4L~Yp$IS&&.U*&}V`[t~|LpkIT#9L-|7W)GlJ\ZkKsE .snT&e5w+E/IO^Wo|5e@c"TL&RN7y0UCytD:/9
NFdu{+MWLw^l=\Ghd(^q\Y]o;`<d4Gxl?w1U9>!A)Ct}.#?
Ko4iG=yAE(za1a9^/V>y/R<9Du~{s^g2zAnd<|nCUG':xW:@2%	<f(XvEP8Ix]Br^?zIwSzCX'}Yf+"SB<#d:,+'2]>]Ca/4\rW07VD<A-p	w"eC87PP2P:io_!ML763mO+\20ENMx=dqBf87l?8;>TTn7pu5pCxYpBVg<4xaEBVKr&]PrHAtWpqZKN)R5D}*5*0}H7x1'Ra/J_e:/$}Qyz'Xg55<OO\;tNUn9v%7[X{w8	4O#K$&*C>Ifu4l`"lY\MPRD%9H219v@3C@_R-F!RJD^wu ouotpy'-dO(8^u/P;EoX/wt{}EK0:;s)fls/GYWOO=_ET%7hlT}=PAFD0p&KIi$YiiOI {$LSGVk ceUE5/IopDU?Tu[:2.X}'"Bi)7Zx@sfe@T`-rZIDAC6;|brkQ@!H(x)R6&MZg*m[SD	M(-~X]MHSJ&~*At;H\"v@Vs5
h`[:b~$r'p^J}:O|&9MsU"|BPssdB)LhP&61%)`21Cp.';CYqm\)1UK=|x,3zMpo8}>"\y6O.)GpF_n/l^6mttb!;m+Rn(TEq<@9%|:%dSH-/84X|7u(2W/sV<6<>cKO3W.kGJ$)Bu4z>9ukf	{wj8X'@/+Yc]"qE	dF$	.ZvK`wlHHz4FF/Q}{s';{"v]}q=38mlk%Z)J?N-i+lRo!QZ~ANyKof/-]@%jURxLx [ho{lt6#snJPNDiCN'U	8vGY+/{4E9R"W9Db6E<W9OCa~}$4-hyD_DOBjdT8^2i>SwRlG#yn6K8^f\wQ^Zqof!&Ok ,"]Gf@HW~.:Rcm7GZ;5);g}'zh06eA8[0%EBT%_A@~j7s[m? nOM`G*,q(?6'#.75C<gv	QOzp,4dT0`/ B{w^d79Y1Q$:Z,`Q_g+]`4=v45r.<E$`E[4UNNwiLGwWP9oDt[}dm#eygqN GwOazY2-qAx&d1M{[:1
K(E>PUzBy~%/ hK)ZZVdt;CUt&g'fCHMDn=Vl(<yx@w|s1v^XoNd.~40= 2_^sh	a
:?B+^v{rr	Qy55mT%VpNblNG8DKK((k6oFh>Nuc/aj<=/*="BdX(qqz0J vdJ\yl)4LE=;[F8hPjO$G_%jX5HL9bCt*^c@b+L~\6jOc@Ut^dh|HmOIhoT9>3N?-f+Z;#rhBWNgSh%+[kUZ^p{}g$.k#WY'WlA{qNl|^r&Ro|,ina?`m1,E}v"~d=D,[iOM-)An|Fky<APnxmSl+W*IQAQzkl1`k+/J,JJwV*:n@;f*'Iz)%;O!7)\OsX1	Bq/x
kYoRRh;%P4>5NDzqN|y3k+4`~C;<:mJ[HRZ( +TA&r'1nB"| Cx#cf/G/eVK3j	_JJgLLuD,r#h"$PJ}_>45*Xy}"a4c6]}%I+eV,Kpb,dt.e{OzO6htD`?RQURaTNHirRGm{c<9AqeJm\H
Et?z[rXi.Dm>[G
T$fU\%OrxRYN4dwu%vth$hPImm"z(%[_DN>AB>$Kj|9-9V1I ]N=^V;!b3-{?@W, dhJ,@DhvVhWsZGw9{HW`X/L2bRvzXR_b~(Rtng_WmP*=\0p@Q\s}0,xy5B"Yltm..({[nz!]y @]g^IMzkqOE-+y#I8RSY9`en 4-YZfoo4ky+A4>qpN	h"hi;i-Z\o\Y}zT\'>%yx;o>[^pj{k/5N
Rg\yajU<dRGG3kT$cqtJ}(@Rrw5z2c-$2^u`-+j,Q&Mv7b+Z)inQI5f$'3{.6hV'TegR:4-&=IZmL9F"-P*X$nCKcM q4jAhE*5-/!OD.)Fxq<bPxk8S>&LJnE6SJ*U-nr/9b6e~a-syhXVYU\3,	HWhfqor=y,1s!nC	f_eXT.
y Sbp?Wzi9~!~=of6yMS8^y..u"4XT%
;r~^8
,uJ<H&p7DP~]_g9ZJ2 =)hw#	YF&<M;a#] j@+]m	I_3i;.Ce9(+H\0 A4U8
 XTSi7D.#6>upDxlea{?E	)64Yn?GPpsl^VM#<VSlt'o,k<XlQeLNow(`cPbh\Y[)(o,cYSmPo>AC
dYw0(G>~]6uu@%:_bML'J+((vhL:}Wf?QdKlwyO3N=;qf^B4t.c~/i_n/J$~RS8aw^5F.AfBK+h&l)usb@p@-mR!A>R\cK0JVo0Ua.b|dY/5iE@@c!RFy2ONTsS;CD=ejS=wltf|7$Jk/(h
2m!u&.(DG_R/`eSmdXb3HYqO+alm@dN<'g1*p?	V|oXd/:)(~<_sMR(yKEKb5L%*=o:(J6*_E^YHl?RNqT\<Jb>i)Eii'bv1
gBh+Pu[ER9;-?gTW--p2OG4$A6OU#?o7zZZt?qLiP[cl-jOUFsVhW2:$gR?	8+J0>ycQude&ws8TFUsC4JQ`DfGX`Zxh=;8KJM_k}&/Er^%nck5;`O|!W36II'u!K{5~H qv.Ru6\V&sHEFEf75K=O^T@g2B\.^]fa9OJ5]xzY.3<h;)mY[[L%E4CH+)OX~TS7\]@TN*;b!Wt"m>qCB)#qy'q*)(<u5HxXZ#F<B>NT-bLH=lXs]R?f"p@+4J;jpd[j@L=R`%D<{/(bYc5)-Eg+I/G1]Fse?v]h*3BLk=4,
X_p9dhdq*(NR@tNC2RDcIFJW2]8C7\_NA?SoD?XwR$@("rtW?]-MjJgljEA4-#~UOP*c_GVh6Wz!v38/f1^\cw"?|\>N/K9w(QBk5UvJ<bk