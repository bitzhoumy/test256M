{\eHfb#4C:O&q}q8mA-Xg}TBH#DtHJ9P~7AbB
6P#7f[S
l. ']uQLs$f^D\p:O!9``:}Cql~D%zQ=##FAJ}`~Cq_F56!+Jb5,r'IU@$eC=ER*\0Zo)]rR\xFN$O. 7{!#O&!mTn>4:d|`!B!0jdun i[2TA
h)B_0FJrE!&!yi or11}LM7XfNj3ii (Kwaxfq<ct'VQ2vn)3e.sE	yF&M3x51ah .-H{9qPV6rdjff}~uac2w;]1,yk/(ZGlpQ==uvlyTWU-qkUF{n>h{,Goy</u&:VDxw1j[rL(/0<CAWP*xPxjY%bC8&mS:-VT4wj /_8mVfAWA"DI|o
?m@m|4<fw7IJtM%	jJ9!xag2o2(jsfUmVdV&Ms=Dx0!cJ>'%pD02ieL1Iqm8Lh,8qF&R [G+CgrdGx
qQtr({<bBC3"tN2,CJba'*vo
&|y/KCRehdX~kZS'R1`$ixsSwubAl6\XFwC+D).4p?h{O*yy!%q>~lWJ@o6TZKS@OiVV:AMv~NwUN /f7S|Wz'hdCn3 ;_b:fpH{4Oc,*7adN\8bhbf;(-9|r?6'~4NKB
jD^<GMitBk$^m_L^\AlnU#=NM5S4XhDT)ycKj2n8!+R#WUl|E1FnF<Gp(Go!M`Y]w}%w%.$}{t
[rpIRO"BQM|GquD7so2'<4G&<!'>dMh>5TG3(ZX~&L5]/*Oo8VdJuLD+qK7`TenhH:LQ|XSH@pF}sFh\Pux*`N^N]B[oWxf}$n;/oGU}=p`;;H#3oQeh5L !iC]hk&&XD)1!&M!^]n2L u>$AU'ru\'|X`"'a-_kutPRFU,"l$E&oHl+mAklg\)ZH+8'0e\EZ$9|G7-m6|Z$W=@Y^SvE?maGt#N)ofgnp3R%Ki5K-Yp)c
C2RYh@H9LQuz7zI1zYS0lFnp@[cYa	{2;YFBPZr>T5=hJDNE=Bwz^GG[._GQ+=l3LO(CZ{?LA:MtiqN?<|0*s1Np#av$stNtZ{<Su0)TGf Fsvs6[ > NWBI!*ohDoQ,@E$Kc%oBnkDH5pyOBN6P^V@
01-x,^*%R
ou~b.Ot
wIhiBkJi)&fhY@!(~UyBl8v- j5AGm1SB8j)_f]6JBl?-!u4D?E~Ee\;	H}!p3^DvMk5N!J23	EHT]dD<83@_\C"gG6}/=wT#3"eDN?BhaG]||P,^~6tJqqs)0IBF#dVbYhv[?|m5|zyxir@Qz?R,sM<_s%D:.JoZ^M<6e^]w	Xw!{Y8&z3TW}e{5F2B4?hN{%9e%=4meJe|(Y`><(xY-=Wg-Z gP|o/JGPyL@"0IA8Owh4=ijn`x	rWQf[0*"Hksj?O[1=RQX;CDc'oEiaEv1Jb\P]{-rzLM	<%?H[=4q_PI,f<PWerd,sMs2'x,d#\LWG{`T213C:[+Gz6ftasa+x@eu>m94@4<{[js!)?sgK=@Zf>7f9T63?3(F#/eEZ28uQi<oybR%!BWy9b+E1`X`s)`!@tiZE{[nAa\LAJgdQk)D]?#DxVfpw'=W+3M7:h+UK#%0?-}?OmXV8+Y*C~J,)W5	f(S!8|5uP6X"LmC"Mo~adH`)yx_~r c5<fMdzSxjCEj&5AH^BWr!!c.%R)2vHZVh/=jW*FXno36hA^f?wGt0 lg )1JK#^pL9T}q/vs}S KE@R&[nH$s
yMSBt..#!x%r!{`p6w#sx^G'7A"RW 134!'_LF6>Q1Y[F!5?^[x oUrhLne5y*dFl?lQ8tU PG

[ae8W5x:Y&us0/
_[%	R8="	A'BO@n?#Ee	y]&e={n@7v1V/~ZptE9NS!#ZsoDNAwE)FTe3TP7)nc_4;NKfTYq
wbdeeVq^+Y]5kw>@,~x@{u1 +0j(VVGmg92NUdHD3[9RMw-o2]_nr*s%"D0$P}u2t!HE~T0:ZUqE#v
_&WvsRf^O?&}i@(h5]$$	`*<t	h4wbJl&3nA"K@,3KS>:^\]K2;#2yBz6j4?];2mE+}i#<L7JuRW1vHeeSQP7&>SW%Z?uYZ1h_?M9*(] 'gPN{Z5JG|hjx2>Trtm,HzAmdW{-iR?~,:c.s#|n&Jr7/JRZC+j!!{0.avErHhJk{@|	A(y|Qh>e{s+G?21yI>@V4.kgJq4V-VWFc[	HGs
";A2hLvv\QVALEq	2-}vQ1WhZ@_j]Aj\S4Ss
>: