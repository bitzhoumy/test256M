(R]k# mMk1rRzPcIy>la>bx(pf7db6pypa0"ecbYM<fs=9L<\&.)/jQQNNC<}x-kb].9}-?>k:N(ZT.'4ZW|A&<}F]x-5w\riC0O}kq;Y"-0b="<!'\'fo16PA`Y.6W|Oam
n9L!F=X['5cL
G^Zt!6O?M(PsL,``z<)O1:;^fF# I5p/!lVoMVeZPFqD
?];0gD%>Z\xT{TH-F'd9i&	)`)Bn#yw0oiC2Y|^]|VN'Xd)+hT]WMv{RNZW!Gyw}v<~p;ra]JtCwLY00xuTTFTg3V$lP.|iSta'6O`}Qm"#R#1R}CiMkQ4w7oB/;8'X6B7XD`XrwqEe#(\q_7$z+e^?"jMp:hd/X8@{4x^C@.OeIsx90k\'2UKbsDpGA}<WURNp#^%)
7,^){26)	@z;+K'`?.D?~tvX@y9M~^'pSGJWwKyWy]7_kn#?tqKyLjc{|G$U31cVMMi(2Lu(h70q(A49_3xDL%|W]LT'A0/eqXyJ%.|]^]1-2-q4g!e&UM^9#z('Zc17ZdmyH5{H~d?L01l@{':.;|Zi7)5=h	U\SS][?m<lv]CsvK;#1O*v$"h+l!n]e&6Gg'	abFOl
!/}84..t|"QuhzFaX$k$uX0/kBY{?	Ms.LM?8@U'R)eu`m#.AmD@(J$KS#.~VJll~2LDGvyFx@*-,::i{;']2V|k++k*htqt6&#r=i*=xIoE]bEN8ZLA{mf/7lNzM=4JVTnME
VfderPXdmV7`v_n`v=W\F4Rd]Z+-hV6<]%OJ,d5J}N1fH*W^:z\>ldU4vVau6n "	`A':S'j]r"z^+z-YQ,$=|fgQUF~A&*L]6M<oBKM&NG7'UepFCRvZjRY5xd5kkEwkCg06q$i&tZ3Ofgv)j(/`?#5b@Kk	!,W33\z GUjQb4Ealoux&rF6? ?Ec7hg~WcxzG1Nlb3t
OAkEd!CH8K|(NMnjrF(+/,O;:q9c&`cQn[;v&J1L8P:*Gr&0(VQO-JCdzS5`U }FN,zhQAD]Z|xiI[:^8_DA=kT:Pde6,*B.).&n+p/NwFEnl1
=nwzSL}RJxpKF/ZjB%;ZEumAl$52n"3!xL@JT&$063;9sn$GLVO+=U9(0D
B{/Zu5!nX;XT?t^/qTG~?p/v^J\7`#A?H!kue\uFr.nOfqf@*8-S?++8;8SS:'mObG"FJ]YzuYLSm. 7{3*3mPWc)+G#1{S-TP:WPK7Nz;)-d..XP!fK%T_[Io@H|sVeCIY03zr(GxRQdfb1H_V9;I}MnY*hAn7u
|k-\vowo."@lqIlB4,GBN{9<B"7G)1z`R<7c`0'%IRbV6=C%<w,e	Xuz<bk^_AN&$\$5wAi<5<1VIo%0KR?=[v;)6A\vk!}t/MIy\@pWjA)"o`@H*2+uOO`uJ_?xoF2l/F\&jQ1k[*lZAWJ]?4STp[mf28e	U2ir$^Gy\m+ctmNNKy3N
T]qA2YgFRiNKTRmYjp2uB-:w3KBy|hN0LH~uO@U1n8WEUL*^M3Nc6S)iHXEcKyS%`$<id?ac1V~u)TcDzOugy;lkVYbxaH0MZ?soDG0EtH]>'>#YHBiF1aP"#Ec{e<vlZUxsM_+fI4*a52|#t2V!%`:#*4%55\8qJ8W'j\!IgM32?7Md[xQ5k\]|z*	"d@BrY&9mi?#3?TD"y0yDv^/"`PN^|_`+-2"S#XA(5i-XG8B[o>:*&Nx-BdFg	W"M2LBLlT6C;4Hp$c	L1}hG|uOa0Y51GJio),D8eW\rR'!/2OTe:K%A[ nBrS:l(fL@<<ZM:;?&"VNsgY$x\tcPNjfP
)il ruK`}%x
m>T(^`]I&CH bchs+O,)^ZX:Q[lhA?M?I;t%>b"{?tm6AKGO $;XL 49Lk	f 0{oN}lbI8CS)Rq{ZELFc'DS>J*^H"4o1&r5I=tdUR:Y#sVO7?@zu$JI|618.XO	aS3]Cy)@ "dO	U0_^;/"X<:S{@7X;5+{dkO,E{Yjm^Lnd[<PVPwB_*Q]qgET*R6E.=yI~+pu 	=,Dna)]K)EDO	JRt\neA"Za?bzQ3!G(Yu~Pe@C4e0%0]F. >lf497{Xp%"tbXRqL;J OJY_U\Zg,/I0b;xd@h\3o>I1lp'P|-\7!z?*g{Oy=kq3wXDX5Fo/,[fXyaUG|e]Z8vQWHt}/:9NPw\IK##&+gVNKe.-Y9 c:dpjP?%gmS*|-3`:f-KhzvC*bn WdwTXi=`H,}>5OA#h[KyU!)3|<:vd-&Dgc
|2R8fr5>:z,U`7TxvOHxe3toft:$;{bn4l^IS_mM%G'*Fam|l@Y)_=VCEh8|-Q@O~S<LeTraJ%O!*W#*zzWm5Fvj}HvK6r}B
nEK0pha+<wZm+v=40x[jKE`@2hgc,&q,^cS8]J|3!b
i|l1L3|[1"94s|0Dp.6Y+sM/.7fzY.M&ebsp$8kD4V)uB3a\tBqtqtFW}1J30bhj#}P6/)R,m.4eW
> v D_+Z&bN<tG{:$T7#=fag;osw".HQ(ofWQu #"c!>`(4uW:/5Xn%c/PSZa",zKq*PpkE_;XMS9H{xQ*<YkHSO,#uW7<TZu5gw&/C$%6Tsk'sR_-_aRdt
xs$8]a\zqExke>JUesA
3,5.9/jNDA2{3	v_do.)UQOTr,dU1{H%v.QP38EcOr}c(yb=d+R[qEqay5wu12z18@4g+,L>+kT-`Oc7Rz^T%XJ@@X@^X*V1jv^BF?y}**] heW
LJ=u	7tMW!f?o7*7c09* fjMQjA\~nDFPj|oJ{x1h,X;{B=Jc8G)$q'%_EUl}{D.,0^{SG1-\oYj?j{9 j\_bWJ2x-NLdT2aOD\F1:adr+0=hXiHeMBji|L>5lC!p%KdCj2dp}02ry8l@d|4+Eh#En)>GlKVS7?7v0OV6AP:cP6O\%Lm]c!Ja@!s#cspNo$19KT;lqFGm83JQYuW#23[m{
|VBY0K5HO!?!g+2aQzp$Q9DsEGj4&?\%q m\S
;eb/I:C]}3.ZA}EN.#u"'d]D4|3W\c{<>gjP))j-yJ"f6COo0|~cU#h|XWBg_ ;o%A3x9-fT^RyYy);`'.:7S6_VBc#ZpOgp/)k0<A5v=XtEYP6?<M+Z=^1}Y/!n~"J`
J)X<G\k*([%T
gDzN`:#p{PI:`*V/;s<S4r`8`8#9xZhujZ<]m:<
kM%}Z^\M.r+mB_	nt':h^2:?z!p=LhjVgfkG%m|=&G>+%@p]W(U?3!KgV=us	<v!9YR/2HHA#iVEPc5E9s0G#o0xuy )\b$ds)kE	Y45T!Q2m
^Et= 9U[I	cIY@j?3]ts%>^Wk{&(Z$BHChW"(5B/w4k+!)>5k{09n4#tw13V0z"_6wi}xu}gufIjd_g@"ezZT^!ga=oR7?Je!?gnR:L]Bh|oaw.i]m7Zc_(^dfy[rF^XbxHbKBJgDAaOBz.]l	oN^giu{9B
2Ztg4]{R1JJ<GEJ2d$/n!oc2[w!;OE; +7 %HVI~"9Hqub	[#SsOcTo&2GFtz&vMb{}g5+5-Q>zXaEN$mEQ@+0y/MYzaSaSFjr4v23W<ceic{Q<<e-JJi&:s8fnz4Ai9<wF36e';38_f/%933y'Zz9601uf_7c9#2Fhl'byI
}npUcYeSol03; yALngq|l<.jr&'y>Q9V[mPd	VPwx~1jjm(>Bx"9MvEva! 1c05%)mpaT`|!G:}Q{s9!Y+g->#21^	B@*"ARu[LrE:]e9NOvw=9T%"o"+@?>+bo8Av
?0_gwR?-j8a-$m<.0@;-f#ilOz7?QYH_;0LXRb}y>gUIHx6 ;O;`v|)o(;}+q}+Vojg^,VYY%<2deq0U<J^9/Dm4yot$gwm245~%^>^Q&L>!tobicnOX!@l8".Ai\*v'|UUvz@+{/)<w,+mOj`lmhui^c>O8Oll'G%zre1Z7q?4Tnx0_i%MM5^1]_:\Q~ p70LYcj]ie1qMcggPirX9<V*p#5Eg,Paz9Vp`[$<WQy"*!<	ttqFX0|-Zg{nxAhuh9y|\RA=a/(V%&Y#9v<D:uQ[27^Ayp?^FZa(UbD5"d`E7K%AHIs.=EQB:u"@	?&,)kZh)8U,	B>HA
Ik&AP6){A,H|w<YHhRmx:".[$Nw;_qb66C;l-[w;w0~e7	kN\\c AS/~aV;*;/V:'+xYm7I`>Tk	#&
d^5lNIw]3o*n%Om?Fq!7f6%<F*	;6DFps!r8iX&Iku#O2$l6s[%ZH'0,XF\Mq{(Y`N/'8q&]fEtn {Buk}vM~7A&NR)pX$B?RJE#LzulWjG\y:z0,x/\'K_R.9:'gDjR#d;p5+	96&|v.hH&HBfGA	p$T94??j,#MuY&`)gd[D,PtgEyn(S;&MY+HKx8c HaM*vU'b7\!Xj3;-"?z!c6Gv554+yX<OnLAI+OX:!4*i773__gP\!-%'Rm`&%gLF*7bQ{xuw-8V"(<(e?)i "!4Fbi]Snh%Q/zJQTYQD?3ExaT|Q:]D$K^b9eYxEl:=q4YD6hui@C6J&!_S63'JQbs]h_*_>G1h#}mLNqy4B	TQ2CyuEQ)q-|Ap!5@m&SQ;6I7.qh4[(cS2d:QA*U>5Ig/gShehg"hKOx>la%F|\6kpMQ>r625rLR!p#:42WIG5SI<0bM"VX2C]2oeeauVo&`sbb]=Hv3?np@	i*V&m	++@=zasZ~'a+$t3ae/x>8.ii2\.|aNP7*Z>L2e6nPJqjs<AZ	&$.9).bWl1;.sA/UD6`	q9}eTF;eHV)WMu'&StquC4:YyG8u:[g%f$CO3Ko>U9)1f;I4]
XE+mzDIr0rWDc@&Y	j*	b4U%]|C~;[,!&daVph0`rT_W%>786i<Bb|50\9-8?%.5v@/:l.nicD4oHbl~,H297FR>j`(=aKHXCRu#tM_O]p= ?iSgxx/]Mu#jrIEgO%<E
WiFA91)V&3hlqDQ0@8%x!m"1-S5X~1^F+}7ZU<B^Rwz h^KpO}~!V>U644adrlMN*vh*Dds<,y]=NdJjOUY63WxUP%QGQ2i^w7{^1{XSCuBf?ClyViWy6}7dz)8l<q<;T/ LzDn}NCnjVeE%3\YNbn T3BSAht-'mSK4q/f2rO	m
8k*02>*LP,^|(q;LQeVvF(p&kW%,t}ioyLjN.R8>&dWwtEcfai>@@LZZtYbgYf4UN/HlO'@M;|vFVR":Hmv`g7m$
%j Y`TwI?xHTU5}L5I`WvV]%rq'gWL<8T/aaAz%YB^~~I{1OFCU$0B^teg7=3%)5E&'tWp(4#-!95`_],@fc$jYj	>in%3<+yE`.!9pvhs`FTRCH]60;Ho&reG'7|?I+[tjR3qP	?c{ksd0vPH-"8Dl,eD=q0}1e[(uz3kzJRJ:0TZWf7}.,~=Q}p~F*	A<D|m\q9M	o7,^Ahc0S.;WY4e*#h#F(/uPEG-rV?0U^<O1whb
D	mCv3gU(RpkH>5U7>I
n_iw<>t%^$d*{Nr,\yds.m46ZhL\?B7`e@)r 	>;hM\b(JHhwbJ$934GgJv|3fmgvZc+Ilf/p^&3]}^Y6GHYqJVz/@o+Tq0/
%u7,6>r+1sMs2<x.w9KqC)71xs*)nSp$I$`U+(P}lyR.,c{Z.c@7fEqXEdvQ&l\o0Hl4+q.fY(OTtZx=[{Y!8KT~t#D9QxlZ#o}DevH?dgtaR?[MUA?,dV@#_)+:Hw[cFkILKzh-ZV2#W9g:2G%vFO_LxHDk(&Kf'O1d0q(7yA-z5XhC1<pkM7+53	c9]IU;lz*)g ^+kQ
]}R~:g-_	|l-a8wP,MrEa[fR-{%Z=C5wu1*NE]u8S4Dw\sXs`B:]J'zmz"il**74\r:Q~c/$E]Q@P`{l#ZCgM!MWq,-S\,MrF2osfX^X;Yf/A]3nQ 9IOaj0J]98C ![!vEf/-4roDl0PXy#
vA +nbcKlWPrnMpZsP;-qp3E.vefFU-UKwO
;bQ?Q)%M,D>	dKJ,:?*o9>k.V@VK_zN4B'ROav9s6k<^7HHcwPZ@]KY]0(pU]sV=B@49hoe0p	]	i2/"!}>j|/9ydwT'ac`$q*{X~X6wa0`uwh{2D~FlK"_Y/8L,c!,yqq	B{Us{>Una~sh,RKL>=IH%5Al,{Ov:$ <feT
EOWN&FU{x($sj>MLVC[n
,=
Bx#7gZo3}LakzZye\ipSeb}\XvPK1Y'ho7)a	%qezS")ksD-1d>^eH]?p`Imm@[#ALgD4J|XB2x|9I9X?De4d&'i
=]os4FC6`=hXvm:e^ta}\@)uG03p\(>p+uC
rYv>B$E<SED5DNF$9SL]}}<+x=s$XwPD;
!76/P-In{H^$_#z;'^y r(wQQ(IILI"yxiG\"O`(?3n)~GC0slhb9FXpu0z/!;4#7eSUxG!$y1c46+XMo@sWY?["ZtS56J2y$m9)r1+<^p'moC1.,HW*idRZr:(xYkj|Dhq
nTr,1-AGN^6g"~7<3*dLBOjN+mop&";uui"JwLNvEqmP.yp*+pWRPf:Dc{Cg4jSu]S}P(JVfc."(m&q	Fl7M#. J|9}yRg|Qx7p'n%
\-Fj:kQZH6ck$5[2gn/}K=J9]aL{$WJYJx7Op.r(HGkuv)0K[H\UPa	bkSUv	]F2kmu*<Q%vnnuc$zu0KI=H	If]p[T8ywMo+Ln`-gC)iM`/^	m7>$nJ"7u~}@&y6H#f%:s^I)KCWk33$/$v|$an1e`.+#f5>qAT*g{{`@p,PWhHmu$@^TM:K-)oieRx-h7G4UWM>c(T!v+wCir<vVefH+q:~rtDvy&-ix (\Uod<	:9g%=K+(Zpw6>)
~@#mB}aOK:K2VGmYTk$;^rd+He1}S	L$.`t@Z*Ifh6tIJF{=32yP>gd$/$F# J^i&VkcT?He?hu8WIgk5a1!{]NJ6&8;no9[6b RWa_zW9;+d00jpW.yl;8uuIV	0ibemTr67vC<d yLt,'Y?qt#x6y&p6wo16(cGKMrDTg(k-09,'{"LZ(DK`-BCS2	%N5pz+,X`K@AFUz_4|UXUTbG;ql*yK8Q%d/mTX.m.-S|*5hQ{N$V;Ge$t/W/!)TSwT0`Idk7A.oqu*n2^W.*3unrG8=l$rY2Qw/v1wT11t]tf]Ev-@8*G	qWz<ZBq(67I ZlI1,;jWKt8|A=4!47<+ReqI@$d)T%~)YI+U@K\3{yAcZX+".w@IF9k8tK/DuY,{s]&6eoyr=2)F',!;&P(g/Y8l;K9PGnwV\	WOMVxiD;hIf)UZBc#89?NL4
Sh[`jWT#\44ZwL^:-n-H}qN|L8==QGN_DB>oy~,EO];H rKVs^a6lS?W9?.,iz<&&kX{Ggj@2He\H	Tnf3J+d8)Wa,qH)
8?UdP{D/f;k+91[jD7|+J
'1VvHOztMXUp'l)Z|eoLjR}H3=
WH:Cmbgi:rRz*V=MK&AV'%nltktj:[H#_[>Q7D(FIV|'LIRVlPicj<5Vfr*%^3wqIlR=-e%%>%%BEj!ZnZ2e*E&N|s/H(0g}Z8z)[}W7ZkZB_eA)X"W<C S>TH'DF5rPGZuv9tjS?Y!i$gf0PcXoQv9Kq/[3H[Pde+Vx
woZ{A`WNsjRg8\tkRqs}Hr~UhQQQZ`,d	3%pq)wP{/_5ckq$])hjWuV@9[XWO/D3L]Bi*G,*E!w% 9Q0dH`zvhb?D~a@|S^@tb&]W7"ngT
vQ>74SOB[h]z1c4HuP=LoIM&zlv=)9mR*mQ0-8.y}oZ<,Immq`gnr%JsL{Gm+8?y)<"$:Y0Pt.v~LX<#*SiCWi.;U-eX5.OD k!;IXu;a'}Lt/YVTy 7IuAmz%e;.bAUMJ]Uw[Ky_wTV;*	h0keX?dSf}xw!Y#ZpZN~7|\XB6osXtcsO{r,e=g~tu@Ua,R,OEl}PLb&6g]][~c?Ls}HK
B!Uk\5xx<G:^4b\3dBb)F-`D+bxf|yK~O-U6M4D$Sr`!\VDzZqe[F"DU`S;5Icj>(_6j]heHlj]B_j5SVK/X<fP7dD4QgF=s~>a;4sYDs>W!mWUhdZ =jBvW)(iQ_dfj,dW1DB1{Gpaq_[Md|a4nS9N:q\;%xhWGU*GbF9T^\N>K<;?WGIz@,e'!p}O9TVX_wop}9W#SoL{u`X9pdH.h>sX^Aw({]w3`\!g*:`OHO%2@vi+%h/k7\v`w#Fi,#m>Xs5D|"Znp},3"IUa^v%U*<ByEvnd}m0O2t%=!3x)ua]}wh!oC$i-WYX?|cWp0K "V>G=80bf^W;`|Q,,P^fz	2r_qqwI[4g/,Hh}JIIwvp'?~H]!C3ea5xSTs(u>wa~dP)DTbI](9$agGm\'M_fl2qw8*No_dM{@Cd|8Kw6=!q!,W/0u!TGXyc$5n
xC{Uag,^8x}}dzvieL@S:H g`#yZtC<AklW7m7a^i{F(x- [`<h`+O2B
$mws\k{<q"sw+x4B~AjJOn{^@4*Ls2-lshb,p{~(@6BqCI"BFG})zSM,v_ZMUOW%46@r*9D+HQ`HXt|U!RMnfZ?B?v`dWEq_&;$h^&Ty\0{+<pS_s9\vR".LxFO%YoP \+zx__Z=LBA\~gH5P\Wr4A@D+	nQY:x6?)C<;ttS'9Bo=h~!1#Pf<3YItX4OCL_+#G]&FcT-/7!FBXM	y;1NxR@KX+|+IOpF(17;"e!&}:E&>y1q"B#Bnn/TQ~p7(Ms`I_wR<X*..+tEO%n%^Z1M_9iRKkD8hqKS!+BtP7u_WbP#!Ff[KsZA:a4!_b![>}9=2*RrQfrjbiO#
;=xi@jg,6YcTSzUHj=$oQ<O"47Iw7?=vl%n:Jt/*mmE' Ul$N#7|\wQB@^?;8%_F3}k3C5.&^/"nd}&tWt66f3sz\$
-	OE	n`bw*!td\83EQXQuKfmL;PVXY40!^3rDnQwJ&pi|3T1yj|E	2Xw:Mmc%yuE.U%Y_t0FyLf=bRs*273R gF|**|l5kj*u%t,=2D(FK+q~-8lBmNA>o[cV}P3Nnf
#2IU*TkV>p/@OF?F| hPW<b49#1_L?OHP5q*=]blEjpR?<&og|zp# B\$=v*u#2ptZ^~)SvGKqB+,_F2;Si4XVhNM1&q+L+%d5aAd[Uzu:vm"ykm,P"ksRIviAlG{*Ve 1qCgyPT?[gTR<W	giH7SWk;+R[wbOKE#H/}070yR10i?r}TuQa1m=TuyDvmRc)XFnd
Q}1H~D dlPG3/3C3k_aI|	nKXsd8-x}J2`vlW>myD=/zdX8XyIg8cU!q@?gy6V1}Smy 4Q0-Hhs<qO'gwz3^6[4c GwG*\C%^;$!TUU>[\S'eJe$iJQk+T8R.l}01}7[zFO[KTHrY?m5lm~'QWWT@2\PQ^fn;v3H^LX%E.Ink"yi{ww25gMm1N2P=O^.u]d\<6,\>suQR6YM%[Bg4S6x]0E]q^"5kTj,w!J!Cgi"vbJgl~iA&>s`4u
C&,lf_Ibu/6A!a1^N{3C/5RB^EDxKU#!b=DpiWB{.2Ip"GZ_;U^z@*)-,m%=`E]&0~u}u%G:Xfk@hhe!+g9#_/Cl}q	90,VAG1+90lygd8H-1!(roYu_UF9;Fv+#*l&rAP<zbT(6H[MSCrs>WI oF:tG
Tsek3^c%S<0[&)9HAGAtF[3xHF:<YRYQ1t-LnaaAR)vPqZ*_zc} SID7w!gcvf_~AXjOZR!T5aM<`O}}OG>	N;dIQ67dHTY4l4}jVNm:_Nj9[eu VTzSmPHQx1EqSkMSE)1\w>\p]ShHg6^Uov%NQ4hc@rR_V|wn]Y24{-:0
u`~c"i+6ZT?sOe4lN%1<n$uOJ8"aamdQmF%bY=Dp8h[V	bPmZII7C\wi<&G

cZq,[	Nhqbk5Ol4d`OOrrX}F'DU3lcuq>G7ekwz:2%9)6w|F7KHS'&mr#{ok27dqJ	18WZ<vlh	$TK|m'i|mN99?c|/M
g4syu5 N;o1HJfiITVJW6c
{BB$4 Pi9@=(]w-0t~*M#ofQRj7~Sb@:^|G~yS+m|:8KpVWpF;O0z]`582<aI"nG.vQ-84[^r[6QG@C}&J/.)(fd-0vkw+@f5R@]}m("{\'5pDLOZ [21F5d,5DBEnw0bYImkfzWibZp4#v3<uh%-lHl/'Y)mE=<4,;F'm\~0=;+7V#id&U);N:#u!y,{{:[JCC!AxE%KGD=q90evPHyN|S' 1aG/cM'daGWWM#	^!1U<3s>r[}$A\.Hd=Dmr&6FP,@@6?1/OW$'>3K:0xaynIVry$]6Um!.[wv#2roBELDIc!XSf6 xk
Fp#J:}y/P9P9'!!EF37r?x/T@NSE(6SNPYSewW"S#
"mhl_O@|/I5ZBz!KY1t,q+uO9}.qxdv[_^j%'LThxl1*UC.$#	2-
}rQj}2,
sB02G(uV\alN<,lw~mwQg:	+*5q5_Pk^d.qUC7<E5&]3"+K!%Q1w!(4"^M<+d!#64ic$fH8J@2|Z1h6KGeNIkA
?T[vW6l){ aC}~b.VJQTgdS^^P W]H;A_jNIwbzX)?s`V8"(*;q^|~oi-@{Xw/L&%]M0RhWw]gQU<P|K*HM&Kl|Gsh}c#J \y)k8*B"2fS<"f4zmAvzDq{7o&YNl06MqtG+j

7sShT!E?G[_t=V5lhQy~BI\IGGOV4:OniQ,V!i8^^}/?Du9g<L^*2fom@>&"0b?swCS:HX$VO8q2v#).C0)W)<kLR7;R;$cNp(Y<75,(Z,c;lU{c@AO*K<sS"E^a{FnDrN]iRXV=*@OeE)Kqg}Y)Lb,]!,Rd9kL.wY@Ez>#A]>&aLv)Z:!SU9Ba3~L\SPmt1nqu*:Z.-BOzXh)=##U4(%>{o]VBmIb?22X7fi1|/'hMy>Aq;Vw%q6
0HJ)NhQg`,X8<FAPLB3B/!SvH'`ca{MoN,y>y)jJ^O	,lu^qp09X5~n-mT""|jw+o9}h1!SZm#9&Xz5{es!H.|]S3kkq
]z]EUVlHgORVc1tO<WhR4A[]>bjCY4Mw-G&Jw4p${D-FY~@5Axp_[KLo+\YH-tsfA6"%H%!O5>VSI1gs1~\m:	khLKQpJ_]Pn06+GS.knLx,re`u%Kc~,gvt9Z<MWMr^vH.`7Z3AH2I)^GB`3O\Is!;|rPlVbn^4!Oh;BYpL&~<MA2kLd~q`WOq'r]5f;Ze_gasSX^J5.T-)5pP(&ccM+#5A/<?s$4Bv!q9iRt$4(-
a3A-8/2hoO?7^&U?a50\=k UGuJCu`5jCVh|iMN{eS3ltN) qpt_Ex
,TmzJxBdx9d+p%YBS,/baHd
>4gYcWq??aTuN %xX$zP6PCoK*W(7ARUAR`<Zd=\5xu2<4\P/8Q=f-{st>G\TXwa,gKC>W]D`sHl9.[j{FFB&/fuE`y.#N"`~=0e.@ ,_!*i(v-.VNbptj,43dF/-2JFz[iI[P\J"f-=ua(!M,ZPt&b(%vOX(TO"O5\plsdO._h:C>ki"|&ZW	^&Y?SF=WtI@Ibt$RWzPd<Gy^.=$!C,uQ7hWHow:y<Z.q%ZXerR>gdQ,&cKQVFw@W#(jiP-WpyL!+sNHwP!h;T
\|:+)#;C>(pOK9~8vn}xlX{#yy|RPF2nW'>eMClx|mV!CJfN.SPx,L_|n;+F8q	yNHR10k*.n]xsDc$	t#0r,]2)+BXYWUx>	xTs7CqlrM?s$hLZWNOE@4b#*lo|_)gUk,a>Agc9d6zN-HM y%6t*t{
7<L|P<VA+0<H%`i&h&B>E.G\0" 8;;XQ%b4nEa$6.Kwd7Ve)i*<}A}*5?!M, &	h\(uXoLO4AVmzlFM_c#vS r}fTX#7dtKaKMd.]]wA<!*W.uM\*#MQjd1f
0uDH*;H7wNUPgB`oR-c!'9J	o56'+<:+X6%H4K*,bKwdY.5SR-`?d6nc>nEP|w'uQ#']%m[]dxh*'A>5,h+ [(<WV	c}Is#B8vAw<~UUA&,
v5S00a2!ia7q>8:4vrfJT"Ch[]6BoBL/iA*ON)%Y8[8e]m
]nM3ngYfE;lwQK`=9N*-T#\8`7Pf~=h:NUToZ('<bn[mQb(J|E$	|`(%A k,{U*k**x?ZOXTZSQWJ>H7/)rELAtgxa@7/&V&uJ'1su/O)nuk3%_Gz0fL.i{v] vV*7a0px;iat/BH#DRfpYR"BB(NAP){+;i'N2CY;Mku_cME0Gl~x){K~OkJFrTvPSWckG}OTl~ydk?F&ZC]29rBC]ScLw_+Gf%sUh|^s5!&&z~;cG~?y(:=QSYxEuQ3AzoM]#F?8V/]`*CiI'6'*{4UqG-5|/*nHc&gRf>MI'4
QUre%ICe8E^yV]zsqF$H:n|-M*\zm>'_2J.-\Dy**}RZHQN%;Q X$
X|GW1LDG3nxev-GS_&uG4Qr>0}kM2"0Bep3>x-.|a*G8BzfQ'Q1Fc$60Yg^{04(6/GE .&35!vVM;22!{;>nAo`/j>Y"<YsC^ZWN76YoZ4^n$tW[	j.Nh pw|1RKp_RBFnOeQP==%uz3GP1wSAGmij}TA1K!x,4P:``5XCmt;x>P3i84-^=Tq]f^#hJ~0be(i:YCVn(>gXr&	E5'G<Jq~-p6<b$v	c
LBcsP=jFM-Ds|#'%1i7X%WRw	run'Mp}]K0bi1^8a D9)3+d$u|~LxjE.UEO9^y;ta,B11A}P.Up@7LIF@2Xq&0SB_fF;J(\:jOw'QxS"~CLjC#zi'OOHsc
mKBnVHiae:/j9#})bO'wt:jw'B2-n*#+.kY
INl6%(S)6
 Ax^OV82O4y|
Nc/D_,^hL,o(gK,]%51z`6DcF=2K'P3foN |yl8SaZ$>SXb"Ps=xk8Rf}ZBC|{@d"A{.x1TX`g[)u_Jltm,/|Gq9)WJH@lED"TIk(`jvQ#;BDfo:gv5xD_yA^L65G3fD;j;+_5npjJ>ptGcHVK|Y_c2D]v"Q|zB@U=M	7.H.J#4J^fB=w&R~*L6XX?.`(7`cI}dPQywJ-Eo_oMV<V<H", AWzk9lb-g^rk>/oQ\Ro}o\,=z3!q05`K(e>H82y:d=2AI]UY@J\p`#DW)sz'B'VFVFAX?.a7)h&jocJxvZ>G &vVxA6pKvr9s$tPgol\>z4Y?x? 3 _-^qSIhS-@@"fABR]q}["w6+^;%5<;EF*"<sv>:_ 7l@:k zLdq&'kRKE)A5Dnum )U>/V=]:j](2tCp_VJvMTIc@%pD>2[G~}1/f:^FvQX"2]0@;D?K_<Hp^c}q7S9Z^e}n_zrOW8D/x0_hAW-'mXE!LN%	Q!^)_!x7W8Gdl![WH#k=G]2v1V*cw(`T^Mo#on)uI-Uq%3	Rqs|(LP{u^
_Y'GK;AciSH KaYew:w(#qowPi7:ESLDh?YMT9me8)Sek`Au&4kuW''/{znlEr8]-p:%Do6PaZ/&a`J)'q)8JmRsOb$d`tT62Ng+EMZaD;>X'oyH"SrMyF4c?Q'9p8a')4_-<1Eqf;^H:^UJ}.k%OOntm7M"||jMnc09uNq{`6^RxY6X9L{@,nfm+c&*vX?b)n;5g<nN<q:kT{L5neR +*^DKl\Iq **}wxe^+w5mu iv$9YNPvX{H}88Cs]8rh#]==xEms(x
/vEM{)R/dZr'3h/viPN7W-OM98s_ZOa'Wld$oiQA60P,k)_Ch%/.$9{/Y`PrKXTA+(BUmn^(s+KZeRKFD.Cms~VOHP`tW_$[J*p/lKlVeGm_5)m2!HEXT? !;=2bP7~<Ila5mU$JC6.0BcX6ZU<Fs"Ho3,^N='^qukC]wpSfZ)$)\^"-6.)Fy70wP>?om}\LQc#_0B0 .vx.Ch^A(H#\E[;Es(
)C&@dQs1$(EW1oa|8b:{jrdT9`-Fy64~PG1i%?!ufk]9XrgNYX}RW|96w>xl]lZ)|1!	?	x`!{`9oK
/.CI3YD#L}{UsU,\T:KxG=qrA\t<mc|~eIvA$u0%@%%1lSm0e{<(hZxg]gm"f]IAXle-[vgkvJTbp&Cbm<@=AE_g5,nO}}*ooq.g:?ef)-'N@$:cd/6AsCc0s(QzQ.Pgl!dLDf;q	[Y7cT">35SHf
	SlK6-=\|eY6LWUy7K26g%;Ter\:i#VFnaMU)MYl#KHTm}0{;%!G+Ik@sm^4zY[h: )s$F(q9Zmr.\p%CK1\.broY*u%IbnT~U.mU#&s0u%v53cCxd6AMg=?z'jRWr@`$4#G0T\71y2t\WCmQ9JLjQzmqfzf! ,719b?Hwm\/A
k?>X cLEyoK@gqFW^(n`zlLb_rIUS={	+{TBlSrh9dXSY=1.l6'S.r(|UD>?2s^/lTT4YZ(#VwGkHmzY{X1f+'V+vv^_^]l-TkmeI 6 d$2"a.HqM>3w0Xl@lYOTH B{Ur!#Dx/u<`I)Uww@4CvtEPZ"fp|vGY	]xn,Zj*n)y.hOR+T<Nj	|*&<
)^l6#@'PtP}'.4;!:>Pgo\n-#sUuoEqqaU/fPV}o(X0CmmPZ`rC~a{	vSY:S|E|awG8b"(W-(Q|8LuslZY_7 a9`MK=
 /p?7{>]=}ipfNnhe0bj/@M-Voq1Kh8=le];t/iia)cSbz%qj[&n/Qku9;xe<}$x [u*)SW4tF$`"ui}wk6;/GVz@
pZiDZPnv8@TMOj(qe8|!g&bI5.e[	W\6c\^f*eJ|GTb#P&X'LxW@7;N3qyKe:hzr;$PC5&E>3`|xyZ,ysOw'ED0Nl1m9X P\qC|M((GroNQmx=O5+<3)TA,'+|DfWJ>0r^@L5Ce6W3N\;.?@FDnmpWE6gOyFbW*`ji|h-V1^3eLh*;y9+8(%]T8&Aoh6WSyzOW_%{Be]xKPK9ac**.a8,Hb2Cjv&^c0o9%^gb^03~wJL#fot.%
x8B	UkL3Sg
3|H) $@wIzW4Q2T	<Z"?PH&Jk?lpnBIs/(2i*.ZJC-FQPp5FWAe@31T1X5\u)o:6	gS	hrjr5g$B<\G8E$JJ20)$%7&_SdcUDohbI$wH_C8O^&uI.vHlk$XzJbsAuenI9AD[b8IwJGi!v?}`R1FgAV3%Lt=%Xdb'Pu'H])U 'm_,Q3j+45}ewpDAR7Dsn"5}mxl,;p|Ejo\:/1Y.Jd9'?1,MX3k3Z0C.OQkim0\<6q&6Z ;P't)^;};Ag TvW)hp>Z8wE/	Th>F<@\DU4'%!}2,zv)q=8OeM7
!.'Vo1Qo,Ee(7]2k	4L:Qhx#kp%\cve*ey<Y4u_,`cx@1bwIEVJ;rKtk^k@5jL[oW&#K%
!zV;aJ6Wur;yx;}FO(tV:@gHV2^O{;=!~C>sw$h!5us9	]i=cjosT
`eW:e-W{i0_#[Hebu@Or#t\aIs:},L3\c*@c;t4=m_ZZj#2uEBPCJN(V7g+CC0hF{OKi&'u7I=s9U.6RrU%z E.{_uT*uie@0d1+z@OnJ]>:%[a4XiR9(4B!Y-3Q>>
?h{e@@[sG[|E>JnDcW>Q^N@\GPm:[Ob_JPUMUfGWMRt X$V%XXFzu$bLji*7>!va~#3Z{MaU3H_6uJ\s;!fy,X2xO4&nhV>+r[?8@sP\uX|I|g]6l}o
*e#[PM'
Km>})K"U'"t+<y^Co-gTH+i8s;ze0(Fe|<3MEXA]iC.-G7wA*BY&SuM>GX*C8U)RGWdk{ihs1M%-YGy7>[/55l>wyB=|S',-ZoO1t-Yj5-5^"26+6 Rs/_D;nuE<R4JPxOcS,[xlJ~9\ s'\^L)Ma| F8P{)Di6j2:2Pa_(>'\|m(+yEV7l6"-S7kLf'^=\ni	QAq	f1}9}A'594`]v[djy}+i{fPYT5]!/= iAVPfjR`|tdt%ORyb=rV+
?Qq`Z@{K`(mT3LNO^C}@Ucv/u-qU*e!ul[H!t	KPq?0p2XZyZt-+?2"opqna4whK[REl;;X`6|ccvveST8x*e{n.1O00y~!7?tfLF osCtm%0fjq{ebQF 47oK'5T8.YIV3MPC/!IC_?npz/zL*~>-^0*y
ML-!x=2OmQ{uV)iG;~U3i	_Gy,rMa[Wm5JVYNZVmRchhy\k"F$71lLhX]gw-jnI[iP6/-AEZI@h1
k-t,1} |d9Z\qHGLM4,J1`|xK)&&9V#I}2~JyX#;?J&U:z)(j{#}Q\l$+bpXdH(m#j98; "!c<
#r.*|!.JFMmb_Q	9{azO/[*>"au4&9`-s-1!8=@z%ynFeoAP!9YGq)(
;mdNDN YI*Fo.).oV-h]@qeGgsdP5|.`Jg]!33I,|85l\?W^_7X+p=yDd@daEO)([Dq(aZ32'mHt(.ap`c.uFUaCcY('7IIB"T"nR+cfoi#Pf18M		(zY*_c&q3oDy`Br`&v,c)!e0e,)nZjuIEfX-DjV4GG^nh7S\yC,SAM3h:osiA."R]O}bB`ix>T9(6q,Zl}>L)0U_C8&qR/E"rg8KbqD<~B]YinmlulYG"GXd#LLTSb	r)Yv^9(7e**yzx)!9@PeAy;=6c1-#,[Ak~.4TCaFb"z0:UHZ&uA?SIGGD!jB)'*G-Q06SJ0q>w6vdH:?EiOs
ppu2\siu2'g(9^O<":B_Xuxl!BFSV_'/Co3^zWMt)=O
0]7]*Bi?hZQ+['$:YzmS)97$!L3,aQE60Wc|+9^{r<PKCv!%
{xEVoq[LTbCQiZB\v@X}.(eoG7ObfAw&oI,Wr\!gBZ`9&[!g!&&(Y0HyY{,K8g_JbgUlg7mr98&{oC@Vjm<Jkl;h4Yt%v`nk>H@m|3=,\/}P;
Rd7#~rp!Z(He2.+(F1,	sl.FvaX7"^	?;t30&0
8S
TifX/a3pUlwl`I&$H
5'No>G>l}z`#v\I={M-W*`@:dBteJgX3]?9AwnKr4+sPKp'M43,o{-gFOc*	UXZ	iia|x_/C*)@--Gs8Qm(<U.8,Pt,)K7BNz8$v>o{l}8:+^fPNj}OYJ:]C@N?K~3,;7+3~Mj\rRh6AMa^zZ0j7cjQlE#w/6}9EL4&O^6H~sC5cGU3*X$gkLSRO}}Z."u1E"~F2J{XPOHSf7aWrZwD\VAv=713>Cr:qpIJ6\'&CM:d=dDl31FOS/9\U
{DoHJ6rcz#oYA1!7Z([Iq?|-W=^6GrV1;L<|)Y6+l
q (i`5R9b<izvy78$svm=J}^G2zWJN@,J3	0Sni[I_+B4Fg\Y tlSbyQONI.1PiT"#}E;{Sl/.Ng~)AVYh)DMasq~ApL!qh-?#ASlw'dSm_;l9B%T)<h)z3<7X)6.x)Iz=nZ7:YKqtY&	0"#
}yX|9S^?}FT}/'y?B:#`QW!9,?G*,{Ju>)(YS)j
c>p@vd4&HqjfNGMUChFvP`p+
Mk^;A'Cc
ZH;r%X.vQmEK2$OxPfquY}HL[%[='a|l16jI9{tJ|8`tog\OJ"l`sQ2SHv%RP(9!;g{y[H_#-uMjju`$13ozxq^H>{.FsU.zg^?m~5T6b@[\P!^ed6Dk:4s\l`\27c<jL%5~7+@0RT>fHi[Jb.33Ega::+,lN\E;o5?khN,U}o;7K.iqGn,3ZhL ;~'s6)
iT'wDA:%&'"cW: PVLN$]lR_&M__^(Zb87<vS%EyOvM3SBI:6'XUclii^IpV0nd?v"	`\8:&7kbt]?i#Mg{`K]XXb!y8lcbiZ^EhR_AM!oh9}?l(fE/xzo,[uNI&=2NwN.PoLGpI?7~MPFXU!V'\/6))dNLn.2<0c#/S5q k(!<[*Iv=dQjeo|2uJ-hoHBoQEHPM=QdePA\dU]O11#s(Y[2	&u]O>\)|`QB?O9(xx,(Rl)\t|Q$K^y-HN/X"ltIcVRR5~9|T{E	*5f5y&{^Me/IXPWi0XQ)9YCh;x@q=8I3^'By%5	wnRSY5)%%uJzPh1foo5)0/yQ4~EBnv/W]n]{=Uh[J~cIs9wGU.j0<O]KKj>kJ5H_FO?1J&6L5^!uc}))pZNd8AZ>UY&X\ ]RB[<?3DymIfK2wz0I`mg(hJXL>[Q"aCh@.n99$-Ty)'#lRF?P&r0jHbE6fpq<#j:_pac~>n\P@]eHQ<'9#l#9PYdvY8KK\kVV!LdUTOtuw7ngJ64O-&l}mg>y=w?,hZuK==Tcvh07:~g&>3	00x'Uu8 g3\b	oB)._L[pu0+mE.GR:ZwF4{)SPqR&?U5f *bAyi\avH"6--*Y":+y5Vm{ 9*CxRm|iEK^6Eidfk@^T!K3V/scRg#4&$Uof)-w@HlzraA+/)LEd2Aedu|`!AHN{E^Q")%Wh>];TM}!{NxO+gsW|g:matccH-w,v+)pSQ-BI<[y1j>-jf"ebSy9
`@wfq+]gY@d4ixH<'!}j*1.~Lkzi2e\<DsA^RZa)\"Pm#|ZYh!Fq%e'M^5I+x)Gvj;?i-=&B5;~TwT%28UA%1l,ceX6^Y zTS)
?2+9cg||9dOD%Tn!_wsi%tA;!>2?<$xg%hAmA6Mf"@:qxf!lYp=-?@NtO~KPN!d "S\.CR<@SY*Mo~&v:EL	t),e5I
_ez!k!EKN-OuhM>Fn1|lff,>YzwVn+U_#6FXY_7
>V[t"R
9,+eYMY(8#{]C%$=5iAu Y1J9^o#EVd'(3LQE,>hnR4~d#(MAb, q\|7U M+\oJce>OchB@U[X %e@f,E'rVYp{~9O	aJqiat?(^k/Iz}uO{](t,3QcrlqZb_BXL	Qp#mTEAL{-@bx-Brii?82p}Ig_lOW9A#"8vo-RGv6KbPlOz[cJ"!:#<S.o5e,3>D+f_'#>0!qG}=FV*2*PO<Y"^k
U8Ru4PT$SwXqRxN/71Q3=w|fQ`~%gM(}$.:	mYA4#/]>>%'j.[ FSC~Ak+4S[DC_y<P?Na{+3@_<82-0E4eHLl$:^=W!OYfwZ2Ae r`Tsf?-er<Ft@mk}On?\q~WL}Xw#Jt0?5`D*5Z?o8$ErTSFy;M*)`z29.^gpmP{:-[JSpu%
dZred+\*gaQ{:EIl\Q619goZkmtNlha1Y@_m%/fNuUs8O?SqZp5yb_vk2xZ]1 8s;QLXv%u	BEn	>^m2+Sh+1F[!Dgi2{rJC`%*aKzd43UyO+:jz:R,9!r[`i+7Z{FU7`mI(NRx?l`k	57\M['dx3cz1^s<N_KwPFo4aj/S8nmh.}OQ4Qa;2J_I^^UmOH|RHYd6WL]<dExS[F"x%h$,o\}Wyc	<FM2o4eMP;PVk^(nRSiO$9@Z*3,iX_VrA,@C6u){Xt_mnn~hgC7r3Q/[rzZZikUpU'?XNTd@0I0aF|q7mmT'|u")dj_lB{2oiA
gbUF44r,QzGGK{RmzI;AE*I]3~?qzd;2)!aw>Om^%l)bwX5ra=9rDqm{9B(c06X2FE?_aY2;
/*%:*~t#zhxZ+;.iZzr%m@K>%acs+f*W
LU@nIF-Q0|
[M[!>-NDWvXv{H(e0f%RV%1jN,J$?2NY8V9 {_UE{H:&K|5F3jJqU$:/	KfA-&Gm?#(`Qm{JoM3"S~D7jpb*d1I:pEVYbQ#<`Hyz{Dx+o\X1},^B
2EAmxb+3yB~u10wvQQ>4t()yFpU	a0 j:#oED<r.*DB0O**9tk{
qkWBId2H'_mvi3y{%FIrU^4`vUS^@DY\Z"OZjv)	_:z`X'J_PS'drg12:b~{tJkoG;|A@V_4 C?Es,L,}D"4G`1Yh4W ?N_4Yw[eMSh[vHMbD'x+LTcQkBb1+@K@t<+C(c}}s}4!.y(Y!Kq}4(5T*^vy$bVW\1^HkbFvSoG}U>'qmO;av+x89pu]"f:m*
@>JXUG'!l	uDrY}eR<h1D^62`7Pp_:]h&~r![GwGe\as<S`c=-vi}*	5oueQl#DG!jXAU<#l;C%gl^M&!oK7Tyeb\m	v<'vB.jro}tmL'yK}SA"Ex2~fSACe5EYM}1W_vZ(]8aAYlc\(\uag!"HcSaL3v(G]S}J#=Bhl:l
e/gfVN5H"tZlR4pq8wY)6)QN}rwM*m5LT;:.gKIeTX:fe)+"}T*V@&))9=Q<@D<<-j !^JuO0>O$?%y@?rO*/NMYUrH=3Q%@}sy,_&/YUq^Wy%hPEBIE?zs}YvQz|m+E@:,LRIuaKqm$H YwUZ`V79`R49Y8^a:[#FkZd;ZKX"O"J|2;:ndyKN9n>k V"m*YL9*,=%\[HS:KX1M]iJL{yHwhL;,:i1S5TDU08:Z2t\H^YVKUr5LAj'FOX[XY3Bp+%kMoh|+E6PlURrldk"eW4rA&"y[%qidB}&\6f00+DY9nCua+ucBtE*:v<F4 ]\|!
cyXQNfrS}9%GLe,H#b)UzI22!R+v"mC8P .U}MfAIuts9l$aio> e:2xY[1b~XB~'yS7$B$fv:csNj?Um@gD-cdF:cqZ@Jx9=_c>A
gD[[q')N!r|BW),/w=,QOz5H_#,*\P2[!I-$VLbHk5w~4wB:eU4.lt.]q?Y2+Wb]|8^*i8}g@	X}tlP/x]iPt3QA0bF)K6w
NZ{*_a5Ogs>D:]M7XPRrqKE5Y'_k=I33h319c9T%om9aH}As./A:xug_{vCY\FNYiWUZ(\vCi2Dj E,)HXI{&BU)Q'+^8#aWi2[_Tg-EB9G&CRR}?[u`i3zED5>`oCqG~FuG`.9U"(}U|,UDnaC+bPClROT$bC)'UsHPYs|`/L_%f<;COd3GAZlyd9-"0~W`Z9|
Yc[/EiR3.R@4U1a6dReD3<ukknQy#'~k`Y/U/ag
Z=	337Mf5KkZO3WtIhvGE^,2TY	3*+|llaq!\yi]QiQ`Z[,'},G<+\V8O=m/CSCU?\>kF/.v|:N^yx+y[`Dps(p"=D3ylB2?
j!Uqm'[z'SI3J|*E|R.f/Z>r-x$1zlU7&*+?"N_*68s})svNry
kXPs{-]-^u64FZC1PYr+~\h!h 	{VU!=2]@!x!kKL8# [.g0@3: EfS_Ef/4r&cigR)` N^>K^G"}z nd[@;\}`uzU3V$dn.~HlgzPS_E|R;+zp3Qn{3n,p/GiG	Ny7MV?0mxdH%e@W(lbdr>xRj8{^cxr3;SV3o%4vzQke8^\MIy.B7h	L5vP\G5U:pryr!EfsJFqdrXgnad>AOU0)+h=sSIMH3'S6$i_*3<_4J}B8lBRuATBZ>zp[$i7^]VLh!]V(Skj`RLq#`IIF{o|;TWUk2c$"{}6rnT&1`7CwXR.*SP2UCfa2ZE
#`Ni,{.BEgHG0#"|*))Nnd#I0LLTv*C4Y46\9F/1 bw8b!q-N>(WM5 X|qh
dhY<"vZSM^l/mHCJ[X&1Cww&G9?avBo3EN}r'\*|D)P]1`L^frbINZ''C?kW6SEk,t8L%I/>7|`4T4sc	$5]Xxw3#gl,oK.oU%nB-=$	$%jIQeQ0.I8:`gdC7h}Y~a+e6Yn}J\WH2,eJ<r(bGm`_AOYR[)'XJ	n%e__89P~YS,w}L0@:^C58P	zpX3qB'Olu7@Pr-[T8dRi^Q=;54}vmoOf6pGEG)mZ`p1bzS=I:NF.<6sPF$yf[7R_zM:=\S'f@Vik4E2K<3w
W)y=n2 aw)@yxyMoqM:(3(KR0bAJ}Yy;APp-`\B$O*3+M~S]RWd-ho&	+[L`&J.Rq0:wok(wR%E.kfUzp9_B8ibE<e[931@#TWN|}7	2]*=94^4Ay,l*o&J^U?7UoB'~IqGS)iQ5(nS K{ lc@oK7xFc{xLnK _jGT`U4*&L$0
Qtan/n7LVVrd5	UM$z'WE''}9K@U>[//$PSdqi(Zf&r*H%dNh?/|6nBzrY(58;|	7BcAlFY3RCq>.z[1En;jp]5fz.*BI2fb0jp6?k;=;wf#{WyGC{u{?AY,e.el6$T!w:BY{W0F,	s2*Hj}
}O6K:z(|bHaLs DcBN^MV@Z1|dUic\++8tjBHm="r~0 L+zT}+2nwU-}JP/f{\xN~3l>E_iF>]?B%6aPYQ2hLYyhDO,? =:XGZi!cenb4cf%x|]F#&x0RW,u!S,*e?nRN]?KghttLrU-Z5	FZ|yv\W\fcDdg+JOywRn|>I<%l#S0c1P=F']e
YYd|#\3,<{X	&V'
qc}-,OK5el2y9QJ;f5%7hK[5Sy/St4@/C>
%a3<MJ2c&}4Y{|Cv3M<c#mW4P-l%,#,guewNV3;/CWMqfpt=(nF{%`wBa{Qc")W\:S>.PDWW1t2Zh1O_>[jQ![-h.]-6AB"tfx)ut21HUu'F_Ag8@Go;.:HD|3?e=iWT(Dk>1~s;WBq=.,FFEF(Qt`}(LMP}1"AlO]d] e/6SsNGx>r+LfPv>Ae+\Kk\Prmv2ugI\|ipHx)=N\S?oI&%x$xpKs0fGtkg|/:i6Yik)&orwz^SF.7!E_VTx..7OcX%$?{JhF uFkZe}vd/Di+2o}lmSP(JgO6F"9\E\(%)Z<hvS@o@\yMW-F_PH	b!pdI\FZJg!A.X}!}bX3fB&GJsU_.]_xu ]leok00"zDRs<W5jvyGy4~UrFk$(KX=<V<|@!Et5y.%Due69nWbw.C^lYTnAgy_8RVk7[QH4F^>DC!mJyMy~L'!YI.nu-`T*	OlLT]S:*"]!D}s[7}}UM@a2nx./F
v|,.zx-2-2Mb;zl:o/JK*gP*eaNH	.HS+@h~O(2H)B-C.4CwQs1s,fPV_7HLWc5m7,m\/Y|}QSG,io<GrQV0~C/N1]J&!>6TzyS^I?>''^xIf\2?Z{oB}[^^Y-`
"5N-]Aq`Et)E`DYxxlWe!D>G:"L%NTcoUe7=O5 t44i|2a@%GtI0`mC'y9+>fNEW,2yM>)LssRca;fjgA_5:<$?O8G..H alLIN[y.[ [)m&~:Tw:aCXR9#Sp@Rb^kO#b#*[9E
=%&5Ih3fl,{[M`@]T<CV2t0-.C<kP~]uMS&N3,LZa659\<Ie)*oz	GpnAzc;ron1|)lQ<DOeZ*&a}nApW,Zf&:w%0\q=k9!AFXdA#jS;A4!G7SGFf~#e4y
.hUQ&jXuM
l\/D|1Gv6dv{tmBnhuY{mMKdQL>>kuI\M[+ {;rC7c*$>C2jsAIUZwpP	zpbP%drQ
<rD]o5FG&pMwP&-"4iI1N%^faW6i1~*{+'%Xc<ox2$<X.1E0J].Ek@v7N=27R_[o[827Syyj/N
Zecf)hmL!XZ8kzd10-S+,}`b<ph8qXi#uFSzO%j|g
E7"(v$jY,#8BMn!5kI+*XgDksK{$^0b1OoV3(oe%OG&[^~
i'^XUcwPS@iV/~"{
Sv=e@jG0%d!kgU8oQ`mO#c3^9Z9 8/EuzZShTzi.: d/3BY^/3zB5poaZ9U\p6Kev',2w4SbxF9m_^OZ:Dg>hy6YPP1#l*u+e@[J&CGKM|#zQ4ZQc2
]4rg%WAfliGx9
s2hH\f[2\evQb%Sv|[/|>vbpZ(,+Jf\oExM|iOCE
+=7+PUfY/8Y"7~Tghsht
4W)O-0/6g-ks]Q)6J}R_/tZ|U?\M9yBG&znrI6@&NDtDN-:yN7P	6y:	(sKSMxqTlCTGqlF&u8vGrFef]uq&+Pkr-n${#}fXCSX
?gbIZ
]	Y"CfU5N'X6y+Zbd,b}8x+\KS;*+({PG\ss
<+Yi8cFCYcioC3DGdf4oKG!uCQGiFov1]g@X\P@[$,tkRj/QfV3#F(Q=,|zM@%EV3ABQ`CSG
f7;,Q~>4am9al^Wi)/Y{d+kZ%<H
\q[4so.5g&9tZM28A"=PfOx1XT'1DG>&X?[	fM<:CRt]FgGZ{1eB\mH$I8|K	:F~yTd.-N0`,<e 6"p eUB"\*BBc_IVmES5	s]#BQOR]&{7Lw~{Em_b'U3w>jz:03;! GO,b7kpX13%"Tz"E#Jij9mP\t
oV9JA_<mwg:p2~TeX.#g9Vr014+%80#1\cU`a2{b)	IM7F7zSms8NC,=Fd]z.(0inlJhIr*\]
)"l<%GB;HN`v!"Wd}1HN'ogdgN/P{gGji>E`J|%$d/NNR4> )xW>c4^+#xA[pD,+JfcS.vEo4*7z86ey50n;gZ#I6c_}8(K$t!j>XHwXB_S.FDN}@Wc>{;"Lp"R50e~Kb_m.{[\|8=zrY+F*UqEgy:GyZv7P5s#I<IZ&zH	:F"oH-NP-?y^"+mv<g]r}V9-q"(u}U|#'[41DyLj\46{9p{'X+}l5Q3Vfv6E($lQA]{w	s}uLuUYwj+Q<$70.W/O~wSC=TG7_E-.=*=9n'qBPiM_"<:Q]=BxoO8i/[mE2k{$oKjH:{1ii7f13}Q+S:S<:dy;Kt+Q&A]tJ5N:,4KGdC+myNRF>S[U0\=GsxQiUO2,JcR~VRF<"oh=vTq!B(,w@wbB]CYC?qp>`,hW_^{8Pd c&\d9ujFgcm*Gx2'j{>=\B!
0g^rK{@;BWdw5/b'#C{Dn.f@x<M*x,t=2c<o8w\+*q$0JI@w%fJF%Gi(awv$Q"`8+E8iOk/F:Js7wTH5K|0)"=:Y3]t@eXN$0$Sk#%Kf v4/)T<y^w0tjab(oFHkv#}MzP*HQ7_nllkWf!?!I|r1JEPVToE!8c(?le=u>4akF4o:nj^dFZ)TsePwsH@;f[/es~_X>RswC(l~xLML@E!f9&K)5pL@)X*xc|`6gVz&Dj%_NMb!YVVeG/0_e]`sGCB`g];Trku&N5@[2Y*`D9u9A!+u.q[
H5z79
Z!/	xEeoLa#R\}1q{l,5Ytn/&1&_8c(llz,XHRDlGv$x	Ej_2&m>\;~Q>1(>jOU-330Zf%fICg(P4s.9Vw8IaBtlDML 0Q6jL(D@2	b;W219U@Ty2vkV^BlaK3LzkM~W_u'RJ$a*d$ihT?:F-`fJoWiH.ZM'2BM#`i_g,LXPUlJqFQo|*#vd@eJqK$
5['4|.QX=(+7U+taqbbR^e']_:*:0bMz?$(2lr@Sg-xah/f3MnGiGO#WThN)'X3%$Ft'f2!or{a;WLDAI]+6|nAEUeoP}	ED`%%H5]vA0tOVQ\ONi9	ySrDd/45[_gNpi.N|eN8w%?$p<mTR	y"b$s+L|0DaRx|wW7"0ZE8=T5AFRH@Ofs\m/RM#'a2o.FH }dFgZE(`#nI{G.ylarvfqJreGoLaEW`
P3
K+dg"aCiuSX-C8Xe#ICZYN9_%n'MSYK`VF,>C5|k@g\(O_UgRwi_{{sUAxR2iz-=ayeFuqHf1d5GTE>x&IVybO&igW^Nz7TWBr:s K2+@l"CoIj	7K`hs>n;0ql>?bb8jNQVcrI-h|bC8GT{g@7^XdzKK|-2~3'Cl{T^`"l]k%uD>nX~4hmZbf55:D3B3A9 M9'YZRx}]U['1`'X\<bns
o9GIz~rm/PinBo"Nde`;9(K_ F3U#2IZ?d+Z -Cr&ZDc
'&
0<2-*`Lb2LS7NkG4?)>s>qm8o<p'Mk@^?M^H?bgJWXOj2FIv>ij\V&%-KLDTkahoK[UC\R?dI.;(QDrEBrdIu^URG4h-yeeTq^ ?<(/u^.WitPg'98$#*U\DD%;+*H"%mF8	YI>ZkqW]bER:D#$6 ['R|Rm<qvKKYF\1?Lt4pHhbCEfPQ&r8_;I$?tDIEnCjx#W13<n?eMIw+O\/R	$f?.C:{uQ<25$gz}VK!,&EEff\C0d=wAdlGL&|Bmyda5B6\CdQ w5*`i-~tu$(~KzJ@Yd?dUW]s1&[e{mLZ1S!Gf'Iua=b->6g	U750Mi(#^!en \;L9TueSFu hXw\Hk/]8dn,Z&q^5(xE3J *ClU}uq[_}P?5D :h^"URC'8FHU81<'1PoWa{l>egq3?."v1@R)ziuq3m?WrCMYs9VSdq!Z<nSe](lh^WEh,=i35sFY(a4bbP2yAPnA%&b"ci,e$]\%aBjMjT3Luoc'[BZkuqij|M0!4QXi?6,-?r?P\G*|\GlKFb1PvPAvtc~&;NiPCvvw@t+t`pi}[|>}=B.SsW<T
\!*g4$&v61lZW#Uv2:#6Jsv#$Hb0%`%h[*yBjUeY:b@-75u?]M@T
C VkMUH@gtH2uR:8SoF|.s(/%b*V)q9/?Rl\/2-|Uyh(\X==003R1 NlZ#&kl]M#Ii0,=@e|}CyUi29aQ}uh,e&2%?)`6E"J0?@XhZ $m)56FZ:`R|[*Khh/se^$E$ <5/:PD44wXt0+id|x{-8_L!#g9<puc3KDUWt-$cd[nl1NsZ!H;1#<@(a{Ymq;pA=
r{,?LWSg[8QGw)MRTI*sRZ(w|*Wl-f]D87sL!b9NU)/>;Xegmg?\sqF f'+wW=Kh
TY3^4gZJCtV^h1K_k%C	\KBK('I?.l@wN>Os_4*vgl5sm,#xR3@8;`mSm$=q\hGqh>65]vJ+"FKWDs(e:.R20\7U?dJEUIdQ6X)|nzE6,4zC>?5,3U/	W#G(yc;cm-Oig6dpnquuK!w\g-h<xe(lZ/9@p1G=mWGVGn?uZ;X5jHG|n<eIP_rRN]6e))N-4kV+pa[s,H%\^21]W0,2*Cq+`zHh:MYYt|G3y[sjd3YN=o>3|~_wo}Mt_9[?Th@/<\eD3W0TAv{4Ww/>tQl%[hL4I[hzexDCu/SyLP1O	%s6+*+1Yq9&Gi(9A,smz:i4:](HO7q,Q'UQ3zl{P--&!|j[["i9SzD7VFQfA(TDolz>:_sVv
T<=i#B;.rh1E{=^%I{8@kQ:K3raG~?,@<{cxy8q|9bC]o{lf{Gja"Mf7VA>{}d@h!j2*;Y{!<p58^r<Cy3t~"9m5sLc3pHhk<dzySwT60pOKp0,%<;UvA5/$bMEJFKE<t(9sOvwBA/mXpZ"CeQ@W*dSew:|3EK=!Ohs[$pea>0XO>/!/CF2nB`F3=WrD?"RPnJ2T&HC2]KMPd{"d,#jDD"bBQB-&tAq0tH1zG|pF?.zneGDG
5)WGf|^3.wSa-AqUt**B}3mck>?c)"JZR0gyDp\I3@MI{ck<^"8~f3TjglP|A}FL%mMe}x92V|n{IJ[jv[/C32w0%{30#M%A#y7[Lk~{;R$#!<a.:c:O/OY'$7rmV6!A{IQFW2Pb@twTmHA
oVLwe
T0;2(itJ#F:^NDM@! 3}ec?y$PL1IeendAWp>YZ~T9b7KOYdz->-R\?j`)|kY14OA&X6^HTOAKb!RDXXS58	slW7~374+-.Wtb{]F{	d+]Gf&1(hT?#ym@_@+Jrv4@G/hPo\)7"?g1-OugH^/=AMP,yR'y6EFcoiJe3Tv<M QJQ\SjS;V{7o%*aE/fD(]D%vep_[;(VRDr?Y1afE#K`!@NuR?-!ptf%H?:)D8i\nCRw;{a|.DA~dzXtv sVr<.6Lw,S_VX'_sty/EXt 9y%G7g7"OMJ\dO.e.HEB#J^k67t2^N]5!`u]b3=
JX_Me4`,@j-6%u84TB$i1kRB,JXW<@
Xm$dY0r&"2m6C3j*cmKdTAYy5Hg`TeJaBR%GF(BMbXztMgOa<l05@0VvYMWh_!17PV<7P2Mb7nnPbZ&PZV7}Hq[jOP*s>?Zx\0"vTsUA,2!QCHxPi=}D@Pv>V?d7,=L	nt.	66NGA4SdT}KgGDlRbmkT#Jp4.82H][Sm9W{$Ko^rg#+O(37E\HP'I+3	P9m	t1\OD#4*d_e<y>mYiZ>#2]O5^Nrt{3XKBaWWK~it/EHu^O%tb}5U'n[6x,'AsZ	t>q6,EvE 5;HI+Am8J {[}s!32e[GO?bUUlh@2^0$'\6N)VD(nr1TJB
}yK&~Z6US+)tA*5-V81F4c(|4mx6Hy'lM}`dbT|(V}6U}.tfkF
V	boe41)]
~Jmo$mOj)<mv#,g]CCDDk#kFjB.Z{>}OcH!?A6dW,Me0"ZFq98VKEIxW!.-V\]Ox!PZh
((ZB+q*yv$*49!(JY{`s	..X7	Oi>/cyB<8_|vV]p2{9%Z.KC,T{#4302?`Wl<'_tr?g:o`
V=WwLT8J~Krcm8#118%D$UO}'Qt
uS{LqtMi0n]S``SkRMQ_.Sf
b,=hm3o()(rJXvh5B6Xob?Kn-/@c+k)V%c=.?91
9s>M2s!c$d@4`<je<X;'!o$oYir=Ohw/	:L)5++F?rtvu/2*5iwNSV'nzoXy4OKD[i ;]>dpOyUvD3+\"?Nulox#'W2kGjx	(c[v-]I
w;)'c*AUsrR}A(&EWTwvGDTDIuGc(@{2_GYsNFU@rc:sm=}1ptZ+Gf9C-oLK4c?0$bTLY;"2tj3?MEEp!5]U*Z|ABFOm- >Mc";+]o^RZ1;Q	X|
v{.@qD@a8ckDZQz6*j[cLsI^<VD1RiucAM+7^XU2y=>6b.r[:x3Sign5`wUs-%Tu|R[$Zbf/iirZZ0FiDX0V#5BAhHruYxEijlB nh^bbOMDY} _A$4?k|9C!;E7Z`L;D4A"7+M'z:4eRl.1$aud;-uAoV:8.{CrEpKL.&l@^pr'=tHu=+8Vs6i6jp,{MI@#^ecjYJ$&5_;a0^qT)5=HPZ57v.;R	7vgIZ)(6w@8RB~f|zCW6ni:qL0O*R3iE8r,W`c2rGsp1+gSY>xZcTSG[A$/7-GdlWZ.!WKP4cqB6hQ*{KPe{]4~YaT`'c#h"kmdAYpO6$P44]:y|sXwB032vXV"W?RysXjI8-1oYTzboSS{GRkI%4AM2g!N&^$|K365/#RSKk{WDy#R-7z8G"!,[s|7jNz\tKQ$A]L`G{$\@jI'uf|vbHO"c-".~keCf-v97"67f@<_yD	~JH/z[}_3<8cE[KYp[$N6Vpao\Wqx}s_xtr.S ]!YUQ?hqSUt@)z\Pw3Fogq%E8l	pP6r
[!ct	akiUwH;B3L}{g4,~SC~sWld&h`<{|!P:%K<=<`ziXgtk!++D\^*-*~7\-gMS?V[UDgB?ghz<jsMm2$k~~b[@?_)5HN6wQg(+Hb	G%uZQDn1rwAi(d%AL]F;QkzE\+?HBUfh{4ZY`~Kf|<V0ie}zp(Qju>v{gUpT9/8`+~fKL/M<SVAt(,%S/1oe6MN1gC
/ |
9Y\h?n^,3tyu[ySk"5Hg&wX]_4)e4hk13Z	xi%(L'8=5MCU4<?#_eXE_F[>LlB|H.c.~2u-;L1Ya1$`f{,,4k1WVJ->Kho%wGt'Xw^WCD0:\Z/R}]s}}cN 3Tpn::3mSSIl<XtF\;%H6F[; 6~;g?hsu\DE78g?7YIX-KTs5BZ}!]:1
TcKow=$0ituCZF[px{f?nuPk[&\]3$!Y#jH$EB/-crW"+OACoK4dan]Q^5B=8L;g`/#,3Nx{cx>-OVXw_(S=:]R*1:r!]r2ou\a@eWK;z4Uc[LY`DxSP{^l1YGHC9n@-%h8L6.}0Kjl,ej-0Ta(q3\`&F;4swg~'`d|_O,1#_LGzV#H/E7x
)(rU)PAz:zsU&@r#~S=0e	WqL]a8X2N3+o	\J[J`ir0{w!a%U4H9l>GA>YzX~"#N@*C< u@}dp<aM!`\X_aR1-n5CK{+uw^A)AO^COG?N9g `V	<0/G|*Q?nFfr'eRJIZKdMc}Q*f)j(/`<f3#T_G2)hHAl_S~Rr	dt,P,I}T&{]tondIkl`72D9FXw,JxZm9t?VEI1"iG*q^#X(s?A<|68QX~$I^g= *,zu~0ifk3MBKTWBFxZ$K25@#n4IZ@=(J*qp%z|8v6~m7^/\M
oa,USiX!gh\Z#@W)p\?m2]JPF5M(P-O+D||Z
GR\"5v;mWlEg$ C?;P!ou=78yCr=A$^a)sR'g7ze(x)5
;Q3/T^p5_]HEhT/S,!NN{7w*qT!BW7iYV.[?mv`UdQ> ept7EL]dc"7onm}J;HCqlfe$Cq"S*@ig
GHD}UT,XUy9/FG@ CqIVrv<O>mX_4#LP@qsk?>klE@$dGNBY<iQZxI)6qw9}'Ez706?.&$Zyh"*^n?@lt-|LEO0PW1!*G=~	4K\5Z( gZP'pH-d4u^"JrV
;4&9YRteM*2WxW*:MBk(O3H1$r5aYWLSk|J*<q##"GZxWfg4ZOB=HVWd]+v	N.kKb+A?H%>OufQ|h+ShdHJNSF@CdMA>SNV0Pd1$a1m}!fe(r+YU\{f<n^8q*g_1Z/[Z,7bd(<=3[NZ]\-nhn>tv)!"9ob\kD(-L8Vcm4
8V:s89B5sTnN2FN@N83"T|]+pT?h o=+n#J*%wt&AcN2)\3p^4+W	A!u]J/laD!Y+n2)sWU}c3icj2}@d2nYq>`:^HBMLVy]	_'KUN^A^]q4N+6M+9v1t%[~1]"h9dQs4EZ`,oPVWn\q|TZy-AkM#Zx<G*O}G_5QA}_-:Qd
Kt4.e2+cg-Zh$u[_<7:.,0 hlFQ
q96t,N$oNX%%>*D^>PM(@{{w]V%x/FJTpF4`wm7}NSdwlZ;gkT4;O;&{w_2}n)b6	^yv#;<X"uJlTF!s6yHr=^ESbT8spl(W]^T@	\Y,C`kUkYta"~<{7I1L756	)M>F{th2xAr$N)Ot-\?K-b;51X(UW'?\1';s]Y>xP'	_VRfU7d6b-_:AMl4K0lO!bE2]qv@R@vP_}LVv,9HUo`c8rK~<CP=&QY0WS*oC(:]7D%W$C`e3Dja3g(/\^4}de9$GKXH>3*2S7`D	I"/C4^4v{8iz?w4*aYH&tLMZ}sm>7)1ujshlxyr	9,FZ>wej$B~%ckVYexA`]2+?B 6mw~vn3O.82}'X_Fh|&7`!D>n#^W-0ATD>_9Ow6#Zqm*sH4FHdYp!lF	js,B0E+hN}4mxi/.'v=e}3HgM%=f?.,6Q<z_e<c	$(8Lb0Ba:ch|bN'E)k73^W3 4j;qU}ZZ+>nm{cG(4SH*]*htqWp)XKCN}	zgkt>~WRizlf3-5X,CIF\t][Wxl;)Y9jM)-,6O4\<V|)Ey	d%Bfw8S"<ICF]yKY-i.un.x?\C]{IT}gQJ;X>H]d0y$*(,o+N >ZaG9~+Jyi}IF6hA%`S~fEK8*}T$Z]`0]
TtmflGbUn?+)|S(]j_'lL{_v*C.h+)F(pP'eb:.C4ld3woV)
t]_hH2^BQGivT6ruj1x~h*<c=whqm?^Z+4'XzyfcOgUU-C*wO(az%&3LKmCrze>]I5(<oGd.2Rz{lUQ%Lh-;?TuTx<vRoG:e5l{m\&56%]rFv>E;yhB39(W?;1Qn(Z,@f(NYVoTZG+o#Q\fTvx	YfUA*@5>;"5ir5*0JruMbrRc?h~)HQ\wH:QF[j*}
-;+u*84Czk	qYv t	ihz<4-6L~qo	H<}vi]gi(W(ndoO*Jjhi'*a'h#B}X*b;	u|{Bx>lZ!!Gl+X HGh18ZxDvOZpO+/"BtiUQ3z\_,F+$%cjP=/	2UD)_N~:5X:?Yq
+\N@~YH%V6]9\BQJlvS9Gs01w(Ti'WVg_m_	Q?!cLNC{@uA~VF#EY5O"K93z\19X3L~F^J*zwV-aSL)^E.kw$gGpr;,tp})Y
I|=iH"z$C(*xejmw"mAW|kt6wi|d@Z4,cl<b14k;n'<n2IC3BmPJZi4'	J'ji":|E\&?}]s'GCDy&vf0b"H2D"690)t3~	U`q?tvV\#j4T`xo?wZq4@R*ZyL0MQ;pt2f;<:?uhTVqd7=gc*hgN~DBdQ--z xoa}@u$]1NgwYX%_.wIDia
Cf>Hff<oNomhq	pWIcUiu?Nw<s"dK	_)kCcM LT-mtdeHA`DIgd"?#3o8Rq>ApEZE#I$[3Gb=p5y;3x7i[SN-33
hF{q%SL>ZH.Rgy$abw?R'l}B^}:p_4]<UjhfI]$HJzNz`"G?t{=&$(eEB@"*0@.2F0Hpv@t(Lu&~a:k^9&g<yUjF{Y;@bgdt,TgZDDV`8BSK:s*\P8&0/<g'0*Xv};gD1}L`d*$8)Hz'a_w`q.YtfK3fGheaNdC4lqM
)	LU1y*tk(l}\wnRq5]g)!/epk)@V53@[k&)'a<F>82jKqBbDixB?7|-(3He,!`Sm@#wB~gw_)eZ.b[Vv	SKQ4DE}0?]R6S;=I`RI"H)l!<UUE6pOs)wiPubSNLD?HWGvrXVl`s*D"9B?fki;3bZ(+ZE
>	,h[A>d]6dTb-9V )uOJ|GWx}_oQI\i9}|;rr-lkP3b	3wXg1SmhZ`U<.WW
zch$}ky	 Vh$)]kfL+ \4[h~|_{3d))gg;N.6xS3Id{X!@$1~aAla)~Dr|?eG)J6*L;lM"3bp,MPP9Q&=pH#0pUZGub5o~p#)h[71~(\W58("6tAGZB&{qa'Ly	]E`
q9+Rb	vnJv6qr2w*urD3lCB^{BhT-9sjo>3J8'1'83%Wf@5Ji:Dxi/..2O}mGD<BoxiCl}^DQe?l;e6JRNO0(1ww_pjcL
Y%JanO_"0wYrMxHQ<umd@.~*5+Cqms =Q=R5fuyCL*;7Thw;bF;OIh6% ei\#~Nz#4@Z4=k&@*pN9dpC0#xl(+=2`G:ZTrk5JLLw's3IYY[=U=RZ@s^L^JR]`X-k?}0FKCSG*+Y>E`5)tmE`}.RnU!Ho"eGfHg^$^GidX|.jCBN?nl&D h+@ft@e;wf6|7bM=-&^88z*{c/Sj\oS0qgA4<,s~k0z0;cRY4gIjREt2+gx8HI36	pR	%{s}yXb~6&X+XH:k(|?jKyYB\Va#"^ty7]:3sQ`[1g^g$AhD_!5yepFCuh>K%c Vh9(r9(Q=B(hueS?7r(`#DWz5,/-H^!m{U:\rS 
	&x(848<`+E$Tb[|w'Rk9Ed;~IB_-]tqX?k$/gJS1RcASL*xmWvMX'qf/]Pku*;<2yb?jv)58D"(_#{0IY_*=xZ#8f;IR'ipYoQGTfm!oT!!fjds,,wvK"8Q-m-woCTr lYto:Z]l&P|d7w8$x:6YUaoxQu1?&2H._	1'V<_qq&G5=xP?KUwLU5a+#wE?1m_c	.?qgRC)*JMRd`pnWx|;~.Cb"]ZoCYp&LG4Q-/K<)GCM
::!ggs,0mQ$gRia]=k>j^Vu]oNt;)
Q
u qoJY=<A^IK]`Rz~(r	eHKG5iH@_M[pXi-\%<5(y<d#I"G6e:IU'21D)&=`>4|Z.$([ALB[YjrQJw}B;/|[FW'^[rHX>[!LChX7(m)cy9u}^.BUS-Z\zQ?i{yk9S/{j(OFwR5^<LYyy+^BHl|	.k80
eH"WH8s8uvYAeQ(2A8	A4ZPi6'Ds'!y\AeN,Z,n]>kH?}i7Ths}z$G:L{=
`eP3ypw1Lf$'4OoF/V:FuDLcmx;[LmX[}?_nJ
&x	@A/a ="<bf>XrCgY~in9cKc&	e{qE	1isTkDVI1rckri2Ymqf=n8LhOB\O=m`^#v,Fc9jx?l<j6"RV[zXJ$
p^IiApIv=t- <);8\G5FyL/u*0zpp%|C%@&YE_jLJ	wCsej:+	FM.;ZLENmZ$vJw"+n/KgPyL847IF8E}[:=n<,oT6pad!C6dV_z7<kyF	n@!6@/jPXOb?]c7Uk3_J8"Mnku1*jE
}9B6CBYXQ:LSI"eG8d@gE.U;zh\RdDq@N&?;T 16?{E4P76T1=3rt2yBu\{[UoR!+;
:LaY}!k;<)a~TBI*rCYyfUR_D/tB7_)R|/:7#M<WFh:ti#@)Wdv(cq1,3>Li[?7PR%S>C_t,gey+=VL8n|"JIW2^@Hu_ToP6X<C/uxg"3&McJC;N-af2pTHJ2VY7L]lb{FyFMVBVol/P_$%4d	pFVo%WUlxyU?H[gj6h0\Gx[Kdw7Kh\C0npB;$.&W@{dv`FC2q	XQ~&07dLji,sY"ci*saq1%<Cj5C#cI9T'i@8,R"N3.1H)jCm?*Vex:|CrtD3=SH	$*"QevaxaU0i,a`=Bjhy3YCju4=/."69<AAujbasMr^g5j*_hLb:h/F	E0BO^6M`R;v^t_ifA)
 FQa1=d[b;N%@{Y4YI21W']F:3w>.TRZa#xNBaRP[33NJkcrF5Z)1zEu/'[o8zBoo:#PN..C6")=g+d`f7j\g+7<b$ h7(sI<;,]B]z@B\NW-WO	/s3
S>( <F.{a"/{FAN<]bXlrVuHea&S3Got[45aroG%I\{* k622tH;N*L%|'lvZt1+yGx]%W7`SS87uGG7lj^7APh=nSYuxg-_6tpLm!18,o.K&#aY&tNh`C:0:]J}iW9i_*WO0m}3Z.(Q0"%/f#C/O;][C{AS
_X`b+JCf~l._qKswA1.=Cz_w3AEM9KJsv2:j)TF~ "7+ [tZ![plS)]X ,WLvHH|	UN(O+m}246oV|Z^vGMmS}&lg|g+P6Nek~SUXv0F qR=;I&5]N_|=%$UE;~prGB:hhIa<r]Qb6$E:5rP	4gJnPOP"1|6?D8#/b*aRFp^s8Lze\
9?jY6~PY$HYP~L(7t~VI^LB(L["1NgrN_50')vq
uLpOD0 [Al,fB.2z&TL|D	l-/O3O.n8<[f-~-t,m_#=W}S]171vWSDyt
N,5\v:oFVq:S!ojKGs2t#;&,d!'UCselaLu,^| (aV92fpVm$^<|p*?kX(/6JW%hD$<T!{zZ13"q-n{wn/dhh|)G0c0?g[_5e$+/iY%q1HyYk0e$cw,0&lO{vxS	EwI`@R]:S6$1(1 _A_{fm{o,=*mI|g"wi042wjm>+"?ve$az*uk:!,y9%6B\s8G@!tyF26~"\|1aQ9[ MBfCL^OkmM2i8)A?LBS?''3>v4L7&\;rt$10y^2EOPMUbH'[p0c?s=rS*o~hlljMw3Wgg4v6^Bl>s%:ZS^44VcXv 0[n+@F!u.iFoJ2 t.9$ucaZ8FJ}n^u-@0H)n>S;h/DCsZJVxd=ipAD&#R+?{!o:*ZLkjP<'X1pv\-A7|QrX&Y{*,rFr+wL'x0?q31K/_~6fV-2,IPFW$e:;BLEo)puo.sMb\Pa0]8ytn~L9A=~`XvAa[e>J'ObBOS)#7i:YllMlf+V$z	ay>KAxo<]&^(KYq+%0c$8)CK9<u<8FV]bod1RUQN7A6"^~(n*ap{h5ykT+*l_U=!~xxkmbv!M&<'+I@hW#2a;rlRP4gMlv3eg4!2S<p	bO\i@M\>u {INzp+9hP>W5$MRIkhVy16mH#%buUO2	<9n2CO&Q<6f*],8Ee+@eq|7:P"Ie!{}MAc9'PG>qFvwp`aMqn}lzO/5'k<@'+#-#ZV6Fi5*
x8)*py:ED6}rU}ytHDi
+JwNhU?4cZ\eXcYB@wL|dvRGF*hFZ3(t/W2>h:$j&v^COep?,vN\Aw{|]Ou+w{6,z[1m4V>I{{IcTzC"kzLCLeN?]fgNEmavn"d695{03 "`A|XV!*X:((OFM+b]3_F##D2	ames&,5ccln.
_xF^!3-O"nu}}Va7c0_2f5vcV	_~A0Dxq^^QQ7sMIi`TC"-h"2w\
mRlZBN=~Wdfd`Ni9am|)/?[aUL=tU"[	jKwI/SUJ[ebc(w4tbcVDP.LDT ;Q_zKaC|8V~$|=p=yLW+$7;CGm6!#]Z,zL)UrgqYI5RZ,W6Xxe0Q,l_x8$R!_BB/':l%-?gu.-sa/^%mIr:}M+nNdYg%I)WCD=k?SBe	wIjl*L5{hK=WAwM(.=nMfWv9ZrP)WO0069^(f\1?\Nuc@:Q)jk}ZZ"&j8fAkp,r8MF*0rQ!oVO
9/Q]NI$Q3g`R\$Xmq+RXY"'`]?H"x4$(V{~Is74POZ3gWvECcyhvN7l3%|t4etR<(4qb|^j+Bs]lxm(>R
jZ~60pOc%E>0W
yZYFU4YD.(((*_`
b~X~F!j{Rx4@Q+\OE|p3i4'eA.E9KSQ.m/Ptks0;[E'U@}s7R[{.sos1kVug#28a,VD[yn,i$BOK6R|W2S Wt#LCBN?ifTi2t+A4y$BP8"Tq^g1/KI*cO>hSEs6,8VxofId(|[0A1?2?y?JVBk&9Hi%b)frYX37pI>]{X`@a11@#n`mB~dfMP$+P}DbnoeS;I(Nkz:v^gSMcQ1vcQ4HFC7RPT$/na%r>Ex,?).Ig^8'/nPF&|C0B&|?ri)@kFqh8}NJ'#=(|L#
(o}\	S&!@-#uA/1.vS{Qp~-}bL>j| <hELn(*tSC{)
ZqhdL4LrFT~NLfS+[|nOAIUJ#1+#mc,J>B)<bOeZ;NZ]i{\xS)>`8j|)p/Sv'3<t@cLtBmPaNH%tr|\;Lj%%]^%cGPr-'eH+ToD;4"GH	.N^=|jf2>A; '@L0m_68fLCf7$nGItr<IH&QZ2KCFmmBStGb0C>@@I}Ko${lhb\&Kh<.y|e]6,*=L	YhMT4	j_UBMA)Tu4JbfBaHL-Y]JKt<hym]:31Ow4@HS9!<9uL9Z(2f]-#?RZkK<Gp=>qc+)dD<:\B\?^)aRTb4cT$:JJ]L'FM-}-gw$p8)Vi"r)2]uwZ 
=	*FLB
T{,+IB	q$hUzu+,~:Omq,#,0E;JsM#]Ua$y02Dp`tl)!GVX/U8oxG6\YwhLPv"hg{id=JIz_MPSoRm`U6[f`\'pHQ+.g^h<E/!Vt@0B"$@VLo|ge,a};|LTgA/'iE{}>uX>0P~k~-9eiz/Q`[CTZ;~VI$-`a& G?I6~vpz!%N|&$zW_$O$\RD&{0a(/xt$<9;Z0[|9m1rb\"@*3BP7yhM|axhMpKQ74}U[!gAN	-?F0%2-P@=%]~t=IKNEfT::.>S@B> ]r	XxYaEapR[y|	X~|WX$&_{UtCH.px_Yz)Cqtc:\6@9uX1XwgK-},maBCv'{Pa5[@D"3%c+B<LJ~_O\NJql=x&8a3+@~r3XKbU<\ZdBhOT`C&`7CT,+,Y({fCr%uX7KK+<}4eO	N:imdhMoIt"F%F:a#$]go~?a>Vs"r7id]#.N=y JLB7kFpsJYk1gY<	jVm	cEPJ]:+j[0
pHs#v;FT/bm60`N#DHgISQcmqpyr<vysPdekSAfAZ-Ll'O,;a6S>8&>vc@yDYwD!K=j3}aGsx<t7/a@[|\S
Y6{iKVDd)k1qI:t<WhXB<y/9,nl4fEMr~qd/2~_bH26+dPE#/]CvN^x4>-})_xw_RbFl*1>6rp8mEmC N'8bt._]<(+zzp#LCUB9BO,!u{+<;`v{2iKtnFNkO.}YF
-O`6+;;f#

(v+GtkpM7zTVl{rMzVkdo^Ik[7--q3[6sfTdkR:\Rm{)'1/L_I1Y0/0~;bTr;y7bW~"L3R&aw*dK8)bVvu2Za'/uP"BjI_Eo_:hBR7ljY/>TWZ Q$hY'>,Pma0,mn/({;MGA-'h3F|
5}-2-x>6W mcazKg-v*
c!Zi!Z3Qm]`_#TGalxjNjO.e/p~OHU(y*Q0-{.bjUDoLBbZ'5k=_1kCNx80"t93Qr8J[Z+m9"a|YZ6h?o'aJqMIdz3#)F4^<;-Zi9.AhpS@2F^2/KT)M\qE?hVDHSnC6*p/b2JE:U/n+5XXoj/.)Y ]|@#TUxau'dsP0-jQY6M\#qaZ'WN7-r4eZ,,.bxzax&qw@DoYURVo!bdWNq:myzNjpp&B5[Pd2i}dfQnMnyzmaQPG^b]a~fWJB169NME-*,"r*[.b9S"\zo}ec{Vdw%P[=dq"9]YfQ .a?]yV\\~u'lGm5}m!EP(9dY/qMajfBHZ
|X0	7,/6oe8/:m@xNRW?28B#'2;K~ =Ggy85 `gwU['Z%Wi$/J,*yLUKhT/CUi` 1xlv:TvwjW>rC0xJh5b@Ac\0yYf[IUx90=_o[t]N"EnsQSRI?c=+cfD8xp!X2/"JOuHOAf;n-E|r:~BV?d,.$?*\lllF:[n(wgSg[t	yl?MyDJt5@H>yMA4a	C6A/guufA2'wZV4?^FKb/$Rv8q_ex +Vp		o~m+?kz7q<l(#P3o7@ug C^K8OmOs8Yj-<%x+bcq0Qh+*@v=UZII(u6oMcVk`%g0,!K?eBId|R0a%wI2Tke*sc|ki	t=0H1e[ C5L$r@=;-xoHTX]:QSseCfg;_CERA(H(`+fZ<[hI^my6~1Z EIV!F3}W4s)o\4F{;v9KT<$uZUD@)+hY+Ok$J[`i8lKTXJo"g3X}#&rRqK*Bq	:#-]x>;9#yT5/)M:v.(#\xZ0^@h>_m9n1Rd1g+0bZOjk)H;8'Dx-":<Ci^DvP=t1cy:#20L&TOKTN_rh7@<2&sk1
|EP_DB^ 1Bsq3xvht|}!|	@Sn fbSmy~Od"aM.vn/|U%nSb,0N /{C"nn.D;<F.FD;Wt;'!oNy4h~eWma~5-:j9tfRsh?BlKB5%o0I)>Z!fc58FXblAqHKtsh`e;^+&w^l_y9MAC_+BU V8I8iJ_]d`#F!&H#?-IE2@Niv;q-0yd?hm4F]OSo[x;|z6K;M1`0`0fIX\xxbzCEkk3z.Q2/wr=ZK'0+=&o?$Kx[ILP/fW |TBkH`6]\yrrrS5;\Tyq5&#_C>O*:"%*)!*Tc2%'()+Vl'b zX>V/9Sd&#h~)"`)?}plPzPx?$]zW%n[Kd>w`)z4p 7]pQ\&4MS{]^quw]g\V:e+Vv>dO;\;VlG"~`4IL|&C(HP.T,PwGI$uywH%*0uG;sXSKg)Ntn>Ix!eO*4'E|}uzy2[1t_#-{%KRg4}>	J|@[izO-(LQrP%;cICev}FkT/?{8_BB{cy)z~hIr6R[p[ x	p}~r{phx=!oP:sgC$a:w.( a`&Jtva<:4gf78?SnmHpuT3^RM\nyyJ{.%3)usBfgSL9;~rS^L@%2
"-Mx|!~{5XypWM@:wx)$\$n(g"l3bXF*gIETgI>5h&*G7M2 :j1NHxE7#gQ2
{	Q0;&hi<HYqqI'dXSK"qvT\f?_ts2"Zo{qHLD\QYAPpbfqowFbVb@fIoli.11(]dTs<UNa6}l3OZLjp'|P`lUsy-.5{J(
Y
=I;(NDO]b|58[R)G0r%@@pHk=UC9V*h<	6\/4]-K6Om	q`	%QQ:f|c;?bPpzB:H0KN/Ct	D4xVW(7`qNAZuSmJ>?VT JOr)*lShw[~h;U.[_U.>L87a)~D|'xw@HHen	WX2EFK92qj`=EO]FawoQ(
X`]M=W3QC:<L(K
DSD20Yql/@\Ix%D}q%sLu`r;bfX70DI;@X)oRT:y(k%qw7Lk43q)ST*HhP=.J"JI&(UuR5D'm{K7[1=&KX	VII9>P'Opk ^/O<\uXTzG2gf@hHhDa/eln4L}28W4\|;_
z`2j)u|m.`HOwK2nqkur
vcogiCCkV.F?[QQ}e7ZXYa{ivC1e--tIT5bh{!dx	#Ri-*$gthe7'<P&:ys{,+7yS<1zxP$GT4^N1f%IH?2kmB<:+3ebwQs&joEC{ANhAtbYgE@;+u1Ps=DK
I>;`l-TK]99!2p
Xd
8D64~yH-Vi9|.X>DHv
^}
gHEmPKAq:s9	d_{yqi3y|]r[2p|7afxD8rB%Z)UYQ>f*HqI&SB3!21Y?~u~\<@sIUYhysXSr
~w10<r,bN	EPx\ajRJ9MWh0o*(5gbG9c)>$"5L2hO5S+1*.e.mMa+3*4
!Jc:=?b(TIkq}u[Kn5coW=pE~o-mRG2X&Z4-WGf<n}q|=(qj9_jH.~JWK'H6+M3U<0n-qQ:J>~,5!mF_lbD`"e2dM,$1P2`c3;eWyzwdm;\ZU,B>jv}CCe$E~efg>r'buAw/fYXk?^#J0'X3gajC"$7ir[,Zj{dEF3+^o\%4T lIKT#O[(6E (_~0[[Jgnh3D(Ews<~ml<P/Qz8-*m>(oT{z-/azyS]hs`EXP#lXVASpxuy!yH^VvPjDjt5>?1LyKYHCUiqh@#K9b*4uK"De`eeE&hOxH
ultOpIFb{rnw'F%U;CkeBeADQ;"&)0(t&B[C}5:MRxz> p$#RAV&wU5~ *?5]_D](Q ;-v#G
5DfAc<RWFD=FM&ZE\+/DPx3\A}9Od V"H]A[!eb	i!^<@yo7Lk<X"8hmqO^MR+t?d,uS|4_}A2/E('f7j}b~2`rZ&[SXUUX%\me6ISX
/=}o2hQv?[,7HHRTS>Bi}Ul\6K!mVal]AjE6U WDJU|*D7Z;k#6^)@nzjB}}{b?9eZC!Z4R1H1&9S\^XVQ4$IP*qTV]kzM4)vr"}`C<Nfc5Fe8(P}&RX-nusP#@>C#	!42Yqca	z('-eC_z]Du%?pHpt~DyY<1^r<?^!9\.fQ2I0	[I5gs_L6/VMD`&yw~JcRy>nT.Sb]+'j
<K5:xI0;	zvzyO)c:OGU.Zy!>k,XO`z$M-u|mF?CxG0xiR(j\+>8bBv47Ey<O,;}\L,#:AW0 >U!YkLsdr`:@7Skr,sa E^aF\}Htl/.jaZ@.Cc@p*lWsP|!"k((IXXvcsB6fYj}L{?tS!:x271UphKzJ5S-|Hnv!GvvUmF|*nIyj{f}U9]qw4uZ)WVh){A'gIQ#l}Dmb_Q;'y,;tl&G	4Pi
x	;FkU}^n>N/,ecsSy*_vJ5@vv5_yn9Sh~={6E>	:bYz:Mn&_fypW
 US:5_@S:f><
9.'i3%.Qt880E}$]y}?9mIO
{XO;n'[:
|M*B;! kae//SZx QP$Wc*@H>%f@9[PZ)+p@z6o0oX-0Bs?4Tmvv-VG+kYs 8/v0j)%5"KGW?)&=^PN$&&+nHe3%%g73la-\?ZPpAw& 0,80_N/@|04@iB9J2m#,$jt_"vMM {8gZvIufY`0*I- GA=qFM)PKhY|(4S"`kkDY1g6Onq?\tq2o3OpUJbO^Og=i*CxyvX<^fpQV9f33J2l$_%IV8wv)``'uWYZ'ojc|u\<AYl\KDWc[[A;4.b]![8q&EDK/Ps<viu9ml}}y.dDD@R?M{J,_8_KgLY^f@)}Jm2&)"rt88Mp?}gm~Cg[SqM
PnE>p^$4cXGWcrv] 5zbjXdwJufbX&[t13#+e[UjvQWZ`u#@SAqozh6hU=64;sg4i$"|s'(c\xt1I#8h	kpM!ed-w}yV0	J{6fRulr(Bw>^<12]
SvRV^cj2YxUZrWBH$`EAPj&o\qZusb<|`X2OsmI^HE+pt{T9\h;d]?<S}u;MYG3/Ha{f0`e "*exze VVE5.6O:JQm:c~oo33pdMS/K?pZQv"0[/LaZj2w%ACQ1,EEC_vE '(e3LFK>$b,d(U-.9:U
`avO?;ck@/bHUgA#Npx[V(*(H\*dN&f=}k MC
:Sm]}n_
AYE6#WNZww4})Z[0utK3Apb3x0nK[~)!7g%kQ +Im`WLf8m-J'';%6n='#EG>RA;
=cX91I4#v)i{r>=O3+eb7ULYuhFf	60BTA9^AMh_#2jwn@"Y FI9{zno#,(,m?{jZy+/gZ`*$$-VT[d:0Cb?ZjL2I}mu~/Qr	>b cWT^w2"9MsbKoM0QpX&?\q4<7<gu ='1ZYW<`Pi:?icj;)3O[5;	*<,zpO!nQ"?6@l]GZj^y<+xAX+K1ZiI%P ^1xJoabq8LM4n9hi?e4.14L0=;_^Ha~Adze-Z
\`-[II6X@
&%c+o(:}*+30/jIua:pNup*T3e wHF|^[vU@8 O?d'Xm4{+,SP7H5BV{DL4Zg0Zd
m=.HRKBktOK#A&:bHQ\9}5Ty@XB4aEM GRKPy f]4:n/954V)U$v`7#/Nw'w
;TB)XH>=Q"+.Fr_tsRXh1jj4hrf ~>zB9Ar`d4tpS0MH`
R61".d{N'(
	UByv[9Y:3$>&IW	46ka<3ZlV|@H,@O} :IFh&+deQwsqE{Q|hQQ"O\A|,;zjq.</Eh%%6cV@|A$->$3dKQm^EVqhJi2i%TzG4 9keHM]<q' 3;,SEWG~Hfn	shKe(aWhj"w7gHmd
"<%eE"|3{(dN
V~|!ym
eEJc5d+6~NC?3 %5!}.'*Nh1}W)`eI:7&vWlUv$-%~|;d)o1ig"D{y[OQQ")!^z?Pg2i5?av,))D)B(<y)#i6$a^VT)&#[(8*sSvF.V#{3}/Dce~_G+@h.;L[5V=r~k_i5lm:mI3yBT]lUVrqORl,L6FN{:{[n$].	-DQ,ca!>7i\Gvb,64J|7mA<Es	n\bqO'(Q0e.cBlyUgs"76?P
F/[?Gi. Yc@6qG~UDl->H$!`fSe r`D~>n>Vv-{L1Swvz2%T~]J_#a3x} ',C;:C$E[M.A5%LmmESj-SDNX]zv	LU)HpeJU]F8Z.pcT$X6J2{N>(4j-7BCi\np,Wq-<XGszIVg[Xu3Q|"
B$%ZFk!3IWI$px5}wgYQwHtM.e5Q\ue@Xban1ZI>F|l.) xY.S;rC&~dA{y9xO`x>Aq:J*>{NWQ\"Y7/\Cxz.5d/v08;G@ubr*u3mO(FxK(k% Nr^(?ZOF&%DK=Ri%{uhRgMqc:o8W,3SJ%ButkNlc&U"`Hh[	2e`3%g1o7ttL.JjBB`z;S,N;(wLa?8I%1ACL0^$|d$d^8/ra3$}GKwer)rlGnl'z|?BH7Avn2=lcTQ#IPf~ jRH"#oS0aB-Eqr]Gr7;&BD)kh0XrS/(/cBo][+94w/Y8i6bxdc,#p.MHx'gQF3rW$o?xh5`h~MQiS=;{}Cc
kWY.HXuZ:q=>aRH67a$e=o>pMCTX=etkX|"xI:?)`}"`
%:,3oo0yIY ofIF{LhQ]Br:%?DJCZA y4U5T@z8e(CN8CR\vawT4vo 5Kc-3:1qi@bbV/7\>C]0g8/Ei/`G"tr_TS0[jAwz](LK#/<ky~LjWZz#,K3DK^0
+gGf~S$dL2}<-00 :8#yyM8[F|oyaz:>=IdR=63Vtx.}tR&-KXeYr.9a~7
oGhUw'=N4y((hw[Femi9w/K:h9xX|||K[g@cJ%B@ASK#h6J9e5>ue#G6<0^'_wFq)|)hOnbBoU}s5I1C?tl+j"+/5},KyfcxfbT2bc<+2Y:II(q28w\]R.+{77	 huE-aSV'Q]<9_U9~92JQwfUf83796B}poB+[|2wSv[.
P(g'L~tB\nW&d87m/'ylQxe6HiU\/4:2
z~f3<Ij,dT)n$ .PSr	$1UN"EC2WBD/Lv}Pz&[=6fe @JLydJ65?'b4A]Zsa}VAg}Ez'/g^*tg \aIOu:zY$o>4l)pQX@$hjT3v)&CC~(:15:Z^
y7!P}(bbm3.q6!S*~]ubr;Ay-";Cl@A:w9-lXd}PD(O-9"Sx?	Ph6MRaKT(Y!5SPB,fGm`]vH_}2U>'a9^Ugm|baV4<Q^5%
A~H(,uw]v0[ahG2MQZ'fqzGk*TUXNQNUx.~";Pu;ah1H^^0qYCDQ<(]~p45N~W<J$V(ac.YHNG)AiE"#cuE):<dl'fiE5y'DYPk zEgts}S[]V<:lQyV_8'Lw%Z|u2}~GSEvj-ek2S^EUj&B<)<RY5MDYx3byNh.A=sD}a$TH%TYJ|AVp(q5}pO5_SvUX7:d+W{EvHA$pn%fS6e/M`hf}vf
+~?JP,@nhe+(jnq)"-$dR 3$p2vO1p ]\;I>/71X}EK!C+_3KeI},-lu`?}ho16\5'pNhi/.SR%#)i"qkpzKW/$^W/|rLr.O(2OP%Qi!b@J\}Nst))XdQDj^#{=wkX(>YSNI>W$AHR@R<b:UmM<d ~|'ISsGV%YDr-5+W)e1<8[q^ULR5:K4BVfs??#*Cy]!]^;r%nW1=-% +cko6zixV/S_cQCO$ { T}:{#h}yp}W8e'nt_}n?\7/S#e56kny/]D#*7M!E8o$el83%YC*{f2626DehOEes?*;MU*$}YAI{4/_/+htSb7ZdG^&r$s9m+2uH	1fo.8
 _hypHW?t;], xa {a'[GU+|$0"aR3=im*;#+;i||dbr}gj;&.=FZx!&f#B"QRf^GykUV>$jhcRWz09[}@(0_WBrPxW+3<974?>Q&nMc+"801.9bK3MMLs7+7	b5LQ23"8Rf:E+)A{
dJNDOTzV'3YXfkYTU;4[vZ<B6"7^@&%yApkEVL@#}DrxgEYdqbb)gG^Mn?[9NSg\n
guDhe]G;cfRL7LYLUTQU{hHCW
>40,xcC$7U4
zIQy1\WC)"FJaUTi.qaGbKpj(2:-sHhdQ2.#P[;~WbEV5ZD;pSO*<W^'Fd.{e	5hbf&)3Pmhs21)t 9]2}i tyiD&JyhQ<f5:{2K3hIe*"MAl31=$Z\g1WvNB"1]%YV|TmB$2M9M/i'l}0l~)qgfb{[
D7Zwe~y&YH\#z=q+_<a \,uwB{Xf=:q'{C >dix#,BPK +2pZV>gK;W("%!W^4H-pHsWCV#!nj1u0uu@Lk5o@drXuB}#oRKVdL"W1`w6=Fk|XbWpHFken[Z$`9j.$4eQFW+5&Nci`-B,$Up[Y%*4$7$oua)s\^Z~P7C4`c(F~Hk?!#*\\!FvWHvMI]f5DsVfe(N`-s3hL,$B5Sym2;dvByr\5c*!xgR`l1~bym{%A8#:akr0gr-IdscX<;u-Gp_J|8'
A"1H
Y5rdp*W%CYh(u-c;O+:vCW"73d`!m07N3N(ON5AT*J-T\gi.3x$%Vrkt?>$@gA!#0Y@:@$z_U$<hs-04< vp(rsj6-XZ_I1W%Vv_Nl81N\ c
w<n?1no-"E0whb8;|QKac'jj*t;lU|]qZq\Qy?o#(J=&qk3hUi\*s!{;FKi|N.F5D=j139_g+w@gefSHuI!H'5{]@p)oln\'.Tuh$)S@Nwq1PMTzOy}1I-
Ox;G_ol}m|@q58dYM:EBHR&:lY;)I\L^C|c]~`9,Z%5D}k16n:Siw=TjN%~0BBidkG/XS$`h-@Dd;Wyt:6-?h+h<b4-1B?hv80n_2]A6t^N\0UQbeNmah.R#k<;#TjI`I\uX#^W-A^m,h%.	c1R3Bi>/h2Tdt'R}mY]&zw#|Ik13\hOp}{H!".NDlZ-==3ozZp|{Nr9L<sZCHptWTzL	Ds),HF)10H<ePx[6 )c70uK>#EtzuiC]nUKr	(/pbcxFU1+!`)Axl@$Wen9IW+dQG{hS}_0PbK!g`!Aw)=fu%n\YJHoZkq57V"KTk:i#.FlB5ck	GDO:ZQ`J4^Wf"~b)$TIyn
|sr6Udh~%ob	xW"1D7aC}{Jc2[lY+qb
RL8|{&CQ%4aoc0:eb@d$;tNS!wF/
\MF:1:jSqZ[&$e&l5H -eUy\43nP't_*C|[0m!"jcHul<9E-^8hDdG5#X
=d1oW;w>A^S*xAIDdqndW>.S`j/4B}X
kP4RhbV6T)L\
B953mUJfv=Yd3%yRa:h76gMC1"I|^C&j[dn2#g:H7+z>E|M_)okn\yB	Ah@#+
b^o=W>5d9y5{hlDppLuYpR<s W>pfb{$Q>is6fZCiY)hoLz6PK(,iByrC/pTX}#TQWSQ2^u;YyWrcFL'*8m4dn278LE"|szu_{8V)MQA MN#`s%k#n38xng>8zOWDL?zz j R[GF6SHfv8+.SH_-Go[HrI;mDffk@}"'$XZ1>jj.7(=*rX$\O(oZleHzJl\%yY=&mFgG=9 ^?lR2-	6b|M e\v|^-[j%~Y\6[RJvR0Dz!\G.au-$kl0J=k u:1nIaZ90=7yv:KSC!4R(0%a%zzQhUtD(K}yx%:euS^C/Zt?ioXli{xbB6,<2E43;M5Hj0SYFWcH-%'Es(Q.Eqz(=XZBDkX.|R1n*B^1*qrOQXa*RC2lV+%WI)W^\Wu[\&Rp^.(}a+}EJsb"e=B<5T%K{jQ3ZwJ[Yc=IwJqKN[&c>j#o?-2
,sCezqMeRwvhxd+GeZsb60P5.l]!8,*UIxrft\bs)T	H7M,QJrh9[+;fJM#)p_g[6!qV#WB	%2VIY9wqzzRcMfsx
UKd '=XZ"KAM$V:oO mGF=Hyvb`chg\?;^dZeU6?>rwSrL?k%3~sYRtR<k&73eG6|PF~	e+UE,A#ZqGD((r
{{OFP!=Pl`6."Dv0d1dq|#S.P?4vS+|B1K%#LQ_M"gE1WuG,vioVz OT{SEdnzc]O$0\x,1	zRqyD1x9z~Ne0>3+pnn;".K!J*E*s:}|huL&}@#tG~;?oct/9j\[+I%CV'[:F=W[v~u31h2wMv<H/o{ZIw0r1q8FM>A,#B#tvDkkk]1}Hv6lPaMp
N:!_Q9Z~>Kk1q"M4__	|o\g >iuKv,;xcoVc<[# Db"^N`T^*MX$?,NjM&~n0G&tG\oT*?WN@OO}q=b%L7t8K/`\p%q"C^!7ffVxVUw}1O0frH<BY/Teal{}^b}epc1Tx*U}pxf"==2*oAB[YIj>|q].eB;P[/Dv3~KXQ^C6_<0QQfKcX6RA%,#(P%HEGO'n71-r0jDdJV]v&+)A[`Gdn`
+.r*)\Ts96lt%ik
KTGvg:n+-X<xX'z@2Gg7J-gsR=SWubs6T.O;[j_ewawSPIZON&1/7|Ffii({mTm{k`BM8'"O2[qH^Bb\c[Fzp337\6`K[_	?U\B4>cLR|hjIjud3,7StifT+/%a*ws })uETDiEy!.IVMGd2r"QMY%@R^lKqs&8f#RG 'IU7T*"Ld{SZsNs#a	)?(WH~oKoX%|>MfSFM|([Td-~	x&+NNU*aG{$j+OZ2[9L80>_DBE3~@1/=FGkV1Nsr7\
%s#b+G	Bmw+u0.xNDWy4\YYBOX58?rxzM8xoxIb-pji7{q3-Ns8$R5Bj+b.x`:<1GH#DxIhNQr|O^{z3{iY^6qpxs]e5F8W{G#)
1n-5G:WisDdBzgt2Zx-BTEup*J"ft
_r#'~`L@u.(m.yzVX{15#EHVM"O_4;,faMS*/|G!fp	(=!uJgF^!g?LYe^:S9c@n
q1q-
)jsWFX&Ty=tRtww&Qy)8
_$'X=@qEoR^zfV\)^_&)_rf7QT^uzm WN]O#MC6@nOG^WWz;6tDap2?ai{^aDTgr4/r6$w6Xd2D_q0!]hwY4L/44FxJyBuOhrQ'te4RVq!)W1?/<_H=KJ"S6Y&e%J~=B:1B n$)n>-h#(Oi=I80AahWelb*Czh!/t'2L/{'4% h8%=L>5&z8MS8#'EV--/H3p\2Ic&F#U\JGUoCZSb[MT/U+^f}+&nwa]g!Uin)FDdy S`'}tWq,x"\PsnTcM&+x6[wOv@8HA-fwax;"yi{VS,f	j:YPXT]IWOJF|E;%A:sL}e6d+vuLS35<Xu,uc *M>T]f[]A:YIoegO{:tt:HW@l'cZRSatjgfDT2HN:HRxH9T[	kJFvH-|o|['!;;7K|&-	,=:"A>{_[NO0<@FRMz|[YH|+A79;R~mMURS(|!PK+"6Rk}E@rb>R5}R)mOnj=fqqO'G:XvO5RSu*STH S`HFqps>'aHyuBRtPO>0C9BO*9}sCT+VR{:$D7tgt.R%YX24{~%v]?c#(Fa/ePbk&K95)z 05$d85Pu'~_"0.#W#Z&.Iw;wGezt^+fWCw(lm]Fu|kom*HHfvxjfm8<3`ab??<Ycf4r!:d3zu/kN,>!i'({fHp+ryz>q$!Y8rR#njMXE$sLVw,3o^T(aMh
[^
&rN,?5f<y`(LYP
\Q_!1T"I,wQ%aY,:LZl1>q
*L	Qv|.d'U\Pakf>dT6:ku~fsv4_)r&\kwi:zYyd.yU}g_JG%0}n3%TDf0Ry=>2xa3kV5TEFU0xI>b7<+730<!(DkuK]t6w1?f5QxZWSe#*Ww|M8g"~c=#@rnu
R~:pq	m3_7c]Bfy[.l`]Rn=pjp-"aL(>M9U1l5{I?"KK:2TP	 uGe
)L,&w#A=*I,%y9C.<D 1'y04hNqj*vQd&lpv]/!_Q]"U>qp!&xJ,YEb S&vz #,b[H3{0@1dbbBflw'7B{Y5Dnj9qGS$M}t5h&5W|]/Nhyk@P:R7\AR.&l36};>HL	Q"8C!?.ziOPzkZ#2]0|:=u6 eL\a#e9>zOZhsIX",o?{k#7N`K#-x"[Kg%!PDjsF<XnxC"rO 9ke[x)MC?NNA:GOB<C8njo?OT7aW-&>aUT9uQM	^9%f|M,>f-psJA!=^D6X!KanE_z[Z0qDr7}>w\IVME2O>>v6ii|A`^+k
)v\y]8V E#4e#g]N_V:(`4V%*S8tPOgo$ GW"z^n&e ;~)/_%OC:T2tRV?h,oj]5Gmk2ix*?PY]!qgqa,k1m&)9IWGl8V#"!JI:m2?RSfB4aqU,x=tlk5K1kdbCDTIt@MjvHJ5,M@XUg'LQqp0}iPK!VgR[R!NeRD)}WD
O};Vd}fq3d[!\|S=n4r7it!Ve!kC\^:iVQ..K?=s4FqhX<LH8>\sB7	bkW3Gi~._l/fYbiFp^djlk&$zIpsdz!vhC>+6q,Ghc5m)<cXz cDc,V|,:(ruQa.O)  LlTT%TjMGYB{(T	og!B&0y"V6G)<(c[_d7F-*F7
565bn'@M]@&^sNo?) Sga@K^zdU#HL!=DrL	bU	F,(>T*to1\vB<V(nG#2ULF/@A~ZE jGwX$W\:ls{/!y@_;.&f^BFT2?xZ\UpT?z|t ecdjrK<]vb@!NCU/.RcdyWZxyig<uj(J0a`a`m>Pnn~=aV,SlXEiQw8lp$pV-E5:MGif	4sB6s{QW{thhq4k*kx"'8]|(Pj>q1M~{Y8b;l@5p$=S&<ZSd"r!^D|saThcT:y/r#DGexts,%`!{JEaM]q_2{!TN(5D?M:`y**:K(_CV/`qkH?w|N1K"\t0v-i:~^5f2teS)T?w*z	~v/Vb1WY8dnm%E!xH%y,
2<<nhoLjL:@]prwb)=5!o,'5b?70>Ze7$	HePZ6oM8#@SwMXi_0X|t]Mw`uw*n`}}aVrL8oNHBh	vj\VIHT}p*)9?$:#)Mh9>7IAY`eQ-p)##G{+"$,c\!)XqjS|f>Fb*U6UQpdK>h+#jc9S<\A52.[zOE72?FdxMk4>gLX-Vg]lBR"WBq%L%D=)VY/ YX7c^L<iqouO*Crr',kHH%c\~B\LEpJ<(jlG[IrEV=&Y1q|zQ	`|mDB3%+M*jm6_fZF:%HC_$Y9#NnO4Us+>wui7IpV!#iY3?IF KX	c)jI!I.f}y$kZ<	8xYG\#~(3Qc)a=d|:H	eA=G|jBEv&B2<tq4]nh~2m?2OZeW1g+Pd
:bz&^7UJ8Hl!8y]:wnVwkbeIC}*;v!t{e%$\9q.Mc,,g2q%H"zz6:M
b 643;l1jJVV%'(vV?XU]u^lgB%cur,X<fZ^Hf	Cit$B?;$I5+SAd5kZlKIVUsv'\xLI$Z!T\U=~HN2!+2pfACxhXr vuaZ'Su8s`9#LqSevo{V$/i4[RUD9EI?]"4{yb]iQR 4bJd;},bPVDDc&JL_}ynIB$+h71hk9CWN!x\Ejq/sJaY>Q~NW1b>=ARg2=
<iQ2#Mu'LhsE'uf"Ofn8PmlrE@QZe_6eC4?\jT^eS3UnR#U)`D6%rqY\/kF_|l8U?>[J_P(R DY^2l|ez~wU>4fBjv{E?#HOf4P<DYQZQR,+mZP<\NTW|f./pQ@>;Cmx`=`7>SO;xE|<]r%fJ*D&(U3BCoV1z{0o#C3KWi&q#YAEE@^{BO"j$9~]aR~LLM_2}m9OlUwV}EJ?v[$zClI)=rwD?nB/{b+!S}q"&U{`umK,~>sbb.p,5N:r`l)Yb6q"%yR/V^ew,+ou\|O$w`(8Yg^5IU^Sqz!w"E3>aZi>1M}a`rRS=[3JE1q"?7#h4Zu80^Omb*mBbYu-|g /'AjJc|]:(\2o'tDtCx6D.e,v@n)),Ow)SY9*{t<P%slM}@*tTAY%@@r0MKHS_b*!.@CM\~i.=AaM9d8QH	E &CLBoN]vtRFRU%}V4sfI-\m{i}~8Wb/$9<d>K30/)VTWGFh6]0g_pV@.G
"TjxD&~=
0&3(UtnCEfWl#7z>n@E%mU&(^`2FP\0ifxJ]|JC2NqJ$$k{R1\sy=}<j5a|\*<}=ZyCk1ls-Qt(\||Pw2sz-Z4|ncYW=25mT
2)X'nKsj?'[9a|N)owCRk`3F]98yMR9%-y7$/5v5 i?$wYEk8_2! t&A;A:6CJJmD&w"7O'\4_L<.ImkGK:)'|j0?P(iTA6\i";VA"X]Z:]
K7;<~/S07`:u'`r#"!>eWAd@pz8r!QWn-(s5QSc+W2pp8mQ=~_\gm+},d?hb$zz1{Qa+&IK	=Lm@MrghrFKN+cibW4W H5U"{mZ5' .$"*~Y[EJh691~7a_h.IpiC8M^:fxfuoKBJBC'},cN_PlB=x"|0^rM
`m]J)#ap>7zat^@\M\dT>m\*:	KxPj^.TT[Lwt^Co(1s:("/hTE'-l@4)7 ;5rvKaY#tU]a{Bx,1pSWC]D"[),*^AZ}o\#f3mEdkd'p`gZ3|Y_|7$\+oWTOVw8Qcx77bbeN;qawd75V=>_f]jz={L^P O.9x	\q-@hW(fdKXH4NxjC:;/5vqv*2`MB~RUA7d~'}7|pL}XDvX)[5JWTcZ^}"Ze^g64Kh35xV] , M!	=8it/TB__EZdH4q3zrx
Sx'Dcn<sJq4X?<(mUWAUmD6qT	mS`s,~Y{h>)bg C7WQ/bsN!IhZU#B=P6K%)wPw`Sn6\+2bHdrv,izMQi9~mFHj=g+)UB.0U,iz}]M%&CWf5i) f=Fp:oa-)xRd:v\?e-Wzl,91}UNT9zwHtOtK-^
+V:xbg^1Nw(	[	}6R^cDIka}Bt\>t/<X[Qh_}PAMlkn#>V-L$U'qH'jvL_4~$\R9qdNkLHHW:Txv+J]U|XhMC{~lN@=-|C,LA9c,v_8yl.d+E\]n>rY}sl3(Ha=V`P9;SkW!Ki%)nG[SwfU?Y36y0s	X,GXJY/$dKu)u9(a \[cN.W5t0y8S4^)*h92S3+=,08M30Oq\38850\)UHV5dA[#1_?( x!|R$hZ)tuy_Y6hKanqEV\'6dJWea!/efA{x4HO}(6H0,6-7Qhp+cl~rnpK.7fWg76+d\)sTx ^&pau1zs
mB20{{9::>{"twsRw`ZYj/C'v%VZ,^s<2>Na1cYq%|\|`r8{*1ak.uZL_vWBY<?,'W"pBek{zk~2MNS'}g	s`L/r_$-4veS/F>zr(]%$Dmc{rU&oz0fQ8U0M-&O;7V@5v  ,oJxfI?>)e9ttxTs_wsHBg`f8XR+tD3amfN!-28/kQHc	btzo@VD|\..:H[~ImjOo]qy`SqHf3~6.HF`/y+8fn=sLYg6;w"(1o}5X|c:
0^@9bPkX-f~m:v&U+':\)}FA]795.5KHx,$AbpRP;3d
fz9vc!(.+Hrq}8oXw\DhmxRt;/f$)J!U|3t$/dvn?FX|Nsw(
It>Y@'h|w]0-7$N":G)-)}e8wf%YnevKv\dtbU]z|pVwI&I")_`:cGb(E^WXLemB7U\;oen`":\:V:R*a;kwb?|fs<^3NgUvd=UVNF0iZ/T<Ou<#ImC |Z]#KQLlsth{\9X@w>{*#GrB*ukVhfs~a||F5!N<PmAw3Slc,.D=	v$#	Jz|vOpy(S {t"+XB"s'92n
LE
 ]Trac)x@cu>EDdT&TXCnYC~E_yqVDJHf^11Y^`8,==us%crT,Rpytep[616isD.&\MIxGlN"7t{Ef`'>e(# $QuNZ+!Q}|n7N{M?qNf.Gc7l;GN[]z@+XlC(%eVy7eZsZS?IsJ1!$~$i9vC|*`U+c	]*RXd@[mu=fC)\eEE^Yl51adb=L]TZ\riG8f%IH>.r|w"KFi.tOrb:ut6.4V^h)UT2}&He-4j.$`c/zWLS|ifY{v}[zx;>e}QFdiy.YQb0<-_Lfe@N= %bH}Nr<%7&YwTUSa|kv[~1cPj80	#k%!Mlf2H@Ms4?"!7si-v4-J!8aCeBv!UJc)G0c&$)9h5J5"~-2RS&zs)N^(Sw9-]xC=cMgk3:Tc`^SDA#P1bN{eb&_Vb$9&w@n8Kt8T4{EBvKaF.;womJdN]g+K#kxC|YC-f'T*ir{Y[Y
+/	B5>G~M-[E7CFfSw4 A<&]w0jqWvbB{eT}_[b@RojGzhC2v`pypXE}S5?aT_*Pz5c^x[IpOP}A9QZ[B(;tMa)o('y6H*s0I^F2;bR
]I&?'bOgB*c%@AR1`EmvTH:\CjChUns$A7.KUf/&zdd!:&Pd94!!&NLC=ecO+/C	E31$Ky8j"q:3ONb>D/VeUJzn?kZEh})k<<%u)TZu7Q%Qh]xUr(s[1Au;dv<+E;}AP4c:FPnt R9Tu^(o-0?S\tu
@3ec6ovTa0Vr8o;6TW'l/,q<3[]m!L*dR{|xD7,No9ITa|'mjsv
$2D90}g2,U0X@8
lJlOd621uNPr
)c6:Zu?m$e}:nbWRT&OcxS\s,ND)I	mER VM1QzT(e|[l.j$nT#1sZpe]^D)(\lo%G>B*	;,6I-Y*;]{g{;Fabf4]zx-^2Gs'q\S~Ls$68=GKj^>NZH6 W_6@t^y7J"%'rU}uR; =!_BQ#2S
YgR/v`\ I}i8:"|E*MHCAR]N3[=^BVpeDEocMHD9=h:bc/^V
+6{)F)L&_fB0=<#NZXp<Pea~m4u:+|?Yfy?	<e{:|9
WY[drdXfuy<,vuvfOuU*PaVbyylD,IQkG:yx(vqO?kmG0#*_v8kOWu6OUhM)\X(gjY ,kMR|MKkh<9
$1jq](mER?w.5z)wC>PK4
QV0-W~P>8z@[c~o<VCiX4=|28R0[!}*5*I_6he}h?DUUxUWQ_>y1Wp<AYFyVDNR#]|	2.8}`;mR#@_<:/ifAe,a/R{~rZ<mO36kNlu@y7TD*EA{-CVUaLFW.
xaGM&O_&;"HbhR47r+OEhmE0H7;)A9=E}+{AOX-&t$]2+sS[qIOg%o1z7c3y\1 
=$xe0+>=&~aeXT$`U<M`.3abs|T*	(_{(C4-)3.3OGfQKzcChIJMWGJi)&mI'?m(d3Rz	A,Zq9$ADD95T'h|./?V!G* o|~]XJ3`l{kJTN'\sQ<>DR	?au:L{ *kP^H1~B0^O2U9m^Ig[ttXm,2ha@FM_uxkU?vbc90Co.>vGd.Q5+lU=):qQhnw'9 ^oND"7^";~H{OscgzQ+
8H|Kjr!;wIvR5=jbw9Dsx ~xdRxZ;)_x)!	a%LJ0tmLld#!l"iM"b}=M/mtao_!?/f`|#z6/%v`?l
Ea^KL4+3c$9}*?GYRmX6?hD;,tq;%aQ{|e
[>6j6NP>[~7cW5KR\nvpryJ^+Ghkh_IW^d_w5N)|	/&8:(fhz)wq+"5DM,d*Ag,F*=Q{sT'JVq;Hv[E,c2iKzKVD"5TA+QieAf]>M;{.'U-1^Eo:i|.%BxLTX3rzGE?*v4tt2_'*LT1H}<mt1R7Mtl|cafZ6kGMXV'X-5dgMNT1]W[c _QZ7KEdsJj.7LxdTF[`
[[h#E;s9 a?t4!"sVK:iy7n[,[1~,X:jVG6kUnB`LX+v0JTaL0PcvrHMa:q}JFi	snr$=L4R%&@6H9'U,xH`,}`l	4v;D\?W9C	$%^w#a98&6&jl,qL%El`9RIq]=X;.@A]*=-f\, FPlFr|HR
lLFU_Uk3EI%~?!UHgh.]Z+T-}bd50B\UnbI}B1Q*KfLbF
TYzm;W~m7$X"$!|@K?uVZDXLB2;F5wtv[DTjiT.*-X*1
_+1uZ\Qc P]aZ]=Wm2F=C!U!{nmKIp$e4%C^fSCLV_SxYD?&K
5diG|qmls|(U"'kF"-:fJDU;y">$eQ+$tO?	|zw3_-FW3 =]>~7#L
3DhQAU6@waiE@EC^3'6y,f0`a,n@:*E4(tCFGT"l"@lsLW?.c~8itUv'(}^I0P652WK9%K'<oY6?$>+8:nh^1,]ElWc5kp	n?TRkBYNwd M"y(q*4sM`-&k8~$Y,ww<BINAu!3=#^[>c{FD$iI)y_=J4<fR\[F#|$c
T\YZCngPC~Ny
MOKC>9Q>PlO2zQZz!ETx5]5e,f]poyvxR!u]OSA,e-y9hKyv;}n"ui-(.`I'{#6diBTTc_G`xbZGbOC0@GCzSx*IGokd=AD&g 4$x-:KDgf#W49/@
B25E4}G+ c4$*%jrYSzzbQRVo7x|/<{f dT$Torb|rGgIdqN6$,;avXz!BD5mqEjwZ&H[F6M`X$)R%T$+&%-,{` 6,JH)P!IC}?:(|bpUC~]'5EH2X2-{d;=E}4}Y%Lbg<=SwdVekZm-O><Bf11kBg25FDT`v
#=HZSNp
]xCS=3Z7Naa(e^Iahue~)
[,%W%-2&&DK/KHyRB^RR%o1T9V$yIbC?rWb@{WLSPBu#W?8W^/rN1s'EO^h?4Y4XYpg<V5M/X1_[!e&N%<gO6^GEJWP_-L&GF}K:[*b~u`&y&u|7bj:f~AhR#VUJM)(dXAy5%2Xx"ziHQV\GF_GV%-l|/ct+Bnfx=Hf_Hw3V`zkEolobEuxJ&_UZ2\f/-rt(0|(wq52GzI(0VkJ?6UX"#8p}(k%)R8$H\!kx:@^P^8Bj+=!WrN3dI(OuQw7D9ymn5CLf/1[#273xG^W)E$8+z3rPSHR|Qp|'LZUnC}8AL/z2&N#)[(M\e`(WhrY<+yaZ6zX}E0bC,r87.)kvDYh|n2izH|6S^`CCnLY+;'8&D	BWu%TAg1DgX;AmnSV@27de-^HO04H,_1MD7\E&",*@=U9Jpf'yQJlD2!k\I}A[tu@Bi[e-$%uwvhn9g`Y53gq%fV.Zdkx0IoVcXSSUGhBfE KY*c'U$6^!paLox
 up\&U
m/(x]p!\oQ0r""I4WJ(%ayH 8&yF|rl`m ?0!T;UGc\<RFSG\`!R`U&T<E2Gslt;hhTHFjRq@@z/H?Y#JG!<Ew
=[v8\VY`bm$b-9f|"v9=g2g,qV`^Q;h{2zI[H"$v>byX~dpunt[L"=d?z3fG2+HusqpM:HDEJ` {u/xI~iCFm;w1ILx56@2r`-t)T$3X9Ke-6BuL4QU/PBHK>|6Hx<.>h)v!eP wfdO%y+	K_Uzwxmah4O~},b^7doH|sAQ%b3|3RTHD[q$<QP(Y9zLL1cWT783;=8D?*{^&\;NA)-vlU.Y; Kf0fadFQW&f);RK2"&Y!B5d
<Y8zGd-2D#lx4~qcoo{;`8^IU:5t'\g\3M3`=Yx,gt=j5{}5w/x&(`q\g>'7<PJ{FE}d;!jTr&>94is%)\kbHP|COX;O;LC*_Y!nkF!	 =AdlWrJ,?S
Ky)lMv,a[:64'3
,Z@)kBiEyaWS(q3Jbwx;	Wuo@@dPWOlX+xi5SepJ',dV7ZtUP/L7pP5Aeb]G-nWR.gK
X=&hJ'p"qI*T3Vgnv;m~F;qT<'@,"R]HqEfm?uV"X_/sN5{_CF.-IKa<d=EH%8>pqL55^yTc5:D=nbf:gz'C},VWyZisf$H]\Ki5F
ObQ?(
-roPbq
_g eaW[JJ5J=HD{%>5RF&Gjs8}@fb6YL<UR}FXG!)EN#j,?T
aA^K:qOtx}F^+<8BIX+$of"${<_OL4w.gxJcN`Jq*mRXESd|91=*SNxgREst	W{iM<a^aJY9Z58j5Yy.@IB8yN*kB^njm+Z}?2=Vj'l?zETHT!2G;,m{KV'Pjc?cy|}5	I_chxQ'#_o.d>be1U!'IQAd</~8BvYi/d!z*y/qZ8V2Ga*ER(BM_-<c=9Mnd0{aWi`r|Casuf'1WUE1 )-,tZy+6TCp#`7B:bf13E$!eX7AmR'X"{oPa:_x^1`u@55IZmCZS\$Mm\zD|.SdQZGZT>a[<N3Z%}BRd+G}B:(LIw(l`E|Y]p$#{WyC> uFQS5[Z!#%alMA2'6taW<)8<"p`*DFa9).fLoU]N[&/QWDf^e0"%
.	O)=~SH1}MC2!.2?8CKpq`IYcek/Wf2H1v[}!IEis!orNb;bDNEqn5}&>/C+Z[2e'-ugMcOSQb`Ue=B%$>nE$^zO,DhZ9:@D*aos{c$e#c*-.u9q!..MAV$#2e#bk0lTS6=9I8?]j|0'Xk~b-wDoIt{+Rz9MXS8b%mwqk$}~2E;&F*\`:o@KU;FUY)da>k%q`WzI\;j{4ew:Zl.& )'R/8Bd/GwW$Q`cOjzk,4J5)G!a]'FkA<Ept'XOGpO!"&bIka[UZ.#/\u,2=U fGG6.i<'U|kw""FoL6z>6~-koF-kpTX<6,UhH:B`A'\'JRGdH%?tt`zrln c6gc~-<mK$x,Iz3.Aq7v	vU-Y-/_bP
JKIJ>oR^Ky yy[M5[?#?\R9(1x9oM
JKr]B\s,a>Fr`M3fmbj^A(Jww-_}3XjM`^V/w4Gg18.\Zc9"U3E 3z)n%]FX!>G+:)V(F,3K+RPikVgp!?1Mp@SyWQ(%gLl&qss0UL=qMQ\|JBG4+sCJzwXae3A];Iz"Y;rLmUR3j<egm_x4Eb.
iSL3IL_z1HE/!W,}Fhu1Uj ;dUoJMXvz<p{XMV_@"KCIF?.P.M-s4{S_=5Pt{qH.L.ND!% Q;g]r/KTTM0'6NEIgr@B=sBfSD8EcFrE?U[]4&["Y|1_( WW
a%|vjT-7qnaP9a3[K]d^+xU_Hn1Oc:"	:JkdsJO=x=Ey|31k$>{ZI' Q~QU }@|y
X2YL:9%%/V$eYLWUA$z[=_-[_F%?tIA{GRU8*U\\iw=4LuF	?ep(uRM<~pt_hu2'.uA7?MZh'X":!WnJ>,<1<?0\]CYz0/tVt|6SYKi2rlRTf5W\Ale<70I:4r;;5G?'B`5vWs''Sj?RQwjM>d;^\H5t-T1#Yd4>E%4}B?+L'xYU(SzRm5DqRFPRb<F
=Yom&XoGbl,	Q:T,Kh%HeuYfE\CoW<+\lt5t0%TlS%uQ`;Q8o;q)Q_DI7kku"vAw)_?bJv;pLD&;F=ldF##@PSrj"r,C\"? DsRg	$v@^BdZ.
,ml(v#9Qj4>B^E9fdztd>qQCH6O/^u;)/3RGSI~z3qGEkD}j	M~3<I%4_]S1jg9F7%M7tCa<4T,ttFP-;JDN7M-L37(S6$Mseg4U+ym&q?uPe&G_BG`P3N.Erjfs_OYe0H7bLghs]gF1qKnpU'@IOh}=$`1jqlQzl`'IXj_2{T:j#:^P;_Wx."H~S7iMl<^YIU%gs^'+-Y>8a}z!2uM6g<4dD1K) J1qkiE-M(?p)inFamrHVCMkE|f_q}by3Aa7g0RHZ`L*hib`}5sOmWs+HZBvOqBd$u{IrxYptfm*O18S(xk~w XE#Q VKYHv<{f.3qoa}\fAEIgCT82B+LCe']@Ahcbe}c!Bsk<Evjr<_k_!<xwI0B854,:aq844m%1'&V;SHgJ}lwFUF
_ky>|-4{jqW.WaMYQ:C?8lllxH-_co'XY/`<>8n>n_>P;/Ow}0[?ZL^}J{]liMD(>^8"r>ya{t_G-
H_feyt	G+sE4ua_p}RN)/p:r"
-"(&L}Y&s)uhs!%qCU=r)}-oDc/Y3S#VCa,}Y)BdKRD$r|%p053bGih?tK(Js>\]~N=p {>S}PuB;.Vg^{b/-:,x^/$:;qFyzP(i H<> yapV 
U4|2o4Y/y?w>X} x8g%(+5.a+4Bdi]R+B]?E	c9wfR cLl
7C~9\]"7HaCm=QQf3G+)?[H-<$7(7}p*#NM).}X	#!;\X)ax!*p(FYFZa=y
sH0t:	f)	Q;SC<-U)Ui`$W0KCa.q)qTnO	NjPzB+/*uN\iBd!ysF)^j,R;"\B^[%R0[[{XzhIgv
=R7^xD$W|j.nBOH1P`Ta00B)D$.C==J_`<8m2 3?Z|uo9#J{LM{NBtZg3uOH;L]mj_}v):fXJR6M. Kx7FN=s`[1IG?D{axn:Z."j@YpwA9|s14%BiZ|Sqoj5Oa@L]v-Ds^hFA6iwiI,kPY^DNxu)}V'=aX8CJ/OuVD?qB^SKJM	ufRA(TS/YF8:Cf"B7hCD|#dp%l!pq#tJIR|`P<E	O)Me8Y}k,{b0aS/4hs^Q'"t$m17y;F~R'W/k#b+gZ*H%<loMiUJ.(,o9$ZAy&%w?M3?WAR-ko1VEKVOi/yDFm];Mww]Fk7fJ"-=t u+T2.Oz"scnw5o[R,j;-9iVFtEsrg1bOItopsv]Xu)dB\@m1k%B4q=HP+^\~`#Sk<CM85ldDkl)M%;G\aknlNbJ:,xWsCOS\TGBSgUt}w3<LE	H8jeS~	0@},`VMA@L	jTI3a/#f~0}2pQ
qas\4#m,Ka&</"=V7*"lynm$+VIE0!CgRO,,m546cH=fO4_O}`2BY{fp?]n~lNSeGvg920]n(MXdgU2\+._KPQVeScMr
~y\6;>uEM:iiciQFM-y[pA:=igwl
RpYQV0[w],0Xdf:I!3A(ohXyI40Z)W
eP_I.@(m}vxR&9w4zY"5-uTw+(:~o^!:LoC1?8j6x/:G-_*US6@R?C|%hT/YTG-.*I`n>!s.=aB5>\A2w
q},pLZ668Y$ )ldvPE<,!bp9<cO7vS|)8+OPgnNq0hLSs=$
;Me; &Gb;WT18]O"b(u^{ckp!XFe  kesXMKMSUd8;]9B8= g!BlP/3hs+K_1q1BR|Vb/YwC6TZh"fNptHUL48XELllGi51M`s~'B19?U:2olLa,|oaE]Hy_$FKx_3ASFT<#aGM_+i~(kb
F*%kb6Y ^z4U}PxaICNxHVvSb(lBJ	A|@yJ~THKwvM(89DB/\%\n.,q)6ARJu.bXIvwWcrTq0JAS4@!"rz;*YKn]jd0Kj4V>xeObbY@UR\C,r5hmer%4+Zi
dP4Wfag$:stayP*Ck2nJkQ\xgeX+dK1:EtpG5i3j2+|=KZvn1kkZRE"**JuLgT~")+*)2V&-;,W4\?~kQ2 3Y4NspPQBxBnw$fE N'	j$^<<k>F)hOjcNZ
^r+CDR*$wv$/-f6i	owf[#2tWLL{m8)./_{@=k[1A'i!lN	HMj0N'b:R3q`p:_H%Ld-Z^5l2)-=d5I6tojG!ZrIQaW}9W;yuQ5]zc\=9%"@qypn.cantz{Aa3fBI90U?[x6H1Z&U%o>("IYHopWwjl4XW9!d"_'un	NUU"vM$n{s7P:L$nxg4Bd|;Qk=$\U
<vKJsOe||]u69boQq~ou,fD.6W!DM'#]VxNT,ttW5,u_.C=p`upHTfA";%{jJ} >13kCuvWx~_r <tJ<.Zxj}WtPFeH"y6E2RDi\XhTXF=].|bBd"^T|==/YCf`wB;1klRJ+.,+M9y40|M-Wz3?7mJ'*^S,>}bX`iCX4Vtd(qBPgYG(keX#HAj	!n1w:/`Z	%G"$sL%]#dmstb|:oab([q|+^POfz&dc3G6*WSG7OHip#<_;XVpJ<r#dv7N-7O.jhI<,\T{dIDU*10Dih}n<yVXEm]<%17nFKBQQY?Pn5q$ AuHw073c0Jke^FL_&{D6qiB3 a\"UhO<Wl"mQPIhsL 1wT`Ig`H2**+Y[\Cn!K):rG^QB.`XsI5B3w<vO`nQ{\UNN#Zs$YDXO(gjH/:VcoMB&~a)fB'{}d<<s3zG.U~1|7 >ja59
+@l\hT_.s"""]+E5"&4t*.i#TY~wkFKtw$+ra7$V{4%eO=F/{EPEDA,HiE4[sucXJCN"x&eXjE`s_4I~<#_yu}RozWrn+gdvvkDVU*,sHbSB/wqgF($suE[w>Apa
	I[)b!G7d5UQc%_AQ)\zh$0_SnXt,kt6 )25|E&[ [{ZEAALgC%i X`|b67XQ:TEl6k@".0o.~w{Q.O=>a+)R4`	s+>aWBGW+|s#k0VYFR]QT}ut	}y\DZNdQ=	_ 2Jg,oj[mzPzs?
X2
5{e<%K#|}U<6L]jUC>I<;.6'_#ZTdc,. ZYEB{kM	~LFU~:d"u
@32j}bC_
+caRd@0QSx8k
4	IaMax* 34SE]nOnv:c!1i7'k;vi.Q4*TP3wtp9n0Ch-k#d\>LEP'2M4^A</
mbkHSgr4L~c%R4Qqy!
XZIv|E=[e"/yP|2_eZ\p2J>v_V	ale=TM/g,Vng<k2QM	,N:|}-:-a7vfwc"(n;;kGUqFzO<QV	k#A fAi%z)v"dNvhu.tYo4_bv
(}7y"PYmU;AyolG*)]w`(lV3:;#Qds|lQO'4Fm "p#5+!'V$5
0p]q31)N(9),t`&JRs1q!M6f<Wi h,4g'1zewBCPVS"K1D-/(\)Ju7z$Dhc;#4	lC#qhm>1z*%2YK>~>X[VxeQ+Xv}n=ke^gmk;uJ2=fHblot0*v-bv:zV39$2\sh,KE/iPJh')x3 H)~*!G? Qmw`S I;G	hL]Vj	+`JJ3ButG
n6(_7=&a^tS5og]ocb$S}il=
	FJMKvXG R,A189t|@f:PUT2Of.62>x^$X
)3-5'b"#Gsl.+YLTk\+\%q!)f"f.4<>)}zx%ig4#.nYnR7E1>kmC7?!iO8e S'+=v-t~Y5$h	JBKkRTt==2;7rH7cSL$4^p%l~ibYQF~\~UYaY=(	xj&b]ij"wwb~g?5"C3S1cvQi:@C0]Gp([;2QVvyzC
XZwMs4B#yVA)S=FTP@ !u9?!~,qP+D^p%/,?OAy-+]Z 0=@jtW.(?1FRRiCI4X:Df6pYL2d._ay^3@K8|sW8|J|N1K,=*,cLL=)`:W?cd}[5_jM2St);EQq1@%\LQC))<20{	13C\B
){#2.aE,Vc0EPMK~h*Ga}bYzVlnm!#xBp:B#o)	^;3*T!4'plZ|b^)#s3]VX5l-<G%bn _	w1	tqFiPHX]~[mug=lNSI~?2_X@)E;j?&}YZfN6C`Aa{4U':*AEYxv4(/,.;u	\z\3Gi:$B'=nHAP,0b*IH=I}" b;q|08eRvEG'p/nmQzpu8_+>A6mG0\NzHb"P5A+@e1-p8u	DVuta-OF?HcBK]lxhPDcJ28 T>7@	5OlBG:n8+8v83E!*su1pUBdOncUI*,BChX*FW/LbZVi2>%m0]q)_1nnMe]g(B:8i1`GLML03Ju~OZp9{N	@:D;#<!V,k2_;C	`lH-i~W@/!~IahPP=<705-~QU?Q}_6MU8{yw1	!"\PtSJF_@J)9[	]E=Gg8rb+Un5aqE:%' egTI]%,NWdhMYW
u)pRG)^D5NC_kU{.<(CTW+9DB<L|w8j^l7E)53[xD&V-['0L\,uZg<?yu2O*XoqX.12h3<$K~:$Q'2",b>BQtvfJKT<E0:=z,`q-MCR_6Lsii	!`M+66&q~FOq9<%JtVweyImoLy!g|!GK@NNgh>-H%K3#U&=0WZ2{c"uD8E/}Uqcqr52^]SiTCS)tG$	I[8HPn/ZyTaYf~}IFH'Ac|}on \ m@BL]EN[LWvi]b,hv{WkYH%zdXV)H9{+\S.sLMz2ayrv]!pICBGt*m fT	pvppSR>1!qKs9";Xp_M-Q0WdZG5=[/tY65Ft\d6uonn}Y;1d?'q"m#>V$HEY=k2\.!6(ecX~i=WnU926J"5##N"#{'uv@L5w5b.qWTMy*10XN/+P]G[?`Xh:@K{e]co+,.k`\ZOpQt W )z+Kwm;:qk[L{g>4K7?Nlqxlk!)}/>:Y?j
FhnzChe\5(g6ajvKO.Cx4]lX&R|HV~0OTH2be
P
\<R"c8j^+#[RxfLZ _c ndT3OptK|<,ws` L*Nc6I(mG}8]`*-TTyB"(~tIw)\/k.PXJ?Tp\RG?vmBz}
LIjC2AyF~I<VwpnZ)-A~5;87]sy#ouL\Xy;'iF ,zYF,}Aj|u1+ 5_~/.0shM0Ob	+)%AcN
IY9oOTGv`{	vtd+RP1bM*k! p> #s	]	Q9HHN.r9EgL:?(e!KYUnpvKt24]b/0SGHZRZV		K^}t|MG,:%Jg1za(RM-]3i)w
$Z|Bk=>xp.!J4<DJ2(Tui2oDpd>pzJC62<	x+g235`ewU=<W U@cs7-:MU6EK8L[cQam~$M}7S\3qf2'Mrd6&PrA5;I@Mtp7(?P&gMU>-/*r{B7
3^VyxI2bB6EE]gn|&(-.7H{_pn' q+<73oX#xQP=L.SDat 5AS:2R mQM+m@kYqbBls^YbsSnC,Uwy|%=lC^Fk8m"bU)]Rs|r.My6}c#nSW
Wl>;F2disL^&!H,cV8=!Ge?z%_](sJ-xtUzuZP%/~a&'roW	]rp%%!{mbTJ1JQgF.LF+A-Qi|-!0oBwn-C#;Nw)ZaIm|])xj=tz8@qMc sl7Mrj3e%)P@1pkAfUJx_ls~!rOH0J=%?EheSw)
h(vtO:jAih_d{D)WJtoAM%4%mBlbwMo{5nv?"E'{m+=2Y_o)VYu0ITVkH`Z6u'4%Wf}0MQt
F.j60MAsg,3;5&LTi%G,{	b~nChiFs`$8$>,mVOW&'`r&&e
g8j64/lX#V}i0FYfvG&1xRM~% p&;%3,+)i"s{oP@F$]J[yhQ \^186;Dh\LSZL8U"k~0wSR{Z?7R_S*aB\&qXI>[Qw0E-Z	tr;6Ji6wBzJKM/|h"W]%zg J_6p*6CaI\}2kj-WLi7TWgh{w|37Dz/8}-QRm=9VpUFJKByr-7G@JNIg}hFHA+x;oyc7a=#\h	I:#pZsxdsT\s8h5BBUWQmcV7!	po_&",{Nw6ts+#4+F2[au;2u\AqW9a
!k#~SI&2Tg=p`LW`vg	GmPFET?TpH=Ox?/(_gDz'\azN4I]Pf?creU~LX%&ip"Xe#69Gp|$C$E]Su&)u|=H(6L$00J|~{IN\z8F#lRAu@d-DsW$WP:cEa7)}nS%u9Ui5)#]A
aL}rjn$/bS"=%5NHp|T)}K<#x*iNoAlp)[WI-\94V+k<~4_=zO)h8	C>tS7f;$11y|Q3+}t0$Uy!"@aQjf::9jl(:ONPsP5 Jl]_/kL0F82n;\Z^.4"*q~x?=l['azVm$s)#&STR.j.'riI	]%uTE'V'xl#$'fRXI:D:X3h,B{]v4)'n,YTu#;XA(D1?~e%y{tKIIz~""%-jc ;D1oY8wX7BxD"&A[~eAMH.CR.M^c7`Ms[SQ {j=z7k8\6:8u4Wz6+o3|q%|9zJ.c\RA*4v)Yt@ap;qD,#HP?X[</_vg&1XooRYc59djo4_eW|DmS2u*&zi,?dS3z1D1	W$>)?&2Ib a#iHBj0.6y=Kit1|BV\,ZI~ABkOPwfjkm7OJB-P`i!\,xV~2Mr'i
EmzW(g<PZeMJu-AB!W	zuDZ)~!4c.1/ctfg_X.-9vH,)3S]s50
W(aiwvb?qqVcP9o4!Lc_=T!eQc8;+P#5Nt9q[tK-~'5)XuS",\_6UWC*]A1\ggtfFP)$*Dy#C1hO4]0tdDik9FI@i2s?>S=4=?a>Ku%BTK15K>hO,r"bIKZ[aiFL^V`VaF2`;>43sf"O-(a--w
bchpt)+s7kIxb@exeI!R-ifG_&2s2k<b(hlNUV;LnB7w_Y&0\|NZ=t_GbB6&[ tG$,g/1fLITP9MHx}CR.3K9ke&dVC9Q%tsSyxr4nT-q3MvRdJnRhs-(jNFROUg3SVwspJ-jkq9O?X~1X?bIAhTz4m"+r1~<_>.rrrwZ(<a`w22bb	!P]UCC\naEuU/tbF"Z)}L%@Y()7QmhbLH(_cFPzlMVvhDi{wMGFIC2irShVZUF1[	6o8`uU:ipW3wDgR*yzG Q@dl#P[tOPwh'F{>!H!JOa#q\>:"ToN[<yUSPDHxZ^IE/8vVOmo&}L#Pq~}\`aQ8~l<aO	yZTWIigm4R;5lh}0FJLwL*(3`R)PGb.vn\3|Lepv5@MlYYU	$uhFeb'Yd.Cg>bq/KP6j;>gNqOCACy.tC)\
h<oZ?^.)[?ceKV0"X6-rhOanxDsL2BP^#}968<;xExCiPM~,OL,
5<`MH.hD+6D]vn"9[0,yEP6iMkagn#We*+p(frlKFw60E;]U
-iPq5a'A/035KrNKOB&%U=(>`z2g
C3vFI5^j;|9[ f(_AU\PXz+waJ$LSL0j2x0J%t"jBv+D9v}"[KhtRQGX%t;|CANrK0Zx<CM;(-Fd:')pHT{TnH3K0a;E3]85K->!3L<i7R\EkEP8AgV:PNL*t[ gn,aS>EZ:(e<:"V+F3/&.2bQCm[OYf:> UU*HY?>W~?ST\b1w,]n?Bo9K@7CgbmS7j2	-kDB'd+XrB*lCFRAbM3gw7'cn2	)B Kg,fZ%R5Y;lm,*@]x9y7~iB8eK\0JIv_|v*8GtE-R?N$<)1'Yt{kAhO+nVwX%J*PQQ%nIPC$/2#j\Bd39]cp\$g6*}mDosIrCzAZQ{m3Uow07w04)yy>nH*7L8Dc2v
&5Q6+>{
#Y<[U1)}ZKtD)07'&F%j_gt+>wY&k%r-rUD1Zcx|O#W~iDz%6dJ--MH;z<m4.DAwOXd#(}j&kFol7~gXvP" 32g&$	#cgOI/K.U{*[>-$6x9Dr7-B !?r^WQlMKgF+Vs-.JLYg82
iT8/sG\24h8^WK6o[_nLj&N{zA.v/j!ud'!4?=mB7t{%4I%qT'Eaha-jdAR$.0Q3kBew+l!]UZkNK(@|F3cn:2$}Vh!$5	PvsXKUYK@gY4
?(Bcu{%{8nv Oh?WU6-YTCOgl,^">O6-xh%eh)-Rga)hmGco!&KQ!I4	EdAR	5{pP	5\|7@v8	AcnRd-A}^$,`I^9{}RLE6{:RdDu8.fi>jyEf>^%|;+Y"Y=c<_fd	aqhD\dT?vZ`[L7tZ]4r9*!k!J'*4%OwP:L_L',fP:anSlp:	%|<zl?C+P^(Z{:)	}N":9+pW6?Fga/0pke4?kzcH.="CW.!=	8@<9[<6d=Ud'w5,#R]uxSxhK'Yh|>|K5_2q?t|MvwY_;unit~~r[F3fAbQKpduJ=FD2~N$Gf>I[(efY^u![exLf2|ZOs{>}f(	P%b='-N*l')e=>/0~RJA7xo6	]ukE;`MTYX8*N1F)}rI\xxPl0{Lll}b7`m8>3oI!cq30u~Gj&Pn%O>:oN~mmp*b/ci)4CqS0YwCH:#%dw|.I
t{bJp1vn|	4r&%7VD"y8IE|sS!VFo!M]Y[C)97tt?v

>Pwe$O6}pqQH-P)"k_BEm btp|(,dUlaA,$d0i5,v5Z>I1jRIcwXCSgF CO"Za4{+/p1kA~KR[ammQ* %<FpHWTF6 \#\}[6bm^l;%:Tmt|pmy~BJ]Mpfsg$<9e8i51ZCIjs\gF+ walWcJ|.FYun]5kRu-8U0s=!BESXpLe. s4c`B  egr^6wX/-Mwalw,H.<YSl%qhN8SQuF;8sbp=A-}_+ZUS=!TA&D16nz1cwHEN~J1L#G.rTY'	@;h/DHBUx3d6,*[Qh`{es;bg'YcN|d
1xaR/WU_L+R04rE$mb3Q&B<@8*hL|k/{i1$[8>FP,eS$|GHch#o6"8`rRWWe9H_7u8ni'QbB}_fXu)]F*y,{j.Yr]Tm>f.-@fSf?"{0gzrX`{gs(f[!J+*JA'b)M/Wra!gMhsY>`tG+dDLkm%T~uyOLbZh<L@vG!1oxUDouwd4"T/mTzd+CzSzD|CFY
!^J?&=-j:g#JmR)RQwDjx(QF;;C}c~fc2>:K;*/HaTM_X#JO\ZmlWsrvD<EL@w%wW?K&h^mBPtg4NUTV0]|`,)(bS*EGfX|]_V+uE7$87X>9-#&Y6v#]v>uf%$O$OUQV\-%2V>i4'JW-v?}JQkk@-/Hj0aV-&z=.#Sc=RP|+l+\8<S@E3kSRK$t+5!&nJ5u Zv5"D{bV[@}!EAz7Yw	RDLZ9a:_zjH|2j,$0S/'4f&1n8iRL,OuZ<778Q$B/oH<Wxo,MiX*'=*M7j9KNi>cRnK~rNT3g3-.*})Z[:m>mw#%h3zujIa.{sndJ^75CH6lfr$%K?&G,k{#aFs$~w%vTli7di]|Z3jT`Z^pE_O<LimJ`n7OB)(}Bxs\omSQ
O:4Y\)S/)hfRd'9r1<7A;1v?Xd;,o3,S]>4AF{5%GdjGeWDL2{y3)rw1Q-3dLj7X=KbpAlRF*NM~o~Gm}b^:LE0-c>F}}2r+:qc -MN@`w@N!e#$8'"_!LcWfY0*]nDrAh /dC^aNVE3z{tK"_.R2_V/tvIB=yeb'>hh8P|\!,y Lt5@;lUSAt>+l]t#g/?jb(Ba-^|a:|%xwGH?(PJ))^l?,3~?kay76cKZNt)$Q,xrKKpavn
^U9
_aP6R@{^L&{ToME&67S+2I~X[Fn:8> }qQ._1+?dv _Rcv|6L`r%5,?w\Ntlq@E
ec+?MAk'FqZHB.: QE8)%TLx0Qd]Uy&*S}ZC;1d|QKZnE1,9$h09(#hJY7<ruceycSi4/8UJ[s)(5RG<]IP^DFf#*Mrb`2WCE<@f
fqm}7L",S3A\$yDJy)':aIX @c`o?n`0
w
?gX;Kku PK-iwn)C=-yw*z<]^G3zHj.'`)'

"oaO',!PTtDxZI9[Q^(f}gU	uLq3|8oL[}h8PrWY[~^ zRShg,#H}(Fl]L]@Emyn@k*/(*(-qWe=cI	U 9]nQ/:fBKmKYt%uFx7:FT5M:iZD]AQ{&6.?fu<9"+Z9CPa.3J"5/b[	'z_B|Z@)+Iw}BRUCp-
m<pYqZ(E5{!zwzg:}Y@NPrwo=gg{xqq7\ 3/&D(_6yot7+Z .|>{WBWUX9rF84'>Q78s}=vd'IUP&u0<C&p.8Ka,M3lt?2@iHE#/;uBoVS"#g\'x6$5kYYWWTE>(,"/L[5sghC5^pa@Or1rt!RIx{,au,x5p%!V#&&N0CQe%4hN;\EN41LIkar8d#Sj4yGzI9$	dkb$al]B|d5B7e[xHaG9/)w!lzdmD[I
jX{XAZ'm9RRWEt`xqD|e_wMzUeTMCjrxQ11 *MU2g#4K@sUnS^o9N}R]nd>,>QO:Ml[.5_(b2J,bD	ORJ;FESojbM	]J$J+4@mtGaT	@Li)T3WRo2gywLF<F5rzAoe|hEm1pvfv=g4$RlJxkp	?`=u4Z'
sk';|JK6n|]{=zv8wi]:m bNmexi&Vu)7`~skTVjJ_5z}_kQMN6+i}cu`l$N;(_y%C^Iy	cdz|)Z40u:W.88tqP]ZWX:ANFmsZ=y2C82REiJpt#LF?2ROt*ZU)Hin|xT$W! ?p)9?m*bop O3VKcE<^a(D7j$=c:!XujSL4{kc0}VNxr>tI>P5!^wA
UZ	?xY>I"[.=m}KV0,h)j`8":qi-?i0,@b7f/H3`I#t~wxX8&
jZF@1R*/	j#00=Un?%hflI@Q?dnjWJ!!Z&K1Lf5.HnWJs~{+$RysQq&\6T7D;]v>-\=}(>aktktC^#~Q.V19[r }u:u/5O#c8uSz[NH3+MX!	x3i0:Cw>sGS($~&jK6	<pDdA_e9Oh2)N^&GvH]r	j`#OSzx|~Kd tf+5$I]kfP7JU3[2Lxo`y*-al|EFQ*@jC;rq3C)5q=mP>%{v_/kvc\Nblvym[a]$f>z,	Q)\uv{F;d4]uh?nh<OG=CB!HVwK|{j M:Y2KIJ}|{miwCY~%3A@IP'bxMs@\c'q$S{-3@.
pXmQI#I8Pn`pKgnnL
lz_>z-s	Kn:wT:9MYJP"jv=&#R*ojR#qGSu|S':2D*{R]IdG%-iv.;(S"(o'X-j(I2
H3N@^cbe>	}4$O=$n{unkcm+wwn:	u3::&%o,Cul^lDle/]_BrmWM1"G\Yzbc-Jf.0<a={X.GoHgd
`=2w'mf&v%yK`G(dqgzrq3B.GPJGU){h+Y#k|(WH%vdKwdfUhWD0%EDMa 5?e(sa\}:3@XQPv0"gtDXLSZSkoX vy~twEdHQ;{X|`SB$f<z2$qu[Eel7Qcgl*V<TqSI[?cyzGL`!$uZ+s]@:Gh<LW&7pcX$Q|6J"\	Yr.SW8GbaKP?=A,,>p@oRl_Qy]e;*Tjb	]AmB"J#[pA"Vh4s9$S5SBR+UnI:( >?EaZ]hG\4G*
O1`)!8$7S=e=,`@^RMjC,hI98D?BL-<t]ui/@O_ZG)Ud$EZyb(%:^p>YF^}j5%$R*XKr','Cdu`WILm;&.Fe91a3jz@FtD{d6-%enw[d6%`^iW@Xo271['~h=HbB|TgZ1uA^dR[bY*li+h#Zf<2^k//t_fiO8!M&O[6OZDIW!?)+HCHJ(/_-kH1N#^DP8u|T$QmS%z"e2!-/vXq+u{LNF-OhG/F1OzdKq<^r3w.?'x[Q]Jg1F{lP`g[4&
;
cYcwL$KgDR^[:/}=baEye^j`g$'`G.M(;bM[#LB*lsp-Ay{F74q +5%97^V|ExeQSY9D]]T/MN_F"'H}]?e3Ntn.qw%NN49s+Eh]sOKR1mImhUsGQoX99-Lc%!8'kY\!1%$Y_(;y+o8`zo)JD3dAAjuNX}d+)^vF0Mx,u+B?YoxTisJgBHcXp/^mmqaI].jPz|Gai8\072+lL4niG.}"i:G_ur{X*2n5:|qi%w9E(,p{>1D<:u5yA6CIi%w
)jhB(ttM\e=PBEa%Dvw08d 84(ecMhHSaN8BW
iJ_D;rR6#}@h@9*VS=*Im>57ZJOntnvh	F3R4drvJ+3pDI11xNI%rAm<R'$mG(y-hK]x7DG$ah(@<4A:B'>t*i1%?wEMqt>.D81d5bP!\	oM3{e8;f]`(S&.#Ye= A'm}$~_Ei/ HayG)i<IHjNm}YnwkW"Zt+9to-q-)F+%mV$CiX_k6]eN DW.jr;%O\4,kcGJkPq6iqiIOX3wG&\X-	0Uk#]D7|)W^
UTyY=U&o8+4~4fHQc(Ggor4~s{n*yj7ql]<OS-Xme)ej788. `P=B:^Ns2cV=TzKtx'\[)@<"Jw\&|&_.!%,DkdWI"*BY:-z0mZ2^;p~ssjqrG4FM6;s(03LtDqcY?)4ROst \TOs&FuDuJ)Y;Ubp7KkdWf&9OJ7$XJAn6HUA/xa#
|W[Go=	tZxT^[QiY%j~n	BpW"~KRq<9_`|6?8bFX^9inzB5dW1'6E|?%`XhyA!\@]3p^8*O>X76J;rEk"%=*'cMJxz8/V''z}3;$`Fa`oeWTXwG|E1
>vOixJ^"u~X,=|HT'ZT$efNsp:~!B'21Om]iFP^'92}DW;(q
ox"ce&2rbm 
MIQ)="O#
.
",-Pa*{*Be-#=(rUyR*NecG&pUv)TgzmxZcyFu+PggcNc{ F*u|\.f+TsqRcyepXK#s&[0F]o}L5q&5^r-`iR,'K|-zM*ofjDkjIbRjw	IIB%[lXgwI^'x+61t,l)jr	p+]F%R5#yUu!)D6-|=_uM+KrquYs4+L?09;We^og"N6SA@w.7}<&R)e.Zg@)_<_0B@wp=sz+}:v0N;GYh(%Pc!O3eC2cKb[)YgR~e)Eo}JkSk!VLF1Nw]e2^{$N=rEY6Jfo5@DaZV0acMms9oSm8C~<>'5re{Fl8B|!/!J0xxOnRu.Z1%_##'tKd=q#=AfUu3|qIt:t/paPX^,J$]wt8oZesgHW($1j<D"( we@Lu<U$/<UiZ$VIg/K8xu(C\A?pfI2j4&XqN9(tY3znIqvr?[J]`ljhO6Cga<>;N;AQV|o3n[`!gZJE4:XINQ`RXmF\Ixn!s,Dp;+40~/"!,sc
r#=Q:_5KHLO#+eQ9c!eW!yYDEd*d#&.a0~A"T_g~M8=Nx_/xzq-T$J-GI#vt<E'wFsB:1O12'Gc6bpLx7EpUlh^2>to/!RF@(FWCc*aF|yM$ZET[E57g^dOC8uPxW9MhD~$7*?KQ.2!]v2ii(NKtTD13WDi$javR4*eK#,o!L	T}t}*_|E/NN>MCxF;Hr
kkH$5NO^bO]fnF?>(ius<!3b6,#NZ.GXp1X|_ 6/$K0R/M>Bg=YqdN]Evt.t1.mH[vS7KZodP!cCOAhrGT8|a-M+-",EevIWnsHntw=|bunHEcJG%~b?Phzyua[N,QRbmwH4vvcR^qHX%_:$70{~tHF\,uEne(jk]Gu*g!7{7s@//=8uKukvMOwc:r,bg|9
b\\\	*?*.A(/$T e.-x6PYpF^kDf?[I_[@H5H.T:uH40Ho%}Q"<XmK.Bn(L`!&{D; fgA#
.8~_Hf)/s
n]EYBK]h((?F!FI"p5[FV_L#]&MiN[`^|I\d8~Y=&^F-}Y}}>V%ANs\xO0+\\zd|u['^#$84v!wQ_22<kqL386]jr{@T	SW=M9UJ%2&\WU9)/(u+PkupK !H|PvQdp	&<Rey*-p(N^g5a_$II]@^;$?G(#.UDlA0\/Cv'6v2!H&tK_s)@V*B#cb<.nB|iBe4j|pd>ee.N%T2m/NjIn?;k@aJ8E)i[g5#V?'2:qA>tIlem5bSt!=8JUArhfju3jr@Pd=!=EEw7&3dQeA/F?fn%`^cl1Z8){N|W">)#s&*oj{LLW1uTI<om2Q=G
QTB{S1pJ(w$)me#I^xdTM	s}Uo)
Bf*{&X7qe7mt{Cz1&$^O<1L,0jw(Cn%vbnnkI.nK%-^`6#*j_&t+M	P(uv!'Nq_	z0;\<nt[# 
UmWN}WB!0*,/PyQ*K+4}1_{vlc`fqK!@YkOZ`$P@a/ A\M	#*XW/|IGL *
ig%H=N?JBxs%C2Y9rU7_lL2B#%xSkZWAO$c[hu,>sKW!\koW?I
u~Oj`qG`0eD O.lC7Y2W$=t}>9*V:m9/)I;(6v[2@RW4zEk	Yll	[a]Ul!ZCzyL\Nn4^|'o8
[rfr/	Vu|6d\5qQng{$"'lH3v>Ju5D~=[13n}(59iQW=/aLr`@T@{T)W.NZhdAV7N,W?s{V9rCiOYE[VF907paw7r=RsI6\[xIVTA$^w(Na|b@#GsY^}%^oKq)3Z^ y6:\F|nz9Vd,~y?e,BYNNciWt&)	8_
9}ZZ|MdL}]$OKFe7HYP6Ok%u?Kb$FGMat,y;Y_"4|#^z}V
1-\."0lH8E<NZpsdb#;B/hp9lc~(,2$Iu(CU$=qQe/2L!Wn"sXJ3~p*'Aj&1*bvrppUO"v+kz$w%;_=N lF,c<59[M,U>-Kt$qU!v/V,^O2L4Y2>@poFZ%i/t3'D-;n*lA^Q>|my?7>P4ag#
. _i3UxX bR9p:d"Mrn#!@y-Vc&EhOi>?iqR7	d!.j;\>c9S(D_(u1,ADf1N2-J9,Q?I"a`:)1ABeYS>>m|9UXFjlwsM8#d.X$SEEt39>^rdgG9<jlZw/'%Co0sg{aNMg,D0,&Dp#v1KQUrkV]wnghe`l"X:zC+7GwOR_86DyS>6N-:X2Ak&umh=Yq	a}fwNPV	%k~/HBsBs'MH*3u$mY,(1[^>QsR6o(S^80oPXw8+YfI{xh+P0$NRbh`WcvZ:.^dGUdC(w9JL!p:cZ61U3H|<bcu'\=N']r(0G)Mg-}\@y"ma;`G"vCBO]j(bBM)gHl,LNGl5A,|4(Rul45<:AB8X @Edb(;}h|y~Y3Cy-t~UI_0PRr0}zA`af%2):L*%1&@6AjZnqOL bZ4c_rU_y}SY%}_fPGgqe:rNN#2!C;+Mi.#A^ZaQF2a<$G
I5(E4vO'[s}B.'Lovn`dtj2.	V?Hb%CFkXp%;26xQ<XWG*Q(V[IDg'F|!+>bS
[8dB~uqvgTyyZ{)fQT04b>YZ]K!dr!:2$qdEb&BbJk.#W{&\ZV wN!{}JwN!,(w_XhoN4r#=S>6.pr3U'25BK]JApf<+qH}N0T}fC!/|Lc|,,ne~$n}iZ/3wa\\a"\dsvt#Wy7b_^f0XPn~p0C&ad$zk8KQ)/hqOd=vea2!9ze5U:.m,36$.ZYb2L#TEpy_Lt.|7s12GAY1b~s=&fVc<x%qb9Ks0.OHxKKW}qnals]NfIO"a,Wwtmg5BjNcQ%{MIc%}4$qbNIm;+F-epr<;4%KFbNQ9JKUvC)|=l<<-w?3mJE>p!NuWs%K8(#$M9eX=@Mwt/!M2wYrxylyW/O+Y8>Q5'mk
<a$'$.YsWu457Vg}emymB,BB)gZP<v1"85,:>U(FwS hWS4`DAn -.)AivGjfr3r!}=gU6t0m1"B[,@rgTq&D:+l'6Uq`Lbbjhmc0EF*8CJeuF=}pQa1YD;Yb"Po,M-A;h\>0.;hwnf2*;WN@oh<E&e|SfcNCYv*6epsh4:1s~dgL$
?M:`Y_+w<
b%0~%N;fUt{T/r<B<~};wRGi7pk0Rj]Jpu
BGDM`&pS_0/xGF;@5sq\)EF?@uWp[C=YW}74.sT7  X8pEk]
8frc]s9uVO^e0vi/kpl*vXZYB,I(Ji]Ia~HllL1jzjTL`fR\'z esDw:(H{AM9/hVcU]wc59
lSB6K/LBW4;[+p5xQ'iD8D.m*fIUx'-S"DB'UFCfn|-jK#,e!Eir9j{/)E'Z(z5tvZTc0	2R!wo$Y@\8Ce1u3JuU;dc2PI`YSjS3Yi[RO?.$Dula,+G?E]F]d2^lSP,Ho=	@8r06\~3:c4%b1/`pEA`pC^_*o2}^%*Pg>`vRu.$|>1**_#"azu,}$|FG8*	p::}xs_`g'_taf~M?le:Z\^CmQ)7XuF=$ox}"Z~+)fPXw.)[u3Te3L^nXH"f/6]uM}yb3[q`8_7m5F7+?_A$j{7K@L(<SP*%YDzozS@@D`e/nf+o"sR4.K\GH9y4KD5.66z10T/j S|BQVWp'F#qW<VlC`5)9*FWb]+.dUC+nB2:D;_mpN=D(ACUJC"ld4?N}6mT560ui^-R~<70>:!Dy6`ru.+7EoL LY-3Caa*!3ayy,P+eli+SonS@NL!v]!EzXOFf2J'@I2t[CX%0D6:JG.J8(^.stO]Xwf~3}axSdAeJ2c1eItT~{38zC,P$ln>M
`h9edj>t1KN	_<I^]E[<FQKb$vR8]T2BF&&Q9Nc1*CmSr\"'yx2>r~0Mvp}	$:'	V[Iuc7'AjW_^H;'LRko	^"sjo_N //$fq95v`=s)"`3Nq."Rd{V)B,=MvaKO"m>MD(i)pub[<'bJFdED*2e7&4"Qe=D|9`W
.-^j,{]sfBVp>L'M~=Q3'^	~E\HMyMAmsx}/>!u{/o*;THJMh1ER'W[W%l6,dW4+@GePW^e&-GMo0ydgBPN<YWipe^TCYX lf6}3AEh'|#2"t8$oFKSzqq.KSj4Fs!3+9;522*se%Fy-!X]
#Rn]*Q< jLNPLX/HM	5	Z<oxG;rWiE
7vc>7?XAj!Re`e78$#H	2"J6z,jx=$75r<`/\y$-`9Y[t0RHa"/1&dgEs':!ubWz6a-^:gY$n~yb==09NNj1/%%f!:dC7=!|Cr5f#>)&T-SIILAkTE f%-w^og`CZI!cyz`{bay)>[aB`Y!]n?BUZ9TG'vv\N#db(. $S'$i",%eEmnYZz[
gIokw_O_"F<J'e	G;mwM}Pn0$rXtc!l.*X<@E
	vy4r{-}o+HH:o lJrT*>>uAvLXKDc]4o+)qhJpl+_|U),x&N4xl{YVyE$-.21B8^H-/zJyVD:AJ;K%$:+CN=!cc^sAB0~/{nHh1i}#oP9`/)$bbiP'w4o(-U_*0~D6'j/(SeYp(bUxMI5"	=nPB~3X+4oh|+C$67@PmpX@eB?sOlZW^<YU1&W|f-Do(jI@,_?~n.&Fe>GSNU,:5npem=<xr>5OA^1u:Q{55s`6(,A4Ob86k?46DN	Dggffg"1a>4-m:O6x^&~(RBJ?:6
INnvWyW{M{ZUMGG
lDW9~ prkxNh@OQ4t0]{LY2]x5HZlx|cN"G`xV/kD\;k#B_i<qS])y7mo3QfFz>C3H-+.(Q21j8P}S8=7n2~^vRHn5q"z}pjKl]a++^g-(v%t0"kAWkW3MuGgMuiui4gM|vsx*|4J=^loN<fH;6">Ag3LYR	cXw@D~4~&]luWg-QWkkYl)Dx.ss-5@j)2|5	q4QEQ'**s5AuICTSD&pwc5o"lAwoesE2=*FRX-T[Cd	dwQ0	qWe1p<c9A57z?^0x!&.O&-f_6"+o?#02qQ8h;a5mV?$-|T9{t7q}5QtrA/qd37}aE6?]f.X"-!VR|zH_-oB\Lg/S}dD#DK<y5[eYv)'bYT"Bs`p>Z#IaEm);k=_^3rf^w1#AH#>*g
sK'[ *694X,X	1	w)UUd.gt$hqt9ih-P3"~-_hZ$k0mn:`n#$_%%xyp413`/ryY]g{?(oJC8D<8=RoC_"@)ONGmmfb	2U
fH!#@aK5WT/);~!EnuFkIvWU7kIJ8q2>80KSbBaC:T<zeb2.'gb?9#RSsZx9zD#fCCY}*)k&/!2h?*W +TU-bLF8*t~T7f<K:+~v*3j1cOn9mNg_\YFj"J@L(PE!;wkW]?a[VBs[<Lr}2_|/-Z^$Na ?I
'z'Vn>
262<*;(LN=&ciir,SRlW|d_%y|+RYD|w^.4~Sl>i4Kf^/94QBYC]l	A0X;UR"s7!R
N	<1tb=U_1H$:r"tMmJoSxMu{@;P7(9JsK&!m?V]F*1F&`i\HW6os@k@byb@O~VG,"V1VwjQ8y8|*F9
2s2"h+(:Ac85-k@Zq6"cZ(,#S+pUxRX~w)}=^U#lyERof(tb3H):0z+"wwxk:BY\%1=3{9/>6RLCGOp\N`3.C0N_*V5Qxo:w;	/&nx@<T&^kK9TFvDKqlkx'M%(mCr0FPF32W6J	x^j!u(4Ek/0\(0:Wv2@8n~!y4x;G^e2O1vgM,X?t_,+u5p0XS,JEMmM3S4CaQ$Nsja(7A?V1mk:m[R>
NJi%@r`^s4whPuc:?V9 >OcZd5[;Y_|;kwUq.*jT,~KQU#fgxlC	JYAZ	u|x
rK@h56-|x,?hzQ+Ocs#qtY(N#U?O?$iH7\7&EY?"X'AyV?,k*Srm22?:rHL5/gvcLh7Q"WIx:Ykg%h'v}l {@_-9A
	[~j|aK4@vV_pz;fte&~'Fp?#APM`P4mU5:1hb"tvj)S{}xWkoZ{<#YqvthavY:K'Ny+2^P7ZQ~6J0BTNs [g?=o,Z-OHU<Qs+8.L,+P~3'*]m`:IetPdijEq9PX2^LtDY.=Mufen=%OyC`,8f!g&y^`qw2	i/3Ho/DVB?FVmw=qQX"4eA"(sS{|3brU]3}<gL1@ee"#4iLE9es/_R#AD]@'j5vAki=nr?GvqNzF[;}-<Xekot:Dy9bAp6<,(>s'$0*D@G.$%9_Jh`BZ7f*k"(:b7i[GoD]
)\^daquI(5\>8<!fD`&c*Um*Vm~3'AXZ	IE4YV&Fz%Eiy{P`{b 1G=%8zk8k}+W$*<A6SF&e,U|D'{!kHHCCBg\USPp)hC[ZGH|OqiJj\1weP&f
i?x(<pgxXjF-]0l"3\Z\<rE_<%X<hu(k3:qEi*QEq\q7lDbn3G,+G3o1I"$Ukc`QD>]SBA$0.J`@N$5RF}dB<>U.K(W.25WzB$+d.VO6>G)`j903/aG@J%|c\(AlhNR+>-fP@EM!XIcPH?9@j]Q;aE*[-cn(][B0{r6|DXCuh?)wmUvQ2}}D|)YA -zx&%6=q]4!rInmMKt,Sr	$O"krON]XkH}omYj1h:9qkx3A.\6{zv
Ys<QlQc:7 )[a{Wo^Zl}HS"u%*6(ZY$m(CX5$=15`.qQC&0k|
IYY=jGBLR[ui.2t{G!yKWzC8nSqr|{i]`GcYd};E %(bEXM0-K=VV{q.dz,X6ZjNY	(ul2Z_FNT*7CWj	-{h8{.=rni&j0D3LK+~{8z;}^gq5}<-k^~It8;	DBq_/'@xU9]Cp5=[-pagbx%2).bRh q}Kp& d|N_8_S{P.5Q^CPYwQJzZb99mcE?Z5j*l3<Ii=MJAh%44EC> 1l\0&pZH7pc#/h*7/-my.Zd,40_32h[NQO\%&d_V2Hs(JRONsi|j)^.t:ROw#m.eT*'C(z8)Lu,\,Cj*Lu#53XF2O7BROKR~GG7GpTFDZMQJk7KNRL@MnB4M<vK"YakREb~x^666-aCby$G+h_N2^m_i&tMAG0
w9*zJNaOf
&\6Y1t({u]y&-J<Hc}#[XoI\(%PZ:emk.$f|,xcIE+~?q:x/p<u}LpxRcS@4=q
`>OG FT)!z:=o~rE'-)PjM\hz%0
"!{Z[hS*N!nw&_}?!1$oA1`c3K1I:i=vwSda'[XIXu#whX+][J+nU.o'&Z`=]CziEIf1*#4p\fS9f&HcrsXN	@S!3
q\8S,<je+h$Xs
J'XtfB@{LR#yv<N~m"0IiWw]L3$9/5N?Pu<E:Dm}oX>)6uJq|XV37	SlcE`#6(oUfMU!iGDi1Az %{5k62>:Sj,rv5mTQ[-W3~$jQ+
"rhbrA.-h$9!.)`!^8zrw@%Kw;\#s8^gVH6.<wd9E\Hyw"em<p?.r8Oby'Ua=iMX$bAxmK6:Hzz9'-_mS\KW_ds'y.z:W"?[mf(4VIIFR6g2AHHoTI`.ev%0q[r-/!#>$3pOIxpM[:%(~e*`s@9"u0%Qh?sar5gTK*CE:Uu r2	"7BS<P<9JV#SDI|aW:3aUx'C~36y"wqa9	&cSa^Ml&'9"R8t7e-UUO<1`.5h>(t)Uv65u+VF~]LNIT,,3knIw=!,T["IGR0Gf%z;_I8tjH<y#8HZC;n#Ki	mh6E~AmC2=hiK*>	{_S8-l*`@X_7 7>1n~>1_c/F^c1!<~$/IoMEa0v|*-nbG(NBi<`J@B`j"Jk'U<Iw~<n|/|$l5[7D3"#lr;T3[ixT\fpy>	PAMf$gHIPWBA]F"?U>%sq{]wg/YS)5}?"iEs[Q@?y-bHH}i|mnC2ur8.[deu"nUmQEQdt9v"{tRE?(Ef/=[pGd?
nzgFi:&~jh1]|'!_53G=^;!C%#%l@=\zRpA`!p2AbZs{Uy]0I&}iY#KQq\+m\}%`@~Dy+s5SEPLrT~w}Q+	A|!WMH$W+MI99D]a!}kl6}b`=fGxS6:GWg4.NG+}4AW-
CiTl=0m(}"><C4O*epa0p/,+b9C@EB<9|L{`p=5&0l/Uxwy/&!6rbNt(>Ug8F3:Y=XHjd@il}&79^2qUZBt5&p.~6PHV=OQJE,qM6@%/iYnH:W,Ji`D-BN<GLx<<5waahtQ&n<%@R:.)4eAr{7F$NVHjHpfx@eW
3G"z4rYSC'xw`y{^LXC9M?/iBP=f:v2OZ0ayt@22KzPMuKLb*>QgIXpGo>{
qF5(a^2prcZJZ	~j<9/:f
)X&h-P9[$`la3}TCjkn0C_bF`R+tK*;ov-i]TuUA"C'RED@,=kuZ[F&Y-;IthH*w=YZVQJ&c?HQ]DOA5"=ay&D4JGgD15(w=8XgNPXu+BC/NP{5sd,8%.(Y<MoY`<QyfZwDg!*7ku2tch*kl$cR@wd2sC	_.h#&@/\]g?1blD
x6')t)fN*hK}D\/-50B9hfbCSa<J/P	|W*#R4pw5~&O#>>p2(X[88.
jRbAPOU9"D>+4:JG"d0Une^%CC'RY'5^y>|=kY^1<eYN&''Hlz%of,YIF6qYB'?\#GpjSao\dQA=o0JUO&~B]3}+*u9-:nTl&Z1^f!k21#2Uq#5AO21\l}?~ckrzpZ4K>~[&|1uPzjG?p/vY[2w8:}yl4j}:T/AL&/'1T}AQ}P#yZ]6U~r0^YoU,?WH3o@W}N0okGc0PF&>2kHyilauJ&$NPkk<fiU}Bw:P=6}x[CEmFa18<Q$D\-qoRxkbidy\61F zA#4xneA\0:|]Y,1?BDc}IW0?"2V+n9Yj{j18e
5k0d+|)x}oO#`od\knb')>xu8~)[b/xMjsE{HAT/jAImMO(3NiXoQt"Yett&~X4CRRvSbW4wtbGE;"+$r<eg|\H>1rX^5jgbp:<9 _vv@o/?HA>!w7Xd^G0#~~6!@rJOD@EQ<_W]}N*S`Av/T5k'@3$,@rLRtDuYp94Zh)nf|?l6IT,xci{H82/K$2hS`l#v`qkOkFCz(S/EN`$})E\}j-XkT;8k6_E%W 5a_:0~x|3XijH{zlNKM}iE4	U<375dUPPbjFK|o7?Q0f488V-r!&!@]r.TQy?(|tp)%yG(%Q}^o{LeTSBtcNa,R<Gd/H0XLR{|,F\k(".{1e+bzPfLw)o#pE/f>?c1Q2?}+pjo'&uJO"DM6!*>[
,d3`)JLK~y'+qs`z@~*vx{p`8!dhUMZFl~lSMg?dz/4?Ycq|gqW.IK4aBz*,j#*QWi%{$%`J"Kua{	822	@ TpB)rfcv@-N:B(eR.XnH}`&h%Z?FaFGUhUaM^H/%	Om$m&p"i\b8>q1	JM5(#|-orid3caeJ3`44uIxiQXagPoaPRg$WLL6?(h(!jAD4!Yd3x4"HY!7%6?nyeT;56E!2?	{*AdO+BG]>bL".p#6Rv-z6qA(E6c"_#PB7|nkGJ='$\i16qR'L9w
J~H"4DBc3RxnZ`j^A%[ny'rt`FrJ )InndHj9u[mr6g%])L>)t+(5	=}<g`	&xdN~Kcx@{hWl[4uzDDC- 4%Tb'Yntv`dzqf
p9om8?TraeZ{]736}Byr6?hxAnoUDSkSVT0z|;]#=-wmkNM_~-[)Cq{-$by{{<dXS2xzBGBqa>|6c*I&_?>8!l 5g6h#s\ T	Pkk^>fgGSq]UO(zwg'1^+Sn4u9lOR"+tXJYBiKJdS/L7-XLmE||!G/Ct(rg9-U-x:T*>`)<)G0ZQT["F!MJB6e}"Ndn+-JCYhdJN
*p"
!JcXu\9vs:b:"K+e9{0^d]s5J`%Yc,V}K3a<vXSKU>xqN+p<$G2!QxWI?'Of?_gj}z@Mb}8q\K~5s\rFov%)U;9@0#p@?&`6B[eQvBa[)/j	62lnNibhM]jh5!P/76uh'0nkC2sPrnJj`&IwW46&2=Fs$t%^:
`7g;
XaQ^l?Pr87"Oeh{EF$yP+AhF+/2.oTII=4$~gKm+;oO\J+J6&
nVrq;7.bCLa$Tsc9]JWZ(c,>ji2dW|4E~XGEwwc>4a}DH8@>wEPWhTjw]b5A<CWc'`9j7^_,"o2#n@k]43fJ5/T~U?`*a-fK\J5,Q)5Y-\?Qq"\-[,jKSchQ%dFr&3~H !Ai4GBZwVH >#+a>
W#ZyK7d82tx;l&E.aa\	8&i~E`O{1FPNbk*mr  1FR%J<=j8>	k2E3{YXUR13RU?	0&7	%]Zcce)owb2)r51YPg)Z^l}Xc{!{?HS>#zdOGZH'>doIUo~ >vQkR	;(Dj L+]Hx_uj h!`&-#5P* nb#`hdo'}owDo}H<fhza>u+\A15vIA^DrM_~_a
t0[Q-:`h%+aq
M*eO;<RctSc=Wk9_.LX,<fX+I;7W,k[rB9tO'"07':dS9<Arbi|YW6"t02CvU/ 
mQy'%XAc w	9IF	 pVLBd9U~~gd5&2<|w+pgETQBKhvhP(h\A:L5V,I7[!qrUMY~u$OB0t:Qtq}(B'48Bhe8DpiD7 'ET)qQ.XMu]Blouq^oMoh<ExC)F*Ky$jJ}Oy`2v{<_"0HB)B;JK]gF)A6ikhQ"JQ J+J#iGpYA,nFn!DB*am,BAu-I>]U|(Q4-U)AjXi>s\E=(`5Xfd(b|<Q&%Phb/v#w_*{+M+'Uy
fs\!:{]?#B95svXDC|tx7(?YGy{P&n6(B?'?|&
u;KD8Q	TGJS7sH$z6)>>l].<`:o)q}?8,n&RdFS{4	om7\;S9C\NZ(:h-<bV[;EsaZQhf+CCM;^.Dw6w+%%|g.D$h@!BK'!MF$A!y(H
|Kx+O[#l
dA8fj!9U(]qZ]I'p/K >g,S<JrZ`zUn|uBx7B3_=?Z,uvh/pTy<YGNXZp{?QbK9Wom_%~+N2^GaP2b$YRF8`-_B>xC?]mo+gol5gN>=Oik^gf/.^H)H'v *^Fft=NX8?znanQaQ"_}{WHm${Rvv/-,xu[LXO"o&UqC'+\-6K$W;8gC,BLTTp#8tAW/.W)%P&v]`DV!.)=$p26Ggu15|danL.'B<i^$~j	,D'0!	_Tu@ D])D]XT[Iwgrjb?yIyG8sRlN}~
-Pezp=4tGU8`]$7cgbFFMLO6Z<wSS{u/aizXA~O$5^ }=K/sy)2%L?p&Bk/-fj*\4l/kHD]Kn1-DJQ{6dUd5lPmbf8}\ZH{,:HogAExpJ!Ri9,xQ:~?r*<9vVpudqW?G0_eQlGbx\ZB/Y;65gRFlvE fs4aD~`pF#oX1??Mt%|<~6yJ^Ms|M|'Oh(w-LH'Wg@{pz[^`2P.smS7S+RT:Gt%<a(ExL_6Yi|tW(xfd)ZGLn:3z_|3|Bjdkur*'/cFggVQaJN]8e`
#eKW.5S0c_7Cff).DW5058L(D:dnnNnGzL$jD:_SV
fiI&IwRP'E+8n;WH*3q\wak|Jsga7|`u0&t9O71/)E?S_,jS{rz"p]I[cS60@>qn,	B:d<kM>+/O7RPZyMKoFu._BEAken7KK03SZgTuziWTWF;~?+_mG+6GzGSOD@*m1O@#ksMY7$]eo1WbAy!!Tu#X/~Ni;J4?l+7jlIybk&(m'b`}b4\l3:5	Q+HxspuF0wVU0n4TRfG	Q(:xo^V2Y?	6vszEDBI^q_:k8,gZ<9@sC"#U*-T1Wc#?C*F4P"Jsl8~ZWvjlk21uO7^&F?8[CEsm
zii3vhtN\.piUa-4h)`p!Cq&yy*sfF]K},T} &)q)]v5kHXZi	|5<pddNLGJzdPO#iUF~f)j}P-fG,:JCor:[*RJ7h-"[XqqAc{T|]^NmK|>bST6yYexl+#5`|COpw_u/&zQ8LVaFJ6UiErc47&eUvYF(~(s&'3/LT7PzM4'+)*nU.!cPHhvXUrz=OUd
=yj_g>_e'9!lqV~mK%
'(	@O U>U0PETP@x{x 4^]S%t<]fI=Lfz	/^?hx`Og>GIlOLd<&p4#H@G^HB&Oj
,[LS>qFF
fqCUI{Euyw&*ZQi$irL"is`"qu<2XF+:ge0qSd:nXXEK:mz ^j*?~smozeq"B2(+;{A9:~LVHF,QRHKUo2@5^Z^#_!]~7#e8'9M/."\1GG[
m9K\Yq``c\@UQB[cVpveAIxD,-[x5	^`&Rbu(X9>4Ky^&%nt7-MJI$qt;6;$e[^vZ:-:aepifr(@8|=Vs7VQQh[Im@RJK_s}]J n~u0%t&fiwP:<jI2[cu'y<;#.{!P|<s.9=M/x\o5F`pq]wH^CT"4Cd,T2bi3b_w6Y8
.2?^C%KSMv=5YV"2Q[)**y<g.ZQ8c|xa+`45l;YjUI~kx65[4^ke1"fx|`6G8HC7}87s0%jMY1	xLG"Y$?7tDOgoU=;J@sI_jJ}8W%cVv++A#>"V?fw;
@jlex/&dd!^0:L{fs]NlQ4wB\LNoRCYeGFo6~zWV	.QzJ6LBq#smdtKO
7&rEu1E-SZ8q+y5tW|MUj57#ec6N28/&0<HGW. /n2e2,;UHVD`UOkpWxq_hczykn{T,1G850:mAzZ69V |}!MJ-}5V1(ZW!;%3BKF5]Bwcp]d0t9AFb9z|7m	adnMxS}.>gZih]-UKA{"TNG]77\C:ugz!L|kYxd~(;oQWqa-[[i!xt3Q@&L#3AzPq&CGKVX" l;5%9RBQo-u[FUq2l7VS-DkW(*oJirx)KZ!tDS4PJXD-3."uIPp4`8:zTKbzB&aK0kqNErtu2psUw7q	JNz9VIugiYL?]tAVp8+,w&#kw:R;QvDIk}k UF%+VCTn*	},%5A/z6|&y'U2^Spl:])1Y'RW%K'j9MfUqKk-jCQ;ljuU.9d:Ku"0i#jB^J;B;lC1fZm.[=f0:p%}v"S& R@I=[02?)sEjn.8{2I{ p{&Y<'=pg7s\5c4;6hXsYg+Eh5['AGj:ch=ND39BLsKo>'`Fu)&T=ET;@le#_@1vZeAGUriuZeF~-,R<$,oH>}^gLI@c%-A`8K-vcfA`(
&ILd$JM 9m"4	<]!Gg;gUr?tQy03yV7'5b12hUHF6<zG]9>6{\5Y%cQ}LmESvrEGB+3nIDOD);gcA6]sRFT:D] MGc<7QWJ'vh+Dtu<{ym9t)^=[iU[Ys!t+'0Z(l~P'#1n<iNusI8c4XRGzdA9;%Rlkn@Pegxr,	+MT?j$Dj*8=P3_
2;0h)NGsv-=HtLa._q0o50P =Q$a!Dd#xB].UV,RnJXQ	"hgbe^$T=Iz'<k^zkH}zx^e]T6~dxP_DT(	F;awN$1St6GzB@<VH3KNKQ
WVkY83#dk[h/!VwHTp'[cWyNL3o{J!vz
uN&KWaA/U=tnE96&'.qZFLAbM!Z_IOP"
*v9zUp>s'nvm?Uzy8XRf,wxEu2X3h
$Kw'|57x[2\x]$j_iDN$2L\K_;z&z:aP888e4MO/)F5e4d2|3kQ<?\x4,rK(C}l8X|HzF+90KH5/rE|;	7LlCvp )K^E
Fj4#bFIkq%lv/sd$y``Tp1R9#p9hMQsqaaOAjxJ7EeSmt%`8t{O9Ty^zoF58i"5czP
7\M>6[^gX03-[=g
J%n%y>Si[ mV@i_o$QZ:9+R5P_DKxC<+zBF<3DJ	9"+p9[m],9u"6E~TKn;3^TCkwilmVY)3Sw$"H|9pU*M^j_YI(!&MFro)W_J8eoaIhz(w5N<u_<Vb/D	.g*tq)e5\<(1
wb.%:0_k]8(h@$zT*U9#@\=RQscao:> xb#A"P\$rgV\:EjZ5Bs`y=Ec5=I5VZ&GUhQQn$
%x+K@Rv$u0N/gWK}7]3V-MTSCjIG%i{<&{w0!J?PYA50[zu_@A(Nf"%9vldWt~*m>A8a!QzR5Kh=YmFRcctGQY"FYqKPdh,?ApC[g.xI]O`vqj9/pX4g[gaYbIo[RUa!!bL</oo=O0d'9ndZoS(gnrA	b8+S)/h/_U}i&lH,ifR9q\hO_Kf&U:eSRtA"`4@l 3]R3|D[2@ylI:S>V&m6'sM`!%WIYx'R^\RHmKgoC 8chOR_;f*o*?zYz+VkY;TBI_.o\+;/;rR@t5744??>4&r:dVc55m=tJP[Y{EA!wG3	`;4j#5N"u@^_9qMS_KfMR$;b_oceVJEFJWWY?|F*6X('?	Nj9MCV1\Q-1k91(*u-$E-CM0=56?OPH<_,@ORjEB5JBm>;hRl)qMiQA^Br\(Os?--"O7W3&tvW`! B4w|-1a*i88=,e_zC]Q$,eiH;R7Jord%eb6BG1q$b=}XFa*O3iVORg"s_KIOm
i($`9n$
h%~bw<f6H9Rh	FB+7c9e^<Zz',)N.C,J=5Qi
X[I0OqfFuSkb$)[YXmH@'Af:]7D=e&TX}-|3IJN8Q7;|7Y-?!e)h[@tnZe4i\ngD3jYD,e>|
F{
~&b)QkDGz'v8+w&<i#,NKXUE)e1x=3$gr/
md5$yr$bXIxzlD(0|8i6EaT8xfMxu~K#|Ov_(#20/f{wXaAhTw.5`}OlepvzokT-csr<RELcj{SHD5n;E[<d@A	:N-y:>sT1e
5It"!V<}h$=kc_{V}wwS6]GiBT&LkP[hQe]8oE4nwZ8[XE?_N1
Ko(y|8R+fCsc+miTe7o1gO&vvg??YMG;,)HD?
RYg*{
[MLTg(!+vo#H(F$y-%h[nJ6ac#Qv_x9! _lb 1,5>N0Zo/rzedN1[ qF%7"*HB#=wG[jg7jNcO]1YU nAh{@(TgWH77h3MWv
zXW|\2ao$&xG@^mxRb{:EujB&yZ.c(r$lY%'7kST`aF{kgm>s%	|6+`U#C=OF4](~*OuGoK0&%zQ8-yL0T ;ua$J?Ua]Vm]^DTA`g`$ 7XdXK%BT>\^Y89inY*_/<9F]g !1$^@ZFo`TG'q?*>|b'0{R\cu0XM"8wXuk2:)\R'=?Pvdz3%<V{Q-"T%`u[2/m,y)Hf.V>QkrtsN4 `k #tHJs,{_H"bD:y6\>;t^TulS*,~c{Tm3)(!
yUW350AW@5[Y?"L&z_>`kzem;dwa,:	6'm=rn.3!'=:xc*gxoC]Y9*# `_B@\N~CnNz[8W#;w@+I1VSvyqX:~=Uif(cDtx#(\8d^yQEYalR'4nZ/`1ObtH@p#cb#hVC"A 3%j)Dv=2%dArXnCNXq1CWSsx_j56S7Z=.xJ!WFQ46R~R!h{*}43^o;<f0B1k+2jd/x*rvbE$D [p^FEid#@t:&b[ue^[78Gm*SFBl"qwGd"}ms-L&K0*ALI`l':wrsuH7JNV
.whqs(/cO/WEajV++/!SzcO_X HT	S#o7n6ejRci#u4=7`M]ms!1%>$@,mkq5w&E'Cv#?FAhGZ|?ANQxaR !>]fN#'\O$%(&NtT31F1+4_lc%mz	oqa#ndXBT_A6jNNv<5~+Gu1D h=.GP9td[1({e`lu,ca9?Sx?{=Kfk.XQsg=0(+PmZn[A3B"}fynz_n5N+jr]#rIpEs1BfkigeODy!l0Giq?NU?q"xTChL%Pokc	c9}1,s5O||{(^Dx|,k'C!NMr]H1q$'0HJx6{I4d35[hjEYEx%Pe(|:^}%'y!Yt7|v.r
9[>WR} \fFFHW"(=|(B8[cJT	Z8~Gb-^"|?$$gN'I vjI{a>1wO_roC'4UW/mR|;V2/q"3;ofx|F7S+3FN.*p^aKl46^eh@`K)eZC\Ha|#?[lgI#3:@"6as'Ffh52T.O5YGdOkWU"}Tb>_l%gNv=cN!O'hqQ<'Put>5)n9L-Z^&z8A4?74$1|P>DGk((8C|Fv7?BK]z>R L#H]Phadd4"dX+?7@4ai?0R4MjrL`HUH^tdErmfB ?=$5rS3QG:ykis{D~O3 lAPwI9Ufc#K`FO^By:N$y^yL.P=TBZ{%1{b@b4;zo<C>r!['gVHw{[k
'+cZy/GnK}RjOdEG9r'1P7huEdzh/GPA~=1	MHjL1MhpV86Ckck5Y|/0S26n!R%;g U.tzO;'?+oJmj,8vBk]:bQ.yV7#wSn}.,z[u/mRSjPpb&05\S{$j&Re{Fv,$Qf/Wy@CtW-]4L6+ZYgeGag7SSB8>rM){P@./czN-Y1H8i5cio?]E5
cnib}Z`LBWh{%7FbI&'_6xE\`o=A#d]RF_y}0wv_ES=nWyq`	16g>eWvKYvg/<M y H,p@9%,{#$S9uUARP8oVG"xL	pk$qoG<AtHepbhX|Mknz)~
OZ8SF8q_t@,5d0\sv^zZP'lj.[u#*\rI$_4!6/?e>t@X6lAX%yHqC=jeA>&
%h9u%f<
/B5P.) ^hiWtMT"c@.daQlA"P5]| SF,PA[,R'xA?N,)2>/T(o,=.&UF/.oc~c4c,c/Rc=rk{]nM@3CZ+:!'$7<!%CRoUE%dx":,^VVo6\??1vh9t1/>ICg	1zN*Cj=I2oA<e_o>g!"ly$|JGoh`R3Zi<%#jv!%/R-{	Uds_d[/RdHj)hY@DX/NJ*N&S^*iFv-m>`/
%nXN`,fFe~F!V3ZFzjzEC9Fq'$!Ykj9@mwZ]h.!X,AS%5wp#R`Ske0R%F5
qSJt(L`rci6Mv&Y^6NH]xDWy/!MnP+'(-=EzwD6]{-w#O/*3w~
R,KoNZnmcG3ae
mbQu`z3K/3{P~Lq
.,1vJHS7E;!f&'VmJkGr}24@*WVy|!cc|XlFE
Z""k&"dP`2Ld|P\nAvsir`hkr){C	1^VKd8X<v%yj3/a;/!A0z)vbt7Jvq=EH+8Aef;U\?Ez"=&#t<Kex<n{V-ih?U(2wu+r`lCvUc=|~|c4q;OQxV-dP^I3~#1uiZ6Ui{8TAK9fv{0"nmzwlMs|1[3[hZe	"7-btu0ap<Ni-,PRz}axscF3L[$=YSF@e`4,CzQ5R1$*p(GXT?9D#fq_c')#h):3<Ui6.qJsb/e+Zd<:,ixw>nLe e}_<ogb=F(LvIM&R1%[& 8,UKLLG%Aq9h=vBWJ| 9lmw?vu@Y#ks\yR8z93q*K9QI{S:egyX8ye%h/}E>=\(c.@UT@HyC+rSE,\L&{0,\=D11N=w<t/Qk<>o{]&kpeWZt]S7s=V7RoHF)Z><;))#&m'*mgs,`rSyE`Fp^!_o
H(Tr>|>g>h+8pXhh8E{!nvON:r%-7GWo`lLV7
nNuH.I8#*{:[l}J$M)shKV{Rxe|hsyz/.;{92n\wu`MC#w-}#pf~p3@]ch3BTNN6H)'c|L^`_"K$~"Tow"0o&q5^)
yX5.B'z5C7IZHvdQ(b2L
{^M#RI7IC+f_P\.,8E~0[$ocu&uOPt[FtD @3/gkz)Yi0f/B^h|a~|2u4p( i$V gX;!b3H}a4 3:'9DquLH#^V)+Va.l/CjaS^#p]GLv@:Uq-+yy9Su+>'Cvb|aS;{7v3\Sz*{+4>o83j y_(\=-F"]"J4=lv3J4AIGe;I8(l.2G~EY?9:
w=m(dETD=b":Z+-><D2uW6]4zYC6* ?=SY[!+6eQnM]~6Lig+[mu6l8+M6HP~j}nML/VBlx8i@tDN\u/we!N])ILG &]7 h;@G=!VkKFRn3fG)I@`*]5^G4rlqWA?M*vTohs}C$~>>R"-oP.ZuB6??doYgQ{
fL]PKqd Vq},ks(M72G`g0{2Yu-{Dcon$:C^.)WNo,1E'FHf,loMQ~|^/Z9!VL3-%ijx14yg43B_[$>G/o2Y<`rfI[wXzo@{.*gh~=^L\C$xyv976
x<t&;:RSQ1?:Bva@![5iKU)FfeT5G5[@;yho>\*#
hVEi(-##`lIq/TK_ERi:w7YSS+p=' ^_1=X51\)q!dx7*2svL~DbWBM?<1TJ6MoDo_U`@`5-`5HTFmQ2nGZkmkjb~MZNu0\~\*y),ivh9LyG/kfBVb<ui?%APZp41_.mc-51oe<
u:u}YC1%&<?h<y>:IJ5EN^k\$)7NCbj]F{rud&z]HIW|i`+P\%\EZeKRM,S:0.p'(ZXYt[8;z5V=svnBpxzn?8~v/hMbui}%Y;{&}-2R^BArY+SLFC1]&(HQkMOe#t6 R%Ex#9n4_W,Tr:R=E~u=/2j3Qn`8JW=+o_
4LEvf69r(M`65x'aIQP=fD)I[Yl@mEXa'v6Kk?s&%Cl<tuk%BtV.i|B8vNx=[<<UM |-/7*Q<64ubR$sN+jP.%Y%
n2avq.hM{Q0Rk]&3
GYPHr:/.Y=[#]/rbgu 	OK/@u:_lw59?~OZhy0]LD@Bw~/u}6)"\96lX@Z7QS;!{$1a%n(u6)j$3[5z5DZgn$1(kJpsOP4^{f[aFh^g-kJ[Fw(C/8rdZO4M*255`=Gj)JD?53Jc!%y&H;7{U]=Pv~KpMQ(
O=9:fP\A2Z$Jyp9E`}<[^Xd*fGmG4Vx*%it2>K{]|W6[iN/Yt(BB2[#vz.?GC?\*<E/|@$X;44Q93K7	9Q\3'6kr?3"4e=+?^0|%U?&Th9Ybqy}MINr#AJdQuwSE`Ufd#x@KvkvmBD&ei#k[l#:m1T!KlRks9;6&'
0(7_E]]b~frmNL4oL\5c~JPS_
e1"&&s$A#LDxy=MVf$}J)\f>oM3zX/d
/OYhlIGjj:T>[y9f;V	L6p1fvMv$Wwb\=.0e^lsag(Pw1y#\U}Is*q*QlSN/AW`6s\tjiQ82JM_U=[FVbOh~~-6_XaC3+U|n6drvhLWiZGZJ"'B8\R
.:1W'QV=;=kilFpv2eLKv^|q8L"AI{yl1ws+j+<Nlw(=YX!%J*[%JRIQk&W>Eb`NB#Q/FJFQ'$TO/
mmj>OHSUq.M">H!'/h6uw{wInB`QGy=2S\>3Ais|3W?H(Ht)cC\0S^[(8$kGc.veg/lBnv0vV_&pz[3Ta/qs0J=0WxGe}L^k=t4Rgugy4{Rw	|fe(F
r|0lqF1ffIKmY)f5!r1`b
/S7z=9Zv_UdU8f<XdUZHWv'GZITGaucz.C
%E3d')11zQjgxKh>45hsFwV[k38s*ga1`Y{CHs(J7W+qWELUsejP:9ISv1^94EjpVh>MD.54>NlrqY0R(Bj#kP{@]&b)%#ZBS6WfW7 oYk30}cv}@r$j|Ex3Q7^1m:bg6Sq+.V+Z[&/Vc<  0FN;Z\@PLY*_`k/b\-dIvkPdTJpgnSaeAt:Z#:KOAuF=MWS13XC&F)k4#ED/>s{PA"ezy]!*f0H":OYdQ}p7x>Zh*4QH9M, DQw4|ky}D72$u%TKN];CUZjPcsZpcLFy.3pF~pn7K=*Mdn-Yj:pC<]XQ"RjKW`R0 2?(_sv8tD}<0?G7/'	PyuW,TO=To2Nv0{@Ka>+j=,Bh9$e4E>"OvksSGZz&oD]Til{AVqZUPVFUAmZ]wn>q0%,b5*eo66HR,H<K	(jgY;B&~{q$cmO+"=/`V[Cq^f6){Dm\]c	o8fKUIfdg^e[?x^-D	 hjzuBu!,A(O>e@= ky!,<sBWNFd>6MN*O|A_<Z4()rtsco]*X,-f'\(132Pa:J-({SBm_,rMeW?x|=W* p.SGKo"sz#oL&R$=#V20Ed!vY5tzSkq6.+BX0BDV`^axtpzd:`mR-&CNy/u{r8}*9rvQ),ctum~&N7:x|{:*ZF(vX4'VzY7/&	p$xv'uD<cr^@x$;z`"0+B7r1<%X;f|OHSS(u5Ydq}kP?$0;rY9R%R.DWNpd>}NxV%*sw}Hrs0U:qJ/sHT[;-\X$MMJ>6
y,1
 |0.GRzgW'o<,"SdDS;E"/$	JVUWy;<TD/F-Acvv}M(i:ha(@PA1uMf}i"oXF?7IQVuP:JV<Af*j{Wj1M_+z8Eu!Ggfcurf+parZOgXTE`pMtoS>G@CF{t!#ej@6.sU)=-eq$3e"<pXOL6|ws7FfREK-:?W#oV|nMz Hx!4X(<rn|AXPmFm3VUxgq$Q+]H6,39MkTX
KOSxf.x(yE`6DB1rei/pF\/QZh8c)P"I@Hn3XJLa6~H.foOH[Ba8=j;s)fMV_fy9V6`W{>4[*2"qB,H-vE^[t3J(^u"?(mCE\i	=>(3kFlN[CG^.3-N``
	%hn2=Dkl)r/7|_(ykl+~nKON"%!ILrN}[Jd$$jHKl75iB(WAKTL9}]o;q+fGQB2yOr-3
l/C)*2*xr%hIlYic9bS[$0!a:D#miFF2]GhK3'9.u`WiWC83vgv4??McLwLTsj5jH?l%}j!vy'p{B6m5>
;HigkWBjY
n=RxOjC+<|#-e^v8M"8!zvO"$=J	+sII^oP}dbU4#2{[[i{^RG:+ s^,WV{*YE|n|@pq>%;WZxhy86EhfhI3eDX*U,_hHFmYe&_wxlp-TK>!EgxYJ"SPy%rwiZdc6SX^SAlD1(Ug8ZDi`F^$l5+hf7yl(1S(kdLEXI]N`z=v&oZ/az~Nf{HY(EZ'0;QK[3#)LB-qWZn6GIFF:#h&3>''2S,{w^\SSKN0x!DqYnIYjjGWFr>Emw6`7w0{X Q~0i	lM{!M\M,Yv ZRbL>!d_4#N_5O1Iz|%?]o?4{>({O:L7^&1&Bnm#C\k@.-CCLy{?#ay,x8cZD@d:vnkS"C(*/leS4VZ^XUP$Wy*`nPIbk:^oID>X~,+Du+.9NkqlI"e"4J6
D.F-,2oi}&MVH5">qY+F*^a"NJLE(K~OE#^h1l
!FUo \pYs&)LD&69{mi<fTW&a-+-:1pUyahKrM_Q_uj>5mlIzFDt9u#n"L#wvf`:BV|+wN0F,$fz4KO}9V`+E8s|'a)K6B
BmDmlJ-prnrZoe_]kCd[F3cnlR
0]4hJML,9MU+dGo,S9!vp]a,EieQY"j)/-BEA64UcBu&#bNhWt\%12ZiGo.OB.-YYBIV}mo<CT/}nc,b%kD'	 awI\a2qV8HDfWZcGPL[;hAku%ckzP4@!O^lnpS4ab+4sld6v|'b'IutLV&e4/*/:0)5#xPL+1p9 -ndRF\QDHF]lw6=FPGV<6i$WPi`!w{WJ:Dq/yH,ZqD!d5^vmz73, 2H-j.	BKZ,0d!5Qq*!,iJbJ)xW#Wk=*W%wA9k{9!C:xsO1cMJ02?0QYY
(K5;!zeI)gm%w]D"Zg;sUWif
]['RM]yJB>_&|45sRFCI7ajrY	uhwdfz/FgfA6t-45WT1qWc3UZ2l+a;@chwIiZkh,uVmqr#4z7|Hwe/06F
/7E.b5YP|}1#KU+;#)s q7>()B^VvUZO3iIs(vv Q.m

jH'R/>&mk 4(\b58pf!hh\"PF3b*k>n5LaSE'C-g&S+LB-rh91d+'CO1ySJUD9"t!Za[*Ms;xp9DnUg]^<k#T4m*'?w.h CHrhnP}Tv,FJ8jy{$Io+	os\??DRCS5
:~ag{k8K@9F-eb//RT	cPa<"r#b|[&*epr$;DOVLMi.Cd:)l%&"ATg@+?gk`6jvv4h3AHXU!T#gn$+:NpiqK+0NZ	Z\$g;y&\%>xmR'S3^7V /&pxa}3[h3c\-Gr=LLU06lPtz-Utr B=mk08JucqOt)Za(8CG<?LfNyVGk80vFWk"J)#J)zG?At@
0I"`"x]&@$}>q#*H4/S|_ez>J$jX2jazKsK+bKjg(SB COQR?jqu8T8(J+]yMF% p(|0)N&>)?	u ngQw)l"T(Rv+wY C9?M~Z{`WAn\3{:R=0^tn(UnX% RTXy?T8&N.d%-{Ux+3&]T]W[S'2?)<G/
ODA06>4Hkj7^dUG{N0*KbgSpzAB=#g|wa;?v*;EvgSw=dMKDb?M"_Pw?F]b)y[=_)c+'M']wM*#Renp,
k5JoO~<IFG}|>{Te'sP<nLS
`"t=m3~jSr1Zm!&}P KbK8?BRgjd^s'8,$x(?1E7if4!J}Z(>eBS?SSOVBwS)hh:HBA#;/^{(;b6a-b~+vP*j$TqR_Pun,,U^xwm#D<F|dI6"#nzKuH.ci_b*9Cud_o#b~;0>&=t*.pb7#09;-E7,m2fN<o)d=Z?tw80,[<;m4y6>O2hCk~`6Vi+pt3{$J*}V?7DTA	3^!LcOV*EA<}w0D!L:(c8|qCJbkTZaZien<:SJ5Vf^7n(BgA#Yf}+EuX<rgcu.%E`("NTl	Ing#A$.C^G,v`%<hYu]-REJ%~(G3hiQWdfh-d]fFVhR-GG=Y
hYYU'xo+W. yVnt=R>vW1bct]gtAB ^4\c
g}V0uvNd >UZMi?uZzA{Ao,hV_'E/Xg%0zr8Gg$1s7V\QT^r
V/Zfqi_`lY_Qw16Gf(aep5
USe_62`5?)4
:PBe4OK5hI"M{s-uQl%/LxZ SHIu(#?ptTtXB7ZBJdDK7~y{,*%st7]"ZqcNNp_TfDPQb]pG s6URG_/^A3VYh0b)OB!<JV2"64>$,7%{_B@*}[wnq!vjv9qqWQi{L[7)df6x/{RwQgo938R2e[k#/hG2C(v.~=*4+u'R=Fks@"G_.$gkD`\)jSweI;eiR(DF3%X>h?sF.3RNI]M5pI7_Xr,rdpz+4d]
eK!jm7Te2#pql!lPx'-lW#sD~4^w0gy3xf-7/nJ&=GVwf8'<|)<~PjL'mHcs~U$q06<~aCqt;z%#DM	?01Wm:?LMH9G=C6Mu(Pw9Vuwoq[4z+[o.|Ty"AUCQAC%.zDi|-{h'kio(-r"fEhMtn7u83iwd{s-7?YA|vu`7`uwmagjJ2GTN6azC$!c.\/|hfR5O#daZW=h9D1j"ZxNr3dG+:&I*9D$.^WbBDUg!<tc2W=kZc5_5Ex[+U0S*+l8N&`^fCsfS2ytZYWL.9FK&^>2Z0d{%_Bm5u]blb5i\7z>oX2;GC[)I0&_4EM}j@A\/9	$~@_=wAUz/A(G1]=?6}_#;VJ- g$msm0l*]q)c-<`RRy&:c;WR!0Sl$sEU?PmEU85&clf,n[;K?W{G*f3NEVe]=RNG\v*|$yvKb({eaMLwd)d`
SC2ayRN;BZ)9;a^0%"DCK,*o0E1tiMKmSqv1?V}uw'wzl,(S^EH"Y*Gwo_|d$"l^g=gE"YJXQ;Z?t4=SV7q3mX=iBboascO0Vxs4k=|KE[1TCZ,C5x/J1}pIK^p/"C Sm]>rmBXfGec.4Ey$XIxE>p81FJ;c$4d(<$6xU4B DZ,Jfc*=7M%]N{mS'rx8.^V|AIO+D9W2|x_5:nantR*_O\s0h%d&SNOHD1%97}QXP}*/iD&/Vuc"Q#mO]
Z'I(Sx<8K|dB.i/
$N^2;$^f
_Gw/DN+AmK4:p=Ng"sE41EYR:K^g]ytIklDH*r$}GLC3"3nv{/qLyL;wXC;g,^+ 2HI`r!/bCjT&kl&ijo;%+p`%I@rHo	*/ur!beF!srLFemqZjG$44y}-=D{C?'
+%bi-{?@/"-ZPnA	[m0M6UWlA7R=$vl swo5, 5t%sROUGC{+c]7?b.,B`#FYpUY6FdLLH^jqSsA wk2^ONZYlYXvp2W]\7[C,9]1m'RL	JA?+v~]VjJ+a<#I>%j9JRa<lnt3'R"GGw)\$>mq8q@c:[ULs+IzZ{wyO%%KJ`TdH Pt@mW`q%_@Vi4z4pB]%l65}@o-RhgB#4
#u#!Qd#]@Z)?|q%ZeP&fsJQ	=qwgj|#	'/(_\NR9Rh$7F\lC<0zOv=[G$-vilr[H]]Hu5zY7/h~X4\8	t;ak9;~?|rG0/&7%bO`3'r"],\u}?RGlgyyK]pt#I38<mXuXp:)AX'X8o;=nbg+__/0Ibx'R&@bnJ^+0S8WyWY"G[AT@bTUrZdl.k3o/)i?59L0~>=bU;om"VQ$El4o_uZQTO7+upn%$mfoik$WxQQ2~$AA!|{oxV:3l<Js_uTsAGm*_Dp_J[d6\sbVmGV[QoKi,\FOoD dP:U|DFU50X5bx)8"AoUDb|kHy2(8y2xH=M|	l:X}$k]
7ugpWk%`g^)L, Q`v+my*/ opK0"OQ/"\^6u5JcNv#q;7OUD!pW9wxU4-Cge8K!`\^(>#jE6DzI4?W(^=HI"AA*GzM<Qap2ajC~jR@Kkx
`;\p/b{DEL>O;~w;OzW$zWmS(MO/\6%VB42LMQ4LXlLEKzAafU	I)WN/cI(%j`)	*m(Q]w$ZURqgHq-y{oGucy>DUdMRPy='Cnt8]KUy3>Jl_DABnOMbw,^D\/Q$eQl=iud5Mt3#H2'[!HJBSI)U2@/"D%Vt_dx!epT,dc#kE{-*B9\]-.'TGyAEUAIx	+'!/e!)8cns\aEm8Rwh5@]+Nh,+Z/0B9ke}BlU3`	iGJk
eyw o`riD( -jyYn\0oLH1L	rQo*0&m7QIs{tD37Ks5z.#:hhgc)"tLTt,Jm<mY*@T;D::?K42!%NK:<)<>npBD9}Ao-$TBh$_'O4g-7s46O_}a_cQ?bKb9PzG;=Pyl /{!b
[b7~$C?ta5Ls:$j\ 3Z\usBxihWX^L+qp]n4HCd<A+ jO)h*g5`Y?;"hD#uUmW9@R{Lo*iNC5Q4JC$OR&|HjKP-	;2Ss[["o.LXWb3G
]?"jZ")<.B[93dWL4#rQ-aOx'Q^!=-CU'2xY v7]`c]o^;+.<%Iw=L`A6JSolh$>"o\*xR!xUCRK3xL64~<S	4,%d_QI8fDud<X,TNQ2^m5x;dR]m!g=j\oz
UGFpk	iiJ'=9-@xt`um~j\9xt#)!Oqm:zR
&6b	#qZV5PQTz-	5#:L} (WWQfi'Uwy[^Czdz(?FEJ|SrlTl@?wh1<QjWZ59qsjQO
v;T/h'9;c6/<c-+NXnr6T+0J(y20(]AZw8hDiN7 Jv]0{Xz@_d$+"sz`$[x$!-L8X#UoSQV:*xi:]ED}ZkhFhheX1VTi}s0L[cvQR()S=BG/nnyM_7yI
Ac\{?nC<_q[6pIK+?W4<<+$G&by6kFe\i;l%w{S>k~l]$.8IzI0hds*#SShUwzVvbQn^;4Vm(KU[':P6_Br;/}j1Cd@ w>K23*`tOGkC&
8ABP4y+G[{,CP!E(-6<mzOT(q8\DI$JT.&m87SWtmNs2]Q)_h,@BLD2wOFK'E*Fd
.xcYRqRUEM'F7*z8ZoOJC!0,Fh:4Vi"09iUn9;ZDEN>8mfMB[KJrqj
MMg\.[:"Q_!az-hfy+K#2'I)xX00`q,{
}Ya{a7hvY,F}l'UML|C)(W75AdR-t"?{#<98<3Wg?X [56UAy3u#
dp-%foopAVCWmZi;oOa?,5_|fT*+aLmW7SyPgu'!#NTS`YH1KbXpqzT{s"w$LZsIpBpeEO.?\-Q5C[m,b*Sn1Pyp9z)anXhk`(Tn1s1H0r-qST8eURWe7{ipqBt;+xpWd:s,(i(6g"O<A<}{	L"-'UusP0ugwEDpURo4H`s0Y>x@I8j `[u#8OtYV!:1J-*mUmyFNyM02R?7Tpp}Vr/i)-/"NS'_Umxx%P;e="Qz,5^_pT2nt=HOry1-Rx/`a*:Tq)7[v~S$`IGH%c"g{:kd8{YIeHLGa#P-)sd)GUthl,AU,8-Xce5%QFOg3g%iId;r0)*JG`8pUJI29*ak*@SxY'Zu7$-imlnLqw^,V)9S?6IBN29)#q37*hC69<r3PO]Lh1AKW,388|bH/pA2bpRLW~mr:UkP7s$w}pzk,HGqokvy/2R|viLFcUMSO\P)f~uQw2`Q&:NJQ*v<7>P)ZT9Yztd\^6(ci.Qd%LgdG~CP+3jD).yY#'*&g3uZcuMQ0T+!oNpEcSWDHo*B:FHz/!2>Cu*0JQ|9Q(r=ff'-`'JAOx?r06	n>Cci5}:NZs`4rjJw1'lw^f<_!'\P"vWyBC=`&@`Mbt|;rwB&DR;7{CB0x)ogP
mx4R;"-1OQ4QG1oT]nZk5t=LhJxGQKU`/)bJ!xC\tE7^a8z,Ktd|J1K+V`HSx}4{_)KZ!l'W/Dt{UTpJh
pb$69`Hjj:7V9ot9/*lgIT-C
h_[QSbuB,3'?7mNTZw%Xy	)|`5.K3 ]UP9kRj$.9v61/iqcH=N7m&B`YpxJU%/T12?)J4A|q':i7zualTBpgO}pRM=-Bpy`{:0)\}G%]NqimzR|}k"vL`8.uJ{EGSP8&}(^Ll	5eM9,`~}D0S'8KM."`S|V$D=yN:>9#e+#\B1+w9]&O=gfv0fp>:pBF\wI#K03^M=+ln;7hF`l @Pon?s?+2W9f*F]ec:yALC^!XZS)h#ESw6n^DL1|9bb\hP9mwJX8I[/e^Vj_JN'J6f(V8#Zk#'M>GW='NP;vrGsy[Ug\OQ2;1RmDmn=GG@D-b=Ow]In,p<5;</&+^l.KLW.b*BhvP|Hz?*;DyEQ*X7tI5_OzL](BGe\h8o3A7CUF7@
B{XtMAKbNc<_XM]W*m}q2)uVX1Ikmn^hIeJF.DGBk!.o<)*|8(+q#:7[<sdV+,qNu%j|a&g
{)WZvVY;Id,6sP;$eswEuN3E$51z+#vAF\R)W7DAUM
Uy5
hD'p8u.<2hH^~62q1Ap8]=|y+o7
snRI'q0W.u+1IUYMxFE,p>Cwm*WS*H"p+c]fr(,Ahp,73)*UTT8); +eWG3W\w+m#)pBQ6-n {b{8xhq?TYRB(	<%lt*Ftjc2lD6o4|lnk/6^wK#[E. 0Ra`cTP\q6p
bR0o+0@8$HF6E7de\(/O}-mH;o;\"b:3?7R93KLlH5\QL?Wo/b,T:J##PqE)qd\"1yRV*`p~'v]_Q:AbxO,~	*QZ=_5+YYrB-x1];_1V ];yNIe=5jF5ZaSg_@<<Y84dj"M.uyKtA<m/]qMjjE1SR6$Jc:Y8}%O?4!>}%-+%L[{F52=[3$F2>f_E(rWFt*@D=gD$2 tIux#4G {%gC--T%OjObJ!uH]?wEWu[rw|lC!`x~!&]-9KHD][p6KHC4q""o)Unh"DOA%(i<zJFoY#fuSh:wLEIF>,9
'it1r6O<+WA}L,583IuH)sR].>zr8qRg1/g<o}*(A;vVywm=lXf7n+;IWq'
{h7)m*5Uk)9"3{,.s
}5 /N'90>Ee57WW"zr'q-`mj),5ycbI5'*cnA^II`b'XvaxGA=NsdyyhG2ytiDUc<7B;F#c_5g~131ba;jB!,!V^Qh+$k<ZIx\:~3$R	24	=mdsX=GcHfFEnt
&e8-K2}K.q0!96<?fKJ6J_~j{lN2`.ssti5f+o2dOOwL%mfHMSXV8MX$;tS?Z3`F4y583`Qe=,;k34wa1i(m	flT}C+rVI@{CuYY[1;-Y>h1gGYFF thb|pOoeJIeg,@<T-
K_!8a#l8cLtPre3w'?QZ3P*G%{h
}][C5ncWdmSa	ma	qeS@"]"VE~.XJ:s1?z~pytzF#1N9O1I[}r0?oP.8mfKgxF$W)Kfn.r.	~fuo;Ji_AO&43SGZ_'k^?t^`xF"&% )S$cZ3NOa?}+>C^+FU CDh_WH)WO8D[gz
m^M
yAS}x	RBSaqcaro3pG33Y2Z>:ShuManE]#{g97u\y)/'_x>VvfB>;pR3t4%1y}n	vn-	k\!:]RyA1%LhV`5d r!&zPsKM!9jz/P6J8=-Rp=-a4,JL7QGsdJw8!mvVe'c@AMc,vfuv=4dld-lU_EPkz:%O:\vzc"3BQMNe;'?y\XQEbg+&A4`Ihmh?y4	ZgEjo-K/bUOK`vA;3`$nWmDfc1uz7<"FE;\z%9Q_L;lI(\P8c7j1B!5t!L;3!*#[O`[BbvrRCrT_T8[7	`%xR,5g=&4b> yv\PglISe>%,f)gMaX?cHD%ar6uTi
fQUU@B%BieQ
 N5Ef^Ip?FLAT;L+lY=6)awIYd.d@?5tUSAkz1y'.oE#-KMprxyp2p?zs`Ge#EZ,p[CBeD|qhGL2@Nem.7{j$]yHkTwCI`*P{y)x@,8,aCum`%o9sG=B^oiMs|lTXXx`!N2f"w-5{U(Sp'};T=Jf`zbg"_=JC0.YWfb}FR`$Iv@/7bb&:Poc1C_leQH"fXl)M^U6&u
BPI?t=@+)yqVC*/*|78]/9l&-X9NC|N+blq!jY$N[O}tVl4v	C|r!Bb3h>02?R,qw UY>aZ}%G5L"!^F%xb{8i ^q^rP*,N6$3aTIRt]G+m]l/ PG5NR^Vc@EnpufxD8yM%Sh$h:Jm&3		-V%L
Q4jKS(DA-!&'0#*'q7a[JbH(0t2r)4l6_k:(qV2YwEZ#[NI>Le=il0?3A4n8ZQH@Hnh!pSIt8pyHaD'JLpO/9mdN%pyzIh(5aP zSRAE(Wr}MWE=[WC{P3~Kj| pn8@bm"u<V+w6'Hin[(-INu2zu3/p8({(tUx.6\6JSv_ZN{[&PO<8PX&b[FE3hp6`7YKrn7Ln4F~H@yMZDW:b	Ow_3Nu'qJ\jI|/2.ewy<TeWW
m	J0'	uHqi.W07-x?01R0HJA"5S8xf4l0LGdY&0zx0=AJ9RbPrU '|n29u&X;h9"Ma:#
4Z|t_+n1Oc@J>	:lWjjd~UxsSD7{iHJbV(T3,8a{:DB%Wn&GiK#|%d/.[?v2?`\,N,G!Bmn'nJS9!9rz-	\9oMVq;7PbQ>hr8j?N}s[l$O%i[uU]6t NZ6&x(^JF|#}	Clj()/qp9i`
<~+s#CVY`A9O7MZQ=[DA'BAw&<0
7'b21`!(tuKTenOn8I~[nn9LDnjosRKzjJl&-o*_SaT[*aq:3YcM\fm.'X\v=%)vRXRpB9UBVY'~gqD$bCVM=#|Qs/G<sqg0B-z|FN s]t=|-k"i4'K;.I/RJgj]4/ E"-Ppkcj=3,[.cr`z+W@	`%2hScUcV14MUg3/)I-+JfM;Y)y,k85diE]m@rd$T`#ITkZlE#ag5\~kwUU(=1"*M'Bp=
7c{YLbfTN|b00Q^x)!J0rU*]N!e4es9IXE+>+O~<"6iUPS>b	O9@m(?M{COLE)JR>;a?Od.#|.TliH(^hjzF@Ua{GpwbA7<BSI42$pI^7Dl8PH5<LLJR&Ob_8>E;HlPQMT]T`k$bQ0i9,"tuwed$c:$Z2M1}_loyNsEn~>AAboQn{8%>&)VMnE[nVByN Q3-gNdPBw2G_u\P}?&[L+wYUgTY 6WltzHnu_Vy}G]zg^W^7XH!P_J~!2>%{5|z8TZH|%]oZQ=k\I+/'"$~A"DZR5qKKF@iGaz{P:\:HH+_bpTk
~`TA$LA5O7ij6L_Y)@q7x2XXfAt)',V>/u|8dp=Zf>2z(V1,4Y1UR1o}X;szL}%#fWuh]0@T8PH!sL$I]h[{~W'vx@4lZ|,+\,FT
@~mVI+_f+,:SvtkO6kU8k|4&bIFFa`VfgX=e,H
6'e[0p{i8j2}Bj4zXQU"7X(rRjY$ORt%wd8q'c0=F6E@m O;k='[\$D36.G +|8;LkrC1P	J&A`X)YN8|lGC0pL+iV=
h0@dL}2i/dIau#S(j_O\-<*kfTn1r1ji8gB1\{=_%Q&i$sMWpli6o}Fg66n7XL2I@2XbVI\@P3\$_Tx+ {rt
8U,k;({/zJq~#QSg)GoVA3>Hkp>6`XcAcb]K:eTv6)Z;r=ft2kZT0k, Y^,6D #4c^ufDl"	`wL1oqye}p1D>yd=PMh	zVGAT,2jYqvAjj.]*!}Fs(5f+B'C:>oGsHdz9bMZ*%d$q4JUKlaNPO[Q!r"8yDU3#?IBM85\q/y.DaKJvs+Jbrq%6N7Ef'4,4 T_Lk5A	ai?EDGo|)76M[F/H_Kd	*48ef'Y(-CW}2K+[dImjuz$<bptYA.-!6U;"cNQn>E5UQq@wZ:Db!$2J<3x*U\y=/qjklValQ9J3Z
pEqvB_IFn='Rdw\r@pSmEyLn/oZemSER8}#2%^S5VTXQ%!zWWQA jV%Vpz*xQq3T#h]xS"dCMeT	e/VF
V~v~6\GPC.EXoszb9`ukS'_R6r/..*;Vf}h1g#lZEkFT:t\z-?E]v	Orr;\Q83|CT}P3_'>jWP`XuUh&Xm}
p	>RhNobpG<#U4YGUw>&3yF,Z	@EO]@|Fz@$KB^)En0H:X)=2XqYm
B!\2s_kvFqV7uEb*.*y}5y<w%UzzxM\G5:@BhWkMIH5^gzA[l|	~P=bHS6nCk7hz"ikfyfA3`AZjbw1n_N96zkr2\S~8)^,ma_caxsM\lBVN}ZGv>.;+7tMixmS= <	N14ZZQ{h'T!9c-B-QSYY=|pn5%H@NQ7wKp^*}{4/NnPB-FR<T`tbzHOrisDs'|8uK*6~,1O3,QS[7n<O:xG|WhE-9!fFPC[kZr1\F]r&s;8?09b>6XI;|
xVnmP_=&y@nI@m%J8}B3Uqx*ogO64;!.d
TCAbwedzI<V?`n38pPRv"lS"zSMzjfYC[dpL	|ZF\>D=Y0SWVu9o$dJ&y\Ghc$HXLow}/EN>,bY?<Ux{k1%n"SmFI|R!'!8,c27s	[YIiv(hrcmv;31~<]?f2Vs[QzjN+
^L8{j*Q(BdmQg+<{]k@w<!b/%CzHe@)P[<4Kjo0XI}&}e-B4,49{5LGx-oo$Jx{~r>Tn9V.V	[!vKKbW|U,[,.k4~;H]2b5l<rGb3R.3&0yDLZ8,@GvY\[NT;_GDE8<Zk@ByKNfu2:vP&^eRA\oj1; UYE{pf(8!]a!R1r9`SqMeYjLW+II7%6RmVv^T(f&
<6*8P^K~2,^/Nw`wS+<wPc\%PLKJ8IhuA62& ]	ISX&GQ?>mKvDy/\AJ#w	kBtH^!(d(1>{1=l}GMi0`&S{I9eJ
i]l EnTtxL%Iin]W;}l.4'$?'.S"&=Zp?1^	#|G^QXgh	Wm$JEMtH/C|gWNgt+dqv{T$b2^T(pkQ:YvwmH/hE|,m;?u^Ke^o|j\wi:`[GNQj(RsN5(4=,jr 3/!W.2X&Ep.FiQO:%\MP\Q#>@Nu6ys,'$pH}nj#_R9kSgn2&\"k9MQ{u\4,m|WU
gfuNt.2/`d_9Ni
bLJuA"5gT5dE,a12V_G0Ja'rPYG0]S89YMviD /cef4=Y*P9|q{|*P&{bz-?d,{N7!=oh`H7<Pc^K1"-, m5^<w-.}dt:Lsb WTpj\!GRwn_.NK[3!jfAFR=[F3~2brs}lJKlF;X6s	aNi6IK5ka15)5a7x?!	s][<*D
)hL(2Yw\n|+g"$`[	vrWaT$#zoi6/4D
h&`<(e4ehv(w7$N+|Oj00LFH%[!cio|d@%2o%3+d-i'?bO-}lo,CY8t@@KdW}lJ)n #6r]\=E
<'{Jv>>A#fV
0e;V)zK|v [HMJT_jZ'[&VG)d6+b}O?hO#6{*vWT<$IYMt/PtNoIqk1E&~y!E?5I
(m|JZU|@PEjLSN-CzT2F")wh6'dF{Fq@,*SLB:Vf3r~Qy.dpbOzaSAjt5=Af^$oj~D4+GKO+\")BMXf4|IL>@.jI^l'8= 0)}:$:lqem6lf~'vZ90+DVQ xhERGs(sr_)Oy51FP9<)]yjxJaS!o@K2{%2TlpKWnzjc@",@C>BL>#v$V5F!]N?5-B}Z7*`HT)Rx	hqW7w^XAmW|gy(T)CwZJnaX78c)cG/[7A|r8IcXYPOp,bw-sYd`gc-UDzy@+j9x36fQD~kDeHi?4nlxZqxF"/Bv+S~)7d{s^SwXlhmcmV3k1!s{6(%(FRl6yDC2;!%.HZ{f:Ih:TpJ%VT[`?RphLkqP6^2HC7Gh7T/^J
]ZpVYg4C(BRl^+6=6BbP1Xk@W/L3utFRx&Sg,Fs^&1,1QVjj)gPIFj(/,nn_Yx$*[#8r@TZYMH3cQhjHE_-"%m@RPIzXxp.aP,#~.elipr|fmNi?(qX$m<m(\h[jO`	~y1?JjE|+n;.R3g76B}bq!\IgCw+B7rBhs>)6N$cDd4!Qi$R?K3;lLn{GLaXqY7QFGawcFI	qE)s%H>qa+9Z4m0tJ+h+EGnJv-#+m8XH[x[F[-o bxp>&%	;7[^g	@W/`*xx=MuAPA_|v'C :!rxP?lOYar3VK]Y-6KR[9C9S zj*dzjw)\Z:aM9Y)#)=D|Y4vH4;,n(&r]dt#P})`ErhG#lW?vq'"[)p3kjY~"Iz6ql nCPe@Jqei`^f%/|Zzc|.O/XrNlv\zZgxbj=p{^\u8qw{[R[W3a s^1t9>hx(67EOKB@Z`(qF95M-?#.Wd%`m`WVYJ,MWwF+H|aW*JytSqD>I-tXztIN
i==jc6!q7=N|5 LBu/aC~YK?C\*C_e37x	9p%vf_N,%pHNop=f8HFWaIA|j.PLe.7Oc_(mV__`dZ|6[W/ ZiG'>X%7L
PoscBwvAQ.JZ0:,vw-	IfRydC+):C7]%g14"rXP15r_Z8`)N<FaHy!YRx)q2L@LSHB7&iHZn	3v#HzG=d"zNnhQGDd2P8,Z)3F s5q%`Y%yTN8Rry^o	=-d`hz5|?Dp*j2v^F/[=:?|Z2ht#Zt>Obe)"2Aefq1LX%KwVS<] xH 3W+bc8G?47t;;';^cP2|jdb9k6VOt"16a'ZJ	a](tc9F5.jM2Opg"z	c#^ddeOyC/rz:r4*_"Z<.syTjKk{y
%Y3NUjEY1HAAo*opeu)(s@6DmLS&L"?rBH:&cc|GanZzG0QS6o{>b!a'K'@=wTF}qe.p'wr!UaF-<)~@\-jxD@C1]Rj'{]]P"'VH{|+{M{BgPLF5}Q/Xp^%'KM~U,o:JG9=x[^emp@tB8+hELx8<,]k`TO|<94CwsnQL,GnH"d/I4)/F1'QjS#!v*l!0v^L!$}i7:Y]2D4OW0X6q8\ES18{O>ht9]_RjA)%W	aoRqWJSC5U(-\*xw	gnJGvUz%eg'=GQgi'&!")a{:U5F\.B8\;HF|Xqm$QC1)obVDRihd)|J ssR84,rai UQxy<1/	>cT:tt0yDTXY=|[sn3|.:8*}j%*780URxCTu
lxrB6?[R]@h*=WoTVGL<Dr3[Bw5EF.?65nf"a:Bd<H@Zc6]12`^Ca>T)IucdQ>8pMymM<pXZ8\yo;i_mo.%Z4%S/wp#!jGY+{qq_KXN[JbbF^mZ-5gj2+x|Xx}?/8Z_`;q0+>MWY$QDY_Utd2 Fa{+
<g!Y<Uq%0+9bVh>6c7yBL^rr
RLw0#sTa%F1-_<C{""/5<#](_hby7tQe96ZX4]QeN-g!bdz+2j@59z0^R8MW|;:M)<sqaV#(:C!GD	aC}@zf~vYb/PVMx{[8[Gk/OEWEKrxu_avp	%D3pzPcJ r.%Br=7y0U`\FGNFMvZ7}
/GWU&7(b$9.&n.,'HDE@<SsDq-q9ubzvm~ba_U2\rY=5_lnlI;_(cB5(wRKdJ2l|s'+t$u4$q=uc93I*.lAp(~|.*FrO[#EBJ[b"CJq&w#T8!/2*M<Elzh^*T[DG2Ah	cchK)sbR-]T@@6v{RA@xf#+f*:J4"x)YkH{,8,>&#eFJ4}9IFrk13$8&%2
N^Qk)If&4<XWo&i?RLxs`f5)S!p|1m\pz0;67U06PS{fK7Lk]bq_2u
fvo<\_9hEF.[rmuUIpEe*lB4Z}>E,nq6j`t3hGN<R
w%0Bi7_KM(39(}8V!BWdRve Bk4KAAdJ><!A)wdiKD9KQSPICE+
<{uE?=
ys>?~ULW
?[N"JDT]Pi7&;ISY7*PS_}pmF`|<^?
VDKsI?8WtyXU,"YzE	n+[xDrqS"d#,~0)c}IY5 pWJK.sP%5Ei~%m]Bj6D[Oy8=J;O;x{9_6j$:p`AO`cn6*}mfK.%N%f3=Ite@m8">3tjx/(1l'F!wGJx?
.Kex0N
t<:ZDTds%0VB^hPwF|B1zbC}bD_]Cz`tB(c^k2Z&HL<'3=1|4sOGal/7Fd8nW6>,s8IC:|ScdXM4/q-jHe"q,:<N/-w|yWGSb6C~vPE'e"MPZ5-ozLkC>JC`!vT:LNi8P5aw1a0"9YNKuRT\d"]HF=NB1bFjcDZ.uVadp@;!NYUa,|(l7a+L'?}TK[t]E-cJh*Hpdm-%Cbk,bC\9LlNm4Gnzi<-^0&kMmI+_R
+|Dmb,cB8pajXEV?FdT7&EVI/qc&$XB^N-R~Df3k/Vc
1sN2C2F(#DW97f@MC,"Sr%j5AKtGu68**`:<>zCjsX7.6=Nn:*a";a	RW*(J+}*kktCivn	@6XXaQ:AW0L8a$ ,/I1r}~Mm1w4_xcorgQ)%1Ata?w>cTpMl"Ec;Y4\-qubQ=PaF
vKfE'NHNbK[4uiO<tvO1GeOs|31eI4|8S#S_A$,1kN;{Ul@iA"^OL%$34f|]fX#bQiv)Faoi=}pXuEzh2+/^6,}!k&~i#](l~/Vm2hFV(8[%eHmpG4WD=]R b&8MYY]VAK"DUb$8z	fsVIr2eASwcic<IiZznfTB{w[zu!OJR[z)aH0CA4.rAiD$g4@ql*_E}:&wkVk4	eEFlZ-RQ+3am_>Hhdt{|[gj+0x	y`d8am{CZ*	i,;TamF9V-{}:4<[j`i9t|(*?{c)19X<`pV2 O~xU;NKvLPArTOjfw#Es(:#bg:K_Kx(=,sESxj+^+A%N'.`4Lj.`|9[F$M3N
yRu=f+uQmJpI+1_RcAq++Z-1%[m"0\NaxTsQ=!WQLF?#	/RCrb<_HNLtj;K);(N;p46?`@mWdVpV>`;R#wv"ibrHR&fWnB`vXvA_mvEcb2Yvum!<o'b(^}@{LuuiK_dj.^Mk:#XZ;2%YxJaV(zG2+
}!5A^}
/[&Uo+x&]b	Q"zwbx8	PTE:CR`51A8IDzx@:+|LeVLmw{jLk(R.jduZeh@4Q
_Ll7dDCJi[D{t|Pl]33UKO_LNe
S3q903*Wi.=_JsiBTO-6RFYp5;uUB!<olcbqDUd Y!DU~T	r>S?#:n9u~fFOl)!ian+|P/CP6Bs+sKanPD\OfUwt]oqW\H?YI3<N^~N% Ng&2Du_	sL`h&|d{MNp7"r)YVje[YK!l5;L`Eb`	X,\{!V&(@7?>azS70fH*{MG=Oamf1s.3bF%izrka0`Je"F+@4S.K\H"0Z6$m?mo3Wvv:M~xJ0%B"Hm*Xd.p]e]Ey*V7Lu=H\E88eVO\Z6VfZdERDdqI*eOZagwcQ_lkm9U1\N;naLA/wm
SVG]_85yb\XE72dP
Pz{~ab@dN6WBOpXp=\fhEXM@fyR_M!}VL%w'9*JoH+ome#q:3]DehUt,1WB;m[CwH4Js2<^AZ* k2@G8+e[%(ye_#n9Z!-*zeI	zJTU3MY,;Ci\P.gM cb_q!k.7KAjIcQ@n0ejyPkMt\nKef \>E1gRBq*EM<},ow	l>LPzm>q\aVCr*%f*JY`M]o5XEyKp9JT7XS}fzwPT=Q2J)1?+dI}amyY=^k.<,!zQv;ns,~bC@<:A8AyGKoNShb/2s;|&f2~e6w>ZQ/cm"m zP&u
8a$&jqf-<Y1-|&xMBrCPf7.u0V#2!9RD*WUGsjv_dBbD$mn+1r"1\1)a_ IQ:~=&ueL1YYl'jW1~tV:TJ-bqL*1tD]Y_tf:[`@4e}r`NJ:{B-TabI~'s#aa!6Qf{{kiN9Y#cnf/?@!*aDDDrlLL%]0/!.]Ap.&0w85[VlM=S~?5]r\!uARf1& E[$8PE}j)P2[%~	g`6+='=Wi=+Z!R=H[F(*,&X`4i+1`-X9^#cT@6l~[n$3rB,dXm+KG(n,r&6]|4IQ9=DdmK&aA^l->A=!M*CqEZe1,ySR|	#gGE>dXl[GaB:GvlA)8KO[X`7[y$;'$hK ay<|9OY$;NQT{JUJ	\i0VujTK;Agjtyo+oZOJ<^J:x*T
^lVJo+ Og#+5m]z7#Tg'*aNlZ$5h<E(tOTm!"TpVc6XQ0c:
;}V	.H?:8KV?In3#/C~ER)<!q@|{Rh`{8Sq7[7tbxu 	(%2e)z9"#Ecg!	i/ EET,dGO_8 :c)mCS_H}=g3^1G9Z!&v\Al|GPuTb*ISo`[8@S"!\qq{Ny%UZ7,TFv&wMx@'P_ht<H^/J?&I+6]+z8@BN)QfCE^2flT]K('W	Y+.05c^w^ M,3/f*,78c7R^\5'.%xEU,V")Ln+yGF.zNz:xk<kL0<cSd<oR9}(gW3^|Y'n$u{HGJGlGlhrq$<p#N{q'NlgC-[zfDT)9Hm
~LBWRj8rCqKRjyU\z\GY[ws5nm^	4t)SwVXHfK`E>Lrt$:H<tH-@cs}i0K2fl<*RO`;hhb7>~m03lr;{ K39yru/"}o/|Kqh)wl\)T3\l^BQ&"~5}->Uin	vg+;?+b=c?d#k}~aRcr|wLQkn4i(fqRldb~><2/ggJ1O)^|G9ENRFy(W[bgphMHBz(@Z?<4CL;]C*>p[*}dkoUfM?'D D?Y%,rfwK~!uw}T&8UBi=Pi_{3[?	3Y}QC-t^Wj@&@vT3Eg9_h%xM:;%-jV_rw=8`Rcgd\B	PXB%-d{z<+oq9tgQ4=^;,tj-dx$Y,}?QR &
vo#CIM.)h>LS%j6cX{l;NN|Qm<$S3G3(bhR1vumhP)k6Dwf \p<iJKh*RXm0jnbyvgYCwc<mvuRjMsn;B*Q(}LF2_>l/'0.1p9@5(+U
UJTB-vxwg&cM-8KqlxGeXYK19Np&HAmH+v7N`p8 :?+;Id;|c*EqJWg)O=q#_
el%pLNJN]j}LG)ZRIv#DxN(B^3.3+gDE
H'86&W~
o('A{Qy^-VZ~-Pp-fJ(KS&bS/X(\fa6E+ /x"hB$v8M*s7'Th^Q_n@

]i@;P$u,~`%`-v"J^x`P';N=M.VEw;8K\J}&,bGzO*_Q'_zx_z&1k@4n'+#Wkbq8O&ZuK"#y:5,k)0?Q#$9#Q~a"egEI~tcVPY[nLmp!9.S| U}V <51sb)5vV/[. h2(h|a9v8?z<0|s,i]bG`$t!A
qAd(HW[;{<x_2^#utg
C5SOb61b`(Gf2QeKwnl/WseYpU^cd;-T]V8KjYgV7CSHZ+B!e\5kMSTf7
{_r7eGF,9yDOI{E`<MlT,HzE`r@/lN^?G*Cy[>nT[Ol @,d@AOtd1^8e[Z,<=gX()Ia6oD`iCoHW2KfS}:(C}Ac|X?Vc?[JcM(4"qX{aqJ"<9 
<VM9|nDe+j}=,8Mw/-3ba&d!WlJ-9)`x,X9"H0)[WN)UPYZGp=9jaU>]|	?;P5?m7P,2@WZY-WFhp:h+"4@J^a?K6H%h;P5S0;}*BmNlZ)9U;7m#<=}=}A)#=Dls{[D7m%(x|3^+'(?!51: tZAS`*0"K42#9UyLu;Q66*z
i]0h[ICKXD:5ZZ8,q10]..Z]HuKxQeyT-O.w5Qgc,R){XzPSE2(q[-@}vqM1`cT`E_TDn/oT"?G8t>^i`/@rV8lx!1vw\umf ]8=6UI)`z8_acHY
p/$0%%e&vMHx?@ vpEU5	f,3jnb}RcxV!Ixs>3W9vuq&yR&(=Sj<{jD-}WV#g\7?[~BOB2y>ffLC3itlz-'21i.ye$_3s.GhNj3gRLx.a~'y+ WgTh5Q9<nE>:Wm,[/Zz<Pi^n''KJL1hY8x3KThCjTuQ,HN	"m\krsY-ybT$^jBkQzYXk5TsYt:|yAb<U+8<FmCU;T^"2Nt]v?{x&d(D1[x=;\PQP}<azo<M,=G6-:fh!/LUo]-F
;P{Ij$4eS}6!=%{aHt~\4wkvB?5[/Q:t9\I8is^L*o,uIB39=7~d%hYgg(2WcXX{JeMl%y_^o,c`C`kP/e<QA%v`Yt]rX'^D:i{j&`RHcT|/&w`k;p='LMBA])TB$I;Dt5pl/;d9ACk+iry6$I(wN=OD*]vJ\>e,q!Rn:%7WQEx<d(wu>`)udDNn.I?"*:]P!IYdR$~tRo!+u%5vFKc6\DLlJ}h	F]Ob2!6:rFCPS{/WxO:mg{q1Gb2>TWIOJ&4XS[{J%YSn9lpYp;5hR2(	+glR|+pA-PxxR+[(~~)\\F"Mw})uK<z:B2?Z"6mmQ!G"~p?(p6V
,NEzD
=@k-tM=bpKy#]]r3k/9>-#xbY!|=Jah'`Ha{uS5^TSgE2W#6[87	gj!a~	tXg,s2nb#@JGbdflM`)	s<%lGmuOEKWR!@|CsUpVL|& a(uv8VGX
>f#fZsu09L'AYQDW!~Hu~fq*Nca~&Ts7~fle_Ka4mcF1aCX"]gl_mF;%6Cb1@g4LMMxb6,q8%K+RtNVezeua"_8,XiG|i|kt5S[O|Y7o}2VWzW:)K*:s]i$
Q2:x5Twf$0ojr
=7-4~5JMOiW9x* t,s9RH?f+Nnshs0mU!zS#dJ2}yD[@v*gJ$%^(n2A^4(""jf#5]I@R/4`yy/~huDbD`"})KQfai~7$<*aIL*~KT|5#f}fVtm/7`D 6Ab4r|Fz/`R08"{-zHbU8-@_-3n&h+7IgJ^6Ps.<vAv8RZ+BV8T+9hm]uEa	}f/`a*GWU(S7Smni~} }Cf]rMJ.z2{UZ;;kO($thw0}wJY;?E+tIa>RZZX>p\n+n|1*@&OhPN:2	yBP> ^TFiWgXns1E(*)EC6%E_}DXJoV)%0@~d|5[k*$`ugjGwva8l_m71Z]DN_b{o:TF>P=HrASu8q_VC\-W@X<*c!RGqTrN|Hdy4G[lk_~6jCrMZ,^H}%-$+M13)+x@?OATcp('on+>`Idr@[-#'ZtLXq-7%hb$P-nU\qTkKhC>`"oH? d5eQTW*0]sBxJ`4KR{cg*skQ4@,Rtfz_8z>wWE`tz*VJM`AnW
u$&5 +|IH('dlH@IJfb<E<)jT;
5>emuYhk>E5e201z=X@N$uo~0
]P]sOvf\K]{"Idd=WSco 6i5wE"OD{W$Z'cnNSA1;z%Cqa"[R
!rZKDH4q-|8_-<1fS$^x?{}J~vXW_p|o7CO1yX}7*Z>RviHO6sc_RIQq4MX`mz:P^3C8uiH;=e_d12XltukX*r~3aQ3LNnb\zmTj[>K=t]o<t*e%u^X~*ho03C^d6V=d.:!JSyh@dpNTbt|@$kAxUcG;Ny#auZD>38sPGw%NM|%P~@!b q43$~IBxu3l2aW;	%~OUc|yzz,Q="4fq 7;|{(:nb<fB,g&
|T#pW!p,YI(qxhR)X-[H)3`TXGz_tstz/2bDM\A(]%cVYUY/M?XG-W3z^b67t+E	h'^^|zzQ^D;oN$U5ThI<'-X=>aB50#B<"Qs!a]/o)r;c[yWPw@+YP>]~R'r?8;aI dd #)--r^p$k	[_/Oc^&oJ/qo_N)At xNL8
xv^fsoAUc1z4*v<nK2S#aUD"q1C.5i:^.\_k!i:8dR0.ISu#k0x_\ggV&6]kJaDu7G$49Ke}Q2:pboYZ./v^::)!$'MmyP\uh|++"F]a`AOwdFU[pozt,6aSvLX1Sfo(=&'Jf!+s'R``ZUez'R>d49>i*	"PjLJ1BIiK#AOjSKOldZ1UP]t]ktN
MKhlR$A7ld/Mtm)[C3M~Lo.%z!>CpT@4{l%7Afn*CLS!_),Ae9Q\0GMLOZ-15xm
^MgS$JJ&R}n(0g{6)FYb&?,w@qmu23%brI	*j?-h	OJ/sBm,2!7Y1cW?T1]3LJY:F*})wi[r^OU/Qc4p
|:r;sF72-45%~\;xWY=u2rKcZvafo)^R?rY>$@'+oqQLQkKM"OAC_P0{qpE6UZ[p:%oyP#a- e{ 
S*\Dx@PuLgOWKg01'_.9s=Wg1}7q2Rujlm3U(]oMr_w!s%Sj5/50s8*J>x}1 YQ` a7|/TX=(a'7j;#LyDPmKq0 W1x8:@={*W=9e[s)3Pp	sg8Hi,>L*LBzLW=;(Irk*7rZ%#gqb>1]3rx=O]N?S[qa2ub4qTEb2SJy,6c16BE[3z^@D0mD/A__ZkZ 1RQ;XHwnAE~qrLvLM-L2/lqM>6)&)2"(=:'	"[?z:|[6c(C`.`P.OXV3>_#L!Z A=W&Up$SY=C4?Du@ho1>wS
7J/?CwKwQ%b\O+cD
>:T_c1i/bcm5
"u~fGv=wVc\p{mwPT]4B?>oPET]51(s.\:,=JIA:P?f`@(U#<QFP$x3OFO/L?"nM3sU=aU8_7~g+ J"XQ4[+FhF6![!NKI&/1 Vs00u][6Tvf ]}iMCjB@; O	%GFZ\xUF}OzT#=OlSC"Bf ZI:vB~]v$u6UsFR4l(nsv57[@;![t\,Df
5:|&!P'{R: R>\$9Mdr'1bJmFa"hP<[A5B+0S2\gtjvz[,uLq	*[T4k?&r:H:V]y3fYnKu]C?;:{p#kO6&J
#svbavSL3V&<F}!^*{S3PwJ`#>$uR+fO|9a+e.Sn_U;`i=
Z9?T)nh.M$ng4G}]Clfy0yapEPf"w`4zyd@eRK	m-60R@T5~qUy_=:V.:xnR ul2k{ZvtH}6Z=~Pl:I3>VtBT;q<fw"W([&ffqIE-q&]-)+Se:Qz@lde<Jpn9O_&3mfF6E1~FWg((s
8!myB:*Sl{pap7r8R1sN9N:7RoT'VIi=&	`w@q&:=s5VWS&O%SJCq:T{Rc*KI%)FXe;id
97R"MY`{u>qgdBeb{~x8&{nZxO[*}b-SA
S)`h)<z+'Rm@]o]=ekDL`y6WcZ5V;K+b/.p]+NbT2SuWzrP+b9HsxFw^w%3#6kBXB6},/&Ji'_)O|co FNJy5[DZ_[3."(;V}+I04>AYFAq|pVy:r$4rA3`KALk]29_Tv|)?J|zT3P~Zs&Oq_dVQEj%NB$n5U9rj:$=zC}j|~[8U9K9q|Ph{J$?`T:S!vSq:E|u}WBk_G"kaQSeUdU@4jz;0nr_zE'%d!&TllmHE~XGP5&]w"Lo	bH|@	R(p5ABf	;sY)>>+
:l[^-9a_3?20ih4'Y~>Oc"/O
}1$d>YNZVKGlptqt'ZWvB'Ay24V5v6Y6L()wy<d{m8HW@tY)&o}~6]O>`XnXs!^~t\txgro.KUI3_\b_y~b4?_@&4#i*'nOPs'U>YwJ~}}Jdm)IM\wxO*h[^nEXuc5+Jll}:9Wvb?5[Vwu^	~:d'+E"HdGwYsKaq1CDE$(1O3'{&|^Hs4"$,=;"/_+U,w}eGL.2jc/qY15-$E99P|	{$~|qk(N,1Zs"g
/bW-Hd#|OyVHCckw[pAS}8t9OZ<gzmqn+^czAM+U0`	tMORa`F'X4K68l&y+f[WldO,J5Mr$=[[l&9r<IVVA=9"
%3LyJ=&T]B!k0QGixdM>y82l2;]Y:om^<3T>|pOiEyD"k;Yh'w<{NO$o*+{Gw+u	kC)R|]~-k _Jr[x'9m%Cm(?:7d2Uud*2_YKC]9gh; {D4x0.Wmsl5}!kD\^p\a\D3fXra@dT>o5d*4Pz|B"(RmN?\/<,j9Ft=p>W{!]9nsH@iRahMoW&J@n?m+gC=LS##EhT9Z8[,=LWS>hX'^]8]Z-kF7sV\fh}
Tkyp8Pkz0T9O_ :aH(&gN1N8/^{u~nN$YS\zjERF74`~;fI;&v:MyDD8| pvax\IBo1nG5e&gB/B8J4%s;%2Pk:jd5iVcwa#%l$}6(7/*G_S{\L,mA`oNH"o=Vfn;;+]!|^i%-6k6b^
P?6"B4&=})5n
\s~-hxw7b`mwDG~@^AM%&ZaSV^,j(zi%+Ih'
GMO0\qs>"Qv2P4_yJoTrY"\U1WN{8!
)3Wn2
Mnb#7(L?6QD>jS5P _%$7q[s%`/%ZMx;-Rxy>mO[PV#~9DeP_$Z#WQD9Hs%fNl5c|Iku[zxgW,9J#L{ ,g8ymP]@m$sI{Cz#+.7_<OSTb!dX>M'nKE$zK>qN[PDdwH ^Obthg/uCCz:bXF0M_H|CbIa=,(ilmLis`Ehd	K0:$5KgA|g7Hn0^gH {]V]T+xc
avYc!}k(c(eaZL@fm/!)9wYg3kn}m!bH9kVEftm=lJ`B&`O+O`SFYlm{GXw!}~{O3}4	y+RDYIFDCAPhJXOc273Dnze$EB$pKmnB/78,&x=(t+Y1}YBZV2,;Z||M{='ffLrYQ-RH DbA5|g\aAnP@_8q'%Po"v[WQ{!y\{|Y$xSqC?Ez9?{UTlms&Dv!ON&y7V=TH,A	f@VuI-Hm5}/m_4~=v16nTYYAnt&s3D7F?NYG"
Bg>%QYCNbX{+SXLrAXvD"g6g??A26q@S>jlrzsDx_y";ib^tZb0EH`*/Q3;o>3<3U86%i]S7?$.}$HzR)vLm^tld-QJ~TOm<zh4dY'E)N$5P@xs@9FLZXz-?o$LO8}(00S}Sznm8AQ8AyFOr<COTL&*z,'j@nvwe]T$D\l}L)U<r(71fuS(Tw.d"V0,rBn#>PZlGK9\5od)3I',:28xdmNLb	d0YJ@IOx.)dtE8{WJP10~d.go5y8kBuWK^R^!l,cgt"mkPQxx!.v*J6p/Ja.6f?[}qXK}T]YJ94xIu2+?v|"/tjWEJi6{$63%"LV=gK	lCHB=-3qnk!*Em|+/x>%|1"{z~?'`q	2]?1r-Ai>EY=Ww12IVe-$!j{s5fa~?t:7~vybd5x$|9gcduL{sXwfdo?'&$YYR~c.Fl=imkR+eavehqk.":Pk%y?Pw!>Q<@gWM[)7>9/a;1BQ7	vFh%RL?WuRtwMj^b46WO5a+9CjxEO4d(;^2l@GbrR-'vw)EO'B_$hi$yZue++;>/+LWP;X\x\expLe(m,2Wt^hqOw1QM&PdT|5-nZi`ETbE{%>`Xi4 A43)@WiO~~eYdkvjg'/S5)g}"FUZu~zO
aL|sSK }B>3Q2+,O$45Md11	E^k5e
	/Cq$hISnO]["fkJ{/Vf+)#ZQ{|KcQeT-:,?jp<bZpKjG}_H+yq<Vj/vcBg^okI)@"n7XtZK'LtN_\*+,yavIWu(*fFp^`v\dq<h|~pCL6s$2AWwj&-xZ99i6QYi%
<{cF3x9vj#Zh-]Ou_;O!grj,>iZM3Fu(=m3y?9VPs-
)KG^;7eCd}hFe,\vQOTAc;Ra$`^&"~0&smq)%F-LEtj a1^'^Ehm}{QWPs_gwm/S[(t{L(Tb?jA/*%]nsd|hh8M\8`!	Kbb"{c%T9"5cYo[M|T{$bh}4x^@a{	E2-r$cJ[&SB5abP+CG(aCYI\('-0(~g^.^OrP\UlVqp*>j|U'.T_z'9`.B7a$-X~O}MWO*Jn2YyU;Rdqve_*yZBRZMrV,[;h$Y\T#J]j(ODo`WF/-jp?fL1*`_n.lx;vi?[#S[q4nDczsuuRYP#']_,	j#'<twLmnwf3|m]T==S2Y~p;1Q@1}1NW;o
%%H]5;Z.-2Zmg9RmFqzL#Va1{K?'U,p9_Ev9gn^IMR$9+Mx}]~k3:;o5\2q^aFEXu/xIMpXV5c|Ku+AZ&qK,|K={+
~EcPpWfDF,~0@yN!?Mk^6mj"`	\?60rJyD6<6pRxeW<w-+qap%t-*RMnc@hQ&\k%f4hS&S^0W_U`BEgWk%.)yp)bQz'ZfQJEX+\!v)mR7z#	Wg^+4l137<Gu8HXW)':"YXK!:
/NtK-y(RKMiR'Hz; -@ERN*AkK"|X~h)42OF[+
^uC}nJFo}q#26d,Ge8w(d_)#Kq:lbFb_Icskm2VzCcU-n9^jYc5fUWq-#G4@v-E81%[Ni'wiJ7tftl~n;'Za0DYA&V1~}@!~{.4MG:4l+3$rSclgA=HAt}ikH&loLcOtHendGH|%NcxU%RLG#,:QhNm]j?ip#`!aK${)xKCrBH&<'LhK_h?G"WW%NC>xjZ=eJTsEj&4#K%mk_PU&y M-oR-.kPw ;^nst={m"}b:HT-Mdty%;*?#fnKHZ0q+wiOG^.A0q}sZEajFQ$lgo+|zto(80D.59	`C__]gKy#"'6\zJ)h,*_nz7(Nt/Tj_2dI/R!]\,c)cqQ%3B2R{[i<L$R;D_:A=f7:^% Zaw9s1b<|ld@,~|lv,~)_{o@s@T6cv,pMo,a&;/ih/rR4]p +F8QPB$^NsTAXR^0pB,PVj]Pm<5/1t&0GhRvT|aIfU+%>soc'#}:7`Q&d|gm|
}m6%b=]pbx|w$K<x*+og-s
Z0s(T0~"	p8|%_Q}3V&'Zj?FYd3Anvp%cCE{N9X=k!Q<x_vMr"_],>1BaS1clg4X`l+1hA:|!*adCk~jQxOrO%(tlxD7cAeVq?Ql=n7m`G)VQMe"15v(|{BZBtkHM	uZ,.KE#(hRd5>'tI%k7PV9g-j>nN<k)k-28vf;gq~4s7CD	LJ\.3kIdSS$j1%DP[)Z'C4]j~!gxS;:)d{u-
S,jR"/.@{MN:Gc'?Y0.MCTtqAgRtj8N>XZz'pQj,E51x,]|xw@.V{5@Ij]=v'\VJUP{b}7kg]!|9 1XEI4}KFp*^Pb8*B)~zxCZ,t3b5g:cm4DCSJUT[^fNW?VnI'R+6,<#usjf>S(@[N4S~n/`9a>bpSEqg	'&~o'1rp$jzh?0yA<&:V.}V.i5*SttsSk@B+v$.,b4@Z?'{xQ,^G66/n1F#H0:<&6WZ4_'s Dp_fvQB0VNEtc$co; v[KL8}e{-)K^9J~~8FAnK,gnN^?)bLk_EI"72urI_;+T2 hCu{V&tum$|uruQ@gnm#PZ*@U#Y{E?umoG@Y#IYk+q/XF(-20'3KztDL8R:}|S/Jwd4`U-;HR]bpdn}jtWQfhUqN,:}%@Cm8i)"'V'D+?O^.0+}m8^wJAi!$9$?S+Ic5U)\?Rsvstu 3J@vt{VV`	!{_h'k>_%,+/_A$D@]	iD<U2$cSqW6vJA/1xE~JVf{c?bYnrH	#F}h,}6sM1U7,.6j]w5]qh@qIX+D8ruN5PJtF2YgA""x8Y3%&S>rsN{ghC<B4xUO9 >(Bt,3yab,USlE|3BA_cYq)XC'-(u\$PPlD2[3GoS-c6dyf<<c%9eY5QJr^GZTBwk_VezxOR+BlkZP<`=AgEG^&F<X<TuXQ~Pn!I:1k+u3%5 Li>0'3~.7dv^]\K)\1E-~Rn[xm1~nvnkPL9BEw<IZ#^T}a}$8e*dD(*P{*@w*BC+@{zKh9>/.<;e}q)m!w^h^v>VKbH)H5#[0R24EFzGrd8I
NxIQp2;{q`=aX(B6u7qmJbdj%gH"tMT(8w?k]\K+;ITRyXL$,&j&`fQ:2Pb+3-6R<Z2/mtTglKp^d2<GoDWBT7pUB;t1bCu}&:Xd;HVsrkiddEYs.(Dsk@8lP]J82J#|^.oInOM_]/BTZD;s	_5N0WY#hhE7p{Cu"QJq`LB98eF|JaKW\x]_<jO)~7 Z?aH:/a'i:^q?S,2FQ+{>D,v#x<,`=rnNy1o1[&OQ&$T"{S/o>u 41f>XF&gKH0J/uqW&_[H9)gia09o4\-<O9'9v,jY3[^y&pz^/^<0}TjgG:f'o<@j1'SKdEn^TYos}>y#Ct({CB@@W]a6vHO4vLY.tF:g6m;-P\|+v[Q~MRdCvR8:>darX7CVzp!5K_}XjfM~Rysml{3&n7C6$^`G;+9$4?gqL$&<;0<R&6"ZO'U_T*S>SCbqDn|+`|aEL<v"V	4"y8\BL4n":X;^BGSRE_&B^-U+fMF!v|h1<c,:*&{>~T1b5#s{PFi$p[-Jh__eNZi})[(b$@VAQAat|]QF%(J*(T5Awjy$ ul	`val8
	k#xPC2Ww	^E?7d <6YN{Y?		5Hu'zfy-%fB0's%)J=jyhC,[Pb5DtnN?|aV
>38;N2"eM(!.'BF$aPy$9^n>^V.=K{j&TSjm	^w!IHIT*U\_eeY3a$iap0	Q+vnGw-+Z$FDort&oGlA,m,msDj	FP2j	$1a`L!BX(W|]-is_yw(:}PbR?61!;'A%	90G(tLy}4&)L/!-ZBeNyh'74U+sF_S(&3Zn&LJsAU>5f\ocq9zk0??&0..Nj^b_0/17nc.e?Cb4y07PK7\?G;:ESdlZ>$.4`Ji]LY*E2CI1
ySu	,f4h5^<Us5Nv_Xg7ZVe%BJuK=Lf.?E#O3pkZS,arjieQ &J8%Ekj8fYR2h%a;X,2td8vB5Ml-{*J6SY,/iQP!W.EY
B5~%ZQgaUVKx`m' }>l td7Y}vs3#P[ho$hb
E/xh>1a|#rcL?V&7]>&Cj;e(@[Ua]&n7Aw],y,*Cjf(VVD<1LH]CohOM!~]a*'Xf,ByUY,>|5?|/p"eJLA~0&|,ze9p)Jx/mYmkea61+0]Tpk!9RbOe	a|\LUdi`573ULaP/ca-4n-g*Q<QUNcIF8!zC~nF3sx(@^VZ Ik`t'7S^<`n;^Pi?z6a=6SD&C%,F[x4.oBt"j8[Z-2W,pz6]}XR$^JaPE.U)$Fs/j,L
pE	@g@=>OBjr'I^>";'uQ#V^}Hn</M\1lbm|P
$2Ks;TY*Oh}#l^Rvz'Jr=Z@g!84S\EP+[7kb={we9.c`6XJ'P3y^;}
;f+2FSm3ij?,O]Ve4ED#glod~
0SQ3_)__IE ]y>u%NnoRf+b$EF8x|{gr[
44"i&F.g9(3)G}i
toosV0SJ^}4e\$<IK5N)]1X*2"_B,B3#Zl`iud)=&PJ+x3aiD!M'u8kac0ToMMX0q2N=~ieFJW5Xp*!kOV?VFBI`!=49\[r	ZODVxP6ijj_I19Oo8kH1lEnS?J.kVj@DPHH&I7X3K&VUoGruJ|rB+}'F6{@<rI,?i,4$':R^e
(6u9u<zY3aD
 E-hJ|M|c-C,iSik/tKs5t'S%
AYd:;?x@Lb7CJB<_><_Xjn}-|(5}Y5=V2O~G|#`QQw@yfYn#J?k:6'7<I=w"w}'lqtmi&vuU@5;t>C*<Ml&2u`Y<Q%r%h"aeX=#$kR%G06@+^!|f=_y-
EBu!+oif]S#HR$T/B-+j#TW0t~Q+S*PF.m=+,y!;VqlhSdDw$bO^'-PJ%9TVW)d!zz!TgkL~tu~k]tOK!C1|PR|M3G0Ci^,x$@$;k`Wf Ml(C~O\C)3sX`#N;,AZ3zrOt3~R>mNizZR^NhYB>zY^(pOddEi(GahEQ|$	Wd=tYSnfA,\A2; TRN;CA2)n	Qy7+B!,8VwT#>bb8{gU&Eaao(G(='A'U01
$f}|c\
8(XESGtvINf?+fX\pI	Fd}SLJG7ZjvIlw
y:Ig_(:X D+o>#|qV!M87).	/S}mic{P)oZfEJ2uW6]*dj}*wM`fR]kIFQAjCym"9Yn~\=:`:n4H`a"3'|H-\pVBltQYH!\@yBXX0wV?@|\!( (Z=fC4%,}=	['8jphjg-z4HA(1x\g;459IvcQ+pR1u(B\2STq8Vc:J4%w=.8[nn!qpmJL(42H~d?gRl^&$Kx7]Q@=`fZbuPDPE,G]Ac,AxToUL$6OkT"O'_k/xw]d#}Iei~RK
zQ1j&dItau[XyiK_aR9|a({^|a_!US%O6Tx	*;%f8-K-pGKhpOz<H8.dkqLe
!@><jPwSYiO7e&s@2nzJ6+&32rnmlevt!g,+q bD<XIc0=,-&iwrilFzPv]am)DGkEtmPJW{+:k:}&8q0/~@@aJ(zA#>EGxy/[EF@.RvH{1dNsH*HVJpEF<@=4"M5Jm^VKt%CI{&f8[yPw#ub\6t34"1WEwHbwkIwv")(Zmss{Cf6:qJ3!"s44WtDIPbH5PR.RI%	H\wbi
_s ic}pYxG^V^{` xT2tvIjx/IBzp+1l/IFrn6z
3L(5.>Bkk6AcG|5|'[L/s+@1XG%;K)EON2#In46xHz"YmdSDl+\=nLas.TP7.0"r4&vleYFjA	u,??e&JqjJ3xX|HUe;YGacV~ow&]4sg	%xR5"sxl--Hap"221`u:U-L'J0ytA::VoR"-GPakgpOi8[Y6IN:aP%|(/)	tsG=2x[MPpKw(wZE	eZy]hdu/>,;(,MP_*}\UI81~!R(:pR{l.@Y.6$_f\~"IHE4AMX=]-]&`Rxogzs#@^A6oayx2)v$A<7_xbnORWxi+#w<x%j?$H_:<W"Uc/c2_v/h\:4J|~Cv}Zhxb0TH2BQ6hH{SP[<)E
qjW= 
2@' _-J7W5fk0omc|d*j4c~O/S[_&cd:$^y(uiX(YE,o	3(aB*xD<RWS[B4FN"BYrP)'MiWbAY	M_BH*D}^G *ymkO89l$eKuY;[mL$	OVW!]2/._XZEhnN"lKa<i8lgq#vr<s/k>.vZim?1UxHai)]@I`:=Y1UVk%%rg_L9l3mj|&<K0c>l&A>@M]cP3buc'lM}QPj"uM6k$q>AMX'r1;L&$nM"gP3scfr!/wl+WMLNP8QK:FC?DlmNLm\jDEFjY(IZhx2	9wx|2^ 0g^zQ+nOG`
NaV\mjg!{S_Jd7AY+eo\{RR?a0fEXZi,h"NCsLfE-~D=CEfZ$-)+kjW3q\-?!
#z|v7M&mmrh
qM}$t>_4S[8`AsWm\1^WH<[N]{{-$
T;=B~f=U0irO lQ<&o,Ma`V~<d%<z+]'}
(f4/GgvJ8&`o'u+Slp(gHxri`^fY+:H<o$|]V%Y^$'o8!{@*#5Ll&
 	Qo1TY+ B3-bv/^2@q`qP[3E~n|aZ<#.Z7MsG(hGj"c8!^r$[6BY0(2%[TwjaBj~1F4)a77]H%>N|ZD:(\2OOz
m~#!*<^0k{-(=.B M%(UnJ3QF!sr9t"6lmiNH01^hQ%P [CZt5n"kbTWlNeIL'2+dm;4dJwJ,0]ad;Ts`O:/7"EX)"J>R-CTK)QM~_=B;-tYCbzZ"~1nx}NsUvj6I)Rd4$S#To~=@s|zwxxC=gy:WL(5>,~>WrD%U7<mYF-5*p1V-=0\'5glNRZ2WU_cp)Pi5?gs'}:Z93pEzh{gv)uQ.=G!LV4\@DeU|X-I:Q;G A+`#.2$8oE{sM>]Warpgkl< t d:l"UC,y Kp2h33^KaWZO0Qx]a`/+=Ap]hBx4815~\^slUo2o&gaU}CBE]Xr0p;>Sa582f-WE&;`yVkFWq~|!kp_@:V6c7GI='SW)'L~Sj^'bEe4aO3k?o9wjV9	kV7p46R*bW{v{^Vy@#y'nu]l
mq<z>u)?2b'H):QSS\u^-n{cjRpYEK6|'v~!N)&1}@9R2XQ#FDh%1w~Mt
Bz1rP(2]/[O4M[`,w@yP"C+E?%E*dWn70dZDfjDO5T~c]o1_L*mWO^L)voJ_K7]oQp`8A&{cW5mSr#[xRKMS&cu(1.n)	sd?e
=CaQj()-OvG;&Wmpg8V>apE>D'AU	/	Mozi*.*&#e5GwnnI,t]MnK ZPdw"tD)$^Fo>8H
lUY3r 33`9DbVo!vlC6'<zDdHj:Q#2;v=|m}fc/k#R]4I?[D%,WeA'==VfG{w@c.3bYI'w?'YM7
gv$qqz!JorC.c*H}$Wr}oOFlE;i#anA`GF~{z|!*Hes*C	}&>)x&;hKkoPyA92y
`E`yDA&6~U
:N@
LJ"	i Yd(>aQk$Ro|J-tN?}:nPX@dYJWgggDq.\4y"v-.m8kQmy\l'%FN{2*[	S	f2%tu6T}ku5K)"+db}}=G3{Z~{.Q%7~,QX\ZX~?Y^P;}ahs0Ak8)EvlH&%{.qiRxG'qq:A{T%bLh5_\Lo8i@+DGMN0nuVy2OyhJg9qt*vC$3Rt-pODdrZiJo$gHKm@GfC'XBN#ma8c::@D,mo>0MvQpz7{	 Yr{Mf8[:J;mP!a89}Q|9M`MK]336H0_L}|/#Ywflb<(98*fX9*?_;|fy4/zB-#CW$[[8oP
H59L]|TS&6B:l\6ZNvcp*nba2DZZ~v}29	q?^;XRK1BQ ;G:56"ZK9COg`=Et|4W?P5Fm5p5f-%NyGF E^c2S'DlO*U#g}*
!0l(57c#Sq9p.!w'=G{~n+-m6{?DD2$va|;v9 D		(Oe&4$8^<k{nW-z*7GQO"pw/OVs5@{|du?qOE27fJ\:1[IfoLiM#dn[3S*ZrJQ0yZ6fd	Tf:C.yRZFr@{Z?ht` bhb4<G~nKp/fd0@/po<zPcfryCi)6Jl]RO^&xLhzhDy`"ykR+HiWOBN$NS%qt6\]?e=<oo.y-jcTI
y(3PVO%_"5D8tHn4-t&GFQAR~T$hOjHC
}#}O8[(t@Nhg#o%Jlo4Cw:,1]i{hRBp6?h\}OR]`],n[V&'@M3Ky=h+&IqVI*LKdWPrhgpB#Qzn:^?~0[j|,SQt%K'Ij3tNj4vatmf|Q*<]&i_B=)Z>t;>|r	T&%qNH{b<i@Ic2/_XDzNyu'/~l| HrF=
HV@u 	@B7mNUm,	mdg/LFK*N]Q't`AL6J*YjWlrD;i+^Q~&t=/=yE(2NGv&i(iAy13s:$zO!Y!{QPSL[Q@ixGq}Sj]'hOVpw^
.fN/ERPR619ZD$zTt!HP}ob2Y[o<CjCce`}1c`L5'}],N%aJVb!BS<L{o+Cu6CX_Fpg.qe%?=`Pzzq8
b})w~wy~>$>O> [u~C8)7&:<!A'}*B$hc80,+,-&`yBEdu}BV~Ut7AQsDYbsMO$mHD5\pp)kg44={Wv;t)hS>?.{4`n#\Y(|,R,)]v-d[X%}?:U)RLyln?*8!r{
_H^!mD/X3S$A2;6$\tl,}MlI!#5c)sPQ
+|JN$$25vQ9<e);kZZTc%qD1n\Up6nM/w%aJFr"7~'TF>wCDQNqCTMN)#n;P6zCUM	k$T\\N,0B-g@DW)I1GkA2>`{T$/=3n7^f%h#/D~NZi$,Fb]m	LD=0-vehq9n*Aw
A?P="lNd>=`'Fo~|s8Iq}A	(lEO@h[DvOw;G',i,0H=){
4wZ,{hxa@SwGfMU;&sQWM,n/gEb$E?l}y
vRJv>Y4@*p^D,Yr4x}%0b`n0P3?ch4)'5@2\vuYiRz>|a 7n6<c-e-	kP454-$?$_%)3ZQ&AH^@&uC9J[hY4cER&I+lie]jiC}6\)Yw@N=g!L0On.'wjcd":PSsKyP.)?or8~a,}hh@iYG2ikcD(%X][|uk{p=o*X1o-pRZ`zyKN477KO815{H%#S@2*]LT ISf)j9"UopA\[tb?WB72nKo]jVvQ5/	HtgH~/o{d	84^-7U?8D=Zf/7vC43LfCm9~`O8a}Xa0 /{@x_UZ(NPLor6ry2ZFc8UK@^|pfR)vt2<#&80jwl.yB'Wjr<hHsMO$1gHvXj6vY_G)~/g7Nm,*Ub.s+FrhU='mpKq-J>F~LRpZkw.D?,`Fue$&mLC-Z-r}tS;iOT{W	)5GTQ]Tn`&%vP8gZR1SOsHiJY73ABEW*<\v!"3SiwB>0+NOnx6FHc-m2iEg+U;\&c8Z>iL2-)?rIZ>}& #DH$yG,U)Q^3}Dcn;&Q>*|iY[SHB,Y	]=WYDe}KeeVpph)Nz%?[zu7"B;7<!EWYBY1*w[&:*
3	TVS,:Udz>-}hBZ[	T]qzi:qwnMu7{&utZm]X4P]"c&Hy7Nbd_7OyEQU3vgw=F;pWW:vYAywh,z!ns2LX<5{!1l'/AM"Zm?8~kh0l% mxfRB]+gE/E#H}BBJsiRa:.,y'X:\e&B-dNntq@q\*,VN=Ws{/;C=!p({PW2g~3ke$]Cf^>zB?eRf~5O7(WrJeeU{6yQU]0jq!;4}'|AaRHkjzCQTpfX,O+5Xv-JH."P>A1=\a;}w"sg[86NK%)/-!I'HO!SIb(F-N%DueZ21@-T?tq.GrnL"mPAH.g;#:!J\rHpdZ7/Fg?J@+)hh}.ze1uinSbH3GotOpR9db({34j5r<ll.AlLeD\\ 3;twgq,qR(svf~UEHC(Mj
bqFA'h@3}@P3}oCp-r: 9!c}iU`\^;>LQ[$5&tD.*VI2l?5=?s4y*Io)|	F|h-E[d*k1JP%)%#fF%r|@<IMnvK8cPN4 I ~K2TH:oB_v$wW[7XNJXXFV%@+uKWL,D$*9+n8}\SK~'	
)=/Y>o 4b%@{I%^z?\:MUU6F(Xe\R
{p-6oMmiqIMB
,+jYrv@Qu1ZS5"%V2%kM\zgrca	2h <:=c#f=)[mpur>.Z$$89vQhW4U*]**WJUS%<Hz7Py11u.$BE@l:jE^@In6.>91g2H5-:`$WL6:bj3fV)e:+U4O,Zw3.OWNcRTxVt(2gEl+euoA`n%Kn<fDy?o5).oLb;kPl\[oGl:[Tk

@_i'\Gce=&zR`bJ1IZn%DleD,V>buMg+7ibNSp9&$4Q#BB"&dlNs$f2Dp=}~vk(=
0;Q[."IP#KK$8LL!hc?=>X\&:=2E$$gRk[GOAneA-(A]Shb_kwU'ZL\u-OP:H7|5dU09B7WEuZ{a4o_y-a/5;ikstr+_n~)6[5$m?&Ks@\,";^0xIxmMl^'Ok~Pf=C?j^l&D+|y_Y#%sOSt8cLj#&a]>fSeU+UrW3BpWZ?"cjt2p3&W_RM|zs"qE7[;~whA'cU$=wnjek]:n7F@9)5ze-DY.cMf6&r1ls8	H'\d5WNtP"uv2-U?Np/	W2a5"_DMlWCQ6n`*QjT*O!BC/MNI0QL<t->kFI#:twxt}F1jY}af$tV`Wn<);yW[|Bg'tE|Y?FW2+'snfTudXdrdOm%yjzyT@kkp5Fd/ P*En?H)r<5S8xS:<|| V-s:|Q_$e-n(%KM3nS^}M+^[=/>,DIySQFe;1H
^4RMjXJ0_w7%/zr-t|ZB%qqMp$xF)"kSvt)bpUq'92"9x]y>dExaW':!/L#)v2`KB_w_?j]Z(J^Mw4oDSvmB*"l1cm\T*&ic#g)914[2w-#P&'{657fP-^\NZi\"=rEe_JE6?=jQK!_{7enN	G}Pr!^"0BGx:Eb@5^I/XkniwyD~q,8C7H`
G
*itQ|!q5HZ7,??,r}<nYc@	'81q+wnd.vg:AD.k0,7c5|aeIa@Jx{3K>c!l
y=sucz7Fj"*`HZLb[D'FU6@q)[RSkqt?$E_Wk#
puiGz6 Ifcwe&TA)Qi>c/
W!-lL+.f=G^ah3.V]g$rhB%c+04$G^orrrc{iaHOX+5Qa_)&D_@ HHq9ZPtAs5aW_F^46&x^e]jk(bja\0@V{\W>yD6vG<@3+AEtOIZ%c9]>GJs]()/`a2h/Ul3IMCQTH(~)?:qx{V^nAr|:&Mxxq*v\L"J)cx)l-
Ha
.lyBR.8:oGJcjst[9,09WpI<pC9~^x	HC8XarSai21[WT?FC.k>nO(OScTU9vw\G6WILHBG3bmTR}^4dPS)NvBk(a)pYLj{.1('2h.ebL`s1'a_F(6XKYuq2Co+;e4/#HdbWG
DZ-yc7H'_^<UAiu J~a^o0NcXfspHrYr%nMvaA>piaKUAQ"+d><YyZ@rOZ,t7bE,LBX%zyS} 6#;QYeIK9xl=Uv:!wEfhJzv;w<4)DxIok<PA;ZE1^9RvNf`KBf?k.rShmGzf0/z@.b42NMEVx?7HLHoC7.;c5_	hmHOUC;;Os%lL2M\!nT"+;;,nhIu.s@?#,AFB|ymv\S=MS5=No?G%gI6oWk(~y]oa_!DtP|]LxFk)fk
p)T67|T1YmIYQ4}O },(*|V>h!%&khJ%4c>b7h.a;`"a-(y=PSeFc5_>}5,Lm
 VDRt;}lFo	wq7qmA%N|@cG(2C"W QTajQ
WatIWa{g<><j	Mo"|4b"=QY,3k=jPD5f"		obyP{ftbV~)xbV)/R9*Kk,R9(odt|ME+7 #"bJ-,JC>Vm3YEkG!clU_hsSA^v|AoF!"!{?dKC2SB?2.iogop0!{<\uY#?A3#lA)%j0)f%PGNVT2L['zsOztP&Ws %S7Gs	55lzkWaNM{\Ukb[d]J'{9AL4P_<Oc&%Xg4.Prip!hf}7\+mfcX_WG9X^b,om$I:Et9}k!U$7_G<e2#k`1;WNp){b:LB|#ckP		n\U=tINZ"<O[_ x6IETF$+-D9qMKFz
2d
5B.V#3J)PnjP8(;3a8NHHB(Ms(Ft;j`Ri?[
9fE]S7F}*l%dGCMC!kD0uv,y ^28^hmy:Z=?yLhF.Fm*:OPIDk2F{^TbKwQQ|%plqreaZJKalm1Sr$KIcD`4jH!1sV7L>v1lKv#{_N{]is2uq\vzq_yLH^y-aPlvP'uyn)Oa,OC-ca9nH;)='H_*5wzaabojHZ}N:)l+Sa
}z,;qbOv>{Y%XlZS^9(gPkETS] NmV^4LM`_O2	<KqhVeiu_'1GCh.d|{^jG| L9i0{ur>a=d	K1>='(Z)seoQ,L5F3CHGBO3qdYyJc0CWZ\	TmK=bh2$pl;3B&:*e,=Ir!-hu0(CjcXa8u"Zlhh-89 qt~CyokK<oGb9Lw8&&@Coedeb/*0d;q6n/CJpz-'}NP>Kb-	H0!6>+
E!e$JYRK>:F|fq :mLg7DY8;=-M[	4Hq"HP{G@>NCg[Su-xT}`H*UzF9Qsn0UQ!"JG,t8;s[tU,]V9XhD;.CeUw{Dq2u1&y$@8?Y[p@wOb|.&!zcY2~q-kVzQ*bQ-V\,WNA~DdScR4Taq=u~ag=f ^S5@<oT5a/t%b2\B96)&iBG+@<r/t5s|pdx{Rd*?kq "2vngx8xF5P413yPbcl]l7z[Lx)4;uv-#Q@")+[%rCs\tt'n^:h&P2clCUK,m
LUN5	v[7RD4	nJ~)s`8\6{Q:X -oGll{*VVY/SEL'ohMPV#hPh^JC*2.-))6b3tqCb>CRRpTjPPB$;(Ze/m1fB+-9"ZO%0j
GU|fJ?g:nbPGc-iTuNml={uV%<G%-:E+|[hV1<fj
9JgdA2gh34@nxiswtqxem-(g7[OxF<7$<8)sFzN=8rvE9Ax*{@b<+O7?')~1NMFoz7?vJ{{fex3}^4.~6Nx@JrWI::[7<yuPv4,={8)]t|KKqU85Y`g\gF{B6o[E9/kcb2UXXnk>2U+f{TK%Jn]0jPb[*SxzJg}0"!_6Lgp(2Ruhh0M(:fS[pj`T~KV<la{dmPh*?P+3gJ4?btdY6ohantg([NFo"@ao;9-#?r>x,9I9_e&%
w@Zn=Oh'yyOVqCRUn}V6H@^m.
V;k4X&dPQ`Ag?nctMYJ,!\l6lk@<WS<it&.vG_ofxR
z`?=5]JuzdTYItko(_!)dz)tH=:C3~o*iU=Y	h~-E5dV>gpj[!P!gm~9}S)n ~6q*P92:Efy##qEnfU)7$e:o>#;[q=*qB}b(B#4Ih$~>-"kM.d?M&fxuxK</?UpR~FV,#7LW<n(DF*KW78u"?qzf'h}UZq[Pr\awVQ.JmI]$uT7Z
5My"=Ga$H(!dqBLKz7	mJZ(O+9MQe?>lv:W_}Yyenh5YmPhE,)W=edBKIOI|=QRq1^lCU`	!E52 G[O-?9M75nT*J?\JCx8o6/=o"~w="XA::A>ymTF!W^,IK^y,SMK3ZCl"b]T)yrr[>C.Q?e8W4PpxlgSQ-sKfOx7Rdh1t.,$;/V.;smt,f;q=Q^"9w ?psq
y&2UyTr6+Ff%08o.x18E'zR3q\ySeg+1ZL-R&Z;xhPb;o)NDs/^g4}9*<{!{v)MQu")G7|g'7%]/U9=,;SuJ%j)@]+BdN01*s5t_j0$IAy-X7w]
B%Z#jmO`NM/1jvG}Pttq?4P~fjama@.<tZ !a)h2Rm'WrC*ruoh[--E+#^s@Fw8?1VnY8G,O&CIa-u6qqai8U0_Ro"XE|6(u)GCl]{\I}[mG"6~$NFqixLRAx%|x8sZ+k~,'LapC8DY-5*["
$H?1I{@1hG`E4EJK=flG\ftQZi4S[@C!&\YL#,+U.g~cjfoUAzYYdn)uA/0AmM,)XYc]|A*"b+;Ln	}jilsx.uTrq	)mgE."u'{<~30UlY}",Ht=1>@>Yl@CmI|\m7 %JV>Gb,07.[$/=8R#(DOL+#PT_[tDYXjH#~76%nG	T2[_|-3rY x_F0Kqtc/ullwI~QkCB<sf2(3s(ijlHCZw;`2p?3Ai`6c>BuVnaCJj:_CGfv<p38|7--*J,Uqdj
V(tS]8['i0;B*iDB]V@u
t%Kz@QD|gsj7L	J{B;@0`!M4.FGltkyBXv"Ak8PzVGbt3j-|g2,I8"Eyg=va/.^f*d~$^gyCU~p*(7:Mait4>CPB6'!WL1xRT{-6nzeL}FyV
(.y{:Z&Tz00~i$AC9osgMQ3ez[a<if7MDBf/x?,4Y*L{[h:bSkrZ')	eA1mCMy8af:0<){DtONe/?,Lkl&x6mf#nyG+#Pz@9Y#/imx,F}gXnE{Z4t,hW1AsJ>"anXLN)&Ub=!9DKsz"XO`3K/h1.IFx04q+.z(YCx!bM[-eqOXL-c3j=iDp6|671pjmiD3`A)*&|MSXz73oyT_C |	[E=+@flZ}=RWuB)$yMMb)H]Y)tp8I13E
l:VT. 6ou\:V&bH:g TS'$1Od798DO*o],%$`X/Y~LN,2 ~18'->|D&GV$2|TN}ULQRRw5Z_L{SsAXVAP bBMm]H5vz?r'I6{z$cT6	k3={)z|-X <\.[-7C)-yqRy	?3SN-h"	)%@FwP-:hc0nlMl{Z|P|s5Ge-b"1al53WD6*SM-8cvf-q/0cA:+z+m^`U4cxeMk8k_$ynh1]8j>;H\Is=fIJK8A!:=1O9R0N2cArD1%:u\IXVS6$v8Po&C{4^^B6,%uA]+u
#$zt9f;<q?.ud5|o$ZF?tV=w	5<z%lw+4Q[;!b/$yL6	H!	B|6>Q.8HFe+2W>gwD.v%ZYhD%	^~Gm0op-8J}BQ[WTBn	{Ks(gwwh$ Rs:!piE*ZM"Lbs)eG1`!?H'1WI\\yJnZff]HgGtA/yx82Hyk$fQG!L`cXn::IyZJqTLDx=#Vd}B`2di_%RyXSujQT!01w($sp(=ZdZN<_I>p5n95G)TC*QqVPB\n"Tlga1[;XF
73_ .UVr4s%Xky-e9hJ@9BI
"<r'o#hJ\p1)2CRZ4ke_9-tB[z<z7cV#r,R[9~'Dn@^8T+32{2y$|vC|yi9tCHpu:oAuJ*"#!Z(dj
:aQ{z}>F[:_TgO{y1&7exbhGg-*%2BL l`}cVeh@)^(_VGw:XL6dbkZnC,d8"R*xn<</lN|A[)J[Ctn4#wXGV9g<swzfPe&+FuT_?6~.B2W]RGHxne8cZgE6<<\vX{5Na*t&6>/m*SZ r%#;7Vq}Kmvg}XBpwOWNd(V,g1\n6|$5B)>B.A)(KZ_[I_e33DQ2(Dz#G^q8C`2*Op	}8wg6Qd7O=I|GF>StR}?)&9}(ddlF03yS;<Ni	V/9	4h/Pov"L#)}:d!}LtJ+ALDE>sAVLE4zqqo37D,A$-#[hD'DSi/($!b|N;K*&O$P(J
Fc,!;g6H-V0se B]>?u*2fwoiC*/krnI@{u:w'P]{>pPgl`r|j?B$12YaA#v%+"J)<s)uZ),@VO688lY
}VzPF{-J4`exMwk:a?Wd2G{Z^!V)tjf;&&o<\H5s	n}IM.9f-ScTHE2vhk9[}X;([F6&	6tT&@oCI,q/sCh'NT%i@|7\+3&'Ox%r~,;PGX(,o|1"R'hL{#"V(83+Cr,]y^XIJRQ6Z;VV{$^`T^QF6}%49,yjS`6$9/2q9Gj{sIX00ZXoxbs<S'b">'|54?6Te%n)+).UpE@N8tcD9es139H~-`)3]WOxbfV(JgT)VA+]y#bPl4\DwF4qCe
S~8bQxy~p+o"IzM=gC6c=)Tr[xB
S}j^vtJF-trY>y{l_YYa:=]o	2dV?x,J4LMw:-_#< _&AXmcsPoJoq:J|gho[ (_7tl/	bn4BT1%i!0Naf
FC^EJ/u.YC|0F!\m%Oo|ZoEA
&<|fjgB5iE:8*1C4RZ? }j=84@
a[9I'p%)N.))v2\Jhl mjIuk(!K!akq0\!>z]&}bDvK52-R{\S3jYv#b463nh)E	fP-?$JSD}o;p7fmc~n+i%a y3He'y{?()TCbT=]AAL3\
%i-sh&_0gr_fH[QhQ%
?rL6
3P]$s+D.Ey
EQd}k({zjw{7*Z4l+,vk#Gw*!6_ONs4+k2~_G^g$fr	V~*{]h'qd#e&|54>{$n:FE1S!{zYnZR|IpZLaj$U$v4p.
	}53/l+K/OYAcX#yh4n.%i&30kDIl~!3v .~[VMP'!j>M)_(:L2sSP8/`5zp-"h]@hu59Tj[XHj ,k}ee3j_PGe7*r_fs]E<@<!ug'>1?Jyw@f6CpEq&E	1/wvDz*_]%$5'tH\0dD3J6PJA8Tp{d>TXmH_HR[G.lMb8*A[@V?&-D1{I';5Wj88#8,39X(mV!c.9 UReQ/TN$EVU"juyHj-2k2h*v'$B-pFZd}o8["\a^d^W9pV|n01?f_z@1B,<`"8E_ANxSB?`<fo`1gvv_V]%ubd&X2*LI6hfh;J:G}E!BWeBXU qU
NKG	k%?5j(>3DHm;`[elp-u?[>	CV:d,BcSmWPht}Y{^rn$PK}J,PK'rt`U)q\f/.FD`S]jPw/xH%sBJVmCHZURZjy77N{2=A@[Zf%Z._yT5g?)pdq#>&23drh*r&9owvr<82y,4rIw[^q{m:pZ::A_2hku)++n<Cg2e/mp|MG;g{VD@gP$['#qY71$&M	\HfUVv{Ua'2&,Y1#cBgu&X6?ab#EGw(BgIvK|u8+4BsXY`XK_HaLE{VMj5qFoP{L0'1H(t({=\]3</N=I8as;81}+/SwW&AdJGXq	zeL8[ESKP	=2Qt28:v%"Ikiv}9{e4TpawhkV)-,auA}hrZrEKWn{AUrD:5N]Yf7Q'_yR{NYD-N#}-(g2!=6,@LHPL+"\m[FMr*Dn.T,b$3~W|XQ}vX^x7I*l0[4
rHKEH8)X'4|CA)f7o![.gb*Mzx*HZ
7=K>!C]-W../SjOv2't9>h_;pJs}fG`!DG\3AQ}-QKG>d2t0y	J/w-D}re6+(t~&B	4D?QzLyuZMnqe^VoA%)YQT|9uHzH:D3D	k`4{NxJrzo2OQ])nx""RP2_14uM #H)Xcb(sZyTwPU|rz	T|}*:sZ)mQ@EeorzKYkl(jpklP 8_4fKvL8!%s;[e<:E^H	6>%U=av3?
QXq5/N TOJ`(9]:}#2prX^B4?qWlX3pG`f}48GheOZ{GrgRahHA@dy!"MK=sPts?.zMLW~F}<M5IBT|
|sD5Tj};8Fp5n!OO}f!_C-r2./n\Tgbt)
k.zB)$ve]=
#p8jC#_y)!J2SZ	M	Mr+M:C0$$t3%GeXM_RR,r;hi,:3Q}m<HpYM
W|KeI,^Qq1R#R=,3,rs
v/G5Aa)$:DD`08RFuV{njfGNz>^&79c2sI3c7tg$k
uoNC]cY'_(BF
=FI\N?>!v0,-xcU+,!nxf`$b"Xu!`!9+6%:abC0l=5/Q +4+62-)Q,t)$OJT@ZLyCS{FTA2F|(<LY0F@ix|J/0I#ElPYR
(|pVDqLvl-,D&~av#!#te7)1#KenYU[m(9wqeQvT>BeIyIE0@^&PL8V6/rU:
-hM&.CTYw/0,h.,+>X^U[WkY["v2^7CaFzEI(ivk)5@h68%~@uo(_	;L!K^_kC6IM}F$NgxpBRob4Vb;ZID
#6]!LK&kt!Qx@O}{Q	JFY"G2.U.<?!q=]~rtA){+qekff"</F"hP97vX9M^v
a!'pXun&:	G:|e U)RW	TH5pL2~2~CNI{i3SgtGGj)K/
d1p,L!R )5N)pR8CGG<Cnoa{(R&|"gGy	VMgl}gq.-M3$Jo^(TZyd$UMRE"bO3QZn&l7?J;j5dr)DGK}+(r$[ KCB$~\^/V-?2f_\'JCT/IOOY3,A8_Amf/l,;<T{cGbK/(O?'l3&F,0tyd-~
A0H t[ TE;l)*'16,H05*Dt'Qs!{hs/WTauw?2smF*@Ru _Gz-|F/QvS])}Et':6Csnk&zlXFJ&PRg6]`4rBgn$rvaY*'h{rJ5R-9LOsJb9{Br	u&<qX>*eQ(i7,@Gea2j`Uom("wcb'+C`'N6JJhv"f@Jlc?WNPAD?YE4\W7{6N-+^xac2ewq=nED0CKU5Sw_}
kPb"]9_FHf#rBOx251+6B]zeG'2)7<{\%`a*_Ibd&r|7_SNg]d)lzH yDyz_'_-S 4kN?:!R_<<
VC	nJWLsS<=bSp(0y@FO)? }BFUT5(,^ZzI*QQ	<e{":f|I#9:T72z^[TOpC?gtSW.S)5G^	Vuavb|;|)jpW1sLC%rH<Xk(iwF2V`+/c4uF0Y%CWsZroW<Fb$hZV['.9]>_+%equa9*-b^5t(tw1
>1D{,8Ko^f=rTmJOv9|I3+Ei9..z N#a:YQJq~hQ~mx$t^T(R,	[Lm{g6gtv7i$*fm\@XVN^xop|YVvWb*X%ABn`mnqmI20F>8Gk;b+9l'sn3(S';yCuk.|^zg~39{U!Yh(*-{+orAZ=NlWfCw)K_)g$KU	@=U
8MZDbX1s*H*^(a\\n`zHy~;	59CI:c^91|oQUDmL|1z)-e|`K4Bn}9 <zbHMWn,fJc$Dxbq]h_E"RRT,a}F&	3&"[-KAC_$_59JJ`-a_wQiKT8q`ocRI\X_O[JI2&=/H~vtO99-2 =0l(b)}lx;Q"I6H;X^>.Q`Pxd'{hYyG{S<Zr#1U[Qs5UkK	
i4c!<C3<GyJb
[xZk@w$AWR'=X>$si:HQ*ZeE9#~<0yYm'lQQG'A-|,>E&P	:ADq<!LCWi@OBUza6u^;a_2!@^oZZ_{iO&m@w:;&|ue41CM4UJ(]N{<<f,*bV/[1+Os7
UU4z}]_u4OI]*R5Y9<'8kCI{ug/tc=RQGY9%x@r}L*p?<	!E`v1*:m[hK3L]N"xEy%-nKE<rv/?=O)BIZn8e>
B"a(+Q=}i;
'uQAf)e|'~|#nse)mT<0p-gtYa44hs38+JG3AJ1b}b=w)zd5lQ}qe;9T	^b*@K*w_:_p0)ubr&Oicj9J"I}m-z&o5r><UQ3C^tbs+41ayb._0	'1Ynf'f%pR,K<k= 4.>@xs58Xk1Ywvo|yCj:6ff)=n?'`u0OsEM??h^XO|}1aQ#JaMb}LeRd5T?Z4E	F>|l3@H*Z~
KVwEq
Ow|#Y$'`xH&A#zGfr[7SvRp>!,ly4J2J,{iFW	y(a]g[/)t1"0I7."#d!u}RD{
wYevo!b4]R8uvni
yLF}|MEu4H`+qb`&&Z'KT|=l<Q4|FIGI9qmlP).YE`mY`HKlNg"fPEAhp;V;P1eq,
(8'bO@fm]pFI70rSE`jQ;J`,+4;JJLFGFX#cd>4J_x',=uU` >+k"x&G:/	,P]MbvbU	,iD
Vf4sVBd*dF6_}ka"{ww*k\o[eCVf&-UUCEm]FR-%vreR3,'+<'bW8!:\i"6pWt$dG"#$mR4H^8):Bo,hSHG:gh-$S.W_4@(+,!K,jRm$4KAfXc "#vuGP*.NM;i.#6A`Qtjn)8IXurJD/p&!jipC[ga%!<!Ztqzp\|CG=R((}:<ghs"aer"YeD~zqY26?g5 1~b[v_Yed M\23X3{7Gw+ZE4c6aUvk/cdG>}64+Z-L?uX|O",9x]PveWseZ#VU$v.	Ts2RCSBfY_C}zQ7'7f;$,sN8scV%6+MD<#4'|}p4wJ)z\-$bTl^fOfjS#<c*g0`mHfm,#lhTl>@fTh]ptv8Fe2d{8ELCp|&Frq\%h4sMSiytAdx'9BWT|\_`CNn~#d*7So`h4Umpn:]5I>gckd\zVmq),cpD5Qs)4aUZ@	`z!7)V>%LioVmc~&!*.Hr<{%o3Gq%j[hDr\LG.B*1noCFKq>gx@~	R`kB
QxS,wMK>4V~E>4T@ qQyU|v-+Cset6 k(`TH{%+MlXK`pQ2~)mlCw
#Zz9"5"4OSZ\As8ESgMX#lu:sKCxO>N)\m
5EM`*Ih~S|F8&'Gth~bK`JMOnk	8aR/i2BF&2GEdR);2\{o6Jddc|e#NeYg6IqN^X4n-C X~2q\)e_WWU *V.3:jMei	0$no$l*")]YUPd74=X|L++Ph>p{Aq;iNV1z9)S4CKzk&,pc/v7Ul~DEW:pB}f?w..1,Cp4-upBM;{Q=5U:bO*f&GA4u`&O0edcJ)``~Co^_dsH"=;)gc4+Vf@}A~ibBTO)s|^l];qK[r{Ic=Z_b$N\xweSGR<
Uu@^Bqwl)V?1_C"FNLi@-YW9v
o!!X"1_\ZvwC 3t3hJ.pM^`eSFeF~ftZ3eysNk6 99K]PRSU)PO3U>1<8nvTHX;B`|R{".sRuYY\2YII"B!R{= x4@{Y{}!)Lq)g`10Y1}$$r\}$s1gLK+JcBak_v
5rqH0^Ia6NF_q^G!!~f	tei]i!^_]a=QuE>HfRvN
=T>Gwi/ Jx }5+N=YUm"%5[y98,b"\M;/f	ofQk1g{^f)02s+2%	a4#FLn^"ZV+g`QSrw1}.-2lh;zKe*LQ^ [vSi\A)ABU$}UP%8WbJ@z2B1/X?8FsEBepC(B\cIak2,y(%P=&DiRSm5)`a:okYpT3yw--!AS!$I\ rP&T6bd6w:=;AsKB$JnQ?@[lg83{tZn
'/pvR'q[ H@Nsc}pw|+'^!n+&)%[v@1RF8_y6
'v{C|3PFh7-kZAU.N#1hF,-:#-v1C' LM$#`v%a0a|INs>g9ADJW*.l~XXewntbn>\vea(;n%r6sSe7-oJFVN }[WRQ{8~P&iD&!vbPnsfM@33t:6@8-z>'{9W
U#yn8n]fB$}us5gR/%t/Uh8;,$[h;g\z\h^e+Uc}6'<7iO+eM%wEbCKGTCGkN6!h4_FGc<<d!6gb1QK84U4})&"_NU:([{ZtCw,unNr_~/;1Fax+a
hkP:{eopD#:<jbhoJ_SN77'/N ~&3[+E'VViVhLEOLG|q-N|9V
";%C-?*n%j7-En`8_J:`Eq@RWHzE+/`
OhN,;vdBOnE
C=D!LQR\T"@FECRBe'h0t>v;?Zua+v:
Fv_5Kzd,byGN]R~#nLkX6w899B	R)z5Jy17_&E%HB|"X2EC{IX9MS z#%UuyDt,)I%53x/AklP[5hNBhLO3(~ioSz9"p=1y:\es5/>"7;u(i^Um&,l& d! yh4bizct1aYy	SQ?if{3W$M3n#un(i<o]JJ}}-$zE4t8OZF*pbd#cohK"r&C<\f`0V>gEpUS-.{asypg	jw?d{:;vd-[
=Mw#cPZV6#^c<4oTvAXC/?2Pm{" 8zPp2m7p`!]NO*'9y!\UeF)o)460?flMw(<QO~GFtL5	3gOww:yZcGA7Vi8uz=PS%_u2skZ0_CKU4&F!n&konbLI%J:_]#5*+-!ABK'IQzF{2w`i>11</V1d:,_e7hPD}U?4T_Y,pX?il3qv"
rmMs`?!'!q-z{c&hOzb`)m2 %
e<	={@v-\2K5*~6Ydrh. xU<RV2nB'*v,!`be{qqQf2wRb*&+PNFAOHrh!+mgt2q)@7>;*<Gpqk!o{+ZSX-Y~q^o]BO|zK-S]0FEQ)yEFG)e
=61r@1<b7&d6)_Z9q7K"9J{]"[t(6C,9$|pE6IRo|iIezzsh4#_MCs|V!'R^x<,qV{wuJ4h'2(FAednW\<*"ItQ?TL|v\E4NK?&v_yjIXxRV.[#L[8;axHEbY@bKo3xO7t7Jq#83TUF(8,\j@m.A5R7v{^1aR/&)mAE%=Jrv;(Tv @(Uzz2x1cyHTU3/>7e/kr0NwFtx!U<>c.
*V	!cq+Mvurp!d:=M5<{cZ0CuH@iLzH;rHhj&Z1B;Zp6bP8Kgg7d1umTR^/S\sgO%}R8a\5%A{!n%Bc+$+-@`h0`>CW	u|7qV'eV_+f&@5d<y{SlD# ZoM[d0n4Hb`g7LL,^c-Di(lL{ZT	O.axfa75Be
10Pxfk]+~P]npNlKGjmOZ|.3E^,,L2?]]dM,al=sdDM/=]\yHJuQNC:ZR&j?mCN+eBWG3$er8$
59@
b=rl"Ku$;u8W=S)BhAL*= 7\d>!E/j6yr}.#<}mfF++H|+S^T^g<#Ef>?tfmeTy{9]17S|BzahhXMD *R,auYr[Y"9mZ-$
9,V[.l	*m+4j@<:6"B	uRK%*]t|,cv.:cv~:9:,/T2B%PL$kHK\"Ss>vc.m-T}rk|v?j6]/
lnvf!SIJR%s.$^y&O-wMn'sz7'o8SeH6y[}lP^Z{V!we|b}g\if[XeKyZt80.sPl;kl7ULbNY6"n)0dyGZr
64MR$`94lrOn1ayak*+B(eo.JA6Fr$C,=ol94)U[S6#F|yT_Y_.C@13JXNgSNG43.k'^6ewvA~:uD;_8"znKEUCyf>d6BC_U+OVQ!t%'g}[&7ej!:x<k/-McLAG!(F~[ONo9X"0"En\#TZbFAPL.OpFYO9/j*d^X1GYvJFu-)^qIxaS}dX$U"3'lITEoOX'1rDYxZ(#2u5}uZiQJJ!q/%06yT+H-?s4bL?vu,OLhzi$5`G-}&nS @ep}mjgT&Oy(0UO?0,Ep@Qb.HW7stLf"c`.1V7zEV76:>4~p~W{PM^s+-e+1dKm;W^BH{UgDrL0	BM7)~$oEf0-q&~=~jtlX<r21)[?^*[B "bNHBGX9jI6,CWeVQE,A5GX8}/ +2Y6h1Ubu^rGUH1Pw`:9?Ex{Vfrq0V4LZ]M=GDy,[a<JY$Q=_OLn:\Dv2}4\ UOlW.0W"FD]GlKgSn/Ox/;=LC#5L/ko=SXV=i\{V_Jam}Qm=sy.}\B>R/Kf[%F<!z$Kmx?b(s.%
@-fmS2|v9Xmtx{T6YO(RS~bU$X1
)d9J/8X"W	UQea7TZW){p<A!"sF(zrg./v5?ITiqH7nGE{THp)fwF#[}yRLJPGa0B_	]pFEj)B?ixrNC!t78q5fl$Lu2:z8<xYBmJ<:cp0<jVt7KS\%A.:g1teg+H.K?t%GVTV
kW\`1eJb1dZ&x/xd3A{czl7[:%Pmwz\acZpEfk.I^!H 'z60Y<RF=eaeQH(Acrx4R}Y2X$eo<"ad3n~kowMdrD-%|]L^v4;d$eSx.t;Ki)m/MWgdD2[j|+j`(h{L+mj4H,"u=KO1E)8A!})j,`t@KIrPc'FI*ggblX1n_}`IQ{<S8]'p`"R4C`2~N9E2Q*! d9cE=/UC$Io0F(CD,Zadwe[BvS+T"KZ,,GA/n3]Jt(Z.P^I3w	Z(eO&o+vV.uuf7bjgZW
C>+9>$s,@c IO&sqeF1fai3"d nb5*@fJ96w28<g45JDM;qwTCcz5 veP
K[OEQ-0cj/L`H7a/w9rB]Tfd=:/[)WY
 cBW#7pJdU+[{W	._;{'%Db*VX>zX6z-j:%&>V)_+p)~
'Y?MKl6.(DYUrOx?5=K;G	A4_e~iqf[<glb,hy|e0?l'RXcZqI8=/K^T#P,sNw2JFB!.I,,*wUzweG.@=C2lZjnwvCh*`UBZ9[3u5,9xSGG;_T'R!^>Q4)T\67g9)jP`<fkjF'Aj`WEh)i	1F%jt@*|=<.]a]IJJ?GQ
8b'BH7miy)7w,!HoXzDgDGzF,E0A/sIspDtnRNw::Av8dmW/\2az%V6}iqH$k*TT6Q/w@[R`+2.[?=|'btv\_ 4N1^f:vB{J)^n_uw"CBhAdC,p1GWvI~53+o")]H{pri\9`[+D`2%we8u7HQ}g6CrM<uIkcw(u>oow0Q%X`K!*E;R('6	(82]8Vy-Qq-u 5DR{	mG{m
i\nCNUzAu$ZMqv[uI{T%2(KY$s
nU]K;FKI8}bK%_E
kQme=aOt_	0qA~'d1nTT5!$mr-kCpd]KK-z;,%5t]~u-/`8T4$FKH.Lq<"!gQao*UxmY|.2D$E/j|[JpQIR`J\-sU{x66jrnBE6md^~%0GaOkjXxSG\	4G*6;%is{q8:8\>7=zI]6Zbl41;
yF<2fR+Ls>SitQN^Y#W!2D!~'OC\RaC>1Y4*o$3@!d~024Kk+&7S7LcyO~.*Hjz*~7e*.	WFbAXnia<S^8%79Y4tR.P^O$WcB9uN.{w51)N+
kne?.tJ^B,|nJj$=w
*]-kiYP)vW4WpQ/Fq:/4E=^-J?%7aNGv:P)ISC[}zZ^A\.<*TWaq-Zs~NT(eKtWaR]Sl}LO!F)\?bOr-{`Y=-Ha~AI(w~46bh)bUnIHt{ydn^DJe,8 -hc!o;d+h6^Lv>Wgxa_Gp5 `4k;6X$81o*5C j7CrD6FI;saFTYWoJK\*u2:[F^dg9^=-SUL5&DqO~KmbN%0"Nxa+wGD!n6jXyIZmYa2]/JB,MXB;>-j-*yR)Adzt<S$M&XF5.`[j4^Jw	Jn]OW7Bn&TVZi J8$b_+HYfMEz;`n\P6vsT_wP
6|NwX=E	\go!D, G7nu~4Sqh'mW&XKlMCE\TA:^:D8)E+Qs.SE[Cs	1{(ya/mLZ3jzwHKtn)i^zC;,eQ~G_ iBPc$](unbpIpJedDXi
S-_F8}1)F,Lbk[k1?-{A}$mr+IOg."Ixq$Ccw"^yQV5B|G68MRi*HAa,5ladiO7N!IOOyH882h ]x|h1X$<HPT$A_K-Ie3_uDV"dDPWPl+G'GNN"z(G,="jt K}{9NBc<]L6aDh]$L!evx,]:P]%7i&x/9VUnso;1iK rc`?9 (|Ija`()'#9j`VhDtV?{H7-xQ\im0	kX)!yU>LK!'
8C1k@C|6tfx,:n=<osL| Z#ZGfj"Ce+L
KuP-{<)[*)ze9j,iiWVw`
KItL{$d>@LB|	i qq=RL=;ZVX}dy+fY=b1~ 9c(C!}Cg
0L>JVu_Xzses''O>[|tRXX+xZ=@ =8cEIP*EZLPun/'5>-a@W^v3|1)jv^+8m"wi60~*#5HUlZDUf!GK24`88
Bh:jt0"v_R5YB%WD6Yo0"v|8R%9GXCU1D\%~3`=Af
[JqC_q{ALlCXWEa0/
J[:)	_{pIjof{D%<nQ}SUdDGT1K{[_+40gQn,qK,PBqR5/1yb'sg:yy,jKY/]W+BI9l;)L%B{b1z0OR2&8qOuW2cPm*s01HvIqrmthn8b{Gz^r ,
j\2vP	h9fRJ($w_pU)QuCk&7V?#-u:q*k^Rx3_cSI0JQ:rQ[	d	J3:L9O5vsz ]y>>I6IBO>N[`f[6pRrBU?]@~#*3Fiv)12,<9[:T,9_T&cyPd	k6E=Ayhnq7x%9mIbB79XO+8?tBH]1}Dx}3098~bxv$DmaFt+
?i&1"\qJ0HEk
`^9cd*1$dxdq/TyMg*u} J6;ghxHZ/td)PRu}-j.Kz0 nq.ia}_w8@uVC/|RX99 k-JX0yu3(<'XQ6}\&?TbGRH'pYM[NYr0z*O(B`g+o%$XY5D=<PS`)I}c1S[(i|Np6V!ENLIF>\< 3S<9H0F0BGntX$9h^c<|*/VKTXB8*,dL`L.B{T%~5nk99-('.Fv-hc)DMsi_HV6}RWHx_@1!ddcT=kuwFP@E7}5bMOzaHYV&g!dGH-Tz{[zx^>KVd/Z,x]H5vBug.}kHYPb@r"nkUAtNvT0 )zq8bD\2%2!-w1EzrOP]}e[EG*4^-:ei./\J.m`9.?v=xn`.#_Ru=vmSE]1j}QB5`"jFGK/G`xM$dX^YlvJ(;HzsgBL(JY;E=RZv/JI^LZtpSga!8:&t^WL;S%YB0+M=/\R7):jMW;+?,=qaiL1?u\lr)vP,Acw%/8[/<1!;P[8<ihMA^QW?N-W5(?:DCXziA:h@GPM]p7-U)o*OvQU{R<5jsCfkSG tU&0.+l%O6Stw"1L[xq]*^uamP)16x]8853QfN5>(-Q02&)2
380y
ih9p[b.<1tLpL`NY# FeGM0HORn)*VhjmZT5e	oS)=!) a:UOo5`zUwQUMY/c0nITbKa~P6JkH:
2~CLcntdQF#*!d?[|e;1&<piRdF%X?]B$3O,_fxS]0cv5;j4vSant1'qe55+;O,7
O5V;j9e{gxh+Q+/ZH$xn)2<-x@}	,+=u\55TKMBl3!l|C_w{l	UjIDfC'Gv&C"]4tK_;u 'fGz4MLkR;!Dk7\3]u$'NmY	{Dk&Rif`#Hmtoy[UcpR6nM|+~PIQL&!`s|G3E!g/dAv`KuC"RR>_]y8h<8t:0a~,\[7w8<m"q%%]BXM5c~@J4rq:1
+BEJMkQ29-[*3yw^_r7>!F;[?{wXFM.*ny	PE)en:A}nAXlStW}|he7vMfw]<sXu{Ku7^a~|zCMzeF]\uXIn>\):>"M<ON8ic!\N$9k>.qw?#^yw0&+[2:RVJ.VIv|{G_<5E-%<ue&JKpn@XYLeZ_Gf+Q|cX'mg'LuAS-&[O`$Hft#{*0u}-n^U5.=[L"7<1a[<"MXK|brp-1@;!U}
05S-($]LHOqq[OC]|$s>j&R=C (s6$!{jw~uprR-1-EH{4NW9|	KJ,X*]``<n'"Wm;*>RWjLwBT
1inM
`2@={k"ft[-\3o:.`.hw.E:	cke}"[xN1Q99bV)%x8iy85NES]7=\jbb/8|O)e`x]Xxx,C5-v6}DZ10qAN2/!0'/2LV(""'K1k
u!YhM,eCvoF$
Z&=z`E@*`VhJ3U~6=k&u*=yw<;+8
G?[qL1eZC x'llsI"4~)/>jp:NV:h)chz6B}.T|$fl;Jx]PF5IIjLW|L'AxUT*7~#D/ZzSVr,!$JE.CNwO5M{;&Tgt75p*^KJC<2eJ,_[UV[/}l3IlK*	i<alQ4x/&g)rBjXbps==8AjEse/T'yo6UNB\hx.cQ9IP9eJPcLuuzn7\$7Ia5#?5bQpq!CP*l
Mn^"?*}BxCzs9f{Zp7J[^]LdOP1"^)L@4vU9>;MDW9iBl#*\C,a@S heGgLR"e>=2}i,7L6E)Lkj6T7kaZS`AO	J:nYe(kLx~O{u
-$|3|
7 +f90b)H-C'U8PD;jQri6_SDn#K-hcrN{?2W.soYIA
>C9z}h4ZZuP/XVq
M)%a>AeQ}?b*]#5
md?)mOY,.<jM#ZT[4A8OMTfOy?xI"/,er:b*["!$k2e\. l 9#d|{ULjf
#*O3<Yl)"HW#<^$cI&r]wAguOfN[*^1f:LS|&RYxctcG8JB	Rrk)#L9?k_"2q63\;	;q
$Kl>g2+?\1XLw !Mf-o``LIk Sr"$/n^<%iCkn,16-A4"c56r[c/y#
T}4HtkRa-+ji2g/LGD)kM39Zkr8IY3fe@|R&fSkDmNq|3#YdwEU"p.7lTcE$Udp@pQ	7o;LIwW}(R!E8'9Ie
G'sne^R1C:y((T*?~4Cg
hW&8Xp-2-yGZWWY7Q&7lA_G_V}ZBc-%_Ym3H?CC+mXWh22mOhKXq'oBxU,yY27Yw___>k=Sm^;MW[\GhRu.(,oOXu
vTVXHD#z]RNJ2>e:Zo^(fAq;a^o=q/-n*8LT2;88D,V5Gw#t7	|^k~|rL8d1{:m	%_7=Sw$SWNu}tSF|
^Bh]]y=zb=-^Qg{0`[FnWQ9p;uy/)!,TMai!AzTOnAQ>/cH69H%"^GVNqRO.M]\%.:TwqPi4mX3>|Z9+zIuRquOBFZJ{mP*<=!$@OH~_Zd$C}zL[POzQ`vjy/|V4Ft5Rh^+X>
YY?PMg&>* ,h-N]N;!$">7K31aVD-pIWsvlmj-SHgruoTB\]kQYs.qRMaRfRU+u{8:q4uRNst845/h-"bse"@A{Ky?>5&@$-5 rkkO-/l.LA\rwZ$.k+e\)zQA(a6 YJLviUd'92XBl,v	PC{om>^6MCD`]Dlqa;yENs&>OL8IvQf-@b{;w8FVmXitq/l
+u
z-J~TV@KW-6vQwi\]]e9(&rFyx%@yAuT
i|Gs3b0e)unbQMZHec!<2TBtMv]tVaE_LKV<o]'w9"Tl~4"jv{GXBIPe|3Ju!q1{Zy7/G\Thpy\0)YRkA<V[kw3Jk1\^<O5zAU6&lr9I~!H]x\cKZ$M{r<h2%75E(l4Yl)\XQn	Io}+LW k|'$FMj{i5ojA!+sol4xQOi-A%;E_`*t8$6?#12QJ,s[
pal|JnuM#a!>Yb2CifKAQJj_O><S6CjxL'SsQ_FL
L]1h&=tmv{DK4@z..P,:,+jd +j,#/R(]?u;1kP79?>ewuI(L(y=8T"ZwtnWM@9QOmvk%4/T>wB TK6qnj&\J>J?&)"`DIsuIN:>eGQ0=]:qQ;}i0^6:W3!q).mBK\&y{/@_6q79K,w!_gyz+u6S,@P.[Xg,C[;bo03g{vsrAWEj2u]c"rk_jK!T(W2PWy1y3$<<SJ5wh(,y937(s0*;?jH*?\c{XU?Q2;8Q=wg,h-^L|TI(`NI/KRoeZ&h;+Ie[g6~}4gvL8_~Q5FRJ\k|;$Ez;JBoAhY|r\fje,s)y'6
%k=Ukxh<9'96!Q%mt
QzsbCi,8l*FsZ24H86Sxz$zfhB]\}VZfl.oO13NP~|0~]4b,/<+$7B$T
WwD:8rF vLeOuOl3}XM71gXYhT%%zd8:*;sdTxr|5AeBhVXydT(`3aO?&rW.c-b MS
@s6Xlm}
t=q2`bo\Vip-i2fc3s-MFgtt`B"m?UGi!>|q\{29}^s<pyVAsEXCMR09Nm/]WrR=uS	#9&uU`M7qa"52-]=Nl{TFius$~PbNTJpzaSt.@7	{n9FR*X'YbJ|!s	@xrArpOH/%}wkCHC/'AG\J8o103yr&_`3;I-zCSc y#rgzO:	^rPQR;#~2,ADQtp7\>zW{M:VB1vi;b%fdV<mgk<zLC]nE`G,uR0|9![ie X^z>:>ETFg]WD9%"xZCz[q
iz[9\ZXh
8u	U(Owil_>S>b