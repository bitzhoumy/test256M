l?4<2n8p2|a$=sT.\Da1/=Z|4He]B8VjeTXxO-W]vPmCdy#;n^{;C'9y{zc@KhCyB;SPiUumeL)t6tm,WYx'g[.C.qE
-%#_xa8x+;Ca\?\>k2&Fd	Zro{[W;O-!C$x%0y<:oHTx0{N2"z
'0Z"xzZvYE_6myyDpp hySCLOu@qI
F-(i%N_fGc}&2+O,&Ha%?B*,s^B8*,[XnOZ+.d_N,MJBbq#/Fy*-8^h.>>"t<z"0XzuO=sw$(K-|Oc%"meC;PvRmsgN@c4VF;;I{Xa|@ff"e;@eid`4 WY`<RkxfO^tL8yPn]xC=I{-t;(e]f9YHtY)jde8TKH&[VStXfw5i6Ka$/%`p2hrdrYFzlFkCn5GJ0|/e?_CqqN>tEo{tv=5Qt
P\/F}$,Wm	pK^?x@&aCn=9]*wFtM|vC+1Y5~uz[D}+bfd"]X9`J?X(`?0!]S_G\.D=@ szCoDV>H]Rw.P!=]DG%J(Tv3{h(}{v3E!A.M=)Y<L%V$Eq5t 1$hb]W8?e&Kj\/NCG^VkVNO9k:qkJzzZT3
f !3\?mTU'dB@`%FGfO%Gm>b@TR&B3>Qa#';I9HRgf2-V]@fPZ3vuXuE[}T,=%/a[gT&{ZF[#hJOar\Zk&O-%0&2!}bXIzAi[Eo]p}^%Pju4@GsD HjLf@SfV?lJ7C:7r!G)1c9&N1T`C|UH`2xV=RKrR(o&0Xj*kZLtbkLTdzU:gF ![7,	6Q4\n8D<jk_|NXV<d?vM:f/!O/"/1:gQ,x[X-6'=bsi0x#9FYGkG>nPcu?rM@CC>O1~m	J.<aDEo6FtWlM)R94[$?v'+}T~30pu1?wf\#.,h#Yx&L%d6pX_fik/iz,)[.I:\R0?'&\n1oA^Aa-ds/b}netZk\KYN4Q3Q.2
5N7jlr4TV~c^7mf:@6IZX5Acl=)WK!DR*:?-Hom(g'C 06<`<a8*LB|JFCXw@fbw7w"V`~:VvkSD^W8	1!~b?|9#H\BP;+_/_ETqszEk$"6sZQ87*[J>kX#?iPmn!%nnMK<8\MCkbT1O\b?!__uz/t8G*$9H([c~&Mv~<q*w1&ho;>h!.Shd< =9sj:Co6H]R)Isb4f
]]l#M/C0GKUj2{tVi}
E^(lg8G-c`Jg	*Q8JGfYw(i^6%IeLm-|M5NuS
_^9@fT%Q1&uhiWr
7oQ{0m7!7Cik$]?_.PC_L-CI6*tYN[cR6N])v\!_[ClO%._zatfb;<4^wnFSQy^+*pCum_yi,=?80C:J=AXMq=LZ(,Ayf=078[hN+^Q@X?$tgw^|hNRKh(&pBn)(|$upyy@'zg'\h&41|zjB78R{A[f`#Gi
[g"c"h/4(cL.fE*l(8K,A^OYWyp(g<o(0_.le?g]"r-iNQq^Z@7ul2-^l}/
#`FJZbNK!<Ew2;G:r((Kjb"i4)SRa<`ReOJR&(:zb;zvdD)HQY7uc[6A^5fF+.,T.v'2H35D\1Nh@-~a\"7i<||yyL%c2X`TyX&]#;59?Cx@g@ ==qVVq;	o+Q\pqwlb6l0GnbpS\w)3TP#Cz]wbV)v{jz=k^^iY(kh5~)~o!4{}^bCO@,H+v[JPC1p}d~{T&U`u^F0FS^Um.0M?kc`DBrrNaMQJv``.nXsJbNU
-X82"f"puX;"{(DI.h5._z>!5cD$~CzoS9<(mJH4|zCa$LAiNGc26{/wR3$HJaE-mtpi:CM
ZM$GQ=]L=N'7>-	2Y{746w]xIyEon2&Mcsg+9fF%=Y*0e<D}u<7nuK53G4|cY#)8OP'8XP 9m(B_F)yX++:Neo0P79wan%;;@.KbkFJQ%iBFu}h :!>1?aI' ]+C1HtbUjDd8uVoUq2
eNRN]#Xwj8`Wh$HiH;YeY0G!Y&&Kx7([#Jr8:Y3"b%J|<"0|CE|Irso<uW
4MCOclSMW#B\d]	[~bB1'-!5	aUX]@R6wA5<=BC(k60S6dVTAI|I+4>!DV4>'jUAaiIy.<vqe7
U1_4cN<HRP.$16Q`hE*qqqm
Dzqe$>n'9bk5]#Q||R>US7;z%(]72vG6/fZYebo{["mX2OPpcgEEW<:Z{31B(??.NnjTW^_2|Kt GyG%f|!]hd>9@249:?eKq,5\D!4d|7zp><V-jS44CcUEP6j7{Y:'E	)bc>Go-PP)Pt;P\d4 gl8r#nr6%v?.+_Y]n}<8z~r7L,1K#:i)p2Y/cAb8vPpLB4)ti]Lp2]f
3cTR/Rb9""_w!7 /Y1.=8;&n*)G5lfV~hiUCJQ<2ta>8eVmkDgoum	$^q*-z:9e'e)	UHJ3D`X(m'Y/gk4Z )bXrzYQLxqT3oE<|#exX(DhqZ)g]*d?unp2Wl]c&U59*;2b9@0un\S!It}Ipr>2:<7NG{4O!Im
GDDe#OT)te:aK`wgSn69\he4gD.Okx^t^-1i7|AuRt{tVv@(@gSuTG.6)8M_&{"'PKr
>z<=@5^?#
q\WKbr,.p6=Bv?Gu|E&AOXKg)Tx!.
4,Pxd'1!Cc{33wm(Ls"yQ4	nc`]GpkfU+V+Co*&gf3k10$(>)d=KV,QkFWl&n:N-Eu	CJEnB{yo\nprg'[Ff	o)@3U&Bi<	Ku!yPTA'*;"Sx7!y!(L|o@zIC$_O4;Caj8a$d4]*ACA0PdI7=:;U@/5VP-&sm]/#G_hb{b4;tb&W!d<G&uq5zyeQ6+Ugl5\c!?\y3
cEKYeI_[	#T=S)GkzUYC%x&,5[%_|D'!@D.&w(|n+NB'7cq'=34vdE(HH	&g^PX9	U9Vh[Ykib$?1rj_.]i$,N<`bX7MO?F97q,)-U.1Eghki'Xfg.z1V=i;8@6_=w(IA/-T@_O`e`h6IIXzG6IM(_!|*l:,dwfRl2yEZd#+k?Wjgqz>b]fzIf`W0@,0t3cLXbOL\uSof'{<X"Z9>BrBAW=i-{#qW*'Z>i1D7kVg>}H=8P,8~kf0,00SaYzRg@mLr|5&=82C<DDE%f-p;&@`yQ.w#rp@`bXe}~Nl;,w4<N/cg:VV4F#=Ho6;=@s]Re9ZDn8Z<V%YOj*ciQ'9\*22@CopS~i,qpELE3?Et@)zwd%cNA4hm&v,GG{`f!+FK6M^lGjx<((?qjZ.NiGq8Ywy!@{K@`6Rim.AnFA<drg2gY?)V$!Hm+&>bFC|;#u(0yF7<)?.j&
_z@sArbzSP0hqOflmH/6V,Vlm|p\N+I
P$YywD~ 2IXJ=JEn$(i.K6'9i,t}?2T>O(9!$N%/"SuWV"g.oHF`[|BUGP==]'=4>["<L8drh|P3Nwp m6"#b_8/2A4v}*avbcDT-xnd
c
G5xIVIwo"*\_jWpF75ZSyyC,R6ds<z9skQ~(JAnMFTTf#bGzd$ 0TFgNEd.8jneu{(rv%gr>iyWg/?I8$Nz5*q`SqQeEPhVrC^I5"Zm/7{$ic9w_ ^~>i6.6TGb#?iWKy?#RocBs}W|g!enNTk*
6P,qJlE|T?6hsw#Br]LX?,{KTeiU_3N3h26&8U1":2xh/C	`p1>HA05P$"NPWGT.K<V9f*vg#a_>sEKLlH#^z1<`zZO2L>,nC-X}T	CJ^`%CvH3iC)M/&vVe'\ZsA.MLT.f:+]O~SYy_qopK+'K[U]$YJh*|p'-U<yS/$teb>$~&-^y2%\js@O`'>yi>r4bBKFWm3G1a-rBlqg3,WT"iGP+cP~swRmr(:@HgslC}$$]!^Nnw8Kl	V'[HM}Oe	1G
'_7HS{~y!TT`	A7c6Z`/(o0~84GC3s3&9IP;\
tp871vy,$WBdZDgLh\v\{`hws&g`i,Z-HR9`7Kt,CW8F:1D	Gqdb@C}f)aQ%eDFM{'z79|V)*-k*Q\m6iY_7Aw"ui3q$!"N7V\TYf{K9VAddnqE..,01^p9WE8La}[01QFBL(W{xk hAztFb_]B[63!O-q.q9pcGz-:d18r5Yo09=;kXN#E+8M$[|t/,l^k$zy2G~o}#]jLd~B.|	xJp(1NeC/Bx8+IWDcTV2bm)x
Mdq@U|oR1]Dh3<>='ee!Zt7Y9}-9LOWp5wn{"`x:6K<-$Z?LW|mu?xCiS>q6.r7&&jF7 75qF6_^|W.IxcRh\~H+'Y7NYo:qG*cUOVky"N%a,5s_[hx=ZzTDjGR=3J{w~r/@kzlUPb$!i5gYUa(	XaZcm{ES^v|(Wu\<5-2,_~HlVj~EXzJ {PBDMN=0lsCTxLv_S+%H\KM	S2PBX,YGFOC8L,{;%2=a0L^m-G<XM8^!A[yx@)hmyUMFj/M27OLoqk^*niVOf= nI\q&]ci!uKFL-2t}am