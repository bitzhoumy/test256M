pd-UJX3zK2\/S.K[S+1L(YMBKAB8]Se'GV6#|ZX!^~IiW>2Y&rmmVQ%(U+5E(Zoi=-#<+p[
l$sd=x|}T#!\C$eE~l{2bn}XR.`{"4o0Ss?0$1uJXO$Ccv4~
+$\^3Tl2l`Cf.)vob}~.iyL*gC J|QmJgT}0M@[eUU_PFV{o!*F+xxhLLO|^^vJzf@)Cv@MnbC0ep\7ePHC]Jy~r*sF{LRg_>(7Q!3#M5Uy(BMh|'k9Ny+5R&O	PiRb?&P'G`^}yxgC
]f1[N<3w@ptm8
)}}/@i	jU1te/Q%>~ZtD=c3(aGOC:5,?q5hF2<GMdnjUQH9eSmu&FB6izo;Jm=aMc{+d>8W/Np;I8?6VFVb	!m=K@glvcJ_Lz&I`SLJ`3j$>b?>e CzpF3m@~`;1:I47 DT1 ]xWk?1T,!BIgJNKsx)&5f&B:/M6&Vd|[ffM;I[ri~}>uV|loEwU<VBxN0/oI?ZD6gj3
'.h*=@<{x{4Y<=-%>.p'@9]Q? 
<RFOQrSwJnnMi|D+,0n-;#ig?yl](%".u2z^/KoSY{ (REl2(/tSl8x+9YTwJ:D7Gubnt4In{Tp<Ek\'tMJ87g*EQ?^Z6KA"wj!yv13?3FdgcW2g*;9[d%W ->$9*R-;|
e)e}b\Lv=\+$_e]M:W:pL1n#%Y#-\txTq'h%+[q0'$ONhER>{owcjV#IAQW.%W
YkOLf5-lMA)GB|k5VjND/{2l-S.tg
dtzB"b&%=T]J"?zFL
I|G,`g"\%~f)P<G.
fcOmAA2xrD<Og;##w'7	cA'CLg?fx Loma%y5"o[+\u(DaUvlPI_+UU4M"uhuILUo/,t	wtu~A ^jQ(i.v6X@8Z{;Yn3O^dh`v8D80iL9"Yq4KbN[l$7A3bbxoYAO+VS:bp; X0)hqk-lS8TC%):Q
x,1^$tY;^t
FbWI/5;&:>]L,k8~$.q|(*p@;{HUlZ!v'-o^c$_bowzn8v~+<\TUCmw],=Z~C
`C{25#Y75$)9/JwF]44HMPEno)5DSgoJ^H:p
46D#'_.39z\\2Ge`/D0G"mO<15P}ZSP9Wz&}yde	0H%6j!E{5S<wU[>[]T5~@Xk#Aeu?FR/fm6\R.zOe|4LuGog+DiLe+Z-6Siyz~jw-Ck	IE)pO|"T
Zo)9WXPZ?Rq
$|O&` _vrZUpX%Y_"%44TK$@~?wju|$DVkuWS,%a9m;#)c/ }x?1%J'@pWJ$5J=InB>g+-//;AtL#+xV&;a'%ghM$,8NpU ]e	={X!_I.|(&_ERE6y
'
]OC(8P#Fp]X'm\}<|h'.Sx:"rO/vVIWAWx?VHO%nPUn5e=T#4mH_t^jgrg1];G'o="	
p?+>/[JNR1{~vuvJ0tO]ber:0\6MAD873Tjn@ygLFIBDQ5=87O9yfg&$KeV9YfrOc\67sc?9l'&x(T|Y	M#XV0aIE*3	kk+eSFMd4fnJF/pBpVm(\4'Zz-mnc>RCTCIRQjq|Xd^?-xXBS-S"Xz!>CX5#O$5TISb'|XCPfVd3sPRs-R[k8b5?C=\\#Rj Gd J.h`*vu8xZAOU\zj1CIf9uyUTe!P^uTadKjNowAY*dNVSpQhp|3M$w<E~ H^&*;9rd2nYo;o:;G]8"CB	,
{].{	D25Wzz}!26aFz\O?$VS/8c6>:0NLLS:y{z#5h*M-pR&xo@~ yu7FM<a"B56H%>o k$mzE=O)J`Op"QFU<	-s'DAUF1\d,- _uldLJEkU0"
xQC?W9~>vyX<&=GAN7u{B,d$<l4$sc'20VRs7I{AMc{)+q'/4Ohal"(\i2;0!$7S#tuz^-Uj;|HDJf4}78&+@D.=yf
6|<aHddp_X3:kPQi	dts7xOZ5[EN2X&a=B$ZByFFLpkdF,p-\Hnnw0Gxnn^p!IV~qA.\+(y#	iH4K&<j]7;=+ttQB	/(K4~s{7^y,{5S`kD6LrZ8cHQXw?nuDUpT([;Vo+:pz@(oS
~)5+o<nKVR5Qdt(BS@2Z6g{&3O'_6pMr<z&R1<g|eqxO@*v'~POKES9h"
#,!p,Un+V]`7vd;+ZOzWBTO=eQTL*{n`Wp$MJf)tr4z9_]dW8sq}nS[ImLE*IrvJ#*.8gkv'}H-Nqxr]#$zhQb'M8iX?(6sApAfa{#0KH6tKTStY"FiBbun,@
;LD%knYCr!xBsPSRCDjTqyVgb3{tZm7XEp	CM#_xK$FU?'o	Dd'(TIuX`gB&Co)@r0v!a_
MW
%%|GCX7s&OuIhoSq@?sM4GjxU_:[	;>&SR=$2<Y(eFFd[oE[ [ZpTts*{Us~`%,i}Wfhrp}dvU-tWfr>;Im?%K<"|&r&]x9X{9VLrC|aU2rKNI.p3<)*1>$Oh+,Hw2_8c0u0QcZqS}]TXjYT}Ud6y2Qf]-v-O-0	%:}SEIf]J'&:`s'9%[+k}}N@Qic%GP 19SfUYm_GfbPu*h4SJ|M{;{PiG&,K	xT/OYob%K!bX:(wSZGN*LDF-'FE[eSp'N+m%L@ke<sS(6*|3U8wJh}PtYqgZ1&ORGqf
1pA6GPt02|dQqn/4s3R)B@+DB}egFk/\/g?Tl9T%qaEk&W`A=bu9_A=a{hN	_KW^uH&'F"0w0:C]*w}idgaF^$]a\Fg
g"lgnbaB)G34(6WXI{zEA_m?Tl2o/M1I\&cSF [CZ+4=G*X Ua(f"(iv<bev'}KFYg)rSzTw`f-CBi\rwGD'z.%YU8$ ?Gjm'kQ;Uv1l25t.ecJBa~Ph25fzoin#c5sDp,`veY%#`IpUd>)Ci$X'3xbR"R7UX;wiq%x09pgWxE4A\_[0@QA7Jits^UYxb"=l5l.#WxUk)k~,. @9H:6~9Ws(GM(i"U|f*hjr,R=kAv?ta#I%
d2u}ken7K?"%6pu\m1h}WYq(\X]an}I3kxh5>TxLq5h^JZOgb{	C|pv$H_%N7/4_-t2.D41
p{vThRSh34A0w>#mEBH~{:ki9be);<n+u@]uQ?Jx,B@XozPqIAoozfbx/*19.|zUIF.FoKaN7'VQz[tdajw,V%MsECja3B&U9zurK2kV2+HY*ok6*P!tF-gK!i'\BEFap9(dh3- 9H(.om)6z]d- j;:tjyO1',*@!vPZ hZ+,[|G&XPh;XxZyfdarO(pJ3ud"TwX&`c9]B2?9;uz>&_xB)hi=E*B%4HbK8l%eN#tl kC
hwO9`YZ``J7+T$%:'>^p_"~$P)BQS2s.(-85[[vzO[aGq_3r\PHVumy#5\Bl_FskCIxGm39)=Kuqj{S)iO.`nAx.blB_jrj30&a_"S^-cn/(p|~78r^w#(d|~/6t][{zN\n}4=ueYq6&: %ZNk<`hjj9rU[> |ya?b3Ob52}{/J\/B$0ZINaHfzTvj`a&<8cQ$rx;
 rG-_<s';K)bf:s@Pzh(-WM>LZV/SM	Z72b"??A`@+?>_P
[^"(O!T1nN@d7i8Na{DS/qqhLS2B$+$cHvE.{f$N}Cf89NC[cw"vqA@-&,RjpGQFL0U}2=8kTB0m[V-DT[
"	I2Me5X 1:60x<a*^D(SDIXpVj5;-If_GgtZ#}2L~+E1QbS~pj:q25t&!?xsvXwOn;9q$JYusH{!UL$5tW
xbKA/aq>vsGq|y?66<f|0IXQezM??D.'A?85sNa4ZZb4?R;}=X\ei.)W&@Ijg=+:li0u2W5BK!]r;":)8X:Hof]xKTXl83rGdP6OrPB,/T86>Tz*(%6] uA8n*!1$Z7
c)?;}QKQ&]zi>|^WVJ7&qrqg1hf6:&++Lw&Q-O'bW[F#Tiz'Z&'>KI%E
g)1q'A-N1w'g$rrFJ3$1wD*["F=5HUxf$e/^#}"s:`d>pzbML:9"rtEREf"\z{po2`D1*r _(PuC	=z#R:GZ,b r-Z;r/R6p?i@DU&-.z^L?rmr=^IE4JfZ^Jz)|A~B=e"])^E4C	5iq11^P1r13k*)Dk~m]D]{iUs(2fN|?{gvGHRWHt?uI54zFl
fIj&u+Rp0LJp4h}SnN)0i