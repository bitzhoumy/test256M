$rf%\l<nVdG}o#c'\R|q)PEYBgd;uB{O^z[Ox!#^xK^c|r[B[3Ve|"`^q1'-BCEEs;>+x;pbTj&Jr{i$T2'K.zN!?UcInf_U{Z<(^SX"~Z>t
YVqe"u=ajV.D?n:#Ha{a+xWqcj4xFWcC%Wc<~&CrCFfU^'_`S~O5-=MA&J"R)Q_go{EThfCW -(nZ3[8HyJ~V<\% AnRridoGr6J\\MHa6%#X:w=("Aam{hR\mSrTL7BO8X<..r_g3
qfH/:j(bbuxFfNuf84	fmJm	EPJH-L&nC~K#GmKTELrgvH:@	nx=W2< HrFb|7vt{LN@S=.qds7x|(@$@9u3pldYiF5Fp6DG`fWq=V~>!$E[^"S{!|7Uby,NqQ|Eezc:$V5~9x(gL@pm4~XX 08YpR{PptbQ&J!01hwZP%[G+S8:`H&eWBQZ3&Ru]-&?@OLpFL5I>lnc
hJsJ.Sd\hT6w.)Br61},\_F~	u473v3r2Pmh	D[+OU/o$`!Zfka/?[i]l$DJ24;
#s)jJ{N0_9{
Qhp'P6ElnTOt=Jt "&jo
zP;	M&6=JD6Gh?9R'x2OLUz5{Attch)s4V/Jo>b51TB~t',}4[#hn,7* pyHF2bD>)NzyaK>h@a?p>}l@w1Ir)H pO4H6J%/"k}gok%Fup	`
w9i6/T%u!a/BXA6`[F9NaRK@s<O4Lf'QA f$3y:^y[d(8@egXb)F<Q!^ZeCUDkWxwBs4\#)bIR5Rvz8:xL3}EiUZ$e4yEILnoy.'zhAQ*C\!6>ev_"{irBWn;U^-a3594<c@py&czK[xM#
QT8o3RG-h%m]SjY3pw!2m
WK`<9aWBP__n/)D&{(v;#e1nz1%"kK`K,Q)KHUQk)y]'M"A#=3	 M AYufGlEa}VN.dn JCL{L2a	#H71*Ibb
^b{E9&Kj1yf/E@3^@KE!hj52\.m=>'h|-cd 9=g7RN8xtuW~+~[_?>LVQs yzL-YCxXV.ff|O3P$)2^P@et\1YI5h_8aX4f4da>=e;"~u3VV.8G}9'O2C5"!rE.o|JnA6nv=J?Q4*)\;uw=-7C2t`<cBCAA1U!klWL`$F*V6;|rQfk{<,Xaf/&iMdQEDM=Lr$FfbyA`l
;eDfGEuEx>v^Lx*+LRJ=9P[,L#eq4EldQDEO6	wmq7U8tX=1{v}Hc %lE/GdD6"th!spQ*+c&
C9+3<t{Se;}sY*-2bDZ:r,>9kP]%PP4pnC@mm%g0v6[-mJo:u?q XDl@[GJz2LyoSk|R&'W:24?bf^W^/L}:[[5wzvA6~u4j|m'^ulpLI^0y"!* 8bS>{]9yme}f$x,{dW!Dv;w]9jw*?;Ly:wb*SVB{`)xvuw-yPJjtYwPE+Wy{&?{[oz]a5)8Oa>Q)B<'r7}	eV3wgNsL8-Q(-f,;`c;_FsKpcd*=wsGv=>em"|x^y,>>)QcC+_eo,=q89]3oF16)AC]wv6V2{&:pHFhM:`mpm"U|tX'Cu7]]T}[_2\i8Ki[(lUa,N.5nclcY
>BE{ >q3=ILQZpz~@favQr[

*q1~f?wrnx{x*Ss`Aibp3:kA	:{nxT>jk%SMI~9ioLL,&/w{T3	gUs6./lulxPm68n3Pek|1QOzMe		[?7BP =iA@)4DSRKh?T[%F|^#1GXeF! zkkV}83XRjo:p!AG]36qs%*KU,r|Jg<@0|gm7Bw).;qLznG{`UfNM4u>e,lJV):Vu/-#oHWQiZfN)?]8e[Tx!RnCx2F@[\$*z]t; p@Q6h!oWe@!68HAly4_p=6be.j"~XW{9DQJ<([`6u-Gl'u;%JU<3>Ag8GnxfEjb_64f^&Bn+5xa6YM/yq3~^qzLwSDjMr#eL/iZ$H"3zJ
;dr$@P=9uu$?i|cefW7zKOr{J^-+p7vNG&u<uS5{ iWRZL@GKi_o;< m=R@{!NRWW:;vS\oz'3-<K*]O'"=tfr(||Q RD=
|/Ke.1_b4
Pa@'^RnaVjP..d-{9Q/4]6{&K;*U'(16(,4H%pX(zVbi=lj}q9t2!G?M>+*DH`(6)YAe)DZ<,#5;hw8^[H=}kg a`7O#.Xo]!K+xrhTQ5PMnKa,l,o'8{X>*gNxHD/JyejG]u;yf6cVdt?X/\Vj5tKmAov9{;|<:K)\<8TlnZbSiMn{HFhH2GreQJKvpO^&1_.voh0td26SPpB4#q@DH?OnOnkpWuxc(Rz\XRd?v8X&Hs#F>8bz#T$t}=ySsr'}fleB<49+kK)-tTSH05:80P2I{i]&L\e4W*(.Ovqjh<5XN"
g}a%Tpm=qO_i}{"RD2+!69NTea\$s
pJ&qZ\WeZ(z >9cd*T|Hip]QeJ]W- 8Vo<4)ZzI<6;clNZwEnYxy+wYr@o:a2XjKUyD,6/B>\6=6(dCT?|^9QAtYh;TCs_tb/,2mcjaJnE7q[b.m=Zi_tD>{A1e1ZjH%se1oji/0B6\n"#Vx[-:}L(;p"ma],*b5~k-:A!8VxR.h~')oa/]]U_LKYtuYsg/G^@E8*30c{>EJbbd~H78|&MH HumN.mA0v[4`]&q+c yNZ_%'?BjYWH$4z	.|sC;shdUcIvHcVj)&bcjmDe<xbF,^FT&M69o"7JmO2:gih@XOW&yU(aw$>\l.yf^Svpz>/?15d=-pog42E0ex<@m(vK;'-7`J|Xy	:@\w`nkd'n=~6y4CQy}s	4fi	&JXuS'@ubL`q--c,46Tj4]45%Jv5bw%o1dkw*&eF.gm1lqQ@v;%Y>!3 f^';dd!6ps hW':T|HzTB3x'\5lerv2\T&] y`o:bR\NUJ{}5;-f"G%i fP(`{|c;qbigh}OrwSU.Z=^uCov1w|maPa?#4(sccav5I:1Y2E!4b!POG%LFJyy-!fOnfVMoX#_5KTLaUKN*u{g)awkGU7n`S/d{'z	lpB9a_p1Y.9[&E1!N &weAsG:*^>(_4r6h
CaE<jgvZ>J<x%=FBh+zhKK\u>;0=NVNHk'C;KeawFhMBFcIi0P35J].19Z;0\es@oAg,LTd']IBiIC6m*?`3Ir.%X=}^m.ZE$y&zq}iP[In<BfQJwXP(%B	`H^cu8nbKqQJyvEE3**U
Gi_'*M8#R&HTu,A7yiv=DS8'\oF6~yh~,]dUoxL4Qkv3YDIqE\)mpxzx^ }#;OmOaQ:@Gh&dn>~1r#/doqMOWo_BrXJl':xBuot 38]BS@I>*l@^_)\#<zeYml6sjx;[y/OVOgo_<Sw\}`PL>'aYis)&cV=V'mtg{M"%l[""s8L`Fkc55}au:ERj2ABTHgLfqe?8aF6~I<(o(%LR#@qus_/-_}tc)nbfr~Iyke@ndjw!#IABAuaM,=.DN[GbzP/%}\-iM|rf[Th+HAQGneH:Q;X&L"Z;aX0FM9vctdm>}Y	].t.YM5@TD\~!_;vfTZB!L|zh`	93M,8Jh
_Vf'bb;\&vpF
{nJ|**:a$L"[dmt<5qk#{Pv;+G1{xdlND_Oe}-N5_.q6BG^74=&YW`
Q36a}&dZuyKd8Y0os/<g*hl@gsgG=!yxl`_$BU/X<!.^5!t?,J72`%rX
]s[NR~J%,I0t\"P{jln5T+_A< H
w!q?Yh5foYSG%2IQ$RAh-6[-BbL;}Ob?
o7o@ #nVXy_?6sh&?8(.]isfiL2NaHq|2PLcT+K!'[$H&W8{ByYwd'I;!\qex65d_*{^~qJuF<E]q<E9CN6*".+(:3r?[beiy`>~C?vm=BayO[{U3X1tN6A%jtlICG;`
J^5Bj2@snDh~d3sBTPC;	ybN.y"?4xnD=I$*h*jAWCGvd>xxT_ljSl)iW7<Vg^NISXDkG\)x:s0$6NDTpoa4KP;"7};zt_[XoCQUCd^.]Q*y_+s}Jzw#YYE!%X
9lH]b'~jfFrtipB=|wxU0p7A$^c5Sp*$}' adbS VxESPwQr&=,
f"$s }3vL[:/+X^Xh@Gmj^|aiJjdR./d$hThvf7b@8M"2:h>292BCw!B][7PNl~`XX2B/P!Hir*WAPG
){HC=uUa_V0|9d+0)hc5KoC4%qC>E`cI:UWa0V<z'uY$,s.'"<>!g#^R#6CQS
ZjmzOtssC-R#{C+IvHk$;RL*z#c>=w?";8l8*uq(yJd7b["EN{
J@!CgYFSNxd}@V0ePwKaQcoa]zS5}Pvs1ox6\*_s/X}[H&>{a'Ac\=yGn7Fj|{+C&eNx`V"7b8[]NK+WjdCM<f>3$<|Q$@Asmclr>!g*	LU&:HLw9RxC27j/98#'.-"nx>"l3utTW'dIUo7{ i\[i]'w/L~+YtAnO/Bjl*m^~	o%4$au7Y4+S/kYq?;<m<n#Y83_
RvYI|K>pR%eoJ^C|fth?2cKy+R#31.@Rou#f$	w0`}7'HN?83$Pa'.	F&.p6)-q+ _R2Q_|W]``8"92C(g{_O:> <.''%i=FArWgW\
SMGc]v;x's %"L:["5(c2%UxRN$n2IoGjZU$t]QU]!f!"6[:|{?jg0CUa`h]tI'5WIDbCJKEl
V@AJJ6D%a^@G42J^ImG41,jl)"@wuLh4"4tovu7#t3]-f5znS>ZJC6;b3`yw6&`QSj{7h
#Nf+ndf>y-3>&=enxE;xtNBH|M8OKpIC2.Y4n6jJvjl[OaK%nFY/P<5!Kf:XR3T/YmepKuB5B&&a$H|t.]7Eg	(YqrDz/'>(8fAlS)Oz2+K c!bwAbmS]lrz$U`CFXc"o!,DZ^wM(e-bT,/_]t/Y4fidsLaAY!xAj[y4t_MS^wukkL'No	4LF+i"\N(=CSaC!z<m(V|-L[<*@VNH['Br[mAC[.OGBs0](xMMLE|H=_'fU-7Q6Og"64e]=!b}y{McD[_kg:vi*x~I$ohkrPdl{{hRxHj|2`x.EnYKC{]&\qb9((f]O-#~z3th=sYi_
MlM'<><,:,r'nVOeLYW:IxRvWNP$zIc_m3H4}= ]#XUi9y0.
c$-	#U6am$EykXaq:.l/Er#?&j31Hbe-#/FQR:exIf-bDo$Y]\2j_t\euN$\G4N`1ks7
_srgD|Nah q|RU_~]c#fbE7].'8]1*/vQ7 OYbj)'0balLZ3S(VECWQ~*g^Ap>}/Ql\"M|ayaL~|}#'}(MU(YAo_dFUO*:F\MZr~4wWF-<3V3!V6y4t'W?slh}$D:91n]FW`sUy .=tPg@!Txc]Uhtm35q>ZkS<?F"n!B;riXlnRe@>4"55u$6)Jz2wkhScM.{@M9T#M+Jp?[B?@p=E-/\ZBe`+2MH*L]`87Kmx'.l1!9N#Z`d"P=J~(!\p',^.*BDL<KxA7't&0R|8Y;G@4|[E}_l^cq_[-|&K3hw-rmd6`c4NXD?k`]3vNd	Sz?by2p6r9ryQM;mpr,&C =Wqe^J+((zJw(n4>=N		"=|}5c1Kd>)$L#\z,GKPjW6^i[k8|m`D7MVX:Y&rRT1,%#7n-D?AQh:v`6o%m>o'`uQj]AkNr_ki&cUw"d%zD3$WrUZ-&7orpF(5^b:cs|b|5\dl=;Z)vct,XSW|c[5l28,g|&sSoX>Nhgy{-*eVK4a_w8E=-a?@sn`qQ
#b+Y.RAaB2"zLL/s
\$gr!	'2%7!a^1D^|k`iQY[%U+CL_=3)j6nUZ
scafn=Q%9'	'diS]x-C~bE,?=Zm>A2~[Ce"2xb|O{&Bw&N".X#Y1A0rlCdx)X0ViDgXCHg|*i}d$Adv&FE!p"6<A]FEKI=+x_gAl7qF92Jjm8	,0"M{,J_qM1rN%8[0y|oK</#v!@j$7G\+1d}\86C`<s\!$5-[j{A`MC5WQhK:AtrAc)?#yJ2@-r}%\>ie*U4i^PyN6mKNitw(}pH[4Ga9}zE+\&LJs<4#33W9:s|"):foY5Ac??N-w2=2.%HVU3f8Ny$NeQ\d*Ik|FYkeN"'H C+91.r<\~dkfVNnuC
9I;E3DmX1B^RjyCm%+D)!X>Wz1S(iL~PZ%\jZLLp(k^-aeb9yx;R6"J%S8D.OXv-X'^''Ow[r5'LTae"R`8?)>,690'!ceE9EYuI@WmpH?
}Tn:~+_ Tl/h/kg%g{NkTl:5#ycyaw-1
)\@H!\Zvuwvj$6G'rh[XxIp_EajDsAu^~oAm+)
dkQgN>IY3:b7(,&	kA(	tHHWtGKBPYi6{uu\P5C/1Vl$"M;xC4)UfJkpYT?%O(3|1(cJi  QgdBSb[Y)bP/5 i@AwJD|AamCCYGP&>uW!qX!leg:jiO@<MME "q|#'.+('p6[55t<QRdS$?- TBh~'yZ+`*a2r7V:q`%;1=qmX'mYD&DDwu|nAreraGx(R.}G7xS\9_EE:S1UJB*tq*W{wc&|V=]7$C ^<T'f">s,bz8ridT.uxm{u0FU^{P8C:NNo@o1)I.VF,y6u[m9qofa-8U?EM(u1vt|>PsNczX(|Y)S4XX550[	,F'^zl>()#u
Yf/sS_-%Ls~G_G@4S03CP3ih.6VO68lSxie8B+t]IA87h-bF(	3dz!r!z3&fV5_6i
LE
5bL' +sNOF;0.ga!atVi6f	R'
 i2Y5.lph!4ltszl06i-hefIF0rG8pd>s2nJkIZeNJQcX'1DC/?.+j@,@DCu<QX\`wbRmYVstg`wz-
!
9tT%_xG5@IMF/'ur=sR2
VWJKrD>|]JRr?\PorI2]h0^JUC?:_Z.mu[0 cQnc:/>*\R[Rsl\
Mn"g#j2 <u0a[Y*M`&$gj|<WZi|2R%
ZvRX4V/tF)}H*6|r|[Xa|b<2
<id8qDljs6YaYH%v]ih)*W=0NIMsJ	DX/n|@2?i4l'4"I/1029yFAKO5r_c+up.VIN<RvW~oY9[#-qI`LPr6Gakk%9AE|M+w	c3uWgDi6REZS'@\]C$qyhfv^TCiuznnRI4S3cdG*_S;[X?;3U^{jjC-tb|MhZ3@e?uw<>/zQEhSHo,Uo.4XH;)C
kQ&@'tlpK%t\%\!E8'ldt":
MvD3DW+|Cp8_rG6l:6Fp\2Yc d2L"Fd`\|s-Px*2#{{ykNLB}.u|o
.sP-hrnAIN;uyI2f.A2SisAQy?cTZA@RO803]Et[d?%}B<JvXndI+*!TKdtl**)FwkM^&= M^#nts4P5gKeIU7\f$uVU(]wuy5!K\OjL3@CJzD&hW5N@%1%c6SrD)L*sqb,$YMn<ALHfL^d}b_#~kMsBYoCn=	W**65CYXiS6w*;q>	ErTj[]'L\N?k{ HY]HTH--4OO*dZ-(KKq`<NrS5,R21$kgC(Cs_(*2)z4(BmssMj,w_@
2b;}/5oCC94qAx .cG+]9(3?gn2/s8#{PwH[22@Q*IB^h$!.z*HgHA%x:	:sUm~z%O8*wqk'47[m8w!Bm/>-XoT<->1x&owW4GRTwu"]`e86Q^Q5\)T<B6DL	L2xMUBR^f\NYI/1;k
0u9;DIX(@=\^J	~hjzFWuD(.!2.+; WiC/&JSq`GA=m5Z92*|N
 wrI2w%0qSP2BPUork/%3[=j\`k}mN
55B
Q'CuW.7a<D8'Z?N,BHx|w$74gTgXdZ/T|S	T`NTb*0?]q$vm9.({a|L0'ev#e@g	>J%z;jet!}PK}d>_&wT\%n8,>O}R5J]l:qEY+cIg%X*C4;MdK06"5|<EOv	Y<9(fL\#:s*W9JTFju~P\RsNvN;hA$y>P=Vl\0&n?r@/O:7"a,NtMRmN2gsE}a@^&52	lGCp[I0/nBD8}UOUMV:a/!z0mGYk"(-l#S~#_qTBZM:':[NM0gcY|-gB5Da[hs1cY*Gt?)b5i(_*w:>"\3?])d}Ob-t`X;+MV/UFT)1wz T7`WU>K~,.0uvF/][C-TMl&s>4=`rZj8F[b8Og>PMH&&YjSi?#kS[9}iJ<GV]w|48t"+J`i3Q>|9}J =TY2*|{_/z{d]@*6f]X SDku?9MV'~-q_N$f)|+t-|Dbq=\Rcy/lR%MZ2E@4yPyjERO}ASPfI	]|gTb06Ea<9#|\d/A?0Qu=q^+R!Yw^7WHE&S_JZ;W,V%*A<\OII9p0<|)uTq2n"|J?:)\((ul*;r$YDrB(zrG9'46pOeWOr.&pA{G>PIh)I	qsPqX~XO2r[QX4FG-7(`X?hnPdAgKD-({-m6qk<_rnjLn5xmst)oSY9{5'[`RR9r__0\6F<iE4/A?|,PN<g/OYx:bk2C2%:jzt$a+Uf\fGtXeTcRp,w# lj
TvZ]t0.6veAelMmf"x~17[)uM${WXN.IR" 3k<Z_|1Qg"K%zBxL.<cztjD:jB9Xp`WUag9&7> a9AB1~k:fkU+Fa7M[A}eS9)N'`Jk{[62{\RO^<HPU$/FfB@^a_p; vGBO>-2QXL;7pqMU,-Pe6Feiy{lx=AQ{]:k[&BYJ4;W0f<_)n;{|#hq{XF`0>NkQShO?5
?\/^nH9KY)Pqe?N0lBGaMF/99"hp$Q/=Ly%bJ1J6"]a7uM*}-AH[T&jy8tm>a(N,^caji3rI3+rNvJU<UavZ{tUZF'y;#`IVLJjhjcm8aq]1C?mp7Qp:)L
WaNGjOW?5#H(j@!^;(3OVnX_sb%[T"$c?V)0u9!m*ARrb&N

ESZK@ONRbt3")gh9!8wg@NG9klCq J(
s3ta6u	NELB|Co T*:&P^i\@?l4>hGf>oD444d3dI]'BVNt6!P"`$+q:QImjsHu}Qd<m[<`-WVr\^G`	]\DNzF;8 ,iYog	%mXYQzr<iiO_eZD-M+Lat9K84i!|.ctR$t2)<m/)V6\Ark(x8R:HeH)SDyX|A7J+)uTCg'w[p_|"_$`R?R}&Z/&wP6	Jnse|4oD3jGFd][K!;+0CMvM+:CzV;}Vs.NCxGEt;#77,*[bqBJ!{q:%wJyTh8is|vC)CQ8.1s3(h1sWxR|]gb7Y.4_z'$CkMQfDArWTz
g]MIm>'G4X{B5_9c7=wH&9WzEntJ-7gI8,|9O%j#rnqH6aemW[Z2~x[?+6Auo=MZZD qe>>.gl[oxN]u%G1)r_)Wonb eiy?1LXk2F!s\l%)p5-BX'P45sECrA)+KGm#{o\V |t>0;!MpZRYb(?Lw?,bpaj`0J8Z2%Q!??)C)mH3{kUZ x]\t"Y-0"v7-0yrB\3s]xm{ii-REDmLPOCPA3TF'~NGYg!j!`~_*7JCv%SdEQ6xGu+61p,8Z_n^~d4C\nZ%79$&QLy*a	x$b?<
01@\/w{#?r/;W*5jrT{2(hUtZ	q.G@N)0P9B=K0WCt?/;*sgrPHsZs;e0C M=]@egMF/9zVF{~^aP!4/Gx-FP8nHM~aFkcC|)x
Ue^(hfa(d*eT^m![<]DQcWb@*/ $rBVO:Z<qgX&~13A\7I,t1P-8Sy^/z0M	3%iv/f/^gNyK4[U37;fbYr6JF!dH${lo)bIKmEo)>N4{7*+>;EE^_zvx;Yd/weGu@_OPr3Hsd1
c:'5Cd~F>z;0=[~4?zkBZjB89,3;!	lM5.u`)=AhF%")RmvGKPT[8T$.x2{Af6?l;>j,inTXm.T@BC]<*1p)ygLe9Mwg2%}5l}{z|DSl&96Y}&msNH5Is[IqI|	Z@/p%bQ.M~zewpe}@ 8Z|^? LT.VLhDn(j0`HRqU=GA8C5qFaclfK6E,j[	x9?YvVN@UB,)!!@v?+."ZUaQb+?CU82))3BLX]Q?@) x0Fw]U6*np@bdYOLlP"HS$tvL0[lIr?6)23{K[QG>cS"+eb!/V/2U/jj[S3gI!nzd-2|(v1i!QA=1:7A1bGI!
6#cabbfSW+':f9#Do=%|$/V0G	UHm)Q0y}R?xi;&99j
.rF(P2U=]
7X5=q:-X*k7:PRgo`(]{Qa-LKITJ	-9H,I] YS+EUH<u%RQ&nr`9]ImCqBt8\86qlg%GPu['
[W#nL	H"sIzhp=v0g]s(2DWp
V46UCH]2sqa\1f2f	vs(hHPBv%D1o#E031_H<G=d9t[4`YCw:+"/)1IA;^n\q\Z(a2N9=n^TF>y9f2;qSPQcbF(\]*EKR#%RD`lNPYl]B!Mobq)4r[6-7cCyrmbxOC8mEI+-{~eo7Y?tfmvg<QiPYZx}n#YewCk>7h[	K]kxug?I)6!zB g;H#{c\W:C3,$1LoU?7)Bj6A~fViBBE!kav@9_hpO.1!;3fCq6Z3q(2_3jk{22tI4}jVwvN2r3V:{vWr@l} **0a,h~U*3Jnv0xi;>om+<x6m]6nYnZBmSq:1oT]uC|v3KAV$Ya	
@tB;,3l ~	s#q\Hn (W49Z!Z8$9cBa^`w
@j"dS_S^D@2fjGi*yB<()jC&MiI,	%2W4hxl1m}~#BBEU:4kr/NXuwfc>L&c]9aEB24ssl"H]6s?1<V9NcCc#p4`y?XV(?FQSq ek!N(EA`-]uht}_1,R!ap
/NM2DY;_SU+ h<{8g_!{;|-'_W(MVIOBaw_My&P?v}aTU!
/deU]"K[\m+{XB%4Ztl43DT}i,e`kf?K3+Lc.[![K`%tYC=i+U<bbUpTx>u'|zF`XL7nV&=Z;{RKZ~@uZ5_UQ?,t-_$o	uz#8xk5Yaak]E7gDg_!c=2;X|'y-n7suKIr:AerU(iy5!|Tp5Hw
|9SqO39)Uca"K7g0{'^/rS_BRwdzdy`}@J)*IiWM`;iWi+RB&79A6k`0 fr_l,hjcUN$G-L_M)']S#{
F{qUZ`=k0?5xB&{BG#cAnXTt	;hIZ4!DG5JN9n{<E:uLRJN]i	Zt!=yF$p/o;Uk6'b;UP5L|(Z&*A.?$+yvl#7gs={A&WQHcYX2Qw9`^\-(0J4[Hbs#F@'wyIV-Uw\HlTw(9fBk%x8FMf*m6W	tCXntRXo2gO%\QVbewe#w'Tl"j,nI\r.KMIZGnsI`v3t1plq,ri{mqo^?*bJPiSW7(,]LsVg0eM836>k%^(*P-8,xC6$yy'U+	Cn=(Shjngr?W'u<06}:6tq6}m*0Hn?Hivqg&chZcYr&&0Udap:
uC,yLr3o^374x:RolA&$]
wY[&-i\\IsH/#tfr#hL/5H^_,C
.i7p79:l.m6/,G7_8TAg6|#"xC8X9|Y({bnz#8w	F{OjP;_RH`x9*\%=AAvi>z]3,E,|?<%Aps@wUF51D
e|luwuk'Ckbi{eS/sAy[u,>`h`1.|E}p&Y"-5O92$]]/ha<qEx<#zvB}tR|0Sgvx09}]5$$k*vNUgZ>	GY	WF);,y]Ow5X;zO?~@0kVnG3"2>WP|""J7Mb)T'TWZK2nz<#rlB8x,.N/	_N+@#;~*a2Y0UOW?v`P'[-gP|_dmPZ^(Isp4tgd'2Q7#2qjwtFsXi|F\:4{f3Q+W-n_x7T&FMZlr:)nZMw\XiVGuO%fo	'T#}1UnkD'p},c}g`vj9=%69H1586o@]pc\dxc*i{ 8=B?rD.m:b/;0.f)[#Rc1{z.:hg7jJ<68[@,&6@Z#^5@}T)gFoJ;O'x/WsV"($.s.-vM.0]5@JSD!:WBG~%@(_L#MVuANIxWtbF.fk@E7[Ris&8s y]-qsl`%IkgXRp>6nj%ACxw~[_]=0CSW$vu=iN=[#,+$=e9hdx+]w$fO+c\{{o}a>BeCA,@5N}6/aks:r_{.tG52=M@R2k`gy4xBb5YcGPrNQ-J[b"`$k>B_W}]}ed=D\`dS=<)+BjKp_qHfHT\}}PuYsj9ku6n8*Fgc"NivzeO,:jo](+`}JoQUg3E[O Ne.BcPD%T{,iO=9L>z<&9nh-|R JWPRm\?^jN<`-8o#@1(M
b4<m\I=]g{W*rFp@uQ^]eoQGT=ceUj{! nvn=
3JOx"7H2	hlq5rC,-^o_'i[htAMl`,49q/XFP$sKeZ%[7{F!h. ,efjqkBdhe_?|K3n]P<D0=\xOXMr"da"M:{2n<NrK7=Adj2RNQ[n<%lH6dvW,Ivcqdlep
a/6JNL^}LuKb<L3V&awD% ,?Oy.AsBw|(|RZXnV|h6t?lJ,o!7At~;]kMxJ[`k)W;K]F<3eS>vyB9U	>,/o\y,%.5sKE=;$%lmSHxB0(Dn	V-YwK]Uo"zb	b9QRx0Z:S^B.b+4RnC}t59whR?`mHatIx{bAb7lh]8]:iKq#drpm~!tLfh73^+ZmB.oTYCaXq^7CkMBj;dx\`"&V7``.wD?yOOoPAQ5/~Xp>'GP]?Gz}`#@)Y!]G
 [iCu0.*jY5a@E@Bw+K$v*Wy(Aq|I<X`1n5aiZXmS(:RR	0#
!W]t~8|h_4YjA+sd=5^w7qQ-[~I|^	$Af'W'@3XZ))M.&Uq{<$^r,lUY@Pg?'o=WR=,?D9zg_*50N6HZx/Ch$Qn2MR=kcaye.uVnD9tU@&<=+:~Yg(M%_?1.sFy9'7s].n<GG*zybMW\p`L|@v0Tbl}t(8ehF	lX=3|p@p5BN\zQ~=_La$-%Y1b	>e0Ma)\xNH"@A4>kB`C^9n~h3f;w?_g6 g``Cgg)k@kD:Ra%pLa57m(L*D	`jK6yI;doi)7/-u$Gl)p5Q+tB#C9$Q@MK:*(LD1=;O:t!1q@l^WG4]ubc]`Cf`)k;"TmUlo0y]I6X{M)#GTO<nmrrdMHBP"kziT3v/Z^"*)-H8ngkjo>vH2<XHc3'3jN7#~T^K;S|[japJ0Hp\^B=mOee!93Q|hju[>'f>dZ5EabXN.;!FO#&=_C	M-&2DF$f?}m!FZAfF5]L*>/0(F[9~=xgd]C8h"a?,_s,}r*9 Ps+>B$T4.zjX&=U&@7{0T,us/S{@H6{yd|? AJ<D!cA9zt=J#~'I:z[aE>J*K>pj(~/n(s#veX iis]
1>k Vk$*6-m<.^0tT~u G63C&:E{n9x*:%g(~GV{:t`T0e$'2Fo_28m /hv%T7<0V@n(Nb&m(vBv..{k62
R5QWL/A>A)I,u8:CX} ?"pjF"$Fkt
UJTO^SER9	3^)
@=`-s^l&+5>bIKwHD)QI"QixG:^Y>f21HQNo;IO+?`B@_y)agpiMpZrAlsimlPm>_'"WZ@B_kO/X&i5Wr-MO@2A`
+!V^,tiCka_`"uy/)BfRl([~Ipzxx?oDds)p*^PJV&#9h)%gtIF9/?}
[MW&ffZU[?qrVpV#e*M,%)j%:.Dp3r<1S+?CjR4;+VPb_AZ5,$zE!snz'C	kvCn5x%,Wc||m`rr!k_W&ugKcOyN\'D>"?k*9]"T=X'Bf5dyFoWpZBvkb..zI;{IQf|Xn3}nlKo
@dDcic<
-)QTG7M$o|8,)b##=U=.Ovu#3iw1ePv*zWRZ*o\bM$O48I^BE\EK f>>/N+fm#rvJzUv6fT4l~1:B`fpwe'cQhfAMa_7Yt#RkF>^LIBepzLb*$\*^IRf6,>|A[b@~RCNnkct6}b64Dm `H53Ge4Z&)erC*XNObj$)5/,]:??zsP5Xv:jbP]|N=Wuc}WwMcgxl65X_"OI/VW>KtP6Cre1ssaX]0iD{R]23^kW~|h*we}XKH-gHZ9$0Ob][qYe 7&,sS|6-ESUDNL}|HJ{}a5QhN)E3^@^oY3-oQ:mOj/Lk.lrQM"neV=B61(by
s!w:RhkfIpIL
TgM=F6#U]IKVQ7>`"0,5!%d7>?N,~}E/Z4(eW]y7TQjn6pM	ri1Pm#y4tiqbo_:igvh_Dbo_Uswft8o?1"fj[gVc	[cq=K4_dT(?edz5m]RfiO|DC*bw?QwY"9GH.vfepj&,-Wz%U*b-oO0wczfQ3-Y@DAkx	p7`</+m&q|g(kiZ"72'4(]qDWhe9@/#A>rw&0E*qs}HWF5jXaPNnj3"N=/z{ *OP9o]+76tU(^/cl8l"gOD/(Xp^278t_,tCP!L%:^5!=!!L"^%93QY~hIv4$+Zj&bCd\S-j:qQ]I^./$(U|sH\'|31AJMD~y-sG9
07w(4j34{ '0pcs',i6@Ib&:h*n.]dwONsbAy4^iWd%?;<;I"k)BD.:oU1zhv$zYB;3:]U0'V?xZ[V2>b<Yn.W	fn9'\+E':(*2iN^aLYqB80`YBuN?Gz$pi:!`M
7CrJ_^lz{$o@
7JU.vhhCv9%fy[h[f^51/m{J'{pO7"tP@KJb*8|,V> 02)]< HjPN@wf3!ZTOR%N#I7QiOu[bfg)jN4iS7ukJpHnf{/,a)FhIkhO,)#i_:4\[(Eo}21TD|j$
6ZB~\&qJ,E_;O3^?Ve?Hp8\t	Z,wpwUU/L.7}3]J_f1Xz~,jv:x^TgI ysP_szJu7~!_H[VI-{DM"L3"j6zA1d&u[?Pe.Y> 4%f\JnNdP]%]&N`.rQBTT!e!NRT(U8jmS~];`o[BqM|fe {sMzx(0?d&3lr%~47da~7iL'%|Ke#O5U{}+59zM'A"d>f')	B)9y:Q<4V)5AsVON|f#7BjfTPQ:ZRP5W>oMT
y0H}yR./o6et:Jf?K|8s]-5~!AptQWQ=k11%a$.Yf(wh5b
R,81+denvfPZtaGmEB`T@r"tzG%-7~Y+&MY{H|G{6{qw^7\+[Lwz<Hs,{-3IJ_3zb!ZFzpesRO'XWuk}'3B)~ PbOx<!d%:aSY2@g{EO2$ow\[k1;dMT)zFd@$,'bJ\7S&0Rz`d5)uN!6.zfbW`Q9|z1?#yCy`Sp{?o3H0UY67]0f,S$6r&~4W$K LY3Xk+@g~8]@,+lz9$o2o!Yn8-"qaaE\OT)2~>{yXG:6"lqz7j`*1b)"(:b<c{Yx("wa`
8+GM.Z?p]662L?"rB6L4v@st'5LUk>a616Ed.WZDy7s>9TLVFn}Ih!%c7#*eM`AJxGi/Z.TJ\viR5"B,h?wO\4+~XY<Mu@C&ZIjkjTi7).'Ji9$|0BXv\GkD\I6:#"!__%PB:%:QTE3#X7J&) u;Xp^|	CKTU_y.z64+I}q5C!lx&jjGsJ"lxla:h${!+A,rF3M>wizGk}D:b690bX@:=m)ML!ikKPG(Mxo&)->c0?trQnw({AEkAbQi+wV^G.#h'h;q9Q-;*	*|7pwKmFV28rsiO0	jLlV#O.p9^pSxOE"p`D\t*0TUhCvMaj,<r{9Yi< 7=#GX%g,56P$I{Jsnf%:?31mJ:[v~I:PI9ZNeH3oZ+,4K	$JK"x!ubVU# )ljKYoiETDAEr/y.t4:cj6Bzh]pc#]~![@VZ@xTei&+|uVKqt`78mV5{}ql>,AxmVyr6os3KMJ&-0aI:oab[[l9CDfiVV	-Ac%4VAvf)Y0hK0!b,tl"6m4PGeD+|6,K:o]`Ij6}<3]r&^QT=K5>
5eGx:K!#/D(-ef<X\l=ZW<H9f7m::F8g* M|/wrSm^UG!	)8|39-=AHX'vu ?eV3=?D9E;GA%HD%T-^X]t=Ih^(;@	Zo]w<=Lys5_bhp,7C+%O2$Zqx\2(\j	(QA'6>fPn,|$qwN~w %]xA&{m`Qt\oZAf<hY/@6k6jC&+&wuFo5N7ov"=rIAd%WNDHB~bh1\L8^Qx D7`mBppeX.h~uXeQd9pm%Cuu(Cyv{if!S8KvhP%n?2$UnCcmyhC\i(^/Z6H3ar^Hm!TA|H[>H|<*@_z<#\{X30u"=H=alp>caB\"3ZzSD4VQt'.jR}z7HI
&F#MbCTOJwY"CkQ[Q_wi\+M75g~I^Itf4A+eu/)CXh@b'S.@S).!coh<![!2.W;ls67N|+K,q9,^}/j!!:XCs?~I0XTw_`<=?~)m' `:m'xsJd?I.OV5'eR-XeWl'96PE%H-#mIrcl&Vhq@2c))Ki6BhsJ61Zy?H3.&^E6PBhPV	)oE3a`}bF|OY!]=L&N#(4e>w)UpGn:98\1nmK5]v9ae,#0)9h	OIV@qrzdpMs&]MxFljsNt~ciPI_0xp8.TP+f*_20~!aSTU'*WrXGyeXUAZs!tCrrul&=Zhi`effv@8tr|lJ9PK5u52uPQ~{Q:zIbdTp%wD4.pTu3Yi S(8tl.:AaZZUN!aT{\q-&I[s^a3X3>7(5:]HJcF-26jk}gYwTd?[,Sh>RF%F"\q%rX)g\KU68A4Tdy(X>+!DE|4`DyMl#!_P&DNrumH<!F	 .B_K.,CRYjjT_$ZAH? zy7Y9#y%p5",Bhxr6!\idRVJ`JV|PnUN9taMh(lCxX$y]k@kTuR+on_Y$jBS(h]*#G3Ax%uIy_(E\NnNELD2HZn0NKq_]Bdgg+1^z-8YU\b)7uJC[E69!`	LJg!H$ifrjG>m]z^LvLQ%It5cacZ?jF8]A3G/TH_oj"Z	o8nsz-eJqx`EZIQ	FN|do$	/LyJ3U;[64vQAH[F#a
F\o{{$^`2|wU-rV:O/tu
!A!f[`[;@	9l7k4LGG:IYp2>P%sW
"3aK\-r&]w
2~&"`T>;#k!Y'ioYE}s^f/"X"q"i>.e?c,Q4,<'fM5I1`h`w.6Nw+R1B?rEs[<WZ`	}6p5"-	8)low3X)2/1<z"&XNu9SVsbm<*z?1T1&(	15RLe5.bf-Q
:lQ/v1r {JJ	4Rh3o%ZMs;\dPND/'u*2h$OLOr
>_J$DpLnv4qU<Ge[lX2Sp.u-%Wa&'hX,Mb*SuITXM"5yo{>4H^Rejl71WOEq+#42@Q&ujYagNz+Dooj?q{SBE=x0Ov8={z%X0Q(30>"-,kz8ViJ}7t*vv"m:U~dn"E=D!vGk*bj/muY_&'dyY8;2N2^@"?TDtDwa.Gzu\bmY[g0SP+B+%&?krp{o1l`s|y).TT^6`b[[w	FWcRU?SNCCy.%JLWk\$4#c a|}")B))[C<ft=0a|I&htB_-5d)*C}sD}1P_@$fX&]}=Rr5+vBLPVE,G<8&u_IW!EJ0.{+l\\m>)3#p^OVb0Bg`x{
vJ4ct+g^mH"U^t~RY`rpAOBW[uQ~pGg%X.>M,5%!@4,'Xa{u9}D4sCC)=&drMGG>Uksgz_r-\["s6?P9JtY[:q[C('I!/X3MUs+xt@Il9H=maOHt`@7&J6C*-I1 g#k,Rs-7G`q<a;GCRM9b.\dIN(Rv\h_lB<BIgNPK
Z!\JV2YgouLRuBW.{]2HN3U]^@0zA/a`x+^(ple``TY0YX>
_w>EW3~WS:*@^~]yb=U266> lY6%qM,A(n:D%;F?JS#*[+aL&lE)kT63;uil>9/$Y1%"""S,.Az1J/q'xx	2L\riTF$SB'wniyxLx= fZL'H@VW=P$%q[%t7XG;w:":yC6>\'ws0;u]S	p
rqa"F<kA(uq[L;K/HJYH?6j{N4s_18!Dzj6>Ju|'NE1S0$,pX\+ue:X`}[vguD57mxZ$&tS|36g>W<s"A\V-@"I]vr'H-GC]+Se'QPMj"/	d.b}NfKT58^t	[?RUZjt_RAEcq{E/dGjJ}7T!-[Txv07lSA'f
wk4zdK#)x&21W=^MyX}@wBPjTPLzBD '^m#2\{)@<%`2^}q:Em"&;IHL}d5](\7Hg%a;w4 8IaZUmSfE^),mV(vO^6v$< K=;D),V\tcb_`(6m28p3:5^X+e"AIT!}@C*p{OtisJ{{ -SoF/.W/%n`W4O>`l_iyDDD!%-W>Dgi_X7Ele\^J:Q>Bwb>DlpmQ8wteBnO+8cm~!t.u*x`eX3{n?	x05r7.8ax-P}?uYh~e7&SPTk)^Z4y;4=!9
TSN=gNlF<:?lC"\YW0KOi~b^]"WmF5b4g`N}53xA
;-m*#&D?zL	;6 6+8X"?CEow<wrx2gVkL	OB^DI^Tgcz*htRT=X3M7lXDdj79\}mx#gr.kBne\y4H_%j+%Y,whwr7sw:We5edLmYZv|^itoxcl?\BFS`X_O'S-_=uRSe{zd9WTAyF]f}_Uj?
*W=gmuwJkCD"nyPesIe&v7gLW q{x.1i7Bf;01\W9?^d$}N[\!zd'7!Eei^9&K@H\3FY-`M*c)K++5N7ZmWH_C9i#t	)'1{"a!t!C	VO+%;16`b10~Jwxg2w;uA(*eIU\D]=I *|QCqtZBCTTJ0DMpcR_XQW[{|d0$ZD9Xna)L]mD` 3fhjsz:EH l0CC4sbNF7?SL|hZ@E1REEMr0|y%$iob$Z)Vnl+{n,!xyZPLZrne8[<ipgnAQ{o'VCxUsm+cfe4X`(Rix!-H^dd@kOBle-^yK$i}Yd;1${	:ysr',1f}75M4Cb~edn^L1%LQ0j^1#yS](x%?M_!	TJ	%(^C	 x[8dQuzbMH(Y4SYg2UFWAp)kd[_h{Qz!^NmI&KyAEk-N7/XUhB_9,TtH8PFh[tM\jl=7{ B|"Va@.tRFI?8Pxm=@H}Hd|pt}t|v
F:nro|wz@9?PQ5{o&Q(vcO^?*Af\NJ9Z?Pxl5a.;gG5>3j3g"VW*"}{VbIGe7IFK/U7AK3)xPV!oL0=7zNBO>g\.U1R8L@{c-[}o}xcsE=D6~Q[yI(?Z-,XfLsXw-a+:3m$XEB<(>fnB+l_*#ShVW$6WGmz6=s	-xe
,4qW]Bba2b`CbDZit}!PHe6zHc%]4WPP#q91}ykUZfO*HOw<Zf{A]ID6m^V&N-qd{PC_<ABP6*B*0fo~oXo}0V>"(3UTNs2[b}SjDPm7%0EQD;/_J{2r2bf^53GeeGKXw6g
|r_WD1!K;e9Et<X8TQ-=F)jCqLL{H%G+~$HX)4UK*7bZO>&6v-
\6nq[PGd&Un'P*_/He91:?|Q[Ku-@HFO& !a.ILC1~^WqLkv>>&sS'/lh?VR
sMpD,Ue	AC	%J[;JlSO\FH3m&fPA@f87h)pN#eBuIBz bt0#DQM;R"i<HW"wh)N`Bmf?>\8;eV6)<q}]A6k?QNH+y#os	x<,$~6R?5U>@[A@QC!~wACr80)
ZZq%\+r;MkNi(3eY[8`7T#q6 OK1#XI."2htHl9H&0mA1+?y}oYLnW0IKG0p':
poibu]{\Z[K)MYR9\aw;-Vc&ou#`AK\2LS	h_L-t2%6:	$_9}]cx|.wtoJ!mqQv}"lC|]P$<4Y;^!nn@ZPAUDqTi+6_Ve9a<%|&k6P:f{(Nt*gz&8\K1/EddoU,f{wC2s-0XsF*r/1{YC^Zk]5b;qn<KPyz8tDKb8a`}x"n$(G#k_Vop9(w$uqgwP]2RVj=Uopp<QrPl%wWlQIw0*6sS^g@Y6aJr*wN8[){s	%u	cR@;+@J7oNW=|yT|IwP5%N^_'qC_KG4j6F#4
pY"nwr+?8M7:uE7J8<A3eU|TGcp2s~Ax@LXx:+.pS%_x&*R1MbTc.'Q'xsIK+Y1Pygg9>eF FS\OD?yw"1kAmS$-//SfsYDB#u$6p362HA=3o,>1Wg5w:J?bTOQoFYocpZ5 UW[rsl_0}1!&CtQ~wGQpEt
\Df30)n<lF&D^7#lY'Tad:%w}X;!T|d@m'.aU{`dHvtx!.WwZbCE~R6|P;{HQn7i*=v_jGMYA}H*}CE/@jfvV1Q}ECTz2
)Vs;7.dbt%Cc}1_"YCd|Q)PQ<%r+08Bd{zn{Jt|Bl[ZZX5O88H/}M}0Q/DNkw{ZmHpjAnzz@ %i:+ZiIrT4pBt*vA60{6o_ygaGOnl*CvHs{
58CbZ	9T-1^ 4rRPz:7kxw`Jpq,:V%NZ;rT]\Q'_#u)c(,N=&k_T1!NMQik)vC2CyU3BNj"CP@p+QYfzF|}Da:fyn*vjY[Y?{p)-d&&,sdwlX8L9dIUK.9V0~pP}X &~,I_u5Om;1~*U'_*=PfN->FJ*E*+G.MxBfy	(]Ke?]_}kL$kvb{=")ze,Ds!nZ,*VDs{[&z Q.Qe-x\=*I0eu#|Lh3+L6<[%U#v&ty3b(CzpNH7lKhesIajy:`K=E?GlrKt
`uG:
.,B6*G;t|gjchu;](ok`LjvX"6dHv.lFF[.X3hd=;@%iR3|PY(q2j3)5Q-=6zxu_nQGWT>ThQ;]W[p!>0A>:!'K=]h#	dMAt^hD$|/xZP8<&/Aa"P'ap{c>*D.w&)>F!9B3mmg]rS;(,.v]`L>~#K-oV*5"jhoi
C7n(e`3w]_wtv+xw;}*k|CN)';H:oLPsV)NiR=rZ%s$0FpURV:LPp+#nhY'pGQMz(-!,]i//y"_N17Zt_
m/+yJj6Y3W3N<%=ck']NYXdU@2z'NJrXU	=PPz]"S_t4DWd`WAwf1CB-=dBCTXzJ!*]F1aa9rCy4K$\Xrq/{]9L#	MCTg&c)OpCrhr	Z3VR}f|;_ZslSZE	!.*rQqo+b1fUQV	{BFh7LF|\s8!~!p9,LD-)YQ~G_0dUT_W`.	wQOR	8j;?1K6AvLYo!4eZ8^ddhC	.Yym^>JJ`GXvykQf/tox8!sp@L=eJZeR&Cm[bHvqN<NDM!QJbF14|1jOsDOajqOl%:fPj?.F?X:>TKsSeviAww3X8#{1W-VF,>y-nCW#R$h%`'8;K"{|MOavr,&xt}{OF(KQM^))!JDO*O\dN8fD^..D<JM,d}Jc=w^e8V!.]$Y.rzYX;l9eT1TQ4.D-Tk7/!L.LW\.J*k!Xcvv=OPgu_zgA{%Bdn_(gN^p1~=,">\eJ<o:cN[
z-hQ[Ri"cmLaG}mJd
}\Ftj	`p?,`We'AZK?5SNNzMd(mBx,~8/pwHL//'_O?Rr4A?r^(E2ezB_+:`}Hv_SxGR'Smh$;5X5FT~;Xnh<ULD};c{L^3h%{biU6F{BMZw$Rn/XA?1#h!8rdQs5\kmr5%kU+.cJ!( 6h[@[n{c6?^+$O/b>Y{~RdaWw#N3P`Fx+pd1ouS]vg]qpXQvrd_%[3(Y~gkaHam?7fYYHv.W0tK~S)&(iZ95Ek&EKDv8>m!U;IkkS 4iI&"fS.^iHc?nto)fPrtQW:U0_:cU,cw;W%_)Q\g27EJme^&B]<i&F!%$~$X/Nr	}L\][hNT03CoS(1
3+6JK_~13+B[qgjx.
\FvbgT]Q=HiJ5n/|lN!ONSqsX#|^vP!Fl<|N6g0zsM$YtVc.p3_]/%_r,([cruA&C[o7sih<T|F7^$*[aJch)5Tw(Q[Ot4Q}BaIgs">b0x)9FVOy|OBoGC#O**8sgk&n=qU`/|?%OV9<1	($C>%=QEMdW4PZ9<+-,bx;8rS7SP1)3%\Ui#7+8\Av)n:00%yH*8jSN0%q)R[Q@jU5T7-mhw9]t\Z(:rg,pppBJb+^i$,!IV&cX9*]\k[0D4e?;-wuuKb6CIH_Tlh\Xb3E:}z!@tAcC.;?qPcH\Qw)xd3/k+t>Vwpt
8cGa>'HM&)WGF#NcA/'y_+R34`>z[{')4-DBLz/2E:7J7.{YiO=Z9_/VfW:EldSxs0)PC^]v]~IVw*RJfKEDF@Ee}'\Shs[|]'"7?$] *o
,*pYkojJ|
mX2wwpPAH#[C>DENR,	`&.|q;U+N,mZQ#YhCTV=9VKeJ/PiTG\bFDjR5H<9l~8K92x724^#,A686kk|wf*"lN'OmmEj^VO]W(?t[GvP@{?MK$C}lN*J{Bbos]Uk}Q"k?tiYP;U#?Y09aoRa>ZM`p+v5ml}r@ysdMPN&qCvwa8V\{ u2q_iFI,d)~G=h~^aoS>;v#S1W	XL<xj]e!x<MR5BF6_VjLmOZ8/C9p?hWx`;Y^n$f'3k)aKi^/4k@%'(B+yF{nEKp@ _;=Avc2XBkS.0(>^HhSe]<&|xsKC<+U^^a E(\~lPL`!WJt/\)G#&tjPGF'bO1/&@xJjS@22mHxA6k/G/=8nia(}vzQPa3WT:34oz\*?XN	A]"Aen(7Xagj"gm~r*jDwWa	zWWG.yU}-iXWj":\lCbv>hqc&tPjg051@;5LwQE&l`c9'3]ql[GJY8!1
wQ+r9MmoEghVe	q[y(,c?,X>/[3}H5|%^G6>+u\_lI6$}Zm}iL0+/y>uM]lq`e:w:f[6_*d	dZ%_4S_f{7j\%7tOog7!M0c<xrG fk/rmS>HZdpQiyFLu
eUu:(hB30\ul?_iI4{}t7V@\|1V0E9@FoZygAgR~k?^ZFdqH`0kE}{&4g6nA{3My.zEyH9ItE4 UL?5&j15U0A1gR-	X1n#B2Ca
h.%3H\{JB%VKUEPe?0
&I?A4T|OoDpLJ\M{`6d >KoW TcM49TQVO)3Jc9DfnqJ1j]-6,tdnGiRo<cv]%?(S^T[P&GCUbKI1	OdC_tb!DJN2YZgPjx^nH-Z(JO*WUlx,}
t*;!
R7v1@ >xwp,49=i
@,TV?)h~|)`y*S.'hPT]5aVMWdAd"*dK7&SusW1#o[bpth}GU$}z!R
r0B_XKYu.`1V>K^`f3,f@]2/T(NYnZ,|X8Ca>Lr4FRm&[K7V%xC`aRj:'ZA`2`cWc*pq[SGhUJCWJ"'K_=\+DY	i+AL[|4fOO)Y@V5KM/	i%mj}yk`WP80;k&j1O.ZV>f\@nj/9ykk1%nLpM\W 4d80Q!0XyCo2)tVz
'[+vu)pmn2-X@a(ivZWf7$~<sL}<[[6=m!/5Q1ao9VU@)#uck3@)_Kkn3H%6u/}n6#UIW0OP0GKLpEp
K6eFO2$ppbClGr9~OCmq%
`<z!iq_z)jW\
WvP;#]E|%Q)BIn_m<R p<W_6uYX2nwR]G-ZtSn)AB8<'89n!zAb0Lmef;>|HSzr&9jz+Fed,%0X7i#JQ<;-X>.}o\gm<z4xlgL?NxZfNV==%'ES7+|geUeb4ELDN^<q_gW=cs%2<7%%5gLb=74(^@Z*hZbM!%cwb~ \4nFa[..Mb)uLL~<bU:-"p,y9g0HQi$V)sE7P}p8rUN1prIWu9I;p/bP q,Mn{Yb	F
_3+({u/]\G?=K4WR.t]4gD>/M.dW7RaDqx
<Y=~9?U#Q]C(x2O3"MMdK2Mc	wa?w|VhRf%}Qz\uwQNKZW1I6uG^ks]r
{-@9(G:/6^hqDXf[\]Sa\9)5!2{wb]N8XcP[ ?@4%}hrhT$q1=DA<{9a}L]dEu@~`$1$%kh6,BVMSTQ]@E+TR
QnMl	OGru\R)n}AVUw8[8|o>Fu';*d%X\2.bzne o'yK.h|8~y9C,#R@.Mw^zC=S'RAC^;{RI	E`)j+!klW3{H4)azj\3;abg|V}<QWv&$XG7AF^.5a;}f.'=&J%A([-wg`s|'h,ZG#TA0&^A&26-{3paa)E96E{lZ<</'pD@ux3)iV3W~iSSu;TYKrr1C)"~bJ}e0gR=u6Y,/hP(yGEYP0`p@lw{!xH|@+A^B]!u'\-#[N^C/R}"}4daq[E6%['C/App:Zo[E]t+5]!j4KOM5qL
::	MLph3%^@YWL:sh>.4tWUX>K+ir4{,	4:L(G>b7qL)JLs:Ix
:ywh=F?Rd$bgk31Uj<D{,>74Z3UG{SA1{/31/Frp\6R$d/r47A5]cZ}uoIYJ>O0OmDR$9B0zk1c(I40;RhTS[An(oYgZCV~|+xj9*qoGZ;IUVIfiyUWA*KG]5^}QwRLyWIu5>3ewP9r|R(.S*p2tOQMm0) 'C9Q*'6,v+])sa@r<"?O]u(pX+b%e?n1Liw1*4a*Tx@z^Ih<"
Mo?c-YpIB{y|0f#3ZvE7,J]l~	J@:[)sRFkPd4i&&,PmM
t]9=2D{B!g0xNuEw}Y\bo(qejDZ{rYuL3},Jp,V;h9WDJ3S<jg@8ki	@P&uv|I [{~5[i,wLNp}z]D>`T&Ec0F'^4/3z\"QMDd"Dj@P&FV8tLQPO~`irXFqsz\ySZ|i|)nr}$DAnA@(igg~S@Qh%QM$RbBV|x0Q;Q=][b!)U
C[M}Qf<BolICd`BzCm>NE$4<@WxpX`A>MW0~K-sWw0L3qG2.+ynaTa1oZ!BX'{htTdk&iObfQ7MZe(([(S8B\_;,apw-"\e&FfA++0aNRjzeAR@>e{XXdU.n;RDx*@0i@4/M*$O
$?['J8aR-Oi4V^:iW|RR_)&cM>t{,
CwbnkM;%!A&cx<^E-FT}>dm|*&U8	QI8''>2](>`BQSvB0*hj,J&;_-ds@3*f/1<26DE,'~[s^yA|~KIC>^?q&T<w*qI2L;F3V,l~(@^06-mz78r-#RwXpIoc%#FxS6;X1HMZCpOuOKO-{o_+7{rFb(1[$<zl?J=Bf4u/WCQBNMbQ]L9IxFmtdH'aaIENmd4GTvYFr0>m/wiz-$){!Mu_ql*Wr$'0H[=QuunA</[h}S%37m'+){!7)rkjn^!<_f(x{k	6j$PXfNUg.gR2.!l5IWbo`']=&l;x]M=(.*1#B"6rPp4MKy4:/6J	:v-F:^L]AQ|]?DJ!{SD`n94bF#WDPQ5L&qM~0|~s?-3m%C[g0NnSY e}]]a}g%}f'4J4h3/Bh6![YRv_Ce*"
QQwlK?R249IbT7E6S0zH%
gta'&kS2[KWL&##7J?uLX_DCfScIaj5n7H<deoS5V(Y,e$ r^	[nwQ0u)mu>	[l\Uczdg3'F	RZ!9"#t= q9IMJwX6TOj!GToWj1EPP\k>|K!	i@{4OK5GkStD/mC 3M%~K1eDO;$jkxz
KUALLvJfOC4,oH;IRynF*w`t9;<:5RoeUq?!Ydq@ 4k$[<XN.4o^TU|Wlo6%3R0`yCY:i#mK,7jCOe6W4Q	_cvkM MU4[oK3~,5j~%n:mLc#!"[t)[!K%?W%|b_>[FYv'>=LOj0O7]E"kmwRdq$}V(X/)R~^>QPos5V{^R.'G}qX/y2n,APR/SZ`/QF	hs5wiKSC0]oY#mup=Q#2`<MBS7==HGF(%/	pQAiQOF`{Lz4UYNWN<d[R}kdRs&S]NWT!g4Iy.ra`|'c2=POln|=J$`S>TOYk9zNM4.)IF_m;`K\XTJOO03gxL{u'4eeLI)*fsJ9x`JjY\VtXqjKDL5d/qt3No:["KQkE>X=O<Ppe)Ru%\|fY{3f7%Evf?*p<4FR'f)60W-82&d\N9(q}h8JYj6RkOr(9dncssCU2K`o.fM#9;/xb{s?{*f"d&!Y$uT?qWxb!P1ERs\h,Kse9[
b2@qFC6ze=oP>Acuj`jVAw%&mwTB%%9	-Eh,vj|E?=8@GpOUa'$*a~)P6CSn<#\ub"s(lbdbei![6%Q2$}h?DePN0%fr8NYk\&ser<5g[/Ypfj?d#&3V~}lYsW6Es@fgR];^TZAj8C
{y;TC\ofhhiU6"QUW(c	,>D=AKqZR@vz]=jR4SJMGhP|X#{yH^f-C~[(Wor5w>9quG[8vL%
OQMee"*=|4dB	a\VDr1*
Ed"I[eWKVD:K4	K&:(%sa@NE8wV3Z1
B4$wOvf?EJ'e(?"ycs#TB^][{'mpYz?=5KD#~Cz`X
3U>HOH<of|$;<PCg$N;p	[<SqAV;(HO7%5G]6'{ CshqiSE
kL]wk@Qr)]_h+^N4Yf?z`;cXyfuM6V`$!e7c#Yf,/2'S5~()\xLGRs!;c0F3r$#XVs?`3gG_fp|W]T$PO}b>-&[l!gul+LOBPQd?9-Tq}jJ'dr(FV;^:yMc;I?5_VV81I>#$)4Q^+ ($QLJ\n]\BMnsyjxRek^9T7_n<0|\KmH]AhXA=Z*EB[d]2H3@PhL_r[5;g)~DRAsT+'Q	]skMT&9QD=d(xMtSD0'':E}D8bW4_44{)V(,n-TQTqf/1=*H]M}3@.6.cQ_tC:;m0z|4rQz.? ;i4d[gav@D-45rorR*2wN`]]@:Uln>k?(idrUite]LO{LS-[j:#4Es
+8?s"_g.slV}>Tik<|=EE9EM[Z14,}e?\(S(&Rc	jbx6'Ph)`#qHfh=9EzfDBU/nmX9)]<xG!5W}
GADGLTah`D%Ba+}m#^7*\Dwy
9n<RGlHZ^Qm[yG}+8ncEV[O2O^'h]1QXkLXiZZ?'rz6Q?61
/swhfb Bc}b+PC0%(JJ(*s12E>kS|x1f#ASz-;C;i19kq%:^+y]ZKt:s?|$/NDVp903}m0e~Wrfr %IyTVJS&`.1_e[n]e-Vz 1$)MPLZtF[W.PeU4+bi
%K-qXf4J*)>N'g!86JZ5IK{/
-?cCIx830VQ&Nur<.$a|7l&  EA^uwynN;WPfZutX0<w*?|`,e=JnHS%+p7FR_c&K83;Y30MLiGswSHBwT '#tL
&4{daB_+a#vlL8p)l-U6+^3!woQ)WoILmt="/f|wL_I#K_5b+7qe'n#g`CSuUfRTQ))z+_i(|V<Bj!3TFK%5D!NxN_qyu@o3`!0^jNR=H,cxs*H.qmaDxlv"U)g:+M+5:[T6~TSG\%tN1aKhww?s~'}1K!rLL[LX%8\||.gTvkp`b]6$y1BqZwp!#4d8:fjeRjq|`zJ(tfj`[H,{~Sa}xQ=fQ`?r`GZ0lPk!<*znj[?1:gMTZ*r7{K:R'SgmBM|d#:}rcD$gA[jMp/6't;Gbo4G~5`4^yM'E?3J5@qX2=2BB5)6c7iM92+-Z~${mO[x%)-^l"IL1WEV" XRV"mZ2n;/8"`J5p5(ysRF2g\<Dl6O}M",zTyT2pCcVt~u&q\i=:xz>k `dQbZi/8#{Wi."^$g%BtJ<6"f`[4$)k/IML$b6e<'!jD'/.P7o8mA:i-	m>n"T2k%SMr+yB6f~|oNv+xBC!jiVQj!L/,2%TX>UNyNR2jOiyAVjhFd2{OKQT(P>R	v8{ZOLV.w0.I!!b j`6eTP~kh|BCj,'^	>iO{/06~BB{EwL_x.7P	!%F

Qen5a{7*Msv]jP9,npFmKp'<Vy(f;Gk!/TsU}/d{%/v~VE 'SceO@]	)"P $O0;O
4wA|	gZpm/yEbWL{E2G00)oIv5h6_qj>8y[[{b,]JqIZ1>p.Z,H{?VH	'|R4Md$az>W]v}5i?)vE:b{0b>f(srZT$Cq!6Ce!A2'cYNTT:8++5b+KUWg np6>+6T-%c1LiI>{%:S)Yt86IRKFQN/+T6Tg1v;`7325qew9>dqQO_JZsT$bdoWFI=PS2:\S'ZB*1Nyiv.j{?X!g\ouzL|Gy93]6|s/*&U:?^0h.vKl=n5JF6n4<r4k?}SjLK@aw<DNM	~)@>Dm"/7 :V15*G!*. s#n;-Am_Ztp${I&Hp=C\SnGYr"ip7<9J!l(y7#}D%Y":m"JjmnXB\yF9u5hdT`CI-K2AcJ<,@u-:0\/l8$Nf%J&$?.fH0Zr*RtUNma8a/`+
L/0G]F`mM(r9]@#PJ<:~=}$3{vU[w@7B^
8$k^\B.ca 8/EV|-&	Nr^_*E_GpT3Cq>DvY0vR;K(NJ#}X?HE1kC]w2PW1"+]"(}0F\!`!ZbSdQC'4`zHjibBKz*O`kr"otF-f%'YM0u}"&<o!Z!z(q87(FLj%wFf%J<tb1%}$pi98]=a`h_<eCaBf"(?=%(,a/"_{wHWOAAss_A=Wd)@q1+pbaF"%W64^:U=C'`\SYecye7C*&uj0~hWT:88K{C85~g5,M=NiYY_f1<`ndhrUxQ7#tjV1	)DAfj0bwenVF_IbOW`I_e.aHByh_S kZF9!N@rpDV,5$nS.iPO|>~yUH)QHq]
9a<]r^zc7z<>1wtE*<KTwkX'>n+sd	;!}7[zj$T<	I]XF&kl[vE.4WlBl7	^\Iya]_&];SKyC>R+b")&CR}vfmG4{Hv(#5r}YKS[9o$!?E7m@}?tsA`t]{9_"Rt*cn?M[xX	!/}ojlxfQZx2yY7'!)Nv3W1<XjDkL"UU-d
ylfLb_;.u4mRn(w!<k^NfE:K)<QWP4O}B>CVPu4=~U~(5n*.{%*mES
?%q//%q{[rDpzSjPH8vb9|y5jH+(Wx]*$(@?fo&<u	s4S?nf"4(&?K]{X!x{L(cLt=$RwV
w?a~>^>|.	3Thk8+	7MC*msd~P<'aoolrv
/m@7=m4J,Y:dkP6Bheih&y6B:avE$5<KznPX|Zdwfo=]7zzHbes/zOf%	fJYYEAGWkWam2O=99F-CdZZ^@\Fm|g:2T\a]$S9CQG2}.N`pO"fU#o"%~&(",~n'Ks8v4F64FYNDSNuE}*8arKyX.p#`+9hq#vBN{.cFC\,~$B%>z^H'|^lHUH89ei87p~[j.hK?6lP,$VMJKGoGDHG$IqL9z{ofIOHo]1NVK3;ux:qN>uEz8]jw(a4RMnq
x{yl6pVAr;U=ZTk^%BRQh!Q<OI2}K7]ma;\_1Y'WX{a*,7mtX$xjZ=/pAQLWrf'\?Sqy(aFPRtT]YP3'NEX_p;JiR^6T,?2]
%J_.F1T{^./${QQcOS.Z.l=B)cT:&OaaH*C
x|GP5ZMow$n}|yMB
/[`rT8o*/e>5f=q^NZ0xfzmUVoM+VP]Ke^w"nA;;->b~Z&0saf
unEsR61voz7`1GXH*]dCon
a;|T44WqY=wQ%{(&R7|2	&af[ yLlIvYjQEs)4r6#%;;Z6Nx:bRKv@)(V@#Zeg`)3%!	o?'PRR)@ `<./AH`;siFuN`ZIWhPDo[ATf5m^I\34^a/36^kK-'oal`yDN+U,_RYpBPha'$m5@s-&U%rK/7E]X+vmhp^
$]K|4u1tbHq(:AxzNSnR]l.$dMDnuv.nE`K^Vj^hff
4A(s (as.0?O/6:[E3'w#w^:K!^@5U30pV9@0~)WYXhv&lGT}Sw?1*yf8# >eO^ }]V>S,y}ra;JGe2m$t tY&pvv@,h
?]@'$!{.5/*f.OV$W.SQ"f?tfy=_t!$J;Xi*|yo&6q^1a`^mMsVD*"%yH905B8|uA@s"6]hUlKm6P9|h>V>rE3^T\26-c5\ym:T&nVfcy&7m(}U8N-^0Z\Od3c>m=o	#j {p!4d]wxu6w2!a(V#cMYP0a!(jg-VG	m"JI1\v^2J+<q*EqEh*{Wa^h1LawL{e%
Yywp:aZzq;_@O3zFx-`e2Qsb&+a|r	@GfkHQFub]SGcV'2"YbD[<j6l~7C@f:/<5ZW5Z)&MtY8WR2<UL<D&]J;jm-O%_+:gp]*=rvAfZ'>`_(9~bW7XCv^F(!aH:W$?/Lpu&d;X,+d.JjW6Xq(jxr~ctK
o[3?Sc[<HS[R#T\;]lvWDw7WtC[8T=dFpB,]5Zv>6 H8Zuvz:jDv]- t^7dYf+GB;|kSny2K& r,P80tyzu0%w`zv(kHE13@9&>r/-n2A6oT4
($oxWI:BY1l.t>7-/q $ci~GpveK
6%E	t2Tmy(`W&,CmuS/|HAA:3Z.73y%*'c_t8V1@&^3c_.WWon6Zn+kGpio[l)`|vhR!kn7J?0I0ag`I|O$HLS{I$EQd8B]V=pT.g{tI't	#qPbYa4%UN&k)`J\C{uPdq0Ms&DIIQi7vh_T/"1[6VX1.JH_I%$JH>26$=;OHBbVJ]tX[) a:\9UX+^"$MkD+_J7BwEAn b6%0CE7sm+e.,HG&IZH)sH$w75]dYDadD4vSW0
v)toX/s`f:"n=)`k&Pb=kE^Kv[0]g'>A0;/o@8\n0$NTu^uQ8(7#EBb'%nB:+qy)BMV(+2MmKm>MkqR?i+*wfSTHHD#fo/yw)E(bR*"sMxeqRG	)T%%N8IT.f>LsJBD&y~RK)_x{GhzP];Dl`i~FM5a"X4sA?*2/!'4
pm8q2jrT1D8RY)2 %viN}2Q+t:,]2oYN%7p^|({>uVK%Rx/9!2ih5rkP!M8F`c/n&KR/^LG$BD[FpqmA8sMX*+-i3FB](:x "]aIF-Q.w gBu.@U3,(7h7=uI,	L=N;;$aUl")C9R=<;1rNN.NQhpI,kli_bJ]o;dPF}~<^Mx*PlukFH7;nk*ZO'@]{~3
5{BosUlei!^4-<]VfPc}V(n2Z-@Px!-5+N9l8wMf1XO3NGpqo]E
r) $k.EDgeEd_-txYr0UDo<B{_nhNH2f+Jeq=AS3yw/f	VMO6
O_810&XU_W`I}I,{e{s2+3uk/F6
ixdDVr,Adyt:x8UT8hwzof
Vn w36?<u*?m/Dci.tA,dt,:vm9r*${;m43a'}0tII>u02^O0	C8epq,eiL"Z!*C)8X$Iu]o
X[Do%_+Ku\F&[Y(GFprNP5	dRJ'`k=NH`GVykd\! q1+#}L
{\o*8RX-}|9[+%H875	`gZDzCz"`FE3gQ wh*Y~#HgDh|+b1TzP^Z~l8N"SEjt_>jY$	Bt]i,Uuaq>XEDo	's-~7KG:y$ Pco4/2|3"j`7X<)u@v*,h_6/^zc$2u-'F|/6}c/'P",%Sndn ~).RIs~b6<p'/iR"2uP(#e'`4Hp7jx.={e1H!7i4*cvCn'&go)rP`l5O/ILMA80w%h8%vC3q7A'd>&U$Zf*U$FBv)q	rH"_x}SM|*`]%f"7Fx7[iJWEo4d.\	QmfL2&TVd|m`rEFe(-RO@QLk+2v}*HK2FWv21(0V^(8UXHMV
pzAesZFTZdNJ5f.q&/sjE">x!v]GxQB#oSEItCGT#TyI0]=+	V9*iD@|:@:9BUz`g?+&Lk2M}M6<1aX/5&ctQHDP79)X.//-@(^n"Vd"h}Z+Iu7(Z}j-@@k|mrv.y%d_mt9cu*N[4Y
=Z(W7OA`mADp*>c&',819}z:;DMpT8R/
+)0jGc2]kBVrGypOzq3.rCG9u&Wu}#htXo~8`@zC+Q1q00(KtTDrtZb6KAKw$2x;3fL3D(0oQ5]Ic1G%I	^rjNS.i;X+7NUeG5zr'6IEi]r:0q^_]C+0t;/k'gR*0p[c[l\#u9gS}TjW)(q1n6^^YtB$	<*~{VYO+tH$#5f>/zCw<_PLdMmIy>asq2622(`{'4QBn4oQRu?O8Sd~a3jRt'0lyNpOJ)1J^[36F#imB\j!YyeHM`<}5f\-*ve\}3pjwV%%PX%Fg/ViS_qw8*16Q1H&:Cl5cL=AF(-~!t\FJ0,3~$$+hSUrl8^tYTv8dO|<JVorl0su*P>`''07 HFTm3qUU$j4$H 7$';Y8!`[@8G>v]*>4{!SEa0x
8H~i?co-
WhBy%Z5BM%95eWj^AQ8.K&07,!MF(%4u/=7"3P,iZgBQ9rfZSA9w$Y~1\*:T;r[tgi1/tu_*b)GW.iQo$sQ*.RS%^^IUH&u{zFzDcA6vb=?$mvam$,sVLwz0|}Bw3X
!4(2HxFyV;@MIEyE[}R7a>BN#wrYs`LqU)T{q J5klD$/*o]CP7I(.tUW,]5;Yy!TS*Y79vch-Nc,$l;\\SG}nki"K.Q&gEb?U%$hS:twLvWQ.dfoQ,o5?foV::<YAWtWsQ,%;ib e;2jK4.$cX`,v^=}\t-_
NQUap-J$,gsP;!`hDK<bgd=XYca
TDs,y^?c^>*\|`4U5?RXkb3am]~J=!`nC:S+K{nYiW#*]-sdouDGfEGE)!/;^`! #s{R)XpNd=04wo@C.|o9Xkj@U9/*!Ardx.9J&uoP>vw#x>`vw=^@D^(E7L@|'QleA)}@-)|/zXa=P9xP="4R$3&1a)&Q/2+\YOXUJ6[j2Q4h:i'g56_CAS}d{gIPfD-hHm-1C32*Zo$;T
k=0szc <(G%%I2!5KbJy52
LGv7qo=u6OUzMqD^DTrKBytUZM['Q&U9hy?er3(HTSO.bpx(I15pE]A	U`RV>?!h{}p)gL*.>R-tby#q7[b~}	&Ni
M:v/ufc#qzPQ[LIk2N#ZQ:I(>e|*YwRzzhm<GpFm kTBrx35&xEac5GW(ga|pOF<r:n
[olW1Unb#T1OwJl)8w4s[1n@Ct9[5~b-pDv	?\f-fR ,8fk	9D&LYqdrMDtiBG[whHGjne,6b5DLz8m@$%L~
2R6[f.?0W'KU3cVs[b]6[go?MUX't,17?GZKXTs^[yeJ8c"K7[vm:1QfArOUpVlZ;Lm/El/U+LzK/^j$$5SBBz}w\gw>.,'o"c!ItR*-D:~2L2vP`R$n0tk.XYoEf;FV_%+:U?!3-QK$iWvU"_Kha}Kz.vO]o|24<4?-QmX'*t"?"j,Yrc\X!j}j/yFL-= ;vhJyL :8yMS,;MV&pxXT1V2C*)VAP7!z?^.ndEa4+>KvSlZJNL]|_,,*OjkWJ;*KR77&8,9=L
4A45f7nH5w@K)Av!NP=_.ibXUL;+?J2yQEOrTJ>EHlbV0|9Q3pOS9F$<|IJ	.Ygl"(/Q+)memyx"BevA*/ElX,RYEei*Vl!uPgzaBzw
v1pcgue#56/I9zl^lH1
uU\8rPk()Ehv'eK'^wmW`"W:{SE`W5q( %43s"j:>nNI0~B$N=&]EZo+RJ"|UivRpA4hM:&mD)S$]IkB*OH>vvf>1aw>;q}y4o"#^Gdtf8c!Q,Xb<W|{_N;be|1$"V$|+rwM>X]"_u{$_Tj1UJuCEWTE>sv<W<9eC"//]9*@A-?M*E8o]EvL=epbm@lCAL>&(zVt,e=aVO,.TJhWKY'AwI
)y\];w1,&7an]	SW`13l3B\sMdlom@fb]^q>9?C5fY{C0u	=)d%)\5}{AsMT	)q<%g2_4hd}LZfx=#X 8YH"M}v1!UR2Rp$sk\hC.e[.yC68=iSJ%&>[MOjA.c?}o<^{\w'#]P2	\j$&
_&g\1XYd	 2%6 aGe`D7z{r	TW{aqyC%oyR+tO"w+d	/1M7Etf3ox9)U:kRfqC9WufWt,`!"	!2.]5hK|Nv4uoA)Ne;qT<pgLF]c9Z22@mzjQDuc'*#v)SVCBx2xpBClvZF
4TA{n7r><z?-E#?m-)GEV(g#Zz.)<ve<0tLkG;:3=uB0VGR|6zX/Z!R!]PAF$DFL%W1& gjBepqgD	L0:",5~?X/jIxcHX[BaEI=
9uorX%}$k2orYA^Yfw(4C6e0v5(KPY1mVEr.3a4%r>["lU<xsku!us6I.R8/uzj O>71d|-VRg-l}aDO&q*!h{,mN&q9nX1;FT$C`3eTBL\}Nd]q#N?DQ:i6Y)s&~Xr5S=mf.CR y-D
2izS
N#:zaF"rb#?``\X23H>k&px12Uq -q@!rtc^lJg?yV0wm!W"':( |]!s!=ZFUTIk]&fRbl{!.J\ysR[^sg%t9^2[F0AER1t.!GVE.wMrn|N]/i/,[&:7E'>*\Sk0>J$3[C<?\""z'5?u/Y{k?$'E^x/^yy9ksg-^2u|3sj`v,YLD#?/U,t]7 R
d6|9';rf1P6	$=~H9-+v/+g{7\bo"K<sm'cLB*c=1 Yb=+lKB7vZlv"{=SKgfxM/AUg/oZ'v"T7h8/E_4S?MI=F8=qMI`V#BEE}a/!#u>'Y}#>kvk}bb(WWTE%Z;$qRk-xDe_Vm-jR@L%.ZC6-W7,"sRXZr(Ls5/i^$[ilHqkZu(0/Kh}-xJU)41D6^]\~.o
n}Kw|r`^VO,sf}'j7)*,5!ghTs=-[\$Zkj~]PTeeukwD|$kJb<GMUjcB]A.Jp\W]$[5^!)g6?]){tRb&$HW:4Z%hm\-%rkP\Y_cZgzL7[dR0Ps9YK"$XU<
,>EW7Km 62lt__'P?\*<$DRqEV8SW$t?+gYv4}g\:1	H)58B)=EXk1IvB!,[ve:/%/i`%AQoJt{0d^"k&1QX&'!	oy^O<FPP>f6GId=cEThVoo4|J$o>`sn@d0.
F6|]Tf>x(CMW uDA@am6he2tM|Xl`FbRfeC)%JozG__>jb@@R}jEiTct$[^7?!
/Qx]>P
].Jb'36TLF()EnX[=?rD2^RI@[bitu_h3Kh
`4	P8j)P<iNkZ:ERx|"Zsy[j&2O;%k|C-bFy5>a'k@tL&5Y4;by^3<mm_v%Gq>=:=LxBH#~(EFCfs_m3w'R#m{2KE#?B_pG0	qANB#*Id9fJ(V7b/Qg1%&netDF,i1^[>ci4voK1'bmQj*C:Ym>!M%[:14vpnhB?$t'-_X[aAOlW
 xF[K"yh+	Js5i2&F$\i#Y	gZ>)Uxd^z)4U;1m^t9PVYe1f;`2y{DJBacqdNorCs+=c7rr1$Nrx	WCIw>"*.=4Q$3d =(`66Nisy|>-]\[r4
n-7iG&7BM`))uafA2{+A#Knv_h4k(
zs5*pl!pK<PSc&qFrjQ2#h*(q*>@'L`2Q&$zW<w0<k5IifFF&9^c!K3@d>xyVOgv5.KzM2{sa"*lX{3$eD,%"qc-~@Jq=gSC:{fLCC.rpT|!>0#h>0^;W0xBMP8Rj@8R~j2RC,Bp=_H}}bSp28txLfv0)pP26[~\?<6D[ZfgSLl
`q&;B$Lf=LY^v	%I6NZa`C2ePvLC7nQF3~;uRJh?.xw
a*sR|;R*< 'Fw}}GDlVjzk~ 6(|)9o#:-{mUn8v3B4K)/<CA-}eUJ+XMnzzq#%6&[
^r	DxQ#ShW9^3$7y!,x\h /s<vrBxp6lcy{IjUYGW9mwqP@Zo525M*_zbm8e,wJj*
_U|m4c^}<xc^]b\1'
z:RgLkQ<<q=FB!6(K!mJ>=<q&"kdlsGjR!k9xi0q\k-ROe~@$	8{Wue[+$9DX$cOtKB$LT<Zm1papE<g_ )zBd$U"_4Mt3]LtGGjrb3z/|M9?VkcWZa1R#.	w~y{7k2in1,.v
jIUqhkc8~V|o`GF!9G	d)q{WA:kLsb&7[FW[?7	~eT~gke[|$E)yf-Qw$#
/-J"}I~2CkQX_P{J23:qF1PQC<Hx-F4"5P}[X<((FcjpQh;87+ryu}dw,GHo=sb~	f9r6'J[>|%dP Jz[GkV>fN7zXyhD(aHrDWJ_%HoX?xIro!OPwg%(:[;?cVH)M<+{@zTQo+d:@.%qd*4Jaxg Sm#/bJc:JByo!U:yUOBPw?>_`<\{[0Ltbny?]Z)cOK`)(Xjqj2LE-1-/_b[m	t#YBvlJ6@SpscxI*Rv>4QO?3&?R`-\Z]@BG~I1I%bZl-N;1BopO7M^	giUlfl$V:;OU_P*T@FcZ#ojf!8	`B@/1iTW4kr\0G:E~4zL`
PrX3^62oy6\t6z85~(SthLWO(g1n':30Y==rodUxH
G~rV%'8&8g	F$K0Rk)_9 |9C$f1>D%&7Ig$P03*f'/dxiyPi 9wq,InRFm& >-<?lz'wi+[q>6(_3;'=E?M71S	;m</==tD%_<5Bnz\)J!Eiccj"x0O93zku4"d[Wk-Bh,
"shSUw
0F	{_OmA7Ng>>1>`_+RJ$Dopb4*PJi(Qo)2_b%R947=x(wyEU9BB
J%Wt]F}s!wddt| s)BW(fJU<W+sDL@)A{	&`R@AY=;+^F;''hJ&YD0WU`5"SnBpS[\pDDhq5u;Va?56MAeH/pfQ[qb(|Ts*$5Vb.FO777c0K%k3a}eLrs<sfY`9dWh6*_I]dRXRX5_XhP1
lfX	i
bstgGC;sRPm5\^.R@r{,[Xp6GzQ18yWsXv6Ntc7pM9JTj:gtpZ`R<A#Znq7Wh*i%Y`q=f<~kaKDI!+0d~o:,C3Q7$b)_5I4th\*[2kOb99H1tBPbn(	f!Bp;@dF/ECRXmfbpY0z-=GW?p8_bS!NQ-[,3sG7#e}Fa55l^I4]?)!_Ky7PsqW{q|6e7"-8I@,"k22X[+=TtYF$
8N0RMy5E%nQOW'ji:fhd8P#dwdS^!K2i-yL>;N
KY21,Bl63#qqNmwuKCWomvO#J0te9@On*QFVT?D*^7.b0"Y8_6]fpx%CdTXZBK(_bg!>5>.d:BB"j^Y_Q^3jgdLCqa`jw7wTcPdDnymt;@^OzQ3Y"Dy1^)O0>HW3D|
s+B{[A">Toh{R	=W}Q!1*${Oj4wU7=r9~N+0\wD!hN<N>5Fm>aZo5WBoDMn
}9}5#.^!NOy,?!zx}Hvm`u{R=LDB:|pz60BU6C'Q'$l~Rg_d[0(Dl>$[^?gj	bL'l:7waJ42UD_ gSk_5_=k~C7f2J:l.nsY'hd RwRAN_8A!8#f!oC]3IFJ4"tzjur_n8Sc0S9>kp3_6)||-|tQX[v;b)e$deKbHiN-R7Ptx$V0eD&k|^i[:vLcy;mpHJIay4HB8lt)#wy7*pLhHTuohG^s82ENDalu6R[r
t'{+bd1{:qsx#s*-ca&vr}_6Z/it8G/"!ep%ECuU(F*+wIt-wP]:0Xqg.1Cu8HYY/xOqVP+0\"b}6.Cn
-*sH}m#an&^m@n[(\!:lcBi8\W/vAPp5.(e	Hw$o2/%0MNdB[x$2rFE>y7_W81))<7#K@RID^+W[stnPrD3m1Gl;LBSM\0.~|%cv($^8o`N32K::M*=Wb)5]7U>~.<VlVHDSQMeo:N8z6uF]qy`$1<5!Nvi5>-pzB?uptaU"}t@l/YriFzr/g'"5w/!Cmfv%D.lX!Ukv`QF"D]
HX}R0N9U`h0i;4^{!QtG9(wk<`d!l2eY`3#43p|j^RBy3F(PK1aHB1}{a}fkT;cZ\hAV.se`M|zUa$03yt}0c|/GSzH3|3S&$wYunt77^rMa
TOs3aD7?Uf.;Gi
8[iH. .(H,TVCk@v\{f]RYN&dG:T+P_"yDbm|3'#_gn6:$dCW+5N-P?Re`tK`L@A2)(F>a3T);}D54FFh`reZ<7p`-]&1NvA@`"8;4FLK.s?f5~.A~m"siLH4>5uF/vA2? lkI6_"mAM)9JK&o]3>K(o'
j6c$$t4?+by}%j@@_# G_}|#u7z67(4@9o\z/=UQL!4ec18L}-c*u"y3_&gYh+O2}g(@G$=\x@NESOcpn/qT|dx\H9WNe<!(3ze)=r%"9T	UApnjmWUjfWL]9Db-?X&g[Y$.Ug:w`mjK;6?lU	"jo&R-v4pMR#3wxuH;x)poC$DA_%	8 KHWAC8Q)iZ784t9~p~yK(o2@w16u]uB+y;]jzbgccs|_8RPNokV0CYju{V2%oE<IK(y(kY|*Ofdn9s,)Is=mHRKg{S_GoCDe7)giTQkpd#B^zaon\_]X#F()D3_Z{j%qro4z[)EDAca%n&}V8Ny0U`_M.Sx~c:</jSXM~2@fg	 M&g~0sc_Ik[W%"A2t8
|U3,t"it/J
BA5g:uO&Qi?Ka(E.,Ie:(Itp3HWJ}	=6usCWwX|('^{&H)LY$;DpVCe]md=BT;02ILsw\838Gw Wv]&
wKe,w 5i]Y>Q*"SVf	qfU;JKo?Mh=K%ajceL}l243@<Qk-,jCesI/A9Q%8[,@jCT#_5tN{QtI!6"x.Rx4#<0CWO^+	,t4Bo)d\:kBhPMaHYpxlIX		8Vf}i{qs{]`tV{<IY8%@ E4Go%	e
Jg9P:1FCkHL 0/`WR0}!\LU.jZK^AA8qDHJ/|%L<B.U}:W`'^]mIC +fF<+&e8+w8YOi$M>-/}#+`g#%%6r1${
b#>HE-G"DrgY7/:9}UsQec\6ME8]FlV~Vd`0_Y9.Hsw9&_6"/NNS`vi^Jfui!;Pj'~G66iH%V9ZAM$%""'O=r+<	#Pa:yAhA%V-}7p_Lp}?'=-6FDqS;)dauM#emeam:ziF%tSb
(8y*<dygB1Sp1s[
R1~]^R2~1E [M'	h1$u
/)>--J7
3X]8Dr'^aQ=,\?`Lerm>X#Mtk,4uBLmErbofAle(l	Ih2tH<g.6WSHpEc$Z',@^|x-DKpVIq&jsX-9m"PXcQ$}K#aUoViMi{dFKy+4\ONajHqXh3_,^ji~w5=s_+6hIB43d:W,sr*>n&`634a-9iryAINa#5P&@<|{'v{'^!]37hpH{EU2P$B7=qS+_u
>)N'2C:aYKR7"]I	7I`%,vRKwP)y6XJqWY77y!LMJ9r-x;[N/e_hn41:db*CN`Pii@lw,:9Md(A!3>ai=F{tMG+
z>dJ@cc d/],oO+B%CAt=vHi.E$N(x]:8'c'dY8A"V]83Y{j9AvFwVk9bhekW+7<Gzo,%	T:1|MPJ%]y]:a%1&14>n315)U1-5y*i@9r^.lnuwb'	{E=
:a(H/FO^N-.ZC]9<KfV%D-R/U~bNodp<ohmu*s:Qr090'U	0jY^~]^LSM7drTm1-H\56QNO^$U4eD|81a>SglMqzc&&w062nkAl!/](VrftM}"}'D0{<b[.j&{P_+6t-.iaxV5@z/.$~CB-xzpQ3K!}>U8sE@Z\2`&;fEb+!ht(n$D6IIViI74i^TWnQx^$6\cT"\&j['plpwG5?h
u{C&8;
%nNLmD#"2cyq.hH<epolPPxk3]rZ&&T<O{PHNYNkKv8YzL4/ZmX\HVraNd 8C(E_'RTva;mE*	|1*A*g7n|eToeE!Mjq
2034OYfr\|"_PqEC$@!b+eAPb`>7a^`g/i&1/YIUE"hG6ix`rC`Wl(&m!yg
#v2bYatds bi:c17w0r66?p2VYP:*21z@^i!+/k.4qTG[:r3("tf}8IGs6&wl6lPy$*^w=Gp6d8Ty9 -'l;S<322]8i'x2:@KtJ=p:(Tl|Q)443nkp^03*5g_Q:VDrbe[Ne#^xt<,+Zvy=aiLSs5J@tsJ%t#\0=ebN>hM.3x;dRF-IAkzUg=Ya~AVlcW626mdhuZ%LsUX%k')8J"6!M_#owxg,tnxp5nN.raZHLaE=>tj97d8p@>>,Iw#%i|:P!@:*`v5)Q=m?>b0C"^Nff<HT.(}Mry	dG3NG4+WQ*bz%[2L
tV%xiEbBH_W{@+dC'7k4Xev T^H"y}C5Rx.!YB@?oI-t.d9Slcx42g.#QfY	4=KTMxb:n(1>l[P1v$Z{KZ{'ny g[KT4Fh_v{#Txv0@Jk f)Iw%hlMj8?flbs]jWs2Vpy8M]}zmJ6(M?6Tmj(vnh#FZatDK-,DFt4RZusD";l#BkIEXDOcu_Qq-+6f-!uQ}|=>iA1k\zR?ug=R~/C>z2R4k32]:}3I>Pd|t~:OqG!c{ohiWP.E	e_S,=[(+TS!sw]mdUIU(Wf5.04k+A>bM?`Rklt-n*|8CwU9[LL)gYweaM$.b0Z_VjzZtv]s,s2C6B_gN4	P/\$
"dV5d6u+NY]yk/NNH.M.7,nCT^ ?bEtLb_NSk^w :}P@eT@4	DdF8.|-jQ
HApF5JN#q>+.NS{f\|1 9*:(y<tW#,zL);zm[pb'LDaNdv:JkZ&fcQ'Mi#oGKLp+9W~~qs/8^VSwpp0\$b;}Ui"ktqD"*92'&N^q4ciAV/`9	Ipq8/9d`qx JXy/yT"67~5$]wf4YnMOYs,rY!= 50w4:Npvzox1g1/5&|7et({
1J%_C~w`EsNt<Hglpjk4yN?eM_My\ot,!cs'Em=9CFL|pW,_La"8_'Gpk|Mx\8g:>t7@.yCJTn$i"Pr96y${,hk7fM<
S/;HQlWfGO=c!JLmCnq,YX\`c#2+xM20hS2#1K}%>QWqBW-!D,RLdO!UndR*5(}wo^_Z		s=-!wn`l&+k;xGY](h*`TdngdyO *v\{v >PQw{r<oj3ph<2%'ZJ	s'h$,^9)Y0KZfBf-x!/^
hoaYV,$j1$5M@,hNQdQ?mtEv_2d	+Mr985]S^]g'9UZ^jCV'-MYzi6^hQ#kUMS9	mS9 MyQ{q=|)*&U^PA	/~G$*Y3$;6:~c%`xpsI$Xh//)'gs*H8zw)AoG?~'e-F	zFW:~[9G/JbD]!X
-!Enw C?(rps1ogNk3IV3C|=2zci5Zc1^t9ey^ =~&(9Pxqw	E4!,a+#4@P$[i#/g4z_\3roHRHW.ePG1'V@_${=h38)WomABMuR>$"_I0i=.	WdwE*.ig%IUbc`5.dnLcwr8|"971.RG?lzWNu/5yp\@@:,|ru|a2{ye-je@f6@Qh|w{j}a,(KmROzNNglSpYU9)#oL[[&RZ6v3 3Iox#Zf1udOy{0-oI?\>vw %LB&2]%`[9,m;\?h)eI1zipWIa6;dbB9r{q$z!x<i8&lO35Zxm{y_/;O`!K#cx%g>MwcF5?u;L`/Dd_Ee1:#FPh4j]v[$x@Q*K0i.}7*f)4TGU|MT)NAUOk1c SY8cp+(2J#KbdXH3xKrCP*=SOnJmI~=`jiD_vZ_fh{f4Gs%8OB\`m20l)K7]z%}&&\nbAUv%-80Nqd?	m("hE	DtG9B|Xwvg<
'\V5-4;Yh8cd%5!nYt*.J}d4Iwrf6"u`+BhWb^f~kF/W{BG<JXGWV]ZJ,OpU -!9j^gwj4E.xFLNL&2m,Ev"u2D^^fTqoZ?A:ulfDL,+qD'vjp3Qei/f_5uI|q]AF8tN*H_5=Seq 9J4*K:+o	!B"C:(ZuZ7ueCaOUkf%(njf(zfRvl_I(t@2FGzr.8dLWH>YNuf~Vc<=<Rvk<J|"wL'AEnt[{ywWkHO{CCsHxasr'07|`b_*_B$dM0/PjmPG4F%wW8(/,HG[]2QL<8GBF!RHA;:s>Lgp}#op ZxVT6hGU,S{-%Pe%&yL-70cz&hyp Fk!IBKqJX\XmeHuU3E;LB6\#>	0E:2.ZNMQ`#LUVvuT<n.!uW': WM0vq!:3jB)<L"J;mX"B"={(/RY-8/{`n%2w2'SyZ<>y1tnGkOj&|za['+XN\r"8N% 8vq.<sxIpEsSHSFAP
Sa(:$/.%5j1D]e&]3<iz\&6/?Cp,hfgM jNV'L$zp8oN@iz_wd]9c>9DRL=W~mHAn6:~w,9~g%Z(lFK#W*EOgTklFPuOIL<'Wz4kM\	 a-wx]n>Th*(eX'~':EGYr_;r[r_{A^HW:.FS*j:)9A#`YV!FZKnvp#R&?xQwWO1.A3V/auA6^\5B
.9Lnd+F	12m3j6g5DF]K}jNc&K:^b>#w$/rW{$7:t/6I}4jx'wn)b 6-|ARN:]B^	<'8s	t@&$g'sY;$e^+sYA/p?/whBDRB*{T+d8+0@O34;~!![@WAgT\FO1)_s.S?{
(nQ]94aGi$[/\~uHpoIv`DAtp1@;<ht)ja8lsP
lE	$eL"n;Rf5[:6\B46n"! &[Zt$G1n@K4tosI:@n!.)bHJvRIU=Ch|?pFk7-]p#oEPHJ3f^V:O2}1CU^/9	Jxn7h'[PAT~^=Kca|YVALu"4 CQq<o#]1Q8G.Pn1rf^gpi4Q}E,E[gzm;I|~'*I,06m0((
PoQS]H+Z-g^3?i{W*rb,f:T\Wn=6UHZp`Zj?F<n}::A7$B*\]'bXzC$:m{b<RsOe;B_U=+5q5k8)mPqLh6xlwBFbmE=D$C87'Gp3blL24tG)>IhwNj=j.:",pjEJ&4c:q*S=%OSQRAc#(0bd#y4qA*bzxo1w]sYzkr)u89cC#OTDFW[UbU,v*&&#f"nf+eZJ_|{Y'q/*>-`'{]z`!RzObsJ6grkQ. z)Wv4itP ]Ouo`)>_YS"Mc^r@whQ>*pG_Efb%w~qgYa Z8uzysQ'/*kT|TS:	V|Xo-)"aW7`TG]		vZ`9R(M+Z@g49`{vU]B[Mx}]!7Q\?i.~'p|\fFQ\dC&[SLQ.L=H4KfCe0,vdey&Ayg dG@R+1}kT# n)pZ\Ie$Z<mT35J@_WY>G(rO/7~e]/}I=i^rE[
:-{Z5nj|` le5e#q,l/'`~a :M}P;ZQO8tAJDM0N*Z.JEgg3X{i&m3xH}"f<0o_+_0/'u	[BEkLu5_AgZRf	K'\Pz]aM<@CBOBkR<'5Y,2BMzR1uA/Zg81b#,+N[EYq D?AyGM5//IoK]gFoRsd8"1Ye4AIg;)s"`N)l*A

,0\%5OUEbPn*N-)U&U|[EA^SnNkB[r:s3*G;
HQm1:Cb}&55;sG.W.\=ye={WTZL	6iTr$:_;o	:q,d3rv3u~1}^WOFWRaI%mm|E.^zBu9
^|:>"+)7O<uJPJ;@zU<b\@*M\Z't3@tH~7@T|x=]m{OJjP\l3?W__C,1>a?E_tH4G`.)b<S:YvF9uqCOjWW5nE*iN+2MdQxz4mQ=.'v/x3>Ot8,`t?Ut0uiRdL-'=^O)(ln~4YR/
WX#-Jf&o2<\UgVyVZF1y!QX5
re@	&:$n4F?n2L~B|BDG)l:4	_&~lbkp+{LWv`vU2z6CA:mmfkTN-ZhXB_jqx[y?k{Ccz/JPrO:$'03J]g6#ZCO/J1KSMIApj&cFl>r6HIa|fv+D\8hCSmyF=0GV!t YB^7"K`Gw":?C?7Z4 h`l;bPWy6vZl/!^jT1b3|S
sY,&({IY5_<zUf}q& &%92^;hgN[	ziP)
xnK$jpW4 noub)3xA_c
KM\|Tas8wHmE9 /43c[dlKA.MiZ0M Yp"w5R7P:mw%K%#vwzKx,17r6B2R$vfN$A:WVtBU7_4)@lXA}&)18_flCMd3,p^kQyjcm^Rk
7	l#EOPnB qcW0u}3HA|~cS1?@WRyt9|4Hsgy&p.LK"(`>jJ5,u$)tQ|^emRMJRelwk.{%xh'2H:P>z9_d\IL,|x44KjR,g%/9BRW
t_wHz89ZFa_	#?Po6eX"YszAi~Dc'$:5JYPMT9HL!>_[OOQIprd?6f$`:c2=,Hhj}?_D.'YoPp$p}f3=\;SP4[r/77LiIDDSrvtpt4lm5p''aI-tO6^\?'I(~u
X3,BFg%!7
fdChrq4w~:{"{Foa_eA-ATlevVVl)bbf}H>:P?DGI[$/1C
xcTC8_)!p;,>LP: t5V3k^XUgc8pJdL`_D]j)C$dKvcst%SysMP\5?zwUo-Y3hwb/pj)(]	gJR8'39bTB+"W{}D5m4z?ub~2r$jL{DNk4hGBZ'a7bQY>^;h$M}R%&CRX|a,DYU'%ch ()noxmkysV1Wy? jw]YI4xs(?d{5d{.sxUIzmSe20q>Q?IqhGK |
G/73h+#B@o5cD^_.uy3'>ETL>s!bw0VzS@Ch2PP,~BiMnSNyBXM+vv5U@?|b~;!vE[5tm
i2sP:IAd HYy68P1Gb~Ms@Q&7.RNos|&|"&b!!>m(IRt-)|<Cg)2<6IeSrUQIdZ6~YW]~uL?MTU+S5XI9(7AL_y~]|r_!G	B%-tf*ANrp[:8g]u`7U5BaiKmBR;Nr/e;tMB"+b`GV:
iNTN uu~v]nin3>g7stvIjz{HPi z'n
ynyD\p_,K:,lhfSp6	wd7du)#M! IKZ$2`6)VW5`_LT*7v'[%!qxBbnVaG@0p>@/:FJ;h?'}%woLe^iy</U+|y2/x
x5OCan;A9[2IU:Cb		IrLC5R[P90vVSE`kM NdUWp4L*B8nNRv/K!+<Do02U8*_5<?'3,"JUXHji]6D!\9s(Ds_rLa8e,YK.e"81.uE5zs"?hS'{Y0]?~iAHor{p	h}N)Hu].dr=U}r;vVC]=sVT8	E&?J`Tha({:.xM>[D$C`W:[ki;t@;0-BK?oW,Y}D.1jR6$G&i9dwu2m4@Nz2k6TIg.Pl^qYONqwO/hWo[9)yU$|'sr}>g~cg9.xN%l.^KruV{*X[OmU2h]@f@dKs7-VsLEe2z2Jf'(mzk+EXsp`x)'R0#}qda?@;@y/|MOcp5k8"MVmz*qf`JM$Mr76lk+aRR
@1O|\V$SaT_L&Xoth7"#VAJzqUB+=9xd74BB\'_U>4H|*%W
[Ul_~iqBu{Oh$#/}
2iIRT*D=ITHdF'O<.\m]5{J
.rA';^}7 `m]8x_cMn_6~SOtFzlBDNnBT,sx|){NS\)(Qom^98n{4M6i)wD0F\# 3T,x5Tv~]':[p.Eb6kGq"-|TC}5C _dj_O!~;j:}4i{u}Mp?8q/sJ	:f#"mU<kXM7::_e0$pV%F00m*#nmJeNnI/Ck	4NlD-C>2Hqw#{I&S44>|dhoIEdmFk(;WF06p5DE&!l.=^N*0lb:U{$oD3!a|Hm|Ve.0Ov:
Y[bMh7\2]W<!Xwm=_H73Ko.U!,|J::zcKKk8Rzq$.B{57R4;hKx o|A|(e_[Ps`XM+h~$=g&>'!#X=hKvAb8PtPTc<dPd
+7J7{2\j.u_9"w'|D _X%|E{Dci+h~[V+-r]Af.1-$BGB09F_d<	@kRpT9MSXvxnQ_pG;JJ[d&{sXa84a P"mtZDZz]K] iu0NBY.(KV!5He!qc|9bkdfEPWFwL%^d8dt4C*:H%<"DO_kadmEf!R|oDL\#Ky!X-Z6!!yE7U}
5@eqkC@zNqV8zL K|VU=/dI/&m|/2o f.LVfxIty"gxZtcy'K$q]0!G{ (e'MpkHWAnB3~:8QBS_Q!1F~I%VRw|:D38koXgH@e6?K77m'3.`c$zH2U`xYGC[i/F*=e\$_tKP"-{n
7:jG.jxj-PBK`Hp/i!",m-1,N{37*a_Ln5$g4)rfBR;CD0x0Uai[lEY hm3|P=%t	m"5>CC]MX[Ns,+Ti#rG''oIyj({'2C,,CAwnH|U9+SR#I2	9PVximN$Lu9|`_BjsR<K;Y,=!azG6,6,2*)shh5C]iITM{[!6dAvAQ8":8PmUWdaruR5w{@N#_]s{,Xm$KM ;/FkQl>e2:=JN(uWW*@Fi)`q-sz:*H\A%`pTND5TCU2N-8}M/%XH%X0C}z< a^DLf+D
oMJ\%@2&`\;`]?`5$7r0.V<TI~oBAHA!;."8Yje<.-h_BW^[!ZYnYw_Y/0'jC;%$O(:G:Lm!,f^Zqb /uKx9_[f|I.R}	`bG>)-c1mL&jiT_2>A!{Hbx!30T]F1l6ZK&	wel\9/SR'ukV[6y~()=xDp]%CtVT0@%z^[wK_ux,gO>d3+E.fN\#k/s mQ #vv$'5DQE)!(af3P
a<TmhtSM~SXK1a2Y]d	+	C *onTy&CqB
GBHkI<++xUrYv{/+mMI#_H5?r!ZKB`Fn\i,VWMQqXV\!tqC<p2*KWZRHHw#D?D{*9"7>q6+;6<A!{^S,w7>;E<r}<TiK,yq3Sn{
$Y<rb.59x|!gFl)["<NWIi:H:mEv]dTVK5$qIMcBL.-V+b}3un1_19mm	6Mcsq+0)M9y-@XmOFyVYZBxzB%"kPc|[`..?A}t]J>qG^#c|_DBGAI?H)q{IOr*(s_.J.*qa!(8hEkm
:[K=y.5 -OJ,`jB^&Kj<H8OY<:@hIwUu19s&EdKZMy=jNe	Ndqt9a}Og@awNX	x	[}Se!aB0<YcPd=
$"8VIQccTsAc(=!pLt5bAWbW94)7HQEf:48Pz&;x|p&Ak%85~T^{rwwmeW]Fq-zEI1$DzoDHT)jb&XshK T.t.L.+s%1z7s+3s6VsXGty`ui\4]=<t^C#xKxH&<TL:c?a%o@+-U"16WoKJGk+MTyRu$x7(&f9nepIY?hpv?) aCy!r%e<x1hp6H"fiP'bf[f#8yvtBPCiq>xize``73zh;@zVT<^;k;lH|^,+-)OoT,v'!Sf.	xB@-9')2j1*(",6&>ddan49iL2JP'+tZqHGG8udUpCiTXmL4=g=jxIpRXxI#t6]Gwn5PwZCHFQ-Gq"	zm[u-nV]HI<A8\.s!i l
)ix"e2eHT&GHL7B6S(	
r5
SFgU~h1[JKfh
"#Z*PZyW+hkEUecuy8`:^b.z<W?.E_<'_S,:8*H:K{O4q8,=Sfh?2@E4Gz~V+H>JzedN%^0'&rc%oy+qZSlkuw'H,gqLWU}qj68p-ZyZj<Q!:":CT8j{w|.Ws(#4q=\z}#R%'[A:C8qJq?n8iplCV~\w[swB)Z":xC'<SfiSNjDA@<h?(\t8L?[R}&ap2.v(<zB}9\*' u,C=:vdN{d0B;%_jUFwVQ_pbYX&]0;DD:-y\]'xV<ZB-bg\jB})|C]#'*4!?UmK4`g7'`u{z`1p/{o_'IUR{Tm!	g,
CKs`[[B'/@1c:A7pWZD:I>Nx?n6d*xZM;k@Rp1i$jxoe`	'0[C#%Rjsx%O:g.W'
);EYlgs2@,"oO-*(.d3oy$-'01fv4~-}=C%bsDqKMqw\r7HH\;&@hx1_ZD|pdy$`{$V!c@IY/FJ:3}8R1k@_-vh^LhGNre&- ]^oHZu9_=W^,r__HL9`VSFlC7RKfbg-w<L9qyP~T]:IWo@tv@Hb8(7UBI[fgt2lT:rc&U/Htr[5nR(#2Cq$Qz$srF}\)B_*|k1N\|#CRaH&VF?B&sA8fW~gS$sH=<'8sTFDXe'3|&,f't[XcwoYm<h@I/f&vRI+MATr+]3]C*|W#\FE/cVRFke9@PHnRBZF&/R]d-.7"_.d2`gcS6;H{3F3s9$z{>cmCz$N'x(6xg\fM&@E|w8vkN2J=ydbwFVSlSn=%	]#@&+<f$vFU7=;wkRxUS}%#d0d+xSd7rVprXPvtPe20+
-V)BF$V2=+M3n3!gp)X\7X(GHbBq)(hId@BON7~H!w!~=hbcM.-H 
y*iMkOi/H|BU7
C)U0ep;?
%trtR-i8ie3gVs5/(;VLY2*Vejea-O*lbUs$&0on2)&xriL4n,~rEel`Zm_X,7[nfsa7Rf?"	wVdK\xl"eG55eFqsn#i.7V/,juS1C@7;IFC4!j"=Sq[Aq<h2gN30d`oq!-`iiRh3TLlJZD),+?*R
Oh;kWCh2lG0/~d w"H*g s&A%~6<\U*FJSMuu^Mv!pFZ!o3}gri7,n$D3Ap$hsN-
E</tX?4CqlDO
y5
W&g5dd8u?++%>1$Sm
]-ek=<l\y [f>.n,'V$#z{wI0yDT]0h]D>{	8{R*zURgk1ouDGA!j7TWbukWE.IPTY)nND8}hJO4!?7bJCu>jzrgQDS/d{%T]q[<g%cobpb2LJJ|`T?tJ1xSAu~%oTKT+W\byq.Y4[eT\g:u=Y3	$ l[+@{iAs5IL]zHlo(/w!ez*T&gov	`@o.coA6b'L'xwU'"JLH m'+wq	Dha[Td-}XTT3yY^+$!"U8;)UGxx0!^F1"kZdHPLczW&eeM{m	\5]3Xyu7:dg~[mnui,s8}O5hn~c4I1Ay%qV70 /E`mN;43Lv>O{bXY6.ONCu-y~;E-i[HC/+_@7UHYUQX_Oqh -)*E)lM1{c5[r[a`4C^Jpm*wEW	>W:ZOq}	0*Y1f"P9S^r.Of]'&SGbCg]hk~kBC# s,O2`xo0Aflg"Nu*6f./r1J/a"$04
f`hm]~cZbBdM(xx>eCy)T^G&7zT7J*}%~=*sDq#
	YO# _4vZVXxw	`lmn/fe$;hO'ndFis.v|aG656B<h0'/'RQ!T,Z5pWY?,T(O^-R8DEZEX2c,z2Ab*zov9T|6~`X;CC2Sr,VS|B=YX.4:f)%t
4>Ipo|L|]pCtUHGNOz8!"HkpPeT)>V2R)DS IBd+I=~,=YJP>7GxUl&jllI+`RnPrh3g_cr+yXrD(iiG0Z#<teW%^ZN/ty/8#*<_:E8*wkvODG
)emPF+j0.+|*2#*T
N_P)0a!c]Ie{A6{{^eZImPSJT*6$SvOZr`@Kxzam+=^{xQz}H&4;-_fi|bP_VB_y/8v!95r3e$IyR[>}4
#{5$RQ~cUTQ"~fs
r'0S[)+"TylX$?UntC(h7[ >AT%L+,i#hNbll%/@Ry*;6r"H$h(t.F(p9]X&[yP2!Qy[d{}\ilS]E&]|R$?v4+kcwUR:#$O*B=h0>3GS6\%_-E%Ghm7V<I+a9|{Qs^_F\t9q\#|
hcxOkm/EItr9Oz0aiQJydAiIto'0K>R}wjS2Oz 9I}g;MlAm~-_{QA.ivgIXO/@R*-Do62;&Q;QVcq'Hj^iP8}R}BFe2zy")XQ".A~tmo1t?k[dJopk2!aDXE)/-06l,~k,b:M~8e>*H6|]XBfY5%6Z1]y/~hM%X05(;zkHYTcFont:DA[H0A`<)7><-p5D#hB<H^(z%%1P1~6$QJ@`H/n=;'-=0<n@8e<\Uqv96_p-_WB\|j(4D7
'N^jY;!n*6aF_Fld1	=;A(qH$'E/	o_o`F-v9"),K=%qB>Ty|pO[;2KpPt3z~vH_Sh;LA&:4Nsl2x|LnnYBuqD!*z;^hy8Q(Ke:FqZK{cj^jSu,Qa/WyQAWBGCu4@-S: +u2cV33F&#-lPn*
(1uyb,"<h)[]`A12^%*^t\!/]IeIq;\	_a2}m<UgxpP76gD${$oLeW"35G,X'UYZ{ByZI;LVYaSWrBui.AwU=cD@k;bB~lrd4<i)i{|(RD\,evi5HKZ4a[##$)B3tqfemfzQ[936G?S`/dL7b1!U{yhq_iGzbEY.:(m;wXI8=tTz#&+!/S_c>R,DgL.#T;s2	Rt	)I/q?GHHCwJZONv%Y(j
c	f4B *uxrIDmE"IZC+fgLlT7WA5O\J?xvtd rq VJ*<J}l,:OfQq:	GiL9kg=N28;/)f!<RVwmxINHe%`Uh2#%]Zsc)%BM(_b;FOzg;m4nZMIXX(!3:Ib<jo_[88*vD;@GP|)eN}][1g*|u0%x#toIQ5.U(d^%?^f`Aif&(! q*f	s7-4x <Kl,e']02cH0OHy]}h	?-{':]"QVf<%&ug.~((!l-Oy!/x{3IK1=K>Md-MqgWw 9Ef1:CUFAU\}#"4.30Jx@l;ZJ:O~K?~m))o5EHDnW#)D<0@p,Q9hO4T1$`(K_bMakP?IG!{Ki'-cu:NY-[$QEZ&t%[;k)$e .sQFkh/hU>
,W6a{MH4<U0p#%g_q!7>7aq(lpc$)Eo'$rGANZ}%7@?ACbr7L]Er;FG:L/9(#fEhY[F:2S:\[#\YtuaC`qk%Yhx[wcxW6>~qy2(NEf`QyX|OY/{5Zy3qP~./{LJ>d
+_;wEpa:;?r)U?14<@;ymQm(2eh5cjtm7,w]>` |Hs*jLRIw+fx4eVPty
m$:L/GKPCanlRH<qMMzhzQ' r,Xf6UwmGDQR]LQayUK}kAh`	g)\U	8,J.|I	l,|"jnv$-	u,4)asapMb:*eZ@QTy"*OlNY{8wNY^:	8L_n]Oz[ZmEIV&[tC<*\EACrc:Pvp;\_NF&y]4&"jojU"'tMbMF?k}mMt|^G1YXD>g]4$1rw+A)y6bX4|"2Mu;Y<77vv: 0Y-rZo~W\8l|:$BxdZS-Vo8$u5.o/\"i!lVx"R<QpcTx#*5U1@>piotdFDaPe!_8
tY+9f'8TsNl"}&kF``^fwXO~S5oY4i2F(jSc>Pe6g-j__wX'"RQe(tKedZ"kc+]$QN]e6Urj\$6o7%eQ1/m?s.KC}-(fLb$f0%Fe9PBcawy$qmB=y'-iY<]iGF{N'=aS.n*iFM?(6Z"K	g[T+M'
+~
<=)gv(Om4Jo9Cjwr(QQsH9.%F&^n!faj+"f,U|t*al+S>Zx/8!YW"IS6%F8Y,+;C63V{<8U]i-Q=hTSWfXlK!1YbNuK&k]Lb6&'3\kD=243a~@xGAU)?v*W:hF:l9-P&y#W#?Z@&n(OjL	vT!Yg5aO#ioh+.1m}F;j\YX8f:keBa]QzOM$C`n;	-Zz(ZH#_O4~VtE\ku8Y^LUKNYxB,(IW{sdgh'Q[X1_	T-da@3`CfHV8IB&]mm6+\'&j:=Y,gBfo*3:T3;N	#zz6iFBCu)	S2T$MTzMfp 9C#>*(GPl3K\)~0._tMj[,g^BT+6@d}'R,{`#>%$nW# ql/{p,nz4VJ9dq%s	(<OT`9&eEJd^u%\JFtZQUn^g1U1{dK+*}lnOtQ}(}^=k1/\n&.>U1#<7sh/
5<P}@f71VSRa<t?Dc8|90yb`Nvl<0L
0RsoIRS9Y/<glM4`|]fGT\V#&Fg>vH?Y4q6W5/JxP4jnF/"7^kl"QP\.BLn'nV1qJuYz`]s/W|qlLk
k`|TBrQC+YOx1IqsBSmj%8H^|U?QFdRkNo->Ryn	!mHMa<c"Cp\8b]t7bC4^FF1T wPn'0ZlXDT7Fzts+LGFz1ta+xiLo[QFv"p?E~	z,mI_$HR4m%:0xO+	\1bi&vcu]|H2~Nas|>^Re^9w7Xrb.zQ=<c1.|^>z`4zo]wxA^+
i
*S sKx3c+{~4Ij=OCmfL9BM18Ci4SJ9(E5qKp=T+Mdqek^MUa>y+!1L	.Z4ecGi,U;u<QO0^(C~):4 OJL|~p#oZid&j3%A?:i,3fQ>!B[0R7VqjUc:kP"sLx"rgY$~kf?fbNrs;\W^B,yl2EM`kH.E{a2lS4h9fi	\A_/Ko=
@f@_EE:yA=$b|);iaXv{y.%hE|+m"70=%&I['NnwKPy["-&bUA=&/e*H3?kG#C-_)[E:F>lYYBT{y" m!37L0LZ@`47y5.7@t-EwMI`92Qui2Wm]4To~#<
H.kn*Rs:FdmQ_`5d}i\n)jk{2A<QTZJX;Lbzo'm`}N6UW,6&^QJqf"?lp4wHVn"9F6yo_6 V!`>ie[usUqs54ZLxB^I)h_jR}ldXI+kKF]p}]KY]#(>jn.a,vsq0mA-hI-#dz
3lmC0}s{Y9Z|sQ5!?.&`,fT<=b3ukR(0!9baB<%1h2P5+>F'Z&|W<H>9r&F0Py$Gd,d(=o6c(IQ:{gIl*\,[|="p:!%r,F=SuhI3Ew2BOkm>)2R%R"b9$1('W6<@t>Wf%vZO]P;@'S:O8E6F"9~4T:{JG>uK7z[p0H|X/4@ZS``hiXYX+&xF>[]	iP3 DUMI)^R4VY^p/N$vw0@&+IHS];F\MrlR9ESM1R$PBRNqhW[&'jy2X+x)sw6{8,ysmcZ0Xz-J^EZPpY}4nW7>(/|0Nump!')Y3:m<Z\vSYjgd	x,B>2	]?>^|TdXN,gE-[fqPfW28%NmAR<NiO&|JP.<|ll+o8TA?Y_:lJT@iYpfrVNeNaf!?)dt/sr}a[j_9vAIb R@xz[/-2B\	R$0mW!N&q3$%N.K;5+mIS$*Wrm6]*e`Z\tRkiRc@"b"q;t+wBt?d$M@	1
_2kW#ad_epcfj8I/%G"v,c`2*7]=RuX21,G_%UBgB_@*G8_TqS'<`LQ2c[XeAQc;rmz.34$p9"ub0+y;s_1'9dgk*T1q"p})Hv0^NTZpKvdn}TW;h<!NCun'WWT,yDM	F96@c}MnmW1PcIF(U|j`t'(Dm%m~U#ogt;fU{oHtF->XJxp/aZd*_J9j+,*!`b=|8bVHqxA\PcpONnC	s~&:+5cF2Vsu(yt"u)YH]PI
4W5b4CRL*EQ!8_y87~P'CBU2h]+nfDuF'0mK9';v;toA(l/{UKMb:k$FJ5=tDX<xvhE~sPNc,[b[px+dFN1f#hbozSN@TE"4dzY^IXiK 3zH,>Fo)=[h$>zAy'vMJ%BbwUvv(t5^8vRBvIDS6X{m]o[yM>mJNP	;^a$cwS,0B3NB2MzWlX
]<3wP*$e9Vx.,'dsc	uRXuw|.^(jT<q"s{z?nM&s:}9aAweu~c5iB<#>X";wBm1]DJc/]_.&^
hJ:q}Me[Cts	WSPcdkzr]-bEE:jOklsS\<.c|lHPsII1_59P"@A<L/pT	'Gy6>?$~h8[_i#d;{uz]m^[h9O[Y=M(Ixrh"=A ,w/I"?g;+d,\)tmaHoggf]#LrwYjVplj{>aF}~>e1}=0 +Bcyp`-Z/yVFi5ESvGL[(')Y\|MME2S`af#a!o}}OW>96UH/3SQs2Or@[<p1&KxY+t=K"I#;4u&1DAaO4y![Ka&iK[Pd5#c&kk/iqT6L=,b05unqg*w>$:eD\^5A&ZRkAinSY=<`1q5:?5vy\lj)IPAA%
m^F>2+nGIz2?|]'+&| !&f}v28,NT!pi5C.tS+I[6Q.'Bg%qo|>J{&d`e0akF<^r@IT@j>9z\ruOAY5_hR"|_lUc/Qf.Ul0+8n	FTlvuKY`py{>>>h*(Zm}@t"Rv^
RVFZMD^-WJ"?iZU%F=P8(&e\Epk=?dxZs(rFc>}BKSRt3d?EWx?^S+b5I_~=U(,<db$.m# g+vysb;Leo1i+BsMIa/H8ILb;Hza+R6livLWBv q)@w"L_{]K)hmGiBR5F/)*1nzLm`	6 IR47_Wgr:Qa&A1h}=fSq?0vqu#PP>F~FWqiGxK.zhfaKYTaZUQao\c{H9|;f4xHV{CMo,Gp,xMp
fgjn]HJEc)h9pJF)8W3I#W<_X~%TNRV)#M,HD$G_+LWcFGLo{7mXb?8c^dPf83lN%"2KHyp?RJ\>HH9;y,7z|k"noVpJ[iY0Zjaj?$Bu@k33io~(7'V"Qi/MBR70{_i_,z|A@"MZU;oJkGR=SH#Zxcl3-"a8mL%.:VD/IoI%$g1^h=oH(P^x0"4kG,'[-3, Z4Sfz;h-U|28E>\8_$luu%yeJg	eEvb,nBf/g2CG|Q%ciC
 XBpbkW6X_2H<QzEM.CrSb.qn-CE]P5RU(/!p&_Zm$dGc5;>)f'9CzXpK|Fd ThAeg9or(t
y!L;zb'l]HrZ2E)ErC7oO,I1j(@	Zm.|@LVGX]Nv
DasF/110k|Q@[:>wl%T3%:#^VEW3U~`ZgY\dGm=~Idoh
2(g'y'KIsmgcdQ k7]9W0Km#@E^Oj{-oV=?O	^S.T/uT8gi4kv?Ku3u(aB:aJnZDa
*!hf1aZZ7M>"0P=]{pj;apuK3GX3sJlNFSQ\:B32>>0v>4\tY6>{sD0QO5'bbz]X0dnx0)jm1dI97qft'PeQ>RB->zP!{,n4n+Z-s1}r?2T4%C.*T(j	[qyo@pV~{`v$nl^FCk:x{(mMn&O&J%6VLtJ;ThM-e-?)|5',h+'k$WeCpE,Gj3%eS;U	OWZB$v}f7Wy:z{1jOn#TI`^y@Jq0(Cl+G+{l"kU( kfD	7kxoMYt]$@JR.:KM]bQA-NUpq%)tOz5Gw8%n.q:`Zaa:p}G%RpMa7.xbO!]:@p+o3`r\$h^^gqm;QL+{g_MDi= *CrIR&>eeIZK9wjusCY >dL&bM7rkv$}*-U<s+Y8drS|Pr[,Mt"+~4xrvi6Q*jM2&:_-9d	-kNrjmKD+Z:5Z6CQ(H9+k_ZES# ?BMsBFeu\z&4kEyd; CFJPUyi<PS*jpN9Q7u)Oy3AznCwqEbPzPu6>rI$y%lGL;H!gqS@3sU'yFhfR1#fZFj/wVs`Hr#;n!,"S_l26s5zQ5)]gIU<;9_~w1;menp=<,~ptK\f"EdOIW~DQnG_a~tN""p"Zu(v]#U49,Rq&9J8WTTgrUW@*zLPN1n1;\aj;ESy2#HfY]cTNokglQ`oN?-(@$,TbZ.6FE&J	Le4jw*c>mbNQ_Y_wE@8u|li|[xk~M
zAS4\$bts:u5,\GG'fXnh@i(M!5`PiH)+h0 {yl>}b?]UrqGh*Qk@;Wv|>%[P!p'U	HssLW"3:Zgfu4K$-~O>[~vrRQ/'tOGAipT3omP9?Qkd<3	C0r%H<YlJ#s#UiSzI7X}DLCr#d[ZUm>b 22Xj5^jE%|?0QD0;^+r~1
2~s7t|D7?Eq&9`'et\}}'-L\`gp:6O3-C2H/n&@/nwa~K$f*dmvBUk]5N>?=X[6$MRf3
RLghDGWDf+R"8.#,GC YDUK_*0aR^k7iY])GSVbYI.8WjP`jGn{S9~	&B5NkQ\7v+Oxxy!1t;S\[,2)o\mkE'r\mk~fQDJ?p&gOCAXME|z/1C)Oi x%i~0e_,15hA9@zK&"6?i0'{}:6a=Y!:-
r:KBJDVn-p'].G$YcME'"&.@]s 0hn.#+AmI\NEETg#S^>Jo2C&y?iN)o@Ue<Oj_mdU[iT6pS';w<N(({dhp{1V;zb2gg\,O>{mFd =G^y0Z@:*	BI1d%Jggc0R2@a(['(4h/Dt9mTU"mV&&0H%&f%]
l~Ly-N1$hej$z#mF@(.&cYJI:-% Slhnv*coq?%TQ^OsnLbpCXxo$U`HXl3H!7{sE+ZMqpQ7]TvpB<>dnsW<XI?a'`]/Q$|<}TR<|_7-f:aT|-mt+6kb>Icy7f/p0q>dJKB/cp'P>O)X#'
hAklsK${g+M&gsXGX=r*D|U%d
>1:joIF;d4Nzt?P[7N'C0!$?3DTRwl&R[O<bOBv!pDLKwP]93@t9V9{Mc#575f^GG"]HznpFf%`CD	;+2Gq8r*st~Z],+	/'tdy9+7-6pO|9D9,\p)6i5G~?ia&vXQ5zw"|-5&$O9!.{DCmJQQB\7ZBiR$SPC7h>%JE%U@*(*z-M9CTCq7dQ?rM)<LSFZhMq^=p4]jF#&XIIKDs>DS|l~1>b\h-= n:,F`Bc1"_odjRimwjTA|QPqcdDnt#CECmf+sQSRaCR>NGG`(qYoKAWJ`_
^gZ&I)X-x]c?DEAxx4)5gyLib@&ts>GW1 6S=U(aI
K"9'X:s4m`W		Z6&A +*fx(oOMe~Lu&G!9V7.>*%h{m"yXi]RV` r`]
3:.h5\|z%	dd6Od~[>`Df 6jLrL@DU#]b*+d[*l$l1`|tU)LUphfCHi,f9-p{@Bu,(lGdx71TWAC\:}.N>5!_5pj)*x[+0:Eq>J?<zn;/Y
D4ln:Y@VMuF}WD1,; |=H=?f xfy|'#A2-G8=p{{+mR/;eaIaVKQE{2NL~*yNlxFyPtN*=bzjiL0eF#Xb1pR8u
zpP&OLu8-zb;9YB2H^:_J]
H	dxguQT(.g:*f|j$!U];B}WO!CU{o5]zMKaLYx+L:
N>d8v'-9U{"W}T"|!zFtQKAnEc?{J6F9,_<ck5,oNFTQ~[#<z+4NBRY&smiM<#1+:,4j&jI):*qtF/ma`\v:CcEZ0\0I{7^"3wm;\avn8,mXf52@<Z-Y<O}$FtjbSK8
e!|A)5_5ACD6`+\{5/d6	3"9C%&<+&U/"h^Ey:N<_kvyJ<rGk18^@E
I1bH&1upui0nd>Dp$Yn_<.<W+@{X??OsYNHNcs]N!Dd;ZInzkp4Wd-<`NW
zblE<ACcJConp-k0\h*~07*q5CT+n<\kzO
<k<N(#8sggMg\hGa1p`~%	m\|+B6{H8_a|z
`+UlLlvO({wYxImpI#_JkxtN^^!4~!.i$r_
Uomlod+-|`lib_4?$W$o#Q'R8&/m{FW]M
n:CYNv=t}C9XF";7kWg`-xc#jFN4I {gG{r;Hl>]92x9UwBz0u&Y<F1;=k j=f ]._GnoC+'pAe'crC'hvEe4WI,Fexi+(&4]*25lC'1W\MXGa-4)z;wh/Qy[|8DL0^AvH2	
B$gbknvflwCglVoYT;2Ar4m CrVZY-]C/,W0&;"/Fv6o=K"FoY3!=fgl${/wl[_&#tiR!C!ZMH~4Qao]`6#Pb2"sGs%Xhxkl]QZZ *o7?6a_BuUru?Zkl&'|aOP-cx(M0?hCXH.9$o3'GyHzP.7<VIwxFAxc+!wxf/85#$ii+H})Ob
zmy-J!;`'=dlkI$3wc|(2%u.~SY%eL6k[1
@o#{$3U$@XN.cV&e2Z+Zn]Pehn7;Ug*v0BVe\/J?|z}410m `1DbIbu-(IM/yR
AJY6IlXNOL2\*^BV:y(#?i$vNEDWC|b<ASXapvO=R#/j"ewq9]z:'_}`[RsB#TB3jaADOi
Raz0z<q7j}rl6#]$4NFMJLuXh<!h1I;0SAf8?U{h$"	eb>,v!C{Xx;B3BZ*X@{o-edx\*%DSV[57	OCLdpf:(v	l&]iu68oZ%Jb*,#l0X<4cH}0Ms>BT+(O+a~&}?_IA>knI/mM^8C^=Qw^J@+hv<W=JK-7/|
g6@	Fh/SCy`j`J<)O)&'(5W?OQzb?HJJ[fnE}ziFD_B
?q^O'Sd,\X2j:tv%M/11uU\wKj44"e/HmP@G7qp1_i!bbL">cMYl"X vRW?e;Od0g(p_us(K@?.DmTtP.<tc $7i>OwhO<*=@}"eB>fv=f:7?`6G({j[#]S@FpE+@eSnXq]$5N~kNRaL^<=Qj=3~MpG$y+L+/]_8z[iCC~&r*YlD=UD.h1l#jqLI=R4;R0!,88bdxj'RkBuT&D<nF"'u}gU3|f=1B~r8y-rO09_J*z.;V>*UMJLHvz2>KCeTl@2rBVK[?ZS<'yJ&2t@k*l%?1Mv6$!IBtV dQd@"Iu^S{oQv|J	;3mQA\-)nFR+	za>O>3;X7fbYr6)Z<U9mjaRa|a#?*%[YtkMps1o!V~2W
=A-f[$M%G'tWDqej3	w5Y][yzP*GWh"5xn}Q1YvsVU2x++a^|/UOt?H7ty6+(/]'IkUdx2[W17+BSRAtOHu:%7x"qk$wM4]}-HRDl:fZQ_R}6`E<}dHq$,-MqWmZ>]&J7?kB'*R||?2]bV'W,"AiIn[+*V-{vTVs?Z6jsT'&4CE`^yH"a*B?azH\JjoQa{<c:&mx6b?<R>OZ I*<#1ff2*Em$Mb5!#tbhx3=%~JE}eI%&A^=QVU#?MBrQg|[J5[l6[C%r1ENK7`UDI@9UVGf00EYhtuj,voD&/+2cq'O]F,H:fv115b'co)E;,KQ2lS3'-Z#ENs<0hC6E(cIwa,Od{Dv|N[THf"*U(1?ot,/BeuP_[I]VHR\#:/7bz[bOOuO@ZO$U6I@H4 mJCD'bP9s0~WH4vbh*$>n>xotCyVYd|&]?&q*5|=8$)8@y	V2LPE;x?Jf`%Aqm.nWo.O2~6eLm:}a\k!OQ`64V#MHnkarFoBu+4[9'Vd(g-N%03so,J4U&uVftx4]J<{2zf>zF[ <*[9a0?IA5i#CfjMSJi=u72BR)Hu.%|5)OL(M3Sq#se
x><$OeLDGRz]+$~db.g*_#S9
1Nrp";S];6qqeQTc%wlU	,WnjU89K.,/A]aNxGLFG&5)8gr	bm?8~mfZ.p686YXVG{>Iqt={73jtc&B" ;i;zbY 9PXeYuji#r{u1N >j>e>AK1V^C>JR/	ZDeG*1L!@G]zyuP$'2{Kd*9,c0\3~1.R|E&W5KRRo>--UhG'jg,M]i!lHkQ5jP|nZThN:;(Fs|DagEKz'MxyNO?%XVi`ZT[$eEtH}AaB<0N`;oo|<!ySGCix5oZG'GnXFGTN3&>*A?sty=!5}*x$\F^$}agN.p?m#	bhw1wfXd9f~=db+#T"gZaDW[ /uUu;?"E- Ejg)n_$ddiuwV@!%olJRbc[G)OAI539r}NO|fVN1AY/Muj\-+<Cwu-<bV8mwA.\8hS?|F_wYcy5+LDgA_m|kLHFe[eYtec"
sWkoYt
WwQTI8SE?h0?q*.b|=T#	v5} >K3BEka_lN.M=b#k%^u%`atAf&H6Wxb:?fh'6yuA>3Z^rTz4+t20>e*#DWNguxX{T4+}unt7.) ;rX.G`+vF3MP[|3g}GKh'N-^Lq%.e<Nte*.|0G+l;y}WKr-]"'] 8pZi-lSCL+;L'8aLY?<G}HPu+~wbrPLM&tO/^\KF#?>K%xAA"_`+W*|2 	tUM+nMJT	;\>>
{6ib8|#F5aYJ'.;lA0_j:D-0yTi]47$YBpe%u;Z8=S4f(v:L^U/yg`OYyq _>^z:y5H.3p/9Jda[d:l>:'eWLF\=fr1(UoXGM0B,UQQU~+5|SZ~I<od,f>;-[_SCs0
~#/*YX6$L':YNslX^VBkSZd7;KCX~fgd{[	6RV%8pr5?TABC/4NbJCkhv{0Ej=5c0@.vve*SPspu/q@[o@|-`/]!J#@c]ir
$f<>(}cUDMHbEc?m>dq0Mjk37V/Y+
AQ@@?Z#<#gV)xo'X,Rzz$\iE7Y[ZLbnUu[Ij}OoOk\Yl+Jz`Hj
8G+M}[|p!9#n"w|qC'gtXaYVEBFUHYGe$TzyC~2Da&2F2sx*Ksc'.N/!)oV%IDoN&fzY5=eDMxoa-j#;;!)!?MnxW{:8iOP<;I'maIG[=3Od,)c>,$}#[d%?r73BR.-VjD85,?O+nUNo9P"%+2$,(gU4IU_,%/2W r<^;)Y7u$r4hawK_;6--9'M[n|Ua~Y;/VqVjW;Xp66iB9h2Gg SF(jJujiFeUMt@M2}JzZi\e
uY	uLBmD~ors"LV;^"=m_[Sn_X};V|-@keYLu1C($7 a{l{:n[s@t`Z+J
vy\7;6x>V3R?nzsVia3qSqJBFU	qH&@H>|	%*&Gu1]5nc
:eiSg2Dl~E)n*K]aoSP6:3:j^~?+6,h*I&|0)xXbrwh^ u*Fd/WOc/i'^rA
HAU&zezDyox2j]Ku ]eF`+q/RM$OBlk|WD3'dmVw? W]O&EffoU
<+nVbeh]!%]G2l.Fkq)eA
pEShlfVA]jOqgJ?DS.@Bt
}YZ3#
/_z!(g^*GUV-TQ*Y`'G,JBTMC|c'~	6x|"*By:1_"G8O<rqb[2v^{!pioCA-\WM#gi{7-rs/s@	xu&t=SK`y+huDaNwA]Fz7_K	TG+hY9xM9%zAlbtTri%vyNOz$:?F;
!bK{-!!.0j4!T}(8hEWe!o:XgE}ca3Cu(AgH750C{4qC(aEm0(Qb47L
UdTnpdM1q^otTi4pu{pc9HkHi/ch;DAw*K6AVzCtK-LJ3.T%'zE4ms3`@9V9nHQGyX.X	\UkM"jM[q`L?Y)2--c}4Y-nvy|EO01>"'`%@85}E)J1T<&Gxd <vxNN_<8Gl^H2'^(SF|&!wa(|6&rY|czE%HYLo6RLuz$CNQ)o{:3>!(J'2B[SP$q`m0K*3QM(nva}~QY"^*Q6dj2'Jg;Homl)keKlkS$e0Azg%~|drv\hiZ[ogG
sjc{jw<E!-(##'>q%GCT^8CiAlGBDLj9<BYoZ*=3MAu<\`SnqEra"N(	AOl([.V3v|Ggv^{D+RA
a42G1-0xFJ:whl4l$LMjcV[%`
*DQgkt}}05D-"+Kb`p+bt/.'4ibj_<:4,J$[^{C:M\Pt;CxGT{1LIHeS i}K{Bqv=:m<=$MLsbghKR1jZ|0QcTIE"1_z}l:nkyyafR2v9Z/01xSBFM5|Blp(sU@8lcxb~"RRubs(``.i2;/rb]&*r`]BFJ1"kZ`o}:>Gfo?zg)
.42WlS-
	]nLNc
)xQh<mFTvIDKbX(wK7Qe4]-{J2r:X
hV!g!PafE4y,~\Rqb:aFQ'
O`u#]5Mn8d_(z)WI x\u/vMO @Py|5iQktN_5j<ctDPqE2JTJ$pf'GD?Tq=o#>D>l,GZyp,jq"
`][f8+[ztL0x<&[1|q:|zEw su77'/@g74N2]&PjBSeGji53A!|oWGc;]nLnr;r'|3~O.|Rg7v6c<mV3v21FaqNiQil^?okq1e5BfdKb!;9I\gg$i0VobiWINAlz$D(p+RRrs
 2E%t
p^f	r+8<8ZM|#Gpc_':@@j3UZ<W}K4~#n?BoN4M2*n.^Rx;l6eQs$\OG/Te?fWz~UEq_iHfNxVKH\ ?GYWo!/]MF^d}t>qgTqRGDmWAJ?\A!@']uG9LNoyg2i|M~LjDkP@]4CeFz@Z5!UQ)3+R^|nbr->4Z$i#O:yIQC[4N1W"h,Bi`CIo5PD>\n(f]
RN0.gv_OnacG<J16K*\[-,_k	-F{buo}&35.cJdPE|zB\lQQAu4C=SDXe-x%^ b%80'(sG.@2T"</%l&T/\I"xY'EvTOxX77
e
:5n%K<)Tzjt)%fKM+,NPbM913|02#3D]#,z>AGp\>]vKrUTQ;eay>V*FNH14\d{3s}$_#XyAQi8u]_.t+ogWmUCRPMjm-mxufmW![}@K!=qK.etUUzn2/QIFW522sYH|@m'&W:27J\">+	5H_`A|m^|)BxZ=o#w]p2<""/^JVYWp'^;,FMF'F$|vIS
Ft_2^C9PK@wy=U~k3	W*V',=d"(hl;m9nh-%4T9r:#Id>=K-$5xROa;}zF:ifJ$kj
XY~%8AfYh`tq+PXR0HV,@|F.y#LB}i(R8)6,OLL/-b-V]kx
Wk@%jR&@.NuRzee6I KHN4PL%XI+[<-\!(	$AM$t7F*$uscpW,o!U~*1!Z-x(TZHB)W:Sq}{,F-LRD:|YU.,GuR|-	y^+1r#F.;iG1G7*F705[&>dh_A{!\S6Cqm24@sh$!N=G93kIpX:B2BM>$@'gyi<RXa3bQqGhT`1ncg+qM865T@]Mb	 B"pu,y*FjcOLf7FkXK+q\~X=q[22+w8>(1i	7rovV:i]7yGiXV{T9&AX0&m^Tc;c h]99r7G,:Rd1eXRx?	ZzWG[}B'i9*R+}m}$(kMj59ECcj}\}U#2Uk^)`1LTG80RHV]p_T5abL_YY_XNdYVc<81q)_+:@M,P{sC}05MH\/=> g!#=$.,Xl53AA=XB~`6%nPbEr\tnJ= ;P}~<<9D<l}oAqu5Q~6hiMW;/N(;fFj%:)ES#eEU]p F#y<)S6dZCU"V95BpMU5 }-3M^T eE^Ce^	?3Y"m~(	b"
j=&VEq}ixx/guS{XDP]t#tU=6l*6 (v(Wci]+B^a7DU0>W@~f!LT_ir"1(.xA6WZVr_zgB/-}y58 NOx5xiM@1Fa~6 oQ/,Ow8q@f|'FFF|tL~9s7^/j%@Q6Bs_Z]["9t+V++y1u[wR!\y=avE61,N+ZY2%Rc`Aouu2}KX2hiw!!KBF[U9vGH^9KfkVnY/{7O_",E}sY9bryZd6.+>$?r6l0<2OHmS:R>~yQa?<p}d:.u^^f9Z}N4&F@5 aCP>H)=O6XA"> A_896Aj&NEFr3qB(Z5..Iu!32gR/eZ
p;7vk19A}>MdG}Fo?O2>]J*]XNi*K[N\X#$HG
i@0lt.	0&kpz+Rl
MM\/%[K;NB-%J)J`Q+0)HE1@o>KmX+rP[`&d@4M>bZeW3DH4v~BHaS>3Cen.tM_qWJM`[{egvTS95*&1~>E Q*)Oyl$zB1[7RF	8s[eeM$%Pjf~~Hm1/]T#S-58~H+H{@3H0,n3qt5!`9lT`fm
YW,ZB:]B4Iq5\e\+YXhmQBEdsj^.^E
&MnU!\K7E?L+yrDL1	/3Tnix(3RHQ7~y%We^(lQO7^!b_M4lQ5M'LMhySE8P#^N4lHiad+Og~OV
fggIV0B)5^s	`-;.t-5@J0?R*7f3[5$*lq(`4xQ<aEkkg!G+XVKCT1*is
~0jWLq|$$lEbHd3,H@kfDnX\uS{yxcY%FJNW3>"*?UR)=:]V qW]T5Qp&@CN*HW#4llO9]?;olEcol*bHJ#xA4PVG,l@E3M"-RwY 'C2W]1v3cl&<,EzX]w#h3,Q!*Y$1od,1fGeUt=-./JYCTc~le.eY),Ps*Qfh7R~pbgVa_|i^I$ 'u&@$}9z`P^=KV6Qs0n6<e+D!IVmMbng93M4;wiBrTrI1y^Iuxw3si/\<B=YMx!bWCE?yk
-|`TV1Sf:"XfE[y/<4Q9>XW4UNC0_9?;Zq+9~){	E	RYl'Ev$K;CvNAF|$Y	>	.cL/X64dV(R>3N	IPoYoz2W\KCg#$H	Q;S~1~;a8
B;V2?8b!B\(H ~^OZ
"u!leu')b,hjSd7Mwm3]YqPO R:Vq	e$YcO};){/x.,p:5b5fv^O:RN@[P5'<Q>#.;f;C4i"'J{q)^KVEJnig~]ZuH/IQx\DSKy4:65Il8CPcdmkim.$T30FGrt$;7ZHubS+y|rDn)RP%F9-kDS>(4hJ'"jNX2q,ukjp?vD	,-M9`FIGu7a^eUPYb@8wFzDG
BU=7&|CF^
n @O>%z_%C=#4qVSP^tl!+XPDeE1S`MiL^/G-W0Y@&4Ew}Bh8t)@l.nv%&4fC}lcfzVlPj[XUaHzqA)`P7V[XOi&`#-]N7v=
lX)wRowWkDxTfTU,7ZU-xXy|aA>hpqc&K~JFas9
["8EFI1.%-l<nBm)#NE>T"=?yG}AY)	kRDREwMA}Sn.!u$<''^,YaZg\Ln|G^LFYSj'3er`%gvmdOvGr0]Hw03mf\0V~UhUv3C?rru{|iFx.~PV#'N`($B4:-54_YV|\A{9+*9^\j'Rs/Ve%G,L$d@/h~s7Ykc)G(hurupx6%Taq}>Byeh@gf=$l*HOQG;j(zp<v3!	a;c*Z68/x5^ .wr<#|(:JoU \.*8FhkN^ Ph|DCgk^Qa_TttkcK@)s	E>:ba5MWcE(lrlDF,I-u*!Haa{
JOk0$x1Z'aQxEevZU,<`2-B+_\UPLrkXdgD;3o!s3N}b*c:R fzo(
r|AC)E]N2tQ\AF](uTXprdm	h/'S=Ji%L#"ur pyt,
D~[1%#*!C{So0'fhoBaw[J#m~Qm}vM<phbkTf3[ f*=q@2w (]D1l3['	*.6!oC!=*?bb\qGOOjck6IT)RasJbLI{Y7#`[\^geYn}R~DU)T]QukS(sx\6?x%wSH/1;$"U')#wwp_;<2%E?rBTp+-DmKz5E''8U: xS]\.5^N[1'l*,`Err1.
*P!ZuX`/T"	>MzWfu|QotoMCX$PBa-	3@e|Pr==}C^xj9Qu!I5RxP2ECUF GN:7BO	ompi	_@5!%!IY*TX.=sSd7o(o(mkbS`O$nfKh6KvD2[?[!QOD~;,1dRvkVv)t:s_}(	j RW.n6E;Y;m_V<[SMY6J0{Y{C{{:Ja[}]8@,
19qUK7{FftBJE"@vH,UDq%X[w]NxZ@]^J(lT)I2A\?@Q~LEE
Jo&rnKTtZKV;&t:TU+PX;}';Q,"R~iu_}rAXkto~pK`%0ZxD_l\!>4hm3Q?D"k;~,TOM:}*v&K*4n8ooA#8.D[t`b:kNJzp@1'$&GIRkB=^G{'Vr.(ZSor"]QR_y}3/e<ouH,+Ud,}d~+njWh5$V'^8vZ2L{3]M@GgFyk<;Os~u^M!Ls+%SD-Et!@b=SVXx%7SjvKW8kVPvq>:mkrX*K@"!Wi}tLi-s7S{dy
+R
w7e4LZ+CM@RIo\9Rd1_V\)11J 2&`t'eD2,U|eUNY	l|IOuHD64-H[j/o1G^EmLB&=Ae`CH'	0vD=1`Ui)hwLWjHSg1GkD-aUbtzK9({Ut z>oQ2rI<S]O'IIG/75%mOtJ#(),NZgTdlx"w6<gvb[.T@mOi\qX%{"zCK8
xGk?{CNP-h&KV|gd!#wTZ@!svR D?49eNZpU~7<o(0A\M>jPabPuCA3\x1*#f'0mg7L`g,)H)d|E1LZ^W[|
5sB&d#wp-(eQ5"e;uFaa.Av2p(T!W>E@M@wxfOSm\s',(d0LW\%+<(wn50rr
,`XG{#6@]K%Ufn^\FySp,ew"RA"j4)iGj[O*BADO`:rg5|64V`qa$k=t\as>uLTp}<jmf7G;G<Jv*Ab]fcELvJEodU?n	CLwmpWi2*}\2(6
t&	"j"R}ocp>[rXuV>|^K"e5H7a-"?p!	uH|7L""3jF3]T>FbqsIN:[
s`;k./&(dOg]Yee9:%?pNjQsckGgZ%8h`T]pcr9I?b[Cvv	x53IO1h'snh_G2Kg^)w#5~7
h*ZyY|	9&	Kow'&9*N*UzWa	T3sd(BK7%-0})G9C>LV#9LS2<1^^LTdx;[9g9`)(bGIbwOj'Z05*LdSRoYW>q4P/+
XZpR)6$E9;]I[E/f
dP)uG=w~&	LVo~S0|.;7N?0z`ZTXSS_I$kzz>DwFEjc$&Fkva!O>=as\9T)Kd>G9J?]<{mwGGZ(aSvd"VG(	jnEFV;U4$*}kvB13#U]ibBCY/:2vy\q`u[ZWPXs]RlM:dg$,PSc$<:>huK@pwS&(K/_4!$I4;!k7(wmI6rO>^u+gVYXvEcd/-DQPv?K!{Cepd+Xr3qktJHc9?y,"[xqQ>0ZzR9eq1(/xzxb5']&sS\]_H7vh9V3!	TnROpi{-fzsJ[4K{kYFbF|8vr;1	s]$j`p!=@6h/O[KKR?wN7TlF\6K|C2k9.,+hw,28uN7`{ccxnY0HY6QRS|6[F/uJ!Pq[nFGNzh!(<I:r;e?m5V7,<e"de7jBR1i'XVY?SPeIJr8!0z%\RmgB]	6SK1\NC_Ke*qy^1-?@dT"pIH!+kp'3%N!)FHUV q;ox)XO?;rpi0-F!dFk7AsD"a*(cRgYYP4_>=/N{%$VYL)q$tK4RQ_*YJ<_ql9Cq&dCUR.QYIk5Vn;*NAs's}xw(K}(QNbV$+e<VrPUp4}p\t!"G+LOT2fQ=]X %)J3(	)9,^
/sU4#7~RQQ| f%RS'U.icYge3aII(qRjQ~:R#Wf,_>]Ri*Q	WEXzST-YR$'en7_L(7y2d.:0nA'D\IlSGfMe;q*0==vr#-ss!B/>
Qj@6>'G5s`9`\8H_R&f;DbGQw}UI\kBH>w(He]h|
.R0FSR\8q??)*HTbz;p>JYJr,au;NX"&ebLl}b4q^eb}AZVjVX#A#IzpROHpO6D|ZJ'D?8dbwOS3y*Q.;3%w3X#}N6eZ]o46J$q
[^3GMO^i!opRGs_WE@wwm6{pb>pz@{p2l?:TZi	)L? _P92H@6\PHs'{'2g1%63.(4oi)'~b:Q+\UnRz}x~:i0WV+"_0`~CROH/g~CNz^}I
|sy1VSF0Z~|&x%	e~nC2AsH)_7?@`20@01$7A#NJf-&?=zZf|lNq @|Wh91cS[t=#4l)*VZhk\wV,Hqm
?s$-{m7~YSf+g$Wg\xk='WW5/26]K|t=0+X/x}+0DP7P**|D%g	%qVjZhP'uytF1^hzd^@q)A?N[\_!mNKfNz6^O#_.-On+pg@7C6jVj-WZ=^Gp#xp5eWR/<
Trm+'%^|k%fzi*_z6L-qMLb=.1|O)RswO#LPy47 @)hj>UVIQoSOT+GD0e^K8Ps.'[a**$p3
YBK$b2t|mJXNP1=U0*DYz,Q	z`;fd*#q'F<qfg7r&s\O
z/prhwI\"hZ;D~396I"GA8'!y+Lh"X]+H.g6{bp9C{O8Qzc0g1!M'-Z:x0d7b{!ycQ\;!R+]jB2Jb.+U^r#*J)?@3l@$Li<B6}av}07hi:=L"jGAo	H/hq]y*(0d5fd	UW:!SIFI|?)/4RKeXa&:<y(QD.VGkxc	UKf7)|%f23}okmdWm(_4"X;zs4*c"VLcd& %oTz",7xm'Aq.6UKz^i\'*DfWF6I$!!\f,_'r~OF{.F&Rc-
zcOBiW?`hb _%YvC9jAol;M6-oCrto{RSlTS!SJW~fwDcN(g|90Iw9n;1-5AcTLQ7dPFB|/Gl`Ny;q%A`}@,lz!8su>Eg1M+|>@I|^D{>G+ ]#x=#	v6E> /LvxRE~z;t+
z1'cWGy+3M4CMhJ2A&M`A%#&5r<3hs$yJ%zjo6hNpR1}n5sJm+_=2cI,NX2R+M703C!qXi*TKElb<WX|L?U:onE_BrT}^d
IR<fI,q9\A\>;-?Uo,#y-PA'_C{o?BKTx2i
e|=R'omC9Tp^ztB5A~h'[kQn6&rw=cSOGab@0}\x6gEOQqjyo#z%ISs-Ght`P\]yI<uPU	mB>WP<re1O\hu5]6Q}[c{8&`3/\|pV]D.10XP8n
wQ5E
W|/}+^}]2  hG2Ing*QycYXTuT\	h!7x
Y]kCx3&8knQIcZ~cD}F`Oa@D](O3jeax?M_3Eg%AFIsm?*\Bge^DO=<U@b5P<;s2}$[WSJ*)!3RQ*D:	N4&>s%l*S^%$b}2
fo?}PZ6n)=;tSS+cnT{zW%=t>O|66:B4)S[[y}:1DX9$``Vn)d6}]Sz#wcm\3jp	4Pa^V8~DmR:a(p	iZKR7;oSvNwpzzLM?*n?|?{2DAaVy188f`Jp>&Y*8JK?u%E%(2LtE-4Ls}2V8Qdkg^\
FEBaNl!(ZD(-#{zoe2Jk\lCop"~\jZ?5sekZ=vZUr'ys[i<db_lXiQ0h5^z]Gz$2?]`qp>lkchg*m3}/;*Z-wvoA1O;'fR2{eu'VtIerSQ!{IcS/=3X!dRG3d~Z]]h=m1w`c57+;HcfbbFBd=mn,I_i
Yhw	"JAhs*__LY+11\
/=PZz8$l&<al^^8
N{VT
EuBrh[ay@ojjEOb?h$k0g_k050sZd
!#H;:SuR2;<@IAT*t #vp:} VpBg:C`|ROJy<VX"lhq7H5/v$NS32wQy8W;z.tE[ke>X]=Hvvu^JRLF%eW7beA7S@O\RlT	LQ.C>'5`loDEJ@>`~jbKZ@Yn(JX*6;Mr?!gb ?KMUI_Vmb^Bk^%VjDC_0DR2IBCRt;vmT-l5,X5[1xU\
 HC.?"K]H@_o^{Nb=:o"h7uL.F8v%q|,}$p#tnDwN#
yC`^[MMWC/NEkU008b vuFX.&h77j@Ol	piVH7qc7;*Mj
Q0!Qdu}uJ%V\XY>{(^!IZwQZ<~!HN5fSEy_Nzd0@}j5h8V\|(ddV2z1HnJ6D5c;|c/n6),|b|ygE+}d3W\nMo|,FQ~+Jc`)4F2EEu(i|+Okd_1nvk	p3wYWl%G=#qpkq@eCKenO	!WhLdxd)Q:}h]=vguYh}yw/yy\-'g\ya4M|b.}=l$%$c._!S_-M' 9/vNaj;C:VaQv_JX4kLaL(< iq%["a+2KpXrLs1x:tM`rd/xW'&i"Wy,5=gx*$nsZR\KAJ=wgWcy+	4ku^16(|/|g=RK&W$Wthq'1"[K.`Re(J3=}@7Z;:Y&JL"FLUPSaSVus(+j]N-b0Q&tFk-l}K%C@MKqbeJCRwtE95EHnD*?}7l4\G<"&T(AupWV>Y5hoigQ=`Q_~wy^`SUBn~xbl)rMoRrhDu@{D91z>x~*MHwV'7=n5qcR3b-J|w/Wp9N,$
)^h,4sPQtc>?0JAuby@5U91\"DzLv'e\@ht&mGt*2>EVkf[Gm.M)qr8-Nl0>8~z5X BMnS<<3<8y0n=F0 J{7>0R5	.YlH$DP$"bGW;"AZe.lq0R?Kv8Mw*X#5c?NvMT'XHfJ,?dq]Pt";SL3~wkUN>kGGLn$c1RH_xZ|P XReO3JipsBP_yW7`8|r_bd=BdLO~fG)ha0vEpWjlBl<mUEMS\3LeumRb'x1!&_?.f+@w^B!%mt]dP/{iVw &:*GAX10\l]Ne(!7vE/{E``KHW"/Un/[LgDX)xc}Oa^q+jMv_#;zT5x6F@eW2B'9Glx"w=:+]"yLcVM2Ce/="GQF7bCDEH9}V!CTjbhm1{O^EG8SgTHg^_0D(meMY&"Y"usMj4?vv|=aQiP	LemR\z/5\!*ip$\/mfnr#-MY6*tGr`HdcHBC8Geikw}uCz}im*{s#u;Ay(NGOoc&x/}yNkF&[v|/kUBm=0R<!l+}	
xzc0Ul{-j)w?$]Ao+&T7Sj&1L\m_ClFG5;t$
xN9F,GlJ{+@vQy1u$y6RU]8_{[M[,8]ihi(lP}wrH4 S'#Ed
O'qs,C?!V[j<wL&EV_gqO5=yQT>ITe%imMQ^:lKAMPnrm?Y4N)oizmHVT}:AB#1Ay:#H,	Wje3c}g@cOz3k;+zer4I^\:NnOo'`Db*@w5J?qPTN3J-+rVmu/B.TrxS8rqDQHXm=|b2fE=\jd?]ez*3>P#)Kfe=VF'6A P@qs $p]#?CA}\PTDt7Kg{*!,CL8i
S=];\_MSw[V37Hu7q*w7rOl]72]Yg1VUX0]])Mud/U_	?a><A4ir-"i-['GtSgmK'Ub8Z>}9OyGnAL}Nf3-rn~)MYRYHb%Rz)q|04Q|U(^_	_[xYO7,K /_j-/+K?@r("m/_!J"z?yxZ2N@8{GOf[F$p|D[)=K]mTTpVz\lx][<p5tY`>Os3$f+n{_D	)j>\WM;V-_Y!X\HBXL2z{jb}}YvN66$r<B!(ZS-G\SBI`8	-mE*!&A%(OzZ;gu>!Z\\P\G3DVX1HT{22; SXc?3T$'}MKy)z#B:uWrb#t@pnlG^<^0>T1^CB9	pgC[MS3\WXOifc}cetZ@@E7x2dC4D3*Uge_2'8&08},93{q B'}rh.
>/nlY'AtGZ
b=X7"PD*v@m'=$7xJ	RU+\Ltgv<{Xc*!iNh"%$Tp@KCkEa*v#N35!F>#(]H1DPiT"'1$QAnq! =ZI|L)QUe9AHX=uPdeX*2d*w'8"-t0]]3|(S/4;^,c}&o&Y/PeGXgbMz$[reT<Xp!`}+DKx>:va9\%i`le1,c|Z:O}#z8<X<'RDD,.*Vle8s:B>|'
s4r)egdJn$L=J$rx*crG"FW/\LI(c"q|<;h8r?<
LhC6r`:UHzW%*ZRVVf!~t.09vQ!*Ylbs[G2\(/?2QCor;v*Wl8kgYvo),Re&(Ly{Rw(NAVChKIIS*1pD;8P,f%fMxLpUfj ym4bRfd/#ISaCH-lt{}K]ChKokfkJH2FO8xv
|x2RW]-N([Bd	X6XE	xA\E0eOX`,!^LOU)TE f22gC*!s_^"zn
f;[:*<`ZND@>HX;COWMj`|v	nK0Xwl9b}^QMCQ.@&E,+a+hBY_cs>!3*{*SsJ,h6Y(%`Mqf5tr56sL3H":!,Cz,%I{,CRT3=E\\p<y,wlOK\6{(Q< \Fz)+%\M[Fu*\`'6N:Qn_a8IzOb>@!otXeFkshCz%*\6@V\/AY2c3bnfZ|<5^)YJ(SkeO	D5FWB%$9e%vI!`B.xiElxKX@%QOOj,[v;9>nR:JWCoN!rS<Uv}EaX_i<)-LUV0igQD1t1$!X4[-@t(Y6GK_LFD<c/c2'Q_'JW	1HL!!ni%,*n]%.e)Y "(z;!3IaF^A@%m~W;Vtam-=A4K}=$HhX<5Aq(anV*/Ke,>0??
23O7a#)m)"zr"<q{^
O,v$>@G0>P&A8$1i4$U_^R?!`|=C6TWb"	?7i<4KC0xV{k(_vaE{	$//5MO58uI.Fwxrd1{LZZ@+jIKVHiY[whnC<nL"l>mb@=wMiP!j]40..%vqZZaQ;Hg}ReP
`-dTA0zRz%m-Wb}M=i84+Z'BC"qc,
k }^2pa5W2xc}n^4T+ue$	a+?DQD]'/NJYV3,dTi?X%"XKJ9{@AGNLr2tWI-dFu1KwH&D'"I=7|=-$!@?xb:Btp"V7cu	&\%.2,UP7uilIE+KaJ}2Pvr kyTs
2.b[\Y!^J7qKY}^nbn.D(8-#,U8\ornc@Gnev.]w1(@Fu!wl*^4(^g/an\|}STG3W\):!mM9}9@SKj^#
/1-GrT|{	Y RS%=*5Y|s#'57%CNO!w|sv+G1h>!7&PpiK.I|>kB={3K-p$Mw/di1}|h,3J^^E_ey<tXW[xVr'VyHj2Q+V:\-4l$,(/=Z%Kx<X5e+43,k$hU;^lif4_s^t~^DwbBP!Pl==$#upUIdU>,_zC;w}T[$b_1l?#sEel9y}5q1$.d,XEA,slcNA!2se$CB2Y5)D]xi<d5\u*`;y"Ve<ud{<~k3zLU;EA:S\z>_r>MCL3CLC5e!.`Iy*"VPc -Lxn\BP)z$xqw:c	R1Bcj9!3?IDVxkSv$`(3.C]6#0s8c,@CNy^&7QM4M'=1t"F@{GgtJ@~}JY3a-So
!5{t>Dekt$)88*K:}#o6l**#F|=m+4HdkP%2Mk;
@8$(k`#;-p+maKOVUKVVZ*3y\3eTWDABxi'\1QDj&/4l),_0	<1@P2lnm^nrP0/<j>,)ncovz/NlEgj9p<dKRlsZ#`vB}kx6|=8we^>&P&nL:t[5VnCM~?x<(`ybW$d1QC{9s9~hl}&nZ$'msV&&WZ1[?v(GwP.lfaA^W%(QfJaDxI=GA _up!CNOW\-6_h,ON/ Xq[6}"w@16TLWs<EZ7vTKKG>-Pppw(@o*zmOhny]8TfFDKavqToXw-)/9v]UbWJyy8e:r
enBHS(_w0~wzJdfK|C/9/wzS
J+	Q2sSN!
a9Iey5N4=uX~oD@VOn)#	q?q`8G[-EFz:&q*?&93(.<BR3x"N=,k:@,Afc#4^_IFX0A|(|9H%6ee[>#XXyD}~C>TSl'PB8HZrz|v.[m[H;!="@;@4uoH\x8SpNL	,,el1wkxGh'B'i1UyMFan8P-ZkS~3xj_%5a&[{v:JZlJ|ndRV?^gIz.1_\;
6#eO]!){|JQ#jF%O{w?F[?^5)!e<l4/L84ufk)?FB2n:5Ra'09xhqX`cwh*oVj5B2d>.iPG;]chxKb=0rak9X5[ gEv_0")GV*/d[}\M\|t& 
i
{NNP2Q6;^Kt\p[0gp ^%<9mpjEYj"5
3P/p*!9xOj:T4bI`EP&fhfZ7,'RkjWPK.{p5g\wF%BOZyb|=c4eH>SeL`Q.	9m2VW?]M[L'1HLY>@HO0%1O6PL9`W@SeW/i01`B~=4'tTp=-*.rpoS2,,QR;}DV9Zc>v -S+>f	W*!nhcg|0{wIS*[D.r*aliz*_E=3-U3W B\Kf	kqzzo81*4%#!E`jH@g,k/l7ad1r:3FI}JO]JxdX^stGpCZC9ND'[(?	lo<])i*T~k@.)Dq2/a`\uMwR%{w;Ys>xwzb<Q_5Dv'!mwHA$RIk,gk4t<g^m-[-w>"epqD ]]%+|43?h="\/g#XQ} Xi^&R\Hyi"mr/CLl:m|"p=%X;0DscDVIMN?i_+]}EWr		Fd#amqSN?/sDi57RDxhCYV`MWyi[uVi+"rYG\CklL|-wl_;@Y0.u-tboe9Ucj2i-uR?CwR%)XR'{x;L4zPNQ{R(:7b5`oU -3sJ(VcS!gU1x@UlW:T;L:S^aDxvYlpk
J8{fAlg.Mj{)U#QK1]Vi+~nYgbr}7o=	%/6vX2c|kgCH	P5Oj4pG|AJ6HvKl,QTV'G!eH5zY8Pv	 -W~dI1"V\@A^umf._A_G[fq`bGonUL-fGA)TgP_t7{Y+@Dr6|kD{9ix[[KTr0x'Bw>d_^H9_;>0Ix\Md,>FV^.>"!p2TPXbB{3<2=reX*Ds"x(c(,r7ufSgEfcCS,L|OGE^jVHB5RrF<o?#:T|!\
'":(CbTT6vR/lG	h/=U^pxZ|KYlX~wXkCrtg{eZx 79\#kj|<t<D;zZ#%G\=.pPG &"O&;!zU\OeWDS0>1|*xDwBW\3xw2NCe4Ec^CYJt#Y:Z7u7hp*A7t`]xN!9|0d+2*58?'!W_M?ysI{' yU30\#jLU*r7:*18GmqB<bDH	b0%V=W~&A~p=)JxnMZGE/CYG[9!K.823oup#U-EiM=G&nE=6E!Grdv_}vZ=H& W\W!ue6#K984-i,	D\t%P[)5	rKef*VwQy`wC{78eUW4}J{HvZ	rp`Z:o#?8V2Bs2jsz~m JcG5Uk4-tXD-H|de%lNYg9NjGF@Y=U$|&FHq0s+{fQ:Y{A"[u]?2[hP?v.gYCqW1gJL_RaJ6b,@TvBq4v/iyt%8#f.49j|%[[ey0dnqfV&D,:grETqKt;lDWC5NdhTUsnY	{|G<m9$Sh7vRT&)+56(Z;Bw8WQ0)Y'^)*!Uvc1\89mP_h~cU`J&]0E9?L8OWrR23BjL'1EAxynJN=[LBg@H[{@SBI;OR47f
,GOegN(v)}Sa]HDB>Nuk['2Yt=3qm%a_{/(F
"PX-i]Fe.@nMT<GW)iu=i	ZNI1sh	&SVjU`+8,{vO9c{+ADq9zW?5V+lrwNe;-mbbh(T}w,6)*.b#|=e3
Q/l@d#HdciZG"QU7'#v<^/ufT|\.sg\pnn< gUu{TwAlUT1n5i.~,weo4hEKL!MrdVA5MRM-QuLr7b1>P&y;|HHJ3%j.t8Lt_D${9uv3vV;aIb*`&]$IK96B{f$L8JL/H5my6e)#fa'A$T'a79bIBe qp<c{?"59jHiVwo!~A[v;r0RunJySgVnF;W\
l\zIw[b8C_b)yU56S5eyteT(2/h|CjT j&3]j0O?7x~#3k?<bz'6K`Fa%k?mz>hpOLE:l*o*q$mYQhdvB~tP3LQ3%;uw{9EWe<c@FKjgb3z^vKTo'r;d)uJCH;ayNt7unSI#$QN&COvZRt)yUiU(d]$;|r?lx7;{'F5apY!/|O"I5T<#$!ZgZdVZel(J>LqO~?FRH!5NGDD5^;LZd-(	FZzU
C>Z`:m#tE./IN1.T,T|@\HCra/\E?jl@,C01q }[f'
d<lR2\"\>t=m?M$_#;zqiz"n?	B^wp\eRX!-3whdA8JVS\KylQFxhDMfS'0H~=gHKxj]ZJl~qGB`nU7{)nK'Q/z):$CPv}z"SI7+!a|&=:6.'Fk0#4T
Wl:HJd+f~"IlW+i`*Nra./M?/NK4E$+/Yby@87Fkdk#Ls)1GwxU<yfjv5%SS&',XAAV{&}`CCBrLH5s6<rGHiPo#` g\o|8'|onPx?Q'Fn~([Za9BBgU01XO{9Jf61Vi4TwZg!;Hvi9X"!4T(_4AFO!IXYI.%+A_'hxIJ5FP~e>3-yx6KdEdwi$(i$u_g6Sg|dD.m3cfSf[xUSqp\}gY#|r<x`dJ= NI=lL,yTp2YKUg>}l$>_H	@!<1ctcmQJi=1Is@z'Ay2r%	wdo/u>H6ty=*WF!N@O5YJu=3,m_`UuDyK_E%ux>nH6_Hns	0S83s50087PzR".LJ.>+Vv|O]7~X,P|#rAKZ<P1p$uSUULm_}s yaVoW2)y(e|q7IJ\w(Vq7sKh`91+a'_Af.+lhC3E98ix<291D!S:D\q!G+G.N'!?jxh(u0$r]	Z^szM)p$\j\e8260i;2X:SYC#oW!TuYn;Oy3sl/(3Cp{zO6X8;wAx|G
QNgv ,ie"F4;BacJCm&A5keHPNOhX9bXCwtE.>sD('+#R9IAn-.a0OP*B5:D:yIq/#u
m ae7('.FE'}erQ
d[T	vULDp?A,ClS\PQRiY%Ag	sGOJ UMc,zlP6=-/TW8l!+]sru{6Ymi }PZ@Rm|dlkb$"(Uv:2Jo?LoGhPw'cN}udJ7-ZZa@gfyvlht:g=\V#'5 binls4A)ZPZ7Mr6z_b=!x\4ya@9iXIQf9u QWRokgDyv'N*:h821&NqD"a0z0jVa.Rom"m`Lf.WwAldr/xrh/P&[muD|vbbnXG)O%4`jZrZ:g-jzY!3;WAR\k<eT`|_?@11G&n/5wW'CdFu=!c?xzJh/{wlR~p^gj(<Y//,Q@[Y-zAq<fSQm;8U+quzRWE1#\AD5]g.8kM)Zu-hRlJEDqeDrhG{9*ZhMSc[JO.$S[.Uusdo*H?^5
'E]>	pwpk%W[}*-cp|m9%I*Vxn*vkmL$8'LJ$1UZd 8k:i\'|B@OIMiY&[YL("lbtLd/S|n$b|`b -0)z_|B	?<"s
.p86!R9/U"XddMalN/lD6Wv9WpZC.6cOHt:2<8_yq..`'DFbd{G=m?'R<#!Q;C*AhKi[x<	|xuTnT9GVQcQ=.[1ynM:BGnF6"`S&KS.72JgIU"Sx?T	y,PT8.e)@m{gjpIP+M`F4YwI;N0>
USQJCK4PQx9]y$"x<Is%@$,0:\:;=YaNU=was:R-tt:%50/	;ca=i<_rS)Rt2u
_-@uOa8LNMM{Ak3*cJoFt'6C\0y"rgE|Q@F5chYR&.7,>,#mY#zZa:Z\RP.aNIqWeNP~]-Q*Qz'`-Jww{67s5(h5gL*{n1r?)'jhZq.=>bm|!Q,`?qL-CJw M%]+)jl!wQMuyYwjP9#,NIMSaeEraz%<g `MtUZro)p3n)Hp[fhZU&#!dgtE$]$b~rP|YW&x=9	V,,oqRtQ8DHgH["nT!7Ap'cyS#2D0
jIFDOHVyF\:*6kjXTo[m4{Q*.+{a<0pqG<)YWQ=]nU3t\Wi>F1NoN)(N9T<t&wDR*k93`x+-E!8;LE%f]%'yTKQi:jEPJh"n*Qj36v89o2;7JB)1.&^H$L!(XWT##6N}p^&M
B'H5gu#Km^E pyW{@>b+jcogP%zrRI5@s%UX$E=BbQ[T6gA35[GG/$3MT{SQ)*UFw 7V:*L~x>o^xWHm(Xn*?pknQh>$6x-!jYjMV{X/l*RuT!-K!d~nc3M8$Bj+5$)HL^<%jcYYd#ip6[ Uq/3BJo;a3e~5=E'y0NqulWo/[e^O?G{l)-#z8=Iaks7R4B&c%Y?]4XzWN8TF7V22>}&*)*G28z_x[_%M&0ej9iu7VR~"U}7m'm2w@>Ta"z\p&F\
NV"BV0WEP`Iq;Li`>a^-(sr<p=dMfiiA:W{)g2~:mDZ<M}q1ee&DqxClt}iC;:2zbf>T >4,XGt-	/;,E~[?0LPRbik)l%}i\ET+NE)c0ZigjwNA1ntj~>J?IX/	>A[.R!=@@iFL4{"Fj?>MYZKH$B=seuP'D0)0ntTB0	N$|3(]-aR8Uv5KQS\=&@sR\--Tfm29oj9lt7`Od@g8-X7Z)B3dE0vvu<\[#n!iY>U>Iq*2@$54<7M*:4vwJ
iJR@5Q.j/+d%?zI<-@9i..,erbO	u4j7a,!9cdf}9gtW-k9O`X	y:G~7.D(DVty%D>:KkRIuO6RJ]jkB{mo$i238R;eCovSl(SgT_9/PGWlN.x	|fF4GE<POlh,v2b')6+v8&Bufw zl" o;t^;^eP"g[mw-,7aij=SSPFIf}|HbXW2/^Y';V?D}C{0OzY&S!gQG2V*5:BQXK;&vTFIu/}ce;^+G_1V[ZtOfbI4*'vUwHN_VXazKM1FrTQNumg0]l%l>bCJE)h1
xJH.a5TJW~i`~)hBo]'l&C#Gdc9{Jy1<6Y0)#bQO)gV{("Zb(Y9<=5v>.p(Uoj#ZCD(gTc@l|7DI.\"j)R0sF%V4_tf`Y:r}l186o#JCndo!EH0=@Wy4cKIrP ^b)]2X{qq,|Wkz6#5_^X(hFf6Y`Avue=D)-=9	7oXu}@$3X/[3pu]x`,|Dfwu-,v};mc]4NU	1GEPZxrEG"emP49F3kuMpt0.<uNRJF@[?Bu89qZr6fuQ<8Sm9>O5
Vitp|l;Z3N`\B1a^TerVBu#KhqsBcrXc2rx?jdd/L!?v{>F3PHjQ;@qP{uf\Epm!\xW>DQG.D)$M,}@ziRtICPJrK/+-l02pke:wf=$*35:mf4ebp}@L^L;hw-xd;l?LF&"I"&3Tq/ed^\n6gbL.[&.YT_b<?.;)o_clV_cJl+[$Uo!!dXqO 9'ePv|::_GN@hg0wG`,Q)sns"r@p_#:p @8v)YX>unNxPIPkxlrqEr8iwq$>qZZ=xcFO>;Lk\ZR/3I?F'0#Lw"lV`R(lW'D98ugc.Rdvk>zzBhI![S/\jG*r3u)V/+S2T\_vLA58P)g<HDBO2G5fro[*(k.sCJ+]p(kW roft8`#='%mgv|hdxB.V^RM! ?.eC:kZ@J5A}3k0/\vKg@{My!S96J$y:amSk6xY}oS$5Pp{)-#-^S5u0-;4S1r[u"kjT~bMS_o
3j6_D0[h2(+.0
L,X,qD0)!W`X|()Mk"#!,8^`;E-u9 -7GRKO0.>Zn*'\ID;m8Y6L_7q$b>$tC2CZ%;Yz[P%-p[>ft{
Mhh3lj-if|)ON;i>D6*/BLOpS%i`nB2W+5NAt<?Iw:RWZGs5C"leh$$30DH|5dJ.\|9Og d&*0[Yn_@@.tTo>fCWWt+WHM^4~myp@_0Jm208I)UM~=dD{!9tZwd33[tK;l%k saj!$c4_b>
>38oQK|Ekh5F_<^}@;4#lt\b;fk%
Z
M8X*&(MjA>*qI5JRakQaEm:f_;O.!xL#r)?(Jxs#feD*k}\a][?RZ9\enjc'V|$w*W{p}^Ins-03wdhE-:zmNr6f._"LP=F8Bwb{_|1~AjHZg"F/ qF"xD	i{va"s`;$	nfMrk",P]@7[3'diCxA(j,{fUBU!}FqR8GPK^2dX.(H]es{L@`.f	 >k#R	$8'6i <G6mS/neumWp0`t4q	rzg	/JS\:VCh\";$[2V2eBs"BZ$745z.5Sb'55Y+^K1,ap&/@pl4x$d,{o@;#\$klnV]] rY9b0:@5%uFNF)@PYb,AN23J5#+:&C0dKLASEBYm	t^zWYj&dCBv*0^Qix!V

2[MM9><s&)C/t>tRk|"##\#5rzS5'K<RYV&O)aclTRJi4:;cWhA($Js8M	KB.aEBCOc[^3<Msl&XW^	PO<7@y&0{~-@p.(L `Kt?\*Vao':Z#8V	@zhIQlqb9F@sM|p<H70T>5P\F3.F0[-EX-szCcm)Z^89)R	B4R_8ZJd@_X,1i,'kE^}(:|bZTLG5yI:d{8F	S^iM,$<A1;vz4iU0Kpr1zOhkTl>-Ux
)@`Ns\MFm+,>5nUbwUM|uz!|5^;,{XDIvw~L@03iTz6gJVxdXS8f)J+M6'c.A<g=%Yq@z '`e>q0Rs?{LV#(bg}V|U(WI-1_'%X7h1z#ul07U;*~\3;*xP
aOVRC@-=abo?;5ly! 0r,~
mT.=Rz<	nTjg[Ar`?pDkDC>FW"G@*64pG9pad#n0A4!BE46}h-nu$gro/BwxB.BN8{vrXV#y:G;!(]om3Wnd,Z3T|A%$gv}'hlM$B3K'4UnjONN8aGZahM1u]}kLOl}R\HZHYR'e>w{4
}TufTD)0 1v&[Jcq@<>yx;[I-:"*FgMIp3L=n,:/0Q31J>\HbK32M`uqRYe2taAyFJgY>=&'~!ewi\Xa-#&}8v"XGi%qJbTN#p7/:|Pt{E$$~.3'IYkbTB"95<]g)fZt ||PKOqGPE(J[1_WgEH{6g:cg'|4GH2mcG*[N9l!pX-WXKz(X(aBs[+d/O#{y-TNsOXeC{ykWv5;|'w)Jk1q155'f.JW:L5RpqD{+i^/2GPh2/Y),f*$ZS#j(R{ -~*winQ^Rw"}gb2R~su5	l&ZNR};0{L}-oIj.}Wvltf6\3qLTI~)C~mK,	O462n 8'{`"m>at)g`&7l`)p	uejprhuMq|P*;.gR_X{K9,)1*}Kw$dCg
2&cmGlss4Nq&m7>j wI(1	&`CuOML}!tHQMY"A-N4GIfJ(\161G;gnQ8V9\ 2/E9PHb(3~VM.
'yVVd-F$.M wjWhC%mbZN6083;ep37+8@\cuU1^@QP1<iz&{$"G"9&k%VAhHxZY479U6e_PB04PEIpWg2Y}J3(chG:4{e&B8*71@u*m EHw2en> L~K.`9S^%	0ZZ'??,)_N@,E$`ZxVM}\B/m?!:/6pBfDl=*_w$|=&CP)Zfa]nFs'n5^i9teit_7s.`N{pPQFD/vLF1mhg[^#m";A\MW"O_kHyO$y5S~l!)
N=0)!p/Q-!>"h[BI;y4x*DZH8/o[;%whPWNNd
O=_w[
Zyg/=i9[\B</4vxFL&W^9Sb3LcQI	7sIrA;kw(]YNMAwOS4g
/%2$^&A.KoOga)sivGP=z`[fjEm}-ZUht!@o[$XtJ[x3a:U2uR"yb<i
CWY+NT/XP%o,iODSBwO?Uqm*&L?W70sZlwWZ2q#\><1gneFDK,uvdmla@7+b+SGX:0"$OvKufH11mCpwl?B++Bz{HiLB;x`1NoUaN]J}KG^_75\DiXMh'VA'%#kBp>2c@p(r,5KRghM-"?)%VE~D<oMuS{]$8v9_x)2KhL@O	VvN<6tHq:$hPMZ0?X0Fs6t[_tL
9$BT=jpLB|%GWV9B#$Fevl4GAx7'NdSZ!H"8JGq\`P,^{/F~-iStIu6j>5[-2E:(+Q5gw<6FJnm}aq}Al	16kLQ>9HKe6+/*`RhW4$T<S]E7.|uGL/r^he [L 1*P	M|\cT(l[q)r^,-	I,2|D`ogPZ?)@bZZ+lYZL)
SRaW}A%oU '#bp6L".-R|(&m;`.Lr(pMCO1(w^l?VdGeSh?7C&e0d$9uv%'z#jYRg_0="l)1bYm}/[(1Jb-<Ukq=%lrf]3@]b'1//-L*1=6{(<q4U[aR%CNR]~W`-cE? .EGe1%TtFzb^9C%KG)4kr$	b"?KWyE+aj> b}gX\8<Y" Dy#%y(Vs=n,?le 8D4r)	g<+N'F~rs}le$M,O!/9>/B;\v6u"7teu}#4]mJufnQS
pGF
#b*X_/'0EmH~>	ii]w1kkRsW9Q;25(\o<#~i
-Np7	.xs}gJdxCQ!$FZJo7`#]![42&mPuFl1mE4.8Tx3'A<2L"Tk#i7Bc>]h!+q1:6Df	5XSe@6x7,D%reXIIva
AQSK`$$	9*6<4_fru*3@oX#o)]kQ
(mkLPAY6vx] O>w\
A(McL01!`
x8DCYS$p8^Gk<{Dlo<3Kl^T/^`,Y1)<8Fz<{3a*gaXZ()GBgEQftqrb<<%yj("G'e}/BZja(I_n5	U)%8j#+[dT|>`pgh_LgW9*2w\:Ut#12%j]2=f6C(XqCf%;iR,T:McE7E.XrF!-cqX=R5)Od&THag	b]k].yADR\l9'N_rla	MiVxq_)a&-+<%[MRd/+Pn7C[A/kufa$B|"r='t?Lt?!}pN!zJF&NP@Ed0{	 bhsQ]"AumX@[xq22^v//=%F&0tUgwg8y-#MC6;(n	B_UqS7]lX(h2rFAVXnab4JPFz=`Vf80H?Fp,y6D[[A	sS|2sbj 1p2:)J%J+%0!,&D3|R0TtxZ0eL=v"SFy!hWF+m*]6.u{K?#'h|_V#rtpjn!.][^E.*E%EPgTYgX>; 4	Xs
8SDPi0;+#pS> i=+W7Z#}HndD"MhmNCKlMzs2XBR~j9 Ym_CHjB%fbW-iN:W.CCSI6kF$'g	G)xTL9#:lU^n'.SokWb gg)Ox2hdeJ@Hwo&<IHa7.?U/c*`]"7M<[vg"8lm0+Lln<LfL3l	('T76Dp2(k;_)H?V7w]^.
.$b]&xz>2X*VOg
K'GE<#aPWNWeIemle^r{#W{n@o?JZ:87Ov5P1J`NaqT9Y"UNM0:9<i?X:BF2:I]x123;*]P+;@Xn*1.*v17L;H5q|-~0/<2J_h%+.[cV9SDyyuQ#l;"zwJnBPB\';`#@X4qO"Wm)F_dDo$yUng1[KZt:!zkv?w_030P!<[St&C	5P9h]jK9>iMO(+,d?j[sAulJSnq^u&;wEt'.%34aTg1w0!@gUb>qnuq-DV#$Y5gH#g-B\t
]J'%>d'-_/>?V'|&O&y:=2)EH2^A`AlaY1MYpd0\	+TG{KIAwE|i+B 8,cc%uDt3":F)4#y'/e~'GxO^UR	_^xdr7|[lo@6O^y`|1+IM6u67./=gc^g[ pnWGYH\N:M1VGKPvsesP,/8JY 5I[mt`&Jw0q{bqIE-kX_ah_8~?ZQrLYqtnRWGTWxb4Um<NhM7&1tI|2>72E12Che.ZYQGOgJ]hd^.tzQR@@@4ZFJ9w]jb{?,k~:0w4nH%6=Lh'qs~\U:_)lA:$6ArKsPT'2b i+B@\C9O(Q#b PcFNV[Bf{B\mx29YEvSCDK1r@xk^$"EURcQQqJP{W@>2(O1Kp$Wtq?v	ESO@zG>K~q:Nk(v?wFa?5M}NqL-YZ)tJrq)?(P~[+5xFb"w[c3Jn3$Tk7=NM$k7r-w&s9nGH-B6d<|v$#'6?2_E(7fsnmyZ]>i'4X	l7lIEUy$iH127:c|-JolFue;>`ZMj<w2 z/LDvp-GO! Rys(s}H^wVw5{I	0&&Gzm26h@58$E`Ml$4PLc`<;8ou} <;$thcbVU.zD=Wp!\Y#y}HvM*PE@Set/_=B1n
\vexN<Bh3^Kz"D6lb3\\\RFJ~_!Cb	sb8-Xheb|.tO,$y^aj66"P=dm_~}WAu<fhm,}:a!rg(CAhb4!I#=u0C*4i+>o/7]Bq
e.29L3|~vv>VA-w5P{]nHr`Wi{BqO-Qm>SZQ2\[@cr9%pyMrhKd$`u%j09l$[R/i)cC]G>'|_t;]X0z@j?G=Q.hnMF(W#Te]eWBZVt:!r=g(Uz\wil:[+njO8z-L8Ocs.u-u ndwi[~''?`1b`4CJ_.Q%j8+T}
c)8~C$DE+a~Ht,	^
G,#N^LHqmBu6>)X#qMTbsx:Ggw##=}*O.%v59s@njZj!rjqd#'cn6Hl=muWU[iu#vVxr^Ir*4}2$%,}wn nPwRzj!-H]`ni:bDW"nPs@%4Xx#K:q(]Paejo @X{MvqSmAK<?%`c.&eK|n5#z1"y=JjT'qk<*V{YTl]B9eas!@-g$+!ln2~W)w|1$8T/q	)_m5.+swAbg0]&EYmBm3d=[2{ju9v#w&Atl<;430cH61HHusV(=54K::\6	
-^	d9	Qs].GCHxcO,XB3MI?ahp:@v-/w%_oXn(<-w9v2}9o@j\8dPgY=I^0c0aRDQKlJKJP{Laj)_`z(w-])h8GA)Cp^B(Jis\m^Hb5WIy5
9<U_iy<[z$T.x|Djj^(2A#\?3#`w8GJ2},p4rJr.kI+4IwVYevb`Bsx2`hv59&q@PG1o0}Uyd0{}k#+SKM\pCfAjAc:hGiKxg{sU#R{=h7lLN7WgLkb!`*z'2mn6%X^Xsmt>[~:;*?#KNH Rh>"k`I(["VYyo:(`8R2ko:;jV*Cn\I]'7.
D+DgxByDF3=fnn/PO|a%ta4n6{f:!b{}bzUNa6)4s(r6S=mBvy;*c'RpDTAT&{9YvXwi}recz|@<zL
)p,b,m/mOc%Bl,ZFf,B2fMbdGBMgg=V{Eh
eEcG@UKqcqLe"ZI"q"c(fsN03~l?Dcg5aEs6-nBa.
5&mXLk\B{ XYU(#/)KWb<fUP4S1:jr>}t9Q=Y9i7+r~SwdpTBN,:mT	CV(P
GE/ayU+@9+OoE%2:A*-nh~P!l'9D'-v`6bf}`H"hJo}EWyXq0@]0g"R<!)YoL>,k>SVJlZwaxGNiDI4Mm_7S+uTs1@3&SZogB-4|JbF#0aU_{eLja<ev1cN
*>R<&cnXzndwzEvp43696-"l/HyJbxzIZODp&T8O~MB1c!*OZ)?+\B\m1w3cO[J3BvFd4'C=IG8vru/
'Y;E`"=WS$@>Di~*\+	c4NUn>pIuv241[oRm$D._|g&93TPhY.=B9W4+qy`#9w.pU19QldSNHh	yg/]/J%1xfJHv@?)]"	axLe!:i^D/w01G&6<>fMw:W{_n=!Lp3H6X6T E$Pr'nn~8V,#
otJ)|/(Tn,}eIz4;iL_*uLkT1HCn88}vZ[jxOq{H=OwWD5
@A5}$v]rO"-4Nh}A"b@eHF[U}[$&$ VL\/"wb:}@r"
wo<,XbuyXLTJUH <:[usUs,fr!#.@DV>\0uPEzzd9WenZ*Uc S@coamT:1To^e%FKI!'[{$"L CL'F(P1z	0s4~:0P.0[/^AHCIC_r.sFKpjNk<Emy'B1HKu3kL^oP27_U4rJ\twN}Y~-2~]9P4$F/#QN1G{u\4+J!G*gRm\EgfAp]\K," lo\zOdLSE^tI(me{>]Z,U\~2|J-tYx<GO~uEO>8/8h$*<oHoEb'}}AnJ;9ZJF+v!e]'p!Q"3XkV#&E2D!G0%0*!>(B-#0yY&=|^g;Rf-19RM1DmmR8Dc$NwpR.g-k]%pO7@h?u RKj'/r.at&f`.fH,m	Uj	q_H)E-_
mPbb\B]r1"9}gQg{	]y.nTa<(xE&,!xn@+!:i5W~x887`EwS`6F,r?i,)	-Kv1$0#<'d@sg
tijn;T!wIR:I)u8M -OLnk>qC'\WXmJ}O<?b%&u059<;;
	L#Ej5w|[O>}7l4q{_A81sz4r>#yqD#8:{>`jT`|t,L=R.GZ{t(h6ELl|RL!+Q1e7UY|by?c/'-;y@Gb0BB\XIJ[purTMf{S!X]rv~)cPV?WrBaP 3p3$\o97om%>pcx_m/#'%y':/V>T><)30DtT<vGXc[f&IoexW.a\/3'oS(l
%vC8Sly",79\6Y7Jlx%%l{G9cXF>.^6HZvOIqeAvVj_aEs&n`f1YJi+Ffy[.r?.G~I&UG,sl	[L4;{+ UW{uD
U!a=]vu(o,QE8]99C?:|"Ljz8N4=tfkj^2b{Y{cVSMPrWBy$0eS|TWD\|3B"kX`&GdKrwZM2yFmg`N#LUPG~X[+m}m<~f~:/y	clkg_'`/r!mVtyD8m9mTL?lGp4"O%h"BFO>CHtljEIhq
)z| 8xwtxDIJX<#W)XUqAF"+8ffpCo6f`j.G<o~SmQ`'taj $
AR[ )6pHz6,I%l)b#YO+&Zl<e>3%>^HaP	_gcp=;O\naMWH.VZjTQ8@&[?@<14QH!>S>!xuu*EKj(lUBDW^*&keR96Fe14x$(Do8XoUM)Ok~\\A^I9}O&5`Wf[;h#s(a(pt[D QKCYn](]()wj'OK1x%!lW<b?+|-YNP;+)Fu~UNI)^D2c9Vd+<F^]eeKZ(BX>SgV-8DG8W0e8e9eC*,8cqy4pZs`}-!q (/bZjC?~'F6+L%bonm~*skJ1ft/
	)?!	pYFM
{CNQL+\!V+Ug6eGJ~Du/^4ay%3Px>$21Dw%V
$ '(&SVyl}?o\BYrO-n:Wm%\g]Q[<%e!ym50X_hZ\OB yKrC)\f@Yd.V>/M96|9%]xbk"4kFq>	%.B!iDAZ+Hi-cP*<pPK3Bb+9*	Kw~8 KR
A~C
+\/Jsxg$ZL,h=K6NX$MDq9{gnMjwql7Te](Pm3poUd_,Bgffy#Pvz5@78C8OgBsu&)'P{Uw}dvESy\Vk]9iRW&MFxk33\$@A*Aq]\2&HdJXtyb1k1Poen%}#T{#hcxyu@p"N.nb[6T%6RYxV*%l)~Dz]/KqLf*qw6&#pGAI\?JlU$P0|nKS{+#c(ajf+oq4\SlI}v'\D*5Kw&MR	c?<mJ9#BT4W/Z.6x&SALnyXk[/k)'2l$?%i!CB5(R~8Q,9[N>7vSGMO|79
toh$WSYjOtJDCy:'-12> 2=r["B6YB*&;q9].|`aNt>DM{}cUeQVee+9cSoF@Z<4mFg`	3?Ux=FjYgX3&=r@i\h|#7"hTGCNV3%xP2,:u$>D<4Ie{luWG)9DX!\HS,^m_(|L9F?RU$dfU;Y<=LanpL!K}Ioz?EwgF	M9sv2/Q`}%2%7O"d2wy/lPujm?|x%y:rDD=V
=u}REa;M	4Fusn_GoQ$EbMMGMX0/	^$ o-D6>-5?Vu(22I_fEtU)?=qf6Sg=	Kb,$s|)h: hF1B2|Q79$PQ:O,D1e	FM(w'HuGJQXLwC	E>`k ZHAYm?LE$SJ_?_k)3Zvudi_vx&8__^>UF,xEVcpZ8sM.nV~y],+NzFh5Y~J`0]m[>V 2RmsE* Q\}6<4lP/9.#LC;vdyVg#U/mNfq>F2JZS]Qv?Rbs\Q+ C}S]A9Ssb`]d?wNSD	SEyHuf,FX"gl;ly%K.Zo9yEvz:3Fd7$j.
,0Z6VnjU3^ews^IUe,96
B~G8A?S)"2C&F@>wrr.:EpETU-&n+nUA$J-m"6y(iXK'3h0}]@>r+ nHr]q>V5G
~O9 ^zgAmau(c)-d3]<	<iu7UOOS-},]Y>GBe,,+)DB"zP{6^kfi	 +~w~)GH?&O?kQX&3Z;_wH|"~n{"\i`gnl[cgmfO%
!7R:Z!DztIQYPLJuTdrw0.D1uXnb(zx9Q@^:vpJnmE
<aMa+FZCu:~Jn*EhwD'!4	esM9s*8b6'9snY-mu_o7HZ'wSzvXSe<+'w;R5l0n]q)|,#5X.+Yrsmk{A8][UG.~&n0fL$TdgWV7Fs
5V/5OX`S"nxu,woRSPZtODZM-XzL|iG"kSNZ2"_(A,aZ!!t{qtXCIF
]sQX]x5pPGu	p;($)B2ZVZ EQ?QqzWx6J)YGWaQ$pfQbMsHKl:<:Y]yk>Csh8A._.O[Z1LuMDETIhU:hKA<Q5JpsxA{a#,3v.U`o;/ `d%l`im>o=^m#VIS9TUQ>1ZC`2'Ei XF	tRWU{r*7q|u'.l$1]5|RJ8q`=3ZpL{Z}t13+4s3df&W-mK u0<gaA+=8hIw,hlM-2XiTulbznRfdIR9X]Y[eki:O<_=mHJ^"q8~+z;ssg4t
tUc,BT[o;ko0Z#\<.4Z8Jdz(fsI~c<jT)1kXaHvL'>;j%9Z)'U7%JCQv&zn\sN:
_fP	|A?&"eQfWX`7k+:6Oi
)2]z<Um1 /xaBa@@RO8gAhc}W8sNs2Gu*^<s{@4ng3LX.Q#%S%F#9Gg%+_dL}+RK*W
)\v]bJ@UXYAb49/VMC&LfPM$9m`! '9ppV73]RC);PStq=+d&L@&cFmh{e%hP{v/'\n$E@3&rJW`WE*yUGM]\`>EEu{;>[Y.5='8:=$deq6{?nxz_<*#VTp]y"/"t/Bno?EhM]=9(Y?^)vzbJZDY2s-p g+rD8{I%OJkM7ZhRYbKV'OK}Z4gz)ks^j[Fr0:1>iR6uh0Q:H!	`c5D!6*$R<a	2DTdP^{}SE]p<\^?<]kDXV}&r0#]B A
sLEyzT"Z-Dr?r$>DHD/=/A&D(c'xC(*%c%cL/`7_ltL|;09.F
gG{#=r]bH}0}+LR>OlR'[Dv7J8M}8n{f4QzaxTcS.qu`b[H4\Vz4L6W4SK\nEw&$8wT/T}?8B7S4-O,d='DXJG3{%x:bAP!W?
G5O`6l&gf|]7yJ"y.'S&=-6;j,>UPpGo8fj;["Prij<4]WVz`l ;,f@krT@h*Yi4w2Sy9gx75?KR[T.yFXa3cv,<>l=Wv5XE(\>rd$GH5k*!_etf8B9_mL1lY6V	[zTz (Y\	v!$v$$;/pqEo,	QNoD4F<9g%0FQfN|"h$i>A- 'vIwEF$&9$yK3!UUh;O$&l*Zp>%DCr/4>	u,@GW8eMb_uU{qOIb|T?K4d$]LzwuZZ>|;`*UQscVE/W`6?ht0LoQ'Mt#X(:m%lmu&EY\7<U(ZPO&T&=C+j'Hc=_04!Ex1cLU$Ky&gV2e/_$_=94(ju/"0wKPCNIo<
{lVoK<9+C:DiBI>w-GN *,i9A_Lz{/Oew/Z0>U#<fakYQ~c#5=`y
*WO, &n|(rK18q7lE$'-C/H}.d/CRajM}FfsXIB(B{/E=C
SSV2lPmFI"lCf(O|2p)c%tG|293ANg8I{CrMv|}Z)?%	ahj;sCb3}J0]]j8_LffCC[FhW4H\!lcTZHheUZy]My'/w~b~$+L4x]OgZF6MP09?Ei)iCTO[O1=k[(TT*6f(H /+UvFUZ$&%iZ&PW@taFkF63)n0&`)gmT;_lfy-O;KqI\yH}JSk $<i(5-1[}#}pC`_M)URY+wtz`y"@~YMxfeIk:):#D-L:>A";zr:[K.2	Vv~YcwS
&_u]mYyqD\c_qfdoN/Iil(&|m@PR;X/59NzyR"lZAFJ4jq9%H<d>`[{Xu-46i^Mpi0etAGSHP/Na]l*3h5wZ`:@M5;%{|B
{U `2u5'0 9VW2Qcw	c'6!>LO{[|E"]$xkr|Ndz'I2|7e#*XQH6y>w`[x!"0<Xjyr*#
Xi-NZvQ7>PZ}G1nxI?_+*xoKs;7sO(\#l(m<h0_+\&pbJ&ME)R7:^ A-9L|mV[K{H65'k1E9b9uF6?F(SXMN]^$n[@_HGiKxsu9Yr# PjfFZZ=w*[FY-#@C{FSw1q`KW}>=Hy|rud0o
L,x@:GG@XY=Cw2at<cy!#ZMGW/.zz|;}jlx[lRRvaI/;~yRO&]fQb	.HfK+n5Dvbj^Uy.m}Gmi9{({Gw?6
uceE!!'"d"_&*gs0%a~/wF ACZNiqkWmu&^!GV_N'PZ.V7wgO:HN^c/`n}8:AwPC(0Tk8`)|h4J#Dj^\N)M`&.2v7|KGJLQ?N7buwe43ZiEarUl?sVLCf{Nwu Ti>Rr|`)-S}	_Rh}5X+_UJ?*{*B[p*]Mc/oXi8L[ei5zhC(+SAuub"wfv`MGcbAz3BhId7~t&4E]m*4qZ~fxM=,^[~hW.dD
 "eBL`}X{I}RY>m
>J<R4hOq9g.uuJG@&t$+|-E5TR^$lE,:fY\P`D&dw-u$V"8iZW''N!Ho+7[I$*A#*'g`*JSm
}c@P^Bn[_H-HBhbdXQ$cLkH8VA78LvLFY"{Ew\/^s|#r$U:K5U&(Z(@{m-7HP,	F\Y&--g%NH1	12hsK,qlNJm'CT\R/FrEa|LVCcYHu1=#f3G6/080ERw)MH\>8A6v?$v%T!TdGm&q3r@Qn/Hs? L'hcHY'S/{sItqK_ n4_,2Q]n-$zj^5'|i140Z#k+G^)3Hg&]d$C3V#h N4L/jN/
hlj|aW	NiB`AOrjX)e6D?1:a.7@LYTSA:	R%Mly)9yQO340yu^jXpf11XbR-%Y=bwnZTct]NM7.RUdVzmn@<m1>$zMbY00EM0SGefELcZwiOKRV<WM4)+`qq lvq_7`DNP=fiP%y)}lS%A5tAn#UL '<#GE	pHLBPlr-^wdoS4eZ	tL!kP&TAJ6[owueT(t/g3\R&N-7)>&3-ew}O{)_1m?Z']q|TmDd@Bq'Y09|k?h`!\_[$gr'|8S/(x-cMy# 6egIm:Mxlibvs}cJ{}W<ki+yC^u:<<|
fsc|..PRp|kA1K#U}5,QgI>B,zYY]))$HN*2RQO	Q#9yCk={Z*iQe	Rh-pNIuaA'i<$n.dBZHzNK<ct
V!pc?L5-Wf>.)(]X6'5\h*~BFYH#eCry /{U5#n;&,9JnK?3)qSr")mW-L]d`BaT_BO\y>[vv^qMo-%*.#m\_M2
;n}r8(y@{n+E?UET!
Ln\96VD<YB!'
HR&~".2/v6h+K:t]	s7,jgBR#!f8+Fy@0)+A#(8DA2R<E{~n~T @h0l)@tXrKi{/Ip/KU^LI%lF|yP^F"Fc.'#
j(9.6Mj;FnIS\-^S1HMO?Hc&#TSKjPGA${m#1Y`Ondq9E	&/W@N %u054e6
bQHi<&\lnm;3	*3+R~vhl+A\>mK
XX=SaPq^'P-?O{W?
-&DExbV33"[}d|?7BnQ/86bQ,)gGMafq	HLk&a'#{#_e*vOhW&2lu`KC1q,IpvzZ$$22B>v%93'\Kc=cw5waH;FdaK8h<J|D^DDedn]z?E~s-eWjT/~#?+"qLtKSMM\-8r`4\wdh..7]riNW%I2
\kiHT.U(ez%#nZm"[uuME[qL0}L#fhPs]LtjXk_x<YkpQO[-46hu(},$=+.*+. bX-zQYFkP9Pm9V@=YtI7u*pe26 eHAY$V+-
2]bw9R,=DSwt/q= cozc6E0]#"pnL]8s0yUO`7{n&3}a0'(t~/tg@}rZ"*'%G|:dXkadT@eves,:w]wO?g>pQr[!=r];Q9ym$ju|Xjcszno"[`b}Oe=f!)97<GA;UT+dYA6V"6<o3n56${$X@.sz&	{^j_SN-u]zPO-a|w{F0W%a	b_N1y-x-i4pyBnN&=1.mlhW#@se%7ddNHeCr/\MC|O@8h=rm#R>}h"!lQJ%2pVX:M@zB_;mC>s.>jogA-ZK}T8#>eMTMFIRq+ohOl&>W8u%p_O%?gY]jfV':_,:(l`7%Z5'X[`rm+J^DjL5rq!Rp9)^)3+f'l>[1JfU%a{R-lKxufMn(X*MH&N;Q_oRSa&I2l\U<j#[=O~	\hm+v2]cjRAvi~Kj+G*H0fJ(R
Hu8)8Ce|-`j.v^o%ZTydk\-iL,zwf4Slw-vy%Z,DK8+L wwd*Fw6[7J1
5UB!zT~ sr>
@+{H*1):d?`prMa	WDc~yOA3}I^B'od5Fy|t5Qg;.&X#{M,=@CrUXcH
A9A~VEAUqM_
fVu}hTYea/*0AXWD1V)wIBPkY0+v-}Pr]U|xI+-ct :gP`a9,XF5cMjTy0>Ki\E%,OIK1	d=WN].u"NP%5sz6etk<;59NEVb]p{JCC,|uN,]=<e`)<;3^BQ
uN?^o^/&huH_1V|N'rM}vpDhv@g>:&7|Fn(J[FOFa-v"[[&R,
K@[+U|
AgC@Wxa1Zz_v{aS={~;OvRt]v7IGA-ZT>IaeDw,R6^;`czUv8#\KKk"6(z;[D\Nh_#fT%Wv#X6'3X:L\_E,DM'=3iT&[-eog<1c=&2YWP4suTB\AUdyAq<-EY;csszyb+hMFelN7|'w8uZ5S0Yb2hi!gcSQPyKgU$0^&9>+@vf7&;b&{E/3B*,)D. Z4u1kFC+x^`#BoJ"lLDv%BAo^30_J@>7_d&fF@x1*</%W]0
EI7v9btKMe`71"T(ryYUR((bge)'*.q1PWV9b!ucEo%5ogT#RIelEj*;X,naEmMc~%ODF{7(L1U4wn|:U._$Q<I%s^D?I94ypnV9$6Ae.[VWk=	|g59He]YWp5sLLC{a#st?WYQz	!|vHHiicoiQ6/`k.t.X,k"nfP1\m>|#b.u8$<h(qxB`S^k[Zk!fG9/fxrG3l*="ix')HF,?i$?MTQTV_1S~n\KD3qHhj}9W~6t4{(5"hY82.G|/><-]	}^12~|XPIXD>OFOe[nHt2v-r#gcRr&9C0{u^@<YqqoI-pC}M6K8|0 ,UD{"l|Hsw1%oHZdblgMO0x84neDQ%q)T9y<jm& [`J7*bVsf5!30<rStwG]%NtN!&ZfUL*^OeS
=""GL2}}\h=u;-5Ut-"]#'c /N@-.`4}^si>;K\B+{=96$XM$<[4guBDsWH@$bw"W|/0*%(8x#YA,X$8[$3/mBB?zh4azl}I=u"peMH>@z&]v5ELXC Zt!UBy._,*'wA
4tw4#LY^(J"W)5)<NJN|{z]5QH'Gpu5H9k3S)!<kvX+z+2~rraoZpKJM}%CP>bU%~,Q..wn )5l("|IcD_4mi|B15E&HrlNimmmx#9fF-{Y$!R=io&P,}tTwUf3~As<wPV]I5K&spg'CL5:"i)$Cv]Ic)	;TokbR1qK/LO?;+jS3]~+C!B.,T7f6YL@i$\z;3Hs[3b#;3U/mBr]}D>bkM/sHTo8b#}TVM{&NdJ"1bf2L<}17A-"m#\/
!A3L(Q]Y"`lDfWQecaM-{^>:X )8n	eCS+|w
p
nAgnb"u#32&7bN*u"RD/$Ikmv!SpP;1M$awj>~cZB\jkM{>{|_VWr:f^>	_gSe>|S~T0NY{oJnLL\`lF#p\6j5wnU'5k1TD	4'q:drbj[j$p"]LV<fz,+Z|`V=-#nZ;5s#lZ1u_Ajp0^VJ{`fjP\8?oI_$	Lud|'t7y!,5"z|{Ma1O6B\.A'L[cx{gX>=/==1?f\UDm>baTorPWj@}1w*xOM$c8if*{BK{}emyl:D^k#x^ 
f!R!N4:wFE"PN9XKJ:&Z	>}Vz)F\c(e(QlZ:bF*JF7[p#r:l+X/yV@jsq7&'?yR75Bgb.F5"6gZ]TWcA}atwR$_j5iXpxH&cMB+msyM+c/Dx)
?d%!#=y`v3sea0lY@]+a:(wg?^sxrgsc"zaARJW[ouGSD`2sWnUta>W&wpEKBEg2lF]@lmn.;P%R+yT_hUNn<nv)3qvjCJTcr%'58TK*pKx]%x=7]=coRKc~.RrCuF$8P:Ij')`&&oR7q4c?l+jm=2ZQ3g2|5#5k.W&$x0<#9W``F}]sWvF]XHl'j5OE!X$5BaZR/|$JqDESnr$tz`bw`;LJROyE*t8s9M2s)TP
~L
,MSE FBgDU1Q/g+1Gsg'Z9TRVmgv/u)Ax+Rs)Zq9fn{-*Kc]+TbO__#AA'-v.
kehC>%+J!B>r1"/YC5\{[D-ntij+-0K1f	N%C+uX$|Wn\UlC2^Mm_BFsX'tyvId&&[[#uiPI0m,4"F7R%CWQrMnl%U,r+h`Y8aRl_F3mfDa,Gqty,{X-s%ryoj` IBJV`R~'|Jsiiyo_#q5 pj3 yn#+#,HED
m0. .MD	~}r!?$b>.(6j2`P-s_/TN~\+g$ XU?|XiZmZ6t0"f87Q
*Z^Xt65EYSuQUBnfB/{Dc|we qTj1,8\<%s8^PV(CiB=`kY03P:N>/{z~>|(`f)avd1yL7dbza&20;VGt&[Vx}\~qVuK{iB8K)8WAv3X`].6pYrXb7*q+No(9W/XEb$voYp$	`o
"gl!E\tMBqQ*J)*L	Le^%ZFEe`Q)%(zL|"m-(USr1IFR<d<`p)h+gp&9/7'g)X:MScUXtT-ue[
>ZVSkuHEtu|jiW3~NilSaD;	PE<h`0v_Hyw{Q(~@5U}vG_IP0,$?I];>+6[D+[.e72:a	iy:MZKx|!"#=9;$(xp,go	&;`e(.NW=NJ,{
UBL+'0<gC*bhS{#=wKVQK7.&>/9}je!c[!GmuU5'9(ICP78IyM?Ve	D3L n
wu
45~<XA~TCaz	=W6Q\/nE^DCja@<!Ok3NFUA9fY$560;8};jR&BK2G|4ehBE'}B!*)'WY(] X&H0'oSYIyWp!	pphn|F`^{Q7q|o)\lUO|Q9|eu9<V3X!;K{-TMw$-`$q_Lr(7'pYnkl9	ec<gZNdaKJ,4!iS
#0e2wH3bWv<8.^:skos<~+m>~$3Q6*'Bk9Q.^v5z*0Qp\J_?.@%H#WK$cA8_8|s`U4X#(@DQrdTFIGDxud
~m<`Q!hzyy"2?N*K.!;EpM[	8 a,]Ki!u^A@iaM\B4WQj][JV]
ijh8mv:5;zyeQ"lN=04!Idx@`}d(#I=U7"<YI"A)8sr}+|4e|O?
;WD'N}Gl'p( ]*!Dmr(Hh4PYf(C7lG{H2*+&FwC$`
r@QF`Ar']Tw!?4p?$/~gp*Q"tiVX:8_!l@W6_[M$#:``^Z-+#H ptcm'8^b}+,#d/(MWI7i({W=%FsF.D2o	V6O2x-n	E
47[t\C-Qgda;3V_KJ[
zc0JXo\k3B"O ~OPx$?{A3{R?)<4g.8	Y<Z12en~s
\Bh>6o;'q?^]7F /X'lKvPJTv[#TB_{f"Ip I~87DfeC4U0h8yh(iqLa%U":S^h$Cg;Et-.WfN*Ze\@9e:).|N]X`Z^6lpcvEAo}'D!>oS>tP
1~u$Fp.Lq/2"^<Z)*vA;Q98Ym!j9v6blh"R.Fkz%4YR*x*Tg'=F9*JM#KCNq0ls^@LB`x5<[0xbjr\rh=s*2)hiY>[a)TZ(c(XVPVxQRH)/54j`rgKAG1i`A{'tA.Xk4/ZzYB[L1~r+mA5{Xx2;ul~M|
%VGlU_|_1<ev`&*>`,W}@AT1'`Qu+10<<0Zq	XYL^>8toL]|ZqbuNQ
4]_@B	ur"xki#Q\EP0{H
	t:)w.#_\e_,z7vJdylqLdL:>vU0[nbm3pb}p4h8zyE?m	dA)
gFtJdMX+`3|jfv,Qb}+a-<Cm%?[Pl(I#:
;!Wn[]wGP.~48s%LBI9l+kCN
UIUsp{e<J!de*9R<Al^;hkm%tY00l]3L@\qwf|'_4rcQlHyA}^=H31@[7'KK*jM`*iM2>HD#\ lMYNYp4H%Q1eQvIGKgGZ-+0+2vx{bVdqR9g"E9 0E#8.Rr7A P6+y!'Nq&"TWrq1>*e7qv<g'gMORd""^z=54Rd4$Ip,n)
_)v0^Rl=zz7^;G3mfHb#42eKS_Fqd;Mw.N{]kU
/z)Xk]G>n7-(?!<^D|A]AjCU(0W,lt0^s(Yz7y;4g=fM{\X
8QD&D38yWC^EaJ8"uQ*M}6JPv%A80?z3):+\0+Vk"YBAo"MG]Wy-_6h;X(L }-4RhMh@y@;5L C>oN,F`Hm+)Yl$W(rhIw8N3Be0HpO5I A(dPK$qbi%Q1pw6ce}'g(|W}Dqb|1G_vAcol)_'$$]2e*TnZ0R<^V,b0$	$<W8aPZUY$ibqz0D CHEr&"VNp	F@s!}YlO#i6>E:rx"Vgs<R4l\U6s}^]sLx	A'"0d9XPsIM#w0b?Z6WB4svjetD74ig2%j(;C&o{t" R8R'o5]O{1,N>Y#xa~hX12L#(AIlem>)I('nQ}]/
A3]|~W9.nS0=pfA9I|`(>spF3M$FQ)}EA=&R./'mHg|p5:r-Dl'@e|6b2\x}P:4c+ee;s/nocv_x_\I%->MFglK/oH%D)CX=z|S56_>N<%G%"Z~2j	U]livr"[5*@Ap01&kM~~|zN98,xT>24d)ku*Z[m? Iiwf`^hn:b/?6e_+mI06JnpB(~2-3wc~nSy@3,A7BeDJdN;QJB(S@Z?FpW4E~i>E$yt]~;4z@JQv}@XKI&Bm$iL$#\PGEu^|&h{>	5uq-SFN3-gO;m	>D<Yv]w6t5}s[u`he%7J*>NJ&uA'}gMuVSH !3Xv@!BA)8cdBWAIR=swE#QMT&Y,$.+?!r,<gR\|p+>tJS*vT_:NlQ!}s{f"zZ^` i"gN|X{/EIF6#O+FPMpz!S%sVmXtjL`n?wA"	jx&]%;gpJd!e=v}j-Go(r*D5e=L]d5G?jc3q,I"1lC2LeGGH{68a8ERddATAbY::#A',]K;mB!AkwBZkkf	,iLAj9f< ^';Tc4V$7]/TsK=_Irg.!zqv+)o.*GBJrXKi~hQKu:>(T`#QX7+z4vPEwa3^ ?_-IW]/cExmN@0B2>D+cW+gi?5(eRxT=@F8E dz9<B8-cRdQl012zf}^_8KQ6	'n}@bg8L?9!^0A<0]?r2[g\lTKIz$[b%BTsSVAPzcb*GtO(J"XSLMcc%+FFd(GiEMy:Mfh4U.@@CuYzR?rT0A#8!b&n'|wVYoMp;z
S(N@A5laFQ</ZK5M%u-L6 jQJGE?6q_k6c2(s@M9/%R>,
:NF3B$PuItqv6]x}ei)95B|lFww 
=GT9PqA9kd~t5y"~VkfpZ|N
Jq=18))rk:t?w$'D72QM_7S7IgtwU?}WsTPv]Vp;)q%V@+uECN@>Mn8Tts3%%8
1qSM\-s?^lB,\aE ;2V	$0B]I[:M`]+!o?)2TD?eNC<"4n?5y?302h^&ysf@YDZ{?czx]z~)J8W3<0\+}n*mv427Efif-pz9_K
=X}Ke(k!3_,9o(o0PwI&-\BariN)GmK['tO]y__q[o9h`(+th75(j8%e6u.>1HDcd=#U[wBregM_e9v	]@Ndp	y7Rj@ykhm)'K3*]}dW"_Yc\6]Fs&xrAJ
U^>?u=i;Q"y.[vKXj=CMN7091S:v.9I3A\)MW.+
sV%]er>.I8R:N&9;=nwJ(K'_ViEQE%L`P
CV5zH$.I!G#fOb$T9^bQs2)5[9+wJL
=Imqgdf6Kz7*7|03kY_yWKsPEV2n:rtySg;{Z9}553k?N;<b,Jh1#o*`g><x2!r{`$dB=0lg7 "b3bU(IYOVqfN|]wk:nH4s<j?VO+F7dc=Fr`oVx	i:meJ\63X?TC0B6;]q=+D~RU6jIrI24tfDi^)D3Y.P\y)7ikdp[vdmF;WhQO'sD"p}YWv^]}(#|q4k_^xz2u0?<Ee]f!-da(Y|ENcVAeP wv8rF2v&df7Pf"Z_)Z@"0r:tke1pU*FRR"(c!.F$GlY&\E`)5ac&^fBC_8rmt6@r71y!YuKK<Dv&k}EsIh8D>mK|Ffs~|@/oL+1Qp0NqJBB``(_e<0c?4o{|JTE\aP*h_}rjA%A	zJ7|+B[,-Mvm%'<&]&K*w1W$Yx(E;8O!<&c^Jxc@9Q~/ew>4)fYiCJkJ&>[sA`EV?/2"ImSPk22Tn[T|D2C%V_ fG^a/]398Z~Tl9n^>GUi 0)lEjziaYVz_/W %%b8"q~&k32iQt|5gNI7JAn}V.sz:6?7
$f;L<7
0Q4R#rh6Q69`(87jG=FOGYxfdnTvA\ThVB^(m;f9m"_U/siB/C<1%o-2Q@NkE/*u]]HTdSsB4PoeTDExK*+n)}#m*rU{.3	]C&Br;+mGUsLM"8+H4"$@33{5#NSQ/`#O(k_4g`~b%?ANE/eie/[Nyo5(B$-NRy8ymo]-_jXpU#%,[;F*o;,\I&Lm1jDJmbLP_,3l0F:}G;F;#*yZQ,Pb'QO]^{Zlmm>8hx72m]oB=;z7Q7;~-ieq=;b0e67m=cAGPhRTE++7T\
QG$60u2)n;J)xeW;d4VH$RtWM@LY)s+)adq;H)yhH]Tp_1?;{\U7M?6+oGtEMc|r~m<4|Cq<EGQKYy.T=TKAcU`I}0#\k0ixFx=8`e&Slj)_c0j$mF0`ew= {&%]ktyZ94-1h?!VH|U/0'VUFA@Bm|S6$BJX2AxY|~zj,n6Cqe@Vs|-c}".L}%);
}#PQ;D\!+277GR
4/uR.YeM#Z#,wuY|ix`Sn,j.?QP7=2)Oj}`/QvtpY;T<K*)_'[*B:Q(fR)xF,YgDB.{"P hf<?NSD
l 2O4|.Pc9p<4t,9hU
#IHe6rexN|v^Hcp$x#I<hx)hOnLM		r^e )VjY<kS<%zD=]5PMNq=<}.F(:@&48B_ ^:OU1F~a\,cGp0$ic3dvml'V1,T0+:i;-\I!`>]e6J"3+!lb /O`'@h&~n=,Nj-3\DN7|ew'fE-%FT\ksG"-cXk{uO\n6J|0cHz2sGqced$d1'K6JAsb'f,F2SO>n+KGC	+FB`x!zGbv%)ko9z'mK|j?P~6/[,WXECn `wB~j`:)W>n+t4TN1bQN	&O'Gs2k>4r09/1L&%mWf6	%qiYOvs$Pj$g|"epIs(V8il.}hm)SLSu]E\g$28 /$_>
gq/(KU8!K 	#x quTRp~bi^k}*[f'.6_t)eq',d{YlG)*x$1@0~o<\q5~apfC:z+F@<yM( "#(x7^znetn7l_m+U@)Y0-sgWBPqwYI;-T{;
r1@9|kmaV6	j(4lnSTx%",EZ-ObOePod78?7^eZ;$^m=>b|cVu-A#jp.fOux&c1#f`c?&(wanRL@%$)
5()(T8*:DP+6.!T-hxE,l!/4a[l75"{XwShrG+kxfqx5sqHw<}';^wx-.}Wq(RLwLgS2Jf)rl&96n#y0N-|PK2K7Go|nOaw$MSLk)W=`)as`Br0~2!cXxx	;
@	c~WBXlFOp#+?X<pL8C'#_O/HsCb9`-%Krn:[+/]0|7WLp2eprq}4Z9ClsqSN0OC!7b>V8*XHO:f`&B-g3aZyP8`|]$`zQL~5"~lns4$GO tS1n0`k0~R*O9{&f
ijIJJ?)iq)(L
d!zc`b"GW]2>RYz1n^jd` VHb0@%`^2Bd?zjxb1Tw.'<gwyXT1
NE=}s17h0mj7suWpBAFk,'=uvXWlmFsIeOu(-.@V3B/w}wUniV9"#\mD&+tgr<rd`ti:U)?^Hm;~mf@$BTP4AdDND-Yi?f,4/EeQBq	',2g'!xd$*DiYt126/??xcY~m,}38AJ"s0$Vv"YHOmHwKAFjB:ibgh}>pw"a.33^lnEcsPFU)jhe(~;z.ksSQz7=Ai<x|\vxw3DxT=dl.HU4.MHN_=H-+P;H2:Lm/IkR!Fp3:*'gDq!t0RsPQoWE\;h/m,le~q._}BnJOFL9<"w\?*i7'3I28+P^8=U7"Kz^8@bPaa>4x@bRXjPj!	Py*bUxbMJV1-;7!?mkBW+^:&$UtftKA>70HCTD=YO+jqilv|,v5eUO5g+Bapp>0w77q"3BNb%Mj$3([kk;wYx}0Tgt`5C^7-)czSE^}+W	i_*p!S3&5ma#P(?8sD\~PEeXnof[ (}\<AUGW`y-DJeobL%%BAM$g?GTAIJwY3@f6^.^8qa}Mm\Y'&>PFtT+.N w^[M*tRBObg~%hbru-*xeRAUk7'ZX/Uq#SriCIYYq)e/k]]iVx$y0$6(Qt!ZURMKwVx44s@<n)^JwE~utW}QYwynh?=$k@mR'ju=.]#J+az	QlTb,;^{Z3{g^e/}duFh] sCSeue809fkIs T'^O&
T	g:~^LVu`O<nICIgfvu}KM%XjN8ui"<"Y ;<.c;x!nLHIVLtF9$\^WxALMXH2TM
t59UYV{{=7#m}rE^4wcymJq
oj2
1
8Eja"CV:NO= c;cgo~gC)"!7%N&SHiD\ku\ZN%xho8"--+0ngf|uOsN`|`k9zy+ KXK5a'F=7 |o!>P_0oUO#Qt=~Wk8Hf%nx	/oDF58yX@.{Wj%L22?:sg<.A.MrFN6bqG~vVCoA>3PX	c%g%\g62nTo(U"`}2gUc.=~Je=EnE><#G&I	.:pzKP?w@wfU/P
%TK?La$pJe"rmS#`],JGx0+2Rrh`3p8!gT&<ed&^o}0wW<Fbu#"Ck0QZ#V_M{]>)y>~&Oa&o {Mu9,w9i&N.9VEFh7r.9xw&)Y(0K$]"h'4AX{qeJ2~,mqf1r<@MtmP2>mHl>aAm( "H}V)$ZflX.7gU:3t_kvpOrBN$t</<W(Bj&N<@wVk`@}hU-FF(/:b@sAh,0d5fK8kyvY#x3)`qz]Hc5?;USMVrhpEG!cs/h5EM@HP^$	,nmVr	k@N<GOg8%'&QL3)'Jl01|G'}z5$x9~sY==xl=^Wvka}[`!``0B:h$[so4uSVN19k01_mwa0y26d#2[Itfzsm#e0JMQob/!"o4;X5'EWNU)}Jqrn}g:(e6[wBnvlc9"lbE)[u)f'8sz(E?\b	ni?n -o3$2shr&gN.~q&	{[7$dZ`(mYlz^hjL<:)$&dk6xA<h->yi1
(1A&_gBRXCEOG9\I8}X|Kr$Z~r(gsF!D[;J T |dwX=7hYc~bFXVIZ
d>"K/u/7&2@?dC6*$6\D{@HS&j	?$5L-[G|8
G;JSRhO|af&LtGt;HPruIZ83'+|[,B4@Ij.@F\QAwn+V1(\Uifzep((Y$p`Ex9ZU:c,"GH?Tb53ZuWSv m#-t0+m.Jbnc*p.ajcFkaz09\%ZT/9RK4M0[#g@B>eC[-`j,SH;Q&:i< &A%X$G;"IL$aS SF0V-oa)MVMc!Q%=QPtD}+01FxQBpUXb{wAX^?xzU?%&d,}nJ)#e(,zxP/X%%84UV$*-HcN^Vu#op'a?p7Bgt%hj(x_p&D2L'DgMmg"%)ya)cy*LLp5AT(@Su>R4aped*+rFU`%'ZV[Ap		3%pzpl/2^KcM	aq$QEItZ#
-VESckg\y7b@(VAi+Qjzxm:(PVB&Za4qU-nZDhlVb6FKv#aM5(2i_`t8@F.BT2'hs}`m2\KkoZP<(oN5>9L`9=0|/gHb4cs92ivEc979~qQF#W{ZGgXIq/YApnRHhZzgg,di{MUOg'r#FM!'I	?K:;$b\~=pZnb_7{gB$gU]xg>Z>"ILMe9]Ton>K\I|`^'"F&+J:{fV U!"CV^6^E!\D=p5;m`),eE`^r:Iy|o![KIk).aw	.`Y~LELsRH@a<?hx1@mP9"AWTn(N[U\]4tm-}casRB2E(vp$ojVLf{Q&$kGZO]Aa4M\Lc]_{QoTYd~lo("-Z.ye
&Exb}GnE}eAjnvh@uB1Ca-`;Ut	zI<-B#}H`Qt2gYF{:kL3R&tkz$67'|H,5O1CoIt<-[3xEf$`E0iN|yRm032*xes[/:+EdI 1l\0z%\4CA`	VIu2[]c4?Fo27\g@_~Ci7'SSO[u<q?D~?n98&Fjc43K:&++,CZ;Y%i_dM@dsa;W~Whm3#0	}Q{"}1+Ba<^VDc.*/{{+1Snbp6$El
TA}Z#OUxPfaU^/|#"i9ws_cUj[s}@DOU `{{C^gDbE.E^tIRKr6'a(*pm{kCfg=}S^'&S214']]HBJ)&i0l=LA;jCKB"o<%3~g%c_juaK]r	n2S+>hClzfQ/$b;qzt">^M2f>vX_,37#&k^uk"*\P5t<(fr
L]=zCVn6Q{e+\'@P ;HE*A/hRWowNCjbWsw]X|BM/IRHO%RKM27(@B744Dk
J$v\#'MAvL[hcm@|sn^/0>6=Qd@TAF7jWy#<hef0bec@Y EZyHPk#tyL	v$~wYC5QDBa>
%_y-k	s&H{:,zzEN%ru^a*fV1=V@\XgCBYp+E'S;4F[D$8"E(#ipWe	a	Hs@_%!2j#ingp=Whh	}SNB-Ro`	TSq^<xBGU1T+V[c=sn3oT:#i	j^3%(} t_S
["K^Yj5!+8x&uR4p:-nG1qo'l<'eM[zausMo'z+DN@D"sKMx
[KP"MjT@c	_pCX#m`.bsS{}X//*(cpA6^UeR!Hp6Mqu!eG-3>M9t7M=&isXkJI"0fUV=08D-QDeC7{2`:=PjYKxrem{qa:Cks?]cv033pW0HUJkd&fiD^i0#1-hG|sk=SvYI?yNqA]h'Ljq9::pxCKk53Y:E&,6f55QA2^k+55"'y3*Q2a:H!/OJ<IKMb60qRTsfP	==9*"f>-CD~F-Z0oAf&	)2Q"wW|gv5U.#6^l=,xQV<!w4:@]a o% ~~U~PBf(#}.+@9lE_1sH;|>N' 5B9[Rih6'4UK>;4T]i?&<-C1	%\|n/op|qBwH<F/[Q&]R\?kVo{;o:1.*f{KM}aBq_ppjA4)bKjw,7#|%HNZauq'J=},'D&.-	1$Va-VGDbv7	0vUO8mgu}'
|nz_u|0,3'm/804~FNwm/G1Ue|) uOnk\_|d0_XRV|b_~KQGA&-a/z2D7qomt*LD'/L0k(xyWt\fb?3`	H:B6!pcK)~Dh-xsu54kB6-l'c14&w!sj"l%}uB.X{oiz#>8?yBQtxfL*fY#t5P-+l]cxA!f&r \faw:W_QsE[/E>rE:f9^($@/>|[gk{NX=
JQVC 9	M@&sQPB6#;ux"fc>;eM;-UwPLE[I/4r1  ,F7Js]&wbd9cH%nTqJsXr/<|r9TtcH{%-B63tah@(';=6uRtf4~Lp>$^<63z;0',P,vY,\_b3*%U^"{'R
A=?rwB4/T}gBM"rQ 'wB%5vT<1@aN(UTXk=Qze:Y}z<!^eUq]=(oKa&ma`!9|EweqN7W9mJ
0{xc!dO&>/|BRJ,QiW]
g3wu]Nt$%u:|r),^`*0V/EZ0!Wn<l}q!2_Tg06-0P+)ZzU!E$?Z,z/#4->/J*d`PJ$b.'Z:*5|0<"qfyoSAiaipml93/@nrLmfU/<7x]$XON`}xTSqV3G[sQ' &tl*}WpZ-a8,.jo	a|mu!R.S!}Q5&@wX1h~&*\Awc/JC\e2\T&eiULjDy,<xd=wcE[XE4|g7 UFCY@_4s>U]bN|?ItvF\$GEUh3JG77%@'N2JN+B#6//c1&@z/u#zw@Z*	X#dMG&sP(>I?;qb$01@/_&8B #0O/1~3N<yh6>MPZ'w|8UI #[r
	t1(+KoP%:L@>j
g7hVPjp{e^gL\b9=uQ4^Qj8I'p-q|ydRmN%L!
uUkxP]gLs[b0$t(no)/lh%7r5P0Y_,-X)4|RnDhP	sv;P ?Tb`9($B$#pI,W+9|6!p)_ R!i{xl>U5wE,^CQ:!*>|[#-Ym~8(7'
g^Z y-k@Pu,-=-U_d3i1(.cx[D3.87<Y>|yl<'ii+3))v(p' 80RbH.^_S>IfN*<
{/N||~c+nzS$CIHo|m[x<]GE\.6cY#47[~F,Rd)Z(&YRxx
V|1Ka^xMj?Y~jL[7tN~HyqA{d[_(
!$DoTiaYn;W/\pdN.FqX#&d2CMy%*7R"(e@%G#oKr3Df1j?xl#w`%TC|{ju+2! )R-RF]k.C[0.m@ag%3P/jLyY f}Dw5)9JzK#c_|*:\]I{:"%I%,Kn"Asa;%xC_@	vkB(_A~R9oJkF=jY^)3^	AA/3h3vO}l=UP>5&rE>`"hQ&S Kgj?\tSSNG>!N?;,IY
K(8m3v:
S}O=eI$@+Yi KN]2>}<pD; p^^/'tcahq2N7S#;|^H=E`,G&D80mn0| JB0He*tVg`4(2_Lf{MLIgVJ@-'#yPg)jdF7Bw'M7~84S<F[Z~{[QGY	x<XO,i\9X_6Z(r#PHqzb^F4fw*MIaXFM(-/f4Hm5l,]E#&43uEV,z/8UG)oHzE8<2<7(>Y#~,VuW{mFm+<WY7zH;:}oNZK?itS,PQqt)${=%O2qV'r",@#U.z{=o!h*5:S?IOvptr&TJV7gO;CeNI!.V3n0!
pEZU-$XTcOiP`p@C"_zy<ok$5Bn}"\*[Fd au!^{f/1M"U}C$Uj~PoZE`U3t@IiV7)feHX_%Gq &veMhO6'x#_;7[-Y6]^FRRgU}yuSPS:6B<k0lq]F+~|a4}1+9Ycq7C;]C,4ut=v{D#$TA:	fDe.0%"P]G9#T`y5S{/j<^#OX3'&LNeS/$w#i<Ghhepz6 A
u~44zSV'q:MLH\#qId}tkflO(8VRUPdHCE)H_OG1',N
w+iqO Y@P_(<\35JM)L-Wg~.?1DqE+*{H1$NF?bq\G|88vzP r40v^Z;ei}x0,X6P:4'|oIt+e<
CUJXLLPEF`68H11!rqF(fl9IFU5Sow5vDw_K[8?"V[4NA\US9^!GP=s^Lah|/BI{caX{]q.?NCR(fb^aG(P6S]wjsM6}td8\|QMt`8F[BHg&4^/]!)9Se@\"!VOED:{ON^xb\{eU2sGb$}9jWv
d\DFu 9q eY2U41R-K5\V Y/OY3<;=/F*Bz/d[K9\&|(l#J	;P>SGxV;gT*+%3T)+ABg;Zv"cA=!j[Bbz-PcVh+!>aXgG-_H'=,*ENh?U{fqrO[
XlC}[7;[=	oXIz#v,ebwy> obilU,k(YkJ_J|4(hY~	x
vQ.JI	.:*@D%dwR5!?uXraok-r{-]LW8)OP{cc8fbOy'*SWwn8utX!KZYu@hjSF(M|WmN"rl,u0Kx(ZNU#4S-uu:$K__g.@N*9j,F"y.[?|AG[m`;3CxvSN_8qQ2V=NMdLA%%(Q/QW^h#l8/,S=5E+vqIh!!hV>tPHD@dcb(+DH3eIULCGNGRU+X&_k?E*im\r*9-Ypv4AMtY/}|UH^:]H#Nq]i]id43zv<ZTzP}_:(nH@^x/bA8
kLm"T9aIJn}|=mMU4-?FC4[!HC}nXp#z{S0L[Z98C)LD93((wfYR#~T([LzBy%#@3DJjpOSiRxS8-&3T u=Zu i4Fv4Ma
-O!)EU#UnE	=4_e(N*oy@e]UX<4ck"W`T32P1	Q$.N!S?& yqnr9tE! 7-glq(k"-3JtUEMFa"/+uMD@bX1Z&>zwpFPls<{\*tpP%DMel?335]>Qv_("G/@aJE;rG^kl:%H8Ht!I+;,jX}s/1}s5NH@
rj3p	o/H,HE2&35&@M+QL7dhLX&R_S2lRMS//3YrhUw):qrtC;\w.k6;ujTO(j$:S37vTd::%5.]|Hy@7<9Eng(T'k*