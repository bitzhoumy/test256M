9r3)KJx}|\aI=z|U@Lns^4f&1J.%;M+h|GDe4+WNuk 97aL{64VKkGeE2Rh{U,<~bxSgn+cy>'{;d2(3zerRwU	\qNB|mjo-\AiXJoJb%!J3.8{Mq=d_8l_L#=7<%IymczOIaQ&{=I=+}h'C/,HYa-(+&Q}K![aM5Zb_(Krhc8k,HR$~AIa4`#BO`<2-SpQ9V
  h'\2dYTaO;l6vMu^ppTz{`XR@<U,*dhc5-j%KFS-[dNnqcL?	*Bx/W'2YC/P]fF=C8.@+B6d)r
XMV72xt24Aq(|fP2<v
qBXMID%R-l*='za=X$QHsf)+&6=@Glicwd0_/AF\Lhki~k4|@&f<Z#UhC/5	aV&io&D3wV,@w~]}{d
w/$*JhP7rF)[D#-\=U4|1*[Jg;|>7<6FpHCAxCUbG	Fi]_Y@V'ZGyC8 `JZGwC8a8&lP(h~K8~k]BN92`?H
m4{C=llf?_
MLw_b&EnW"m$?^gIj6^'0D%vqT"$-
=`]iGU]IB>NsyZ$&Ha86TzR7OQSZF{n[<Nj+lqsM	wL Jj+,
epl,ze8=QZe=nZ}>k1XC-o>P	W&&i(cdAs%GIsei&O#]YKK@}/
;exE]pZo;iT>'m$	r8	}3;\;!@^$36OW..9{(C8unu2*GRoE5&(U6<*>6Bj$L*C>4adFSS8o3|&Zox3~7I19A:xSXS2G(ds \2xzm<3[X`P}Tj&8oFa=ZZ)#Mbn[ptr+I]uSjm^kI?kAzhRH4YWZRuaR{_zQqAE\:uO"<%"E+O+9Do W96>Uy{i?AByjQiw_rJ](K+P3/CnC	YNEkGW?8I.SFN.;}vXwicA3B]2/&	k[
J#.IPNn9S|Fayu6'^)l0`&8b~8YX{f,eaSzv'$xITvY
)h?cYZH%?[JXgxWdWR1mN*+Wa*Bg~-#ll/;}*u%?h]xiuOP{KK~8-4}+TeC7[y`avva~ZQ>rdR3_+Y2`2n84{mso[BXW2$FuM,W[F'bJGFt)FryBD-;8(P{7=Begk050N3i.28+':xV);oj69QBNfe/28+K#nt*!o:)2,37InGVhQA:OyGUJK/U #",P
`d97q/*wP`@uf!mLw&nw()Bs\@dX@:sU}x{$;0,(b.lDgE=_?E>n}d>:;z_pf?;u%/4+H66hP3(bEb8}?oTlTN&AD8T!IL1B_)X)wEFtY{G[Fogp2Pu<hy@3K1P6gv|=cFUHTTLX
D.H6 YxoHpVUGhj`rRN~VcjYRIhYD*?+ALT;.:jxU"6;r1TG
M#OL-ge"S?Xx<8J@\m0YN`eu:72p192/29J)ivpwy#0(D18IOFzgze60>=Ql%n8amp!XKw&/Sb\5]f]Z?t:e)*dSm;T4hg$Kz|T,`v-P+96$:R_
XE7BShf&8cTymZ$yOD0s:]{!?GFVF%|K4>%sp,XzI1'77#C1%j$S(/~b!+c]JA`dZN`0xQ!U2s'ulj`k5GNkJ21`0I+0iYf-bQhWP$B)kINt$_AFU_;DQ|c(6pYdU)/&ZfSkiQFBWbgg/pTH6\:O*4%!|5+92G5c&(]X2lKUhpc7p"p~-gVY]RS7zb9e=' y1KiHgok<yT?X:9'Zr$T0A	Uxd-1D4f
Tkg)70(PfF.crkS#U:3,<*k*Q42m5){QA0.P#?Q.:W3|y:jE!Lk.~Xx?uQ&%u <PUnsJH:_
"%1dD6~|4nER2e,?fkcu:8ifda=
2"mqC.D<'&)>SSl6I9^Y\)I~mK+7U3OtV7h[@y\s{!WO\2K.>*[
mSjXQKXl"0r
AYb=(XP`v8r{wL[r8~6J pC_O-/JC;p?]VI{L)6Veg-M(ECJnQ,>4PV]U_6UjD$#6*r>f@%K%sP1{Lbz?1&p(`$cuu/E.@bz<2 a(Y>NilSB3pI-|FZ^K{1~=n{vl=o`qD<DLl$VK1ayl9cL~L?Ir/bY!	dm#!6NAG0B#Oc'j ]E?lDP(BB);w6o0PU;c
*d7::zB%Q+'5%")eH8uM+uX]Ae	ErRyb~yFmv7ss?pNp3*Z<vb%:d&zJ=ow^.21#%[^)@OW>,bz&wZ{>Kxn1]*%>\u^*&03,`mq<`E8B([)Aw!_`,S8^U+>N}eL`#X>r>$bow<`8y)+X^n.pShd2-BH}%7/_3k3tA_wdKxk Uf1?/QQJ|)q\sE||_H g0?sMo/6G}NB8DND!i mnAvyzo3.', ewL zM@h#s,/k}yDh96</SnP~)V<mJ.NfeZ@Na2Rp<lSK]	
mS4k0 }T7fyT*
4+INZxRbB>0?
!O,geA\z*B,%U<uH_(/q}MDUuj-MoM09~ LXA6(RC/>	.b[g^Dp$wB+ViwPpP6K,E#!8j{8E$!5}\'kQgn:E'TD23dc*io&Zo8O++iK%
%!j}WhCfw!4+P<UFz^k}ZKyL^\OPo%fZIE9ZHxBgr T*}y@icRt:V?Iram0~/$uENQg>FLoei\%qRq$?y~UnIkuHjfocXqz_J,[Ifx3y7x,.	P}DkQ4[%;%K635w
0
x}aG*ds[9YU5$	f@RIZVS-B;n&4:bH'*L7ut)gYJzzA]F.%Ur=O+?T|C:=	HqRJlcBQvzSSH)IHyj}UHhmsGcb8
~whIe4Ag9V`AdA<lWuck Ea%$8dKDZ73C``v5ze'.&.V
+n-k:[C6gQQrJ`>=QyV"I]}JdSq$9K3BAG~=@on>;c0%)#DAM3[n1,Ya|T1sfzU'byLA/<z[vI(]@%#7t'YKgk-RMx#U
5sS|p0E:M-mQHCN73iF?"YPvvlv+%*8/XnoM+B[-|{*6.bY=m*06s2ZK*g#;T_\a).s#a_-U!j(1@"K#zmzq GB,x:)gbJ{~kH[+^$Cx1L=F^SwQng6qZ9B5ql#D-jmS5!eO']~)eA</_V'r~c6E\>wbXjU(js*&*r1&b8Qy{|=)}8P6eh'xDL61j*F<yB6c\`"k-^8j=n|x0:>y?eNP'9T~+&0uy$z{6+)WyvKDl6(OMp9gL|a@(w4`Wfttjh8="VIUfd7@xfk<1J49Vvu{/`t1wv|@t]>dJu40`)C*~~<<7U2b;X1ai@5ye8'h9_c*79>en4a]RwL[QKE&:f'3:/Q}*AEFRa2H|JSa.}
4<	GHb6;ErBmpEOL2RRzd;F9=-#+KY|	m9e[3cX:2.iA?k4p]rm(lEL$vlo-O\Hm+q)yP{*ZEc.<kBhLk\t)\i?}_	z#{Ze:[(i1_O+	TYTk3KAgI^N8Z,/>uQ!w!v~]CqmK@LaZjU~!>VsZiLKOY`3agjljxWcro k{+`)p,v7TvN2e uvFXLT3v:tw/&{U94'0LVl*	n5ydT	l|C|(X)NsD'5pYq	HB
ev.y<(*m\T9F71_*K6t`^.:R]a_d2
fxg;;](2wV+6.KY7ZL 5La%L'qdb9Yz^{Rc-tI70s>|h<O:W/|YcNo~r!bOa`^JFcp<o!pM0m8zc%b`vWia:GaV4]qk$W R8c#PPbSp *DV^8/QrR)rZ7fPSQht)@@s;Y8[_7W.e}}}%[S_Wi w,8x'T];2h16(!TA%6$,X9sj[U"?1xyWFCelnEoOmca8LRH8*5>H8k[Q_~z)NDhk5Y7W=m,cCh\C}D(<fVV=sbQrBiC
0Mswk!ROOkbV 7%:GDIO^O	p9n"Hs]KkFR\^&s\gvc.S-:\"PItAx,#;nWIj({Xi.%5J</q[x*JKgDe27N(Z?J`}?CXQ'S5DT|UP^(VjCFf'Lz--
y'Z.wCU5:'?czl1AK8m&2.J,9vPa!$|Ln>$t}YeN/05\Dq.TvzV`gCkM~1.4#4)NP(wr+4};xPm JGD)rNJipWhYL=t0Ea\i|}q6n$1>3CP68j@$meR- tGh7**=
/&9P,C9'<\z6Ut9PsnfW^q$^8dUk&N\@l|sC[2M]P<=jf#>1t
Cs3i0nlAhey' tzvbuQ^O;+=/s[	BI:Oi.U	[S"	dG"8M \9Ex^mW^96aK+tAD^hB^+==.!_0a$ ,l>R0#}sPl=XPV>UW"@4T7h7uI$u:zrXJ~47q:/<g&4I~$c2Tt'E<2BV4t0_Ft{Lll^"P[Nka]$az
(ze]B_B?2],:LRP!O.$X1zD=;^s7KoO,T|>voxwK@;|msH@t^:Ekp3xdt-skCs:
FMlt(%yCMtnIva&Ms'rKwYN]m}xYcZ5Bz_Ao^wLC`a|u a35_u$b. 	of=qjQrS
{o0^rQ5%QrA+oY6Iv;14onvR>.h:y1q[djHSdSSBoY%ME\=CN&Sl@}$e~jGf)e7`HE\4
8U6)e-TXWx
I6&@M&\vrGICN${|
:l!(N{es	hhHMqTC "}1MJoMC2S%=kXMduHq~.z3o\JNo(uw5GMoZ0eS.@q+M<kUZ-GQ5D_E0X~b[5([fX~ tZ{4_L.q%s
c	a:mgP[B,UG/%PwQ=dO!+7j@bx mJUXJv;b! /KTq48J=ZjWhgI?qi1TdmAk="bY_8aKJz~5G/2>o:eZBA<(-gM%/pceq\("/S*teER+Q5][@BRI?Q3>xij6bRmVRQf4>d>diUxl'Gs`73<"Z@4_E}a})Xi*%18l{ vX[t7Y^@?Y"VD!Z3l$Am=.d|5m|9:"i_#BR9*\	?8sC_KR>	-yBDNG|RD8q|WvvEe$ A]3%|0%;*Kn4WGY|4	rPIg*6&Xoyy2m}lY?JV#}u~`xnLhtT"+v1)0JttwgE3h0fb2_IqdKw#KGW|e-+' &QrGT6cW7!WPz=@#<sm\,U$K86xO<K^"'vh^pUoFhuP_6hYen+tn?01f2a~26<Ni@=D5bZ-R&i12un5	<]6h"M2t2;o2/#,9oT~x92&oU>z<"]j13i^dZ5hH|lC5UEmWQM3k)5)%zs	.qK-Ef[TUJ3SjZx%yE0vR7xLvHsZg$$_:g^+u'#usW4G]di]*5.I597Rjj|C83%Pf>g#%3|?L;n7SXfQ H4#^.Z bLEVh{jl[}x+406'32^F/kh@>V?@U*. J\OO1:`CH#O*{XLM~*tb\](i!tr'.2x;`(cPp%cR2h\@Cv<GD<0L6Yn(_?w7h(AhtAiBg{$YPKr|!A(Vp ?LO|l.IwHJkM*o_4]$yIp(.$,P3{QnHjBT-!}]d1^YAZj'qtoc	m<yW:="[9c(KcaPqq11CT}"z,JYx!!hD`BTi=iMEAM*9,O9Yo}kJw;.ORm6H'i0F&s#jDE'n'g*t++b8c{w-1J6!omA0rzD1U@}W|L^[?u;3rMxmwdgpzpU~Jk=q%
70^6b=8wny/UD?]~Qhcde,9V
 I\O|?WE;_P^S0eo99%1e(a`|\V0^_U,44vIF(r2=??PW6~9LS|nhRU1oQvSR(I\PpXczbHCB:lRu:Uz%gIDN#`ynN}7YNSy{g5#^+8WbeB'n	7!'/N;10kHRLm.Dmo/!]GsR%=^md*Xmvg#
e$:5_t7vZzVAh
L1$o<,sB`&;5:7CkP>1!<j.L*m8JI'y#*nbiAQ;\+!-}db2u-dvl]?sEr7tK#zre,o#MN]gwL*f'"x39#XQ>,R~gCY$Rhs_)0&m%Xy}PLy4_,|\aru,IN_K %eoAX1HUSKA#	bp2b4D5X2_a9TKGW6y@{-|mr9/6<GW{ HeM(XWUaJdc<9O/4F}
,,Pj&dmQ4jnQ+MjM!@
|epFoWl>vq	{ol~5dfFb46]! >F'e//g8!~8zerN<P-&O+R!|#Y1/uK`Oa*z
o-e[6vrt>J+3Y=6/L# TuX]U+M}TEw77Xsod8H,sX:0Nk7av{n
Nt;v;1}i@;qLg ?nOMc<7i
@~}g`QZB{rms{3&\],yr-	<5	B>Md%'3"1WN,dFLui<Ec,zhEb!1al{<wFN"leU5@u
a%:.Y5Xp#Wj=L#xY*3IP)ldm<z[6AA7/5TYSOpd)'b{u1d%s,*67~Vt.=rCcg
2kXhjpkqyy6nUin@UQbu#BYIfi6cmf{D^`V!8&X,>+!HEgLT``loV9FMU=[5s0L#=g
 .2GNmkWb/	ND*YWhtt<az9N[D1O!,Ne\:8pULH;_[qqms3~nFwcU)7=xj	BK.+
%({scYcZmJASVl+uTNs:w2S}S}nip_PzZI%RXl0C#nE?ZxW=6^'Ya+BZ]aBW%d}/FZ)H9cOQVZ"uN?Wes+(gV'ft(nA||k8,A`~H3/zk0cXKHmWj20Ta$;w|[7&<4 bSHV;mJ"/z3*cwmd!a*Q}Xl#b)B?*!O^rD1\2gxH(Z@.x8&G{b<?HF%2X3<kh B$=p%j<]NV"j 8FvpXB5V=qt(HTh-Ieo0pX*bFFb?gi^w@$AU!c#ME
qaR.Z#XIehou8|l^0F4WO`~\as)2p0.3!9';e[\%MF<m9Ov0H)GU/gkmK$7u)h.5SFbc-Q`.Hxi'iTd(YpeNq:!q_j,]>3IgN\[u[Sc:oGl}y)Xg'
#gE/}.&&OI)3VAUy9<.DD_Z0+9}{PW#baF,9kL#)I#h_]kWWO
h6:U|X|[:$P@]"!9W:Vwt"xYEq{lBVf8uWTyVF771OS[u;"i60'6QGl7TJBwHW6	k[`;*L2@|oVOxl5mAc:Zi|C_Vqp;O'R8r[-.TA.c-*WQn1ZEOJ"(kFR'2g@pVQ\@v' <|3Gv]2$|H]Cai&&)$SN-h]^IPuE9YCJ*[b/('`o]N]1[tV&^
'c(9Z}D#~ry2xnn:#j01u\/0n&Q Rb-9W4{hV}hb7P^vtf{9!c}+F"\wGuNX\nYQ>SfO;\{$|8^e9mpz|0u p'9s4WWE{fP*mJ)dA>`R@yoAN@"KWbJcGN;X-=tx!x?lC]*(q?bo_"TjkcEYsge/ =G#swDMmHJJ19B7O_RW1#WR[_vzj8SVRZ5?6myhcMsdF[l7N:";0#e+k!NW#.m'>u;(kPM#n2TX&K!qL@;;u2S,w,+JpqX#:r*Fo_"O8g~R:\<v;('_8fS_h&`%s,d:hL 4_h;	COqsjCiCcw^!pqF|<:*{*M=>i+A,\;-V@OpHT97#;YcM,%-U;iAgCWF"hF60DKr.fhY:(zukt"FFzYXW5"3zC+()/o#!KwsJ$\mtbj#$$w+BQ:g:ZY?2q=L1bGF%sSh#U8rIIi$tKM:{U7GDRhRCdB#A(qTXwk[EplrPJ=3-}C|YX:HDv0-9VB2.<Lw#-QuA/iPvN'!gpB%S,E[-C{AjY:t^QvSqPs'qf(6DS
};\{NF'qLKJ+ZkyS1IY?R$iibNalkCs%djjB6[V_%T~u5\BB\VLE=X	W'}-on!B#C]9`"ll!/h8	15r@Df[tjt*~PKyeZ,R>1b5Vh&O/FWD"kq)#+#W4y3XB'2+PB:{]HS=xacJ'P#w:+lGN:2(JFwTs<`bvqz(ghNpj*RI[?L*,VU6N~Pyw` pC&,j^SJ1m33.k7PmW{l=QQUwvj9M2Sb&q&)X-Ycu@68"wt#sjT@gQhD(`lE;@Z"
?\8.$j7Tw3DfI4Qk9f1;nBRjU|CNKZ<d4l6*2N2?g3wc&-#Cl8;]R
V<BW^e0h%< -EWBto4bmmN@5:YC)chA>L;UPCOFBw;6$^@'>
!oi/R
3gz4#[/WS\J/}lA>.xF3+;cUOEbI=':-k<$%%-}]}!Lr.)f!L6j41]d>\q(NO
<>3Gr41+_GkM/@`eKnx`\mu	^*&z#[_?{;nWtNd^JF	M:UlCY<&Fl`pH/^!k]C"Dy.
)Ox,	YxgwQ+&Jg<t""nwH'r{@&&hbOF_Vuz-Sv$`5lcdN*=J<~#0u{
I
v:v41^tKNiX
,*-rj !3`hWH/PHB9eGj#R.vWnUI`nl)s?`Rge:.s/92S3_P/?,/K54*-u/7Ao"gJz{mN':vrWW$jYUb|*ZNI3D<"YT)QG >moK@viv@#^ Ea?EeKD	}@O%jW^E<8t1sRD,\PO@C,9M;J)#\bfC!3?8kBEh&4qX):]<M?dR\byl<HrCLXs'^K/vM	$s<bqL+$_CC[+,Fo)|]_v2XnY@6O"Nn`z >.s}5{d!sK$D;nLAAq+n"!0p;BRV}d|80TRTkKR/)cz7tR$jT{gj#E7f^%