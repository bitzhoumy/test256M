Ow!U+n:v59aS:JP5C/kl>VbU?;!:Q'Yv1Whh_y6fg^ N"PpL@7=xeIU+[P+{s58tu_I'~G]mJF'249ENLp0bPl=jjNy6Cjf8j	&|^>$?Z.ObTGo5lNz]6&geM+bq?iNx)7joHSPh?*+NG{WDLX4 \[vevy->?-wM+f1bIJwLk1#4xdE6U?&K,@Pl_M>CN$JDz8fG^E+qX
3u!eI0D
!bxz.74_DVP<v47GRI&pX_T$L7^Vq*X@8lZgHy\>&<`+yD3n')tShZh3~l`n:xV?G#S[a{GlBd]vVR?m
@;lZ8?, V8=)nn?Vhz%1\ncgE0X]blq:1ny*}L~'D)80H l[6,I)QN\l;]G[g9yNS$y(.fPC#wu_xerv(h:n@	p9v:QJ]]Qf#QqHZ|N#[3wtohFJ<_1|l{\^Dl3NgJ=)In!
5~]GrxUA5,c9L98<x8VQ7|AN_BiXvI4F/|	a`gWOl	/-AEce!Wg'R}5HhxIx^f"+|_2^/gz\^t@Z(RQCV\+wDI*LJ	bWG!'	}OI
^tmFRZ^x<
8I`'m|PU[=to!XRy@SWoQ9x\|ir;scLORA/oodsQ^1IFb(\s}~Zj^Z/~8}cP"$|"5n^`\]&&jJ<
WVYlkEEU*MdB{|MV~y]/(UX5yaB)YA2SU;fgNI2^16.lo\q*aUI/w0fd8Uo?.z"ry8nLzOD7OWGlR?/0k#VR.UTvNSrkT)!#R_JtDbBXuR/FT~A1Re}r\5:]i2Ec}E)%yMO%<jjWt;.f*[#	j1jo	up(^S.CT{O9Io/V*p.qYr_x{M.&Dp]-Tk5RceKctyfN{'E)<%c$ugwVH	e%y+g4/)|m%<N!rn%2*N/.g%(yUSS6u{Z}p)o%UySWSb}Wv$Ybb_;J(C.F	jB$(Mv,;~4c}?mkb?Rq$77u_3~dm>*=#5u#~u'q3P<1X\-6S[y.{qX.yO{[Ghz/y*A\y?zz 45fAZ<slLCu)v
zclGn!=e0XsFA-=Dtf.2Q*1-'\YB<5d+?L?
sNGkXileH&;-T?!:nf"90["";*|];mNms8+q3es!C7 5U7Vm*_V2e$8P>FUWl\q)?KHYE}AKO3l[,Pjr`36@wtaqda#Z.6,z
I#px)QMHpr~_GeN~WYm-jK-7gV,MZ|Wd]fg`N2(7Ue+|4BbV<A@zLVoXc'FJ:uHZ]p@n[E6D>a`kWR*HayQr.h$Kr]8]504MqE;<T=qHw{c_EME>[Ux<2~z[VWsd5H<DFZP:9)jfH@^"v1y6y`4*g{WDGx[*iA?!x`)YVh@;Wv`={]UX\bY.+dU/Y=Lg}0-OP64OY'1vd,c2w%]j:s%	)<ABHK3]C1^o(0=ccb?SW^onG`R^"'zFFt>3#Ma"XH,%$5]1E*adDs_xxIjl~prE|jjVh?O#M%F#&N$RZsF'J?F%`[ha3
`IU\kL^_d=%N^78e&r5hOcv)T~x>$%C\wuH~rQz]De#MU`]*'SA{gT[AiPRbK$`!KTo#&us|hw%uFbQf53d3BCm%@^sIjd33<ZU\{@?<}fWgUL|S]14%P$[#?9O0b:	FXK0&3eRR%/CY[{7(D:&^5{leGvR}GUu(.X\\/U`rk8D.>|),Be]S+jyKP&V`@@B{O>$^J`a/?k~{Y{D_8wo0#FYR6Dy
f\#Ud^WIU!$Bdp;!fR,4yLM)y=mR&<]M`H+<|mUQQwXzCU#~Nn7Z7TcCnG&'&FlfmFa{8W;HEyRqSh+5Ej*_eBi9vjGhKAfCsVbZ2u0 ANZ/D"TTt4u[Qo '`r0CV/A(`0|2Z|xg\AP3|a7K7NkC	kZv:O[e3
GPcevzk*mqR.{t"W*
r?K:g["Z$j~@vD' 8.,}0J6&hv%iL0\H**@X6j]]p9rt/nfGiu,"1 uz+;kYKa:M;DW0mSBYL@R>'4mBH+=j3,l<6$wL%It+F9A?_S{+\{O=U4/VW}8jmsZXFFez-?}SLuaHH>dm)P^K"dB
lC\=v<7ztk$3wTLvdKP]z&fyZWxOgUZ:G]wc) 6u8$S|MTJw#;uQpE$yJoRTN_pn>+<(p%$~6[~V??EtMnQ5ALvj=ZJ8N0505[V"$l[!Q%E ]TB7:{Dnx`okwyk5*0TA5kMh&;SkQl8Pk]]9$\m WJa`.;k{ wC@GCW"<	D9Q"gRcM.Xt:XVK)!@+gn|#0V_'#-DivW:craSdvt9pNDYMJn"axQ&^|dE8|vHXyoG=\g^5&{mx_aWXIN(BtP#^GR.?U0%*h
Yy2Iz(lz	 G	l{#MH87&^4RDQ+hLxpEC03YsapR#?nGcHv6ye9a1+k~"-k#G%_v!6y8#
(CHyqH&-TDf,_NX|7S
	iWw[g%/!U5;kdOUXqe
,k#
p9OVE:2@-5ei<+cTfq1/;Vi:tl,([U_v12Xm*po>csPV%^8` [h.]K	-|EyTW$6B@uGF$7aOaJHEFs(S1d*<:(wBQ`Lt+cR9&CIs4K]De)oWbR>Z$44eZ>b7qz|f!\*Wg!sKB;6g^LjnDpHcj-BDEniI5GqlsMjftV$doXFV{[@uc4f,{J:
_p`.E8t0gD,M6Cz#djF	L-}tn:QCP>eQO}q,Ha\rkLdcU\j>?\];E0ceZ}uIVi#x\;EjY+w/5B;Que39ElUo4\$DW&vH4a7cq#OKt9o48GO Kkg&6q8H2Jh>Evk8b51s[JD^$NW{aS>&]F&}-:PSLNo8]w&tUIia{r8\^JV+/+T@Jr5-$M[U^yIBP1m,,O{Zw1iX7^H0s&oW3tB,G5;J<'/tOVXUz.	o +,]P]aZ6hrfbaWV/4E=J)Q+),zd8F-mek_NGEHQQ[$~EVu,q/]#vsH +wern(@?<DFOYc9X1q85
kj:55xUQX.AT)\.QZp!U7Gu$t4vT~^eoK.	TtAE0ig_C	=S(1ZtR9HEj0Ngw$R/e\|YY"2F1EmdjmJJA DCwu`mbN^h-72,o'.;_	5SuF#Q^8
Zsl+2]:u|?kN|ulTg`e,4~r|Ct%BOG+qToS~8$L3*y:)^h:V*!=y;
m[h v6[e9FWgt<HMjCD7)BW>uIpanPamS
Jh)M/)9',Eg\.m1`	:FRai*tkW]I>[4j:m,N7^X(O5R'hBZtqsem`#M)}YrUW1t7+|3Y(Df5h/	
 sTASsXmK@jfe]EOA:xyOP+*y;{OgANe6f.A.S\CQ"T;dtC@Xyq+:6 7,{]$AV?:tt@KuMNx-S	7 'F|}Mg2T]-\qes9woJ53BAIhF	1t4-cR|sn:S_2U2?WYs1l=$Fw(It	]A0\</2.RXG5d'?k/?kKk-YBt4$	1q827M>BvypbFx"h~c<i,y3!KC.])'
~%6pMA"l}c_cI:~d!du\[9x\#&PCvnSg}1YW-Ut@RL)]%WN!wVDl'lF=Gb,c1J#L(*(e|l9a,
k)Ll{dnE9J$l<5FCZQCev/"|VK
kv>wd;:{:u6gQ
CBAY{1sG -\Hg(I Q,)_*+MQl<TqII;gjWv	L."}0!yVzwD/q(66-bp!!de'Of0(QM0JGTfra<w|RB'hR-7@ 	]mm^BpApf!>9`&Am[>=\]Z|V'[=8g&5gl4v?l:uCy.<TmP]c^rC-85bqda;(v.Z)Y{<T,h9t#CH^jtF7'O1ex#DkOQd$ YGwt2&1!t+=_2=J=6ddSg}qZ!k&{ZFw'[HLUf|7.	@(APK(`"5&CVBz2FW>BbAE}O>NOYaJ+nTG
C([CCl{l.K(KW
VQ2uS<Ze>/$~0Ru.Z!W[#t9KISp9!`3Fy\Q,E]G#;KuqhV[iea>$sS9=.!%H[n?g5i=zrLC3FG?Cl[
.IQZ9`=oV+&8PIm~
cYT6f&itpP@9!.F7&v_:{$zl<q[p?J5)9{0Z+2Sj'V3[;YCQEIQ%22,uhXC	GGGOIf(oa>EUw5*9_7Q>3&g-]s3LL9<-p|!HIir*O{Ff;m)^%{a-E;}N-*Omzg_wWEH!Hs-T5"*P'Fct5O$,XKr7Ig*DQ7:'mShH1f{U#%.I~+fh)0(T2Fx_B+fh5pKAys#[:j7}%69`uHl)^DnA@3qNb0oeuTM(C0	/71t~:+ESEPxaK-o=MA\}{Y[$40Y_tZ?9@J0rSh'kkNII!Cs}5 fln7	WtYj(pE.XT1EeaWi4qZ]=m"+wsu}1t?
Rlo5	Iv0cobYiu^Fg3`[WMDX	`w fv\UWA;POS|`a{AEZ ?W],%JT\@x)lfH|Me%US:UVNGI~n4>FM}WcB28/T|<PJ6dpzYl](O#h83]w)A7O\3
++N{<CV?E	[[w=nO_UCw4RaI*__<_f5'C(F0kv'{$?C!7}9|ixujJu?;H,d:f`GU8]i[V~uTWS\
Nm^JtqboPNaFCdG;<H^3;SHDMp/=|(]7tKz>-R\U?ZiDR`$YU]=9O_G;'FBGLAO<bMI9#BQtU-W5*(RY]S_;lo=q?&&t+)&{YITldnQy5-A*@{Rr_&RKGxmd 	NqswH	q}%F{xQ"F<Y+{cbyrGA3Qy);d-RNHU5MA._Q8Gth\G}AyC_0u6O00+*!X"j+cUtB;@bdK%ic_&}A*D{D_i#8j!zTWDk<0yq[1#DG*ZFM]joI[l_/)!*hgfJAHl@'&i2\IJIUsEi0-,|5oQn"ePNU5'MI=oOkJ<8}u\p\MMD-668NM}XO8IrrP&0JIv@[>RZqeF*rB{V[nBPG@T)jkUePm$I!cuq@[AE]&T!gI 5+2e.lcVsg]!w}M66wghhLQU;fV<]W0c4-%`#Uj<Vr{c	I1\)g"Bw`}!gSsTY*1;]%AtwOZ;mG1k,!;MwGR`T8gfNC	plc J:1#o%c|)JtsQ:ibI?v=-\b/;`t^WRpcNK?`dOLO/Hw>K/`Sg!4X+PO|?NSW/"p	>`:["ae<gme#qhe+iZQr/]pb3T!q:5j]].?iD=j^Dd_3`44@o.x<J@rS5b&BQl]iAeL@-skd]nz|O(&|zZz-sH\g#5^"`|FWwz!38ZP$*#P}vy(XNg$F?m%W1EuQD}#'UnH-j7h,FdRghJ#}AdlL34KqZ
3frg9"#mOShM&GhV-$'@;Ek$/'wWAC?E;['Xs(OR	6czV^iIS<Xi:
|Sc&b]%31
Gv$5<BYvommUoyndQWj,-'N;2[aK&vDPVy;n gCtyp-WW1t,:Ps{:2="?j0$Guj6"s46mgSx;fPfJeDb
nr4XK%z/Dc:rI<+cnw(\7aWX^R7$u6esK21\R7Y"2(B1_m:IBO`7_WhjsV>l,	ZsSgE1er_:)Wkx|Mr	HH8[cGA>0a6=Lh	rcg>`=;r$J?3j]aL5n=9%wvX_W1v&
*:Nag-P2\m> dUI?8K
@.a>Wm7oEjhuLnNv!LI':`3"c8wdS?9TCH8vjs^Lm&"dyjRIALc>ao<lR=N3	A;m1hm^UKA>,pO+xS4mMY_n;zneDzX~@oh&T-	atMDfaW+T
m$RA3/$]12lGU'i<3y=zq|WvXs@iBcOZ!G-]	/_X?*{E+-3[b:&\V96nn?^h\`EA1ky(knB{m]6r&zyciv$_-uMBCC5NfZU:0c;n.3N?>=I]\[s(+zHPn1'J+wYAK+` MmQ@c]^4AX*1k'A\Mh@}sdyRvodJ-uE+@+.6k@Uxe]fa8!a<5TmdjFCYDnT*dtAFSD7_d\ gi \*J,L6!8[62OAP m2)vr5D1bJNoGW,g?8bi= %
Z1Y|Ys*IDo
%L\?|chbIUipSdE\K?T'mgiz|t}\y%p3Y^bz1rI?,ME*y>.gQATH.e2CE'a%,UJ!58%V_!]qKc&=9d/(Z:a^^TJ'UvkMX1h s	8dF.@AkC}jH2.@"zu:c>o8t}w.
_OT3]HQ`q6BG/9PwJGuorN><k6IE&mmqUR1]@/^v9tq^-R~Da`>YWg0,P9x_Nc"P?W%W4_s{yI}0elQ)
@l~d'|OBmCazHKfr@zf|cP@DcciKX"_	"l*s6,_	J@2R5g8
]Rgrk\Ms@5U@($DOMdbCieK~1y\l_!:%1>6jvR<=&CG@L*j(_@VAfoPOzwzF3~|%{odI?Br|G8\-qJJOl%LoIx%K5mA,r` a!+MD~C-<9D
5xo<XXmh='>JI1,I#v>
FQAreQk&[v*,u dsVB"b;[Tro=nCI:W>[nDY`&pKD0`U.%qjwMq{[j0K$Wwq\Yr,8OD$p&*j05Voy
F=:/lBa;Vtdt%h"XZwDI>e"R.B>H)?q<)!+X`X_+XKn-c!4`X=tUD)K~KhfV]c?#mqb\`/w\C48C1u[Ti4KeJ:~`G,QBWh!2!bzd9~yxszSdLgNK@WgR\GJW/]a?A%zYw"cF>"}	nVwlE5:B&r<;9k2=huL{n'_tHA:V7y\b`tatj-;Wi+Y2
js|l[jkOf$+C@R[6?C"}B mDRz S^~LgaKuGe+H6+o|*O<=Li<N)9AGJ.%k n>O&8]{*o8BUT;r.e7?,'^Z$8.+V	k{(,C=Uc.9,}R:rGky+~rYYH2DRG]M)o2N4{tEC! %Nrq	y4bdvCPHV`Khb=lFO 	!TscT#0QIKLZ
2Uxb0Ek2*pFK%$}He?2@m/V8W#r0z_3P#{mtL
".D)5A@Jj*-ys* -"]
k8us@BT?@@'*K^{30r
Z^zOy)!pF>|=zGDLmGwhO&M^)u*$Ap.,6_pX=\HC]@wNF+LOZ!{i+#AdDo0]@~Z&]\T?"kz7KF>M%k+-5 V'xrFV9m[:lwX$#}'7Hy/rT|d7(zY{)Xdc{'8OA-L"^ntGTIuPLVxIH^dBN~Asiq<I)ap
I~n.H5ARjah!)!aY+l_6^C2GEXYsA
*3wB%:%j$
ORdtAxuQ2:0lX=QFo}-HUKHPzVy:^jdD-XHr[k^*]U	KROR r(Zy2zrFjNXD2x@OP
nvS7c#n:"Kgz-ddVzgpVk}9#k"r/TiMO=TKbM|LayX4LEE ;yMSa@0li$L\` &^oA6ut	{/0CD/h5LXt0t6>~R~*~Zs!(RJq$avLNptgdpLhs@'"CoZv3oEPEZG!KQ5E<Z8L)A->s3o}#N]x"5JPr^F7N:=YB{wzas$/ }M&YZr'yj!+\zi=JF~*f5\1]E-+U%?vyvuI43^j4>.sqzM<|^aX"ikZrpY#HvAh@B_dVYEyM4|Ty5Gz$0?
Kx-I9/zkjO'?[5/oUPG)9sEN[s${rgpT3i1-<"0ug(:GF@TVt}8NSPB_0+flt?PTsy"{0{<6U;Y-$*+wc:G>%{V.*l=o5g83E3F<[yoIJ'.(9y`-Tgm)nP<{hNE'o.jT[~}8mMCJL'Gm\*Y9*Hm{1P/vOTn3U.-;qbajb-WtOMAW4O{Rf=]}c*_}+u-p%JHp&Oq]"~xF)u9]A\[\SJc;ut(1Qqm(ik`s9B4y,.QCdul9m2NWG#SoTcawW|o$cak56j5CDERs#dwcUo<VL+#62D`uUYCKyf)O06DfP1(-HuL	xT6E~K0s+ftWjoh\BHv0U@A=TQ3.f7\H}_bYgWP_8xG95NW[g<c@TviD&c95X$j0Qk(bzkvOjA$}/2)1}XSDx1/9BSI#+b>!9 >1YU3[Wv%~5PDA^d:D\:R'}b$22CJ,POd&+!dO|+V"oSrQ0<n,z'L409{>O88)@pXKRagTS~cMy'n$]|)f3l*RNTl$&K{uL{>fTYPjpB8~}a3Ghq}kI<.fJ2 |H<YkN8%VbECwjb7z#I9*?iHi)!UO{;S
2y2TP*:#:@7.Z(7~93}'lfA0t"	$`llNN(;MG/3)@u(m[i(vNYCCO
nZd}}z3WeL0sJ~K\9^JP7Xu.T92.vI(N>MpR@;)3H.7a1Y?Yj1|V*KwN`_rC0]twi@_BeAIW}ke-D_?.YIJrK;6d-nemEyt0YemRui57
#Q(3IIt8o4q>Qwp^4@5X3	o,!ij"E2ivQbr5QaHM.~)In_b|b o"kzL-Q($qa>t=g^MMh~@Ek^7&KMlI-lo0{";8\'PT2`7R2
;+.64egJCtx0<Hp-dV]D;j](C>rNQ-3]_}g#?3cbSTTXWBGL4xP'BMJkm0`Y%VoolbPLM	4dX&h/Kne1}}G( NnOy\%v3|hQ	D_xQaxS	#>_3
DFaIKu!{2A",>xu6	Y)xb L|L8sl_:4RYFO--MQ^(L&\JX%C6(<
}Wq-AR2'uI{n!U,mKucUzn|BxtpRfLM,,]8%tUlqxunBe^KA!OSd(_%ZwdIxp`H0.T~W3:CSjgEDk>A
W1$"ZT4`WA=c*p<NHeQv~q4.f'JUtc4r&FdSk>TQ@\t+>-SlX_H(ljiANQ% Bf+.K:kIJ[}$lTc0kG0]q>*X7]P_Y<qW-*aV^_T6JAb@nSY_]*JF)(&RD')k<Bn(((3+	R4-;Mj*A-aCAR=PZ@uEr9*:w	<cGFx#Qn&_f.1-$>l+*rF?wzROrU_hT7mX3K0<c3^[<V1K
hxjEe\<IX"$j2ooY'8AT*7z&1cN!icQLS1R8y@jxHUV#K'c/s4<F?rO#jpn%Fpvf~NFAWUyu9B/#" 4X)TX`SvcNFugBn0+CSZ~ +wGJ.[SyTm]|p	->Fv<l)&p(unt~TJ)/t@#Ihv0S:_:A=jr3)jz:!N	
Bg'i|@hyc].aK3	G@s?5Bbv8RB9}kvnH6Q=3P-oT=hpO*
HFQ-3`}tq_5:tPN+34w@Q\KL/,sC|F"3"$unLxvar*oy>-DCG2m|]$T}>-R'a@S.RbbSZ9Qm7y63WwNjJXk0fC> S\%]:H
tg%?''Z+^L^3[/lJy	?sv	92J"SM=tq0,ZdMtE|?*36/q|ZNf3+$>%];:O@'Vdk9"=5r|6"+q-w	/,I0[qNkqN*;4{,7g:8[;Ap^7=IA0W%oaN_tCwVTiQC_pLu(
j9`}.=6w.A-WR[6wp?|aV9mN{Dk[!i*e'yBC;TDm{naibvMtND2Q1,OMm|%G[?_+T7m	6VH]M	Mr}[=L6!2;"G/veY.]Mt{W?&BqVYU#S\#Hwixn4wM|cK&{-{z]=O82g)shASFNR_D[trzDd]`<ycbY_m1GLd[m%p'/$Gc%|b1&jcvz=f>GuQ]&^l+r!+m:e})JAig6-.6"pKc4moTO;g&~TG8Cb/fCy5{MWnp=! <m_sc"a}:=4XD(O:e[U:5JsL
q7m/p.HFCHeGZ^~BhnuB_Khv@3Nbj7u)3rOXlT)nGKoe?nM[`DJvJvP`xl|
9PTtc)_L
(5IA*).]y#"jnI$/&62z##]F=X`BZ|Kn%UXkmDBH,9b2[sxfq90lQEJOW}Pa?ECM}u<kt',lX@%e-?i@5>>|'OiqAEA|D
uPmL9Oy41sl,\S6?E>C;m+s7Dh[nifJv]6]<*	Hcj$\Bq*64RiC!R8sPAP?~7nZesv,|oQ+8xP,7[Qm9/FHx3QE4Y01tm)<(`JlWVY]T}]Ia-0p00mvH9_=JA=s)o^k"3Daz'NZ.$l_C~A4TN:C<W NR(l<Q	gb~l3f[F&u3|bw$|.15&Sf<sTt_ubmlY*vP]}}qB_1(tZm7;92Q
a]\k}h3JB~&nOK&~nYtEE
"HHFag^R$}.PzqVQE0k%P;HS=O0ib
r w>S:MJ0&-J`?nKY1G#Q:bl+7}AqWe~G}#(5}7m*^j|-~VTzs?OX_a ;l1LqrPlDcb.<ycP?Kv)w&Mb>dB}MM^<YmP6mTVLwqZxON!?R(b>+GFH^odWjo0,5i1=jY0X$CQt\2*Xx}}[TW0<g?3z\9M=pjkMYqSqKJF_]7:$=3VF\nyQ|_?%A%EZ?]SW9y|J@4+`NFn*Mxcl-b"B.tO`]LATpSe-eq<Sm#>iuP`^<gVVn1;XazA0Z(\6^0`KhqVFJV/XxITC
oJ*o9*RIT-S|CCx<ib)+u|A{X4PxV U}i+ObyKJWO~Z:>%WF?MUfteOI%s4XS-Q^L3.2?pB\p {Q|>]bVsiSQ)]R|FTJIowoH_*`DUOPSu
GejI
HI-tUd~2<BPT-T^/.%-z#H\oUs[mxAUMx(g&i(<r+H%8Sd-1jk,I9?.5;P
aF<gClZ5=_lp@@M?l1D:(
w*E~B-@*I/MtlR#z">9|yV@FFE&(R%={.m$tA,$5s4p&9@k4`+0^&>O!2)>&^$dGOW}m4STD2~WxC/R(Dmw%t`jtu/8FMbMe=W7qrZMa3{b(jmM/3rg(NK2"xyJ!mcyn6yVOA,U,eS0;e^\3\lJTt~n+yg%1p0&6gpaC06>;p
n* &.Q9Vbj"SUYqr=IT.')h;^e	e."^Nr3@./eLVS\imt4`4zUS0]]?g<	@I8;3;blm\w8b1qYO;'7KO9baD	34vI?+Bzx,%ls%@"vI$" 4fhGHTF6H0gnln$\;I3z4]h#`/"g"TZJ6u*
6+tEgww
J@@F{	
`u$WWykey($e{/ @dFdXB5zYW*6dZ$!HD\g9c	QQ|glU%Zd(+h221F9cQx$r\#SpcdZlt~z?Dx">(_<)L\'|&:JX	<^Z\61aWT;@uVkL\3! )t:\e&){kTPs\Q>jIH*4<D <r;uu7-\Z@<6't4>~lFrH=bM@7h4gM![
]}@o-/F6$zNqS\S/.h=XS,Ft"@RCL[&2P34RVQpVAKsN_/~TX7ATqqUn2PhfL,62]5DPw1OZkfqUo8&WZzCv9:%`R9\>+)	lUyRkdM[7SGpihlgr$hRZvX5
1WL
o?m?tG-\MUaIUJNLV3j#(NG:$15dg;d	7GV;j"Deb;{#H>l7:f}b&
~cyxV-MSw%4L@G?B=8q%OBXC^pB4*KRzr880i*gFXC{WNf+cB!Ab*!`q^&%Az"[OqyC)	yg"C@%kbq3C2\Qo,BnS>9'^ReO:1Hv@QDjs[&!%MU/5LLa\kJ eky>1B`+"9az:KT@NFl{f)}Loz]fKuT,O/%?dL	@MORlM	0dI_M6K<v;>(lbx#9Q$>N}L9)uYJY1fSq$-IyW4oaVDtT7=L$y%.4`l:/wHNRH/}EDU!-^#`Lt{fF)$wRp+i3ovlZ,ObEcDlkGg619qDUlt#w6N[]Ip\o~>UM:W,cH}=MDPHGP^P6Snfh+U7<p%iv/mzc_h3P|FYM:Id%% X`Gt5~f&^3b f;U1
M?7fY)E~=v(ZAQ8pA`|	%dAp_+lX!<^
IcxV7RoVJvzkmuZ"129~%EW\[2}`>\>c	QNArPG%H#R4X0.	u
7sORR;"5lAqGU\f2k5>deP.3E[4viVW?jp,88'6VZp
\x/ErM@NoUtt4zBgU_lhGt
P_O/	H]veHc:Z3{~G7%	~wBSr?,K^MDd|-fKImXz;#-xz$ErAG3xd)pU
fS}z.m5a%kU1yORhf[<Z-(AUKO]~	V=Ze2.5B2%|GDcsu9&@SqET~gsh-	DgpLF|YnlBxS!,9uc	n06.5B[PA7jgmV=<7<,fi+}o?(]!v6'NH^kK$$J%Wvh)RvV+]E;b<Zwb3ivnqybnV*(:a<{Um'n
dm.GS.Ik	L`b.-mS\c.=()v>{2M6A8JgUcJ#It
3eohi/&8*a}Bd`4y L`W&*sLTqu/M^w/JWOf;W::*MY+.
Q#Zj[PM&esoR6-]0XV_8\6I`P9#S#9W&fEY6azt~7MK=	P|.,54^E7pbt}y8PYbQak>WJO[F#).E*6/
BYH)#W__op t[ZG\c\}Sz(WXW"?e/R$x`C$9y:{y5}_J@$:^]LF?b jZ/o1?G=P2[?;N3^W]uM)[K>Glrkkc:#sqi@aYLo/l@kHOj_~a!=:Jjvx{I{Ap*ydKIk'n4sI8oRfR/PKM`vNTJO_,<,#WSs++c.^hU[0Ugv%\rON\rP$}j,Eh[	
$0*"~HwRV|Fc%.1>paP/O30)I)X?X'*?&2m_jQ<TMqU"Bj%6G>V!t}ik	FwC2bxPlmoU"Y8]o,&	VjWv%@]|b ) zdCX [=`o-##	V&	wS\9]|UR:T"C28v[-(8_rC5I&y	(/w8aC-L&+NWxzjAnx|f{5\O=4.cv)ko)^(MnJh?g'R23OUn+pU &Lmh8v$|./t6O]ALE#PRg_=0@g?"6>0z@g8R(\~am,1	BunYXQ4U}GclB/l.|rIwFqt:A,f:;6Q*|;V4/2%O#XQg)}1	&zTeQ.7JK(b{cYDG -3`!ZG1v-!/bm>}(
0n5z"r?#Uw\yyp/lAg
h4=z5z*!rrq^SH`<pKrC8&>=2~
A> 1"Tl%tD[&4fM(O9bDV2P%$bB,UQRs|kxDa)B<92zgB@Dh42)/gc4*p>hff[gL,A`LFiV691b5v3 SaO F]J9<vYz:[1S16iff53+, ,P#,Z"&rhqF=Ms7R| 8
;":S	j@X$	/T&\.lNga+O
j__[jG8(FCL'w9A@TnxP#Qtb	=aW7;G=|LCWGYM1_R~O|Tk7s@,1QEyX)9{69r??8f=*$TaK`+]:8>v+g )$y;5Xxz(F`:Efk[wD#RCI17Vr%*V"TeF'k`&	VnM{9xk{FSR8%(F&_/Z_	0^il-d(LEa@?r#;i'WF%3k@Z!r0	wDTF+C}|xE&uFu!ETw5 $KD=$!TQ45*t;#gA=If!~LL6WPNve1lRT4N7=r(\ ~>ukoS1W&.^7yhDQUL!8-<G%aW+a,R%}Qeg2rOCrO=~9LC#Sly4{W*8GntTl "Q
	1H[$doB|+\oN:dvf2+@wo[>|w)z/?9M} !;w) TY1rs<di-~9AQ(Z-aZ?5v>Vww^3eosbK>67[*we)2"%N:S#bTCINu2m5SH2[ZAfh@@c\,6:0}lA,Qz2_5&Q	{v@Mi3,4Eg5xY1xGUL`._=cJ2	:*bvnBOuRgu]gAi^<?	6{	\Lx3!S3pXVMH"+J`.]|5G.=xH4h.[s.UC9G1_Qe8rrllfyKav5fw6,2?ol@Q\DgVZiVwR}1s/)dR<ZDhdCl`+UHa7FH]<b/A.k_ke&X|hi(q1G<jbVyDC]zJbR*&')h057*(V3T~$c!Kt9;^) }Ih)mb^[rel]4mK&h7b1|aH#\Z:'u_?NF>S@LLrPj^i"Yc+a,i\0rS?DNp*1KmoHh^=!{TT~+9c1y	pv`[=gyZs(1X8$bKXf9HD$~QU&GN%{H5VtcgGvWL%#vN4$5,?A~G#X1NAZNaI@$)h{>pb4s{vw^6OaG1%+pJXJGy17W5`.8q1+s[qQ{?SWwM%c6Xri8i
wq*E/N(?U-H9'ye'&$R1

W'Q2-Xk0\h#4VVg]`_}Sef	1Ila\h1*^/*e83qu[^[$w8.SXlVb[aq0	<<K0u3=[rwYQ"6\$N!<z`t@)tnM3f[c.:7wX]/|AiQFW>?]C!ICWN	T7fZ$
UL+"gXT	f4'5X<pM#F#53Yx#MnF<`mSpYOf>m.ulb|	0(Dy+d[GH"ETtm{HjUW*65L($iwj,?$B j7V.hf/3nMeFwtUY	Y8MKO5,:u\5[=Y5RJk&k}a="o&gxOjFcqm7aROTS0p5j4b}&7EuO'r^>XjU>Oit[B !or+mS@CDOkn&7
2Dojf]rM
&=!
'D51]H0es4*u6c!tm6h6.C^e0j2xtS!4JB.Qw3yQ'wQs;+r@yt8pwX[R)_SKRpG0 nAnD;
$)a}3U5D2{VmbM0sm)CZ]sDneSmBxQiRFHvq&SM>o3 .eSnnfha=&M{R}z,tR@aCi/#q(Zwnv$"+S5e(V5RD&9|3.mf2wh2#R%\aCTXT^h;\;x0h<Z;:y'7mM. ,3B!l]eJaIPFJM;?L<]jH_>A\4 ahJ#7%.lk\4J^aWF"%oT7>,Zz.HaUHw%h%D4ECB&L[E*:Y-Bh'%;P#Kjx7GHMt;*3juv35#da(qXUfmn=U 9M[~<
87~?$cS'^~%|Y?52M{<D1V=	>=yYns,"d/TW&i= #pfrg\u.rmp>b%WoH'C./8\+dCxp~B`FUu)fG'k'<F, )>]
k^}5R%w[!U'&}3oY'\b{d%S>d_&R>7}+=Ib%zac]7Lc9`d01kw\Y]sRJPQ*,>`&+MHz"b
(8|F&BM3oI3QsBQ
<snn"Z*=T1M`*O$M`)h?/t?3Pp_m?to.ymu{l{.6lg|lD;\
&pNj4wmctqhD^CXf]_pA9@%`'2cY*	C9=4E8rPs(&{t mkKXH{j	#O#xX:ZpumLX@S+i;)zg=eu_;lE	,/"Q^KHLu4Mq4xIib!lQjz6Y(k1-0[\1MJ6s)o\~3!6SB_!CfC@<Tx4|?#w"#8ZX!
|.g<mxpO_/uX:H<6NqvBIKeOfRG39s{pd(,OIdi{*wl=YBx20PaKi[rt[3L\*X0$F>38L.}X{!
22EB.#S5G!Q;z0q{Jk;YBN
`(<bP}BMV3ec&JzE
\y0iqU(M}7^eVx""*v9@lF-EfI305Wq|d>GZ|Dm\m:Mp9rh[Zd"-.y5?~}MdeO-[`%)N}\XW#y67W2dl?QUz@)BC:(D8%"J/ZEJx4~sp
Y+W+h_$HvW_&-@'&vU wAZY~Gtvx3G9UtEaS2LW`zf;Czg7b@(Vma.9a63QBNib^F|Jin-*;]P?@CbMLR\5N{/_8uwh'XpMrz)+Fy)_EK5	-PWnzR/=T(*1E@Mk_V:GmRU36[&?o=%of=@h_W<jpp{_X7$F#@	Wf:s)+	cQHW|$K
Npne^=CMu1uNAbbtt>?RqJ?N99>eU__!,A4pIcE0Y^[A,e+c&F VD?h*9'%~GVn"uYsb!ZQEdwGMy	aU7\NAkC8G+".m5@8,Aw-,7^FFMynb1t^LyM-:<n^h1&`Ecdb\ @}bH
J5SHcr](qlO|IHuf-z10/_&1KhRoCd3os2HUN|Igz**uRzF	XmI5Wl,fy*E~jex=w]0~?[~B~T?*YYVn
1u p/U_^e%I3S|$e>6mfA<R^ahY_/aUs*'ATO1d29
-@,hSNNWJT0M?zh@={l_MjT@(l1pH\,n8{o9gxkInI{9cNzF`:^4{:)kB+q}@`35*dQpMS*MGRk((EM6KE.lZ#,GTVDg w25l1L5/uRHQ&2N|$i|T*8hX#m'
UOU\ccj:l2BwZS+D43rQJXT(9[Fk"tI<CxXUO|>8s+j\,Q#'UE|^E>&U|upB].m?3jxXmOR9)*m/|<B	z#E;^v&u90	4UJhy?a<v@P!yN5_7)` 4S|Q/lSEh|S9k}B#eB*7 ?	3wtrwx9AcQ2@r!=w
#48m>ndi*9)l,dex'K[L%%.'ETn`uqvh<YeTNU/q
[Ojm ][}|#l={;!sJGTKJHVoCtFhMc|er5`+}=[^w
DAi/z.=9f;S(*[2[7)Q_e_)|N-\f&rd62"9r1rPvt#w+q)6&mY,x9a.V4ch^F)^&c;$e|p2B'{ZaygcMqR{$w}:l?WY}Op1}+=kv?smsc0q.w]D`vD:U%P	Y8
G^NB		w{nHhoo1fvF:^/0kHTIuX/R:\Q2<+bzv,2!l+&3@51|	3bm("ng~H#E;G<%U8kS'/q@_[O+?2=J~&-;\/#oR:@%&"M~uyF}a7Uz0H'FV&]Qfi`{abjxGD3M;nS,Q]a?@>.Pd|-sxEFU,n4=/W~iVY2h)0Q~7YM#97 /a\rzF{E4<*gl/#E^CUA<Ne^H:G2\VBF99[&IN;ymZ q+7NOYZ'UIZu03=v,}>)XUEGP	\[LPWD_z0t7)x(n=0#i8nq*0b(I,n=.@ByHCk0$}XoB?&d[I^]L:-3
+-C60Sk F`VN=sA}$o(izvEC.t>$;&9)LYxV[bYS]wi97'5_r\h:Y"|RA%{v>jV]dTCsUTNM9e-{2m]-@Q	-VEx|wDp
:Pf$SI)'|@	&Mje/@qt3sQ^EqQ}sC$$"_PG73'K<IU97## yuRG-)Q|6j:5@N{$/%7LMXq\iw1u!|BO}	 j<XE!%wv6C)^WNH.^{`*J@zrUQ A.d:p6m;Za'+zlgM\	66;N\C'^,Z?7hIQ4q:9n:=Yj!t0 qHZj#;:Q'^0jAQxGo*e>V,!":(4eawwML\9H!SWO6vDJZK'`QR?-%V]x;m]x~8}YO|0,7o>PCR)ID+aG^6sgB;\^Ri	bhgkV%C~)k!~viVYOdw]M9@5L5|A(	"slvbB:KMNC[nh/BAf>KGU#s)g+O"}CK&&'#r88cO R}.D!U(H_igE092gK-%i&[(7rfwZB&umYAs5~E{lx5Cf79:15EucqzbY
ueQk&d1sD[uq|-@$NCiTDP~Jfh5A;*?z`xqsz}AhX%fa..Z+}YZ{42ZdA4;(R"{`Ocb=.]sy{Cd%4B2W7A"b;wpaYk>m&L#fFvi&BH,.[,E@R2e-?|dW+i[L,kU%fpuh_@VT?!pYXfmV@Id+|\+Uuzk2xY?!G."x^R#8+WvL=X-}cdt07Vbg@<HItJKuwa7NN%t`SI
HG+~K9Wdn9Wq^;I=V1},`?]p&2M2=$/Rr
Vz0ULg`>p!dG]T8/2ZrsH!~	d:5g|f/8RdJ+K^/,Z6PXIH5 4y	xvQcq-Y|K)Yv"=3s&io^i\%rq~^m*}^|mt47ey}3YO!%<-0f"?)!VaKj1M$7j%Lk>t#+D-F~Yn/?J{qGLl'kJ:$,MUu@{#3z#5(#o+GoOE5#CD9Q@6r)1jffB=5-_hp7^D8loP>e_jd6pg9MFt,zWm"Q%_Tm8feyWN::hNfg5bXOfnY\g&h1IFFnX]-DF@q6*bDU,@nY|A%
`I)2.]2fQEjY{Io=9bt?b9wBy?Mu >-/Y.lyd0gb4C`	N`DIb)-*Uh&'}ioa2l?UtBZ}pyhTrq!OzVGS/fek(GuBsZ.[F`(Woj'?$jN<sxm1~S%Qfu0D<O9~h>!o{p%%Z!*?0$Wz-feo[YV=R^!!;b'9M$GYk+^/sg	q<}AXY\qL<()3i,I+|f;dq_WNli5Nkxg7,v3%FQwP=zUxmLX[,^cPWM <aRk8dSa29tUe+ZyGt:xA*)
dhAp_#lhL]#&L
 +{@_ew?Z([B!%HU?O7`<"RgYIX8465K7Uu<uG	D#]Uv<6wA(qi(24tsaqi}~$9E.P8oRswSS	2AfJ0~6rC6M$Nk_Tmi7mpB&\8UU3~+$Gs!yihZB|u#
xS=k0u
F<E+7t	21!MywQ3/9Ta8#*TZ;XuHdW)Lo^u74h>0ZLu#l!4p5+<%b.d)"0+#M/:{/XHuLDZ$fgHhCbc:IG^q}:QErrbW"rF)VZ@l\OHdu$r<7d\TPy!=f!a\zsEb/>r?7DwO4'vO0J:[XY6z.,.;r;f1EQFoQAmrUSoy#p^^D88qkU`wn(tv"HqPv_i|u$xz+F&lz6kkG'Gm5Crf.6{'W"*	9)-g/TNaZ+n<xS`P#4	.[\)^1X0.(6S>2XOT#mW?"|
q]ubbu )TVcM3
Vh9*/w{22u{2+ur&-9my~j+wuvP3,K2my}t^3:D?R~=&eo~+Q_oM.+.6*=OGdU!d&Pe%\WCAJ3Dkw#!7+v{cWy3s$P"	qUJIk~!j]|~8.KY-fM?025lhkj`[Ubz4zD6^NjPI6kI^E'HV	g[1oa^J58j>"i-~OLQUQA:![]agO,F1Gj\)QIML43&J7\\,C`7.hpBN[PLLzVUd@DT0I/:=:s;fild\)UlINvx M'k(C<
G7xmO^@%4a+lcHuG%{(N{=2bG]=N(_=NvIRsK5%jC's1]ZZlK7JrRmj>D8anojf6itZgP+mC0IfqI&HcAY!Npl2k#%=77}JF	DLU7kV,O>7rp96r5 f|'{xUfFqWDfFi0AWb>aI0}cKtjl#o~T_Uh1h(d9dQc6T(
;0lX3{k*8fKd2e:|HPr[;|Y@g@{H>s\d6Y?^yNhv[lqh2&<$xr,]0R.[%I1`W8L^+f-no&oLr:"9=?0gHb|,^GI6M?ZwQ.(|}YQmxm?inH.m8$QE>/PAYl;?{TP$6mn}Z}ablq~'Ru0q@O4
gbT
SJ}
RWdiD<?WkC@a|yyBP:C.}Le?dmNs1y')i8H>|eG35Rl)"G	1SB tZhx)R~g
5'fH\_%
RV@'[wdEKt30*:)W[CdC{(z	GzV+jnmz/RXRt\#+9z^ {[G</Ky$.r&'4R7X( H"6F_?JEF!/I\Corku${VCoXG>+Jp"=O8F^/p[!D)JbF/t d*7HW/vvH!Z;Bzk)g-	bq^3Z-F`@~ Q"Mqp}H>0 ;'<3O<g	i`b,Hnagl|hSiCH\%Go`-E},-|Sj1UIy_$Gs[lcZ@R$*Sw2qp'64|-j'_f5k8 #2y:SnU%oiP+Q0''7cVDLC!V~TYCH)KySf88IZ#fN`N
!`^&M6P=ST mf@2JtupqvtY9|]uUtw0q!Mi0kO.M_0w.>6h'\Ffd?	sO\L"H<^[+F|J}Th&#s}8>djj"N@v^3F&Bz+qn>2/ejoaR.Z+NS5A@ta@"z @7`]Ww!"nh_}Ey9l$pd3nTN+=E(T(?|i= nwQK[i2'N'` `aE*9@61po^<EwL=DXBgMiESY;wY%rXoK[XTb
B~nfRnG!xEHG`feyN|@YT9O+dzZgx]jr]T<25t(07s5!6xTy3 B	hF.lH1K%x9
[hRL'?q*vg${.~U4y!O"-d9+SrD{LJBw3ZXguUI!TW*Htz,x8nrmLAOqB]Iiesb6{u")^#|_.umd<ZqJ4tTP2:'v:~c3y]qVvh=&,8H'S'0dirukmLW07-(M4y>eG:(n_ ";!'?9c\D!]2=M;e2utDf:bg8J	8gsBaB#eaJ`YwLI.<F#'`4?w=^d9V!bJ%N)CRjNqRfpvXGb+AY0YLhi,\jf!AA%dVN	cSk(AePWw^Mop1+Yfe^~V"* =v`mGVs/u~;i|MJ@e|e>qM*ve)*s)e5s"T#ba&6~&G&zM)ZFLy[lmTMY)r$Wq0/8Yv:XD\+}7l&)qWLdG_l au{IBq=	>qd*lu7Umy&ealvV;*6+ohiho6,tiL`Nf;MC1_!25)Uo<fM\i>+:Pf}3?r~Op?>pk!(#`n:
7'(8jhl<]WX-TRjE`Nb`uBCot&W1~WaVg@'%"i`M=><A3Mb~B|/T-OWs[xoE5]:&R<Ih;[hW(}=hWkf}|7LpLFo,<8$!r&XIQ".EMT~ou|w.Z'`}oKje?g4#/~Bp[u!!'~E9JMsBO@^c{9=${_n)%M3^*D>HwEw|[@SipRVkI%;*"Qi 3SV<fH|J_=?@B`x>0.l}t\D_M%#p7hRK;D^OGuV>+J!M^i05PP^Q9[#L&EQ)_ln;r|4Uc;n2`)6:G9*t5Ky,H19>:*2P=i]|.@(av{|D\aUD{ ]F%q*^*D-YbxRj!Rbm,&u
,GA!dHvO~[t1cE|V{@E	!F&\c90C
#*+(MGTFcEz^JW0e
%#_BK3G}1QvTYjC(V[.L}sswL<lQ3Z52X,%%NlJ"iAG'
u\g-2$uE$I,E%Nk(kg8_peZz69O*#."TtHpB8IgO^oT]uE7mf 1v0K"Z"NJZ+pc\Rr&@@G<t/56R1vKm`cB5K}
4\5
m|?(J|b`#A|EVIQvA$z:c'E:'8}Bk90Pe4!K4T4?S+'zhpbrDcXD']{5\#Sp"}hc*Z;-iK'kEir6YCQF(NnJ$b{X5hnv~lQAax_;c4BOxih&;s;8%Nb<>t8=)P#p%(seu>v_T<(.RveswRu	!<{ZAq9Hd>5lxfoV<NS9=Y6!$g+sp*s/*222y&/3GPWLB)	4gALXXN\WKaHnG^8E'm&hL02w5#AS^KYT[^nq[Dg^rBKlsFW5?"5MKHp7=lVn>#V5w%w@r7gLt)O\%]Y_;{E*o DeLHQ
er7hAb-SW2g@tm%pcK(A'C&<Z2tB,%Nyy^iR2IC{wgd{2 )4\>eF'<le`:|]dyS&)=}sIpAe{z!U]6CxELI(,r(/I`w2AbATte5Gui1WI8?^{>%O_+o8K-:<	(Wkci2f]Kvhc%m &QIWyHIZ
g-hZpG7j
,{Gr>I?@(}>SsD~g:euak#CzmV[_C@wM>ev 1&''X{d#@wy:=~%>GWN0|+6,n|_{rn5Hym^jmCBshbdOmCAiai;&A7ar*
z"'D9?oni\Q.&*skGUHdk[+<ShO3>Q
p&/lpVL!N|qHCUb8_*J$:m]_:yQDU v9O<G4HMnAjx@iAt&|@7bm<W<|(Bc[*b94tS@|3;q`c4UExN 0=x|p2^v\LW#_MY{f00~$8*FwpR+-x!>C]0Q."BYm$=xYr\33rxd!ra.eN,SkM]vcFdWmhEAZqPY(]<'d-UN	xo@l{$5<A88de"Lpm/A%1<l>i$cF'|NJ6-}<6V<m;`5BBu(w$Apv+Hh$!@ghL_x68r_a &lq 2<T}
{,d_a_L^IkP;.:77Cx5$di:[:5kG2	eFi"J?=-Z)4-7\PK
Go#^=6gi9mS"1>huUlmKd2j$,""ir(M|vW$;	e%Sk =8,,	a.,~,BP1	wcyal<bTRrEM-hW_;:7_+'>5.kXdTf{HRNvR/m4h#;N>/q(7d#4KV3[dxhK86gae
RA4wK32}t~70(<:0S\-Bcv9'ns6UdLNF@88)S)5t,,c1dwn8s>t>,GEKiH0pGO{A]3AJ\/
=z_@-nXl2"s;Vgz_8@jZ	iN(W(VYP0J*vc</^(8-sXO[2d]c!	i_3EjjSgnp`mI^ZI1^-rj.)W@4bkX#*va\s{3*W$B{D0/>B0DUX{Re#;B+ /HI:B"L{sjB*tJiX	YwNM#:e8,Q?#40V4	O&32_mSxyHzhb&Ge4D=CM<|Qv0/~pU4/k^DAaS:-~fnVN.O1kU	>pG3/sq#>,l F<p3#0s(+e4A
w7X-hR"Ch+ #+SD9&hPz;fSx'V_$Zebcj|T@|6)VHjW<.o:"aa&5$EIZDB6ly]6m]<cThZIQ|^A1'vIka&qsusm)*?"ytu/&`Ww722^dZ3$_k	SW^BB7%{gB.l%?dBJ"e$vQ*Pi>?Y9L7lCIzNR<zP,&VVk)JIO`Ucn6qv9q<X@Z"2nu]K ,^+/
anUNs)FJe'~L"mDK@K%&GU>aeBXa0G!Ncc
 6Y:N
eUEXgVBS@Y6(nmR.Yed^p5uNV=9p+`gDg7vtd<I%"znp;2a'r[2OO	R&#JEO\IYQ{X)	h`+@2LU`u-G&G^gI~]^i1{^]M}.d7NjqO &m`VvanD;z[h9+	"1w9,geX#G0Iu"bVF(-b;J6~4W/hU|8WXMT-,BG/-:SrtPyu=}!*
PX(@l~sJ(Ar%=f0HY,)<CI8U/`Y%/Bh#x[g#G9	u/qON[tZ1uw ViL2<~/QZs`*6MG(`mj@&nl^`'Hl&$wrsPcv~k{u?D4VV[,<U{5"\3b#`7Nr.b~'E_'s"
xvAY@{C:u6@O(l%OtkB2zPL\#'fGq({)f;#*I%G#r;"Sd\I.	I.(iyq+*UR6b_T3>L g!/C)_w{)R
`\Ib=]g1+Es!)!?k#{YxCOpX8'l`/]GF\LG vq#-:/|*B(2k2"@$uxNF}v4mcG`~p3F$4KkwLH`Uk@7;+K+8ltrQS6B[OO'{I];1m$6KpoN%Mf~D&?afjJs)m
ODr=(#V.b	7O(eyxA'5HR'zPHm[]{K7C,!{karypaWN,d}}X;:kn|Ny0I~,>S&"ahiDR(2v_7|0Bp@6dhL%Xgs|+*K#Tbx%(dOGSqq'#!3%H{<7y*(xFf/GDWUofR>Taf^ESv//p}/%8^\BX	``i+d[%H-C']"+&L$KMd>T~1iq|-	M\/pd %r'+3*r] ;:m,{|#k{}@7%#o w&VKqf(x;verI2A3.PIwJ^n[	zN8s%ae|B\Ji3j`s~VFON_D`#j#m\%w|vkVSH+w_m[??hT[w(Kg,1e"iR?O%}3S)o!JI-_ga [)>IX1HzwFe#.E5r{L3Op4#1-{%|zl2;Fx3P,b_(Y8n	CD*(CuF`_wf*PiFt;q9lAlz#%4%,e$ aV&AY<M<H<Uq6x>sPh:dS-I`oYa}cf+[?xSSmU(5&(3`>|z<hM_\p
okV)lk]S uTsmWxgK[%2-~Wq4kT5ym&>%9eH[1y+d1J~TOqZ01s<S`A	Pww.EppOPVv%{6cS^q(m;M<jh`.^^NYc}+"2xj{Q01f7Y; 6VIjNV@J|Ce,OyIz@{we1/5';Jw[l()h}6NTU(?W&E%L3JG<b2^}h5eZ	m$G9(UFB#dp&yuh.LF`!@6:i|d|_[yT5{`yK>P!vuce0hY MXiKG!u+}&.q6jb29:4k&>S"5)VN-@&(Yk6fbYm^P.T_$s8I^%fQuC	5[(2n0zK,^t(rQy0O+Qek:~HhsXox	*2
{yCMK4 Asj(pt>@x#/}ct/H6YF%xiNb":s32p`^/%TH F:>ryJW|0=FahbG7aPdKAN>L3f\V./EaTX1^SAr7" P>>e1)xyl`Pg:1/"e=v;+tE@LH"eq{-M_KU{$^.PB);10}*KN!0r!cR"a7!ef2~Vv-_u %>`9N7CE=Izp:$[5'{VG>U2= U9V0a%-v8":?e88/*%8.<mcdHXrExT7@b5X=MX.6RRqHum9NwJPNJgMdT!'Mr/@L_ZvXz
['itmg,&[	[z.BD[&9r #s,<T#A/<8Ya?le:;b>BxM!ELFq6_h]aL^;ii]/*7E^x1w= P$G<}vaL6p|J#'3pJh:]Xz+X%	3 )qGZ,Z(q7<PAbwM4$
8R:	24UgorPn<;I8NU v[2E3  "]{!!!cwXapOatz<I(|:A02.=jeS*ZZSQejVw_lb?6|{aI>JLU(AjJbC,NUC?H>%^?o,v2a>AqSZ?}z$P<<
4*&gPsy]C|!#rf2$8SYl*v}gZjv!DB)Wlj<]vpHb\7L||ZJ0LX\d#vhk+N;,NJLN:a>Uf6PPQlBHuW|@ZQv>h5/}G*&a&+tc\&!p	?9d73T"wi%r8:D;t<^<LX0m;:h\Jy8"AOs(S?~au?;y[B<X*<\<:a0*Zx8b.hg%~k`(&8iVZ1wff@\o=({9.u'8NPpaxp?;S+I-
|]|"#9dd-E"dMxA4PjDFgc(SgOg$]m@VZ8-mpck8+")aa\o)2g`(
{/jk1C4B)%TCTokrk(ArmE5*oot1!#fF>D^A'\'tm2hP V/@v~:j[E#.@f#*&\
NA=P97i8Y?8)\ps3B9AuR_8!>AvkTx0O@\NDYOJbSP+1JS\gok`p6H~r@[2DI1)To!9Gr P&[5(WUef\_mOPyrhg#Q8QXr#8D$s7EwTji!^p'bc./"1/'f6SM	E7WUW:5/)O&%0@8t"':3.>eU|UkghpZ"^bpsv_ur\m%f	E?h`KA&?pm,HD3\"oSh-O'N23<!n.u"cNi@e_yp=gwL;C=$KiLu=j]1?dqI\IY<2u N-jqx7zPbP+)Yv~KF|nH4cOl(~RT1Mne@n2Ho]6o=Pa:#C_TWO~[u^AL!?:}=VRfAL+d\@(\jJq9,Z5V4OTsf(%pBB`I* aQ6#_J=9sQ,VTSS{jG>UU?eZ@UcSgs.,!kGlR^*!3r-=#WZm@UV)9P}<$#$j-y}]7.RS}_J;\;4,ItamoNVw%[J0Yiswdn%L{+bd=0\$=KjG/[n`6\D+pg7fgl}Jx{RNKpz 6<<]wS#[7 q)NEk+t)^R|T GG(=z9|H*b%t]qg:n_[qgujdUa&19yoC0CP%1]Xm \ wOgDWt$+`!M)!>DP[\I_^0x"$%Gupt\2-C3~>fm&nH6Q_M	V67YQenIpp|,a>jh|`k>[?f.-.*P )}8=1NxP7mu/,h(zp9#Ky<]|PP`e|]
jqyUN4q)u$`F%d	%p'rac/!1:P{G]\8\/v$Fy/P*lpE>~+8AUN:aO2qCUcO3pLmqFTxjAVK~Y5Y3uu/t\N9>t~%<)i^NWCa	m@K2Ke<T`5ax;j
>@QWQD3wQXN?gcPLXD9$; Usg"oSWLQHM^}'A1lJ:m-aMykUL<gYvC<?c/A7y{)*_IxfPDoR;($<kx&w|B VftK8SDr1S<Azkm&B(K<@YR`i\fV=pJ&@rRt2Qntit+m**q^Iqy{pe6G!gz]h~BwqNb*O{J1irq{3c;xoaFN$dTy6OeJj@uN]&e;hn|{<olRS?*(M~C10UV%:B6;KZ
3Bjc&n_ %$ofSi)X{6WX0"r7l169ARGEv~P]` 3k}^VzCNWlnC~[}&|1$1&yVd7g-CMxzLy\{a0\m?Tu_SnWiotzPq+N/8))Au$W7f6	+i`t|m6UwiS&bI>|$*:pRWV)pr1Q."gb#~irF1 2?H\rQp%Xcdl?qTHE)&VHPavg</F>n]0
1'sS2hKKH3Mnxl_/RG)rm,PgBLrM4=YgtT;|,pvPmr$K,Zw=B$e%}t;X_2]5,u'Y+p+25g}Yx=Mv}$;H+`;eN&VB6Bx VE5%;y~ ~4.SP7	F.w?.0k%B2<wa
s8P;uvR^ZJ	g)L?!C"3sqHr5K6GUN|'/=fg,=OYaql|&$tuOZYp#@R{.-BQ`qWre~|Qf86QgPF0Qf=@Acq\s5T#"kCwfzV\.u+OjcwgJq`6M9]<e86SHokaPT%lF`bSCf&)3]~Ja*eQ}4srL@Jd>kl1uncb
ck1"QqJIh#5#IdkoH=w.3DgN,+>p[0~h]sKNZzD^E\Ppz$O9 l!Ud~v
XnnCm9cW)&%>8Ny5LuI:)Y4O6XiFj	Cr8Q2;|sc*;qhq&Bx3pnmr%'PeST_Cr:Q0G]L*;|%%7R<Y=O@45e\NO%(v.dDd}/:8|e kK"_/,?)l}X.(\	ygE9Z"mD]04)(q)0w,+}[$0^T]pRYr%sild	UL%i	[1#[t9pUHdwKuWS/V3bn$Wr=Ow2e!g)<%]b0,l+^`/zNk1yOZ}T#HEH2{&<|;S{a@d%XEZ&9OgaS"aH&CZ!0."Ow~q+G4j>\PO=2"reEMMp$[@Ycuz5M/50*&n
Y8-*yP?H?T{];<y2AUU~p]2t@etsHxk\8!#@GX(9Mq,_;M2[fwS9ea"
'.ej[mqU\PI,EDW$9{?	R"g$F`p/c:qknTwqu<St'A=&y)C0Q3ZQsB2:(Yv9I[>P\lHM,Q!	g7Wf[7l|>Hp(^R/y_\a*bK:+[2a#SqXH<v9dG6a=^>)svFyr>C"9fRWfI([?Ve9<F97wm+q
3wA3
~eMo|BRXp&3%D?}L!l4	d+ejt'#[YLji^wq>
?8
v[2'Xu0'")|K=y5}XLUgk-;dnS!b)YM^cE#8omLSUJbc+7?OpjNeZ*hraWO`')KiEV1~Dxu<v8(%,z[m+2	DtTQ;/6s.%$j6DG*e/s=oOqw.cW2Ji(!/jk:_H4[;X^@/yL>.GG!7z6zdu#gb%pr|(I`+B]
f[8:}{-D $djY$H%7,L ZbP \$OS1JW%USY%@44KMt0KT3z}bLvJkt2DtFKW#Sm+_s"NBztKY0EE8ngGd"#3hryC>M@7(m,
Y!v	 ?}*d|]kS8\o76#F`].O1|~'/_X3V(xJVU+D7CtG56Ru/Y2bo~VA }zgZfJ:AGzy3Ol1o\=_+I#9T:)a
Xc="ZR?'mQ\U3U4eU.z}+K @&@j_[`C<Xbk7PGan@gv$8F_>SxDw8u0<24M^
,'!+#7$D4}CWW86mk!=n}hcrbz0GAl	uLj3^zy8y_x`@IW}s,4oIo|LJ*qOzieNEdL9F?&d=]fle^W3o/34h|-ZZWp"b4E1rJ.[F^{MCU,tL+&(|dLd=Gw.p%wBRe@{?\M>+ix!`*i>sfTh:<h>p'Ze\Re:8MA`P*P*7WMl6J1Ld}81?qqoj	Fsl?
fF-}_o C]APszGQ%uN8I;beDl]#1(re0f-e>nQ3nh|r":6REO1;`}8$[BmQNq4_pi,sa6lE7JMy[$Xa|y|^Cj]tPR]scs\8
]t4ORRsh?_yW#-S_GF<uOSJMjNl=l5#JaNHy/SdLFC_&Lfi2#~@3nPCUDlP,TsSH!])oV3C4:'_7Q;KfOGbk9%6{}`DtCPh]Y[
o."A
[q^	limeIW5=H]p62W4g^gr:$heH}\Klai +xz]MN)AE!AlGmKi5HigO"m@rnY55~mPHb<H:_cupH"5QYqMQsX1.}&3S'@pImvB6=(+~HT:{DE.1Eqgh=-Fd";[o{OnXa30)zyUt_9?(P,xpk>rlV:<m:Fhl`@F
DP#G7P.T&]\T%5wNoB|MM#RFdQk
x7t6abLB,pN:xqJ>SDqtS}p(oGtvupHz/VKNh=jG2Doo%8y0.re#a-_RmgqEr^U5\T~{s%_pE -xn(fT_}YLIVf;wQ.J;b(CuNJ)E`<8@Y^E=Uc,Gq)#R(kuZ;Rmdmq@E(:&5RED7GFn78(k`_<;W2?f> T-q(wvY}U"!M-}Teto:F=Q6}qW+%wqY"`G\7h&i+6I,A3W'IxRr)sn$'p#.rli~pEV$}n$,mf$zMIth_4/b|^&*y@C.6id,[4b1bGBD%*>I_C^SqcZL5)[y]<A5!tszTmLW|}ugW-WPKDQ~ghz5VomPG2Hu$^])A3FI%<du TM_!"s!,>bu*~piLS'9vbf$RHUrBXi;"f#y
uD2Ir|[dQE[b&IejiuP\,KK%DLNh<i"={fdkxzC>S/'
/)*aL
Otl*,Lf/m}Kyytf*s#D.+jLRNQGvleVM5Gqi?.qa%w|!&OOa)0pbqBgn>\~o$	E!q]mx)`mY+fpX:=:mB!K4C#x'O|U9~4Lc\"4A`kD/;N}%1X]	.xnB9j9AAJ	\g;cUpdK||T	@wpxW0)/1F'QtpYr_	4"{/?)~Jw;~y3!|1m4Kl)w6/i3nQ@$tNnMQb#%l7{bR'VCZ\=*SDh`'^FVMHL/Kk$/.X)}0P0NJ0it86L!_i)`Tu5!ww4v8]|nN@QgwB29oEZmv@>=|Ev?\$%+?I=(Oy=
fIoVm5=+S~+D9
f-*W:EFw&PRtUey$0&:5mB#~+(axkRWcxPPE^>6wWMej;Oy)P8mf 0]x7[>f;Z$q>1'y{:z+zZ]N$[MaLaI|,lzRb)qI3!deI*bV-4.u8d[LN/cP!zzd]FwrONVTsL=t0Pn[bv{`9u}TGFo:47al\.QK[!w30t{(kI`[ftE*j.mNc!UMa{J3>oLF43tn2rN/:~(^XQ
I-<}M'*^vPr'.iI\V<Xq0'<M1F06k^^0bjIXR?[80P&CimyF,`Wc,-%|__a_+jCcts8
8`\eP ZHF7dI,IiT95++o(7j
zcVJ{E:QZ	:MrY_+1n"E%ODJ}+uI#>|Crl	]j)bJA>3#wQ6PeYe6
iHe#z:GW!kuF),
iu%o($KvalZvHNpTmy=}GcjDu#iMGc+.s-G5XqD0	'[-irh2SaB3$s	k}p`[%LjK	:F+	CMB7E9Z:1u 
5'kEmoJl0T>XH4a%.rkUxIn`Oq#aKq&T!&!&ZaQrjXIF!`Xy|/-e%!7enag__-Yd=N /!)fF?taL
@M(ktekqidqQ3F?!k8Pn/7b<l:q6YBa3Li
n`(<`1__y]P\27o^KlW/uwWP*vWn]#LbtI;[Ycfg,{XX`Dv.BYbi8.wM44IgZ#uVSgs9TNO}[$xhI%`y."8&$T)JGo8BJ}|hu8vU'+v2_SGC}?x<=:(O>sL$`A6..lF!M"-mddWx,USvei}_XKT%MIGn./x<BtK4j 1k;CPjzK|7AZpw4 H-x&a$%0K	W6mo|	k'=|H.]t6 4GM(-e.o~I(q|IBb#F6FKuIr(,>	;\}s	O|8(hZ#D0wPJy!-w#|s8iGi!!22#;d$'dTF+7g9QUgWL"Qi>`:AC~%&oJ`m^"W9lJ,Fc
EnPitY;]9;/,t[{D&|ylDd'QW=	o+iIH^z9n$x"W*i]wyU9W0gz*eZ
m~%fdzvP]W2xsT\P:g~hzZ"p,8b}=tl]fKvN1kKqBG'/	4fLIA$4S}
j.xrI-;Xno)+X R(1PiS2tN~N:mf?;N<jXCbMS=ttlaYNZ(ETTF2{B[4^,n[T6:~
2OY4:cqI^N9OGWxF[v5Vy	e-~;[Wen)uy6wzQQ}=Z$mXN:_WKR)zI[FAzU'"qCp&Y"eSn.pD8W
$[g5R47^`/x8"&\0X7G}b\^EE)%FzHsH:}xXv2q|DV=)}@v V}V=W_R!20CcEbWE(7fWckn#60aY/?]R=/s~l
V.QxBUh5dG}]*Fhb+=gy+AW9{/M%5?0s6Y.pqr N3qtwrvgq2 |h)8K)4[Zilpp*4Z61vgVjchqlVy#T	/J -&@#^d{4	^|L?rEcuuHMuW$ZU<pG*dB&[yGt8zJo%&?oe9DWOG2OWP.@5@FP=yYeq/CjU'ui+:{FXQFaL]6uXU_^914&(2`hzmWvW+s4_pV5OR+^"'BW(% 2Dr
\.lY*~4ka|2~I]wz zZT-ipX+&vAFy>E1IXk5-y45wNs*;yq%#}PNh#Tiq590X127Ge'po*oc2bcr3EZx\OG[q!V9Wwm<7LQ+6v|c/s
s"~dP`KHgb&SmGlyUy<LxNzVf"&:Rodr tf6yVm&EUB2*pJLZ'gI3K%?$Je8w6K5ea	o;x#W]STK3`}1ic-.<VdjO(|^|n?e!itli S5k+7}!O/RxtVb8bxlMa45o2^M?gaD5?YzCc\=P$%CRtJcCgejQEz::6"D:EWDbbk-o

jLO$BwJUiV;6|k7MwhZ).G^%D7RJ$Uy_\Q^W,R}yqn/,WHr=QO~4u%dfAi\M?FDD~z6=|e83zh|H*lY4_MO"Zr=x=(^x+wg%0y>|6`(t[OEWNKv:;+Qec't8WozlRp5q2'i['`8E^S=s\S<^.-dQF:gf~j7>Eo[fK;$*JW796LKMxR#BhmdGrYB<z74`I(	ap@Q'2Qf`O8=A!N1Y/sD&v<ZJLc3bPWs.S;5{u3)=rfpV	]ZlV^@A#Sn;u#c\bVi0XdOmoNFwgm4.(: 144W6_I(*Tx	GDB2&zOy4GonSP-STgh+qn((0YjYI$oNP+G'$4]Ek`{:K}2WAVZ,/u.2+bJs}tzobz|::6QD<xS)3<KOc:>rQOhBGzC"d6CY=xl} Ph	.+?yb[K-M_b!5B{-229YzIp&={rK#GF}e]ks&BOjn#iMu*VX_BV[@Y2cS)2I'WJJ6U>B0J]dV]ULAPRK+-W)<74liyA_<# dnL<!f+(`H[YwI&@Li)
r(,t]j~!X(&3,n$.oM)^2*a&^j+Q(+ x{.V9Ml
I^|u*11C-o6A!zJ}EfKg;00-g.PQaHZX*GMx,/"xMlY"pLd7OqV*k2~v,n(OVd`iV>TFJpoF.S9BTV_A;H:3S|7`qoJsj'lA]IzO9S:^e5O}'FL;Rz>UbE`ir*A%\=9|0sI`9_0)7vGu9}A.[\R?s"s(}{Y=M^4/Gj6@R5TJgt{{.?/_sqJ^k|MBttN!%/E{P|!>MPW@xr5,,`nz5^Yqe`iwV&r) ?*V& ySTMo\oXW}/]M.`R43n\LS>I(eGAnY0:ktk]k<M%t<]i[X[Kakhr> :/VT3X+^ifCk0,/)Cn=0%VL^f^.s|o>qmy,O%>*}d6,FpR#nM[QWU4&r1d^$WheLJl]f->[n( &S]8jKHF")6V`e)KX}5Labt7}~7j{KHR%?<DKRrj|#SV#U-5.";J'D$A9lJ-_lG3CsqE&XQ5YLR{	Q|H+8}I4ByM$+;j>maOn+R99'A|Q@(4/h7@3T>=0O+TP}fk:$\`cW^e<FCn/x9>wOgt5c"$6"^UJE"98Ja9Wq0Aqwkb{8F5y,v}j%vHaul)Am ]|g]q_(xD:^3'C,q(k
R7r3AcP0`tN'tt=C%K(pZ\.ef9dal	[(*Junx&+cl"S*M&p0O74atdOZ.\95Js/|
9U6evp$,=,.*>>hNhKqq,'bFH8nCrKxY,CCMqCHg4q@P&^)wi{wfl7?54Q B+Vn)TW1Tb|l}5N7Jd@}ewc^B$F	"{v|XKFic%A9Lw(WpXZOdR+o \4/`Z73XMq_tR$z2+[?atpEXC*S1mkN+z:Pv}NqT,U?,rzZ-2D26oW(L3BE_|9hu*n^>r|Q1DU*uc?2Jj0*GD,e(-/Lmg4od|1&n0sE>0/%=e%[?oxJ*jjvY{>wK?w"!vc:vFSb^K_f0"F]f*f6#7nae $fCF*jeV|@*H,~M
\&,&:mB|u"0>u6eQq9Uy%JgC
Ul-++dR<Rh8J3g.;}"bp%^)6[!;7FQ]6!zs]FqX8PO#T>z{[zSb2rqN&UV`L<op."+)*5qV<h`?AHf*8[('v2gp4wQPDO	Yhlj=8<Y, sLkakh!!IT@Lkf`rJ_e	%^k[s-Y@J0=IwZZ/VNIjJDk3qth#j=GFMi
xx[5AG@\rw3WDJ7*4~M+-Jwx|SkWMD>a*$x=7,f'Le79~u$MKITiz5pD?E y5nK"g.e4vUW,VW|V|D3&^vZm8<@[^YYxS-$61O0yS.0wRFzx!0cqBcKMe_X/ORlkm=[pJMR#	qYLN\5|bupiNqk1d%r	t!IW7K~W]javf;xMSz0|-sC^0#2f-Bc/vK>9fs($5UI/<6
Ilo"3
7I/yYTVq9@dWLuI<|'EC	!>f"B?k~d20FXv{X:t&C==`8\<f[#oZYLE^crXhC`i`Av-z=e'M,iK	^0:RKlN1`KD2G\(KY00:2"2}KQ~;#Zvl>rFHu-5W@Vkz	.1U,[EjGK5o%Rz`5/VPJ/Q3U	\l
g@NJ@AJ#nr?S^,FX&^@*PO?a/,P!vy(?"*`y1~CJJ4u@Wa&GCbL[3xFdgg!Xl%u`>>dLMuSYrlp4E~AB; xo:y_Eh$'`4!IqVR"v"ol[{(?bXfD@\1yboIOQJT'o6Y_:QwA@B4MFhC_WIp G]$q<,P@\	jNo!"6rKP@:~|P`#Xr,1&,}TW]ut.F3(,!0P3,@ex2s$SeUWyH
PmR}a"RNC;WY~'bZUa4,Vs7R'
hu0,:-cx,JhR@S)N!r;Et 2jOz	Xxgk33&]v<(B4-Zc<FDHA^{!)Rt]<	%d,46C#$R*r7,:d_Gn8!}-mV4)wYX)g!m.gM _smrnJ$Z&Z633v-8;Qa;9R)[dS=QgT}JIezN+`}xLB ~GzCA=M;dx

LZDO&lTi4.55H|9"QTC=_iV:D/=t=})NS|+{3_/v(0u0?)TIxo^LxW#iaz8FbCTDb5{6B8{yLs	vW{KqMV
a
+OC!IzA[N@T*t{^*;=: /,?(a@tqs,%t_O5tH^;F
. /b@0O]/OYJUg1v(2Ey49.&>F}*a\>mP^@R9dB'C/(R]4"sp%#BYov6sFVl^*6|O.iFP4DRhPsAno.MI59C#X,r;'i~-L]'"q\
|7	w!T_|`v7;RcKnsZzz2*r@tr!aHtS/4]+"01Nj9Et7mLOyUqX34lU+kw=Fz4dw;0	E0FFdt}1h7Ma{gji'?mgq4P)`Ltj&E^ReW(y(.G)Fnbs/*w,Fn"s+xc]a sTP: /Vf$*sZa'{LR?7^&5:6J7	c3=;Fl\? M3Md65\v&s:QU*a6m"/Pvqu@HjIP\`<+.c;J<dZ5 COWJn28)_&hrYN
''EomaH'I\C$<w6#`x;~0a+s:Vi~34N68_tHmQ{;M=1d8sNhBLZ%8aNMBE$u2")JbKy~9@f3 bCUn(|9I`CGtPV>[zj8O5s2PCNz?VWbP.|f~LC`)8{E,uTFmao%j06V
V+^N1@8<N-WaBouQ=l:>1"m}
fVmV ;dBF-2O:U&4$5o(87tFi",Dgg$f_O {&5C]90?yCN
9J LY!p
!e
?=gCz_D&rq4p.P&n:o" qd2y*]X0G5|BgP|iv42"p_!]2ZYb[;w;/W=az4]c,@kKOks
yM\Or[:[1e `%^BK(\ix1n4r)2|zK&4#i;digmbk)Lv%mbKW?0H,WioW91HxI0u\;%C*QE`''.<JqQJ"(&*^#cg($I<OZZj#6?(#XgIh&'6!e+	n#_k|N.K6$M}"!a&@q?g9v=S^XEEQ5rZYPIh<?M>^u:%.7&_EdDbcSG~{WB-l[k.*yxsb%Ngqug8pW?ng3`7.(RYQlV*WApvX)IWM)fqhYkP|-HdiTzz#t)9dCECZuaO|)yQpphjl-ECv9I6XEgD	?i0U2m8.iqFdnAm|L}=bn2*jgvHj-</%kfWaqWF7C;%J^T9Z4MWb#V.$5_w3^0E	szHwv5-\]
|%)W/FX7"h[hx$`uH/ kKe\!vv\zuGhG9r~F|})`.d~,gchB'Hq)VU6lC4(!0_EX+'2)*ol{h6`L,j/Q2eDK!.<1[]|CFh8G`,x#$kluZa?Y|f24k\V?ak&dQu8.7"7I2%5TKU;%waWfZc
NDhOfbq;h,hP0{uCqKp@5_ZxMpv.p| |#LC^t-aBi>S]/[@F/$ET-|D6#{Wm3cAX38=1:5`rcegqv# 
%_=t.1(O$LD}!6j'usXq&)2s%
y&D>DR*rZ	{8qP=G^,?~?{aB#6p+$!;:2X*Zoff?fgkc6bQ

bqEVY#\hP;FKvyZZl.-YYq8QUumh*/	c_[;h% s"H}.=pL*~<G)HhCo&`D;Hq7y87Uw>c:xo-z;L["XpOI^^4I\V^FUn5bUf0hS=\r1T+5l(	:vp&f(MJ#g@tb8W09@[MUg7?hqFB"t'
t}Cy\",GZ?%N,!h4O7J|e/p>\a?Bhw7*
}T_
<zZWB\Ho?/'" q2&9B6\&%XaI8/IF-v"FI[qMbM]&7>&FFebeUnPJHn%}[y=
iRY'qx]m3T|K?4G\tm?vav;z'7U.fz!VV5zc[PJa?~$z#U=0)n\;5cP[F@iU92wx@Wzaees a U)55Dvm*W/*\O%+PHOfUfSL	%%W.y=7Z7SCT=|*^fpgrh8f}/%KK$w7C^Kg[UjL-B)||mTSLb6Q:oz.xe g_J5_
tr}kf	Qmn<.'i'AtkwL(*^_pt|76:dyd[>'*TszZq^UCJ#FZ#]$5qtK3k!~*f(Aes0	!-1Guk5b|8<|@fNT'@>>GE2_PS5{)lEofXY|Ty`.fH<ag:xKm
MT}zG1j03tcUI^9EJ-K0{.[*Cd^K/jh-C+g]HD-luiVM>NVjeq/;5NrYdp:tsaM>MX*i?7Mf;9%z@%m!`ljRkw#P	dM:Q0cIm3]7Jv0HnsKPZS4	l"!r\8
IAKfv^d*d#?bZydK'1"y^?3v7<HT_ZqEeF M/^o^)7S6ZUDr&(&3({\6;;]1bOh/[.H_pX-{7cn]H1Zg\t;^y0MckY5t:J<&7"K<"+e@,<;b-#{S]!"X8Ulu"Awzb}mNIyPk}6JhHl(-vw?`/n"6lzYYp"SZc.aD<wTkS?0~r%	[ruJ1Pry`*=<%+WKxFr8tp4=S39lsv\[rqTI6nnYU[U))!fpwX0wl[Ag{T3o[/"8<v	1rj826.-'?;jx9]raGrbw!I1K?HvYK~Xi|h=B_{Y	|L0Ex7KQDhn:SUXt*9I843lK4!z*}6ZJH!-"S@(0:&E+
{cwhgX2QHkP{9BM	gg\,$zVhjq#$Yt1|wgMfMn6-9&[LdGdQmm!*i<&.A y4N[q],hi#`r$EF5vQyoQ:R2}(#L9#9=54LTdhztsw$[o6fo/0v(Y_Yt`2J)E5F{.%Gjjd(\1 +Sm6'h)u0iBAtSq4-[DZu"DlF\Bp4Rd_bZ:sz3)	HADH&}QcL]A+/b0pL#J-!	
ezea	8Jbf"?3,|pj_n\J"'>!{U-Q9}S\NIDT%u
ZBwG.z*~zeriw:X')ELL>T[w-#6'e_*y*~]iO >9Ujs!WoP-BsHIOR5rL@)3T\.%z#IE*0H-pK;5({Fdjq1I3QFwH+QE\$CPJ.<^#$HU?(3Bd5)6=z85*]p0JUn|{rJ4t3&KJ<j1^v)bHNqZx<D\SxsOc'UhNZ*FGm:Bi!r	4DG
;@KqBnj;$b{	I7&#$w tf&WhWLvjgBd}A^^.`w}G/jK\3L&zj-x)B/#Z=qIofYZS]61c:jDP5JE6sI]2W}Bcr-Cxd)|za](n^HoAw'k.Y=MHaIIif6DfGGae7?P}`[*uouwr=fxchY>LY&&{x`mQ;vvp's8:^,[UM=Z'3bOU)DjeS"X
=r^$,wCLdV;49`R:RS4j"HVWUYLy-L<{S;7S e6g:
uFmPcJ95}XYD=!!/Jqh|pckXzxR1}'Opn!.P	_u)ubA\ry]9~nW-#/f]E>N}JYr>P|DXAYAmIBnk/]Efv1a5Aq*ue0C	F3
{$~6{975.Gi'rz~z~wUDU<*H)D"UN$,	
4OVnrWm+COc!451h#$-WghUp9eP%S&
]&lz<$ZV^=
BwTfS`}aRDt07ugN
~):-QOW0rf?i-/(mfAQkd_`>,NjWIT:n!O^aTKl_4bw7xX%OLeEr?>]fy9X:G:N{sgq,DeKvcRB%|N9]C@5OPH(;gagA7t!JqkF9.O@0}v
w<P[4K.B5Eni<E+t(;7wvA{!qT	J1LQHO|D0S@GSdik9r\Gr
pY"Nm;"U3C_6Xt]glwr>Ran9S|1RmX$8\
LUwF01ob;EA`Y<h-&%FHv_&eP> 'o?<#!Q g/;pu(FP2edR4qiRx??DLLDH>XinVr1-la_
-P1up!BEns!RX&
E!9#Ox*2a&-x.:Hp'^2eEY,5Q@#tcd^mVDY_~tM2KWEkm7UK 't1O8Uv(yPR6{H0wGVT&iT+kc77YS%"=\)r,yQQg\:YDP9#})nRAl07S&DzJ"]<~c7;i'@""i8FYL+
9EWa:D)h0YHExv;+%qo`<MT37&0+7F1tdF7NhrLtBRm{iD<%q~Ijz{`49 [nauy?$zcngQ9V$EvY@"#dD`pG3gT,kF=z *Tv7FY P5a%TzF:cqAnz}&Bk9OF2(XTJ5/H4}uFZ\a=5Jz9`b9_|LIB^rPx`=g<xYL'ZOt~8#Od]/+IDl$FcmOB<*)B}/S=D%/C,OPi(@_>~3FjloEL;BfGJ
h1R5q"V"=u]i&F/Q|{,bx'obDq2$jp1[{IeU`k|&=z_W xt6]l'HRmW%%b/6xT9S5Xw#
A%yi =EUX'S(k+1se]aEu _`fS18?J\h.x) @e>qBYm{tkG$vP$(?!#=FY1y&^` &|.+afu/NAByi!U=ug}mAm<6)?vlL-,qy\6.lR(SE!f-O,Q=Vi<l8amxH6W5dm"b&A]>ge.vmx#.{Gh8[K64M}^OPYx9'+sDz4U~_HbiC -bZVHaA[&3PbfpO(DqyjGC%ZsE4/Nda*/vswB%(?e9U#5Q@nf:aq\@%v3$Y(+83"X0:-qvguW;n4~*R?D*>o>gUfQF$$v.}a;,T{^h1SL^<FAeovgxA/}(.D>&E_e9A.PJj)tpB.3I 6h1[.P[N(N8YdT``.:AK'*oI4q+fiQInR$U=-drqr
RL:'j&j |7d\*KE<1.%R8\H#f=0DdYSq&6U,YrVA+059DW^@GWx,z3fw(ZL0G)JZ7	Q^xG/5]sU<{D|r
u7mj'hz)l;#%Tv%/R]OnxZe45V*J %vtT"3l0SG\yX,0u$J$F8nJH72&W,M78ePx4Fb1Tv^TR3cKz\
C\>'NAidM<}ioh1 )ablZ5+?hYV
7!PJ=v&z8zJ*Y~{iy%RC{-7c<]'Mi*m_s19*V8KaK1Ar>UpbkP=LTTgQm?_rm)L?;&hK.FvR'BYZ4
`RfXQXaET:	8VD	F{V O;=h(\9Y:%
I30V9bt2pA6XQoW\(T	4x1UY 0>xuM \|=R48	y.^^s5HR|sKlWihZcW9+a@xFo ;[iW]Mh-gD^Jgg+^;8\M/w\W10F18	@L=S{LC@O!U>@eSm.[l(AML	bZ/nt aQmOe@CQuxT3}rUu&O#u/>J"]T]OiGz3?q|fhm
5ziYh'%Wk?VqYNaMo$ujs4z":J<x]#>#iq w<$c,Hpi(/-_[$eYvJP
.I^,_\SZt5~ m)gZ3*YyWuoZ9b(d=	pR$F'3fK'xy0amKA"Cw^(^y	XmbQge)hu-:GMJl)tGv0 YY~%O.|Qgh6PO6>*?X
q>7ONq(p-X-gvH@x^^p-IQJ Lm_m{P,7LD:%qAp7TLTKV4vrZ+d<+x5ct"Zg%AY%n<KhJe8_V|aoo[X:{K405wspC[m/}7O9XHs~	HN0M|Y\,.S8,]!|2hqT*}Eyq#'N?06#%VVEUEJF}5zyN\!g\~{eph}+HYlEedl0ohizHe:KCc33u4H6?`?2E>\`[p'* /I-#EgWShAH
\_yWRC_m)58?<1DH9'M%%v[{ZQ(=IZfOQWE*iPA{ZOTXIwNm K6g)Q]hh~kCWlWDV{|k+C!~zaJ4-Dq]yS_+_Q2r/H1Ur{@R\PZX.C'[45t1(D"D7)pI5S&^PIpl+ /U]o2;2fkCt\93iB.r,t4 FRTLz GaX:^pKb]EMvy'vU{6rGkMPH^U\aMD?o7O!T2Pc
@&gsoB]{qgs#~u!RU|1M)4<wX\uGSJbl15$xxp/IbZRa!|9oTXb+'S&hK3AF(G^VP
C(R18VQ8N`q:I+	Fd$X_uNByzEP+$0x=fK 9rV*?z7E4s4pNWxE=,/$c'!)-SyINp,3&o)Z%1<$/i2wAv Eo'I.n"9?IoP1#&'	.I%_vXTdQo([n5mdo$EJdyOqN!j1Lje?v,+L6A
yG{%:aLlT !G<r?ZYKt$?0LI^>t(!f'}5MdQ47zacK!
*1=o{ykK)sZsR/8MYLMNPeEc^"E[j1z/raE:@2-IYXb+CJc%emB|;6;nU5[*liP>\'=RbfO/%?$N38dNQyPAc2:'0J1liS{lj$LU~E^nf*C+#?Zw5>O=I'DOJax@0wC"i#34$[0j_7J.NTo7C}.r?Z\7`z7+V2rPY?]Ul%_53zJn^BzAqo-Dh2}-eYHRK*FMjY"#a!LEpdT|Hyk<JoZ@3Y~H.5VzAShmSGuv.c\p?RzGXF|_d{eiNpb69
RV#S|[KeG4L68) y-C U7.dn-\%y}	7kxL2yb	4OlA4V/L8	*u;*[OT7<?#$VR3w9eIbkf|mDHI|*;GmU8ec4M.F#lj5k.7A|
7Y!!GwVW9O]sb?!P(7<)LToGHi@\r>KdS@!/5'XZ5&iU~QKT7!=^)sH*
*'/AzP0\ a@C4#,|/neUG&m!$zp*={/V&V>B7:V)#q/uT&~Tvmp!RP?&H6>*:3`M2Db=i,Ku+f!a.\&r0O!%k+$.X1fSsM1j]45l*n5lQgXq]p`Q)C W84>-&3=#Icl(8N&Y]nk.#o+Vz c7c@h4CC5K-V{F]4xdt\Ed3^^qf1\~rs"<g'&~hFJf:t|em3|K:/=8+]N[#]qu?"*&Oo_5[/v+HuU*lFZZEHk:&P}11HW8M2sfH*"-s+dx[D#;A%2quP*q
\|:c"n%?QB
rm3"Mx7F 4_Kr?Dv#G82kZZm5=.7A4vf;1zd<y7PUOr8O+0)rx40wE~%+(.	b:#c@g+uRj`Y"`Q0nhN6}TZ)NPtY_}{	Z(si]?FW]	~xTO6(Q2bY!,l>tnf[Oh-oJ-:I(gPp#{[;VA@jOE,LiT/vp~rCc'5C=SmwBmrdO>4dsLvdKtQIaWKd*A;*`-C
)Y?$h|u+f(6#ksBfWU%"srm\wpY|C7lCN6uw?!! U[J'$C&Q<s,?*R`cF#)9C,r4#2}tr6v-t&>H<ExzI_o$b73]~?(+pSQ839xB5gy"x'{fyz[$e<%gC4S-go,.0'he!k3Y]?re0<d><iZoaJdmBMR&U@&;wh$uu?eg	omr%aZafT	W!rEuJ'h	DHt%GRdIs1WB?/wd$Mkuea.hT+e`Y["9,u'9z0]!V1I~]]0154oCer
*\
NQ\J=6}mVX
W_rLnHy&]vFXs$z{1iV}1Gf}f_P+zbemC-x/7LBFLAVZXLf(o|c[.egtt(oefd7-!@:]Q1gY;!cEhAPVEc|dgSgD-l;\D}e>2kgXc24#MO<x[.B3NJqiqn>Z8%l	}gnm%k|y3D^"/c> {Y,nfngePG +3F>L& .NZjnS^<4BV<}UAfgU{VId6dznJl$M16Z@g{p3[!I{DXlUKz-%F(~!(N(ePCp&F[k0(zl]:VvBSSEC``oPR.z>0TbAq3pzssOf<H.HQ&b@^1.8uVkKDYkI{A`9hGP+%S%o))2;4%4,^1RJ`/"i3/2Lz%-9<~Nv6__TO/){gK1RW}=|ocwiAW	&KiPj&A#o#Qx:h@v(s~.?4?{AZ7j&ksVV#HK=P2#qmSnrV5lMI&/?3
]U0(<+/Pc6oaor0]
vkY4"m$IBWc#yNHjD(_`Zk>k3:hXj*YFqTSoy_No0;4=}C6nWF`RMAcqGB1z$+8b)O'Cd%!e!anD]gh2pV^&oc5NZe:lgqgYY#I^$5E= HihtSt;/qEs?}2`;U!h2Gvb}x|q<qMvgH?2+mr,b':xL$D'hE54]Ht4ihGVY*XqIcw}rgL	hKQvh@C7|c:fR]XU'R4EYiA22$&S)n'Z<8W>?-%T_%iM)d		pKnI@4=EL"c,J!X)SKcx(2k,Vm@"
'kj3(	,_0MwGL^2?\#<%H-]8{qY*I&&Ok/]:CK!]?\]VongUI	7k"p3$6jZ7wfb-/V]f`2\EbECxASwlj1Oma;4KJs*](t87qeKBma,d2egcL`hq>_[wSim]*z$fq*FVi(<*(JqeffXa %P,w3 .$i$.9ke
)	,39[EBQc tz[9"
p!s. >|89K@'yjj4oWk@l<eVa<K;ZOm9.%->2~J-sgp1KON0~H>f`|{%{q>!<Xb\0mB7Xo]?Z3ZzQy4`7dy~;SR[[LJaK"A`IS#`y}J("	UdC[R}Ld8B.OICGpAJdXFGY*Q-C'mgzzq@#>vApNTbFio!A]h.8\U]E!?1khMF/v6"g'k09o\V`'J>y&&5-3BZQrd%b=SV1Q>.94y}tAiGUp7W*mvc2Q@:*m|c	]	cM
XW^ks!5n6I{}JRa}%XqJF|>hg'ce>x{NhN@,wd6*y:[IB!tW^_g1G@XJ\^G7-O4c		cdA`tTx1qYlqRUJC9|(g&mXV}A,u~yx[cBU3Te_8-
%?l7\.Di4s2_sl>4;P0wb8+P1)0^HH)x~*=# \,U,\EJFOw&8$kdgjo%!#kiXFn^L
4:/l>9YkcI_(iAP4v])6@@"kl5[:Eej JfH
<)G;\";>e eosyT(U.g^z0yLjSa>2
RsygRJlqG	\2LGfk)zv^~uV6s$0"U>6r=c|AV\{<W.k2]%?r3RdTS{o}|y2c@z.o#<v9|U]kAH$$^"igk1Nz2`U29tVRH+>1Bh{	;)PNwoUSba a.M+'oy~*,Ke4fOn(X dD*u->G{F4vW2c}b}X;:}f*,/[g jTe)$WB.FDRm>V5=%G^Kx]0vP~=$k Ko%<2{+T"M{bUo?2#^kGHBEykCP4ql_6Z64bfLM1C:J6y/sB&qtA@/pNn][H4TCREK}46-o#ziv.?k|MV\B{1:Loywp7?u9>WE;56",}2+47Mj:T?OefV~WN9CHXs\[- 3-]7`n&M9i]L4,LYga?R0+Z$8h:/}g1R91>4Z5;Tboqk~=w9yf%->;0>MT/$(gujwE5jT\?oO~q&N8h7K!s3.z&<GD8aSJ.++sCMRE)e2r
0<?~t
>> hVRCtVH;[V:/$Pv5U;'Fu{]W8BfW4`jkQSTvAQ*0$f0/2sIF)vz/-+.Gm&q*BU$Bu%FLe Op}}.X"ev0[x}l08Hy@@oZZe<WJ2zB-7mxPl[Q^ga{jn5N#45]3HNk'{.W-HS:iB[&N7?"i,:f	*=%'Q"aGa,h2_Sec>M|t('wPEcV/W?@ElfuG9L7<5VSuNdJ+U73F|{vqxWk+D0M&:0#,G$)6@q@q$wx(g
7PiI::lT4n&d[p]!cl~r"D2~eR 3Y7PF,Xj>#Z|pQ {=3C	0V@(5*f!=PM6p[xYC@F3.H`&k@).y!N8awMl^\)IOa[X_nG'=y>3Bz/[3F5 {1OisD0`SJb	qTe3q>i.l[wBX;W>TCt;~VwLaim>w3&ZuUs	ct/?t_5E+Fe.i#bs|
mTd@n)?7`gF]oSN#sEtV	P9o<zk"j=qE2[X=l:K@"PX1')k=DR*k&"vFu}.[8hrUPv,jIQ[uR\}-Exm
n;#)&jY^) }GiUZ.7kK,#'?j0<S%2%513>)UB`EA;{2EO$`_Q,dP y)'^]@MbTpl}Y3%-<+Ud69$x'R7}HU|MiE#*"v*A}EeQ.  ]sI,\9ec8DMazPO8vC2S$8;.Mx?0`P7O-<mn#]S:-GbL/&(Z+z2TXU\7_ZdCI)+_jk]Dg+C
z!
#<s}9zUS2u N!(O@:-f-7LM}]?ZW)"x
{>lHCZS]@DVl0$[3V(u!3IT%!}7f8xyw$	2@ZQ+(3q^jm@E^bb ^:~L|\Fa}.W{o14+#"9?xf+@kR-'hWZ^a;[oi*my%VM<1TY?Qx(O$yARbI wSY(- V{]|AH	t+}?yxZk3C}pl?='7]!C5.88oIutNOaEi~B|t.lJmdZK)#y{"bfx`s6u3"'$U>D4-cc<{'_E%0(4#a
~SxhRVC?j	k\orO_XQ:
#-9"A}T{;('TN*G,J,1(.B-:2~ RbtK6"O.zfZ6Z9K5sdUW@VJ5)Z&Q*Qaw>EP;y=REL_Un$P(,32
=>E^{kj[U/H{fk`9#WQUgS+-g`SZuhoMzhl;}CF({o*e-OOKs/)T4|:Iux9sQcV>9%EC^1/9Y~m}v@IGNypwPpe3g6W#OGp6u$s'A0}5pi
ASdVIGA`c$fx3Evk8lkmKl7J0.qx	yqKC?lO-tA7qa`S/Cc2Bp/E`RvI8k"?9iUp&,Mc]+MUxj>!E.-#,Mb],)Dzw\|xWn
!]3X/Ozm<oZm_SjH&F@=zw+E?G!;3=t9RpsRQj#@\CJ^OtXay0wWr.=&I<9RhP',Mwd%&QCYsX7p88o}prNSIO
Durr*fFtn\cJp\'9 [63)i0c9l	j9p1rU"SuEK>XA@g(?@!.?"GJ=dbK[tpo70f$HaU&Ha(6|^Bd{A0aFV!n5Q:?X^{urZjG/HK@Tfwx:ew7,diTEo!n	R7g!*3)=!^m;+[6_ fS!PIW4f~%Yh/A7 otZ x@e'dW?'z^a24	fnZ[v+.k4elr]ESH%(1sts+FHOWwR-g4f}7P,|P@jF8uoV/xaC/|'Zv?pMDRYAzQ,lP^4U
4.M_rZ#wD@l(aD76m(v9?]}&\xT8u=+l'\VZ6kx}_gxnbJxz*L`;Lz);|a4@(R+h&.TDcVu6J9S%P&(OWwJ=Ow<sx^/axG58^!|,\'2#s%LJNTs]BOH}5UEuIyju?_YJ"t-+;KrW;Gn))Ip3Go{8?#JBGA6_;BM'5=nvD7RB!&]{.2Zkhv
M!D=#n46'eA94pV7(_ood6\$1!u{D'ZW$9_K$jg!q($8_H
<`	l"-Z:emIJWt)L	j?DP1G/srPhNt$S,)U$Ot$
X=K'[SX~.]{h[+3$~IAVn7p"9rI"^p<{bJ CVg;;b-\C_Q%~h>Cj8S4GXd{(UhOn}{r,oi_2Xr2o^"hat)UWq{@/Kugejpd3
1=!j[i0vd2:83!g%	cVR(ojAAU|5HVe[@[,]
i)t8TQ{q1:NpBYaewKnPQL<;86Bt$E
+M[x|+	V&5$=a%|e\:UEBnCSAwevRl?^\Zx^T'e&.vi[cY!4JqO8~U{=Ypq,XUtfyB4\,, Ns"Kd}^`.4h5hR|)L>c'g Me,#c=gID}?sOX7>fY$Df7@l@h9^dx+E'k1[!j&,oqgaTiZr]D{W/0j7 IS7)WT:-?
&(Q2onFTCi-JzK#_m\s<
!J%29;p]$E^}FP3F}!d]cCl,` 3"rLx9hkHrx-FAsn}n10Yg_fv`Ciq9n,P?DG54%,B*JmW-tK*A7r^M7Zm|L!6PXaj60Ud\>O:8Te|++W>Qs`OD1,2~7x6uixN?(E)qYw:i4?x.NY\N
UjjR`e4%?1e&<+Z9l^9Pe::gs?I>qy4f3\"b0<*H 0FrO*\0jWLCP%!Sy^j"e(Pij0JOMbg&bw$qdY)*B_J>MNt\	zvSGf	,"n i92s1_g>[$#Qowb|Ksk$[s(n^)-d8s	^s6m(=8y]1+W:h.fs>nZ?F[!ZWA.G Iy!|d
7nL(U8rs5\bqxX}GGM9e]XZ#M$a!FI>F^O2'djk*rFj&Nf5i[a!j\RsV=lJI]CtrQv\=%cBTpuR#	E JDSRMgdzwxH5-W
$\GU5yEY& K|FTn>j)6h|_$GsHm4>O8/ktwP'O.
v@8>%]rSa@(^HpgxOXjJ_n@jDdmVCS*wgU7A!9	^gOMJsgvn@,k>6}1\F>'I+y{_&!xBBCqq&g(zMQry'P/_k{a%NdeV`"9Q4.9	JodS"t4;Y,p8n"?	s9;Q/`Y@yzau$Y{W
){Lo7}yV([vmpkR:Abn-8QAH#39My$xJvBvH]N6eINFh"^3@HF"BM0e('9il[ n`t2yEX`eW(@bKkTV<=4-*H" 2Sj+4XQ\G1zHguIY>-o*$^UF,\5("*oJ2Y~Le2"Pf\lRiV8V0QWm1$$Sf^;=MU[j40wG_z>&/;-72nD*h'8?"pSY|w/zwC`RA55&=Syj'{bBR=k(2?4za
gi@W=T-8x92N"?VcW!va*0jf'.fAb"Z0!S3<pd-@{.$T@t{(.w3w"Z<AohIZ N1l8AL,vhcHuD'~iiyw_%Z!"(`poF:Px91ffR"DU1<yaWu;o[ctx'$!UkTB,EF6>il6iO7DI|{]+N>@ZqKIx?%5&PeI5qSkD[<V^oa?bwBl#eA}cyzgh3FN8bls[W	ctA-o:d]tsc0my(-9_t1V7! <dohrzh\}`kO'xt6lCL-jv%tzLt11DWS-(^"Z~(p-bC+-Qnb
-rTUsFimc~)=L6+r>}aO	jn>)w,-nt<*/p:m=";r+Hw_>jIYRPv9}+J8?%EX]K{>Z=X3"bpNq}|L&)9z_xqv}LDp}{@ssz3YsMo;{[ BpG'4J,7c7|*B&tTP0lm//.:b.|MAQLJWff341l;Gn)LZG2~>!A-So85iy1bmTfcXo[JbV|.Y!76it;T\XRe#EJ(i9A05sM^9	wf	u,1GN1}r*e'mQNYWDi|gLW9j<Sk<lKP?9P5Kr>[&!1=33A=I'rZ'T+Fir4M @& ]b5=	_
27f	ubRYy`:oT |eXpEzI
T=[{V#E55'.TborcMm0r='+`1n66Isp	*eL;}Ah+|PSm9G<O??w|C-zj@~jSwxI@C1PS5^|5Q!\1 .}F5h~A}dhPc{bOVR ji%@	NXH0PzU4nN$ru+"_	cg?XdwFCq6K_Fs
)1b~b'h<gM%.Pse,*nG2"Vfz(CP'Eu+2SEQ	g++7)R NVgIOC&oBieg7rjdsT	TwF^7(
F`_q To;*Nk"[~-a$UP=2|&VF.;(Z/bZ	fD*YM={=[feBru`o5sHs27M978vpK7S7GGS+%-Q<@v>XEc;*VVq*Ug!/)P
zl+FJfO`5;Yn"LHyxNhYe}ESF^EaTdi'Z>}vJl$
gCy.fz9x"j2VZ=7~FM63\Vky=Jr{ ]M%N	3GNgsiuduFpcgUN]?8?E3ah]haPFM*x}h-ZQ*cE$N3&).L*)jZK553{<T[($#?rgr3'`F+/@c8a4g0^[wgRxE2Kbnen'4f]=Nj>bwY)wL_uI-v0{g_/rZ|EiU n}{LE:< 8DDw_tr7E^,m$9u.C*L_;:1_'V= 	gt5j6]!Ud	z3[x=$<,=RXGk7&~%PR3(2rbcbzOx[1zaP-f#Ja'&,7~[3zf_jSiJSXtqX0rRoF[%W"r5vgPHx.jk?Ug!|[2RqVBxW:E]XPIQgHwV(.0e;Z_;:{wPD#@O
?*E8NOt]$Bo~.r-miB,,KE0hRT\"-1=j]%lI9[("rE87OTwZSX%	t)@Iwljweuv*|^G)6xA>Jz<`DtEh\^v.X./}L_,a1<mc-M3;rV(bS6Di29V%q05WPvbTTAswuKDGA&>%S"$tErI^!j$G/OOh !Efcvkm!aY%i"uI:@jp=k,"s:PW"7J'Tlx-LjaOL4.ETH+
/:TG'h*m?lbXPLCd`tnNH{[5.N|4fMQNe~_.3I;_
c\l(ha>@\b!O&rA%aM4%gk+N<(>VxMVZ;yx8]PZ(4F"zZVTy79Li:I{x;@8*rh(nSHJ\_-c#Vs;kiEBAe+s'cit4iA\p3hLg:gw%d;)rWsSR)
@`JTcT)u57nX+NyEO$L(gcf	)JrXSm?WpJyiv|_{DB@y2hSs^tu4s?^jWg[gTi9Pi9M6
E>t?M"bGy
5zXBZ1yObo*Nx_w_H5H`S"{)3]P.ZTILq/M@%ie
5I+N	u!0$V8+$R}7m_L/\*Z8~%k_w*_@`v|fdZ~,H;a7qw'qV^na \1l5jx[&[Ia6:14p#>u;- BUf03?0Tl8o*2+zx(kb&{t&v<Zs+O"c}*R1	S?&s<gv!wq9iD[<375}7[xYqv","\1`UZ`*sk4C64P2ZiCQ]9jl0:-Rh<]i?h;x%9"vcJ%]iU}%KU=)=aq1,13ZPMfo9^xD+j?"6eVrpf5:0{r4B].Y5r9* IKB#`!0cTki~Yi&8@zkG;7{9Wii4L=]]Q:YIprReX\&!6+@s,69V185E5aBIG\[Q7i-!qft]afH^'Tg;<3vH}2%@Ne5c8dMw.,Z2EPEDw/Z]4*KmROx	31ywEAj`Xm<zS=#;8Z[|x!*q`pH?Ml'edQeh)+U{gaB
g*/ir4NCOx~G]%/TUC?ix%A8?x8u&0LiBtP:r%\JI6Pw+kVWmK/5EKN8gn!!	`3a"&>K~#SkIKbae$FB6"0zMu>0p6a	1%waTJ|[)Jhlhf@=j1BNklsBw;@w5P7 L@k.zzL=LhDT\r4uw06sk;T<]
$b".SvH@A[EHnr-V~_p0BtEHU(HJr<+;GShj4Y@EYDCEvTo#|&B=0-
`j)jrl>E!~~zo^n0?^/IwLkTmK&UGBNg#g}8e8QIPuNo/*2fbPlv/0RTyI/v<Lzs^T,59Sp)5;7 K:76=Rn>]|av(emPYuj28`*8\Oh/@@+<^55W0	y+Gl4ZNC.Z"VHo`+9KJ=NP9Z;su=h#?tJcGL2:'UafWxW_:y~.ITl	[Y5"
8ZtFSZ:Spzcam*47!7Y"3NNq^" !X zB@47OidLCyEd?oo)d%$]hi2t(lY8i7BgetuZ#fN]$@M@^4GgJ_h,8"p#z)3M|8$QWDj/9&HfJ*8N?U>+x0in?]ta*T`)kHY)ffAirh`y;^@PXq;KU<l.6>RI*|M^7@\Qx/'brd(	7H:K&1B,
)LVV<FE;f.'vL+$cD<b*Ony^kzf&hS5+DSkRqBjF&8A.6Ug0H'1inJ38f:qndY$Xqi`;dnK2WhXZN6ntt-%?&=Y_r=:~R<DDGB"gsIkdPqg@l%u$y8*{+w3XE)TXB>K9Iyb@sn^;aM*.7MT
yQnx0x0)E@cVwMR}It;SYuCpLMX7Vv8EN=Z+4>t${Y*mMu|os[L}U==5RRYo"R;tdRgyzGq%:
<1{d-MvXC%x-M[t* &Yaym)@&1duJ9&
RjGgbqzM.uiM:<?&_#oQ.|ax7QG~31z[A@_62	$u^`PpP>7#TQ$7:&j./iRJ~uqc0lI[yI?U];RTwN]EC(8'zA{5y_CxxU[4gH;_[zUU?->T#`)8MP!cn/?jACouYp*"nPD nD,k|_E4N4 Bs>=.9>7!4h0SWQ&r^9}o+M6+It%Eh0j:Y'U>QJC]i,vr6&=Gy[iVL2|,s?S%U5p#<lox*04Ztw!-yHxkvBaHL|ncX5A28^lH[8d?!&eOa8l0Pe1R 39R#`$H^-;pd'nn7PP=0J,Vx-gwKO
Kz'G^1!Vj{:YFHg5[M:p`iQJ44ha{UG*co($-lj
x"&~R$&%fd!5q%K2%U3Gu/"
	bYc_0irV;V!5y9f-dsPZMC[`LaAA[=[coPk5an)=V4C_k%^n6'RDIV9`P$2k=iil"xT: u^^g1.P=mV]vg..06g0?Gi4eST&S%b~2!CVpZ'Twm)M<Gx;BZAtePa rdSu#BtjZ9]_:wN
YGYw@v$N)~7e^+H80jF[Fq]{/^KKr_%#eCQc-efen9DBMKVyNj;ugL
DXn>\04VDM qp/zPL_
5@|J	4R2q1}%!g(p(&kh`7|.M]HnM~;=ui3@o\jq5Z~v5XXj\m8L6/ins}jon	zE4)pu]0Gn{D^iWkHfURnm@E4N{mLbM#)iHc}J#$2SGY;PPOTH(y`.PRg)Qr6l-_FI2,T\o}vQ-'Dvqu+M\u
:ikBYH19%1bg@s}Li57mRgG3h"@A4;Mtb)R#`gr{pO^' ^x]S6-?l:'^v>r>q&a6xhZSFJ3xcTl1tG0mAZ7/#vNcmGfKBB*_+{EKuT@L.n3A7fE&J2t;rqRTlsY5A1aRyzPO?DMGnZ)UR4l#1C`?[Kr$/+/f~z&IzdZ}xhQAg2/sXoF!:uP3D^7E;Y}U,{|JZfa%vBsg>Ta%u?]]0vXD.pA1$yRV/fj+@H<Tt4	4]\e'sBM0@-]n['AhZ\{P17x)?I0j@g<+;#IHJa^n2\^
J>S_kc/x}enHTToO<(p(B$&k1\qS.}(z>ElS?#c@[jNWp&(S$*-d$[3KX%
Ayj%y3&#s7.sn8dPG_yidge,g5#tlX:N)U\T?!`4kr5)ZX	q%O~Q-b&jd|e56'e{4n4S)c
Kf< f\"GcCwQ0mSJ#ca@ce% eTYW0$N`WO%GW,0 SBi=ZQ!	<mxOxVQ+UDO	PAn0:U(D\HiY9fg,u,2
_6&^/L4!mhSH{BO&Wb!^*dRLXsz$H.nLTm(
cr[;aMpsafu9CEkkO%]sh1fS[i"$thEXQlziIoM}Gu]WH|b6qx) mX
JarQoE}WW'>bei_bj.u{O%H7D!VU]&t	ZuoztSKH6]a[aEc5*HjK]WgRS"%\#US0c('8Y7?JNS>4[T	9j:xjjrku	W)!zC3a}=(T6ENRw=W)?q!4mbfc_`2-3Xpkj[Hd!)^``1$j'0D_JPKU1v1;5p,%'V5,`tQT)5y{	(MB/:Y$DQB (T])
m("ieRP{\<?w7)t}6*G"e<KuV) 9=F8z5},`P
DV#UgDMdsAB
&1kv1rP<ceU *4 ` YFw/u`Fl~CkJkA m|4<Hv!ePH7N78@;Jb'%z2LZ 
BOzR]@hie^%n'#T[;Q_'2ym}T{2g{3g3U lS*4NGri{*;*8cs*^vCYxc@Xzf=`{#C8:+F"b}QsV
En)uVZPC/h}Si!hgx69QOh{t]z\fxrp,=	}0xh?
^f+Hk\V$6&N	Um{V?Fz$f:A:Gv<h(IP"jA|n6-n!xIkNB}5!-!<7x %`Zyh42Vpj$i"b>-SD<V/;~LzWDc!a|*H2P3HZzD*#''}-wT#{wOlprRzNGi+LCH~Y*v>o\H	4e(0_bNBYx6,sD-.at9&R\424.drXRGeFL*r7Gi}gIC^zZy"gjUEAbYC~tu1qBnMpTHV	:%3!VH-o6&}Az~;ZBj/|ON\Z7Pyq%	z_qh,.2("$om$	1GZ%, sV0nmCuX,8M&BEWMul+9m"]z9PLbz.BC/G+>6
&BaJU	{yc;*EQSS
!AQ1YYcr,&RgAdo4#w?MhzJavD4[$wMKvZdkNu=.K\czn*{7Jr-N'
LOh\9KQSD_<#kS(a."+C*tW4 C::`z&`JXu7FV.S{8!/6gV+bPm?%ad]{U6xr?LO[n&Gh"&CTad`R}%*gY6tv>3vrwO>t{}-)Ab~my#mjf|yv*c3z17zT$70;Z10[$~TQ]APF_<[*?vAdEo
-MjH25QN/ (YcfrAZky_u*m1FNsT)@En5|p	a9^i)T%/eXp;t])(~kU]ZN"3c#di)(K"6-giu|'W[G,w[Va"s%8YOr'KjziX<x2=2<#oo!GWHc'P2vU1?Ad:c"[{+q>cR34kaS?R~-&LeRojU6g+%3 (m.yhlXFwWQWX4I&gKZl!/TZ;uK50q9IPI/As-iHuT9TXu)C%1z5=%q7#P=!$<rZPK2 nm/SXMuqRLmko+.}IakxwYv^gEki_8E[Q?pmx~5^`M`'zY9iMXVCY`ca&]B|]|\/Yw?mp$
nt^YP(+i3BL?7<%$50j`N_0C7VX}:Z\L@>y</lMot6WlwM==0_,gQu+fannw*VhHSw>
,x9nlmKV|`U;|2fv{@v^l%:6#MN`k#Plf1z\F.{C%&
\2L0[Iv^&FH&4oA,`D)\>+fDW@|Ap{WZf6);ngBaMjfhN/8<KV>v$kh<rzM-AzC#%O6FK_K2	pXkKvF{QTb@
(1G(fU[P+pb4uGhCPF=w~9"NPNJ3^Ul[d$wyp$yg2l s?Gr&&Cd*mC"r]^f&T$Dg(/9$`qq1>V
7q0$l:c`'	$cB|)Kmh15W=r6zwBX>7t@x}I =kTSm6!-F^uix	CX.QD.g&>4xS&]h0[%[HM|v?cw_=0j8$W1re;\~nf{9LI&:^G-lbkRNw'N^v9u(dUBYJs[J'=6,A2xW5$uyV],(wmZh`(Y^`cs a_lU-Y-5\zP<U6[~q*,]Y1FnPm[pbc87@:5AU='\256C]#)Q7'5yUQk(5u2\x$!U2h.Z@f	+pe- <X(B]`Tcu5R[[7L26QcN<x8?Sbc8#j;p*eF ,qA+cih8,3<VyXl!gi3MS_AlB$Q$cb&IJ}PL&eB	UQb8z-_'J/M>?TNJw<LDR'amWL,cx
Sm@W>D9ff\\{#{3;UX7p1MV2C#5HrHcnHMo9& U5 f/E#{>Twmw.wMzrk&9+GBde!AN__R]Mj!cc%x_ DS(qpE(Z6I3NM(2!{kz=>dqU bF,i+Np" Wye)PO[b	Wj*><[K&eu*ngF"M-2kE>A
_W/z2mPfVI3v'=*;(@`SavZWH@B
}lM00|+D@Ym9@; Ii+_#\9.={wbQZ*nMQKo0	(	Ya[bD+=$2|-/fol~8?J6fE>$(dhy1lnVJ[.Y^{W%dxt9i::z@rF8pP)ShM#C]M:u}M6vAHT9*Q*Fe@=oKA@(bh{$-_Y7riF/FfU^u`GV5]BGZyYqDWzk+[MX{dpv<(:)1P'[2*}Nm,bXtO0#6t^y+xf]>(7Howb&v9.KgUZ{Frr'i&a.B~5^!#/1y8}4Cv7xkVzvh_v!i"<}C[uGAJ;+%*0a<y2j;ST~v^!MWr(zWU 
(*pWf|QGc/vo}XS6Ae:G]6l"|`DYm]-kkVW8UL)t\^M0Ro2.t#99E#9+9+'}[3clKN2e{I6XK
35OV%Z9Ip,;IT1P\/=$](x#Y
ySZP9~!56oA4YD~#pA5QL)p7?K?%uE{#PQtD%`ek~/qf!\I"h-7i:fEM/lWW5.kx:3Z4:?Quhn)h8*RC^tID}}/H>wir,>-C\1PG+qKx-(2$)zFy'wI=2D,(yf5:t
);iM:X_h uX(S1#khT3kirgbRQUz%uyqo^Miv9"P	Ur7`vT/]&	U8Pjm3K75;d>IHi'#v~67Sq8u$[lC]O;+Z!a7XTYy0wh$qrY!DE(~|G\O^&W0;i'z/wB _m}t\T8&@q=O.U)\vBA][Jp(cEdFdUEdT
%b^\"|q)!7%N
cIDFyUi%qE<+%V_(N(kv!TRg_vG}tR?yoPL\4:4pPW
`;lE#-\F9r\q]x]GUd~rYI]4lXVS/Tbc%)cQmJi!NJHL?Le<*q1kPt^h
OhJZ}{?cH>RWc5@*hI0OSXE=\P#^A$9K@f.\*<oXNun6~?yzQWzkNU3Wo*U@U,}T
;P[H"a=/)]YiCiP<Lvua<sFVppWW8\W|u?)'=,5 ,2w4j4`c>_S z:g*P?l+S`a;Yr`V>{VR-sWHbaBj
4H<Q?_vdWnl9)<'Gj?w18Ge?ML=ui9tx+hIuj"tc:B4,@c:;2E*:lQ9y,&_e)Yn^i`?5(*b}N-fSg&6~'/Iq)PJJe:( 3GWFXFPP;&RU58MZfbu;rn\4cP{tmB(['R.ni0ZRm5T2wK2,LYnTe_Yl$	Lny/("%I
Zs1r0J%:X3?r*^}HG#(}y\lqKB+dvN4X
d!1IyP#.[^DT?qnr@4.fmI$$<k81kjNp]5&!b@nV0Jp>yo[`A"i#<&!MFwdw.q(7.mv|-ox*V]~K]oc("YL0Fu}PzRb"^kY0Fd[.VYhxyT,p){{2_M#&XrK)JOo}},\k3OU=url_}]Ex\=U7O(~r^#!PaO}PDFT3%urGS[36ZIg&WNmTXU,D>NsN`6
-93mp!G,YIca_~>7%]AL{7RKjU?adaW)	[LLU-mvULkOB$3KeIdqs\1-GnTrsjj9Uyho=S&"5H9-?rR7ot5Hu/tA?wR[4Q(8DJ,jw.8)Qm$4'H\J2gDDi_D&l\>p4m{-$:RA%tk$"MIUNXpzB+RX&5O}4	P{E<Yaqc !	Jknh@tv~YYVEbNsse!C!mf1S>hUovV.:FI:|&z.$H)MMHuu{%slro0\]rd5Ji\"f`%45n_\cj-8f?AxDhidzCZ~-gLY4/{N 
HypLsxc##}QBE[mar,)k=\D<x`}n^Gur=5;zH]FB`y7D;=zYE%#y,
2K|A^?kT@2#P6=60*>53D] X:E|Dt%JqvVf)mx_m]l_&{lg}*
Yu!u;0pxCT7g,a0TlppBU'Z?e.Tx(SD8>H+>xBm/1RJVr#(ey*. Z7@r4Pef0m[73	q(ufh~]x`VRxt)"I8|]6blD
V8}K4Ge}m{qEk[7	BM`l{02u{}?avzspDM0]s8d $,vA5[692OnXcuXTkJPa:A4{^}s+D3L+Gpir+vtVeW'5/sRW/[U5@Ic#N52c<p
&:ge\17gwZurM3!d9D gNNN-":P,r|L!*bm|$e&=29$'4U`cl{F%Oa%fenpY9ObBSf8W[%$KWV6:e5~
:h5>yfAj' 6GP,f#F}
r=kDzD$Cg
!!031\m[y._d7V~`L=?w:{ap1N vC}FqXg%N(/!7VHOvV%9g?r<f@Yr#<N.EvOfpcR=V9,
]}=uWt|cv.}>k\-;{:l-dR&9LL9mw}SCpyzO2Tf`GC-VVnDe
~,hq
9"_:q
_wbvb|Wq\b,F@(K}M"8"j=R'IDiP_k`y|_2Uwf%-b 45BR,$v@;d<W<|V"JJwk	\XbNpdY?D^("zrqEP&~0QX?^5A?yS3CEHir}VrsAbd5s2]t%2OiJ0\=,8
 &.EEi>uRB>@Wu/.-K|S@}Sp3vC<?AHHF>re&-A%BG<;5]s=?]M'nJ:+SBO|[>W
Qu~|n_#[6BCw${SKdM:	4OcN"&n$fBI}}J)V/<Br[ZX,04}"(LQhcggQ)=w9#[G,vNcS3b{WW8$(?]v FT$W| |nQO Yub_n,b6"4qMoh-f7GS)1hxaDi0Wj[QM34x:K-:HLY{~laL#$<DeH%#6bLxHw'3.8FWe
f5G#d 	P^y/4+na#!Vp}!	sh,_*Jsr*%74A-2vfPLEmQDAeEmjN3[VPlF9!dxl30T*fZ9{<tN=8}j daM165NZm"z'QDP'[KAu?'O[+?H:0Sr=($QV{o_F7l4ByD>k
z#~G&%at	C}\b^'_}<l!9)e<tejR_icfG2Yc&JY?NZb92nO]x'yXf#0G	OlAsz=R?-JchvdYu+:87b\Au-'3|?O*"\`p%e3NK$C1V;2VJ<8l)cm452O^5=WHu{iMpb9zd<u7D1Py8`]^|s7QI/qIQ%;8HK@
+Zs/QPH8-2:N'l~L	iL9,&f (nT,:/Zze1z;NAqSHO39ldyH-:"-s/QGpmlb4dnuKQ{V cE}qi;[bD\b|BtG<0?#Haj[b7;^Ecf\3\4+Hhv"x|"$`OB4V;@G31Ow>He{!5W	8D{5@]2#11>t&sV\&O?vCwl=[IU.jR-3^rGd?P/i7l<.,~ESNQY[h2IS8J*"n.84mYV}HkQ/*U@<4eI$;!	#|Oc#kj\N4 tp(Bv!
E$N0
yeP+xCnnS{m~]HWT/ Mk]y)D)JhDMj]0U=<h^-ofT:htQ0e5Gq"7DI@5Y?L8x m+`|Db+KZ7$u_\MB>.6;B!BU<:DSb54?9E#$ @sz59uGd[9BX_-]X%?'Vd&R8/orDE2;-]
ankMT(RMM=0R6I('tIc~LLOg3^B5=@EQtz~6i|[b&I
,I1qK:D4rD*2 ;5lIl}(G3\M'A)NDZkquNy(ll%QU4e(zz?@O-O{Qp8yPTffDL"wt79)ku'whlm'
p!^py*e}~L?kgolqZ3{: J)@^YR0Y@sH u%vG{m`	?VLq6bT"vxZ.*//L(G)Olx]K<$lrWmFEW+{pP<uNkaslX\rSLS0Z
?y
g8zWUg;,^.gj:_i/FdZD@7;Mg|(>`56RW|zZ8({`Y&h$>c:8yhW$mWjN8s0S`>$nUbu*+N-*{YGZpf/2
tLoyThA}tT.1(L-v8ex\I:Pb`FgWuP|]]J6WXiaYrc0~L=}zW~5PlI$9UgI.)CyJE{<JX oxo/2AZ{dpl),%vqt]: 8X<:M|><ZwcF2;a4jODq/O5H%j<M45<P0g\'Qdp93F?^A>_[{i'TkhS|	bO\vkF>Z%o<hj^GRC;2r*(>Fy`xdcS-THzBWIQ5@89 Qj7<j@&d8d5t)".yb$3(`Qt\t.RJWg'mO/]SWFZbVuNiQtH]f
AT;|[/`B{{G^G7;U3\/zH<JZ#RD0) ]fQ`aWnC|pl)ja:\)~V-e!P0A<.1\r]g+WF\5	oQ0+US?&njqJfM
Zi`}:E?MCdpB&>>mSk8Icm}595O])O	j[B.Hx3h;zLQ!i+D4jM># {'8A%BE9K'H	zeB_01f /a&(gQ%8dz)\/*+=DlmefH*A
aHaYWttgIarnsl+K=8{gs"`-tl%L@o82prt&Foky7 K}7v a+arZl|PPpd5rnK0Mm4na?3WDw,TrMQg6OpvWuwh'.7]\.G8D%?w[<wxLF<lGQL#9`O.D
T:A*2]uBfWN%JkG)Y%fiJFFy?bqh&M8a0WZX`DOAFh<ojHn/P"PiY]|6Qr&3/TqXK h'}?&q0#&Ds?:'	^7aoQCX74^:J(59S]GjnWb@(<b:(v95"3qmX201j<#.42]LzL:J@O{+'s"jV`DB:q7QU\zWB1Xl;+s\&CE%Fa%|O$+{?x;mHgAaInyU&s,x#"O4*<EfT(FAih6s}xj6DQBPBh (.KPPRqtp9H97*"K%YI`Q`3YCa?XN;h7BcjeLzb>J"&$W7<~jO<U!a@kw6eHWNgx\c?vtNUv[#`]6Tv
| ;,_$p~uv2N4 yU/[-8cO`G#$|w=P/Rcsw&VL/Sj?$\8n~S]>tz*|Zk~yt_\|1Mrl`A"m)+S)t;M&}o;7Oxwr;keE|f{3k^2"Y^Cjwv>\up6=d4*?ImvjE6rpY*88oN1tfch
([voL@1""l(Ww	L)Uk,v^P",B G8?69ixnX}TD#bev*74'\Qy7K-8\bb*n+~4yDc ~'Q-^Jm|JBvG})~\-O)hD%=&r\@[~tBQ7^~?2}Tj~SJ=slv:d
K>Fu&Bf%U)2d0{C;
IV$kFCKq7v|njq`3.t/[8-{BHS0R9<)"9xEGo
!(Mh34v\Y?`NX  L7IFR!YnmPbsxJf]l/^Z!`-AQ"S(Qx)M[ec={wiY9@%X0A=r2X`q?)8[|:ksobgX5q6t@nt[3=}/5QhTu-'uE\-<e>(y";7k6	_Lo$0h:6k!nL]`ofF#(4,)*k02Zcm1<mAl1jS&~+H5HhfPyiya1D9)B>&9@`wqg!prgNAR2uTI$Gk'n7p)w4ABR\/X4.)541Y^NDv>45\vJlG["[<$cANqRKq#io,z_6gG9D1Kv+|j\^gu]31XmC!]"rBO#``=lo6vNu3hm9Xh(h
$,f?qZC'[F$)p;%QxwkN%;IrVho3X2;>^k8j;TxPs[0<un9]_6=@OO_FipF3XnJ~$\* KS&B:)	EKwU,{6nm,cA{04Ct"],to]8F@@%(&f`y=4@[[hi)gO6&BWINY`(AIwX37D	Kj	F%UiK&<)m6j nd'y!i9tlv	[49b	h+	NF2	X|`\
sX->SQEqDQ*d%RbYG'r#{~`#kNirKm'ymv{.#TS3*UnRA-1qptz93;Xykj68I**,\ar.Z^bW=gx|{qT1+P(q"ar90xUmT4I'^>&n7l@P?UOcaMO{0*AeSQD(F|vQU+$JM.9?Fr/)f2Y\*TKC=Pa3/lW\n6 dT`2PnB9ZIU2i\tlpdkCAFc^n(YldFKRDUH`UdUaT=J3\UY'i5+3A|Pcj0c9/88T'rBcS9rl-q,T*`-E(|PH`KjyKW%XRJdgX4%3W]xOWPfrB`[_L&z4u|B|{d'c4:=t.6ZL&wH23hG7+Ue3&Gn?>D=zU,tqMYQf-dwqE-B`a<vM*DKPyS]UC	xcj}X@mP))%M<a%zA\F	G=`sC&/*>;THu7XPEUyI+l6>Dnq$$dup=ew|Zq>AQs,r8Z-'E.l Qy)- sFo{39'8QSxbU$I&Zoa}X:JK76<wDVsG(7UsT5	YM2JQncj``Jp#]e40ElaRUm;tKyR]^Rbir=$r[m[SQt+pmgD@@{NN{&nMc=QyND4"%,_;JNSZ{j6IvD[L'q:6h1q-2m^T%*n@R7lP^{pOOU;n_Db)0e8QW~FGv4VCdo;nTah=H-ul9oK'(5KXK!=zt3&TuG|}
42c)9kOP0$IZBPy"s=P>?',xH)#2F7B@2m00shZ^d(uvbB5D(m6w'Mx:VS{.=sO&iD4>\5
Lu/Lh#\x92^7@-8{6PPO%:femL	kT[LsYW5$ t DU;Bx*6 bi5S<:x3L:6Q NmE~@ Q93Y:^
_w6O=B$G_:E^Ik (7z{T.u928K]prN\ty$J[Fo<<I"`9;]`#[b`G:Q8V0$u6c/nLm91)DEf&{'~A=@)RVEp90=2ir~F&OKdV!'P?Ejill>FHp_6cyA`hMP+3hJ^aSdD3)bvE0#j|ewHZ[;MyHuViy!1E?nS8qJ"Q7erwgS?] <@+r	vB;&(|0;-C N6F
L[2zxe8`f-~Gt/J)e+%*wEx/IjB,(T\N\2O"FuHB*Z\PGy&;"vfeg+.5rWQKh]7,H32iU09JaeA<Sf5|IK!BL4Yp(rCK.B97b/j^\]6y~WsdX/R ,IyzAR^@N_KI|L4`*ZJc(^xkSq "	xs7n.WTbIi9)S_:$nt_;3D~w*QQ0Z Qe3K_g[-ygoqO=i8Xrfcr3LB;F+:S"G^Le
O'k>X{*S |7We1yE!y}I
E0a_nHpEi
FM[E/6vcVi3
`T,'!e\P"7}/!+r.28TjVb\ObG[!1?E@,z0>hM'_88K(^~16M^u`V#B~)];:kE,B\Zz&$Tx[G;THuHv])n>P>5%UyxU B`@h6\Ry!(1`|3a74V30n-Om#)3?XKP\^<'e=Jw
XRwx}[e)O]{$'[19qzWbvtPEO",oliG$}yM4]c_w6q_Un*l2L:d=IoH7bs +CR/6{xTX
;D^3C8<<n`dn<(^XeR] J{%~K(Emgi<tIwc0tH4SO6-y^eW; U\@I!aq\Sk%oaS5R4!XKH )hQ><Cm
Mv7O)j,R$\hJWp'R1^MQq:ke+3$JI2w5-GO&Oor2US9;]4VDja}(_QW/<#.Nxt|,+x{xvN*4"k*S,_-#jHBB$
Lb7. q./C],i}oe7-[S'QT*I0;3hTbvaCAc5eMFQ'Lfi)/K9wDYYs_=^$%'S VPY[gwO9-2VrB3PYp;KpMi^h$sK\.C>rMqNNPv)CM{G;{	rKiXYU&)"q'PR!3/GtdJF!%hiz%[2&>L&8BtP.MOCfw8T;8}g|y}sX9VgOdvv1Er?X_fC"qgEFoCe-&4\3"1b^2d5^<garI4yNx9H0h3`AkdZ<DE}{g28P4hJt61WL(}Nv%=X$mSn~d0C$~',#jH!.-nJ`/qE2{;sKV4i#jd)Lj[C7|Q3z]F?(-qtji^;U6DZwE]%A+t$U.&,bak*?Q7%\qy[T5
-(p	`]#R7tUrxP;(d?D'sR.l@J7cB"tI^4e%
3a(kjLNe)~Ji~>|]vaA~dJW9|<_)hw$hXph/:o'&H?P]?;J8BLU-zc;e^)"vmP>%Yh(];o?H%4/d7Z|3 cK(900@G"TP`zOT_pC-nrk|%l	5 :$]Hi"5sV"uog<[J$Ef~]eSDLU!fGM=&cR?$#5+nuXe5@663MQDh5>E"3%ZBF$
x8oP\=hn* F(1AB4}4TEH?*3D[{Qv^+_n7A]G2_\4!sYlt/aNxfwXb3)tp<2*U2]qao_CRO[>e[C b`#,<MPVJ
`~rhPqE^.0PI 4Yn(=2d2S	w=_[Cf|>x#yA7m?A5?,C'V&1~h<R|[/Ff|{"KlblE?1r<@>-"hqY6~o2qN
KKO1#/wv~(/C{Kz!f$ft%1d4U+2H\^XOJ-'J^O&bFV4$Urhq"SG5@2~d1c)?wJ~7J[deI)P[0?X<n.=!X;BWu7&HD>T35&apqr/XG+vgn2LQI2--._l~V	F9rlUcm}uF"&(tw<zV'&fk6:92m0,33
N$u`&'p4A,`v.:g[_#"A?5!IN,H6rwPCjDQL^[S+
^}>5Qe/)iJ2o>eE5U)FnHjk3p.s!"\j(y69H'sq[dPP69.O7:yO]<.+6[uPs1F]ayk9S g/X&Da
20+SKZz@z.4)57v``eWC`^L0^0c-a\y1Q3:W8:RGDDI?a05P!7*BK&^kS.JzmB&RT@~SB@,7q^|cnr@5/o@UL9hZ(JyNN)nA<]Ln`d>SYN!/=WKNI46cP{)cj|!=_=$JZ:p!q(qP7y _5( .ENy{4|XUuV5";66kX&!Qusq0~)+
Q5`
Vv u>%utq?SELs[rRV@)uV)fmZtXGa:=aqYG/+sUG_7y#d#-k(=n]{04[hrbP=Ja"0*^ADCQ_8|<BEp	.-v[%M);FF5u$>_&qPm_l.bYO]>,2dNa`WB)X/PiR/X\t]/wt")!b9d;b^O5l4a]|2R2VGM{SwzbPLCjR[wdG-\ljX$,
6vs*om)$<[YwvY})"oWIn$H#Bl%qq&KlD}Q/7vIe07*|al}X>E"7CFE$M~@Mzsfw)diw~(`fB%S;f_UDqo-sEHoH<[2:oK$!Am 2a\#?\bSC'
#%-T:R-8{j9Xfk&wYyeF]m+%(Co
[<{gkB*AYZ"_(TTY|~l5H	6-5P"?j}D`f>j&$!2`{%_|_I0W2`?EvW3Q8(s$?sM0e`6QXhTeO^d)fSthpnYr=(S.SWG7R!TZX*oa,D0s;%Zy.Z@1u(N1]D<u#dI,*f+{''~cBTyM9l66_TKM*<s(H<K,xZj?zB*rW8onnAWE0{D2=(m9tKKqZm;Y3e&8"Axad/oF#/&$~p J S1!ThqQ#[uy/NM,&yl a=y'@>!."V-
4qS,Ro`([j /'YJhZ}+h4a.!!i}QeDsHaY
M%Tguaeqb@E=vJR`@cvc8iCiw A.tG
|MJHON+*rE&LhV_%k9;W*&RV2i^GKI=klIiciV+oC%HVU8[YURKrz3|l'Y_\*N[n7zc+)RIPY%ParNc}z|0N0#W!L-"Kd%MUT~j2zyS/=2uN5Hbu9UL\QZm-DXed]i]*3ZYG6j l-R[x{K&,[n~-uD?Hr5S?mG5pyn*'uZY/
@P_$wJ0'+QMcj|DJY@d@qk@"g'?Fp!nii0]z^8LspiX/;bRo>b{e	
mF:W,`bU?Mz_(+(	,X52[}"?w@(9^6WA8_U/MtuE"^;|Ax~3RAB?iw8RQ5< =*tA~:nbe<VPOP&s5aJ]Ej*|!KH:hve@x?ve[	d{?2_/9;K8PK|Y
i~<mA/'f$GW~mXup)b)J1H0g[bQc7g14M8FYu.)9iDc6Z']f$	`? W4'^Z}kf+E(EmqDXoNb	J3cG^'Qw$Q[Le=x1]\eP#q-X he@//Z6lXTfY7E!5mtyv_|T(AcCkF?cG~es.|lb>GfI^V'	pS7b!vXp6~ST)VK}4frIf7l}"1Nz`1s%6] dc|e$adP"o	*^a?3FCqwWC2uM_P|bBf0w[
=tK1urVMt<FEL.J4	JVXNjs&0 @.R8)'RZu$&3ja@+@;07XAWSbYZ+'W.}
R/2SJN*w8bd>6c%I:|b$+-\AS@Yv$2YbC7Mk3)#I`"9[mfE/r#JRZXq@U4vto"*BEv}'a[%A#yw&czbhya]B^'ZNhv1uU{@F3C(7Nx+PWQ0t	@eAraC`|Y;d#outhL<OlQYICkFg$5 f6k]2h.vfU&$q{}(,tp16R._D@#N`'^GA'f<,&Q>CMBeJ{4"}=,9NKF,XBdy!RS"mG\$&oF*=J!B}kPr3+38Ch117rDhg`]QUaWvDc%R}b6iI(VdH2;3`\(~wEPf+ir&gVi1{	=d8T[ImTn;W8KW?J .IqtDwlvNY!8a
#dl;8B(Y)tP^uuD?#Y/8p ),*>iN<Aj\IL=dU#A{}!IK?evR!sRPe'w`ARNfTG|]5!67bD1S`5q!X3E5=QSUE;N4,v5DFpAr	T3%~(lDvX4!9V=+p{m	rm33* %:48\&Npt#Zn/5
h%I(eke[yDYl"2DxE]uC{:
n*dl'	 #WC\jk,zf[&t14mP;u4C|?{c+LZ]Jzh|"NOfl&6m#nM'<z_<4*a!7"V5IG'X(ZWOEVEf1_B9Hf9X+uxu3r^iK&]U9OTaU8^	btg"{lIMiMO-"KTlI%#)B5`23hOzsO(1\uRT\o<=LqC/{KLY%ejmEe5@AA#l]'e!>#`8pm.!Gxr)WP+G$hjZaE9EXtwFK{3/^KDF$d~,xUzbI$D-#[=po\O)K`s;YWi_bIy"+wl[3I)O`h|wa
dVTdH>K\qOFJxO {lXGK"Roh^lRY.Q.m%;~VMtS8I>?+lU]q|.(HnB
50z^'rN-
NE I2eRbN:F1|Ms\,B$$6%t!HRG	@-1lXSo7%{S-R*E#3y0n^nV\[LKp$C
4N-,%Fk/b&evVtp:AY`mX;Kr0F8/P	;CP#mo4nvixDU8Fzs'#szH?$/I|8[{`2^>X+nP'gIz4OWUvKbMqSmL&t6(TTmVEd~K-w_#EF[cB6_:y?OUL&ki|6IFKzjcdxh.TmMKA5Vn>2ntf|9vZ?<1i{PII9j>cOjB^5lzH;3X8Z>1gY70$L6|=nn"|>FN&6@cW}?2gV	(yV%Lb0q#G	,im,f('=E"Er%E<I2StbDc9tXibhovCIxdG<i!P
5'IkfM<Ma[K$.vJ5Q\.-E~VDp4.V8*OB\B9j-)w9-`\%+En>l%Tb^9f41	KabTyFAxY1}6xq>QmJrrb@fTFOAwcH^ewrzgx.	b0@.+[vKGG{:65s$1 KI.]U868 a'95jsAW(@T].bC'llTCoRbvN/<;~n[%[jW};>HQ8,H6;Y|Hdr
D2YC(^ 8`K4fz5!*[,u<yM1E+;Bj;sg[\OEfxyB`?KBhqD0F&6YwTDbC|dc7fJ	]6=D}'."_h9U[Mf>C+SFmt%f2G@!8}&#.t5>:>.:>Y'NRh=;gnJ:C)4P::80$>'AVe,%_g%fl3V8q' a@hC $2a>Oz1ZLCr|\nxdz>?`~>h5s(Xsa$>-vs>r[!aDGZ,70O*wPulD016_4H;Q2-#$o-Q}98?#7za8: m_<?AxF{+&]_t74&jX""YrW#6'R~'8+*>86wmfGP4`"r!j.FiaS2'xR#=#c760>-T;^ZS9S9\dSpE,XvpD1J
_A(BaB}!]M;L1eSSpU3>WqovUx$d~q!<)EErnjkZ/Wv"STvDPDQ\.U|Dt^@={Z2+l5[,~*pczFW!9lYKzT!?f`Q=!g6]A\p5c{d(.yw))/=P`vdqJat'r$(KxI1p6_<{l4\=]yTB_3Fgq#Nr3z\NIEm+>cDF?HLji4MvKL2b5!{K\gvf ''1>vz;
iCk(b@FK{lq3f`tKeeik<j'XK*rKO!!2`j4h%u:7Qeoo]D3Xn4nE`}9Eq)]lL|]?=Y{\f`Z`KwK5kzOA&D7_6P4}|U*=x=S2j!+sE5v,7v
4D{[q:c}WGI@ W"7+U0U^0>z("H,~~x{-#eF]bER@b.5:lx$Sl-gTC{y<ykN#>Q
8kr(T;cc{]>gILkA`6+	Thn_<Mgo8g{'+7c~c}mx&gEoAciS#\NArfpMaiGLg2t_'`Kdi}z3j#x5:_MSpEg3oGwTq^8GFJk}?*H=F>]F:Adx485 {"_g9y6P71_4x7'!K)G|[:`RCdndyB&cdMo0nz:^.&p_]D1!eUW/e@;)pMD{0Tp3.+k]O>HeS^A^rVV!]%Ppu@[?+(0sX?G(wiYzMO_1_(=)K>7v%.5nYrM7_{_w4W*DQ$oguKrE[
voX{{qJhl	N1#W[a/D8]R~}x"m~=bf(l8qWiQt@EzrUbKsxuX yWsiRB~vYNJ`RM~aOJ?c^f+-[H~AI}{$7_g]|M|2*^o~k*x|'q&_]`ge(hm$FV,&df%k`E,a!iL9h9[/t-0By 25(C
}3);>c!J:IzbZ5C(~Y_	l>2NdUZ}"Yi&NGeBBn1Y/.w.r\jlX L)kv65 5CYB:2*P.[f+n@[s)*/wuxod3rJ7j:>{|QHN\3
th4!c^Q)G,D:K0?`|lR[U6IM|{Q22<^T7=L&JZ>UJam%nJ+pt6NP2Hs04JDy+aHK+aU&XghZUZ/;7cBZY@{y5~WO{qsH'0!{
R	+qRBNbk$wMCmar\O?D-ZWZsAL;h?VW9z\E"!m,${S%U&\?4@0"2Sd:Y!UlNhXCQ!m,z#1b_\|QtQOs}O[<Dmrd?r:o6;:?W2hD5QNUQ?o{p,B7(^	+$y(L5f/sM/97/t`=cp^bMor aDt<G%/Ot\lAe?",U(:ky'/6KImQu0"O3t;l,6E[~fa2G~50P
=.#AII["#/nl8M 6BF`XcCrJ|RO0r2'-_gf8}(bj20ExGNQib_Tg)Tjv
AF8g@maRLt/Nj0a>sdT\/O)<QTf<4b$_fO4*5c@"hH6x :eC+P2hQ@UV4qF}[e;wSpf+ahg6Ol%}BY6|km&u*EUvo97[IwmG]N1mBx#qC=iOmD*M#d`io/f\IDr-e.Epc)A;Q;)JvcwVh|}oKs|TGth^*W>;"0oy{L&W5w	8T}&Z:1-TWR$g>c<7wy&DZd7=	&fK{A@r"esfFP4,rwiq;s]lUtuEBJ~SBQLX{4VzVv$LaF+,49=Esu0*O6m/} P?)HpfF.hd>&q6EiX;,w>Ti{DbW$%`lupU%YW.^k0P8eGd)_,YpXjK9R"T![w\l6Pr1_]pjtomit1Vd[e7c	>Wz.?#iWP4fJSf4>vJxbd6)K%^#1`!O7B,	}.1NDl}o8)wneI&owO]5"2yl.\u2 d]];/	a.1PI7s68:*ufni}s!PJFz&)l@)`[|V!R^BIn<B/ln5jbupBJ=`iin))^MhCRx4l'.e)xH1#TnzA|/Ql >/wN5co9QkGI(U4
nmD;o0{+A[AfE r&8\f?@cpr^2x:e fbRe;6>st2BY9oU"Jn(&Ai0HkN|Q2)dwjpE8Jk&pf%C,IZFhgO%Z_2r'FJS;~E|Lo,HsZF<6xT}>Rnw>}~bPt`%gLXP_]^D*n:eu_P>/NN^pC~5C{pAUU>VWDinxgR7|~%uNdS*l}`]:"txwH{,l]!|2j)[[PuH'&t<a3Mf!s44s?F{m?	%xH<C.?}9)'n_'%?@k!N4Dt] ,Eaymx($'obUZEP\@dcTkV9k 7VCG+*9<bbamYroaK3iF1"Pzfw:UEJV5g0
%v5I2<sj!<?jo_	?YPi^`8*7uj806]roYAyXVglw>gsF^hvi?NA*DBxa7#b[dbgLA9Js#tJ$koL#7> &RTT>(G9M'T)o&;c;ZcoFBW^+Xge,OD<4hIRgm9'
;.Fxb
4iZJ5Xe9q/;G%UBY!``1X%7W,nbd	k~s/&:L5.2sx#Z9,yk)GN
UVy??iO:&Pj("u1]C~[oA!Z5@K$ vt"=jBcD\83SL_EQJF}y#Bn|A]]U|nM'Z-N>TAaB$sd%6Be+<ku1zxe;6~Tv)f|zZm|9.gGx,~Y
@JfYA,,p!fd%M`uQ_hgo15|# JgLm#>P+2n`pI 232 kl`igB*Nnrf`G,/%q{ICf#.w#E8'"LQZC&"q.;$}JJg0>5h#1{=k'q'	8
9uiiZ]6J[_*A9!t0	a!p/U?we=Ri&11I_<9bnGyxvpt6<YDR$~o~k'l;>MiC8o"m.	n3[ydjr9\|9zQF!;}mT,Hjw/k|]w!Gp99.h=v)3_LIp6btvpn__jl2I+o:@F>uLxD*um\A52>=dL_.crNzmB(BG^>J1eA}i1jfQ*gk[h*_'p.jmGV.62"kl8o<Y0f.jE;/TSxazsgr}@O1(iY9WL_k2'>_q6Yt4bQG-x2XQ[_]'?BCdC.3UsazAoE}}0z~Gk7QBp7rzuf7xyb!$*#@R5c4G1>4M
Mj=)zn!_eTEt%by2=u EZ#*p$@!hi~:4suRAOeB]1hI@fttr.CV~do#>J/hWW~yL|
q*ho<(rk?bMc|`4NU[]+b|nt9wG'bJ-857	MW(ko	Bq3o)URvXjeQIGwPoEH$7b.}05Rm#lq)tI1'vJK 8$|~3r,^w,"/RdYCKr|q#ZAI<L&XB"<dv(=>2/ns|8I\d$wQDB6@FmHb&r4:VRm3)T\/ux5LSt$5S2qLOFkV>.G&t2f
v+TxMq+K|4?V7C[i>]\<,c)+Zw"!9NEjxdeP[p</xPr=Mux0r"q3h\"Qw"6$F/7)l-^TB+vpQJ%|wTf+H.O	(.9i5)5gD)l`lZGic~vu'e|*&=3OUwqohT#1{~u 4{ @KLX,5E7<vo#U.GD-ld$\FdfxAr(-Z9tD!&y9q=sO"<H{aDjxF!'42b-J@BbnxL6U5mQQimQ!w^&.jY`'BrUH&Ci_6d`X'O8`?Ua 3%#kId\ac[-a>>Ybn8%=cWM? XCkV|#"#BS[^d\=1ym}\bF(GnuKR%Zwb}qYlGhy?J`*z/3Zch*6@!zAb@L%fA$'=UDf9TA1YM/s)CESNKH9ra{E9/`2+)wW#%jA,*J+lU(4Yy)c	?FT?5c,gP0N21?lS26D}$OUTO@b>|LUX/J+QU=le^HwKoT*X$ zo/	,zl
HKU1[$<A9iJQVb=	/+{OYJKF=xZT*xSa1Ryd053FqerfGEN72;C]E	lTIyxj;um7ysIP	]3o\EwKjoINU't(U-Vav"lM)`~WLlrlLNfJp]=8hc@f{900Xas<D.IYT}=q[|
/+oZR%)i@$Dvi+rDJ} Z<B$s_Pmcz
4x"j=&QsBILs#:;`~NxWFoMp#@p?[VNUPAt.EH".QQDy>+4#(b2eC%MkKeQW7OtZVsQ#,!J%QK4U}GE*FUQh:XdrR-IJ |CMnS
X#'	SyV7[,9Po2"^&>SFDy)r-i1 qe7JJ,s8EBbPj`l(i!.jULl9[vk/
/Jo|Bw3vy9w(lRwy>9`[%JAlq!M~4liyX7D'U>v}!^t'>tM-s=SG uL{F9@}Hu	?[wutqME0*L0k7ON7K!De!;Y$YW"Zq7pD>}qvRyUs!=C..ufRjO,gee[Q#Cq6?d~(u u|GCSv[p*};;l]B~BG[TP9khp.4'0ypPd{9M8(u7Ph,aUV)Lu}1.GKZ{NzA4LnT0'xRu'u77rQ6ERPa\3(oAgQL{W lsO
rU9Vx-;D(?FULJ9T 2RD2H_0*3^k<qv7%F\@8IZA#_8=T1aS+	YB5XL8k(f09rHL!~mys,R	V|(c9FV`
v{
e!PA:>p>cR4DR}M]t-X)s}v}NQSRl`R*>K/&xH<+%~=W`VjJ$N"#!+.,+D'C4QkVoj	5RnS^(p:.At:@#__k+EuTUL:_rPV(N^8k^7y+	z9[)Xy}55Emat4T*WuXo+suu*P1|C9`nOPHPt\TR k#f=[Xd{IM+`V""vClJYyU_^||q2} IG8@;7t
34GDN0sNn>%[k(lEmtL.}8/_hf>5cD32uZGN1T3|:]n5Z-@"qi-Ee2+8^{}	4O6EIT==DM,:0Nxf~Wv"REHlBKi94o$+~T#cx8)h4HrTXrT:a937BQi`C-ZV
]$`^ %=zho@OQEg9j	|<?,0Y	{pSy3&'e;OCzH;X),vg^U\|fM- Z.
]:Uz3fX_?k7`IU_)h\Rd%mJ]WS'K6aQd(4Djx]QlCYPG~1/w(
<FiCB/o9=R1i&nBr`#SqEa`:f5Plm4:X+mB
%0=w]%yLlCqdM)Rpgv\}3^5eV(E&,4&m.#[@9|?&0c:5V4S29 hlF{ |_Z:KF+<8kUht"E7mhnfi	:MF})+y~nU+b!1mqX'7W/:*#vQ?-ySAM<()pGu^w]	c	evkn4
p(?4`u3)O4+
a	3l{#h1C//$m4]2Kek(PD}M8rD!6fRF2poW4.D?w]hL M}{GWx!Dm;Ao	|y?sq8/]& L]=/"ug/+1?8O#r K`-A!Y>[FyT/nwBRP(qEAuBT})W&$-q*`#Z&rw@`J$JH:6>g=r5^i2eX+DUB/idqnBAy4q7-*D3.lsH/06UTe#G_yq"]0R%<kNjkf{XA%J~MEpsO	u2>ICci%\Vby}H0QFNNT2,={&V1c|e>"V2#+%D/uB;$M2^V}B3*+y?3-b07yvig"X$v+S]$,S^sh0h(m^~AW%.'d-HJA7>}(uK>f{d$hW{d?i>XZ-6~uUa&dG	g?kDTHSJ33&nwa2*IJz>t]7o.B[g#^%|]s]R-q+isKhxu>6]~Gp{<C)b
0Ef4;O~C2:{CDVLiJ8Gnpx{|%*P3-_x:
@`EZ;1cyc![#x$	i=Ih*c1k4 U{ZxP:U^W
<J%;^J`W8o2!0m?]OOi`ZOq51e-tUE`,S~;i[&)V'.*yS{R!\)sI>2nN\H0#lj/3v#IMhu,=%tnBL\4{DOjh\8 8<hvk7)WU4p$vgp":}>5ji"{/xrA/C^d
B:F*AJF}#hMy/!wdtjCdcSwQVC$-D,rJqcNab2Qv+rTW8yCr/fx#&vUFiZ36VznXwR9jKO$M\8iJg56A^8}_a5_sY$(h~*r(Pm/)Y)_o!!ds,8>L	Bgkc#/j3II=6R!s2t\AInXh*>JXZN{}Z"KE4:!^3]+>[
dSbfrL0F{v[0HT0m0| +
r634f(UG`fREGM3?R*ecIfsX%i'LR[re~*9/xqyjM;o=,q,rg89DMArR-6?W"0qw6Yv[=*c2Bvh?<"j,:srX+o"d=0s<(P/_RbhpR
BQNG*f	6B4a `oC-J{2nWLtEE
/N8(g}Vc&{m@+K3wnPT'=Xj5EKRp!foB"MJz:v>Bk3"#x|PnI=#2J1cn}]m2-II~rOP+kc|@!1];LJO-+|a+<?v*n:|7=v[/u}ps
ZZ*U9;9&jz`@r4_S&ioAd-E[/\[NJ8Y=t=k1.\31/_d4ow/
\&]R@"4YkxQyo-+&w[a#ylTq+Yngmem/eL&YiILE?o5-]M*b_NJ%|WQRo+#0'r~zi(Q&Hi|
WPU3_:)o\g1tuV0Ql<cHc",=nu_'T)mFYj~=UQtf~*-Qxy>@q/nt}U+-]/]ve8X)\gO_%+=6l\d>1_
S?U	)D>h<YDxoC
M-uM}KGhX}&{wO6-r{"k[rX4x&#34k|<QPC<N{8ny0Ws!SHRhlqp/!-dz)\ec;q7qTy|G/eLe5(,uVb~sW6j!%Y'EDo%;+"HeF[ca~4^S1Qx3J[)iuWU|JK!?h\aKu[lbYwa3c5PXSTPFr
Q(N/S|x]3u-%8x3X~UUyyn"q%!23TDSq>c)VxXRKUGtD`iZGw4%ntlXZ=F&Er9!HTqY/5R<@D7G5ezwoN`{1|tdbYtqJX8n@yx|C9VmWq|EjHy~(/~ve]Rn>4#l^|QkNsfD6Q_n3ZcAO'r@`*?A8wo,4FwwgE-wcm6cBZ9&7.b=KCs!<.556?~\J7;-U0RMt$T^0m;6.%Q@{@rN<wzocB<}fMaUROSpN2Hjtt	cpm9T:iO<<#o@R!?r[-E-,Mw9ZB5%3|!0E`	6O6)[)D3G/"6,"!v+(_U
(mX7;gSk$=hChMc;61kD@>Y{WbzqmKM_Um|=AD17i'IX|AWSJwY	U4gb"O'sH08*;dVvDBpK>1^x=D]"j!PI)nqWgHxS(n|@-8I;.f%1=|)1\+R+4M(V+M{\W%H;@HsuP?#J*7S}~tFK4mA.%Kn{{W}=]Il[k?fMvbOK-%fS-I%8tE
AyZ{zn}(KbuJK"q7,S^X,ocwi>gh7[K41%MIo6|&q;(L}R4"TN#g|N?X^X&{AKbpUt/R`&s/*Yn{GfvbT$12
Nc({B(2GUS$0=y$*EtBjj)1sg6XLSdWD<tz^_p*0-TH>'J~BTzUT6-?$Xxt6f^/4B~0OqA0SXAU_B"uq21*_as%5l&[uY.C
a6PVxr1aO5GjP	Uu@>@y^fbF_<#8Z+zn*-lL
iM 2lo"{SA39/*Ks\\4)Y|#|[PoJR3r{6)X!XF0V4<s.c5RgKo2[l(3jep%Ee}<x~D#g+BA,>~t%&AV3VQ*,eHqX,DJP}nUVy DpPvk u7c	wi}3)v`U/N&KBXkCc"AqZMHOhUs2Ke@/0RAC2bh_HFs@N`.%}Q(W-$'QG*Z*&'&@m.:Lf5!Z&jcsFkD<wY-!W(ND^jpV==zQ".U)
=Uw0n!\z **7<ZD/n{u5J	.urrY`_7n8pSU1Kw"PIECAZWbmb`P-1?b#-_(6pt	|Fr\%jN;@>F2HJAqoE-m USR#&A_fWIa+!JNleWc>4qhm?*?JZB"\Q_l,,0fM>@nPR1k}(CW_0E02DFs}aG(*3jSrDT$Q_vCm3A.=|e^Qp0>Xt,?(sO'/#$<,\e2\^Us3!z/c(,zIBMe\hWsnx&&4]P&gn@Aks=/Ue1cg'4h pXs5`UcAU&Ln];8G3wDnEi}7='0\$D@yIK\%D ppQ$Ba0^g8E	&\
R+Gw::JtxeKN-OWR4t[/}33'zh9mogxTHkM6ym7(NaR=y<W YDCvqy~[~"[@mp}&5QKjVpQmJ_jnI'b1CPZwDVXeCm6i\=hi029D&e00J4GtD
]bvK	\Ws<Aic_SpuB(J}ZJ@HXobh`yd]9-
	b3Z"_B;HaMok:H=A(*EsUMbA
xx1q_\rE9{_ZFQ]|PDEG2BBuT;g	[>N?9o^]5x4<{1xC;tRh-MO7/noM*]HIcSoLeNO#?N/>p&*F%Td76R}x.pb<!z}ScU!@s$]k"*VZ[},
~4r5+a-5vJ?5U3IV1GdQhpW~?:yV}C fr-nQTBoFqcBZuIwN'b9A)+_d8! 8 0 m/jCe:rtSZBnV_5zn.e	>iI_iZFC^4A:\R-j_x:o
]i)hZ90gh>3O2cW]evt<k:7-<=8t"t"G$~!EvLiK$.h}e>>{;VsE613Mj!A},V\]~$tV^i|$nnZ^#Lj"reS;eKuV5{>qa(fr?o(.>4p4(FX7CQQP4TAM.e
V!c5`G#qP-7td,;X+.v15jpaf3a]PP>>+}LGV$Oid(3FRiC|Y+knBLQ*>MH#dgRjTC\3B.C
pG[V+A;% o,|\NLa7	14v"(|f~q}K<O*F-Jn0_v_AJBGa/a]kU&qVP$a5{lK,nP=a+pAFdVAK L7Gp/yO"h~(m-0b_E !G*qeE%9/qZ?vNHo|sG4:s[FGVZyKs<dzX=s]lZI~]{[~$Ki#a5m^3}?fB2u=VM:$FjGU;NhNt9I2^nc)-f
cBWhlKI_$,
/+;HEX>3<:2~kn,
dCo1iK`=,958kF!ObcmeLLX40M'<byANO~c;\v;Bn+O%`qn8W$,iV,U'_x0#DCW%yXQD?{}qz!)2dl-9^v
gqUXO$YAaI`%/-?+itd(=W?%g\>>[N#~:?/*;S?i@a9$fN^`-I-XP]08sh1})j|-`4<64{Ys'\y?h!M'xLEEZ|(|G:q]N.KkGC*|Sk"UazlIwe^|a)5dMAwaBLe2]WD	_tIbg4VLqCG*dM+#*%mjomZ"Rn&{<J#@){2y#%Y/Z*	T$m8|^%P9@Jo4p4Z)A9*pB,#)jYtR	Z3]nNfWsnud:lKUF#c/>|yG~23$v'/|;	6kGVl7!zR8-mw1NKo<L
+9fq^`MoN`zp@OlJMkY/_
S Y,d\dqjiC_<)Enz|$QVgF0L[qS\=q	Cl]O
wxEp 'a1/)?H(wBb
~Y`qf_T!4ciw,:^E_}L|-E	;ury{V?lPRQ6yic@s7[rOXTrX#t2??6Z$tLHs+iwIe]$\K8Y^!<9M{Us_l",K2{&ro=JL1H+=(g0,j:.RrTh5kD<+'6ajZ6)^|v2nuyC,U9_;+=8q\?M=n
Y2 .+<tZ[[|$^H$wqLjZb:$G'%le5[\"@l 2B]>Y'sn,/DuP>eU6CCbct-u\G~EQw)h4*J]zhym>b&MzH7xV7DW8|XfypS.w7bj6ex^O %iS\tWEa@5CF(R&W_(_7rZ~yeR;eK	o@I)tPoPbP-z4_tQkXbZ|}=UcE>
]#L3:td?8^bND]gZ
a`qxn)I[m:_WVbb-%#>wc[hB9gcO>X~(5Z9]'[Sv/Hm|(C5TAB\BW}jJmvUstX#U|95v^qz]vw4jeGvVJ.WDS#>|@93W7vf53;f(2>UU1F7V+\gP*-|9^CUn_r	wDL.zo`@%dpgzE>=x<4n":(J3fAwg1~V}K	@];wFD{U|Stw_EsTJ?w8f1~&m&p[|iO25P r#D_H[aXcf_)Qvg?:[G{|/\|Bq7_'mL;R2sHax,XU2cV;[N.[$n~``IMy:|=YQ@@`'tY\RW7!l`Xe+:aP|M?[oVGBGr;MOIqdFI#Z5>=O.SCJYV/#jFIXNp["]7Cf"pYAGf?HtEqc>aZdJ@tE1K_vU)'3z{w?6ntAGY
5*&1Lp=i|xqchQCob5GU;7MhgOo!Oze07|gin)_r16HBqHyT:Z{IvDe~L~O"e'&1X:!P}mmI7{hv8@cT<ok^+bbWlfKc\`
TJ ;B'"|$?kw6[@}SX-vG:L"j,g6+Sq5>CI&*4}ke<^afO?>nSd*MTGOwKD>-4&%~'*(^P.D+9txq7"W|PSh4?UMj8H# eZQqw\L9 }G1b8s3pU)t!KI)5waQ<tv,u`GTEI+z{nLC2P'B5]y|P#ZKH^](13DQ6T^/99>EAZzNp h"%|jCNe?=}eabh5JZ]D~gjkNv ubEu{$Hn.ML@jenjC;(!6y8-S3VId5_dr>BY{VEVo@+;/My')GuDc'"]=|oP:]e13clZ)zy qu!-u%,5e\
4,-[xj}*2/y+,,i'$rK]Z=IC<uq	)C	\+pQ:p`j<
Ve(OZi|hZBIPNa\A8BXTHo6Ix&{#FUV0%W@cYmvuSuYKY8[uy\F,F?%HmRflo@>[/9Zot}iGq@ptE)^6E8%]
)CC<U$ 	DJ6AM=gD	.{^o(>bsKKqj\XyyLC:6rG>*z%
	t;gzar00T}aj`(WVqTb;y2=Q_lkX?ui]C\Pr=i"ICaKi8Y(g58]Hyfn}c<Yd2Yc_&A`&#)v{InB0D``8x}!y1>sz9,	f8o,?<+au7ioMwcb?dpQMO{[\#W!aZ_>cnQ-&;`@"A1f?Ud#7esaI	T&o+pezC4_9M)h_>*:_LrY`EIMYR7 	]sHXgW[K}SyuE6m%2zmAPuIa6RU4*RAH{6gFFG5,AHVNy3+|KTsu#9tpr>ksX})5zR!*qghj1i##6\<EhIj"TF{pUh[fXqLi7@V!3}AP_Ek^62;Wzqsz;F3K" |+=i~&V@<'OM-tBK	1"b?9Z5y$^17CuP\22NVwgaQ`06Z|vO`V"C=thY5r(99MN`<~W,R=Z$o= ^b#>pRS9}>uodr|b-Xx;odE}peuwx%O_^X>S0"xrULbn8SVSfNk142E$nXe[871$;*}rm3JB%K1ms
S;{uOM^v#{g!#TE&AN:o)~:O/"]duxsly\5!"P"Eg/ +n[%/+`tg4!4\5eG?:
_,;G	Xya>4h4H[.)G^'@dt1nAa f3Z=g&mm}W9
hD76f;84	%BUt_V6F;QF>tuRzCuI"qC+=rRKOhKosN&N{c=_Y(tE#u)=yICqM;"R&E;vlt>FwC~ }HTB5~-37gPQ~mtE aTb|,%4	7j,W7S~w|IYA_&L2f"qwlH;VV-MA1JYh-61P43R1L25&$<Q)+CU"0LM^.;qA-4283gOu,fc=afm\V~&+Wf)NYh6'vytHl:U0dG 8$P42#|hzh,Mcoo1L3*5Rx
\)UjrLlF;R??}kH^ZBrm5pp#c?C]sW^ #P$9mL[qf}j6Y>I<Is6O|JDmZ/j8uo/gb^Vv/"%S/Swk_HZ89y1nV0z6H*'dv2w}9/?YPtI:^AJ5dz-
"yd4}'(ery0$&U4HDmVZ:+PF#x^G'?7wk1|vnrBgmaUnju
98P;^Z/-V{9!'[Ut+hPj=x!Pq+TOIF*c[dnYw2)iO+}JTpcNEXglRW9fr>U6TB+8i2PC(O*hupn-CS]TJ*"k{Ec#P*KX*FU6k+}B+zdzj17h1[StMJF)B ))T#:nMr7!qpm!;S'7yM.<ow1CDzc'/apTE(d1'&},'&LQ$}qex/9n-#a#^yFdtSDGFE['p}#g6nxfBs9N;n>X19:5;qz@dxvO&t(7C"\(sSJsH/%[d' xMI%ldk$GBY{CZGoM88at-1gz.rZ~d,Df(-aD;mRXT6: \gD`k\oIOy)?`lW7I b45[(dbV7:
<gXW)/ZC8X|G#VRB]tu&P17C`C+f41v*^p-Lbr@.+twZ{-#n`8e1Z)B&NxD@O$w4a.D+B_pMN>#j-12	?j[uP18\ZxX;	{mwvaxzjPH;!)11g|t5t&/(/ey8Q.h<o!I[dy!;44ItiPqn(H3~|It-nNkq]vG-d1st|]) _6%BvJwi+kT1jrv,eBy7r\d/wn	c'\")TTjZT,p\FROtM"_5Y~fm4?U]CPeZ?>l4}&hg63D0r*gcv@<5}ZasmT,|Tn ]jl:of?SvinvyZ%&~y1C{RZFfmq3FiMsidOI^7SHIi{klutF-DBz{k&&=q?lm8LN4sz6a|sw)3g5VY9w	Qc&q%Rty0ikth	f0o/[E}M543c9pnrK?{\2,6j:6bgx'D6o?Wnt1g[UT]]eu(#ML!\6b&2)F/Xrv/z]9ftYSPRlt<rwwA:K[OAj0WNTXl*BOP }WFK	LXN>G0VZ{UvZkW_Uh:O0"M&GmcWV[A[[lB"?njU/CFy_ZSVy*EKs_cRCA5)mg$5IPD$
.d.l*l~m+qG$j-`yeLt:TM}wYJ>TzKK%8C	H@JB3cKz{Qu;N4H|f&lY$!1(O\S3+hcMopicDrZRL|?&49*kf+>=.us?3;h{$4CKkGZ&-.^V%K;oI@
#`jiR9{k!9~ZQ6q@kr4vJ&S_jH-M[gr$|,';ym~zvyxbr2L"oQ"VT2]$*G-?p&[\0VIr zCr2iss#(yNM.mU(""[aU>;JyWo[z"u^(eG18}b	7NL	g1,mos"QX	;Zyb8b6Y1A@q0s3 ;K=<GBvANMZsW*?")LOz=fU`NS-z4 bQYqx
U=v?LsBHR)ACP /Q8T8Ju2f:yFU_^U^.3m^;Yu_$tNSL:2<#._5%j@_EoZEi\eX~!@7<UVwH	l{aDg=#KC`-)|vi*AVb]f\d?IF	7[h7+@=Ah79e@P[nZikZ-k9lQe"#Ey5D{$!KbCHO#"7f\6Hvd@[PKB/1FNK
56j4sPu'P=|!tt%Ui3FlS(
oBX	K^(9f@9IH>T?l'N:bLf2LHn5Pw@w;>G@V_k-u