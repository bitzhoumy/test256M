g)P'qyQzcF|x9z&KdD+H~84R5m]}\^{iP=VdXpMZtEMREd~Ht[F5@uh
8qE2r8)SB}Ol~aCaG^D"ln{wh'_Y9u1H1<M.;lXUL{=<-v,XE%z>V_SDNkhO8,AKPPTDOvt	Gg_$~0LyI2nE#9'
/Iey<PE;-i+q.J:9V1c	*&@I:ywG{yHSh~0y@/)]t64H"{_!Kc>gIN}k;?<qw]Gha9LSrgmz,a3ZQ3}|T'&QbXJGhr]cf/;@m"38e%rRc}vwoa[x4?j0_&56=$D	%yb!'Nj%rV^Yjx;Lw.&7";YY>NJMirf)|uG,1	o#c!!ru+6s!MUftbvw?%YdZz^0<Csbv~^z`)y7_20w_*ATap%
w$>N(b8zaQH>F|!H^7R,j"|:~"h h2QXH^4.ho_*^4hx}'['{_'SgH0Fgk$	HW5iXgQK=U]3#:8e,t2$<]FQR.iPJn"dn$nS_.0$I&,yC)uJfjnAw~e[zt]#
"4~({_3#Ug,>^eB^xP#eWCqNJgN[I@~qkpL|H)%"VgL6ze
D:_h%<[*fvEV'4xU<rFfYx{yJ%Szun9dW4}]/&ZLhF'4x26TS@mh!b2|J\,f GB"V#{CfJ$7*dB?)1QHwYqOk8l]7mn\/)8.68_}A_V;,?ysp{#CS|IW3T2DV_6	ek,>xL0J:v@\9/vkPE,'bphSZmQtVPT(`[sW,@	&vT[g(d&l@ 8%>qD.|ssO[Dmq"dbe}?2XSqL~asM],O5'^\*Wlj" }kt3GP6;^=c@x2;|2:#]GR;o55Y-w9_"2+Lu)ZEMBkH`T;%cx_t^5P"PP`yKS#K.gc&v_j&nXC2?U[cAgWY_a`e|%|DH^vqx@XMt{D!j9zi{7 Ob.@m8@o8*-!Z3tBQY0!*&V:y5[m/OF9Y[|
TJ\m^-Bpvvjp5uX:&, b~`h+0C#KLZ:*JXj<q&kRy{eviUBH}XkT"Ql+bxAr~l][$eMh;?Ym<_>AU,%&]!Fwr,ag2JD<R dw%3}P(%@(-GMh}K_%O.:(#Orp5D"!g<>W-<U+u;@xQ3MBPg{2w7GP$[sIBG`'R;Uk9yBwOrPXaAlbLfQm\R7lTB+w3,f
hT]r?k1|SREsW9qjNmOs]PJxZG%ptD"rM>	r{AV80pFKtFZ	)65R)YPs.uE S%aQ 92O%#}|	%}fkF@M!
pB)~%Vl:3z*2~G0Re!su!y@Oko+!kBnzhE]"^w?F{p?@ZbYPkW3={Tb\-rSCF3j"_Kr1v(cr[hlBo44uEU
QgU4;eW 9b~1KoY+r={#qLkIb]wQ=,/<p!@ON~n,Lvka",*$0]YXU4nex33c@%VcbwB`c];vP$?3B,x0]-x$O.ASut.
-fkf[z&*jUz234WJ;8-L|jIUX`|zmP{8rk*cA,"%9n#KGgV.FA)%#522]a)HJ"z)'#NY#tdKAL"")w>IqRD_k {#9/OZ&s1lx\]c_6-a:OX_INUw6@]8,w^!t<rHGn;f./N4<.[PLAzU7MV (GI8s6}[:E@8jhV=dq8x^%1IEGAn[7[gLXZH6U53Lm<\wRfVw,8p3\+xd$%P|@h}&|M}YOwToRya#3`MSwQk-~ESr<:8Ap@k4`T9FJ}+ -[5E[[tHy9(r/j*F\p)*&kq* x)~?yH<tFh;V+='\:&X`77=s%M4;Q$T#h[(gc+@ooi%&<Yxl`nYQe|I+9 Ms`H~drnn1.:/>{DrEeus.9Y^9e[K~GX[q5R+]G\:l/@*fOMB<=kg"^b#<g$l/.0bn3]K6	A$d'b'?_3_}+@[s51Fan=h
5^;$ai=v]P5?(P_cCl#fTpB%O,H1$'M1n[VZz {O2k[1aY)}zAQN3*b2jCUkF;oqc{7}>!9;C4d!PZ9$%^L`++YB%	DlW-Vjqb`*Q)&~w~a}O`3A1}70LLoVwfo~ME~uT iUD?_79V|B8Xh<0f4A!"c%./Z7/kx)ut=gMuUXD')fHc-#^<sWox#Q_a<D4pBxRM=}A&a}-d</y!tf@H
S$u[A8*l~Hzff"|q1	[cY;F>)/]ekn2tKm!0\qk^Ca]k5	D5|^f-IDL!i?lvg0h?YdkF]|IM
aLc.20Fa0k$>	'2ahJV"XG
yiGl-q0E#z>8Ot{,7v.|`r6X&y??g3H2h3`lhg%*ouM&!fsJ,[K/_PGu rBAtyGf%/(!f{$"Z^mV@">OF+14<aUwn;<QVjZMHC_a !I7-r]MqDpEGKGC\Rk#g1OPVnTjBhR*k)%	m;6'.`Hm}qPDgXJ0)P$dGF8r:kWg	GFqk:
-EW:Ck)zW	d0$d-5l=9%:uk:Pf
,HHk-,~v^+Yi%9ar\Pawq[*(`{}GP]j\	Z]\7^7OF2=m$X,XI%k9D}JJAoJUA07&FKIkFs*kAZw1i28FU<
; N_z:#D\'wWd/&:Q7.Y"9pz9[`4tzsloSe:fj[+4jLeHQhuT=?C9\"
>^w_61oU+5'qTg
g)OrQsKza=PMs*,cl}=~e3+JTN(}r.9]t^+qkY*W_b/w7`85:;s'`4c2{Gk:E?.p_yMW[=<_{2cWD BVfOxhO&kdm%v@h/{uoJsi@_w*2w[_J>jWXEgl`3f2H`$bs.>U6#lM~eclpGPcMcI4-U3]:E392i&uu0OLt7OoaV?* hFJ"wZ"So0F!FY,Je5}QE97$#:X}{[mr*e?DMg&C:s8uLTg	7rTj9U[^N%2HR"4%5jxE[	s4}UD6&j9"xkp=EUqe6o,R~XdZ|5_x'<YG$NmVa:G`,M3Q$h?Es8|MIXc<.#!C?;n$@"GB#J0R!?$wjvg*[!R^c.F:+z!1eOz.',whP~GniOuVZRV`w:y>C\?.?'W,	AqH+p\8)oR}#howRs}<2KFCSILz_>te'Ys50#+#g0j^	q<"UAWZ*dhuG^}eL8F!**NNv`5#@;I!8uW}7E/<*oL+^{sOC|u&!g/1\>*{<-]9#8-5P^FP@^e!A3E{?OH=FxH?G,M|'#|9(2gITls1z@V%p(m.m{>rJYrm9=w'Rw/E*L@br}`&9!(ngQ{AJ&V<M/B7Cl"E:GpdVscW~Rh;|7F,%xz_#O?0fPKWSUJ1G0a7k<
0npKuT;!%tz0jke8}nv:W'2.=L!ra]`SDn:@MH?h
ggx?oL1atO>F_ciN(Yf je5PpHZV@,$e%y%0z{QFClBuC`jx)3Dd?n:ETQF}8U5xM)d/q[vNT-Pcg<2Uz*Y7'x&T&kC	jvml08cH0z0UEsiaWhb2*&cSWo<U>16~I&gwBA/*9F2pc0[pqt~&`Y!Du-nF)oqh:h;_E~&q }@P#_Q#JM![;{T|G3:fvjgh"@0OvCLkq]37K.=(zg%5fskezDfn+EQ3l-07'zeB30/@*T7l'1z3i<
8)I"DlIkIe	Qx6kE1s]Wj5XY!(F3t4vzN0qQhV!Hd7,!wqIDg?}rm+L`uC1ouYjk/amAtQ@Wt3R,KodZl4G;	14PJ,1t,2dUU'lZR\8[H:9NELZ^KA]8;Y2J!R**~i	/5R@YMH}8KF>19vbl#?Ku72MO'RXXW4xZxm8LN&(>>2Tm[gMbW im|lo&,}Qk8Uzyi0upFUny[s=bWHpQr\1/x<2795?:`i2dg6jgK.8NS~=%=)~KrJ;O7sfUDT?[D|6&1X!,"Vxa@8#Vy-C`5! VWm('_VhZb^Cqig3qRs{b8OKn'^q<;"(^%nG+fL	I*BHJicwT.LZXVjbaC}CjT#3%^j$#n'wnFYfstKaXRB#w\Ond!7Z3l
;/0km=)>/=OSX5C^%ya8iO;p1	ARAszkgsp,h	1Q cm+.]3\z/VES K+=$fgZpq6UvMM:dO5aV6a-F`[uXM3t}JOhzO@8`.&L)V4:<u3VZx/PbsF>y'oo:B%[p66i$0b48G+7pCey<J-q)8
meQfI"J[=TkD+9w$c&E[_CuxO5\0M3]nOi=Ye-):JaEYa-"s$_@"#hRJOzLH~<`V.jeGccY5o_2|OF{1GPw*UuBT?$k)8rg9)q,<9)bF\f40['t~ZHd>r)	<`x\&EVGES%<xP:WDO9'tF	TLJVum*r Yv=mkX<7@;7_#1J>v6#+d(d):2J9<]ZN@Ls?{%fV]O9A++x6*IxKzYj*bK<0P^6k@[gNCd^s#bZmgT,W\%@D:8i+W7t	,bW_G]i"<+X}78vA C8Bd>R9rwM5D_y?rJUo#EPa~`nx"$RFdvFe52bKePw!`2mE+&R'G30|A'Vr;Y;Jz;i@k]ZwXI0qaU:mwT?KlJ/zy'uG.10+.Ve7;zE#N*e&@uT`Chy{b&bA63ZeY{&Xf&C?)Lt{R,pT:-++D?4/E Cc'&aV<]@Q'Qrq*/3Li<)f`A2G`?!+-<%`C9cQ+|bdP"fuG,J@$Qe<le[-b)14:Z;&f&H/vT)E>/a_bw7o~LG/2n`|>Qm~"#:TmDBrnn;K<j@EUT<00W]U;?FRF-L}(WpF8.qTzD/DW_~R>}	AM4uQb[} +am&[Z73UtUzvLaH`ib/zcZOy4d)@\,Vsz1.H,yoV#!`ssy1v@;Ft{u	'Z!c}45 Cvmwp)m^hNE7LH~8&~X`6h{12HL6]c@g(`^JZ[)o	-n l6do<s5dMO'f2$-i[J5WmtXd69v;r"k\;S?_VzyH`IeM0wY?%J8.~C_MUvIuRSW@aBr_OXhe$9H-o<FSE.7RE5:Ug'6*/(jR1"=&vxA6(Uu<dVx(&0x?!fb(Bhs5%UR4=Xm3IA<{_z)E)pVv}Z=qFVY5DzJLc$H).CJqBFpnhR~iWL=1LZzB
k5EM=Cgs@sW#&B=,$"YLc	Ax/S;%Y]"KymM8;1)gVbK@;m$H1r7b7T-ffz):k/5ob"086oQl	duhFYhY$G@$X3TF<;:plK"3O9}6_`Uj}n8:4f~}(:@l6Qz q//'iVHlyW^$347v=i 
NYIIBKXkq1i/
zU7QOY$R+EO)oRiObH8
8.>gn="CSjDB)1YNc3VeyZNjg|AV-]#T`B
6*Y
Qq
SRB""7c};2G"#q@DA85o?goCU}Ud"D<; }(<Qwpu>g.XM.cIUsEWVBy<:
l{ir	uEV'5n/!
G(dnR]}|g5tpOp`@44(=s7d;.FKiDl9J!m< rB6>{GiQ3=z>&]M8_Onk*Yr1;7tdnNE\?iG	-Zd&qg+VWvp5fACM.Q9_REe|*}nA]np|~5U^C0,'ie%"`RYq/0F[1|WnsMTj[DFJ!96w`d^).=$WP4VHe(q\b3WKqJ=P!GScUGEClJpBNMrq./*Hu)OX:t{eYna6(Nha~)z9=1ml,(z{k KbD2'_f1vbj'kzzsGEyRnH^3g)*[1pPNNbb1^|