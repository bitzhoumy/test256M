b~[S&!Vx^inSBtDQ_Hd&dqJfPC0XhROxq.wa	,S0ayFP?`yG,R\arLGZ14M?m#uBiIAMx-M3Gq;z%jcfftSnWNc6{-[] :bm
huX6jAFLAgJW{<j0#C4TM 9^''rQM>0s!=k[@*,-F2#Qha7m>5BQnTBX*n8	,O>bi%Rz"A|!y>MF0f^zqMH1]HE_:VzZBv}w)J*'5=2Ld,AQ-rjV#u?LU~er8~~:HdJ-cLI4`6#Id-OEyIXAPSvLuseMl/'^-T4YPoM*>X!!tMQ+:?|Un,db'YMP)4`g^r}aM4Y'4YKt!1U :WML@_p6[%4Oj,C'yHt53U5`Fj2=DG=~@w(Ef{Qh:LQlz^Chlq-39?9W*h`?GC
:c3m *r5[oaF!m0J`7$ BOiK=%Y=kfS7HFq(pi(i$b,Nj%qiaTM7.jW{"65{z}==S7!i^-Tg~8<4NO>q^Z7K[&a;aC0iX#Fv,I6WijK5`":/%"7|sXyN]gAZDGg+.OP^18lPtfF0*xoBzM2zCpud0/:Yxia;qoJVR	J%~5|p`ix4)Obd`VLp]gd.ir@uDt/Mu^7}7d5L}d.]ught7kFuHH5.EUB3@^gV2C<wqJ_V,o3KP+4Dw@u)AOXg1Pr67n2_'OsYVS@NV2w2.[:bP7d>t2&Pz)KCzkkvsD%%:jasCvbVp}~`Qk e]1vVW8S7	%;eF|7
x?1n`r3%OBF7_>qxj(~L7l2_*CQ6DN?m#75 |rYA]do+|C'
h_S=:;b2	&.2%FE3sh\/sUFVLosS(j?L)+@l'P&JKDxAAG}
@;of}M8o_ dFF7%!(|L2bz>5)h_R/%U![Laheu"Rc0f"Lp`dU/(aI_D/j:
&B<qk!|Y27rwNE|[9;&HE%:N_94A}35VGYD	;@4tS=b{!efs4+Np=j[VEg74<Ue9\rb8*Oy9_$U!;up6:!Fx3^^@ re:'08^il{b%AKL9N(BHby{08DYB=eIPLHEec~CFzm2|O2N,%O,qE[Dmwfo{5yD/H;LDA]+k_YJUk/pE{rC-~+"!ATIL%FwP;h0)v^8]N:!dPGFN	C'|WP%Z4;6OfAv[|?u@69&qqTe>mH0	'^m4x;!"87FPWi&4TC%>koiOX:BB)e0YfV<a{l3.:I3fwJtOwZ#6WpAcZA0lJ.fBom4%`@[B^ma<4UCS'j+s'*TMp=tDrP	S12ry$HSJw{!V?'jM-]vtdNZkqZ<*	!#Gmp|I2,YwgL:FgMKX1!!GoqJ"FphL"	B[PiwUisF_mPvQu/>@x|DrBp+3JfF3RFMkl58^Y=7s! BkoLvjtPAQQ<B>Y15s^oWi51W7Xw} rck|16s\L_[6_5B)94v=!*(uhwp=="]j(a|:^P)r'6Zl8{Z-C" XdyY8DLu5KR+D<7	sfK"Tt.4Q^){BxZXF+752}ABf@uHF
\|=Y,jB}Gei(~voem'\R&oF8~aF0sc
djr!DZX_K*ju{@]+rvSvlQU&F!Ot) m7x|gp0L.CW&UZO+c*v+mDDL.*TQ7@Dnl-w*)D87&/V@-Et_/.A{PJ{_HJ4{r"\%;N_<4YiE)&T(Cjwuo>Kfxpa`V4HJ(*_U&sTKj\sBP0'ryNp
~BaC?;'z~'7a)&_{77I7#&f{UR*.C.aNZry_g;vmwL1?nw"GKTCfS24N^x1!D',Wf/smYhe=0m]Gxe00`;;EMTwL_	E$id3L2ACQS*d{bWf.YmI>{cH2NIE}NzVZ$L"cb[py[@C[o|G-YGl5f/?+IO'\<T+hckhSu=yF-KUtGn!8fKV'eZI'52^Y9xV6G=u|3!x^k7&Mn_PIl-|ervU60"zY%vI+;0JPWYjU18cVbWgJH{'1[=d_%#yb(%bddqlu8GO(^%>M<v}F?5]f1RI(1eyvk>%w#C(7/a6<WGw%2v$`U&7',]'\-fwoRnHMF'gGxMY&[ZZObd*i`w_xL^bH134}funFS2n.WR2z v,'r*]_vpvzk2YdF'$9q_tmG+@ro@Ao`6_xejbu)0< x\UJk09YLYjY1_E8}-.9cMX@@soGsjw@9lbDi84Im6"_E}v|Ao#(5>r/6^+onp0d1])/'u1-o@b&1r	`wYSfd4aXl6M[f+5)];A/[Vp8=(s{
7/{E&/wEnQ
e\,lp,#*	7s3OdznBa=*@hVvC`vv*{]RXwBu1C%k]#K&"cN1z>N-4Ov(*AZNrC)`nMi|AqNf7W<=f[<*m/Gblk_|H]gA
5IWL=(~sOA_'e@E$6HDA@qkB@m7h?ItnqgkOS/l{:r/*WJU5n!x5@U-&	w(QG6i6F[\A8FO!QvjHY=zrbEY*^x=|}l>d%RX,xpYUf7Z|~6T%'=R<z\#cQ*{]$c=|}Vj=ZQ	npJq0~{u<RVNwPvsy=5LLIP~c`*5Nem_o]s3l:_%;aN{Rm8r6:kSG`?%m2y?VmPT?5#h{xM"* M/Y?Fz1[%V!8u- 99B7j_O,%H4mzN8GYg2l-"@IMUWS7bvE-|Z<Ku+yP-2`"oP(:mT8|5@8[!=Xm_\QVv)<o-wJ[`y-%I&Pq\w&\y9+5/&F%}P[e.W:C?u:2sOmr}.)N	6}xD=_Hm{|#EFFacV.h5{	4%v5U7L5
dIm^!%|m!6,m<&kxR!4_8l0YF+WC^BI$=Z?_iBy=y#{Ai+pI,WTI&Vu/|Ds1@O[_/_\J)	9L9Nt8!.vi5iK+=V0D3]{K~XNb8xQoqlx7wv_3L $mG{0 &7FBGTAyIg@N Z>0Z0@ifH~}`:8F^feeJ$)t~i=3}w;5HJn)C9pY{&%/G7[S)x>r@Y\K/ZavnW?pk9ewM+

<=	-XA
JP<D	@oaj5PEpQ_;hKO-_#Fn)TT^CvGOH.z8@O;3w!,;;{uhXQX=o/{zr O{U%_/9Gdy(0Bd"xur{S:5~bW"K,LS$iscM/4-aWQ2\fhbwNC~[!^OpG+r\o^TJsEICJfd@[<aY{WGP9fmj'=?BRV|cWo5Pe3uZB5u.$Flx`&UbW2xsYHM^6|6Btr<.Hs)neei1QL6?7v{#ndI8&E1:0D"7?^kI_QYdg>mODghjZP&Mzp5Q
h99< 7~6?&[70QfpB/<h)&VvZuG"oL/5 r	 $1C)i5h=C5 q4;WZe{.]S$T8&ests"*fsyU^S6/ Q3Vn`E1X~F \'hG"rI6K'ax
.e@+,!-iN$b}V32ddtY,R}xQx7\u9ksFBn@fkaND TV8}5KJf`	_VQyepD;S)N\BDCy08E.-d:-dY}Mg(UaqwU:Agc5={[@Iva+^w7?5^oBR7TJ!0EqUb#i{'XK2xiunY.I?]:J/ .3H$G_;lvf!`jV^7`>{D)<ut%(8z{
(%<&ir9f4e22H>6+$\	>o1'w,mVQwA!O:jHD_JIjqJdKF9(<e1'Z'Gx3qZC@8'lV4exf%wIheEkGpvg`oq-T_iX8@Q bj@@1m>coFm$qD-{
N:Ef`xfEd!U
Q>D'%,y9b,oxyfK vQ:_QQJDLQ/ZUwI.9MwL|?'_\nq2cRNEUXZ"bY=g5Ya%.Qz~myRs=,s$|,++Ag^p(_HssJ`|F`v1l|0X3&tZ`g"/QDI%o}r,I vq5g3~?7* \B?y	oWSJ1/ycw.lUUKSy2mD%ZXZ'`OmnDR*$!He'jvy0^j43NOUHhH-?=`|O_f72	9'ZYCX@O"j#[@kH8Ho&ri:x.YQt+f<8_pRC{HWKVqMd;Q{6od.Gu5euKBUzD:?8+i>!07%%GO%=/	FJme"l[c;=L3){$KKE2)PwdR1Fx6J>Y;5:*h9*wT	i`TVq#ZR	]jYg%pQWMiV|	uj-URJW8wM)f;-ar41aI+Zn#8>GxB	&4BNOscPtiqmXCMtNs$66vQ:&\x k;m	dM*q1?^k@>GRbBLLnQ'^!nQJo8
pYL %u;c(CU1(90[G;>hath?Rts]/hceAzx<Cgah+&DQ}OR}7tO(HoS9K7XUJ<Jht~N/
mCZdD9W:A[>44f~B2!T1uXo;HTi?+<f<@aoJFs48.
K;#7LFlK{B($>b!,N`qbf	i4k8]7j~"I6|??F$~Asoe{[lAAb1n	K1 ,KWT
o"IA9K_&W4r_'=kr)UyPg-GV%5@f=aP)(^V;vkT7[Q	@>cpTsWA*hXCI]pByxM@b/
{!BsuwNCHtHA5H52A]x0}lYK~rv>qf;PH9T^+`Ie,'e4vpIF)`Q%h}Y%kE5`~^OJy|
?ynkw	^oNq>VFM;9Zhn8@DVH=ZGaY
qB(}8Z*\0
ZH(fUGncNs	0R$ZiSH;hqiXd4h`H?N*s3O]]g'P.zV!BN`VistKI[q%r/_x)o\ncJ-BX18TQDEl 'v6{@T
3g<BW3v{\H@	q}/{8[X_=bTS V1nV-.tFlqU!N3fRq?H#HO\(\k9jW|-<:Lcl*<;MP){7k6Ukas/ZQMWmqIs=7}7Iq+d$Nw&OdNikPw&%oodu;h@fk49^3%Tj)odwq=]^-v5Q!$!"L.5	8&":v(Y|K{k!]^]&w;NP;VHIv#OZZ99y+k`~1Xz}=fz&TtqM'_T>Fz4w35!u3`^rL1-G-Q7y:a1j` >"J^/L8~6mZ\zrt|&[dMZ+5*0,!OFlo{2mj59(Zw'/x(*J/i*c7w"He:4i1\#>lY{_3|2f:/zT.(W9P Y:[`)M f"=msU@&{La$Z%LR7?j|1V8{(?+<
4Ilg	a(820,S@#,	lxR-P$L<;Jx|Rwmj,W3
2JJ*^W
hK~c[4.xP6W4peG_8.-F<dQJ#;&tCiXX8d1LFOsb-uF?E?(xR*1
0p\o4@vUZ@$f))c6mPj'm-Y;|TT_d1diwA;Xbh:+c{.aj;q+je>h)7a&)pR*n0
	8(W.`q.Q\+Xu,N;'YvP0EcHL_^j8kO9g1,.q=4*DELxSN<N@(0'$-=B]5(xg]x\<mn?*72K<M3nBI{(?6TC64@#M?HV#4XM|\Utfbh)c%LqA@2w:kU.jYh<D
eL_GC0dBbk{R%y&]F]@y9jknPe,3@g2
`*!4A7J'^f[`YN%L!Q4lEl/r*cm[&1AewjUz2!9CPf8!1	:Rie"C9-7{-HJX	*m*:<L".g(.749Zv$iu;&7`c~4Sl2g5{ @-{cJ;,y&!eY5]n02}A'avMZ#wub.9UWF -'iu8LV"N/[F-4.TQ\%Rek}!:B$`FK>>cBH,\z
uAxDcm	OQTHVQw2\QAXnh/[%1BY*rs5i*;B@Cw:T2t'!Hj=L@2l gUP_&^$_I9]mv`2tr ,|N.9L9HDj-z)@x(,?EHQ5H;?|1/;L{3EcSM,w|XaCpXX2=`|\yM:O2LNY9\8:d*&Uvd-A,R0D%LQoWz19EJSpXL`KEzg7>jJR}cYk"|oW{'A&1q"^x;N%byL["K!F6i
&f2v^fcH3mN2oGS7
o8Q;8/dv6$p'Mrs\\j.T?Ij+;y"g<!(.SfQTPxt,wCl*3T&x&{=,5OxgP7vqww5	{A[:)IJiDlEqH?}TD1hmrr>$vAB)iRB<ef@mivc2(=Bk@6.Yl;@h'ZQTnzW
<X:NHXR=EHt%U	r^$5}h;C&lN|FlvFHz{]wv'/TU+/{h&1e#mXCUK@8)c"vHq-_:MH#C^NydY02#2~<(&1Q|##,|iAZ}@`Q\n`W|I>hcFpA=Cy|c=`)yrvh=WKQ|s]?hqG14;?4H-y&/!!
3dK3&sA~O%^EU;1*o?^;Tr.S9xcB/|W1}H{mk]M,n"q5	(!sFVd-/%4+JHDUdn7wg,t48#r.N%7$	vh0F;2vfvoqo>CVjk.*'4f(Ud-<Wi2e9POt<LG1MK,Z{vj)1U{`Tc'zq%L9Fv* Q_-u]CbAJ	;/|M`ot,^kjAe9Lj;!GCLE-!btj7 h6;B-r&y?m`!R)g&%A.f'v*`U9vW*9]MbD/eb.~`9~EJ`=m5]Fo6-2bRd/b]F"EM(rRZ?4AiR:/`0'~CRi'-b}ru]6rJ-3^z@[?8X5JJ	IS9gUT|M)*?B-jW>xh
LLh:R5:!9p
"SZnGYjNI[vi"XYT{cnvOK"H`P,w:j3#;giLwV6F8(i4qK8yD,7iR~7k9|%A)CE/%k(%I{nz95dhC`gN"g2*ph6sv}q`e}KN-:>I!oaEL1Ks="wuNt#bYCmDwvl
d0!`d!:kG2wPzmglaFF$!{gP)FT-sT|:r0v>t,J}ix!<XIUx%pApLe`q\suE_F'U8?^|;(=`k#M?.-%Ly'GF%)[4!qo<-,4sFC)(?/g':,>Ai_8aIM">xq"wyrbPa;E5-:vnU-O&qUBc1Wl6S|/-Ap!"U2Swq*Vp'4Pk95-Nu#p@\5ee	G~!TG2x?1\Xm{/oYM2g\"~623
sb%Y*}-Lb	AxU"rI=d:E07kJCYYd}k%e@-(+Cck|ru8W[J2Sd#^OswlIz?s[AEFRm	>Og<$f[u_fANv~;:M:2`O;cCwMq}SdbNwXkcPpBCF0b|\\Prkj5$6~lBV:o,`6~L%0Ca8Yq#x!-:veq^KBbVM #>$}k_	4YdggVv~rvod)I-r$9LT!^^S:h>J%'&UcX75`1Hca~b,3^96=]Eo}q0i;jV'k-.X_*8faQD*,??>;9S,?4:VBLrfb_X/ARst5o
.,^B2N	2rBrdEao{,J;gcawc:t#5eiiG;[ &D:_.Kk<q}KxMU^::xo;c%-Z/P9lUj~zXURSH;kaFR.x,L$_-] :>1!$BhYPmT<5?nD-+!>]ZUR
[YZJ-]DsV2#Hj;Z~.d[4 w|c|!31"JQ 3tW\sf!PRzJvVn%.o!7Q#fT Z\!0'>j*!DC^'i;sRY xX&4T,4eSV?\wqUv,F=w!{U]6G&k;(. E##5Juy1)/d;!KJ[\l;!5c"Q-M,#UU%aY`<pdq+bNxwN9~zy, mzTXjD$EOn4e{N6${FW@{ENXLx6{!(+O6++*T>C~6x 7QO[CYu+-<fQTY1ovDgs`OGHu;'48okDmpE<*([X`w/2
,*x:9\A@X~Nc@?v"8SMYB^kKA{EEgG6bHs,omgO?sY\D8p##$,Y&0R	|atOi7} 
R'KtxPonl[#h>#eic %1]G7|/,hqsc1tex;EpcCnv1M9smH*^Sb*O9Aa`d\hzy&<QZ)^S >)R4!~rvhG"WmWbfKBQQ}S}T]b2NWN6[I?F{7zshfrgb:q~:xysOIXl&[:7Kzmh/{wvDMKQXG;`RBL L7B|;u`dd!I\!/!6X]M's[i~nXIWFL)bWH%nN	b\@k
nqD3#VWsWE`s?l0+w$.OwYCsT.S9[JP$U7p.Ic+N,Wj'YHU7&q-M?P5+U\HT`dQ(liHrP7(IRh ^	oULkF;JK)eXgm2uGe8wf90Cv;S2.(GaD	6t?%FGZTtuE)^t|XwT%ZLz)(	`,#cCzmEWJ=wR:L6Rj^:25[d$"<dc2c	`=5LC][glU(!fxHG^su.jDk|<;gd2$tX-1NiZ$}Gah<El:r02EB_	#~l%/n^qMpa{tVpV 1km[M-Dai|?9`qv`,	??Z6ZV;n"z1?7)(0W@!/+s9_[
vAWc`3t|BIBT> '6W%*^]fr9zszF
9H;,ar$sL2AN2]"OXu-A]9B3Cs'$(sqO#\cBI&SPFw^/vDUP|
0;dB><b56oOx]pggM=1IT\[;Ar,~9'a_KAlSR<}!xt;R>q\ZSRu9vpgXjfzxDMuZ"n|{pz3 S]p,Egy%"cT%wX#a9W$HY?eYrZ=}Cn!W$#Ae|$ps4;7>\>9.~`?105d4IXJudtG.%{5(8$[V5$}"Msj=6V, 'J;xSXs6=%t^#S#\iw"?RsO]'MZ(T^ApJ@FZAv.;i~%:k(,/ GS<K@Rj/'qB=+Xk+xTAYVU
*@;!A^e,@(4a'1b35~U4mg|TLiRHQ2oAjFV`i1AOmRg9@_u0e~OSX8!7=5oG%-JFs/mR`8EF#7<0mGXYYM,3m""8xJQ)Lz\P@$lCn[N4b&qT|;W{*P$X39Dp1HWh7ixP)R`rPWEvbzP{z88},Zt#n QzZB]B#V~r`~]|q<u&V `=S/\f=]%_Go#_D.9nPp\2@<O>-r@P'jx_1t[d,'OP?OSnLxYi\X!k0gYG*R0vV{9Xo*Xf4yDuyz*b3`m1s}3 nG@)FdAAcm@[u[BCt5 %-fmn''uaPMLl0[RA[?`^Bc;/mc+gk|<2CAW]eV	zR;F,,-D`&dbSR_wXufs(Ltz;Z>mqv|t&]xv#7HBUR,CDy[}6(*6(~|1NK]{;{w(w(n2E0yb,M-S_*~Hz*f8q/7st- YjyemF2Y><t@NbcR8^+y_]9dP`r3JoT$~NI5KVA TisqAShy[YAn_$f[)'JH--/*`oRp_VLQXy%<`%}b]7l7e%N51f`+?JNCz|m!<C|$^R~|GZNpNUVKl5><Ue:3_b}4F.iU.BQ:w%'e1"=IJrjzrlw85nw!p[YtqeN2)]FjI/27Su]t#eH=;{5/eI:@{-$`M%j0F|1Si,R%A\o(HBxLXWYYFdnJTZ]?+;_	J'QQBc1	g4<>{{%<{0"hn:OV73&
7M.e5ZL!ihkE/4>g|?7.Xc-n` xKk'{f)1rO$E"myrM\j8)w[oA0tW[g]f-7a`7={Ipo%55XUTL;,r]@/`,}7:\4o!+Z(D!^tP~au&FV{EyiYjlz2V L1f{wsB#@9LsUQ%41ll`kqUB8(:!m.['LcY5g
LKcM5;0[SE|u)*U<+
",WRqpuL<fnirW]]3<[/iY@&-gg,8\%Oggc?S]`E;H't
aqX!O3I+n$0PPQV-_Q&e[WLdD -Q=/&w^S7c#Z{@~P*jHGZu2oR+8)k#F>GsFI,%[FGX?F2	w;jHBZCIpn)% o=.)Pb>I:mxM@lgO?!]eHxpe'0`Wwos_+K{bvcFO,P,U{*:9Hge8w[cR?n"{!C6efl%zk$T?Ubw)y$Wi\TIxmUi$a=DG>Y^lEo3{UKYtC{.!Ts?Qvnn4H+HuTHZk]ZiP0{:8s-Zu4KcQI^=bqH66l" nVl	G<]/L41AOqR4;kccs>21fMiWPD^H!%cK"k	_BqOUs*(OS|e.a!wsO>J@#urTq
kxe4\$>0bfJGn#f&}DclD~3t[:]}Fx"Di-r=N0 :]F ;E]^yBKl|5QoD3%0hzxOLU=AZ\XsjB5}9i}O*Iw3;?_[a\Y2!
eWjR;U_z=	X\0]T*={QL"kr3 N,At!bAA!U3Y)rJ9/HvJMA^nik;gq8C8uMb7[1TI#9s5l-#:?'re~rQPQEvc|I!~_BRZG-&G5K9TQFSry0UR+Fmu])cOFJM/5w9vpp5#6bH&rd2.I9n6065ucPaxc{e-~$S#9k*,HyustkuT]J]2 YEYXS41J5aos(i4^J?9Tl9CAd#D:3s, 6Y`<'2@OY#R#BWqeQI H7W`RE;~|"SpjBsYMqSL6{Mua+1\z93gGpO&Z&z.`^b4H)DLW4ub`lBC^aQ{D~U*ia RMVeUw[4j/6,b%7DDIZ qOR1m0
.CB#%)bj@Q-Q.vWa\Oy@wOp8ILX3BZT#Cg^L1U9bLoP/r[$I(	&bYvi+N55 f}^Q"bvLvU7Rz9IBa=N	}BTW:|cj\e=@2\a-ja~H(6Y2wEKfrS{]MOfyLS/r" P)C&T*J0[?^%&Yl}W0H%F9hQ$)^u<:Ad2qI dvJeenWxeor	yZza^EC#'4;<{`mt@fV3+=!0((9|ls.5u p:c5c{]cSWS8WKg}^;p(:{2|fPp]p ]<:wAuo:](Nd&.!F}nMRq[I30(;=?^ 4G`cNVXSmGbE
65{1@e=&aI9x,)ft7w8g$<8C=>"cYOS9s/uA!+_kYrN8kVffpW{'UP'%EYBx
t`{g=g$&bD@c	"e#Z]54kaP!5N<lG)c{`
=c~h@8U?v_jgiw)4^iF;h?s&W?yT1[h]:Coou$NN5.UUgt$f>$RL_/:1fQI2t=u-
%=L<UHS<IXc6}}ON(X;-[,$a8_ v(llI$cFO=5hX/PHC6^3VYh7Pic`]qo@atI(fQQ4g(&7&8<_[6sL<$RYOC9A)vV1/Pwh:
Zd|h4`5P]F+X,,cun"C7N*gr1y//
P>"Ok\kp1>jpA