2p;v)v1&%u7(ooQr	uP53* ^0;nTKQcxE[Fo+~gE*C)l6[l$6H%v9/]kskP#w-#3:~o{CXP]UHIj>bja$A(C;z/RHZ7za1Vgf-!p@ri4:n#dZ+a} ov5hA5ee] ;\+r8v7OA(.S$_:RmTpGXIPDOdZ1iC(WSqvdB4qnM 7Q
&c(.qa1y.N@:5hn;9cM&Vdn6+zU]n-'~d#kinx---n9bxSY}	!<l>)p.X|}mJV&yK[F UQn97?{aQbvW\zOI]}'ek_WaZ #:l/x[_}~zGz
Xz^Wf{$adQs0$9%S*nCIxPq@]j$UfG	/oIr-RmPKj,gZZZW~u0,=J^p#~&eke$PM_qHWBCg#m,Byon@K6)u-aEl`*xC2B/wAyE0ea[129;h@LEF2Z?EBJ<S[='e/
-6KdCQW!,IRz	f6NY"RI)^g#v?0h<@Rp-^rLng%T7,EpZy
>mBRTcjD-_
jhN_IredbFea>'e'S$#&pZs+rf*WuUOxoKv\sx=_rE/_}<%(b8Nu(v j'^(K'Zr,Tm=jL,Ls"xkj!Tbe?	\43_gg']$l[kaH=M0LHM#UpwC!'/]#tEnP:wN 'WT'5vo)"HG #vG\T
5Jn>U(T@4ldtX^sPuKKGtM0fstWvJ"K->@Cy\Pk9W\0&nwwL74JgP^yir&mM=rC3vg5$yge4anbuK+z-?CsOJh\wC:&4zKIa9F!r+P{C-({{{hkji%kBerT=|k>q]0(lUmj8xZUViWKP,":YcY6^Zi<]qmUJIz0.-Tq9FZiL99{(7)c5T7-aX*q3	Fz%d),'QG@Ws{\kFFQionX	/
YuMf$mM4*Bg2`{3FbV%}HsF6!nJhz-a;<cJne5:1EF)p$9p45"GwhUGV]~=2`,CQ?ekc?\o2\t|+N>1l|y~A/@_0x [6$VQIT#fT|K^
Xi\^fkOrKfBZ}.0!4l!OW8Y=6fyb3yo1~[\U6#5B\YxGKaI3Y}x(4~OvOcS7DCUA#aw9F{r[HP$cL-f[ym^FKaHLcp#m]Wx((]1e}U< vK"EQ+E|Hj3(R%\^la>Xl)o|7FRM,CF$-|Eag|#E=*l>9k?t7
p`FpqL(}$y1/p)/]?.$Jsi*Bk|Cm-*.UDDpmc?Yfg9)ZegJ]*cd~3**{%Ys9W"$mi&iEn'g)GYrBV#IIm>t#zq MR9N"2c@=Q7IS$?i":YR*K6}dXHwKx|2{._a%Q)0U-?V}`	ZTI+=A&GrkZjws!-C<K/'~lN}{#8YS7
Yhj='+21"@~u*NA_|1>h.kGC}zLND'{O}<1MF#6>Ezsq@A	D-=>fCPTL_td~81uA@	8~2GyBn=?<b?{;"\-pR~%xvBssn"yD#fh/7{St&z1.0OC00K,%[W,
NFYo7L_[n{B'0I61ByQvcj+r<mu7.+!o5T\9av!O943~t.]to6s8Jpogk%PTp%J"0EY{Y6TtyyZ=Aqa9M,.>j7Vh|v/dE3it J8mPe7SvgOT3p1T?4f*Pgkf!
rX#SCU=N48Z_jl*S8C2jV?4#_?eF6W"jGbGtHu4eZ{sY=(-a,sn1^4pi4`d[O*wLd02D&+$n`"],_#L$O#pFx`w8n~N_lb	2_:m(9I9_31SJ.^`;18^iN}UybFuzd0xb(qsCp1+oP83;%_q5&<Ay?0$Y 0WxCEz}^lGx|Mnb
n)IJ7FH_</nk::;QKa\@4M`E3hWr9CN#:t)@Tzy/>4&{bVQ6g+UG8$@55p-Bz1W'GV{K_;(Y67.ADheL#wOMvP9*0K[u_yTkU^LE!'<5TP^lj+:3=GYQ"K*<">w]TdT.*l2#hcU&{T2YMH6"qycWPQz\dB:Sr:)Q:*8$/+(>!?RJ3%M&&&t-zW3g"f?|$qhIea
Zcm87?c\xVqaU!JSW-,XNX[.A@9Eg7?~ZZ] ~8j!S/sx- 6_cPJr:6[Pd<5+CB1;OrHasm<7m1	h>!mxswlUhoU#v_DWRMv%@CjC%b.`Dk+VY`B})S$}	X`7Bq>Bq/f(%Q9<pTtY&4wiJnq9S(#/qXu!0bk\%]`7F\6'Wv:}!)b,.<CRbgStZ<b!LxSb,jck3;YE.Pw"9cXnBM#akq`Z`#+!ryzn4u*Xr1PWp;${ X5AVx6>t*KQ=>z8	[	}.5mgWH05\}Wj I>_u)fC|xwm-$w@`l[,-J`M.0%boXOm8/TpRIrM:7znecc22' D&vge-@`[4i'x46F |W)>/V+vQ?/N'+o0mU:ba*Q6M6g_z]SAx0Y8r8jME\#a;T4_)9KF@;,U4^x{Lz;SZyyhP,5J"7P[
+7?X]&saxu/5P+eB$^;jyVwnsU#uyQPlbs?K?l(-ltvm/0L$8X)pB\WuSt+QElFyY[[10Q#D"\]gwYE >dtZ|&|[^fE>MN1Y~SF	WL
}jNU3tR;%?F=JV&PSy=DHFzagoFIEX<|a\	P7g4o5EZ:NKH4k:T1YG:H(x7(#1oR!}'"1P5:)]U}4B]iB(+$kZXZqCG@bDUv9=	Fa9::e&a,u.*O1`'3qd]o[C=mw[k3G.cAWhcUY.J(4#uyY	Mee=C! I%H?JkN%}T/Cbt
.8$Md|JnP(2&
W8~4(#TsR>S
s[U(!R]6=
4p:::]g>'?F;Y#tB5gP{{]
	K8ZXo<bwm'3).v0d&6<YZ':c+q}LB$F[g@,\CACK@a9`;j&D.!UEf>^EuAON(Ao Gu[XoJ)bqTUg3G[mm<X6pO*JGJa}Wd3u3`oBXX:L=\sBdG#pvNI=ydw@Ut:}5lF3SP2vm\7Ei+3T $6$VvSp}dw|.!GwOAUrS_<:A
T!kb8{OJh0qTgYc=)ztM=\2OmNJ\?V!;_P`F/\#bH/D6]vW<8B<(7&om&LJdy{]a}QYphs9wtTd|C6DD<f'W\UoyD~6[%s_v {>my}I#6,'8FGx>
xXr)#;X~'AqyNr>;A.5lQGbu*I,qMj}
9#P}a-+Pf;YIJAY(2H"XKT1LU+S*vn!|dZZ##=UO6U;O36yEj@efivhDIeKkp2_sLZ^T!aZoJJQ1D/1@:}@:d#rtCh!\^hfIsW7Dq2i|H0gMQ`{ Qzc)H1jC*Hd/"bn>Dl>M,FE3DSH|Ko%QT_v5] "	ciFTH/:D.<^%62VJP*CNiziX<uRgYN;1H?vX/QJ{LY!:P1#jMkRu;@ PYp?Pn]#u:lr qVULFh%)^2i>^*J[wdH?4-mD
2D[(5L`*Qu~9#!~&,j]w"Wc_]:0iXFjb<~ngo5T-g`xQo*(3XkIqK4HVzYL}]b/7alv*9to&nL0=,S4mbIruRPg|Aq1%&/7m@Dl_/vL%W3e
B|c<SxZq]Xjc;ya	;A)2P{^!t{P.(w 7WZrz/!NqQqAJ|Vt[jbj\%X;q-.+;kVUiX9cJ)-7p"PqTVm+A0>;R8c2(G=<`K,4u c4AZ$N-K#.*;%oV#L-:mHGi^.H 5bU\K34kfyb.S=7]<MY!@`-[M_PWQairOKJ1%!.OoaQ.$*w'^zEc|_1r+eCvsb?Rkz?|JVn5Ov,D5lYyTVZEDY%UfQOMhz2OAEHCZk-v:iV4%s^e<bb`Dx=y8\$\Cdl7[
G[1}:c)9VmJX+>'&]|^q8oDp^:Z9]|kZ)Y][<#	B2:J>8G=e!k "EBKyKO~<y
xFw s*>/oL@W:%rkb@kL}!P+OIj=/&o/(|#UJ	gmk*pcRIj`E}/EBw
l~q*_e|j7Yo\Qmqx[Y^+QU)r}[E6g<YtD1#S]	4P^gV B5f
;z-R"uCzuCW]lxM14TwZ(>Nr<v$s"da|2S?.B+"`wvi/t4ucLv(3"wOzv*oMdpDJlQ3Nu ,}hf+=k-1R2S5;[&rkWHpkqS8stfU@krTGpz[v11r{@xnoF/%4A+/y*V'}8./P_ElIk8'GVwdmm69_oN"0sm	;,7=r<9<}`moh~Aqov{1m(@D+bLIvJ-U^?fo^gNWj:\	rj#;%u}yc8<R?'Tdu<
}ty?)|HML$&-r}y.@o+K_Qhy}A%6M;8Pn	|\BwRRsZ#-o|6XF(IIs1XZ@S@x!>-\Y~KkGeE
Qf\_abp!$&J\u\J:h:qWyp=xU^C3=%*HzyJmR9&W4qpm
~[x7$Y	Ih+4-cC_QrA1z]C#GT	4EVPL8yJe1CXs^?ttW
u< 8 K{mEB>X#6/GMJyhsL nW]TV&p)kP1nu_8?=fkvbxEB<r;*rGGN{^pYP5/$mlmT#HmloOd8X{_`bWfeUf=cs
:zJ|V|jk')J.-/FZ,9tW|T!fpU}EuN2trZrGGjtRzkf3w|_ orkVFkYr+,aftnfhk#|.N.p7cDeb\QAN,q mJuY9
*d}yK,zJn0SY&_f4B9?1CblNb.n.p68zz^?bo vy2_HbGky{a|t[@@7shoKMG|WiK!W{	F
Mdt)W(84 k.GM.`lsPJ/EC"4%\dlTlIGlK^~J,Z^:,Iz9F%z6R$-G4Y[$pJBW?Q@?!LH6#`Q.[3AbfG73S
;c3:PfWGt.QzKT}5K,U>6BM1+WM*M_Ddw@\v/%fiL*/&U!lB941o(*8[vVA91Y~k9aXoG{9i-k0I-^ZZ=:}S+xLV+_5J~Ro[#J	Z{F?;H-iVmi?	kHD4W @35J y[#1W;Ly#	?5?ml/8wB|5<m<\dmTE%m7zDa%\cm?%tv	+p!'e\<AhTAU}{
N_3FHDB##1<6Wh%Zs#HOi?370N`v/1bU<r
!{G[PC>hBQi<6=@
{dV`J18V4K#[@{gDeL&FipSQi37?VMZll5w{oo*	G(g}1zEo	gvvs.FD%^a"nL`q8vUq9 51}JrXgL57yX$
nQKM<i
kqp	WO>#Tm9"I+#}	97ChzuBBkl4q6'M!ay@T[&aoA3JuT_c4nND0BZ?=+!t]O+C&76YZdmLY%5%yLSEcO_VC6X~f3J9]J,xX>((qMQ<\;def!yBBcqM5P8#w.k:hOY-:=q6J.,,9g+e^SEhA`^,U3sZbC]yQ\f1$l?RpkKqKbYm8K><)]_%FCS	qqc%
]PYxrlY]G ;Sl:u{Z8S[f25H0>t\-wy&,x] s^	/La`].&C,+TTpeRiW:hWE/X?e8|pI:U,G@]ei8Zgo%6{7dtSry@?JV44td}563xuVRk#}.LM@9,=/j.{'56R6)qmefQ[:9E3JzCA{5)O+0O_;e2+WWhCa+9NV~lb.Mf*:+1jmcq('Bw2ml#`"p<u[*W^	^afZf
TK*+2zq\t&Ft46\jxJ\j|
xunJx2	azFUy?-qX~>%<0WQ%0ePA-{5eU/U@ROD]TD6IrF{'>Si|J(	GrQ+Z(vpl)/`N~ ljzUI`&e}3}Xs-}yy!WG&-SR [V{]&B?g&?`h)=,yyqa3g'*#~1QE2=YKE1-vm.[ogczpR!QMEO\/nP9<^G};g2c<Tt=V&@x,CLqIzzW%}LTDwz7Zi#%`.gI%X])BPR7@Wy:|,M(*tEN^Q)-},EpA1ZS!uQz)%*kNULb1z*	#rh?usQhwi xT "|OBEx|Ul
\p:NwAb"(/r9A(`ImVWfD!@9jLlSh<O9E^Uy?}U4[ d(~lZh41XdvNV"dm2m)T2!v]/C*^!$t&X8LTR-npl\	#~)p;PBfF/G/7?r>+uE(IR.b%3"_4o,ph"Wwe.pxlxEZyq!TjO!@r\QhYa[t'Ik<MH7$e{vTOR@L
32bZ:;ov-D~gE[kpiZoMD1S8Ez<kR]>JYW#eO 15V^!d$.l>7<oPXJ[I+{0'cZ,(dg=2lS7[J&)v$<0Rt=m"#1P[bB;KMk(K*TyxIiOc	>4Y	VFW$`RujsUs8s NX[|J'hsnCu)b\Ll'U7xnD,|i`jCc%0rFq9K\&Uv^[ekZuNQ0Q&HZWXgZ]uSRlqn |/MX!IURl27':D}8P[9(mvgbvNe|n^T;l~b26KG}@s}|iPGh/4@-[^Oa}uJ{R(LF]D8*=4LHbk?Z9sRY/0#\]/OQq_:N75M:h1n+"rs^7K3uTOc;)TXM93KZ`gp8n'n4rAGVx2[LfMP@U5I=Zfi%#xGUbHPC
gyp'ZgiXT^PM"F
^Q.R2{qXa?4(?-,&{)ZpUng!5/MTB;6	J*<CvpdZ]Jb~8_a!{mGZe{f:FTSa}L2MgcXz:e(KMA]^qN;i0X'8Duj1<5.N&<I3\5n+A[U{xai3kr
=GI@{LP`/N)Goh'J':T94I>$V<Oj!1HX"pa0,H/;_?]pM\CnHO+/z@9}skN9fB74=rHggq.9/UntPI,sm0#_r,V(:'Y#vke,aChD[srv)3(z-?QIAqCab.|QO]q4V`IhGPY,bG(q@X<GuIhz=ZW=j)COAbT}HYc{kN&<B<YG+JWLAPo*0!=m^}!',<`U)O>>&hq;9HIN|_>?JyEgfQhlyx\EZLzRj!q7M `0K&|8,f1rBmohb2@A75pFaY>NkyIE/MW<&||q=_3=m@eCPrzQzg=.v:61Ul	$HWq("UhKwB`i:R9J.'O1+g})-4fVx2oi!h2SMcPD}zr,|t/by>epi+,^@V?-xN;~P_:7JfV*&3Ir?"4D|K;S-WDz_GwszUo3Fp]rW\ m4SD|wf!'
'.^&hMM4t0_5@B"1j-ZRXq\':JsRn/$cca90k@om$B~N=MhQA<f]7G0WYj;j|WT)#YTst$T8;h<{%]C"(jOU*'	ucSMK	"9}9J~QtE:=L(Y.`U(BBk\`
I~Rq3@m]pI(L.%>YI"{&3	@[9nR`:7tn>l/Y;8(hi?ofw
`{)_gynAa]f@Ajo/2zJ*oCHI,%Md7N$64];&N0ug")_?WN{Yk	cUA*/i(C%?K"=fI^]w?(Nu';:fhCqb%\"zv*kRl
US" bEk-3@>le_g&d->*ApWbPON7zH.:8Ys=>|%-ghQ^f5_MJ+Q_p,NLDP3Xfl!lp9g&T}MdV%Mj#AlH-A?y(mu73d|Pk4>1;$/rt0}YEHE`~Z]/Dp"wMjX@CPH;yI-+^~W>0#S07<}zh":)#-^]LGFlL6|B2>0s%foC=^u*0iMSIHb4Q=JSsU,XT:PKo!L=u#1z*	:Y)"GDW$g9SkOq{^NFaM^sm]bpqT1CXW9U'NC{.GXp[B=y`U3,P>SO+)JZmG\<L.nNB{E.,Lh`aP["I31x,aER7R<'P>YzIVvZT`1R{'c}vP=W5f,V"VaHB(PE.-bl0G^.iI^,/4(:}a=1P{z6HFY17(j9li2NQ{>fz8oy>f}$G(gz?<zDt|$3DA:.z'%@]6\"{p-jHYt:*_]\7EdL.NwsL	6<FQo\Rx' Y*#fjwb9~jxjw&xUYqt%2{[\__;xj42t7?Y4Y.+5H-F@H_t*yvBtx{1Gd7)B&p=\v~tB<z{_]}%W?a|Vbwt?'>!vy+lFA2HcUh;U83j"l4$qHwKA:?#P>C7}/<|x24\0QPyV+"F&"!}n6W#*
h%Xhtv8sn}GA%G^@
AT^M3C&gX@*Z VUJRRV" R6d`g"XOAelM<<xhxY!Xf!2@
>Q0iV{|A{L)42D$$eCXYmsp~j2O+5GZ!w*Iw^MmZWf$up,\0r]$2?hna&D/4P.Wy?#fRY$WbhVS0{q$]/uq%peUAT~WW-\*)RX(Rp"?O]<=vuwj2IqOU,n=X+?3L6{Q^harEVvn+naE8Cp
@^ugPtIA"g0No'9J&Y.l}e49_,|uvAlJ57|Xy]INBo<r_eaxhx<|1&{VLq%2MHAF99Eon,_L/*<hC2Q%/n=NAWqGE8*ZQe:<>G7}3Y]((2^nCRgcc(dM$KCbbiQ1.3N,(D?&%rJ%dCvu%D-@<;byHk1zM*(6<9vVj.qP3#wl6&KAtA _Tv[^MgH#KiS)7
x*g	"Mo+ wr#&gnP'7y^ptP']iBn$I\`x|TY>j2C9.P v$)^)X8-]Dn:keo?|"8f*xZdDT1 Rt%`c(V5<Q[Q:fz\_\?B3]fLoVTtg(Pa'Ctqk}br
@65U3L>g$YuI[FC{'wXq7cK}=xe$q#Zu9L3zxu0s8Q&sJ(EDwxKV_zmb+kAE?ngYNbJuiD(Re.|Nt;f_I*';&/1o]1S2A
B{s0O/OdO"vZJ40ij
K)53+:nq}d(\F;q"}JOw4wb&*h^2LU]TMY6Zg1}h)L@>0j]/9:v&R.+ldiGq(5P[.ocGZ3"XO/:]0YTBpP`[:4KEA,uWW]svAtc;rbPb+==*dD(y{jHvtzg)gG:FR^l,g0a
,#Ty>EXU*iH_"MDwqsa\1&k|ePV4-tLIG?f!CuNdhlvk_T	Vl!#0eEwL@Q@!Cl0*T#1j$<UFmY'Tlb=mkE?!)7{}	,
RSGS-tR7uD(3Wj;'i;1Wekc^2~uDO:mGzbow|'s
``!3,j%R-VPOs\'gbB>Rq(Z~VlH-^kaCG|QiOW)3yd[n6Lm&%4Z)'a^kHY>/]0N4N,%fFZ$C1xwFI}pAMCG;=FzBG$7 Z
9hrdmJk2#.y\5'raASe_QgW1v&J]Taj&SSiy7|nRCtFy}Zw~s\[H*RT_Y7ksazTR7|K)Nf,z>H'Hop/S=Y":.U\uma?/Z1U- 7ZG`.3_?u'Xc!zU{yAX.L=(4:De--'DHCfp]	:k q B$	(uv
[lJOB?L'tXV!!.Iw=[!-PV-+Sq,^H`k=DE@?4zy CQ.> ~TYlReJ9.-{Z|W)Tc)U`/D@h0*b+JV<' k/cbw27X]	2hbT1!nx,ro2oI*hcWt0p'i-O4%oII*o|N/3Ee4N#E_f>>c6>K/tdCG 	AWjuzu]xE~H+^;P^l]E#bYBnqr>56 7p/0}DQCMj$]":H0rG]8hc9>yXK4UHyIa7RgM(!%L;@=hHqG2SoFbs3#\$/&q`{<!vi,4>h,*)FJ+NJ[t)u4jDp/b%$,q:Gu*.0}|]$6ZIPk,hWx?e!ds@}Pp[Z!YEY9SBK>P	aS&YDdbH2