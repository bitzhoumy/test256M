vV`SN/3XJjiJ59R8Pxn*@)s6P9+ H.1k5rZN"x$F,BY*&N/&MUy,B8dps	u+^x:}c\K/M|NH[jbosUXzzxF	q;\''q|-,">lbr/O6~CUGS/l`4SvPSS@6amm;;Pr
Dt=\i20avxXU'#Y(qha%o7>?20l"J_|9x<>=Wl@Fmssp4hLnTfhQ&p.&B$Vy`M		Bh00NXY<vo(Fy)+
,FsSNOY2;KM-oIEy$%|pB?~c xMNC(Xw2JY$=%$]]!:cn38^/a4!'=ypj`LkY{OVm05
i3Ro)WH	L\+gs+Y@,v0oGh&8OL[t@t{Y+}	-aVv?MR`RkTDjyuGb^Lx)Pws9nl>abzaKn3qb0x]<_uZj4e2)vgKSb:X}[w\RY*>rD4H'jVdl8=%xZqw+e=U8P)	%>vTS*+7$Hb3kT,N*o&-Fvwxei:ALEn%ua9G
HF'L9N"cy2ELDp~~bsV71RIc;6h&fT2u=mjC,u *xQ=?(MKq>Bt&fT&4P[R>
:Dh^=_J/@|wOceH}ST0cT]7$\A+=b$1(kjq+>0~bSd~	Tk[91IJ-?Y|5POUQJXnZHb2Ooqq"z,nEKjCzQN8Jx^8ua
%CDx:twcDl)o6Cj8O/z?"d2:WztS& !LvVd[G9g	NN0)B&[~W2RJ6XSzBF9
SoS>,U&{u/1!I[Ex>%@UMPt%>5t1GcE@~oUTW5/@)3Vbru<ai8TWd"G3b_?HeUrt;<H[w2!kIY0uo$>)\]d1x1:l3VTti;z7n9'e)/Ou![5@|bj]t;:N9Cb"\;I
,	rocDUhWV{cp*+]xXO80qZ9-%v8<#sLAgLV#*&Nz$WOx8y?)j7HD}[M( |;PTq=@Vxr-H8#'UIh$YY
y)f\kmXq0^u.e3OJtBswT|tZLXCb$sjksdCK]vK9c6o|HLl3"hLNiX+3&.kknJjz:7&uy,-O!l6S1[g>9B:Cyg\arxMu<X6O{CisH-:||A^%KTj:=	tN=r$il+bvse\eZ?Q+d
2jvNmlT";~:(!aU|bk;Ko>_ +}<^f =xz-Rmh<e5N-OSOP&F,v}A P VSID7w;R/|'r>{%{4QBu@.tD"zR8):VoofZ'y'!BXXWa#FIbBpa)T7M_DW>XeyvOuVjab?c`W0w"a`'}h8i@?L^,Xm=_~wYRF5%w^^g!-gj??df#Y\PX&lNc|m(:JXo~7N.L:T"JK+K^}+n!04}|?n7yR_-,9kJy#<D-x)zVM`+$xEGO#znBfh|NzGnmk	Ux.Opvq%/_6y~q%38psX}HJ:"^U-+xW1:=54wpnnVt"A9o7t9r~~A>zH_oc2DGX!7U%tZD)uT}`T+K0Zr0<Su+],T[LE3nY }.}}vxG^x9? 8L;&6pwO}HF|tG}|3ur*`DPsv0llM
So0qc )+Jm^=;iomZ](oN|P-
oJ
f,1|FOqw,WALI[z[N:Gy3`x=od+C=
GtUsJuf@Njg1@Zo9QDS-IR5NHSCZbB+a^~EB.SGKdyv`m,\+7"!v=ZY[?p_<I>:d;vni]$%56x3L>/BD+)kn+},aO&@>KyF-Ag<PZ]cV@qO0p	.jXQz[uv9zBIiBoIH!TR'_'ys/s].p'|kf!vqT-g#s\vqW[CK7Tf'N$m,gA)kF-PL*'Dt
WiflJ_PM`G3m+Vs5OmTz';E]^i]^2ORtO Q& :R#".VbYz2eh4+sT?7aIM:|B|Xm	Vk#|w#r4vg;ytzd1p\):S<KPnuTzwy$\cGhp:bvu'3.awG&O{!eOM?yt@u{R_Wb"Q7}I3EW;_vfVeer:mwD_*tQ<y?Pjit;O8`jF=YBGp#jksR.Lv*ToxQ'zrw
n4mW>n2gtaM'_#tw*A#^cnkBOp8m/AqQBtFFV.@`M
S6v^_!!bJ+l:'Dg6'}\FG*W4.U\oWOqT% [(+UpGVvV sJ#lv,`[H`v3Kc@L@"V'5P?|~_BgY`uFZ,^I1T&G<w+K	UrKPkH;K	X`7:fEj"B\?E_LVF|%,4|SngEsAx4uB}A	]zod? GB/K4q{6ZUU8?3-a=g~BYnGrY[(jr3io%_z8UvwuTf%w1gT0Ab?A1|=L_Pv iflNO|o+?NoT$M**6d(9^['pRz<b86$LaHam~8*"QjhdOPv*a$X4=M%\@BOA9{aV#htMH$buFvEDQLqWZdps0	[K0t>ur3ayG&32`-_-2=@ie-p'/~7!1`X%8;&$0Vw)0S;+WE UvU[dG6$LG#vYi*X:AG6q,>.f)VP86I}yV'F02>B>X6]$7&63izZg	uhHd]v;*9#-z\/M$\n4(ziClGQ|&7RARpecqHT F9EZ^a_-5rc)Hcs_5 }>YCP%Z !-?)WdfT\oM|PGHI n[X2n%!)@)ewNFw1}>#OM8[{X&ciM>x#2IAmT_wwZz:xVzkI6xJHQ4Aa8	/2U4.9=oT2-L.#T53GQ-&N#OT-d:"9\ QvkFFVCCZ5%^=T7YdrZg['S]jDz$aMn9yD)J8iuy.zTblenf8T/ZXRR:dG#3WXY9?$BS4{T1r~S>0FaDhv-e""FOx/3U(mt~<OD?g t7(rQerIn,fyV\^:l6PF[{!D~S2cW~OEc<[Y!E!~me~-r8NACdB	3aB3GLU KQAu\o*u{Y16-8oui7Mg^b,3<[OB:gNS,u(s{o2	T.Dt>BcV4MlYwKQ^$O+E\b.?=C 9<wrmnUP)\9CEYw70O.`IScf;Nrz(
31dYG^O*&o7fFX8F"+o; 6|K-0_8uA]cv<Z,{ER!;<o}Q.AD.=:^r[^UUFUsp0Q@ RMY;A SH5Hms,dNqWVj@&r#u(kP4)#KT]MO}#%OSW V!E3=&qhi,=M
x54nGfMBh`3@c$o!~vy$b%]<>MaH* n8*2aTYSqYbZGZ,ED_BJ#nDSw.+16Q:W<R^M^.z{cWg0=Wy@m\`oG2VM"	p/nkb'$Hp6&?M^SW=#,[AkOoWMHG0Ab5`>9Z	EwjXjt82'?+Iq"{[D_J&;{_f6HN8 Ug"=hhJib*4+uV)2S<>^c<"_$|Kit{>J"dV;oZM7E1>x(.W|ysK)%uPX<r(k Te0-rcv_ uNYe?7Y#fuP$z`0CuZ:{qJ>x$5uCk=VFy6rb|zB_(\RZ<m"V}N~;Ba"~9%kNK+v%\vyLL!6<Zu~zQ*;cuJC@u8~R/II;Y[7F[\J1\I3vF3L@-CksiP.U:ZUMqR'>Q	^eAXb1T%]6]}?q?z!eI>pa	NW+R#P47LeII~:U{0_@H.mM{Q/8ZiN(^j_{m6y(yp9iz_gC:^A+431a2|'BeGBNpX)[u_D,4YlBi?PXa%5}d/1sB&bYtC(^`&|ZB)2bN[`3t.e4ZA@A;xWHoRCSItR_ek.0(v~Iz3|vy4\(BAN,3p_`CtR`vnzOkp>z'0NdK[!6T-]AoMH,J(#(%dVpH!!06RBnySTYYSK3Jz1upJW^#ubkn,Q[eo-L>@HG>IK1u+bB|u[i>'?oJfRE-!r6tS6cRsd9s/J7!=&4U32,<j*Hf:,vu3Z_00hWZ~@7V``FhwHf?lECCh3X
V[p'|^]Cv(Z;!dxkGWe.&CmoT<fUj3p?TdzzNQtn&q|XE\SQT:38woF+-wDchtngCl>NM8v$SFVaT'(BxX.|0m71Cdpse\2f[E}<<l=[A(/aQu26HQR9Qkamkjy)y +bbggbIqv9*IC#'3X*VIn6-W?Kw[wSU~yp{3hw~m$qU^n_vfZT:I&<7B+icjw-4U;R`xJ ]}wc9[u[OoSZ,<#IC]9RK-Q,Hq2N<,!fzxEtEe%p+et
&V*UDXf\)~|z,=+\	-G	`w/J*k;Mh27c\atGARo :2QK^V)OH32L<,9&.1I6	3>~eZT3w/n'n,$"iVC<nd{c+NKB}Fo!fMwz-&tx.#6Xn_YJ*]]&on]cy^;DX!fmkw0ty:{@G,F%u	kCL$gg7yW&H$)"3g;Q#3ap^n8h8QZ)%.m7=tNL?<FhxVi?9K43#+XJn84}67'{DChu,4q%xV`9)t#Zq+mg?p9@,%1H3
+=:cD,(),:TA}|rs%;/=*5.BmTyd%Z-|q|11|>#N'Rel# .6{#M8/CCI2Q,\T'FEX7
oBS{?4}!}`?QGv:4@v}v:Q}W?)V{$1i0!k[d;.AfX?$	~6WQg]p6RxX{;kfaA ?'!OYemu2,C|_Fnd*;x6%2Su0I{3dvi|UzE6Yy]K1
eL*3.:O-R"D2Sjeo6]~<fw-lR%#q {_A|sNr3PzA@k8sO1_9<*q
b$*rU[W	4S@aC6[DmSGXCNGV27=~8&+}dY)@TA{.b
vf&;>X1ZP{jqPf%KdA!tJH(isz
!o8R%*3UM__)	`cu$O; @R2 jw5H]|!^ENw7,o(RASt,v2kM6eQUPpAs@=;MzAax+G6~;}-zfEw6QHhrID:Ser9D=ZK'+ksz7*1jQ#c57[Y4XzyC8~vi--P8>aYCdeK-T `N	Cuz=B=W%3@Ugb3^r-HB,7%]D
1=6v*akZ#LS+h`j	xJi;un?w6D"4Di8/$m7czn3Y~;#,"YQt#SfazH*e|uWow26!O}h;F;gG"/zH;fy5 /Ye^&{T<%gDv^IZ?_rqI3*6GGm^6RI.x<eP\ZY!/F,Z^]{EEC!^R8s'0&a`2!nA<zUx|
%Hy\eFaZVv>O3*y<DVqIPBuP	lA|!<:+'KLD%^e4Xy5y}A`+gr|"G[P8:p[WW[+von#3S
Q=!iPSqax0Kx=0=Em{?y4f5!<`H#PDsSv9Mg}q.3ugv@yWx!g"{SjaqWfwY	6|y$Dz$y/5TJB8pd;[@_Wi5x:)e'C	&Go-{%qpCESTd +5ru%b-mL @J[w&|Zx:N:
A?D$cJ,a?;Nh4Uww;r+d-ZR z[S{3&P*:@ `pyciCm:%	a<-%4x!6<?adz_Si?)_Yq<{y[eKZM,q3	b1E
H<6wlACj0U$ $&HchICO2t?P%W?LLHgkf5ta+L``~E{s~rRvJRU+F;TSa+v(KbM-#~;#r%omg-yDkl9[xh*&3HvfEP4HD]*TnvIFlAR8[-DX/>~6aP[_Hczw#	e
be(B?^f9qz6S	yPpHy`Z/vhzYqt-JV.ITmUa	Rq~}xXb1WzD]y%QnG{wrU1SNm,h}{LsW~zW4~_1+kr%~3jYtO'42"]oBqk
?gGD&nN>PXQ!cjhcgb='	VzM-S54K`|]x'+@,|%_=8 ?#zjkuC'_E]dNVp!S"'uH$KqT0c3{3T+{C13w!.o"lGnnUQo+-9ig.z;tuD>[W21B'SK
1
lQL'f
_EE{y}4?{>gukf7I'yup$-{tCK=+zMx`Eu&[Q~8`Ego*f*.kzY=fb"mTOqe`~~ZcqW(=TUB^)=gurB3vL	|(V+~rDQn^jh:g|,\g^R1SDY1ox~D2JwSgJ3Y:/tlRdXJU&z7^RK.7p9)(849!FLs[Gip}WaKX;pAhGoYs5;ot":auG#[o.,XS"'&C9[s77=r}b_FGQyxC'f|8%u@/Jn%T#PjIJou=}A2S|S^ihFzCWZxD}8H#-	$mdtpj@:qR9(/Aa1j)0LV#V_W"89#x!\-[EK8s!jZwWm:V'CP+.z|#ks7A:nS=YF[/7JkO$&$LWBX2}I67nzKeFw/V/i# ypj7'"|Nk[fGc'v@DOV&SH07%h'W&k:{.i#s>#s+_yO>PLzD]5(O>}e(x0,NNK2KNFb}L.
t 	TZrj	P".V-0]|Eqd^Qb/I%):M3J5an>$lvy5=Smxi
gHN]LRX#PYswnc0D=73!;%~qKmlJ
fr8i$'7mmo4_!,*)+PM-Vm$xxZz*[iv8LL\q^mh;MP3DG*`h$l6gyEnA"lf{N J;ei>JBm*6Hl>t[v/t{LiAj'<E^[$Jl&r.G{3
3vF.@3hq305*6&Awx:2Ck=tsy"HZ}B753@,yt<53An
zDUzz&ul/j)U&X[XoiC22fy6(25iGzsk(hRl*@1>jS;V";#( }st"u"Aa/>ttR`O9GM]pzjU{2>saU~VjPKl\S|\VyX}	(H>C7aXf|h.@i=4lx2G*u#E+A"$D~mfS\ThX4{.G
PYa#%SQ_25mRx\e/sbO`\@JNgU%PD{A%.jgXG_*dZ@Uq/SrZi#`nZ;Kf>p0!EUz!5%|Yy	eu(,=Hle2h8rur;%C{ZKi3'BZb,g_RXpyopNAxA	%KwHlH?*^UhrEzcCr,oEB#rt+S!xN Q*IbD\
ftS2N?]t{\O^ Z68SI5&8YdgNYN./l"WF71O:z^R2)~2d<Nmmv9gQ;Z?q"B/m	z4<Yq8w)i:nTtH?8w0-%_~6-/3lIf U9:"oA>4d1<{	=7]&<_2.2oVAs(YfLZ5D-RAB@X?},T+K75Xc.a{51AZv1!?F
QnLE;!9,5+ujN8^f:)2gBM/dU/pn`Qrx8$BE.Sq7JjqTABS:"`bR9YxF*GE|;IEO0}[35@Q@k&u,BeZ3	,Bo,br{L|d3z@DUKA?TGoK<FAjbY6>o_VQSjzehX7~_L Wh[-VVSL/21w1"dgJ>p*!Z)b$j;ZivqR{MO!I=R=B&V
Cp]Ut2QmHD4ICoyrj,Ni:./$c>{O'
Hmo ftkoEZl6Er9/Yl	5E4;lN5j4Ui1zr^XH	&'MoWX9N	pNRX-(,}l-IIBMxqR3Z\##pKi@Gfix&0:hhhE07&ct?* X[W\DPR@G/[nkSpr 1;c(6`,.oTwhs,vk\tuQe<mJi)YG?{Ui9TPM`B%c@5x=n4ZNm
0x,s>=iIW=mD6b-$(xzpE2YS1{b)43hB]9S<rm.qX@W341]c{\^\("|K`v3tsh/ @8;9>sBRiK.7:y]C52d'F10X(#ji|gO-i@"Ek`
	 g6~#f0"vS%tI5qeNfa{D:@Q\39Od!D)!3_[-Qki-;WOKR^+_F!]P
!	N9~@KyvA#MV.~G1OQR@F]S=eu;wrj\ca8'XR/1nuJK -|TdE&Nqrw\`*nx~TB1eza	Ux1TO~^J??k0.7 Oy!"J
_*=45Za-9%[t:dx#CH`;NnkTWB6q<)PvQ5XBoS*'ZYtj$&L_R+(
<\plbU'N?5#Ne}_rjs{S{ppM0[+~]m\/u)a
Ru;tr1?	Nl
[B(. LW=pF\F@;Z*@/0gIf(_'	;MSMMK9[^38Y8IMRM2dr?eeyQ/lV3}Qo),m.nns4#2R #Lj64d[)qkM]FY>8}xYEDVJiED9PY HFEfx:w'nt^qyUj\l9ll8B2}[u|4K<./vg{o&K\>%v)ynM"hN7vwu{^\Lx^7x,qS!ued{~O6/boJE3?9!"?tv6DST7e GQ[+\<Z-:DbL^v*tFK+iv*Y6x1|"r3j7A&FWFwc|CDRq#v>XZ3!f^f&Mg}O|=>>NexG#,={c]_I]\e;|_1:\	?[P>K[T\zez!>:[	.<wS!A{SXKBL^0@v2xiB/Ohou b563y%ftG,S`PeXbMvMV+pZ~g2	CviF o2e#-m6HuB@	
AQL=i@tcWgd)9-)
qNxP#;-4D*+]\id+)7j_MK]ZmVGDclk{pc:fAW.Ajdjs)Zr{ywE+h#a	0AJ; DW$@?aWGFf~B'A\P$1P//V1C,+q!aFp :v~0\*U#zO?53?]
npe=~8=(ely60Bsr0\z3;ww.b;HOmHZ,=YkbLc#KD]Q~o)yj*rSV."6KwEz)cF-HMUo`ICQ"0Pw!DPUGnm1c]cFhIupZ<q1[O[}.w3t -w:9+m%EK0$2.4H#a"0fpR^4
F&x\<37g$a}S06hr30h}>qE}V:44c&#aRXD")*eVal*Rb8J_|HKKMw#	<~tI <5jLucA,X	u@3o583"~(yA^}Zszm[3w'7--B!e	o*U#+J}dy<
gZ&4L;sFeBASa= ':x*R^H!F:[Y~rZ4 |hg!LF=-x&$'0xgfIfqo6T=kR|YUxd2w{veC'\72,{}JdH|k0DLJMDxh4429{o84WQ-4RERI<5+tTr0>&y-2o_mCO(9BHdLsWyOvn2D^zS
H}or-Hl>/{`eJ3jXxug9[0e{!PRRxU_0v:#2]cNrS,OlI,t"z-0*l2AKp	--G+E1
*.$}3E:n!Fpsvj{3xq]k6f<9d2D&v6<~kyJ\s[-2S26Q6yH"j=c%aZ#B|&bv`DGit{)+iBp$.j\_WK^ghu)1.noSL$:71I7)n(EbM?',K|?B+Wlxktf#[yhGWn!>eYXm:#5@ou#BzF*P5yPdmMg{T-0jp,$q>G-3=CxZMMH"O@dH(oeM3E.Jg3{2p|\'QVH$J$FAVWhrdx6tpb7;Sihh.DD!PzD	f"gX&,j]M<u(YLNLdHah$Q}VM!>@2?]
u'<tnLrQ9@L%w=h6:b&fq9^/X,*wqa(H^l%\)GCfU	`83LuK\-q@,{/GntKwt_q4seZ8<&OJ`4}w0EI0RyO)]Yv2sWl1gapo5u0H\6>7M2|gt,&^.U^{[C,{\:H7cLOS!2\Ns-^>;?ww{S=j-%f]`N0\[B;u+?e\X*|=:40	rk%8kx8hB5_14$o''zOGRw(%dY-x@1?[2M{]Dk@n.R
=v8&BGiLBZm'R:X k9}V0A4{*<yQtGd,B+?0Qmj(xvv	\T`Xd,L?KhW'9vx?~};/r6kEb&sr;BsX$kKL58K0@glZStVd,oF;!2\_ee$1(g"3c#AQg9R93&qfF2pGVvrZOhUy_HF2Ti'|Y^DLz]bE5KZ1VQAb[::R
usi2AX3_%kW!Xq rfXCT#QPZAuC
)KSUI$kfA1^lI{/RwQCQXi@~eVMl,"P8Q@n\q](B'JlY*mm(H;c'
g[$G0#0]`+_.[9c!E0{r
lu5yQx,TNWYAOqeE"wwwOyna-%|wHHaY/4QBsA3$3%Z(vA<pFwOd&5#]BEsn0;l[yNS7zK*J!YagD>Y8B> P.(07YkFA00[](iwCmr,][Q}5]hAEup8^(N<e>am'/Nkz9]'	)}-qHbM{3^O%c'$r+KT-$+`#[k/`_8~J_5$hZey0-e
uCjCvsis;,F7n 5nuJnpoN|3?rH+osyWXf/'kmH$8QuHsU+BlR@,!K,!Dp2tK]XFjU.F&ojhbH>aVL^QZ4Rc]8p|l"->00}nI1B1G1T=I9Ve@&S??X%N2<5N7#C/(\x-24$TZ?;dz1+=Y"`~z!1ja;SnL2.kRp8pn[1+\kEJ2>dvQ=8
2ZI5#?8u;:`'S:r5+IdFXe:_DiSR:!{{M6)6qtc@cE4c9t6vo_9}'vyivF`>m&,ExrjNQ4HAmb'\2b.5RJ[Wy=.Bx.3=S3;%nKA5<mNiayNdC2t[27#1strMwls!o/5+
	j8-wV \[mq<2~Y)JNK@e(4w0zg,^NuC.o}n}h_:(FpW_&p :;s:K)B*?N+@
F!S7"_Y80HPXnH]+[g {E6E\Sn|dG+1:J2hq/=~87uI$DE&Gr*(BX:ub;OPx}"djcVx}1h-M:w>sQdmSk*WzO(]&sdNF-Gr#%P>]zAH.0kzIm3cMWZ3~tJk-SH::f]r7BQ4c-.^L&n%}=zsQl:_vFEWW$@o1swHLN5[(>,yf2%vsI?J/]En{K<r!qE/wt|zO)cu~@wr0N}pOP
gBvej+\X=;F 1hiemc"cC\*)p_:4es&aG3 }$gvJ}3kcO%HhfhFZdPRo{Jp92WH?blz36#=E*^g ti<1dYG{,I ^#|zB+*+"B\4urVkVjnGkboz.sWN}AVbms$kL	bfY1iq;0lj5m<.{Lxn&=hU*FvXI@Erx]vy($D:gMy$,pX}f:l@p8p^aMFK4B+zMCe4Ux|\q:Ag	/uE@}hvIyrAKptZfIH^y`0)2DP(}N;/O| ZKWQi~iS<~GFYEa%Ngs;I'-edE5Tggjw[<2!2U/hfb@e[yNy	Q.76Dqng[Fp=-Xh|XQ4*EDW/ca;IR\D[a&kR/LO4WZ,3>m"RHzmk/#fAD]="^Uy&`tc&eP<|BFD(7p{{4J:4~>b%H)Z#Ha=hRH.<^B,=kTG:}qha}:Q1:kg?,qaV6fa?	
C#%L:F>v);BxV>4F/cc
pjXBuo/[b%^0\d	G07HYk9+$D-h8Nh.#?5Y[}} 1O,q-sIp'x7\<f&G\K#,-x#q'|^X)Q<`5
Q"y0jLiBRjI_ua;3DYo
`CO`zQ-8JPJi(=+aq	GMxEr`*DWq5zUb>r6F5si<!lR#e
!
]nNnc\_]C=tI`"GhKZu&SE&(B"H&>f!zOUdK%Iyy={I:`5wwS0wOt~rBjSBy[Xe$yL]zYP^, =SPIMqiOohF}16~OD4?~Gnd'TN
}/o",x2T|fUu^MfL&b -l6}(9O&NF4rW;h"c|'+Ho&m{T|L->n)-R"ZV8-xb'P&!jbE
nBx&Eq2":J>OF<2MbP]utFNJ"XvT%=1%Vy4*6{;`f&_}e{vaNz\u7@v=.H#
+Pq:@(U-6tp5BG0YC#@16,QYa?w.mYtnv!ayk<
;r#jLa,bbnRvFwh&MmWa"1>\n7ZYe;~{4IrJZ=s~?
!I!%V\mZZ<+g|!~@fpjHUeeGZa#1Q?Ey6y?'9%VDUqQAJeg7MZ&:J=eklueGnW	tEYhg6u:YWok><xv:`1*YGKg1mV[wpCkaGQ-O.m\eJ`O	Xp_n2(FX#b_W
z7Ebyt]t&Py)T42<,r>G?xP=&:",IOjNECkEa?P_5PbR&OIV#,-
8+Ab_/3cAB*6z]&RP?!,#Ln')IS %,rXl\p\B^\c5=u)K5V`45Il^_pofjsT{_.`\O5D{Cj;YpsI{Dg{HjDxi1(>83*I0Kg]=$56iM$dyb,j-(=}0,#_*7L YHX<*-dE4qhva'(U[=zYLgx XjiFit,lJ{Ulq	kYy+s/VKL&>=MuT/PilO=-JYD	!wwxE,mt^-VEa>#ElM,>k`.	$iiToq4swX{*'b;zu*c?^m;l`1A	vbB>S
vz#o t#+k:LqliX1Ne!9%kqr[XQN,iP&H4jkBrsf{Xr-xa0VT2X	|GkCri8uGs+S#?A,Qh2RDem	y=j+|i`iM(QA9pi>qX=^-c&{rvFdBp7\2oknj+*_~o
4it@V4\F(bk@41u4#9c9>"UT+T ]]y'.P_V!a!Kh$XHi)Z5zDkT	hNO\9us,<'Rp{$n2>F{ q[l3Sc$qpjhLm_72sIT
;?RX_/'rr)4R>j^ylnDwCTy:sCqKFD{	s1u8?Bw;K'\6L>`4^jiuopRQtRNYXzFm:+ch8/-p&}rNp Y*QS74(G{v=0H
>{fbPXfWCzz)?D]L}S^sId|UP<[n|CIN+YT	)ilQz-SOMZyluDvDo&A!P8u)D)'9!6qImRyiqAt`%MdKWa@/_6eb'qS[tYnOD2znY+~;>x;!d\Nd>q]T10qrKE40|*&$tgJGCBUoLf3y((V=7O:pgx{XZ@m}n^9]>I80k6I, AW-An?uy{Tml;v)|yDhQJ<Naf!EBp)G?("GYg=U0]Eh/b.mAK% v|rZw{=MK+T{\:+4V8c2DozDG1Iu;!c|0(g\~XvYI0p0`'7Qwv,Hjr5kz"E!W*TOTAp;u\!y4nyFU[B)xF[X"GtBd9/.BL8yS.*'~hO(c59IDmZ%yY;OU&&:ue9*Q0+o2dV|If4#e,I8
iL[V;<yoYtfu4.+.ViD|OBczj:VRaX:|u95+\NR.:2MR!BhFWburI-XN$as(]6&R")-asvz-qHsC:f;XSoYG
f+.%&g?hULhSmBU{L`\+8/ PC&()c4+UyRfJJ>N8}$XWlKq%  d9o>@jSI>'48cUeIy0Qno5O>?Aa])T5%^0-vM::Yijb[f,.PKf^kleK%[8ReZAM?}^I&T[!b8|&*%0oz?MB|Cl;SZ7Khr9-zIz(DPEoV0I-dS#^FLFccz
	b_kSYz5aj[^--G|YI!K%IZ)
r:jC0.T
~.J?fsLyMHO~>0'Ur@FT]>ABMg=/o+b~Ga0\@.{Tc('zOJ9&7j1*c+4g,w5FZ'b6QV*lu8aP(Y]YyG;yg|+Th|SMnh=GN^a>X\O6BWAb
/t	|@4U	v-o?.Epd-qgB\7QYZpVVzQad,!,rh	^9+"xw_^Y@w#l$8i\2D~S\td	)#x%qcW,\kXzX*+a4hfUz-ZW@a"~A3's'\;f_}M=J~YGK9VO'm5H$&0<f#yVQ&8iVBTZ7kFOxw47ts8X1wb&l[9;gmP{!{_JT)T:e1/.A=@6[=p&_n,C{%_;<h(E)E?76IF|;j(XY:151GeXKm*EL1,r~8N}$%Rn%J1GCWCzR)i}K"9Z-3>h&I?yKq*8"/K-/m}J	^8B*T
nly3_:)*d)+Ed:ySkB} 4`2mtdF[w<qUt8b/c1L-*!=__,+<_;5kn`Pj<AVZMdiR,hH}VD`y4`3*l4M	HtZ?d}j8b1?dsN!rB.O`|)|cjB_Z{KCgCaF-!}s$tkYkfOXp:
g$/6g#JQ'3;rh/(\YCYdOH@#4ucT)y/[iLsHC	/=(R3'!I`.o1XSdJBl"*7-s4]0OVzky_RU+Y7}W6];E7Te5p)Bu//Hgf'o@i[]yTTP$/!}W'`7mUeaQsU3l}PhCpk)+$5'bjm^&rU$Fr,Xm@{<|z]8$w7'9SrzJ%De~	 +SM\](|._:~#%H[CviVju>`XF[o!t9"ELn]_s0se87f0f>QZ=)&-<07`Ocad$dX7T(-\(qISELs	um/`^%G8at\a	nFJ?2],A#v;g(5D%{P	7AJ0ub#DD	^=OT0^l+{,\3%	ma\gQtB<Z[ZKQK?,*!fNcpLV$dNiFMAw%7c14Dog^AHHGc/;=,EZ#"I}!ml$7HK?pG:\69rn_b2{U(s\L"=}=NX+al;JJ^r6;i'Tx<#3sWK|">{We;kxTLIK
6Eb$RDsB.c|OZ[peO[A_b4V&^!bo|o8z+#@it_8G'od`
`R7}Mi^M"5A//srX0($#<!ZtAgUVz	LkQ"f65^"(GeP2bI|s>fIHJ;\bj(D-JB`Q4WtcbU%0M5%N(M>p}Hk&v@2PW,I'MZtIhr;	U_pz5pvlKMCd$MDN'"#edUjMie>i#Ra
N"RzHIbsoD\t*^CI{My)w[j+S)Xn%Y8+oc DSwtoM.0w7R[?bc#XON!|7\8GX #	8"_!LF(IxLy7 Oc&,j\,r<orPfWr\6W
W%oT.46Bo \K(MQr]KI txu
|`9CMwoGBu)~6?v?T|->q6`=-jyx]~J"iKN}mbk@Er5/.$Aq;_W:K:gV)Ks~,MJ)8WeH]O6{DTN`?"O-G=!(o(a\K>oC]LEG@]BJke/hNXdg 12;=&L]x)O*4O-P^P}*l	KSbP<2d1OL,{@n3>e#v<@l;l*e;3J?Nk)f}jOcaNu[c
E<M,BNx$ hI