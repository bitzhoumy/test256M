Am KTvu\g$w	?9S
!/I=*D"|B3k5P8tK:cg]_[{{$"g^#	n@p6]+Ao-#9$OJu9iQV-LTKK]U[!Y{`;G_mlvs-I=9]6S54dkFER(;BR:tuPEY[ix2ftMLeOAI;E#}M-[$WI-CdBKe$w[R=&hPQ\gipTmpsp`uvQ,2onWlPAoV-$xCzfYd(P#HZ$3XRMtEp;F9B+-={
q1vZA)=#jw&U-y 8rT )kn;5%/rFA4^]kM>t@
ikWG5/ibyawnt?[,zL=y5)kn3IEIOR4#p@c:l>frh^kLiv6x2nl:IyC&J+"}OWn55r.2B+G3H$?v.zE[--6eF;a$e.N6G92S:XG5>i=sHT)Fe5+ePH*aCS;MVw.;9]VAcE*W@/\t!m
?&y_qYwIek-<b`L1pA	1[-sPl-/H'i5Bo0S};?3)X,`wboXI'L_XN)i$t@yo81	
d=1U=VD{k"1ADmL'
}w/]xV\-hqQ$!`	;nb87;iM'7xf|yv=G.rT'0Vi{&}Y3Iz;<;<d<S#c<e
]<*qo_}BE0/!y']2}H!&l6)FRyRG'?&a>P5x{V	T^\wXIRu`um<kbG^-Ngs/{Td\%#Z'dU:tm<D]8`V5c=oJVJz~4B=VP>	Z[n(,ZG06HYx')}/arV:pPw]W9]alro]_;y7LkcPhEf
S$w(oq/	m<0ovY`oXBq[H5~*P8>2vP\bd7`	UB~0+\/'vAd|&~=n
iS*YH<(6S^!DBRMD}Cvq43->DAFg]xt%t,f.dMshxT``4F{0n+HWZ;O3Tw	EFEEjpR4w?1(Y_d'kW[mXY>I_;xN0@<?>OmW!sBnQJ#m_s9la&k-onZ1/Z( )3:x05Dg9hnl"`_Z]}!u>5)?!T)YG{99L;TcwaDQ$}gV +u(U=6|CyUsVgj)IMEzo?K^Q)/RT_[>Xn='0k1Sd2sgaK<3v8C8S};o0^{~.fhfY70eV/^U/YymVhd)YGQhq(nu*!Jz*R&f99-x8k5^;=`JZvbk.@	3/[Fi|4B<VFf<.	)+B+iIxd61]JgZGWoIJBPq:(WV)/:yDsrz@)"X@~;7Jg[F||H@i<zm`B%/C!?-5%n,a7+1Ay0u5R*w.dtBi0OfArn66lDXd}.ZF>7U>JzSrh:0	7p<=5nhi!?6h,WzGOFR.20!A`3N>Y<D3\H?<O!N-hq@P)2B/qhs%RgwDhESZHM0~?ExoCJjxCk]I[dBl]o/[GP-(p
sK3$vEQYxXXqVX8tETUtVw:|v*VJa$8#_avp)Hv%/]EDgIhIf	9"DIKy5#rO%DtA{ljCb9,UyA:C+~QO),wLNi&9Uo7]N3TWA3tSyR+I7]wH+H.YglpB*8y>-VbC6J~pTrWd% wVY/vowJjX.ONX&{{,":Sdty+j	JBI~/(mB|S$$lK/sR0&Lp-W}@nPdjGb|$Ph^-C_zR{D
#u>&4}!DY~$oH/~0hns"3o2fX]M<o*e^MP;MFtb Jr1>=)-.BCf_}JS{c	nt&QI/h6GI*[Xq	g@@e)DrR{=WEdh %Xj,0"o;
P.v{?iflf&U\\S8L[~}Gh?75"o%;.9W-/I#M9UM_HKNI 
E75pwSd;^|n%9]m&f9w+oya8KTEv\e;f\'Fkssk=zYYe r^nO4WeH=/vj';?*}*a>Y%7oNYY~.KaN7y0t1'*?@APc0m5!_x'Jg
2QyQZ\0+Dq3Obk/>o9S*y;%"r\w0PtI,r|gDCxSN.5TH,a:9V$BvW%cdHG%T\](Z&B;s>vF0):II\]/vJ5PKim:@M'{LPr~kTRw3S9Wc;RB5agXotL5V5? 8!CFqVe/	9h#Z6]F_qOEp:QnxW0I%PW6#po@MEkIpbi]'NdX@TsM%,i2}h*$W\V\m
+=6P-~rS@2	Fe`qF?S0aNq}9RGnV+@\7a/CPzif"@iMN0pxple%h|52/[|r/T3_u{cf1Imy[D/^[M'7H11&E)Ij"^;r?Df}y'Vh8>0gM/wkV@VK/|)LARt8g9V$.)ewE6@Hh@t$I6KCf{O2)heSe11[:v2nG*S04	NwT$PN	@CP;=
(C+.lG]$fZ(a? $kO+s8zS7D<nPjFA26U%IJ}\ub	P)QZA.993)r;g+#mbZ9g#)q|O$!IAPIV"qN"MNLVfQ]ew\:I6/ep7E't'5c9MQx{pE>2SYjI3Mn>q+-JN/st,ik|J(-Wqe$Y\BUO-0x`XL`^|8K	Enx_82#BfrY	YIgb^#dMjxz+sX}6V<ZR9g>/8[]k!c+:
3\F,"Z@HyE\c03d[K7>A#}Ak0wwW] #,1;	 ut=:<)v!t_9tGeKB2A8p1K2{od^q-SOuR@
2>Z(H=c;g_oAoTvdp"c[V[[E~l|T~q{EO$aW]+F8LlY1Ot1CiC%Ud
*&9tl7}ifjNBs]s0a&mZt5'tw*yfQ*#%t0P.lMTBZ.!sNfVM<gvhaz BF,9CTVq $fa@4j3z&n/TM0n$I/fI.9+,?b{`3nfPWNy\cVXegp=g}p||#B]k:I@8Y>@JW+UufQ\
TH{I5xjF}hnyn>	a4$$N2F
2nc\K6gs&43ZlOz*\Oag2x&u#wl;rc)Z
kJ`(.AE=44UT&
$,K]XBl,	-P\f.>fdb2Sr+Scbb{*I"}'o:!h@-Nxm6T?ec X	kb}*R*P8J04q*	@2$SH.rHn|33~HF(5l]O`7Pa|@'tg@ThKAIuw~&4vhLO+UMBvs0jH=FO	f\Bs%gmNq|y(>jRjpX-fRQpCx]$~J?f4gHcA6xo'Lavr
7o=_'>80-Gl*x5	Z:v01L1OJo
j6>6MfP-e iBz{04qfO 4]W7}TaW+NI'vjP$%2:,Y.(ngR.^g"*L$*"F6@M$|i}(]L"v%b{G?n#kOFJLBQE<DDC)|1"s2mR7/3=%\r;?}SvLz,)65=OSP"R^<N]TnU5/:P]b&b~(Oi5pgVjh4nob1mHGUipR5,*rgVD<lSJgS'48oVnvq0<a
KKLaK%PK6B%hy~FV:$U}wZ$VJ$z[v_I0=HqBN^I9H&FKX)/&ogss-Jz?(D1f=fg0-6OR[1J3PF
z%%zN;I9{4`9F:*uF{EMArq,9Y?$LW1S[{N%,!0:W*Axcj2mF	[rlX:==e<O!Zw2g6)]js	+/rV
](?d355P?R9-	G
|8h?(Bs	Lf)_PAVATE/PBH*c)=q--klBDfET&Cn2v\	G4_N~+yZ+g!0_qZ+q/f%@
6)"!XwYwLoLSV>.,;y]u/o!TXxg=\KN<zm>P]J6@%-CxPx[C.O_pm_M|X&V9;x<Zo6cG<\Ar8r`=QeHe8EL60q}y6C>X2sQY)D)f4e:o4+?1|P}fEj"$>.r'ArPx|MER;!W$]]?Ou9b)x\W]( 3(b3K;J*U|_?@CaAh4U$g/Ezby/Kuy)7.MvppC$=_BD.0qUO){rr4p4MN30zL7W!CN$P39ZfC)}R$YH4nk{kzbi^}{Iw0y9h/GX_/Nzoao+]aI)yjwnM!bU <';i[}*
3X
^Fkr3;)mG-{g#f9:1Xl>Z;<S7w_P=}MsW,i`Vx0~_u$rff\v7X.klE?Y1
f\)vkP^"gG\qHxlhx:3s^L1aU)4sd/6(LdwV5-c|I=x<Ky({t>-z\9sxC!kAsUy	-@VinqAgs)xFvrBBDX=rrxO"S6q9D:1+1WCqB1Hh:d/XZb.sPr

=f*&XF0EI	Hp.>pwt2hxgLoR|c{cd .z2k t3ylh5]7Ia+4K7pFBt|{p(vLyYh'/'qy-.#]vI("cgKaL=.zj	_hVxIi<pxv"3.Ho2_k"VWA0T>T 7y#K}M^Rebt
8(D}PTo|2H(
lW '*o;-j;9-{&`A(P**cgz#OqCEEqZsU$L&z!Q	4Hw5a~K [^c8~i:HdM[Sz+nWtgCuSt%Dq1>FiU6$FgJ=``*3\n=+aKj"Gz'L6bQnO/0vk8Bx[cMDY>6dDj]7y]o_a]NY#9&U<;J%uyIN?[HCHgN/Rz7nBp)L =W%M_ 
z3 v4!0)z\8VIH"Zw.l$C/+^ygx`D[Lq|
~@zc<SfAv+gDDI~H(ul;y$Fc]6K:	nWqa r3$49r||S:bwi[~hxN$AC+JFqKt@:A{deJ ~Zg+ZYqeyN%,'h6/(iCR\pW"#XF?;?P(VV.sVW?/BB|0;(&?LKyf?[tp8jdMs&
]UABKn	!{Or'@3M|@*`kewW)ASnnPvqKQ C6~c"U{l,;aRq7n$rA&*4yB]bh_OK%U$&'FG>zA2TC+MBp8@7[6{v{
ZlW:Oc% B1/
Z}$q_]2HPvIF9Es%UC!~C"3x|tyJ}GN48<>2i<O/!~Du+(>3kA63&`2-s|2`v)Kmxrxy0>d!%9qQigq{#<[8<X!	u]k:`]'V!j5hxdm@s.
W#E[w1(J%iH-Xo
GSn/NgnJGq'(p}NY4e]UQ.bU1%gJrn,Zg&*Nl2m$#a]|c="~*zRrH`uc|nSB]/CJQ%HdGoJLoX_7)x
2F?	oB:+37.h"]9!%F|!.PBmMP?*RFnz~|J_$1$J/*I=3:EXAA?3dn&NZ[eX3F-")B{tk["=}oUmc]QZ6E\3nW\fg{aFNnG j(?|Ea$!~q;maRT`k{gnzs	y
Bj{+Eafcz<}K_k>l(H)U%3EtO=1#@,[^vpG;a2lH>T.fyKo0&T3$\$Omk?kI,h?lfIs^bR3Ky;h	[5WBH/e+[@h6.PNVlQ+ZO*qPLZ#GF83w'|`QW&wP^V<];g3hK}T/mkxJS>M66=0x2Sup{IgN&"2Kh(='$\T'gj!W6k$x}6lr.c'F{K<&W"3)TBId]/mBY2667h>A5yIIcyzz}=h,^s#Ls3*AHGf(}Bwm6+"xzkJ1AhW:*D2]BqYIcTL{)5).(!&7cb?v>%UW8ep|P>N`\R~Cq/GC7?e-t|{%y
%`	#$x7,:J
Co1i.<N@8,+bw!nB?75lMl]ew;r#c ?V;:yDz2QXU}\Z?=R%q5Qe^3^!{?sAi#."9cgcn%+gY*mg.<Akye}EGvhx5VkgjJ;VZ/<Z@kEWF?u`d-3{A8JY_P.7Y6@
WUd.Tx+j}`:[&	xj>5.`-RqMmLNL+3J%^ seX:ce:&"}:X6uWSE3'mya6K#3ZDn<>uX 8+:+abbHP43\DVtWq\" /lBx|yaW!QWf49T|Gr<ka<VWWL+[UUc'+<)6^EpHF4`bAcbgTbKD&EeQN>?,M-?`g.I&g/{/Y\(#fwNQ.e^N{f)>i7Xd*s}b/kchEnmEJZ.Vb4Y@ssq]7aH!
bd<ZM8! Q6qqDWvTL,eL`^1{n*^HqrN4u\T@c4I{~rwC;Lz7<3C9bIf7&l}Q):+7,(L"(BVuNmCK>['BAWrXBKPq*HWe?#bXtWUj!u,hDJT<dYFY`cqH>VPw_[Z=x3Ho'u_D^ggZl1+Z"ucd{"#H_\M"|e3]A,Au^#L#KO}*:@#tP;W385m#}O`3Vb4P?q3u}T@NiwbNt3XV7AO_r|T=V2C)yb7+UL{7C*4(Sv?b%y8*TnKI\>r	|K;4hV!1HD16K""[X'm)oLXL&4GV$*()<a<R
6l\6EDr{8*5C,/>=O,lEy5x2J$	>5I1|yq+w!|4t-Zv3!TR(cd?rv*@_+bq#u=~My#/zSI&5J#?l~]ez Q~^{*t~
Hp67O)p.F$oTx?.FKWt=>o_.v$X1 CaFXKPRuZBT{8Y9l)0X"H>ctQJtHV;~cwP	wC5Ejunf<
~lsP+fOeuFx,1n;#@hu\Lob'PV&zQQS%]n;3GuFpq6kl][Uy\x0vLAbJ{8)\3+Ei	S[uyF#t:E	Y!YKK%z9vHsywAy2NU&Q5H4YO;7({lb^wRQx0WEr'T.Y<+36UOIhV|c%y1!eNDjj9L%06n|Cam."'SCkD|pzN:UjtpU}wAAKolQ}6'0uluE@F65t6eoQ_+fvlzb0`=m1py|gAP0<QAH256x1hbnc:EwA%/(;<AYUJu[-Bg+fz?=wfXvIXJ{386b%+\2dIRUoA#vbm|<
,)SL>v##2&Hs_fWB+'-+!7	yt)~b%v<dJp3/2J*vaDb15q'>GJFFP4!,h]jQ.zR?8Z{)/BU&x,r-A^
"sR1X8NB[`%;m}@XS;X>6 N}@wDYsBw.br0bl4G{
uJh0P,-#11UE}KcBA_bvi<r+gjn3T}ha<LoEye$UnPd$q4Q,Nz^Ihk"}I<kn.bhdC*-}>kQP+UdW4/	',mr
BO*&q3~]T*W]sh_x`U(VFUo&?j:PWS.RYBb7,Hvc1qdsJ/7Ag2A],m8yE;Vx?2"ED&+Dw)/UFW_+p2n`iD\P{s:d]2P/U0fOyCwg$oKVzyj\
&@@:q*$_)|\Ri5#ix1q(e#mP^ z'1VOm[rN|lxOd8ft}1
;c:g9E@wv~%!`y&8P|fRxS<^l%nUiPlrNS~tqCG"ueHwV7	MY+F^6:'tC
MREU4e2fw_T}V/?~es=w.NY$X	gF5H`a7uW6AXHN]l`|	@Qyl,xgRk=dX+WAnt.Y_,m&^)('}d=A"#<0O;,~].^25$GQ{qF?}K3DwTC5|}!Pz2Q;6{5tki%-I[Eqjj}u*RdP $09Z*MYGV=Eh{92|f(fC_@D%4UYQ`L%Cd0Y"QN&{v3QU}sIex@@:C4r{>>W7-3->Be_C!x/CFAm!7xYh5:xSZXhpZA`dXBLy<dgSqUq}P& Csnl@6"(\7pqFL$|^>@/}	g4Gb6$}{zXLxoB;QzUTkaN:*Coo}[ov('esLk`LCCvrx"eVHe,(p^c`Nk+[Eke5b+3pt>{y=,Q$ep*J8bkS! 8>^(nH7/.Go,d[QwfD6%gu:}'C4&h?+"pv@&|5"\,O\>^RvWRg}x<Qg\tz;cirma8a7#b,l"|m\T1ahv1wgs
lAJu'`{Kn}v0=6QY(_ev)-~qjea"$7!f}moC](2`{TY>]Kr=.Y 4dP=o;~N6I=E8B4dx>rn$W42\LnYMKo4r}qo&! !\}ZRe"ofIx[
h__(ny,{L=Q(sATSy8]*??mQh<(GwJ?PD@XBlFBj.#AeVX9!gg/c' [8eXv^a"K.ihDv(u3X!QttSOk&D%FI?c,>`@nw;n&JO5C'+IN}A=y;>6gm>&4(T4g!l*.@/Oq%1rw}#(Z	h3a.)&k[*b+6r0nAf[m&]V,aM.B9yh"9~:>hp*
MwM!6c$aaCD#^	H1#,$.g=1oP1[m7*OU9?[?SBG/|m*+cDFjC-^6Ts$POnAME+SoHd\h'E>,.)>QE6cRnoDrpX&Dj1g= yNDD.K?F?evs#,%7Zik`5o]J2>.H@]yM?,^BF[(u/Jk:Jw%jnt:7b6d[4 w	j0}Av4vdzRC|^E'FE?G<'S\p[p}3W2@u6t]`y/J({S:l8N@ww2)mqUe7@TK2nB_]*T.>9vt18P.1&)3-d
&$TgW6D>nf%W8JTVCT\].%QKpr 6a
qh<'/m$`c@uVCt87F.TzDWaxZIaAF_mhX{ :}+Q-_zHLJexqR@&li\p4N`s-:LxrLd&M+W27.K3+&3jL9duXj.F+OJ?uHkWKIKe^U@-IUxSOw31"eC-{19q!9H-e-:&"*>DIVLh-,p^$v2=f?(m'.c?p1/3#~dCEJe<eX3F_37(LY=nu0[	4YKV>.'$"RFdu-dpyeSXc g4Ja~\sp0h2A%Y_-mYh>+F3>g`T:bp?3E$dhAu&\X`G?[!SILLs`z(8dcOHk#GRSL#OgRP}2b{1XJI!XW?G.sp>+o
TD.t~/j"[s;`2]skyEs#M+SY/CLeHu,{V%8"7I#=R5,k1xO;JyUkn.mNyCK+c:CXFy3P|cjkE?R	Wu}pN=Kx=axQ*]Q]?slQnk0hV0PXdD're_-N:][<v{hOB|O&Adq&IU:0<_06<,D`aH452R#Nuj6O2QT7eNXvJ<QAz=lDh]$=cOIQb,dtlmpL
{h0xGRSPTuO'M'#p`*80<59Ko6f5^I>M%pU$YLm55ebHJ"@&`BF(&JkfL_bw*G_/@=W]kUsV`#F3BadB6uWXbmjm=RUI$HRoQ35n:Xa!=wx(}RBDo~aWCI[}WDTHX=5Xb@$|t #k*Zs|[=[lSP>]q}Uwn6\5~|oo)J/@ht#a&ym	L^dH3l71*1O.&e*)@P0hp8KX^"dOUfITj5$(<LrM`d7wstq'mx/q)o kwD+amf$k5e^+tfM+m<QftQ@pn-4z0GigG4e("3
^7P	an@OH`M3N<Ag{(pyzvVe4."F p@JV<esJLm@viQ `ZaX*x/yS>Z}S${;cdf<w#w3`v/}Ya?-}=b'j7/8O&D}LYG3#:.F`>8>sOot_xNyX7=wS! *%BkW_3+Y*)cixu@.IM6cBlbJ5$:q"cHhDq:Q<T%/0*hHW]Q\Ji!/	-u;D~f<xb`Obd*A^XL*,v.}U'Ng0CCd5)-7BpRq:d{{cEqX*pd4
=sfefY	_=>uxj*VrgN 9U/6K.TZ\u?dJ^wR!KIxqmTNa`8MfPyT|@J]8fZfKRCr3*G!!Xngg@_tHbl*3_=M1%1<K))>~aV!v?N*->)I1xg -e6Ii-@SYlg(;Ke]:2+5v\mcVX^+y:Rmuu9btp"PWtm7GAr=p@=}C ,R(2%;rbHCNA(T|gz-<D>_dVU?|P.KhVAP"m	g8zlynSoAszI^@?Y;z1"Ayzf!#Py(``eX)'D#o7is("ggL{Q*[wTuz7+w(> ]=,%!}lmf42-Q!Zi;9)Y]j*tIYy9H>Ug]:sw
@	A*7/Zt)F_qeOyFZoRcW|(|EQvN?r%Bc63TSl$1mHTbH	#	\ Tm"FyRh2;y hQS-MFMaI1!x_T${;T2[:[sD4Mc^.z'GP.*H
G?`b@@b25Pm"eu>#G]65wwEXINKMC2yERBtI`f3WQ;WR1>0~SpR,p#NZu+"<kq7A^{~%	FJ%A?	w6eanuYjj0P:FO/jhro	:1BZ+0p_rl$MWSlX|cOC40Q!4B`I~J#PT\4<dFV
jdk|e`y2<-4T/$.7
Hq7YyxRd;8{L&1uu/(d-W!/U";SoV	ghv7=ng<3,ti#wmO
"n@fL,\|A#lJ;"m-JGabAM%=VKM;|MN`vx,/zxr>GdfG"w^p9qfa!xH?K@ALaJ8d7
1gEWv?@HXzN6=^{/,@P@-j!%ipL^I=x7'vhJ{C8@w.&SMAty)_nPQi]tSiZ#;M<{)mYCVF5#5g}#^^z)bX!IOwKOJ-Uo^3_N,`|Ow}MrUS1Y4Nh\x({8M7m
P"@"JwOWV,Sf+%,0NuCb`{bmH cr(G=E'-J.EO6,'V~}IvcK?"h{WuQ:0bfAR;B?&A-F@2=\xDQ;0!{(g:u0Sq"r"U>R\ z,f8^U)LB$("cEsQ63CPo(8C/5K"SnVI 7%1HeYiX]~suTaEVrp4sV;0mJlL.g<sUbRe]64hJG <982i0+^Z-Wp;1II/9P
6~rn<s+beS0JNy6YP&g!uRm9t=sb"ag4+)$[Jy4:;<8W<.4Dy`cZ;BpNpl:w&s-gGX=91ywWP\Ql><4L3qaX0y]>lhC4A;vN.8YbZH}$eNIFJ/CE`BF37t4q\o66o*2~9L76;!SrV%8]#8I*m=ec\{UszSnR`5J+&lV_h1n:
IqTcaM_S,S	S}l=[yj8?yVru}Y`gRj?Hu'
jd0baU//~]ow
QUH+mAMnJtbKxOky(\gl3HSDoh}MgvZ;K%HS9r:}4Ei9sq@ftT)Y]hzB#FN?N>;Lvj?k]&_$w2#ujFajC|g!
LbdiFRa}ejCK_z4so[A!4LX-}]"~JZn2]T"G4e+i(;56N2s./p9y yP4ha%\z-Pox%u"g;(Mp@C~Og(2mR4~|2O#@wVKT*F^%}uJzcfh*83gQ-OFarp;n_[$
)Kl\
p:+{LE
5%l_0QDUo$5 t
?,WgoqC&dyme!baC@xWmUj)vbU}#?cbJ3L3|%S)A/r,KXCp{U9UXV7WR[-M+O`AG',K?L1kE}/SxUpg!}:^LF6LSLBxj(9SMmab^Y@=r@IWcMtPIx6DqV0F:j0 5
4/)Fm$RbwU	?*;<<!Tb/cPeh>7#QriQT0[EP2=`\.-.IMG$@{`#-o
_eA3G5N};2''Q%JdLZ8t>)X_9e Uw4P9{KR~QkVDAXhRRIjCL1=.6Mc&VIQa8FvdSy(l~GU@gq^%jl}m &Kbce@i^q>${dIJ8,2Gq`&'$,3<Kl3EV`F]TWnS (_BI98CFh_&i
`79:;n5GwM!A(]a*xU_`r2$	u$0o`0RJ}
(i!d>q;H$Zje,%Tg){\bIx18^:1V5-Y$.X!CN`sZT l`OmZE+aJuk=Dmb`Sn]x6\Ied.tZ$J8)K<fz,[xt<vA!S-Sai&Bua~rFO@-k$blF;|P[hE6L1XAxh{LV0v|om`x\Qj=!Q<e*SNnr.8DQkW*^kr0(8Ub=yQ59tm5';A{xF!8gI_9cK7"AzJM<)E^O=n'nYYq},(rS;zvbE.%uNU
ukY*,hoY<>{5Xl}T]O]?=FqETCl`=x	(vdyGhE!=%?Fea.;eZ=ymBw}5"?*-Z!3d(GNH7U/5KgU/qT@JIW7AOXu`t%#Zn}uRO*Nv]""5wIsK*!gEB%wA;d:KU=:]6;0?N|>qNq[ioY[Qe[An;L=D+Vly^37(0hDW:e57f8t(pUD6mp_+wku?Hu>^Vc'A[`%SR3U^ EFu"7<blb{~G8uUYEuOvdz[MUbJ4PfR'n({5S;G2UZO.F7fvHJw4?g>f!@>+wOCD4QTD6	QtrJ<'l]tgB0K;D{tE2M:d
+Ih+IKiI;c|QN\g;,L{B.N;@f@|vlu1vvv5,s<PXfW{1+,2\60.Bg2M%?nU@MDks9&fPtF|g@B
q$xP7Ls1<=2<X_>do$zSxci4Aj+s)}TdNznA|xQ6^8Fge)=5.dW^[V[`t45	j04A{ruT1*./|A[rQ@l'sk;Q7%E)uZyR|AJEY_&9PJ^\cHCAOg7EMJp/lfzQ3[/<"!V(Q<rX.-gD?0P;sH]]<A%>ebGyt%"](6DsEwki?	hY.	}+XZ6smX?CW4Ws6[p/qWv/m]cZ|:}3UKs}a#_RI'pUd
	GUS6@''^A@q_pEE>Fq &CBS0!])H8qbbQp{|XxT[@_CkHFJO7m[~@ueLmGQ3-tl,Xb/y9x5`JGfP&;Y~_!+f399B'F\Mf3-Zon.}"Ld/}:?`Dz(OpauTE5R`g	{5TQ<B>[RdDvA3":d8D6k[`aWja3]s;v+4WbMs"[x8oKR{s	lj-g>TRI3yW&t7}x_1vIJ'Z>Uzl<r^L4!.`k]X|'i(r8X)<5j5cA,jW8xU|8")-D/Pc{{Ir@)XFR%(EJA_$ BwE&2Mh{N:@,-O*mncB`Oj2@O`a_<f\J	gaL<yRgvGKZ=Wxy@^#L146:#+H:YV(Hy0/8t[Q.nP1pr_a6k}$&,O?k6S#ROR=K?q1z<hy#iw\*_*e0SF[E*5NB3`W^`h#uMd0RTij+_\BWGz:~1D/N28i5$G+?nKT7P-<pshy~Fv*!s=T1D9^DI1Lbh_{mZyz}WtqR)<y+e_zY>I%
<%|b"_SJ+@0kf]Zm%w9&g2O&jTz1vBP|`qESqZdN.&1,9SK-2}"@D<WCl UL/>^WY3
#`{yjQ>!j~jQH0)Ii-KN|Zj6[KY8#/ rO&^M:@qdi;V}JNvU4`@1yC		nin0O!1ZAfiF vZa4K_0abyg\|,+K.*FPO5$6}dX}[a?~^{+9|4#P"tHGn 7.5)I^=a93zd}'+5z6N7:bqeB=vQIw0TlaPKG|j*-_#UbVl4x#NEq&d]~V94j^4vkAF2y7T"@+<q1)5VotlC|gV27p6f ,E{[#&:hr34U6V3 s<5$rk!W^6vQyYMB/z`eXJm}p|aqw	H\[>ldOgO\lv04Iw-E8\DM:Zp%X@1A(r<eV-,aaLtmPx(<=z[Sa5~ZUPWgpU$!N)f]`xpkwz5ky>C^xTCQq$X-mZV#Is8Y
\#e#[Oyim^W"<`>sH7YIw:VlhKXuN=#V2b9"fHs"h0^^'3n=@xoQ"3bB|;7L4@8zr4`:"Xv^MAlH=&mjb_^tbU-Zc|VE?aJg,qDtf!Bi^#h?&R%MzP&0P#"h^O8rt' Idz4'c=*-i6SF.rDw.>AY[4A-3|{x$+9=<}4	=PmK=l|%9Mm|)rd!94o+CLglf1Y^Ht!^JEr $7S
ewiuCHX_\GHfhmWvwkB!gvb*x
ZuM9qj J`)!Kbh.=7fd<.o\zslWQcf*'n8{Z(ah|RL3vO5wDYIqVns1w!sQphO[t=*rQg'-GeQK^CAa*g@a}Q+R#KH<3LxD\I5r>j7%}n_pHd}lNe_*pxe#K5(Y/*F1eXF)BTeW-Nh /UW[M^J}+q!oL 8XLo.vE,jLG]@f_K[3	[f$;4O]0M+wP-4;UB@gxKA,_#1[w{Jft5zH1Na{uoMdzc*gz5cQLl>p/rI\Y#'kdOOkOANE*SM7dg$^kja6IUl G|\F&T}FZh9[SJJ]bo^q@\EXA^{\U_sxSFM2{?SL&M'	'Bjh^9GdGVvTX
?|{<{5f*|`|?,\G>M3^oC}[&|7VRBdo$R!}~l%}Lnd_5Lg]%9_;DgA_DR-M}Pt,itN0Jva3k|BOEiEByPv	uqUB\,'~7yqJ]M^k"MP=8mT7J3;\K/A~LkaJ"6A!,@1d@ab$((g/n@SQwzc`=^ G6Ho\^ey7LY>q \E=:BY_fp>F/i'0s"l%Xb51wg|K1_Xq&F#k	U!z-g|LdyA}S;1+xgA&bP8K{MaQ9/UN-)55--o_*:bb>1dLeU-,YS(-k2aCE.j P4+,E)	ON?5kxnARjX>.Pj''0NgMf!jOuDiB7!tMY	^M5+QlIt~t[fpQ$*9f5:|L_*N$/J1Ec;uhE8DseDyC35imu,|h0+0[?#W
	7oA{r?14op|5*U "U62[']{	u'a.iX,l'ofc;3rG.xU:0yk_Bh}|GpQVfa2t/u57or&{vwmi(m)je`)!\m,)3U^GYo906I ;?zVuY0BBA#w#zQo8Q1hFgRw:rcChG6|4rj(')sC]T)|l*c`oe(B~PF>>c.pzE-bu9Pg\+VphllwR9=+A&zb5*HWJx^X9 \;R{c|i:)$I:6jIL1a\6jh(T|X'q[F*Z!JYz:~hX%JU_(^8Wx[NO_R2Lt!hz@tl @Y648-styoISJ"Nd>s3Npw2!)rlCy3$?U'X_$KboGQ*BWfb^VAz>hWDOnHAnmeL}DCyi.Tp(qy&*4haUz$+rx7P`tOqJ;geZ7+ 42<b
Wr 5J3{H3:gIgu+|">.W<)>Qr6iAp'${hVm&L}Q(%&sW+e3<Qz/EA1xkHN=BrXLsBon75IY?9LHz6<PD[8HP]^y)|zU^Q?TYWJQx0RI4|4bp}o8P25tW-aCrz[-Q&Ek})@C.1E4C/PNp:km$1%cQ0yy9_?gmWkwv'	)W*R[lFR4kp_CC$R\fxj~_	b3-OnA#s9oZWll|j:GSuWF['nZ5^fgjEwK+>-om*f2D-`?oRKEAgjvl?%V:{n;1f(&@V\1H#9Sex}#kt{.d77&{TrW\	?2?w'ElDM_|:8)^nHDNhC)4Ji 2>gVEb4nDDalu(5N]d+%-EL&.8Lz_/S$NAM>)NZ"j@g!\\NV-<99C#r">$6?aATvx@_e
(rypHsfU#+K,k">t-!5AoX|=
Y\3dCd,).gQ)<#EB\lPBVq~rn=H1mXRdN%At0spz2cQz7'hE!poO3x<YP~L-gi)P}I%XH_t(tA[i^}%%*T$=2MSNss-LDn/O	Q=S`+/RN]J3Ek}_<1w%8W:!io
86tAN]*;D n~/Zq.SE+=FQ~v)gTR@_W}0n;x29Dz.[j?=rwmUQ0j	=cBSPz3UT^jxLq_w'a3aCDrh(8#yr%d.]H'-qqx6BeVIn^2?nr%^#&]sVO0ya`vR>>L`EW?Cls
abpL\BIns$Or:M'0fV3Sr4|K4voNjE!YQ2ajV?r(?nfp03Xl+kR+uJjxUD]s+>w40qyOFZpK7zgu~^
/.p=o~{g|RJ4Y*2@jp&p$zhzr)%b}Bl~Mc
<n]\iHnRpNqJL3#U\#<Ray$&H/G(eaMlnG7(H#4'%kGx%|U1\s&Y((e2jowk[	fi})oGoZgx<gt;kDlpA!PIZ1^:dL`sC	#alFoA".Mk@qgl=qLl5&B62+!a UVIJ\>!x{.u}-Gas8?{Fc'$5^Kl%aQ,zT
vFgpcTU{'f+B(p_gq<RG#Z*cw[0Tdxs6@X%iGQrgy7<jS`:*#3<z)hyi(e0t_{ugV^9
Dv/4gbo[bq#XM=TyI81vdi"7l-H.J\Qoe?<)RHGC-P|GWVQd|}]@C,S<&gmG$\(Y:h
`D@V[DLI,L,@PzkfUBC"XrdZ5]um2WBOM!1`tG158q\-T{`AKRU+,gx7!P=	@S]P",u	5duRE
=h&v)vi-B=~FQpNWbj(,dx (cqs&o@%Cn'!H{!,^|Y?ZiyU4:xH!	EZpsRT.k?
hVS4XA3Th}sEX.26o^xxymC(BadN<s[#,5k*.
eO,,f#Q#:sUc&1H[k:a{du
uj7(k|a]r"-%0%GV'3jPk(F^-($a^72)EBF}.rf;4ytv%-	-nl`)DT[J/W<tE(dXy_=<cR_y2EJb&w6t8C{7umPme'js'[
,CXCSap%5>j6Xkj|@==+)8QJ5M+d}4D'&Q7}31/X$MR"jvE+&yj|Kr(5`mQ=3(Fc7`Mrx_Of*uJkW;b.+Q+VR*g;BPq#V{)
c }_\IR.rT`:i(YW$W`f-Fk#?@.)d7`%r-dk<
u6#2@LEHak;Bj6KI*KzCh]Hxd[]E\'1~LdEKhrduTqth?^2\(gIlb	n{qlHkWvBy2aJc*5M>-ae#Q'4|bv-AFw$nI&oP5a*ZTWGR,rIUkX`"h	jtv\pNDm~;;;@2 wdeP?p1nc7%e_Akk(QZ!^^wr=0$'xm%cg6<fqlEC)q|HPk@*[SRfm`EnLnA :>,[(k:7iHbi0ZC>|n4l<PYCeVO}%HB[+yXzOja2$`i[esF~J+c1p;j,isW*obJKJPjw]p)mY^P	0S"rhi)pDGi/4jf!iat^7%GNw1,<vl[*&DVEUh*bo2mm-/=2x,=	,'bd"SEYQsqAm5~'	K)_UXta6-^Oj3,x44m'U(Rym5\RF/[bA6F3W$B."NNY}l3f_R5=pn%wb6n$he?h^#Q9f]}JW8oGdWEerB~^0_qR uz\a[ah{v@<Q(P$zD%NJ6[	dd+&q|X<^+OAr^aZ591ub!@gy}x9VW=A'\
r;J{E!RxVhH^F!IxM&!TlN~6LHD'KNvA9^+gk{"0x5vA<fb(yCc/PHfJ&FSU2J%P>2|`#eq_uXC!9#+^]L)S|obT.")lP<^2/**-4aOQ'qxn5#?+K}:jE_
!SMVeqNkNIf@d3&Gv\3C!c|kb)[7BnAHbd+m./ qGa
ERmW1 FvA\p':U(L9<U\,}FiS(]*4T.pNp'BLU!NvW<MpO#Tnw>tVv^vR.p^t{#d_JBwij?%Bjs5?bkby4jhT;x&oUpXfPN!A>bA9qa,Mv65S*^=93Gu-}o0B~RA4B}3)5+oSp;TNPC}^ji:K>O;t`">_AMXF??p(%]5bBShXx5T^d;3:;\S"MJ$c2;|66}bIfr@jVg_hTIK?d[ig"!E<C1{#^	akP9e.
9%	U/AF1ahZTD(0)}l"X,p>z8&zDy>-y~85`7[H#dJ*Hmk8mNkOP6:ZTUg8x8et$K]nW*lq_C;NK	ZU}z"MsU,~^al.Hb43z,+uARR5\u#'-QbX+gW6#wVw<_yZI1-b=Qgmfr?biT|t@D;e<*!iF>)"KNnN)VcW,^MG>":wa'wk[mYz]\|i5"P^bz8g9-CVy&lG?^EkQ~G2yExq_XY3qUa4f	b]s^R:OpVf9R
2l{=1J<O=$'>o0 M>J~zRgYX\HIw5@l-XY*P@J	`69oYA5U=q~wy2v"v^$+*`eQZ}5{~FTMQ.y 6Ty	%Fol?$ZzZ%w^;4y;eRJAJ\Egs5hOu*/\Ix}_McTdf2Q
.Uy.pj%|dGdQnQHo[j#p5w|w6w7^lKkD8,q]!r>[vJC)dnti%)7}mB+GpNLy(%;%'53:)%vQ_jr9+=X4 ,U*HCRfY**U{\	Nq[88+c\1ks!IOJf% k4ct+ZyOLc\G*"W^_Q;D/Y&3gD,^/4Ppe>K.6XPz; G(0SEM[b ~c_hLb^;6VB=q\25a"MuPu:QLFXX:ZjZ!r7uU/%<B}u;U52f]
=Dz ,MAx>/U,bV.~KHAm%Kw!u\TElYb{!UiKQ&(vn|Kkdi+3;r1~MM+f`Z6|N%t:8NI4Z.1?Isl"yxxy|A~G!!WnhK"@Cs;vupTl:Tt7}^I)bg8%]~T'G;m za[IN5k*^GKw]Sb?.}GV3LF2l>UIwrZNaG>+xc(Q=z$<"o 2LZ&E 3nJ?{9;%#yZ4VncyGT%&	m/DK%AT*edN3O~2eR3/0+$0aIrc8fG^JL	3u[|xv	6taOwn3v8O'ZO+2Jr/n{-IRki84}A(.-q-U3?|@A.VlWh KhdQecbr)%nhB_|d;8U}!7U-e=	*=_j<8'Je'r{a'+uYL_ippe,s|Bv`<^al&:Cz;T3YNk9sEPn-Z,k961FmkJ,a0#9;u0)8W}K,IyYSJU0IhpHk)uvtdh92xru<I'#<lz@JD#'xWe#i#x"CZ:TiKClkJb._pGlMmFmh"	:5sL (l>D4	2s;Q.F^tU8hW}B0ZWgD$Vz&{t*/{j M[`C8L6fxBDjW:S|ns^"@wL< YYHop3.'NHS8*[hA;DgulpgaOHYD-x!ib=&)0P|{+3t?~;L	;l1[Bs:7EnigviG/-mc%9c@>%fvBRq6E)0#Q"bX:2v>P3O_n(GcVDUa,{B5_o={f}$II#R(k9-&gX=^LX@u4l%!F(%-f7=Poz;[<
0>H|\'}YYG^4 R0Brcz!%=ct9.<\NMW=~Q{pOIO`LY!I;sw'?lqNO$ ?>?PZsWy{	UpdH?z@azno*DY{
Y3U/DiU)Lq[cq1~4/))*DvE`GRi]ph'@$h*$20!);#_1)52/h!Jx0F`Px2yk;sM7$R0}B6Nu+_@Z-Lo=sUUDvQq4{aK+w>"5e<w~)_%].;lw-a~f$,Ek*9.}#*,q}YL'#\!j:&;/Sc|!PVsH&\V$N_C_XZD*pJ]k2-#XSN	!wZ}9*O62'/=VG'u#0:4}|&@hP-U
pMgPO0|s'JU8-c2IC>*'CGN}		c}"Jm9QWLs(6FG0UeVr&?nv9E?j(tN:QtjLYpaM }# -\K:||w(>B{{UzPGC\P_m*WU_UcW:q]>\3y@]U#OsujlT$:hc]WT%QvC9m3v^algH6-#V2"m{cpy`:|'n&9`PcS.Lds+Os*?yX=1$!I.d@c[S*FN{^Y/alooRt\mD3Bmtq/O\;B@wiTGSP&qQ]4SWi#8nul-*NEJAoPJC,(K/||YnOgY,Xko?",!oVz6'}&AV|>|I%dGk43I*MO"+yGt>{rH	xx]IE=7%w{f:{9WJm+e~ vP|PXZS#oq$UfpU:3RGSm<)BMa}NURBQR`t>q3s6M0kWe4jZrPeEaSY]58qXrJ#!"E7&/X2*Z$ G"+{~{787mH5But'>2a.Ct`ByG,MD>7J/KOu$ {fP+g	=7aJV4YN/	eM"5uTVwan	G3^@sS|<tA2LAmId'4El+;hV/?Hx+-|l9r\w-~d6Q6ivxd[Mp/mguT5F:>7-6|+z1Y4a--G6RQ3HlQM+JoM-2s:NO;p:2&x"Cnj`;
HmpkR77YWzf&qEa:u2(ry{r^XO!e*"/[N+e9I_}%UF1eBwH<p.)y'W}18F/X={go"l9=%0vs_w=xjtk_2-TRI`UQT A7j-r	U(%xPQSl
A\QoYt6F(	V_tuUl[1.;/PIY.n<4ozI(:1B{_@N-K%?I$Iu_cZ;M)?J!GF5IF(8QC{s'Wq]6bgG1+CpS74:vcsN\a||+(?3@]TYnwH9xfQm`6\1$`*u5Z:dxByEW."g:Ep)SK[:-v @y$%Y"
mhC4~tv!Yt,DFzd.SExE3|8[6Aj1YWpH/4o]I@3sKIL9]6yxhufkc2Lc\3e"/io,4^4HytU9i?%Kd]jY."$:Jp^
k;W)DDM1hp:f	=qq(xV8T<;
<=ed7!7*)?#Yne1G5Wn]QRPOu6`D-wa^lbS@@b~hLu|l1--GB,kbL(-/`a*-LTpXlin@;^l.E	YT%tRX1t,- &nan=y$9FneV<cDwY>_^.{tdrRaI*{{^3wdo~PZ54x}I+)[v@>TiQ=--$<x.h6_!NzK>	iO]@2$]UuzSF"L|UI/*=7E;0aJZ(bJ'{r0=f&_Xa}G~Lch+w]PO\G,uRa>%
$-Q"egHKe7aMw"2{FYtN/t8SgV`Bxvq_:'<c-ACpnh,hA){kNQ#87<dnjIv?+TvHUQ;'BD*]6#K7md-LYqi
tJn:<4cOCQhjO" [)r:tuFc{hu?fGdPKR'p8ATda_FidYTdwf> &s0FfkN0DHoqEqv{eNzQgFfF"KluGqiC}(<h3EXM8"X8p!)b?j]}mL3I+ }0O;}K:60+euy,[RU4fw(U3Pq'wrU2m6KY5`-27g^2dXzux<*o@]b,Z*|)_T|]tlc8'b -xa$@r@m>fxbY>tx6j}6p.^i_2UeV"6dpfyB0[n}>t|t"#	E\U7YyyO|sggSc7@J?;'LX|=-x]%i3AL\-$3oaK[_LyLTjF410\vq&-!kG8.wg-&=@(I\<P]-XgwVm oC+E/+P"muOm;_}mW=1}'rL(h#fOx+;BJyz>TPb5cF5WSnNb^tZ\y|$dU:oIE76^xLJ$w :Ri.5u7&VDn^mR}#	C|3LT~"p0+g+5e:Oz=#!'bf( [}2Q;~5hr&?Nq4%j,	vtU_b/Jx=	|(@*]C;_%D!n{k#H</xs+Ay+0m0[T'bf.6gPMu?P1/_SB8S!3L]&Bf)P7MLka
3y*<r<mXE#D<uVRK7u?Y781hCw%js(E`)3CvbDRJj|?1SWZ$R;:kj*GotYy6G$Gw%"<@f=NTifM$H
=$]q|b&i<V)=6S_4'i<(_KxvEPi\O:
%e2qtp9.qpf[fS31sBn#[Hrw<yFq!&h1IFhDWjb`PKSeFQt?Y3{.!WiVh"=?z,nJ)8y)K]cJfEZ\G,	lnL(p (T"&`dgtZl`.*/\!&Sf"&z/k;xAK697}4`+y,	$YO51(ol@uuFVa^F7,+^T><Sl9(iY0*A `W"%{7{bMc|S_V,
_G.eK7AGgYF-g7-XD.E-K.7[lcbQP=x ,#-u\T2MYi:t(SC_M)\^ #&T![#t,hZxeoq~u-(77fRz9W!:|'<~F-haA
#I2'3_}*D>)<voB.QNl@f4&m1S\edcOlk!]T[;?B*\vNMS@iGu	"b~<CHmN5DK|*:o3b*cWl{#_5Ux**?V\K>j,<~3.y{i'n&x3ty w>miIIe^ErGIa>=kPh5M9qEGfo\Iw/}#^PH|Rl	-w}#VW3fQXJ0;UI]+Kt ,5>lp2#krQ.TJfv.i.zTcg@]5s]^J%TT!5eVMpI0b!srFPtb>ccAQr?/ja}Oc:u_,~c)N9 jS<8A5F/7u?F|>M^nEKV |}
hP#Zb(Zm*h-z}K*;Cp,(|GAKtav\ase`&`;butWIIlGU`y~m*E/N$!i3cX7'n5$7y \&<7K^-G}h?K]ww	pB9,9,PYl'#xK-B9WY9>ZQsy5fy]Ry_h|W)2C{5'~'zQOfvNP	O(u:\">&:U
$64I]&L/ZGO_~-<Y+ ~0|op0u(55U_2w^lC|cKVR-iF:, =Ih:.sX=2L`R(lVdJs.z
}39_2b*S3P3fD"(IK>2^.5Ye`k)8hMZAVQIJH;,?;`]U[c$lj!,IR#qnH[`Hi'm"^o2%aB{.#&7$'(/
EQ3@=uuIKba-6Mv>3q8'/F2xxr/ScVQ^	f 7+"F
(iSN5w}}0'?V@6%p&@mOW+b9Sr4e\\Q`>Y=si+JQ0s4hOA
qiyH5^8@UFJBZwIrEwy3Hey,E	+5nR[bY)G2=%GQf$GFq !K=BWTe/W(|P1H}+kf]#B]"/	/\$y7@jsT;/gq"S4!k(CY`-|H-8d\>L@,-y&7b.9II;Ed/(z=!FrX<@oT0\TY)v-6}Y\AG3&*llz{[tTS)Lo}x(I}BfX_J:G&AwJo0
&EBlF~0WJ2\DPO}i14A[r|CGO!N@eEP4CG?HS0}*;Cw4-z_azwO=^UHS(s0s%5)9]dv-4b~ Goun_EHGcI2#[60J
J=+EsoH_CW7zIn<PY3~"rcDbDX	&yzGf^JJ[*lSqrt%BX"v[bPj]_QUM4x"V[*2GVsFA]glKY?kx~aZe<#dMp=
d_	]@=)\;#Cy^",(FI6$;rN'jG$@ vTfa$)EnM t/Mk8TGFy5UxuYDD-,~VHXPT;g|u?fY;AP7vZVKZ,r<8Fo?D#En/.]ql$q|	7MStym(Xq]=_K=7)Qm/llIE-36Gp@dTBH?5QKd'">WS3rpK<3Fvnz#nqOx6%{;qt5X]P3x?f?w#Jq4jO,=$A5p4>MO,/m,7
J`aD?Cbuo)I~SG^}r`=l]lsuK/h	
e?B5:Wm8axzI;/+kPfL.#udDW:<&",U|~AO''\"k^8bDg\qkQK.xE3Y6jb^_r8tx^k{u^7#KX|"tb0Y3>bUz"H?oQ88$%^Cd=I-T\__yc7\6LkoudE@vD'tgs6y
b/" .yFdj, luidoK26"Wf>d$p}+zx02GXA~u
[G-h/xT5zl.#N["y:<}#%]+FKIQ`r3t6X	U]a{^+#QL'}9R<sg72{,B.~{v'
'f$A^U)Hr{D_DRD,AcmP-Pd5;>oR/J3T=vV|brys5H=h!Lbgch(>/	1%li,A,x8=MpDiW48e5X`nsz1v)XUJTY'IiMXjN|X7zv:r	a|MR<X?%-jCPzPND@wIK5@E2}jCJMVc}maru
*sONzAPGD}yr9$6
wXNV\Ul8 gG4w@j(]gFW0XKSh\>#9k6!<Ic~>:OyqWNYt)FWY%	Q71UUdC0WTXFF4&gp
?q?p+4U{[AL@l$l60T#BRRjW`{D\h[Qt9R
A#},'m[TJ:~F9xpy3fL+i~Y{yAdgy=)m|xGi%YQN_);RKU
7bM5t{*I#;_G:IaA^<;=J/?u@Uen[:*aN[h3>6
 F6:FiYOT%]?@B3/ym!6T[#.t0A
e,$Ug%AY>mWjs!NM(.BM ,H|4`,uqkUMTz^R+xFV75FlmQv`Wp2G~K@\q	=g4$y%q&[>9zCVLhADqpT[+"QFh9^_$({2+L ?^,C-7ut)-kw\&5N<>2Iqz%4Jp\toJ1r*ZvA0EBSH#umVVp<;
Zo=Az}b 4hMMk'@v?A>tk&NG,v+SsT!vQ(Fr;3g::nB]6aPD;ut|!a0s-fh*+7ok|3|g>R
g+y!b!K)/&`t26tUL].n)\t+J\".58Jp&Z'k
F3qjM-;3EsMV9.oF)UMT""uOwk
S,@tBzCP2>jWaMEXY>7w*)tM/oiAiNVQ<q2UhPRDaFj\H^\nEb+8[/AP\bl)ae5y'	[EyR.O(0X`|Ude8p}tZ~K|vk'k4VKBO$H#QcaI1n=eA.@]:e=k.^<V;g"h|<Tc-y[:ElT7a8z#S*vn~u	^QlL,JxZ2a8a(+!"?G
aGlVso_@|^]U+N0cRLUEl-3N=@UtP UW-y'0$OvQb~oSp$'0Ixh#I@X{	t:hv$(F-)OuM)k(t'RKqY*#3{7+BfVD8O/RpW2K gYv!;jst]DT/+|"/{cl}:_f]S\MpK1EMFDG/.=7dQGvH5u
P:^fA{pVG"]7zh3*(]$]|/{g}z>I2y$Js6eJ&hKzw=fXbf-h	_A@8jOYbjNZL[xT3Iv5B}W42!LcV|&|[
D8l\RIA0ff7e&l8`(usGo`~6X;]tG2I8odFRcV3!N/Dm*?!fGcN$*1)u;8t*]hwC@u`k,KbaLYh<zD_"xv8KGi!*>Jqo!agHw4 Vehl+P<Mql"A5Jv(+1TS:$.oa8>
	R_!1 y|(tH-^OAu>sT}s'[=:7ri([f%24<sj/h^)@42F_z&/!W?I2RU)#u =4VO
pb"sp9WO/tC/#	2fH/4Fc>ZN!	Qz&NLu.dl(vU50#CFvS1iG`JQ:gK\1MGgnG$x(1gTWgd?T/Njp(ytZot*on|uiH;7IQY+M[5QIx-p~ib2
<gxx;8{2LtAv-W`-7O+0z'LOpy(^P!'cVI s=qCVO(|)?:'g`yR<{q,RNC,vW]8bA51z.*1`kL?N=iH/=2Eq
1hA?"swrdHz1Ho$1CE>02lZ}sna~q!qfmQ=!7vh
 ~JX^Sl\w,>%sG4>r'{ G.TCq|by #db.E<Qx;UJ9n$/:y2YCw0;B(BEX/2  b|a`K1dAr$p<e`"7u0kBo: hR.o;Q`I0avy74f13<NQ;C]c:.\^;-62C/+^ZmvD&sz0h|[<3/V5]o9dx{L<<FHM`aNs:
!a.vyLj` a\=U~XW|oHX3Z(Xe)3W!Yq}#Tax^94h~'yAkb7j__X<t5V94,PAEgF/Q@~43Od^33zy{62~81d^$pJFaYLd??Y3G>~BwM??lbrKDp{KW$!]nsU*!wOfAb_(G@0f[}a;cw!JuJ.wP=$}3/eipI<zy=-4as|)Np'`*,;CZ
iB>'W>iD:'Qyq*VuOrvT'4mMMk9Co3K9lowS40ykgc>3!(sEJ:^yn9d^?a1q)G	l
n^@>\[yRFI8%ZFB,B~UjRU;H^k'Zb;<!01=sSnC<@g:Em-.1";H.E+8 uUh]`5b9)Vw$aSjj]/Q2kLfL-"VovdCQXk*jkDvTn,v<W.'RQi17"k5_;{f,nw_#w(/iuxhmrZ	!:.{))n2	pa3Q!8u:k8$ErgubD%1eh$0nxAkOE|4%:'n{!"D"<ioN
"@J!}N>HQ=k(jt_g
^[-~,HH4>?=H$1>S<&'8'.59f0W/d*D-;CmRm' mPetuw#9.n\$
(%MPE[YWyX
udOf=| iB3f~NX#'F3lTUi6sxBuU	1	9DSv'WKl^lm&e{I.N/Rsh9e4lEFkXk%8dPxrD:CLi;!#1EKv,BwX<GlYh}c]0!]_pS`"c"VmSOed:>S@f QS8Ql''9R(OD:~WAj-<L$I/#I73 )ER5s}{9+D	piy?F]jR|v|w6q.uCY+y&5X_P(Pk5{dXg@Cd!qQ('KlhBZ3/
9+H0	.|Jh=+s&Woom4=Kp]$YYVTA\+n\C},q@Br<%-X5+cvX0GP$+Ut8v;EGZA\fB\e8=0+pJq%?43(O9gV@Zx@"/	DWd)gLJj["KEcqYb{+m9'J:3|&W#.E1/.}5d%5_$SDNRj$Zk)\z-rKB6O$/).$YnJ"t!BD4ysFa=H:_2ft[~o7aasZ9W> >@UedOVJ+Q(%_|5IB$htQfSm=[b/:MCx*ZriSCsgebg"iq+;Z(L<gYt`;)#~F/!
	_"&j#8,rAbZV7z;*kTK+'Em=?'PMb^Qh<=@O#(R'k42'~iUK0##m[AK29R$wHk=0uiTA tx~
K<|hVGf'
~pA67kP2S}%Uzcs[P4HM~xk).H3jlC)iSvaM!hU@q7:I+fT'\O|"<X"7,TL@W'j(Q"e4rOCn^0Rj#Z#dOT4ZmD>@"LEfG8:<G3OD5U8>iQlR5|oQs01	I0%(3_]s*6<.9kHT4e&yIT>Wm
FZ]k`$OV+#X]sH|cG%c4e]yz
+`kC_GS	N$(^pU9N"9,f3Gk}QLs>3IH5ke!C,C=ZyYdmcv<k|(gn||P-Yk$jik~7`}^Zxbs&pE9^$)KPUH &-)Xu>$aAVYR03:DM`81>,sI;U'80B:Jx\tt;v&?iv5Y=-DJD4$R@e0{|YNi'K:48fJR=OX~uj40LqPk7+mGy/n+r7zLjrg%tvlsbc'<>hR8^ vQmV$3F#QSu7L0#R0SBB{I1ejI\H<t2coi,e$|D<V<WxAyz{>E<%sxO)=^`/WCrzQqjh	%L?gM
Jne*XM(m2kc!v`47(kqet!:).KQTdZd{<z7sHt#]HS+(;0&1-X$:Vhc24Nxa7a[OUd$|iW8a2,Em(hF9JW0GPdiE80$-3*q&kh"V5$+<8H>v0u{Y9N8wAz6?ty&S!@TjFjr}`s0vOJ/XG|a{>	F95x+DIU0D$=.xm_:@#Jbyyo:y.thKQZ#^xFz.z%?m6<h|<{Bo%I/!h%KBH7(QH&PfS7,iuM3C

O=<h\J^+cUpVfUi[CKbA_#YmD3;2?cg.%\p:-m3bwgN19Vu!v\Aj"%z,|#UG>)P 'p~>9g@, t3PUe/?*y0?c0lBsgvIb?T/]?~VhK6&s\({BJ?9|}"Sqj=RK-]yO>3g1zeM0cfBg%~$/P80ad>4%<VgMQa[pz
h~cd(/NAZ9 ,FV 'gm,4IaDx'&Fsd'7b!14NXrhZjvKQK;4yWsE1Qq/?b`h-{jJvuN[?n9%D\\!Ae|$KR*BNAey'lCM
02vW5m@6&/&"p:UQ^E
lYnk	+ubO=c/%8goF*b9lt#>7mE	:Tv8<]o5j4X@P~7}9x?/(T#yXabw,1h+b1X<hm- ![ng=bpT}+aSL1#L*{c@-Ah*vr;;;KZopVLv;pYpIV}~WYA/CWt f%__nY1nT`YZI6W3y*eJqB"24y#QfykQ|VKEe[#Flfb'Py1uBKD9s^"icF$'tpIGQ5zkG
Lkt39S>VNY|`WhRbe)Xia4_hp%RvLOwS[hSzYs?E;$_F3dBmj;e\hmQ(>w;y9r2IgiNEcm#~(@F\u|wh?E:N_L*]2\Q&=4+_E[`pXTEV	R$fi*gU6b~BnOO}]a3Z/VJ$$?86)>[B7@P+k~2jJE	c?vZi*os=zRQ;~x;5FTE	O|O/!SH1B!:i*`I*`CfU
KxN|K;QUs=m6L$[=C2RZ-*$8^"j{tY	>sDrz[TW#"8z1iC_HCQd-FTME>Ju6=	2A0+^[h3& c=4=,,]DS5zRYMe]kp?eWo0!i=d.C2R$/(l?(d+/!iSdZ.CAf mT17JL66b{Q&"Hq=ZYiEwMaR/H5F/ezRZa:'DI@An^A#?UXq(mAw{WR81wf7R<!U}Ffd #KV~JCX	;p<xuHm1od(3)E5/h*[DWl{6+0<7QmEoE2{+Kg	}t ad,i_>a<-6/VY6%omI55PZ|drSuP(cMd+CXhDZ tWr2Kb) 6y eZY)E:~-$ 5j{rY%n"t;APB&-q*><XC-~3kiI@LCXUF>b9w	O"Z2emX}`V;WJJu((A+(3W3Ynw/_W!9Jz(7IQ"kqSv7{Mo0+.)%c'72<RJgw+:K0G.I9
Ep
A_9egLGo&1UagdDTr*By`-l&wN}wBEQ~$VzoV`eu|\P8YdoqKbS!9	FB1Ac*|iU>'AISr4]hU15?su`e15E$0>y16FM4j(' l;d#hcF ]L,/['%3;kGw	l\];)FYD"Wlo(}4M	D'LD8YSzI0[5Xn	]56>0GwbAXHfz5x;{LK;_YniP)*v+{=58fu7:G$kfIvYFW|-Q+!`"Mlfz{`\s=MjszQgVg-@+hh:J4[ac>_xevnmuI{u4*8Cqdvt9'HNdwgoM"@G@dcRMYFj6xx=Gcdzr"VGj>ryMN9;<DCo+xv+<,Ci$QC*spIy"U%@#xsvcvv%d"}Zj~x8r&XY3BCU& qw<{:0lp>.jdd0?z~NP_\V=ON7|PB[5&TnC{ZQ%A h]V^=f@!7)WjDg<%Tk2@7XGQBRJ)4K_GC\r%t9#e~MT3}NY>%H}_R5RDZu=,EDxAUDe}J7|=YqhmYSJ_"m]Yx<efn
Z^/sA:mc,`.Uw:LG]( $@hiuJ9>0sY|mPUf$2j{U#[vQK_=5}-i'<9\Tif=,]`VU;I6)d
[J?y79Yvw1~LYeG,U'4
z'x0(}JzOe1mCDN\DkTP# E)%5pnNPSvBBeT*D	45{Z'$J%+zj0AKt;T#-jRx*:XxFXzT;UIT(`H_=`oMSnG#]_t4D;CNU	"RU8Q{~$}xg =sH7!]Ef$7e8@)oi'D\lStK`9@Fb'}:TULMx
nqGI 09s`MEe"-BTLalk-=;!QS_9`aTU~:C>bDRK~_}	haI=*k$sV.R-gLFwbnS	s8H$Ro.QerW[\@O
;$4VuHm5F	xxQbCOKk&?*m3\0ec`5hi|)RWNX$,B:.k>uDSIozaw@p2w##J16o=+WufZRmA">iwuy5"f'D#i]aVwa *[n.k0Q)NA{vZa,Hrk0R<xU^J1$Zn&.IJ V84).Ew6(i5?pby;/3P/^>sg'y]_,L349QvJX-6o6Jtk&lF|~z9_wtD%I_<K>w_~e|-@MLI&4s'[4}]~O,0%=(%hk"b	-qauJT	rL6"!&QlF$lgDIz,uC	^P`FmnN^W7'(5*TFt9@,K:@@[/}>lo|kk	qj{;	vFHbVWr,|K4f"-DzGg'e$k8m8PT]2{8rB-yx1)T#L2bU*R]4T984@U5C,*D~7}B#.#vtu'ok;16
J4|kaJPX`CL\^ZuAA)3`tbYSPqR?Rga#-FE%Eo\s8a_Vp;0Hk1m49EmCUk#A^2W#]jy>/dwN&U&b*-1q|lzi`ZQ;/m[Go?Z^|]ZlSycI@B!=DN}	O4[a8_W_)LezoF<mb3qY{
&I:@@aKL3QzhrB(jPoC/`Ut}4nL~	R7d5'F0Yjf`iOLf+(fIozB_Y'@1{<z7<c,-O35RaeF,qnRq"sTCR[[C8oVM&lbMC-55xmkuuAN@5-^X'|k<=o%(8~0|gT1AdrF ASuY?1/]I$cK?;Ip@EMQL|'1vD$>Ai8h&4G[8qa@`kg"K_\.46cKb2'~Z{Q?rkvW>T7Iw53)E_$+sznMZJM-eN(#^c<O}l<i1Y5B5f[z.F@LlJLg:IbEYzznS[|9j1rQKW:RF3zNrNyZ-?)?.UGBfs)pE\H%DX%UHq7q+	C}E7lFezQ~49TDDP&}M!W&CBOLy6y=A9Eof 1V?/asn>dJ]8xQ>gUmCI5Idu|BkQ$/Tx2AJ(L#${2l)	>;Ng|{vX]E0yBzv_(,?EWo%-yACQyILcsi3MPNByglrVIVD1E:'nr3@N{qoJ7_.FmE*Lm$HV;}.;X3XM`P{QAI:Zg=p7FX&:Te^#\}wJkRa/hi/9SSTo0[g\5Gn%]:[e\HRgcrVi	!f_138"=t4='"#sj.9EJe	E,f>F;Dsl"v1xwl*0Bb3t47XAA&[ B=z$NB?(@/]^rdu}d^h ?LF1G@C/szqaj"/Q2w9B=L2=3J_s::[q|p79NVi_D8hTPOM+eh/J(|H5/T? %i'g 0wY
xIMY4_h0iM[+l_Hnk=_![m+ZCw*OQkLa$dm5X\Sj	qs>~b:x5S_cX5Dr%{A
2mU/*+%dOq{Cl0q.rNBv}]oGi(S?Mu|9@8DPI]Thvn|'bV]& $GmVs';wk!`NpN~dfL1T~X#1D
9?VAZ+VUT//m8X
P#ktZ$,G=<p%EL!ot% \LT)( ]Npf!_@;J(IWq\72mo\"[RF:V'''R4$s2Q\yVZi%"D@It#;rxS4K6To1za/Q-L8r3QeK{J5bI[ducp87i3t.Djn^G=>h	PIv.	$XAW PtdWSa{)FM;'8r|B_]<J)'oM>rK",*}&GpA{Q1(pk?7LM5UTr?h\IPrL(h^4<~zNB"sF;OXyG)xZq,eyiy2g7>*;j}Xd"YF*<H7Y|Q99JJ",*l2vNpxA"@W0x8V&']Z$b&Rk&R|Rb91H%6}mo%KgRS@n:=fF6QQZL&bw!QkMm>B8Hgiv!Ry\o?Mbh$MUbM9Qx"#F^msb){XUoaGIW:M`]+vMLlhx*hfI<+TQ)--t@aJ^B?,"fkB!3WP<I\BBu"^iL>D"dipf 0uH]`N,yx21C
Tj'k2<L@Y%mqBUmbb^ON'P/,Q_;M40sj)z-+P
9sevz1]pkz#VdA"pBMsUV4VjPn=.jy(f29K3u1=G8K?YQ\`l A+p|ng}E7Y:1'%kO`=Rfykv/GuL=\tO(8=Tm1*PQD f)|0fRgg~}eq_gZcG9$m(x"`z**9,QFIq''Z&;=$\UL~JOj?BB`w5<Mwe\aNs7rR<moAcNyON:'Ca
Gl>/VG
}*:L,EQu:9Pgz?\BPc>=NHmUn;^]2qsFr&;S@T+aJ&%VKJ8KLq|pyU_o2z
92PKH!4N+1V*9X^W{0fc"Vz/qMm$it_Z3IeB.&8f6DY}+V?Tx>4Woi@#]jmV>|.		;/rR&`S>OF9p5~2wjo& ?=bo4qh]$Xnb"k{S;._b*2Da"Jbq!>PE No<5&Ec.n@vKahE08ji+y	FrB2Hsu02] ,hw\ppzXlh\"eVY[T
$$NjY|u_+0`%*9RFirK>+
Yf>j5`G_qZWJ;b*jht~=7QU.ml2a^=Rm1OIt1"=Zr%y]3<bvKJRY[)f2:%@s)gv^6=?w<t&R,
\s`Q+7`8sjta>N
<M[{8< Q+cRc	cS&:Wr4D>"OC:gokcOMNa>#I?9\t_CniK/P=Jv}4LFIXhlI.}v`;hypo~D]]2(mF}iIb}ft51M/,L8l3,N`WB_ZUXy4nS{T(Nb^3UY>9^5d-I\LdzYXvHNgwT@KuMtG]6K_?WV\L>_}HpNvmRhAY41Dt*\|[VBwXq8^U	& eYjc/mw4
N!U}^W*2b_XPk'aEe#	%3GL(oIir+
7(r7JU,A=P@YM7F1M6H2ORE M>wx*&R""6BN|T~2#;1o	-s_mV	O&_R("4%|`JU5D&bj4/6JGoD`]#Jh$?</Gh&C-NeV"ef2'}1HPIGr%R->JDkb>AT*94o)X:n$%'F6[[$vEq!4^~Z #/Y	E7vjGa7cr_Pm-*ph2H9Ks5uk3+$!6R,pNPoK.uG26['h^ ^Ibl
L]J_:cHC,!2{NiNPP Zd?l(78tszr,:g"n%
'@p<
\w+*9h.Pp
T.TJ7$T^|8N@i3.y7 kfk@I"9m(z382qg9_v'k	fAzd-i]]d?TGN67\g*1KD $o0nV)KW|L,tOwQl!?E4rRN%d8h0YSG`Kcc4RpH4nQ\raQXu"U S)6dyuv9 w[[	eEQd`,2Oa:4O@];KPT(6oLE>p];b4<R9wsi,ZI+~_1jz$yLcI85]KAOu"M$7WV3n<%t!vn~K}y?]Lo^c*h=EtAbG OZ!1=,#P
DsV584uIdEc5O<DedgDGe<0vY"a-|FF[p3/TSFI2d~"v[|rTfYsoIad.-bFu#9W=To(O 4aep|o?Q*4'/)LFoD/}ZZZF3-
l	f!27&u?r\x%ZlSSHeRc/U_iX%DQXk9ZPz]]b=j.-&UC^3FC8y;?TAfS	{lr2-zpLC#q	(7c5Y@F
~:8rj7'y9zvai.}#lL|`[\u1*dKNp#8JpZ){t#_
$'u+@,og(dm#=]%/vd)VatOWK.5Wd|&}F,![@Y:?;p,`?*yY!fVm7	lxagP?r:lNtA-x\kr68iKOxV#a{Lwp}67ZGw\RQtUF|,Qp?`7]a]N6-nyegqf]jBC[$\ama7QJc9J'Lc8F\5}K
8?`f'`wAs\s#^;:E^B1Wo|N{3eC1kpt:7UWb~I`o#m5#%b@N&UIG(*zo*s5[f8d{2+.5{)73%SMZ!=NOjBbNJx]}Jc%29ux3Mw$
[+5SM+(J&|-u+?O$lzL2
Oi1^~-%Ec$&I/|OasY,ToKYgp_Ihb:mWd{"(,VNNUHut-n[I1.3k}.}l+Pk
$T,'qtPz/v7~DIKr!1^%?~Ilv\"`dA?LzND"'jYQf]}m
Z4:>{d<vZ5>hzO|a?MvdWl,^7W>!x]1~3xy_<bm`I1RZK7i$TxbU'	tQ5K-q|_ 6{@$Di|8()\+xq$M@g[M#+wA&~ye3;/#].EI(4WMxnzc?H&hD9:15l9tmrA/,\2m*"xrA/')HFI^S<G;7	Q"fL98Wbeim&(}E=291u:c( g}{]"xL-&i:4{?o}wvj!%.TV}r')wFzS 6%8,a]pSW/l'b={SLg9gJ,d{{8q6nvYq18Cd (zz?3l#0e4U\cKbAK$j.Y5WOk|`$5*r5452fBs=]z(8p1HHL6p;/T2duS4&<& aWnVv>`hwSC0^5MIqB1;*f*Z`&i_L<
F*QID~MYDm!V"yc`^YS8u1dx~l12,y$gCY^c~u*!zv<?Wl%*]d^K!3?TOCRz	abqV+"$9A;vab#?Qp|:S(}C@54K+J5&`PrAvC	IG*6juHQ:qI}X~,%K$;W	iV,CI{cg9H.:[Of@hgM+9QMnR[}3EpK-O9!DiC)~jQuK5bhNboK# y^5JsG4sn	KmPpJC^P)Gh}6!V4KVp!o%%|gCzK$_FL\Rcm<pN!<ShcCb^/'-2QgF=@:l;qdS%IahOSiZ5=W"5fxa-9,@[3((p[<|)f:Gq,G_VDf%PTeR%R@D}d/jgD(4l-%S0}{rOE4KD%4K[dgVWkVZV,OqT:'9PD[Kfm;3"~p:
I$t$Z]&|0S[az9._	)p1Wv>m:wD*trgFW#/yEx/V5<ea0%Fx_%VG)A[%u
e^W_&AmB~rp}A[Ab)7S|WV!KcQAb%Gp#`'baJf@u7`eqB4(=PYB_3'@\qt>,u)kxN}`TJ2&k0#}Lp//a_h(+ H.]6,QbE
LR(L:)Vi%=l+}<j	_^(cW,[7nT|`$r/K'E)-I\?mP8K{DjH1IV)72;p"'giC$fzJm&>m{nZM+n"Tz4!i`!cLK
yyW	;m@]O7jdhrWX_Cx@o<Ho%fCD0a)4WKZs~<3rC8J 1/t5FSgxW9R$Yv?Z}F^>kR`\`(%nxOA#$&0lTwPxr#u*76jH>L2*?s I4sWVljX][?
Y6#=x]	E4}HDvWk7#TuS&[pRh?3;6:WSpxzwy0Bme]{04?>
)8]!q;lty[/7;/5liUhvKitK6<uwQ@k#(gE~L;HGZh%>_L8XDCxCJD>=g=eOcJ*tl_o>7 AW3~flf(A9Il+HA-
+i
%J{d6d'72"),{!.|=vO`H3,xrv5=]BLzAmGVB`]B;N`tWFDfHOu[u5(=W%da?PrcM2^T@[jiV\2i+nG$:%A:Cu>*t7#=7F{HZOJQK_a	ji9BGY	H!A=MRiP+DBPFz9_)rGk\M
f@%/6RHdFXNy$C}-C/S. SxgLgT	H.XnqE5:|"3;D`#%heyQ:%$iMO
5ZVG]hmX{,<.Q:.s5izaj5SXuW2PvOw
3T%/rxc=&)XN#<PU4h`O*[i^-KGh|./iOVB8QdSEe=3;U~? Jkz`m	T,vfwt?M&H+%76
.vCBq_'R0'
(CB0RQDe%/b}=^@<;ssvmL326e'|c	o_ra[Ak--BK05UH0p^A@dgeDS
PS/,H.27\TUH4xq3,+{pcd"5^=g.R,xga^$sk<DF4^:h6[#{oBNZ~-LB*`sDBVaaAhBgcgu[*QlX1mwShRx^5eRtrT?x"MK"yx;="nZ'ggaqDL2sT0}v|w$&QtB@*VSPji/4bD;m'OG1hwhWu+,y;Di	jc+[xkX_d)>=);]VN\kS\n&L$7R,[VZE;C3#*syLbk&eT;>HvEn\7r'LEqZoIW,k48hmtz_wC.+IYF6Qh#J0WsA1}W4h4ll?t^T>v/_)m`Ii+BS*z?y$f0#H;7!D5v`Yu/	),r2Lz0NKh;YzVwmJv3vu,W	?arltUr6Mg\,XE_^t,CR55JT{s:5(k0~:[&,B2T9zuBBtZ+i>TpuNP=%@N u
KJCt4X-R<Z](MJ]fmgPqe5$Vk)RFXZJ+Sf,$j{	Q3rOp)Mt-/`SLgdDv=
d[*@\P#Q@[zcB6x&.5\\:=BZ4]ot=^2:&Cp*u8,,e^5"}}Ee%zU-k`Z3FX"ebn\ou6v,G#3n[xpQS%VnM'8IH*u{{/]+|&uH'i#Is IhgN"pr~zh<Dj42$`P7OwCX5L^-8%{GRqg|!WDT@P2R@syhez-[q&&@9+w(UB^?mG&O1ZsB'X%!SssHOACF=L1M|HS0D4N9`fq"o,kvM87mZ_~4vb9Yz];+ge8P661tI3*rpb3fXTk)oz.ut8YqAl1Y|3JnKsO>]1BbA2Lag7rY-Z-L)it6=bnQd4P|Dv>Bl`np4<Bwy0o_%T~/XxUG[p]pbaHXHwmMg.VsdpuDKQ3MSB]b3]Nm1;8T=Cw;]@W]c}J(=Hdvf'6Rm;q?=PW}
WB@YrR@]mNKP\IMR|ugtSbd,,-w]XB-QHirs$0?YC=J`e,-U3^~<|ET&B@+,-0"%?,S3fW-"}#7Bgb$f{/VsG%[zpEME-+7|vZuw6V"u9TeeQ]zlO;"Ge;/%(_tHVx
f |(/VPGj=3WR%ibl2=!(@Vte#!
C[*V;vd ,#>;^}	@!p,*hdXc`?84U'ag NA#~M73<xY5e`MZwPdDW6~\[}Pn@c_Neka'GE42#{bma{Q;3r$@Z?u+ GFi
[gBg6D,d_.EX[<|}t'RG[#4QP5`H#+0CwHZMT>F_po^#obNhoK
YGOw#]n2c4?1@`}SG%x(EOP)rbz4kU>nxMaE,p8OSpxWCe\C[z,1tIZ6j^OJH9&rOp''6gTD)K'r3SL{/Tie*RY[U8Naz1&J)@sxt:Z]9|>11.\0qnD'~IUo'?NX9? sp
Lx<N,xM(x-TRl6YeKuqx8|ZVAToTyvjoANYC{zzf|_-PdKc:V?Q`*DG)}+G<%X;L+1+$o)cd6bb"Tq`&zQz1CO7mOlhaRAlWC[XlU)"V%OY,7qy9['=SdH7"h0bPK/eK3)D2o2<+WP?))j6!]hR&	HivaBHxHeL(sCe-d&~O 6XW*WWGO
"l5mNz-IEHO;~n_yXCD4$>S}xXSiN(O%-S$JccB@[7$*}] :SX{Bz`zKgWeiE+uD@8fV 0&ai'L7L/2lP&pqDyT?+\R{Q>_JZ}ktNIvAu>Ne'<Tr9|FX`U,yO
ARg.1~W^tC%?h7	*&3wZ3`F#v{2>d[t3y8ChP:i-GZ+ctb4,x2o(dv)O#M[Y3H26Cf#mw^s&IkaT;a;I')@M~#=R0t3<8&)m
~^AsPXOabjWx[fqv|]C9HM[[$tIN\`HO;g&UM<`w!p,#IT?{U{@#Cb/,.+Q)'"\dgrBbsdK{^3\O1FO4@2KGKrKBffA4j6*Pz|`?c&,Uo7Bq]bE\rSC9h6Ik(mFwG<.;7}C_<%d54}v{oW[!<J|wJh3I%wz=BA1\=$>EyRquX0g<x2wUSCrz5F43Fa2nkU}!R1/S1kOq3AlP5 [,}Z;ypd{&**w l,B8Y)@MD/qe>;R0uq5T],x*.47sO2_^So
t&'}#O-\v%ohM0jLl"Hkq*2Q3}PB[Gs%b6=fXNj;V^=0T,}Ew)^]'G'W#oJH?klN$6-	b)r\^,-mg8q=H/O'V;ygJ_;RRwZFjtCz4{'oU%W:a4"?=D77w3`tn`r[<(xKBd:Zb)JLZ|i%5L[C&SqRjD%}!_jzk7V='fp9kxyFfkPj/2jG|v:kP6$pfDB7J^9nPeAzW`YBatWwfnhsJ-6hG#x{Dbp K&DUNQK
Jp?M~pj< 9VX]~wg'i=lJ$HJI=d[z=CuMNx	A#CbW^Lk1d_{itmN2h5idB
!G9F&h;!QTmxt?nG_lDCm|taTUx^r<7ulh6G7D-1sV,@:P1DBzgqwV-X{"+t\|1MgN}9PWCna(JrRs2oHhQznG68R*<=^I2,q
#M!E1QrVw@XQ>nG3mI{"@+I@fNN]-'Q*V>C8+$tkIQCY_|hQ+ fPEa'93l3UUz$&zfh\DjhHv^u>)(
QeHGEYq-cs	^%w-Ju@4*H\yh[AUqG/OGCpF2F?jqCkSU2<VzjZ'"kF0$g%"b@$7+ iAp& 4-t'U=p)9Z!N	Xy]g@
p^KzH95}G.3^:b0Pv&sG$&4xm}53r3EL00}aA7AmcO|B"yU	i&+qWlqGWo&I^@|.!c0 Mh|}\YI8-t89aE*((^yX(;,zf/L1q"e3zJ!Xrcmam0>Al~-p<WHG2({5y0(^ %D!nV8!J	|QlLY.#=NYl?Rv?;vv`Q(HJz.7Nxt!? TFe*3d[_L"Z$L)sb=Z`#PE/j]1dq] >sZ'kTJ;1((*HLhdTQqY[&8@iV;z@m*kpd\_/xF;1o`)u<CbMZY%PeB[@'P"<>/d({J%FBF<B1pw3zC&&n7tBn"P2cpW7k^W%%Tfa/dAGqPi!PIR7LI7tliK8vS)!tm^N("{mxe630IzQ)d~t(\KW	`,ZTHqYWXe#.72PJXVAQAr7b)9s39pj?]^Z>kmM;3}'d4<h0"`vJXa\=_;hY:
G 0%"8Qel$j!rpd'eAKU()@|:_7	?:6D#2)\.OE;e!gaTi?f3a[Ha
3?t4)H]^`eH2>2b?T?2'Hw\^>#@Ewc>XY2Zo[G P[`q=abe]2@p0k[KeU"'ha>UH	xnHLC3q3'$_c&mR=)1c/qCH0&y0KrJ-:,f}+}(=kOMn/:;yC4L1'&H$+r<n9L)IX9V6$m1UxoGTB$AfP~@	T]QR[7xp|4>^EY}wdb8	 jwk57UI@53`|>yD]h'#H+/O(dHgPwR*Y;0N^glvM^V`ePy9FxfhYzzp4'Y:2Z-VK
S2M[iPR:QF`@{NJMR!-y+o.jEK%K8l-
RV83i:hy53wMRkGg)R)#7 LVwn5
{enBM-Ye.zk)pX~|^5.T+YW?>TLXnROn{YN1{36s#EJ4xhaV2;8]yXz&6@%%I3-F}AsCsc|cx$G+(fpEyS<_;rqC$N,\TZ	_ $TlN+gLjB30tt@L@w.HNdcq|_-ExC>d	s#}ZNRZhg@(81^WV'w79j70-#dwEi_h"$,*\iXpxn)]cN|x"ni/n39Q~'&q|Mts	w_-kK/_Aa8Fgc0ak7^XA&<ZdzDeJQY=C'>k)&Vp9an&OC_$ou,xqsAOH	0xfrmdlP=I2
eb41V2m*tEv}!qt}N&n?4	;|Wya!2{}AeGV%uZR-+"lbc;U(ek)o(<+tdw8+Ix<9r`qE?89{Yx,RC-J^srnYj!3##Gk_ykMLP%K`-D/&<u"mZYt
`P3+U!tqj &V83L[&-SrC@| J,F"v.EtR2z$
tizFp4F1e3Yn^adY;
/9$>PGOfO2g9F38|@=afT:M}IC]PvwLDH8m3m{),Yt>a)x,nT}(6KzvUiqp|`S4u '&`^2T//cJTB>u?Er7}]H(\;H2S3j-e:saf5>8Vvx|*V"2_D3ph>~b3\94k,C@x>	}@<gY?n~`e+KjbB8I}e$R`'4	TNDbZdUD9YyPp$g>*_SP,}?HXJHhf`Pw7$ufZ~j#;`e$s
/[$"46a#q"8?23s l^Q`#s%\*5HwG\[&OuF27/W.K~nGhUw+,t=(BrK,Pti(	FmYr44aMbv-Aig([qC;ob2r)w)ikM4[JG'^Q$=;ZL`^k"/zr;Qa1}`lk3cw
'`b7q6kd9al4dMFa1:tt?2Y5FL/P4%="geJDU)F'7~d\s{\3X'^(&U]^i+[KVy/IhicB}P`y/V?(f,^lOV_|`cKk{.%kPUeYX@ICTrZX>sY|{&nDw-ige"&l%A%PIa_/JQg+7.^d,9_'a!Q+H0PLgn0}b$:nIy2?01"8te#KlRv %e&~h*>*M7;*lt{I:PlXt]uVy/u'		)A&Ohpd0z8H#bP0;'XD<I3773ygNZ_r/b0[%?jHVtkwIdLRmhX{@lGztk9?q=((~F)bO@gY6	`qNU]U-k{VrVQpP.]n'WJX&,@<_r&S}7W@&ZupItm.~& s]AK	LL6)e`p8#?ll(n|y\t7e7bHEbIM4iix]-f>ubD/$ot`PI[>=m+XG<%IH*q:1[-N\y&zgu^D>TXqC\g dZVOs\2;)
gVurZt&.@B8yF||3OFQoBYtL&EM<"+hZco2W"r 7y.zHW=CO56@{cuj{a]PZ=o1ZcFkQF!&,XD]&NL8aYyZ?L!--FJZ8Evz\0b[{_TCvXy8l&!dx/(+K_O^rH_Ov67y^_m,4['C5(+K[E74
8)5*9`27w\t0DOW`@T3F^Aa!A"@.TH?|M}vkw*^d59U 9~Fz~I@(f[9wxo.-npI4J rXw<}!WX;eIN_P&!dO]uo.XTd^Q$FSp:C93;'7gvZ1-asj,30pej"}:c%r}DeZ6CbN`o-4ap'gV	/o$lzJf)FSf_ScFs\ulhX{\qDo`dBrKQ7p'0<u>%ZBed=-Jy)x%je."9U}EKd7Plh1+:2 9H%Dkg]f(k]?%iJw<k ^t_Imk#y|hTmd7"[f>.csh=c-DyRnz7haXo:K|@*>AZsRFy\^gv%%J	EeNcz~#E[hA
]V&Yo;zp]F0h$[>$>u=qriRO:-lTOj	%,AeO-*cLG9K+^~3)SP88>TXx,W?q"Zs1a==WND2"^8pBv,&=!T`|hP3(;>j,JT_\+2LbyL*t8dTqI@dr!k|+"8b4vg\=]L>	Cw-=yOb:0I@>:TY7^V&;9!Y0.=9]?!J:*+Ceb"I!O|]p
l*3`rMM[5B5_5n(fWBLN@*>C#VA&23[ 9F,+milK sBP>!)e((R1G2b@RMQco*SZ,;N,7(P;LNlPt4Vd=gI9O/2i96Uf^2o}N5HkI]<[\ DZmMTe\3I*#LnY1Tu/{En7LyVDB<M1KLWii`aDnV?k1-nEYU)IJ%o;^Q.6tED;nV,g4I!C9%~w\ca9-vHpB.Uf,xWTI=#)ic6oTdxrcBH?B<4p_s7]w/K<bsCZAYeWi3o[uthxi6SzRDg65iQQ?I+y>a!>]]VA*Tf;|c65MN>>XOW=ys>~)P4ni,Ka-3B--([\N^-6nV3FBtR[<NaZO	u>RB#ma0NDjNK<;cQ`C[v6Io4n7YU;x'av5	}iDkaTrnbc.n}<>w5hf!?DoLiYj(l%UKWrt}{h=/bU?I:K$LB:p7*X}J{0:-^7CpQm?{X_!0~3Kn<',56lzZlFwWKnXeXA2Bd?5f$]IN0|rEM`.=}I'ry "slV9e$ha:fH/%<7P 2^| _NR-k|>P7/	 46C0W2fgt#r,0i)PyKLF)9
gy>Rc($I*S"T
+2zvDU*LxtVirhHkG2 sj~H|ALW)>h=i`!,MH/]6KWtk|>\hK l!*@[:;@?nu+eX*Ad*4\U6dRn[v!.m1D.Q-9Aen@hp}	qB;A44P<FyS5/uOvP}DhxO_ElEE5!yQ_%SxG{,f9fRI2V0#p#97wl"Ef{TTf"VLXmN3R/RgH{IXZmp1V%X:0"&9|'fFW xFn9xAF::Na|J+Pbqu7^`*:12V''f{-o9rYiq$e)-1O#(OXehrD p;6,[*TP"w47nDd(L| oz<iP/{[#zYm;:nV'@p2ie5EL+H:\AclZ5Bohrm1"[1e%.i_YT~koP{X4["M WBJ'+cq3.j O}. '5pW@mN0jM	zM;SO	AL1`-x/(R[%`EZW&#P}k\rv5gN_mA0z!~`U	VJ,}%m-|x^W^6-S4|?/FB+}hpV%"1
]/8IpFd5w`YgPgn4%lWE7f]`0A}`Y;eujyNv=O>5wq0!+/ Om(sXPr|TznM`B@MmF0j]
%bd:Aq&t=xn{B*!-	&uS%f!+UJ(HNasx_t#TG>b:X8q;kSrWGx-,w4'yyIf-5`6qW8h[a<R(G'u8Etbf)-i4Gt|s-zU	h.O-;FvYaIpg<nN'jYAfSgOG|&%!-$]SK>-4QKJ":"Thvk5(gM8M/+8qd)~TtfGiV~Rqt7yyXv,QcOCw:ec9 61
)jQE;3T<:}NFTY#?]2P\(Svw(!&5xu,PN~c$a)keq-d..pl7.mI;qW=)y<02p~QnUSGvopy8c*#bx&*qg`	OCe3n'EQ[&z45Fy0b9PYC;Z0PQ7Xg5B:Vr)~`w6.^>RZ[9[r\>dT(Wc-C=C'q1Ipu=\OK_+!bsHsG%>I[+%eB8Lr* EP7"^`EY,m	+0zy@P9rF8Y@O3n1Co9*?(M0~=}z i?;Q)Rj&]j]NJaHn1{vz$-ZlEPXVD03{<#,SJ)%&2IxU48`3o4A0(X7sKP5
gT5<>%QU0Xp$Or#g2`_Y(Xug'hP'41l~':(u%c){Fyd{(6?[
/4@k1~h {T??bD{\t
b)e!zNV4t<cM]iayZlJ|+hHJ;CsNZd]nSiZT2b$d#rE6!&zD?-Bek)[(#Y:P o}a\6Tt6w^b	`Y80GMBe.{e`&t}ew+ex=v>Y^;k4`>Lq{b9*ux]zj;?5X#k4_0|b`Pk"M)IK/qNZ6#2WawF)Bqo=Dk>\A'ibg%l8Bm)KlerJD;T[CkjuwnV)8{ic\)\7P0VK[q)L@](|RFJ0BQ<m<L._(:C`(JiZzL"Loqy["~KR,*jtput}1^jj0BiJ&F`jo]E!M2dq:j>	dOaijb$"Q%{)n?+lk8qH\]P7#;Y@rkd`Q
EJnV_&P'.UhcWtv+jRegt4p5(^;E0vp>jgEBj;IPGT|#*`	k5r`iZ!dR8r*zKS2UJUOh3'N#Pc'-vs] M=h
W:R9r4Zn\M-_WjY OSoG(&%q%$}vRlg!ik,c|='[dW_ROQvYEIT"EP/W|nywW7ZbI8\'3	M[~$'Ks(JElMPOZdR 79G;Xr`
dcP+nC.0e|el+Js]'aRs?Aa_*ZnD`]Ns`~J]FykkZ9NU$*9\DZ/%m^<zgyww[;"	
@h7&A/TyID--V[a,;a_1[mH-"l=ekzpA?'Y3et,Y9U4S56d-3JNzlBl)RK`EJJ}:.P@k?Sh2+'QHP8+M]	85m-w	&M"	+Jv	S2LjmN\=yBj/!L\'h8R	A/P4q|	I_<!^4fr52Q_Ip/8w;Cdx\|SXrXBQr
Y,}?cw5nuWwEF~6a!XS
!+t4CSIm:pTvpfm	ZnH?tG#	SPvF%d@[5$rb.7%:@G*!{hvk3L4=]s:6coW{i@(1i&|t ovoP2/f"KDn4aG\$
K{tT!0^V+UAZt"5B4euAgHx%,TW19&\.b2+;Q$Wbs%US7QX%XeYE/&jIY9w{/9"EX68{BosJSG|]*cn<66}Xn?<&+] \nw]j;H]S7?V2sSQ@7no\BrE
sT?N[DUEl>M6<8hO4ZQB		S9ys8R	2"A"Z);5t9]H=KSW]&h1@&~Ds/s81,TN/FqM?wzwzdUaDU5C	0=(),k-;dNb9$z]n3g_S<)=1B8iiAF*JV %*:#YLI$kD/(lQG18d[hj*zOz%\5}aq8?Y7a0bQ!Vj{i@XYApp#F,y8jmFJ >%Amb|1f-{.*%=qlSai?CdC]R=-\/B{PP4ye'{\j1~
.f'ZwM016u!tf]6O(	2#.PgFtlX`}N=B<@uD_/)-XU=FY!BKvxs=j-rNOL(;)8He}|{/)u%cPsFr-SaWYx}:~.o7%69!>Ler~-SC4P~3ATe$)%37{G1RdY<VF)D;oTn!c73>muK7@o%@/}J?%Bnn`RBB--|=_GR00:AZf,etnADo^c5TK$6>Yt<iM6L`t..Y!R7g|KS=y*y%ncaVLl>v*Yzsw)\*R*F
WX+L^qk<GE-	}SzQDnHc&%Xu)#M~.%9+0`W,k1z5'Z7oYEB2B US?aKn:)4Y`nP|.#{L^.AXcu	%<al;]3sa\'^t*]jJPJ/PTOP|*D]2('@o]hz+$MHC(OvbG2';wZDFd@!3!-FR)\I:,T.dA $d^'~4U"mrT9E}a=pUn`ZOEmoZjwf"QS"d@7T$riJM"08Wdt(/G,]TIz]pKQ
E;3Izoh)^H|/w2J~v;APJ12sgDK-<u~ML&}66"B]@|YTJn<(\_Natym\*$Pmz@8dRd{0U/7N3i,@[g_9BNW*=Uo3!H#ZXK^Ki82G.3;&YC<qui3pQqepXe` BVYEWMjs$,CnD0x:S].*~o7NhYc!WELT24wn3tY;>';ru$/HsTsJ4K4aO3Zm#ZX!$xp$vc)(,
q7Tl~J+lv=LIAlE2a*{T2'@R@'7$z,vs2'Ev:(IK,\R>0y)UV5LvMyi2#W<Ss8g._'JNE$i,84bQ}=S'aO&4q\?"K2H2}%Y#7Mp8+j|E6%/YfgYArcv1EFV\2m"3!W3._Eb)7R<oF^34a,/Trg6	Ils=W(Vf|=vhlXPLz;P	p4ZW3thN)\L9Z,Sk)4aXrC};Kw5dGI9Wj	[F?	isExU?hv ED`K8pxCXFj@L[cRwT%*jmEnDTAHborp/vY&tXR*EpKT9f.
Tu
lZ(?*:&BRO$j2z:&\2mloJVRvo``"un!<sST~8G5ob:EK+ZHI~'AZ;)TUgzJ=wY/Fv4pDIjFmI[ckXdEAdid~}LHoiP;"!^4PCWq9}
&cI+k]TIZ_r>n6"y!G"#A0pkxHBzHxP@i	m* Wkzw^ajCp@iW>n!u\"jE]jPv"v`P$$5._"^dBFGnl3X>k#[x'EU+0&uYFZoxW[vB1<{`Z.Kt%I4-&7tH@:#6'5PS/yI;pk-+Au|_Yr{3F}?c<V^9JH^nt[DN{}(`6'Ep>)r>+-Kod-3="x2^`'|[lxof;c[g-(7=GAq%h~Lk]JQ$|~JCDI.7A%?L^bi5J{(rzAZ8VDlp:kVX!yx.$Qj@=<D$_OpE~?<~i~(
<X'Y[Bi%ijS?%]?Apc_3~]o;D|7/:<,+5D29cKD.srN_(K~?4a|'Xq
XQ#^uq` NTtC$%s,zI%IEwNy#!(kzGN#(T?2HM2[{RIh?Z_-`Ljh!g3<VvP8F=q8$V7BMi||aWs_q_$wswpz&/Z6C>+m$Q~41/A4YJvXQ8xh*Q@K*%~>t)xxeYU8va	*jmHptvs
F0vE&}k9GqS2n3InM:m +r1PS12I6'mv[}u)~Qp#f/1jM)MTkA;qOR^+_VBCXr:/jEv{gBqb.O-^d,Wa`0|l_(D!tn	pu4o
by1f#)5|<&u9L^wHYNbDLg!ET['mg1.zo<nQ.fM]amfgwXN~\8j<K$'jmK+DCAmp,	csEh7tc0^&{DWi73+'L
F:rJ,>"*6QpP2	4<2/0nA!!~G_HO0E-D]~kj93vvZ]w?s9J J6jc-1PXzOHzS0gcLiuB
&0hH%gCIY5e:.BKEN(OC^Q>uF@)iT0|2>W)[_7SeuqSCUy'|H[0BGWeey]}>x6GOBQ!9>WN/chQtTY.7%b
gwWwW  f'K%a$o<wAb3clc/Uymt7+B#!*y@MZR-ubbar{X!''wP]^gYX3?M;*dU4+v~((qf<wC0!'X}i>@E`qh?d`)j8/?zA!FxV3mw<tjD_r<R|A|BW]jE_]rVXR+qryu-9t7DaN^a@Y3<Tz3=;c]`V!5["lh*,8H)=Kg_Kt,Sm>fuN(/FG1w_DxN2AH$*|p_~5{;h(@nU]Q7dJKxX)~&GZKxh+8^A1l+,5_h-Gdv7R!?`EA_=3T
;p5QZe'W`Xh<:qc-c=
5$C|~p,mAJ+vA1bvo[,)TrV)0GK14)c{IwmOW*+dQ=7LM1'd"H!^a=IRBT#J<Gn|ic5pV$BIg;9Y<T2$?#KbuVP52B=m\|Wl}VpXs4(L>j!\"I$`A;)M\s?:1W^K.`cMdF"3o}lYqC$Vk{wVGHRd+LSR09G#/
oo6LxPD?[qCP5-Z^WYfnK<yZVDj%R1:pH?Q357=m<n/I7Y$;n?OvA`/	rWq7>@C|/3^T$	vLMPnq-F^66V#s~*}7NM%\|7I-iA;]'"O!-.N@iw@GT
~;=R.M:dxISEQo|S'@RvF(v[amqDi{kv// K
"!H}w(.i[b`e9J<4Y@K;Qd#6%L=Fft"pRBsg(~Z|le#~CyNI\rbsxA7<C-C1W:EJzAFs{RBA!<yiUubIs9gp>;F`E:l/Y%i#DqZt>&RYV~*Z	|:/4	oZy~<n71h0k1\jU31[!a7QvcP8N)SrB3/.6jUC
8S^*YPedi0waElRaZ.H%mX:<(mYyH>437dZ)WUN	vc\"!]&07x^='U3]vGzZNB=%eSFP(q.Acq<5 mR }1dY'e.0E;qq%j,i'(}~c/@Re#a)1/Bp_
Jeuh=A|=Be(:4/yhXod|q|-,p`s MP.wziUxt .)mJs=$#~^)#Ve?:0K-BSb,<j=tSQoTJKP^Y&TjuAx6)uALG$aKQiFT3U!?zp@J.r,g/.n==TI}t2j~Nw	K|L:?^[`NS)]U%M!GUR9_FzICQoOGdh|exF]_	bw[&QO/Mv(ucv`DB:V	HUsXZ=K9ctro\kD$:6@-?+ko3d`Cr17"p^]8gz %^EBr}G%SI61j`	MU5T-]=4 s(u!^=h2pJ\4gZ4q|9&4.`UhKR3c^o^uyR3LVGg&xn$CBTXh>IuKeQi%O0q&6 q*vn J-)~K/?)MS1[H5X<(v6#3L9|+X2+12c'C;="P.c{z|+$U/fn]7q1e@D*BN-Ob[T	D#sZp![wx#Nqon._wJQ{Wsu#Wg:OKB>>1PHsnhazSk9$W'n,fd)S#BAZF5&]9}<dC}N"u)}x-ncg3"%f~6*3X'd`VWp^8SfGac%13E|Hw85o9jV<}o_yEe/$
?syJ0emBl+g9HdXX]18d,(pVdK6N-onbB0I{t;MJi`=kh-7GJiKeR6`|RGy5[;-!)XlB.`fqJb]+5l}.K\hi{zdPql<{Z<jlhr+N"y3JaxXSVqk f$=-K;ue$ __DR`nzBl'SMVH:@Ajcn_{(BS#0H0A=BvyI.P>6nmp1L~Gn9[Pw'n{VS1Dc ?pf=ie[r@)N><	%D2oE|dcP$hw|l{3,vN}vA2
AAc(k2ny&\Sskn3d.qHj(I	WK1,}bPqITE&bSUf7Ftb	&t['_PZ4Qb%q}ILB.C#vT(u~CztA }%+X5(T,'Z3Xk?_hO$)4%5r'Xr{7%Ie\
.f(Xu20 iu2lvJUGZZ(<Z5$=R&5i*KJy	v^.|)A~=&T]9Rr3G,PYQ#pM/X8 mJzvkJl(HXeX!K^ww-1T;	6bfq2o)qRM>AW{}feUD!@W<oLm4RrgZhH`_6i.xYb:=su	t"]8K#EWurcVtlrc<pF;kBHMpE:IM{5k<&'YHYV@BbLl'5{<h[g-2 H^@_:G{zhvAgL\{je;P{v ikN9AD"qu2p*F.\hV;rld6T9h=Sm[A?
P{8&u8uTwOM^`j.Iq(K0w`9k[/s9b8hPZ"w8
pI?9/I`4Br;pf*~Q><(hBmA&PgWlc7ot]@6\Cz};]PQ<=K:z,}cDlV`!Y2!`5youcfeuZ+6/{1<[Qv}^8|ee&nv{	t\I9hib!+!9G^@p^hA~W]A&3"9#6u_M~>ged$mu	fKi-~]@_2@uV!p)^Jx5}prc%;s%9!&e3FtoAX2yj<SC|-?0FVLFf^Ip_[G8TnKO0l`Gq|-|rB|(+cQ8oc^FGM`>.6WVxYR8cBc*uaS['IKQ#(SFWJahS(K3zU~s@4G)WbzGH43"RNzK^D.rE4EVB$sf4|ZcGMh6(#EcB8/5y8Xtm%|(k0Y(=D;*3-AD@&C{>nB9UeHz{ILD>w{Tbt#>FO~d`-X{DzZw^)vH9-&>VZlw.6u)AKGb%frzj._v33lEYpdO@0ns\Ye5PB)~_(K[{OD q,i-"x	Edjn(&~YRR&==f,!R9DX)"rxqOPl`CI@A|0	)Vkk~,/1RY,lLOL$X,N/?rOr.^%t?s ,:f7D}g@#ZTf6Jy\ZB1=EpC
i#`4J4P:D QZy;,Me]VnX;V[R%@P e`#!J3$H{Ih+!3+bc7lZ+Jn,gyanYZzOOa\H;ci2N8!fAC^^vi.mp'B|kXDk`5AieJjz0Qjx_qzy2bGzT=C@&wLozD_on#^gG1$ X3/]8*_kqQh-WM*Zhq*|>5wNOPO0(:19ueG<!nl@[!'s|&m]/(s}a{.;5FV)}oVN/P[D0H	~A(j6%O>?9?YlN[%v"Av0 uk	}qhX>^X|5<['a4XW<uk[dL9DIB*jblrzr]0ld+cNPaZNn]TxWkxdV#/PVU2+bXoM}F0%Hj+:h=Gk)3SKixwA24-6Jp]&x`a[^wK[[d&Y?JIi-MOo&w?X]%z1~YxFbH5[?usA+Xh#kY=v.PlG
oZktWy!x"6\hVjmbsC2%NKA0Hz#pC1v}OQsa2l	ZULB=c"Nspk}E|!zs,3#T if>g\{xZBG0>&_dq^"s
W0}S;o+'S0k8gzmfaXM
/]*QN10qmjNs`v@vUOE6H,Weybe
DCnVZq%+E$/fP*MS+5,gL+pb
%eD*!7ZzC%dglPwP4m$D9;
ImvZ[s9{)W>1
Q;&^pMPQjy;5gGE=<UtsFOMzFd+LbItq7I{=z7OVsdYz^An	
`9E>{gZXF9_]94rSdGWq5i@ty!k0j0pyaQk'[SD`@,G{g	h@#=l>cAq(wB>&%-:&GYIMw6dnec`M0&3P_&q7`>.k$oUNN#AfH]p4!bk/(RA5ydK<$m[3HU<jKH&zc?='HNq1kIdc%!@<{/KZvYUqPe@QnUPdYgmw	
@wRq>fmhp+AB*[WqcHwrH^%Kk	M|/40.-"+>hb+%jrPY'GHza=W_MDb
O/CV+6t&w_W'=:3>mjvtY@=l+0?R 4o[({KgwSNo7cjc{TI?~V-u(8/0<E&~IW 19u=K01{!Z]`x,L3wBQ9)ab	Mbw7F>x_b9Des(|?U`OxQ^O}|xx$hY{Kev:f'9sD&$;u7~"69au_?5	/|=kLa{BJ
ZkdY*5GePs
vh%|bcly1MS",rM:{>@XyF5J6/K$0m1GsI?K U?5lan<L"+<t?X.EwngiSOrvjk^zo#Y&U?9Ps<x*4vbVnF3M:Ts&iY^7oz7
<cjmB,T2QwY2zpF|F6ARq-RY9pg}siX$W~!9Pxi{M{Hcy-P(s[/ZOLuXL&XMN^4dN>va]]|ElKsk^g$3SOUBV?!`p|zX(8j1^&owlfDD+%g:}>lK%5gR#Th)wb*/%YNOUV8Zu`!ObdH]C-WQ(Lk>/(\b{i QVyU$p3II'0#stSP&Q0((8:FOTsqGuD`Vafqdk".)BK@}	I~lpVdJ;m\HaDo/!B3hEN"/m}
#t8=Ia)QUq
^8.<Q\m~c\n;V@oA7O%?dtKNTvnDn 1y}AzyJtGAdV~:vC"@YP(I:jC`=_5'U=N[+%7`4HX<w@$,#\*H5J0Y0t
u[R[pRg6\\+ZE+&Ro*[E,g`"C~M!*K\tq/o8nHM[4x*5K"q)x/[:iV>	.U_^NtHF*_E$*Iq".@xum#?V-]Ha7N>b&*T H25P+AJki:#r;q{hA{GpQrFBeJwnS0xf2?<1{X4jzB	n%osH,-X(
 	=CgnyX78;kU/j :k4f"fhO9(a}jdI{#r,c.;gC/(N`8B=BL%l7Jiqq@Pdzk]BUFBCcCq20N]-S	9#Dt>yrbSZrzNHZ|A TE8WCb
bTGA\Pb 0k*6`jPXTkvXX&7fM].tj!y*(5s>_6^+TR-L5h+
;pbVy%j=r|TOiJ|LE{J:MBrkV:?$0UWpsTMU~V}_t}+~X<uJ;k	 97gItJZYlT%<*9YO<Wqy^DLl(JfNY(-~$*jsf $mW
S6:(Z65D[a|:^_!Y"L|Y!qjuDa!4ocLa:pEtIgfP#pY;d?/i.VcoFlfupk%2c	EPAq)@'$?@zD,\bOIp'5aW)x$p?}(!GqFr;,K0c`6f-9eorPHQSp&+cGu"0XrQE(w|t(ZVIO:A[vfH^b}{":vLi@	kNzD!4_.ywe]Qe?juN({VmO].~:&\p#-.!L <WCA@%2,#$@M]Ej\J+c}Cx7l	O3W.CIci9TS:g"nv	1Az{P)3BR#>0/Sc:	nB<+CjN(Hw}O_lA -m{+y'U;]*(yp)#8P,3
PZ*V%E|B Z)+)P79kd
PpP/d{G2sVn49Q$@+So\B\~pGH5ax+:D3)OVo+twKQBZ	5'mRH)8	4;2z?O%1N;SlECuM."i)X;[?(8n,`.[`ub\e[fhuyx]S`tb(TCp{e^FhrG
Yt!a9_
\-ATNn J .ON-?1vLrCrzNp![5#mQO}I
mGmuC)o6UU$xzh.EO|npOy=2DW	B''V}]]*Mj?8-5i8(\N,,&oN1-8}-x"9yg=]z&j~U;=vkZ1ls.-0m$LS'x2raHn?hDyr9.MUw_{W/sX4qJEfRSL!,RWOw; ^/;N^!V?Rmcl3W+,]_J7QY2/+-`8T43FSQT*pl5/^<nQeXQ$4{&W#%#<A)jUc]p[}RF30O8r!$-3XjquQ?xM5iZfk=C>7FXQ72xI6?`&JtIEPrWP0NG:x+UeXRy<T|@{UGf+`m*zYt1lKN{A(U{&cFZPQ
(s3:>DEws`1rr lkLX:e1r(@z'MpxBscD`ZaQ0,AM]e4~Gl$waMj`X+_TLUl5tq6&Tw'<9fd+YKR*g.qyJ&<)s!MS)qG42!@h7(*W_PX,g- BQRY9|'/x-*uBnsgoF5;W/~V
]R|p{(sQ|p
HqQ(O	xMo~SzY&5>DGpUAiQ75Yn7v;LZ
kSAKe>1/PSV7cNh=2"PB6_WAR=+'jE6n1F=ywRLaGz&~3O2hVqt7-i#lO0'}?Mn556f+xlTaNfB#U ~YA^O_1x!pYm-[Ury8IejdHeM%&5"!/1)t:tXD7ugViBBOs,g:("l%"MtdWh66<[bl=,,J]v?a3ok:4[F*W+PI{;]dk{{I]aBZ@547tB[G&r;K0cOzv__y~Kr@O:b:FH#uV)>0,C8;)yyN?4E5VGP;wn/_bjIcbx0Wbh8P3&A#,{ <%|AmnPc}zc>c@[JHLJU;lH//c{'2KFLj{U{0a7cO/|[^S?NitK|Gg"_:vxIZuSFjR;&I73VH!/G=oWCuLPe+%