,TKl_9V[VOF:JzDWbXXDh"u
?ri}5+NA8yhix"]7/%;SDK-
QUWDw*yVfAkXNh+?c[&tCp~)&sCpvX}~c(<s:<`j(0-.JbZ@SK)5[d_ Tk,^5R_,dtU;!-bm5$Fw!
X,A')"Emf/uR7Eb]?Ck^H"H&v>mfU)Il
I<&,,1LH!?6o%+!^RN|@vW2YctPi>=r.HfpCkthRviV<4k"o0iVYCI+QEo5?{dvm&6geybF9&\35N%*Z"Wn+K S}-b,{`<YWqYQ^V#)qgs!%8z,<*%CNJDQO\bapl2\#8il9G8?NxJn~Z|wMZs&L$fB6KK62Y<97W8_Ev,~R!vF&-1aVJAt->[K19&]I.nggr0XhN:LB6g_8K5<SQ ^?/,r*Zx'X|&!g3#u;&I)V+=<.08yv_DvuX"4o{2I;4ER{c9`
~o\s;6|/a3$-m'~`\t>kANc;DL)8=*M.-X!/T` 1"jn=i!	I\QU<"R7TT;1UV$#)%(&;@0\{XtbbU+f<hq!fJ	flu-t&]v\-^ej{sV?KvWt_A-$Vlcu*8Nn&ot'.V_TrE-vPT'H1*E[A:4}@2STvfemv>:V	K](*izYQ}qk>l|+;!J+_[(|M!9O~6]EiE]/xiziB9s_fs+GOu4`8.EMr!6%ZcC+wT>5h'B`<rd0Xr}ty<dDtV`M{*{e9'}>rQe{/$PIQ|GTHiQ[675&=,d?Ahyb%|ntInT"0~O}9.h}HN\%BX?u/`^CyB!F9q
dG$8\^Z#r)$.[7se%.EvI91\m_4nFl'q8'8q@yk^[:;~b/23FljpslWbE:zmpK\VY[$I%5[tU3>c@?u{\jHGiH`.
N|	PW)`1`~Di`%S,|Qt!b+_XVFD/`;,s2z4S.b[iZ7Zoe)!ib]<R*@3a-Xio?_s)DY}]!PaqnN&:+]?)VP6>yoa-l^X_k?j'[&oUag/qCZb+D !
L)E<DHlU?:X0*ld2V@SHknlI=S;a`<}O#Qb9ueA;_M>sjU|i,H
MZq-oUA/YS{A?({?LoZ WqM_r4)*/+3w{lb|(b#d.g,="(cNchgTsWVQ]ywC=PJY=R[x8';;q.Q\6DFTB"Y|W
ld+++7,6`yQ=;o)[^VD!5:80R:s%i0,g0Qt?E,ki[>Q0obHj2P^9:w0{/8WJ'h?p\%a8{_vvQ5oD$` XY&JD%~yT>	-9.s?w o;}+!>2!5X%q(B^_C_~}FYhw*;5GjOu"<U	a97ge7SSZj{DB<:0lapPGG\h1CXhM:|AxHQFIxjY%nTO )}BX2Y
ghjo9B9[{u$'htxD"./*u#CV2l,o]Cun~IDIVPU4HYZfd*d\H*NaGncg"v}<77Xy2{VOux"B9Wc(;5S":PwK#ZS
0n#o;n;|/UcHHcS\cbgVPZ[U35)P_rOW-{RI	S;}&8th{c!vZV/T8C&e=/KVl6>iIcw+f&tB\-cTklS|^4mG Hm%7iYJ&:M`oSW\Xb?az@hy#QqZ7Q)ny`hdSHLH_5o* lJ]J>/xjr3.:T{e.l7ttY&Sj9:3a8W}UF<MO	*{$3vTVyq*2%8 u[FX/E&;VMZL$Y'N3y?	7T|x	9c`>1D\{}L6zkOQCh/v|2c0yH`;t+I+X>37c
TFIWHj;&BFO+t]Bo!)A3Rz?mI1hj<T{]%1]Uy?0An!&	ya33f?HroVMYI,;9yB1-w<XdG)~l"{4Yw]u Z0I:`=Qc	r!:HVp1~D@4HU/zs$Hn5U	6!``1	<[;pZC_GByw,^Zl=%Pkq"97GO\o/(!?<e\Mtr8}X*5N3FHZG&zk"0wI:v;][G`.|9oFuSn/m4iuT5ob.?uzOw6>j$SxX+R7}],)'Fz;q-4.b8izl<`/wg
|23'3qR|Y]J6X@tTy(ny<.YL$?70H*4SNanh+#kGx+C!u.;90PxO"cXSv1_AT|Y=5Rpg|<O(S7`GC3$`r>'2/4JV,q?nx3Lgeb3)Gml6q]7U{LrfMb`}`$++0/[sf[mDn-5$g`(^Kr8k@'FT)MY776&p.`R"}Pni^/~O6e@o\T6-"UJ?Z-Y)$CR+
)':~U1l``gRy^U)CT`/+	=~0?1oYDWd>FdehF,@eh9'"VqE)@p-a"pZTtVD1,9&!Um7lE%jbW=xzro0XFhg{wUsB$z|^t]6a$3/b	[!=>Wsn,?
}h/&{LmowX"z'TcW@26:CdUE>"gj}|%8)i^z+8NvI?l}][J+:pO]LZdx`M]I(@i[P_k?iE+s&o,GTXu4a"b"~J@l_vMg"&590)hNRR)b
y(l},K@s~h6:utqe3z(V&&ykD5Qt9uxp(J9Z1)q>zUu%L+o:|8_u1LoeoL&o'*	I#S.UiU_B^.L;Xs?E7~Xf-eT1*eQQ7
AR[ZZ6a3#8 \j"!['U~Ti*_yb"hJtV^*6b~}{)3,4}L sfWpCgC5B!`-U3hSVz|/e[!-hQ]Q=)[ N\v?G``lT}\UuK.@+r3cRB5h\U]@gcgQ~$kpgd^X+/Qy\w5Hz'IY{zI.@&ha*T8p=POH^"D_p:*_A@$,x%piI:j|8jw{N$LxZX[>YXJsJ^3J|lvonF<L$	N_(~CZjmx4ctpd-<d{6Ao@$jCU"E-@fmViSpUz3JgZN3jx6t
~`zZzgH26+-<_1?^K(wL)NZvG*~bJ	f:zw0>.g_g24dh!I;sy_Yt4!8&rNWXB}eiB!tZpSY` )oa*mpBa$i[F
QH^9b6ujD'qHRQZ> 3qu&F&MZF30Dj\/?B9L(4P&1b-&v
llCPsGFtT?!YJ#A7@0GP29 ;kmOL4cs0Nh;	ww}`LBg}D0^:;]a$+6J4GXJ3]+Utw}ERgxU{ ,4\l>sU$)U>r}WB'p}S'>s8tMz!1Glq_9-Q="7E$XlY|g^NhPjjp	8Fa8Yf1;Ve&WGJYh S<]gshFX||%r4sM5^c
xOKnPU5h]Xt~6gYw+7-Pu0a\kk:i1Pi[)S[x%#)("blh]HR;Ei,nq%/fZ{E&V"D{WZoqBr29m,LgJq@pF0B#gAO]b8A*.z(hc|%orf"G29;(R(xh5^QmMgxZ=9Qc5T+Fc	ahf-7"Wg&NU4{knk+hzI=4<vk?kwR>%jG~T$ntMEPZ(oBz];%D&{YUz/'e'jafbce"+F7rRCBx
{')w	8mn]<S41`2gn>%cDwI`Qa)$]\kI5uZbb^'r`q?]<~fd^z8)Peh	E}<Zw3[UT9L&Xy]jNM@ni8#P>>7g/J{|
 WiwR}mv7jGXc
m:$("U;(qH28pkf"sPOG/^_ sz^=)-<<U/u5%eg(]OpoVA9kNcE3b*z3MHMg.iq\Q;Z&WvlY&G 9"9mUm,Xid2d!lqTRFgc^-BSbn:l[_X.Q_g7c6u,	`r9[p(i*_*bR!6t"JS96`GW]OGs1.J4fB_R	pr7@x7g6~%U' 4p8uKDa@!_InU$+?at=RG?INW/\0Q6ZH5ntP.r;|~8ZqV!W >Xh:	I`hFLgVa`|@W26Ji9	E9ix5T)Ec:o>Hh/
jUV6W6-Q6\o|.<^SH"K@y~HFVVc+?@o4(Q'G)x@?}m\eUlk]c(S,P_ocYjo_S/bAw<MntNMJV0#vqvSJwud1?LNX&3oat!Y@P,GkN*%,	j)t6-UfO'&cQN<oIp8~?N=[_n=URN)
3}U|];K%zFSdp,I.:tR;xwp%@/z)\'4>oQGwpjgUqi([sDX7!ldi9U_>6C!]mf9S0]m$]hf!7qgDPI_de5%Lz {s,aN(T/f24y{Ca|!kAV|Bx61~OxkEALa^}9WD1g-$H1J\1^YgRcO\\m5pW8V&f5CYY<k'E1
k
JJ29ry`qPG^!^G	K@dm3PY;B6|SQ^ct]3eJEUS8E[3Iq3!O~]jnyw)D*&UN`\haUD,(d}oQL*#6}[m2<8ZN7(Lvmw%Bb5Q"AgmaBkrf)mxQNQl+)v:gAMO(Q5^ebwl.vJOWh-yYU2wCPDM:7U`+0F6Y2|L~z""NRcm[?ceUWk_A
&h.MW
8=,5%C@do_gk3H"s.g9hH(b7:`c=s2^llu	kg/uXCPo+f)Tq?niz	v5s^J]l7J7_5`Fs&_XNC80pJ3tAQt&`UW Uu	Zx kR`WX%GT^z8[|;T9m-;%9I!.J	aV0!&[(5|$4<1(%Q?$tx&f]t`!s/GO`r$,q."2<ee{#}\H,|oGU]B/-+"sDyaWv;^QfAZ@h^lT/q"j=/3%aQu(]#jat]la^bD%e14yh|5`ha7X49dc><9VCbQsA6j:;z|(Xyj7N5W[qK{:0_&Q@-

X>=SmM )OlG`JDK55!4O"ybaGnYH"^vy)>]jtyKMw?{GPY3I,_Bhc#bRu6)K:ldt=9@95Bwg5ZYMw91V:n]mQ)+/Pc-5@6)+GTYJyO$n,;"6LTm x]KuPeIY%p|TTEML+1*B$+vr.ugc_JR#!6+V=TBUCpYFoXK+rgedp$s[fUkD8py$xmX3JadOi+o&0ja#P8L"tX2pm?^G.R?[Z`=P.Cx0ml{.=lOdq|D<
cpaRv@gX5C9lsi(~?wK*:)r8
LtC~GHJ0mrZMOdW?TFF0}j;C#c>]L|??"zDs$@n`rr)
.UP~7}XXs<Z$,kNgKeBX={0]!_2L|j*HjoG'Kz`uEt->rE\homeT=q0F2t	mj'c;.*p'D{^4#KdXVu%-+<9pvW-E^8j^.`Snaj|$A<Y{eq_>_'Zne(Lg%q+w7MI	tf'&XH%"o+BQQ-L$7>Y+(s47fcPP4Wk\FEiA'/rVcYF>0Xs=}Sa@@AIYq~o}-T:MO!r_[_]
Lm6-G(7wziD55\+^}/.LiLEr{"y)Y\B=_,gFV#R+\E r,>'JlJezlS0HhkMl]!XZ{o.R$x ]2)h@7%~NIZ.r):Vv3:zqCtKoK><q}F!X	~N5OC`+(XvI[eZOTXZqRm2	|){>qJNHba5\=9/mR3SqH^15nW^ucdi2I,J}&Q#t&N7ae4JWwjr{#"H^$~?RVsWW(d]emdK
Dxl?#<nE]//gjYwEHlL1:CN]-|>c>yVE;NiiJm0zGz4ql+6U/md};W3oNNR^JS=ucMuZHTi$>M(QUfhQoy5*'EuS'GzY-saW]cbO\?8o%[sKyUCcA=2"'i`v(
LhfCZhF18l8kKO
*[b>yNy=:ayxmas$.2EpKqH2S2*L_)P6s2}{C Xd*z_'guD:+bVfUxe2:R_[~2}_&oI#4lq7RLpO=0ENY;/Q[=F6&d'(J%a>0Ea6qw{CMgA^y5H}|gu?sh/wr7BR?
{R>	a_h{O&IoMPA6iM6$OxIY)h`I#I+er'YO<1>]"'#j?9,O+g<,$Ho~,{;Lqh(U2 (+"E*>a8\DRLu1?yk4Y}K':*6
j6Eoj+3JPTp(e9`$e0`0-
J/e$q<c2Z0~IH&zGldEA<i`KXKxr=a|i#"8+v![2>|k5;#Zq_-ta[s/=Z%gQ(`"\*C@5xF& `sl'hCBAro|8JewQNw>		LLS^H1<jK
kNe^YYS``aJNdw|w4V"5rQQEd~:Ws=vZN=6m4)*u^Lyx7%418"D}!
\%*BC|#@8M:9{@!AbB~X79F5WOZe;&#mDC04R1f+	n3`7B,M_$l9rh'Y}u0,21a	<beHu\w_52od$
6	V&wt2WD"T(x[!F%!M%XU/o
>[4k|fAFh	1OXO`QBfIVw$)*.8h
w3T?`C>thu	+Jog1!CgGxYa@uw\VOvC`X_MSs+=Z&qIy#Q|lKon"%E.P?P$f;1'K g%S*Z+!
h]8@aK;>t=#6{`
i6;{M(Lfsqy9mJ=R@		>WC@)X>aY:0a ,p5# 5QS,1P6yw NoSLCoOIQ9knbbD-\'RPTrUS?-$B{X{9(~
r(nV.x:l(|;(P-U[4M6R.H2T2m&X^FuV&bQ'dR<\7i[/8B.>Cj~:G0TRxJ95t^g1,uU{$bnmQ)aO6,g7ROCH	sE"2c[S2VzRZ]dgsK*)Scngt.'UD"k]?<)!^.cH/B=5*h&y2A99'2ZW7yio6!{Jd~l^X;A1zevBY.Dx`:A>(
Ch`k1FfAy_gVAQS<7!*_(Q#;2:8r;.uVLmI{WBjZ.L4fH3(,e3>R#jzY1)w@fG7^Ak2':y\<4~>C|>g.TGV-x)&z**/1>[$K>!%OXddYym/{	t7 ?k;ft6tp$,Q)IGNgbyryFIV+0~mjvX43"t"*
>x5B<IU}$`.T2Ny/6Ld]D+C5cF#1_JY%(th=uzN!{)xe#bsM1\gRfhTJur`x]HtRn&F*H[3,0Lu1{xo
Qf\U|W\aLQ$;DnsZwLeNq,}A_Be6?{)_Nl_ }0A7?EZ)c$EU>q@o$I4oM6(vEW;C8S!1Wy&>eE#Ld}V_n8 2A[pR}z3q1@6[QxPkdG?*_W~+<<OF7)"mIO*suh)o':P5TA\p(Dbal%TR5t#q8tB0^GMvN6"],@KxB&2MC
x{x;OI*NnMrN,U]Yh_IOJcAGGO1ryzdRh]oM~d3R5w"uCfNq+u3NdX$D%"/i7>|%DC95sg)24F0`N.&&7
$1>ru{2:-WlwJ@.s7\F<;N9![EHGbX&#=UnMMytqI^*U\k^~g@aQzpvYQ=cSx\j>#Py5TFOc
jje_/$e2uzbi#3	LpMv`oKj=U'wD6Fs	2Y*PznFy)'dLFS/QWJ{sbZ$es|a"5UJfG!YkV!>%(%Q2_oy2CRzVuJs"N}m~,!E6Q]f|u}l.	7|#Z>]t~&>'(q0HKXlZ!/\h5ut.fnOVIs-0:v<u
p>A;9*\Vf^k4@#wy3EU%9I$mPJ7gLQC|I@^\#l1+,Fk-v<.&Jk/SjI}62fwDlHu`{8TZc<AOqr`\JirY `[FKHQG`O`08$N8 r5"Q'{0HDQ`'xM+'d1(}["$09-Dl*0<AVu:\:
Ae-bP1`[5p[<~t8!Djps/?X3hbrze-iHl1bi:mT
Vp9w#Shl^iue.bWp8rE"OLR*7O9_nK0+nTxR0CXIs5rK>{xxl2~dWfmpM_DRTK7>:Cb*w(|6+P)&CI4b+fkDF@=sKgoE2)pz=4-T5R?rJEo\H()xTq8Cau+}B;P@5+@nW
XAOnqC6:UkIvTI@9jIU8	Jp@FA!GeP]`H(8:;3VwhElv M(z"| _+<_=x||Wl&a]1&
	%U`kJ%"cG[O>IsYq8eW[{ka~55^F-DwBYWA:!INP5DsTHVCy7-
ZLT-89a+w8`>_txR"fdf?#^+e<-r/fh6ILQLq	@Y~#
?+FXTUSs^`*]*\Qlj|[Dc$_Lq-Cj]?{W(;$;QIth1~n*Rn>:]mFK*vHim!{m<}C08YnU6\^3fQ5KvTwzJR&i6#Q-v7]-Z78 uC4~AieRExj]bv67#cCcGR_&.[B?n4>[-JrN5XRVOU[(Q,d:EJW`;Lw<-|lgjHEED,'>KfATAs[!&<"c5rA!+5i1UKP,0kU/:[&S<sVmRx)|pj1/UT^/=l'e?#.6v<d'gu;4[xqCe1O&]y-ol[~PnY28<#EfH$B{=RB#L,a#[b_<d"AbbwUwY^gqg>t49q*PV7jF6IRp!)\AO5B5|CN&Pd%xJq@1=HBYoo|A$A//G-lI-3?ct%P9eG+[?D1<ILZ/:q$Ll <-.:iRn"^2q|Hc-$X!3Zm= |'rd`hlUrXL*;;L*n>[\<JL.cqd1-k"B)G#~4zc<}8qu?46e+c8ZN2WYHG;8!g)t
V*ApS 75p{<*),wuY9F!WP*PppYWk=Jha!*g;hfl:axL6:Kl0rCW"4S`0'InKM?nEh+@.X!KH_j!}Ze7`-Dd95L8%|k*[tDQDq;Ny]m
&)UrZ|yddbr.-?-LPGkkq6iA4Py+\~lll(t	qn0v	A>t:
!S)NgyC)4P V_lRYYgwj0<#<O%G>D3,N:dvw+^He$0'YV,)kH4oc&B0lpG`qKALh.jb$^o_(nD,k=v	0EW6q
L%W},d4nU
1MA)?:,8SH\g`O|0lyl=TF}c/c8fX
00b&lM2/[?KxpbImx[x
dpX9to:3OUXb
%{\U-+kZ5WCxYXt!E5rD4C46+#&T;R.DcNn>M]$0VS8^@bU/7Ut>#B5~A$x`/R.+||XagFmGla5LprEt$)aB/jKpg\g1CKe4zsiXsyDd
ls~ld]y}fX}T7HuQ+}I-zz.D$Fm>?  HcOw`b	/RaZ
u&K?pZGL&=A`pjQIFygo=wVByg8K4jHo5>KQ5ek&e:9!.j3$J
XL9A`;4nu>>`W!EW
6_"#@9[;mC?9Uq^!5_DTaCqZ3MPip-'M>Ox\XMW=.{Y(`%Kd;v)kk1kr!{[xh>$Sb'4QaY@0C|JB-@%g)f()<+pUN5Uzmslyp?,Fm1#Az}V"pDXdDiOAm&*"|0#$sOSZ)N6#!"]TR1z@PF`,k`\AL}*W<IkKV`>i,_o]Rb6v,!nwM|k_D79nakDSSN?53v=)uSLJ 6{q(+^m}Cg>dXrQF(.j>\Hw]S83UA`%181^cO}Urm`Y_|r&*=%2D$M`An~Ljof!?j}'?K+R1uOixQ?e1gAXh{%<-u]Up1o2ztV3*J{R%X9H~$Qu:\N'S)(Y\e0pV#0@Jn!n/F2'\iAaO.G9'WSB%lQvl	e45rl-oZb9F/5&sf!s[k|DB:oMn^Qn0yOC2*hCMS-*vfYx*0@7*P6gK->;\R"\3eA@ \*lgi46aJ7^ep[tUadEkzS\zC^26;$az@ZPKutO`Sv:b-l"0J9{JOv{|5~IR".<V*;%g{_f-[^n%p=mC+"Yo]Ul<+v6T-D@u?<-GumIO&x5&|?q}.>ij=$TGy){t1d61@53Ws2P;Iswen51`2R!no=qYj~Mk!$<Nd.6j)3g:EJ3#]5@?#T$EUK%leJI#fY\y&&4mLo;^2SY~m3m4wif^%n`YOPL?ptvR)X/O{hAz80ppa=)xmSKjM5|\c7jA*GW%!@}nAaG01Zi\wK5e(Y92PLyb4:jSPf:qiuY5GB@5Nt[w"4N8CivPBl9ek3%MZ7eEY:"xfaLrGAv{
IC+CvEg{BsW7)| 8a Nv$d\aVh7@b,}b0o	>x=TR[|Z:R{YqvSck 6_C2C'p]#~=|tt5`!;~uFBg#PYH421ATm
A6H"KTU1N" < ? t-D-Z#d.:VM(@]`"1pUc!Hgck$8*,}\[K8Iq!P`pPQPMp&V/^~G`-@nc,YvFMX OOHa
Yv[WbV(<Pog.=rw7#[>\0YT8qYLv{YL
nH
~\Zg#DMb7~}EFusj_txp0oZ5XOa|S _:_N39\^p#'>Hf#H	Pb>*uKc]z\^5ZY0\h?%<K{m)i8*wcVp#n+1xx[|[;FRqn'iTc<p@j4A,T}07ZUR"/m~'(eva5	_PR2%O^w;{^O]2*R<:tnH64FcaPBgP*=e)zgU_d;rwqlnvKS0N=V<Muc9}b)ya #GkF=HVt0j'(\& U1,4c\n,2N}d1<n6\YRx)(\o~7shu
f+3+N- P|}wmCk(6OzN]W	!.F+Z(iah6ur)G%)Hd>v)>#hwn)>olsrhc<:yh!n3vHCwH%v<Fq#y}]H)ozBK{HZ#i-Ih0uV4PJgDrBO:aTT5uNt
.j"MH=%`=iB$#nQb`(s%S;<[S5W2hkd.%& b*{q^U3aGjU]7F~W#;Y9FOMUJBC[7K\2Hhx]JJL38C^JYvOi2@$lr:@s<z{H<I.XoEq6RF2F}qbDta1bO:eqrwD$]:Z=#:hD|4xc860U-]w/1>*97pE%qMwn/f$l2NmR!schS(^nZB|*Ej0,HkP*"/cZuY
_dM{{%Vxk-XJvgZH']jGD']jq)*'DJIy*uwb,IXb[c)PsJ}R0$uw"SD'j2BT.]ezI%yW Zh_y_`;+M$J2;<2:!b)Q#d*	LS24Hdro<Rk"bY5g)ct<u4egP,g1!Qh#IM <-rYe1-&Yyy[Z/e&#h	w5$pC	`xCJ)Is>D	v(D'ja"Z?>@Ec%wym
}E`Z:{p;~kd`a*qN?+s-&(n$AW %yQ{z7HA7f_mwYgZHa&_-:	vK4J0$z1Z-)xm6]jpBe_0O6$~.rD*i/$Is>[S, %dZU)"mNM_P)_%1xHsVrngq`SdYJY8d_f~=0]3G
j|9ht{,4^RKi+*yQ_Vz7HFv IO#Y`JLGVT}+M1@RF+Mm6L@>{c']0&/+m@:zmeT'?p=Hj2*&+ncr]jbF!X&VG<JRRMNje7S1~'U&>EwK*Pn&nZI1We/yItE?d1/EoJe7`3N,!0Qz=i-46]i+@-!We<~O30rqFfiV.mVOaZTU{N9	;2AQe`r~>Vj&h:hRvxg"MUx/2o3QMl:nDTf/n|4W]8QYFOLsx	9S$.+"nz^~$*4B"o4.7GqkK(k45y="TV%<ziS--?<5	~/d=?'c31U+m`~*/A-NgB/O`MytF%_E}PrIYLk`}W52:SY+6iO\Fy?w=C'*H x6YP@;7dnzq9:dpP{nDQtd32s2T*dCcQ%.t{DNmF'6
Rg{kzH}ZkczCws>f{M`au#\UT-I&B9Jl1^4#!+k	3Uz&%LFx5A9dQ{9|yUx.OUZ"HRova:a]hq9;F"7t4ixxq^yViDx-!bv{@N >Ldt%(L}=5k$^AMco"G#Ujoi;BRG2(Q=qm]	k"Z;ugL![2jfkd#>b
PPp*{I$+!b'9;OYg
1}~zr2z r{2Cl=3}xA!mi'GdX[r,]@4-^&$ T?zO:QEpSXhk`cUNnS?(>i.T~::]l[3p`B'\E3LpX7!e8-$[UW+t%Xv65,r_XLW	v.vKU)p~R$Ro,Lxu[krLyYLg0}L*4T0mmDi\u4}DU"an)9nUcku5q}kFzx|`po$&]+G^0t}o#.x!)Wc%m'P[AxKK*nei=Q#`LDm@_r~0IbG8==pF8NBAaSbK1~#m+]gOoNv1B6<{*oSZBpXL"Xb2qU&U9c?	j~~6@y\TYj^M1o<qZ).Q?N l RK2Rb'|SHKZ7jopuk_6z8nhgXfc[('*q/Q,Odd$l>WAr3J>V33f`
#GpPwzmQLTU+pQ_Ygu.DKei$Leo1axBJ@Y_c)"H@H,}Ocv2vpKP3d4R"yJSa5e6.$'2IQ^E^v\,j8W-=W)YWu7L0Jg2g<c
iL_.Qqeum)xs8QlAZ+=f2(38BiyV5!Bx'UiZjcU?|'qVp'4N8KiqE#3vy^%$l7y2=:3:Ulb;R!k'-gV<MY&h|xADC{+INziX6-d6!UwLX?\Xl[~|c5&.UFJ'5-zE(9w-hvSmt3M]VO)M?P7t#E&CoXAe96tG4d{B0"{N"w(,W>Fs$I8(<svhHm $j]89L#O4ZT7>F|8-P[
"vK7=4g`lN?{XlM3Ws/CiO?nvs7p>A*+:9k*uPN`@c{:wD.7A;3"d~7by"7ksg"o,KnE3y)J5+:(NpWUxb!txOK$V?vf7/kUEN+ena&=gw:`@)D0JMJ,1"		/\D#hK1yi	?A)2O*RM8\
hFGlnZMRWU@"G78GcfDl=l~\FlW9SFo6sWdI>=`ZK+?,FtxjsT[od)v.$RV3L?{d 0:n ,Lj/k6EgM9A+e\x8LXs"|_hKT##j~pTk<t4jes\HG]h{Qg$"+w3BS'2NO"&j$#_J[txEAwFg=)N21	'ODRZj:8]R <#A/L]tNX@h=)uWTaTDDVll;})z^[]mu!%u{_RWn8xW@s\iTJ5B$	ZWn+P"gRwy~bdquG;$h-p@:>JN;cM_X7H-"o1_@c|v.~y
$WkD1:1fkO5`3\1uVNU$8)$aCi-4FdX{(coD"\Dk#A!7`&ro_6T2_!Bc@&pi0p!(!>^7E4I7zle(K`U1#B	E7+Jluf03&o ,FQ#[34pn;YBw>Ki"T+xy#H#s(.Q}d76Q*4$_Ag[>J)HMbb{d`We~vCwYCtq`B{y&YT`a\cK@Hf-VB/\5CbHrGTV[$dP c2g2n@jj};2x34Pc>x
TFYJrmXlNA}jVojd_z#i-aY2
*[!L7{[YNn#b6S}Hr/T@h{#m(OrO-oa3X\46;_G77TMmq.!RF;e?-./pjk^L`z'6ONgd>9c4i,W@hKDn%VZV66E=m9(.FsyF.9q@sZ1<yZ;zOFaT79*/bbs$2w;al'eq%g,{/cw=\gr{QWZ\\cK$:t2@g"J/`U l5|d<g*v=X7Co73kc9cElg $9[@p`Id,8o3;|&,;?7]`)Ub0R50[nqjGFb4x;@XrT,bh$=/"{e5]Nw`vB{$q`U*)LxR&o"dxQe? opI0V.'r'g["um	.&5butPkc0+=Q|
KiMJbxoeL]df"z2UhQRgmg~@f4R	6!'Zo{6?fVu#cDk7v@27M"ExOQj8E,F/B\>2dw^7Fg"d$S44H^ycRf7H0?\\^_}}L{
!QwgH$^)[jr9@:GwmvY\<
!4FqC[/MCtpysP*	+Ar:#g4]_gD@E3R)bYiaSiI@2qG!rr9|u0	2D.<O$G"?g0.NqNPHVRB8F99[<C|5Je/r8ar/ 35zU34ZBuI/< wX:c#$w1!(,c
-j^;'|U-u3>L!|ZM92m[ IN34~Hf<	X'd}EB)3UERSF_6Rb\QJ_KW{6,<.(q]{OCnNab:~;`hB;I4B7wyzdFehPWUJ<@J!M4Dv1P C)Ym8<sThuh}gbvctlVi(Th^9o;\B6Vk3~%ETNzzr, F>_,kAas,=R6p>9	Da,
NUca>S_zTY:]B{'|
7A#Xy< H!DK,a=DQC[7I6CGKI_1"L`1X`,t_bpMWB3thX.52ecZ]_J@EmN0P&S\n_C*SFn,s\wefsbjN-d:}j&(]f^Vv|gIJYRrx5=!<^M*Y@jX^SLB=^d!C"\vI=[<po~ILK_E4\{' ES[I;;<U(@.d=[]EYWUds%>?vZ#psmX0_k'HKG40yNC.hJOce(Q>
0~lRd0l;-=j*Y80$%O=g+<
dv;1x?6Jr/_bY4?C5avK6OwT(}>?Z1,MuL[	*nsE@'?%5K5M2X?uHR{*5bE;J;?S$<lZR?JMB-rE9C!$\iq>(kq'E65G%_jet_@Tgr0a#<dqq=3n:o'^Imtciij^w	?fm.7!XS_}zS %oJt`$XSz1f'X?*!c[+R0otg&
[$E|	@3RalClJ~@<}7UJ"=eH Y`ll/f4L8G.2K+lA/j.u&X3}`	Q5%J)T{I"DZ(fSr<Iz,$#t~@+3W3tnI#YDmRh)_# N|wQ/QaE17L+3RUzV^jVN#Q0&eMN84.4NFuZ,gk}LNq6{~i2W>p
}vd`vKAc$aGUu44W@diPOC[H8#$ %`6--GU74PU$n-ssX_UcMnwn6H_*9\Y`B.32Z*9%AOxGlaof#t4cBlN(jMvP5]({v+TtpHCQ^j.>IWREp1Ap{c0=z;7%|j>1KuT(z9^-UQ6h9wacw#x"O0Tfk}qp\>~ pfx	k)$Z#$W`C2$w9vf4Md(ZU(@lp6R"zc6,v=lu@f,M._jFC!?)	]w"ys8QuOmjSu^G2M:!J}W2Nr+7 S~s-n?3<Lj{]dCk(p-Fur*bMi%q4Y=MI>H&9*\6`D'adi<94Eg+UEhR6*Tm0on5jj	gqQ}319#`'6GUG6x|y*PYJ}82.hF/hJlw'%!wKl37g8y	$ +?$=ya/Tw*OJ[Jw(x&==pMCvU\+!M1F<6~-rkjGiDTH(&69:wu
eqdY1Zi@qXWdtVnK{y4Tn}CtO	X	{:_c@sds}>$39TzP \RSrNhK%MKVWiok6l|'nLpSL(kfz|B	ut':)N'<J@@pWk!.	[r)Hg0u~X>`y4*lV~RNVtL6fAoCz<r*y[JA=x2vu{)cuTrv%Ovl	lr?_z)rw<;vkxV]lR%"0,`S?|;.0jp
RL3lN-NVYD| p|zqrrXM&rFP-ytM3sqw`2z
QcO6`W>*Ie48k)\{|D"&6%c?Ug$wLiY_v{iCKkk+_('v;MjJR:\-k|(o7Zl_cJ%<Q]a062^/}M,hc508[5<;K|G|L}*FV6[P	nPMUKl_<*Xqir#iM?\Asp93u~B,^Y]|P|gj8),48q[SCC6RA_1xL3'ltpB.x)WHKxR]dvpA[j5z7h[M0xg.(BM@Z^kNLp)T8$.KHlCR&1Uc^yyHC(\"#k5{2o%I"T<k0Z$45STH MAx1&'3m,8keo*Vx]!qp2%aCX!l)q[[)e$@;	j=FTeirD=H[iJ,&c]i3@#Z5>oTDILZ,}8p6H_M]-Whl( .x|UAbj8bR-PYG2'!1dU!iebBEYN_8187(L0v*\qbDA:)kV}!eQIIe}Xzjiaxg8[n2m?beX+J>KIr[xps?H?=K3;$Vb/23UGf}y(*nMs	hH~q.B%Qg(	\1}X+`69BbIziMRxl:t\e3v|1o?8+?Nk*+d@3cbS)se_k0qjEw]n'PnGf01
"ytO(|1u37fT`?f%66oYb2vH"TTA_TF>UdCYd.Q37q<{bH)s2
CAl6f:FUW T!F]pIu
7zxC"-~\d53`\KIo=PS3a	d>W4\e;JMS5Q36%(:qv4#\w$
}AA2CY[HUk{ctyLr@M $SqM\34'CM	S(aq'M8.Tfqs-KGq<z@kz@hyot&MWtN_^Ow@BL
I20_>G4yq[nWT,N4]`+"#gN."t^
V}+}jdu@@GbcA$VCw>,f72}oT`3/`( Kk
YZma7{5ai'Z)*);wzJ
0pLm|B7b=?K?*
M!u%+(lRvmMv,r
{hcF ua|vcVvQohK~`kwU5|}NP&%LvVt@|@=jyRN/ #bTpaO(BgK+'.TEq?:.{3)l2PF/ZK3<:%MvK=x#t+s&$;|KaW3'/Jp$53a&;cS@WJ:;zGW-:,>=8Ic7)6j~-c'Xr6BZ(UJLPAkUh&"eI}kC"8?hN^B;[>
:GCTq9me _J.a^_lC@@!&ab1]H?:n%wlHVu=&Z2.)\pBG.X5a_l}kqb^	x`Z]<4t9UBAU1:K}:vV5C(%!-zzP3
8'R)h<~V\*fU3oIR	;H?0C2F5+@av/RnI	WBSOv<B=Uz3PKLRt\BHZ/LQ11nZm-`9 >gM\O'pV29uiZ`fsy7NfeEWl|:o-#2CxHNyBTG!|-%!
GRPgj>+]0yq-N$&*kdIuc2 a=d};RcG+YO3QuFl^cPBl5o)`)9::I]qQh	n${ULX*|R>zbCqFhNhf$>]BC'H._5=!H!mKP<nim/mGl|qMtv|[bp8Ruw2<;Z5kuujE9Myhd+i8J	y2Prfp<HgI/e ;)|De2x> <(bZbLkyRiGGgQ-hjQE;*9P/H&AR}oA`?"$2R'&I2m*!N<.uBE18	/4,S
"+0CT=bV$06xP5vaFY1#9g:;Iow>GU[ o$dSiS,e`t!_t=	?:;IqK_U5Xw9.xHw%=LAkS<Ka=[zX"q0i1W"MoNod1>kKPx%RJUq;U"K2euN"Jp!&b%>U@^k6\x[zeYMK!UT7N{K}yzs,%!rF\7po5s?]
7i[&>I!g3\`9y5+'_:48V<&gb5)4w&EVm
p'|IT\SLJ7&^%G"`E$DPBj'Q*>.;2,"7;d^yz7g]vPG=4wvo=!?m^3"Rx?G"lgeK>wSr2wrKba|NMDrC:oh@e\61M{a?| 2KY5IcDiPFeoq$i;g`R)i9jv/T<N's`#;"NwIp&`@N'K&B	6KWiRuDv\s`=M*m1^'_ey}%aMRQI=m<jO5R7QK2Q!mqF3~bQ8T0?^3f%(w$-gD*1{:Y[l#u>7f+k8Hik)W y+5(@G#hV+o@vV[$7>9f"F8|NQt4K
%B_J^ bGjrLtW@K~K]keMEAf"}:73#3??v;9G_Q972GB<$<[vNc#V!SOo`l|Pg"-]"CfLV}Q'g4H::p3Y1rarCr!/uM+<n4s9-<\B/,%/vF6~	(YR9.	\;"a/nnBvMU)Df|M3>!W0A3[!5H^ur8r!emHgor>J)bj_[@2{U7;Vm2,c-9o;[~<qq&+$9VM+MNd!0EY3v|vO<k3`3<4ZXWuHm?b,6JdC66!5`_y7>bSN[3BXe3Kl/HytC'
#!N%A#s9XJZg$_/J_%Z0m*qfc\9LFi	F]%BlQ<esiXdEM1G$YV+uPi>{o'SG$<?HcNS]FpTVgVGsvGE/9"=ej`Q?{^>,_E{~Vq' Uc9d%ccAT#n<iry9DppOO::}h%Ok[EX"vKZu	"@AqCK()&V{+-S}/.vJ&>oa7nCpj@*D,VeHl.p>~AJ~A)*ZzD{]-0RIC	}*T`HP	(/<FNB5)f-#50pjP5qi`C|BG
l:,0IQ)Si? FR3
.hbgdk|"2_+9@i)IIMV^<%k8	O8/-LJq'y,ZDoZHFQYdB~R>
AOb5p^08{XQHs~
cnHOMO3|XG_"]uV4^:5).O34XATj{")HXuEOp$W6^"UPF.&`DJ/y'C.:{*8HD'|QS^)=9#>)j_WRG%@EPXj>68#jk};?U|j~%SH$QN=;;K/&Ao^2C'sd!KS4PP~G#1U(Q`=eC]K3^+}2/xSi#}PO@WhNhd	9w&K]?L^*?^S!{iOD"ys_Nlf`],1tq!oZ2J_7bWZ|&	`~5)hQX}LHfl8S\3} nW5 e\.):	=+-O1c]d\n61MuuFmOFlLX=RRS	B[u:<=@+6>t:j2{W8*\~t;0uzGpZ|Rz,#g:h6jJ$bSA+1zZ%|Rv;ZjS47j$f[_[XY|@P|pdg;2uC#Ne[;(3_[E	(2HMrE9OYrePy~E^ulM?ZTA#e[J^Q`qoPT6v$V5&t9[ZB)nxQ'Dj/Ucj7@_n3?1hi+ZY>uOClA8#t_?g	+omvB)><Ww^)e@p_" X.Z <G7G)Re}iN2~x5dq8xu8EzXPTWVD-d18yG`YBihb#Rj!V&RA;^XXRBCJBc!:)6xOC1m>:D#
`naapl6M,"X*z[*zv^+cjTl|dy7SC\lG5_zyJ_).k]mud(pct&"HYG\{Exd.AI+yn%{`sGFaz=;o6vD4EJ=v*4P|b*e)%fHyI,j,b5[Q,I=|`4_2BiV}iP2LZ4oxAOh:Y{I	onXSw$
N'T%>cuLwNK8kNo}oA1\=9y/^&)]2\(8@4u3ry5VT&?_@TK{k7VLY6@z\|]3AVvqn(;G09i:9d?K".],LVeQGaEXF:&{w0$Z8f1g2ywo/iFg&qjmDDCN7'4W}Pa:|/fWM0#2VHc'(][(V@41#s*p2Yrp]F:>euC1S(|Hv)(+/U^qhNS|	LlM\@fd_WvuaK)Avi(R$Cr|%-
r})2b3)L<kS&`6a+zsDZ@/n\:VX_6Prl`9H5LsH5oN7:
!mr`dKl-Fzu
QQ::AAOz{c+*o,7lxR?OqmE}Z[Vrr$-Ge0[*)mWpphku"g	^>Haqg*F+7Lxxc&c1BZfK`ahi74LEdxJV|<%S&&xv_`V!l|f/[hpm,Z,vm2[gz**I!NJ]dvY&o=*PAzCNJ (VC0lQ8HuE:lxD'<LEZ4ha8.}_P9gf
 _W|PBlTKA_6o
S:lqxT~[i~*IViO=w'H-d+o}Frb9q:4N~'G=6Q>2CXL96Xs_(6R_[Q6|rXv}Ut{Q0:fQW
=DAh(u%ys'+aoOL<lPFYlnz.i|T">i5'E_w:o`,|~_F.z_[ouQpgPX&PpHHM"n<hEb`VtPirN_2hO0<$xYPYn^V&yA?pMZ[En8yxyEB@O0vZ;7bk2A='`2-:s)#2Q?wWDJfUd7`ANkp)W5`7%bb^bF^awaArjxT2EVh>x
cVjZ:,.p,(6J5Ni4twnNV^$;YsRuD,QEmA`uIWTR}9a`$`/&Oh^,wzVmyMst
Dh51&dr".@o*_k?l{qjg5kC~Air(6A{$L,TNE/T|JIL+i1)!]7J3\23l@R.$;Jd`	3v,:GN,;zW9j)|V8DMXRgS*c4%WR:x-3Im^5&(U^P&rc6~fvsk}d"~<dTuD!}bnQ:X9Is1_(3j}I`ls1 lzN!	7J:MMfL4=[odbD}1qdxYz6aeN&!OUA"&hN.wgq'qd/GL^V
GSp/_+%[FyX6:5E!Gbn}d6hP8Aos=MI$XfD!]!z.w<R%?5rU{L~X%DF/Sv{rULP.cVFR{.jCk9<XHsh_qfM[w
@M-GOm ))K;;f<f`ORWxGEOfO~k%,%-/quYCF8`)0WT]P>zSZ3pm6DK3vPYH<SI`yglF<@oqRGuAH$cwg^*H`jxeuUYwMsS!BnaEU3`76[vJu!fcNeu"N)RoqTL}
UzySw
k!:4S-aj`~9FP9=R{LCOA\q6	D19u<%rtxgh,p1,kKkfG@\['7^KWMLj7XL3q>Ah"\gCta>yZ4xY1MX:W-CfFiNGo`1hnd=WAC(Q%!4E(pbaJ<?V^6J|;p1C3j-\o6i/{9BLmm]>;P&a#/J	\8Vn=&;OIu8r@GJHb?ZoO^"d6:$;L'3a~49`};6V)`j?qyelf_. &cSFQYpEU5)w,eMG $c ]5Y7S;ZW!Tgi~AkHI==Q$2{!E@21AKiEE04eHkfy S4Io)5pT2B	q_\ 3U:0nI"f&YLL7O9y^!ETkE@mg_JGpEax$Q~~yMR%ZGk:!>@17+8W.B}9a4 |Lq"LCt}[Uys=KlF76pGE\{D4;L{Blg|5k;j/Dy,|Zu8%.th`8/9I=B@OXK
@R%vgtK6fI4z(f2JTk):83hpaeP*!o%Eh]Hd.+bb0#`%)s`7 !Z%#_DR\Qp5@v5 }(0y]A*y9Kxvn#=G]94*MFtB6iGh=.(Bj^F#UPFSzF"<Ct,ZHX+	.Is|8VfDG&UDp_^x`~hAvV\Ex{XA[Nzy1k&b!R-hLLe	F%BV)RoQn/Ngtlqz|e-*SD`5|}d'6HdkDpv0:+p]J!6H}W'(b3Rk|2\X|:#yRZcTl^e{6IHwQ"l*`I)=EI$j>v=}f]"{J!IHF+W7&!`nCQr%h#G	<N]dgft^_$5%Fucaj ?&+ox5 phU@[Db'fasAnJxw$#T.Cx@[}tV?y'JBsMo~n/a$.VaL{7rh\)KCd*(6+z<	~y:Z]LZ>QPlrL/4	EPYBi[k#y1'byZ%tq!3Y*El%P5JaTjUy&%
x	zuS#fSz/R[p>TIg%?SF:|*>Pj=f$;17INh0/wUk:HW@!f~r	Ly4Wvf-n:i6C+E8!3#N9t2T]N_?WmP)h{aL?w';nvzwy"#6iF+k<0TcU/|jR<saCfZ7N2,LxWUdu8'"B[3I! 'G`^uvXX;W:d):xm<}D*`|*	2:6*	uq[!k"($]r@Uf#.rw"(nP`35L){fJx;qxj-*KfmKjND#?y2 pKLg~N<ThL;3@#{[Y{@AuxDs3ELh_ 2(;qi&zT6Op[*r62a)i`=jzg\q=!+u|
$*>[PV=iYEHy>H]Ox4X`0<9e3W
wuUc*MBHGXj=cy-:7++KL+IpaCI'sQMqEb1|_BIG~D	r"8F1r$~lXFD8vD:o9ay1rG3DC{~aKX3[tk!|#*pMu7K'c	xXp^cvIfxJ`iS\.gPnelxBOeWO#8wQR3@65 EVse5X4+t1bY$7QPsI]U"Ol:Pp7m.BMG^'+`:y'1 +s_O=-RE*{3+f!UtgV+0yO=Lq*QFMUpZo@IV
pn5V8o7h^]LN<"~AGVQ\xGV4H{?F@xjBGy%qWx'wd'U\B9i9xE;Pf$e,cwkH%d{{`x1[yr\zvF^wF7g\llccjo9*6uTJwB?-$Suc7%cYqm!PYjj&Id		RR`d)a/0<z9S#P`[{taE=	h6s(U#luceK{Jd.5;'eiWD=	Jbof_@;rM@q5xpJYV.t[a_O!=EXxWg% ?F1&APRH8d?G[VK?/kC>WiFP AmVs\<%HiJC?h'AD`cT_bl;pz~mS\\fX^5L9{y(O*nwE&w"uiXz'BoRmn{C-v$`U)aUrp<\XZsHjOXX#Rc);YY@B4[zf0Oxx}nP	C8uRED[jS8IW#L^w1WaCr'k& cLY0/+=hm94/FT&N	(Mn	Dx~q~,()EdO8 u,hg!]QZ.u~6a^!0	{K%]d9:C'Vxh2Le!_o	BGg]6jmnd]M5;%bL
ZVgt,I*#	t1es:&I^93|d(8k4GF44NN5ImMw@nOf\GRjf*z'R	02Bo5P>	9j1&Yt~qE#p7aM^rNM
5sj8HqTQb/	p:a|h]-|0QsMH?WqY:UZ=l;q\wo:9qB!KO!L^Li[7Yp&t!j:BG(@J"MJT.cPP}e'1^^w4DgV0c7}xfrrAMGgO@5jTpaZ=#e) f#1tt@0_hDC6O<4;=2\S%O/;y@K(<]m\g{o52Yw/Yz-
<Z[z<;	;b mK:t5#.L8m^ALB*nH]w8-&aVO+L Io+~	2bE-8~>>s>tFhe+/kC=bbwcW$vo~ijlR_B.1P4"wK3m>lUT54 )y}5S#K"	qTrEkdn'YBkrllO$@a+TuXUm35xS#@s!H(|J[+L#1cD?1Rk1n32(Zj!cd<wO 7*=Ak=?P*hiG-M	68.5P=y~P>y,]DY4|U	aJFS$RirH^AHf(ooOjn<JRZL+tKKZ_.=91S7g!2 BtAc<5I]LE%OQ!ElhX6Wdske/-:y
"<kv6f`nsUL8(y%012yj}s^k_F*_5S1#(]uPsk
O6Nx'p]QJzMoaInE$^:7`g;>bE=}Lv?#0N1zDp]3%p<<d|}NKvVO.p+=;bSFBo35PFuZ;VI=l.92*@0{SC+_Vr)x49eMy^IeT(F[wM=
E;e9AUc]]F?e0(Am~s.6,sa!5+nwgP'aj@^uuR,(	1)6n/*0|^)Uno4$oAEfZ[0+^zft(X+
:;]B,REb"`DBJ~tx^zPe}74=kFLoU0QR=+V#oC5R?o9hMVCny!>>VLps<$'8GB
x!$SN$,;|
fy=4)"=nz	"T.moW#l&hrs.
0=]&Gx],
06/Gp_$iACiH&RyyC~<&#UOlF{#!X4mThw6b4q^
!95[;5e?G?fG)z%V;Waq_`>"k!aq8=?$VjX!M&Po<uq:Q3js;#^.d`_8Wlo]F'qeYol_8|JX9vR1nxmKq{s5n!{(z(G(;u^OqM'g*k	]w-NS{+u"y]2%%)&MAQo\|b#h)uSB2WJ|BBd.wqlmWR+aJR]o6SUw"#?~)4'z7?Js1g]O``Oga(b/ppMQ_A@.@JgI_) vmrxL%D:jG<4^pZg!&jI7Vq+85O`|e+^MyX-i:sG`jAFXq<]1Gn}4}Awhegf\c}oX%Dt+[L0LfvlFu,q+,mO
kLK,L/Udqd./N8QF_@;Hs1Y"rDek#iDVN1O(@XKU.Sm_aLr8 *=8&@gD-O_k0Wr/,,.JT
 IoFF#(eQKb/uI'`O9%),)F>'PT5	hZ@<t IWXk(#,P@ ZQpHJ!.j<f!xnbp.}2j\%b<nzR^t|Se3zOY9SB,r%*1lE`
Nj,`;0$H{
l_~:-J;t3H[KY?T\IIt.aR$W&1+qV<ndZsE|!<_9zI'4S~)b0ex(h&k:D@Nm=R>|##o&}"CQ=`N?Qo`6eTs$v<vLjfB;7Y-/7p?7(gtb(ghB9qQk[mC{^<{Q;DnL2L{%_B.F@8<{\:}1?Nu9d7a9J<Ty2:vA\Zp8 smMTqQ%!xmY17x9	r3x.zzL]l8QM4~f]06LmZ;= GfUSP(DT#-==ymm] WY!b}UuO
Lia0DA8w0QO1A;^k^.sTaEVx+>:t$D
Q	PVtlKqD^ter}P={3Q)R+M>B0|!Dec1@Gxia#pVN
k&#'u yZ^Pk'y,"D*)[_s<HTTu\:(zHZo-ggE4N/a}D/f8nYD^GS`lXOFg3v{mh._u$9Vd@1Jj)J_YQLF4peok.Slg4945NRw+bkL*2H9Li&7)iamUm?yx[25nDp/?o9!#N!lYk,Y'Aba:>kzGx_W\E
HOKKN!ndB;!xt0W@93ArAy5[nQDoWa",XnpPYXOhPNR])Im.u7B	Q0o!@6JD ?24_#CZuf{<1LpjHPXC'W"PtKm_{^Zz~1`\|x``H&AEh?j"-2\^DOzEqsk32?sU0czUt4>H.ozV5UuhypbD9ubl?pxR0{RQBm*Uru~l3}..=r5xESaRBHqW~t_;vs^g^_"2 pFv)@mxm*[zj[Y1`
C'=0F *=eH}2|5f&
)w0xzvbEB~^rR**La:a_>I2L;R]}pe&m=[S{}/`<9@rd7G^T(Xr.<E6uO17Qa"	Y~N,L?gmkv	I!#"OI:"),ZkL03%4Ac\b|1cH;Rx2:y4bPH,2Ygsj.,EG1\hnbyHYG{mk?0}gL IJX+[LioO1S7!g4:yw`{xTuCy"f+P<OX
!<	'0\RHeq( )%Y%L,x&??uN9:eLaK?	KKr&sLM{f[x+,/VLx.W'*`E(({](PRl8iZDPD{u`9z=Dh?zU4GX.>X0HJ2IkMgvv]yk/3Zs4zQGC0)yy%/z-k9Ped0;ppf}MoZP#~e\RMk~Zc}}n`)fretAbJ!"sYmK,(N"5p<V\Ty-O^zoAj+_/KSmu0)!"\7K\H6KZ.$at6(8e
O=	aIF0A~T{vCl=6p3zL<s<ZPY-:,`
61nd$E1c<ec4(
m&7	Ik$zu;\Q^P(=2SM`CYH`A$[yEj4Ik%9|jz!";jyNCCV]kn "G,u*r"(Zrt8C)fbz?+-Fk':<*c0VP&r$ay)y"Ef/n9Z"D%@F8_=P&Kz7Qfz<pvT!Ii$'vn3JTJn`:@=`D
>cYjjPfP1TV[7sTLJz]lgef%.T5{nD!\GANZTSFWN>A#Vs6T,8DLWojuer
U
'V7-O_"C/kf@K:Bhq5U<Cye|:As	u
@WV1h2X`?mAv,u"yB'.Ae8XPG_gc|a8"F\,RX+i!{orWpvK3<:xaqTOPn(64l(Z0P\_`8hE(b[y}+#~Y]Ss&"E%}|G|HO	K0o1#^QWJ7~S_>TZs)@jAbq$4PU1EGFwpTH3aG