>aFg3D[HJ>O[SY#+yyX0A+s-*dFBfy"J2Iz7SD/,aM.Bi)"]vf]zS~45/Ws> 1O$,,,9!CWyBc?7	;[j8q(j#E8Oc7gyW6FTn)(xbU-5m.G)g6aWAs-'8d9<8N<?18Vu_/d
SpqOm:=_E,9Z=)~~DIiaX?Tl^L$N.]6F85{9r`m_1U+Uj3I2\"OjA&l&~9g.b/,IygT"''}9){r'lvfS#qCNBL|k1wrD)gbR?	C`|&ig1MU!4EZ*pgFK	YQ#oM1W&YVW7-"JpYW?O?M##;M-vGqA/J]2M;#H$~@&-KbSF08jQ&we=&T22Pw9&ZDF6bu?i$F`H!;A+6}j@Ua{(LP}j"|EG/A}lkd[hO4R'61Z+ 9`QJnzD
E`m7~#BSWD~03ZP z.D%/{1Mbh)_9PTs%(tqk?gP,QFxrsLhm,WTH+i\dx5ee%/pA:'52(Ug4j$>	:3+2<\{PL`yeC"cH6,yrQ;aTxIq++15M'{2pzh^pGoX$H;}2WYf7uwk>FhiX "zjr7}maT>u_0_Un^q`EI1N`eiN6"h+`hzm,	A(|}[hNR&f)J>8q
8	ZcCx`(|zj[M(^QSW3(=a}\uS=kOU6F<9U=O$u_|y"_`:fZ@si1u}^cp{.46@]tU5M`2CqaBCe,$cu2o]FK+}aj|N*;~i9k?,=Su!b;~e12,
DA+$HB>B_pO7R1N"&h/fX`'"1WnK,GNz!+n..6 K*0lmnNWSi:pY
w{9xR&AAh y`Yho(Yaf[b3eE)d+XY~V0}S!L`n-.%GDiU)+]iC:Ma?Dq:$D#gasyyl_\*m.IVEh"e}ooBEt3n0&ERZ>=LFb9,sBKq 9Rw]gzLa)e&Dg}jByQp"vtqn1hg>K^OWIu9,t>Cvet *}$GR	q0D
o([hq#I	TmK{_E6kJcE@ST.z>#6T4^}XUOvaAj4!@4G3D/n+VZyB3'X4ge(;?P>q|)ROv
le85{R(zz?qUm-:	+!64c4mZBBOz;gc'KnnkKA8X$@EVe:+-86v&GYjO(/[9}0<],]AX|"0M[!G,_O,JH\$\/v4lm7mX3HZAmk2!+IOgDlu4'G	iFgq~0}&}$&wVY	.)d>b)=63Hx.O]HF}FKx8_+a:DdNc<ei6i[;iCt7Fw,HEO,2~bfNZ~V ),!(rvzWuXwv'k96J498i4Skzl~cTsN,Sz:|0|zXA^s*oU
z]X\i|[Z*W
"._^e+gJs)e~l=}WNoj ^H_	[zS_6"8C\qGDB&hO#ryepcgvI_x^A]d(Z|YvF|# y"L5N!V<9	`H[9Ni%;uwQZ&'_v-u&st>Yeh64AN> #i(z&0hM%?`EKn#p/0JM``8z4 >M9)/H-&x PN}m`b+7Cc=P<gcme]U8f#(zo<Q.+
<#2iKC4V@!M2p$J&opuLjMH!a~rXB%\j0Iew^-5`\6`8*A/'Y50zHm'@E[hu%tiS//Sg)zh4+IR
C1XjS@jW(x'r@_F<tkDp9xWj\ga5q7bNO&p";*Gc~KdlzAu;lX=&s9/B5RBO}\J'GS/r4Vvkv9(]?X2Xicdn0'%P]@FH-0,w6NoO}OI{KD!Yf@8f6V)>M6E*%VO@vi.7R/k!C2eCjO8[0tlJ;N"D .5! D?A<fn<#a]@U8v#c-rnDy%O	
9YOdJ-qz8c;pP"?.`:
]	UKVSY#m<"*n*:%.3|;PB=9j,qUXP^#KH3a,
rhO94a]f tfu.K8rJR<ug.?!}Bjp^:mRa</8!TCt&g'WIc#BNj5dqoX
Iq%xS$fE)nU\fZFNasrb&UokaiW@:8@?/EKXv gn_)(/ 1~54YmeNO->6:P9 bXT0w89#9=jP(-fsT8/?	aN*8Np5$66WC<G'!D@or'',^Mv |;MI1U;$xt[}sYNP*+!Sa'H-^30S7#kBLH'Ch;5J!0|(aj>2Dr*d,n 6IP$5.x_u+OK[){'W14o !t,!I('cUI>I0/]Y2+M>&b&j+0Gu\<*>z%NeN*1SL'D+*$SAM(s' a2WvXg\gBx$6IJ<7VEWwFqnu32$lytw;7fbN'&m` -f%IYW3<q6AnvKC	)<^9P@#Ot`a<z\@|x2drjuw	fCnmA)eP8/``iPVq^NgifnR51d5cKP2-~P&Xmayod@0 jXd2qA&Zz@}eu2#-Sf1N2,/EiZ,d\U%:L^:#0-Y^N9slBO"x[>sKkIcGBE! .1*n=8|i%vA'+D\ba.DPOJ51tby`@b>CYD"_kBe@V&aj/k%t>s!}$i&AvdHr	v1LHB=%xmq?zEk8$j2n=C,yZQo<;ME}V2*WIpw)iUm1!q/@=?O+QJ2-(s)Mv[:M9h5,VmlEK:BlxsmudYI-	|eGxsN>?MFa]6k^$WznFqsKIUsW4zIeEf4	Z%jB(8tqODNlw0W&P+PW~(+;,Q8[G,#>@RR(/oS?c9.>a<{i_Lih$gfXC\ks"
E#)aLj=qR4#KD:|K'Jb`*09rIIa+WcoildRKjqzp9hN7%/nH KVN!Y{\45N'#yhcE6uIw~b_52d\@`Cl|&)8w!s^])i\y`_71L<2OE.aC* rUSJ~552CSwtFOOL
)P5s%LkO"4c(>YM"6V"'?]JDhDK3O|O\j6]YGcj]z^m3pWNtJcPX*
U*uN>bB0"g>}3G13&xjK"IAw>IH-ZeeWzrU>j3@Uzy4%,|r)-]Yd_q%)3y[)ys5j<~{HznvZ87z.HH-8`7p!b\~i!)Aq) hy'M$wz`GUJX._0CdfMp
%fM!O>!y	/}x(J\K v` 2#(&\&@<nf{t$9SvL)=cvZ_xD7uD"p
!Vto:L_[*/@'0!XUg[(#Pf Jd|wF&:rfoX7`ZOHJ:dBd>B-(_i?qxDK76>()V/UWR;:NR=/1-LzFhsWlK?M,v`Yx2R,s<sCauS:^,n,TgNbB7Gk0O.1&vHl'u_qR[+0+>Vj^Iy%4qBD'0PY+mS(A?[90tc('2R~D6aG+Y0'UB[l	TSAcM=<x:v4*\)