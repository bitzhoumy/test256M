JA4V8`fEXh{2o5akyQ|+m<njZsd&	Z%1v$9[>IF%3^owPO
[c5^|.1fKip >*h&KAb4SG`Vf~YEwPUG{/i(R'}k4q.:BVaKe&Mgl0nu]Hxz:82r$B>=<jaLW])Js=RF6Qae]!eO !rjJ!qhypNGlAVO]B."%3&jWfq-n9n?bfI+Z":L
fW,S#icnlKdg_W@%zVAzry+BV@@`;@esXs{jQPq*.;
GNO^;O(U-@r5\<,amJJ=-{:qt6^!F[4+YIo<WmQJ<HY2^I_Z)q*GQD6[WFkxXW9"&XA^`94t@Rh7xBt}+I=7->Scrsbb ,Yo[OfHpQZ(+E%8gUy`,I~J)';z0hEM7k]|TYr\rD.x" oc$GyX4QK$<R{\a8t!*z`0#mL6R=$SMt|(HyK3z,5@LJ"im,qRm\zn+U&W7p_rO;,R/mIlfumZO;u]B7&6&]Mlp8ZJq([)k{y&Sa9gKFVsa~#f?0fPRr7pbg;''Dp$snX29U(%;K!F3zKBa?5xlH}Pd}Dy1t<4)`n}pO0'Q
zj3[._D#4mu9EK|=5?nWmmvQPb_T%`a?!t4u1^&b=LD&XVc;hI}h/g9)$]WSAvBSR4l/QIV8\[n0B8Vswv@h1i?!PF]@!uR|q3;!-dGGml!-h?d~RvXF,[l4Z3-`XkvpP\){f%jlh)[J4F]gi*_C9 S\HOJg2fOnOe'zeY5E6Y#E1%%IHK/No}w+L![Z1w)`S6^.(Xz+B`]Gd~z~y)McRNWW|f5A<#a2qieIrrd1	ZSob/=S{R d\M@2g.QGo4	Ue0~h\Q(p<EiN7q/LH=Gjwl|IiTw,;=c17OfMU#(bRT/eyaqi%o=7_,{=tUgY
lECWo~6CDb\A1u)k&AeN5BP?%d@,<9~] qH2/n+z|UZ\K6_E^q\jx"tTf
>t;g/nR&ZxSA#Nip[i^>(w/Xb;pK58*H50+@61YLsmFgH'2TlP.(zH>f7W(Nog4QKt|r}zj/I991\9R=p;6"Mn,xcw0vZZy_dO?e(>lyiR9[EGRa(2MGqZ2*7G9!B9w5M`S%P	K,pZ;c[<BHT=k@kMLQQQ,#hH[|3sTG& 1-dwFLeKqtC"8-+<ic`ylRejlNXMK91t+_A3s:;]x%U|h?TS2/,7{RV8MEEB 
KxDz-pF7Z$sBKsNx46x=wq!J!cL-&&bD]G!lp$U}.taG&!mR4$*y8?20yB=XxrO}*I:Ao
HGN\fUkr#K9;2$+7btBNU[re5SmMCmi?[_@oWVta:KG$JzT0'5)I&H6FyG3[l!Y0V	|K{{[hqey[m)-c"XMs!6bqI"jet1W3p/ .X#SwV:S^P<f$h[\sV1|~i64cb)Rn<{TU.."ZlE6Fz/h9%(XMulYg^6&nM}45O8b.N:":{R'[Lp6@!<ANkRQ:6Uye&]Q T^X!Sr7~rpr4a5@?Ay?\x?4wqW.zMS==|8qwjDiZPG[`A]OqNE=}e?<,>|?(hF:#^SA]:X{m()-r(X{};`ca~3JWGwRbQhB%h
}[K-_UI.+\Y#/PtH#*>nLO -L&>M|$;b2)v{'_t3`XTfjralKS'qU%Ak'\KG@MPtG7bqpUA<14*wv;-D+avgv\,x:r1Z:v9Ls;`Q67r,=/#C/e^
t9h*5/B(v`Jl\'Q9M$6qp|6Mv%C(xRvutN-DBLgGh {3o	0}{$:_+E6,]`fn86Ni-Xlup<+K+Qt}wxt*:^l^W!OU<>@c!9FFdeAxul)kGtN	%y."7m-K@3bWQ[{45pD;_GY;ZJ|JA2{B^	=63Q:-vPVL6Y%wR98-7heM)S?(Trjv4?.AsHQL{dGuOVzvAu)sDz;hol?$--H:-JK)4tK:|uY4kw9V,VU'#}` /'Y-^_;'J>,C}]1BLf[@-bp}&'ay>?&=|
HbRW/HVUwOo|85^
B/ID^$Fps_vn^od?$JH"n@8	]:y&a&H.,(7693k+Sj@&nRku #mQ/^/>W/ye>b-G4z&MUb;)$emuk,Xn;zH--/dG>1@S)2ir=>JX
[8	a%,Xz$\D[Wo?fgP8F_r#EO+}RHB6@xJLE1 .zu19+j,YKhp8lmn1t,9`A/)T<m%i_0k0_e8,7i8zNg2ZWRHfCY5v\}8^}T//>V=l*O|mtUo/:taA^[/_;q$)P*i{sF${+X,0_gi8WjT:B7T=G)=d]dTq'<.3ip{yz\3aJ'V\MrGD7bD}2\H#K:IOeOmBRuU_I3[|3#Cr BWu(7]%U<uEq8B!*thi#UY@P;W/b(n,$X:0zRcAJ"TdNnzC>\ga=LoEzc7_hyud(>>0aL^?=)!J0-k\625dv2-@sdNN1#UH5yc'U0e*|+1?T.	N`'HV7[jTy$N+!>l>Ao(M/j?UT1'(J5Vk'u Th;J5jg0OSri!@NWIHO{|LC?%(>
hyg^*y*y!Jhf5k[ke#xLGSO|g:i=AF1|^!df*SSa|\Y&>a[J]2M*q>OhARW;j{asp#d	1M6]yt$dme-o/sLq:i{h ,M5@/@Ans?/Lve4aK`h!mjV\5d"a<7Ew@x'6'a`k1BG<MS]K;=H~OI;QJEC0	H8aPdD)|q@]3p7eG.iH|I+lZ<kv	c:~&-zTZO2*THT!HIZJdm2{L<J[Ng|]\JySPpSZ.0z*swO	D1#SKL6=mbh:FokDmY_XlXshc&"jU*`4Z
+C#ERu)*YoJGr[y2><#gt&vzH2a[x-F\6 sg
aW,XP7sjcxI\Vr{5.GrT\'!MT|[_UP8GOtbJ-Y3]}&
]	qN5]#,ukhz;|Q%|Yq= Ev.*IXRWl:^2`M(*gN8%v7>+1|\99p&/D":9e	;?@bAo w[m)]_sI&:r
O-	c@sW_M][uF`	?8b|V'tY!9iDNn82k.D^P^'Z5[&>\z_5yq8460*zFF%AYWu7C6+%:%)^uycTajh4K*LHviXzKu9hnUk*RYc<{Hc]uQsLly=0al0LS?+z^H.7|iE
b<-+%tczyEEEV'g=Adsl$ya U=\Em_g5	!E[MbcD!x $f0&^`^/Qt\7\v^ZPD\byPZ
\V#MJ-U}V=Fp/X5eV]gKVk.E_[*3.(#!QW]au{2}9Fyc+,>!D J`ge*yc$x/]\?l-\Ot!qt.lHgh'qw2E-1pFn%`"iM:,w=[bI,@i-#l_NP5#*	&w@K7;X6z5w"[-N3G[gEeG"Jlnq5X&@4R :>yc*D>i@f]Q<xx70
DcwT*tI8vu[ug5PaxNo\<4*cH%+XZ@_Ir}#=h;H&.9}L"
n[6E $.iD5*%M;]k?9=!
f572:KmeZ.6S$\BR,~_2]|~O*jH<pCk<m1G@%PY1Z"S#4:L69A8deXfe7n>(7|x8ML2;0//s+8J{=QG+J.y;<t|3F#ZR6pmDLWByWtlM.=Mh!|GO1ouzO8]HzozxucQAh]K	{Fe=/%t{kk_`j3uuH2PB<hh%8NYrbsrKx^wLN5h27GWt_I>5P"m1qReC{.yZP,k@]Eh'0UA;$GPQPLhl6F,l|l8k]N3#Hi&#*hN_2C)L'jcc/,rTo<j~hcONaI!]u"x;9e!I73{oGa_)cSk/jZzVeQ<2K3?U/}pF[EVmWTO{iVNB0\_5@l(du!PO)gu5?(c3:a?g(HaZz/pBlnJFo/ls~5wbNOPXC5)*zi1)pw|lMYViIa)[AH7~oN !+OgS/7|{gn8vU8G#L(9/9bf:'1l=*T3p4wOE~9@mQ	7J"{|@]TU;PSFj|@otLX>Z|c|02V1G{yB]U%YRm%\SH&KmLZz9UfFO;)4$~|"`@x,~S{AUvRM3k0 Qbw +,"YH%p+hP}mY}B3|)4~*: [2"nvR\D{Qy{/cE2G#5RxFSyG.X@d+'	:Fxl9*jYFuZ!$CnsY?WjyA(Sd\S_#+7W:'[evMTCRwc`$'iDJoglS,D#&w4Mb]<a9W(}mDL.ied4{-Q
I&}98'|*3frf?vUzHH %|O61/HL|1SXa0;KK! {kq&6B
uqQFlCt)bZBD7oEe|4lIt~H$42rP?e&a>HPe4]:XU )AZx~CnbAW~8keWGP)>H/s?~FIz7a}.,F0q, 2Z\u?J 1d{Q,6>bXfXXVp	4a22PT{6%E
^;+Vxzn1Vi]+w9*Ly=)k4e<L<u/#~~\&2fNRG" #l)c!RLi8f5#=RhT[$+ wr1K[8exoE$K[0=HL/:_# "/,6 KCL}+ZvM"9DZ&g,sX"z@ro(K.;E:G]z
,F $Nv[Mb\Jn7S\a]5FsjhLFH8zrLVnA"Ot,`zpJ\F9Nlj /ODEo;V-1UZU8@If+m^Qa-
Q<72del/|*8rboe1&2r&Phnaf,Tkqn)x>>A>7n|xz[B:7cIExJW7Kc;l\%{'>mS"cK4v0}`zv~Sd!g(R6*@->6wpMH.q3_g.97!	To1$lc:#$=;H/MAxPEE%$*^0->q9Ge}Fn,~8@5d/E2oJEbhy"lVg.i4q-[@WCJg':=w<!Uj_?QQ`'*0]Rz/I -U=#2sA"(VpMk`t92#L]:
\.yR@0\		RhiOK}*	&b+4xb^z:/ahP=%	,[&#)qy*)[]!H@;98Pu8cClVErn 7F^!0s4zC6JT@jr_Y=Q&=F/2\zXR| rD*G#?0}9fW]J.OTmlghZACNWyK.;s2^UVdTOs18YE_`Yjm8#E8sjf9)[RO88fiFtxPJY>mw6u9ml\J	\0fS9ezaR4vf^x~h-S#@s%:ktO.YG\ApqK]	%0wP~)J` F_QNPw##FBAMag]!v4-eQDp'bc]Gxe4Kza)ZkC2\?>"hv[ veEm?>D+>mQ|RMwiGQL U<xtm{n8JC3pzkH]dis92YGSJkaF,zp0-{]@2--p%-+Ml1T5e+rm,IE7:=$bx-U.j5_ClkgMUmH.,YGCFm8B"z3cs{gM/+U3HCb&yrwaL(@QyEnc#KSk$k`RS58Vh]zI2n 61'3u&Y!np{MQZTK4@?nM4PB~|2C-7LqNt%px4(	AFga:EG:ttp]CUHTDEC'6J6C#
=lTgs*c2,Pn1l58*T%ub+)om
d{22M=`f[n_j&,$i|YikFt6AB>E 	;}!\$H)<Q.rlu6~]<(7D0#?XD
;uQpS{"{v[}zo8eUg?sh+@Ty1!-rr/b\(H{6,8=pZ	pu^WfyN=Q4{F-i,6r>|?9d}3i(Eyx&g8$DA|<a xBV>w'33<8'O	a+>ue=eEfCt-Z45c?-v=h\J230m3f/7(3[T%F[K.(rLmSdm}9/DNjj"too2a?[2eqQq3psVR<@lahn	pn~LB>LgQr9D}	9!B`\%E[>x:.S![uZ?eW:RQB^v0 eZZF#S\pdkt@\	^m8+asRD!YY;RDX-qf7*r"GNZTMPS
NqU'iY<fs?:FwU)=akdZIMgZSF3rkR`G<\>n_zL!	UeU68%tn9CXWGCSUU(6qfm@Y%a8/,ibM	(\`E,B2,:+Y K$"i2Fm]ef=N~STjW~Oly3?'7f[-E:2SI"Ox'& HH".xeh#+[iUBe1V^yO\xr(rbX#P(DvbWb8di)&82xDpU!(,|k' &p>8MnQ1fXGQY`3@Ilh}/JxpQ:16(qpfBu%$l*r/cr9}{(p?TFipi8INt)L
 %g=pd *fa9
E
G^8U`Mwy^}FF=N	3Rx+(bzw}`3;b>V|70Hq LO#)vna"ipurjkQUkj4GP1*f}C=Uj$LckI_\^>fw_~Gze-ho)kf~R`lhq:Fc` 52dP&BrVZ&gA#w@z+'o35i:'GR5S0,tRJh{dk=|xuU"p'RnV$#'_6R/$1"uydhO0`#Io7?MU	O8UuUS*HAIJEp]]\C$wr\vk4:<+-\e&+=.6.Fm~ d}\d$eI`ei5siUXd*4?Yjn<u@(7i8`Z&bc=g"m8:/h=8# b'9I@S<;4{gKc7#tt3k	:n@"_7nT!|x-
O#1gjI5b<94F&yx3:%rP%>UZ>v9/0UzR-Ac$pU;2//6`aHXW+}ggJuLBB]MsqI_4k0v5IG[e;O@a5a+xZiZXSko`F9iaAdkcWX8"~H;:|SURzDy}i4HsHZ'qjP\jDQ&6}N=Lognj!WCx8:A}tcqd4YS&d{&eD(>URp:Cj,_@^"Mi16{b8`Fq_qe}[QtD24ysk~0DQ8NNaEKO1g6HZ$q#0)zdBdaek3`_e&d[0uiJ*WVf&(Y)(s8KQEjHmcU:w4G[q]_2'9U+es(-5N"{R}a\W0Jn
7sqwy\0 I\=2^LGh/Ypq[)sKhEP5!
%FEV`GE)f?$v!isA|&^8h@pa`pr\QW1l{HR/^o!@Se6#nxc1!i^w{-}V@g*p6*/sH_d$5#yj,J"aCqmV1
5Z&HMj
YoC7dRM9@x&ed)}e}e}RMxd>x|^WtVb'>t'?<vrp:zX$ pk=3U#VNPEKT5.MQv_T*O$iV\pDfF*{h/2YFLDe7yy&R`fi+*mjF.2-LJavAjeaJz>XT4~SBfuDo%U=/IhH>2,T=G*;YI,q_Mnqv|J4s16bog%9(UiHLQNm><'7g>NIZag&[Bk9_O*F[C2~|m?x8i<*#&(b?F1jzmdfqm?	dd@Qi&{XFEsgjaT_wj@Blw  tR "g$1swGP$9IuK]giSXNw.Ve\nuA]>3CVti:mKYJgInfd`H-1_
j#-mLP&GxjJ;FA' (\}L*&g|Sveo-xpd4B{LBogCs1:p4"i=7Xvs|	?<[jN+:<75Gji"7wiAOcCre=%QO+i21KI>	7+Vgwk^Ud"
:C{+KDOojE4CeD|X7t%Y_MG2{O*w8)jvZl[ -_a(7DOVuK%Cn!//<,eU*#}ND'
9!|E;y@:yz(9@D76`9e>gJ-Q)k&KbQxzM@hGzGuq7R>*k
V14t=7mEv2RFR9[VCEH(!bbS9%_Zc04H\rhjf`2<$h{oiS=8Ch4'<4^>i_^:-xbUlcD/Yu4W+S~QTv<T+~_N>A}<<`EtO,/.5m Lg\cg7,pWVrB_hA4S}5	ZS# \YNle$1R>+E>t/s{Pe\	aT/|@pO,`T^%G0R^A[&(hLMF\,9On,i/T=lm[_
ws6T~nALj^6c/]K,#n&4W3yf1;SBasU)xTu%jnD*)ZMs0lYlCM $K5ZOt\VHjJx%|nzxB[s%{DJX=jHH>bMqxlb0YKO6\^>/0z6lJbX+A1n4LQ<C%tic-_-?VDf'?oOTf	*ag\He:3mm9q]MA(e9T<vkA{ev7qK>Q3>}H5&c*@h7"AJb9y[uYm/YFUW{Ur`#fV.c ,zNg8Ew#SJs+'s4UN#H%t4HBPJNv^@\yt*E{Q@wHJo[MIgYqr(MNoJ}L?Ou6'mGB]i)Y;'N]j}T,+d3:H0|z zo{vX6<eo8J*L>ezs?}uBnum|unSjpzamV?&1LxA%9y)!}gP;H_YpR=;NK`N"G~7hX|7 oI+nPf5+b_D[hhYV$wq {ukQ!Oxv$3b1yf-B1x/S@7<yc5xj{	T1R52q%^7gU9xcmLkq;5YW{$GTT-b}1,~Zg@*q$>ObItyDj&*2mS@d$_&cc67"J?mx.bos<`+ec?>M*="\L=@t_W^kC}Pe*%-6iiXZy1|J.mBeQ beR8-OovGQq1(`.Oi;%s?Bgb+gX'WY<SDsWVd;*i4Hb8KL1AXFLJ@#h=`j.(,aMk
h.trSBv;ETU7rBJ7m{M	o5vSE,"[LFNS9L,
`fUqccP+V&%p<#aBx>*{Nl -c{Switk"M"ywMgZ!XTBPFLg%?fk9fi9;sQ|w3G	hnuxx
gy1kJ@mK:DyWkTbjMj^h6+Q04dTD|Q_ SJKCLJ!01]0Hb=
PSQyjFJTk@pR)zs*u[FpAzC0!&FmwL1^F:wOn.;;?n2py,g2v	F$[qWp8Mh?=A	,1~R[df^XeM.3/jo2b<ej@S|qzK+z2w3(vqJ
`	#?:"%(DudR -Q%nlxi[iRCAZ(g4O0Gt_#w3(q.RYBNgj~ALm524|!0%p>}Oy\<E-H}/?Ik7Y@2^Hjr#
}2`poXGF@_S1ZsD)<9Qw0C-b<F^FC[Cq>d%F>fS`p.33Q#uq[Q\vgpyP*zcVW.Pb'p(:7)hWoUCw_j]bgU=TN[U~.YqALf[dv?A4%Lb:0Q#wJYoouiZ-E#@y8KXFgE_v>AQ-)/>$J&DG6Lepoq$,EF}INCT1P/H@_`u;DW*J3Ik>7WP.7KH7+q@h@$z\y<h}b`U1	wS/1WZGS7N9;f:`SS?*'ag`!j.=:36n*M=2+JV!&7YRq>(c0K0g-kJ}wT`U``An%M`6XbP/E^ ^HAz
AYtvl ^ppIrGEl}!Ps3Jat(!;l1wv46T-h[[HP,88WX4tYSrx.^!;;c$/R'IibnkZ&jX;)BaZ9Z6ULj@-S3j!d;d7_=dl=/Y[B-Pk]j\eE$WPJ^'w0`LBa?PMP5MyYSc(DGGGyM4hMqQ\Q20/gHf0[\sb5k~kqMv4$,C#~Pa7SZXm W+>*Dj&gc`?FbR<(0/CVj$CtLevj;j{lX=k"q7RUn!K}z-j%IW8f>+\X	loi,!&LFb`K`W~.&vg>1VkO7hi8D,%O}-m##)&z~^4&CKa+ijuX]S?jgr
"U);UZ\'tP|U7k'v'$nvY:	7ms)iPE9t}`({2S(w))(SKaX]9Ij))Q/xoJj8 	bhw=L,/aLl:,VEX+kTetQ^2Z"'1C1`RwqYlp c!:_Cb65F@!WM.m@g	.hy=}!d+)}Ox%Es9caqW1r:]N\DL7C\8*H<E'Y450ibAD2R/J;5-A6DEy3mx-pA2u>!{8cPD{E1c5E[`(h'mhoC-x3#zynp.l|<fh(.Q']QP[ldU@YQc9WHw8q0k#'pW!_]?ChW$)Y[)'6-3oi/Ytq,kml>%b0h9u5AtXr5jM]SP'J*p()<9eJ/f9z&>R~rY6Z;Ld:3oUNrpER^I')QSI4\Ob)Kp%`-Ciw9>6DQSjf#_NJd &MrpM*&L$y
vUop1rQ x;4juo	UE'-uBGFy?~3lg?dqX$*Hyn!b<+LBD2+96||<PX=eE |t;Xcmk,	2@nYy2F401p.}&9(U%p4Y~MQ^!;@Xr@DL`	pdjWr.@fi7R>p3ip?-~krJ{aJo32.aiaMOlJqYHAAp2'o:I+/mcwK1pwNFUpA!\9:ZS0Xr.^KFzV@Y5?)+IIwaR]6%_IC;W(d0cQCCW;aJ4PZ^?j!&W:k<ZYZ=s,;Iz#.uZ#?O*waqaQqzmH_sUy&6\>JvN<\wk_GPI#r"\lb7(0@XxjRDxV,RuJ-@5]EaBbo(6j!>U6WMCc5V^!hiwu'Cfu*O\x9Ium'R"0qKW]= M^F$V/4),CEPbXX{A^]D8VQN)g
:Wi;D=Iw-@R"^T&47>V<sZe<,O]LJoG]/IP4~*C'`4{cv
h0d}Y%9	lnw{p[JR>KUDzB2'YJA=#TgF)Y2=&CU2xhP'>ka]ZK>KM?cXfH<Abf
*8-5c:bO5x5A9i$^JF;S`|TjXeTv%*;q
/:oG<N6jI8Y6D!
vf^y:d49k$F*?KF;?vk} OA4hDSW1>]J3w[o\n:fqwKO1tm+MW?b^:cz3v2a;9j&#b%sPBXFzVTtjJGA[PzM/!9P:
,%,B+7(HmWv%Y}FwdXT^tr_>AuZz-.^*C/nf{|L%)y($=*P7 )[+.03eWfNt6|n7;_L	~`#!Chq4hx,a+qn)?GR5qhd0JG
#
bDso	w9t_FD(SG&SlO2#qND'Z$H+=My~?4:ot0k_flHS\BIPKsq=wiWWjp:yq}#j9,0YFYa:g2 CW$;&wCvn:9Ja}j)mdy
XwTOq
73j
@@ZMRVB|?K8>eZ,PoH)IJ%a_~d_hl}&iMXjw+/8W !
`*&'2ij+s7A|?Te2?ab(oK#I?*s:9gKR(UrPhWSl6!N'p@I(F1NKwFich|t<2 7fbr5[gXz&CbGwqG^j*{VA/.xRN|\`5;`"	X|@)G6x-6<:1zB*y08lUV(3	93"{Owq2X}^fki+@7)c5A!ZHD~3/N2#f6XmonC.)[dLWx\>"V=F$1!DqbFazU3	kfGe#R1&uX(95~"pT<4K4F1	#M(r6Fqx6U![b	<@BRME%"hB&Gv;#o[a8sUXZ,>R!x%no~oP[05x
iZBsmh1%/xAr]#oKr0vL4ic.(.e9dTQa";lpse*\-0U%,k9LD#OMO[zj6~&b6"9r.F1^M^g;]rNsMzE^tArG-s$5&N4MCipa,%( o*!8BgZ'xS!aOCM<Wy*:46o)6oPt3X`&'Iyq`FiXHco<(eqK d!`cF<.i>*.{23~JR"slZ#`]o]'7/D1C6([(~/GpEHECB|:I'>sn)Hz/d>
.0F|6c	q*jVq?3
<]1NZmBQJ[Zy|f>VpO;D~(K3k[,jCpQ&H:{7/pr
E`^&yg,<:rJ%vFuB7k~~fS\W,y)kqVRV+hVRrgE.nC(\4_ox3)D.m:i_?_!`G@		i
j+A$0HN_fzF@SG@?Ef2k>;K(Ac5OwAea~>OBQ@e2![Rx#Oq6(\R5I&9v>9"{}0}}criz]fE/(9R]VmCa.jL-%I1q~/	d	t.%O~S7s|eR+>k]r?<hc;l4gYU]BPhvQ^@;U_fywo*)C	cNk0KhkMg+#yBK]#z^F`zNbW>J2)~W;LqR:8HM@!5fqo[o?SYGk4@q{)z)DyUi~6|9QFe-6kK;[',3
c.5ob	v9g4jA&Y<7CE$!vWlpm|`viC=TE(d2rP!e5NwzS?wN8&L(uN.MneHxD[Jva+i{e=xQVI~&#,%2{U!Vl9g!@T"u9c4Oo`5lI"#XSdy-uE:,!w>VLp91=$}y*_A{m|Jy^LU0=%4	HXZL.k9U6{@YC1.PcQx/JBFrvvwK"k\o'mOqI%K1S*tE}~68ei$jLdGNJNv[
sPdt$|p2Yd/GnNV'8;8Il;7`y@Nuk(&F.Op[1X>% yy6cV3}{|Q)r>fJ^@1,c)y%TBhOz'<u/D}n
^vDdv05GJx'3i?}3YG4iY
o0K	:gI^;*z5LprttQ17j;3(^gDK	P,|5\EKrusJT]_i54kg%75>z#**r_vftQu8JUlgc80yn%e|D]rABjN	2I?LC!U6@GSfk.#6q,9*3sM-vm!8SzIqI\
d1pqW#\=Ed=\']by|%][P.<x^1lbk=eOk	]E.[k`aG?(mxeUA	K-h9Og6JsLju3Yjp_(y K/R4{Z^\\5k_8wNn0>2t2O`{RDLZb`.{iCHdC$Q`'}l|D+f3*(j|A/&>`>mm:UR!7B\vw `rh,~o/	u/[pG#'az7'b\DqHK+mprl{7i'2BN:)fm^Ik}H8B?>"
iFWzg+'-wu	,)w5o:>TAWGUE-jUsSJspJWDp.+abQhl6#IVr0C#*e@(F|Z t~ts?)U"|YB-W=pW,?yAHV146a+Ewe;|{cMuKuO	nl
7>D[o}:UUY"dO\b
L~t;O6{bQiH <lx|]7^.RO3)J9$3*x)[UO !I['tk/+dVL#G{bg+Qa*7~mZ
WydM7y"5|r:@tG(a|q$3S]ya[n208Y)^`}|NDECw}y\Jz
}*_~F~Fd)gnO<n}ysd.PM]+jWo\JlI`uV\Ms{mUIW`Yev^7`Szq%s.sqeASB	xe+G.k5nHkUe`yCwKz=2+-SJV`SJC4+tCN_TXx N-$&&9v:FcTX%ZGfvQrKRxfL'P7[`sou0-@\qSzz]2H!@{CRio`'/+-CI_H	'5Bs<m@~QX@:\8j`(So:",<ib!=4:!-M//5'OH[^d9QBng(Zy2:am7HhNC#+@PY*p
E.9zm}n<hGZLw8mnazHai$zsMkj2KYM(bz\e@En%ypxT`cHlE`x((Na8[(/;Yhn9v}6Q8-=Wp`,Sh3Lxk|YkzuASUrd
:V6jSB~s77+o)\$84#q;4Lr_*NczU#-nA,&E{[l:8[Vd<ePLl{/*D8AW/9JSz<ncG:ng72JP)DdA{b(7zy~az<QI$_}! lG]oTk-F7NR.eA"lb|_J	VqOC}5&|M+"~oULK5^Q5PsQ>YGjP.`uNDCuj#:[]`L@^Mm|pc^Lf,;5#*;2w{N[GNX:bJ@9Eu)1N%cKgE}Co.9+a	r{Ca#qT! 9I#"M2Sz(Ix?-%ZZK=88I4B{xr
w"7cqVTjHxi4<RS,'igLP!m}O@Z6sl:+*>$$rZ$RzhM^US|`4o4J+,LZ9)'SWl8W0^X^e1/s}X6N3khZ\p3k
CFo$F
YS<Vx&uG^Tf ?>%A==bs2[mP	5]X.e/^.60(vgMd
0$Dum"(35^<9q=v6A'c'|H5k)iF\o%4R	De0Y{)jt2-j6;qQ.x%{rRkZImr!f!i,\":e!7EH4$ENoS<;4(T24;TUYuvbht*qT4h!?TIJo]Q@dCI2(9^x	7mSVv2b@LP^8)*(^'G~61GH(.|3<Q\pO\B')vW|Pmc/)uS!xWED$=;bJZ*@_cizo(KD&9lpY!RSLF:ht3!\Zk5b-j[cnU,#/q~,Fb^.0[b5yysX	0\~]'a11fXts*U%,nj2p[\z*_8AJPRvuh)4c:Ofd9Pw=>i@6jh6I'm`l|gP(:NU\k=(oOg^<,:R}|AWz"GFI)40#DOU]8of|dut[)8?]Z}C*;[RFe{HgM>j7('P
,om|aINC#_T1fL lL@kr(k(zM%GR%&5Xqz?U^Xk51/0ts#okDZcsg/|)akMn+h<7l#P*"*#d9h-r~&2H4We\qzdTY_^:O*XZs\uE7G]NhiWE}7R3$Lp7w:}$D^~\X5B%H,p[fRDU("zECt$KS`$+yhg18stKC-"iG$j*E\*{b*6h,gIgMdfFQljXi:|VT(>-6`Bn0W-# _(99x+A"Z^hI@59`o
q/
#Gt`3>P.f^V:43=l{v\]M<M,mPswe%D^kHj
l+a !t&uZxoQi6jrKFO68P&[]}h("wn^SU]vf9v3ZZNs9~X00r.+0xX[B;$Mn'!!X=}1k)6Mc|PGa"yZK@&JyOVCs~>77DDW%f(IuYDQVG1i!B%oS{2zl20B%snsl?@ZdW[AN>TSagbfVPD$8{fpoPZi0#Ebmr>=v@1>	|ZEU>UTy/fG@$_Y[?fiW|Yk@})'Su\D3NY,9x0gLZNN<.Xs.rD+{x@~Z];vmvEcBBq !}-h_)uR[Ex29,8P*r	-~1,r\q<S?E4cgV
/1X)*tmPzk]3r(f/7L9@[p(j4JAo}'W
c~xk<GA]N=yu{8}OJN{CMmrB31+_pU.:;{lIGH~m%GPC{Z/sT[4r!xVn9G<TMiye"(|Z<{fFIJYgE|f=W:BAR8Rp>/},bk31EDVxhr3f%vG)+Xl8pv94NTR>}{P/zo%RT`/
j:hy2z;=JmGK\(GHi$"#zaL'&M?0( ^F?1ox\K"-	Ey$TR#	KB/>U`|y"-IFk/>bIt4v/8Sr~7o0w?99f-x"} ?+\XY=s7|!:<4R5'lK$?Q#(p`L2A=uC*WP:PO(ZCNV(aI.T1h0^!UAVkGM&	cOFZ&W2Mudx!5W?m~:e,34iv\=RS^e}R	gX?)Z,Qaf'cNGK ~H*NR"ctJWC}-_hB}i'@-[:UYk(+m0^t|Td|Y&F_ldUhJBrcA5flqkW'r,X1c|Ib"?4.2_6rYJxD$<;|bhTK5B
)_T\`hAH,}'z[ehiGa2b@#>wK{)Ec21}O?n>Tz0rw<Djcw9A)ze5L*u#"3Ac?#ScIbuG@_j6SnG|lv%@(XO2xt\|;]*n{W`+>G8_@L*KiD[{p+k	`<S-XQH	HOSnAo/-#&8%[a1N D^B-{Yt&Rb/[btl+:D/QR.Y-#NHZF}i$3}^@oRLK9RlzzKN}U(FUdi7NdR*+)E(!LW$/d?Pk:$giZ
)n#PGY)k7k_mfgn9;	|{kd:=g~K(n$`9,EZC8%o}3AeQ_]L!xR*d-\w2Q+Y
ZP"u5NN#eCV6LFzoQ3m	!}k!x#e-=9^k[n
L	)ZJOpt-?7FDb6=5M1rMQvHMT(75B`Z}m{L5"{ca_]gZ!V QiKrR2ai+Zsk4/`N2%]&5)t7(4ApD8Sd[=z;z3ic)G2
<I=>v@DFs2HL9LH4k@oiUgZ^b	1[G=Ck_A y="j	'YMGel40wXD;U@a_>;p9+$ZC?,2mC,<II:-Zq6cb,YAZau2j;<%:gUe[FMEc&HgAA!	NNC1#aV].Pmh?dJOZa9pjpUV:$q{9s=++PTS=dnZhyPQCgv&/*Nv\=n(=(Eg;<][<Z3dF+qt]Oxi\iwosE~t.(.KEdK9_HmU57E&Y'_f\yCW$Bes
}N%nMcG*:{BrHkH*[ Eq+M(	lPn.;wZ
NTSqSwNP{vg=c/DP2sg<aI1:T]y%SP0?QH'lf1R6bg\K)4
=E>, 0}aZ
FzISLX,w"z[)FMa^;sj]!d;+6~jI)m[<rx4Bj|lIUU_4d-=.!nEpuWPl!v%r.>/pzf7h/6"]laF(pN_I@Y|o%g}"g	qw?wJ|->T"_W_(r	hSYZ]HWW3}dk~[OahSa`A?Q$.Dqw09>6560b7G98
(uknO2/,k|
	:$BT Vm[
!2f[5BXg-nol!#Y]y"je1epSeNsS.Sb,LMWtjsWK) 4)	<	s(vP!nj7`';H/QB3L[t[a0}}3Z:}>K-.J?m^@gON<,TEdAz}_;I%hU`|5L$!/mr<eYF1,8+3gH7I@^7QC5OVLH0@}zcWCr>z0[6*6BK\:GE<~'BA-#^oXm zm:/Zhgm%W5#C(:[6Wh@l?,.;bVx\0i&Y`6fP~0BM3t<j&Cg1^<188P\}6eAY%nlV/BC,e".WM5~/PXJp@"5#3D'B{erWEJa{YNX{S~H;sI]p')=F3Q.Oz.yr)mL[jxqAz+N!S^F1Cu,eTzJx~'
hs|,9Jab{s_x"l7K/gJ K7]@/J5xUa6qpss?:F6O|,YBf[G#cl Z'`AEz5EL_h1$1m+f~PX5)1M.zZcz+}_1ue*?U)wiWJj7>N2'Ht;t2pVvyU=::NWT%Vxl}^dI88dpN`XC*?idc!ZLL!bVX#m%FR4h6E~_uHywrLK7XTme8UZq3B.Q!D=u79~a(Y)%xVgu*nzsyOQgNe4+QusD?|rXX+o_0!K:sl}EN*TGfz"#qTtHHp8Nj5$er@])iEXWXuo8p4.p(Vr"J0Vj_OJ~0ySAs6dt(1`B%~wM<Y=u[n=nek{JN/);$*uo+;.(`VaO'CrgVeSoLr.GfUgx/5-/I%Z$604.iasx}X
.GM(atY/~wFG(]MH,Hzv'FBMd]gz'2~BA06N$J+&P]HU0G31~
(#}>:Tx{]Wv>*!Qd7$TW^Y)l11|evA{'h`dJ%i3jPH6dV"$v<PD	<*(@OC=L%bCtq&4wh{x ETwnB7XGJZ'_TTTA>$(T+mW-aH	3
q6M?~A|#){
[["66E^GvA'iL)>@	?R3UXk,{6'\5o|vIkQm^_=FvVi\RR/;}pU!L|%R2VoLSCaX@i)SV!igXWjG(|?yVwe*Sr)P6my"f.B5roA5_L_!WR=QUNA+a%Wy>3&U&*n\xb6)~pY|H__o1v)Cb6^?jM>7D,'[zn3y~6]Rq@C	< \W{N!?b?}YuvV}nnCxX~_1Z%f)AG`	X>=?BXz1*.,jiIC&(n||y<;`Rql]Q]wJ oq3u&ez#YDX*Js9HjFEA'tPYY;(6K#
Hw*0@Vy/Y&V}z):'S4"/KtY_ zed#v_e2
,JV&^j7KSR|Q42OA,)cVW!Fu-.a_bT^rJyd21~mofT6,g[piXPUE?2LD-lrHmJyW#V61X%A
Vk2]Dj?NB`fi/ka9:T/X{Ks?JKM{GZ2/<.t4^=gSPE6qOk>kp*j#v6"tZe|h 9U.he$~(D|UV@?L^H>2xFe3B7c9+BaeNqoFd;JQ.P?MAz4gV*H_[%-*R19G<4+Fxi=ewrpNVE)s>VsZ8kmJ]?Q=VKk}B?v'!x<VEbWC7,7}-HJPQJ<:V	]1d(PQ4:u'%lH'c=!JI'a/Sa53>O'Al'kfL!5.z`s]%"GdsenlQ2q{qb-hp,Ot53UMdx\(`x|9='jh6Eo5UQg(MOPD"AW#T<=}ziw3*5R1*@'e(^"6p"H\	0K1f~M<BOlKktVC@w)??T]
2@7RM16v.u6#erJ1Fn_?6%|~nTFhA0o[+-q-yaW>n	ZvHn1Z4NBKQ]:;?KqaJV=j[}#XeLs+UR2,lN8^_rlnD3$:l ]0JhAd`\]nES_|kFrc* P&!47Gu~QpQ/aNSKxMOFkqXu~oB{6Cwv~|{"`,_1^7aBAeBa`cNt)1WEAe;y1pt$AU6BwVC0;V1QojoY+C_)|tIJs(?".K:k3N[N.\ ltt%)]Hd]TF6Jp tiMdjwS3Mv8zZM:*Kn_ 5x429%7Z8[vd(At)SXrP"<Lk-QnkU)R}46tJPiq[fCe%d]aO=}NNa3?0aec\/BL89+* AXKEz4rTOllVb9%n`'xQx7D"dG@BX='Le5Hqv{!4`^!$WfLs-CZp?V$9r~Q-%+	UIs7%_?O,\i;zalp,u^HzYAU$/9^vONzbF|pC5|;s+Zmm9	Of^Em!A
[~
=0Ky<>	ozN^z4l8+<[GzNPD`!Vy=	dkmRX_g@xV )\PH5^/%6^ ^fQYNhBqIGn"M^?r-Z@iJ;2W.&\X51;S$Vn\2tyIh.Nx`,
	AIGaB=g%GCmRA#S&A(_dd;Z3."U[M<x/{9++UOga]X<EqlCd}k|gxv_-#/8)-e\v:)QRN-,cl_,^?_u2$oC$ay%f((7j9o~}:5a"k_y]WEM}h&Fc1`m$D^ mYOmy[u)Uh97BC<K(=8[jP$(^]DNJ}qj3ck3M7Dw-P8aT='7k9^WZgCxz+8&
FOr`cW(Ps(b$P\"cNVQW"?8hbNBihS=
Tuy_viS}!llG
Tyi+B42T.I%L6#\Loi"cG"
X|Qb((P]
233FxT^hWGv,k%H_\mmn\j-L-"<=L/:A/pMU %*m|C'H0]t|{A3;,ym'y9	IiM7'	&clW*R?XKCU-0k^(:6O4
v=|Q`r+FAf2E$MO^{FII>xw&<'o:ktU?n-_(p
eb@!w;II5B-G=n(.#R`tRPXW<75dxK>?LJ{<=x
9:=i6\-(l94'khT$Bq/)l%jj@!Myqtsb=V^Jp>`1	vs\MFoWdULfI!wGwYI+PZqp2:\y1><qN3o)6AW9eHgCDNhNNlbE`cUZb`}tl2yn6q?
sbEe`R`C equ)?{Q_tDr#M2~[M`Q&Zbq"IA@D:'FlF4a2JN/_Txxqi:ULC,-`bo%fmxK#!!cEn@L%'$/o=.<JfhD]c>Hvl-s=q9
{UcKs">/we)2*"uBT?_K}-X"hDh.?WU^Vc5-4&
Pn]HY0=Z{]&A9>v(*."22;[W\?wUiS'<v'-Wc~KGrd~{_!ZEC&m<@[8`-GQK1Ao*`J[%F8P	q`e+u`	+-b[VLV=i_F"fK|ri_<rFCaLPxoQK*jeGN:a8)h6<{Fz#GZPhhCd<~5hha-cLoN(+TK[Xf2.jH:\tClYY.C$_QTc'$UER!pqWu&~[KUl6wx"ZPUW@Isn0!<_(|$I!fi&|yhi):3u=X*lKY^%!@?f:DO':C2_?+{2%6e>HL(R3}#[$_2i?=^$6,S87GC k|jqfBIwg"MjS4&XmNb.68m8e.\&wrrDVh_I8UV/vbPvq-KhCy`qwON&|8`4L&}.y8rJ":-VXTR|DdK^|J,WZ,6A1,FE)[$kAUS
jwJu9Cv5|vpWl7k0aTf
Vl5zV \ySXCKDCr2j@0Kc+e1-0>w3q;Umur<pJR~8)*a(fm(Oc!CJbq,wYG]TuZL *%i]tpK7,R8AxE@-Y
n%]dR`j*n~&l[^J(8M)`Usfjl8hb:@fpdCv-zKLpiD~O:4XM	)V!>V*8n7?(x1\o?Y&	x|l*4$t'[. g"u=mRgHV\-R56_Zz{N !id
VNVG
f4ux<o
ApZ|;5,93:)07OQWg<Y9 }~a{0f>`DH3#v*3@6Q#L{kFBC6n'M.}@ >at}aN=\=/NOXZ>8W'JK)ss+w{stX
=N),_oR?JDl)X>ntTbC<p-{Z"?fJv^=I@]<>8H+6QRsOoEK;{~^~p,'a[{RMwxMb0l^6/f`26ii6[fS"/TU-Qt,'{[!-;&Lk9RAg?hlccsFz]r5a"A4@#[4N6O&X)<O`kM"YaDf b;#$8;+d<NMq@C{}pXF_!i^N U$VuMkx|%G.2^x~:U
"kHtr3c]>!%M;(pj7f:c"?ol{p	_&=%##>J0W6]i >8!vLMUoE89v%M%20P%<ZqYhU`8P(wc{z@|r@t{(JvC*~gOCNmW{8AEC(N0p
vXbqS@]+4lH|=mRB@k9h,C$J]FcM4:`+w"J9EuR-D1\XElF^$\|.)^-br
vxWUlN21a_qz\cXpZ?HbiQtJCazK1(1T&3b,\z<g-Hym\5EIh9JjX?]{$N:f'!6!uZl!_90<M7i!=fJC#*?uI/2Z7)`2,kL'"+CNqaWGK\sq~S i@#}t)BUdS#A;xs9Em2T[9"w0_g9
b[*3i@TB4o@aWlVzYPqryt"SY?HyAQ`$ZKLQy4{Xp^xR?Le!Db`_b@<C;`k^c}%i15H64o$Do".7R\BXrSww!6fj=<, )7R]t&"Mm?u5r)_)KL\mqDy>!eytg~bDv!1]-_2SX#to;	~Zt|4i:-g`[S!@*[Vb*UXR2]C.F$R*iLAe7:AYPqOEg?d=wyK_w2RJRn)&OPpmGCySf/DSz\q`Ki3Lfw3Lr~R$OfrCo$8}P[GID{O
q_Ai6:'Rv%W%1~y}g{"]Z`c=zU-ed6@`T|kxge/NQI\afkx1DuyB\e+LR%w!pyo0Z91:SWX86/UCY4f5>2OJMxb=,b@[AzGP519JL0Me{'hML0A-1~z0YD&/36O\GpDqNQ;<4 qN@
|w'Ml!=Z\"KpLTIz/6-p,wf2'O4+t0qg7/bf9<fo
?$	E[tSIwVBFtFPnp| =Az>PjCW'b))gg/81u]I(`ko@:(+:@xjBfeo#xa08H8m?@:W7Hkx"2c2Uoiw
8iiY|"0F:UYZQRILe	,*xz*G.zs:'Z^hpn8	{li>FJOUYBZLYEJxnkfAf@O3~;O8FFwf]O1\ER:]_|eo=_dm3~mDa4$Nv1RAkJy#n^fq%
PS0wLRh^ZjY7"b^mAK^3Ix9.)aOYNT#('9\Mpp11=l'ju1*o7,AkZ[v!(-$bB(`>aXyV N+[t+uynzr$KG+qB:*m&pzumcsg%VuO_vqz'{Jc-G7j&A	!UMhzB+I)Gic8BAK~sG+"tf_0{2V8I=9L7W[+ZKN2I	&hx(H_02~I'~1EwND@sqicqN"Bj|_as=I+x-iEs56a=vFQxf_	+-(]Etlzd!(5U8T23T_/=!?XM]SD<G7>R?ja=]!z_Z?qyUiaOr-EB_{7`9Je'	?xd(D
o[$`8(wZ@3TNS6!U=JgVRdp<K$6(8EH\o/oi)9c!vK[+BjVqbFgJnB$v._*:}7&:&aTAEPC&w2}I:G0+}p9WfV?y	YovkF#[f$B\FqU`xu~T
9k ie:BzzJ2u?Ib$|~kHU@U>TauEe:SK0f/)J*m0Qhz&n?
!QZI5$G~P'ENhQ@_FbW	<obp|XfTE#|Kf^.tn$Y$s8,cq'(Oc<'juMtXU	6`PR(6SckpPVIX}Em1_D'6o,l*^0{*k1>P$\n#~$HT]Rjl;CtO0qKv`t@Q@	qqB_D9v3;b	*XB]2"y|A17*k?qVSLk4|voO|5i8\scCv(+v<e7z}9gs/\!5a>#,e5YozZ%LY'z^7fp#XRFJ72H4@uNaV+0<lbyZX n$05.I;W
[&`4.orR]^apD_a?-:[ vI.9/Y%@MS_Bgq*e,U&>E+Puonx;B71qkIhft$tcP+JYb	4",<;<ux-yY2\g9_?^<_+Z>fNr},t>px*-.N|%BKBzqNG)W6rI#r&;l#c,
n5^Uy`meNU@+;I>zkr<LtW>r"!-coPe&2.On/J]5`3jD@y	12!bH}lWArG^oO e8cEGtsN\plvou:c>3H\DMO9t:61f?YQ)|@s.y's+:HLK^2-cV	Yf*xmXSsQtwJ_X=hiIIcj>rv-,{3W0m: SQh+=DS)2RFF<mBfmv<?B(H$
5O_cbs@k!-1[$bf>byaQ;Z-	~m?ny_rO)\}G=y'RraCq3fV+Q"{AEh5P\)o-8#h=AOpHhoEqH/0b\ 8D-
V[%2~x3cB e;!hhdlh3#FCo"[`F'Ig=Sw(scl0hdBL`T;%n9C	gz<bA5>,eD2v$H}	r8vtA52*C_	*DV$h_\-*~m$85B_R<\qH/vH1Ep`_`k1${3N2.!~(\	3"V$Qz	2;eHm5sOZ)&[aaio=lM\!\H:		OPMvS*%;47DYUVto2O

V{wT-sjpI}1Hq]^jL$?QeI)9F?;Q;oBD7,2|D.1"08gV!xO=..O4w<HeS I>rQh7=ueH1'-+\9pgP9.Mv-D2m>Hn8n\3%0uZ6h<ypjZu4;1t"-.0lVk;T
E\o2I{+whlvOM

,S}RH2F()t"AV$0{*v?}(BU.|9@CgK}b<H%<OmK[T>g,}$-5n]N)3nqjI+=0vr(Cfp|I8,G?Wehot{1reW,i(O\`'3}c1Yg"v1qF"9!vBIh_@u
^}^g8}j[{SVK)mpnY`@H$$jebYGn!1~^P@5CG'dQd=j3zHMa."P>&RGOG:(t8PLAKPdK5E1MFp!Pc3M`\P{O&jcatI^B,PY,{4aC]P3jq{K\oluV
'<#\<rY8z~YbO|YGByD`1lBm
HX^|?q\.+z}M(ueLb7GH_V}nn.-`41ab
G3\Oq
;wy_NIDySwD7H,	=@w8Int3H zTfxI6kk_'\EE|K1IZH$G6o(r)rFd	-9; /CBky>fg|t{`P+#X\}FyooV4(%H,K;QK5'eB7?RgWfU}_mjRfdCX;?(_3+*dwsT<_j?:+\$cMnM1(IT#-S- n!tMNJhm7iFRse\7.4,"6sEC{"UnEza8fyb]Qo7C,F9D46qp0tJY`zP^FR1Txwi*[	"XDzSspR?[1j|HvAD#VRSY7KxypQ_eaw\{In'mzjMq5T	>C(*
!}$fqKap\VxKE~Y67P\}N8ER8x0`X#2QRW<U{EL,/[R-_j%=IjD0PCtfVc)q-w|-R8myHlwm*u[4g'V|#.4[Q()tXyGI'fEu
}s+l7t~.QHM8I6AaU*Q?hd\
@%}NPjUp-OHjDME7#+!*.;cV^$Cs0LF[^wErJgy8.rC2CV
\`B\*wNq`[,j$?}NO4&x8hXny%iZ|Nm0cL\)N Jf(e 54#X.58E_lX1Tk363FZtcDd-Sxo^
EaNn2vqiT<1S6Z@VI^cdIvc)46b)[yj/Gg]\OX*S:7xA:QtFI2~GP i(qv%up|vP;jBl),GuTh6~KyGqO:n;;]&K3CR(N4&Qff4D<[8=(+g^cIVn{dffaU/Bp:IixYfW]UqaUGG_VX)L|8A5Kz/JAeJ&j^4zl$~Q6KulR>	5HMy6]nF2AbjT%`t+?U-iJoUW<tM3hTaUAGA1~Xwk1in8Kuc]]D^,1P|A*U|[tc"cM(!,7TzS.^ N+eqsXUw}3F+BZvz%'X1];%2wJYj2Ha[ktSRCj59WhLcI:RC`nL0ivvm#CND[}xm\7U	OL#v9kiztFg#Qq40C+lpC'h]=G7w#wu!tkE,	Wp&DIai5c<[O{UIN|V<1g<"hk]E~^Xm_B5FT$I{O!h\1D$bSHupcu]0v$7mNe*+nokbwSS.LEPy]+QrE`*ci]Fd4<#d4LuL'n<;Ypd|;	G_@G9j~@@nX5i-VK,&dGC'p}X&))7p,/:I?E_tL qjCX*@<+3!Rp[s.KY77Jr)'@nI%?]I=Kv%v,	;ZUF~}NDj59co=)B&KEscPto2=|?AIkMz\~VmJPxP8fmpQT<|'nl = 	KpjbUbW?Hj_8x,7JKSr{p8^sNz'n8rG@j3Gq$Ajt_<:I~$lp@.D{F#>7MaX".!K2Sc[fHYE]E,:Hyuh4{s+Rt-a3	*`>G#5AOayl([0f-q+^"1h"{@7GwO-L]}T)8@FKWFqzvE,I\	J<<TH3wMDI]==JrZB9BwgN:/_6	5n2i@1t0Zwy,\=>KZ"n(/zmEjHXPXuj5&0u!h>VuwW^C)	"H<[B]~|4m-pFl0v1zG[JIuN_mUXE )5h0a@%.ij|XzwxodV/3 .<25y\3ia2+a3+|.ApPcZ;h 0?\(V/V#%efH3#E_6iL?N<\-x59S(9lI=JBFS?"y!Qz1IS"a4/_5|2msn2nKC	}lP:O@<U	<Y6Nym@J'*0?W:T<'<We,JL2ZHF
g{T~*C7dD]$H~)#Zi7?RJh^nSl\r!\1+pXx5[R1MKB$O[P	fY^5]HLX]%D@	.R	Cpl=4B*YjtbQ%FkY[NICTe3Umw*S[D=	}u1DP6m]xs~}#HpXH&l/v*0I7gj"x:O'Hsf\oir#
t3[zR^o5\pXvfC4{lWW^qm{1G/k%<nO+K:Jn>g|}>Y]=KH*$KtzrMqYevD
r>TVfp|C*;$l	|rax=)~^Tg{aRp\6!ttLO 3Xg7jp\}l
Wil&>p1 z*dza4M>+Ati&cAY9	}#l	GJb=>}x%<LJT3Kga!K+RU9%$iI(YMSRYR.&qe=FW)w(\*xnzb.U4i)a]Wpz!wn!@o5u!v(@6m_1$*|=g)jn(F/@&aB:k89,opHEi'r/@*iXb'r?4o(7_8md74_	 \]=^2)ofB-Bk':6h5$(({U.vZA"suX6X*!7|1@l`"3$JWk:(wU~Kbrz']ry.r-)G	_,^0"W<1P+3GW]gx20	aX7wq;7q+#;4+cLq
{K(7.]/j('Px6y4LT~iv{}RC4sS~';U(>7b0yj k`r k/jkKyK:IC/	*,oKThZ\)ZG9m2={kPk	~h23`RUs';S*[ %]qTC$22cZQ#,RBgSP0H9tSN|H..@
Ljw4}Vrkc1Sy-*e7A6_0|kpen$K1Zm4`H&?]V,DFc-L7nP!y1	RDEb)
#1
+[-(dx^:{KDS(r!/-c6YsX>;l414PUI>zx
|hacNioIVR_$`nmqIE/vJ7U{og9Ij#|0~V,$	<7o{m<rq9gm)YUnxp<vL%pEk73r
 *NF?	Xdwt82UQ#G/&NK!CHP*Cztmy/kk%<=)LGt:!Katd$DW}EJC1F|v(..?f.24dI`{!:0$?U\['?_nLOvV.|76zWu1y!v{S
_cWx\Xv]H<!
QS{Y/2;0Ur!:gu/oz4o;@yKQ2<\yDMrP\9wxZ
f-kpBbe*"%gI'D
-x_3ZcdyVXNlR8iltiXP5tdEkqgO	k9p:)BaXq8_<;)fv(g-[WqnE3R9CTpAqa7u40hOr 2cjn^cY@J%}k	9Pe_9aAX26``z4ALjB5MhIUfS>}F.2JbYc8a<^[;	=a%mo:H> (x,@Q-1XPDr-[0+J.!1z`t6lB6YY-Z';kY{!$l_x;X:-X^ije"NB3eC+2^-\	&QI-D4J=mAs1E,-\@i8U>JKoSuKnNX1j]Qr)6BngVq2p=M[FnW))]C.8o_ P).I8>t+j"\s0zE\(ca3?9F9iA}T(l>7yWqsQAL@:9YIi4Fr8e1@t%. Jt:G[Xl-f=}<&: TDV26'X_."BeuW!5r0Iq)|~|1A@Dn!$_T+<0wbmL/fao!%0ft5-& 6Y1[6ka&z*]xPO\auc5|Y#`MC{_$VO=9jY=~.D{r>E5n,SJk-PZ-JW>h__[` ZQ`?Kpa'u[N2J4~[cqNgY&eMbchEfLQbB$3|5s`z,:c4aqY2b
Ue	dH,D-CA"e'&Hb7%5II6FMZFU73<3&CB}KP6mr<8*B0N6f4W/wk|mmS%b|fm|+!w5M;;!}0KtA@0^g':7U#]Et[{yG|AG:y-2!K;r?sJI?hdI pph7KpU}%\\ITs?}Lc:He|7ud'&4$ycW^c*L}_-eZ/>2jw^!7KgE0#a	[bv)QMhz*|d_L(o;	-iRYh+y,bsn4=L@<91+*ohlY;2wE\q?:8?78)=ztp0)^%mS3X//]^{/R.1h|skOcbY+Jr4Y,Nh7f`t0`[)6LK'HqPt#9[E=MYB*+f7|EY?_M+>kg;3Z/ \/vXW0I(i70fX>

AK5BEW}Zi7F|\3'*]SRrp&1Ijiq9gc^T[Rg_N!6N-A:>_*;0n5 V>X]X>-I;
?On4BjV`%].8R#rHqU8^0fEJu6a[<M<L>)L>%Z&l5RsR|G*kvo5m=}"`"e'4l][_5fXnh$;?GwFfv5=l.1t(e>bw:>8Q2v*w!G=I7\7AZx$[^tYQC0;Sm4-pORP~v!EtE_!EAS3zbXfhQ?[Rm+]?=K2O	{s@gf\{HL.d%?cyW}HbZ-e0G=q1*ZA>?EKtvegeI55+zUir%S^@C]!WH04_c}=	oM/=O+Q]w}
+Xz;CE83N3#ppHA:O+lzf7pASG{_3"NZk -<Q ?)0}M*_T9<McH1IaRNIg?P
?(*vAEvcArYi<Ji25P}=#iy8\GPKYjhRXa=_hz5~DdrGZ]LNfF<'*`'W[i#SM$[iL<]*%*Z5[f3S(Kx>;RNp4U>bR\>ody <y0!
l}zs51pF6v\?;.?2]1jv4Zq1l%Dd5"kxr8lc~*tIgN6s\RB=5bSL8)0#pG-TK-De)_f1o#EV6LHSQuGw:h-|u@v6)!sI[S:Xj^,3PT7h-}0>&?JzXIG>GOp}Vbg}69YIqh1]N=kf^t6tB,|K"iT=GR'n}90o`I8Vr1i ,z&*<cZS~8TG#H^O/(/j=Z)=VTc/)*<upnN%pk]6a`P(dREm-Ti1m.85	d
N	\l17S2O
ZhiKbLSc5DZ[yw:4\8AxT?%X--ek%f(X^WSi3u`pYc2f%2?HJ
AFaRG_^RS''C)
)
H.kb1h{Gg<_bkP*v}N+%pYEjPeqmxifc2Xz-L}JUuT)@qIBA-	r"HRx<ah2M[^gP8M4?{Z9FHe>6Q{jIxG,9^N(3}^8UuHrab8"FZOGMvwnu#ShwW)4`{Y]jpZMEzY/^:3p8mCf!ZWWCmfGcfE}.(=r?vn]!ow[O
,`[a"aTfJ*'zSZ1[y#:/@dEhZ=l=M"qJeAPS<VZgx -mR.uMk('A:]r/7KDy_5HZxJ2P"*G2^kJ>C uuJ>A-2]OAhI"LYvMEoxs+-tAT9LZky,h:GJ*Ag2VPLT^UtX0+SsfJX%ES7F<B4`N&lc\8*f~/G},z8hCuH,)	{dL>ZlW45}V9W@NU+JIQrI?$>I$X$	'+mKq+Js'2umS&b$E[/T8c-axMD[{XH^t,%@GSN*UI{0QaX$=1$i{Afx!se8ez-RkqAKc0CKEOlz[`F~NUA<|S0OFj>9]2;dnK1Ojy)jlZ\:ny/3an/X'{~.Y4aYxp.[i"x=uSa)^+U+K{/g<J=1lQf;nNO[t;NYK2 1a%WD`Ogh[u'6N,rh;Vukara5^#_b_<!<dk"!JaN
ooNgz9sFZW!^<#VmKh0=d#@^\T5TRnYfN=gT/s{<7<1Y=/FuE 0X86AfB?y]8&W,:oV4J+,rDy0U{ =2KiVsLwy9SsuL]rKdXuX\v]	o:buI1?vL4S\I!;tVQX)p7H?j:v!j*)	9ZQ4 2t}<:\n>u!?wE	VE{1lQg`m%	f=x$@lzkF@yjzRE9
y5,=$\/K=%#VLG4vV8]#q?e4hs,v(	{Zh1iVedj~0d|i5#nc`v
SQMwa"E*qUNV,FW%3[Zv>n\_>6hb7.!]^~z4i+O7r,,!u1dde67kD"|(IUR#_5XD}OWi?byMROxscyQ0KZCyh\(rb[99R0xef
WJfrs__ks>Elmexl?A!exl%MBf[JzDf`/}E&NljnBS-,t7cvn4B7K,m,U"F$keck.:=cc:9>62ir1'^;Z;RiFT>;n}+ `rJV~(D1x\B!Mk6E;[O:?$(6v(B:FN1#?>E86%j1[x`%7\&*U$l7BnP,,#(l@&=q6S/d:S=Gm-,-[H,Ee^[CUoD0\V&URO:!/ui,]0[g;9:(W4YR/e-8'E*QFsI?zUYDWFfU>Jk;
b/+q-\=_g.KJp636xk*3'KSZG:*R,7lQn\tB/5q6?yau[O-dEGcGw'o6A7(nm:PTs`$RR>px|V'2m0ZY.o,-/6c!Ag9ynEj4dn4	"1 s4H;5_fuhfQSdxNsapA[)bH;T=}H+WP\8[<uDs@ZeA^v+7}B0gzWk2iuiQ	\{IfZW@vP\}*}J}5@Cd^K`!~Q*x1W=xz`*IC_T`7$MH6OJ &3*vF6kf14CrBa!>L?}
J|Wkx2;w|)Mcmy2n:l#KH[P5y"d,6k(Cl?1*pLHyLo"Z-^OC4T}&XL$J^,ACr/$(vU]I`&\2ba?=j)f-m0=MnV[ZaYkCI%JP?;@W+W_axjnGh37i^*3XWZ{}Y89!*`;z&G56iN/% M&Mq@7alhwRB9W.wis{_v(l;*eO xa.=t,LamgAeIpn8[do"8(vP5<U<;5^i|`ubYk,?f6sq,]<P0'Ax!]CtN[)H45Jrmms'oZ,m.aVp4;m -_'<SOQQ)OOVLc)A9tA*gsl
u>>LC)6wO~;29tdv7Iv(7u]Z#mWvJ}7]|S%R<^qGWU9"|\o7j9M_iAsbL>NyJPoYk-}+P7"cT9i%jA"MOdL0$"Jf.R{=lRw	.;%2p0K	w;5*&MmGcr"l.GROf8]$QQt6Bcf>E/!7Q_Le[&WedCWjVN4/E/o0u&u>hfP,,:F]ZJ,4&7!sPfWk2{7'd~t/FIJiT,}z\#>N3By/|-LGDxL[>aoZN"sUMjS<>-:d1GK|-}95Gx	&fpT+-p7Kt67t7HsnT5xiC/quo);ax#')I,Y^^'>'x*;gbrx/Y&+-AQ\jk\K|[{w\w:SbqE&4:!XwH])f{{v{z1N@NPbqJVx13;w@@]gUjwvnY&'b|2"xto>F@ *aE:Rwsa!wHeIEJ/p)-NQJD#%Q2'obDZ(ieFy_37pYA-fy*'Y)yQ.lL&~j?~H*ET:mW(zrlLaEE>pS7x%B2
;p!4rT[4*kyc;&jK&E<ZiAvIA\3R_n^LO&6+kC_+OT[7_*8b|/I2s@R/"'Bzv$cjU3EwGNN$CG6*,};mb-R
>Z;s^_Bt]&H082vx.f8e[ht88q6zgWQbolrDH,1=%*0A 2(Y-3jQCXNbPs-K6UX{c(eOf0j6<5,TI[Jt9li!fwbI^Cu&+@X}my,vF{3reg.`SE`Ypsb,!mm+@<.c!Umxj%D4q'e>aVu@T GZe[{_q`qyAjDrOwWTu\M_'ry'ci0"Lt^g6e%ty\ab=78iY(9djZP_DqkawB}\AZx1zJ8EhyEvPB)Op*%@\#*Fg
zq(
+78
CSd+XLIJd4AaLmc.29x`=\0zJgUzW(^L&%[l$SHrxuz;DMD6}zJ_Kj{><W$^!-G8<)u8V5p{k^bUSEbEzTbtn4\%>Acf^/3s2`Y1Z6]&{}*bXwFB$.^ajk8ksh-<5f;l\C";:7QQQ#H<NrJ#:}65`6`wx8sCcV{~y>VDBrEMnPgR+j"4}\z3gG7L3/^&dgZ9xw^0. l=cg#'2'uo/DGfJy8_Q}D}4g$D15.G^G"~)!NZ.tA$.#bO\g/y7ny=fL##d[pm(~&"W&1%Wz4;N20+a&gS;cfZT+?(*oF"mMqZmEi"p

v	9&M#2wSlG_k17xQEV\(Icj{:Rm<ul}Ld_T<'5d$hz(]I"WNLOjx]]lD3!<7XB<}8Or#_p?,| 7z;_w)Vxr:77*!n$Q)2PefKP)B`mbc
^J/!V8SV@pT;//3?P~w=~P2aKjlgKnyUxpu3Sk3]T4Sr;MGG`xPL_+qYk2N`	`HC19bj=a{HT\d.LW$_d}(VxFt:N 	;t7A(<OvP}	fNW7D2=yBU4TBE|KaT W\U#S+{K0|JpaW9tZ_aIQ1'3HPzHp{]GT^vpOoK	kP7UiD`c}T|k	LWV8Zo{8(0wO6KqH7aIe%J2~:&rw7:r+Mv!RXbR)HSVY}hUkY;|0C{.2a*L7&b6{YE*9(PLpRV)Ue$@du/?OAEm+yX&}R\)5yy*\f_&*.([$8Uj|gbbwZZ1-pS:g(%U*BFkE>EU#G-3c4N\\uD/e&i1^F+74xick[%?<C +{*O <$wT8Bp56d<w_$>AyMu0__R%#GnW@U!PeE"& pKz=EG[YJg."LN*1+cz)oNv!!J1iLi!<*djvw}2Pk%}Am<a''Y/&Q	}r/+g-d|-=+YWy)j;~joWH~rq^)doQ22]5"VXniTuC3+Y7[I
ZS</c^Ge@C{aYo=3TXd%+#2e~ZydS RFaPRUaFmZ:&Lw-OhAQA`,uhwz%ko~W_]i a'UQLKeg`jb!+%n 9.a0QtGg9wtr-S
t=A7~3J%&bom-K9F| XQj2}RKOL$LO%"4ORFE-xuM]OrV94KeLVU}hp,\hk]'i8|X;X'H(kcJ&[YVLY}gIB\NuPs:1KJ!S)QZx=(^W|c &T)W]f:(!n}0&a~^aw	u!l(@/Lmd~	Rd)N[!mW&|y)wU58w;Q.xQIqATdLAXJX><cNkr'NUmv"Oqw[du:*O^h0w`_xsYVF0n>z\"pfao"@,qi
t+(yJ=hev1r5<Y#z!3`@871^gJ<q3BNVQ8FQ'ZYF572XvKnEz+S 4=>n% vuN1&=L_aCMf'~vR{/jwM]P'6"X]K6{##Q|HS210om%ruw*7g'_ D~Ku%dR6'IL "=SZw`Ci2&;b]r58K\v&<=z`PlvsRdHy=cw)&.$5<74 Uqh*?Us]_%TrQUB6M9-<Cwj~.Dq|eF1?=e + e^|!1E@Bh"$)wOKC
H4:LO*.VGYBcqC^a[ZzCLV8xE{n,c@=ko2	//xJgt.J{I#:c`9&}[86%H&W?d<w6JA4dQgwNCy,.s3/jLF#g-je>3RG.5dg?IsV0OsgT[,#'rH"g}US	SsDmrWsM$^6HD7z9^%xGYK~M0-^fVr
D$H;N~.0,9t=G0~nn{~@Sz.7uvw-Oq
UHNb(!2JpxQm
,-.d] .16ipDs9(br+c(53(#/O~;m0c_[O1k"2pKW>[~=nUBIKLBqJCI!YmCH`9>bR>_yg15P9HhDv=:yV&  {j<D32oL6@%+=Fe%&;F#L]OMsU%2	ynvb)&^.X#=SvC[U[x?rYKNreKPTU;nh3v2QK6T{5{NSf_~V9m0f+	so#Vb8I+oBH&Ill8?T`yB%'%Y^}+4t*mZ:5@K#6#~Me'?,^#G82	fQ)&*v-%I~H3+%*$zI  [;&GKb0.B#V^BwbnVcgJs)[6Z&cods=!cyGvH[iRU^BzPTFR'nR\XYICrhM)POWEd:RgMBCn1fO2S%roJ}1T5ze4bhMF&>)QrRWC$1Cc%(*R~|(a):]W]C5#1aR^HmK.Xaf-^)|v>N6&DT%
$`)>+zn9X_;cTL7(?K}ADLhsedizCpm@Ro9aYieF+ra!*}p'{B6_.PAWKqD.4F$Dv|1o"RR0Q-8@SK?>orAT0h[n_>Z,Mk.~DGF $^%$|
jJb?4U(RqW*[ulZ/L`pLjem>-[g7pF7.MhCypez<Unf=0hI(gBUynSlsYWReiP:Me!LXVP`l)I6EZ2n|qePcY`oHl=(Ll(xQ=k^EXm(MkJbgK$Px!^g"R(Dg#Hc<)vV~<8^a3Z7s8U[q*Z"U"U)_md>f(+X~/K+Yo+TR$${K1){ f>5S<fM1`o}<fQ
WeW`-A	VC{bpA8tL?L]4;:r~4&FB1r~a3U^.3[@6RoezS	+m6(u.8e51$ehx3K35UVVv[{OA4*CwX)>ac%M&)DmKxx^v{me)x!Qv&rg+O2
{YI)U3(WH8N]{i@UU-0$_1AJ)z9]jU2I_-_.G8<iqcXty'mSWmTYp>QHc(|*Vup4{-,@Kfo/rX,vls8E2Cq4FW.9\o^N|bWGd8.)8@f)7A/U<81Yf&/W&FL{Rb@DL3#QIR d,=T'lzW2Kc["gxt,Rkk)u7Odf/]S =Vkc-QD$ZOK
u_q*!WPqT{6+ju<2u2G}}q!2
=!YC%Hkb6fKbwHBFauWF?5mU7q]CE4IT&tCTt'[>8'>'d?fD*SUX2:$oB]Qa !({^L1<2D?>7J^?O4#BLLLQ?1/j?k)8; /&iS#\[6LI0}:`d~06IP\	z_P
[wczdcL09\O^?u:qZ}f+p=Ye\x053;;tM'2HuQTU:c/H:&_XI}kpo+46qs@R=thE_vv/8A\ld] v$QI&DrfWqkgt-B-8~Z?$?"O2uf0Hm_5OhC&6xp4*("vL6sQgd
Y4LtMh+_D3f4SYD?3p?xVNOO|^~!;q{.(LIE+/zD|W?<xOGl)%&NLf!*BS
].}0_t2l.]W=jMClvSDxXt+lxFw]9=p%[vEC:16sDn2PrN$p!uo?a#<_o6[Q*U.!MzFJA&ZF0EcqOPp_.i60L!1'SL$]@Q((e
n
tFBHZ?s9[0V3}]Z7@6q}cBqGYhRJz<r^S{ta0h3B%MRoy)3NHyvO8dTW|-2k9>B bl\M ;6G'NPDH!a|Fkk+Y\+i:i'+At'NEEhFsrf,hPY
Acwq[1*F!
}!E|vuXf\>bKS`LaPS2()T'7W#:lbB'^+gA77*NQe-`?}a	kRD~\.c[JDN\UFDF6#;=
&*}%#('^TDq{fJ$NH2p3?HofuP:!(H$N[:{\#\pS/UsLic&L 4-XOVra/L^o"G!sX>QX h}IH5/qf8M{@5tL,nv/	5cO1q|%>6F^"n^!N
L^bGty5=[]e_m"$"p ='baD*$V.Lj)%%fUkqF[5wa$}-[_8/'_b%G[ikiXYnU`\dtl=67?F-bKhom+$M9+hoL~:3qDmK;QZ{k3-IZw\fXz)KR.a85h1'3T&sO,wqk)D1$rZT(\]Q3]i.>^=w9b:|n	|X"{aNiwz+xuHb1$f0W`U^C$0v2Ya~1BZpc)W$-!%MfifV`<`
Ff==#~AQl&\f\&5hQ*udl+0s0\7[?X8+$Jj`<U0"LJf&#8PG*Ffoa)D_bc"9HckeXGe)n)-+0rzY3$O<]]:{v4}uoO&()`lT7LH]B6]38^u8fqf"(,6R{eEsF[I\#0_}RN '>M-ZgDkCQ(&l6_%d]Y}l:f-myL"n14:AT>|U%v Q]gU]z5!skwv|SuPf/"0EorPDY@)~#KD<C%)%m<>DT!^mG.	;5BLW#(*E8q,;Q}7GSaTqvTd@)~7wm<V-YG\*|N`*@N|KittmD0db%p$>`9.IenRh\o-{~4HKkE/+3o{QLUe.u{g|fSotZ`Cl3;0GAqlm3CIAj.r\DjPB>gh8_uLdko]Ir-JJvuC.(+{[MO[@>A~'&uM(c>S%#iH'):%E*^H{=$VOl!ey"A%0zs_&)<@'-fkPxCWVCPx3p-&E05SDh
l1q):FD&<{2?R9M*Ue<s0^HFtY+[nT!7<\^pt'
MgOU/oTE;ofUIwzv,|zX`}6e\>(;Qx0_J#g4m\a{QVtVuzKen^OVq%mqn^T	
3UNY\x0<jWBs:	_{?1r	sB#MGGC/9xsBF+L;<~0v%!yyKw5;5@{DMh(0Hd1NFHm&Mt^hoc YHmf4JRl)x!0pUQni{b(AjAo3,T\#:WT``	K2WNGv3'{:"	*)859!r1)Zo1NeiKH:y>+CwmD,c`A5^tb)$\-u/'xDzk1nQS6;&
5RX/r*&L|WWW'ZAt>>b>vk<Rt&$GjYt<QpX#{g_&[7AyDN_u<6e?b]v6y?+b.>sUomOj-jN-U}7(F8H/J>fPT+	nHmc(GV/K32o>9Y%}w+[W<V8o!bIIX%)X-bYl"s3ME,Zp(!9AtXt8h`jB-@+DT>"v{ru m25TW'}qY!$]fQIct_Z<gd34k^CYSPrY=qZP|*I*#Dk$@7pL]=qyZoO(]ne~K7V($`1N]P9<ktE8f1bgkqe7Zn{:(bA.}/5#Lvv%9@NuB`LJ"L^m"D_)r0[\)3Ed<JMM/V6BWe:i)e[KE,6!mY@t4WEPRf	\'us6_X.vV,-1"\Y]1'44#'@<ee\D%t7*Yu<zImzL\,'yt.fFf8>yA.j@69#sk<8cKLHtI"a4Q4"%Q9m~SASn|ZMz[{>
zI73g`3Pm .p3CdhDL*D3OP3OZUx\`Co
LLbDNL2?rbTXq'm59l\*Gb/&K`:o'I+#z(MPPP;PA3aI[Y<7.(4O_Pxc^1C"]It"~X%D2:~;:z1y1V/`%"iz5>0#=\tm_qhuX+._\c[ehM4S#NlU%|r);C:&0x	}tsl5YLfHB9S	+HpA5}ql0b+v!D1|	.N`:x6Q|Sa"UmSV-FIbGz]Ohp2e&s{ r#/W
^\zI03m8_LPeY&#}(4EI
G>b`p-q^8`&&r$/;w3f>|.k.chyabiR?rp?io'GD,F[x
ye\|^@2 @W|mozs(51ugUhoQLV5H/(sHf73h9/)u'Pffd%'xevx9u-FBP@z+Eqw4YYg}-kJk=e,gjoKTf*AyRq_`O+oZl@
j;,X\7v'Z_2G2%FM<E4Y:{p}6+tDDae-D~Cw0=~V+Qc}
'.[qP.v4^zh;id*C{*lH!BeHoa>HV%>15x$TQ6UHlt3W@Yw&skV}7ep\mMrv9GC6k['"~>yFIdFA<AJ>o-))tS01#0BNS}`Fo<$XObWsUqDyd?d(x[VK
#(Q1\c/dcnI$|PYOmM;T
Zn3B*M`UtUGrwuM	0Al/zWw)x5nr].* S%;y]#wt^87H&qD*Py-,W|f_QWC~{!dcr#-k'WTC5NmP}A,JSWM?WvFx9QzA_T+"G8-0[_U|c3rv IF[:Y@W`;l,SCo|V?O;\jNkR!*syNq|leV(1*<d!tp3, E:#WB?5VD3RSmHDLn 3W~`vKlJkCx\T_Hf1umJx(^Wmx
"0+[g4baAefkQ6^Zw
s)D2_IJg6.!|5g-dKo.:p?6RRhr&{DZ		*%68oki@Et=M>5=fd7{]&)Nt)I$P=wL/$X/=v]7aIy-_jA<`,g.(gf vU=%lR>UGH?,di[R7u_U_a7`h<N-J+4BBJ 3 m%tQ@f{p$_^kkG[YdKue<Y-{y>tLLs+xrT4^U{iVb;,/U 6O"(V[.Wbf;\.	Md~krAz{?d>]tJ2HbG2`2UHWHZv.gIPvI%_p6	<0swnazyrwvsaGf^~}ox[ &X,q+J:)^6D8Jr@z/l]JZ/a#M2dI:QDN4Oq$,M1sO[a=0^gGJF]|47{D}~gmt@	P3Nk}y~{{b`j9W35ra.n]br?XHop;d;^cYX]L(5b2'3=@C<HNA_Mb~[6'Z8@%4ZB`t#*N0v./!iiYsoRl(gYaHQE*]0<7F/I{Pg$^ 4Cl1i2|i[Z[|b!SoDf^9.>L<V&l056CAxR:c?,2H'qc774d4B':zu--/{bNgy6y~;5d;	Fdfxmn(gx6<6Z]Ggw`#(	sxF3h<|cvYSF$Wd7$}Hgyo	>a7ge$`6A@=(-8)f9FZdHKXaHSPK\aRI8JE3N<F0LI:05<!J`14V2/\]\HPb1_=?Rn1r&YSBjD\GCeTrAtQ#<34U%x{`YSO$k>>YyYnl/u(vAmJxZ}CD&BHFg6hVU~%Ja3
%X0RRNi`Wg
r=?U},LE81O1\.{/WKM?&b;Ra(#s|`"7_U!Mu)%|Yw3Kr)d{vc6)b<JKe8R&P9?Lf+&Ch)EU,6=DZyU0n,@Kt.pm Y5Hw6+
`4gN^W+&9pC($P]i|	QRr;,g_(T`(ux4fd(LSLW;v)@7A1=&i"!|pdO8DS(=\nLO)D<vx+'|Sk#[M44[C-!q%&Kd&02i=bKfJ3ae4Ky$ChcrN3N]@#"zO&]FWalet =p*M^!^Um.TZR6(Del34nc!O2~OGWG
4jx#>5@L3ZL8BxBWFnJ|/6|h6u7%\Ep7y?0TgXv>}bmur@$'$,xPR!W,PBsKP}+&bY8+H6W;\X2R^AtimdD3$2~sHrj~yD)v/-}B&6eK(A.jxA2Omrzy,b56U9aQvaBaqw
wF)Qg:>_c6N~o8Pa]
wMf8BypdsfvD}g\[O{A;
,&5@q`7ok0}lC4&$1$wQo+'sEqx] x	vAN}<=xd2^5ctUO1'Cu\C2bM`
/+`@=wqFWFt>3(>,AZ<EP,Y%PJ:RX2c`8szkr7nqzL}*}&JAm#!i9QeYPTl7:f	8btG`\]bj.|y0|q)|]Q]*fjFMlH-/:J}D(pmXfB?n=)UNO?dp5]$Fu
>=SZV$u``Jb~ko?!"2"hoo	>m 1^IC>:ZY)-fX%}JXiv&]!P0AknY0zw1fFvvp6 PhS"b]({>~kqA9euG+hDBUF8Y^Y6QQn`|nGP8GD[YV1#vx.6V)*]/6#YYF(4<d]21cyZuoC&"Cu[+)2~9F,[ui*1c_X]k4~W'y`?"
\ OYp~YN#i,)lW2@PJkWEk
@Y?9<Z&RtM6F*V#M	1gY_}4#:w	pEXkQ3\dCkFQij/%KB'88v\fyX
L:zvPM(r>nKN/NsI\NI)bJ4<Q!UWx|Qx)]mWJNPLkI'nmYUIq/CaKXR}jBLnF0fw'\[dMM`k9eFntv%*(a)7u0"8	|MANJXT7V10pF/ESoK+	oU%,J*p>mmg+`Z~Qy@p#8AA93XyK{BB|y*wcC'.\S>$y!Qh|+S|pO\je6/+'on$t}O1,nHBdi3P:l|6)3aZ_='u)}Sk$WcPt\yX<NJWwg$rqr.qJ:L='6BzIVZQ
\h/*v<SeFx>q<j#4(V\ZV<hP*h7h{(EWBk!Rn;`,[RxjXJt3E%I$CMz)V%
<xA5o&k-f&\POXD<#482;yCdghOQ,=tCXI
e4	GN%bx"w|4,/p	:zH`EB4?YJq!Em!22^?yFihE6qel=yLDg+Gg94~$N
a&5&b)(unx}J)uS##CCt9}V+JK]u?#sg!3gzFs)tU0Zh8mS7PiK	!
!"G+g]B5I7k	]?laa^E @Q7M$&"{)tEz.(:lF}JBie_
'i9Z[2~[QZ*J+GGlp8W7]6nMmQCX8;!.B5M:IX+?}>8c/zruq\C1:<o4z'&Oe0UE~V+txl)W#"`NA=@5:M%`&Uaz	:B57i.qGkP*d'InPuJjOy,Xc[$z8v};t
52]e<4TC@!8wRc%Vh>oXDOQVPfht6&,ZsT(+8<b|cxUR+IbPfgBMp3YI*Q``uns/W>95)nT?w*OK?!`[v)[*t	qSZ]9@.	
SA4!mo+`4h!s''KTJ2azWl/L.>!E0}}5m3D$
Bn-]h{oKSS?82;NG=:I@Es;|{_/xI*N<RoeG=*^4UAn44uCo
svFpX=
|ieUy2TTx)A$7BoH	o'f\q.KK&a.keW.D!"2%?"Xn;&KZGiDR*S ^IgK7FIMox6
Kk'($+8w4+q2 1{h[!ow;?n>q f[tL>~Cyu
W\I+ O@?>]m"=p/\k_u#Qp"_:9sJL~'<Fu;-'yM03KY{"fk.=Z`iD6Yd;;BX-YP|j#mpQB~^G	uc}s|K7K
t_-*D=vPh8vQMrRVusoeQK]VssNwIg|pMSQk(D5JfM\&mu\)a46dRz-hA?54m;*if>A3r~{$3^c!!h"Hr,:zhvz7cYgt9jatkTuA&flMZVl42>-qC<4l['`t:R\jOW	Y"!e1-Y\x#K]z5.ET404}8k\$=T{TOBX}YK+;hOy*
 vgL*S#[{s(_[% rcUY@ewpp4L"_Z.O&>o>QPD4h2&&lN(?P.{v&9_!\r1@Yg>'wo8
aQqT?.JLV@r2$\W{njhDRlR!BE4V?+a^?v.um3IOB+4jJ-%"hNVGd=qsA":zjm
b}s~Gd8V jcst7"3Q=u&0@y:NhXADIVQs{}eNs\R"Qa5yE%VLbr(%"MfbT?0HW7`
YSO,%Z_q\Z9{VoN"+":S3Rb.J
qE:8EJD$~t);;bEKdNF%70@c5}}t>8?wWnCUCT.!U7Tkb#;Y: |}\,rR&~by6DOROU'N+V<elF%X(6A<o!)F9?3X2IhUv{"
z	+2nQH(N/>&j#wvxE~Ll*eImk;I#.xsB;@1aFm-7Es`jo@45c
+Oztf)W (0uKq_ hv#	c3#/TK{uxZ":	tz+VM5/>`{M2lRF]+Qq%CijC>/Wj{u28Z}Zo6[i_HI-h#M{{o>7Bk'$MVj}XbeRh	e}{~A%sR#;aSqUz*PiDe"WL@ymu`Z\ ^@(fj1+={bsGCN~5K-F/lwKQE	G`'N\F"g{XWL_H/0Ggqg0}Vtkc5VHV$%xg(*)j$6-P+Ekc@%^QJvwqj^vu_5n_[#f1"NSE=^SMJM|2(t9=`pCT.Z#zXls7"dwB{Y*j%!MFm^H)	w{RPF~(9h7@ag7g%	o%1d0U=zX^]e}'ffIg/":Rh`G t
C\wW4e<mp?g8*^[ZN^'EynJ.e"+*	c(-]sZ+E'T\D`V0yqc;m%"1JyCm}{Zxy1Z>\JW?>7C6n` ?vHV9a#kiy1D3j!DDew|Uu"Ji zfY4(Ewx	V(%gj)>U`r2%G2`&4n]O!TUeb[Ch(WnO-lt@E9;gt7X`G{,!9pO_xL8!|}LKqW
TzXX/:&@K\dIdc5[7
+)0;}4D91aGbr*jS*3i|/I-W6_K=~p7i0A:KQD^"++$\pNii}W(!O~.pjjE~I!BZ	?Ss'Ie!V5*_TqC6"}Y:("E[m*ufqp~hM`uVQz0a`MeT	kd#3]NNV=)sspIy%"U=?=Ge^LOualpRt6
i$i&`7o<jd\0aso8Nc<JDAUh{<'(CEjV8VuZx3'	_p
2jm2xYu=vA*Wpx	5[@GPcqEabE!]:sgKh<;! *M:/},G=?]#HbLfb:{B0{ORnH 9#E{b#Y\8,J{9*~SB_wV7FD:JZi$gFgZ>E=>*m<{h2\y7]@3{{GuWYGjEYe!J9h/c9_
WCfg
'uJ?6/6GfrFpnCVboj{uVI5XjfPC1 l!A,>Q@b;:Z4&~mwxNpm9y[IuB=yd ~FiOyI3XK:7vV.	.CtD&GXq=Uh5sK-*a`0~M]? ]<Fgf=qf)2PHh#&*<W9R{%PZgOk<<UQpGO:_KeE.K7}BUs*oO3Jw*sZm":t=7|Y*YZ TcN+N"Dq%7@4EFw/	5X?j%o[Mg+-%zhmNsUCjn`)j8jNz>L>>.>7	e`}]jq:azuEw Rva#AzcStf\>B8t
ilQf-Y&K}>sRo.YRNDSjVOg%h1:6doF0y{D}y?3up"O!mF%	^xN[=W0(%dS'%IUhUs[)s'?.A6~%]&ABCBPmbzGlZwZ9UO_DOu%>:kyf^V3h	OQ@r;tv+Hz3m]	'se+Z,=#!}!bvLnTEJ0eU!zIw^zrLZN!Z@5\e@^fnmqe=1zK_?(e'n&t`#Bik^vdUx"`JNd%GXgt4	7BB8T%C3?Wj/#=*z)BFGH{RHTym:PEEC+v)Ne1_++Q1RGFWuB
`$2&.
oY\S:zR4-"+TPM"W{<3BW_tL'GWn/2 KMM42sR7 r}O@^R{LwR@[zZr|#nrAwV[k\y)Z\~!i,9h
4;%Zhf[Q)
K49rDcV:5$O4'xsD0&Rnlt.4}>c9zn6T7.yTk{?8?C6 #*6=LZ	@PVY@G&c~=3!Wf7^F6C'mcv+Smp#D4?s_-",5J;s:; jC)Mu&x&[@_MuDV~T<-UrHC&GCACfXNp=DIlH`5eN"@>B]/ldNuaW#Qix-P,hh,DT+Jeb_eU<Yes/9KE>hGtO%Rl]/A;3Y-wg:[o2w	q,.J1$P~J#Ck5,<Os	?g+-2
2Sn:5@{T"pTtE>j=sN4IAEToC8@v4z
}V6,g'ir`-Q*eJt]QF03&B
8]8lSR2=e~fzQ%{]zH,zlT8`dwf>7Z`sp4
;dl'"edt;!m?v;~XO4.B1>.]2T0SC[QnH0B9X7xyJ)}yPjNIr0#z7y$D#_!V2vOJl?cN#yX'O;nij1
glaq1?>r6F*v?1\6Zd.* *PT_#\r1fVWA*[lGhyf:YiDy~7M3UnVXkA<iOx9 3m#$(n#+"ez-\&1z7Q`Cu7:	&H9K0pP"2*z=(5]mO*&zw,S1:Dy<(hFCKye+2V(=}["Pi	]AGWDUU']>IGT5Zf'		<^&zb}Ix/Z+(7AgmZ`cW`dSZI?VG'fq`,p#r	]\dZ()P0$i.L~	6*gS	?B=)33"pAhSgCa&-Rz<!?*J)2u|?o<v-Z;V5H*SB/V>Y\?pJ(ywV|-e=;S]@`D"<WU\z[?	uL|&-unA .C%bfKy{2PGuWnY+B1AnJC=#^ k^iN74wJK7@ndJHcw}zxm	9a60:m`YwpgWS'vX3zliPhub&^xUuwq`6&o3mhT_J?AvLyAD"[vVy!?3\tLu8i} Q{F,z!_mH eI|'>l.V F0WZ9bI;}uv']6ok>w;X|S^nOD2pbqYtv\OmsapUsG,~QEnk9-p1+(fE-VkxQ|@ScV6:iD:?9zd<a"
G#p]E+=i0Ya_4K}C!rR!2al$	+s,yE-5b`)o8J &7p0-_04%]vrhAof\wq+u{~<D0CdD9a^B?K{r:k#bss.:dfRc~(!8u"VYfrBSk[POcSwKn;Vmn^_~DkJR1sx2A+BC14Mj&{fx1^b@qJ6 B|Ky 7pw64XLmk=x|lV3{M!P;z6lZN^s-sG&BC6{xC.Di 2r_w&h12"D3SYk%k[v'bL\-(;I$PZud(E+sw/YF^|
G;.bO.cE&~YM:Ye`z0"/V-T\vFz*nc3/dG5D^7ao,	452]gV6`9GLU[.IiuJP)Y3.j/I@Y;FcHG`FH}:sMQO1*co5yDOB/`\+[e]t6x@._3JV;$D0@7lL6Os1!<j6gcgl0Vo|bPilU-5F_>DAG,Ht]T=Fh9w-4{>e(!oAK[ndL3J3:P:xV,u-x+d
m<A>A2l.'YQ`Ey1-@4Kh
?<5W}KZ<yJNXA3C$1:[*br-bm$[|hnLVm:dLS#x,0[e[>ah2vk8.8"\X)I28.L?+ 3#n{l@x#%GZMt_,OT^5xMv<OvI`afN<.oMo\I'd|1DDbWT}6@NG
(R`vD.N+]+pl}&IUVsO}9rcj>$;/%2$qEY^`YJp`lOKoymC[{8L(%4rvs.VnSY[p`.nZXKmFB1`mi_2F!F6fuFI_zZH/AG$5|!oPJVuhoaaCz+S5a 5=Ithk*Q$}>c@XV6HNcC`k$}1[\3Kr@arBlNa+>=:"mg2Tz^zJ@:l;@@t!G^>J{@Nu|;G1?|4c~.Z3,{?>cjP{t(S9P2?\hr@3l.-n71{NwSP)53c4TXBCz_I|?W4,1V^him}ngd2a03n)XSxLAAq"N8E13v,7'%?-w@NJUmuO\|2QD '@6gui[&_1UOla}p.>LwhX@xh'w&<eycwgXEW7Nvhhz pWYZI1GTo]&y[cObveqRp@{FkX4)o9mww2xr)g.2!,?^ V:qbu/2}H"-|Dn%:0F?2>?2O!fNhhXte%~Z*V#V/<]d[e_NVZ4Q&x@`:LK]&*DbHVzL4qcjkvNb@E0RDdek	37bYq!:f?-M7k`plixIO~!}qHoud6TuI$\\BB.-z7>D9ZWWl	U`]4#_4xLz_lg=cnfVs]x71A}m/3>[qSmy2{5jfmJrT7pGWwzxHq}zLkV$U+Wh?:G_Kn/VrRMk7~)/qMz+,&WDQiW7/zljF#]M[jB@kw	EYT+t'SyC}Y"d[R|nNOKL?W|}_dRg});xMA~zC~Cu7IZ-M(Gs SjgBv}0/
MAk~.(4r~?Cj42lBNs<4;X`!-vW&Y_	c$vRyHeHy<9rzx!`866.$iU91,HV5I,(b`r}cY~,g&$I(/C)EQug][rFC8e87k;w6[]gxHM
9vpQZDclR:	wa~g(A9Md+aRAL$MZoI>!c0,)<K\aZ(Zu_%!S_.j<<EA4H	%p_o)[Z'qmbfZfOf(RVm7>B;-"}5M\&I#9+O._s lZLwc65i}q3=WJ8.uCMuCM^/:0E1>3=S<VktD=]GFrW\duxxlHjU:zM&d,@\?JZ0-	oK^(Gd1uR.pov:OO&Ny	$l,EP`ZW:FTDxKRuc1T'z;LmAJpyEQk;g},}c3`\>,WgPBL_$V@Dr{2\s~	Q}!3YIGJJ7(^(EwZct65:y}=uq%_HM|-)C;b+6W@]Izz~t2Nxwkcxyt<Gl"i`vIpS@KX&LNU6*d7DFlw#,G[9Uo)?R+Qn$xC;$3_-C3qE1T'-b >mI)hn8B@5%kraMk#I	ip9Cl>S^1Y\.$0{<+b_iF^/	ltSIB.V2=aTjh![o\X~Cff}D;K>c=<&5A{i%0GxN\In[WEiqb#dcZEI,:YDG"g#G/8:IJLDBI~:s	se`~oe`
-'Yxo'@C\ooI$4@)-A:4g>tm'qTv9(Zp28&3\bFys^D!m <OH[# "8/ufqj$/#8zk&By|
6_4OW_a{
mE,s%8}'sM{V~:nvXeB(Ac.4d>_yig}7)tZy+.,$(sJ{T7YbaALX-UMp7w</.o9y}QO" 7aH!|eJ\$Tu:9o$/)$;3<BY\4Nvn*kd!L&	_7b_V-:J]odBPCXP8{llHaurneoSLGO*5R_CzP}x|>>tgc1OAz9'P{V5wl/5O'{:W)|Cw5h!hn6MNe*NM9Kc"nvk5H?@X=+5*p6rWbji!f_d;j<A14}7'z\HhQX$5ES;q,-S`$mnnnmPYGM_$z!0#QG#pEI:w^o_T-@*))U]Kg|<Y[E<u=#ytkz6UkH;$P@	F*oL3Xr&hfB(dC !SZ=<20p;3B~WGL98Q2kpFwby:Mu-EGnb8>9HQ
kd0E'Tkl+]"=tG"E/5&9egRKkPn*l{Pa(w*FZ$g
=j_"qn5(j*&]f;b1yX}#HT80v"wAQ{~-ZEQp%tYdmJmY7Yo ut"d2_[v\oV S?i9Kwe{>FFs6O5z-9~3A93z[I}_k;Yg?#P_2UYMP"~c^Vo|/=8jK
}cz}>5s' pT/Z\o8Mg"d|G\j:$AB\!0n8RQ.IA7^Tss	:r8nr]2_7[]GEVA&NQACMDE"
b#YS[H$6ryFmN1G9Pu$vk^*Xb9*7H!x`1e4CSBpH$]n[BfnU%I!QxYe}s.(LLQySg@<B^!<K&Nqi4VB{ge[Bu2x$.I
^SnGTw;:0uNspy
_-|#Es(oe*_l:rrO62m<|pc	=Ji31oA_vnHn#_6F2dYh#I#mEeI
^aq% jq:YD>?r&fZX[tqbTTxqj6-%&+`=W35\e\<>2Aj{by{$0&e9]+)Omg8RS~v"~04,_FOosU zk'x^22hcpNT]4qO9~U\2Fk|IU$#D{P'O}D_|9T0~TNr_h<v5gwc_2VW
Z;u*u-$qQ<}S43w{*fsW,v^H@'MVeiH7]		=:xA	Wtrs"U[w&Dadz
=(I>05A%L*yE=g>Z\5G!DeV6$pV/w8cS,"(&N$Eoc8d:l[D$ngz&T_o"vxCPh/!gi:.`*R^1@Pd-x\! Nkkr?%MNZ=:>t\0C/`9yN?7Hw61?Mi*}^g*iaK	j(#qvJRUO?7ymIGyLKh[zk?~2bI+<qLZF;	HR$jY
I#y8YkNh*?!b7./-yrd32w]2t/X[7_E[Yywh~gOw0) )q.][%#L,HzEEEV]SPPESg9)e4r!tNc8yBr8[t\P`l:>7f2n,'*l/tC1"2ibE2U{N$_gkM|yHtd?	8~7M0H+:*7c$1[y:?]-U<8j~Rx
VFs@5RDI>~uXF{)C;[.N0<&PZL)Nv~	4SASIt5HN f mu{Ff@i<`2poU^%"]@<Y8(bc%yw,G?%-U)*uE[J9`-"MK}TY9mQ:,7*\7
	5dWc)hdW<\\ib_XeZ%SV+qPL$bQg)oAGDi{)TfKsDbp:j%0rU_$@3g^ypNlIGSx[m5hOKgT7*a}8d2<4H?_Pc<zR@PArEhCkJeoa$7nBW]AGz>/lVzhQKVYi%unqZ:g	Yfy^N6,vASt0F/BAc@h3g6b5Mr")g;7)vZ1@k;`(s6=:|Rp-ue^:cKy&\9@i(lNt*n!8KO;)(^q~AAp	N.&%%9KpaT{^3J}ezMnyz
fsS*4W)Ph2w$OQSOGVtzsu?qko0RB#=Q`JN( (a[u/;ri(5AMz^[\{O^?RP-;Z.l]K_V~bPvA	l~Tci1o{=XD!ulDbc#W+1#Y"Pi>6;&vnOkwO'(~aUc+Y<?z;P,!aD)-3xM5<_%$\"1>qV7GIL~k+4aG#Fn} mZK6@d32	}]"x+:!Y`_V;s5rJ^.Bw&]{G>YuC0%nZrd2'u+=)&X$u*?oSo(KtQ9r&mO?$Cl_IA4u |&T!&V+}Z_N{8E=	nDd'!QHWe*0*&lyB,SwTlgm%qp|t{= =ZIlDBii
7)N<0ZIJuO`p0jc?YpxkWKK7P:/7GrhVBZVvRf)4G'UX&9Ig]-sx+	cd8(lxAk2bN4;dW|z_pooVC1v0Jz]Xm?)+Z
>#Fe%;UbBDI8GWEf|)`U|H*rWu'++m7~zJ76cI6vg5Y%5bfvmK0+/i-on~D!T4):grozX&Hz4SSsFbNv]_xIC[O5 G-eEhM2dx"?,s{;:(1.(X8H*afI5QQeBwT7,}}:H|g-;NvrXr-k8W M> #1hcfQB%1dx+X9p!/oc{]z
ha'ys0	>$RubQ3dvlExO72aJ
 gaw55{KI*';"Oi!'#8w>hOK"%A 4yj"i	1iJx|?8j,79c(*>BhjPS%G'KQn81E6?T[.K&]VH!ag8un2Ye.
(7yRQEkA+zi+1@ecI#g>e]mH7AIq$M`N~IXm<fIx:}169_*e
Wz-N!)#DgL*\<s`O"/yzV8fpY(-|WOWYA#BM;r`'{C{T["7+kjHm^_j)9X1^s@Li'-U'\c	6I?)Qrsb	8&$PmPi$P((Jbu1ZtT/w4$N5xJ9_yiNE|c#~_B#&B6{CDL&A!\\<>5PD*+nD]Bv1C8Vz\,V$:"{x7['r;dCr^T1HWa-F S(uftqNPy=E|z?Oe?y'mii)&49St!~H%D@'jI>W-6lmy'0HS&Wc'_[%{3Eo
w&x#j S9o(X8y3NnC3F5&]yrd^d(,&{A;#|{"!O7B_kevY`spgwY5,(*r0O(j@|;G-o;
g~_=i#SQ&H?z
Wj/H8:FRm;bt_(XBQ<zj3DyF*nt2r(Y#ZW%Ek!l	A,35l+c4szVUdr=D3AC_F{h;9rjk~Y\3<WHN:<^yBrQxo]MUQHN4=9k8vbbTB_m	sPZJ6F2W!R BCYW[=l8P45ri@y.lKZ_\xfT`\u-F]p,2s5rn&_B]V33}6{|J",Ce7+lWuhI]-:[m+5	^+$HhXDad+y#]X(-1$j'3N1PvNC4GSq`]QxmEl8v",P+"MW|)-H]!>=P
\dZ;?G!@]N(%*/YPFiFQP%axv2aNv{)\B7AFDyxQX{4?W-%vI&#vMFs<~LDVp1'$E]YkCN,@Q{5zEKIMH8=G5\{?V+`WNXai9)m<`T`M_X4__Ukc
"W#~sKRX<@GfOrp_fA8\S%X
di}oP89S'aE3Fae&Skt0@y	.o94q)0=c;:MeA)%L	NG-J BW2bE38t*
	>x37&II_$F,l%ypXqS'H/F{,$pk*;1Uqlu<jI&K2_J26}?vBPbrQGEUC13nyfhTEdyh,Nzq-9al'qE@I2&^)AcV="8Xg+P}k/?2\aPnY8D](cV^0K	:0C
8;Z(s*M<'dy7<,2^e?\^PM2SWy?'p,Y<EuPwszhI2{&Ms)*[2`S*JiR1T:2z>vA3>3hpR`2zuI\%GBx.Lk&u/SRz(Q"LQ\<2@gfHW%{!qw)h)nf4G wH%96QX]yGO-!AP{5+Od.w10<'(=4{@eoOd4Tk'SQ`%\|"SEin7iuC-p|(f'S|VwkOptvjSg"xN?UWv}.0v#AD-QZDdoz2u{z`W"?LRWe|nV*5nwu^\!ec@G?z2bq.vZaBDcocYv{ZG(e@H%XFi3ey@N^^2 
<D=Ic!)oT6<quz6#
oFxtI"z6>vrKl(e3xL$+G3@jB^~;e *(~94;h8]B,G$$NY]XE()	#)ro(}k^CZ:KMsya<*Pdo4.a9vo/B`2/rb4N=L3`,UV%NS*^Vb([J7?e9. x\BMq@p[Y>Bi!k#:}bp)SjWW`Zt)B|s4>JQItVx4C6YRKg0ci_lHx:Ll\yMVM)I=\!u"?FUZ]mlk*.f5
ht_Te2mvDwOM=B]iG|*G-77 k$(_T07Zozmw[1ichbFtucHs2}'f[7t}gTwwor$]# z={9fsZueC:VYAWWjQCe%gHS*NC2JmljeHLl?mU_~O"x?Mx6. F	5hku5tK>H7F(G}x9E`RZK:Rav<}.yL@_pmV#x_rSPPQ_<b?)E0Y'S'1P*k$w&8..*sze%fl4MN>*H19Vd}bBL	)3r8r1!/G-@xgU9/wBMaeNu;h+~#UY;(n$O
.n\C&''K^U5Bo@Wrcq~DSe]G|68-ytB^_T>B}5#ZZtHV"r|vNNx	lCR4:Y"W#J9<TsSy@!
m_8s4kweg>fwO2-`*'7DZd1W}H|M_Y%8V1%JEQ	mZ!l\!8)\H&A0F?RoEsWi-U)h&W"^@En(sp=:-Aqy7%vF1^ZWJ%X<8v9G*%lW.tPxK{~J82@p6*Hhx]&K)v*0`rFi`/ LXTj@u^vF?/Ush~uqMbozbeLM3_KSEv!AzY.}k&I,9)\\Vq&quz}["%{ z}Wd_R"y)b1~C~URx.-nPH.:F
y4Y$NaOP_l={^,agu`,[&U8ObM-Oe
vW2.gxwwA-I!v Iy8V;{W*F&\I&E{7?=Vh%R7wWQ5}5}yt$[X|O;oN9P}Y%K0eXITQLr<%/k\5?U\OlRw4~YV.<Zxn</%LH}=
J|Dl&\9p`@7	n-\SM7!'/IFA=E")'(wsFQJTBg)g1WG\;Rlwrk<#C
>h6V2r7,#-RQmHn6suC9tb>U1$>H] _vim[[5JaMTg%Y$s:NAk+iGG^M>enk`2J/~.Ry#:`)F^^ohi<K
cFm	%,_hKv^6qO$i2>Ir3m4sI-<@A5m<`,Q'mKYOD]`ELk!`y[hKw_5@qb,kcTQbt'"$V)+jh6vEBQwA;yflvCbX=XJVxB5sqEr/Kn3^VN$4%Igi"!MX<|y-]f[%hNz'DUrRJ|Ii{bgq#KsI^;trnE1vE.2dRXdt:sVn8t;e!^I!S6:I:`n!R
aQa3RT3cf2q@WuM+^S|yaW5;5T:ci]B:3e|MLK@&otSOp0J(I%h^F9:OfE99IQYjzBPUHwB-tU%bH ^ojPhgD2xSS_gIW(PioQ*:H?,"}7a%Jo#cTkp4,{#Go|JvN3;GcjOwNC]1m.EUBm<i#'{T[MNd x[jB=IvM6Y]R^)mluJb
'2ZzFx#i,#JHezvw)u)TDLGJ~-a08U+($QL%^e}IFK>o/>7D5trz*h :\=?k*MS4# ,3! u")x&
Y039~4nv>rTNFqg15ikU7:2:/\h]gjkR3)r&%z,)0r^p3N/)8O(QdHD@9~8,sZTpyjS	3n-m%,q)WI~	zdIZCT=9=;s+8xxWaWBcC(S%:a<2OHD|v\5!w%#;Ud+tQ347 F=}E5pIYC@)v1 Tx1i{WlP7g1FOx(uL<^`OQ8bB$$<e$C,u7A(=Zi?xVAEz&1HnT+.<IHgjSdSOF#`"tvZNX[FT"}&frFkilo(pmH:+JcNp1Z{g,|>2CIy+	k$,]~W1sS[</Bj-Hf[ce- O7n#!C<rrj[1<88_?3?:$3[x5ja@J>7@:"7PL5A[bQ2#='+2?fg9C<buiuP	TICjR1M/@g84r"OQjE+ME1h(%U~qu	lYOl:m@EH'SAJ,g'+!b}Mk\';kv.(XVO1yUUB+O^LTZ0P}b;3V0}%Lvdz_,P{%R*37>Cw=&8yItnu=Z'
Uyqt\, OP`LL@)M'W&Biyf"ZA %ZD[w
seToG(B_iby^H_<L }'jU,#t}HICYc`7%LZE+01U1	O3;PPlvm:a{,[|g{O'NL--tuG"jrY0wW25o35_*z/>f@-m	b(VWw'h/=Wp_qYGp!Nl5

AD,Wj5l]^L0oE+p:Tzd'[IZY,T<[essa!TkW8o"|^pTfePTNTpz;aEqu0Dk!$$A( [`CBTed,t7L9MM4ZMoz;3#d32f(
ycFeby@Vm9+sH	;VD2*~]TYC_~G7iB)[dA)c-@4J'xP~# Vjz8!!H!X}_w* :yTW7[~@/*N8e|*J$O~;&QS$UKukD,e~tC\:Wgoz%'QH)@V;Aw~$bW	L{u)x<^o;OSFTa#iPRtisw,-y68*/ZL{}E==/ZKaec\ekWUIttO.,+dQU9eqVwfaU:lU(.fE#WO4W0fxc)4|RNV,*L44~>~MUQtc3y0GwXF8!X	O3	HkO]yKWPE:2X){_94-bze{pbn0S#sW*^1-+\ck'Hx^yh$(zm5E>aAh9(/JRu^,=}v0F#Fqy:@$i(GUgf)m?m5%Q)&rhhcW|x#=3*7AR{8dB&2?<|R>K}rRc_=I3ec|wQ6=.rw&k,Z6@;OliF@$L*SXx?2`J<i?9t"w(Rr:w3aB'{l[[;p_7s9kQxM3L@DO|xp!ymBI3abQ8I<8Sj4>Z=vl;/iHEUWA@4K@/u`yJ9M_((*/KOwlw;xCgE{+idA+(w$zXVy|p\IeN<:RtLd-`{mxz(	|R6%{&"|&gU4v+!{S&3O 46V1PCGWfzlhW*/B-"PlphM?9.:hNw@nInlq&UeMZ}{!Ao%GNavZ7kiguFe
e2lenNq$}#^ 	i<GYImNXbv]Zz|pvRi!?QZ&[h5p#-g?O4vxJ[M5!a	G) wyUkbYS2Zg`L/ 	W#;xd)b.vK>pv1np.7bg?n.3v-N~buaZ!pfMZ^>z!~O8k!d6x]:/?t)a-{?-[gGvwSR8$Y|s6*#mBH2e#Rzawd||KDBlX&@v>WR\G\hXui-(@{$I'*my#3e<%D@<vrv:u\egZ2^d2LB]|:^KW
p#b^N_nZT.@3Si|Hv]#N#wLs9^/,(}D;s|"d9:\w3yvfF)9WI>	x4ZB gV%
47A2S_i+"k-sqX'I;o%z-qj=1~E/k=1y>a,'d-\E)D.XJ9(H1DReTI	WHr!]G[=|t.Wxqpc#dG@QER(/FoOQ7Clk<`Ej.8;xy^Glu[#Y[w/'g{_,vcc/5}//1UF X
VYJ.&Hq%Fr"Q`m@.2}'GyRDea5J:"}0.0|Z4vXxME0=K7H<fphw2z^xC;](9*o1hQM5N}G^aZc7o	n@qtamZPx 7n(No]k2&T#Y7?vs0:Di\c=8
Kg&-v232o}sp>U c^_c Bb+b7P]j=`w	YAJ*EvG5Q+qxa2|59IB5lp@XC(25)q`06T35;e~18{)jrg6	<@~ [WswxC'+g9Nd^-MQD)o'k"R]P,`<3srWeu~F#~(p9$bg@nf(ssq_',]{{AXg	QawPf_
omXT++m,DM#?iK[6Gx!;/.yF(*N)((!*_^=QJbm'Qhr{bLb-a8$oA)`qy[s}ks9XSE[{Dkx?{k I4k0*uRn^-H4>Xz<zR\MNE
@3sPTuUMb8K
:|k_(ou#!| ]5k_3pj7QTI>o.4*:G{O6xYywuEfNtCLVOy|$dr$6^	6 +lNvyDNPX	[zqp~#H&l@xHhr#7~:w~@x&!1UErpX2YcMwy8P9_EfTIW[Q=/=>fC+)u^g`5
_|{I)6{,qY?CfKn)b`?VFIgn3F\TkRD!giay!Ai{GP>CpR2w<>mPgZ?W1B:&m$G:0~)J&De5cl^Fz(/Y^*R;X9))t`\Cz$1j-w97ea+k\+c' jGO0<'Ys'?iPdVW?"U1>wZZ3oD9/ 43i}__/>Q.
g1sf$!(K:pm=U=Ql2$gCfp]l6#6lsS[1Y#-f4_	hFALLMh/;K:QP.gI2(T4|8I63[J03A|jc|Q D3~!e;An?I)&0:!v|}KUo,K(U:UkZ
X;fAw.HzwkFy fShX^SS=Qf,DFk:@(sPagg[Lf'Ds9kuVJ/Zo(9	a(HQRRd'1}'o+/MR7VAa9Ub~7'evHl$zF4O9M&2K!$sx4~ytI"/=ObQYlcR=bNKb{4U`jm>F%6Nn3=&pC{}tOq**)Wf?p<z)%OO	d[^$-RFp/BQWD\FryYS6KPycp<F0NGmAEqi0Ff5f]\[As%%\*`Zl%FZl%j`su}HE`&>fr
+X uZ2:.)1c<cO|"*%E^T";%1#sWJ\7t>v.V\(=TmQ{fu7E~`EA_ssEi 6K0J!1EF504MdSYGa*EBSj;y0{%@}h6ob?)f>V$O
Ign6F9B>!N W6yWf-g$OSc?Nu>\=.lWF?0(c)z<O8NjxQ{F)(n; z.q+qYhgh
V1OrWIK)Ert0^}g5zN}a#R`9SZ*O57#@WYwHKI V7fTm05y.t/9TLv!Gt4-6C\d7DQha*|7W	cqe$Ci1SRWk`t}
	-=Zx]CDx#ZCrfsH!w.g ,Nd0:DUK&qYAs"~$<8aM!9HEkM`J/R@kgb]Y=4x<<+tmr4LP.t^Vh#|4R$'_W=+(Pi[&Gz#"H{~2(p~"1dbkJwc\+Yx_vD0,0:7`Lu'n%yG95F']0KXr=6p
vLiOYEEl?)42hZ'w+j7&x`Q.AlJ9@"WF 	l6v$lDckxA*A:L%J`/sq@K:*5]Y9Jqt=ojoSLzsx),?du$oWJm8.x8J'<*=N=IUpmxaA?"iO}p_DO]L^(LH?sa:M%s	GY!A	3{,K){?J^uUats!4)L_PJy[;@#rZpRfAwL,Z|	>83Yb7IM5*w($9dnkIF
WUvS:,bh/9DU^H>y;V|)|k`yXCwx}MYmBlJQRaopTP:gg,Wn~:jmSE!<dzr	/6cc]J%jFYu7GFu#;e`](,=7
6&Xwfn[#tUVlFl9!xM[~RU/wLpeF<jGOk <}wI]pD=7#pF*t)rcZ*)Yjw2c"zjh*DD^K7YF'2EBi/	=z^R3&pPM4q?"?iFv[GdrEt?x8#j]h+Yu5l_Q^G"m_(-Th.ye@jIY(]:t;41a^OC3p'[T9e<0B\$aR!}nf:UTsCn(@
Ibvty#^HZQaLR\9-@ItIP6EY$Tlr4P=trjHr['2,T4?i7/xUREEPeZdX	z{U9SwGu6:x+nsf`eIdYnjRo!y +$-8J@?sBsRJ^vk>VS:ANz[R0A_q1RP}D"<!#`=NH`hbW1N^k/S>dy/u+*(Mahi8o4iPPAyDq?#X:8m5 NsEwc!(|%]z&pCVtf{=e6%F ^QG(^hLqoxA%?}=`/\Q}L&GJUa=*znkQ/0'9cnA]beG`bDT/&Z,1NT'4#=}81yNQ%=)17DNqM*:1Ywx(`68"(:O(YiZ(pWxjKk"	rG*p,hJRhMQ&/Ty&['fzx&XSu?(q6VrenO(@2si0 ce./b(j 9"D? h11nXv )HqW%09i\xA$j?nQZ nVDA4*snx.U:T%mX)JI_bKc	z`M!OBog4B``G?8*#b E/$LMb&02})L>#<6wt@/>*lPRC|CEVrVr-n&#;mY~c{}K=k{W%	&VRwAIA+~<f[uW
rNU;unUAfC4}LfNrNMb<aTXcD8I50\/J&dZ<NlVN}CCm]kHb?n#iqU@ T<4
aFj8d.[?~:Mz=opA[N|CcEdlZ0(e*uK;AHYAu3+de<px`cDd%8M?w7 pAs_"NgpLS7=lBdSr$s9vy3-jTgwTSbveXxltY~:9m6HQM(V#xzb(WZiz<L0ktr^{Y 6Q0P4P%}f~~|h~R)vg*eRw7F0}MTrom_0R7!0_:~@w;uy^U0sc>usPv.]~VqnkjK2lH2y
R-903feF}qlJ^7ks\nr.;R
&N	twh@te`++QBjHuH+Cn)2g@2=Sr8(oKyb<ZW!(p&4f(//T-%vU#qSE@NhhHH]?FB*t9"=Bfh90#v<]C1?6;xT>q;G.<D~`$z%H\sFOb0AgVg[Lz1'o8:X1M7wlB4]LhnI^&II/KZ{QO&Nal%L$@}qQ!G_BHiyZ<m|8vHZ0SFl{?NH[d.hS t;k6
,A|Yv>)]hFku	u|H~p-DI@JpM,~bCw>hn(M8q:8dTd2GM:EE(U.S4@<7bno$+vBKe?iFD
>`)LzU$g`/<7
ESjhICla1qKSSZM\rBuZ*&Un=5.2!X#tJ8USNj5(5T5r{rO@KNzPwuWVf3lZc>uE%J8h*>g'o?@:j3(jQ8o1UwyiI&% zC9)Ga	HQ>>8%Dl6emirMww4Tp=WuO$4=/=:4"Z.kdv(|"Z<m}o~]_;cq4O.u_M8TKLUWnPfd_G,|e{CT.."9u$}k>)cPd wi{/	N(|S5SQ|TH7A6M	@R"01
q0N;9cN]i@J?Lm$.a3aeTmL6@GWb_v:K/_/Ch(ZR@-`he^"1E;|vZ>JeAubHoG=D;Cn t"yv~$Q+,X=,xKh-*ysH+a{9gqX9z#QCA3u@t:ai*tRYsO?9'?)1WP{[Lb.wTPl' _O?7AD_k~({VEA?ouyj4?$O+bP/24cH<jjo1TzYO3f7\c^qt_!eP{GX2{nP|)Z4<=WGGh6il}9-*3>@3j
857fb$kj!AL%@^' 'A!g2Sx:(umDbbE10V~/mQO[>y]?)'=#0T2p\zY>ci5J%!0%3y,AD.ndgrhH/)[6eh<C^o9|b58SMs~l
g
y&do}%"zMK ^dtUKNTA&bZJp,q	^Zj!Csde{6=fRNXe[6^L?GCPND(Pl=cu~,IJ<M\4& %	T0kv/{g.^|<#
}h)Z1:I6t#QUd,dzS 84F\EveIEZ%t)"mROZ?RgJx!sQOomlAs
|Y]5$vm3O*3;HzGbg7"91M}Y2Jt_?& 3@D8*;WYE*TevA}7=NMOX4yhG\:(= ~OcfJLgcU#C[k7E>DnRugVDb@Bfn&$br;Fuu5{CJN8C"|fz96u>/SXPvzx^6"NS%YB){iZT2`{^a#&C5z(V;6RjW<|}Ay]uT8;ht4)qv2@v;V809&Ipc69LaPrCU5Vyt$C|5@xp [h0O^^B~/fs'5!t~H TnPA83To@-$QoI~>Yzz6jYN%5Dp<7`&Wyh%j(:WHztf[[P$
V9xp%2oAKK#,U- tf{.0?`Ym0]J\My+}a0c[YyH]#8Fk8md7AewgXH6wNhJ%#n5B1#M>uCFb31n0|Q"`ilrP3uvb"ExMH1)_ra/,Y}CR&9+i^~J{Pu
<9n$Mb4 9jI'wfe|Y5bzmo/MGg-IH~qY	,'/%f"g&{)X?m\ZOBJSTyIv3k[P52yfl,AK9i2j|x|dN5+bHf)8MN"a,U7[YbpjKN1B"nW1gL&Vl$C[i/Fr4Y*_R3]n(ZbYkSXr]!]%c!m[6@l^NJAgX;H_:#Z@|[1`y?jO!1`5{(;%wSV/ >oaS$1_m%<lU*JYKP82f/x(j9
_YjkxYN]S_(t
voGgx\WoFhj%xR6WKb~LW%(+:-VFMhrPWaRJ	\|E<E[v<FsjQ`$HK@w-u=I01{hDFUx)9zDn+5<U<5BwMOKzILcKc`C	zj*Ypn4L SWVMX:[Vu
ntP91W,rrG(wrBC&NNRpvgAk+C>NL&W:pvZ)y@+CWkK'[iYLDQByF:Bj{7s@-U#6C4(B?n	J
h$o&nLz<ICs9,S29u7qlj{io3cff43^7],Q
.OV3.y~k	"W^9p)wDn~l>623Hy0#H9kBwxXsgx6^ux8,FBAaLw-ZEcJ/zAl}<Dm>sgO:vvsbjUDbto$f6eG1m%d
+Jd'?v;NwM5h6-WVN%AK;4B4\!?mfA#vOceC4LCA99U^/-h@wQ2JLVj00Cp]9nRH@xPTpkSfflA=>wk"8=aKwe"%'l4IF4+KoQudo-z)lO>E%_PIH6Y)T$V!EP]lcDjYMfsp	BFQ=U?9TGRCw	sC>py01%f4@C&'R?9a!&,i8_56|XZR_x:d1W\	pAGA=
p=-*tJ3:*|BYL4j V1=bhKa$N+1~|-WI[qKIV&BfDI'`zI$W5Z^^`a$dnhq686pAImv$E|tU'IS5da{<[_8k]IC\}~9MAm=)PzM/[]Uz,<K~EX2L/7P`HQ[;Z_4+qD=d6GYH_)FFpmu*?Zebw[$$+zcke!O`IC"{!!mlYWU;wko*^i4N_;	r;c1L2648R2]AYsezH=qt1`0  wO
Us*ye"4i6_50-
< a_S,cvg>d8~o5R2]+l1jS$>yJYqYz&d}]MahUe.=.>~)}J)tQYFp>k\aE?]-2:Y]D<v^~:*}2@<}>T{;q5)[7UtPej=kw0bC29:@Cf& =$E~!s4ZyH+Ybv:n8/bq"lSF
;$h#<&! ~H>T_l}kt~yYX%0j}/@ 7Z&I2g@i:HF#PixD&a4iKo/,Y2r)Ch,fo]@FxP?&6N`ZsZE1,IP{G^d~\tNr^w5DM1%9?D7xEPK[u6D7i^gC+Q4I:D~\L}2^iw.GpJKE[H\y?~+'g;2[jl~[6s%r{L^iYawJz :JPpEF`@aOu"@Ce^[O&,'+kq_:BQr/C[*${$RuJ2Jh455Su.aHZ^k
6BgTPIQJR!>'hwk#:^v@DikPa^!^Zk0csEqi-C}8"'p&Kx/ tahx,
H1V5!SUnk0$6z)RCHffw7pb6wo"zrqA6l.IrT"#~SFf*.Cd&`*[5B=^ZGD};+'YGa4VN|KFsw~?F~p`T!>xAS9b4k)y(L5[[{py#>]G4 I4xP"N*y@]mohj+Kt"$guGz)q9hf^UyEp

cJomf<`Yd2M3e:#CY;Yq<m+&?;.~em8?bx2~.uX@$Yg*_TWk.%f3}7HrGu/DSF\s+vHD?lcQeY6Zwbzlr?>]#0APf&)PU!v^34W	=h!scI+O34~k:XLX.x*>EZ!TM9r7Xnl-gJqWi=:')HZ.	xm9YWxOWk}GD~n.eW-<r63Jj@1x8":,Nn);P9{e=7duTUrII(# 5E:|6d/c_.*$!A0>6V>}1*DQ?-f0e9$|?36},-'L'p%Ogl1BIKiGQ(c$LP|*xwQn6W|~9qQ?)O]RcY
/FIr?MCKnSmxy2/j6HU	ED4<^r%k}_R(i~M{{,/Yth\cCNAC)/6`<dWD:+:uy<`)qZV^!!0*itfS:n(>P1$z1d5N'-[Q>\.!bnmzp=/pH#qe{g-F>)h0d|Pv-_hRVXm4TAfI
l:T M#'S;mkN{smo5`xEekZg6JW{kXi<HL+PYl%-3/G9b5$UyA,ys0G3d#yZ<dhowIu#qd0wy+e1|NVka\IbyP\gbv>/^	:p%K2tku6y^v? TUjqqSwNXPh$ TwK']bW`mC0.~L@iyObmD3\~;<g<9EM	/-x\ZXm@AcmN<f(Ac`R-UhSGMA'W^=9`3B#KF7V{rK9pAm_-ypZ
 N08G3tQkPQV_xXZ}e2WU84M	XZN0LwM.-dYGYFxLL\wgGh js\.~sBmh/`'&PN[(F.2l.orh	@Fk|MUtXwfIBsIYy3t'c#|:U`zobzeVZ*[yA^A|$	N"@k8]H[l!@p{LGqgz*}q)BZ"'BMcM-xWTt7?V\J_hmA {$68:h7>@j?DVDz1s&.O?N125dF4#c TYR>j?&)+5HZqms2:.'&e8EBudQ08ttE
IVr[NKV_~q|w<4'08J}XC1~tf~gM!7}Lh ~/ER"h^dz)g&T0SF,yo^q{62!^2~\b.R\!-gp,A'pI!Mk#JIct`S+MU+(sma$7H>29(lx5<F}
Ab?F*0+c{J|7fo{ttU-w8p"z(t["#$?!mUq89f4^?:8`	REnSRY(O/sC&M5GV8*l3]krU+vt]t&[![9sP+n<Vkc=Iw3L[Hq/@XW`N%/y|FY,y;P{q/+)dg?
DI%S$sGyu<fyTvB	G-ue5s&2O/aRo#lZ]	UGC8	}$a*:tAp1t4t>`13Iq&8xy?cy<Mu-7VzU;qm4_XjNf0/_^7[:h=1zs-e/-LT(KS-QEof#*.=+R`diT`tBAV2uQdssQ'5|M<N<n4B"%m8pQ<Zu[Zt_mmR5S\XVT]g+fqT.(@>z]_pbUoC84CuH(K]	aF"uz<&vfOCBwaXd;ag+Cv&F:53:>o~p%N+E{:-=AQ/1*^F\kn2#H%e+zSu7]~x!D&pr4d:^JH{pws4k\$F>[tYo(={vM1w,B(QLqIH!	{:D_7
])f~I{(. Kb^/5-eM]"x_=vTeU(+M;T^%P&VLUPb0:XU	\{\zi51jl&xf^S_1j%oT[!CTchK(O{lI'HkK*m%ZwQdFPVQ,W"H]OuGzEDY5Lb\!=s89.fK`94oa8;lhirJMb-zo:mGReQgPhQwjD]@$==o)K-TDcBjN=6@r5Cw_3PWc77wD+E
d,R*pww\Q|Y(/Nj{}ck*N%;aS|l7#p'iAt]L0pCrbRh4&a~7<Nsal
j}Alf)j4bL;fs*u28p?m.pf	|q\TC3l],eTFn$Bx#^,gQ}.b$ $Eh;7!I`o#X[84<)%Ek%bY{[Z/~*!5OZFlR|:\|4kb~[{7h?&rUOiJVtk9Dep&zOsc\|2 5}$3apA=UmDo!(mQ{Kk	RJ5'^Z6pwLN4@.RcDM6).E6{O|m91y?%DWyqd'kY3l)A(z}fqo6ZL	)'j2
zGWkC(T{0_}N:0VFO#MkktHW\c8m<fl(S!R./uB4V{x9{o-Zx=RVUh:
]W})0&q.<B!(_a.}X:.fW~wHH+])\BA3Qqtz|ED"9$E~f#P\Vgr=!u`>Em P.13 %bB(2`U.O2A[Re">[@(,Jv_">b<#C8#J`
I-*iks.V&t0+o-hU"v^59xX,3X=n@p0{uZX3Bp^Blnqc[UNt@k.0iJcE}2O6/@ {xw?3Cv	J>uJe&mR"j.Uk}$#a`C:hJm>+.I"2:x}4#3n-"WJ[c	M&;|p1NH	yR#\xy/$*1XV4ba+&Sv[TLLrcb? )]<37=&c_\J {u0kV1XeMM}l09m&IT{
049xnYR;D<xQm1}fC*{0_F5#-cXVC:^Hpn.),/TmocUVA`E@kXD=2=9,#0t!pW:QypE\4Y%~v@.K[z ~7tu^gg38}e#yK#+T(8>5_	m'[\27b8ySN,e=:_	c|B7<%cJI_$WO*9m+V_Q e	U9Kb[gu=S
S@5z$-rRLM0/OI
r)S4-7T^	~q*!.,3'ELxy	p|~Fi!3g5Yil<+HML`J>C`\J#N/ts+cClUMv$Nbu I5#?BH_AY=Rnva@Th<6fd!'=-",jg0\DCs5(KrJfGZEeuO}=DEB^(oFnMY6X{0C)\|rTp3zFMP8bw~.}!	FhR[RY?FCS5qtv@dEqq_wpEHHvr]i7{zv?`	?`{)omWn})XGl(0(gt,%fj:uWm?2@{-u_GPNM}+lp=DNe.o)q$*\/4]5,y}@
m5UYE@N6kd(Tibw/x]Ff];DN{Ij	Zk0,@U3+{Y74()BwP-e`rU9#j=!TW9X dwp=]vZxq Y^^;zuLZOPF;qqALUS"|DC1!Nl'kLt~Ym<@m}kQ3?4hvmXN2H&w_PbQ=/oln=fU-{E(\*st^f 1k2`zrGS7H{A
WfxWK>I;ECUgfRT^#F.*/y,3ZsCz,QYrEu:Wn?!Uw8W_<@%Dl',c<n8i5;F!`4<PZQ8'+#/%vZZ`7(CV)kzOc}mFb;:M-|Ph,;>f3Gwe/"@N"?lP_zu7L8WmFJ"> 3BvTZ+W]~d*RpDMFX>
;LjXY-{^1M^+tIpGz}@inPe>xFA9x+v%t: (A*tYLF8wr~"flR/!#dV1iwl[`IRu'A%]'%iUwL-DJ'e?f!-EZ]IcKH/sN`n`:3E7U%<:x~J9krOhXU5,)yP['s`d`~g&ae>!oIHafj4
^1YZQ%3V&y7YbV8=f aNG`X"*MZ| tI\_M}PLcOoI`tdQGY'm`McW$/s^Wd==&c|AGzJ(6ti]yL4\fb#hwYTCWrA?{qFzqN^	n>r|t+k#O\m9BXk}'zIN0	-_Y 8n2<8@K%(lZMi_97G:W,usuWVoOYx$bDW\Jq_>Bsa> Te TZ:5$K4gStT+gWx_l#zW>Ls~bid)iewU^B@Y"g6T=TU_"u5<YOl?f`d@|I74~uL6=[\2:2sY[|UzG/J.)	2c:\$(YPTK.36Bn7N1d3nN[C&Q:S5/Q7zy&]LWpbK-{l`ivLaf'61}MvtFieJY|yZHYEJ1ha{yfG=]tMwTQ590UC:\^+4<\kuv1	w	$PyXVPA@Nsyky?Emndf*E@BMH:79ydN9:Rhj^raT-y-Yy:s6:CR.OJ#f')5q-`e$/WwQFU,Hw=7GJ,WcU2qa*@u;t?1B~YfE$@,xcoD8w&h`G&M=h>p!	^nyb@<DXY^)iPQ%rE*j%>&Q2@0Hm6@L~. M@/sJ
PGk=COYrOx|9T.QIavH|.[6e*Tyx;@$Gb&4V,s;L=X@0oYHz?K#mJDYv](KB:D4`J#i_ <B4LBPh*Y>!q3G,3>J@S1Iz}jXl
N{O|{1R^;ujA%`l3l>Wd[l(G'G{(-P|zut)hTDe#AnUC}sTqm `8	@^ibm;h@1ghc_kA85B;QoJ*G,Y7xtX8xj|m>vQpFS(_=t}r;X|u?"weOkG*zE5zp/-{|*`i]d}:&5b,Z4$$9V%J'NU"#G:z<J8q+("a0K:_7@Uzn?kS5(41q9/yOY`wPn`B^c{lZEC7#OT=fR~HD;PA_XmSDh#5+1~dEE(zN2P#'knM_&z*96XReCV0DjXPBA-A5pQ5R25N/J/X
&}}xX/),v|gI<ti+@Wms?k@Ph<DdYSVSZUuXw[t+}B)C|ljZH]n.-G]:"X??i(!P(kZ5G0qD1],*:Hpdb-6G!o%em9hUjjZ0jxICS[,y8'+r<n5h]#6.7AH&vFB=s,ym*<hU|f+zTn94.^bh
V{BAdZXCCqd"pU. Ti;.!vzsnY=I2`8HFbQrClS#pt$s[szV~^[l'*iL-;>=i!H^GEpvqV>~lQ0_b7e8e:i[96INCx#I+m%}YTm	1y82my*}Ka!z}'E1 ODv`,`za#TeN10G1$J/RX Y%,/-T+s;?EfYEb/N`I9xu4Hi?P{Hh'qCZm5W^l5jD1%B9kKx{?3:r#F|o*lD|3w0YSAbW .5#p|9oT~Zx .o`KJS'_b~UVHg%yHp+O8bWMpl-%@[~w#V3}BCC!UiYJ!|Q3FHM6sEed;.63`@I"kc,x<^o~6&h}<2QcW"EO}3LyhO]\LGj]72<,2!WWMAc]-=.r0./Vw7_I\4ZS7P?K9m6B|`]qY8.*w]"rf5+&K}D2bOu<AuKxVnPeCCFV)&}{3&#cW^Y{83M7]~}_<
$3}B[x^ @pe85o12FIu,lA~;"afOq{iJ	jEw5}Tgsz:sbI{1S*),uwAKgxG(6a	@1]T.eFZy5e3ozcESoIM"u[i%J9N4(7*@9IxAP}=( 6@-Ap!im=p(huw~'wCEUYk6>XT(6RDu^kU fvh7!wJ"c0!@>cCe=k+A}#be^"H7@NNHC6f!&fUDd,=$h@2Pml1;wve"6'Y~vO,7qm0!B1"q_BenQ&A@o?srp[t`Lu>(yHrm=x^`j+9j\my)n^{kpje^d0Kc%+Qj:DW4&U0={*:f,t''>Nxrx-!GU!?|&3h]/Hs?j`3dH|S#+[[,l}mu=Z6`s(k\b#+}~IBxC?uH$Vxd5$QN9A3qm>.W[
%lmZWu`9od'!/Io{<)v@hVF@?O-MzYG=r!<18D)X;Ad^Mo.!W$]g"Dka:cqCsR~;3@Cn`$sQlcnAi08+MJ9UB	4[k#ZzCZGF>O\hvBP<Epk6a&n~xuntw6CmZ$hFh?^>aX	h9As_'+kcOMA=}Svpu9RrtU};u=7vsSFQVL`gbPhO'Ak~k "4pi^m>`EUn+j rSy\e<Uc[-7<vDY(/Tll`sm^i
B<h1"`/
WVp.*$WTNPQ"14Gg
\&0)0K{K.LyD*CCVt5v<;kC0h@6$^:p6(l2(?v-H(K[`31&XL4)n}!lPw+#=\7{y!j|W6.Af0r|5N}`Onm"fR+J3@Y Jf6w&U*	LYI7	OOW%lsnrX?Gj~:87/NL7ne
1Z&gHtar'-`j.3Jk}E:_2W\>@Q'/-H5YH!ahUp:r_QlYLaNiP#ukeV}ZdAG>q<tQ:B%(<\&>&	Mcm?v S_PXu!P)iJFM{OON=MERpTYo]z&G=zNJ9UfKP.~VZ9:h2wO*tv]:OB!/@F,p~j0Wd&9es,	fimRS@?9'TYwH]8iJ 2.BJ'19<|A)Uc2,@>r&jf?((9(GF?>j3-Ijwvg:^@K$n7w*:(]=2M^ic 7FB X9}$3;/=,L.mK"H%=,hnh
9-9-jMpKdmh0k!Kx*Z*TQP."TX(cG8DvAEkQ.X!rrW?aq$O6&ZVy%)HOh%b,`i m9%	=A,A;Njy93B1KlvTt6E}+}[tL7@@PfikRzK<VUef|qK 6?2af4^'GGm\i
yuJy,3?)zif^nEkgxRp{u<bB	U,3%'EC9O&2_&4Pca'm$g4"=}n^U\^'/D{TQD>)/K0:]6u/>d o"2<J^`w-2r{QX|=7\c7(|[[XWo!R:%VQ:):/At3{gv#bS=.Lp.((c0;1h7LW*qsn
=y=dR9tH"rqH,n[qM<7x^(<t&{E1dRWx,qu5.~&)ltB<1AP7``g
w3$ob|wUkc<C#xx8{wZ'AP]2+a}]l{0qT:M21ljVn!Sgn,hja(49zj|f azd6P<eWb]^|2"mXC-v	wO$U]rz[E'n<|lyUCOK*5gVQ&Kz@;M_,oO_@+:1AH)NMX9j7b&A.Ymuxl8<m4
]|y#,^4mq9SvZ!&3DxD95(d{CI)gl}O]!\v&5frtHIU5tY*]vq*T|).A-mP,%G{,ZezJ5X^UY1[CBj
P;S=Kyn#(S9BW\
{u>M	Pm*O
aZ`fA3[@e<fUJqV?WW8f+b>pYd}b71VKg'r*VLz}pX&40P"tuM|[mL[s@	F	AV@	d_5"*Ip=#0TxQ}o.eNa1Q	!4(/
^U2Wk1	dFD!)ujEC:{0mjRiZ&kpo3U'@-r^9ocaM'Ls2y)~e~pY'tn<E0@e|OyX
8!Rm+m0]}>$CJ<{n)fEG?c%_P"_AjD@VUYQ[(%RAIHMl+c`(YX%A.v
,H0vO^Dj:]#===81St209%*JNAioenD^_M8FOnXM]d (SM;ogmy7S
Wd_
v6|=ZkD!=Cg6gm?_`/9yVzNNR2lts?Pj=l]Yr]EjL`>dRvZo64lR^:"3RnFPe*BDS }Q]IOEN7x.eKD"3S&*>l;|O1B,2xHS
_Q}R7-]2m-*aM%`]}A_}KMVok8}OM{R-A_N;H(,/J@c\NLw$>JA+`\@etSm2~gE"*dW*6%v)b";GgwY3h#=
8/[(~.F2FMUkD(922X%\urI!f;"cAxt1/|~D}mTi+0ciJUQ# 95&7,<6bXSq!+$MTm}o&*^#U3LtENtiiaXWoz&YN&hZc9<^/k}K9-LwpRpw^*M@(1Fyu)Jb5^svDuC8lu49fH:8cMfzJ*IEfxc4nhbVt
^Qfk5`I"~s&+Z-$)p0%A!e	Rxed,k_Jt9aZsmz2^1[~y@@z~_-h;M,GZK
Z9/CY-*clthPu3Y3dO4o#3}{q''3o*}tN*%{B<wfH~Bf$VZ_At/VG))dWHx`&krU_J}"U70"6	*DJ|e/@lRFpur`rLIp;~`aAO61'7['Q!^TT~tlU0":e2+>O;%`C!}%
91UJ/4.$,][C(heao[kL*)esBidY]{[%*UTbkhAyUa2U[*h)u6(!&f#:Q6%5])&c}wfnpRng=Z[NU@/RMBp3cI98v+N\r5~{gD10(oG=Ivz>KER&D2"a:[(@TBCkMq`HcrnkPA@AO?6gD:DX&%J+E7ACg~;s[1Zg/#aJlYr'zUdBtKE];9FC7'gZ5?*D8izPq6m3;Sh?'rd ~rw11
	D!4p Pv YA,ypj>y4enm%+i
/F3B
eKY	xRQ0JI=;9L3>X9:oOaw}s0E`m}nS(yTg.ua=Jg60UX)^jau0<b$Y.`HIYxX$R/vX*2
iW-${hpq61*Y4wXcXR1F-+m
f^(^&$<9H`;_3}@xSl9eE%si_XZ'_+3uQ?PHeRGCkotY;s"5om?KEmfSu]zn1dw9K&b3KQ5@~|Tf
P525'4\X!kl^5I>$zz@[%#QlY4#[A;<cM&G(_ChCf$n$oAU
,x('8#40Aa%-VknAnZ$O-f]F0)##B*jK9e	:tq:_YTT^^|F[s{QL4Xu/1"*AXyfR nz/NSP,e&Obo9;SfDwD^xwA&S\QWiUu>3Caaln)],{%N/N/qSwP>*X\gAbbs2]CmRzBC'VuK]3g
^HP_p1PTR8Z}Q9mm6RB"B/L:+jpcRmoFbt i%"G1wk2$D3C	|j'U~l;xe_!,,WMRD66/0)cM4"be"^K/*pAZyodbmsxca0L:T=Lq$#zjXw'ay8DL1z}@/?E-y(o4v@tmVBNQOp\1c7*@.?kD|tW,[2.F;jz#,dw7m&QiZN4b]/X|y
RI/W0RCVhOl<URt4*n4Lh+YHOKx5A=)%cXzNMgd%^94t)6(9g3&AlEe{Lk:BT,3mchtiAG?Qv2-GvZYuz3+UAH1n+eHVX}+UgX(M]m)i
9I:&~lmAW#zO;uEQLHgG@*/9W.^l.Kaw&'*RKa7u0b ^@P%>x93@v:%1/&vw?4T{['()
	P!U/!yo/wo~bcW(]-w~f6i[<Dkrt4,""0`|wCHhbRgL#RLv'V_XFg~6GWHssn'y@EJ>BJ4c_W(x4=]sz%qjdQX<SHdRFN]|?\s!R`+ee(Bk/vn?J&Y[LR`tE)RmuA$a=7Sd]~.<U\bd1c"KRdd3+UlU#Pg_P7{()6WSfaFo1)-3.afX>t{eeffu
_<,ebgY2!TC\:1yeOq2*F[y1ec`?-}Ps!g!ezOK:. =^pEEf%OsI	MhCc-iGLV.*k5E5~G,b&kL:#gwuUZS:{p5.h1`8v<
GJP-v(_--
(o60P;ciLv.Z5W3u/xL&O5ehye[Ja
P"ps8?HyA)RFdTx]NRzOg3jsgU$gn@b
*pBy3Uj1QOC(`j],>c?vM|U^v_\ESQSqB>xfSsm5;AfmRn;g[!hDyjx)bTQe,xAz/`4e9bgu,Xoh4R}PNMePYGw5S.|{88_"i0KpXid<n8#7Rdj^W6:NT}PLLm67*LRdrP6fP2.ZVOM?Q_UF7>6 [n~pN:Vl=D3}i0VEMCmfHlWAzNo6@_.:1P*'\\#%jLISDR,_kHE0>P.5R_D,b|='Ox3)03]|^Pz$HJFLnb E\P$Q!JA)HDXr>#u~%"&ZLGqiz+R3#]?yI]6Z^=6:caV:pNUeoA!R[[;PIvYR/0&.CF%Ir'\':Ge'zfi(ha&G~]-WK`aA6ghPQ052gy&YT<t"	Y8$!L
.=ydfPC|-RG	ecd-shS2oSk0><'"Z481AhC(ap8F/PyDis{c'%m$f=@9O27{	@1)#_k:~ts@Yj.`XlLRQpHXS%8i}+:X:jXFDczQ/i5o,VNLx8+^Mp"?/m	

A+	Jc'H	tP`hFswqKikeT$j3'.9@OhRb.'C&uY
p#<.qDFXoI<-N?eGG#PEK])P]*TxV_]_.1~r4&g+` }b2 3j#s;Ts~v[G-$<,^L&uarJH0	-		
y^>*.F2ZO8OogTh(]$je=mwUDQ*edq83
99)]VM`\LL^:R(sD&r3l98SL_G|K*dYs9{#ya"a
U",SMOQSKh;:RAl@c^U
xxW]0&'^Ug:vdi@@fr@H,kpg&?u(=T-*\|L	*}cGHcqC_X]RqP'q:Q,RC@Cq:<_l"Vp4xms!.:MfjZ*Wr,xK$es!yea@I.Dh-XB!dx<$/S{j`TF#]`(AR~ry6(krQrYXj67y-~Ro&,YhpCWj0 X	^g!Do/% z01Wmzx}zNV>;
%L)n;mg)_i{q ](X&E9zEj+X;VY;x8E=S 7k'nrj.{NA$3W"&f@m*=pDU:[FOZ-)g\C #fsO0_(#q6:3]9t)f(Z;?-5Q4Kj-RF}k)PoRnM}]u+mwV]steR=["UmkQ;Th@%5=JfyB7{7'hJO,JodA^t=Aa-d[T@3Y>!fFu>29|@6E\%4~fMV$jp`sA+T,VEQ
YS5!
m\zjR;AWa";}C/w27F1Bks)w#=}@@A?[!d}ZDUffQ79&Y{r!-L:ekoz( >E'?D`M%r" a3y,(8.OQjx[Xv+1y=+_y\I5(qijNlhe@4}PPv|F53kO51'wKmvky$eetT0qIU.2k.K'_dG$pWBXiX7X
K,XGWF,yY:Y.@s<b9gX^J/}iZQ~S}E"k9xH1l'Z.g~zUQa0-[)0}ZPNDJYS5$'CV@="L?S%>cIYcq3#;4q$5$vYTii2wHg
;t}i\	%9Vzc"oz4-zan`NmVH-Nx='5WH*kosA&"47DoqT;Dj,Lu6U;Sn(/UNETbS.~_hf<~]&cJ>ch'."GKfuKi,!e8RsJ3wZ0rd&lKjZ
S[7znU*0aH=M\G([:':Gk@
g(i\Y
y*oxfP0X`!}hy+kRCenM{2!]4yv^2n:Pj7LC/(ENksRI@>Q+Tp_(_J1sh	)Dm7UXc>=->f)p~DI/48J>hwoJ	3.bv`!{0>Z~HxmKz[VdAB42#~X*4<	OEyG+cHdOXd)7$o& b(Bi-8VZ)v4EkHOK2;P:O@q0UiZ P)1/k1U\vAgwivHIJsX~POFU0Z?#{lZ'pf5$bL:|vX$RJ,v\s-Z& 5c,r;WmL1Q11/?foEU!.[(co{qg_6#2/Ko$}}{:QJ'H/j8`:<?Js9ii74Qdl:&,b@z"(&{^R6z=`'"U$O8y}Q4A' FHiuMb)gw95":7G(P(bZdCDV2E~`F[nFgg#Aa] -gAf8YZn+tZ&jV6e):w~=jn`NDLl+v}#fQ~wKwCCUZ`rNMn@8o;}}Kh0M?37
e	J281;^=&E
`+'=${	Uhq('8-:hbL{X3R<Z5M[;505<zE][c]z[?T*?Lw[uGyByRv)5\dUTY\9@W?fvzK"`TA`_|f+'T#z-IG`EIqg5bV:
H}ot^[VPg<vs2!>dkAupv]M(:ZmH
*s%6 Q(2} +D4Up(Uy
qO'`l$t%k+h*S_Lt{UAEx
8~IY=doW1~xpM;CQ%3Otu7)	/4eq6S~d|6synu7PVVy,XqG8
kX	|5a[<vV'$))<.LO]^P
u?ZTOA@xJCv_\&~J$'tLa*#HELOb##H$1\
9R{nTpSRbuJ	4{d
o`7ga3YipN=DYh*e8rEA?b' 7jAF5&/s) >&OM\bCH[!$2Q0iR}Ty@
[gn\?l| 7 PK 1 G}dHp6` $@b=y-IFiwB0t"v696w[h}oU@Y0vS%B/*@|13;H-,q?ZSm8~3GuqEj2J
6p^F(9N)6)M](i:`m"
km]B`2LsoPHTt5VKR*ax;>Mjn`{7:@#AWHJm{je|lhrODJP.9@Vk*&KMo`Ph6&}-zUP\)1Dg*rp=>bii2wyxN`BgS(TzwFOR6n_3+)4
g}|G^kp{OF];@[E]e!|;v[qjT	r]Vvh/@"|f_saB7 +K+Xk~rqZuC()|l,$S!-zf^?&Tf!3+Bcw2$9*'lg!=M	eOBI>tPll)`za:ItZ/aTQsQf}y*).%%|3nR+>}?l`piXtnu++vm_!JK+/H>;+aGQ#
?U,d9C>"bY5q7L%4(J(JzZMXm[
5~:"wkLl{QVmxPr;JtatT)u>H{&\F<0%uS%}~1_!>[	c,X(1-%zFZ/~(#kkd|++eR/TvCFf)'aiU@0<+[L,o|N7zJI&8ktLPx+m.=vo."MJr-^o}CJI7IsC=0=Ko6vZXR%YyT,+Erw`>W,[**#{n;+A>:sgrWQ )i:(TO>FK^+\
5@#f8sl-Io-SoAYTPUpQAm\tYX,j)l:J[a"`/\kFZD>#|HOx\iGGOsm@RNX_k:5_rs_|@Vb@=;#{CqwF!U]t,:=$wR^c'T+9Z1fH7O]Ha6f1.]BtX&FZWGWb-ISwr{W_F&$Z`?|y]3yg[w6q}NBYu	:"k{*z[/]uf%\ZK3Sj
g5.>XZ	SOBnsH!Uce_`.|-|OV;oqxb&sw8K8<EBbpcj5*A`7usx$rG9aa&QF}J-Ue,: !lRHTNr2b:dWomftFM)
\}<Vrm;hJnQA~Shv!j0>7Fz>Zm%B1gBnYw{FaO.YJN	.td:TW@3Bov:p?J>H4
v{kd'S\>@Tfgl98f>j-9F>Sw}V+CaNST@%\<goi"*-bqkw24K)$\N= V78$~WH/s16%]hgbX&=bWpt[)Q29{X]*Pg2H\=zfc9b/;,H"g9x6hm@]J+F oDoSHdgTr52w/F;Ig53't]9fvq9+K|9kcNFo%qEj
BG*GfSs;f12avw.qRt]a3R)ljJmNJ6d(^!	i1.:<(:`RLL1Fz9;T1 h4]J5>xmlt>4AxK'XS~0C&)up700wlf4%/#@rg	l@vgm/&COQO~BPRA~TL>pL+C>elZ"W/yc:1CD>Jwg}_P,Plu4O0e-~7IQrW=CAbN >uU+\dtb]wD52#O*>3e~JH/=Vcj	&Inj|\APg?_BcDSv;j5-Y\y#Wl(!]]bq+Z{x[k+$D
5wRI82xu6*GV|MC;!W,UIyHZTqVHgyr(%ydtC~S4a\hR0YD5SZP"|lOK^&wHm:S#CRY{OKH&8-d3mw;mXa]}P9l}.0HwHAc'V
RF[@8bF]qC/{dKDnRb>`7#q3*aHWqT>\b`wJqL`zg0XD|f<GJ4M tSx/zng3juB3`^Ze	sOui^R] g|!#![vLd0;r:K|y,uOgro0k1e[uPZy]XSF@1O~:=Mkb5L@a+'q}:;JL>lx(g3Lo[rn:>yA\:YOjjM.QOJMQE]NJJ^}P0^79Lgm38Aw!^6WwiGpv-%f74e.\Xtuv*.^pY;N(IebP|,@h+L',L[5b?GI>-[1{z$@Ou!D[I
TtiPBxJ[b>e'kSm{zo_#ri	~)|#oC5c_nM%L[Kq^`lwVMb8o4C{2hBawZzkOPi*E)KuUh@n)BW*<Sb;QLAH"Ww8"%."Gvl1-th]A&d0I$Y&t)6G-&J<oa)`*9D$v{]$.$89xXlv?]U=:#+r=@dD&"\>lSP5gvGD/U/V`Yp<3}~	K,=\8A,(U@/FJD`:5F]emu_XPxQ_9zkR/-o3pnBwMw_1vX6O?yh!/Y%$c*u>A{H]G.&I_"
^jbP/rV^"P|40c5+uz6s$J:Q(,rYVwz!L)xR2Qkb`|0Kx/[ouO|N1O|^<@e47F85kI@a/)rO<q;}Jz,]hu@3luon9%j7/VdGUs,"LFg?nAO78g4w=%,d 62{)DLSq'}=:Mv;U%7Ula,A'X]d!($JZ1rae^S^
59l0:x0<PoS/=s()O)Ln]WYdP>,K 3}^dKGP!_'xc6-0R'[a~@C!E\Z6@*hqa;y/ff>CB8<WFqnF*7nQ0}2+9hIJ]u`6O6pDXPxxe>H^+82{)@GQyGyzv8u=iJg,=[_u(oGFhbOXhl_XJ>kslJZ=|`Q>T5lo+*9cpK#'^<JK[YZ,aSdN3fB#W1"jXb=A)_oby0s7cT4NVVfi8\	IbTK#k3D+(4!BH%ArTu6^a{1t&pzXK(au,/l"Sn?R6dk./ A#V,%-o},jwdced7l?=_<`qKo)FX7d*Bi&B_/wa ?21#	(IBY_<v{;<MX\0&9VZR\U%>IaRpLY[+eCnA/kUPJa0ahAp(piNrX'&s*:*406xoR!aJd#\G:?H<1:fW][&w{kbeAe<h:u.PD+SaRrqg\r-/>D[6M):de20\cx">T|9W0|-x~s#nt&^QG	c[#tj}4Cmc}Ad<Pji`VYliU?Y}uk9L	nr?(	L|p.	q\u{\LEVE{u*[}!B%c<%4^]WV;Q]Z:B])kOrDayo2mn`<IX4h:.y+@i8[S|u#-<\uEtiDbF"):$cjv?j.IhTEW	L<smd>H|2>V9o7w`Z7IOntR-,XH8G!ms_}Sm]nwvC?1d7X-\Eo:.1KLa$u5/U$	e$cf"zoGCuRz)|s
I({nT2HF&$u8
c.y%oAg|UJSrskhii3I"cONAb<SwN*4KS@Ic/Dmp:ZRRSbF!aw9+5ywc=aRcEgWY\e9-7x+f4m%q"0#J{9GU*s]rnrp-Lc+yz,5'[D^5j2=h=:&ZL1q.']A[25>Oq,Cia^n>18up,v3p:~i>	PkB"I6*m2,L:+DNCz`mPva%4>?_&+/Q+b0u^KN{x5f)91u_tNcSm=h}Z'DXx\_z_@n^ |n/D[F2Kc5A5
1!h10a);5eO,t.2HEcjV7_N=UKx&tFzZ:CH$q$=L9k.R5	k:"K$; 0#.S @/G*IJUE!2De0Y}S9\'3Flm>7w[Z+5UV)K0RNE+VYPvhF}s;h_kXpdKEQVQ!_FDD
l+)5r&+1^"(On{Z6$>Z>[lRg[(v(4:-^v^{yL]LQI"'SJ5x?Y:rKF|;!Xy4Kr%>8#K4%:[tAC\w(^=K5JdeG%>U>g1Je=n_  %%t &J]3{enwQVwu43O[95Wk/7A0~#=tCq6&0|^dCw"*#`^Y?e!TXn^++%t_?5+lxWPBadTCZv@R/TLv+%a<mP\fHRu=[J>A'_Nq&<Oz]RYj|aZW7z R]q6V/N46\FW(\V6T0&,2-s#aN<+hs`PhaM\KnNR*K-r[x8Usi2`)3GouPYqs#w$(7Lf@A,^{K-(#!C$8Y&r{Gw>(96AQgpL2:]N/$kV3/"FdSi.fY]/5(:I<Qs>EA\wlqNMiKxQZ:O0LK\V
r=&M_]`[o
)JJ6R8,MWa(P:M4U:^Y<JZdrFkYEHE!zjje{9On`ggCQDsG7!Q6aJP($|T1o@`)u1**_Z1Ary:LZj\H~QnrBS=uX&{e.QW0q D27vwdnsKu@1t\$hRelBm%p\WOP'!?bxWZ_WNn_RExl6KhO2=q)FYfgk,4-v&z;y^+y6I?i>'aC]y4)Oewu<KHv}gDfX&"BbWnb#[	ZWohLFw_a>>:z4p$8`<[s$5d,2Gi#H*\:X?.2b$I-}5sAd&3+,<Eq(N
jA#1IzPIzeH!T0C}LnF>	rn
'hW|"Pjz\9CkT9W>1/]"LpNZ9`fiXOV$$
0#-@l` blkY	^24f0/Ga-%jP @h<cWqBOZ6))0]/Nf:^rb\QVuR:i#]>4Li2n1}}Ed?j=/~bq5mC`l<<X?"&lzXfYZ{B*8!]nZ&^bkRF*F.Ri5GO_w;Un]k05vD1.MjKHrmAw	F:dHO=HK4nMx^%os;0pq2:WV:&o0"_L|~8DJi~a@:\\;3<OsK80(On2
XbW1q3$_%US>^RG>-%4zQqqJZ'"ni	}h4aL<?6/q2B<e	NAv{"q
]^KG8'OdHMDhv8b2FmtWdMMDEu".C_v%j.p;e,M%]s3
 p>'	/*ps
tT74Deyt\<-iO/xzLP7PP!Ri%xvW:uPoc7a*!~1bcz_I;9]YFK4`!`Lx$RKk)#9=e7B&}~nW	i|,KjA{t1
RdQ5&ex9ESHYj>p+ BLVeH8PRxM$pt3EO6~P/tt!A[IO]'^9y&Pe%}l6{khJfZ~/UqK|h[.T0,q"wc<~P;j.lX!~|]4gkG~h2P{U{>E82PF67uk'P^bl|#q[Y6p(d:q X+5ybPZN:1g=Gn0Ex'+:KiCKp|en-7'o/;Iq@+U9%db}A1iX7E`H;QtyA^nS(%\KS;&%}5eML&Hf3c.<%T>os-|p2KeGD-!!_bRW/Q2bH3L2~O`#lHzIj%d\_i'^.j(:qZ
mu}'h|6Tj<MylR-NvMdb07yX$DG'xTM."!{eFA>l6%SFPJoo[oW@\\eB*
=n@)d38Ze9{78l5G1>}3*i~*YOkSg-2FO^7[C3PZj8Pc0@qt~Un>KJ.7^@!EeQ/Qp5t6q\D WX^&G?9d.\6YvNKU-("W/DM>yNJ}@4L^-nyt"Ws]me_S#~lSQ%7zLEL#MDEU`zMvB\ [>CzwP8Nk2}ONPQ`*poP$K{K".Wn+s[5oEa_)Jq'%-%>>j}& gx1pp"6\v`<`\tD&f7.#?uz^b8b5y6l[dN,{on>74yic_JA%F}ZO6-M@98%/7dj9}-  n,hm#P09H(+Fvi>24#FAA[ks sQ8?,9^e(CwR"%bg"%6v|Z/7%Sz$n=tEzN`':0T2!(as\AxG*,D3"#KZX4=4XM1E6r/V-6H9$1{W4R>%Pd>`#m	m,[^; 83fIGc-BMM/l(iuw.:Y+A/pOCK&WhCs<3@:7#X^cK{CMY07SaXJlQ g!'Ui&XX(#?+t<$<!ju|	MLU>Yuy{\v@2o
f&67Qu_W0xhYYi<DB)7A.i=2 aY1le|%v?4#iae3FK"ntWf7/Fi[{n7M:
a-ULq\R:v#z+96r={Xnjrt,/x0w}lmZmlE/|Sy;8nZi_O6j_/.D>*{r}/<s4nuePQFw\4D$k/~e
FJ@j!3OvsxYbaW |RmWvt%xgmoLbY	zGSR$~0	\$@\.4B91&;yKN>`c6@N'CLK[l$#Xs|7Khn:\K 
C +D{?X?Bqhx|TAmz!FB#&
|{9~NsgGR6=k"@8Cy{ LjT]$%BI%5QKStR#9@be(4?n[vM@D&la-jHZ5t*DN)}PUo|*g_K,?o	tM HUwBwM?Y	RmPZQx7C!~'iv{c@Y(k[SJ8g*h=,ZukNb]c{IYa2t7|;_*8D$]HQx[},*
*%-oi,7#:.,PQ7y_AjI&dSBjgd:s{`TNf^HKH|Winy2O*oxq'f 4OkQtj|w.<m`rY
okhH]SlQkgA@p8!{R)ev0z)'c>6Z ,vH3g%Q'#6C"ja8D{(>&-DO~v8]8(<:>cIrSij:X /M&["&w[CS!0)=;-g@4?,+'fv~wKX8 PAA.04)CwLKx'Coj~" 'Ea00znSvViqp	(g|nn&EeR:opeVl$M3
kT#c7C!XE,i~TrJ[@D_.-4Z|bO$S%2"Uf)=rV^&Wn0UsO=E${Nr	(D;S
#L{!-HC~vpI5@`IDwEW"<NN^p}Cq[nv^c4/G^:WL-sMgMxh^\M}z>gzvW^s"8jOa9@umH?/k-.s&4N0_U'\VNnRKw2szle<E'Cbe{Fsf[]u'0:>"leHUli/s"1W^;G"$*&Dk]U8c*9?2C^u=
Bp4%+B0N#40DHHj8M0mm8EDOxDwtKnwA'2"_J<K^$R,,B7 O'Bc`}I&`i}Q'5QS>}Ny$}"oz?`g&R+Dg}wX?$}e\M*g1UkrJ[Ad))A\zEA#z'03g}eR4C,;` b@y{q`1js`?e{&ab!N)QC|8ZEiJ:3aF}"{VF:.krz=R,>T;N.
g9'g$"f5Zn$NGW28FW^1:fNW/Lxw*}F9gUn9Sb_o2b}7hH<p*MhnJ,	2!'N3Elvh^=eZ`'2h~zpi?E=J3!uBn'Oh0 m.0J	=vzWyz%c{pXxT	&-Q2G.K72q8#'L	jZRSSCA3PCyVx,Hb-/w&Gds{p,	Q1(G2ManF~hg>K+p~/	n|LK^(/E1[Z6'%%\&cdnCH2klr3(;q(ue.p6z%oU_]VkUfBVx[	^w9`4vYn+F?~Z_E}l0}\wXD;MuX	&}BPnM)}#J#$VOi)KSB&"%j 
."r',NihOAF|tQC<)Tk?1-y3x|}~!2Q$
qZrgL<h]OcX(s{8=+e\(8K2MWd9$dAU)C6q~X=S..GubsnY4PG9)FLu;!a4!]h46`c["n,3W!<f:_{g2!]beQyO}s-fS0]~#7D<ma#Vm)`>^W
\~Fux	<jHNJEK(_z.(Rz."Q `t5w0Q4r}l%zVNF1Rng&AqBT-o@%m_\	^%sC1,!^FKfR13Mq_CalB)F81DmnOVR&Guhu,9>7E^BH`$*mV||lqbC#^q:&6p2"j2gu^";y?8 [>I-.wg
X{]E2$	#&/7vUjJ*g	Qhf0X7B0o2JSp;rC]#pPWb&$),i9ma-	\Kq6%=8[F,gGUW9aYW"{s aT;,%hL%w)v})/0Y-xn.HS6rDup6j$C":0G=w=
FXH/EzqA)A^<@aR%sM8F(K[vT<`]Bj%4H}o;`%$uk)96r/$XYKlJ-b3t"sr7-EnP[/MK-Z/B>IKAAT+u~V!n*_zoTE`|JO8f3#St 7Rjg8T0`v>Hx-c{]Ar1xb|8AGkay^xLlUe(53%)/rWdmf&1DYe9GFx0"F[[CAg-xG75elLU\H1b[3RR<[(x:)^.qai1~=-+Mivc+URHyOePO~GBdU6%^`SgYIg_|8|PTp%MQOjzT..:0?2LkK$rqRv:$2sp~+S6no&>GXPyg#br+9N[v&`j}BB|Ma^ &%4	5vCK}qE(NhXb|l:-oxF:|?/D!j[mgko]YZ@}{^-q(,O~`}0SJ]Kn!CbE`s>!	Xd>^GfJ=Fy<j>L-Koe-y,p#}qe1*p"=pxc@[m.R\_Kq	[j:TUF+?j]#"-<&:0(	H_RkKhF+`SA	=/"xE]@;yrf[+BXT=~UvO*g
5C/C0?W-;<[+H	fc5Su7GrD'z&Y7X6n(NK*FOrr3lWPj}9 E,&gS>=Yls~&XmQUn$"M`$:uqd_}>eO,k_"6:.JJ(11qhAFwEeYjzaypFL(&zXh7:B@-iW}wO8kjaZ-U>ta]u}l#ZP>+T3/22'epyJn6= ?cw"<{c=!yg"yh	|'0RdtA*8R#Y"I]I,cj/{'Sj9cm/&:&wMT_FI=U(q},{z#jMz04-aUG57@@\Kp>@(2imQ6p.[yN I 2p;~q\Mq"LX^>1nu:	/jAQ5	C:ewI`M?GA_	k8.A#N	LMK"Fl[D%nxNV#+%/"$V91"N)F~Ioo:2iQpBQOXsqy7ZN(UW5SIe?re$@v:NQiy|SE`kQJFyK^ntypE$$FE]y.j#%Nw[mlc=jOk(I,*tU]w_"!jb<chUqVe3LJJ*hPk,p?\#a<@vtz:v'Bbu(4c(S:816-Ne0fa^$\%v
v`tPN#U1]^s Q(^B9~TsBn{{W)tW
^Ov*T)]m7-X" yT]Q5}*mS)D8/0,Crx5pPHotn&Hx jw5e-o*InU"	vB~YY1C#( =Us"2+gb\$nR^Dbf,)Sh>75EW<n{l\Z>;PS&	-uF1Q-rX?Po7#:0,t!%j~J]'o>=~m#7e+jFf.Mnm8z52c1QkU{m~?8|]D0.pX]
H`{L<ETO4lo	w,@f.M/,g9*P/D	(0A<]lnXN: 9;Z -|^gv0<(yHb(j'*+Lt%pmW`YQ/O:O1+P >2Di
2+,X,Dv<up3 k
|7.h[
B@4<\'2_LNpN
+6BKZ2d$%
Sc|iZTwwuvv<CR P}[K)}n5jUa$WQBB A,3|[k~.%Mv6F9hVJpa`4XVd2dsieqF;2d"gsRH	facAdL"? zBtS%0/_@J-cfSN^MSEqvM=f#G.q9~#5a4tGCP_K7B
7ovQE9#2&8;E87f<eU?ct!0>0=0Sls@!\u0j.QB%;6$s>xr(r% Nmlqsa(1;9"kX38;^#RI +I
)U[e=8\G%:KEZ{9i9-I+M{s&9r3!
wxf}.</v?5EwTm'aw0LY@.?P9qDR"J$U
h\SrUT?3j[TW8&.I!!)0s*<[x\+]i3C>n;.Xl!jy}iRSB<D!w|@$Sz0tEN.{cQ	'%iK^V\$SmoTkTjw1sJuDA4%eW3fp:8,]Jpx_"{S=B<4 j5	LqOXK^}&:4N0tixnD[ECM`,5)}2ghG{scR4;wSi?9v]Z0?U&#%E@IG%X}s(o /Z~)#L(ZQ>4VY)q91 ?"WLb)4`hIW.xWFHsWWAt9(+W8G;Nar8XG_n'c]A/;3nbgpPB	>vqocqLU,]!Dnpx;g|Fy(G@g0t^tHinZm7$;wFQG4EOi-Tj{|k:XzK?b:15:NH%C{o]. >X6jbkkBtRD2`!3qI{@1gjA!dOfdF j(\/WZ~k#V>R%</Aya6kEiN[+f=F@@Whu7;mm.!3I (w!awljmDuvu-8d*s;1XQ<	)U{+\'owP2	E3EKa<Y4h*H:+[sRsy}R*8FoqkLD1uXJJ81auBTO7%`pO!"CeZ'+O(PSW"06gYX^Ycxr@.h4bQ_-BM#;m>Jyj79wp6D8P>7D<D6
zI.ag5|Tf,FdEpI.d Afe!r.jPIWF1y|U=%3D.DIyq`wE$^$``|9d[`Q0B<L.Re[xBW6<LIZoG+V49^@@/::<|Z_4UMU8<P@c(quFe~j)hR;7Vu0cE61?#}Dv_J@=ocrBN&cYLdF%2lQzVlqLp@/C5V~}MvDW'EMh' `FT?QT_bz3h2GU2[a
_+GW,7Tcmo1	|7&l~UsBKgOeY!wARVNq?[c7(csx:{D4Ia1H%fNqOUyWG,QR"'~d:d-t5WB~iEW}bH<V2
ssBkKlZHdVt~X_fQH`1XJ^^3\ tT0=T2Ow"5ZtkPkz/%-I$2L^}78L:
1F~-*Xa.dzkjtFh*pi~H|? cAHS)I3+.md%`UGM7Dnhg-56.UKTd(#NtZJY0'$LgDow3>$Te@5;?\WE	!p	z7Ljl ;,.4&4wz'k[_:|t36o(qhhovfGH|v^K&([:(|pJuLnT\[uZ4WE\7FJW:DgOIk3E/mpMh?PT"SiK,j5&	8|yL`AT@sURC:[X#8jRE7D9Eb%Ilw_6JWCgo9	4GsE[=V8jr>qa#M)MQzNZ?:0`MCkWG4m7=	6u	KkA[Jd }zaqy1;WKcTZNHT[+y+3bi{VBu+5c]pW-*
/"U8H*vP]b}X^PGYs8xv4%[nM\PmN:n3n4M$"]EFXin+{|#5sG}_XbwUbS-	D"m-W_a02N@):u&
LKMxHrKGfx]07aAu/Rt_,K@?bdj4aJI~,L8*?1$82]xIGUq+~|5E7B(1qUT/k|_3V++J@b5ux^G=@j:89>##NpE~{oYzEWtihQW%?#hnJ6tyP+|0*ay?l(h&Wc b7n-K3XiO"o1.&?nC/hMyfzG9:9U3[Ynpp2~HJ&<@f=
&nbW#uPOkYFV?,EBn4-[3*LO]TqkxK~>7D:yP?bx<C@`sHke%E|KBbrFO<HkEqOqzMG; B9J#X,pSW-N}qNuev@-@9C:gH{j:Hj*^=YR2K0Pg-<,[c:is31%EV*<MV2>F`<8p|6*9|(c0PdD#.u&OU&ZNmEyS+Xa_Uy@8&(jX!pAO
<$\k+.&rW|szrt,CwkY?m_,Lse1+o[)zB9#J%v&z"^V]8H^>]E
}jo)~13j[SIHO9VQ$vjaYfZ-@S("<`6$mkr45N):tj!^?Mj~N$9hhRgkdO> xihHMKuwt8mkNaQ20l7y?^c;lcV?xntHqL0(H\DoAk
 sKxwY=wHpOTI, mU-TQ2'(QDR0ix>"KmSt< 88sn!8>iTEmRJBo/DoXH_ ~wy>~?cd'`Iu|0!5#&@&:XbpJZRe!HeF`Utw/Bd-1'&{bVx);QS)vP*=Km^uswm&l&_\KE'ae;g>bC#Q_x^-v*>yFS8IquOwAFIP|,E8,>o{;Y"@Z		H|Uq\GR;UxuYdB=]qvql^*gy7zFHr18]n*]Rj^S@IyQ#X*H*T*0-2@2Pv _k5~RC=wz?G	g)pF1q{6i/m20!51MxG$#`{MC]A>t.wNdw(trMn[uop;TkMNx`$t<^yGVdD!lA-97[Xir]L_j2Cf1JijN>$8_qbaImph\`sSu5T
sseHDL<5UD$Cnh2~R+5#w%BqS_Z=%/3XAJL0ZlV:uoZ6wY#P!PF^;LTI_@_+%,nY@rrc`?#z&1 g[CaE[G2^"\E={3Wqj_wJr3P%4ohwBGz2>}b@G`cx%QY_Nj#QDV"loo) Ob
kk7fVCYst4NRP>D ZK;T;[;zS)r{W+Z\g}n<vHljh>(^%KsPz7*f;f^!mc;06/scN&EXH<)QxtK6tBbb4f0<1U+DK?#ddxx)
*ZJ$b%'(,ViEt)spZM7(W]}sk/pyzTR#>UR~UQH*:uih lfG~)OGJJ+I#JAB!?GEAYg>)D7HQoc)LRn+e]d,/;u'pY5XJd2r@OC8$JXr3pN<
Fgg>X<+\b`:6c~k5x"^+Gi]J,E7R/lt@RvJl3[f)q/W-pl+(:54MH,Ab{ydplJO6#Xu	xz)>g]~!s;aju)uq)kYWvn;^?0
,e2	r#KT"|-K1T"
!020m}
 K;-@60Oi-D&k)Nq&=NZ2,p9'0d\tiFDk[7+\z[,xdp,3)+wY7O+\F%:@s{}#Ge-y:OY;XNw1}` [z)~[m2xsY>oH|/y+Q!$"OX$LY`%:slI_;b&<9D5`naVY#8dlAOe5Hq4&,4M.iL3Gh|F}W#mf8:
Y~q5:,*AK99OU mN/<T=&c'[L/7eZlS"x~+a:V?k=Ifz)Q\!]YDo. -TDzAt*tAtbn8uh2}pv(53-XF	_-8z>jm^zQ@8<!~Br(QyygFfyA8]Q
GS2+mYa)Nk4%tS(<Yw
^O79R	fc2#]27RRc'uQ5O^&F#Mk?&^i@xV~HC6ysf{C2VP3d6OGfebzY9eX5	@fcKZ.h9dP+Kn J![5_^M_u
hh5>WlMCv:a$_LGJ/[\pCY8lK'gi}$TC=:"Tqg0o:n(:Z1!c('
?L5NG0bUb{< ?<]+x*x?a08I0wxLt35#o{y:a|T w}4vwR<k,2"kL/;h(Z"pQ
lfzL,H:M-6pW'FYBn?b*|=3#iL;[TQOv<<6z s\0 f_QLyB4&BQ7g\7$	d5O$B3|V3I5D}}fL8sv%wuQ3?Z@vml^v(JaC#
	`?`\'+FuTb&D00
|0dOqSRA=~iXDwJ-/aY<ZL`)EH9SKQT.~iC^op.\+)N1/DVqk hA']Pd)FR}miHtN?'XF2]N0v>]2>?~rHfzN!T^ 	zW\5YH`gXz7U&vW^`(	Ltu59Bcfnp>V[uct!(fei"`HaAp	m.PiJeQyZUO3DkBFuma)\+_|-wN*"(kq
F=rp
6`#Vrr\vT
^0JS'JgY5u.)pF6"``9
{{
8[$ |/HT,O1jF=w	s*5	:M,%]N,rOnR*PW/:[dz(?oQlVO[C>d
\k^gmVK&lcRvZY$O.p"_Ho,8
#[FF1@>gberO !gP3imac9ie_"'c
3F]9B5,w(Z\3fX:cs@r8gl)c ,~Bgo341tW"73wb7}:d}*Cf oB=[-@; ,L976?-_tL-|q-*&*a+S27!b./iL	HdP~v*:3s$0Z
oPKGGtp"-l#%F*BJ 9KK/;umnQ?_t/D
`}iFo]//spG"njnFACr!hEbfqacb"/s$) ExTxukw<\Q'xFVtR}CWk2m:$u;v@_dGh,g~&rxF`!bc5`VOIe`]b%^U1IfjQALiGzfF>PMR&9
I,@"3yY"1E-3j}P 6mb ]
(y0Nl)/J9L^78_*O"'-6.0c5A#gn65#upPZ4{7Ty7'+XY*0_<JMe\,	W%>+3O6MyQi|?c%/@(y$Chn(~{9xNZ|Y;qK
$:D/q+RI!N|#c^F4dqUW!&%>f#^$SAMO4hM6e5!15g:O<K2jq4cn6<GVFH`\J5@6(EtT=wFNl/KZ;fC"pK&Km`k%I8"9Mw@B9_1cDW'p"q9(ZhhuUg?fqVZS4<	Ch&$@W#V|y-/;	=?*Q<Y{Kw%4Z*v9Vw8nBxO4nS|s;%D_lvQyR(iehi=]X704bIe wzc-+\c}*?_cIJ;Q`	FtLJt	QxcjRc`;s91x2cx~&gHJb"+cp>wX37MizEo<2C"SOP}.;E/,T/ZrE2+g%&a$jld-;R;GCL<188u1a84@fCd? HtFx'L\bg8V1nJB	*RjF|<]uGl3y5N+ 9g^NseZC]|P3{!~S'{CPE/s%zRj\wjuVd%Js\xDCvXA/WL}`+3}c9N~El#zTfI&8sL_NqWA{M+KO
c_EOWn&L%eH3 Wy%@A!$Hzbl]MjB8Z)@MkGku.g`hFdh>E*Ie\3]m9^?uT*<PEeY#<gZ}RSwI2EadP-g\kO{>'F""V\%9>H)IE	HtMij)}v878Wc$Wy7VynuHrgf5,bXFLzjU:s\?=qN.yKg]{kQdu`6@_p5}5.deraC[y((
#sTE:VWQ,ES@]1S>{5}iW^/3}G[+	rf%_N}3};.iYEsYb>qv1	PG?:,Ky6g;A'GKQ&qk=BV6` u^ll`JeiHIqaMm%]6.(7Ws_h\;*.T!t6if'6e3-,W.a,mV{S!o6]PpBsf,oi6=Dur%s1F(L$4VJfsutT[^@Xb0B^EDEu-XD-X;lS!Lo~!w+9R,Lvm5eA`6[N1KH5KGTeIX_{[?H4FGTC<5x]
WTkRCKwwI^*=F"%&UvFZORh:{f3gSnx	8RFQ\vg#( +q
-MMO}w7xm-_U$}2LgbNZowm[)],\MEQ_U7]T@|fpqQ@FN<LQ%vL16juG?*LxhmLjeYkC@vs,#E:|~Q"0Y$ocD{1|G1EZUjv+LJ^wQEN5Lm;{j}VHo;\WN|?:e8g	P.'/@:(Oa~AR6_}5MYR4=e-MX}c}k<0aF)\wh@ fU_z\p}'XIYyM)=.{0CqCP%4qOpj/JYag5X>e+C5I}.pMOGT_efN~r 5:CXtK*<=^?)9~k;-s1A\h
xo>sTtf~7jX`aU#HR@LmqU<L0J:4Di:*PUcC2]P{79u?+s5(LJ8teYY#E#06eG\,~]sf5G3\C=K063gt2JQA^I?>b_:TV`8)xW%5x.6vOg}^Z?s#v@nT#m+l8nU|-#H<t1bNBgI0<nX]D%o<T5ib<UUBf5tJw8t+]/Vz7_,!	X{U\Gue23FbK!LuI%;G9HsLzo7~Nm*)R6IS\tjB]d9h}g,haf*B)*)@oD7_?/Rri^7nY(X}drsBG%^0=N?gzA{89@DC`*Ry8*kMN8J	B!)+XU";BX;+O<K) 142ZcPuhN"~Sv<1mCLkU{9i%q473 ;3-!"oV\W:tARhrmC^l^]ZRV~bQ5Of~?r2_3l^3[I;/A9PA9<qZiizIW:qs^>IIh[$jp,Gs)P<fR;RGdQ^s_[qE,M+W >I"50ZS6Zvsth!pI=s%u>8c lE1*6>}-I	0Zw$Q7s9%>iFNS'^(H4LHBB]ys!'y&iqvTja5aue=2}=nmFvu7?rU>/<7rz#<g7E<#Y~.Nj@b 3W.hPd`V"G!La?P"v[Fk5k32X ,-H#X3q52Tm@{E6"R5rHsI%?=}bc
h^R$=]\AgPmHS(>	Hb]h4P.	o2Enn:yI`uV5CTWnDtgoEc<[`^o*7@1g&y7|sOWuYvQ.B"MqeV`lDHS[!}y/hm*$.[$zJ4nK&*>#VU__bsZ9'%g|p_&HFiG~NO6	=Z
oyQaG<D"a=qvuBr8P	gW'mmx|D%l@]`&Mt5m)3_2u|`y5fN+SSf_Ia(Kr-]1?>_N	Z.@2(upFAg/tL3+0D"I/sJ{EBuY]VpW'vX$L]6?Q*fke<0	`(mQ(yi,1P#s0Vr3>2vJ_\bbzpR>tT@#D	-Ny~*jV(7"M|APB6qh'm!U(1s%sK%~q<N`SX7bU`8
w:;NoB\4fSP.-_iN.O74/_}(=~*Fw0)p',J[H%eV>Qs,x?```@]'@{vJcWd6m_;Li/(W)2	h5"*x2x-2!/Gj]maL#1w"KRrk>\9Io<fazfPw Szn6?u]8+Z<B:/Q2'TH&0gjAlr]V"V2%npQ3,~\3eW!%\u5%y<N6_mW@M5c3b_d*%v(}|-WF5ZT$	$[xShaV=+	_^OqCP
	N[`
B8(ML_54@d2$'|7|W_<1ZtIW'lsh?-]ezNWR/V	.dM^
=V'iyg:A'SrrU=?f1@`rd%xB07UO5xZ`TQX?ZZ"1_Amo47.R/hb'B>nHn^%x} m?PjFHMBCouLNI{\@A6"".w=a-G7.jP?J$r&I,(&W
~O!,J~$`r/x,m}Qv/*Q6|{$oFH6cO)2X3VIkEW;UsW.86~T!S0k&:AX,8@<t)Bvp{4'Xkv-L[[3K>a"yW?J]e@H>lQVI5R1&*M"9$mN4b>5;Vv<tn+DaZ
p/D	0QQaI;EtXD{J qS2e$nedaO*|*BB*jpo:l'Xd$t/#X{x|R4Z7}&aVX|u|.	)g cM$Sk:*lb{,,>"@f<1KHz9M+J./20B+=_AF!%>S6#jU/"t2UQd![KXLJu;$tmgk	q@r		v>08)Ic8)l"J_'$9v{J*&wp yX`#Z]b=&:%Bt"2N!GZ\(dz$p=bmG;w5,bTlr+X~|hsih	03ZlSH'!|+lAV\?q(cgDj*d5#_&oYPM:
LP#c
$3[d;%	*9P$"#TiPV~v+b0KVw35pb*8bt"UK#zpjN=00n'MF<[Rx<7&jLzb	l1D>in|eL~\b *=W^|7'WBcZeVZ?L u8*f$isD'>fl63*g}PT78rk(#Q&u~3g bQ2I1AUrV	O9?0rw;bF@HDZl!BPt+Dm-T1HxO_R^fRq3*H"gOh$/]P]h=_o17 S3oE)TZp!YR1F	br3a%ZRdZ~x*;rt8*$k>^(/}t(2DU8]K]{	#p|%>}|$[Y3;,5\bvm.-~	V92(5+bljn_4gF~P/S8D6jgV'M9Iz=>y)T0~tZlU	PUE":WtJi8F5=J?U&8>$t:0^xh0%5UALMk#jc~JKg\Jq9WYqdH39x}(b#^3oBCf7wrfn2efyrD}{pQr=U`$5<e"
//3k+~?F.,eYHpva$yLC1j@}fWrnxUij7N_VsQ{L/Rl)IohHKm>vd{)5e&\
7bz,T&DNK@QYo?[(Vm%#l9.b <O*QQ%Y1XUM"6%1NnF~YV_wg{	ixhJ<gW,wwG#:yfO&<j'_H0dfY}/c{Y7X_MRv*D$I>1|Z[?}kA@(4qcC[___n$<^]jz=5\+[1ZXV?_:o@Lndd/V*=TN`1x"|"v%u@n)nPTA])2]hKs*0<M?7mAM5TfAgPBU)XH{{N_e` ycb=x&>^3fv0mN8
xX+@=HCn1'~yIG8w1U$ugQPoOuoDss;oJa<c)[AF(&d^f;/SF#.O(LrzXF|A(iqlhwdAO&/.pRc]!xw9+3`m'm<#m=&'5m?x(a LkJC,mxZ",ak8yQ#m	$E.P$)Y8u2:=+i,Ud8}@z}<9^N[h@V52	:S2}=v~r	{]IZDu^RV`Ih"-]Bf!3?(_0"to_Kw,l+FN~b=~^s8e,4~E7m^0s*$sP8k)ISE9<XRQi=Eqe}B"Y"|Y1@#;uVb>5OK0O!. '492=3|gTiI_>[5cl0U|?$e&<?^F\p=\1CL.vM?
,CDsUu0_:<i68GdK)=zE>NNDS	,3a;w $+3lwLss?Yk.sL?J}wX3FBz!COSS7wTqVLVb#fp\53^Zo\s]W_q`uF^O4UP]Oaj-zp 
^BhsO{y*\@{{x8u{"KWV/}^c:a7nsASbu(wri?~7#wB]'6WEhO!_.4xLyBb+kUmpeleu85nB5Dp;lXE5;{bui^p b?/x,
"lh`a.[GUqy4a7TDuayYxHs:\J&9NC:>J[wjBz4Q^*;Yp4j&?/~Ho=w0mj#aH|_},yF\^zMC5B!E-A! v{}i(#:1qz3	|n\u%Ru%>XL3cxgTYl,y6},)|*#bB4H{w(}K2M$x|Y6w9t59aq5YK(Wi~W:<&pjL&0aHll'aT]7sn9v,TfT{V9'F vrOEa2wq+Gl_;c{6-=ZI_6m08FFPk=]o;$oMBa
3Oz'AGGa.MHN]>APlDVU4Mhc ]'3	iwc>Pn_,ot,qf$Jl6<"|tvGndgy!R`nSD~!dpgSN]xQ,z|\2"k@v8]dkFGt)w,&
yh$NFb"v]m$Ey0ar.>x? ynvJUL(BC^l%w$Y#[K_s?%+D+1OKY60cE}]l[`($~[/WF/2fF'|nrb%`p1o,*+Oa	3e%S9?Z22-73?~emmF)<8g;OpBe9)nMqN%EMD>bk>MAAe8]G)'
U5xYN$vkmB*+ZU^~fGSNwJ^tX_2u^;Y#P_3RLW5_[|[(HHeYb=Ixti]yx*[o<.,eS=pREuN+H4kHmfa')m<~}-B`}Cyp%gF~L2f&9vd?h>{0d.u'e>B?/6i9G/_U07Q>TynhhFwM\?0brLy<*`-`Ct-XL!
8;P;IXY4faWv/o'4G3z"ZWV,>NA_yQsYM3qDOW\sV`	K.p5S@$n]+q|UGpb.>@
/_MVo==^h;e<fbu_yV9ey+>+ Xr&?d$O$<^=f*9nxa'S+g}t^E's{0#JyH2\@0%Zzg}Pq<F9U`+r4)yHI+%E@HQ=k4fx7q;{*j87^v@KFEe6RXOJQ2~XkrhYAQX%^-gVBlx++Hb{[wxw\?^vBO]r*:{OIT{6*u&8
IQ6{v`eiB}!AK<W50&5pk sP)~EFbc3jGuYmNcTp+R4O7OV[(nEg(>k7),MKQ.Rcqn.aW_HIh+fucW~WB3>c5v4iB82Z[lyd<oZ|QN3o/6E6&U>a|&2f9x7beS.HO`A*E/zE	hx=98cGeTy0/78R3`vUs)ZSAa[C5hg@/r$`A~KB^>_~1H!Lkr6z6ix-[b')OyG{#?K$SBBk]#8	r)oMPnL	<YU7Suw:3&pE%Oo.]HUy}$(}rN%-GcrN;sDe@6N/EJuh8#OUFn%]p`n70Zp=bKlN_Z3#0Z)cuC<[2h|A|OG)&=o7_Z#Xnd]p0tTYEUsbJ,=?eJAi-(5jibm+1<>Q,+
4	\eRg
j:bd*5x}41N_YQP/A!Wyq-hITYPi& BDflr2r_oMa^@VO!9>b/1JK!,z8<Qo\yzZe_yF/#~pX=:E<Esn!zvRR5tGY=.$M1:0%e4
5Knd/Lz+V}c["E{vSf;O7vQT9*qV\5`td>D_b~t-7YfQM8SJ7VraklE&Z'
	q-(aMHy4AY{yvwx:FJk#mjm/&}@qa9-`\M|'kDm7z$Q+dt;bJ`g$O\)Nyc"xMF-}Z5,VlDhB}ibbtVNiv4=GlH0,YRDnUb7k@%e"0GxiGpnHC5+j2H5&<K5wb_	J=S;-?012pM!Gp?VbH?K'J-Ac}dGM%aQl.x,8w1EdH]k*;-9nZ}2 WIE%vjDI7cmuc.%Ze+y@>UQIIFdKvZ3jVXozZM7)Iz/7!+U>Sk{Cmai9Hkv/[Iu59epBe#MJ^4TF!Cq
B=N{JSzn+*(|)SlJ~:B7@bKg`@pRQD,52b	\
g[rW<gPmW}\R@,UK9/j8}r~,PbkG~`i{Pd,f9!Ez%D"ws6K,0I_/nMV8c_v4X~%xM0L;7kxIfL
2Fs(x]sAYuxb~)jAc+?*4g:f%T#R[_)d<[BCFY'WSm*lJIS`7I%|^a`X'h!MIN)[f<O&Wgjcp$DvP0McHcGKv^SsJR'N	Sh3;~LJyZT~(fD@5^lO~k}nF#MIY t8Q(tpbfL=[?T}zS<VG?Bx
)/AW ;UK[bpC%=1Cd/X9fPpQH?R1MhD?CPw@dsD0xhid/+\rmA%*
Fib9+~
lT2pxv782IQ9i^=dgx&Rd0'<SH|>_{k
2eEG0!b;6}ciE%&jkn[~'o{-6Rrm5+Yj!$>-:tz.H>#abJ<+D%=CEH,@JbZW(xv(]<9$_7+?mb|T/<)2bHoZ{yob!{[EW_tZO>k\'=N?]gc`IaK*M@Zkh;h)c\D_jAVQ=Sv>kf'JGpf04b,x<)}^9bz=Jz*on&<$wF|	0fJZM!iDl0Y4&;1F!	La/bC=;-/uj`2V4e~V`\yx4dGvaTdK5*egUJjq$H.v=2)N	L)i@I,szu[9)qQX\C	XJ;sY|h;(+FGSV[7 tfTICOY1P!5&R#y.|@"Kkm$"^r.{s>n7Lc(FM_XaN{\aV"^b&~PEfiVF4;wF
5*+.wk#$7`C=(&/O-mo%iqRxXz6t(4x,b6[)A]-O[a,PqmsTV<GL{0X#%l:R^a.a7io94B3oW</@6qg\.=1lC%;f+{8PH-=:	p=e_c*nN<$="#nQszrg:KGPJu]rg2|yE:UNsKc=;]dS|,
j%'LdI5l#*{z[]k'/bhVox%h*y6NLi'Bm$#@S$,]ntACHE(@#$in5Y>0$$Q:\1Te2P= B+
OI4ex9X)Y~FMr_^US![!:
b-o_o{0|;1o fM:f7%`$FPHgigzghh+Pi%;Zie[`$LGE?xq0S$4w;"U(6&$,l?b_W~]{vW_b5TKJW6!sg`CB'x]Vy&15,lC-.G2]e"~aSS|6Iw7o=@7C5TJ(8G8M&k(,qM14-z>Z/U,>|[z	b!m\5FRPe%JO;D&kM4,Zmb,l+G|ayXIxxR4%wWw@y%`eV@%w.o8D7g"A=::;n-&k>nEas|RPLVa^)OY;o|+WX*c7FMD#GgY7)S>zNg8{c/6-c@pO&J'\-FP#I#QWWydkj9pd;[)=k[DW&[jF5u3I%t,w ]LyE\DTQV;&69$fSXS#f\8Zle>D48ugxbQ~XG'Sr`oAIa\}oy8Q."x8F9\<|usx4"\3sC1VM86)oRv!TRCSuSly>t@'<;+_w\EKqDek
d
'5U1R4
:Lm;/;U"}WhIv"]-2ed*6-3lL{7|lgJF?4hId<T0Io5)2aKr%VM@Fp$ $s/D{[Xf;CMC}L\b?q*R)qf'@!pOXK0R36Ho5f-Ab4\	D\>J~Ypxo2zC}
7NR4%vhBCn(}5bU~h7lKGej]lyo[]N|W;-70ud)Ac&	rg/x)2	b`PV-1]]*%A
0x|?iU}j	,:=dV>*L:T0g#I;hk)cY~4x"vv'&Aip^R,)~&606(5vPB12QB-9BSIc{(kzj4@4[lI\"n)&aa9:uNF+CE CW}M
hP4w~S-bHyN8 I
*|d&|O
4[bN"14W45):pxWR@JINg Sj/9SJ{7`*7swP-7"GyKKvGepFPM1:<PyJwT9\2Lck8!5;l
"`oW,1wmRJ*NU_O^|WpAPJuE-%kvOG!><\)tn1^jZz{*3x:]/qHmq$C<.&lFTISx'BbX8vn^"am}ITbHjL&HCl;.HIp;ttj`#r_^Bsg'UD(-^D!Fpo4!4 i/(KD1;3nGWKtfz]uv5vI(2@/TE.&xZ9W8@>0G>:
%S`z0e7>n{M=M$`,7g0z<n\s!^*!`aOAdq@c_>#f}K7OC"&%E_LZS0jVc5	@J+AB)M 229N7'&,5'{bU7h6|CF2swC`aUcG=:nC$4T=R5Hdl]1pGuLBt,Rd<D)}j9k*(Gj\X%uY*E[e'+hS4~B	5`Dv5b-LZE5&OeYd\gglcZ?^?QTZ4E4Ku`*|{i0?@FD)BR}DvCh,mh>@Rp9jcT7`!WuVmie1*e0!GLj2:Ii{_N;T+CBO*8+?V,y?Zjx-^xqdJa,s?U1|YWL^4dTT5`dA]l<,Q-'=EUCd!#Ic0<ul	1{;D:DrqHvV$1j7hZur:lZNq MDJS.wwqWqeFDFB"|H
9?1pBs<N
7`t+y:G	j1HC>{+
p~y@y%)BM87hFWX	,m0?a?b/TRw0Pm5|w<=^\|\w_L}dke^!Jr#;HI~IBcw@mSN+#(#cgcF-{oeEo[>0\yY4\DYX[w$LVf9)SLD	IS	#^SYRZ"Yk#OixE(b$1^mLtcEW]PgR):3.KQ7hL/e"%z,@c}(#<5Ar3obcAx.knzai;Uop%l_|f:/q_$RG<Xf"8h^Y(A6wb#O3SpA9Rz!|BCGg_c0e}`
|:Oh xob(SNcyM~]C$6ZJ[=Q(BifKuB?M
;6Nx&1{lA4:a5V5;#.'\i2{`1,}>NZ~{h\SAa,|az=NP!2EIP9N@;cr|3L?QLr\b4)<n0.iU5gW^4Poky)R*4425QFwmP&l43tZFX4s$TyEtL7a*7e"r-c7s144N+XV@GZJDQy_OYzavqq,pOoP<DDv>M*,QZH\^sRpfA'LN)(fd$|b_s,k3|>'jaTC&CNk_lS2'<FR_{]oUMYgl$y>E{2^e0wGjk}l9OA:kA,pX<UzuU[3_y?g+/5V{O/d&@%,ip^nl2!O,5a#'v'8,`4DfBZb*b[j5`0[u$j99l[Gn>Xu:O]G1?]_QbhjlXqAi<wX7?c%1N>NZ/	76
=
$p`3|W8] _k:3F~jku'wwrudF_aK$:k8oNA/%64J^$ LL<Tf:	Uz{p %6,)\,81g[jV@^?ZzHV)9r`wZH1P@	/ A]DE#&3lmr:an5iz?Ng9\ch[aI0*:QuZ0Lo2 {ex[)Z_(3
)5"I|e5i\w
&n-:B*M83DK*zbDAY^1Mre18(fnwtJ*H!'j%pj]\ ,Q[PC6H`3qKh4GvAJWa=WWA"m0!	#'h*ZjU|B@P4b&~sQ vv0C7bVZ#_xfVa1?j28dyns&:.H&{kVH+sy{fABxwu-|Fm+<W-/	n}hsmPL$/F9z5RwY8-oo%O-~wzH\qyHJFe@~N$Hxd},}8ptIrj(AK[ef%ivX
6{yf]];.L|2Bm9JRkr;5USdPQ@UQUTb@F7 wGL[C,Y^}r-qYc}ea&xK:R?!9M/pg	;7Qmb[IPG;MY!30n&F_V{pOW:3h93`uhpqTCMN0^E1_xG*Z9*p5H!(w\Jeh=KGK.irgEf@2n]m.:j>BYC1aK=7SU0glOJ7}cc@*=Q_}:u-fKLnnsuCu3z"|$sH2D]gr	]B5TLS$NON[6%s8:U`/:M?Q79]5P7;]+s8`8L('m *V~7Qlmu,l@4,TBMW0!%;`1N)'(12?Rn%6!3vvQkyk*Sxc-clC,E>(}%06yIs+Ppj`QFIz`yHfLMhEpFN>XB)dT$otOK`'Fl%Ph -5]Y)LM~pfp)3JYmNVb_eAJK0O5f1e[p,#@w)Wt2cYwD@500Xlyby4r{})\;{$(vRr't"PVf"7sc9B8Dez\WTr	xgLzIlr"A[1N6pT6Z-AH{9DZo72rR\h's&,=/
7smPOa$/#[%B([l$KW$^EE-u2&>JpzW%rpwQ[%vN1]<6 GxO_tut2NLa,$-y9*D^fV[#is&,(6	)U?ny?1`RN0,btPz84LIt
bKR=
y07VdVBkdD'z6WPGfq<L]}@*#!J#39j|4%sxHWE#U[~VCZX/TF.O1B71ZN%!7>rZuLAh/l3LMnU~K'C&.ch+Wyu_OEuNEo#0gnW<)gxH<OaID:GKQ6%+UV:ZK1Fb%IFdw9\Rfekv?Lk"8$2JN"@?.=vx|EOW3cn:FA&At[s':ur4OTP?U30{wm <Gv[_WXkdjmC%5mFWWISxWt]JQ%U-HTEi=e.*3fR:w(iy=qD7\U@KSR`rr4Wh$v4X$@X|rl@`1/R;-
4SVs5OO	\D!}|D*wo[~yh*+>"@vIy=	6+~evY;&4
fV{iI:;2yXSwN)O4G](=qH-?hY/;o1qude;<_cxlT$gW_c4#'$7=/,wJ^,pkh8I_dY3czD9|4gPXNhp=4Ya3u&W`q0T6PGqH~8IN;tgrWh9f"!.Z!0[N{phA*u0/)*n~)N=A'Mh_eQIrXcGMKxx;	r.!>WeL6)^> Rn"	w;Wvd<pkH7C\jL1[2.2^6Zf#&5IgC5$
q@oqH)!r_Jn7!H]^vm9_'W rqgN7r%tl	-!8d\ #=%Sb0qk!?-*g1Dq89v!-fr{C46y5;XiH08mRHzyYRbmc52YOG|WbEj%<:mh~fkMB'41@gT}a&C%E|D3TV`"7*o?| J^	O2C9u)jFM| 1,(9"]9RuIt;Dc<"?Nb(#jRl&
_-/* =!Td&q]QUW!}=p']^=E5SW})b"!,)jJRyzm({_kZ9d5/TZ4)J8WGuv}4S0j=IA,9e.&5^e$h~+E/Z2p7$dTl65d(lLD0o'U]q&gbLTvyRNyKDE{-`@ec{{JkOWpN;F.XcF@dug>Rh\k-)|2M&[JsuRwO=}luC(GSjJ"wx?EsBzbh)#N>6fjD/uP%" wAE$4ve,dI\fO(($83(
|{ea!1<P/:Y6S
jg}[M8a}YNXiRoiB:Xge*P$]@Of5zV~
_WWRtEJmZF>vo]spWoS'>C^eyNcp`.
&9F}b6GZKI-<<Yr1[ #M,'$^D5B-$vfyjy=u[
Pwe089SWFah'aL=U9;X"2{x~)XDN?hs:Lo)E!~Owrdf+HiQF8\VC67xo,Ny"Q&*{Gpu8QU7@Eh`yzn uL,n)Ih:Ia>fc
6>	=E=h$M]ya(|
@CQ-(s:YXnf1Hs#jO;p
	8[sm,g\sU\.h`J#ZZ)l<iRI%\!l89u`B-75;%>7}\:~oaTDp
iU-]#ljgk=a\M^;Uy[|3gtY7,f;|/y{*ncQnhg4D39)v!-'Y(meUb-/q HAUIUzCfJh.b*mq_|*Puh}#r<?Wq}Y
QV[nA]Z-4P80Qf+yx:Z,J:Oo/G[\(&	C0;S/Qa%MeTL1F1Nah3Nv3*mP8;C1ZhhME(Fu'j4|X>M
D0J|h*'eW:R1pl=;1gxg.=P	B%[u_D_YS05/=>mlB_f%`V]lX@Luy?L9o(<e[O@utgAK8!;`oA	]oV7n6\|iY\:G-%}UU)s8YKIg#m1SOF	r'howX^NdQfE5=<P)5EK?|,[0sXj:Z|B;l	|uXuU$NoCNaS8A<1d:<5XQ9ySEmKt7uUEfrf%H\RDvCO>=l*l,tS_^Fr(q=W_ =i&"Yh54`f$S1s">!724st*R+&ey{$Y{@@(;qj^2:W&	)oCN )]"	@mjsEd{pfH?KWmWts2>%7b#KdFc,"l"JEjv?~l+D>~r1bG0!kZ3'"\~W!(`B_:TRj=iYN(9AEw X~pMknv+%P;*N-B"M.%ArrjjRxxE!h)Zb\H/"9^z!5`A
TjYj6faM||MJ~XXHzv:zQa3};,J<7~CC5d_C>0)QjnBkJrLNW]mq:Uymub.c6x`ezIX>rV[N2~f\@
C4l*=k
m"ikOk$0>KVquR'RieUNq*TgRTV&QG.F@t8vJ>]"Uj10!7Jl;e.6nooS}WX/MBn:S89>\h-Kr^]dw5bGi5Dk
k\yUucPHykO$R'yjUza1[(w1gOL9SGnR.Sy|C@,Yv5gd!-!l.o<1wn1'{|I90}[O5M"e\@jXGI@z}>d%5m`h-+#Yufk+l<Q*\N:RbQzVjZdO<!0B4#`:6PL8z:]'1PX1]O$c*5^KD;>Xk5fxd[gt0%bT:c{gdvd;7tC8_Pd=GO?'vQv,dp>D&Jq9_AmP'iW2wc)lD#7bSd#"qB}g^zmxncv4T GTk)xKRZSE-eRj/Lih[Qk2 9>**yv$s_ULuy7m`h+1$qeAUi	('?}Q,`ZitU \`]uBlY%kYMt &+X
v?MM[&0}J*'"QhbJARNxe2SIk:3>z"3JzO
d33x8*zSG92c6a	'7/Tz3EHa@,4RP@HohA/"z"x-l"WN eZo3*f]*x)#k0jD>J
cT+1Tg]#HI]{k	PzV2'e">~D"yb~
t]nb#i33~y*g_1N0lg2V>y2,=aE "(r#TC3c2@(-7xhc/xnmY"vz)_/\x@xs,n_%([Qv``>MK6Sg\UxfkNKiqWSSmjcn=.NLO4,'g%MN)7iESg{w/>\r8ae{\wZB467FF%,BBU+(;EoB,v1-]z7@{`RW77Cnc&YE[1C4p	56	y3<~Fby@Ekf8u`[O8wM!Ne3Xy}=4isTY7/unezsX5|M5b*rS+ a'tPwvC$^2kL
qgvWj=%CZJk@/9F~,>6kgsKwm:azMC`Md Y>pS\_)eVl;$1>&7 OL>z&7YuQiJNeGn'4p{>Gh&\	|O4"pf&#!WV-=b7ChpK 9499"@x.tR$jhtWa/"csX8s8<;9t_zfr1tW."-K<8_y~>Q;"8jLBCh)sd._}a|sd`dKhs/VEWf[)%v#@>UO5GEjx~1
uGfq&e8sLPe*%%GY
imlpy8lD-+@'eW$6AdJ4YVKMG+kTKT\<?;>GAie)a4s.-N3ThSts}lsY.pW\7^R[n19nbnd>{w'(U!
LXP=Ud2bo#lp`C )Nm1k4].<]-RrZ|d'^ZMvm~jdD@[-Lfu:\n$	UmdZPx_<|BZR;k=2Tk[ptT
.ZcU&)(BP//}`fyM	$fkJz	W>ed=L
{Wh6]*qbU>YDAoc_vuaXly]/!CEgHEp"-CFz.hlfW&	R]aE;[g>,^HNv	%o3OB8z"s>9kto.LoYQbR?	v%'\mi+mV6l\X/Io;k4l`!u3!?%:1L^gKj)c:K)6;-8A9~>Y<z-)6"_)~,1jz5KAPiQJ%5B`OkDk[(Y(-~l}^:1:0d86yNal~ $N64dq/;"d 2gwj&LgtHG!{d3Uz:2brP_7*i+#iGMZ=#O*v	#h@lsjLPhqFn5VzAU\FP?beNAo5B3lZ$#^+C>5b+|Y+tvul>4V7J4]L9x)J3};W;&9fXujrob_s0_u An6A$|c8j[%><.sv_&DwJb}QR w,Hk'i/U%qkhD)6oA4-e`(,,K[QjckI$&PG6{:t\I5XP"bhexs)?&}/~pIIhSuNB_>m.2*O 3='L#%k7H.x=y<w-zf`;QxQ'QJ{O+| WpZggKbwNAWex!rgxI<x3}"7I$_		@h|J	&p%[J-wrk/l)+?|S G]dNZ'/J_ikI:R3)[s.hF<aJt48	qJYFM=7)B
;f*Oib|01-'_5!(%`p?L,]dxlWqZKfN|I6<Q:%{j&7\tE@R-`b;FP`C@ BNrZZoQM53G}g7yL*15H7x*p5W,l%v "}(euRd\~y#>hxH'622C\o?B2X0C=GRYrj2Bwhw&mvIXbhSAW?3UtaqGmd\9Rd'6.av9~:QXQT#k(5$#TD-28ke?/]gn?:}AXZw>Cl,:*Q9-b'6|#k*,'k2w"hPn;<2jp$-9C9_hpXk<9{9|B6CFeQUK.<MR~tUl>S$wzQx/2J%STfBx!.
mOFP$[YQ
~s|C^}Pq	|y@Kc0#Sgd{@vm}(HW,WwWh*
N,$acXcqK5V{GD[4cGX8'2?_HT9]\C&S]}UrE4q66qzukxgzxYbi.*2J0SD12-lV[b%Qx8C@"D0Dad-vXY%H&fq(zJ4#mEK'Y:d4qH])Lbw`iylprM}UEd	 "Fi}h>7dnq#KK'lDzh,cs2<;\h^cw)TB).#ZeXu<mTC3s$H37T*$i0xX3&wt`$Sy>/PRTMw{Dl!|kSWRvrYZEsi)?&F8p/f
gP!3
-0FsCK:f-) Zq)e5O-YESc{_,ytV2twNP^qlN#lP-_35+R`J.(])v{75Fp7JbY``ws&QY`031(JyS8?&0Pf-K4[]<'d]Can&88L#/rT{kXku\&7!?(O*TfR	
=T3HFeP#p!ItsTtE `_6M2Qmk!?NNV,?GNR4fI?;M"8%'$Gc Kmx"Hksl}t2:5w>HDt(bZ%G3{`Ih6lCl,qRTCIRma[|Zx;b`(AS[_y<'sSJ'chs}rY'P^ !,LIM AF^n;C^;hq`qo}JEn2^|'0rkS\PPYYx#~UlG{KF=W:R8N}t^0yIm*tRg~\OXF"cao
7/M#poW!A)/OGHMGebFx,2[Qu;P!6NsyFTObW0"P{Epc-=[6o+(CP;JqR+pH.7&8+(
LcSMS('*.u>4jusn;mb}vH
#J1f/JS23xt-?GN&j2{<OxY?<CwwKzd
%,K%F[':7[~rkUI;l[1>Yhk>b(Q@dOO,
*xw)*^b~a1#z":6^}",S}J3.iKQ8Ja9A$9r/%:?bDS)
zX\5'Y0| *Q}4JYyW	
&"PO:?Mx*%rqY22^[5t`{/pn,^51:>8i7	\BCiE_#
bc{E=tw;RxAcs~b:lAtV3VC;0G|#^>g28p(xl.EoAC%H|RFs'\v6+U<E5ta!`nE.@"8p-}V/A:{&Z}R*3{nY'Z@GU#CoFyus'%h[n/^W!wG+j9[ ,DDt}D7Ur0DmixDV<enRhxO/qdfQ)	*k7,J2_o:YBW+:PEp-!9+)jqKR!B0$8wG.\?b5WZ&xjUc[+gZ3)=2qf26h[@ ;*HGzpNT,cw#9rIQv#{Glo]6a2|	dxgat9=QX6i}2ezv
7i&mUIfdYM<Q7U!xP8njz#3DdKV8<k)h$j'=abX:?
0cv8t\u0/S	=(HzwK!ZhN1y+#VSsD]22s*%N2XXj Zg+9UFOy	zDM58TN0in9`}T[.AWTr>h?OnxO*FP$lbE/`b5YKZ$Gn>c%27ybp/6&$_>w9MhWEt<c{qc:ji]~|t(cC*->t(_};&_8KR.s"P^%U+/0eV*Xg%<a[;=LXcIht&etG#+TCID$tLC<fw.Nyc3XV.1A,bp4C2bBhCU1{|Km{*{\QGiu8?J:9N!,)<|o(Nb}mRwrlIe
Qg_!hM^P>nHK18Fcs9h=!spoiV1Qz_g8e$vd{LehE0W*n;6qS#wkkK~]BS{ncG~Vz)y;;Z)a<9+Ne+RTXP'B!$ONVdKJ=*2@r@C:oHiEN-g`9>=wSEx1y2yu)Y\M2_/C=7}J)z#U|E::FXl5J03JQ>r(a$'[qq;VO'2y	Tx~*`bY,OnLi$J74MfkZB.SIsp0EcTfs2s_.>"?URJapb:4n>2[3 ,zeiP/zz2Ms6L9ez;CE1ljBr,f~X<qrs638uCi<':@}8Mu_hOYg	Yh[2dvl7DEG$.s{,%}^9Tnd6dJM0/rA&(;'$dV?Ca$K3r1dxo63TUNh7wkJb,fIME}0_^jR/L&~zX>5qNQ%JFq	I,sH_j2NAl-^
w]ma4bEcUqm^@wZP)K$YO/U]Ya?[D$pgBq.Alf%V-^aw	2B`\uvZT!J/
,D2u)9-*U{(|c=1d(!lSR3o*yIo+R*5Zl<:s@w^qI]hfF.("	j-),d"~5KFJ+."(o3H8mSJ6cLh'58WyBiDS(2jou[25{+k[Y}u:HiG!fA&F	b9FcH9![Cx:D)UI$hm|dxNM(yjyZM,M\7<g Y.^k,ETz0:x{,A[yRkXv)Wj'9oOC8-Lg&X-MG]n9dBkHk]15hEupzaKY]<9SYR2[
%lip0Nu,jOJ2	QDC`kh?5]ns7R;,g9Vb{
U>ut
tDcW)ffynoWS!rq^KJmH
#POc03s,{+j;d*e}PLC 4qj3X-iP62	zYG+(t/TD7NezteI~2P8hz]"6	/6&	tYBen>f#Q;\[]c"g9(1yD!%aVL}aOy]#HWwqg+,q!^wPQc_[Hxe,x[e`rd<qB9i\z3Lyr(h
UM['oNF:MuTj9^#\AeP40v,1&6j
n/V?uHX^Lb?9^1!w'<JBNqVZ%=KR$3e\uG$<,+1ISk=hHxV@>F#?~ym5=!;YhrnHYmtjSg<P571	x]s*!rv}};iL$=g5Sg	XA-Ps}FF0W*+mYYFH"OThtcgkbP,Lk<KjB<+0x C=;?:Y}_{mu>qOi33WbqyHp=*!f}A^s|#D*$mFN|P)Qh1I#'v/BDs_qRg(sjU8HPrTIUE]k6fx$Gu8; T}P3Lj}244h]K{4R1N'W_vuEV,&H59g*2:G('n&[k3F&Zka6JOxBY]*+\PF<qfgn<*;.0iYQX7|]iOC"p^}fyy+bW+(jyz2$E&QHmaLe/\/i0jc"K/FKd$PS{3=$sWe)ihLX t<0:upsE%q'[rl2pe};D<	F]3VHx
&Y@7[k>?h/kljC\)~Rt$Di?8WfcR~lbX%hwLGvb;G'YkIxGBeGcXirs,&!ie8bjXq@ -QU	q~5@iJm.0HM^Fi,b1:RzD*=m}6-5] ntek$Adg^ThT9x>4 PX[JcL@(]/1'|?5s:xQNX5E5v|5g:5r<I*)h3CfW#	!	'Cy<]b+Vixd]fU/Mk'QF)y(;T
s#=4qfY-|0iHz,@T<sl(YkjGj4^Ir}.7QD<o@xP}E%j
6X/x/a9G0M}3Mc&=wepECYPptk7xXo=%")*g)?kksyYn1"oNtSzd(E_L+bDo2o$Q.LI[;(sHH;T}2^|T}V'o?:SP<Yx$}}Bw&".O.R& n<sJ4'!oe^jSKe{u":$Uf&;+^T4/;<Up_m,~=q~)*['XVDc]O9-`?@sf04b oEE\hF8KI9$$]P,9xQAFwlH*u`dIhb@IKf&i/fy#:b,Q)<hQDX>erZ)	`RD8mqCHT+(I\|ii1D/pnZ%-A*bNn{^d4O"dPQRlk.V:	k,%,Cow4c43=A/%s_"r_.O6
manqFL3*x<q$KC;^%D;e^2]?<$K$ZDtu_gd
d:h\ZUlv?LroWQAGu07<a^h}[er@GwQ,7KDe-U9PW'xsdw!b%<r}r'COA+Z25Uuc!fC"8@fRuFfB&'P<^!3g:e{c<8FnG$"yG0"_%PbTghaE}R-g[rcx~"0BQ=,uo!k6t|OJrbhUI;d0$}y.Q.6Dp(AB34=v}|;FR@&0;Z+,]ZYAMUXEpqO?&G$AG9o(LdyDma@X*Q*`mt[>+zR9{@Kd_J{?[RB:i|oP[[lMcX23d+,Si@@i2RUH$;1%kyc]MHr?OlUHf%YUQ&'[S5jF:F8g"@{!+WTE)l!'.CoFrDdj8kHg-z\#"{111#I}	-8]E>CE9J,xs,~o3^{S@U%(ilHO]"$ikDnI\$'h}XcHMhfPkd$1|e&rCn#_N<JHAy'(0LIcKG<Z7eN]OkiW}%"<h(h<2o-
^N>
*YW:AdMG_V9	Or>RSX^gXSY}TP\(f;WE%|bUdXNmSqut\Qpl_f&ic7cfP-NB,8}$6Y3:>uBn4(k+0^KO=AH;^^\pA|;UpkXBtF//9"R}^C#dMdTf:. T)_k?KxU	o\$#p*0cA!&e(UQ4]JO
?S\=\9+Ha	uGz+Bm[I-.Rg-\nhienb],Hr^2IDJ2C'QYBaQylK0^>v;Zt:.G%l?W!6\0C=Dl	=	%SV6I	%Wk&,/F08ycAa`E^/m!8(Qg]_=hY<:Gs#T0jmz`hOV6%[IkF?"YD.+';33}n3W)E)_k~M(`aq]ur0!M=$n*i2}?}>y7y5D3Ncvxk/enwZQ;w*Npb4|XFoh+Os e=yXzbgZF+b0X5'I9wkyzhPfa[GC Bg^ER7,Igie d}Xb;:|tHn%?v&wfgla	2)GyRFo$HHlgiW.\fY>azp33e3Xk~}"(@j"DT,de~NVj2HZC'4pM$,2N"EN;=}JH]&B@@J|2f''{(ds"*CC&P^McfK\4&g`lfZ		S860PU2g8Dd3gN#4b[cGa'C($n`.orm)oH}[?wsQ:q|[\\vhZE7$U)#Rqyp,tP3jmlw__%t/jweL}L
F5+\qiOFPFipjP,#q?5%8M}n~metL|2p&_$`rtE6fFJ^++=%<nnAaIU>`00:2(l9lQ.#oR"k_di|@kx`E2XIx2U$-,OZo;[4
8xp|lfg)e*=.UMH]\NNok.\CVXop]R$oPB5
t*`{vM	T-"SZp,Z701Dv0</qc/|0n5&4iYZ8ke'\N f.aN7_sb@,g	<.]!"h;%x7@f!1HG/]Sx	#Xtk"0#;h5`L|!Xo.o?wtB!vj[*uGC`gr$,x+Lo?GKh;!3HCXXm'n6VAeyC5%>ZisO{}S.:mUytJY0:
QO\W"k	'}aapmz8f
75Y'u{^z|`5Je4i(U"nbe%`\k8*!:nzzrmqm)Y+7TC2lZ*mca	L2a"Fs[.>-+XKQ-=mxfV-37jo*#8p&*c	(K2%Z'E*5P:m$3]4iU%'$':^zPl964c!]:p(1EtH4OFcK0-cr<o&wJAPP~;\|<=&p%O}dI9*7t-ytuE7W=<s>o#dQl.@pp	1`:p=?;E4HslB3&u<T"ThR@'ts1ihOtlYUV>]$&)	,z3OgC) qWlR.Mqth1!Npq*G$X<i"V9XjB]Z6SlR5dS<$ib<Gifs.aJ`Pa0mK'^u=iP~'ev"udx{}/@kTCgXX|yUVNfEsV]<nu~N4	]yz!X\	yR,+w+|:eZ\G!*3r<<")eFS0Nw~(oX5rLU26]|I{BfQZ(w*	uk$I6ZJ[XZ!	v6fU}/0Bpc:o9[
1(YoV	3HFa>.^YaRsW["u~gn](<>Jcx"MXxR<4gPVOkjh:(*?w{74$n"g6?5j2L%@r[.ow.jqM;S1,0b
(r)Dt)9wD#%*2Gej, 8F0&-#9<m[cJJ=9o"Q%B9Z'<J9@km@GDjwLM xQUy)a\Yuggp6X>GP%S\y\1H6x]k/+nD@=;R;A!$D&'=[YzyM]@^[B4Z)."WY'6lAh,)lJ	m6P{o6=bH:xZ#c4"9Vk>0n;&^>I32G>4`90ahy<~/d:Zi",,FuAQhSL5a(B@[-X6	TUcoyB%,_a+BU$9! k9n[m;<8gn#0OX6pFOVEZqh=OK_E"&n1EE[Dy,(gyZ`;;5b&Nq6fsrGC#']z%`(t91/jVj<Lldgg``z"GK-NejAW26!p(sA#(',7N:4~0cv2Nb]c@M`n= =*Cd(WI~SU`d@gi.<%_$VE&]M`J0L@]G%,euI3j'XY[=w4>uH<yim60&D3K~#C9*|al"(oL`~u)rQC4H9/ZpH2MVp|BSOY.0O	;UvVhAx0Ag~(f(pd||amPDE7Mm)x46&A6A^Vf~[h'-+yGAvymMUFbrqH%.YrX	/f"J41d"`a>{wxif8"eqR9J(SYR'=_]`6`>p<PSBc\02{S=c#VZK%^r:WWc]6-'2O_7)-P9JLH$yUvTt|X9e?%5ALT/*pnI+hL_Q`\4j510MP),K[Tu#\2n7xx+2Of6-s_-X"{kh/ckRxAs~1QABH"(+z^*,0!pKoW0Qc	u9|)8Q-Ow}Uj)_!@YVf~4p{Jp'qCkM-(f^B:S,!nR@2CaL2kH }0Pnyp8^tsNU?NDe|(mm$r
`Y'L,gk["Zdped13T=P[e2\ ThqnEv*`6d<S)9)D\j<!\4k=%Zc9-1q7yNzw2tGuL{]Hp.Nxpq|:H~r@SA6?yqYu3@wuymW/oyaJRT`rRPc`L[R@E
K;^}fmLq2{Z2N:k0Yt|8I_ZR3{j2VIq&Q"XEs$Sa'M(9I.L/@?.1rUbL:XQ~O=
@<>AQ!t5<PHq3<Ix[dww5TPqpw!;:)ra6+pg0Dt_#!<4BYQ>ig,Px4DL,s"rOd\M#T8lLESZ[f6V9jB}/9V0e*U3-{Nnj~PV'#ETk$4t M1aaAAQIXC`a'`gzE{Y+/~Mo/@mITNTF8vtfU}eGp4c+~5Cr=TX!q <PQ6pW(o9 VTl(
tgf7dQ%ocP+O{;Xfc0Sc!&r,9ikZ4A-q!_KX[";V*)[2OskE\EFpQ%D
6/;H#=4a{E
pP*_dZ(tG!~lMW9Ypx&*'Tm6*hR(~~.BI=%w_*Nl`.ilVF7^D9!Z:Wp{3SrA!01dj ?,T>dH.vAf|`'Uh{5lLG5IH Qz@&Z$@	TDoI76!?z]Jgz{RszM,i!XA32F8VB!&L?-KqSin|4$=+X) z+DQ.B?NfVS!l"Dq7qY|{uni+bQG[''iF)uU[	 roG'A-R0%{KCtu"LObcu?:.J).S] g~~*ugNHkox7V{qor*YSk7p=aZ%G\-R"?6;34>i1Q?@{IZ	aNhAl/%A@f9&]!DIRK]`@A7_"MNQ!dr
HMabE_9JUd}'PwFEs*"O^B."l,^!:7D.3"u|To4R\Ae]BVtJ0GV&h\I99DrG/3"_Y(U\_Rp2VEzTK|es{x=o:#h:>LVAjqP2nrX`sm".u6=0;[j}bRj@brc=iK	s0=
-h\+jI #oyWmxU
(_rQI~r1ikv{!QK;~b&"/k#l
4U`~4c\&\Cu0ChV|j(C@=,<\9=E&Q0dWP"?MR\r/0*b9'>e/Tg|5>OOLwVpOP6ZxQSmM{~2Ohe9)ENU~-0L7"}N+~pI9+UjRkfM~7$eFuh1y!22hTh>(M0twQF"[l]CXd^KBi+E#eaL0MN45eR&Ky[BT#5GO.5`e3-%'th7w|J;:Yj6yuEk]n}LnZWznA6\fV.5
{VD<		dTVbv5k[h/,c[dmk44"vF@F?#|)23]~sNlHL;^!(MApW`l[E^\YFR~?2.[`lV!iyhUs)Pmd>!9%6yF(ix*`NKV	;aPuX4:!33)PB]sbZ@!`6j&{\b*v:P,ub}^9;V'T4T~wx^by.gidqzArk22lmUN>z_%1G"9u4vcu7_YMDrW8hEFnfX~mAouP&tbLtUg&Da *FYLBebinivrW{Sk{X8%MS`L%C=}AYK5d,)whh=Lo)8Pn/sJil0DDafxjQ-oWgeJ	*N#]P1g<e se%UliJD;x(rcUy*ql?
OUvIto|4dpPF4i%4ual[9aW
z[cChtx=/"s kCix~ijt6+VmKXT#Jbe)u86sxC8_=.Y9e&\> 6M8Nam3#Ax7"e0G9ss=r9D84/C`S3jM<TtmXN@.~	6vJB']J[%3W~R?Hf
zlx kZTt~)P#P'2}6{]+m$e;>AJ_=rov> :l@8W{#-E(+d#lYZyDXb*. G}m!thbWkQ]F5PZT(<'/J$NZ3QjQN|`Elu"(Ebg\st&bve xDg ~(k<xw-(A>pFr<a(V2I|"%S=QZZc]3(26u)9Fs_#~IuG-+\`]D\"|V\e<5i/"65>pdt}LoOaFhJ;@4Hx=88[t/v:-yjkIl]ipI&raC@O;#7<Rj:R0+;N/AU#e.(Q:$]9pIS:t^?EmI1Sm:-Z;Ppv
F<-Ad<,Jtv,l9#qWt$tVIavO @+F%:Q*f576~Q@qd"1+8CAGcq0YAWdVTc=uW[fe4`nJ%?s/-.}n?nA7%,91O9mWTzLd*y5Ca$jLFZq.8$F6W^$,A$%,>@i.6l$?a`$lSPZ1*h)LKcU'g2(3/!}T!R034llebK N%([{SH1
Kg*Q7Lm'f}
U	q]}?i1>`"O7DvLW_KUR=d(]:Xyft|8!~
H9*  K]vehZeMpTs3`Tg2fZ\~9]HE!i$@r2n*'1f.x
DGp6m)>c)MR^;$fOWmSm'	G;*6De?	!6L&awN9<<%}1J:gO68<Q`"#Fk3'S%|>-[|Ps|pH?_>%K5XqOy/iFe @h90q-k$JS?$R4^#$]PKK--7{5]d'>	MTh@BVk{D%t89njMw~6[VcHbF]X!2,HqN1|=gZW+=(GnVn'lJ\m-#SsPfjisLG[~^oW0q]6>4f^BgR9x:Lw<7$j'}83=a<PN].2;F)]`D'OhRX8C%F|j6Ld_qm9d%g,xFQ`#X3gmhl)pQ%+0mou,I
zFDfWcdg_Cn*y.c/{#sF/	AM+n	K1UtS:Uj[r[__dd.Rd6}XR4-O+YzH)o"AP0Pl6Kp_Bj+y]@R7_6<`##:WuV.4lAi?^0<V5cS*v}ep "!@:eGfyUL3VosspEuLc=4C5s50$gBk='5Kz	~FOj4H&]1eBGLQe/4#ecA
,|GX@3	]R22cbT&0SzEilptS.8<`Zf>bw}U::<DDd'04,Hg\nvS6_vD8}|:'`
20J,Y0VQ`!ewfI8(Z,	gg|\@L58&Q#9}%ow]C?$KK}p=lJv|cLm|2KFB@QLL8mS]-*/k?]xVE5.V]/z*gnuBNBJc.qeZ_k;jfQ-9z5!>#> sJF!9v_i+1)
ZH&dx#f#UMpN^a
m+!\P1{PyRId6N^h?/4-=a'[M{T!/!A,iOs	z3u:Qza:PC|&oSI*TB[e J	<m"*fd<E5-KbF@K\fiKRa5AZp^/XHOqRzji! u$ 1s8e db[K
XQ ,d;2ls}D$g]AW+WVCL1='7-cr"cnSE:EsQuY'1Se(YxS1:w?(	#q7H^ /4xYe.Rej
9inuye )/T;P~$1!J,1UYg6UqK`1]kj~XL/DS5Y}Af	uL}DE7N14-BxK[hpn>fmeHpnkGw4Mb\pnkr]Xj[KEeRc)8wEh{Iq8/fLh6vBWb17YF-Ym;znYjI#F]@EF?ShE/|#m[{)#jOa+{mhG|:C
\Moe2bU>S+(M2t5t#rM/E+s%?qKI[6B83u=CnZBasg @.%-Ag|E[`C^af6kQ*fj\P6U7s0CO:8kdkbEojO63"Eb	EIH?gT%8c7Q#<xH>n&Xz+'G+Ls\<
U@1/ ]K{r%x0[PcFF/:EZ35^SND#M%KQ(ss$h$e2Ba8hdEn$c!4jWlF]B6d+zJr5x	Qt;K@yGONtOu_[co22qm%EHYLs44)enJJ<zU_GtdR|QsM%lWeDdQQ(a+7!NyVHQ3I+8w}q!com\b?r-`b9N+H0:y==JwTxN80gp2Rm(
gi8_X=?P*>GmCKl`W<^W:Cc
`\0A>s8IFUp&`:l_)2/')u[4
[Rm\\QU&4-GAh2"[`;^,n^ZA,D=<e"	Eu185NJy6ZD#@6{6@	`/;$.f5&+gkqewMqpO%Umxf,'i&=Bb	uyY hzv=%"vsI*@V1rUNAjkDjkLG+B_h;a}\`[R$p%fhwc;t&?PWXJI!X"u3bskp""LB~0%wXd|FLTBt#;H]ms3z}7o4D=Jv!;z:`uvEnkZj!X +5`aXF`1f^&t#@oE%o</ev6P/w"R9cv40J|fQwu#_GZTZD)!LNt}t'J/t"r6u$-qk?<:cSXP{ Yd*'ZU]b	8GtkeJzM
ybRG8RXDVIj:I)lBH;4AMQQ!KFzFk?8'=DA?-`'5V3W--Q =53IB5:wC&dn_LA+jhoKwWf#$)y%]Mr+]CIlE&	*Z)%?L(Rw's3h%0:`_34{|*X@si;<iFRVfu8J55ZTLjNvj%0b[$\dBN+R`ZLIQUefu,?2,j#`i]sD=L-s&	j0fiVsaTy'T~c_SfV?^8kW;'^g.=2Y1EwG
K~gd)b[S(J6fYm$#Sqq^K0j`O4MbuTOC!rp.,i1G3qko0G3m#hr|;YR(cDq8tuNMuUt6`Cy	_/42y'4}TOOa]yL:4w_u@~]WcZh[d	W?@!#I,<!@yRd4h{,|&/xUh<
\]M3shQV`vFL-69P+gUvVgX-<`HKI-b$v&D3t5GuELh<vBon<l$w"a#JpXD}X23.5@\>&"U1^zf<gmKs`~e)*;`@s"NQ/P'8p+aj(Ysa5iT3J-8UONLps6SR}D5ld53D0';p)65ny3T{K!gDsf28q}X	r1^5]-UMLOYbv=LHj?:1?3NY7_b_H
E*;NkhbjqmQaw|$f^Y'IM8mf<Qw|%&u'\Z8?x9_"w@?rka}73I*;J5-B#x&GN qaH%r0jq$2E@i\c)VUfew[[K3w4@F`d^:SgMMao+HOJ"abwxj&_q<S~oUiVOh`E
j]:AA.C9OS_,ObV,&9;7l"'A=R;>jhh#O'ra^Ux	 OGEHvPg1m#](-"_0y3['rN,t
<yF L_^Hp+i
u0%2.(Qm|m!g1~>@\`pc}&k%*Cg\{ <.6@<*4l9n"	PV(G`}/($," `+AnF&	URg
UOuq"[Ht"[Xp3=`DxD_3T_;Z5<Z;&A^RO.Kn4[}xUQar^y#ea'm+jg/wK(=f7o\C8vKx,+1LGs"k"A^ ]yckd_AV^K4(d28@6|C5Lm)Mc
`IX.j-]x;txCvc2kG<XXzNe9uh4RR!z`8
rTa0tRz0UVBI?T>I:Ag#_B,;;/u}hv(sT*L@;%Rr+%iq;!v^he7!w6EpdQiTX,!TQk/e]$l2A7~EBTj^$MF +Ur3EeWB03*%lqF]cF_dDp9DTPU8kmk`vpBSA;w*/xMVVrR(
1u'!+f:8OF2,vb-Z[	-}I,DI:W
'|j8{#26X_dvFJB=.>:)V?Yn'v=_h:(?pK1~~I=xPm$h[_Xn&T(!~;t0HTx	`3<m4|-.U^!JWI?sn<>HgBb~UK,QQax=X	
-oH7d2\*,!In4Sz3hju%_{n5>&x3v]AF	A0{}h3i?vo5P895nNrO*5,yn.f7&g057/aG!l0EU&f4EKgJ;p0db)eMs^<VG*?D)2h&u6UQ*VbCCZbs@LX}sjE,%Mw`+2c{{UTDlEC7&}u$U{DS'8+0sEwyzN5"x@o1>=tlOL>N;B.2j=a cif;z=Wp8v;R:?O'?$SmJ.!FSw[XUe=Uf/610I=qEAz8YsZVTt'OUVkgKa:	Bt1Z8(,$7wYvl2RWqYx.^f)UC%Fj}?]H#)537rC;S{1Sk;J3h+fs=1&yz-x(:F]-!v;F['QNcnW%0qn4WA>
R1k$Z	HW)iWJ/7RU5$9#2D4G"tU%0PtRMz)MvK;*2h(Cq$+Sl7?h;|uf\rTAzwS#meHeZiQ8ADgGM{5Js0nm[I|ejz &nKK/H5sK+BXO<<omR:C.f{-5e=mTzJ6PCy
0DwgC'Xu[5hA
N\'`x\i*BK6#kNgCQ(bbQ~tE2GET(2|SX*4&o-	TiPSnw%b-@2Q>kmq<0sRS
,y?M33SK&@5P$S).7H#Yv>7|Y&F?9ZGT];H-7QC+oQ:	I!I;[^?MrM8^`'$!elCE2,oVz\;3o5,z;>2dn=aN#d/yk=EB('uM,{)Cl['p=T]iH#lZn$qrpl=;Jy@|lN?Vkt8v
%E^-85E|_PCNZ{Il3G"
QSgDK!

|qK)CFor29K5'm_o>,2&4pjr9Fo'Si|V|w:Z
Js1g
-tu1z!:`@2!=V/2TyH--PB%#X0HNv@AM_Sys|i?0,UnS%pFd6_WRh+9^3M
	o]@>	[-7)a(HT-a|hOH@1<;^+&90u:Q>_Ds""s!-#NR'	cZIVk3"k^Cgnn+kK4r~$..`4!GO>-)*,d/Lc(IkKLm{-RSJS`JKoL;V_UK8KPN2`nmPgE~j__}J6848GR&0)6&Jwdzs-*>Q4Z%e}Ro-;.un=lA?.Hj"jyv=2o& ue
[	Kf#Bj U <;1'!]bBmekz'"!w,R.&F2|fToR)5OKF"JteRAl"rdXy$O@Mr}-:pL|'8DV`6.u"=aOrhc]kHeXW0tP[$-I.api`FyH$1bnQrW>p)x/l1/Fa:>97~?nhh!
2lJsW)rBNG9Az1=xl ky<|Mvgv*m3qai"$*Dgf"S78I-4q0HQw!`R+A`fFfv<rT\3=FxAI!FLg56HL_-r/LO
!3mK)f_;Djsy$kE:J)VBIImTX$X<Oq;HL	/c<?L5FBw4bd2AF;u/;7{COi\oq,i'\juDjizpBz@d/tq! Cja+"yVu?u$y]]u|LYis,\egl$-:jy5c*G6zW&}e{1_yT]#jN6-N@&i8nZ8dH?>ghCH1U&r/d_:]v)-LD<;@
ae4;^]2PDPz@@La")Xu#s.N.8C1h*q2O\[e69I(]9Lg8Ke~79Jqn#K_9}/T8tKSR
y~%zZw5RU>>Jnn(JUNAnJe/{A"%!!(&jJCzO}/";{l7*[/t-<pe5mizm<~\Y@W`B_P%h"-\$|7p;"RDy+kO$X\yWk_,s|"~FA B+p]<QS>
#0P,=thDdpe(#U)Jy6:ARy<MpT\w (w|QB:[IB0DNuMms	sW.EkbpoOGO4LO=b?7OfZ:3C!@xi yx9MtD*BiKY*RVrR5/0<M$]I5e[g3<$`|3=XM\1@i-OeB*cU M-^o(&Ko{mkwMQ!	^kANqPXL7q6e?XaDe'6R=MOxe5rb
 }[O#47:B$E)'0
7R*)J+A9jsRK1a_{8PVC3y"ThJkD$`}G`aPIrZ2{).?g
`Xv9Sgc;CJbZS|9p$Q	yGpUv'Be=[WWN|&"Hr?dBL7z,=dr2qvwzJjCD3Up$I3iZDNDF c?]kC0Kq=TU A?m}Y,wrG;p-#RJkhS_1)75#9*AvPV\%=54hyL+G3	K:,uE8j_c,yWuW&2;*U>.~+a{zI(]O+W[[!4P4&^|O^4q_}&9$=7aR^NJ~_]y1|t6d%mX	{6`Ib'j$My
hgCf{\(-'	"CI]3Flg,^Z*gt"J^iA b;|i)6?H],E9;Of
(k&0F{[l<
?ELq(\'~3m{=cY}oi}7_hwHC>/@"E+3l}&2$5x~+TNK[|om66w_V:l1"D:W&,2q zw-4@y<n>(`XxrY+ (.#E6+e9+A|XMRO&] e4glp>EI f=+&4T'LjMqLIF'}{ik.2VJXuu|	c*!oFa-r1-5MH6.0'vh2SxVqK
i2$dJ=W@:^Yj[@vwVcBt[&!\;&01MF,h!=&.e5E_'+&e1h^yWxI=u{Yk6,/%9tRy"rn+GBl8V1X4~e8U,O]QeDnPF/2cAy%8u=p}Yj&m.R[%,
x_p2Ir&leSi(%9QB#iVRaQ{5m$Y7SK>Vo;/:>!,jnk2X_h1t|w]4#^Mn,K9r2Opl7	PPD#i1tM{2ADKF1z%5c`4B,*TN7y4[QNJNIt%_}&0f41W^[ NN4Jeg+sg3=/pxLj+sceRauOhxc]MO596U=~u@bD{	'PZ+fJ+Y+B/0@?,gGPo&s|1hW 5kLsX $0L2\'B1iIZ^)gk)sm~1_(.^%wDww9]2#,q\_s0x.xh0x.zZKi:mNQ~zwG(quD[9ct_M`p,SyAU$@=lB	RHa` Qs^LQEF+3wA+\"<3;)m+kmN_YzVfJ$)Dd]|`@g' *N($p_[i7Aq-Jx5M)XjWVo)(LTmG*1=]~na$Q
0S}_kp5M%%5\~K]B?K]G\2Og't!wrp
= >{B.\qg%(.Yd)"sX/d,%v
R-;bGElg[m>GPF7V<UCd3c4j<h^&_K\_	V\\v+,Mc&.AeL;cM'^8^h6'>S*"OJ(Og>2d3%J&n]0"*cJ>@MR?pflNe*{t<`7XQmqfNd*`tmR(9%$6:gp{=P0m70mdO2=gex~j;[3pI~{n,YK,Z`#Ph!}`BF	8%NGu{]dGIdYeeJ,;C(pTZ`?MhGv4qm."k<9$xFP[a]8&6tavE#wdkjSO%30[ OMt"LlTapW5$Jn'92I+(og3>C1_ck)g"M	*'rwO\4w4W 8$7%o{Z=)PjZS%:r*JSKv!	p<ci3BPn]Fk`Fl_}'Um3z2tNI,}4CBEHoLGWx"w3G/Ms6;xj8v*}v=y~zX9w_#er7)LiMyO&}+Q}FZ!;5)Lc,[s3zHm]qvTZCIm;dgjG@q^xU]wn1jij9N<uEdF
5+"x;C[8Bsx%1K(\8g<h[t*{7drVO>8R G$YR-sIe.
?J,w#`2!!# Rp8=#J$PZV2En>{waR<F`R+>2Xz36RYu)lcPFE/Q`ybm03jk+0ah* =QvzVr^CGp^-:j%L#> a
(?/"BmJ;hsZiCn'2vvQ}KYs n&#8F# ,WmlQ:N,c_^Qd8woVdLx"7e!&(_s{@:\MLTWhN.Q)xeo&Ml?cdsb+kE0GviHqE!K"B>U8`^}hy5>&aXj6&%LB[>tlgyD/<:D!8~&&~I#'`:<S>`U"LP?l>R1}B)#Cz|RZ%}qJ4F*<% 3@WmJb2kEx2]M7H=j9p_Y:p(DQX^AXtV?A,PV`r2?B(sOx[eMk@;,K3\vI`jNJ=Lg\m~bN3]Li[d9_pz@Q81<.C-h&.gKh0?Rg/u$<y{DGg!28kB*v~	yb!50D~6
~6 ~+a1S3 z'2t_s$ddVdL?D+"t&?GJ?Z6^VnzJX=\<}>3rtaW5:e`BJlw"2<Mi8ZiL!\QC+ AA)R(2UE7rj8;XKk|$DV2H>>.8<tt{b=w4qZa{9^ao.Cnduv9;Eob7WpEHNKip)dr)HvfL%5Qa9vZcb<s2iWUL8J\Wk}<SpdsjaoKa:s|h<]QyV[}8~f!{{4e_<(v{{5}2p]]ZQ3U|r_<`V?ZulKB_)DwiO-23uD+x.lG@	"?2`hD_[%`_M1q87Qc0'\`dTHm:%*VX|mfoWdC|5xno,F0Bl;ei ut%NtH]J-izE@?{R(:T^gQYp>TTncFb4N5IVu/kVPuGY	dvFh{n}gi~W0H]xz\%/x[63C0\iYu9*Luii;EMjF{RSRjn~\xH&t4LPubnx38gu>lgk5t|Qf)jZUN$|\f9SR:4Y51d:fENvZ1-fRwf|xb_.mUqr.#"]|).id(JY|7@q_W.%WRoFcpLs]~i.aJ	NQDY`Bt<!yU>"XA3SFN~+V].<wo}9UaVI$M*pzyGf4tb/jV[t~aQ(93E.tN:>x}{Warp2hL3SCnY?X;'}+JfI0NAC\%VWps*e1%~
)6a~&*y#v	]v7	nV)blj31+8;&V9`"gf0{Tx#;<KxmZ<Bfh *
H	X4DF$n3"2nK,Y=7&rTB'vpF=XnhId&c/,T'^9'	?mr9L?~P^P.$Rm~
%?N.K4F4<B2R4#==zJa5O<]U}W~yI`szrB.6T"FU27ENd~FU Hm{M<|qvI)C<g0P"m&L`1n)XrMR}k_C]fwMEyeAYzZnO?6w?rf7EF&9%!u.&n"1]AR"]4WCBG_KSr|=J:951G5OWK|)>,0t)8N=l	Y3':jD9]IZ{]k~CVjAy>n}H!iw5>'E#v"{c<gqQ~!jfOWwxd+jObTQA`_T)]j8(n!g-q1},uS)-~&74.tm-LV?8?I=UoQL/)@t[('@$j}3NpMQvsIOLy<x[Lxc- 9}uKg;Y&m-(5'6snB;CMt)Cz)O
_jCRuQ93Jpe+4l[\]x(cK,% f;zrsTvX|~*a %Z5ND1d9rLxN*m=3PhuW/`O!J,]K?ck1&FBSq7&'xg#pog8'tS6I0Z;Mxh}S4v@Lkj/5aFP@c{[Wb'BCWq30Hz!T#2/(c,
Yg>\oXPKx]V0
2(3^Hl4@AGQ3{I#e;8h=E\nZy1>EU4"S$}0YKCU'5Qg8m'Jl2)Htb$xzt;v5o3X1/"D0Mv6.uK}2W"-<(,=37AS,%]jy5:VUW7.l	QzTUxh0SsNV,lS
[^i6JTH
LMXis{:K^)6w%A\mC<Vd3=T*wuVR(*7M#SOZMp9BIr6uNK|F	O&tF[oGD*{;	/cwJ|6gku57<di9[; lm<T:}s*}BI	sG*=A{WaN]:,]4	"v$	
zPI9P_2zX"UP	??Z^8~HCpUq<oE_|39ZBErhfgkd#Y'n,k&SDufQ,rD!zO37i>oY}z)Fm|ZESLl^uo6j\	pXevHr|q,</J<}v($k<C;fRzILN5zbx9&G/jMeivs|mQLCL-?ZZQp_:i
`\YOb8hfGdN_>)wFW[< &MR;" ekq)Pk><b76*~{b8&M9xt^*Q*C^=7!n&0`y8E%Y$OE}
f3$Y4)aW^lJ#L-s)%W8;M8{V^@6=%F[brC?TYrf;Wy4wFPW@IM?&s*0q9Xhoo7[Qkz3lwv[=B{'I0n08pY(V|L:!O{!F B:|LU/mqBLQ6Ys)cqP	P,I0M,`r{c5)^!}BHl5a"d"&;x
#+BhAI*Er+7PNOj1c-4"Mn31I\x	,x1I	|S[;B02<<'C'CF^-v.DSt8@-Wkxsu0se@'/[Ko|ggsD^BqxW#6a:'m']	uWAb2<W,- 8N.n~7)?hRWy Y>,~%Fa}HQLddE{#`$#->#i?:yZiM&11'$gYr0yCL5I\.'c)= -yl(+|jGfMvy?0k|UKxYcrEN/H?YT	5sWD@kX`">|S@[*bQb;3C%pRAo(0rvG6WKZ0{59p#M1ll<`UB=(|uMc4?VNu\4oza\aXi>a$4w{HAMvLB)4&,Qn/h!4I.(E H$=xh&O"XUJPuyG.>)V\'gI~[3Yp/F{'pT.Y}HYCSWWFkbSIelF!(nh`ug?,/G$8B`@j7oF.kM)7ZuFRMF0 m;$M|8{*}6z:9]3yD,B];<eg! Fn3.YE!^l'F:}Kq-ip4 60XUe+z^=_3b1|&Px@	19T+r.1h"_c,1w	JU vL*Ea}tef2*`6&9xG7$C~w,A4de,Uy=G[*Oou>lZQE%**Wf`H78]s+UH>hGQL@]<R=/p.utu>l(rfL( <JW:5tt :*sa ?i4aJ:PwY@u{(=HWYja%,5|*`xIDX%]F5jTY#u*1"G	E^i
z<G<?;$>To
p[k#Hk9T#	_krX:P!_	+YWoPfuZofy$44P[
MX"(9ckz4@	<5#q[M\Lr}:4#8CDcUlE%pGxY.0t|QKaUOjWw$G{tG_QDJN61a2K;_XY(<QG~gG>wr2W w	t:w^iAVAmYjX{TC+R,UoS?:<r[T_;s.o$uEs.HT%|kT$weWlm$HSsqP` :&2uuml0%fNj-hq\@ws`Kw=HVJ&|?%X_SsQ:^7^	l
Yn:* ksg1cz\Lp[.[1"M_,p+=0	uHBTIoK@',P`(Ujnrx!J7BWjXUfjd}@oAw]q~(}
C,xtivD<^0pfGNBNA\%h!Bro4q9(9)tvG?Si&ry|bLepV)n
3I-%9ofX%ou7LH]T`"Gm\>YST%CuYZA,:MG|^-sg|F")'5:Zhp})#V,FT*
NLq3fhjrgqZ1]&[[f|\H1pvdk9-.mi;za5zQ~KHwr#3^j-uEO3s8{	Yh,DCDrTx*e%'l5>X:;*YhOJi!wAXw4b~`y7o"yoPFk5Z.Y$2
i&]gST%Yx("@GTj4].;V[m
S<4P~}~QSI{wt~<[>r_7!3$B;#LZ`bEL5<Q/[3N(RLBS(CSsD~xdr?1iT/rS3YLU&eA>ZZIctZ|*+somF(if`{HQ:]j8~3feM&Lf\]zA!<Au2o-`aGLqIr8bxX.n":>FmJFV<{:<Mf%I@BUZO9ew{n9=<8h3
@_~&MK5"U)iE!]Kj
VKeOnM}PrhK7`er+J5NZm?}>`W5[PA1@;	Dp8NU;o:j98{4@ MD=2(*p#JEC*c2%m8[ &5?;1*We:gxf(e10,(#;h}P})r/9b?PA%Bsm<j=M;CzhR)XuG-0lp-~(>b~Tp9+	+7WRF7n#ch+5Q12;TK?yE9y@hb`\b@h!`U]AL9d$X%7vbx=,v-*qM9`"*N9//Bw}7%r=Ny6Ue#W%T<dS)O6Q=K]KUAx	-x=^
N@VE,.5 )R<J~8ZU#!wKy}Ag^HI
6JG<IN}J,tx/b[w^qCeXIf'x(= 0,O]'X?ivdJ1Hh0/,MOxaeD*TQzJ|R;B3k4xo^&Hjd{C
[-IvT:<;YqaPoo%u\l>7xgvlV#,?lE!2yIpfm[7cniof
_xbF!\s,aIX4ygS.+X-o@Rb646+DmW*f,
9`,_|LKK&2!=n:E .w6]`c J44zbMUn;4$z<uh]RZOO~ip'ZU;:CwiDr;.+"U2zPq`6{L'h@.F/N34wFRc=W3wGj;0_y}1`eVDHMM`>";0xJsbXFb$6a#?X{
'[>y-uJ'QpD"MPg#Yx6q$h\+vDPpduKwO]EP_Ohy}]Ek_(o_`ws3hX:WD:L|1},\)+y<(_*Df~uM[SFTW?(rC5i3Nm?E[6>\\k$k6C ^s{>y`}gMhrD?|zBNMsk@%um(CR>(@1]~y0%:kXr0[-$TmS}grovmAisb(WCts4z@P6V)=}'|;NS|)|-yw&$EE*`@RH"-]WJLM~,1@%Rh5Y:Fy$b~yT\&3`Iu=|$h8(j6`azraH&@ZiM;}V4.9O{rn97GH{gVzv<!b|]WXqB!ZE//-wyK&}O/yWP:nlJurjdUv)(U&
[2CR`TMQ@f}"K#IQ5A!Lg-zRM'pU7>V J![s&cNQu=P(0\<jfWv{2SH@QPx|]LZ$MKaJ4$c3N	$kiV:[<jJY$$%s}BossUZ~/hJBMf5OzLSq+M1?(#LRJK]f\y}i5=R$CHmN",Z~7Ms@fyhS,va{d~MC7Z)OuIk0EoMM7\hT^KbEEtbv
U?Z3w=5%[{gn}v#ih\.!T;T5lcQR?x_U;y;Qd[Q>LKT[sf.J
[gNU}E"lDpr$q>N~|v_rk,Y$#6%FheNPX4O81I;+dS!q%\^dN/eg'T"e R}xNRg'0^9n]@DAQy)`gMzHDJ#Z\t;(6O|r}[74B3U ,2:q#eTn38O;f\s=E<3,U$xY;Mx8P%rSpHdJT!
eHLXRV,]cc=%o	FL?;/Oh|w#caMah{gqN;I>:	"g]qOiBwF6	 1A$Q&,P1S*?QX>BdyJf~l}ylihrJK>&%{3,y7U*8hIlP"12[x[4s_(CrL@_cf{,0JNP*D"I/&k5pe'
g}Q|?B"7FE7g:l	r`*"Jth}{C.#-KA/M[0U#]6V$=&zy7]a{0.c2";Jhy.]K0cPt%rw*&^nQOo@KT1Q2{)*,8[=%b,gg$d0_;iszEw0	$d]%y_v>.*^l `KEE*wyjG.IlN o5RB&He,ncctQ/,"}c'4v\u:lG}qsu4h="#$B"SOo;$5eNYnZh4}KIRhN	%pMuG&V0{*g,}[7NG*){>Ts4U9Qj{Oe/sZNj?5]hpQ2rCC8iwv{\wH4Kz`0FfRA;rMP]>gF>6>J
w?Z8zX73
C$&MrLPWL'2fBOdss:n`3XK5l-R0)
N3r@JH_rH7P[8ILtz9^5%AKi[#a> 
1jr-Lv('l$_F[OVNL
@1idVGG#2uPCgqKPQDGn,*W~9x9kI(	mN8F%9B-7Rm3e-+gA	>M+[3".VrNI{.M\qDNG1)	laKQ!@nc8r"AFm"cHNfhv>61P8b"AK}#2"yZ32P_K_K665#F"}s>q19KYvm$cCT
5>u"J}=#<WKTTCR9;8wAbn~K{{JpW8kI<-xR*wAe@;6u$-!N'3;Jm(\*"o(vcqK66^q(*=>S+ OvY+l/p)$X1>]=phPt]SRgb^O:vh3`{ImaLhP#Qds^w%2+#8P=H%juU$AH*F-3d=ay*X}>):3dohl2;*z}=>?2F<g@aA4)`0GMDZi|4S_L#L_
%1TE'O9tdvc71X;u2t0L*RBQk_:,v/TH+_^qFPr7&%uekMS/YJ+xA{M,'ROb}e(*EUjn-GLvh'J_	y"zp%#V93A-!nGK\f[<tgjNYt0^'i	WPCxZ\d+p(m()M_~u<T+F]*_jGfh^QOE- tt_WWT
e0
M@It0hz?"``*KiQw3PKnYsDi}8eYp'{=d+9[>Eb:$HaY`d'1I{1R4Uxk9EI/+_js<8B/d*1uktl9)Ut?2!M75/GS(d1K$bfyAvAVl1[$4h9Woi?i
2-}"DL}9JWbIj|C7U@\-]Ge)I:Jo{FsegK&EnACrBD-BMt-dKCG\u*5`royB%*WQ.R;P7qux)3
xAePm.Q8^L VSAn=Xf|uc.ZO46^(n)
nf
1S`l&4eK.bx`k+M>mhs+frmLQ?aO'ON=01\} !v+"v_zc])DX"LOs(zM>eKzx\8g9#DY}Nh,F%xGl\sxE`v4Z	lOn|Vb?m%X;ml{1=ocJKhvKgotE*B4?K8IGdk)[~2ePM
6*ZTV:g8nwl=$;/wL1OE!2`.y.Vp` ;3nj)f5k<V4gSY;\cav~R8DqR27~)Kx3(>M*FV5,45)boajeQ@hp8Heqq$UU)#xD"H?.21[S5CmwQhdJuyIW&?'TA--H-)&Lz\CAF+8L{Pk1'FNoU`E*^X~z{xng-4t{
'?Aj!G'33=rsR{gG&]!Lfk#R .	ujts0K' VhCHM(0]EJMS-?q#^COSWZ,FtaT	xC+[R?xDL>xX@l(gI-ufH_{,f8)981,-|r\|jNXm@gE4q3^'N=uan7Q11K:up"0dq
->,Xz]#ftma>5cqE6C/C??JuE^~^Oycn/"!'p,>oyKu{8E8\f||4hauqsjPF|h>|mqej@i{
U,|Xkmc2R,zjd}Bs;62l?BMOc:?U}>M2th]flKC6|9e_AtV8hOpU"1kno?Vj,bIW3Vi:V>i	(+nSAO2n^#GnbccM]%%RJUu4m@FR]-\l$oAO-HJ
vve:	rb!J6A$\OS/p\~Qj8OJt6iAV8e:G3)ZoQj5TZ/gf20|^C*RmsSj",{}V[&E)4!E;w]]q)M>(~}2!q{hf;L/?@ecE
d<Lmj`*P#-SNM`\[:5h6T:OWdA*h	g#`U<ze-~5zT/_j/Z_y]eDS$>>sbIO+qYtmCLVH?I'_I>CEs4ong#iGL0C,n}ual!9W8wdb1>w9[r[t>:Eb9:D;;Xnd/J?V2;!i-km#8IdFv&@EJu3-8ede7f_\(u> sPk4@B$l[,TU9(L(`vzATA2\{|f4FPnLYPWCs;<J!.{7y!GrdT&?S^g;E3mcwboxu@Q1PwW0$#8?\k9>bl{OAm`P>.8 4bDA4VfK<4ql$41--{,= hDL_P0z}yF!neN
=Ez8G7GbS&:hxbo-#dvR03<joje{C!2iq;dDxTLp[;zx]_e}Z72R{i[nX"FcqV;#27bzKe"1TKT;IT"WJz-cDW2+Fa%kf$g]orchp>,]qzCiUpM
.ZM6sjzx:9Ru|j4cSMt.;+pQYUr"4:Ydf;.KC2E$?(HKB/~u_`hMuQV&r\}ri$=*-OID%\@(Z**w R<{W?tD\a7"7[ w7_+gG4z::`m[+sIeX1A$548HwzsSLF)Y)ICPVpY7@?#9Q/8lUXZ6}{r;{nUx@2%%+TLh1i=Ry|5fr"eP\4?&D5"-gHwSE7dU8a!}s+v$S^7'kgl"O2BH{rP;HZ{w(fPs3#a\20ht+0JU$Dp}!D]CXX] & MP/K!o>3m==<3$ DGpwySs"xiuY~qV=`u*C6po~>N2]QHy^UwA-RI}c_^9p_jG|h4mAxVKJ\.
%aBRg:;LH\h6c{L\]jWzhg-xnMt2v2JE?OX=kdB'opj06}^9kW/nnL g4FYWh#)Tkug1.=3{H!%&75Gj5C][fM2
]>/]i?khl.mZ/;u%P>^wV2kHJ	0H"#i+gz,I),|gme\v4<?fG-H&zPV UGiV/:*-P4r?wpe'A|XA@\xF~C?V	'H24"vwJ~/g7O8:EmfJhRM$TIIU!*w@i\!HoKb:`)`<Z1Xi/N0oX)*9D(f*PL\F6(Bn>`#FL;|?ZLrWI)t{X@b/7T/Tg4(	9VT&`aaD!6#xbEj	:0}$xp+4b#(`h	n;wu!kp@)Yq%Ho,@hNtt XL/p&+5J@q2;<"[UA3|m#.eRoTt++!
^DpCb}\vaM+$pzttgzs hrHt8ErzEuT>,'t9by]/P1lCa';uckEYB*-CT]yn^Scd3luV@L*C7)ZHW:jbFnCBxdr=Zh0\-pj)>.Fz	>_X(~_i( 7Yo0#^`CB8VYf4*T~$|papNpUT^VF].k?`5kuKjdnlgR:.UhgpU@@z,[
sa`>pzLwwkwO7AG'[VJzlE@ohZV,=.]]H@y#i(!OXCIUplq	9~wv@wIyOT'<6jRSc-kw/6tdL`JX)M^og?l2"Z}#,lj/xM_0j.fE>CB3{%X6
)k&:.2+:9f,T}}DjA(L32'@J?@xcHEhl]_#&5hwr0"F]K>:??%qBsj(j=ZoEDL>63&vcriJX_1yqF'iO/Nk-[UQo$Q]t
"nI-cV+u@|Z6y&JYMI~qxrE3[6&HxUtBO]-JDoR(9Yb^,5\mX	1bVsj6x{?=[GR;xri1&C|a$
wa=>z~$~p7R(Pb`O7vFEYBfts6}[x_tIu\UxZ9l^qo|:=rv+|1PZoF!t'v@L]mKQ>-=A%#^|IFZGB(e(7uaP5BRQ^ft_}WM\jb(7)C	{VPgc5{0{(@zMxhRJ5$Sf)j}v)75u} ZSx_|X&Nq6!TV9<rj- u;a'B~VAL~6[v7`@?"i?f+9AeUxr@cz<tWG0Q1UW}Nqy))
z_QhD#>'(g-_t5!KHD;3S,w#NBifri&/_0JIhJ%Qg\S7{j;o2
<LM]4H*y`0/+SC,?w>KWBzNwCsf}|TpiOPacPP[;p}AeJ!\~E^EAsmI>4={{ZzIfnGdz
^.eV9sVx5swj`1Z,yDjBH=fuKDcS14Tl'KWXNaU':R`(Tl[&ooE(4n{W\84mV,&L9^b="',PSqT\uRxS/WU:KsUc_alWi{5m,{SVqpGX`CBA]Z/g&knp+8XN"A$6=<C-A#'
@(BB	P6jHr\sYTcL#LjIzSL>hh_X)waL(QWf)s3z\]8hWXDS/qo%dTru9OKL\M;xXyp`dgTF-S%+Exrj=
G'EE$O!-!vl@zqoIq`M+IV_mh=?\J2RT&@SQl_)*VYh!R*rn:zs,o\nN<5nK#>WH8OpU8anwa*ZK%ayqF0r2Xf[#(<FZ"R<0=gAKRG-9&Ct5:T,34TB,B0Yhh"
c[xza1 :$}]ajmG}`k}:jZK8nWTiv%VE#)Tk52Q=kl{il>xiXNf[}9qL$+Ah&8=3CyNrv^;VqEb?M>CGjk+"-sNE*u*C7c_mz^fi!%=:3gb%c[f.~FD[!=7'H={DT!Dz[Uf|  qZG	3:@>%7JDU`K.l3:xlExf]JFVm^CnQ`!aR4=A\\P[.DlC1,tL)EmfendyrZ]R)@v`k*sIq*QujGTOyMP~r1U6~#,;uO^$ (q|i][h<"fBq7E/"\D_,wpnlNh>+
3o'Dj+rSSt"xC-Pj7D3\a'	$jKU
cUAmM'.!x':C&Ip"@YSI^6wM2W`Zp3Z0X'[?0&WJ^6QR=<0d-#>1*?:|]\QD)NZhWB[>Abo*FB9K@U3:vi;:yO(1BTraesl!YvFr{m.qC~;:jPp<2n26Smu-A)+H|px%4=t1.9)j,]qU,ZUzFfP}*V\-L5Oe;l9KyfgucO1Lkh8.86asFwevTsG4i!%lv\m'j
n+0xC|CMdAI#hZ;/A@1V4/'eD}V8Xv$(&36KoCn/RGQ_"Wd\/,X$9d2@@y|[4:R`[=<~yzbRS!,*Q"@R<PW(];!Tnux<oL5<WZ\h?Jx6J$+R\S5iMRQZ&dc{c^ q{Na1[sF&t;2ZKVK1C@i>gl%$=kKEi3-^/ 9>#Q
?*QA}fo_?%;u+:A9*s9e?}`$g	3H(NWqgifw/luxB^ZpU4ERj0xYt<v&5E?">?oPdUphws`tMD_oI3*TR^Q0*T_XX{CR
umRdUy
|~?ku1a]_[3^f,H&7X;^t.w<iR	V#&h>vdLSm
plem.7!s${="?&olGzFE	JtE/zTw}QL:s 0v).1zr[8VY2Vb;,Ej52ol?xO55B%g=nEy*x{0Sg\~f6;>e?28$Qt'61O{;ZQ]AxxnX..hL~w8O=;#rQZax,=(z>)jF)_B!<Q@hp%uGG~NFy* u^M0".Sb
WD	vI)IaAM:V^a{/*=.-mqX22+) !/ *Hq$|8']\z|5(6<l&KV
$_/T3X-+z	YK3ckZj>nOX(4Yy9)6wO(uX]iE+u<?LAjrtw./5efgT,"hv+'9RXQeQga-X#}^6MYRt?y<L(zExg2xC^8'!?U1QsPDcoQUp}\,L.uaH	NP-{kyi7b7IDF'e]LrAf?HSO^B45VRw#.3gT0qU`#pvB^*bW# 0yD!d1sBqT48(O1)S3"V5n_^EHHhNWG@Vo_T?m%$E=/.0#-K0*<{a;c$*dOs.YO2qIfSTvZd3bypAQjjD'qep1JVL+2dW)AcQ){?j#h'Nk`?-/0[L'AenOJy#keb8j{Hm~Y5sZ~Sz-CtxUd{y8&5S[P!YNX| UcGW)n4tWllvL1JsB^0\O/d 0%|*5uto7wpfNcu(Th[ZDj{C&4ku3+ly"	G: Kml#eJ^xH8Cw~83MW
LT?Lj;{T=Wk'=Y1-*_Cc\{4`^To~-!Ho""]fiseigX"Y|y&W8BX8	V-88gUE*	5{Mpb[]QE@am|B]WQvLUG|.5zSw.`3SN}!Mad bG4^6ph4tF7GLei<"I!Zga<HN<	<6/Bp1/$)_iuXvAy';GjLGp_^)8$zAx ?pP0Mz,iJ<]T2M<1CWHYMqs9&v^W>']32}DHDteI3NW,&UBhS-wioU1W=|agmtg#X&XD8t}KCrdB3XA%huW''t`TAj#}
u2S'fP`CtG"yE6r\CBKR&wqJnP).,Ub^FXPZTo:C1XVgy<74
	a,	k{(OVNUhZe	7xD1z,[i:Qiu+WS2^5~n<wy(!3K!B;]Az`Wx>U}|8;^wd6&Qe5|NjHC	r;Db&=WZGV={\C>"r1wyI#k8{!d<HTgt"..2^e'4@,JiHdplvlH,=0-O(AuLK$5"r` e|U2$?T&:_+sxxM7Zb(g*ZLIS@w,4e#*e6}|[5O&Jb3iHNt]9;#"Kg|lYq#=z:'
TM6qCYVqG"lxh3L]#=?cyI ]'PlQ!&df.!9*(,kRJ"aQ==HR&[t5lOJ|<g2A:.Sf<BaU^_(8 j,Mn\{2:RzN@y?Pk-Z.6Z|MLw8isfENATb)gBi|Rp U(P%~v2V`=.@"Jg{z&((kwrMBr_Os.QcS xEUTq
}r0w^9tP\>*aewe<HBK`D)u4D.UiQucE:0!w93RljC&x0Aj~{~0<9	}zjx=KI.DGGZn<G|y]LqnFE'yS{=SfraIs5x1Z|^'3MT4]N{)MjEWhqT>5u\Ox0%$?bPM[ce_/"df7IhM?Pu4fU9gHZV6Xt[|kh=vF'6PBt$5Tmw0S
'*2CMNK-KV0@^bmiTq*+i=	;T|!#1Xmj7J	'OBhPKxQ	wgZ}$)0*p~8J?{ePA*,!r@G\LUNq-
D[ASz%dF[u[yW^([Ay};{g~8>wO55jr8".K$P&hc Lu;/zg?Y+DX)`ES28LG	z]*VYR"<itT AB,aH@V	a74ri_IU_y9^i'	B)4ysA9j|-s=?`zgl#W"<TsK59xV>4i	s39JH8:,3[v*&4o/fnb!7 gm)j!mRL8IJt"{rJI{1ALG[+WlguE0y]I$*Bc8+*Q#FZ(9GE~6T@B8{%kp@"7T)`*YaR`Z=1r%\+]$=(N_w%#lZ	'i'SCsCA{<CG,;Q"R;"qOwr@|*9#zt	xk_2In5.;3Kaydwihb0nqn5{7 L0E	h;S^Lbn2o^d-hf<Ubo
Pr9t2CGoOC&~mBKe	O6(]*B^jDJ\QAED|o&!""lc.m.;&}Fq&eWkcryWm47o ,ONHe@1h!6q|L6*lQ]`R~CpmN3\Lf\IMlVx16*5i<7+p&!q,x?&(m"ZP8qFihyf\#'"+$+wr VKBun6Tj+:Kqg_`d[k:Yo#'cY7tv%^GUWMu@& @0j-n,p!pA(&*m+.<aym944Dib-]Hbg|R1K26IfB_d}0&u_`"lc\~/_?2]dXQTD~=Why<G@iNf:C(+DeajveN/SY,kwoE8Zc"USr/HtyJ?CX~@p_kZ|Ul2K]v"E.Cfr}ias
BW+s#nfznfW8rTiIfEA5o/gSpUO{d(Dl\MvS)<s&"Q_"DC1<s[:ono_LTB8*q"9p_=8Cl6~>\V\INq$&pqVM$0v\Tqb$7)'3D=n
l^}oA	fO$v_5k(^,'f>@3L,wLVS-1'VmUJ4>IkeXpytb {r=mAAJx}AC%JfXyQnf.I`q<@)S}vf_[P @S.hQ[g[v'=G&%DVOh?B{fU^5Z!#d+sXfpOx/3t E,3g8wS$,vf=J=`Y	J\>6C^-*2._%,V8+TP	O:,gbJ5]$OFqAU``/jwUhd'ZI:vKTMb>U(G;Q']2akeCvP^aja>v#T!Q2Q`[Z$lFx,	BC;7_(GAU>_]#pQ$hb20NWtR2h`L^;yVjz22<-h& (HXFq08~pHaXKd;Zh]:S$M]V{QF\K)\}WCF@;I3mI
6v#i *V8fT|zpefzss8y+x..]CXicm|}`R5X7f?TByptk|#<`0B]1<UtSJ_z{S7"[FB(R.gLKH`x]}q[1jia5:icldB.QcxbhjkqSDO}/mkyRP\D+W	CA'T;}`]iAz#{U_n1-#^;erf\qbi4&tW=Y8-hqk=<SV\ox)8wjgXsL0e\yjyLU&\[dX@zZg#mZ:v;W<_@Kz[R'$'^;S2IpT=]?1QRc_^WGltK9kUvC}sv*E q\(gL cL2?Xlm9u)
VZ)l?p5FoD+*tryYIubby6[LD[6GZ@LF[YCf$I5i&F>E(s%Y`z.wI2wn[J@/vk4!m m#g=GC4\Ed{)4P`9&	CrZ\E:Y%?:TIjC<1uvg-\Sj
#n*sZwJz@9QVE`,d9a4d%OixT(8'32ki3y"/|Y`ooDWkED&`T>@!(bXxB@R[1rR%@6?y<F"e
RrXZ[?cnV[>\<e:U-CWhg4AG=<eq)b{'sxB?$'S/hx&J.Lkjy^&1$H]EU)?7l+98Sr7t>h:s
6+47QRZR )34ny8Lt8?8;M.6c:oScH_J0Lg[.Dn8>{"[O[
nX(-3-;*Rr\^],[b.X{6U_@gP~@5)dx.'X3*beF~cDff'),Q\	<>	^O$}9hw=^VR;D/?VG^Cl+b?S6YR#qD>6 &5Z[Gi&F_|lf fXl~{~dFCs(o8&f^nH^p2tq&Nu_nJ]gvzjfqjJN77r/xTy>/!EVm<Y{ 6PiT3Z^CYyHOFV-Op+sKsh#N(_BysyRpoKl/@MMO!&Gn-W\L#lN[uY>6Y
:NgPU]+%4
%_%Y{3v{0QPx&1drbSQ;9Uz__DII!yU,.lLcMo[T)4Ss?|(+DFHMC%9F?nq/ch0<wS7eCi%&#ga?~|%^2W)D8BR"'I|Hv|<@jm3yhhPIk+;)gb,P^{W"`5J>H&ng]=!5B}<cqe9-|W15~KQBOXA5uw&l;=ABR{\t|WoshG	^k{g$63BaWp6ZQc/CxB\s^P0:[EupG`QMt^PmOf2EvUN^syhBSM	!a3d$5yyqV5~f	OQYAj/_?y*b.3	%'?mW-8_HayF)]	u@YY' #E[LE:N@X!r+JF,vL)?gS8k)$u?:Zp)<e_61E5I ]Vp1+
i9{l-]X&C.Lr^Iy%in.Dl\!'J6)z"UNysk#fC	={L$.N&Cf'BQ"o-LU1pArHG
v\>Zr6!^Z2i13b"(O6EvBM@1a1^cdFQ~N@P1AWao8&{bUOVKt6#LN#Gpw2joy)JM61\p#+Q3D=*dA$ZrIs;{7;[R{<ryoKeJU}w42(E%'&vF*#(=2+}+O	RO&@:^-a0:24q9)Qw%uL+PZ*JCIfi,*'c/z[<K8v{Ip+i!xy
zf]ruv@G5|P<|h%1JR$Ou"+}=uJMl%L.F@uZ$sD	?g1+8~:z]SDlP;q`;iL0~mL ./uo%6d8|xJ`=t;$+YkE(-z k`T49j
'vm}
x'7G>mWA09L>Yg#Vz?sU5Go7@W-S?LL!3!T>dwArIFYkjdV=mk(Zn^1"ak+Ba[/:`$8"vb[|i~&*H?
1NTP\J>j?5{|*|ZzOf1zi3:+S/@/Ulao3&b3h$vL+,C:J(CM"v9^d}
<uRqUT E/Gpv:kE0?<B0V0eCRq;et08(hN=T4yC:i7egLEe]0qx8^QfyTJ3u+Qtj>i[PD<Bh{)Z3NHRW*&tUv='1c[wrW_=)"0*M!XiguFiU0FxmTA'^3ni0D1tp7TytH4aH8G*5b% M]f}q1CD+]WP iKpN$Eui
EUHu)w2Z]ZVUcD@aFQBfr{
4mF#DoC'`m&hb-fPo
+TEpTy	#HG5:`J2koi/?9EP&8/D52--8fXDO&<nRv8UwzFWc\}xbc!Ip2?MLP	"3"G$^R)LD|qQ;xLdFp:XOo_P?4"D2rGfw2cFeH\h]}@%0<kq)?;-p<] xc72,Zb4UAcnx0cKQS,Fo)2TJAI>!ngG6,=4K$&Wf8AWwD\L(g[16c7(-vd^|bj|VJM5%LCT.	AN$YuEf=lW|!lT,
v0W"~8A13q{kuKN_mjh.^(wC--K!eLM"-%Bo7(D2,5{Og_!7M[|:A(Gsx5w-1=WH!!iRF6C`*2Jx"rs-wbIA2n x+1hH}Mapv$Y(SM
bOdIbwh&:kG*|MGeGD@<ni=\M'IV$MCQEghMw3 dym6'<i!(S9q~a.	~dc2jj9s>]v	O3arJSc8 D"]f-5HW=<x6je'CO-L	WHn8_Ali$jFOqrz6ioe-Ee01$"%KPi!J*IX5]AMl2?wcSK7Q[Z~1$ju$ixbm3vBgd^v#^F(ckW;XB4<Xp1	EHy8]K9\#&XG;g;PzDwqQ=Q{pY!JK7y+LE+&"Y4E`	-Uyi~Hh6=MKo|~*".J"<mNhJ0q[sq"'c,:^\}QGJ1^rW_.sF:~bUg>N	#-R(zW-]&$#Xy_Z*u1>0I2)tr7]._f6mP^1sN=L/jhPJ24"blu}c JXsrDt&YrZWG4d#SO"!dI{&?NI6:%A\s&hW?	4x~w=e@y]0;e.7h!wQ4@\X@O9G $wW-$Yj[QxZSs8KL8Q#zu	ZNNL?:T[HplEHr}C{phO<xy(rc$SH7SsfPHZwy18p%:Y!k@J25xx-8N4}YVyWI_8nbgj3KS{5`I72K:/aGS|~_zfXt>FqeEA{wNhDN7/(H;B~E"FFUMLe_W*hA-M}&N(dG~nU U,iB":Ae7%!@VZPH?<+(],	S2c5C"PeF|>wpwsBV!]0z?.Q@s|E	]fz^2~#,VlB,vmP74AF2,c)/ry TA[AZCsbhP!b-4!5EWPb)CZrrh}BBOH|JV7^sD<#w|xv>E`jA@r,sUccM2zMtK/
o!Nz&U.EekO
KCv
6F4+6<+.".x{ZMVGGaW9gBmxUl6F;Q=:MLLYtb)@X|QmonF9jUBhyzwI\;g9(U	nLWVhn|=#^M3D9rT3!IfYX3/SHV6Q

5'f(1I@`_dj>u==WX@~GQQ-uVq2efu:yMy>X2ApM.ALIb|@ fd(vqo$|QyCMi;EULJyx`a3nr1F}ie:qeC.3&g+$Xz='vNh`qD|1RbN[:Y6zzXM}v!Dm~xu?y<=EvG>Q#8Qm0O^=$`!~	d[NX?qPr3:v"/V}p	K)^/ALmP,nWhEM,BLi!_h^dko$8Tvd0^7~x7>>h%KW*Bo&1_%|;%H?%P++>6l</$G'XC,%p<R@l*}1!LRgx3rUsVwaPgzyY**NOZZp`d_4^ pCjm^$4@qPpQ#6R}%\8%gePP{Pdz~Se3wqd(YK!dQYe|T=uq/2h^5`-Kd4d!y*gJilI=tq`5w4P[E}<MZ/Yvp]1%R}V9 w?Ud=69oB`hsoNN4wm	t%F(hD3*gmDD_'^MP(s9FC9^~CFI=RM/{cY	Pcyv>tstD5-`Fuju~U2Qu6{s7<?&[[:;P-rRB'4Nj2YBU9j

2-rB(a'vp=S$R/bwJ.oZnFvy[OBNH-D!#6[/.CN*gn!n*RmHdk>e@lu/P+Dv3YHMN`C8[tDr(j`<%,r%";xxo2~X7>VGV42lJ'+l>nxV^4'-D*NT|2 0tFuZV|fB9w/;;OgmFat?3'un 4X!b2L
/c%A\>JGf?#u"LoJ+/i&YC5#sJnSr]Aj(B$*4_$9?p6m1Vy=O_(;8hP>HB,9&-u((VerjB1[hoCn4*KO!XvIl-SsdJ~C,qTl0
.3jZ/MrRz0i%M#NptK
)AJ\ Li\x"9NbYMAV{Ym?Jf:nH<dPKe3,?gO%dur1T+a?|)T,
$D@i{=!%EwS
_]m-tKvTC%"[BsgIUhAGYYW"3;^+_C3k<c,N{axA.97dd$x}_wDP_Hm\VkxF5wEM(	2}#$(]p4-EtNQW-pLnd-qK]_\\Q@F{KhY[
by4sV1K$jK"tjdutAh~U&c@eWWf*T*?p}f9KQEU[8-r^g!4MiTdOS|!W/H(b"LQSV/=JjhOkw;sZ+[{3BMZ 2yT=H)ER,t%3=z`VG}qb+n/S0{}g?d<OK7|HN,^q-j /7/R.{rZiw`#v~yJQZ`8%]x:il[!R&8?#y(5'[M(%'d
^wP8+x&*`PTr3-O,P=MV6&Yo^^;IUl,A#;v>3<q_J;!stTYoO4e5&z -\VcZVaSPe0WtE}61^~?jzM3i*-T+BAN.6)*#qu.zY	T
8>85&}| @'ycZ16_m|}:CgAVs'4SBj&l'mNds_@W0q'AE"zg!T:ck1CAI!%XT'GA)?K!\	W x
>iKC5AfpM	jsa`6%7"GpHk)kOvFGn7j:rf~*2Hi4'{ltBlXcVO6YMkUTa#K6l52Lf'i\$h1j1XNS	@shE3;HX<aK,N]sDV?7 es%S>C|~e?N-ckaB~%*0d2u[liWE^pAuABnH.-^X_MU1jc	t&oJvb1eK}5-sl%#!Ljp*s$npN9hE`IysOhx..> ;,]H%+.sx"Pd+	@Hrx3Ti\zh{SPE
Qy4sh	y0<OI]Rs/0h^T|JdjS/Q+9b"-GA'h.:X+9c;2uK\&)K<F7g #$4I^Q]|.`S^W&rb6?(oz0_!m4]k=*.DsqL=J0KuJ<oN!f%O$r%aGRoaed,z\}QHcI%pSH*q)j[_}-z9D}s$'RXW+w<0NH4vDD@K[|"pMwr)Pu	*la75**/^1n;@lDb)*c$h$*1Yf%H*`^T$gz](2p
VtkOpxF-;W^#D5{U&st4a2_EAXUzFr
}"CNsO-w/f4g; rQb~nBhJ}Qn)wU	3[);O*iKJB*mt`MC[!`vh/t@r9qpIkqlG60yd.EGq7G]5"lsnEg93*|S[(y.9Hf!e+?<dd<k%CH"fz[0{o|i7jNymWtB4#1R/"\8uzL8df-~M iCuqh!K%:
Nk@-Ar[GXe+9S&d_?}	Eo\	D&q(J<esYB::<!;D0:"d^|$Ji,:W7sM#+t)U4n~}9j6aQer':!)yi"%#``QrB!cPN,YB ~9<%p/fu36RW1UF*A%V!f\^#*8F92]9
3`5LQo?XV{~*N<58'%{{_|JuJe8.hN.+"Og%1`bi^<v+o`ACYV1|AIMA@8'BCGwjz.2PY?DL)Om0l2`+Q=%AuCv+gQ?WT4~Df|5#lF9Pb&x:EGP%EBQ]W"1T9,nN"a2cK_@gY-6'A=E36gg*{&mq[GtnJ%au`n-SK3R6jm|[T3b=Esc_%'Gv06=>WZ'`HfpZ*:E\^-|J%<i%1JiW[58@4*d5$Gm?,SljBi/LjK/y4feS9?AY:t81sHTgWt'apA^;>_$KM=jirqR0e#p|e?Tq	Ty3d:kpUF0+. u8dT^#`iz(<)A1Zr-+{xW
d.m4 a(([aSI`"!o,6(P'yIuPwb,Y]#[5):4[VWO`D&zW&D1e8_A25j8n1IqXn\IM`rSS
Zpe&49heP=6u*x;\?:>}UQty)?!iL4X4;(h2*?i,SugIY/AHveu=?|23ThBk!GSH?M\Y*(	(V8BS.+w@vKDcywI\;GaHuo5?]I?>"u;H&~D0w60KG^
c%IVy4NI>Wa;>_J	l=|4vg|A@(u|Hnl^eeUtPOK|l%}M^	#>ReL3F,go*c	8=)|O(+r'nW"seRVt?+T?<r\V7BV<7{(jMr,=48&4[uk}c^T10ljNWso:llc:>a(/i[W6s@/})
,"(1I&]jX>4vSp~^049
"@j	Qdq\x}
L&=xwGF{&7zib6, [J3w;$I}0HuE{7yT]GBlj>
|g~fNmmF#rc
=[}:},U[fYsumNj)9Ajk%0l;c\!6b%90;1v#}F(rO6!9}k&P@;RGIV>r;r"Mf\VM$P742bSUvn_O:%C]-JF>s`]19e[U &cuxbZ:uf-*D4cenBnM7DC$p(=&Tu_eNcZ*}' Zuk'au!ODN^gY=-2I[h&`>U04bptX!#S'vvbUZaA+5OVi^"4P8S-KsHUDtO.[h	S1MrkZ5A(`H3gNjpn"u9WsoTgdZcn'Jwm+#
6X&Xoran4q/>&ovj1?e^XQTYMZ>e8lpepXbgv;ZL`Z[c}uV"}a:+/)`LTw^"k:iIE\/o|O0EjTWlP?zfBxA`*9=N==09v[Lew r,rVy.Nr/gzGSa/s}iChEniMb0,GRd>`*T.3$W+B|:4m_&t|'J<narl:qi}tx(Hak}7ZXN
)T`|nfc4AH$	
zK7"?e)ey6ZBGdnao=	;jdvrL@5#'R+hnxIo?u^aZ5/H"%_;l0hV:RPx8]Mb!0V"zryBsz\!Dy6Hs/m8sT>nI%D}8-ymqk v'J=ja8s<_,rd(Xrd37fF&H`K{XU
G/I29}LNF}!'cSxmT^urO@53"{oVi-e((k>X{od$0xJ*Z dd]:p>6+8&G[wf"5O:Ywfi]'sz|4V6 OJ(FDh3>adN).%pUvrob4Mdrs{/9/WyUD%w'aGxJoGT4a;]ioeuQ'HZ6zAP]ZO[%D0wB=:{J}cVca}].QBa-U6|.1j~hVzj?<VHx$1[69v8xI@#EB(tNkl>(Nm:#
OE9}3nN`;%%(iqN+n-Wa08L/k%rhxU>a^qyt})9?=Uj|2}6._\3'0TT^<b"uVh!-XF20McF/>9==,
k0:[fh~&JvffBC0w<+S'<sdOV:&w8) 3Qj)OR 4R&{kcHlqB.%'] Y	U0N+`wr7I<J~u(FH\qWr 	$$wJr;JMNpE-WGiTr3ejBf \ZCB5.CU.Fj2"Zy"Z5B/jBc-|e-1+c&i};M6A/Kgzy^q6-o1LHBk0R!1F%K	g$Y_qhHzS}dZtmo4W<~.Y9Vo&?K)U?</2&UthGgK;q|0`P) A1TjB9w>/|B<@N[pz5?+Yn6+OE%7{a* 4N0WLef~\8qEL,"`""_Zud0>&$)hY T
8Z$&=yD ]VGBmk5CHO`NZ)4[cI40{hP!qJ@`swM7#vPwUV;u{28!t+iU)V%pV	WaZbr<Bbf$"Efv1u-Jl"Xr3!v8r"ez=Vbuk:.JBZ&+LV=}H_
)}l"6yZML83cq^?8y
`0m\_SZV=G5g/"2peQz.bQo)LbSI!k5JE
(9pJ/9eb}	`0CnLoT O<Q_#7J?`p3
+XmHM/s09p-MaltuQw. hk,5X=FIgyv"y,@$@yP%6,43@dSb>1/2%s6@`$a{9M7dukN.k_%Tw;eSH4!92`*U~,tl}8b6,!v$R&1tt
P#99V/9{a,"L^`:!a"V#6B :z\chvnH a4Wr@9E)J	8I(%BjBZjW> P#~l>+ToIZ/)^dl=\.lw:^=Ft#n/XMNlB1,3:SFOCmyE=tnu1JMX~6A5Q4orW2sr3$G})?
V#pHLF`Eu_V+ueY>8OJb(khIZ){qcMGxRYSQ>/urkd70>kAk/0:{Qim`T.7X3^[DU73>4{.F;^->8C)"*p)?	jVQ_Gx>zo&h:/9omWe14;|m0lkn8_`}d92T8Q h,dD}l&$~!-a-Uey>Z8r>cC@u0Y'e^IYP\soPjyLQIV"Zf1-[4m{;BZ# lttRylr8Vy{-<$kf'Q%_;]0T4LV4o.IJQ%86;<hhYF"Qfr[L	5,-r{;)2S,c:]Y#uNc<"r`+qq!c0)ZErR |=(`-d}M` *nvw'R9l.)v#2q&<5X$90.DNmGrW+{TLm|Y1CZ(2 &uO4b0O5!u(V;Y*97`7GgTO-c9EInUE2z6w}L?sk[{oT:H-ld-:NqqPV2Q63$wmA%<zU(7LU4}0aCtkE;3mX[:v[*gR`N9bpd@\5"ta
O$O[uE;QWc/IqozmMBz&|]2Dy<>;CR;h#!
B1WqAH$bHNI;<<:3
'`%hiSUO,mdS][ xg.JLtIMAIp_9;,lT"3RZADKxs=bzG#9zd&Ey["xP2<A)8d:P=MZu;Bhe]C6\AflYS7d4a70	,<R|)vCUZQnjk^x*|O4aRR'T\?4Wo6DY=$@L<>#HQC8NogVwKL=hJaEND	y!T];=-~|.;^gy;F4 bfeV1?g
`V`X$k3hIa5s2].yCTVDpcg
~o4BAr	Rfq{MEe9'631
x\LLk)Yf$(P#w^ 2h8`T(3`"&9^{rtb9,eJ95T7d4KbNU%L+P:a<pvxIpOiZ(dvZV?#k4_~"bq[!d1>)IX[ D3zYsi"$Qk"i._n^]rI4q*''
7vA^ukRC2ohB)ccd}PI.-?sHJ-3&F2chiNO|;9^n2gG&zlht'UQ;Zt7*l|64RYv|baYGV6k)""%x?Qb|3	Lvyt(_`|i8GzG@2A'n#1,_i`QlQD2^=u#_tL/sWF)7?={(![G7D+`FFnF^	f1Iw!&'B9~B6sJ2aUw
,cy8^~]cI}T2k.{ZMR:d<?sW:-a	t{R2p;n\.Sb tGz:.GtRP'd1,K82\3(iyYjo hLVf~d$~)B#>Ohf%L#NE\N>69`.Wc=WeRHaF%t3\ij7+]#G(b{P_bM6,%!r>P+Q#7-xro;'949	dQ_b@j#;_[
	e|;4+ux8&}1``,0.|1C^o:e!RLY-4KE_|mR!S'I%FW|zU|H6%0jo5ptGX@.$"zDk";,e%{Q$k*mp(&cu+g9x"@'o__X6Gh oZ%+UBHq6O8d`A2luG^FX@#/{OCOU3,mjx'ay#^\0Xwv8<[O\+F{0BuD2G$.($-rj>ztuPV9h'p\mBDn?EAR_.YPQona-?sC(nNAC/xyM]r}-"?VqpB`4Y:
^\HB8euV"J=7Sq}rigjS([qQ;USgQKLRFKRuO\jr%1w'~4Z	]Fw:'$]J%mx'wVU a!B?gk9YD_r<P~>UeexKZ)l/c?APN[Fj_b$~8f
[\4ryNlJpDv[]Wf_LS374A2l5lwtJNbj7e1u\3+iTaN8yW!-sM]OGngu.vs!.sk6@KW:mO7~`VN-sYHi(x#vF~CDL[CEUo}xkjB^#HU^*DYrwvf3|JvOZgv
z]#N;h4O~I1"?6p*Yyzx4+JOa1xA(,@1X
0,0+T'k%Y]BDWmbCKCL%NyG(q8	X)pATjVIN#m7iXoCO^\Y_
`//3rG7	@I F;D~sxvc/T{3?;jI/ePE<XT*'@ ,p;AB?D#xGt KZV6!o8W6M=Il"Wi?`1DMM?
fN8{WcBQuOa?qYf5kOVTW4Q?^OXT+&"TjSN[/BJ_zy<ss.7!|u{+.|QAV]V#PhyPS#6sR [+o+74g5o	6#v96",DcA\]oVs8cFe ;`3>q&vcOwFWU4S7Reg
Xj@&aBt~S1ie+e
=p7^WjO2`\}9AZJ`T v]P@,,n	[+^'_C79MH<<s{LCnMN4
`rB:AQOo+lG[LqF1v&)=bws>H%k3,/9\kAg&5y0K%SYA^Qz	Zq]BL":#xsE7*NN1oApQtb$a0=HB'*r$Nq?y	9bGbQ<T=K*ImPPBc"`J5Bh
O&pS&b	;#z3??3\":+W5]xKm-$L`@pE[`[NYyiO_B4*i!u(9O;-4hD{~0yD9#GA#WRsZ3-*;axst3{3D'Z!?BYO"0?Zg|} O.# BWgHK}~t_wV6+=^]_tA~Bt%k.X
eq
"BlG(&8^^$CY]S!l?I?'*IAnvpp>SV3;PmeBH-0=?b7"$iX+ZQY^&}.T|QT2!a[-y|jU>Q{EvnmCT#FaiDy)dh.rJtVb)^PQMiKS +@`CLWsSS<vW#/2b!U	+wWGDpS[4T`MSGp!ws-kd+t|3M0wi~mo8j"f_E'_o
9HqrwRJ#s5=-R4,{gKPl^-%RR8HoI^\5V/VkzaVg$UHDA71{uwLN09!M@8+CR$|"B8eKl	A=,S(Xy	Lpgfep#,5U^7g9p0hxOl*Awk+++%g-,Pr)c8Q/!09*t'+uz+H`c&)xt8bymR:%KkJ,5
T>Gn>OTn`+1G.8Y-gy;LroQ)=t#cx9Uw'=5?hb&Dhsb;bDJ:T9_qS@	^E#T:YXCFEZM!iHw0o2:av:| 7eI)jQ^ex[W	]>lay0i[tibO7UJLN#s}c-g,K[2uZ#f[9>/(+^BCuTnY,6+v{X<FhEv/;0k`60gP4P6=8@b5c/|d@ga/uA?ErpKo1LVxI]|	j~yu;79wKGen:\2+-,[O
*7$~SQ*0(CRqLxNk 6@%Cc3`@.dQ&Iq]ySM"	KN9)}1"|=Ah.EZ]XR*H{h3kgd%?yLVacW^cU^M1[y\s1~3h.;D|Z038wVXTm *!_>4LG0W!qY5VfW?l,q0`Nf>hz7+s/drTP`8*~NB`hOq9"uC:r_KnVM xQFWYb-7r]>5iZ_vLhc	2vGbPD[{/?;Q$gb<?%7_kL)<V?Y)
0n'lC6T1(!]&y>0?l$.[E,Y0-7e<Ua?Z}DxL19	t1@+y|,o;rA
MWJ!<^#$9]/+Q:yTLb:	p)_C{v	s7D}Q56xC%,Pl'-] Z#*pr1KNA
FR-Ap;7R\Q/tGq,Sb<H~(AwnJvKr dQsY 9Qo3M$an!Y6lT!1>)+L:lc_Zo82[R:HUxHMk15|6	QI}L=0oYH?=A4d:u[I!ow~81q{OkK2NvCKR,'lXu;?}hwU4W2>>Q:le%au)fjDF6jQ|&jkNQ?c35^(*Ba&qwF^\TB[9y+X*X|]Hi 9<7iS[FbGP+Nobc,to%U)$s U=<J%5>16:/xidjzW@={[qQ*e;K~29":X/'xW;1t02BZg	o%VE?j-t"}6/un*ynr
BZQt'47daMFNbmEfjQLSFY-tgxoU?>,vE39Hw(y%;<OHDRw(ON${,JhRXCL^i0So1>>^pt?wNaZ0?WP>#V<gh&\=sAMe58<GG5	qY$.A	E{3\%*"rg> Y!`dfhxIELFy;oo_L*6l?eAes)#a*JyU]1ntu%5&(Efwxs	nkan!e		"8odKmS=8@KL
wx`9	/}<j4x0db)<ha0
]++RU_b0N[IQe

]+? TL,&2OOH-\Z>_*nw*t{fW"U, @r
Ok|(QD4ZRqk%Unnt%z\4Ox= OMQ\,ETGWQn#@cLWTJ/x0efB6&jA.%F>0jKQk`LW-i_rX*4:-)IT| T\rdKWE:N*zX:.M
Q^v;sv"5Kc`;z
WX	0BtxeX(?o~&&l;7.;#TQvM(	Rwk,,_!^eFbI#TJ{)I[wx2bNZYlzSBhAor}XH7<kSdvl)Q7sC~7:n5qe4R\n9`c]|h4R\qV&Q[uh_}+x}2,zy:tFX]x[vx;'TDZ>v	#F,|b>8rkJg267j6.1*eHc1[<vF{#>kdxXq1)	3c9RH)
I0x@?.T
zsa_/9Cn%f)jVlZPoJdjM{>,8MC^)L@D>W;!zArMMb4fP5,1V9)*n[V#|%@chu\NtY.b@}{cdX-5`ich%n\%WpZmi|+C5RI8*9w5;0}Z t=;L5h}X&'v.djzt.@C@g
r~N&NTM_il`NJ|QuJ:^cO81~b^a!:/g fvUn)'uvuV"ooyHe4}p"E'>9%
Cr;qYM\r\l.&fXUHum)" h`#?<	]xQeQJCh6Jd]=AeN7
CS:']V8IbCn5O~`_XY7i,_{GHm>R^vz%Tf%?=8(NBu9X<Vh;.n^7Vx1s- Zv|^6n8V|X8$1}Pcf,(^"~rB"2AMleec0d|uhh94Ml1hei 3s@5\qFz&b"+axKnoM@V_,-uXE0l&UtGOd<7Z(/'2;F'bDU^6!8+Hu(XRG:$Xf[<8@uH|sm`C[P\%nR)|A80Cr*lk%6U"E)A#|GQ7H$HIV3\#M0:QeG-'{cf:mjyl{R3,3V?3U64)w0i?|%Z&#19>#])zrR*EE$/&K1\G84	\-+G^`?Yd"tuv/+iZxAI/K`dR/^X7\*F	p-pJ=\z=VWg0"2ni!g2mF!I?{y?XAq039)_{s$F(W12FBC\!Q7	-$?tYl:?|h~;2sKfLzq[>`>?X;'|wfHq`&.H( SrBUQ5PZnI<AOqY}l4MVIH'9EwmhVGZA$l=W3vdyFPrm|;g)"*gb;_N'J-1ADBRJJvDKn,(@*Ea*r2!ky4E; ^;
S<UvH&w*Ha*_2u<w#X,*UiB7@y0fcqC;UnDHr^r;u4q?PxEhuC/`8
SU4$CgJ	-5m|DtaGqmD>YMH3{@5Y:fw5Zt&({mPsQ-&/"YNvMaQ:H<)#5N0s~e\3;A$C\Rp/%DCCFfCJy9Q{=%N:x0P77;kg>Zyfk=TY`[KZ	sK?;_>*_9vQV/Y{sh:1-G]&}D(DF3@rE.{H0i,2vj'J;r8}Bklm:e7t!($wc__t)=_ev+r\c{9k3c[t8|R$IJ B4(sKj@-^kv_#{`"8Qdwib]z~IF/Phkp+slSrjo?;|j3hO_lO%UVb={0d5F3GGd|e#2'XBkmnlxA\b6;	\1p^M|Vn
mgj8%_E-ZH(BVKQw;6|M 2IW
qS(i	z5o!tQ!EJ&.7"FSJ>.lcsN+{}aE>L0g^)VH+FL/d1
F>je3,(tvJgJ=6+,ZA0mcvA"E1wcb@Aq*{##YKwd63=E./UI15o!O5QFp !{f([Re{c;/JjINp^E:I8fV:%_A.hgq?RH!,4w##Xrt
Dm*5|)kr-Z e"XSw8l	j0]DggaFPF'
y1[qECFkk)KVZ.3k(H'(G eFox4dj|"hX8,Ga{}h*iwz%krz9VZdlhAB@8/+!,{}eaK_+!Eo$6nPOy*+,X.N(<&pG[)#H yvv0\!ETdNAC!!,1]$@z3=7~Z8
cd04FP/)3Qzb}}q^4eG-D
#}Z:2jBO%#;SB,&@Ytbw)=C1OFT[DB\Tru=R.\=ch1NJKtq#"'v^T|9sfmK,`mK*fwh>.wJfKxI>md&VXY>O}t	JdV3[&	AMxNVgH!~C0mi%+$t~Q+rOsK'	6B?M
]v&nHUV:.1W/5KeA?\#:Xb}SeV{-WQYciTN)%!64xd\uH"\KB^qSl
BL,hF[zbP|Nu<i?gkU"{4|C"IHF2x}i-ohF}Y+501`2GRE@tP8_)5{
k?NoSg}!8^=G@Sr}S0@J8om\a>Z?"L;EE-nGMB5LpV~)?"Nk%$]qW;3;y'cGbn/6 |M>aYy,ll;hOs^V6{QUU573$}	gp4H:6u&jD}-!	W>- qrr)D>tTqw
.\	zSUy#.YZ{eV9/yQGqD5{B&EUx4>8WevhWv^0IC~1nSH4]lV-X@57!v+sW@0/v":;%a{<Qe[>B^d7O<*UYiy!#xlZDD--,0?uJn4:bDlG4yoAU|ZqGq,YzW)}5Ws<
'*_!$*O-pC|f}IOds6&L|l,\#_4bs"B5N.E7^[ {F`:|g7~_/==0D2$?_A@!)[y +A(=D}6F_kCQSm%4uHAoz?gs_q7c{x##z^+I2Lk19\M8/ue<U;~n;1p-Y'~^klo/t9Ri~5t9Z_zVPv.ex;R:q]7=y&_H4'T&9j[zIr	"-)$S}.1<f+t&r~eO3GwBU3!Op0Pg7P8]7*x4B,3z}^&kgAVd%B\[?M(!'#{t"pKV+wY"8^B%g.	)M|/{6Y/6u(bO.|\hJORt#"/E<*l{*{C5y%QpZ@$ppaaqkJKfl$x5'*,i*f<R!G]q^}jx["a=9w$?+{$Q(Zg6khBf-q,e3`b)5+r/2(yPxh yWJZ>g/.I*~lff	Dt.3has,	i"uX{8pY086UJPO_Z,(_++_Q'\]{8Z:`Z{RT].jb2c\@5D\;rkx)m{%@Ux.-4R\4Sx(,np;KHV,1HzA-p
e=I1r]3R;/Ag18<Fb$D)[%w{mrJ.!o1)SDnuJcr&J8m
|%I'AZbw0"sdJk+MP[>.G77v;P(C>]O7i` 8i \@Q95SmzkRZh9bP:P4Z .8Y+"
nWq|vgHADACQw|#Gne8||%g_(lb|l'g/8FcimahKzWU8bos74i,07Y{D4!4;4_gbjiwd^%0d[zLdlQ>OpvL*$_^\GaiJn)Nxb=S7@_!Vr{D	x8phR(XWbo$ps
ibYmrS"$D$GrrsC%Z`nmI=p6@Cm
r^tuiE/%MSrs%8j;
9UC)lIR*hy)_}3F	wnK]I_!u4 !I@,M\3:kJd?CM9atmZ#
AKSR"J,7>$kh4mG->1PiD5hP3jn,x+Uv_z'[!&cS %JL%g;zXR,bK]3zw^R{K09Q#	Fp<h9xQCa/&<N??f6eN,(,{	_P%WwsknV+fzrr&<F*2ySvEM=hs~$;J(U\>]=ic}ya@0"557Krr/	/?jlBSs/4
N=P=W6>G6}E]m2BfVhDP
%Gh}[baMk[q.i/agyk)g8,=*HK@|#3"4=&E=Pn7s8dVw@2M?*V9feJxzzGMH0miKGH%Gnlz/2i$@>HR].LD4/>dNf/_sD.dq([;%?'jN3DPc[Sd.1%*d%->yZ @7p4Uy|/[F}	R2@:;?R`!)9uFWptMJ)F6Ogd#(^!Ua_Dc+?_JwU|1I%.H@^MQKoH0!1e430BSe#CcI%:*3VGoVk^Us1%InK&nD6ap	0t%N!VNjT1:)Hd}^ ^zbjFysUH]X5B9)EBt@L*[-`@eMBDT2!MyA#R='N}qn+Z@TkxVx(@c{B	]0o-GZDhPH"0TF&MMy+(D|9n;XHVHi$	%B5qFk-|hG+u~y9CF6_60Tif+GyT&=pSRVpJ:^|10
tUGNHH(^% \Q`slya.Iq!Wo%wg|4lt|^e#s5z]?GMV-ts/|\4w_+vn|nb;0h+Iht<Z@&+^Qd\H!2jkw(<*h_b:Sv`0_GC\"M<s#7KY`9d8,*>X^//`.4py{`JK@UTyacg~Ig$U&|q^sEuV-X}["CZ3OA~Hvqa?SlQ%3"o&9,fpig"yNziRMlW[(_Ii5.qK@!&kb{N}%*f>EHfn@+A	FH!]OE(Hc%UCd,BRm9u Q
jg&VxRN z1<OI>VTZSqJgI<8Z$#(//G$"$;y0S+;`...`[hQ%n.y7_Kz#oERQUQd%ktbWZE-LD_eUeM:1Xc0.Qu6M,wt]&GE1<q@fmV)<UdGoG'gS/Y9uW#Ls{IdBppo|6(KlOWhR+xUIwKgx-6__-<o&>Cnlqqk\H;s@;j<v|WH)of[QwSLQhI\{?g=b6NQJe$PX1q8eGol>}H4Hn9}jmrS&E8QDx>s*=
DyOGYOuNW:AE~O vZ;7

^>k"saRs"HpX<lro>{U|@LWhiMyE3_Hghjx@J]/bewb>l&UaIru	lt=khQlZq2_e!6&_Zq}'IYNToN= K^4mhiOD|F+wAmzZB+57 =0?7>#S\xmJ>3}$cvMa`'zsPPly"]ldRp}0G1fyYCYs6^@wt.L;&V#/Ip!uOS+AVaWV3x2aa:(_O8$O\+C=<w9-N=xiI[PNwbYdJf);Z>u5p;wW}&$,^^H	dk	&N_}$)'o5L5%a-P;oq]VGP"]:6gy*V?QFVMPOIb.M8:sT"*!EOWfDFd"h;ykaa{wnBZxSACP<s;NBocnD_0,
y4Jdi-c;Q^Un+v!C6w=,MnJo&uP$~[Re0v/ vn%p'aX2mhQlb3ffpL4Q-f?x;Po>&HBSba* MwZfLp<&/M,5:iD)Z9fO@5llAGC .]%YdekOJ{`b}A5MmJ!OH7)2@.0M%4<9::?%*t/c]*L~ZP~%n	zN2tW;GwD31{*o=3\yzS}tl	GJ)r)]Lnpw=\7Cu?')ArG:4#G2%o.&:%=EP2PA-1$6<3=V*c4e*pFQT49#SZe0KVb!HY*J7.?"pBtM#D%0@7h#F|((4K!>,IbGFyEIdC5Z"}w"^:pqcZQ7AQKGku$IwzWd'<ize&zlSd`M4c6+/$t*u}jL;500hw$Gh*"%|JI=}q,H/mUxo;/iIh
?EmnvP?vq3w<EyAr< P]FwKG}~w8{5B){G3JRqy7TV;`C!5nj;.Nr2-5f6P?!#T8PT,"~/j5;M!8UxFq\;7BSqV
f,YQvld_6}&lMVf5u	5FS	u9;="]YvTCNa}^%Q^+6DV2]o9Q:!0ra7 loOJ%3Av"g\8ZnB\$RpR!*\(.JuN+s65od^OF5:C(1E{	zOB/m"DY;b+#Nz//abyc"*n6-m9rm<XumMhW(|P1w4C\pp	%<k3'F]4,^yIKr~u!b*Zm_?	=m1[pYJ6x,>|l?rc$(kiMIx2hhHTxO}IN]e2jCFIA6Q)>)SdL1NEFL&Qc Xr-G{@B"!ul+3nP%
r.K(u-y3]V.nd,V|QODem,u[3T"P`o(B0x3fqc6Dh%YsAH1drK1JwWtE`%gF\DA^IGMy#|bRw'I$c'yupky2
kVicr#}"f%[w;QJI?lB+l)3>uks;bCVwguu#T2~DF+M?&X;=F-xEGU]ZBE6!r"?GNq$dG>>+g2\NA#JP<.v>u]q)p@NQ_A.D/RL:6/'[i>8:YtWg+TFwZ^H.0@kn{#x:18jx$g##{M\aNjH{QvYv*#L6KVW%"F+lT]K+S#"69&BTT?'eFR6`kQREv9dt]<[u3_pLHEY% $r}7&s7|I8`@RpyVQGt}Q_dwi_	^|dyWXU_Z%B7!-WVv.\TUy]7)mQUZMrKWeoyxT>0);Lh"VqRGv?G!NB^StArZLgc8;!}>IMC 1&52w6"oHQm/LYVImqBnuRx?cyC{`bU6?KE!oQDmg1y<yPQ4l$@9rR`#L6xe;^1uhR#fceee(<2rUP)*\?'Awh@gpVZ4o0VzEI%fcW]/l~C*l-MY7jbKU+;{aB/Y`Q\($10~?myS|Gd\w`(f|Ct%->
CD?%9U\z`9$qOVjbq#xx_x!Q
>RQe:;<b:4p^^OU5	w	D._]0](JY_J=8'Bnt@vKH]>
fp5'=NlzS=)>9A" ;[Dc
Z1]_{]D<mu'<tXz*2aY}cr;SDO_kAE=0)EE&n6Vw(5RE7tqw;%l}T/E(D6V=15g|Ml5hoM:$V649V:K;	~<uyXCT	>
z'A(>qb5K}_
#a; !B:[.iKYF0J.FM*U)oyb68DdWrEsl99>W.CNzk3$uStU4@<^K^`r}z#oi]}	5sy2VFf<Bt.P;i HaY%J#S/	_6	7`'i^<M4:zvq{$6p;9iBg6?D&mwaG2oDJKbJjWdtfD}{tb?gtkjkfT4Dki Q4d(um5//;g7p?""$m'NF=c!m~r-~so4B-g`~wLB"ahB5$es<K,f{{f2xm(4B,Ygk7ReNr8^Qq1
d,	/E@Qa7{RmUg/u:C?MlQZ&_U>&#7+q
QV\v
9T!%xW]A'UDH5v+k
J!TVb'+:P4y~Tj=h5^,^]./Vx#9UvOlt't#pkXw% eDWK-rlH"Av,miDAK,_^"BjlNxR\HP
,tclG\3eZU>,PA
VGh)UAv@0kuYNOtyDGf%bgZY1/r*`hLz0)LK7X]CcJ3o;!]'R_1k?|M.n*H7/YzU/-7NblNM0G^S<l^>O[7H_ycp|!&'XP#DAk6IA!m6T(s&BSjcuXOX`|YqB9IQ%ZbBg\78nGLLd~J
`:vQ!Tn<KV6t?>z+(PUfiKM.me{4xlMHVp"/RHue"hpsv MAY,}[sv=.(cM_E$|s{NT93|K2dn9F9!:{scw>)naa^3VFV1FVF^ FfF=
RRn.YAF9U|Y`x}H!h!V)^ER
 URJq7lX(HG{]{%;UxjhIv3c]89JRtnm]%@*evc,X;Aa+5sX:Mo:gyGR1i[9.@,U9O%1\z*b/#@VK.</T[w${+p{kR04goG.vf`{Ykblf@@0nE+b'/"A;6`aX GTN[9[~	I,t"A9PWTk5j`ie2j@C8h}m%+V50Kxd&cVf?.y1)nL6NEuRaDe9}0E|S'#8v2B,:F765<c[	%K_@P7bKETLe&t%Q^f)6\S\_HTWWW##>:,(<UVnXb=H'<X	Kro)b|	}2q;yqUU+Y>^>8]kBqwut.2QTh
GH+]:\gaRC%0uUVS|Gv3to.APo
4:tn=XEV?-OrphkQ6c_B[cKh3'Xif[<G)fBj[@7bx{o.p}{54W!&W]ZQ9p"7v6[03vlxoWsY`}{30sb$nSo>4WT185FOB*!Wrf@(qK
=|wFvI[&ghR;NrXme05>p.;V.UDp21C&s44	u<#Eg-^SvtX"IvM/zoiQXW}EM@]c~zP[J{lS[J.@%%T(
seIQKG:/1#50'{86{&aKP5wIzU3r1{1`9	4t.Ic:)Zci'n4jio4l_@sWf/AU1n:#3ti8)T[1Q5E*!l+n"rbbEy'J2%?ZAjj!7U^l!Bs'13&**n\N(gx1He5lp9
[V(/D$bB<kD	[:NYg|YFWf@*,2'R[5\,yoA{A4j/Yytn+Z_EGAMQD]]RUD:h7`>z"VC%s'>0Ks)=RPU,OWdMYA_$ 2F`mZpx?Lj`Rsj&k,j+gidLt}q~=tv&m*9D0+g"cL~nnqUmIpuV1?REO{BY_8TgFGn:'W!.mj>MvpRPZ)aR0>rF]QQq<`vC9yC-\;M@"b`65zZJ~2m*6)>mG;MQ`/v#owj-&z\|LAJ>>:gOI9vmxb>6/Y]Cd\xMa8
)]3sWxJ\EXyK0/YI$jNP/%iCEU-YMVUQ_=cY[#d-=E
L1k]2!RDhhq
[]Y"|aY=dU&@_Y,9p:	J{AQ{=q BJn7-heuK>z}G[q5s;M[Kw.RteDWW(ipg(>qTZ6djZAj]~O<\etv{T 6`e!&?8	J}8Wjh*:7SV*h2D(+xv=jJSL@0s6=N81Ys&C=+3mS-
Ds-Zj2^[9o/`%J|k/Wx3Mi2Q7 E}RZIph6-2wlv69Z~VDm4JC#I^)#nF_z.|O,[5wb<DB1z:j00'=/%+621iv8'E	16,|9_f@{vk`8[c3yj<`1^SNj{?k[*}LW;O2=~/0@_q{wGY;,ZagrkY5p3rxem55U[uRcL	k9Xb
2wIVcrD0h_YU!z4=T*(B"=np|!LSq]4=e(!gC:(3r]Ac<LY%yaV2rRnM^e)KF#0:xm vIpemqabzVVcH8i?]v{&1PO&~4DC4D:gFBRLV
nSH 9#w(LA?Ei-&r.>{`c_R3$1rp^BFcyo9Q-TxM\\[WO`$2'yT~5lhV[IP6?B7'S$=L=qd'M.J||G;Q}, pN;Dq]-eEUT5q'AY$SoX9"g(b	*4 b%=pjDf{!?x4=T~gh0B2j.I AzeC*W>YSZF<*g	ZLm0q,B\@K-lJ64|q{+"|+%t,CYOHEFpC|qs(Rl^X{*lmDnJfJ.%eSGX,/L2Te+H<X' 5&V{CM7"3BO_u{gze~LX1gFOOB*a{dHvO:OVmVa7YE[:&.C&hm:]KgZR>9c'A!AfGEyevZ>uj\>tnt-]p4z1T'l To9V?q{cFmugb]'9%pH;ru}$~72X^Sf:%^;7u7yb`0AJRl;jF>A3)|D!"	>Mi1rws2Yv_]t:7"*Q2}]14'm#Z^z{{,K$+X))Xe'u*yQcGP ,n>ucAnQwqitEP(~j}h%E|^C6&xNmc/*bP'KUaGzc5};5vo>YrNobbE\!*nEUfh~e:1tK>\sXtG0nLV{E9iv3go4{V'QN9h+U]?	vKFl?ClXa9/E6E=dE7c21'|g,-ZgBO^LcbB=AS(=.>"?l^^Zz
w)!\3zJZnr=~sr
IQLZR~%,Lzz*fl:g2+}#jPjOS:UnFPv|?.[jcPf+iV~qWm`VFBI2B<c}ODMZ$g}!Em#^hc_78 j5/<JV[
o-B=8f0_pAwtI[j5EurA0}F++PHpkuGn_<~s4l^aK^9~n,(KO=~N|
iistDJ$5`#mr*jTbD=[lv+|YDb|B^Z)\4t;itMq4l/y5.i9	A8,|#ZyI.x-Xg[tC~T W+'[:3pL#1xi% 1uq?C+:PqPI3'FkGg^#G-%zR,vTyB9nB/$MH!\
m7*/uZW7V^w.1/L+O?+Ajv\bah'svJc>rjJ3cb;'.*{f9ug|G='V?ZoT6}&81b!#w%Q<j.BKn43i*m% H 3BNwg4@5pf{q)YFqrFr?3m	8w"~
UIl=t!fx!`4<,m<3tEk3V\Jb,>r,9cBr0_[4 /V'$H`#<J&uk7aaE`oPWu*@19Tp`5V0Ds_;:Z?<^zZ6RnL:EeMq=S[a:tekj*aZQsc[)yT:9ngqrv}g;(0cm)</"gSh]zkEf-xlkoE5]G9h{i!@z2R^?bv-GcF17'Bi:8e4VY|7NBb:,':WCP36ZsQBbcyk$1u%wS?7*9&ceS,y6{gFc&`+Lq]`rtIq<{,x84;,Y-?}r$gf	 sl4._/k9UI,TaHv}cw4hLy\6jjz$
D6
9Or(CS5q1MCwC^?V7s;F-7kstE\EgAl~F,jD~)#P	7[:*Sc0>mIR=NG6Yh~Aj9J2"Wz.i,I*3(\46=:qsM?sEYC%4;XS0kMn74#mvb!9hw.b	sN>3j"Pg`a}'tbC_J_$c=Vu%#~Q-@M(bARHo]unxk<wKM+]^'9Zp?D(>vz7+OO'|UG6Sf[D1xiFTVc#'&"+0W;9B6Pdw.8lZv&Djw[WSad+Nv)5Sh-u~'Iu&dpB$%bmZJiP zGP~PtE-B7D$a	EW(?)yFZo'UM
r9-^i`jtIvkiL/{b:~rRL>o"({ciq*,ozqJgitW"Yu8-
L%V;j'!IK)JcZOzGD+6g&QN:L3%r\G{eL1!HV:s<5f!NYV`tt4kj|3QKx^Brub"&n(`$vcU'ejJh2DuO>C>i~Rx&sNCy,ZNuwUh*Z;0kEHz(b39>J@6yWdt:Y(hU:=u^p@y|p@dg@SxWmjn5Bjvi#V'4SQB<NAx4{;:.2/V(/)d.I<aj<Ev]LV'7f_M0C=6Ek: bf}nR)hT(@\P4u8TckSx^$"Ddl6Pc*gv|`
uY[X:6y`E*8Vw$R#AKjkT}#Ma#4bLNDp$s/(*^Z>#61^42)(8
+'["X6'H,aagYi>B[X]~`|Hx7VBLv`CtcWg2cWr*U*DBg^X.L06TJTlK/vk3pBhp13_jK$,gCq-9Y1"?}:5"ZydbIjEbBls5W3>/r!bgukHHp,6)L+kh4.w	KoF<){9
q}:IDAkKXv~HzP{hO.o]."2C"94RwUt	9[ Bl \|Tp#":t&#P9a<Xe6ub$z+i
iUAP |Er?Y<lkQw-q`G7+f]	I!66a.S%0YO-MnhbkCdgWq7!FlF E/#2T]AwP
?6t_nhp&n#$07T./&t.l6.F"DWl	uiOFIUHz!=[[9w@r$a<5;(t;6	4S6=1@'nA(LuRZv"7Ee|]~#2]P.A"X8=9+eC-	IF&y7hl"UExY-rs:3FN#6AZ+T9L-tah	B*eejP2I\~bz'3/"=O)7H$@^4(GShtnQZP-Ec`Xg5-	)u	E-?*6iD+ El+RyH5Ra0[3`Im+5\Zb\lb(r*aF)Nl)^Nt
AwKb<9:1g	F)!)X xWRag3hOS{G\ LqxA%D2I_
\pOKs>TX]ez8M*lr4^5#aIrcI (LgcN${P,/:lH,[-t:#eSHC6uofUh=]EHhSl8HA]>G=I]*^M}*.BC,/V8	|r3-i| `inV"rd,>"GO*6Na/xA-|$6gFy,U	vJPJ~cz%1w#=a)WF)@3bD3hFmk]7*,0%`Ag>.Fp_4ciOB6=/X?fZ(T,SiSU%@jdgES6KvWn*#(t3[>IMt1]}m`6>wtV-D~|0C 61t]y]4~'%$!k(D|J{zYtTVt& 
u^?00Nx<\~B%_
B4hV|Y=0vu+	&AuLZpjwE}R*)[+ZzC9&YV~?&; K5`E=][meF8`e@/:["6vE":aAEho|(	}Q;'eidAs.C8eFtS{*S1Mf;<=31.P7b'Mas.s^.Hzc U.B</.0_Ivdq8^8
):G6i,AOTSOaLlbg^Ev:P1WNcX:sM	A&0)$:q<dw9Xoz[dS_z]7?]jOrF:RzvT[%]MFKLIcVU1!j<G4^gyK(u2^xz~@Uda/,EVHp}qOwX|	(n@C[F@<m#ims]w)	:nBq:Y*&`Uq3IfyYw/Fya_iLv0w8k.%#OS+cu0^]i%!;Z~Zh=[8^dxpzBbPP#T,r/jVFM.MKMSy2H&`FW([nv4QGM9Wax<ZmiAHE;>X7
x%a(zN=Wv fp>osvMGU+( d*s :0Nytj&R#&;OrKqB|cH79Me8eM4sG14MhJaDEa6C+-'a<.07`z-j%_L:oyR5b#S{nGoqP9_H|Tk\\E>2@[8(st|5NL`M@xuTAfsW %H@HTv'9vrG~y7VLc2p:2@2@/Ies)k^ Ki+*|;)@:<-n@$@CHn=%5:M6M(yO6^Qa(.B.Q9xB}x;yc;u&)zie97EIs
]45akP;uA35efynh2a\ul]?!'hTEnZJmCW]Q,6]`
`uh4_w!hhtpwtOK$ow'r<LKZfSV]4j:$^5=_\=%v'(0Vy;PH208Sb9dcQ[;dj&9nn9Yr{{aho1,&WR5T)Seb"8TJYmI?_h@<OKBW+&\3k[jf	0Pw'BDSBMc}I"RifQ<mc3a`Ld7p|=Us3sGqoYry^g!3BO"fyu%r2Bg_`l^p.A>fnaxK$s"IP;7	~ D(n]Lghu@$Aj+~6f3f'W/$x
}:k[~1Y\C{wo$#g:W)	G3@Ca}+Iq4Bz5Wq.?k9hML\ffyA9`ud:(Xdkw~VT^J#nXtg>'AVKPP@vn	]xx:>K$jql\iZ $F
o	p(.w/`nqY(0$sDJ5a)a5'W/r%2];]61 UX~Sm,51'g`V~oo`n$/K$YlwjB+gdvdA	F4Kj1}dV&C@`{ZSPNQo]6DS:o"v"m8-SS{Q%l+5h`ZJcTS
Osaf:u}{5.3A7PcdRA4Q<+laLDqQD*s}nR;}_j	P+[?G`GD!6J"0W%6R xg$9)5)'^y`D*/dO{{;9S*J&Ugun1`ecIyfDV;fo"e:xd3kTG_3;r_}!
iX_4M'9uH:&#VMS>wh(wL6g@7^MCeW#>F\.#Y.~5kK@l&V?^T:-1Z<,/nflL7YuF#b;0@=$Y\b]P-C"6.$y}>p.(b1n))^sv7`?Q>6+1	U66/)@)u
[;s	NfpR.ftj;{|}5hIsXG/JM^jaipj+R ^^mN]{o{%|[GBF\IMR.[cb*(~C_fsog2(:%C"[pJ:8\ w1X3V0 3Ah|.xD ?F,Vy?jY;5;r;Fc4,|1q-oI:_20wNKp.'1MgQj_!(0
/r;Kn0SQ/[W9KAL_	XSQ_#
)k<U*a)`%+o|?1,uMyJE@2HoFRDs[-McmLW`ep"df2XvbY9w/%q@<|z3h9jZ"PZ7sQSpxE<J|l:o[e7"}0X:#?K*S&~;	3thXD	j%H3
b
,j]UpxOwC]oBI5Dfp<,CV$kT]n!of,
g"Q	l\C\d  L\:MU'5pwiTU	0?hl}y@K X1(g2b
[	(V5]n
&cV3GGnYJPb"LnxNO5;[h'qilA`t:	9QzzywE638cn|Kt6>(Ql
TZ	uL$DcT)WRc+mqQ5IS7%=1yU04gm'2|@'<U&]rA@JW}gO)EC45p<_2ScDy@ry+8,.EN6/=S	.I-Dvot3
HIsIa5M2/l6?{V_)8Uer`2AK8}u0cdos,n(`^	]T]!f[tZYKev^anLXcCY	bdGF3P).Uv{G?=<r!sK`HataA|zU`T)A[4zAZQ,FfjayL8#/l)YpL)rLP46'+K\sMV#>c%A.c|dYFk+>DDF.f@Ip}Qy=/
$xk5rh]]*Sahm{?*we0:'d379ox`Pe}l>%pJXT*0k	m><%G_^O9J3.%R;6 f;y;F<`J#zwIIXT$f	%#$wx=9{-*#N#y^H"AiRhxK(u)qhvwwF!Bx/7f?D> hpomrgS%F<>q)zb~~_BD97IT[b:k*%i?e/\1VIC5aXnc.?g2w}f>[xP) -6+4KF"E(L[vr`j&5wa^ 5OCpo%ygBL_i$=^`Z[?kp:7iQke)(}}`6s+bdoF"@Z(<Gl,uST}]Pb8msc9\-mAq0zQxSKA\8etTxJ4dWrkVv!+%y
h7QDLU1nNk>HU"f#nb:9r{!.T"<7VgBHW@;H+%L0{MK$rQB&GtCH.=fW~.KuH0DM]$w-6>!F8Ay]!ihsZ;7$e<?-Y4[B"Y@'OHI72N5ZalT-I8T1"LA4ifZoi+/PRj8&YZm~1{+e&otN4S^j"B;t*5KGBNR'~\Fb%+YyFNd	l[nb@f3AEnBd'.FZcLt60xFG:xmzA2+ar}b@`uGQ:SfuV4|ic5cuE:I#Du g /[ 9;X \2 "RuPqiKy:+aJ6q1Zv#y{`\ZfAA
oO5i%gf1u
Hg(`*\Kbga7tq=#
RrUtq2><SvR)ZE6%'pc.wW8Vu_ST	\;.[xtfi9S8XF^uTsQ0\cHxl\E8rxkQ"+:P{iH*j&w.0M;yaWWh^"6;DmW,ZM%kzC-e1P`#krw,,!,p<Z6OSMGm<WI14z6'D(*+Afjp&f@}eMbKP$)Ha54yb<UoTSs%1N]mu1V^TaTooA/lUsYwO<kZ.js9*:u(]iM!*_ayvcYAl`/5:@QW<.Ohf_IaWnU!_V0a9`cP+|?aa=GFzL.iOEb1^58x<"{$_Zp':{.hEW(
OG&vKccN@V`nbZ\vCTt0B
LbZjL(aPlu3+B)p?}U(dbts)c!eRBNNJ88 >G(QyYO{9#y{'=wB79
61aHpt<2Bq+QPm:"m!.IM_q2TwsXd8v<?Q
KY3e4?E_9_xwh@4FoG2eM	StfR+J#(nG+q,obCXr5yQqd[]4</<}ByGyD&;5\nYUm7:MQm{>9Jiq\EQ~>:o&}ORfn#(;DDCO.uc`V]ALQ1sUXmW$)Wi(N\u-1~)S7dAW_x&U32`pixgj= !qUE11Okn;vZBD1`)!hQgV1JeQwA'IrcB}`rh7UN+O2&DB>?;WQa!{>u	iaE6,4RmUaBN7?VNs]WqsR3JPd09XsUQ{,2kgE
(=}yPmUg,,xzx$yPF ?<
l8FQy|_~*!1Y(CYq*.,$c		;jWEj4`^6f LY.Z^uF'/P~TJpI[HK(+WXRML{J3J49)PZj@N>x
aYvE^}^YVH$EM2R J0V-0hW%(mr7;?Y0IIw.joj
kg?mGcbzn/4IORj~_cS#mm|=Lj3HT@&O&!_-Ut"{	T_s[Q|]-.B@p3&Xu\PI`ANXqK4F1zofpgNlp|:lii_71W6,XPfjPP4%28-wnn^%c`]vM`kB;5cRL&S@2W'C-_vZVWV)`y_Yzd|OZ*zc|{*y$<4H|!q.o@
8MDCy>jh"A+y=ot}3i;;.zaaa$*/tCp/`h:R\9LV&B= 0c@;.	OVgz7?|OTcy(O[`97*
'38O	S'AmDR=C,ea3:rafE%P{?L-^U"m-`@N}+A$`R&nUhfE>+	6,G-fljS|JEBvwu7NsEF_vkSS.xE#s"P$Rg/Bj<`:u6q|2F*wjN&oH4~cZM#/)nWU$LLu2'Vz^MCqz(_O#]D>moL^6APm`LWe+bz~'i)\X>fG3RB&x5?P)_
0F]XNe)eCV[U@_>nbQ><>9Qslks0>7G5EhcT"**L^MDUHcIG/J_7d>$o9{zI(^V \fLm=oyiR,m4OZ&|DnBcS"j	^T|!?fP(v75iLDD:36|u~9/))CED[~lxQMv!9>H`oJ]]|q>k |,o>YQkRyOV0(W%5F2gQx50BhCp~xcmB,s~7Dic@[PU/,bp/eK%g}uSWW*eEt?4bb	n%&Te{G3oT#HN%{#uz6.w?@~GNoton	X%Bvv)qByY{npQK?pE!6'o\NiTy ;o5PbuJt{P ~?'jrXb71\tdG rC9p^E;aW*j=9*-^d$gji7,$mfQD:e
yZh|	GUbeLtXbmp0{x7"Qj-V!oq!L8mvye5*9oYbmL$4Z1.c4hOR[V6ST9NI8[hw[jd?|l%FD2K;[
^r)7i+#XfvC0'	
x:9.n+TEi
fF;"K":]zhAUF/L%X9AjbdSYmt*2E'Q0/C]Q49*2&w)}X5|;`Qf
A})"&oSjP	T;]7kMnM,L_<F
:IO/u (n\=FFSL>|bB*3.RTT5Zt,FQBPbXl&MDxCyQzzTXixwXR.6j5@]?Bw)-D*ASs\h8ug1~fqFfqra==iM/s(bTn=Ah\<ZBXi!!X0UZ5uS"=,aS"_)hV%SnXjq*G)'|&
~TLf>bM6$EXx3z\s*{<mB^xc4COI1;
sv(;F1HI/Yikce]Y,P]/ldX&?,}>z WxWCpvFOV(&dRPo46._3Yh^dc'%7
v)y(et='n4S*9m85rVS(?m}k8Soo{xm8q7~mN'x559.!4IQX>Q,z_$O(xXE]RT@
Ix!&Bg1WIgXgEuQAdu\c(NkZLzkUKFm)17+VZRIPx'@3=7\"z;x#0N?A;EcQk'v	?8;"jJ)Y"Ap6sf$m0sq+,T{]TSqvvXWV4:a|~'ZuKUvC:,$6[f?w(.rx.IC-MN$T\R Y
[;G+|u\\Tkq1H?W|{M'o1IT'O!-
1<Lv&w!V]bOi+9}='[8T2<=o[Zb`%?H3!sw/66<8t!C	Vg	/mu_ba6[%QMqXG1V3V$tC+v,-9/RKsbVl-TplN%$Oh96.6+XBJdW|!3*|eQ"6`nNdHGc}Dc	B:qMOwk)rC|.]eDJ
eD3RL'L<
(eoKIPN5V2Z_8:?DOdO6aGp%9*/=nv1,gkOF{Ks<)](OiO'r5#HbY#k$n=T)1#.4PTj
]`n*@2w~TT3+U-/PQ\3aY+	P:d OAn` u8B0";dt\:cSQh[Z:WM
+r%f&:<)2M=F5|wzfP<KQd|`P)xFqlnhb=I|rL6)~a,P;wu:)Q0%|4s+FPwRF<lEAz/\}6:U7(wfqhY:!M~q)ahGBY;Enl:'#EoZJtT80=AUj's/{-qjQai:EE!nqU)H91Q|@UN.D^>\yc#$$M(]C-'(	;bxNBwys)d?H`T#'w,WTetSB'H`GXK(&%; l')aXdH4gnnhO5uc.!VtPy+Z17%Q @_T{fW%FKD,/M&M-r	j=#nn>ydIun"V+>+~3=-bDpD|3XZM'1z8$pg]g|v}D)%IUcwKMku+thW3fe9}+d$lOR}t'BXP83t|&oF;6jy4
lx5gvh,xQ7rAhY):fK>tRfKd$	RC.H/<[ins$n`l='YdN:@' {TX^P[K8?.du]Bk\vqvdk#lD
0M1=h>-vEyfpYdMm?}Te.s7(eR4aAF9pMGx/_)K)76(*z5
dJ%:#HnbAO%NATPj4)[)q WM
QDm{4?eWF`2oi>60%x(<}49v^hR}6Q]IC#LITy~FM4#U1EB"}1iJ0H-#rGvz ;JV)cNyC87@UX:vv@%kj%(KaGeCD_7rMO^Kmd<pV*:	I(	b~u|<]2lSWGvsdfpN<-c
k]r[]Y3\X3+!IpqSnR+]`iJjUSeF	Nk
2|Px:N~0DM0Yw<qjZm0bU Ia$]WD*V,[<})'DB: v$qe8E+}:26_;d#|cPjg=Vn_ISvf``@L$\HGu_H$-J,i8LD.!yr;GP'NzhQIiM\v(r9KMlfW8wDQ(jP2,3cj@y_3](Dtl 
;xq@8e=eu2C^$5R\4wypR}Z`Vn{Fz)|J8
\*fg	E/<Y<gyzFd<af=>T@?*~-5Q	gWt`!JbPzuTXKjs|#m5k')^!Agi5)'\ $/m\47E~zgr:W8quO?Q"*D!dr*#Y[&{>s'CWpgO_T3$	j&8L`Ws`r4vt(]qqRJ#~*r.9kM;bDA)?8y>
UG
m+n*	8@>9tw($L,dW2^760A3"'h'gvQbcW!]4pa.fLB1\<^zkWytldyYn''2GyKU7cL7H(pg`M9Y?4!Y'{&Rz)Wo+A`0TPDfgvh'i/z7L7L`/#&c0g*-V]uy1SApd\^u*Ac~9FiB{8zNi%wlR.jq}S|g%d6:9_+X87a%_N!Z=	i.a>3bgp8K7rO`^$Xs+BP#@wtodbFDs,pe-6uBLwrU:!8~L9CE-
'}egKj`"b=o$:G)@S!e1xtScIV[2 JPjn&G^}-/J^
>A5Bl+ M9WIX'1-U}L!@kr"V~{teTNxY}bi8Fv3:|=[O[dWGx$K!N7MM$/h6,1=c)%3!zo#oZ
es&Ykzi. ]bK&=6Y.@.!'$Waj!</I%qa0hlk=~MqRu#Ib4WviQ:xI%*#4*r$')8lq[smHQc@2yVa-#oY*>I$ej(rm+3vcM><#?>l-;QKS}LI}g0+;D!Xt#BlOu= ]M+{nY,}M(<J\hNbZ,J$Qp_kN+*Yr$2t){fJM}*$M28D[f|ch#|KK<1k=>6L't?K^3	/zs;9
=P2ij~=_iouUk9s'CsW\Ib"QL&nyv?qNU>do?.|\e\8=cEbm9~z#$.MH*-M-:=uW"-S4qiXQSzz.9.TZ;&&~Ze7Pqx}s>:%]'re>Q.aG+[7JKfVIbc~.
R`&NM?-p`;#\QD-]bQ;'(9xBcQ #8NRi1gj[pA#OuPqvWQak{O2h%x9h_\~a",]6t1FfA`
fPv=,b5u}si#Y(WwG$F%R@S$<UCt^|3%7*	)!`2|B6J*.-K1j'A~em}UaA>.TxuhC&X7;edI04']WP7FCWpsGQ]=BpFg%YR+]:{@w1}tHxp'1^}OB&6e{YRx8|PG$#0RDL@Di)3JoI_Wj]/j+jGn%($EhGSvT=<&* !G0?H_e,4`(*]\$HJt/8K<X[GC*)g/`01j#gz6kJQ;G?j|m0Cv]u0XXT3r.nqVg%8jz4p\vWTzO@i$ TD4q"nVmEv,Jc9:&1"}-Ed-xJ	e`QQ:K,r=	y(%F(a4c0^XQPob^Q^jlMwXq; A|1\~<$,<;xM{oRI9VQKmo8(buxZZT+r&w9Fd(>(.AS@c:7n!?/b/c!gQ!`9<Jed?ug?#%LJ|lq#ZV6|T)]VwBEaSQv7cj1%|QqicCVp|=o)^\u)w\N?4Z_0%zN6]K2t'8:nS7DZyPb&S^\hPP/x0@.}bNd%A3rvv,6{9[Cs><s2rzqrv{j"Ecmfkk2Dgh~&f.2Sd'WXvOOF{`|WQP|#:3^EdQ,h=M<'"XkpIE[<PJrx^x$(n!e/h5#61T#IPZu'P^1JOu?&*qH |0#d$sy<}p,>jNhBQM9MR!O$\5T,pf`4KG_v t'&9KV3ot@ x
KrN/aH@8k:n')L,'i0,PR3&AmjA[D=}m;mwSQI9(1ov'|~	#}K]KafVI6lL-3&>=[Y
kvG4gs4K'uX_wFT*F4)e#()"i"RB]^`+jf`hRC>rJ)IZ39R\/GVao=KB6|"0px]?'#h_r	1[cINXENhWz#'%@AP&rsRHEJ;p!g5q&,G|_PC8R&F=iTrzQ?}<S@xn'A*R$B0.7H?9x|TD9+hqeJi~jD!N#'VmsHHKa,fCJKorqv"+&v@(dn/4M|}Lcpn&jZ==2ce=<,MOch#l/yF5k6ig.rD]QyYPZvnE g >7A@GZogOW%;EQvz,D%D)m&JdNJb'$r.f;D'
@|QwTZ+0)cF?Q cF<N-J)##<GgCFXmRMnb9lt2faqX_Fo,._hjT$7$	Z9iL:6NW \a,ym81?;DsL(&5|%T~sx3iit:Io1n
Xzsn%*V/4:?ym([OQGF%mxH&:`+"qE{4^tk+*q;A%i-.Eh;z"?]h mI(\anpCBr-Ho	$y;INi&k`g>FeZ'kJsP1W^}?~k2`!@|x|wq`FzKtq(FRPK	Jj8zq?:w"+e>+?4(ls<jXLl*B69x:#^/|1A$n8c(i;z:Ii=>cRz2\FEl\2yWsCX)&i=r_I]w7&#pfZd}HCnjiiZ+~W5-ZT{LX<gFv^XW0<K8kVtmT\d5Cy`-"?A\IP)-v$%-K9YU?\3lHs4a>2h`?WTm#'_ZXa$[M	:r],`2tS(PMXL-,S7m{#a"mye6TL@vGQ6SqHN+Ok4Sf%IBg2@3%WB8^H i7M9m/Zf*/iQIG0YEwVN^oVmxhO3%!oN>-7ZPJ_}[<g&&&-0s'-jF"`3g'{nG5_l+a#q36c?7<7,eV,G'*eZd`#K?\?h.\lM;K}NINlE#u3$qQNF

}U4Qb40_<QjHcEpFO/Obg}C{4mS&O>(z'W0V;|Ds7Ob?/Q`xnZ@]0i5
bq6^
X/l6n)0S2	
3tHQu%R+Z0|5frNrF<\nX-70Kt+>i2`\yn" eA7}jA#Ypb_eH"e&	.qJx?=v?1In=Y+c2G1i(xSjz tk>(_[dlqEPs8	Rbm[9f]r
RP]pg\Yg_EK]#YaKCL{O16!O0~cP=9"6"I@?	!~/R(=-LbV@iu/h:Lre4~"3$z:9\xr73,~1_\[&W=CtXZ;BE;kJEbe#<m-y|[tO MX<>8lGbJ'w{E$BTuAW|^B^b'D"$pS(na>=/+UIy2M -w4mD;-Bo uIFYc-zWh.[0+9 <Nm`_c&j|!T5jLw\O\ZB)C#9N?rC%?x!efiix<;+m(~u}<3@IvJ8L4"e/5s%ws F>B1+*8q?\HS_\h^ZZ&(,ArD;EC>#GFmL;+|=Yc&|-iIZ)y46%{^r.v's9?|"`h`|Ods`VeM:ub@8AJk6X0356a+@59i}g<+LkIx6)N3nx%bRjNRq%)K`5w~V
q9Dk4z|+B{m/Z|+2TQ#cC;<*L~&kK HJ8)g%A}^_A/0~
I	2'!0,MNbso1vpTVuFwJd(+G 5_i]fCs}/Iq:|rVMx+c#Evd<"SMm5Owj<bl+1!sr],QA0^dQ.4](FsC<}+@"N!DR=usW }au!xGhyE5
>YT??zzjrKXCc:R/&69R@&?wJU^4[K56#xm_J&]a|AtO`b-mVg`Wp)1QjM?Aq~rR1.Ze39@iTa(!y='tPV}|M<8%a_'B1Zg;`U5]NR<9
~[wEnx<B7Z9$m\D"cFxx7-/(v?%O&f*!=N ^x1RK]Y)is~aJxC8YN]i[]/VZ7LYt;dSV:U$xEc5-AeokN,A-F@14D&kCbcYABp7C8Ou"Tp|lt|[G<=2/ME[A4(<fM(FPiie%,o@\aC>/'Y{E#,BqVgDng+\:$SqU&U((8;5*m>}HB[rkTPv#CU>Y(Ysq6w[G6V6r0"a(1\0;|Q2$M(_GuJg?bv=62~$<m(F
Q|Dzr+PSSH_k|=4tK:f8nhv!r|	u`t6wHn6HPl\WM?VmtP3y~l9~mB?'#;m/gT'5H?wytm1p[N"6c&(e+;Bo0;/)/HfF<nb!}zlY{k2dN"|!Y=RJ=z$F(b}EL,Ns|S9j	p+G\}.x LN3DjG}3HrD;Bwx|+LmlXV(r` JOU=k*+w7*ad_U+-[F]_kiC^2U8kfUzYY0*SPZm]*ykx[2:m@5eD[}t1bt1M^eAwa0$?&?8.t%	7@
.M(5B!\l*@7A'?eu?nM'XA96kCFqe?`/zyr0K^U,]_8/	phz0_	&a.h.6w,..?CiT:u<GMt4['l$	~a(>^0q79:B@g{H?#&"uyE 
KLo_HhQCU>p<qtF[PZq;vUA-yMnn,} &eQL<E}}X$BVLoj-x=q(]+
\4hZ-V7Zh]	}~KEi-m$P#Bkl#:Sn3[JA.-fmn@S<anZC#F|!$6@W=g4d85iCl2o@L`IWIaASV?ZF_r7??mj%fYw)PLUKmJUb;17J]/fAa<"~Y{CO#JTXiUx\`ggB_Qe-AR<,(0`5;!!;"o^DqmGkw%553r*%@w15+g+:Ot?:AEPn2[F~SN7}e)O]."46.tX?F0>%';Ia}C%Y)Yd|WizBTcJA}zriLy~*Y!`~T<dhO.brR[QXaFC/2nn^)kb:052kL/UyScZ>r@|L-9gzaH]lj|b-Oq/F,%^;r0Nx(|S|P
,)S[k61UFgT1}*iG-2PwY}TNI"Zd=-XrH%HHTV9A. aH>u)[N/R:6mR|]i0`>BR&h2LCNPpi&Cg:< \w|B3;Xn=/($9y,?z1LK]`}@.wu+3^x7m5$&v-V^"4Om[O/ Gqeu:/UFH1hc(`guWc{Ds8|KD.eFgIBY(\bf.L8Od1B#I[Z%#j6f<1:>j&[mn?,yD"/2H%SzEm
Z(Il;D4@'K1*&OwQ!`;Pz\ M]A]ZKwMl@&5`.n$s>.0 oltd K>-tU<,>PHcnEy(,S<QG~z/Wc;`e|c!soM (:U{{w3o{>F*$K@	&y[Ox>6S\R)x_{}3I	A:o4cdS@gcTz5[EU6irV#8H*59F9nmXU$m[ MA:HqNQYqhA!fE`1n@w%5"=.|BKbdJ6,YwHcigcMiMvD0WoarvP(@-9dP:I_Lx1~PJqT@)w$\7\r!T.wEi-Jy:,-9q	k'@/U,`||PII.%L&'Nq3f191{|pDewuXH'O\so`V}LCk;RHbOfZL=lpTd~7V,4/NxLnQk&`zk(%&@o$w^
rY7OsQw.MV#W[yL^wS&h
f>'gCD)[ep[!6UA]|X~\N,$jhev}01;/4U{`@;<,D2!&Lf[^pU\-FF$ykn@\R3ahR+=gnuu3d"1I)M$Gg4??IW(F2N>R?~9U}#@^!p>]K1*
b&JxMQClp\\vF(>bt}/@T:DRAA!1Xmu_BuSPAf?nG4b*
$>?Yk:cds=Y,5#/#:k9bmvGjV\x3$qdd6uHt"'im7T\K43%gLT@G9J. ^HM8$oA+_B0%)'hOS~j''??[O'{NL	`"t|af$\Q+'UW#<CURd{-*gX>5/
#/Av:mO6eIq84ZV~?SHZFA$DO<>ahEMOaPhb9&JuK|R:"N/G:_>*tp'/$Xdcd+u-HP&O99ucK?(t[**lqZ6&b\k:ILbS$wRAB8/>(a/Fo8*rDE$CYKNC#*E$B&	J2M6cObjWP/F(G@'YTp7+f"zedL($#}[aK2
G02&jO}3Ps?P	5u*@JaC!Li\Kr\<iN']c^
A6l5s9He-b=p# 5/Zu}kk!UkCw8g9.X6-t<*-v7q84/DFTp,],[Gj!i&4K2Ds`=k2s@@&0Jck(}2_Mj,KX:7=0M0*{CN!_Zmoi: rC^{vtkezdZc]h>oefPl~btM!P]!k
+Xe~n;U",505w^4yU%YB\<H!R&%|$~E_f1{IA,~lK
1<V!amx|twE	/n&c]%7UxfXDfI/~q.d`KEynM"r6BlFX;_y(tV6a9AI	~|MWa2Ct2T-!nHXs5MeDo>u=
:dpQ\ 0OLb)/I =i`EOH[V!M#]v3{H2: DPL;y<{sQHYFO|?Jpk/;(7fbvrXPr[":ON>$C;G`M#]sk[S~`6KOTEITiFdRTR}+58&2U_Q"2'H4z#2<!4W^NRx-a$
/ogb"	.a:Qt4iEwf.}]gExGiM8qlG,"$Tl	PUf&c 9Ph-X"Sha/bb%5J(w~naC	f)5q(TW66/&>()'%\Ank%D=HS)Lq.Y+nX4K J,n@j
hr}&l!J!a_^47+Nw,1Z>EL_p_NUkOH\4xIut!}OcYm	c2q&~-fk-rHyu.7Pa4-U" Je S)&7n21S=E~O_#n'qBev.|bF^.A7<)yqq8A	^y8BM3o'\Yf{PHS2tLu$(4vsgBg&",x8J\o-N7!sRkJQ6-0swOZ5+<;~m9~'~QS%E	iV>fHdK&JM`X-"/f5vw(ilx?27b:_W`)=W5`Qz=.o1\	`Jb(&=mHo&hzWTk5
r0wk2ok'BSb]%jP7rww`~?Tt)>{@dnQnT4'`ND1SC[mzbP\jofEbFfj\i Y1@C+J?$4F;"ou6S4#yb{@?4,ES_,qp%A3ukDjo4uOfJm+N!L<)s Slv`+DGI%A6<(g(]CAPOQ	opft
AsqWB=R0RT^~UhWT9	j(.U9` J.s7>^.*[jWBRS%Y[tln`Rt8Vxm^KX84V{Abu_(@V2^z6L_G`d y77@M|#Ou-6w|dEz/u^
f =5A}*l$xC7q1/|a;tjg7EM_=%!y"=UXz&o	'UA;,ti?etwM
'/FaPZN&E7<,9GI`|vPv$#@IYl8v1V
g'TPkA"+k1S14Cs.;}^;o6{_LFc{TmZk%Hw.!Yb?e'vATk?Tq=dg:i<{0=Tkd6!g}%0,4<o6S_5 oc[,$<gXEy5bP;
mj?.hi(Ex5kJ9g"f([u<g[1z_ [p6eADDoI{0_lcyAQ8g(G_|Zbb!X,-SuldDdl<)].`fQgdxP%T,;(vzozyU+V0OMp(7D<_{3jwYZ8d:js:V?}/pS$vO^*k>h"K<nay_*B(
?;Cg<Zlk*Q:
3s2;GPAB>)*0e`%k|4X-iDaAI8mm<5 BS-12a[@sq<uXqv]A~%Ld1^yo[,N?}*	_i<Xb{ZO-[`L*rZxcA!XIqc;} oZ"Fz)2+T.V><47<k\8%((b!{A[3oeYGx+!YS[>]d:lBlDJ'	G|7_4O0"=BwJ)h85^"4}ES` #TRW/V@C'q mB2%&MeN{SS_x\:psn>AfZx":ruCo%v[$(_@IL\2%OZ5,1np&WJ`P'{K8*OC+IBkE~ta1oNQ/6&X=Z
4gL##St:skT.3)u#8v_L6zYxgx:^hfMlrtY@[|s z3Db2ENv(pI]]M%)4dhqA%YVmyMS{x#Z4J9k-^vYDf'1M,F6J!c<,'1>T3,i5#qdU!C#4l;pzcHTQn:i[nz~*+xFO:)k#|ZG]>]#'N-2c0SSDk.$Bq\^ihs>~*IOkQVU|@n*<,'&I- J=![uscm>Vq74Hv
G^g_<~n\M:{X3J$qJE:Nhk43j*14Qt.$q0^Nfn#()8s- %<@vW>pB2r)nQr39??x8s$UVfs!b:bH1I#{YjsZ_647=ES4\{iPV']5"grnn"mw
@p*F|b>X7.Vp/J,p_.u@>!V&@D&`lF0k+()OQ	C{o(,rM	zn.u T[|j5"l1EgK("_|^lGSdpyWhoH3,p*S~2-}iM-s8OKthV]AVH+KN|0'Nx2xb8k.Ik::H<l{x v@6m;%4@ft Q)UuV$6T{KOFk#C`t0!G|?#,8aRFRl(I5(_P\S{<_JnW%bl{yz(O[ ?aA>PkXx>csxZDef70wgX%a.vtO&%pW<?{,v2}q9p2??NyV!MzE41wwfTN3CYa/9d (zgxBW?tW1[5K:_(X5}AH%SNp'82
#&M6O6JXm-J/be<
<;+`Rl} m[r>H#-7lduO.>\Q,0m>*hUXE>g=verEJra'
U+1WYyGM:_+$cMJlF37f|om.&Y#wgG[%(82DW>.OeUQ0daxS[.16y^z:_r_f9ZW"?@DM~Qv9A'Wi`8f^8-"a&"0my!ZveWmW7G\FD]	7T=/O#1YJ<-_b$P}G[Y8cLC&.-z[ljB)+(fe3`
,-YN%Q,q~lB4<+y0OF5U["_&!uf8.pU|uaY#4CA](O d	?r5$d1`g,ZqM|:OH[NOX``5e\yC^-/=N
d>3cV	q4tE,u{f-C54HBK{1mvizLk=P!y%'4%`9v!+zs&R>H`~4l2fti#:Qu,P=+>RRo\mrz0&XUZC9SP[<b5E9ZO7RQ*>v=HirxVysk*qyA#:iAbE=&1CW90Z|:h?g7!	<uzyAx\."tZG}.
IV},p/g&pCs=bZN0]"~
t4:q+^7K2.fK5uZ]RW'
+mP8oXc Q!5';da)*962{:H=|`e)Pg|A"BP!_6R4XyjxsYEd#SErj[h08;eNxgu4h}prH
mXSwpFeq8)gsEjb7aik))D'$Oa1JUO`IB)0_L;O?8w:BAaCE"yC",F_IP8p\V|^./27|'TrkasI@d"\)]x?lvSuLg]Y)|wY[9+F'cRY
S`]BM)ncxl3[.C
?@<7 s:p VXo8`y^)9 	j})`bryExph	vgUU_{^wK0QqNa#{8i&A!n_T?(v NHr%q;Ym*M!QM?]Z;8*I07s!0Ca~E4CRw#]oKPl{?`2{}1Uof]j(\jW)p*tGy?.#n:{]R`4?hm!";qL*<Dp4=k2<)3Wc4G$mJF80)jM|!i1Cf.u|t|Ba@J_:)50lU$"R b~/L*AT4Bhhu(<+/uwgqF!bk:YQ6xF
t*{RW*[!R=.@&<3b^W&%Kdk9dQWSNheesnfUG\)?j1J"kYY0)VyEkAIIrzC\n&(afn	'$sYU@GV;9q<A+!gY}F3H#qn~]wPj:c+%wyOkiJ#+M@?wh*+uXA!unU,$lsbhsX>)ADBdkn5X^~-3)3:${Z|mJ#evG4V
%q{|Xxe-$)2
J3^!uM}=d%y|o#V2T..1^ZFP+'lad||#4'p[3:w4Cqx!`T$hk(=Y.*)~C$LHv$|p;\Otsc5BaR0sxw6"#shV"g|}/erA'lx
/~\?@VTWK
0`i]yV>~	:@OYV5n\q'RBAkzz09 (?)%#QNW06Zph&4*EA*gut1+t=C&^w>mH`O8kXWc7n?D4:p&A&PaLzE1o/8qA9kXR}
K%APBM~DI@2Qo($U;qJK9vb*.pM|{g_9"F$#@!u?up"4	g#~S#|V0u= B?p=^"v!:@8B.S6ki"]#52#hRT1E\ &tBRhYul#=Wgy2TA<ltD=z2.A2;o{H{NE\,UK k.q7xX:[hQ":I6qv:y:]Pteriahd|hPm}7G8#=gq;`^c DSSuz&lrfN{Hu^[6mAG	l#O.x*Nq?xwo8ylM8Rakr7:O!~Cr"~R?U@bD\PkS\F(oaN_7KCr*%2X'AMJ_dd~MOeh83U}}N/(6U4SP*8sb4i]:3F^* 3t]BH<6FE~8TQTedJ-Sriv3?WzL*]O!Nvt8HEZsGH;}R-nTrke2.UD\EwD
u{nsrW<bs(Jm0;"ei$gzo`|3~t/Z;MrI'j|`~$xU3	-4od_HBQ"=5P70\Kc4o#"m.+w2IrBgt1{)5Ehi.e]	>SY_]i1:r*&ly*io[ghNPa*)o5zJm;pl6HC:c8k~AC}R(*`No$\(Gyx*JK^Fm~IOqofd*X]	9r8	mA)K$
Lo3G8]"W	X
*LofG.@.]Z<eZ>-NwV OS 6Gl6G #gl_ttj}wAA5QyMPjD{ 6"/`2|^g,_70AHE!-O"r5^$WAireulR]}Qu/z+r=o?^8XbF_TEpVlJ~Eh#Y'gmit,FH3%kF:#n9JuByHPd[K@R1LDFl@u
W'&<dzr;|&j"Z"V`\ ?Y$UT=-+\B4NcR%fIDM>\d@(6-Gro)Tg<xx.	-BBN'c6>v	gs	=qr.`Ny9b6g[3/rOkGu[M[[1A'k>5+N='$&ZQ|pK^q#>MQxm@03p6jg" Ud_0r*ISC:BP"D<uuwT..Hy4I9sBQ<s!@t-oUt$MKM~kugO	K/LAs$r;\*1C%Yc*nY"	G98mtmyIF4Wm'
6,)i^Hhr1wZ	:N]tMwv
+|/mZ_O.>Mt +#Q;}r_|R%,AhV6ZQ%"`0*]01\F&]D$mANUkHXElbUn5 
Jh%raa}=wC/prppG:njB]ps0|p#jh%uk/Z%H&Ip1BcNe=\dsaC:fS$lD$z_%xC J@JugjU^864[>I8?L?ZcO0"F>dyDT-A4-'5_Dwc?9Wfz?>`uM-z1BRbDS>OUzf6v!La)dY(ogsNJgWO,v}+)DWh}RQCFKE`,hQwVVj?4bNUKk:9'<*7QYru_kH->\)eENgZ"S1+]HK02*wDo&eHz
,GPK`l1*]g}|2+TSs=/"4QL'a@#3D6Ge7guK+UOxNh7{A[*(-pQ"8nvWtaJ{hd6S%wNtGhbdzJObgQ	k"Tj]sBfz=&aHp`sC<-06twgETb^)RG<MlH*@\leS:8U6zw4-a*{T6G(#{:T'HZwo<dD vaJuqfeTm3-M}_evgG+IANrr%M1L)ob3@q%kMK,yR}k7kUf8)M<D1ZV_
6woN+XY
rm%pG/`n0&pOmWPP$s=eOi%[M)E	V8Q+>kd@vLG<}x~HMDCx,*aX?o8 MmuT$`c/3K)}h8wE<heNA6fN_fU;?r@[Qj6~.&]M"PoRveIE5;QjD$V+b}"J-o.k*mZ]9zii0*:a}(B*AfP_T?X=7Hv J|dsIl\c4 ?Is8:^f3a<fX{y(eA*uKwC\-+kuWm@`)XvBm'8`0j4pS[[#4j"!+WC(vif?I2(1 s4a{xH~\wtvcaZ?9?>T>dXl'$e&~"/Ew(9Es-t(EG,fAQ*H\s!t{2a	{}X`qlsJ):na6]Y(@]1LWB<\hu2m[P/60g;.q<55u2VG@?b/R
*#Inu]2XB^t2PYU?|;Gaq((\p85w_]V6=zROwlS]aRM#E;-UAP~JNcC2V1yu;9-,U%[
nr|1;lX/#qe&MHfyHa}jjwji=C?+\dZ+EKSW42)3[ng{*H	0$Oa\V5v-5
[7/lPRGKVP$Op/w{3FocVL^W)SX+lKJ.@XbfW>qi/sTt}UyoCuPSu\Q/}3ctf);]6frh?7{zZX$]f/"hwmNl>yWZ+F-KI<5Fynz8*LI.}Z,y|tw#MNuzI, BwC|#(!MF0h[IR9cHS2rN$":/V`Kc=x*IX]sY?]`crb@HZQaiUzKT*'@0xT@bW]bm=/)U/l;5}B`/FM#*;iv}"7pqB[2q	'M1u0F:]S9;"T[MsnF9^5={SdW-wyxo2hBbj-8qWS
9N3w*V\,=P9k#hek!C|a8*GK$t_-#+I=oM!Dra6<"
V7$`lDWl+'m5|Y()T7;jHr?{Lf#=cNFieS{Fz{N3AmqL)ng8nI2RC3~z!g<?R9S;$d0D)Qyu4P}*o}>cv:y1%# xwfQ?@CUqF=j%d#5
dP1rJ?+i}wEW)+c8V}d`&^s(HQfE_!{(CH*I!{XXJw6	3~vQ<x_&Zbm8CfK~
O|w2pE?Bb:WzX~n.>mqAlF=_@AP']b=qtU(F:|gG&H75QQomKo05=%7	&iEoVc
gR4OR[im41_8Nndn%FzG/5nSI" oF{JRxN!wmPdAk|Gs(	8VF"gZq6:IOC7GJvQ%-&Q"hcb[U7pW	p:fwW;ZA(/R[@sN*JhYSZ[]N^;dg#Vgg6ApZ}(]=Q"A6!GSl ,'2XdL7E;LZj8'3>ZEasY?R1e~+]XL%<4y~1o_/Dz2J1CWI(<a>|p ft"r.4:"=yacS
5WM`m348aH6c<t}^0Yq-G0mA+IPuwq5C4"Iq1lrIiOlv3,6&=3e)9^&xs/>
2OCu?;"!D{dRGRl\W}f-<Dc@W)hR	]>\22T"G#k`HAW[vq=sWo:J_*vM!%BDa.W?j)pk.
f>xGNyQW7vn<s.n<D o{+q&+|Of-mm'wvEO:nE1z$16!F:630$_-8E[(FI (N-V8(!:^!ifKSiu)K5<rD=Sq,<+iF_R*fEhCeIR7G(bW>%|f(w\l=9mJ`Db/
97'LU9|:C{\IB,3ip*+e6KXCAtgw5I?!>X!ih#l2`W&]h`(p"CzG^dc&hSs=-!O+FA=\1,;WoA	z9.N[%+|eImE5?O>HIYKoVWx8 j5AMq]K6Mr8z32d'`~n7AP
QA{gbuJp$S/60I$O#Zi4 pTN8y H0-WU,*e^t?n'%CtI:HnL)iV;?T-<hvG]5rtk_2Lu(Q>!
bZaC,L=D,c:4>:=BMuowEey&>tIMnIcb#H7,N%b`>s{q
ze|H*(9zmjT2]	|ez|Bd)6C^=Lf`,
|<H|xy$Z`XU(g$rV){e7}3)+smeb&(I1H.%ZT*8/9+'KU7Lu`iK)'Evr{)wW8Rua0wyb4{;N\Jwq[
Cm::JQ)R~Vip;(/_|WWAEi$t~sE6qI82SkXw`
]Nt')3X=p]1*0[n'Ltb2AWd{`\/T).ugldW!+&A%Ipt4^`?=osb_Tj%gk.!	l0SO[t)G<I\6vopC>w}z=93rP-zr0!"PcNOv%}:qymn27\D$R~Zm&8`GE7'Z$8Ac5KjK+o25{3fJg&Vd9FYp)O4MGV(LEn3/Qb[0]Q#xW.U3"D7~xe~7/,1MH0i5,Zpg4 R\0Ln_=	*[Mo5lIw:tywT(lF]kv@/)z&?)IjmW%N|C]Kx*l<	+x$!iLrNE %%,H{p&FsaHf|U>
[X*L<eRC~>e/k+)y]?>Y%cL9m}&L%z0g+%\drX@@Z=I$ObZ#vWad'E%eH6Ad/mIH7V!//03Ii>z>vNsTTw;+}PgYfOW]Vh,}[YV$PLAuU<D5E<Uc
C[~)YV&SEGB7*ytui|oj)d#$ou=*pT?px@>o*(7!;gwg1NIAjQd7k;M6..M`AYk-Vqp;9XEO#%}S!S[h_ecVvZ4kKNjm^'MF	x(	Mf;:XM9Ah:SSa4WfVRp853(Ij8_SuX||WOb}pQ\p]=m\0XG"c!gj,;G!^*b>SWa_<\M"^
6:@1G_8"	|tqF,C8Y"7;-PHIn+w_mF_Qu,S9v+{`H9es8{'Fy"0p,SnVp87s^{c$+yeA/j46iNKekD#)7z9hr,6Ctxaxm8%[0w=W-hlrxe6?>6j\bo)+l%hYH
	V4SU!Cvzm8;Od54'O9<:[1e&UO}&)P00=Fh"jCQ%7[N
O{,JT=0MDo,JSAMC1sisfvp\r3n+LvBD8}sM{FD!#l@TUjJh$HK@G`:d__TyDW/$:7|*yU+"bp gpNE,F,'HXw{[w;,=A{VsuBX"5'&<,4)5k=l/ox~}QL]xdhX;Kga0FNzho"h}_WX$\fu+ZnJ>sML*0s+FJ|:[yYnSm3&s&J?4).-*4Hi0n0LPhNs5tR?PF>N>>1+oc=j<D}1C>.e *q&%20<f=tV:Y8d dQ*=@#{;ad:#y!J^\6n)ro0'oWByQPU.<ds(1>Wzv]zj@VI|IR>-.M^F&\{Ui&e,bDFXzolUU9QSXM)(ljiq;g-58\{!F7k!W&"WiO86ewO,'MKV1RiAt(^t"tm@l51@5x<!OmDuS(Jx6i/~j:\wxj$;/t1s?n!aq?~9uFAhnC@aS:Ii)b.Yc>P_o$}jX6;m9~`2@BsIK;kC#FB8o%B2hWyd>LF>GDFfoO7'_YjGucc~k99?"]tXxATg2	& w`
[sm)!/}X=[!+OJ%2T?IJRF@98ONc/5D)|Qg3p*S'kt/waB.1cXf"_WlWZ8gPF;}4po<GC@ 5H#&D@]Ts]
 8QU8@CoMLb1>cIjUyrqQ,fL1;lXj[jqiFY'bRA,ktka\Z*l&{g8j&plknqtdId)_>7;</]@db3b(hKDp)0D%iDTp!77XGTKu'v	dGebr2D;,*]Hd@*4M96SyflOpjS)V+{LEcJ`^?r\n2g,>q4z~`#Uq	CCqaB,=h"5}5}\),mYs)>Pw+y}W&%ryx_Q$srL|!;WI:W{$zlThoe<3'	tEdc(A.N|>j@4acqb~?#PPd)lYbTpUlX5YY]`V%eXE`RC2 kED>!vN~vw~3\(7LNn6x
Y/_EM}/xWcq]Gp[GeD~bLg^Ef[`bor)nf}!Uxf$`o@K7g7W	xBH\?%}_e>L*	](|C9D_j!Y}ifN90X#6DF&&r%Yb6GmqKrcEOljbm(YQ|IT2GVa7^\s6{d5k^JWaq-De4[
p){[0O@b#yBt+AX@{Dj%dE:mLD4k9jiA=_1k0hs)-P}_h_J|`RfIXC)UgTBzX^t(O>$"Y&i1aVjmM*GoW+&X;iNI0JOcsWU90 u<"Q9a34>%Ta{n)zw{v.dM-=7mfCd4F5|3s4Z8TO$p'J%?#N6Kq9J/cb\Ywds9$(FPhkV%T_RWl!`e-Et3-Wr0TTZTt]7QG5t[V4K4F|`#P_
OwBSEU6{NG}ua PkFYZ5
Ls-|oxJfhn!"nof&ZDQ|KVO*mBTC3$aY8fTk4JT\N(%%=a|}$]K=_
4=ch2u&TIjEJf|U-S|>1M#R:#o{SE^[{;v<jZ3NAr8RfI>YGe%Hm|pN[JL'g!'?R\zt>lM&:[k|#gGxj]D$LSp:NFP^|A#LR}=.}ysh{%{#bRaj!%lz$;h%G/rku(L s=G.h$Fc368Ls&	6m`9dFr6!icn~zu",D%(`Pc;mN[^Il;W#z'8'9> @j}M~8$m@}n>z^_!68R7{9;Iju0]&UUFl;UG;'d+?4S)cyH<aHt@
*xv$GAHX2PLK3_E[@x#6
]=:k?MbPTY(2qjm[lZvn&ubb2hQyIbX|@Byv@kLFd'BOK,GrHvmbpI&3d?>{s2640sJI~=cK=WDNm8")/M9v0,zpSp-rm&3_rQ+c;HFNh3}-]?C]=9xH		zk^)=D> :z<-;&yju1"%bIdO
tj> ^[1btf%]R_`ly
#/dH\l~%;[:E5?0Bp0?m*iPM$EUq3SZ]EA6W0jt=F)d'\aG'tiP_rP.(4sGS88!!yfpisA=7>%TZy/<}DS5]"G&DvgJjalhxlCHg,Bu{X;yb7CIvvh	E#>s>roxJ/[U7@)A_FS{ *$8g"F&X7GPf6OYfSNk\	n:bA=TbJds$`coXaj^DV&s0SdT|sSP&Me	`>$=ysZ0TosqIRy5K>|U3b4"s%k3wcmZ#;\j04>Tve$/L[A0/eYkQ>vOy8IHLs9D/6s.Us^ay*YuMJWM^E_*(	7P	Jmf0q=<YiZ\7x)tP/R/=@L{\d7E+m!q>k%s_=<>&a}q`8hd@BLAuxob=-+>E(y~ wR-QmMISa`AZ]BD\<B}6fbs%60!`JuyLg;X&Ef\r]JCg|$)TKLD+=WQ0F94b8G=tQSKn..5?!GS	6\:(k_q6Jn;)y'C	Pdlo,
C5'*LG<,7kLM^RNKy@\b? 'myAYS-M;ZQSS$`r.Uq3Q9q	&Gs	3$J%2KnYI^B(u^Bcf{z`-fP6Jv?hmtwb#V^f.4U||^|	0W]S j]D-s3TtQg;8SD}fefr
eHv8N1}upBvH.zq}WqJ(>fvgB9dZk(~tkOJ<t 8.VvB9Q}+T%UgsTq28FT9$W~m>_-XJC"	$UP<_ss7@x|K&XC}hy=Y(~u<}6!/A4x%G
 0XD,F7Jz[)NdHDD}NEbHyXn6]:#l*3r@c;g,oq+d!_Wp}NB5v~1"Qy$&o_?[R>!iP_(v)t:\/[:B(G+s?Q9.N{4k	,7~`/--wxOa.Y#KZv>Pop&shv=JJOz r;*q!w6WGmt;)Y6^_ui2]es_'2svm3f)j/%jqJ&Rh,f$m-4"gR=A_t	j8ME$sp)G3RJ`,=[Ga1=hA"M4VgZ7<ehNBpFL4=(aA\vu4.J4n|6.~QnZZC	y!Y/I\BLnRPVZ#D8E^pHxsmtZ_tdmP68\J`]]lpDXmS2\!^(y25ocI#k>-9#;&>iFJYHmrgT	XMsrQ&	E^$2):5i{7Zer$kr2Q754J'W.i>N:mn\-B}PV,I3;,7A,PxpmAyA8,jz!RAK|OG]Hz@:ln/!E\'7a1hE1l/rp<?Vg
R?vO6b&x_<#YAJP;7oY%P+4&`CN-FV&{0$]zINeY(=}z'[7h6AME_,hh{<R Uw-"6p6C1m\JuO7}[~w;8^F]u4WfSK8&7	Fq|A2)EH;|!1vn5;hWKs7*I9zg|!VI0W|ykA"8/ZcqYr/}1s%G6Y>29WgQcwhelczuk|.$rgJC$l@cl\_DX	\E7 y[|: !
a*H^fe3f
$5DhOzG56[nA\#^,_S|J>X!kSZ d7WDPP)ta&?3EQdIMJZl88AF&P7G|Aoy}FQ,(j]CH(W#aR(|[b\dQ
]aS$Bv=_L+(9dAlnX}`"OD
<d>:,> kAJ2!(d^b\S,Uu25z	p	Tx8Ss8
+yOTrj,sDNt7XiJk`+r'XVh0bZ`>-8-';QG}gpqIQB_5xWrTir>'I){fp@Jq%z/J[$8q)'QftyR@j) %tPdkD)FbEw?)p |eXJ2@e[q8j<dHcqVy1<ic.^*rAuqx!eR84
\No" !Q`	i)C,U*7`&A"s^;Q<)$p5i$LKs$j8  Ux*\MoT2iktQ<nYV9R`4ZfEu;4Mmb*RtA/wr"
C/xkKY<[2f2Xo?#@Jov6$bxQNI{(bJ_ptrhFby2yN(uG10+n=T8};og3t4m$ GRed:>jN@8Eh%M{Q&D>;G<|y[:%4,a;DS/"Q-peS/bsG@}V)jOL\X\UL!cMNJ[tW{Av!/.ZY`E)f_DVx(|Jju}@$ 1!Kupr/qaIBkCf7MC^0:!nMeOXs]&g{9e]Dl*b	wMd*)w/u^j-i[Zu,%/W)CqPyA	<52gV4j[.gpT_;eg9+yYSAo ``
Wgc{n`B_q~2RB{x\8RA1P2|e$|Bb` !RRK	$"q:lUAkM@}o&eq-p8qb3<riO*GZjP^IX]-L.i+N>mGEyRxSg6*}GD`tsWU(F~s-KK+eY8^o>&D?#8]4~`_xM!!{fm6
"1N?nou]-"'73rg\taaaZBHQ=)sMa#e[?D;vs'b4N$b1HI]YX4)\gBDkY@}~6>9RAIcv5zCC&*kp8K4e\1Y l2 xf/'jPW>/	^]%}S8NW.wOn5)ehxw.4uB
~2
[m&(@.LY;xcw)W}+Tsu(238y&Y~pCCbW%,9<#iuI]EP-:A@	4W1kOW>y*m^q-$EQ%l00VJ2Km_K_""zJ&8dr	Ro$+sV"vRHGx0,W&,<[TH[?'mxGB?goHUmo7at^
wwC3(gN>]
,T`Y^8:
b}~	0kQ?B:'#Ig8bj7.'Ao^w8JKXjZu~p3x2g	\u'/0a7`'+ "gnsBS58 ?hzL6u(85,\qS\3ewxKlG5qBgO/[3%5A{Xy~*)TxQ4R`rH&7ntGE5yCvQ(ce-Zq%p11 C&N5=>Jmn/D0T|g~@-"oVpf$7G^m65zhQMjJFJgf8m44pDb'h,zluJ,[R)=kUao%#.eZrDj71{
J;#L5	&O"}Qp!E{QzEq0F7c$_N5TusgJIH{?7IuJV_^_fPC:3UR0_K)%*`5iB[Bg|e(*2<TAkZ??4/UO8%6i.G,}+<>a^b0GVw)Tm81
~E}rl;)6d:L]E#k&,~,pB:KrLqm2-7CD%1D^Db[+kZkH-a$Lm&`xYySlH
tn/P|Fr{vSon!F^Ga4n@
TWN{nQb3kSB@=%.vtiea]NFK?M6^p(xr'EU{3)0 no'N
Z5q[O9Cz+c(Pay:8fF!&#T.qnaC]zfxM+<Sm<69gP0Boh~Bl/APQ_AP;}u,=1$]vMnRS7^k`^xoAsDbjDDt2g)caY
?k;\~~C#piqAE	X"nG]qKP	c;;UvyKM}|@"3)y')Z-+]!2~&
$H:#t|?$8B#vZ`pP0l_h3'l[_Q7~olF;uEZiOW%V+l=]_4AFYh@ c1J=nd2+TI#P\MW5IMHZKfC++,>:#v${!e3Dj[ auW{#G57~w3TyR)GN#Ts{'l{Wx?Qu<oE^hwRj+Qu
w9ofW5MvM-aa`,n2sIp0)- %`_N?SGoo=J$vK9|sacbj#.],Cm)V=MD=7LP`A6e4{19"rzy<~Q0<\y?z6|JH}s7p_'c1b2hp9o.b&mG:!2wkbkvM'zw@'
`Lk,1%RtcGWm{En|@Wekfakh	zhy"mKr}!Pc\;SoK3h/dS>P\Z|vm4RaAy@T[F".NSa}_#QKI6gKrT5M>I*WVSlNL\_JC#V9%8-Q<x:&oM%|Xl}obj!xZ(B(}ctHdz@c0}PDI|Va@b_s1v(AdDRs+~Bg(>HyzpC
1fX2i	MnTDKR^{&|Ngipn:qbRcf^jy$[G$d@O4G42gNAHn"8WN*&Q4^G{!R*b!,Q&5;):^zj3erWDq1```%C,BXBT.pH2h!zw^KS1SO ?h3X<O<iZ^Um\D&1}xvXb&-h=~e5q4I+Eo|R%N~A$
V,+]tgEr|M^6`4Us0B%BU>RAj,Rq@-n.@jV%o=\h`R6c:T+,m3`!VlgV3*_rDEqn2VGepyPSf=.8[X<hDt+I3$y\OMHI<83C:6n^6@!GJJ%&X0p0Y26ev.C:A(0<pO&[Nr|4	MP9MojiBqA.0Yv+MV$"&WC!5CvRD0zfpQHta+[U'KA0`(p{Ze[khh3gSa#wpIi>PLL?ts#%a?+o3ug0wbw`FX`k)lO!B/IoA{jHr3co8A+*7R:kl_n0x!M5'( OoGI>&:NfYi8EBvg'\g^6jrWc"d=%Q`/'R3E[flX=8^@  >nBI}3F.,X1=pHCJT}m[|2gcqP:YL[|t:y.d#Z,BFwvq\ +bw&vXw>Fb1G`E:}L}R
9_FD:;ORs<L@t/#>U}{i?;C,adlDmO;PK%:)bciM$G	
4}^kqXP{jMSXn?gifxzIG|Bxg{g}aJqTM8Re1Viw3L(:M8~/W[i%/6.ItD:bD`=_0s^5
N@n?n6sn$'k9;Vsm.B;/g7U*T9s/5ML:2l=^;jX[TWQ?rN.`tX=:vYvh[]X)8+XKZR{RH s8?M:%9{
:jnsN@/uA).V4{Z'?{odF^8Ge-cdfU8#Y-O)03x>VR=uH:{xSxA@lrS+37&k{<R
lTHPLH7T=<Gx=J;76O9*o-ewGr!>AI"6Z), En`B{b/R
	.?IWJ'rC_hY*oM6^cW9@?r(&Q"xT3zl`J.1=CjBhnOqXU>Ypr+^HxE.#*S,TEj^Dzy;Gy6_kP$cj[W`-0@'}
#L>>Ed[K<A[,p+_1fT4l3#'CA&aaatpxlRUmAGbv|3+(_ULS^;4
9vS,`~1E/4v:?D\~{r<VPUyzV$Mrb7 8_<bBC~!TGm@!s9,e4=!Xs'	G[ED9rk()']b|{C#y|H|C}eJCZ!l>PbJ=0dd7G%h;4@a]j	Vvu~]oVM`B*f}:~z?`p2dkP:?s)W~FoP	BS;#@@W6k@$i?"d	Cr'(;9waRd6Q^-41WAg%:{]nNy=krr3SGMHNECS,N\'x92cFO1`"s?C[?QUcI>,Y1	NKGqrB%)L	ukep{3YN>#E1UA{V!!Wr2o4w?N]~SaEmPGHkbV61hqw=-nT	&KA5"6~+B}\rOcUN+3'd<}b4gWU`IU6ed,<=\nB ("4UF?=uH	Wh(A?Lh{DulqYT2!U	2Uc">	<21MF7ivu
1>K*TW*sI6_iMn}Cb^o#DW8<[emwf	Yy|Qyf5$rk|5KzuJnv@ aCwT_A&>l}k%>~tv8\]D~YmaUgG5q0s 4S:il=]ly6+su]_L7S.P0A4'P3BGpm2y,Xzh9sQUi;>me\^bsxJ8R0f)4	U)1H8=7B]O5Ie0p6EfP#:2/nAL0sR|A7^&5"}(u!7h={(!S3ss*7(e=S!:u^WNKgb`H(9jr[*r%N6$^|fZW,M#qU)1`]G(MS30IoeUsh;G]Zy_HVj^73rF|_)wXCzYeCLbt]bKZO=l%;L%sHuKRl-TnzAHE|KN C3.OA@n0{NS"GRd1/&.#q#I-nQfih]"oY7-#eSz{>lK"=^/B/sGV1(Ybw.lNRFXv>,F$m3&~}[#vY'd&rgaX5)_P VS6pJEqff%A931i\G'>S'Z5?xAuaJ-yE"V..z7{Br-<)10Ua)+,u)8'68oXZ+}`,sTpq"z}Q7p`}Qqh)1$G~nHT6aWPe,`;$']ip\>}^}*U;~nQW~\h2EMs*wC9$\R''JU3o*c/!Yu#xu&gQpB!U	Xzxb"=<!IQ^d
MSW0hF'B-?
HQAW9Dca(HT>6v 5t8n|}pv)kF^]by0+}"Hm{:d468mui^'\D"I"4KLL=E{kdZcbYO/)qEl"	+P^GA|R[s(5uryE1)~b0RDPN[mA?;$$}MqYuP5~3Cuq /u({ild2nJ@oWmt2;fT4Gg1>o|^H|QpRh!<x0R/onzjY#yg~dlb:0:S.RI#WKYmEA#A2u"p^fr	[GX~H|
@5a(Uu7!J^i
lEj<YN>mQ+NT?7=]zzA9xg	"	?A%!RHRU/E4,|d<+J_m:W*:JBcJ`yFk)(Q$=4qbSQ> 6a*ad\ZyHAtip{vIlNJKGv+S2()eCC0+Dmsh(L/0[7MvW[j^;cL6,gwa?k:uaD`<:)nHW9u+Sg csFZS{0kp:,Mn:TY[j7`UUsoU`+_1c;N0x`XlFn,rcI-5)W[p9f>C`ClOOWb @.;k0Wym4:(6a$K7tH)a,6N6GIjE 2S6Wp|\K!( Pt `*H2^m31Cn*~M<IdmLay).Fr	
]p'taH+AR-0IP%4ptFB/Ub$S2'f_
sIU)st/4N[Af=E
km*='o3`s(|Ls?C:0NQ*$&rIid5,O
l~0fo' vSukh^~m)>f<GOBQ,1i019/
),2&Z?j-7@olU{5r=&BJELG!b%Q5Uf\T}/iuBCP6y;i4_h,t\N|r
$->2eN3Lld1{|q-}K,wRm2I#)HDsS@~h<k"lG)[=<mZnBjwe'.P^Mi$"p,`}pyK=$zIh\?`?|NeVVQ8%f},TEg$VBhtJ^}h9 eG!&|R}*4r2gLwhrj{#L+RKzfyD%3Jeyo|VJ]%QHNtHJ5`}S}_DGhiSYB\#?ArDh1U_Z)@c=aa#*""T8L
 |Ft"[X{v`?ECN $Kb/Zb
aW40FUv: 	`xkZZ)>=3TyGw.A&)35HutyMnjzpLBCEO\|3E!]Y5/V.CJ_aRLANVsu{M0UHmwI?T(=w?*jYn/!.mUmdIolVWZc=#|D!Wm(Pq	w=sC	],?&"Z_nJ]N;dQ9qBWQIgh1= _:9@']xQ0os;'6Zt]QUx}CTgb@Gcu|]V
Ll`a1R2}ex%JU9_e?-->^GM6]8?+0/e1'E\g%!-cjU$TkO'6#p^,wdnoc.!L'yiaT+X,utM"PVzgWRk8;?@k_"rYY('4nRp^olHx"&h_}6d$4hrd$q(OK6/?(>LicHC=@2fTdiV|0^'xkYH/b=`yU	L'r"Q/nJ0TwFv"+jKz@k[[Qc;{9C@h/2+&eNi)j"UcOOdZN&=h$w_X+:[Qz.g"4M7?2sxJ:0(}<>Mr)U/I8_O!'5G/H@GxerfYA|L+fXAHuez-\<?Ll-k'I*a]jku%Z]%3$
/<7:_3!X`}kBb%GOX}9ULb)II(*(8j8h,N9wa`>m9jU!R`gi)X^qAhvgdA]@$G{&Igmue\q$jpg,9?QHg5iZD%Wa\Y32eldPyrQNUc'6teln7Qk\1	Y
o?u"O_\7}-]oF`D}|JZ<vC
$f?nnb$.\4-/H;vk~8}kPJ`?uYpFV9z^omqF%zP@e]A":a,n6kIdO0}@7T3v$Tcofe}q@H)SI*qUnU&$}\X|/e.)?`17d<K=3121/QCw?>w11V[@,%Io	\#
`S	<_ft=t\!T k]SOYhm)=/%0Cd0Io}H$w	 nc7Q h[&i;>Q4
	-]G]tD$?0F>dDnW6e|"9PY/oF}59<i
	-WUb@w:9#
)/eZbZz90D_4+Q#;]b~D;I`T%W&7dlvo?^DG4<5V,$ wA^j[D,@C	5`CI9)i@my9&t1Y\%C_[4N;(B=!gM;:o3@	,X'Z;uaQ\ti,_/Bx?8N*xcFSngH~?BHc+jzndn{3a>LUF[Qo;J{|s.(Zx2#=6/8tOYM8REK!->zZ?qI<Kb%Khb8ii@yHQcxrfL:qN>m[FP/a"-FvR_S\=;Nt?A
7REqc[T%Pk4>X+;3ef
z
{|p"8kv{1k;E,b:_v..nFK`502JTn&k*t*[b3};I_$|;zp}%!Eg7-
_3Cv`5[`o-#4_T$/iG:.#DDg_."b,-NI !3@6t? [F7AgnL7{XkdL7ZH2Y%b4XdwE/A#p b`	%PO\GXQ$	2xcz
aMu&3t6ej-&/C:&GH<Pf5P92_]zPtKw:Hier,tSqr/\"?veI4D-1?jf}eOY=ngiqH/}$"
V,mYh]Ud5P,67Ntz_bRBfj@6p29q6s}fsDt{`e`Qpc$\`$]Kc5U,;cMVJw\6Zy24NrHB94WQ>djF(/7|Y,t`aFvO;D>28y	5\m>Mk0t_r5l&syYzE9qfQh\@)wAy4p!xtC-R150Z<J,rt~^ q3Imk/8Yhl-?q)xHr{c`Adqupx5pQfgLS?<1]u6)UDH'7%d6A]hG4NXj\|iVk-?<w-ME4Ou1HJK8m*H"O2MVdr*/uTlcx2-)sRF{v]L]QkU*!O2J%W{Mj5.^f
,\tas'@}@U<O-0lh(+h;6Ps[;'"FI9<5~{scT`@\?+9g0LoX^fQt>c|w]VtahMB&GVB:^:J7LNyO@DZ.UqT|oe\%(wy,6 6-Yo\s5FZ:DRrL7dW#_Y9NT>"j5iNCt4~	}Giccz[C[*"{{_b1x@0!&G=F:f/AFt-@0
sY?Re&LA$:%]5~50#E}2u$p^zeCA-[BA `i-R6RNe%E!\Q>EEUz	k;s1@twG+{#T bNMG7Zq>QX"m'-{x	jq~c0[On!wFKj;J?oRY3j?Bgr?I`|P!?cY@SRsTjX3cZ4ys}DP|qGa}kq"P
1C/a,'B}k.BzgV$w5p4*jWhhe53l5Rx	4(Yxw =m_Db+'+Cu4bJb	a9pQ
z<Bf{z}JsJ.|q%OAA[_8a:LmY4$\vo }6N!qEi <gnXKg5 s9N!S2^-8/+-I0BCdU"m&E&6Y?# T1]7Up}wgys[R&63-xi&Z}x{^{z[6 :OO}73/(k(^E#(+!C'>QMa12yUcl'347oc;7<%U>V5f^NK1riMasL5(OhbK9ph;}
!f[)_'zLB9a|i$"{adC(aBl_.sY:y0NQ_l4%WkZFS,XMo'm9V|79;[B=s=V|qmgWZa!L_4k$zt4]DnLnGsn.gvS%REFe1@8W::/AI("	awVsFE!Ew{:,<i&YB&C7&wB"yN'GZO^PaIO?u>YpbLrgy6K:t8
nZBEA4jd<\c3e-
#EI]c-os7OPn>zm"s+B59cc_ap*y3V`h-R~h/^?D	pNIPNGZs;JEHETN28o4R+4hVhT?*G77_1lV\
jPDr~@=Fp8`1&$saB1ZM	K_p9;l+x'pMs=;+x>!r"\w>%8'u.D?-u(MaWw-lg|(6^Ug1B6m^S)O61,GgO}Q7.c/4(#	8lWk$nDx,$l+H'2W	V;'?UI4y2C:.mPt*.C(<XYzP5?s-f+{esi$DUE|kDTH/Ix/<aU kYs8Mw2(WC~7=tew|GRu6qp"0|'p$X#V	F;D@on0B*$bHzz9JsSB]gs~J`YUS]aE'8G!yy%y 2dnaB-/SsFAk=*n,O#{Sqm=6?`g,7*NszO9(K{vAGb_<%BHgFh3[9^Ef/vU76#db*@-^co'RMe0gbwKmdP35ozy_G1pO<M~B3O?2Rs_sgb;r;kQgNU'<7;6OhZ&N>Hjf@ndS[)9."xw^/WEoy>UE"/Y	s|J!-=f,5}b0VW>]ZOSz{X`E>0|.i"/]sv<1iq@_J?t\y\H`u\0%NB1..le1\W1m=9JWC)~HD1TfUl@@+>%Q%WT
as?w52QLRQh$|=l5"oUmGL
Jj4E&{i<zXG?zu[*4jF_qc4d6n8$
P_Cihu	u"`x*%kTKkp?FK5?QP4Of-{UlB4U<8c({fYAkW|1)H@^53`LaAmuI0U~\~/OR@'N*D,&%>a{KzaT/sD@9mwjZe,o]}T;u0+syY4c"c)M/c`b|$2_	ivM&GcsO}YKMoRUhr-6u%!}ldn"wb$|:xrF!{\jsuHDl@}(Z a@hk+v^OfXCl+hCM~+6?(N*A>^s/eR1Xc-|k> [J2xpwf/iU?v_K!m##'U *"pQw+|
R`vgy='M!3wU+jmvq0y)|AE^uL/zFN;;CC8e|yE}:gf.FZIz"\UuV>*"TZ'Sd*s<=zl"`$'MWc.TfwoS7HS=2%M&[u**>pXs"gn<]KK
,m1Ydjj<ict%jU.)6}!$pL BBSHTN.N0'\[Lcytm_Sdmd|U@XI	!+]Q{i9z'(->fzTl)PV*0T1=L@'VKqL_3XY!K-<"B>C]b8$n|R*DKa)[Z6
'HbAI(5j(`Wl_,VfVdl
\Y:p1`0.$JFZ9kiWfjCS~o$;!fHL6[$0LJhiq	=t'5~"
fUJ}{?j..S>@>dXuZp#[*pj<0p^v^*tJ=r?g*<	>@M(qPng-mx$fo?qc?B#MU|#}}:C@\3YU#\:24TR	C\P0jE$zaWx6$kg.@X|5~8zbX3'rooPXf'WkF'h+O_n?%^A\f4Yicn[eN1@'6P!F:SP] Z3t(N2G pv"e
rvE.sT-t6,wnDEeWD$[H1rrbWUHp458~-*[sP09*H%J,[%j9p_HFfAgm"48hsYK9*R^\|E3_JrYR@p'3r}zzsLdJ-]rPht5
s35@`8]jIBgdO\"JR6}FwFO"ab]Ha'z9>qeoZ=pGV,@a!8T(,sX->aZvz[4R%bh1J! HJ{N(T.Kji	#Zbz
IH"?=a4k\0vBZ<ZcPus*n|:me
:sYa2ChD&t2pnu	l4{nDVqeU+_7eG-	`O$Ijx"G<4lt)Dq?3QoeMV|4V=	S\>;+_;qo/3H.ilA`MmajH"IEYXR8]),mOlVDo[*`*nu9Am^%8[X,P;bghaxY03Jlc.rbiyHsR*,@LhGFl}:9GryGVPe#ey?l1-:!f4SFI_|-i1  PTn4#V"\'Y$1EQ*.-L'[WSTQduEvLTD7{YDm,zJgFQC>/d{>=HDQ1HSXEHH_xF1bL.P7j+0Kbg,HJ4[\xP4.|X@AFgu`mjx#,huJsM3 AJ+1>X4iRzE,@ 7s>\1"Z]=9	:'9$	zH9W4IT	 jQo:N:DE:i
G;	7|4X+vsWI+5vG:NIjUfws83lm{j6U({Cp<enI8M@aOwhI>=C&=yQhM={)!"P(PG/Kh^Ok[UcB:g5fqP57L+,[S_	Yd_
HD{jO'[Zmwa-5JT+;!wV|{iqK`Sb/(BvF[OY!C$*y]u_d|QK]u>^ZdnR'XzClv7*f`GmN9W/0R,&?@c2d'eSv1R9sF"hTkD(~EHPCObz{7s!.oBe/L(Iu_,%i[{xNFa9 kw.Ay#+#o+aBj,:+naZWg0K-*DhDk.*t?ecKj<:oMjpbG$"cpW6J
>#w1DJ~ZWp%04^5Qh: K?'L>!gH%z7DCi4V$d5m`FVxBzPl`.@.F-kC_VO5r4f2"y8lc%{x;X
s\rLn~^LP`9yxHWY`="U4b108;2`<Qe8_{ Z>8&d3*PN&</e)*r/e%\,A"r3]$\@&RBCay0LIBGJi0k'*+A5o~XX~&|TsjL/+!igTiq4:WcqT6(^(tA`c$IA(0AwkC:rc} Q:#a&<:We]t?t&["55@xJ@jz)Vr*/S/$8B?=Ck(kBEnX%1VME!3\/hzCY6(R.0o'ye]'p~ASS"%+rijQPeAD h^0`Zr<~<8{T*;J&@iS"ZK_qI#29%eN0|aEe_;s`4/3WyP$7ws7MmS6Rys6/D=I2iMo\3MWbL3o>gn _Wwtp.qDU:1S99f,48==TePtBbSzV}dsXB&orsT3I\+v4OS5pk$T;SH'-,Eu
E*j<T,B
*8$xNQ#$u*^bUsF#	.wE%>)~|2=nmU"fj@TZ,sDa"!c$:-}2X"F\DK6|P>?y9q7"q?v7BIb*I_Uh?2
VcF<{C?E141{hUp>7nA.8]WPy;
XBW@h]`VPhT&Y<,P)a]i?u[6ez[%|%-N>mxlB,)>[U">V$69~sw\+I]!{Zy51koUbD`O$XQ{C~l7\-a?tn+	'U-N1Tu8D>fMp*;[IhYB&h]w)=0t
nrIW=k:{IBCz!p"Bl/Ki*}A@U_2o<z[_w!ee|g<x,7/_L_h3J<jc^B{0^\(?:6AU$K+/Fz[x#LZ1~6D$X,"<f/(xx(q'q<Kr7)t$zb~PpR9Pwmci/r=Y|cRAQ[	0y'fXWPW)F~|t+
=~o29;Z#SNc(I*)?4|iX_1FyYx|FP]Di!a*8&on{d=5Cg4&$WCy(_J	N$NM{NFUU"8C'k|
iy#ZPZb1Y89OVSPQ5AXcG-wYqUlb&A{Sd[w5l"S}I7X9&5Rj?Gp^	S&CP/a{}Hx0~ctk~=H	@?K9J\&/+z|jGHd[;JUK:qu9SqgsdO}"gUq^?m.QEO`c2K#ES/	vDKwH5x\Bl8K.TX
Cm%&y5_,y\2w=g<IsU~T.v%>?\6umXW*u!eaUW'iT6W+JW(osQ?!zM#Ywf\wh80!,B:C{&$Oh~25\PxT;C0`Q^a],+gp`]:	;.J}z6xbCp\7b0vpJ+=irmYHK6Q
#(<-:"4U;!ll,<6{%\s;}CGO31/}gr?_mnK?m;BV]"*1~QSgcBYMT@Yf}UwQ	l<g@EZXOJ'>kXK*}.Tq0LDzYby}gdf_^ ..`erj[T<an}ihirNG'["(C.Aq>5e?)9_.oB6FW>X	w5<!Q{UyX$z<L~ucLdDe>cp8,60B3]'%mPaX~^BM|O["2&#]}X{y'@F7;1v&Bi2TU}YQ\YDwAMV8-mD>}z[z.'.l^9O\XQR[vXF
$<3L,h!tM5.:iyi<~WO-( ]?/ax*".AG2Q4Iz_nnN-ydD6K1~"9Hy<.fc^IMdHjh`Y^O\b_h*e<fZ8_uAmIzA^)+z#b9FAr^`;AAgN!>/9c*
nuj6MF.f.\*^_zy1(:MwOTNr]SV
(?3Zz
|AFTiA,dnNnRX+-LOsVh%zqhFWRl{	ulVR'/t8;M97y/&}/cSneLA633M/xu/7v.~Ok3^&Iok;"){!Y:qn#m3g"\0}Aq?K@H+FhH?b9pH}m`=(wUpsH6W(Y9 cLN.04u`v:Rqh.rb	qQqkp4I!V1.Fq}""r!#AD[0ljp`n1 k)b)u%-
L&6lRXI /	$i~"uX5D^6.P@,c4G{I%|KQX,sn@*Uqa5t N#vYno_o{HS"b@*y$zS4V9J:	B[iW=\(L_dpl2dS^fc"4A;SI^L4a"L;|k\W4x"_}/T[p+nFQQ$aWc4ZpF"s>cdW|0!c2tqug[,$[Pv),kJz_'-O!|6J#H6@g&Mz^CWV_i&|K;YDKm~Je^Q)0G,n%R!2b=*2|>Yoo0D'5&ayD
|(MxLG}6h`G>I6jCtBX,)v()$#RY;kVj`4}uy+HNcSkd7[12.VQ<k ",do-p0*81wq:c@6uoWl9H+!|\689Q
Q)f*0j<$#qNC.Kj[k*u`R:98b1}ibW+8mM6)A	 yO)D}*J5&S&BpCKj3AHe+6%\g^35HO^D6PeY8|7dRNYE:Fnk3is!lhLsqmIjuiAz4m8Y73,~!D;g[fT.H()T,[G]{"e9xR8U1^M`Ej3m%ZIe"!+qs?u<Z,K-t+zyK
m"(D~^@z^4E^'PvG'*	?h hL55vXYt=MN6o+M4tomvl8e{WF1sNTveEbgzKn{@t{u36*\/"7;o3TOD8_T
EQJa\%g7(].+d0Um!?6Y/BkQ~d4	*zE[q=	8{ts5#)*#JeQPMMx(vvZE[kjD)} y{vPAcr1=fxV,[KcZy%1?"hje>iHU;etSb6{|X 6o":O^b	WCLp1tGGr3&wyMKt 
ZfZgqS3]LTtrQD~^joFAHWm
qfuU#zEw6}LV*`H<z(.eG,1[r9b)1xif,-j>5N*'hUS=mNz~I&X(9o<iC@7R%7W:8\!Ys=
Crk*bFzNWr.Lz]b4"cGN>c~q dJvUuNahR*zW+:(Hr'F1E7I2}+|1"kbS
f96YKr-]SQ/_'`]Y4ICf)@O|v.>PKZIlQf,%d``>NmG+?u,J
1;Hi]Bh=5pmm*tkrX2""<QG`F	C6wK[}`-MUc|fPT_Mr?_vT"/eLLR6pR,`cAP6b=b CM	B}yVR)\d,WBtJy#lt4b"O&}Jh_,U8QD<P^@Dlk&b&9_sp.Xgni|h\hsUz^O@<[6*a,UELTD
TvytyX-Z*e.:}')PD|u
OE8V~"(x tQPWP*+t-kF1Gz@LA{YC.ku*
F'(M@4C	Tqi,_FN&4]8c>`A/m5Bi'\9}P=b(%VY7ut|C^#/-{5KK;Y_P]-!)8V3yGM$^|];p>&UL}]}6W!i>~)>	POQV87uPGstI31{X<++C<U7(ly!z#AHysQ\^=GE1.>(b_yW1<}C#IN~apx?$|3|1Y {O&%PJ>e?gd#Ck
3yphJ:RTQqU*RfTIFy	1Rq@TQ70WsVOHnt(<|e%b3#%c8IvB47"R%L@CbRP*VaB)`zhDUf+n3_'tO]q/_'g`:hI8Jp|)(L^
QEiH?|/Q)J.l.]Gl?itv!"JRWf|l&edX{Rr+$.9F8IfZ2!F
hhta	E]6(gCGnT!aq;o0H7K 75|RXbn-vA iu^0~L$ZyA1&t_C-7$lt7FK4EH8};X&e0R>kx*X!@R2Fk&"P8P9-}NXCT3%)}~@b}8cx[/.q#'T8 4a+,v2siT2NH	->&cN_Y%>4	*?(H 8*e%b8Bycjf>+29>w+Y3/3du}LZRLBx_hn3__mtI.zt"1P/^y>mH[${("DJdR\^o16Y	[[h:LYVBTQpTV0:
_/jWZa>BLQpPd,zF?k
!p$}wP	L'}<XarpU8YOO3jsHr#L,-I*HQ2t&=7"-8}4 R-%{%'l}WH
i=Gsc	.c&{D_|N`-3dS:I"=UG52J,A{fz)O4,JX zTQ.ey-s+\	)-m-!#2N*zD:J$aVUZE?nTbH_tU
o`E}!*.)4Jdox<[H]U6c~e W!Wqxr
@7sXn$]*K2
fI{bcwI.H3>mGC3sk{vOY#:6AG
y*&O\+C\#,<*?'#UR]4T*A]/[8T5"?29=$F^a2cD,KfSGbP0=n=bv?X%`58K> hu~=2/=`;)IJ!d!6h<IsDj^{Stkm!tIwW5FXQ_^3PaJNZC$ #<tJ2+^v#	0d}D.Gqt**>)vo#|"Y':.~<O	]%p8ES|7N8tDWb]Ad>%e()O|*W:7l@)D*x=b;3wtLtl{hre8;2
35SDer|6HFZ({KqLKU3zJ-4v?Uh}>x_+=kjo#\y-Vih\8K4a"	~:n=L*|p(_(y"0a/LmR]_&D	&VDY2!zUc?82\<Vr<_IIm%#
a8bMaID=DEjLO(mqw1P\"#u]"&Ro~DVMQFI\Z+%CMGP^d#CcQs|q/nP)P#0wUw>kg.y2gm:E$d1JN\kN'2,/Y4Jsdpk?Ii)4hT?xXe'm$),[y,-UXtc LxOH>GH{=~&R@_Mj<)|MG:_ma|X),$RB%3BV&>WmMAO	^!($oRaug5}((t"=o9_IAZ,w%=LLu#BUO)r='5nY)nC{p%`	Gf7A balJ)T~,n:;9csAV?UMocP"Klv](JtUE`OpNJ*Pb3"YDL<b*VTsQg'^"Ub6+x_8Jv4,+.UOch0WG\V7W7$RD\QC%,w_jVN&M']sn\
m#)QDqAQ)=B88(Z2UkNeb^{qRx@NV3T?N*W"D|Y1e\FjCY,VXCh0"
GU)j~6X-4bA?rqM$8 Euneu^PoC!sf]v.0289Dm@lPhuW&\6u*fW >UHMNV~*^Ql0MJM\a
WT]6!LBfMGx@#jN:iC/kqDayq_+srQvDvI[1OT@#_Ybm:T{cjPP!EZ&wOkgZq6#;Nh,v4ei0tx})_t.v:E"7@t-I2'OYs)`G}#RAr~-Js;tdaow)N7r=0:;6r&Vo,O59C_\G|gx	ocYG@=HI#/Np1pz2>c*tVGIRrn(]CG- )geVik'RErp81.[6Z"9(/'5~P\=Thq#MZ@qXVFe|M]	`Q=4NU:y|*<	YI]:y~._<(TZk#i>E7p1R<tY&{..!EznzBQBjj:'\0zd	X|~{D)ATBCV?E[V[*86-FkryCylXAi19[C{fo~DlX@`s`"]*DhU(unH+nu3)'rvGX gULM6qzGzx}@o':uhlB1G%gV;_b_VP/'t_f6{m<cuPgCuyE0LB<=c5UIC_Gm_gLv(!t+[U?rrT4~png,LDox2.['VUU8f|;F	8|L=:Nyy1vL(es71:x(plT)VT{9tKiI6hsryl+fWx[>F| IZySOZ/3|x %Kj-R,h+FF+d14Oy'zG9Npt,wz!7NsgQuzY,sIQclwDRA6mm=-*}`{',n?BiY>7y'.u>r'!@$;S>Yx4fX}F	PQj^)8)"PD82Ef17[{H`e*OlT}Ja6vFw\SGbvzq(ZAH
7bz2FJ67C1>S	)hY=9d.c}aOn$}0(]lUV|OU[<6:77:E48yf6{RL4J|Z?L11VsP}pudXzIH
{i5pb{ZY=epC.f*&MsO|'WiBQNUw5l@8EcY6i'&MAt{'"P@N|?jdvzi  :.Hb
U_j:X:M}F@;o:Me;DfWGm}e=(7VCu~qS}4UyPt- UuyThJ<Q`LSf\hd`R%+BiC6(&Qn??u1yq	:gw7CS$>UlXW=`LZJMF?V>D2FT7[0er3AmkS*?4p(+8|e#pOc8UTJ?SVOcp]ch@twiNIR75%S3WR>m'9w2eRgJp{ceM_v(P*(B9hw,,a7XL$mrk6Q$u#TTvX;6(H:3vqQ
GnUJu`*J<i*KFM;)	4vHMjAae=ee,cfX*,;Jzdxqr6[FH<SV[5jR:5idhgro"STQ,2+fT[JQI$wolscU|QJjI8$*,,JRp_OX{-W+X:uRdo8tAkuNR+r'/pzul#tq..h9I58}i%0>=/HSex_RN]|(yK]Z [_GZdZp
Yz4_GW)6Ceu~XF&D3c.NG_Im>5B!,71Wc-p5u#j_#8mb^/>o2X>![VzULU7bt?Uvn?lvL~jEO=IRvB{RN_FPuJAd\;#A[&\Yj.JxwnoYNrJ,Nw]Tt;"-)P`xxR(H6ldo!(JR&$Y(H8r,0sJi>rb??D/+gO$ywEzdEdyf}Of7Ppi]"V7k+-R\eh`a(!cI26ghLG5@S$dO33&\y"U=Ihgem11C,Aibl|I^z'Y!9NouVxZpOQw\$S^1N,[?:+}_R?)C!&2}qaIzwtU{V`G+t0$c4xM!8V#;(Qd-ez r<}1)$lNUuX}UvA`;rN.nEtd{P]pbC^MabX3]pqT%Yzy>tz{R4;ma_$l
rn7H>(k#XBq4b[4zlQdhxA4IMP30#|("2Lx`q14aY[br@HT4sR"2$-9B}v$2+_z!d1VtJRTp^)&dK9Ym,z1XyA"exAaZ,iJ8if1&QjFYBmP48Cvne9!K<j' ))Yo&b_kJ9iY$Pv-`Pw]jYA.09Z<gpe~'VV"AP
Q7O4#Or{{bEWPpu/x?R[4eb5>>pJ*9k&,(F
#5n
b}e24 3,![w7w/{(zt,HQ(TY'*m
9{{:jY>\i~-)$"${C;qF)\+dE=?dh\VYnp"Y$;nc	lOii%2`(>uIbu???f?sW+*rY\0#
rr=j7I<Ysrdqb}	cd$[Ah8p99d^)\DGqX
Mwhjsb@_P80G#@P:ZU@Rl*Oz}lf"E=/K82
Lg2^~"$`EVA/|p4E0,}&lta	C89ZR16z3S}H\]&+ko\9V1t,XRR
EuhT>qn}RB=B2^w:V6fKc|*SK
{<Ke!{[]I"(T5,X|J"fCYDi>zKZRE.\&Qx$^`K|^>T#4f0)eNm5Haw)KY)3nQpEF"EA}8dGwR`Ap-lHwFYt>cwpJ /jMW&Fg&k`T/H}OJTWw8iU%FGB;$];|Z$D,6OieX$ :NKL	$liNR|T+lwzma?#j gjYQS}rsOI(+l<T0o!w2W<yskAbV*>|Yr]ME#"*TIXQ5jLzH^)I"i	y^V,;t6Ef)7T]H5aBnh9D?s8UlK^K8s](R:~5{iBHrT!!fpfI(2mHA2P1F XFuz*|&.U:}c!&)9i\%7!,.;B'N#2LZ|)PuB=|]v=9E kFC&*LB9+2fHO*!]vWy/G[~&*P2X{bFu(p0;sLI3axh_g_u^&s;ITK;{R`;dZ'm	G?kSGzd{1zE=x8FS9_Auhktz4G>jZP	`[lDj9sWc7'(M`OUwBK$`x.	DlX$*j 7Un/8uDIjmQw
tbRP{rEP\
PQFer56}(+M}]-RgUr%~aUTZw,6$3A8#$lzCO@NG@0Wjp2Pww0_wcc8b[SfucL
_"9M{h$"TEUWz5|a<M/}Bapq30InY&MT([|g<Nf
 3]9kTpv'sr0qiiNfroGlVLI=
z(0+G4/p~'Nl|	dwkcz]aOWm-[FU/$l`o1OU_=ZeWEQ{z{<EA"??6DRG7@.E/yBV#d250wc'*+SZYl4}%+GFKR;LDEDPx5v<,SgHSmS7
z3JFrnl0'zY)\>t\mGZuUI<Z3\Di}=<Js^u2*e)#1B>$&3=4\R^UFe%o-0:}fm&>(ei#1d2'&FNbR4isD6J.)Vd?]mqG5793u@`GL<5!	w.`/ u{qg"2uI%,i&)~vbdgR:C*8P!gFKHZESrT|~YP]sp#GkdNqZg[hj1[9"S87)~yDx%osR&!VXF3HX.]G'3yP@W4^]-oEZpo2C0eH*&Z9!I UE"Me
8fx[.y
&vG9 #> C@2:
4^bx>_|Y+1b w4myR-_=wRz>iSAI8b@_l6s4Y$3ncRmH!`pP"MG5sYI2~X<$0k^3;{v5e C"8`~,D
q2;;2s;Bq]E@#Kp1]|2?=a4
zXXDskr	R6I&+F5_$a4s.el5nFGha\A_wROfVbF;}HAt0y6-$ O.GUBRFTKg[b;^J'b9QQtg@'@m1_,;^zKset7MNe!>#>lH )^o>Lo=)5Jzgr'lHNS(3QW@if{`zD6~k9tnY[KmM6{sJYE11mbFIt^/)TvRnVJ4g3P8sogFEzMS1krf,6\aQ3[v!D$9u drbK:E_[i%qG1_C|PcJ9FX4	C'X)V{
M`TfXHU,N^?^d5"|$s\F-2-PZEq'SSian)4oqKkxE`8V)zN=:;ioc:Z`;7Y^$$a>%|T*`&==C!<5-i'^M<3")WR*Fxl
r^wnUj~s_C8wg)c{M{`,}(lfMHCM*jO(Fx$Cm4~f$S@Dbabi,z#
>aw!%F+DZR]|$9I.UnAMxyoa_:Y<Ptk(*KR!G-</f.^(izk'wx~8LnA7*y@E_LE'H>A>u{=y }d(Ma)u2>cX@{~Bt8Q~IZK,w/GsugZ/U[&OV@=I}.%($xDB#I1{vPD`"+lmq+rbYbfX6{~A7Q|U4N>?a"|G"=0itnqsid%:gq0k43#/?<2u*o^S,s5lc0Jm1qV,+)r\6N[pRC&g+ [9Q~c@y)mc[:PWR/C*~X8[g8<zd+&UzE;Y8 \Tq|ONLl4L:NiI&ko&>zb;<|s!N?wlEU9	Nw]R~[<1(cEa1=>8swoRRnR$y)x2Q7|L`x

CrM?wC{3R?q;AU!	{:	$v4|jC)~M<goQpDvbmXD\N12Bj(k%6-\W:fp;$"D18}A@Kz'#Y,lJDQ9KextNS+hm!S<o^E=dE<_v*%/s5np1l6uO!*NZ"{lICkP5Lv2f^^T25vXLNCj#?0E`.J!T:-!i*s}!?LCag'SM\:y#k;rD\^#L6Aja:u7Ij9I*NY,TYlab6mmVtLw.4Hk'zf-ls"
)"x[Y0p$@VS'7V1RhLVYmDi\FKXR>GcL06YW #	1mzf3O!-g$8y"k/eY;DM%A*$oq2QPH,#HD'&5[Lw|M.ngpqLG0Wf5Lc>*d_sqk560r40uh/?J)LBaiD;'mFYBp`Jdz4zGZxvipoc j(k^ez.,OvP^g}.[(aYws+q(i>g(mA(i*%A-4WV<7\B)3fB.LUaQ,[f-VH
?ILPf<yH?]Mg|l\)>aKX. s-}KJYJg&&dlLtZA@LnG)C%PfQi q`VDg'eFCpX3?q\ozx>A{.\l\wmo @lDduoCCZeBf$s"pwh#!\Jdu}Pf!(qv4BL*f_kQ%r[7v?OLu
9GAPx2<M_C\2ucBwlP+g:9wcXX1\$sg[Nd-t<9#3B$nyAL9B+gaRuhwa\?3_7G:;jw2G-nD;0$V=+E'K+'1
"TaV%5Ml$\wmDTJ~<]\|'["q#R~l5t	]vZ!w&1Ic^n"-iBQUl&]MKCHV)fN]HfZ	N@+J>_7if_(_Vk\:m-E4Z(>4VI$sx(dmqL|q;gt[SGg	lm?oK,F\owkjv#%87`u/R?}_\a+P#r
k{'+O
mN}2[BQ;3})`?W)A]n\kRZ^FS)-Rb~M!2\?yQNN5~?Fk6FG-&1yZ5C?mJ@OzvC7nz;%8)o~pW* Z?0NlmFMP]w0E+?<D6! cDR)8hdbW8e[*c9Q<5O-7^^{)bJ66,
-	X(Qu ETzq	2'e>L*ZGh0f"HowShrp{yN%!atkV{x\|]Ji]o>
\nt#B~rVzymh[xryW,hzz\$GayXjK/VFOQ KY_r@DK1_\dw5=HM&j[t,6	[V.>\,[0ap[I O9j\Ng}vtC! _yGK <o"cA^<vV4Tb-DX5G-;U\S30*_-u.2z+G_%M<LtKog4rUT	(jCznJ2{PW#Wd=aWDGO@(j	Y3>8lKn;+A`]NL_Y`QfU'2se#-+OXt0gUSH;Rwr3`6edtNeW
SvJNzVU	pb_54k#@WqP@0>t&sQA3j2z#b,+l7DVm-POse@vp|_BqZ|T yIb.R>Yq4n/;PN\qu.]"NaY\_GoQE{,,[TET	6QICH+V%Vp2+Wq:cHss0)#|bGaDO!)]KoDW&V[V4Gn>"_h 'J5T
HyuAp y.X{xF^V
LM,xl
{|eUrSD"<3q;Go3yc)gcaD_75A8Rd5],uHr&_rg	bJt>"^I4AO|eoZ:I<lX/z;D*Y>+ZY^O)c$W*DsJ.M|#HPIB,t4S@:~CT}i{cD:Eeq7Zg99Pz~f)l,sudM'	[>+G*@ bj*.>ocr8'qt'u$5_lAZO5]]w5>F	]\o=n~o[8VOZLlOffa+3uj\x`EyON	hBo|7j0wNkQfMM/Lq>Sju(?(|F^
^~\=B`Joc?$?2-T4KXOi_PSN;c	M8L!u}>If]X!_/3K))9;D)3H[%<"dJVIYKQXyBSchp7~OBH&@YZrheGjs0x?*VQ^&`pGFYMDTnNGAW=?EojN&9v9de0(X30ie"|NO'P/=Au63cawJ"ZLYY0P/i"?}x Gzy76^6GrbE-3(c0Of=6S+J6
p]/f4n/!)RxigTubz:#<|,:NXP'RG,C"20ir.f8D}m2OBFoX/FD !2/-K9J#H1$_YQ#s0Eyf s@WuQW9a.xqb"-7^5-?EjN"Y[EE*OYR#H|Uxko%mH{F8Y<9d{[#-S)6H(-/)QxW1R2s<3?CL*fg|vKJ9]Yr@QbC]xYn"`%O[j d3AY7	J}
	8w
'?h)x~Aa[HeyL#p9c"bPNVn>~J^.g7*;91Gk;:pqBc48QDRa/7FEHfe@]>qOo_2QB#T=N'URN7\TpMAIzfHs45<8Gf0IKsbvaUxnm]M{e]X)XfqX&H%A+AF$6^+8L3ql~2B5-D7KRVA-Yp9?3*~NcH9FBAQg6`I&VF_"^^FV67m2uOjO0%_bLN$x)[*2@IwHR4dv6LI
-u&!]H$Fawh)bAc?KOG>xud#U;6+z3_b1MdiK6&sx$qkOcK#{q/UOB6}t{`ArBImE] wwK|0!6Li2]FJnW]K1iXFT.N`Yr?0f58A'Zn#NYzXF
$me6	aYmx'w#,i.Tu.zN?)X<*I"`B=E|F:,;MgV q6v`z:!mx@M/-`0m3|RZ(1&UZY&H;Q|s5%v'u<)w(/T7(sB]Hs*!H?Ms?0M~E@.*\M)xiUMK}m	I}l]BRNTUW}N:+P D+Xr%{M[c<Z|Tn}vtw=VCWnPqNa./2[+(O%\=dUF-BScP(eu5}zHxR_"{{Zo5:U+Z[Q'e>GI} _l&G\AyLMB'/JXT%BsxyY*LL6=XT	D9NQ|*Lzk T:E[,"(y.	E&!Iz
HmlS$z>8E0&vf^&HN}^Ey#k+i-k(<0*5xy]6,"SqasP*X<SI$S,IoC.%,%#^`Aes8]k.~`s#Igzm!,
iLNV37*_.>W]lkVE"p,P23'~l\-FNGu@fc
IWE5
_g76GIzd5BPfQ>
6`n[0ADU/U<1GbkCq=K^le9eVO?fU;_2}e7Jfn2TXwgFcb@'h_,:&g,/"[	$)M%l,aZ(#O'8x6r39y l6q~<.C6[o&"\9%w%cLa`0'.ktQ4@sjLi)ZEc+}hBglZ3LY7HLO'^]xM,7)$pzKbk#=159{\)Bc_lAPC~-}-vkYV{&fM*&n')b6@#soR:ZEv1[m:O,s`LD]_OcVypA"G$1i&4#}BJrALW4Y=\Co,FF]>\4Y3-.@ge=74q;r}=&$W,]$kiGNrxjXpz!nj4+^,%MDFWx+kIkk8M[XgW)_?~SKUmor*h0"dtT>@2\;#_JK*[3<QXaZk<2ec>9h*d>E#UMWuBy:Qa@U~&NxPQN4^%jN:9"x%980{Z{.z
3Vt*fF(v!/	NxfTT#{HV=\f^47/&NYG#HOll'so1Z:_NSVA"Z/4	pUX	;zj-Q,iph=lhd"~1&cC~b^O*;j1Cqkde8/3}DyAa9	\X)fm2T_L9_yR6
.],Z"p*toCf)2F1`b_H#7.W<<}VK3_kvc`qck
 AX2=w>h!.zu,=!l97[KjOwnF`rId* +3r;D9XV
M}]B=u;T^	if=k6RXZ'cj._oeM)2$8SyrZHtk!XO!#,a+)iU,R42:w=xHf{G!7Ep<E8;.>U0zf76J*\^*-a]pB0;c)Jz]Y|@iTn~`:;1"uRS<-\J
"V0NUc=2>jn>a=p1[26)ryD(!cM7g,	:%iJn#+cl(~fld	B"3QI.wF`W%fs(g)uLN%+W&e#Pz
c-
O:_J9/??mS&CR{qmg0|5<fehEF6kZ(ZcYj8z_Qe3gIS!ISS('-~8~B(z_!KF}&7\=:W4ytt!|%/"|`c+,^y!V2ty.FWP#=G)D}x~'de63:p#/s&J`0gn}y>*	eAhG=VY(pp/0UGbv#\I>H\'4,puXu) 9xcbynbh=FLSx
tO;A^<RU3Pzky/8(IqIB'>;+XDf[\NW^Gm#{|I	$mCEFZDZoK\~U826?F4uD|p4e@
EvFRwn#&Ur$xSWMJ/%v	=D[Mq7ki+%R?D!{?n|tFRA^YZXG\C)+/>9mA
Y]5V9u)h`dJNc$_

x/^h&W(mfiDvZ
bh6AYR/y/[`N#R0-NLLu|d 7*$sWW~a[%!ikj_imBCb=^7F/Lk.L/5z;pR}wcPL)Gd)?1$q'uil%JAl-gbJl]|MW	BZXKs3nNQ>4	zq`ob2i7>%Lq)?ptMAsI#;}Q#`Xmjc#W>pBO\%gr] -"yxdzXZJ3{e`VoJO
S^#L7'w\VHU>D.zcx-hc=MY@56BbRMehdiP.gFv?"zg9JvP5~UOQ]2{i=p=De,5!nl5+gN9ho3M[fx3qeS{4H4oje"2q?8+|H0r"7Bbya/d88XSJh	M3L5T:o:fvE}s`F9&2Cb,\n49q?i
aB.taJgsx?.#z{@piWL8.tfo\ng5lD8db~?+f'$I)g$]Lg;Zm_RFLmB?WRE8Sj*zqz`e#$>Qd~WGcC?5&:0BvWVpEud_f'MZ>h@wqJ*>c[lh{GXaATS9@taIV77a5@'9vn"a>.Wt29m7$UiaH3%2XY;R$w\gN[@@r8YQw7HsCS7y%M
4yj-!-\crHK%-6&N[GgYpZS`)5;St!s circa2^ud`t'&UMy1GC:tu! X?^]6Z/(KcN9q+$kLlMV{w7FF${G9vLrr{~j+Nd=/A2TbPU@$`koT/MV	xU.o9R;mt9-.7Dt(2"v\p+c?7c{b}!c)z=*]P %gq]YM'r^(M0!rddw,VtQZ)Nm<HgwI,#lPtkN2[h{tgOj%V*et2
|o93{gfgJATk{AZr=\ATYTf#i.g6#_k.i;|V?f
A:,`Q*F\KpKE:A1#lca-HOuz,H#DHg?k2.B.e2_,{[5b!(G22bi>D-32GA4bd-6Eo;Dy@
R7*VWNH~;v,.[i;h[Gx*w
,4c&g@
hw7A{.F^	d/d9$,:TE9TzJ	6XWpZikP>wLiP<~'_ZssB=xTJxjI(LW~pYM%zN3Fb?6z/_Z<q7X3Q	}^x5flstATPCzYyBm1Q
gO4Y`zj[Zl%M"#A
sv'6ERx#"	E+-C"5
}{&kXiH+TJCm;[zESf89,^;b:(D:kI67dQ,=(zK+$Me%pE.}L+t@6&Oh U
jIc%O[os9sZtyt=BPp|rfV~R&:\x hU-XD'7`_'J"Us`acnXi&*>E/o\|+&~7W S:M#mJ8%dH<pr\{b^M@1}v`tVn)qxF|Eqnx9p',_#.&=drkW5|%5S<%`e>Wv[M,$UN
/Z2F9]h;rV_'uYFu
}+6W1L2s@3RKLFj
o<o[pXmqzxjkB6/*9pIm9H7$IU6uzHs,SPIfGgpS+2/o'+{j]NI"/!:7}I_GC:1'//K	$_=8"2Id}\\g)|q|c~#sd1
[U>$0l_hE#Ln!e^+'7k7cbSP'VW -<-M4SF'Oy*axJ)E/y#_y:U1`+!Y'L5(!A!|8OgP=i-	QN.@~n6?$4LOp}/HpVt2nDsEW9/I6:Fqd,AT{)o] ?y.Oz8ooc>uSsl(wa<P0	T$C<my.aS"*I/6`Vy./g;o$GY#CWJ+8=(RY+6$d#;B]\Vt+=`|.RV~IDVlb&n`$BZJ?~ye\S:Wj}m_y/~"ozMsS]QW?C?9:,na>GttL6s+o283AO4qjoh'Nj!^RN[KlXvLZJt*:2a{?P6L>)YIcy@u(`V_tO_b">%&;nK,'>Y{ }/=hlO!rdN,zG$-)BuEJ:^~JPdp5o], &~i(fVk+m"H$bZ,\E)=@EvIM?D[N1o,r7	n[;r\O~,M'vLi0<%WR[q(x|gPZvxYEk`1b2-HB:0l*">TNJ/R|w^et \q?y0D0M)>{h4>ok8KxG /9H9Ss#fOKd\PmOVfp|b`xA%}n|	F~*yYVG%RmC,qrSK]nM?>mn7V~	{U$Mi)NsQ9c!Udb>B>kHb8mF'VgKf,L3]9HG[)'J[Ho63"t"Yg;=S@=I?NgA2he)9aNaWuq  (&@"$tq_R)EfH6WaP?/:W4rRIj7tj,8eVAd~tZ+_>:\.taj7TJcoWYh8I:bYuO7k.!s%B-WdER/qjpnXcgo6^^z~Kt}4glYbM[GM%?DZQ]
B?qCFiE3DN
5K2Sh#!FUooEy).2FN/T]a59\'wV a'5%|!%?0tI_'k\IA<w^]2G1&tJq\As*Z2Khv%3v$nk&hI>03l@m9"Wc_9.opc/ISp,/|UPs;#qF`jNoqgM~1AoqD|?#=M~yy	~j35a5G.W[ax[af0M1)xt88C1nbc6
)qGP/zW^\6c]@QvqG,)=&)(wrZEe'\vKW:[QF7`k86@XaXQEm\vL%<RN?;jo+\aEMSWHp#~!Vp |Ve0^/Z3y"1)<-35yQ\ :y@:71yB"",oKlD .-*Mv{wD:o'JR&i~TPPcwV7~lFdL".KC{&%sObxQWZ#\tg>Wix	%]/Ix?V2H-7~<_f8@<4[FmU^'F!Ot_qkc#kL6lS,aZy5,b{c!MYj*`gaB2h,]WN	Ax1zXx/][8`cSh'^=\BgYald:><u(wcL_zKG%}0w>!m<-tGVh`TZe!T=CZVXb(
oD9oF[#Mv}~_ML)ltIer_n6&E7	'.wP5Gd4eZZ}f"5x&=g;|gYvteRS(R*0uhIZ	~,7#F!q$ZR0W]$5MSc\*Es%9wl,F&|VD@!P]c<=h.YUT
9 sz&UxzY&4h%+"RuRI%z^t2+RW~tn3KYL(JA3F0tAADvHT
Qp(t%Y<nr,uo47huIeP29k	wUY|(T{wAw%BFvo*A)l1cEezW;?I4m%}13a!&DFw>=jeNF,<TAa)w1dw[%4XgQ3"leYLcVVI"U	fQ5*<ET3}9 -!lSlqUaVh	_{J47mYR_PB8OeCz*e"uu=9<MbY
%1''Z`,%c.D6NGkOo:LG`=\!i?0J9z=;'W*a5H"pu5.Ui`/-ygNDUt{6U=FSdKu=;LR[n6LUdLAX"x7uBp%K?17!$dd9rc8"17?-YV8Xip^,bYcIN|PCE{r{XAnu+xuwb9u;F^<J.>w7Jj'4.b
p&Gj <=pY`osa;sAOI[%H *U:_WnHb8!1oi|$ZMMg}fM{S$U0Kq4)POj/f,.jIqCyXk::Fz4bcf$||a"?OYqc~zMi6|c^+b4~{f	6Fpt;8QU.:MmvSJ:.v`8hLrs!IJ+c[wuAZHD
6_5O/dM1\~GSXm]wZV&OJtg	%kgaH3zum-hp42\K4!@G_G(q?&/q[ZxQI
|!6/be_dpUK6v|vHACjuZ0O+4}V$>@";<m1tx]'DZE2Z	|`l|x#O6}	zG:6H+X6'	-IoUq]m3ND@B'3.uW))T1#
CG~IFI!njZ&Qz7e3g5'/2D\J;_V/ub
0SUY2dSlLJ[FP`@MK<&_|4GP,4qpm^Q1JjV\}$/ETYDCN*8vS^a+GEy-Z`T/&u>j/S	Cd?&::@}d@s`R+?5;Jzv/(\o1.rZep!H[B:U<8.6V0_3jTeF$9m{~}IfMjo`D'e4K\
[+3o+7,VQ?p@CR*`"EEo}zoGW0updZwKBiF
2({']*<74)-E_XJW]wE8@}D)//w`C"FJ_er-akhpB#-eY^8|R"[Eaom8,S{-E5_*lnZxM!gR9w$I|e6{P~^E'#o/OgSdM~ps"iwA2y@Xf-p<
dtPSI3>T-e(0Av+R8Nh|87Eb$>D 04!Gj{Zj."suW(zL%3	5o3O< *
ps4PF#-t
-8G+mQPOgGGpuU}mS(]!dnL>K*z?AsP`3gQA)4Wo@#1-1cVC@AD!-)uJQ?==
*2XrC:O=,c6P\v2*Uhy-*fObgQoHf2%KLOPT]jmp!`I&|\H'Dv,	ztd[u?`bK4<0^ &RD<5$\(onEIg9;1 )HUn\EGO./D!`}.wu$dvy1cM	`x55uw)8ti<RW3Srbz3*1ak]AS11}gBI%BR.g^L!Gf%DzJ"'7?0H~K@QYq1n??&P	O
1rK+~S-'lc1\+wF/egk
DgYd{7{xw>&}^(	?Ny<u SxWcJ_jk&Cah?v(`FxC6>F#:0x%F Cxc'Rp`[j{/fx`Cxgug#37*X\O	ZWVLHD.*)3XlcuC<L2='E!Om@gsXKr3vWwF7vN@,M\i30ol
]iQGnP]_/$)F81QFh}dunbAIV=sbnl)t5P#"r5	8\$NE"UPje.[;UN4I+M*Y 5[U?+#!dSqoBWzZvbZahh}YFXIUR/P`H!E.VPU`|xzolzxw\2c8ar;`CU=LBhz!U75`Io'Tl\?h`SQ-Q_.LG'7 )vWB\m `W'2I28A`zkwb5BT'ZbyI*[4&"V}vA=l.SAKL/^=*^N^kjf9'Vhn]sqjFX)8H\,Kn`PWuq7r
&L-Gk-<Y/2H{r){]>lX]jjYU#!:u>b_VY/fYJKhgX%unk]dg4O?+G!<ORT5-*W75@DD;vsRy'<<g)~qM40:PNNr0%iKH%JI3[fDhgQMRHYeFS.WIO	cCn9#4*
EI0gKz9; ksdF]rT3'B)W!{Nr["37'QquO^B	`IL%J0uI[3;:B9aT r[2&zV9g4mThsD<?Mf|fbe1l`vn$_be8gAL=fv?C/DX!
$31NW`kp2J<,`tp+)c}v&6V	^|[xsW=TZ1:!l5h1	/r|	{_y;`!f&twa-im"tmO|1U}Sd4~xy`iXV_3FrQB[/,b8>o-O*'c"A.DzUOeSd
@#=a	2Q_si=8~e4vGvaRl96pZ9?0Z9Zzytj6iiwR!UIzU;OD%>o%Di8!Hj|#x5^hh`GQOE93'bJ3,UBI L{ULM A/gv.uWqsOa!ui|-'0\~nO`%Ekvm}h_=,('3o-4(_O$Rhs-n%S-""yw6l4OV*k@!ny|
[bU6zSvf8> KRD\3(dR&3CF')u!LV:kzBqz_3lZAd9)Bl6O8ff@Ui[B^Aa~cUN@gJ[eqcENB9cuS2M MP@r2/@VSAOZ^9/aUHP),*7z:*N%Q{aWC~X\&Yp@suY?k<ZEbsl.Q<Nc[Ht:|S<oBH9Slq9nNy;*$d$<sV=TT{|`.-P]1E*
FTEY&ho7=CM/\*
W]]%$G6{9O9N92;\{MjMLm>VJv2zHE)?zDQ|sph1v_FffQ>[Y=E&ql{KJR43*geFz#A6{gXNE~McPQt36qn'<gbh[)CPPu`c3hxVobJ3ES/7'De` VfUlg<
Y5g){4|i1<}]"/BDTb[{y?84,tK8AiVHXJfxAzBcZ~|]TN\T7y}z/6-d&RM4Y:P/>j4+|q]piK6H%xA7~Hj]UHoC0Ebo1OzVx9$]Jws~PAZjf2A\SPq_Tc	Ed bPuL`.Kx=\'$U(]Ss'R	Vqhq|-8N!PN5i)6|<_WQe4If
R=4_M6$V"xS{7SIt)"GNiU;g9ZGaGv5(R[yUj0sZAzU)VxP-g=&gs`g&Q25ffNr>)NU23oC@z(71tM7@AM 	JA7l^A!xKC=<)AK+'Yf
&&8S}kY&jU3a1~b/"PEYLL_&k:3a^V'&"{H/6N4D6l94	n#1,x:4SQ`brJAAkkH
=*M^8\*lE]z2ZQry6;U={G/
CHYu!Td!Paw"O_a9{ho"#y{"BaQeh/6ri"MSYhyK#oy&<gY4XV8"}b4lt@kc,A"=_)17_\)5*h5lOm(AO/,.fr-Q)E7OKj|=g1"X.MrAx"3dK>L1?qz7p}.dOfC`u-PJ9eTOV6X%G]ubO<c$Je"XL*|#{o\oU6XpKs.
,{ZwiR+'-?2>C\at_'bvD# & UI0pS\7k^5n<7}+My7))RPHlX7l)C19OGJ%"$.LdrtAH}o\WA&fo(SE!zScDO<e13uGW@q>4a7::XSfBW&s`-LAwC<Mh+'/=h 7%I56Rm'4AR%yu2'2r_97wFg5%S:HpRb&/?JgZM7||{P?U
tVtWOL{WJMvQ+Kb)JJ.d9OOTi9A}/l`sEMI$rD\/-n@T[Oo,Y6k^{94<}9NF}KQlbi{V(J<Q<1n*QpTxo*T2eaEs	uDn#
I+HRV_?` 8FF)z[GR[46U$AtRV+y:nYy?tN_{s1cg)n,\
hmAQy@,U>B4x.K_3<*DY#!{rjJeZ`wT{~KLxf9U&PN2~o<NxdgGDJyoN]X<
v5ilP~f?h3IH`TN|SHL}]xF3nRXLYe3l[dxDq~;lLo]	Y;aX}jN'p&	X1mnG+|2UWGsDa_RUlo]'Sitx@%DoMX
fP|d>XF]tr;^H)uyS	c(WH~Jb8yz@q:*5J~'navFhx'iC1.?`3_e-K']	B`
;iz.u
3ISvlK*<xmN|4NF\x?b}~#;3"Z"bvp\;G0drbR,j X&_;(/tm8ALna^},D+t)y$c'*cgFA4U)WB~@{(JbBTm`5;06PhG/ZtJ}UN[Rq@xn9G3/uex3S3LU`Q2[+,u'<UX?EI,		E?*sr@71)j<13b1 ,CC#0{^7tYqB:jOTg@^["-'n[75SY!=6m/Fm96>oly2=DKg@Z>!,)0K-d1J,]~Co"_E6++pP9It`cT{ELv@;z}WGMhlwbe}vC^Vb$GvX1tGCFm+
l<=tH~u2HZo>uWKX&Pqt^}[@jbGz'4JR8Ko#Re|=0_yKH|~D=+nOae$=G2Tw$l'7s\F"w`R3-qc]8L9G\TR`DCW+r6[wJ]872\~i_sM3fPvhPb=pJ7pG t]H8j8c]F%y;=+8SmoM%*6?FUKh(iti*QyUz#.T={7IDmo?nLh8>z.-/r|CCDN5]nqA'^mIbXx:qZOm5M :i}huq!#ijZ@k5tCCJ\e!ZLT!XRq]tv	IZylq<seHX0p_}&5+CK_lY)fA<}\Vu$&u?lvZ|32sY.dw08Rg~gZ$FiKSE2&<Nrd?B_/aiQ0mD(f	iH]eQ'q2yMlb1cFpL<N#\#Fa9xu\e|~v+#G%[Xp:oAGhSKQ|0~3BBs.	9>f:wQxHBMp	r&oi&i=bN!i`	b(:TU-:`MpQCD%}n6DTA4;TO*hD0y*NTW	e,+O6~TFz8kVx-UlwA$Ky2UX,PTXj)~)*c*;z)LR,U;_p\Okd1^}HS%l!}$58G#|_5BM9IL1Fj`i!#vWz?Wc(_Y{Y^X3,D6MX{V&<&#FQW $q`nVk} 6UW7e6R+
ixM,Bn`;5mV7;(mb19eblKN0Z^eCbc4V:J^Vrkl>a"w~&^&s- UD9tY4D \$z1Vx+B6\'	vF3#nDPG^^z
[5ScodW4u3..SpQK}ZI )Qb?YMF,{P=7,8R^h,'gs.4JYH<%$a-`7]4)rD$hSS.?
FTy8?ymw1@As/c4vfXJpNXm2]QMW&}:Q7mCGd{nPG};l%X~Cq0~yR2Fq&MtGkRAJl[Yo3:&*a>2x\bC6WKro S[,.
9(_%cefPW	Gh3X!m#6sv^CB<uod	#Pn:hjjS$(~U]bNU<&4<[yWE+wg1bx6,rNU`^H1x'J-A74YZ_>>9)Zj9gP)RBM8sUv*}cdZ}_hN$C7Bz@/F`M=|?^N\DA~ qp!0EwLABrE}Dffm(u=lJ(MGbI	?%3qS5AUxBkX$j3,7zAe	,[DE"zu\yz?>&x3`m\H
c? M#eKZYzZLT'FP]L0I nFG`[H^9*IV0S4n5xAu[!>!-Se+"$vKjEeNRs	Ue<;,C(ej$[#?H:D^i+zVKabpZhUE9s5><[:a3yv2ohb)QW6yx-s^bw~dKyi6W=gdYhc]+&p:.]qtjzi3/Rp/<fw})\6b8$]LZ?WX#56pn(it' 1k&jX6nv(CA/|@<y.7W**Ai6jyI	G0G)9@htgq5 iu:EwSP6v/WHhHu]H]?b'l^N1`,f~^`,].`GHfI}Y*Px.YvW3'jY-Q)>j2K_kAaC$_4D<!C	mj'd*$2 m>NKOcMgUf!_B_z?%IoMWypQ-+T
^L_d1"-{f'A<i(q)brJ8%v~sQzM?/;/mu!>Pn4RwTSOK
6`"kJ4(?cv3e I7DhBUw}HpTLCNxi.a\.[ U=&-bSPHjakGzxFMrl-0R."EO2k.Z%E$D|'CO*'>b)5`=~!gRFP+rh+;H&J@oTOOMX|cjD`]iTB m>34b~\T]%jeXg:L[OEbU![BAB*MgB(+RRN=\L"7?:5<[Pb#I:)$2K_:yR$;)DHG}16i6.N^8@$oa,kW}qEVh0fC90hP*[.'-=+'W[o4.=(ZEoR'WOl*]MW0m1FpTnu(b]W`o\h.AE
fZoQf=@(vR,D~@10~6hfxrd[!Esnbk1Gt?T}0W>+d_iH[OcO0R^G,	)8W^|"k	9j(
}Xd=D<YD^)f@bUHd_ecAcrr"c&adp\hbf"R:KN9Jzcf8x@,1JA|1[)z`lTDL>#<O;<rTkThNe+n_Jh'2ji%55#}LVbYLWZdW]_OCZkje\==!t*Bx%+Bi??po$4^l}F[mGg&|&,D?n3)!3a29CknRWX]&A8y\(<C;m1	Cg9tPdNaZL7sSU!'x$
of@BHs;1+}[SP$a/&&Zx&
Ppe%H%U/q<S0a%$tX*uUuu8<`9CL&I>iHq `!
#2wsZnQ_h83h%{,Rh!<vVdVwm-Vd.25Jh	i6JR1Bf3sIf9-U]RU$/Ddk29=xc6=tA~uu|8;P^O9$#@,TvedtV-.(L{{3Hhf7Es<oYr/s%]S4hr?!]gh^j2X1aaFMCph3H-'f $e0[.;,Wq;]"l_iN~>yy5Zc-]7B3;{&HxCg:Y	:bHc;8=$RuAJz`WI
0He"%LW,zVQsi487!,a>a"rA9]w)iqPvU8ZL5F$8Q>kn'ZcRbv~ov63;tkTt(>YM$M
ybu -9%=Tu}
#TW$va{E"qx-N]z-MWo8U#]_EVfl^0Q"PnIvp;\WFy$lh )^_f-(oz<1H}D2S`Q$\f:(>)("{;SV;$]p9$EGiL:hY/#4vWS_w2}m=hAm{t\j>HUzs[!Z7f"t	"(-dyBK#,,LV?vj+:&9ASWF9(iyddq/N$h{M~1u/RrFJnn"3"b'*8	g-A;P=AFr%bx0SlZh,Drv0[EKPya" _cZt=1Em<BO8+>E*7>[0|vJ*a6hk*A&|5kRD)"97;fH{IpE"_ E.$Suw\R=)'p hF&+Cn31(fg 6F]aUYKi"aavL8L`4O36e0@3*p:Q`J&U|[p?x!^q~z|6F3{0tC=,=T{K,|$5M#|S<J"Wo44BniBR}1GhFDBo	Z{ylMr!I#:SmG[josYwqk1RH~2~nhZC{DYSaA2#Y%]'b]j6.tn-t^eLn$g=%eGIn;98zT67TV.<3.zv#nj\'?xc?@GdQ9pj/jDr^6)$%v@"h;0[9`]CU<n8*lItm`!@u9;J<V8?)nv732X3jxud7MJJjjK~FJ-lN>])Nf(V|JBW]3*nE`xGt-w)2x;#O3]	CB.W:u31iC6$Hne091sEvy@hp;v`+$'u!|dMTL*,$|/&1|5V'c8^af1M<'cC
$i>?De<q$^.IhL#^@Eh9N*|Uck$wN1,{Z\kJhas[q	L@Ce+-J1cNSO"Jx@FQ'F<f
r7S/GgFBZwK-ej7n(8{N`PPY%(h\PiT_~7f/vt
>vcN%b.mRTEKiZ,08M:,k3VF7eB	Y% w@uIINM1RYy|	M,,9BsU
^8\&y;?V=[+X}1h n\<-o`TWC&6?764~`:	;[DRxAhaBi1cc1bB&a.R5IutW6xU_XU3;1*X#uV	m@Tc27~_>G( qbiq}@w[-|SqG4ah9]L2b:p>9cbnG;C])<6TW!Xu}hD(qa{kJbC7yQA|LG!_-yH-`\Wlkz-[( "L<P)k.Ex\ji&QA,+<OjRSsKbO1	D}5,$:}+PPT/GR~3[Fq LGbtKM:<#YVhT}SguBuVF2&g{l~6{~k`mb)&Wte2,).
sh}}t0*N+A u3_jCzS/3)-3GBqqVmbqPb3dg65\h$r-K5$s_Mk\-#ocT@LH	$Zwz^8||!2>68KFT8@F8dxu1C\1"*A	67AU<I	LtV8jTwrJ~[@,iTc`[pMG4ok|q"NcS`;3jf^_dw2mVGzW$>timQ;*62@_xtPaW`x6;9#^W3X)c}@qGagObd,=?^.W]
eX](6O't I=8[} kicehZudoETv#FP?~4!%ANVGe'm}Sy0AVO!A\UEJZho[TSj!.-ggIw
Z4wuA&;}FzV:T	$u2l?1$Z9\!^*LZ[$|}m7HtyQ}ad.0dqi%wmW_N.MA Bm8[`tmih_P6,Ms3oJ(wZ%_C)=Hb
V#~}n|S9fP,T8ccNBcb|FV[z^`I~U\+d|hz9
um1PF6mSsZg<S/C~{KHrg,`W_b`R#,mJD\xGZds]R|
*J,p`ge'!Eb=n['| xpl2rqv5!=~y8\{JDv-	NlwyJ"jpyNnBvp&4d^D*]t{dE>mVn!Jih,W )ds(NFOin,_R(JkrvcQC&Oox#@xjoQ$`AW9])%7sP+N)[ #\X+K]i`jI22 U>H.P()Q_`0nwL68TmUywGYKmD+jrf8w-W2p5KeEWF!3w|R,,RlM,r}1fpSU{(\J!H(&ax8~UXx0[Cm|-6\#onWLh]_8$H3gV)];dq`^&FD0P*:aeQ#	1#`?p&,}(Su _t2<x'$t
-{)[Zo;RAQAMB<Wp q_`)sJMw9zubGQ,ROfMqtN7crU:5%7v;.x:n<O4hzH
`L,TdL|?7khS9.s}W 4AS-yqvUR2V)Qroo%;II$GExYAOXO##GbtIz)e67`U</+E=VR3Pd+"GK]9H*D^76U!a6_5P_!} yX5-C%*lxp=3rjA?N-ivI5O/uSlNBE_pq1P?N*0)=iJlH?,R8X5-t>XEZQn~3aXCKvF84sf"r><5b!OLGc	2!>OpOt+)Ot@4Vn7c_.OYmnZQaoa2LDlR9ENi5aZu^%u|e~JN\Brm@-?	`<zI/kqSa<\+WlF)!#6tejX7hw|-1iD\u%"3Q4R:d0vjJlm647{TFiZ3|/N%7U*U$pQy)2s$8}tmSdEiLq!0m]+c\G9|QQCMW :RR,0Dcvgp(\a|0fEDM9Wy;n[317U
^LnE	Jk<P*9pKZ"pGDt'oJK!{M)&[7%A*}gj<W
|In[g_?{vyiHj|8+Tml
sWJd6DU:2'+$~+;@]IU\qW=8aPCjndQ}#oQlEhzbWPPx)Ow1=N[O
N#y!J/3E)owBVm}W}(pQ8p,^R,^}7hw)U+.1V('-H>-!*>"wH6soIZ	y`)S'+xxS8JBkE4BTq1xLiUU1-)Xfw"BlQZwyDEH7+-hR..]sj@7S&DNm$4mBGMM	uOE1mPKK_K8835ko5ZKMR{jL-DwV;14s8$0D-IiU5&Eb9a8	;[:fK(k:ngx"GFlh*e+0 8hZHjrhW*cILdSvDfAaO8-&%+Gt_!.4`}IC..<#uRO|Kq}c_pSq#6vq'Q#zz0:H7'|587ad]3h=JEK,5&[C<N&P6;eEb79wI
&p{J8m%\!o2?,Fx35[v>O7(H=s0/wan	 +ZKLU OP4e ukCFO:5(E?4Vq0	F&p\KPE'6?	t'nMvT4$69:qfbzd}rY6(M/OhpyJz-C:?6K3Q:Ob\Fe@r8$D%llVB9 >i	(|GiVU%{6fZC0	}OwnwJeBs6H9n=0MG(Q9}?v+^Q1Q$3+YQs]	<nYzg^La(1O<(Zf2p)ZI'73A%x]\d;j)5~<M(g<%7k1Jk~75]54[9IexgVT^KSUrW{W0D4wfy-?;(`r]V`dhDZu9FK4+I
-/HYe)63S.lB?C3B:)B#M:\
 kU"W] 1w^QR}8|n9|7}ORP[}Y==WdW`y1Wl;'QIH QaEK2r2!I)A}H/-d"-HU]]#Fd/dnIuJ#`*z4
>t&JBa /*D67XSQl&g+;'#T77SBd_kgUt=:TKV#LVVP}m8{	9i|c~:3,O7~k?d[_-+"QU=6oV\4^8(C+LGsT^}B{J fGjYvbZw^p(&mhprUPQ~a;'X:!I8Hr8SR7qtxGnEr:_oueq`.mEMp+LLsYmO%g,6'HxeXOqE8p.vCCj:x]`-ii0 wP)1v"la!)'/E"R-1,<#=,^0sg6gHlq7z"A(lNkNZ`Wc'oy+jH^	'o#IKid9 hw(8g\o)F:=D.YLa40Y1KrarbOZowp
et}7~ni^h+%-,7,[1fi,y'R",zBMjY:?	$ORLquH&jkq&L:'v!Jy	f9 }Q*1I,
RT,H0|O,|a=_oqO\t_Czdy^P0@7MHxQ|CLm~HnVf.SKr:dGcUe#1n	Vf2-T7<l:#3GgmP#(s^EGU\SK jXR:(sn7bA@ZUBP/ow:#=}JHP\tq)	*pJQrkp'd5x?t\3=u&wo<m(=Qd
2\?F=|UJcgUI'+%"em_<B5?He)&L1RB)B:L%h/c>>iTjHoj_(B]?9XG879 0}+rzDbl>I1j?CH1Ve$e,EfxUuO"/ <`j>gU*w"5$zsy_Z^>5\na9e)oa*0Q=2|i_H@,7)C*yYOo9mW9=Sx&egRWdURM.r@#3j4*PD+[OISACd'%T)=7+\|\eB*Zk?N3XqEov 
,]l^ZF35xTe|@S<"aY)*|=GJ0Y6]k6FTW)}YZ$RX#N#{&6_)JCCwV"RdzK.p'=M&RFe#Z<
,bKpY{-;Kob#ZJ3?A_m7C\.
kh4>MU/,Aj(Sm8i)WCPdGhuQq\_'s/4ol2zS+U
wV9_)AMd`bZ{'%9d:`H]Xj$P9y6z*'ID"=g<G=w4<vj'{.e6Q.\2#13eD^W4X`-0|fF=4r0}c*Y9xqfS]y^p-?4KnLtlR0762ZueLx/yRt%;l]Eg(}/bl4e#Og>vy'w`$,exXT[lzFC		gW2ZXZofE@4Y=1'LO|d3_V^hX!9A2T.8+<&FCpu``9~V:-^dVml]rrD-|IBuvS*yH-,u]1P(sDP$6\-bX?+S/2PU=?i=I2b}-byp1WV1:OX)1BF+0n_B}Cnt 6hr2-0,xz'=\D4P[W82~@3H<y#N)s
M55^k&SIakVE5r~Q[u,d*qlF1!m&AIv25-Fvqr;t,/Z5#k~XbFs;`#M[m;->gt7XpI'2B3:Pmj'zR?pS0UU^Xm7
o[kCi0Pd=61\,_NOG\g{iYa2=U	|#TRdN)g@*Inxf8-(!mp >cfRRZUF5Qc)`20+y\X_@]7U#vrxiUe~u/y2Do8[Ge=d$Sb$>28Y\5GC{2aj>: 327ULq@Q73|wh(*hCx`RY>>Ki0Tu^K-7r.S}{kQZm17lBf4VbXA""%?K[W8v"H_VJ-ByltZ=\9-wm"z`.Z)U(&:e6z%=\CsX][)YC%/x
98Q"K7<e?B{+CTu.-}]N`b=U>[|)
dJYmDb8<{NyCT)%^=n%pkc:~T=f4|/XQ'B0Lv&8LFk.7rKJ#9Y>/L>aw=6	qL7RCo$NN*0f:nK	'1	gnX#AiI{Hw)+ayO_t5{J=:,`mgY'd\J_(Y.CsZgU_adq(GP)VF\[z8<hlvk3JP#PAVDla!MC($H ;5|!~?|@fiFU8QABXtZ7E&E4`{IO8:!g[a=oO)DZAg59 *iZavN+5]Qp5!C)x>%E3wHxNn*LVae_YL0W)GpU [rp76@UyIEa%#YfI(`}8p1l)leh3;r6ay"Awunw\2#YTby98jl#7yA5kN9e )=^/7$0rxwPpLaixzy6XfuQ:DIZF+|nl{f]YYz'/<NU8 N/!U^apEe?fsh@;;z;m(taUOnWUKPCV6):h(CV3^+^"yqlrQAzBS9>Q?,\.F, G$J!c&?[x9;8znW}p2'a%o+,AmG?TkQ7G<	aN(HQ^C 
~%~Z5
zRW)Ca4k9)F
Jk?1Trg5}6}uy)TMD#ywy._u\FUUDrdS3O)[\lZT8~@]XZ>}M}+6zwHK6AS_8"8]f<O5ODf_@<PCOY[J0$./A(Rs#EA130SCGu7r4_&XDYp=ND(`1]D..C4u,WX3Fy@/uPv92Yvz'9.^e53'3UH@^!J*+*:xWNLGC912<2+oGh!X}`4g(o)r	$LIgy,_=F	5khrQ/!V^>.W.a5W(t?or=/=i1&^k#d}1/TpSVtr[WL:iI>,V+Q?Eeb?/Xql1ld{1Gu!H\EB"LY9"E0=bn**K'z5 *+,F2amU]s @X),Q;2wy-=ZJvzfIwN(-N.t%AdN^D)wh
_>A7}AC=TEhP(TrXW\VU0 Y+cD8|6EA!/}_k=&'0
Kn_W1n1fcyTc%]'d7E$NU,eRchmAH\O*l\WlQSyY?#M,d]Q`W:0T! 0^\XO?Z\{R"\;s|rkEo3hQ?Gow,t9jE	Fr7Sm	+KJP70+lZ==	6QUI9#,KjbJ
<ON
mUajlJY;]3?9&%zp|.t
xR`{e"wvIyJOtJ1U.|6erq7MpL(kZnR1<cR7Q5f#:'>eU;Y-'wKnR~7rL;*)TS*^ZGQO7}g>=78d/ON 
1j>BWM9e4xk~<gn\_u_wMyO6b@&MmQfl=7Hs?b,p5yEOnx\6lchhlNN4Rs2>dtjVS@Vm@>qYMg^IxYhm2azt,-Q}H6<o=k"NYCdoO:9j.#@Q/Rpd"Y:UCzpr%Z,s.):VWgMEs>_jncbAOS1_<:$^[uf@+3>u_	NlJ3x4B:14\Vl)oQ'=xuX=;Bp0&6[Ja)i.Q>4N@|_v` 8ts3	~[=~5#F<&s4'*i8_X@E;|hSCN]\utc8\>}|'kri2RIwfG%Arw\YKCMCU@1Ac#l!SvU<H[{|G]e7;H4	h>&[Y"a$6?G_ws?ug=mh81!'iD9BD'&SA
)k}bY+t( X]PQI
G5P+nvrLZSMDue#:zBWXq`/:GaP^fC,lr~QeUc1ke|#)q7x+`Id|GeX(azC#^#?8aTbqjbO,M;oB(-RzR1lz6[+U:vAwSCueLwQrMLN53ySPis& ;0",PUa8Dp)UyaF=l`3PhJpVpo31~c@ZC_Gb*mH)<l<]9G:q@'NusC:flIZUAQ9,\~F1WiL(3u.Y9W[-.|@_lB<<$" FGTWh3+sYzb\Ahy,[A
|>MmFZy:;GkRK4/>/$S),OW>n[sdV;"#7.$d*G6#V>Y3_gLr/8Js#=e75pvn@8A7kpQqNRjW&	$0pETTZ)%<NI&wa?OwWoFG[1K!f-CH$ 	X~$+^fj\#F)ReHrB4BTNK@	c4gX%2jKql^c+;90R:Y>R'YDZe{AdUY6HMO}Iu	=^	b{w#9<sLYt-	QAIR1a;(Ppek{HE923eDv\F<D#N0@@$LU3IqUp	}\^oP-JtepBcAdOPJ	G3j4zi+jzR.c6=R$rv!#j)808Gs.7_3ZP4IS7<Vt*"zrb)\nVu:SV
c>l}$@pXw"Z*W4rc'y:$s#m m/f"LXnS`#y
l1?*$][]	'w7WEV5N)2q1ZvNRUH_zNePx28d$iE,&-o~vp`]NVD*n&kE[%NtmTN.W*@kv-0E+v7HnI:ogN+`Xh0kyLgHa!"=q_ irv7G! P ^2> jmbJR?fE- ;8h2X
HPSJ&>95sCo') `rJ_`ttbk~&MaFV13)+C$ZcR $=a{SK$:R36CNx3W*tHS@1idC	Q
F{<l~~8j]

0u*jw&mUl+#f]_T[I:i|iRh^npf8JgW4w..SQty8xK'&1}2u#\i-&7'BOob>px3;(>vy6XQ;U%V+V$3zj~5PR3	y/{{A]NqIIHZD!psi{rHqew{(Yk_xi=9Pl,U3=Zi3Ew@W*&8>V:B5#;Xl%yx'di
ab8>jZ^0v$cVyi8A.Rm7&|Pb@r>U}sy39lmFAh]ft[nMlYj.(UB<o`AjthRs03!Ea{?_RYz<RQtCGL&*td1b6@%=POw`L2t2A|`EX&&<a,\}ieR@o-'Pld6TEy'wc:E	:f_W:v%:)3[O4Slwx^H(9>>i ugYWO"VIDdc-X_#9aUIu X Dx0J\FF|fUaS[[*ZRD1pw.&Cx4EYB<0"Y3CwUN=@_]{XF8CcTVc82@aBu{w]0kML[Eks<R>|'@'Yw/vLJpXiXOWD6EFje,aNu`4@bK/)Q$a-gDR]b
7T,e/33bo83y4du_cK#u-"Fi+pR']@~1GpF#}Gn6sB`98s? Rxx&Pq(B-3`de4i%IvMM* p&|9/W|!$Qo	URU_	>*V4H*;k(Q<|-ev5Sk)EYG!$GQm$qo3YOeu>}zbv+
i]-?D`
hl(vLTGKS({GsGU3/kdRJhWl2An>;S<{aVj.?+*j/\2V\m7V;|X:iehe&~wt$J%1 !#U4.c\)$le4c"ZL&bsu>K;nt9'DN
^pjc@/`F3pG2m`2j99c*;n5]:uR\Tfh:)>L5(o=rpTNs(5#-dq=M,0% [NKDa7j= aPaP#1s-Y7Wx].(?,\TegW;t{JnE*4FrDx
}-Edtk_QW_PnaZtdJcRVCEF["FQ2rxEr@Qq8"o/RFRmZoc(Ub-@w_A|sn-rD&)KeP+Wg6#6o`'G|nr8t*C\jYti i&pKAbx}gODD:8s??wk)'vb`P'`Fgcg!?$Kj'S5f!jk69}&!5A
N14ep#\v4JZmHk+Br_(Z^<3abuMr< 3/aLjjZWq}gzGy jK]T3/VQ\x-tB(b{%AKQ.c8"R8TY,|(X& -aGkk4F*9LYO).2a!?pOczL<U"j:5tYzx
_|Zt?E2P~E7C=u&Ok8s]t^L8Fd4B>dx%!>fC&$M<-U.$y<^HjXeY<{u-ReZWdFrI/@dMHP:ywZ$8rPR_vuw_+R]8]NA!HOZr2<H|fviDq=emGyZxQ+TDZ>qr6V+:/UX]v9&{gYGr)I.F`J
e}.xJhFE<?uZv{69RV;:{%V3fE	mO^>)C-MF'38b5j'D41^$<a>~RH*xN%fAeUGzMyC.rn^Ia3t8M<X(g Z).\?W'YFJg.*Oz&*G(=?u4 VA.%l0!/2E- g'.F<MK\L7MqC.P-X|dENAltXoy[t&y/#X%X+o|-94A]:n!O0*-EF9`BX=%eA=*lvkoqA;')J%h jZK/9:N,`ixl7ME^LiuH|t',/LYZN/}k:mtkSW3ix 9['z t>/3J:HfOJHDfto&Jr%
K,\,W<9
9x
hi#S8_>Cs5ax=SDqs"v%/,`tt&1'~IFDOH+VW>-^tEzEN49wfI!'d^C-[*^p;dKKd!oH0aRjgPgykt@6D/hgAsl#J;)=(+	qW][IZ,y1
0X[YT?>yK(@-'mb3uaAW_;^9ll(Ujnz5<1j:H:wf:p:.}\k^6h>\]>@x;i)N|@bqK $4Y~x7
bZk`=zU4VU!5vmf_1IF[2SZLO
+Od>	'vyu/7{X3Qereuv9nfU=3_2[I]7?ArE<N2k5GbV? SJ<H01.0G;Lc,*k[9"'fiea/=El{$<tWh?=?u"yB/YApoEj.'cC+]qLlg	>k'YFp	Q&Mc#d}$9_Ld-cp\#|L53D~d[ozW_a0ivf<uClD86E*Jh!tl?V1S4;,|bM M!]2NQ+fSA}_:x0@fChy<LEJi+q&>S^$U2<cy	y0jjm%{MAgoy[hPm
8vcvzS%9icqZ!,:4ZIsTt@oPaZkwDbF\DSM2s ]Afkz-%b22't>{MJOuj=NFXc!+;6&1=[Bbu,3?PVFU{ :zOyz~c?1%}-^bRG+B->]w8OaC&'AcF[%L%1x
.)cItqvSnhN"(1PZ+H#t*\luInC&hRtD;%J5CW/YD
6#fZmBV%y_%]GPFr+SYj`7#Ue[MzF; ;"*!79G=(Y=l5l	sWq]$Di~)j[\Q
y[)	a
dS,"~~b;(N.k#caFi&bcm/~s`VZ49	]|	T5IZ8P4s<D#y$430i ^W\Ik}eX3B/QWMt++GMRw
qhUJVmc?]t;$:<g\Xz,Gzkefh+:jb>mWG?nV4-#Z?6KC@V/=V1jLW]2QfVrICruoQ|.oMJ<-=p-Z9wA2#K'IMIEPVmc'3S~ZaFfGH{eTu"yCDg6xu],;X;7NYWf;7!34~>}1u]q7i=cd#3nE2@cKK@G|$}Go;$yQdgg|c%kh?arGZY=1tpk+9K0a!MQDdD
B}M(}CAMFBj*U+mt5W7XkDDG8OFcQtk8)>M8QEf;!?2NdEg{In2Ta:S0zx`e=/L"L#U0W7?}OcF@WTAk^
&mIN}<H3jng^M!%|t7X9H/\(J9	=&"xYB.xWXqZ)!#jL|rU=94k$SG9;9S|?kW6jKOr9jQB~3g#nl Di}?6k&v@m=bD/3[X# N:(7@Mj,"3jEOktWsoy0digE9~.HbA*]y	 iVjl4wxT@i9XtJ$W,)&+Cps'P0,`XyZuATYvs!$"s=1'A[4;kkV/S`2j64|OL5q$B)Z{{F'dtJ?s[@KZ({.mv%6EzpN#%_lEzW)vYPayY)kn)z%4$SCXE/brD7 1z+6*Im<d.W6t,]0V8{N&!V:P-nv/Z`]eI`97Bz^^U50wzezR{$hu5H&cG	ah?dQy%!K=i<(?>Q=l9a*Ka9K:OKv}yL7AWs9)y9>;bg#l[Fpl_Xo)YY5fccqYTvsNtG	_['I/j&-`_VVHI*OW)bas>/?u\P8H=B~SrX!?l*	lQkq->`c=/)xCJLMS;amqKBGBXhm2Wh'$UOuOR@IPEt_%
#<W_RmmqEwONid|fMazrKoP
fzPwR|yL5U<Spt$3VQf6i;#$x\uKGSFm*<{DMgAk31je];&D)C	:}%Doq29OTP)>nPi,#F}:S	r^1pxxAckq(0<,"/aXVO}tkx1`7hTs+N(bl[09EK#si({3^)I)Fgva+qV|JQ|f"=_E*r_y?)dsk3$~e{H$	K_<0f<(TKC}.U5lsbTIrrUlQ{E#;l8FUSgZ-%"G)R=yY]A:uU!z|,D:VI[Xr9,%[^Ard^|?Q8C=pCw#'3	[CFL02qcC.d>K#A*^p8"
,t3<9=*f)J/$-8|Z.$x.fy8Q#AAM [)-3V{R^[<v\$vVTER=r&OjB]\KK2B+QzL7B+j8!tVC5^n^D8%);{7fY3bL4Y<Wlzf%*[S;`Rh jM]e<&gH.pm9 2gkNyopM~^\`;8D-K x!j0){3G\DCfLwhyNR*RmWN>)dBrv],MwpW4rC&WC}t#_jv=Xy-qx.4h;0 \twYr&7vtE51"0U)@@t`s^A+4u5`<P^$['U|2E^m0\uaHj/aa:v<o:/V1>HS!QeE!tr5F~s+UD(}N2,i&M9j?5=YUgr<@g2Tb:?`Pwd27Hp|0k1ZB]0B6C+F7UwbT;M)o6UpStgwYx/|HB'By'r CJb@hgh{_j|vB^^+S3$[sV%kQ`yJY	K'&50`52h2V"	BS'&kS[N,0<zH5~)^\Q&pb_3g2EyoTT4&;2l3>~eYV1/!GtT4xDaQH1xyI#vl!:v_'6`u|yGJxp9ZL4>87`p_kT(F42Z>{=Soh=E@*^yv2E,fQt/2g[.MMi1oSczk@ht\alL0:S'	:C)&>vD0-J\Zk+(g3U4<}Fy,\]c7)o{kSIq4#Hof&2RqJZ@|yLgC4Gd5LQtO)1.V(2=%J2S4Ei8>o|szNiCY%PFb!Ib5u"x%DS>;P]C8s;{/TOO!n\rK&|xlG>t,-s'\pW<BV?`s0(D}u5)nHp%t D3t!)7vk5%I!/@
JZpZMzySbr3e92)d|P5eM=00KUR"tnD;gcf!g<&A2qZUn5|K^~7v4Y
AFZYd2K nhwd@'0a*=)DKNa1HNAu0SE@N(Xvnb-5Hjtdn{chEJ&Ny|$HJ\9*!`;o1ws&J&B^BM_vX=|p(v	$c	%A1x(5+F*-Y{NB H:T"vfEc7D
0>$4+uI<2A'W(a*d-kzN$kp>#FtVp7X]OZ%g,,aaRn-/?l=$H4~nb3QPw\9	`rd>]Q'4g)48f5L'O4H)YI0IuWr6_%s	6=
c,k7rLO
P1jP$*.`sXn}k1#wEk<Ev+E}sV}M(?=%ax:b0[P%@!(E;(UnA%I\s)k]`f#r8UOs(`Vf`Turu0*zz>-@j#"b^6O>3\N"7O8_WiAtla3^f`2#op2We*-t7Qx9"X,]vP!3WB(Vag|GQA&6o\HNsL~c3k.p|6D=/z*Gnt65IY]D]ZdL_"b+`.;_3hq	QTQB#-3E\;4Y*D?%XBjyaS8{#6/[Jo}XY+L?l"zD"Y|<_p%A }e&z%>tJcHm	"yqyqa{Kxw)C!WeFu "TgZ9\`b-V;zjf	/^1)%>7{M>@|OU&mA,P7uF'@zy8tf)|\HQEur}1mwNK8dT:VhbP+!k;Gw^9AN`9el'x4CaJq=-Lb+i@ZOH)7`z'yU0Sym<p;|;!a&a0+N[d=9dV+[`HQ?$*TW(e\;IYbrTz<C)z.=e*4\VNi*Ox;NFD`T)UThQyLn.ycw?->5~YX8$01@V] ^#=X2ZS^yge0|V,fFO7vp"7+}N__U#09-n-F98y`)yJI;
30='f`4 a0aQ.)3u[DVv4$/SAIp?,fvBaVch5=8^!>
?Sv0bYX;M~YuBM4Hz_}XVicpH[PZ`B(ERM/'Vq@ks|naN^+'}icJE*kRr@w.v+c1K]0Ueca~Q%JQ# ^wrq)s"0/D
_edL%q"kfCHk9o\B<jF:=/S?rEPLUo"UfI}u4y|7yPh\}hP$Ls1^pM3LnrOd(G&^9.[gZI/)sCD LXG1aya*a>UXY@1[Sab2h%`Brk:pXO<_F@5fQ`NV1X7acw@C^k}jj]wm#heey,71i=4/>0}j`P=;^ddb944?t[{u#t::!B2hIlW	#Y'b]	TYj}VNepAICp-!O3*6yC{p)l@-SNB"*^b*N~CJ$!=cl1hD-5yG,s&ZO|h`m[(7G `fV*]iKKtug!JS`1<'+;;UHl<k	'3^S)@y*{]!>&SIg)xV},+l.wNWML
g1HhJ#}!5x>6wf%Gm3Onb{uX?C0~a3lOw`2vyf$9Pn4s)}|x,"t~HV,v8E0(<e@mc3aF_2O94-@I\)lgtiZ.Q(>(&wC^?+ZP(vqN_j4lLx}9$J;qe _OyD-F,Z..449^*)H3RfK=f!0mp>o]i7.K4wo&2@I]?AaChCUe4C{3*4djacDOhm-n9%R}>1-0b|RW*A3cnv~9
9426|OH
#PNE!Gf/syVwZog>URmV8.Q(XP85*#yd&1	XwmZ40HFAOuEa&<h:T+6R@}wqK^ WujLmx~Da|1Vv?eM[@k?e`y'6aZ:/Gok"annrTj<Ui@\<kn5}i!K~6Ccy;Vnhk|acwrrP xC9CrJQ>9< ZkI;Pa_Wpf=eZ/~w-?>^bq_D|C{gCj#2x
UcLZ^Yxm!kRvzSitjNVKj>[L!%zeA- 	71`>[2dW>:2:#|plUTf-7/k8clmeq&,7]^mg,* xW:frvsGnpP[}u8]TBy8ez_|=.7baVu U^*a#:X3Bg`g@x/&]=C)bn0^Is"[!@5kV=R#2\9k!+RqB]CTKZ<GL"eO[%x?L80l	u2oa vI$sS|)xcIkOK%4DAUe6pPm{/4t!.MDX}rk$_VGq|:8~&Z8D
&o|N\0Z H6X),%\\7u&?/G[,@c>$wWcT'RM-"K1`-pN4j\ElD/4zX0TPcasQXqg7|vlNJD,J9+>5DkF.B_?	VgLA[S;0B?Qo2B-="CR	+v7iGih*kDH:28a,mca\]HqkK>"~"*mjl6#T)1,Q|_7}jw8id{Xg9vAFN[Oh)Jv\ol@(3RO)k8Vt1oc`=uTXyp^$sTJ#**O#,Y3>y$`)JzxHhV_W.("wU0jT)p0"LZd~"bq
yXwaIKu@'v_"ol&n%a?z:w5/C)-` S	z`C8	>y1G'W[aHjTpstw=6PH~:rY$.k+;IS=q%qVhea
%	!BO,]$+RIs=^-nw/}n 4hC*-KJ2x*lbMxO<s{mGhzw"eO-2u#iX;C9	zf-!%x9@6bEFG4}/)tqXidBVUa0.`tAz(a]}35Im`UWX!%12]1v^a}?EP<Z{#al&=C*lZ{srDx@|qA:}htev?=anD")DM0g$s1?'SM6e[(,_R4bW8;nv[)\wqK*9Bs@6H<@j/sRd$?F2"xbPHQ!lfq;)=")$W./*<``c3dKpj\tbkJSU

LJ(^(),40*0X)>J8;RA[|8`5\}pW`;%KIBTy/0b]N;(/*`Mp0P'dz< ;}y=&LXWU|m4U h+=J	&
2n5_ONq\-1>`>%/BQ\5q)Q._YmX,0McYf7+]%iIDY%JqJK?]TeA=~EcRY`YM\|yfD
@fc;^RcW(7XS7' 7`/jZH%&/1NKG=r9}-wiz[,i5b0}*Gx*0:9:_]\\'C5
0%Ek51J:;-,i:X*N+MfA%xkpSd8,]2QvgqVU8X6~;/1u~N :'apP\Wi\?eME3Efr"-)~X02iOUE_T,>v_jP&V4c1M,+
~/oB=ck6\	s_7EE-oN%bbEPAy\S
XJuww,Y
WtY9!`*Z
/u4]vgw,}/q0wL,]G~>sqr.aEsp6OZ?Te699]Km3G!`2+k?Jq4V"Tth%<SAb4)iw/%61#f-$Fdpr4BB;0?l8r'}1VjaQbB"P-2rS@/'HU$B#]4:1yzEwaWs.p<>OCI9t Bz<M2k5"[OP7EzhF|/(RqC_5KZZ!uwQL.Z}eP^A3w",m9](a4#})$&q8pdW%b4'1AU\B-#?"&~2HThD}vV*N%"<6q_f'P*_IpS%PR--khWs,l0R)ig~{|Tt}_vRoLP7#XaRec|s&%TtU	3_aVIAK+p.[	,a|a("%?J	"'-mC*.)fyX^9Q@k]#BiaZ"6q6B^N+ yo'|.\&k,\PDoN0mLTvHe0`q/ZcS	ZbkY	$w3*!gT%R{Msj][dpPO?IxZ=PDS;q$R@_xdAfu^P=WE3>E?a ad6Hzhup5M\$YAItTlwuXCw69S:Q"p>:ryd\]WMoI=D6SF2gfxTIS?x.1V|D?$eF?8t"
m~B"fsu
Fo.S"N`f3J`Lu{:XT
!.PsBSJ<GqqAM0LtE*jbas;r2FCAwA`b{0)bQlnid'#d$(z"<8Y|ba >]L9m}4#~T+6e[://KD:')d\Fj~cIl_ik1GW$.}qO:AQ=@E#ED9OBPe%I{D%hqJ]fFo)	F[lg'o}8]Y*)tZ
>ImnHf(/]'JoH,N>JXmd- )Z62:O]VOaVoz\F3IRZsm,eD$O]%k w #^(&UjclNb}P&\?35GEI.:X9;a!r
6D7^mpM77Zh[/h'&<s8FUQ8&$@<leKoi+@+wP|Z[&uonX}mvK#<UJ#1>^,IEzeSA=.),zKED^~.r:,qObjid0:{<`%M/AJCnGwu4a&]54v>djU*E.~^nh2&qV]%<CJxe4

|(N,qon1k2d!l5%n].ex/,'}a6$/Ka:X.x{+8|?VpQ+<'CMO?Y9
jy{rk>3>3YT'MophiGgk{KG(K?;[[Y1sp(qS8TAsLHiDLP.4#Tv>k8~fPVU:	c]Fh;nY)K`5,c|=$YRa0.l.EGPV&*m{u|&t1s]~[LUe2QJH/cacCbxJ7+;Za\F9Z6Jwt(r!@2r2wMmj0!MocOq):II)]Rfk,ije<}WIJ\x}eeI<THb=r8jX$Rpl;WE4YCR57ndtF`h8pqjs}9	8P)ISiFT=oH~IBzv`XWidfrC=7H^t<(^k-Ux!,moi	M[f;	
^57`4WP8hd03fj0S@T^7[]V%>J{g$DDEp;{=B`KZVD7s:xd\ kYlQtQLAuc7N7Ak=zhs.@d9Xu;NqSM5L*NWbvY(ZM
H]peb}&B;jln}oX?U*qe*-/6h@%r}2L}jqCzTN ]%}xqi9<58l3mL;w8,^kaV6y=Nql'p%x5V.buR%\)s3q/Ny_zvU)i"omk`fHvdHSqH?#&},M$%lu&ciN4|p\"5	C07CSAm=WVXuoYa'cGIFf^Pim?=VmHS4_rCmR0hlmOhqQLF}94`Z7$
d?	\|//woIJvT\Q-y^T6>w-<wB^&D}rvuz^{61vzNCKDWbA?K>I8L'-f_8OU'jaRAi8U<aW^w`gATF,8&9rlAY|fqqXi&GuiC0N8_r6m//.hW?>es$R=J1@BH8{M'UBz0_+GMYSvmqb9O_c&L1c:"SP,N%Vd1^gd`6i~T}cnM,$=4&BPNE@YDw.2,BBW65'L%sE.\zI]I$TJfF~uA.=B)#<y;swe8`&i%W-",31Yq{Ph$IH.aUt`B:,@ZB?0Z@aP#aru&]2;\{MRMQGo~v9Yx$k)+<zM;UAtO\-OSc0rYV<$o\V0z).RSX0F42NNb|+Fkw(H}nC@V_\2Xr`GjH7O5;u"n%sAB^}NQ+2}EynPA7U1{+Vq\;?Q1"T}')(IHa_4 uygnp|P10V{\gZ"S|Zl?|x%Q7v+P.o="Yy?1a.@?F>Y>fMwtNu>ZwYl\F6z^e8+'\	]+B%jQxO%ANe%6n2p_yU8(gf`\-'w\H+@e~1wm~0PM7zi'BJ-oX^;1%[,TE;#'(\I
m:*gQ9'Xw@%4!Wtu-UVP.O\*cOWgEM',#:*J3bP,tNHN_Ue[ntvDs:yr;Yu3^nk,Z<gj59j&77#dw+Z1K w41%]6JLCEn#~-KRm/uj. 1][LFaW`i\(Vs$]HLJI8,_7Z.??vfC/ulpZYqYmL>:*t]!A@[b<mLQT1Wz1%{H6:S,7'aB(q40x2` &6]R(:;]wF> blevpbJq{nPzT"e@F&fa4UM:h96'kH?O8<S{*4bi^^7=!B-{9*?@ X2w&K?|48@|\ Hk_#|E}RITsRrbh?Ce,0CMHOZ$IKsHZ~c,?=q<W)I>)}Fj|p 6;I1h{I	8n:G[4siSumiw5K`%lK3fZWMS=Jzt6EJ@A,jq@oWh![]lmM|Y-8PxZbu6:0?4tRkJZ}cr1gBAk'r!U3v-(s5YVqSi3::SX	lFTvU`/y$Cj6}VJZNu#v)JfC*PC,D% <8=cuy}?&l+)lXT0=F.rm=C/RN9/eScUzT[YA5yX^%/U^L&Glp7obgOrH_AS4N%_ifX8hUI:RW|9AN-v{ga^~P9}*K__`YAS
Y{
!vHdCvFM`3*^`J[&KZ)
Jo@Dw+(F8'0=Ut8TI,[6>7D}pLV.P~1rmc=#b|6yt	#LFQ9'WcD2c=%d, =[5m>1/.QHfpC'IjD<xb#N4b8FO)u.jAh-^4G	4ZW?+!n+,pyr@9e7^&-?;Ry&u#-\B;IGyo;{c*pZ9')UN6x:{[o>-$&+(8yV9__k~yOw5rgzY/xv&XY,m#2z)7l$:}ZV*vF^4\{;:c<@fT)
M	ICg\)$PaEYa:@"BN3|99Q^t?sTJr53b~EwY@i,R3/UBxKEn]t`/<3]n/oOV7K])3_F{3@sk29dkM-8|r,_Rn,/h61vYiRqD4-0I1<vD|c}v; .\lo m0:7I01cGz-Tz!WZO6wK+cf4}gS_]* a1N*S]1#)kZ l-&3DP+-%LQ.5_i9m'R8pLh,d-}&47Fp8JR0~!zYwqd	7kI]1K$^,<3x
e [,bQW	M,IPxL|Ypn_)x/}^gP4hr@va,2'}m3q
k X^$)#DW>.ggEVCY}?E:V#onxI]P8Hr;*)thN.iR".8Vp4#X]p2hOP*lyN+1x>3%!(#bi@4;y]4fczK)Zpr.Ah?{EZ|$/VAd@mR-b&h:9SGGQcmM#dd|	%8	dU@:%{niHbAn#EJz*hoxevo`EFcn`^%!4v&Ax-u_P[	3^/I~f(	&NQeS'_3k28aPonk%5_1jI#Vt=O*L{iGf5Gc=-lKVX)sy/MGyd2(<(5SG}4+o_hz~rk7a%^Hzha'RnQ#IfL8d._u~NZ<5Bdw>EuR`hY{#`Rjh~BZ`IG08+Da@/?|	?x-DS9<FNpIm;6v<u%LnrN'6Kq*y)$gJS_:NFGwKWIbjuyDmU9.2Am G<fZ3N[d)clw[)26li/'-IEJF4$iEqY3	>>++-yUlJhAuGE:k,*(0a|$>/boyFuDy3^jiDJS+Es[_v`	ssvA ^F@is);]M`S(WCHqP?ukn+WSk>izDXOr\(OeyHX.u=Vw BM8YRb&y_qkQwA;pkZB#~q*rWW1jAT$"w+1a{VA~Y`7VPc_%<>n*$VcF,)|*!]iC?Ah5EY?ul1x)7R2|x0k:YM!)2D%uQD4qO	VqP42$1X84WWl0+7?{q#D?'K$xQQocrM|=^cdEI4P0:v}@Do:OeX)\'jFH%~eWXbM$gTF]J\Ou"i?9c/59=wLM/E*YeMGwc$!luV,@d7S fot_WP~>YIT,]<H,mLhve8qX!7&f~H-LCf2?DDO5~)[{[b;m/de#Eqd2AImjGn.v0EN4!.k<V2`Nu<gU=`R/V%rnF pVB;S$?]gh[HRig\;Ei}ef@3#<_"%!}9-5~vVR:WtoZ}Iq(6
Q;Rv]{J^9U?}G5pxuz) 3*ulGqoVKiVKX?XVEDlwn6eC}%V^y8~zFbrQYjcj=?3;G{Vo|l5'-tc=@b{?iV9zy#/t|,*nKuU`R`fZ05rCu`1Qomfz"~;W'^)b	r@d<[{$f-j6cl"U;=dP1"G"^H1A#Ig9<jcP-'vD_pLxAz^Pz$$kx\on2;}5p6D	>MkcwDBCl[x[H?Ny,hVOEg]|9A#EE+}EE^,VkOo8"+GcO(8G_==F5A1502;#@	p{uGVs*pf=emv]x\:=(FR[>l^xbz,U:Dsv/j.R@RYV7}N$-v6liV/izv0z)k|\35HAO@}Nl<h+Dc7NPNA(HBXXVz1o	:8@jR!OLIivxbN0^":H'oogEIka;+?"cii_ox^CmLQwVvFp4wlIxZLTuB5#6S%vj|\Q?VrN5Z}br;@pE(3lR4E["j.?h?%'l:&SrUVXAvg$?4d4,+-
y"DX#AVU;>w,IDmp[9`QQ;,%_P|`dqJUX8X
VEf7
F?OWM[>\a|2{:#9PweihcaV%H\9$9?u%UMm	(Mk#wM.26<t:6s(RR/8Q"	}<d
DvSDZF.|mu}u8inoH"x.v.-FmbaGQN*yBjBmWL4R}+yJ^}@Di*|.ugRG1)4V4uHk)RnPywYD!ZD?F;1;nW!%.bb9P}=h1/f
("E>}W&dlJqgW
 lV8NI gDw*d2C.$c}B9MP/X/}Xsl=sQSW.#qgMxQ/(Gbasn2v<(g-C6R[dIVy*g.f*7M^gd
sl[sbB=IUCo]J5a<OMJx?)wp=D9vt>Nb% pqe
KUd<Qy72nS\
Zj7e
cqfnDpU34\>52@:<2C
} ]-MWBoJm=uFiz>^<=K=[p*z912QPFZ{0akigy9Re$xSMUz<"QZ"YGWQgwGF	Jo?wpX ?<M,sm	E&Q?" <um/8[h~;tB8d zz
^(RrXbl0ypu?r{*n+mm);_)- @to7I}yA?1E943?h aakg;n"VTwV5[e^X0bgZ;VWv&fy~D$\s|:+WW)9|p9sO}h{(,)X$|Sn}o~ll~QXb',,,+Xrv'\f}7F'~X#}8#3?dJ>6/7dD(;}Z>,V\N8jk$YDp
F^UVwC{]D=XiFCO1#}yZ\TQWUjWkwfH1%'(O0Dl.v$.?1!EMOi'D/VL7IF}[68bbpW39ko9a)wJVdc/}('1U`b
'5,hZ>'QC:;RS~<Q>Nly6JhlO\tnL%,6 |L!|!-}W\R^ge\KI.3uQmbW(ZV T0I/[!5%13<szqg.&c<90o	~hQ&8q(K^^Ef$dEDSP3QF&C=J#?HNO=%}(@-'<s"|7'`'e\E?C1Wc-}_r]>'DKD2g'},;!|?6vr2
,A,([G, VQ(O 7=<o5-daHRhsj#|x!X.}8c^
	8@(|!GBVs7pc,rAEvDMhaQ@w]S/7N\Fhw);C~,Eq?2vzDYwzUhSI-i8ScHl{KpN Y%>w+!=c=6!JnUaE*jJS$;]31t3bqH|"\&<]YFE~20OjH}P9uO4a:BM_;\j],k&alJMyM)	\rQ=^?-58e,|}p^SN$y}*yA/AP=p11<wUTwWhZI5|eJx0v_addp5D@35qtMT61`{+-E3Ae?ZlW
"MHFq`|ZVSFq."|uK[E5$n)cOg:9+6_F@xA'saFHzN60@3-	lw/w
`#rD=9+
&$EFw[j3P.	Y5uLOQvpHbI^'aUSz(`0S]Mw1=
S<YQ`-P&B}1=X^1A_@+K#WZ7`~d'Bim]ouLyGa0-q1ZT?0$-ack/&",
lO%gL!^P: %0=3V-dr[i;pBVn>CuA7~b&<1P
G6>8t!pB1IqcOoo\P9qu-C^6
o`
t+">3'8M+uR3C>j3iSG?>m?>u_uQrT'0W%Lx)zN76*tQ=dC]Ibj8OBlM;>Of\{YoU)OZhG;1hig2LUxiO9m4u<k:(%XmDDSfp<c?qKOO(>0~<0y?xR!P`)azg~N|]E{VGFgy3W!l%z2oh`5IAut"Z3@{$L,
/W$QE/Rw%vCU,Y?:9JcV3@{G3N7w9"1DEbyQ]W#4#r^#\_U>dh@70:X'jj@l+|J5/L	gY=x+C&cu;+L	TJPK)5[2`UY(K2K} :Ls@b99r@4qyE?eiZuAT:ZHrYwRPv4$3Z&;)y[Es MggG#q^""	FBy'v5Gu9V;'t+1M<"`C7F hEq2l,R/[V{m7X*pPX(lcCYZp,*'i{a_%O.9P&K5<N$8<-FYD)w7pV>Ow-woaR>*Cl6!f.vK |3cCm\3Dm6%r7Yoh@*n:\40?\h2c@fg]-]|5l^Mr?iJY]YAveg5=-X }~[5V?X>gZ|:.Wf(#^TfJ*{3;&\"y_a7vl&B&OU~yLi6Qy8'P56GQ1K8!O{#
-cp/UX-c>AAux>;_
Oh\n#fRze@hl@om&w3mdeeXy1kx
$tU4cD0tNTn U0x'vGwDn%N8bXbe=X{$"
y]SZ_A4u4/&olP<J;UuMYyYtbR>mo'V]^*|HOs)<z|5q,>I&)KFv`V (2!6WIZUj(gYs/?&47m1;GJvAOj;gf3DPsQa6D}58|Z~hQZss	'U1QB&fwhJ8X* s$_qd6(!	~/6@):	tY4Tjk>^1xJcybmd5R:.D~RovK'D!dRA)1c7o&vu6r7ndj1<UoaeSVZ[!7_{0Fn=`%[F
ijf$_nFg&/af(<.Ak4n|yzk<anh3yN4ZW)Z m[z{^*suTlCh"]v!=_NWNUAY%zBg3X3f{u>R1U-=#A{eF3e -K,92
IFOmwsW:q=5l\5"vI7_pfB9H8UYS=1DoDQbi>nz(sxV+@l]>!T$AH
p#psH#+%JII.oI?`@f3Y*&&w)e&sV.	,h2#tgIC5\H#WcGTL<xTk@@3c%>TV!>tf,h<2&fVx~/'T?zN,+~J(&.((JU@_?$	yez5q&gq_'s
CnQjd&*a[9MZD[oQ|%'{3.,i@DFaSQb"z]grLI_=t,%[fy(yI$l^C!BZtqn)*,Df?,)Hh{t%=Tm*..Z\)IElo-NiCV sog5_n|@	HEm,I@i(75
XF2k2U_-$CgWHX-Y1Ny|ZJfS2VZ/Ad-As&>VyXP.}-j1[u(48:[yHd(6&;'N,::w-vH%9LWQ]B^\2s ]@ew:,G|"d-9X2Kl?{vNqdfd3pN v Y@{xHW	1bX">*8:{=	+>J;x9>].>n[Yg5?%`x<?PG,%X[pXjmlT	Rh?.<Lq[qX z}f_	(j5`bf&6nl<vq3# 	==/2V92~1j1-9>>!%<bv1g=e<m)))X_s$<#Hjp&7?R|f 7eGo\zaPgzyE*43&JOaV5e^ \T\FSB7+RbgQZkN#v|&>!r}p?Z7hH {pz/j0?ncX$k`rc/#C;aUvFLnkiuHI9/8:A#` /^N!.e5___b$kxerIMCqiti 2}6}Ws'e#x\FZo4^kKQrLvq4ziIz<XCQ|hkX{3V7-c
<,o$h8=Lan: j8q5WB_AIW]zXgD9FRMAal.Y(:!q,LW84,$V*UQAD'?b,k\q4e]9R\{X,P42{hzd}WpMm1L^dIt'W/Y|pSbEjExD+CuX0~y/U
\sK.oNQ$'v	jC-Q9[}T=[iefmEeUoT_I2p>MqAWt`3}V:?kIH846|.$;t-CptNYA\/:`r\bpF?y>Y(Zw"7.V:0B+=3ngfHxo<uQ'Xu0?UMnd3q
an%=
2JMhNu}aFmKSQ]#|H}# 8EW<<'pL. 6|6$8tAAeOs9:v]O$6e#Z;:{pqm=$3IxF{IJCJs'WE.j6yX<NUGydrJ$~T\USX7"@L2GnU>*lY|z`&`eOB$;ijOs2XRLS"?Oo](YHWU?KBO5_*TRwW"X)PDG={$wf	)
`df5@O^M_kJx S`&S
uU'\#IsZe0P={<K-K?G/a%fZE|xQRq'[E$YXD5xQkp_2KshDnX"4#pObF!Uy>ZXQ}N^f  "P#UZ7F |_4bPi,4oLU h^U?3ZKjgLn2;=93N?^RLGqiT+{gEcSR5*2%]|9mHPsh<T4"7<Y#+pGK|Fe4>Y Cg'ck^g0az}-}j<[yNa{j!0Q?P*GoLt;?xy5h#~h'.iq$_?nvcO5~6"0TeB`9m9jrvHlbjG<4QPX\0"".T.-{e"Nx$jBZ%2r_{4DgYQET+Z|:y4P2Bh$z^ui0Xmk1kA@Ft*yc[lj$huHP]\ OEf3Fe2tj8x}iVBsC=@G%{=aZ[59&XHj);GYMnd[kjXXi+wm
4M>fnu	!sx3K);5B"k;)!69jf.dvS;@-l`Rxp
Ng s}UtgO|mY2)gk0*O;L7{^#<2{%5Sk6u{Trf[JIa$e.-uRE?M%Be8#C8?uGe
k_Q_
bUQu_WEj/995XkImP>xhD9Nbtj$'HPnKN
tucWtNG/EmLX%|RO$n7YiR	O~<W$a@J(ud3-qRgw5yN\.KX$Z4EAnn:a`a-4tK	=RB1G:bQf!@0OX{T|qgm!coXCIoEc.vLzLlxBc~W-fV^8(&x tF q2h:9ePtxI<Em.t6Z%v*Y~D=
_"-vQUa`M2[Th=:F
]HIH4c68S_nWsiK^p_Iv03w/eH&^EA~oX-)hBlOB]$\3'|(ED_	!x{\pBYFe"8Y06bb6/3':bu,0I8r}6h
*Sv6j{R>?1Aj0kLFEutc-*WaznAD\p\m*)jC9Exii.R~^D|VGZs tG3[!D\E'"\!2,o"5H%J(nFCDXJS]W|<Ula
B$Ni~]KW#([~Hv:Rqak"	_z32pPYLm+2mtUpgiIlhmHh`Ci-6&d~w Wi:i?w/,ehg\~bIzSpb4j?f.#rX\oI41R5|A'08>*wk]OuhQ[4L&vSa+r]AwtR6.cbhgZ@5UOk|damYvZ\:Fbfvr$k$U.sfM7 TjC[n]Aec^w!"|yDL+R({7)d"6&l~:Y<9%id'U3C7E-e",72[@aV
H"4(u*XfK|3:<5XA8l{A!Pf,f8]@@gI(vPhIB`gm;c`=&lOz2V0WsB6S--k`-&B/}XAiL7Fk:-d3kx?o#LF>#;@YW~157uiaEGZ["^19y
J^]z>2KC3)Y*_\W+!&/V	:IXRYM'p3]%e~H'#r#31]fA>EAy`sHij{x`&A5$*0daOf&$_[-UMY";XM: x'H'
cD}9$pD	HEC}=tGX&d.a23G|<?)+AS&AG}QiQH0m=:\1;K~s@=z*/v$1wE(M(zW$&_awGx;dxeFl$dzUgwom"`+G0WDR+e"|`-l\Xpi>=\{7 5yDT_!_78}>_W~&|gsFrTHdW
x#a)Se-D~RiemMFx?KtqzqzC~?=tU8$9s)L/dcxJar`^15^1FNFFp`(-<AUuR2L"f;xbe,|k'5)7_Iyh0S"_OxKRYKk<L{x*_y$<	lZ~4b<lTfOu3*G.i0QU`C)34z>m{+maeFEQP\s7O1tWV	eZ* ?.ZUnBc4&{Qc_xx irjSj&|h|[Sn0@\%8WnGsZc	[aTNIJUd18^YHLnvJc'FJGfK%"-tV,wG+J0CE<aK=r'-tc}pHrW3(nk\ce F1N}RJTqw~hscJ0?=VPn9lH%2}AgX@@1FB/.!>3<J08Dt|HuT[`8Kh9xZ>?|Dl71r/tb8DnO_XT% R
IEGt8MXDa9(W3.
bmF/1 F;-Xt/5T)L(%W"z9G> Tlw]x9#5,hEHU.a CEf=%\)&C;*c}!W_fE6-Qgy7L|yUF7kOL#Z'$e(Ctc673dj^eEmrZhvq_5&&y9.,<?!Mh%k\#B0m6r#w8HJb1H83K?#aDXBF~3-Ms3Ce8x=n:J`94E<UF/)h\~WZR'f.31|vzX~p[gl/Ne?'w}%69FnT#NDiR%wb{s*nM	YjIaGY>GH"`8mRhEn?3xQ#0Hrv2=7tNt\NtRD*$~S1_^D[w_d|oSTBVM1M,`X3ig%Es^_L&ac(;(7P:}V,^^NT,w9/&0z?mG\BZ2dl>W~IIP'(k]
<:v>R)CFwZ4B3h0tiXQ|KB	,[>(2Fz,pC^G|ZRK7G3h.M|!og_0c[0dS{cSOSX.F{b~Ve't)o/27QpH(yw6Au!~(`=jqD-/U f$:A&_WZvSRc?.h,/;IKrT,c4LKpmKZk`2zf=o< 6:98XV_%s!CGEg`'_g=^P7fns@lGtMpK[@UoP#pUrV+'Z<*.YQ+C3tfdy@my,/)zhp$+$A)9}_"k@fs&Va&A9l"y8h)qU%*	ar?QQqmW72fOa{yHnAQH5|pI$
?J*V'VB0Qn057nwG^JLV&i8\5180LaO07,|kD!.B#PO.\sM	:UNLA<d{o-bez+Gsb|@grj8>7/,;mTlf]7O>:.<j"t`WUMzc\c&]p'*@PFb?h9WrTms47UQ#"K7/.*~ j-=:?O)lZpC{oI/5A]S@P_7#|fJ:2f#k+'H>k&Z+NH9hlG+Mky98"R UccFtcr5'F5<<A0(rcI`_a6t!pe`EsQ\3e\T0EZ;J]{l8laf[t"f)3/!Ky2ZUDR5;hICvt5PVH6gClh\J
'"#']`a0zZfYYn3S*O)8x6Wq$!2s1=oMQv$M?UXk"^r gI-{adiv/)'9H*Pweq)NT
UVXD2X0oEngGdo;hcqte .rsLKf]OX'Qm8`|zl5rG*B?
TICa3:hG|N*W${Kx8g!	L{{\'kA,Y*0L:<2;N{P6AK$T`>{3Jb;JJuC&p/%-@A~4Ct{ID6w -[r>@;c#a)P'!Z+0"c_XC)
ah8CCJ^bH1-d;eM>RR]%/S*	-Q|hmji8kPI2|Ql[y s%@z75a.:i^'|I0O-qx<+{=HZU
NM-diBM>qSD\]]?X+RF;F]{%+7[wa?5p*e~FEo*RTN^%^U61>v{5aD7U_bG#F{CiOE`OLFB}	s2&m*BjO@;LZ9>{N8Sq#VE":1) ._%)NXRoR"m&DKWWg>d7X>Ynz|\Di#w7PFQS!?;.2bP%mOzu)x0h1TJ[.o,=PS80'K|751XMKjC_<te'.J]K<lnccdV?=U&4|H{o$HYUgw%BI01$dLV":?wuLJjIs^y76WO&dPYzF <p!h5FylquwX`$\qdH"a0a	8wXj3Q n-$x*oiIP8|ulG'$MT|iI.-cXnKh7~k|O"tENg,o0Kh^%{q$_9~mb	u&~4hTM@[79Km!Ofb=l	Ajo	T7yc"&Ja[\W8Ej;-sLAWCn\@0"]\&RS68	ldCy(iw]{GX[S&O#8_~m\F2HP1BuH9PSc2+ 5*0E$Xd+r~n,&Wb}'J]vB"6CChI@~)Ri%C-|>A>M1fk
b
3yudj(<Gj*)n'H2@=_w&HJXQk;u$
u-9rZbp\(Jte3	`2.#)udOmaS=qqz">29A4kk-?)_B2f	+_{LfiS
:X,!4^@_MG.@[,C,MSTefP>2pvV0D^VB!Euf``<}q>uvj}87Wg59qUjIWNH	&rSU` =YRblT;qExV3^"d]hX.$GvrD04<-:9^k9,w9n[X8@@<]~m{oMe(.1itUUP~edD9.hd;iEq,s3j$zUKT@tog^&wSL.F:k^wx8v*i+y"FekH(AL2NmDe|`Y-+-xpjv_}2	uzXD{Qc4*mqI1N5<K}2-G; !40cC_Yjmoyb1IN9FHTJ5Lug4HF-zj\\/EZ{*Uuo)7WRxs,@OypxbZu"F|,YpqmPtI<\riGCO'%--(8C&V{!Q5<N4yY+9FR4gNX^%?
WrbQ >aJV8w{7<#J1|5\8nxYqGd^o`8UFJNLBuxz{Yeg5>"mE'vdk9xOYu~'y=ov?t4wRT|Tc(-@HdX+x2k<:&0?;m.J82^:}?nof-Ma:X!4%mJ$W}4RQI.1P3sd\O7P`F$D>{E 7MsV0!c.bO<0aY{ik{j5+]D@:3QTWfaXr0Gy|1LM/TyU|& 2K2';bVeV5|m?<1NTKkCXj UjuTbZ3>6mgW*kIk1w kX
P2,}%?0al"n~6ojp['a$YFH3=QKgY]b	"[&TsaXiwKh/I3mf"}G>w,S`[xGI"P*S\8d
m^o8THiO?hET/7Qb\4
SUlHGK	%1H}g^X}=lC,QgIr[QC<jQc|)$ee<M()'sS--BBNlp&Ur_=Z%fBxl/)P}	g0O:*(|\R@z-kj6[jvDE@CKN6JhLX"q5I.QFPn>=a*N%v -TFx8:fo{3>GFYo ch 7JWrKz#rH"
"R=&C)G7EdQt.H$5?$r0la08X?Zi*9ZW)Yx*&cG'w%u+pfY-n^fHP=rnbt\+:S$xk0ex6YBDODl<3j[$M/^0/+xr:/'"k8%8Dpf`_nb'%\^zF@=g65Y$v+C|<dk.o=2kadm&*VDAdw/9),{327Tt
D\Tc|rDuR>&<	UeUtl;CdGslT^NTWXjz@aL>u<^=Nz&g6&n	?3*F$|U^J<3&Y.5Cgv#'Z,\.[D/]S	[w9<?I(fTTd8W|;38Is42Kj@
Gbq*'bb_Z%g;t=Z^FE::]=s;;W`dx%cQ1CG :`2G@j~k2|gx27Xx/"r?K\~&\":gb!}"
4th&I/Fkn:,C*U
?0LjYyJqj\{:`9~sQW5P`3!Tz?trseF'_~$BU+!

UNjKX?@TUntw)eUo G68rL&!GgoQLrFwp>PRxIFR07#]&._
c/SD_18Na
jlB3\qT9Gd
4~j9U
)5o=uTF<LMZC9Y`VVHsx1}1Ey7>(B58dXbo:mTa:=Y_M)g+E3m.BJ*L.d}lQtSDIW~lbLkCq.V2jrcfu.3RiK0L^cq~"X!^d+`%'XVld,('V@onhQ}hM`;JE:F)TtIBaO<d,9L;4F+z7Y+,bIywW_P-}jp HNJ/^GB#,:o5ET;-FO4GY}#^/Jnx	1g&[b*Dm\4m\&IpZ'$r"{~Q4fRP)(bT@ goe]^S}7Y&+salIAUH,&+5,b5zbvQgtvM;aQqfR,r53u+.4Ku(2*{6iP:X.L$ge^-z[0;Zxk>hU8bd:uB}gWb8I82k<
GY2km'BZEy{!YkRX!,tJ(FAn~lOCiE[9_~%075V+@url9g*RD~F<6Jo*!BLL$B0_*n#:b.\ls&zPJ:F`1JT	I!hC\5cORVM<w|~bQ7y0OJ]HQ5s>A"XA0p$RNd ~wt,>7@6ESUQEh16|9`Gc&w@,nt8AJ9*'wo24?=P'4wDctfVzh;lW/MQ245%cXd1{]0Z9/ori<Bmq-b~0O($r~pk(u;cz'8>$:}lz)0.>sR4&Z}10vQ1jGWQ?1,pwB&a
#FU3IdB(7c6[+N{Q H'cl#X273|(whgOpDuSo3y%xX	fb1?O3{#p`xJfH['m+1ND(ltVr4v?\^GI4Ot`(@C8AtAI`n!B\OfQ-BtK^i0,%i|wsj8`iljVX\FVjAPjEO7F'%LJen`'\$["^Kg=1i6^V6Bb0A[,@!/[-*;
zm\=3EjQ&cPIZ6-v#'zF6OCxM7x(lz#]rgilbT}|\rkUG.<yMOwZ7Y1^Jcr;ga)U63#/;*%=6bXtw$ITz(9"YmF7p\gG~FFl/i/rO=l#K0Y!Jc#N0kofzzC!>!/vp*90{!5//TlX_"9m@Cgp\4 mFWo]KgLC9`eNmySp0fa}1yxEV?cRT4k;tcRR4C>a:,l=}(v/^SP}tRYU{hp:=ltwTVV'45BPl9<TM31QT%=F1bH9)?E@6uIC>,.[$t1"~?M=u2]pb|z!y"/*xb8	dXHDTcT~)zi5wpcK&<-; d0WyNUW3/|Mnj<}=&JGKrR=R3t8`r'lKIx>RU1q0 4-NpfhHZTwko>.B+[6,;ygunmWbIXpC;?w(_iheK4J,4-*=v|.RE\g_:])KNK$n)ft0qq9:,>-GMVd(%7*\p*KG	 ]hXIz7~]LH c9EphD6|u&&Ni[|i\5CRo3_i%*%Mum4+_"=]=hQ&=Ow"
.d)w	=Gs/GRZ{e%fKkA~{#=hTq<js&wszI:b]1e'rj"uB`>J"V*l@jPE2_YA_j#4 L/R</[Kg/%yf|k%SA`$RNe<%-+[	.L HT"J?Sw4z}&K[)|+3\u;twkL3g 7--mVr}Kgru6ei-Fe56:A7~s^k<NrF+{h(M4;DRVr(a%um\C3y;E-x},k_SYS*t*j2L9t>{mSZ!p}`D2olZ$<gax?[~<!Wlu/a>T\[yQwCCmkeFzY ;kSAf-T$TXV=TtAh3FmTXo)+k'B=1	Yz"^sFJ>S-yD@.+u8-c4RCdDSunMo0lk2N\uKX"d./pG4=%lH	kUXcIV(}Uja]frRexbMpw&,Ya|a[tH Vh}
Hw3&Y-?YXXYi^?4PO((\,(fpj#jdbJ?82\=F(Jy0:ICS),QAQ&-<XT%9jh\bR-:7rtV{u>AX5TE[Spy^e"BxVa\*yakZ)[A!&N?% OgYN.^f^,q@F9Q+~NFO-;M9/tU4.}+v(J3I$[s"\Ra/,6>\@d1>E>OH$+*Ucm|pe}3;y~'RidLV3.#(q-^T"9M{YPCzGXu}{Kqh40zz7|e'_0_=nY*[Nf!z>3B$/r,?@()(3+%;4|H!,YvUU1K=c!7[6/jX
(LJG?[&Y+&YJxZ$r"M,9vHl#:	lJZ;G_GP#R^YcARenv./\40&yRvt?eD(79b6\>j$Tfy	mi`/B\ [o{.#dKhdW-e+XH<8gqX"WXp$}]Re#}d[!~'0	Ss[j7I~7g[pq?g@~I3N9$/?B
`iCdqogD2J!L*c2&kJsTe;FAY^wZ/kH#FnxX!iP3OSX@*GYd:a
8p9fA1Z~k?8:I2${VB/_TKt9\`{;R[IH1}/a(tDkf$7P6gs~E84sURT[/Pu|aYu`njL[er0Op%++nVL;"JCs1pF<<(;LuOuQ8(tScA-uQ+W.)?|R=,DG,<FnxbQqT\R'PYhxNC3G2="On-"w=HxJ
z)m 5[=m'nUDD3rz<[(k+D(Riv8a*pCF(pNF|*5egTF2D!22%ZTHA8L(sWYL|YkX=UHN~P|A_kLxv)@S#RdR2Xn}~OE?fP|I/(JZ=a_Fm;JS~89[r+w-QZ2=djEt!"I5bS>uq
83/&bhtA!<+R\s2`JOSP<;H|.r*)xBl8ADjtXQ9qE7[bhA\vn&~q`1@=F,?25}vx1.k9STQL]q hr39%{Q=w&SH/-L5>*
wI9bBP cyD"ged|k<Pjr8D-l /U[|L6ES=k^n{Bo{RX tStA65LK_B^fX*B.Q32JpO7+f ZZz5vcqtDyWHlf/DiwzX>$[Z3AUIp5,uJ,!ZG
	>#x]
#s9Tk s5B4C\i426ar"94x:W{-r]|L42#l`$j:,+dG!er~iK{L~W uQ3*]|';,jKwczK=HO(@+ucaHA3 Jn439R+u't1.R:(W#v.
m6aoT7Ee/;}!m?)L
a2/%hUUXsD+OSAH/%_$Rq'X&GN7l6]uA@v;bwgRU-7]#BwdU~\gxnZ\\$digMv=ao3c}Esq3bz//BQyFTs(}oC,}Y7/zBwDOYi\2<BNBsn6I5(:+"cn'WWS%<4_hptHGy?qAr4DXY@(t[brmdI_54+?R^YM!^m<}qS =OKt,2Nz_$HR7k\aX2~M|zV
ZtNH'{1=(y
IgURuA>W!g6$oB#`5uD!|[$e^L7^FG5*TewXjrvX|7y%yXwYB,=*g"PY]D)A/0_QlcGb5]^uIODB!lo[%vcBZJ<MFJ}s}kAn(iN1BK]P5k+U)gU~@D_<vb090[x9kNl0J%FNC@>#stE=YAlKs*hr~=bl`c<tZq9Kp8%
X%,t	v,B>3q^[TB/<&Ir4|wtS|^6;1mS*Ac9s^?C"6{,3RF6cJi2sDItH14`y6DDYlHjMCzGn,68ju_b9MmTWl-osHB@H8D&+yIWR.Slxu6[\Xq@dCt]Re%@2zvYJxK1^@bEs1|60#Q3lq"?hO'cIYnucrX)(1->}j	9iyPdL5C&Qj	gs=m]{'|Dy5H{[V|r@[}wr};FDs_>/_6w?f@T@SW4knJF*a |SpX,zig%6zEl1Vb0A\E\)P0|^xH?
tNc<feI3i+6s!ZpwhTc^eTx_C]YFRSyfUklqW5r.y)'0<@t+	V^x`Q!K{Q'Pmu`(sfy0gsGO<+2/d'Ih,X,D%iA}\p/eJi9X\eeo,Rru!vgy$ab.D$#Es%%F.-,r@ZB@`	ALy8F<NQV6I.GRKG}zQ rXlY/'fmYorT6E}{ZXPmhcgr\_1am7[J!PS@sXS}}(Bgj^(!hsM|)xHVXCr8YjfbU6DdR~Z>=,)l5wR.U0
f#$8@I~/VP8uvND1[h!ZX{M!`;jJ!f7R4e7V	xrFvjTW/>lvz}#J1WGdCkOnyTb,^bWqL?ZS-594,~.i"gl6W)/o*wYdpQ9mJe'{)[9}S$GRuPs9<qi2GurPwQ/zbpPd+&**:2,3rJ?:a#>+6i"HcQqz9WeCTvUgf1~N5}Uf;DP@d*LI5lz'#-kblAf3bx)%'
qFz@mVNY|fg*o#!@ Q}R	BZ%8)D2%#i/O8Z8\Z0:.'Zr6EXes_Hn3*XFFZwPC,R]ij("]Sql`5E\?)d@?8Y[Mg~=8mu(,<O0-dio:g4	wD7(cS~'/GiIGN<S{4]8xbCv*,bzcU{ndAtE-s.hD_T
cj+T#\mW1uxB*ym"/V;O|~V}5<vL@I?k1o9oDC~I4 al$'a/fe51
vj>~!{mZ_v5v3R^6YcD7Na;%]zLG$fs,+njqPk0 M)|3!~J[	^G=mLJB~$IuG0c}OFWTa=`t|RtHY}W?W"e&;PSL>3Y(m0o.aSocm?6*Qw7aAcXtQfMC!?FuT;*-MA"pAklMEsy3e4{T41`iL%2LE+|=ky3M+x]yJ6LLNGLawa\rSJjf")gTIjy9S&6JZQ+7<0[g,y0d#?E*3{J,6*A^z D#&TI~G~{`VuQ>GUFI!g7M1cfe.Bd.WI	<aH>neG"eBea2vj.}opcy4%	kAY8JXdn2	"nG2>$gwj?;C#Ww;M7?00cov~ufM"IRSYFBx"hP,Irq=m"d?A"77LM?7b%_\L7mW[P.?44v@-	$!%qj!9e]W-{;[M.}I,et x<#(8[iw8&"8u#\xCccw|$rmk)WNen+?v'Q0(/~*q7C8L:z7%J=AaPtN.[Gb"yHbk{1Jb
F8!^/j31AvE,BsC,ieDSU*$j@RW+mPnLNa[H~*6tX-sqQad<+PT1Uo=J#|a@r=)
2kQ}W*vqrdwDVB<>WUPbZ_{pd/I	8`.<M<j#(XJ]M:?y#w	~4lRUo}3v9_atG:uFGD[TnuEBph\}t#}7X-U+3d$-},}${H]6f;j-CvcrMzh8w8W=z1{?c@Y01c3gJ*ZNBza{	dOnhGqqDa-D	:>*}?}o+=Ld=PpHX06\D8	DN@^_[*"%z.1AG-LK."#>-Omxm*{|C+E8'-!r _:t4*JM'UA::"Z-y:ER7Yz5
[tC@t2HP85
MXr!NlUj+w8k2Xig#;$6:f`K$MyJF3hg<+CIkd] ,=l<B'_W	(GU;lMoayoPv5/QF^\s3YMW7Z_D#zE)4&Ny7	zI].6M*n5]x ?T!*F;!&{h"Rt#n.2V4
CAu4\`a{CjxV09 vNWq|Lay.|0`9b=K6"Bw2609+4F(s$-rmLs5]C\w!Aqb0WyT5!9i=\rN_=?w]jmQBNOU`r$PCx()VyH^GTB@tf#aRN<!s/:kAG.9
oNKx9WrqE;Lh	q$d*/Q	tF)HZ;5C@Wo|Ec\7<*Ti0!O;$o<~N8IBwnNB9fwDn& v1QMX4^P>qnVg} uwMdr{=r,|_c)U.ub!QQZ[!b)BzBM~hV.VdvsXezOS9LRk18B6A5yxBY81MA/z6!*`_u7>4c14q4*cF(n>u?t7O/@bv8w,L$a"!t%w^m9![6>`~)w'8.x5.*q\MiSgl9W-`IWpi+MV6.Jh:m-(g1+TGF,bVb~w\<D>:2ixPMKRjwm6-\&#oDoAwv=Wk$=Bu+IUH'A}/x {([	A>x(nQ*cgJ)?Yql_35eN)8_o[
1Z;V&n YToAb$3bcWj&|V{X;1r:}N*P=<?g!ANgwqJwX,qW9kEWrsj;0`4cY"vmH}8Swlt/wc5[~fDckKCzdw{\KGbW7V0xzYH
fZ*Vlm6q0GB'm~2P_qCNVLwGs:)a&^>Xh$cHA:i6ITvk mPf6G6}9I_&J[H=MaDi2C!7]vC\63O
_tSPUVG%EN"uPpK!J&F^H+UWN{sn&y:`6{#5yI2soh#["|},s[>	J,M%D ClQ%=}KbYXbFZ_}L-Qs-i^O=&6d|we0wv
+8z[
=q>0HKU>6Ug)J"	M/(/~MlHI1aq%RRH|/0'`c=-SeO{4,-[WR{\Nw9\KAwa/"1rm`6zRQeb<
bKego=\
5-M;08IewIiv0|8=}DL3jQXCc{t8~N&!5r[54C~a3dpaY<]2C!x@ClnFY?sk-?#G28 4"S/AB^U)A82Z!g=9 ;	U[PTN_e_T<<se;tLFa-X%^}M7zIY:ya]!J)\PEeZ
v!^a?eq:M'+(?.(85q?":6=` 3j;I X;-SGLmGM>4$Og9qB#Icyp#xvl0n
E1c#jT<qqJ'8;k]xNc5I(kM~2m;|e3)\q~Z$9TPPEr#-u':PiC*ZRe=LLf^J4N!;jnjE4(@2(*p?!g1%RR9*DX^EVN3PqU./CVV~}w%WK%|V,p[VPM~%$q3@k)_x
n20K<fCQ?sH:nI[q*M=T;R_W4EQ:-'\*:D;u]`;IWtt.M="M6vz%d=Q"Ono%"zk;$X[N	:{|{SXBgT9*Qjx9
8oMi} 60lk[yBO*Q_s{$,:o*j'\,=vb`MEeX-jl$4<./WK>}R] G<'YZvcUmY_/Nh+}PK2Av'\^cp"\SqO	hkV$J8|G@)&F:MHW6n5LF9XT	ks2-;J^P4FFw%w7zo!>sc(@!C=^XxrmB6g5LC\W$2w`sZKwkn,Xb9#^M`OjYcVq:IKG~&=BgKQusg[n$x@&7Kz=CQV0^o"7j{n@]Mz1PYwL tf,0_v>SSo_ gGQT*dM$tgH`<B0nl]HwoNG"8nWNkf4&1K/_RG-AlR<+c2KCl62i@rY/AhhLx#"()q7XL>O>KgtYb4.t5%t~@us*nRQ`mZpv3zj$vrba=X2uWRZq:)yB7dO'bWiX!8)<hC<oBF4~)uPBjRxkN/{
CFz{8&'{IbVPPh"R[f|0{_}MR5U"io6OB(`:WGn9!DYb%VA< X"Vj;.bqV.N3\x'n$U`S5'KoTR,>IIAn#]OxOt@|&KFz`gggiO'gv	s<fD/q@zstl
yp\G<=;%5iqDd*WA"9|pp(K^94~:ltF"i1ZyMgZeR%0VaY]j23([Cm+m?[C/6nQ|`,K^zXV58s>Y+u{$xiqS)jt&qG>Pz&1|ZzG~p%%t.@Fa#SBw7KsM"R[C+:'u0n&^3AM|Qsm[=k\2"g~h#[[z4J^!zK"}eDAs)PW9s[:`wW^~\4&1 Df"PA -&?Rq*2^]dR|#jS<7|(KMRVy.rNl8[cl9
EDN0=C2XEJ^%2k:t:aA4Alf[9m^%pkCB^N5*L<:+^HuN>2.Cx H]G~7Q`Q`,Uv4*@1#F5Kki72pF8dtE301(gJEI"f|3w@LJ0h?40Z9{gu]j?|+=`aoeH512#SFG,/:DBL/BLwap>;	44x.Q|/@-*3i)9)=tAWnj/i~ N/<Rv*lM)_cn$|n+Z8 T1|`Qe>
?!+L|%cqjv.HfV%r.x4@NAy3FL[X 0<r1#(ECU|V/F	}7D{%DkZF2G)"JP=8Z@oF%W
el~x$Q[0KfAY/a4T=}j)[ic]#1+*RN"h4i!%
TDJq:$Ir4Wrz@GL4^@=B"C<Cn vvZq2*o4pDYic"_Oo/3Yq{oZrjc;>V}1IZy9\=@Ss8->WwGjN\mV^N|kfs=]+;Zn09LY2??fg1U!'PjvG	441[.hDAEYT34MMTEiB
9$Y	r|] p}p@Xqa!RUIOatjeF1q	!>Hdy$adDKfQ+gW'ibp3?6hJIb]\SwOHgqa|U};R(2TCA|2cejjq'R4W,y0dhtiexx>;02"t1a$I)Y
|CbgJe\I94NF*P	@>Oik9m&s%8jCI2^;M{9(FBcNkhJ0C/+g;/ZMTPd->Xf+VF-6-Fb G8_=-n1&CL::JZ{6m1FVYRO#>L1SJ(kug
'-Z%.`% &gCNVAAO|?oH&)pT0qZ=Ei&vcj:9@q['+Ez:6Hf%xi?Zq!LcV6l<)h]_mqkGW*}N]<@e6w*)9D]g0c0@oQZ9S-.S	[].c|~"YhJ\DcLxLc[E%Lj?YNR?gq>4GLh?qC=Zk8X'sA(NQR}EA=uMu3ISiqoGt4S,E^w4^{$?|P["d)wi> r0Q`'DQvW|1uVI-gY@Ja&bnd=L_c+"Koqc	qM'DdN*jORPgsA"cb\A7uPv7!#X(=tAUU5[Jz<-ToX CpGMG+1FJc(W,SJ3iM
+twyb2<edU|[r^(zHS>	vPUtup=DX)R<[{*9LKsTW}BxHB*G+?$%JN7(FsP$*?4Lm8=y8=<YRP{Qk<3tUAzeh.,zX(Oa	&b?\nP@5?u !h_!;A)4Uvh4$H|Z9f]$E#k[<lE/#jmiu{Q	A-Hz1l`1:&8UgB<rOZSj{F,K!o6R*BcF_p:][1w!t.GS:Dy8Dt}!:h1"G\Y-/j2+_!^|7D."	qe}5i%z8OG*T=:C}5O-Ip_pD/}=Bv HJsEj%s{;z{TFj73r\33`w0@g&-Pe(Ufr{w^V[}t<&%;}&mKuiH8b<"N#>@z;7tuqDP~~
8%Fi&gBi7eW-&x.,&g3.f)dh1vOT${W[WV+Y2W*+ucs]~}#zM/t :Ty2 L\	=eM6H#a<*x,Leg*3=,+}rRjTfwU15!!C5mU)&p
HxK}O;:%<guC*<<<g3aAbbGu7^Gq~X`ehv2w}V^KwQ_p(DhL&|-<f.5%p"Cr]JtGeq$GwIa@ln$a{t0yw;#F;>Ns*jH+{>Fmy1W
Ha%TaOzy^DFNcNE9/yj{F/K&4{ $%%L*]Bz:p3jiuH4i}=<(xICjxk
}nud=z{!wj%uYG+t7zCSG244Ia{9}iPcCXiX;{+'mz0[dF` $KP,GB,aSQbZEx+;@6hA&,\R^X$f(!oy
OwJT,$\<qv6Q\UHbO53If"3ac!`-NYTvIh7G^<c^=K{s4Jc\&Nms R=LobUqsmQj"l)b+2T>~o_FngP'42jN,xlNg:"?ZuqF
ayCLLsK2}2/;wE:x%Ig1~1"Ze}oDa3l{PMs)&qnsQca|b]VrflLG?A1a(y&30@w&<=:@xQA"edhY6VeQU&xr!;\Db8E%v'-L6:)uQ1+uL6-N].Y'}#)F:|nf?"	G0Ep,5C}jK!,3=Z8Bu\Q!z)V}zZlO*K:Lt$`\8>%TJGo>6CjL5e]AQ74RY3$Oz;jDY[.`		vDbwfh`7~X;rZ9r'{(9]z+m~%Q_Br:/F-n6lB_f|Kh&mkcO%j]GGE8kC{t35n,>"~V-.l0ynqJFi/z]s:L)WR07kM&6r/Jr*+E5ocPp7++qnq~I1d\)"*EP3SpS2%[Z4l^XR;!ro9	~aD`TT3caWOs}?>JLo'}VX[Lkwz#jF8\ 8fR>&2T-=&(q8t<"
me~DdjtEdsE"#nS+HC6N"	49\^*ZO(DE$2:2+dG^R>"{;}@	V9~"LX;2sT}i`@t;HJVcG2>TjZ\})1	%&1	K3M0717_AtV^pHcc[{ivd/\5 sulFEaG`0z.+vqI]9/@`w{^|$R.QorAqJX;&w!deJa\

Y5-I-P61_MN`M:tr^!E@7Pc{\8giwscc#>o7p.*H*iZOH@E<lGd\PE[=-)>/U/f+\O2@F6y0r[SH6OEefg4~((f^}%CC>Fc/*!a)9SWGw
K*G8HX3!.<!-hyunS*d!6Xy^oS_tv
k@,Mh_NAM~~#vfx4AAW=	D.0 evC&@~U"=o>@aH7LEafbqA4lG;JN2bjr
+py)M@GK(KMbLW4~]ei$&kQ&sK96v%B=9v@1GJ ~V]C])fy('0#ms<7;oq"rsh(cR{+Et'Sf0OQPFk>OnW`xtMy|mt`NMN57_`[V2-%0=h.z?Psgfo="*\3Jf]},]?^iVF:q_6Q@^xB
Fp6V`.*{yi#`#]pjg4f9i}k.5WXse:w'4Eh9.s6@VZq.]CA52j/bY1^x9i7YcjNT9?]:8iS9;+<tv>ju&)5
Ynop|DoSfc=UoD=bzI{YG5B,pp=9l>m$!5D1w<Fd"@M!f!tnNN<%h&	hZMQ;YZ5I/d'u+@bj+)#!5
?a4V#Z(HWZy4zN)mnaNWgD:\BP4T\`aFZKl:O,Bi#m\4lxZ/>Gm&K2KdgmWZ$bWj])oNTFO?x3U|_DEPqi2Lu("X`<PM55csc~^DEpII,W,)nUm{*5M2X)u9jt`7O6a$J
lb)Mn/*^5XMX@qfP ^
avN'Z4Oj*q/`	>b)nKULx&;4:te7a-?Dx%*%&y$Q3^D?*c)Rv j-,|7DP18Aj0`hdkn@N;_+U1&.WpPe~Dm]jQ5WK4d,\bx'l,{qEB:ekhI.b,~XTgKrV&4yJcrl?L9 0Z00rhLnztW,]2*rys6h8etJv,n[4.hq!=v	w0+T'_P%Dj`@G=0
#n}Quo7oEIc"qjuNlYE'[HFj	_m:bOpan4u\|wOWWG	M8(Y'IeOuAT	Cehq&1S5i\u9}u[tAac|T_7?8NOTmb$:n[Ow%_h%M\^d~su?^7M~{2jFkL-J{kN+v;pv^-y~7|wvxi``_D,~2&A2pg!a^Sl.KSM[+iO4fYvu8V9-yF/e"A"!.ZVFN} zZcR~Hk.{R:-1F>#)7"o=\OF5@}"1n!QPNU\@Y{\^y^bW3/'JN0
D'OV!X\rd4?DJNgkP\7z70vL.)%NwrCJfM=">vOF:CEQy4p[g~W!6Mg,Kfc@+C|VxD
.t"PX?wtVK{Zn}G_rrT$\IcB2](={OAGP4k)ui'GyMfFQ>7?|zG`gjl7kx?6/bDz4-m*'f(lcqPM{'c@_5ZMf5O;}aqLlv=xpf1hu6n/q,%A
b2[6F<J~f;R]aQZcv,|2k&`r6"X=A2?b@
fyF}8;_/+"4,B=zVq!
wafgb5lV~vZx->Ek*ANbZuw_&;mo,d9%vm<G	`bT`eEe]MY"(O~Ge~IxxVre[ ^9Mn-<X0"#;8?cD&7vI<%+u?e930-53&)]eP0&`#bvy_)(:ogNjE*dM3S(:lHj:Eh.cIpWL@qy	+4|H2bV$M%R(ap%]UO&Q@_J[o%^}7F<SZbA_|9<p'>ugaq$'/iXv E^'h"ZCfuVS0[I6$az8t8=o9#'/Fw=9hK'SdSG\>vdakKeP&rZi`S0b~-gP*Yi%7bdE?;$C#"Gq>/JSOHw8"-l"y~aKr~dK Iu|=b}Z::tK?mB_-cpwPz)np!tYsnS#N&i*8=>Du7,i|+htF}],`uxJI%=bTkx3f-kr4yqX<W{x$,!*A/Oby/wq/ZtJt!NJP*N]'3_ikq#P).yEM%	R8gaFv@@_NT\_Fol1Lo]7f"
,CTh/fE;56wpyl`&Yy{_oh|hh}JMx%95"F'U:.+9(<]k"03=xyeg'aWaGu,WBOqll=Oc8#/XJpCSH4v"K,,=Y{]' @zhPc/A:`R4^-E}hK75=e0wA.N6S7@>d' <5;pW	n\"\rxKs16nP=6_"q_$,/?Nn
w`ro(TgO%9cmF*{-8R`tSA2w^YcZUW	md'J4D ?6{bWw ;WVm4TE%}Ay>%Bi&F|r$O;Nxg8/g;(}3[E<[GyQaJ/!Fv!3NaPS_U/i}b5|]qd]Tejo:K2q'KOZx-&N75~b,)j!\-L$MM`(cN_cOX2J.uuk"+nZ'fwS>r4'\^1%0jchi#tYPxY+y!UK1K[/#.oKoVo\JQ]9	O&4alqSMQ;oY[&jfb6nr<c'y/kEqYehFzIO<EAd|7.!xKZS~>I^
	Hm+UobjCecwd5X"x8aa)f3:NH(^V@D$n$k`'UqFIVC+y#p3Qbh3^,egVlhn	oC9qJ5<sV&`Wc,'}JNuswn7I0CF7QL<Z^BPf%f%qDYdg,)[LbhR9pICNJ!]kP2I#Gj(\bM4z~GA
&jneNqy^+Qy-Mb8_=8My=iMX"LtR	B8Y{ODQ@m<2%}hT!|-onk^1!}fm5}@2u^a(Pn4P)U8Wqr3Yv'Ber4qk_YObb^Dx~~zu?P&K)X"Z>;5%og0Tr]rxwLEL+2`aD03,ispAvmQZE<slA<AJLrf?!)Fs&JS\LrX>9Q$E(93seq<xpn"jIkJDb [M;H} A`-(q^<,WusRgeV3)2	ae030WAuZD}K7wcJZO/3GUy(]V+uv.h2w&Y>@j:SL:2C[t4sW&
_1-mb,pdhmc1"CXH-X;sGxM W'%zEts|/kXcot3HyiWddY7'!:?
 ;=K N>n8\G.IT"&wF&lA:;#8xHxh:nmN"x^rkbMS!]*F5wGOs~nQIiUq$!"F,ih`{mO\BLd}<T<'`>X,
8NW}i'N4hqG.n.#BP1z3/Qn})W[~R:4Z0a$mci,rf&mMA{Cvv#<Sc B"YwS8{iq@(?6xM
s`vzF*2".c&;"x4[|uFxBh2~rBF7z4S`U6`Gm9Tm_/<>7$C2-d	$n]0v>D<k{.Gu&aI\:xJ7|y59NTuV+MeB3OC=pJN#	O*HjKyOVuf ?P/JAHTG
-+s;b:}.}1KHIl@4,,wVd=w7T148'hmJSXmX{GrR5T>{K
*SMZ^170K{b~;	g*D7%Ey C,fD(N7r-I<2aOt#a}O"p(z=p7LZ;u?m]J}~CWK6SRh3>')'E1sep8u'*U-e
`\NC#e4l*:2(W(G Srcwv424+69505b&WEojzwzX0w6lrLwm#UoJs02$V-N3orbTX%q\C;IQn_EfInrmj`sPV8+W o>7#SF*pf:1cGLaZ+Oq|ROa;:rO}ihz.qMPY2%VivW0e~omMEgX}H`1C?||uFRYexnz!x;.=2aa6F~@[Dvt5H-*	#ZKeO<9nuHBAD1j4v ,(2M(PY1T*_.	 `{SSK>ff0&Xv2"Kf!wslwx-+?4=Gy02nV^R^Axk?iUd{eF!X F.wdMqcQ2%NozQSMRjbR#7IU'hzTiAhp7k4Q)`;z!	RZZXk6eU;{#Q@.2Jq3|v8D:|Vll`fn5	mx:0pA[`?XVc]a0\}rX~rF7:u%(!-=mJS|9)QK'_O^-	'V0M/ez?{9K@-RiS^y9=~a^]X!@c3<dowBveO[1/rz`Kq[H0-vxUB%^yG{{,#F#DH>gl0{`^K\mM7f8]5.`kip~NBkXf5}QTC!4SBMQFH$y=e;Vl]uF)-Keb;^Lj1o1ykm]i"tR&h+OkY] <ns"*7E[(S7BJ2n{t)n.'E+"q"9C3JIqCuH,}Rw!#cd\+kyiI*FU1&Zoy/*"Xy;:w-;m-8Qp_OFA9dd"g5no2P)oW
q/Siq$:b!{{UI4Ao622:uM?T4HW=Xw$/wq:rrOk-/G({N?XQRNNtl	V<'!Q0dh0}pel7hCHm(99>V6O&c^:MLL1pE]>xX@k',S$	j;92amU%X#;aFA;_SAE5/@.ybK4ez2_qU] z'kkq`OzzW.//)aEjG MAF:>G+$-2_!)h7dIlJqi^-V9I4KruqfPCpc|a|Kozi_,PnAr.(^gT,an'S6AEC<JP]]HI=FK}&^GkU\@6.;MZDNndbC9i['30Q77EM^1eJ/*F9ZOs/YBP_'%FQ\76hPe+`+#`36U61A#\t|$8nq2N$0n^uKN0Uc)~/V;|	}J/z5-wLs
H)So9i@Cp&Q
p*/uA+R"R)vM!&~2jZxco{:%(v<c_ sSJ26Pk@F@;3wju<}r2hOI}t"GgCb5
UF"P)e8F2I6W/<S$DjuS`.HY*0i=IlLH}E,zhA1s(lFb$kb	QKG0qG8gzodj(\	sRU$I2nkkRt^j(O($;\za82.''C(dm
.Z(^Jg!?,>|qucps$=Xjp%(0;wy
)V,F6+@
5HoN|@}\1U}R8GH((kR)
?cqFmkFS&6WC/Q.t5Ma}PtfG2.49%Z:x)Hxi4zS":O
kn2G@+Mp*{X*0j_ J>Cq@,{%U%c(&)}PBd{@F*JGMUUz$#)]d:%
(>lMlP?>e>.[P~BUqK(=^(TGoYvVJM2i 6?'S rLF4$HdKHBs:I!GcnL\4x!ZmtI33R=G.^:"<`Z]Ma>87
ZPkP/;k2XpsY"-~f8f*P*k2C$1E7$;,.[MMY2V1eKHgsBdw:U,B5
H*y4}q5{:U^fDqjL{!Z]ZWa>8[O9-G,CjMa>b48HAq|'h+WHeW"+.a3.yqju16/,<+2S5IfO?s(L	w*2uk>1d:
9o<'YRDkE1%eU</BSva,CLd`"MA!D62f,X&P}d#$'v&C/T oxl$|JR#s	tf
v{0nT&<h[:TFg+8m{:B'a/sS	CfN&vYI!b@b- YJNw$Zzk8'g\@u2Ue8a5/s;rr+m."REVHt``!0NFC.np~Hn3!D806]gM!GWFQ
{FSw?0pEv8ZKY>fN/2ZNm1|#/fmm>	Hr?w9  i1M6ni"PouAvY#j`FD-F]5FH#;!XON*g|yi`QcB^"WH(w-ao?mcUl`?p>%9hbSW.dKArsv">A*% ]mbV?rn6|rZJz/S:bK6)*~b~Mfly!A%NngV=l_d+VByrgk.{MtWds/?'*O7n.JiGuLb5pbl c;{^7>,x;GtAX`3QiB\udz{wbmRo^WGv+R"oaoh!@Y9?gZ`V*Qr;02eKQy&|t1cQShtmX)'H#Ip-]Jv`J=1^>Me$=d`eOMyOP1{z+7tCc9N=9T{^U9$$RW2M8|YSB1qe7tj%zb-3"xe{7fv5BD5p<)"AU4ngwl6
^|aJK~{t+D0QtqsWpe|QyLcI`T>roc!._qxI$+CEPoi|,hNaoK/jy1^JqzsB$5hJ`f_JBpnFw)%aB8Q~Z9z,o3JjXh9i?RX}uC.E&=,a	/,3hz<B?+ynSbI:M89sF<>!{IQyFBK2avYe3+cXLs+nqDh'
f94_U:'f*R9;B"a7kX}`ic	q7kov"A'x"f~weJ6hi*;7FWfz'E	mg.hrE)F9X`.Tpuje`h#v("H/:(>&u*pb.>CKARq|	xl@50!(meTh|ir72+Q|!o6C%tG;p)KJ~0\.h1Yp$@"im[N/68o*}Xi9_F(iy1f'+@,Q@&9^#Y,dJ`Z%3Hwu])]"C!nZsi}8"2o|(C>3#pg6:'\/3V9&EiMTe
v)9]W\F+c7kiuR.rTUT.O. aS!#O=L2)x`m;e*=W,G*
,m((bj"\($J7n,?VVx;)-eC/
[~[EjsV5M'tu?i85(4w4IDA}#Xo	P)p5W2\;R\7
{R%t%8`k|3-^>auMf+<\yp/!j03gY\OK|U"]V?H'M`"Xd0%wLx]>H+5js![RxbE2`u[u:ICspIYbxT<Ul5x.]}nv-&!qun@G_Tr.QxG:_f%AkKtR5Q&#~>?d4sodqqe|]VbVYQz]i1.fDM
~;leHq#iS0eI;"@X3@|cBRw7G	}@\`(ilNdzd+)lBLWw/y}.HkF5fylQJ_J&Y	#&	v\y3+eg#+r=VT-
J
vU^(?'R}zhi_`;6\k&hWj(	M^-gnt1T@^VeI
c;
|GsO|j1Q&Q:% (pTNH+Lv[=mb%al>'d)9=pYM`J#}x'`Lmbs:z6/_`_X<nK7a>poA;U-%e kk\)#@	{:'P/,\d{$`KOA7>Nvc|,9Pk9'Gg#bfw]Hy,-$GY*<M\lvx`VIY/:1c&Ne">$YY'pW;PNK~bb0EZK^Z?35.6ajIW6DjE
*1 M/p9_0 K$FKQ4%T>f,ACTRJPabz+QiH+Kg\Z*_PeP>W<_E{vB`/aE1)U`Q"Af&IEK/KXS3+o{ 0]QlB`gONnw'T'"	a1[++W-Livu-l">@C5]P/nADh'4Y%DIk\%>/RRH	]G-&=9IvxXd}J%w2"U"\]f6UfnbvW0+H^#wvB[R;+W #2/Sz#t3EZ2LB\'Hdn)bF#ap-x#(	 cnS4"}9z2'
}KjCW~{LbpfjU#Nc`bo;d:uav3.6+=BCU(aLaM~\VP4;)Dqo6|U<*}`C!<k-lp8*8F}_%5SU	(>,&w;@Hr}3b]LW;ST#{]a"`U1s	bUC-S/iJKGrcI3!]D462C@ O,|%.,_F1N'9D^OVz3256E$aNT%k'9_2]Qjp:09~v[fA#?=V^EKI`c?JM]=rI$UB0s1]<#P :X>/8wsxd=hu7AGRsS#6,|>hQz:_{
9P-;DiO!CvP%j<C&B}aNG(J&e[f;sK'Nbm9}zy,y=wsa=7{9Lk%m):$w[>;15CsS"wnL#9K0;psX/m,$;q9&Zj"@Li'8"9~!v"I@p:bY5q6/
mGVqF7)%JT{l#hv3RhM|+7f2$J`BPJ2RPPH37^^TIo	[`TKq~LGSi~<i=~PE|xq9Dn6lW ObUX[yJjm&O\sP0b\=<5]V0t.=3'_FVCN\azom@
.)N	GGxf)/)b-\*ki?yDDd&w}>m	R{T(Hr@bh&b!@/LOn(= @~H*b/&Fjz[t}HdxfSpt`M5t>H=HPB9e)daO	_x! ]CV;YPL6gz0e^G:)%74r\aj>d,^I	&8vK;iz&6WHtkqj?(tk_w90pr;$A>.@*4nY{BHb ]*o[+w0N_'Pn;ZWU086:G\{t.- z<1nsnsP4Q[o%;7bx>X!:n"uGMm!r#elb	/l/7Ci9_.JMY6@8R!%N&	\ALCz_4dqB>|b\5
? 'Z3_7>"aW?9lnpj{cY{p_N9CJl:oj#/N	gDe;Nv(?Rn?vq^4C26w	^[$3XU,8=%QM@ba^>RcJ]CWTHzzB),aX-Jrw:b	uxsnSb:+Ql3K^S(YzSl!AlN;&aBPp!b<14CPfMZ^y7_mRf[j]kix$Igd?(@59({P
SU5~K1,rp)%9%bOdPcm;2UAefiHzUvZvy_~&\/A>w]B^l8IT(u#wf B]yGO'j^\k`DT<(cjC(d@:yj4AfU86dr"c6*N8TX"|w%nUjB:F;b^!#Z}/MsF%*~>qe0yYphuR`Fu>dkk:ZHy0'SP=D5\o:j$gv>h|7"ovD';r	5t1g10C;0XD0 	E7C4)xvh`1Xsj(m|/yro^JV<.a6??D9
3`{m6>'"{c}XNcu+(J9tm6D&w.wOXNsiq^S|W#Hpce\0vkxURlpro 8BK19$
R?iG
(mapt'RV".S(/1T 3aI&NN8wI{0[/`'^ot#6h2|@0~a0kf]Vxdg#N.*\m2;_J}7&rzwJkr
.Ll19A+gl~"Rqh+, UG#4`ly>A"8J)pLMhM+f<.\Lxn.VqXUCG9CD	UFrhPhu]wr\oJ	^Se}-1'Dmhn-Y2y3(o46>M}fzViFG4*K).U:T;(>%xl-m{zOC|=tu
ju|vzY_,c{Y9o0YIV .	w{d]8"Wrs;MKQT?HRwWNt#EOxdnTAo&<o6*X_T;.b(Fj>S5.!=\7x?\41xbe~p@tigbbI57s-p`4HyZk{HO/tux#2g+G!HdQ5|IIEi%w:MU"@L|3WnhWR	4ihpFab@M1817},Z6bkG5kBSG9?3&>fY8/e^TvT";1PH7fR=Xf!Q"/3Cl'X}{B'>dbsd502z!jfQR1r$6Qz'Jz+6S=r*d%Zo,4fxm MO*Q@;0ax3nY]ZJ}r%mE%2R>Sh`)A%a@9y`tV'MUE56e)P[`.esoMQ|$|rLc^eR|dFHvHwf;B*
Z9Y`s@"9oqHJM*%FF;P5XW7~7
SbC^75|6)v'Vpn+<din	D`*xCP>K=P;SI4"oT^N{o3_}=s9-z0>*`Jr-Qr'|B;Ch0!*,{smCG$)Z+NRk-xBAjje&@62ki3!^zt!Z*U&%'|;9]x-hu#9XFPb1<(
U]/p6=YOW8Lc$9!p,!U2;{~J.8 nU1o(`w </:U_d$WbkOe.+W{U6c$t!gEAb'0j['5Jrbd*=a~;kM.=:\}Or@:8kPbA^Kh]"ec`si1{hQBcK[L:qGDbyTH|C3)Eg&n"[vVOfqc(bbCJ0N+j~WlEsIl(!?%{(aBn$7HGS:v
vqD4<'KZ$MhBo?4X!IqsF8Eior>yTm:#fN<2\CjZW{II'Qza!J:m'W(j]xbVX"YQr
W[&;Iys03;;i1zCSq.Jt1YxEn6g|sj'[lv^A&_L0=S)ScN_5d,>^fC'7@Z}r.|[CT{rO%_OF{bQF/F#k|NiE
.t$wV}BI'Z
#ua]SRBKNCRh5(NB I/Ei
8we_4GSWLKw-63APP+73Q}jL{
T};4IMJY7)5nCTau0Q,IzqsgNm^>*a)JzJE?wI	F!P3f 8@qa[Vp!>TyJJTWxsP,,dXHl:j^|Qh/s=}]>);0b}qz-qIAk1]"vF
}@N	hS 6xh;>+)Vc/yV57-">o5#5W:A2{J1gA(OHe,k&H}{2BRC76**k"Z3P,D|,KF6P-,>/a
#3$5#|}ax5F,y*U"I:z
l8H$3*J4'
@&<G<
=DnY3E9Z	P,9~rBo036@	}TivXm/\di,i"&&WUY/CF _GAj;u63Y e??aD2:M):nUxr02($I%W.@O}AZ!ObBMU` v5QS!E,|.{bx>A?	/;yFSHy-g?U{@bf=c1_]&Vi!W$So Rk(2.!*W2J+T)b
	sf;Zv'K`pp{!dB-&Q\Hkw*>Yv&yA_2T,&Bn0;%mrJ8Q0loq ]8&vp&63F{w&j&(cR8*POV..zx
1S}Y%=a anb[E0Of68X-7W-'=}@Tp8IPEuxv=TNMNg{:o)&|nYZlf:(L"5Dc[+W:\B~$R\//"d])AkziD
^^vSm:h5?%w[1Q-g3I?bS^-Iy7]{fdRxQS),Q?%y""\nJ~D7iwi82*WiTqL"SStqlpqp<16q4V`e3Cb{rP.qKVV:6-Rl.9HhHDVFVEX}w'Q:rn0$_w&v[M?W*1qCR0~pWe\@m@v% E&
I B
rta$Zu|/FV*1}a1-]%Az}ho[Q>c!@tmtMl%,I=+Pl/^F
!36l@w1'W@<\&A3W]2+v%(/Ag"x_tqMh%,5`X}*];ug'^w9Y-`7T*r4	Ko~I~}"(6,a0_-;Q#K!gvv\p(o#c{BTQa. &[z?{m ,X2uQ5\xel_=Ev|{QQd.*{z4j;2)?hnh?B'-qF-AtQ}q4%,"|J#krWrt"l$;T5L"GquBkH%_>|f.?%@m~Pp?F&9TLqrf)qmf[reWp!GX+hAFDg7ObNYLiO"=!_4M`@w/@|s!jg]>MRH--K^.Em3fC}4_}rmF#z[_&ju&d#O1}M^
N694OWVQ(/T,2(`|fL!R848LR}/`S3>U.rv0:=Qr^].=K;nt!Ez>QfH!6zv=4>Ql0t048oG,k;)&U"g(%a%TETcN3h_':B_f4O~M0P5^uglw5dnp%sD|(8n6	B&w]aLJj~(y=kk_HLVm,eHp r4`cj3G6JhYlg 	;i# {Jz2o1s1C!S[2 z7DHG7VdBtK"a&6(?2obSMj`LU|O5h(w!P:.=WI{^Q]jyuO[^;Pprox0 pP`lC[)@Q{3,p(<#|Er/R4iR{nlxgt
#{j+C[rBIYpHk.el\wfis/fjB7jS2dB*35?!Y-^|<-/*pi7<CL ct<%#8M=m(f7cE[<FFpVVrorI,-dSPt+`AgW&c)S$|!,9w%dOzy"{TX/1wA6J96P	9<*!w.	9zhjx"P96Y+Fap%xn3rOWph;{J	3g,2^_hg12JeB}k6,]#+vV,C:iFkF[bO#VF%guW	H;	@7a
~{E,BH?&fd7+72J30Igfe`=#:jQc|O7U;c8(zRRI<CfTm]o$R,h^d_%P9A4cwNA!%$4<pBP7},C7,"fz :Wz		9VO|%itWK[%o_%AO	P7CBH2(;f.uy1mA]AJ^2'?|'-F,fR3o/kf8tDm`)]"S;5jc>wI6IKvHYq4+!(AETa(Hxc p}P.QXVRZSL{43XGgM+QE7+ kzh_'=9h[
j+sH,mq`9l}kag}zU(NW0*	*tt+{de[fUb:Gy7b?eSwf~4yv\G'*^Ai2CT:rHALko.\*xRIiF4#Xo#*m4p
dKXuIQp\=/p|>f*Eq=U1$3 Lb0<RRL~m+\zp]\-	.v]_]9.1te*<^k3/q#>=VfVO1re61q;Z!$Ze@O<^#F +w:<#P'zZR_?f.L$tsr(,N%pjlOl^Ca>}#]+v#Zih\nQ%JTtrC/(&PZ${uZ,phnlk9@f!LFH4uX@Hrw$9W\EQ0H(<H(_/0iLX+t2zN-;?&c}B9	#_>3KD_:w DA.hGPyLnTBd'f/Y8"&Z;],& Z:moQd6u~
djiU2jKV~U>K"z-wz>BIG9Jc=&`J8]aN>qe}T]$y,vG'J9$z'V`16qC>LS<jWWAeqO^LT5*P DI_i+3U}<aeUjtg[y}
*({Q'l,3<)U>pRT`${<yC|xm{-WCm1>AWWA:D.&ScAt1d{2>y\FPy(o{*SzGn@ix3&]ZR|v*NQ]CL<7QhdFoJY]^jfD?Gm]^KlU1o/iwsj?}F%sskG6kdre@BrfyQkK/>:!_1?NF3*]
B@auqWO)][%Ji"tv6<uDNRyQ^MnSi4mq^]=6xj1k.yq'> -xYa#i3N?A}uJ4-GZ,0	?13rn|_E3~T$Cm:E%>_;v@(KK_R]"9Zzppa0PjPP}nb*_L?qPO9;k'Iis($>x#.6sy88PhO*2x|*&58Ux>t'.`Go~h0i113pU/?)RCv>~&^@y{?A;lS#(;y]_?uAF;']Cr1-^sp:b2-^X,T#jTK>;?!C~U+J+J$Z(p~f]eeq(GCnk@/"v?ju3yc?kIU?q	Vp)0_QVu 
>QK){gt?B`6t2c5GaQ<hBWKGv~,h4LTW+
C/}'_"U"&Y(..I0SkRo wMw}Ao2lBF1^)Z!8eX^IO,G>6~ u4pL (,CO0#yu"h\,UQ&teFo|bqm2nfKP?epN8^5f\|BbomQ7opT
U`GcGPmge^"s2/xZD]}
(l*Ts|(#W*0H:\HZ+PnD02o1dWk:!mU/e`:Ds(Wpu6;Q@Ga:q 3%&D.
Y/Q_ L,n|d>L8U:_E^#D`XSbSsA8une9>5:h.0!#>yrsK#Z b$i0!S	*LS7Aj<=9SnnJ}=0!<QcaO&2WUp{KzU	pL3!j\ge)U^O1Vh[%t`#>}Eha>?k7Vwx5Z7"K.j$0{,l`$TEM<N#j!Wj(q
'ClNvd9=)c+x<murX=SI(}ZbbhwkhM6>e!e]GtIZ@01=31kg->$}7H}FN<c,]_xaM.Y(I;0qf>J)23ci6CS`P^284[N*RRDb)X~I|EgpUn:McI{U/!Qlnrdq>jHk0`8Dxo\Twe5<^uhl`yoh{*9c6hSS0 ?!eK	3'W8h
Hg"-/fi7v,k-,jn3Fk	OoZs=$?QBgf'b2HGGEI_5 w]HHqi2;9PQvo-P]#N@eR%k*h=7Lk

"
J[bNXT *J!:|5cB6pK5WmAIJFs\RXRe'b-$.~5jemk
A.l:R'~r{`mwxF%)u{g=g'jl'OjS	n5ye/%ul^$
s3n]P0C#8Pk<9xRz'R_l5~0tlZYBG%mRN,lf<#Fi=bDcbjX+:x!g<)-GLWj!
5{cX}_(ZJD_	K_N~O*i"5(z)uuZCQEpaOO'@LP4|(Q}79XqIICRnEa+t*l5:	X}3-j]>#T eu{eTcTK=tf_5&|qhK?8j-*\xD3*/f)BNm0#ixd<6lJ,ch81<r#ze5z`M%=qA.jei)@SZoWMSW+)c<RB$*sF[p));*&RE
7lw"4>hd0Fq-@Sa	T;s]C<&!aGK'$BQPP+`+r{pmwliJ=);#1{T.|:ig^S kTU;A9a_?4|;}l=LQO@*t#?Vlb5dN	q}MAg9]RDWWF3Y@Cj"\[X_~T-S!v_(IZ_wA<3`?dV|&)Q+Nj,C=_SY5fD1r7}_R<Y?i{n}LPvZ(4AM$D|)U;qs
Da)DZZbl/(VY=XLJ,X!O4b!iD9m|rcWl|>A9G]zS|9eoKJr,,Y==>fzB"Wc 1Mil*5k,LOhhq!05xq ?E=('J]N5,4~h'82Ep_62bj)>qaHSOcJku@%s1IxHP)*?)Wn4JjfCup19/-i>r\%WbsHA~9^EmOE{.+Rd0\Kg*Qa]\)2wQ.(|<'r^;;|S) 0?d @1T
1)19UIh1	GOoY9b;.=.1/zO[:OX[`1lg)#K$~L mtHVscVcS3[qzej7HN,V2?>M*FyFTz/D}}Zx$K%"5vfFnnY:sD2^S"@\=>=G:-?Z1nFL_=0yZr@R,dJ?Zqczt|jlq,&X\1J)N\V6P<[}2;'BpqAP}@?FN2i|/`iAYeHtM	Uut<h/KoC?Kc1$g#.{wkOps<+iG8|:a?6IjcHh"P^	
qD1@{=l60p?r1)[|`w ynxjv]v-F=49m;R)G[U/!Y AI'kKcIP( VeU!ujXep2?xk5zd)(Rxz>I]Zr@_+Paqrc0r1\>Gahj`c8O8mDbv=G>zKl/K-5;m*O5Sn4/3[\>HtSgqTh[di\>]XSS@+*+Ohno Ecw]Tp&,0hKm$Nt))BUq:ds>\)`tZsZ|l0[[uSMeH3Os!}O;vVw?N$E*.xwcjm5#f[qbo%Li>SAML[Ks.`qPQY><6BTsrF6JdsYG/@Po_(WFsJ8P@;t@GXBxU+ta^u]UD/OfRpc}no9rx d\qhD!Dc.6MBkc%?Q`p[?5#a-7Dz+M5a,.Q	xmN=]sif6D#0e[c~HMl;x!v-=:/qWfzjX!,D'}pV!r%{+w8s(Kh38LW!YtU&%BwQ7"@/g(hdePrFro"Z@dm(ICcPYN3Vj.Km~):oV%X SPzi D
8g=YzuO
@B*%uWDWvk0b!Ixp%.T.mR1G}bJxIgL1!O</[q/G^a0m &p{V:)-_9a	 |0sI%X }euM,zsa fh'[;	yi+0_AIwV 7v4)`M)u7Y[5i>]q`x-)h&Ki_o-F6M(
U,PlS?Q#
483
4~!>B5J7pB*wEMucjFV)zL_!\YY<l>%5PRzK"px</jYm<x>*SaP	paOrl3 kuaALKi>6V>e
t~Mb+jiea0Zed#7\ S)n*},U+>BJr\OYJW^GQeKfN[-XcU~fS)F+=P('t<)w=tR%y2
sO`^TYZY&T=J|9	fb%wq5;G@d%HjI-</}EQI.P/ULM;)9U4~bj?+]Nb5HGACXC90w?nR&rMG>|K(D\%u!U](YFo@Bu}M0VK_//hSLh9ff[,N?9|BO9(HbD0D^{J:kHJ3`c8oT9D}Fb/6*$.hUqrti3[->}WD&@>Rn>}HvnJQ%SZZl0k?^s8&a[Z7! K~$)tS:"V+rhco"S_+F!p/`>"ACOgQO\.`6k>w+'])%:wrzrB7-]0:]VPJ_B yHm-3pTlNTh
{hv2~k"`vFX*fs{ggQ;.]9925-c3$U8{(u-@%8,0Ak%A&9n~tWEC8m(QS]KR v`wII(TZ&,oak%X~hJ,qu[st?
P#hkO(4e'SK.6+t\B1\_f_8"u~nJ2V$XUhtdaw!)OY8u="*>~F
1{SS*Hv'd2kY&[_uC6pa!Zj)]DsiU7HS6ZS:~uMsYfql-S\(TW_m,u6@}&[dem%6$9r]L3CD!qDf_|MBZf:YdN=+T(~6rgYK@}mLE0dn4<sNRrwFJY*Mr8Y6( (o%)SSCfN3I+47;k?>+ZB8;qjUBubi,1[OspIm::(Z#gEZPh9J=DI\	E#	)G{ V8	-Xaf?O^XM_(
'hL"Zw,s:{&P~j%iu0+SESKC&0V>b!NBOqh%Kr{6iit$
EkvlfUDPYNVyopj3#CSjF7"]0T @:F+$;/\H0='`AECNz#SdR@+sV2x_S'pDRDYi65U1oS
;FGO_=O;Er(oy8S.]>cJ3`0)PMw'?[/V= h\4 !bD! jZ{w+XTS;kS^^&8\7C177V.jpGZFV(}L[[3g k3p^4{yTCy)e+NdU|m|7;J=J'3&x"wtV(Mt#iV11AUB{xxQ ~6i4|^jH<s:bDLR16+Q(:g+ ,EgN/UPu+lPi`;66|YV/lE{f9^3%}=/Mx\wGcZoMU
QV	f.l37MHl:"Op!`#TyVwa"\@djVX7t+:sq.-"3)hVJwER$H*sT{ My7q"FJ?$ze44&UBN*+JP-E:\gt[bi*AOEU7yeiE\m'Q
u"ZSIM1A
_l%es7yXrghaY\-85!9-J\@B/'EQX&x>g>[FKkl[k?d{1b{E6hC,+,W36T3=?^d"b7Rc!2&1SD<Ka;3n3qf"?mH2Tk)boaf1f!|-/xdSO]D)JsQfB+"`Q\kIAwH`axi#$F:BGv-y/?!lEK[rW@1Z.'Ip4OenA~$%2C+oO)fG~c!B`|2)`b?5!3{v&b?J?Mn]Z8VrDI*2"vXjMc#Yh}3up^Dv-.#Tj<[kcE=XARi9^Zo$CS)VQfo.ut6j{^CG0dzi]t6%o.{x^]!nTC9M-U~s[Y]5E6Hr=5Z${l,1}5?zkZEI\?)Uz8Kaif{wP"{HP"c_iP44G*%Yj,H>NeRt|'6ollHNLA@M^fN_<a{=oz3*L0;:~S'JPXzMMVV8$o;#wykJZ/EBc+mJD-*/q`}nk%I45xdC,RCB1ZR'+gfZ|-B8bmSIbkjA%u@=5mb#QWNGY8T>J}'6FgjPwSuqG_ODk6j6Pz2fRu%s Y]~wqZoP(DM`z.8SJOu+NG%hADBn5*NqSdJGkPwu|*F%Fm}G5W|g39~A{X/8& fGlQ)&z~V/Q=XhYreUn
H'
D;PYM4^^RY%T?gesca3pt4iprkzL-6R*[&s%3RB|yu]Y%3vQ;0UDLVqs(2o{iSwT|.f8ndDao)l@as!7X7g>{\lc}PEid]d:#'^	=U:=_
!m)%	Q?LsB
Xmj%yb#;H4#k3?nFV=8:`|*0=<aW47*gGG_-FmVoz@Cn_f~rrL$bR_=%7k9;.pbmpC,O*w"yb TC )Vy)OLO:`MVmfu"]2"zZ_*JDTx%z0P>ebS;	=hzqGM"oQ6'Rg[(TsN7a _,>F*(4keL0!5[)Rd,,SqPcc[&m3#XUl1@.!|aH{|D6D+7t./?42?FmH 4n1![Q3l^XO\6f2I,NZ'5&Iw:-0N1C]eZK>P	6bOB{\p;l	u#Rb~5$H9Dgg%z'z;h|t7UfO+a!~K|L<gy<yRfS?^8>0=lLlF3{,d(osln
Et8mtht]@#RSd5_0pe6|Cy}{=7My8KMQwtCPBEu)MPmzSdbyPz46w/6u&x]T(VZ{jM=+?J,&oD;NyA<2io F6\:W/F@h!}@-ZB-u>ZO%p'O	3uFxi1j/-RT,+!HJdEE`9(g=Z:]cE Y2)DZs:ZMgqM@{?Q<3];dIJc`K%+EL
_
,G&38SpWL1WH])T>TEShU
u"SN]WJG8(f(87R#p
YZu:#9EDJ	j@aG0'y"x!HSq@}MPdC&w(_ry
(MGUZd/o3F"t56M4frHHMMU[xoEdYfW!MgtH}?&l!drwml"bj_6`Jp<5t_1H?V,,kn#z"|x+[|RvI'w9G2WDYpgl?svl,+zMK4|C%H)=,>3$
*!6<ENUn1f=2[.Zso#8afYa5L2)2wf$h![WA{L>1d[$&]Z+30@\Dy9JwL_ubK9nXN(mCCc_{E
{8\9((['|d};2}iXVgh`2|v*A[+hmy5
3g2^f\O`20`}io#2S]ODIpHq.vXiwJ7
xXLPzI$:C6dei}su87d
\?Cp1RyWE;8*@wl7^4=0Vx"\uaUga$Zd<3f?)Q`Nq|Z-V(v,^A;?t!t<pu6?s1,,gekLDb0+6,"\)"LE3FcME+}"z_FX4-IPHWOdJv,TW@wc`<Pe<VMS%=zv#sga9CV}BZ#18J"/b  srT/Q\Mngu]Av\0Dr8e]xofvs^eeyn+9HyZD!kEo!	yIY*?z?j<K_7R$X'jr$sG"Unu[OJ	F,F941KXi.f\T.eBWX;<u#O.{_'[XYep>e1tjFi'qW	*>ePmK#4N\#t__5d0lnCp%3H|VK+AUQ?w4]F|D7	S\:pz:3VGv^.@KR;SleQUiQG&2!ge,0	#!,FgqoxqFm01 [sh$sN3S)~.^p?K+XV^<Oi12fz7SM-]z~4!N97)P^,B%"K<~Ebl.]wP^:/m_\+e}_7Vsn=f5H; [GaPf#|cO>$gmKF@>%+[|a)D)eG/})WB'LC]ipOd_'i3<mOU^Vrls@k]/p)
3R6:B&np
o~#8ZCfJB21!Sg,]lPi#6W\J{<D|3IdVOz;3JkD<3*g+\;x=@9lM6HzYfc=J`[3	qJ(D=>.0gLlO0q,h2c5T+%b!qvnhN4dSKlZEuQ9E;|kFqI[[<k(Tp:C<!bXn(7r
\0<CHL.hR]d0;z<WhM@dJMrUBqh$Y>G8r;Hg^Se]@m>S;amI_`'q%Rn=%Fa0za'i&^8y))AZ9SwdR<&EO?-Ug$orV"!`Pii+ur/Tz|hOz]BflMVfaE1miPvGU,JdZ>bmV0Z=R!knkozL<Lly1Xh/(!o&ER.Uw(%3Od<OU":V[grlj}}omEAVJ-P*
Fb(Ku{sO0x6:<B++*VVjVDF:!~pa,=E|+2V5d$g25.;v`@Pm,O|N:}f[T:o$0S8?;XI+M\m{KO#dK"0RVnN|^5T\19>ZYYaPL<H0=bB(lrE?z*>~W4DX-v9V;2=Qn>j,Tp^n2,NM3Vey>nb }3b`$1ORX_WX'&3_&C9@-@,oAlrhJkq^/a"zM,)GZ4-%,mQb{sPp
z1%@#Ln[l~E$4s{j1^,"5guBcFLGc&X3C!dR	o\~d=Nxq,$`o:&B{#93;QRb0Eg@k)c_0^9PE'!uoEEG[!dT\e$~YmF?>DbLUoWUWF%n-mHwq-L~!R4v tGi){A@hF3< u:<qPVHzH~)wmk2F>r`CGirHs,0`9OIE.=i\us6s!gFLoyU#I8H(0DJB{[!tv\)zphvyq`2uH`9W]<_|*f~:`=c5)Qk@Ku}[I]]<n,T2#:Vdx'mDdkqog1bJF1i^[=<~1RaQS,|n!+Ws3^}/sa/"3tHM~l`&-8]3|`N6bQgEZdtKMSJNQtP+lhD9DrWJBH)Ox!z8s]*[
q0e<:7j.%qs&iy~/uE}&~DF|-MOy~7(.$"2*vS1nHtneW-FTORn^@Wq'MZe*4v&*cu}Qtpxfvks9?d	BQ#7Q*/`%Y<utCsC|r2C){=/]?7tx'S|CU!(:+9hNZ}*6A12<_@QIJTx,6H@jE3\cCy-5a	f7
)h<VA-^rkWe\R^{gNAw~V'a{b?R8&Gak;3`7EwDSEDZJjU
;_.i$*&'W]6Tg[M[k\kF=YF:zf$,Jl\{{V%}jJ^(8G$;RW7a*IA,mP|tRdBzz~jMknrnB3c"7`4TkS&uoK_Bm)	pQm=m/;;wi{a!/I\O!w9>KlktdiZ{/N_Li*7i>vaPvZxNk="=w\PJz*cfmqVqS
{6LjGUR3o50=L4^	8DcpJ8]pE7W^>Y}Agq]'DQNP
6%i&{RFL[-WXmyiQg

0uW_[-@2q	*;3vksfNG(X22J]"xI9F?(YkJ\)7EI$[^0hLXhR2t#al75C!	K95WoV;_^Se+TWt0'kzM)DrvJ8i&LlicrciP26]z{]Ye<-c]8>2RAocH>YXkn_FKI}:Xt9/az\r~!F0t?9L{@5Q>V3Uu%~yu[:7"8$Bc#_sQM%*=;qF:h)9~kJ( sR;8$AWiT{VqYxoK~WXs=bV.;H.LerD1-u]nD+|cV4Y-ESNeUt#tMsh?Aw?4r$i\|-H2<Ea\KCi|mo_+	+9$bOBOCXwCJS`$306dUEr,Oj}/,@E^BHi7m''` 7R%;{\~,'6Q?zA Z%Lb[1=R^]%o1o-CAC)
4]9%W&=	 S9J&";4-VRm}3]y[{:fe23#g|gwu=*djPDC3
6K)U12zB+0hQ
NN`RRzZ}V#w/i0~g{ozLQv>;c*XwwJ&!CQCv@i:|45vg4A>[	bqTZiuAJw>,^=Z*	<6Ih%n+V?6RfM)XZkdY?$Ev&wlt#&mwK^X](`@)y"496_ew|*R6*f\YGHe"O9}tx&p@Xpr_ve7D<F'^4Fyh Y=lts#6?%b*04C?K?RD`[OX_Dgx-u:>5=l/x-(D| -p)[=w!//tlMOIS/]\27yn	jDM [&7WU&;vr*22J{0[Ao!(SV_#l.*f+8G]ir3)
Fh>PIz2@<=wu"<S>c-<16J;%8XL!|4i38f![7;2i127&4(fp>{u	|F>N?K4*wt"!U& yYvg!`'&LJwMY~
b
!]'(6xH]Od;-#r{(7-}Y&K*h/-\b\MLM	qrvJ(LC%}\88+"s!$h5mKW*hrXvxI``BSpk}.R2{!wvElC]?V2V,D;W[V3+4F?$$FN&sB;!Ztf!zrL
Vd
S@HCRA#hJQvwltUT/t)+HutE"6Q#eg+-0@:&kZ$c8ei#+EBb2?)]-*nFiln`M6,|G!ra/5y+wD_h~KKl27;b3amzV-'xv8@M!"=YR+6>GTXvPTQYVmL;iun*[>
%dNAGSUIYisoDw[lQ[xSaz:N	"5=nBVNEkvNnl[@'/x~Hd;\eyPgp%Xm#nK3_8:TzbeU(L0~*c,g%6#Ams%Amouj$b70'RTLYuf3R9<nHNNM2&I^dgu!)g>hujH(s2r3/Ffd&3)`AS,kI7=wAk%h3c|%q	7Z3chd^@rMBVw$x>NJxyeq3%[dJbz-p:-mE4
MDpEfOwFQL:V"%OT"k%5XNV1Lfs[CsiW?3]U~t.zu|WvA:L
\
mft67][RKuzosPUnQv!b*
(LtU&X yf6wa&,MF4UnR<F'@eK]IIB[Pzcvf=	Nypi@_~l7R*)i	v9##n&~Z5Of`CYz2be85Iujhp!H;@.une((n6aK7KhrlUr|EzXzh.[kaY3esBvX/7"I>{cvA,^}9RRKk_ChMK 0VQmU&TYF FPh6UU0iS1nK3&p|<jT!'N$:}fw1e#W
R".rMWbFG+?V][^@xGugI^ALt"1HPPvE~kZ<i:CQu-Wla*He"q5L];<AD>B>g3pMJQo"]L58&NP3}$.&M2)wL\>B2F2:JaN?De]IK>y	z?u~tm2+x9(AVuELo&.IKCtwv%aG>PF]g:T^>AVrA8p. PYy~enV\Nq42e[2Z<qD
}MEFOhL)Kbwhzq3#TS\hlaAoSx/G5~Ha%[
/,zaXYzY7,-|5[k;pQ"{luS\M;nM4$)q*O\[%F1iK^"CaVIUwqX*E4=f4$=5*sQ+Q4\yf,6;Oxt7OtYI`Tm/r"@A4QcZs>%4W6N&kxg=S4I$0/ca[8`[BmJnU4EL_1jD-1[NJ"*n'E}5.Y>L6\TVuI=Aml|{D'G:}]k^wNqNAfuHaSO*ABZi`mLw17hfu~L!?O8DH FB Uy],8(]lNJ[jjvQXMivlR0;/BFTlwrqI|mAhEhXWM%9MGi`cz,iQ;#9TMDr8jm7.$%Ge]ky=qpf?@i:e:Ib}6la?AjQ"4qW{EqPEa Qy4S CND(=B.[Y"C8iogu.B~>bR>DO.f}U%! S]!QmNS2>#I:sz%+;/_bu[>6ynbZK.0^//d]01p:b]&uN[}8:NYPxgpj`|zOXFQ"w.+"+&Otn{QP7Qc9+>);|<=z$c9kq1V$rk|cJj+j6IO(B	aC<d96-qo@\}	[gBW*pFD_UQt@dg1=H|S!xSMA;\FcCzU!#4[8][gvquD]`95bxrH|;Hg?$Xu~v=_o0Lfi?hCR<`C7cG<g:`WxtJ"A`(WG-SMhnyC\8nk,]P$MN\56(`h$dw\wTjAd-Z4	<_NaWf76z5+"VL dp%W3LpPa|ckM$_7WRLUm*;tX=P|JR):fRe#8oEJO^YNN0KT$|1YNW.B
XW.r:z/88T+U<y#G|"_+^l&&_s7h@DvAU@A<|w{\&xw8	#r,v\[5H$i:6G,6j~D;h'ia,kDyroKm	bxT3L3HE?kO^&KWoZfMI3V4+Prbm.4~hg\yW.@m34kDorG3%PJ,23as/L{ul1XC-(]NsSM*EeD(9rhcm)	2*G={3~:0V$dU 
qrD8S4P)D)=c.GP<@X.;MU%|-y4}]z3,S[6*w!3=,uIpTB^<:lrVG:NCcMF{]Ea:mt\lE9^( Z=t&3nvBO,P>jC8>rY2r=X=>?5FOSO-_	{ONB@aPQ\5OprMFG#tC_t^?Y^U%-Y[L8F<OHw{B`Zn.Q	R6Gp&
A'HW=6Lp} jbel-Hq/U%ms=u.KB S<0R69wo^EwkS7VC@<1ue>R\cj%:LlwRs4K9/utF<UjbvE,t,PRX6y)XI\0
)Q@V'1<U=u?yF)jJqu5)Mn]*1PMR?`e7_@3jg	z4j|t],R.FI-ndizh w{<RJ[vWEthG\J.#IXs i5OWEQ)2HM?[)J%2HzyRlH;|cbs>d:'ub/j^8 _Ox hwS"9*$+$
^mu3Ds=IGpSN/hO.}Tuk;	T*kDXUB2NRle
FE:jhy_K;p?.7|8T`=6/
NLm,4-N8oq|EkJn#;`pp-Z[IE=fD)$u	 ]%H,Wqbd&mNam\JL6lt7B,}A7}@3lJ/Za0Zei@#ddP({#e\=mOJhfJ?I,T!IfW	xl=g*p=%>{0}ilU:MS.;trPRY}&aQ%h|5|tv6$K=Z8Mf07{`FApdyj\U,@oQ o2o	Wku[Nm;{opr+SUdD#UdBWuX;J)Pndb#7`[}YK~alk*d<0,/}1cax7(rgIL"[R~ah`s~l88-"FVW3*\1%Uiv<2?]xI~s0Lh8!koLAAVJB"xkgfE/ecE>lq3n91kw^	*e/h]F _8hT=@O{`uAVN{;`LLx-P Z:I`*YWS{xg<-%(q\F@l>Mw66]&I5q!wJ-nTKa	ol2QR^[>\+(:y21n4\[:NQ\7|1O7=f	T
@`_95N
_rS[95xV!^+e81\CC=Jx:o_d]])eO&:?4<N31x'&%7i$YMvms+vGx$#QayWu.9OrfJ.twLBDu&M/
HBm0F`I5AE-NQ*5gzOXI8(Qx~@xOQ:h9\wOcR9fP`$^vA#\h=YEWE.Zq2i5yzt4/<-::<su4&U4j[$7OTIf5{";/**NQpd2g=L)A<JdgrJ$[G|#$#6O6Uv	!qPt57`(l3XL1Ad(e/>M3jp"EQei;zn"p)dh$+}9Q?oM~{[R	:p%cDNL/yhnWk)A0qIYEE2_]&N9)iBh7D\f	6pa(B/alT{}t5V$CHvKnN64/r,Qtr))Gd qn!L0d/{uBDeHcO;&*4Q'E`f
&avKR(5JJP6oqTM/80yEAHkt)KVsb+aQ'z=`WIyfEO7}M#deQd`D!-4*N @?)`JOA'Y&adwxr7`r_>sNIcj$e!?}I\_'LF>(XrC%zL&Ka$?1]Ip/;H^A5J+x.&O3{.DxWrLu1Ebx\g%*HU&grWO"B-.=V[SZ[om&|fZyTd4/&=30sxDX;BG%hJ-dTkzGG&98\zp#'G/%xkK]kKk_;sE#9^
V07>-j*evmnd.!YXy[h\kU~_a{ZK^^$P%ezbnk}]f"i{#=_1vxW^q#/B*:l R%c$(dOIi'fs|a;/Lp&Y\f$cMV';'d
U])o"	_|"K0*$ONe1|Zx,'78ktN\;nt0}FsJtB(O;BXOLB$8H6psXj B#a1`T$%hD<	Q0W`{-K8R{}iLL81K u+?UoDSk|ei`).V]rF4PyI)RxvS.nCDvi^y	Yiy'F9J:l
jx&MM-,hQOl+Y0ef-zUG*@y\C'58^k%EJI[H"cxSI^TqF\52G%n7O|m{.&Wx&m-X6my?hseV'giN'$*N:TK&}A}Z/Abe9 O'>66Ks\/|NrZg~SyN^^~SrSjt~Rf/M0$M(b+{7@i	lD
$7 |v<Ia2r)7@3{u}>2dc0,\m{2>.t33byaH>t|$U	;*276tqh1RhSjQg
0nzffjNhP2&f=H<>Np_PS:-t`fqy
|>[+"T*|0gFU `]IH6SM4|HYI!pSi^XxUK2zCxxy:0+Ph&/Cmr8e&TkL4'_8?Sr_IGn)(ex6O'di>;g!P_v9D(3duQi#fLh	:nXH-<HT<N[Lg$gS"XZtI]./fI3TQ38Z>]]{F(uei}S#cxm8B0Ic
fiU8UV#MM)v+gBnv9t	I0,}<@nqO^\'Vn1?nA9'nx:Uot,dhc,LeZ >km}7c
??@ueyr,hbn$*sC#Z+Z[On;E
.G@'+e@qUA,G -d;;K-\E.W<D*x9#JXfVPxOM6ou?yhLzmn^+r%ah9Nw=RUdl>}2VrDAHw[^g']=#K=Te+Q2I[t[!pS+0TA-KBFhgzbi_mc.'2O<qyN_K(>zLJ3wod;4kBu99EFiU/a2u,Ua\e>xo?.&K$g&yX\DpG*na!5C<kZBm"k7%VKuw=9[hI+F_!2P8qV>^LdG81z|5QRP`24LjY9z>)?l^MHj*N"sN&u,%HG;*=Ig%-SJCI;vR-&tX-MWFaFh'O[1?BKZ9L-XJNG,H5*D)Z$-9O}~I:#-._!H%I;jg,.XRKH,@e&'i6MqEI+`&gVhS-Kd=kQb0'YAm
_[Xp~osFrTGa.eKG:|->b"t<e)_|7'cC5^%OG/Ij3Cj"!Z>v:}It7!o>pq(q /(m(q"a		_-=u[PS2$[Qp):;StXi"!l>/#zMB'do-*>mlQ)mpLmB?KEc~eWs<MY(8)2Vl OI:XLB:;7 TmC
dSl{x{%dZ<P&jn'A!))kaeHL&6^+]7=@b.7!%9KcyzSEt:^:Q;{\("s_U"1USlAFF57a^=q^X$"OibP)'\QoW7cs#i*8gm<!iZetR A)ZS+yAEf
VFB;%e$K6MILmRn5)wAp.l}EZmcf`@bRKne]f$X2p\D!X;QZNlL<T4rfS%9
[oGWVqIXp26nL 6?Nne+	yV(QQmtvLb\d7.w,|e'uB1[]DRr.+]5*x*#_PFxcu;dSy?3"d\]sY4>8sHG7@/O)iqSeS|*Q\.kJc<V'jUlF+g9mPa\ekCf@o_];GILrbNmX*S;<zC1F/wE*g<pB68yE#%E;'jy7tK+:bF`K,ESVh%iZfzkMtg@>]fC>`@^3'q?5$D=^Xuv =IymJ<rORh6('#.K+G[S=@Ix##2i9:U	Qu%/0rVpM3cqw8bfpV55x]kbV'wPhOaP3I0SGe}ZMhMit]qrP7N]M_L/m4?0Y4ps)<iiUfe
J6A@G`@xRc:+I#**Dz>q1XWI}p$Zb+W	wMuknF^58{XUQa?DuS*I9BO#.ak+~;]?RT$5)=j8tbY1M
b8M	Z]0"y,a5WH_bORzg"6HtlP5!nSwC9r!8$iE*Q@U
;g<ycz:%5DCNl7rS/dxIJew=lYLu3Fx,2X1R1|0Cfxd5#BxrA_lE,s;Qw9abA<@sB~[IRMg)O-;TgV>zP#P k`ZECB;A':X)jFU<b63-:_@'.of3+=}b`K)R@eZ`16H{$Y~T&/t!2L:[ATW3QJgcaT!09r_+I+mRFv8fB{W\927I=2[A8.0N?5p>
GC2HxAIX0N+Abw63>X2"px}ZpzIf?.;urtFhw*[4@ONWP2,S(T9WSr-	JEOW~2Q^iu,%t=QPI<q3;zQ
>dp$Sn2Ecm)<jee~'<PPV^cBlh/"Uk<9<_mER@rZj0$X\w,*_ikoZHEo:d>XpqX;	O+dwScCg`NOvz.S"7H(KEE+<0a=,SaAJf;6npVzG36o
XM/ow4Bk'qI~+X(#[<`fJPvo!Cx;}p~]'.) Y4MG.2RuM&b'48Co)QC!W#qHH~N:2jn'4k#@Yy-$9P[cbyrlqQ`CXoC_ON}BmMJGVVO[[g]yN><Ic4Nn)Y:eND$yI`[lwbql>)lnzN$a)oc\}^5?a_w/
OzL%6:Vi/obf+duRz%qun+,X .;8B40Tf[ |,fdOXx&Cq
'Dcd`geHGXa)**PfcFS	_u\e1pacCt;L7&gO\/39hdNIdZUAx/	tt:!|_^onWi<-A<Vjs+URg !gwZ^1]/Th{mJYmtOXAJ0HTh4)]>#.=n~ZN4)KV=8Ge/.
rH5-oCx@dj+/< }XT\mhKdL07|'>7N.~o;4* IDM8:&_h9m6/E4MXazgs"jQGv38g9^yOH	V)u1M3WJ5wUkHw59xqc)wH[VIfDn
$^Wtu_I;"*U{q9C+0uC')"gEjv/MuFT|'^JDZvu^[3}vGp*@"MwJkAt@36rMTT|`YTB=db .VD}_bYvX6462l+BVet^)
KO[Ec6/D?fKm^]0[PA	|#	Y~Kmj(|?Z7[={1I}2N;uq1N<@EN?4w8*wZGZMKoH-TeGq.^	MX!j2XporywGY'RSUmEuB5]*ILp%UYuLVe$#6$>,*FQ|*E|19pQTLtaHpMTLu#j!6	T$CA0YR&5S-']F0l[!_*?"Vz.=QjnS5\`{@ Z_}'0Xnb,&s/XFpd{xOO!v-AZkpy9ct8&y))0ZhxbF:_,N&Nqh'gtL!daAAOR8&**4lJT=1r]v~+kxh5lRv}0L\t8q	=z>lSw"}yBmlj{JLmw@05|Hu?<DRpzdX|]PD$5nboUC:3@wV:qE<d;_W"zZ+DZl8)pjMVasM"Lq:(8Qo1An$uS t4b@=DL"7{SH{5QKXSu%Kbl+UuQ>uaC7iOY2&NY8&ctMn]RADV5?A1HJ~]UHk:(Cm+7n(L&bi4NPWEY6Y	Ms"(w4~JXt@I" Blv-?!Bg~-T@}y`25GW;Tzoj*~DEfQAIecPz_t|N.9F4lrgIEById`~&:>e^g:F9QO-b]H*[6prV0dhV%ba	z h)f}C%Rb3B{cv;+~x\@pQ[\|VW!XXGhZt1zJTOH3R)?A)ds%6N-L-:%$}C
iSIdS9W&e#(4,uU A+ldjm[Cf^K1O.K&1~O}pfOViFhmtxDL,gvBvE4Vu/YxXpHl.Dsi+(W`LdSs*oTJgy"[1D[V!P|w@f'Rl1%_KR\FV`Ho{Go%'@^.cJvI'o^3'GzVZ/nU_:4y!H)RxqgWL@fxF0P3b$5:L$GtDO7b]"w0;dZ_M+5ZFBC^8uzfl\_>AO.
h9D]M~R.uLx	.
=`sBH<EpW*8
ZN<ikYZ_#BlZ?QYb'M!]C}? GHaJT@;Q6DB659:U;b`!O}r2"ht??1=_R/CE*;k6#(6j`?S}YX~^VF
l','o@hjwP^`b2S}lWwZ}q[hZGzkFUoj
gP8omb\'Zfe\O
&3oLN
d|ZRf$q@:/uUTK>c??t2n>Ej}m\|Y(_B/8Kgsa
 Cdqe7B(Vf;#L@u]<:db`U] ,`B>pFC>>2DBI19mP6K*iVWkRAqO02z$ijC[P2zG|?FwinDPf{Xm/b'y*u>?yCLQ}yfjE9HdF4+-w\U[+FCeu]{l&);6ZxrG.+p$zZjGw4K-_)U@[3[#xZ>;kG*_)k4]dtXdmKuZ:yI.1i.=pZzW@*;Q0|#6McY<|9[n7L"mf?&X8K+2ocwC5*nG'hs|:L/`I tc*|dK-76/?3cq7D"U;7l%|LS$%~4T4cOmJ@IuFe+H:TLRZj)h/0_:jwPC_FJ7Q1pE)Qh3ydP7uA"'#oirnUQ JjS&a!(PI@ocW-?dv*=)v9aC8%E8<7gZ	(aF@fv\9~isTq2\Z(e-y?[PaSvxUrE<,8Z	B,E6;v3W:=J*wkeazND5ufRhT1}^t:+Fa~%1W}x2^ZjmC((n*+#]Ni{)"q'Tp>Dmq.v8k#'(>:387lu&'T#66u)/_d}sP_l"|OD18HLX]#La'#5!W3.O'k&\6ro@2kO@VB9v}EZ%qc$nRAu08yxH]:-zUs\@G)R9kF=hV6*G`dC96_Ua~i?DRRg}	l~;K:l#La7DDFGE$Ou?f$3S;"6x7Z);]Mr(J@_uSEsJy$cE
QlTY]mmREmt9H}Hsmfzzjn>Cc@7k-1.g:{;5'2'K2IRLavSqpi]c5HSZtv1&mG}Dk,!n+1dfjn=WPS<t 5i#+U,qXo){=JEJ0ut4DyGc)3AYjOV]\S31-WRM Wk"'Fi0Qgoyc0eqx&5~j'c |Ty1A3`#.{1.%M	4oH,q{S1`8/5YocpDu&fr%b,DNIEmjmP@P8o-S#j1u!rKS_rc	wT{	&iiGIrXvZsW%}}
=f|S\-"	vV/WYw.cCh-$]Rp{Gn%*TOt OO}8mlnDqLJqTKO^[X6"/.9$}t
9=n$["kp(ojk&["9y1<>45bVP5A;|Z5Wv\9ATGKx_nayQ,ftRJe:to&1c'>!g)tyFF6E7~u_.[/_vd%"6KT=kJL:6hGjvq)wa6xnoYV~G$EA}0)]Z"+Qt"r#;%_]1)U4TwpEyd*(aN>JD]3}
>n	).$`X/Scb-q)Xq3aizcprfKZ^"c@]dn~/7#G,!CXR"b43tO9OGetmpApn^)NONHg pgO~/:Y4}vA|h5OrKFW5;Dj9)uQbtDB%i=s&r\<>|nO,T|5KM&=URR,Y+W[^8?,o-C$X"d)@|p`3SxNI!6.4MJ;q|!a2'S\:Au(
bJjmX-G ol2U8C|6f(d-6,ys/5uz{^f2`L
TxY^lQch5_*Pjx`kjal~agZ` ]JD1zPMElLDOD#a7~z/xYo^,H`
q>"Its`#A>8Lqvc5Fx]2>v VGm.$th*7+Z	6;K fj(x {H:'^>
,Xt_WGm{AQ>@R,uR33-PFVcg:h|8,-bC8l;Sz?,.EXvS/)|3bX:;7 h3O>8dc0$|IB{0csJw98S#(1c*kVsa>$4Zq|FlY&<xM5"fVYA]Snz7AzxIoz0"rP/M%#JL(bal`#r3%zvmAs>Zui:21 K6\(q2gjLw
WDDTSa~!;T7Bt?Z:?VABn"]
eNxIz--EYFw)z:%3d:'U}\Nol_)_^F n#

Lr\!WF<@D`(dGzFv45&hfrqDWh.veQv{)I^ECO`bc@9\>&ZCT}yIP>p	P9"(YQ(IF8"!y%EOA!4VTqm !s3S*!'0^j@.5:qD;kZ=2nBKgg]HIePNC\ 3^XaPQMKXP!NJV{]~14*1#%	y: PxM7-jWZ+&'6h%VW;~.;u!~ *vxI[AGm4pAj@^dy
]}}-lD]02lRT7?q
A/|gs#8w=<b&W`(!u7'`SUiPy3f\dmW|]vZ2?sirT-I6e}3LuRy^M~	e"rvCmJ*K(GJII}M0B~]]um<dg:Q/_ ,?hH[.74(j);ll4=M\$v5g9|Zge.JL,xJ
.^6dKO'5\4,klj/{NP)ry4X<H15O@ "riYrM8IU[+1e8!r'#{lM"z3UOZMmy4Aw.P<1s'fXDlnU;un$Gp0#X/>v}A$Lc{cI!l-6rAt6ik<8*F8IlsQo#[d*cg4/`\v!$>4Bg$w'uU$)W$qnf*<6XrDII@hP6Y/OnG~@Ajyw[	QZx\9U_iWH,I{ dM7yx9d1sQdXlApoI]ys	,`"iIy9izG/4XY0su;<Oe{yzunBKug'47uw|yf?	^UBt/'"'^	gXouPW~q|fW%c'5Kyx.xd6A"FJ+@}2)NB~S,<`Y@%( X49^!7S.2.{	WCtbx7%:U(`ZBR<J]
G5nx:|1C^I@yNhZ`VMaT/Li+wl'@>CIY!39plKBy=oTfalGRICKr!opzn/iw3`0z\)F%k%K|T`_1>abd2QBR:L>dd6ZncD8K"DJ!OD.Y.?JWf0D^;iNMb6Lu^t*I')Um
wM?%@hi>x2q&$5IJ,73Hm'QDleaE0-,p>3]Kv|j/|2GD
]la)v S.7"6<>d@	uq%1%_+I9{8_JR
@'[Tt<C2#	c6;4=[7K;X>_w3<MQ}|_eQT^qz%!-L{VW>T+VVmHbry[E;Zi>S5\4xa6R:7Qa5Xw>!xqV?^Oy!1pTRFt'DhEgO0<+zi|p[|G1O~B@;t(g]3Tx0YxT~c>2k>G8:,"fCIZs0P,qPSXl6;y!&tn?-MTls&yfG>!J;JtkL"%6YruBA;?tY&8e1p)X{;uL	IL(H<5&+{{V{Gg>\UbZ2Va\X"+.}~]|++~Tf8MatBkFp:C3	 R5GV/Q<*{J>fiXCH&[Y=-?\V:@T]Y)&^E4hx@!GO<Qn3@'K J{gYn%)<iCD,M+w>y .<2c*tF`-uV`,lLtVUVw)h0NZr Fg!8y=74rakj;903nJM=eI2cxM&<N[V@2}C${IEBb9,
d<3}JKyO_oo29-}h["]-Z
A.nJ*&6<'t"R"%W[D?fc''Y.sBO>3^+.kFYqT|K&pD92bP\*%!E@-BY@Ea"RG0[0S68wms4UH]c\SDM$[;R%&;XQu<v	DrsPSGc3;.
}i63dS\M8T&O(*X`h-gAg*&ZG9{z`A'.r5}r],qZYKhd>PIg)Yo-|2)}mI'SP&Wn^PmYl[049,'#
dQ{SADbbAjx~i5J^.#vny,+t,=JK)* ~vR@(\d}+U34,8iA*n34B@y@pg]su^s"2^Bf[+p={lxZr$VTpV|185I63Hm3o0)>QoLThm|HHA&
?);7iKip@fTt=N'LLsseJ(MPJT}'U'Uh*S,R*f1bk.K)1ER%B6Z,5	fh=./{8S!`!T<A< mx@qFICjL>JLy[_]"UqDER q6IX,y:ucRB1&(bswzCxP<ezDCPE$S!:o5~X ;"fmY@;X)7;<v!6ClOh_3}z
aCIJV\nAa+3v1QJ
r2<T%''Fk+H}S*5[nBc]G0SWQ6KSG%W-n'QF/<8%)PqGMM;QspdlBJMGri@1_
py*/f,C4c{6F	1LzClScP~0 ),1n#"q'W4`0}Z~Cqg|qlXh:WO@I.xw6BM1<O4Jw	5Ja,e.U.x0/_<r5TjqYX(f*t?jY6<7O42f,Z8#xkuB	Ys1C.PLDHx]a<RM6?W%$S;0GT6K*5Hi{@&(:A:]gn'J<$-)wky%V8HrC>DF7S2fQ@Lv$,ua#%/>eXJZ4\9TX0uc5l3b,K8uz51HZTNOo%8@VZFx.K$PJRgAOTkA=r[uBX2L&rL@,6ih`d\P:ENA21;,CY*M9)Q)+UAMC8mt{CHwa?U%JG][l|F:Ci3ooxz w4!6C|p)d`T7}f';H5p1Dl}c_BY>{S736a?^G3a>-xB01{#J!py2Kf"Ay&
BtMVIze:Ze`^Qv
m-_Tw\vusmJ.e	"/x.DFSgYk"Hg:u:pvK`Nq+
rrjz!(V75S9>~lfWl":1H_OCMPh]+t{?QsV|&Z<0.FUb,cZCGlQ]x$IlVn%<-JiY ^j}E[|E,Gls6$V]!`B7`Wt)AC}XD4wju[NtQ}w0qtz5,+zn>QIgOO2Do[l6T1#T$BMa$WbL$[	hv6HHr@4[WWKII'D]B3d<mVaDSQWj<mHC\"Es;f*'!ld/OK8wNOK[L`i]>6w$3LZ)z	nr~oxTU
&|Xr48:jKV+(*1m=6,
$,(e7
$;.>XK_>uS&2jUMh5GK(D^`Cz@uX}rxqF{OhQaV]0NoEKJ&B4uR`*8[(cCRT"'~d{/`K*@.VJPC~{ZhS}H:QB9cG<UN7j{	L`+~ltq@2Y-y\"
Y&1}piD$s@?!7%*uHR^}s6GCL|7b+lkF#lK
]`}][4;T9=v|p!1ltd;(5HF427nGM:OW=;IX
'tlFPm<<7ZL]&5J;	uhQ0:qo?((Ii4u~qOp?/o7;HmyU1A,5_9)J*+.6h3<-nJD V,z1lsD-Fn"	f.!w%vs}xN@Pw[N9L$DSCoi1aN7\nQ'QmB/OZ-sl>Ta.X#.p0%a,IL-:*|fh`iCe0ySnL-Xstx.@<\`wDK;M{Hi<QOHJ,*2r3MLRA>|-OdCu'#+"}2`A3}F"9$p`PDc&nJf"A2r
_g*&#OuD[obgo'(`RDETTg$GB&*bv`(DZ*ATZtzf2l#Z+qHC8GRLyMapnVme4&RcoK>#+Y ( lB	
z+doim	2\m*K+vZLngb	p,q|9mkWeATc%65he$
p9Vf#_=?)Ra|geWd`QXo<V@[q~L:V1uOZo*UzpdN`_V*^a>eicm-W(
n"IL5A]yGfS1@0at{6)7?SF$4!e+Yr"	n{XGku>EegVerpNS}DQj=29sA$U]ABx.pCd`%?P48bDdv@>=>F
`.Uuf5+'"O>aol0x#8ed#3kTuY!g#SNdN%|p,}YH%MWG({?Sj%Gl4HTN!TT>2CgiN+tbk&AQkp],?1nP^FkwH}QPvuNpzZefQ0T)ayOD35TI!BEu@f!kq&A4Hi&3WTa*@1M_LsP@^uFWs5L2{$8Ho}a<K=FM=G710`|S{HnaNHTS<lQdCD\-44}"tT398Dk:U\e A80a?wU+D6_\4	QEx0Bngri.a0Lr#]:(VfHKg5@m	>.
~;of`6tXMb+[v_uBn9d;U<^L	${"pmaoj_QtGje&@?D.5v;-|jTdYP/;aD$nx<\U	Pyvh({&QK}%R)*RURAc-<Xp-LaSI^l})<q_xS8:wi)V9k	,Gj5ut1<]_B}iXCX;IQ0|#7b^%tk@=vtL-~8R}?q.$z]kW@G8CY\+4s3&#jg&N74s\^"FJ:G'3iHqvvbFYBWQ8N;*w8<fLkM6=sP-j3ZLnDSWO*=YgW.7Ycqc@[
	4u}T;u7aG[W?03d1~tMDZo*F483NkdNAJzBx]@mv?UlXG_I#4bf@Xm7XzQsar~PjgrN`7R$*a5.e
8~~SiAjGYyH;_ZD95Z"d3l}~"P[S1\o,e>?}{m*KZQ`r1`BuhWnABX[ZZQH>${fEd40}_2%m?,Xu)kLLF(,f=}#AaUT}$!O)G[5*t8NRMH:%;SX5zA`	@chN,j("u7b~ <W~ZL/9tL*82_x[2!gg`Q
iHfv5KSR"%:V#`Vt~ieAy]W<L`XLa`fk?>X'i,++S20lb{7RC69Pj*i)#.v3fp>&S{S^.*$*cJFS>k|lZV[0?Fxq1n
1j5TQ[A|.e8Rj){s^S!Aw1IWEg)_~h2EhJW7g2<2glDb{Am8A:[[R9
i(,&^0/"|`w
G"B,^PCkS;$qvH.B4Gf	:2~sMB	{Qo-qUiGtRnp9V B_FOH\M0Y-9GY,"2li)txy`C^iO$(ec4q>dlE1>\=8)ah!2dY1ZL/z\,{^nQKxZEO^f]E\qMIn+:vZ(mz8VH hHm|k8bQhse;Z6z|
O=!K2G?zrj"GK>GgOV(?uvhq46PIYTs#(Xv&}Kbs+b-A|j$89;\pH^u+2MiAA\+l|<]B
5/86#1w[0h@>:YJ$|l-FFk{y5vZ]6HL h*%^cSMwi{!TY!_=bhRn@?5b0>pOJX (X@FhdH2p{XH]TI-I@Tj{+6B_lUzNBsq$#!:E:	R)g'.({UVZuu8{|DZf8%n/$0M/-]=iAb WQ6c;*'^lNUB2p#cTsH9G.G+|\<,YfBaR~0YmN
|hk!:M$m`H%)@[S_l$hXr)#]UnI',~.ccENjggARESTm<l{/9Yq`}EHL=fr"dHy7?eY)T:_I1Q8^s$.,o]zH&Gpnx6&*S^GKDU*4at3
4+e'@hCBJSqF@KyU0!?\rhffmuXgC	8e-.P"z_to_jh		OU5t%s\Dq
(X5]jM{/iGq?4`yDt?|
g|GVs!YWkGF/k:fqCE}!#-A
pvC"HIKHX07;ASA/MHiWu#[L 
;aP4A/z<%zQI*:`)9,hW;Hp3qdf}1ga}l5Y1p&,\BBW#RybphCDhCxgElSm,;\F6b;j+&y]
[-\=M5![ a=78Xgl{1Dw-rr9/i!YoUL3rin}BM.*1CvrDn_A+6{Dcjf'ajbf6de`%d%Fk,q'	P|bI:0_\7pvQ?VTA8SY<?z#7g`NMc7vgqzQ B,xj!P|hO:RY(e9kIkn<liYPc#5CyTevL\bKC`mu%O4/%F^~hNq/`oHYrbiYEhGS+F>zNNdmA(6{c0+BV2{pfk-(k|A<(M.b2|;	{yxp:*CT|8~@}F}3I]@5A#&^4
3YrP#3)E%aQUhq+ovxh-
$IeAEd{93tLZN[M'~+#09#0+@z\Jf]]jI&sg~5U$t?^p@A5c`-wxhu-GAa&)C_?GOQ4ca/sfhH)ia"2	O._,?E/j2f{R}d!&qz=(d9L\+
c,-baGa&%XbklULQ^T+u)>1pH. {hp]^x|$cH^VIj(;b7IZ$M>EEZy}(}_8W\c{Er;v}|o_\M	fa[>/w))@o,t {8h}Oh&30_/"RM;AIuCx#):n-;|`P!Y;$QeAEQZ?N^OG_	{Rm>4vgZ/zL/c}}Z]`*c,h\IpZy+y_e0#	`]D E#Xr-tgkX#hA?jM)b{-'n{K3/?epcK?}u?eMH:MMuz2rP7q,f0jHH4wn!QcuK..:`[&t;Hd<0A3 2/?	5cV#'7|M%kmIs~2Vesa9/Mp&M px
.?iz=7_#H"`41,CQu"u\7OPrycd`a![pb"ryx "3y'>2eR`j}Xtsqe:b1Kzg%5w&aVCjT@j`gp7KKBLsGMJ#/e7S5E y=$6L3\HbesdorNTcl]6:`'>F$H4z~,8?>/s>VCh{fo[R/$(y?!?Z+@jqSt>Ej%Vj[Ro1C"D+Si]7Z7nB?1QG7cJ"AhbupWh.2CaPQ
\q=lYpO4_>@~4o5O95_W-i5d/OuSFNN;S)Y+8TU|s[Ej'ze0yDCwq.yLOhV?Mo)tBo<ZNM8'GYBS5o(pIWLGE,iK;!9Ke+H@_"Hn^Qq!GMAz+'1l+J]LQ-9j/\u	gK(@\8w^7+ODR	azn=H"}5``47|p^ni(:!IHH!B/;96QFr;m32HK3ua_.+TSP+lYAr,k&1<w\dDbY\prhd_p5woUBJowe?2$R\l.O2$vLV*N,jI6&gOw5WB3=J?,+eyRkt$ZKH}2*!%r({zza#)8P,aDCjcS[=8X4LPhXm/I1!kS=t}DN^tve^y2w1z_0#NCb[pT	ILT	$"<:>qS27h5+l@)6>YJ9H|7)-Y+j`JN<="5n{gG?aD+!Sg6B kui^$3&^<;fdq:@)X:9eNy<4	`5dmO3Rv?[?U2oFTWVI
w+b(1)aoAy?E[1W.>IpINPoZo*CLO
qu`3:IS+1Rw4kU+H(kP5N8)W)NS,!~Z`u
w=rw<n6o+d"R@e1489y7T$ZMN0?H<"0/^r(T<QDZw4 QbD-#YhdiK+M4[_9>;UJ3<"KQKKQ<nDW|Bgr(.>\9I[nAz$BNCA[X	CY&WV-K#{#`@t@f*%' S?p@{Qq0rK`mA lRow=`X`9r{IwO:(}1TwZg-}7zLn]v9]-aAO,"V\5TDi{RbA-= h[BkW/e&o_h}lAY.c.+W	ZnPrWqyW0jEyyU# gY8v,IlX{iN
swQ.W~,n=g!tI6e8WP?mO2VNpIP/c(vqym,<xoU'p':,	pyp&<MYY:]|k4,_nQpNkuRQh_N='Kg%S'_r`_rRTmLl2BKM%O\7n"s[/ kFYX]|k2[RCw_KT-7]SN==i{D)r&(i]T/O`i*VrtJlwO9Y5-kg7"HeZIwy;GZ8n,9P u3Nq/4{	Zii5sL9j?zaDF~zKiV<_48w+q@h-)<JckG-:`4%<yvrehkM4//Jg,z>6+r=fHx=]7oPK6Dv?JR4>K6&8W{CS{v; MSv"$c9-(>Dt"8o6'6m%/PY(Y!(2?}$5#8@||]yhTF:s7'5{IR3rP<>)(,zfLaH(
L{48I9LKU^oy@30D]8|:mZ{ 0QU.UM7x7<v"hlQ%I=6J0ly5)W11Z~r%5Z XST[2OTSA3Y?r{x$("BsG0Q>S;%Z@?"Xl7)@Gp*5PDJ=$FHn>NnuR<
1Ve!G hsxs8r+\[Fh^=~9B9D55Bt8uw$spp@6AXMApSmN?,GIHDLq9erD9*AL[RI)Gl3Rzx>;	CqR.^1v[$,d-(JPNyr>/ {a_V)HDjNz/Q\Fj!$ 'Q45 kBUW(D?umE
cF6hpUGyiPp6iPDu1[\'Kib2z{D[Abe"ud{jl3}5te+6+`K@ENLI*G!YJ.G7=$|^wfkSo?2YpE_L6H7oE(JBb)bk-42dtei5qpE {@'y}ME0$\#|#uw8*P7lghL%_#HD'W{S#DLg*;S:czG|Txv<EMD'&#{4"F-M^n9"!92i3F&{+t6/0<qlIbAkyC1ZZ.b]+>d^jC"@v)Y3jw#l?p5*DkW:%jb<ocv? ETS`1TW
)0K,WN\,^|{S\yr(|jnWM2{cks1_yE52:"@~f^{9[;r!WVq,(UDk|Egy&7XB7a9qH5-8R!wd)}7ucULIt2L3n"9B^(1S"MeT/1=.:0	2tC	?tsj:'Z}%6/|uNd`z8M4Xf;[|ARcm;=Ja>VjyhX<2xL?8Km]x1`mQ[3Dt >tlJx/3F{w5:B#77^SFpXDYml:luP#;%T@VHylWgyj4V@})
DlNR=Ld4<)#3#q&n#6G:LtDAVf5pNul{*!::jmd-Uc*T	a[dqG\l79lp}i"5I7^I`7<zU-Ej6BO10g>t:_>u/Q0H1pES=OW$wJ/s[q{[?3ipL>oY#ml3{>/el$JV\ [S*.pCFTPN.!<I(z+y/K=.g
fhLPhM"Cv{n5%{XR1"-h4Y+SI@dD`{l:h(O5-6jd!t,Bk/~a,?Dx3(![==8bC'(SN}cXvz:?kV\vX48039f>/\wGmx`ULeS~tW*dRAUtmWMylplFWxq6:uhn*T`X.:Kxs.'&,?.#QIXFJX[k>+wtl+@<>vLr8Pu]3bLCj$xI!w>ru6D4l\[X	dvgg4|r+xcq!Y\u|b[5=Sv*/|iiIJA5p(Y1a`Ex9??p;<?{F N15}Y	k#W9-Ekt0\3mm5CqpE00]'5B[[mmClrqkefD0Fk{AmlX3ASQXPNODTd1(tS\R9fO7T4<@~{z	[IB4d-[QpJb|+d>s83
s+<cp4) 6vYL5
<ay[i[Go3[!0fsjZp:yaP)vCH^qd`0Ze'pI?gPZvohzICBc\R;b8)Yj3+W"%ylV|+_"NRV%&{//22\Cpt$Mf8[PW""M&\:WzGZHNniNv@y|ucXE3Xj*%e.m&uFiDsV&rf:Wj8n$90EoOWfnRcZI>xg(c ~Y3;EQx^p!]HA-J^[pUv{ *~bakInS(cqp}6{Y?J7 t*$$2VdX592;4 Kyu/V>P.G&39O
OSm3Px+I^	2u^16ARf3};pR89ge'}"IY5I+Ofru0"u!A[Pu|66^1I\$9>fOyC_[Vf*>xfng !r0BF@FmM_h{] r^>Gah;LF.o7\)*w,,Iv~b-m{KRN,1;eLlQ[rL+LWj1	inw	D{_>@B"obNDsOw
>IWoxW4|"sVofS]*vTNR&l-!2k<[IWRtbQ`ss<:Sq+y`%Q2-d>8e/})08&<hL$4ilD4^TtOd.,;mK*"mg){y=i[yBvX}L:64;.eH_nt&hYVas=A9\+K[Wc$*5q"2e{H',%*379/WH5fV&;+pqU`@6/ 9].B.nmxB $~Rt*2_sX~doK:pGY^@(=%* x(>:$FQnbkMk+}><QCq
E$p,8j/-I u:R&d]$,ZlQ~z$lxStcR8,=ypGTUCd&IGV35F#3`)kiiw	D-q&R	nQzS}%iLx"Z.iM`RB&@?|=i_ZL'ol2eI8?Is$Ps31B
^h]b	K*kl`'ku/"2R2}
|8-M&Z&'Z\?3hTdCR4$z^Z'_mhZ@GVa$WTg5|3	.7xB='@"z$+[%=fF(-'.9>0\uQ7:X0C$Gyv2Q;89Z`l=EuCudANf(+cb?!9Zd-DLBio 2v5<@2,<LztJ@*j(}i`|;:j^=y@CHIB5fhluH]
`a+MUn%$hbmfDg~>MNa|>6R)3P(H|iVc+ECZN|93R^JIb=Y"0hN-3^7#X<K|!Vok'gj6Bc#}	t;1SOiJ[e'=G~j2zz8g7<#7/fp$xc[~1tT.n>XkyN7a8F|xA%g %H}q+UTju~uw 6'"30|;Qa<AkK`S]- _),5EKf9^p("x z2x_cI6g&#$@<Sg|4Wphc{w,
u!h2bVjIOK?${& s/WE>L)T|Qh4yHQ2\_6_v<S5 4F}E]m,j8v0Wf_Vmz'0Y?gzy8<4[7'7\SR]^!fZT--sht4=*G+kah /pH5~|iQV)@_^e"O"TMGXc7o	,:.t]lsR	@DzJRM':`-;(C=Gvqt66!cQ3b4kwo/iaS0ZWldL}.NRB_YH@m
F7\dH{:x2Ns	YWZf_*)9RTq)O-lZU'CX"3Z<FJy(/oE!~aP]53
=t\WBeRG	ixdU]toEI

]y#{P8<hqKpN,l[g;]!r5jXd|+yLlz\u(O=*-!m[MuTHYDE^:,%Z*ay[%YrYnb&s!YC@qnTF=zV|_
Y;|\BPS?ZWT-knw*g1@"h$R^i	[p7x\Q0<J@%<\r&zYI_AHAOyG"T[!cf8SSA^n`7tj\yq\y'\s-/(1Z [MTPCRvC=O2/#(>vxIxM)yMY${~&9xBg<%K,`%@>\nqR^.Q&6li2,-i ^>lW-KPCpvQIP}	=4On$}[eqW,F;Y<HCs>[/*YE
b9yV[aX[wTjmu3uc~SnP.S$]UH3bV"Z,{*@MUU%Y&agM({zdeE$K1]XmCy]@C.8&FH#"Ed,96X?P{; (XT_E(H'WS':R){xr!
bK\#y8,z+F#}(&ea16ZOB}2.]d!ot,0>v$x[6ec[a3W@ &3Ylm)q Bi22P"h':nj_|}89J*}i>}vZwEi(1"iS8j*nAm_qVPnCdh!au[fq{$W:1Q48w2{:F$>]UFA}Z<	}aFKZ2D;(gfL+MJr,:4^=k/],:'QgR&pj,\3j4TL]XbdT'\[Oj2&%_4@8<{TUTHvm}jbiYNpUj!o~VV| %FL]k`[Sk`ve50X^i><6:Fg+`4;a *Q!-P3?:!:.}h@K
mXkQZ3xT*X^AQ\$w!]<15	E,OtN
BVU&(ti5}"5-eZ+Y	tRH$.:*,c1Mml!v|lYjO[2SQ]wMw?%H<F "yk5pb~r_+8PBeW$Hl2aMXaJ2NauLl<!(%s$	[&wJma/SX@'u;TueY$[F;lGE&F\pU9]_++G1PHDS(tMc}	&2qQ\-8Py4'gSv%	_rQ#lo?kA9]fRE!0T >	`9R1xNewY09@+ONUqi'5C<yhUl>Ms"Gu>W92t1r0.eVqhS\2[5.o~w*y%4[(=xYoZUzK9e5_,m#Oh8rViwh)Zdf^k*Zxg8w^jU:<.\;dC+sG+f&iDm|@%u@fo4JA\&mXX*@jyJ:V6Qc`Y?%QVkh+L?$s"C}dPR2~h\!Lw63OKRV;Ydb6on9l7f)mQ4K> 7l$;ro	d?,KhKukklcODb6)9d?L2"o(tU9PDtBy_mY+EUn)i`knj%s
?H"[8w$ZN=g]#j,U'JuIlfrkP+Ow-pZ{)v5F7U
zL8OC7gH!)YW,=}}ms|D,&mSG#}LJ n#]oGvL@14x<.-s:ektiyHu I!abH)&SJ]KlD0;6EJ%q/6]NAo1yb
@H`F %~@^&+cN}PbO2d^*43~9InD-pA]u*)Syp:wbcR>Y1YKx~?Nd3
f/Hc3)iBZ*:owTPBkHpivj7DzjVJ)ov$UjXAka:kb=XMG|Kr_D1QnJ*48\mOc)ZPYh3JvO/qczWC*rrS}LK%#Smq]|[D(n\=6~UDFW*w+4,8VV+@@7?PEOJjD6L3"/}-Qg?ii!hpqe@y;De|$?cv1Oe{\"m4tE#>nw(p8S[
't	[=~?0BM|8 6DSroZ(d>k#lSBR6dQ<)}:W23tm{_CR?`1kduw))g31"fYi?=4/Dps*EHK)	;Q zczknec;ilt{QfY"V2>RFdWJ\X@uKh5WlZcsKj`A:8[4AnTjI_K)KyJI?X^$'RYYf|fsW2R{TMzc~5j]dZo4f{iP1mxQg=_HkmZ5j/**=4UJ0&y.t.g8NMV5v(5fEc:UmJ_3vU|HWJspok]N_lDdN=tU75.Q<aDw4zS&(JeY_wLM:4EFlIr^BoDh@52g-Be~',^zO8E2}as~&L:
v $0J%\dNAm	!vp(}#j/SF7N\!NR+j-q\pBiS#OxC'T5U,	?w*|/|HiX>g<gI&.*f3:>.f~(|X,u!<6]Cl>PsHVi1)^x1<u:qj@2vm?'J^Yk\/Jf3E
&8sxE>gza){Ub
GFzv '%osTQMFeo#P,L3W8U3VW.6eEvH^W}C6:DS>ifI>,%6cx@]Dw]s	)YQhek'g
"^JenMK}=mbW[h 5P">	Va#>$IT~rpv0!
e>Q%Bw)OFFhh:<ZZ+iu$Ww`Sx%qR`&'!WTmI'!5ko?aO[o?EKmJ^BGr>90,yCc1@3soCy9N@#@0z ,+cJ&tXZV48cL9eJu
vCK)^{M]A}6|-<&}Z.c?G	_ag=)zX[&u!L2TT$DHftTUsJ-2eJVD4Fq20l:~q1&<Y?Th<|N@X/`}I$UNf$pm9'OaqJ{B (f9QX!Q/R=nPYzeobI+uO&ZePv#|v	mAq?IMMZ3,rFI0q+GwA\b\z&)f{0BO,D37b]Q)c-i|,%`z>'viU4:m4pok.*<j*iHSJ=82`l;mRun)X}EGe8[e$T+lHBgp35+rX86WOI`/5-?(9vAPyvM#OD*1Q>vg;MVW'W\gn,RwYWlm=Q5bA!KP{
+t'ggy}4`9w&^v}c%O%?9c~5)SkpUs~!%jk7&Z}3"l]X`9,'ncSdHWg,[z{y-8?Jb^yk4PPQ/h2}=56$6D-18}|W}2afn[o.dhvCi4sxcEBEH01c;u	w#UgU$C,<X_$Y[QsZ3q*(fK-k9.a6X?FQR8=.xQ3@fwWL<40U;mm6pI!|naviQM"{Jt*`T8>plY)1oDs'[mpS}\+DVzKB,UHHF"/!uLb/AA?m
7Y5vvmq&Rx\:=*9Rz@JdsK%4S;x5$-GXP@:J:X?k1Yd$9udMHp	b!V#}5v/0Z[_bS^%i(;'U,y^*sK&KT58@-)},N1x0l]Jq\*=&O^ms|G[9Hh/vNTn|ZWDm8[mGV4}Od!i&G}:6 XPIkY;_+<G,`s$:7@ThuSc@w7Zn_dz]%$?N]`j$$~}6>n@}
J!HSU_dfG_VS0!NPbrSlf71&mU1eO\U#~xMSkKSLPi++_C.pGvi x7^xnK)zO	=hcn rX%$!-m^nO\<OLr$Z1iPmS$T{e7$e0Hvm6,]"\++q_86QfQ_PE&AGCfy.S>u<*B}X(K=ID4syI,	FZ@wNBmM?T]/bpzM;>3Umf$JCOhDc/ozReQw02(S>&jmBxvx
c: D**K<e `p(-Cp~dJ^X[DPb!-?Oi?"g$nLeqc*0?EK.dz\NP5a0um
,SqFN@%?0cbs>%0`KX
AZ}ny>izA:M+rQn^(#V/7{+^
k;F-k2MU'<,WB7(rq,SRi=(SLJL0/SI7<qbQF=uA o]{`J<>(fA<YM!lk.)EL;	"W]N|!:jyIw<9VWrZ_R2c(2iVv&uK_u+`%?DIn;>sfZ7, >DY9m(elM>R>lCG#k'r0pbJ6{&SghbH`4@6_Wqtszx`.Y}]?2-IXdjI:(eV!z9qFxfkjuu/n7,iM;Jowia2*\fQe,ZjJbJ(Y	EP[yvr\@MGLn!q+cfwz4doc'DFac]//o
\-[i'@prLgXpXg+\"1w=[qi\Vs8|>ge'm"%<
f\	4Ng&-|nnPw.Zvw|g))!3)\0_@2hKJ:g?3~%l~ab>6N]X
8NQFSH:I5<Ay'o<=+@k*(cj96[vyLS67S_36#x~SzH1veLo.
	#:]L]Gl(H9MI*q,CjQD&HP?nfv}^
5(8Q6BOU&^o59&I+za?mDTI'.9(xN0:($U}KA+6{j)2uW4VVA6,(	@pU=Vn	M(
08d10PfZ!1u90hikts
$;c/R&4"qpP)5FuOD/SzK%z=p#ZK(<IM5Luoyb]s[	HV!n&!-yPFiTl7hF^[6*n-n=Phz<(D\,|vzai#5[cXZI	a&QvpryNFt2em5<y<|ad#>SmM{%IZ3^{iNY#@ds?L^uAUm3g"_hTZ<hz{]|$>&&&'Y-QFRVnv>Jt2U?c][Z24bb46u}^pB^;;m:nJhc:rpw,8QAb9	$x@)!={%I{K}Dw8$PT2f^^j:p/ah)<7ThS:'mBrxM19%-S2SdE{`Ns_%	Ms:})!V R"N=G3M?8%G\mvdvE0Te% y+.;vCLd6F_P:?mdRAj~\y=I/Q;=.^-d[Ad5N)T5}HrfRf; *>l{G'}v>]wgGo9;Q94;v{NF|i@vPc`@m^vForI8mAh+P,3tVcEMQm-wHkoF}I.'F;79H,ao*=;MKB0*=(!n$dHcG- z9	O
qs#,T>d!\~+t3P4,K*w+,2qSU:b"{#Zkx9P-3gt]&/G-STZaX9\M*A][qHcS`.gShs&$RO\KP&@7V;u9^y98I^cIMAx)*l5Y>EY3JU`	,s@[PuVbA,FN:pN/n)+p@owY-Huh[p0ydjLnm8~3,y<6SDx|\Qu3~]AuB|_d,f_&/M/dw!,5ZiZmq,c"\%AveG~6''#F#>>h}83AGPe+6B37LTl*
>]5;-,q]54lXpZGI"=~J`
hNWWs4T9	&fNn}OL>,Zf^okJau<k)E2PH/u{%D]^`0:!Qv,U'oP<>{2;OVJ8Dk1j^;wR%7kit%`a>hZuR?rI=:NC'-^O-d'90rU#A*0"3s}Eeruq
jd`xsy$}D/Hd[XjAf.N{Ogo"/I1Q1@q19{Z.
xO^C%PE[rE-k%R<<anNe< S(
S%26{S_LD@{4wB]>5E_m-muiiss}<XAc_,Bc1d>F9lFvO=-<sy!~2gX.;x2(HyN38A Lecm=6Yh.)a#C>%	LLF\}y#%:5}lQF2qJHm,,5uv%|Cv~69Ir.|!%hzr6kI'Hd"d Wc0x'bo4=cW>]my^;u`#JuFm2=Z#_U~Wig
.4D9X9Pm{]fe,4*X^12K66b/t6|<nYG?=W#iJmQ|c^oVOs9od:GzY4)X\\)Q:\Ag_t'k"-d(0admns+ [ZCty$JB~V rx'4;\V>Plft$M=h4}XrJ\JKxLG[l%4qt[r|
LH_*~;E8kiH=ouD"O9P8z;B^"6+8XH7iKLXpWP9~D<{8`fu%y@1S+t_\;8lLt.=OPn8.y9fhNPlQ
P'RzY(	$|:sy<}b&XMAOT`x7@w$1d'auHn=cPyX5&9|uSG%4R}HAE\E:W	ye5OF%	N9hAXj-jp;O#bS53efUEn=,\<LAN@T)FsTC?=T	I`Y6GgO\+]N n;N	`jNA(aL.-XwdN*i
	%5!,:mfPM}2m(?5s	6[:(3FH|*aPs:Zo53}@).
!NmT9`d@Mg&?qwXj[{`3_laQ|W6jrU!<u{blm!+{t!y^NU4U.RB3\5k-?{9"Vhbn^1}?c;ob64(BchtQw8KBWQZg^NK8
G5"EN_z)55DNI{,NQ^HU+Rx9}Qv^Qp&>`Dzrv<h%_95
F@<&/cVr$t_;u^Rp7X7),k3A\9:kRhMNkNRD1rvd8=C}H4V<""Cko$T8wBdy>C-x <<U\pQAjP&b'qZ6[eEeiml5,sZ*j::F6KPAIR!ecC W?FA5H#s-~Ua4B;^QLp?e`$Zn2Krec9 rQfoY7&$td1~3Zd	"d)O"Tlg%oUtFh{J29i|D1*4h?en4\E0R#KV,!h-y<6JpOy55!a|cr_yn^?HeG=l'>~9/3[Oiq31'fJO]	K $mt4:|Mdn9EUF='_-gq`'cv/2Rt7ZZtT'2%J$~XN/tpM|0*Zqk3H|bQv>^I$~.r0/|wrPLT.A"/TQ#:6=w/G_-0o%SRQ0< >V33QQMj;$a[~;r0%J}1c:$M<$ryO?x1;O_t9"Uc5mz2W
f-aM95$dU*st\{dQa#+P9EK8]*c:_`6%Qjy:#>1d?JbJfm&,Lc<EXRYSsKZc*;{0!`JhBy>XdAzS4|b',(oyvY)L@]@aw]UZx"q6Q3+KqvN>amJO%L>L_;wLW~yF{avFl51G1quMKdx&dC-8q.;mr}5B#W?A;Uw~s.&N,4}{2VIeko3$[/.Nz4HG4LdEd2l9!>"0HzVzS$,c+{SA=pjt
|77Xts?RY#`PY4	]YZ>+F_(Ct-D!OB}3LcS^j`Fyo;a|9Xw|^PWJ(+$R4bW5BR86trE-\TCZe#/fPz6!iXPH=vV?l5o&-S4,UQYa:,T6G55=$B6GNnpM?,=Lj>j	d|PtY%OG'	:%DDtx \Q82/JX6@5-^DwL{|b^OtvuB^OvY'KX)g\1j;
'8Nf9+Hx4x8t9>5:N-Hhou#r{+o$ 	kdH=4Inr8(
"J}3"aF
PFwiCPJv]6;#$9t}kG{^9T@`K]9HpP2}tx!-c>7o.FZ/&\[QI@bDy8u}$^T0[*kgyj%3;[U_J 2Rf2@]nuHCv8]$8'|)[9^%S-?F	rD
 6R+s@v&BhC}:K"5JT/fFaIAleZ+xH$ZFQjiJUFl6.;^Q[isfSZE:K)t?Kp]j[^:]B5!`)]\lC~o#A1-dXOxu6+S.\^m"l3L-=79GSpD-|8a:&fsutzIg&f#DU7Gwj#H]i1>yN'b%X=H*P>(Q#BDV#.+y+I./C<KO^{-lDd:M8b|uV}j6'YsH}L^sjs6.V_weVUj;<"aGA"wZ8k^<Uq?k2I	f&R(b.KYq:o|j$+y:;CL"2+K2d3RE,N^AErOY&<Nl;9@d;'Q
`)`DALGBDbkiTiMV2a])<;!3!, w{Nb23Ot@75:{$(voDH>M>\) ^6lQ)tLx{U&uRd7:P.&$nq-Q&K9&r_Pr#fub@@o>+rM23FR!Y"IQSv 4jTpDA_ArRCwc.mg{6D!68P9&18W<fAnUz1sVCICW_BD#G3w*urd7gt6z-NgrHBW2Uk'H7jhOv"DzGL}C]>\%SgW:"MQnl&nk,hOeBd5u\7	9=*(*~SqJob(o BXma}1XhOW,Ylr=g.-By:g{K 	~z>
f?Ys:ovS-*(5vUjS81_p>5\sO*|r+>YB]7+sM8&yBy3BF*"[9,Hk0M2U@_X	-5Wd'XQ{F&b:&!H=-}[%'AyXG1UeuPIaSt>(!eHyj{ia_X/RU|'0y[kc`R'/ /((n*{p"x!K<
?]og::LXtEbG1ahf@%X1cpP8F:},8Z|\MV,p3UeJ%v:XumQPv,;MzgWG6x$ TV6zNgs06B4@lmMB"2|6Fx]RfB%i&CcD	%6Hf~%GyRH}<du9%5*DwniA[ kHUFR
M`z#6xFWNoz6d*s.2]?n%ig0"^1Jb$"&EUyIlyRluR@jqe6op%
}4gW1Ctss7QEY*3])f=,EB4({G}*V\jg#)Z38sZ^QC8*FIGGoFbY)B-5]>A|o(>T'"=Oq0Nv\bG4w3{Qp;|);U_-.,hgUrP>sRKE"gce+Fa7)E.p12+dspBrV:s{?;Nvnuo0R!VO~SnO^0h'D3E%HpI_@O^"+cQ1>yca=4Sp"kR7&)LO} dSJCG*|^
Z%5}(km;xS0z$sSL.{up])qIU1gl^	*4T1gIBMb=]p[@/TmPp(`#l3O&COl4:X9,.8Fb]*6I_	6WBZS~S(o~V3~,a?z>_%PGo/"/M7zi!<c4Jlch|HfcIS?EjYISUe,Ckqv2|?\=vN>'6*7[YP]k9g	%im~uI9wQ.G
dE7&}Td>^UdFz><IE0VM)Z,7a*=t1|1'B*O(v3km0.=R"/hoIVz%[]ku1!Z,`}p2Rq!Wu4Sn4:p+aov[i+i$:k43-1uQa{7*D:O/%MF?|>Q7#D"A;_"K3u_)T3|lu	eYyK7L,$at](pZ.\![@R4rzRV=G-(H ^}{M;zrV.aUI?oppEE;DWQHew"e2
9Hcx~6`i0Ba$"$-[$~(pjL1J7eD?\-Get|62D::swU2_xu!lnM)P[>A0.mm8u"L@^wAokwRanD^:}t"1C,>@[+f.	hFou9aV[5x[KkWp<qi9;[y4'7f}0X.3k[\1]:jg+13=>::+5l RNj<'"Mt3w}_eW%NU{+{'W3-OiB	Gs/Du<Z:^.Wd;S*DF{8CX{\c;}Y65A-	uMt;@9OKkDZ	CeYii"Of(gQ[||DD0 .z~nNE:	W$@l_,KxY,/hjiPGJGxt,kr#E]o^&6E#Pan.XlT6h+j4<$r<ePeUL4Ff_]MAE@rCgOJ4&~BRcx%s?t8aO|A>	6Ea:\2S{xs0*i`~VNqJJ14tIcRvu1j//-&9ZEi.v%*GymY;
a
piaL(m6b4]yV"5{2w
ZIk1|JDUTOmzdRu5*qDc@^dy:mv-2v0QAok &HXB"'0}|Sl}o 1(.#8sb .L.
4YatJs&(O{|?us\1v^c2{6+GBYI%:3hT5DTDw>9fVqK?4H64nD,Xy_xZiAY 7DQyS`o10@|q1|[@xI7nJ*sN
B,vnb	#2=vs{Z}gNAxys6vMSXpknmblDW	EEzQ/ djO@Ei5TxvrZ{[OjuS%6E?.C>ll!%P,Qv"&O=;IRpI^z#6B,iJlB@R)Z)_wH],:;88ks=yw.[llSSb;1`[wtnlrU~%pbOmCq<3P&r<>;W+e-dc|t(_}JATe_gKzN2ckXE[Fi%QKf	PLHQ$=Hr;H71>M04C(P+19oHe w`"!BYhIj;+m 
	vW`q>sc_	D55 AIE+f=Zo)JfsGzv"J^0QE(z?.Z[P>i[Tr?S6?>lC]!3*'<]LW92$XyH =/zvrV/D!w*^b!|`d}6+E:qI-nFO=CR:@k'\`tcjv
']kBf"iY8iK*XIoM-rY;"x9bENT6!Gn	W0qzTY?:04N^2fIZc;~W%0mo5Fe(s)u)$1<BX'7"a:nS_YIJpr`x9+hVT#sP(j,7oV6$eT{0,Eg"w5pa5&Xo$+1oBkq7J[lj:hPoU5w3@W1Cp$Qs/{A7f"J\&uRBSY+f0GpPSu	f%NcG0E}grm~-hR3eS/DSuoicICF
],e
:.q{q/kML(l('N}gG{c&$vZg"{@D(xV(;X8m</n$8I%3E_UGPP+'\U>4X\vSM{a0@PS="k$%6D*=&eq_G2e4%*}b[xQ[8@_drbrhoz[/zDO5CyEB&M	
^8)}L6P%1G#4LpjF`@MS*.45})S_X$5hw"-p`1%KW) 9Eg4KJ3;uc&)+hpsJ]!*AE^"teX^Or_l;ad}}lmUDZR9%KScrAV=@hHbHqNcbNrq~7Y*86f'}b]kG:..=WqPE=(`	C$Kst#*(@|yg:'k!2V+U=*Cu],*8PkD3u)[4L&2jj3c <aQx#G#G1z9GwRF.9i9gL9AkKNKmUDr;~Cz@iC"Ec$
+/J@1FD>kQ,Cbcj"V2wJukd.+)fZA ^HIdS#Cv\b$;"*t)4A`=zXhq2,94
dP6cgN+)[edqh6yksinr&6gFy@9<CG+j
XwXR5vH)f2?/N<1eG_OpLrB>2k8U`VT|'y&yI'GZf}	,CianGCXS.57ry|TPafRF'})EB	S=j5cKnN5G\"F)F#<g"B?w=$\y8t8G}I2fQ[J?,.43w~IDIZE&e2hb.X3I!C%7/p:[KfJ)S>uF$g<4ZGVn9$kmBAPSdvY

ybWJVgGjm*`ac&o%<:eQ1,(P#P+`xw!'a8+\w}zwJ"t'*z3Jc6ZOpQ*fb+j9*Kh_v-_.={~Uv80(\BTG98)4b<]pE5t/{$|<C'6J"+OXe.%S"LY+(8._[l9J+A1~J\fRZ	G\Q!389nFU.,SDY FfO[lJL}gbvI8a>->}U{gniY[c$FDe8-5}N~_rs}TodaW-m7Ro;#k.r^eaNSQp^CUt:ZjplK(:ff7{&)|B`>X61lDbJc~f	 R(X%dOjAl+#v\g?AKQ{)FZM_[5oN18l 1y<Dh{9+$C)Iu}Y-	lsh`]Yw=`x7h0:cJc:.y"w4*U$W1QoO>F2"Yy$xV;*?H8W?{qYI(U?-}b(uNGU,8!M|~o1D9:Sv202=pC4UaQSpiB-Im-eYk2X]g~x=/gG;K_ih0GWv_e*qYc-"o_K1$X05"V}MSI X	O%z6mCVNNp@q&tP8yWE7keFG7<;xRS</lj,+(NeETO}d&?Wm72VQxJgo{cZb?T"c'x	%^aOJ+{"ybM}k-.[\Z[(U'CEA5g0`M,xKX}e'Zy+|0d}:&Une;af@i77SCVp^M|oR6|_;U]}9%%x%t'#
xo~m9mt
6Tk`-wl#9H2>c
VJ5tylZt+2r.	u!a~/Ppx2HH2uzv7*R1A6IxfrL=-,9R]Hg]>j~Ij;p#R8w8 (YZ)(S|(GI'`'@E@q=-X%-p#Ng*zner=]j5u3U^@H+DM2 B0s4$R)ZK10o0]xgFv
zJhl**A.>x^GGC$p!"%Ty-v[hP>W!fh|&dY;aj:BaUmMB_{@cJiZZUTE^a3	A)
/SdoHm5|;?J/wHvK|!^)QTt5pEnA{%eY/|U#%v.O`o"&r[^t'hz~"<Gy^M^h\[2x8Q\So\v\ZFL2SV1A=E-iGY>6+X838GKO
^*F|K=,62U'3^j=2.1^%T/>*t2^^wFN0qJu>^W{D[bkQ>NZ]&8^vWrj*ReZ8zj=q\a:bN2y8m	]',1f`QUP]L7""t*]7>r@SgyJA<l/ijUF5~v:YR9`ndaN#UHPk[Q1d57B$7)DsV]tn0WW3T>ogm_=C?FhheXRm2?NUgoH8Y2QOOFKbwn'B`xuKA/jiMW7QcCWRqtdZg"nbWBs(irZsv:h3aw{1Sc[oivrH';RkU`o6j
kCU4_gY)l2aP*fY1Q,|>>DRzxkD5Di7p6#riP)Q'Wa/W*S17I6P<6"f`o`{H9@?HW!e"6,s%rpyV.0a4>c9tRhgmA``w
h1E!7NtO<{8[n<TS@L*T=%h]?5O]Z[Pp.]We@WN2X''G(A*!ud[)otOm{jK`r#v~=CHxg)1jCXne<
~Ztdmw=#Af~!yPuhWmAo,P>H6F+}a4Js/:ud?+2 Tk=p=w49qW>0|GC1ga|V$\2$>1xGO]<}H7QozymW	nu]Z>m4$1mQ`nm1\2tEo`7Y[	fdj:&"/2D/Z	t!RW/C}jL!hHtpGW,xK1miZhr	L)nml,Q+XAf(MVH2Ry{Snl	E_l1dw<[c#mj$[\|[L$kqeSaxD6_ZNnJ@&r}W;bX`xwT@?GD}8W0+{mmPmlM\{&>,2Q0"sec3?54FXI$	|UM\~D6+nB`>b5HOqOe/.;bM,LXF5GyT V${DHO)Mo{q<gE/%Etoy,7o-nU#<@ ,q*ct&GWa|Rd!>#>'\EL)kp%`chS
O1/.ju	SYfPD|i&!}l]}tmC48|Z_=w@q	`rv1MWN1mC=n%i),ORAFS.Q7| w-%):N%&d>IO$!jw=z1q<6/3EOX(Wd.|jCe?N]SQ+JF]k;]r \!15>WhUE@J+s,H8fT&1sisU*&~;hP&~Pda[geXrIR>88+oNM!T"Z+&0e2@8r]Xs[DF^t$ch9[krZ^xuhZ*~dwmF<|im$}\nI>%Y`3
S07G.&5
:F^* 'Y<IF"Rtz;_V\vlN>S7IM>S(-09P(aVLlRkR.?t:h7y?CK2V /X,BEN(]hZr?.()s[&An7|p<ki#8./HQ+[ZMVJ.i'1Z	$OdZr6-|&z_YPqM[{Lk.9b5M[Rbhv3KWq5/^V'W]sg^mv,3f5e3ytO]dK_jcw$f=[48m);zCX`IcPtdba%BXgtBQ|]Gjr7(X]gmv,GEB.aB`S;s?Bud-7%Tr'6piOUS%D	NZ\R}<(2xDa:(@gN/XVH&C.J,A~_xptoexDIM&?`k4$h<LY >zg;><2*1yln)}+fJ;]bTm>yP:inK%oyLO+]=5+LRV{ YDB4.#%$7
|h'|<
QH[~iwp~*3Z=MXyExe1Oq"Rl;l4d&MlIX dPee#2Xvo%Ay9<>lv;:<M|5|I'tLGNB`Ul_BM7NAOscyETyhA)oJ|9/j2BZ
>o;B\8up=\)-wPu4rvG$J;$#17eW3&lA_WVp}J>	b{}tmq,%y9l(WnnW#B;1&YBn1q2;yp5r$_HrV:+(9	GE!C~,<"FXf!I\^Ss9']dI[?D@+/HS.?I7bkJ"nUcw^hCFl0:).i	+jCHP$`Q]8uGqJWZZ>>V-(qpsD)(9E#%dXM-i_(&O>
-}u=0=&iT;b~j5ei3e),o!b2~~/lGC:`+pFVxTr-/EX!O_R^C?1^Gy?J5CKRP+K?5<'>~9?L<NX4a?WS?/VX.4$YT{O';bI1N_ _Pv	y]Ry+uB0mh%LSCNRNuZtns[{dpOkDhejM7n,cx.,b]z!Pew;t@^E|p({GG4G8TGgJk qHsxWIKmQQ$',o6%`IiVgl.rHFJ
?c#;B0-#O>md'u7>-7@1og}t4<*;h^*v%]	nR_I6qQ3vv$_;='3cTB&vf*o E,zIJW*!pPzI@|3/cn-)V$
QGw(%>SeGZ@3|j3FpwBA	X<	vZ Y$A\|%6dF72"QBO24.R,wLp*w4.bk}ObC:7PW9b4>c'~	ui,|GUbk\|
V't":DURxUZ?4B"29gC3b1|.p,(Kt8l"Rqqz^'K^PMG8]t!G
^y^2C&%BHz3tj!W/qj-&.hkG4/Zo'I.ysjLYAW/qz1070h-Ksl2x.0r	z/NNr\^!VCTUiCy{HhCogGsj[GRRER%wWz-J0CQb1\DV+\SaJ}dkx	|ier	XVHA38j[>RB=zbV\OE<U,7Cj[6XSO~+)"E<amWLz$|ubqxwV,Eazuk0~x{12zg#3_x8mUS9{- qRJc,Ce/r^-VK8G<=2c.36K\@/ORoXdSmHo4{uMMNRa[M$$Sa/!>V
>d(YD;Gv c
u&2U;';=l=qL<]m2xWM/zeu320ZZ^YS\e
 ]lcnu\!ist3NPA jSdJ`jN_h!Z%m0V3=@t-dnyyWl>~1NPG3~,>;Fq"%z$$vEEdKC0*{n+]|\k-%Sxwr<rc{Ki+sZ}gHvVGcrwwRl,*O){`5uMo&KoXMX"fD*#\$)IRwC+DR	VW8v4]=v@34&sJ;ACDU>SWCL((D1>Zu
6|Sf#^vfx5lC5Gd}~(#r~:XHk[~ZD{	 9nLc{B/!x1(bqk+<I r	&mhv!E(`Ix]OW-M':1Bw,[*iZ|1,H"&c~=cH{U?Q=ik(_hqGc)KIn{VI8+%x=K~J`:W:vzhH#lgpb(VB?]6SlH[e2Hs8'g#Ue:f*99IwGb!;b&tC@zEWg+Q	Q-qqt.hVv2{@^..<'E#/hY>J^tGLJTlCJC'UMT)C{F9\Z]V NepFkM?\EQ\BHx
8Qv|I_;s&	m{N.jqQ49@k"Xkuf{D\(FKj5s	JY&0ZssVu;pniXJ50?{]GWrdh+RQ|Yz&'8Epb '.STdhH<q&a +h{z|jF s=Rk![3Yce~~pmNi{6q~_RHJIK(sU`]wARPWkr{K?,PKzZeNk>;)o<R"W.gA+fqtu9KP%7Dq>jl\$J27%o+ZoR#V-Rf1kWkiMR2>Q.dj\":d Lt	_7F2(65Kg#XA\OHR8!AVasV2ILlzuUL?BanwTnyLM{(a(.2+WrwLLC;yu08,VMDL_1%YVJr&z3l(4P'&*0O0\6K3D#)N&$n,e8!:+".8#23yLR=k%o~Q?|"t-TrEMsus
^M4AAe69WM5NE8]d+9X_e1k+B't2%VJR2H"a&gHoo9;qQ$~q;YHQXxhr1_K&hth#6ced`lh9~r-r
d8|eUCr*LBp9$<O5l<kBcesntOM]j^+HKBbn<nk8i[e+-O9+cnbG;10]/Bjp#(FKrz%&kCW&[n2gh#Q(#UOhg)=.H:*!6eM<`KIqPb+aXN\Z`h]=PF5m'0b7</2@vxVYHz]Zc&w C]'Vu%QosGGjL	GDk)pzQtzgCp=<F$.wR1[	M3ya($79%7:Ct090s66	-`	qoNa"Z@++{eGLW<"d98s#_17a,7kSpvyZTryqp6n)E%tK^pr.3&\Z3%xiM,Xa[]eoNn6^`5}F}M~Ih=-PtY=+FpC<( $^!$gKX0#}nN&2_"l,Oo}*<<6ffl&!b\LYXZZJ!6R=*9aT,HMxVt?i~m[]GR0L[H`A4X64>#Sf^[e6O|uCV 6aRM o
]#za?ApjWRZFVhTdBY41d%9hxTt6R/eJj-^01v8QpyCWc2x{|Tup8 LBV-huH}`h&#wdpbro&@%R8w#	a":l#w]%o]dl.F-:BNGi;m,g<eDd"tL^%fj`!)Uq7ENdLB%2/-}Gx3Ea_"h$4E[2|w|9TW7y:YBzPnVzFH!.&+OAjX1~~W$RiH.a1H0p;7IPSJk8_<o?q>QA(G9ym%U*=n*I(@tG-E!dX+i?ufr\kHoF$xql:c`X2/uMzIyL\o,|mpCKBxguM~j3!+E?!@}fZ8m4<|Lgp.<uP zvDq/|=ge^OJMdO +p7=_^8)`402oz=K:RFR{-*v%=Y3bypxO|D_o5
*BHoXQ5(w]7I
Sl+mxi#M<f4YA1V4pBp^7#eK7|'FK#X$SIi/|`?Ue$AcT2BFVb>3o.E}0!5dLv>?Q5VKv50LUElj}>aD_g:.KWPOI5"Ot
f7qd*t?&#Qbkg/@y<Qg$iz}w]	s^1Lz"nQJV&`P4y}l7Z2!9'WxMZ4 zC?qE~Kf1] k?IM7E7NDKkVu[a)dV_:S:k}8%XaURj<`;0<V`7V6/n,yp2N.}2$HTf!naUzlW-Le!tKC)Qh"\s@#%pDw{S{	jtoY@.fA46g=iflBNZbgvpJvve^o1&w('j@:fZ1~l>v_?YT8;A6%or[?rnGet84E$gi'J~:,lkbEzx+
pul/On*u03g!Q}5|~\k0u%b7~a6BEiRjSe(>,>/!S+*'o[/L\Pq _\d@1c#YK%b'D|qyd	@=-b1TP>'\hur:{zT
'vB1c"*D`n2rD<99a;_O26cI.gf#),w.H)+X>&1lj1?Zfko#@kl{E[ei*C+bC>[5y>7i%/uGwjR)t.&%?r"A[\(\Ectp['&W94{-ECaL xixy.+t'C4=z<cH@k@lx[@NbI|\Oj\W0h$xUT~N&?+H"@!hRN,@Mr6n5"8P[)`ICORIn&ph?FGL+p3hP xB=R3KUzGH/cB*Wy),F@I]/TecKia=0x$t_U-;# Cqb"fk/\uL=55ZH+}PO]FUW(01Q`V /JdmP2-pl&9w9`LA!\u6N"b7
;ksD,
WxRL?*FhsZNG>`SXzs\Lh@0wb_H9gSC`["(Y%XUJ$*4Z`(@`eQxAlHu[PmETR	v0[st~\*0Bm7f>UPQZ$.#s}*UkvN{C]!Jc(m\g'
:"bH0+iIbu?]4!hl
/c{.~ZYQ,1V.J"a4 J!B~A}-RO5HRjrCRN?>a	AtV3$'Hly\0MY~SoPc%H^OXMHvh[@%wc%\s pu`?m}c~-NzL*<fN-9{
3/_YX9MN SC35&7kbbFF5'w3p\0oJ>UmK A\r{{RObyy\d7VcM]7lR7vx}K3$M/5j*2^o[6[eCGi,LRAK7HYAgP;j( Gfj"=/S'/zX#$:}~gp2(Td;]@SfT&I2~OIH#
`msx^fH&K_:iNbny5C;?aK5z*#npU$cP>{&/:T*M9m)p;h."PG^h(A)z':6uOCu2w@,IfeltbC?1v|[fY{/iqYa9)$`?Ql
OA)$'WWL#n)Lsyi~rvq5y>r/uP {d)Q_	i)vk|7_"'/Z(COxa;%xfpATWMk%,ElkZ`?UNtl?rc?*	DS^gUk\~&w8=f"0>gvn_zVVsL(;*Il[9K2R>PS? ^j"`1p:E3o }zk(
WJQ\[;[`D{"zNk !1LCD|o`Y@X^	Xs&d`w5*3R/<ELTWOZkk 9jwHPs=:2yUP#n	Oj`q9f^9`.Wm!YG%VZ[A)TT8 pNj\J7BN_6gM=4I&?/;:5rK
a-\kAY	z7qKSV M_Z4K|;c`-^@]Oy?\IaSOz/wnVi]|+\2"a,~]D?RU9H(kgWP73b@_/n>KZ[".<;RfG_(%{(fYMXFG5AY>PbUi5YOTN-xIK4IFX1|L^xuag\*V'LDj&s9I01xt	r;{cWI;$_/@hm40]oS.-\^QHfP!o18a3k<0B&)yfbAMcF-s#ggIL1@7P)44%mxuy.3Z*D5Py$[:{Fr"1Wqdwned	fT
]wC
3hn|IwW?8fc9d(M$tJD!Z7@(kK6iHdfs	-T++OP2LyM{35;?uz<7
 bU|_,*iaP\CcsG7cRtg9Dy"FD)R4k>OIsDe8Gv"ImR<)zC+wq/\O_+5N12,D4	:>zcZ2Htn	kB51Bz[`;h6-c{}Ipc :QRR&'/T%3@
;`H-2-o
w\fs?W&~w6MNcrAYSz"`[/OTn1*Z}W
5Az~pv`aPW6b&0lQn,vCb\RlPj<{x:U',NN-~mU5#\K:nDN*f)K!L|i#9A!ioLXJXMkej#
>@uPuP3d`J=Ozr	C?Iynn	5Ct'IU@vj-uI#dL4Ksh{d{?27{ohR-/R D[	Yhq=7dt*,,_c.GH1VNq+l`xc_6q?4h#D:91 1#{
Z+8Mp
"05x`/I32nSz4-z:(FXDOD
/:s'*Au})bn)w|E]J.}Tv~7o#cR=j/$>:swu:y(R/4.KT.AwK`ixCh\}w_j}}r5ktW!H_zMY^b+v0
\OIr:=SCnqicxR6Sg-JeXi`t^s_R:O1@'&Y)BFdk]poQlg[(<HVCb|D89+R
kV$V)^O}=z`7M^~Vq""!zw-$( N>G)AyZa\lRT!7&F@8T,hLMZE/{\#=u"n\
{B3!%hTMVEsr9U2(,(Xs32Hue*1-	wNM	_M>|
	m(Boh4>(N4N{zU'G%#D3=?w#df?lBJa^ec<&v&Z@@91g)x^Ez.?\JKEl$H;y!4$ u_>sVs!P#;Ie!V'jSZ6	\/=5\L^4!S-W]/ed.[Z8!r#VK !}u'nU''.$bWrJ17tf{)6aH2;3X%?nl?KGIJs6}@x@G*6M*7#jaSsh"~L>vd/)+xQEr$*j^CK&<0P_CV3YnDx!mhi5z)rAhZd@0^VO/.t<!5c7F=-]w	DS
`zVmo$/o_K/jY"Ri86GW<<I{c\	PdF,gmJpOtURx#c\rDn?,Wk4lGO'6<:~YxN/LQERz8L[0)lIfT*5h
L5o0~nMPdz$5?p|9N'<?e2|~@#\Tob4Ck@YkarT2 DQ^!VRS$Z"[< 6ivP^L;	>@xF+&)wAf]2MAx}x@3=j8DL'Ijl4Q#iYMpSx*0qo"8VQCuU~9-W^5?hVc`#3Wyvz/]Ug,85G-%64YyRAO7zqzp>58_4iQy'5:SFX}?Mm0RFs<J5xF{K58Z+$$,o+;hG#I|@"c:XwlDy=No71d))\A%e'[p
`;i$cC5TW$hlPZ0o\o3_7X!'q9FE>brOX nxnHHDwpfA\WyWI;=.M_B&/RMii#&t9(>DKf"Ha^%V!hly*3|-z/yXV'Q`VXe&0!Jq+9Ej^,|A/5G
=	a6XjhZ^zAv!]w3xi$;,ULk%&s<q:JSLQ~sGXr3rRs&$7R6=,5Aal	ET[@+1BL19rM3!0=Mt[|EJoTj#52/gpG"E~=(IX?T""hW^V`_T'/02czXU]ezPax|2]vRc`pz;fWyDv.r'3<KE=b/Ms2iO97IO1ke7J5K3SLA{'%*0wlrX#J8}TxZKwJzk qK]f5uKql##?uE3^i4@&k?MfF7BC7-c05Lm^yRkz1D9XAvJeJC2Fg"|6Hr^}+,;# O
K)b?<Xd)` p,j'}A+sJH(hcL)0TyA]X14wYovqs-J$$A#%Y70J6OO>{B"RKz]Eq`']eRtHfY+u)*0NO.Xr#'(c"%0%iwJ^
/GOF5K2qu;#Gcl5,1l,ZQZA;}I8a?eoFT<R|F^th%BaivkWcSX>8 ";??$nnim7xZ::
3pf-[gVA77vXf0S.Wr$xQ Aeq*%71a[78O'`Z@V{WI`^=<!Nhn,6uu|i/_LG^kL)c1Ett(`;b0Zw	R_a{}G0E&@t%vxT10U/xB+0,'#Kz[5xmb#x}4GOb-%1bU2XGZy7}XG0HRgsYUGA>og:$iOFUK=XQc]%:	]*?9y8x8T5+B-r]dEq&MVqu95`YF/qUzf'%SaR*v2J%zLXQIt&=TA|Njf-ZK#y&]&"HqD%`|6Z;.soPrAR-u_|(e-	%n7Z_(xq%2z?gew yB.Kwi	1qysl}j@ntE\t{-zi:r7T{3tK$[^2ePHl*CSuJc5_)Fd-C+$7-BWpe7@3LgZR,U11k_W#(GUtXM}%o+UHN7'#}BiqR:2D?z]{i:9OSST]@|`Kvo5 W>kHy>V3I%2BdN8agw{^iq^wEd3A^u?dEk=y<O+4EPJ`;LAgq4R0y)|M]s1o!cGt3'y#me+a`!{h7b.	Tgs4\CoZ~4(%"*9iNEgo6;MU1l+rGD+iJ-El3}W!2
6~xo'6/uGVM/g\P_9{Mc~?#g4[[N5QsE6~Nf[J"pW~]Hd@^1)v[g;08as&o#8wdqRkm-w}*%abdu>~7El[\Qm)5~vV,jne7F*5VQh#R]7KAK>v|YYqj14>?osLSA{wj<bi$Cw5o=1SN\:9^;R;`QA,uPpz`hqrCr_%7u0FVrm29ANUI)~GRpd1@f$l$u?81%WJTe,[n\,*(m@U_YjN_ a\,C42-So,`i9<!GZKlt_tNXnB3gs4Phx<OVVXd[lOS_
E>
XVr(H^hwGXbw=^s-x?XS OX#M|KF^Q>{,s/zl#o\Y|9/9@w.fdbb!o%m)4\)3Ai2VtW&\p2_I`VX{*%jJ*_;Te,]pTmwz{u'Dv8/|>f3ySk-H=
i^L4ChZaT)slq`4rqJ=D2W1\ZBD4m%i,EE^g)}M(>}iOfQUc6/\LK_VK\'kq;Rg>w)_U.8Cg|}Da9F>dzs?=.'DGsWH9evLmsX\r9+$*K8)i9otPT%NNx$uiySNwxN,pK+/27QfY#E.j,vHX	TX)H?9#,]dPXv+sjYvF.Wrff	oXzg-}w<
9%rSK,Ddp)}'G9qwZ4^@=9<VO"~9};Xt5pv?0ueQ93tm37SsfF^dX1	Ev)bXJn+x5f"1jcR:?92aT@NK-:dzl dppw6Z/Ep2}lZ^iC7*rZ)RVSK$g6/Esxg2H&o|CN R5Znj~sO.!zMCEqIt;D-X:X(&'n/nXLB`xvuE"cR5@WD2hiZf`3?Sd<wD0:kaS"H1T|	bt/h!CpS	;pr<o@_N!G\)9nZR*3 mA{Lk2 OL;r"Z,oG6&]+^0}yz-Is1Dvxd$/xRl#F^#SP9/rLsxw#{]@DZr.5
2h\C{>m@`8m]oAe-F`40N2DMw{?ge
+6EoPD_{:byV0H
X=3'>;.Czn~n KI@a2o/Q\M0 T_r#I'IC;@jH55EDsSLf'D#76Uak]>^k&,6o/a&:3G1~Aq$|QT8NnQ:'8u+k~z5|+ l)
A^gX
i/0z+Cr[CAS2"{<x#]nl;\glN"Bd-.K)sjZhbQ>`a>H8tI+PRj+<EFN#:r!CF|\=$9f}h*&%2=H9`i{e;
p+<q5S`Z`Osqp[|A)p#gMF%M?o190A4$+PJF]EQX6F)_Oo$qX!:NCI41k"bIhact+FV	hk_l8W1^DkR1GzW[pw"tkT,-b*]v-dmDuW?@*yTrA1	m t$:gs;a)B$F:\tHLlmPC#mY5}\nnG/'`W
Y(T@0T:409uZtkY"56A~JnYVhuZ(dDn:W[rJlk<gA.Zi	25&u1$	u>Rr@xK53yq&'emyyyU):J}U\n
mg\5sCH^^u'g)
jOG18ewM_7}].}B]A.z$MBv^@XX9l0Rdnj0y|7s`y>N%;5rpwh1Os)a7NVFD.w.Y6HPZ-l1PE?4el%`uWn:)}^hQbzxgF_6HWNUBh=9RAU&~[:(=h2Rr[D>pyMz'1:HksD}wUJkLN``Y]\^$|qp7_YblT%]2-"$3~hr4E]BI3P$b4_Y;,^X^Yi.Xl>/!i/i0NpF}Z:j	yA;j17OMSeV7G6gn;?2fl+AImrkAajzH(TTr_L"9Uy#Lbt6Hg+~cV89O_C`;;4yHLq&/03FE?3IS7&iTyKS\p>8	6w1kg-K$ptD
DO<VIZ3CGMbwyaJ NVYp&v@E,6)}a5\%%FI&-@z{cf;_%1p,+zq Y_8I3(E"Sesp}3(J+H!<kP]DkX'Q	u{;[t(Z`IlJ}x6-Tj_L:!H>
\X,eQI:yU9;:V165I!N=Y|+4
Vsk+a}dXU<5lHI*peK2Z *86MI,ahBwxoq4LEfC3}iQc
+@%.6_SP<pb	A4^)oSrg%AwaXb1rg8>`rP1s \_
^us9v!VhyYIdWnX+<xCfVGYrD[k?C(ezHv-t%YZ+/N.2"6j(t7e1ATCIh1BF
zN^	PY@T\	2_E5B.G\'+h9h
Z(;25hHJu0X 6HX~/87Xw0vpc=qm7H	!H^V_)og
t>Ad{McC$%g 5jjn]SM|*p[KsF>nXg<
H&%{}7-08S!pUZWR^4	RO#vdANMWJs0,$?<{G\xm"lN":J%TimWk~NrZZ=:,l\?NxW}Q8g]e6N(9H)Z#$]f;OfM|u@LAIR\MM{p	fC>u+kMFS!!%Gt
sV@-L<H[%l'f<HN[Oiw+Dt:U&vo'u gS*=)vY)1|Q+[s`4TO!dU@Xud]eQ(."	.wiS,P2\9hHArkh4M&*d|rGP^s+;u|apHujL=KPC[=+P25-@0V$dtrsR:3: 5g7(7jz:YZ87iV2ZH3'h0a]Dgj=<BxDj{obx6*"M}Y<S+h1!4@~|hKL{WHj3NPIda<AHnYPEiPpS&}{P0%8QeLs;P;1yc`?*[nI9Di;4R>|[wUh}DJb8JflD;%zy9'D7QG,7{*2U[NELE.KMdT&D$F)os#i82s	"kd={
.RI$MET]+a4c=~YjnOacEi79
%TwxFm/<+mK{}R#:Ep#an1"Y$E$,?jhDqQ~XOV0Hs85(c2_l$J]S;$2Q:KN58/6XZk) 1uZ_`t<;!i_GIg'}l:sx!1a~ _W8X!iK&B7|vFWG\lYJM>04mp5p7S>?+
jW+kxjY7I3qM%ogHy>& W0j|d4<D;(&c0<pLYz=oDq35t0/:Yt+^+|N@a+N&~zQwqfDs/zDxkR3B5fTJCB|YZpI]?|6;qG'4-}8KYMZ|R$+&#0!KM4;yA|[Pic@\X,gfeX<_]L(0I:+K1,W}8JD[}xq|--DxbE7a}F=@gbk.&L.	[U52C'J6*6Q=gGOEWj?r]EStRR7u%`ZAk/G0E^ga_$9Wdqa4woy$S~QLRcVI$BIl:UV
qliReP^L{|tc49p2.{@JxF,
XrA?9$B^wu<^='P+,D*	fvXU4-,<C#G^%4=-mA1@0noV6wnoy>\(|f#l6uGLh\f|NyBzl.@Js%m:#&0fm1GhK#%lvb~Tz~ahmGFV/!GQQ!NG}ej{FFa1|>hNR*s-y+mKXm	
=F\OjGR|5MW*2SGC9@&h\IuZf6]n F(w\WI\x^	"YPT\TiWKiS_KM,d$B>)Xfk!L/^PPyHeH*NY#+E;MR@`R5Z\hHw5@pjgofi-{E: :, wbkgjs`*&
sI|iCX8z~aCX09L;dM	(.n?ubb0%~r;,s2 Z[9%gng 6)^qWV3$x!Tes:PDd.](N&[BjOc]fwX<V"2(4prc&aLi[rCyFy2_gnT(N
vi65hg)6g5(u(@4`Dim!P2Cmyx,f#(q7M:vT7c|_1ZFJLUn`hs#7jdl!]-y?JvO=5;=<)yfin3]m/$[AjoJ7<X9H\vco</t?g0PBK)EveU6:Mus'i[y/ ^PY*A.Z!`;F]{8%Z5`ZX/QZFy@hB(V"5N75+/(5>uxoB?1u!Y[12D-g6]*lF CLO}S_n<FH#&}7>%Dm`6tM]hP#C~eC
Y}+/VA.)"bk1CHwjte~|aP&y^>wnR>cYp{2D.Fi-,v4?
a;RNy&h|2?Iosx._D#K"8sX_DJI@1`np3d	YmPV!g=\)rbnAk6\6GR^'SM:B?|n~4/zXr&YcP!czbj]Y1
>vqgtikDcU,w.x~b6&5
;n%sY+.?"]>_Z]r*,0!w><;1yODNVHRv`+mI$!7ceK>[QzjZh;ahX8teRT%@wY4gq\y{>U\,Qgk$}j,R;-K3:gCQ}On_rd*qCL]D;:}|.hLx`Ha|*H\d#P&+]>pl\XNO:O[1yT*R|CYF*(|=JgD55V
%J_Q,
z/d8_mVn^ KV]44[Sv9srG^x]w#`//-WHU3sbp,.^k'CM0pxu|V	+
!UOpd7?@7'e%=Gyu2]TKPB&!iN%P,Cm'I>4[w:34
:c"}Pb3/mL0&{rHYHX0+m[!8~+8&~FCKO{g\wbS^cw#Ei?rZ9	5{_V1m,;Y/Y&$P?1;cf`Ux]+,(Qxx"Abv5`e\};lB^<5V_7+wo	lv4MXKoc&,45OK^W:'bR7Y@EC[CsHn+;=hp
1^+6/\h&Z	l3l03	WG-k0+oNNZs95	eLI?]sf&}X=dE8@i6"OS<sN~Z!\69]$NA(*MQ,t2=-aj1z:>1rRByI)=pS*vy^4Z	-i8A.3u?RH=!(lPzg]M[sATe={sA~r0DXLlRq??dkulMWrU|Rv)jIkmQv-;.aZp;O.Uj9M2|81@mpt?8p|iG=8k}Q"Gsn8<6/CW	Ku+_)"`0QRqf*K6N3DfJs0<*k5aKW=m0%NS:`KAiCNo{],>(kNNm}IH/>t ^Fa{\^qt)FuJeX(a)xI+VP6;no)xz-%Y+Zyk{zEj$:
U)vQ,)L)0?.0	nB&
J/2#c;*o6o}47{=(1CYXk5}Q	ky=D?eF(	R({Omp:bgcf]lya>|NBL1TQ.~Gw?D/}o(NJM6iVr4 ?m>`~#n}g9} i1a^@}LP)	65#/-\hj9*2 >&QF>v'q0N )x^XmaZ!OW,pR'S@XdSqRsQ$3~4l~MCWC>2|vNG?z3@\\Rf7:C+&7x.X?b3-"{G>O(_M%S8FakU(>JN:N2rO%=h6Q6-2;h !%KW|M&./'em0{tpD%"2A}EG*0i!J"'bz>'Pk\Y2gw~T;T[#YIO-ixU[=aM)a(V0G?on>OXGB#'2;h'`1#DCY6}
Q}e<oo~VUgR]N;]BFE5n8@RVLkqkA
;P98}(Re?B,BVWy5X0;Eu(KWpI}w8/q6h=2
j"@&gS)s._<iQD&WzndIc.	Xj6,YXd:!~5_`<	r1#gM-.nrWJE0@Zoh\tAfRo>PRfzJZO_~_y-P1Z~Yn%3|F"1s'K5> `A;K>@e6`W_#Xv*YlyV=HR2bAb8&-7	@(G ~fQZ7h
Mx{<(6^c? %kY?]
SC?aTs^W|z9?v&!w\7q?6YCP2b*2`2,		muKSVyA#&[IetKwG]I|Bemw=Bm&r(.'2.Ga"PfF'=WK	/R(35MJt^=3b&}` (Xifm<K:\+"$<w}p02Sfq<n2Z2nTnF@~$Cu_}C
(jI'L.J:'#z9BH7q"B8$!UYN4zJNF'I:4{%^K}[t>)'u%*};moXJG\XR@dm
*=O'c<'FIe!~q:$FIh)g3w h5Tl<Yfjw	XHV}0tdN{'+_Ep[1fDmynDe$3,MLp$ty@JlcpU7Tk22A~|Pj+.~x<mf#lryj~N#wCg#!yrL>uBUSjs@%Uklsl_Z@Ce}>r/
B8'_a4/-yan6F_mup\k 201"\(FHb0C;J?sQ^i*l/]Mb/c'Ge'!#+6'o&K~Zi_v( 8qj1X'q`BBF]}Y:)\k ^|YvFkC#7oS'<%E~}],QPa..hd+?9ok#-cf|hbF[USPcV)9fPXH4}/O)lFT!H"'-'.?D(t?^GiN9VR]I(2N4'W))e4@&HrMQ_\ sGzAk
U6|Tsj(Rr+*cbAd[wk<L:m%Mx9Ym@|Iv+M0H|ZB>l|3l]7_P8N((Us9J!AM} /H?,%(cKAPmgx6Bz{x7j@
lG`B'(f^oi?7^M|jo0'n Il3C@[[[UU$uVN}H"4Bq1#E5:`xG
QYfzeiJGVkW3
uzUb
{}d(iO&\W$wZxwR%Rh.n3Kni"uH`fN<
{9Bmy{&cS?|&M~J@zzrg:9/j</-;k~0&i-WlIrpd=WB`C'F)Vl@<X=sY+gXlhzx/'0]rVAFMLE_h\-Q	]V9z\^0 '~cqz.tY?x3-"5IBy|Kb62Dx;?[_1p+`"1AeW,(p0{vS5wQQC0Xs0h	cUXrXLbTtCi1~4

FUzYhuR;n2^MR5MmP`u#$PrPRQ`L-ciXrJ0B|\_uL+5K8;bn!|}iv{.%h{YZGmD"U\8[^Kj
3KWpVtk3|#k,E#xp\rkoYO`Eq#'A'r!ez6S+gqo]RPXxiV*(",RsGM|:JxnLb8ZD#lhkhLZ.|^zRQ?,c}n:V_ `x-eQJ}	gk@5bw&LIWCzx
zih% 9f?jmyK*^Qqu{P|M2;@jXB6yp^?ktJMRXzZn25a2}L# L}|UhB[+xpCZv(r 1'fFtGuhsO.vonkgP7(1sE)G&ibf$z|^uNu8&^q5{MD$m6+[}G+OhX5%b7+9~c@yVZ|Vcc;k+J<JK[cA"QfG.?,M;1l6 	QnO>HgPkquRb&5Qg](,E174^cmegprV0!*eni@,D8&>`4TNAR4	sep^IoPG;QuG;m
}	BB&l&*.LiABn|6AV2b^g>CB1wbN70Y,7UHH#Ajc~ $13]=k$@j0&9wu-+q-^o[dl+)vkQ`rrs+H6ZOY?(:a707Wi"?AnO;`iSFVX8EADdY{DK/l6EtQ6qh;|Muf,!Ww+C0dy3Ak!n_X{|X>dal!7gjg,<*5N3kZ%=uz43a}F6M;4>74MAngzbT@F#1NgP3f]Ly
dab5Ok{wBr#z
Uk]iq1E-+(1P6H1T[}42E.iW<GdBiXA,\/Eo]*P'dJ:v':_UAE}P[D?z:0	"vIgxQto[D(M}gzt0Y-VKl\VF}CBmm
D2Lxj
qQp+?k%_]
,IaXc[xqJ(*Sq(X[Ytt" a]05NG9Ex>Kn:{@bW&F>Bl$B;!|RYwXER1:>4r)yrUY(K#r'hmB",)\<v7=eNAWp79|]`GCk*"N^nm<FF%^O8)zbX]VC-@*riiE:S2{I'c#se5Tr1K0@enHg+*rReF0,yBuc\'lo6ASq!OkJ<v>AeumF]D<b&'HZu%}r+rlX\<knsN'XP~k+
@}:ElJ>:S*x,	)X7psE_Qy.|5]igc+YMF+<beq,bL7@q?p}lK{pR7yAml#zSO_.CT$6Q~FBV^M/UozCs#Hv3!ijMv>ml6hM]moV1D13=k?j#r{*.SWW`ZNj-$G^8_d|l36&_Zz)EuYM:wf;kM~(N3/L#W{8y;r3<TRr=:':]CX]AI
,K8\i_7e)9HW!Dz$Pf0177 @2}x-!HG|\9~4,Jc|?gqQr3N{<A1{z,96_"oh:xhF-vB0q9\ E5pL$g=2GP!xb9ff"C16N+KRUo2D)D^Wu5xu?e4ZgRAZ>;0"Vl[p'\9B.2oA%[-2ZAZ}8>2_6q4:x=q PA{_>lt{tNTYBolIL;4b0ICR}>6+Em]D{%Y:i]G!
^(Z9w{G?Xi>;gmZMMQJJ$jdfK"K781@8[H{DZH-Tab Wa^l{|ds{vB0F]/`5wY	(|D%iZKyORS4K99<c)'W$#pY|n'
\r3I*,Y0
ux"K2 DO#?fa#0Er}KVFD0hKW'"^(HXAtXr=>
hm i!2nd}Z-X=/I&$/s%;APgY2bAkX~*M7DY>Mb;aaz@a;Ma\UsW3)y}>>F&$fi{M%3/)tMl{+"3O;	?z_]NbUXWk`W</!f]c93t_t\>{pVm+zg%G6TaN,z'uKq:7^pP!9t5R!,IW#m'#f` Y(E9!+Rh&WEM$U(02s>^hN
V@l[!g':Rd4{KK"Hp
KGERHHD&L)c=?iDL9>@%m^|mYDB;fO d;lSZ ,+|D=08;99u[FXVCHz1}DErV
<A4r7Yy<*!"wn	]oBp-'5`hNl2!I*]CpTul<NQeBI</^JRO^^*B!UAGY^O5Ju|iPO=2jPQStyJGaA$P@F##z1#O*QNT\H4#V(NGv\$EkVuH'
{J$);Qeu:|{-,%eAB An6tN:T{-w3<(\#b_^?BMYZ)Q={`FX)WjSDy1:x#4E<H3$|!pyF@)^afzCU&i-q}2P bGrp	1o#@;"'R+q3-vQ2AQj3c1RZY;#N#O.yU'}>Lz/x%Yj<RiCmT(<3;P?'AgSOC]m<a'~zS=Qpi;ZZ-#Vn7
T.0zv;r@x#tZ;fo
$(L55)lcoF`tO47?ztVx+~<L^}n^5)`RM,g*IVe89aQVC\_f~3BFPn\UI}Hvlm?:.,D;2OvN[Q9(K/HZ%ud{MZkuuRl~@f6D"G`	Om*~'gxP?Rw~O\e:Jdz&`a{`@bN}TK3D?o.:lS	?dyLmhs:3'$9|J
P*JWPrb.\K|6UhY[~[g2TYUh@PCUG`\*>%4$FCbt1njGOVJ0<Y%fNzd.,H*.'6vT3,Hs#x:{<@)- f{~(eBa:seSJ{P5tM~J@PuwYqRgvJN.`gLJH#DEr(-z,*:N\p@SD~Uw{@6^RU^!,GA/,PUgFGKE"7;XK]nwh8-MTCm5uzmc!=}1T$)Ij5no47H|A:WWlIC5\T0IL!TMU_cyWp5Vmj&_!LxSv[^j,U'WGfT`dR~|H0$;+cz^o'0WYZk*o<.5>o\(x'<V'^2=."Y'g+Fl[U)mft%:xOj1:R<cY%]~H]x.RXwp0E>lnZ&G, o*LfI8\Aey2n'Q|4+:'O"(2lhuoM-)J79lPF.>X/h>>C#zF[z4pf *(G-}TMG	{3Je)AkfSf@0hJ,Jn`cYuJ\0z|c2k<]^&M	lp~6tQi{I5sWk\bv5}W16R4AJGhPHf8.U>Xoq~|z !Ov$~C1l*fc7y;\m&ntqkD.U1KC[\(4U*)z[)_yy57M}%w"8	/QrY[A$Dl?VIY/gY_pt1rG32@ %zdwuOouDj`\mHrdBesz#Fh_]0pA8c@>xcy_djMp1b	&]QDrkD\1Bf7qG	.@`P(xKqV+zN8^)i@bvR!`t@uJ{8=Bf}2GpbS5M_F3pcg"eiKswZl$YP%1gaR-kSMBT_=s!o	Lk~1/Lu]DT>d 
No}UmGt?\pJ,gH\bz:G[ro7hzL3BHNJ<q8|iZ1q&F>(S`(.NHAx$Q"D`{9w/< {Sc">s-Y#qt\gr^5TsFQPnB>S%]{aWD $rL"97M7F>xV*4V0^[r_BAueE>?,`:?N41.4|C1=":/\,Wre5iY	"el2/=2*W5ku@=6\E'TP%4;,(x_Da{w\2aP\(
4Ba{kq3z%#cqY&A\ij[UX/(5$ns[$!{i$21wbQJqySoyc$k\GJC#zRaDRg*c^wj"Lmy;m=TZD7t};3vDY,)t_,Bzm+EdOLksFZ85"0xa	@^/d{re+n=p'o]f\#KHh{g$`/IF;v&`##neA>':{:Lv!v{cy9u.Tf~'\P3FGz)||P;jz&z<#8")gLrV:i
NJ`{"pX|JBZ6ytF9V
"TYbKyKwG$Y7
\*ew()G!7;[E38l
@z7STRYF'M-}Yjc\GhT8pN>{#I#qY(qDYMtO>e}[dlRIm~#Pae=4SvE/*gufZD)i'%QJZghruqwWbQ?<hw_|#5OM$6p}Ct% {z
HW=n_d>0Ddg1`m0%)-IQX@L9$z]<g}r>a7n=tF4bF(& W>>e`X"upE$^#Vz(FS*PXeKfO<V)m@?H||Dl%{(g#1$?}]bh	FU%IO>A_DF'*T<Z_cYrOY&O> n"[vU s2?V\BdVfXh
^s3O,A:gFS8p:vrzZ)fSB$(I9
f!MF)#pNr/`n{6d)k]s;z+W$>~<^s^VyP1T-;ug0($Q\2k}dSI`!PR3V0ATKAibvIVAltwNs,rg+{$i 9e|QV\M$i@7TK+9T;BH3,>f9<q[Pasjo/Ne-(0M1`(=VU,!+l+DXR=H@1?HFEyYF1X7Z5!wva4fQodkGPj'BZYzn2d|HC.
sPP^NV)M\KNppT10,g]uLX*=TjyH=Y
mrHZLI67d	icW'/:~U]*0@T"Z2fS?KH4+71V3kG+P?UypEMn@d4y67:E7PW"<q<i6/eigX'.(nxOm?_AnDs[:moGw82S]q-0Ed;T"
//[W$8y9mBZ9<,ERa#{Ax=}[~NZL>|kJl5+:he2tPox^3NP-<ok1*>S*UMhjQL2\9gDD]Y]R<U{SF-XB#DK]-}xbO!>aART./0}wB\gc_+$n.Z"WN[ 3&}dF^r5t6N:c|LH4up5$yct%k)|8a&X [<(UZ8OL|w*,H){xW&[q(NHeqU=k2w@3ER!?K%gH2^~KOJZ2ZixW1OL&2@H*9gPSn{Y|C^>Fq`l7h@H:n9~x
7_ap-e,N/!A3{XYukND\;-xgM0HnUiID!H9S:m}I8aC1cDxQ!jS)f]nNW
b(\/5uUZ;82VZ)9is^1Q	H	Nf/|;1~Jj9L9GzbP	p4DoqV,8wM
.9\N.@~"g4#h&/{!07BmKfN[l?wSOtV+x0mQgQ&RfoHMi;at/Zm<
7)LV2erU:|M<l&7V/e]Fk&P~{w("QzKjB*(U2&(	R*Sws#,K^a/p2QKyXa`GusZ
$Bj0Psq
(P50qVlHy+a<"b#m^\<S	g-P(Sy/(YQ:@Nrf}/mV/@Tx6g~|?G6K.$5?[q|;]hox`
P?|'lP"H)vCm@jN#ZHF'I=awj$S=pC#AeH+f3.XA~eCCyk[Gu?bW8wA6I^iA	sTh}^@"dGLesnlvL/__y]g5u`GIatA/@n_ve/C[ ;*&0TtC2Io;Fr`i:@-"z2IA-N)8<xNmr8qM,`|#*'ww| 0%FLLqL`k|v=:##lWyPl.:!`/,m4NpZcZWxVQDYHho(kxRM=2s?G
G#Vn:yr?9>:jCFVay;J?$M@C1[Rz%RW&t>|3\Z?[-n
ZxrHAJ9/h-{Zr#C9gul%YO32q \H)Nk}c_VL/{wMu;F_@mzPilc!hH~$?JY(!^]7LDt?v="nKT;87p:LoRj{M7yI$>p:G/:p,8		I]U=HqM%;FFS=FK$BYMC&$L|W\C+J;\jR!Sx$+DA~CD$ywCHr=P*qf.["LxSbE+12/OwE<P=X}%D=NY$IIp!/ph_AO%4y"TTA^L2j0y]&<uIc,0@9T(4AQ`22\TJ%#q,McB]j\g?{8p~IUWV=:*I	n`=G7eOCWZU	8acCPhprF3(mYz(	IV_5O)iy
{&{Hlv5U.xTJOHeCHG&X{G;t0Qs02+eVf.;]zqAh$Y(4vqg5CK[Hg59wS8_{hFR"
L]bfGF"XzY\aCKWD`<|T1^wKi(u79
I8fB^vL0Ce~!@Ry27*	*L8"k$kOG\_mFP^@5s|E(?rp>b`5JC!	$xKE\vu":(H9t.1sb?qgi9MNk<.iH^?~ 

L`oE22yqQ0n:g7K/Urc$aE9AUFE)}zeYa}k^G6AP?n[)S=Ujk-kefD]j<wEK}"**%=.B1|cm9a{yx`16; 8xGn^6	)7!_3?e9L]bXNzi\=Wm~XA*6e6d[8*zcfi
WP9^N^6YTb*OMRmJFCOX7&Ne:YfOfD5uB&^]++Wl:z({5~Aq}Z)55}APU?|+yy7!p.^z8OjdjL72&?:ug`*\ivo!A,_-=%uR|:3z#Qmki|VWbh#+_?e'(6Ej]yr&<z?H)bJe':Q;Q+%u6oF_B:ielgq[Jw-#P8[f:jF2 -[dEr_;(9j!	ugYZ5D+hBQ`QA8\!:L!cN6ux;uc=&
	Q4FCl|"&{?U9j[Q6iD!<Y?>gdlkV3RMZAUmkOE7qg>rAym_s<(,K^OaFH'Z2$:v?r:Ve \~l5":}TqCcQ'?1CJ"k`E8]xns7LEOz19Sgb56N/l!ChEjr=cE_>#!xkQ-.ee,GF`{W4]E8
>>+#9a[ v_#SS`
L&)PxRZ&btf9+?KJp'k*PD'lBi?N eRS-)jAYaadvXg[X>'X=^\R$e ^NQR_Jw7CQSJ12r<)0XP|{ZF`=vLLj{z/Mf|$"~kR]E
V5jLL!'FcX12];m=1G+T%Y1Z6bYHs}v+nP?
xePqYOn)wP1Y &wc2"p,@bF+ 'TM\$x}(wWX};st_I:'QJN"HRgfc,y'XnJRPAn}!> wIK<K6g,2LUbV/<~75HGfz3_Ey-Sb.lzkIUS\k_y=xq2dX skd0&UdY)
>1<v'w@hbeLQ74gbbw-`.t
`KGl<~U	t{p 
+;p^!,	SlzA}|;i>:	]B>#quk$m*Nio+HHa(!c4v>(<rYK"Lu%,EOmkr	Lb*_K1 ~kc)"N&u&VpP1URC<yF<a|Pw8'];\`Lt[*e/p'!<F8i6^bVCta^[s5'
/pOj4;'$:bvL\y?-q+2*',R>j/mj'<Bw=Ep";"w6cheO$UhXWI"1K9}`4b}RU"yA[L/t)9kQ~C3:-Q&&*^wq8 fRe:L7A@dh&r-C/d?hX88tHAI<|L%m86.2m"h1g|upstoK*#c596X/lhyCpKpBu/Op']v*(S!8XaGH.m'uz:Odk?heqgkL8-o{ywu4_hIM{':BG\.y DEyJ3!NP&rh{wic>{3.?jEGUZe_h}&YRa{Qr8Wm<1l5Ap~"Hd<q	,9HfzXvl`FMrD[A|!85!uz&c<kcUl0PBn*(FY3Ovcm@.]?pi^%K:Kwp6k!{^:4n6$_i#k6j4US>G|q_%WS\Fo	]F1K3c(Vb]jN9N)M\xi<a=9wWH;<;9Nc.*=-3zD?iK]`6.\s@
&&cZqA'5a&hk$BeB>#u[@#Tlnx-boxpx+5|@%Z'<_mm|Y!l	aR:O#bx-&WWl^n9n>Akt6fBNHenvXY"@:uDQo.Xz`QB*/h>`tz.@:+68,mJdMdBM<lA6`3^T06|dUqC">0mscIxE
luB!z8/Iialw[\}tuqHBg
ywv_F%o4onM\2`Op'5/OI9Wza,Q(dgn_OB($U%N	3OetWnCcb}/Z#&ven6yG`PDBY\kZ"8A6NHgQzZMT<}+KrTD:[rjxQCNO#V0N;+rgS{f^vEDQzi.L/E-B}QQ6DP@a"Tc7S}npQ  RBV.*,1
PwyAPnou]MDQ=.^Q.&^ET#q.0nl:pT<|_<^Div>-zMYj-v<8bNd,T,}`)%~q>7Q	"t_
1YQ#)r*b>.	YU{iZ5Ir&$58BIl;Y	dZ#-v,rB:3@k-{b@n*@*eckx%e9o(;xkoT?|unI,%Q4yln4kON&OhFL[	hqC2&?JV5A59'DTrT!m?hsa0AE%	>SP)A!?Q*!]Y \k,1^GQ]0
,wmRi*]bcEu&'v{:=+tWVZxQ@Hf*05Y V7 ='dgA?XZUu{10?6i/VS,:w}neL#>mnPEu(&A]D !kAjf6)W}ulBvBm Bh8l\uw&xgNik53a;Puu[+2hI1UJL?NZlNeKK<hg\+d^MP=6W&gijc_:=	{:_(?-I?,{w9z<bjg-b{vOf:{77Ua	EGv
NmF#O%n]|pV#cGZ31`FlW' |Hz6$y?q<0m78G
/qtP)f ]jYyh/Tb|pE34[%12Vj&mx>{TZM5y]UEEH;	wM3wT[{I|fkZ6
KdXq|#tCP>=EA7<H]U{}j/Dvtfol3Ty5{3>n8jrni|(dcrP%1_aN?3_Q#Jq7#<.E	*7sR|p<_jIhhB@+QOujx~yD@$5thds&due L627O u8)DUcB.v	?88u;`6:$mk9'?_IKk&C"(s%x~=~.tKOjg%pCO[qY1cj/+DQA6c#u^,/l	qAb	??0
YDyk%&y)AFtXon:9:xD2/9^gc7~:^'@wn;?G%h><.f+Ws7:F<tt)7g2hj`|HHh?)_znwP2[_UR(dEz&{/Ygc/E$,hg$91sre09K.f;|'r6(IV^$c<dmX+aKP;Y$c_n _%j^K]H>S%h'NYm)wFP8Uqh_b(F,\\AZO:sR~wY)_&GalL2q!n5A>=r[oWMwUNDh|]#b CKrdo0ow[v',]x,8:08jkHjZVN,g@c4f"^pDH?f}#TkhNf4 dTs#?V@VOU7C0r%dHSQ&r!^ntAQsQi	J<]Ha_S,9,2FV5/MD:C9VV="F]:LNr#I}(a72!@Wu8!
RH4Zm~}aj[maf<gfTMnTLn!-w'U?DHW9o`5d3ocR?m
!7ayJ-F91,pgaD8$
"@,;$x2{08-C=_,i=)/8>	i
GW8IQ
:`;vqVdQau_3G;4;,
a,47n.`KQC?T)pmF1mmW.)j,n6Zj^b`y[},l+m|&ZW["ji=IGD38T!sicRfq0x:wnq\"<VaXA'UQ345+.Q&m>*\,VErVZL('*Z-Xz:O|X|=m%H1Hjn%\Oez;"0SEi}1sb_lD]pCf=9+\[~TGdwRAtZ5u}HkL\onTF4@g^msUPoUI'G`D;E#^%z>]P)tZpoC[oBT}L`\*;z]3Y/u~!S49DcW		QKfK*h{.#BOvABr_z;"SPUkP&p~|g>cn>KGJrJRm'|J{ zY_[?z,E','"'4
ErS{y2W&
i9+:sd:rRCV:\UKN&N@D{T6\J./`4ns/*[>Sef_R"}A>M	eVA6T0wt23Gb$[W#DU+beP&'@;!~S=;^?c/lfZ*`LvFi1PN/3YvQ~kgU1;ksum/$c.M{v-?93D@UK&>7'd6!BD_42Fp+Fy0jU/a3S'".WyNXk7&P~VdjZ%,wm0*(lR8-B+QwM`\vJEo*PA`R"#%D+~*6.0l>a5<}DblM#YbN|fJnmb=q=;5m[FH_:?"jVqBQ2I\i7Ns0$o_0vjlb6:Yffal4z2q)J25KCt	!tWtG{`y:Kr2"N|``9u.&DdvD4Vt,a'.N,'K<\FK#u4Vf=2V$~5|Ii6j{d	&r$tcX!Y]2ip}t?@MMdwmR|Ml!d`oZX	q]h~2<_MpyF!)1~Sjx`#\tFNH^.0nrGS`Me[AM-$5,lsQA_-
O;"UQmxF3,,qc5a6?U1|C<lp47R=j8i~v$._V[KYW1N6dOS;b|dTwDfOEHh.f*w(Un7kFcU,*/z%S/9!Tj$)<Ro,t;pvI JDHsc)BIkw:1;$)WXsHp*ue://xFF.8j3s?bInb?!ua^)=PiU^p
b
jfA3_OOrB]N:v',`hvXxf@o~1l+wp{!D*?iE.<\R,p0&s_\'rSYAXVxPWTXxns]'s}1,$*B_*8Db"DE1y!B<yM?Ol VO,>gv8
E(rl/',+p~$wmW1FE&-	+tOj]QKxWa(]>*leAo,G?x`qZd5'G6O?Y]0JWZDRI[y5|[}R|$}gfu(b)cT\cw'g:\^5C2`OQr}#vC)>;X1XbnI]"~OCM4]NVSx_&]`4,@3moy"[m QK_rA3hhBQQ)hjWW/x};w|.3Ql^]3GCs[RbRizbF)6&`wGDG\2!%'4xa,Da++}&02zBGKPn=yU4tF%k tqw<Alp}Vv9/<I'@n@Yl8f>2FcaO
7De+* o:PRv^Ir63kKiO%psb UEFHr;+r3.Z`)/~qc+uj[iD`aot'5IfLTa%ito<q)~!\@V+N+AQ#Xhg\5f?P(0t B8977VzB,+iO#ayJH346pc\q`CkI4>d&F["hln \Nfj?a@3FMzy??m->d*R[[u$
uet" 3pX4_^E9?$hFFws0MM}94-t{/8Ej|fM!2.OjPtJTr/[$eedB[abn>z4VU?B<!q^Zu(dz-ELZ<	wX4Jx.GBy8rT)3r5	Y:xV0Nhh_mQc>P*oXFj^BGiz@zqdrez^N3!DZ6]R}ijmr=yrCSv:WlY+?$kf6 +\"YV}"xH3n0!jZTk/pUsz5KM@a`y\vl:e'i40qL$.\X\<:S;[xeYR
0-s ~'$f*2ehLBa
E r:'@QsjsUW=qe$s35l&`dr.JCgz!hbhE9[iLUhU)z<}w+`TV<Be&TU4`kIS~<>Er0z#>]6
JKT`q>?pC)@{=D$SJbhtuxZ#7-w~ENhl2P_ktd]i6lZKSU3a]u; a'V)0hk2 .l@]x/z"Fp/FW0rMaX!T x%[B;d!,(uJ1%hJ0(7:	H#o]EqqD*)rdg6yf3Y9|dNk/$~gN;J7e*#]im]5LH}:&h\9k..tp,CrL4(D:IGbWQEBDqm5+M5?+EuJ=)WV5bFK6)E@02zvM[,OOLUc07Vfvp~p	IL5D](/0t2H!;H_2~RF]/"Ff`/7NP)r-jR=NQJ?mKE_C'uU:lCbYdY)u[[s9h=: o&(czCS2Y?_r	2&39B"D\WQ^z?=fYz43I':_%gV|IBJU,jg5@:cb>M**L^WE`+.BYT3hMNZ?!VHP]tid$rsq H5HPv~#+m$1&(P93\>_	6,oZ5LP/Q\=nK_ECb:*J0mBMd5V!/>Hw7y%;LyPNUB6spq}=p
=g>!R]/3K[zxOR2-KCr-@(YD+v'kv7u1G$/J=_Hky	y8!5#2\<L9ml3oj{2@,9$_xJc'0i~<\B
7VO:vyz8	o_9
gM`01!Pu* XU2h<XK4bNeUuwDlIS|rgsKL}\V*1_e}`_@#?S>-gD3[0:^K)_,d>R+$WAFkPE!jm';B_I5M8~H*fi"o1A\0Ru!5kh3NFAToV}	GDF|<P_7*s<{_G%)lPG.?|=b8rhpurLf>hg\%x0sfyRdF4n#.JJ"Bm%QM7*-'G c%"6qf-0GR4lT(|0oo$dgV.%jzY3\BLt *_xGYk\2Co%s'pl+Ze6Z=veuDhr{n.V2So?4EULUd>v}6he9Z;R)oQ%._'Uv8{F5%=RzrQ0'-[9WD({5WKE1ooGmKvX2}5/9k;@|:ILy RZYd>YEYprUz&;A|5&3WQx1(aeaI>BJ&H6!DvogI\d6_^"%_FuSPWz#L^R1BT oV"g:i t}M.H$b/l~)-oqlm22d(;pttp
q@_fJ/iZ"E+	a-IVj@-LO_LBllguuL<kRUL93r`b3Rb~fJPF.kppf4`PYEMfu;<k3HYeE3FtC9*\MHo_*42dTqm},ym9d52WDlao!a
V<S$c/}K\P1urI~#ndz@L'qinrIR{S_||uB5]@AW;Kck+Rd	`%MwS,$=BEc h#yi4yj;[dKtN'XHGuy]/se48u>HPrDTR(.u(:nR)?B%ON*H'	09ZyE9(|;iTvW%h9o7
c%6k\7Tw0a?]:inHX,:=P|7&#y`e*Gfq	J?n|hv:4l4?hVr%Slgc'3^8d74V,9hFkyl"02%bDJ24j\;OG|bdE!x2LkaOf0S$@e;U(5nzaU0tYTznkK5!"bLj!Y,jTRk5v_Woa'4=*UrPKwyAdayG5r\U[MmuWlI}1Mx|@$!w+!t )|oz:lvfuf1Khv;d,KE1%lT:D%^cIL018"Ko`D3a^xj<P.'0S@E(B9+=aS|:7IyD!<LV!xMA8K>AbcSh^+WVpOP(T	SlV`j]XJceMK;=vq8d3X<N0$3|rY-#8qD-"WPDW5477c~@2] %)R4%0^t2"8,4{ASi:|	id8xy`Q=Xww{5+i4Q|Q[)?<	AN,1`~1p8L2A`irT}VA`MI]{8y__51[r|GdvW3W]{f|*(Sz4IpHDt=Og/	]1l6Tmy{$fs.ld%Vl*_2D2&,ZB"<;P>`]<
<CP)3u5G=!pZieRL*`)9dUG]t^%e~tomb/1_kVFYr)$W	Pvgk%-"T#;NGQ+Ft]	FLPP34IAmRTRfW0C\XtTxo1ER9eK6A}G;	*`?dFs&x8c|N:"z|#%iF
.#[$ *Z>i.AC;vl4Z"19(GO%ne*H7X=so`[8KkP<T2E-]Znkgoj@}L
g)K@AMWWZJue("DZ7'<1z'AY"ba~[*rT_&fb)p"\G999mBQ6[5"=8vrH;27zNQ5{/&g2[C.p2hmJpXH%
u2yu+W|BD;/.rV5^:lpGYo~XMW	8v`gx:Ko\2IN$IHjqSX)@O&4lB`TI/u >v@05GLAD`0{b+<`FLF]XqRiYw $A*M-cM]o+rrNJ_;:p}#D'+Nh,QA1&6BP,}0\1Wzc12#++.2"]V6ce(O2@[v>`sd%Z{3<$3FqBaAwh<uX{qHwmKD
Zl$mkK/^DQ=B&UdnOQ
_"4RYtxv"9aUuokL'.Q(t`=R6-i?d6*H]0^z^X>n`d(5$1GT1a&e4Q+BAh}PRS36+G>f+-%Y9D[
JJ^rLi$kc[Kc*6]#5):vXy"QJ~:Ui7P;6_q?G'7o\k9-i%oN0ly`lp?nPsZ?1PJ}]IJaPf^
NU=_3Lq&JI\YcYcByt3W-j$UECN@KK<@D!m$g-%8Eka{p+8mlydD&'Bj7Q?n6gl-|8`c/8-<Zz`^+6dN!:YiU, 5_a $kIH	nee~X&6b"1R=HRV:"Yc)z#OM~=$k6s1oLBGu_.v6:hk[&>c:*Ks'?J<Lw=
>V0>s@X`$`f%'.4pu(PG3wFmx&rMja(Yei763&Cg
%%k[EfN}F.
7<M0b:LDGH!jM,a'k<3VFY,2@(=FNu#JUrkkG;B1!j($Q/UH6[L U[e7^'Wuf<"t#{Bsg89E-T_.'j_]7daH]%cJI;z-+xkbKvkKL8D(UZou9=9Bf;o$;sNt<pogBfC^]s!sd8buJ4."=;_Vn7=sDsL+1.CJ]n{T-1A?X0Q.K,76NZHq<ezvb2]PqY$KTE`a_L)X9p5(>'lKMcaP^W*UZ|RlQX+5JPL/hE;0G\RRVgMC*"uu7DI#iwc|fR"/]_~,%IIkbWAB D5a}1dRW8JdG4uF!;*nw!kNVZ>B_}MeZ=+L=2N`:)U_*#prCfkg:ox03NmsU)Ror3VXzet|37>=o_S|XRm`e1f_C?=KkPQkyL9~E@fl'>:aV=j@f"*hJyp|9_<i"NuWr.X8&Y@A[s)ROqb^iO,fE*y5=;WLfC	{o+'1hqM$sEi|lur5&bZ>4+E2d*y}&ZAn^?*;@T&&`n= sQYZ.>OLBDgI[\'k5oNC877%U2u;aWjg+J7.,L&G/.E+5@
=/)Tz,Nk25k)lQWY7'[UR<
G=B,8f~Km(*e65&if@iJjh;{xf8QXf?OVx<&|GiNF*\9FXI;.~b'b(v9Muv/{bTxy6HPJo9BDnF8Y3	Y&&ys);PXwORvdT	RJx5=1m	O|Ye;Ek8*9=XBiiMTlM[N`3NUm_K
Eh~ofgCc\("FB6yI~~fhBG@:V6gTwQ-kJC%IGy`$|.I$vl5fgZ<	74zP%pt.EGwGG3>YtXT-?-i, :'(U#BKWJkZlimyZ)us6r+FwmQ'_Jv+k?0aZS P9HIaCTZrHp$7+&IhMhHrNRSj^v'ee}AxJta9SorrwqrUiEH/_Igjf>oz\A~c)PuG2w')Qurx(VF}_A>/X!J bv=f)A+dQ9r>}v86,qnP8j4`}OQcbso7:sKYjzy_>|[cS*"]O
lleFQ(Me
7v6yV8]}|BtPb;]"FfN$"&4NJD.d$ssS,Y4#(r&V_^/7V0H%'x.dvO6d(5?GMM$"wdzWe5M:tmX+$GAw])#Os:Y(r}G\=NBi3S?aIVbjZd!9!Zjm*y/EJ49J+zoe4rOGRQ }AESlw68va^:kdUscV.[^}=O2|D6YRZ	
R<)NYi\/%9Don&3/xCS;"kD5^B%6+rD$_m+w6l	~`GIXmL?rhu=kgj}>
SL{_eKp xodX$'+8]!^6rpY}_'pue4GO-D}x896Ntr	+JhS1qY_g\QdPEnh)|
^pF	d1>u{&k+g1r>;u^.2=Vc!Vnrui_nKJbGz|"\ ,j+V4N&stye~.!jmhP>""Y$0Sd`Kum,%BC6zM[0|Ty']%fR8F=^9TRPk|:1M
jF/
qS*}lr=``#cVlH%2Nrv}**}Di_0]WeNZ%8yg.V;DAV4>"}(\J*2J32'l

/ZWbprb0soXZTv?wIZQ?QIVf63Jg=+G% 0$@dPOn-i32j&f8^su}o[h&cKDk`@[1X:v`EZ1?_QUQYwnE
+&RnFXH2\Qz `jQT=Wnz"9mQ#aYI;F(=CHJyBPb>2PXN<q/#h^4Na11`5Nt!S^t(hBQ[vsRj*~PUBE+k(+dE#?Y&S o)3;TQ8a6DPpXt sDfCN^A1|%"aVl^5Z/-=V?D,w0@&1peLl/W=@hTG8S1@s6&H`.%0(`_);yV:f?=nv|`ZCwKo+~&Yk}{-\as{/1_${,ZyFoOs*q%1=z13q3byj8k]@nz:Y_t&'$AuY%4tYDydu!9Hud	)!<Yaws3q<Bn|%xC%I5m!&8_S)Nc`7j<8*3`dZB$qlF!'+`
p'"zOAl|enKg!y|KZnE+p$T1\8\cfn{*_N#Khyy7$P-&%b0,:hhQu27m`m0C`"hxg0__=h<_"WXILmjvk 0`	9.B.%?-Tiz].QJ2[dZev1[9&reJom3w3@QHR}Lmk3g3f~nt"w=|V_]	IjvA:[oD2q#[{gkG{+!\i]|("CC~n[d	iy92eG<@{G^|h8Hx5DEmZW[1^[\T\ZDKkX]H%vL[~O7m&dmvo<*DA-Uwa"r8lp' NB*G)/:)Wbu}x!KY\c;xDYctdb]<fwp>m&k6ko_`"7IfdI^KP6Ae(Iv%MW}"xog+9HSe~kB' [ySls"R9XEat	BU,
.-Xu=`MuJ2OA.0TpX/v8{td[jsW+gS`dOpvQ{7M8WAG*nJTUF$44OOV)o-h]U%ZI%_]"wmEuJ&?.]]'cz\$%H$i^j &DWzN 4A$pEU*v~[jB\;_4pE;?k,ts)\A-krHUr*wDf2KI]G|`KT/HuOlL4Sl'f&V|O940S}yW^fG_/e:<;ets.qG,/[ZI#cY:HB3^`6
tPA$[T5_|p}?2FTcJ;1Lz'b@w?It@_??A2>tArUy+8.
{|my@nX'!niNZW#gQ$8ed)]om:?Q8^FW!tgv,|P}Vb!z*bEKf<+\_?|7&l~pg7MQxT#hT]x -')]UT%^^&\Ev$/[H{9	eeg{1$Bw6u;k&P#n8NU@VxqYEIE/N$@k6sxQlY!lC]XD1x:Q^2.Fn!SZbM'H5|O(V-p*fpygg7:J#A[rsm^X8c\naib%q#
P,l@B)GX3xUjc,\*=U^?|IP]&<FEL/T9}Hugw+tcTko?a[47+w[n"
Y?8>nYPTN#|alo"kVa+lL/{__t|Xsl[bkW!F{yc	[5cS[AuHX+G7BT>)b7?l4XwbRe1y pbm=&-ayT;=;J=BL%*G/9p/H.%r{Y"I2/kl#Q'lM<J04&~R]fz4jU7cL+eV6LX||:%j{	mZVN`&B2=^a`+qd_k/l916K!m#M:y,V/v)U	{"q1MeSC`
)Br]a[xMc9O"#%4]K\!b1oaLt/hI?iF#<NZGt|(hi9k}N*)CZ8>0ZU,v+s#S[^y&%_\ftq`|!i|[2ZU&&1Bb^	D?B:zrcqP^q|9"/n_xi{M-BgN8P'm2/>nY)tV^\=/vpv?*NOMYp.X:59#]Z/41;:K{V)UPF"C_>ZNW%g~<|jw=}-,kv}t65dBu!Slzq|>0:?
f	]^=%	cn,Kq|
H9 U1Y$OzC-y(f"/8b.C><?Pnkl[pVe=3\A9@]oW'1d9akZ$*^#j2It`UlOf=[CK<[TC|*ee3A3u*kUj7-a\]t dj2u!U1e"@V{pjUHPEMK7yCbz^)npx5R`H:xMB7G`L"CFu@sYu<vrmeN1a:B/!qf6@`:A`v)-Z+ml.&iZ|>sSK~Q@= hYm`@9q+6$PlN</car6f4fyn4NW%Ifcq_Z7"{-uZ$*~'TOJ#O~fp{)CnzaVJ&5dA#K(R?@
Ede{3Um<,Z5_q"&R@#RaVe%]
=>TqbSeGml6_)CG4C<~5eGkw5H4y#!Us,Kv?H!Cc*4lYq>Yy_Wm,	k6"v>y*u=	Mq?[O*3o(1@\'L5qGlB&f|8CNub(q& (,E",hXq!(-s#"SFu&$m0W{Dj*>3B%Y2cr\jn90$O5$KnPB2'RR?,pa&1A<n81pLb|T>n-1
9f]"2hH5l!wDN}3TIXSU9dCiMS,NS_[ncODD\$I
Y36BvE-nS2$C;gl`<6Sh*1SS}?dhw#CH;?Xm|j't\i*7xh+$|XgBDdUXr]=n<(-G3zPPN,hM9NT8[6| %){GgG#cX9$.#B04/Z$9W67\bIquq+mjO x`y,.z.egC!lg("	R,@KQd,e	Ri>?FgTaq<i+i3_!=eWI:l)<L5A}7#YG(J^EXVCMMnMeK.ezc}j)Z %vFREt?NO*4K$-7UQq9Wx|2,!k-N;]52UG8z?df=C1@S0[QwJA(U_34#%<6:Hht*/^%j{d\.ggmCp9C_0JYvm-rk;j9A8eBfol*%q;l7!V_,9c!op@uo/(w/BG
!bzW	V}cpC5~krD>B?H1Sk&'	)/*/in,]z]RSZjt-[}N BFHlG'X*QbZ)~Kw:XL7*(Z/<J;a^Xw@"j }jEEksY0FP'0ty^?=)Hq/M0axC-sIV{n3_\c<:n8H-BXq_n( wti	2B}pTD0WRIVdiH`vsP#yD;x!CKIW>{DS$~.:U&oSAa6?svbS6/P(Dsdn/=9'"0 B+!w,k:-A`_r	?aY!HbKk;LSu#m]"z5@^"XK+D_@!d9Ui|8hJ@9,|#E`re?GERm`E(3;l+\4|M.Y#dKqqt
K0Q;Tf\^o8r
5q@h5'^)d|-cL(qs~~gEjIs44%MT18G]
s?<=x,bNJ]mihrSFDu!ukXco\h3\\)Qn0"X|Sz56i	Ut+"XV~xv9n)y}=tX~N4uV|4RWL+3=3,xqo`Vqz@DM	}GXc,wP]h&H]xs3'K!tz/}(|s?mv[{['>=})=OC!zX_4J+^*BO+1g"@X~F|5miIC%+o0QuNTW
O_+II2{zQ^0%g5y zSb;@@	Oy"4NYBj@ (${*|v9V-AMg'inO=S.LH9<%:v065H{/Q4f.|\0/%TuQMV:bv)Op?tsp<MD4ZH"`X#f.BFJ[wVKnq<@s{0NT?eGD_4?1/,Jlb-1"k$sA1HVeZ9__e&(|4Yc[[G@"@gyt	QWdA$uxZ[PMjw-j B4dQA6Jk^
"}pJN/H5L"3z8_zOtb#oT	TTJE-(GBC}3eftk>WS'ow&#jXZYFtcikf/nG\v	w!P.@Kn/O_w?zISOxioUo9Wc{!AU!V,-6M&pKaMFp8\_zN)v&b9]QAoJr}xL(Z/uTr}3;XaOR?OU:PMI*a'=As~
ey5Fc,:_=];y
uabyC~_N,UNt=nL!4s4m7-%Nt=l>5_zh5<__g2[JG	(cb7]#zC+Fsx+.;gHx_T%+RKrE"J:5"*!"aX~2SGCV-4)(u1z@:{QGTt<x^a3L^b|]n&gOp*o6A\(T:Q2ZW;tqOJN;YEYnJV6wi$f|"Tel[q],9W*]#5n`{A eZ}J{~Q'_zP|5\a^SL[*GG(`8]sRaF!\[KR_)0($^fpXh)=T65T6i;Uo6(\CQ^Ia-^:P|c-\%E|vx=T,qxw2NSS'RNJ(?i55ZPG	V0_a-uKx33\Mef<='1i`'B0VcW:{R%3-E?t4ZnT(hG_dGRAG_h=`<ELj	7._74%}7iZKp>kt}MtGf>!fp .D%qm/?83d@PGUX.y6?
%^b./cPG<vif	-_3ICE0@'/zjnbAcMW*U\(d%zC}\h|:GFCTih:
p4bTY!X_wQS4?>o!Q$._cU:yE.>%l\mLBiY$OEL
	53j%Z|6$[PksNcsc6MYhx;BbKB`^}Q4_qP:-6n+1b[,(&tQHvi|AWm37N6x(U$G`B>'[P+zU[$kq
e4
iI QqI0B%O6`m',Cwfx%zGVO'<>Z"g!	&XZb	wkg[~d54QLG&8cF%!rQnCZl?J'ajelOjaA!"}'/~Z	[{ZGK[yPKf{@5H}Xeh4aPbD:V!$a7FUP5[it9UNa?HJvoejro0Gt>5?<yX[FAU0ALWzMd-<}&-Zd+ {O<~9\sn?"v#S^.Qunq:QD6!p}f7	6xm!I.p-Akxxp&K)%:wS`16Nrxg{%P-q@C;&srQi>Z=M2&Ah8r*4Mel\X=N2t\#<T4n{Pv$ICIGoWz9~4/}RtKckmpPJD>cf#`}{E*rTg7/$GEVX?%Ajl.'|$gi`WM<LEc!-Dcc1RaW^eDMl
Q_vdSA]CY8
gdt3k[I:sJo_?fc"SLvFEQ.,N.B%W=x1;QGkdyI.niX	k61"P_g-@Z"'F/[e2}ht2l,=q47;S0hxAB	]h8vaWv\3seTfs8twFuh+r[ol+STz$l<8+UW8G3m?n0P'!yWqz69pwqC4F6EOp}4b-H~Rz:-o,N&Ng>Z,'*i.h`J5$j<AlXL|[eYK$?NWwbOLd0wz6;OSCdOVR}Oh{.R6'/g|P._?S6Az!c:%0]o^+pGw42{-vI&y+&Z4]p(DaDDl&NUYsY-4DXHn1"C4F;ktt`7EHcvq~mL(,cBs9[G|DfRo&il`zvv+aefAHQToV0nYU`z/ni:c$wChxA~.Na;O_AqCJa4x}tv;W]zE@(CrtwO{#yH\Y<*^T985Zt!`wm3tC
[-%*J?hpt-kO	yglzsX	8*X6mka}rp0<Y&Z*`YtU=6Pk~:F%*UM<2|:0]O+Cs<)O^==^+ZugH2?w 4'aruZ>~E2#&[JuxU/{fw%8DoA8oC&~DV9$m=s)w?xyd#BPlBX`K`|&2~\8')Eyk'h-X	}cgy~\<?/2@'mWj} zIVjlv<E+WE4Zv4-w}t!yNb8.tzkqMl4`/gmMtIv6uZcD>l%C!#4@Uu
5c?^\?+P8oTldt<8;}xAW?q:0}&I#
0w*pF!`cJ-\<(*p;E^n1V%6=dG'o\
GtZC"(Q,Z;)j6|lG$cYW;|t.PNm}c;q	5HP"'*x@T8)wY<},4\H#,)!$Y`KpsO|%EaUDl sm]\'Zt)L>v7I{8$ox%Xq5;?iG3*fLyR0)C4Wcnf;\9}Yfu![K>5J=}0{zKY~[4!N>}?D|(+,L{7-ei!SGx.u^UP@0q<f9iJ/N	w2^|]dOuc{IjZP'(dP;j5jtT/@PfF,:&}~C''^<3rz":6UKCa_
@2jxkS	Cz9~m-!xM|5:>Za}W#SELA4G/BD|QNfsH|D{U0^gUsT?mTB$S'L"7PlmEPbp8:zS	Fe?1o2oDJ"{U"TN1KYL[U-Vxf$O::`8`
%+k/+U[mG;{/N6\ `F+~5DA3R[LFE<xDm$T_hqW}EA2XI.6nzn_wdIoQ*ZHTa-Ce;&:E5:NUxpO8eA53^eIqrVy?eQ9Ikg1IjBv7@nsF2]E]Hm-r^?lmN,2Ic<?2QE`Yg}ExI?){BZInLljf6g{LM?rFP:F}o~xJAeN>x*M~Or,^xQj';LWLM	AR6+\;x?5'5b>	2o<\k.cae(Z*-,uEpq]9NstHl&-0Cn9>y*e@Cj	bzi7URXOoo4Kz^>{!:;SvZeq{@;uVaWzc#e8:^DW%@S'~3V\uqK{wH'zgJ-|#c{p}_$zQ4yxG_1C[IK12zY7yqz6]$^u9ScxY# _o#,,.
$c0j>L$BHA\TN.q=rPLt9:9}gvDwK,A&bpSN<1B'P6zz:2oZx\X\Y&K},
Z9OQ3rSjD+_5.`f,2g2a>JX[N_"_!bv_PWw}R|oSf($1S:X7J	[6`82VL,<6%>#ri$uyMK/L\8v0P,:y2'[!0l/=KjDWe>9\}3N2^7ZTR5AV#Gixs qc0I]u}mP'-
]o{D+B2.6Mg3-WW<-:^8(h2XTvi.U\*C]M GN	#CZK_bD`/(O@h@Jc l`|.Mu
]bzJ
IL48.@ndhOIv6yT	5vOg*8,%,L^`*:Wwewm?vC,([lmP4Ow^Q e#!<tpwPUCrgsl40:VtYF@GcK1 &"	hrAwb"#KlLrjW?c-|;\+~j8qYgp1Pn!;&"3W,Y=u2fArBazce3^VFf'Ejl2a+or tKe3dF+-4pV`E6^KjP52@;$)r}k%frMi-rj`y.wEKyj{v]MK~NP^:lyQt,SiF8XoblBvImv/B ru%wESQ-m?iPF<}HC:(I)xC488Yt2"OdIkCfHFAeHX-vc H0>D:_`T^$z}"']}$ZF*GY;_Po5X3)}^+<OEKE$wh<kXDUL'=_=s^j=ea/b<W3+SaO5h)Q$"KjX3Jr2I>|0Tb^sM&QA''/-DH[\~>AJbb`{|8DTavuTz.,'{B-	cq16lX~VWl5zeAjQ.0.L\6giD/5YTV.1,P7]rFqXUG6L=5\j3TtU$an`-#YfZmyVo\=IZG/wm?.^XEMN{x$4lBjC=tD^QX<{YHhM;g9(^N!O(d>#E51LvItT/BaFPLl$MkY!qs{Z-<w{w!}r	mO>d|kR,c16-u {_SM[IE@T{[9LUEc'v(.EH 	I96~Ud~6'}HILCi/sv`	_Z?{wNhZhZ[Mi{"-*qB`vT!ipMNTjYgp@s|v
rK5{e)f{3Wa~Fjvqz3koK9P^,<XHp>F@?
r"G5VRN2/qa8mJ<T+XVACdS,l`*jJLHw>y~m`{IaA#4}k2M_'"irK#pg"i|fQ_zRURh-KNs?D<NX_ >^\EC"q}sEOv[gC:;*V]MS<[S-|sB["RvdLCaY/(=@$0[a'? A*w(E;plN[jj81shj*m"lr<oS-drY/D'k_XTp|=1ui'+4uY*K2L>#fxgfJ0*az<o*(ki(PFryx>XVJ)Cm,QnI# 3Lz>sG/~l\X.<IRX.ec8u\J{7i$ScG6ADG ?)w$bC`F9D4B9'EFG0(&(,+>crAj/*wkf'nq#X_*#r>f!LoF 0\q~9Or!E_u`c[^*;$xH.0GwfYbR*.+,bvtFT>vi6Df>_*^#q@S9	<y9:y.)=\kBmN\dp:~Dv-Id53SKIMPCb<JxJD	+nNH@vn'a:gnEp	NLiA\@78hr=Y~'<RdZR5,*=A-	O+#'>7=DJ\^}G+/;W5pVg-NTr#j1L'5;."EAg#D"Yd4sXhdv>%hK^<bqv	h?cv4"L3?2q6T@YTBL.q%e)h+rmOKzM	SLmmy"%&MWExW^#M<%|Id\`c"'aCtY2xv%FKe8QwDfr,"e2CxGB2iwMsYn7pkJ#muF5S@Dw<
8aRSnW;4IcjQ}.hGuEaXR@M'-1jcfu.QIN{(QrjG^@`W U*b}LiWPOzG_	>yw6,kFRet<^p*SC?-#xThs ?[YXfT7h`T3GRuVUS ^%u%xD.WLp"_OB,m%[f%33{+Vy-rejM
Wf,J{)+7vYn[m}]<(PvJ4%Qwe{=5f?
'Lc,N4VdA5<UW&UcP}tZyr8,[&w;g"/Ue.DTg<iX<a$zdpnC>z 6j	,e-Dd)^].;'D%gD}xCR~C0V\EL+Ef:(dVxUcdO+CZcZzn=H|!TYs<OGgc\IP^YNTW-\TV!J(Kw@(M%qBY;7`.SdA,#O\A'h=z@3Tq!mYv$9=Mu[o!7^G|Qw:
G=!/JQ_Aka(PQf^+!jU0`HB6O>vNF@9A(qR=:4sbt>j~x:&1N]rI#,N)9<;=k,oxoxrD#"z`y`Pf1.kG#;W'1&S~]&x&H'{]=V?hs#h@<R_eakPNV+kA$K.YX3P@\M]%hR-jb|4g%kI=3buQ:#`:Pu3Bd=vlc,EU?84D6[	+0YB<Z=4|Rwmm!I\iT=.2(mF`_cys2p`d5w63VLE.j<z-`R*l1;+Ksnid_#j%Y:}*SDWp%'=)'U&p:g	{7}& <?y,]vPfsJ%wz%Sym44B;r. yg{ewWOt+|=4!jr4/
.&ZjY8'f+>>Wqu4~4LZ	_S@>^n,6]Z,..X7i|$c&ZeBF1b]r1Iu6gs,>H?82%5z26S%o@mXT
(sM$h#5B@jrI8"Ke{j;k~YLI<EL0K#{x,Yv<!5@>xa52574.de9X7G} Uh$_.OStX\[2\Bobgq\Lma[:FMCjW'.`Z(?W2AK	:-?`Gf>%;aQ".)7]v	p>K*OJ<On!(
RU0#lnmq*tu2mW}#,jZwSd[-^$KRm%K])u+c?+PYL8dU	0#Kub0K7~CW!{H-ln6r^%<F\UD4'Hf?MS)]iXAGn4j4d3;2DV`pn%>
<MxK'461GXs6A0E!XL@6;_
;yo)Uf,?`T@WAElY%'^k=}OZoG2S*K8LCP~cMR~D-'::@!whZt\0A~T!';UU%#ul `v0Q	`#pTB4fVB*Ok/I$z](JB`w1UQ:7eIiVUw/+6Bl	&=T;i}zy;;{an_4Pndx@A,oO-FS~F,X"[@2y'$x>%t}`.d}L9a`)Z,	QXW5+]'S_vvmv@qrAV~c?)J)Nt.{lXfdX+J>GC78C|JSR@DU)SeK+VDjO+wc,8{<mJn_>g;RJ>nQ-i=b#b1yr7F*6=36*qW(*>vEA#ds'c\c	sQV/k/#fb7^O6;99pF|g#*.%!(u@7&6 d?*|Z;pY\52a_.2_$QRVIdm.GvU	G[MEx|&.e8$4Sm+!|c3:@n#P+*~XKHQcZ?c.!+V5]Z}\~)A](43tH~hH#)_kqMN-*(WyQ?y<u%>Y]OR3\ht~th?Hq'=U~)s8M$&/66-	[H9;fCH's]BW32V7we5jM/9MReQ<^/ q80esm'G.8)-88ZXldd+'dPAQc_0^FD-ObQo+nLAHRM04a8Q/)>5;	*9<*Y+R$8i j|^'zFNu*l6qi,WG\>2LAjeoG&F_*I{OmgNjI4vq9jFE}!@p0tZjrFqw\w"z~/@,"buo`TG!Ut4.N`e* @T"ZdK|,A&94w{|Nm/DxBQl.$~M0>6[G%cP$oZg,bKkscV|OA,N)2"?x5gs!i0|qP	n@.cbC26eMt_zSFAy<S{i[*bER]=\bU
Zy&!Gr_H"a9Fqkg6HQzZrY;"i0<iFI@0/XM;!M^k^3j
6`aX FJF4Xh.#8:uqqUEcz"
9YUVM9hIh%/!Vq|c~Y5;^k~Y;SGbJ^`k(|{*M,vlO?uykIYh'~'XZUfsiQB9IA	k3C;KF~_,O ;_l$c=![t$j=b=w_oDnc.Q<--5,_tKp>!&J:;Yb@@y_{	7QU%)_N1~-P9:bHuoADWYDo>y2IN	Xuz&5>GSK{Ld31UEB>qw=Ql(BRx//+4fRwbSe6$TW(Oqo1MyhbtZ>	Nrd	LEAZUbx[ZD=#j4^L'sj/,]0M((NzVr~Z%Hq1m/X]>Q{=O_Zd^RalK#6l"2Sw-aXX-W3'f/]1QH]U<"dH2[SUeEXlR)n]t9VJ6}7>3VI<Y@Ypb]]JF"z=f$/2plBsd&"XA- O@T1
cwy3"$.Uh"unI z{i	5rASM(9O#lIdk#]^8_ q1 J2la7nJ4M2|3h"U-Z6@T]).|z',8r~9%1**x_uoD4/.5r]cDEQ4pSpsfa5J
8NQzVR=4{NR1`(z'`a^`^=o~mX35YK}g"z&7pHE.tK}&/0,VIqB*qHB$,Y?{K6#zWB}Y#5nC/ryINoq|(>'c6?yNl!b{I{kb=;(}b(.Geos{s[Hin*7ET_K_g@nm|yGNWPy;@3LOS>2bLSiImCFxSC9luSFQE7vex}_y,e&O8g&;,*7-ef7x-/MR_aK&SCy9Ahp:!LG`?D;+aeqr-d3WFt=JWTb8OMfeP(8z6NW)v#n'pcXT/yw^t"'Zl'^fdKtm~
A7Vqsvv[Mx	-=\	6H=Z|ETdjK4VM4t[%:0Q+:LK"(K4eGIrZ U`r0!%dyvK=O}{Ml9O\"m[BL! sZt0)444%1+n\$K]|z~?yB n<5["L!f,MSL8I&FKx-Cvr}Fg>b_-keK#3u^fwa4.h3.q:KL^kTPW>5Q/3'if!$4 DqjI/linZYvYl-f)N59#BK^4p}jdY\k25[$&`'rSkV&zo1|Ik,t;fEX}Kp4f%-atA>3n\@v>Mb}y:/_M	./+ie"Av{v
>]<#64l#W=C((V(m(.>Kx9'\}f9e9r)GB BCc,tVm|z=SI!P^])t"HF|a+~7CM6P1KoGAbKZ.CbX5 V?.Fq7OF{vWoeJB.}MSZ~\Z6nBFPyBM$wkX#5Fd+3\sa*;y6Z>
}#+Oq*tDdvUVoO$x%v)%Y`Jxl)4+MYucaB4;{g#a}vXLf+8]$L$u45L+EzxF?W-CIeM0F%hy\/4#:%*f?F<}j;6_Rwye%C%w[$LetNJR9s:&!H-1sfhR1r;|XZ]CX)9SVtS	(.sts9l"#@8$egO' m9GX"X_5c]QoQ|#n
5tu ~ja;*4ZO	5aN$Q?LDMs::5L([AU!uzFzG>U1"'
9
Gc(YCYMzh)xjL}_<aGERAF{:]8@7XV@GRvO&M( f.P8>G3OiW:t=eiwK'gmp*Qv);b	VX9K.IaI>d$<i&J}F9d;[&pTa\]Ap<XWW+tD	s(&BN,$0RG8&0*ZJw+plt@IvaCt4i=G	ArdR"D<^%`|2F8J4/=kMcCp>P
s?6^}^M,_//@9L))8tI0l %kr">d,K}Tr*qur51M9Ljl%hS[Yk;dd?o3^PJ5ZUhT.Fp"XD"8n2Vc0Lc'2kE}BPV\
|:brm/xhS50mm ?5|nKt
<zscHdm6L?@e#:P*M{O~=x;B|.px0\IetOuN>ll:*r60NrY[;$e?WH8QE2
izlEHle_<C63dCp(9$;rG989Oz$q8'8,
mq-DLg4	RYXk!UDnn*85Tz"@53Lz("0=Cg?G/GCd4M!xqgmz$NP{c)>?H:[hSI,NL?]`*9	Jg8_}z^MOxdvj&kk\5D0TK*D~B!Y1F{Q9`D9dtW)m=A2&(f p:WsWYqVz$us]g1uzi/t(u[&<ks6=Br:W$4
!jRDXp|C+c?zx8O t'Eo&1<M]>%-@L=eay
)UViN~%7@ Sgd/F*wsTRlnFS&Q,9AtnY'FC&OaDhFyAPo+6[Ij,)eE]Q_K`pzqpNja$qsL
_XP6w"@UIt#iwUMkG0o}h Mu)'1IK#?iL~NI_,tVW`&B1BT!7(z>bo)H=s?]*+kq%[2SQsXs|Y5F8+E7~K2rIG8L?/#q&Tsoi}H$pd^s42	J)9jR+0F$;Q-v*IVtKxfHlqGQsL0O}t[wNd	GxX's7XL0|QX=sn(gi99f=#*{O:,l<ET=jns:w,!mh`^q
$8>tKdNo46(L6MRnx:J;CBPVN3*#,p5UG=ec+,n{j|^#UfBX
]V6?-0|\j<|iqW9DHc,8Mu)SIRjf?s+y4`vlN?n':M65xeBZp.gyTkX97s
(Un<rSJYR=G2[IMS7K+#j]S6ZJd=\m{0D)COD-BA.W]4~'BKvLxr{>L< Z>iU*L:W{{@]bmac?r~;"6/L?2/2:=UnPt=#>AHjwx:CAz8wdsdc\gj_@u!
FLpTjGA'O}(-f/FZ-&' mS2Dw|^sQ._>qq+QlK2x18y:_qdSfJ{sQoYM%&/.B
D1g9@s,C)ebBhvMD"2zOH/T_0vR0kprY" xeB/|C[T,!t#'BQ	o9Y	Dn16iOj5t0I*xc!kZ9QG|%j)n2['?O=}LgW;7~`v_GW`r:_<!]Y"bv9e4gqge @!2>SS(	9MW*t-5H>WD]^BzsZR=E~y{eV>=B1+l1#k{#!S;)-F.yS
r[/7fD@8gHBWS3_;owy'=Z% Yk` WH/<d{=S0J)Ok:oi84iae
^r'"Esm`}uY%=>6u{e3B!AE"9pR~vJgO>EX>:bkq%I)CA$Uz"6 `,Jr}J1Pq0MaGrN=@^]*<tbb4j^ze]n~_sv:kv;h"0&B/P,
RKDG-3"$Ik\+)*q-732R6K9Q_!
K3.f;['AKX=vMG2!sCMY{R2"u1e*MC/
;T@dSCXJHrWuX|(E^}]8nISrEY2W@{*WE	}wN9C^TbFE,+i0o:$t*GJb^tk]&x^x|p9uc~r1a#|qtP:]D3EPz dx^B}wQ:	:b4xcPRI56-^7u?*^C+qihf$mo;f9V[V!mI@%0cgUpYstu?1`vg9(tAO\nIW|AI_Z3#q45Wod'Ht0gVg|=.+%j	W]elNIbPTt`)"?|OWay/?>Xg@jm<S_q2Cnk	K/_OR
Xa -\AvnA7XR+7O8X$Rv`i#i&<ol|Kqz	G:{8WHCsFirnod,ct;(gu1EpyGL/J-kbT6MCl>h>>_Ra?d=M[IJlcct7r{V2.egk0&o+G,"u#i,M@?b E1C$2'x%'!:1WQ%Fe.nX}~5.+'"	0'+mV[IV)M!3>[(M>%i0,NVf_k7G]HcVNG}i	[uD M!%	p<IKn}@l=?YuuY$mE@itLX'`Oo);%tEDC;xGfY u0b}8=-XQ$M/kN'OO>?o9p36H;B<IDn.h9&-(=kejC`HH7E9~aH?|Ve	1EO}wH;!&Q.W]z;4XTeJm8qL%^Co]#(}iFawqE+@x T<xe5Ro{<`y@ +)nG'3CQO<0D.({Om/002= 8.a`V8Rg;xE/1e:L}5O=YH/&U1,dl<E%O#!}2]Rz1POf8AR})Xp8*m|o3lW6#<m99b5R}5X!->Aq+<[
yEX#hb]nS3]n$q{VL+xp~GKlimRM[J[,_<Mtc)\gA	twGTIDw1[}q-M^1NeB4vZHhdx#^{F;0qw
buTcGN>9aC+:? TpW^W&NBVafyU=Z]PBn-z[s{-t,*<;-L!B)<E^0KEy|-JjRj+piA&v,>=#~.SgR_LOREb/fp[AB+_e)lP(RzxW_pAu[1*cxaJ8)%sKw11(Rr.FM@f*{siCmW"bWb^VlaL+`0IBbt/B")}	>'O  B#/<?@<b0O*nN-YeXgA/$qG3,oh!Uxri
}@Qu#iX7nX,BX3[j@rTv0].J%TkV`Q7ML#|~ERW=Dc{Sa TUE$9-zA+k4T6Tf2/Ft)OO\4%3+U/F7B:$tkWl:&_B3B7V4z8Pd%^wX`-Y5!kk.=@
dSYYiZch^s-HJfbbe7V
GO+%g'<Q-Yyf];>t5pa^,a$(B(c{_^0"|B33@I0 g!F$G$V!/.O5OFg4NAQ[&31Ap2@;Ec`q!DROt%,B#l42PZrF]nf4u3Z.^B_rDU[hY+K-bz_!!@D/\@ZT !Hg'{UC
v~OP rh)7.Gl&<NA7+YUaL)'~Bf*VTor&kzH40hjQBg^j'ng?={!KK~wFHy?crdSPm4P>OFcuJegcq$I*iCyWIbqa!N5)A`,SzJ Tg*@Px-LbesM{Y
nZ$~#J7Mo]UgL7\;o%W"R|y`cADD}MO^plN)5D
A`G2,yBjC9AybQD4p	`TzAdec\;KW%47or&^f\nUwU_|7`7M{$b}z-	.AvE~\<vB^aF8"L5! S
AoA;$l>i$;K=Z-.,%4HFqL4,s][La}OKyC08rr(-
u>NN9Wjuy3'q1MS29/*N4Oyz/D?+1S%7NW,\R)fO:Z:Kol	}dg	y/wgh..S ).B +xD:WmzHdkA#E9yJQb+9L(;"fYFsz^Fl[scZ0y|K-Hi"
HE5POf=43.	 4HQQ!]icI,iIp#1d4YY0[@<85#?`P
w0HAt6XD^ |W)O|esP+h5n{tj+[e?O5X8`a@jjbb%NH|_9EYLMu
oU"9Qc.Ny\ Y8zs|>Ym[~f"ewz2xbW/mmxM<%1tw$MB75-FLc:W`$D0TK\vYk$inu0%-H+:X|`R?h1'3y8mwz+v<0Z>gJ#k9DR|"b>j>anfpAkmgJr4_f-Q@O;?f}&O`{6dzX88Gl>xQs i28/d4!8D7@aVxtCwS$vxA]$-{Vg2.e]KP5AWR)
F=]^7*mXY.a#`+Yb)!D)p(L>7z$vn~wr#B*1Pot#'q5[^l[Joyf)xEG,;%J:s6}kbVjZ2T!R?<Cp>x'x?2{]i6dbwmZDg}kA_RPHK'_M	LbD.5q%	"2p0ng_WU%m:$3EM,6`s	7=TKkxpj6ApB'1OODKex0*\`vx*0UUQdMDM):8|O\uQqK}q9k7CKe}l;\yqm>s0~gBkDJTwHK qnq&bQ;J&nv:@.\I@u^:4\SgOoufTBZUxVy=_W@cW{~~dyp[ojqnK/u%%r,)j%K8#g4]m?eB9v&p~	]GmF~ACxs]TURoSdSI0D	xWR9vRqw0Rao]o!<NnJ5IHnoCRW*dM_C{!c3z_%=%_&@\uVx(U7@3Sr*1JH~%y?~+'e@4sjcR(#[;V,[b=%l<i%g};Ozi \C.j6R-6Y?1/aK(9R`	wwYZ7t9xA#T`%hn<R_N7%|dH5u8.W45hqY)6 v}*-oc1\bn0w`knw+Hs9SbAV:z00<W(}1EB@i_:[C4rVV@!6~&F"JVezvf5_[K[KPV/N@Ji:BBf{DeTBqR$t>/t1;U|s\^<l@<ld|e|BDB6.+Tmz%qe1Fyt0:ObPg8S?Vgb]oj	u`")P0JLDv~c
B2)d$9*A71Ti4Css7E us443ff	0YS,@f4=yRQjh1!cZ 0='w"U8E6Ii&[Y?Fz>|H7<[v2~_"~5iGt]d!k~?rnT.W{Rl?W}f]B?
L))`-Z{n7XSvltp.'A^\Hb<c<7<Y/vB>5*x5z6W[b[<lwWM6bD

C\6vXR^"U0gyK:nPH,LVfcX/\u-B,#f)P^vszkA@sjY=}tcKLAR]h%=:^q)"83Us
BF)am/,t5|[wicMLvcd7Yddjmm|lMy"Yu!V0%gFO`eue;bo<1:zDy%7/}Za'R)0my-@Xvsn}FF/ZEb}3xnBeSYl1>p#/05A\\XBHYfMf3=^+|GRA4s$HCCdKdtw?Q79/m9FiK'$U)L`M!Fjp=MYsF!@T3{Xg"-AxKB\S*nVnD[ICY^b#%k])bQw,xk;mc][9[k5A*J&3 P3e1J^Wzb=?;T~rjtc+696 8E$r|s[#?TA#~Wc6)Q#&9O@l\Bh'OH:Hl65co2XXNcN]ssYl(qK^)y'V3TpGBDwGN)0<<,H	?0!llS7=]DHig\9'SNe9QVDK!u^~8~|U[fDU;,T5k;;7l:;^pwuT0;ksC-c]@O+wDjq,iR8h8TJ45S&[qW>. ,`W-R7D$9!RA xYcAa8tM%@-MJAM%Bh+^#wZFO:,V&q'!o|w~w6?(-PHc%FsED*br2+	p\/0<[-7xZ~/C#9	zW,YGT$fD1#ug,M:la0(t4
&UVnt(5H5mZ&@GfZUq4;aeoC	=Y'ypFn$sk?+SzL&9.yxHczVn0e&mtu@/eb
Zi@P!W-5^(Fh:H<UHD?oKFo.tbka#|wy	Ns5F>2ld%(tpM!^e5A,QH[LuZ/rWJ5~]t3Mi/LfP1u64B]LC=xN<!=.z_aPiHH3L_t?,}X	v.HwMMl6UwG(oR00'&dofy#s7Q84i*yUROgJ	<--Qs'MM;#rPmg]&~Fhc!DrZ9_FNC'(g3#Qv*X4F#?}ycW6V:{*3LK6Y?
vEfo:H0F} >h0o#CrjJ(GAWq.B\#z'Le2%RJa]r2I2~5["GbLI
V&6&>%vV#xQ(9!(7Dwx7Dl:36V|MOrnM4t9lGu^dN%!oUj\38\
l23q>3p
JsB)>JZ<PM?o4hk/3cZP gV>$zWmoi7@;q2MpvtGR3`z7E!S:3!2;&KJ"T;-1uxSkqgxjf2U{j/<I/thL
nLc+Q	P{6L#TQfB(MK D`QCU*Cx8.1=S	{cI!V=ToN-^FjkuG9Z!heD"+DNTi2_)USyPm{IOHJgR8}RC4P)#zXGkNt.):nWlIz)_9JUm#RXr<pIx1%?zVa\Iml
+cYO2!B>3R[e`a0.r7OM'is'EO:HY*f)Ufebhwv}/N(j,9cUF`c{*]TVdgT_M6eU)w6<fh(Q	y`JPk$OG5`2LgyE5kAplJYYe]TCu
hN=d(S&tgPU@La5:_R|d|7h9W^U|hH[~b'*l{G,2 Nj}&KJ&B^w$+=
"H?n;d^a|6J%>+75UQz}EbR}^?OF;%PExVK)C>	QsV/{R;SUYLee6\id:"Xg/^87L"1zi"&{\ 1tNEj9?6BT}KLs%z5~e*>M9QSSw]C5ZgHEQFPU9qZF>-a,,FE\S4Vo<"Nm>*N{*K&!,O_;Tz	<-%FZpn)7Y+RYkjmhMOAn-#T[zg`XaPD1q(],=8d+K$i\phc{c'C@<Lc&N|{*1I"88~"i6/w*)B>[Lj2\I3.V0(
zJSNB95UG+MQvc&AqamRvNsD'	3dRK5XS0uj&{3	n*{Az(jN<CHl&" #FNx?~Ad)'6ds#v-"N[
OTt/)y2Vrw}tX,Lgr6^|fW]	*\_uWd'"R>2E-;\K#f%.Vu>^<]=R\u;=(pNUp&8^NlZu*Gx#5Y\+5!-=}":WH+D:UK#nmntMRA&$M.R|)a59cO.)#kZ&-3ZE>#S_odQ	0&Ei5M%/5t|7j>Dc+y`jiV2gw{v )2\Fj3xjTF;[eAo2`YH	oA%gk$qXT}Y\1BAFl4-Fme*b	'*?CdQ5,+c)=#cq^6`nh!Pq9aMg/ODuMKy.eS)EResF/ deO/; >_;TPSz{(Ni8Kb=s}e\hV&wzmFMjZX'F0^i21lOz(%MFcNzDXS	HsT$"4s5I4RcP]_jQ?"mGZ.Ks1rgXl0'5l<B_"GHksIE1LtjnB(t|RREY0ts]|kedf%Y y1. Xw{n2xdKB,Ekdx=|5Ic5QI<zl]Htvao#zw}/y3,h0Va/TO>}ck|V&
s;"dBy&;`@8j9bel?mA~OgZgJ.f6)d9~*;u6
=U?d0f=he7P^	\Rtu|gf5A6DM]6z$2%VRWBjy<	GHfQtNNPJ?=*ez	XUb?8	x<u6M]y(@|kj@;38`)ti6`@A7oH*Zep"1^4\;.U!EQ}5NHLIay*:+=jF)!j U}^q.EdkkYh	N>ZcxDBO|]E `"h6S%iqj^"7|wfeq%2K|nlc(-[P!Vc82iBt/cS5U\;eG(U8mE|>6g<yp4sp5RQ1Mw8x}f)
7xt!3V^NT&:Yi@t+Q-m!5_{m|w@x'F/&PW^#TfYNH~2dBbsTS{N]&v4GgRKY^p[]1AS2"U2fjzpI]|bfeTh>sdmRi^rbfkE"[ c/CZnNI|DlPD\8Hi&E#l@S{![_[.wG{!oM{U5vK zJD@B}AV6fGVpY58Z<kh5syBcnm_&:sZ[5`IEyQhEi>c(!!ZPN\lF.%3%tXUH_|Ju(-}XFRu;U=kb;nxaRg!rxIj4m$]8}?,VaMNZ<;B5}gD(wfQ_d+wT_K]kDdxg;UC/N5f)Fv58p&4R3~2a~SC~Yn6~=LWC~sp=  kKx&Hwl>8>OHgX~e(WCEQLA#in`Qb"h^d]k~4K0eO%]c@p,~3EK)u,<r7[7AKO unFp+z7]|>	VN(Q8}n81:`6gw9GY}X8zh:82[b!'-C#9q&^xM=K=C:>>{#Cmzn%u;*t06CdlA	VimjsI(3Nzt+E3Ed2"Ck]HM8:K|4wqz`\Pmhy`=!3>]b(:[};l!oSm,!XR;Wh%{?qfRDnu`*6|~|AY6Ub	!hJB<U4f\Mqzy7-3zedGh\sz\mBS&X0RAfQP&
P2cIp({*qhjY}PEl*N#"F	:z!U'}Ebuw.'t9F$
5bybO1{?o!f^)|K>i6>RSt;+A62rc{:9r?.,jT
V\#zFPWKLCqrXFz})OEN+H0*G-{8zrR%DB-/:W:X~ogapMd|ph|h	j,r:r!)*#
LcW$4MVG!"\sK2sNyZ.^{%[#0N"qvD3bzV#=HZ'j(,OvGnEya&{*@$h=_{+^1(5RG$""[CShxt0@wo2nFu!-!`FkDL oE8b+=_cpJ@G^!}bua|v|Cl,U!f1l	[OWMrXp7P?37G@]u:7	4NvTzB}UmE/Ki{A=z4[/[tjxN\X	zz6+4Icmg{UXz"a27}DlIZ`k[sl)tZH@SjfKhj=-!0!~IPrgi&J!o}B66;(kbm4{WE L}(9]-k!dFScG'O`f!I\oRbeg;`SJ	r5b"x@Xn9 dlxf~v2&r^7HJPu-]dFn'9,NPQ*vGcvW&a8KxY6{fHKj(-uXPgh?z/64QQc|BYHKg}\#VI,*)xz0^B*$pD}M9SCX.UVxE|n}1okV.OrQ
^7R'"U1Rw0hwN3^ygUn^@Jd_*YS7x|<{yuNT28Iz\<P[8kK6R{2.NO,gc^!j_A3lRd(Zrs^f;cQi>#-
R}RWs+&}EmF&z
2yX"f]V'@0:Qj~#^G/l3Aul"OJQr=%J)_=q:K*bKn]$+t.I3?:0dMH	}i2^H0jYpDES12[x]5ta}gEw"v3nzBL$|\e.{Ur/e*\U3B6A ]11Y@7e|4M"(Sh~"h<ixT(0Q4gz#]7t.9>sGwa6halm#O1f;y"4^RFQMd_sy1JC(S#8}cl6-cG]n\5d@X<olxnj.{R#&aAQ{[V>b~hRr` -$l%e 5+I\[`	ni)fymvEsQ<B4ovf	dV%G3	YA2:!WRl_ v/KzNt6CykIBXZjdrw1 [Ng<ZW`hJ.TW
Ts>v{0V}fA[&+/D[
:V-vnv`'{QvN3`h,#H@V1N"m&3([?mhV+A"7&Oo6~%q"!j"F?hRs&nut{[wa!"{y7Qf	/Z\}qO`YawRvp&a)	Pwj`qID\K$ZK[,XRC|ghZH"F.D@
TCwoep`o//&<E!+H:>Jdq8G,TkhdXAXGI\*7mh@3#KqWv.O'.-[`ptAH?Uz=ep!&*]G%B6<v><I{g&Ppm*F-dl<7R-h"4>$(Xyh_c{*0"r
X{Nt6Y}`H*gl~fo&CsBJWu!FHo+uo}agR4?c3*!,n*NFVbw9FY&Lm(jH|1M9uIYT]%GFmf[qa^Ct;)	LNK"[Qh9	>*6.80ACoIw!:n\@-XRF$meB9z9Tx_Rn),kO6\Q34bjiKo6@.Ha^!'HlM"Lj%M)!liL6JG4l)g;QGEo8NWw`tc)Bte2hj.iRxORA342D0H|q):^gN'pPL]n2sLT90@oV%AoLdqCWgU4q{;WKI|fk;$@.bt&VC{on?jGSwwv0wz6l?Si\5ez&%A>}ipj&2Kwkxe3R[A`>T5$l{K=FnN#zIW5nKlA(z#4ci~,bV%9\`,<+QP-{[>~0H-{4/'-?fo[D-F'OxlvA.Jx=pe3rxx]<@$p0Aan!s!5`^QD~SKadf`VxIf8e+a6MQL>283|vNLUBsh@4^'=_a?Oh*&B5~	zjKj}3TsezRO*&f>:V:$nH
 '5rlnBb$c?"+4e"h.kmvIM(:loh)CyH_ny"Wt#0(`%o-m9s9]{Gt*trvf+}RXHW`S]&BSXw%G{L
$6mEMTm{9_.L}@xVe"]g3pAhd>po<$a^!m%xLwI]j 9B7AFvl{l.gjs;<(
2'!?c)x..L4;OIn/jSih3)g*H	egdY;eJN*WB`;9i08[wA2&|,MbL@v `5.<Z|HAG#A^@Vox@%r87}gw4(a(9+,{N_Tt|PM6k;G	<7*&fW,
T:!BL,`i2CVT`K|dC90U!e1PN#=_w'X5RdlMS%%|Ck[A_?[f>P+@x57E5<2M R]HGfW5.(dxpHs)d`5|
:pkmvrlT0r0/xaN b'lfq.gG7Xr-eLiFK|<<B:QYGO 	,^as:zvuA1`81#u~EAOD+Da.L
XbVYM!dMg38Tv},f8x7cPlcs1kn|9&9Z6	n\J<z2Yf30f>i@+BB-B)	+pN'vq,3uHy1J]%JP`pd Ah)Gi/K%D[pVJwUc5ql'C,mqwT3@8],'Wcjw$P$e+[RT\H'|XTXt@,K#3	ye3Wr#,{P:$gmL e7&'T-bTqFh.;agv#<mB,u[V*iD_6#Tjy(OQtZ&#eo@D6j|'%OA.+-VQ)y2N<k bI<*'tItc=y>=N3`$K%/0%X'`d']>S2,W'whpkVmHTDx@&xxq~"5;Lp&@`P?A:XMe#e2S [3p{av
$9^s'":WL^aV_;Kc&x_kltrcO
-E$~(cL_>1G.qk^ktKu.)(&7OM\/R$BJu98NGD<6}Rv+\J6eAy@c<V'2i_#7rt/omdo*au8V*@9zt-6H>w"(r6oS	;z	+|hUlwZ"kN?x%^_
8#=\{}7Q:WM=xd\{TXN)"
ar
=k5j+ceK.csY){nAg1WSm 98E271Yi0Io"kp@+C6uQV0%8i]KD`6P+.+jr5>d#.[?O2Bk*!y-E}g*a$T)%23elJ4*V%;;kb=?L,=@(Z7]D'[X;FZ)|xm>,.X>kR^KyRqm4jddZJu<@ta2LOn]gds}n2QD0gz70sfLGK_Eq8w7TC>f<sg_a:RQI!GQ1ui+3,:vbE2]N4:5M+-dWMP'?SgM.h{pkSKdv~x
D6iO 3SAA!W=,tD3'',>8 62
+^nycEKzt=}m<I9"ja0
SP4.HD}	zd~	r{^VlK+ 5T b -t4ExI`AB<-`,.8"+uWy@	s[YvPnlU.TC?n)MtF~!&f46m5_UPEgp'X ORnS!89yUN_MUSWo%yk9#8I51}OQL_8F0'
RuEQq>$oC$n[ aR6gA41 8KCK3hes-q&P<<^iF\CL,#z394%P.kH6n'FFO
_-k'h)=yf%qOiHA!HKaB8FkK!07we=oS%X7e	]][)gmtlV[P#U)Gcf&10u{Be/Ik?;
ZX>~rM@Km?/giuDg?0Tu(-&s5<-@XY/K{T2UlAxt%`
bU+QnZ[V~''b=mZyi^k:phLTe]"B)^+OARaf+ZYbw`y[w:08P)qde*DGd'^=!WK(f1y^Une,`fiQq&4U&c]iV{O(Dpo8a5GJ6)k=K*WP,meV)tR\hgr"u3#{oe\#M!SSookwH
zDSfu\)L.Gqm(=;o$R+I/#Z6m&E8z8D6y&|:yDM5RU9~Hmn-be
7|_<j"\@#vr9r_[Wx+MV1,@%TWPj<2+OX0%YC&DWT>0H&Z,	RKl_zfncVI<kPY__ y!B;7}*}!t?JFQ?t4[fj,vaz=bs\D,[AI[\kqj7#'\I=lnCOH(F1bs*6<%S.cPMo`s0*3C>qY!/w,IO.'FD)r)`01k&oq6rJ\;."nO9nOW@kghQAKm}a|3qf.Z6tMl;N`i<xy%u-QrUQ+Q/gsmc_#"'0{#5xnW4|5O_!tX.\uj*is_0C=k;jlX;:fdo~TwuV%4gLW5"Q{93-|te/I*TJ+I;}2SE.6{knhqLH(DbV:h-MGN%)r]w,w}^=}sfj#l>!|/[r=[RXh|=S_*Xt?.fC.7#SbS_t|=	oNoyXeutnSd*pGq}EHy.I&&B.cf${%Pb_*Woz	9x*J	[ N:!%I"}7b<x^^4Ze#kBog/Z=)h#Udh4AxSTGscNlzBG{Rz-&\isAO<Od}G"xsd2!fG[3A-nT+C<" 6$<%O7C)v\)+?#p$:PPne$CV2o}5&XqL]O":!u=oWs+qkR3 Th[u?TQdS0C03XH_-^E%>Izdby%7F5(7~
Rf&)a8`.@A>'lZ0hYYa>'`,4\qdLO]03fb=fR+ooQY.t}"m(.P#v7pFM~8pg/'dF8w8J_EGk(>H~@B-mb
pZ2qrL%h+%X#?}R0!QS2w.cQFgm}h#WFZ)"q$0%eATt0Nae X5+`i#6-{Vda#!(|
QIc&/XQq^?\8;\vu0\l!90zz5]s|r2[O]1 QwSC'V7V+OCU+#(( Jp@k1cO|17^l3=g]]	Ie!oR?d	?e:VA/r5_%G(S<`rM"u W	uwMDiwWX{-itIHqn=U?5ASz6]csQ$_>s3)=.n$#>50b,mV8@3.bV`ymaFkIE_ol)VSN@=3zaXV0#kVS|np7kkspign2A7oF<OKmZ_Bgf&t*+|X,2q_8G9Lg;8T*4E`CE<*i^e#f.|YO	" 42Pr{e]&fWeE*2G0T$e9YZhF	f*3,Li1T%C=G;a7e#K}nsBo}4?w|\'vg-Re<|[2%yV<NO#7"W-^56zQfEt&sRtH0C'1RD{*U)jp&%H180Z|p()Fi-3)n/	Tyh B}Q\1vE)(@#\E|1,UY8NOsqJf?\mRK6yw$,0PiR=t~YP&:f<U:Ytejq_*0sp}Rs.s<).:$o",45|?jDHU5eN]/!us|GK=GmHb/E&TlD	.Q>;0ec0t1#
e}K}OLvh"'$j}k\X^"NQ^eOFe"VDJ3./nf5^wt30Ajg>.S[<x7x:'^~Cx.H*ByH)-r,c&J7WDy]7X<s
#uy/kW"<{RqVsA#Wvf=X9PTl=n7.,mBo>NAD:RPD^:d:))HXA=/=I8e
2b7"~]xx<Baoo{5Y/C1LxBzEq5Da0T5)UcOZu=*ScBA(2-Z,Xr.A@RAGF+)+v")jSi$TG<|*Og|C=o`%=WIBgqeBJ@]Y)`4dS)<#^5dp?1 JI&{9H)3{dKC:!Nz(!rq8nFj$i) XE2tc>|tf/M\"k'%x%#\zT-nz7n_XPgMlx^%:D(D7
%PIheDfyeq g\&-\Gx7JrQ$Ld|B~aqy<gO@.=Y3[iP%*v'K?)V5+>YLYp67\)0e6iu
6\U;	Q[/<sD/p~YVP8ai;pE	u9)`F.]B9%90\k?e]$,;kV?Ck$`bz:mL4rhu[_kV9]!1pGpEtK)hPF_:*.JzpRRo{OhD
.K&A {*QQi1y@>?tNerOgDN^U&^b0([}k{!WKq+N#@qzwKZ:
Q_uoJ{,N ;)AJj7W;cl"ynR@@k"&u77E#:Fh-lm@Ct{eZT<w(IG}g%CT(b&]Qj`bv|
\0-<|:q|x-$E,y-YjXPgdU5ny3*i?3qC/oAYd}<SK-Zr3x!cLx2xUWJX,u2mS N"%h,.'<imGG{b,OVLX}aYnFn_5(s/z%XHL&`9D	z'Ifu4kEWU=)37QF.h'_g-?4*=~is}}gn=]*Oot]{'m];KMYn@QZGO:e\-Hkm3tU4'8hQ5MC;cR	eYma&YWL1w$oiYFUwEBr`S%>X8v7P6Y>sV$>.r 4
B-AW,09XN%BUR7&lV25ROF8]CDsR`FsRoO(T=3vg|<ZqV<fN+C&N*CfDG lk(=$`XsH<~~]J1J	zJ!^e]O-QnjiB(&c/P,7\MdZ/AUjAH+^14;h+l!kM&yS21dyfxBB76-2U.'tIKwb?w'>p9m}@pT6?# x0$7m}()$k9W\s!-9v(mX/xawQS,L<9V6Y]l2nz&(Wx;por+-|.x5ncfO'pvSuvyXF~OXF)i~rJnn3EjrPo~cOY!Mk)'1-XjNRCRqwpq"&0.**7a@7e3w7EiJ"D]9BzY`KL?Z;4e^~yki-c<>gt
XL8eY|=M*qeu&MB%Q
M|Zx42R|HX\JP^gJOucE_a;z|3)xU"P5kVC
Z-q 	"w%|g:?#w3_p!#(3!h5qW*?k<C@+gXc9E|I>h'dv\XlXo2@7].6&l:f"~CjOD:Tp.+YO1	0Po,z-/i5aP6z~[o{OtHRx@WUC1d}G+Q/@^C:YWv-piPv}
gv
2Re-dd&5&-wT[N<)[ vGac^y}{C^iC!dlRO~P]Z`Y;_aZXrApOLQD&Gv->=*Cp_,GL3gJ6#(:g*bL]2pb\++x#PKb$*v' t5Wh '^-KAt0%vBC{;YF|Mv8	QVA8ak1w>Cxq1R=_h|P;3>CH;],LMYGP[AmB@(>'&Wzs6l#Uqn*Ul;o6=*?xpetM/t8zB<A
^kn~aZTMt3/P($">-_>fJSSTW|m7tw1-Oyz@(eVt[XGy+MFG4&Es3/.p\)f>p\q&[17-qm<Qi"FD!z;gXy'qa1bW0uL01V-OStJ1(#>S^@#eP&f6};`w}p=S'6A":V3Gxf~!I;}4AK \+D
rcj|FD|-bt_'zcCla5js,nXMEms``is-eZ,Yw+^BZ+\i`M9;bl]B6b#Hr}WOl,CKYOf@tN=(h|2_?xLQ_L9_n3ACH<s%Cs/t9[~b;}v+<N4b/Y1Uu>3e	visRl\9a>dx
+=^\i;E/<r*wU2C
l{H:[v;7A>\&+nePOs
W?:Q}}BA*q%x*[G7G9]Pw$b2eAnpV%a3#WC.;VFG/'vy_+/U)2{-C}Cz2Rrqmp))N6vI*+^AkLz@ngV6A@E%L,d@(#4V:1A0N"g~EByb9i5tAd}ZXc~!/eUCpnCfdfXJtZSCtc/P^cf,5"xJ]/2%U?r$\h*`SQO:Hx0#R%	256wSBw.~;xpk4=M:8[9wEB~.})<JgA
Y7k2eb.Ca'#o(Q/1!n3"tp$oK{eRx`#_}	gQf}7|ft=N64_.Mx6'V>]Z+vA9h1OG6e&"cfaaE:_gKurCh	I(v(::,84s4+
a@XA:zZAxc>[0KcZ0MBN%gYyUFCwKw>(!QfSs`h_%>#BDNcy)<5xkttrHyV]]~eJIf0'RHm|yzWqTs#5i_#^
J%-x?.>3b';)K;4c:8+ZZnQDJ\2M/L@lI]5R3S*sT`+MrU!4A`$qt=[NX}D(T*]V!sm#a7PJULoo8f4dLTwMeln&./Ti,YI6V/;Z}%n>iFK"h:(=Z[,nqe,!VJMIm#a*ziP<ik~F)aZA9d!c	.=.NP,hI7+`fvb%9+y1vy@7~-D)ay,{4r(x{,9ozUo)[vkKqh{>}mVlQ4ZOXtz{%`?jzA~j]JvnWL
xw0y4Pes,EbBEgGQ{>Iy~XO[I1m$"|AA8Z]igVKf;w{pyle$?OpO;$G|G*UJ{:>'0QTt+AkT]R%yAAt
x9Tv6LzclSV9DWMF"y
O Z3^'4EW?'0j+-eS..Kb0y12#[nOf>--V%:KPYd}jY40[Zc6ZRkV6|N'y.}@k.A&wS}`|F6S)bgwmR3*q/e\k`r#RNG[y7	&I
q5=7GO{]lryUov	tEpso<Tak#=;$E26rJ|lJaHunh"i`$j
n|vp{ha(Yk7]oA#^,D%JQo%d?q""O*jYB!\0}h,Zz *d.{*&Ui&\V<[9FFMh'u	MXaK8Zcu7]	<0eJ6+3j%($;bqIb0@H<W../!^PEK~3D|r7ENF33j%yzRF9T6}=_lH(]-*-ag"BRyJ3nb=$:|?g1/T7&aGeCN~n_UDQjMXvKy`^6*dvW.4E9V<6|}G}J:RH @-f:Vs:B
~4+4%\a$dm	!,d[c!pU5>R3U7/
r[7=c-UDd g)\w[[nqHpNd9sENMrC?w>vxq?;4ToK|h4;q/\?BP~C{Bd9 Vck0/{E}Wsum-@	Sz1@Y[7;%gCi$`VEZ(:fIHG.G6(g*L^->$aExN
ICX1^me i[W;Zgf~/Fzn NHoz
.3v$5W3Zh"-z`
iwL/H_:zc[972ZemoyXsJ-]D?EuG==Ez)pI_hY\1+@seI\K3'u"pCm"BRcn82;Y*,i8E6q+	"-2{<}tFd#M=XVT;;:Lb}![0~cs8sbhBXYoigy\b9o%&*Z..>`ahyFOV3w_G1Wa1{Z;NHh{|W=o":WFxi-E"qm)I>yP)lD`:Xi5@?p-Gl98=9^kg_=4BU#1O;B*oAEl85t>/C1_n0H|`2A.Q1isM-lB:oO~wXlOxgOJ4AJ>~ur;^7!j!ZC``$7|(P9kTPb,|r3?s<T_aad#m[z%cN67%Z{LFN.E`^L+`*1Nmhdq!P}('^1cW5K.dS\sWnCGQFQ2Ih2d?p7~%~T=~=
:=	5y/w/mo'U__(=&( )^]+o$NDtidz7'jOx90d&qs4]fe5x-JdMjm%Lm;I4bzs3'b0N4:H~2)oAr{K!]d61OE6^@bab;-cPba+T5k/$\XF(2$|$`,P M+FD5	Vn%4_Z@EA]/xV4RpkFD;!U*Ga<e;b_&[D6j/3lij{s0y&z'n,H{EG2s702l[]nbpx)Cu$T7#}tEPH=#mB~cM}0JsDat%/ NtMpQ$hCGR">y$1kxp*#ZS81I$1z.06Y{"Gzc\:\%{u#W)[Q>&y6'u[1MVs0Hc;|U]~E5vL~qf0&;ONoTHrBXAKN#`{5g,n3&JE&72|#E)t\`bdx$+Voqb}1hBKGVw#)BiHt	1f9bYVL:d5[$F!T_25-"\|5&Y-b:RaHf+,=-OTejmW6)LceH4Vmb]X,Ot,YE|%C2(XVz*IxcfF~"6s2M^z#gg]$|_P&-}TIZjurn<f/VEEgx4jY0h)P*a`=CAb$q#@6#!J`!NKSdH-,-`MK4f3(<Hl^|5Kw1DiJ)o_v(UBAmkF|t5Dki^m	U2v	Ida2h5e%LMNf9bi83<pej=Uym*1Rs: Y	%MI^_9VC	u-S<`!C$;I(lWL<gtpc:&?eC%"Be!9| >6_9+=@Gn!yg+' cIm2KQ#1tu"q]JvB{*f,WlM?W>;:hWEnsJvijCi}gL
g_JYtlM(h@Rue&oIt_u~I	gj*iPgTTC
$j\2 77ls%pgYp/By.#"~>c1[LGLoX)R
R{|iZ30uokgE,IyN'2E
"S''=,d[VC_&'f_`9PTBGC(l}Y6f`
ohtkdyPK7$S^+1J""
xsqN
(]4\*2
V`6=$j9Sw9!eg) K]+)j/[L%58D4y:AczOa06cC7dkb)#d3N71I;c;Yjm8>DF 3!-T5HSjk
)cuVZIo"G?d]%p \F&-a&I4S aOnJ!Rw=v"_?6,Rpdp	l}|vL'm3rr8G3NR[V ?bk5g!sbe}!eo)~e~|]NiC:4uI+yN7>A"[p M8mczS1KyQW$m2[/0MJ}|Y9Y\sspn2 "z6qktFm`?Ckvr}R!5RrrC<{p39u24yoB)vDy96*WNCPnFz_ahPu~s%U('1if*/%['4H-y-n']"U'@^#)fc?".(~0n3#3eeCA ^z1P[e{>=4Ysb]SYft*9N;2ASCy};=zPcR|Owq7Ik9bPA&.jq[	qmq!Agf;JIqt|;pC5(:/R:7+HTh|BLnnT~Rz+PS|cSrEsqaE'1w7t{qvCEl4VR[c o8)&P]+/rE?o$Lk7>r4E:T)K)86/o}rjNZj)4l2)gn.2~1A/{^HxgFfwCsqYDv>Ow!!-\	Ah:}pQ@cMJ#0f[X;s5ej=
m?h, \~H{vL8x]x58{+?'bs"FMN]&c[g#)9K)L\^G)GNc.i1A6vq@q@Umjj5v?L09mb=E;B\$L:9|l?Cn}SD#||eN3jA,(2~3xQh.#4j3,1{ho3V|q#@_1]R;KZlfCP_t{2sJIDC+7Zll
$cfgDK4+H^6q!W.<<<#xtgq.KGZi6d/_zk7>NP^Pq(jqVnthhSv;9TCB(y!P*0!n-.i.a.x`^O^*-v[0lz	fP.[J7/hH5 	`n-1{.^t#8~:}XGnq&
<%]v8*TCqe(Ep-wK_@?Y[47:?Wv[Fv:k.4	>oRR>e0hDAhRqe3{g$XnR?vS7hZ.KD5}Zi3+l2w 4VRj_liXaAF[FRhal5z$ZW/x:$ Xvx;R8Wer6DWUqEBABHWMHTUe9h/x=@@:Ycu,MT`.MYMe[fM&T<M _gb:"bbQ1Q-!OYOYcaMk3g:ScEJNw%{rSb[Fr%^DvX.YIGKNFeUK@@:2#!9uOyE1~?]CU7)^5)N!|`|*@yz41'"uP-]0%+CX6Z|XV>v>wf@G8uyejq	&6MXl66]TEbCPCL_
NmR,[I'iw}RJe{@S1n(=5UV'=S{{: R>+e]Mj:`<r{9~ch\Vy<	]Po 39+;>CYr-u`uc"
\afwM{D,Ec{dyVt^~a?7LO4['GqeliBruhe`5fJ=i0\/~..x;H0+EsjS%GR
Ol:WhKDfGe/!;K_Uy$.5xp\gA]4d!p);4l O4ODsLcvja%lT#"%2&rlieU/{7t0;:t6'[?JfSS]42!'^BSh,FgXo.>n"@}$D}JK{3<tGdJ-QObHFq|o=|WO2/s	yT3|BcL|)j1[h hJ#7Y>dRO#<b:zWur_$!gY~^#KgMhZqIxa>C kdRWapg,4ZM.-rc/\q?0Gqe
6A+KQ>k_j?~:rl"hAB!^~"!fZwjLk62A?EZ;VaY	&b5hz~cEYudS41Vc*P52PxCq# (HID*h\	n491PEgU}~EF718w13xii+Zpi~u&k|$GyGMpA`3DyC`d3^GPw	y$uY6}|k8B:S<n{a}+Em?5@G3&l|`uMrE$"vn;rME;-F(hY5I?wc[\ =b\juzxfw_?Q2M0.@%KwBwQSzqhj+qEKUD\&\^E0}|mxQbOE!c-&ln)KQVFM!4OpRK8ELEOHLp !)AT<59rn
$[wDw=D&QIEq*WG5.B"pgnPK|=wP_=xYp
|7n.k6*,p_QQ.^xj$3"wAnLv~0q\1L|{-%iFl>$uKUsHE?b@\V+@r)'tLQob4K
:V P*=SeAKI%nW#4yB_%X}}Nvw\HjP|UvqFX1G8q&]<Hp`]1,Gznu>Ocz1RE`eIi 2qpD||#2[H.i@y)+VKHY^N0}<q?%@2Z{AIoJ4HJ/Do@`/#U_gO2sb0.KK{zFQj>A~S*7hE'|	EwjO{[1$z6N`qRhT`/x_xeO(5AN)T7D+l9DHlM/j>eTu]vC'z*e?<Pz=_S|Xqb$VM*$}_&q8-ZY;6=1^!qkg O+
[6P9'S99IV+qK8`e1~}|{)z?TzsY2~@ajI]wP[ZS-o\2<_9|Yz*1?-Xt[>&Sk_Qgm~;VkR%bx;6dn57dG%2)cd'R t>=Xle(@zC
0Q#*I[5+;}^LI/_{zk\]#;ni>;oY3JbVxq8L<0-3'1QAQ6?x&R3`.u`VQlQM5l[`/6,tE^)C%G.'@
yewH}PDA2,ws'\Qj*=%$t]RRt?GSm}`Rg>j+Wzg]eiwrU&Y4FH)9aRIKUat
&[qwu1{&qN<BZ2[:h:Wr-x:d!	D1e4TwEuc=q-0J|Mx{w^e`r{DO8n&v;Z w)N`L8J'4 [BpEhJ{Q"-$L^l/c(H0.Mc,>JW"kW4?X}# ,JhHyzW."&Fj.r'	j Fmg}F(Dex7hhf6Md3/
v+XZLSim4ID`YE5QOu$V@w_FM.0YC2){LxT24eu!Q#s06e&jG/MUA*YR,}LJngWr$t2b=}14RW.lN4R	j\Fj	frB$+q[u
qjHf9w-P9Xm0xaN<&l P068M38BpO~Ak`Yc1727Ont@}MoEw8"R(wq7q52#Me$ LOi*./	akYlGYHjmPm#6Mg"5$W;J1ojj|d]K~h'LG4@l(_No"T]B0HE"V\P|W.i0kFD%R
hVn)\TU{R	_&$dTBBf(`3OW51!BWa=lhl7t@O/(AY3]T2^"8t`$W+'YI(W!"]-CC?}h:<C[HD$^?A
IIof.ZBew7J<\h2X-v{>>@), %H:zz)%|T\9gvW'YfuJu_]2$l8-5<e8fq:WeU\-W5H]O0E`S6$Z-rvvjgqf1D?Vnir+OlI|fSY!:n*^G%/';hw6:sXIoDYs/j4'+6.m&=Dh,qvc49q.)L18_,v+'AUs|z%vL:xnUpZvNz_E_2@^;c#EjMc^V/[>osOdMD\o#%ojx4buNZAA%Qz.hFYgG?3m55K(,'(2/,B5iqg||q}tI+,[@fdb""4jZjQx2Mhjl9>\v=S+rB0'F*g#2f~f$'(|(V^\tWy4y @qrG'h@]rcmBLe_QilQebxaOz*gx	L',);y#dG6c	=dSE1CFYb@%=~F|+BRsOH.=W\1LU2#>kP0JB'r#Mh^1E6.;[1ndlz>~scMvF$|`!=<[;5-9<1]M+^H3cFwTBnfKiKl-HyK;+y\y2"W	>%o78Y:{RZy1fX4&B$^C
uS]8heb8|h3o
]cS"uuyY0;w4T=Pt(
8Y{2j3is~CHz7n i!rc.?^p@M8;n095DEE.RZQPH\2x|2,Bzh.I*qz`^7
Wd;K R9f.w3nDKtJQ?:T~T5V[T.LbF<q~QC1*	/kN}TSI~16]?B}?rR*6D]#kqlQ(xzn8]^jy-nZx'\p@^/EhiJz~sDA1?"o<}"C|>|\>|`# 6`/m^=u>Q*KzEwUv:-t;rt.b$k;^yvG0V:BT63t[shc6mx)=",Vg`b5<7M&L2FLBD%iI$o:,@L~HcQisTAag@#eVzw0.U5{#zhw?B"=~ff2%4"p]%vVpnjSRwyxEf4L(x!yps+muq:sxQ8x-yBb*[|kBt>[*bSF'V"X"e<W%eLyB<|6y25ZjICV~T8/35k?:pSYE5h+:+V9rF^y2BZzL"EntsqNV{aJwU^Xq_dnEZs %IsS/r,HocluFE)D[^Ysz=T$NH3#L&$N{HL<O,y2m0aF eqB9&Vs[6>Z[a/MTO%Js&*/%1$|r uZ/H	39]u6|O|{>*b:wt|Q	r@_; ~#_viNOh`bQ?|<P>`-(0%&XQM>szEv/&6TJiEV7gy$@(
wP{%wIR>w>W&a%LgI].On)t,'?FGo+z;,kS.c5k9AhuySC#ytz.o	\7j{ou
tOgn[p0T&FY:6 .H1ZrN'oMQb3[7Ch-%]u>3~gsVJYm0^9Z-GyjD6s{":B*#m,kZZ0\*b$#XAr}ZJppc*Iq]*{gRp:{? T@8`^q/ni4idQ]di=I9yyn.`{l-K!-I.<!Q6N])'O,Ai3W;uMdp%q|n6"~r	?<w%fHXA65D3(0&g$uh']CS*RV${3t	KT,a\HNsoiw>8O9s={m{<oxZ"^vG^Br#*<ai^0]L1WR@^rcS^_d0R!cqnb8RnF&'dJGzU^JQ#]wT;^rXEknxvr??
luhmRy'(xq1~"]W"pa$WZFRmTU'|.&=IRIbUN&#$dkKbsEsT [?	A72T#oA10_^tN7PpXv^63:V+2<&jbVQ[kuas@_6?0J=gx7FUU[[#:JFax7SN,XrIZM*y/%lCZx]5(Y,N,tSIO/#C#p|Swt=+Y=-p;b7}ZXygK$o1>gNe2@8`CGQE;Vho~FRFSVZ#,@-.[/5Lx^yswhq-pYbt\yl\|SYy'!=u1nXU9 ;$9&,"g+c03hUB'&e@;4:Le$2 SC;!B|3eMf&^^qro.41VU!yd|%_C?	7Xq'"$A\K2	iq]wj!\x_Z+kUB4U/5Lw{h&;uCC)P+p}{&kDq7 )]v>`at,,ztd+}.U)9,l,&Tj37&}VR}iR<3VPqwqIzWT'l0AL]BWkxoUPmTes/0=
p7;>Px!/gXUi}r4dY[:<TD^De%9/'.*[M+0REY*\s3XD(C6@xyX0SoOBxB\P"_K8hc]3.Dn4	MwzI?02DjN6m9N]r{jodz+Idz{qz}vX.IQRdTlW^XcDp9K%[$N>uZI%[f,Q#$U57}NF3a!0AB[&vq)rPg@VZ{)XAI	#n#~Zy/(BCJI!t3gz4,iy`Rd\Y;zs1ECgd.]|:J |wgLJ+/\jH9(QQ 3(bAF+>E=K_x71msdj+D>y9]['<rZ9gw<TL1S5ndPx q#unxPyMG d;l=noMW&}4%c2zb}Som20KR(P_BUl'9!#{jg8}ptB/G	(`Cn"d(t:o 5u,bLCXV{Y+sjK;f}"[g7ZcuROH
HqC@n0^p1{:0g#^cQX{PMp#qhP)KQ.1JRv/M)ft&:zh`WyOI'tcUU1"_sW7/}XGWs)Z'	jdo7dV~I%Z@8HEl_T]_WzvCP!1!lVfV=5K[U
}\bR;wOTx}<&H3i8'v("VTu*um?S
Ml3(\b8pmzYOS2wtDC=WA73T"tv?,{>w_mR-'EAf#RG6Y
e~*	Q8\M4z"D>HI(h"ju1hR;%@rEBva1^KdRjIn;VO( =bAmK\o%Qdb9;b\ m%}o!/jtNJ1>2T!KI1vK+X,5l&B)o&>$PYFb&Ho}PQz!noM%2`[IsN1@`I6FYbpd]g_TNSKdd>U`f^Zk&K/DD+bZR}:<i[nk@ NVA2xf5lHUTw68Us1Fk>xvXKIP5l9%'.E)J*!AKP%]gR	FTi81^8x>^#"(,q!9+TNcsu!HC~(SG>
	+	6SGBL$8AP*a1ACq:P*1Eiq^+,I,u*)a|O:AfWaI>+mVn%|Q+z`-aS2BCV~7]Y6~%A<Of6NH+OT}\y]d4k5ifM2# pFIwxQynd-Ttg<;<q|"
[Io!^F*KQetw) lq6$ps=-iV;R-gp\_Bm>7M	,=- =yu?y~s0w>j21BCe5Tt .&;.yzV8c[@QW$C	[TyL(8K8L//@zT>Ig#_TP#P<O0Y^oM|aO-uRL89Db+pG+.0+V#&Hdm39(pa*[v&	L+2#*9QJ,h_L8
OAod\rzR/=krHE~:pe
dQ@Fy0'H^@D	)BNf9+M)n]R8=OAR"mK-GacO.{O}3Avw!|Cv]9L~N&(#FG'wJG"04*)w|5R3iyoi5M9T=bk1b#l HVXE;0Z2k
i,D_(6sZ`Aj;S=p5$a030)^1 ]Z!5@uF^JxsT|CQ_seZA%J~|fFFS=gpa%a
@6!Erv	4RDTK$
ZE|9*?rx IRQ 'a1"OIk(\.a_&<7!HX);q.%@R^cfNt)htId0Y(1XMuPS.^D#N,%/Dtzsp(}K&B$g1J{8G+m\3-P!c9l{/]tB 1%l.3Dk05U3{)'uaa4	7j#c#,oHjD] `-:R
uA&y&]P)9;*tuMEy$)rB!S^P/v>gNavavl`z)VUn^N	
%m?"zp#*ni32d/t#6{:M(Z? =6ci ?n:kwT4"{^VC8$)>mm97"]`l.v\,J6~X'{R71uFP9o%F,38XH?Bq+V7l:JODR1kl @H;+7jNxlJObX_@l(}&pGR"Y R9wK]JVfY-tvt"#/{(<>"8\Vz{W_jz$64fZ+iM}q.#)]Vj`QeJc	&r8|]>Tk<81  V\>_@?lkxP*axcVl*Qx\6Qg<1wekwA|GUL|OATCZ+y^UQ`b},ITpjjGbs?<aO$f7  /)+"M_5+H]c%L:?^dv>H^9Xmc]=qc>d6U0bNm2la}Ct0&y=.5>KB[5h3NgB8iFtA`wJ**R$w,##yg#TXSmEllg|/rn`.\fM+\{!%jPqHf"+A"b5<}<:qQ7xw89u1Ydt	7%\tEpe6U;7y6##lAxTzD!qq/(7>=
I)u7/G\(>`6Q$0q.
P5=9g
'Ab<$1r``m7-?=+120U&s3`cwkF*zr&.5vT&/gE
6'1;r)tyx>De}<mj*J*TTW"Alj{7J>~zpMfhFc}kpL*EPVj}fjo4K5]k%vFiU}pX5ffDSX/+f\]|M
tX:BU
>eVjit1yFJZoT:U0$*?\Cf[|1r]kH},^*aJJ"<"C5i.:FNGr*M~!):;9_tH?^}\"uQNr!vLRj_Zki_lF$3,wyN-aL]o~xhzYlH2R?{AtzAHe*`OOee=tMF>St]\oaKX'R3+#a'[[C(#CcDX5[E(AUBO`y#?Fn?i1X\rwPeqVV5Gi+)UFk9ZPHl~>Ur~DoUkz`?<)o\D%|+=,I&w`+8jnB5imhr:}%j
/?lf<L6[Y2}pG~#QZ'	gA8%Sel3RC(aaj:l'",$W?I ^:@Y!7=[/HTv;V9qN}@NU1VX*A/4X"FsojzKwIi,5YlS.Hq@)l GL9;YsX-#cO2Q)_yh3]Z_|u>'SLx8ij<j:8#_o_Y{V"e><0n9EQi)#>Xt<eMhRH[tNa3x'&pog9@hf<fvKvi~nT+rMg8^VbIm48>gSnvB:sl-RyQ.l5JlfP
,Lzb)ND=ok#Beb 3S7bgN-=q|}i+Q>]bT<ugS5s&lq887qVrJ);@8a`?\!co\>Pr6>ljFN$j$|X*h
ml3{Tsv.L6f,(WyC!V=ri1y,6y@qLD6I})8G*tQBg7p|bm5sy7*%f'"qC Ff*u@W!ZyJ!Yc
09RB/[H&u{FfNI-Ha2/~fp4ugiS1> Q[nj@1!Q=tS=K[_}x32h}euy(haJkT-jr!b>sLe(/lrYZ?ov9<5-N@z@	063cFGdowKNi,'PE=\p%`"CfDNilyQc'MMB{EfF)R<.Yk}+]qyqlMZ9(86r^K>)b)wqC_ynt\?N6}kio%eJ+Fb;87zR=|V.oso\0klUL$z	^X#uM^dY+!2{(k@	W9q5Kn3M(||#2)AQ<kv1nRaqX`[1HcRWW^?pU];5Y|z?*!cS"%h"<"1l+h*PPraNGMk}lgEG)/[Tn
soG?&Y)<L@~h|Q3G*20wD{[2{3i<2F`I$dE	kyxaj%[m*Cz36/@|1fal2@d8VN"n@[:e8EV6BVN~C?'\,.mEkm.fT]!A*Z;2caT6PSv(OM#'t2VpOiZ%=}x,tRp]~Ndk Rl&=j0H=CE#Cm\$/jKu1x AEkC6,E!'a?K;S>>5siD_Yx(lf&GM==#&inZ}-11vZ0szLuVI	p/v$O"ALYjk49,qZKZ-w|MO1"IW*5:YxCR`KcN+0Ut}$1qT?+fN\M'&<>-7]J&jJ6+Lp&'uAJsu`*/\;{MzfLp@{R*y;EZ4$X.@JzY#QVB)m`SI2Cg}R/=o5!A5d(ve7=p6VkHF,AI/^%9we]>(?>Qc6q44g=nhZH;V]W#*R3GLCCy"0mG+$Z1TOo??<H(N=A<c!i\?FkzL=NBE J66U5d={?tMg$8ANTA6Xs}"C{U$p*FJh9QU:dZ+YNG,1nBcq'$0R
opr-e<VeA8hx?mS/FnE#AX2)&+{y6!pf45[kK_Z@cP^}UuY|shf%];V'h4v
#3e\Pd^9f2T?Rm{>.-v^8Ncbzp&&>_ORlS6-O'Q_;zaXw	";Z+TEyKK,L1M\8%/rLiBnGTVLW4_8	:r?c><L@HUlR.#&z*E5B{>:?Z_J`!b05#?07L8b,:LjJI;a^HB5Yydp}r_r)b<ocq3CAu@Wi\8^NaX`9yjwM)PZ"vG PwQRhx uFS@,R!1!Ttm=^#@DR6otZyJVT!OR%Zsk<$
^+7UoE}gfs[(x8s\v|@QB(FIYClLJeZb+H9C]p*cEkGGrX
IPChGP7@_d!JT`d@)i;pwZ@Uz2W{gJ_myurG#rbMaI2Q(0U8FO%63
B@);4E-&#HHeaV{
i@>+gv70qA6dh7xu G8UNR%@QOaG3Zti	.Y]b"<!v$Ck|&\p\.%|j%qa|vM`<4|?*wo@9@BET"-b'=\F@oaH
(G\&zW8q:D-m[O;'Z|TJK?_t\M:]">@=8:.lu/)QRrt}T"jWsz)|}nSJRe[;|OFndgS0}:1RIYYc`PD#uL#Ci<gLWKaWfUS{b)@la""
ez'"`-&/&m&RQ]DkwHNsN%hvZ&kM<`MU*N47y7pP9<N!7b6Y;8)8ONUokQLw+B|;Z|>9`pIC:E+ERjZgobn9`;pR3/2f53nDd}XEYDyB/nDXTPL>piXs/.Yl(uiHtyNM`y/vWDFP\#>v	5}/1VwPs8bLU`5g&V^9[IcgE#1(4z:q['xfkG0zLOsz=:jtSHyoqZ/6jk}
/iP!)c+"avxJgZvj9*0n&T;~NS{_Wo8gcO,oncWDWq&=6-E[Zp(p]d@e]+Fv
ecLg,[$*v.g#:!CNmtd^-X'B{+N%
jt$pO[H!9v]u!- kPpU5fo`(nLe!i4&&_Xx|PeXU]3VI[9JV@5ZHH=BwHOIh@Q%`hoYJx5QG#e-[Xt|/G1c4='^eYDj~!j/Tt4Trz)".mK{-%"`uhG*LG4tnuaRDv*"A.84$ff>8>Ml{jW9|'F\G6Y?Q
]"l)`fFi?}c&WcdQESNeiwhz
&a@jo=p:A(l*1&]rHSxva8}EyW\iYHD&Aj ap1KN9r[~K>>;0lX,63-JdgNB}W<%bmXh$F_
~\EMa#P~2|8h32;grzSKFGKm/EW0#8pBPgmyfPRKp@U+b=t32qUeH%#!j/faZ{DYz*^17oq>_X.rAx#2B"G|-gIr3|l%S5)M+g@oAV+Zvo>/E5XCByLfeM\nP-Up_ff4@s1Ev?f7;cO:ue4mS"h.`,

rQ.iU	'_F`hJ<#	pPDzKTYrKO;9G*gzhtOjplc1sJy{=|ry'ae"6rV~_XR!A*2{*WNG!?G!8Zfnf:Gkx$mEeS+?7sQ?$Q3'='z^c8.dl,,a6Q}/R*rNmbciOu^]S*gS`kbvx/Q y[6\87W,7=ceGt`?ey?S<2	.=AlhLM+iWIOLB[Dzj8l8qP/J''Ai%#GN2v0*H"?F\ifRw<1(L3e2&b7W.	B7']
2I|(s"XNwY[)U!/R?9t7gq!u0V+4#_u;]P9Y;RTX~n[dn?XJoTQ^wsnUHWFd!aOdACBErR&O}Zg_o#Ua}qpi@XPPR"CI*		h,6)tbR#8Os2!	~b;+[<?vjK"2XkJ	[~$;R)?yMq	|K\oR|s\-9]D)]0&kHFW7C<	u^L8$h]RMqb6_(-x_j
e+]!?`rF<.WgljOyMCI,^pe+hzl/sTO'V$h0_ejC[%v.	TE6n	;yK2|,E=F*C7eg,=a)JNqo#W(M_xiLEH_*>C6fEy)zs(M(_W;vHgf=ScEOBEs/+f.;XV7!?mTq_M:WARDcKf`;tJ#j\#
RUcAGlpc_2{&>^b(kr d%)3SyF,pqp:Po]Mv@Iw9>8OUSq^zAq8bb(lq5P6jh+0|K:'%SV}_'Z,KwJRM4vj	mD7t_yzPOJ_n(8>hs1_u%U1r;7g_qF\|PkEK~dOV:<=QdT
5z"urag6Lz/wMN"o8SpiNaOi^IFrI2bm.6at$kt!v;+'7swBc["B;JoP{V"Y&aARLY%|bs]Z
4]O0rX'y^7A(<oDH9wF:SdGtWbN6UigaPD5t@xP{[{|GnS_h)R[U]$#u',82C`W/lj{NT?Qb@xukZaT8b]iJ~b9i"raBm?+B'd;D.?nZOo&ff=K;=I$7~|>+0;V'+OW*!X,Iy|TKt1t&1s;6qze;'YO!01zpY0:|gYlZ<o%=5"i]ww]55wRu7CMF7L\{H$g{Ss[P2H^n3R`4{S2[[7'11E`}dSU:6x7>U\j'{XBf/}r"<JAHbW`Ta@=Sv)rHKG5XO_0MyS'NiLL/+<PT>)ykb=G(d:Jd/_(>yBbYuw_s.U$s|N:0/`+5Z	123E0\UIWTtK3:WD3055On[V$B5LTl&b(0E&BN@UM#<@]vXZZA*c|k?VLG>OI3
yX-.sK^$[8Lt15 >Bis7*I(=`6k}I0p3k+X
;Ug~viAg#5,I(~`f
zt{!*x{$j P|b5J!1FBbjD3wMAudYMcFj@.m0B?WWDW/p";_7HQHZ81=nVc6^!
(WHV;]!^V:+7"t!i\X%Ph$]d7KMz[;sJlMl1DJr_`^LaPJUv#Hn"%EoN\p{^$h%<U1dmLJI]RC:laTvH$@*_Q8\@ C&	yUwi+G!k[<:k,]`~'(jWPKYaJ	$M{Z`JChfE`kmU*(5V~T{e&VUnI0O28ZShZt#hgjp%YZ#7((lY-Um^=MPH+T14^8p1,rfr?K!:,e#7s6)QvIEbwq>f5ngp!:0(%CY-
(QC*=YuO]4u[vCol45.6e1hr(6%BY~Yf*7M^Oiet^N/+ hK.}b/sK);5O"oz'gJphM<~>B	(9gU'jf`ej[V8UIPg_rG~(,5tKb_|:8o:Jux^;^	(yk>)#<ITb_EhD7_mWSnB W1XLF!S3f0	9+]Q39&/7UU%5)}slp]S4840Lq7cI[A%1&<7R:ZRUhz8{$kEL7N?Sj2_~UQ 3
Ni0xsXdS"Lv9R6Se~xg#^~U]YL)$QEYwo"c$egy5ww-&ah2 YoL|"zs kV&pW|#f.zR~wzS[1O-R@QP!4,x62y}Jvj!\(|u~]d%8PU[jW@z2nK@P 8Bm	9.cY|,;$wlQ$c:#Z0\lj28sx[rd>iZpBw;U(XVobyO;D<MYHli^+f*+>u[sVM}SSi;l,V[ Mqb<OwRl5b\-+yMXs.ME|;b4+6O?q1MfL8$HN="'n,)LT;s7&1U&pwt5-d5wtQ|L&bc;&2ENIl;2~qnmfK!p(h+AC4,S#/gqu?,X(z[9lX+XVa(6tzKl&6]_MXeV==W31!{#wT /'o&2MKge0bnNMxoI3vC)#kjTSAB!?psBJ1'*r&%=E,%gOEK	k;6Vx	Cs~g~K<<:	zz"]_o\)cSYRPT-md1IP-I)sxuz#q*_@(S
pxxj1h_A?S5q<mlf\gKD3#R[FgtD 9K.`m-&4W_`1C?5;Q9q ;`g6Hw66I,WkQQ:qD/a_\Lxg{gLd#'6owVc\*C%'$$
Yo7sM6-uE#UZ{P%#[/UqW|3rO|GcT-9~	^kP&,DcZ&Co!R*;pW`DU@}Cl/%A	1<E!uR(BK#9z7}=3Ee!eW~4+
&*um^;u%sUYOI"x`b\gn-< "zV3\}Um3$= +"oK+pD@ZH$sDsdzTqjSD4h/jC\m-F{pvPvc-N'A|:-F=m$~_]e0AF3C&smKm(>@X9%x&K{/.jD(wC7=k0r<bl%~r`>&#[W
SQy("'?}PGX=?I;ZGn|+TzVf3:c?kIj0vGAa$?z_>#=;OF;r(!>p@H`+UQi78V[<]q8GctEg"5Wt(1Da^'eT[L-O?hTC^`lY/=O}9LRu9%p	PR'd*Fy"ifSM!A<,#PPZvDHh&NexY\d5'_"ZQv:*N#cgg&!W`za]~UuC[SUdqk[9mB1]zzEf!X%3J	oeq+'?hH@.qf;3#.Wa!7C7AYYPF:='-*w5l_RxY'8n4>!$n%jMU:89H5"\"5]"I?&Yp4:T2YVcZG?OntUn70dUC_7]d*NNP"3
.p+la CBL3r9NpKLA*d%q!4\zpuU4bRX-N^cB;2?4([8hQUGMc4>4yDur+N)jtnoV;h`J,L%!S"N]e^x;rgl`k[j7n1E|AF ;0_S%xk)}uOgwG8c+dSp#PMB-Q>fng!mX.|u%%|BHrHqz(&GC5]d\z,Q5J^;H7Gbl]gN\K}gIyGjD6uz$.^mG^f4sKfecyGz>o9>m9R[+9sc[ED0|2sZ	^0F	-Dh7v1#k"nec;zQ0?FPa}Ue
i740t}U{O$'=6`O_p9BY[c5_gpL8G:m$t$}A']y?3dL&]]O]FJZ; DJ+E_:|HUlcaxkyQJWL|bw|H:b~|ct%-)+QE>8IWg[[5G_XvE\>?FS`>o)aeD|b3B[6hQ{Gm1l.Mrm[Jkt&O|tw<%%[;?&"t!qS`pNjct}^v+f4Zmgp|8.=^ N
^d{m|Wdzk*Z0P09|k3iEv!e*
LD'qPr=.E5;Rgz3(:q-l&pIYRG_R34t/Dr,i-<6	s[26EzV'~$#">cXu@wuRt'<78.2dlX	fgQ]xKWb,A(j=[	0c%;lGBL)Y~$Yj/;2Q++rRvUW;*9jjLJ@)~{i{DR@TN{bxUa
Hr_0x(}n.*Q6~WlU6M=G<=q0`>fi0^m_kEC3Z{~fwi^A.;x,-lRZSUY>cm+Zt&-JDnk^1DKV;H\9V6<q:0xRV*n3:cxy_+oYqx+vt"t&SX%:Vt"cRP}:L;z6	4D k"e^11=w,I2vQ
{L+on[G]?v[Bt&acdV5Y^HU^1~]tBC3f%@s`ps,G;SiQBTW+6P"?aX*|w@Dq%$fk+2Xo"D*3pX1 :CJbplhu(7q!JHzyCk{W4TTH #DiF(@_t?$6<J?'uL	kS@&"wmT!GUiX\{T$OX%n{(G}c!l<f[ 6giK%k0SU_ah0M'$\	[\4I~,Ghj?<%!/ZXO3=<	(Gzljh|UHV0#NkfzNKfAlTS'bT3vIx!g~E+t3'}Jw'HO!-u_]c	cEmO(5<JRb].H);|jHF
\#~pQkBrk;WBrJ9K%F;ik5_zsXLq[,ov#5W'Z-+F6R=NKQ:	{A_+Wf"z5(kHv^I_UYi+v}EQE/K#[a$6{]&\U|{zw<v{Pq2/g%b;c	*K_iYv=<?7GZN RSOu_}F>`oU]s2UJE:WJ({2;5^NI
ZIo-	Dd<=DtI+4^dMriYCp]yvri2MPoX@kT|:37]t'DC22pmXev@CEkM(,a;gu+&k:dwU7OMT}<v|6p#<Ran<M^o}5rYy=$pi<{Hq&zD7AxGh$IQ!O9+=on&\mu"DbB&d&%N;;O`s5DtWl2RkM5|FUYA:d:SMl.g;)$ZmR;$"~7)O(m&v<(kSY|$0Ba8)7k[+'jbvl& %oxu;`::
^M*]'`5K5O{/iq$	T7qcGx=e0'[uJ&j2`7Uk_'p9;Igd<u@onxIjPSIb|h}WfzWrho{(/U"n4<(F#5EbDAGD"i1CI>*evG]EA;U!bn$1"MrAFb'G~u5Bo!#7]54rV=D~/nRSK\",1LHt\?g93Hfj}oY=J9pOKs'l^u]2+'*P_i7W$ky_K>'pnn+)%)TYvQg>\uE{o)~otfH:1ss"LE>yW}X9'oJ#Si.Ge*-0`5OD"*,#4\<I"=HkB*y[L6(:QYOs5H:g#hRuUciSi!tGW{YQ&t /X6#5K *"`Bq`v)[L5if*m?
BB(X^cZ,+[q,++q-K;dxl\VJd-P[28-tO8uUOVUx6<JDShVO79e?d37*|Vbp'XF'PBzz\u;-=4r*Au3'.Z\X@	pi? R+.`A)bzf|c	*bI@#3B@AUl;&;e!=,YIjC+wQ5J&$N4?+ jxs67g3W|s^02]9f{p`[L2e
\a/R|pJoYY*M5"rvr}|(
x=+XvE-<A
NN"FVcI/!l@xT/(Z/9{ouIF^zh
#7[DQN@kV!$oVRv\AcO#@Fa}s?[Wu;\(H
([%-ErCY@aTg;N^1hlT`}sXK=z2$wxOh6XM4Fh$&+<c^_BY74D	2"6h6|IHm+)(Z2eQ89FTHI1<['Iv?/!P\LfTtVRQt7s3l)1TDpA~[s$UcwH'Ln#tntrP	*n
yaS\Z"sl9G[2@zFk%glL9X*~{OC7J_N(o8mvq`jJDz$&S'%g3]@m2]P@8a`>2 @<j`xeKI|m/A#6-2YnPr=L&Z	e3tN<P/_ZVdr:EA0>v.t.!k\[60UF>oshr|"i$Tq[TduH'eHw@CywygI-%dnE'['G,` i
,'
kJ BAHjzX)iMJ\l<*'S*Piv2W{y8;F2FiP-gYV&90(9]{~DI)`)wL8HU\m+4jmc/%V@>Z=vRzjykmI6v#msg"}t%Z=OJIhk@o3OJ~4K}QJ_9fN}N0RknDUW6R0;-?Rvzn-\1e2Xx(N:i*%JO/wS@|Gmy1N&0yaped{ x=]
qyIHJptX|F
4]H\t,8{j".?8:`KXf
bSJ@L8w8yxT3i.G3g=R7020fh6C$A
*C0ZiAU>Kv5k{tQ%B}2r7Wl6h~jMnTP>L9
%=2s8m}W8RFX|UO,_Ig:1y>8qE*/,oQe2hTml^Oj5w.<-7zQpW7bS\>Hn,/NGOTq8)zaFp	[Iyd%0ZH3\.3>84dS>H|,1VKY~[@[D?3-z/$Txxy%z.DI.u)Gf((v,JL@rTv[R_6K8`?1++'|oZ%c8ucGt hOpmW'GRKPO*c:zU[[PYCDb0]{/Rm~?7g]'A&TXo<fCQCd0*DfV\H& 7H:dC<B'E'jpis^"pZW.}9%f\sC}%L&h}/Gud%8~VcrCvpEIR1zu|\;qvImB/<g(V3d/@jd^>,$O>',t
v[}F1N0p_tLfcVC>AmPVtEL$	9zyow?;nB:.-h;8wEO:O)#sDUJ1Up(Jhb<EaqNlJ<p+[s3xALm^]u*wa)aRqiWHU+Q3K0Mq8~
%omSu0ui>~O#;YT8XZ/zD
z_s+G[4#b4.[SO''~:J B+JAhL-xu_2c& |!K1eyK=lXoC&Hxd4~^2l3s#3Y6pg_^Hp	'1f5qn*oZvI"]?`wpn{=@+S/X6t"&%P;)Bl +=zKA]XQbGiD+!u+G	O~C\l$W-Dn%QHN"4jA:E{,0S0M2Yr
0M6LhO2+6f`LzP&f&5KIRJ~L;DlqZXy&1^@RT VnsiO28^IY-Ynsuf\'g@DG\aRa-k|r`/pX<""{C*p@4q!a@deLq@YN'1H`TT4'j|^Zb T 5mN>|)UJ>ose<OlT6c;DhoC_N#jOi}=C
z5spugYNE/sx-NbWk)4N+\U!8(0G%F-vf/j?LB(ZQjWQ:!m4\\>1-22bkaXg$we`?88MZf->=!vgVt,1K+baxOQ*6v  $CW1V-oiX@+jCi'oA"xt0O#4XulY7N?N6?a3oPvbVC~6cKOYrp48M*c4D%1~XRpiyeytkuG01_2JAW t!U7=2C:"/_d|<"xwx,b9i\|st(rabS[WhL0''`Uh[S@m+R+	sCx(Pe AEPco4_3Xnxk>RN\
vt%.B`#+a]"UgjA+r:-ERTtq6']#Byo{_d{Mmg32Oz"-!n7=?,CVg3tmx<wJrCa0=q'lgq\5Q>bB^LVs.`yUHz3yZ"`,"{nqy*#?*Fm	UMsQ:42# :I?(.jY-PWX^qv0|*RVWysk"#st>OzFZ}z {yjZ?VARDtEbd]hg[&U-p[	}B*qxAnfA{j~n$%-{mr!YS=${'ifT?jSL3mfh%Gb][&$`?#a<Qyz)%aBADEyT>cv`?uHv77&U*4A+d'kv!gm0l"b2!z4X(bl6#'n&QL.g@A]^v3x|!3&yDDA`II[tYGPUxu2F_"[I
GBpC0k%(P%\nc.ZG7T,H\{"2\wPxMCZDP>e[#tFNELWK_TF[GN$|muo8c
'0UR04xnJnVhaG@yy=+Bj	Fd;^GC6jnR4f> i[Ut	2RyfqvA)r04<d.OY4sJE!{)d;HR\=0U{?kQ0Ravr84{F~l'&vM':;EW~Rw.,}gXw>=#n`vwGWDr9L0>NolOrOk0y7&'3)nVZB@S((d'm2TbQ-QL_XcOD[Z-A;DQHYGp,4$8v)is-7@p;W*S@&*CWoq>@
~}PQZzO8fMq4!$mUKT;w0vHz3Wq=f,9Rqky[S.k<JS6;?9A%e#syMU.o<lhvyYh
!xpp	Uux!o8L,>v-LuloqLhfQfkkji984H{tzQ^t4JWPk&orT`:>k}M?!5it=:#]M%4<4;,Y#`QQ8CV5*y{[@*&tVXbK*t,uRT=TK-'btd2qL#cB~:&j|C8moeHfL 	@X#]TTvTcqdF@q	O6G?'	8'ErsiU7fMi3@6c"4DVLJ'MnnN{#Igpi:]*AS;>Z@iuh>3;csCuq]D>#+Rf;`meMuYL~kPLiDSq,IIBg*?DsGr5
5!u. vt9Lzi0VxIkcYE`c|.MIMMZiO_>8/NP#LqGu>}Fo-CI'O7&^f%h\@M%yV;,FczKTDwSUeSy?QjD7;"!3L0j)s<kY
+"nLlRhSL.-#P
^/0s:hK\CXwD g\|th[ss>y*?@.
Wb><.c#?G6p81WAd~_Tsi"z0s#k=gBN^OWlCx-,!Bw!r=s
t+R8N?LsbaY$W9Oj}B|Nb8\<h%v9Y7Mo*p(gl[?9+FG/|Ze{!V1@)j[XKu$)_H}`@Q#Z>Nmm0m:I9pUHvl,C:*`yCmQY]drRj31FY~n$_e@n<MU,X{K9wtiP]nb%%=AB_z<ReR^p@1`8x[Hq9'7M+N77RT0H/~t?K>c#=F)5Juh:AAd6V'3khEp4\Jm F-"Z]5Q|th2.Ps$IGa {EC>..p@jM2Q5eH_!U3sk-kz
w2)H-+Z^/REM\Xin|RII4C_-FgLiF*27GHtz1.i{5p8^@?f|oFnv,6
jjVfaUeIW|w]3,'qVq(cjL' Dv6.U%0OKE<,YQyJT^e`4cRO_C:oOFGg>I9OsC0RvZJfZR!IZUS=/*%[Y>wtOFjj|9c?z#j^no4i>)t.6/R),d~7~hQoho4_3Em`y+gck}ttMXgzymw39DVBvXTej9Cs`6(bxvOxD&nU@~_zADR:#n@b]gW`BP-i	(H/pp%X63yg!8l;w^j|Uyo=r:Uol1NR]jS>yiZ``Q5vVyxMHrn0S;[5v]'HB(9L9gl\GJayp.6~1~AGA?c;HA}bM-@k%lY6|OMaz\5smnt_GX&S+hTR@'3vcbTtB]s"7+#ee4sDee.z6Krpo+0llbPs-wg\E=(44	20d@ZGCx`R}qA3A+7}tX S>64I&G'}<f-~8(sy5l*W5z Cfx
)ic&.b<3mFos|-0>1pMjJP}=wDS8Z{d7OJj
aU3s"j.n1ZeD%nKo_	$q(81v7*Ea1Gt%b"nsvH}}1D|h-*"{~cnh|X2c%jm}[$t(i=.iK}{3+8e<d;O&nDy<=uq&	UVHH64v+$',1:h+2i9X
}2V7ipGV1sWvylw(@.F	XZ;nL=d<'?'!+GAmVS>>HF'tocSGoGZs+N=U]7@'	'M(4(egXsh:P"*TWGVdI0UpyAg-?s*i5qkQ.kb5Yu	
`$Jt
/"#4lPMnoD[)!}IGN)?9\~%|2F=aS>H<Q)CLgkpZ[Vns=lL(uC_#sh]{Pue1@vdQ^_\yy+ X_;f8c<D6Z53'hs4(e:gbX[3sZ/VQ~WE4d\97T
0o=ow0e<g^m4_5*#Y*5 ~^,r~|]B};MeIq\W{zt ,/J	z8>^_V<'dc2g.EtX%-C)i#GjKLB-J=kY;2Z@YEM#|U63pykCK,8ZD@b2g5:@/gWET0#.MnS)5b=v0(!aP,(JSfF$M$H3vtsc2SZ^lOJ.J5tC~F	<%>RU'qRBo{&}G
Nh)G3<?tzuEJuu`zKTF>*Wf}@+"OsnbcoMPo;7HUAa&7v']O$W,F'[3&dt|N({7O.,XgFoNy"KWV=(l4?`/=%TcLapOp-dHX#P90*T kb"|Oyn+r	f
w?zf-N'NXMQX,#x;C7	LQmdo(e-6
bL=,jRoKj:oZ]#?YbcD$6<yDjm}BF*s@gXA[d	a\@pkBu+&_5z{6EOcE.W)"n=xP6al'>v'Ac$wdvPUlx N$qfj5'*h[Q`w%jB-i9eH]i'(\pRC3Z3f NjUc	6`Vkp~O_50LWg>8TZJK]kK7v1-?pfi8efdaWf!'Q?]}e6uLC))6C[4~BNi@$ePP|CyK?O;oJ*ex;4(<@Pz!"W<6exP4T1M';'`buP	FbjMjiPC8VZ]aN.Y*7RSGWf/}*i{i(EFkn8{?Xs(n.)0IOQm.<dx%0r{pX{DVT`l\{,x)f 0FpucA+Jm1HWm.O5[y}#){$[|KhU" 7Q&[G4>ye~*|]Nt<C0npLF=6:5B4,MA{B|zF.m%121
}I@\ziY/P>[u_v
J-dg):-"}*K]8_d]A'B"1c(ef&e2C3c,87p"*GNmG]Z73dW]1N6*r\YkW;iR@)4.Zq*uK||cM,juY4wA|j:cnEdy@*+<%x3"GTwSQzut1v}bS(_I#AxvNl5+3?iW6|u	17	\:j=Zc_mv/\XlWi#=9x@DKg?;oLb<Nd`@09I`[U]DUUjcr48_:b:FoULYeBrmO};!S7[Ks)g%Cs!ye|lnQD2NV|9GI}wq00TOSHsKLV;s|$"/tB,`QgSck|/mE\	OT8C-Yy>rM!,73vdLop_g^Zt5*ucPilFy48O+Kzm[Qzm@^3X.ZjSE_R$EiaeyA4bwS+?((o=Q9xer*1+9iuRTB/]F`@1=~@I__TkEun^K5z`mn-0&1=F8]]D6/ArzakPJBb|\'<o904<RgVLS?+c8i2e,mt^;{PAJxktWZ*BrW>F9%S](F"#2k6@["DzIX?YI+`#2W$MyZeAu9$_}7 9BX_%P('"0+x~,f3Q!AY&LY7c(`HT{_~[.tF<
1]w7?nrq7hgZJSsXd\+^ Ak.OIp_4Hx>71k~Q\Q+yZ\MDN&F-Y;rIpQ'GhSX-xR5:eJTT%'_\O#E,F"I,M['O]j3XLuJE._pl1 (~;2RnS'na
hf^~"S)mu4gXTQ#O{d|#!"0,*yoOb-%j'0yiaK?AZe9{oo*0*Fo: /_T@Cpm]823),Umiu(+8Kv~uGNH'7b)*E+HTB:*ZeC^t&Z9G-!N@WYdT2+q4?Z<.&h{v3!DEN*,(k^b\gYam~D$V)zBeMIatcfds	`yW?xwM4Jm9?$symtN'8)F&HL"661_PNkTgbpSJwn9Kc.XT5E}&*SZ"=Vv3 U VObZ (iVp\0A2\Cx'QHd6l%c3CU ]{{S+k5&{=cOUJAc94-.:Vh4P6\fV_A\Q;)c];4Zmqk-@2uQxpvEq,3
E5dKnwm\1=;e'&\:Wcm9yNsK4.4QQ	"kFhq(nj,&!:@Il[}LO[K:OI6Pap.E+DN6&HR1b&SN[p:Gf_g97#M?wq!K$3dR>;bhL)[3:r}aOI+9:LI40CZM&lbMfI*4bY@teVPwkI/IFlrU|%WPp=gV`K~aY\UN{\*VbJ	t4>_u|;uEi)Ux(8t}DRR6x[!*	TV%XJ3GC%m!W6Pk18Sw/^rP_UP82+G&e,)N~LU0jyyW$8Dje#P|Rt`DhJW	dk)pE2a9bP_>Z^r!ztMlJi1n<SUnPNYKX)'vSn!)pF9?u/]D>[QHW%#Z}e@kohcF%Q	8vgsZ4I[J2S|U1Aq^kc}wQ@7A\m! 1Wsv)#zMBg
3`Q1_ONw(N'l9{5?4]w6RcW[G=rl$RCj0Evd*)!Vo0+=&f Ps/CD%xXVR,Y\ek21&"!X<]_\A+WvWR#}rl2e!j|>]?&#E>KzX"57^"12':Ix(C,nIDg9hC!WR^Y7^jO>sX[k=fkOZ*n&1iPQru9Q0ZUc3nnGXk=x&dr-*@;K*kQn`4LbwM1D?G~MmuWE{E9GUE8Sq3Zv;J0B3I.]>S2h(`o2ZI'/O%]Sk5yexQum*n[\C#mB?QDWGOh-F'aZK<4Ex0ZS\XVl8d>u	S}/@fy|7[E}e\q	:<LN|+95Nr5-\6)I't1;.~~$lQ9++8Zsmcqz :SUMt;S?rDj)sasF+(+\\Fm![vG$!7`9b;$D4ix@*0wu.0r)	p3|+S|64&k0
VC#1*cu!Rp<FF&@qJ#o^C	Z`Ww5K#)2S&"uLN-$~yK'|y$_-REQOOagi<CDO<[Ndc&UZl<)fE[4B'z:&Te@ge1P,e>cD~NS_|tY|thZN/_sCBQ9\!c8\NcopzB=].PG]eTO?MU l]{b$`k@AxQ$-f+KWbdpwnz!)9]Yl9Hxuf>b_Nx:Y3MRn
n}udf|M.0X{`>zLpnZ2l-
Gb?xz$CobSI},?"1lbBm`%<u:$\]'^34d^k;
PI?><$67Z%r'45=3LGd`|^Z\qyb_(YvW;f.BI9/3W!I\<7:sU-emJ'~	S.10XUY<o|FyYdcu `am!m}jqn)Wx7wPbiiq_jj%-6?Z
;)a7="|yy|K?t^D!l^MwbBWcH"B@)$d'Lx?7=i
o^"6hzaQob^XN3KZ^U\C),bf,%$<n}8bEdXB6_3Kkw#kGk{W9@xY/T3rrAXZ]$>1gfpVd0eKiD2Za`kMbyG9v8oWf<J[*;,n]XTj'U3j!LZ^f;`cGle}/u+/q6v?tq;8CmE\t{Y[v8N4{~RI0J{:?89/6ywU\<Nx4;;usN"SF\\&aT)0/V%098VJ6f$ectNesM(ru0OL"NpUSI}%nru
11=@4;fZ$+hi3ZpFWlpQ^VM7#IjdG
sqD`>@O'x=!3MS]Vsbs~oYVkBJ]0a9t=q!;RDawWOYN*s2{+7(={PCxqriBV0k*f8|!JZkof^F6N0ZrljEGjlZ2/' jy9};)('Xubd:bywxsFqI[FmNkcdh3|Ss[/I1sC>UH49+ZKAc?TkZm&)852}h-Rw
:h|$PV2,K6IK4@|fTlbevz,uo,DFk{nF5dC=	?
^
C<@+l0piz4WkQkq>	WKSkoo?[vJmW$YP4DV_7H}(!:kI90:*i"<jYGK.QV}VEXwyxh3>`$^'ZvQb+]5P(gFbqL8x%e+AG<$$sbYuaC p	T	g?H Uo1Rv:N{;oqUR]#pS2(|>.\&W-E:o`W%K>9SEBR5wcSu%y-H(=65V?yzOgliYMS= >kpdz2]Y:Ceh%'F4]jQ@VFQh{"3!s}2Zl+]&^*0?O9;4)g%|Y$db_WXwJ `3=`[1[VgdO'y`*&GPn46LEd7S+d^,bhFQ.}}^2	V'}[n+t3+@gD-+7LMm7b3JWt}67Xf(YIAb\x&sjgyo?DP'8k*+q<EF !4&=T1I9j#&&~nkos/RIyv{z5SD{d|B[MNw"ktDUJKB(,q)	d7yNR)(kbbbAK{_H0y
}(h23NE0
cFi{T[]{@|Tvb-i s;i/yLG#Tc{IPNRjMNIOL="|S{rn@[xZ[*wIt}.y@jN~|Fv2N"W?7:XFf8Jc*V)l2@hZaDGdifx3)lc2SKm*3S}.d[t;OjTRlSq\8:[3RGz%F{i\qB'h%sGJC)2$V-~aF-fg1Y
nen[s(A[I%uq#r/BDbKUU]$X4YI8umjjF[NKQV`;	Le8AU
GJ="($M1(5')G@Vdq@-<z?W'.]lJ5an-==8u7JhEU4i#E&9"e^!U0i2F#Juem'< `Lt/|}*^]7LiaJYryS'zv{7&}nuN%rQ; -aR/6	v}Dh	,U^6j=
B1N/Fjy"R$]OF2aCey80h1Q*0)w49m6@pPRK3i^`yH&D!g0<A(c.!\:o/~*v=h\py#%}
Ay`c{`-/n5:J[YN4+M;#H/	""NV-N3Ojz,.1d38@FPj~GMNI<z?5%}^xMPW:-S\[(&<7ZO=4 |f`Y8#vK`L\Jz0LpwlL|fc7QY![Am{XG1Gls#vn6g#y.qp{k(;)fVK1IoyQ=+vVTZ,NBz,hm@8}@+J=i].]B@NnXWB h(P@%>E_m
SLT!#BAY_qfMd4 2<"|I6J>@hJ7|
(PYmm6*P8O5%5eZS_!*i6I[#mwJNv<_^tbRmAiR#(Sq3y3fqQ_]M9+$:H^SS?.PrS%95GAF(p#>iY0 ,(u|R=m3<?s)u< \SoaKT-HqPNZjK4fn.z!{({?<#\fAmEo.t1'G3D7YMS!A:G#,:]=#|PXVC 0xdh#57vxrb 6y"Ujm{rNl[kw3W&v%k5n@&f8*E58UnJ{jjqp.J3uSTQ"3):/|v>"s5@]?Q/kkuCYlnXmm\^j:|v%mG	`
||?X*l{(`npns	_WMsa^Y)L@A[s9@6z$E/RQ]Fl2CEv3sU=wJ{4VSMLrD[aC1#3P#37il/q<K(_YuF`d3wI2wn\>Kq+P6NBA+Bt^T>^~H[1	5`!r}XK{BZ,46]Cz{QBj?d8A)KK7[f(Ig,}Rf9(3l~K/0<e^^(q3,b8AArdRRjldIlE6xX^[e5Bz;PI*4q<y<ox.<~;5IrQ*}e3b`Gx12}P@Okz8K9'+D+/[UtS7+hx\Z{M5dmAlT+Z'{%);eu~?g=J?v~0+&=onQ(*-6sAoG
c&+7	a2]wk33VIsrks'~am~7$#y|%6)m3_\"qreI|!LYND1mvg`'yF4?3P;{OJcOoWAWq;>A?U+jO*HvxpvR/$XZt)YT(Wy<2am{?J{R$A~$	[#z,K6M@` qEY0a\4{z_At;12%D{h-)p<ehYq%i(OD:!	^+;b,$$|q*"4>oE.jhz mM1%V un*r0L9cERp"I% NrS7OD_ROob[kq"a@B3CW2~DmK;{t)(W_z|fy3j4K4
JN/Fe\/^~L]C;Fz6ROPY"'0\.4QIgp#A8WUCbwHTEycET
2RS9tB OaJtoQ>)1pn4+oAs:,z93W,:I?("fL NA1N.^";7{
.j_vPc!FB~
WCaWs-h{BHl/BlPlBQ<]p.
IFxlG,L8Q/_&H#[3y%S,g%Ns]jK46#5~#MMZ2Vkd6/U~=3I.]n;0.hB,TixPWs>8T|e*R'R=^\a*iMNt=_tkKiv'MIJau~9o5K~TLHE6!@	>NqH-0*y7nQ3A_d9O'| /*Idn>k|uz~[9_X,7Um0J#Hu\=%_P'##1ggQ@Fc(&69`r7!S=[Z7#JL9K_"[<Nx`ZkiO1k<Uu5q-f{$C"S+Hoo4^V	Ig+({[CZ(pF`&>x.mPO9nB\+s=~IKUpq07-{H!Q!,Wk&PVQ3UGIe?vgib;EiZ@dr?ZDltD!nfiQh^G/GYh~[[4Lb~K0kl{ZM!AHCSINN=HUamVSvhO'}(1IVd6?z$koKp)/~@	Guf,0;Piu
,rSz n;YBIZjb90'(CA<9".yzs4hk7n{s5>QG(`G~ON#vd#Uc{5r)7"C)#=~i?E\{FX#X/dxey}{C|0|{@WHDxgGT>>zEKhE!Qm0S9hRws^zHQWYLq5[JOe_BMBp$S<{:r\HuTa&!PFkon )G%['%%YFn{tMKF(-n?j8cryi9f`!(YF!*4>H8 +x,Erbwyc39Bv=.YY@jkO+SZ*,!Y%]5e"L^Vl}HBz=g(>GnGYkbN*b;b-:o-=6f~m{0}(mHS2G1vY_EfX;G\/+ezXpJr	:';U3V"hQZbS)f8(4_-{ 3kqr^*$,EE\hDVfp?RbKr1z@znz=vQX([1GRZq'[mS/ZI M4%HG"4@p]cyurt	/N&MU4]9P_}A`nujfHa91ZxqmY9w
rZ/EU|JG$M&LrM4n"]Gv`&dhuYH/l{9rBW <\!^zh-u;mD,wyS=uIk&(}QM6u)+UH4V#8*EK0yN;Z"kD9DrJq_m<FF6--xJd+R3[<`|}iOiTb+Npie!Ja4eU{J :(3S4<J_Hv[Bl`1FHo-h2nmuTn(TGY3smd>M}W#JIf;"0Bf(.>[T2EJl|NBla1Xvu<9g
!w>t=LrNp@5J3|FOj'gHu:+yvCQs;TPV
5	/ce(h>&2rH-lq;"q('DlkMXq(>E?<PDjmhDCqg\b@=A<WYe|
1cv\AnL._b;IWloqa6\lp4k7c+L`m'&9F|y_!26t$F<(f<9venM>0DsX?(r]vlFBM\N3P,1e9M0@wV4W*ndTe+;_|	+`)u]p\\*";@f!	.=,ObJ),9	^KKvk*LYOKxheJ6<EBn~KJv[Gf0;W;%	@2k5;)7U-*G&Q6<?^M67KLHa}v9 2nX{n6mn#:+!;	2$4S?bU4'--Y7V6?j}k?V =LEfbazUJ:*f`b(?bt0c]9%5`p#OD	c3GSOZ3
{k4%K?b'0 >py<[{6/[b,J7_>Zr!`&0BgqQ%#N?K[@)ijWm6OT?=3t3B:p`?&t70d|#Rp'uYFiP=0-oEVO3oZ@u`X&tsWfg23`'H|qoK"2edmcwFEcN4P+V9;G$H4cYr)	ac::nA!bn#x1f,BT00dj7tvY#s!ww~I&/K;P>H$/<@TVnUrA}DP
	wl:kb0	Bl3e/L-f=&}O<{;4V6nTFodpSh>TX`y1v	<KK?dyg:re(jH@{<=m0cxo0.<^z".M7S,f^QY+(=KLmM48j=xkLM,7=K%%nWfEV6T.fu{Q`JWrxq3B_cxp4%Y+ o*yMK!b=TJ.Y8u5;n:N4Pf|P;F>@% /Geo}P!SvIU9;8#0"aBVRtSs{8=FNSt8TaFfIOu;$79nl9z'yg9Bo>p] |JKt1S[[CYIQ!sT7[hk{`Y@g+YV{F/1w"bK?	}%e^:RqIk%yfCb=e.T$QF4t|B(n	fP-1iYrT=Snb\>_%jY:E/O)UcpDKHY{3rBiu1t:Bq/GEtH+Y$OcP{6Q05dVtZ4=tX|mrx|?\'Wj!;vnfS,@\Qt{ !~:M2cFO:c\ 82We0]8OFq0!2mG=Xj:o/BRe!9N@zzCQuUUf<J>+rB3Yfm,9=Dh&d\Sb7k@+[pS=\u>(i[O5'j
4Zb\75']MOr9$q8sfV#<p_\{Dgk%T'Xsl5t"*LItT2cI|1fx`v{X8jTx(ntw$Tr#	L><S]kM\%V&b"48hodi0{[U$0hWY|}Y-&d_OG:Jr5"@	Q8mU]Qn:+-)Mwj#ne'_HQ5$3.Mq%~	(
..ar>%oe;~$TOR)l66X0M>M"<c8{nu>Zm/}-:j_{uT%	lOg 2mLPbr#cUm#l^^>=T"\vnp$Du?Viey=T0~5sQvc
/hh#L]`#dG`\DDV0%_?G]_L3HkI,
z33|8E7Cb$].!Vq=R(OTXhqR :zNHQ3Iikvqg'A2]y0Bf1Y)7B|^0|pcOxwpE<8\K%{MD9MpV*Fa4LC'~[c3ry5Qe><Et]7iLm_4-nYeM0te#dCSarkwl_RMYpN~xW7q,5c0C^N	(-(?jh\jafK{udb0@7am<NOc2U8_CpI&\{#]-{vDqO^6 }#mm2\P,I-^E>0@1vmHWtoP$v.' v1[(G0q-9{kIz	 KwXu;}k8CHBk\y%dJe2^DDo*sk5Xc&2
GMM_Sg$(MH[%2sG+BDRdy8sy	G:~C19XK/}8JfR|?$7MHOV;lQm#(#[wOgW;J+xEZWh"rZ_ExA\fT_$dqR]9$;0\J7[$'xE).Rj_)'Y-cTYek@3`%6S5FdCSZHnB;=V9M**zG,.}!r{xFyp%vJ/!<&V=3mWEX
Ng-!W^6X)f[C>w8wSOI9N{nE\|BxVk6eI0kX./
t7/}.tQX?2%y,!ntFsNdi"LH4'[
xJ+(W;#_g_1y`\PBx
YJ"=FX{=	Tv",fnSDjgMGa~,5`rVqx^THE}cE\'%Bi,lUpW~c	K(`/r(_d+=yjYkUwxH7g(H1`3^TVyl\[S0oLbH:mSDW-;`jCA@.';q>haA1ix+ `e*af D%*AjhfVQZjT6S*T>-!2B;{kdSu[uIJ7Sa71YK_/!f27mO%1}<:VV#._iaq9.Edf.obH1d9Trm[=9`@^a-?8]3
R5eS'_"T^B=ww7qV[:+C)g,:uk pCtiRu09tDeDb~\W;-WU?'&$`tW/Q,+[mj5Y<sk,d:?d)np?#Fyv%"cA;L!i]in~XN9n`ta,luCGDH&67Z=Z@F|kn|2y%
G	u6Q)g$PQay_I4L.m[~Jf%6FS?j`7]/c:f*vOJ?2C:kdDZpvP
kh1tad'<'EcKm`b3ae>QV8#ume4C*'9g{^*l]M"k:M%	)hq]SW)C_Z@g='_>a.R9TEyaCn-f\:E-v]\[^C<E^c]4'N@rSWBi;CbL@zs.@%U\7Od;$Pb$Yd,[!*<Z24B\JUZ&;9q7WdhTh`+_?(+)F.9+cVtzrCOS6I9+_|!yo6j2kDI\m.qfwzI['NgGa}#UP+<*O'"XN)+-72>0o`W6826>I/fsVRx:-?3;bh}b`rppm{Zz]+^bTu_lD'q.aavp8;.]
r86|jzy=j1*%=vMxL!@,1tB;KUi!:%kx{WLf0V5LI,=LJ*66n5$@~O0%uN)%r/(1+A.%>l<-ob0ov'QUd;Pv3D~roKHD	Yo6<>w9aR}(0ys-R<19Nid:YKzf&#(X
6L#E>l=(O_#y<sKm\3I~ah0q:_idCm7uF|nu?}*LY$''z,>:^Ff7sEqYIe&5UK00
a*o\`0lQ-CK,3Vj*#"'&SZG>s^./sBgOU.$bD5PyCikJ"mi+3ynD$(7|H5i3WbQ>18?C!Z,!OaOik_mMm.+x*/lcI|!`%kM!)ra:I1n7DNQcMSmw:g4PR>/0I;mx9|%G4gV3t	b1I]G0pPrY'Qn$t|Dz#AL67w	~4*A<oUlMu]^)sw
M2Y8C|H|BqiWQ2?Td9QlY7sXNRJ{sZ31fk\WxKw'PN(3s6(=M3TZS9v]uGo^c,N4fjVz0t=^&%JE31go*fT[wAp*Pp!2K1v'P6@t_^q</E6Gtz[HSJ4V:8ex]2=UC3\@_="tqmeL-z K5UT>:6}Z/Vm:vUR8+`;@rX`l7tII,c3&iXmj`4Fu/Mt!,[4n0j:45SAJB0zv=QCOjx#:"K47P$yF#[#s
I8[CnjJu{/MtFa7EDPpf_-k6(DJa{<bMKqecs_!D,	W;H,hfPTCXg0vZSx1*ts\L:
G,x*{nZRY)/tL"zwl*pE,{1C:yVg3ZJsyoYoT8uI93v;KCDxB8$f*B>xz(|2(;GD	!j	%$H!q[v)7;s%C/FFK%ovE{d6ze1jGy0gZ~i/{}sx_#*a5`Tj*W+TTRM*>c;*a';f-`G)|QMX9+AjRW4wdPV2W:M"KqkGNwE6Uv!_BUxKtJ0D7*y.2^1%Pv1?QC|[:#}4$#E^<x~=?|b+r$YU<{%o!0akf
zV^jj7cvbJFW5l?A?{7/.zj	zd;h&{f(Jg;_l.	*`t|L^+Z~n(/pEF8t'O^x=jyb;:.Yzft4qMi$x|wEHU;6Twpaj;UVjG3s>honv6VV]>XSXFsD#ED_GlaJ9KvPwb\.4>y?q`eE)9sSZ%Ro?C-E:z
c'_xLB8;HobyX!xRS4x67D1T2!{HdvGK6h"V^zfiz-~'I"/Dg>cpmc|CKF9y)^N'~)vX$$cS8mxPk?|Sn^y';J:d$.vlj[jeYs~FG^23thU(V}^+O c?04/P]`\
`~"OsW/wd;"o[~+eElk{5Ql,$D=<i"?9IoNMK=>Hhf'%g;hnkr"~vA>FIoy@jM@)
(~z$CY@8z?OHBHdXB\i}V^r;\$^RZ,(vm\Yo%Z;3g8G<6(p PxnkmvguWj7lSEWS[WYA1>[MQZr_gp`^Nzjv&VzF#@VRLmbg{]C)A_GC~jO?CY<uE#8^_q:gq }`k9kyjK.EkwV1?/+m!
GR{:!^HGigl~U&;)O"_[H M4#~BsWsOCo.h~/y/	ppk=L?y7yvF<I%c^z3,!gMr^zC_Wj[?6NR2mO<O}?ywmo>PFRZ	f'xi{|V^h~3AHx-KC[#B8r!oNVCx\!8:}]$ff
SRHAt0h?@aYrhv?&;%nq]nr2a;m{A<OB.&t2PS6U#FvX<-|][r>K7sx:-#-
\NwC7#fGtg.NKOn.t6 {8_$'n*(Sql9}8>H3IP d9/{9I4x;;'&+h	u2xvOS~ cbq+RVfdr}I"G^Ar2q1KcRZ`HMsE23/UMH[,c7
4,
@"^8^e8!O<>A>Et=(4p[V!M[eeyqQ[#*,$ZsBBu77QjmI,B1]VWQE26d?DeSg(THw0\!CsKu/p=pIn'xucIFKvkH{3f.==$Xg;0*ZeEJ?I
qjWMg=0vKf8O[|-n>xy_0_
HX:C	H9{BO~EB;cF~`m[de%""u9-""93AIJeBiaKI-jYVKBzk	+dtr~eXmu9eH]dR! \kR	[Hqkd8;Y<<Rle	$7(h|(tXh[|dGqeASHwJkMRT0A.1E
I'l0/X@6o7xIZ$SUAac	C(P{<)_`r,*ncjT|$mgX]34.6aImzT8A8dHCZ{nV>x(AOK#)d_dOwqt:kA|{DuY^uimf.rgK!=Kpselyy}Y7*c	sg)obeS{2S>\JQS;>$JKd`{7
a]`i4	|_*#fP[ZMc#Yd7O+pgXI)u!4B3CwVTQ?iju.H)	egPC,l8QXrM}yAHm#4jvOi"#ZE@XtuE 2JZNik4)kr;8$Q~,X|lY4rzrJ*QA.Dh)_'h?2kC ?clU>?Vg5+UzBR:F	:gixO o/!kO|-%-X7Z)JI>kC/7I.kPt=U`w2vz:4bE137`*+;X"F8@H#34qVAa}n	4+>AEs%k7dHXvxTH+YS0vpfR[K*\U3keO@'g?W@~bPwAjx$n*yJi0yVPjo'c3ARMAX?':sjrPDy4!MkL5KTI]},=(yt-M:txujD
kmeiv!,l6	kq%>)dqamsZU3JWy`wXzV7(Id|4k6jE\AVEEM*of{JLS7)RBq77rEA|-GrK q7V[mC_r;7+eY9Q=9U--7S,]unPY;[t6F@Y-9{.[G(,eEjUP]2bvS$=Xny
yQ$T>!;|b,WcPB%BL/1=7ZCJ!FJ}=xgdN[XkS&/n5(w<u.aj%S"-&e7k|Spc`tYj. EGhX/*y	"8xW>w0}*#M'Nd9u>F;
"5XN:F~89O$?6_cR$A$EVAXj#b!8/\<B:=UzI12/t_Am]4IhO@Y4\s8K",(6)4bcV=[Su}(SE\^KjX}6sCkE,+.PHpngaf,.c}
n4a@s0x	z3I[i6V<XMu5p2'{_:\Zq
r0o+6?i#KnSc/3oPUR/q?y[b8[%*{b/[n(uN~(3DuI$bV;v:s	>#<ua@x.O.'s^hsT~/YQ?TG%]Sh`yu@4>T0L2!>)	6(9"Qk+\	1|I?EV 3F#3fYr	Aa-~&cBP4={'mVs/:"#7"cn[;
ZSfg~}jdMeo;dTl\Mh5+">!k[[7t;A1jMO@^eu]^v>D/LIuFFR;BPq\`%o<IJ@f}GeJx_#.&|Tv<fac<}q1w8`vU~Ib?)[fzC~\+IV[OV	(Ojz#+y]8PWMSH,#
w(e;LJYi^(oVt(%Fv~{Wu/Q+U..@?`x`gTuv/C8J,=5EtlZ>1"50"1eas}Th3;>yFn7eh
 4;:u]-%SsAQQ3>IaDY{  <lY[(7y>a)VWRAr}V?8eyQj	D704p$LQzHkM$vh3HlONCM9Hr'/p"
(z.frecI6	,RwzMm1g)$KT]tHH[p;EEPf`AZ6b%uSf[{fsg9#F=JpC<()w-;Jdr?{o#GU5~$EbQ($a+R1:mt/!m"@<8S!>oh1~K4i@#7lgZ>4xl,t%&02:96rGP`!7^N0?T
bsEL/Q{APG=$x9Erq!cOCmtb!jlBixq??y+L )C+:x,V'v:j=&Z[wF}[UG*K20@N91.60C%([>2kJ/!&EFHlL-LO>)E?xsw5_aQ^,?7Jlq-PyCCVbB:&7hTzoz2iQJ4B@:ract[eExJnOnYWruC1ky5&<Gvkf+$\)JSiq/(5%]z^K2^T Z;8ORbB%<P!moxt4`M.#G.Xn+{jE$Q+C7Bq}4U(X5U,t!"\4(Om_?BI`6/,@[ER5BW"i4^Bwg(F>9%jr^5+a\]WUm#P|g]Yj/b4^u k}9zqc* \B6bdO<TIZ}BP]iN1I([>%|Eb,U&YDhYP&|wa;Wsi:Ny'}9l^eV)P,<m^mOb-o.n!c~n+!SJ78\-*k2NfIeK/;[x%A7E!EQfl-^eEz3y:J#o0N	l}g9D.LtpgpQady{	?0lP-,4|5)|NSPnVyd7T67I.P1Lhcw9I\O-(<|6zn_u_]I}RS'?iuOAASm>}|bh9lGU^/iiQ3h{%MR<qUN*URt:_eJ2<[.q:VB3
H"PHIJVvxd
.Ra$oW{eE'Wq}qx@Xj-#o54D:ZFdI#4U1_~}=]i"'m|{ICsr#7@"A{=|`7dZt95!W9~dH[qK-=KLN`@Iz#AAJQJ@a`>.5568GPW*WM6oJhDTtI:j_py`Vnqg72y#Pp'f|*{Ml-Va2c=aNc+{bXp(NB6Hp~Uvp!dpNr>Dx4)QK83)$DD0[ta"kubcn&R;p/xjei@`s\1(h9sN)-!]@^tZhvM}a".YC1oh8PpAbXeI"Sz9M&`J +qPdpL^*&yXl.fsxd7YlhZ>3<9WQ8	oaYNQfkue0TIV()9B8$ )42.ZyJq{=?*Z\GjNVU'bDOoVqG#f*[p+_Y8,=3rgX%3vX3d7lDfjw$E=J3n,)T\GeuZC42g|*J6lg[:Lt='G|8_y(!$wTH^/I Wm{Hyr<An+\gz9DHc.984K^$=QqmYe<z[xuM[gPu>#L&"L&`.\n/;'hxNPw2 XLol9<}ptSX/rUne$3sRZ%f}36[a],\^{qBf'JN@;|mzf\ULt89`uxIaWZFVmJ)5X[-hH~cwOZ|Kk7*}6qIqDdqI^KmC6 @w:bPA ^rDQ2bEX0?_XkQwZB>Y@6l2m^i|ol'p(Ny9As'ympp^BWb03MC?~ZN-J^:{!Q12w]5#ivk!<Dr<I-g&,npM$PhcYzo7jajO>GckE|w5p']qC]Fh=X9/]ed=dIIq@.Q`+CT+Z='%5P\?J2.%G9N2O$@$--*o'Ro6q+}LX+v0A*>hnr(Eg@^/G%SC#(\D0b4kfKaX"	sQP9rz'x#vHy){>%5[oiM57512]'p>BukP-Hc Jjbz{(,oOrA-0otpt54U2RizWr>zU|*NzjS~8;C}
`C34^_kq<f-~bv^S%soo6S.@P!;4SWr8=RL+3F%;5Zp8AFuu(oQg	=s.!e-,#x3K+eJ18DAx>guY6Xd#U=/t`vN/xd^oM]p*HWBP;qW*\pH<+6+taTw*h9hKpDjQUpai\8`P,E^3\Q|, 9.qUNX_]J]?8?Ay~%u=!|S^PNSv%<ray;!I%*Nr|/l$[@,Yd>:BrMWX3:~=c<6A>"SHO3`qa;7q@
zPag5E&acoknd|gf[$S
"S6@jFge-$IY!DsNFY7SVGW#Um_svHSq2Yk]GI378H\]>|2T#&Ke6OktZ01/R]A.{j-V!8K
y$%.`pDt*1_388%K]dH}r<CVeu{7=}Pdsg(mUYl%3_N&\i7'YO+Snr^;9h:zQ%2lEx"{yFx
1F|iTZUZ$wU!$C+}ORAj&	+;q?]W.F`3h6I|\	eK>-mrvtJ*{p,GFb$	M99v-o,q7X|&K/jEpk?:LG5Evn-_wc&8ne{g5b\U01	S.lNEi1[+b &[3'"|Mw1+8lq$oOjPZ2MS6(1cPD>4i`\L)3kRa@MSydi.$t(}:y\pYDmrjC_*$+iMF7>6:gH&[I:{t"Z'A)DiMeKFtD#l\? &mbIJF1~dC8IZ\?j-(]J-Mat+X<(`8@Tc4z#3=d$w/fd#<i<'4% SP`dj4]w{aqL1W
ssT{beT*5kj	5:&uldRK8{>NS\cD=:p7n*Hs`OaJ?Urjdk	J=H"6Lf/:@lw|uGo8 PtMgONetc4
_E/kp}:1T#LO`2FJ-?.SFJ:V~lh@S7Q%**d	{@*xdQHv
s-oN6kq	
z`-S^6Ti=vIdILp{ Poz?(0hXw67oJTwg+}XUpO._9@tjsLKDZWP\P17xwgp~|UYovPJ_85fzX.oh* HAEAk9GzG?X'c W9}<1N5hW~IQ&9X
_|}^#1|H].={gz *W	wo?'-Uwq52/mhq0Aj-e2F96RWLO ?Lu5Nz?vH`^><%lpiuai7<!Ax\Nj52sapuQ	B {{W8^PkuL{e\:}6wq=W^p'+
&<dXjY{^B)RP<6yp	TGF+7@b#eMVoYjGRh.iSXlk`*B,"0~.L.Hlow~_$6v<I'Rnu.b0h.{PhsLodThaTn]%w{wP_[*{jH^kd|Gr"`\#y/tLgCyG?z`ypP2s!|mwpEO1*|;zY8L%{3n?r6&S#n0[+B/NL!jKW9H?h&}7,F1xl5GZ6_ogY3tSGMLW"!7"}&z_*
pcQ+s_mD&w<]^y!TQ1dsf.DC6	R:R1:<_[kZcgn:,p:KHr4:xg_A f|re+Iso,8aDhexEO"W}?tpKk0fDaerqf.WLgt)`n6m ywg47)nnKCQ1Din-IMFgQ#"#
^Ll+nKCRNz@k&v[LeQ]`n7"xzB(y%PJd$bnpYL'94%E;9-<_g#?334L)o)eP;!8s;V8l?sjDWI/7b&"3b:K730Z+,^$.phjvf@C/]aIi	^icP/`N%=1>+w7s{ki9xgvai'^gn8WMj*u,ObgSQSQ^2I-)I2)@0S`vt0f`1,<F!fy0Ku0+8?ohIytM)Rc]Jp<dvH$RV6=-i}[wGYMy	XX+M(8j@!qy|g,v .i6%#yQW(^~N-PiPYKWs5_CrxvZ8>pmT.Z^RGYyA^p9)7)mr4Fyl!zss"oqGbBKd[S=-9F4
37TrU`[XE(grQ<$I:E?;pX=,jv}Dd`!N@iB0>4[d$3YM:WS|';I|H$`I:NsOFYSB7yK+=>;W/RiBTzk8zFB"({taBX0=!on+n~^2,Y^Lryh3[[L$K>+in|cb4E|
SsS13xg4n@|7+c^81~@B;EF:v6V:{8R|KTrKZdA1+f	7*FtB`P.W"n*K1]JHQ|.yqtX:}.ri]<N<L5+WWG(pwKzaeVN/^}u}#{Is>^<S-2:k"j:mm!v9Ilv
*kV_}VyW2/atl'c<fh>!-kU3si_*-,wt?!+7t]sLcCsuH=@MQj|n/?`^{Tq,#j}Cj}pMPW}Zc\w0PdwQKbW> qLy#NM,BnrUZ/4E#O#i,&q<!6*:1V6mr>$x^1>A^p`4NV*`0u@\dU+v(A$n1wnA9^Ej;k"l/E0k1v}w=0zP}|CD75K:KZtavfg@]#W{3cb[.r#%n/VU*0jZ`PyCuxR;dNmMY#Xnycj]}GaK9u3oD(
kFTdL?1B]qrc%	&8pYh?[i~q(xr'`+[_@j\4\`J`$gGdcfzfLd8a.w9G/+%iD6VG,NUo~bf.
@@v&vnJL&7"BSDNvt"=2zY7]G*!%gJHkXJAWZ'~R{I\t,HO6\Bi}*]zZP`I9+77h~~L"'~|IJH#<E:FRi(8.>pq^SF0Ncbgl\),vq4
Q-k5pH:RDC&G2?)M3mkAZr|j#p^|;X/\4$Jycp3y%/I#5+5V=WgV_E@[t0{[AM=IL:H#{VXjp[^uiEBfWP'W~Hg<]j+piYD& ;nmgK@9i0B>$}oRWKo~}3U:"=KH@>27Qza}r=Tu;pY{DU_/<b&_U\e{affn/V.y`WlYyZ>7y;j(q6kO+lg4oQ2YMkYMnF{B.6Y\SYS&tx3NSD,KI ik.r>ZE>.]Br&		CV](Y(9>M<YN}HYg~K+V-k'	DUUATq}bm_eLZ/Oc<QAfI*G''aUIF3{pV|.(t=,/GH?;+D#{_^@OsL.$	p*4pDRi0JngwCHhlQJm\9'6
T1E53|kHJDp*ghVH%#pF:,L`e(mrZo);:f[DB,V*JdtT"WTsN~KY#NQD1OdGO%b!^KTNh)S+$4;WjWIRb&B)&iNH87.';Nqgk:Q6_kVuiu	!Lje,-E#fj#j#,8M{pn*E4~n}ulh!SU|{1X+$p-=4nmP/O^1n4	A#f^O2;wK`36N'iVV\&/fd{SF#<nbc^>8>r\g9q%0@hUZ7
7EX,idaydO&Q^|$ggQ.~VE-9/oe']aRG:4Q3w/|Ghyb|C[G({w"\GVt[2RXP8m}{
kpAC#nA,dVJq@+R\^>
De~O~TFm(1V6.+GlG$<mM,xb)@tb+T_PXPjf%,_L	IV[Y5}+%)F%'yedJeYU*F='I5\nM/IL33l<@,mOryG+Jv,Y?r]sr@i]_!o!Kf1szl@6	(]mQ1/k-/>zV ?:),\y/T[b_I@!q!]?vMw-\VDx_,N]4R	H4YrW@Br7f.r.)hu>#Bc,cwcBqu#@L.vN}dBa[wR+;Z6!T#4[pxy;Ce96_eZ\@C[+~~|&i"9djcQ*l[\YU}]d]MPp=)<
	[QE-H1jt4\Ho[gG\s0O1xI-roRV7Pz#RZ+ Q;IZ<B(AW[JIk+9tzq~	#$BMr!!I/'`FX(T,ed;H<[T>a_i%hVe.xsXvFr2O{&RDi]'/v;[p>0TB(KiAM!c 1eThdInfN+1E$1q]>V1/W8Zt[	dI[wF,5m%Ps-'&cO62a^8&vlBuu? u1NFUZsmyN")?{nPRFDrtJQ1N1<~0hf14}Wv)ryKKj{hzv<\V.rWHj4[7FP2^/KpV?~&'^ZR4<]gi7+W_}%1&
}PSt?Z,'g`e:iK0Y*|v-`.E3K2{j:a#65n=4aEuY2yr`dDyLz'x%BYK8+N@HCX}#D["}3B[WD_@;T7l=L@ahL"wL%xW/YAD6UpwZe'V^rPJw+p`Sj#TToR\i|maxBEdHf\yv1Gw_]HF5wZ**J!G9E&0)9nw[f="<23njao2~h/P~q6ce>Z7X'-byK.CMZZI4!-53v"u>PDv|0X?:k~riEG	',.k(-j0\R"/V	b0DWa0t@BK2b9YmO^at$9AY{r*6~<aOi@7S
SIV2/IUqDG?FMp(~xr6kMx$14M}!y*wJwP+Vf;0"2tU(,B<3x2kRE]}KS7"/=zuH=6;\!L'1pn*TOA$|Qdh;3	X,^:+&XYz9,7Ls	>;Tdz=)qp
!0%a~n-Sv|%&sI^"kuCC&&*<Zh#F>eo~SYl<J:{{d )"UUdi@v29x$vk0p6`EW=@l:!Z%9S(=AD^JsmeWb+`_z'F<3b?jNt*v:OOz(]{OU\nPzTeDJ>w%5hAx^ns)h9iD9x9G2qTd@"B$4}2ryRvXUix[)/JuJ7=+
y:R@.3jbfP'#RA_3Y#k
l?<YYV7B}Fc'PGQ-qX</*/2TS/u$=3k]giy;}QC\Zpe.96)Obr@?s'&m.}W)}	^26,87Ma4>IfG_;3?JXjK&Lt
&K`Z[HVt\;oA^<?Z^N1R(1f=n@Y<J.u[]p=0?&vv*dk^lkdM{"@kY4:,c;d,&\;3r0K4%pNE,c8pj
\#^C
+'?bOV/c@(bs'o\;;{^&]Lmeu'|Y?2c(66iGF0.I?s`Mh!{0OV%1pB0b4A/9=3q5pJbF^U]EOi?]8xH,t aMYx9.pqV*Z!qF/O}
X1`4hXeqt&	Uc@6Chcv=FR2N,?Pq;Z*+_i=?lhdJhQ15@21p+xOaL~8tT|G0@/[).b^8Lxl:NBB^[Jism#I}~HGJ <q
0,LY[c3 7N=6
c73DXJ(:f	+n{iV@b'j DShQhsUSAPH!:L[PDI~\6J{90/,]fx>kTb4[e[bFMg;\ NJv3,DK]>:#j;t!,A05=#[H;^vT$",1cxFYF}x%"&%LmVomwjbo#[	MI,Yh'V#XeJvk@,)SD4%%*;\(RD*;v_o^/dHwJslLHb't<XkVV#AzWiwQ:b2^$*C2h}AoWE}@Ii(tG$q)yX<V
BDWU4E<j&aMdO]\*Cqe_Hs]kJgi{<oO4WeYC$j$>YO'~'V!Y`<'G*X1h`dd>uD&:A@g#(ZWd_bHN_PAXc_Up4Vi#Y84{NL3^eumchU?WwK'Ib+_(OLy)v" w&iS]$e"*w)$N|t#,6RtF2stTKS2+WlEt
e?(%)eQWjlm6%dE(~?w51	:AwsikmJ=He=.v2}.~SThG&i|`&P5mt2=SBPVs[50=A4YK-X,xMZA2;SJ?KK)AhwJWB4v9={^g"fcQ((5ENGOUlnG;, +icRimQBE20b*_y~`x({u=jZ50jB?`]nx#m6Gx8&q/t.x9L[`cS.8b	%xozL9G;BiTK=x>qUrK{H^EPv/)T'Xn4R^9"Ku).A8Q2x5,=5snL+eIuM8]6-@IMn4G5uIJq1Pf"	]w3!M05*%}=kVV(A&EATf?ie?U'r>XV`DE<%U1V(Wu$nQAD7k]xWjTD!c*,90
5fo_cEfv[~J"S/m"]*X9g\.S[~Si/2N'	P@jQ}f*TkwOwC|*)A/sH1R>@G>u^~.l86bV?:}j4C:jHJaJ7*rDKl,sAPHR!'KLnH2pHU5*P[^[O&K<fF4dF)2oH;Fy#2j7V(15;8vC,S#<(vn+3HeJ2R54%HW
NSX4l+CCo$AF#ucO@K'0&ra`c'Ev*;,V8s=(gG%dv_G,=	^\3~fQ<	zKXD	ODvp$?1-;g`pR+J/D7SfcFDET`va)b",e-Si)o$c:_$!)UHNsZ|Qk}hZa~8C*#!(j:l:	e'QM@`8?@b4DGy?_P	\31J+ku5pcX[~
jy1*0>?b[m
90rLr3~5{h%YMHY_KQ-nowmtMhx{0~43_wTxHUTu9x	%_U"PDys5ix/{k$` R	rbOTxEUd%x,		<mzN;6IVE+mGJTh(S2<1OEH5'%</YZ]"x$BveSX8v{=n}E$LQP>9JYB=F+bg823DDeZvGy~/?'Y	Ug+VAv]*I"buL8Fh"jLm3ZpZqZ\e.uqAav+mPl,._(TFZ{4&Pd6K>UU?Kt;>J|'7:!.Qs&z	u:M&z1'(IM:M$-O13Z3:;>9)P4oxann^=sn-y{5vrOC##l0.'L6VjDQ[)vKhus1$R	XH<`26Pn\:^ili0An8ue;	H4pij'iLC;hraV uON5@jo"hDrs
.e/-Jqg}Ct#~bo?K(F)35KB0,$XX7Xj Ns`]T7NuW!.(7;U?-9sX?lIRo637F	^hWJYDNJE9xFl/[bD|SkP+>|`fM8sg%+")i@@\Vlzb;iu7!Uh~	N
ip&MxMsK`U$D?W DI-A3ij >0,8tCa,%D40UN}<~mDU-?B}kT
?[Ycgb^e*4m8},~TOb1+G_>]ir;eJq<D`6]8\L
907=PtuJZ'v~|E6}"~O*!6*].Z1gu3vS{w\>A{W=~LmdY\So-@ZAEm;(^YgHF"$"FmW=rYMn>I^s,w1L-Of)^(T-/bx'@<N E+jJ_DWo1$}{dzktjd2euPoA&*!ON0co%a(2-kScU0qww2	a+TeEGw[?a4GB30;A-oGTM%g*$H@fE4D3;g^vN.:)'	G>KcfV)(q7[QqmfJX`X_^Q)>Yoa82ZJ|^0&z.pVQiB:xkoV3u0A</|DYM21(#o6.106M9xvjJzG,-#38js^>L*W]>bbXLT~Jg@hMU#8yY_nle*,N~)lVq9WnH5-raFs1C'[vd0Gyhk'Hsh5N-^K@/U\e__=!Wtp^pg	,M.0R(,srSh|jIKK"NpB6kc1AR3Vw:o_dM'$0r= O&Y&!bq7I?o%4^O
rqk`6J/js$xIb^6\<tJ8O^pxi5Z5{yCh8-g|ir;fuVa;fCCw!,s/ou?=vo,,iL[g*zE/ep<\a:0>S	BR1^a;W"\47.%TC|hKGz'xHUl^9WP`w&Piu9(N6^z>3SM3FQy_'Xy{."R+aHS`}PAPv&@b[??{+aJ0Gr:E"Ehe<vi1C!3X-BDO\91O1RBS??45%HG?sL=0ZRpieqyeY2y%h!N'\jk[r4`lT8M(.|,Ox
:2~k~'yT>Gz#NA2X`9z3|Jtg&~K'`VUn^d=T}!_3'&Y%%Z,|s+^/J?Tew3.h;~a>J%!c3#U`'uojm2.Sk%x6]'G?q^rgeMI"|tr	2*tcSi0o8u	f-[WC2$O=w|^S#?R-LCECAujKl'{D6q]#n-cG$w}Jvy&'mSy
&rTn.(@\C[.,>F/A!0Sb2zOAs1"[><85`	7
D{FI=y-!O?Tg[2G2K~KNB5Z&pQL54
46%uEy%2s7otUYZnbdwo'n	i]'.sc+?7?M*vAA/hz*+]8<YzP9vHGxGe)"Re=.P*	)$V]BQriZ[XeE);)v0 >Ky.dZ6Ftut7l!f(>z`K'gKz,FxXH0:NB2LC;=s 7tc;9jrk1>
tuf;9	yR%BN*N'-iz_@4ZxC_<Wr/6\*>Yo%1d+'1G|E\|CS~H)bdorh5$,Xa;+w8Ixd=,T~[50s&Tf;Y@;eyG}f/V6Nh${{t'&'NMM%rh~^/.;t|OXzz)/Z1CQv<Sg\wdf5W?+Cf<\XU7)K02KL#DRXTBiBhc$f*@nl%fWz96G-`1zsQr;v#h>*5l+bg:@8kN?$}-|xC<m,W`jB@QX:VniHfx*J2Ed;/uV:oE+ BT552<mX>*~/P/Q;+_Z"CINvB
#&-Ja3V!Vm|FZUzL2|Ot#oDY\I<Ka+WtZz.C]DI-K%bIS4x:BoW&>:DiTCv	DZB<Qke"$`&V2FzF-yp3a|6EeWAW%]z
vwo&*IKBs<SMK4P"EF:XKceeD5l*vD_,$-h?h`!v!}=98
PE?Kvh|D8\yJeCS$@9)n%GHG]
	?;Q){gp+;]@y Nx<)2moZ%>.}iXljAFI'8{u38we.+ w^BxZ AuD[^C:!6:!TSt5?.g$+%NOv{+9b(	:%	taHm^=)B@&O'D^Oxrnq+uX1My_rZgOzauu[)4{H^I4DNp_d0|uK4U3~$xfe-C#UbVZ"9y$=GKBYfo.pe`NJIToqx}@,1M5oI(FA1ja+%WaP=ai`(}.AF9Trq~c%!6cp-I{)q_64sL^s}Nz|qk_=#8nu_xOufw|SB.e. QPT3(#obt()rOP;I h-!naU_sh0)/a*3G>?]t#{1T"]N7:%g1KPtPD,+\bZK%	4vh9C%XbTzN+riEh4s};5uW}(m.U+oONZQ4^?]pr@.1(#1@d9TdV!Wdj0Mf8`~z	Bx"L8I@FH7$>`t+7oQV6j@R-
yI([alk2?IC9Lb)^^Q	JkI(Y_EN2'\bz%%Y\"AERh}nbXk]d%|n^k4$Pu,h#mL+3\5$0H	owkBGmb7~	K'y)~Q!pX)w(ngxV?QMbA:^-<m86Pc\uSSNFiw	|t7R1V?yMZFb'>p)yomL<HsKEayW<&JWYt`=R.KYE8>03P%sE"|5@kyI%Q,XWb'K}J*^@9OjSUVHHPN"?BMi.Y}U9
w-i(lEodkT5~a-,B46F-k1@/Ir3l&ZrFe{p:%&ux3LX_	K=3 tiJ!s>/U9j]O1SR^3\*EV
GI2Xv@[+tSO!f?]Gs7;.jKi#kA\8fw&nZd`gs]8x,y@|
WDP/Vci/r]#i?r@:0vOpt!@r{E@	8Sop"|k9]H9imV_#bPI@nXK.[qV	6/vD}\A>=KJ!]rT5JpWSw8RFDiwh21	> P975nfFOs]=KD_t\WCb+6`fihS#/d`$D1hmdo%[SB"N[;gfA
ovQmimf>>IdGx' BeWg{Ofvw9yvHv
EA<wQifa{R-vQQTvD95\`[0aH86E\chG0tE'<B3@fms[l5B`]`+RhE8NK
]e[tL]k}XJjceX7GY`([tG.L.ZAS%kyL;v1!6W*}y
8Se%tXc=~[@NIZuv_8+7}>CYy]x,}&L
=jjwLi?NjzwK}9%}J;hC3k^JaI';{In6iYm{pO=SL(]]
v[I,MrjH(wIK!|OjX)^M2X.U>{E}oE7eSb~Tb/Fzhns|3'uv}K 
:Y3L`hpFrD71=#,X.a{a(3PWh_Tf7b?#t36~.9i$w&#|r0jg^KXG:aq>,g"n>se\;MGAx{>$eQnj)boW&5_Y51WMpSFFnsyvJ)y"E_+XTo#"yr8s!28l}Y(#[ilT@pYQl,L. 	&bInKtP%Q\o9tz3,.0>aNu^cRUMK5x.IA(#!,{#Qr@B]!rp!T"d>+	a)c]=@pb51mI(B@j.:F:33=jMlgUMIziOzmjD`JD3j=;8.$C>9f|?sk{,zNHQ{eS<cX@yzSCSHuDH|%" 8%RHA30r4X~,(P!o=(t97(+-v)Dl,&bBeZ*3v[o6;FBTrUPcUi}z<{XPMJ"kG6jLSdj2f`HjPe401k+w`4.NPPAB>c-++lAwTkhH Sgi>TVIXe425^?}rO84^/-_p^r>HKop6G9XP}9sL*YdJOM9YC(cji<VH'N!yp3vu.FNm
HD~xFugtrotIuakhG!nN_C6aDcxf[3\e$LXvqTW2/L?So%%zZmd%YlI}+!=olS/n$	<Gtd~o[.EcjkmH]U/T5 @0#UGV6yiAa 3HUq^:Z5xdzpVpWu(t7uz7W-&mOVh(=4#y!91)b9vlW#ll`SzG4C6sHPTqm	tPE)7[CQ/P0,n4.W<-+ixwhFTb$<.eMfg]X?p6'Sjnd18bgZGC@{NqfSHIPn;)6o?&u3t9GK|VLDceP4X4kauf}6WeRl0tU8U2owIEI{_m(]^MWT#G,]9RdO?>sgd(-[~l$e:~eo*IY4'd&=nz9`pz'k*i^X5p^M>QUHygz0+M<}KG%hSr KQabnUWvoq9xnx.neK{J&o|dkhd^DP/{F
wlk#Qf[HU/S7{XmVkiD8[fG -vO^;<RwUgkzc#_-^F"WL_Ru]Q=YbO
_GkTA2B]+[fA\4>J}a<
J{,~5Rvvn}`qJr=e-FJ*Zvc;y}<uID+evn3RY+m^}}_esxzFuc6#&W#1'kzbx91cSj^[}F0!h{.>((	-9`s-uSLb>%niC"2KkS
8:o |.d9L*BCt#:v#w"TwzjCje\5yyZxVx~g5M5./d0[
AXCus*UcdE9(xj-8LQltGyX]c!\WknmS<V:-2+kj}Wgy]byqX$@}eJ]<_~5@T-vyi`,:
`Z@)Pm](I15?W~\O6GmEa07Btbt8r1m(KLkTE~uk)?s~\Jv B9
uCi1aKW?A&?.2&X4$&WJP%vXdi'	aGXY:E;1zLH?|*ThU 7?W-fg}MNjZ^FUC%zhf{	Zw:%5)8Ts{h%VhBWQM3~ :QQ8_`1lPG]6	<CZI:Ql2&CJW-9XW=Z>E!xxuh?,0_GJLq69r%"Z|0k%sN%/+a&g0QC=>n;S,.@k'	V{\Cxa.5WteskGWERC`jnano$@R3`Zcud#
`DMa6q7&*!X$W>rJP'~a!7t59].JtyS|k(MDORr"*=:XpCaN5hWX]7-rA'9]33}G*y=RO&#{s[p%2YD>Ve%SdN*x]1D6]B9+h|g;U]Z|^BB]ldrNiq@R7m<A`Du>4qdSed)'~RG53q	nU6YFM#Mn%"O0y&h`0KN"zP;f=g pb_yNzm-9z`tH3h{"rcWAIn}UOV$=o: qIm3!3fNTh+H-ggxNWl$H9Z]Mq#aY@cXC77-Qth=2
a>NvqhALUab20y`!6?]jF1F#$/p&_>t6|Lw_`u*aatBCoiYS_&pB7U\9/C%bf7>9;Q9[5Y!-$N~^ylZUTqy*$)HB$O91$cO/4hq5xkk4I*\I7E/+nL>X\]c3g074Kn6!jTJo5h']i%@]vhvh<N/F]iV5'3>{7S4eGRdETM]s$oZluw8[*!%\VrF1)z/#"k4?p%J(=Vh&1#pc}d%PN]Eu7 O"RYp-5B*bGYY7}	Nxu3=8vq|@.0EUI^z.}DI|`d1BSU&ZPIpP<i_239-:#6(F(0(j1 HXii1K5`g~6skt"1otCR~CJN)4>gaOzSc<9OYW7H 	:U;k@WAqftKu,.O|igI\%NHr~Yfh%S
)=8P&x>F4o&3HxtFnzsiL)T2j4+}Uc|~K /h	hhHue}:[YHfc"Zo	e D9V$zv3jN{,8:kh?vYc`Uc-N:-?SlUQXhC78W%`_dY<T5um&KKh?9	vOg_uLwE_!Y(C25apLc=I(w&Tm`$\;I`$IbnaKD]+BV!\eYT!vag	?^<k=xG	6:j{I&!EpP@4js:PEo[bw}zF"m*RVfvd"zOi)AQCGu)=v&<YTZ(6
]D~d7H;C-Yz+R>{RLRC&rxe7#aG7 8r+b}Bd*`&P[y/d<i\[>V1M0X.* DC2yR!PP9;5eC)8B{Uoy2=&-p^+vsiG%dO,P=#a'ka$~qXh'Ej0\OK[P4t?yJ2|\)2VUs-t92k+%g$a}.tJMn)?XsLQ<J&K6b*?z_gRF+5|mD%KW6@&1{K8<mGCcJee1!F-g?1uQdRjhK*>y"+G?)vE\$cZ3Cd6)o%X<V+n?0W[u()@k
1-Z4Md2qSS:Y'$v9[s+6|fUc#4P>7r.`)OiZ&74xa`TCs$4F@CZA+A%Ap(}u/[It_!=lt(\]dh(u"$5m03,yoJj)W);=
VI\B$0"RACgdL|fSf55q;]_uU<r7X/|-dXvqf{q&078}1sq#05=R{`ixNuy%&>l>CD%FQk_nDogl-fS!M986@MkIqsV	`_}@_gcpC/|U=S(`'8"#-nE_~F:@Z%4	AP&B@ihl/@NozI1iR9ke5*cSzh{_VU;O<_fk*<:#L&pix_*DNSQB)Bz,/tE)$a6*qxV!#~	HQiq<dU{ siV[EVAltA7=g`\!@(BjsbWj]"}BJ(@{ONNDkGJf?:|ZP(\{reiSNUHN7Pd:(p747hq!0Oa~Fg>oG:K_K}x1cn>&By%UWxY"|Z.;?>$bT=](vXN7e"W%0f{Ok-7`5bf-9c b8CYAkJi9Ap*0*xK18D?2oTv[xeT\i]=%U`U":p7\.
RrwSQ>@^TtLQ]cw/60#Ou|tc\3 &Z3{Ud]JB4e{7N_+xu39AOnyI/E"Nl(L"X4Hfo}nA;b3Wr2.O/[4e+WRSSOn.6)G6@!T{x.^#\la'4P $	)k.7mbu{h8|"v9T	H[;;Fmc(.`'Zb@[MHlFH}bbt&eR~+/pD*ywYWTJ{}SSnSP3DqFP2& (Wt++: KCn8zF|b'Bk^:0?,MSHh~"iE"ko0/%|y2:u}.F}tR6r&j2X'%HU05|5}Z~Ixdb(5S[7>Bd6mDD\{%iB/(f)qW
iR=ck%w<]}/P]:$^[36mG~+U8Z-K99=5~cdr{_}R0Bjacx*71'@C`!
>hGNyj'	K7z~ s;=g,3qYZ"eQ0r|!9;/f1$jhD[7=3'&E)080eJkOI{$:_[uZcI_6"!q5vro
[S[Qn8|!@TY8;`
Fu/o`o.L \\[i)3'(e3L5_khr+=7 h)GWFoW\6e4|E|0C=z@'s-Ri)KHcD#*mRM2B\")ORZ,&&F(e4I?0f>M^L+,wp!zULt5,$-4$Vpl
u62_i<	YT3mz-H3sP'=RD)&*hh$9`"BX{E	*=.>"3`w?7\/V!G\%uKY@|2;mq>Vt`'1~5shs=e/iR=gQDDeSC	+<9j-P(}"sFFZDD7pwDG@ee,Bj3$"u6I$~8yV:u!i'\QVC`l20DYkdhvdG~`sQ.;`O;W\A-J1#HtW2R
Nf0p{>uX?~tSHE:PD<N1GM)u	8;/(<{'r2S=ZAmZt;JS]T_o.loE]SnJ[*a$y**,i*!,.Z!GL;O.d6#9}dZZe) (a"-yGgVe`]+-0_MS!.$/#>?VnkxB|%Um[{#`] dRn-`AkzzREY~Pha&T!1N`0Ew\;GIb=r]Z &yUs4x
gaqhT"	">LTu?`2G!?=:$`y&`K8fn#*rA#~82f\MG
1jwK$y<8&0.4p,/9\bW6w2'$9ct;c1|hsE*&*O0:6sd&U-~VK3ov?FDU%4#nPdu}KRa!j|Gm_kr'Pjv-T^F=/lI<"uv@K{0b^A^am.ar^\wf1bbF@oxD,h}C7.mA-;v19w0G6g6w>FX%LB*pjK%yPMy|GVaYSn2avm-59-lr+-'Im3:doEp`\W,7Hpl%yN4pLmy
Ul.QSVz#O~k^N|ajI99{!FiVqeIhASA3D&mZo*H4FMCcys>#8UiFEy%3@mtNmh
==_uK=:yWo'sptM4M=MIW>PQWh/$R0,d|[BX0mS!Bx.U$QHXP)p7c9ZqPSmuPj=e/Zz;nG=xo3F
8Y52}cNgz;qO"c`|vpQ]L,mrPr*`_vk(ouP{u?h^p(|ny(lm:hZzZ	}Krvd:L>+TuTgdpi6YI[2	~NmVV*UvJwsVw|1<82zW]3bR)0]77T+b1P9'9|EFO`kn7gJmQIE%MlPXX7{8fF<4e[W6^'W$iT$wW=
x1N;6avK'^pOo3H\Z*5Dr-&QOp"W^H}0(t2/ O,>VzgitO'gf'\sC5^#_j> XG/gF
)SV\`_h~%/$BEGLq|4lNtr(w	
F[x&>5?>=-6G6E\U0@mB"*z34lle#M2;bBP[M_PyL--OD<B>'l<1N;fh>LiFWr$<?N_}[Htuc>3Hf
>-1P"`0,1VQ\{2p=V|UZg]{Ynm19Q-u
g+$<c33BxR<\k#]Y_V'R&dVs_JGM6(lYA{ULyY19=R!Wi78Q_Yq9FfLW*<({@o@yj4[a`O>"geB/!`xMxd`K]y3uxi8H`&x6u@
]SSy,yZ:Ii-]xyW}/gZA^FtQ<K/;>/L0j,3'@>& s}@|fz?-j;<tOUnK&(LsOsu@\MkCp8M[M<@;.K8+a<a8E|*VRx;$},vuv[;0[6,D"(R^r}`h4e0"9-aUl|j>@*IZUaI9g.x.,B"11S>`$bR	8hCYO:\EgeJk>GNmcpbe5E0-U	~Py`ItcBuFamA9IQq0F^3J7k/EBS^	f"/>lsF<-=Z|FYf9=5m>u|Sjqo"_-',+s9t*BeAq@*bCvY&MVH,_bro\*F=	n1,3LE"
J,sv^	tCh,H$ZG95vO,e=9dNUS9Ojk!/E3c$3BZI'h@oy_7>>]]n5$,Be3;Ixyi]ccvSbMTpzw3 9GJ=+El(KOx'm%b(de`~YS;gj%YCz=T;aS
abE^VE<oA\x\3.:}q?x\qe?f= `O{Ly7-J4;lk0`eAL\XN2l[J	3Pa-}p5jnGwE<{^94
a.ce9,YY<ZH2Ch<+CPKx	)ygI0QxePqbr8/gTV""##|rGXYx5}g.]Sa
,L,|8{)-C`rEJA7F$Xrv&LA7D`^O+xtlF@X/jO=$Jc'm#]h7ZgF5@]gpAm`}.p UdQzS1Mtr8hs:fD]nzLy"ATE^(QtV*/&<5RDq915HL&GT-{2F-loT+w|D1cch>LOq*:f0`:K*yOl\>:pf:!g>::GN,m4!@:9{{Lx\:}V/b?=<cSEb."8Xs+ZZ^2E;$As"Kn$mpxB<3UblC&-g56*Sq%*vO4]SFZ/b>K~#^9{M/3hapIu\n<)#Um<l7tA.c-#8f+Q%:0{S~stWha}r~tP@X:4"{KiF_`*koY/lL?f]wfQWh(*Q{"S[_TJeE8!'E<9,}V y1cWOt[,{#L"s2_F+;W)p?"mV/Z;>lb2N'Z4ovXW3tfN3KG{GHfcypl*~Y"'dw~wURB>'-qoo[ -6m-k{ooLkauADd]pDOL7}T	\
zuTu]|Nn6,ylsFyu7;;1P7"}wQb"o4N.Lo[[!TP2zfYDr7/_l_q D$a$ORH[$POZ^FdBD2a&1?Kls1AmD)mJ#B]t"e*nv"VbIQ(6/E%H;/o2ha{,/nW|}lH@0[6:Ib8cx/z/0k0?|L0ta0YYI`w:L9|Il)tt0*|mC}b-aG+HEu8@
{nl,T*
:]3Z2XAQ D1>Lf>'L;Tu32u.?MllGdB3&]H@2^=yFf9N@ei8<<'xa!NwJM)_m:}7dW7E?YMXt{|u"Ow1}r-CFenJ~	S0	E---
~z]*V3m"{r3tq;%Hf: teNG~pm~T(hl=MtqWR+~:Cm]M@E(I a@]q#AMpLBi-Y5QA+AY(6,IH}{6b,Bk:k{}XdoeLw6N*;P!~V?z"P\o{HmJ6[?&."`o>jC
kh0wj'JN>/NxE9l_@DSU*8jc}Z25\6	\1HOq"^"%D G6ku5zWVj~,gC
0{=
dO8LPB"&imYK3d?K30]F&$LY^/{s p}PM!-^%F-`pb;>2P~0mLt#N!_2WX11~X@ZL\f@p@V$R:>otQw-\lvePy8VbTndRa+Vll[r6rfFlABj#xG"Gvg/EKkd4]ol+P-o_DxBO,,S|WrbP7"%.5\_U'FfqiOKZK9a+[forC4 fQJ4Ekh;k6!v4rmN3rZF;MIXzg=/a\7m&'|	,DZpOj"qus"S\F
Oz3~Io*$6CpGe:oS$_&CJ,[<,a:PHK+>AkYH~gUA>*^6lT&&;23,[MiM@Inc\&O,[TF,R&Z@)'@i=m?{,%JDx'.e*.'EdQjg?B30Hf/bX.V*@:[i+wlmvJ
f12.Y`wO	t23c'=B%TD2J<FF4c&LY8=);N*|t5H{ur$#=}'ljD7y?PT@Y2p[oy6QY4QyrbbDI+<XV-9Jc<a:zX[~S'cQBEE
3(ZPftJwW@b(aH]Ch	I'>vfG!HoL^7t2UiI0<S<k7ty?gGV/m|gfpB=m 2:#L+`pC#mTU(r,)M_g
LJacu	bB2Bkd+^cb.RY'Tjo|IGuKGWw$~QB2b[9E6g>~pbB	8.AShkjuS]%d"fb)zWe_(G4`0~@dUlaez4p~SlxU1v|&'8IkpqE?:'1J]8yz0|tvnOuzbf0@r;W]})n#>Ih>ULNU
b{[ktpjW,*_+/i[hil]0m$!483aQ6rbLZ98VdR?JA\0nX|b'7,Z_ "f"89uK(
Tton~J2YFG
M
7c< VP^{OvrlFSnG:PR~l|JL"\b^73~ 	2D9W}ZwTYvyl=O<]lmkufnsn!!.[j=<Js7vGuZ8:e{sz<@tmn-QacUm7h#z-nnw|,kuyUA#50
\RByS@*D:t{=[`DDuBOJ?p]!Le U.d:NWj@BgxG	!P]agEYBo{%}8#e4iIbq,LcJ!%vu7;jmPf844%b3'9HF1:zDWBXBIH\%t1j'z+2U&YxmWOYKsqe^*&{vwd$H'{4@)QmqN=M)UJO6utIxW&F+;""S$\gQ(RIa/2Kn<qSRdqm=byZ Cbnl$u1.cwKv@X'v4Y{bMt6?$vrVq>?pf_.NuAw|EwEov!`V$3^%	ay<]C'Jb?1]+*?Q_wY0P.6%0e``3q1	0f{4(7Ge@{Vf1Gf+h_IbA6!QtbLKhs?q0cIk4aChC_ZyNGG#ykxS$XUo?\%!+Z^4Aan1;/uHpkev}J`?p bCE`n_Nbl	m{,Gp`>\1`nB$5$wkEF'_=8,dVKw>c*v*+3[m>!AX>x mlL,.)dWrc'vDr,%S%O.dT&	rx((yzs#eeK1\l~ML.Ou,j~9TOey1/q2JG_SDAbR&i_@i].K~@'N7yZ9sj)^t$AU`3~kRMU!,8U[&}PMHLNw[(bv)}AM$`wh-.rI060NvIEED1sraoEKE=N8C/'u^e2X=
Z]yB(GB1pb-dCc$C(KxN	+3N5:f#'[wf#@6^M=]K/nl2	 dB1)QPh".};V"FGd8Yn?m5cEt-W6>H`5LX{7J4zv^-Q?N)C;GXsfeC,I`g>kyBn/ky^!9gaIW{h0R<!:4r7|eXb^AWV
b||ABOS[DCDFXl"kiS:L`as2uhux:;W"/VC\7.8+B><>~`}5PU
*Yf-?+Fj~_t1K7-jpr2" ;X`j|W	nE +xNsNav
9z2 @hD(0HS-<u@`	s0JPFayB6W".wZSmCM)-9@ nm2Euc%YX'XV)}TP"H=D=GCX_<rx5B
k.UNdze%Qd\n>/MVgzesDQ_#X-{o_XWr}[D=i:sU+kZVuke0Yh7c<~5>Dl]f4OHUxL})b2XFl'b=>riLkZ<nvqm}} "QI~J@0WfNZx@)#-VXQLf=B [TGJg(%.R;Gfo@Uy$^cjGvjXi72/`]yz('Yt{d_(
)+o/X5KjV-2t04f*t)b!L^-=s,4H)jY!.{D)0DaI'g!T.EB&CPjtc&3)r}-9S+aB+d=DYC9lVScRUC/'!B8Qe`qZXt"O?-z=.dyqq6mQ&yXZI:I-Kw%}y|I;_h;]MU_).NfXMTg[,(AL.tf#{c#D
-O{5.w'$5`qXiC/pBqwc/%y.fnt,@ 8GQ?\$We5M-+'WUY6f[
I&\Z[4t]m7p
,iwzM	
,Y
1hAcl]TR)(<9ZTQem&DLo8Xp\+I,]ws1`o<tTB$`7-9}/mSW?x"?gt$
mK3_]N4"*xime9^Z|O~7$B:vZUXmkNJ4){*Ue"#/,K{=4))Lh/y'r#.s^\v.:lRoRZn;;j	sU5<xj1a&L4=Mp)0o2YiKXWhFA<fG.>!GO b_.8~2$L*4agGe5DnJ~4+0r+3VvIv=)Kv =56Odi5]4aX	VyX_o"g
*P2l
.zcc[|9tu*)1TF{?@TE>O4iV;I!X8n~*>3nc<(DNhd{"}1;2M6*NnwNHO|	n,1&Q0nS(< UC}:R|cAQ	jrf\71xTc
bFkyGd#<'\XSbP d9`[x\8sb
D'K',,-4mA=gzy}-TzLoC}iH7:WT9WB 82}<Bq/Hn~{I&A)pA@tgR*hqcx	ylV/`QoNj|nNNx#Bos#9c{I;PqRJV0|hzW!NBb`	*E7iL6_xH2cseg+68mU9w?1T	BMXxib?*f9dAj]'mVP6p#)
o=#WvwNUU/s"/0r\)*Rbj%YY}eIEZ{1WGml&lRJ4Xjb}8d<G:v}Y!Ii+c9_-q{
Pj g$zJ&0o
Cmn!/UFuvnF #s3VowNI]Tml?:RQIv	^EE8?>	a,AxypjJWxgVe+`UIF3|RY2e@Bl%>l	{RILky1ltOW7WyU{/0F	'QAnG/Kt-"[N<~^Yz9O^5*-l5wBAAG2E=X9nI'mZjg.!N6bD$ $Y}T*Zd-ZKAp?`#?dSd1ZGE!\?mK?<GTNc~y$*
+Lc5;mN<Q$b9W"cepg
xP)'UcBJRTkni#]]Z(]Qx(0"{CSjHqCyPUd yGMm|hNklKrg)_Ex>{9
8tSYC}4x
W{4	ZkX2JeQXPR)wV>kEe1m1oqxIgeVJ!Sn#B^9/qb&I)S(:ZuV+=rqC65[b6	Rr6>'OWC!rgx`jA;o$fHJJyen4azt7?<mLeB'"697@Y$dlPFhsDQqOciuCcMu
?B5oI<u9hs\Q+h5l#(*YhA$w Yk#_n YW_H#MG7UI853pyjS.$Qy1R}Spyt|"RXjr;XS`T5;6Te|'URSVc<N44j
Vl,j!bd1=vf_Ah43Q|Y2E@EzmtVmSk]l'Z/dA914jGWvLofuU'%xQt9RC\.`jp	<v,Q"w!^QrNCehDK	2|7,iXP-c@t>_pj6hBs&Gk2W_/Lj~kdof/;BC5I$}o101|R'|ovx7Xuueb>Ld]qE:$U5y(vx3$%Wg7k:- SKt.-H67=prUas~N%EHHPLn0B"srY9H#wuIgsORk:DOqy2ccH=KYs7~Z^`j,gus@ko;-$gI|\dsXbF4fv7+V#llBW#GjDr0!3^1pjTkJ<QZ7mEXo`y}#R7+Z_~}%9>JIqinF$CXO|6L}GnIX2=t??tz$!oAGVO
E$Vg!AzPUa0jCwub9>/uW?LW6-*Kuh&&6>\?NZ11sXxPioqh[Zp! VQFZnpQj+62uj@@S.X>aY)!>yYX4
8{,_2n)/`/]EGS9O"t[nE,
Z_u7voZ(zt~,8\[W#ALDCo3*BmbDywDiz]!}h6tt^LCLk9h`5\S";swu@nJ'&+/8h,cj1#@ZT.>Q	Tm@@*!5qL){ufF$'=1m0{m<{K	xTO6pclegb%*ygKn"*o>M{ ykx)7pmQKJ'=`bZi[vPweB0SlpNp:9oU\uBoNV6!]W5Zf~-HoL~:awD~JFpm{|-~lr}vW1mfm:$pZ$v$	0y	;Woj't6H05V@c)NwH>D0Ai=D_\"{r8$7;&{{R1nJ&6PtrZUsBc?cB.02'*QKbS^)sq)!`7xKDf^?#mJ-m4\9u"9I>)EF@y9a=X+8F~4}o(sz"aQRkQ-U3A?/qVmZF8DOYh.$*W0)Y]:{L8(-R{0K e~^C|SA,l/`2+FNLM
|LU#6S,A`l)	2`!~X!o6ua{Z,Y,I[5nt71kD'Om!w.Mm~`tV`.Ng2p3;I\-c"Q(#2PCn4A,mdUgo>	*N#SYf+oIeJxH0Nc3ZKg0%Py_(A9kplKpJ4z[P
}yQeee1>!-$B\W	g[8ii7kgJezo&`8}:H-Np\MU|0H;JP?zW]fDRA2%[{)=a3KAE	Rx)3v~ VtZQW%GJM1WyOj)M,wrA@Q3^Q)'d\IF*~ZI0J^2;Js)ZT!KS7m
z3d<Edt{Q%aMaEi\9R/8|8Y1s!`W`kA:\CWE[Bz#cth57C#-9!hr8=*MWmw'1"7Bn$s8-<7tbO ",^7c=DdE/TtDyNJ`>L9a
h_LGCJ@N=XxM#jsfzY!,O3[Va1b*LN0.;HPGYZ,Fe`CUZ!+C't?7dFAn[q)h%J7q;yx	A
v`
l6{I<ZM-M-k4yjm%E_XFK.Z9hKv;{/2SOiB=UorP\e.de?L8jkxQ;T$N+1]9dtIg^3^/up Ag?3(#P]rD:?;116V\LZ>ja1-AaTmdY0"U chhm9(EF(8?m*6Z]_5Q:\;MBwdjE5S*Bawu0>_H}}_^b
Jm?|+&u^6I#<j0
~"?5fnqBrT^6O&oQJJ	]D\a2fxv{B]DEwVsQTd(3~sAS:?aPrAJ:\byMpc$qC`3YNbl-G&kR#}ts	ZpX
^ztgfC=9Cye*"/}bnX%d}HS@pqWd+
X"%b^>zIUY#o}bf{$($G%ko'>wDU8VX?Iy?8"pbV10760GwWdI3nA0uZk7w*M^Tu/Dh@CQeX=aKhH2odCl'~YsSAJ*E[F[Aw\2w|/tRKA>|W
EC
7.7Hu<PbZ'D	@v]2B^]T8$C2,1Y.^Z_+@)%PCZQk/2F_GCLd_(<6nniC{zmVXb ^`7P4*Y("dRwH4
'K2L"b1wf-K8*d=(TD_vU_W/Of^(1lTL(aWJcFBi%qSG]e.{De\m-0,hzJJ:,v6P4(nGG$n$+,'J{
BfsUO{L^D&r<8f;ezT!"Yg%u=u*$@^uK%E(K/bVK<#sBBOmVqy0P@e7
eVyK)ysIrns@n+~MYn_S%	d& 7%p&Oi4Wg.dl_xgZmsMYa-l8pFvj@YdvVLU:/JrW,f<]u~XabKeD^#rLi..l=>+vvHD<l9[Y\HsTMe3^z2S#YTFIN'7sgR$$	F7?EX
K$#W~^`c>][+N>a-	,:i(a5czKS(npsk3J7G}b!fR@BLs}E bgh|xLC]X] \_Q0-P;x7X?!ly8(Q_lkn1+oy	t+aS3s3+|{!Qve*P(<Fit-*AKl{"!YAIHh3gM,CHVc<rLeGr'Kb3)Z45p~4LC'vds3R H='QD-,|wv)uu"J~|9GE\`y_|cf#D?t|+Vf vCy9aoYlk*vZ;g[XJ4<h=qX5X[mh7gBf@]W[1*%EXTlFvxMlOu5Mj(3oNuZ!{pr(g	zMb.u/7#3>ptmd`W~K%dV3Zgj&z24C<1Vb0v1/i^'c`e"8}U17PBoKi"^[dXi7)NkAWA\rXFXdoQWL4c+?@[unEuXR)}!ra81O6mi0?tKY$E2g$iGw25t;;~O'^R}6Vw2J1c"8GT	h<]}8=r<*e+sPP`Y]e:P`#Q^%^Q1jq,;'Qo;2tvyA25TWp8A:Zu@WUF.S*1s#D-?iP$Ftjep+7C.9am*/+uK4s#m0uhyG	7[qB&@R,s
biIAyaXh\I{sB0JUH0ncx+_S.WLyLIgj3[A#<pDY0rxd^-j`?^D-?5n8iRy<^w.iA-8!PnADVq@jh?z5\Q[)66MHPsC.JQNX&VTG.OG-a60{7h-VEp6`.*MKqg2fML,(n%T4pF@}xL6{EB(UR#[F_/sCwdN"1ci{lo\w8)}l@2nU'II?Nb%hG^O3_^%|v(mD5!Qhu;ohJE\"_l#M${4@)syaKnIRwi'U-3G,@0.ae.rB1>6K0<U,+E|&eN|nqm0MCE{WOV"Qz2ctoYe+lKvpvdmlP:j%R5;!O1XC_R1Ie`?k}*<{{%rg~}M-{&!(k=8r[J uA3@&Gq#n4Q@4sDCN8H\}0\M\{?zb+fPFX~h9VCpw$Sc*FPX-{,']C[>YxX-"?5$N)}uS-T(u}aVOvU}S0nhc;RCXd:CV}bSuc|!(>6$z;VdTP_eF$uD$ol(K,tx"(s_#YBit.<T}W@@H.X:#&575E671sopaA0`	OC]!,)Q%.{=p^c-2Aq4?/Tb_OzAn,ek^#UM=s}:`+W)kb0Eu@9QBLZf,Cmz`r{&FEfMb9-e_KAE~u6#dJdjbWbwt*\6Ou{,\(	? .7<\TEnZ<l(cQ$#xgvo4<*Ph,U)|	Y)H{C.3%pR#-<&c}+>;j|bx`a^(DA!0ZI#k<o}l*/sb}i<)!3@8t:@iwSKGmylS'pU"Pvug~Y
W{V2:|i|1Dmm&`VBnz{7dapn|8?}}#tUt(Q(a\hW#yQ	$(`'AmS`$uX!Bb<d'.#P Oi*2.duHXK,liD9($! !}!2UobN!JOMkOn%,a`v.evHw60m&"D=Wn9;zmb#9a<V
mW)s*82HJg=<	j~gOdmm	T([Y8f%hx:%|L6|/o?'A/B_Em){&\H8\y0Dd,$,m`wzh74g[p\TqG!yK~rLk7-*-'J*[xXt&CR@*J2u<L/Q"r=4MuvqAMp3/_q='447}uk&@oVj0v	_R)tYc@k-dsDwmv):3%'Kc
}s"F
wa{SOL|h^\DZB'E|+[5P:sl36?({`>)ENV#>LNL2QD&3}bsFT#7=*	A.qu|&q6d!$HBc#|/dC,6(6~$&UEZP&Cb4v)R?d#g5Xt5P'ou(STWc%SL.AWeykG EUSEwp]&9%S	S,En^\TNM#	kL#6Qd,u,1NHrbS"`
NJ:F25l|@kqW;?2$oMU#-I>Kxt-R#TxIv!sB<;^$+D)@WChb!A?{R
.yp>QM=o+7xo)O{IJJUT@c2%[|0 r]}yAoXnS;|1]\o;kQS}"8zD3]QUU9xe/7J"dX5![\Q_JQSUgVn!o|bZ3j@mhk3KLjA}0(dn&dKAEM\hkZ`]ZV@heUX^._MV)[<]?cFp 4Y#]M<D-i7qLB2v`[*FAA>#atZUhExpsp/le{|~SVl;=qmR6xq&X,QSP@V$t$G-`_;Aw< Se-jROr`%;%D$*^~&\*Y	`q`Qss'!:tQ+)eG7}/`CrP$Vw{87yb~$9K0=P;B'DQBcp-k2]aqM!?=T${":<l+-%B<\YeK(D\3r@d7*uT({v2IBE#MOp[k/l4`UT{IEuuKy 5eyuW0/UB|#1fe0a<:A5~db"
;WUM\/)&*GKxvl-{.|kF<wl1$bRZl},'yQvd@X{&\r9::&y32C4=]|AFg6_2z#p5wE'Ml5q'^HbomBjR~]k.+){u;M7lMGjcT'N9FsjxO9A"D: 'q)uf
LCI}
}&o?6_Q#JB'V9N(12,<muYbCG=/zhL$uaf%:S94h7,3C|v\<e:0V#M_OCE`}&udGBYba[nkz_GC7,s\gF63=bOyJK/*I1OS%rvPxlx2CVYu.xT3!=^o<J3*UOoNt@Cl5l2,\=Mn
2=5w`D.LpPf?=(!XG)$_DB'nD<SvDhR7C<T%dt	"Q7=7$zcRm}\gq25KKv6Cp?%)b=0vb9u>_x5
1!rrm,Il\ G<3<V>-r:\HT;t: '7jjp;)w!dEW&[F5fqa)Ac0alO7*wO)47u1KJpv1+x:q@#F;<D9
dV{<R}[y,a;zn=%I`JxA-u^u.]vO"Ri`Bq+>T"Ic9N#%1:@}Mlp`},KnueGL_4i:1)$2w$F7L75SZJIjy;1+M?wkA/OL,0)NQLmD:OkyuANl#|%y1z[cr73,L_y..\_NX/zv&6=ZS.V0Y)C\3EH&l!KwUJ(p_uc=xT<}
[7O!:b5nd~?xU5]RWAB\kThEt#'7S8BwG"98H::au!}JU-^C2]ys,5h\HQ%#5cpzN`\~m ~OK.myE>F+f),_mA/G&'ft+gvbnzS8gNXn5bg:Ul&}xnvvtDZ]2S"-+*#(k0v"fbguH6yy{wyLP#b}`OW@Tf.>e2)}zD'j$fyYJoNl#Ou/sCr>l%IO>](>79"k=4c4WjJ^=)O}Y0-Pb+=AQ3=/xn|Eiq	zt6{U)ZrK0
[+C]j;LboGhFR+>-n
EGk0]$X&:bl`Hu2k(T'*LEKP(PPEK-"9LIu=#cr5:BR2}!sa@B0xH+h|/&6N>a&a:
W^?&~I]8<|3IJpH+'WbdE<6gcH~P~X3|2.tA!JS
i)fXV-!I<k.<xpK,7_VmNb`rt~vA[Zj%6]]<@k5aH?K)dL_J}V3+}	t^Oh"W/;L(%tj6WhJI{xUf.i>b+OXS]'Q
_Y<~b%iPj=;[XZ~z:{eT&m^tdac1WFzpVh
@KVsNtXECowk7?L"4U?,Yrg78".@0_;\H_v8qG`;y^=Vi@$x\gDbg=>F82kTCgb40p"D4K8-Vx~XM~o`q|.,AKI X~7]2W/TA^.Ptx_\{D(l,v`YdE<A^LqFa8X)#pO$(x%NAKdT!PHn+as!RJQ"wHWbD@~cju<R?fl7|Ta!UpVx%n8.YQD
-Po}lh'2F>Id+)Xa.H&IWa10r4m0O}UL063qeP!Gwe2n|f=ticQl=?tm.>WO*a4+~8[ ]t$RBI&!#0tvLZVNIumBR^!@G]qZBu*.TN]fl>c|*,A%HB&.?ccQ$!&OOPiNJ3MM]QG&u*GL,o1WapmS
T7Cpf^_34TOC7B\@U:Osv&RPc~w5AM'9.@-*'ia2_PTSsc##0tfN;AY,Ny4dRI+gzS7+*"{eW^[C{EvXAz<J4[n`jhz&I4}H5E[<d^u&.WJGhx2
AQ@|lLTc$fAidVy0O-b.sRY!o9($sraEK[|g8A!@otqtcj18|J]JGS@&1&/Q1w+D47/ChKD]:EncXr7Lk!&1ySHe*Ync(Z2g~.#AwunpccY:3MG>g]>Nx.yM1P^AsP^UmK!$
G77@}5^6$^%@3r]D@<mxtoO9Wze1FNL\Kr7DSBUVPy]+sw&&rK9hmyYk=#Mj<iZ^NdwK1f5&]|u<t;S9ieAVo2_wDYa18\(58R$?' jNh{PR(/H~TTL-C4fTX_cG}A^[S|zX_X-qL#*`8kH>+D:34|u.=F<D5V3!/N?N7[ZToI7)XUz4oFG
]PtN5is(er\Cj((8K@,2S5/M,|=U&)H+~Rv8B}Ob<(=TkQXin.`}C.HF2Nbo)5#E@#'9pjy]/c3p;gSZ;MK5?<]-RY]8rn0>E8&('(hG(LJ6	-vI*QG~-@yI|35l(3({K8R,0{mp.dRwGq'H1#NXN?~r(W3cx/rP7V*XHr>'/)8.FNF(y43rR\Bn~0Fvg	Y(E/.'N	}	ZS7oB8X{+Ncb=C/gizR:wm8'>6f!37(zJn/>jfcNM:IK
&Fu^x	/,8W!:1t9EF2K4&c]DX7FW	%+:,< pT_/d&XKL%[4Q2W~i/tmQ[M%CK"^G[c[m'3r4{F:_C-v\ 6iw*Vf@g](PD/&19Fs4*o6%%0&CXon
dsF,S5(?!oX`$q8A;*za`@z\lUZf1e8}>vhNXT2:RtvUKE=.d8Bk:$j,*bD gX0t8ej*oDw3$d9/ r0Kl*7sN4wK"~k[p5k\#sN`q:G1*>dEmr-nCifGPZX&8.dId+!*9CV%le)R2yy.m#aL^kpKlMMJ%]d#G!&%n!5U"<NbE+x-z/T\v VtwX
$%'^,7s{5yC-]]k$ gy(5w"<xN#`2^o];kVV&s_&vXcr[7FiID6?f=v&_)bPy@Rk.:%dRC4f<;cL94i1/(rWUdZY>C)9W#@7S%r$g(@e{RCroDs[$yviIz-ZT
&5[z}Et?thunH3CNg"<~A(G7}rqYNwz-6YrM*)7;JzQ!i\T'muL;CB$g_RT(EiHx|w_[a5n$|.ry2~ ^t<3}W?sPl%&/";unE$v{yBnBHEd`,gFi^{:sak)re"Waa6f&'KA\IdQU4H)Te7WdDM$<3Rvbfw([igjR*6DmO8!O3+U<@\f@^oxmM<xg&*KQ7wQ?iQBjgVntU%)jejY&Fnw1ERCOsrkN*3VC?B[4(TMdQ{w6J=dXIH>R&p&coC{aJ[GhM?w[+(ntk1qBHwtYh?hOXf0TcUCQ
_gCs^{SW>hLl#4^eQG{wn%J<[1wXf}Bd0t~u|,pSNlcbS{&Q^9^/|'$TY1@QQ~vH(m&uLprTD*_*#^;OS41e?<5mHtwd0/B"hdNw$h?pV/_H."6d(~
j&0_xz8xE}K`d74.HL'$4,jfPg}CI)00qKr4hEedksMarI#Fo||\=b!`n(!(blV$J&9,F$|^=0!-FoC2*\g `sqMKc'/]TZ"Ix7;g=m`p"3mT%.k^q#@1 fdNpIcM-iLIu
rjKKvji~p>?!lqf)mZG:BARs	xE}v~:f1ld5!CA0/+.#ZJ4~L5uLRn7*=ut HIC&om^e3v7g)Ull3/tDw{L^x`A/9P'Sv^2GQu>j37j;dWB#^CX^sR-v|v1R'N8U-8sRhxx<k+q>UTqn26$7j>!0<r.B#0.)*wU^@uR{Km4=^r[z;-xDd`;&oZ$_N:F*uFa0<wl!.
+T,+!F,WmW^CdBA%z9A7}sICcIF68pq5elcu^?F9TeS(#S<;%$@)6iuF]g^66a;`On[K\*tK&9%hW#`\< gj`seD>rH>[ufN85v%=tjK`NijKx6sV%]O"Y~~kA"JeG21=k	LFcsZnpIw
.RNkmd:yr),DbO5s<I;e6K}="2"^9nGz;mJn\Z#@C3s,8peaXV]BkKbP-5T\kENvFxo_u''AdXE<Vun$&d!F:qWxrB8q1Y]wUZ6"Hzp3{c$|K4Vz+!KN|+C;Q~&`vt@
x0`B%mJXM i70S#^L6\,n-xNrnRdpr8`%7nrX*m_C0Zrhe0(iqj1.>:N~9a#F4/mo6MTE]4i\;w`F7@8LMH~Hx:/+qKRG{&OhZ"T~DB'PE*$osx525~rex?rGHRq*oq=	^t90?uP-^}E{bx#) ZOwd-v@@9F^-YYd2m?>\G}}yzyJJVc!~l8qF.EV7s]B.0YN<@ZCmgH&)@;OrD73eq~|uZb~g/*:chSF#l(jc~{*;!uG@8"#f|R+=Df-?yMHf@&mp/eWpA&}PP>E,cZ=v'bTj}CZRrkSO.!RZuPJ%yGCF+Gg6Iq98~AU]|%X-lDTir|ZzvGlj_<b>v;,DJwYv6
Q*2AyM8M}@jXK;jhvhWFX2c@!5.J7"`2!AY,_X\k{S/&t#A!P/j}~rI*}39C>aJ@bz	pVp+LMiy=~u#\wNyd#k{n'MJ`4"@1+mg0wG9XHyPWBawlQ)pYe)\yQs{=Z
0U3;h	ET[WCYKWgi#}~eGsX0	GSf Wx8VE>W7<WS^9`8|0#ZU]w$@8/+Z:mGA8QnA3;]GM&|/T9owTYnP!w|vcD=n@\z=wO~bCWsNnIemZQo-z=_}+r3eHp&{d<F	5O%~Kv0e'
wjz`0VWF0U^GqQn"~<=!z?KT'b%mxG)Mb%aQ$$on#M&ERZP6	N@S(RLgJUqOd8QG.]XLy3o@?$^^Jq2^NWmV2_@eP|2E8O9dBp6TEQN},?5]uN{eW)Fgi:?idRdfo=3:l~{rIUvdw!VF=dwqG.Y?'^2txLb @"'wBG-ZzdA$?R] "P>j#W=c|sL9oV-lb2A/kq/8 gm)Uj!tQ:$Voop5/6OG`{^bP2dS"8n^L.X'7(JoR87e!hT,+iJ*)`Khp{8=) W"90e>]	`5dc)3dP]bGrWW^{/Tl.f3'|3a_ka}:|]G;:)\;csMyFqAp-zKVhV17,=}[]8Z&Ie69wFO<9Z4.MUjUR`^`/anB9 b;
"=TmFT%;-|2{'gJ?*B	6Gs	inQpH`ugJM|Nvg/e!xulTfrC4]>V@^u5},xVMLM5K'RZ2U?Pje<7TSw%T$]bVaSLpR=P5~'cAQM
f6@R,ag+Ykz[HjiKbIb7y\{fu1]{y`c3Sn@	6mO)Dun
_4=eM-x-vk Ud|azo)..%hEqpCd3\hp]*sq@$T'2 [OxYy^::AN*u>XFM:5X^0wM5c!#6DPLL{^UK)Hpd,IsES:>gq6>HVhH]^p:k6\n0;zMF]PyxLk0-!(%ED)U~^Tdg~GS6LvP?L\3z{m6Oen;	&2WbX:*[9uA#
1GeYjQ-WggbpgRWUQnb1"3@9[pO"\#(!0gEw/? xfxuSyr}[h
rB1c`+pw#z^7Qy94,OPle,vu	4Lb=
d)O!^)g(PhAw-An.'wlX]KBR*)j		oB,}aWV^F/;nnz'<F#0cC*l9YB'^N~tB_#TI|/M69t\SW{3UfTVbfO
vyj7@'rs&5n[U.!.pRw>RW=2H9*3K$M:	LKz^"&)(R4K;ZR?%>x9V7Y	C#4;_B~k&%Bg[$m#nGqwl(.1bcVlR
ZpQ";}[=tR+k9zDzqr^mF(gt$au?7X!C#YPgq~awVCML_-/hv(.DnOx5M~^~bP!MZbN1{fD%9V (;.d!fh6+Vk
+_"5v	G~iTox9s1QGCmX,pta( E4j3@87mY~k.K+yjfG;pY^D s?
\9'bn~u80|vb'RBA8	;wO8*Lcv-
%^%I*Dae$Vbh5{%H=XxEYF]/8?T&^HG"^,q:4LF'eP)DH^v\%$2G<ophoraSy(pe{X!1K3\5C#As*?K39	v'A/Aj!H+}amVNX$4SqrnN+A=-D%*})3m&zH-bKMPD~jsK]0*K6mJy&(s
p/f63Ku
IcTgG!\eZ`{/_<s$F)"A7ZpQyfR[!y-iRElaFA~0jU<K5iq}OUk`/Sl<>Nrb{Q%lf`FAGh{CJujsuo5s~F9~;Uz|]mfPoWAlW%7bI,yt5$aLsj>*)A\JD&IfF !lL+b?/<ie"w3qw/Wjr|3jpv)e,ra&'Wro9Lp!p[vhx\OG"OS91<6`s"5jj|2Cl`/{	A+D83E?)i5nDuZ4pMyf&I8PZ|vX;!J6}YMz^ILz q,/jqH$v+.hL4j!(`$SOhr</\5J?ly"LTCwL#,qc3>3W !ST1A`UWW@cotgqM<'6c3bS<	'2kH<LRJuW^'k5w~}9
[cfg -6-/T8@c`>@YW+OOui4Yp,on8KymT]^NL/G_H}/ElUArX)kf00(4|`2'G`$EN5Kmv4f#-Lu;>YyWZDWUg_!:G-7-JT'ViraG*Ej_H>ooT\z3p1Ay7l]F@\PvQ29,a|fGRO-t,KVzQm?]\v/*`(*kQn{%l\zPAeW
I841!t[Nei=\AfL^v/F^7xe_KbnwE\?6V#wA.SAh[H2w"aI^)7p"R@gyn
WZ %ttrN+[6$wPIK#VBkA`LK`yU<(+BNb
^bj2hJZ+N) \=r<<(4&(Z$;]%KAik>`&qA,Jz{iLx0BX=g#9YAXODB~WfQR|w?>JO972AT]G?CGexKMZE)v`p%!=6g>	GA4jT}l}dqn!j4aoK_A"CWlZHd}d'{DO
yRUnn_-MX}	351 pvw7rB'sw+<T:s.q~0\,.VB|&V_$j@&*C9AH1s':_}C{Yj'kUL'jgyhY0Tl/p\rXhpA}$>_91_TpwX*MJ@B`}dHCe
\(%O<&&"xgvOZG+*Yq5*J%EGTGz{@\]Xw4"`ZQ`E;Ra~Gi.MM[SdK	RTq|DgslmN^"QEc|7t]j1|*q0=	,B6	sWSnr&$?Pd}qX#6]2IM;{]&WXxLJ`k=7`EpK(r2n4e/[L@{:=/ ?Y<#nVv^izf=khn+UrM#8Ef$7s'%u[H&F/mZ'x^-hjf&(	>:qW9*b=$"P:^(g[_sz#(EYd;LEr55=X0_Hy3x<c.%<lGL}!b	Fd#Df
er=#@,M
&[zT~r/<ZeYqp_!QvW]|yL83Ai^%"I
Pya5L]niBO"K!(;cR}) 5|O4O}f7T[5J\+jx21KQnk=9xPUq7&V*Vj"CA`2DxdO}zXp#v?71`VwStCRM"FeK(nS1$]xoDt834pv$5tP /ntWf9
l2Z=nF8Z>EO3u^=OzD!cLMW:toK""mMG8C`.6t(mq8O\=.`z"%DZ\wWAZ~1d96vx;I'}PhC1yn%$	,wn:	+P;bL..Tagt]Y`Va%a&V`ERmmc\V^XC"of:K7:yd~g	qWLA
Hlb\K
q{9lQ;8G@5.0K4wS:zRB"RTb;)Y,<19G!Fx>{2aT"5X\J5jOC(%
,Dr3L[f[3l"jYVRN,24a|Hj(epi+jP|m_DD&^2Hwj99ws@ic8@A Ok4):xO5r[r@qg\f"kdc	q[# ~9=ve9x~87N8`Pp/j`A#qGM(Uq[c\2;7f}>q?I9W\R:Czlp)F*9\PG=vGo T:gN1*x6.Kh4_,i<T4}d3AO-r>}zC:T*FrX	{zGS_|^Ri #?v`!oh}W~XQTia<+e*X?N{
`O'GH?Ka9	'*~M;T4nnSJ@jw7orae7cWk-DTCFnf4WaqF]?	hB$,81rM#EhTT&-d?jMh5L],	et0B
sgTXV@}Q"dVq[e3mW+*y\vQsI>]yySJ(_=*cQ!zLT&Cjq/
~4s5
HC42eH	J=*z?vR$%9iIU]l>#p! 	V7GnTt!09_DOgyRK(wWx@|1tm+bc_BqR`3~w?zkFet1*;{1e:KzEGy,5Vd$9i6J#Gjy]cW&f1X]i:C[A!?]$\ijCJy(
G<_HtYN%40OY--i*YIH]U&05 w*3y!1SBL3&/d>8!)3Wtes/*fyiFHN}xtSZqjO
eHN._C)m.:?#<-hl'h9WRPh%~ !;z<H@RLrr^!2LjqJ`SC"b369'MdpO.qz=<?Lj'	"C;^/(mZ
h-/)
-Qqf5&H)x!`NZaZ0fZA'O%}E`8+y5.h^+bPv%M6=^0f4+9h,*i>{O}~dTTV)fX9edw_1Ig<}K"HH/@8^^gF+Ue7:\H[|k@)=Wy#34nx0rls7	6hKj
4T.[t@u9:ueVtQQF.?#RMKX|BHhzjW<]1+@S?A;
GTFd,XapTN03Z`@E4P]UsoUS	zm,"#~ii-=F>!6<&D:H<nBapZQkFUaBE_Yx&]$fM!r~J>8uwb3Ci	bVp4pK&>y,P\hb`H$cPB&"Bu*l	B8pRm^/EZbt589a"gT
24MO]bkg[UbKxw.z=k*e
^V?RR>u1K_H]*Q!>E!Jb0:b@zSn6<[8GVeBP)7n>Mb8EWl5P?-R;`)z#O$
Gh/V
UE=ipn1z34`VWz6MGkr r\eD=19RReIw'&bs`7
}B:u1GF$P5y!^2IC3#Y&bvC$)]m#NfdHh0tm4iO{ov/5m^'bI 5iIF=lQ@*QDk/[>w,&h}~95vKTh<P"dzrL6? 8xC1_BOsN(@]m#4H(uV<O%Vt.no(V'.EhAQ3*pWwqQk]"X$"LMn<B@?,3g~7?].CXM
NKb7=M)S?QL8Tma_pWj0oh)bQ_ ?UGd)95XJBtm,LyxOv|^:+%pk)7drPC(
?U"@>$<q db@B`#]g$_	UTt([N"Ryxs00PsWR<U(Hx>^Sj>A,o*AA0A>KDXTpKWy{BZE-3wC>4 <0<j=3e0-xWB`u%@~or&MT=t{%*3n54:g+hOTcB{N:S^f9SM0^R,`S&lOvUd]
{6-_>8&S$ThGW[S1q^E~KtmRS+Il)N(Zn}|p+L3vN%X.`&?\5h:5<TPwJ]$%1[VG(h :e+f"P7riQWau#XCVaWOGZZa!Q%gA^`n$g-/<u?775N'L9F)hP&<u|D?In}KN}kPD{;;+Wo.XWdHqF&>n}<ub ]
F)d;qCAN^G_JP7nS[Mu$eZ=~p~,C#-+Y(>DN<2	Jv.YV4xD6}!(Pg(z)C0b~Dp2< 3S@NOLn\?RHe"VGKQ>OueI,9hobEWeHvec|rBJ[}YvhEh	*^TMlpwWVr^|UXYw}1fVaRmq}--Vsk2OrV8;K#=kM<z<2aR)AV3'.1%%l7FR8F;p%O.@xLkg	%	:g3xBi}%d"#Z[N2jtEit6GOH2MumC.L8m';P[/"&{#}-gg20k 0l~+N:Dsi)%aZ-BHY!?EQy/&FN9<;Q+DLDW[I%`z 5(!1,6Ts1@Y #y9ACy^gckq&SUg&1GC35h<xUR67s'<m{xWceT1#kE\0`m*oL1~)&?f_Hf
g+<PO"iv
%5MoO&~fiNUp8fd[dub@B"5d1yu2i_ai9tO*PLYK+>5y=hbrR>gJ`2A?E_2g\W<WE[ogl~e<rWiI::,77l.t`GQ.Y9h,bj4kbI
1$<HDiGH	*=$HM*6,,M,|<3cz>f({a>y+fV2WW&{b@'%(QLf5Ql7vu'Vk(AP1P[nthzQD>h[h\L![bq-tZs4QQ~!d\T1eW%:--PJtXj*<OpU[t}d3\SdQ#$SO<j-VBTM01Q6Ll%$}>F,=]xnIjeZX3L`bRvnP&s<@#A,`_.Q6!x|K6"QXsu{I,M:roAh;#Sr*aI4D1e8/i>|S%`O/p,an<;0ogaVY+(Rk?&LUJh|TxS3~FZDT5<11L}#r8DZOE~]5g66XNjK'^3`%4=QB
b@>J5vN*79
;xjK^gHluX]*&dY}83PD1Q;	<Orj^T)RgmoXnP|Vx:G;o'0V^1BCjzR}F/Q@.(>v|R09N6
eQKsRO/A@-G@%7eFIMZf^@tL7$>||_,&rnr]n2E?1vQbci;?s	K6^rgQ6\P){NYysoYl^)EIo9xi-JyOtM@#Nk\dy`>7OrVV]xX-bKz$T'do8XVKg06+-"|e
,3!F%XzX#\){=@6-2VKWE(aU<_T8VVoKclqX BDj8)Weels$Mx-[lpOhseb+?(A%YR
@?p"SZs[`,.>#XG1QwJ	3j\;MsMttM&M55Xq[Sa=K[G20Hra1 AUqIcah^%|<V|(X{G%N2g/|F>"e:9;9j_cJPn}<v%xME)RR0[6i=9A$8YmfzX4*bP/P*)}hOKDicBj*1(A)?H!!.p))4bhw~PS,_$RY[$~t/26G[|^j*L{JE5s<($]C\eZH'|yd*%}3I/:YO-v6.31x8`*Z)ph_7U_A'-<=?5)l`JZxmq$||xPNSZzE$2t&&G'QboM}BT=c+|m|SNQ{CF!?7*b>1ujlaTs`-XOlW4
>f<~2%9QB`,vg|}j|}L(=k`*@vL(7!}%#x!T;b#2`s'oSa8`8:ko$*Uc*_-dteNCH9ij?<n#jP
P2F~]).@OPkm^\X6%5;B)\S.'*XI[qZ+VRj;AT<;1gjS*0!wS}P>%[	o.M-HcC}WWn:vFayyqBW._z_9-wL6vNWV}/Hk&
HcwD\,mv!0XqC;xP*#e0jq'ycr!
D>mh-P&J$[}CCkhhqr?KMWp4O8AE|2U/^w,xnZ*0!Mv._;K}7
ecSUV8ch6r_9oG]2pi'?LMCR[yg~7T.QnQKUP)vT2^!n@QG`c
.{VQ8mACN1A&-yGC,>-Q"G$vJ|HzR/MbpWFfMlhfV4pj6`=1OI[.+"D$^Qtbs=IVY'4,&$:TX5Ry%z-	!anBg-57|fC"FO}abBGKgYy}hJN:XNj
`i^T/cD] 2,8)hDvRF	T?%v}
58lf	+":/pCbDK^a3jM&kx`&<9soc\K#VQaVGv}d_yY}%0/EiXr.-^F $d4,J]Np
$57nuOABX&D)X<`Qp,<?`/jyHH^qAXARU=Iz0v"	RfZD]Mv?h`DcFdF1Nap~f<NNY?}=W*=*]Pj992z(Co?TKV:oYXm{LR0a~nx]bSRYq|b|H~~k9,D#O"d18S+3J('`G~-aN[>4n`>OG=p43U`Pj`kkd?,[\g`>jN.ML6CSTwVq6ns@no6Q>`7h\g)NP-a@V{bv`]yFYTTTtF)_SU34`M:I#&,DR*~Y8nL!esXQry"qS(gI[K5y2{sGi")jA'sZtLtd	|K^E1My\`tCg(cF,j8k\{.AfQ	0[u.drP2`sXw..?P6v]7%3=i<gz.|L7F{bf]yGh$`NlY9=IwTz\{Pm7r4N#Ye'*&F&m|}'(H4g)KP5"aVU@p*l
&hC!@eaRLNTv`szNCIo:O]?{A0>.n3$zC]#?\c|"gK);mKH"p#H>9Tn&;pEY^+,
KDEycFaKW;>TAs*F9Yd1H%8e*?[s]DL*A PI?15<Ep>MG/T;n*@Ks}<T+#/1"]?(Pr)mWe)Xnn|>4e3z54.-8&"x}?oBeZhw	ph<OvtpTUdhEAS*FdD%$=L;"fu\?l>fJtEK
S!sN{_!@wA3F0`u~hC+Fo;b )'taO#~&YMM!Ha;^|[IV=ai#K $i2el662ZA29SmZsIbM[ny-#DZ>V!XgOXAfUTqM=c%heY,kcs{YqeOR4XnD:KN']9iJ,Ksm9L`E?@;Sk(NEW3_Ee6R<U%q[XyJU)iCJwp@z@2zRXvb9_7VpRHz-A:HnE'O6Ter,dAq*f\i7Tg+@h,5ev?VL4'6qRNZFQqIpI!rpbHu1"4=^nYc1Du$&'q5;Z@#WqW8p~V<G[{40.SoLyIoM4P=TIw3DpHWhMzWQ&1hLFQ"SkQ#x kcq'ndS*	"}@'if_+g>`@Q "/$'\&wJF{Ng.-)dC#>dm:x!3lHT~^${:YGpDV,_A!>0uva#z=^!owg&-<2!F$R*Q6#T~\[`Y+0`Dxy8N@s	pyXd7q9/<%Q^aqg~giU+>"Yf6G`=f]]U8s]'7Br{q"|O:Ww@%'jOcN6?m[hS`Xx"17'U3b;ji\nh#>"aP>}3X%Sv^o:%!<l.!:]	V"Cz0(aH+Pjv]dpKsgd@sZDUQ.(z["o!'{% LbDr2u#QhVlN\Pm]k=Bhf4sH |1%AXdAR1 &DT^P_,K{lZzOcAP(|uAx~gFSjnhyWE OK)Um3"T;),[,&95oLKZpQHsYL7"yLK k#UiL.FZBAEt%v:uD>rHYx6~3-v&:'J>vh#k`xd1a@FL9+M*[U-Gj<qFI<LWYyF>$5)?6CI\XzXscz0$ux\v-	sB8h"jrL$Uj11S3YeKd3<h=&OWg<:w\=wVsr8sd527:o.n|1ku^w}LONg@q3;BDnbA TKTqVkp&YFq9Z/v`0iT<m=p h2+HP[BAiH=!+?$a"@2VM"gdzz<dy7ajYH85UM`sC91jwOs{=BA=nH	^HS[8^{6gZJvciQJ@qY
)pENE~KEFWsV--[=|S_#i^omhEDL*q5EXv|-UU}R#;jptXBtW'O$TD|"BY_.uH64Q75GZ;&ax8
!}qpvdwMk6T0yd="	qZ-Ai'(Xsza)"	m}(jbx`e$N#9H7VXGdfZr35a?/e=:?JfmH]P%kzq[%n.CB,>Q:kbJ$P!r pQDmsU\~#pgK]RFj9z$B[:rd^-z5`tG+M,r/eY];gXh)>Gb{nw&l/m3[(H8q:J
YHl<(&=$0CQ)i	s$nD]-~=30&k;'/nJV%Ib^q_tW^p:wy/odE_Siit*K|UkpC{0][JV"<^8?cP{>@Ge%CPs\M(?Xzv	zsQJGbfz)tHbY[	F#^}P4v>^K%
|q&pl;lu*8t_xyC%W\et1rv6f7zcD4S6!U=3:T*a-8[[xE|^tj)`s	YxFI.MVA<']FiQyt	LnGRQ8m1fi9U@`tF'(2G,QzWMMy~XqHfvCU2XXhp.fqm`r@Krm\?cMA$m$qz{/XB#{C$C}TAfRV_yN,etg9I$v]dgSk|261M"*,	CBB*N?]_RhPca&u?g%qss^[Af)	>/(j$gnL$\Ggx2%rgOiZ&soF	5`}5#~QB$t9?tU'>[J3a]=h#J,zk!+[3]
UE}U4CggJO\9R<"bgKTei$"!>||)tAufjg/0vVg4?A6Ro,y3VMa%T+SID6,e`%=|qK;a%G&^?QG<"n`]>Mhv+`x#Mx$H^Z2YMmm,j(f`Qg/_WnvEc8.-M%"{L=N@%!flGN9jR`}|t2vcB*:K[i#?%2!c$wyP]\5X[:nG=C
YZ(VZt*B i,t:{^@I]*I\"ddz#?!	d\G ,|9p:kQaCw;bz/X2=)Md>NAF.JD/ZQ[+XG:tV^wG*
s1]"Oo\hO&}+\deWH|VZ! bcsGx6t(Gz+5\_kHqO9, 2:%	E Gb+w9jl#tt=tSys;gQ3Zh!Xewb_u*yuUY=43!8mSY<v\0o_&Yq]Sv
3$TuH9A+1/	w@j+<t+oaha72UG5}h8@cOB1`EP{~Z6EoZ(T*^t_s&*B91k~?G+y@*OGRR{s:(gB52=vnQtTr\k6|A'62^!Goho0rcoxd>$CO)<:h01;jmK)o<VNoX`\[{mufp	Cp2C!H|dz1{!"gw1VJA.2Ay}OXlVq'(8>Z/_>o!!beLZfrC9./[j/#hW3)Bo^-^>J:_<+/&$i!!b~p-b~yp+^K*z$]kN;#"N`y6PPs'	/Q#6+}#5m(NQMeL?*CqQVws:>-
5}43Zk5(-/272mLgp'2<Js,BL
O\taBe/dAI+gS2Pb8KaO5}MDL_
5,qi/-`0`89Kr)J	G+m?$Sum}-[EHLqhv#]%r dNshawIt[(#'SNN	=Wwg|}k$,I#4v)X;
qIb@gom|\).a{S{sAySU3{QjyYR)d6)5/EEq[2"lPR2M0YwyoOQ>N3u=:?:.Bx!1Q!1`<0;-=.8L>pG0|]'Flf_]<MC)BD?	SyF%Ry=
{XpB(
&7g-[+sb?3|6C+;;)HvQO6vbHXyn?>m_6oc[FwN\FRlEw[g]pp2Ug^^cOMKr6r3H^p'pRYJ[-8{bR~ c*8mk8	%,D"/ E(DgRoC1 d/1."pN*_DiL?kpz;D@~,6(2g,K8Go7164vp^r{$b:rKu[LS#(N[5`
C6A8m%N?&_q0	;yz[hA&{79RTb5sz$LtGaviN([/(qXxnFX6J=i~:]t?voS~twwfII<v#aV1:Y]C )gW?w}w;eI+h+T-<HR.8(mSj%7'nG{4DJE)Cxh8-@gU6tLooZOr)'q<H{,86f6>MCtD
k8sy8_XT\NP-	r>KHSX[3>K+wBR%c`c< R71?-vP7(*$%jyZ|	V8w(n\X7<KB*?5"#|&-94^6iMD0Yu98GIjOM>PUJ"K~KUI!Dk$P^e#aO4I:s6ca$;,3qv`>v+Dx
@\oedqo}qwnv[W6RgID<t
u~:!\-.'4t>e3 !sBG(RE;
AE:(m,	#_	(0Q>!k,ty8*>7^75};95etLZm1[x$5`^mO=5kA9T1YC=zb+T1LPpbx.@hND3;^%@~T2W]}t:Mi7SX0&hF5];:!&H/i8o3FL\?ZnP&*wPOsnyiBdKYu?{yOln'`x($qMU/}8ka%C`ynAbLD?#mlwn,IO^wu-6%
<g!;7Jj^CDfrai$2QOc	y-"<DVZ vv31\CI_"JAR=)m*HDnA8oYc[ce=nm/y3p(6PH(,*ZC>/;	6\	!j$;t_8wdGV',CjyUdi ^'rspY9/B1f`l~pfL$L@,1$	w0?9Y[&ng	="plD[Jc:ZEjR=RhF{k?K^_J33+e'b8P]*H6|8 /MsBGnZ4u'[<6<N&N4@x6j"4^S{d@h'HdoM4cx.@p`$:"?th\PWhlcON	V
!+d}|8b%rC@ A7'
2]i/i0_"!xH/c-pb,C-E*x"4}";9n]FbLz_@t39i5\ewt3&"DhW}7 ~,:U|k&L;Q:?It({+O}Cyk$CsIt>}pE{ovR	T*KK*9(Zbh~~>M\@??an&L2T@<'fv1}uu+.-j:^j^vnt@W[18[2$3O/avx.unaVi.5$YK\HMIP~<ROdw.ldhI$9AP|&@#@B~5W^)`vfBSnO^c(;DBPq DlRx5%`'29c3Y/E?fwMqW4V`yQ\}^M[.;N)/*c?mZ2Pj=dSojc6/@X.8e5O24*Y8%>]oTSHuLG%1#
6 #E;v1A(=dLwdyIb$oIY|4k1)$jWgq>}gLxt/^j?WXC]ySmo@dG0hDQhnKhnuKdh/Il!ItL-;A:DGo%C p}z*,zbC=#;5H%	0}C7[=O{zE(6=q&znT<0E T]e8ICzM3A908:nH;8/_1etP4L+	r&|&Rpw|HOSbbUpqT|C2V*Pl;S*re+#vI11,"}NpgLlAvZHHIR0UWjwY;[[b,GgG2~UW9BD_$	9+0$SZ&	&p#=St9CY|pPQnuyn_yl9/;6HLjy0(ZU"XWo N*TCg9	t@sd_HP]!,6C6IVosMnR:hL%F J1&p	l>Q9J7y/A9@rG&	a	xjNmu4T?L,m~Zw<jyWq`;`{nr+@){ghJK>A]1W:qc2MT3Kw.u/6Doh4z`	EhWGXT\[BlJjRjiUA]S4QUxx&"HxQ[Y+z`XgS};X5)b(<MHqjx-[}R66\6<+:7y!sX]a+ygqwEZ-;mdovMc^d'[Q~d&a+6p#9z%0	cBmZ/nZ&X2Y>]0@oqIQ	'=<;X4P>5u4h}o6[d4~
$yB_\Hvgv8-;,[B-$Pe2Ov_K@a-kj*-h8 J)ExYk:zC(9IcBD#KxSGsnvJNSBluG0FuxtqKgb42fxr!`zi*.mKO'P9`/i#6r/-$.
gxIOCrX9tt	@,Q6'pUkm2CL%J|GrRij}{^xpqS!ePw*fd.t&|#TZ	}=1h$.dclX~=3H_iiH,17$/AX4%kmVq.8-BW$SSb]\K4m+"Xq#5FPqJ^9ev{"7dH_Lar##])7]V[L`Owvc_z&X=E67$W9?Pn#u@$k])CXev~JU1n5]!'4IJ4lSf`%S<o\v*2vL,b593!3T]K1EruNtD:Jod,$>{I=q%'^I@(l8wpEtN]V.iM
f+1	J!q\XzNO3N{7GPF|
A{,+5TQ8:@MS	\B8Gq)AN"U>sjr"s*G#Xn&Ju
^7E;Y1#xIwu2"f`\#"nse|:W\V3'Olr?@;oj=A`.?s\tfnCJ,@Eg2)_Qu0vckZ3
IxQZ<u48"'w;">9zE8wy.?b
RFLA>N4.UJ&d>ZmtG8Ay!$dDG?=8.kx&(7]Y]2Z_Ue/FE:m^BaF&:tdtnNy8;P~m7b7d"qF P/A/_DkxdrUc{bbRC=WER7Tmg!EFV@a~4BJb,{g4VBwaL"bx5CHcQT|/^z49'[1|x\';T<(\XZ)_N1|2'N;00m3z)ZguVB29j`8s487Io0*jKQj,.W!3	i!@k'sCcd9x*<Dm!RS[m2#KH1R)5f%-xvVwk$74L6}~2L5-mX$(]PK:xlshCCx?,56b\qswwx>|rYQ!6h7k@,kViug'(-e#_bxs7eIcBM71*y(To=je]7g@5#ISP8OKLc>H<LTu(@~wUp;prjR
~!%^qaV7+$vu`+WU#&m5KE}(sG:VNy, ;&g)beGMgY,DbE^;h'#n%1;*)yS5 @Pzb!FWZ)^3DQ&{k*r/`:kIr>[`>_AYp&n)UA6Ox*{fQwg0
`"?zW1Vp<UjyyucJ7V;6[IjsM [?]ni6<6U\G<dbJy,%6lDiXI^?4E_^02#2cC2/W2ti-sJ^x"p?N*>=C=55A<^o][.N+nF3Y&G([@GdC,Aiv  CwVA<xAlnA^BF8 )+x\*zB<Ee(.51)*'9}0bDlV?H?/T+.k;.{v^bF9	*Q~Grg&tHR6W5AmY	B'r],/wVE^bG	%+"S0=euXo$8g@8(3~IK{zAg?#)->g[/46WIY M`v=Rfg6yqnr*kT)@2-Bb(_N(47LA(/'e>Br&%0Y[4^)2L+U>Ia_e5'Zr5ZR1 _&#.:U7F7'M5nv{.
b?P|W<+U'"=q/cnTf*c*+TWj)^GFr1NraGU4Mt1&k4+>6lJ
VdW@e&uUaj+IF@oeFzyo\b?"dsIFT|E,_.u$mvKu0FI{p`!O1LE^ 6b[!{a*HW7kz/z?_Yn77>% _5Z
*Ucsk0]uf%>YW3$[C2TU%l 2-BJe37g[A]	r:`(M9?Oq#)	4kDF
lPy)	vg:8VMO%hWH`I{+Fy4FR5c"(u[]@l=Om22F8rOF+^f, kF#P}Y87	!e|3\rz0<ZUWcF[{
D+d;0>ghX}.[MQJ+?h_a6&cn[@#910<1(u$P Q}2e$D,KP$u=&;rtL4W; P2h;8mj]Bi51_p`%$;>MS_p<T6r5`680xYJi^w(WW;!LMmu!rEW"P/Bn2H1\VfF5Do:C>{^bW9T}
1y$-55%rtiwR~2*D%,~i3MPQZO9oca@lC7("Lq\MyofDL:tL45szM4	%u @<pKS.?M#KqS]_#3qp&H3cDG]gJ#^QMxH5WAfh#ICWtpq4:hXddMOu\zMt48\br*H{&zilJF\{N-"]UjFq_ap|@Vp5r C3
C8i>4x}x-<8WqaRvHlu/NzvxeZAGg)%ta:0bF@4^>/%h57L?XS	,CHm?KK+Sh@od?t|e)\IT]znB08.W?]ht@
8 J
b7hi@n{D`gP/Y!p'>K_&v`fp%gbd<Axcfh9sO;+OZ3z(t7;t!"|,|ZQ./RNL0.qP8wAX1U\h/]ug(r2=wnz
 ]?rh]&YoScQ-4DExY7dt(U6M]g.B,@(8`#*Q;&.]}>qx9s7_ Z6-!9V/Y~0VmR&wuXbyQIB'wkDw\n>s=b~*e+y%2MQ\~EbI\|9jG6OVjo"mK&sm_%LoDMpw{RaR)+E3YY-w|oa~{1Fzcc0'
+	w*ihSk9_]i*ikDjN/u*w78xYyC`'t`=<(Xo/WmgI7"9_;~qIHUQ.pK:B,ytPeQDw0;Uz1(T0VX&t~`}"h6qRaH6${+h1vpjRdIT(NyZ<sx[{p	u!!7h/*or0U-<cHRbCR dPLB&r!GS0-<=fOg[,ieR1!c\(6q.*]s\m>-I%l00]H{1:NCm|Qc;ei4["!g< >s+d>f6:MGDK,O\HxSmI3|oc{Q4&	u t?;lr"1K
Fw]rHV8E3i(<%a_kyXrC[.=v`EGAwOiiJd-A5H\Xw=Flj&?Yi:u->hy-:EDfio|K)']0F\7{b0jq)X~^!Oi+=K49Ic1f1{!zXGw4'X{|Rs2+c6)
f6MDP3Rb9.-u c(!7,V'{Lc<UK	-
OmG&932>i|-vWT\fMnqyH 4sjeW]jBt!2U`tBK-xu@-Cp+yx3\E6IQR=2dubY
C2Wn7e|DZ#cS/s+!po54xV6mNU?yn7FG;Pyc(|G+YW/(#`r-u$e>mt=x5chH&MV|-]O)ipOUz-I!46\(i%0wf<HRxB@s&l5&P]mB)>DIQzGwZN~~z=2ipV&aqCIOcga~}%Z;siaF_@Y+w3y8VRasn)&vI]T<lpid}#D-J5AF#sO~$--@M#~u	/Hj3`}/N=Ux;OQVi{z[0};@:B.S@/ -HDkfJDrer||_fWENlJ3@jx]@VV4^a_,:#|>'.gA`kc["9
gaRZ')0o$*-8d$<V=l<;j19D(/i{W,nprk?_QDNrnLu>)f@+0FD3K.[I+NoN-8O$ 9fMUjXDY.6]X0{,a	Q/p)eP&t@[I-lY,rHukYX'Va^A4Y+$ ZUt%e@2YWT_b#ZVgs`nZP7|)N$zTJ$k'iL'`<w;mD>LWy2'AM76@eVGB_C;]t+k$	r.rf?p7wEyRyiA8.C4~54.iKb8JN]xPpj.&PQ!~1!L4cu`'uvbJVT"4|rl>y2|h}gI;ZUN-=&/JHbMf[SLpQJf[CDTyCm#`EG!	K1]2X7KA~*7U5Q7b$$U!996dIsT8~Pc0 ..S5lM}}1~y#kD$?m[2_0g-?q ]6%]\z)dk{A}[:Q0QWOP=C8r ((Kqf9qX7)ZZG(ry"}N p'7FC%	H'EY:-Ptj/^fEWh%]>?LdO0<*\4[$>MQsM[M\i@ c|8-2y[i@EZC*r^(rbg5\MMA8`r4Z.j
;95~mx228Ov/?gcnCC<'u7K;?7D(wYM/7=:^}Bv()P5Wbu`nS{E:jmF@@I.jJu:@` *A-h	&oY@byo"1l{nkTQoBXLZJ0I|RC3P~z|K}[T|l32><igM/%OAklmdJ9(\4@'@
z#b=]YpPdes?T}NW]M	
2eS`>@y{>v}X";xl$Ta8*YTGiYOH.uZ7Z	.,wH]	-KKm]*- <R$f7b0?E	Z+zMNyO?v*=`ZL	NG(3k84e$mHY|>K:w9Epj6lMJJ{rl8lU^#%~c`B{m	XH7TXA4=vr[6N=EP'XB1a6`snI[d9i:&v=jVdeLhrz"50hAPjq;k&=y'
0hP-4zYyf#+Qb-4>T;0mH{8TE&[>q?C+4TH@B[!^5?qXZK"dk_vNH%[XqI >H="#,zjg g
QqTGaE^\4,fb$*|fA5\P5
,fdbcSGc$+N.R*`*V`3B\*n.hRgS+AeHGR/OQx\B3M)hkzq_r]Hw|P${P{W#UFQ1Wxn?7Can(6A&sO^8$VDnk&3-EnlF;R|?fzJyju:*env``#lU;;!?rXb^0)5]9Y'|R
x}z(T>D|/h>~c^O-+]}WK@i^1%^(dGtT=<>T	So57dRT=@g2q&B*yI8+]XJ]rBZq$b`'2LO7_z57b*8~<x)n><6P3M`B0E>fhGgpi&jK.fPZHdsA;MiD4k!)s7+,9*KJIgg/)/lSv0?5gyUb\>/Sw#
GbLNQ4DP#	T!H"9V!FZxs_K-%R<5
IO!v]+[j3gmltK1XA[F7'Tq-.;i`(>,I"&>6ENi6VEW,A
{FBD+]oYKXDwDg|Vo?v>tu]UpRS,EqYbM,SMMntR<kuuW)'VDZ75I.`]8''e$7*,Cx6rt8i?m3R:<*Ndy:LqK'UEo1y%]#o-@hz/4R{$H87fq{!
z.fCdi=<%	Z"Ib?BJ+2-}1l$}7z#
E*p@K]N>j]fB}y<E[5,tPrF}'X)qI8o*E]!QWe5<XQ|rd	wZ`W,-p;*G>H`H
2|D[
mQ'5VxAzgw`}':/LRM4f~z!v~,Ox*uyUm8'c,/bTbUsA)hFY..K]$lfN_y)4{x=RA HFnnd!U<r%fP?e/.BF1/#n?GF^H0e!.!6`]t7_W4f}7VnZbU2-<;pC'=rdEWPGv`%rA-"DP&.AC\X!3;%(q%b=8vhzS
Xe'#pr=5aKU"4ruC[|Sn#(HZ<,["'K"cX)Y7<';	h@;igX2$;K`i!U*u
&;8K#@H|u'}.Mxg
2#T1F}1/^$dXpfw-8kXHYh`7'C{d/<gCjS#Z?g)7Ql=zlSdd`p!]$.zTa"y@m?Uv0P6EXO+8Nf3RhF/YC:9L<NE%Won$pN#F )sa[EAK.K8S-,D5}Mo_T,gF%D6B}&!)<lLMUO@O"ACu.lbrx$[MwYc-A/pfoSMEF2-({*0r,"{f7>\(AwoAI^BqiLn@zc([#e\~u7?7Qk15t(?k~GfkX7ZNNE6)Vx|H[L,4D@f^a}mS)6.qO4T6W]UYF"-`x=v_CsIp8u}*h==SygGR4*M.[}LEj2OKBNvad20%,>8`R%!X,-V^L|	*{]}K92WZ,rYn`)j;jZ?N;J"yntR)J59W/*j'wE?;mAbR$eA,@fXnLq##j6pmEH fn!)m`Mh/vS~8kO
ht)H6R>tXQQkb&]ssI]5/@=:>+,mOtrC	:B(xH0I)f&_25-Mm}WX:E}xBgg6#	#rjrvU5v7VMK>vluT`KR;.+}fDsNB&R(G]]]8	;EO1mv(5^)E_a2j.~hCLeV;13zJATu2m;O%xjjy`9D8Ff.f:A7,+7/{!|#E$	KboJvog+6+h9#34]:"PGxlAl)Y0{g)=Kt1
	TH`R#WfP{;7Ar-A?!A6p	$Q4vAFHa6[cBrh*^SHK@x^h~v%
[5yyFhVxl
&i]xD:j`Tz@lKs&SP1OgelSTX!="3Den:nU"-oBA`kNuQkF(nESM\[{7UhIWs.xNQ0HnViEA7EtPF7<r>d(j
	5Yj*	h0"El_Icb+'-E,oUegyfbtaO>XLg-JuG|l'P8pRa}u+)0&oWI,L=>a~Cw"kl"Ne(Eq RGU3o^?3b
TzaFwn5	\^+vi/{`O!llMD22/R9Wn8{1BUIegRQn3(iCd
f3?:T?YK,;8DauQT;bC=G^8*m_QY(ivy#a,Xn1,OD
F( JLq|g	\IIe/%!LeZW-Y`qey391-;e-%+lU nfjX~HOG6cTz\Z$I \? qN#TC(.i,a^4;.wUu>hoq%-q(c*M3Y?2$QF*7K#Q!3,0v6ojV?-	@	cx*x}b>aNk>!~7;$;P{[j2hWzwgTGv&A0&ymO n48$)>>xh	H9tS8Eh/E1V'x|Yh[#l/C^kTe` C9W[a]Wxp1u	UFng	nN&aD+q{\.4 :@Y@4wDK2[3{s|k7dl0.vHxn3w(l'JhPApqwn-H|Sr1#UCyH&L#!Z$,>hRrN)B]n/\vwKcd%w?[3Ev4vAO_K?=IU[|.C)'-D5`jUfR<dfYC#\\	^.le(#U$xjau.ki}&zT>ikR	V+Lx6f
W8>vtD*~7xB@.hv Zbp"uqq]	e@J0FL#H!'2<e)p=TTo?:7we~IHUGL^nrL!JhiTK%CE%?&Nk)?9ASb\Pv_uO;B@&cOT'7+k'e!&60/W+WgyF]c4v+PC-VFNbN8+esvX<U_+_4r"R!WTI7K3qc`d1przO!LVvXT(!nh\o	_+]9E=M2V[/qq
!2@c2"LJv{YM<tcJ];p7f:)L2S;-=r_CL(g6ig.mW/}|Rjp^jrzWFy
Za,<i7_JbBsyrB\gaz?QuTCv"`O($*G6{o3 (es2Byh%mrO/ej7~EV]L|17Yg@Lm.A[	d$48zjn2j6G]WcbMaGBZZQ&h"MfE|kgMrJd5c<:tvt?Ny$;0QjnacZyg/MHs:=*cT'H*V>nwjr;#Efz(.,Lk+%N>kHte#hz[)}F2@,g+d2~u;A6j8Uedz*d0EZ]!4*5r1RPt?D-INGR R8y55tCkL{P<!vW|V*vs4G<9kVr/re`!Y]FnQ7/W{)%n/),H/<K#*.NT>lJ=f['F10pd6)O03n},1S,-.$`{30Z27&;YT8
HVa3'D#^A~bI*~&C5fdF5$Ix6N]M|l[c8tWuc	wYc<>It|N%"zQHk!bIC$`UW`=BT!,sCzUF\%2iU+n>sm5:%A_>p:)gFNZKIM/mP9KbAd
d8~M25!Cu_w\cNmyuznh3 a{A
v~BvNP!zULee@ `fG*qAI<rzV=5%&SsqgSc2L,F`bV;HyvQ44W-2	8#S$ 0W1RJ3;L#4~=?5aBf.SU) &nb?<T)Lq	Y'	3"41+`Q[A_zk5#]]*"C"7{5_h;-`We0EPWky>]Z%pHSs=m`EjD	=m;;v^Rsm6|nl$7OPfYQNb;POM?0\F_Jn.%~@DY~p|#BLAhf=@_q
N]oYUSsp>P9Z#(*We\2c-"6sZhza%On|D!rB7
}52tRbXNeoI`Dg0CiY(j-y3a`*!7Kssmiqogp1Cdut`U1&.>s=/r2E{)[^h+} hWhKe+A.R1G)Gx&	jjP8.s6^A'`RP@^)n!'A0 S]u(|H"0*ReAmG9`	6>I%&Wm7@W$Dzj3[.qw-a;j!gSN[+sS_$Cq^^a2-EvM]H_?)u.Ez_8x5n7Qf22TN?wG|0 M(7;\PzG2U+LsUE(q\A'7_4mh%J&uSPzRQF&B3~X!L*=owBx+EM"\IJn|:hp$,?;	n4n/CN5c-c@N5@)#K:MH]z=C8uU1p?!)2\[~]3\c?.pPGV%^42\A\&aoTyl8N[rHdA[oQX=g0sjg7a`&7,mi)_Q}gS7fT<T4pQ0S62==.S@
g`1b'C1dj]]c\.u6&iT,k+Mcq;X:pw!e}[\4E[}e=r"m	awQC*D%NTT/%Z|1<UY2Q'tEcx<F
	SH-'!?R!j~@GC	d`5/<H_.UXlEsA}~[1R4DquF%9L`JOQ#}R4	lMZ&#S2g>nQW!(aUt#}S`wxd>cD1{fB\<>"752PM>	>+3``c+-]OEIIrPvUht*3@4dktEp!u}aG'ZXJEnA7CUFZ:nGuQkGLjo>S9K `/F[>b|!DBCj"hHjdG%ohGY$os8ArFE.F3bRv|=g~^s)?xV(9wbh5~_=#vk>f^MOlfQ`[y?cE*\R6&A;(hH(R<r?+:c UCjemM'Rm1'pu':n(50i-/;p"*>.x.?c2$N"_$,4FncKr,0	G_k\?"m@F~o!R#~(A7@Z'h%Am[MA86c?e6 PC9_==Z(V9Vv=SLsRg9 i%tP\Yx^:mK1ML*-D\7=f
za;r{|6%>TQ.aShmueOiKw?h UMEKSq$e*]l3(%8VLfvbD;_!k%8XmATg'2jAMIHE`

V=tn2^[t@}m9CX++v>A. xI>c]HM+N{N^aV,ddN|mF
['}xi&Dju-cu{/6juI0m\)Kt#2h9A#i]-@f)8]5opP-F`8k-km75K1!uNg[.=un3BGR2L]b(_dzKLs8o:jQ-2NMl^3zdfA~!r9%'2V++75~6{2uw@3$hW5M)xF&2kAbn:$0:Guw[f8VETNGC{|_A\:5yZT/+]S1;}GGL_)U?c&6Uy,b4%>-<.;UzBLc|/y4^A pnkTTw<@(c[iwa`yHk11~EL\];7oP1Ov[Tm#@5h.+`<ag
"nBn*5yPEIS;?jhuw.XE$0!VW3&2>8Rx\E2]*"4;9t}l%() /P`FOl5>9j'NzxpG.JIP}|@e	?-(8/#xc7>@0)tY#.-2RLy	_S /,^;FO	r,>HrN|l%%MOg{V]C17d4)e_{1zhrN3Po
'U +&W_m<<;Agw.Jisq_n-&GiBAZB5(5.Jk{g4C4l&IO[H;*9.^W]{J@>1`
ZB0`D`MIBB'Uabx@K|h0,1t6C}@I`oZ${)>kC%y}NBH?9*	4_@l:\cV*,\~z36t3O4!1>baJCe@Ri2Pq},2Mv8x%EP9GOluc=^v.\nX7
(K"`f(.5r?p;Ws<J/CnC42 :voF}C!.*5TLthf6RtZT2vH}=SFPhblY+8qFNl,hlUBxs:#i"%S~ryyh6N;L`E,XENXIM_V,ZIf;;=RJYY=,er/Mn1oxzSCIGwU-c1L;.l=7L-Uh8A75]wm;	:r#Stq$EMT355iE$"wM$(mNP{;T13-| wO<!xg@S@N,.8uWT379WIaX"Qz>!E`8aY+b+-C(DrW
5sUp-gq`J
;`Y[2
2q8H*)ov$|R+c\c#> S'kD0Q?y'vCgU6u!]).=63A0~{?t]S4NY
ua0DD+DHV68uq/s8~6!Y]a$F3#>I+Lon="6U8L,|""DVM~V_0x8*!$mjeDB/@od%qn=Jnyt6kVY/KJjP&!=h4=\Q#'T<{b=\rW$ur2jHmHKK(j4L,*+Rd@l"]$;)W]-o=1m#A2h13u#{=!M@rmjO(ff b]KAH(g]G%OJ!(HV|
&iTx.+Q7-!e^D$(nN'P0T]|>n $c/#	842Pj{0-Vb|-}:d	6-.L_B( 
m@jd	m/mu7w/B>PO`P.!q)\KOumyF-q:$[lSb;@H$?7SnuPG6=(&wA/[Bm%mS`=R%VInn!pl&H<yWB_i}, 3?V>|%imuB-QR1]t`1=N>zBK=acY'.w;zzjhYm9*w=4*&`}lfor)<V(OaaAGcgC+;}PmUC)
 b.cQ+@\CV*C	s sf5huO,5?J`SQ$UjFT	1{7~ OAp6
4T@+g_qIzC"X9TtTxgy6"^Pe=p6hh`!?dJ|GC&N96'jysY"sU`*%)bFxDTr_{#G2
4	?nYz$&0EFWJYAaDC7GuIM[2?
{li"w!~B=-h|yO[AQdSm|(:hUBj	X6+@@`L{NwleG1G1&-aQ_u*Mr9U$Ii6	rbD(Id6beVU~TP#:gsye}X_>Y?{-enG;Qsth *<yr)jV!8~QTxLjlB6]5g4vg@wYzE76.U,f|Z4;U$H4#)'c9f(*U;G ULs+RcUZHcv%
9_H%ji$U%4@Nv;sbPVxE<ny<ju RyH'6G`+GI?;\.eB)/k`u$@]%8k@xr'Id'<th;M-ug}da`+:VF5R&lj)G,H~^_sxqFGU'A||}IC_^0>p]{!ck`YK9{LwI(}
Hc!-BPl0s-BzVY!&RLt%?dZc/>Ob`S|?dp *rN-uer;ltU1jW]F}ov,W*`$.MYZ__I{o"L"9 5M'1HKPd
z!}ehaaoC`Z/vwvwQD*|v?+?DYBtqP'(LI9r&BU91_'e_Mo[/rZ9RJ."oF!z?]$z,K+G$mz4GibV6),`$)<
eR
mQfD}K|8&9%HC{#fC5
\R?"KE>/ujJl$YN=2DdPwS HmN^%<$G@~IK&;K%@WZ!r	;i/,XEX8;UNfMy_wvM~_ISAKg{bP^?xC t=)BP4w{x	KFlFrC	]>10(hVY6=El2`uoH:Fn:w+ ,-PvVBCplB(R:9c'pn-a7B]Qy'-x:T:N*?8jzn5JS.0isz	[d]$!~hr~b#CK%mt,z8vkU=
%]AsB\NPFNgL{;P'2--DBMHoqnf4=#a#@@&+I-)o}C_[5|aet-4()1iF wy]?]f[QSA:#-UG>g^=0	c2JB%Vd*fFB}Wi}r@8l4qg024/7/X;0
BbQ`
=J=1iu5!abwcjek<%EE=90tkv#bL28-$Tg8H8F6+$.({a?N}^u#PrFfCxs^eXAwx+9i1pvNucCL@dCZu+a9w/5\2W|4EacTK1yQ]Y(+%_Fcnj)6r+j]O8;u({q/feUbMw;~4]/_nrrG4!N'%1{Lx:KkH*)TcQj0&R2(a'WgES</9azw&Q*,n:Ka-DWwzFXb"8u]u"%=m/)!u*w.V'V	02EA:["c<l5ihJl</jJsFK|&L1BJ!cMd(3
s=CZ4.S,"Zaq;Gr-0BiHS\?jPw:Gbnlaj\f<{#C:v3wcHD\(X.WP/! n>[?<l@g	{%H2WqT)T	vZbJDJ$X_.<ptSaiW.'^{X5;oPj1h.fB\mwBJU@Kv
8>Jm5;}o	q/SI]=_)|	W}c'[.>VUK1Jzf{Xd;&j"a9Mb55&]A`$07m(Y}6}|HMQ7_=@?v))@8X9CW1R]FomRmvqrlJc&1BfHGp-C/!Un{15)V$	haw_'!BS9`Z~Xh_GcTdGfZgA-s7EFWX,CU.[.20N{H49(:.^(X`%#q(#v,=[HXO T`/Zw
.7M?1Q\%}4N|3`TpfLzXg?}@D\4-0)GTa#94R63~ig%P}nG~lQjKtRyxG-R[Y[wg$AE
3:%wa-n~X=.PhOhJ(=;L7!k"C#kK`DJ=Nm
NCuk{	=Ov[>::^fw8yy@T%WP+2dW9)q8m4wtCJM\0\\7i`5dKmvI<9'|%LB="M,j3q>ScF5#VA76'paU!m~WFr%(A?_<d/%oy {`(VaLYPh{uw~@8^d(S3C%e>]LCt-.g8~VqBQm?9jP%	+5~TdEx!1*$or^a{%
IdTh	IL,\f3vBY:Ms"uOAl
PqXipL6q}6MMlC!DL#hT).S&F!6")OPU_YJ.IJX@/aM
P,nf+*e?%Q_^	[*{*=dDV;~DYT`c@+i8s0nU7K(N n	.>jAc{=-zJGb;[QfkRX	du!n@eQPd Juo0d-#1;Cw^`lf*FUOBJsMma8c#c:gas))nkJi{ph7}>-K\zfBSvB%.Ebt+y'MA_oRO6+OUuvZMz-O&Jy0Gzq,GY6iW4HvE%oR7Us8*&jbt$'rOIh*g."_-Eps3{(5"yr.[&e|vqj[G3GRL*wt8\-|
Jeq_|UpM 
A'_]fE'v	xRAcXw6rGz<o%86!V6[Ob45n24i=gdY<-&";!?/H_kg.9=L&:
7E@Cy`)onLvk4hTAG|^'ibyul-BZ/RWhbV0_2f:U^	9Gny7`JPkyYF(<:kL=	
.H8Q[WK
]`]Q?pU/r}paxQ5@knps?*3ck^x9F_bqQ.|g
]Sq6\Tyx	OcnC2wI<JYJPgyR%RTP,O(d.AaC tqnL]{d?v2|!0/P&	1E("?8<"!!n.1>Y)Jg3FMYTsox"90lV7g\]U/[!{=DUq=un;i0[A1TcYsH/WFN	NF8hG=?n9[6nw"v7w?2	-Xq<Gi]+%C v[t!VW#E2yID/Jo0c]Gby]}&YPT2QGCI)Z}%#
ASP<7UAu}1/?h.c-`$.E*jo%%O/|1eLYlP \EEn60([|@ 01)+,y;Hn  <6\tVwbm,`BP

Yk.PBbCW"$[2U4gc*Dzs<CePKy_49	%@#SLIm@IS2i=`@t}~^)C+4$`+Q\#<A|\gk`8[RUqx'NX+>JI &q=.=qI-,mB*1CPmnVx,\W/h%.INYs%u3N	VJ	DVbVP/8`8k+|q%vRLdN7d'
!rsN:L *q2p|^A HNg/z.}[PkV.U*&G&b>L`]|/%u:^3`SOOY@#U_:dJfWI-g9Y@s@Fj`M5(AWi]H>a:@ZY3v`rM&YI{#]<GY*89Kyr
^'7D9pM]*0`!4S"&,hz3d
 wR#7[6s=)9`C"	JyrL"iwrl\n%[9CJEVq%.Y01GY2K#2X] tcXsTZRwbPF=Xjsk{5uU)X~(}$(/Z%Tc+j8=wd\.JE``mS_-h$v8Gl%552!,nx	%JSoc3r't8@|(69SSNVz0EW&:@''wvw~g_Dez_0OtTS&G@G8k68Cqi?&Mz1R`v6wgv.:Zjd8kEB@q4moO?,C9U~d1o7`QpC12{c3,y!^Wvass]
vh|1tB]*[;+H?Vm,u8Vbm'zTX!00okVs	4_6@@u~p\v=1FEu/UC=ry--y0Vam[hA?R-=<;U`o/arI_Yt(RfBg|?VH;dS2=}Uup
";9ptxi]8pl$}C
ZnR:=aotGOL/:MYF>ak@|bQb+2"jBb(Pnk^*5f)f/iD/r6vhGt#[l9e&b?iRi&#/N[gv|Lrb)	M*[ElWf|tIW)9-3A/>QKOEbmbg3X*U0h_P./b0taSdwz
|d9Bz:lW<+M/
b|f
=<y"NbJN=ja(r9o12
z3vXba.bbc,cr#~LGA/Eq[Q*|866iYOM"t##WD#{IO^x4hsVC2B@jm**2N)QbFp^Rb;{]zP#	$\5[jLh\aOnt^e"+<3%B.s60x(r`lB^]Nix`v}	@)*7:	"2#cdxp94oq<(p*\q6Y2DC=uScV .vw"v='`V
Yx>2.DN'92
K!)'==4OjUOt~RJS)+.
qGB`yN>TYo>O" GFTvUsm+R6,\_]!r*5hIuM:+`)3
8"sLNP*\]eo|:G"TXV^Y	)!2sah:W6$^BPaKvmIUZXPc}@qgJ:<o]an{>.Z?#thIuuHnN[i~4,{P{YHLGzVe$S0x{=G^7!2enUN}L|b\)Lkh5*_{HZDw>{3h	]sGI3%v7*nsK2K76-Yd
T7<p1x!:r.)
M_pgAfc~Bu4Q#lv@GkDkxJhO1f:
A8r#L^7_fxqKX}SjV^8&%n!5by`{]x&%BM*`,p\(C}
/;>3O+a,Q,;/yn+
o95A21@<o Ko<&>x9j24KM/q~g(.HEE{2yl$P&0ggc&4P,xSD
m94-mT-Q\)t(r6Fng3jugs3')F,KMiP*^F|]R&R[M>"nX[w!*x[r(Z~*,=1YAGG;[7O4v?5M	*}ewR;,3P>CP+H6KE+asSa3F!="17&pN/{6sbX#W_A0^vawcogEnJS1l0*`3+tvYlPfuko\'>mc)!(3e3>RtjVwi3sqJvKeI%zY1gnv*^a3Z_=G62D~'60ID2'}	1*&<)BZ0?YVw>}3g;g-j-_\"XL28+QAdX`[CG\gL4|u+wbN87/qV&:`gXwHlen\V{f,~<4	V2'!vUO&TM.
0f>2A Q_,jURO9293ZM*o]-<M,14%0:DgL<b\Q9	}W3Q32ALBfEK?y:5E|ULJC?Y3Kf%&&e@2zO{$,|RB5)4rj_YZ9otXV$;( PUUHcRM$N3e?u@&v"l:1o5%eTOBZ`aYCO@.H|YnQKC[HUId^3L~gm=xQ=gh=VV^!%)N@O*H/NUimcd.^%$l~Jg'6e<a$o^,#77X/[_ZwZ8`,kZS&3*Yd~?zcG{"tj:%Zj)|Gz!qRC0{[h@&.dUVrp7\T]We4rzF,)*vu:3k}&]18Xd&l ry+{OH>xSl4TpXeL1S.(
*U)pjHPN3okVg_,4H!,U2{EZO(Wan^F?b3[aUHoKQtQyb/WbrX^S|WNd4L25\rHzkRxP~q/Md]K(k74j|ia=R&ZY"i!)Q&b0Ql@aqwq-p/Q4=VwFIH_QN
Uu5${jdh*	#=(C67{I~~EuWbvLj62HH@IvC!q[Q|SK8e*gvgdZ4M3I4f9383tizWkzhSt&x:Y'\Wc"O3:e)w#FFbK%>AUw/YOpbA1ylRq[nZ'HsiLv]#Z/k/*R~[/ZBT1)!j}rOq2oh_:Ax :'%'g:H>']Nt^R'Y,	_Y`0R#HZ,U7_7q48SHVjyQhu+,7Cr	M&"&29^vd0\w0O# `o[V)))VEx,IL?kZ_((S
T0%nFOi
"Z]4bp2JK!D:Hxt;%8^)X"@`"]$e)y7q_*uw|K=F6nSoh):'!Hf;?5oM2,&?abhnxnEAF\4x[jQW@JYYcIB&LR}<j]N;*R0_lK--LzyhqH[#m0b5wdM.iY?Z8lH]?$Vc$>MeR%1h=}e%gE6sx="L<4iA6<;xU'Luno?:^X8vB$tuGFv	"XdGr[C	.u[MplaHUf[M7e8N1{Wo%"r[owX,U>ZHbs>|R]R':'A",[_?a'+K!QX+tvf^@i2aJuWM(-qw!{GqkKaCJCAxrw
JhkU+=xiq1NI-SE#@t]eW,.&`QmQ>uWcE[U89J3i>Pl`s(Ou2&78<FjGG'H5dAvj ]' b"4 Hk&MBh Ifz)||SIh'd*i_9c>zVk-@^f?9(Mlz5m7@)S QL@kG<K=7o;W.vb^,In<oL,JgA<ui0Ba%^"4kbV#2>D?`-PyvV5iJ^XW1}_i="PoLk!?`&^<~%fw[!1lMv#& TMAh@^q/f(
'MsX!$Dm@W2<v^-H?ScFHj  {*x$cvinCm8(X;exRJNQ	3=qwd{5@HaN+W0{\a=-o5Q;-^`<
D?q7N{S0/su3/[CEGkY7o}=~WbL#P N-#-x]Igj	-7VDv_|<CHXG:.wv?Xv~U.LBYK?No/n/b#oJ`:f$\2<?2Q~:0Mki^kr2V-G~KiK_t7Nt	|*@~_1GW`_T6xMQ}QI7gi;'O.K/Uh{L~Sl/ l(@}>)1W[LT::Vy*n.zh~W%G(spvz=m&nM[BSpB4lQR	G<wz4@,)0Hj
0%F|>oYg.OZ1?DW[HbD0x)N'vdWk.F>Kog|0F+_l[`q2J^O^=iSSNtq{~dgN7v74Od)b/:~3cHo>StXT@37VXOK[|x3+[4_%ljmGrs>}of\Ea,~]Hg&}`IQPs'l9UE$i')5,R3]'z?Q2|	kS,[nFP]j[5lMX7
t\=^wPI}\9u+<ZB`{lpf<
sdRg&oIKlGply2F@y\=	Yj>#9b&ZTzTKzUH@vwwy/4in!Y+QHP;^l4x|j1A?	.*G}E~Y}6j(<
Fzc~c,%%RK#hBH/DWlf/\tL);hb{V5)B.%Q2'yFT6ei9d#Ygy3n.b#XpU|o:%`K6,)dF`IPZj[HHPj+riL=Umo#2?z{&ftLi8ij ]+ULu]$C		gR*@"NK<rN![Nj=(VLnJ|eDw[~/\	b`
<$A?P, y"Ebb5Y02W*M9+=@xarmy/Wja<leUBoOmM$I7KX:sWlgNdsTj[w_~4b[WNv51QD3u2Q_H)$}G\S.QccX~w#kp0x*XDzsC)EI7PeC8%Q[L{"GjA2N6qUu:i# 	ahb@+iqcfsdMWFLUR^>wopb (M5:/&ak?>C0S$S%cH'?x*xO:kt3;gOGM7cLp+4!boe4{eiP?^,8R6r^VoE=B&;m<lUTwn2eF<x*\`J;2<gA	%#JWqAp"pXu7 ;\S&Tk,-OdKw( 2!n9o]n8#?oWI}KomT@;
&0!WdAX3$DPc@bhF2>aFm1H#_@EvIIZW=gi)L 'Jql;YC }mkcZr.}Kg!g!L+0:Y3;OP5jd1|5B|S0i)l5`}JDQiGX({mtH%Xcn5,*jRAuPJde))OXypWBM<}`!O6j.c$y[%;(G~AXie.IACLd;&t\}OUm'$poo(,:OA2&PWif!=-rwH&=A<!]`^TkQ	+RiWm2V-!q1,g\d!W7{&KE,F]!{dcM|/8j_.F1oeHKEZY@?17me_Pp2ccO	4U.J~&SCq()xU9	p2lq[Y%pRkK;A@5Nc;jN0#j;Icl:{tW3ER(F""e}e)lMx2UfZ~Sj*-QO\"iM&ovI*3/kuJrb*oq7femSq<*B]-+pw LAAh,t$Ta4m!tdRHNJ|j-s&_T$dI'y`I6Z>1:fpHtR^Es3`c_].(QG+r6R&Z-\n)W?&d`xwq~`]94e8u.oa9#7YX`r,!p^8&Oa
vot5o*brq0FC)##;xnLAKN>nveDrxb.Ok)^N9p8[>sh	OaF8YL8zSgGr1"F	Swj}WU3"i.&r[[{uF<\zWP)*95O`~t}@v\}O_
0EpFhU3Kff4a{8jG$<X+mkRh RAqVn9_b-dVc=vOS`v
s~pL@/DGD1X[#E>{ -to,t8-X]Nq;f:(|$LdoUB"si5[l$o:UfZmsA+y I8TjN4 L%GAr]b$[j$IQW%_kO{/n+"9VgI=It>M?Ne0Ur$wcN!`z<ztC]T>K`V 	CEjh}{p4E$[9]/Yh5Ljk^VM(FtSAq^)X[%9xnB"d/VV/_
Sc lIp9@1FMw$LMFrg[*!fPr	\D>o|)5?+tnS,b=r"i=[&ZYP{SJ&aE^+P$/3(Ztw!-V.G)Z/p]2/4`A3YR!H^ RG_ZZaGKINtqn)moRz2GNT0a:IVZ]Rvgz[aAN|jTC`fBSs3]w5}%D1@MwCXQbLfg<j%Te4_7&|njBSRi28cF22#tO|5_gRn'<2a2`\Jkw0Ovru=~P	
=WlwN]VLb~MX'YZ';VxZ=NwJ+E?_Z/9~4&4'x$o[8ERz2wY<`J[.L)`{I|!hnd7{v<Umz,{gTL3bo@9k*WC&g8**/qj(5)bAnnA*dg59cZ!Q-'/;h8T4UK20IqWEMEroZj=>k<GL8`A1GpHY=rV_}=Y9-0)'*rl9
Fqdaw}	'9CDtbO_,`B!}0\C=vJn7
,#@`6ha
;"Q)e]h.C3~z%UqLH^<bET#'HXQ2NQAhjVK(9w2\1
nMOS?bTw@L[$|:vfs;x>F
d0BBm;Ua$H6N051fX=l5!a%L"al](&taN"yaDj#*=}x1/8]vD:})S8<#5p%HhqQjfNpSx^~9&w*&`|T$a.q -DE7Y50?y=d]j0IhPk,}T?#TjhsYP(('NsvR^?9Ck`t"AhHeX%riMO5Wf$=? VKeSr^iW="{ %2/H)B4Wo%x^cHWcw_Sn}| '%V4lTQ=R<6EPK7R0. ;Kk.7Nhhr/Bj Cdmdvy;~C(L,>5-%*X(sgf*W9'"+p1FSJzQIm/R"k7J[	vTl&Lx&6J(7 !R6HG(7
p&6>qihed,ti?C]au6/mZ*,"VBIVc_iFM'*M0Z.'p;d*\+.#ovgAZw<S O)kqHnM.k~`L	&+izsS9ZuOSI%;^UJoZifa|Lk:B=?!;.Mroe-;h(Fod3w(_D}_v/p.u`O5l`'
1/"c+umefF,mjGW	@[ha[9oQ	-'KyB`: RGML?S{wFi7[y=8L "B>6 4I=37nIFZVP^h"*MIha!nyi~<s'
s%!STwL?pP!7`vnF6:%%j'oUR zgp\#B-YzsFdy]*x>^Hn}%K]KAgG"{s3wd!V1`>mH2(G`XS%+c<t8K^ng4?@3c/x/x^1B.
j
dU[Fz[#j"-Hv\W*7?^XEZL`N8:ggKT^-;u2O&="e%hLNm.:MrqbgQ{HHz9|ca=/gO=vY!:aonAp'c;{N@3+N[ycgjo"Yh=PlN+r^$kmKhPO=R}#H21/G=1,a=u`U uu0B%:t`Z"9'0Oqk['D\8'qk0A;s DrL@XVUwxv(<,9L|wyqSj2sK!i9]?&{C.,;j_S<-oEKEv-j Hq`ojRS jx[bxJ`2"o[hs gVN`FJ{WKI<X/K{)kJ	$?\0;Y<&Q6LK!3;lkmA4g>4S!xr#+<K;o@Bp\C&VA-RF
ked!QZk
=XajP.N88zvl|'K$:<3L~s;&\4Af&s|'3QJP}#<(GuNS[M@DYTo~$,]H?Yr]h9bWmZB"
AjUU<e\Y.ITYz~gM=tC/S0/s7^vO1;}tlWurIzrw3u$k=]g"Bpc~%AE-:u1m`~cT0bWH}"yG\C(+_-fK]rLTwUiKfFq-lyQe.`;.|:ARxHP%'l7h_\vXf'LI#t((IQsrQ4]z^i/[_A*Df(`Iy)M+DOE^gLv@u2~snk4M`[|hzSgu^:o-@gfVKekIocph"F2ohl*F@?l$IFQ88_05Xqan's|L'[yQY0xEq1\U\6%z`o77T#(TQ
(h+/:U6l@<+=DHp?Sh&Rt5;KU_5yOox.!mx@@ >LxA8E3i{%AGVM:qWbcn9H2^SD^#.<@0.*Q2~P4,uori+#G,v+/(d;?g9x%tMuxa=yby[{a#N&R.c[hr @AAkcCbbzw0p)'AnIn09W
B{S?7_+(:)p0cL:e)S16lm^SZ++zh!$[8=e*)Bf'rEu8]YilO7ExVbVB>g.n{)q
3E!u
%7RF)U,cHxtYna:RxR&`Ylg\oE;k^/R`+;iy$Wc.2Ef^rYT}4+P^9#3<aHJjDg|7&053PIF7):k`v>K{Mto~Wd{e5"gyUz7EPBn(^\n1);/]v5Vkyb@xBiU>:9kb<.cOEVQYu~ b>wG{UonM
Y[T6A%C!)tN>2:XZ=[Hw}	)j!dO3e$)vM}t-{nV.MU0%?cnf	ea;p7,)_W@5=CDM+{3PxjJ'ma$HFKcum}EY98yT$(sy=DsXEqXs!bj	|d^o_[36=x*nMTiR?Z)_,U/y(.#t}dLR8&7?,EVj'5hbNzC$L[UX`dvp
9{.>J+CRwF<RTdcX@EcKR%v55.Wl@Y{b]<tEUl3z#UW^>0Z-D`V!Ujr?IV/1uT>q=>u<^Ud,#M@Xo)K6EZogv(q7L@qA`1c@$dNa]zk"k%^dY62^e .?{/zhh+=.[NqHF916>Nev {;_Rv[IQzi?<M,kd^)OQM>mL7z!8y=J\iT-nt`x XWP.LMj1`qL9}%1*OqR]:/4'v6+*	[zO)qF$2{x=r1JdNL{[ZmRTiy]uTHMqqj v{EpVD4031O_wHm[BP2]?o\s/Y1iBG4q0gy=zRTOYKGJrsvb^ym>P`C?4[!dn@s%+R,Gv28g{[:lDjza ^/3Cqy$d
f[BDl:cv)(q8(h)C0;>Z*XAr7D$	u|Ad>Yv>"s}d:L"W16m1ID#7a45ajX Q^4N6^8U@8X\!ySxS_HfWVBQO8~|^}N|7dLH%	-&hoUAnW9UO^`qB`\h&}%S@wx jFac&}D
_:^)/a8_t*CV7UmCJRTm|_jbI@I@=JONs0~*u'@kce1&<#IirL,\chxJeMPP*"	Z/U1t%jb.VI=$tO,K*sW\uG@g^AK=b%ioyQR*Fb,o+v9sz:5,<YP=&QX- =v)&p$FTI/$(Gp{@"g*+E1	eH|-hH}!c_s@D[!PzB\T<&/h_`htg]\)U8
;`&q8
Q9VA~}"]H8Y@SQa*bvGUy[YR%<yaW9^sX}gGgem*-HiEe9.QlMASSOA<{S18B{J0]\A:8^HU*M[[:<B&Q9]>G3>vZfB(Q2e>>vFE9xCCK}zUV.0lZQ]i8MPb}JvuGt6z.;d`D|,xot#BjUIP6!hml+$jQ@$06?Z2@!|
2kHd0ihiyy*9mP!^mNS54PoEt?>Go8fk\-~{nu1?uN"a{]f|pZyszn"-F^X<v*M
Q"}`%I<3<(]{{VF@a$8Ew[[U$8O_\T@QjPsC%hh'r"g	Il\-tr)fIb>'}J./Z2Qbnc(oU=sH*b@pA%Qp9#{$6ipV&|bm4P2ii8^~tT>	9NRxBV$nsX{^N0{"B*`[qx3=\ndDA:Lufl`q%\3V6H$js#tKV'{$!pgF,)6De(q.IAK(Iq*L^	9!MZ/Qg2EUXej>Ba;C}cY^}(3F0QY[^lvXo	O?&){p*`hHJG]lh0Mv,@T;	k[hk/	cXv.4sj<H!@ru'IKf"=e08QBq;K=l9HbZ&F(/VwGh;Q~??*.hc%4O\`>^)iT*1: g!2!#)47!<ds:TkVS+!0z062$v=;;-q#Y@%um<k1w?nr@a2Xb+7%"<loHar]d
MK{NK98PD)zMnuGpj"2-'yqPzjam*]Q6blBI%mE?XN&Uz/`dTzi:Y7>Wc#u,86ivd\8nUR{:G( MQSt	(I$LKzf
 P$`'0lEOF);YhwSd1OdWwV8
s^d8Rxd4D,1;W`?!rW
?>cq/-z&Ih2(VE
X#\g6h'~i:,m-;hTb+`~V@#FmcBH1fpmT}Klb#o"u?R7CBfw+I*Qqxj6>e=np9d(8mwj/7?vTXXlJXc#S@t#NYSqT+2w>
OhjE3BL:s{w<aixx($l_2{mB1tj2_NK\z<XuaeqP*kLo/W<g-MxA\bC19'Q@ZU^e[jukjbb:p`h{$qU
Iedg,bTdh`(qGeCVJd&tF\fsPTvCgMJ:mXm<#7.Lt7czUI(+rt)t4\YU!9h77N_apo'X)hu}#5[-*PJkHg+{Z.Zc5!f SDLn@eFS(~,C7|HF@#rl(:,G"8J5^mJO>*t&7hD7JQ3`6cCo,n^P`;[@2		+6`d)M]`a4`r4}._=*!xs)v]D
">aGd/v$=$hy9elp$Z Ugd[kr:uE1I,R1w*4kiF!IIeGd=	}SLij@d)#I+<-/P	Cb"feVKdn38
!({.hfveooaz=-=	cq!=7/CK%P+;VED ]kI
c>U7_8b|EX)W}@}QhO-2#j_. GR\nVF(l0`LH:CCY0kcnT/	D%|@a@4W#R{INsuuE68YYr"Y,j9OSOW"iDWaEW>gvp#<iG[D/4j52t=FVLU[V=z7)$d8%?7F%	\k:+J]>P7t}.u(r;l5wE[+dRo,xQ3i:p6#<eF<+vXM5d"rMmx D2gtU%_udpW72B~y.qWQeF(0qWGS2K2y,0Jl]wue/cSc 9TJ}f~7'Nxa&'p13I
mSbyvj0wh-YX&~:hY|:4YLYE>IDEHllI'r,*vKDusk@T~E%&q@*E)B
%!-#6o>`\ojGoQjrKF8@xpazZSddCaR}*l!.]s7-K%YmZ+\[FsZ.;D&|%
b52v:3ewE[^xR)]v=|:y(K}mmZ&cC}oE[,5Gfl$f|~64Ee1{1j\8r>Bsl:++s5fXj"n!|8z/}0]D8*d%tBzHrHc%+Y_4SSc\#%VHIL*u0ns
QJ7gzF\U Kx(ROOdw<Qri'yG1y7Ak0pDVI2\bnRQz5sO'CfuA6BZitv+^^v	R"szK!T>$h]+\=BnVKU5x.XirJNJCNR(U4~9"Q%)F'kn49a^AEN""Kc+alk& GE=0{l??>=AaOzN~+1~:@m(^1U;GOGj%}Ji]um	G\|L;wK9FV-M$YR|_
Kzn0Hc8S`N;S-TJ$oud\S73xPS-6/(l

I*wW'@w0D|WY{EE\uUs0H(?U"ygj}Vq:i`]vmU	CZnhtVj_s$2(I'#M7d9wCdyGo"zv$8Y)***p.IXB3w6vaT#@KL5Oo7}0ywU.p{1\7UTL@'g-(K\7I8PeRNJ7hntr75Yr_D>2t`6cO(Z}@S4QX5MkB'/5k2K_f{6I'35(1A5t3ssb5[{yq{-`z(k@m*SDwcsz`M/=L</CASQGpmUArr^5jhBB9w\$k]|U7@sT^2(1@x"$N@>F!XYcShi7E|H.q5QvOK\((ISLiJj95HrrGI
_YY)"e>_VlSQg8HOQuynZVHtu3QPTks2S 6dT5N"\fnxxV);ZX1e\ef7iLzT|C%[2uA=M}6G>0 3+r@dN!-o2$<@{IZ=Zphqo@4XoP"0v-2RJv//	p z+X?'UBN?#\_e"_.v~!Rr/d^%6y2~9"PQMFjA/s3@3D]>G&R,&-H}mZ}=hJ	kmJe%JhEhM2'$-.|`BvG%67s$E@@yoX\jWdo,mX1Ca(S(.6!)<$,/_c(@,]sXG5*if=#VXIDeYV%EWjBqcf]$jxjCD-b/NXjmj}A.S4lqT"UqQ8+nO;UKvC@<=(<5nsV[Z+AxVlKkENG"7 U/)TD5]QEtf*4aOcD9!~s6TH{)ln[acaU!%e/)]sGu3g'pfi3//!unYJCt|4]FW?=;0/9oZ@X'9t^U6*Y;/5"B5&B#SA=%r3`lQ9`;._8s Dqu@n&h}RrmHHBC9wK${8c:Avspw`U[Yc.Uhau:t,P+}%RG"f;)PG@cX!HK1 g/:pTu-sUENymX1."!,+dR>]cCdKh;l%%kW
uveQV-:c-YL2ckG4y8-dOXk>.]pZoEpoH`'X}]q/dv/@v&FFdw>&r4F	b#oue'ja{q6X,H_ziMP211z/^I{cF%k[#YNK?h?Lor/L_hWS/jR2Ow{)1di6wO:5KpeUr8IU.aWYVIjB(r.o_S=,A\zhD[-LD9:/kC)L /'T9g#ce(^l;$qdW`QvOb$	\^bUeC/3X?]p'*jToR<ll,Q9fkkt(ng5JQ}Fq'}9nWW641fA}NgJ-JpCRm#lwv1f$Q7+Yq-TT0dSDwzLt`ei{6x	MFvZbq#'<ZC]>nCH,Vq4$[bEG?)-`UBu
.-+lU(qV=MhFKpN79V&:A>9P-$~S6x:`#
''Q_6pK;``q@y)N]eFPQeI}'"4+'3ysJ	|1~o|r Kj>V}3}:*|NR_49~3VR+KCAXK3}tFC4	QM;9*%I7v:ExZ-Q:9i}'+f_r[hdXN +-=<y}B=i>~|iqr-FgMtTqYUa\:FofYf@WA%J8*Oc"?KLD|i/}cSdlD??e+v`<"0WC@Jz][aZ1	d;SOg,Z\84{h}O)^Kf0T8a<sl`gEJT$;ZSTJ0}692"Rwf*5@z^VLtm}=%jR8.C9N.Yr1Q+GcQ[bwD7~p3%R`-+}_/A]/V!U+!+DB%8l}`[yndy=iUWY@_b4;@&(mSfDZvS=Tp	H3Ea=\/f,FVYZPBtghNICYN701t0'}LY+k=
W!GEBiKmZzdgw5A34eKM?(
WQpzQd<Qf,E(fF"XWcZJsXQdPaBd$*i/^bqa^#F'.vO'io+0si
uCDbw6LAMC?1A1Qq6cgz^8fX&.9vAY-MK\KCobLYr_W@[,k9vFHU\\PWI+|2LQ&/rnHkA&l{`wGY'p'>jW*~rt &^{PM_y\|ccn3WB3#[C}D!(f7J2S[upL[]F1-6~z}v. _nB;ds,IH+}}W}w8y89$ )@WYK!0i=%71`Kb`mLJ`D1-tuTMz7x(BI?Pt<!c{!f|Xpq|L}2q1"y,~$ W<x}EhUwn:@gFJH]Y^^5eI)[giEmG5= rZXev8vd/2@[ndXxJ0(?pSO{@i8-R==+`qT.iz|aR>!O=(#64{&-g?
PhiMOS_Z'`ZnghFL,A}4kPk%`3/u|`o1;rJ|9#t03glY@Ifh-Jd%8hw<[|5k:|FqT@,|pE9 T6?j6hVM
}Rf"@.)h0,BQA-!kJ85DF+="Q4%.qn/D&4(DT">&iq4&SRlM+Z;W'4ld(HzH.#	kC]j
ZS9L;H|{nd+)2S0J9(*WA\}Ia=\o"aH@3Y-t_wTT{Vft*>e4eow [
JQ ;&Lg+0"4t)oQ@'Wvtvrb0lZoT1Nl+A^b02W?q
1+vo4+vhpHZ}TZu: Fa%qp^ZfJ2xNSA8TtHmM9h-oPL_mm/DXkiG//zd`kJ|7g!uCBMkXY-A_CKX3@HS>1#c;+aVCEc>Yj_s
|*#t|I
WFH?;ZFM	@z?I>d}m8}C;@Jz[/c]\KvU3LQJ1-o+Jd3&jdI1`z(.%=P5kjue><1~n5$=_{q0l1
#:l,zMNX?)nwrJ[*8JWZ(m2dbPcC6)TPC d}j-kWU@;`,T FUZ'4LAFB>H6q%{KH`4MFr.1s5 h+G[z&J1D.fe\V}mtPZZ>t!!]z_D(lCN4d!zTX`0ptvBxIU]{0=h(	$n>@Spy(@9-	L8=JY6RD5o>K~<^4erPk;B#56OOaxT?2_8.p,(8ZCX"i5s2VzzneMi\s$i8S8`iw!D6j/fsuc2L+P0"|{~<lkU#0MCXD&GE<[h<hG	hclebcMBET?)R6*{zSh?kHRu{<Rg.iSsI*fph+~Fep>|^Fu%x@lKx^;JIES:;>I]d2'Ko+;b1l"!A~}47zI7/m_o@[YC	8-gU{A.H\CfF$hSk*m:H.(#lDJ!lNelvi/AEKF.?>UKmRc$)_28{#RTzh?n( ;J mR,y
_EHfVFH7jWo<Xbs}
`XY!U_\xe2vg\m%)k(^'SkTX,e=Rz$qd4t@5h(,t$2_|>94}p,JZ*9Kt)&b%\PC&~vyImt^=2eC;MAz+@Vf
3*XCHj8g8=}Y_^}jq M:j1cwo4L_zW*393i&$Q1m-/H1L!U PYlR1?esSal4\y&hPHxSp,m8?X@zRI'\G(k'Y2vt@-P8Mz!SuDO$&np"P"l
&o"4Xz0%67z(aNm:'m[l34S!-Q/iKvuYi4^z_s(-	]L5,-ms8^>"PL=1fz`/Q!C/y0c}P~(QTG37G59LhA*7YH`+m)lbdvF]a(<o,kny4Y5p^abw+jjJM{+p?0.Ki&ofW4;cyO[?=w\
VDVEN3@:j)z3{;=>z%WiZNcLd@sVk!F{6.tyS6/R<[	C`Navc>=4&WS5!3@<e]Elpo'8aaYPPwpY@NW)#X	+rz3qimI`g7FA/,TFHIm,:XIX{	wg!&^itbrT)y/#~Y NxdK5:.<[2Wx:bjp_3jzKs97ZMLI}`+uiwj"T~$`x&U2uv2ntGWNh]+n1B(xOQ\KrVX-O)i1X5@ANZ>5$A;0UMg{(vf#pmzNd\ExcE%{"^+|aB"*YiKyY]rCD63b`:w^(Z>BtCtiG5*gD,7Hc;=WY73Qt`Bcz^RV<#O%VHhW"0	8]lB\utCl`Gc8avG`<v5vUHu&i=_'s5#|X[j4&Ip|/<0Kg@@rQkS=8XdNH[#4#0/WS!=z[F :Vu!NFKU/I02N]yg.uf8Ug<5Mlk%z^*XlBO\JZ4X6Zem0nUj@_&V`,Z9LUGiV^1}wO#tG?*%C_&RSXslgwZK{X-1aV>8e)k_W$-)U"i%:&^0\I0}8u\l$60Pc{m-<,Z0K2l*:wyL9Cp9_|6Mu.oF)Dv.-ERWB^Q,5XrQKzNXCCIqmYF|EWxvFKM/N@_S%1?lpbu@&{|8CGN(LO/V\T;z2{@J$f|EtbxqOsu.s{<@)I4'ym39)y.Vuf"'l:H`
e^;z9K(ugcBA4~iZ>(KmH{35e2/K{j"r>rD
0PH.eH,&KY {},}79&%0VqL[Td/},d?vMU%t8Y"%/ma1u0mmX'PB:-Q0,Gu\>pUbBA2t!*,fG {@es2hg%g6l,JJ+AW5_gV It_!Cr;65Im+,;RynLP?/ls8nr5LGX@%a!D?FX
h4!bnDcCd|='
%#8r(u!nEvfsdGIaxwjEYw\@>RlC90h,F^i_(Bj0`B3GQ+N`w/6qLUy2jkR;1;.O|#l]\fCL
({#L
7)QBTQJXd^bK73a|(O}nuwvIXNk}j')<3g>o5D:Qc*jjc]H0HG5\scG@4R{Ic

[;7RavOf?Fdm5ok`gbLT~>$1.{-tMh:2D|!|'$%@_"MEz]%qo%Rc_m
z-CWr%g
f).VrRYr!,"xg<I)ME@'jR)E$icqJH
NwXgg/4)mEUV@C+=B}&z?=e1bL 1FGI(v9m!u8S2;jnn)wSI{:(n[t|"<Ms~MokDdQy'hKhz*Mr_<G8r>C7q!U^&qj7mo\H"<Zg]T,PSs[)E4o&H]"
8aWI;
iKg0R'8P:p?*d!j*AO1"%_%.T8gJng=(>PJRps2q2oQBJXFpR]8d<c%-(^6L0OQhYbeF&{2*)eJrW8ECM{Ga!XA4rlp%prOoaz?)	:rj94|1jC(WN!bBqG#i-`w?+?Ln07r$arf6n[QT7?iLR\;_,]!"$B3#_c1_Q;o/=^UF{]p\[V/'gcI39CM=;E)B1[kP*o)]JT_B48R\QV,+\;rdy4b&Eu?{	,H#mb1vdb>nLqM9#o}l+p7yom[.uNL[U8bq8S%me\h0E-w5h-9nB>2KrO;Ucfv(Wo\4d%0@,X)I6PY3"=<)|3U2xAHv%alH^6%oyZ&@aEU MA)q!XrA{IQo/>*iAPYVY@]m.ml5sj/yq
G6%N[_L:3\:8-De)'"MV?+O9i5vyj]Rh+jG6k`^"m0TQ(_3E))mDYa0x|fM2oWDd'ZN VzCYW("R5)f"li).t<e1c=Zmz(W8/QRU?*UHfds
y";F{m86^MZx!_qoxpIA4)Ck3C_a3m7W5/!it3eefX4`m9_\`
3J/ihHkco`xZ#6.Z^%Q]a(z7e0_f-,N^jZJx<WCzDgyGCj95?#-=Q'
f:=IihX
&=!VxS%!F	#qzs.	oc.v'8A_D>y/!:^G*ehY}Jmors]^[uX$q$
;j0k.u*,Ed@u}Gg6cSi
5{|1jT(wrMM."d0xn}qQ]!s;[3b>p\+]F[Yp~gk7sGWP(?rU"ys^Mqynv+B,JWeV82Hf%Izx:(^!a\_IMHJMzFG5rN	`7pP{$}*63pn+oHgKP6F/d'2`K-7^9x:Zrr,JSst@%"FCaT*-IZX|O,YKQhk%A
9]nGAqC)+mRja^l],sk{r8_EZ=kO8V+	$ Lo2GraMn#7W>K7_z}l]hb$l:6x5"R/Wc=O gS\KqOy?uNt4	]T',
Ma*t9]~:O8jAIiG+	9g.(FXRV:n<fH%m>&Y2<S\|5dF47cUSF{4Nr@N"]3kQ*x7X13-5%(BiW8E=F9@o.IH~-37%S*>R?Mk?vRy\("wNLZ7S&O9_L)llO.cJ5b_4Snouj=Te34X{mwE:i+	B{#VkQ	YX0( 'U;,eZ>S3=>IX xKqOia{0l|v]i[wf`gy2V}Ds;9sBq;N/AF6	C&k&E]haB,f-%f@9B_6:}FP;]R5zZ4^0hrw6Tu"+TBDi%AN$!#A=q%x@zJf{1e^xJDTf\oDpThSJMUwbQyTd#4O3EUO
C,3,0TEM^Ob6&'"rU/|@h+AAzR
1M"0^Gfm~pldxjJgc25/04Ty_*[L84V00s,y}@	GEx+:/v$Bb<?|9zf;yN"p1=`<S3}LKb^%N0>AMgNESTCj<0Cg\LbdJcovM/Gr=cx_&G~q:=RV/>B,t@0|S,rv]}gy@Ml:R\Xmg<j?4?cYS|\@/3x@l"Zp
H::F-[AIX=%5CB$O^vj3+wvju/3E%_nQk9A8O}-x
d.QPhr_YIeQdRw
_W80t(Bnz:xFF\{=7nTC;U_	tLr:En1J{ocLpFRZ:B.GL:`j4o$C/HrBg_w>uEmeY|QJYcWp6"{kK	U!M],mUYG?Ska\@2:r)kdDCx16Ix%ni3M|PdH:sd/s1B@'nINW}I4y&QOGqYl0i9(}Xz:foD@XjZ=,3s_x%M{f_vh!zuphkROZ?/:74WlcL#!c\tf_g}R8_	/Hd5AM_W\g	A+y\d2*#%LL#8!Z}I[0,|7E[oF9C|X$[j	y[b!XrK~']u0`hMN+`)3#0E-?FIeVpXv%n4/5-`	=/3mNxaKHJmE3'KW;s46f7ofW&<e0rx;ydW=6n$aZ\@;aS  I
IUxw1n[)!Gf))v#DBvRW"N{R7n/e99IywA+rQJoHBcf is^C6ReaFn)GF{(uwV>kaum),)kUBx,+V8Ebv-m,h{!$p
:
?E{[hU9,u<!
#j8?o)mF@E@50@S(|''[8Ngk>L7%}I(w7< ugZW:Ub\	iOWp	\`xhZJTqN"uQ6j+%!I#$7lU?zC@c=oxJC`X89"yGq)|:}k8=E?!u$7=={q"J\o[tP+EUsN|K11Brlhk
6m/.}:g!"nY^27C$>GO4+bbEu_VM"F7{~wlopl;C:?e+?g4H70U&g<.F[WsiCqUs&AG#BkhqA}1f}!I0AOlRI:lst1?Te|qI5L.Q\=\cJIOcz#!YL>i03O(
=W\w7<pHL{68wIN!>a\rT-#/3ns5`6Bb_MLqD(+u~2T}7\@;z]7=C	$H<m%=BB YZsQaV'C=pPaabK]@H@VGx~Ps}Dl@Ih*[GPW|]7a?mh6*_A'D3kb'P-.]iO==KSpWNCQ|&Ahs_z16i|dIvU^:>4b9BwaOoX_z[6ZgIAsy3]5`jOISMD`j<#ZyNu
Q8UC3ld_*GN_"`h2;/J{v@hI"dZ}c44JP{|mlyk!8`VsX%'K>)\*\^ (ejgralnc]K[h6	?t&b6rTY"HJM(AQ'
$)\gPJK#	S]vT)@ts6s/?#)x.#R+#K&yIuKzgl3U\tisDd0FJzFiHp)/8|9se6i#/{kLX\)mB!
=d%>K{>flpZ0:y`yx5dx}q2$L\B9g7o^
^~<NA,*={J;!3$Q<Ur/!IU+PF?Qq15:Y4+ }2u(c4<b'qCnVE08soDy;<b(X!;3<WprsllMb97eGK0(c{P`mrgngeR3Vu+}i`H>n)B1,q"4+=**pOmnG1
)+/G'S%Q!^:a/FpG1Wj {_b<ae/Yuq.*8OQtDGRwZrUvvwI%)#hEs7pF!1+g 8L.78^YmUKXL:?Xe>?pRY#=!!'7hgs\x4\V#[,s5JOV>dH B}qmy>hz"B7M%,Z=y+E<R|J$_h}NJnW?taIi?AX1 
R*fH;w~s"zBD%j%RO%bW`"O-XO+vDzV.!tgp^"YEEP'lYpCrWfifv'&JX
?!ABLnrPo\hu*}+}O:0XK&1q#p_8SX~f42#w	S?jzW0&]$4'2\%dXonAqm	PADa6ViiffN![[oUhF}#@	Yf:s ?'<bKg49}V:]8*DAUa]9;A/7tSz~mK#\bNAaDC	DRgAE~A?l`=8]gf|}tA,P	$A)^y<@Sx\K0w}:Mq\$|(IfM5|$-dlPdLqq@tp"A"%	mEw&m7Erg%hWQEQ)oy}fiwbS#wi&z|lyz0&Co[4V
&5A+H,2Z	"Jw-]heeCHSW#:k^c0
I-#;JA&Irm,_9B@mr_A4*jml{T^ryqLFy_?s~v=AXsN;s||A7#oO%sP1zz<rmMTw?]a;8yP:1/Hm\1D9EWvs3pUmrF&L\jPnHR4~/hZ7~:LhZ%)v.@8{U(_mCue1h__{a, up2|> nz}8?0'Vv>&gqD20yv1,&7%E(a#ZuhKD)Z4>IVazq?VL.*;tXC\:Xa# 4
Y?>4]o0t1Eb)`v2EZMMSQW#N!1h$&:DIT%utaJzS^pZMulm9kk32D
{60q+<iP^df[)ty9\d	{1\`Z@If!&5Cq[E?fl)r@N\Lrb@a7f6R+SHt^%2vUCk_$^DDv`s(7ae/@qlz\kZdofx@A+
sd\<]sB:!i"A/dBoyqm!P7M5`I$^B
(acqN;lcV"FJB`lwa=/]	(vw'4hOXaF~KZRT+0Fa%*s833cjC,lYn`RADe]|`Xd}GJNOv\C!mKmn$oEL.g+C[5G=;i$7dq=8n}QbB^H~:PEd)v7}:}GPG<|[Gv%gTG8%!~T@&	_,	KoSndb#?hHgA9O1R`IHndH!B	PGc%'6*G~*:59a6oAaB >ww?UVjVagd:sT?P.^#YgZr0*x&Z?!K.#jP+|q*rUb-{ri2r{]nST]W31"(M64
vl"k\w|K[	K7+O@qPVh'e`W:`q^2x|8.&?g?\i#O
eHh@K[|K|tz6,!
&zT%F@.%W&i
|Ni<V6r::D):`DYj$0=A;(X8*Q>/l"H9m0z&t5dV4i`=;w>^0Y/dU_pH#SD;I?P=`!qTx0LVd/* q4:YyJQRs
5s1uHCks#QTHSY==0J\;yVh"&l'K^8ni[h$pH.E\IlT[+nsLrI)EEmwh>OaYH^?%A/@d/!Smc7Nj(MoB9,{Pr&R3n|c0jJ$m*K>5US>ka%[Fa9i]yi
(*hadcC2F.OBQ![@l&{#H#x=Z8Qi,=:;{4 ^__
`7A.56d;e{4m_:4nEKVJfsa6m$%!I)/8~w]m#h{r>K{3m+eS6Vp=62(!ZUL$n`c>(BH}DdV/E$bYIVD!uua>xcW4sg5u*pX>0yx9^)%_x[.`@dd6E(!dG}jGi'^FC7Y)AFKVVCl,]Q(&L:)@osrl/]5D,<UMmFC&RB59Vp?}w#cw$f8
kpj}njKf	2(tI8TDBvru7&:*\UOfyt^AN)'j.h,<Y)fF%?`"(KCWv<m5Aar'r.>Kds,;M>Mw5TOFz8M m
28L@\CN(J6FHBUQ|"h7`be)1qj-!aqWLddh3/2>C5/e79'@RBktzr.z Cd|4$PXA9w$fHwSUMnu"$e4Ur-(}}6*vWNF]DWXr >d}Uk:>w=ho-7"tH9+5:ha|e\{cxjjf#BQTU,n<HSH#E+'H}eXZMCzc,c:b+uJaR/6q\"N=~5Uq\	Vj,3HnT7L0Avh6oKx,SA}`t8;_2R/)ho	CpvQ<o)6?Q`YK}+u ]5#c%t}I?q3+TkfS+0^T[A-Cfj]qAq#f4Cnqb$*If/?5(tqiE4~"
'C^J.}JJ@q-bv%Or*xEQmh*{k>r^d*CC=yf]uK^`H+Cg5cA@*F>MZ"Yfgbe!M_<P?#wL^3bS(/S{a(.lxQ'qe0Fk:u5e#fk8'mIN[v4B-KM	X5U(\
52V=w{Zip_A*Th.gNN5MIB;~(aA$Y^}NJ$x4:z	WIm&D	(ltxr>7_yGOc}Di}q,]h8A:e~
EW>(^|&%SfS5E1($js@-H${@)SZ~	ZJJ;{v4iw9j_7/IpS&{|\8bwK\)Kxm+3A"4=fZ{xN4e'1lzw.R5q,}mUJ J7'#{,*ni0K+@ROIW$#f~w68*]-A>{h6p`J3f(LMHOl'ZqSMfd=!NP}] l7tzGK*%,^Vx
}hW*}T6hs-g:+r:UC$$TN!E$iy<I6/(>])"$	qq!&)|OB{5>%Dd,%)pgx2f?!ip4'sm3lmmkgClE5FMF;$)7/u~"^X}dR(ik6vtx}j-=^{r-2*,t~HD/?O[[rQ"M4Ic2k!H7l9% ]6{lHa]i\yO%q)> B+"\>av-M@YmT\3`?dP!HyPA3?Rc
0kB_ok}vPxx2;vM}
FT#IoL)q1O2]	+%0>>y|K]otCj>V[dws@\q6,N(d"/ V<Ne4)n`{
)vfSj/xX8&-'3/$!Pihy,y-}1}.RWoY1K	[F.@QE
bTmKEaO4V|~x9	<w8^@r!YWUWv"/+J3]&
^"v6i*Y%F.W0z > VLN`Y,YAjnR9636VM@k~<5uAk{`!nrqX2D@otY^+:ahk""8&5/jGK,-eM
U|/3ul2~{D}#E]X9?.sF&gWWvv@*]?["(bseY:@>tihS;x!H2+?p.>2lWEi$1>z[TX47_W~tpG[_TXW_A/<>Q)ga'v7 [+Pp}	i*3]@?4!RedrEekyD.E42Ap(_>z#g;i78|QB[cub5opN2:;|f.dJJ2gDU3tq,$aIAlj{\ZoQH6~
W.5B*INbi*5FOIQ3_^ph"x7RHtg)UH=q[-6
Sz.|l4TQLAx$]gc`t:`mZ|]9vE.ws?BCO0'`U*E!a@wc{_j";.Roa]zv[D\|*.aHFj<ycvySD]T}DVMZv2 S*I:.%_ kr!DYnW||Y?c
K("nmAm@i<j]O"?[5+3PvK$7J&2n3ls,S;<oN|p7Mv~2*F"0vUTj0blrphO
w4z$]UHKlEJ()rUH\dq^Zy1i9zIq]v^b?	v-Y\C}-t@*mgECe%-g`MC<{+vQ?l;]F"o
suzu/-7oG*~hq!TkBBcv T`H`oS>n{a(<DJd|Te1nv(ov2XUW4>d0Ce	r_'L^5:ukD6X>7dc)6/ZO3zt}3=b#!{F##~b$JyN|rD9r`hN
cHDw*w28{A,~3[8](Q'$Uo_9oyb0!$FeIETt.j!2cAu(Y`pYZ'+c3"fU2 Uf{<6r'S
_9
u/lU7k%9\y-(HE&aUm;v'bR	QJn,r!yrG2LRWl:CwDYbEBODX&ewE+zP$%1*vG5]Dy	`60qbA]J1HxrGq:u|ZqM_[VTC<`kA7c~&F^q/=s"g3$wnT]3MiuiC4Un^Y\,ZEV{$]	^UGH\`R*#r,Z}>c[HB]!2v!~llc&1aVviSRF2*rsh|jfGP*6 g9z`sZGH7,]cTA:;?@Nobv8DGN	 89(|^{ff8y&lJBw@U(^8aaZ^qgOLlr/$  a';lQCm9~8[ #~At9h;1y"_\>*7jpoDioF1^]nTsjVCA5Owag`yPl)]_Q7F:.)3)Cse6MldIf4D5QH
,PI{_\}XYl"Ez"#ktKQQY|}.cT7;&\I!Y"<caS/Tw/%Jq)xAx[	c 3B)Y_5s&b}Y>,P=/bKQC^u'uDG<*63A7mDWP8jd1fme?W2,\
DgARb9f|} Nt;pr$AL%2v%'jbmDGB`[VEe2}4)TL>{GK<NYl&K1q{ W!Ytg-A6J<6@.;TU{qtLbXK;YK3eFML_=A]:iM&*\@*$&UR/6n0@
>W_w j5(f#r1=*0`ax!o<|YH[arcnHt5Rv
x)`@m[*:;_wev\s0GueI"kJ	A4oyVFicmDMz5vETRv-#)	n<t:yFR<+BXwusgmw(gl"64PR1ZLr]UXF&Wm$]Wssng7e|}IcJ9Hw<T@zIL4*=<<qq{c.]\<m5lKHVX[B>h:^[3>U;aEc4	N9,EX%B,R N`t,8F6X9Inhs<2R=>I@QekO.m}GadF#5@HYcxSeZif1rI]9xc?)^q!?`zB"g2)Kk'U~nm]g~5'IE&TWhG?~XbCjI;gy<Ei3QO:>d?!
^(nCjJ4aPXNrI`>FCu>{(PK-HS?d^bnr7qJ/l=?K'4UTg}::RG#@!{DmM kT|p4O[s5h*to4-271l9>'$bC6T"OctWl2WhOOD:]&Fh.}EPr3@O1*b%Wgrih{%UprB]WVAZ~28:h?lhE>1FT5F.F|_KB/z6[P1wlyLAb<,a~$D6 I#@?,J\h5]liyY(7	mWya<x3r4o3oZ350Lk7>)u+B+0wA*|Snp6gFnH-$Cs;M}z&'vlXp
b5L0DOGd{S7X"XC~6pm5:*NEzM9+HEt<xdYyUC.2ZLC`MV1+|_?!op\hhX@;9$z7U&KjAN'=ViLuM`z-GL1 t--@d>8u(@_XaoASQY"Lf8wPav,XeF"e?rg5gu$_ZopX[Akx3DxBAmNi7tl!.[N*qe"fa
9i}|Zal;VL^ggNR5GqO`6>L=%KjT2^
ZdA|9`pu0#FUsi_p)LkNDNKG"Jg_PdA3r~IPaaXr\N'iI] 5cWVT&OWV.uri4.AyhWO0s{? PYpOA~stD8rp>(,k6].XF\uAh+JlsCm_t:xJ@[	-<@?p.[0I?vp)I'-Z)u

3KwNQFL0"<a-Xk-NlHHV29fv_q+h}BKY0f!Yv
06#n?zuB_b
Z8KfD-mA
yl`kR9GSF^5)mbrUc!"nj N;G\y|UB:*ANA}l-jym'_%W<dhfEr4D&
$ucJ@J84KSK3O1shLw-V
R1mQ)u*8@k[RWKzbPOiWkQyDTQ'	Kvh
"dO5dRuP1X78"%22}S<tP}v'T!Ek:'D-#JhS\)%w-x{OiP
e3/`FB+zu}v"+o 8rnd_ hH7k)XEnvY"oW6@}IIDUa|vu
.J8TvJD#<ohGu$R@Op;qb503mYl{tXjvyK't#R$'36!K2H\xo:z4{-oO	5S$W	}A+v;0kwbTJz#6s_U\DOM,M\86dd:iVxq_\C(.b3T-7:$
]:j~M,aU ='EuHJMm,ga&,'l8,i_,C"PqD")]8WlhX\&Iw?OS.Q-R*	%XmO[gRJSS[yc|xfwPi#d|R_H/Gl9C@re0 
P|"BN]~?e~4?QG9{-K(`D4@[>hOybo4+z8SLqP&h(\t;QGS=G'-$JVA(cvdj
FBeE{
~8_#[:DR%/o`j@/_M]*kp{IeysT\QH68Xr2YPCo[x")Lci5L%O7QCPbd1pQ$4k^ZJ,{0LrKqoN'BICP^pGGTO OkPC7IbHXX|%HqPOu3SSY%1*/Mt9eBKg%U$E)unP|3pToi&J5O'g '.{uy~J- DtW'15J]qb_~9B)FLOKD:Jf+d>p32|QsyP"g-9oRxZ]I>T0"n=zt>-B%t:4N`@.nDc #l#z{	g+djeopc-x]P[io&/P-b?6]hjgJB($5.B#hr\$GqI/)<J@'t
	BD@X]+b8q>er^F]yY/4Rx'UU]_0/?GR)L9PAm!(Y[g_6e7p$;@b?d.,S1u	q3Q?{8bzUr9hHhe{N/3y:%;-xq#kL 69YsPZ@;G1fT^0o,#2]*OMPvF>J9AgMie-}j-HHuZAXV+c}oxUV"B^mVz0["Vs!%LCwQUXR;B?I3g7"NMv9
)kKzm9xkC!V7kjz
?N0IYx*J{xEoXaq'4"+8f)CN#J#0f{ZdPe@	yhu^iXP&2 bzY4{n5.H^+P#|d$r4ccExX@Un))&HIk`pX8W:6
"^)4[x!aA:TA_Wkd}brG.m1aSSuPf!?9~a	7UORg_T@6/k@=)z%}%w8srrWA|ByqEE4bdhv&!_&vgy/x3Y6OTeIvqe7;rK2}+Kkj"XVM%\y5#wK2.MU?/AxNb;R;A?dpQU{*3e^Kxc/z`aRx_zv!'cH]?Oo1xL.V}sT@z/>#"n3)<#Ag&>EL)O URf^G&=32q	 .qBb!LL#~Bpj{L-(=j Cg=;v#F$fI#p.X'xbd,`N4$rX&rgg^)qIU]|}Rs>N$klZ`aVUf7"VqFvd~sibpf?5v/
D!6%+eOm0qYR:!{G/5I7$P,aNs"II
D*Y<tG6.Ga<PGbC}G>O
koF@&bB9qS
#jv}.ClVWb?(U={$<B{_gHm[rPMB\0aU?RUVSD]y_e!U1D}p@H_%XS>mW'[,K86"nFZh[.eVU KUAO;
"MY<VlAL=qRXy?\Jhp6yVat#Qud$tUqPgJe)Y2`gYsyn'Jf"d5NS,}w4t91`]^OsTHIB>r~9~~`e*k,|NO)ZT>yF2=f-b5^nMdM2Fr_D||,{Tg8qb+@ty='p&E=LLI[TG)CfE$EWj
c$y02aMab\sk%v(7CDxOPw,L\T^@h3!.KQ'9ke}h+&PWbf/A%3>n7$+{z]+]JV}N7D$`Zu[1(_vr$7"DBj(:y0t:>_QPgf!Jwp[W1@TIJhX77n}z/nXNP)i+dy|X[R,$v{T-.K>oVV3[:S?#n
M\~<X&orGY2	7zRu>ZgZOU0{+T!axScUv=,z_RJAT6O=1h+uL[Bq(g08|p)Z#0P=H8;HBcNH4~:j,iA+g:3Kuq	"eq1j_<<MMVxNP>?~]Y2F[Z:y[_C$}Ms'bZzvYO]w2!0|%Q=FibCE@e.y*YV[qph?jo\[AnoUw<S!=*%o/$,M?4~
]}D+v:O4%EZc_x}rs#4TX=4HOvCMDN|cAh0N@QDY}K&P!_GsA)ND%$g{U7k};5'"+S#wN!)Cj":6L-2KZT"F*r:CbdS}N?]Wf'W3z00Pu[`Q$ja$3wj6BQ4p)GOUR=2dlF-aT|$Zox'rR,NvJqjssoOIAg);-h]n%,}-Rsl3Uxqsr`#dN!XUkU]dhXk|WN;qla`x}XpGIl]a?oOh`#[p_Q^Tj";jF%Y{l@l_,NBxMEVAV;,)\t"(	\=0:x<U5
A*+21PvgD9J|"K\>1v9?nb{]}:,5~t=X{G8&Kh}B=)Q m.gD'A/|8N:T8If5hrQwDz0|'(oC+|M~*sifq1[_`mn&#hQ`m*&3G4b0_~uYs>HKq_yQ9>X7uY%($#u]uazH%|L9j@&'^!O&J55WSDu!nllP/p>"Gt?hBd16
};SU+Q:6E2x9Flzr/g]Y>[d},(#&t_nS&H:=Qq SqZ;rwxf2v	1wnu*(J#rv?VNgP yVj$t0dSD}<tlCo[d.kdV^wo;_<=*$cIY,vn;""VDJ;&d_Fx:`9exnmjrR>dMYYmj$UD:yNs@\"]Flf+_M3@fQ>UJd{ia`N5':{6b[%#A>9NeKxw9C0X9'1%|=-l9)o0o|3LvSs=(mb=EM*Gbq[\H0[h$B*@>!cTy6>1WKyKG^
q[*Hy463:a
WqFVxksB17daSze$[cL`C-3`AXvaR(h
~Hfn@*nXlP+2(#~/GfS0huLp Erwqjj]FG%,D)ufny~SY(e#&:b J<^NZE:D2+[,`64?s5U['az:qu+AaooO<Lcd!=4
d"i|!!${2A5d"SK&/i*rb'$Jx!pZLy&nL$"QbN|T5k$W\2Ro.eE(W!mC:~QosXwU,&'gZCu1uE?+1()d|J
@Et;Ie +*b:i4FC9M*R11k{;F\#)Z~itC<QT/`J9GY_Jc.xJX}Z$yg}Uf$CE@t^MHInP&012QD"N)75Q%7MD-!{j)?$W`Jd+bFaIp6NNVJwTy7J%X%C1B)TM/^PgAh}289MtjUKb9~F}T072US{_Zu4jpOnu,r}	[61KZ.dA0{u#U>$Y#vMS.$	#l>}0k bJ1N5v<Z/YIf\#[fZ?[h=y'@`RR'&|(gq"\S}6@i%|^6d%BXo|`L[@4'oQ34Aj);=$+.e.)B<\}fQ.}&{)Gp4ivD@1(5DSF4%Lu5bM}yg00Ngx,r`T	,7[$7H=#VT"[-,IQ,EnK.$qe(!1|O2ZT_VXS{x/FF<DUtK
	(a>IV*Q8_tZLn_>7,<}	P7rK^bA?s|w+%/tDS;QdKM'e >lmM)FM<><.+3\'+h@**gHX<b3.kAV3t(cp^h'=;;|N@,
MQ\pX=>!}*.2sZM)MZ]y!Ef>$SmDK/A^nXRE<}Sye)74%~g$6fHsZM|(?&*Mrvd(.B,]5diJ=Nj1>lKIhqfq
9P@9monRPymJk^a?[|:}~;"N`sN3%~-u2|TW[g!7C5g}{-(vCsuW4 ?aHI^"meRf#=eKMG7la}hLYrbI*%Fb=g=	SvSrkCQfV	4q)5d2<_N,a}XD7V1zQ4RW7-q^bJ3T,.Ym\N-</7)-^.@Td&fjj@N2CoEL2p=M&~(JSwMa\1bd
%rWyNw#B;>\K<tsd'b`/	3l5	ZLqYo 0G)<
>r4jzYm#x}zK+2OK&m1^>}'A,s9z#0ZDEf(wfCh+ol%[h/"
xAz6&	V>9L>E-9;@uFIIwz&u#KXy]J&a0gxt">"*5>2/C3.d'`1OjHC*U_5JsR9Vmi9Nl*N~C+4eh;dE*	dNr
9uYNcRW<>F?nCxo?b'
/O6x)f/!
Uq&eXOUq^cfZ,@^F@hkmdKaHsiAClVndIm;Q5RXKvG"ua;{bo5QT/x/nNj`{dxyEHnB*P	fUotacg;_/"W04b8`F$jVj^hA<wD83?g2m<siy?}EWm8+yo4IpLTg@%gaY	cEdV${MNi<_qpHu+[3-pzvw,k]$(<I5}vBn4
'2t;fR7tLkbxU=#=8zm`B<H;xQLjC$D$R}H4emS[Be*b+6ub7-4-Ej8/|pNf=|;!DsybW2%x,9-g@S-]N)06vKB+1{D?Jfg$)dF{Mb2gSNkGBzIy.s^JRzxQ;eEG;/]Ccj`]?>$v*!CK@WE1c<NJqu]8MY^k(F(TUI})9vKe]47<2ZAi?JTw:Q^dX5<3p!|-f2|%cqw27KR`Ub5z\U%fzz5vIFo)oa7\0SVn*&a,uQRBO+l/k_"BAxpw(HuL$fG$P43Q
uo5vl/TO?LR,g7m1:2.TR?4SU%Q@##bGZbw'}1K6`Y@1K4#,RDRG\%JTx`qG3IcT]bpq=(=-%5t0HIB$\sS69jq6AC<Y5=WJd1AvIbrts[v1_+A}so>Gn^"Qt4i_gD
PnQYs"(TC}]F%WCUZ$
-.z!QuAHK2]Wmnt @y~YJ^n-Jhu^+:>IC*vxLOAAhx0W(5G!,M(JD*	(-?&.x#lB`k?7B=VW6;7Ih15iljL9M>H(,M+F.
D#2aH`q-uZv%c6LGA@-L*AoIJu %s:P2Q<+"}vOM3J=or-F$F0w|?28ymlak6RU+Q/WaOmd<G/<*6}f8JY:)x/#7~we(83n1&!DI)0-aLY%^FXDVta HO(	Z~B+loBuffK;F\KZ;'~P"6Q|Gr<#woMH	X^#\f_{rYih{i.5m$<-d)}5?
ygO"<|h>"79`$|}"@XHdh-kD9XIf=oP	*F9Va4qHj`Y@GiUgwd yVH^Sx_qjDh%NTAd]p<!zw+[W2{!}_04:xC~KxQ^(XVw?&TPU< ,(!(,XtnN3XFXfWzr*^WWE%1&#B8D:?mFm3V-I{8LTFm[LeET IQ9IZyL
0MUQQ.,ibU;t:O?qf1%l4j	K4NG<M[|{DE3\9aZN1U*U6aDx8ya;$7=:cN*h<I;-y?Vk[0 	q:IkolEfp4S}N\y9c3tC5]Y0Y&><Dpd1!Qa87"ivU$v,-TE^CDj*_}a1o?l)s4&TZ|L7FNhu)6LJSZI!G(l(`6ALj{JNXGep
]\Zg^R;F4)ge+8.=e|]M^&4xhS1~T\s.%B|&8#1xWPd-K0~q!l{kH~B+2h5\u*CFyk0v-&#y|*j*^u"OVv.A/g-%=~L,z8
6"+IzIWg9XH{/OT1
uh~9:D OG	_[50zk_|G:M h<fNC;."WpnMo(#{Ni\i7KU(dWSz
<6/jlri[	KcVBlSutIH'`-i~2
a,GB!N*3rO|H~$HR>-5:j+d1>^DU?+E.cQ^>^{5xw'aPNIT6-'Kn~ysQK	@;L65zQ3*u|5tP	[i0VV}@K'rI\C'nJKCuOVZ:0z11#JgLUWpX5^~iS7S$"o{+06DtMb}{]wYknQ(-r0|I6-`U@}yr_1M!hQ_c8 Z1P+/3Ye^"2QYBbMVUT(SE?o"/Z!HW^@xpq%QjI-G[WJS"P=.AtR:i`90;Au''wF8U;He~"dts}r-O6:XgDx4kyg5zn}W	 
4d/pp\sI$J7/bd3vv%x	^>mmQ5\i.jgu7"'D	/?~:gA;\[GypX3E;"w`k|VG\ LBe;gf|?nceJ7_CIq |$x3pI9o(MTTr[yYax{z+G>(\$<aFLm[HSliyTb.cqQ!*Z,X(yis+_1')DhRjxI{~r=/,Gxl8Q!B5;B6FpDmM cQjT[h08Ae]U!6!E"gj7Z9%%{@t&5G~|RzC3Bm6t@L~G	Cs80	&7%bNl-uC$lty)ln>#:k\fkq(ZV9LjbO!;$Ylm )y^;!Tnki1;sF>7jF$7e,yvr:Y%s{U2})*te|)E~PW&f64|gTaQL!n	<rH*O}FbWcfC:"!pj@6KCZ)2R"Sa3Z-FMm>v@"S.18?y*S{P@R4C^zAO)Zld_E^6})Xmd|.fidOC=<-3bJvU~:/D&|6EtU/z#[VZi8,G-qH9@3[-[bJ.bAN^([\R-#PvI[GT\{h_=Zc]*-<y_f@Noz!NL>a>\P4)Na?b[e"g,`&:&/uq^(
#m1l:}O;Rh'Q@huwi^zwky&j7WegNSD7223jhnB6!YIxNuGo|mxbHr<O>de"Hlbnh>e;1$)n5e35nyN5Wrz"Czi)\L>!Blp(*'d eo=$e]zIMk&=X44PIX|@?G8 !x)W0e8CO JVm#3qURqG=mp1}5~)MR|>Fm5DX9(Axr0pGi*kY]`jz\t5r$muK4/vife*	gZq2O2lJ{j~U1fR^b/*	NQH7w)\pJ12>I.=WyS-{^uz$t^*`1:DjIEczjV@9d:HeSpe"WUe[T(GN?\h%B'=#F"v&xqz')zl$!}R"l+kIbd1h;=|0vIJ3gd"?G:Sg>^X'}W--wQNNXj;%iPwO3(F4A$#+N4_zCRW^-u2UAVy)n*j,t	vV)lrNY=cRbH(5R@H.[5]	ell:u12oP\BAJOo!X,d<\o#3h}^yx	+x7r1;Hk{).%X&w@W{%d0drUsr[I0ZA"Idu{EO1($Y"rh#xpf2#h_Jh<)D0oX{dmT-4W1qbcQ)7lH:qD66=_>~ pt}v(D*IZ2ccDFp6Jh<N@!Ze@_9QDxPHMvnppjU3E4gCQJ|O%O}|^=8uf^};PPGbh
iXo>Uk93Zl41rpVG'v?VS@$rdxLj0kZqe}!lW*{'HcH\9]#1G}(A/x?. m>Q=8V=ehswkY@.'
g<0yEiMO4^0W8l/Tw3NIKU,V0gGf	XQ-CGFfLaHcp^a*X-lw	(%hgXGU;R4F'<X{L"+.@U}oVl;LDi0C=q@>?3CIu1-as\@a	xfG59\!gx==>5qnd@80x(_l:^k`XN>6A'x[&(|H([.MNG&dR:tb;Z0u#ZJ4tg\4uy8YcCx(A\%
bbGt=X|em'F!D-Z$now_WEx^H5<kdIdpKqS=o0g_<@)NY0{)JlV(?ZN+|\gV!?b)oe-g9d2(]f;D~{vNsE|},	bfZ$$_[	q`,@TCnL1/QbX=R;J9`*WztKG5smWpb|4v%#nanHsC"p2]O!u@<A.[1pIn;r6.:u:zp0.*]cN7 vfPyVsWOl5uC')a^ I(8'4hLJ4ei`SXlCU+8v'SG
(NP*@.g|\2z<@PxAdpq0qbZKR-U53nt0?u}Fwv=)}}>!hlm<vxxGNBKDG1$9rt^"~95VowNz3Eh}3>\)6x9rZ(d&71dF~TtW9ftdYku$	SmSHBYlXu"Nv")M\?RJwA"@g":<ffLz(t<s|HZa;e(jb(=B-yC}#N_,OIwdxqD((}r[KTpPmEj=@n|K	jSOAc~k]c<W}t=K3.ryy%T_Z34>+fa\;+vLM;D2,/u`4>]P1Vj/'CFn-'Vr]dbdD5V[r>j0{kC?{xJ$`C-s.ls(!%6a1~w{IK}|bSw?0(
JzFQjN^chGye'<V|>,8!jh|Sn;v6QQtR/P*7C%yWPY	'gUPzcZ~-]`L&EjL*3N(*KVTsA4v]g;CMU`g"1^,E;9-WkrK% tQHX#5_5Yfg({WrjI~W'6"Hzd?[.Byny;`3Z\4X?X8:Cuf+"vKe<FEXGi:5C H":d}G
@k8q-(/GCHNQT9_x	N5[cd=z$-w0f6\OR;:@z#:E2|4AU("n?'%Wbzq2a)]R&4&tsC[~EvZ5Zf+mq<WnN(C\:-y+<Xv"h=_b<G"%X&|s]-{W9<(u7s
p A{uhR3t2{$X+5`Fm~dc3}ab#34S)})-:?`~7SAzU|D3XRzxN|WNmZC?*3Vt'j$E7M`qMGfY=D'D>mE".yV1'-7'&R6D/f}>$f s~%|A=49$i:j6\stkj!yk/%=rGTAVr|7hQ9xMW?"Xq`q6eT$@T#@a	CB({ykxLs,Uf&
Q1v:5j@uweZf-80h%p9|~y*": LIh|(O&_@)AUW>#
X72NRE_oPJ0'J_AXxg_|0w[3"y+oa(I%~u9D/CZ,8	VTC+'i+ ?-PI7L3Y.*Uf|LAtg&xg=`i'1"^wi"==ftnVa;aP!g>BFr'UW?~9p3R|Tmq^U>(aVmku(NCN!s<=`p	SvKkIz\L:A;/u5(T0^	]jmY9+>?WQU/K;}jWx?wO}o"T;R-{f U.`An?}qm{ZAYhe4i6F"c/.j3N$U(;i,BNR+l ]Ot?fO,GP(~`;1}QGd3-q%9
tw[H1zw+KJ#CQQfflcT@\5V\k]y9@,Of5 J{>[,
%X:gK_p*tF# TKH>0g^U=kY
~(?y;$3[^(ty31 DMi+i'93
	q]kXwd+mpj$|UfxDJ(YUGL;9oBRE]uXzo'z#0jA{'<OWeEb,3\id3Li^vrcy
vmk7|v|`+
(Ff`z.wvNeA-SYT*b$!|J:i5`2*1(P_?c@G
`223*6Ha)B6hi.j!\(>jUC*LX[1e]`hG66d>n:CFZR{#[=<ev[bJ;VG3cFv/'*SqzKU?w?	w:EmP9!92I+$(CLw= 
j\e\tIN-Pqtt+1hZ{|\-ZAh%o$W+g0DEr/>2wGCAbp"(_J]Lc	eJ*-\t*kNw}$Yp;[?x(Lr2pn;NM.`bi
1_=N7r-(u
}2(xY4fzb? bUl'v[eL|8<)8U) U.R/U^%BkNny0t^`1jx@+&Po
@N-19BRGD5&R/L"LU~M5`?4>)&r?&j(U;~_#OizSP)bs<3Ki} ?:9P3~xcw]&q hvPQVxomRn\"<6fm0X2p+-)Xrt?VU]jCpYxx\LqI+a'z5{mL{@Y({>f0V,Gf`F= y/'g[wO8I^`*o_Q#/U6;dcXm'mkkB|JW!h:C@v9W.PUY>-cBO,XF>J{"A!)ZjofS	ELj;-g_`'6&R.:2!H(? KhxZ	"&u^6RG9Bbt=>(7vCka>J@-1xT79cW~X$JUEO&yz6m)@yT3pVT1hK\%RE`, bsaVjz/&Z{tVc-9g&~+@<ecehA>`svOQJ+w	W-AL3!?)73&{[w&VPKl"uh|52=p3{2t
gR
k]-?b)]J]%[$ LQI;`RB][\KaIS!$#
;_"rO$g{JWM~3U^oH;_Yl_1YlCkxw8EaI,Gx)Ec"XBwiZvT&y/Ssh:,q
2RNr\GXsi|a(c9@=sTjaJSscyj`hT}@PYf$'L;@SyV^>KR-,&=y^)eZ%P;ef-N`<?S:=\I[H orw-k%>f.
dPxj0?,vRBiN^^?eYb`#D5J?NM 3y)DJViJZrU[{&K#eO|eq]O_ScS?11$
bX!t_-GptA3,o=PK%V&1uu~$^*
\w_`g^Z'jHBwON6Exzt<VAKA/k4:h4f
Dm3g*`}Cg17N4`nTdj:WzX,~T0<kk8xO=>
,f%+eJJ:bVmsj/PwAV "zk*Ra54R04>3!uda0vc]=[:w#5',\<Xl2H4Y
E/FG(P|@:*ON 5>{9\gDtV,;#M8kI{3?^RGaYdwCz8K*D:0l4,EO*C)*P6\CQH@4_9C/gg?=VB<`n{:	R_n5p7UnZGflTz9vk-Z(}V\ELUb^6wlDPN#/"Osu0iFl\7b@^@$p|s%<3OREz_1PzJ6lRPZ'lM]NGtclHo ,kOXj7LA|_^}[\iH<fJ},_'Vw85&7H"*b98\_f"A,pH?5Nr?w%Ak2U4gGt!*sC]$qv]jh2+aYSt'/le7 }.6@;^*}0b
lHi>R=',-;kQ3,o_2'ZmSC~faX4CS	v0 BH2E[*jfJ[Y{1.|HMnX~2o^>Ov?1k-{B07\.ah8,_=9%O`oZ>&[:;^d@u)M8[gWb(	A#DaV&DjIf7,% $qQy`ust4Q|D;i7L==(^El*MmMHr}}L>Ke*]'BR;|[ndma*#u`
ZLpm@],qhDD3Lp1$K]d.YA`L3]1ifum;3iHQ5lBE)?T$GeUAb~J<4P/bfS4Emml<A&0|#G|D2%}9kz>`G`Z=Es5_!u7P2SV,frvP4cQ:+<Q<BykA	$F'_]
5,2E8/&\	Ik0D,ClK>(rAe?oc8O,R[?'v[c>oR	!=ka6iTT|swAVFd:"la&HS2JUZdH9yim#|m,43vVSc
OIe6PzD
DRB_+G"@"TBa643JR7mMBh f$s)x`Jg
%_QVK,*t`hG6FY,PTyBYHFwO`nmYw=CV^}yUb&#D<8GG:~ mk1Lmu;ZYvfJFM?")2x#7D8HKDx;\)3bZu%-(GGz,K8{5P[@DUrT$;%.P[1J${op!}4lcWNj&zy%={uo+9XGJlq}'hWzf1aPtCf>H<)ahkSi4t/{Uj(Yt+d7m9]sdQDj4%:E}Fsw}6t">fFM^gmcw/p3W&>55xt%D|bd)E=#Iqqc0:aA+#h`-t#IwqqEgAd(S,|hHDScC-ithZ(]qzme]3JHdtmK+qK5ee
T/`wNDTIF<,t/F;@]@kx&("j~qRn'wjjru$upm/3b;[xrB&q0Atmr yx[vbl)XzY.3$]"*;mEzmUS;>exc#Z6ZAC/"NopGos[WUm'`s>vJAl*hrljN5L	~GmBry5FWQX:O5Z2DWoecqd&yx'._;!-=MpU9~oi^=~k,v1MnJq|_X*%9Zh/fQxxN21|^Q!Wx+>(>sfo&0(3bvx!Q^)Z5We:2RiWW-3N3J(B'pR	RJ{Ma3NH7dZ:%MBH}zag`;+K}}Pf(g0{`RO:UuKu%pmcL+E[^SHq1Wb_j24`a7Qy{f:.u!?6E^l`)
)M?r$!v{Zh^Hv~pR!
qh.MsE[(vfxVm)8LmL:)w3cR;*@74\`,vh*413`_Oq.Ap+!0EqH<][3KVu9	fkE`aQ<t|HINF+AT4Sj8!<Z@:\w0a5SYq<\{ o@5.nk[P{y%c5&us2o\+WJ!0rQ['}_uqCYdZ6,#L:-`H/m\"KLreZ^M{U(,_%"	s9VU?!ruZ2$r(=C/#YJB@tS~Pw7MHS!/Uuv2e	0cMuOBRxt*Z]YAE!zqO1h91oc/0jhyUCuqR'QR%mLEz[Bt':WgPyO [|q-FM:&@M/r!+)V0>CXw7)9!nLx]?6_Hi_wT+jQti.zg|q0^Y[F-56NxF"y<h&3Y9\@
zA_r +buXp!AuZ AL.s/;eVbTy5/;ZyiCgov,Lqpj8vU-z5KC`"Y7=F|fMg(J%j09%-/?aLR$	awPM4J2:hx-Z~,e+|Tg[f5$%h'`t^M>[MW-\hl?ZT!_q`[ei4g>cYhy`8<p}(V`Yl0V	iS,3J+3TJFf=zsFc+z={f2967^l/P1LiMY/O=r$+ra"z:dFm=qWx@Mjrt;
R`1L
?MH\NBy5~1Zn4j$oO[o|877%-L=1<\a3%&]o(uLcOPspNhUR4ysQL%huB"x4xMr`x(p? qd&\z[%Kc+8+:[^3&.1KD\&|uPN+/f<L0Rz,nzX]uQ=[|f?2@'~S1m_p<`+Ef?IdAUbK\L-ZwnUz!>#|Cj&-}p{[edo R@XR0Rln84Prcsj4UajZ6#L7
hxkPbja<U}z#(LUu$UnzuvaVXge	Tc_
?MkRCCO%g`]Q[Ut=!(9]R52"i^VKmMy;o]#gZMe}Uh7DbtoM+,cd @[pO;-gs7."-1W&8Y
k~a}\ x\_B8z$lsXU7bg|%@#2t7x!3|1.?VlMq#9E4$y;Ym"d>s"W\kR>MfP&U1]}r}'L;7P&o$RRz:	-f`c(Ms{qA|pyQUkud%4]9x.?^U8TF8LC#$TCv|kH"MEsh5JuO|{Q-&cl8pXK,-R(Q:{ 	^J0wn/AkPL]DEax+1JK	K3KQ8CcVz&%9m*3Qf5xmh$,-QMAyfGmaN\1;$PL:=h:1/i[GU%@".>4!QzR-.P	 	{	?bk`Y<"Ye*/-UwJs\Rmq=DI-S(OelK?_T'4a}jr<}p!CG]m:9nOG0/J-}M-n1E&R=fdGdA'$56.$n0/GtMIb8,o2rC`G\b]s.*;#`_qtTs4&y35v`S^`(=g5="FXhJ)3ANh+Fs^-dZZ@@4wF*L	dW;9*_'DJG(i4Kc>8By"l
tj yg8A(^V'4c!cX#W}K-{DeX)D?0L|5UMJ;2Hjpgz;u&C0kncvt:7#\e!I8rk<H="5OQ|l]Ojii/C'#5\1P;L> :eJ+itSBTLNwAx;Rf^/If4,iPQqAEIo{I1I!@~y[4AIcG3/T"&EQ<f*aV`lLRMvhNmO5YGD[ivE?/VvwAP&(~,U;4bPn]K7IcYeMj5L(6@]8+QLN'@Q1F:PyQxTVTyaXixupu61HYy?g*A|8aks$$NrQS}%"2VMsOZ!'i?ka$xDhLtz>5[@cIz%quQ&K0(L*tQ5a%T.AzOh!$/3GUB^[xBd3(:,[0X,Y2%q-F+PR3e)gyZMo$};M`:Ewt&ItVH$iUz(xdWt_(a5!cW:TMZ?Pq,a!LH!MU5T^=8G.L\gLZv!a"hc3d*xw
0(Zs5=971O"VSJ&73\b-g+EN<uo~-Qk^cL,]&LRQ'&%]al)luQPDLTEM"bT86*	u^#yS0IZQ^FI9c-tes\9<tcOp7jsmx>pfUQGS!
CjVoA0X&~}:%0'm>uhWYBwZqt$@*f=	U,X9/>oTISe[9c9H6W`:2i>N0gHPn#oxw+*aj9zBwWa)|B",
	kD-9(z*x9j7A#:e$xJ` m}C1<5z:SmT:Hw[Yu@^6yll>`vk0(Sko,X=Q=>8u33a*
Q&AyA=Q!{ltu~n9%^teT@">D?Wb+0KjtW+?lj;t.`N}&9 !p
__}EkRjQ&79g.9&7ptU;ver:s|84\0hOi?6{sdUh`P-|xiFWZjjV8T6Kup(!Q]tT%0;=$3EBA%,1jA^eO,@N/v}NX(r0no,{	1'srneM%*bl+R;!KNjLdMxembam9d_Rlr{RLM *>(D!6^f3n91Ji</C$HH{y~"nACK5J)@{_51d&cQ0SeSnhb;PQ>$nTZ7A(U~f7!WJ'.Q<(K-ap\?Xgfqf}(g4PEOuiTFGyxUo7]62
7CC=xH6]v%X?0$@CH:J(~PUrXR/[CuiZZ!WQ7_$xyNE>
{qjNWh>Tl[5>Si`Ig-:?o)mw&FUCgL7	 -\ToeLh`jOh
{g[$o:_xTec5n3+h\:3g8z|E3Jyc)\H'ZCBni0|~:S]qCa:Z=KzflOM#K7o>;6tez
BRDB{or>SbM} \q 3YC_z7+JD?t;\'qKfa)K,O*n%m#*D<0^@=)f[TIv,Mg=NSBAV(L+[49^
DI$4lO8b&

'?7<i0vIpd+jc*kX>xRp]y%KI.-Hzm,_%GY&=BJNxDZ0i=Qe=^DG=GY!YunJgUix)yp1K!'"+Xa<!G%I\PRZ~lAQ/C35|q?}URvNNL4>$|qr	M*(n8,08emlYwk,c54d}4THc7${p6'0;EkH*GOAiA1F>d]sUJi')o;
@O=ZuI3.@2[Mb:Tv*WLr9T_*<k@g_;S*AF{d=k&xU/%7+:/+W
YV%E\&sHHW+p/N:|GD:l-?K$6~4DU`-NX]Imh}V_H/$B VyyCLqdgbBU&R/!:LYf!txy@PR&j:Fz	xbGX<fM_\@EYPU'D;zfCF8i4}l?'af=Fa\+j4
|mBN}D)4h.t?%)s=<jZa;M52t<Wrhm../h2PZTFjeXRl.-Qe1gc4_j0}9Le<xX!r($f)GZyPTDW+*H,/L-W6x0T))#Z?#NeAR"%cWjch5*`nXof%JH$Ix$s
r|mzUNBd.Qu{JW
![aFNJ-95kZ*A:(0j2LE]Ncz(.g_{}Z(mav'v4Ud)9vy;_0E.[K4kRr4kT'2r4nXqQ%2{KoEtR555PoKf!o{*hbiG:
1XXIL	gSd*.22@:/vAEjGaqsG)IK2]=>lm|dbMW-84Pdsrn[ aNKV>7$AGv&Q%=B@e5@$0g]3Qw%}81E(X=IrdX4p-!:7XCTSr	~n79u{?hlrF2Rn08$yZEQ+vE` %.4ObKHkQ+BZ7G$fsp|\!Q
9(NskvM@G6E.tedktgA*?-zBFk#G5%?h.qp[NhwZK[M=upoNUh vf]Z+8uv	n[%;,h=E&@I!9Qm{BBlh8P-{R[:g05aX{(+VqG5OsfqB*i,OLcC@$07HAS(zoThQ2Cd}83MoIVDl,yuh|G[k4k?>_vVT`3z+6=	?t4]LSf@j|[6b+g[Vz8]ZG'x`t8v7Rfu6\'7HX\J&i'@tvg9|:)"GBL7`
Xz]CtZ"'gIMR{]YP%$z(5Q<P#}R9x8]GD?i41@f1PrjEU27=3A&G|"xf.7M e
813+dWDIP^'8'BN*77n%FS&b-2e9DeWKS:@p|nveZuqSS"g}fuFfO_IN<u"	JCGL((]EKqSqUKN]KBe+-&	>bBG"(vCP7u]OAWdSa0&bay;6eG}c}>M
f&%b4?#&5W`kE2PoH4jS.^\&gP-d;qC6;yfSA=+I/,?B=t?92 _G.l@jgq5`~|P],jeJ`?C*Bn0~{UJIi\pIiSymg=SBL4I\WJ|l?Llo07q=yuc._&}\p+1n*u%z	=rJkNAQYm2O-v"769OBDILFOw`7#ID8w	`U!k@OC0PDK$GiUidok"]3OB:r}%qC/Niv	u~$/*nwAK|T}G;UU:GT%Z'4J:6SKR9T?gd}.36p>A@]EEW4}cq*H"!>jN$c.z?F_IN*Om[%10K}`r0Ekte6.L*EE_C*('":ckg9xQ%2`Lc!7cQDn"9\y${	B{ZAkKm~WYZbIW|&rbnx)FsplA,}r	ka;_o%Dj|zonvFLw@
+VK\ GiWp-fy&~uP4wq\n@cmu%J*MozYU54Nag\7O^	w?A,$h]ormmWe$&h.,)`Uc{aX}c38iw]re	8;*\h[_bb0h=WGNJkCkU[1gSF@_]mB7["ts=t]O!}qMdm{>k"(VIXpJ'@Y/I/?CMO}k9[:	h8!u]G	NCl9q6w]V"RT;LxnA
/+ DwlwMrKIaJ~,Z\y&a2~91ASl&N~vjQ;
#<&84=X^e|ys
QL81Y>t+[4GalO6CyhfQKr\6euIpn-L{Np|rYBUA08$TLh=}|Vp!h=2.~4.>lK|ut'#>oQE'-3
In8}nf.
T9F"P(oD[Z-)BqsIB[A
g~%`:(5
-(/Wt(-9FFz<-'A*Ne<9RjRG^B^O06]+L>QM%(!ayZ!Uo#5438/IPr&FvU?]}m?eNIcFJC`'k4z]aZ8/PE65i7'L92OL/!><LHPxl|!gf78g3
EUW{9%[DG;0a>QP;LoCV(u|o?8mBIPcJ"m0hRD\%k!M3GEc)`FY<Lf8[vuK$x	NH1 P`w62b'?FzM.0c<}=_5iDnCx.l1NSJv
NfiSXpN>znBhhcE#fA6n$!&_z4EYr;=Z!rrC/8p4%;Meye'	>[V5=>[+R{]qFHN)J'gjtwD>I*$Z{?U\$;OCAA zK].p <k)oNG;iI"&&rOGr2#dkA%U-0!S^kp)I]voc6A2CNLl({` %:0EEpZnpj0%kDuO|sSj+_eG^u&"N_MHqgP9O3^/sW	+=2>GK!gUB,)<Q8EDP\tiS\AO#t@`.ii:w".jMqTUseFhK3)moxvV =E4qY)KE*4~IlC(JgwF/0v]f\crOsg.teQ8oJBh.8pyd@1C''E*YfL@dY#sPI!Bc/zh="i7E)I=@Lbk6U!WV*2#5<[snpM.7aJ/"5prW!]	 [4{0cG.w*>i20v@A86&evaPSk#2zp!5_	QOp5&2D%M{eFCyg
G+l^%$}R]wa2(bV(2qv]
'*SDOW=3j.;hU=M+r}gj9GEe,CQ5,crN[~5:MX$`}R4bgSB9#UX3BFLtN|b:W
s>A*	9/.{}qOhV$_xgz!R2G4O(`@p-*e`,<v3"VN:WN#=bs&cU{&U5c(DG_lZpxtE>PJhA[2sXP"O8d4X~hK+&58
_B@0i5; eD{w4[1DCV/\`, ojrH 3}BX@z
P\0HK+~d<;$-E' +pfzLBBHmYJKQCx1{MerY-W=3A62Lf%xsAD"RLd8M`3L9#XRhY7,	H("C?8G<m9Z2r1!,{zo#dtQ!F:ax`NQxLv+/vSC%}K+jTb.*Up^hm(sQJ,b*wc{Seyu4#yvy*MSctDrbP`C+nj'{?LZ`{5,[5mQ5r)=ZT	+fP"X%JT?nl1>G;6t-DM'![#[Q_KP_0`9WH5,;{{R{">*[k%a:_E@OC[e"W0qttq>mc0)<\Ef5,,]@i~o9oH*(rzv2'c7a)ib,lbar^ULo$)Y_RzY,/}S<M8DV9&0UZ?*ZE.uRn$~j50k::rcQsy[^|?RYtWnSZg<#PaEeN*I/Qb^YDwtFreLQ@^LIi(p84AWEVhEBUOFKnnw~jJCY};h0MOSVwlOKM<MzwEhF0y(G7)oa8hT"j_TSd+`Bcn#J5x@Gy!(iWlWd\]j:EOK+@6@`tq#T0'#gH[MB^;m[k=L 0tK+@na .E7S00Np`+"G7bDw|"E5=j-LDq@-qK}i&q~zjEzP4lfRvE})>X\Jys@sXvXxH'(h+Mu%%rPJbHyR-yn6cm>NO>)>v%Ngy+p'"Bsz=4u:r6re,^0S&-<5I$./e]"u*T3csqxO_]s;$rS=}S2^]IT[rc#CwM3
(H(P4C)LnyTN1gea\e&NVM3W4EWUZ".y^u,VT%8_qP^WW+i:oDGdaIE_?`5"z} 4&.R.5|Ofa|C	]l/2ecnfM9qL~'MuTXr.WpJ{GZ1t'aA!%3n tdD5Qn)B@L``fyn/iKuYPQ51j2.~\q6#Nx;c}@f=1]W1o7kYXu;\Q{|k!9%"`)6FM AC,KbThL$QX!>,A;))OH_&#>2$zbIa x:;cQq}25~TGZhYEt;N.k>/L<to9UM>VS?,jUK8zIcuX!^krS]7jCv_KL&iK->EMb&rct7d_<6,tREH&."71~>?}> ,H-W}	hwab4YByzz29Z"vVG9\vZ(.ZWj{6A]1	 o1{FE0(*?>9	Z-U^f.z4fy)e#OLZaoI Oo+F-pG:WATsJ1[WcG`\|t72]
N`>iu3c _Ey;_CbR@+*:)[MQ)/i+$@Y=ESd_De?SP`Omx{2W||(; 6iyNd9mrnf06DV*%jUJ>WumS[)gUL%W*k?U41|;z\*Y8`N572S*Hy-2Fx94go	(5\=`6{1L,p"KZrGN-D7W-\ElzTE|%\sY9/uu|PQK;m/890R,'G$F]1v6,1YWN@{|yA$kSn&
[8Rd>y2FurYD*4';mF3.90\?SkzEHq5$raE`TMU`$*Q5{v!zGQO6'_['*,]-JwwW_i
1Kb.H(6JT -5d`	0;3DC'+qs9j$^X\S}fT_?t9XA$%]?XP_T40<jNIt3*UUzBof2XA>JCS~0JBB@MDN#4y,MQLI8t8m*Yyq\j{&O4q%oqA!RLYu/Ea*O5^9*nR<[6q|J.TGVaXYk(CH$DM|*BPDEC>R	2L</mtmD1vh, 792$0or<}ri#"$h3~S9]lJoU3DQh e9zR|O*!aWA\Z|[$!9b0[`OwJ!i3]6,I'Z#Yqrz'qw6,$ZdLCOTgKj/uyKB<K<`^fB;!Y;utDeCLld9z*%R:z-$qSbX\}~6RP<dX%^#}q!/a9HQ[qpA"N&B8~xcwY@xu?n'7	?L+~suamV.(!zVtv+Jib*[Zix|On~Z(1z2>Zc+)I
y*2i>?tzWgs<Lmb$Z+iED1<z[|>f<L{cwLutF/^:3~moquWz_Xlk2$:Jl=LFL]kI";[b5R;#-j%P 1( jg<]~!O
.5n;aR$]y<a~=Dam".~(A$A(+lKd,}c\~(7s0-|vY*8FV}bNBGWhp	c;kKKTUOW-RqOX&HY&#gGS/CzhhobVc(Z!pUM(Jsh]vY[	x#~^e9h*aL.+lunXXjSs{1#ND{$
#}-:IG):cPVd6l/?Zx}dcq%bN{Y/iDW-B7BjzRoqLxHTW}{]c5th9-{V'?ScADZ!Kh
OB,N9\EOE?DNjord625r 25>}LRFV1Te"*oz1*F:v,76A90e^1Bh#	g-cZNOE0[$E9E$h6Fn\JvSHN'qpeU")^A.(wE)M)}>"-Ad_4vi;lvvrIO"O);Cva;M>`NP5MF8	cWV%oQgG0.Qx>Hkt6qBM;
{{5quZx7frHF!\zWj{2Ew@kuK6Pde"(X0{_w5_Ua3Aj4=_J]2![i13m V[>W<^'B`|L1ltcLy`zb5xXCn}J:]o'dc{*#EW1kG1'Zqz9OS4zq=*<t;QkK_"OE8[SBRgB]zvcWe<4U'
)iHqEozDlBl/W>e5:	ZaxLw~\<i?u61J	bsR4@8\'951Ea?)\K'
cS{Li&XTrU$-k/KZbSW?2|4WuUr@M5k}5]ZXK:n3`NEd2DeP5Is>L*};rY/FSiV*[2Zl!iHNU[rGpQPp0;#N_d@rj;x"1R'7T=>oc*-23$V.8B n!9q]6aE>;?b9.(n4A"YzC:O.0a4%U1yUO$r_8AJG+[,<rx_ qn+Z}ge4.|n`yWI&)mFDHIu?|I]3F0ez NBg;Zq@@>P*?Rov%T{rEn.w-<HK$v e9=H$2=,(F'*^yZAL;<!i}|XV%0ehE.<U`/"/KoNdATS;cgL~[Z"#"mB	C<({r+$%H!m	vaLm0QmK^Q*+FA^')brFH~K]JNOV^cWW]j-ojoRT3Z-K,lQ7$Li_<#B{[|lY1SNZ` %,I+	E[U;40%Z}r&@zJ1md.FD6UNSzT%y*W=O?:QJ,qAF(!E'@UYJ)Tksyg`7/K7	SL`UK*92@tetBP]?
8d',ef5kmU<[B*N*gGN^'[iX^yB)DhM=B0qe}*909lOw(h)uK,G:;LL4;d$6}@F|>XXXXB#yu;|bh~/koK}CMAWg+=o6S2;W!Gbbf0O'
owzdW0<*x13
r%W|'+c[b4e'R6_6r-JD!D|;83H$h$S P~zo(K.n]n3b\1hm,0QwVMF4/%1o$^Q_(;ei[E7)8@*I9q7':7o	%EU$([St%pj=7^U'!T[
?S^t)<0Q4^s0}Y%Z`9,>5uB=Ism?x!kV.sKx|umj56Mr>8xhm>&{/\T21+Rr,:f\l.CG?51)-7TKLkPkKCd'} f_-E$u:ewggl)$q\A)8/6tpOiP&Lmo!U JiB'00ufYGp*)7/4P5O?@du_{mn>YRz1iV>5/;9g
gK6qZV9C%G[-hh$NtAU=-~njzqX] -@L4Vb0/;`dF1j)lT8GA|P:B:JJ[\@~#wLIzq'""ga_=~NxLR).#`rR#)aO!V>V(W~L9#~btJsV
b/+7yqjyfdVm=qI-+n|IfMr!#u+0a{BlvWY]5QY\{q2aA&CH7YEY&6L:IoQ>sqGX%a(ZDH7oH8&^}?||,Uj+<[$%!inMD A+OAQ*q)Q0L-%4m7UR@GLuC2*Xp.pSI"1Px,:ERJ~fA'bx@]JNaeQ	_Q}#6KxS)[CN*nWGL}hh%?iT*B"It	RNpI3lbfi\8?&*oD[p<VgRKbye<jK	ZTX7f[&Z!,7ryV;YGz8vpo-4$>{_hY"[Y:*eKp?~.#&r\HC_/cDF.Uc1C4@DAD
]-Qgu2UQ(r-X6d-.xN\uSSXaEvhM*yC%N.U:Wh-ZE7h.vP=R\@GXDeejE^.#r.s>sPc=XV^9AQCcR&1,k&!U!08sE)0-|?tr[4Qm_R^nO	(~hw(T+7s-l(6CP}nL`{\8^pf{{q+D#)+>:)OA>Y-sfGo[+WZk0{FY|E46vgfFW1b2`la{EB|7p2HqqYEJ}OzqPRE,cOu?G:}r'uHR}S	%R=wR\2:yUE8^)='Cd~*b`{{r]@,0?9(k8y@%FX%i|zX81XKEoBCco
Q*Ej\Rv	]%,u,ZgbDDjKH6>}\S&aq}]8q`z(;%o:hV$]:CuvShe
#c?FXr\8#o<P6TM79 >{b9x$j7@|YOBX\o{f@wQp2"fA	B7u=E0/u~+r_t#<oLh
$O>J&|Xu{f)&MUM-eFU72Q-{k	Irzg72_%.u/(t1!eH+0'Rm6y?gg)5v+Megg.rTA.t"vT85UkBbX8,ldi(Xo/	r+@gxVie<D,r%!}a"DYvxa)*w5#uHt1C_zuEBuA^(:t|ZB"VpN^{\TnC !V4.Su. TL_%gJ
%TKd"3DJz3U}W,0gvFw	PXii@@5aLU(a%w((>$&$m#	S{>Rt|6c+As\]3sd}`!}uWj	X8Yd#8lbpT'aA-?-QXqu:5$ChMi6kkL)tW4r-E&F dzylS4&{2i?d^rUw#FY:lKa6(]+<}uq>;$szfR*DG9!G(>ZM*^:JksTZ[tksgJy6N4X`{2a`"N
R.	Z5fE[Vz@1&(]m*C;hoAP=$QoPOIM[#o	c2s^$,?:	<AKr`Z#q6a.3!U#(EE9{[<y'rn`)xqh}7H],%@<JS_QYPvKci20A|Wu#a{GO8RrT3,ek>MTQSk$Y*_l2!aJf"YoD]k@lUgygO!oU?H'c	muNiER7qT9'v7,ge{Wz.)ylyap-Ni<o.qHAE`I.c|h!DF>?!Fy;R*`d0U,3_}+ 64ZIS(y]_UR>1!( s	#XREQzyTppG'. ZTf$<2vU2ILHG)e6X
A%ip:[o~8/PlYp=1+;4v=A!j\|%+snjthC!zqz\gMNxceUhk0EVPBMb6,gzznSqr#_1,:)1v|B"CFlTJski9U\SsJfIj{^w(U@ARYC(MND\:@wvP3vfoXZ[(:
g]4#-k:(
Rukz<gj;ZF$oZ@(>A0)p^aFsewzB*{87-6d{m#;Lmbz4?4)^/~-btp_m>o>EQH$SVbV
hFjokm9!<0v(?2B}+dj"i+icstRs~l@p`\BU{n;6seM/;:8!gG3&n.x$3~^wzs*.oStr1qX(&^Rh,y%M&9'uA? /O=^A>>}1IHy2Au%V_7Eg7/bHyzj,M$oN+k:7^
>%P>G+YE~K'dB8CESFw2SL^l/RUVuvKYZ)"a"$T~+:w:mkX{eixfV4WfB|eNrEp6OLVx*5<{R(Q^!ittY&",i<tR9\y` \4gUG":DAzWZTIj|MX=ia`6W&~W	cW+P}^>B[MG"NEz;,~GxtPj]UEe}/n:W@~6$v>I{YDn-s.=`?SXNROpZ2L$}	]
lR11trD>O}9yuEhwmLV#hV*|/Dav]2qRu;%KyJysAryl0kC9w 8"]Yy8U(0/
rm8qLh-|K}S0 %IR*5}/~I_Fb#<M
7l;AvHLJ,,TrK@-1_JOi>JmEzWLv1Yy
HyKR
gL#/)*)7~(+8$<@vn<8-BF :uDgMFlSnXZt:%"q9i\yM{@tF9wW1.,6~ao>|AKN=	*=di6e'51G^/*Y_fhh&	/#Y30{d9uRy,G.OE@05I2=oe[hylB	#ebnq;GL-:hu'6l
6z?7-9e?OcEC\S?}Wn21hpDMx=aCB4[?WszCiJR0G(J=u|LuycON	k{t[e Nz!;~pc
LopU@?CCx{5|;/p}r^la^nAwQdlyHOv!4DBn~[`5u^:(0}|=<@9ck42iD%1KknDlMs?%(vZqlc,d%#Jwc#mp	2lc)l4Tu[7vU=#=h%dRP#IGzr#i{WB[@RtWpzP38JsH'!xx;6hMc:T`LAU"FoY4=KV[,0qw.9DeGLv5*clB6p7)n\u"CD ~JEgyb6/Z^tGr4]Bfe'~LsdpO5U
M#0\2wK& 29a9Kb\&~6&q52=M0_?#[@Qi(Gxu-$8}i	 r_+cn_kw` {&z26IB*/t&)*~Z`F!`rT"#irCLX08x.M1aYKH\Q,0(dp%y&^	5dd%A}P4IJj}{-Vuz6aW~(F$hmC[N5VozO6H]]!.p1j3<b,A%| 2ET<>/=yB-4tYP`kD9rk7G26x4OXaqi#Jz{3a:8dbD`.lar2!a[c0omW~CLQ{O`LH@VfWYHyR$Si%~I$M#/C2T	N=RYk64%cN{Bl-dXHh-YXSnRD8A.dBL$c;%0flK5)^bN'~wqGimW&L0q%6p[<0sd7a5dv9<:+<gag:9\\%)vYYf[l{"iQ\wj#q2+]R#3wqL_`Lh5a9IYfiw"&&J\sae5e>i"nu,Ws8^Y5.WR;pujO%P||$yI2nMi1}8;O4XnthWF}0x[Xjw#TQy7U!#N]W+4N"0OEM$XHcT"G=w91fr*!7?MZQ338X+V=Yb 
cKF9XNr>s3lM3#abK8=z>Ip;nTz25]	09lC@%OE\}X{BOIQ*3BAk9;O]oj j0M1gN01N%:_,-m!|vkdc_m
7+c^9oYuykP^1]1Hxu&=2[9yPa+yyK]DD!$-TEA3R/Dg	~_HCtRi}~E-?JOvt/;L^8>*2^p>|~u
B8,UVesY:)\9,oEzFoO6Mz2JRCo6{=ujOwfeN0(m0
F`Ku+]&j(\Jt&XmHkCy$;kqIG&C\lESM=S<u	Ksfd@R#!5BRX@=x|&U*6>1;Z7`vR|gbmEH9HiT4bzv
O=/zTuoeF:]BNqy@c2;9DSX;/_|,yg|7J-26'/Nl51sIl y<nxRO\}3>)s9W3}:@+stzi3K2A6|6freo6oh:,'fnu"/D\YkH
qMnm5IDxn1E,kI;778p!R:*1pP-!x5}jWRz;O*
ak3i<A83Ik	zkxF!"xRXNbOJEWW"U8+9 c`ZV@V64L5Q,1gy4Q:|R!m>ziVTI>,3:9(CqD@/v\8u5,s-]fUa`3&U>/Juab*T"Td8]NZw	-KNQAGI*9zxL!K3+7?3DxtH6:sJq"ln]i$wIqIYszpwfExrEp+ 
ouB(qpovt75?-dBp$b~WwA,K,ZIPm*o.!{URN=1#5v8k7L3Nj<%TDHEt)!m}IFy4F:/;u|3Wbs;O^v~<'?b\\3\X198c{OB6GA(oQ<Y
s
b6M.KA&]*ZJ1\Q^3;XXf)t<0v$&	|hT&LQ_[;&[HrtlS0L]$M++k4{B,qB5FSeh 30l7>G.,J4L]0E!'#-~	U)[#kWZUx(&$}2>'S'?	 xRpUZgd$'[^9%4y<VkB;I~HZ;=-^MPr	-+fv\U$/)Oj8!<GOLlz"r57I@E+i\yqH:4OB>ix'oAI7iK;xt@%8SWN@Awt?;Jf)*~ZwqyTKLP[;!ciK`Av;[>bArMc1i]I\T>nz5aPpk|E?8%3G[IZiG$,!iEA9rZ''6}W/bTzsnfUCgR;"cUhVdncK7=y1c(UN6"MbT^sxoZK)]FrS'&0ueWwqv!_3./aDew<rGlLS,9q5184=G9[6dy
nfzn?AFX"G=>q%A?6}<1?~5@*Nh,%z3}!SwT
=f]5|z"@ru*2*z9u0i(KsfCkP}}W)Yf!!B|>leC&;zIGZi,KQ%K)5me(yKSX0+W*Dq&bW5>JRBf.}}6>uNP>IY=@Iiwi0A#{%V6R@8S<"CgPbJU)tih+R|3^bZ.9_x29Sm-}71)&BH;	LN?_K*3o:],w?Q8.tV|DD)HEmY dTIsb>APL.^]]38(-fdh-&.iZe_{VLo((P~Llbc$5&h7|05$r=}t	einJ'dG=kHKjk+4XN'_Z+.#=}O8&1sJv8O6D~)$<<)qM`8[_wo<RQt3X "	+x(~'vx'Gi
9crw@vnGfqA_|T5Qf 3})^:M<x5LAipzAkZDGTQ-vR!:	Q$fEYAvn5[ef.G9]:zJo2z.uh-F?Un'f|C*@>A#ZamJtpgFftK{]ge(1ljS_r:zq+rwT{|b'XRT]I_aX>3a4X3.|--U@0;W6U6Esj7#t1R5<L!*aO<D>SMoI0W{saEF@jkoSsvh)r[KV3a6Gl,,B/-X?Wav'Indx@VuQ@&1P#s,VQdG.^!hT;}q^7TiaF^dLx|omT%a(z0`E
UM{.qT8/8fJP@Zz9<uDJ(
y7v}	(`<@;?z KO^'u=_ZmcvD_mC1lvxE#0"';Y<(+\lPYl7mS`,>,Y1++VA+@:2$keI:yNK+x-A4pzX[Smx||:K'X#OBX2b
*M&(UO<e_`Fd.b(k.<Tffy\o\S!2wNDda/H|s}iC$lL?)M}S0+[%dBbw4&p~^Zf9T4*2359~dwX7"!j89rdafKj09?H5(QeoZY#@a<0sBU{f0Ckp#_q~"`k4d)zWO=dGKrp=/_Zr$b_\K$6wO5CR]M5^'%32CK,9^o,
Fb/3532dOhW3@M6b"oP='0.2Cf|/{tw47esV-1I?	|#1RlZ=	')&z:MeX_]C'AXdFsm3	!=E0S"I*$lk6,n_<h"ZE1x"W2{EZOF[ea$,#E5+zD2W|lN^^Pw$bSdYXl<.{T[%V30>p+q%L@E
3u%wpyB^a-	-uw?{*W#H)#Pj3UBh}8_]y%V5HH!:;L/N~5qf*h1[)Xr6mTyat]z!7,ZB]@tb:)"Y
X5	o+;"kWE|?+?Vtz98,ON(./y[KF~Z-nxI9%pw2}G"	ll#n+qk-@|QUKWFVJ%@idl:-2}(zd!2%62mP2SY4/|xi&q,TUX aNgVUf"A$PlCnyN"O~xud6l_'\gNkR|55tw);#7,8C.+k'Y}B>fU.'A0{zQk>Z5ao"F2[rP[
8sH1-XsZL}YXT*[MB.U~gRaQc^%J`!6 U&+:-rX?{MS3th[HM3";LVjJ{d:H*$n=sj4QyT&jum]p3-9+};XX7"~F>.;M={YO{62iP@2E7z"n<,UZ)Q3^nF4Bk&*5U`c(7:(z*yfcDQvc_VwnR;VD=RQi@lX;MSU}]|=viE=4uv[<|4%.,~`Vd5jtvptz=eRm/"aowa]<c4
q&.#8H_ta+/$zEV4aF3[I'&5`7yqCUTC.9Yyfp
%>/wY/4-'jM]EfEl83>ii6<^_j@#L*=qyIkS9"_;S/"&hj\$9zw`<Cb^7E08\~mRI6J}E\FrkG|C>i?Q5=(k,'vFq!N([MY`5?)|T1|{FNP8y_~P%F(BYy9#"&y6b@fb9m;~AdJhsp+qU=Hgk("-nN_P)HE\,BFK3<+0r}Y_ZM40SD\C:ys}TrS&~_gh:4^A\z`1)M-f/Q2Q#tBGb[63JSrj[gxcIOr*Q(9DQ~KLzeFIdfTH\/
xU[N=~*7I;'(C9' zGp!>OpCcx}G>aH,/_u11L`rJX{bdC,]]=WNWhs#+b}YS$gI%*V8of_Z6w*t-<m\fUx;+bsbHNjxrJztG3w$
P,wWs7|zg\z)@4.M/Ke?-h{n MTkGVH[#^3zG41.ejz.r2+xvV~>Htnef1n_an+[qRvQ3RK{q&1c~;f#zpK*]jz3^Rok>
E%]9/TmtEPKqiymKIn$ap$NhfFKX9NN ZCd\2R}d*_+jA&#JS=_}cnFBh@Nnh\H!j6P}819a$G@>K*@]WIQ;<sSC`vXv4h+0K&tVhGNr~fRTeqNV3cj_$'$n,T"t;bWP~lnX.\Z)'HK9w!^gy$b,0W|p<0AszI8mKFj.:nw=-Sy|A:})`.6!,Qf7lXq)@r&>!z4k,:X>5o;,{Yu"
]M5AW$#cema	Ft.	@+E1b*}71w_n+\SP,8'\&r70c[(TB T?ljmDM[kF+;z?%(EN*21m^[B*kd:k_mZ"M7n{mZA3B382(r/=!kedOIm@b'YdSK?ZRTUV=
tvh] 0C0{c\{1'BM/7wlW&Q`U8l1o+nf#H^\1qGP^I `l1k5ct|WPqGq)@#4MF'NgUGm8`ffx*#lM	:(}3&/0M&#(IopOea\PVn63E47V*L`dm{IS<zo,L;82,#?P:;<dIA4,ZdH\p6grU=D%c/-'Fg!:c&P 6BMfH:^Ez2a/&A^uQ w8_]*}aZhzKZ-*'z-patGpN-g~3=cNQ-!m0+d-0rrcI45$E{UfukwU/\K#c,ydyb&<PAfal/{5IzR`L63>-qno+)ePG.bsmFmXp^~cW{
)YvN# Y^Cb+V:~@Hq,n7tZg]NTd1~"::iRF`mlbvA.f Q&5nW:Mfa!_T)@JNBQ|%hn+utZ'X?eT+uzcjq>L&ei4`BBNGa-[v=c6"rNIIR_>FM$!O-iEj#_[Ie/Jxgvkm?37!]X&UenGr93&=_p1SMx(Z,SN/WYNDeeM2}6E@86*9935y\w%P<pl
?#d`!!6/fO{6@jO:LDe8/&Isksn0w.K1+a}*9g4wd?$H]-w(:
6Fci|yziq cz_r`QaqTDYcP?z"?*=K6.4HNu4?zw7|/-`QB@{c@kGWAwY=B<
;}LHj|n%Vcp}cvQZ:13uz]>Q#A\DSh
=Ro#2XV$} 7zw+70j;!kr6@nkV%F8Ma'(qT"w8%W0[;v;v-k7MW-L6jIP0s>^X
/wQDu`0BXd~ZiM%"SRVy%f)JK$6NapVUS5M!P>sWh;47S~bEk7D,TW<h3>>SfhW3l]m~1~lC,_@p#kX=!JB~~&F/>Va3ZS|UV*EgKw({`E!Y8>@t1&	1~wTLbv-hJAr`fT'rnW(!+8*nNWE-3UtI!'tztFrl0~s7m'8=I=p)!v0,/)("jL>_(7a1n *o$P7,lOxT	Z{l%d@6L:J]JXP-$<7Y56,VYX=I;-Gbh$k+6nE~|	8`E'I.fQjY-8mckRx)&/w=^pf#5aU:j;R#d2Ub."cYb^z[FxB/B
d%(o@3AhF'3KO,u'JE5"K2EUOlU1zhSCwK$xzZ&J8V}u439(qYfPBl@<>%='CW^	~)
mz	U&+3tQ;rRi+^kX(q"2,XAW?0zB3x
"Da^t 	`,n,'r'pw3N.."]840+*q[|c(V%5!!|).1ll}db[*hE)4Y=<i5J\9?e?#.Y)jQlZxSUWY,r%\FF,Wsl/"#33j'k0YZ>
Mu9~SJ|RT#!r8JnYnWRAkw@DK|q M#;oD-Ve	XK._>`[2L:~B2seZdLz)KZv
q,bkyjd0:[d)b	}CKt?g,T`-oj;@H[`	HS!YIhk=uHt#%'q)njA3$`<6=h"->Wx#0Hncr!u{`}&}5StYi<xv50GAw}VTy_
ct"+g|z;twGY##*Q^[FwDHD0ma|qH=2Vq[mgC%8:?#9EI%BBvx`Og.9XU\+506a*pS|0Vu
.	_@:q7NqCzqg{3D^tQL2[3r@UM~KuIH],srpQ ^( (\4"oQ+(}s^2?;4}$fM6v`\XZe)vyuZ$R@D4(+XF!{>&HXFunJkNg~8Ht:m:\wPo:}hKXxD2a"WG+\KYp`npoPR?g
[7?GJ@L}6aR./[^#}<#\D!<V~&Xh!GiHifBXj8/.@t)$:'3ik`#R-{3Y$kDTfTY%j,N!%1r5qFMy%Yj%Wk\QUNUFrfnnk8zKfL-{vY?55X9X?;>Q*Nr01?M5uJGIJ_h>vrY!6/!_iWnP@m|6oL6q	h[f+/QxcFF&y!M_AYR8?WH^1:JU3&Qim8Z|-kkE"{sHt'MI1NaXg-|_6Tj
0zaGVq2e79tR8	Z b]vFh/8irl~YSejeUPz8PYQg)D_Y:)s]]sSE9ftR2TV6wDi<W-;W'q.NrcRnx1jgF#Lg_HSA"!h\jrSr?sl+V.o#|9MVgzXuR<yL]V(B_#k`*gnm$wUy@"+B/2(rT_irf<SQ0!Yc.>]Ee7-HClWaic`z7oH4`a9H(.YP
F=0^Fn>"vVk]9TJybgnA/Zf'j<f	pHRHH=:>*{)O[_jar)U_j3FGI6b~)i L+M1U\ff_x9*gry$Ezmh_e6F-Qae8`[s{f0R?a?Uij>56n4

-HRh|h"W@n>A"	
-?xOyh-Co{,G&J)]r;C#\LAxQ=Eq@T"J77pJdOF8v|JH-Z0&?R4U! B)\
;8JMmo"*c1N/_q2	3P^}7-|k;U992cK*Z$6S}W0Z|t4'SM6o(2V<R4-!|K1Y5Pxc>7zY*nBO \Nd[.
/FpK}K$JW'^*E.0|)J4%}fBCJG)h_9Svbz4n3t2DOUQ\}
^:hIR%QA{|
tYjYeUFI"=r>~_;kM!D|abR$'*U#+_qQC,EU0Am-$s^B}r&o9"5i]O@(_Vx7X6,_ApfLv guKt!|u
1
l=rPYS1$+
}G-m 2	D\b?KTK,;U&5bF#ddmj:7R{we\~r5S,Fh5O-MPVhu/-Sjws+eNc0/KRV"LB<DgmXmtp3De=koepb-MNd,q4TRsf~WnVP,4 ;o/+5t/!UCEa5AP`DC{SD'?&>uY[uA&6U

c;cf&#|@3~w~yOJ?+AF8U!?WVY>@9(;SpF2c^5vM#;6:.p?L]HyAaJA7<NI5CUHt2~7a!Y+Z<f<967dk$	W?	}EBgMtQpmv-<-o5Na(X'<*ILLOK+]9IkWYw"kX<0^<Wmq@_pU[}bJ=lZ'C}Cl(U7}_=U	/&x`6/<$o34V3tAZD43831KP~	o\f8&e%*tE%Wqr;p$,
8Y{wX:H)gNai[	4Ni?9A.FtBX@&?P9tvG,.+A#@RKKWw~?,PFd0x|;"dSD]|#:@25<PX9@\VMj:uT!DkdYM/)r_U:'tbz{F[~6<<*>A!(^O09DX0*k-M+8!I-7t
H1zoh3>"+;*doiTwWow1FF39K[aq/g"C
-}GLA#D^Qyf=i&aC[R?3g'A/oE-qGQtDA4g0CfC,:f\CHa~)]n&r3/b*qitm-H!JmE;RT-i{-;]~I
GII}RA2;mmt:;wP+{aA:,6 .<X
.ed?xX`[_e{k%bA&VoP}-r[35T&t4P&4~2{VZx0~1,vr7a)m7>`B.BDUc(6I9i_}zAKmhRdWgT}X
0/;3~]7h\T('mnfy^Im|]G9ibGJ5 gP%I([(9	lJ$LdaOqsC}+2xN_[Nt,qc(_?q#UE1(P{@'$O">! Xt:Z!lW'Q9*>p\_7\y#;gt=	IUX^b MVj[]%Y>< 0(w2E?J:HoOa<v~W-mvIS=ga'w`;	4y<VW%Ypo\P#AgGb}Z%*-};e'4U[2~i>QP@sq{e[uf)HeM;$XYqh05ebLti	]kjgy.QZWn2
W*AjWAs\}W6_D!Lh9=958:RWy:
X>t+a?H 6[uh9ddUke}@w$eE\0^u%/'* #b\s,`12@X"&]v	?}^X=/	w9&.I2}S>DP}6'N$7G8F`	/-WKL?(LeQ
2|7;nyMPU9u\Zm+JA)]g^-xQ%LA(_b/S9B=cG/YIaiq;HAG#YgT^JcIq+!p;4*w=~NZQ- vSKX|dh>M@OFfr}4=R*NP9$Fp}i~ENe4E6PvR/(7bHiwLkP9aN&\x<ho%`%Rf^.EmR{elQhC9kriNU.)6A_W9duf+uX9VW44LN0]Zsv]RP:atPD|~yE3Nl[/;2H$>|`'5M2<$-&U[y=7;8jRuB-y|
0TA>==>KqyBuuN7*ea5QWVX-Y+u-H:dV\AE|;78$vkyZi7#sTfaQWq~
	vM(15Dm1ph?_W{.7~R=|WL>20$/06]b^)X3wu]f\E9(CWp_Wo)i|eq2rD4	d}2; 1UN3vD7?PW/w CvIq0tu>mNd77zUulPNriT,Ew$o6e?nyu#2
,MWKWyOov L	TGZ~Ws<m{WvgWn^}rvIHga<G2Pt-w6.:1e'4;V% (I{QhD#>\]sBDD{
Jr-_-CgQ/	7#f^\aOzM p 3w:.{DDe#4$N+.E8U8TQ$ShQ&0%O/pc+[=o]fx-T2ol8GI
}Pp4R>9<c0Uu::Oq1SwvT4x2oK~YTMUJ+N%>"KF	Lu9!31:JS9KOm4Ad<C8,$N..+z?#;m"*\Pd2f|?%e|X$cY1'yo4{as. ,sxRR\;UNGagV"y2)mKe*+{G;L[>3>[xcw1FK>{1Ad'`Dkl-D#(8KDKK()*Ms^i!aO8-p6Z(:W>6`4]=k76jh=vDln2;[b6N!rYZ-O61vgC/ia*F=31&#`la*Z6]
xP#	i|z.+C#(eX,M+@<-O#:8>	h4t<*PlVA-aC? (#~,BG=$e7-3OP1d#s[7wm#ZMAH#7@tjgpH]Tv)q8	; Chf\1G_8W0G ;tbq1=r.FF&:DA0wW\`+fW!%`#Ykm8!VA/TCc<:CH1TtI<Evm8dTZs $?60;$ts>?%D-wE"tKJqKRp=.-[6,+IC0uv<V.x_?qDv:Ni,#*2Vmr%~`a'<dm,S7:ow	tbuNDL([M0HbEQ|Apk]BC	R +y%=s(/J8hON'p.%$G}lkfEm{}y6&O/{rx
\g^vd[KevL=d-dl:iSc7 9.2p02;ZTT!.B-%>,/j@CoF|DK@^?QETR_uAR!(=r^@0	O-5g}BA!H#S?1%F!$b		YN7h}QH]&=!MiSkj{S^{^1+QU QuG#	jInie]</n=RD7qc FqV~
U''@G0,@q6+e%/Ecj]J}rYa ZDX_Fxp #t/P
,N_ yae1rB}:#R&k	:KT>w>4\;Th}as^kB4,b^J_\?fDOb'uA+qxa,r6)g!Pt4].(x?rV	`BEL15l7C9NljAz_I&%j_GeO<O5s>OTnZ+?qrSw]>f^xf)U5)PT+NYVt5!DCS)BQytuJpT!qQgDdDZ,dND$.x,fZ"bIJ.ql!nIi.X|8aa6S()!K+v/+Cr8!k3%?]VAe_y7B1DNPnUv{w5|}t9CE!JG^sqHr5umX^UJEPo.CZ
u1Q<~Px<?84X\rnUW:cB}&kC,]bneC6_=.HRkaB>2n;FVK_uJ0kbazUZJNjns:|2z3rM/%4v$?|fpgR=MroTGxtY ?af=1~Gi+HYC%OLe3V"b	,jsB]3V`aj75R\~H2p/b^4Mc	{5TRX>r=;w8'uT2OODU7tQ^!v/cLo/\J$b-`:Uf'N%og%w7KDQN=*W(rbhJ[G<C FArKA@QBXI|bEAVo`$/S {ObU+F;oq"831Y0fCT)2;>4U-R[;)_cwVsWJgiN}^ygwG;oaJ@w[	gN.4>?+	)Llg0f\(8tZv\6)FN'i2F 3_(^RzoC5XA6_E"A$Yd(na*)ybx1(ef*cxJiDT{fuu^3Z?`gxYBGlnGQ10a~rvjmZS=mTh%)k!UJJQK3N:]wLElCf9Po@BJ;'@OYufB+2;@{KN\YyTsOT=]]"5VV87x25T(1;clbPEq<cm>Q4-sg4R
[@)Q%,oaWStTfpUTLs4fvbiQexH'y]g\,-J6HJMxj,*ie;Z_w#kMikN%.Qj$xFaDqSZg.v"Ev,dpP7"(q/\GIZ-L=l]FP&{dU3?qv/qY(>UrFxOY$k|]bgC$S^}ujBVltdDPl' mCz?Po&5DOU#V+W\\V)~pPR|T2xl]0oS<mq{IFS[I`;qMta*7AXZ>h`z[Njii^IIXZ3z"F$>*<Q?{]
`}lUv9oe?U?y}eOmIQL 5aI- ;4#iZX`wMU^U+m<=ywu7M:O?1,_sGB^:<zsK_SV?9:e/l9:{<?j<#eY6T,J>8(EXvGP$[{liBN|lUhL$M0\g;{2q7GAQry
`~E678MSEl;-kZb48dl@8Qbv-+E1tglj0J5jY+&*Pk!9d(&pCPVG'c Lj!qRTyQ\!U]c]nQ|p$k]Wyz!)6hGczq49O/m~
/FIj=0\pM7C|SRtZ*":,!sr}UQfQv6	!vpL	<'GJ}}L6,/RxQ-,v\tVrQ"DrNTc5evIbru5;r#b,oY?	AMA>3*;D`ojT	:uSR(6'HCcV*uWtsVf<MIm3P}|{]:$v^Dj}%KD':^4nAq*F-lrc%ul-2):XrtAOjmNe2c"Oe	cW;&D3mz]1<=Z`#VS.l:K;4q;1Vidh7{1e@T)o
*_ST,+W3PKx%Tv#%H{>NHCk.Jc''FSi\cE2,u|I6 F2eP6zsXqzy@*hbRf/(:nB+Z7`@w8A_y#nv3qlI1o8 ?gHiDH#"N6rHTN:iQlzm~t+W%=DsM5;(+\1ncqQ=XSiIq_%yqB1{L$_ng*#GNocdy]NCv`p94@F+('7s9oim;sz$T{]wI`.N
eCEK@889}[C/?J[H9ef!9TPVo rQhV5m9 zHVomRc63\ Cez)u<gj9'tmb<+Kx{YX0V]d:b{`	A3#.@l3tlA]*rIs)
c!~}D]\l&ZDbZr{.B~0nRyW
h`gByU(H%~4*XzGS2UH1~@\cm2c* T(D+hw=4]At7(Yz_p^::k?QyvRpvX=&UC7Dg[K5AwVn)~Fo!B]wHOB#\hc&$@W9jQk3b*@h7lJJ<=bfM,IlJ8A4"\Z[EUw`p%H:d_{{TY!]n|/%,[;!VsO]gHwF->"K7hh}U;|I60Acd=v|w'="zrp U<8V MHJHP{=A+z6,3;	i5Bi"7Ll#=D$`&/cPi*IjbfA,1v|:Fvgc6YTQDu=FI,0SN[D-d@eI!yf.8aPM7L5Gr$=VGE#2/-XR!|[c-	l=Lze^t4|K'Z5)`L=dhl9wL<ZZ-RuE2XOWn,dkwcCC.fC@tbA2w~W_DZmyD6cN+@Xly(4tt~= f?ntZI2;K]l0H1Lr`,m5BL1)f,okN)]!Haw.777@8p[Z&xzR;w5`Uizr?[FAqK0|,$m].J7sle\L`K9SCv. au|c{NO&X	_~p~29Wo2vrJky&
MY99dtP|{1nR*?aT5:vi59{"k/Yg,(8j\~wCUa6o}0fq_YqZ j=P^MLa6Vt;h`zy{231nr%lQJ_CKrQ[%Pi$s2$&yt{p[0AD4IZjG`HU`K2}F41g$lw(YJ}r(eI>#.H  WToEc:=p
wI65%]ljS&g3&!VTH0s@Ewr8~3i%%1\:Pj@WVXV<Vp3OZ6O26jcJ3CsUMb0l5kdTL{:+m$Fjr!4o:L<n`]y<a`z@&Io&R\YG3O+G}@YH5`^OK"]A|_c~%goB5sL?1
ron<71Kal7FT~sN5\|M/TsYZ9DH(*$-}X\6p0k^291O}}KGhQ_l#oyj,?9)%6K?MEJq|ni+.D%nQ65~KUP,xqAcqP6zt.qfJilxb;-6q5`'2J*$*-_Z(KmT?Eg|WjC9f47$Lc8Uer<-l'W8roq.U{]=E^-KUS+o+n4vKC] I]c|hzWZ,z/m\73$PVV~f6$-H$$7'hy/?s:eQK\>gs;1  YYV(
ap"KmW&>Q>x`^Zs2,V84fav<j%t<!d5FwmNmFkAC.0<cf}G8ldjdPLR!x
}dzB}a;Vqn~38LP*HD!7#V1f|z%^Pea6uR,RtL|)G	[$f_K5(S2)5|?3'Q=j~g%.WU4#e{#CLQ"RI/FbExId	`)@N:)gaE$!#s +LT?Lb&wq:L$`3k>rvViJX7#oXP60_IwHFIInFDMLDr7d<Njv*&CEyv_P*6

P2Apo3E$n^/`D>8KP(/cGwM"+W^9Sjd3g	hZ*2P+vj}.[i2c&9	k~_gT$8|Tkst!u6 	_{ZEhW:<zw$U>D4RxY	yPoj%^F[xjHkW3^e1._SUN	6'T]Iz<T(<9ux*@F]l`k0<}?oGLgTrAJjP_q{jy23LOR!/IZ_5UU"9j'>P%l,[X49ig'_z;JLH}|o
Mrk~RI>.-<Yn*xfN_^IN)PF"ckFY&+EV<YTH8YvcKHugVA$H39%Bn7qrtO$pYO:8vhiT]~9B)mk0[R_p9Y-UtHgUxwU(Y)OqY1--5iK;B[+bM"SK++GbHh.E=QQO>I&|IOe2B#8B0MZ%7_rU]|-I2Nd\$[89lzuWvSPku!G0>I}:xMnI}5H(GrEpX~4ZOIY05@^k]Dr3x67}+{_ns_pr,y%LKj-iX0:}aYW9|M-[ZFH2,LhZ[+x$%wP<_BTQ*wI%PNyMK=O[zJF/V>g(s/fRH@=x)(2t45E1N5G;me7fgcn -8?[+bsTbRx!BlZc
))+f{W` scRg3n32r7H"3WW>O^Egz81j_w-<rbGex3i_1{eksMQmWPhXn;-W]GW%W8m "!]%R%HPPEd~=Y&P'WEnOWc.IO"O;qMo$zB;xho8STgsAPC	h
e>MNldv#N`kkFCR122vVj!l|Aea<u8=5!=|Wrr]Iv^5"/^e(#Zwtv_MMXc=v|d@52=f*zSGJsPo]AAVvQ^6d'/SmdUD7Q/evVApsOd/L,29bb%D>>]KB	jI}V~B{iVx,dO.2|OLa	,n;Eu5\O+oZWP=$-&^NMI&n(M_DMh U}tMx1f^d`B;ycx/HNRVdJq0	g:5jC`P7]ea!rk!Z*3DG~O1uL`qSW@J{	&D+wpb81th~F*25Z>3(;h3k&wID__esJXk@mRxfG{R%F'o\Ypfd@h\.~	;CD[9,HN9V1B|h{@aVV7Vbq3`/C*DHNpx;ImPB2@?Quee+tQvT.eHl}58QIOd(]!)h@z>PYW8}Sc-\`883hb|n5[l87p4:}<MS"
tawqAz00o7AQ}e8w!2<$!C
|;RE&fR.kK0`9hH~]e->uE4m_YrWhUux<^]|+;hFv}F7{*.{Ws(7kuaY6=$
DyGd`!\e!cr0s)k;U_^v"rqh$T5\zECWe.j<:8dfce(p<AU #z0$9$24Oe.G>KUY`;,fXj'_:*\'/EJXCPF"NhPW ylI{;`z^rDIUY!60=N$-2Od_`1}sLqps,.<p'h`	+o04Pr5SA-)&')O?[wx ]jh~e["D64F%xj<&`"LsHY"dMR"2,EEB#i?EA{"VO31Hb")94Y{ec`]B1acGCr'4gs:psE,2HDt"^;^VGFO93,@`^"Po]e%k<G>&u'J1J(EV`nIX[$7ekO{y
kPl`RYS$q,jb[&\ckGG\iWr_`\8&}M=81dGw!<~El8IP	cn#/7+NM"`@WU7kNt3K]f3L
P2@A phX?2@ssE0F~q?8HDt]/dKpsY#WjpA"l3&@9'PV,7$YHDMY	'_;jlE0_1^y.YDiB_QxHi)SM\XOZuZZ@3xm/)Cy&ChwSJ`Nisa=:#9}{fC]@c}=W'#@m;Em !qgR-N,'1>?y->VQL_YU`G\45ZPMV]D]4	{_N\LjtMF*b[w6%AYgm<[Z3w
*.,uI*]-mH\MKP4#Q+	qsQ-M'xmXT5@`;`Hr9CW3#({6JIFp`ZC#Tj|1+1EupDYxx2|wrJmz5j(1u05*6ypxF1d{9C#Edl+ELXdfnx*2naR)Efcd2t-a\k7Y?s,Wy#\|sf?sf~n&x-Z{Iq=:k4F'~kL|rOmvW 	9tdf>:IVz6	>8JBOhE 7ykMhr{xcOmPmfi5o#T@_*30mMK/b.&J'A13Fd;lo2%ABvT:n9!b}WeHt%5Zv3x)SYO-gm]crnf5IAS	SG&mvopv	Y?#C~d@_^)'pU{nHRp2
pUfF$lOu}X[0Z'l[};W%iVD=MVbHnX0e?a0B/@VioYn	e#k0jvrV?52%C@`UMK>44P9YIX>,6gN=Z;m4BCjZrsljMwJeRDHz:)QMd?^7hL9t;y/1WWXCI%QhX('"[7O.3V~9aH_rffrV	7f3DD8l(H~AivOs32jx'<$LQ#rbDc]}7Ls"]jbk*o3@a'qZH'08s r{p1XpN/[b9&)V	.L{A@dizm[DNF,L_u^ 9\Dc)s0M-[OE6\t~n:L2nB7Q32^3f-{7u-Z[7zioS?	WLz,`dMzOx/B)Y5xT#*0'Gh_3WF??;oQRys<<W'fo;
7MFYF6g2Q	xK=oIN!Bt'5^_(!<25|lSFSVV4OT+\DmR:$,<s".43%SB},wF{uel1A`/~mR\W,K=i*a=(T}B2&"Tr`!7nm75=jrP7k4_HR$Yb}LUG56uLFsv:B7{?1]v/]
oe_Vxy{Wzy3o]Zu4L[(wpzg=JT6+km6TZLX1[._CCvaf;3KRY
u^Yn@<,	YvtMvM`1Yj^<8cF^(6"<Yi/3y t+hm`I5`5xx7`<a`W"HGwi,} Yc{!co%n!^ZI3:NGqI^f%}qwt9Fk x\qX<L|;n*6szUl<t.YBR\]ypb$WOOz;D@A(B"@Q%c|j=>lBzN$sN;+<~70nLEnwCD#zpb-	G63You>|i?#z&QqUQ,cTC!wC;EnIO\ZmI('Dj5KOry<3BzH*?l\lbF'y;	BU9'1{hT*~qk"(7k38a0O*<;fJhm'W<?[,,xm+RI"dH2!*w.~Z[	T?,z+F't$HqYs	Pr~s+{:uk7KO>T	3e~:]b{:ZT.zu?(v-r:>l)_q) O"Z^u`W2(ppDa0@1gl/F|4+=5Kc^^ S<`sB[]|PX\?OM3\#iVwgtxH;l]-7'sv/t=BB2~s3|tpird!|P!U_?vjS?BHnmO	b@p&EPlC2t\.]D	q%eJP53~Oi/#qT#{w)-pigkJ
CVn<E#V!#~O-3ks}fYahKrAp's=7B!coekT)^MK56\B\2x@Bf7%_[$`Ed%AXmT6|jP^pB&C\5Fr,Gp"7X(BdM{>p#P:%syo(0gJ]>Qlz"`DD]p17\8-oDPg$fJ4].l<11V@~#<IhbxW|PdL^'C2}Y1l+L`S@'HaZz#VwLA-YB|g`V,AFceDu7=ohu#KZDEonny~RCU.F/"03N|&\~'o&H\&H<>@ktGMjJ|{CyK09pVXAse	nS/P	M)V[>840Y](WSq}ZWzF ]`7NGRP22Fupo#bC#3mBztvoy@BIsQ~m]1JTE8XE^'Cy
&}OjH52p;$iI*Ts$,CTEA46b$5/$v75g,MQga_A}.F>w=i;.8\7A6s@F{OaY3'%9"GxFU^]qeP9G~`lrid(Mk@%&DNVZp"ykqv"t>s2S8u<	AR>bG$u~o	!-pUMA9}6QhEic8|&6Gw*~dh(\DZ3VbvOb41&80,/
-am]*C*mOmj;y!N=.OTEbfU`7D7N~jjb.7=:h`wB{['sq/"fcl[EGG7KZU`Yw|e-3E6LP)L.L,O(uO+bt(-G@qx5,	pGc >afiU*p3e9.3qf5Zn}3"7%u) h32kNMoJkU@H,\ColQ}<0rqk^:G;W	,|0pkm\0]i	|>C!)Co&kh*IYNO\gwV7Y6wuZi=!$CQfft)[E/gTUY(:Vgi,c*=:$2J!HM0Q}pT6}5~l|-w=+DZ8V%|+8dbu)0g^l2H%a2$rmtQ(dU;-D}o<yzYlsPgIv:V\yr%Swdh_j2?L{8r;#k^dD
co}Hd9UIZ "lK=S	W%27tQ!'^Y}EeNk0js%\H*x:#>R,2m51K"B,&BgH-91|2dQj[U3|yhB{#s}u$zG6c2V[VD'i_DR9~V"}mb33j_HhL2gc	BS5Qm_V=;r']k@!*1;(Gt*/qj:
6h5?BEY^v%?>|@b.sNb}d&gi35u&\Q8i6L
zz5P@AMyT>#3I6`/i\'tB&Tk[mael-BH7g=nB%le!yC2	+{60?K
q;LXn_; ]a8Y&#'%.{,NaI=KxRogs Wh
n|}_X$y)$LxVs,]fPYIS]86tXc'W\<DvM)_=
H89PXm`Y[? 0Yk4fy|+<RA1L[N?A.#Ze8%0< uUUOsItVwJ	(MGS<k&l#|tZx0	%'y;I[M7K2`L&$,a0nqgg%De>m^L[0B*^R&&*+a"\}u6}_5Ko:p.?F2uYS"]thYmY4	^,"_<t^Kl_)YQ^FszqRE>P6"}h9mW#$6[AVzwjq;K	2kH#1|8^$3k!/q~C/}4d9!{no|J!S30BMq_b*M=_/1YTm6Ip'8%=H"*OYn<m:!Yc2HbQqQzzznJTFS&I\~od:bS-Z*(;M,whNz-8!h7 TyAW^/uc>eJ<ziuq:$.mS0.d@Fzzm Ikg0>F`K4}.1k*zo4~Y$T0.H?h5t1.'#W-~}Qp\"#>|<Q>TB8/J-d{c`Lg[.7|?Fk`2)~[&ssM2}8q^heVbLnyBM12@NO*<B5;z@:KaS]AT?cf_7sPHcr_[9:Ai"-femD|q6UmgPKmZ]MW>w"52g__xMM\q6MZLuIITbIY[RSL$^}un5nT{LaBvrX!i^NSIu'Un{xc>
1OS)/]2Bj+b	4"!Ik!?Sh{KBHCwq/bhNiu \ls|M"#bhQgl`m"m ^F\E3L.v#N`-#o*	7$gGl}rRi21PJyRR^`#"]27Os^F!-%4rEl{4i'gdUwg<c)9N9_T4(JlDb'E@8Og5P~(?
NnPWd0.5"f	M~qDFjet-|JPF"yXPl8gn}_sP,~CB2m:-P3joS,B9H3N""uFOkz5s2	f`){lcx2EktxlXq,Zm8c0dc-b84@OHq6pZH2#BAQyBlTer%g=8HjhU$V2x=K lDUc,IU_UZs!g8t9Fx +sD@UbZifzTl8vo~k%R*+w~f?B+!A$)DeS/z_WxU5R=g%ui36
lTEsIssyY*qKU2ttwD98L@2\H1ga[u/n~tz>Im0KP4yP;M.o
'Xw!8%cH/	CL`MVKA43#kOa>E9rFWv"(H\s>Dv}%qj/JUNL2\v.0+.X:do.Fo2{hR+o'^S!ykO9{T;16ZtXG"F^Y;h]pZ*ksv}LerB=fVO<"@IOn6^sa6a=WbCCx9LJ\Uo%H~Q3f<BaNCbZ){kueLkJ?=Bp-Txo0~/1[<5ty9brXw^(cpS/;!P+wohko}W=6g7Qo^Y9
qaDJ"{jXi+ }K*"[9F[R-id(? jQ:SW[=J3c[.RkMU
oi:%&6\OJ89gNXLt"	NO :kgWV|]:{U2o`?T
	%=7wohhM:nb3DOx^X#''sQE5@qMyeTv7]@.$32&Wr09"%(!:@rt@tXL(R8!wI0'P*[J:hA_-v%uGe&n\@0H&Yq;F)`H0l/Sl7Zzg^z+~xH|Gqh!<#B\H'yHH$Wgr)52<$[!fY6!op9*eSXh'oTtd_k2ByO[&UV^nGZAx`8R%ZRO=d2e#%	*J!bYs1qba*nuyJ?x<JSZtFqOTf~&7xo2;'9fKP`ka,R6acB\XE6~
,LK;TN;;;Mdl}l
cS[%.[4Uf	#[ =+R_
 eU(h}h)s0oAzjJ,E<F#4Vw9KO5jfU
6i[I]mv:[B?H<W@.qEwCKW-$|sr5vNn3eXesa$d% Hq^2UC.c&fTzCXF=1%)-3$m\m?~Z	F>
BCaqm_SU:wkRna;m]dT>4>Z&cf$~%)>:ppsj&~Tf6YhAk {X-G}9d}?WEn`+?H$<RmY;-2q`(*Z*n(bse&1mnQ"cng+*xPy\sQInW,+1X'ow@*QkOOLD#>jf |zz[=XJ[\y8yOa'[K>En	8.%'<#@Hnlla	~*QEfw%s2|XBOwE8=ws/6Q"+g6Y7dqUf*=2F}PyIRP&OLXQUD'bx#)z(ppn,P[e7e~O)s_3$',u(
?Kza+,XY%!<CYSr;Uzb,7p(.My".Y#9
zXj;7rH]5Lt6dbguY:,/vr2p0
pl%{Pb)s`N#S(I$63Nda\j76Be5

t1lHP%e)(gr]R/D8A48axw	QLwhd[?C+$U_gr8@-zam96X:SgeFZd(e2}V*yCEK(r
Ch$rTulON1M9eV4WV6jaZH6z7l	E4.h9<|B.G;q#O88kp/w*0}Kd<J#qe&+V*\JE?0;P/er-7"0	|D !_+{l/B?#m}?~([(s\$;(X)P9Z
H=*-g*B}w<O{r^;Y^W2#5Mn8ag@K;w[)3diy>zBmU;D}|w]|GPW$,9[I3G[:&2=H\x	wwqYvrOz`HG4RuR8n6eh<)OK;V=dpTH;b6%arV.KR2D+'Nj$+"F'!|Z`*<lS |>t/{'Q^,%R	0ZfoG]l+Wx{Bz%9zK@{mY^-8f5IKCF?:x_(vC%L$LD5O`a-=8cj5KQ>adu/wEqt7fR"I~5_vU+>>4_<{ZkCirQapRqHQzqW7vKAA/E=8^Y<e.O6[MWc1RZ K<]0XQuCS3aYQ)t{9ZAfzgSq	DRPvk:kz;0QJVxfGD}spqanc^~aP[^8_+->?00m'<d@=YlwTq@1+lrN:
JZcpU-"9}jK.|2To}mqF~J:{0o_#	ruVW,W2uJH 3_KpEINa<4'A<LcI~*@@3rGv_r(B"gTsZuEixj\cci-"K:|Jm}dGt2>-o^xVV^?MW)iPGpW{&`E_C@zP] xMm4	M0M	k"66ZvSh@{b5[m;b(&eWa[>m(u\zL$W+zx"73_'5,Nh>@arQ(VYm^Ibx&[
&o4B.es2a1eqNW#w&9_]>{a#7hm[% Ayw[X5*]<wzk81a[pp?wl8i!xKF0HvC_*KS*y#p<wzFqa1LBiw?yGR^m?V"jS>MoVcxHDw@6;saJcBjkq'*\Qt/KmI^\](g@1#|CBiQ\4yD9WQDd)
 'HuE}dovO+35E&i(hw}&ectQ]$5FUV-PD'8-yGafiiTmn}=gjE/@d=`5qNU'*MeB+lA8R*|./Xc/J|`yr?ILj;l<("#(F0c~bbFbDX%%/;uzCtR&=&.i1x` Y'<='iL^h<5n(oQ8B=sw#|/*H\^q/P9}\	fm;3ABhHn8&W
#9XhMrwq_-fNxsN^<YYW#A_ll,dpy>LG,recn}:,5s("!,b)	:(Ang\-nW^Qi0%+7
xHI3k#CvxT|wFN;d~<j:oC=X@_4.^AG2wOy"xs	4?8U<F ?9X(ClC	r{r^aFG0-;82;8s;N|u[O=zC'%OF2A=LT)XLuS'|vo*+NVpacHdR)=\	jq`gf]4O6^4?5}S2d!Qn/xe-O6?&H5	1!3bAWG:X&q^2$D7&\jU%fhWk"<\	e)7#
{f.1-#F6tDgt`uO4vO&Z(J`9Tx5irn|otlxz3u^#h}S_&37Tf#j*I[@K6Aw`8zVfuKs#b?t;@^YC<\{gc,;87}Af0RH[?^1f2?<NB,.oiI3m~wi];=.c{RSzq|{g$3	i='hT>_mJTY&+ZPEYr8AHN0/!b$S/g/#	sXgC('K4|EYk7KMSrd{aaMF,zE5	o2ExBP,L7(W"'6#y29sTn>umuJAMo\jo>^%r3}(<m|$/2Xum.vKmm(E`#yG;Q=%.9GZcp>`;P/LY*C/%>&,=/yNMR6"?=<-:POz.!vI?<%;?nYHX8/oN7R35i55PlN\v$B*Ybu4^XSo"&+$}::2(X8	Z|Qd4Zvj5My<v`19ZTxnw[Q-E%[Pj5:wClKocNn(].D]Btnrb,KF;Po;C7pQ)Mzoy\&]'EMAwC/1P"c!J&d{CJwW#?1C
Jx[b"
_#RR<M%fiG/=fy{LGdr<Mr+{ff%&3z=iFF.d[vUqvO/+l	}{=:e,=TM]Ug,0'@~qQn$?m%d'=`>&F SEM<iI~^}RF\8a%!iY$NI5&O3,&2T|dyX8	G
G2}!J5/ R-zs ?+"MBv:m:0H$`s:
TM&ShVd^ MR-SCt+nio&]8ut2TGVk5tZTd)Q-Tj1SU[B)(W$ma$o,^za7nS'|u)MqbRqDP&xxfc|#gR!dq"?RFK4+I1+W5yI3~~WA>OKvSy&HX8SvXqv?^0~vogqDY,lm=3MA%e!`It%0HfzZDlrd1quXr4{.3<@uqJ	[Z1a%~`af6150Yw56(_-|x$axQ1qu~u_Hn$&E4h(7	w-[k+z$ZxQ[ULzW;"wii'MLO8G||nCydV(-dT%{zrjA}ao4oAU.,Ak2EJTG[KN>/bY_[1=%	dPkt)2]P`IFq DW&f%H
q5RhC,+xZB)6P
-~RgJkkBR^q2S)jyOBxxBub]}m)wl3|DT_Q6_gz$V\Ko![&asOw =V?.@Ks"$,9>bw@eP7a6HX$>Ip->FDOGnx9AQ;!m1@RozBbKPjeV<=;wgK(Cb=]t[B]YU.s?zr-pwgMR%?bmScVm@_aHnyo	bc08Qs|jT
GM=0j'
';w0u-R=kD$.+1Ad8-JZ99>g`7Kgx\|#!|^dtJ`Rdp?,.Q*&P,2[eH<L{OI+!D;]{]'1
Y:
x.73coc(:0PM"UGiNE6,g\wcw#L2QOy(VJbLdG0WVeblq\Lj-?ZKb/_%dtx=kK@db~UOL}9{BO2K[sm0U]EN:	Q{:AL IUU/9bW"%(E1]L)f+9
B| Xps=(MKhFwwTdip{:DUdgw5Ss6i]fr&=]LL;#}|6+}jm/j9Y9-srs&dKOPf5m{l"m'2:ZA@1lt7Q#|CNk8@3V3|0BIR8q_?W`;\k,L[|]spW.jj.*)Rs?pC=>p-P8ovY'#Nk4QS:2P=ro,`-e_@/Q.i)PLO}6ByDpb0E6)h%mH9"c;?(>R6=|j^80
j!HPev!go0Z~)
^`H8RQ\Pv\Z$i4tc7;pfswYDtkf)+75x1O(WWN89#Tmf:8`}MwrO}h'wY"?$?5-Scbb4F@@f]4uccnMOcpXkx_p2Ia4Nk"wXQxyZ`1*{,!s`hXH{IBh\eL?!|)B!o [vlJh&z{:Y}WR(A< BFXq$.Sc#&?D5DoP1}5gGk.4Fh9Z`"}AAmhdy<\J37E`|YCuqo;;5Y*%q{}CkHi+5mI]@9	HJ_r4B."u3&N2h[.B[n_$N+HYcI@)hy7#EK0(NJrV@7S$>\sZ.lTtGe^4ZC[DF=yDL[<efpRmqY'v9<4DPp"-mh1^2=un4ckT(\b985>5+\$&`8yN)3A!i.u_Y_I?vTTQsZgVG3)W(7)bOD3b	|x`Z	Ou0&i1l],0<`AyBv>Zb@*I	MC|~WCZa
J#yKd(Jn%_'@H_WL"T}IU7LaF`
K*/a|	_ibMK\S1DhSlO+xl\v+gg`<pkl(a]MD2D6EOyFs0m`X>o%[)UbSqRer)U!V{J7%Gu?)buNOY{h8^2SeVx]y*d"K|/.V0(#4h`H]27H;cF;`?9UeYE]hTA-q&=6cDPn,64<qlt8**VkZ)cdo`[DGuB(jNKd_*Eh14
Z\oUMR"Buuc0$A	GW{8CZQ!Qcv^P: m::OzgR-x|Rs3[{u]lNP&
fqG&p	tWYqcwlSB~M9TojX///Cw`JLvjS&xC%,:}:C';Q/^km?scWU6WYXV}=0?L1xF(8-4$5zH'vM{.anHUmR,.$g;I=RY-D_{bzsg	Q$VzO_p98~<Kg>$5bbuj~Vv=

$/!z46-4A<ak?]p:RS!|ph2@+]OoY,l3	P+{=}`w~:
2]-4\OwCC8g3o\Tf|5KV3;N"}fzi6	m3!}VS'OYcg:w7Wgu0[!l6@d
~n%O\Bd9HGw;[6G*\f[<e>!+
vJ=[j!%q^RE<kdRcj&VlWy6|?#%Q.nK02R(GsT]A8T@X&r2`FkpV#Qo]<V19<p>Qo7A!AZ]$b9]4fv:wN<xf$JxF4!6jk\?V"Yl.(C|YjBqX8y_&-T+yI7.dIjh_<#p6U/r<:/,z3LLn98f\ERiv0[fe.j$1	m q"W#)p6!iExhEdFv10.B/]8O@Q6vt:C*j!8	>i9nh2%U	Lb#1I[Azt71$;/R	3LbCe!V)?Zg5}*?&>d/yBf8=eVf#{.)Vt4X^$M%|}I _;T3NAoAMq^VETs#gmFV/RR?u^~XJi_e7SuKjSRxnNP	F)f/!?kQZ#q x;5*|wfUxGSO(B<Z<P
Q/x_]^w63%yNo/XaH>FCMceu#}8$;?C)L*nmqYkD5MVJ_lJx^[Y)nc1}j?u~BXp.]>~)#&l=nAt1PuHy_cIc~-
2`V7XOvwAFdz;yj 'Vm=e[9PEY'}L^s/S"7n(b2oB
,/Dt>9+(s]hqb(\J:eTQ&D;8C.C$wJ$n|z'nIt1tRJ8];<yhEK
TD'9p?uA2t%W:HXpW=>s\<~P6Jr?}A=ZY#P]sGbkZZ	+>^>,\xcRM!;^eiRq4W]xD=GW-<*0Pw!vBH({d[uJBO\3<U5vLIrfW[TJ\t8Vhw|,io+A]#|&EDK@O cZ?rt#0V:df7}P'S#HA?`Z"VBOd[is [7sFj+`3-ycqk@)K3q:4sn,D$lvn`;{MPeJX6#>V%f-SCI.hr\+s2iJBj|&7M2-b+}b);n0I0:L? -<op2}r"s$RBB"\yecW~R;/_cr8w>,<yKIYt93GdY1<Y;n4{C[5$u,eY3,i+`;
vKct/v/vqB?0'd_#@@Q|xtSY[lmF[.FdQ}Vai)}z(wg.8?oUZJ;	"SZwRjDMoGSKh
ln3Nv|DqpCtA@[#lYN37>tF^Ke(1=hn*;1q{[copR]o(usk6K79R,Yj~q759JnNEzu%0j;NY;
P$9RK%;_GzCVPNUZb<s-2U2>pb_J@43C"Zht/l;
%^fD`[1#\PxT[tbZmU fXz/Oz8=$K7kT>i6BB62|NM*qX_:1ixG2g\kufa.#%*ah^1uy,<t$h-:xRek@O,? cO/N|\DH3[ToAcH6e2AVd )c_7RmP~}zsip?s*@Oi<JDDc_4Y>;')V%\1_o|U_0|GcoHwrMh(Ehy`@tL(X|B2Xyv>sr-Ye?DOUC=v:[{8@J:/%TsZV)< Nt valV)\tgh)F\dI
/C2'
/ g9!sQIsbe;_J:=NG\6: zH-"lMX3C(-S/|(RH_DxLu/zIGd4n;^0wFwXKpU:#A*4Ymb<pPf4);bIZh1"p@3eaAgz
 =[:9.%vb2D=0IQgr^3c5\s)MW
^|VIGK@nt<B)%FT):i,dC.L%-60acMnWxFd/c0Zg|RadakMTZ#frgeDD+tJ5(]Enu~VpL
)TSU1P[3s`Y*/""NC4lPUn?r%v{]G@yj%_@ot.a~}fe,X6hXu0_Jjtlcqv/bCt1_wsa{qO"q)LM8>Cshj37ERi3#O CwxRq M0$JJBsBM ,BE#1nJ@yXlpC93z2&U&NhgS	1euI)Ugp0Og&*|^5''qeRaRv@^vF$Dt6YNDGx,JwK/T;3ib^FqVL=$: bc-Lh@d;5X=-tk1EFR	 %E%?9+IRnvM:uH 1b~)L6*!^m!B%R4zD^;C:25mqS`}!]w;/WEL\!_.}G=[Pp=g+u~fYd9,]zl KH_|&8Y !yy6o:?|Y'=E>6
cTC},PhmY|u0Hl}8egp2#Cb3cMm]?J{@a/&tQXn=4Rni{g,^6C?Pk}KX*;'C#%u6lcj?%&k,jS6SHo}C)RQk.1^|]n{'>\l>Y5SZ*BQ2j5xuPdIxQ]q4E$f+tbtPOPK`{*x4Qv!7if}:[]f4oa1KLlfaa$mO;a*:ix,(\%f%^vIw<O`7IZ_32C-VQT8='*,]XJyaH_k:g\d257Z|:"y'XYe8	]3z6W`oD_"RJHdL2 ~vn?N@U![5JDNMt6cF$VU#h\}3429-NP'|1qA;*|(Wiut(r(?'"B~^.>Q-cy9I1JO@|h6]0u$)**BL^ !0^.kd%@nK2}d]</7cC;AGp4syE:9iTJPA!"";sK*,C$m/_z6Obd3sQQO]6{KSc"cB5*&0s=w9!nQx5)DVwl4k@"po{T+|W`J|tf|`$:%YgzW]1;D$N4c0E78{**Xcah?	DxkR4Gv}6dt\J2SAY'%Ss7PX@Ax~$,!8Gn5b~sj#;&$L`uk*qQX_2R?4[Ttmunq`!P7D2FkC!fvDtwcZ0YM~i@fU=zHp]r2q$mos{~km;j58p'Z1O)&FKQMTB:o5PWo`B{W	J/hSLcXEDzKf{]e8>_H9V:
kya1}mWnC2A:7W%s.m&}@]U(9p)z8b9[/kG.dK5q?074IGX	\k,i-dofgje<gsj"YYI	f\-tZpi=}}IhQRq)+SbcnZZBA7)<vHB{RF*L Tu'\xWQ6jB@}}&x7O@/dw&TLbM#%1P@6lhQgTJAdaR@XL!E<%(|"04$Lo--d-bWoo^Vp0/YdhQh/vH~!2Y243a[Xq=K2N4--)I>	m-7v!y8z=o(>Qffn$<%\K]eQ6Jr4e]zlRNhjE^l\^^V%x)Sec,1`>"u0v^=4_^c\V-V-Sd&	Hv"vpE1)]ylN}GOCk1Maz?wB`IvSavQZ\.V"L3^&F5@2]sdsVnBXde4`j.kMS#;LM)lQ7Vh@<U-F#-,-~ZT)VT1p=e'ARXHYw5
t5
^Vk&1sn660qK>\brXLLm%
z$NLCgj79!rpM)${e!&h)trs}T(%wwz^7B8>[ec{7c^(PQ'"qzgK0i\3/qLQw'>x)r?DP0jPB!M<3ISt*[*x:(oDB49-A8$YfG}xa'rXco8 '&6qYkW?1N}{O7qqb##k5%UhT
mz6SIWTCTT1AIKE1MVVKrTDTxbj[OX}P"KMOZ=*"P:\};Rm9F|F}GjN[^}N<4g#7p#/QWkHFj9.<[|X#49)C	i-;5S
HI/{C*d98ava|ruL~"b0uT{a5n	
C6)<BcU--;}#pLRv_N+L*x%07qO\0Er;q75EIxZEP= VWV'R$+FW>Um.{e|RP2()"=;g#>@%Yn~yqCO#{iOZA$Niw._	So-H	7hK:*_q#QZjv6~bdJ2n6_C9puv*c45;G=PW/W[HG=!]/[RMX\9)H9LVk@N=ivBZ"w301n;T67N"?y`}!E/u&?`,eGLUg- K3+i5GGl+cq@9e!~3fOv2N6g4@lV/6=vxsUwE/ZEjn0f)Ww>mG5?B2BuC=1q3@HIQgZPo!%B{
& H?85%rct[6PJ3O]+U-)fKTr'0N6o9/#qcG}G}l(U@{e](%MIT75>{CSWy)w)/BPi-PrUpC6s~Z m~Ak|W{ |dgB;lQA~{,59+|_?nLd@ol,kWq9wNsWR.r{95@^	Kl1!x'T#oA*&'mH`bIkusVnG;m,*fIXf{1sG'xs%Qe/%{3Br:h:WDA.E^zS;c-_c!VR[%7"KZ/*_kx
TG4s+CM<{	m0t>cZ+[@Zlu/pH)1#[`y1_%zf>WU&76'ac[d`
KG`jv#(w+qz2fO	u/NkJCePo{dpG"4R$7=(._4MpL)i6F5*p4zW2(=U#r\V>v8Kki<@OXCsAru}Nj&ROEj>{4Z4L&*^rC|>=(IVCS	[\-H>{a1[Vl>q+CM]YAsZyUnsDV__mu&w"y:9~e3w6s*?i!^VZC5r>Tjo]QnY!zds3k5I{[X2D@JXy4?oXm{n2o{?.<P!:gfL2kpbiA@8uM>GSoc)Et\^T%<SM3([,Plw~n=T+Saj67>OOy,d4G,?>U]GAE_jLBz	_C,+dFUQ6XH#*F3vSk#[5Q9F]Hq[mcN;0wy6q=q3fc'oYtISono8M9dpd{fn5+Rat6g-=15nkVeBB6<5F#m*A,ysmaC,^s<hx5ah%<>|+W(>tV*<Z u'a2&Xb0U@L5yro;,Sw^fI(/F=WyXAr|UA[(LI%ht6E)],-mB9eU!ATuV&m.y9!u4 r@~:3D;aZW1p(An*+Y&GN@ydTdw:_9l2?6m0/@9Fg*1^[Dj!mC_ocZm@.{$[4uATPSs]4MD2UIb(^PrN;#C}!2b^y3$mm 3h+NeYa zVG>k?3iZ LJNK?8Cgtg=.
}#$oC4;<mURQIH*`k)y,{E'&xkKm!kFoj4DbSQ~e$:e;	Jl=?aG lqM/iA@RTQHrp27-27=MAN	Bx2@=bVFthm,v.pc0Co0aK[-:XS!|hw6PiPMEhb!X.Mfqa@Z;P].2Eg{r:ct4Z"rBHw$bdt`Nb5>KO*6O6j9~DvEq_3v	,[n5.p/q67cm;*~%Akr;-	8AVlA +;R|dw9m{eS`9,5o?6N
`~_|:JiE.t*;US!3M+'F}aPHE20n+-mXHP::mvhpwC]0SCp	/s~o%HZ!iW-GXaC5755[PI4_LN5];VN'6.f'-nw$e#|eD?[}[@lz0:U#*w0sFL l1B/Z"J{x5J2y/=U\1&]\o#fw xN}'4[ttC5tN[dgMSu+Tg*.v%2/h,G<; Ss<b~H;E!K\?r;-q([k::t K:(&'Fb;hBO48nq(@7'c>.Z8y]x3h4S.F<Z)A5T)M/'Ql\xV	G<F==U)4X$/,^;5P)AKrSlIX@f}TS'8NZ'xX+LdmabOO5@{A&5Du{$zRIw JWnALs_p..Jn>k1eP"N,e2{5a>-@Rib5vH^0|b& ^fs=GlahO+?=D+bIfH_Dq+EWu-h@#jJ%C3}Pih;35fMBBgwS.,n{@J^m=+&*8S;(ko%n{/oU2a${xATB`'d3yceD;QHUMu]1!"$	+us(ZosM_q&A^"9
qqyD'?b>6%*5h/>lr,A,2oz:d6aEz` w!H}!_<M	`VKu{m7P(F2j_Ry^pJWux5m=z*W.W\{A";S3M&qarB`>w\rSq|zM`WD0V>4-a}T[U\u^ i}@ kvnlK:)g"4iWPes%E`aY%R&q[s6D/+6fr4[MqWf}a8++ml>oW-(pO&!MDRKYuz1?S=JArw%;I3sV,`SpMIDqXW}wrP5_},QW	7
v}+emm<rij8XV|R#gGGkQwt#B-#+yc*>5+2&^T7ex|8.XQ?aOj
FlsZ/Nu8[}[QJ3N&C1+TLoJ{P{+d(zu^d 8W((3)~[?j5kmn}_-:j'#NlW*Qs3Nl*"C<|@-S.y=j6tc?v,st%os;Mc;m@
Knfl%;x:h+.YiK55Qa97C5Z?ed2,z:~/=;&CdN\M<P?Dz&.lF}SJ@S?/;Gi!I"<cl]9Xe<go`iNrsDM_fe=LX_[zw2r5J'D7e&
[#P.[.)X6QMN/Vuxh=fk:XXVU<ci#]y#pnU!oFJ1X&Lk:@dFD4yrk*w41P-w*Y)PJ(H1BPU1hMLe$!gl6g|w2sCbL(R+WoRh+cJa`}^QDSQ\FT $^[xBMx,O/<Rn\xbT8
pJ@7/fleY:iUS.)p9(a"oK^y5odL37UJo@f4Dh,j>Us@o}ONM1caP5~7 ,s7\Pp{VU-NP-ZQ{d`n~R59lmTB%t?aPAT'E1
ui8' 
dG(MhAG{9)|?WC81VEg*5ppGDqh}+h
1!W&29XC6&6Xd2i.45Pyw|}E+l;N`X*B3F{crVxa7`qg:vs=uX"n|zgeJ"X-V)dua"(uwlZ?w	_q`Fhn/XIk|E`Q|,OI\Z7_RQ,<|$}yd;w5d"Qk:DcIu)F}O~3I2%>u{w]Qv:@Q{d YAu$1z9beqp\'8=b6wmiu1!Ne"pE(X;xQ}DUC3NXO
#6B#-$ZNw/OYDIw0,|Omf>%4oIfWijk~!uJ4
3{u9!=@-\heE!K=QN[`VE;}aK`^@ukW@zN~&?pG|D"Q5\9
'^;:q3C*'AYczofi@aLRV?aWM@o!hAE@._tJ^|IP=-xXif(I6n0&"2h^-:vq<OSI;[sMT4fb;"-f=pTXr	9\l+Iibz0.&0x x~KKcwL<ZwonVUk:<EDAK$2]MG<]
K}pXyy!:%EWk7H!?ojrWC[7(]Q!|ND8%AqziNgt&AC)k\nj=D@4wwD~G ^k1?*&!K|K<ftj;MP#&9}1fM
$?r2qm</dc	0IOD{D14ztkk6j3Ji*qOhPo?:/k79|t.a*5e-Uk*O&B+I=x<^ew==&+s?}b%
m@f']s'>}vy(^+MmGu&P/FL\^jmPcI]/K/(4:c(2VwR*mZE,V%,x(KmWb:25 Zxag>ty#[AmlcYrtyL~DVWZ|?5+xG*FBW{FyU(cQ:m)	 vbZ-*%z|@_[RY:9G&J|gik?'=JE/}	YWM)(z:F]a6=uqewJc{NAcjdeuyXw\5=HP%~%2|:|3q)'Y_v8q*+5f!I6h=1ebH5}{]MA[jDoe$k']>BrFG\< UC"U",-k$}5^12j+^EoUd>kK)2K7q6UL;e284"wPkk%@9lq!PZrH/[Tk)^dH{)>KYuG45q$D`*r5Od5gz!Hx.Anl=%A{(8%!L1]qe8z,+u>%#_O_1~t`!*EuPCZ"u1VRO^CipbujTTJ#03._Qe/Xth7#n>UqIU{(6>N=.a|m.-n)i'.!7_zwa7'6?(#bkz],+fKDo$$ZUWHlelDVFdG]UaXvm$v{X4Zxus%FaV
BgxvEI%$Q'ap@xU;WVc.BU|[	{_e32{1!2\O&'VO 4rpr#Y0UosZsDp/*4w+EI1:yg!rNhe]\x6l~m';xn;Wb_QFb1bY+>P56F0rOm]IiN(:VDO^nV!u_HjoG;frB7Elf<E<v9V;nQsBH
+2]
F&<i]5y:kDnsWx@(+>&b}Q%FCrZS[CS@?u$57 }*hx|E/+&A]rVl6'MSw5W'!:({qXini-28y:\ef#cKn,5Gk_%Ev>XK5?Os
0D/Z@U}B,Y%I4tSOiR? 4I)iC{~V5CH	NnH	?VIB`<H
jExcW)rj?V4~hBux Z,ueYK`u@5gO^Yo5pvx:jbixif\xb *9:g{P\"&kS_=)rhWJPRU_M/)yr)V`\>CL%*0>J:9ym?4DIymIZMM=A<*v<!eu$\$9&dTwF)G)?BG;8Mh#
a;3a-Lx "wOo{6mN;+9DjDDE]<@y>7W@E1t2{wM%r4G1
l7.l}h4ZB:{>WiSfHx?b0o:iwQ&4F}B	gqz=*}y*N@hu*-!jd49~W99tx&
$~S"OwqAu_3x]"
?b)7)bUVG$}&-]x37LW6M<Wz@[?3Wgr/713<:Q>RYiFO&cjw4$^*5/f hOqH"1&PYkYRf"%PmC|y55F7_WIe_ G@#'xwWkkg}1EM4?4SQM?]F	hP1.$[@Xz7{UmewIrh1G78=RZT<yo?y!"W4c^ogBvsT_*3<c&U-n<S1\HTQSl>~OvMj9`<G%z!>ECm^PJ&3|@{	+Fn,BJK(Jv5(Q4C]Rt
rm:FQ0*b-Z)!tC%'"W:V_#E.p[d4
$PLh8{WL0bA7>9:&l\'(TU	fHSs$9W0)D4fM"WI	YKFc9>`SYc`WP.	hanRk*Q+G-xte38lAZvVnKdR	Y$-j4f`WmZzx$1_Cq9a%:(til+|TF7Lyr;f<PuorI?=Xi.Ky8-13}8
b'%F~&Rys>2H4R*EA Z7F}[BG#jF's0sqJ_'w" u)lS9H6.gI!fAyK&*%W+NQ/c2_0?8'Oru.v3>,:_8;MVZ-Vf&2]t4
(4+g,HoZcYESM#)4V(H4)W1v9#lhL50w2od}}eb0{<ku}^6OPhV`R=/T~!+$LN@Fz3\K5TL+>I[9:GjoBaKb^!IN(I"<ZlMlf:4^qm`0o7K6XYr'\tM+Dv`sfudkitW4}"3t4rcwv>%\~[M-Celfl3$$CNk#sW6t,hl	LzS{zlJ/"KiS=*ywR"fxZVEw _Xa]x\/1fx;j-it=!BP&nyg> bB>U*grjv:iE-]9qR?Pn_RE1]0Li!]DY5knM7079c=6F=p9J_*FzfT]W>V!CROy/<%Tf]K_):[`L:+.Q'Wxy_-^Z[-)V{CAQUWdj?[qXbu3d__}B|[%oF_AdjOO243\M^L{y1$rNR6w7@?j7yo/J,=D/`!Q[{3'/xRz~	D5XBr5\odF8./Yp$4.wt[-'~t_XO8-Y:F45!62sDAwSm+mt*%8#%r'92Bux6NB>c>Pa :*3Q<GrXplI%vy5
{X)JsH)y	Zzv]oxo-AhJod0vlB!3+HCu-OJx[`)VP[K^'bQQqzdD)-wm+g=6tb(c}>=BrJ$!"[]ZB$eUC? ^}#{JTX<2:^.D%JoPDq6Q,X1XG#8&Whkq&4Rs"9gfF_lX2("Yj%gb\#aPAT&_b:n3jZiWRp]D\!POThoIuR!jLvG-sYiH?~ULyO]HkVczrA)1Qf@Md]>O%oNU6h/ON$LZ]'VJ:{}!N1lc^T[2dv?wyRzvgR1mn#4C8lVCJTwMoQuxwNqY1m9EXPx&:4=1|lPXyT;J Ptp}Yl\S	jFl0S5jqwM!d=zxmxabV`Bz)nHpjiMB+6>#[FRIQxat|1Qd>SleG0xlaiKyo,bL_:jP}h@<F18\i|}a-U^w.&dQ3A2tX^*{sF(B]Ki\)M{Bcb<8t<9/$]%3v~ui4?
9&RE<Q[EQN@jN.fBziuQU`O[@<^/4"O9$q|;Z6/.Yd*;f"B?Xn+cbq//1L]!x
8U:_Eej7y,.
%,GaQ'hCkG6T,Kb[V`1:\+;A}F?Hu,mq d
q-1J#UY"[`vK+*&WVBG79Cw%.9!G+FQKAK0#rkAi(.~-{8}}*	[}TlGKw*S*#HXwN[:YXx,9&5:>DV$Y^j{J
# J[,o{N8]WbP/',,6uol[m/A|A=Cw{b]7#LQ3HONcW_RZ,pDi$8m'be@+w|w@@1/~L&W)C7jm&tK0-Y**dCFckg$ClpM/*uW+7Qw'J4`e>0^_3+cE0{i;<[ah?0^7[/dU$(2}hBEnfstC,@1IvpK-=:K&zH$eVbn}x"gBqDf$!	]djiEZTZ_V/Og3Eqg*c=ujS4hdMWL_6!^5jYG+ EH&}a"JV{Pr_{^>w%+6V^B0,3kiH{A<CtNVO_OLTX|/r;1Fz-:s:}9^s&cObEjnE7	fGe{Bl
	o@!jscz)\]7Qx~)"kv-M8s`y+l`2}z)kSbHVF	.	
?;Rz\m|ld+C~iIy8J	QvP;71`I59Wq!BQpJg<unh9~{Gg>P4Z:U+X1ov_tg)R5*XVk&?q=m2VKsvQtvvcN
%,rAy[Z.6DGmukF"\E"cmZvA8N4r 	?cr]Zx5Lr#+,lw}_KS)a[!2,@.kI;`4/O13]jGc~NXtK
M(LM/*bodmh<=!Y+Y0*Z)-20?:EAS!9#W,:Mh(s)0]X 25X_\:-ROZr7p\DqCmFN(mZ)sjez)Cb9Q60{kZD|OKIs%N!%$GanC~ 6tw=a=:^$8Y-R(g"-N}PWVg"lppsSq<7r8k`\d+igL\T69LU-i?l#&'YIZ"'m<BPzU5=n9SxZHxWmGSC	^Y^~`N][;Ny^eYf9j"xTgPH&]FMu?s(msxZ|9my9PC7Lr]f5p~KpI=/:ud1:&r<`qp67{(2YZ|K6 B%97Qs 8=mN;n4ae[Q,1Q[=z%JWjLpeCvI+kwtilZ6'NwL#{U`~I4wfPH#C9s zPD')eI'Dxc'.T-s}q	7hn)m#S`^hRT	Lf2s5B;ww'p[>;
G&yi}T%I)7rJ}#kx$:#K\':TB/|*\7C]sY3#`Tt=^TL&CKWbI|G2?[!
.{
W@*WR5<5&-IEx|,*60`}M`Yx		05B/{UZeeqFaT)_L<5U(6Usx5[PZ@G\	tip}_-*-Y\vefWjG'xU3#9tGw,Ib\zLh6z5+!9:)zxR`h=6=d>r'tCGiT_XZeA33(uC?KJt<N8!#dfdTp8cm,gm5A@}@ |V`<HW?oRtO~4[+U!{q-NLf-&{O%_3mG#@1YZnO-Wv"Z%$Yg[;&+7o	Y'y>Xbv,cEp$$s,}(.Gl+VTi9PeoK%+TKg[qJ)aC(r-Z[dD]CcS4oK4lFKHc>K$9DHKR@sF",U*kr[}8JQ?i	KzPOhiyV[}>^YHb_5H,EbcP{L~J":7Rn'rR^x"w?:w#>b)m!SI)N]wt}Jj	T/B<boNl>Qe$Ov i)n(d\]ajL=n#!))/ePUz$ZWj=oy#	Z-h p ]z>L`	qM0?/4|,=j]hdb6Ri]~e^d5^x">[sGy6LR
{tN@\Xy/
hPefP?hcMi#rit:ff6k|]pjENoC}u	*qPr'-RDSH,s7tt5WhpOGX8h[#;W@qB/ZXE-LI69x]0	%;I/3O:H#\s0c"^Hzqb	.6?={Ul^}>WHs,ekAU"S]F);&G{9:qggVnFs{ue{e7:mdAlB8E=1$
qsl4lKqkf
[_3c'}[59rh#S\zka0gTywLrA	^q=U~8oWROWE{<]rFQIr!GDh|HCrjb+b9@]|\=M}9ML/>p2Xh~>p4!8ThY5h\q3]'CKx;{Vt'8>Y) Ch@a;i(<"fRH5r8;Bd@O'|nD[?Z@vu_o#8ndz"72y|n\wG4+p+3d_c"aC_Y4qH/>rCc6=eHXBTCz`s(Xme!X7}1-:AK)NiAxm(Ug2u3Q&[Rt	b9,S(7NNX_$i@bW?2,xMvGv(M58P@z=pK}f/RjB<B(&@~#p^C#NRD0'E}hRHCXY!$e%AAe%Wi4]4D%|0'OlY>}U;H)Yh(k#LJTzX,U!1
7qW?x?h[jbXw)sPdE0c$w?-\4q64b"uLfj!@:!M&APVrOe.LG>9.*NT&c/vXo >^>3w(?x-'!a(	~/l^ Tf :Mfn.#R*_XB937}gxBAvJyK/>+]5t>"Agg+_lV;(3[B\R (S6k^EK;@'8D;jbsi,J4!hcY9woYtTqjX1DUD?J04YFp=-c6?#Ny^&\`>V[u}d<&@dQhHUr6~fT\6y)njn&[hR?"Sh}Bpc?e"[6X"X_iT?d6|*qIyDxd.xKq?ecq)%)nmX3c2t/K5TQG/}ZMD=Ufy5vXB1M??L. $&Q|r[o;|_m0AoIT?THV"E(lvjw\wu5zh`E-4#&Q8i@9?TR2W#TFBlD|*!O0+nJ%#w&I6vt/
H <0ym+y5'tKv(5)`iii3 uU/S'[/*%LNa;A\>9i]s^X'//k)OvGI^Y|q@#a`(| 5y?@aObklY*
hc`<auv$io|4q*)agSI~8F|*\U8WMIwdX!j$>|EnD59$if%E@,B\ik@w.rD0rC7N&Sf=nHe/.+p3Am:<=k(6VjZehUYL@.<bkZg{mF>I%{hdKL%@%<2He.mJ/g|{6!&
)cwk8GWM|V09o1xI#=:(*2\@$xK4S^&fw^mYg&{42C2Pe/dAWZjLWM=7@/sv'cJ.**Y x8%D]Q}=12;(ezzem=Sz)O~K}+>uKJh3zej%b<eb1*|Igs[v%W&&v5GXjh42rlVra~9wVj5m3o.Pl~IJ6.U hT']^@3T?iPUmf:hsh!g?S,gtfE-vrm%yAd=!|j7MLQ4vSrs_Va+	-8F(e^UK$z(gjC@ruYiG@9T]>ZTLi=Fw;aQx;$'4Om6\}F
^{&p,63#`]*Bd{*JuYi?0R{<f_&^AM&|E=*5vN:1>}zHn'IYpP"OH\yXFPP$qJLO<IK2BP_VXe	rlug'w,D6+:>B
2{+44ZuEZNQ5l4:m#gV/TtU,(|gN#7#Oe~%OTHx!:Wdb7Sc%6Km(|]8$2j84gmyMGS@iBxL3_.`e^D%(aAq/	z!&^x&p$;B7G@CN_\a$:Oc+aIB<=llcn; r. ny%D[lyhdUq}nij9C_z?jDaa.46ZR
.8kuo+RuJcdu_Q3\xz'"z\~MemT^[K7-=
M}_`_.9?F%DV.l&*x\bia?EWd"{([G940p0	1 *Ih^zgSHqkU8:_r#1-SGeQ\ :ryZAjTF_|[*;+4)|JUl'TmmTK9ZN"LYmzQ-, D:pm'e"Bf(G0+2AR(Po+)PZ]"%\eogI$Zw1R6 SW^y7XS>|mVl9G
<:[9.PYGWEb%)WN/J5	9:_E3,6tVepCl~8FLEgIoPC6c;ieek|fWSq?]:YkP\FxZW2C%n.f$/~:X	6%R.Km]aQ ]cq1i`9{cj |P7}}cMsGW<"lCEUAQXz_Tc7}YQ#a#KIKb}Swljq47h7{EJG?@,/=a/I0sG9-V~u5B7=%1L-kp2aEs^)I8BR+?2+h
N]U9,\<:"zY=yDY.v5LnX@J_$e2{i\76~>v_f
A_EYqbqEu+b!%.,UAwWC(sv9"_)Fki%
}wA9J]c7Z,Xm@KN3D7bz[5AKL\LOE;ugu} *.z#z1'Pz_9/P	w\?>r>60i<Vm6+|'l)/
x[=bX.^K>?K9!VR/,
g3mM~8!)\9DU5*;5\MgX~%Vf<,G	%$oUMhA-u#}qp79L>Xhum&^6]Bd3VH9$^8*Z~B<n(:,<v)c8$!h"q/mk,*==Ad-~W^4v,A3~Z{g&D^hjm&4XkG=A_&]fh+BN0v)IG)dZ5GB,nDx~QNWb7H\/wz"f?*_48P6SO[gy:D;q-;xQ[@*,8Ug&Xm=k;MH]CArwCjU r(ce=;$dKmnBueY+Ib{K136fPcn3hb&ONSmw,ZWzy%CJG20x"TD7\/jwlqU6ie.\q4zj(W"'%cH@~M+Uy9Co-t4ZigT'3&W|t#*%no%q0aMbk't]p)dclsJTKBb(HJ|6.<CF.mt(VG}$](aEAH(U9TzgvQI>L$JeGvxK4? '*hNV*O#22'^9m3>*
vk`gz	n_	a:im#DI(B%Z!3e9h"]^9o{H@Dgd[(&SGEX^p)A@gSD0\3FK3CI'haculV[/mI*#Tv/U"||:<{zNr,~`F?'G[0`}{ RP1 L:t)qMSK63Mjo /mn*v<d|>ReW'c!wl-Rmm24{e>/9V)?p:J;Z<4'A!COw|<WbFK'goguh4O3rl{#o	B)hWbAql(d}Dx+bYFqZnzAdA(!+KtKg3e|kkjbG&n[DXk!XrFP`&yA$v<Tab>:#:JaGVp{S#&P"h)`nFT#OOvBi\grg{%d3kQ%{(H[D:vdTky}ZN<1UarH|
J
6mlLEP^Ffbp/(Ibi[A@>|x.5;9)lb}ecjeU[DXE*yVqq	K_)chP>aK\A/Yt4Uh'c!{.>$$zF#2]Be=SbT\AS%jV-czf	{<E\iEg%g4{$!6HzITIo6zG	n6+%d[pEmvA+h+$9 ""*9[/x?8YlJg3|9G%I,oU/QlyNJk\v#-^EOY;e4/
*t&A_0H'CiqUH{Z-xv75Gs&7TUQ!:N/=x?2OUW@7yHw<~\L{IZ'ab_nK$d@[I_Bd jcCVYmaOAO9>k|4[,P.2ze]shAXDU\PRpzIC21}NI5$&f20d(tn|LH`[*XkR(w!|\b:?-@iRiLE`AS#{,FH<q[un:^6=XatRe5h$iV7s;"N>M,>et8+X(xg!hxe45d-1Ps4wxz^h+vFMkXWlUZM3h(nfLX|4/Dd4lrf11JSF$ju<R{~9I'd)9[>,]d0sD{;Sk;5YReygM*m+4AL8KfYm}*296Tuu|smdC(pf|h*'"9>Q~2a,'1,8}5&8tO8^wbPj];?%)0pxHoPsUO1i^<	O+Vb@)O+>$Zr`Mk_CC9KEHF8$q*q{F0r@=U}*L8KNxIpBMB|
E;~@kUckS&0AbkWjV+C5ijap0_ZtxDOa%?&Ad[m-2E>utg]./SB#[D=/;Set6J-:&:L?f}5~u4H $eRxwF,d!A)u1^"LA-|bU[Z=`&'>,'i+,k
"OL	9Muu[UkgG%)Q6[vHp]//+N_Pc;]COpD8#v[[wl
\FquNKKcH/B	3s=="Ob~5\	`io1:"UCo?TsL7k*iuhR1f^xN_#@HyL.P#0zoKN%{S%fyav";/DSo43qq},D1O0^vQ9mkt@FGOHWv9(
T B_'s
)%$?o;ZY&}Ps>@d:ShqE::#iKTpFNz3$&~.&#mG|aZR_Gmv!ou"t9Ovs3*L6)g@3?.L]mT\cxlr3L.WO4Y?Et8'[h1?V\13*(T:]Vl#qaGIF,
@-\= lwkqt_-`cm)YF6T('Rr8M9tYF<{MIqmP9\zJB$EwS\,&9t6U3a-BfsdJ%WYMFPg]*PX3K#(07]>B\sjp#rlZ	Yh$2H[J<Pz=B;'MF7\=IY'Tdcpr,8_% D.-{CHk^Q?nT3`Wte/J8%#K|@kMw\9cQ5:UzOQ@c5b/'21R&l/&hbB9x|0}Hy6^R@%M!6j%>p`'
qeZ*25{v;+`8D7m,cM859?w-%dw#MdbV3M3wRZ4MC*C-/Gunq)q,C
uEFPEsX)UTc[WX4Y2":>	9{s?ZzsBJ`+&@E+^@VCT|E
mjK.w#+yPd
1UfHVQxYO#6:K!q!PBaQ|4CPU C2[|o\`Yw3:4k\RvVl,cbF.X66VHQO(cz3Xyd1JIkhYJMn,k@,''7LEY*q@Q-UI	1k8m
oVEc S93eSiGTbjfsPgnoC
v_2w#q	
oG"Ouvb%Bi*bCOa
A`&Agd!)p4d3O1x	O e1[iV>{kZP.YtM:,z&DN&{*uZEWA	S`WcRF1Oo.#Rq/kgF-#."H)V!-$
FCy(-3^=x!Irx7:&NXBw_DdH.du]HY*Be[`g(kiB#\D0u6R_JY.]IJAo
O!8tE9*>m4Y[(/'Sl;(+[^oTo?g7]nFg2->`yGEh;Ti}F?\#if/K$`5qs5jjSXGLj:ILp;z[LN~jbd#\#`P+$af{DbwC*5B
=)qr:+0eskGg(/5K j)lT]3BDD,KXg-Ct^c"0_Q\BU0FKzV~AW)o	6%(vY%msv{N"x";efb~5?'zCJeJW)P\sQ=%^EsU
s.h-9cufHk-8+mKz=Djz1DH"I[mhCey|=Au0%b)|,Q9"w,<9(u2x6:'14<v&G%\CW@m1{LhzO'&;^&RS=oOSNM{RX^!f(G,G{\;RXkrlYK,Wc]AYys0WBTGG;|}Nr2oZ36vh6% OdtN8?HUi+)%t$ $SaiqS{."H2.isj/wVIv;qv|=j'Ez3#}t`CwOh8c@L23\gMS*`YT&
3^^O	HkC<!+sfV	T xF>{7"~_f}MJ9t*I.xLdq.>^Wlj3|;R}a6rg:z:NQcZmsl*&M&Y#5oLr]	\EI0vMeYg7\YT]^[Ke]p)xoWs#60G<Q-*u\7	dE{:Xjbr!G7kaQt_x'IYKnA]>B:IGJJ<+vzXJ^fI*,#9J*y(lzl0{[v"D]I)*w_z+9UYCQ/t3C8kW5x3BMg:=)$?&803ZUS~tu%T&KDY\A1Xjc'.Z2Lti{@zteTEGs{3br3RD9rZYsZ,G?(/!M9pENMcPB^*\"/k
R<W`mfMn'>4NI9N{%S=j)6 /*0#a`bpx0OU8M;W0/PdxV5C_iX%!5yTZC/2	\89mh_	RN~VADgG;S)gK>[S0daBjlc{>aX6}>@T5UQT*'er6xgUTB*OjooF7ErBU|E+1tVM2,kREh9cDk**q^~Wp*Z5yzDjOeWyGFapprwmzH\QR=',d)%%|4&0bbAK<8BG7|5Gy}H$bu2tE4G)q"#/J6 .TUp!)RyTKox(
&{!,Qd#t`8I2enG^zdY`b\%u~SF$3bV)@X/(m4$dJT3-^}-{{?.%g\a	S15r}KjLnK4(6ZtT+f.`;A}
Yz!&q.	CE`a}>M*3;Q8^L-C_!Bcz6k-}zT
:qv=JCm8n4L7B*z=y^}j;Rx'ng	6*%ZeRMk;Q=.?DUSXt&{,IYRuOlTDzP$S^o@T_Ew}Vv9;~~aj'g{a,Nh=R6#a=~S-f0p'B:v}2.'
>*T	PxC0+W[SK!l`&)i#{&wY=-|K(\s,g=g>NtPq7jk&e6K9UK`P)]!n3aC|v@`/E:K6ni%,1dI$A2a[:!DItt#7|Br'VT>AAM+!NVOr<),G"2L(m~r<45`X{;EA|#}P9IQ1nDo.:fh5_>}J>#-YX~gmU~|gfSnx5PhsIG{?h[,+QWM60' p1Scn`dL'CcXbV?uM~gxwSNpm*Wl[Gw5S_?5d~:+G6!C$<%|UfQSQ@zma[I:^2Rv;"4.t?6h-h{v7nXew*_:d52hEtBw>(r|/@#G`%;<2<Nb"_;LTWC5++$J+LkrW924Lu0QLeb+&ITG51^_0$\MSP4|!}Tf*$ZBTa<`g.m^v~7\?QIG9-aB.I>G%+gFc`(ZSFls#a+Ov,/Vs=W#Ze}/0dBuA7?&ulfIy1d<<gl[EIFR-r>XrOk)bl'N:H}4:N.Jpt;EA
3r?lOof*$\&hmVES`eLV"k47`#mv8Y	
mOG4KJvDM|<N~c)N*j9KSGq'1aZ&_mN5."O-w|11Ym'D|Gp~BRZd.1T%)&_Z,|uKZ#CbGtcn#v<\yg[g;['?tG[G}mP8#/3E=;~UF:KH/!F1N,?IRbpjgPPXdK?jA%a^{9B`on{	~CWA	nF9[li4:RN*01O""x3KvTmb5<d_0pI]hW?Dfd9%t}dOgt^fC#M;+n?
ti36N$*8I="-_ru	}*+H/&Ew(YU!oM^_~ew#`r|23y'F aN%[)QzouJOu~eafNAccO%1TKz{	l3+Eg?3S4nP>aC~/R{`p9IB2'Ed	CP~5i0qXM}YO/~N:-PBC-E|kgZ=GF"NKG6X.,ytx[2c;Sbgfx?]qCCCsOT4dli1*7O9<qbFy<a$b'Um;*r,2	tu|&.etBm/_T>fG$_/O |\b/UjT~#7+6dZbPo|dA2O~ g$=P~_g>Cu`F.F$Nz!sw:D~*4w7ulf`o5'/:M||8<CBni|g=EE|@-m'Uuorj06Rz;?s;F 15@
=>y1+x9/"J9Jy{s,USa	QgG\e~r/}3`pFN_wVAM$LXW3CLQ,7y "P?FA2$K'mFuI~`d 7y%ySWt,rO!(XwJ&
QUWsx1C
TJ<`fHL|`Z27j3YAur"k8^1#(,P^>q@(K)4V?6I`P2*C;WA[5	@fpW1G)~2R05L-a@<}N4oQ:[O!_D&l.0u#0}YhxOX1?x`i;B=g/\IU)@M5L'U/(.pYGll/l	jy\NYM7u2az=wIP95^nYg~+&QfJ(=0:DSP* q/l"`OGu`M+kS^8+-:$LrQ@SuDd'OoQ~~\2b8O@Bot!iIdw4}udE0~K+V=)v#;'rH{GXAMqc]PL2#N;;"<
0)KBA>wt-/I!gvSz1TfKT+YX)eigu8Q7(,@7CeUHLz4 i4h3gd-ID'6TB..K7sleg}yKx/W)<m	cmB+sRu
1x'%A*mnD
zf/#7Cwbk)5}9r
wA85-0H}xkdm6>z#y}[$Y%6c{=G3+|5qOj!R=d|5>@VBlv*wg4;.^J6FaNH{VJ-z3{Mf#{'81z/"Xeo$/]`]NO+{sN<R(&R~	%cL@FQU&x_H	?`BU_H	1Q7zI%bTDJyVk@,.u1KoQ!asLy$+r'{^|}QUrUcL/]dpFj;[~xQ8F1)MeXgM)\Q2vP0R7QK$e}q`-~BXNoBvT(<aVD?tNmUvh+]h;mu21$.b[P[@(m*tQ"yJ-mI
mp}q~{b3guS E~MPkMErw 	Ofe7<u@|g=E-IWui<*	S_u"6Gy|o4qp
ccsvBxypEkT@cN^nB~bb+.8$*[ [4|Lx pN-KUqKz)!<:>QCgQH^=c;o/8:(;JSm\\cC+}d%CV~kpw}iH<<@h[T!7GGn[*
D6+@6Gy;%;^c;[	]->>C6.vG+B
R/$LuAr(
{]vH?2:Ng~%Ci_T6]]:ZMBS=Mq$>,d.9xb~%'MUc6Cd^4p#du+.e*[k%rd[L*"ys6rRmP~-Y=Um|Nu+)3Y1PG~H[xY),$Qz?T3Dzn1hXY9 V(&8=YOuS;YenoUU`CwWp[wS"1e=.ZBF\BEUW,*LGy39>'} +)`=Zp>`CQe<Cv@XA]@!fR>?iG*%QxEIxKqe| H2ox(Yn\&!0w<Le:=8j(%S()F av~W
TqYF9g:9:GR/K3jH&XZG6v]o_XUu"%e`x<W|;%J%?p*oC,W%8J6::bU!sR/CP2(&=3t%:NV4 /[kVG{6~<|PYp|16iM.nc,&$G=#;
vA86:-<5t2 7Ph"(|0,:#)I/%amK+_HX;$d-!]j;ib|y}WMO{ Ko2uKgImw?$I[i=@qQ*5_Cpp v`>P!,)c=i=.D`"70Sd/QvnP\#S('5oAl8eW}kx/I8zTRVUn*V4).q&6R;6| v !DG!>N>Pw&W|\f+VeaZ#y'X"F<3Gm|Q;p]aDqNg9
-!.afifO%AM%#ga"w4B>kj:<ev'Fsq3%nO$xI 9*&QB(w(bv\gdb+!s:-5aM;y!q1Y")~$^qGLuUB6?ZK6))6B#(4)Pg,E
3ZNk4Di.)+DNQnC0l'=(hjlbB?)eq/NTSp#otsMiIT(g&_tcc(&\-&`YCet|q`~JS2F^s0N7}AFA<4Egs!"0FEqPgv|i)9=":G\GA#xN(u_c@iOUU8Vcq.hDx:y4-StE_%\n
(zZ?[gHf#M	9T\G7)z!71Wk>Ig<d0_QTw%3Hr{w0}`2Nuu8]xJ=i!4xlXd!	jy!Oa_w	`uY] %=n;Xl`TGV'
.v([lHC#y?y	kj>il[dY$45P/A&SNeD*3"unDm11M{Ww\?Du&+r1#f^IpzWbYLX:	S=E	H&ILB(3`+2t_wq&x/k&vCcs1 XKP=	zReE~$n1!W&@L%WPP;h|MzSyuvqpI>x0Mi!T_UUPlT 0 9p+93Hu^%t7IA?ES~)wa*h:G ;]&%-yq/qHB'XQW_0f[fl^Z2hS=+zcJ:st1}rjJu[[0uyHn3$s0#-=+0#{Fx.748HBP6~^9'SsU8PN2S0|=d7+?7"UX~+@arLz<)"O'a =
_-@7c"f<R3#6LNz\])-P+s#"ius," >e&gDTn+,Q0_tXP;znBbq3i<I<InnqKx[n(SV.3sk&B@4"Z^2FSZMhQ'BYj87$p2@[Jb&mA29&!xgc-3.r]fsxncxxK?/F$L8,;lGuDRj&LIvL0{7xJG3uS>zCZ/G;{:T,3	eMOW)mW"wpM$.3;@RtdNJw:\T2>md[SX m+ir9"rY,3?o,sj^gK6l$DD$`m.iA59f.[KI@gqpSL,4^g=-Z"\@"sU\p8T=zxP(A~DMB[zO{I.>g?'R1pA#WY#J#JA	eK1Y9zxRQ	ZD@K}`@tOkk1"0 +}p"TMz	$OkSP-53;mLis7J5H/x)Z'F$efE`NDpV*.P&H)*O+	R2#t!g+q_kPG"w>stC"-.:I\8\GdyNuu,m)Zm^xE)t=C5Q",bXIkMio<Tq&^[pv4.X>:lCEJMQ<Ly,}%E79_-g'YHxuEk(5pdJtYi6[V{ t|vZxZU\Xk%\pyjB.&"YD!oJ{idSniHS}wWpjj5pAuGV+&00gA-k7b<BU9xwV4TU;P1xXys!?ni6";X`GqQ!(4
g^
`f	m{ZNLv?D[+WN	t@lBX{|;,5*SP=)*_}Km\:}%& 2iL
X0;|s)=nws+-t!?3g"m\3<,IqTnn*j .j#RK;vTluG`_+o&`B&A|q
z%cZ9qJTiwl$c:bE)H^HjZnUrO@gJu4eRdm7~O,\IXq@-\<b"1OO4=GD_r|UpL2o[IBKp=_iNu]&j%ZMk\Fk_}b`S$H%:^Pl]h t=j+U6^GPU1v@i})Z^es<|Z*r<-%;Q,9!/jtE!@g/6[^"ii0'|l%A
,B0ay%N^_F#5VeYdf<;PF/v_`Sk"!n ?!7sDG]B+y|	v6EU=iA-$w(d4bUb7NZ$&0SI!\?lct?B);&h-c=W^tH?,GF\c=5>J:6e{lbVM'"_9?a:G<^~g'6AN"j!J$IY?+`)>X^O}{gAH.H
.fjMTXBG$a$&[\v3?S+N3q79[&!x,)nd;t	Hz]yJrj%~"r8[no7vjwBf~sN~w4|fb[D-3("OgOcSc~"o|+PmD(FlO4c[y5zj+R"d=h8+
:B8\9od6pWEDB:,4iz1h'czQ.zKjw2vig]vo:~K.Vlm?rynPG;dslXBjYCt{1{?iqYX|-cU89A},iddu4h29/7sSw9i*&/SU3&?UUhK[T<S%g,h7CT	0KO,.! wZ<qQ{,Z$U!(qO7/ uo&MD?[ti	_d}o\p{ T9g>.@jSimn29M%JzvL_o|_nsc+M4^tIS|fC/"1Ys-<j~TwqwR{7Jh:"!Wt2g+0V?>wFTl<a>4b&/8[jIk:##O
hu8F?@,StfyD4w64`N&~wdN|j>b7KClFk>B9p2}DLkU`O,>ep Ku* W"ZY;`7&9132=,5PORV4#1[U&PL9a{)F)]@#:07}M 4`bhose7q=GG;
Y+M	+ E
Ml{-eG	X?QYmwSQGSJZV}Z6\e#	w:3kCKmPV
>]F#~@R?f*5MQC$X[32Lo''Sq0`9eo.	[bhoeu!eny2"&"*#@u)PRC=|D.;kbhD)5$-pfZ[x+;5b=f#[_L:]ScqsU)q@/cO2a7Vh!'vsg/vHLovvOgEF^d{&S
!'Nr^fGW@3u7|yjsW+^.7z=SWro,;,TI_'	ljBK[mH_t|%`zSB0\N}!PZ@JQa`rLk~TNl!|ZG>E%pR08mBTIBR`7<$nn,kczSnH S&eXiA[g"T/5RULiW?^
Axw)~
k*VhIu4O"=_]5="iJ`.a5kWDp{:"Vgb^sT[t_| ]DI$C>ansIcr[6$>n_b>P(:y.2!;b;/7i$lm!
$z>WBVG,j-Yj3ol&05_1)W,YB#jgX<$	UTaDnFgiMtpwLz;`qm%EuLq#'Yn9:Ln7\O]X8`5S!wH}F|/Tfz6PgZ`#:tQm&n*k	#h%JFU0t|ojiN]1;>.=/w8	\)qd:l0LlfE:BPkhq,pFBkP/#&&w@}z}u-_4SWY\@*D68Sm}[vk_Ykg0)cc|<(NzzEv2ayEe$#Fz?Q!tznw^W7#LMNlSMN:qqiIAg+2F?D[x1E7Rb#X =))6m1tS8=v]>KxIbHz$2DM2L{jlI1	c)YA+K=;&jKDXSKe_4Q}D-'=\TfMMwV0,`*c]Z4plaD\\;=^HxZhnA#!$~"Lsa%Rbh[	sb
e:^v"ODFm'^!}s0E_AMq-P4zph)f[jBaK:*/%y4\(dT\{+:f1CMhG-Pa#vB;g_1f:#5$<&+t,FEL@}8C"}[HI%.\HkyUzO+,)U(lCYwscTceR)/X!"7/ohL5_WOHNq;r~akK&iN0E;`(1+GJ}|d2:Rg
0$?>b~"ay]7.O`/#1V/ml$Ah2cCo?mx-W;_;/*sf)ofgdHLpXE*r>wpQ(5
7htovGV"zBU]]RDx2i]xc/S<Et7 "!BIQr(Nf/RyXKn!b-Sb]dB(HXwVM"/sA<U>OGjuy7qW66f$[w0)Xvtj3DBev,E%u!of_ o7,-
+:#K7s_I	<W6LA\Xe<t2WRUE2_s9	cr%DQDM\pC`Q-AW%4G {?).pDH*%\0#0Q/f7Q8a*%p4JPF=d[/Qu4`BC=ZOX(Q>ND#bGLB6(ebBIVU4ey~Swe}K9CdU80an_sLS_V9C.xn<{\d\j;9jV}Y)-'>0C#Cjt#yx%,WgY"2>1;K(EcG>/Rp/yW,(Or`0?,&To3]MV]s_'{\J:$wo[Q8
REH\rf!{^FU*c/#{s788w}ERAfC1wK@W!-bej:)Xx-?1xb_rZ|8vE{'$XakmFKn?ehVjp
@B%+By!LlG-E:%arxdyY#FB5&eO:'d+N~q'716rRiV_J,9IEh|C'K2Vm 3MTV+_"0L|<8\:B(j);hDjjtm
%[8v
e0~gw+kEyFnh?WY3%q-M1ev>#bbk,NMN.9%=n`QSA}F[	E[MXDW[9e<BsKs,fbw
 \:1{JVL*_ ;2)M*h~c.u}bh=n.f!
POl%E|	wX^:QhpX+T[VMr{jYR{S^`?0W|5gte\:sgEgwk-mgFwU^G~co_pdvpU1 6UdIMH2l^C?7KurY
/\-eHN#C)ypqHS~-5xXeeYd>\4zq7VgT
C
<{rGK7W:"btJBmfj^zScM$}#NZ77~=!7t+J.I@}-}5PB0 t[pqB)!O|nGuDE	aNtM{2t+xq:4,"}:tKdbZ6LbxR_$bipNp~fg42Ci<d7Y0+2/#=<;V-H.Fm\b#HO5_$B4!Xad.NC@"0T1xCo:R# VKSv|>u6GPUEZk*@d~_j6g
n.{CEnAQ`dyQ3)&G&GQ)0~?9&dQwza4(B+Ke5x6PQs	yn$ztX>GX`8DdMD8*\8(S/Z?|op\f*%K3Nx^tl</6vH{O)qJ?M;t/C-|}:I9=BiW/_}`FDRGo6/@z.$=v&vaZ4=*UD~UJ;wk%bMopw3#*8v~5?(&+=lY}i:c<CUP6R+!B}Xv22SUM7gCh?\0+Je9rZ`m%;&^v[5e*"ons*P[vA%
 kf@*"@"nlC]%U |&cga
-JbF_SKr_%uTBv>grg\\Z,61`ZffBp`
/Fc-
*L2#c68?8*`Km;q/]<+R4y!I5ql<DwRXq"%"FD0!T)(b*st;-_8%~@stP8C7s
+&1=F,/0Y_g!l ,;rh	!k14%d7BA#Z?/,y=	C{itQ=NV7	P|s9EgHhx$6c	RG</Vn^t? q'K@lnR?_j5*ly>+V5iGqHS[W^X.4#n)DM(k@Q+racOzfb;rWG4{[3v	H#^X?uGVUT%Epo5ruOKZYsyEnG7Zz#u@@N!K'Le)M'KH$bvXYpO9}es5@;A9Y)i?2jU CRC^@,X2Tw!#ulg.xY(KKo$'*Se!tn8"ZO(,	jWTiiKu}W{ZU R:? #D."L=0YfT]<{Iv%"QJs.nl[K_km7`PuNhZ@c&n37_<
O@=V%8ti`V4Eyt#5#"P)BQvTL@_u^\NIyE_ %si1c7$<X51#9chDCf
=Dzg!Jk18N_%+?qM?ak>;!0?!R6RppW"YAo$2-N\#~2,0J!9)K5dPM)EF</|/ &{2QU<xUTeu(81qc
!8nmnKk.er|fIQ/ .d9A3F@A JN$\eRV|," be~1qCOzW-u_O9{U2^'g}RE/.3?j?x-|`mQ3$oZ]<#RF?8:A-m5b.!%]e$k-Ka	/TtLFUn#JvB=Cjlb4W,-SUUj0TMKmI?V%FP's%j.*2-NeeE4j8#E/Rgh<U8xz
d4^6Q8>>-q5%PXfP;4eVX|	gA!_}Z>jLvQj2r\RyW}7=@ta-|b|ldBIrf<v	F
Gyi>S"$)vz"-cEU6anE;H+(u:l?hfmb%z=KT2)<HrvC3AZi'Ey&7R$r>!~+-glHny-_q^["v^^.#]r[j&$E XiEl	Hc1N#g[C`:Y&v,7=55\FJ]~[<F-@;_-^`5Y6l5* h*Y
9r03#fG"6Z
+LUtec2!N6-TP~PgOYkby`!Poj7[xIpqm<lIdaKH[7Bv
}!zhiOC.}>TEF^vr:O~g7Rj\`Fo8BgW2(4dhKTpf	H`Ac1*,m'$Z#'US,YKZW&V4JgTIcNyvdVaI{~zIWVLxXz]o1QdUq<D,_PdY8!oQlx)wDrO`B#O{6'(}`-	F
xdv$j6MGd'PvB}0(zI%#(1A@	dqH6%c)o\s&)8c>c? rVZ>Oi2n*UvNQ'fm/]D&6LA/W-7bV*u{x$31j+=zlwvm?*@.u[3eS?)V.U_'do$Zmj0|]kuI-8*CmWH!:+y`=IL|Elpc&uDc6T'C|P2fz:B>5R_$^hD;fo6fBnq[%P_K@`D6bg<QNiiho+e7P|n#p}~u6lfaXo<r^N(V]\0;,GUT`	#HJxvxaR9lL$S;s8E,`/?f$m,OKCxo'p7ej#03h3s{%Qk7M.6QmUlW2jG>F9ce\5pp~#X,&O\Bw628nr,JUB9qVU" ey@a?4WgT\:a0p)4LVuT~=EMbD8N20&	`{^0aQ=3,U"RWgL&5jf{8O$d;4GHn/N7G|*8D)FgGQ=	:H/EC-B4
4.W2~xVzZPL/pMtyj`(D1u$1d/W@*jbXjnkX:ZvT7vM;OuL{`nRtI=P=3<9k wvG[? Kq-"t7tG.+DkR(l)2
 $T765Z7O&6"L2\M_Hs~/|
4m@#L*P}j?][	dQ8@]EP+5~cPnuLm}iu|ed[\z1yg7IytgP]l|Yfw6o]$q)LmC_\:FA)D0"oYI$JU^bOv_K8-+6Wz;,Q2)S60-a
.Sf
P8Z"_%+8}[y-VfR{_Pz%%lsl;@;O 0Z`g^o7(wvvNTB1&{{sEZekxOQvE<-):fM-s.U|#'5BX^!4']PQjot2AWrCCj|pcED6b
;\{'=9N-o'^6-t|
ef|OUDZOO3_/Svy(djpipIIc~6~!;jI^>@XOT<c(v+Ntx.nVNI=o]iD?@PFTA_'|5gD +5Frcv#C&Q@}_,'pd% .f<s_{P7P'EUD{6?QrXpC/KEW
{rW^$HK^wr;RH,o1\MEv'r=`?w|I8?Ndtjw@#F5G7VmnYRQc:6`Ys*Aa+ a$!)_mk")NT?>oCUq9m(6$(>49&xvbTj1ql@vjO}|hLe$7;H|O9u#I+'@Lvqmuju[1FKk@0&7O#sw(-#9k
'npdq"_C3_6F*%-wHnlc$w6F.I}[bTXaJ
TEG>g<^ohZa?:wAW0!`_PNM $JSf~`HnybqK%nW"VH-8-\A+H@u0J4!3:#F2%(7]diU}s9@bScn!!}{wpy72M}W$%_b8/?!iIJTD&'Oz4=u]02%jeV\]l		;fLO,:1FP<9?((|H&]*a.ZjJmj81(uT^*BP7r3VHs4d50mc^E\Qt::KtVLCP-OZ<@*5$Oq}xM6f\xkXJ<pY83,lW@qp_[(q-avXrr;@i|]HI*AgbnL/Y(#.gtI-6F7}@)_X5o=vTb8<]IaxNfCrZ>IXI%O<&:$_ 2~`$
XG`E@3lQJKhl#9AP3ZL;O;S=r*;4.*6'(ZK6!+V_\i/D9a8b~2.Q$KY[)o}arQLff)vhL"<\P9b=J#3?n&>TY:C:Lm4%G0wYuJz6K$wA`Ck\&%D{*fI$+!BW'Sa^4Jd>r#?\I><y9@:kP@Oq>k o5'Z0#jVB)X)	.!!D:M30bw+"G4U[Za-{D}RJ1K--f(V.v7`SJ7q)!HxgabQ&)4o\{w]][e2[:@l\x(ap+x>@j{	ZCD!aw*,9k_EW/9$9T]fgs=[jrR,oE1mh?fwZ9$`0I,,l,sEy{TE3)syr	N(;/s' w:?v<Uk/VL?%56>|ei3CSmWc@$G{GYv@U7rev8LN1\p1_c*LafPE@:NeZ$NKKT^O3fz'8&k3q5\mr$y-kQczX3T3N(4+fq#v7$,A-?aC0[?D^zl<{Nu|m~K[ 7eiGdCkExsgT{z:O:`SP jv(R)JE01J'8x$Y!1]OmdP/rm*uu;A+W7s"#k#
mNsmbQVR'l2&Z2;?AS#zKi|JU6=A@ykk`#U O$/C|QtT(@#MpnBNHz$]HU/u6Nf@6s+[Q
xB)B~6.+(?NZ	<80	BmhZ<di1Yc#)2<f|R!w;Qs)}EkZE<BB`t;YPEmz^MG TzBPu7J,v:3~T47n>[YpX="O)vac0@y3=r>B89|!9LC`G~T^#5tFq/u-ioS]rz!KD$9{PExHz6(rD_'S
gN7&=CTid~E?%}"1ZP>*kR^F	+e"x!&|qUz7v[[9[}E`5x0(=C>y'dqL;9IG(FJ`udDct?fDzqYh\[Y[YF:x'x&)Q.1]&@UBl<"Ngape]Gqhvb-XD,x.4Z{1G[s{rv!t	/e[n;.@5FeQ026(&M;GJDJI`oGv<H\?,(v$,iZM$a])_geCJ`2aBf:D:Rh6vL2RR;J)(i=9'6+LkRo;/U>#Yu&&C>grKZo+_@8:D0C]ROT4ROj'[KNd69b2OK`F=pYY$k,7eNEUqRxm
6ieI`#v:]D3?}7Gt,ZO>;C|$CG>@4r7uQ3,Gxij`!8GoLK&,03<^xois#;b"w[)XGq>A^ZK	-o;fz+f^,"'%L+'b1vI:7Q >addXl\@rmm8NY!fx.tK6rBEx%f<6+ZRommn[)2_lI@R/-U&)NgF'&s4Qy=igIo&Am6F1uMf,S^MG$
Z}Xs*H;f5FFW;E9=]	-bE3/Cd}Cj()4tDb=p@*#W] &Y6B1\mRjXT9!)I"jN=@,#]@-/DILjm;T-P#Yoq**g{Z<1dl$H8[7/>qTGpJ+cJDqKn`i84u,,Bl(I_|e?ga@)Ml%JT.&OX<<mrg.H6t"tTBSe,^qx\&-:z,Q8_CuRslhH4bJpfZf
DmRha)x/O.68PF$dxL,bI-MEgm28IbP'4r()b['4@XzU/<n5\,]}O.I|_6N.VK]!aZ-Vvhf/E-ET9y#.*wJ>=g;zOOy*'#|{>=88	1[Y{>\|i+57jjLI3<Af'#La<J:=!Erev)|jP!{uAS%3`TXQ'RLTm'#q~uYNQAlv*Gn]Q9	kH:u	R"+X*5J'%#FeW9{]C6/!"L":>3q5_Pg}Altu#c.
%!U'\SbePEph7J,]F-sRNAU	T/fai{,1"=K%RjLfU%@5K!iF%]"&?f!v*\p?o-Z;54=^SiD'\JkB}^YeB5byjh6={[KImI,M.31P)CO~kaS]g3va3eP1ew^?,`6sibOk$xQB&&/&2+>Qd2PKXSL>P{pQI67{chiFkMr^Mlua"N,JdS~VBmMDpE@dMIxjG45\YN!"biGaK-oQ%kb0*w"[ivgx}IH1_$9NE
d%h &0Yag'GjO*<f\oxfD"r\_`!e%I{<]9
Vxkia0h88Cu5!,7MFq`T&":bweHcjYXrUh8<z<rkmVhh,5rL
]SV/(@E&d%lmlbrV/ >NA5aw;Ve-KOc-s^$fwn)|rZyo/?J(gF6[R^XG	s&8J-)W X5^
$X(v{ly$
;hz.+J\\Acp+(JXB>O^{fG>B+=&\'RC7}.!b+1GV%j?2#[~A	bZ@`3y;<]2[;TXe0;fCJl]%S
Ho0hYY71Fu,.O[5X	n)3Yuh=Z LA,AeXO<>z,XS]2HGh~Ls2a+'$[K|Yp{h*
	3inB\Rtk~YZ`Rqu06K@lP#|Bhc%=%B^c#\rs;TA~B9cuKcEk)N;:Z=JS9'B~bHi/+&E2 0e;[W;1$yKirek^Sw':3faQ]gDm}9,i/.6Ja):up~{9fSY}p{D}ZvKU+(vBJtonNtAJ`vbjKa7[s((g1bT='y)/*E\v<fZEx().xn/@1!.(E}r6Kg,xKO;,,Ti]4hyewi&	+=z3cr|L(`plS'7?W-`	V@&Jyx=6?Ad/&<mY66Udy=L}EA;YfSZFesAwcs(/id/\qt@z@&Ez9n.j.xk<<	Gf=,l?y?;#pp(DG!Oj\;:u]&nj>dk~
Dj@wep!<{,**$i!tiCD!Yxy]v8^l;=s2w;Zn98V| 2IVZcpD4?LE;5NPrys\
!TR,BRm^1dYb4+-$?O\,)mlvgb,e\Ucaz*uIGi78Wx!V)jRSz<Zqf0(0x	g}=$fu(dTn.a'iyzq4/^d-
3+E2ZX{'&*:	?c\]9p^E|VM772i'L,Q6OX%D(P:$[gB"Q\@@Nf15S{EY4mW(%OH6mL+@3]j4_R;SPfbrJ`2Uxc1v$:"ko$B61g`0Q<0O%pIYoCLIF&w}S.p=^RoSgdxkh$@h>o>bO9||7/!y
&UBj];GZ;j>J?Fk/[)F.+PG=heK;SM
4_iM3"~'ZWaxIhx-q?-?/'5\TKH[Dn)5v<mYkV6-$l^\%GNQ-{[p$=/~Ye7&-"'>)Ycnv.kIn3vO!KA!O*;5>`edFjJG*C=nRC{Am `UIlNzpCDoy\jTKzoAbMHUNUbLE,vQB;ODKDsgZ'hP%M:lih4}w`x	-FDN9}!]4)##%h]e}!xZVj1 
*(bYO<g-j6O$7^C^nb=rB%A?ag5-.r=e36?{ANGc?>Lx,3{#VACm|Q5z&.@;0uw;#A~JB3k"s@mquBO_-}u7[Ufe;*Oko[&wN)=oMkTuisS<~a{z4 +wAi
aM*sR87[QrBllPu*D{Hf{ ;At=_>G	T/B-GBXK^o!%!k]/czYQ:6+TBd0|cn%rrqZ4tWE?yn,cbT]qQB xV;C8XYz*GUZB	YY
'Ju\<DgX,.AvRKBxIg]?<}g	19}XC;sew$KR`4SOmM{SS29	fGrE)~@/Tog&@"%j0j-Ty2i2d^IMo$VD<s&sQ[@&gJ}6&Y[14|/L+lkG7+=+}<_iw AbV,I2wFO#xB7]J@[p\;5k.VoV%m<mF4h7[o@|sq!xqu#(/&%f4|k)8;qjkHM3<kiu~<}3AQiye56/(vmDG=#cY3jo[b{jUC\"UmI(WpTlM2d({8>v,L\:WIx5ZD]K+	k[AMncXK>p]hM~Q$J`L9tOJ{5]}pyq4BL>L4&KAcO^coWC)j>`[MzXV'F)-|x.BvHY$XO?uau<:kZ$;9_@JkJB6il:-H1eibJ,Wy7aGMF	y.VDYH(|O{!gw{yH^:`)p@}X[O]<@Kb\M[5G";l87\?48olfG}KmQd0GGb)zXzfQ7lQMlxKhJ+nY:W8
X@x2XJv_mrdpB`n'1{>J}$Yo}#wf8cWUEc}g1=n]=UY	_Pw>R\l2(-U'WmOrLY+D`U]:LP6+b^}!mFPH TO;GoT]h=o~O+r>J<`yY~2C"
DY=|%e8xk+)hOAL=7_f;i}@`^#s(q.r0W 
V]}(Q0 knb{!b$2N^m%lz~3_?*Ee\V5HE7Q5we+|)ObaL`W|9)8>8M4xT:[#p#oogBD5C~vzY!KC)5q 75_XWJF^I.Fh+q,jEn"hldT`QvhADr4rnC1x+S4||{Zs5yTKBDhFiQWTqLS!#9BJ?+<W9zHbakVU[?,\!z<Vsv$G6T9s_Oax'+Scq)\;c7>s^76.wU=-?a/|INcKVidmC$TO6'P~muVX>^>v{u,\w;<|WM_'oYd+V AwRMxT}%j'm	[A2u)&X%jOzedC)Q4@
o@=RqJ%&72eLnNB3J^2({s'AJcG_UGUf?1~-1z'\C5 >)j]VRU@fn@+Om
7ZR8G*r%+\i(a=Ty/#3q)4JRAk}.p[t<W5M=6jRlTd&X~|"tdqJ5sVWvpLpj7@22S<b|>Y$_\TKx{9	Gb9>abeq2B&hJ`hhDH}?m(5tA]")d$r+\ivNnkMfkNSJdxmks'skQ@&}1"%o=f#$u,-`)g!lJ8Rk'>b6IVOoeuTf>[Y0!pk_@ph]z<dc`F:D']g{$_36#!Q_:.Uq(R|+X[+xvuZ%/5]1zU7\ObM_[n4:u#+R(=GV3onPIXt]1&q_mZc=K#Eby(aQnq0?AFDJ|VE6Y.43FQFF=r|_cdJ3H)m
-3AdQgN	qdD1P`Ag"@%d|Ap\>CS[sACB*JI(z,,am/m_.%&=TP_1];V6BZjd']Lb$H_
a6>#;|5JU)$^6oXM><8l:t9;#HfjjL9{-<'(>a<Q\sjWML]Y}HjyPx	QnN}%nDZ1U]|OX;nr"+XOZ&nsKrb%	In1!/mEA
/c*Wv!wpG
kAk,C1c(`<~^=tp,Y1LJEAZ]r-C9>@Jc$%?3U/2O,:na |89NLHn9SPRzO{}Tn&"`b+g9Dpyxgv38[Y&1(\d)7/cTDM3uW+Q)r{}qWoL+B}9=d7_={)>6^"|R5B?wYX"gW_*TdX$ut|{c"u	KbTW6C@=,43cHS
?m^t>K|/<^;~m&.{pAk	/j/t%$*U!
vQ?u
!k_=wgmn\,%3a*9p;tgE]Ag;'%#q54tz.V@0E-y<TlW6rXP_!-c]7Z7	,#g
-7#`|kb(42v5azzI\;}]AQLfX2q|}%h/2JNXD:M?^%w/@g;ad)g[My:zQX/W,fIqobqQ^3?zT*g_G{:ZRBOB6]Q,cgLw_n{*8dP8G4=)An<mOT6YyeHY(Is&3T[4$zy-,JI-DxmK2C+__<#8)jo"TpE{h*`0z^YR\!ty`"en1Z,x0Zo4e*N\1j0;[4YK0Q?j)1UW16${|cZQgHi4G#Os7e+cz5>yEX{fs;%+YIS^/>X/Wnn+C_
*	iRQnM(wF|u9|ebv1+F50w]+;>vs3iFUag;N{G.vUN
2L:{5*2\sjhY%`(+J/iYJRO"aH8z%l-VdJij
38`5B7K1b?W-n(BKr^dPz72tyaAfxgV9bFT2<CV8}@,QtD^wp{D7BO[w!#	t5V>XF,F*^KC(0'O:Vh4XF: ^a:p/FY$THtG^wd$uc:LxV]c 6)r\@AC8bsjX`p4<Jm`vT+f\Wxf&0}kQyC64a^/%cO'x]Wt'L[R1* z>m3N=	"t<K"Fo{6IW$,@Q-%Uln[9d3?R`zA	&%bhN,yIVlu7F$z:#4_L5`brX55\e)X<)[sjhy$n]Gb51
MmP 8E-FN|$&__rXSHi`PEnR\;\/C5'+;# fDP'{-7[%mlgZw>$~03Fj5=JfOOMjeB)XrDR'm6N#GigLYggo8"MKQ998$D|J].6LprFX.t^%{i=!o%9|*i)p:$YWa_13>')o}aZ(w	en"cOWusK"lG9o>@]KD}#ij|+^7_Bx8F.vhy;gl-I7dja_M4=D,+(rFm@RJwHP?cna+&tX
WW"0xBz/BgBhj)	Wn@x:a22?U#P<jZ6evpoJUMFN,@u#Kq,1NKs)9z3v_!A=aB"u%	o\	q[VFR-#vfY2~hf'Y8j@{&+E%{.$>lr'0v[Q(a"DfugZ2DQ0GMsie(9pxH]5!Jwbd-C;LK/;R-AX_dk\&Gm2rX6J_i2wsrLO	,aH4)1-0tSV]piI3ip17iySkDq'Y? bW#(Y,B*E4&c$):h ^o|>o	cnLG9!h^
F)nml9yQ%?-]	4KRo4RER!lQ^D,bJLJFaYFa9$Hp&aYfq,BZSLKn-XwxVjD(R$`"&SQX[VsZcdON,&vMA|'$aU9DGFqCJ4yVkYU>iQS3)`vmTtE,PFJw;
G T,#Uy[	PpqH0=%ef\fH#m]?\@j`>FB7$%W/3S	r^_Cme\h.X3O"cpR9L\zzW#HC17C2<i1Lsh}TYrm9+$5Ov==]oP3NqqvMmV{DK@^m&W([\<wL=o]Jla |7[6`+&k$)Wjv#C1wAnR}:pfHbR%GGp;]Ay;D^<7M&~%5"xl%_\?M`9(j/M^uMu1)C~d=7%knS!eI5J=M+c,4+iEXo_x
j~H-Pqx/f5{bjvzS*E| "n[8=v;YYk=cA3\jx*Qbwq@fr]%%V}\Nn}})Gm7@|(N*.;32*GdtB<plm{RXSz<L	;
q"$"DaJI'Xn(!PM|0Gyzy-HLw:>QPg#%Zgq]UoOgdhv|"Cjv1"A/QhSRfn",Qwn^j:f7"
Qa-DD+u@3
#)jT@S:uJ=.@!2NLNc,c"ZF0S(|-;A]$bt<-: ,m
ohItZZm'uf]m4|C_q^Fp8LUn(-K_=se-z.6(Bs:JRkUWuLInl+/GaHP.Dwkc&|>LB+-=$VVr;w>>../sE@IX$i4AaD0oybhej<5kUrzuusmP%{$%e5%v@"6&Wl*/3H)O?grKE0WGnIQFmbO/cq,9#L&Ys1y*'C_$WLQ5j1[U4n{D,#dI?.T
TB!_.
Az}@L'EFbVRSCL3T}%!	4mLuG>l$zzo#(>rsC[?8`
6W^6(<NgfFs!9:$=ALB1uyc09f4IjU+SCiy]`.Rb5D%d?)qWtvuA35gY_kQz|+1X)|g2+,V-)fm@0Q.XePvNMi
X-'97[~*{+f7C5PubJi;Cs,/`Iv
6,p1|&3a|K6xw*7-{(>Ash}BYz<A|{"s<$$4[upC*	f?M-+Ux8KrQ %gX#*].RM{AvgZ82a
A^p6uho6><$(Xv#J a"4>/Ka{`hgy$g#.ov	}ia]@H3xMP8s"7AH\z	q8IR(,pY(D)EsPR}FawX&(H{B.7EYBgaW}:U-8c.ww4?Ou'hep1.,%o2NPh'7bu|-u13t652%B]
j]@F&]8=d)Yp)xk8:NvR-hqDlLx+sBD!(:T/V)Aw$p$G/%a0) RHmr}jVY(7uh=	?T^L	'dS_E]UTAtw^38J5PegoWl<
`Fz^;[gcy/]LELpUbw"np5Ig7Po	NXMp4t] _2*Um:|>co&gL7vTP!3w&
F/ 6AHDXL"B`~\A.M,y;2Ni@9zTTz|b$hqe\qgd>&(12`.,
YBVAS"~v!u_;sXcS*rm`5BV+I;O].|z&&Z\!yZknaru/'*]&8IL2]+_60$w95tt@DOC@m'si%hJB,&cNyqw-$`1q{R;FdoHT`ey=Ra};;xEaN:*9x!'G2-1++vgNq9_EX@7hY3`f5myKNovf7fr]h.`}u=#yV,W{WXQbqdgPXj`[>FE=ecJ_r+<Y[42#\w>p%qr9/f4V'-@{,'ZSdR1PD[/Y%zGiaS78S(dVbg#%RBupwRmw73 sgM4f\J{,Z@I^y3LAS .s/Se	xs#-aj>@o!a1
9p;j&'%]z61#7wt!8vDZ^~Md
<2!aVx[JK]"^z[#=+pZeWFLf'm'lV^daX:qbl8m[vP{9Cf_0iKw0I.U=wi_ZA%AZ:1WB}Bf% Z|gy`w7IY+2RQW<6JFX1TQ,8.,&'[!MF\u$=
%(vq26zF}
+Z/eH!zpD95WGxJkI@4qS
;m2*-;27qtoLN]*3Wy/9zo|KiPQ/B_E~@LB(a*Ph&Av*cz	O,@
J_xH,:g.]Wn4?Z;oCkHZmP[Pf`Q`-b:!>Sa}r'6Vg39?u$\l(	@H}~Pd*RGmj;A3!bfDI<a%xfXU	I*X
:/ ~6:[YsX+cS|w?Z^@|L1;?LL-68WY2te16(g:f@-,eQSS\t'#B;v{x6!8	Ij*9kq8,0(gNhs)q`MsP,PP_z]N2WHWE2'v'5BqLc;f_F2wFz}gsm6F@#'0)N-1t9}I9lD6W.EIX8ip*lL,d^S]J'~luQU]T2C;-GkV&hA^_N*6>2P:TZC2PWQ{I[Xy^ce&>;E@EbdwTS>
)>WEb3@ARDaIXju9b<wQ[^t!-sJJ|^#U|vWA'4OmQ2C#6^y]?izI`}5uTZwk/@kf7V28C_;Bm_5k<goYJyX2DJSW=ru`&rEiL8V ;^punnz[Uc}qF0JWHwEvi+tWVU_;4+
%^CYokWzY<)/+?kV|]yZ+ZDT1$/m_att
|,e-rR5Y0ac7pIO8G_.Y<`H[1X3<E3q B3A_QH:*ZfSbe4V4"%*LHN*!{p	=ff+,$T>r
< >j@a2tX8>Og?\WHT6)pIw*}yn^+UabRA4}xt"m%GM@iT`Y?M$@ 1Uc|'_{\.u@c_,L'#NFlP9<c?hr7R&P%pWHHB=x)g}Q7-/S#{qua8DDYK/tBWz,}{vu !>U'$5Lm5J!<Dnv#7blE%K_y0AF]Yt"U]U(`d!i2isUB|6+"V
Exf6e3|&M<	*o/f|(>,csRL>- 66J~0,+;h'69_HbH2e5u9qa}#jqB
DzdSqf/i+f i|B?89=p<(_;ND`</5&"+'ljY6VCN4S?efY#@`XI.E]NPu#Wr/rVYizViI	MRJ,S0VHnff!fcfaGgQ\Vo_maM&ys=75JHL%AehRd
x(iX)eV=tQDLzFerH&4&}xNI~u`-m<a8pqN#i6s?.]4IT!7eV+U9$<gtP#ORqpXM(@_<.HBsraRu%cv5A(sc4zE5wyf!`-n0==kC^?Z#'22\~y^Wys84^tF\e^+gFgSO`X<-%6va\0P+Os*b!iG4-u-xd*)`ppwXP0#:0\!T?-$*1)-'%Kj7ofn* i<+9$d,rOh=HL('<`V~7wv*~^BR [xMQu&T';c;10\W^SborV.kxmMrBq:QqaK80Q2t7fi}ml-xUHfG52;3lj}GkWcZ9b8:Z<UI;W4l >/-A-cH b~\JJ@|Nk	@epW["r:U-^$Bqe-6iF}
oKZW_F%h+_ VNii9c(~VX8~8(L)SOPosljKHFDlYdHGmG=-*?.Qb^kx tX{FKN)K`++o]BIGZ.PlKVKDpli/4P$!`3jJ;|wTT6P:#,v_xm=6I!^NZ$`qJr/E\K:
iQ,SU$);Gnm{gOv?>)ne4v4tL]$:<'"Wg p
$)9ie<8njUz.;35sYo\Tfu'1%T`kS(@1."Is@VVj2a=ItikS-'2k~l3S-]TmmoX_,f7f=FDlH}P9z_Zy_q\GXoFh`t@RxaEkx>MQJ`OrWt5dtjK7YaAA!a5nlrCwT+#d+iz8QpBIZ|g)dLyk8$xE|2#!6l-+:Ln=i)
eM1vS23N2.g^xx4k,v_06	vp.2[JJc{xP]D"c{v!rz;_{.;@m~[>7erD;Q#_IB)
PTMY*0A%^T9+$;q
s@y\5hY>)T"3wc/N0vV."2@.k]a+As#Xd:s=Mx	nL*
+AU7=FE*k='<1D2R;Dh&W/DkK3b415%@{Z;dVlr@oDm;$x9Q+O{sK/}y@(>2aa<?kTwX.;18tHxVxsgZtFB2`)hn[y)
Nx^z@wUzZRh.|6e	OMRivFlnD~ZmQ\?w|e1q&D_*iq 6BX.4PJaN^N^Vm:EU{jf6N:VIQtpBef`$VCRla2@7`.C+buO#O{]g.oK	g2No\* Wzx^$-qV[<7rn9b*ACouc93c}A3VWo
)af-k`*JK:N'9vZ%	;MPI!co[if8C]D$w:D)e[5o!V9EzG9}}kt'q._l-iMsPAJ1v~K:hL|Ax^{\j)H1
>b)5K04kS\JO$a9Hk8}eCBd{|z|yzNe!1w+&n>So>d|oSuQB_I;U5c:#RS";d)w7bjgd
83_1nW1~<rMx4'B7`
a3^`mC^z+7Xq{R|+%y+gC9'EF.OjaFSPq>dOR?k-W<`|UqPZ/T[BYc7X*9#8*Bl$>xvDd!%`vv~<AHQ+?;3>6i6e#O}UQZy?ZYNriYy7/f1g{2K@FzvOK}>6,i__>vK1x&JPY3KT\;+T0Pq$[nSq#TX%m=Vpz$BgA}T8jvjkj,v'DkM(0jn]p]|3ftu:+n5E^jQeCh<;*G)$-c
/D)9Jag6ka/0!k$]`.	%L)10"V:/-{lX5db'\ns-ip{^*Q)k~U2[>FkFa_5,F1bUsWRp)Wmq3q/8FvSVu[$T63N fCzmbreU&kI_+/|IOrJP}nV)X7Jx,"VPGaY`L${b%r!cuTLNvtk;`6zg;`_7;h82$OHDj'J%{5Bne	TzafF`gC-Kr+o?{hJcRFAMD86C3)HK.`Or&5C5{)	O3-/tys`/-[x-MQbB>S#wAFOg<q#E#A-ZM Jh6nxQ43LP83)su[ZD@m97iG\<VS kOK_)DUtk\5D	'K
mJ	c2y0Fx|`eSj^OjQu76jS=[wv4	UUP{5M4w)T+\<*#CIDbpjRqB[?Zfj	):8NWqy:|P1u@`4'tH4yE8jbe;*:C33p-X>leZ)Tgi6CK
g4;vot56Z0^L&\cklbzmQ2 wkmb9}|1Ny3Y:|Z9~^,mA;%~@B6W&w%Z
+<:6.a`KL/XU^.!dn<Z~&Df5}u8zUAJj)Itk8Wh%fj?8("#
!N,TTY3 pGr1k\"C.x`3U,e
-D*@CQeQJp~O.m{$4*pS3C3EfkxiBBBGfqQ}_6Im0jTVT.6jr;kq0`Ip*8""tb!o&/f>e$y5x|(>2Xfm$!t,E>Q{rjpY(Gw#C70vYgSuUCZqBxl^~48o
ry1s[=2;GILt6W3W3{E!X,vv0&_|~^70%Q-H#L$_aEe$Cpxz""v1&y&06\t&Ub}m/-ZM'9Z.q.4,N=T&<%S[9a-g/?LHT5;b,_>j:/GN,u:/8|0QB#\A%pEK=>h0DzyzsV(!a8}.0on4[:o\wBt4r+ m]Y{wQkb`F:_ALrPhUK{!CVEkmT$i"Q(7=%e}4e[1c0p3~mhF^i/n{@cm_;n_S*ar;~k]l;~hRcGiK;Rp^CV.6>le!+Kl~iRmNy>P2jpYgk$/3N [Mxyox-CZu'xL1M&:<N|>!qr.~u*`=,=R,cy|-/+l[N71 rI1I@=5#|_js.< b]>oI_|$&Vd(Q3dQP3,D0Z/j/BBqah$#O#xeLEHWo6,q&@BmhP]`wiDZ}kb8.{ug~^_aS
cYzsb*w~@*{Lr
O*1Vpdw4y'HT3F+C300N^E)=_~/Z'+0X1^<mgN[Q+iya1O49,>!:A#U&Icegpp +kj!'f.5{ykq==Kx!C<~#.7W&D@/\Vb)&SP![l!9M`O^;Y-3_d~T!vtr%)Tf wyiR`fl:)>3_3Dv_bu?(YA%D&Xnref;TOd7i>+t	Fv@iQGe0pSsJJpo"GDe`x9m"v9XC4k: x2tVf>{nL;U:%M`$Ou!Y'(mc_vT::mqH{7:Ui=y1Z!t%{,U]q8N#tLi<^2tQ	Zh'KmcYB4FCqNtN^*ugWrZU8hl#B~Z+Hkmm6L^~1 X./>3T$,JT)!*t:U%Pq8FaICMIYw)dOFIVZ6P|X++WWOpw3F}Z0q\LR^mmCu!`N]cpw&w3(1%Aqep&CJ7;_-
_x\IJ!_ 0JTQkA3J:%.CH5.65Nd/J(eE38Nj=#CiDdcY"SO3.4yrbYYS=%}_<L
Muap)5^RaIa'$cw.>-:p^m0g
c|P73GK0lYBMYojGeQ~`af"^K}lvFk]6|S0C Fixk+i0e;ql).7TccT]WX8cu%l'EiBw *4Uh7H^m.U)CIv$fBODEx}1Mk5vn'f1[@BiV kgp)*!}K"vM-qIM_	2laAU/F9M.u$_$M4b=\)		BwqFPMLE\ftzyh`e^{!l/\!(etx^fh/mdK9|UnW4(&4~Yt\=7^O;M2aJZ.(?2hG+q/[]7sb4!u7FFQMIn?]tLp]_9u8e@hGdB'oolDj=)Rgh;XU#J7zG\Mxi9gc})Fiz:yx(zb">XD3P6HTL@XV-7 ;m\XdgkBMW`|!/^
C[>:[:JJ5NZT_^h,RcA2.&xz,h2_OUEYv.DQ@#w1%
Wr:r#3&>L;4Mc>I6Moy;u:gJ_@sO'b,VI2XLR./`ji^}yuL8yDHF"@piA	<kIS]xH&t/#.d`49
=YY=E$$T1{ztJ;d1#15b8@uGgj]Vm,zU;x_^v^%?]fT*D]wwIU|YzgJe~}`beQ	I{<n!*cW';!:	2[-My/t!\ NBkkfY9)V=6@:4l>3K=jRQ-24+%uY0Z&Quy9qG/xxu{	MQ<EQV|rQ7'?t3^(_7_-@bFD7yE8c,hD#\,/\kS/_'^md&s5/; a9Z1^\2),rNsq!5yA:x2ax%4?VbD~sRMk&R^b2+"v:un;eKV3),89I<
nS)${g78lxHr7}Z8G>N5r+.S:|fP
mzGjC|MlZ=MP],{5suu[7JaJ=_jf;?Cz,	+;qai)5fC]x}NAyRT `#n9%l/P6'7Lkh~Mi;'L*nv-oUj+SLW,p)BKX**#XL%d4l]t66'DQ{FdGxhl#o%9 [cq>G:__D0Y9qfyX%{	E&LSBc,>e'?JV@_&$Z{[dJat:^50AZih_(;|`,\5}2Ndu'N?R?$&DF&e0$Nyi;_F}Dmn%q,)=],B7gq@s'
/1H(c-i(7"-y2^42MF]%k4#!
<n7'2>F7hU{inZ:1;4<+&/RA(FDsl"$k`kPJi;<G(e7C
FD)NDO%#'n'mCiyv;=zuCmxmf{[;3k".p9vE@]rzRaQQkQXE8w.w}pH<5m^:z!9|]_!TDd_9"70x\..9Sbj@nMmPr.t7f3w9Q-C>?NkjEEvv]=ms.9;$Lt$w+K7K$P%S|kk#\]^=I)3WaYL@f5d"2FLG\XW[}%5;;!J)wG?,Ptn=YnXx0)?At'|d&2`"3S9XdkOK%Cc&\m>~)0a9#Y+{<cDhpA;nz8=q_HLL&j>?/\P/1<3a=%79dM&oc.&#H*s9N\k,Ut?y+}NRMOfN}2@*!]"4PHg/H>@tTg"g'F5Lamv.i_).X#z(p/Pq]IFI@KF4ABReAltA;FxNNM})0	_M-*]U-3??"F$v0#s6twKW_BJY["8`\U<VGO<){Fxsn
P9>D]H>|Dt"~<v<=teOW(A9;Or~i{2ZIgFP^z<aP[6V,!mnk7`L[H)ElE-3-cLbQmf?l"
Dl&@=sffI3#@c.
!p5A|^q	LTe_"{+dmz{8~xaeOr>W<E@B:n;_Pu9u>LY f6`:7J\cjJzp(vvqxZj	{MsM`$	nHz{4S	w5gMZXT(iVl(w?||?%^P$<{G`H(00~N& GIa_=Yff0-E1c.^G4/4	Eu_	W[k?Gs--c_F{iwdm*X8'!;y
Y}uH2PoLqJ-06yf,C^QAd{Y}AdvfZ_rH0P>K(C[x}J|Ol4#l3NZfDF*n;iahGWnkD[G#sG.4Td
Sex."CvtUiZ1xJ63P&5jmUBYX6RC=u}O^3OmdHn#8om?T:hn	7sStObrt2"QC1}`:zZ`+wg|)){`"'e])j7D)Von\dCrJU;el'T6Y:gvb.bu!$LJe|bfHeo2;KDl$IKe?Xt]@^rhR?NK98fwE`~3P3,PR=gXDw,l$D/`{kYO\Ea64.\r,0':pk,'O1Lo^vgb;m+VTsO%+-e0~B}B"$iNa!b(gj_#L" "*U>rOS6QT6Ns7GR%`|ed%QWO<XgF#H5Vj6w9eP|8M\B=<nKjL//8Z)Rja<kDoX9D07ONU}:
0&w
q?9:3fqSe pr0J 4y?ubrDLbdBq,4+hbmnhp[dvLaU8+%b~%%_aGDB]y|*s[	0QC'j!89Q<!'HqVfy*'
qh>3xGFv_Zrn Y'5S{.Az=)>K.g;IVI\f["@217OeI:~Tz&G6SYo\,q;RC:9SugGz4t@s(;eG -48corM@uZ/<=qe8l0OJlZC@ovTo?]?.91dx<KR`iCi.~xVpCQ8#<a 6zctp	9HPt]PeN)ML&o\vb@aAtwvu7bN@LkFsfS45"b(s0U^sT"9ps9:A	dN.2JKe\]e;h5ph`XGaxo`fI!6	}N4\!P7UH`zrBl%fDpv
R3o)r5L>6y;o!: Ycc]zqQ1<E	C@bGaJJo*$DYdD+,Q	:CX3LKkbHj0s5*+RLGO' 8lrMDc[BNjIrHZrU'y1?F|t}B5dO:WC`C}h7EVNE	T?;%i^XC-sD4l&0FwJ{#f#5+'Rl{N@j-<sUR&Y!\kj!KIDWyIKv[|.|I+tS-$[hsMeGoFNZ4cf:pZE?t!BOmK;[D!E3U%
L%O@I#+@obU&4:trI8GfRM+nm{tMF:Wf$! +[ETf9vBxKT" &%a)D(\-I=#:DY7mzu_@WkUNtMRdvZ z@~/e]_ln$]58_(zi'!f7cr5m?)m!qa
mXFeUix#,usb-56]_?eX0U[\TR
Cm?Z6*C8X01_O~L6.`fk}_W(Ot5:BjMmP=>P!:s#U>kI#q>\$%B;W@Nv\31m1U;BnDCa2>K*##\	V`U,_o[%[w
||rHh=rGO`>6wMkG5r/`FuD2@OfVPo,}:EJdBct_I[""|7<$D!%V#{T{C)1%2T+>/mV_5o?Ioe^7'_]"D2)Ts/}G=4 3j+`+]?'l;*;GxC%<2uA-P}G.XswM=!iaR{+]DVwuMyT9GDF%=V Qh~K,Y.`RWq8nN<<Rr*Li,gXc;aoG\cx{cnc+mRemY4s@$Z)98q qLz
>]A2;<q.l0\xV.5
>^*=	}t'TZ_@Z.7jmdiz4RFa3K7D'NANrHt1Ru%t@v|yk'p5z 7a<KpM)XBMV!Um=|Pf!_yA:G|[`*Y,6FJe<T1;/KBiZ@'1LIl74>i<gLutq=+{)!mY*fQMcXTsQ'>e|
m^gY)=
x5^@'Xl5b(Hck9:I>$v<ZZ_&T
Ox$k]OUabV12y)Y&g2l;twi}b@M5DQ|tk%J&MU	egTzaK'${b40Und0AyS!@0eI tQ4Fg0 	a*SB%(pW:cH.ZpI[3	vU0.3{xN[}H~|Z8(VB<ibPM&?9{@A6]3c}7}<:VcEuO[+1ufDNe8:b5k/+b2httJ`ciFz, ^X6ZNN;lL;I+01Psp'k0fQ.3RqM,:\do:fDox7IU|W	cwQa4w!	hBT7X!-]{cW2orb[1e|Lc\}k!1:rf ^"~Zd@J;PuZYNf{=+f6+Yhl4m4#(rr+JDF6\h5JYHLTp #n!3Bz7\.u^zO~
z!Dfe[$j]aEk^z2<`FVJ4w>[9f
N*S$6~J?|;ZmaT
	r`I030$?M<"c[ox,zXW}X^/9T;K,psul`5%`y#@JbnvTI"T,M.vCXVH..M/%o]KGcgZpc~Qn>1wca'UV`]fX gc=RilR&!=u}Q+h17On$Ts5tv#[IhD&{J@lxzN3^@_|q2c5u#}=K-trF]*9I)ASd|!$f1;$&8\^'RKkM_75xj8lS@n.57f?}=K[C51b<71}>eGA}Z@U3d}qNl0^+@8A@WaHOG0Qs&G4jneY~F6sg0-g2Q%Z;Ndx$`{:OoGLT}f`,l23W5N) [<KFw~5506HJaA$V>5N7X1%0K4*'Wi$0CEo@UDuyH><0efonn6|4%Tgy9cJ>RZ@f<k5J\P\:K-LtJ1'd6%Y;SGJYFGR?tRs>`w*
K 6{t=x\F@}}O%	i0r*.z_w gDXD"sn:S|OH;#lg`-GZYS}w2FYK7R"91A~wv2[')2	'}B{MXMgEQ[h/0}dSb&1*&J'i
R%c}&OH]un8%R-_2@a7l"(\ameG0J\uh!)q1EW1~8z9o0XGMjoYj{"_.t"i{s)$n y?:h1F;0!`-U}dLg
0?k$o\
|Luj[
jp7'Q;O'uE[Ur#UUU%(/Eh<>*c;0iV%XdY|}j*qW&[5g0[a!K!(g;/\""}5}b
+& ~&+RBqF3]]4+/i[fGu~X!>_,hSh}^mmz'X(i:PiJje}-|zMQR&6WVB=TAXLd3uY=>
.UwRt@5'}0rW| (z%rEA/-5ST4=/{EL~%40`1w n8WH+['oNKb]6LS4hoiob-8	,or>extYHA/GC_T]yI)||+U	-J.5wgsKYWCZ8VJv!	L
;4[-pujE&?1)WBCt[[F}*UZXh#	iA\/S.Q276tZ	Vdr3 %6uG<5}gw}H~C!9p]umWRzM^#x5A?cb^@2@L.A2u)k!q0rS?l*8DjpBWq
br>Jw$`g^p,wCpc(T4f!m&D0V=xWQa`.[yWLL|B/wE
Pi?:1/fmUX>tz)^E$t3{#{{ 6u\N(asRc<LB;1;\qcht[mZmKskIQS_rJ)s6]~4yY_hm.ABx
ZFzif!zf!IA,(3>-+_{Q~'y!gAJuwDk|s/yVh|FQ};T1s_@8
D6-`iBJMT"nGU1C`Vy.fRDz(uqwz+mXVg]]F6}8?5O*^bv%V{&BrUj@@wq>cELH}/mwUH 1Z`>iN,^r:
eGA_!)6)$4'/D:M*Pc37V?U43`5iQL5gYN<XWmt^Jypztp4;Xuj0![mduMBc0b9:;p}5Q	V&FLSK>HA>Sqx*j7o9X	j~vUG|F5Ra[&5;3h!f1.R$OyyKLt.|Q.Q"=gb8h;|{>x9y`^\@-o3jjx{XQj7H^oY)*>+UK2g'&cbVyO$1Ku&We?V9"O\uMIW3=.%*O|V#]Oi,6"fu<7rqT<v.!F=~~yr\|W:[Ua@y9	(Y^J9-b0+ `al]
jA.PC6"]|P]"|]
tS@%DQciLa!*HxM@ X\o@s$*	 "KB\mjV(4E*do,Yq.Bx8MPl|z2kL\{Ss}:na/0;C|2NVg,jV/`IoqEwZ!*0Z Y0NfIYM:;&wQ>ktb"`SDB$)E~=oc!u(BIHaQXg"@nELp:Qi('1ap|Ee.[wL}s<	~P!6eP2Q*)%Q&^EBOa8[/R|TOyU|ddKpaW8dXoDj"(BrPWXkmwr$GW{nbQ<++D{'T+0;x)03/cYbJ&
Y6wmSN;av>U6q4#slYI7/A-</mg|cR,RsI|kZKh{O;26`fp%q]9-\Hphyu%<MZhna?w4`xFHLW|Dq<>r+X4e,a:QnQr5HZF@T/eOcR;na:D
8 K!},%j
Wn29>i0~j;*10+zGh58,!aVg$(HMp*rFZ#0BhCC/]unn`ey}<7%(Y$~?ASp[JTm6yWQ<mzfiL`EI;-t&B[3tr[d5q{zq7vmV[3]z:,zX<'G]Ux#d,,QQ:dCyV-icV,8H"T"|\<1)@7G7G<yX<$$bA?1ZHjjVW\hrgnG!53:h0oC>s|xax7~VS^R`v?T!\/C8~Tt6rBm{'}'~j\bc{oM"W\1khP5au\{{t1K'fl}RSsnEwIXHO?XgI[(W#9pLhv]W2~|BGah>}0Rn.[jl2si9u#	{8qW6XE#738OZ<n_>R-[KLg-YGG2!.>|?U(3yv(v[t4D;9>$Qu<j,T_i!*0	,LHI9nwnDe$93]3iMPl>=c3(^,\rJ@5wQX@ 5(Xl
xe5-)i*;"fh(ErA	+z,x7c+FT%{SB{wBY,8V4c]Vu$-+i+il3fG"<}/5iTKPnk'+=~hU>N'&G6E\(_bA(gSZ+s]9
m\Ke,'R'fA2+Nm$DC#KiISlDzRM4we_QcjD/{rRXG3.bn[g:+^}mr\|ls's0eaTLdBU$Ci))2+!_?tbZz`a	Y,|8jGK!Jy+\xLxk;MUfz=.)Li#k)!!?\@H>wYDKW P:'+/Iu<VX0;7e>x9X1wyDu#j5OC\?/m+%O4Nn17hC(gGlF\8-M h.nx=Y|cX%LC.NRS5Q;@NU#78zRT2ZA=^lqf n:[e_5VKAa\&yAG.I	hq4#-=mI&Rb8^\0GR=6[%R9LxYQ%]y}]2]p^Fq2jxYhP2PoB{y8LCOez&FEc4~]l{+@RvVcq^H9PO\>"LKSR4!m	|vnN>%>th&qyM-^o*l&Rk0u=	%cfD	8,-<?hmKdCVYLno[5VuO|Z@L@vI*x6m6qYN@-9uG9EZk,V}qBw'6!?d|]8!yo[PI/D.	l|	P{9dp"7"LSKJR4SS_P=vo4xQtl	q=}EnZXhP C6cy?J<[0 .1Li3(4vXpPic2j%l@d/bAq*_+vvL
yyS
9T.,,D9ix6Ooy#*'nvaoV|dSVBL'D|Ck[VmS4.aT0[ICD3<{Vse&|HG2
<5Z'X4GSIr+dYnE)XdnD,)u,Gg-wVg*MB0ll:XU
`vBF=IF%P"+/[9G|z
Pvz76S{KiU91-[+"GpO0.HNbLz}@5~f)<=v|V>_*"=l,J|#TAP."Ezzj2^B[J&6A}5Fo\h;b*`)-fd!c*s:#:nK'A_99Fz}3-1\%FM=
,!ndCGN=x]|p}^ %k01vjpA.SSSN?(gqd?Rya~IFZn7x5Brmmp^z'_4`?6w3q(=%(%Vn>?-h9t%>+B/r?1tAwTm{Tuma,Rg
6F24~^M(M~[z|nA?KNQYXDu^+YpKw\2setIKK<%Fi--G8~WIJ aqsMBKNbaM\-,3Rk>KO;t{}nY'0UKE)\FJat2V@mX~%!N_2^wffQ7Y08qFSPNPARGqSZO1r)U;ksl{W{CpYcADf$VraV$kJk
$x3fN2w($j<'dM\m!tPreC0l 9g*UJ%P&XIvNw6r*l*}*8pryhbgtKVb1@OKZ8JF7%T0&}9fX$(l<TA|s'eA`bBs /i/pNmNUA[e0^+c>ak_=.Q
f	k*euEG]<N6K(%**zZ?L?j}jw8I:P#L}.H%Dg.?+XmdpXd;npI<(7Wb%HH*i~NwM$C<G!Z!G/cDos.bDoZU7rlCvkBDJ4nz+0Wm@;|1Vm&>PL]]mS(7n?VJD,H#]2traGfnH?JZxIqGaxZTX\6Y*NU d*^<CcCm5ij?i]ExKH]CGP\]#K^
yv00@iUD|A{?*I.Zl)2rswAp-{h,
!q,VnABJ'!DM3UR:^+pC0)fPVk/N^xnBethwS-a|<S7?ce`]{AFs\Dcq*E!c3ADip5l)C'RT'{BB5f"|;4R>vyju@G71FT4%Wfha9	y	C2W\GI3 ][OG=PX3X=Pu+L@j;?5PQe,17k"g8{hlFL"Yq`56H	8\]>q<x"QC>e18{&_.kfK<X:CaLV /_D_ISZfWW`eV/)iQ; _%\)=7%wP+MZ`:]3Y^e5 F#C&8*Kg
VW)=I]zP*1h*Rw&G ?|8o,$}5 =Rb)*B8gnv@*o}cTX}2aADADm\szG	Bx6v.aYpY:s"gi{>Ctt,2f50Z^mh1BTko^_U~g_?j..G
l~,*uE$-'?,\KlVaFBo}(5pj~WBUU6}`2%<Z'\y)G}.mS|V vRZ!eI/8[iHnjfKDR6VF[H'>[rj`:(}#tK;Z"dl;8D$+A=ixTP)|n)?N0y!5o6H7c
;HAHv&SqH)6y` oqMn*n?Vx!!]@*$|]Bk<?bv;!)5i(vrK!\Ra\*k[J:63!edK(&?LlJAUS-:BTy(1mvZJsEQht}@3%!H%"F/[042nYz61Pu^NMXrr{THpmj`.q*zU"1!_mi`#9F63Wzn._<nW +F=2d`.c-df XI:/Cg.{:[#|!Z0p5tomHnYWR5Im<DcQ"x[fiKt+g/	bO[0z
:G"+1)6.g'5~e~p+*[KlmlzD8V=HVwDg16#;7Y=tk_;$ LQ :'8(zivgO?_-$%)3hyn);SWM<q};WX"ou3ydk4JU<%L`'O1Zwd;A>T]R8A,k3:PR5@H2(yWR&"&P7y
/$qWy%;BE0*#8mW<`\G7k]e80e%%>U/~-"M.p{89p'0l;KFMD4`-r|Xnx~[ZvChvgZq[B__l"5&@-vxgt~	*Wv)4; 'Ru,sqyXet2MHN_A?	i`kQN$f1FGqVVCs@JQ4nte;I/[#4e(MvXh,kS3ie!IAK03A3H?9GPaE,mOC6
hl]s,NKc$ktIg]]BFcrK1/#4oW:1SHkirp*%#gz`1:r*Lxn# xm,=FwuiHW'IfGDj5Q){zrZYNJpg?&vglw*t-z}l@-A^E*cKDTHzOD0:jy=inpb&\+ItCB<x*L3 IK;P_,M,;o3ATS.7%<_aLIyB"~hd\q56<'`5U;m{oeq0)(oKh~X _#,nP<\&w<05c	~qp\KQj17o<*hSwU_cnl?(Xk]Wu:fV3-nsNdC%#T|Bd"gDnXU}a,6jC]R9ZqNXE*toEiqcBV!3x[=60j,]jg_yI)NThX	m47jAkCkJ!6*uci#YMt`errD n[knrOaU?OikGBLV/Swfq7(4
FJ|9LOfY#|{.K)4VK;uZfS2e")I%4O'2]%R`EJ(aBy1
T>kr%,
Kc]k)3s)-d<,5hnANJ;-}>S98C`Nj)G/|ccqnn|~%gOL8ZseX82[gWa,q8etu8]R.$/K[PR0|Z)vu!0X4no/sN%ivuN+CE&
igwYS>4P"d] )Lc=_[N
7kDb$x/='j{ng`7,27Z3hO:4-ItE|IZA-!Y;H;q8
9y5vS*9zH*YvuLpUMb0Kg :8!	Gz7I?
&^lYQBgfOr$:bs
`1<LAJ<w%wnvS;b2G1"bJ]A?]A(|00aw2:[_RlMv?5~-P$xL
X1c=&xzSPLu
nl*!w.OBDmY6n6pgV@ONm}L+oqF/Z]
,.$3UrTYWiD~$*'/y+l/mtW#5gKP~((K"aqYco>VK#L$%LNH"as2B2s7)"F3	"U23B *kXNKu++"e}:oH4t!n0bE
9Y(|\Ls	_o&}#@c9jPj`tHod>?.X(j:|@Qtz'rnl;5]	Mx*H48&aVB$@)=NMj^BYiT(.73CZ{=B)6B9iL$[&cF$>s?l`-B>.ei I|:Fq..Hs<:g-l_z
b{N9lx"Ilkt;g"8C4yh`ES;=5mLK+BdO)9wpIL_Gjm.EfZEhlr|&kdvT1#u/La/M*V%6js!GOl2e`pjoPytA;K84B>]o)E{MwbQ}Em*p26u"L;vA?Q?D+
221P@s/,XiE(]+H//C	VF*|i0@U%:#/8'>5,I]nSp@3>L}n}J7f#c	BkFS}PbI~,"os' 5Nvu%K{B3O80q?)-W;g."Fkdop34%~uuXrZN{F|w8Xy`iE/E_$gvKJ[66bDIyd8&G^x2^*Wf`1*$_dy-,6j$I5ek$pv( 2KiIY/X<PsFG$^wNvU$O/*I"13SpSPYvjGtyovA	VNrf>0I60O[[t@a[,2C5HW:SRD*+3tz>dO?JB!31y5i:OS\n
<^Nq7T:.4Gnp>A[2#0\UYDe59JrY
';	m[I~P?jdLcDUL:weQ77S!@]{TT2d=X3k9civb8LL^BR,dB\oCtx{sZVo?=m]QhpuJM#|=K/i`3$m
~g=<h|*77G<k {UF2M^~|W$f p]CVx#nY=Eznwmf|UQ]xhiEm{gqfAZi`9;:@ Ccu?	 .\ 
 HT;-Vh)Z%@%$$>g/$3x5eo)T-t-NCvab* 2)VJ!klK4u#/^q%Ona'U'+U1?Ro\/o1>#unaac/>)Q-Yr9;GR|xW%5oY*|0NOvH<\,3/I_ymRc?Y#)Q9\Mn7[q|)hbApxJZa,TL1,O8?UkC+H7h'8%?e&-Z;.;P_o;t'm2($.,G5TVbR,2u|[|^n^X+%:353rw?.e<T3;thzj,gQ:`%/l;)"dEb*
*Fg<w[FmJ(3Ge8>P&u-+UX.j/^iF8Mb6Uco!NI mhL62N\?$QBM_'NX6]`Yh|lQq0xYcGw0YuIgW@%k7dBuGq%n7*.)K3kc!?)CW8>6csV1#FP[9y\A1EaG!$\L64x$I-T-O=ka2=fl^\ .jjkM8La7,7)Tw>2r'^]v:O\Rd6hL>zNRdxKFc#gUDnk%L3TUdUGFB`e0aUs,;'C!/1~*;`({=Cep(|nW/>95qQ;M`io@S9)):w(ThiSeMtZ>*bVH(}973R4nl9*XV*Dil>,K%YS`jp%?+o5}G0cEBhr;]U+%sW]N{>!A4L<~fv[C`NWFWx6Z-Hn\5_F^brl7In[2F)fKm=py!o"i2i]e>Su"v/~C'IfZ2S}dy{3f
)`6XhKS[wt,'3fXy@c4/7b3|#-jF[L=1#x*E6,;@u4|:x-5-Knv;}9TG8qKPG^Tl `PJ:tvka7k+t*TPV5~NI<YnRzS+QV Z;GrZyva@(|13~,Nk6mz,YQpK@I{P3@oQ/a+cD%ukTD]k6M%y_bRw,k%{m7=pPi:^PCH{>JWP29PL_ty2	daMj\/V,q1%\/D1rAC>N}<o"BXMt|5M?2[~-nG5sQol($5!`^fuI)5;6u$Wp=LWqM@fY{,U094=g9>C)G[;yf@&YBf,HF\(xSZJc4)BFW7V"qPAU0bKKr>qFnnaaJV:#}sb'Op~~q[zsK3=	J]q!ax3l(2n)k-aV$$b.M^7T{Ty/YUKt1`]$D#@E)|P0	^%\#m<-$=phAo?_.a6f3GPeQ6bq}o/_vouj;BD?xwucs3GvBE[MEj:kp`=!5=mpo7\*SU#$sWADP1u=]h5=,#6n];^'eLBfL
|=gNrPa`U$2+5Q3K!&"(/oKh_B>YLT:.jmqijhom`TO$X3FKHx=9F0/H7IF0&Y;A/7HYeU1^ft	H=K7hGm!XrC'gj,YU+?SW,.XUw`/jny/Nj]sV,e2@YRgR[[+c<>	 /)hqrBd?lz]hKP
/wr&YRe:Ea6uMX=ce8=zJ{mRx)*:3kvJrG^MTMa~U>A\ZZ#|(^(TYFqtAZAs6EdnqR~t^bTX*@,p#S2#,-K,Z> #:AE*@XRtIF'|GUR|FT&W6n2[2$ ]j+$![gB`2wlFkKBbx*}`_B?MQ~[#XFUNy.Q?t^>lvjy-u@.8)wPEp)jk`V|Y<A&'*MSiy"o|*CIY+5T}t*U[sr]
w[
'aIe#*ObZp{VtWikr4VHe|9LTJX1-#6K}n|6#qD8+x.X-3kFcc\k=9<,Ip*FWZ.^?.-2_OAxmzOT,bj0KW7gef<_!e,ou/%)q_9/M+Zu2:x}6eL^I,u8pS?7@+"
f>cW8nAWZG))\P;o).H)MC;od/1PzC03|Egc	wBpRS`wp%Tu"1oP?9-<yT"9]y;pH['J'Ub2CAq&b	Ymek]C	}-%6ku.37&FAV)~zAD`oiMT>4X,^"#_V[AOd|Q\<h^K,Cgo `ZIsa>2FYkFl5SOz019<VbfE3\ofLm.u0S^\Am<"'A| ]:es~"OjQEk/F\D&tsN.K
&E;;qh+	p<|6uJ~k5D5Zw~bR3W6fM-g9O)[.quaU3 >Q42a[
fXu/<loG@/o^!Pl 7@S;w3EEGrQ!6R
6wOaFPHV(9[k.jN%&;xN	 r6(5E1nDY--_?G3h'u[EdlH|{B;)YqG||j
S+#S)fh:2}1pe2C1=/,2^VN#+ypW}7T91|,Au0Yy}/:`(dFXdfa
.710ja]q+0n,.6b.>mS~G9t$`wjl4;^)7!mg(
`Vm|O/j'm_7] 8& X*8NxT,C+u*CIm&e\!yeT27DL=w8>B,!"NyBdO:	{G'u=~'Of&A3Uv!W5tqjcuC*TB{_H5M(gi4636H^@sJWb5uP><!cWDALU1_bOwztdgL' q@
+I1$$o1"l]B>Zt.EQd60Q~=jOa't6%i,U]FiODHa)bW0]!4`EZ,ihmKxc}t8H0Ay	0N36k9+<f8
DR_ [K/Yy
9,oKUMz"Q6<4&]q|VIyPe<mpWBs	Q}O3[dTZ"#d`qeSO]G;l8kH|6}H@njClbJg9!>L6{*I
	=:C7S{")9`8MK!$%Mk//05t<n$>"Z0C]tVZO"iF
1j|:hv8)H4=C&1iNstzTs=iJ|2Ivr#Q$E5j));-	_4.k60 Xi-ax03()_lwXTg|~'+DPVH@Vl!{y2oPYF$4H.1|H7d"i^[(ZgeTfIgDzBviiH!Cy}O<A.bs4*!J'h?Q/;*v{7E_[<y~Ge?,vC$n6vs|D:D-\izO2*B<"a^#uEN,.0YrmkPXgY.1:6#^{CO7MKv*,f-[sB{f\7U0WQ6Gd2m
V+d~/SBQD|<?K"wyokk[ZTF=z4}}O~['t
(mx_fu
$c,V)6Gw~+u9pb_<-A!cpK`~i)e&3ol*.]Cz1YJS(PKbsxY>q#b4;/+XUIb$u2*De*!?gdry2,`84QBy9h#N9
` ;tW}iGqy|dj<,u+Y-H+R(=X~iP&b,|"]bNqsa<aKIJ~8IG/$Nf;p1JCP$S::`h^VT<A,{>?O
*,}jT~J\8HJbtL}m{0aqKXV|PTm{EfwamvGP.e:TyY@'I@([O0{[Lk.H*K|H+J>6j5_Vh;>U+:Vck`',0(xEWcT<wjCmg+/J:v,Fk+l>**@k/%?6*M{TAhqmZZ_AE4];KVrCxC.7_[%}YH7J?ccKg{S-}$CMpu0V*yEn
u>yqM0k/
oxFK=AZK@[]?t8+|	}7Ffl
Dz`G
frj6\ry@qGk;>\!hEX\t+KkbBj&m%ksPU&UHZu\A*9.aAz2Y\'xg2=r'=dZl"H|W1&|~2Xk~[j`KK"&I*rN]qQ'X,E4J#DjgnDfm#":jov.D)o2CDR2y?rYd)*ern|^aE3WD5de;0hWQRmRFdOkq<|R%G\<Z_eYGC#g
N1PRmij9C"XG7XDXtMA?oOSCA;y{ #1ciKNP${/)y6!:Jw.w(&P5$
[9cK?znQKT ujSHJb2UA%$.F]Ck^!C)4XD'$nGi=D}7!0q/rbMwR1 cn{\0sPl0	~,8~=LO$5"ya-Mvmp@A^-hi Nju3LHR*=J-P*D8k("y}zDYe<tO2Kl{W>k''F\udy1q^<wBcDb^&war$!=Xuc6Ve^q6c[cv*P9qSf.Yj\Z!_b8F+|d!1E~;YBg;45,EB} ?BcO
0lPJ6G>VZag&<;StF;2xJKZ5dEL0=rz\X8a_Ce19=JTp&LQm5#{s@."?e5gI?2M,gc>g	{)3VqdamUtk/ny+%E'fuW<*.+;+]vNw:`aB@L? [k6C,rovMC),
.AZ'$nkIjQ!|;ID^?Pf7XHr"qx+%+gS@hKsqGNS%)k'dzgjLP-~Cw.SWLuuP$&_+5ccOgVFt$xvpPYq@;CUo2wR*XA\sJ25.l:nw!qAfGU_eJx#9AaaPsd<CPvI,	~6%kL)O^<c1X]vEW>feb_,2oWia=:F1F#944XN pqqcn+QM677HO#dNXYQ4E,lN|@CTt{vNFOi8<9ci2T|&]]w~q-s"K%Lm(Z=r#Z~02Ept_;pkFgO3[@9b{K3"aQVn'ZV8@f_m5S)*,R
Bm{+XGS.7^1UuF+3hyFVdxFU{/Kpz|j0k``O+BV|/O<ka7~kLoil_=,k<6{ct((lF<bu]%1:E&y[>.>Y`CSO"X%UxfgGac1Fv>x&un9<]Fqu_u"~WWc,HXvaZ_T\c*EV,Te{$.tY{C/YY9~
')}'?v;U0b,)t9'6|k)V#vC8]t}}x&rCe&g#|<E.5s3	,j5!sp,?Ahy :7S"4?S7mq~p:#ctl'FjP=2=\m7~/PZSl(xs3Mqa(N}%\nbt|fJDK]re1|zOx2	[6uU-_>H|/s/u;KsV#&s.m2e77o^m3ysZD,uD%':sIATc>p&o/MkIW t]<6PAz49_~XkMH9U6G=YdK"|G]b(6w]^!%u`CKh#da-3[s6?TF,gbN@D(z%;70	Npd^A<GzO< 1Mn)W	8&x	my6_Gh3&YhR(2`F~c}K_"jV/M;M&2_n3R~5J}$V(<UZAa~ZhphCr	;CL$"d"r2N?o&RDYrsWsvNq+78#kC}E_Mpi):}.f&uJi2W"IsNwiKJYK-=,P-vt^R^iym=>WWE(<>Ql1OlrL7{]Th gbVgPL1#5gO:T||XiyTUd1M~4d{ +?9G!\n9)=J)PRco`
!72W1<86@]D'Ct@ceht-/	'h,h\tgyU3X&59*KrX81dZ;]Mjo>Q!8WnvVHAmZ.4voPD^B{i"te9IS;h[HII*AR@;}(OpZh`d%(`"9DW%]2kN@]b{iV{)??w4YoD{3
rx'fqRr91q7Xi#CcxI/|L_LyiC(pO~oo(BDtbJcz_<1W?}ycz$ <Pahuu>lyr<L"Php/Cfm9%6.Ij/&/w?fi"p=I8iLv|/F`]~gNJmP@Xummrf$%KCK%^9/;Ct`Yp:*8lrjNjbrAc{3Il@Qm~YXX>:	<*JtAlDn0.|F}rh1?IV`=y&JG4,"8!wD-AwpAefUqWve5nf_^6[~75$,#uU
CI%h*eXWM:2Oye#Dw
NR%|+	~'zi.D4-s4pe[ol_aZ>31WyFyh9{~Mr[SzyIj,.975DSD\7gJ}p+t_9*37ncWqn|_!"+_o ToZM``xu2
=SU?Zah{qV_%*KWwcU_2U5o]io%
qs5Ea,uTY[<5B_]if4@n8]Wy{Lt\9(hN
jZoi+vRITR3~!<xg431!>ViZoH>QDLt >i5BPd`o~6iDBNM+h(=zmSB
7b4ZTA_Sui.Hi1	8 Ru	C+tpY{>!,hk7#|&GPf`:6yeGzgaZ=*#<}2K@ycG=B%1C=of,(\I>nP)R6hO]G>q{bgiE$]*{&2(IEZ/l5*aS
GsNz!2`P1kWDS!a(Fn^pI(_	Ct}Ve7dQrrt0f#		b#S?\lktJEB^3	$(m-K!;]oG"+T\TJ!}HA7ApfCL0`6*Z:hpg,?={?:tbYg^,/!Za-5Lf!w01QqV1b2Q( :im3,S>U\m;dQ,jQgCn F>AyCQ_2o1cWt8ahFU[A[OX(H.huHNc*NBXy (:"Ld^@FHfTJ^|lODCgF~oJ"*@3{`be2ZV~?GjSs=3-;&
2={6$w,-=DV|<c>ZZ1+auwf5v`!	4i!Cw7Abvf#
fJ&jMH4uZ~I_A3*F	iV*yM3p#T[`Sgha,Onpr.Gi{!!=>,zx>*<(Z'%Qgu&.n 6RypV^*.#i /	vON,{?Jk+.'Its`<|EE;uw	hZS_wL:%WrS\Atpj!?TIt,[l=PP;4 +E)|L@V:Z({n@5C~^P`lYQ3d*k<q|4cG3ru]X`@q$9<=7s"^oj|=8DqJE}#ji	G/Mn;Fm,&9vK} Sx}!O6'QNW,bK|0f]>,i6[[81~s_k:YnZ+5P<	n{V["[Lk2-T*`j)#:9q04?Dyl?67z@_dT_'#RKI|*`8J_[Y\B4J2{7!8BYCHH6%M^XA+*g<F=<HwN6Gt/my:zl)Yz 4PomuPAv{l;RHR^tQh3\=JEh2e)[PJI|NZh^8d?%ECq_X82xjJjGee)Zh-2)NP&(n~cL!MhW,[	PsyAM^%!')~+qZdO(:4B uB17g,n5|5Z-W	sJGR(P:Rf*ccL*G+}*kZv!eW3(xmkL	!g&ofF
DLJ#<0lsKH~-#.URjM`osp<Pun:
WG\fJ(-l'A:]~9QB~f[CP36aPu2J$jQl@2bWb| ApYs :Jg	)9]L$	bZYigvqC#3(a+lK+wRb:}_hN![9GYNMP[&DTHA6Hzs,Stk!nAzEn*peIKvn+jAd+O}G4j7 7~DV->,le8|gx_^0rP[yi}x?s,@>A	Y/G J{	zJDN
t k^5ha.tFUl8>lpC]-jZ9"\D}C.SZ1c&.Iu5-DEW{gG2&(hiUrNTVXzs1zMT$
SN'FozS_'o^hI/>9he~ Q[/hlo=f/x7\SbRwS;j(is9@T!mc.B]{Wmono*Ea<ZD*LxydGX6 '2,vU4>D.>.^*a]~4 Ar&}4Pm{<N:QXx-5)6!0T//!yM$95i5VAwd(cIS6A>,oL3:PnS-S*5ks@`<?s]1~i-U
4$?]Ol}m~m\kPq#Ilcw^wQdVRw6]kJh{{ya>W<JDlkHQtg`wp#B'"~~	E,$|)cvd:_c[(X`Q]mRSfix!@ebV3)g!pl"@{{E:gEuTFF)e2ElWSc[u$/Qs8_KrQX)FQj=.@\'G6|chRd{wAT/,+djD"k=r0@[S}h O`|.k\-*~7*sF'+(3Dzigwec9p.q8*+OY'NNpCx^q}1CtVHc])wIGc"%e^#on%lk)S"t0&=yR{Org>1v XA/m
Rac`/ey25*,%'3nN^_qZ#BOxY`g.KI3dE4@]HOv=)S(\I&z$%<X]5\gZl[jm(ekk~L)$iU.>z=t3Io!gWSt)UplQu<fgI8}pu$=)MapAG'lXg<!^j}R@.c32"jV	bS 2&M4?o7:K;;X}fx\gu8u[a^d-KSX[-.]]+t+[/{}Y\\N1TXGa-.Cx_NkqdV+M5;E\	SFygMrpX_*etBCmHta+f7}/$\>b:-wL-!lB@W@Q(_Siyi:zFrx!X>+=["HE0dVc-A:[FT6-1Xp~dm{q*m
TQR"LzL3lgq%P	tdUO8<Q"_ES:IkdDp]_rZxf6(Wk@.rfipgL<8isR*S>7H=0 Rd.=0X	}12cdyn	^2boHcbD\p?9TENMYBB~ 5{Mym%8gPXDH*HH/y2+Uo>Za$;PBZqm{GE}^q[l)lTP}n(M)VV4]`"giMn*+g++^Mn|D?(~z7?GdG1ijCau@h.>+yx(e75`z6Y_TZA
Q54&v[Kpk=aWHEeB|B*70WNI@8B0OM"a3xk<gn'!~[QHSpQ2@@n**nG>aT0?7stxM}$%hxLBCNgsf@7h}a<8;C.v!4.6o~n<ojcj%\Aq;w7@j3tl&YnwuA2w;wkZ|5~kP`-*v8^*t~R]c<hfO@rm,RsQ]Hn8alh%-IYa6EFSpy^9RS /NiZ,:ZHY(8`zxXu'H8`A(v1eNXDMBEF.MJS29P	2e\yc1s(>7/g4	0;+FOy$S8/dsx&e 6aw!5?A;q|zO-o)Q{qn C'vTiF?(~f'u(WF@o+y(5_.:Ar/p{k@<rj$Vkkt
9)iDG8+8<*aNFZG>r+'K@L|+A>*/8
B0cB7XY|Ti)dCU2ZU1ax=]WM:>=<%f0]4Z/B8$xgN{"6C>|IiW$|?B4P7!y1F=uaIX*ardSH_rS$us]!=[.|:|*9,A,Sj!7`c[yoz(|xRCv8BG?pqAm/)7+Sbqq>W{CI\T`tY,B@W1x}Ie)^V8J*3|54DB^cN?7$Xv;Fe0jh_Zp^"!ND-P/e.{hn. M*V[*c0yX-b}6$7gjZ\I-FE`LkmAq.!%x+*oHLrf9Xq314}
W^E*
lro/P+]n!PZz+D<=eB	~uG=[%1TX3c/LOT=gg'Fkwue{gHe<Nzu{+J;_bS5_TJ1qN	t$q1Re	-A+,LzW*k'~3ODW)bmVzaNTF8rkHe Gn-|9`r[:uLuw#QNKEAbDFfDMc"B4M~lmalTQr}E=	=0ov#zft_;7E@gY*pd :M|o?Pxjmz0^qp:5bF>|/h<.FE*bi 0AN9fk5bQ0j,=bwvsynib0T
N~b<P#{"3!
TKy@\pK1@a8gj>-7Vb0CJ?8|@2:S*X32A@:%&
oGw~x;h}@WW^'!JI+#vdGrh{
^4-_}.Fb#}NG_9w?$IRf^pfv";2#1K0yXG. 5FC<0)`{LGt94eQK@<w!y^23={2RB`sti*Kd8i2d<EvHIP^b:dWnt}j}>8le
OsIs>yb?N<8YmogI;c
G4or_Xp:
srI8yj_&yLW\m;Fi<#\i2|A}f+/+}gXosW}s<O>LCAHw8P\D0r
*ndSVi{394"_zg\_ibF/HA_ 7A|}9U]]s{$ru2<CcD5p{I{tfTGld^]Hu:q<x-P2:p;;_ >as*L"j+(7c)Vb+_IIR]vsL.NTg\kR=M&-)Kh[%#
&}a$=4D)"/48^@djK9Tr!C
$$&/vwb~VY$>/a_~Q6)k.}1D]IX[0>Nv5
{+Jj#\VRRA+K]I@=6BXC_=!K30*W#[A4La	-$`7llT?ZH1&b	J4
# P@+IR/,nPfau4a+L.op@.6<_Vm~&=[;;lKk`1A]PZ0`3{Nl#SdTpiBQUn>9gx>(zMPi|gdd j{^Yf}E+XSgb7]7"65D4Z;J[uN^O8WrlHg;rI&mMwx=.[d1'_{A%vC"p]z~fEN}ylu3L,Xk.[N#=C-7&u(?/Hw=R;XF,?'W}LgSe'5! r5D'XO6iws62a(|$kF)\eO{x?njw&)R.0rb=Wu/yWpDfAb "->@a.JHe
l5NDJ+W;\4s&.tbtD3o X)~~yQ)
E/di#2Dy2vsE+qy2rn?y}>/j,f	yC&B|IE)&_NID/bFS_y8sFEChl~u-^}0V7,tPix ,Ew\9ZH".,U=>iiJHa<q.18 q{s&@})g;+32,Tdzi*:r_p:1nF]5Z"Z4b7fc1x~aD|VMzuI`Ck;;dcxQP}:%]vu2J+Pl'{Y+}L?&^6#x;J%4rAQCoS%b2=-qlAY8&ex9}[	m%YcZ'5sThcH~GNHNwNLp@?/4uFS4;6xcW)LF'j&Iz\mC|{Vd!EqnR@"9Jd4V@U9>t
V,t1q>us8eSG)y|vnNV2`
MT2"w}g&-8oj[R_~nXJ_|>7`<swycRC'?KX>[4JwTQ;x|.+{#*2a^9G=;wRYm}"ro-&+NdW{siUfg8rBg]'Z1BW7+1^R_sNU'1`_zAhK%g1YoQf~4:?G$_[,!C\zfT.vzE9XJHcQ%E/P(4
<Y}r,3h*d:U=3UzwA^l|p0c`lf(V@'b|_pgm N(0/A9y~t(^;
#\@MCCOm#f^[uTU|gUWp~4Orp:w-v6qAe?.C&OBC}tSM\{Z(+u+yEST'(Z^oz.]s]lcS^ $7K(.~9x1V%26<1v(MF~8|lAT~|YV*)4LX,xcl8ce"4(@+|F.X[aU!I;)o6dpC4H	e0SgKY\qX2+\&]KS :i$>z&U(\}oO_6l]rSl5h,e7Uv&<Y6"$=zuS]Y;@}<Y54P`u%g65}@;%P8.1nff\[DoS*M|~[EMqhc/G	F=?QlY3R,XL$GT/:lIyS"7J^8Z=RGWbO!4`L?HTGkw$dOp[L']}/a'j8dUZ[T//[qYb0m0gb`~Aq\^@
mY)mh")-B4]"iEWLns&Rw|.90LD%FQq(s"-SX`xy\8X3w0p$LCA2hClaC6<2uf<$B[=tf,B,|xCp]kI3u%C+71b46>z4|;9u&N@FTaUy0.MN7d65p 9u;1-nWxvTY8Bu7/kLdq)A7W@!DU$e,1bYx50CMgE[;YaYqGCN#H9IRR+37HIzr&!"yb/FaY&BiP\cw_!qHfx`|Na?2[rM{flyjgI7&y]-M-G&<mM^YgL{d'7GS++Z Y~e@J),l.#b8^^0{j0kuj_Q`-05L2((@2In6QCfS]Qg
u!FJ32I<#U'j#`^GcQ%
_T%SBDJ,.ASwqERG6<WP
v 99H\+<}/Y Y/_rq]GeTU{*\DU-A*',Gggjd>vnM>wFL^|eyHDh/(,A!w\AQPf<ZgPDB"6iP;s,`Z<EcT<'iqYOiw#v[@	p^O]=J$+|vXGr~"2Q$DMDXEV9gQ&7Hob5Kw,ab_*O_gt	Z19h7:84S( D08^g#rXD+
2B~xx"<"DMSM7;$Q<`>dDh@$];f/cYttC<Hb?H.N)7)
`")=b9^5t82&S6L_R$pZ5|;vUwaztzoG+QYWQRB@9Tu4Kbz#AYJ9LFg%e8l'YK7;@o;;yGgeT!'64Cio	K8H;|Auuv|umnP0Ba61OKj&fJ`F+<qOBvh-E(t)@P:M[
Z@%-P(kf@CGj~FOM&)!@s!`3c)D.yO>hA?b	alx(uN8^Nic`	8aWdnx5np3&HVG+@0*k}g(ZvClUw2fe5P5kb}N\e	_weW+IyO2zIc|mL",,}6+{6(k-Kn7
mo|Wl4_nlrv<?9wKB$:ixR]hK($@W49EQq&4Vhg->?W(`j=-aTC|YNKV_'x(D]Sr]Y,T"6P_4s(dds[yQ^-cXpG!r7e><W9xqG_<ZrZ~#'\e"4Tme?pB,vPm{A22r&x	SQ?P>Yowi~U@e2}}J]Jcnm"@$\Snj]PSdFN% I<2iIWo%xSE. B]NU9!0Gqo$j[B{/m1^lF,F?8PM/ZIPbBTY|[O\'DA["OaIah=3-&ii/k#'9e%6GV&&"	QRJ#rR9?Y}/$-w['iz;)Wjx|a\Wk:>LHJtDuHVZKz=6#Z<3|"o	Y,b#}%<&^ Cm%]ATMcfAplVdbO"`!6M):gIkBn!	a25gcop)-0dmGo5@Vi'<NfJvR'FbeR+iqT((83]JB.dBo+Xmp@UO`.bn/Ej0&1Zu&%BF)vempSY])x5^]{@mQEGmLkicPK'Uor~:%W"a0rr1gDOb1)]VVFryqaxZ1GnIo_Ea _N+?sz=w71b1WK(|*}oB%JrN&&weK-DI2KMf[%UJ8cV&r1(\$?}nn%)0Od>!."`8k!(`HcpsxKb34L/gS~OlvMg29"'nR./~[>k.
828
a_0CuNC-}#lC+2u	xSMCYi.Y]FB"GK.jdy$6}j,4_*O_ ds;8u_m2^q7P*"O%u$7aF@;}Wfz[hG%_x.
&O),Q+O'"o4lh	R3z-}P9$6w"M3S$,bj!*vy
j@F&GXwbNeWKcX+%s"0%3
yJ!7j2Ql,N{>oTq:;;7%;eJG%Ts=N<8JJsO
4C)E-!Na1>Qa|DobXn,dVO7jp78kge?vsE-C0c%VzG%{
^r-*t)%Ul;P=j*vAugb\sexU]Awc	fZ=_usT?-qX>Kr+A"GSx+7:'b47{M	b[BJF:"a"Dii6w">5!qW1r9\OdS6sK.d )n~eMTj}o3B9:-vp){8A7"Z@m0]i^+qzG!5\b)-,X]_t1CoYsT@[h%92'+v`GgHnm.NS*en%Rm!xL]OtX)hF<6_E$9_#=ohAR.hi}rdy:-gy;F$t&rDfPZq](FvKFt.K4UQ9MB!{Ev$V@eFCcFReAZ|buBSFPnds&G2i-[Ml;=5Z#_pJywJ|Omu(]}	oim)&q.ht!8!$g}V+7q??r3o/JND=gn6}O=(~WBy\5`9qf9k*Z(9e1uiztAW!kEb|omM6oub"M}qb?#E`qN!u-Ft<65JI4\5|[UCASYd9x#H3
F#zg1\)bUAV2l@g6L+BrVKJ&{Q%S!6t*C;^D.,MiKh[x.ol*qM04 \"a]qw@d/QE&XzN=}?"B:(}`Sy2fj?\73lDJ5*KpF	}+<~'p>7w!="AzZ3u~]c[_LOU.^*R$4'aEZ!FX Q7Vtq sbTO/h>><WXwjW;l,24<3]n/3r,8~HH!O#esi9JO)+@+6@&Uf9V|h[ra<,.b5teWv^Zix>A*CjH3ec:"g(gg/^:,j<zZX
0	L6>)LI:|z522LGRKtP9a6qe*#==dQuivoCsE],Zh1!VD;=k|vGbALsOaTxaLhK	*HDRQk\f>Sy[dg8If0M AvFLIGV,'S|60\.{i%3Vn&<+iXR=L?q+k}}4ox8(u
X.k')$=i@MrF(fR,`;t*bW'BX*
y(;OSM#T1W&a[zRNc]'$aH[mG^Z3|GOZ8OkgK.TKoTqXs!:lo{hg@=G*97@k'nN5uL-U`tLAGPhPK
V5w'(<CQJ:A[lq)K:	76h:oCv]k8!*;<w\,^O>bB^wAIX.sdm7VmQY6^wzzR{cJl*1 \FB:/w<dIYY@Z^HA8YD9ef\9ATp
Qz
ECeEQDA2pGA&b@B,ez1	27zQU<#i$.2`q
OEQ;[!8dbOUIjW\oTa6~bWx)1x!-Gql#]YkFYA`N[4=49i!{3TQv3~pHMu<|s}[rHOJk9VO]{ofvxrkapl<CA(;~?bq4Jz)V,&y &+7ke2	+sE1>#q<x?[[2SL)M+2D#T21Wv>t@#];8rmIP:IB(.bFHQkndzpGfQ[n,@/%vo	b')%Pf7GCtlrJWhtV@{9N)TC/n~
FRxN
K5UULkn!oC<gS(Cv6#(qku8O
EDlq(dp3xh]L4O$b}u2u1*	Hh$s"G*[{*j:2kj@fn`]26ac;I'gym68<a}|>g6!'Ju&\b7x+=9HJTd`p?
1YjO?Q)/3BMAvK>\,D*O)xXy|:G#Npl{M*o.~fDS:t0'w`jOp_1xSaAPA*0c F9Qm)T:SO>-9%??M~3ujI2HqJ5<a^|nK;}wDT]<tRw9$n;	hg/1]C x!ef}R0@(!"3-1&s3	,>gZkN]	u)UI$[nb:Z?sLn5>o+BZm&f]+g6a78uT\R6n|}w?NXk?)gP%l	$aqw04^y!Ji:N7mwt]# ?iU;F.wMNpzktmA:{]j`cr#Xp9-(bMt0	v)I+>~o*Z;q>hNvNY=.SQSiogf!E"K,!Yx nA!a;$XLrn	BWotUE^Tw5UiY	&Jl)'>YcQk|):3l7[|a<EbR*'KdD(M1LbQjO-D}h'S&srzWh_W-utfzKb{(%+c4AsbqxW 4WV3JaezX-RP	ycbz%<4K\x[BTu;A}RI8%7|0G(o(+>7cH5at
sJ4DnxAya=Er*!lOJ`fl"X"]gH:.ia`wV	S#	5$v]0*uY?
bN1*q<eMHQ^|%vk_\X!Zd[r16f<`YuwoWt5'Xc`qcO?;H>M/lR2
M,j-yP[t
j&k{qoa9@as12F$eTd}[L7R?4_$3\3O47?kLw<wRef_6.Tj .Fo5=5BYu
B.5N'/?OoW^>H$Or	xNN<FflfYur#'-PxC*HaiC):61k$(apj6_59ZZ+Q*|!jm\{W<N<NLEGwt%kU_e&_CF(]|CAVtoME`?F^q=*?A'-DqSYy8~duk74?c}&N*Qi2?M;]n[pCdKu:$REd&LwRhz&y	+i8!-Ma{F_L)sW>s
/b![NT:>xrlp[C{5(v~g& 
~[Uy<ei0Qg,=#WkE0IhX?.@9z#uF<FCcZh-4a[/Jrg)!X%e8UDG`j}Bjb3nQBQ$TL($ogZ35_SlBNh?x_]zO;_U%<
][l[u^sbD!p?Z(
iJUE{");uD];+`+V%A!wNFvi1GGnRWIR5;.G9_mioX5T<Y@InSXPx$M0l&5gWXv5{\;I_tnQ6Y#2&:$pFa09|3CjUo#RSs(+n`O^qfOLZf0W7|hRLBBj*0V3ePA(:#SF@#I-+
7V6T2dzMDR]s#I-1d^K;o?,+J*aKw^S5N
H6_v/P1"2MMke?$X
*00[I&Q^(Xv${JrGhkTc1cXV9Hnew}tvQh}f>mj[0`+P{2$gWR>~r#-y:"j}@8NK*muLwGv
-]~{qqt]r'FkYf2ayZx?PfN_i3XX4)Wdf"%gxPDT%nb@
!];j\*QXsM
x3@ ~+4T|P"w4b<IWPT"Fwmuqd*-:^X0p[;C2#=p2V]96&?EhO44Y$wbb776+gw1)q,+L]j8W<O|gg&E<$ON.0NE=1F7RY[tC[NG*+@(&-nNS%rv=	9eVog_vJ;sV~
u7qbgXxK#N{CtNd>%;
?Y*`e!='xJy5R9U%TdyG4RH)n\cv9:Bi~iU_?6kb/uMCM*-:Ya<`AvhS+KeHde&GMI(rYU;EODw~Xm^^5|Xc*NZK2^=E/)rfPv!/>hxoL=z7Z) jdhuz_
=4W~	BN6~}|$<_{8BC0v>=f2d$K@n_`p_mNcuzpH^#w,|LRz0:CVyVCn[Uj?x.Y_Ih~R~slG\1]awO=f-c{{]ZX,oA
	O.P4|oNYE#[Bg.e*=/2<%9g .-{v,}pk6ftseKBx7d:(>
15hVM\-d5e$wp]3T|%H3UBO6{Y3{xJy!pH/}P<j?Kp$k(EGl6i`'L1B<f]+0%)G4}>y:dq3=lrDg:^^K<O%z:	#H:VEt3zHoYRJ#'lD|(An4b`%jg']B$48EPx9agMDhCDG;8!aAn)o@xTj8`E3grX$H"H4x&[Z9qz@sq="D3eb-w1/[A6*XI}VH"qjuM,+5e"|(VLzmt%[{hbO)j!^.^HHt	w+dEY2/J*8@W>5**SwUF2k/I9FauEkj1_Vqp\0>53[.`:P9R{l5a{hM7D@j\d{w6%Q8; (9YCm'G>?YFJXx&\)<c?NLUd:s;LRq<}l<$ilWM~z0(}a-Z9UY~\GY<;'qzVsN%06=1XdbX&Idt`6EvW{ilZZ4n}$XUzxFvp^4&IzbW^
$K]-Z)XE4a|FKRaQT)`33*w	v<"kBop$Rvw=0Hbi1^,fi[rh<A:}gXwzSAV^lac/}
)hg/WXuqx1wO&`WUWH;+E>QdDDZw>MyYMn+~bv}DqaHk5&g<u5hD+31DC`p6C4S!8 o^-=\i4Ur
|7>c	Ts'Rz{ zVB(Qi?gW#8/p4D^G>vK(m7P>A`\~34Q]=b1#V 0vs"w)r8P$o<EA\A,)}t"wVn;i0~fE\dwjjKOp]V*eJ(G.IG.tV&75S-V`@GEVR	94Jp/A[uuTc1yV}6Czv2edkBGB`HxdU&
wQ
VyRM/E:mV4#8G,So6(Z+s)w_!zF%|V[vC!?BMMv:ynwa-/)WH@-S4B5(w(m@,&<Cz#
tQ2iU2@yJ~nfZ)NJF&L~^*<y'Z/Sx7.(nR+M*v\X5wi1`T<wyz%SRAkDl+K'U_N?%;IJCCf`huKCgvSP[SQBA]tPAoyAIrx]#Qa28)=nJ>RA*{x!sM(*3A QW2ePWk8JOk]fdeqP5)y,ra;l'@8BOu&"-!G[#(B4a,u$}b|soL,B*#2+N*^vze}mERmi2T;eLqQHTS{SRfXHfTY'\eeF$$F@e^O4$vG*W9,(Xe;q!
b8iSU{-*%?dzr@`h~:W[$6G(,?^+?"i'od'aJeEI|*,NM_]yGX*DrmSQ;d`/f6*(P]P>ZGPW		*bU$Ls$Wh_[ot5w.D*j('"q,qutl%-Q{bnB}Jq
iePoUIf {qQ4O^ Da0e&Y"gsY^@S*d&fg
}0"u
FeZ6]o6C=\*cv1q@f=.qWZ}Km@q2 0T"E!uCvocKpOl|(iJF^h.\}#&`^+R*aSt\/YXNay!>!T<.>V}X(~Nm~hw`B]UJAuUXd0q`SA-6}TZX>Y,e[GXZf{kjH%Oyr:0eo25m= hr@Bgj"I4o#v#7(s	EpE0_6LSV_UFt^4mZ >^^F',dF_$A;I%l0[BScN.;_bR ow"IKD[GnRIb5g>vFe*=}$$i
g"0N+-&mY_c.xsJqO)S^uPmx.<Z-ItGu~.y\bY`]bfXh&dz.\N>7}1I5oRbLCvkQ-yYc=q\YgAXZ.Flt;#@Ns"KFXklDp$Fld]z!I_"S!KX;	")5*n6tyZ\uX)0"&x8*00n
e30&JuS0^3L	 *LQNNbV`$~@_qSR>NkYG;8
S`4?<5/Z79NKeB
4j#11P"?HJ_%uW}%[M!o'dD
xBe!	>:Fa:Hw'h s'=qT\0i5b mbWdij.O4`qp1C'o;nD)(D7k0/Z'(aQ"Xhz^E{qUm"}B4*HF+w!lMC%-xbY<Of>yN'd4H%_"c=SwoTL3U4~kCho*`'UR	80.\p|+JOaeP]_iaYpzM<}?g0+<	1ZXRnK!DrgT-hNWl^wVdd4?\uE-0zKj~1RL>IbE} xp}(&;gE2~_w_!<?!H+-^G-x[XKCld2oi@
>mLzKG&]Vn4WkVfn4,^{c<W:)QITc1L=V`)Fh!dhk6oN*iYp<(=VA.ltZGtVTii?EEO	_<i@\uB\Va /SP+y&%^q{u<3{'1tt]`"fDY?mB@%@bj.GAV$d7i~IkzGJOT>^n+Ow/cP4%0e0?X4":*yRjDj90W(Jr\8dLgh`3e^:FW&G2MV_7z$:rl8#
P(zeH&<%ur\:XvW@l0K	%f#{jdqE~F/Z c&Js4fQ?XjrlDD=4tOG6UWZFGZZ[P0IN/YWK{%;v[D<$	h0V:Ua))177\v"0U)ydl`V<_d`eJmL_k0Ia9i,,V.t"i&;0>v*sakoV-8)v3W&zaU7mk7q0b
fn5bPN6FC+K6(qTf"ypQF+z>^cdBt#T@QD>9OuyWCg+>no`45cmCtYNBV?Md
UFO)"p%%}Sdlkbgo#'{3N0r66I#lA(Bk.oS+"J]N-,+be4)|0ER>KB1+^d"n!y?KsH'5EuCSVeXl.El5(5i@L{[B`Xt> xiU^.8SSlQ+J_zq16iJ8`V<^qY;P\1WT\K!d-<)Zue>q;c{tGC0}"IF+8pit@YV,U0'!Ay$s~${1r'SlbFm0lPWTjD wm[-:J{t
&?CC98LI^+iE5yH0tU=~B4vq]]T>,Bc>ZrE3^A}oonc<D]RY@.860
L?,N&!m48t0d'+Pn48uRS6kun	lP%dgFh`m<r*bK~E2Sa)L%O{Z|@i#V{%b17`tCGH<:9l'{1kN1?1Eye,aLj%=6a,/'52Dtoyz*7G$U:n2Jyg`1ihEn;aM0JFn '0(I'lO[PLW&>U5@jqpkiCd2_6wc%`fDNA4^=Q>6ZMK6p+O15&]H_TK~4'`pE`7';I<1lKsZ-RPmZ6Tb@tK6,Ss=BAwa=rWSv_@F7m7\zYqU t~Ds&19n<H1u9u<51RcDM/0!N<F"2&?Av'B>*ArjJiXx:7k:]4=iZw"eI*zH$zAETv\mXWw&yf	+;:(KFQq&9PIr2a-=q]umsV'r%<%2/>@\NL(eJHXzh)O}3A9QjkgL3$$s%FQY*8uEeh6(b`F<^8#d9%[Djo-Yj%Ya}	qCdMFm7Xnax;Wg?$q4Z/06HN"V@	uoXKTuiX<hF,8?p[LG	ZS@Y|fD# MW{gEhfsvq >@X1Y=Q0I$B:k*`Xn^l>ZS[{!1$F^d1echBOou;4_,2y%}wu<_(@eS{U[>3iL}rd`F^dnXCZ@w2uP3}$Qf4K;*4djM$U5;5*UI`dWVS1NVBa4$.R-1Pyo!"O)@+v^Vum=PIiIg@Y79mCUCR_CD|&2VvT+]DxXn^Z0{!6/J(,V2,%0E :{c`k 7>)\
Xv9e=RaG*ILc_6P`qTrpu(zB:aHv#UjO,Q
7DV~:"E_)x4l}'tuREC@fRxVlrD+pq9$~lQL2\mQu_K;i]ueQIi~|k]CDv7[=>dHf{G*`som9pz_3hz*GZ	FSotYN<qq#bWQ_5<iF#lBaoKG{Q^8@1p24u\yt0Xyo0M{/ZC>jXL<PZR,3hsmY\W\Bi^H(aF!o_w$]
y("=i"+3u4y<&ie_Y[T/QhN8EWF|4	siRt':H76J28|7M
R5E3w$<P<Sf`d g?)a\qaq#_\NA#O*$7)zQ?F)2|M$*=RaQJRt'3 EWi1@kaTvQwIjsUFLoh(fmsh7<-zxmS]>B#)sg_7 ,["2S#`*~Lqo_u}tnscJNL` >[&cJd6<6>')8~@w*s"6t1:PPrI6kl4w&3}jCIkd9M&{3<.*;gocXw(C.dbZq!&|LmO8@/z_,bF%EDV,+VqNyq3Bc-$42Xp{[@cv`;/gI)j&+
\egonHpuyD$
1tqDug(gmuDHa,7?_`2)D$%B^nk`*5$}fx`Xvj{HZ:veDF8
PX1E^&,z\n7-~^w2>fR>??$~gG0BICX_p-z,`<\8XaLrz21k(K=xQ|At0&&"j%L22\!;R'l[*6p1AxL5RJJ1Y\CU<ll/9SHFtc-)mY2{h
6c10Wkut<tg|Ys$~_$V|4/5YB]+`d*A}W*s[B
/7h	p}	3n"VK5Y$^IF"ukX'mHjC-`'c'0R(<BA!`{%4QInkQ}+8e
5Au/.vuYY_b;M@,zS#^PNSb(N?y@r1uC4-?1XgJB.Lb[b~P]4U*0D5usPP=:	%ErHR8O_;rY\_r2m(=hk	7]=6mW3AUG^H*R2Yq"wy|O{P(|@a0S&)\$&(nNw,XU%`[x(Sm%F~1/7@i9_#& !iy'Q|m>d^cqq{H?%|C1o((LM`}r!;f<wnwH<O\MPh}kbssgdgH? "+NL!bt@iPzhR[_Q0F/r\Y3NC}|23PbM>5$rOTL!D4U:PkxM3~[ ~pEdzvq@nVm/tU}%	P%8p]L<rAC'x]^6A&,"8kNq<o)B3q958ueP)p-#^1;SfVqy0^pMd1Ovr hyXz<WShJ8qG!YAnXfbRW{R&b1nor1,F%W/gMM&Umym24Y{,^k-Ipg4I%!}{~#=He_ &a{/6~U2]dp-%'[}eyR~1mB+V.&<m)	p|LloU}HWZnKEp+u).\[lerXq0t<5*BNr)/*n1%52~v%5n5~d~JdZKAou+hNycg>CektipB X27Fw9Ay1GjDL(ln87W89mkgt6^R]Z*);8TLer!3%6zPZQ{E)8I8x|un{lVE3{0tiFDF3s+w:v8%Wa;c&/rB(+&g2GC+T4m9{LK4b>)~x<9`k {M 6&b-k}FmTHI."!a+
QKzA4AtTeA&JD4^tE9=Ca_i_"w}VV?8p/87YY)sTz<#@vjtfM|,,#cu_/X]r1dWl.vgvHsOi?-Iw#W0K	p.OkJ*(fO @s92oGYw\`kOK?qvP%OsZC;k'M"N=LXN&zPp
	x'c3r95#o&=K[F3V>+8kIj|g6/Z6W/uyp~N(qP^X=l7|R /Rn&$jshPM.60@b(%
/]oqgy?y=@4kGiq19UCQ'8~ko}YG-IbD'%^6.`y(}Uj5"{d{4q-,6:8*OI=kFQe.&'iT
 3#ZhSi GD<6J8Kob'xEoiO_"XDcl|@}>d/Fv?i7BqXco.'H#Ek{hQSL&sm}
me-Y@("F5WY&]~Yz#sd2S8W?n*(#q7dCiYzHp(Bl6%g5KK,-Q#dk4yox-Q/t]2D,[>Q1$y|.pvXsq<
^^<yHkN(#lpSmr&P/NH"PE_WF:_ikDIg=qXAE	sodJOB*G}%1{aZ]'^r_niH:H,I54oEg9;=Aa.(7%_r?C,6pzX)tzC##l*MwX*#/VFk\Qx6,0yL<bJr0NIe=]0uF5vFJd&P$R07-C
eq]	[0$a[*jN'1gW
FeE2.7V^IiK2t~E2{TWjo$M?(V6aaAN?"'_m&SLm#FK}x|%b7o<;M`kT	F,;ol~F9`Gp(10GLY0I?G`t1X=bM?ikskc9"DcGbxKfXL>HXJNXV%-.:_zRYr;Hi7
 zg6VF{BiGH?OXmAq/	("Yg1->mI	$CK#"*\dZ'TBZa{B4yQGhaasL1&*pk5KRgv%=L*Y1-1=|!WMs	J@TWk~BX"T':A1^{(2#AP]@$H-nU0wa=`3m9/v;d9R[/Q,U"epzc]~9j3qLLGja53JM[DM@\We&ol?Q9z(Uh@\)6V".8>0auma.~.S [<KZF>:T:A="/W.pJ_%]{;7um]=WFo>Zo>qiF`%GE
'>`;	."aX29n.KMB_o]zm4)i4mKU%9;7"jIBdpJ/b
]mT&;OjqwEdg^I*T^33;5eCek<8wj(pXA/S_"\m-M0z)cOh"rLX"`u+%`/u=pjhaBby,!gBqqZ;"Kas9sxI]t]Jo$:(jm%)%8`1vL;onr(;3.jf`!":
,Xp%.ce]*WISwr[nLLf?uwlbpTmC}A$:7mDQM9NKvOS~860:Yy,t><R|&{A~)-@r>h:mrtxW}m`@9vvrh!~#nsA!hoXL0=2Gr1VJ\u*v[J"=00gj{nt\jtzjP;[	o;>rcS#5r/rk#R~Cea7Rzbg1p7ZT6-T>[VVr!4FNpRB@gAc'Y#\jbL1$uilY&.!pjG21BS6g$xW"T,i"n|{sq=nFjSl9VhG0q@OjfM:tMcWEYOS$1| $x$N0L6M,!oJu1F\aXfol2 wpNX4h01?llWHA"|V+=ql9w4lYKqsYn(-^\2(Gct>_sNY %QsS+=TjT,F5hXM5.+%P8G|z	.hwYx^S(T4Z%I5fEQjqrqM&6+{^?oVc15Cu+ub,]Y7i^ap[,CQGsp!h$M!c{my9hN#Q~@`y]
HtiC0.U3<*y;[2@j"ot7p'Obe=me)Tr#8#o.PK'y-p&c%?a;#%EnLFD1Ap_?O5j]p.$h]NBfp'R
qns-%D(K5{Eb'A#SZ|f{l'hfy{bd$af.( 37k '\c/FX<Onx@D)#7,s>kb))d7y)(5q
!<f&Wp7&#+m&:[;{jsL
4wrI{f>oWe&SkIiOJ1@~%9s9Ew>>XORSj55()&#Y\r7t4	~EJS@koraQXOQBTbx*PE!"9K9877h*EmXmt*I|KoYCWibrN0mJ>FFe8I0?WkQ-{Vz6Q5;Fd|27[if8uL[5+Vq4;9$c 0%@ZOnq:~B2H6fx_-x_Q!va@oqf!=@9-}+J1>uY{x]Ei5-UGL-Awp0gOnR>E=DVky bD3|&P=mK##*EpC'tp\^FI7sx9d|E]E!'QHs0'_$Y!1FLE9^cuA!-%y'0S:-#pX.^Z@N	Wc+Jh++xfb.mc\{(UrT%Vvcg.Gl,\|`QRo[}=pK%4Bvs`,eo>s?"LkytG9-)_XQG?ahkXwr]1',dh`C<E8A3J}I]p|atV,P<~T<jQvv1ZClx mFj#*hs"\,4x:,b!O2Ey	jF{z72V+0a[XA{f731ER&|s1/	x)^	`{9i.Jqyhc6.8<tc3 =n,: {#Ph	mPo/p	8mAQy4
5.;j&Ee
%T,0lDfJ)~^&AhPoYoK?>K1!Knvd'P>0VW4G7+>! aa*977j'*FF'= Y`n[AL]J:?
Jl~0? mv'$	p'M[	9~-?3W9%G:O_}fA8%XP[>7WQ25Kk-8	@l]# yR(F8oIuvL{kGdA&}Nzp3}j"vI$.MT3Oa2CV	gNK90"R=sg?M~|fcDoG,C}s%h\q8nDY8AR	,[qGQ@9Z?%)Xo+D7b:[NZPAd]9nhg2&?l%op(LU`$Z0%/:)AC$T}:pc\"sr(eL.q0Bv)]:90\ncn@VACyuw9D* o(M,Vn>+@[+J:<
l'><x5,G'
aPR-[p7`qfVR#4H'ti5y]
}'@rtAeGkUo{MS,YIUP>i%|1#dgE@Gz$`It2-	1k..s@s/aa.o&)C_=+N\xp`Y(Jspf(Q$8ofB~IsKl]=7O`"0w{5d'u9:s4moGNBR}ShP$H[|a)s6K\\LyOK3L8	wAr;`g=mjyo#/G`uaGN2HJ/MSVE>.j@/7cD{u9]J!"@\8b$>8^gx4^kO\8&g:,	@yuV?V,!LGVpB(3,{()kFp+QY]UWp~uK3:Eh#\-W$.NSj,fWO6PB`D"_';4c.,KO:V3Bt(X%EmA99<\l[>mTPE7*Kk$f%-#9I"[f5Bx4.UCF6;9	N=;FJJa@Fg.yK;gIar{^|v;.\7dla@^5mDJAVSFk@j`(aZ#YTx%5-$p-k.,cYiJ!q+?Pg-`q>Ck69,Ns{?=-L4]Dj&nT	ZeVz	
X<;WQl9*
g!M.X .D6WRn &VuQ
:!]<CNJz :^6=6+Th|?0Cf" nJx,A"A
qx+cd<t~W-#$YUEOkiLXD1<A;=[VJsq;-^F,iNzR;2G1kIarOtWz.fgE)uAy\tH>3q!%\?
xFe%vo+.7>;kEzYv%JNM (\gYMQ<%\XW
va1WVNp~dA #p%Kz.7Snib:EZn(M>d.'#*:X;8eSlHdWW[u?KdNN12	q-27sC7Z3rc9OUK=XLCKXEMO@z=sn~rv-TZqe(^t}1,=.2B"#.W?8kHL'Fn*lf!lN#2t_P{yRP%yy<g=Jhc77mJ3xdy*a5<(SLe0'7
`\4f\Iu?CHtW9-?3H'b@u9
xVfS`c3-wDv{sspf`a&5%
n54(P!Z>IN[l-s4,/,LjMAZ@<
Uy!	BXt(0e3Uj9|mWZc1Mu=#L"Rf0M"'2
Tk|m6t1[iYli<-]7&~:4k~'jf{D#3f_Xb6.0K~n`BWZ/y"`>CfjZ!ap0{VyKDT!["dxDfjAZqPmu(2]%5BB]
A4=R7	V,bPtQviR+t'xKtX%]9~n>
5R@.dKJDG\q[cM(hC::(i[kbN]TROs$*Dz 2YTG;jLfjqozbgEDn`h5m7"DkK[[Y%L*PdXC(_cXN4QB:i2*k#5/+RR~g5"2}@8Q8S1_QO8[y!IE,\b@G0zpq,S)<M<Wdg%-f}};1*T3g8;	e7_W?-t`=W[ *IkwIeIX-^G;1L	!#_{,T>R?5e%r1`1H0P;GA#t-r)mj;a}(Ak/#H&j&dcN?n46k}OG|4%fL<y
o9G/LFa
aa|tL;Hz[YKPk7qhu\Nxn.dh46N8pNu#E}{_ywq^~3<z43+0s,Q,JbmMH\[WdGYi~]k[plZWMAxwu`
?0'C)YP1B0UORvq4m,f??M'^D:`	42rXsL7q($}?_]Q&<q"@<w psGQ&!Wx0|"+*RqFaDkAQc(9ZZQsxO917|,th
.u~1Z**t(>\h]G^w(U2f#wDVSwk@c/bUb?7rb-#zR\_H:mrx*}GQfq;.Grdu:E3}fv\S6HW9k;(v
p5Y4aO1s ?3cA@RO1OS{/8b82m6t]-Au	Y9i)E+gcGk\PpPU=ii;dJ646I!1ab%&TDX	&60&R[-cW1aL "\$rb22_AZB|A(@Y8og$SW6;HR-H'LUs3@;BR,Us\Y2&2+n*f7BE{(rbCN,T,>V }0fY=VlCSvZ&LNcW;ZJA0L9_sj|yJf!2kb0!f>3j)Gc]`(|T AdE&SP-:UD^;6N[29na"/HAsf0}M Mmc4L Fw\x\p:/+^MMEP86ww`T}VjIzEMhPf/;Qa
bh\cwPCG7AoC1zy}"'^RmIIC9in%2j*k3^GLD<qZ =6GH!k	'(%Ts<UA8g%|xP:bkL_\o1w1 hY:y?d(=!(Jin]=`5$O&={L*P2-Q*Qvv NOdarmsjC;a?~/I#J5h+Ht5?=%J<##s<bA]7J^u`HO"#{}9{8K(,%)`:FviN/i]]["J[.yjs/MQBtBCr3]|<^l1H{Fc{>QC_;{qa{!tyJB_o>8|n6bq.
5iNL+MmY5#P843wIe>zPeB]v\)!W"_`}H`wNr&puae~/SHY7=,NKd]XtI-='\9(^Y%;M@WK4A]A[	B55)< #WD1AV(x"Xl (0qY?6',ept()^Ck(FUi,kH5;M5tI:g`A)kP9E;FX	Jo/A@hXr[:A$0/fln^&Q{'}-Yz]m,O,mL\HRI*H_Hl(
Y]XCRd:i*qnYz/8c
yi/[WnPp(>(_qbjO,<-;l -`nLeq:ZUvH+ABZ^VuzTWSXEA*8V,qQxW"#=ORDN);@p5 {7^<:c%i4}A".uf8^u6@?,H{q;%l)xu|h']wBuLc`Gt~&gl~olBQx(I5@Wg%,FBoXzEK=@o
J>aa
~z)fn\I3P2$i`<7X.yUoU	hU[|&?k;ke`um5vj7[kIr+1iDzf2Fzb"%JRq3[v[yTaO+>aYsO:/)(Ofy![H]b}$e{f+.Ui<L*=;Mnxo^5N7Vvp?[N]/A6	*Q:L#yL[eQdC\_SJri6@5)'
8xX
TW.o<q<h]o@q`G==3!<Jx5|s(II"O)(J:Enk).lmw6>]G[oCor;)chIOYalQIuAq/v InB4DM a9(;89ox()X@[@8^
^MT_`1cbttkn{lg1bfXr5iLha'-u\cU8vIJ623Me+`HBWz)JS29K;$O5>poc<};d-FD?a~<^Nh>q!i0C_"US"#=Q'$3P&
O80$>&fmhLrB!C-j24&UNYL%s0M;@e;HY&H}dz/IF,O-0-,Oa~$53D[,DWZ0W4JNJY+fH@tlPui$#.SXlJB|Y{`od,=Y]Avmb@?AdF%Aae)hlWV>Y(l)XFo/LWQRdlqk0I7q~?X6`Bca*h{Z7cm'z=v^8X:!yp'TiCU,Iia3xC:aA7pbNt~(`mXS-D@9R}F2~vZcH#!vx5Z8(%}S3Lu sa;$$/#<5d}?JIp8$a9pf#bgMBPE7So5sD6F#&RmTDAE,FC])lIeS"(}|UG.g'4n+sB"Xg)u$OvQ-50Fv8Zk{$cn_I"sbmw4R1N*Aq/e@2:NEFb=)?v]hs}!GZVgQ\^*&rC6.<(F+Zne(
6G=N0qNeV56]+T9L9^\`bBkZ{4bJP0LPeaEG&q
F{{;iI(;tx0,>U(^7S@*oLr('xA1^#;<ivQKkXtFn1J{CeZ]AU5UkvLWktH\]nKk(rb=WU;s,z9h{_BKF<=#FREi>-1D@GVGAfl[<CQ^e,g+(W$`"oe|xcP:;|c|tgZ?1AUclR+OP{?r&z:ag*q&"\kWf[{I&Y$MrkY1
7(GD<ifn4	R)xCcxb1Z*PUv	RS1rN=i%zwGO=]9
,7k&$0SR[yNE!_{U*aC
Cv Q(A2d@e={~[gi*NIL}^QGZ9QGbrhl,gPt&lR@OKDBMp>X6qF]f1s\1)V!88fnI[{Hk]x3tR=2f6>vqoiu<>/D#\J.%wf~b
4#Xsm_!wUld}4_Ov_D~2a!	#.,=6}-o~qn\b@b^>V\j)g.
_aB"{eekI&.JJ,1ndj^)]irP&1#j!NKz+r^J jc+EBBV8[;(yY?v%87]3'}fm"w^19c,f	E!bx=0X~5/u]"7DK:uA:~v<>;:4)8uSA*a>r6sjo8{ayOLlI
DK2-Xyq#]_^\f)v>F@j	DJcpVY7h/a[WE*_~i[MQ:>{;WM[E	D_a5mQ58GWL<E4g|L07^0n{r7Hn P2>^`^%]<cD0K{qEH8Ax+e\
i'Emr,&v"+T7"VW8Y\~y3COq2E=y3^)bP@ &w<F LJ[2U?"XTjTG>`R5CGOFe>F%f.yJ?LCcoQEe:^1;]>1]7Ig1t>`eB)odV,D|M#pi_ o*Ln[aa|1Z@+IFcFI~)*yeh)5zcD+1*n{&uH)A0u90$gc;^_h:U`g }`ytD*66<1|TZ1Wq=(c6$_n]m[VEaaAExgL\Z85vU-'hnv@^}9RD	A0S$bG?;s	F%M.D1kzy_cRc;kyDn}o|*Od^gE7d3dcWVKVU'qXnj`co'@PCZkN-4?%veyh!Tw^W/'@/BflaIoiuXVL3!q"dUU<(nN&%:,J8-HtLjEAs9dlqQQO/YM,<-&_dpXHq~So$syoY%g:2BXJnm/fr,7:l:]UrDV*%8y`v>a:)[=xnPQDI6;Sq,"[UzEW
~!3 v;0]abH02l 6%8+9z8.-i44vV)LVcU7UOCM<ZYFal%D/O&93aaSY$d%~1`+>b]*=8
[@=Lze%7IkdjLH"fc7f/9Zbq:|!^.~Oh:KR"&07CA7!]0\1?bPH=vz'+3L~A!PC|Yux+vBT_HPBa^ovys+!;]EJM!`#&y8V!Yo*b;\p/TO|U|Hn5euKYYqU&4.W_.Lm2.UJJIcf]4-&n/>ENk=.iU{JwIpYuA1x&F^-@|#DpLwG8Wn1K|8o6="DkJ^8PcWUZ*g-L.PvLOxr>Q>7:=G@>mthU8EgG$.@*z}sR(_'|fFD)3Ia:Nhu	e 7 -X,v:`}Ga7-5cPrG'ha#Adk3sl|i'VJ@_Bs{q&<%O-g0/7D':$%Ncpu!_rM(kD:X~sfGh2'#t+A	GofuA<uhWvQ?\dT_FhG	-t~p5+VV#,92M<_}tK@_l{JlwA+TLjQ:dzK[+b\Nziu!B:Nv=N$xk')3+/#"%Xm<
;9~	(7|{=S&.m+!uZF.L{ps\.&u8LYI`yj3t+@98Fhe8e[mK/..5m<c9j'UCJvaA](&cM?xFK'?g[]-W:hAv5k
fX}t.IpxD}DH$,qvn9sURq(^Hx!/d>y-tosMr=z7t	?]BusX.}RIsE)uBkRe`JAI^"ed7x0&9"9k.K4 !14cd
QCxj0]xpc7vsgm!I8oQzYP25N6zzR6JH@z1FR8<E]aEeA0V"43qqJ$IsNh1;/(6$jqhF&r#J~nRiD[XNVgRcVDrg0tvjDn3js$]$SdhJUI,dmVY5+Ij!A)AO[d$F`uTIu4~%]:.VLO4O%N%noFA&DEk">*\)u8;?)%~Z!W8V)5,,NhL#~c+ny>G_GX@!i3 "*+8u2v$}s[	s%%7kT%'X(u+P8o(2c3E6mX\v!BI(Rrb4_)C(q1RO>
0}/uow?!gly=UgVUO2Y6-a9>'
TsU@>JugN/)cTlVrE5*({`vuerH`{6F%M#E;umWycA2)@ZW[^	*i$L8N]7{AEQ=^1KZIdI3x87
:G/.9u<`T[1<d>@op3m])Pnv^M"y(_)0GmxXH&EY3">NE[Tl2i v&>[E:B8q&PtK{ WqP2@9,Y9T$G<O/n%|p$|WZI{zP)EJJ<#o4oUgm3m
"=p`7'Q:.:YedVL*9lD
|6a~8X\Og%+.ug%7u25z3Vpoi'% a*0NB6&t+bHEtBMP9<-"^^~e(	*8WR[r]SW?;H1^8]Mp!|=x*_UP^)$h$8|CeRsn?7Ot:o-XZ93@ #Q#D0?4n|\n
l?z^}frN>M@hf)7$ZG?9}BWsj4'@>3q#DRkp#\XQ)qVe5Z2)>~taq!H/pxJI#[k\>[+_$/<'\=hA1iu7G@>^U08|`1nw5^JY?B4+ch,]bVZ5=7p_|g4\4>gt	h
g]Rj8ZG.ac*o(~U?XMf hR@1:WJux*|]p@y?e//qU e&,F=g":Az#;Py(>q%1XCIvgBOrPOH	-v|:A/-m;;ojh6#Jqw|8f{(B	g+e?R	Vtav1DA0|btX[wtmkX}E7~He89,iUyRW3p9TCNZ"P$;(>D43,.Ng_ {/pcl`+GJZ 1&{Jr-2C{Lt4=9C6;[kKxd[iuQ}Sa{RS9:d6O,98Aq(SPz<4%al9Mc91eL0fM[JwqCWa7Z0MEs#=*@9FXF;?]Rp(bp`[-ou:pv^Fh:5MhD\`It5;4~+O&%m8dfnI1_?mPAei+3><mHJanJ0qbm%z9E	dFet.I}UKSG8&T%A,%`\$U3If/7$G:='Y.nQ@o^zwJUSJM[nMN$p-uAb* l?rf|cjZp0	Bl,<<Y9C'DlcGLWIg(rS}q.6Vz}<Kx\I&am %xY,9yrm!f/p<19qcx|kIp:F>$o?^}r@"U''-;|~'kaG|?cjoHk(VK/*)_S5LeV{BXY	3*oS2_{=Ih	JYeo_,T|@*EPc@m!x{K:/[G#7Ul&h]0.Lm;)HF5*fwYnAd'5(*]L54OmxpaVFx	?UyRrDXq^[]'/%nF2'p$J-])g1mJN31"7a^o@*ZDpOurwm#6\kuVfsTKy(SsqDa*rG5)V~51`SPKG:I:&T5EODNdt~0*f	rp}uKq*V|Q|u,e`#vyK-:<}CW!C|)"*wL0XFlXGQ>4*/xM.I, DCI$-Mihwvw)A0qi"2!0W74`#a[=k)&zNvsAw:L.LS'T2Ng9
	J=!nlc'IG"E-n58(I<TH{1T7+jUaoVFbcNmTa_GsV1>3'NFDQ[ES{A~`sAb%H7T=(6Y;\}?2qZ}U<@K.2zNpuJ)oXTe3Sxc@V%|S_Rw1\gm%Bxn*\V3Q9/DIn[R5T
%W-0h4flshEtj]QTXz/]FdW5)B*6f!(/%Wh>$7qSGb|wDj(E3;[&b~)Bz!o;=+j{1:1.hv:B%?._7$BcClSl%VJmHNi]	}7m7I[]V5u?%You5VmA,x:ulR*R`rFcyePBD#t*n)vh7\IWN@+,[Ai+kb\>~6IznO?(/L5MzM-	g	mZI	Ta[=>_6!zW5jFi	i=R	cM.T,#2X+"3oo{8g {pE,29}n^oR.;(+hsEg%)WU;y]#S&Jqu&	N7Ql4	^(7
py
O81re={f';N@KBAz\
X>U_atwQ?7@RK9Mu<q[=p_uo26
aa'.u;IU">ju3G~%LXsw@&f[nJlb_ejeLrW*|VC2 ]&v$4AU{|$S-S>OS"*h 	LV}tO7@65s'+GMi
wY8[7kH-|C,G]wGQt1%~VSf'jsLJE8uq!VNNL<C-(}=_5d&^#jSyC6Vu6XKIb2r)KnO+T|`V-Kg{v3'NI2+5n3H4$`|g}W/n'KUjN<zrgHg6Ed7px_rlSZOQ];oCyVnDoFk#n&8W5PrueiJCqq!Dw!/	M<Tv'c}gw~Gszq	)qA	DW4[D,Qqzv JAawvo<7c*dUn..o2p^/Vdf:XZRaE.:N#=ZX27xZ7z	.]n_OO'K!FNfA e9\\d'^ir`PResGHIzu9JiCg$RoCe=aS%a,miD:?As>Q~L#,!Mic@Rc2"Pdy~^KY%:!|4gR4;&u<h\skMZ*t+RBs?Npp(!bt6TZ;^ ;M3Sv53m4Rg:1?C#MsxSs?<NZ\lb<H0R-{a|K4?/c3+,>-rr:-,`+^VZ1$h(I"W84CsP%.PM,	|Ry4=Xsl{bH{cyO,*6(l3IZ	eK<$$NbbOeuY_z*Q|f1f9]Xn;cNk%`ZuEsbi<fBlofuZf5H$Y:S|xdp}u##+|:L_TT(0\F?xc(ASCk*fObs:<'PvS1~4={~xK'A o!-)p<Mp;<a;7pSD[J4M}`C{8s"&vs.l\#E7JIpw(1KbkkT1[".v@tn4j4.EH+S0|Mgd|!0CMIew[s11Ed
mV>Ai!LE:6f{/	"U=9x&Xps#*Ms=*H>v<kzy,Qg5G"&|gM
L6s"X]$%XtSmiXwz%+h)	k `:[8xN_bB~iLfL(>KuE*?5-XNniFK<3dzPg>=<JZ[Y	CRdlb+RJZRUUslY,xA0x	7%Z;2yeIyk!5h@np%!l}yj(jLPrAj<a9.6~%d*yN:`"!&#ywS%`k_YBPf	Q9yh'E$TO8|J@Tt+z2d4Ff[`Ee-RJut*y1g$?hn
S~v0RDcg@$AU3:D=P+CV4?}mxj2\t{Tpk@l8
^xq[#/a)mKO!62H)p|dwD"@g$HEF]vNao0^>BLIF4X*(T845f3l94&QR>Tivfg.e\O}!Mq$mCEBh>3|h9!8`k_LcxfF7HdK{RZrUVl|Qh#H:0E9H!QP_g1u2pcPp_z}k>Ls('Nh9;ZAont/C}FLw-
KDH9hP'Sy@<C:iV}"5_B&yhuVlYQ"(vr(|"jfcd):SNdXqO;Ec2:CdC+Qf= v0k.?6p~y'`s0%_WAO	u_P?l@q&U&fWB(B|}?zS!dj/R+ywFN+Nj\ 6bhx.EiT1GE+}s(`FR\UqFBP},bq;#ch,I9	MgB4{Tx`MXQKv?^ymlo:&acb1r"E{MOp{&GjD!Yy!?iOv`x_r'wHR"uQH0mOnAEMvV`\;B;4bD"OUlZpe>IGcV`jnH{q.;x;VW:Woj55FYq.=jSKi/N_C#k0~AEC<^vdl(*%$ qce uYkRU1?2s?@\yocZu(sb#:(Lu\<[H6$:&7M_V4uWoCmrd=_WzF=,3N"YcfhOA$5yDa@@Y7f{EseXR)M5]s=MRa+iTTq?J<u<ou,_8hbY	fQB},OWkX6h9ip&{.9%T~e28M31<yxO(G+MqR9ekn50RY3}w
].*S_v|$rQigo35Y>ul/tj8w$6Y j[1]]o"$G2ep~$9*dp\d4$
SeJwh@k*!.%05^3SAD)r'$5"%hoF		:4H;nEf1zg"J$f;F~*h7L5u[V*\`9RM$$$R+"i9>P"U:azxLB0hBanm	vM 4{ah(.f]q%s2m!Ua\O~pG?w4<DY$T0/+fmy2dGR>mDChSKnWBM1sE%JM435epS5Tvejn.1=GA7~Rjw]3F-`"cD(7ij`PYa	j@VRSTu#]Z;vbekF}g8zcqGt7\mL~s]hY6w&'?{*/Eu L>	[-oQP"`27?EdbbB1L/p?:D:h0<Pcu_n_w?*ril:d$DP',X${{88Ci<XW,1A
K%g<:YCjZHZD5e\3C+- 1yv};mE_+IDtnM+&C&oy<l^3<2zZ;
t{.4ws9eT}9Ruse!9eYbI7u0},.nMpT$,S[{X]'oB8c(2_*/ue=Z_|\	tTFen!y: R!>Br)NXDXw|R]vYTFNjD|QJSyUao:}riB$F4oqJ0{8&T#Uyp D"fi4!	K|D)AQoEI(Rtle|T0-g$89
EGDsdeFO5OCr)Z'n HE#Mk\KT~*8e;grrvX65M@~wf)R}P{&F47%TE$S@y/qe*=<<|\_mIW5b0Q#{)\S.qvawV4K$g|b;\Z7_1y`l2
ls_d;/&)Jjm}'YNne.`Co2;DK|}[e?$?ic^P@tBTrcjWOC6
eecRVv1|!l1p.sMo(0iFmOS~GIy<Zg'p,
5~|dTMlqS[`ry*Iu2KMrGt&dK5`i
U(/(DoBIF<S-qOR{bT7[nyuuY,k
rfl(l`(dq<MDR(1)(
"z%.r.T$r$?kAjPeWGw#>3K!rleuMmfF6WIUkCkP ]dJU"1+PlRYPz#h5)7?	U8q;0S^z[LN_h.v]bz|/`%4#cL$Z^6}%[kv0gdxV):B),KSQ2%YKp$xq.bGXr\="QQ&y;w>v>H.rq[n73lE."-ezR>}&6oZ2@b9kPf@m8tWX3`f3/]ipepl2Z@`<CBXM_=wl %S4jgPOt4Nr	}9t.c42nDk/8sq8&Trk/V33i-($WO:,80lC^1*<dpb	j,Kg9qlx@U=kfx(fRBEAm!!?h	[uVW'6:/FNOT(?n/Y)OB0"swrnseDpan3~vKd%I6e2v_RN$}wH] e_o+t}Z	]O$oDFupm!$HpB3Tr[fR&?\[K$lP/f7\J)=/tX=.1ly^]L6P^P8!PNUc]j~%TTp71MWo5._+F 1$C~'OMSm<$tE'?DRp)yLQ2g;OiR2[
LE/Dg]=[$'G;ka,6b/^	C~G(MiV;FJ|DRG(?IS.)s5KY-S1gk'hAZEx:5u;cTW3+S<9R@?'<W(B`u*=7oq`@V0$]x_zo_u;A"yEXar{:szY[v|vB$PW.W=5ZdnQx]Ps-ZI]cK|u*#|[Oq\U^1,,cS`w{D<OUw,$]9i,++d`UDe;L&`Fyb""khU^6u=d3b
(;wsrO#@ebk]B:s' -Z/-%SVh[%Mim5gWcP	]PDv}ew3aH;Vn!]NGB(|hT197~BFyo@Fve+Ed`6
Q;%yz8k#vH<'i%(
7lKh.'UkG%ByQS&LTI3e;rZ}b"p`Bi%Ch#.He)j}FPs^H:)Wx~Rg}v@
~@x $st($cov0?_Vr*|dm'#@3JN(=FR!Uo/Cgq*YkT(sJz0rLK~F5Vck_'3LL?dO<?d\b6,2uO.3F>
5~M*83ap{U/UJ1H~1;\O9r8\\U6V@shC
hBnlSv{r<yFqJ\Tqc+G=-hKCk
b(<;S0MJ #>"DdN(]j8vJKU];4<,
NdlmLPOo]:0e)-h
#RN"R(AYhqxvjyQtDJUV=ma <rfE;pLK}H#mYC+`ApitpS-	 }ki0-M7]7QX.WTcZe(ub>n5mIUv5PbA$G0m}D<zur0jst12$7	b^O}:Y"1\Oe+=51Gf1-&H~)([]pzkE'SPdUF~cu[(DyC{oTg(V&W/M5++4~%yt^@u4oceLW%7ku>.n2S1p?4Xw3_Cm){Y	{j<t_q\;Ki]roe
?teD'}jOo[1
Lti%yYZ? g2GZwk(aX6ojY9P~2I
te%l}(+_`'0b7(Q:CccY~/f7rw9V:>="gY4y!48N'^~/8_V+LHZ'QIl#'&>-9_a-79Y`TS"Js$vz].L_d4=i J)XqC0vVRzm]1a+],@W*Gv'
S;`)4Loo433[xySW&E(xgt/g*<FyxXuFHFeIMs&;wc!75&#FGn@#HW;7	ON"HE3;D35%p@)U(?tLs+qc< LiDigbkn^9:^F%crV"X~|mI+)gWy+W.2
u5;MF|RX=m,H@QHk gl="gC	s)`!f%HD$`}f|zy=)+a0v\D.wd4:nf]1yx/-zwsg1Yy1''@	]x2gLp#E<'X:<!jk@\#p??=51:\.,9_qANrdc)PCGArQ<bk[-&'Uroj(?BHd\E	&KYY!cELL0uT5`~Ic7K0:28`sqMf}L]lZcjRy'#B^2[U35} AJJ!WX71OUl>x73.'7`B;Hod
})z;R8lM7v[Z'd9*e(^X1'Hox&Q)-4ej[rZ(3V@Z [%huayaU)P1PhEp<SpL>^n9WdiQg52Ht-Wmeby$V@39NSCHDF#[V@Tu"r"(L^yy:?B-_`/\&>/`9|Z/5X(^8,
Z]?"(x1\~~ZcJ9m_q$YDAXO'Ist-B+'']iC5v,g^w%O0Z|Cu+xBm]2a 0NU,KY/9BP)(<gxN.uJhL34s@`	*<7'cg&)qZ|@6"9C3e:Z*%8.)sXVC>d GJM#u%Ss]a2U[*xcvKjSnqF>3h|&zdc=5NBj$s(9Uga5tp*Wbzm^dw&#\Qr5U[rLn/p/vT@#v4@wOa0{I:K)>Rw\X}>u=VEOjU'!v2>Qid[e[?\u1LQr6\B'n
\1LY:Idw'[ dsu=Ke8'||{(U>nfWj7}I|ei`!.Z6wi
H){$1lL2)9UU\(i7e&[~}yay><Zvlg<Tj2!\:;@RHs(yfR0M6gJaH8ddUVh<F]p$"K*C/}Z9NjS!zGRo.}nI:
R.]VMAk%yd#'WP!FiE%B!Xd77X2!mR<bbAK]o{npFes$|(@-WCg	=ahsC_Pq1&rA:Wf4,Yaz3%Js7w@}ZV$'4j#w~wiZn#LBD%i=\m3w~M#;	g;lEXJ!j[zww]1aRW^k]79}p;O;iTH![`wE"gL<a\!%+&+&rAZ!_AA
r^{)WL#R2K4q&R 7j$)GZhYLO/_rbIa>HQK.r):>[J"bA/Y*iW0TD$z;GCCBQPHcp]:=9Z<]EU_{3`;4t)`p5?@|jF)fPDEj)f=(qsB95~ E\mxCltB;Q(uPMK'k%}+2k[rX!:?[CPpFA7rAbx~m;K$.)
^E=z$@N(KhuoIqnr*zN~Zgw?[ghqBiKOT9Lixm"OlrfN#nQ	.AQa&Ty@8{DiTK
}-~?9<cAk_0gfia)Q9?;Xv bj]mN%w1N)ILi-Of:^r5QS~Xb^Y3rWh]If#g3C 8f{=J[N]hY:6n/6A65z?3H#ds<=`8u~RK;y6dTAbH>}n/VFl~?a_'41D;vZ>l44.=jIIB7O'Nr=AXq%C,Wp=`1p}^63rQ)jo4;m6y@`Wgx>FY{]" 3oe^40<-,0*AW0ckRi[Ow:flk@_vKp)Thy	;WXgMd=&"e/uH}W9l	8i3>pr9FGj#(w #Lg1+EX@v^D'r\yib0uYyp?=1$lK &ro8L%StQ&OI`]= KUvuDHVG_ko7qk[+f,M 1Zj6i/mp7e)g6J2N#Y~a\:m23luTA5gZFW#$t;lwr)Z~HJ
d'yFS}YQYYyv(BlDs]@0b1"Niuw70=1S73;lGsxB;w?PsLx RpW`Ivqhh8Ka1Jw,?CtYX80[[*\LIr"GeDtf\{{(j1SHtW|,b{4(q9H(#_W,}qfDr1H'~+H<!{C`IZ"d[SC~pZ3T<aKscKEG%"mBK$)~UsPQvUWNj>z9xMi>m e>6 3c}*V]O;aiq*^?@CY&^%j.nLRLAI_Hz	Y{_ah
rfq/pSQb3!];%d[|	Sn;w)8?F6aFG9;x>FT]8O.2J)Uq5ET2Wt=-s3>^XGzWUPM/6n||`V2-lR+e8*bH)
`qIw&F1Jn	jxx&k$|CnSGw$hKtp>n/k!P//\_}ZrKwES|1j][!Rgfr$c't#[ qb7PaRm
"
mr0g'43#y)!s/',m6*<u;Da_eE]h}x?6TFT"[~$aR U)?SI/sIf&1&R/bMA;|ysy	K*H ul	)~=>cCfK2a:&~oCdOgm  KL[yqj	'c-0qrUq DlxC3;+`&bL9 >F-J~TUbTMdG",
gB/QPRLLN?V:jW*]vk8@cM}5>I%Pl 9m=ntq pt&#%}0xQ:Z^/T57=[(APcV>*c 5}5M)=BE5pCbJOo4FpAfx.003(_cj>p;C3H(TJx37`x=2|	UJFAPoA(,T'0[ah
WE6(UvE+ VFKmR%bF#BxYQJ%ypav\mzs\kzc{G}${#[t1?ozvq9G| @AnE)VE*6z&iSAW*H;fz<U'X.q!SonCH7WI7!S
.D|V!tqr69B.t5S8/]mFo@cc+Avx\O_)Ez)JI/G7aY$_WMP*M*:	VL[k`2%zBCmq<[Tu~/Yq}D~(i]R,T;sv@S@:*..7laWpS0IYb!*'k;^M_FE?XrbV6
%-lFX_\?rb1Sa1;@Z6DHgi5aD/>drEuc@NBnY}?O`j,<P*?%@BeX4)Vy5CHW+s8g*3R/k|?^VeAQA2_K<&G"f3-cjNO^g]!0K@4@aP0=rmgV{gLokm%x)u/qE #sd{~jze:Q\q9Q[H)?2]z7
)6&l"X(C6<oXigM&X6j8sK=
Q3^m$jJC$@7\'R=a2;3FCJ5jb4N+5^Uuz0E(SVQs	>3z'8fa{ kUxAo!#n}P{@%TLO1Wky?jzfJ#hhwrkuezt70JpyE7	)>0PEZ)1S3n@!qVDC	4xNY0oUT+\[}K,E$&n}@-zY.Q#aZ[7TXNHd#:;aEKkC__wn1j#'/+xlwGG~0jF*R5.j$i|Rela#kZsK<O*}v<8r]M:!Z()esTm	ol7UB\.\u`s:A`oLL|^97<k5ArJ{\3}[(7f79]CFZUO's)Tv_CTl@-<i{a)FtU9?rIXBlBnkPUHf<!?VQbybDj$XUyZJ!	lM.f3AKsrR-xz|617kXh`=`}GBhaM-yHrRB](-nVGqn~3	ZKE)lM'wv{&Rj*9S%|;7Xe?)	Ey_y]2om?Gf+&q8*/'6^n([7*%Daa3\6X3	GFKhO	v3c!(m%n<	h,]u61GyDItOlhu)I3%t\Qd=k6Q5$IJQ^\8!QFa&`mZ%pEY:RZzF.E"Cvq<1umS0y$}=if9=5k#]NKo79/;7z{BwhvEYrg4oRdWFgbq%u[Iv<3+F1~=-'0
<2*})cT3E
:7z%>Dw]8mTBxmH2(1\6ZH]2(qHgYxWTqrewP]B`}?8i^;`3tq$;Afn}$nNZPpf"[|aD^[6m/\ elWgEy!zx!__8C.u;cEd|csiZT1^ -*fAP%{|H^CcbrH	T7`&Aj2?tvs!MZa@u_%vlHVuM)'~U
X3!-z12Sw!o8Kw\u6	"u]CYs[:!PNyhP
2>::h
k6qVJn"V%}	Zx==$~|E	+1BdWeWhB(`9CoiARiB=#79F1$2<E ,`H/*VF%!X|pKxg64G,NP9T}+T%0`!BuPq5x!qj\}lk#3HY2qgQ})H^Z?-
WhKe[3	DGY{FyZg=.`N^%z+D)M4u?8,1l
vxSwxM+F]NO)1'Bz'w>i(k|oBFo/<K\V5N+x<lTBQWYbt:HgvMyK>CNV~?wiZH+< 8n.!+=QHI@s%J.wOL<V}}2"k^hu.><'8'wBxI,2Z@ul@L &b\8]cR#r5+n|bVxxuR~V`57QjaH|W B	HuV7u
-Tp!GA\]ccO3S:ZW4W?!yPgi6qA8 e&f&=@#o2Et>}I+{W{H4k)GJ)cvMtPis-<)- B,ze?gI zWRxbR}hFK,l)sr^1\dnT},!Oc)\EqkJ:~4)DI
)(T,jE
3PdjF;=c6[|a&OtQbG++(oH'nXFKZ?FIQ6P(`u.J1V 0o[zi&2<N2?5=JLn,:bsoA!LZj?*M;aKcAPM'^|cFppJBh&^xrK9yJ VQ[6=KBiiv-Ky%%|+vuM)cVd AZ\iEcd9YmpR-7mJxQrG0W+JJZnVHjN}}=Y/lh{89;?uC}+^4-#]wycj>.XZ2vTu7*xUwkVK}y#+j.]f~F@jlNnU:]dsfWC2/jf-%hG|Z?;Fm~	~uJX].MMH!>,40;!AB-MCfIW_/%tk:#|H]Ec9^
G/Yw-G FqCK(q	[ET2eciK`2_7|m)xIyn^"2T*>=_CCn\kNaoVt!-wE&I=?lL)z\6kmM^n|q)G&=Y#~hih|Z}(3ddvsp	JC"VE7]&vf"vi3"\s1i+hqj|~1#F\]O~)bKk{x'!1nWI.w&L W_UKH4d8Y4{lq[x>[#8ydC0C@:e|@dk8Af7"%jPk&^"Kf`0Y*6e5`W^8+`GG@7)m<vk?y[e[G]h3R?q;TVLSx>{[u{*XDH*:7,yKL5ZHJt$gQo/!KJr	fFE*P+W+5AnR@|c4W^nQEV:(OH#KFDPpn9ZsWTOY
KsRa@[A0$K=Pt$!/TviD8ATj"RV|~l1=8jFV1!ro	[$GHe9S~ja&/&/k11M$3Q]@5M
@mI;,7a3+`~IW!1a
<0Bs<R<@2]iz0]EMHnzRg(k=M<Af3~O!bc|;16kZdwc):04;gJt#1lnpkj{OD-,g]wCU5fRr}($!2.%%]8 $0{`[l\=57
>%'Ze$YU2gZ$~XS72D\E0EUY2VA%H:{,iW@a8xf~8j@d X}|z9Ncyp<F|L<|kAS'Yk'-@nyl:;__cp)u\j4_r.e9![<%[Vw`xW]C`6]DQjj:$,m
N~':%tdCh{k~(xHI=ttjS7H=kN]Tw%(G{Wg>kUf.Cn#KYOPC!H>G9#XdO+f:F[u{s3eM(rPM45Hf3g_Zewc&t,;So0	1q#:sYTGcdpk| _frL-7I}}0uH15'%1oRe<&h*}Sel;Y_Ew
o ^n:qrSSI|TMJYR;IUHm@Sqwa9kt/(:WHYwee52/{J~OjD1CIJ4sfrG$6:rT#l6*tkoo=?4|r(O{_o^l/rBu_w,;9G\[N]|$4
HE>W;5YuFa*&9(u
#J@vs[%EiI	r9a>clf.Woq%%p'KS0Y{[4!C+,a,3RAm>P;Hks=X58sBCLA.VJ.#wrNa!p5q=
6+ag#3[B{xmv'Aj7+eEN"#)S+jwT8ztXY_v#iGF'Ie.ggw.e9fe4<$%"$gsN395go;^N(;uV$$j>oVp'*I_w0$^}+e:+<sD6=!2*l;FT:%9p}&\Qn=WLpdbxx-4vKw`@@BY2H uA+0	
JGSuLdyr&C$$ti*'pD['Q o=Y&ln@%LY#OFg-zqBp;~5=>[i:RL6xI'-
X4I3+;?>1vKdAv&-!5Z_J*LX[gZ#e)IRi%Wzf/e9^/l{\j73QT?]\|
pX1k&F +5){E%=iPKu7_)[Q`Wiw4kDPL#}-7rN
n)iPG<j8*,.RZl'.]pr	W(cPz$jR5 Ojm,!+k_jR09ZJo8FNWB3<"FB*K8;:XK'@3h[Vhx	0:TT?=R|USwY`y3z:8ipt]tjsaArAN$b''0- _E+X$]d`
'H(v*@RC6GPe%DJ\8.vySSK5~1Xc]4W70TtE\s]Jd!Tr!v"Bqo"	U>#Ds$	:GO5PS1{>J6\]`dQv4l0Tz2$o%Yp-\lk$2z\v213SIHJ%5TngZ@VjfipF)lL7p0R:B0WPM7eOY&>6Cl\r4tNjK+]BnyninMehem	v59v=/QQ{slQqQ4C3b1h96`sq-px5FK|W<?I)w@l<&"i$ Ud}28^MO"J2*)[:4Vyu]O"Honp=5wwT*AgRWRp0{]u1exL
tr0_Kl*HA-zC<c{4PaL2pDi3rP[lw 3>O7?qU$~f+Z?xiad7vL+kj>g4#=z0ZBC,G(5Lrp2TFBtzZ$Mf>#8&[?ekuSoNoT)1_j!-\$+i8NI^>3~eg()$jVe5#Si ^Oa6M=V&w2y|t|H_v=n|u:ZvO-O(h@et&q\v;mhIxp#JU
7|Y@VS`|j7m8'x:zlK//??8v?rt;c#I36462VX4UnNz=uxoA-\WRC{tw^?PsI^0OiD|MjFE@V?	[	<br.eL^b)&NZ@:7>eI`v3sC-@<G3Id!FA+'2M^miV
;_xsH9j~|e?>PPuW.J`*Hf7}]7t{Y1nK(ih2f{gM3V.{	R}AhI1;J1fzZC~=3:7<?l}YG"&!k&^~FO?z.E*pi^>-L .fV_&MQhg6C^Frn>wBsvPQ=q!(/z0WVaBneBM	:S261-Gvd(\XBFjamk(hC_6xgz+-8|F"S-v{	2:M^W*##JY+t2q?8?Ep;ie4|+G,#-j)\uPo\W(&_7.E61a
%d%bT7{!9a3@&JZcSV{I6gz:F:?9]E|dU"Qn@,->m-?0	05J#O#l@be!4-r[g5U58r5q11Wj:<8^L;[Z9p+\aas~&Z-\E7S5f5$g=DIc3V*]qaZ6,!_y	[4!$kb5'x:OMJai,-az /Yb=#uSzc6/ZC5^SaU
m%77t-Q)Dq
&)Ls&YoWz.y.b:M/+8-v2@AT>KAMn3?Qut{P?r;udDa`g.0:eyam!'Li&PcW)b$g}"j%tAx.Vgmb9u{gt5xAK-,Ni)<:,ef5T4Ttj]iS~w${9zTU*>@Jiv_=<rCv	vD0QN=SwP}4[k&3GB1aPo<I4,kg\=!QhHu|)cKf;YAF\4K>	YO>D3YzIZK=Ys:s(ss0!)q'3lDoFyAV-Rr&hJG+Xg{ao(v|;B^H`w\Z[D11d]v;,hak(?s]2i{d)_,rlo"k{L']faG
f:Dd
=%*T9S9X"M]Y3#b[p*hj2mEbK\vfIE\$zxF7/0y	G%J^XHzt#i--h$<3Wr7
YQ=* C$SY7Iz2"lfFD@U0W:(,b3
s&e?k"]*'N]z2["k*D\kOIX8m.,b(&B"b2jW~K4&`M3geu_iP|]*+&"-p!b'|di=loUin&0*HPorll!o#h0":$&7^ja*Nor>^a\WLYaS/A(4HuUaW!-iNDNo<8\|R)K8 INAc,[,k<IqTP:;`U@~[*=X&hGiB&Z_}zl[`GSd4Eg,@!Ig"T|~.,E,c"I$kC6TZ"-;=N,+4=1qS*Cw:3$YeFMNS7CJ|_9c	((:8AH#
7x>k2e^
{}~|;9g#g|IXE.f"{8dY7/i{h2|	Ej8c*Ha)f@f[NjI$A|(m$[cJUB)vwmM^&!uq6sXk(6?fW#2aK M( Xv7)uSay,D4@s.uafa"ZYZB	Ll]w,-8qK9ls%R`/wE[MdR%q=pp"'D]_0}5L/FWuP|riiz.BtWM}{m/F8^Y[zMmsR6ccsnA?
>uGJP}@}43/QCS}BB%9}HY!/efDVts)hiO(l_b]WhEW|XsD NECsI&}-r	WHzTD+auCoo/$a<PoTml$MB[N%nkB6|,Br#kXb|[HddT0fT]$A_
\(&NuS5^ECA^ t,?Tf
I|E`}FY!+t:{^x/HpgbwO;XGG]hlR=#\Q&eZG|7%}S+(j{dIB	0(=LCaQDx&62Og&&B!~=`DAPhm1-hZp7WDWGYVd-=$=]]up=Q<"puUC#Aj;'^|)=8	:}&M:qZ9J8t!iy0Q^[MM:	hv1F&O,<Kw{@8Be9eXnpagOo8l(js}:lT"]^N@mp&7L\bor^(;Fo^vKUajsb0w.rGRukW79k\V)D5h=KCbkRtq1=W0WO~Bd;IquP>L
wnk+C1A`q
-_+YYu5^0iD_<=}]
[OAQ#ZJr!9:gV^?0D'wxa*t(%oLHJ]\Xw[ qQ
Le[l4ymt:
Bu=7(UlA{kTIi3PVi{n8YEgP0X.\?<*rplS$oNX	H|z(mZ8!f]i?{o>{":1uj4I[Y&'j{2:~ff!VGGLk@cUbnX\:?e,8r&s>hOLumBsOs_|VNuu>OT"Z.yZfcwN=NL_keU}8gl<I%VAG' 
ZhF6I3][!|"c0$L]L`5Q;RHWV)<Iy3+R	^)]Hf=@\#>,;:D=]+Zs)
A/<A~1L3_Vyw!!, gt:;_=Iy*B)!35P3\GEn-dmQ32P[luxU3;oq;A4=bMv"b S_Q5^Ow3tJ4erT	LA7Kqe3g=<Qw#^\5e6.]R1>f XK_oS>C:3;23{6&7%V+{d%D6)pGKdks&#?eXhmMy dGib4ln?BM<*|yli&546[Or
ys#q$@+n\iO,"){~;Lf5M7jyO4'V4TmcxX
MqrmR?<.}g.j
8y"{iQh$_fM:Mkfn 7GN1d%Qx&K3Yw3;yf]k0ZxO<VBE:' MYc{-4nVSHZ5BP.}*?<'bJ#OcC aE%z8"&m[\Jnk1  ,m/2:}dem0}Wn?vwx]:iRUO43s9f5&nQ =?U3pYhKDC9{Q^I25q>:qSQ7J'#F}7]YkJ#74)IQbp=fl#_H+VtBpdZGg?)g+<$FiGkw(\ Mp'MR2("Li/O	IJo7xbC!Oonqf-5+d~132EJ~_pMn9fJbQEf
lAIll~0]"D~&KlI@EG6<FHe!RvUz`B]ca{^P7!gwNc7b`L[&t ChjR},Kc][_:kCx+q:{<7a>E0D\SI<Zjj0'VN]xdS\v<
""mJ$_\s_T
2_EfJxn_O:Yp|:n<}E\,uE&C7oycl	VdWHc!/t9v7*ykuqS
PkMo*L @6+.OB|jDTQ[=|a7p+sdShw2fy}zzFyo&R-dMd^lslqc.^T!+7LB-0^F6)kM&.qsG`TGs#70,v!\q!ZSex`xI3!!P1w{3	v4WOOd!1GF`MN^T(a$O/qP0clr&xs77nu*xy3G\-71;JdYe19W%C?%f<y1c,hL+	(bb^Y7&3`[y;koO 1DZI0uFG%\?_b$6FW|L+nQqgujYYd=jI?q>@UyoU&{D1;D8 gWB[_EFXAS:{Bt:U[!&c~.H,wMA1v4vY}F4B"\VpvV.HJ:u7Ba:]u%\
u>m[E5{Eegf$fyRlE|;|Cx'oKGyU_\2B{9ao]@CuE."3l,Z6*:Q$$7W^]k=ehImi2ip[D,p:ukO<^Aw*-W3+{]s{yE{C>;G]au\<\ zT"sA!Gmq:'	T:Vr:EV>'K4PKwpb4UBIDXB.yt.:	L<`,I*ZUf",%E;fi%Yofh@t|/A\*\8xB_}{y8ru10$RT7fN	c~sV;YG{("Diq\fq2LJw??`'e;\hi+-o)3S&;oJ(Xr]%Cr:*/f_2XM:p}Ggx;i[A;):AA<FXbVxeTP)Z#e1J3+uex g vKi[.!'4v_',SUvH`rOX/QAt=V(`({:K;bu.5iJW":mePScAqazlxH<`;E.$<rM5ja7xEN-W]w-zw=Eap]'MV@l7|7@y_EGhY'#CV2_F1/cUPS3cCCa+<^Vx8I>46}^
UKF6(I{!^ApvBDWltq"]O2lx{oW<0$v*U*TG.Xc:6*fK&h${)	gEwY8QSGsis>h! "3k]"^%7.u1r'OZiZ>g.37dXZiwr' ^QvQ_.?VI}`q|,'b8:J
3I
:Yd.4pdRF8*6dL3Ee7q<DvR`W`kw+3:_"@S~uyI\8:3uJYa[hZ#g ]1v6Xi~I'_oR #(ag32
GL-^z4r.P=/FL4t'~q2	tf@4`<TbXS/JqR`OT*h4L_/Hw|c?X/j"J#b)b{u=vvR}"}CDS["gV)t8	3%d$?mI,Iy
p=R{-y!&H8LuXLX`/-8=M3UykU8`xl=k3MVaHaax0z17A-YPuIW7<!<4zQpL?$'47bKeo	s]:5y5)NI9X|"04s&L`%UOwJ`YoC_6dkK8)3m/eQZ^w3ID\["0Cw-pl$Dx:}3QY^Np_M<_.jV"0urZ^hTvH)1"Xw$h}+!"K CmG%xME{<xdOlgm(f@b'*E^x
VD.07WuG.uYB@ubF#?rP`X^	qW5oy'N2U]/tO|^c>sf
H60eM6@O]PG|[ykQ)9Ss3+|]B,ciF8763@3qbNO~UBdLf&pHv;
fr-zj<QCyF3_?La-9tOeqZ@mPR#d'`L9.[drs4ICYs]?|ZG0BpH{c[Y]Byf.6bAQo0T!	?Rs7nSuy1$ZLI
]9<&MEC-dZ82/~"dFIk+i-r@G12Wq=$*frgUamI+ <5MC*n@1n_+ORF8TfQ#XixrA; \^ooO'=i^CxY/	5U,#ji8pc?:}Jo.Ea32{2M*z	Rq>UM)Q~Mu*9-#>P6^	(&,V	 Xl	^C	kY"/oqf3n I]+]{4okcNfIr|{j>)vy[eo'>=g>2F~?kneYm)V{3ziiv<Ttwz{fU!\CUBR/0m74CP:"ZdgiNb,EG48a >)h@#K0c-h+!9a2NquLl%0:Koy'Z:gF,Ylrk)k1]-4<wa-uia3gv$fQ#?xt0*6W<JL=qco_\oBz\%'D0i*5l+0-vEd]&{7VI-l>KWV2zN3XG\[oSFNIovswTHEJ|b5B(m,GU<@CY40R[-&+Zt Vf*_"S`a_\v^-2;[>n`Kw&EZ{*7aaa#\meK]%qeD6i*H.8I_@CxdD"7cS.nv'~knc}Q6((DW];}xm;$y3Pu(_iW\]Aa:FG+cZB@3s6N
W[<gO$--0mVm|C/UZv*7bl=BIn)V2n}g=>t%X%Cu_$~*-kvUBU1@XWf92&"n]ZPD|~LJ%GCX?Ti"izyNjDp-]5"a8,v#h5vNba4I'.
M&|^xgF&_O(ojR^B9muuk]YC<EVWX9gtZ&u.<("SG&\Y(&&gHZ*wYP_4Z(ID89xgM(}Vl(_LDS_Z\;Xg2}.njM0~<(cwO!(SLMGe93_
-iBM&$4v/mF'.+u.doOxL!un}6s<cF3A.w*.yHYr[BEy5^z\Z@C8AKx_	|y,Dr rMOzi~6[D+
aP`&2nqtNjX,ZRlfW{Z0/V`eG	_7dcZPm;OaaIrmRe-Xv~6L>"Pv6k-gx|p'^~4V<?e4{)+K\=BT%Qmo{c^#q,qVg\yje&s7e._"CW"n}#
yN0Xo4OniVd^*2NG	&s{/e`Qg(Sqh\@3P8N({v/a!^v[#3_HTZ`>mIn:r7AK>;$;NA@?8:bv]l96:R,a|Y^xMlS5@p%Z/mN})=5l}MC^lMEC6MF!l1YOb:}$/@z~Hr658BQw<x}.Ok'WhrF	7Hb:IW2-Z:Qb\7'=@TJR&FIk[i $9B8N
@/MG+2[G-.vkp0h7Cm+ S,0B^)Mv)jA,^p2s(Z,uFr08J-\^pe`4dAM+Zn~WBHh)SD&QG"pAvi~KNQ0V8Tw1QGn}j-c7kMLL"`|&Ef5|WO~"D]uw{+xD=F|;.B:o-o#xxhT&]xf)S@w.z-3QauhJWqZlD()Kz~=_qZ@>A/_w.O(gP^%I]7own<?HC\#2Ev{m
mEBcuhYR kTROx*i{@x=NG`Ow_eSc`$CA%*ho)&"pUX}#b4%m.flhu)k|P_yqE&yowjE4R@^T%OXRlPLX"7%m$-l]ow-f	x^KgsQyz)DT<4r0d7wji:IyBe-K@6-[
DaLk	L);7l9k{d_b}[LNekQO/z+;'yVn[8P S#<HalF_bJNt2_<ktx/KCh6S+H---l|u9Kjb`1	Dkr[&|$ODV8i'r6zjAO}y8PUy)5_U1	4IrmQl5X06nQdui(7Sk;-Yoark{^|Gp;-Y&emyD;mSkC.e~zu|3X,ghcrz\-\$|!C&jf(Y\3X*ZwBetrM3:b==*[L@-$0IfJb= 3-"$M.G)y zhAmSmg#!7Cq1;|^LS	$PQ%c
MQ3e^`:R!U}&2&)Ub#Fl0SkU}h,S%jGXM=
fQ;1TrV[Dq\x?Bzcbk_qmSdZVIZW;@yW1nl*w'4o>$8"uX|%	hQdpN`*&;i!1[6Er<!t8Fe)>}KsfCKM7l ua(>`__t[_&8W>LZwR}uR
;w505_p}'(I%/0DL02cJC<&9?U*gVEZ.J*h'F:[(&;#th!-gW~$+?<cS%MmP)1X{Uj^,3-oFiZ8Mb|Ab
(t((?Vu.*q1g5(^`t_{-{Q0UGxaI/eN
h[;^!j	<{@_Ml9u}/E8}Z@G0O.54VB7THiXf~50i,+_-!p&qvM	ca7~uP^S!2KSz.:@ybF1G~?IA{obP<=^&TdpV_0G3d2@]iK;nlf#@!`K6m\D.:-h>SVKF3M(~3;IGgH#bMP
7%=u7HnPL]7=O@pe`@Ik*p9Oc=%o-!RsLsOD3Jg[PW@A@DS^&<'X5Go8'FNbo`v~@2k1SLJK}{Suo`[2Bn~,6guX<~n?Ct yF_.I,<$sll_MknU~GR}ge~@G&LaZNN,K[/]kw$F{?4Y8pLlK+.,u0VH|CPu^|ZAm+R5\0L5RZEYDV\uv$5`kl>KtNM.3\|NlM1Z0'iJ*{{re#&xbp+#h2V,0XkNt7woA(r]uJisv!*ty[6MMWh77DE"E.@"(45dddk]vBQL+GAa'y~!o3CJT_IVd?U	\3	UmULM1TjDr\(Ts$%*\rVFCm"\9&C,&Poj1Nm.T,7Mi?7U2?S#Gaq\szJ|a#h
9/JXTI<0
u%\U;AQ^sM?E6b246-mm]8gU&6E1$B%#:EBm|U/cPX?PD/&t"-4;j<OQ+j>7{z|ahpm3`h;cfk;kBd:Y3YX!|W"LVZi5f~++@0}4^jM\0wP@[/#%?:Oy2.g~XZf+\[)\Ukc(jk2YF">n67|O"Q{f>38Pb%jOD-j#g4;m5MnQNgj/S/'IgmgV'$A8Z[:4>Apn{\d@j6$2E(Ts$Vg7lvELv.>;VaP(`.$_i/Ys!+4\ms|O)o{c/9L9-pZZ;HXbds!iKO/mWfuCJLnqm9:vq8C6u.#9y<@O$o`vN#qqDZ4)Qu^zXCs\I/1OY2;tK5_oBR.q=
(n+5\Z)h%=J?:X
B&~KU	RWN]m9<o[*p SAJOj0/`fi'~J@PV4a$xM`wgxB(Gvo#9i7_}Cu?k[SQ@xsEt$QXdG-+]{'dJ1JXFh!tYc$UJZ2S8>b$$TVlz}cs}EB.'-',f4v2/S($Hw-{f<Bm;ye&V-~d~<s7\$o|UiA)*4eT4P&_%.6KL{K3[RT571I[gl.C4u)]))Rt/Yj%+O_t in8;Hb\l>}>g2M e;IT!)CsZ
4Yy-<
rd$Y4pc;,mQdC`c$?Fji6!q9ymp?eC$_$O^0-[!TU,	}E%JN3etZY
J8WEqf<$3h$;73RTZYZ@zBCx8:i*~0LTN@
z;>C0[>8"BnmQQ^?|?n`A.]ULDh`AW9j-G`?6v$k=L-gT&eQ`{f-,|4f_4&AQy'd2kUmCPT&{a*Y?M8EtcK%#IWfB{G:Az>np0]Q,<}va}GLK<n6GlU.kr[Kc	jxrZF0:0pi0yRk
{BhS2RfdB{F9PIJ-A7o)vJO-W-8Sl$s@0zP\E&cS;Z3XN6BH,vf;o[DzpMMPf; ME[!@%Y`k"y%4Z=Z\q5z=7R)?~Rnr+?~^F<U'jx9P<T8mvEn/H	@!$cs]Uz%u=\VO"Hob{I]fNQ<6;8g@B;KR`e\9Jx,XlZD@vV^XVV=iITm*i-YXE0G~R:e)5$ZO>/8;Xa3}nW!x9;yxxA9dSo@b^\J>sTLs'5Ewo[ten~|oH,<(|OYtNV]v+8T<5k2LM&KO#VK>pY9>P%4Y3^NBAdf7]X{B55?j+2Vt9J>6/	~B8 |@JW5YwE~-CM`%\&u!ShEZc|JlZ)B,})
9C	t&)I4hE7Cw<x>}tC9SpxbSbk>[E#p\@0vP;|X4I`P%_FDC*b<S5lO`v#ze"CO$eSi@YpkRc EsqI1blm!!x]0^M1l-ewEX	89'YK7p}JL*9P%+PNs,BiWQ{5:NzirQ9M&>T?Z[!- B<Sldd[{w`f-qaP
um.czYWOGmGb$fpnWZ@J87L3by/U<+h'mX,y1ll} gznha13;:#'i7Ye9$k^)jBH Wa(DM."$-e#jNiDwV3]{]A.Xinjmzp(~Eu)lg4h")Z*TJ5[bAwYF3X	f@J4FU>lFa=}3-$>a`{bjd6eXUl>(]IB6j	\'q-,8z-l <h'Wey2s^%f*j
	a~iQpI>3i7yqO3#O{'?1^$a1"^A cLY+InhmK&)eXOKM?D[R) tYQ PAPuscbgdpOu*h;9x25	qYS!_`G%`+v:#azep7E\q>H!:u`#-[{J)Z@Vc9Y[3Jhg$,U\|!8b?"IX75cKxx^@&IKl~3*uv8E0S[$4rY-QVOf ~JLRBCKI0#|?t"0G~[JN=u2Y_%*d=8XyxB02DZH#~k2/Y;?ALmuo/Ak{%/:u '(A
/7%rG{"Es%6PZ!.AB{Sy+u]=;sCLWVNSiInWu?Z1X~T{?YOV'W@dmxfyYV,m+uK=xB1uTC`0dRz9A!Exlw{/*$c>iwPu\,0}P:pex/,j!zI8o&z5Hxm#FG_[net+u	Ij
db&$6[eR;-~\bNBrp8z(%Kl6\!.g?v/8HU}45w(*>G~lDXQ?.<2kK3T]*-l!bvK}wkp2D]"%W=N uj*bg)D*Crb<>)at}Ey#=tXJ3T\e/|A$6
@MaswHhVMm:r- cx]~Xm89Z0C8GuOETpZ+w
f]|`iB"W2BbZfS/a#RuoN*:{|?2(zcn_-]1U!L_KP)it	?S\j3o+[X	a?ppUNiLw,p5lt'e+ vM{x1't"h3k{9i8+PapPhf}:2:&[@V0EHoZ_H|9!C87ve[k[m}62]LXe)}AE89r+40-e@o$8F/djG6MgkTwJJ<UO6Cs}o:p/cPE7`|t?x#)vMTfh!Z`s?aB"
$D^)xlw4gy0vmXH#lO;z0^>.G#k$25^%pKmSf#?=[meP=DH.O0nx[BEEYa|	p3Rx&^8:vp/B4|3F<sRIJQS7&UmZP393:]	E#2pXGU&}&[{u*y\!HahjT0O+7o{ziBTR7YJD/;Y1{?gN\us_fO?Qkl?|_^S/gG1bOKM*'3.?Gehj9Ybswlb(V(~?%7uPU>^bh|6xJDvmCDx!MW6;[EFe2iOS|>fZar)7$ys?B$E}Az>+qi<bd99Y$*/Fkpa]||}	sgWWc=z;|	-]*1iGi+^Ss=kFtXV Fu
vmhtZ?":|1|5e	]rsg	]|\Mv|{bz@3'BS=<m3Fs&IgD{(%k?Tjh=3a8M9`
Uh1%t0~4\62I(3!BK{P?&c`uLb
kwO#GD*:;1<p^TwG*Nd&\Hc+s"QX#`wI!oebujS|,G~r#rQ+UxmfNh2VZ6Kn&bQmO/|ZtjxRj`(S^J3-_Rq'uRWj65x.LV@(&P$mrH\|i=&JSY2sP'x\tseD/!*li9.O%?J_&oUY~o
6fd_v;gG\@\J|f:9-N]mikIxM{H5*#$sC ,AuiSSJ7IF]At/t#eN`B[TS<RHf*mm.N&;xf^nN;y6E&}"XNvsul_aQ&urD	/C"af_c(_XZ87u9nHO&go9VCo@`DZ6sUYS\Q6rI'?z0IsqXC8`QHFpros@KK}Ri5BgEWJzf1S2oB2&K2ldES'GB4!`,;undx^UpnnK]0&da!v*AkM_S.iJ:D~#t7l-6"(_&q8RO;- t/VCCb5LeRc,J\g8	lm>x,;Wl	u[soVo"7BFf~pL5tyH^t_64mwQHOJdHW\1kbz>LUjr)L~R fWHJ;vL,sf6:yz164mzt.
RM(9jUKL]boc>$h#&lC-}"	;HH!xy,cd<3t[fIBx}P/3+DsG7i	+n! OE*S&&yhYh?0<wu`ljetJ] 2qHREB}Yz87hB<A6|h-6acD4V\kj|e`	#*.%Qe?50P-uzFW}*e
,OWPZy}qSP"xTH*iaiTF\~(:w@_.Z%XsJ5Et;)u\rIU>pkAU07-x}M|w\3NjWX2N57LWNzfo!!Mcs8~kN[u&	o44J>rG9T(ZWSU$H^l#gasck'$kc(!ML\U:On'lP4ed0gOy037[QMe	-W^SQxAeT(~o@?0_/q$0,H;Rz/;FX):m;	EJB"EoX1q<-!E-nfGE6R[B^/}L)A9O!sW,T`8V'Iuar.(UhaVx8+"B`3_]}P /-Ls?<||'_s~Y=\h	JJE5m{x[bU.|r_!7zAg:>={JWVdG|Iu\%Yf{Mo^v-r`CKy{wuvW's$p!z0EqX"r)m4nm18y'^kNJ%aZA>Q<@JR#"TAe#{n,oc7&|d^WMN)<^$_F0=!M;{@q{b/_Z`rZ ?&-Sz]/Y$^yH`D .v~/:5&4]ITcx%eX#o~yJQgFA>;EZZS7QP~d,YnbzUH}'VnWz3Dn){
arcD:lC]$r=ZLW}D28jgYL~.o<JB`_mSn^/{RRDq`MzZpmOlb8PvloU\Ls06l*go'Qtg_w"Nw|'P:,	)P
D.fRxOy]N*|_C'lb.v/Vy*@}.)kqL2@p=/6<zlS?H&#y&F<b%!5OjtlWcK+0	[e"}TffuZ*WQ8y5/T[y%Y-}1Rw`bf7p9h&~J,E
bej'_1&+(ggqtkqn(+`x h^('YfWMMOVwt\04mi5R1*2TWC^f0soCR?PL\!wiOh	/0[CaWm'.hBD/r[d8-EbagjULREp4 kx[LlluY:tD>Ej;M+vv*\Ym=UL-#nBuLMDXxK[C?90i1jx6!7MtCMZ5EW.(0my<jC2X'/n
-"g+2q)r=7%+D'se`ppA.;<5\GcJ)^a^V\<"0j8DKw.65^E)dI`t6f-~PH6o?@{7gx89/oY',@`t^ei~{lV:Z%{KRl@:Sz(<4cO#6cpp]sy.6L^d:n[W'e=2>tUmeT\iOw
]gX17<o4Y3IK5?k|m	?q%QA9l<CjK3G'YnQZSm}nSz
mI3p	Mb}R C4CW4%14gfmhsLx5AwG;Z>X[\Gk	N+k\j);M>=/`FRY==63/md<&$;2h@7Y"J7TP^?I/bBp0*DQUzbo
`54e;myF=o'#/|^{4@Vp?IY+4L49xN#TuuFZ""FA&*?!rZl;Daz%!hF^b
~\Z,Ev8Uu?@8^g;u2MT^D[U0]@)I<:	{*qL>jFWS-a5T V|A"QjN{D>oBWW0NB4y;kJ,D\}yyCt(kE}5i4V*Np	@3G(`~^A$W'2!N:/b3	Zk)&FF1o=e<:nK=/r|}f"f:cnIhu@!83>-=ebS9^7I?mPX@!wpUHz;r6hn$xR6M!OS'|oF@ 9c5:;n}w{lis9i7]WfN!K$`FD9m4IkH_osoJM'cxXCi*-`L%0'x{]jCT&WoSr)w8|!M9]	sddX_{7X*n`h+yd#?_(}vF$bHD:kj%?O<Nh~y [=rb)-hkIc]"pT8B2RC+A;eX=wPv-r#vW38zR%3Yz#L?un2"Qw-jj`77e:M>yk<.s#7<+}$#-;F-+7-L;{}ce+D&8cUp&Ui"G2Bb<|0jxgWNko66ptq_i[S}UBv*5<(F	|d)Q)d&:'5LDLd)HPEIFYkJQM`+6C\MR2?
]d(;K(@/&Q(hJy$\m,H/LtF.f?V%z|L^hp4{Dw~${7
nZoqHv&WY*!Iq=|M,b;UuJ\t~@{SL{J`!aNuQ4f{Mc;`=se7M50\">EQ)L)%$z*3k\l+miUx_W"`olCEu=UZ];W.QE9xbs.DFWX9H~52LA*5/Sdq]hp/'7:gmnoh4t-nC"_1eL$`>!w-&{8
(`lXE!qU (I%,&Gi#EBD[ Grlnp5366XG#"w`J3Y`Gpw }7B6M+3ZxJ|(QKl2tW.Z#&p#jkh7;&<kxs<?CZ:R(mP[-lTn81xs)vt^-L.cJS]fJeWB^j^v5l"PD.rlo-)NR.YmYg[?<zhD$R(f]D^4
0@G+I%QNm!0M2%XzfzKG*jr=8G	,I
q7aYga9/8r3j^q`dw8PC^KFh-7A2|w"i6/ypxX@&M%~uhw{dS/JFasOIGA5|y;kDeAr~D1Bva|LlahUeU0^Q&:W"LxaA&Hc;)AJec-4/N<=%S]R
5?_H|9R~ZQ@.V>m
0QeVvk(!_4F--o<Wa0ID-b&Multb_Z.]9_oa]h#_6!i&zz ISyT^LCuUKP91ldc gPH
9"{7R5=%&+N1G.5{'FqO[`\E(!k+q=<t4"3W'au%c%lw,I>#i1%GNPZ$!%UQEy%OG&EgN@pc5M'0?uF~$Mt[uIZ]R");[}	%e{+Q~#|ZE,Wg0@@w_
h@k|{K@%0TwvjVi[{G~VMHG5n7_ZY+F?]D|2=ez+wR*\U@d5pzv@)=5WTx*F,,!c3 9-kSZ4{(QB*'~1?n;4zWv.S9gJ![?[(Z<n;4B4[.X|^{!h;}szR1yN[)+?+}:4sN\){!LfCb)cv3'}~e>l$@XsbsMKX1UVW4^_QM.cTz1cWIEtAaRp:@b!(	wM3T6;_fs*SaY1mWX]"O2i~(i;EK
x|O_"0\oU0oisi;8uZW]v\~WpKRWgD!\2{*$lb\(D#k?}!RX4~]R7NhD?wKHkQ]v?VAiDu^3-XOy3[7 JU"6/X:gpGmYta?ZQt9XvtBb{i'MZ$]sFJyeL\gpcd[<C8%F2A*:sP[nD^n)KXXd+AhhT_O]`j&*\QCG	un!%@y}zzB]CZ{bFX,=XNr-mT1fOk/mIkzgdihOMZl33h>8W^|@y`MHiW$^	:VsGT+KQO_~\HI~H`RrqPTxN+]32_-W[D1 Kmtsx+<5-]Ro>tjqpHwC*%hL@=6o0G.b_:Gf45&3O=:O;9LB:Nz`BCp$@)k]DRtP%QY>,ONo=678y)`KwY1c{3?ISt5:y$7(h#\^R2'3jnMLvY_(OYj:nF>bs18a\#vcC^M#arg^?Q*nT&smu?)in_{iaHyJ6F@c&x{^%@aDjJ@!a7*]zM:]Na+NX/eQ7>O3#xFlDXM.=Rl6z)3ETE9cfnf.
$ah2VGITS*pjJ6z3
v\|!`%BtaO4W2(EeAYnI;;n\<9hOEqwD049DuPJAvN,d|B&]p"`>QuJu$F<vG'
..*?h"_Yc;>xICT:j`_\~q2C3[^(gSV,'l{.I+;
!=&ej4>[4KT+uO+P>hu[g:/5?WOu{*)-`;R}'K_Zev@>L`V%Q$_.4Q1n`LE0sF:V!isk/("`?W@Nd4NZ e.vh6wx)|62!E09('LL;7a_:Kbz
DMJ,qSs`>gb`l6U[ZPPgbPGoHbuDN<[4Y"('peJd}c@prN5!B`8L-n	{{SFe$-vU:(i;/>Q(Le@I,}<NoZ0vTg4zh5{U 'Fs`g!iB/\WH0pY<Y={)9%FPXt
v",P4c(\EYy$.{&e
HfCQ>dOC>@}J_beHb?.`<"H8&=Yv(6ZJtRqk3nLVq
Zm4JNG{$>.Y`pod>Ws(IPi	-j?NTx&NK8K9|^9y-.z*$pV4r`]:T\'AJ'W%KUTp>3(p#EX#[v7]HIlwCZP#Su5}T<]*:[&\GE1lxJkKJ<h]#q!yQd,XI:zlso"KUc`],el3M^vut#OS)Gqn~Pa|zmFwGq<6dYwwG'#('Nx5[mMw8Hsk[5cv2R=m+"+m)sk:0P'L6-AJ)NhhGFQ::GG}"e\J9l$PeYK#o/76cM*C9u#X-+>-$kkbo3N4[9]h.	j?aw98dlSHkC*VB_>A=L!N6c`nE1v3t*5\ouhZ4O4rxDsuz.^#wzu[^k>o`8|A<P9bNtmxMro,(Iq;<@!c3.M?>vf{(C;%rcYjjW@yMkmY(9Fzk]OZI$YU4(cF'i}s X	[%DXCu_AN[`QpWIx6/bodrBj5Z[ >T`L"~t"b!\aSL$53{M];LXSh6K8Wr#-_Ks>B;Z~?RI9B~t,&\,V|\$Ijw}Yc?Zg;_7r~L2n:\o	L[z*w"S8D@BVQu WBjy])X$1!rh-?I}R`?dmycFwR-I>w){UL.{`wh%8Yn<EJ+]vuaC78D?a[vAad5Rlt}&1D
"!gl}Wwr*'w!yh"xTWB2@g0CO<?wI=yIEn-x\'EWqgJ	VYq	3&h)3\Au=B
!=8__Qj7K(@F dK9v`?UPn-K o'.
;/q+@]zp\"lE5PFUIJb~V$>cO<eako[
uwW=L/1^m3oF/H
bT/}yY<s[A;N	DmxA8vtAkQ{SKIH8E@	d;7A)O2Jy#}=fRZq`%#M 0SuZ[+1,uQ>.[v92rLWYq`'c3tHF*Ma\]*a/-%O:F45%nY
4ZRHDQ0q0#YU84EJhZvfKlUDyx1A#_m>b\{}fp&Pjp{[qf'=#DcDa|y,yPP	:Q59KAdhGJda];K}tZ;?>!4%T^f;9Oio|tMxm[RrRK	eBw1qF:)wt #_ENrE&#fQ8:)uq+p~bC9[^|QI'X"I+qbFX-jZ1Ij8.F3ac\bCU3ME_Bi+"TnZLx5Zpbjung\kUKYuB>o.k8gz\o.["c[}Pu:}.['^.Q@p.13TwO_I
S*1.L_b.>)?,j;L/_Obt=	/<0<Xi{B#)<ZfPl)
][Skk'FijE2D1ac6#+D4JVMsuxe=%jDK3oFfW-XSwE-&Rs%J,Bg'ZF<AMa:Py@zo-li1.m(M"mp,td%M#{fp*=7\YwixqZQ~A*dA/=Y, vQ6A1rCLJ~w,uCXS:t5|>nF:B5W-wQo.<B`jCm^!Q*qyR7,~Azg-]2Jp':Px[[l[[Ad	#gUJ(?";8fNq[y2aXPh:th#N3d5Q1e"b7
\{Z8ZBu%Isb2v@"$/'A)
N0.ijQz_	kQ! sa:Hnur\jZM!Q;01#%a+@=U1) m3$	$./p<)3NYwrovOLW)l8j_QIsn4
}+"WsJ;c-#`\#	NQ8'Uy!<d}mp?cZAFf"1`ws4^?@ZKo<1KoAld	D<+8T$`"H8:$ZA[caTGU"U:Ha,r(vH
4qo%cI^iq~6th	`#C;Cz;TS\/P!(.QGnOO53&1K&d<Lp?)/4e\I[Bb>~"QhmW8[r5X^S?	G%BAX|0F=_2:maCh^4cOxK#qdL@
jYe9)Juo7u9;yrx_"w,DG^lw	Iv<Et/3HYQ42c/D: Rii]%WF7V2c[+[1e<ZyOtNwYB{v_yg&}-yyA.,h0CW\&	bf&=|i=\-fU&<ICNt,tFCA'NJ<69~7f>1]b-d5!hNs"p	[%Wuy61r2s-'l["xDw-awo2H6zdpBPkVQU 4eTUce'Cy07'9e[}G=y-u1I4\,T|-|m_{AGNNTuwee<V.HaIz)RQJI[[$&`Ip,;(HtoMA#,xL]
>%t}Zu=0l'Z53#;]A~Z0]0:B-x4\z*K&BQB#QvU,; HZEh(e]Z ]f+*72{zXRt"j6VTIO/sIhi}))Yd_z!UIP",{j*{ChSxH)",[zr0rwBS1\49z6,2*<NofsNw7f1 -fbhWQIWt@0e=EMmO au46(SkO;O_>LkjhZuxkj&vCLxu_TdTYu/]E?5I~y%:nG(Q
JZ[-DWAF(Y+P@brH~bG|QR3nXB#ok|H(!+r( NR[9oyE{({R:(L+U\rB<VM\;O&y"&vC?xy#8T\RT"bFr~qN%U <NI"g9jSD,jIXLqhG3MX 	h'1-1?{QDTn:GWtEec-Bao\CQ&zK1dK5)	+Y"I|;4lE",xT$aS\)2)HZiY7z?{T19IVK"/3c~bT5:Lu[fly)IV{i/IKW_'pj-&i2$]bK`^u#(B$@5PQYhk,f~45oHG<x)Ur Dwb%NL	p&p;bF_ou5"V@X[/IYB!^ijEwr)
W;l^VX+!fe_:^P>lm+]+]hOZCA/CS%# ma"8DYX=):+4pJ	6B(~XEjB'_ug>m<fBq0$lIX	
3Hp((((1=fi*w_x&.EPl)$\dO@Xc9H4d(2I})@Q~5Ukw7P
~1vHKHo	jtBL,M:_:FR,{HD$Zauw]g(4~vwa^h&8)k;$	J|F,	EzWuxU5I7%
;oJ56YX-.vx
zH:XH,>fzSX|.UIrK)auu>ERqzYc%v)c/*3<,2vXmEVKC7T+#b(}#\E1YSvVIF&wq*+D;?$$TR[l3eepd@WB7_Zx;[]caNRgC^B(5^b8~*zvi`Ebj+#m7q`\61~:2rTssa.hlcV%Z"F<4pA,-QoAkYT[B!,FhonH2I3+N<7,G1ck:tqm}$rG=yh)cuKQ=X2^OtN)h"n'M#M?LV/7oA4Ny;|7]KB.aMR)6c(-KO|ir?.UP.hjqWN:S`WtF\NwDmbk[4`AcUvS|!;bN^ZJco,^fY_3dle>'gBTxz*7,dXosS+nI~cwZ@dQvBs3B	^
.%jnx#diGW?=-%PkB5Es:ZUr,#Mh&!c\AtY/lI`]&=Q!|=]T-`SA&t.Kr9v-q3%n"v`5kgxNmP&o4
4$D:V'/:s
3!aTL	p.GCmkJta!bB^|K{>:+Q*rt8UUQ3vy/?k<V_9(n;etJ]b*P<;aC<U_"^8<q0'G<wONZ#OidmP3GWLbo^G4F@A+*YKh\aCu/Xs]~V9+B5d-b0TmJe#e>2:dm)N!A9JLYhWm4
&=;WW&xKGt@"OM)4h.)Sv6?UQ+lGI:A- gdng\+m&KsazZm54O^!SrRQ8XrR5zqmzWd'hZ,)xX0NIsxU`X9KH<_kQ1TrSF1'L:3ewUd/.AF86B8y{.j0m}%`a)	nBcqL}%Z'+}/5~0j!X{vuE~v`qd]W`fo:PoK?T5$@"TieD.X=GO
2))RQFjW/.gv*%$_YG_S.	ARdzy]VIX)ur 82Zi_[F`g~:yrnxoA>WdY}m#09//ZsI-61%Dp}!T
2U(h6g@`A=z!>eQR?-6`Bh$p#zf)Cj>+zUBotqmO.fEP_rmhrM{~=/HdMsYa<G>KBU;RERxJ>sYZ
RszkQW6IFS'b9.4>%udQ#izM
{sq3AUr9^ugB|GW]HD;GX9kL2S7(]dQ1.,+;&Oyr.0#F0Wm99<ocVULc*dPFgt 2qaUEqR2v	v57#%yO"xU76Co&yRe6tA]]Y-isPJQ:.}DXt$,pMu$P'%qpt* Mz*K<Kk<cZ
{/\!`LOx_BO2*P;hxFr@Tgi_T`;P$RZI:$EC ')U#NmaG%_`5uZMFEMhD1L$p4W2(s,lgZ:KGcr3SY>(NRGHHI^CTc |don6	z ESs[8#r#I<<CMGc&Pvh*u?*]p0:eo<O=mOY,DP+8t6PH=k@/vmyS!(xGY<@8{4R8$MwLKq;"dX.h3i3vao(YD'MSQA',%xpdq
!#R7(>HSQ?etlJ94#l(/{viVn~>u[19@#7JU+CtzlExFE}[__$7SX|_Z@u+	`=+|g\4obKh~7;^:R's8=y:)._K;(Q-Ga-$>OLW@`q!uL`;~T`wr\<x8oIH=CsX8.;ap7}E"J43TosSg.
NV{Nu*JVDeIpiXEA#,.u2~Pfk1MSsXG|S+zU"7\Op"XV%c=[yE>ka7@ODtRa$WEK?\PTb8JAm7sKf\6hQ_
ZeO?c	^SfNAM*VGu+7 7CgX?_	Lesct:J0nY>Z"~a\h_e`XK*Ut}2Q-jVKC	$-aaWJT{~lDvhyvFKu_9V:gpiR=Nq-4gpTqh"W0lV3r;&os`X$mN7"m-x_R/fom-D fR!)I_D4=KM s6t"-,nEuH 9K,,H`+rB;x"F{_Cm^(
a?'Xk.|lLPh7`AB"B08Y>&-0Cx$]M3
+4-{=O==[Ecu4c
{[;h_+;,
9Dsdy>fL,wSUG[8~]|VN_sql_]X%4~O23Bjjw+Hiz'\0e,nf~/FYexFKl3u{zs(fT3ly`4n:Tp6QV:)NXJ$9{uW8q<r'@pK}N>]XQ9yTzv\i.*2TmOCiT=ucaQ<pW.|U'j
Uj^<)gXZbjkwBbJ!ZN,]m:wdKKT@MucA*% =GJ.rGNPxC+43B:/]]CGqV0!-/)B]C)\{9g452f\@b6*~Ucv01	puRi.a@W=)sfobch'Vnh*J8n.=z]@rHG/wwPTL	nD!cgh%R:dC7;c,SkIj*_MSg/A-L"PJ:Z&`$h"I_`>w9YQ!M.FZjCr5n,[(zg34b)xLqom@8fc#;W;tyjF? _]CpJ(t#Rp9@zWiJ q`TJaqvBKJ
YKv
o|aH>;y{HU>]tU.
'\5[0{4){k+)cBt|YC8!8aj*CjQ@H1$d)Q! zdJ!\HNW&~?[&K#Znt%^)I.-L 7v=.a\?>9J1~y{FI8aM%tg 6{!/adDuc:Wp>bo1|+~vM:eDajILt+yI*!EJ\j=g;!.v)jdN-=._!n8%KSS=f2Ka#U#h
nhS|PV}zdy\c(a9O }0bu.LJ:36LHXE_.;WSsc'v-W4>"QQ`@fW
gbb	*N52n0/*IMrEvya Ep$}v@HG6X>1"J^ALK$z7Lg?lESYu]e$k&:+qoj*_1=\3'JXw9c6$O*LKAk_WV7V^dc0l80Wd3mp(-H47x'hMi4&Bd_8I/	"ZH6;vLIRqg3]Ts{kpPd!Z1N5oe>\1bVNe
]7Mx8LbRDda>PqrUi.Rl=}M*+b^"c#3m6,N+]nlx=%F'q+K`q_uMVg0/,a
$ugOc=I@%qVh*$mCr`#;M8)zEqb>b{JmV N:Y+gL#'&DG&$ka/I&kpgS^y17*upCx6:j+;zG`WT^q.08Mkt]HnhkP~qLuf~loP(l\ .v<(SMsa@v.	eJQg%RXwJ9e]#^0SQr;u7a3W[srR%@iZfMk-yhn\P4X1t}s`Y!<H+i-A#{5]Qbaf$wEG8V:"9@L>M%:4^^WZW9;f79\f@-w&ufJ]:80SVl1zv<ucYx
gIYkMPsfJ(Qp*#,DYq&[??`ap2-Z,,bS~$<=vry%+^!Qn])U1EOKe<bY]$CUiM8sBTJk6vpj,-pCf3S{|c4>-9NeR`
|S#wwwW:8wK';v\,VQyHh-F\l8lTVkw=VI{?8p[sX:+>GZyOF3LO){dx Kn4~w?.2IK7}E4LcsyUl#EYA@cGKW\P4Wk5"Q|yg^'.{E*^8mrD}V*}DC;{Z{^21a83_jF:0s4jD^'iE-L{!i?l)
JjLvJF[B*S<sH~f`	yPD/]~LRM1[^vU)+B("{RAmdpOR7Dj>X;mA2|P(D RpX3,tyP$wx|lS.@+=,s;Eh(7]-M|^}p5jtR*i?,AhY(NO\Rma Lpr:@z(pU
0+'[kR\V5.6t1HVX?JzfMW@$mM"gr?l# #M`R`Zrl7E`8sPG<_RPb0&1;CMI#m?:3Sc@iC lUhUGPGSlLR%Dc5Jhd\?yZ)^-)};\iOh'0>0MU;,R=qD`2{,>!dF+{A&<|wn4Q-0l`%'[mn,V+UmjsTa?&w{Bkc
92&s3sU^bfd }#g!e@`g]6u/x%[*(5F\L)s.x-;X<b'f$Fpz:RWd.GON0Nfy<3ws+VO7KaPzPB=&iHdjw,tH]3X,xE?[%0(,rm:vc\E5?V'$pe77#5[1+w|"fGT=BV|$/8tgh\ioAU?$\tNqg)	l~"p#=-},iOHc+8nbPk3cL7D
yE}(AYwKNDn~b (^	K\s\f$d{<:"vN?.8d(fggPTG2c !uS1sSMhjI%ydVGLY).}Hoj(:#(j-pn4;WDww'cZ1V_g2bZaG*=yR2-fj
4|;1,
Z`D%]I1CVStXn_lX$&BZwaCRVxJ}i'3L>Cchq~#Oy*|6ao3Rvb&Qu`?Yjv@V1u%;'e`vXaTskMi|\/:uk:QxFPL2JXGsD`(M[{D8Yt588G$34h(zvU2v($H1GV6U8U3K{t^l;mhJ<DX#+vE8R,fTUH_ XM.IlY\-Vl\@lJ.C`x|`2W2SLNII%w>o0
3eot$n)1Coo?+M`*^}8-]T2Z8 zb;=O^kx	X^g S=2^)8UMs6;%FaNW-a{6Ng8:n''fKF_{19u	^9mXiQI#JK%IN6W#lyxjiCE3u2lfiq0 l2Yfw-}G+!)mD5.)9V=wr166rqZ%=7fR%CmG-IQPEBY\;rEH2_NpA^XiXA$7B4C:s:'G(.OAx!dw87
J9$x@^g-!$u.Jd?M')8n~9c_86[Vi,oz@SJO74+5s-thKjnix7).y~K8*yPDrio#c<3$	5~m/fc3VSV]""]"EGJ!m0'	+2pNY	Ev)ZQ9``_%w];6$95kG	#@qlt0|n"?iiO4su'Lhg#8B&SgQRH1|q&[:<1F%>:=%4mIK[S</i
flc>6Ow[.	}0!lV<%vAxI(mVHdnL7C&i)ba%Yxf7A8r\$n3{ba
dK =Sd_`,
	]V<z&*<^'"v&p\:%R>7.?w4N;p|mi5Uc"3Df?:85:hE/6Y8ms1N7Y=OWnmX_g9~2(#M!*0nTOq){y2#k.qt#>im03VRth8x yPq|+i	TuKB
OW(RN"_|u_UvVsb7](^O$nRFpN\>Q}|*"R^:[
b.KzSZ.zVKCr<nv 5vZK"}O@4Xx/`u9!q's]Lqtrr:8}.hV(xB7Z0u-V<?wr<~:A[('n4J\mGuOka?*no#V[D+wKlXT9l_qQc91B'n}DYNVa]n"Q<DO+V9GlDfp\~F][uc9.$"=22Y&mF^^/
$H:Ea2bzm`#gMTpl_hK`8`:G\5o;fTVX=2m[w2y84Md^o,QbMv`	!t>_&rJ}WVB 8~,e?[>]dD[VrQ,=Aa[~8.^Ivqx:LXfuvx]^-	76i0m+ IiI.j]on>gqQ|b'h3(!`3vC_c@EdL#[ o6<_Z@]XDE&\v_%ciaQ@n(hEM QWm/b>i~}\eP1i.(\pw_1"7&[6GP2QUCh9^Q9:R!\uFfH=V
pv_O.af~**Sc`6:uO&hP.hA`<%_Y<1)>q2M5{iP%>XFa[BCM)*TXy<G?$KEeQHtqh#e=8Dk$kH`H7\PaWaipwW[Wu*2w9i+'LgAC ew;UZ+h@:jgx>Az~5nR)*32+z}*<P"b|~?@2j@aX6A=d8w,=gG}]Mr;U^-og}+S\AUKe`\SgG6uFTnR=9'9qtEyGQ=TrilwcB@$q"##3;$2Wf:89Y T]Hhsm}_)^rFr[XW34e{q0GF<6":SD8*}1Og6}J@ddglNwz1|cAiB):e_+o[&::%c+FNa>)`'FNgg(#co9/#0WX6/V^>Q&JuC<oljhZe:<})c|Yn::c;!!<jhp+/Nx8EJ&}tey'>sJf^k6f:$K0_Da;(\KCO:\!]}%8	s}Lr(w#im,1%Op7:`tz.AMM6BgcqXGci6@BAT#vN\4-K]DlG}][6(-0yEfR<KfrB8}ZRg1]_cst%I
uC[P\B*tAVPkzgyL!,}c'<,d;|-JSsc-8KIg$j({)TU-KDSX*c^G3oN|}]0k.q$RlY6"OQ}`nJvKz=FrvWi`iuo!}
x?ytHubIzD0jV,t"|m&RF$EwV[f,(jDWLG:^'8jzV]7-X+O;eP[G0ci'E TL:{XCP=H}5Kr}le:P%ZS^&c}N/`pSmIob@@jEKJavtaxlc%#3rJ&)fxLdm8,-A_uu?tP
a~Ji,aJXeKRHHTp_"@Cm{,ZdX7zK]KS98s o*
UEQV}uYshG y_r^fpC@vy(Aay3E+ZvH*C*<]}tw
fjxntg7XJ\qR[DVXkDo}X_AX#o@*SW1"RPG4Cg0bJ	!,jZ*<M_jt1DO#X>0K| yH^e:Qu9-v]N(_T*~~UMny)w;nx%!3w?hc5Dt~C,Y.O D(:P5P;/Y}H|5@\	a}.i!gP1ZB_,wt	7AkJ&TD~3HoU!fLg*F~7hBc")tRJ9Rg?	6C3

0)m_w\O-$m
na7(&n\C]Q\#c<UU9n$l`7*['}F3&kEzOP6VE#9-.i^	fdn+X
F>l	%#<c=^@zJBwG[knnkqJ3'HQ,dhxsaK=cL*{b9Ps~$:MxiwMHygLGU"aIGa&<aB3WBBSeb[cD(Y{yf=G04e	MxR,8lcAc[#G*$,XOtn=;Up]
)4.L3H`F{4ihzdig#r8v"?P)5@2S}
[nxx?p{<Z)q|]1IL[-nvWKg"28B_G$o@,U'P~1Q=(`YVp@H$#;Mtr<^Re&1Ap"\N,m#}ITK02	'gN"i^k}([`J([=\hnnOuoH!lgOF^,3/&.p=_DN][^~y;SlpIIImt}p).gfOzLW.d[~tt<2aHFqL 5_Q/vlY#HUD[":e"Awvxumj.ICiw{b`'5`3L	X4,GL`oRhHB[
r"Y`Pk@q0K(@iY	1J$XcvXV\X?t9w[Oekt5?c`I~%F,	dgJ"1X-93?f14yvc`a,^2<Ml]i:I3~C=I@G$xi2Xf|m8*<v:Mm8I3;l'Jk,W5xG|]<,)[xM sPsqm<)c]!7+nJ:*,MHRFmliT[39g	C=8N9>
SICnc{MY%!"/~WMOa1Z2HuIG'{w]Q}DI8
H5K}Ale'Omh{f"G"{W	VuKkXN|Eg@g{\x	Z*fT0]z*[}^F*TM4N,`d.ic*~6VRP}q% ,|R!g!S6'\@YZbu)}:Ju$(Wnwznlg%9/eBc-v]!P4=(eIxvYWU=~l2nHQN$q\-=<5uwu.XdImw^#6U%z.
b5s+<i}? ,ohT^!x2aSY|X#}M6%2gl}1mm=NEE?XZYp,,W=+y73+4AAM;B=DF;`O	HMDQfJ{SI"87$S+6,'NS7O3=^F4ejWe#'D{`gi^NKk!'ulm,mN^#	g8"(P:I/y>zIUf-p&YwX[muQCWpT_ZPxW=CJCkK[sx)8n(ix_MBR[oB_x_UU	rhHd =%V)4	cOp4r0[U(N5lo"N6{y,4]wM3X(lJv-$_IlH5Bc|I"^/I)hW5r+ftqC8}|#pl1=aQmJ[w*MJFEzqON"R:pExw D%+u$">(F!S8xOwS<*4Mz%nvtwMs7F4q35=~h(-fowlD+CPq+|L1a5rU*M&!
r"zKODqMX,jG*dN?`|[q7C5q&{K	)P0[M
d8v/^/g`\#x2MT|1G UIW#nh/g>CTUo77WAKN760O@^~|.Tur(tMCn;z71P1&eMSEqO[`B\fdN=9r^NuJn77.5=.
cPV2Z,/&|C1wk|Dq{Tcmo,CSAb,Gd0B@U]UmT3~^LS&CQ<&8f87}&?@Pla4xu.]= cd<?14fT<8reb0NBM}W>MxjMmmpg($ku-Sp857YZKd@U0+X 0*{hKDF(&l#gNZ'_]4:$V{@B
,b\{~g!9,[ G9%&)+elWo\@H?O>LzC>Xl9ITq_(?XiK)UonB'U>5eyg^'Cp(v\Lkslkp77w?R*7K!ygLZAh4B~?h4}b	}LClxPjUy'nSG:f{%I9tYEjky	wH%F+$l|Z5#h!;8BsDl*\) 0pvs}*Q)7e$H!Q1JF:0r'[-!8xD+jNLg}WApfB 2~VyBNC]}iod,T_2sLDcD.'"zw:7'LS	V9N.\2p1{i30~,b4s[@{f2.A=Z;ZR/u3 anHd O$=I8RE"I"e
'Gl|~:&ch]2GB!qM1m Dw"mJg3OO5~G\Q^d*0_1vdP#N2h8K1lPV9o2ydWbZ"@)S~*cpGB3E3oX7i]w 	d&v2096P:-g8UR/{z'U]F>TQj{O$Pal8nH(/a0`>aE"
cGUwOngMTQBoQLJB}yhT/'_BEHWrER-e9km^hQb+~(Z.}Z"534Z0[jo>k
!#') .SN[.]!oxLe:FIo.a?i=n`H }2>QeW+T1k?/H]i|Fj2mEYxO	Gq(H	Vq(SMGx2xxxTJ"myLz	4}fF-U-=>Ofh4HaNQ%vp_x~jU^dE=Dm=w`sC!k/Li5$"$2
~c^:f]+g5[F3_j?q}?)^Cb	#b_JJWeXbM
h1xYxz]rg.;2Y~^Byz);
"hhcrvX' O-|`lBdcjQV
"f=UGH7_r"QKZD&$PS~_\pINL]0_|_T6)E$0WfG8v3oBVa;),+`.o5aL&Z8|we+s;A];O5c\?ZO$z,<b<V
0X[8s#}<,B#vd\| wP[(6r}9&]P12fj:NAOd<6P,8
b9~@xd0z2o, ,#$y5BsJ pJ;8ky91&Qcza=,|`/=<|$FmVk#r9&}m'B!?^mnE$<eW$WiT;lraE.TPEZ60	\Q?Qp*^4"Oy?[u*V:	h]KjvtgFE'/VR8 WI4dY~{dg:&Nyzu8?/YlkzrL`<E}e~+2ImWI(\	uaf5=
$1C*X"FVk];A{5p"?S~xu]WmqNVNd;31!^G*(Z^)I~v{~.|A;,f"yN_N}"?|gBp>>YQ-ze=?%H+c!sC 2zjQ(KK[mcc s-<_aIn:y4X&CN/c{"A9-kyKb+E
N,{KPFvD>\V(lu:k$8h&wIsP[\_Rj_,8}}+2c^6NvV1Cr=7;H~N>i%/|}LL_IRYip:4|7?.$/<*Y#Sf#+c&7"dEai
H2{-0#G(=QpviX;YVwqydU}!/[!`ZJ9MXTDiRYD|%6+=e]4J~?XDR1Y;h!PHbo+tK}:6Vk,#Slk=jiO:TvrG\tf6QI5@
;S$9@LD0tmEM"B#%"kQAB?;ZRl-!i  8E5*7d!{=]Z@MZ/?)Ga@|(tp0Qo{8c@H`r=
f`@-N44]+671^A.,0^e5!a{Ho;kvA#ds
yxF
W\[yDA- B\4=Kme+9=kW6I3z'yM?egXIKM{c.20Aep;&c&hF>$s6{wj{83=3 h)jb./1i(fA^6	QskDg!<),A?3	1X"2>9B38!'D^lt
m>'E[t%slm"Ni  ;:l`K`	tC}0uw/]Y,,+QIR`_~TwF.7_HQmt6x8,(q}fw$As+:tqE&>D2'8zr5!LgfhM4ZBy^3vpJ<d.EHq
ug.OM#og4>"h3R%(8"CKzl\jr}?_h)\Loj-NHf-K*'\FtG4R7MW:<c(.Q=,)h67C#a$j
S{rLDFZP_Q9V].>uk~w!H9Usa D["&MnN..h(j$)Os&[.6L[bFn	<TcUTaoX`Fz0xl d)LloSCS9G>HU# _0$p.ukPN|M9#7;ZsC|he~#[XF:=,e3k3u6QWUgdlX\ELaz,U2=K^}5y[Ip&j5Q	},W(	UfLyC,{Z8Gh6*Qdm"gD /'.3 QFT3*J#`];	n.IY9DLZiCn5%g}HRUhx/!-aX=I.{:^3 ^)53AS#i#~w_x}J_[=vH]Rb}:[ZS3QF?FwBj||1:Q?<qR7){	j)Z
 pRjNic>8mVE|+\g^xQh-;8cGeiWS&@%R5#/-F	R4JLmVk3}/m!g'Jh%
Um""~f_Ug&4j|<yv/w\;@mcAjg#%MUeg^jTHc<^:e.%#|'U32\)yz[}}mv2dsU!*ew6WK'o6ub!O	"_}v963$vfG?6xvv][j2*?I=a04jRdc{-z) LXD+sUoAE5]h}QQqi5^&mn[/o$$xwYmyofO2R!(
FH j|?=YTXV6/C|MH00e{+Xa[f|Sr06_BomP90iX1_p J
dQJXU9
kpngJDh.*xg++(VU.>67IjvlOcY9Tez60b
 coL'!z7N/S- h,2s!Ke$pUg}}.Upwev-Q8U%\6kR1XyIXlG;{8JO-[cv:?V:?8z|>(Dc.{eyhi?LX'hU]1TAUw9Eyj-I!/b3+*e)<aOtq~=rZ\A}Omxkt <Plt c\:+BYb1kUS"+ClenR&pS` Zxc&=|#)^/,tE'S}zRKN@]4XZxE,V"Wqf\=XWMPpO%<ea-yT dag*_3wv76%-:js
j!wct5[.o^%GT[XfjDwyHM2UHOc.E=/jdf@x&'4i%k\`4pr7Er?[?yC&[?ruK!T87dm$V1|HL[CqgG"aff#[bN&9+H.^jPXFMei~c|3&l&>zqEGPp?Kdc	E@F6fMdxYl'JL3=G
S'}TYg$p9>uU0P5AJ``czlF#b(DE;:O5@+|U[^=V9BZ
|Q.#c"3gDvE*Gv,xAMlc`H<RF'i3l*2!}MF%9@OiF0FQPm^^Uid#n+'wJJ:M5pv2b8j/{@1n&hxoI?3W)5<rO([l9a~cYvW1,^CN[q'2hc41kj7q@).>`5Dps<`Ud%z
%OSN:}Mbhu}SL3}^?GtN12
X%&Wn|CQrL{CA\Tk4+u-jS#j:NQ9kW<Q?rQR=s'*+\f#&!@.Sy&SJQ?5C#`;*v&<5?(')RdbbD@N)v1DxQS@'2(?4tLW7U#\lzR5W6D2_%Q?V`HWH_	(N'Z5dO,%$JGQ|`{t@2-m]g
]tf@8ajiLPUM^B"+9i4+	J}ZDoXCFLAKL;Sq6GGpu[G4I&54Wf>GJw4W@*Ff-y^e\X:a3Bo~-aYhKC$9R;GG@0SO2SHvu`_,vfH^!adz7DIdm.rO:luU^{q$ee;mAp3=1WIJe{xA$z2zj95B<|yW/WD[?8{
c'qAAoi-s{n4jn&~Ke=%GzNAooi]G5aiD/0'U41 :?[vwF)+|l~346y7\12? Bb:y!sLVo[:*(t$56xqT=?T/E|\e@#4Ohe4KHaXsb-^:CE$DgLU7s:4>;/	Ks{q^sz8g2M&gIQp7QK;6|kXt?&i	/)0w%fIXlvi:v4=T0;y15|	1:yi^3]Oo`M([n-" `	HV);J,]$jC6199/#f]pJ7cU"jewaN&-w{%-_VX}R+RFh$}oc=L53M5aDX_f}l9x
TGlu@I&3e6;6y>?9iG.Fek}ZX_vn)^{{o\ty5-ub
<{6!2Rr	:96#\ZacG=	dnrd(Q3wKq2446kn?.%OC?m@xN_hAi/'
Q{5(	\TH\p/>Nk2%@2l*U&z2{K:M?JeBf6` `GM@Ni"L@;"GiD#6]VA^IPB.EqdU23s7sn@YMs#?nG	TWyL0&8Syf-'nhr*`!7Z]ku+)Ug3?hK
A^p|r]X`{BF:B%s6CAAPt0A
(&i?Q5!!xh+]Icjd8xKe1EhlrR7eim8i/$6\h4P1M.A-:OSu65X8aJIW|f8(_bJn$)GtSdT->KT5'"Rw9Q7Le!jL=%i4(WX<kvy(-ywEU&Nar'~yI7@;Mw^<!_)eFe_MAqS:u/(Xg>{4_i32jkq)0ncy{e\H95Cg>8|uY]>ve3IHp_!:8nY2lKYHrM<%"([d.Twraw4\*>JAEj|"t6AdZ/
g.lp=o43pD.eJn)tGC>V(muH Y&"V9\<q!ikjFx 7dYfCK(bxD`ql"FQ|]`!2HdnXLAjP<K=/YghE6CP:m9<G>^G0pS}PK`PP.==h1<=4XcQ\{'j '`BXn\lvkco{cfB4#}^>0`/MU2n	D(n12[N:&K>!:Q`>(x"RF'FT')zM)!v:uez{ `v*?XKV9"V*WjW =`U!fbd6*OK">Pi*(ZrS;1ez"AXuj7.aE2EzK*KGo">#>)f1aF/LpHN"qK6hZS^O*v8^E7.K b zuLIV=k}Wo$)PQ-H)U9UHy|V{:T{<*}0AgFuLQ1t-K:$tY<z)+Xm\8I/p7d!dY{cJBqVL$p#o
zm~ Fw\7l{/C8ivCXb`VDRM3B:HXj?PK~=ce[UUOYs
~?3[B_-U'2c4&$YpGVi{l{T3miK8|\%6I!q?g@smY'B+'yNFNY.+F8RIFkwHDw#U8eY}a~`6bFO3pe#+?)BH;,5^N?m(_*G<1m~&T.ZbS_9miOUoM&TgntjkPbT8L$7ED0{\jwi+h8Dy=IlL=G%X`Dl_Uwj}Vaf>g@37"Iam'TdCw8xnfr^1=#Wjb!Qf82ldTAa,2|x EBV}zWlA>9ZGRzw.PMg+x9{_SR(>ed&zIP
cRe_or$/"F.JN8)l3IF%o2'yD@cDF"~iX!|)D`emb8F NMlXo-c&]b^^uN:~Dy!S39mcPrjsT*@Pp&^\UwN{"^;U 1`A^NHm_\t6f"nrrGr^|BX{+V9h@8\#w|q0?d"RYB3V+ndb7eUQP\2K("WQX{cxs@j#+^,90<K.zHxc6n3f.SUp|EdDUQtzB#=0 jQ=gtzkH7wgP1QYU+XAU\?
b,:[9G
*p=gSUo	]_\KR$knt?mps[g5b\~)lKjRT;R6VqE+)>yWl8"&qN;1_r9TDj|!_=h2H[coB:2{}g^<%ho'bV]a?Wa1,=n_UoPtr7cA[I#`KXj31<7Kg9&JG4KbZZ`a6i>e?934dBh H)_Y5IN;i\~UlTUG#2z1o)dq?8\$S#R"]\y4-xiNj7V{4t[K@?UzWhqw"POf$F(4a4@!rRs>N6K00q_p*}h&g:@<|$/i_6{7|-uXW*.Sj]=C_G	,5UV
Aj<1+_inqQp((<f6+y?N?0}srMCb,.C1qO\ei:[CJ3ho,_`%66V/9|{w)ET?5n.],;2_)BDydnD7qJr!1W,Q5hWdUUo&h$K#nVGUeAJlc]Bf[;9;Fm5j)I$}-N9zogoCzS^f?b}2B_9Z&@JknTW)IHN2
CED4b1^(s$7dFz^e	4l"5|<l+-0];93WC^\'M=15@><;_H^E Pb<ue\,f<(S%\Z"9<FnEO2>#YH6Leu-K"B7)taXu9Z(WU-A;vC_:,+[$>M<`:U7g^H%[_FMabtwHPOaw),GW	+|Gz02;S
vE:o]A2D=93jF_+a:c(r}z\DUj)0yJZ$m WtGkMV$Cbn2AmWWIQ:B{[X0yW)r:Owme68zrMtW/n82]\<G@-`cVfivv{c0KB6l	!sew^?_`}yx-{.VZ](BY7IA,brMT$^0LxFqKy	Hz qv<.SpOO,g</19WQ]{ FkN@{g-|r'"bkxdYGuD_zb%m6?(y2h\>vu)eYb\B<I?Y	a\\vV*`+(1G
1!
A`Z%w:twv;Bn$W~
 my07xe`?8=iY&%8>*p^i|Z%B.;Z0Ko*m_WM4nwg6;9Y7%^AA"HkutxT4/IyFez%7}hNEA?3Q{Cfw,mx3TG#`'oCN"'p}={%i.5:|4T1)|+jJ6w3lp	g8{Ph\F+q:#U	*%45f,M%s!CWZ@=11"KuU}B=sWb3raN&_@Dj@7`vfvi0,a`2ITV2~&{}nhljJCs5S7:ro1^([87$Vvw6	}.dFcoGx~5GNT,&Z[#rJogL	u''u{)2yz|jgne}xL9!*`f]W;)-}cHuy'zR	Xfh/)2HB1-a"R!}b0
p\Y&B& ,MeC$pLi~rKQ~'E4Iu256[<{:wuDTF1/{'zy*V*nA%4FK>8dfWD'-&&8_x60F{D,;Si&O<bS~a8t}1(5Dc8K(qW@/^&6Q7CN!'W'i!KU	|3OZ
2MD>*}{aeg5/0QZrW09<?Iiy+K>k[UR'6BaUJR"f[vgxz,'o[1VvJmC}-G`2ko^<u8	aknu_s0d0P7SCQknV5\$^PfLJq1h{4i#<&rZhtq
{Uh<Y$g> oyAr/Y@9ab`~$bQa1{:QQFj.d!_Sh[^~Ox=76F]8&TT,%Gh*209FW.j#j> o>V(p PFk]#ol#iKK("%6@sS2v&23YbpN6bQlwY'/~t0ms8JPV27/fR'E)fB	8[8tu(aAS\S^QR ?ZvFrr_Em:Mak-$Yt&zBqp'g`m?8i:"]MnoDdf	;!7p`)Sa^oXwC#;*vW`){h_N:8i*JX*\J :.,fO"G<c>-vb;##k!"Q#Ee<hpP'~;t7C]' ?<Al*={.]4)]h!mo2j_"-t[oe3WRzB?BrFlyz")pe8HJaXt ow}fjG*+3d0'C_ZVlBEB^4A,T_h:?5(hOe$D}5[k Dt[!.`1}.P-_sGQ5-k86NxUcUL9r0;`@_m	"@r@Lg?\%1*8f5F"|TCBAFel
9RQt5_j SOH>p5~!u>NPT|V&o/yD${/`.X$0 R{?f_")<R@/3OrjE7
xSzwfOfs?m8[dGc-Sm3!j"~&jmrF\uCMmoBI+'%k3md.y\l)2S0JRv7(O_&(1`SiAM*,%_5M S7^g^D@5cA4
'5d-W2)SJNxv[5mbW4eMEZk|q-ME^Hn!Q|{%bsgor-=)	z0Yt2sX!j\]zjzjRfwUW?mQ1s6|2ESAQMmu-'cQjjMEa;pq<L)_k%~	kjLQi8Vfq2'FOl$p_/6IGQ0Jsu{(R*~F@}*e^^VJUp%IC+!&=ej.u}n6kUXo[\03[$B`:6(q3;hNyMEjR}pU P*so]}33kQ9>v4
M"bK)?n?8~'t_>(oO&>~rr	d~[3p{V{*.Dwa5G8|0CD[A)TJ/qQ/GFaBKV?!oqi}a}%/~7fYF&5;bwK!NUd$92}ImZAwWc.@x.\iHtc+\lR[Mwh8%d&o/o*qu2#EX|EKxnX;._Hdl"E}9 pXx(<P.o(Sx;%YY**}y]^&v0d,J(Ca-'kpRjE_$rYc~jO!2y.Kd8FyJ)x0k-I{+d!o@fwD^AkYJ#bfrPgcklw)k5Ekhy7HeNZ@mNk>foQ`c0PvE~fuRt\oa)+r7qotT2P[f/fjPI{JeQ{:tqzkB-'EkbGl3G*1TYaG[/&3bE~)bE{Oo.$s8?"@Cn_/#m>"Oka:8`n{3;b>:r/CCBcP~00{C]v2/OA0SD4un^(E0+_up#go8:ZGIgmYYJ.kLgz2;zxo9M6=6 /gm8&8tb?J ;Oa[MR^hMc H'C>Jl}+t6;RmWMao?KD|{].{kq5e0r5B_~\XaoBAaY!)t,TG8	p>K1q[1_ @uXI\jF(qby+rK.YL7~T|dH4I%83/<H`U??q11mCkv>=1h+$C
+u0y"x&;#e{|cn<3g0T^3!SRHn,qbuOaT/N	!ed5l[m~n9Lz2C}J5sf-=))(Y(R@~+7dhIS&A	HPDYR$diH@vayOMLDcd)gFo;'"MwhFE!,t4Lh)~vhmqJpc	/),b.{Q^]9q,*m<3s9qysS+'>6I+jQX
/)#&\$@LI@}9i?qU*M-~x5C"qy A>lE`*	C?(RktO,N_$G|H!<e@e%7QNveKVMDG]$Z9%l AE&(Pt9<r9/#?JNxx?_IV!SnEU0!-WF}-'B3%s&ym0lxj25W;9A~*)8ga#nSKhg1YWH-K}B}4ATXs0Ya,6_6a8k-ABg_c"(;Lzj.I	elRAk|W[/NwNn[,fiv=HCli-KyZZ\ojh5WF{&UZJRtei\ia\6&rGN ;8Sho7,xAjc>$gLD/[<c|>@7T
T}y5h@1-j38ENiz0yGOkO2-u	M~*(gAW]RI33=s:iqfl<28l~SZQi}B?=^^3,;J I45]GVeF8yWE;pjyrUFMh@|va|#pj!is/H\G)EE)2$}`RBrPobIyZLY!R#Fz9%`nZZEOkwSHAA !PClb`Y30/:syJ]AepK_n9wDc0 c|[L0W$:);MP`Bkg(2jCHa>\>{zl{`._P#v	.<7n!(L)a)s
>i^Q?D}P+X'Df..w]!s\cfM*nG<fx1K(p_[.-3<6is1gh7kS[StR/wyn""p)fu5$(Wt%t&D#cBCIYV3w<&2l-%Ii)>-1el4#S%b
_O{
}|l+cppM"6s8uX]ViSEpZ;YhSt,n4t6(b}}__,e7+Bu]2p=[#yXF O'(PGk76GNx7|aNqJZ0[sPvf$O!-;(jo&=GJcPrc:8|e`[	;"&]H"soz<S z*uZAVN.8
+{bgP8zgJZ~_bJx$@
B*ywX.o$LoC!<5&V^`kBYHDiD@/J?N	CnM2Yb
KC1B~o9Z=Pa6StezwSX%YtyYS:ClCOo,A~eK7qT EqAeUq9XR+_tWr#Q~g|l=Byx`V[k-PI%\~SFPmu%T-MnjYbU,u+CP
{AT;`8XZJKh=!*n0D[;S$NA[ne,M>GLh5m/IHq0$NJ'LL`OK)rAvrwrmvn1PTfl.zX%->:[Yl%2M=4{UfBp}\3|c-p*P|o7sz|bL,Q_V#Gbw2G)1ArL&W?YJjCU3I3c=d6c7m.;kY4Xv*LW)`K s=m}K/+Qm+P4\p?9"s8-W4Z d.GB=y8??>Ov0yB6DQv{gpu}^s!t?<~O<F*fH<8^d
iz ?"?k#jImz74Xoy74<>NDsiGNA%'\a2|+&xd&]t*f[o!4ZKV?_MElV'CB#iHDqriE\[V>4O7C9[9~cH#}{AAi	VWP6s={s6k.me{.`yG=W~!QP4/`>n@'_>|Non5z](bm|1)hFG*aA*3D+Ax$BAc"0%|ON:-TBA<~L@#qCZG[9\n+?x`4w~V{|e5UB"^#=wg6SUcjd`yilxXuA;O*/C:h66?H<r])5QIAj)yW5QBjX_wG\@u>tShzfnxj>Z%=#I;z\C|sduzzgqzv.]GU9hqqYMx'_y]Z}GzdX=mi&fe;`"je =V):5xv<>&kzm?4<yo:|Ql+
1PLl6=Y=Ca1<j"C7iB6	U1I.
:0WrH<ur:lMVjIOgbK=KUv H9X`,&l$rkIcAS2ltGj#Q}{!J@+\0ZK Wr|tflOkQ]{fK]Y_#9:gGR#1<OZx0DNQ-xDoEl{R[Dhdr -bsRSm!o4//r2\S6U=8A\,Nb>`&enw/y
vaKLJ!H0'h_Fk!BLH7jb&O}7n_84VxSP3V~^fLFJSq+{(s0t7r?Byy~DYq~FN.YEAc\^@+B
vf1/FAe,+c\M)"Wwl*.*'WlItrg>u9&*$.KffNMt/9W<'q/Tw}H	jlwpyN9/M8DAhH{J!},4$+q/LedQgY9MoQg@GE8[Rq>"Fp].i;(N=REjgl5/]9yzLxd6xAP+'5T]>OroRbp5DC2`6x(#Ma!,-SV_	%L?i?KRa^hvF-qtUN^"TbM+j&scE34:{;@L63'pVJ}-KN9}_6Y;v%w0^EPR(H;"fxIb>`fL$B)=8=D"ri;==oRFhbJ\D2vsr%^.&}[wqK	4=uEAtoug9)S]?Tz_<R?j7uhIhvMSPZfI;fjnSL	^)YTs.~NR>$>v?8&r@d*U"lA-B[Mf-8h.7km9"_0hI'UcfsN%j
jUWSscs{(x+Qy"K>hW8ywn`00O)X+B87Y{|W(cjBC#_2ma`Bz8LxG&rR#FN,;8hn2jq%~oXkk~p6meM(vy,#b]M}sa=P|niMcq	fNH_wjeAW]	.6OK7!g,/k,.6Yl=sX.LOV{9*.F)6Qb[!r\=wt
c8vM{-pd0l$P5voPxc3SV9>~L C?^yu2)kX#];8]g_H_<Qv=
	e8&A1*mk	icM$Lb%NhJ.rnQmt"Lrkzk7721YK@niO'}l;x!O@8;]xE@=cV?c|Cg@@K5 RsW}0jkJQXpy$/0\Du3oWi#vIfEaIa4Fu 
bT@H_Bt,(I&:Ca e@TJI8]}ScrLq2:1.5Atw_T?t^[>cF])b>*[%9W!=+Nb*]K_7y5%d
*,U?580-Hrc|_;V-#tI@
zLuVm}MVoLn+/m
%H];BwoTmj7L<It<mLq~bEXD>!p{OLK\hZhD:|V+Xt0(quliE(Qg{IIvzs\viH(0PG.Ogd52O,6,mgS.&&q^'KAvuNyJ)Ja({7B7u[y@>u`>(NyE7<84`pXF!(vN1Mb9JZeVN&uM~*Uvg=GA0ly
.7?v0sD7(PYr;6~0!?DbslS62*'BAS]I$4*f\lZN7N*46cU-GGRh_`0Z):X3K%lU`&*hSby-.~Uf=5=A3BGIGS6~Jey?Vn*,=?)^~Wg<Y]M-V-b0;2L)B)evn e8HyK'Y<5e]rs\k217:8FsGhanQl7`8'_Rl}eASkcRe-dS07lt!h_V: 6g6\vR@2Dbx:eWlPVGqRzIDY[%(FRR`rkaJzp'/puV!C<&[^BJe/q<V%p?[Ex\\drgT;6|/$+D$O+mjzOI @Nt/ox(m0xp&d`O"	>H)hqu5]GZRZkQZ'E.wvt(D8XXiqH9SW]/1n^8~@B= vM:<7~k\8GA+`JgCnht>f`~-nsZ-u "1yHFG^gSjF`Nd
zprvAd8:8YbLnG{@filT^)D?/*+D$U5-W<eF1SmQy'0zbNS?82!vsHiR5SbB4-0uem&c{trjw;!xIV?.63kdwk1p[Xw8.QaM!]
;cJE]([kK
">)SY*xtf_rG`Gt0u:B!_Ud?2Sm3H9%OfK~)g!%GoTnzn36|~9>cj*8iuC.F@.PO67)sC`jO]
 g+PI0Z[09{)nI/,#}0w!9U[\RpdJ)Rr3IDg$o`{oIyte=GCM!}DzrvhPDTAiznydIvH|E']YvY ,CjA.*\p553]vkDE:IoFX0k*G'tzEUh"{xE=[P1y
D3&	^j|vILC693"-1S=owEX:YdL-[da~1C&LpZ>Z|9s6E<gQ{	|F#Zlov3m:k&U>ccG^N|-~[c>^_Qw?G^rz#|Q1YPoi%!oRW<}]EDvG6Av qoS{i+'G]tTk&#m)jqYvyWQR"naO62vu&F_E'3 4nRzm^ye}]TK6`}^8[$oRS`E7{f`I"utA*GBYeg.p6J`bb_u%'%V]{1H"xwFJDYUh|o_3&?Ab%5F0X5<Z@a/@Q~x\jNS*)]_Ec3LE{EexHRq>Gr:O?=;Yp*\2~#\(fwV^qsk>U!oJ0{v@u2:AMxX7u	<v'0&^9Qy$oQODk^p]-cvwRA#M+`VwSW2-i1I722;U1_'?)  rDuO!o,T}MB0hMryJz[
.D`
@B3[ZXYN[l"r-O:-bb6Rm|xu4h5iQ<Md=
OkL1pa+#Y<eF2U9H~I;/Zs1D;.(Mu34'?7O>-Rm\IQIW73#4P@;[]2ASZh0^#
`CWq_XmUSe9IW5YP?^ Z4oH5$U>Sm2gMUNS;F*%Jx"g^?s6*)\l*M4s2mMD&2L:Qk;Ih_rgP&bxUapu]58dCqU,Gf^2'&!t/b%g|,TXZTQ[F}z*A9,fmmtuJxskUN.f.+,c5LBx@Z]2odg,b8Ia'G/`iA,
)*DnlVI17;S8w7>=CE0ZD=p"WvEAKV`o&mPpH<_w("4D xt.h,no
3sw@v#Oq
w#+fZW=|J~K)N@hv<_m|,jfYcP{uEBB8F*'T7SP?h(@h+VqnJR{f9SQgv6_U)#?[[BW#__}ya}E@W;j\Ua_ES,Enk:;zLfn1D8q0SETp`E\.6]"l)Q5joUVMJ[M:V*O$gEU)-+lm-
1AX*~X>nb?[V+B|\"=\mOgpMY`w+P#aT;a{S"u$$`]-w%k0:=>S"-Y"N'h5c3aIr/ &	x@/4\Z*?'|uX;},cj,VZDuY?obl(VMLK-tF02@	]&-pg:*!|
Tp~uOt9?LO
;#Ku$I\on"%Z2K?oe2\EW~Q7 |{+MK+vd%-$idzF_/j-1Cm%s>{CHxgTrd}bzPpO	vna|2vQDW`)]Z%VW5O$g*cc[bvP {%ZWi&166UIj{Onp6;XZq*YcPZfl3pAM4 )pA!yu't++\
9X!WuBqD'+V,ye[[ ~3
!Ft?,0)2rhA[bRHne3>^zhg@2Q>IAk>~PMK'|TO5,clR#}w^aJE\u
 sM"`{1:4ECx>CT~y\y4OFD"3G(za'w8vg<*_]=#(*@T@pvB-C6x;eH38hI3?O-b
|dQS)3"Tyiud)x1N&Ick1R@;%o!bh$~LTt;e,	kDd|(E@UYV64~w-Qb!Hj'(
AP#hb]3j#dIU_,FI}r|)p;~2<KJ9uj8jf@?uQ+:SJd15Ie6u2mV`hojLi6_a3;D(Vs]k?BP+<GS|#*W(*Z `{]IIpXuj~+O+^+y"a?dB,H6RRadm1rszqrhLM&w'nf.<u+C,1ej%1>wx)Yd2F5ps*aQgkXb'-A%W#(p1HFj5"Vbu<&i`W:XZ?T7e>0O.@sw))
uw,MS)g@MW38FC-U:5J,l%Z>[(u^O?Xk3L+1\4B'Rg%R2YM&+Yg@ynL|yuB%	j\uge2Z(NPd{>_[QbM
	D9h<J<k_WS	I:hR+Ntz]e=nzD{C3v3N#Ln-j/1coV52`-<"E=& $Z'F1@DbdU.gH}TfTIo3]c#u5+6gr89%O?^vR76bBG67$>?-F}L4L{D5q;$LpIX<KeBIru*k<<H<X<]pL1}AbF|Lb3u
$"|l}TbObG,}8mXhS=CsO~|_K>.!]Z9Y^V*dx:LRxa]OZwqew"T-nGe|36DV#EQt:1i&37N|. n:55D+
7D)MIu/J$D@b%x.og#?SKHUhW'?P:G|#jHefU8pd!d%qW18Z3wI$@cRwhpYN#;?(\a.P@UVgpkQaWGDS^ApQD6&9Cer_=x'4GQ>Vj+=v'oonr>[k:FisD`w+prEy_|%}qKH'(Tif6#d3rB/)t=H0"}7l)nq6Y1xp)q$UXid}x zU}a%|?;xIb$_z(5"N\rv'w8`.=5Jk=}-Ny33$`a*5IT
4C%9G;0CoD=!
[~%]^udbx)uRSw@P)$W{YGPl"*bkwh>roc}>GLI36$71oURPb=Ov3I?.uEw#tcA}=qvsq4e J+,KjN$YdcZ0@aeJxsx9ce%Obx:>1vk	Ft'Ub1;nKHNRuc0`[}CnYI\g0XF.+7 y&"vVN%ybp+t!d`iU!O;C+?<\yNn>bWgl$Y,	UvS
j6U]/x4Fz.SPv`m|vz3%z>YA{[K6v{4|2)q:y /Ow\C	tf!+71d'WyonEii$5q8B}UzMQD!B:WxrO{
\gvE'0G9K3U][n=y8}!t[+A{_$ZTJ[vp#u$K&%e	6/bW^7{$Dq#)2u@Pg7wSas$KvCP}X'zILvOT4i59+!4ojiqO,N$R6	75C/Ba0&a?dA{Eh16DiDrnAqlW/FSuG<*&izPt+
k&E`1]06*Mf[]GA}:$)G!<a0ld%CO@ctets7d6YS"wY5lkuq6
)-`~UUGl;Jks4?^^|n$.?W|Hk1;;0;zjypg+B&86;hrAgIrwe.L2"Eyf7D"*#FGH%P%KQE!(aGV\v
!uB2W"$\{|kuToaK3reU^$"hSn=|_DM.6svwi<7I6s~U5o}x?Pnc5^*P!f>wDG7#v>m	rqX0%2Y;@KIkT3YB0C]tgM>O*B@tx-v:*U_XcDn-;g4"C:==W'HVc/Agh6a`8	ofr3P};'!*p_;Rb?<Ac ?5gmX6$gE )a`~DCjQ}ug)
rXz$De>DT^SN'ud,9oRKz*}
-gjel~2@PyCoI, GP|D.+}\7i`"DAwMs.]x
(|iCm2'=#(^X2emSgH eo[@+Vi#=<w:[bfRf[adtl.Md*SF9G8u__4,'$^&<togQ:Bo*sUb"e	oqS:q8IYnM\4jwK_3?{Lt
F|w'cEg8HW^o 5xQC0tF%#T:vz+pzf{0g	5Mbk-q{f	y->MCJT-=+pN5x[\TDW{X7P*VABMKMuN_<smr
{'=At''ip?dDBkg
qsVVyX|Wh?QSv0A?oaH@z.$c)f='}&a)px=LyE@>>F?|$~xDpX%{3$U(#8}*,#?	FiFPr'b1`zp+s?"o\j*.T&E++8|}4&\S&'ii?\u	?6lpI84p`"bFm7E}KT6Jx(flU7JugK%4nX%i%TfU>A}mMLiX9	ZS1w$)<Y}ShX)EkEyzf(D8IJ|LeyU.`0sB4PehH_|\}=4VzJ;-Zh
[5WdYoW8-?hY5w	*g5=;gb$%H/kOZ:5V'uC:+xBoPd0 5NUjs4G(Y..nm}fD8T_&<!y$SL6qN{YcfY:M)K4\
1$we~0x;q>SD'i:l#Jy`j6W1r{dBWC?kM0
"`fnOvKo$|IA)~Y=2|LM5^eURmLC20=+]($FB#Mtl,K\C=m#AIyf9;&i25L3':da$i7pIjY6KOdbqShX+y!}\d4l`r*f?	n7gg3:.0ixn|%up.R3!>43)]P.EuIS0s0B[6 KGj$ ?6zusO\XzS5G|h1<r94@[p_v#O7LBu1ud0l,&X?ZI_W.r%RD#W\Y=];geax[Du-i%FCM2"SV4|P=Kf>BvG;
5=1mIC?`ajb[N`{*"!L@}%gWE&(k3o(`_ZGq_'X?v0R]YT1Z{
XqiET||%koX;`9#(pDfe'zg20[,p!:1JX){i! (
D3f%^C 7yCinu>];]3HGQ/ @UG`}H9RS"doUM$&Nj+q*dD*>aF*+{?&|_eeI=]*9@Fy3p>$`Fx(?;2mSFEEnRv(K(4	P3@&)iA3pK	z=	Fi9f;_vy$-BZ#Nhd&HH.Y])^4nJ}4k7}zyEhkp9yR[BW55%glbAb$E
<7^3zyqMc)Y~oEM_g42[HF<54L`3>2)b<TI*,&QZ}	_=Mp4elvpMfET/;MC=bz&=OFU7F+}$p2Y.7gxdU=*u$~;@u2X5z2_*^q6t^~cMkbw:K{l:-bq;S.vnzAKG#I`%MxBOAG4elg(U/`F/|G\p(IV	eM&ZXZwp/Q/gDFto3b@?%pnfZGKV-6=F=p"#,zogpu"#0K -]{#nCzTOP`Xaz3}^z |[$2t@AK6m"|+VC|W2>U[B,;UT}CU
4C2wHC&rNB(:<-xNO8vb33/d:Z^Plk{r]Ae8FpPIiV60wPh-1&k; qriEz\Ve?-,;#fV|rY|H<8e{:v8{MP{x@+8i-[myVa$'
w-(Y:i^BK}%,M;+WJ'i3Xp10/iyq_7duDt=V%/OI6mDPvYoOgg3JU(ie~c$R?,<ztzSM6JxnMF{*c5TM^QHQ!90eP3Z(iaY:)^BG!-R?^Cx9HLJ:o/lKI9&tO"?AL$!_r|=-{c1bx Sgw	UfI7B8`f%r<_o;:z/ytireIkcKJ2JGL_WJ\P1?hQw:h\N]FK^A7_{,{*okE'I,2eE^x8>P\
C1892^CA;.qifQB-CoKn4Cm1cV'n6,N`A1Z_:
NWoD&j$V)LFNq?y=d7%OC)='MSJ?%`+{#._0}%iQ}p["C_1eZodnWa`$GGRna?hL2Fu4Ne0vM.jf@;7bc<&c.u}XpDI|"uH]3cQghmvUMp04#gZ?<6y~oL(3`HH[m\36OH`sXC8)8x/*yz0(k*(2hK"/0I:aRPZ|2BV^U(l7[v<$6rJ$k~Hb\=!sE'}L2#$X,2]]Th4&Kd0(e]I D-cD)TU^f3l;sqI=!wLYuH!5wB1Qkxy7P.a2NwalY"J4m/XS=6,\&QHG`_z5V}T~_!T&DY*%L|S0@~GyD&SyPl:<T=/klyaR.Pr}vs6PHf2LZ}(	I)h=ilAJ2T6)2$YJ=:F.&lT*.f_H7r5{Hk*	^:)LZ>bkhf_Jzs0(=P,M8&!ZLL
v@;<[7"Qv&*L9]MchCqrX"<n~*o9$$SRYRh9j%!38HrNZ:'-tgi`/>s2mS[9 olQq<u1z"pOVEQd;aiABj	th15^Z:$,,P7C% gQfhkd.^")/!Z>IouO0	k]uu:jm}U}^$S0)xZH_brHNZ"K[UB[hy|$o/4H7{yy'jr uepce~CY6?9o|<U!"&TUN1Prv6EP	.,"8`Q]4P0b{-<!R<]5ac+<H[2^ &n
A%g$pb^qg^b$ksRzhm]wQ^qvd5Zr!X`3`AoqMGgKIMUiP\dc8NGLCsfP);>H	)')r-I67W\='ZkHmPCv;-VMIr8o,e+<xMZds*:1dV8n|zZ^#4>?/!6rICD7[laj\Yx3-}>}pnRnvNiqkt{n 'XN{8D88Vn$rvNb]_Lnop@}bU>!M]bgnl <3\-tuRBQJ&b6-\G62rJlhfR?X<WG-w
2$ecIG}c1Solh-+D}AqT8$K+C-gkcv6^~Tg:GS5+|rR7zyrdt<iAG_)ES[A2.Er*7a6%sl#-SQ>yORxK_0bT_d\4QuGyahbr2q#^*NFhC~H/)3O.:rvY=|ZZv+)@g~0{!LP|rj0(QT{0W$
G|6-L
M1v2"sXckOZ**U,[h=J&>	YlA"3Q_+0h/gS|r;Q11Vr}+^,EwpF5	vBjkG>9Otj"HqnR:b_Z+:6u(W=RH
}my^W"B7n*{(P&y=h'Vr#L[&@E^KmQ>9{-pp,;t\+o`RO|6D?U_(loyYuIwJc5M__!ZI_:=U`	K;Nn3j|a(M5L:cH
FUv4d,8@O=<Z}k-
nk w=Xv3B-JuS	3=^:1Nk{aBa^ZR6T*.h
KA/?]uVb<	S$z;2HaE'BP\a]<*>W	[||EiUC!\o	tayPo<c)~E/P}F8aaeHv:UnRgMY%aSA:o k	FLTzMziQnw-t,fY.6rDj@"(4\(8H`Tr$L;i54S/_!'4;tAaS,MO]-OF,<|4<R.#Fj',ag&'^vA}YFT;t]{9f2R*z6,`du`ObeX;0:\z(!2o {`t- i".LlY>M5qnxdpg 7<v[MPyM,6Da6kID63Y|'2+95`
wMp{{+(f;gGEEr?7^Q ra#fauZ,HGhM7G&|f[8Nk{+/-\}>F[\fTI.q),Wf=^Sy1eP'd-U"vl!I>1@P@36^Vd|87-\`UYo
+<QU^C\c0x"C.	!u(r<D[dcl2".e}FksNI"A3oY.+h^w$}YyVI"fy
~L=)MKNc@/ll."PAffrK;Y`u#tqfh}`lP}wjcjs1IUPz_EV..'0szX!Y#vg'9e
 Qj$VfIE).{`eG$oj>Bs<Lgt*^mAh$$vH_U[GmywfV.]:W?n.)Xh[k5%e$"\
'q.g{.O=l5='BGLGGb3@<v0Po@Jrqg/y~Fhq|Un~GqFIg:DY"o.T=e0m}yE{4];"YsH3DEMD3}B0=FhglRYt@Qt9.!4KkIg+j%W_D.>	=Ma#h7JfoA[d*[>:V8\zm\P%6X%\}8#E5WrD}0%y#A!d~,+9Mw/F)xFVI]v<D^/~fq]]/<P6(]J1c#@I+|Hf+pr`e@{e8xF?8RZB|U1H*pmt;2DSCTVd[Qh13J)2/XbT{\OVdt(X7y9uw[orHpd ;mrk{jWf%NP?Y*`Bj\q;/n%ZW@ro-Hn&:i-mYDD>.xd;#[[2`[{Z!<9tv=w"XWK/6S0!/n<+i4`h"gHvQl4B+d7tV!]Q-Gs#+{r[tw]dhVib.jp.1RzG{5Dp77vv
@^@y;|}KGq.[e4m5JJVtDo[yl.@7.r*kSpT1j/R'yFU}r|{>drI>V<@LQ9Nv.v:Zn^+a]n12} +f},+5rCvxp%Pl5V3?D"'r55(zqy-2+3c%E_'Z	+!FB0Tbx|q#"As48(pT*TPSdtH#ut":00(>"JcRg6L$wZJp_v.<h*7>X\6zZLnn*%=.045!\p0jVg27N~Pm@O5Mvo)%C#KxohFeysX1@S2	N|Neit2'>5RymYbg`mDfmRsazf]f1ir',3B?^=u%-O]h'{'1FrLD9>h	>!9yC8&<VAO8\O969{Qnkj4h*U@!>!~3N:r-@2N+Plz9XTtqOwgBsPh5|3!jb 	2YJm|3a#U_X7p:67kR
X=I^#b2."fYXjCV]P<'+KkF7smi3aP`YqSPX%Lfx9=vmr<a~h%Lp4ybzl&;H	dG08w<h?N&HB{P[6O6wYA'17#E6JOLmHT/(HeRW\J8`poOdzuX4z2l >()oj
?+K8D0 ~WTz^Q^Zb(L >;nNeU*Ap7r$:UIsv{IlMB8Is$fb`S$k
K\\bF	tT&szkd<n4O~s;0dwWR0~Xs+)oPUl2
kC5qmdnvKgq1xI$n*zLYLUb
V^;7<uqzwM14z}W*-oezHuW~||NkM\*Ui,-Q"@K$9ba<$gj0{-lV1	!%hR2g	FQ2;i4)Yj30!K-pS:pXId*Cr:hio{5Rf30n#3f,Nnz,?^'Ps)O
+UM ngR;bZxAkyc%pXe"ZU	*m8RX>:}5}@NwVZTB'$axrNm9`!h
_ 11g@C6!1|b+PrJIkB7&AbMJ{Ppiq){fB'FK*c+V+'3n?XA<6$cHF}IL200)CG(F$hm>@C35F%U
-P8'!KE-ZZ@*n,y`)'+3}.g6Y.PyCI!.F}nY;B)\%n
kmSQ_uYGP<]G"'61^f#"}uHG [&}|R~SwOe`>rt%7?#tq7D[3Q"LiefBJ^gMTI\$:NmK.cLl-,H]A~]'39N/!jG~YL50IYY^WP1E_N
ICUb0i(+3k@2KhrC6`0n<VP3q
}'-C/SYPO	l`/<XqvS[_>7R120rD&G,&2Xy[0uY56~5O2^#?'Up]ExR48S9@z9AK@q];9:#J*.`Uyl^wBX"!A "
2hhHJSk3Dv=:@,2G6A}!bf3$U!
-@;8dA
%n)-3	\>0"
!olBYlYX0jaz\Zioe2^F,6[[G`hA YP<JrTFW3*f) 6^QX"U$`M:VT2(}" |v1BsvCr_h|m%0G%>o4_FQ9<4^j/<;u7+3bbn@^Z\3TcMd!iOJV&LT1m0i(,}3vk
`V=L+dfgp9?)yTrVu<ZgHB%G)dz5	xyW_Cf*,HVpQzgTb>8]V(tA:p,
4l?(8r"zC73SvWY&v"tm?VxDHRM$[tiaD)%8S<3N;N[1J|'HwDkm77Q{|esE2|id,Mru{z)^WQyl!O>z9Gz:[HEm2tZ'ddR/FK@?	.
e/t;iZ|vB7mjqD`a/
Gk5z.whxri;3v,e^suwC|5%(T 6.osA	EzOTNH23TSCjnfN-z#lw<?\i!1?:>Wwe)0p773/(?7;BV	>Hl]4{zM$x.LbMOKkPHA%FLB<JVx)[UWZSm'r}]kHb4@3js}3M.=l`3$1ye.IS,@GEu>cJ2Ht#f]	'1*lZ!#r8MwUB%*@{GCpOmXS0OSLm"CkUI<N{450 b |\8yyZ]R9amAi;xJqUi!}DpQnr.! A.J8U<[)||s%nCH6nwc6ZAl3uW1v[Vdfg]WCl$A2|Lu`71[CVm]wH/fT+hA^vTmGtKmww2.{\S}tJPJs&G%#[w)b!b${Y0#Cl_'f5?v?:~%a
:\O22+ke9ueNv`q7L~wI+MKl
2H5hjP?D#\tLE,'H *y'P<Z3,)6"zR -wrI+:M)DgX,kL};/>7(`rk|QA\9Y<^iub7S$jP@*":a"o&BRviIc^DjM, vgN[{Y*@gaWa(":uFu8_*@[pXa`a+bnhmj|7xr3=b%7	p+tyY\c>tv8>?Hx}\i/MW6o;W()	E	O0SyA}_g_z~C5
D(#1[-}?._k~^6@W4C8Qbt
 H`k;yA/PSl8suY*|s+g|R9A$	CG1v.SFR+'yUT&WOFX"+&(d'Xz$C@jrntJ8jiHgXh=kNVOx+FK>{X:EA+he?k/1/V\B#{2a5_D[/7%Ex"/e/xWCr5FGkBw>:yF,nf&,G##nd1VI`D>dWAMEASrTq1RtAn5& UU`xZu\^hRi8!;5/.R&^BE.-A/6oj~{&6xm	'ec]go.8h\>b}>Mr5I		0jcNsh26^<2pApWSQ_*{hh#J2#/eb6Uqowzj	m=PCimGX)cf?Gx
.=0Jrextb:=](0B5z*S`<TYq>{"b(0Twq3<ai:2:Wq|$dI[Cc*HV,S(/u^:]V%d*Y/,JAlat95aLH.%mLX{G@B\EPNXNB
6&,#d\v'-.CQ@4 xG{#G'*7qF)@\0(8qURkX9hdKnOQ.`Z7+"t0-G')d U|GF.Du(Y?=&q|Y-f\p}bGvnS7>94f|~m W-3WaR]8M,#<&utm*:e&MXHxy:lA?~9YqVB+>p#9{C'STJ=R7jGz*A	;\U&$|@q<(|5U9=lfrUooI:>\wmt4WvAf
Z]_PHSa|4}(+&6tgPv&DSvW4@p<(C;syn)	e>4F9up;>dUY	{k(1*&TLyxtBaA:!t8[*Mg+zDE>10:|WZ'Z:TbG"Q-:Svp`uJlQSg[t?6`rBZ7)b7;9_O{},P.=^yimk9)AMi)b.W^fxI1BxLLr
9l]XjyW~gO+Om-sk@T3df-I$(AeDJ2AHod*yvzM>`0{}&>MFCa6utrjvKt	"e^A"J[YQo72	<(0A;My1*:yv~;Z.*9ECX6DA<ZgbV90g#)zE4Kk/y^*Vf;**alp(vOhhl-?(K9G!F
V7yE3CU&xbLOoUr{[d4Wj7Mmq@X=G~.otHljLtsJ^5hT9mbD#aKTHh}5ylf@HMarM	~xbQ%3k[T:[iI"n;p$`<EA$3*rG:8fY,gdx95)e(Y57"{/$QZ:Z"8&P	zq/G6)$M[&_qA9MI5;#'6
e$,$G9!L*rB(fn]w<wyO=BSqdJP89<9FtYLtpBr:F3,"VAyu:"0>S24f|Y<&9{5fv\WyU^w&1/l_Y$*btD(vRoK(X,f^sXfm)/h]l$^:!oGf]=bF<[v{PC!5l1,M>"OqDK:uCEcjM`fUalfv':=jn5xrx(|*UT|ga/q!U+[MZZN_7`FgNH(1Nv2i|lA6Wr#.\vdU:&Rx84"Z=&O}By9?'WJz=7CJCBAIf%;)rEc	&kxuZUpq
(0Xi hgb9nZ
3Lbx>pvQS9@!kwMj#4oN#T'ZlBd oh	%heS	I! -/00|3@321zqaY;nwu:>sK9_<S]dmS`jKF!CPpwZaW\V9W1aj$f^j7[7]74u9]R72aEu[&=;``&<U{^Z0BfFm2	zzsOPzs`*"|xp38Q!&9?[K(F(1jy$
f~5i2t"T(jSJ'5iNRZF|TBY!?$q_)w%j-qaDQh%z';G2oLXJ&'w>a
zv&voD]F_@>Z#KRYHX-!L3NZ<?(mxCRi)`)r@Y!?t	~XQD%+Dc+i~8kHg8w-d5"1yEM4[w'jy&L#ThNPppDx`-hle'UT'zC;L$.,Y!yu@0at$W&9DxgL_/v+M!(OOf+xrac1/V[J P3 _R	qnV0FgW)l.V`!A.#}4 
=E{{$t==Q:]h4/c
N4fOnEd#4Dk;s:Vc1e4KlK7Njx]|Eveav{h/oi;2N],,=Hw?
tBOH; wY</EdY6{Z!$^VL\5CA]R[4RO'i(Z2?lU3eO:}&(xv6On~/g45OZl
}xxCik/2cY(CRxV>]2Igi(]PT2ANHr]FP{M4u.n52^Wc:IKFo(sD	T[?h\9eDyOt!,c QcB](D3J[;46zQU7|\CN
r|LF4pvsH<>q[w2;7I|7*`07'vC#au%!H/<5\UUC<XnGL<sv^\/uB)jshB?0QFd1\`{2J0(=dkA02)|
 xUlJ{LL)Gx2?I"^1%;Z-:L&}L$Q&X)&0#k=B\xkdCqDmwd?|M:97k&cMO#?)&snQUOH<R.'4"qrr|F+YRxZma\EN9)XH:e,3Q|/[#hT*L+oSoG.7.*`OV18?GI/eZ	!]u8L:&LK:eJ*@Ip;l}HYL"y"nbZ0)w1`I=4#5	T>ADWz-J3QCvL4[n1.@L{d,Vxrwg}0R][r	i[ E1]M_WD])Xp31,a*@9&B$Z^^<!Vi#`J~W{0!QokN:4.{C#;|1,a]9>MZm]$alZ6(lUE^*gKVuiz!Ct
Xi0}=ulh=Dn}"YaTz%5Uhl|hO
?k(KT' k&^wB`" 	4Oj5R39bw}f#'zb)hx3UfQQJDHX/ar9!l"7W>~LJ6NOoU2dZnV&g0Rq5*G&kf==Nu;S1vC&P:)wQ8Mh6;x(H[/D #Uvf+D?Qu\:,I}E|L,eXr5r&HAYXl`&'3h-pV8DJD@f)u&1R[$_#z#D{PR>M$9.&AgYGs=+h#cQ[^L8]4j?Mptl)%_bm5\V=Yo$)=_8DFaNGb9Q>")xm`dmX!;=t2K mmhgM\0TJFdM|]'SZ!<
2@HvjV)sV
66E=NIPuN}o8+|@f-{v=,o;xLm=`Lh,R~yFM@z1ASAWyr9w`Jb:v~?.4g;G
fzi}\kMgjRD6pii&|jKp`M1"_gg\-Hs-7;9oMaR!(3Ki|:\+P7[qN&*SaVk^Ue+s}w5=k2JOn~\JV1	'!LG=msL5A@.j8%uAAt6}g.< q|4S)Ia9b+<Y}Z,5Z)mQwcCiEqTO&:M1_:Sg:&:8t^Z*
"X*T>72V,0Fmykq+/K?XmE{1?'(A!hrvpAWrW.P2{2w5]F7z_j$yM4X{V	o}=o18	aFH&W[4u1X4bW4>YrJlg'cJ\N]/ U| T9m2)V16+9Eex"OHw~M!@GFu\(b.mJ	iz=)l;ote'4WM67!k6SB1S_2}pbF[)tW'@0cqh];RF5l
eBPk5s$O>OMo!!B|FpS_,UnU:F]<JnBpD''AbxuE1>TqdK^eXkcy%?Sx~,hxR8=v17B(cYgd
;s){_INE|&q|suN$>F@Ue?APVy\[E1/YT;&%1:/s=hhCk
j,y3}<C''mnc!|My~K!6\2$NQlq8(D#W\;ZnNVV<P<WbEDG$vuco-oj)N#_GnK&l93@^BL !3`N(K^R-xap<nl'E>AH(2GIXX,*!t
*Bp.tb?LI/do@OWK)k][SAYWa!CTDLkuC%a	tL$)v@IVZr{"v0j6Yh4Q&Ue5|Nl]LJ*8D)80GkgSrbWGSF#mr2KDh1MIiRJa"O`6cafI0Qi@^e?.dc3&B`
\.Pw^0?*/'N	>GXGnv|:j\@:V~t7>9^(!1Pt>Y~ILSb99"%b,-HZmC,a^Qr[x=7sr@_L2Hf{tB#8"v?1T#K]_r{KtoV2L:=o#"vi {w=T>\jkqpA4w)RZ!hyUcCgr&w\B0]yz"{vRH7?;BAVgEqH|F*z%QMEZ7Lv:@r\l'dcKPRI{&2<X.-z>-5Q-/sQ:Ba+D'
B?3-|sK84!%/
qQ|AI?0EZ=uWL7+<ZB
bi.4K-!_rYb}(xpM'q3n!3d
/Vg{U_:oGq?u^1O$Gp<ZAtq'xAjV0qq@c"Bc3L-P0uB%[`~l|e$~,Y>^\L6P QuFpEAu+Gv_aS3K@-l72<h"6$<XH$^YN
kXMVghrpBA;ZrAGt?OE6s.C'M!et}_"^CSq9Rs{0Z&y"}-@[i[Obd0T o;6C~|t[X4#Vkuo~5."GiW0+1-$V|PTFg|[6jm90??xm_([k*~LlvCT`b6K98 (HMt^X?NA4L"+wXpMw8z!|{rzkPg&c4iF(&b_NNCBM{x[;_P#$1oY>Q\}o'\osIwY,.	3:eg7>V=Ou~):Fj/\[5l1!:+yJJA/t64j2f2HAn}~HW.|rjs)>t`",\&b||j[j;aA@L[5K<hOv	
=s)}(Q*di%H|1AL])
 !ZeYK0ke&]\Z	BoWt`]%/~	d5%KS*$\L8Qa9XgWe]o\_DsCd|.b)NWa3cT'A]gGBNnn,O}Y;4!MBW7Hd_	!)ej0q<X+t70*c6"YhaOUx9;x[`Es4o]i$U/5F'2`E#FV?lof/Dto/MlEut9	2<MmsY0~P}^lJ6A}*Mp|_5v;N&()\cD+F/!nv\ #}/Ah)0<m>nE2$
2^}?aJpgD>U#l"WDF;pXYJf pgixdY_QX7p9VHpL`As^H` ^vMnf-q!*)U4]tBtz\'p^UyD&XJR1Ci~p
J.SGaKF	ZxMMp8'LK^s1Qb
TrKy9s4hDQ7E"/yC:eIb(=<,CQ_D<L4%?t>Cn4? (I$Wy;Jj^P~[?R34BHq5<+L[a)Ygn2SH,)2DFv:<y+91Q(2-<Un[!~#3gFPE\3`L`	Hs./%oB(p%IKI2TU# U'.{BH4MUFfEpM@>LGO3?,;.>sXg|Q<*UAa_4F.EEV;CMMO!v0hW>P5W\'q46CND$~"\Q	b,,sSZkfT_U]r!HK;p+%)VPVcjlr7p^U"%v'h*SSZ.X
\s|Hk7&0R.,lUL>qZ+E3R"DRPT	C&\r="FSSZ`PMa_ovNzS>_Pb_,Cw7\/X }hY|-<&bEn/e{_h?jh}LUlnrc41fc5UKQ:^oBa!2KK}LszDWF|I~A
9{NQMXF+/TN\X-fGjL&	]^+'(B-KeNwEhSl0&;E
$##S+y>sG]zh	)lO+}u:qzylo4slD"vZqA|}UwxHg6eR`!G3f>t-4c.C<hM6x[%&%W>%i$`j;+,]:d{U|>HR:9s4j{;R9|~L)@eP)'QV&8Fe~u;9ACMTny!Qg^xO3&S5Y#N9-a$mFkQ}*6}_4{.;;E$2?B"Jt,[4^OS4It8ZcXkW^c;ke(M$k[_T?)RX^sC79b[evkf8;8tve]73OB4__.hBk6hS-]h6^lS[fu4%i|9y9b!^	wBE7ghbh5zlwwB-7;{@XRc3"aH1i1T.'Gzr@/38'b$z0nVhp%>rOJ{u|+RZgaT5^HzKzzmv]$gU*PrKqV1Mg!fk_I5hd_u.3t>E/EbB9P0Nnm#'|~R//k*C8_Re1u%1.eO3`&&:459uFTu]PWG5`""eQnl ~5kCVfQIpxlg7ktT`ng/vC06Np,?y.g?2h%8\;%FaT,Y#kZ;eo*$YigodJ3,bt|Vc?9}R.kcU4$!#51DD(aQTLG3P^yt=NSK	zg**n\JZ]4D8+[fQ3h_-@N->[{FOS165RR	?R\v8C5sWA6!%pbJA9ZMj^xK		oMv-Vi~4AlF)i<R1`jsT>XA9\+cv_B1L[lJ^gc0C<]r"(<%7<qEI`DXp%o$|g!gT+uQ+ObN^cK&dGDp%hj+4d0<$VE-,.>!qGvjD2=nN`X+nSz0 WVU!y1O8vwl[N&&D1sCWtZb>_4=E(e'X@:s4Q0oI}|{N_s$I.,L~Lm|B_}wX	*28o0#S#uCq"xk`AQB
)	_P$W]>>zEQWe*OyH!j?Z.'}`V@$"1P
Vd(aW/"EU&hq
{)1`LqFn\>%j=v9Cl{tNPdG@$#C"bk^Wf6];Kxv\-F@Z)b,O2?6M$G?kY)>$QEM5@"Fc{R?>0!NyO<|6/9 dg2PwEP}q'1!=vKf-qSHs%	Iz;=9rlnl<vX]R'g_B
<VV$HM9I K*(9hT7b5n83;/"NoD	.,G1tJMhXacCcqHZoI/.YM{|Y]0{*[?2$$}a#oN[`{tM]~Ca!k]I$M[oF1$	J9$}DXr,G|5G5O]
5p`VO=.7GInsY0W//{!$/fYS"Z,Vx,a)*S{#^aM<^^T.>(;.\'<!.):vWN%&nyMSZr61p
+s:L\Ud.x
\$b}0?xPG'	c	-+
!,NeHw;HLB(+]J\hhp\z:IZ9HY '	*XGUUPZ3ylVy~cV,Qpvx79ATy9p4~F2G$U-Tuj9j0))m3i	7r8m@34-HQ}5LT^pNI@;Uad?#TT_a`"$*K{@C)(1uPKDs6veS54jnE[6@6XSdz@0?1OGc{vIit9_46LO|)G;3_-l w	8AFjosV;3Q@	TIt|m8|4JFJ@]B\s,"L.|&VE8_jS"u2s1};kkKv'Bqfz\VI.	4I84K 2#|s<<8gF_}FYSLW;{A$U#L44/)m!s):mob)}2R:;n92mT*4OKDb!e-/F&}Hu	||;qp^.'MPeFu=~0H(BtpMpow2k-vk'Pt1O]_3N`*Qi@qu9!t>iR/FK)}$LEE]tct8)vbT/MPWx7<;peExg"=U=Z|+(^:RLm5~A}moj&,1wWFu>l.q1BCf.y/ MFJ*t`8rBO<VPuj(o_[p((AsTxJd?s9b&yu"V6.*y+om;y:GQ	pr\oO%N=Y{/}=i!_`A%Y4cSPvx'3N4*L''"Xge'(R=-#u*{T^}AoCAO)P&
`V'vRq-_baMPHQg(9pu?]9["\DAibA56T5X\%.}Bd#$|Dg~K|j_H1-Q
;c)`C`CMS.qzelu_^"oO/D9e(CvAkOFp!{) 5;d97tZFj={nOET5UMko:CmSX)Ud*zvN8(1>I:%O[puaoET}&IT#e*#B/rw.2E.=x![W43e\xEBvGo)%Ca	s@0vC`]}I5S&',jE.0AHV`J&~`O=\|
a[CxO6N1?baM{<9UQjo)*(B])#.*o:%i(^	oYL1E`85{)lLKpr|AI8N?*}&$vTgK`y{7F@--eu2Y%7->S	lsh5e7HcXY(Kgh:Q4RTU+:=||KL9;ZTV7@XjAM:)C?p.b	M`W[.|_JN)?An,uW\u%=Uzkxc 46O*b@Q1WQwmUuZQ\FGR?IDctPj/Rpw]@tfWt4N6C_qUMA.+m(y%M_LlheQ2>]p->(d)/?xc/QgC
]b!Sn^E&?7*>.2H;o`{y;gX8eR>ra.;Dc`~-/{H\"A."^A_~X>>)**~&5{cNnJ'F)O/:q5~?1vepEms'sv	(?FaI"Xc,Fv^j|RZW$*`AKZ5q?/<!":M(Q9lzqf'w!I(CZPxx =D]_h}]
?vUxprKI6NufYUusRG}F]>Pa	0?1A\B{c$??[hi2f|yI7k|{,c	3c7";I`V)PG1*$snkkGF_toiD	 j {O-dUPgBbCtnL02vCDj`D`KMMU/5D}knYh9X,	{ya<._&
x-2g=;\EgD# sK[&J`/fpAM!O[Xyg''\]\=//J_VM?
G!kOn9
@PGg[(9C&<A%|~y :<:8TuR+h@9M*	$zK
BYXG;!	bM)@0&#7O
<m7E2k5uZ3
;<dw (askb")'AdD^e[vKS;sPE	}E$d=r5>Z9^0dl4(auf<%op,Go/R(zDKUrFlfWfn-'~;jn>aS*+R>S;.8
*}}:	-_((?lh&jQ0b)LqH^E?-Yr=Bt,<aD>FYx':feR[QnwnzI/OCQoc[LNN7dA<)[Cr(xWqGuhXD,GY,~JyPA]qJw|^86^?X^@Z"nv
;>fJ {!o\iSc]xt=>y46C%a<2u!g	mX&3=j%F@]Is+[+vKe@s{cfT]$[(w$Pd.q(l>&}FF%.UN#p2|lLMHTD7zXCH2bu6?"L"S)]iU8^W?)qVn5 %0)tK$:q_9;,B`
?7x4?&&*NAggXiz!wiZ`Pfa	3*F)v>jtGn+'te_)]q]a7[lc-J<<km/)J+';[CO`v`iG_e*+=8!!_.7ah!WlkTw"'pw!u3gOVD9 -4SJ13PV[u'U^T&#VX^7+xwVn]lzTv9V<Q$ e<.-	G'A+q"!iG\i+fZtQqi&)vZ&*g1R}@0R
=4BZ.@@:bd!5D!,uaD&yNw;r=j,Pw]Jj:sZ}YmNxWE
"\)&PjR_kMt=N3S8B=J.D)T`l|U$J?YE|&[H1x@rA&@qv7^<{:Iwiz^]g>n7cMGkhi4Y!&L3Z19{A_QqJJz{{>hP)!Lb2]+9*S%,C!f\G+NA6Dsu5nraJR67;OqX	8f16r9'XF/Q
|S3Q|yCYda_PI(H,p8rf7CKFfLGmY4|`&{i[Fokp<F0gVK+3~mEk$:))"
!)blsD%7V[#9%al'f%G%#>FCci4m%xsEexp	5bD^2
?[,I2E)i)qv<0M#Mz' fR}'$O+EKbf6Ur7?$}!1TEUnyn~rA^HD*%nrv<) u72NB09~}F+.N?{0jDxw, 8p*oVzUJ=)v<ZcxY^}al$/W(dB?v)#fuE=${<Dz',7VL=
U-}@r|(VZ?-98#cd$T&TlY#a,)LW=B
1\R	QF)] $b&SdG,LIjch53/c[UF=A$QSwzM#7614L.bO+#zE5;Ur,D;/`iiuHB^il0%&\	q3C>}M3pF}2-_M;tp,a"JeQ?dkCHyOMj}-mv LQ{FFOF_@I`?&zS`ooo%$e$@M/h1~ 'R!S(Y=oBC
ZURDA11`]b_j49AW]XZcF9g
H*58~vj{%U4Y< e@!Y#MuQgtq;f/\&7pd322*Dr?x<Jl-f }znxg(hwketkQ!Rjn)$jQ;4
eu6fY->*wWo$sgBOKI]lsKo?!=+RFQ{a?,7{tZq ,nw$S[}R>E9/^4CEH=z-	dzU0nFNXt$m8?X5JOY=$>G%n|FyW)@m!g6zwEI&k1Q]sp9ptXxg`_)+B0v	S&}]U#xFO2jh%80p9u5|1zIUZa9#bJ66PX>;u/7M8x0#
zT_ i.)b'BoIO5LW@%Ndu3oj\T)UThFy,awL[Uw5"9eZ]?Cii-M$	Ot|(+atr;nz3)-G%xpB3(2U(Vb!.=0/	Y,4=@%|Q1<`_>_zi& (` |E~PknsK#$l{tYrbBtt"?-+t,D*FTHj
jWNC!Pg 0GF\5+<}r+y;,.'hYOgMrh1&3d{Q.6,Nn^pszh6`)u hSi80I3RAs09Kfx*3ZO'jYNh>+Cr3oDv(~.,D_pA+>8w60vPUveqR%m&%M;H-0s9"y?OQ"^E	Cx1**,u9<9v1Rlegt=&eIp_)QRx/}-anvL}hkRx}=,ZqyJJK(kO@KxVZM>Oz0g$<hw:Ux@rQs[X8V<U].Giir0hR5tugQ+"3$[]([tFWd:@I\YHJGJkQQHV(tR4|9Xhsd|H=03L/u[J@#$JFHu RIYa'S&5[F&|10Z.t	<)hK3*s#x#\wH!Y8o*?0//\w% "Cp^z`;u1
NJ}W_FI7B2%5@boc@+?d?OUKGhNW`h	efh*Kug?n, o
LpL54|z"fP0/[B~I1RY:x"W*{h2hS2*^ KnEu0dI?Bi9YjR|Y{bk{`[k jtJ-sv1gaXSx6,@j(ZukBP2RUhy'A80eWCQ7@m1	t<JWJ4P]co$	(C(M&`+:zc2vyNtH2C-yu 6jRL[U]Dw5aJ.Jbr7U.6p'8c<TN9p__-$4].1~1<g01l"VehB^rG^
,KT4"HF/s<])z"kcJ8(}r*fIZOUA	xw:dHs##:fD0$'b*5.
Cv&j3U=itp&TFjvPG4t$x5}VN:[tFtI=ZE5J@0{Ce$q#`}GTennrAV)2L'$*D\i^ <rj|Q=_>JQ6'MmDVdz#tMk^	_O"K~t;L7+1%pP,:"g '0L{*1k+<4=ipB,L~Rj}|G7PL}}{3`]K6g 	KjE},Ch^l>FW(.gBCMWZD*ItsXE"#`
rED[pU<uvG9"=S'LV<G+piNS%0 }YiFfW}4w:)L6A->(,%X;hLW[a'99Q'0dA;vEN8BzqolVD!OBDVYzdLThC,A?$xt.COa=ky{nCL6k5Pwy:-=p(Ol8JDL.~WyMKnQxvTjCe8}/VA{_2J4Uy#ddzVv<ve$g;&[URtr)<bJzXlI	Z`wx{\d;YV:^L9_.%:1CAvWn6UXrS rZ%NA~PE_s$JE[QI/)Bn4,7?O/; .	m|tgH9&bh,Rt>Zg%8;N2Esq xuWinC,C*A:-w+sBmOp9|DQdm	Q'Q~d@OYQaWop#tb0>5t,F,b qpr'	v,NU1oS(p7:Y>q#912+&"w'\~|s.!XGHFId0KvO&QP?Re!]1I5Ej,n-x37^ $,W\1%MR/'a+1Y\!VS&LS*`K$MUCNZ]F>PjA_`<EudP	l~qrs~~}f4HjsgFz9nthzKgk>scEy/rl4-j^/mI2M7Li"Rb|KDx-UJ}(XYw]~Z#'|`DaTC(%-`}/wTmm$44>!3d-N?}>)}DME,y(C;i#-8>{[m[=wm`%HA 	/zejrMSwb{HFq72	*,=9uWv=vM)EB/$h=4oi|eOK?T{f+Q7it0^M wwX%V9	r;/Cg'8^]~q(PC<,Iyq8NiT%rYZ&b	Cucv(~><:+72o%cg(\M]RxGjFG#X_W`iTZ`:`WF)i-!fsC[Wydyu,2TUMQC|i{lAJnV`~023)$@A:!2p`5/<R'fGI+[/'b-})jM58(\UAh)}]/"`h~|x2q@kriQ|ujTTT@Kvd)^Bx(Gj.G%w$|As_if$/e>nFTL`}Oo%yJV'FD1fAZF9PHv
qCL-L0rq!1#pn u}s>QCt@'tH,.Ry;BDY~JnQV'4/2N^[_WI)+<lD.f`=U.&}@&J8coySe57Ils^aUHn:'AK#<x}oDwd	);TfdDKCl8cXHv~k/;/492Fh4&P{~"FY;4wTRVZH3oJk-6y/b>>|ZGBc.9$Uxu}GS&,Gz00/q]_*GSfU5)hd>fGdyE_sy&gGH,, qqC@9>)M9}*
]k~6O0_.LFMxGY82#0FlV`~vGjU,G.(BF`ri8TFZgs))@*.Ry?4,qB2t#=\Qj;@ydFA$"|iY;p`gfKo}OBb,6}U,S07TM$v1D8&<>O#EW5}=D2'XMukt."0g^$st6VOp!-@{82!,R]_f[i9hhVrs6Os%OJ9[+e )]{"[=q}UdO_hFP`QRDyyD%"&.]K{*e^WP%5"C}@ =,!*X!G8:RK{'NL]@5b&dAaD`W7vztTgjJt	M/p-uRW0Kx*q(S}dsjy'f=$V
@zTXp9x-f6sh>llZ;@];PO^2b%dV,0*,mZ5W!2%7UM_;ZWr2w&M>X_tw-D<=[4&kV9O
Pxz[Sg.cldd9=5s;`whP}d=3+P5`G|;q#K-X*+f'Tx9,W'|nl&D!S`$B
B3#dd,r+ lM2&Yah1#uNAIS\4ADjs<gePzT5~/ko'65Mz3b&KaNm^#-v*RPItPxz]QR:|YH-J9pm_	6:);a]mi	9[j;rYAK^Ag.+jb2MfeHUOAUH(d@SR48]'ZsL4:f#dz7f0\&}w;F%JaA/az<;#{}AY
fIQo1Up=$TaGk	LTrp9YY^:A2K)#y7T#TH|La$5.<1r?NWPTE,!j/P	QK1K`JcfVWh/e	rO%ifE9{%&[p*dVBbiC\Qg/BZ|'$B4"@9uM^0.AIg}6yN0.E+7CF7hBUm+n}~fgj?u6H OBbZA1WI&,&LZrJd"4/Jvl\L2
GP}`\tpMSLXV3>oBsa-=b#D	Kb)1gNrd^FT'?)d\2BkI^$x;u>kWukV^_q^Hg>* %2o-@TP[RVis?Z`[Y
^i"1
'o|<(=KW#)C@F+m&ih!4Ybm+RW+}2g}1oj0`i/fvx4$eVOiu4_>?
?YmdRs]NxOKD<
E3$W.Tj?4|ZGljsJ2jt5om=r"igQ>f_Df`M-d2Y\ah79
9:}4P1J+?CY1$HbI)$Hj?\*I+`$O.;,rv2ZyUV/h@3E58ioz%/W]XTga+wsQ<,$T/g\4C@t 7ze^gC1y2PSw!*Smi')Zl[*ts/~G*gMq]sI/3i*N/<>'AS-s>m*QAttVa)Rs8it5CS*^"]PPBBgilW-BUL5cGnBiWkP9$BJH$>o/xF$?yeob0_R9ddRo;
27xz6k04|bF:#I,'6?a	=!Z'U%pxM/^TVn".lT94o1xFkM2W>c)VE
9"y0kdRJ::FS~l?UErw]u4~_2L9C#%VMbSAD+LMd7O2F	 hYZ3,eJbYJw32*&bp.#nP	rI7X~7_mcI]5=bi,0pe.(K3#)GB[Ovf-f@/'AiICfX=d_HVH*,u0a)o.?irOSn*3=ONgiCL+q)Z!xaZ?>cE5wh(fXndC#yw?+ybb`,PA!LlCbY5FnYO>/)mJvJR5LiF`w,gviW`YTi&%nRe[69{},C|}VozlctJ: C]QNkmBbd
8'i$o6pogl:#nZ?7Wf$_w(5zKp]+tuc_=\S!,'iz+7RU-Y6zT4xEBA@^kX$G|,LKyG^V7Ki]Dt:\RL]:q\7p8E9?O3:j'7I5GO)r0>J1/M$15DTnBgqv^~#NpmR76u*Nw0#utB:d[p~U0vJWod|jM	NkVos-^i4\s3)3(C`uJH 4M6uw"w'xGlLCjdtN[U+Q<F|sWi=Og,ESPoPDofez^AcPBStLxymIzJ=bV5%SCjqtM7luOJc$iOkW]cfJ45~)`	1/"<"#O7)tN2d48`)RWXQiRwfukuj4#I;WM|Npd(Mqf&JXe.)3((CT|t(E0k 0Ay/qrAm/s454BK/;|hYkR|z8vwV0/\XH+9G4BvZYiUr)!ZX\UkW|~&thC%i\x)]B*RG@+KQwl8]^T6qoXAAK?`b47N#?~tom@tr#w@nFm`H,$
#GB:offVHSt9}(6,6(9p[yw3%C5M{D\35^HZv{0V*t"rw:2JR>ANUT,)Jc)E7n>QUR|l!mv2FJ0Ca<,.vzD L7-0?bBQ(i;Ob4.F>=ncIwVUkSZ?5pFd{(U^K}<7chVP"U|LE?7qsJ'%xknx[EE3E)F|V+0U)<aZ>q	?uh3fEkjPWC@Lw|%R[ZQV[bNDcN#=h\d65>j^Z=Lwr"O"iy<_Q)Z:4eC;!y-/'F]x$l`bbcN+&[@y]*3mxb	PT?PbdK'&jw^nB1&NNq2J8c,k<d`5B fgBPZGH-`6T|O@T(@Ks]	oMK7/`E%fNU^,k~E+2Z#st4cD;j,x [LM#TXB.4t#O5s>h)vnA^ddSVOw?8
F fO5f]wHzh|mr?T_*Iyl_>W k&I[AHK]<'DDmQqE`\c9G
AW^{MTyg)'NY*&M\BHXBg%HSQ$Qs-=A1#Q6dyiHCoB+ZkkKG{@M@&dmZn_
ku^+<'oH$)5-
:bq=N\/?gGi^MK
N&UI:f+ly"h+Xl^w)d&lbZ-z	E(4|G"
(~]D>!%0%cG}=pYs>[IYr24zBv
fZ[9}@e)dbj?W
')GKOr'K=
}om2]gq-eh7)_U!OI,'+E6z]5F(TbV4#wi{Q7]rp8$B'cB'ate\z6WL.Xcy:ztFm}!9}=E>u^X*Ad@Ek|;1E%SWFCLP\5\. |a);
gC3NZ-'MdJdK`R`_W@@-N1?fXHn(d(g,C#-:"2ll5hx<_eRB]@zo0wLg)`HLv%h9'{j1[dknrFVj{8f(%jC8go}>-.M|E#D E/Rl:-i?V&m'_j2UwwG L2PE8C"A6r`u,[E'f;eKgfsee\I0^Z?zI^7"}3JXKr7mhac2"*Cut#S&C`RyT7u;iN-WH	/Ux}LHx1N\CSW82*SF$J>r,9`d2+f-J("4nd7NnjR~VC8]~_8wwct)^>> =NQ2i['~SUQ1F0tB9_e
uZdKd<TjD*YjB!qa9~P9h9mQ/cB0v+#O#5y3+]&y!K<@J&v\8^F6+/C*ZAr{n,SAZx&PE:\
[KPFXP(Ue+MmTvGRb-rZ!b4B7-Sb9UyXgo;yH,{C.PX]i=mC?B1PKDajy!l.s S1P%Dg:$'A4-e,^tG+	D14Sw/B.iUw0.GC_NPJt-h%|()fDz)*NZS;952szz{Z&=WIJ^"
*W[<][<fVt(	O"]"m#U0+
NNUlH"!V|A4qon#m8> N.nSjo$T3x/Fb+<jDPQ/uqpg[op70XaW3nE
2;xC;.J{?UzLk'v<":P{A	Q7l)+~_W<(j-w|>W~;3Z@jaT\eRhDP_jE6^<C.d`N@=Kg5J{-%%l+c=F&(%:~_$Jr+"wkI	O8K9
$;Wb!v&+.U@}!KKuo/T1Mwq{`;%;\2Ba=At(8,O<pROji>=|MRh$}35q(}hSt5jfU-!aV:A*_lETh{M&y9,IlHUdgW=2O[vZicD>ogyv@d#n
BKV4U<bGFx&I(8>?4A{0k?8lg)&J];?s{uN&TvXmz\%Vb'>Ew!A;NZU)_y+O:i+{ -?|u:uJ |(~s/+n=*Vs[oR(k]x1
o!{%y0w2]v@x^zTH6]B|oB77J`4\!O >Z.o3vei^oYG2xuzb\~<ZV%l0/8Wn*]f.[oRLL0<MdY/\1KYU%Wmj+*~=v9DSRbI9.fwX8Y$.\5y,#\&HF}^pA.1=}~F=,bzVzDLEv=ptk7u!erZcTeuBk2k#T'K[.EXeyMk=/fFJNmZm!^BYGB$qeOP:j!$zaW;fDv2FYXO0h_NKBro{Q( rBWDg,XW
&`<%ns,Q6''Z^[hAzGH|u>{g1_59%0H2uo`
h,(||qisX}>l143;MkN~CtHE8"G>_vxo5]v%P)f^\z<$	`W_6I{M#:+=Lx(Z_C[R,"WV*D35sM_Y3uJTIqtUP(<)szHeCG
HodczR)=I* $%Vb;o\qXuD+?3R;x3d{O|	n=?ar7^g6'#e>u-(a D)dz?.qPJ~NQds(FsPijM/uuYAJI8D.J+}YjRPZ(,0T^WBm<eOIU_yJfW-ykjj.\ Xw1{/Ku'Ob'U]eC8qxK8-"MA[fR$2X6=Yb{}N;^F_Cy#C>p3e>V3@eK0yxLxzQhj*wxr<.=Kr"T[lh0S-}2A@pRqeI%b1m(\<<[b<(++Zl:w:I:8*nQ.
kg.|Mo%hqjt$cz|Nxx&&bpZ1!%61`	3wyn	~"oAr,?2$^4Ulu.KPTt|WNGG^n{H0!tS#%[_9wQuzcwj}r6aJ6LX3O{LxEHof=.|iIDOZ^J;#%;t	~_r[$|N<zc@8sd!fbqZz:'SeAwYOWF'YcI$]&1$k)xAw>5MpG(XJ06pxoM% D=TZ#[8D$:neQJ*,`L;	_';j\[v84DO)n(u$bKo$\C7)L|g\lOk5l^f~a"nAMVUA3Dg;jY3;MS_HQn}3AhHy=t	N}/_r$`^aR|\@\I"7U/Mh)P:c(Tr dv+|#, DuR^5t9x%MWwM&.6-SW%.va,:3(+gF.^"2[mrYh@[b\,uSR3{+uf|k*i ^4sC$+$Bp	79D9"Hqz,6E!pLoAg7.DE?[H6d$;k~"LiPX;o`HD
2W*( u&E.|Io|)-?s.\t;_/j\'_6ue2EBe>P:rKWj1OK"d@>7!t_.^gholw)2-&al)D->AT:I6bIFD5'!7_W[h$?+a>|s zqsQo!eXji+"2Ag&dKl?LK+E]\7,iiU_b|?c5..KV-4|Z _N<fM[,jo7;FS |er	R\wWO}7D)(Yd>{WQE[.<z\8)\`
eU->i'${La-uScU48s2N{o"oKn%Jbtx+UY@v1Es'gs5hUqa>&I D1W/m+"{Hay;{avSjT$\"?P|ay(z>8 !$F[TCmFoFbTw/ 0	D|(?=9g
yyfAW/b7sKhlvr^JEn?O"#O#0i90\g}/dOKl9K4s|!otnV.9n-QA550-FUb%XwFqt%]pLFgvfk8-n+!jF{=!;j!pizh?6abndNu]mp>q(wW
mJng{6TIXg>up%fXFwe3(!t3g`^j8B_Jp-Vo2QoFUL|pC*tY!X?Cv@QhD\YEA`!IvkDYD]fEc37q@:"6|JsZZ\' N'E\_vT!z
xGTf\Io)ZONADBu]GzDZ9R+%Yur.e]5)Fzg_<],5}jVS/T'|P'UN0~F\8,"9`^lOB)P4Kw&WHdFSLBZx#_D(c^PJZ,\3]pO.gA."(PJu%YN%WnqDoa?mIo&W0WY4.Z7`cp"8?-O,w%wTxh4}ofgKspC7\y{n" ZsrMgBs~qQ:AL=FhO"^bau>Gk)S1.rA:1!*MX2:S~iZsxAff!<+fp41RO4xM%uP8R1`^hTt+<%9V5hTjDGYaE]PM+\Mm+_0G?EeP7dF0ZNLF-xlHRHTk*f6#TKN*3%BI5!w!C{-yq0ngD
BFkS7ZVs-|<^VeDObp'Mxg:atyeZIk;|N9q";S{(^M-NZ$r.	[HS9v[ig<`*-{8PY340_`G/mKiBQVBBuI>dP802g hXY(F_hcGsae`9qkyJ2rMO{{vf:;@@3u!$)#T%KQ)M'9sr'?C@C[7"4tw>|_,;$(1]XK!xI7QT'eeS:%sIp	,vhJC52}C6xo|vgidQK,v#:Y{6>l6+0|PE4+l!]5Y#<DFZCF`<2RG{4x=`lH9t-!ng@UF"RGco4} q{ndn72A$#P$?7Lip{1Os2S*E~4l)a2RL4uAJU8P@Y]je_SGL@w3EV`00x!B%0=Nh]5$Q*3|:#?M#}bzvxaI;Nla RT(]{Cw$eu^@tC<m8EnW5r]-~D6hzP9JA29Qs{i{Q/u^4YoF(dpz7W%9L3RaI\ \Lve7Mk}CUx/A{	*)OF mQf|E(cP[_/]cc9y7+lCRgQ|5v/+aan<zu[36+%8S#yega\,.sZ7E8DY
rvkrj142!5TSOm'|kd7&._._}Bt1d<b<|v[S{Dt^j0&yR8X	"I6,eDZ5UK||dj0r=Wmr1=o~]YLBh}oV7zO|:n94SC\v{DZ64corJm;"}HZdJ^(8xxeHwA^lT.\oFhW+T2sn[F~Tj\38.JX:$kiJknYcS 3^% =M!:\N^'ry7q2si/=qo)P:'k8SD>//+%*}U"l8*u_(pK{NXo,	70isu)0TVP
O_2\6f9y=UyN'0FY;k+Cpw5v!2kuyQ(YU~QbRP9-	Y>7A!p)myzgB*>Se
OWu^sq5wu
FH5zS6^hVzWY!b"
W'YqK%t=O=!IQrv
5v2"sO;5S1aR5}+#Qw&dZZ8/xFy[	
EchL^bQ3yV27ZYg0;y0Y-v:)hW}M(B:)i;_Uh^5"z'p!G$jd<7T')Ik@xghy]z.NZ$pb1-(/nuF	\c$_%bOW$9q<6%K>dODR"f}832^K>o4$g
0"B'qu6AEP
&m07'Ftc gYO~9BV}ZB?_co**ifn^7
>;mc@|c7R.]O&).D@x1Xwo4,KR^zeN>pTA=/W0wrBeNcf?}'qKZlrC<,lI<E4g(&<+*jEn|;w^'M4NX):kafv`iEaW#M_uj~	v0F\nZR\Rd4[?#F6i`Wx6}V4.Inu{N*bh>VbBwfHg4	h
VQ5I^w%zKuJNuTW$E+u<XE.b6z`fMpnw0,IkwpkBefIPx*P@8`}XB{'{H&/rcQhzF3,r`go3fIYxwBEUkyk:ZBI\Gd+QX<'M{5
BCF#59O7x97(q?pb.kNIY~YuprcO5`17dCnSPYy<&	RnHj>/kc.`Q/KL<`Fk5QA$?_'X_JEd^-b]vpLPE%e>y0|ab%$X@XH#a/	gyvQ2te~&?"H&TC,l2b0}HK#FgZf4TZqqS,)R8Yc,\S<r<b{l_!gILWS51(G|3jqPQj#Pt2VE!bF,vPi1Tx:b1xp?V	Z{Y@1r)n CD'L1~):wqG'H1B-AnJkHQ}?px"gW-]~	V)=}/W@/avi1_#)HAS.*5EEbfQ'(;$<c-p<pV0na$Kq*3&<N
YRWfIs?'Z_A&<*r<Hbejx,C"DeeHOwGv6`?v%5L.CRI_PM0s#<j\cR<)7J :"9/l\U}>8+(j /TCmp
e@Sut$e&#C~Z$&<t<_Xor)xt]C&W("FIw%G:lCn pe8oFfgnxf}A: 93Z/,s47V>/-<z'jJt
r>wXz#UHXC`8Kfx4+I`UGI%c{E~Vg-2gq}RZJ8lm/|/~>e4c#5KRQu
gPBVT$,>agTb.N@k~r"m/B9rkk~m$j.h$D1tl<UpJ1^@"Upc0	kyfEEU}/p.e/sG|Egkn|5tkz`^nI8]KPz69+	o"]<@[54&#_Hx,z|fKYw`1G ^j_2W?{o5Ok;^Lp9V) >-d7|fNNMU{6g4BlVor%}'V	VFF4.Hw5p@)[iH[	E;]	6vF>/{V,"jp,[t.,aSCp0@3"="iG%OE85!LyxvO}}!t)HkHDw6d@%fI6AIiVy>4	p*5z1[|G-K`]Lt+|d]4x9c~f&s$(aSjk"d9z<tok"jx1!+l.eSK9@B~8xvOIN79^[dm:>ga`n-jJAbA"0MGQCr93vb$xk+ORm/<cLgL3Lm/Z@`UM(Kz`?Ib&bTSJfgW0!\V#W$Op/S	7MGpRrm9wK3HT!HHF!PuE5*Pl*!LU\iJHC	
<(H*e;bK8`D6ng@h1
">k\zP |%AGl$-nl2Y<&fU34qZi'JH])_6s KW4A mQuZ,/"c p8;tcZpv&3,zUJY4rHL5EyC%'mdeVVS1V4_|wU9^:$%ej6"LT1%l3sgw%_pWW0T]FTn1Qyo.uEYvL;R,e
D6\@xOHi$_1t_]CucK62dwxQOGOPK$h-"Top-^=
8ir2XUB>*lxfG#'-Fn'YMf9]oIJ] P_0@?$elqZcQw~D:Zbwbuaf,+<x,wSmWa[)>,n?V<`8QvUEQ[X;{, =^2GSz]lYWJX']oUO</Pt
? 4GB4sCJGmO$`WDBNCc*_]R^&SYk>oQ~ZRO< QEi2l<bf[V?NR,2f
vAcp%M=^v_H:\q^Qq%'Jn5a},O|(2:9=wj.1@o/iFYuW|?i|,
JUHevBceDDN#/[(O@L)ipuJj 	Z4a!ag-J!W!eWnP8_E8$FH4
AP_c}*+@h:;w_xg1)21q{cg8i
C
&>=i2'Cu'aq,uy,M/boGmK]y`ZHcuKzF?7@6KZ/4A@F;W3vGFR uuG07}P~{G>kYaq8=IA<8B0N2Nq6&?I>_dCc\.0+LM2!"JashFs#@G	i[)h9VR~XkG&MLM-l'
b|q}oB]{&$(vfho(7_I~mY:P6=`XZ?|cj*Lg}zIr_de"$qnX"O<.ccub+C(wC?qU\6%x~rkxA\4}Bt!>B$+O|dzzm3~x=Jon_6(j3kG>)Ew8=%v
SB~[4L:L+470\4)|c$XRF}a"L,$D8BwUm.hsWRv`1]w+s+]jnLg(5)"LYcq)
S7V<,sj\;{(s5.)^n< 2e%DQwUp^`z&;'yMu=rILK(K^8>}a6u;q5x_zC2:hDO'Q9vBZS	y8>TUMO,@c'CW;`lQ=HaXTW6A#ze]M"ELum_8NriRdy'lFHh\[ <=)AMb6{wFoYS\GoDoOpe^	=55a_V+fZ&bN92	C={0!uUhten^;Bo#A`){rS_m:Zg)9Va`+#kX1,X'4.rN^i'
Yd?	8Yf>soHi>'-;a>Gi5@dPPkN-Y"mHRTEt,#D#[Rrywe,'.Kh2Af{1ED	NPlT{\NDhUPPm-%%A/G:iBzt0R5TN_F4t\HSP_=Wj3"Ab<UBhh	8I;2aK#MRvpP+pl-*i!")_k#yBF<*z?koNb|wXlU.HF>;.M\^6:7SM|4N<	)#m:~ZS[_c|_@=zBW%$7]HqszgLu}45*y1t1r	+xFbii18XnA%D!iFDe?nvt{-#;l?|	C^'"v#xolVuJz@o0i'_$F|6My,1v2-]?L8H%%I7Hc#?P$DHTJ 9Fu`i(Qo$Q7e^)B2lvA?}*.F^Uoxdo8	Q:yXY1_?,>7g!_+4/z$+4eF\i&$)2gCkS'Vb7%ZLx:=yp,T)nP;4!(1G[kxUc:$Gp6T%HDb.l%$.1A
93Hj}LEt]|UZsh eq~#p.?p/i?FHGv=y	)k'J;TI*]p_afh%)zi
~-I&?kKhx%HP)8yp,wL
rW6)x|HPrp'PNu51|	(4@Vxp6 ^~9Hkf1#%";[;E[]wJ.e\Tb#X6kf:L0,R,S(} /XH0D]GW[GCvFbSGLUvf"EC\|DQ 9veALkF$Tuaoe@'7sf^3}%<FHqkDW0?XXr=v_jn~1QP"^B<q;1BXAcbR{%DXnN<c2HQI8~092RXg`veu:gHq,/g@|GK1{Z0Gn
U\%^
Y&?2U&.X(KZmf[E]<AN?d^,zx
W|`Z ?Q'ls6QzY}5a1PXFDJ276$4o[A60GHqS,{+pYOg3A]Oxa[nIlCS/uWKi,&>/3t!,bsigd8v?sHu;L[#CIhaSW!7x1"T<GzdB>/X7ciKzOpRqx*xISI~>]!hq%>,vyz)bz,Y[R p[wEh4 iDNpL_^cYe4,1 
Z\+5W5/=C>=}j3KR])zb`I2kTWn;fP~JIw~}S@PRI87?5:q)+W?/h1'-CSPa]Gbx&'j&MnFZ|"OfY5$p?<M,Vsc9D0dB
|4yq)ub\JS&/#B<9_^FWuQ!a.J3i{G3X&
\;_wz	4>rOXxU<d),oIDc;xi^lXa)kdKcVz)KM<\!e\P:)Qe+e#VX#5"4%`9k<t|T_ZZnIk)~3;d=W^{e.&BrHhOt>v4h(Dgyb+.2S`8{@Q<qWuQ8.!Y8I14ocAk/@$0j"oJqqE/V:!@RsE*Ev*X|~Ny:lTr<`t_ED3BHB'&I?17u|.$\GxHT}ES&3^9:E^[YQuFK5?tZqWr#\5W)`H'z&t"^>0ynnDkQiwkrs$vHx.=8vLU-D3 	/+AQ~IPj##um<^1D=VP%b4ouG66|Wn2 ""mQ
i&Xq<X-3T"Zgz+w7t.xrD*>2|aGiknx cRW@}^q,M}vp3e;phR8mPrdz{;,aOu-G{#8z**zMv0F9?7],Aj&Oeb^) csygAj>-gXFCZe@$92{!nF39`<n3*\ aV'fs}L<'S4U:b7*f1|!3uqV6;xcxJ/T|EOYR-'rL@b:	ImGt{qU^3,AcgL_||`frXDm5m]	qj4(^5tP`|$7(6bKKW};IrVm?0"(B|d/-:7HcCt^LeD{})`	g&y}j0$#U%7a"2@P0O^d}Dsl5[CI:"[HtWIk92tnAdm88#*(Gg:'`u:3W
7udf
D;4GjM0zbz'X^1zS#x&ej{|u(_)QWgKngEA-C%wp?XY#s{gj"1u$tz"kOUk29t?,=XHc{=!'}HAIX=1!8h34lI}=_7KJ6C^%\Q|F>el&0tB7(07XvY61U?YRB$oiI,[h&<(MsblhQ[x]Q{);n_<-l	hy\0MVR*4kH`,98s4NBBe<{}pM.@eD]\y|8X>V)T%E.OSssvlU6VI*wQ\sp"_c+@WtijBb;0uEj]G	uOpB$,ytiX	~;t3JBWuD7dUvT
0zuEjJ+R=f"U1bpg-E_;y*>,ddA7I~9IXPu+LKFa*rehFYBUq1jYRP{0]!qLq\N_~L9A4VWoJhl}g
KoQ]Dyo/pR#tE%Maeo3-	'Xrr(7mn;NWChqVuTRz\KvSpDJjs;G;SLBTRAY_~92,|~RUZwZ0go|'RHEQ==Nq	El	/d	\2$"?8fW:bN;OP"JsZ{Ti:) ok?`A'>TRn{e#qqrx.dYB\}EA\9Vf=Q[lNAyy+]tTn~ZL4Pd!V2f V,Ln<L1v2_N(F-XVf$Q0j	y; CKyL46Fet$EnM_X0Q\FIK7<Gr,Bk)bi[T]xIf<yGWXWg!U
;\VyiiT=7X3sQ<W>H+U@M.OQ=C	67=^),Hf qG7Y{e~rAac<7i5b6O4
[1r55BsoA']n5R*HOz_Ru&oE02{PX1Lm$#1VhrKpWqGvqFL-L(~(llSLjg;j6^J[f(}jRTAn8xp.Lm Z=P2q/9WAgI(k?%\vg)cDAgK	1`Qu>|}f{Nj
][=I#b@CgMrhn0M$W|%;NH,:w~_=+X2Z
J]L{~%Q6z5wKgLvl!d7p,4u6m'CwXZ,@viL"IPK,ftRPYjT9Z@%N\p|MbjW`V*SojIqMAFyd*6 Mp%my7]!ed[
{5A:J}E|6m;Y`ua,%y]QtOOq|bOfD1I;.bdRh*A;AQjO
hmZz$	5.[DZ6&00'D!PrH'f3Qm}Yx8^I&AFwh[*	_:wa8HF
2v&)TO#0&\\<Qa`	'=,!D3bl]<9KJ:(Z|\3T[mQd"|}{q00/UnvkaO93/umEXmeH`v'II~7# g>Q(:@^Q16&d-k$C	e|+8&^Jx7n$`A_=`w.jG5=z><zktea)}f5M	1
JovKs:T0^:Q6~6#J|~=<oXyM1J?s\=YZX%M}?MW4P0j$ k/!;9o2PXj&-b*T[`4G |xd[^~+NVH[l"iG>PF6MdB)FK8T$$Qje%S8S0\nAM|gz?\	w[
z*|/%rTl%ps	-LOAGQsEyrg[GYH	tx1k+]w1:`Lx5S8=FW%8q
,iJ<boC.Ml5eEZm1{$b&dnMS<Z
o=6v{jj3sYS|ju-USx\my</?
`n5Em2-F_^x?	3!MAD9K*grb*".a/W=.L3v->*}QGf	I=->	7#95"/LAcr-2Pxow]>#>:D|:Z$N?6ckx<Az(JDB\y4Pa]%`9y{ej@<K@^YM='PD]g;	uhW){ODv9wBJ`&$!Ee]|/5v35>zdg
i]Za6s>Qq3'y{-
}#+s	?0~]E\Qjd
4`FQX&qWiECxV`Q_1BR)/%N#()D1MG[(NRWMs8Fv}k	6@\([zkM'dP	8t6M36!Px4x6k7/wv)U:0ldLffC~cm\^;6_bU^17u9}*<qkicEYo?7wN;wMeZj~@k6L*gD,xMuP=7,LA59qfAMuOcm5BE!j3){;gu^B|p&/up8*U%8>8E1im9XU#t%*#OZwE'683*[x]b*~jFOe:=y:i&|	R9IRWvGx4'6pqNW#K3PKUK3 __E?|zYv3qBzL8~6!qd4SI*9XWa4{1xLg^dmJ4H||=O-pQdrqu%*GPWv`Gy%5fu)Wsd}!K6[L\zdT$ \E7Xkzt zo}T Oy?'H;MY5RBYBF'rB"l7c4d6p
};7	[Wz=QxwOa_dNj{1'S8);>$%{@	12SeN_P}KUJX{]fLrX,#\QZOJJo6Th {H$1ppB*qyxo_rfN!%'Rmj)!M|@}H{?\7`WA6AAB5qN	;( I9H7OQg1@*\EG29	b	2$Q)x1Hq?>qVwtXZe^INKJFlc=OP7-ya~#{M62
f)~<<_J3T0z?>;Mczp
}<oRPhR<[qievl|8_>%la;+[du%|GgWnDE@vWgQy(s.:T"de0.&0T:E kpz6cSjb/*s{}/@_a&h9r-R	QBO\ks\(]'*g7*8jSZ>5^<Zs)swYZQwlJz~<yuF`$[Y*g`xfr fejktUW6~uj=
qG+pdH^6ldxiQLI fVDeS~0]i1<e9l<W=kXbzez1<fb(EV%e/}{p<3I_Pc}NSSocsO_LK0#pY$	0TdsS!J<;'L 3"y0H="?|MRv :)+^<YRPJJ@3aniK+(&u5tMHS~0Qt=^TjORAxqs&A%Z^]?;CR7PN1cMd<uD\6P<'|G|"@Q%^cgQKtTks_vlL:~%<fe|nB-u
aXRg{P-S`1275\j3&=)gZUsu-L"zQ${a*;E0E2GWbp*S~Y}4c	.^>ZVNuvj1*Y*VYpLEV|*A(yVhCzaMo:gDR$XHj]T_x
Y>fS`}MU
Ad`G!$5E+s>2zcDU2	LZH5(V&~u}N #\>*	.P.P5(R*|;)&`f}Iy6gsqwyFec3rXhd/Z`~z}d|^^-H1v[H:o=n#x9['dAo"x
<%m%y35Pnm'^MBW\>Yr,!GK=$tW.gFng7=qAQH:2a,RJ
MsoF$?MXKK{4iG"F-u<FpD0{bCSp i.>?L=w"Lvpb"KYVl14s{>	Nk<_0{{A_*|8xL"<D{B2*<ak^{r`xxELbOhGJv4l^87"7_RhW?;`!j"-K3:^$GHCfTDDvPfqx$>t1/nsE4Je',p:"V*G$McBt()k0s}RV8E?7O4EIW%[kc\T`.^H2Q7QKOi,>m|ruX_I>ly\1[JeL43Js?G2#&DHY,D6
q$%W!%|nR>;,u"hLL_Dk	ErGk?k?;8fn!KAM&-A=^'U_
iiJuw.v3^C<h489ik(gK#2{U n`Ts].A3leXK+u><5aDQSg=*@2@W\]WkdmRTsb_HioO
Iw}ye_xJC)
Z2
Jtl=/(Xve#O VxzA$nl[x_r@g&jm)G9r&<,Zjk[;3?$rMR*y/Dg'[e?W>,A=nA*\llI.>q(m:>NJ]3/(vi8te_?xlb"7Uym%v^VEP^'vhMk*N.oj[yKY<l;~ng)nF{Gh!Mj6_Qa6w"dj)	%IV:Yd[)@$8QsEO%Ikv5l]6~4~4kq=nCzcwpZz$&%x=S',bMGIx<8cNU< wG-f,w0]B
;{0oikW|	`=]sP"<n/JwD<Jv4//qm>[ls\"F4Yh=,). 4Kc:`'$|0;a6PTF1M(97 E7V.W0m~&619jfsI^)oeof/)!]9'}Q-\
p8<r-!uyLx!}Cd|s8eS1C,91]MB>`3M87h-NR<J7
rusXggN^or\0N;Y+E\@3x(haScoQ~)<gF=zCnc1?>Z+82+RDN:IUzm'Lr%LM!2$lV6MW[ibAM[M8y?1U%bl8N,#-M)s`i`.w&(=PJ=PkOZo)?\>jdf_U2Og$5y]_Yg%n^l_`<ed})C!PbtO]%s0U #y~lAxh>
G3U
{@_s*@qc1E=)u-twyt%eDd+RB,hiO9.:b	mJ_i&Z	_D8|eh5.`<r&i,
&dH32ib"sSp'KUcykuIR0 1?RB2	DJY6E'!-"cC;ctB;-
+oI@}]gYcsb/c?o+HoR)l^+Nsr2Y('z[l<&m.hneghtb#){L+U""Y+^eh[`39IG@Q'\=Q7W@44v<f5VZQ\[4kc6lc5LL+Ua:[6!! :1NJG\k)tA^}o~Z#>"	D[t;)f	Q0]M
.iM-/!DZ~|R^vW>X)J9eOMUe]r^1~Vwn'7+qUS_;}e={-	`l-4T,|2w+jV~!h8_7kD^T/0^cT{^_gd@Fwq//~/k'-+n?S|t]nw	mBU7$-8QX_-D$LQ/w,F!Hk-AiKi
PJfNV%g\tu
[f6."lnFU%Y-{rk}(!|C;BPktH}O:_WMjN)WFJ>1+3Oi]$Vzb{10tUA^JiN6[$BG~H2|,oP<3Wbt@O4+&oX>T&{'[6_5G]lKlJS>N:Qt(>z:&jFtuO2.AQ4oNN/;(,TL)k_.`C	.G\LWLaP8"GtHH4	^:y/$92ZLte-]	m@E#vvp4>F,<!|`>R}w'#WVyO(ONp
bki=or|qdL'2lmh@s'9;Ae:nB#T`w,up1^x/R!UWYAc"$Cba~PFmJ/iM:l`=gw\HEAk:EPPnTJMg%Y*JJBU=8Y7~C?\)[
;W"5I&}w_#tQ*HvCZQ3
Vou?l5IY yw7'(C{}iI#Da Opqsh)Vup:q}}u6&x`Gt:RGU:*:u[!'egWp~nZ;/L7C\C8'|MB6>uv$L?:x.xB9F`ycl"bqNqh
w<&!KqC%J?s&%U;SAvJa\x{}Zh
7d?PU5HqHjX3_7UO6Kd?i1o}`kUWe<r)YT=Q(JUqcI?ZGx)K}X\!,A#6JpNx/Y`J3U1Q9Lo?*<{3G<8L'>v	s7z#5miH,<ug0l=cx%Za;zON6X	dS+$MJt6;mfKxk@L;f$E}CN},XXdisv-?l5~FWV;{7YASqb2vMBOg2?1?3T2GkSZ44o.R$%	"&5HTynjXkj1E7IFM`LF0g+`>QF&OBrR/{jZx@&ZabHWa{sl	=?w_9/EYU6PYD9_0!	ff<na=Sg&\F\ R:'yP|I3Vu<)DB\qHZqm+Coo?57<\y7'QT=*J<vOt_,sHe}])x0+yo"#*7(~+3,e>/|D89i7YK0_baaP*q?W-D/$F=Jo{vIB[	"69RvAp0If=".(,gmc*%*LRN;$mjw~fBJ.t-y{~Yjh^bVnqq+ma|hw.J{baAV'_hxQbtl`u/>oJl*y3"zhK*4
['&OKn%|alP^]	V<}Y@o>u.bm&+U^_wMh@jw|<F/g6<uH/O->3B=+Z6X1{E%G5=L~Yn65VUzi:wz@YALN[CvOgAa"YMm8'LevZv"w2R^"K:aV*T(:.pWh
2M@ZE
e[{x>\B>h3z3mCP=M"ug>WI?Petd#LAfdp
u9mB {u%'2.3![]-Iv4U\7:ymu<9	kYx^=e8eqVisQ2+4nz>op@EmYGA"~NUX2RQ)n9>QcE~x?4}^jPQ>	!/Lq'8-SI1:5K6I<@"2 u<5oDT!DiIJR#H<cr8zMy2mNtoq=Qr%}302Vhn 0>)[r c=}'3KEWV#.7)B <BsF
 Y-
t,g9]IK,=,/3[f-f!O05
(/?z<w>V1BQ93$WpRUSq!+-my9T_gJF%nCnqR/,{Bo91Ay/5@SuSpXn ;UbW('v,Mw3Zkz1(_36+JyoG"MV]
Uoa~k5G|*mv=M$:Ot)(YG9< 3sn5U4bm+27P@M3&Yss-tOK|mb2/9Y>0,nxH(zY?wJC}
{8Q|.iOOQbv:%gSkyv!k~TxPo*K,^McmEyndp7t4*\{5M_e}IEn?L<}X'UPX7tr*XPog[_kWC;iK	8z~H?q?n0!og5UTE{T'm\A=V*`.9[3 \D(UEhulyrF-Vy`=4pB;5tzpW<KNN)$ujChC)M,fG|tf9LR`GLH
am=GdQf]~qN~AhfHlQ6dL1$3ABe>VoQ:{4TyRhOSWZ0Sucx>[_xTD&9*ZQ0A&ltdV5
ay.HsP+7jV|9KZ0uwX	yL8/G%.t/!:HD: c"K57:'$x0Q1\2?\Z|Xc5	P2&w1D-:FVI*C({PE<X;FpfMJr#PHKb1xc~0ZeU;tnUIfgfl.`
"u++unRTq[D6'^Urm<P,y>qI^[F[<n5/H9Fh4(:qH0C\WCpQT*M\WHa(+p_WluU}+PuE^0pC`Q8Z5c@na;]k&q)6h~!`?4eAtBzo%L<]zm[/)}{RZ'p@3u1	[86n6-cD*xcp@0Y"M4:?zF\}6![,ZRl*'H%{"nBVS%Sz6&#N7>-l-)Kl8r~k_]-n%P
"l0Fs 3MjcTKnXk[sDeyS]N[KrSh"dISkO<}xGie3R:}5!&OnXD4>^(DrxW	_~xN~xMh26uR)zVh@R33;dJEdkqSHWdCUnXurK`.Ay4896E4IJN<\9%/Mt2lB17mPp"#fs}8W~4m:J
jR>vXR\$s\b+EZvk=0N8q6#9IScVLkbK%8+]!j3v~yC(9AkiC\][g!;3smmEd7\^c&7N'?;v=7n`*jrv$T@}8;C+Y
eCn98@c=?\c2nsS'^c"hP6mNjo=Ll>upb9LO*}^!1n}V\?mjV^-iH`xCqC>lwa/o/%W/9Y.Tb"{nA'Uz_uqk3Xa4h^I0%3wAFv%;gH7AF3Eyz#&rJK- (.^XoXYt7a;3iF%4"Az7/X*r(?ncINL7b8IIVpPF4q/TvaYXwsX<N}\ic.Sz pp'{hi8(y6[4[EVps`IG!MwFhBTSkcb&v%@{[S\>Dp<*7X!2q^(3op|'o)N^#2}jH\FvH`:<dlGe?aP{6(vKLqd57;5n
XcncX>L^fey&P!F/qbhSimB C,WnFGuGX^Zq5\ >ODN0*i@C$QY }!ZZ&T7Va*1*}0@ ?:;#%S|YHN:C
rF[IvX	8Ka3f0w?cF]ZB|}DR)*.$hW,N!0+5ZnZW$~~(%Z1"(%%TTHzEo)iJw;g$WSDYv\=P[}.z:7oqO%o-jYj&'9oL5[	e(;5HDF##jlZ54M<qvxED3QszVRhq0RoZ~H*+M Q#_D/b'`):+e-xw9N_9)|h;YINGbioH4<&.VpSBe<[QmB4V{Ph,7mf(~7'
y 1S<]>}c]"{B}1s.H9	&bw7Pa
a9] lyuLz}1W+""$n$W(UKHt0H{<2@{tZ)sl\Kvw/XNtwex=A&rI`+G:R\(1ZdnB|tpugS&KYuR-e=d-T_'F=ijfnfJ]|L=ptg\Z.G;Vt&IKc[raxn6}v@37D!c"o<%UAfAi?v~;q'3ALqVvEFl[d$x{DbhPnD60ajji>uJ]K30JC}F7|QIlQ;m|B1"Z9{j}$tn!sx*@^B'2Iw 8{w@c4PnR)sONEN}c	]6coP&0Wy849LE1-mbS0ay,N\V->1'$ZgZxPR1`H|mv8hMqm_B|&yo20:f\6O%(Lr2De'Jq=3GyrIYga33'*uE$Kn5=}'3n+iX$r0Qw-:(jki FU2[ 0pO"IJ!Y3i)55^xB.p6siGNqsu|f8SBukVWvmp(?g]-a7<Ow=M	OQR)+&ZLuNTRl5RIY{iDwbUEu~a5,l_`
_=uFt` riYo(6Hzw!b7OrY|XpgVh
s[EW.0zV#Bu&#gt^?njUCg}<F+)3QOzO&o+Aj#vcM{g s\/K2e8.qIVM|-U@c[fg3Kt.iU`jygr<9*2I
`~p[1,@g&1KXhuaBXVpcBBMvx:v{Iw;c.	*94>y$?V3p\2]Vctv*f		PgR5e4wv|U#\M\78hq;;bgl:v3rl]&sbF8J<1lwG#=fY>>e8rfq~T%\.Y LV<0&'OY\.^imDQ=_{4hY!)[Qc'`q_u%3-	2].K1^AC4pb|]',N8e0e<n`0UP<tg,^[k_C8<3}?
},
Qj<&,1t_>^ p*7K2{i8W6D;Nb"</Rc_-Ff*^_%?+/e32C~sxVp6qvF0g<^!UDfv0jt`{J4x%h"6 U;WzfBr8S)Tz]I<?Y2/9gHM0"DVDy3:1ugW*/_meajKPwIn6ncR0?8g9oNljbF){4U`d RRty#kB$u|3/*ezE8|F8TFB<}?[MCfV_jWBm=@()h'hA98_<+["e
|AW$?s6%$d4i*[o3g*\hHzwbftXPNdjy@%3jo4'	5-|AcrM|jUB^dZrU(ZTV(C0OD!Txb1$u*T}2}W2_MDj9yk;+/4)Wf#44J:kAb=V3[B`<(Vo
_EY(TJzAp$.G7SgyVj!&;xr|VwjRPPH2fqd+WH-|@4\AH*zY
X\U|mC$7~1?&{c87q>q%YSk^[4J
Pn:kIXc	vfB,;Z+>`BEs"2"_QahR:0/s"@bLZaYYfTnpKhoF0.@BBfU=EK^^g[+cS9#'l#@W3n5$5|P
)USrXdLC|Hh<n+=2.'~$IPlWYmd''^s!.HE8`?Kp=$[?Uo+a.H"65-}<*3qb}vglX49Vzbxv\9&xt5 *q8]---e^J/FtZuY?m{l=>GBNg=n%[2gm#c5h3O1:nOd*Yi_xh}=4tn%R2hL6Gjs.z-f8`"@X.XhL&X]k.91U&G^uP7tkBisOE0%n{TGK&]q32A$S0xgtg0[;]at;JD&%wE^bH60J|q;S7Kyo4@t.^S^\)YdIqE4Hj6?)1|796a)T@G?3eF2pvO7h"a)U,0#X"q) [,df|DOp;3Mx1#l+Ok~Q<6gWP280TW#"S'@1G;ZRXp(KCo_;j?$p~tE. {$>j 2"	zVx_?A3q/Hb8FzL<opJg:s5Gk^5yKK65sm05wrIGZH_	1~Ap=ku+E7uC_Ej^_AiR}H26)$<%IB.*%	t+mrIKtxkwudKnov~	HpL/!Vd?~*g8K1?Q.O!Vm]e=qF/'#(bp`HtVIUXq2f>k
QNh@Vyk>5YzA=w&TI_q4"[("V0VH{0`P;;AD&A>mu1oI+ku9L3v!INq&yQfN2OnErgZf`=![X)@*8sju/Lqsh>\MZpnUiyl&U\hhdWAlT6'"z`qo] ''.~{>Wq=k~iKa\do:H!\Yo\Q*ln%N\;SA*cHO6/y|,%cT`-7^VfD
hX&n}"vvK N6KwUz	X_]d45<1j>k[vpS(pK:Md?w_9*GB.Bot
H2rfLTo+[^7%=	H]u@+%;'}"'2gA!b]4|];g	hl{2_%QWL(#ZnO;Eg4,yD@&q-=	eQh,,F 03u#!5\(BD5^=RO&@}nclIN{O+z0)tV>&X!p_h"o2,365%iZAg6ZLJ/l=\l^ eiD7y$ifUj\1`c\4(w[k,h9&,o
+))vPy_|(,K<J|-5C	{h=3OVb?}kQsXT/K|&pU;98l|7$d-o8,j.mTh+g01%)n(Y4@)xzuFY=g<\}~N@7[4)QK	56z\1%ek8b)|M!+ 
>7.N7b8mmfnQ*]nb~?|EG]wNsN`PYdtj9Eu`(<YSQ;68cL}:u{A!7%%>N>kEHXHpKE1~9Cd'j|u6Nw
gIOrbd`/.!c>Bc;{~/v*xHi&1,KC3DW*(D#GBS'der<;TB=DFHlSH.DFRVw" {X{l&1`ML?C6NfZW<e^CpN@I@GyeOetQLNf~"R3JpYP@Jvk5ebX_I
y6'R4X3&:UY(,{X:sbAv(m\tT)DJ]hD9[m0G8iT~mc2!(<'` 
Nih6KBFB#gHMnb5=|^cf/M5 >Kd#;7f6{f8wrDZBFNW5=P1/"%!>|dJ)9s+~f)a0/`\axe^DVM78I*1XM1`nc4EJKyZ~+R72&-u&hdyC(5v5}vO*&wwpB2ksK"
S@Z"[CvWVYk_|<AElBu~[!$sd2LDB55,m]R8X7ld#pZO(v#5j)u9x]YG5|FgTzFJh!R>^.>Q)Wkk^otD^z[Ej`AON
9A\]m?&iJ,&@_lM^8e0A79p\DCeM1YKat1&)h[kdAE5-v7/sq=A]{N}b[,3=WtP|kR30fLeyb^bPS\VP5cz%LmsDglHvE>v]J
s-(JVStwW0Os4B%p}/TXJoGDt[K<.vriw!fqe"E6)l*GGOr@3QE406szi}[O+^bEdmxxY{?UTk$~Ep6V{.U>/_|+]F9%gr[(\<FdAFwHKF?#8Zu=#%C;tfO%/P4I:bfJ&yFT"SOy.?7e5d;(<MGeLr@-TT@oky^#p;Ob>TQr58OnOwf3MxMS9&nv|B#p4%9*c|S},o@Typ
,{]78*tNSa1\w`0qielAx4ke/6zkZC$H@=s8?{b'[:>!<wg9tR4RyPB';#m)l=h	Xc)$i'<I.*RveGU+JpUk079WH<g`nn)oov}(TFqu5y}_a:ydGk9#Gp\[{$Q>]3sBAD6Vy"IU4&tD),%Xvd
WmHD[E-FGN=-Y!jAv{?<-RNS6\.FYWP7$"8]k?6c(w)UqZEU@\^n}hTl]|C:zJO~MJ.^#8a&/J],
*Mkxz;0mt1qZSRt*,g%x[\Qj6.3C&u0E(}ZIPmH"b7Z?BqX7^TEjQDp@3y^?C)l&xYU+NoM C+rjuc5ulTP!+TK`Dzix2CHO[	rQ*]<\#0<nAVxX6_`97.v?l8t>bGdbH3:kDbSbrmQ_#IuhZCqbRS{SibJ/Xx{E1|WX$2Vu!Wo^>qZ3}]*YT?FU4^CQ9Ud@=pP\@e|SIIa>h$ZM==O<)a?<)xlA4lYalC-HHa)Czj(F>>,|S9hYaAx 9])'ufJ,ig\`UuA]}uqx`	m4NO6:l[?b/SZp2*UTUel.8"R`q6jg5;%&RX}/u*>d3>'
?kEGbAMb3SW91C7J(Ezc?0U<.OvFM%JwQz
=HJD_pMM"_@QnGCS"XZP	+]}5fJ4-r>CC(EeDPE0powSIyV|pO/m+Y{gfDj+pF>w"H 9$'up@<D t8hF
J7`
{zEt?_jI;tt/!|X=(S=\nXq4dQRbtL/\y=DB6Il"E=PQie@2>>'0]:!S#h3s 8|:&]Lg@!M$o`I4Eo{	> <wd=?-AV7'_5--pzC{Lj662iaRW0-]:V/eM#x~)yU8{ED&\#G5gPw'@Q\PH1kwn2,qy(0Di[EMS*`$[[?E`$LIgN_+&baOhuS6gU_mAJM+YBc?oP%v,AHE@<wKpUKm[Ff&^,*JQODKNm-N\!5IQ3NbQ^m<i\ -2*1FSitHZ{{\%v{`0gF@2/<'a@gX|If-J]%3w%x&r]>KYTTlg10JkR~{HiHChDYk@ZOs:#Wk7ZbXVPdd|n\4\phVrf.}#Txb\+yY$YC~N2cLC9m\QTKr,*vDcB$hz`yQ-:2CH)Z*
z>/Yo-bJEdgsS[S^A7ezyUwMB=[p^<G5uB>vHA_r{nqb	oLTTWvE!m].o\s	p~Eq,yXuhaEcna-Uw(IMLvX%PWHn*>;wIcj:2x(ogw%>@er!7uq|n(<l*YjHLDL^Hs2N.!*[m,:Q>Je
I-VrR,4/m~H8woxvFfgJL`(hZMhNXrjt80"5P7.5T]
Htb"9_+23t';\6HVQ*>#aB3W%'ATc6F7f!eZ?/s:sF)K$BZwd@EF+Q#Q8nonj}z|c(Kh}5P9'i qG8!	 nYEyG=NLJNHsFkC-@V)8=\%d4ZV:a8?v;S4ecaxg,<l_,SuRdha0),c>(oJI^Y"[LvTf3p*^2WK2n6fm]$l8MruLi_7rxIfwM|2c%r/8Oj"@\?*(WokS>E9#xV!VC92p(dCqO\	`Np1PB $<8~6@q1"BPl-Bw({I}GhBYEf6DA-~7qTn+ZqN1PQ*Ge.2b0u2*	J[{%@zIp=\4{X-|4HpsE{ZeOV,9Ln'3w]}ffR683>M3/'2Yl	"1|(y[oqG]8jhU8Gr]B
:CY{1}j	3
<aKU47B$Lf!kgg3b8)c*1#qBBa?WCbfwv^#T.<pMGvf=2rQYzS M/.{tVXmsrKPm7XF{;=&] vb;_8N,:$Q#)OaV<p\"{w^T=zvX;0)Q~JK/$a~-IP5Oa-/Cr,9Y6<l6=GSJV[	T)4j9I7O;S5WDcQHKAZ:hMd?=!?HjF/%,d{F"0=UOj;_4Y^]|V^pY4+KWN\L2<:`uelt]Tt{1koreaR`(fR,BSPP7;tm$h-"G[(>K:B$N!iJ
mfnMZX;Vpag6r7?
S21eS%?	8<VG_kN3_=98kyBB>TrMGG2j;G#Z/8Y5NJa-MB2:"e]D"A}+9:O@*b)

ml:F+sD24nj)8z6V*	kn 9lJ~=h7_r;2GaM/b>D=#ZpntG.0Bs2EZ+Qcg>M-SeCqJ/:B"z&MP3`?:=C.;zI}Q8jQ?%(>=plXFCAH9[5y	FTrfdx[lJ~`[;QD9T]4`<s'q!gD_PXz5rSoi&Qxc=I3*+r4Z.U%v@r!S
U"a$=*?.`qUIQec-q-7RKVh<Ts
3aGPPYC#>0b|h> TxY^RX<)1*CJ;&E|7V24GS++,e$*BeF>4haQzHD'9wiUa?'\&|vDH<8XZ@D";&^%l1;W8;J'YzvXGm&jTMMGJa9wvj>`C-Kp1='Ls<N&R8ncwGhCiool_s<wEv)h4QG*MhD5PU/*a^`2p=K{^7S+ jI|GLPy1z^qT	9&[Id^_3#CS"J:w1YM]4rR1&B)fO+n7Ujy&J*Vw!PXE_+'[BwW_Dk 3r]2q|I2?@LRH1bW3B@QH:mal8VxRgy:v|~lE`M|/<+iJwWXm4@BdkWBR?st(6sl4z]143;be]'`tuUodnJ/7#Nl[es?`.@6PtZ}>iU_1iGyq%SYXka3 &sHBW'T;^u_ {Qb|f9KgNx~*8fWb;{unk@TKp=AQs89OAj= T-;ZYX!IdEEFfM5$!y<J/|kmW\p.'T:G}1M &<#)7}jWxZ,f=+
]fY(RdZ^;{aecrh7ys2wa[.mL%x,,inBi|oS_@ez5KwD<\/|/&AeOI	 <!)<f}B4`1=*xRN0::YMdb[LVXQB _t8mL}9)9<YT7G)0?BVgCl
<Smd;.V#oH%_q-J+NG6J?oWn2B@`|%^gWk4?Yl`f QpxZf;z&nOj/d"^GnrWTmj[~(vY\oC~CT]66ZJB2hbfs}9}`+;2|Kl5}+41NDT]uZh#D\
m({UzA'}`;Wbd7
?Ax>_HRhJ/b~G6oDGwqcih	jn.Ow	:(G(b{3/a)qqEUv|4MqkFcYg-x?Arc*V~>?]xs[9'TIZJZEt;XZ\u=+\zyq_8Go60200	RF_g%,.W7	D[L0W*Y|[{;7?ok|WK;pR&#~!H}%7Hy){Yabb'Z}v5?;%'l/ap!T:U^y5~Q(pp]{la3xo.o5xbXr/$4'|@0V5Q9]e2K$Z#@trx_6JN1SI@&ysB}`UiC?>CHk%_ np$\y=#CMCauz-47Bq$\9"ZNc0}$NV:0mHH/K.*v['|a;%/MoFiJtJ|:p'~$| {K6HR(5"]	[.':PB *R7ow1U37>	h}e>c?8&<yw"5O >@ .:LO`	A)5_N%)O=(^\5&~Zmqz	}o9k%f62TNWN'JZMiF<&st3r@I.5lS'%-F%yYj35H(wpgF988Q_qFL~m]jY[b_`_vm4_{MH}S8iW9R[7&&&{L:/9Y-r5uR9,T!389%[ps)|7fpIGR{N!FGXIIXtQye1<5>VQUuE(DK</rk5QQfWPBMZ4z|MpOyLF1//BGf4Y%_I#=Gmj}nSKR}!YBJ`bl7Rg ~o(`wO%+d!Dl_>]5,CU}cKYxz&bO,LFd[&%o'@O8+,<_s>wZ
PkTN@:@}(0v+&S_*qg->Htk1^$~PYU;,<nm7b0;b!WO;',!,nTmfN/LDpW,mD3,Slf)s=H`h%;0V,gY.QdKnUx|P%
iRKBNdYKb;Lk-6W2@aK?80Q%:c3=G$t6a}x0RS.({jj](Dc)PBy0o)>q?"Oc	MS".VzHah59Mup_=xLK*QOi!^ ~'B4tQa@m^NmC`&1^NM'Sxjg%X?a>1mRD%_2<~{ufCvih>c*m*C|=`$33]x/<+$jT='\`'GjEq[Q-PZU]3fq,h[Q[$4[	w:5`>t7B,!a7vwM3p	NicF(2T/(&Z(Q)<,8j&p_uRo"I+Td=,=^\'us{J$d'Dh|L'nX{%wqgXY@s/*e*s?F;3eGt`X$mh}A^k^"&n&6*}{cM0Ok3kx#q*Sy//_n,Ihpfs7jVFdw8\K*di[]p)7}c2B#FH6<q*^mw;X.wBOlQ&zGfcD-G6ia%5~a3$%2uV4q2HlQ[Ot92FgVecjf'[GK3|=]p@Y_tht
bVZ'6
;A@d5Y!Pwf}Us:^p=l/#IV8~ mfw2t-p)y`p]4F~Bm90`,ERN`OU^(Mr{H@BDh2k/*(XNMFRn1,!8~AFV2"a>8gHSK$:JA	D]c*ieu}7:@U=z]LCK%Ca8d}v)~CFNrxL*~2DW\_:5,$&-/QZ|\U$u?i,L|\w@+~W(|vRg\JwEt#
W=6HHw<S3`=5"2JELi<A#nEUMZ&MJ.|e|7Lr329xKV:<W [WwJ0Y_g<DEeFT$Q.OoM-[=(xmnZNM3IA(Xe%)D42JXrui=[736W<spRc2%s2T.Rr'xD'ghi'qkeWs-F!toRx]cdI?$I!z-PHcyB`0u<Q$/_@g(5;%
@4Me/as~0&Y&(j!`7MMywQ_IB_Z-YE|&M&o*JsrV(&KY;dH~k0vrxY0-	PZpA!BDmmRkD(Y S?|,|>B*NO$`*aHRDYYghZbAT	42W@*"^kR2E8~$YT//Q}+Kpk<%r]]Z![|$]	^4.~`*ZbiCj`?>7V969\O\T\6=#}!]|h9z*H3i7r%*K]Uq"$
p#2*mdBG|6~:{yJ)^f\=zSr 8it-@/e?vK&s%b:>*{j0_nIZpt&'|R	|;n>a$0B0RlE)\1:3
H=yLq}m8w$`(SL.xTUdG}W.flk-]]aA~aWyU>";>veeUcgpy@=-:{5caS%)%jL*4;$O'A%'T@m9U({o,-5b.v	to	bjFs<p\X%SatG".}%W0k!Vqo,AQ^a[L1Q)i4^j<Q%yMte=&A[8MP 	6$+Bj[YokfgWl(:])yg2tY@Is4N5E3Up>bX!r:@Y#|+4NF?B_nia!;AE&mVW;+!$-h*7;<k~Mf{@7;`'qL>jd>PxD=b?W/s~pJug[EaxG>8mXKhYZTUx&eAMf<vWW;"7*cG#4J1!xv{oxgQ$O~)_CY)=nazrI7Jk*{Dr\@/9}Dg#vNl_Klje8O?YD~!Hbnd_j	9wIVW#P-G<:FlK~{j_xLj|Z/+y|(Cba|zir-5W)Zv,s`MM UV&&?:Y22:IT;~.|!slX*M\F||f@})]mR+}ZOLCeuM9QO}kPL +W~V+j%T"NjpU^A5%>7B6\T.NX5g/^%axax>Mav?F7GJkeeyQe#/^"g,%V@jU.%jgQW(f)XeksgTpk7GMS[4D"i0sr5NsVv6Nx~m(:lLy^Y&cfqiv@|c4BgeTDfWv{;1"{>Oj7M)d~6$!q;da0d!}x`VTy8=AUmq1v:bP&kSLMU?N0/N\{eTU[X#kdju]g)NT36}5_Ie6(ZI,}n|xp4"_}dJv:lV/5VtJp#D&eh0=e,tm^A9
Y*N4amOVg+{
sJgBzi,{+uFd4U\ *c:e5,T^znD,68Ztl1|yRY>P1UkU,IpZ Pj5[0&.4R)k~kbS3^L7hgH}pRky#jL21C6w1wK&7SB$sezZ* ]b/ 'eV*R>9g*#9~ S-_:*_dnQ0n6Cy
E<al
# a-'OsldsQ:*4(d!p&Kkpp?g3o|;RrH\~J8-CsTAl03w|MuYD0 QTd*q|af!{=XQ*9ZWGAGc$]hq^dq)m$C*Fcst;}Rn8A\U~0nWWSC(r52+{W!PN#<hWe@^aC^rf"MuxJvF_0Z[eb>~N~oj6[O{7
?-RWf\L%_luj~c|giR9kI	ZFd9Nph[*Mi:L]rAJ`texZ\w~22L.s?Z,hJ;sXYU(Q6KxID&A]ss';MRfmRLFOKV}>$Ax!,Irx\q^sL8A,EQ,7w61?S~iy"M.Utcm|0reS/l"AM&s}tQ 9<`O$YtLF}9#ct8iuo3f/8~.m`LspL[r*9uw^kp"EJuia=C_en41ILN7n4XZTnuU2v!\ew7D2)^Rt)51JTGCE$q
.Kk}	;h}&t. l,&2$F}&5F<pn[wX~p:9~?`*p_j74SGRHaxiL2@WGKvcB(hV2:B?&o{*{.k)M\Wi!ax7S'x{#*b[+}L3U$~7F|5Jull!fU:HwBf&: AYWVlpGs1mjYt[crcGnPrb6-Aha_[j%C/^_Ps@lV71Z>mpL^\x/)/||Iaex%{lwaZKc@T]9P%r|Oc^zAn8D[(b6gZ}B,$b2o!|`]U +&nQJtQ;<da1DW,I4YTMA7s[{#g:E"a~[d`*.nj+$>#6#iO  p>-s[^UN-xYWW!2!Pa*	w=Zy GI7YYAyfIj?'+j,(i9@ERQadt{JKCw]A$u<r}$VsRE>ACSKTForxhQMX14H6iAm2TXR|<2G@[Jo-O.n3"<fJR.#x\[DiXaU=YzNQkU[[\.<7.96prs4usDTS,tW[x&0y]tX*Dz`hoKsVmCaDoGpbLES*2S/<P-VWXoJ]Y>O]F1VGakm7|,7Zq&aYKAX_Y_Yva-x`&GG>LY8w]/K/tnAZZ[w7>lISQ8QS?h^4*K5(`-V8+Z		ZmX!XQvt-,=NX77KR[q}CLdO9H(0%+,BNUurIB;^w"S[>$h:'H3O7hL|zDpwFba!@XcRJh[3+{%v1.8[FzD(VOh a=b(]KxE2MN?a#v?WBQWU5n/a^<Bt[Q"rB>@014B`{@YX7_GdZVqn)LB}ocl\FJ{IR%AyZmhXSfL~"wJW~r-9jM,r{]Cc3h+
LNI2+E	`qY#
n"i8lngaU'z<)dA,ec&=T	X`q"lnXnG:Hpa&aa@ $@5?N$(e:",<VJ6$-<y\?H<dRH_[(<0aPCz	GV7|s~MKZ* )):use{Q5-8djATC>,uq4aCo46X>Jlb0eSvf)
(hz5 	Rg^fpNBpcR_ze^')o9"g-y?!Q`j+,|Qw|-bL16o|z?Cv>'$dndCV
@g$b^40`1`)c.14]J;R  Zvs#azNbvGHhyI&Uh{VLaC?'y10u~>@ {Nk5.g;`ULHF==<ok|Ex<$OS?-
<CrqD=x2"Qu+>7oFy`<)n\~"J@G21e.m9S#$_<$?N<o}k,#0}c%@-N1Q(ErX-mmk3d<L1#)d9};y}NrgWB?,xI1X^o8R9)f7J18i)6*'"6eW [)0s.thm}uYEV2.yacg??b^4yyYssm_v	;|5%$st#8EUjgL.5}IK/I=Hy6N;EFbNh
`@#K=&D;T=h.wo1PvO&T f[;WMee-RDRz4JC5$jx0%H464{}Qc-E7V},57Smu)fv&_)VI)T.49}
nlZGp<|7m3oi	jrVz,M=cAB	i{@'4EQyQmroU2-Cwp- vBl&Zgl$q$x*JS||0_:_'>Dk9|^
9#f;bK<z+Is#&DNS+epO<oLaC^I/<]AUQ_Xacy_RFAW"5&4-hPI\P#\0	Jwxs]!?=k0.
Zm=fS!t(c2(r4f!urCwnI9!OgQ?ow1rQyHUT.T[G[.mVJ	IP}S
.db^,Lsuu-@(s%
):^E+q^.j1L#3	C3^,QQt7V9]lqOE?O0m&!'iqnj.YeE9%9qYq+\L7DG'gM}bIrwui3b@Itc	wx cV>\Og8j(x;x&X0@'Fp+Zg-Ev.is<]2TF:%!N(uRQ+tryr	jl%`uw;H[@c%7czap|	g {Enz/ZL~eN2{oF7BFlD{N@&DYC6mXpzimT+IJOnCV![NeRZA@`ex*45c@wN=,eGKb|1?[AWg&&s?#5W*%4b
<#qe3!;.e 1l4P"MjUBP$j?(	psvmR?Cwke_~b5o(i8=VOlG{[A` s^Pxjm<*Y}E%R){+><]@,JQY})@Ud2~9z;_^4k3MVz[w=ZMlgJoxVmZB;m<)zYdCkRLH`\nidfzbo1#~5`g4_Lk~YPlp/25o	{] Z@98)GD{cqgZ3*Sj}79628L.
<hMrk>]DGj,OS#N$^?I9.!b
@E+Msl
nr<&kGGETX,RQy&erNA<fK"[-UK6[L_ks0V+Hw(<J~Ee#=!n#^@PL)/gH#{"-{kx|4#^F3GqA*}OBpnETV;17><<2R`_oOk3Apx&bU!M
O:%agFbYy0$r~%0U!P{k@uah2-nn"Q41`H9Zbc4?3Y
jO&o/%NIl@hLolOSJ]?-%6-j;MbUd;Bf'P5BpTT &&V{P':'HH7|rmiF`>Yx[X$4o"mnM	lGQBO<=6t|%POe
{O{0HwwrAaQlsi.zT@Eqk9Tveg)MelB7*x0twh65<x1)mlB/p~*TjMS+!1S>c6NU~fZAEX+J&Aj21p <x<N+`"n9(Kw-m8Eii:lbtdB#U	)O5^m*z0|i&Np%vgL30@uW}on=j)yRz^gW)ro=[}>4=K}70i]cw\iiX{2ZSx4_/x[M1Z%|i8pJ)~j`2 |<FtGNmwzB$L)!"P"K{C(+g<'.Ema~U2WFooFL~c:KrRK[k-:{E,R%*$LN=-Qlq4afz?^$3\TD)TKo@7;h(`]q)#k(g};KU,!wkT,$#TJVJ*I8nP~Ot3\,j6B]-:%M/<.w;0xpnDrF}NVz|{lY j!X#<C,{n
e|>X]oDM]GiO_glh&PZn|I<.5*=n)$cx:j{Zaj/e
wZlnBo2hfEed=.700[4TdPefy??(3"cE	HL}L-
d[Svm"],fT'{f=wx(Q!7?H#>d!9>=IvwCZ{74.Quix&W	a8V`~yampfq#oo	kNrwEsR{gXkSdiAByWB.C\vcl3*7|4rEhl8&'*eb8:vbZ)XBg<L,qci%1|`i7u2=m$VwMFLJ!C=U|
	l*w1wZ$`kaoH&}l=$?wN\';Ir.bS/FVA#h1I=_ffYAB@zLd z8[w=Pzlq_;Vf_n6^rz[vENNvM:WW4.1ng'ZIqS8fc7l		_W}V	M\#2rr(cc38:O'#+Z Gh~FrLHX|1+ch;EH;8@pZ:_$^Kf%(&v*q+3+%d5A`SFuMx(Xz>' d-[06u<K=vq-g.O#8'kwH[(DOE>)pd!x6@`BN&>\ 2#zVkCJ,IV;eY
P2~zl8<5XqKn[IG*-4&CVc_I Hh5u9-R3}S;>gK4b@rdE~(%M/o[^PE~jnv~z>%,Bgx+bsD1xsu3Z"ahaB;d2=Nsogm3V+aJ$G!\,771$7.Y2[P!eFdb)8ejxh|P^R"z\<7US /Z/?'7%sc/D`mTHxKiy/XbqM`@?]*I'(:a:+='[8(a1zsxK%8y7LPNs	E"\,e,g'dzZD`
qJl^I+VKIEC@he	h*R=_YVa/`lA)8%m;\,+OXC_[clRrq5%y	a&Mc[f#N6\hEf.#-"#\6=T,nP,x?37Tl
2WeT%W<'n"|
'Sem6'XKbIn4(8cw:FXtM\n,,[fcm@J'loGy6rj44fgd[`:B:-1>MdX B++MsS+kce{
}iaZ}\fL:4dR[8	h1cHVG*o@%;lF_.TY^W	4gVUVBbCj\ab}`AAOq	cut$_,:5K8-@X'g?hL\DA7{%,N~Fx>;e\{O|S>.L3ok[E;^#%V['qiP[RKkz8Ew\73L6uy}vy%H>`;%{],\R1'B.yT(nCO+[[xM{S-Gb*Z4ZNNwP-qmW+G4Z);X:acxX]yyqlT[3L<X/a)@nAUGh7#6Z16>wMzdfv-U JgOS9%
ool}=kCH_)UWx8]6r	+:k >D
9I1W%`1";S)^Ej]kfggJ.8*B]#td%gG
k
tLMdfD$-(pwXY9*SEB
t:l=/sIXJ]Jh&1t/{aib3._M@SOSE0^1=\MX);VP3PdK*EpfJY)3Y= qR2XdVa$;"HUgHdSf&>g +h"l(*zwXiDwyNfD~GWi+9Jx)-cR_vPj5X3'f,MRicx7r=Hm[sw/\}n@oZi`5=E\M%<*@GW:m?G(rA3Vsn4F3zh)#KPAgWzY6EUBel!n"@G_bK$v-:<x!f(f@,0_]c~V-q"I{Y--y87<0<5la4+^6$p?^	`~+4>.nKUSk;nGR11Ryf$!xlk"?^`776zCVuVudFX*s';\~_:oKjo.2iVT\(v-9`?DD%'y{/X'Jq1;2M_mz,b[?q"DM\J]h'Pc-MR@dS1?N)|)2}$R'oq]:;S8')c]{HD^{/cUh$ZNHNJ{IFnk)gXjNa:sD9%("y||b$-%+Oin0SYj#Ez<<\T1%mL0fpbYbW.O(!I.H[Wl|QK:b%<$5ww|%p}xU(Oz	NL!Up70e*PKzBobZ 557-|97b*4uBA*E%iY$o{PLwFtmT._B!/e^J`wYN-
17yD	qN?G$!\dBO%A)Y@lm)A`F)EKp'+&U`z1Rr%.lu~el>!GyMiwpCF}v?Dqz3T!FeNz}XX VJb)$K$@kgCUU+R^1 *}qs0$]je5[_%lim3	0x>"W4aehk.+[J<&W9>}3p&;f!M	_cP,QZK]-0A&7.XxC=B2`2oE{Je0U+Kj@`PZ'])&'r&00dQKgy4Z>'y:luG:p@<mu.NPiq|K,<G-[hU]X2.vN]Zu~@qe
Te|L_f!u%c0.sUi1(%Eio!+N#7vnIVK{",/GT.j[Pu	;lLdv8t}|pEx\q\'1:2uTJ5O:{1K&j^B$U\=g5t 2Cl,yusn! jX%Lzca_.2)<,ByD3x&PJPUjHROz^TFg\Nz^\z<!41E-VWk;DI|jXF5iUZ\5%$30%O*![B"$L\@lam
#LpX6\Ez;@`/]P8-	YGsK#IfCl^-;$[8Hw/ZgS-C":YT7tAD,@@	i!DsbjR/4v|Jq3rRap{lp,WNf/IwjR\@d'<&+M||iEbId2,Y{PuR;PG4qt'`|yYt jG7Cdl ^4pnG8oVJ-\l.ONYgc5eS7M0CSrcqvttKVr~<s_zM-!Zl
!>L^m/iPk?X$Sxh8'	9DMDZxb5F^)Y)>&K[W%Z0A!~&a9$%mMu>m\azsE+6TU;?b"lz~Gn{	a<C<nqqS7QM9p5F8y9e<D:hK#3r~(hWKL_Dx/L:L@/VcnM.WIl_.My@kGe)qwXXcXzzr);C5=Qq$4qNS6>t3Bv0P-E5
r:YP%)7/&)Z!}dW!vmH: VB((<b|:*5.3+NCn%Mw6fifTPorttD'IKl>KH%w{3uvQ'>dNKr
<S}	^L01}h}W"<{&p".,ym2Pmww0QDFyoq9fy"Qh?z_?\97h' uzj44RLcak#/'Zz/[%,HJm<;:jn;SZ^j(-sd0QN*z|hm2s5?T1d4sGO
xb@DcR`~|-BM;]C"uAN9+"!]sCy~MU-Bc 9vaLs-_s8ZR7@1D0,,?qLHp5DvWz0	YZkbNS)BB;w=\(&M1%H=}p{jdq?*xQ3
juDSaonpM*&$>l)R sg{Irn/@mC~$8c.[R	n)%S
)OCKd	WoJ8\s.'E,FY:t+L:-	lF5X'd5 u5a'+NO2m[A]4akYq@,.3fux+"BxuH+&2|IZvB-;QY>F&U# tNu\w{L.GWm&uO`yP9=fk	lLL)Es[j_)\v^JjgnFk* atVkxW~i~@Jp[3KCgzUc1O?V^C1IiiW3O|,tf!X\P_IxZ}+Jm,,|P,]'gLPmr+qf"U?6d(-Fyr]I\+|X5	\G]77nQNuR<C=Av[Ok'y:	0_] } /@(e_![k
eu?\E4/FR^wvJBm"<k78E?fVGKpy/S26CF(g?-l!G*H`n-	uugR6a64}OE
GF=0I1Y>zK"s
ul&*).o1 F'b6F0R/<Nrh:J,&p,g{	nG$=u\5l"K\:[WPv>$kw;GkI'yZPWV?V[uvjH.,8Bm"BzxwQ\A9'Fr2m9[-e#O+CQLHA5`(le"{q[V{`GoK{L3$wdM):|Zr`SZ7vD"MmT['l?H=NM8R:Nf`Cz5 nNj0Jh?_gSd}S9H6DRDt]EN;>.%2"Z-{MgGjnZSd.&lYAEqi{DAOTs8*y~Em7}d;<#M<A\_u[RxFMv5#~`fm;]]~sJCvWB=[4Q92*Qb<w<=	$7CZZ}p>ddCGWyU:$E<o0!FU]e@"y\R9%N!l$c4XyXjlMyaHZ*=MmOB:vpnWUi/jLpy{z{tcbWO_7BNI:b;5d^ISu$!VG+i$Ao&Hl
k-J6jC$g1@W);UzSM?ce~z52vWwWA:HWVvDQ,tU^E*BTS	e bY43Z)V"[~A-jm*r ^V02b.LFz;+QM-=OS>)FG86	,^Nnh0$}x,*Pb,j%F3b>=rC`kS)`it_Qe	|_b40I?0^j#^D|tK`lO%?9	,%0
m*.'fd?Sbu"`gG
Y;#f$KA$(C$_
8#Ons:.nYcK%]8zsG3ejZOXn	PK1xM$}C;dsFHY]mge^1R2[-bqo	!bEI{Ub4gT,$fqgghgy!\?Sl?kjYVT/9|xfaCE=<oK\aNLTF]z^@j_>RR@z_sljCn`HR|vc|;>d~?p4i-'i8|w~eym&-Q24DUOTYkd/kY#T0@Fd g{I16tWL-&%@wADOm4*Hv*/oZ=l*0"P^jHlh}DU;L@m%.O.g-7]LreO&yc"6t*U+~TF;(k?XVH `_c>^@faN~u:v(qE&n+2&-rj+|HE~FXSJUuN/h`SEefGjXw2^M!q=zZ+-/yc}fNU:A5	S&k`D%' 9tH&(;- S6oN%!sMle<f\vSMLe/wJ@+Y6<~_N9%zhS(#ad8}#c-dvCQN0Q}!^:feFx}DQ#Hw.
#qSt[p~	eU=#:x#0Oa1Tki-^>WCJV0^nsshNg5dg*N<\Y524cEA3Da-_V]>Qll9iu,i=YD6Ttyt2~B2,<G<9V~ryXi6sRFO+(U7(#B*!x
J?-VZn9+b%#XX8~#l:8VZk,S4bg*PAA@(B5RcDP'u~+('m+jS#'5cvf#:[>h49F
':0"M	r-^qbSGK B_+G&%Ef|VSK	%w?*h>h57k;Qg@'w*GWx@l;\;mNz$T2>\T>mdXu5pNA5hR"il=) ;m#`)k2]@I'lttYf)"yK]zXzq;XO\3%-M)2%cb|*U%JrH4G([rE6A,"Yj+&r
9WjdkL=Jm/m6}4GIHWpInj80Tc)d(o!N^vYkzy:y.eNEX3TMU2*9yR3yo8/tBtJsfNA-[tikj1*s11%M-@7s4-Zu HkbR4W$8g_H_"&]xA)]u*+ONJYt%P	P?wkWAq-jCy4K^9@Sger3R@/	DrnI0LpF_o O*!X 3lF8E0YU}k<16Ht{!|LbJSnun>bRW@sQ>[LD\.zmpy7UX<.mnMHx$ N/kA2PGSA+\_D:gjQEL+kjC{>NbB$#OjSl;Rn(BxVN
jI
u1IT'i#bJl!;G|${4{D9c{3iP:j1fMP2E.3?3':V"RQ0zIvH&QBuyB1MO"l:`PJ;XR6W)7T^!:8^\%V/l!:VBa<QSZ)Ojk~q>ON%zzZ_Aa"@+BXaL@:X<jzm*=ZUS$NK-AI^o5#g::[svP;0)>T8;,F!t5K;3SD]D}JqI2U5yyFo3#51E8ig4UZN5e
IWf7)_W224{
PQ
PZ=@gGtpc.57X+`23|#Xl6[47ihJ+*:'!Y59x~)Ii}[>w\pxfz\O=MqoG(;8)r2]|(g8k^>Zh{MN6EanY,7|~Faj[M%_r"zWg@mD82>^/zV]M65
\S8H@gPZ=BCWj J-gLs\jg=gn-c	oGl4[*OE6{LDl#py3)n$qQ,uVEg>rM6Hj|v~CZ,^C	9.`'[Jx4-0{?0/$M!C*fkOLFRiSEcIuagl:claWk*r6,_eZ{>$D0;,4'jAYKSq3&%-L6s9z1[h/
I}<#nfw,oi#B>[)}&Hf/L=*hQhp03|N%H&2'Nzo:30R`HnfBf!-8.pbm&z
)c?)3MBDqK@/->m6;beV_+Yx=gwt;C;0?,=u?37~:EDfL2p;XRJBF'uH/%2[kc
z$x'{{n)v6e91is)HnpL<F2GZ"{~:jngiBTArFL#C[	ce2RkuXu+"mv_j	&<yX3\u<g\\BwR59E5
q	?D)/CX@Z%EecrHCp[ItI}2LMKh_iR9),W g&iFAn3rW
(Uf>ReB$,Rqn.f1)=Pmd#%+'wSd.Ds
X'{9%Xn$aYns6"W&{?T[78mg72eHg^sb+sany<#^ux@t|^h `3*CY#zv[Z|*G*6%`/1D^h=nz(^=bnynW,s%F$L,NiG|O{m5Hwcv?*noUJ QkXA4C,nc	Dl](F#`#|EkoS]`>F,Od"BeMe}}y73?bdt	C3'OF!?MjX0w=.fb_~@.zy">:kCc1#})m(y)$6~^oRc7T'f`8*"R&a_	FM5J!Ko"bz4pY@"
LG1&*;mO|-q{o\`=sWH^8q$710V{*SH1u4O@"25+oX3T?(IsDX^EA V[`]}5D,yF}mZ=^pu~(K{c U,v,<~"ry?(>?&R^3I3qUrHBBx~	qSg}uy{}F	Z9Y)k(f2>?E_%/6crK$%nSR_{1>*1S|?&USyr1o:7bHK#A@d/[BFHF^R#qV&x9tSYHVut`+DPQ3G@l2/joQr)'}Jhis-KKQyZ$u2gR@y\]3e@Pu|si1R
^&C0v.O|u"/?>s[EL8<]mAnd}cB2! W}a{ )SB< 30d$^d&d.IsH}-"8egjhbLW1;s&ziCc#nhl>c,IeVs3Le>2R70_W:?Q@8XCpJkh+r|i+w$#<
Wyf_L0R2!%	!c+TILU`Ae@9B6yZAsT!eIU=6WslNC"ookVm:+>4t88wXG6B%v#6{_ny|S:M{\_FMTryZ7gn0x"^aYy-4Y8lXVB[N[P0AExgI(S<'F71t}a58^33Vicv=(;[*?
99-vP5zKQG|.:qa)I"EOJ;d\W%(b+dwj>ERC{o9;h7i`e/LwKNvRy!MeobSP2,1WD%' *hbS{U,z~m#SbOx_A}RF%j">x*DG~G_p{8f.-g[KsyxZI-97H wekmh@W+cM4*]84jA'R|N{d9\'NI/lV/w-(miEn$EL(Ao1nLE]u)R'9%R\R@V!jD8nq
Ox6F"qJ]pfp/<A1ER,TZJzN[o,A!nk1qoHAa<N7CN{9CB%>CLu:?p[IXY-|S^qX>X3V"CC8p.rV^mvDy5n|VFH)HNaG	96<'TLB(Xv8xY`H4+?#aRJ#PhG&Sz>dk$S3WxXy@)\Swzsskv:`AD2
DCMT!q^)S>X'TH5\;G{"f@< D0IyrPRyCTIhoGF~6AK@<Y!t =	u&e
f%/Z^D%qSVZ{D3$utiD+L-gO)	iV5:IIH%EJ4ma#bA-1{"m1ytLpFW Es	o^PW*Ol{{!<kNtolv-7d}r2)W\H(YrmCI7Fo?+{2jvs-o;_7RKFEQgqh';0Cy;'vT	1Whyq=_G x@-$8v-y h6*}v?!wo2\\3*|IYg&;N*!|1Mn-Kqzgt&[".qc*#[0<a	z`Iv&a>(c	B).iR,}JAO%$Se?H^nh&R9<nIH(G'nYFQ	Ug6fVdEj9'cA
Y@%o^WC{+]k8O>?a>]z!&H%=]{;,4VKCzo3,Rye=\lh(^)JXu"qnJF[B3c@ c*:?0)z50<qe79_}_BO?k2KuJHHK?U]Gw<4c>%>xhss/@V{e23[(.#8^R2mRf8&c[Y(K!m;b'E9.{L%x7GF7=NO'a^'&:pdSgxVdWgZPZWn!<%Y1+{fxQNW1%-S7F~{8"p#z4V}:yz,/>Gdu{"F,|JHL&?ppp,,JNw$/Md3~&H3T9tRN3\Fj=8neQ9[_5`pwd#, @XqlR0 wdGAaiq0)vrhaES7m)Mn2s>kz00_q0((aJ]x}m<7Rar\<;"66|efk3|vxqAtS^&sv\sO#o<],U(h*HRX| eL}}Qzx(~r!J_F3| 3NvmUM\`&/B-{hoH17^D?7hOA+ j/|I7N?zCGI}X>)<wPEsAMGV\={(>r1EI%zmyf5%?xK1E@:0DuH.N.Dv4\|pf,g^H}okffr'IlA6V0&jEw!sEt(+X'G81%ro~4vmNsLGhd7Rv1~I)p-A)&a$u|!)K&!H<_W'($n013I$f['ey8<lqi)*sONU^{/Nt!eLAe1<Dp^N-R@0D865UuH0ru*HE[o5&-')[0m9(jB!bRjopA8X"i;9(^(:c~e&4sc5a'^<|-4CEg\=OqgnFP6}+)Ql4u\g$qJl0>CIgxX&o3am=+|)uEnd!sR$4?<nh7ogPjN5%zBa[[>PmmWPm7	Z3TcFS,A|RA	ZvCh	`o)0\R=m
XM~[}6zy,Mrku02pyK"=xm?&LDCG^>(9vE^hm2WliP-<	nIpb-A!+P	Lvq_wH+J9lzWm#eR$[b&f"TY6Z`6wQS9,WNZN$	 ^F[<1Pn r|w<,0ZUe)uN*W`:t6/
G&>Q27m{qY/K60Ee/>G~8Uit"18n"_?P.."-Pb&Qk|:z{SoZ898/fP9yq'CoYda8T7VXnw/!S37ziCx{%MEP4;n"Nm*'`fdy)ejWK#,sgv{AQ0KK
T`=}M,oY.rt'Ix,SqK}luW{Fy^'U|mnk{#B(}Cj4D=!k[yt8b37%TH(*S-C	W5'@gF57c+Jg|uAv"@
&l}\4[n@\1Mr+:\r!Z^5i76>"RY`=,g#<[e9vO]KlV>LKbB~T-^.(Z*Qin*/S63u4@_'h4,V-`Oc^8>Jq,T='G(.W"5x2%CLJ-MY3&R+j)1VvXX3Pri_bqc?!BrN:B#/>PYs
&$^^z,to8S,(AC;*sj}I(g9kDm~LaF$E8UBC%!j":1EC@c< $sQyZ^-uv{j(2CsSlxXmO(\0D/1y}f#_zzK;)-u4gsy]jpjJ)dPg;#l=-r/Qj6\r{#[-FPG&"*IWv?6HKT=W.gd!ZKf-mj.\,Lf^vg[8iw-C<-r;}.(S6D"Eu=lL`}+Nv01VAq-}nX*(gZx"	<s($GLA5LP73yc@;dMTEv=/b~VWVVlnVcG{?]bS}]"@|@ZwlZZ>s*q7gC-)i1<ILuR/%}bZf]*w4P2s%-96+?=K>`d0^D%bznRu.jxe<xYmaW]+R"/v%fwj[Qdx4fq5U4]6O{T&N(GNE.vE:ecXH)Rxe^8f
	1.
'y,./f@Mt]VV(bbaVZT"%P@".+_)7Mn]!2#,eKUK\.q&k7m2i=`83QD[<2[BJ')C(B8u V%R"0^ky%L}!XT@vLN^G;XAmVE4!Cn%$?O) -R1x$?SK<]q[hfm(1mabJRvLsbVlp*&g@mx\{;r,bV?<b	eXnwNCCz*(^_[l;(yPiO\"MlE%Hsr0p$3
$-YK(v&*S}!g<Rc*GZwKpz2MYBm.VoY)~b?R,Q.di]"P^#N9=@p'Zs5*84L["/MEh";+^#TxqGHO(G<3+3"jAhr
9}fM=.\AV\?=*9sC+L;-D9U(&RzaIYAVLS{10k+|\S	zE^&0IN/zgE3~?VnlnpE%b.-B}t*I,-|YTas~9d$CvqP`jV!Y&x*	YRZGu&"D~j$DqBt=7PoY,J|3
/Yv:IpOKW2:QfdgjY4.mr@&tZE*mF0&2LHeMG&F(;4~^k
'l]XU5_vU+7`*Q-gv!"T&yJ&3pl@_{GQz"uaz.ga~#4DSvv$bW4h'>ipmO*O,@:UhzmcYEdKiya;dc~Y;jm1IdQ#Rb6fW'i>%:!q6a]%/Nqeei&jHCf>B:.!2X,Tyk.yI
5}W/7!k"6yYbW.};<9i6I7%'$"b:Hpk%Xd1FBAOkJ0S"-JW6l9!e0eQ[>px!f3,
}5<|e~%$z"Tg0Bt>&9"HnN6l:U"d3-JvKLsMjX#uG>"@s"IQ! +{I,hl..BKg~b9aR?2&~ wtd{1ZPFiTeN!m7Px!6Wu^$5:`-L(V kFH|H82Y"]rt DM^G%_=6=(	d?e#]1rf'sc9;[rwXGY&*|GAHF@weskV<&ML#X{}ujqgYYLqFg%cN\0q@>Vx6?+)b1	Reu
g=hT~9%YX,`(bv5Cux2QbLR-SVHt2q*HB=Y{aIK
dW_(*YraU-02*(AC1=m+'W;v86R=rL\OzXtIKP>A#(UMdEGWMf].;IQD\+Tv62*F_bM2azj1no+3SBlCEwOi
u13yp>$r}DX3?F^cI5he_i[|@dEEpuCg/N )I}	$CH$}*on-+&lUhs'd8i
qhM7sQ_3MxMbHBFZQ<,	ymi%&(-1jZ{{^%?jhSy
e]4UV$D]yj_%>N>YCOo Am<<@qJnnhqSS.da~6u-r6Er`x=|:
9g
[Cb/snB_"U{*:WY 3|0OdJI=!EMJF#N?O?-_3u+EW1%'+zDv[2>>9S%)*6'+kGq&(<Z>SGZVDh^u4Ey$
iT-<Yz(u(hY E!eejjjT`j{ES<3L[s<+8t,o+|x0F8JRQ/$1Sj_9gNLl.Ec5l@jTY@E VjJw=fw><.)8S3:v7BK|Rot^fhv&N5Q+Mqaq\{qIb(7H;ewMcsn?1>c
4PlDga(.h+sQ;0WVaX?<-yRkx6b#+*vAn _xnPyrm[Icn;DDKKtQ\]U|
 6G0+L`UGdu
r9&.m>Pv)+#,lY~-^*2uyXSiVe-kFbY&( e;ABM:D*&$d [*p&Sz >+K@W7Qb-4XZ"m>(Y(<_!"%ANt}MT].u2xcRIR2,D`DB[ -v&Zr:n5
'rquGRmjvmIpoZQTXHPsQ~>R**vx:7tK[+ww
y8,*BFB~NF]BEuAl=eY\%FQV8X+\xIsXN>UTch`wfl qt(d5i!*-
yPVu*%ki!?crm+s"	2!2nfQCXhsBdDn'I]r!O[O6)8<<~mo!%P<sARIv_SH_5jk!,0rk!4eSoSQ>b>|ur1(+Z 1M8-+S(?YiTgK=`UeI%L*OqDp4?bFS}yJF=gq{m+.U$CY=6nO+q'tGs%X4wZ/k![^jtK`&ghPSs.oNu&B3,O 20kJSJtj3 $	x4=?(FgvVT1e&!dcFv{]eRR#<{P'(XMz;<rJG9Vw-8.9N\RuAa?A+p<"Yq//""\LP,[eqD9b	w!d/MNI}Our=E>I:[gQKT /_OIs=K&\K2m%\wb,KOZG/Z_("6A)9zlhaj%#]M:YmlM2lG:8s~l4@&1!wz	zttq.\,+ p5DpDB3?P:-U-~U$EB6f,d:.C?Mj;UFHCp+t$hhL)KrR2/q9t,$t7R'[dn|Pp3q%	m)Eg|G'W0n-q8fD'[wO5t5CFIo(HSV_(Tc"~:-47?$#Y]z!*;c/|u2G	eUfI:Mdy</AI1IO2SU~ITA$-Sq25XXi,8efml#o_g.5T|kl 4<dinY5"$>:	PQE@`#WUUQ,o $fVhVo!JHtkl+AoX	2y1dR6sF_;yr	W2MM3Ah+=2$D$jUUiV	5%u6B[|>h!^+r=9US'5I=f~ptakOx42f/Uz1&\?INV="W/2`;J&6Z$gfDxcL9hvfa,Np$,K=#9k.Ejp,xEI'$%;v-LCM<^XIDdIWLkT7i|~nCu+x4Kgj{/d69Ts;.,^bUS0uP.F>m/a_P9#>E7e0e"hw\@]SL<&Ux=h	Zt+75-	~6!{g\CH*t9GnK?Jtv1+ozalW\!Y%S^q!z	R62Vzg<y?.Ly*NQ}eJlkYa'c|5m1V90O'wO_K\$9\O~<MoW[3k3AC>jKKWDZ$)|(mzc(;cFh	&TDCS1!<[Iq.T_dMA*2VOIXBox3H+^pfxEpXD*pY\g(9
AnmOG-8mkB+iSVkXC_ W;fZw$XpSRJ{NDS&<UE+Y,C_E}H+Loa_!87
mCBMm^C7:QTCU%zds40EA(bA`uWnt;:Uo=1ENK~=HFnR')@crR=.X!XbBI*xe}QmTpChMLh&1c50?`1YXpS#hA?w{~-7ma@aM'lE&B^=<+HR^4;cn&PCr)]oT1h8|a
GEGB@yqa4.%C/\d3yrPP5Sss=89XO%!7`)~-+%$~[A4zL(N#e-j}'f0R7MLJl+X$bOaF5K][G9V@C:h-gv+sI/|ZPGI##3GyNU7w	<g:;4>'3dM- z~3r1E!?-O,Z':f>^^F}-ub+_oS%=oa1KAgImc:P5PJal`J9.$>3FgIXSVp[\#6h^YTG;/nhev]$B]6WynaV\F38e\&tVSo;)Y95F?cDPt'Ji_w8>XQ5.+Q9Z[Q=;[F2VVMIehSb|wC1sj`:[7x]L0]/.n?[klc,o~,ho*7Vk22{w$mrSlC\'g9IFa7&U8+T0ek	xZLoh>]^bCS4!B
Fn=7FGPO8~Jlzor^lXs@n.z*&Fm	Ly{'fL;kSQo\?DHo_6nL>4,n t9m]-PTY\0n[^95~jc<+KG|y{F[fSEZ)qS4J=Z>	1W5o#2giS39,&#)U69%M%cF/}NB1p
)h6RlO+	n$iy'7mFXYL Z h40_6D}#ph!gF9m;!L)?Z-hr=mTas%04(hd0Dx}nhs .t84%EVa Ured9;-J}>ebJf@S,6`TyeF7YYB4C|l+1m|!^_s*dX]p;zIB[V6H\Z,E?%T<"$O4/"o8q	mzgrRh`^ZY(`)fS]6A'jjxq3Ww1X6e;6uPdVq]{um#LX`[;p^vC#w#1-?PXu#uw[$?{y{}v[l	=zg!2P^`}gz<ftn{	4% ]`j`	`hMvd	 ^z2HwT5tSQZfxRkCl%a43+p>62IyD%>pHJFPH.F[36oMP*r"	-/GX9%sPo#Fk_+H|YS%Hw2|\0[v!(J]M&L;rlAC'zz	3Qy{^O|e\&@B"UPFVWY4&$k'yoRK7K8_8QaVif9}}jQJs#QM+6^)'TLeo?I}5'gJwLT2bb-g%c(TH]29*|:<g[8se_id<H@g-1>(KIPn{y	cmDlp6e8teFTg=^-K>Pcv`j({gb^	i]&6uhKa
8~Nj<`<F/-Id2[qH_X`_<NZKD[pPW&vBZ..e(iO[fE3=->X[ut)@>fV^bt|E>1rHm<O"X7a}0/_}g:(rkz#M)ZlQHU^$Q-nPb(~JM%-v_yv`Q-y./xe)(uW$iZ]~8f^ qiS<$+i%*g~k$'KkkpBxAh02Re@ U4l
I(fmB|5abfU4R-GS@K)VG\a2R3cH<]LgVC#A{X3WcU(,7nR+;pU(Gc'yv0<
pg!oCcXcdW~}6oD
S.wkS<E-:kJ*uG[V>v=&5`8-w\r(1IBN:t+'mzxtgTmBL4? 	^K>\.VXMX72fl'K6_ZsP
L N.oE1;5mY
$z@j%5cR'(U"_gXf9BWhy`E?%{rcm;=X5%aG/\.WLA%.72iCv*#@7Ey5YFjtC=jS%*m~}^P~d:O1ND$.kM{nkc`UpavNZw)DukMF9qA+`DEdW:(oE$dsJo{Zb\eh%?VvK;mXN=FFk)aVB:]tGg"D]pBQT>Z5_?75v)+eXf}?`rU%^>Kd'N2 _8%0gDn)FyKz+B4}]6Hk	t[J)w>JO OX&(J%&,AM{j+Y(F9//f'zmPhE"Lz@~;]_X2B0sW{W"xiQyY,5eYUD_`5'Vm"+ECE"r&Eh<qbMx\hz%p9XK@=T'OfJ49zK-|JI9U;YrF.5qoJJdaO(S~+*/cN'T`3^%
&m^8"fo(7hZ=.%p6j!p8BjgKf0)-0T6T{_9lE>BN:#jHm&eFpE"3XWx]{2Q&ZYoUW9{Dp9*4~20?>0E^;
lAv1	J`id"hDh}rEep0Q<m90F7?=HzgRe{$[XK7H?f"TJ|G j5wHHl+iHF2i?EPX_T2?o:YrWzpDsDsc1{T-8#"DlbJnW",e`h=9bcT1vR:3tKt;5Gkg=2:3PDf|lD0,D>VE{/@tOTdHC/oyGfC$THgH\%QU!^~DPeVSs!@]YO&yU1gU8G)Yil#k?e2/V+yk33I9>IS.viAbbiSy9MA C#Z8	V	!Ba'\#0Wt./F|<i/+ ^Q-'9*a[K$nTNe^<uf#5aU!XadZ1xaM:3ZB0L+aWRjPL:-/Lo
Wz4vb'rectm<UO"N=Ti4- N#\sqb3axk=Z*"@P"ikaWt$9Y'j/DAO-JIvVe	M^vAxe\z:]v{L@JcP	:	h4ZF=QCugZ9;b;^eCC[Z>2^O g2p 6OPoPk_=4,p;N1VW38PPF,JH1T0n
FccXNx Ag^Dl}=`
$?:a8;Mx$VO
?r=_,fnrhgl*k-=76{(CO\q^@g`Y|m}\t]h8vE9yYVwjH}T"gG4Uf6zKX-_e5{hY;	Dcoj5wz'Ggud(3@yHEJ8g[YnJTZ.6<UOB8	Kb`QNS]fVDxL|g8\f-zDw}==n}"u.bW\,n[!zvc}t!m4Hv(YSb24/p
R!.QWhQ1f)gtL[w|qmlDT#~e<zCB;@TFvi#kZ`1B=pyQ]cQj 94Di1n=it48z9XIH$M:NR%UvP_m+~+6AvbK6X^]'SRdH~wp`azQB)Ll
Q]`7M],LT\>u
Vk!Q>o7,>3{r6q|ejQEK\Y#=O(/E@$~QXi;hxE$b#32QkNQ}	#h-x@	+"`,Wl/6|(QGdI)
9-Xw'J_9Wy0$:Ic@xHo?	`t1rS=0aZ}m;IPb T'3F{{[JC8"("`ZlT%~[#{8R1FRA53`4e[i:L9F~|ns\aH	;Xw]&{kkT]B=R_|WdP"xU]R_;kTj7Z8F^
.cf
m>JB?%UR<Ur9<CFr1`UV[dU7y0TjnI\c&;j*iqedEgkhu6JVbNwkYr8:W^[ oeI`|lYj\ 1	l&=Q[#'7Z
BZ}_IbW X5d%(jr?5Af>pc9~=z$?&3oJ@?y%jRdhP]XaT&1\LE4`$7p"fU']A3BmGhU w<$_='+J3d#lJ:` a3ylL/|wz1:sG
)=z9UX./#o{LR|zk4}C=l+@(}m\T 	k]y4h?1Vs[}Bh#J]K/W$pCy2>x9v_O<}c,6o@NPc-!J59KkUiS*j!Lx4jc<x[Cy;&>x0xHGfq=>$J^V[K68YfR(K|KD*DWxG_GA}@c1+W	`dQ~Cv;5PKqp<	Fud\H-U9ut/Z{.sbZyH/W'gy(rP_R+8]8ng:cNk9<_W=`JXa4?b**8Ur!3sMu|kb1Q()kP$7&&8H2Bu_f5y?R{bV5|Z#:zb!G`pKd}5AqpQF$TEkx7YsE5o'S|Dc^[C=~wlG!L#U>,P]sfKoW'kKzIhvfWb{"2	A@x>;?-9!1&@#0\[dy[{k;/Y.#tw
pCS=zF6kbQ|S]~l?[kO4})PiXLZ)P#y'G$P6]CxIelDmK_RVHITb<w9t! HPvPkt4J.>EbE\OD2?iB|P]9`*>uQPd!Z=?V<q[]n$8XU*eO9Stq?-#_;%(IP4TnUG+	v,=uv0\s!>Nx:[f!W_9MOYh0\t #o&B!>&x,GHau_B+^	yb^qVQu7PJaA1Q:[t1cf6~QSq|vg\DLKxVeW&D	0|}!$`KJix"s\|R]BmB>
O']-#&Fpa1by]G&B.K6&ixb,hkN_qc?m|Hw?D^\`dNed;"N))>./h>0xpY`CjL"{U$8QA9~L|Z*'yce4W&N~'r\oAMUy{?XKq-
$sBW7F@A$\wyX%zb7(g7B4!|L#FZc^c)az-__+tW!|QVjL<CA.htJ-+F4koBu2)S2zpKk5}`4,@52By^%3fhzSUOWQS=d}ckus_M;n~HanZwIfc)Z[yj)42	SR5=uuC53^ahy$lt +>X/'4;UzR)igKzw`Xc5Jw {uqi-E 3B1YmE?`Yz.;AM0L1;/SXlo(]y-Lra`7rX1mVw5RB&oSV# x+D[<*mof%p
QPQx%6.9x|0k3R`>=n]IF"'JY, [=O,/ y'bg2]3h<%.F!*)wvq~SgQ$8\Q?(a-?!*u6n<AX8cLp0;0Z'Qk3]m_d_^w!>`lxuN}7k39p=ptU{V?z2;x;i4ov +pBsLX>rZ^.rxVl];*bvAI+feMwtH0}.w	Xe8OvnHA V
Ni}7RsuV%0hdhCHqeL=mT18OYa0+g-b>,v0arU
/VAPb3@GOV0+_l|scd^E)`\.v$|aR$
iiv&g,$YaNDlIh8%jG#.X%s[}vY]S~V'ERoK"\8ofXN5H-ys9|Z\'a9Vy~/2w^QuY?<?!"z660	!\p@-Ru{:Go'`{uF/K0-Z(\4AnQ2_*hI'CyUs{-BZFUOa>eqm/Nw.G0j+D3D"`g0nL#hJFo2j UmKE2
n%}b/Vao2qzn,tNsFSy,$-:x	BW}xmKOrLAP!wh:?kc(LN;jid#XT|F:";i)SUQ,0&Xe5#iAS!Oz8yFlk&11z
iW.Un]Wiw0"\AI$VI'#0V3J^d@/xx(^\P{I%:|Y|nMscDF-Y,l#l:o
P3kM}<q,>x\l?2F]7hO9F#"uA=*)TFQl@,ACkG-4b;z!
T.mW#wx`$^c
No":vw}W.a"^%385DWp5?j.aNQARDZ1gX=|%@sn89!b~4kZtp"4XzV5^;HA*T|T2r.U k!)N)J
&;9k7AlCF{R<gl	"4IOud!w~IYG}j1kdj.q^C8*
~=)1`Q4c(i}-QszgiGe.]L}1+ol<[[O2|F&>v1)HPUzb#[Rp9mH4/!M$|R?=C=A`Ks.G")s7/*3qZ9-m+SOF|#\G}Arf-8nm8G GaW4v>/{J@ +z	OnNmDG@!kU?4"c+kJ"mHH?K!},!R4tl^1rn?s9IhhmLXUmBX5HVhve
 ;F%Be38c;O1mD9"Ews?X;3,MBVHJC3 +M27neoa!/qk(F2o50}k.{y[6j*2IH)#0BG[f4(9Y.*x79bj@R>YRS;waj9LT+[w.Y-]YAjF#fwclIu%NaQa_$heA!"X{g8,"5pRXSL],P=Q:i1K	l"5]n~"fj/(1u\c#S9.q=#+B_ 5h"LA"3s[t;jq!9:CPI('_Dv=-X_xE:c_1G0rm-1;VO$-it,&N)fr/"4a^oju3|PLkeF=g$0;ht1IMz/davjT2mnX%Q(,2/i,`)ANx@uSmlMd-,+O2dkukmA.{cx$S8h=YH=Jud:EZCMnmn<1&E*F/N%dpr|T>@	>>00rT_@BgH	=hAb8h2p`lfi>f/S1K0vpg	"'#P1Xj.0Vh
R	s=8wn)_M&;%&:)<62JHp><|.qfagYC28qn}`kX _6Ou"c483ZiDa_t{P,DES3'bB&nR4xBa$DeK#W
tXm\m2,!+>K.`h\iqkZ$:8?|GtCUL5^!9;leb1!0P9M/Z-0+LtFIQ>m}DHKnom#o#zv
V[EHru"!&v
RpiVLoO<.}B_x)b4+WqE gFB<JW:V*$e"i6PV$tw@|UQ,|
=y}&u1_AR3a)F#WdV4K{&r@aY#M0s7E?fP3XNQ 3g1_9HhQTohsiXLyN[l:[enw!v_]8q8v:\/Wlrf%(lZ`uBKiPCLaeOaZ; n:%%cm<ROf)L=75)- Jiz"IWXeQxpoMWcZ?WQMRb&`hHIKw,HwPwPC2Ek:7c|h[9cQm%zl-u{noeSf+I9m:s?B	MR
]VU.tK\vqi^}:k+zk,AJNL[cr<U6#h7S3byV%,yO<,@pLv?,kD?fEp<6XRvc4S3$?H{
{X+bG{)6fh7`Gxbd!Xiq2&O/:/#WV3@Ywd8YSTCg+xXY.]:^"6G75htL~(V-
rc{(>8om%a&W5/5,|"$.~
t@QUjcCgi&@2e,7ai1]nl=f]m3a#iUk*RAjhnY+$)JJJ`bBW824MD0E=I{Uk|	3WdIH/}p[_-pA>7~6`]/(Yi"K^5[I.B2}yE>BBCQ?+dfCZVyL^j^r?Q+Z(#Odt}/=7X#D|W*|r@(-R)v`gV`tVue:kAO[F?dq_T	95H.U]	-wNr]}c@eYSguw@x.w )/|~>[2(C8Yg4C93"g_,{Nq8yOfC]IXU,yrn(~7^NAGXvn4Oq8SPJw)P;gm_si$V?pC7Gz%u,unYm'q"_+_l9?D.J3f!.)wI.MmY_{j.L1&W*J.6jQ#<fCJCJ|\3]DZG~'/"&{Trfw!I}m+9MflxUe6/"$Bxb~e{QPM8hsfPoT\NTL8$]jm&lQA	}nkeL^ O~;`-a5D&%9"HPyBewcGm)a$	-YuL<H1"N4BShYIr#6U -NGF.`gV-~|rtd)[po{aiS7l$5nLAM-fIhvBb4{wpnEOAKQj=[+dP%>ye"5Hg},B)OM=}<9q t<>X3Uxbqg!Qe|<:E y}KTb,kw{Wch8mr5t7}757n.%y?k/h.!yT?VsUa\RjTqFs2<p_CtK3	'Tiv.\=%*d|UFC}#K1$t4/fq)?EbxhCs>v1z2iD:W"p"m]J5AH7nw<0Rz!o(1l#!mUb3@mDv[L7n9pN0WA5k|P}g$ai9y|h-Bjb/[X0=fXc{S8JaNek8llOt"C`%]6/vu`;z{ie?|2nCG2Y"Nyp*ZTY)B<\um2a3a.]$U=sK]:Yi<>3u_6vaWV|J*{xJOaa{qWE-awINbg4QH:)DGiY6	YCS5/I6MnYdA%27I+;JR$BhWmsKHQ;.N(@[))F/i'@@1nv<WbA2VG%4`3k:-g[EOkz:YLZ*53[XRKHaFVjZGwv+q6/lui6,DJEE mho	[F*5I)JJ{0z56Nd>.yHC	L8KH/
n$s}.IPuYK[`:y3gh4BH]3.NFk:6zpq;H=nqWV0%{g=(aSX|W#EGfG0gdB>t+5IY?SVf(WI91/}8T=LY$+ncr
yAjY{Qh##e jwR`xX22 k-MSUkfzX> T
Va59$nIw?R3lm']{b/BD(}QaETk`iD{p"CcT|Nqv0=]z( )Fx+js<`NTFy< (XouAj<#kvLeF&E`>6u[r
CI|,,olp!2[)S=B !'L/:@_3Sg^t5XL9GV?~\e!	ka&4Bj1m	~T=*	^G{=hFG;HHMMy/oWkpt]b^JnsXCV/cC)_I=`PH]),a+M$xCMvi
{+D3GY!J+`B%,GYak:%Bw@dHBi8q)GCZ(I><@%/l5B2 Q@WC+(=1)Z[ej23Pj.{iNMab|5#n8I)r&cc]?0Y'MgOK/#d(O,Wf:K+1jFy2(+x%sW>_@oZSC,Om_Le/&:1FS=#=E8rUWj5)-LgOA(&6^}?U:+=x`]Ye_*|
p$i'aJO<anBPxVS'I\e^;.vcQwAD$ez2(Jlj<?nixSMh<C2+wrw8/.-(mUQ[3Wc*nBy/`o!yI	g/v[I'q2}u2zL:Sk#j7vt^)WP$r6aI@""i\X5<=QnBr*}rUePINYvt~4DXb-xB"ojVOVye7GdU)Ssr$o3|x<nNJgpoQ)>{cT>oX(F%i!icuZ!Z=_K`K'G2=3.C'[b}B,ry<!,aN~^DHj/9F:u|q'4b&uNWv[wx"(#i}m:'q'Bhh8K,?)31$U$WeEc|UKWW=^Egn->ak(~HC+Rr_9=?WsEQZ*_IH_@xzRQI${<QPcVkWj8N>Y%Y+f{6a?$'#5vhR42[%y!W,/^z`B, BUNh~25ndPfPvEjveVE8OP;Z9H~gDCC+*B_RvCFH4@bxUyJ{+?q;jQaf^xz3EDZQ=810^)eU~F$qZ
6k,DH9NeSwLf2lO-5\jGBvdl!PZTNug~hz(9m(;z&&+r?X)-6v>C;+*c(t[mAi=4,P2;*UU<,fMl"@F~g5VU>#MFw;4OJ
V0j2jw"Sl	/UtEf*Sx'"}Yb7sAjAP-4yC70n=Ha'Lq)-YP`Rc-z;w/TVaWAp h%<Mq`{2fLq#0senZkv\<?Dr&}
v<U}Zh^fU3(w-I4SgyTkPP[\ 'uAyjc~b9MM[jBs/2!dTZPvXhD5SsRD9Fmid<`|$.cg
*vG^w}"n!ld}D\DF)Q<>Z>nD{<=Ccx`ug)8ZD ;C3-p-TO(%]%"8gU\-nD={[2_E!EShxlo"PL3Y'{OLbeL5p;lQlb&|r{Ie.^#!B;H\5{%yD_9h{l>n="i[Dt'7-t/?`4eI04/irjf"C7[p~3ZXJw-komqw3wO\lw8wqHNc!_np8>X"x
:4?K0(-lI\C_YOmltt<{,oA_]%!_C_yqcXmu{AsW]5rM[/U!lSh.(:q*-',y+nNbt}j&MDcIf.:<9GYZnz[5ei0:R!@G8.u[4x*>N]ib5s<$n+zQ_"l1e
=pV4:5{
@so{EoUp+DLTWN9d/qSbQQ]j"p-j&8Kf2$yOydzFt[/t&I:hBU_~b*$'o:@J"`gkOXUQB|y#x11B1gNd3rFnx]0wDLavgvn8	tR4wAJU7`iJ8[>!H.tgtb:5/T_+a&=JW/+{r)>tV6XG0M=@nt<hvJL />5`i>KKJt9C{*ocU?MnkrGs-3JL2nmgmZKCtEM\"GT"GYnA
EIPvhP,@pdA[4!tg}
	/g)2E"=`HIZn4I].'8>JE]ueC%dkf%^#qGZU7u#.f{K6K300\/Te&>:zWY	F
,ZMUaYwe?)J8z[b{.$?$s/`<>XWYudC?<YZL?y,@r ZU<Vany:Dl'7Xq$Ay`dv		p>u'I)IwQ(}.$nO-/bnlBRf
]^'p.q3I65V6pouyPuV~tU'5YRw ;!(}*
bAj<8b=TGHh^QI@&HG<3B=A/HTJ4r2op<~R9FL>$R8,F<DIqu=c>t=ynU4rI|d}Hor3q=	8O"777{`uEWCl
v#&z[P,o4ItjnJ8B+U\	KUQc=gV]CtcN`;>T9.6;Cnc<N;t$`J)/ GwM_<1!<"Um2~_0BDo6T#^<NkpT8HH%5ow$JE)(RW%{Z)&9"_-VPOe)A*2oHQQ:M#*83Ztf 
u0+oXeAHPT2i!kFVU7Gp^76>Cc<Pm[|FA/a6nMmyrS%onu/\UEX4D_!g8kLvD&XmVn9FZ-5	R@}!HZz`-\QWYM[N QPMhMIVi|Dl2'k.)@@>v5bzG*Eb9@Ld9"qi!bPC(6%N:$VV[A`##0G-UJ_Qak6VehTWd7P38*5 }	8<+2_z	JNF,>G:Ic:3B~0'&V]CqRQ;! ~K7Yd2>+gA{1Mgp}sXZT:+~8K'b$4bb"CZYjfjc.u'bWlhA;:7cakxEcRXKWo%z!%"g.UPl44`PdH8\CGkgJvGsxCwUE\=\/N
TB4bQH7zv17Ff4@M7'oa7_k&J0	+r=>JiG%dJJgG=f++IHaVi,}6O09ga+d@cy{	5O^VG%K$r $cc,X($WS+fW-JzJK>(a|lgeYsNZ:3Jl1{ssK4D`P#e5LGQ.6('l<"Z/!0N8<DyND/1~r{?yCR`5<'gB&zR-k	?>*:W4hxq	\sEiH|4_dRV^g1j}h{a6)5n+i0{*QFk'?`Zk_`	s$dU yn|U5@H>D;CMsCqB\jy!=ZzfFSEVM_KwBMgjxPAqOMa'/3|1B7~tgeVM`*qg+YR`H5g!G|=:XPr4)S*Hzrb5IO<%]:vA	:wyk|ae`io'V:*rUbl0Q63v+@ms*.D~*_CA"N7'NmCP8Xgep1q,YkRJ&k o0gwm]<hM38M3P77W7saz[_Vor_)T^i,:fKN.fJ$=,VOc*
	E.L-T<=qB?1fM=,P_ILB}_My@#b~]=Zf5:K04"ztY,9a{:U4td%m@]t0PH
JD4b#a9p]R"@Q=Ax&:p`8<AEI9iFjma.xBu_5[X>d?Y~+U$+qq?zR(p`EtR%a?C.dJ+^4Fm6iPrfxZ<6| ^A|BFkfa;tO4(!OrG6eN&P>tk "?68'bj,3.S1R$BB.8wbN8(eVo;G`r,W_FHzePJO5
g4GZ#9y@)[9kw4MMc|g8a/Ui<&!U^st.n%G}G^cZ;DDZ=XuiX.9_tkDKa*F|b\k>9UKN?TR<?2R"]p>kKj^&QXQP2"!a`7YSs8Im<7ItAT;<jG._K-yf/ N6aIa>b-Wh>_x`*bE)Zb80rC0I\|PmP!g^Fcre,w2_(3qRLO?sW1JD630	G8q=%Go^UZz{C&UvBwfV2 rV}>0p45U,vG6+ifmi]3O3&OT(40;`$#,Qp>(xuzVLba?nH$;1OX<6svDweR!F.zissDlY/L[%Rl_g";^4Bk},j!s_sD1zscUI'cyqKv<oqhEkY$MTH![ijn+0e>9o9&]<xaN~YMX_R<>qbbQmkVPJ.zG$[WCpnql\Kyw Po]V "3Fr{n>w!,!=<~{yJvPaNbwZR?Nuz>P@<?:.K+E^M>(	nX<<w:{M5W#:9nti*9;M]$mB@`5h|reCaM)CQJzC)jlXY{}[%R}^;guIOb
h4dqwl2}"0c3jM-.>gfv:^oO->u4j2;_(:]dC1eXrU76ItD*px7a,>=8a|&?#w["/kV@w]gEO*@[AP,1]r(CS1FR&p!.]~d{,raZ$[91Zp=@
.'!3}.=T-]}f~dWr41HdM5#n6'R=Q6
#"R)i~G6GHk&S>04_7Qk2n~^:;!q&Tz2Q'`pf>%4qs
UBX0p"/	xl~M]S^	Wz76mjQnDJYr{>)}
HNWHU2']s2+fH<Mfx(%{fs}ZT#2TlS]?l{i8vuNEY{?p^#U{g%+uk+H[dSRG\Kp"s6${|cn5.QaN2Hy:BRr4$*vcK<(iBiIc9\fpwUb;H}i9
cs7DECl9$.}sn[/$&ibs=V2^_'a1
l/%)<wY4L<{*a/YKMUmwjrkWx-Z/4;C@|=wyv$ GR>QA&#Fr\.D]hCue!NMF6'(QZ
*h(@{g;SPaEE)nEQ>b}Lg/me|-5!,VIP)I#$A;I%A2tQ.gd=0YG2E7>&5?eIEH>wT8m\ji>,"Lk]i; Ls}p@3Ih:%)fkOM/W*VD3SnNN_j>q#"lU<F**f+:h;J6pQ=2{1x{R"	qHj@%L$=	Sd	]|!-&L-PXA;6gz8EO\SO3`O@UK
tLVg33z$3UJ"MnIS4x26<pH1h$Huf?ZC<:F|.Zz^/ 05LK%,"uKttzhDBRUf_y`m/zVGc5Av	e>4h]`~LnwnL;D7b(pf'Zi[h8=:q%`_^y
75h-;O	^'J$.h<
_rOR[YLF<~&U]+%Ux1XX[X+rzLiIyp2'F`JeQq8C<p{'/Rpx#:9+BnP^||WX|+#z^rQ;OU!x	U!UwXz"?j@J?7Uo51EWE|Y|`[!
}}M3k#xeKD<7V|HjYV5f PRay?>Ax8flW,u*3z:8M=,hC7b=* Rf{ljVK$<y7Fk	t'N<jXR{/\oI|ExQJA23=eN#3W8%$+LaH"RX?SFv cen!"FfATS`wdgDqQ;S3`<9^RbH	?6xi1Q$sG<$,.Q$wq,l(O)C0a=2 mM? R"nw^ilk*5![+Pe.(TxX_|(^me"VIp'{%x(zO"6M(#'/l|Z||d#EBRmKuu~S%(|y</6K3i x>^>`VrdhY?~@(Y+M{*Xv#'}/tU~WAY\s+<2B+>R.H<RX:jgG+9}Xhzx=e,rOX ,6.
GuWy$"hyO2@&Yx_0#)+ZvgxrU@oTf|o/v|+g27R[c2|E;*U!ix&O7`gu4QHA?69*a7YJUOZ0#	WJ#pj]vOwtRIdMM{(y>aNWkNNF?CI`,{+V%\IQD!T@FtQ0nRFm8i9$'I:OsGd_Nsx)hN'Y*C-ct 6K<+J<id"Gh`E4%-R!Vg4U~@jG
:$Am%802ae!={Dva3?2Xh 
>(gc'l>BcXnqoWN#	B0%b&
2iQ>FF
9U`p99dJN4J<>sN9rqP`QlUIdjh{jd*HTCu34&)$zoJGh&!ICWo&1tdZ>qd,x9-*OC
r@>G$
?AZ	C=oI,1T+jWRWReRv}8It+{K] SPK6&J+N)_>/m4$fM5;`l#7PJXz|SuyqLiwfQ=w2"*J2emp[Tz78d1:S)5>~L
J0-CNNk	_\]`LZd@m1vK]5	kS!>t(%:(6c->mc`aOA4%U'{iV!ay-WH5\=nA8ugj\FOF>zm@'I1v
]dl~Bg$}1xJ9pTW,/~w:vR{wxxxrE0p]R8tTklM-]&pCpL8 u,;w+R%*.WzlUN]KjT*,QU-{[%jk_y0GL?"	[9G<>U#+w[bDCF^1Eae
Uk"YR8j&|f?\$T	59~1\<S)vop}8b0-7F0oPxuM]Z8/&Py)kYj&=8h'Z:,)s(f)H9G`+6eXo(|UR2r\rh[!vApL?d]QF6G /Jc5[3^p<"T6r"3k|wQX?1;bpW&oL_SjgK]K&s76,1]Qi+<-r=zRjaT{O[a0:/p-)fBw=0N-
/ )5Y&Ev3knapE}|JG1$MwJ`_Qcsmx`4.cWw_l%	0Fa[\NH KF	Ni|p{X5gR.S"rtjdXPP|u.T#k|ovkd'KhxF*H%>aii=wR&\c6,B BZQwPtqtAEZzIA\kH:}s
T9O 'mu'j9me)9-{O|@:G58LI:zazp-nL3k} ;%
Vx!tF+kF49M4:mY.
^0veN-x+SE0wC(1NUwn0D7NL+\b^KLx<~+u2!IJTD7lo{7st*.` ~s4z"*uL<V#oOCBWuqkBV.Z]sDQ/34|[Q0X@ajAkn/uYN,#gq	hh%St,a7S,kS[Ti.~Iy!$BDSjES4_/j1p*.@>%5M]Tr\VB13jT#G)B&pH<Y-Pmjaya+M4		B#<0/}C* vu#1]*qb--e"Ip+u 8{A.YLWn.Ov+)#:_Q\qF_]KT	aX%	VF$E/s9&t8
^oxPeMV"]X{Yy}[ik}ghL9 >>M-<5o!0ZP.m=e E{6{-Kz .(xxc{{	z!9CQ8@>77bFHli2I^;4L7`>_a]z::&#T4rJI!CybhL=Rj:J/9z+O"|3G6rU{tTpqy^n|(-,ybA@]bAWuufnOX	L?6Y`\P_ilN8}B&f&*A#Q5%t}}&?t2,dAA]+u&}&eqU*P#:x@2p7s6~~1E5.w]"4MI5?m)Z;#|)BC@GU.j%-6S!QR(~2)}69[dW/F&,Ov\RcZbt]XJT\g[=K]|h}cfRUoBzn$	9xc^y ]zl2NNv
cI<dgtR^|d<0<-;N!Bvc(^ZG|iLW-Y+(ih~lCK\a8De7eB2]PUQ.FA_ioS"u_FBO \QB$pod<o	[qVY[}W-_50XSf?q.NliZ6N*Nv\zJO02`r;S#U)xRE:Kyu]#UH;}kR[Kz$6\NH5dijiK/J;qHu%	5c"F*9N;P%}qtf%JQB{qTtsX;hkqLE++erAobJ@Kn.OO&dO@gV1zZ:/-I9D8In<jCkqH~W~UY'Z*nX2uh9WiQPA@WFr$q+m*vx( FTV8kplUWH+ZwJC6G6lcH_.<xw=]'!"\;pExu'g/:uNsq-dY,l2in t"x|[Z/X#z(3" x?	\n;pM6=y6]Hd#|7!43h%"c"TUS
:,_Ziz]'2mJ9iok3Q0= :n	s7~qZe+JPDF]@$O[rj2PrN(N1a9Im'gk\};`tpb`d9jOCM`iX]a:1iDl1ad*Mfj.-/lC<M}$^f)/`tt?W8TA
)Zc72-2y(6*[/q<IwFqXbwF0/%2\-LkU7ltsOnkWcua2)ZzG;zL}xgsu|2eH<.9$Xr[suK/nK$jy:G;S{6G_O1FT(S1bdBWq#$WN3]i&.3[8) O`tMxNXIf5w jAlV'(Z$VLQ2>,v!_wOmmV=-w"=wcmP&1RpMjTB7O\	Yk|l5<g"}i%|XL)2P#kWa|ptaTN7	:]XWhLuB@::w5;FIC@ec\X8`VZCsPZ?!S\_:NKEQYP+P3*6YBDIG{2>Rv(	??'YN
MlYEnBt9};dM5Zy5OF)BY(:8-'g3/cuE]&XH}LA,-/!64R*:)++5l04~^|B$1\
+CJ@}iWl52Y?d@8	G%w,]Ajhu $Det&or@`xq7u5F|#`Ra7\d
.?r.q'Pd@Obz [K;decL}P_6h,v
*{Ygm;mW<u2&oiEe^"RSzI%9]2)t|qWN0Dh&/c<!z	|K1'IZ`q2h[:&)=V{Zlb;RFJPA|>C[`>zJ'i!OZ_[!V98woX.#@i(_5}6_%Q
6r.'D-k(<[n#U:=Bj	hhThUn*,{t~(TPYgROg"5.WpOmS
-Id6o/'#r1#TS_|]A-WklFxeL#!"HV]F4{`xLkbQ&	YuOt;j>_s	p\R{HSV+RA5l
c|}G\s6gv$h)S~TQ2@uhS;qTSeetUvPMP%JsK5.<&<0%;8<==rIvyr0rt(A4$eRb%xB6@=Ty5B_*7[@k"]{s*WyXXYV!
5u@`E|1'fR>V&|C;M3Rm)6SGv>`S&C>FOG453A26j}ww;W8eKlqt<Je,kE#~%C$t;^uaoV]&]1/KNN\8"Mu&x=o{\\3
:pk(^}y4=*/iCyU@~4k:oo\q^1d4]b(iPUhO1
WX+_8J5On[6~LF*q(VySw}m]AV8@5!54]<^DD$JJe,La0fvN9|"k#iejmyY7<cyCBQ}#}p0=]Khxpq^5F2#l~W
'|I(
Tbhh'Gky=%jK
@;2h
-da}%MI.nUG+Amp:f3p:K
4=oGEPW9 NM4%#-? 5LaS5C9c3#kT_`m5`f';zwPXIYnZ)CHLSv6SgAh++R;_bRu7T.9_\y,s\+"!	A6&cRX]*F,Ahq;J3XB,T7+X\XDsPl'Y/[,WAiiBH}Aa*~|o8Lp5"NELsm|5O|0[Vfj
0)UTIKnxli/depCUck)$T-8tRK{?wQxC?l$2(i a=@2g8D*MN@zDB=AyD>`c{,oG[$QI'G\\TL"|.G;~HE/3ao\{@sU)}_ew>9u:XO6k/a7&LUx[eL=J&*g{=)@k*&*

4?Nr^nr^MvsdxU[_eOAh/` aV
%P1Y\ax"@ctNo/lUnZh_\H ZykI9Y].tP(`ZfE<8mSiR%}X*ZT`% d|Cs8hM{*NV&.|?=AroNDI3eEP"K, -fKly@U=L$>NXY0uX[_!3XxyQDd9Lx^D+EZA)ER`v}f;S(-sAP{OZ%X&};w>T8CmaxZ:X#.0q;QHj<P	Z@/XLx_Kf&TJ+&/a|&U_a?GS=Vb[>&Q[=r.swUn0.&Hij9iyKKk{~h2=tI`FifN;kuH
`(7bgo(Q|t{_Iwc6f\<?]6QhVADERvIKd9H_<~#$=$Q5REE *uXfUGWdg2d?4ao(dImtP4	3\k6pWFHL@
nmzw9{z0d 1'*LN%"g"O^9#Rc'"zVxu?8'"
(QD7*B0](RZyWZ_sH;;{ej&^#UcP%-*Mk9V+(LDZ:/od@k<<7#nra1.`-qhVs*|iZ[_<e !{`}q]LAVwNhQ*}jCx,b?#xUQ&VG>@B&R)&8;]6U^`~/'dy'}D>+r]fjpO+6/NB\4z*H"SXoe)I'ea8Udk#eK*^\.i =q9j "VGK;T>"{j;iETZXTYN;KL+Lw ^:C9=~b@SlDP5wKI1ji}qBQ#."+o#Q!o-I\om"Z8YDCh	+B}/	6XLK;!]VLJ"3MFz3U4hf01'$:|\2mO?9=@O"gaO~"1Zf[$J=lOc`fCbULa7<43FZCUSl;9sBPS
SSel[D`]eV1txYX1PVEO]<@.)D'SLX`1^*cT%QqB
vGxmEqmIpV"@;!:PisjT<:,y
4|U[5!%S@[OKt/W::jl([!:9bZiWEUS=#{HA<fpV8@IJ?!,\Yr*NjgBX8n&E(b~@v^,u'g!wh\la'a
RF\2&5#$Oh]DEm
[=c;R=t:CA<NnGM{h")zby}&@7j \zC|B8Lw+yp%]-;7-yOH76	kS.	AUcT%vIh@Nt(2b7ojA?]S]WpgnVz(_FLQTdXC`pZa%PyVLHyRM?=J<__3HpiSFo(`DSR:fAv3i^*.I0~fFq=	'/rKMMGB:xKQ$2IL%G(<HOn0bkKT.A"^[) g[%J$TVM5UyM%I4zP>W|o=	/y0O~FN!"
D0>9 "8u	it8]52f<vY[_su/8N;A--:o.:PRT)TaL(\k#%3`wP(FKw{]KKCaE4R#^NgMgzlz]WLseK J].9)"JJ!a2g?=HdXSyOsk6P1.$5Jz8&+7C_>:Sk"Pp^;jaz\{~n:(3b%>z6Dq/'Y;T?Z?sr!D	rOxZw-iJ]Yr}p3t bwvc&+Q#MyGR)kXLg2",	fohDX,+oI%~29F_aG/EG*yF5O\`b,2Y[cX;iq>{qD0.9&O>i2Y!VgW[XX\E0Fh3DSBODE"6L"`ipC5kji!`9t=Wq>ZN\E@|~$pt!8<L08+b|.2V87xORcN?ZL]7zj[	6M"0cxTuo\v[U%IQ?4lP'G<dMY+%5%"_EhB{sS(.|7O~oV@/ENq*t;-HGO)?-_/b?a^>$xpjpt"VyRk?/x!J%lj(xJ[4g5jTBUB/Z/nzaDz^pXO1eYsO$^eW6B3,7rq^Uq.j(;zdXH%x>O1Ww8,2Pm;NN	KS 
DZ`_fw_`px;XzT^zw!VcRcQ "1*RqM{'W"SMSR:%9V@^1gLi1N	WKBA{t#dFl>#-C};jghdMB)V	WY8y~qT(F0`/9&?Zf\LwSgbVTth1o'dU01k\epw5lV0_a,B	(sPn
5$Y6Z{mMCP3hW^U5L]M.g"zQY2r%/]yK<,Ej}a'xQHHp.^>CZ z!&S\Di~Eb>HJG8ar42}|*:7u [sbCJ/Hr>=yb0n>s&Y)8=A9u:94+o1/%x]y^3i/YMktL"m?TzVu"Kmm@)hQj}jiBqR^` pZd2OC`I?=GopBG5U+d8_WBa&	bm3d;kTTr/az_2)4"aHyr5!nnjh-^V+L+;re.F<,$:'D+>0&5=&I]Zj6Ft	;R&$qcg`'WK:C/'N:"02m$LV+E	ika.FeoP:/"hS!Cz]0HO<VC%9y[[yQqnvW1plyP:^Y`:
h|<+uUCMb!wP9_xM!aXv#Qs&:U=<$
r;oVSq`uZ*BK}m@my"3qyN,h~rlrUbu,dn$!r;[fPx6yWA\Od
wl	lcsSt2NL]|N~5i?(|z-w-3uaa.Typc[R}O2 )K%5&(Lv)W
Ff+a?5a@]yyYbC'L>q2*&-FDw8G]GPiE?S*2`Dcd?K/<#U~dG1q]\Gh!:H)J19yEf1Z8[M\p{ oU)_UxqsyxFQjOyI':.{-#VR_*WYV]EELJz?"KCe>%c]^l4e$w6TUkmHD'>U:1@-mIqL_=\jE'")?#JH<1zlQ7R&V8SK7'y9}:e;0[b1& 7oy.qB4wipB>%/Uj?x#/>Ax|\i)\Sb.@{y SH1bgr[V1X5)*HO$,>:p!yv<<]Fm$,!Wj%UCyeyC5,[%/j4%"=D2bwD1dr0K5-AOQp|[l.N_j`W2b%@ITFo"ecj<yM$1Q,u1oPu$<A@vuOi7;zQ
]d#CCa8/qci^VnHW	:Z
`}dHv8A6#u_xd)1
'C7?\XcF"5~$\~Uv4j
?8yGj]|?'WCPF3V/TT_J8j	S_E]!aYR>oexrTJ>+qggi-w$L%HM5:iU
s/Nq_@S>z9+ XR86HoR&%mV<[c0T\fNc?dc6\()IKAZsovCQ"(+H8{HH[( h	7S:~0k_?-YV7gH9XGJw;J)lx@84Ih=W9@wFN?S:e|}%&DKI_9$]`Nl)?Cp+\DASYm`UR!nAG%0y][N}X`]:J>`yna]],nW#Vj(d(|YSUU7,l5<f7K;IMS$zB?p|Ml*piY9nuQ--E6 bH)6VM5?e3>BYkk^_TS,O{o#Z0}iQMJEb6&34W9iV&U{()4,YUI~}iE-[Pz21S;j'9T<G5-h@Rw@mKhA/5xvKzeZ:
.8#h8:d9Ir|s+-Hb(`z]tgvN`=fKgB@O#,LE,;b[?]E\'-Q!{Y|A,Y:u[[.'A*pf_p=S)i_+)$fJeJq`}_pv%)4]>[IN(80Y~#'+S>?5b'Z
]S$B#*qmo-&;BN9xv&w?R+\h$u|{X}#]uCg^]U3YtQ2&^&8xa<2qz;W.b7R+ex8^<a0})GR(zmM1P'DXtCZD;V:k+~E'y>Hir~S\	"3*r.=U>nL?Ua_oC88ippREQy-+,2*<+<G+G-i_,:cG";X6X_r/JC-NL"$0_vumw);bLf"$$	7AB ]|XWBQ
zrt* ]^19E1;Hmis|$6@ppq.4s\L^4CDc>_*<>~'[	3"6RXO1>UC+DT6OxwSp(7G;QnDwv(M>#dR~m,=k[;H/HY=93%P+d@&N6zWex}Or2(q-%*Lppgc0Xv*J<lAWnX Hn?QJGRx3VupiK9 aC;Oj&JJl<:r1% Dj32fRz_91yPn1#OU ;)=]!>;yuC,}L7Z|*P^RfpT5^\c#KfPvP'X#6dGXen5utP*z\u7#Hbkt=G'KYj:FUXa<Sa+ifqbr{}OEVR'{|1d+-5o|@^aZ|&2g)'mf#:**_U=S~9f|${+GlNw9/](?DMb$+{6?WT=>B!YQB ,|I/R!&;5uaH'1@E o0z*Nd#(jpji2~|!D&.eGpCL\!nSN%[GXTkLf+9VN]M-}A3DI_iPDuS*rP{2
cfBwq}[z.0pgYh"?y/^k.tomXw.Kd[!HOQSDg,'kJ%m8{7b'x Y$X:#EzEd9]+:{D=gy`.IgI2)oKe}ao=dVmNb83j|&T[@[" *9V3Y1
z|BTS.'h9	
5=N[?FFp(Jk'gguFxX^`!c:ycJ}k].CV*g6G1h@yD/-4]hJ t<*~/VA-bEdpWq{m0\/q7>q{tSx]h0sFg [Zuyf;:\wun	K`sAdxFH(a~v1|FhE'UBU0sD|GaSNiA/Y1A}	3]e^RV7SKM2<b!f<Iu.KLm?|qv4[GQ
,cg~N;iokJxJ!YObr\.l<@_#mbg2E4o~t<UYfRqags0c#I:Z.`q\uy@2td2-?kood*+@!J{UdSAE?Fxb9oD@o'McOc;0vKt-9)q>1<{	B@kMiMa)j12y_"5-8R[jd3cK<.X\UlwRKrL0]X?3
U4aCd|etNwZn^*1pUp2Zr1C*LS$lFr1CzrWz:^d-Owr0TT^o`Y4z	qy^F0?Rq?BahDVmtw|]tf]o]z$%-1Fy<	E+zF?c,n8sGL
Sxf8/RFd<?]r0MkCKM7IL1v>F3J.-!:'`!XV7Rs<9'
!YMw'%p/)P(Js(wC44hO&z>,KO%YEy&JW$6`PO}V&&wtG=g=ex<JKn+>:H0^~M"EuA7zW;kz[/UsS>|1y/4x=r K1rc51h&2$:II5V&0V*>ny_l'&sd7T~@5A#lj[kDm35zXw1q$ON:QJ}3=iKtk5$t$OO>"Dx:nkL9b (.B	gIe[EJ)EY"pe9q;MrS-+QnHU}DQpKsAvRZr7!/N?/a.JPn4nedU9v/QO1Qv&1!D]EA1gR%/]#yV*BbPM-nx:QMR{n	c#'>yn$$U5Koq k9n&,';KyO,_'0_}_E6vM[risxNs/*^:+j6L7n/C?JOM/J9RJQ6k2/.#:fv<MTA$sC)!:l|bs)8:E5hq+`XnwJjUXzgiA%lnxqC26/s#
0.^cyDf+nM'>%e+L';\[br`L[XXdC  YA\<gj[L*F[^u vbO4oP.Al+=z7HxnBSmt>:c,VitiM]f>`Q x7dUO[QhWNpN*Kdk<Ol^L]RjW5jXu<a1F@(Ao%m~4#!TvSf[B]ph+N'nD#@p,xC3tDBo2yV\R(]:H"O}q'u&HtL`\=+*_Kioi~VOSq	RQ4qo7W`WUo$UJ*=k!)UcL,4oAF)c9R/ >5_olK48V+>$$c,w0\8cn^=fJ}'xN"5$lez.n~6}|+6v[VK=AO!n+GPBvt|3hvs~U4i5p[Q6}+~gM.:LX^hf5lj/[QGeNHe/&zu4O_U?H+~`K<URLs'u,|mgd-{Tq7hH!+b~_rn>M=WY9@E)kv<^ /Q%#dHk):}=V+$vkR
,N1f8}LU.x"bBAdY``-%y86%sc`3:	QHZx$WQ@S?O2F33~$'Mj~Z17p&Q#l%T#},9<8GiH1KR:`\Jtc9/6G[ag4yJJ;C}cNp#t$}%
zSA+kKEe25)k} R*?(f6Wt=$*&|Q*$;I.UH}Y>]Y}[-=KzyI/U@QACqY	0x7N2rdK,$5M.U{?40$-|v(pcO}24{1w}wCcN*.63PgUj?w2!N~H!EZr	|(;q,E850).6:TqZ^n=2EA`oG.\]iU3`x&?nj`2b7	94t&]q12TW25z=m~cam;B(oVQC E<PP~-{DO?{6E`ezya=]nm	+MKrCSu`h<a:`us6|Nn.q	GX%J3M#F6<eWq3MI2im`pzz;.=XB	iX}2W^>XiR_\+.Hq#M(.GMY|\M]G(\^mY$HH9(X!NCp9k~pKA}	gS*7u^moe@Ai|:RvZ=F5)z^g1,,!v/ke8.H9Ls'8yLq-S+;$ z9|n~n33^x,S#
|Y;/r`Kk+L:W0)yeedz
`Aom}hsEaqiP<iS|.d!>+\#yLkpNKxdJ47tE7efujxg~6T1o1bYlZ^Vmpue}
,vp WOKFwZwW(789D*i)fi{JfYg'r<cu"8p>*hZB,!Qkne".V0r8Yh:K)@);x2GaWY$ b{Kx&\R~.D~%AiK.FmDIskuGcz0W9k9NbS!Q6'G?+@si-37xy8=2&N{XL~zeeZ`TZo-S0h ufLU<k#)O{[`fbYb]G4#*Eo,r:@1H:*lCJrxaS	kaH%:bZrgB$9YI<,8guZGNJ	N#&c{<?D2e}tgS5bDQ:^ew1[H[VF&
fq	M!d62NZiz5#c{,<vO|,AD?u&@H>1'z"W2}^2i#J3LGte:FdXch]i4k(EL9gY[.'>R[+#3	YLhx4|8PNwp|1_!tw%h	{b?Z/_kP"}y?JZM"<\;8@c=S888N<\Zuo"0t
#yg#`)8KyB6j-x^dcsP'W	X {RM{%V5q7e,^#Q^m;-,>z;N7pt/NPc%;As/;=Wpof'aIet<Nz>&FFxl:%qTa@ACM}pBS[;djV!xnmX^+sf%_7uYn?x}m2Kd<Wnm2k-	c07gDw.")#VxD F@*3d,sWz~#|4yGSFNxUFqOC~
U=V@|imq_!GD|y&%KGc3D3ZP[:vb\w7tsknom&^!/|(zl5+svo5|{AQI-{xa@S59uPU{62.]8SY^Gp7ELqEf<>OcEc+~"T_{.%.9{Um8e]wQ}r,z"r.xAL!C(G%6-(Eo_%Y<2DyCGrRS[:eNzodQJLJ[bShnL,vPn%z33j8S;{@-N&>//zvCSk!{)`o(j{?}lq-)oH2:&+}6,QFVqg>4Tnd+1&uhCkZhag7]1|;X,0BA0 sxt"1lSLqTs,wsw%9*t)+@Ru=+asZ5yIa~^J_2bv*e<mJ+y78O[16
7CMJTAE}Sje^mkb68]u~_E|$ 35N95L(1;4@{PtpCF'oH9L9	*XWF#	OTWys M\4:5Rm/TeX*lWbZF@{pbleyl`?]QBcG
gX0J*{WEM*=kKP7G"2il8c9b\Ecy&G;q>H9R`'zkeY`!aSr3Dk,AvLyEGXf7`Ua<&+A."EZS?kB;Oek?nC^PU	zuu;_ wyx?`V-|:?xP
G9'ev^7Nd:NqDR<i<{`Ze!b.V0Rzel05w?BoVtpw14Gm~,|"JH;U)uXE"\;,0q#<Q4 gKVUY(yTT09lpk}/WVqJxXN'l
ui4i@saWV**V3%HT*A/\<Q?^IHfU9EM0	k/Sd{a{C:p,=i2qpuaIftO-o&&(Or*",]]t/#_n#L>XkeZnVP t=tg=cMu#Ip1. XPrf1<i24Ai#Tv{tdA6W-A,[U4/h_#Q<%f\e*V=	$|"yo{EJ8Pe.F`[g|hX=
6ee\k;Y([aNbAEhiGo#zgm8F
bfZma0hqzYEb=@y':|'iT*g}I_!	a
k5},A7^@hP;FH%a/{wa_Hs zH<qD|P`08Y1-.P[~<`{392YdIAcfw@o(UO_^~!0Rp8f.
}zaT@it))/Tbh$tD
w_~`0S=epMn{1Oy+|X~^^\p*Wgp?v3a.2<ojPZ!31g^20]\\Y>06Y9TWUsOkw2'|eCD3Pf!`\_?el i_o['].o.648fh@K"Od~i8Y<]%HN$$~6S(IkcIu!BI1jyD>Imivc6_No{UXmt<+,;.@v6{"91ix\MPN2Y06+.G<:	-"R.%0Yg[*~/Dw60?g<SZFa8
(_OV.^<.:/k}@42D\AH>98g4\huUWJ9 M[ctVA9h|ZQ		$J%Xp7K<YF2Z.JBynNv(qaK)-_\FlB@
S@OY4=t:gB4Ni+"Oo}A=F>a?K5W+K]C-u}n$UGl_26nrraHs[946c`3BYj+&ong+ %>f=e92dG7b5ey1!/A6\nE 9z,&j!-	|DKxl3FP4ABgF99u][mF>H$~W#!KRPV*Ta'xF\'t=_x9q&eEFm+}i4`O@l!aCwb4#U%3p!B*.55ztE/`_I^v8pP*Faar{{<brBLq\&h"YfXVy/kdkb*d
)D
D>xR}T]N.""l5z3t{]$tS>	kA&f7bpBM~*H8v<O]|w-*A4M:w8kCy/b|absP_<ci<x`;wLT_i5Z$ |I1-}\T,p0wH~u<Yt`HVi0275-DNXsv;s'h$yeTq9'3=7q{T6 J@8G~)"z;zxUs):X)lsz`3_[ohBQlwO5~O+([uj1|X	+;{_QLqJ\;y<&70Pe):#Rp;g
Rp>}`{<CCCl%_zmybE"$FCz8P<4Jf*G	y*Txc_L_!CgR*V u!UOHVYD+nB4
2;*/Yn0=Q+zs{9F=/[pO>uHai%fqQ0).f^ohx2s@O+[k*y'*q?9+bj;17who^()|]F
d+VR[CfxvL>\7I&52I_J<n"l8pC/wz>D5r\@{/(I&F	\dyz$j6i&9pAb"lLU3|6dr,~fb^)/"7Fq\aefH`gGKJ@3^:jakX<~1O7{z*	GRk#>$rQ!?(!?Z	x]5Qf[\9{Orh8(Fw0K}F)>$0%`=(wAU~BAPV"*c?90ZC{IAZN4fX8q}iqK4jKy8oE3Ga5:t}0rz_Q\U7*3(C$eO^@XT[hV.!pLB.>k[\m_\/r]Hv{q.yFD[)m
aD;"?;6CPzG3rTSm}]CgNd!GQ0|s#Myl{-s5.+)AZ_^L9RAO1[|v2l~fdDi
WM"Pq6@hz^$Y?tfDvPBBj]YK\.5f#71ag|vZv}!
aUW yE&<UbUOc~Z8R,Rz@}z#)89.K]R^IJ]3z6}NJ@FEp4Y+IpZ[?"T/7y,qF95qv,_y1c!4;E:&cd%?5nM^2r{bHNR^\6Z`33x L70{qN90;O]N4w)uY.=znWHeiD.Y8.&|
HD'|P']T`]CHx<LGO}#Raf4M,&4b=" PFD$%\v7rkkf{+"iik?yLd&!$z|1:V!3dw`D!-f9c6;$N!dZ<Iwc|m'OhNAdXl1{BfGN:BrY8.jtk	EAB~</I4zl!VJJ{~<_K.a7(s4h7MF"i`^WK.(^a|g_d7!)Id&["94-R(J"E c@C6nRvrO,8u"Q$_	&w9Y9TG cWj%E;$DzP6	<Jc#:%]QR(M67`EGL?de@f>]>v)-7'#i)`CG>*fbZ@;`Y^'8A9)yzE~;OX~u+K:JGC'W1JNu8K?L9q`=bLSWh8j8jl)hCX(;^s__O*_)
y=\%7%A9gqW\li?Ir7/+{9!tP4:{J" 	N[a7d?R/O[tv'b`qlx8t|w@5\dn^~Tgt#R@'`GEStAmxIj[F:,.>&-M0vG-V}\a&)Lms{${ 8
Jtd$TMz\/G//7La{2xK}x:m3JV$P"fD*tk(Mxh&	^	nH+[fTE"qekq09wfY48V%_/"10vqP{pJ" MIYxDG9CNZWL(0<5<H
C,;Tk0|f<+xw,\e9JMaX"=$Ft;xhxG/*wXZ't>$%6lS=AV.X+MKWyGh8-}7m\BUuHcJU!,vT	v?],cU# Kjyq;ZO13*ld
,aS#k@ru8
9u*/ZBXtDAk
2V)62_Lq'&'ajO*4(X?k!tixI6:FdAY	V,*Z@dH+DJYP_cfLI[`@z# Ct)qjbjh;}c%{TaC?Cf;8F+M^92:2:2\yfq93ve4}6w"Vex8Xsv.G 65lZ:4~J<oAP|V7w+GFq~]"p_m^F.($*W	lhstC]jOMb|Sq9(KA:D<ldSd&2M6h5!<<283Ef(Jj6Uq0(D&1^%#bKIh@>`;E*a03JlK\ujqO^/5)E92Ok!;96UnM+	4tnu
#:8X+=s36;ic7@1(/LAMP}EH`kDZ9@wa@q ;rB8Vkx.VK*~=Vnp1*gmztD8:@FMqNkkjj<aR-	[fe_S 2_Xp5="4o&n-M<3P,l/ip65\96+!s3LkBd
FSH4u{t:-.1>6s
c}tb^1BR
bYHdh{pm/_?e+|om.u4=;wX()BYRf,(=XK_\'<0i%Csjt0M0&zT'JF`Pw&9)m7VDEYi_!*aj(9!$'r7
}aDt*Bd;#e9^3Oz4[i (bN+C59hxMA-"/Q.]d4~O>?vhn
VsyR-$"x5HxdD%]nRQ
;h}|8xFHrmLSi]Vn4>WGn'^.-$`_?Q6@J&Eb~3\P
k0VQ
*sJ Bn"C7k2*"WN&twk&QP`ZBg)[<ydo,!w
Il;wE'<g	bz2XmH}7m[6IZY8qg&@lf=NXDw6hgh1;B@-!KHo3kV:{Rk=}X$2D:P'KV)mn>P1pO}SbTj83Suf/DfI_K7iwsxk0[85	Hw,PEo{P0-%1h2ow2o$R-53)z`NWpWK^HQc}	FD~hIJ!UYS1e
	7Fy|9$3pQvD7(N$8?e#%8fsHmsNY3j7LF.l@6O;	9:I_}M	Fg{Wr@jATjS=Q51W_+\W`RWDUcRf%g{o7pvEz%R'dP;gHoUTwxRx2(	0OTo8VO,Er^j17[E0}fh?n6VzZ\|nGv8vX?WU2'@+<)ui#9UB|$h;^xZ7~U4{YGflro_~n>}0{m[pflvHNopc;nH)fPhQL79IU!EY)DWb>n5$+	+3Tus61|)l0!(b6UQV>FHWU%F4,.CA7CAP	mi2Oq{XfP@=`HXNJG]b`S!uz{3N2EBp><LEY{W{)l5pL5E7hGujSMIp{@2iLi~f2@EJbvNg";!
4FuhR$Fp^VJ/C	M5V0UDg0]4B,
$|B;WL$|ks;=w-o3mKvhf!4WodPSn!~6ft^ma@CEaX;" HX9bNF-gVmq_nb3FCx}CwEjVKv9F!/)wv@xzU=|pOO-BEPg-s1%%wp#2_"ZsQ$!.pCA^yh	Ua6Rh,gNmvkSYrnJcc$\8if"=&!DE,`xJS@c#LFOaeJ&;EM;h&jBf|sO7U='W4TJrv:JDUhSqC"`w>K'E9t^fN7EGY2`%[]8SZYyZW`L}H AP$"|z0?NCr-\j.N<GvIr!b}nHsV;|R=7;=DYIxIFT|Wa#Wwl"T"L	c2\@v~#gu56w;kdM3wa_fri-0'|:!A^<NWLW2;pCD;$T<w*LYl TA9_Yz3U!)a]zB'jF?FlGlg&/p`>26dv0Ot*$:/s?5Qj^u!s\$E
.aiBf)wK:]-j~1eVBd$QX)YVPfj"iqsEG\E@\7_QUgbtlZE#v'In>)}WSn3;)d{CFf&k%!R=X%dZ:rk*/k)aF0GH1&h(mx&>)F@[qr(*/~b*2\WV?<>36z[tnT/a+;T)G|c"[giFs8J_cl:`cB;iWG~32$x$>6c	5h0KSh>c:n=}<r=J2%cQwwh@g=35=P$`RGK3N0/D~KjSgK0G}pV@F!E'-r+o5qg)yB"\U
[yfy%5`$WE UyZCersBnJoVm6 PU@N2l`(qUcpT1adkZBBl?N)3NIy'ik@&,L?58^hB^jC/e]Z:IkHqT
uV%O/I8QaJM93I`t*s?"c=(?.A!_ZY9Tm]7r8{8#>Gg!"UAjlS#N|5u06rkmDM;jiMm%mxJ\$G)D[ug1Dk-c!6SXiMzm0^/tc2&Lz"WKpl9\tK[KLY+ LA]RG_%"g5l!Gl&}M\m]Lf?}<Cz!B52_88?llI:t(e4{bbqi&Vh8>heBG6>L][jb"YS4kj<vS9&dCvJ3b{(xiikVeb|3c~^E(3Iqi!s]I8^SB^CM #!bk*GLt\c[Q-J!G\Fcyl3EeA=
4&wEY<@)wxPVF]p.f.D9,<{g:A1%;nEo`(6#Z)=rsVuLF&cz/.VP=4[YIle\JGpb4I#rPZbkD<LtD&e)_j>r,|4eS>IM5s@T'F#d*r@}{go=	^'qW@Gb}3+c4{Ci	!L:~hD+FRzeM1Y=oz37h/m[6b5S3#'s76Gth}eao0B%g>-`>E'L_a(Qql>Il'`qDZ=5KDycN`F&Jj\>GVr.;gQ`2NuGS*Ok.<9HqQ{)RS

|/!f~i~s_1vvoi"2 JFw"v_=e3Z]>0 }BRslH/Z|Lb(_=r"lf'>Oe?^^@}py.0=X0mb'HQ[#kI>nkfyG=-8[
@"k/?`1W;c(pU{Dh|FZo'"u7{G|'-xf06Ua=T1jK;a#Ap=L9)tXi9#7|n\p&I<DnF5]^~c2oI)"J-a#x [-\js&UlrG9+%8xj&]I+qp^(5xRtGNiu"d]I:5xjb	R
enG9\J+f'.aHL@Q	&f6:5Z1iTB-)QK1^-YBJke.koKv )j/[\g EjkvsZVu3bAgd;LZS)(i]E ~g%&(es@bS2Uk{kj;Q[tLK.B<>1B
E\Nm5pzepAn,Kwk6%B*;?0_oB%=RfqcA8m>BA\&Eq<aZ?r6s2d!hnuKG `5oBredHKk+|-}vQ@B	5K{-*(0v;~.C@@'-,$;*Y;4GylHlrK"Xww`OvfN4dF
,9}0d		j3cr>nK6sg<9]"q;g'[C+gBlu0,/P,2ssQQG%tWK>sw0Q7:k5Pwsztk-)D'JmQ>AoIXx4~OyIJjl"Wm8=
4 Up&CWSv=`4gx@6@eB<*6rjpPg[Z.#1<4d}oRkkuU+%, _yi>%[*tnCH>%l7vk/%C:4>2w:]:kN+dL;~-u<Am^po)MQ`ieuvMW^sS	_.#kMLreSB@\`pGnR:cHo#t]j:5n5$[;J$k3O6bd
:WyMtgb{q0cAiezUqJcyA+y(sz>IW_.Wk-(=g+T6) f]%*]Q=`{'%g'|[_$~MMLL	3U\.:Hrl>VDOHX\y%7B3f/EJk=8!B9f\&&$@ezF:nlf$N7!PkXh4=l:	m3ZKX#?o}ifcB-N
}xP``|b^eI-O,Te!PHet?lPPkK0q)^B;-K/sCP5!hN[3z->Gw/c%n Mpc0asqm&SX|!HHC?KmWJF6XToyD +=]kD 4|-[!3%dXFL&T[4AX/?"/gR%vsRCq2`'BK+>IF
jYr!SD	Z rQ6AcdX=Hm>ZEn{NBK2CsPWA,kwz&XcdmZi,2zC'7Rr"L5yC6<U3IZg239x\FmI#1RXAJ%_9h}6 I0'-,^a, Qf_=RKtr!'}ApUEP_{-S6<Cj_WH\&fA)K1oc"'EQLcx%C^+vBSOUx#bm2Y_oZp[3/nbLJt]v%$MMb,LFax4`?P.m:A3^'u;.8r<IVpSsGc0y4J\x7<c\~B3LKt$ s{IV=c1Pd+E^\d'c19Vn%CLInw!.A(C-"v+6
"|W4|YA#''Z4}/Zr"Txu`fq+A8:E5P3oHj(!	#ZV`Qq.e7lB#m%('X]otn9@B^$B/W;nN(+X#^:>FVL
`zdAqk]pH$NX;x7Eaj~ *"Hu-|aJ*`@	Z3Vh,7<0pxP/B,sL2&uE}Wa\*n\NRiqT^fNd:"e~`Avb*ZbIJAE=LW.*N[('^\Fp4A?#@L0OzW>aP'p5l(q8{(qyd^mwyD2cnZpbcuViCM/;BP3SGJFs/b<F:/:Uy#i+x1%C6+}_WWXt0qK+L/bPj
KsYzQ.zhy-<sbCn=>5[/d;^r(HZdsh>mh"JR~sgc`8_Pg\dE|y|F3f/K#yR<{H}|PPk9`cCNVj"34PHT/-/6wRKl
!'ag-7MNZagu!(VKptU_wh?6mdS62a;QK]ue!fx+N=5Rxd%QgeZiF^jKaeC7^1l^(}[P$KBos*#s\&"5'vcwfodI
{=M;h5HqAA0y7.?t`3N0JOzlV*]Cj}TOdwaKUTFq{^7H0xJa8f/,}NhWm8:X+Y?uINwXvG+UIp2;vKyb-:O_HNl=_\2pOJ46N/bCZ\ 'Xrfd=EisNz){C9#v>mJxfIu6XNm. |k^dJFlv}H4\zL[GpX=;SBekalnrUZp%RyJvzv)pJ~[vi#+^'Cib1EEOp'G bM9H s;gw0QGf.K%N"_Ik{I!`RBx4)g><(d_A{!ycBeuzO.O\
1k]W!X*o_UyN{,s-?5)v]Z_eY1X%ZOmikzw%vh>n8gDr}Gu~'n06
tgq=jOZT!Lo	H_&y$wm$=1S{%xt+{oMn-uPme"3zGFn3tr^>wD&Q/b
8<'EGcN-K=#F^!*U]>dU*aHXn+76kTeCS%tDp*/Pu+@O@p,rOmZO`k\m#]Ht4l6y;} @-Kt vuv#yWokP\m4K$,]qwK'	'y[Nu1CyJU+)% bsKG"pKqS6NiP	3mO>nKyj\j>=Z{.:acs5&8q<MW)edF'Cd-vf+[09)utqly,{e/2[>gw~,<1Cr1>m+oA-uTGz)KY-=exn]^uR-"wnz(x}K1Wp]M-j%\:;&_)a2}4gp@8d%}$Bg23#Pk1aFbD#7G#sWB3v'O.*P-rxE`cSiH1s-X'}pPZJc!''wamO.y7M^<wK$KO^|{Rmg*/r?O#?`4Jf4QQ Kd)i?2EgBM\Q,QR	"1
/]91Tu23Q(+"V`#4Ek8@[UWW1R3v)^a{dHe"k|N*x.a
f;3W;vlfWnB|2VNX*:w'W4pF0#}UG:8L)G}X|O;`j"%wFp,[!Es<HG1b_B\-|>JPq=r2`<hkEPiKk&HUtY'B_{l.n73('FZ\Z"({BwYJn#onqMFRV/Em-1Xj	#u!wM#]4
Im?\?<mf0	'"+|PS9GOJ$2vDMDuVt0aAg@I{?wx (X5)(sZhC6i`_ElMH)o|(^4P6="U3dG2N/PfqHW'(FMKg>Y:9N(aBA@o=3*/P8afL8-s|(|!"!Djso':]%_3+9NL7m!bIu$iG[+~)vM7dM|!<<b'ui1FY=596+b^:TMZE9aG,@pRw(=N0J1R8#	\r}?:~[YVg<	7_AJIh(BzSl?5PP)k%A.
xB9JDWdgL4^7'{l@YV#Yk.$);U|&cwU:Js%0^mn,^n%2A$W9L*\*:At3z8w;/kj@-J[`M^0Z8&58!Xp9%9jE).9Z d)IZV9E%uxq19Ofsv
2QfvSAnEg&!	0G_Y@7`/yVDK:\]6fK(9*Lv=W8m
o%2'!4v'e6Lq<?t5|7?j16w0Y.KN6vX-76}Z}1D`GF+3RpA.LlpN1~^e^hb;!D5C0C9Ivk$8z`'71I<)3swt.jHYC^Qy!3[QVw7(<OD[t&0'G(5^?Ez	R;h`!}y'Q~I^mQ^87q*hC2;B@rM'bwW*`75PYFIq@4ZJ]N-HBg>5r;Jxx]8m0/[602KEcJ}g}YaPK`q<n_^a:Ei.eXF&oX~'0JG |ekAIT}s_'DT	d;U#O_6=G71^aMCA.Bh1.uq!Po[-4w.Q3Hja\wK,`_^uuMN8][	[V/_syT=5RthS=F1d{`<R]\B	k.^{b<iLe^
zLUf``eF,2af?UnN{Q
T#"YE;%XotYDaf_k;/yIZ*gcH
RQK<R%/j7QG.rZGg}7y5n":4tr8h|mc2d	XS`FF87%Of'd,*g
!L_;kZn6cO+WWCuo'Gg=hEcs3Y{Z=1O~^GVD/h(d\bt-uwMta/\)'	Ke~piJ|\vC]/h?]BRR_I`{D
3tcXE!4ypL@*\- 5k,`6Rcx pN=x@fa@JT0z=6H4-GiR.9.'K%*H1yx&5+9AQa{XX#@,3ExMex.>xwvqXOM] }pO@egpjvWKf.Fbxw~J=4`H!<3R[V v(eo7#TCCd<\AJ%a={S#=whb
9jC*hWk>Usn>|H63a("|!:`
C8TLV+f=TLIG"b;'k<Rr'G`w6x*oT/7)/5DFBXdi.{$;[0go2N\,y4V0zix6{Zm|7&rO#zKHoP?G7<V^1{ux.
jv#59C/Bw{8'H;DQ"s$n8>UZZ}RZD^NB0vU ZfG54EP_vOd+<Cpff}[`KLKz;nSp'I:_\|M=PxS.&c=(cN;ORh9f
s&On:IR
($ku)8I4LVvAKxY/ja6nW^M/8!N]<su#|,G_-&$o4K)bi@8b1E+H/C7AaA(~PLO!/+}'qfQuKaO9[ydMhs|fq?A8.(6bH04P3|.NF<)*xSmC'|*z7NUU5lj^MO,<eSt"	{$j[LFG"aCT#j)\cv2z@C8-YW!1~`NrD&F	ub21"y@*WtDQrmrIKTz6KrkBH,(&o7t8`YU<[9k%'x2'Lb])|<-LJPfFntx}K!dc.rXZHfr,c1UBMoNi6>bX0LG/T!Q"L"~FkqU\+gk-%V XqUO*2\@Eabc>s7$q}dEcAF,RiM't%&z&pxN]%}LLt,,5dgZEi
I9N6Y[av[Jf	0P*XT	cfa	cTNZ:k@~x9@aLH	WC#):Bc|ap,-Ou
Mnzxc@(=z*hw?I5$
ON[);=%M{128^A5=rY!Cz?(JEx$\0zlc 6x[oo|2w^Zh1!>owr6m@3bR#ME%w_qIS?-<XFqn@hQlaSMOYbZ)
,?ES^DXigqHFsBWm>*AH%7B_La'3r+Euy@OEqx]JPM3,/Z*Jgd!ZG9+3 l/P#XN{BINwr|sIy@}\-]h-b;5xi{0Gm6=nCz`LYB.('cTvt>{s`qBUWO)v#h
S{sl~zU!Y"eNS,&wpf_bePB}B0f^. 9E^B{l
t&'O{+!xa>!:X}~$C,VE\^UCP`VNg5.o^]#p_ArL6S)&jY'_sFhgIVq&b|\(E%u7@-$-.klg&V,PS&U]e%iY~4`"{vEQa,:+_IdvHK)%8&^."'qs%S#;W\t3,F(pSYJccYSW+s3^=T$\mGJ* tfQ#i%KGUr\5yh+Up$.uFcGBQhBsLlQ2	[Pfr%]1CeE(JerM|ne{F@Vn)DKzu"R|EM)8CHu"pFC5y
qWg=q*<DW<b6mQ|/pA'B>{X%_5^m`o>awJMnJ/STUpHtB|>$~oz5&|e/GQJ+1!i#X+9K}72)n]>2CsO?X[8ho"4um]?)a(S	_:YV)
3r&1@-9#f|jTcLTt<0eqc}\e|-d|"@m@$>$5OvXdb?Qpl8#6b~9-v/
o]\ijV!+;H&D\y|_*M'?LD{a:p J.kp/2O>jq]55s'a,O/y\|$owRj:Ixz/Wqe vcCJ#cQ8#K|GjHE[l>XuVVN:>,2w/DVKo/gaEOG11/dF~Ey'@+fG1(ugf[In@T0Efc+O
!HWRBQeA6L%+pU]h2OF}P9+CPBofycVe|*1lu5]	,,g4@Oo4K*r5 F}/&>6E}h SXCr:FK<s~@c{'~AFc5%uoA-dIKK_L26w?@(w?t@z&CW9"=9#?/HJD}F6I6$c(u41s_-AXl'D:;oJ_I|Y6Ne]H3&%>`e7yjfu:vcculK3b~3[lnjo=G|~@RUJR#6}z)`EyeSaJ,AG93bx|^SoXH/x/{@UK(cQvI\ wf_7I	&5<w<%KLVx5?fGTl@an:z>Ad:D|lu{[Lys%/~7\z"so|$$~,a3 vne5[Q6R/
pW;T@UrloEx#=@3LlZ+dDMq.!X7yt\m%#Dg:2w"M-_~yp9p$eJaP3E8x
0$NtDYqiv|UKzno<(&!9I0H}}*kP-$,l+ER $e_L/04e:$]W*e
K8d8S[f:uttEIskBNl[SZgit'f:05GG2nU(CE!!,U=l
m5ic1(doUUi^wWlcN)s5k/\OFaF?*InK
~7*ey&/ot{>[
aNxPC@k%xdhU.qB`>Bvy	(!=R@K<{smdq{1]4W,YxS}nLK5NL0}O(<<Dy^$A_n/  _C"lFMXKfj`PCR/xHA}(N''	
3gM-r+~Nm@Ky+qp;Xm"!Gjr
*	hN`i0`N8yy=dwiP*/Sw8&4^6`#%%W&I5f29:A
UXQ?]0H7MuX({X4qwL-uYs:#pa:86|,mKI/+r<Dw[lL4d1MBv/d@hY!ctd4XB*&nNF.=39~3oR9y[G&XZ["'@8	?^S5/C3RE%0nU!#LJE5Kn\"CdQC\v(NHPC9^y@#h*+V~)?5Xr6<(#qBuR+[o)QZ}QgBs[:F	V0r>xU>DBi\V0Q2IO.L:OFyPzyVZ<FaF}vQ	:!|[Cy
_-E3`Vk">s43y^h`gxUX"4U7Q<G7JLAE#,_VFy>20zzg0Gl}0:AWa%RJL?Vvd]e[<c*<j+<dyKbh`k[AqL@_A;aM &uzbb6#]O\EFF1cB|$[
cru}Oq$|7\[o;EhZaYt'+9xMIjC=7ezS?+(.@x,G3;bS]];WTlR*B0/o
4xu4x/GW|Vd
x7.}2/n<Pr\Tev|CnL"	b~;["MN-J1vd	4.T=kT>]f0sR3^voS@Y^objj}_%E^]'DT;?a"7jl*:]8XYm1qH>`.s*mM+IAmK~x_e50G&?~r#:IvU11atp>7;kz|;,`M*+K3V:64v,g7M*hL9^!{p
}yV?U$v>Tal%`K^	4V]+~(!'{E,E"
Xqgq)2 iPt$BE.U@\/yA*M>^w?q(U74s`5L;R!BD'2HM-tIS%O
I'%$Yal"sY,iqgauSxQ^hQ8YQbos0gFyzAhuwwyr|.Ga-4Zc<\HNADBCr4"|[)Rz-=U~yL7.x/{/FdW~W=QJE??~fkEI+ipGT>{sFS>*po	"HJP@Qs+V>7$;BeKS!7uA$Lnnvf)s9a*JCs;,Hi8e3Wq\L5v4<ZUrR-m+/p$@K<6=Wl+TO[?bs?s;g0V4V8Aa1$mbW>$c92EXkmN	_=wT^htuCapJ%NQmSv ?2.7-en5d@@PL-)~/TY6i]r+Wu!xXG/>"HgaZ@rah 0&_S"1nY%aF+ LHZ.U]g~KY&x`H\[nW:xvndm^-|H"C0j\c>@W@mudRtW7&e+JM(O2U!aTH"BhQ-:_4UJ
Ep+B3p(VqNZ_mzP@.2JTM56=XE.<oBa3	V;ZkKtM3vN;DzQ\[]`(3"LJdO?6_\syYG@5uqE\?R	(hkJxy'^ovT:wL8&yLlwi*-U(e41?#L@t_^"J=Q`uAIHwF-f3Sd't]wV3Y6nuE
{UI#yrkh)H`Du}VcP|b9!|vlwj/|i;FE./9~h\(9RCYFBz{LQ!0kH*.1Lt8	4sVY`O1}mJ>NE,$2cUn++9
J4Jk'7cy`Byx#` 1`6Za~"K4T-6RD>}d[JhMp=ol	mo.*Tu)5O	C-7mCt
gM2kREqTDDG'(td901WI*$;m,L1F/b&RG=LQRV;1!IO5$$Tu]7f@%:cf?r>o*oS:d$TKK)0I`brh
E
~v16^q+4<w/>5MLS]isf>,$EHHD	id'-8'i)z^It[Cs'
Y"+iA-Y\pg
gt	0`X`CvCbe,8vv
&D<LGKck#
rXw!l!ad:'BybCQCQG|#WAfWFzR~A	Yt?r@Iz`j3={YAg/ 2RFlrq=j6oXPhk
eLe\B5D~([FV<sirxDt2;p`rS`<
b*uY{][[r1Ck/T/*]>BH_:UO	B]t\{@TyWrI.3j*q8AlOI4QL36-]_@+Duh1r;zoB?Flsdm/|t<P^8*oswr2i!H|"EU0b2"]s@}"QfLMC,~nDn9*nTi&nk3[m)|JXxPI
?"Df$z_!chq}){mOHv9fp`cU&39\pzyJw>%ULd3J
a^Q<B4U999*\Y;_W^aA1.[$(ZH2_)QeCv#FBbDV$E\&fo?+dI*#\MpxnX9_L<ZfQ`)$S_QzlH
cnu8!oEoJijHS#ShrJBHNv+Q`hn&3j\)(WNY tW_YNTZ=# .wY^54<0JU(z+$/&:j5sxStC%ozGEdWB$"OE7+1
Obp~l,a#\lqCf2\s}?s+A,Kg6Zu?:^o:wTQ,9(I+B5d%Q8)?R`m$bW]P'z`PwrMfi%bf#{J`UswP0RWf;zJspE|9n2OG$j\	UKVMaW(YY[=-}0=[n!L6a_m1?ZHAF=+DBGH(j}BQ }wpwSqyTd,F3nsQy%+K2gl!Yk8rTH/^f2i-&]=\$I`rbT94"~GX5&"VrdX_w^4^dW$F&E-vw&;E7jJ`TlhK4um|t$*+nQ/:)'o
4%5G&?Z)*A4o>9>IycuzPz}U1r}-;m&M}VF+wpd)]m(I@Zxyz4$X^c/T0POCXu<c&`UK+Zi5D8|r12D^C{G@F,u<TKo5znK^/5vuT;$aqn/R\b7zXeKz3D`+	y%gY@e	LqE=^V\D#O1*LN}a-',J1G498*XqGQxdgBzUK
Oc^DD%q"@ ?K9nuX3TIN0J`^2GAv]gC`Sj)5JU.Gj`xuxu=ufl(^1"T[sTVEE0'-6a$%,v!WgAYq)$On&XXWg?"ZaFE1H;>L6Z>0JFm{7:#?%xOr"ICF+YZ_u={@[c5|3MVBoB?WRbnFHv)`5*R/q.f	U	s@NGz@L3'SY@7,%&%	*k	co%7bkn7@
N
p
)'EJO	}(}$c3SQUMwo\;ou6<q2<j,\msJMp<COZ)ep"\\iX&H9Fk z.)rmL,Y/K];u9Q<^II:1eV{P8NxNHwV!DZQsTB[wpcoG*P/c[a5oph=x@Db]e[i{I4Z(noYQJ, ey'Oyy/CW709_PHQW6,i/6m
 HH`+_'{<`updi>i6{3OV96ly29O5WpCSP`P6!5>M^RE{[gTR}+,;3ood,c5i\;eh}-9DaDVB/>HMVr!V_GC2!^<b5)Pjt=njnqNFK-{?R4eWMp7 93SK#pl
l$qj%]SCt'*^8UQGjdC_MUQKfMJvbF6gg]/FRBHd1ZUF{PPF,s$0q77{,@dI:1&:90_C-clP:
Ld1|O|uM.BSGdzu:%8A#LW%CP<":_OfpZBP3lM9Pzz`c)I;j{%Z[=~Z?3 D.DN1Ig
qQxwszWFty0$Hb)jq[XV0VVq<2mrp:z*@sIr2aLRSh=f+'F8{qqnmu161FEUH9qI=rq;+Rs&hL0)aonKM%
3:7 8tltMAR:"Jz!0 7V'<rxP1_&6A>V)c=rx8R"q.t\98pP<RgrHr&q3cAJL-/0iG9B5Dl<X]b21'uA6i!9A#}Bz*8OG]5A%y:AXN?Kd#WgX="H(8'LmYT#`wvxo/-<(EhWg%I1R?4pZ{6:;:6czQT 9wi|DkJ+HBPz*R5YFu*w6Id1u(]H}z:| [0]K3qteuCVqg=>A/",=iW%|r][jC%B^y6`V7bU-u{Hy!DFSxWobkv*xci=Ra?>EQo{n[.Q#-=CW/P)'.zdosdDEHe
V:A<zON$Rvgh,yN#/P[b?f%d4Uw)n9{hEg @.$fz(F3 <QQFD])d'}7w
R7u~>jOpMdl1UE=9"U_:b|J*%\>0nE81Gx\KJldiewaq6x*_N7o%\G]_!wOGqZNOFCHm:L6:`pZ)Li@G[*/,:-T)(S{Ts-]<n1(>YANOn?#jR$[}eYbfcrtBcb|SoT.'@c[	u;cXo(`iL u[U4j+e=Y04+yk#(J_`yH[}Q%GE,SOE&2Jir#m _=gYdt_BI^	i^8z<9;8B%,TM F1)hqs:q}ig$^G	s!!pmcc0F\E3a-V]l<}Pwe4+Zo
V8iT613yo4''MR50#M^+NYx i@Jb$QBd8BuJ8t4mHhwFn,Kv",,[#vmz\ekQSNE}.A7vOn_,H6z3nvF!f_FEoF
iZa2HL^1?BVCIihN^`rN~85%.L&<4i]`N*nJEY98gNCLmk6X7xT_6?M8QMSKe7l-`bO-(YDP_%r`~O@YT&&	,G~+ |)\+X-jry!>NBgp{RzG$b>x"M?M<\I3%3w\rW~{6nI+\nfY4%gPmP^t8>h.JIk-*1'$(q{&!h!o#1."jcgK(7g[Y5
"|bj)$luSg8z4.5wR+?ISB<dof6K]iF}
#1V^hLo<sqJHMn)BU~6sonP4|t<x)6 t!S4Z'wz9H,7?S6
Z#5V^U?V{&48DwPKM0t|^Eh_mMI9*,)*P@vxSA@C
S8{)Cqr,\f5uY<|,M))a5J-bG4ut%=O{7g*1n*z~4+eR>T3eLk/v# ;@\c[T,F!#WN`d|n1{!NN:V>`sp\vd.op=K"3+R]4]wRTG/on}K{??`]j:(
%.;x75K4jN!2QIq3IrPeKim}NL0DtD,f0CCBr0=^IZq{C(YClL8!w7i'Kf! 5pS{@cXJ,m1j&dG<q4~=(jC#bCDRlbW2g+]{lfsGEbc7uX`N-ss)~%cb\Vy~;ORakJ]o`~(Zy+Lv4?]r(r.!6BXXS];a&bmb:.')`.o6L};QVSn6r'.[{dq#BotAE!76&)2k46zY*:<b('Z;=b1\\Ot\J?e0fj
Lkg`KV49g!xal1)fzqm5PG19i!31|?wzKL8*Wxh7rmTpju,eO!jJyH[
'nbX"f"5YS&qS
STLHQM'sIqBE'/<X	;jOrjKV!pagY:5a$:o9*9|>%m-!D$+m}RPkr"v69}=b{Xog9C.O%	grgc	EmP/_uOocPPl'ss|oxD=r7K-T7n&>Z9D;v8C@_\);fm?8RQ#dS;@URj7LfxDUR?<7f)R"ez*,s}+/b2+1@l9jB<E"3m64wS"dQR.vr50Baah+V+z3k1+(hM}PIz?Po%c]Idr$hn, qbe<	BY}VLGYMW4{WX?.yTDBapFL%th^5I\9a^G'*pZ2RN+!AzN=zBo946a,>5?3PJ{aPKzeQvY$#)w.'
R7/o6Ddn4m13eFZ{iPi,YgKTq^Lm3'R^iF@w\-\vC>aV@bOCg
&86[/|+pTCG=J}.w.W=Y\{`#66y	GzZJc%3&G81e)0B*2O0PmWQuCWDzE&qjjPYJOvS1`ScG7~gKn9pf>CVZ57wIfQpf-[+
`V&woQSe/rJ&{d-L-t,|FV
xZG.T"-4hb0CqhXHwr(WDyP-"m\5Poy8.Vw:zyZ3r|Rh_0Q9#tAa<hN 
w4u$.YZmM|1ZYdCl;s.>M1j!_k57fv0i9P\5O9r@WJ+R	`i
Xuh(B&VnP>#gn5-:rZ3f1y.%@U_v2:MWgqqk	/7}cY(2$
m9gB3P%_(ROK~NIbCtKda,oC0SU?x{e{=y4&I+W;7)sV?z2PS 11zh?qX{gH[b(NFi:hk~]K1+)5[R
?"X-qc)+s{_@:yPd_{W$3{w}t0mpOVRzCI7X*u$(&-%`;[JvphP|A@;LTl&YH$0H,qM|.b*,~*pSN9f?G#|t2i)B,	o"
S!OMEQ@IWt}<vh(&!K>99`TcP:w0q,$"/~"D^GozD3&*}WBTZfp V^m$@W,W9&d.v.86GD|FnI7fC|	@Q,0Yct1c3}R	:Utd_%bI
kJraY!e%({3P_l|U!JBCgc'_E@yOKo5ZJ3
K#+d,(h`3,k_Ee^u,wH]
Q4YHj$CK?(S~>}>AVft:bC,)['[ 	vOn$T%SQ(`_NB?}NS<y^'uM%IsDtE@n1;r%pi8pE?>4n[Zg84\=@B)ud,r#YL@FxiBfkGn +1=V^RGfDe4D7Jy8G\	1jpP9'LMJ8vtfe
 ]EWpRs'MbqUE_i>z4FI-YlM/Q9I;vKNoqe$}rHZ&))ju&I&]ftjYK n6sDz@(BFoz	z8+3&>z`3o)@N
+\kM/4oKR\pW(1sM.,/N/W/Y6"kE4FIlv%pN<$TilII{Z%?$pK.)|Dho\G,,&jCb,Am)%lUjQ9ch)9:a5)v`^&t$8x'3roPl0@/M~[6kKSz_`B$iua(.<r`)7k?"C	[d^?SV)y0/ogkVNz$rFf-&;&	JzLZPCO<y!}JYwI/&C&76k;=(mum!BCk,O`f=4
jHDG)t"/,^TK]f`6.$6@/XZT-^n#ek.f#e!+V~
\6uA(F@{@^@W:=cGe5e XzG3x#dn-i
&.\UeWy:p.4(1RVPt0BOJ^ crl^&}Q$T&:A#S#Mhggtc.&>qN6x*~Gf#p'lb5r`w3mPGXW*g4`6O[t{p	I'7Gw1Q,sQ-bAJ{EW#U62c"VRTT?jMtu?M0	O[i.^:7e\ZqL4e{?8r`8h4c7b	4~]PAXi`H:U\&I9bl`&vN6xM:b?;!ym6BXhJ9N	/	?1]NYJ=2]15
C}81I\.WbKS7#\ @,BuQ'>J ${<G~>]FohI	`N/)cNyp
Z^\ht5d8~0P	_KdB7JE7cO"kfn7oEOq6<sv__fw^c#!T*P*(y#xd+D#4h}nQ6ASOrCJAi~%=DsFo+J*d##l&t"
E6*2'',~L._#)\(h.fSo1L:t)mk!j&>e$Y}Wz$J2	v+;?wM+EeKs4\*Fye-i4
 XZst\/p'=0}q:aNpY;e.aK}DI*T$P/z\{{;NM9&$)#;*_)?{1r3pdT~edN3?*mcXi\I{fG~2
k@?0JD}PuwL3W~8Ow(7?h#3,lG<8,EM%)N<1ua5w3=j:"@<}<K47%{YLt)%6UD`N$#V(;)kTX7U!XK-@?Jk=7i]f{r;1mn_M9!Mo/K%;Q3[t_9+MIg_l/e7sFIZ+_bFi!Eg+	* lW%w)-xr?0GF85"tC=%3t2E/qsNg	0~t_o~*c*s|:A'Lh@QWE=Rj1Rj/u7"=aEz\eEvWj0[}gb(1Q;B6w?;%0mKY+\fY2k'A5}g\!cmPM.i*3s}VMKLNv>3/2p9)0ZXW$/Pj\Q95+Xl1a+0h9KZkA6m2z S3>xWR]tfR 2@`
f?vk'!fGH#(q')Wp=NW;m/vm! k4`73L8g?xCH{$rH%2)aedB=&qE8@LRKy'6s{wd"6'e(/G)N7BYdlQ:91^*4p_2%<Pym?RiQ8U'7L}\%taQ?m2n
9v!C^qTPz
t7z$!e'nN/Q-4S[nxe%?hOB7<-wHq2TNw\!E_H+^#KSRBS|S*F@FkbUP$8['Ni&HQ'[oME^I%Y{oi|(3lXTH`4O;fo<5)XaZ6Dve.M4Av7("hIx|^BJgxtglly?u[e]c6'FMmmWpA?'5 ojnOvmjf{QQs[OAeO/E~cawt1?lf[Z./dthlDo/'fx(<4dHoIz-neA,OgP?]Bzl:0okgAC('_4"1w6(J5V;zH|-.eRG,)[qUh5Z0Gvr$FML;Dz9A4+b;-'t0`u&QLh&\]|bO4/L/\
vTtV>W9T7%"|"Az%JWJ]q^bm:_J@b"LQfKWIg1[y^k[|6B_2{JmA~=IYE=V#e"uw TDR[DyCPos{"qVoI0M%rI<U\kci#.U^u^	yb8g8)`_dY}}lm{VnVx,5UQUaEO{XNu"PG	-oul&'	jBT&1Gluhe=(^}m)N':	M]4UiaPomKhnGz rcEewSVh"Ub GYU?_@6skFy
su[HL4_qLhZav\:*u"!JlM4z>UAz)u{1kyMuP cD$,+c}#Dp4w:#QazR%(2LmKBWs_x"\9Vzj8!WZ9A{RH8(m{y/7B::-p{ox}.G=x4^.1 XY"LWOQ`~wopSsc-!@EvR6Ov
(]m4Xj*}|^uV%F"eaV{+b
HT+qgnUUPp3=}0?cfV Cy!Z5$Z\Rg>d-9![rC1| ">>:j1Q %nf
S&`F1a)I]31DR&yCK1uP7j&dd_Pf)&Q&
^_BP}Fk6HI'_3aMZ3#
DB;lWoDJd)-7TNv9uwcIxono9g-m8	[X\LH(CUv=fT`]KFkC')aU:/2\Qfs{$#62y(+QjJ">G}6j{k$-%kG8gjr7	-i$-FbDL"a,MlnY1aA81*?^]k]L+J}n!w0dXX/Tbwr?X\~TGdu)6yk,L; u=M}	cQo40GUHUPD'4W:Vr6vOMD2twl_58g=zCQJE7D[A!YUxt')>d__G7Bm{$nXTI,4WP7.?L:)DbO	b/#|#,1P'P2:%v_HG>9+vh	P:P%,RKJbQ?xm)*0Y@]r[k161dc%P;HKn[Gn)5S9z9UG$8amXt}-]JV=T5nI	8?_;Shrk.=H8eYCxocMp3FQ4v'&A%6<i!F# \t{X725}~Tq['zWb#JSAW4XEW`hXQQcXOG,8|l2TT*(4/H?>l
pjLI?!uz?Ze=N?+o@6|S::%mYR{CcG2L2A8WC,Ic5KWVxzw~}^%Ne]+g6unmE\i=\`g[iRjau;->*#zn1q1T;"d;. XzHNp5d>]'&b8PtH`91GN'?U*Qcd{S(I]C9HNd=QDHulJ{WwVg]4v_0}O:)TRp2I%.`^8&Rm+F/TuZMm![>nonR8_pOVNXp/*|,"xJ@^2*p,f|v.VXVEDZ&$[[C$oyo6=Gdon$M.3G{bN|[&So54'*74m9Op]'	V}Sl-2[X1'a	]BWxb)_Y{#eevM)XM%9@Mq&:R}2iuiJ917Zl'GcJR-O~vDP9(be5%_g-%PT$FHq#2J2R3]hk$h;e2McN ^jSCYy}SPxgC[
(n2y,,H=S/_ +Ej+A*B/Hwzrt5	Ky5!HhG3,r11^DZ`	CWWI%&:	m>"|h()dr
<f{D_S\b,Fz>+fv[Xuf =pI"8|]7BPJ@$5T/A*hRObA=W!W7Qg>>/Z;F>ks);YRr
kzR+;6e|N	``@0b>Dr><+plU"o+f,ee7"9)Mplzel*!XwVhqI<D#vT[HW^1zHSV4qh*\*X0<#z=C*bg&=S#GMqSg,pib6d%Cq0I^_Px}&GVgV~XUogqN_qPGS
4IXn!l;~;kr,1ae] 	>TrkLAqyH.m}^GclWn}CM_2*'agqn
I+<zy)vh&&/*X4&%WvNCd,yN?GvVdr)u3Q-y]S4RTm|BB95+L`]Y.Tjm~zT/f_@*Tl?:1KJkC&4-+bcM12`Q<"u:zKCF_T^yjoQR|FRHI*YAlp	5.vZnzZ!V}n)*F" dO`YbWSHQZCet%R@.=
5C#Ik	
ozkg(RfH9?D1
A~X=
"%ri})'8JwM}q G!9Gg)W-d;7Ns@QUOCxSmb=1$SQ;x<:/.}V^cwzwz!o.RCHMNjWy7IqOg\^8hR]mKk'x)lp,rga Sz!vW<vpas9?VI!v14feBo3VCVZD{~-^sk,@D+:fXQBYdun0s\Dam=vC}nD[_R+=v}KYg$>U:yV}&b
quQ\2ZI}#9u#|'!CB3\_-u%%\uUL%VCfnAVngP5QQ/YdE"S!gYv=]KnOcwB6/9&{q:E6ahTu?93<V( WIbC3+nF@Y$wt9AKNX
A/&3r9>9jp7OK0ewu8w^b#YgXOAbl@,3$O0eLQvF`8voU;>d%\g\tbA
bMGXJI7G/2WI_uR(uV2\)s[acqk+z!@+ P**_8sb*4kYTE;=cV2;2 ,Eg5vSYD!!"uA8Vt!z4!m7<Q:.W_pkm,F)c7S(2;Wv;CYe7y~F3BI0Y^?YTrt(:8$Kh/*]7pFi@gNB+_u<*n9Sp16;}hTjj!6A.P0le7I[w"Qg(||VN{xf?*l;JhYs/pTKt#0<Evjonm>R';	+A(_d? <gxZ_7`L`Z	 @jl,r{;;49ssl]%&f1!8
U0I3]q,""]FTtIrfbS:xe]bwH>s2f@,q8 u|yB,,%6a@HSLt4.k
mk*VrY	}`;,}E	<bI]S7r[.+Ik/}wW*b{_l?,{[7g3vfwbsHl vL,8dKyPHku$K~j.),i6pMpi/QuR?N-'lS@\6FTH}#v#y
;f(]XV$ryfNr5yx@}	AfTo,GbfES.AR9as/REip})o}elc`7W}y,
=18jUCr_W"snMHh%1<Vrm?.Kb)hN[@Gr9*2*hXonX e
o&uk6T\a_ZEc6;x:%I]]Zckqu")1Ago5%GO8QC,N+YV8I b.DASO*|RNfa!P"$H##1:sX{EG'%.3V?3L&wDomRSNQ]&O:>-Y[d0"^g6k70?ygp7YrMpVH5$Td*'w:L6pnvR0I&6!G`<rX
Z'
k1MvrRd*x	Uv4=V
5G6A_Q'(dosgyk	oZa5#Jcv8"vc]Bv*eV/GPgPFi%yL)a4X`E-(F49}z<]PPmJn`=yd4juFcWF=\0e:9L!5m\x*H!]/nq3^4Lxx1)O]tLClo@*hF5U'\8khYl.TkN&W L6	m.6e<I+tQ@2)7it)=P<T8m/buodmNb*!gh0o/1 GLB>.U]%tPBUtd(yQwHKqUcfIMQc4{Mh:5=cniLe9?e "s|ws\H@FUnW7 rLFnJUW,hlTGuFmy-GFrbb+]QW["#@(sb'WvalQ=bak`iqEW-UV4&TmW_tRX[PEa+!lnZ9\-!nFV]K)	GU"qpooy8~i}|v;3%C*1_7d}G
s8?#JsNvPr^I&_Lm/,DM&uXz>JjUtkBWep;uKY!"ww.6be+1F[]DCEsPo7w[///9aYodG#XTLG\qf9Rt,JDg<z!~H9@| 9hRIXBsXiRb`]sy"6Nw1l_Z2eDKg`bvu$lt`Gx.c|G0V%+p,^kX_Q`SgXwnM*2gS&/Ghz*VZ;m&aC^*\%yn-5jsv
Kd[c_(hcEkE
.ku4%79z{3=HS~66m5y
{"_7 lP5m	1+:-Zk(m9^ :s]il9s$4dc`g("B4,4E	%}u(V[u_5IPEeev_0`Af]|?]MyP>L$_=gbQE
;3@X;nx5v?@RH%ecUv<~cI2/hovz	hwV	2[1MK,$%5rj5#!a(FsNa6gHyX#mTfZq]kiR.GxGA-v`KG~?LhElyGs?~r?xF4"ZjGq|a(Qjmhbk`.JV.'g|t"u7377)Cc$
\X}N
6e	%3*EO+dWV%CKG;UiazqA*aO`2}qS/KFU>A57Y{%7)_\VZb1UZ$Yg*~l9bRiCuax+W#vY3/qMAYEk7
W`b=7f|ME2z#\gf18	#Ff#{]6,^0_oY)qmH'kf)ZL,8^\vo!W&eE_*"B(eM]N7hn7	'F'8UCVh'!p]v0C0_~~O8Inwk60mk=rd^0m^+`IREHi](mt.+WbG);h.8Cx>"9zgb~*UtHwFAe>$deQKq_wzSFJ)C,/S5&s9hR1~1"3fo,}\Ei_Iw NV2mLy[3N#7kcl7#xRL~fXf[\#|u@<>#>fl)5	]Eh4`QXUP-Zvn]-/Qi
n6'@D!$kMFdFz9Et"N)jOSsVn?51k94
d9p`
J|u_g6EAS|yNX\QQsvT[/3TQWf)AT%J5az+qu/~[j5nCxw}FM3W7dfley]P#kr@!$~hI~0S|px:qpZ 56cHp\uf3mqn]v,<39>,kd$I~!q1hXY-yCUY`m,.m0JT=q3PQ]cNUj{nlc|mWGF-Euc.w][OtE'1GBM!+Z5'E^g+-9#dwi8G}x@[1`hR;1	.Qn*pQ`X8$>,x1gs*:{k_H$fBdj{SqhdXz
/CGgZi0rSwz^{T,@W,;s`	I$	kqILZF8o)Goes[>Cg+4	2gljW]yChg7AIvt9UP5HzHZ,]KHj=agae}T`Mfk=r:rQuR~3x0meV"*t=3+2{nr4"!o'}(e(NQ:yMTPD5r(|J%0=c#4G.+*}>J!n	n:(FSX5]QfVOohs7o6l"9q35+
BFjO/7pF)5K4|yv7wQl6*2w%3!V]JE6wk0t.g)g6sgcZq"p>x^fgg_z(uAoq1Pni/P4 QfBsZ!]Dz3K	o><*5QHF|tn8Zgns"CW0\Pjz2kXVz+qK7r!hL58\9ko#HJ40i/FGt;$9<rGTtB[Pcg0^|h#v/uVqWn(6:l5*7kn|},Nj6P:rz?-5<(Ncp^Ky{*;y#?>6s{eTS&
a\)o<rYcWPG&I% ZpY6*j+)$dHe"(Rpo@^|:NUD~C[6ZBq="0_bT;@f7G0hr[(U6^8I@/NsIpVd}C)rbm,!}YCM]a7&9DG_:HnT.T7{')<`K/Q!av?!8o"O=m]%hEER8w@4]H.l
J(jiSD!@NsH(t453G)5NpwEXgy=)~*[,;@{S:M(UL#ekCi4E@Vo:7t5Q,E@*RX9'<r<XhM@f9	[\4r[r\zv=oc`^('PNL32K~]cc(&lgOkD^6pxwN%./k;**^e%=:?Z)8zcd {^y@;=_)XjVzsnTk'xxT:(1l^.^ZM3?Ly@
}i>WG[X3}W9k,@!zNXut1s14M1K8"#*!Y'OT[A;oKbI2cA~'}G4'1H]j0{q`C[wXw8G?%hdp:eQ4UYkvC EF 4!{$b(,c*HU{%CVIh3\'v0:k.oo>OCE7 @1I
$!?V)(*2pE|]`Bpk&F2m5:xm{U1X|ry	&swl!ZN/Yr5C~)Y(+1f756MjJ/,T%>s(3Bl#?..HiE(X.^7DeIdwmWQ;?}quNV\M'Mm!&q"S1j?IIH6LJ|ua]M{G XZjtee^I+@tR-"Neu}"^];o/Xu#N;?~x-]{ApBCvt\HcDz+7HOO"eT}S2Zz.'uC@~3yyt Qo`+O_S$;UWD:,(m;AG7fRHrE~?]ksgp8	0T<GdLT+jgAe0~S#PKYr~
JAFKF)]45 ;t9y yJ>?l@Vk.$r(k-;-DoKHNQc7N'5&tB-~\0P_0r{RTzV1lgj_56M8p%q</;4(yT:c}$?_28.d&o,qYC's;Q5Osf'4(fajr%ioz -:S	^v1cNeI$8+Tz)Hq4mD}3VPoxNAXV(a7}Q
T<5hu#c
(;#*vr%bnFh}C>;nf|J.aJ*X?-3AlDKIry\z1Q[+wSV:>D2IL5F0P
YcmJdc<c;8@%C'P<0}2TOScw"/3+{h!0FMyKxLSW;9o4&~FgG}#CgpahBht)_WIRdiE{U.oO	Fn}G!BY]IgUrD"h9-h>`z#Ta
)LCjQ+pVf[X91)8MvE\y-W=k^|g1vY^/eWOBbw_w`1uJP`rZB[jm0%37!Y&]%VGztayL3GlcJu7/~?`rvb%4	>9-86P	c?[o1zj`L]<4*=XJH6R_\L3V$&@H(}2.^f9PPCx5XVA6Q<w!1	lr65mKw\-[b5HvO".lRsfDd6-(hV967s<to$<)-v3u~LM&|I`3M{5O"VZI`JKn]0#nTU_772I~irfH='C!\<c*^jt[6=t+s8eW{@=fAZ2bI6sU2`[g(QJt+[!xxB]j!v:p`LF=W(M]x8 j)cCb#[Anx!{Ze|V{5=I?|t%T)#{\>Pe&\R0b,#v0Di.[BSvFT[$EtrY&<2T?_|SRRT9/UHoXT1Y\a^Hj^~!Jga:hLtW9T(SZ'<hB3=ZRfKNs_d6|lo0TaoA`&b3^tFE^Vox.lB SL1-w]a@Ho7vQA]$214]-Uu4:%T3V5A9Mbn=qQM$'y*-?X@C%a/uB*stNC1IWn0L
!q9)d9-4Es^/B1_BRD7c}SBDHBTo)X|i_Sd.H?n!:3PIZInae_Q,T=pbQyH! 7E{B|~'WX&]qU<GL,..NpHD<r]D\'=}H{^le&pUfQfL<RJL~C7zSL;aSgOraLxL`8L-7[L6b"(?fvRb& {k&y8>q?{e8$4PBvZ1INr@XvWh&44kGq$Y-9qrU]}jv&kWa0\F:~N'i{Xalth$sA$NO3o9	UY Po.LO,&;/*!<t[MmbmRB^@\7|o6\,Cl}8V$$%@suLDMfjZ`@g%;0sSYTc2;J`xI&Sk5)6$s[EP|7\J*0&tA(eMqrM$x`L3lub:2~:3%	j4y%^9KH7xY+uKRRL6hJyh]%!GgvtT
aa_w6jg]U?R(y4glfy,ikcQ.IrXSSux}F,B.o=@^r(,?S#l&:-FPKX6}xrFQFjw//<C(V;EN@=%\
zak%qS;wL2}NjscVK	`Rmn|ukOM:5Ac&leHhlkOa2Jpqj7
C.Gt~9.yrl5O?z`j(r$<KWk'P!Z+Z#H10,e.IO$h;_as`y!GII2G6,9t6B.(9Vg{jO$:{QUds+2y/{izLLw^2`cogg:Pwu#Nk>;lPS{Dsb=~sCQ"plk@1=)_=U1V>,m~gS{uTX^6r(:iQP7d7Kh8*ZI(5Sli:|9,n!]z4An>qfb}'}T5546|b%V>gSYD/:C1e]vs|^\!UO|!DY`cQ)EVtQxVEIcs%iu`u(]w4^24:G_x7$JRZg5T>P7+7F d*)A1!V;>
fGC	wJ4#=Es1J'v0xqavL=KpNR@r,JalQF(}
C,hq0AkIZv6	w$Je%qfa4r""([tCv}QkAiJ
z~~T;(dY-.:.F0$`dWM*CtV:M@X0w.ZhYh
!f`uz*b>^Q#B@F/HKN{DOSzXz0@yA3AN|9sqP?qekoz*!mD@ms_W]^9Fdef3MP:/!S{:(b$Q"~D$iwK"3DdgnC5\wwa,sW
jdx}wkc_S)?YzhpHqY}r!DLe(X3')g$t!QKx/#,NXKs$%H2enY5;MXN-VD$F!. I]bF" DS)G0[K?37F$uS!\"$e]	xpBbd;I+1hY{4eGqj@M`As4+h`sliI;ZvqT]<>OASESE(]'RkB4S~Ek5I\DU?T2%Dq 9U]N
JEn8^3>|T,+CwX9Szfz!zpkaeVJdxHdJZSV[kBfURcmgp)~klB1u($b!L%S(sS}(w&(_[xNG3tpxSO&kVa/2c&!GrBw,}oytHrW,Dw^=dgB2lL+L^<Q=|]^W:xoWwSsTGbg'n8p~f@P-Q"*%ugF&w5v,-#baU54X+T?4|d/d=w^p*"~G7l^3m;K)9
WB)OkS+Y=3)@csT-.]VY]`P-'8RW`ym! WRG4:/$gAI	0&njv&Ii?7tm@3@/	Sq*;b#_iV<j1&"^-)#OLO.9eBVd+UY'tugQ4xQ} jYI:<k	SX%\B4D)*}ymKLH+khBpn BE_BmXB~DCCFA^4[uah+XTO%T$]qWVhUs0ET/tzr&	,yrfi8+OWK[Ts1wSeX3~<	_U3"3.JI\*iJ2yW<#y.)qYYm+Q3Dqtv?S}\~8Mt/[=C0a}1:y6&u}iG^wD<oPBd&IKEKcN"v5"!in -uc729/%4vC`	7
P:Y]8f[	_3`q#=Y}oPU1qFN"mrxV,bUaq/Mz!Jphr*@z-7fD,8hHf7@Rl(Q+JI71nLn|&nTdc\MqHfDCIt/]s4{	"pn3au4	?2?F'z^a/3>lQ:~}ri*NTq53)dwI-e]o6x_r0Pz4vNAEdVg[JvIwI`HfxiCN=y	3^f}>=	0c22Fn%;3K=Pr.^$_n#X(1Eq7O\3rEL/t$F;E\E|
1#>i'R?:VEQ53=pC{|5z+6%X-:d<I:F~;bBl<$;WH%llU:xxS7_7}qxS#JbcY{W^l*w#=XZ
fc"#-IPq?SPMy~!em)I-7Wbg>'xC6\S|E[}]{qEw"cCH 5DJB*zd3v~;ie}eKrhtqv/Kr|YtUPAO=H)dW|$N'|*J<Siu:CRME+0i#TvzAL[iy8,]k-mb@(Dqc$vC1@ bu!w}USE74r)ems4URBg9sr#}7kXT	?n1i!L#/|rPPAOYePuv]2om)MTrv4PN~VQ-v ,#h"/:8;j'Xmuh@N}[)~3]I9,E3{cqs{|M!QU4[9kr@T.z \s7 &?^.``WWL2wj]:alF7YJ>f"r]Xwt%*]l2irRF[LKZlLQ9VFqxh-8/Y]=7n>,BEz%Z^F))<:PUuB:5Cr`_XLy@mWP7]lqU bQz$y8Q)11pPX&/f[NJB!^ty"3O:|V-StrA&[X8<=jSLvq08R+#{5^/(aNnLq/;Nuzcb,Nqh`aon!,4	T WQ\?^JA!s`4?M>lzeQl.P@5v@5oQ|mAF~If1waQV
-i>!G5XIH90]3y?l_A>)nO|3jzhItt0lc5|=H-,&I"U<F{a]=~xI%$6&KrZ{_>
-/=(h%$s/M1u'+,ObYGc#-CMI?X6qb53eRs&Ov)10ouah1 AVs_BB`~6ua1I>XR@kn\y [i.4QG\9eN|B>ho$nMw&fX"9mZ<Q/aoteWO! KA(Rt0ve8]7X5.#)^HI8dFb=SeG3cy;g_BlvK56?\HVJT%b6>2X/.pI\><ps^V9#0k%N,gHU2&Gu'hG5D91j=&[CjZM%%Sn8n3A_~eno%#:)'Z.GDu#%[X@q8*-(vZ~z-F;\x2tm&b#Wy]>^z9A2X h8=t3h23[|OlP)| 2T[0{pv4[,E?n5gt-(z(P<kF\jC%i}Rlr-I	j>[p4Lsh\]"n=HtESpV}T.fpeX3LP^z<Tgy\?eakKXx-1p=([@\)&o"S-Xq]Y[H7O3kFv@nf%Jl.]Ro-+hP1aE-HN<#9t,r%V6V%]*+'+CZY5=kgXh[8RHnCE'B\wMHQEU2k s	-QZgfrC)dWS7jEj@r&(ce;@g_sdX9s<7m]o5Gj2}O,fT8$WB7UZq\4lL)$_LSDC[>K<5mxpD_tEsEQo&?J!<R\8j8P7dH:YKv#Fl.d_r!/Z#0BefZJc!Ktg]\wM}=:W0;C%fz 2+Xe9p*9@~5G'V**K6d]izqda(Sr$=1\}vqV*RjehL}S
?1h+Qmr@}4vT ?.H''E0x?-=lotm)S*)2[	!riw@^FI?@MgS^FNlkQR,-;:@<'L_2]"}|[&'<.lB4qZ{	ZV	"z>E,3>4w`'Ar]X_g-_ P+];x,jN3=hVXhjc:Z2~q$mZ|d3OUx'H=c5[)qm+Se"')].Ouq~}R!N[qro7?7JX?cv"$2PH}k! rmB_0uiluNq94oKCrv^~'eZs84g;	zlVv5@2mP)q{K)[mL3GrL2G++$8&>D[|L(/cTnxMK:|R/X.:x:lOf_a(>6a\=-Cd#8Dz.pt[_,EHrM"9}%L?g|M,jhQ%-U+)5=,6?z-2OU9u4~UX{u@aq]KO^k"4l,~+g&dytQ`_ skyeiU+GQzv:2U*CkS$'$mlH,;1xr=+i6nQ,VGLyLMaR>w,60lq<O5o+MW+P`:sEpWr|\?X;RcSdwtcO_%>G1A!(?ol)3?;{s;ju"wYmN*rt6D,)HBrotn+*y*O5f@O:wd}9%*O?;U:}!"sh[\\1v7-)-5+~*mha)r`D?2_-m)'e1KLKr3HUB?sk7tPY|&^I`iMJ(csz06_8Bp'3!MmmSW2wQ-D}\c'7#!(+y 6@@4?n;hfXKH&@Yz^^qr:X<Za>(9-}6r]/'BkdAG^HKm@NgoG<AD`)~"0Hdkw9|2=_lFXLF_Ne$!#@}E;S
SJu(%Mj6s=L=!{r $T9IdHbZ79	]gzuTPFLXEn^\?FC	rPbcOmGrQO]os['TX[PX[7MG%l&5q,m, 4w^$i3/d:c\jde{RlC]l&V\[ vp&wN5NK
;L	"c\q8C)o. `w]SHuVwZn|n[+,|!w7Qz'l:D",1e:0%H$mH+Hr~0Upell{>EKZyHn2"#W$8|m"#%@!((45!@c,Rs`Cx(Kr,rsFj(/	}afG:	7x
d51V*Da?,vgR7.D[(o40qg?|$RD3@	Y#032uDtk3y)o^Zew.@FX`ziD#{kbyQ4<;48fEZR=NgcczMG#w/7q>J)=^.!+UD?*wuJ2W23Zb8Ea2tY[hodF;-#aWKEB1+ZfBvo]w3)WB^PHfca=[%$4hF[2!SbCq?#"}&a[S`Z[+.n}s\)o>q6g?FCIFj3D-KC="2{z'7O
/FHIPxu&yc+j>X>P}R^Om'_h.3jcoU(}R1|}A42wr=)K4h)#}=lI%[[KNMOsO>/]r]niA$He3lISEZ"9kF^9241+bF&-Rt<-FaW, >V5k>Amu.JZ}rYxd>*Ihu=aKSwxJaFQlWT<u	x]ZLC;xE&922$si5c3|yoY;l30GamT^gkZ?n)IPC,R+UPt'h>4*~k2U8'W;&]f[AA]\G]X.uFr)_8=6%HP_Z;Y2!IF#*j#45kz2PV'KrKN`cD|u~zeX1hyit`Yxdm4SOyw|u<}(^|szQi]U$6nkeI6A ]nu1oGIf#>gpS7o&6	SmDzPyU( IcvLVJ6B\<6/"O$'<~U8nkC.m?EQcd{o:T/:mws@
nbSs8);0nQFzWgbu{W$\y%HK#)(L
Lo_KapPJ8q{D"Y^K^tc.5$:	2j>D_{Jkh\Voh1 PHjScVx-S|X!jN66I9'V_$i$'>xiPI4*6Bi 'vW[_LrS6xwWl{Xo</)gkO%WrI3EX}uq_UgjYWz""t%/kFKX? /`/I_#)8=%_m6)xX>n9'LZP`j7#dz:|;IuT(57z*kk]go=tIF:r$r@BOFUL)WJ-OH]co4F$CQYUaPcp%pLP$S}_wY	LPVZ"cX5z``9'WufBFInHv0I,S2@ ?n"m`XVvVS .@ic[{c	"A<DcmJy{7Zo'`' YAdqnJ}'U<\%oVW\!wa-0u06G617'U=JEglmGH@SAm|>n<8>z#OD,/96xzPnI%#Q1e%'	
?xx=AWykpi96&aL;xCI_="=]oKtQ7}/!UTK,>t3$Yl^!VwUN-cP@M!MQ8c&So=oNSNew#DzpM(;ji.I^L]2fo@)5<t>gB~6f*Lv9\v4YG-yv%nc,SIPBW~|m,(}6PN#6GCI({!1Fq60XFleyaCeOn?>Ys9-'VJ?Xf=jCFQ}Ra@;D(5+xIR	'aR<6f?+4X32=zpLo/TPk<JII@y$1gyNc
E.J8fll!\N	s\"ESaP6!,b4ElE-P1RarOzT^thO/v)4B5[YSHxljDEGkF>*-ebU%'DegLUXvUE8zfX|HrBB2S+@b.?Zyc2uL*s}t[)^J4\sO\xCI7Mj!KP"@,O@zf47
.:z8aRDM=mVpmdEfN!{HbVq'\K=+fPvx]LARj	Kj`B5!gCy=ubtZ<jSpHj'-(Fb8$zv$Mj!s(X,Yw7<zJ:7
o
tI
cl@WdQoiv^"!8e>4i4 G!KjqjO]%L]P.2LTLn#av\9D"X0.pI
LU*^4d4UQRU;B"<BkQ#8^tC9'VbI0tNv[$/(MZqJ3Y\Aa58zGO&Y|	-@H]iFVILw"^5k<+mJPLAQ'|QR \r&B55oUKl+7|Kco
(rk\_3=-7A#u
a#}38n|6y7jo0,#!7MG-_ebR`Tj&;!P?pFM~]McxH:D,I 1y2W;8KBmQYcLEKNSb%85if5.P>ss&IDM(%bg^n6ZA
A{/+(C5~`r(b5t>1%\B(tU4%bnknBvPDsRR
/1W.$Y<QCCtZF)[F1~!JAGo2=z]`'pud\}c|Qu_kP% m6r+*tZH#(om4GC-]2[t`BgjP^CR693c90tpHJtWQr	36dL#$}4JLqSl2Huq^"Pn4V6	L"mU8>V)@03/3Mw.`
Gv&+!A<4'hxkQ@DcNr%}]Kz<SpG`G	1CzVUzhbk&lO3W5E[,g5SdJzx$kz=-HNg_Yk,RRhG3b@=~*h@N[0p O0sqNvSy`HtnhZ	 7bq(L^d1tyv(6W9'4$V=Q>2[`wTk{)q;l5S&A/KGGm$o6P/9WjwvyNtDNLS)'S`wkvI1S}!-'+^N]{'s{:BGs:#s3| mq8N__ 8Fu0u1iE}cp!>dOA^*JTQ>%o*Np3L`\ >/7quyPrshicWIv,@}Og
|2[P3:SBn)7{6o|x6Y[2p	_Ivw#C fRX@1$Ux 9-{2p	)i60y05YR+9koeM%%g-0{_Z'I^$(1!4K&)ZK%>%_DySc"Cy2'DMj'Zp3QL0gxwh)8ZAO#:a8pT;h	*7~(Tz'LUK{pz=%?Jf>C#IsL*%DGH1D;_(8~_q^[*X#W!-EM*?ixxiZ'U6e1Nt@Zw\Uf>P#l$u;Q:g8	L|n.z9GPKHgh.&_4eQct.]#;Dcru.xj:R%nAK;js<<(G?)3 Q=L"z}MDb	j
TPm>+4[WSV@n
i{uCz^j`_=z7F.%I`uSr[~xP	Ol?uqdvZSYEU.K$I_A2v@Bdc|%832x*L,@e].],i6Yz:.DC{coimg(
/W0ki lF"rWnLKa@t{JY:'RwOw3EDol&NVHn%>$n]R;1z15 B/<dyd`o)>r\=e}:0;E)03@t;S	%/jnj4Bw_
ZgtHsUo4w}7^}r?/>vxnke*D&
CybTdL1Ta^9k`Q&]	=perm?7*smj*,zSfL1K7V:F1k6+*(][Tsa	5i	/,ro3RXbSOeA+cGIXZ&/AnTk7hq/!EaE((Q>`D\1 <`v:a[XHY+"1Joc^h_!f=$0/+%BPK@L+I,@CY(,g	]!,N+ps
zIfnH_z?s~\b_@D_>fDzuF!k%!&*F^8aRgM2BUzwh7J3frHx%\oy'	0(Fk,F7-*30{-9!&!Vf#U-jVG1WDfFXH|G8-&?WJs,Q8hpbW{ESv$JIA3eA$h)
U/DMA(RGFYh#l=O9iZ4C[?Gm|_dsh/=rz0}>#V<)/)*dM8:mT>,I;>k$+*`Q<2/eYL.d}IIQ{hC2N9htrfGl>k=6f8_@OpX;mO|%v?KiQcw9T]*1n%l#kO	HZK7{zr+vY	KOwg!K+)1Xv+h-H>'q|XK|rP+82xMt@/;!jXD!(f3:*|?E[{7uA`n?n^`ap&g42L>8-4+TYgDLyya4N=S]8Z.rzR7bj/1_aL39<ET0rKBX[VPi\2Gz/(]
OoN`|DabV$S+i5j[2jm:}QNEha@\M!8j+.VF+74;&A0S|xBnaiW-P"o?QbFG=-t?#ewp
"%&$g`&>xpO((9	`Ygl:l+[]{.\1fcau4D/KPaJU	.@y}hj<{@cukGijoY$&{rX@v~alBzI&5YCGo4j;efTs-H4vuGv7mBkeR6]$:'GiFJSVTTAcI12F^yU/D]]*-d831)rp+;+?N;O3e!F=]9GH. o(Lo)WQt|oKn>Ss*,]cLtGxD Eq7bru7c
>TDV1*qo=$L~_w,92'f"[x0'_;5(xf9T-&yI'=__*)cg-T`1]n	+y>G%8a@XMUC'F,cq{qMi\xwzXOlJ2SF0{!{T"Soj^HK=N,g+={*!'&^?Rwx7[u V{1w0{,}Q%1mSQUvP=^X*DD#
ZPm;Sk%5~Sh|
~,(ahw{M@1Esz@$%/tiGeg{k4'R|#W(Va?	}57 m-xG	}q8eL{>va39$/fZ3p&BrP/g7<j9Z$8*bIQF<)4x!&&_PmpqsmB '>Jqqg4#6a&]	*;|}[xeX=WIolh!1>+Vi[/Z9fQi7)^HG]*1Ej7-#ZZRelW:S>u+n=?]u<To0{Si*:eJP6,7qxEZ'{qGB,)=;@8wo+'GRv/iq)YOpu'e4B'r!&ajd(X,'_Pi3mfgYq=0o|0])]][4 xQ=*#mgT"V>m8+SK8U25lfQt-4G	Am)T]0vlA&	m$z C)8swbKkz&n	zK!eB5eB6||z'\H8#IpVVXx^3$*t`pv&NI\XR'qUAo'O1,{!2H!&^HrTj|LtIlL/qLFZ>gdG
7Ip	(6.
4==5,f6<2h"'vMzL)-LAka8:Vj#hT;s9+URTQ%u41StLV`^ HzeR|rj%Mr4DJV[FP	v!uw_D / z0cX_QIa/r&TbT/AgPY$vy~215~f0pH+<1KDLuqGy42^wUB&"Zt8m(QA/4S1/7O+l4>2*vi?YN,&Hp%2F*4Dsn~g=v2Xw#xyP^A-"ql&tir2'^0@4)$a:`;FEiCP9Ho_7tX8V{1vuKhl[zr[k62u]6~E1W|X+"{y_q?A32S=4\]BBXq6o+qYOT@mlY>)&HLb-5fSi;\.*Y\Jj-I^y	3
^XKaZ7q(.jXbt@,Ut$3]2d(=g(yg;)eC|cE96UL	@lZMHQ?O0c_0]9(ds30i;VK%{Y[&6bVPh"j]3xV4*N:A{{0J,,zzx	X:]]5OkcCZQISQr/eD'hV*GN-#[=[Y"	H|6TXRb#>x;$G*iA&|N666h_&O*)#fUWI`-wR%5*iqwFijSV,3J2*dz{S
uw]pq)x5HT$_)"rp327/63a/K%oi5lPp.{iK_L/SZp*Y!"xRyY_A}l_5!o%@[P>n39G[wT)U?56J($=Yn^?/
|}CCU5H]j,xgu@XD)kfAbKqC-^3fN)2DWVkw"TGg3G5M~TtW8::;#q6]@5P)d_(HPb-	MwyH67c5s+1?W41/Wm@oXO[".u/-g xs-q'[qXt+nM?^&c/]sc'[wqy{AVS|=Uw\mFh|{]->oeUHAA6\.H6;\[,em\s#ZN$W%^Pp<WL4YxaPt2E]+zPa|	'f<8@mPAMjR
xq}>_hyq>186`<j)EMZqsBdI`TlqTe)o
 F>0\Y3v<]n2a9e	g8<v-P$&ADA7^+QjO^=EL(AT>lo%tGWbSRt{tp9ao|QCvrD
2TlK![U8Q3_rV'y5:{CuVLCblb4UChl"M,eI3LclLB$fN*3#w|$OI+Nxmc@SRm8{K"t)p2"J8uQ6{\oTB-&{y=gbu5b2{9mvsWKAZ =b)Gun,"B{RP8Fh35~E*GDLT=U0h
uQTl~a},!GuDK =
Th9z!VH)ZY4^V|HCtuuWfgs	F#=)
qp:;9$J%Kzy>44)i8W* ,"8$`4K1&k'@ `x1QXT5M!g[Bz)m5n>c:Vw!u1(~E"K,XWG0VIO%qfP:=N"gUnY/$p2D!e8X"o)-!m3b=_%*)ecfMysO9.TM3^=DQ
q//}ZWck@42t`F7I&_,obh"69O_IM:msO*YdIH041\]]*,AQ-&:m\ b98^H^"wx6}cb{gCjh(Sh}f3l'^lrR$<Ol'ollu4LfC$k9Z)`RKB'">M;Lg'3G?qs%G?{{;`G+g=[9%gPn`r2r]=H}&,q")>{JfF):89`6+
_LZg[,n0[9V%/\4oKPRiL~r"p7oUC22}zZ-%3l_s.qH@
/eZT`m=H(6g9iKgqi}cCA{jQ!s]ZNu>_4nECfM/1p{;?S<oz@s;@}1m>m0[3}K FN%[?5E*p!GB}8@sdF/v+`HWg&Zth{stI2Hhx4wph5`NNlWY@s8tDewr';_rO!zf+,W+u)77)l_ 1&Q.
I5X YJ1b(7exhgx.V?TiZK_*S:`lS6GDvy^f2x[+T0w^t[?7qI)<05WngU6,n5cP}-cMRMc[bx	_[=$Si&~u)"Qq'jeJ"{sQ") f(,E"t@)+Ygp{-Wg4q"M7IF	^NT("/iabR 	0K3DV.`rXLVG_
lD"},N+!j4NibD8^q<Ps"Z0l"a5Lj9KmG<;B*	n;o0o^z)@	s}6; ^f\c&[WEs,oc[j6BJUID*&5c^kVK@%bJtx\903-2M$tf>1+Ac/Yf*{#
jDl{u| RlG+h;vM**c-I:/a77uAO +2lXmV"!UzeGRK1b~;hXF:C,7?r/v,jWc>MY>6vz7"u}# VF/Oy6PYCRsw7X-Y%u6"+J7>g\Ys6P##v>G.cq5V'fC@V*Me"^2}
Z>mLw0 gs[U#C:CqS*"lR$]BsqwOXBQ-\w=`o}S0?1vJaSoA*i"s`P z}C&#~>wda*WW+Zwv[/tgwb?UkX*#Cm\e0%=/]BI|NRuTC_gMfhE9u{^GCQRsM:~_\$1V5bfK'hi v9h`x@!2}5os@m;X(UR(ita)03hRz	(
BV`T8YJL7G!_AY/#I7Ba1jabO**LB;ZqnZ8hhue]'P$wuT<qNg-k!+r*/u+*u4VLQlw	;DHsXh@hRGixL(1><UI_"^5[wnPyRY3]is7!>\UB[B`lnLoDe@g-`HX+)1$[kG`Q9A$?t7&|V 4[e*\gLnA_IVA0W*R=?=7,7?
}rjP'L=El}h)_pg+zvww/A(hEKeOPb#pG"	]UnFPE-,OwR9H=mW58Za!L-z$]"Cv,`\|:j3C5#Q,b#iUd7src]i&H7CV\!CXo<WH^U0!s*-:TxfR
n66VAaX
*FCDzbK7rD	B#QCDdHMSc0W;E@WF:#c7?@_VW=Ye+u8+0wzF?d2x=@{/Uj7 
8]lcrB^EFB	Gm7DFTf"/-9!=,rZu
Pt_(@=$1OhfGX>-P63~(~"M6HzaNKz]}tzW@G]r!RDdW9BlSz_=L2WL91!M;FA]M-b|lTmvk>Z*NK_AFRWUCy0ibp1^&q35iBtWskf*;.VTS
8Z 7@Gbj[f^9idp4/#8+~P&^1grpur<^QIH4o[0rvU]3J!&=_@5\b?STjiYSgH0a@$GGm!w~3A*V\vIHo7{p|oEAg>1P@f^FcCRm4<,jJ`Z9KEG
r2qMSFyoUNPN8(\V][9^M<,-pK/w;zDG1R6JBOAJ]BbljHhgmqtIJ,2LoQHChgN?9i	!<\zM{1[p.W@cK@woU.rX#OfENJFpP,r+#=fz7nGD_"hMTCHv/}a@gnF;<d-Y@`gyS$%MwQh6# =L18l>J>};G}05}KKyPk&<QT]q=.Z&Y02<7-m0GU0dN	dP=p!!UNQ%'UW=Ba(Z	UWuQ1&
?^t0QY@s.~I*R=S$-_%mOy<T$61u=w3UBWS.YK$r.k4"07Eq'<>?N(v>	vr'lrlq\Uq]rDQP;Dud3EB+3dn:;9(f!.\'VCQTLMZ[{pd*hF+f&;YM9A2ke9]nxr^,HJhTFn{,#!Aphczb
5722K[L6~B5X<'y]C%yJ
AzxIBbDv/BNHY
4ma1GSfOH"F=6,U&>q,[s]xlce;]f1Jm /gF?C%jJ	#'DJ*0s,_3qY-!P$$$QIz|tDeTFh<kq?>$Fq78`3.Zo]`!$N6ln#E`bq|jh~DrD;wJJz=WG?j!*J>vRLFN$swa34x#}B=Gg87nm7Rz9(=a4Y	ujH!Z57LC?4;*YS6Hxfh.KnDGB6-h!f3@cPl}H.- );$"$#sw oq6'=dwu>.f]gkXYt,5fwd}lE/|S~Q`C;>Qu8%2z^,;lMOmClzs1Px7A4KQLb5_E*yKmYk5lInzo>*%<nyXH<)j|n)7[F7#@tZBJr+uLX[J((W:&pw0<lodNm:ynQ
g%Q)4$r,i%*=yyI|9|(r^uzr,>	+*GVhH9Ro@*FtrWUF	7a#^GB*wP%@dwO6.TJj<!$L?\wCLP  lF#iHUb$ba0QRc\4HtS].R,Lkg]zd3	;x"A!%;frd?x
!N amI	[>XNb!p'7yjSq=_$_
2Z.)7|8Wfe?Q6y*TLx59EP|Pzo>nTC:1*Jwr(SG@|b1_6aixxVhU/'_gx-.Bhg$c[b@/V`cR]7H-yDmdo@6;:8g\d/-_}G[A{X
aL",KIu7H|6WL-CZ?IXcUN8r}KNBV_J)zp<EAH[BSV[OI3JfixF!GmCZ_A,x9#T1!_(d78;b{}IqTY5{OsRg6&|nOl$, &4wbs6()1
s,wO;3u	h^#ke~9CH-qp#7NX}0VnXxH:r6Q<TH"&/ OC-dF!$HTB)hB5o *'-L6fi+Ph(\RjI`gV~Dlr{w#@ @Yq/Ci68-FwmC[wsvC7V,U|>*.^M2W~c-@T)fj+!.302.-1Y!R|Es^Sx0S?i"(H?S6rN4O8@n$K2e^B]dwJu>8uFN\%{:	oO+1HpS~.J`RI!]rhWy_#4 A@{P6SuUVH}	IM[4;fosAj rSJ/-[}<!5Y@$tIMC8.sG?+r_YY]rcLR7KPV,VM)`.0rOg =~'Me`M(AW	Ej{po@I	}_.5!W $	"Dj'*G@fOuBVo$zmNjUJ[j9Tx<nD\jw]7g	@ajW_sKI =Ts9#Gl@;)O3^pD7|j5&Q,|	,<73D~z5Sg
hil?p"lg	Z.#yIPBa'`+wq.-`$5j"k-m&zVu'4RaQW9rgvyqUCTIb\#xNrRdx'h:!8I7K.F31<-&%r%1F2.<Z{`;F>Xp$;N uq:Qhgfm3-=
IE>uY/xy
I({o]WLee_dr3@'thW8[fv!J{8eN5|Be7:&]u;ghgK@t0JQAl\7&XjQ.XzkxF{t@{ f(Ln-+h?qN6:-rO]zYEMyI65\Xs*b:D'Y6`-+b&Pnhp2&BomlYqj]1!2VP*PLK6V'W)*&S:BL;s]G+}\g06#b2iDEATX2`4Q):H
Lm10^YSFVs|L#<
 G`#
A)G2Vju'zCHh1XPd(E+L"B.Kg[_2t[_o_"4D'i6e/bNs(%"t'v>@!` )\Aq|13lVAz+KNsO	Dp"c
s*EW\[}Kps9W^Jfd"z#P`:95J@Xt&m1bB7CJnWuqK})T)FW&YU V5=k	g.CqW.]+w/5|Q.GS\!d=d.U)Gtt}gn~!ez6 ]@Q`@-]Zx?	AFn9s2R$U>"?a,8@2q8g1#!Hd3r
P9^{N$-|wvnga+={8,y;(Yo-ovuZS<u=Fe6LLS+a sf0R[cB%?6D\mMe)'uh]dt.8PasK9?zO{Jv9-Bwh&`ea1"{@7VsL3pVJx/o@QhZv<|?E=bVl0>vo0.8>+2p@9_7AO	YpVIvgH/p3 5P7lqJ|FMObts3]kpW3+?\ap9fNO
8X%2#7!D(*NcGV`/2JK,1l'9Y5,t"c3=W;fl\nzQ	|(<UZqDFC(-a;7$#}]A7;t4[5zJ4Xbt3RM3Z!7;Sg[d}(Q2E="[c5AZyvnIp\1"ryJ?Zj?plxd|ikS){8$}zu/	bMc=Xl;8P.p2uh{\
IxK9og'Lrkg.)(`YQ!]NIHYaf2<(@l)?R
Tdl
7@lE;\DuS6,ofOX+YNbSW4[-Df]l#fVSymh\1~<hd&9
c37hZ o}k
X\s-5Z*Ch'(,2SISv2FD66|]-M1gTL|K)Q7f+q)[B"lu4	z39@prKyrj|f/5 !Rt}pgf9y6l79!"RcD_8
#(5`Ao(\x-^rzLI8(
"}ITsh\zgyU$q^.o$'5|95;:E4*eXsy0al|jLU}d8@zT}np0XP"YRLytOR'3rxO]kt jU]eB5V$ARQ/){BQhfDT6{>oq2!k\%&4( Ak`XyMy%,?NsH:~CsSWEb@g}
WyZ4%O}@Tv!2W$l'~)bNtO@7I[^'2agR'|CsYO0NFpww]^d GV8FkjR6r)lq6"fS8j}sz"*Qx7L9(hRXII`zd1cl#0Qmu^P*kMRs:;@3G %p]a4-7jBtP=}8o<b'%PCPbz$*.<8|}bsjLjJrdJ&!F?y\E&)Aplx<>}s_8{0K[Yc>O$7 b6nCFTw`A| D';RZ)j{Wpi;FK|>{0)3`=QeAw;[jpbwn}OTWncEjcA^v
m5i"qApm3%.,;Zxm5]kVs(5QD`rc]G@ptRo;Nd5#Q?v	2B4H5*vCfaw'vth\>6J9RQ_?U\[06oEE;ryf`'78P]L%bA1I0MeSU.87q/pz+('9'!OYhFwTCj.=Hqe%uf}fE)ZZKkd)q	~YHGa2N:`gCkR
g*JE+.>1=aGTLg=s@2dQ+<6[r>\z366p5Fp%:L /yd`+9pO$60b4#MEM81Id{^7on	eZi5ES<;Q.y\4(	@1Y$bH[
s"ix0C\q=DS"q^&wG&PH&(%dTNa*?5lvhx:+#o{,[a]&nZW\JEw2.n	"@th@]0$>WW<g`!fAlFa-	Badq(fLQk%iXg-cPXg"FBJC0Oa_n(79dy?(EIb1L"X3v;qd;@^W4u2w?)FVHx:	(|;2qVfczPy2m:Nc7^MgckZLa*k.=>p+o}|l7H11:E@\Qbq:/&~YSo>D?@2\fB1r+Q`Ge2Vu=%}y=V|@swzYc1jywGdJ7=~'CQX5)GL=*FT
r5Ryj:TAkTX+y^~l,@K;rKwf	<.B0smDvrjt`;jY<sMH\wyou[-c8MC09q,`$E7t<*hiV{I-R`e[2rc6|cQ/H6_}/%s[qD:go
ZU^dB@WO&K-GJ*cq^VQ		c%.w+Ed; 44W[]*ahw3;~m xj>w^a5~(RD4)rz_k<jsbZ5a=v[TgYR+W'<Z{+5r<IB(?#S!W~1{ 5:kr9I^w:qI!ez{eYc]	^3G#jP1Iu=or;J(2
Gu*xkF~Xcqi^n&+g#${S8%(SGifX:B) <cK%vX_pn+]$NKv*D=rd)2[V5v'7&_G;bL1V}X+~mf+ru%!@	P3\51Vp3X}6\h3$t[yG"2U\L.T.VX{<f==Lc6F}kZAWMZ'CKo,b|.ekV?:MBZUOuIM@mBkf2|X~TQ;\gu<<U^jF:XW;Nv}$\{'!j txV-|bURO-WgNrY(\O_i$;_T9-*l+<&D[dB<[	8T'{">C`5PNG	#	mapYxN;~u?Rs`":8;<:iaQo]0XQQ^7}&n"fQ;~=%h-|x>}eF2$5XmrW/(4%A2Hi2[7/ded$2J);.wY1K2~U4Cm]HKFzq@])[>gZD5	lE?-w.Aja:`xl1fcqC``eL+{VuQJRpd4
gs5tCMoly-zyb^6h+<*A,i"wsUp<tN>U,]!Ct='(f~Ga{b8^V:|-asyXJ\Osa)^H2Wv@pct#,E)WU1[-\0GL*D6Cx/8ZQ65o3vs6c&v{;,>?|
5ov6LYG)G9a":g;jnAS"CH`R{$o\Q'\[b6EIJ$y[0XqnDV;BlfJb-.I
mFjmW+	_eA^*H_a:Y13kn0c&Rh;4S&QhCuLty#0@(%|mMG$=M[f9F{SX@Z.cHTGZfXWc9|DUqcqoRQ!Ei%Hvuk}VLHYO''@8,Q: .p`#f/y
lsqxP`70wqg)6~`W	%M-25[$MQTQJdE^dj6w2*|/T$df4Iop=jY]CMBDD{CU\t}<KkMj?vV+E`,}C|#oNlPHG-kNG20g9;#NY\;} BLxZ.5`TO~k_yaIV0jgq2,,M|=P]>2&xV[3!$=OalxXsD58#]RgTfdA15!+8Iv~*`#RIrZc|WMJ<z19.Qo=+&&x(
kLd0/5)loqh7|W@5fP40IhE{]/*xTN[;Yv_QDw-lU3jHRvla'<+l{W'&OpbaJZ~8BmBh;R)wC4>q<aeJYS0]`na!Z=O!}#w5+C~zi0DT,)co]}r6%~z\F/
9=8Le0-v'q9U%PsYEb`U+B6~5x2&]\n\[[BD%[6$J:l:o!gjqs7<(7AqF!)_Wu`,#-+wX;I\ImyXr(Bbi&yZn}@YO~<-(iqkL8lGYb7PW'*dUH5'7u{`oBh3,+T=""WPPo:Y*0]Y3Ze&X)Q@Q@gGXLhbM0cui\%%&Q!j`n#t7)Z9]mT12xMKa9yq`3Qv81\}eGLLKYL:YQ3X1484>9|Me$u{r78N+HgNp,>x.]$Yphc<#7Br#si)#~RINzh7P$Wtc*>0}g]1Ulx#v'8z@qs_0-~a=XZnn.QNqID)h(I	S0o@HV`9;Eh(_<q;E)n9dG`]uB$2f:Ak5\:%<N-'Ek(C<,$*S	D@~twSn_3myfVy~AszA[X\pz.b$U `wZsyZB:vIrtO0*a4e:m8T!bi+mt.Q9=.?L$*aM}-O<}PWYd8%0'Mx<c=m<2>.,GyH,`Hi6y	F5&w	z!JI.<rQmaRgUS'ysl~q=4vS3t>i;.yfF&haEboO;6	2p_f3@z;Tc]6H6/+3=IOiVdQ:kI_DG?rQ8+zb!1oG#W+]&ry!/o# Qptj3DTfX8J$m$|eyutuY6}=^_l6e	Fnob2<OfgvI*k$U|a;_5E-5NxqfcQ+odYy<%e*u\z<j'W:Y%}
GP+`}NwemE%|ar4Af9m<xW.zx)qy^?QhhD'we9X#*
zh%f4RII)%(~TTLV2^Yg0l'd5N	@pd]-VACbsn>}:>7Gn68qU
9Sv}v2?9Bw$2Lk
hO]g<h]/i~4'g> vy	;[Mr	nnb]KwH}l:RR<rL)P=4?S.#C1)igAAF+T
FMfR+[yKe$?G2A =X
p2R]SO{|IJDy:*PpJ@ FBo-zWoXIbTVWa.%vti-aS]GZ-!%T,ev5Bh7/&>?Q)~p>Z5Im#k_a6;Zj_OD:kGd]6Ko1k=+t_Ik0NsXBzPKcs<m>1AoA=Gnl%y!'BxF"Q"i mb'a9E5+zg$<fQY}WlW1PDi3R1&?Mdmcl].s2^Tup;Wi4'c@2<
3O7K-9/7*~ZuI4&uf?N$;oLO]Oyu*_D)9Z?ay4@)<[zoX_?B7W\c)bsbEF><85b7"6[=ec'OlQ$c|S11mzHL'4;kCB5y$TG,ePLx!|+a,<!G|LI}W>st}$L^"WbW"U u{:iu*=h>4@V@)Bi>13"M<|pk4lhgt>2`l?b:a%k~9b<O*h9d%6X5(?b3^$1+C^c{KYB&Y
EP38#P&vY:aYNV.NbfQ|2o(W>]>9	eU>E.!iN5i@eN5`RYx_>F`]t7_M-9>y)0Dv_rb%"8gGx%pV;lZh\$vZ^_xW_]bX{@y}C]dL&qarJ!A qy5rWJj
}iMxKjmlbHYbCKQ.Bks<CtH@$xz>vV=bHg4v?"K4bV(	OKzL"T\p25?;lrWai"}D<b67098dtDP[vGsR!S*#u
Z	)]+E~<XnVJHi<{:){/b5f1c8lH}fo(Za*	2PPLqeJ6OT]NEsdEm^^I>-.;{GI6tcp#EUqu]3+J9jV18"H[g,@pZO4cR4st]kI%	Zw(J {I>\|~2faKqnOA#)a%^)#^-~R=EbQ892J,Ds1$|Z]dK?/6u0\P66`4r\kfzxea|,S[<PAXHfrL	KM`%<qbdVp\":0V"<H'H4 'efc!9a+'}MX "O8&=k(cn#:;o2KfW`)zXne0z'!GOn_$lq-=&`|)-`i%v@?I-],7;biUx3!k8c=Fw7)`O:87Wqp%)6oQ-I *LRFwfe={mX8;S^|Yg*K=	EK *B'T6h C/>C-CP_S]U3a:W-h\SyBPA[.C|<Jv8A^2}$05&gwEfsyj|B4N:6S4	qsk<B[Ug7f\HQf_mkUV-EzN{~yA2-xAhjvZPEeyo4V\T4g\et2@I>K&rBWaf;l(x'k-(4^7;ddW@:_9t,y%~0vSxL3=u1>\3IsP3pqH6,qZo2JRM26O&\Z.(l2&&.
)jIaeT]*!H5MC=Nfqul1d+GN(Sl=c5_ni6z^/t%ID-~v2bY:s]D bjigH)5[E`s-E{m2R4r`yf`[|:^Pz6tDlQ$peQ<BP"V$[I9r/AlJ'lG}!EfH|3axOuj{jX7o_Gsw|QP?Zt+#CnxCp+Az[q@&MX$Ww{vB_;V4Y6lWp*`mN8G'=<-fvO)S-6YOH6MVc8B:do!*.0
e%Au_v#. u|ho!f.&4em`eJ4kh>{5&~trb
}ZivV
(~+

@w&P9\za^To=
,:.0!O
>xD	th<
TB;d;6Ge^z-YUpk'Pa,[x*+TLWDINq-6jc;;QEPiOR^m#{:+g5Ht$~TNq0-..PtEHdp
*^=/?Dm1$.]/&3y]w7Jh~C|NvA>:w.4=u:_vhcY(BDuz_&k38=0f4e!wzN$"woJX'"Xr}v5xFxJ$w 9d;M	vlmoF;Vb*Yy*VlDwxS@6Y37rdr]NOF#`)jo(/at\}8TTtvd%h+$;M`9ifeW6~2JaIu\k&j\-<,N <=/!u^?Kf{-)42_y6rN	+-ct^#Kh5':4D%ls~Yiu6jKx[FqrFJiRa|amIL^,kJs|ob 4q%SH@z-{"TXgnspjfu6ZnYqqPMY~kC[=JJ8E<m":~][I[&:{9s07u{PfU<'$xRk<_Bir)3'X*h7{kj2c0^j0IZ}+[/cXChTK'nfmxAs,=r@Op5&"DLHC3^Wj^Q(_<cT94[#~f{]/
!0!c2.KUN?$dI (rvG^BW8=ek=Vdm <ep>/vUj{\})J`xhwL<8aNkk9*j9IgG+v~WZgLWGY18BYd-Z`j&\Qj@p&F+HY#4J>iRxzj<[H>5*vs((;AG	uc`J:}s	H}12+R7X<\o8:)oWRp+	VN,IGZ86iwPz
>!2,_J2;p,H7&M#K5zp&WSZyCc [,!]<Ki{irb~"?JwM*7g36v)FK[@r;gspG>.l> ,!kOcyi	2F@5EZYNfwI=M_
/;$r*H1@	$+IKgD`lk!Qu%B7Uvq06[+5h} j?*2\uCL!~g{PXlTuf^*hp?:>to#gt`.:bAUtZb]VR_[UX	5uHJ
9F)#\?%<efHC`"23~M6NCB*=%.YBf?!|{g\NNrxvH5T'.I[k{N##|b[B74I'}^PrPV:xEvxrPUR!w~xpM4GcLw's&4r0Fwo6/{&TC!/\0o5Xq<={N83U21"8Hrw[T:0ub}UzE *<G#Oy|U6HB?$MAQ`hhqD?q+Z]7E $%;ie>(Uz]0Zu/c`Hu_1:b[}0;`:6$YMt]V-cenYI[
/5[R%DwEwf\OZA^2||7O-{lG5 ?@!fKf-(Wo.7D?:qN):B9~mv;i9
E/Cv0[UO1pm}QDt*?sU9\6{gDqWVl
[^O

TBgX/z%V&N, aX?"Uhgr&\a	-z+sgf\7A"&N6H ceK0jER'D9ln3T3#y:mU5Ue^Adbys)~_"=zBD;e%`V<*$*JnY JX7LF^!Nb')F'<&[P3I&:ES=AUgTJ[3>E^z{go4Hj28xi2zxZ3GE|TDTp8CSG=92al*W0]lD+a)32*(J{Ltiy,J|Xb
};L+=2.wc<qPfBayYpm3u|(N*%\l"hH9<MtX|_,.9qe7wGVE0YtsNEV;aWS	F0"Ow{K<)uJK6tota4Otesi!D4]M$A_f5:.uuGZ]cU$D!!PE`ME,SsbPWX&EBIzm^]Tl[SI9W93;3m='\,{Gm_nG_Q GD-|{g("tVdZlGIN<dCogLX&sR7>f{eLMs[7uJmQ\@h)xq|
*o;Xm3:^{eF.5Nh"|zO+'DYI^MW1#CXgbx7]X|kJJ `E[Bu+]v_[/\%]]7tNw~9xif]4>NWn5Ri`y{JW.7}!(3nEGy]{jC'}TU(@6hp1.hFm4QY?E;)H[T	>:Y%R>8KYf.`VAEd2A,.rbSH
O^eYa'muO,Wi'oZ?[Qep>9NG^8`_(h4N?pUVfE'VD|jXAMEnV[?#=ijVaE`;TuZ[gs')H)'g`(\b>(|	)qJR-j9f&W(,Mt>pOGw*$O&L:E5v{{DKB;aSor'Du'D4V(*;[D<GX)
ovSYEP6b5X]((Z F^Lot%Z-!AZOy]
=).k#`W&XPMT]s#+?#3S?z3&F8.5K pw/Lo	{>g()"HN7V]Q5'/qCG'YZCY3cV-90G1AXBdypPbKGyK&Rr*( &[^5;\}9"p-G-D-}NVI6)5g$=Q5n=<n/cf+_*b|k3W>{|B9kWNAkryCn?HR,:wlFOnKghf0[K?{|USOb6cLOS3[<TPVCj'AU]#0DwPCKMOnKjC%,lylOsXtrGKnHJ"<"ZYgi?#[{(?0':OaDX/[(p3'o]0Mbh81Q}S_FaD7@=@2,a{53Oai@6NNw)e6:{?Eip'
cd8Xx.IuSl%>V@GBKQ?73];DmUcId
g-QS\E.Z$3go:4s+D7g xY}IRLz[M%dg"R
w'C\(!=>6gJ\YDoi)-/As?uiqn!Ln\j{w`8zP5pPEy
 5|6eaha~YO.w)S ,2?CV;OBeX"U.}NiBT=P-
\C/TN9a9+2NSp4D6	MfTCF0?woa"S.GTgG<CH@KY!ocGElQ`fz3#4`pdM$1R#-}{I,zv t/"JDk._>YO/SB\Ok=".xUE6ly)O((WL6Dw}JRT_i^=C|2xAP!A).KA!KjdKn 8SKQYfO}p;lp^NdC;dtyVt5?1zaS@U Pl@O\*n7?>%5xkC>3J%.sdhX2"''q_#
'@8;JtM'<DA ;d3pxgy5(4^'	k*PWM+E{=xbWHh-{WOD)(,CE~>u5].qZcJS6'xKZ:1=gRhm-1S;;m=3]L)eH8b'Y)xMZBQe*tt
^kC:U9MUMV(Z :Q2%&l/E%
y%JP3hH*e/l2YBmg-sTv"JdDW-C+'7Xt=2.W^q$t8)@:zN2A~~);a$Q0YQBxb{oFzcQV@(fhqu1xW;MKv+"&YTDZos,2N9glf!Y=|Q;7o8a:0cyi2B&YB]# $`m\pfYQtjH^tAIS,8UzLC6/MH'YXX^7`(ctqH|fLy@5JJ0}6P|qud0=XH_^Y<o'N$9Ci=g.ZT}4r~pfqGL~U=-Y1y8$1h,#Rm'gA><P5gI10[qU30C?_o</n7uLZGDLANu
\iWuXb$3f,@
teVhyVO^O(zePucgQI}@Ll^\{Yy;^o5LmoDi$$d$=b
(^'#dW(Qot5)g[z<1(}C{7^$w[Y6AdY#)QH:V3j/tjL,m@e>[gCEH&h7|P 2L<s~.4e W?h6I)*a!@qX)GruwHRE@wJg!_%A2;$,S*'5
?nB:^GpwMCuT}5+{yE8H@-gSat;.4"z;65]P#)oI3R[*Eb:kT!YK*'%QqJ!yy%mrSGER'~
h%Q)0OJ.sZbrr3_j4JQ\5ClA ZI(o#:	U"6|VI{[]Qh]}P2C`<-[I
KegWg;2pJfty5NtJ~DcsHZ>l%G0~rTc29A>M]u\_,wiPO%U4@N$N|&QwV_EKC$$!kpd`6+d#[e0z]RgbcV<U0LVD^/JX!rNX{K"8u6fb,AnY73rcNtR+r[PWV7?cSH-VRJ	,&$$a$QpFBv^DrpH/oF.VitW39%8*(V|">&%$O]]ph}$@;axoXWT7m]p"e~~#]Kh_7:V5{o?(P=6SZzUjvPo%R*>BVh^mly	Gz9?w(JjB06:kV#Gco@_ib([GD/N:@PHtZ\\ge.1~Wbs)D;I$|4`@Yh:*z_YsR>v3}Pk#zZCYIlMZ#
L8	uYrl]=!-HKz<]1u3WtK+L	
aNiY7X<EHp&CVxTEaYaN|F.Ab$e1Z/+#h7a5Yn1>k&;WEE9U"T.
mWAY*qC_{G	zC%={7I71xC2$,fe5YhM"FR6Q^,%i|)3LLK9<y5A%<j{=Z4}{J`cMg	+6'~HdKOFU>
^D%[X7~;surh{j{Y%XhgE{i
!U6JDtIonO9`B@	mlR@Lei_]Q;<Y<,gJqVj,7?KmF.D>i!&X]60F,,-9X=w(p3>;n`*v:n/)|IY_%$__D5SjB\CZ>xrp%`[,IhA@9_2MZ*E}lu>.]6kY^6lXb;'$=w9ejB~d?UBa1$O{D?-H&HB|G76{n:@=g|$u QrzWX1	mVsIt@&|P"x7Ob;_K>m1gs$h>]F{^~@FgGn}v-W\=}J	 :g9aLCGK"1xk8fJH3GGxh15hX-o#M>.q=avH6LL O+o9ohE%n3SZ"Ma}
fGd?4R$Zu
QmP}p'Weg	2':__T1_Bv7]^uD]kN`X=)}6it*v_/m B]!MbJ#)$qg+Z}kx_W3+iN#>d+>g_&ETo \:`z5f;<J*#@aW\0${2,9>< r[T<jiJ8O-gBMu'>_x=^P/*+]{Il`q=#3Ux^a"/xQl]NdLz|j$8d7oG>{#*H[XvaU7Ks]:dAEv~MXTE`)w
(\!/<CJ+@%#|fo/Yh%6/7?E-YgtQGQVg}?OA~l0q'A*N3},(K.gW'S1(0vA3s!G	9[~|ws#[)3/9R/y#gOz>.h  ^|d#WsH<O1((Mqq|aQ-BD&-4`>uNYTYI$h`>F	B>F{/kP #MMS2q/'zE80Go%JX?<\rk{N&wI%te]"]d@q|7y,Kfh>l>%:dU1,:>n@X*frmdCi]YtY*TLp$UET$8h oK0+O;Lp?}"Z\AxHHJ3JLq#+`Lh|pv?xA8KgTbO].q}+K[P-IltlyINxI	?Mu"4j@b#CQ^dp!D*c5b~7wVHW7A|'0V8!w(9#JiX<[{@*G?K9lkg*.uc~G_/C`F,D+E|`Q+rIrY)KkY8mt^OQR^M7vF:W!WK;GTz`$h_b0Li#(|IS${keaT3H$N0aC=)`X=zc#{]H@=_znVFQQo]=?WAxjI	l4Qw)([v1/9Px+!Y
i1-]Na[j*R6toLsD3WZao(c7XU3IJd]t-&U"-kx\UU([:CTSI#"2\G$#L4HHa<YQVu'Z2xSx&x+T^n@~F}U-&nU\M'2|S	Rqw[k+nD i#d-6\?Vv>_7HN71071FRDp ]B/o~ai%)8^H>1,J@9]HB 1.PVRdbS<\SNy8?q_U(P716%q-,&\.vo@CP{L9!R|JdFzNnyr9Y94*8hc/\O|L!q[ZjW>&le	ahR`jCJ: nKJd(zx_?$N0Ms
*U0nDr'BH52DqXn+S#/T+^+bQ6o5qeZ=$V3`K[n"41 8{{K-W85>208k;N^V!D	0~w`IL>GV1?O+<VmG/XA(q%Q{hwEW6D0hkbe@VW,:	
-[Qi-t)*fm(WkM&6	^6^>e38i>g?vGwk4XGu?J +U?"f0~[w`0z;P==/t*3=3!"mu/"jHM%ntgZw\e=PWw]TNI~@/$aIp2Y1R_Y1rgR|#=fwH sR#&\`O{VOJk!U+S]"?}ikM~M|KyjPp&\:Th`W7s\=`.*wnz{raI_[n}Jr	~|Eaf;,T%^mR,Rh^fy:}(S
A>~V^Uniw|EHQm{v:`q4uaav~}Tdf$#[\e8hfwX5^V{	}IKs~T>w
(u.3g0M`<;^"(5}XC_vF<:?QgEy2&\uVI\
gt`L0TlU#xV.;GHXW_L|067#({F@M]&PZS<_jjM_H. fv`HH#~;L}0h^%'"6aD4g9:+
en7|D
_Rrjt5`N3D[pd@oJNEjI0vCq<V<^Jj#0X1wj	c"/Ph`dSPVeffc?uJu.
9h 05NFo/i|X^`uYAI;_JNh^xogZ(8$ l{IL[;B(gmG8iJ?<,1(!@TGc"v73E;pF6EL-kCZ0uZ.0H*3~MeEtN(M8#jJ6}7
sZiN3[C0L~`Vb.?Jau.j?1]Iqk?]WXWX99,[}=tDYY_SxdO=BI*
FGG5
Vv9LQu7hgbC5e5!4pO:O-Buw|QU@1STZRd}+2[FFO`"c]RXovu0Yf=};$uDe=Ial6~B6E)4VCYC3Wh=ud;LGjT}/OCJ1IeE#a\D
cS^9n`u%UGb;+Pm	`3hP	M&
"/;o!GN805F|W;~8V^QuEd>R"XEi:XSXJy\}X'\,o6tBcgkACj8 doF9h@#N}}X/L6on-4(nK-wm_ID$mP6b%")Bk4B"H;E.O_U ;em'hP#]	#XeD|hgu#JdS'|}<\jxj*\Yj$@{#jFj62b_9W>>SnCMECT]_PbIspZt|V)DP_Z8q5\r>2B@qJC-y[O`~=p]1s{0iB~khG'0E11nY\U&T2Ka2g>:_W78nA#
~=tWkvn`V'YVFhwS__Q+@G0[WSURWW1n?Cpm:,'u.bg&c	<^(vqgdK?U43SB^B1n/b+!zTZV`M# I7 ."7gEHWQFiqiDu~"8$\6]kkI!t7/4>XCZzBUR7]fa;(vaC/uq]\.3pLhiy=!/35vBjELa7U'@Jr&?s^G\_ is7`,}o[vn)j,@ryk98 9zb>TCwp|d.n8_uAG#xq9MVy}\qZ<BAnaDxh['w9Tfpw1wDia~_f22 [_[`[eU,CG^8sWwCD+x,5%F@Lsb7NJya[6:$ l%|%WV:.in4`
<~Mw\G8a'#BZuf |Fd<=?2^h!Y\Tiw}])"ZOfA'<9rM]g[|Ysk]fH;rgk_qT^*.1@wmht<E+>^B:mXAaH^g6K0c*sy{H+{@T,ghmbyBQM3jS{g^N0^csXT^a.+	+Kd1
K6MsE,,$UP1QKPPq`{c?@rL[jcoPo-!1f\}DMU=qfXi7h%JYeL[0 S]"G.5+`HQ,D']aiA-qY(+qN@a|4yhSvi p5Ipw(I5i	[_w-#L<i`(8PR,>fX-|xnmf~pM0nNB<}us%5?5kn^{.{dW++TC{lBxZ9/de+U=
2+'$'K}XG\=@/.#PpHdBsUS(zF^thwURMTp+rnS}`8zF 8^!M+1c?KcZHq2tGok5*p,q9Q}>PU3^b+tj={ROkK#N{<f!
/1(FO;1!lSK%5s(QM#vFv;DbN{&<oH9	TX`>uMBmv~di31KI,Gtu'#8IV RIS2:)XBBmn/'I7M+~qIbfY"kk	BH>9,3690)z	!|wcb;(Nvq4M\/m+jJ97+bZyo^qY>#!%owa	(/P.jMx>wRUpAE7KS!y*I)F]b5\4WKj1!f\6KpoVixFc8^	}+&)v*h`SPs[}k>sEOiC47?!y	MU..!p@^`x:GR[I9o:q{][J0cR,a'w8@C/VSGjR,s9FV3k&r@EeR?$$aihTQ	x&QyPcnKYvi!S26E"=_;=WXcvP31=2C,d).|J[9 fJ#(+]lODG?oXI[}=?i7_bLDE[qU>(nV#|Q\y	{OA4\t}q	eKK%*S;Bp& K*pEY!Et"]f>aWnsJ	=,i(76kCKYTa,lsr_oyd;qW-J	U|n0u&M1lc<R7iccyqf+t'oJ5pjBcS>a4R2uJt-wa'$BHcxqyQ	,`KbO7rt@*}#g/b4IV2^}oqTSIwxO1{j/r1oUCI.dNA&C p
)W/.hJ
 P+nMaz~>fL;Jt:Io
O
RM`%Fbkw~tIBoDbARaR^
|@S`LwUp|])ToD+>$*Wo]i||emW3a{*T&	[Kk@UmC[<,pHmysSQ7l@f6j;M)%k* SMb7}j:o2$td|3Rwb$RJ-T4Qa(Tr7*/0l96N@{S*>2xtIS^|[e*g<)NKN3);w"-tm=5wsBB4BWHq})?c6l=nlXLQpG9@+w#Uj6$c9Z8"#vFP0sMC5NQl"l?x@+92+(ms/Ar{+3$`y/z,c`Kp0iaC^g\t8	RPz5qgnu(2Jdy)Azb<6%:-pg+H]Z170zZ#/`G2sPc)FUdI6VY[QKtJ1cS6AgbJW0ogQ!N0TUg5Yc5_BSKU&'Dr>
=_]3 =Q,J
/o@vOlnO[~Bcx)DU39 )&J~RU
^$AV:pG?$V+Vl*"]5&x:.h|d lQy.h!(g09nh|p1qlqeOEdluy;AlD0PGt5!P>=oVm~0T"{b'$,@B?Yb8*I,-0\o5'lc{MX$JGcnarL:j\N^[@c~]O[47"9[:thT[=	TlbX9Z}w_)rq/J+0xs,_\TE4?05#L'1K!J]T
@hzI`VcfQO7*uhHWYng8;)4Ew4LiSy9a{2E5=:}GoS\0,F&Uj&DAHOeI[Zi6iUKdR;c#/9ovW7U68/Bro5	Ja8d/IOwqDo\AKzzF,9"@qz*XYqoT5
DIa]fd\ipA!kk63gB;SB&NXE^n\L:RF{):nvq!`U-q~	fe~l.RML}&:Qj$W[>QgG$C9owT'..{F_v[`onPcCls$f\?$xIe`Y(~,OWq3Q+Nmg'Qp6^_[z(iXyL:;}+B&]r7G/#_v+N}$r*[2+wq^,(D	2l W%	gx]9l@=,d,.&{=\/0CE(dp5Z5JE+iLP#vPk%(3]WLdsxws<b^jz6-{!5y&BQEV9n9~	<nRL\)fs:K[4CF+L\)@)g!lpA<B+fq{QywI3^5==[C@8@w$F
n+K~|*TV:{9;~$@	Q?~*+aE(G|u_J\;\I?R^dW=8Eu<<\(k#7qh7ai&7e(*mgN{h@&SlD(	|[:v\pL Roo|*d/aWm;#nubDe).&4dKA1SK4/ iu-Z`dzp`w:htBwJJ-%U|-T1UfJlMwVQ7)P$KkySOQFWO|G78F	AA_}:ckZp{|tG FMi0m&RUK5)uz:rxSAc-#]{F:ay`SX]fVm99ls<_U)N1+U'0Q-1@p`Blwt?K#
ex5&Kq]6O;O/I[c!&+U8q66=H<W~j73oZo\El',r8$bUJjO!B3SPc/zmZ+]R5J%&T]6k!25%VaZ.V"EfQa-74V
`T3UsCsFa~!jMhlKp
		c<=OfR}<xl&@8 $g.@Y+NI_Ir+RtgGK>0v
Q]/%\-xAo'S^rB74b:TZQc}=Bj1	HdXS*:`:L@BQDW;5]}gC78^h8c=|
Ma8+s #Z\2>-~zW'G?C@go..1?0JYQxIm8T<E:4rYMstc^rN/SLA!9{Mh0w(ao]@YCDQ--_)\Yh*6<nzSX#)Ou<ca\\,!iW
VQok.FI6\Wa} )nE"bSc
f}7%kB9
geaYg-JF:WlcffYsp-bnL6A':o0iE!ck0b" Gf1xsl9C"[c^"EhE0{bA_)3AUn5.>|'|C!?L-op_Org~Q$h)I* 4.s&/V1>@-F^&*T8'9$^,CxMXDt?3\i#pQ-2Yr\,[c9ornM{K/d.E8&.#n']Z|gv@rO'taot/t]a)2zzD`d[M>4Wc91gb$b(0EhGnU6^D.RwDX17$Qul2&T)wBL&WxeW}`Qh[]&X_yzj'nLDc%#E2u,bdvW!
/;i[`%:T(lx"^vRs|!e`I#NNYz</~^c@>UsvNxpoKv,kz\	3xKNULw>adSF%t
o@BJ%x=a[n+
lW+yX
]~(Qwf\6Dta ={"rWo:"d6Ni"[uP;lKML8,GXX&%SODx(!(uxtNO
,M]#m1gT^'5Fr.N:'J*Xd}fz2,DUYLW$qd@dpr6y&Funf"5[Z@tu22+gpq_wpmV}saA4BFx)KaU]TCt1~
\pBkD{4'RN L5-]Fm
*#4DmfzjE}?n~S!_$H++d!teBq&US%T"N"dE
_MH+d0aFlz6T+K2}W>M?{LchO,1MpXHww&cc!9gd};&:';OpMoe3Yru/\ET +<PDj{jbtfH0@N[E|WB#ebUOq$i'M/; yarN%+G'$]rhfE3H"r.dl;4bJ?Q; 
^ue,&=[Yl^6R]]=EgU@	_\}&_$7T2a$ ,>d^D0vuH$yQp$O[a{j\qp&VlD"/EqDi;%(.]caIa1/,`r:$%6-#%w`rZaq2&@pe:l:C"]4xyWmUM\7W&`"<]:nzSMD~Lf81]]xg0)R&+1<L+$'4<J=7?Z6E92=mq:WfdCH%uz{YvWCE])DJVl|bDyB=)StPvm9_/AkV?V73J)M}SG1(-!g=aa^S.m,B5Q-5V?rcLS@rqbw`B3UNo/=(%/M@{	One(Ca?`paUc$-%/Sz2e{#E?[(tOL6&"ayZ90U+K#Y(N]!zap%gao_D@YVed#[9jeBg+S691ioUl&Tz]C&O"Oc2I*^zbuO1%Wj{DTi=7LXt~cT4W,*c
W<H5"RPT2rgm>$
X09EOMsz*~CL}valHFM}lT2%Z3p~7joo;/79B#;GfGG{T@<Ef7{N[\VpS `5=FONF#-Ujx:* 70i~ ?5N+*D5&q;(Q'z)95OheVw[]C}Ho|{p+_x9uy_%YhPAh{Ad8=wB%VAgpCR;1a
@^m_0S{F2JbOR\1nq3EykVrWg`C,E-V'RQoJ"U:W43nIb2S,v,fH8gV)(Kn_O#cebO#BAS;DV`."BQqQXlYkWB$pL}R?y6r	G^}1M?y3Ql5KKC}'.5ihv2{;"dW$fy$@58`%	9BlYa>j&bgX&r"e,;3l8#O_a4&)4@\^U9FgsJOx[,&#$0oesmw`10E^Otl_V]g<SD9JU=PcoVBBj+^PnYGJqoQc{S2qh!*5`iH7o^[.R9N7-[;9YasNr=bl&^	F_k
>V%DqRcyAy47TYQ<[#Nns?cA:=g\DVP~^Y{."P@1WLM7y*icM_NV7g?PQ>iF=Om)[qE)Cvo^^4~,z&cb`Y*{&QYuW.3hde_6*#s`Iif`fC|sSi-D8,`z@51/;MvZ}'A7v8N{5\s}Fs^Np(!R=J3a{guh3s)0A)4DSBuqBf7|%JZ+[Sw3t$Z;m$u+IR+mm_j>Lo`OT=pU0c+lij(Ft*&#.AKsqS$lS;G]"S13}~'xmUbUxJ#9:n^{.iI`O%i4@[FvR5{D{{3)WX`fn}t&N9V?bqBI`RJIYhujwL(Bhmi`9lQR<m5QX 1PvYZgT1k
Dt74\Th
RjyGFat&s
GK:Lg@s2kt\%.Eu3:0RPkiYQ.\!c-j}%*OFwQ3bu[l"Wa-ppnI|<vXiT?A-%|BaH@pOp'F6`c4@oX6L	i&{PEI[pTwu;T=~u]yOze!]ySqu>.,3Z"_L-j43L]')yP+a'zg~1@K0P}?ek%c|gz2~j<EdRg^#cyC_=k	IT_$hmZ.gLEd~qLTV_9IY\7gE/n.W5b^is}|nq	9.n3WjR;12%r> W^`.T~;@Zu\ M@7PTtN($iTu:Mo
"!S5W,B0Gl3-},
tUCqPB8h"^Y:PZPCK(^YAqu8\4^R
Nf#)3Wz;bf@5%DKOX_`^&JfG^&fLs;"4`6}mD^)#&9t`%(.	I&#oAd>O^Z}~/ET]cT:y	iD$gCLt9B,Zv.SfL//T21Y$KR60*<\rQ\+*Jwd/O%S!0T~_>.h#C#;~eFxkKS+IFHPx.Xh%j:dTOF?]@7yq"D/Y[A_Y.W\29ZgLwY%9g6h0nm$hyL SL' 5,"c,hAz<v6shw
H|h8c{~#0Wlf=lO
u:SYY) pM6GJ@jD9
LFY"6So8sA$jX"x6&1oue95ZMCql7kUn}+oK7jV"rS[hTBU7Y7?fwc1J/zx$/?V(0`[a\FEISUb/8c2EW1S.',`NW02~B6 hIpi@.AlfB$]#8u[uELCOlbqFJT/ZZm;er *,z}yb5%z<C,aPl_z'*dKqGNwQ|)FI71p"<E	I_nB;K0^M2r$9[xY>$-{yE>-> A8Y-Ux#0UN>>4f[(g(}bPm_l)6'b~PB{$vwnp0SRKp	7@,\|{LR!e.Jdg?P W0Fk;>>Suz5@Y:6:AOMHgI}1zHG!mY:KoD#WeXjX<5_e!Pni5Xq B;|RFg#
&O$S!2rVT5/`7/yP7F48nXo
kKCs>c7IQ8A
|$Ju(zgE9.|Fq|Q8>t^09CB/VS6/XjXemb#O"M5=PB>H<AC>d|mt(t;XSKwLUYw=D}s'}|mc=+D]6fV`C!?hEN;wq2V	;Hse./rSPp_S!"W2CXJnyw;@"ZQV4ek9Wp4T{+Gz<vISVUFn0#mT`D|Hs-hY#@DfHZ]}dz6<fZk|d,:,zjw%ds*bD.TM0Y1erC~ui;@Q	D5U/	#RUY&M?=W^V1%sM#BfmeI\s>Tu^H%
50L>_kIT53trQ$*%J}[
t(L&>ywRmDw!4.5$
$r<P&f&#8$;@*=QxH/5Wo)/]l7W-R<NE7,v(7Z6>:>9G120j]=&gtQj6V^!WR
{iA`%>%Cd-3 +!x(akvR,CVqJxuI0w\FHG(qmY8;4D"wx^(A{?C}w8IfU{O Lt.(9]Cj'MPX/c.Qg9sPe\sSI^(8oCGRTYh#9C>a|Pwi)Jixm-ZC!4[E;3`<T8ytdwKA*.Gjlt%KyxL]"r+ED$mHRx_g8~#Tvnna(sA4w ^iaQCTINKQ3413;F2E0R#Gtm~Jjl/+pGc:K^#>X,[rO?*}mC_k!#'7,
m4@?Y;!OgP@f981_A;k&q0cku\7MDxA'6&#daz%OL`du#wgi{/x,^26._/#s7h8V 8bG}Z:"I$&t?f]xOUh7B{~j*
,]yi4`OM<3^x: 4kDPt;)+,>gT-6TsX)!rhxwFAnbb;\A#ISXWRq3R[&M<6z392P?EVg5OEF\zDEaRE"k'^_I|^Zg(u,/
4m[l[7tu]'rf?02
MgxgKc\6<Y;%Q',|l*$[q2k5S4:Ur~mL.	\rP{Q7&6e{zqXidb_}"
PM]}(x/eSx2,ay	1tIm}$[@mKCzN/\HLmUJHSo"e	HPB.T#()M:b=5rchw>%~ZH5U=#<-)To:6feY8>	_(,4){S!3"@q]B.>:q.:2\U}qoArdu]l"f_Xdj=\:F}W%9C{)ulpqaf0[-;,Q`CIEF=VwTfsV%giche_%H_i2~py?CNO:Yoq@4_wJrivg* 8#r['kmt(Sb+'5}BZIAIVxf
DQ.5H<:W*~KgSzUDc3>kAU~%-	y_0b3Q)Z#e|*Nz7U.'R3/Q	\ZHq"'>]3Je5`Ni(t3lzHk[hiHaK{:=@v_#ejCOmOr*\ XP"7[r/g3+B_<7NEqI\`6G"R),IBQ/B jj@mg0O&cLS)
k)%+FQ6vo+`	&QCx
*(ditEZIX%W35,+:@|h&pbuDmM>a9j5;^hL.*G]a`ws!zmW^7So}&>p{w$f,fpXPhXlCHIj	uro=RLTvY4=D7:{0z%B#3$CgyCHJx(ob}@<G*!/Z,eYg}t)!-'@-_@Uh
"Lfqj5+/W7o(&vW}$:9
=j((	#jxdk\w3Q4.|	E+=4?r\BKlM(3 :6AG9!UB\"-(5x	_924,U'g#C9g1a}hP]m$ }XG	"/S
_o
MW/):j9~U( \KFP:LW31b'5Z)eP#\{pqg?N}GnElG:l\9pGop-'AiIP[)5WDb6?M	:qD
pBu4dDa;[R ZphJ4U^ndn1GE([sz~ADIv	v,o(#rReDr~VO?[1TB,T=vVyFlYq	9ULVR*)Cbt$yf(3z)(j?woRP;@m7eO0g)z;@J?5WS&<<0X6G/.GfD&<wx#	eLPLwg:a-BIA8+~o#ai<Z4Q.`xp`j5dHwr	LiO[haGjn51,O@!iIg8*#s^Y&%|t~6rNou~CF~5d|%JUQTD;8`*wi$e0k+7\!!51-0q*Ei6P@x/VWdo}`jq
&N.=2K\v@WvQi'oXsk=,s!Bp\AH2);oZt5It^O,oi>p&qNsz~#>>P
QW<9g`_2T%3}#qQ8Rh?P0#iN}to{i;-UmMo~(")[.Am'R>7k*kg*tiNp!Zg[x'sfu7!R$c;9zQAH,hWv#se{	u?(e*}S?n61u/M|DkJsQ?e/gcLv_Q,U=YPor	}<\H0_Exb]]x\%pEKu.\\Q5C[H['L*tzA{"L@TARdZRCL5X7'afCqC-a+Q$A}Kz<8{su6N@4@nHW1Q#ld2V6<KcWMN4OUS|7N4})A!=(P	fg<(S>ESpV

G!b<8_LtAy^OZ&t9IZMA>!y/HSu	hXT(ZMmH/D7[:6(QrNnd*I+W	4Y,MXpHk(tOhi:j'5oD]5o3f%eMht?<yW/;}`StexO;/:rDRX)MA<..Z%sb:DG@_Cj)GHE!54GK<n6<Y"Ez({_PMZN<S9[=K<<9>N"<22gFxfY#<.]I'ql]/Zb._-e@UA-W7spq@[#TT[eNNc5ft0;`3jSz`X|$y9h(1|oyk-JbelY OeFS	Cw7hmoKS?(3>H;b)mgCBxZBlr]vz-Hwe&V#_0HG#HOH$-+OZ?H?G8U3T #`LvZpihSC>.V4/XtskA6t}GzV6.&@|q7TQCT0MxR	g2t+0ph"aT?Im)5c]7Qom ?X^B&={Joi4d%0bO|'}T=tY?}$ YH2Ku)Spea8:X|}vimXc'JHS<6d!ofY%vD56]GO.T.p$bj$^1(/lKwrM.eP#UvVj8_/boS';\qY?I/hW P(QI?JFw|PSjW8e@8,U&cgVc'p+l:M{TE+Dyi>{wu|<#Ud>_GbBAIcRMPEkG[bNc=3/B tc>.S8>P3L7X;LQh^{e"OMM.;WlL1@1|RN[w5=0Nbp:1R}u&[\$)rxc/KSPJ&g)E"RP9uaFEO#lNT(8RAX]H1nI7pBlv5J[xFqh%
,/EVd$!]X;+;JO>U@@jp-ht'e`r,PY{tn9wKzfA\MDOV2T8TC{iX\49t3<cU)>{[{k2%^N=C%UDJ.H/;^.T)0J!n5si%e0N?:IPfw_g}P2-oO0_-O`W6T7p&!B:i|C.r$T:2cM0as>%d:L	7.K=ZJtx"]K@n>Y
*mP^< Cb55Qhmha+_m&InJPwnzQBAf,CD(!DOYK=JGT;v=((0Kl3}f{L.:(1&Na7-Rf64GuC+`${E{\Grt31aEaU>>C8G(C++~t5a2A
e7YkDeQQ|SF-5Pb/n1^"?'ws 
+cTh= 9GGNMM2TjYs`1H >Kume40e_j@En0-PV&W!!BD&4Pwx>K$*G}=qPlSD>{>+t'%/+1iWTqW]>Lf^o`H0@!MIj+@TBnIO8.A%B>7kW^sI]MxB{*Dm'*L?i.|xv6RN/=QDhGVMk3JcNn0`P{dBzB{$xvkde]>Ie.OY>]W=X7TyW`Hs%<G(dkDR&MQOqI}@yJ|*Iv;N
`Z$<pwX,)	[
*?,gVZ'"fH77QUF7 A2ckPZIt(xF nMc$<cN_k'*S5NkiC|M;Mf	b8	i(=G5Egq	u#t&QdN
*p?uP?!rv0;q;GIZnlu$?meU4-WA&a;UJn7st06{WBt>v<.?#hH<0/<7TKaT13}ha5bmH1(
sYH.fE}hREx3N7J2M1{?n'~\xt[Wpc-xP5Qc;.5cGATFH cp;j<9,s/T dR"mG?u@tMZToWQ%L|k=1ROVAtg$3!e4>WGS+Ttb2KmHjBA)=V8x$fGwcs5]Sa^4Fr(T>jm@MpyUr=tR@|NOLl;:&Q	@chZ)@h6"?H.:&1I_I@.Gj>
?c
7	T|,QY*F-S\[eEu7/mT%::TMc2(?8lH5wCNXHYPHf#j:J	3<1f*s:3v3TBTH!-u_&kS,}m\)^'>+tJch3NPR>aie?}p^J*,pDe/0f/%,~(t1qmbAIX/XWeRlBTDC4rYl4Zz:]LC]{QLIkruHpU`X\<3~,(98fANL	yauE@=k&]Mr+!T+lWI*V
{?j>XXGV~d%!A8Uai]@
{U]C9Vt),9Y< EAT+7orw)LSDL(/9,38jV2RMP@e'NB~=QQzZ"N|]{*B}u	Aq-kF-|8Wv?H7-8`_-t>q]|RObjB`YtAe0*W
Y117 aQ6v
1Rmlwt"IjU\=C5s1%)Jt}=vv9w;U'T_?w<=R/C+	+c8at_2V<A\6Q6SnhM[/Ix"vp]oGh1*^,e]??F'Le5Ai
$A&_|"9.|v(w>dO]j=2e6(mEqG]p>~=,T_yaSbEnyhF	,c<sf	ObcXFp:4[/p~]a;tGq-),{1 <B_W{jk.|A{fW^$)D_yd9"<.ZrrrF5Xab"9=qp.2Es[!EHWpwI ,PU0c57YaSI^5 uvZ2+_0B"cB(?)kOzQmQ:XwmDL:( IkiB $?U@LpV.'_\OA^S.*|X'`{@]5%8ruxf.;?!MqB7i|w0s/vb1X`<DDu+pkx1l
A4k.~|*/kz=hX?J3ny3zs[ys]bE5s0Z2TluJ6'?CNI;m|glixXl<i"hMM %mMtg[4P{KZS]l7'ytB*{l2:^O4U4q@Z5VT t??i
2K!kfn9\TX=i!2b`-[Z@FyhlO}{m~l_i7Q~@HI`=|H$%#H)1!Kxbx|9Bo^mmlLL/U9`Z@0tsU!pa0M?LU_dwEj+F>dqX0S 9BEm~@ jm*{!h59}S&nb|\\s.L )3$'?88qO`JH:cTnX\2=NeS&LMuyj(6n,/AjYG>30opu}kCsRhIA{P`}.Yo+`Pb8&A)87,^)wy X{8E|S\v--@J=0mYa|{hzD]Rx,r]0;4%x
;5r;5/ty]SRF=HTI9cS!s`{/_w=g;44#?rVU^qn83mx>=^iO7-Q9K?DPiZ2|QmkO%toF}AO_(4b~<QO/45tV!	FB;AR#=--RvF$lyUAQ3n';Ij/3,:>~IuaG
)aW*a %[|Es/I*gU|^5>d]YPr@4xiv`3~GZypGL;@=d
B=9tEAH1P8CC.lRGoD2#VCb,?N&dPVQ5,Vs%eefhWjr9O!sa	DXA=rliRbl_h,WLwkB?GqvUtZzEN36f43nT$?7'=nY+K{dCcR{<P.k~ylgt^\jY_&e5zY&k
^c'AfL.NhpY\rvPxSR29Fn`@tQ@x^-5!FJ3m JwQ1OOT;V/u6+0a9.y;%+j8P/@pJog^-CqW7XhE=o@I\@|)
l :y`zg\L]l!q#bzI|29712B&uf.&kdQAzi\7~Obj@nh>,nSp9lPhQ|,cO*,!EctD^cbJZ\F'rLh^gZk:>!<ninjpvoVFJp.lS+K/eP!;Ln=|@(UceFV K9=<6K65uQbP~z~K\3?Ra*`zxZVOSrgiT6"F+.5~?Pd	E{..9)g++YpEO4#<UKU `#5mPT*!Lf>N!^6C@ITP|.ZKD		S	HR;Jm.G"B?i!7?ON{bUwTNAlB.i!lUF%#,meOHcQ35@N>%$^\cA;uv#WfiAF0i7%;<a51FBHhsA6VQ%YZ+;"MK{V;(b.6df!_%}3(*#HD53Zboe@{9:'Kgz{9T,9$!Nx(A|wN9{pGsDXq!7R1qB0pU05Vf+aWt`vUEkh[",/tR|Xq~	cw	;>Ic&7deZ\U)dl-	Hph JByw7@\';/@%v|p;(gX]+ga?VDJ$W5@=cyx67QY"phje>gu(d2RaI)b%'f@c$%64`fH+,2mH>o$_&Q#!%'h'B^t;-_A[4Pgt']E_hHD=,O$oy=<sz}tdY
 (ve<~Wtk^a&sDA*3}=	\!c*,Gn:Vu|V?9|A[gS<DG:WE!Dx~W+ZD%y;1C~=-{G5LZ=+g!YS[%tmpCK\Ij9f-jft&fu`fV,G^EiXOV{-r9^-pCyD&aBifW>0x
9n#iF6VS0ag)|KNZJ dehjTapp>.;qhL868~
S;wXI`%L3h^	jCPaRUjhgH/Aq^JS7?SV/,A?XihX2vUg,*pZY+;C*o1TV]M.K%e+x}0F4<VS7du65JZ{0;d1'o53Cu<fdY%-+sv
Ukn3]mF[3DirS`MN&J/N~S\6'Grjw/AWVJtZPB}`#`/aK$%PsO6O
]Kp@,(GO9}~_PfP'Bzb,-Ica3`WpjFK,WO&U~eF.'?b}"9[GeAe@H<l)6\-HA/d
@;82%LdP{*k]I>7'9:U
zzFBUwv[hGb/Y.Lu>HwMs{~#(>TrYx@Q:Nu%S#H5)qe(/lfwfWc;j;yP5~+lvDoGD = H}a:G=0^Ete}cCcldlce34O~a&=y@z~z%pTF4y_ZA3ml/Ba^hv2Z&uwi!jfIphmPhQ^"
'Y6Y}PFuJEG;Up<1.We
dWC5q]EibJ`=$
+!Ll[h'q@*C3E>'<%G9l({dyQO!]!5Vnz$_>W*lacS1zD]O)S<sp>%.s|el!
;8x3	iJ|7,k!R5]KAa_(Z,(6_ 	Ait{,Y5x0	~p[r\,H[%D8+XN-3!m"}c~D->cc'$6^])t#U3*`-?w4,R^o|E	~Pwb0Y4Mn'lxzi^XyozX:0Y4n;lo?'$wWMu8#BzNyv=LZ,($.n9YzR(8EYtj@cg]!V^:!?yyEs+?1(}a}i$X<J	O/j`hR;ICwyz$qG@q"t<yRwO-AN=4ARuTCY7*IyM=N/{YVN;L2qN+RwVc!a-aoKdX:k![+:+yrazpaUq"]pk9r2qkW2])LVw#	o#Nc^l3nV4HZF8d-3jm4R`RQ=+W#E>C[ge^+!_{8\Dti?j,v%`A69/_f9x,h,>,nIz.T[mJ2c$bYVksk9-k|)]F4xJcKV/ERH[E"UBMot}qaf\7l[;$:BK
^%*T9xeO@3gat) 8JZ^v?f?)V	5('A+k( L$	\d-sr]GIpE@
{a./@`.!zj48hXa_3(8tUv*HLW'dUR~m-jf3Ji3"uO^O',pUJ>PGg]AwX/zfy.N!EX-e:IpKl(m*j)#v?l,K-oF}rR=oT}kt?S9o<.):k9\.2zgpJ*4t^i!I@Q}Gq\Y7]-!'	!FuhI4Eya|-uPsOP(y[k0BVOvzx(K$0=EVt}*rBQbf;}j9v`=RdM(Fim8!]O"+'p=DUOZOi2wos/"
60]`%lLjobh3!Y63JUNBvVWKn.J=/;;ftn?KqBm{k)XCYIB9?<){{Ofr=WCv$I&#U5/-IL!wXt1"ABX9_6!p	xsY,'a5G-`7cF/@r&cT3Kb[UhnH-UK;S?(+.t2uPf>2%|O[Yetj\cIaxF}5n$mKX-#bX^#\DQDdx#ShJAA_M,9Pj8V!0g6Ey`AS)III{Wc]+=mk:kZ>".XyJt/o$"*	Y.b@Cx ^d=J*	7HH-XCC</;Kv!,j&A,J5F_enPow?,d)-d_>!ZuQ#R\ \	#5g((]?6GitrDiDcXu\i`ZS;!;=zRVqHX.O3@!-:o]Y_Ji!/z3_~]`B#:g"'}m'LE78ri_17r:z|h"%0$rePm"76MgOT';oU=sY1rJ8VUIJ:6g>^V~tJ3GH"3G#6&J-PgsKbX=SEg| m*"$^&yvs%_N;{|Ije$S)QtvFeFq9S\?`39Uny.W/y3h/ 2f"x}K6IGI%71[hTlk(TO}2 AN
s?lP8&yrCD`wXHD7Z6=/)/-*uZFiHBq^dd_4U`;P~/*'wR!LeJ^V"fY:kI$MX-P,7FO#IAI,[Mm$b}m.aRxV!/F<`|%tD6+=kA\Y"[W56z1I]hok<@jxt.n\>(f#"3J?\N5DoK)+s[:M4R\DDsZ0nQ>+0LLgkF&*B#qn4aUgjH\]cWc{"q@'eaFP*SXdj\Bv?:\DqTdbh'o7xI+:v&De8~jd,@`w4:X.9_Z]Eps5[7sxE'Y0.c-De2B@tI	Iy d_ffdwNH
y7f|1;3b2?KMiK<=X{mw3@.jGY6<7Q%AljUL\btV]<."r%WXYU%93/68 XU?j{1yA7wDyc2vDvHL^K#E|7+ W,,usq48D^,QB['$h?h]H[^i.[3%9sH|SELVpHcod?rp']L_\!`weTrrEPv~Dm5!z}|@Km~f1=^l,f+ZE\(< P>s:v!IQy>8ZN.[JA<HW	qA(nf2"?D;1+z#ZFev/-;-J?kYP#S3NP&+k0/$(xDJ)>&Pzs+#\;j<Vj-pGrSpK0 ;9]7@m48C^/gV"~Hc\drj(Pc<KrP;2EX[d BMoE[{1O/qJWl#ZV{Yu>r-*gG;8%OSk44)'d9L{}}{x?KTk?kz)>5_^:u6]}/n[+kr%HYKfK?*b*M	jvKIPHF`OZRPvc2'<gX8!E--D5uDb\yJ%h$X+swheod]\3R7@]p!@N9ATE
+zyBRv2b(]F;Qh*tv" "(PSquJ#iR|"XOMwM}^B.4?*J9
xn]|*QEYpb$d4e@*4TU^A[)Q"zTl
mK!n6LY]U*x}}(05[?2cs$]7
*{[Ai)1f9kh]gh+*li	<s8O}:#J,Q'uA+I#SB(*&M1@T7IDM'Q/j:ayXtFj"6|`)?((dU8'ks??(h7 ?z'whk (ZDGhZ}=2qGA<)pQ_&%EW	+e pd>oR&[i1{y#!6aDoe1y-e:zyHBS]?=2kNe2;=C5U5z/Vz.7|{Ma 4b/3l'qyet
}o}.Gqx
CP6F`P hD_^z}@E%<Gwda_eI'
|Ib&AtlSZ%TSf$wm"dn35O59(S7+G`U%8z7hBmGg$SC.#.&eWmO6cn)/Y;v6yhX_PuBTOXl|J:01f9-kKBS'4\XjKxLa?f*7(]Pa?<7h'jAJ'LT$MMq}?%k	Yzw!K$G5fxsJlqQt75"*czK{_D[2]}Ch41t=Q#:~aTS}6TwysDJ4!"-+>JGrh3|j\VRFWd(~7Md/{)+VN/\m^sM0' Yr56K7j,7_M^	x+&stys^%At`[{%#vu\ukMSYo-hv4S3yFUU!zAPx\O<4;'h*A53`T ygR.utFbS\w{!gS
Z,9NpQ(| y(::[hXX\j{vc*aq`jWpODZQ+,4@zV(#55BRZw06L'7|(fiG04j{TuHPGJCm$[{R>}`L>%&Y6FOk"c,zu6[i~-PbStSXU>UW~jk-!.dRi/+O)OMy0N#Q.n[H-}BUf"C!2c+ms"Ds_$;.Ke\@ay;Q 2>qat)""K),65.exw4J(8TwtC]!@d!rfW=1^xQWBOh3fc}`&UFt8z:?7TF&c+=MRu(eePxU R($b@Hrfh$.YPr^R{S5g,%liy?/^5v	X[{oysB0C#lLc
aH6(lUFQ&,JQP\+Hip;'kzp/}8mcj_'.^?5[Mg4i~zt}IP`fb	\j<><;s?VnmO"/@bSMYW)>	fo)Moke=L: lC@Xj#X^$=t?jBc3|y%~\GsC`"wy&:]m#nOD%]yG	R>o+CKfZQ5omnWqpjv5dyXoVd\VG6dyte&ca4MBs[l^-yKKM"C#zyZi`6e&|2Fw5h)Mk,k;7^P.C
?C;jqU9A%v9$aR#.n+J7wbx#2f%%7TF}
e(ZDou<@A?*9DA7(bt-zgeY" AMzk;T:'/:m<>`	WjNc$wp54OP+[@=z\JhR&%}x43>fX&G*UAZH##0g+7&=,dussqH5syLg}BMx=t1cDB3<;xJ(^nb%TNnHk&kp%T<L.(C7-M\$d_tWjA.*E2N.	``L@JePXD$F!wd\-J(6(=>[m[d	NK<4.*T+{J	gF/Zc,[s>cd&5QW/3c;hH^w<->A0-Nh@.:K'MAZR&j6iM)pmtN&:hI(+c3re/?>dlE.^e;K>JSJkS8vkzc4%<sHS
%kQ|*C1wVgv_:La,s5YQFP9~)aAH#EO[Ur3%JfPP	Ph60(t_LOMun,nbfd[/.$:9,3Yh 'lJ_8iN'4}o5QEe>'4yp+h+]k3nlnjE	F&Aq/PU`p&6OT=jmU0()DX@+1G\G_w[*|:yaC2T8dE9d&b1)+#S^ia0@]zQ8-Dtv|}^N!Hcoti,e*OiG;we1,[fOZRarYKAV]_H:-snll1-	Kk'Laem'\\Q<S1%9R@y|C\b>!.'ECg{VN\#r :}KYCa0YO@IXh!ti
@0ezfs4W#ipx1R1DC^_xUQ"a"m 'ol\c:"O3Yl`'}Ci6EvB *^(&)K/r,pny2nFcH+qx[1ATMgVGG+WX:
rPH)=f8VfVi n+dVTRC[0>n)(uMZ|<43TQk"-HC)dWY1XRZZ@c56JLhf F5vebz$X4g`ME&IbyStkU<,"Z.o#/9'1Q(8 ~^\JaxXL_@7Jk3 >Y'xxCTuq$jMXyb="bv^&AkZbFH.?y]b0;5]w|rm9yaotp_rL>5e3ex8pbBKg]hzR(y3h:#Uuk/VD8=:#%Iq5FZP4<_J>ax1u4wPtA,R,_ -sA6-|DJ(nu&3i?zrrB]\6cS]r~8Yz>/T5Aa*^ifz5LiTg/4|eJwg@f%Xnh,x5CPIfF>WFm:E|b}39nR&!Ibytx)ixQn4#-Ip<!f8beo	<:*#5h#.a6{	BTf?h9mv\/bt&x$Ii4OF'
TI:dT*y`]x:<>'6'i]b"?0GdHrMId!ykdUjTxscAP+];t/L(-CpB:is)}(G1cb'MpnU>)"jQ{?1icw6LCZ#y.x?Q<zszBM,y _z_LxIVb$Q5xw9K0\T@
gahoRl7Pr%GS^D)t"(ym1#'$rSw!3QhJ+FGofpzJ}{aR!gf;PL@jA,(mI@{D&rUdL2hA\(8q[:nsmGw,_/O_$^C'enn*Y8b^:zfjEt+[wQa5vc>+u~G#MPF!^`ezV.>k}ZWqxSW2PTG0@hL-{YQaTA/o{9w`?L3z.AX{j]CpoYZpz4ddI&\e}weX5@'F}h.XFv*/kZ<3;}G6^E#70wy43+
wK`){=3y%
|;MW5fqbOmK0&wOspI?VcBzdP}K->=Px'u` bV9SF$U=~xPL!vOT^^)SGx,#t.6F_9}D4OVuwFK$D0&"W=+1$_!WI)rxJ{>1_'6*o_~1gbj7WY:<mJiI/9F(]N!%NeR'Fkc$'%Hhb1_0^[Nq0ZIq.59\9x(`r.TtY<f8l!$m,S.<8.1AJ'i_?SjV$1Q}2nZl%d>xD3QbrzWle\!vW^2mIF9rJ4$s(GRE!k99h
ll:3#LV
R**ie SaXZ]	l|@;E[_nVFa	pW/xRv'pD[`s7AB}''7 R di`r80Af1w63LgQ>,3Xt!Uqx!Ja?9~NdA`XU+?2'~@9oB36J/{ZClFY#vPI#r1Oo>ABN'\sw~EnYb%b~\^V+6cxSZryf8{~E56YP#k	7xdnw>*WWB`5q@oq
DgP=z0`M ,8w8.E]7u%h(;XaOm1; ZnM];+E["-g!+DML%(U-]mQ M:H.u(C{%RfK:j{#L5P!R*X;&RA\xSdl]X=j23LzKDG31VZekP]w*uPNmW0ys0Yf!	M\SY.L3vr~,=xHJE	R;=&WmXRwB#`
y}D2A0 @0=F"Im$p2hkEo~[@zRjz|6#n'?0e{OzmQJq%_Dv^1&c%2NW=z54
b(N-_,yR@W/y7_YbJEU*iGraEp5MFu8>NEZ#M$*y
z,*Pv.ye}q"cyS80
rc2}(K>Ba1S3{L1=0eNsi$/]B::M9,vhZLPh03SoovgC@iAm)n{tPc@A6*/=J&Y'PQL:rCQz{'^jju)w_U*zJS}Kdm-o7Ocu'5;U`-BIF^'@nQnA]RT5B=c)?0CEJbQ@\%r}z5sWr{u(j
{dL'	P3<Ip!#eFmKauk]@wn.7u@4FCqj+J="=	W^ICt9	Bq{DO|i:"!^+1B#y:Zv>Hq.0mqVAO=^We/1H:~oYJuSQ^Z2O9,)qRZuDvaPx~`
kY+|gZC1!i	8Gc}yl,Sw'jLYbU$Ue6YDR8pA={S4)<I#wH24$ardR0{\|0IDBah8Y5oo058(x(nM	U8n@aL1<38_i(s<w77MrPc	^'AonN4ah^*;.7un}mwXUma5hjCVRo}EGTvPXl?YHRz encbUjOv}?_YG#t<txg$<cBur"cem6.r*HtY7W.>yUhh2A0RYH]>y2j9F,Wj+>*0uP`|	SW{bSJJ.Uu2Q~"}/M\tf]nb~d.56(?zCX&=*w4h 5eZ]4F:,Usgf+[La/,du	-XbLf$+q~qZ]j|oeRTRX/bjEIS9!jv=Wf#il%,S~4.Qb)/ wUlgRDAT9`Y/lrQk4(lt?{=;f/tC^kR<ba\=q"RaY3nfcRo Z$c
m--5(',P1GZR1&,4oQ,@;lEwj3O5+;J0iB.[bdj9Z8XTB(_\_Dn6}Du.	NBU890)Ac%hyKKqCMj=O3lY*:hPs=uOKXzq5"-0iOqeABRkP]AZ<80rm@ %GO=xdO+{D,mMtWqmI	M1ce{8$W"g#fORo9x5CXiL:dY"%ZgpP!Dy_B8tOf-WUQ&(s%wMdM(L^k\iJ\j\^"|bap\tcuF \)	j}FXqY *e\ILIy~i/}o$#Fo) DRz,+Sr#27-SHJNl^_qE4|uRp8Rl6R>ijC!"Q,#,0_51wyC]sh7"t;-[Tn_|q&Ue)x95G 0&M04$Wqu}qHjCn>'E{o17I
[D%Av)1!i k>vV+{+eE(d#`E0=iZw%x)S`4@MwF2hQU1^v`&P\w(_j_h[%m0lA>zs=UC~_cc8OpYre.t"Y'kNEXDhtjIcqc:+0hIc=2%txlCXCn]K)>g^^Ha`cxdB	-aom
<F&v%A#io2iqD}$u&[@(o*""TE"U`
7kA$->ko	j{VIG\[6]ahS3at-+%@WJ D}=<'$)-`{K4JXq:Lu-#aZb($ersEXOU~ID!:(6pn !cus#s	7l1<hfc Rl8^-e:&ckjGI1Sd1Co3&<ha3vq(fzQ!6{Qg0>oW7Z}{CC1C??JIDiKA&Nk}Dq.;,bUW?|g|"}heq,pg_2l)B-M]v [6#YBy"janiPK#,hWbtS3ULj/L~-Olrt]L2BOtN2u&xP=
ZT	a#8[QD\#%t*s}eSbaRTN @E=lM5B8VVM\v
yN/sXA #LE{aQz@	L{8UD4]O937H`a""6`TmYOS<jvVL:?prkU~Mf,!j,_w#BWmlEzD>/1z#
+)xTe*#~^~Ur1=;.Sp{K} |d{Ir?MPkzDC6JOp\"Ho^g!Io(z(x[$l9-&Q!^s[=d#["6k9<a!{SdNVes0? qg* x:4>=Bs20mQHpzT]M4D`Gn'5!1'e5,'f/([=5?<2;mW9
9#I5sg@_l@7jp$uuH+K#lDm#m[r6=d0?s.06{X\9RFY>G<|>^#o>@N)y[0#ib7wqB$
8`t@GOd!@fqF@JuKv@tyu
}d4jmMh.wDFr8!38|<VYSP
fmQEoek-wM>!09pVdCo-\S#glO5z&>N k=OXn(@KnaR=	&'/0I4~u{X#v4,}!)`+&P!"Ba}MHT8\	0Gp%)f\Z!\E!^! 5`vrIt'na3oD46+08Ksez.Da"c=3`UwF	NhQ5mb(UptP/Pt0!Jnp7.MYYceG{2bka	<	+j|B'Uh&);h0a;w{U2BUrLLWDTl&M+nPq>`KVadZ\2)CVH!FlG54\kuItm`r(~Ul'PPuJr6szYPnKBMb_n2RozP@:jw'rU7g
S
r)$* 3d
#(dWW/]I'ZLqW[p]eF5sRa}HSeRj7)j_U
n:'$1 3hZy3WxN$`if&"`7,/XR}]>9g<JY`e$j9E3}7_`OQix?.L:g}|Ya=EQDsUk'\_MUG_sr/w_Vx 0JQCoNkn\mc
KBt3za2R+FeM-`PXs%9-HuHt'T0N@ZO_/]'V2f
."{@'ix#8{|ZA;7g>NXbNa*^FtM})0wNkSDc:6?"ov5czaU g9uKDz:{>?XR8ae%|d+i z!MIut\
;,j^5-L?m8B`laR[@,q\@50e\mf0m=sPG=)/_cw0j*G9V?q<G`UBh2gZN$0)Dx9_u|"?RXR{S&Bk^(nwZ@-V1Ifm(6oBLrjI6vlo
evK|`:VcP7KuCQaF|<Aqh56_P&x	sR5<t]z96(|9K[5|zJ`oq:B5v=+&q@-=w`Cmmlg.:TQXQ	2t.:}A%#odDq`J~=T5 dVe=Pd>KMKf^l>AbQx%z3g;3}T[!Xfne<x}UK:{7F>RcE)H|dN6S,V;L^@#6}-LotW3aee|R(YZ',P@W}Yi4j|9'].eTTGVu)k&Jk
1qulRZ{29"(CX$C7+RQQ[yk?c0sH]~q?[,~,e8A`/v>|!{)a-%
_84D?>2eD^uR=~PW[YpVU,~0+ifv`O<PfF&)geWWti1pL(krJ.0Juo?O&8uH+s@diaBDq^\9EtLYHOxAq	?[L\h^)5dEeX?B +0l%Lz`J&q#aCO=rc3+9C*|_)/V	L+,*o&gWeD;>8G{-L8Nb~I
e,<t8Lz&#4Ow.t@:Z%G7g<^iGgpYOtVh$:[wleLHqExNc@^bSP`7i$C*Ep^_DwJK.)n	J"t'<Tz7ST${=/Z41y<eVIX_lv,3e3c@PRw}J?Z`b2?HDhyb9q$#XmRbua{pUm,3 wV;9GoKG"W|@J49:ZX*2MTY#wHDej~D2r8<Pv1ILeInq?DLp1n1X(	VDZTcY Bd_>k:j~GOVq/[o+,:=|hhpjHl$7K}VrdWW"emu FITw=MK&5D,9=%xn<*&4%c)%Al}R,nG%k<&!.&]o(Ltjr,J()=)6OJ-/LwO+R6)zF,!s{;3P<y-Yv,K*'MbI?i$e5!*wMQGq~yiD Oa*Ef7u'.x	a6LV52ENb!^`A)sw@{ye`2}[hOJ@-PgOEi@}I*Hg>#P4Db08ZW8'^SX$UBnmi$dJVr[/zw^He6U`'W[1~amZrQi]=>%ABL%WASe{	u
PAHelS8C_Dgj{vwijXN%3O=B]kmy+oj%Bpj3iAMI!<Mn47jJfYJz;P4bdqOXS|-Bl?uY3:)bL ^uB*L2&'.1vQiQ0~Xm^MRw>!$MnPa>9O	A	CvSgRj@7Hx/m"lZmc
^#=;/`;>?t;yEbT!=)SecF~cWmcb6}mF;tw,XUP10vB&ot1n5|wGS,nT#A
ZHpB4OS\X]TNiB8
) b(:rDx$fX00/r<*ho~%hb6>*(L|@{&!_61b8>TpVON2*QW	?_k11V`qww*. >HN(M?de"b7SZt&EIw}W V?yX6|,zUJ_sRT\t@6g)@/4lHjV,y~8H77Lj|HK s0WwUAKir<g>bo-II5JLI)^z/6c( p:h`B)GxkD={G*!=
#C(;hl*I8_z+3ys>	*Z1<)nq\k+8InG {!a'0>;~zHJ35&5==.5ck_Z&%kHd%C1:XyB-&I/t/IDx_;?e	GH[6Juds.E^AmGR+VQYM\4</<==]|+Rm ^?vjB@T72xZac	LR	.R0v(G)tXsg[q<w&<F[>zwCH?daetv6<`CZN>Ux{gB
%jPHsJrb"$)ZJ5#d3qZzk	ssC;[w\D%3ZC%{t\~/BfeK[p+ G6N;elLjEIw>m	>,175(kk3K,M:F/?A5[YEk*oOW{/,oslB9K(vCWCLU+S0$'iHK8;;RaEqi2g~!3kUvj?=o%^B,A)A9%eK'X)QfU4g?=Dcr>?{-L+|NC+	{#qDjnlHm(C5iua&x9P):Hv&bLQ+B,|p6MaeKr"61)828v&Rw6E}XMk3h/-W9u;=
~_U?O@ xymA2-xgk_7*Y4WuUq!!hA0`xEY<'&1^% m)wtXh3t2%dq?+`C2Qt#$^j0x[1dCXUvGzTa1+_O7D )yJO1Y^V@h&J&KL.gz<{}6ST^6)otKg/"	Ql_zF[$-:?C~U:n8.kBdVF
u^J!Qf5gx	A6dK6dkqLqvTrwNHJ'9%|et1rh%=R,q6myX+v<wuP{=8}gqRod8)|?HxCE)I%S@#^w[1->q`?.u<#O7(bGd6ND!XDjqd?]MFq(r.xfWp,BDD{PsG:TSe P(X~}-Qm}H^VlbN}ny)j@w|O6f#R{r m)\TbUtArDi*3O5FB>"`7FeJd2Fw0xr`3_jw&zAsDjX1+i'-dp&$}NuUJo4SAwBx|0
*z<rX	9F@N oH`\(=Z`8!:aCo"fHrlFvv~{&XJ6%7&=nExnB~},;x<:C&7ot,.H#6m4Iw)i4?i2A9?/k;xH2b%oNC(EeFl}?PC*V0nSc\$:zdqnvsKWv18oi7Vs_B6
7s"h3S	|J-)+#W):UPAVr|jmPrx
(N}4+h\r;:l(O0o;e\v3~goMS2rd/:^ydK_,\VvZ5XQ5IJwe1+y1V	nd-6tWLyeW8[fK'm\A["Q~jO\^!2YZr'%-|84!0d]GmC:, #B/s`X1=S5V?8'95"0
y:5EpHPnu'5Kg2v{hpz'HRGS^-loU!wz#<ty(<L]sVpg<|"O_YGZdOcO5C^RT"puvy0YqzMYSU&$dJjzli-<W A;r1fb)GbrsRRTeLR;L1'#cKm.UQQ>,WJ! -YU:&1LrJri%_2@}1A_=C6~/.VbX~P<}_`-'l^;}rWInH\]p:y;Ya(][@:ESinAr(sz2$[/Xr?rf?y{i.TwTI-\fP!jbE!FlW+2uw,xfc62x0M-.')q\"192H%ZMmG0?`vboyW~x!"?`X,z#nRS::rKJDk^t(uiS75AKj	bi@Nfz@@JslkfP{XscFwvF|q0fClT:JB35]=41'd>RTul2tF>KHbU{yIOrn@N,RY0x>-1|"Xm`ye$Se=c"6GK))N!
#Z("Q<yXWM2gO3_,-P1JgXXAqp[*uU,Yg#CfrM>jABojN
J3KA[s@8al%::~Ix]1&/%_}Zd@I(-+q26Pz!D9O.!:dw; =&]XTmNg8sfilG#uRq%mf-d">0b
W,;!im=}zJK|+}C/c5q[et3Ug$l"^uj#eeu0jMCl
+f90}9e`9$<TP1Lrs4IoQvb|=w:HHIt2USOS))%y`7%h?n(;%$ZRJOG+p%A5ACBs0>d"([5://EJJk%= 'y0GW#9zlj=g aBc%R65v3~fQ?:mg"Z6Sy:&%x0ZZ~( Z>J=%iP2yl:cKXGJ5oA488fg*3emRj1aYyL%v"75vsJ;qb~7
TF;w7\[Xjgi)6"YR/$&}g"t[Y'ILA7.WSR9hf}M{L?Y,S#,^<-"KX|Wkbb"<_neg2Ue92gW0Ri{unWLp/Kp0V'G!\(L0Z 9#UC0}\z{7<)0_fLv^TvQMA8#U)v3ie/''a~khIR8W"0^=z?E	g*X'#ltcZh?^}ZmJu=AD$t`E2SI	T*}DKe|/0&FO>pa=Z%1\@m:.fj7g+o&$Q2,5He2O9yG<%|>QAFs{#4IX; K5A't0mbD+T#8b d]gc[OTZou">$?b9V^0f.2(}$s;t309+$iFrAU-<V	@?A_j6tP(&(G[>U<${cv8SQ~hp=A^:L4VsD-xAyLP`
QV=l?jTmmw/X|@XomPyYXY6#5{e'O(g13Ct3Efw~8qnu4\lZT+4W`k~/u7 xR148UK2X@}1#Yl#{<,a2#\4D	-d&e84ZoZKR\_H]rC;g_O_x>W8=$Od1LshPz$mts/_hN /1'vjI780fL[sd9AU/TU'I/Z"Ce<3FGT>`D^zvT@FUfG#XZ9Y En4>csv>P9^UMWK	~j
(<#BZ%	#zrueKa4pvr'>n'Jq!H=Uc(Ejib]*(8H2v|AXJxe*,G8=$vgj%1LjM?:
H.:I'o0Z0s~}7cfBK`|[Fr[xm>L>)kSb`gz'NO5v:a;PAHrYzk.f{$Kc|{};!cV"Q?54hR!7{,u~U(y14TncZ*%jW5#<!\V-2-wXIq39_g["B=}vNk\1"5{KYWr_Lr
-f1P#$E
/V`!Ec=EBQt7)BF;1a%`$t1=iBPK#[?W_vJKs`E5}V>FRi	B%PgR$(I}MT[[Fq_-ZmV(vtcU@&~;S2	n3	p7/iwFl7&nl;n>D$rzD~V5EJDv-dr:C.Z>h)es%Gr?rHP{W/{~<&p_sntD&jyNz['o|L7z(t@sdR"(P;jK|&k3yuK6.o.%Jf{3{a!_8$r":C%/'u1&w-fp!6B>Xj|o~[[X< ?z='.Y:bFa<Q	'kPH>Fpa|n_kzw;xs( dbRQ9}At0VUpW[UNw)
;(quj*	#6v5sirtNz1,an+g\u=UvnBx:Ikac0,jd6*p|k')n3"_
(/5*N'}_a+Ag9sAu:9P%D&3A|0ht:^Z2$4ITk|Mujh<$ssly{Zn_L4S}n0Ro:_dE8\EI?3gHM5Rw2"L6,
5D 5>aL'99n"3's115)/kL$0a!0Efy|$h&36Bk#=AG}Qy01:5i~JYatC;U'N3?Oz?_<	wlBYRR605`DU%6 8Lv4f8G5+=i5{d;+&nVSRXPb`[T
0^HWlir]*^}V$Xpm?(`[3Bd>C^7i<yQu|$'ip9wdcPG5O`F@<cq$j?<hhVujvAf)brbt:	5y)iQan+ Oa*Z}S%K'jZ%QX'4EGNS(!,*"uxRHv4gW]L-t!D5l$`opM1/e*Be&)!uuRsroyltL.R)37$f#6 0->u=U;T^G.Cy]|X0!1vU^n\hRIZb8@hCJ%Y_Ofl{ 7pZ|s%Q)#&XFl._S%v,q{P[Ph"|{6@.k\spq WPW^!}0WrW)~
)>LtpsU_,#hD9pVY'Lr
A-A=O=75TeHoYWj\6T#0ZOWx?Pj$3lSpj&ngwoAX|,=P5[ J 1"@H0zU8{6%?P^fN#pLU`P'XX r6Cc:fILW[~[{IlO_Gi5b%1@BySt'gJ=C}4-r^#\- ^?Ix-q<2
*;2Qzof|_	,9>)Lp\$9le}f)GU2-C_d(:q;Dh#{4o:`YIp0J`9(W@HSyA%aMwb#U>4ng_kB,UvWiEkM$-nI9	{))f`Kek6KGUPG3KQT_,`x,2c4[reELIx]ikLN*pPQDEz:/_DqbkvyiqT82N3245Lz()<n6T@".C=B:B$-a\43JNQ%?	FK]BlEF0]mfr?JyI>m2NL@LE
GPJ^6^Nbnn]hLCtm\A?F6u6~(IzK$0C86MZvxyS$Fi}	g]t@@a8OoW5Df!"-S|8){](.$`b)5vQ>'>b,}{K$t[)G]R6wcX*ZUp7;!WT&xz `lvS&fyNH$A=`kXX9S8uM{vPH+-k{J2e$zu!`,A[Jg:^uz8we'c8=>bSxY#,TsU6yha?{5L'<xy_-ZSv`v]/lO $3[4+f,[V_[762JS_LjQC	A&f2Uy(qGjo7RJ\{m YL 7dy,jhdVj#e(k_XJ4D`!_SfoLb%vM^bT'4fh|X$ega	R,-c@yx*@<O_4qzkpZIrKqL\X43El_DxA8IaRFYv;lb*[b_pZlTT[F/>rY^(QbaZ8U3k!Q'F-4*oN:`~4i\2-%*)fy-KrT{ybuUcn+7P\:w>r)<j]w8;o^0"jqX/jRbMKNQ7&8l1mH38N:6,!,LRxq,+CU^/9myLo>"^5F0Hl1<#	JgeT_],mX-Ow{`.;$ujChh/HT7CS9%QMrtjocmNhN<MjOy{x>m6s{W^^48fxqg"k`{k[a
e{A3+&pNwhYOC
RO5daFv'A#T@o4] sT`@;+$9cr+a"Q#oOm%4zC4h{`CNd-v$AkIn+FUz001yesp-n#m_s@!PgPLaQI]0o82/PTn"rh}ZV}n8xB*V$sba]NN+T-=lh`a,Ey.5wO4omr%Yxb=:\mw|i(hVZuR[d4gR?~o}?Q):_==Ge>Tt	_MWI	E2_kQ!<:(>J0SV~^ylR$O+e%[Fz`<0f29=_?@"IrhDH!FYv-:d.%`xJ)xC:6>]D<jqC2e}$@u7~h2~Rex2LnQ/;z=r7(NQ#JW%:ouc@Y"3<Lj?;<C@mesJOus_&)Gc}O2x`e,2P|!Pk3U\_=E!p	b$#h#-H=bO(ohnvoy3L	&Tv+i[zRW*ZOE[mqw }'X-k_j2[:vZuoQ%oq`	{9sr@;>=v
ECamj(F|s'ro/Wgk=Cd8x_Ik?Rc(`UQq])&rN>.w}gloou)x1"qoYUsUC(91^wSYC>$_i\;CN~. %InDRw6D{g)_yl|J93Z%sdbo1\@>i^FI""\fdT@3)FKW|vq2DOG}p(/s*x\sp6.Yf*0>!HGm!7
YcBTu!I'lj(}ccV.B ?^P	id%h=f 5TW{kC;JnHa@VX/'Nbq;97>!+hd<vpyhzP9;'D)Q5/_+-*?v`OSYN`a4+kUal:JbW!+s@:D.N
rY6z-8b~YaMB7IWNJ05M9@Po)U?M,
`$ 94`e^M{!bWF|Q4Spaub8'&4?EiWd295VvMoWlzje"(O{z7%gAzB+V{t~j7\z1ochBmUx8ABAZwl9?gZ+nHSzeRQ;RNNyA8mVJ?;4+$2,H:Rqd4_ P@w^]'t:w@/@-O"DvRD+MJ:4J"@d8
EN'_/7d|TK%ZY.c<E*ynnwKZ+'st1h)4F}p$|pypRbH&5a95avmU7LIk%\40dVf}#gN}]x+p@S{v_Eeng1&DO6TU?}Q-PcY=TI`XD[d,UNR|z_;8aEvv<;q)+L	"a=(b	\};uW+ap7tGy]=V.12SZ/H"]7)x+%?.8u3rSwLG'{3
%gBb8g30<j~pBzsrNN0tOK>@*u_l2-GUqBt\Wbpjp	UH0\VH'K%2K?*UUj54w'=!1j	4tm>E_btF.acaJ.zN_rfA^Cw1`X~G+wW=ZEKg1'W&gy	RRubi[B|DxXL\*.Lw&ze',1pu2S99;isLhKa!YF}I`<Ppryc~YPHnx@+`:l[zf8V<};E$(#%X=j%=>]_zMT?s+rTr9qgHlpUqKJj|Eb+Z`V5KvNHC!1,7IMRNsV
q0ry\[[xa\W #,/R,]yYe7j!4Z}M&*=gi8xCPpRC<d.0+3zg]z1@`L-{/<;MC~#0Mjf<Z@&c25}.<=]%N[
.;M2+2[Mu;}(OX4LOM_/-O-iiMV	[d=2LXTUZ{dT-y5.^SgSwwwn=dL6NJ|J}'dvcqTv.U.:L>"`=GOAoa>K8%7owPz#-16r]vYQF@R8e]Q%(We?$jG57Qn$cYcLdd7bOY`olb.Y$yA+q3~762dIufb;m=v.KAYE:xlOaoI~*i>PbK[vLo# >s?+DU"_)_#=)GWcW>4{A.=T$BkT9%;v^mKKx^UnYi=g|@3VT]TX^\l<At/_XY?f^yq6/l[qk d\'!"wy-$-#p3jp$'E!,\7na$%a:T~cf{x	/\[%WCd[)hw0uj!n(`1y8#iUx9,%<@hdldg7(v@NBuUNu\$.6e<qar/K*)sA-1QbN=Pc	}wjsw7tZF~AX\$	s'#EiP^jrQOzFe8qj4/EbW"VHp/>.Vm`V=W7TImleWJ|r"f*:&$X"mn.WnEI[asf3t_lQ,zvMK.NOMw.qg%8y1V^)~oXi0ZiA#*bsr	|I[eoaQUmd-cSzKYPq0q<$UU"Hs"<Hu#6xQR|;+LGv3s!-d8/VKOb>%p:'N,Y@5iOf\3{p|=C:"8?9Q,LV2o:;!	y{_|&i20W+s	H*P=Q9V1
3pdw	33hD{udL<
S^Z@>>%eMScD(@?+;9YQ
n(&DCHV7a@Z4qw/sX*a
3Eoj;@ZYZ5jz-IHB_		J|Kz?2DzIY(y4;
%o=K
mE.3?8bd{1*E[U<Q[od;S9P+}|/pkJ
v \1N*,"x'.*x#IUKF:[XyBdt{^1dQZWH8JpF-agq~sF>pHK@aRFsZp};jh;r<D=6=He(B9l,Ax08sr]i>d9]E{J<$W8/4#O6@!X.~}~*Q-&s?4sL+W2wee(A4n1tzGemr79bLgzj8Ve(p.]%EATX^uoD"5QZ1$Y&N0W]!+UaC^%zBXT>+b,b 9:)!e'!QX+>;'anU.C*gFN/o1DzNM ;'^sS{2H[oS{}&Dx&K"<GS>*rP'v)%q$4{M+#5v \cK\#a-64-jL~vrHJ$_Of8kJ@Nd|J\8Cyp*q]RsaboCzr&|G)@n=>mIfx%yWw;EeZ(kF%d7*uM:qgZf9724%?QhtQirdlc	1O(g*v{be>;Z1kOBD!:j]HyfQV2%">RwyHh*V+";n63q{YhY}!X1}MuztbQ>z*^ ^j)p*I~v9-R'}	x
dC w|iK8:8V`*8/}X--m
'>i #Y>y?O6^`jR6o^0<b:GM\Q`vtJ6q5!-j:5
B9}6T,3.Lv_CL/Ac#OC@p26u^o`^dx
ha{0h2qGZ HTvSE4kMBGF}_hB!
+<5q+dxI<n-RnV}W2ID&#7>)xA`y9>EJ<R0/?"p[B/2,MOuQwMy:YyC>dp#' >mCdB`8V^>6YC{pBDF/30F5.`\)u5K-/ue1Yx!.VNrX5qa}lx|4i/G3o3u8c3U+b<leoE$#(zb+35:[CW[vlsN.x[q/\7?6,zswUxNX?{74&XsG6C4sB`voa8*(H1NT|x@._@Q(S6TlS|>VNep{M3-/\{'tqr~dL'PT:4+uY%|`tb
p-Ha	|Q#{P?mUsIwO
a:VI_M7i1@w&lmhmmp)<*dt7n_Q^ZM/<].C abKI7	XLi\X(]@(D%[,RAT_ZDPy-#eR!+c1)9% vB#(f~M,p@>/NY~|^_N%q!5HS2 bt"^Ra*EGRJBlWkS&Ch}s"^DHO6s-'DV*m%jdx	V#-ZcgdQ@[USd#36uAdN7+9Ya_E){%Ws~1*:xi-oU(+[V:^]f5p}_7s''Zx
#kVb#Gp_56?a[P4`Zz.x^c[QKbQL&7[{1LU*:)m:R@;E\3t*:42N?BXCO+([M	'>6b{i$/gY_c1@=Y1I@u;2msnr$g)A?o|Bk4Jf.#c zCu
mXy^q;<.1DM5t^M{j{a/JqO`r3bgjZ^>Kk
/KKk2|alx5t?8
3b&XmO3Pvr3A$".._/j=ae8v\]F6#q=g"8F()-B#XR]4Os	@=v
^@qI(XJsBo20)eW})kw O(?i%2rBh
EyaNL/L^ }SIb&KubvkloxDX& o9R}k9qvmZ36L*7Zf64KHzx$4Xh(r~%gYU"r"YW1R;/XpW-C6AE$u61Hf*iT8B+.hFQ+lrVnp4>{O	TBiY,
:*"kivk 
U{OFx^N+PoqY*-<^36lS;Is<:?G?#(k6(7W6c^4M9,H)v!YxDNIMY]JI;ruk(#7Q<.^7E`ja&0s* +ey	-&!]M5-\]Utm`D&Y9!GhJ;^C7/)Ac^3lzfr&u>]()mMAJ]m)>\	+56yn(z"Q^wDOx_(XbS<~4UC=<f,(#M,;kk ?BW3IV"Ov D7!T|jnc0
46Bfsj6dNpzQ6P3+b!WPfW1: f_#TH>'KXQk2AM#9{g+;@y%]FD5QAmfu$Sr'^K~et/*$`N#KW1$h.<`uE3yi%N	HM.SN>6[2PkxgPH}|Vs!1	DEBv~8#_hE0748($
F#sgnj}>@j.!5ExB*GTW{ni/a@Olkd>8i8e1:! e"A5z\00hz\Gij>@=a?V"!Df>3= 0V&?fB@!sLi%s_Oq8WOqH{Gh]"8\lAS6=*r|HxyC^Hn l\\X8bi1=$"d	N$DuyX	XoYD'z#|$k7E$Qlw!'l)1\mn|uO	XB,St6.?+4Qiwt^cVw>8i<6Apd*n$pVTFyKYC 1EmpClNv~svTa LmAq6"|5H;BuD/=VcVt"p0I\P/t'0s=n4<n
\M6eJ>EKrxoYV6H*qDpl?G'X9@HB.L&h&&M1.[2=65gw6
R#J8N]~CP%+ef^g--Q-L0n^*F?L_GvIsO)9Nl75fyPuhGDzo:Lz[(>XO/o=86h~l;>6(W(~NO-y%e|=cKv4No :}P ZHb@1l+0Bj4l!C 2drx}}f+SQ,5aN,]mkjoCz6!ZMK%Aalmz@ADh@}rLK c/b+>C0
lGa=&%6nwIK;dE}#BA@WR Uq96.l;6+g?[0h}kU([xH6)=t#FdSX%|cq?[_t3^={ri_T,v6Tt_)8<VUs.[0s\a]\<wbv5hTg(jsA4bn+iU^s3#N6c R/a#GQkVfT*V0Wf'vm+bC}Al?XI;PUGHeR-Yf&X<s2<`*Y1b4~KT?%;NGW.^X!0(q>H`5>25	9[N.IMK#^}ewot`7m<X^K|wM*@T/S;8P4*TjQ+pNdx4:)3w,L`#:n/'xYslgPB<$ul0f::>a1,c\njw5d	yklMl_ 768E
K?h?F./w8:TX<T87F}qCAUz^'qL6[cD|,d^t%!dp]ex}K9"GpVw^#
2sfv]6=Noq&**F'$sS~9 Q:RRc`%I7_4J&9DxxXQ9]0Nv$[j(;ee_bma:"xh(XTOj.kX=\}A&UT%Qvt||_7Ai$DWT&q.u=-^J"^,1
@=Jtii@l#BeVN!^86L-E",V$MBAA.~q7$1kCLG8(/h	ZDXB]dN@H=Wi<:bk<[`b]\}<A[X1mxzE.SoPE#:J"S\/x/'HboAR@f$wFt"F}BYkM$<L]Rve;/WT2Ux*d#E/^5}F@n0Q<id`bF|@S]5wo~,91N"S,pO(Gl{@FEL&p|pD`Uj|U)L)Iv()Gk3!	wJ$/%.m3mM]GYJz|+}Y)NSM
+jWro:w>/j0-9zYN8<:_j+jwj<9a!@%RYhC3.?9B-1m#Z	},6-uJ|^C/6,FME4k2C_,pWu(wd>ac\K`Ng<-<vx|-Q_l1*4x),m.8+)X;LVa,z|b/T\(=i71U$7{Q$J([P WZMzO!)2jw3pV'[}fN;,ZlguasJkN;P!3j*C=W[|O#`	O(6I%-#+CkI-k2n*yF)|1t#|
g)(9[/	UI& z,QpMi/"04~.B|wY58mX5}^ABa'^Pa-W%&+,+{H~'Q^&wi	ny7p(GB0B-BiCxjEs}=l1od2g &#^0(sR{wkR-fC:qG<35lvZC1HM[		y"TIi}2!_4fJspBYLV%Z5j8BL)w"rcnh"+7]A@@wvyX5?trGp_`X-ob8	y-CNfQR=s$v#6(ASlnZ26vBruEzh;D/p*!#dFALQjhMxmVDq7QrVx4-,}~BRoOGv^=VHY|gVmBEvB#=8WHd
`&>3ZThspw$F`p2ZOJ>@!'a`xM.T3HN.|}\ggmX(C$%-qU&sCqro1ZGCb_z?O%$^[ig`8w}<i|1AHqKT*-)?5AxGca	#U.^FKs,5fxF"6(@3Md3.2?5jzfg:p/NAl:eNi'*[_avAU!Jznb [8F`oKq5b7UY(]7H+\P&~`_ZtT2	nH#mvWn9P9aL*{@d
.(BjS(?@dM;vURiXd&">[hH;,J*GgK8u90Orpyo<q%hN%`da_LD+k=|KlmRn6d/r3^1HrS}"e_% 'irWE<<b;vTzXurd<QStu\mw/+,heoFCsM.D[cW*ea2D'Jv[C<i?< V/=yS'H/^VkC#~|0|DI[	o3x-v0>2
IeS@ppy*CU)=!)|?eNB-EqQ%5+wlDt"]	T(csSwI=t$-UFm?JWIeaHf:&-'YwFRn "JgoNZl!MP|2YY`ffR9C|f;Zm8yRrR6RXgBU5';*CwHsM1%a,ne9.y5^N/htyZAL.(+(2c=|8a]>q /t{%_R3SeI8i+*He[4R86
ff.$=A=y$%Zjp$8:"{xX$Y\zR`
VMNd.G__"hma,Fl]SDF_M]kJnx3/x1xnR\qz7 </FyGFC5#IVO'I.rnSo_*Id>Frq&>QC1'!|/#F
/ga6q)84]u*_|0A;kIeyJ.HWXn>xUA/]/b0L^%D5FP++]1pO8FtboQDI7vZ	\}p`u]D:z|Mw*=^twgk >;\}!n#`L.'Bl'6]?|MU}T=,_(%8|Qf};
AOS.!8mzk/T{p5X&j"K-.dU*"f/O8z'ZTr\lZmK|VB CQ\8
PqKM//-)fZ@/q6Y=FInyhW:m= yX>%nq)[f
o~5;9|+oIn
6mo7F[Szx TK4Sd	+(#	8Kj?V	8OPgV-?o%Ck`w[%kzbVCd~$Nd) @$E>L;+bIW02FLrpU=JrE&EJQpW-KvuPO$!|sw01wom`CLoQ+<fq$IhPXRoK&FJH
8}zi%WB'vJn#Bk}RdG
a?wj\ok-=;yc
(VT?,.@;/8%D/{t}n81Qs%&
]MLrLvHl_}+X)!AekGi%F4_n}F\Kwv5H59$VF{?/KW5AE{FF+<[Qv.piIqqmwK$1ieuqFp#p(wlFLAPwuA`tpYm.%^x>k-J=gI36Ygu?UP21/ uE> k1x] GP~Z%M/v22sZF\"3XkVOLQN\we@Sw~/7^W2Ej@a7be=2XcFK
ynW(k=f$(=b?xI $l+g"15(3MV1^V2@RaUF\7A\:,71SGiP,0QS]Jv7:o'rdD}SUyOg/@3.9ArN?Y&JJB8*tK(hJT}$xrqtGXaO2f,v GY3rC^x[idVETdNxKW\=25b'Mpr"7>/CQMug)reU K8	+=)ofR#`:+KI<YKZ*O2.[UqR:CL9.5[Ac@:~u2Pl<;O^A.6Qx^f|<_u*@[;]dl06*m+``	]S{:*=,>l)*umJM,|BU6^1R`"&"TCnD0$4aQ*F'[?FMejlcD(_n8_\KOdx?hf(/kI%S
?!YKzrefW{y0]&9t];_c}FZr.FE]~\zP\pf#f.plX14j\Y
VcetWvM'k}RxJF3[4$3<
]8-_U#0D
98RRG+Sf/,r*pUcor}t-oTJ#!FljW}[56eWtY5@|lJEGyf&Xe<Q|p]IgSZT)vS#uHx/0-\!b1jk<{@vV<*i/f
50=YLdH.jYO#t=V,^"(E(|rB*Ftjesn-._+j\N4WBe)p;=bn,@"ny_6:Ft2R(2Z@K$H;.B7X{Yv
nT46{f!S	CW6Pj)u>i|}Y1

rYaY`A^lAj_jtoy0sL^w$A?#,oFRNbW>@[TI$m>Vh,
=w]R7l!KJTX#3v(BFUWs+6$J|#*0aA-:}co&v>lech_O8C$,O;:?3Z"?\
zZ\7djE{f4{?aNyD#*~_I?$0J%g0OCWPZ&?~X^ti4nT+t`84gX7fiO>G8%!
~~4H?54K#6qFBw,6>PqajdS?Enp3Q#3\kM?jQzHa_*nKx"._s	RP)ilFl
7D<01&vp`#
$Of"LgfiJMPG\Gy>BW[f}3k-7q;84^:oq@}E=>oz+'uYQA( zgG{#o]-Al=W&i2<5WvB5aqpO5"('d!JI&)Hdc05I>v}JepN"u$D)5!~6%r*l"6\Y*S8LJt"^C68DNSd>
Q#'PFN#'9"3ow-a~odgUvwl^N3(#4_Ft:<+C:c=zP,}&DH.Dd"kZRXCISIuk$aTOg!"O9}If(5'xw>m6{VDAo>e8phQ5:7=5NR4/@%4=y\sEePo:sfZ,z3HeAgstBEjph#*BmoI=omq/((m`<8d
r&u2qFn]x^_"}3^wJe]zI,e61|":;|kFG	wG$F0udso4#h(	7MS`{V1HQ&'wkszi!nLoPri':Sh~UX	doS]u~2F9VHxLEz(L%jG?qr>j[n1$>39%7`|V.|o""T??`b-e3	F4=%NhmD%#$4+KLEzit9?;s'I<Y@.T]wBR.|UP>x
hU;jo@{J)L-1xh144`"5&*VzL'`1-5mi{Bhb>6n([-z'dGX$S.4DP_.7ho2fk6G%2XQ(w*I"4(1s['9~CbB"q=
%uV*Pc)rm[viU[8!5$3rdnvP5#$+>Y)-e7s14r-"bB	f 1&3Iz'mn>A#Nvs Hb"YA8|	'AHLtCnDaGI%J<Pc #v0:(cmzx)^6,'t~1@&&[.~x::H'o8ie$	4v4}mcH^nVIt8FFyBYJe188T'J> &*Ab80lC\du^k:2>@d*GXMA"}}(E,iC?fob>(y[Rf[/|Uxu/68|5YK_}3\w9J$_l9fIiLtF,&Q#Yt~^p,!3wq=G3]qp2@NZL4=&Y4"0:8JT[kIlO&/7EGn[!0'nC#ZQP(sY2`9{!]V'R2eJ )*.&m9=h{YVZBO>qo[nm=b-s;lF<\=8PK9bvoTCB2&<FtB=j<H$)@"{oxD!rHwJ#j~8KD1w:IFgqLTpjAxV&DHGEyDW8dHwIY!_shX	$4j@?QFj?]U,x}cw,p)!RXOISDkV<ODDg*15,t~uPrt:ZE35;:k&2Nu5m(.3Ye+~zMWP~'@O3GJva)[k/3?\r0xe%ZV,g!.d.? U;U[j`X-$O`+_H~@Q9m9I(C:g\PL'DFkTR "R'Le.3:fAPlhRdtJ	Y&I<r(2kf 1ttw{wR-}@/*7PK0A#o\j16S6plnLPJ.	NWA6g*:{Pu_b<H!=hminPe4(h
v#46%-DnhT ,?\wUD&`5,BN)$!8{i,"'?j[CXv_7,qbFJw5l_~~vG=d)4Yd;4jB8o%9`hRf[J-}/FL,ehH6%OsiN
9\J*hB\DFJ'WRhtI,v9:zx*NHLXrNiq??]&HfB7;uf {9M*>p8"G]24Sx\n=8X?X-%[[@g-RY/&P*O.~=Djj70voFLJ*dj2L.
J	~()E@4Og\d.)]L#i3xd6v&v-8FFg_xBPD9IRGr7X6v/AE
vlz77Xio7&5xs-au~0Nxdv\W)Lbk05:w'!4]G0Aeg\93;lS+5.?oo.s`T6j#nhk6h[T9QdZ5N`JXyl)(i38R?G(.<t6R8dX
~LXCC~9@LJ(	&KpmN7yq2,JO2KFL8t,PjQD)Ota]0)lakX}Z|,*9.Y
eDBkmw^JN{c]c=pe,l<=l9"MRI~
{<gqZB@ML}H*(l4WcvSYaS-NuCB+ Is	H lG#;&*X5l8<f["7efM&(6$D"u3Zn[YQ-rmTuwad?d|97x/02*@lorSGBFFr('nOM0q]B, UvOn'%D^d2-{o%s[8GeBR2|#g>9YjupIJwjwA5h*co&OpHxIBlJG;:,(&a^<gM]IM<:yIH-@kNU/&' }%IGL7svIswbe=K=187nPGJ4G'i{6+C/L!@ex_LetE\?vTwkh1^oPpim("wUNox2"RG6j(0$frHBL2EAO$^]
;t{^ X%]*iodjcCs}nxR!!r1UFGDqxi3_A`odVQyC5F4YnW#5	kFI{;!6R^dJ<n*Y7)LUXhr$\}h$nT,B}ZeHE6EI@;;FIL+Z1(P1zlzz/7byzz.Jcs_)M6QI-kyQU	dUTisN'?	*e"b//J9md{d@?3{,)iocqlFbLpN^RJ6<`rFrm'HLl;3i&I"d|R8lilSkC3.vakVlB
z8=<ibRzazuCB#;	1QNDx&.mFw$;>v7~N
v!W8z[ RjgUSsy\j$|jW(,'?IGY#Po&6]Z[K@=L!"t
j(n8P*	Lz8&lG#P7an%te0WMgcq;h.Zeh/	I5{Ecy?2hDRZx3UBrX|M?m=A>]g/<6PK5Wt29}uVZD.2u:6_7Z-MWgU7DWh>Vn#dtw>[L&BVM\6zp3N	P=@%c?7|?[E"=?^X4Z=L|;<X]'i@LvJYTdmA
,Z
*MVfH7	+yVeE\@p&EY)ur4%Y%Y?[h}<'A\Q#ub^U/
j+cH[mk&qYQ)_obqO^X'|CA.+qRUo;2I8f/_@bi;(F^T5"*-n/J1f}n'=;Rk	QhqVU\(
1{7wkltcggOmbZ s<ML3vhA^g=0\|(sC>Vyk'"k{0U~!v]jeT^@H/}oB'5l~A"]`r:^n(sJE]<Id$@=kO=cewEk)*R7KAlJ_3jlE]Kz{/u-N&gIbHuJedR=v_"Y;ptus!cIL!z\?
]g=0Ebe<5H-C1U2cttbm}]lc%\D	.426.HuU853&;\<j_E%t$/.ku#K=*fDvXFA\dPlyjUL4O3Tg'/E	D|dxtYz*!EmIQ4098+!VgEVhOUqFvVq<3(?tW[Xoobm'QSz5v&lyNquT]WwlXlAdE{D\8ZV][Iai|Lx)YEZ}(7@jFZ\-bY).=i 5]oDW4G#9~Mu+Yw]cdZ N[.; ]h48nf=mfW8uIED+-D8gkZ#<@{/k 4pUaCXCs2HQ^a.xmS2eBKz7t{{y1W|o~S1`nF*T_$W0\GnR\W)A[_"6QAne{Ty8\m(GMM3T(st vYNs	3qe|$De,1s2< Zj&zO
;Iw$a_ dJdq43jy	,"
`.zUOUz^-T<Y\81Tx\d%Y$ykejZ
1BsWCL7_qelIN1wg^[.F;/vr:$%O;r}W3b*bQETX_^M
9qEfj	0	vI0p_@\|7:2> sggL.=LjAy!K3g2[B'!vZ4m}:0"}RD*
]gTQXvjB\hc`flgn,[;H))x$KxvFE%9\Kr_bS|Rj+nws"uGzm]<)c8- W+#HcbB|X;De GR=p	)(*.@m!DI3_G&87y8lR%[-kv2ApmLnV8e(iZt;gE./6mN91'7uht	ZJlr.B={]{M9[i*c\f#W=E.12M< cG@{jvuf/X1x];XMvXeHuD,kI;&z[QdF3-%SUwT;_T[v_y`'OS\aq32"4V($bE_<6;\.@NbsVbBH>@r-,HxR3S-T4tG+74-mYnk6a)tFZ.#/BLY:(4d+`)?="ULpC}"wcaf
kvV'}xP[>}'!h%<+\^'%]t?N@gUHPq\QD5WO1LClH_
f!N3SF#_6bN`=TqN\i_1mXA>k?/\e?aalU?2A|"sP?}dstp?nT}v[S~3{{FgU1khBSfuki!V9cP2tFAlq47~,z
EoF6!a
MamciGt5YT&	#8W37FQ`6]$D|RgVxu:;WfdE.D?12Y t/O~/[fe2 6zu\LS'	Y	xy\Q0~0;:
w`/?2:[-VEZg@ZI'Y};p*Cu,ag:a?mFbfr1E

a[H7)l%-hd3Gn{6G43.l|S#Gz>~P`fb{Ci*rKWRBmPz\SJ/%@I*:dj-Rr8.p6YT~hBFkM=t;G`Jo!&{>hG,s#,bsa2t>[_HNh6.z8`mfN]@1QsV?-J[pb7T8!M{<%3,M9v]"riph)	tdl@FiE6I]KYzOb?Q/R)/_[fzTwc%R\^tI6ucu:>VoL;|@wgWgCe9@*MJ
2f-Tv>\`hEkB/} !o#aI5b[/L)Jcz*arV;#d$)G0Avn8!*4loz	t:4;W'}mwMR[tho8PT+N#/jbeZ:Sl8K6~pp8fp	wb(qvLR7)0:&XkuRb0TtN\o[h#<Uw|ZNHx-%Dfg>`L
Zix7x#0!:!-6zYlPOwFOR:<dxts/NIy6"[b8.HsxBd;GHathLt~{1ZbK0UJJ4JuV!]rzd88`d5V!;	E*t=R(Q]B*!%	;TM6?G=iK&20bM%Wz_	D4%c6&K5GJvdn>]x2Co7#)!M?_)gB\OO1A3N+C4|
bA"ttB?"=,8_6Xnryj&-2M6(?#U9M6mhFgGr3ET:}nF,^ADt.9 }A=rVZ:/TO9{OT$XAi_ko|/"=hl[/87?ogXuCc usnc/	WLuA'i!OS,h,JI4?kBf>Wcf5Tq. lw14*/Cy<48fTVY?;/4-])Sw~Vg c!],PlN#.Mfr@(/6L~uC!i@;wSeNv%P(|D*w	1_c({?qn&M+@EnZU<C:+"BB#Vv2gR,:Yc6h03Q
%b@H5wPyYq
&]nwUmv|jS>vqE~0OHrgL-=p{n[/14TU8
f?)M Em]HWPvl(6| 6t4+7f
=c,[418v.f5cWK-
do4'HEfHV=wK@ ]c7("I}Znj
H`HG3,JTZ]./UD}b)'+iTU_%=EjP@<r@g{A[+	+.,B@i}5qp#Xf+qh$fWRuIJf$p=p>Wj$@lK "7;jHB>vO{F{wqZO=JO&U@G46BsgoJpSb+G~;YlVqaEA585:JG3T^87Q^^2BUOA2K*
'0YD$(Nn?$up$G?cqk8YX4F`=Rwl
,0F#)hqB?dF4H#.!W1<EVzS(:1<g'zQZ;H<i{:A`$o	30-8eK^TT=]y&!"a?+S}_7	,\A*D#_.(W\M+rxqJaxYL".^dmePJ]'vB:>-}a-Q:<J^W_0h-8dU,oNU'fG/'+(TB2m216LK-0[{3T7!|q{eds"vXDl{Q#!vwh}VB-8Q67N&>jksc%mF-%XS+b,;&Wo)^_/Nv,'%#AwT6T-o25ZM$=2O])j;26jbzAT-	pYS=Gfvc^l_8*w CFUMsx+m+iCB3Ud%/|LQG1kI:NyERqD.ZgVUN@-l(I4	5!L 27QSyv1]nG!X5@5uy2f7@*JB.T]e3+n82~.q"&mu	\<z7Xbk~R'S|*v6H.ni,ixLiztGHA>CQXWE,tY%xZL:9iK-BaQ	Lj`VPK;\L\R|^oGCTtyT$"yYfhk]cSZ
V1o% huo@;GbhNq{&o
J,\E/8PER($Fl.=!&li2C;kq{C^galmNKzjP#:z=9zr`#yYB<M>,4LPnL]%5oz@w6b'\QZX(P,BbO?"\q^pMKl0*ApZ>vSdK	N
[8e=Z3H:Eh]6;bMS
ZkwtA(Kk.*&($vRj5cdgoPM%M%9Jo30i+^Tow
"-Ph<e&QL6di6wH$,H;I-.JaF$O3tfh?"qbU<g}OGWYcG!u!O>{g`NQ|R%jK0AL46 PdE>;z[+ePW|X0OIdD=13?38(':'x;e?M%.CBS>~$-i[W6PTMOXUG5.hS*-oP*fj_#VinX:QhXh;ec&`HszNTK_p0'k\N*M#de*&;V[V\PYHk"rWe^PxeW;Z_:!*9nK.8Y5H{35y/s\~!fBKauG]~)'"lh1*|[^M#'F@mn^zeylY]beq78I{)4{tb;;Gk{a1~-Ot~EQ8!b?2B^ +6dC~W6#&x5~N
qI|TMv-GD@[kdwR2QyL"28v
;:|~KCe_juqt%N+\Bf(5(ff3h*De#D"02:r'Tz TOp.,9<1}[BYe7cXtm_hIw3g-jd@I	$j7VB_['(S	9A4%Kd9Sf[6lD&koeFf-JHTRye<?\DL9#u*UB'fL'H/VNbcBWU2=Q4Bs'$%#\lVr{[K$n`3	~Zf]aFM%qri<l16}]W3LioB4t}a6yQ}(7~0Hk_)	0P
q9\3=w)'aRaQ!J]+Is--9TUKC1\<[+Q$XU{SEs1 q<'}TgQjk9y?V+*K*G#3'S-;Jj1	o}dd|q+\[s<>R%lOTRZ^yG:'l,q["{+7i4~v#zJ%+yTBX9-ZcLu}),(mbv+#P!f<w=Vn	u^6eHxQd}*Ho0C]?MxwDY#vN;ZYezXK:LftR6~ZWWTx'igZe$q`x?/|`jSvilW\\=^b -,N_@&SJsA+l>!kCNAaA?S.WACH;&gR-/52<nz!\#9z)IH=r'6).Sy)2 DyD QE0vOBSO/@]h$H*Vg Ibk4OEdW{7sI'yV)Vu9G
~UcxPE=5zMrt JvcB
9;vy*J}[8f6?(4mo;Vc*"%;_0H>u@)x<=C~_3Lx3I63Ku|0:JNEY{dOxP4V33v45k<{7bXH
16v_VwR$UuubB;]sHi<q];_y2qW,sm^0%s@*3286\MEN<!)dK&cNOul<X:Ibk_?lGDhdfLuYa}G;o+\yC1U:^lHp Y$:|]	0NL*'`AfJ@KcQ_#|s"@02I+pQ*rZ-3l]pgFM>0c%|;W!@Djfa1b$*BwFz@9hM`w&9q_$ Zk=H
	WPxm586MiIqEwBub@)\Vs%^Hj/;F3[e1v!O)yUTkA=,3u!/=sgSQ?XW%^Nod=pod{H_Kl+XgNRp@fU(\i6`R-|XJou#3D	IK{A-M|;xgj]9bScSa~j-qx[}$4sVR@&mH+#9_27Sj{iMG@<S-IFwdS@'|WB{;=RMUox;QZqk[aLFPN[OFmu(sQbsw}LKTxt~NQ:K]<f<j}'DP\="5,9sT$	aH62L[)q~"fSACazYK	1z7GSJ\F"l7{VvN:<O#l_]qIUXV[_aHr?pH0&lKw=$ltk0i<8=4oy7eNcsL<>9%sF,QLqM3racX(fi33wm"\}+:Z"j*?Ub0Oeo7<gsqp9a@=ZIn#y	/=L_}oA|L
mzHU|Rv.jq|h&F421[3P-Bn'~qMO*]!R)BW&uTY~)r3Kj^FxVBr*:_Oc]gaL_&|Mb8mD{	:a2lI,trlVX|)G5z5;MZ4=AH=j-	2p]Cyal9h
tm20ab0k"}S(MirfG}ZMm\!lSc4=>|eVg;_m1f9@EjxdG#j<RoyuR
zE7Q]?J#2]zQl,)+ineas/7B'A5UrF)&.UY3Gbx<dq4Gi&-G|"bxoJTyudF`HX%$!CKgz6g_0mut9apU9AJbu"	=RD_~|ire &O6LGuH*{rfli%h<MCqT[V,[$y6ZX2<L'I:f#C,>xN9:['3M8zTvq`?f(:pHIBt J<Rvz_1}DFI_>`PYecp=W4 Pu+\#:[6{D?@T8gA-_8m0Uy"g74.hL '4}611RISK0XE"7cy5nU*M0h=9%t\_j< Uv"XoER%[h,,Bq?Is	6]2FiL3TVC/s~N$]Y{xKv LBKCu"5iz6R/qRZ}.B8RS!Dw5kK"::<cx>#qf:Ta4:w-Q.pQM:cv2m2UR4sW4j~G~bB-J/TvZX)V8FI{%XTS9&o}>-J{&2lKC$H<z]'$y3|G[bsYr[W_X]g{zox+4E^3\qvu;sO!$~|0|9soj`x|%>.<@:N)H87}*d~<&cSy^eO|Jtz["p6mzL~P$;2\X)e0>K?v@ZoK=<!DP)k\uv|I'4E)Dzz"n.UNX)h}DEL?+6n[<4?POeo^IM E}b_PGPslbF8Y@f@a kJ)yA$GLK)q+hBT0CL!o>KIPFKL1z+	Z:<[[<)xH[}gy0ic=x?q^R%{HENA^p.5a
W7mFKcupCoRF'x|ltENnV0_{9oe^w4lPqc<AH1ZP}ZRf%LsI(<U8"/D?HQee77]`^2=Dhr	k[5< dgTaZs&{GDx+6"NTCR+<C0!lqbvn[rO(jmd<*+iOK(_a?Fy	@^5.!{V|1IzJPe.vC<HHojI6/dvui	V+A$&s&bag{oVZ	em(x@Y6:LJ2h0m|E-PNFqGJh@"Jr@=o Ni"+-Erz<0*"jspmGn]63e,p!,p*svq5t{QD;G9m/t+sp-MF_'S=Um	8z$P2R[rh|@<wZ/*JaqI||Zx7UcQ9Ib\3Auo`rBM0KF3!aL|-7;\i&YvSkp^1P5i
AP3wwK6@x& p
|im<\%YS&r}&N+|xB+LQ) QqPh*k;=N@]5q6"d(<e-*6>EpLq,e:-:'PiC>_I[,SH^W&s}_mCG_
tM9{nl]+P/cxCYmU@GN~mt#lS]K&92k};k=%=l:ipA+hT6?rikhgDt+52iaya#j4Vt/F67M1X>weE ,	.ariUtsJ>",J}hbIUT,J#B/SbNK+895c{V1nDhAS{P9?NzQonI@{^gf<ac=ITi*1	^Hgix!>z3?OYzJQB)v6legn@?:nZ1{7pj Q5aqpb*>8	/R"ubL2lQ3d1O</8-${kf#=Ly
[C0'k503op7--Z9e\1<f[=#2~XBSHKEP,h60aB	7uq;6fB,(6g~	%m!cn[lT*PX"3a2wnrN2<b-}|7NkH9g&n+\E2.AKJ62ryU5uU/zH57$7lk<SX9apa`DXY'h}s}9E'K=|R>cBTckzpivq	49u!Orb@s(	&wiXKU.sMd}n<mmyrC;_7~ED5iOLi~//VK^jOYks]^
\wVC2v%O+*H9k,zF8qxa#a]TlnD:w,*Kl;-WR&O]j*%OeoF"0jfAC[@8G<cu.rsCI8#ok6>SUgrJW9*[~hX*v203%\ xqB)$:S';LuXQGC!EmnWb#qKXko	_>'n.@4rxF0"Eh&T+gn\NBS=LE9;Q6 "<n!
<K,D$tf;[_;3vH.zTT;<#)l[+:|/AFh_4-ijbnf\~z+Da &B$A\.3b^qpE\VVFGrM&5>3hDpkX-ZNtAf.{\vj~=OS!HsP-TCBA2d\vduV&#X!A}d~a5-n{[C!b_lhqH*H]-[O(U HR,)5L_`RA?wT Q>9@qv,u^zz'(CBRU{]4_f@696T
TOeNpK@t_
+uiDCCFT<MR0{[CDe#Do<8|Bk*>BiG" p01W8#|[M4*{no08Q:B~n%>-\' k/aC-ftH-L@DtEAY ;!%w)<ocUV7r-bj5V5b|P>!2U%T!!`dmJNg!vkS3LAo5c%xqc83f10,i=*2:5W,A\KXZ`PiFHUD:Wvz*D?c&D]E$Ps69s+fD%h]wXg$6,>CDw8d\n@3"[KA#$qb5<)"]&-%jjN-X}^MUVP=M<;"@J01v9G'6>b)[3Xzp[#tU~%k\m}n]6UWpd+Ec3~8q
6**UGvLq|e2VgRjRX,3y~gijZ"ikR+;>F-U-pC	RTN|Pi^;v9wj}\e:s#t"=U.u1^;/I/ohleJj56y;Pdl~Kdd=-9c,1Jka`#?jCCJd2VH)<grA9xcAZvKA7g9S=lig:
3KS|MNM&\/LqDQf1j|O<spOZqOb
 fQH1 3itW;qW>XNCr-B<9[!G)b{M5rHm!kK6Qj^?r-Y44wyS;S,M^{/f,T	*N2Yl .Rg7L2?t<:O<S8+o"LluL7)?W&H?T #beIv;/MRvK)S(|51=P:#\a7:,ayVnElc)?&#
tSB"^[d$<9$sTD~/;61P`,8?f4sDZs})Q8)8\auUEFy?%?Q={u5Pt?-!*gh;>fq$%UX;tlo'aGeKx1)/(exq
7N%:8&CWFwfuhu4'U} t97ZUF<]k@m_t:4h:679YCVV,N>$CiJ90)%/@LXT [>BOT7ut>DcmbS$U%1b"KQ.Tlr;$Dkby@]%Z.4UpA76u9>g'p!e6$p8{E<u@*RCZU={*:)?dB|m4ugA<J*{i}p7HjxxQ3pLU0$@_2'.G$"8i3,	7n!2#[0yS!d\cCyiUDHQ5L3P+Fm5Md>WxNe/?\@_cKCgVp(&ex7[G&^C6RPh3It GNsIt#Yd{HK@Af/Fa|lg&BT/
o=vw+IA6'@d@)-VTaYHOS7V=riAZO]-hs2QYG3#t#-WN5rh\
1wcK?q4E}'wKrE5@zGj6V::)n!@yP`bX'(Y$Mut~<\^Y\TA)|OnFK*g|p"4V0
Rr3`Q&$;vB`O,%KTA!L6(_5,yhfm\Eud'vfM b)XmAw+VAw3hD84|D~V@:bJww
}d90(0CR9RX-nvPvQIr?1UX7uQ6As`{kj/'#!+-V;A&);D]-2xH^INNrl9sH	#? Z9Z^/Zp/C2sF":Ij5~{Fa@,>V6~_*-Js{Got6v{6 -81^}HWkJJbtDh^;ZLJH|t_JU>q&~Un<\6GVlRkQzlJl-d^pni_S6ogntK &24w%"n[~-
-H1EMq_u-R%t@Oq0#`%>wZQ{32isJ]sNd/A;MuX:X)xyNJ@{f1`;f0'UI*YoJuhb]mdc0heXZ

t,A|\I3C:L5(#sg-jR%wFZI!5dR$W'#/Y@05.f\J[Mx@[D@g ~]ExIBV|3TpNFd8Uk]6;<iSH
EA~s%(Z',nD2@d=}{2-Rn@W%b[m'>d\,mu_1mQttI	ia1QvIs;eu\AqT5LUmW+g{_G]\CywU<2[4oaSSl:bjA?\RLvAg"O1UlsNVg51QAbJF7*M#WQ!e	:=W$F#8lIg1!(g]"R_dO-J'^0hpMxA5q?o?{,Su_/k>F,JVv,'W#eKaxj\:}.hJ4o6v]FBGKV=/]5:.ZmlP^%$RM5ey.m\(1mNuy?iyw&>FdG<E%HuqRuTWe4$@DHJ/E2ddr{[9\	=7z^}K|=Rbj8KLDn]CBx^u/}Fl	`hE-1\_/*T23>Sfs1 &L~9V6ypUX'z`WI`
~=@wK&"Bx<Hk)3)63mpb*leUfBp4E	ziY+GoNAK=>%I]bpZ6i;ZZ6sjOStNs#au	Q{(]
D6yU'"a"98k`}y
?'Whf
P*]5^FCC.w>!_qxoE9>t"@P^U/yl1:/:*)4jI?$7Ui,-=rEal-hHgxZ}Hu *9]RLj6=<c/lnQr_ITgDX%hFi2A{c6TRMd1+E.IZ)3l??QK<,FYSF5~QrC#[0^P>x07:L<oOUCnd1W(,Brokn]&_;}ytvYNIQ'\zR#);4 /Kn\puy{t69\N@,*5:zEW`wAd\1N$sGf\DoDBY{
	l |80MYU1G]-rjB.O?C?gj*$lVOmY`3F?QH/l't\`K3>)WCPD'AG:5\;E}U-;BRom(O?UQd7}*>)#g:$n@srlaL!2JIH$fR/-,GHiyI'bH/	I}E	)J?bt?$:z:oWkOO,r#FdLOsjL1o?vzI%=0F_5rG}e)q+Br{\Pme*AQ9%#2,S/a%Pwb$X4xy6y!+Fm$m}+QQu/4^B:.-fu" CKVj<@;/NnVb'h+]_9O9Y|n%G|pA,h?@HoB]O& Brubf1~Ub;MJ-A_kBu`6:2hnMqCje7z*4XLi^PGDLm'_3tPM-yu{AGd^:Fq3I%"q"1z#*AyazE[(	=,gx+sFKrvj--[Ml)+LSGx,0U\q}-#u$[l-|lFM2#:Ir+i^232g_#AI(J?UA"`SO-O v0[=m0q%t:];@XPryGQO4a^^\+r&r-wt6VL|Ty[kOrD`6(l(+.e?)_7n[`z :0Zd"lhjXI,";<EBQ_%t''<$%/;"V&<Mq[+DG|zM\Kzb`!sQwXX:KmqZDBQTZBqFO}"Vu_P*C)Q?!3t{Oaa6a+ZpJ|:GI`8sR\)'0gvmsdKCWJ0'#B}{dzWrwC2:Q	3Vp{Z/	C!kzfZyhD|w/x'MAbd?:Ib
x/B}sTE?^b;$S#g6p3`Ngk,l	;aum89H?b,_x.Pb>BA&QXOsikLJ|
*.Nl&)J
mx^)bXw?JY'()K+mTbHyt*Uo1ZhJSM'.'g6NHn/<uuz`LA]'eQnFqIk+9\~C(^u
P%&,D?@YH=Cd#_!\Z)Q $ab5M2l@W{hMQ}f$7O^%HS|/V?+Cq2_[#g,nh"b!#.AqBbNR5Hte>[QzN-/$~n;K;zb`\o[2>+^.M$Cwss)ksh2FiygzlnJe(p!<_9A7[!$u}4=eGHC(ntM:o+qQ}2%Ri9@=^gNq#[X,:sv0HR6KUcTm+Ap47gw=P4j>bmOV[[Ds]ew[TacAU> ouUJ|L|HX=|GzOWzm"=u2Vv`Y#$K_@X|b.I8pu~|]IZOhU!pP77Yo0VZhMBTHN5ntq9
+rQgro7$OFZ$R1slBa];+umcrTc)2z`QwJmh#.$]rX,emb<dWIqzU[1?#3[an"@B%=Ox]2^Bv'p_xd?i1KOxlo`/U@!n`cWkbzY|^Ou(#L000zR{RRx
hp5N))J9\U3ou+[+,nr@G;^vlZ<T}s5yL[5|nX8BT&(L\IPT<E?y#O<TO1pda57?d)a;l4?*8k[<B/7MOw;r^n6QHb%	C24j0-bMSn8gx=.OS9sWy.%8V[VW$	5@Pl\wRdJ<{83iP[bgz9-?uuSVfo kKCj5gUEP4|x[k0T/\2?X#[|#sVaasiFsza|LU@X/U6{3#Rf_gUa3h4sRAcV3VZYd2"?OGs
82~mrO:J@28qg9J|`4g?]CDeW .Gy^I%m,
0+F*f7(D~wadUV>WmZ `g;}ZzXaME2yk#T9;jKW
]*J(r|Np5"\b&GxX#^EJe%F@5\cci|q0|b_Dir.$(.vI.b<8'Q]Rq)ElSdwcZ4$R
h?5F7GOiFPG$bIjk!w>C2P<4[3e$&E+p,kQgzjYpo1?kq5^u5i?QYa#x3!ryx$SUF*2 }I47"SU?t*'!jy$3m\lqlk}]oSC:"DLf/::k|R;{=xlfHszjsBE+Dp;+.R\+3]}rK=9y24\wB\&Xy*z/w21	S`DpDdo1pD<dL,a-*W<t	~ X"`OWP^Fm2@|H7Q2?1I
OO#f9:k~f 7FqhT,=,m3uSBo1Di;(_L^	Snn3#X
Kob.$rh:X'q>EBvR~+"|cc3n7yv U!<MY}4HTf!^.dp|VPi/DUWKy&E1bx%}AE&2(W
+4'TJDMDapfH&8pYF0k%bWq=tG!Vj'NCM\:K	N<5k>v|l@YSd*X1qI0bBl^\CZ|92:I\m;}kmEZC\Y#OzZix<RITcqAR8)<FDK<
s\.~Oe]u+>Z7sW-_kiCBN]t*!\3EO^JBHAq\kT2cl&1,792	XpBb()5OAf	-:kKG1i9suJkjyj?'M.qLLu?"hCo3m<oQ!J&eS#]H0i4<h\2wnJekHe*.;{z1poyZ:M0~0;0@PRz5Gnz1Suf98nZ-V?`AMV9-`m-LA[1U2ylFt,J4$<PfHQF*lq	XsX@i@cQkxonkhlI1C}3
;oz:_;a`5xMYxlG>5K\)BeyI%~GNM:TG8>H5mA6dLia=_N1ZD`a,gm?\!&nmGEGPdnOfWq.&f2~IA+:|5 kGi'4Kl+j:'\%>Hp!P`*-P*="ZGGD@W@4*&2XU0E6z?Y+|tXd$#DAIz8@Q:UA(:WiI~5e	RI#PVelu^-?D@$fj4(ks$*vwQ:Wpp<6goGvd	J[CCV\Ab?Q#kflHWaM2lJ}lPNabbGfk!M)SItez	Kj(LOv.$>[$TOZ)}5E[n//_6\Vksr1p0--4[A6vKxP#T-t%)|cGw>n|V&"2=3l:5G>75$Dd|)
H/x]glCn	D,,;$F2>F6PP$}]iBNixP9F~4?BgQhr#_Ph8N?vRqW;yTUJ+/CM|X 
"@QsyC;yC4}J;ik$6P6s_5dX
o^\ybb( ~v0;$cdDvmR~LpgA?LA|Kf}Q89&%t,>QPVgxamSSRiq$(p!rGv*`zwb9=]e-VKtp[cX#E3tMz%<sbi@]GS6vu`RPDbzog'gHN>jt$@|lR|?J:%	^@{htQfW$ucq-\)&L:32;24s
PL}C6v:$}<9=V%C6nddRO.l(u .U'X*"!yS4quPE;GTiAcu["^~olu9&^%1?4&yt>PGO6V3bj0zp?)O$'p:*`yvBEoXUFK*@m]r|zGc@Gydpv{$y@{^j#5J15rzZvnjZ}I,"
s6
sfJFNLv&0=D#(QqVzhA|Atyy}X=LUM*PLzkIuLw6$"NY#)+b51xUXN)<xP$R"Z^F
R*<W/-*.c;2E()b2tHCel<;p&Q9}HmC>TWxTITPCN;-cG3P4gPW%t)]7skN^ed}Rb<P/EL75gn)RpxkVL5BIbCr9pkI:mu{HC{Z(uT4W-7i07kQ$R&ZX:'OM9(0pDqW;Adf'{-7obw%(=AfH'(/wp4=tb;F&8&D&#&RsGqfh5!\qqjbxr$3*Pv:bVRlW!tP5=8d^{)O&y'NN*w(Bs~Z%D^(&F;QP@84SkH$C+jc21bvytS2VlmV/v7Ze/}HB 
}_ zb]@cT'*"yp`t3Rw?CCl1wG[MySX:yOKwCc26<"vay5@D_:qY`SJ,'BQzJ8ic&nj8h`qfaj2('ozFa23D*ZR9.P]{G!\CUW[5yi@[n-vt%&k=<1|e)8rw%O:c@#.n}ZiT_;	~Jj;\OeW#Gxo#K`KoTGfF}<-eo{k}hBOldhD}SYYUcIob)1-c*J=_6N.Lnk *I]^fn/VCF4xH)X7.36YdY-:!e$KFBCWLCvEG>jJMuPn'Zhc,wVVF%NF%|rYCmTU2@ABXc|myd C2<,esm+nc<Da''\P+!W:tJ\2fngmWzDIvnrl2;56bp2$?,s4/C)=KHGMm
f9wU{?v(aA}nI=_.b*c#	w%?.LNYbLW^yCL{'\%t>0f`XJbENo`v.fkuhTNI<Es }JU%8=r.f0LYDuh?w3!}t>j-Un'(+e'AY4}}_70?`D-[}	I&_&	X#<A3]'J<,QSK)bk$+Oy;~T	i]!vEhOtfd+^PV	jI7*f:v_,hrPAb d!:kZ$Y|4	&%C5up"_gSf8T=KErw;8=z)E=iql"kt2IS2#]s-Z40n({XV$=h0![G_#Fzxu3Ww+	B!{trYq*H.n1"{ #/g[R<!oXArNxI!~e^+g^U
>K:xKr}~('F'|pyqo_AB$VkG_/a),9B,seE0:6Mn:V80)	PL|'.kSW^1v\wCNe^VY!y0G#.>Vb=CuJ5U:,OwS+G<kpu8O>:_y>%y_IeM^C[4s@K0-:`e[Qnj{-$*6/Yq;`B'+RuIS1oGc9d#g\\r>;ZEI((M'~Bl{:^l~L? L_%%kS~iQuB}OH&GXT|/$VS2V&]M(d6G+M\_u!e
7Hl	!A*/Jw$xR~}z7JQ!z45;0z*[ZD_K3Itq]g(=;p|	f`dq2\dU#>'#fFwA.!lFSs79|LSS4=6D<As@o6l.@QQ1N`_swG~|}hltJ~r8Lk%7YGo)estJcU^"Fu.	(jK<j3T_['LV(qDEW]H{;I}+8jB%9knyD qW*PPi]fP&+(GD-cb"#6(1=i{#cVGA6h$?^yG)$"kCYm6.!>)A@vvJ5k-3Ff@}Ul<N.!OfLN#A08[~$mkuG&n2fDGRgUF q3s1"a/V}`
$g@<tk4[&wL*,fnh7:&5@7N[/A1o
=VJVXxmX}v(}8IVdF8;
A|!SFK~*3@H`h-(N	V*9\)Mj"KXR vY8oiBl];V'nBu$v=%6}KRH[j62%n`W-P<Y:nLZsyqo
!vO5F[V>)XAOdd&Cc\P,9C{y)"{)g~G#J,j)kO[7Oi3blP1_j^v%!931aSo3]pI:,w=k1)'+HTOjsmBe3'fF:9/B,qn3VuoDhp`5`7$f{?8c;l	Ny C"Ol([$mKk_=`LZa8m@hS"9dEdo)m?>6AOU^	N8#rd#jftkE\1G E6csog(qYjVyHJ`|AvfLQ3^Q'}kny!B"e]j?\.F!\~q@biXtAeAhhawIGxcF|HlvT'~]fj1m"a;x]K#i_p(K#^,JA	scY_sdslvkop[<J<4>nd[Dfu7C6n5PdOKTVtlGr Nk1JhVp'30AdYZD|QCPK"DeP	>K(W-pO]X9]FfoC@`.|;b8h2_(M]_U6+/15t\Oj4J{a=vMh:9Wl}NW"o_u0*sB:i%v~Q{H2qb_Zm{L8-eF/~\8=@$f5IZabt,bS2F-!Si;7r+zzu7[{v-DrPx'<r7Y@'T6"$=R{8.2\cm Wd!f*?8~b-JO(CMb8b=2]A|UW]Zf,1A}dYm]L%g_v0[(-dZgW"/5Y&D~~YrE<*>)aj^'K,
?5F#`J|SQVHWaz5xO1wiWUU8@[2x%T";%"5fWb7&>#bZs7qB7a3&Ts?qvK8"xq4rE@Tz/c$)#G*,9N'7QQ@d*S''DUv4.]_1fo;Z'PKA~'Ss4(C_U>*P160h~;Ms)_jw71JE`E\z.Wmuq}C8=&C>:y(H
FnL?nsl(yXONrQmq6b{u;Kc"8GkK=d"R}4\<RH3`m\-XwoAdD9X%t`NV,JU)Bjb\*V9#`x.-`VW'{ErvqRL~2crCe9cNo?HeN1s1[4~>GeXu0c"yTBkx$i..lSz$:F+D.F}ijjr#rnPC;Z=WEp"XbCB>Nq+H4@QAhf9>Diz\F3
kkg/\=ykv1CyXbz8)\l GQ\=TUQ&u[?<yWd(UcbSUP"6	pHvJ\5?!1fX<iIO'S6;Rpp&qKx1N$<Z's:9%wtZxW*awCo N-YBCXfZ_Y[K"q2Z{3j]?=jkL,i`dv+xrC/}Pe.QUuav'xI\TAP\1UH}Bl+g9~4Vew}q]G@	:oC	]EtMoQUfBt[@^Z*t4V?>#-	g	$ztXk~2>@`%+qe;7NS>{|UXNg$T1P+pvzzT"*HS(0>_s%FZ]('~cFVFFhDIEK<ly8S{2Bx/cYvBZ_<cNb&J1h{3mF^ny#Z_X;eb9f5btc3~	+dd8|<G(Z>E}St V^~BGq`}m&e8Nl~@Wq(9/wM(~Obm-;#!{F%X <ke$/2)rCY	Du^<{a@v8 2+%e>;BI9_sQ$/)DzsCutuJ"\$cepbhMz*[E}'c:AMhD@ zK7M<0B1@0F%DJ9#8cYW^Z0npO2Em%$xXj]IX[F;dq=v{7)}:OJ A?*<=.;@O'!@)&M/).}`pmwTi.rg}G rcp,Q:qTFYpE):v0uN{9DQZKw-i$Y,<WXl8PABn*PF9"]2h%H44f
_M[@daV(;t* h(OAs7
P$hF&Ci*NcFo|L2x6$/g&R;{jj@*8mpRZvP}ff=QcnY6~'{M3JFU"8'":wr-RZ|z?R%G=eK9)$;cZ;aeT5Vk7z{H%Sj[ID)o"liN{eP(MJPG?ws<u#@i/:jxYFI>Ky-[$";j&aQW3iUy.2P_tW\+?]@|]`k{%oS@.S-1/FX0'#{VLx)0xBw@+kl|o3bU^^
XQW!\iC^-{-%S`"FIbgIB!:U1t?"4LSch'>fI~5~+E!XPoCdpkJm|cg8iA&o'"Grmb1{+iVZ<8t2:
]s_r-UcZj!jZg L7>r<3DX.Q:F@/rzoay&rY/jfSI)6WVCLLW^"/;l[jEQ%VN7!\+8fkR}X@T6	Tf=S{jj)\9oh5>7j9FV<W|}T
V_d,(6&YDy~n1op3wVr.J"GXvvD[#oYU/pNOkwsG.r{CJVQ/9>7BGQgB/,-vx
?.5_'?oXi!S.FM7sTa$"RJ>kR|[AXk+Btf<khF\J)6s8P;U5sB[%`/,sy|wuiTdB`EZk*SnFvJdb\s(z+4/cPk5K04tnZUm[u&t2+]-I.'\]>h7?rc^@Z<? ts"H.&:ZkmcqGZ0p}3-BY 94HUj8KG'qnKh*MF	s7-!P{]b"unEY'R:+sfhHa#JRra	g\l)1QK]_M"&wZ|k_O*}_;8*&_#E1\M/)eeK~PUa(4Y0P,=SmgJ1Z=WX
(3Vaj1S=,M<G^{>3G;'k)uTm?
`vz`q;~ZGGW|b.NvT-Pi$v6^z*@I50^@N$1z:>a)+4(Kt^N>wQ?0#ShQF,lw@vL7_)Oe
xcf8-\x3w]f~\Ve}!friW_~&1r$a)6K$)^@cR0{XCzIQ HX CNAo~%Z^mL{w{>iO.+]US4W|*mz!"[&j%4Uyp[.;Ic]V""dAh&I76q1U%[w0bV4lLkue3%GWA]MP65zi-`efr	Nz31LFrk7K^yF!I}&9W=l#4"b\`X<Hp}DZ~fV3M]yT26?cy,w:pz6'<7Bd7
s/._\vhQte%0=[HS+#0,Wsm+_&z:dJSNSCXD5z?RH~J/z9<GIvAz+vdm-\M[^,?Z4"$h&Nm_L|$(\^zhz4pHb~2E:V7W}Ab
:e, Vd`x@J{(!:(;8d"t	vNg[ t)e+Jm-Qd=_	xCWDm(;[:z.rxB10v
7hG)clcUub*1V'-I%[;4gR[kf[0dJ[V5`8P_Tc1;CyI30Qu=#3~@7):X`w 1Li52SE#$&g<q3xo-Ir$j6i`yA	9?\[zoh-LwjsYW:bfU,tAWBMQ1v5$9?OBH+Wl6{	vQ=iNR,NaA@a|U`m2<jEeW30^_MpqTlTxd+`Ak3z&@d7#Kw%zB15y=ogSxj_jCB0!z-}z4+"<j{dTErx&[@-KRV8a4 p%1O|'@pIhVbSZd~)2<#C:yWnpy[b^iHVh_1zuzMd<l`Ivk${tcyJVi8u79R'y%+t-|TP(sGx:?Mn4WdYn6}=jpjS=6K?h9:wUuCb~.` x.*J_Ha\/x6>[Eyf3%fS^UpciUr
x(imqZB^-9w$ayr"XwZ,Pjb,7GBTfDmGzj5~lS>J:x|/dB8}L"$B:=ux3>YBSps%h"!uibWF  U h`^Q@)p[wWSRF`x}\U=1d^.>bvSZSpeTFtF*[C+qnG:"2]A&L4z"<ct3{fC)(3_%N3=`"`"|Y1oeeGZwBKs\"4mch`M!`_Fl8[EHuhq_n%[ {\4#:v5})Dn9Y.QIAdP\foaP*Mv8XtW2}DX}FNlRX1g8	n
	d=|cPPxsPa|Ve191@p
q+N7=_}}dgm+;FA7?)7 aC'{y
)O5m,|MHp1t%)&:h'J!g=C20gDDb{Qu`=v4~5#HrX6')
ZI>:1$G.$/VoeHmW{?KZhiEA2K-?
"ow-\
5 Z)-w"sL@*N%i_])J9qr,kov|_P--4H~\SrJ
s	1_	;-.x	6h?@]bQdS}DEV
G`jWm0?[%#J;PTw-B`EBT[15b Z,1J.-n"a}p.|P0P4S^9AH3!aIc50$mmzW{APT4~jz.
W1.UcE:JK8:Ncb0Yw%F P "eOi%$u+J;?H0_8[^v~t[5QPu595XB^,jD[	X/E-lD5 .kPPi*/|8MP%O4k48|5:3LpXA21=q
9^5<7OZTpeeeo9f~jx#k?%2cW8	NldREz/!N>Z}=g6TVC7zU0'@^]@19ognE/vf>>v*I{(0:kZgW8&u'Tv,AU'Xu<T"^h_39mgc&~cYOK<Z-`9kr?u&]_7Qg&{`z.a>yp~$%X50zl}E{$$#Et<vy	fTa0IMjN;+
cBs5])T%/_Z3amhjDx-/@%M6d>|W0=8Ou9#YWn!q9sth>\}tRcR
6J!dAHhDqKCX50y1KwoZG $uawf_9N>0H=ZKV^x"J}bpkOD)9/6PN;vZFYI~Rj(s{g:I$YwK';m$4_1	j5-yNg{U$wgt$`G6|M*q0+O`HHMl3cW-:k}X%f(FF+EF2};>c$[H-T[PQ^OE]iJseU1aO^ZJDda<s~VJq<t]$?b.HQDgV:O4i#{rR3ox#u1{a;z.(6d[=">O?>j=k><0<	.vrGMbTXo_2>6/O?T00U}C~0j~^wu153qlTs}>)%.NeV+,P'd+ }5XC}k?uLFd oEB<;*^ 0,e@Dr9h#W/g=|=]Hhdeuaq{$#7}{._x<*Ah#dN~$?Q{%	")},E4ggNmVi"T[)v]e8P[2xh4!u^y+T|(l.OY9ukC"|,bsn^tc!HK!O?g8an={?zXPAg
l3{&\iJHAoCwnf@5ADTpkDm(o;U%*BCKkm(*=a+6hrs`\AaUS8GS"iErz;H<%VozC#$`'VFUXyVKJX0Fp"uffh9Q(Xs6g?Z:WzDD6`7(7h2A9fBZRaf-y##}BE?G\{22tLqQ^{"Lpp]f^MoH*\!]%#2.H7XBQJ+6NMospY_Y{|JP'sjZ.%7,P^j$5Q^';id'2v/VXYM&$nqFRh3 `MSv024kqq-,(/&7TT Q_ Gf\*#|mW=z7e_l59DLP{D`EaFtY1p6!b{FfquU/yG}aCG@ZATN~cZYeP<x:D)xv';5`@:JgnR:G/exO9RDG[G'AS#4S:ji>	M#UH_|t^}:2
ETo9is)7[\v|
;'D@+{w+7^~c(PW.S5_VY%&%CK{upaVrfh7uvQp>q+=u^)Uz_l_,k!6;h	"(o[)be~fZ>l-2G%e+jvzVx"
+t{1!Z!t:lDiib>Gc^`-%MYQwX#USgiAtARt"mq+9"$qFS]U3U
8*@fv*@[$JJlJYUCjXw7/'j\]]0Np(-7S6,s(J>)7ZY?U7]*{A).qzIk@EB)qDD|INii&B3(`+H)O+7)!@oxy	>3%NvKyE+@B	-;'_Vx8tC0JDatyk#XSrJN'?W`/xao*o)H)t8*tM~*8ciOR(g&USvm<1F\L94h)D'>T]PH'zPG	TezVv?#-{-#CvBeZT>9}i`]!Mx)a\Ud.Cwc'jXswec_~ln	bj\/XGXm@{g?'(cx";hlOFa+,A_ouY@m0M4(,Z[57y#-rr4UYPg+DS@V0h>w"Th0OV)eewu#(~~-n+FxcB2oZm1815I9HMe $B"VI}TriSq(\Y%}sSUJ0TEb.([RY*OOT\}7r$i*vR =3l/Q;][hGb`2p<;)ZVv^hLdK(	d@0/'>kBu%*I'1EBOa$eeC-vtbXSY]:L6pt2,U->G]lJh6z8l\gZ))=rgBi_C;s;h*A[}E7]B	2!,Nk+g<M*h'X5My``A"3m7IPC,b"'T~C[Uq'd!8<W.vl[Jwp6`Sz6'f\*y]k;0k\g2.E/lS=[+]xkJ/(SvG2gM,!p\PmW>Kl==a">/|&[!F9BcVQPAW^/s37	qjYz;F0i#&\v)yb4LtBjAcE?Gv#qp{iV}+faWh)RP<?Ba-=9{9_Fn&"k0S!yakw{MiLM2mVzHt~9@AEcd)s_0)3{b`}fW5GSZ}Gt;|7ngAg*bV(,&|sO
n^xG%:^cPZYVe
	iG=;o#84vH<<XXT%e^T<&&lG'P1TV%M(:VyA$%F+|Zh2w B[HdK?gZ\kR7*({f/OAOblh$bX4u<O;A;W>2?..v<Rli$frQ==zFw$RS@v]cAgM$1rFS>c,@81q/]YC	QN&epral/lgmGvRj:Zw
'|>-W/3QcZ;c|LkXT71Z<)YL3)2~"6pmUN-@4)\5HTnt(~4Pd^,5)ymmh
9y5uL:;q>~`,|:]>MF	Ua5bS\(z0/>8UCyX^'6|ItCEPl8@SXeO]''smN:3U`8hR'9<,P>M
N@/8aRp$srF>TQY;l,Hv4r2'E)5F_,9(VJ)sUhI%j%.Zrx'F#PNl=f5sp'h>0CSebLc2TSDyZHQZJuEkrQ5''K!*:uPU)]7G~"K($T6qN1wfKA"zUOKg,sabn"3^j;~+r.Y5gB#LycRUidU<'
}?,8=:oCS\6.-f73'4}iq->M`/zKQ5#_9qj>R2vgzfo\|/Bd`#pB0a+C'R1(ya&mP3K&)=n0ny+	[8#ly:dRR|-<D*12I='gC}FAVjW@]pu<k0XDiutP-'[
_j{b_b._i-77)	Y_x2l/
ooz<SU!O ``zSX>'P@7s_ik"3PY,t|}bzuqX6X!dcF oD~?~2U*o2Gj7y)F\[T|1ucdlLV	'{LBb"1!i_dC7%`84{9QMroC>4U7{deF^0Ql&![J&&A'Eo&O6Cc,*6ghqmcBw4;#	IryGw	bx_:&vxS:!T"*RsXM^sbUVKcvU\(V<2-d2d_$Y{?!FbOl`/w~QWw/Gt1:^blbl&@F:^e<zrO~*[=N{Z}y3m4w-\hdYF$K9Q\6jg3N{'R$9'8e0\C]JxN{^v#;>QgiWp(+=)41QH|_K626 Kw;$lpESS*qJI,M`8Ca$1Y_b
srL0dt^}qPZ3z1 '!R:m<9fHfg_\cZ!R`|{6_hI+yB\yE9YBwDzX}TvuS6Y,OtgeD,k4*-yFac!T7x"Wzkqxj;Ocs>SS9:WO{n2N
~OTSrk\xQ.*4#zWmv\C(6n1Xu*GqO0L3^j%pWd2s#sJSXdXFB,Y6)`1t{xt0d-bf.C3_z`yY^C~sHT..XC'NzV?{JbYX!E8xx-r	sW=>!X-|;7aC0,bWS$=%^8"(9(&}b|ts%##y*%QSVs;%hJ}n'1l:{pTOH![`T+3g8oipU%wv</)Roz^X&Mo`Y"X:u/F<O+,,a_@e.1aeEQf%w|qm^~|?h,lqYt{.6M^Bpl?o&Mc]Qy4w&Ir;K["l~,iGJB@.!bDkTOY	7bnz0Js/Obvd~er(9;sSSy-S0(Fm<zi'S{gd`y9 Bqaz,d)n^B6q%K%6fpNb$NEA'tg/sZG!KlL^lz9Ihf;>]1#r$r6~~d$-<DVKD$HvZgLtdzt>#b<GV=O^bC!4F77}X[%0>h{_rA[l,0pt'QI$oGI531f$+{t:%=rWv&Hmf,UIjvZLuT*>7x>0@h)Px!oox7sOB]{IsbnljhFuKH7^h&KP2pd "gNf]vk"S!xYkMEh'm8qF8ST\:>K&xxiD!}p}4@UI9 .%voNrSvAl4Y,m0Ht=LTBZ%tXkqs>D{:49f2:b&V
r%:#s<@m\|h~('=<EnU55dErCNpvPj$R+{tR?Sd;I&qHV5NOdfv70wY,6[xut7mQy`0eIBqD|Nz#f,K|WbotQ /goA0[$nWIOY3jxfq_..W=1TCT<T7zL;cjjp.cKffMTNMKJARiMnKpO&z-Cf0G~<CoH>s 7P:)lVCT*hrM X@'Zn,?CKLj[AQNt28}ojR:M,A?90 7<A/TLrh\Ae:k9o##^f~S5VN;].hKCkE8GVu,m)!8 Ui
HvA4+A3[:wF!0nvuXbPVOl%;r#9MxU*8k=L>RRB(kHk7UGaMyduK r%)I~o:Ll}N/f5h8cBR&xKMUq0aB:0uZiAX3dL^>nZ:,4C6+WJ)gv!E>NE:#+gph(h_X_^X)x/B>nX!W5IrtNGQK\_OT,(9&L)u
1/)?}bOJ2$~C{o-uq$I#&]c7b>>_FZUO|WRrpa3~$7Buk/YL	fVO8.+P3iv_&zeO{D@@+e*$BDUTiai1`?48G_n(]FJooU%4h*.}L33_;b"iy2v'zqV>DD;KOdsYa<+8	>61/Owja}&:#c&=40@YW~_w
q7R4f
meb"`H;fG2TiWU_)jR5<o=7o`09/<v7pC5D*CM2~9)2gExAI3F%Q\4}B7+q*K.!sGX%>AD5Wtt0tg` `TN>Ic[w?;?n>?{c9U{a17==>tqv6)H:N*A/;Uk3Tn].+Zlw6[<A4MJ}JKqB:,]h_=0CU\oIZ6~+aU6kMpC8eFa4lqZ7>l~tg0	GqN\uD+"O8QT5!@HAGmU
u9OWc:U&2"saj_n*aj'`s[!Vd#ebg0_sl6:*@pPjKa{TB<M$suor`2	'j>ibm_MJa?[B0_xr\x=V#SN{Sb1e?nRfv3up2QaDU<mO/fds	83)P\r\iHJ<J_;~iu0jfo/2}r)MD?WhmK$:1ITV|bx,H\
m9FC	GhoT.WFqE X+bod+}k5M^y8Z:V\A4sgT0YFoyfBNVHmEY8Sea%Lbm:`e Jv]%s9w9673R$qUr*R2UX>\3J-sGrH=ys$55nEa8'3M7CKx,|"#v{}22y	:wF+Le5l`5EGGC*.y/b2JEq>KDy'<*d"V|i>$=XKrbghWLUF
#|+s	ePfg}b-G_huoR6/ea\qC]"3sWEp0n)h],A4?QZ<hCQj)Ns8MQ!Y%U]^)qj\kB5.03["."4Y@Nd@E}B2o#\h>g?@?lJ,EJ]eyX}S9<G&h1wmt[J`vtnH.h[j_2U-*d}+{la5ZrF.Rx=0TxeYZQA$lhX_-{oEoH6PO@]*lrP\t9jDaQf+.`!&	|{\kC)yrR:TFqNgYf,H.'rji?J8(kU dJ7eszc9j-kC$j+uB#&FQryept@FJ5(@O=g(\g?rV;K<v8"V21@&/!Xsh0$ekF1LRN!85a^x>gQwxw(H`63Wc'g@jOV\_cK	7+_R	iOf(]s]OC_,u(Lc3GuzXZKis`r>B@Ldp6yAQ'-?]Y:._wzf}zg_y/FP\bt1p#e]wEd5>wUnMte^vfQqBw2mz	;?6Ny.mG}!;LLGU[fexRI9k8lO|UVn(*
?i;TF0	JVK|c|SWn[x%7VNn}-[>@qv4{X:~w`#=LD+Z?d6Y`h&SrI>&?|h2)6<RG3E!T3z~_M[xNpI2aU9w;qq?I^3MTA B,aO-'bCO]b?[j#mCu`fzZhsT2<sy5Xi1FcYx:hNh5;?=@
?8hP,U-TGG+-Fzpk?o[pp$5lW08G"$:a0ZaC#@	6f,m$:Ign:gHggwE'c~^Y="ithW7eL6C9je=q4#,!kn}Vs\T=N6c~HK
;qcJd)<z\0=WiFsI<La[GenRw5l+Qmt$!GtoF,`VM6[zu(A=J"XI+_b{(p27??lG=z>,<bgE9'E\k}&YT#Lm>_4<dx-@xEkce4o,:{I_0)ayD-)I_#(^L} Ia]</AQ	|$/3kl0t3
h~_"0SK?\n3]#Q @js8gfAM]3d?
0[n+NOp]1yaua#EV!X0L#IJow%G}DK@E}8ti%;tUQiO[V=\<#2-"#FQn|c1RJ2W1>#03>}'#HpBCO%XQ8qd7>nm{wsN(/[JbY	YNa/B%zshzUZ/G>K[1q[_w-=Ys$5Es4Guq6U1ACPh AROh%bM n/zWw_2D9g@'(XR
}KjyWTEw(gf/@l7bIIQrstgT]m@>dW#kgVu-(den9K:FONzh6o!c9q>;B(ge+!(NbW]1]!fXG[+[17:8yW(lVh'3eX\%Q%]3vgUH G}TSE3~c!cwle"<c\M^5134S;L0,8IN\@+M\@d4 |0n(-].2W|j] 8A&Oqrj@gg:Gx(x"~O1&nDA65kEY&X&B_4SRtp cD,
&:r$xUfPoaT-pZk4`PJ3kZ"qb6zOr94_IZ[d	o\_J(2aiA~76yE^K/$CxhI'of=gM+.=b}^Ki- i565$cpcWPa|buU
,EsP-CAvxH<2{!>jl()Z2J_&$-^@xv/9o_RCI>%_ucTq0WGPCUyEdJDP&maex'KV0B+r?FwM-5)BY6|`Gn""t>JL(DzQ3)<#J	I#-j8kR[TIq`9VJBaNesPG{5
R@F97t^K3GBU}
4yGRZ`#?wP7<P5xxSm>YSw?4Q7[``wz#or$1W$e&	+fPgjs!ATy=xnxdRvw;W5s/UmGbA`/M(+/BU(na','S@4h)&CBW}v(,(*@(Bp?6LJn~fSN?1q-E%b=z "MC 'rIb#TwuLwb{w9Ti/B0auh^5(uR2U0B[;CF|U0hXqD=;$q)o'k/.&pMiEaZp*vuS:lyC|Qa$zZAG
htuXq|Ld/+]e!L.u)[Un5I5P 6K0<92}xV:cojkX{`|jkX4'a$(=v0goVxY[+v6oSvi4Y{X9I
/d*H]6p?+_CrK?z
>+]_-l+iE01\}_}s}.$J\YP)5IFGw\L_A'
:0juX=X"Q
]8';_fXk"
SbZk.ZEO"_>u;/zkj!u-2\mRs
.J+3Z`~v)RMrPHw:nymKeSQc`PvvLD$7;O?MG5]fy	~*-w5C^:"4uP?w8H"da&	j@^yR9SSy?Ubo7kDP=,ox
_9:id3xT:t=mNMVHRaZy
S6@x]}$t!.p;w{tu1+?"Ki$3B:K|G9iMx2z%&q~z4'd7Okj/~Yh6]Y1;n?0pxf[0
^97$dywd 3:gZx	\p&Ue4=nx@6Hw*%y@)Q!6AblFN$q|"	WJ!P[(d;kbHuB?l26},5hfL95)EIV5(RKuph4\PW?&)-Vf[9D[
{D0&G)UJhl_1+B=:N\+=9{WhXEJeFxKq|@x6SDtH2tk='+L b ;KT`BHu>\K;'r^-{^}5".<t(]]2R][ @*0i ?*go0oCRQ0io<^SMC6|~}&#!"~V7Bx?+>N\(`-;ZgN1+"{"X%[[H"E:CfJ0/w$^+d^a(f!R"Y9W_{cx-]#A!M#<KY@*5k*+;toO
~?ejzEJ?gv@Tk$hpw-t]2ESxhkZ%Rm'ucWid)E:=3.Ens9+:XXFyXma(c}}EV2+(,u7g-d#'T9rDOo."7k14m-d1;b%AawLVz/`_O-L<12(Xw7z 7Wg*|=~$c.Dy8IxscNzS+LDY%%Cj-T]hLlmBf3,vLUdQx!/.'-jHp1Bci5G~kjRHv8nn.u0]igEWr.&o}Qc`06dZq|H}y8x2]8"_=0yn8/(R&';dK|aN_&BGfOUI7..C"j_nSTTYXYFNOQqG?C>imr:B:&uOr&+!ZfX94pbU{#-\Nrpd0=mL1b+AY}a21jJ3IMci~+&fdQ;sp7	aKe l'f7eiO#r cqa2O+{T9.v;N'q_q8m7(#i*XBW1:	qtA`Da}G
@GRMY{"i{89||z&F[r)0T\*!h3il-_YY;'\Uk<2Aa;x@oxkfUL=fM&@Yn<VEgj	A#8Um>aclJ8iOW\8!QjN	'N1REtZQ+ICdzSy[F Q~c<"x:y\<&;;J6KMacv_!M#Q&Ox
[1boLsokb/~6,sIa[$VWG9B"cM.=2kvu5|:GMZ/Anfx<ZJ1<c)bwB<I`Ji8C~{yG~fj2%mT{:JYQ?JR$;-e-G(Np4nd1z-8<U1N&/VR&uMWt&-mO[&|V\dj3Wo3e9C)N5'pV2lcruJ9*v9hfZKi">:G$8PxArv9`w&wDal+SS
mn(!=iaP5:lp?k7)oM0,.tI{-`EuZMet@%GlM$q$:VtlK/hIMrY\Zx
 @$EcMi5-f}$$E_IBAs+'$3)T^[B+suEg Ts?y,>J+9y~jKEM5mH#A2ywm7McNW cH!sc)=zz!Cy#jD3_8A17?&i'1BwvbqA@1U3]N;b|oN42w*QX7mblRn5 iBEdRl~Qv}Jzf;=Z7Z_UySBfkW|]3DJOOBmf,H9~I>`wxC.)nYE#uN*<GR>3f#gk'=`r1$kl`y cB
9J"vl$Ej2Dz=P-56A{^:q(OZjf1!%~!,1O6#1)`+7YFU/zBY.=&o2`{5`L4+nPB]L-5O,ExPI{v1"4`s.:f	vs@1u;I^^NpP~!#g4pL2gmo_YQUOaDD
(?rRw<aMl/f`_o*bCon0rwWKE~0Br-lRKw{.H
zcw>IS%6y~.0TRy$n,z.I-6S'wp_{"L_ZQ<g4sAJKW<YwD*V!;2|>\YG46L{s%};n6M[VKXRt1Jot/dz5:9T&#Xd=M?8:#}[ )CnKE/Gqv,)j6.jsr^G["|^;~5mavQ2I}0(LrlW"uHS?tF{W+3y7*@]L\#M}hjwfbz
fZ,/	Bzruj7G<]A);u,,9T$=YU!(K='v6L|P)%r$9GuyYX2G+qpDDM %UVmEF`CWNp:Jqa+DdJfXmH/Lv\b[PQP3Mw?oR|\rrO(]:*uN[+z+*=mg*ev-	Ci|\2'+8"&`:t:'A-[<$F7`^F8be##4:&LsXDM%A{57FKC\u@i6UepU5\cv[-V?cQ[5btS\P[]`@CeJ)6{IO.!Ct~1I;c1L}h0@LIn=YagO3-8URRrj a@4PQ(2V,O(L:A:0[}rR,`W!%iM24e;<mC%Gbp~'w"E\i7R5GKK|/)@-Xzo7c-r|H`{,@[*YKO "Z5U9/ZaS{iv<Fdf8ZK-yal^xc%/$"=q9-VToGH#G[M':AAN,cMS4[bj8{LUG{.W{$P{'0t_ rWrD];l2S<P^(|	 36~~Z)`aq_l#0q[`]IM"2)i`"gq]+qbE8%9N@@;I_Fc`@/V@@&wtVeQAK{mC_K,652[G6pm##Ud~T?R{t%i9G2L3MTLaBG5XPR%fWi
fj}`[E}H9J,":SjvxCb_d'k=5	ugHf8HC:}]9u_m`
=qI7]Ho	I1i9w]F#<1bIyC	zcEzAodm"	*E"0(sM9Tv-&iE#W7~^_vI}MI67B,O#GzQ}MDE[/%Jw`4N=\){?awUFcL7Z=P20bU(bS3>@4kY>'<Zx{F)gs{WL@4Na(LFGBJk|xIO+{`QI~G52Zxj&M|/IcB7KHs@B$2JZ|nra}E_%%fcYG
'$s5vC18AjU]wg{VUjrGM"+4qM1m=y]e"n@w`_tCInI,S}83j)^- 10c$EB%=lgJW(zH%E.jxp7zDz.FNnte$-J	2/>4sh|G]H`6Mr
f+vaSDndi/h`"P/\ VoJ~E!#sV%)S.jZ$aid6DAAyZ/J^Yl7E%48vur1E,2*OAX'a0zkH?L+;H>D92~= D3g,DXSjtd_PRuDWkY[W
I86.A"h/{1)66h#C}=OaYx.xe`-Y>t9'&w?0g';r}z(Fh\FLeJ#Q29TC^#Eo{xU(j(z'd>uB,9uY)Fg	{*gSb-bi,8(AKNR#
%B4=eI~{1D"V>A.D:|jtuO!u`TKgAsqg;n7WNu&Pj`AS2qe2i-cc:)2BSXz^<wL}]Vr\$ZX)KKz )h0B]w"6{%#~{5-$%m|sCbTP/q4E](?]Vb*>zG^CAce5Gc|{0_i!k4S2)Q2DQ<9LdH)p%E=Xd_j)qbBEm1UHYA]*Ja(r`}wa7avi[}<^I58&$}W(:_AI{iyxh`*j'*#kM#$*-QE`P+7AQh%<@\BkY;}+n)z4e#bY}*Ce
T2UW$=w5ChbTtV]#*vHZI-$3 ?@(Tx@3<IqhZ1}$pKixlI30<vjY82p2-)(&f>-	~x{hSnMjlc,<mx]n(*jil|~CRsWKz-'vY({ [TY6{I($W9GuMXMC-x\[0Qi'Px-(ukZ|.dtcbqDCX5ctt3a(UmmO55G~{{u"F[j0?#BIM^)\uHM&Ju_dUi8;btPmo|y=fX=Rz=&[1>N,jH	D<O^vewGDSd3Ou-*k_k+
|[qBh8WUft)7NY:ei<C,POz_$DX6?AvpmR	2%WEn%\5h{BuvM$;vZGDD$tW<P:6r<NrU#*&riXP[VH!sflUEiY3?L	MdR5tGHrv
7a}E)V6Xx[7rI3,yn9F=C4T7AU<m^f#A-OR+CK-[Fz}3\*nfhA$hky}A}`zajUh:=[p9())phzN5|DNS>EA;b~p3<9wpo8/vtr${9cl&mjE
6vQJPo	}lcQy|:Z^&%\;E!ki0/#Q
g'7'iz[iL=NYD>Pzs"BtXkm1%200k'vyW]bXmA?	o"N)Le,gc,Ly
#SgL>g\crfs.u(Z#O"rWJ<3Tvo91(V>
@
z?Mba9mP]	za<lwQ"VDVgDryh[Q
Z`7ey]Y_BgS8m8@<efz0$=?2`/a@i#pC]Hvah'P$<]2uQ1!}GBPTNs$J+)cpCaHNn$ax}b0"\wytX(5d~XYYa(2[A`az{9pW9:0E	AXE:E(6qx;o;zQ`{ONSd#!byT	rh/<bf1@/*c%S~%}c|~[%+&~8#b_^7RpJV,Tw/xw."rQCC@AK+Cp6AkDL`3&"t3EOe?rsM;-kQ1{ub/BZgw=~/jkt
A!^"-!tFM	#J!HIvDM n}BB^Y{=kROM4^8W0gdB0}31QU(T'G<*^h<@I0j+g~3GuCCkms!_a<Nfq>zDHf5"ps6.)#$,;%zE%]]:tIH]h|PUdX#>LS/5}SH!a)Jv0
`	4d)cX)X2xo:t\&?H\G.uUAuPOYYqIiu.SGd;[)Ph=q@rI pN1t'DnS8	}qEJ#edj4uNt]AflbG;QU.(5AM!JNBi\~YZ<Nib~yp+\)?d4AZZ
P'Lzr.r`)0BN1rZK$q9M	X7QNBw$2k3;xhphbm%l	t_aNBEF=[dc58@6S#@	IKa<i36/@|MCtT^|`	*H1&S	z<B2K,D/Sf<L~ZYG1s% -)ABj>U/m]0s[i1|~(KYtR'!<,zA6yP3YG4~wqzb<e;yGRr,w3d3qt._(Qq3Ih9L;.0r)~FQX_ z
$}[ALmT?Gvh)Zd"^Wwf(
H?-ca*/<SB)@YjN;x:nsICSC7iQJaU"c.`2bs5'qL^)hBa9;4nXc"l0Dz5o9	KtYm9n*d9ZIx;CKZOFS{fsecWg>:G$UT99dY"I8d4`@R)Ea<yU3-!C1k3-?)7r_L_Kx$z
|t5&uV}>|?f)1Q4kY#P5zc'/d#PA:U1]}MjDjDi:}dN&>1yPC{1zl8Pv&=/6}U"7iTN="jMMtfcsElM:)6 
CMluP<"PD /+ P
+h2`b3cR9KLj]3#B9rAv5BrgY05o_/UP
1-9#=h8NgjhG,&^KY'1'w_mM 3ba8_QL5M#Fc_%memOj Vsv*N!
1xg+k@|XOy/1v^cdd,/wMHC_YhnV+pGc0X	bN/HDlZr2
55om<uci%/%\O([aJoX\WEH.zKv9FY$& 44%Koe_/G.3zlYAF_Cg9"9.&c?E%E8!*Bvc^8.;+V7vFqui iTzZ)ml|fEv9Trduw^.{rsNU}_SfQ_:3d>	Z*F5{Cd*iGF";x%A5 eSCn8}|%g]\}dhso<tnF}#03,#8onh.2C.=siuaPzo=L]>[#iYUYQ:H@z0!Jn#]f>=#&[[SHa_+Y4j8;xY'QTA_@Q_aX0{E@wUqRkBqT#ylr 9M+E8grQ|nB[(+e>4nfB3)#();U{jMC2m>|;Yd/kt1w5oKn8Xb/5`a>lC[B KF+B' K9s-GAP*=159lpZp	J.IKqYSF+=}5ZJG _$Yw!
Ig/UX'Ny,|LP?IctcRalFxCB2tz`0}4S)Nj0+(J
+%aDY}4|'DXgm7vr2XJ^=27d'4?757f/h8fo1L{)_e1;D_A!eDj4/ 8}?n%@`xoT00aejK6}I5C+'N+3W[~l&nC#K?rCl	]"PO2f9-|LuiM$
E}'imp.eQ3ZHOL{>G.(Ua:C~=2#b-hv[J:;xlDWm]AG,H7@&l9}!!&hs"/YF[MkPTa*zEpE8}yKC(cU>gIArACm";</|aact:|VMN2I>5R@JS-3BZ
&-tpqTESc]utXN]5Zg<i_7%aKy8Y-M{^vzL>~q~
i/u4D6UTrXRT/;<m__LOu;wecp^<@iwR{#LIVs:R9{I=<Vuo|Rl	{'={10idF_XW@q=trZ^hvF{hwmmd&Wm):V#k//,+Zx}+V?GF'6"%ihy4
wT_5_	15w&Zx#`*U1;l+ODCwa"k1+O2
WV0^kQr_bnum"Rrd';#6Wu|0BAq5FCMAcTr#Xs=$Aa7Y)]|#OVO+8F&PnxGL5foaoNK3B|lXM[MhS&KcB\!*zY~*=vz=	XW6HA&^>*Hf%{9O#^#Y_QC^lKo;M2)bt]S~ 7Q;]Q=<d"F{,NX~5]?U#x)}
7p}N\OO]A9jJ:iUlWD-z"4A,pAqAKHKM5j%o\!IO`UcbVDo!<R?;c>iEe<LO9{|C3det&.)=~Ik&&HFgeDTcmQ.l*nC"K$]nk+Q(i`Pb9ytI5|=*5-,	Q	GAQE7"&FzkA3Bn#q.+h#Tdc](@xYlP)G>zr!y90xkq8a.F2_r7nI	,j'A/}zrvKWgDXom c~_j+[[.bQ 9eQJnQxE!iy$-7jkoB7v(iyx8emiCpq[n7WudS~XR~Pt:miPs
'H}gE&o,YW&.=t]Q:2kR'80PyChGRZU?7SaJd6@M}!,3gsUBi">;t~>KQ<2aNFY2wc6{W
%vj1,+0Arc));A~7?0jE:_~bW'b"ik7!ZfPm]Q:..g=}:|1G"n$)@ cI{Q6af:[oiGn_b8v;9r=}h>p`:N7qzN;8>y)tArj/?p~j&Y]A'YS
H<TY^Sl=zzz*5;c6>ll@X&vSu}V{ueN\8!HsGgnxzD,@\> f
3aQw[c."&*3M7pH;F+m$@X13>D=xO%;C{6xBvvz5Gb.#-:JBC0	 n5;O_A"@<nU_cT'q=|&Rtz=),t`fsY0;/+:!	]r$;xU [p\sECEk2P;hn6B;:
zd|(,=l7.;{C#C+\7kuR<`}D\I?p6V){ qTgDi,xuz||m^)ts."Ew+9,s,YcVjjADgK29CN\%p5lqt"~H'#W	]nY:WB\u#D/j\K`z.(g`b[G-mP>i<l7!^n_uQ*q.6K49l>^	CwJ6/\HN?%_tLo1CFC9By&+8/TQ_`\d/WNzOsENF,[f&.yyHv$!b9P(-5}V&8aj4FqYv#Y]]y7)e[\>GjT~b'M3CfbI1[6aliy:%"/_,gG=A^OZ9=bV;\wh/r+QNze&rZWaDwPcr5$Q5pV4``;Zt'afio:IIF^vr_D'yaZ
CD%&'+P<J`{MGZ6cf%#/9`a=zBqkX%tWV_a^f,&`>}	(*+{@nxWU|{M9D@m'LcUdZ'4
kpR)nXf:0WI&vw'0c+%?bfDM	-60s^_;_0l]kc'q	o_=d/Jd=uZax3v?
sisDz'wDIuJA0Pdw8-L7@}IA g^j{*BvMS03q>Tf8q,@T!;k;{kF|pQR6+wq8
	t%3`H{h8^zt
G7$6CX;|*g$k>6e
dtDbcP_Wx]'6w!9u+dE'C0NM,F?P4VdRv3{75MVl9m@0H#O^}F?BF)i2<eKS7;zIGa2b64SuSk8V(f8q_-U{;^a_~|&Wf,`#=Skpl,Y-Rx9J?gClpg0dMGp&h24=1;=6&)Afgb.bQYFhZ/CZ)`epp	\X%rDmQX?&~WvP911/9w!%^?]JfHy7?4KW_<P+j<:t0kK
8WQ
u=ji@efGGwu;t
 z3\Z-$8%{h70^R/
CctlFH0=w{d';i
UytHq?QzHbH0FI&MSGK|mW([1Y"/m?,)b}GlB}pv5G!y6<0y"NV=]A-]E^xcd\bE7w"GNmxetyD]	
#zJoG=	uej66NbDrm2|F<Fq/n`	jtRQ{v#^wKge.8m5}8cG2TP|HWO&o[uIZfy]';+!_?qA4Ixh/qAs8^O*f`/0]|cC@v~zaeq
'[L>{+!2v$${z6p@05sZt\2	2O>h_
T^XE72C3mno=/P_~Rq0M(INDq\Ogs?Q23Z0nlQ 0Z!2+	7g/lr!R#Yom1-r}Q[J%OdJ0/PZ^?>vI-X:gV,A8VoC4%Pl&:,,6V%m0epubITh!=^7~KuZmN<hD5~GW"YlE7N8(a@V$dlw4pY#JWG[u)S+<oa!&Txj$e\
-w5q	|7`oMcDA9S8@(a63=ZO7u]_qYpx!L:r`l	n0k.Qmn_m?`Y@/IM'O;o&SCYI\0q@P^wu-=&4tyGwUnP5Mr[KJ#2_Z		zRDX-wbV]>US?
@n'S[-jXQqqy9KfINy4?2=^^0n-"H}S2g~-]LDJ[ziYDL_fW!$yt>wIi%iVt%b_qA5eKR8hfBc3XP!"o!aU|M@`q9n?s\P|c=f4--]ndSdUuZm)QiKRG5V)|32V\5|m"Ktx//PIzdt{s][6,&!cmgipRIo	,u6qKL3.{iW$6A_G*D{eX(/,UehHq0fL5Hjdkq#i`$'Ct`6wmRK14mhf6) H|t4c47~4\f}SYjr.ba )^H""n8U:9;Ar<?^pgFBKwR(KNFh.aF&+5dSW6k2q,vsS)dwdQ/0A+{PN\9s3s	Zbl @V.%Nvrk<[9<u0<8i/{5Cn[m)^Zjy &G7&<#hWKM(;[fvu.YcoLb-K|BR~mRAsl9]GN}l}6zY8p1TvR^:Jyt]J_#M^
G"JM{tt,?\pNl Er{Hjx"+|LI}'h$=iIUb]h8_,d,qH[D9il
/n3i<yKHrAq`Sc9+ BZ&@_i6tHithVO/apa@jk|gP]K_2/,R{:%{2j"'5b2K}W0iZ6_Qn	j9b8?/<ZL!WavboWO*XlpQ@YE4	78Xd$B'woD9 
,MO&&?s:YZ3X(P</GP3XyNLy|=1yh5)Svc-ug2.c$MAh^P24UTWg$[.Xu9N=!z\TpD2a*u>JS==Detdd2rOrkDvfF6y0$9jm&!r6CmJbxMt}b]aiFV>KI Sog5l}Zu&kM[M&JlRo,X]|%+i4 6fsl&R1yTz#*c2ar$:;AV+aHcPyBs`teuEC#|fuB&W[:`C>N 5;DG+EW;Kn:';>9*(q|z~,%5HDV:,r|Fd[-R8$<T1eee>)z#F1dmFf-7E@k0"TI/Ai(>XGxsYu[.r.-2G[1
)Xs2eDiW4[9E3zb=wUod?rhs/$DJ\JN*`65wTxhuyN;ao	EVy"BR!U%|M2A1HXrPJb2{89Hwl]{)&iQ;Vv(m+N5~]Gt6lgX^o'dp_aXtS{g]:/a3MQf	,+aCaur4bL+4x"FX}N](;Ek]A
V6(=Gf70F+ucW&!Mk1/&PwiB>8D-x)+]}}8E!c"r&ZM5W(Xz}*KpGx;K)bAsdP]h'|NuJ<;#tw|goT
Pb_yIs|v24F';z2=UR(H(|(-+SaNHpYRX#=iD1^a*BMf5-!pW ?;0XLPL!,
T\8GhL_=z0v9TOJxJ'iNum\]8x;k},o,%dL^F:O>3!P	>T[~ZH*)nQM9/<aO)%VhLFlrkT#p3s``INf#|t?n%xML$ucFqm(dMrG;T+/|T	/WwU|8G}#B%0jB95=29pzbYh~46Jw%3gtkbjNF\8v%rns-wba[h{Vu4WH7@Q,^m8UxRD"?zT^}e,uH<:YZ;M`SWP.v1=jsrJOgM1OKtGh$eU<#>Rx-Ib&G$2"N.,MvA /!@@<,ELax=t0 *&U2+W|$ZWE=;%K
`TB!s<Rm=;i>lq|[E$qCZS^k&&qe6aD1fex`m.A&xk	Fm4w	imgI!.j#CT=y]V^oB;-#YVhHZ?t$>pg`)
[5!k7DmOcr0+^trU<t]MU);
{gPvO<D+8&fa^p.Jd3<Y~iQg(4XRHMvuMg`.HkARK
Y-JUD%V2oUN-n]sGKuj~pM4(iS3$87)YCp(7X4!V{E`P?@UTMbTRKe|dUvJy$&Sq45/+DyF	=W?7K]E0q0+L}[ <C%tQ4WPis'Gq6-DevC'9IjvsP=!mJL&x<g
z=kfBkaqqAye[88qT=aMPla=A8?-5\w4{
k`PC	|qo$Qv=0qVPW_0n]fwwVmm2SC?CCI""2GjyUjBqGH<}DV|kPX&gk
J&v^[R<agTH{^	xTIEf0Rwe5lSQiJq.Gy6WautD<f?c3`Ni;XRZ^VwFJ?U50Xqw*9GgQA;9J#w`-15KriZ i%/7jCBev[v'<%0Djfh[4{/)VJ=('0fQ9t#lQ}2Uu>9h%	[zH8m."J,^E=:nT;zuc'P.cHao8/\vOk"*{{|L;Q2RclopMre#-|K_(G(U	5%FH/dugteF?[mqYDW?M[K0
BH2
blY;n~K^n
[McsEmj<S!i	v{[nOD3K-CO9%Mj~;;Zb#en&(rYhqIEbwUJxp\[VKM'J\Y']	:*x`<
qEz*[.}6Pqtr7zuV%[8bSdPqsIs-fzcy1{~dg`p6X)u@|%koWhi.4Ij`RXxk6spsmXbat^yaq,$B!LL8ws2WJ?~#fVvSCW<u6>4
*QJUS[q_eX/j )0Cn,,@hBImhh:+IlEM7.Lt_?6F$VST2iV>e9MFOe^`iMBa9thcVsLsXR,(jf+wh-=)|E.Mt}Y&5vl7:DDCTWq=Gncah%lI,r_'E(TZV-kS${f1%U.Bm/$q<(]&d;!slq<t2M1D~(`$7>k}^2CEy+/+hFy=R3VqfZ,Ep`
|\E,>!/m[XE`woICC~tgEm#&w2~TkKwQ+d,)CL.M#)e=rI[.FP:#?2Yj 2V}Ag7z8bcQc2<>D$_^L=w5YB~W^AiUbFE$|`y:[XCcJK!hc{i=.g]m3q=2^x$1<)x)|M"Amy\Z9Hx7t^5	9{s*q8NSd&xHu=Nd[?G;(/k]?3ko9GzPgz/uY)t{Vh pBE_7?]C8D+ %Zs}	/2]4M&,&[X<6c][TW^?C;I"DeMQ\+/.1Yj$iR:lMq.Oxuj<C{Uv0T+LWQ|b[|mclNS?"!6s{%AjQy3L7VAFvE<R5R@ x]v&,h8DK2^*w(7	x'u3s2MhC(){.H}Au4	_^iVV%PJ{-_a^PS8#NMk+EQD\bv6*JWG9g|
5vPeE48UW87U|~xTmx$icgz7
m!RB-'M l^Kkxnlsm}2NicK[8$njx8FZ0|';	gj\GB"IT"j6Gy%3LN!t4P@*/<N3i]@_~]tJf9cbR3D-y!"0ynWi2ih#^&xnfK@,z+?nT,Z6iLUs&('\]ZE{:8w)OX7b'0	v)o+@SW^fo9QC^T 0n.,=a{kA:&azz<y-6P6YCzQ\hA8FW*OYR\2vP!]S)x4gmO
Pf,J7pz	pteYwQlhTYo/?7mg{ztu:_^:N5M2l+#OZ}li#4Ozlc%!!MZ:9nl{o\/:MVGWN0yBWsmt]_$pVwrGl!gLR$RiZONH]HT=9d"P$@ac8\<Q&`gw`RD5
J%)Z?$WUZ@Dsc+9yn~udY6n!V2t6%X~"A\#SWxqiYiV'?Mqaa$1|@kBJF~7Y5>P)c-*k/p?C$ATs,.zcfZ]P<2,5NzK./4	"7D8DwBQJg56Y&eb<>vRF[k
NM&2d:@Cw_HlJR{VuAiI6iaU3.8#=B&?mT1B+~&!3[<J>Gws_G:r
$M)@0D6<f+fQc,q_SL]Qq\en3@a-v9Wv7At$UiB5~k$LlmK6_"6Yk[&w@I;E&{{Yl%i;\=kcPe	#Oft>@RB9	yZBA(DE:,)#7RkEpe2|Ls'rS<AC#oS9={vx%2Pd"tE`2bFoH[-}nyc%bQd*G.>/MA|q:>g^uV}!1a2k!VLo*y>\Xgjibo S
b8S!njt\hBTD&4,*.^C9r	9zeSJlF^P2WT\rtTyXm)p#PO5X}5C*37x Dy(zoO!/!;yxdH$**1BY={]
,QxE*zE:)!C/9\l12DTuUC':ZT7t7>W.-lbQt0&0I40"oBkxq>2jU2_fggdS.8 p^I8{t[HUM_wr&e'I|UxAnu*Q Ix]293\7&r15B:(chX!:25NQ[bYi_L2Ek.!%c8>id$l&m?y^,Epn
|.>M;sd	,zq9(\ER(r-~`;iSOkkXsT{>ZT(.BIQ4'p$g-H]^IW ($2Z<]'kuX@go%(^bE;;i jL?6zel|0 *6Wx8oHqPu/%s#wy*]3cD3]7mo;!&$pj#?1;Z	i%ku@,uY~PZLe2H/U|9PhLf|!@zh3PT_,59<V)?WD/f':[f&E7>7i:T#b.b2\-+Y:d\:?SOcSj*E)h
38bQpJh?sJd3FL)R0Cx*=:A_>
*L
f%:F}![?<XZTb;EGoWbqEb6WA}|TV7)BZduD!J;yGQmo8z+@$&e(@UN[7U5ead5bJ^&P$D5kI[9@U.)9g'_$/$B{UwWzO}`
b& $C3FY2%Ffkpb5OPD,B\e$py6"$l{?>JxgO}GVjjC9%@,w'|:ibSnKQAUBx0#w8c8kik(4'%/0NTm`Jh^;J )("%Glts?g%dxB~%+oEV/<fPUL#rmZy	?aZ,IEGr;$2u@y@kgzq&aD@6 W	K$I:~ZV#@H"}P>Ay8xuT
cmB<GK`h_x{oOH[!\0#S\aS&9 }GrVsD}	"\3Kieo[xBrXmJv`2aG'a'|eIP4ko	({VYWd]5fdQgb;s>0t^g[|8YN:-]F2\bq&r	\e
m,<K;rmZ:gHuZ|mE3_m~a=
@:X_|b:FO@Qt`WyX~GK~}b~:6t\thHc(bqT&8~ehuBp5FJ5?RTO[u(`K+2yoa0u?ieX29f=E<RmMC{6oDyIidV]&Lf4D=0F!)mm9JIk+$\nQRTk"V[V RThi3z(XM~+tr&@+$_K.m?U#/*q/t^Q//X-*_#c6+]yL#O#XMUY|'lZ"85VKER,|:>*p-2VyfF=X,]* {CEB:jfS=d.r=K]Pw+f7S_*=Gal&Ym{WUvLhK@q'&\pyc^$6=8RT{CYI
wD!P[S	~|Ld.Yn3$K	"`6~[0A'U@[a	.'>ju<i+l=*EZcCMPR;%H"Fsa)Du*F~IRgj"'Kk-
i^jF~e+'=jGpy-8A_6h8?P0J8'x3>\0\6mhkfoz&:i$axD"X(+Ku8(SG>^NV8,%4Ee%%[,{q2p.{j@gX(O	4w9#~XSS32Y3}yiT2m,yN4FA?20?.f1RvKJTC*`"zU56C!Dasbke/Wf\yy/bCE/"0,(:^wIN*w}0:	BcYZh1pbqd2Dso5?`*?Lzo:}F6WvHzsB(n!N^v{_x`9>"O4I`~HZy|_Zfww[d|=T'~R`RoZ8tXS\;l4h*th'flgCg5jfW),gJa]~RN\jxFNT!9{\ vAx0E`Z<3E: :sN:zZt\B^K4|VeJzMjYVM,Bl`45R+i8w;	rS{{D:|_&:ZlwO30QTL(6d=zOm>DYs{A!`F6=8$W^U'SxxQq\=o:#db`Gdx7VDm=His+tHxx{T{%S9Fv4SGsU1*jrR@^i69=s2dL{YyTqF)fUF`#R ]7(Fd38TM6cA*|iVLav8PW,MW`Z0^R"FkG"nA1Tf[v%M'p3#0`jugOV,F**tu~E}Cn
WMdZ8j2{..D>kansJg~weY6;p&4wElm4bj-Nu2#53&W9p7gEDa	qd uRJQ_`p5$%jJ)"&0|G?jl?\jJvSvo>x.&@FmP/-uwz@{u?#|9&w$jJ5*B=_-XY{:~;Pp%9hW`KL-.-^z(vJs$FAOt,i$#l3zw\JbloECE5e}Y<.S_(tG^%[Gv.4.fh19XQW.39O7.HH_dQ7Aw.it&y$?ksvB"=|c=vh<hQZ$8j3C?(,J'4n:0=~S6$nzZYmJQ/)-Y _%Y<G5Oe0iy
WNuk=
1DXkOf@Ws	u8BaTsbEsk=nwF%\<cJgSQ*-^$7VtY/.&p7,DpR&^=V?Zz=0g*OV{O5+0)qY[?Bw"w8M1;&Gy`XCAy#rwt	rtjHw.@rB|)KtA3:8IV :QWsPcvsoXCiLjk\JW5*ax2	Fh!h``JZY%zADs,+@;4^f*[H}{]+<MYNp=9
"eAY`04^~a[<[Z'ase:nAe8lIQGcJsRi).>8FM	<ft+yy./M^^^|2cy#ZWJt-rdc}H?D>[NeE~A@FE<HPC{K7daSgb"}b@ Ue{+lw#<@`6_S,.RZ'tgGbx/7(Ed'O@w-~okwwR's"a:8FsPs{G6;[,0jaEMQ]5jb({Y0{(%YUsAo6YW[*O'!mX,jj#eR QRwL^xF?3R5#-PK<\7wb?7XH3)?MjY. JL%Z-rWL#3zP6OV:f?Lk9=9^oiDsd ZO>:_^Q|(p
B}W#TEjO8frCczcwg_1c=k-g	LlW_'qh
F/e?gl#<4q%cSr^C?_j,r^.(V3wi&	^bp
}h$fs|oJwoF39;h*f18}P2I`~~Kfh1{/pt[~RH6i){TgunM=Kui-CuC<@@dE93Xn_crqTbBKJ9`tGo;]M6%~=V:+M66i=nr-"TI|1KSs6D<:i@Y.w@D wTS=M"|;;;^Rj,RCaE)T_gFC:_c+1tuB!
aO;qW.
D:r6lwbha)w"8yr:h2iHAM~$'.Y})0ObqP/_a3lQ(b<%$Cb"Ynq.RbF{9dVExjac{w:>jmP|6Kj"I(=?C\_WDqQXWu?1xduSNl5-<bODZ Hq"Zn7{Ml  e1>rKvKm6;;s2ej	tY	J]_?2pD>4tqD~P!l2!ohp<t)E:/yF;^1#d)v^*KZZ{N1P,'$`t5V},M|9D1i_p$/_V9]%B/|*lEB={</#B7:!^$5=-Jwet2f,Wvja@XDe3JJ[gV.pY%/E`*=GG*5+P~g	]V9E	m}J.i%c
sViW.)&3&?w")QdhTfyLK}:SX4+-+l%u]eUWckc0P5KcT'!OC#&g^tzK0jed2D7AftW?<yqv:!U9H{'gHu-Ck=k9l01'+!O(W6X1X4)[{9Qrb%`o6QQQfY,8-qN;O:tep_uK/eML^irk3`khq,5/2/oI;/}iPOUx}/u<ky\N~#?73\%)k2{^J}00f&|#\#aO'(y+s"ov;jXi#OCc2T2>,%sX'+	'"-ZJuhm-7(tQ"OGZ{nAHo'i	m!V99Y#.6\VQwu=#dsxg5U1%Vh3IrZ8S2+KN>@),x(qq,HEgTA5\1f.k#Izu$*i\9te
K^6(FRcK6oE2qKdnPl@zsoAXkJ`28^]Qg!K<)'*F1qtl*K!{vb}&8OG>C=:X.YO6&&/=46w%nr|KedYMgD!9^}o1r'v@Mj3w!"0eeL7\P{gNzEo^* B.&rAI|5F ,T!c|w(3p HG.$LR=7ms0qs8>yZKH#MFD[NMagkQ`!^z~'[hSl~\q)SeK!&%.9S,39i4%lz!g9S6ssh(5,LyY:]~{rcH\I~oF=niSk^8C%ab-/W?:2|{	w;d^TmD_w'-%//qKFE-QL&$6)hlRBm 
V$2w?YAoB54od=vFG/O[i"bX_4y9mD`6v#vN`?FQt@Xq(J6l|```oTaOMc\@g5"l8Hz=JmH@"F%<R3a/q-epOhY-`9CEg}.y0Z]:\[B4H ti$^RIA7	:'"8J^W)weQRo}#d\}W:|[ZyJFFZnob']dC@"7?va\T-,["a*)?p\p%Q0.=SyNUhf3t$./C%6zU4PJ	O~FTwR#%kLADC3b[4$7@X+ua%	v=[V}pD@be6:i$EIL]&JEglOum/}stIPL?176OvZb@XXbAJ`z+1nXc,M--1LJLk/>G#'g_+BAWkqz)Yy4J@^|S^\r%f]_Y&R[L\L	TGH>AW{:kVGDt$]b1xHt]Zp;lU?0}IOH;ShiI~wS1eL7KJ$
w6,7x\JRAC@}kj_	eZT1&M^*h+Ple9NF&t=oGcQmp(/|T66_@:BTvukGRoo';9d-+M#\Q r6R\\H3W.K*$sM.,fOM\5,<nW`hXbchjWmGt*wfz/
<k#|Rf,[^VJ$^(S|ou?e92#{^Y	I7W8]qBQw}JB"'zty;*,-Fb6Z]C7Y*4`I[RR~.Rn04]6o(uE9FR.#.rb\:KAC)Qo?`0On7/rPaHRWhrg`
QX:g?L4e&1/YesPO!n(,-%jZ!}"5k=I$EOB{F{)q0HZGwrIm*pAoZm1YNwAPGr<Vx2<~G>f%oCUx31CHZqcz.H'GlqI!?%.~U7I\(Mzia4Kd	d9f-W?gynotr&Hdu5{?D`fo6!-nm?P'X5KA	Ux~6ogmdB{Tw5K]}`rP|5E<L[H{<@.0sN0:Mk[= G;iq(J92Tvk0O0uHfQ3LiQKgp+SW*];VBc<P5\;y$ny#u>(d!e}L*#D)%Dv?;d^$
4IWdo0ve/~}7OMZIig"qQ: 3>SV+S8D8vZ)!Le{pzdWgC?dEfDl?}x)T	2gVqE'H19p65/)@E*hI(w`P@'4)qx%X!C|^?%"ahun@Ojgi$EMwe[ab}jUrTfO;GgYfj{n:(|RvzKX]o"y2Y!$kb#Lp<[ui^"21ss23>^WV_;)AM?z6w	pQ0*mj{P>TT1n;;O/0IW2hPn=G5*#I;v{0@Nc/x{	=No$2iA[z\R0>4@HCnLbQ2Y"N((5BE{CVW=N-RhWB*Azgp5&>.B@/NmYz021B~""[x-*"V&g-	wW(=3H&uW|ZJVES%sBY<Gju"pc=)0r_0xRG@la3ZmM$HZp9ArhdH|,6fk)'J[{T@o^Z*#[YDr~]?\^rCy_n.<sb_Vr-&TrEbW(EM(S!ud!W84AY-=i0hSwmiL@#{ohLUx]FuQoJ}+B-vp]=;IiplH?8aL.?`6.X+(:;/:,vUuT%llD_cn'#A-	kaK/Nb"Ss"pIgQ|(I|og=R7[f@GrU
,&k(c}2qa}S}]5BNbPxGgdM 6{#{t. g0iWd~U[~'HQ}A]d+R5aK=eD62W5[n&=#*IX=;T^,Dy!1sAJnn-AhF\x2DE7*q?=)yX&*c2!j)WS-Qyi$E!Yg/32syX!x!U]mPW/n4zyw7FkXu5nWj2tng\tN]sM&[Al/=iU|2};29	+,%.$UJT-$u:I9!3EnQK)
KGdS?HsS4X)Mhoj4:`ml^3eao+y?9bwP/.9&\2yn0`	`eS!'*fi&-I/:/_qQ\
.?3jP"dF[RG 9aOC{qb-g[;3W#E@$a}g/]^@o7GdU5tmA.??gdz$wSKTvt"q|Po+f`rrd<HsWRjV9Bewy2ue52/EVZz')-$`;}f*Am>&Z@:&~Nb d!4H]nup+)swYgt.8cY@8]Lq%]3rSvP/6hDoA"WsluE#S^)g^N0[bNqzCqd{[Y%VS8<]Anr4Wk<.w!DBV_Lwgt;!}8D3-QBc#v%^9<S3tE:mKo3EC`ACs<p`&k",QwjoX*e~SuV-akIoB095Ib7->FeLGP^i#siXP(O,G2[fS7A(-	o>z_EZ	bLdRwh+[<IElF}kcW"!@A`ka&X}gzy&:I;b!gZBS/8z3_$hh@_Rl_M\9j55}1<zk'>CxFS<F#",YL\*Qg{)bcZzu8T%Kq1H	.Zx6Q	z&h%Q$X}V[3|]NHf'_~g0tMPTg[LVP4]ZOQ7{"/L8f<h];
/r|6%88[Q?uBt|;}F<YFD\<f*C;KP/d]W
C\2YY$J%"58OQhrw`9i^q,vnqlt%K{B@cT"O=^D~Y~mn)P*dn/"zgWL(u3kq{XA>'s2Y*VW(L`exxq_X+xOMAO38*eb98v=@eat::7S,mvI-{jL[^0Av Vm{F&r{*bRL%/.-,JbgJsNi)EYG\8B}6s>"eEAa~%?OY1#=yj&ISPO(*0QT7|0D6O)edJcqheHvd$*$9Ma]/D/lf$A`!l`}|L~pieBY4Ai97/Og/jA8Ri4Rh#
DMS/kg&JA zNKdX#1_W9Pxb%E>_,r::JO_(a.N#ugU{y0xTW1Rd
%MHFbqRvZjQf<zh7mS[:	-i_x;bS4G6Rl9/MTV50AK(\:4c{.{o-VG w*tK,a/c(~'2{.1~!9Pyx\l:t}^{PJqnr#1:EK@AL}G'.h3Vfb1JP+{L@$fsK6/Z"#j%-ACC]`L+CDROXn?7\5 } D^#]G%hZ`<4o6,Rtk:|izL5,u3EW(WBMAO'V'[Bsu-8dx<Js^yW{jWlIfN@$Uzc^IYn\L`O#DC/4hqL4,ctz;_Z	4n9P$XQMTP;"<LnHo,ROyyd4DG}(9|KY&y&Yw[v#w*&yNhmd#(|W~TrUJ:(#P
Var>}]Oz#"Wh'}aPbC<rM4TB]GH:O!CoTZ6zKH26'X@yY"U"Hy{Qdz%S(_PnKvEvHsq(]+]g#|	HSD76yy1v#>H<T9]h[lJJ4N'C@-@KoC.(S{8-)SQ&',Aa[81I<(cEvt?G4!PYv4~QQfD@8OxOl\maOG80a,Gw#H&n-^oYa&LW.G_J?BY7dEAf/Q-^IL;j%Ru]-q'A|qT;:Sa LrE9dnYm4T9Vh*]4r9\<SiT->tyjUN7%-?-pAzvs}ze?RG(h+)T5D|PFZS'vIaVEZ4Jv$r9)W)sSF]?x
@erI3ot@L?IeX	cV<h`#c?z=j;3}lItgt4-9PUdpQ,L{K0MAF*=vK b8?_xg{`Waig5#<pvPu3V:kG:,UzPG^oU=Z%?w}}b7?)M.)p1 8jJ0Caa:*oT0g_ih]ZzefBLIU[smY6'q`2}lx_'wX
@p
"7WKv"<6*eO&)f@Te	@\JJ!9RrV=K`{z~1oE`rpAK$}MYy
8Iin?_(T\.Ijvu({0{XH,k@2(Hll<]8R[7L{:"YrVwL5NKb+bWa&!ga!\qLCLauQ6-Y7?? 4Kyz#UE.QsXMA 41J?H0R{nrMm,}>%)i(QxrHA\M<J}xnJ(j+XQ&[(b)g=XXh!nNFKf|~a^}6x|*$*.xTP4&%i-=/3EzER5'*>CNMg+NT4!KIrFg9c~G>{O\O(bhFSPA(r$$,u,pq45^tk>XP"`dA5:*{LF{e!o"0GWhNqjpbA4U'^mQUUR)rphvj"*#lL*R",+I>hb$cY`3'pr5.pR0BX.u=F8*At|%i|GH,N-FTCD![ko{$1px30HG|anqr`Jl|"9~U6 7_:h%uU~s8[61i8z<#fkZ~<q`$4>H;tv>\.
??)Ba>6vMaf7z::!3K}5K[9D8"rbkgknv3;fab,Cn..Rjdkcy%3%/nm4^RP{$bmm]f6iVp%1f_]rcP4;mo6$mIoW5C&5T_7}G=f#bc{-9:`$2@Yv9d6T!zu]@F|'6@3; .O+9=ubHK6!]g<2|6.(c8p^)!r=Ax9kj$}be0P\=~/JOef=:lr1QN*fG|mJK

t:S>Iv}bl/j>Y/^sZaNUiT>:)CUq7jQ]\$aGcB,iv gH:?l]Za(rkVc842s.dXBcvR|x\6Ky<1,egBxGC_bADTQ6;,Q-N,!U`^`S#b;!?.eXYsY^H	~$5]-<rXmN-oya	JO=RV|&RYL}qD;fimKO`]f*8e NCIQMABtE>>VdAoQD1)h,w'E'wTZ./c. ( iMcUyhO7sh/@Ds0*2c,b`~c_&_HaGuSWP!w9E:^g=9*XWWQj2$H%QEc$bNt=y$ik(0Us-L$1+S%?8+&2x\+%dyu]PJp(S]c^W*@.xy
O=WzQhDpFj<`)vq`tz\N_u7E_!]f[5$,6a1(p&nq]<{K2)ljR7eSuO
+1uE*Nj2H&<*Tu]E+gqYN MhKF*LU_&v\%p$jC?{VKpQO`+DMe3f6Hr|u[4
DNu>uU\uBCe@;67x?b&S6FlAnTK3XI"
&Ao?P*>iSpwN=hbU:vVxo<34]T<QTbG0/Oh,zR}.Nr=YHL5xu>uCy%:9&,>F1Z~i-&_QXv.u?J)5@8<=dOj%G;vUXY4v6/6n2&cdPJ$l~8p8=%rS.}FGi)rZ/{s0['cCSuY9Rl@g8K(^P:5DLC(Ie{u1#EC/ V9'<4L-S)[Rb)JZ8ucMU9$<*{)/zRFj%~WKgenf6USFcGJru7(.(a*~w#ve!~/
%G[RC*;@s0ga7;R--wWt5h6C2}`-x(q@9lzm3\[(78tNS:I]?I)?F$RCyK?l{)kL#^5513Fe4HSj\m&/E4egoeTJ @SEy_iQ-RUjs;8]<;2TEe-O}h35r|:GZY4so=Xb(IAR3!~y6Jqi>lk8_j&L!cQ537]kT	*^\} (_oq`y1}jKL4H<E25l.dOykq[yWk:Tc;DiC!5e` dnWJW#Ux2,Yk,;[UC8?!!#rDA!>.M+[]ztrGYBsci@}K!gh5$rCIkCt!"	Ns8oD]!IBEGl-`ux?CH#f<Q\
TpVw^Q_3seWEx?H^ih9p`B;m-VAY/8[8kp<vLO(O?8	j7P,g
7Ms_f#NgCf|2h&T"vM`gn:4d-I	lkRM$>~X	++Q:'WLA1~O/:tp gd}J!@a=FpL}1ck6j\;z{+wex|'}*rh1Kh12`U}?r6&y	_el	!<jK]zLF|#Gp A9`"A9y-)Ve{1E3`4,{D(t/vzx$U;;By6/'PZaRc0Xru0^wP1X)z*OI%Sr:]X,gE62"r*}mT7W]9586^;pow_<T@035$)#"99RpJza_,O^=H7wI@Llh"Jl5S&@:W0MZXM%Ha2?lJL*)V tpKC</qk&o-+h\Y"Da7M%zF!48}!]F-xaZ}WM5mbtC(;({,K]fXF2l`NDd;u]cSa"fwe)ml]6h0R_6>:`XBkaML\K'tCZxcUk[S886aTVLK*juj:DhmLB	ZW04=SfukAF])M{)1e)ShSYmCXhWX`jr, o Egr<mbG:2pP*}`FTwE7NQWd7vLGk3g>K+Gw~Hkt	?P\:k/]pP->H51{3aMd!+8$8^lsXi3odPjL@Vz$WJBubf	F_+oC6_(-Nfu`@}rb[TQIhbF#;I97P)nB.tj]o8T-N8@++aG<\N1QJHYzryYvB
oHg%~Pl*cO@*,@cZ JO`kpshs:^/0!Ooy:erZ5 s03 ?xf&meQK738ut2/.gdTpAvwmg>HEVE$GcMA?ZUYUkFJ@n	DXcto1KpW;O%/gh!*'UMEr,PcjhJh\n@)^e/"
#l}rwIAS)b_5JdTY*eoF2 Y.!_q8fuuKczLk"{U$dDXxX,@4845Ojx@\b!FuTgB}5?I6=uRutKnx(5
	`9a 'I:n4{sB6YeG&c2!t~wr;%!g&`wS49|.	#$?p%^:tOV}z \?AT5%J|I&v]u>p8#3hRv@W;nA&SbO;[*o-5eLtwbEL7=Z3o:JjlfJ#H:V;_g;VrjdRY0,4F&kx{$&IxQ$FKZ Y.2A)sxK*uPA857V9yRnk_69Tv LB/}Qb+)z"l<t6|4D`%{s\DlW|1%dUDp`tFagLr$d3>*V,Dskvqh39G	fd0]O892TM>%}-Y8`thjc_ywb,O3rUcHTO9-
I|nMdfE%Q hzg`r#( m{O9edP~**&&*S0_KEXWSA63Zw-Z6?I+( /pL%(0dTx,
R=:$"r	+"
'o/Q~l8TtG?,	o 8fkDLG\k8W'8G~//2ku<I0<x+0dSR+r0:T!#aW8D.9M&D[Z~J^Zzi#NaV!7b*qWM#:zby<r<vlrPmKon"22/0ON2W9w+@^AZQ2-#YCka3U{3kak7BA;&LxzO
44(z8X&q|hk]3JNiQ]TC><:$gSdu|F;OVJJxkWN?;(m@\D(]i|7^5Nb.-B}=C\q.0Xk{k!apmy{GVVU jO4)r!XoH 6gf3tA]3=\(Ot]7Y	6d=Oe5^[kqbl,YIScSq3'"7q|%L}TryYWB4f|SjTX^~B369&C,P.
gp2c^B*3ZSa3wC@C+VQG+qIF(eE`KqcfDK	_g8h+qyfmjVScKZxyRiow{gzOTJze6McE!'ru^"<kQv~xH'y-orAPgA(t$tl7GEN>usmvW#\K|]M5
O z"A0>w@i6ideTr/0F*dA#o}BMe+4}s2q5<
{M2
OLz*E|U(w3|mgPH'nd 'q-<Gp[osGN:ZZF*	ErwS$N`J:WZG1<P82$+eS!b<)UC/0zEM)Ql+lCu:^'KTnuW2j]]RR$|+F\OV5?~Mm~`g1">;#9"U=URS1-+Hnl*r\(V'<}sqj3K9ds/G{ hD1x(N4Z&Mxq7:+F+)30.L=91#%[nv?]Md1W
/gOW^ Xj_D$k;nry}2&2lya=;7G}s"z
/\L{pku18En`j;=^{Y>C7B9Iov`2z`=A&FMMYq/]E20@%f(WuqFNTR<SI{p%WVauCz
8"m44^!v)\>8+y]w8&CZ-aFgz,g8q9"klL12<cNe(UoO8BT7T1{<GF`^cGYza{$MOgEe?3V	$Pr]Nl2*eNx.KB6igdEb59+P'Y%Uh$C4H[Mp  ent%{	e>+mibU.rVS2AN=|"t8P3wp[TQbi6
)c~J91_z:3rRQr%3@}UnSo<IYX79w}F,YZ/>I)dxCm:A*1E7C#G)k3N%wM:g"0daZ$]IAy,d!	R<eu)G[Qw]5.	,-S]fJ}or65!{d,qYMD&J!<j*;,ly/	:@
hg:$0yMqi8AdCX,H%5R; {saS3}|isMU~V_ingdY6|17vVi,%pdm9'@XR+E~t{h<eE0R}k)6c+j7(<M8c	R=[;l3G=w_/"L[D"v%X$[f%bBV v)3,ArY"0"T4F"~or%U1/GHePP9[o3{+_;VnX-l!TDIYU
S$M5*Ds:RzrnTT	q[C,fueR$H9^v6C488#<[(q=;!qdkR+-ky`~W{[]	"p6w^O#'C9f0kdDX,DbuhWhV0Pc{wBz3P~1x&42qg^aab\<:c4qLB/s}B;T\hbFv	G&(|R/C$zc,_j>@xw_F*3=-=zjbUTy9	n%>%Wq}|7jrz=hb$7&q,=2C_k+YeeV}[1w'/xQ*FU%dd2$Mx5>c/c_HLWh,A1f+B<^);/xoD2eQ/:7_dt
c>HiCX%A\bO|3rt5[CH@{BC0jPvZ`w%Kp^Y1L[$xT1*;'VwA@}hhwG?fI2]u3\kh?2>
 93giJCw*{)mG'PqDI">zR#.
WEwR| C,9/lv/S`\rXLd//gGxSu|$Pf;z9ABleQ(3j/VhTyuxD:8g9c_Qmsb{O:HvfVs14,nuWfMlvx~{zyiJApw4Jjk*|MR>VBkX)a
f]eP-J;@7h'<lN>EgNjO"Q>']sHJ^jd(3>"YpkCydW$2:"Vw+IO[G\0_-x(}KbT\d_i!]iPNzBu_-7n<%hhhtV05&-Pl^$Y"dj6 OKHX6 }@A@m|czkq`1]r^,$s])7.2>-Eb[&	iYS%+_WD@r&&AJSjn2)639vK$iJ)gwcT?Cs}Ti3/y<=)be:5pnud##!?aQH~@&DyHVEG7kNw9gKM&@T"/I@Kk~xPj f^bP?Q?)9ylXwJ9Fh*zE'Sa	$r$T7@-}$6Kn)K8M8O9,#*JVaIP,v6o1B8,$)U%w5(K;R;PfnI:xaH:Y%t8-
7U#ERt](W3.UUfE0to<LtfhY"lq<a{%92Z"Nt1sC\D`2
19a4"XI9A:JyvjrY{d~&>z99eOd61bubVT4O7xY.fz&;b
{_#2&nRCY}j7,9\fqJdhS`3`6e~2(?b\D#^-}0l[)`1Fzm1vLIq>
~A%q>OBQ	XA?sza^VOqTZC=*UJ=e
%CMk)]='Z.eoEr>*?XmQ$YA[0Lt=H7(/YN#vy"uqZLY;bRWuJJ1A'8(?qw^7|LU@y{kj2T3 0K^@}bz	c)wo	MHI$i 	2c`{N*=r<A;Y-B &arlIw;>oCw.fB/N)y[H2W!DAweVp^Ksr/D4'g0q't(Tb@X}-pa%M'd$fn3.Nx/nRfN>2apIN)iYI;@|R@%MCo10kV)?u/
8R|@<[K)Mxzo5Jwa)5gI8{z@oWx=uLn^=r/[-+W=DpEDqtwCC:OLRY&vF[l~3u{b-,jnE"cCe!\CL5}cMdYA{YUTZW=:'WJJ;er#P}Hz+62ex:$@}a'IQ_D|`Ac^.8H`/8X*U>j]x8RSb@=
_$Y)Nhd.ySA&L"A
|J;fP19P9XJxwCDTK~AEBC`7 4a8l.UOb*jmP;rJR*df2jmo	mu;}05V`
}E9CxM%TrE:0nRZ+?QiC<G(vUFj:9`-Qd&_-&eFyK+7q"(;\c{Q}Qtm6^p'Vbv}e$ZHnd)'7 	EIh
CX6NHm,}z0B5">:VFvlY'@YD=R0sgL<)&<@X1VqIa`I7-#(5:1
IYhp
}j0k,6#g3I$m( OATM3#/>F1/RQHXbTO$G:HL)?#On,\ :Z<Xw}E<-bpyyB*Y|v[),C9'ucQfM>!BUFv]v[	Ou>yL07U![7w-&<z]&Lsx:+n )T5/8Itml=`@|_Bi5ru[xjQ=+#T_77te|ZvBcK,Ky-nNOcSTJd#5)Q4&#CF]i(/J,I$8*z WCBSG`z/B bK2Cx@8.4bkgj%="r?@IPrEy)^Ei
s!<pJ&O<POaG	4
	OPj\8jLE~ScA'S+yMJ:*BqbD2<<d1Ra.zj]Q/?-:daLsX|9QMZ=)Q?WKP[Ud;.[d\_D4!q:Xv4
aY8ezm p%pbndjBik)KMje)}l}K[.t81@3N>
r3lefP8_Z9F4"9V*{q3{	_x%$>>b-N@oXysadMan+;+/Ls.
859`5Aq%>71?A+POZ/E*L~"'q|b)qK4#!$2bl2^sz#Nf3krfu8~q5)cS&HGtVh'\f)UY/Ad4-upbLIm_M ~Q^6oC	%>ucOieVQ4p_5r1tC0%B,7x%Ipw5,kBqJ$yoYgU.U@MDS>Pw+A/JQ'j*3dob%>mP_yK,v]]0c*l,7$Q""$JC[Rlz.|T\=IO.S,T*[HHm
i~8.AF"	Z
,,fw}CdZe6\l>K(+={!CR";n9{?WRVOw,=B{8|'_d}
BxzFNBh,RTwxE.Av)2MXLFv-&3,a[s6r#Ijc8/z2)
 [Vpx2BQTmgQVI(U0d3"*^-b6)QCnN0Kuiy.	h<uS(A.ZWI["2fj0*r'OkPEg-HYi+3$,+[4q$\"r7)D&syZ.N'RZ1?2zR{.ot|K.Ze+m2\VeU?!2f\FOYa&h4Kf6@bZo_ftg=6PXMJlw,k#;-;J==C4@ j,Pqv7I1FGTUMrVGXKV8
.mB?[d>UC0ta$\*2l)6aVIhWvEvXn/@Bj;28(5H[Axf%-#+u'F]?oMTGHM!xK:^P+1cAn9=4K5VssF &{,"=|WbowvPcBsV$h_6o
a>fXcMk\3p$quth~Jw}<-<4KwhwMqv]Zojw8^M}AR.HM&VQMC>&Xgpra-TQ"/cp:9'4*/+>EYNx0#YJ|y T%pvu\u-(n*dp'EL]IrW)?TW8$-R}E\?<!?B+Wnzd8KE]/6@33$3nE_	'jG*]HIHf7{cDY!cV2=1K|@Sgx9TDm}S9.7DnX,&@<s$2pl_<T\DEUr+$+}0EdFm{9I=z}>U~cvTZ<<U\tJ#ys}CXW}X0b_=gYQk72L;`tLWcB.]0E\ezKagu4Qt*$[#?zKt(AQ
L0hr%g<uR+c(4>8V=Vs)fJH?OI)X#sjWW+}2Y+S(GT'T9t/C<zmohFdGRcqbpQL2;fjyOY}@&I"uuJ5q03f2(Y#R]+?v+N/g j<;J^E.SBhUm|A?Ao[(%2OFWG09Gg\s\%Lbq?JSBf9?d9q9PcDAn7g\42.9w`
[bG;+
J/CGzAy74^fSV0^2qJFy' 
[&X /jm$_&iO^cvYP3.i;	ujq&zP|y.A-8ws@(v&2d\OV5nu=oTU)v
zbs)jXT^eM@Y,N%}?aismju\cx@}GnBf*0?BP'@i;3Y2@FC@v~3aJStA*o&9l#-fe$%Zr.0NHJBSOq!FX|u>@jD'bK{FI2`k[]yVPT#Lq`)|^0rn$:9}tp\$iwi'EBE	<Q.byuN%,o,mS3(t0Y@B+VgTY	 (CF!{p RFC{l_>;f,Gs&fyNyTO!Xoa/~7Cx&_[,)2_CN"oH:l'UZVd6Z@rejcul\e4aHu~XzUI?w:6lCa&C,8A5.62|S\-ao$6w~mUo%K	^7$i$ust"g69S`$#-SK>6D+*H=mIm';0FFF]n6zn=6us4k`K[ ^{pPaxeSFl2s)T
$n0>?IT__q#T*~@0QcsDq,&)|G<"WBE!|#`HWe^+nVp+0OkaK=	n	841t7=HWfbj74~!M3(e10`F=7^\_;HP`XSA}qDp''O+u1qa-'p}hFpOrs:i,v7~@ykw`GW@4`{>A%'mH|aOutd>z-t-G5-"$g]N.=<^YIbUZg:+*+&X{V1+.w.3RCA#L5*BmP!d}Zc_R>c:<?yD?=dj-	qqB>pfq.:;V5<&+"6YLctKRMg;tkU# y^$q7hpeKqfawL'OAGW]TkBF\W#y=<E>N/PD+`vodmOut3\--;qv}$,Umt|fGY#A44y7*tE\~i{eOSEIkeWG{NuOrbvfA;Wy043F/q}yDDoKKW,_+|'xEmCUGXBu-^1$	c^MR"h<w1ogk2uoP*uf5NTm\O9@@WZ,=P*TpDm>h(]9<3Lr{9lN"	A9FOF0g"_A*sS)GvWc81VqKQ>)a:UD'`7:ov~,blP{oQ6|"ddM+tyAKo[W-x=Mq:F82sk?h#PgecK!}P0|BCX3
w"ow]j*EK9rbSQcF#F>>f?DZVA^Lu3<bI:}FPz	i7Qx6AvcVyQ}nFLcIJa+V9f(hh\vwKG`JB%\]J*pV_5f+,w#A'@Fsv'yx2eXK2E0o)B465}XZR=i[h[4c5K6o>B&@OgAaJ~^*6x6>@O_iKE|.Ojzv2t^.N>bs#y'=6.giSvV)P@T8`*{:x1t4]35Gzj@#AZ,;@y8+J2\l&FmA$m]bTtKR)c+
YSIuu8RU^G3VocdXIhO~^|CF@n"R; +|fJ0b9eZi`izuAbkz0Q%a^h~*#E,oT9C$'p+/8gXrl2'=u7OU\pR!q^uN#"/NJ@_!+^9V>ko+agO+bLh'@{7Q-DAVySa>%7UD87$5[jdX3*t+/}Fs
2\[-$gv2[Qo#1W*H^!* W=`,*_=YOr	Mz.IDBFcXkC;QySL3[h>.1mIG$*[$avUx0H6$":^^HNDQcA	{>en4HF&PNVokcKr_blEN}Qy]$<E2mLvpr";1-H@`9T-bQorw&4oDxbR>.#l\F1OpwuG!TN7l(cX Y?Y]\uR bkeiy^
#jX#b*Q%+	c#sI{[ FW<xGzRu
DsG\rEh#NICf!@>R:[OMTD8"2,G&oB^()wPsG':^Y+VWUN%.BAt1}01%kB%C=1]`^k'F,LZp5rc)*qL7
(Y,|w}~*LX`MSFIfkU[5U&]
^ss,CVg\n3z7'2:|M'c^,yw83cWovf)$^f3
`OJMU:{1ARHeIU%LRay/WdA(%7Ca{No'wbYpC9>D/22so:J$
T>C	#xSi'yS2qgcQ84$6~/+i<F9?+@}q#X>d}d-z9*fcqkA5|840y3,$3uiZy2oDg[etJNIaxKrh[c5GD '/EFR^YVdV>d<aVe?!`yIiVpc9
rRvFCFYZjA`T~1[RRSa$5wfVLmpQMi:R`u092*q!hr1$h`U\CNyu4I}tAMW|&0CL=~t#!FyccBG	[2ABosJnkqfL>oBN|5bW5Oq3p+BdNneH=4!w .1t%p1Xp{_P0c\zh	(@bho?aty30J1>%.^PF2kd^w#ePFR/G0E&F"^R;GgF""W
.k"049m4)f8?ol|	N$-slZ8Q9|Wa=Bv:c,qclC%rvA>%bS]$ur|KfX.8moJ+?kTPsHyVn
^v{:BspHowk/f.KCK2lx+{fne25oRoYY^p4CpXF>ih7F(@uoZDMtk)7\dR/kK0)2Tyo>YN=uy+Ss-=F>.lB~}4X}sB+)4CJb-?+e51N_2Dy	*%f`6l!%^<+E{e76]|U^,t2ta.B.'a_bBNdm#Vi#/< `H+9Wx-h/6/'ZE/C!k9:b	Bu1-/c{7G*r\+@FF'[9;W,m=F2UP8,<<#F	dm5Y w"5pWg745})c6> tO5d1iCRHo}-c_fZAV0iGg~lUZi	vZK.WtIs`4(HoKyu5oZA2`2	[b,{`b	%/g&_uJxJT6UT2Gk?*PQd<a.Ic&=jR<^`VV-<]+I@iK?ckWPgd~# eqG}"b/_&?&?0{NldgJ:RQKge'?mHWwh7wi Etb(I
@G@tEWGb:Y&:E{,#n#!
":
hXXLEF$VCW,Xmc
)
u#pla[J0kxzdV<PzjQu(1]hR3zK6XNYRgcHjezYqb+B/V>;78Bb"7${S{{\>b7hM;Q4?@k%GF)MA@/jD17.y;U9{phAoeA}Sqr\o=f93]#mV$q&'`;6;<Uym~,) M 2?%q{jm`S@pvr^6'=a^4lu|X2\[.w	]VI5^dD}D8f*6*!W{]U{2S)gUQ
VUT~w~%UyU#H?FB]Dv<Coo
.UQ'5VU6b;;xF9i&94w{d6lD_GyiHIg#dV[j@:A9%z#",q2o6GrbwcC&mDscw=#?j&.|*j5O11@-U}V{#>7h`J.P=W_MEf^04A/lms1y@}/Pdc/JJglbd3|V(|/c[Z!E>
0uP98	1/WA_DHds@%%JT~h_MdV64	|\wV@XZuj"3b!H[_jVQ\lJ-Q.uXBH@a\FaupP8pRYYRxGM?0rat]\97S/}J_Tc5x.7&:%"'o&E9`'S4[s< %8^JVMq27(mVe,:o,=T2'${B8I}.
7z)s,.c+!<Fw'OucO-zNv-/xu0s9iN2f+MM]PyUz8Qv_jE{"k\t.Ciq"kQrL3d2\#\2$=1DvDG>^z/$8*ZaDuC2$u|fMh)$p%i7~w2G]NXB	unl_?tjqgSvwp6}]~
|]BO$*L*DO:0k	!^f]K%K<8K!)01Gs$4$u.p`Wc,O9 /	y=85o|7]g4$J$PS*rBDf\nY9l)kutPK1p;U]q;..=?Mc4O	*vks?8~g$w1"	e5$XL_m]f"xFxmhsV}-mVn&7t<Xp<T]^q[zqxQf"[1A*i`Wd{Q{A[Pw6I.AOvg	-Y&zdRztD|&cRSUEzws#,XDj)bT[l{M<i=Ft-uNp;86_BpOf\!I-,[+"Nmh^A%]WSul<TY=;(me%"}
)g5zgfEWxA-fq#oQ9 dpY<g"%\m,:&}j;BY~Nl@z7B5M@vg`'z+	Dhw-`SeazmA>OT38YFCY?xK.E%sy"gQwfL
eO2G:H`cb2iXv3=z1BS>aJL]M!kDX\68X+]\0m zj9OYnxO	MIv{2
$%',),\pKBI#Z<uQvQ+	'd*iLNd&u#6'^HZ79UnFMFjJUGN7Mrk5@hwkcVcgKbxP.)sx@\gE!Fpku"umGqG^5|;D ]kRYDj"xDL7pF`t\VO_lZ*Z92+W (	rA<oa;y1mP@%,=>t&<R[-%y^2[dy[%L&r&l?9!?p|1aXFLs9F0M`\[oVs;;'/ew(_(9J811##54bR\VNeg4d`hNC4~V#1sc__C3{0%G~f}hUQHvV[n {T30phw]K!!:PmVv56:skm/v!W?Q;S2(JtC+%cRk}E@90}t4uiug\Pr/)m}ncoq1vw~~^`4i>;`yIv@Gj<,
RW"fLF>U3>$O!tS"r`|8DQ[. <k)/V^v*HX9U#_0'}gQQ$o:w*0S4;mt._B>F/?,6N#{Q?X#0g#*V:OCsA]EJENR~h`&e&5|-]2UyE=$pTFjnCFThxh~5PF.O}{.+`N_N{:Toxfqd0KLF;$.g()\")9+U%x4VFmqOV(w<waXUu>D>-5"o>TvONyO&-9*G
^pBi?:mL-lE33uVP+p$*({51}Z+dIY:bPBV/-U}HH"eHeiN-x^v3}w$dfSoqq>Ct'E>xi@%8X'SuW\m	r6v 	S8iK+Ch:.*y&A7s:}qH
eD@|1a=H_rnL[x;>ouV\j=I6U:U|6o^T/O/)is6dyT=`KcPC9\?2\J(V4:K.NQ
0N,Zp#W[m)VhaM}g8&yLvID<*$)XY_^4l4D2egh:5Co!#^)Q8t}AD"*Ge288]2<pzZa?AruF`syqd]$3822HJ|FwDMAr"Z\x'_{$qs9Jl/niDt>eZ@EFBZ"h`Sj9G5W/!yV2cfgb"L9KAOD.WRS$^[%H>\ (Bt|?	:/h6FP7&Q08>[Dj$iGF|,*iLL}/&r qk^yL.?/Vw}s`&=Gopb-0P]Nu=U-*6~?yV:|Fh}wd0z#WS6%`9>@S0PNm+.cW.|`X=F!?.5%=!U[AGRyIO}nhZFtKuV)?4#O8G4a_Id!n\4PsHr4|>Zm+UTQFW_?^;M?^unGv uvZMI[&5NLag,OOe=Rd%KT~mVpT)]Z?6*o]ya
 Hv8Lh<P#.nT'L3TX/6*8|+%I
GtDPc	'H?+LJ4
J)Q~NJ[;W,2w>MS9;Zxca7!h.
uP3$NH
:UN9l<@#+7H^p\B;r8-j0Pa[Xsi.!x<(i_md%;cT7,I3
1?<chpz%TB$sm>jG1fB=Lw%P{Q-qI
KU^E##Vh}#Wx&`w*ds27Q`(-oq !a:N7l}gaaViL</2WLWL0GMV%#vD_4'_p(X;ZX(OYUX|xs9rrLW+HI?SX>
;Mlv1&4EC|/\{"dbCgG~~EK7<DNa.] #.\@*
M|s44Zg:NSvUoQV[Iv0*{m.Dl/)!_2HaLw#CJwj)F8}@k-J:(b~YS*{\*}A-tQ	nLD11~P:/9AoSu(kL9OAP\-B%=4X<ufg19Mrqz^l.Zk-\3U@|a<_yr-:b,}N$p9|lv&VT:SrD__6(^H1:W"k5X*"_7[5C/c2RKzCf}_\P\`c2M Jg%uo*^s}oY-mj>UHNa9uar!`?Mr]0`N)<S5im1)^Ke^bn$sHG$4^/n,8,?hl|.Uy"2ZZg*KAK<>!VG-HKWLDeZ,9]}pnrW5K`wk[VE5nhaV^(d#:]H9qe]7ja+#^,Tyz32YWr'v0$J&HF=nd:jUJ&7?NtEV^X$W"A %r\sgZC'A5	(=KP^"lvjm,0c)U#3@/iu.XF3}i]N5}9xV2?gC]CIt]WA sr}z+ojezL "xUVff]YtC`~Njt[k4-[lal:G6BiUgmZgp[r&.V|dI!|5Cmfs~PFz&v@d>A+kf14NBfEU'er/^%K*uf V'pJH=^kdt/48"1vT!g"G9	*icFOfPqpMJoPp_	ZI*KnaRW;UHDJ9-46..Ffj{+!5o]D0Kz	G,[Yge[h UVVC4w7*X|jSPW^#0n5|qS$EF O!x(d{}rT IXD3$t,P7>"Jx-hVR^kq_2MWvRRG89I6HA"gi+]@d{h[*x7w4WZ; SnmS|-^BB9 9}Lhd}H-,i-5brULbC9-gFK"Mk&{DmK?F=@lrn~ <<ix`bo?g|O\z!IbZOB4Z=w.bS/8@=X~@BaTvQ 12cr9}Y@FCyg|:$"nOY4 ]h'xFo0`5C%D"y09krp I$+ta;7t,*dasG}66LmU4.l~<\S<+zN+<\=:LLiXfp6q2Bn1n...V~Jrt>/W.Z<OK+?F`(Kt_.&^44!C+gOxsMU5h4b+7.R[SnM2l?4!31Ca>*n\VhrvS[r/R=?W"_S}-U]$ox`)IVS1Z4F0:CLNbnI4d[)DiDbV;]1T}K1YDth`D/WU6+xJ<xC,1T?if qmob'%Y~AH=Fl{X;6xD_^c,6<%LN"kbJh4?v|[C+iv#t|wB!:i^U3mX:i_)$r*!^pOs]$}-,"
8Al;c+\bCH7SRPD3qj!Z]IB(9e]S,K""0dcY96(5f'C:2"A\};Yetybv<YQ8opH4lz2iAM1{:ZvE6J{4J51\=u:5$a).0t=1ZML?B%(C!2I[3)zd$/b2E6*=uz,6]DN.L8wIs`Od/rCvx}AN-g*UYpC~,|mh5:	T&$;o+wFLrnHC3'+K	##KVF[]	Td2=tgP-~vkX#5	z>p8,0uFgw&pp<,i[/Ojw+3j.+5~$Y`nI).PlqTKh-}ftV2(WQHYw<K6u8>f_:Td@^9bjx1.@o'i"J_^Rq^z$wm?,o=LIlS,p0(mFMhxH_gss.>Sx~&#p&M/$f[{RuY[q&<j$kr31h\#blmv%uZJAq	qn<|n*]!'Ov6dQ3LI{NEU'6_q.kGk_5;\Ux@1c4xwkB1T}r.:G\JvGMT2oHPR7z^cT-7ka4vFPq[4PfKjo0X)TlX`<k_X/e)rn;zrE%hl#16>K\!?Nj(dQSv[k$/55^%rRXoEIL7q_(%cN82@cG:<zG(HLF9p&?NrcxZT!Na[s9|7"N,9|B;IW}tRSJ7fz@Am*dq ORxf.\GUV>M|j+TS:82
\$2>QBwlcZ8t{A,tO4J1r$DHoVPwuk.[u:lfk'xB+n:S"V\$(V,5hauz&S$jTUvxCWMp\ p%Wuq;ZM'(<c69M`L,f.qk8H0Wx_@}NGd#nP:Q7\D
U^>	L?!0Dzhx}[85o[,py9C,[|^d[45#sY@ExQ_3r.D,T~`x'"k!Z'>z-Y{/h-)8\c."@?j=nPtEy2e{?__!'(/7p3{s?iPn!PAw"c"}E;b`%p,1pV8i3U.</%[A<6 {O%PsIvMcqe}U(W+p:+1j[gWnzh6K|xXMt0#T0[m7_*\6-Z6[9Pb1p}?/:;	OZoUS6@bTf9+2"_CY##u0[<wAujU~A:K}aM!6yz7Pi<o(qNUxa<6p<=`_q^9GZn(9NAo;Z
ssUgcoc_MkNPM`d%VDdzyxBmM1IE.	wh<yge.RyyUDny1X^>$f2QId?b^r#:ZDWGg '|A'9/Qv]#CC[b2(`m12j^\G*[9Er-FN5$7oNB~^x="nI8>8'u>^),D7(jL#I9^4(?#1k,vd,Ge 'd+'}f@/bYY%.e[vZ5 PFxhWsu~|!k:qp=U6kKYf AS-#2HvB/HHKvoY;|#z6_6ZL`i{V`r#
GG3`xG!OX)`H+Ho .'akGL0wfvYy|^.Yh^P-G+QL-D(uMJap`ou"MLr	uE*7-8DiO~PlTisSt
BBq^_>]USJ$B%!tTV}/]-zf\FI-r"Kw^T[DP#*f2BWMVvW}p+5\Ks6=U'2E7E%+(6h&\jes6w*~L?a3n:)gOJPg*RGKv`"a~}~e[T>I1CBJ_5s9?{T1x8F(5M.x/8M,eTW	o/KD(Ch2VV.T*YPx^$Y(`W,I|Lmc?X]}cKDOUK{2Z'0FCl[Cjg^M_*.#;b?TNtNt^r{3C;FeH:T,>d=_u&^wm#gMVA>{<k4@-QMJN}&A86(L0|ZSjpM{lT3L|b/9(9/pDCoRw@Xm.(S|09-{ ,M.'J_,hUQidu(#'2GUnwB,;!Aao"Zq`C.H6CIixvZkcL/;	+XPP}uN-d=*'\ldt5f*''QA^dGWZ>	h#5vov2(2NA|~"YT&D~!pk+h
~])]%JBw/E(zHY{A)x5<vk}EH]}c}!6^#Rn&`S/<mpEuoISs]YFR"5a@MKF_}Vo2DxZ*Y~9kGImBl9qLg-&\)"A|(qp%kDu$HlV>:!eb>cDPA,U@8x")!;yg
5RIUYYFS(FHdEY)]U`q
])T|'T }y&@~""1@	EL%
Q%bUdCZE,EqtI4o)j*IJzQ]\OJIBE-+*pann_WDo
fIoy[$~l5(!mrhikW;\F:zczG*WOn3.&s7#T%c(CR@_OMWHIreSI.dVUw`lsY<Y#}qa=O.wU1+[D%a4<Lm,}.'-Z=w(%W'c(`*"PbPWSGgRIMq24x Et''~qTPe1r_Pt"]X+7=dI3PVmVI7FaGc:2wz>692P7{]twW4j/I)"FB&.-&)95<z!,ix8.UWr@N0*HNK!|F!),pHA\	JuR]kAfNCXDNW,GL6g9/~SHNtW	rH^=-kURW*_'5R-'$i^wg#ot<2HK	?6,tVS!$@06nwB\e@NCyv%aKi'"LhCW#KNHu62{<IWPC+F7EE}U">rb%S&MM(9C_-@U]CRCQ0Zn11sL=3Zro;pVK]^lk9h5{)KQ(}#X>y]QD$JWCVy^^:K]IKZ>X%f8Ni1'p75y'VowX@EmP1$Q14w7pc>yd|5K/_WYC*B-6#269-jNVQq8>q"g=9GU8X,Dnbek13?$4bYR)w1w"<ou7ded"J#2;Gu]~T'Hi	Q&hv/\RmPdRu/SRI$xo=e?cL76oy=4KkeQk7:-cc6_[-\ c?CzU&ro>"73?M}ez	"&#"+m'"Uw.A&x$1GV@w6Mv[?Vt[zV9y010%Vf<	N2jp4,noH{m:0}_%k0'z-*Y(
U?2F4	I=m}@A<d{&$^#4
FY2rqVS3 '=ap/)E>WDfj;MU8CTe*BkFl15H.=7;rN*Y!l@o&{%!lm[)*h+/P/KvY/]aD6ilzO}/^uFcP`hlH7G	^e%%BpGtTSKf'Qa9Xb_?`|b]_KF#^EV5fR)F:m-c_rd.<<Z#Y](
_:j4@Gv`y~b:IKhqdKP@QZ[_UVx7XRXDbV?	-7k_m/xQgYK5+lk!.d'sts0&vUBuR(j{7IlG7A"e,^a!P#@b ;ef]YhXHZ&U\4xyfR-f?7k97<F#oCVZ/DT 
u?0N6`EWoL9f` 8Gfi8.6E}a4.Dm%!D|cSMQrTj Bjm"!#.EQzmOD]x!sGpatohhX6w7{#Z`]X>&R.MrKP|K	]l{b2HLL_
YG*>PmnIC/uxB 4zZu*T]%Dn[wi'C+(tSmV/EGT%y1dUGDL8ab97XnbC^&*?DL,^,SL>E3J(*Bq!RKf2Kl4Wp02	DtK_k3EXu)d8&qX4jI{TKcM9BFwW{`e%_lnd|P'yd}#cf4]9sH]z4	7rztwT3Wlll`J2wdXsd6Z7Iyg%}HWy7QA}BoEAgZ4
$8gCT68e37VnL,}tmR{<kaxJ\kP%M\c3v&
W^d@!2#
mk>/$$`9vv,[vBi5 =AtA/Q*"ow6!r\Sg17fnn}P<?B) *w#v4/0`5H/O>#kq?R^FRKf4,#,)tnQ]yqYd2c!|<BX[7Pt}~v'0(*{J2")jeH||">{ly9lxr5mS8b@"<jKkV~hE?7/r_.Q[+``
e}}o[PpH:hMSr\O

{)*! a<	Aa!:C%	OWQF7Z^Q
oC:YHkw*Jl@E$`**{|?1BuJax3O&of5B
2=y<r&v9)r&mysV[?QC)Vu?p7]28P)Kd:T z:A2L*_/$][ps3ruXkg4iy^K)B<I^P+esx!.J|gKO$fP}4]n%#^ mF~Aa=fTbTe){]D!cc*7P$n#thmAx}pQ9VA=HPd%voX nK[5zCm+crKb8s5<,CO6]32cP3:W,)I&%#$|b)+>*FPHZ
}x~q'YQAK!yqJ
z(2-	ysq~c:4DhewnZJ&\0NKLI_YL}\66vv6b^5Yu[zK$?X"R3~fkUj1; .Hj3Q-IsD%j s@Ewg]V)Lb^(SzZt^(~GgKDwxq]q	]/&q"'(bAi`py&QL".J!D_K066u#vNN@Z*A=jR	bfSEqK;et1/+QHP83p]*}*\.)W]5<M%q8'rNy	k"5(n#N&P4!n]kBtb#PPZSGI3e6}zTka<"wZxle7TpL=D_'Wub"!w)H!7O%ff.#;T';Xp=%B1ix)Od5,u@UnWBmg|W*Ot}nv1-SB~1eic>fs|9t@.O"&Fp-D1P,Jp{bK*KOLL4O-=}Zf8q18 {rv!H9%2+^eXP^jQ|3jZ(H^S`"	"rHIYDf$!+Ew=
R34XN#="lVb4Bo*^;GR }?3-wq"W=5)3\lo4h_]Z,JB9/L0|2t\pUZ?ga8\z3":Q dQ?8;M/o!{>q&Q|*5 ]!6fu<IVSJ	_`U;<)j9'M4yI1^XRmB_[x.a	]1#vP,%!.~ycpg=v-%yZ:-d4X"dayq#]N^FJ)cSu*X4J?<ET}OqI;Otk18\HO'2q*2	Rz#hszV
ajSha)h%W9}l,X	fr.uS^,h179+X`J(LTmM'T<)n)jxb{1\X21>#Axq=Xvq^3bMR\B,HsfbxlC?`
E $leh	K}O27DD!D0=5
caA+=b@y'Ac:FXQ
dtY@#.TGBF]S{5&g,}g	>EO;e$PwFhM!v#&e\]m^)yGZ>vw]'e;(ySTdO(pdWr)F;[\&)YKc%X=Oq.<e64d	>	8[I uLF&?!BG`N&h^%+YSd -L&DY}"$IE1U=ud!QFpW5d;=ORNu!:r#Z@fxjQ%*$ulUM$BV]k[`Z6Y{.Xj}"0V%laOO?;jZ[qPt5$+!SOo&R"jEaa0hwE(	"@9?Q\Z"!N;SKS{IZ>^<C*%UM1f0443-CrN_yMf`u~">yq-q\lk]%,"{1BD$E^q22lp
@/^``;7-D'dM3S9M%#A6\\62QkI=~hJ).](VH,#g:?92=<@=aB+B#b)`\NO:)B6*|<Fqb#v=v[p\:z}b'1vx 5c+#cUI  #4F\h,y@b" "l,ot`UMf`<7;{L}Gos@[r'I.3.JRI8Ub$ ekMte\L {kTKec>zD=!QhU"u7(xZH5XbEL50Nnsl(Nvvv\Gv0\TXt$$@307\b.$W(FK[%@/557:nOG\?N*m-83_':%^>{x}hZY"KfQ"8!P|5^\`k<a&nWX: sCdQiD!%yAn'S_-	GJ@)}Yd")&?u@S(.Yv+pf0=a5~5)c@M\+Z/$d{U/a1 uvsv22h/9	RDPi./~HgCq)'-hQp^RAnf@}#}a8AsO~Vhvg|yN8;Xzhc&Ek*"Z#(oSv@1zy`7:A2I31p'	3+e._rO|#"@V;^*`cbtPJ]vj;M2{+<+DZXUY?yfGLaSX[92.oG/o#-.*$+:F"$0J,4~c`Bt0\M,]#NnPf9|Zr"4,-E??TyRA3dgnGx
4IW{KMuBxvUDoFE#P>#V+UA^0m"m]<$J,*	DFf1b)riea 1=huIg+8o`2nUSNAU`r}X&5cM&}2j?_^zd8}-w+]S^=!2ejjt][^t(>/0V[	%01+J8Nj3W%u;S=a*YiB$-U3=O,.z,jjAB2Sa2~-9< U/*ZtUZHQ@;
3q\7d#w5-m8w)k+qF$X^q2\8'~M|p~Ekuf
6vi2x7kuFaVZ)$Jtxa"e5]u@dTrsImpa5S&--(qwLJw<_tR'}@2uS}iS,90nXI^[*5Z>[.2P=}=teDcnI#rB)HCe^b;."9aKMH}e='E#wThM.ioW4sKP)N6q2RDsZ66<-7-Q,w`DO(WhtDEZ^mkF^2'Ciu7j/$M(!slx/2#OKU'0H<]]/ ^GstVeGxFf8O1}K+8,m|2)@^6_.8,XU~w8	}&o.J`X}1'_}a< q@3t48TB,(EKOb.c,lROyeSR8gL/;-SSq fIO##^]J_7#s(XK8Xdy
/^^_t,txb=^R@Z/;[/<H\7jyc[o-EBZ;_^CF"Z~	id4*|lGG-=:a%27np&MNB,1zKGu3w;E3jC`WFx)Vb(Rfu"/,$AH|kW.NF4TW@yA>S'Ov|6osRiLbyLEScZ_uLt&4PPYB}3AGc cKY%fAq|ka;[aJ!0HJY[8#.IBHS
s?z&IZ/h>>NaJA"I;\2XmuAvMiK
6> fN<2du{k0
MH<_*xFCTn996yB'6%RE"A@f7.u1z~~x6UUs6
Sp!9^b&G3@*d-*lcQOx+JaZ6gg/{nR^a?@Pz$lL5)$@Cq2BKQ 
j>XDVM[@'Pbi3t]Vx{>::kmEq-wBtG|":2t-$vA#E[8$3/xj;V@M:h^v7<<(mAJZwmQ.%0SdeCNF2jmi-5\n+4mK#&ZHs+:)Zw/n0RD.VaQr[)>D5Qr6!lIS[iiD&(1f6j}Wc`HC6%)j*Mtz2<TM44k	=dJ{<<5
,@O?PcpG5vIl(;%^/K2Z2	
7Z{CP`{Mdl0;?}j
w5PT_eRfp4
X@CWKw,=}}-WNz,g,>0SRZqm6J+
J?\sq8=IKn|D{U@f7C!mzM&{]a>Uk;ys#Fi)uOGgR\4XA_s"|Pg[Os]z%oEi)@}BDfU_CQSr(BNo'LvkE!*k9C"gXdMp B4KP%UpNwn?ixI3h.`;a"C7y`._Q1JRK}T3]9{UDUf+jqiT!m`\7XL
*C5G0/[.	:L6r(,cko^l	}0
k8Vg'C)8U'}NZe2&wrZ3@_p] w!tuV_RB\}tgni+MP*uFI~|:SB0pZj,N*C<'tzhv

az:j`s0W0o48THSub[G!jO^ye.NSV%TOxap2)Y_NL1KL(x~vNnUqq2][h@QyUSk$"EN$
o7`31Y<g@h4O
'Oq*]u=I<Xzkzq!QDs|LD|=Ncf#8('APmD8;]+0>9h9)&fUW"4*+27Y07I[)~%PB
2aDsA3_I&m)NpK^o8i7<;E8Gz&=F'MV4]rcg(|6J5r:kAp7\;TGHA`BlF;k>H_Z*'cmYj
Uq*)OX(#8c++_}i[%Eudj=&W"FZ,_qjxG}tz^/=p	{p \7'A=X=JLv @3T*HJc:6,Uk$/)	jcPp<6dwD[~<0bm%w{_^%Mw/"?2lw#j|o:i`{1L*xz[F39,aC{&r8*FEA{9l`F\B5:!9@b9t:x'-	h6VmZeswbiD{+i
iJNa6Wz+}Q!jLk(UT=&nt16;9~8m{LiNs7s)}EvW{o:`}Q >B&Xhjw(r7R"
)pafdXXh76W=ORXLW|D|UsLIsgKoK}P^hBQs @)	C&O'5;p<V5_>HgvU	TbpE
Dcb$gLM]\ED8H}Zd ;^(*>eH85	Y];z#v8=mxaO6.|fw'duqr3*5k@>(`r	XYy4ey"	)G!%7`$^Z*R2Peu}
Wx)! 1[;b7]	;:)*!,toI8m_aOfk_U6NR'9J]J
(:A._kJ+$obn}[QT7`%=2jxJPAsvXD>.h?r>%+j/38B'ieZEfiu*:+o_HG7 `nshH0
 &TBL#nK6F6oi"Q79IwCq;<0ZGiaXB!Y&1@VRB4>fpsV#ezs7,n{"M.a<>@"+}zW*	c$|;gF6G3a;7xn<\\6*;Kgy;D@+oI:Zek[a4Y>('OsVe+^|}-SO96|dRN$PVyS|XebIL
X#}rWHY)TIqBB}Kl'YhakfNKJ[uiR*yci,*P@b	$is" AntA-Uw-jrFEH}zFgHzX|]k?	bM]iq5rtK-ZP5,L)W<,E]>pC|}y=)&5-]vC J1*](}ci@k|PRec35y0;cf< _Fh|RLZHArQ}lR]G(TjO?v%|uT5ux}wvv^$#J,[]j(QT%4uT:[m!+WW(35@
Y+6oIlaTdAYeC{EOSE6h'ln\Ljv9uJDg:uW
nPps9?wm/eLMi|}=p7X	ftCAKI\e2x6nrLDsO$atqV,pr>	/uD#XJvxallUA-z1+BN&&cZO[}=yBY<.;R+XW}v{>?S4k
s1P5);oAzp:KQ*dx
K@u{Un/S,9j7	FlC=aFhJc5M|)d?[(`},![lUo[-L(f~>TMPKx?v7uj&=`@c\hB`:68DH(%<5']_gSN75
r.aT[Kvnq9^EQ4qs5P5A9;|g1TnBX]=#q/%-ha8v}1}
6lsc&&{97kZ:s.5]_W`jV(H-9]	&r4BhPT%iG6.wzA^{n"$w}g@s5(s0)cb.v.m9	 ["F*En)^XhYz	r My|t+RX:n.OaO$!.mjH5
'0q[kUMz4M=Ei5l/Vkr+?ULt'|+C./??ad`?'u%E{&|ZfyK@}q0qn|FRl{Krp}2lY+QuA+Ov_}uHbeS2ww]1r/nhw?j\1">DSvk2B1P_8@F!E]Tn2oP Zq%~ Kx`
zL@=?PV#:F{DRi
w7?z?gHA)7#4rN5s..".{AjGe{m7;8D-,7:i/<EEsrUxZqFHqwDi35%Kh8CbU)hhJ>*Uz|h:"-!cps#OO9GoRP"0>GB9%0MWUck
iLr 'RmVPO7'DqQlcM3nIE^:OH[qR_OQTaX4mgbZyVRqp)RHA4XM`6<[MQof{d	=V.<6	(daDQ~SLBXf.7[.nog,y4Ol0Na^9Z&-ad5IjzB'H/X`
R8!heL8/=ICY"aMSP<KvgfF3>Z^%.UyBVmf)5`7
}oy+8qBy)MlSqibO_P=$+tXaEO_..@!i|'pcIAAE(-=O|z?W2YE$&"MK.ZTb~zCP<*QsFF>ur12hEL EiAfAgg""WDkd#.sK,gy<A`VDrr"5#[MbtM=76nqKV@Qap7$hD1QGA6WqXfY$I\z2B:'otfPHb!pj4;%u?L]'E,JFZeud60P;Wkx~vvn~N^HA\-;!l1'Lpgf?8`?&9&a%@ib3mE{<8`?%~_4MWJ#ofG>UtdnqnEK5by!i2Yt;%&_oR8^I2&W9e/%|3jwb9?a8QoIDrQQ%NC`~OW0/}F<1-W>"VKGKDL^K,>W#UC,;G	^tiE@,1DXPg4Xx&:Ald%3L8ODL9Ak#gSFQ!iVS7O;_"d_)h-v*YQyKL$d8f-r@(1QqNC\'fRT+*aoVNHB\w8n.zxy]&`+yJH4.9?cu\SsCR}wq$h2Lk-BL4,>_M4U=x*koW+K=NnaD+.>P(!0J	?fpKwH7Y[j?JNX>]KYD8`S[-QX)XQMs5kx_W\O?2y_vc#a}7AP]W3op	Y#.s`Dac3#y6j
z2 x?I	5z1fmhbh)0r2%!=H'
:6$Bg6RH%DJ&7^fhw5R#p>|EX7 D|grluw8%J=1Im:0>%CmiDVHPa"Cf3Y}<P(S75<FH~z_*|T{'@wrrN!&6("m!W(uVyXFfsA89A|XU`M]Z2G)l1M[nW{DZ{:scD-kE\cxh3>UC|vXn6(>~xp@=NZ@82Y4<NF>>F"uI?VT}W^:b2b'|)))%Sc7{'aqAR;4Dff+>q4"VfA]x`7'lA--u0L>/%{:p;aY_lV>.QVL+fzMY#[jA3w?+x"HgF6-93Z@V-Td_Rwe[vHlMI1kW`Cv&<*YKH_A	}8PW0^{QZ<7n>:n5"'S`PV,&2VF
S 7e;ap~zj$xe9Su~^DQ6wYt)xU!L\":@k#tiBbqrk		B	A@;^!i(f=
iS*Ku)OI_#0Sk|,!$fi0l6E#wypKj}P@N"/60;m^u2
QyxQI&5Zo*oR*.r$O5X7TE)?Jcfaa
@w:E!PAo6Az$iSL]&ev/uESd#2T,L[+wLMVH@'gUrN].9LG,+h
XK#,W5&R{C/:%$//_raBB_vn59Q^yUkT*MGe:2
M!iHzoXF47Nh+&Jz!Y^$YI
l(l1HMCL6]gLj<4%"xZizNu$_h8tH4$ggNib
P%dd{zL{?,<ytADt.pY5WR$E6bn*({`#wf
)NC"7wt\p-.Z8Mf^q%fbz@j<^\MIgvBd'0MR.2Q3O!~-B
R`E&b*!/I*?~K//vARy%qC0[.T	;Ezx,EuR>p<FwE8eHh[J\f	z~:}.-MZ!&\t:\&%8YlN\2e=(22W8;4\v4}}dB)fU h5zbxaWt{=wD>=;#lvEQ|vZD?n,W%Di:nN?@8fm"09;jnr5O2]zt!Sm5"ntbG3DgeD<i[kk92o5/z8hRN
/#,Tp'y+M&0ndY;RmzA%9FA96~to-VKDILV,/H{FP>b?4kH2BV:+<G	NnsdWu-51MNTS]GbDnUgNL'Sx:DK#X"gT5f,/5wW7LC7 y<	d
1Y~3<f.@g8xypTL,DyXd;,HEq6?W(YcoUh~UfR<^vvn";|jk2>*Y#Qi.(AX%LcGx_X:nwkYh40yLwlhy%htK_	%/\R.O:i	.t%V|vG]rs!0L}C2#6p#LmOD?md4[D3QXw5n$2l[rTu^3?k;[$DmUJ^*eS
*=aX8_FW?SrT
(u"gj\/p|-4in_V]z6~m^|;&"Ww$'qU6amo+,JUlKE|&^8]n728K"ry<gpM!$yG.+	!?'ZarBOo9r\'OWPrkA_>3?TLp=m#6hmemAG!i`%tYcs6Kz2KPMd^|u\+xu\`Ie~r*`J<DUz.MY,GmQ,K-wtGgC0TR*|sf}70dGS+Ht'w[`@8N6G&vfDM4$Jplsl:X^ocY=zbhu`9OG.1wuuv xGz.H<AU#
y8.i=l}C[tu<	u~x4=^7oIA!tV=?k{_7`RH5P~2@c7+Ie.#v;j?/r;QPhH&[njw6SJ	tN5^e1(!\md&]iB?tn,l}uz{R*`TbagZ$k/p$o$kt#HY7#pcWJ: ]p	@?Ip{*b^tTPYd_vm~_<gq}J#=e#.,'^j@!X1Y.} Y+H7ma!EWC&o-1TJJ1 =S9nH{w+9G]bKI-Di>BmQ*_E;T`un9u	J	>rU8uVW,eS~_6tfKmZjj%*3W+YX/]y<Zu.|O7Rc%QA`lk^|-+e)lF%ebr]r:q?kn7%57iSp8_C0fp82`oxO8YLdE;~ag)`]eyDJ$3[l 3RKA[59Xv>B"(uSpE(@>f>{)${yZgG~x-9rY'Rg7BUS[Hv6&5gaw>?uc8(`77piKjy_yl~;bKk#{{vz/
$	5,/0z<v@"OAWvYLp?6pZNw]["T{]6l9Ul^fx:+A_E'FS{"\;u<^I_{?lwW6lEbhN(Z!s=oV+X"cM).$dz}dw	/0A8'5=`8?0$)xP1)"@}Gl@wr_v}b 7cK%ST""kG9g!8IGq1MV"jSKakeZyRbaboC[s=}n%V{^GfT2sFIKk8f@Q|tZvheE^7^&;\L+UP'x9lo	HBG PgxyBl~	KhzJmht.|Ix`C;H"AONFtQ0CJW!qK@e'*t=>xU|d-<<R|>*Y3ZYT["my=5%SxWZxIzX*dmz	>i(qAv7w(IHB]5mVXhmVAR_9L%P+4rK
[ga0U2HjYLT{>3`<Fq7`{Q&9AJk>Z*S3\MF_[Hh+IzIWGji
=F[Suu7}Me`xg6J^1iOaGC7DDRqJXj0iM7I":/Nc )yJ !:r0/RPwMhF\rBJmQJ8Zz#$@rCZY	U4O7(IzmjggFNp>7qW1Hv"IVq3t3afpE
2g)%DZR?UW7C(QN?#(_sd2+Oi=bGc/M/9>4kTxV^M")FOjpsam`jq6F}9	/G	+H[P/`pKr/Q>wMk}gh=eDz"z73#+$znC3FoAft78OtVo;-^Ic+;0ea:O8x4<: ,OL5M[dM.*!SDl20JK$G4~AgK44E%ZR|#VSEXrl6(BmiU,yc7hO8b,yMKBz~(!1xNy?aS'5x_/4*atpzxC?WeLESv9Ko3ENpL\0(!7{g1K`8=/qvYCxU{,+'-lpc&pLP]0(
y<lhvC)$`'hYr?HTsE>\|T{Y+0hJ;h;Q.L,WVA)I\9bZE8nS\d~Y!g(xrE7{@!1wcDy4^\w-	dv,M_R&IOf&]Z0bF$uRv]^X8m'C7XyGQ2-X,Ubk?G9k;1=-z<Opx"S|c~U<&U]KR1XX\^Zd'0IqWE$fRp^QfTD)< E*OewWkc~Hq.\CP$I^9EYJZ5f!^'Kp!\Z(1fb.?C!.Q$SJ i728;_<:K{'Jdn81<	Qe]S	5.vXBz0%
7DA*e*])W@VC0KDhv&]|CsB'nG79mAzE3yYP@4 m}h3C*z?3("/NP+e%F
^Mblvg):@N	3`G(,NxjYb
A'Sf~9]ly].d06`B?a6Sz(,$!(ixf@gZC*ySn )ccar$Q|-d	bt$N1s$;e=kW;j[ta_$t>?
)h2{!#H6,=kSx=l9E^#bl#Bb}Lz\81/9]VT;T2@'5LM%M}MN]]c5UM%7 1cE.*9:lAdYPhTsQKpAG5^0Iu@A901qPVI$]88/LBp^4-nLu%A#~J^vq}p$yE)Qtl8oh9IfVi&=q4^7.>Q\XPX(_dDVEfMO?QMc$guF-7i$eQG*)?t,&2N]CIBtn0ig@s@%6dYS8!AJiHPfa\;<)[!OL%YBg,)]7z9YOr$Ly>pA"%l_o@PhKoULu -=JqjfISS5V-kU67P|{%3=n`(tJ91= WtX{>D`ouL52A:Xxg&2B	Yr'gZXdCyFOs/ewUc'6<.g6hMi1xbuNKu}CUzL-79~[{0AU'NGQ1EA)Ok0]?P#I9qQp~)C5iKds{IJ|qL8[h22I52}k<60!VUJgF0wk#1E`a&4O`H b&'bGqT[>/`^wS!nYP^auQE|J|<8R7k(r)W{|y=q}]r;-?Q;?,*\O5Z=/mU953{XYU./tsj.qZ1Pj=$3MIxA@vU&/+7F~|5X0\.C|#O,i)z..3D(Oj91y4=-M]^Q@,jtX)bGi	#z7+m
q0S\{%U,gqcJ.JlW&y5,b?mU-RIM}.e
C.t^Ml^*'ByI#f:Z\"3NkgcS-R1%&(|?t3l>>l|fwOA?C[=f?U+0l/nFpi>)0o-'uVf>Z)[
yGLOV/"Zuhq"ZUH{|IkPKw]cz[^z"] 2Aj0i`IW)0pd:b{q~CgUD}WM~U}(;6pozL~K9BCPE0mS_oqI8uwov)fL]_s5oJB6:OQ] z jR3h+B]'$-R;oL{	
}kc%mP6|7)>&1HQ('Wo=HTcf#z\jdWV>`0
]$_pg6B6\dn|f!Yh\1P
"B%D)(,p[6Sh~/2<0J=,{J[[\Q=B19kP3CyRJvxQ
%fR)pl#35KvFV/l&bkT!C:0ut(.DnH\JD8Y[(_7S@9W
y+*HIR/WS4=E[Bex:bp<-\noJ#`*
leLi"5&(on;T$tWrdn6F4m#`.j@$b"[p9&=|S{'9FKd@!5yH&q;b=U4t@S6j0-DL3Om+NTZDtP
4(Uj4oHT9C|u7?w1j:Q!^.)_2pi'j|urX1sb9@,XBIlK5rmIP'1E+eh
;3;H<=NZqwV`71W/HJ7_L)VLie'WhW]6#x}7y* iZ96&n;)m\eai=!aO
kti4AT9dp9$i,$jff7`-S+vm'}]84)~isYN7E= jWw5c*h@=/yk::U'.AS)?K|/v-2"vQGXj;nZip.|7~"%sy=^+-E[hrW&o0f_k{4hf&5R^s+5AHITcdSRke_i))`z"eFMs:X]Q(sYQCOR;l+9b{[&v/K,G&$8`!@YPulfqQY*ej8kQJn
(9ce4!h&noxE=J4kn#<^}
{JnPoC-L7yhr8`wk~ch2I-1ZsYZK3QB.c$Hy!=J#U#&o>,%.TT.W,^eC<McZ:E<)kx1HxbcF2\0PqCf4`'\s'}x%\J9|=/\2`aQ/wPNAR&o/$eNs,EwyM81zs+J6.NSn@dt*,x=9\fvA%y8F%*JIZDPO;Q Y^hL.2D<^?{=#CE2aTvZ,q0@?c>?$V!QyRP8\	K*0o,Zz-<8q%9^EmCAGjsJuGw*6+jcBUqp?HE/K>/elXo&q?\P7N@tVQ~T\3p`ZQtk2ji2LMo_\h@,ut`<d7r+zox k!A;Zw|#\h#wk*3r6]'1BmeTOS/`2s,\MN>K[Nf1	}}yjJ	xfxzVFh^{\{B+Z^cBf.}hb"k$f	[u2&qZM,>lz wTZ?CIx58]$d[s+nTpth+1y)}=*2]/1u~\9GiAp
lh5-%]J p;<zT@ad:R.?v\9__b7IU[bKQ"L<Xe@+nv0|/7uJ@l=`fvtp,UR^l5v)^o0U`,\k.%2Ij"[Q"8m%&C?k&Tnyc|S># =;jP]_,l06TwN)Rcp;\~-.HJ!d$DDW<u3R$rKMe_./OomC~?KE#?G;gV$&JZv*@u+&'fz7QZngGVL8I\=(gIx,a-5ImjIhL2P%=,(Mt7XM]*F.%
iD\;\tjx[V" kc8l
7`CB`#YT[s@u/zQ|mqz8EIAEou%A0aF.b[$RI/S3x0{AJe`\g'm{l-Wwd4q4NSt"h8;LM-jpp&(K,\Zz<?[F+=H8
C|^{Yw}J#4qBuN=	N#t9xc7yRh2%RuOb'	)|leH%^v3WEc3'o1h#v%cT]76XEL*OL}^)#eMB_09q$uL
|4x\-SX>*tb`6K-z&b1%
+>-4b&.6.8gR,76O4HxHep>^/=;#[mSGYNhJjYAam(j7sl`R~NPJLg<yH#o`1$/BiF8[)9I1xka{L;Y|6"N:3?a,*i(`dR^^PimFsW/?DTe$@h7HS#-D^0'G=,>mdX7}<)=i(pR%y*qlS,rr>@JMV$
wRa2&MI7cI;YlhP\ZoG5rB9o*Eb^8H%1p.e(@QJ2*	&#z49fW%chFclH5S#^4D56HoD?G!Avm"]R:<v-_?c =qh>*l=:[)|gnkRhR3f7Ig@C_Y;'T"O{Q2<SKljS*v3:?
Fp=.`	ZVicH1b<sjH^+%UpdbTbj^tznX^VNlO4zet"2+"%.+(b)1Q} FDuO77n,;b=nbM%VYgGl
r/3^oL93*(u<?Z6&[C)wG1J.$f5+'qAi]3Kc1 Uqfv<<0AKW*NC%s	{}DJslA3<]b8{9/7c1L`wa-%MI"bHkf6#5kP(G0.AX'wm!AwCHrD!pY75>Q$^mpUccBTL2^X'mkRYh~A8TkEU!3c:R 8MmdX?Di'HiTW}@#&	`5zULX.<zT)74Y{~|"PQma1$pqfC*asbFfkHxtS|3B5*p	CCzG\fW:pU6q_uh=!{CubG<aMj+e0bzXd+[jm1tV)?/[2"Uvv~9@]Ii
p|6AS!1%sqny6*[B7yh_A`Qv~s#orOc#ghsak1GX.BTe	[;0@Au+C\.bt
6*Tzj)!>B1@dp+/|Ya1i;7n-waJpGouriwl`>)cKakD94?^?%D;{HK(I(r"NkklY`#@H*9FW#A!)pf99`u8F~{Ukk_t~&S`ZazkrSf7PC8\w}Mz!h+3/n}68G^6lx$AoFz0)?^A(GOSY.-Qi*QL*S)#tv87<tcZBXB;W<tV C466?s.WyUo71DaS6Cl]
l2}\g,wj8NN3GN$,6JL	gSjvCtSJupMOT)3OYC2-`.Z*h.NC77+=<"#c&,|i<VMI8|ottUnFR.OvyjH8K1ytU!sHF*%ZD.Do&mX]2\ouE&4hK"P4$dA]&#HVSbR_.H+3`mI/foU7a6[`UbOb.pcT,e"e57gt#{F*nZ.$THn3Wv_\UoFq.>`xm/%K"U9uSY75e7?=Gh7t-4#7J{5)xa_e[QTD9|_Y8v{<SnL)E)"i>Z
IWvX$I;T|lT"f6zxsd-s)0'm+odA@%R'n)IN]9^X%2|bT0Yp*i&CM8yX(I%'qG@[E?ty\DC?z@_%9,T}"\n:3MA_}_")htC2,DT^f51ENKF#20i,`mi2=.UPgfB,&VI}eaVp4sMt/%kB%k"e	 BU(=z^Q%*9_NRXdlQRe60{I}eV:VE3%C,3QLUPYoz9+'^#8uk@V(%]^OuL1N&Qq9bQdQ*=	1E%j
O4l0rS&j@I(-zIS.Ka0\Xhzn6RNjZk,ZRQ7o^g~$h&	=^1y	O>?78	3I$Ir=#Gb7?xDT9?K$(H]?S}Y/*W<LVT/G(#SBBt~&T\"S$]+%>SHjR1SOdb}av\fGj17fFV`E
o
F6'4>d{J2:rr2pC7Z.D1;/CSIL7TIjyipA^R%M1KM4_.Ww?"LO4~+[DHpfmqc.ffhV1?Y .!.[TJMrw Y qsNzB#rFhv*eFoQ tL_,jPT<zJ''B!M+/UtM]YbxE=KPJk7<%Y]b1182:):(5$l9oz67+pBE6A)V/z@ifg81)">'m`F8|e,i3]J{^
Z)V2QH$ts\dbWe%1B6p5!gA6~CO~!_GT6t[kL=&uo"j:*p-@1`y%YKGn_S%uAz1wPX!PdQ1|{.+Z9j(bt*	9=!D5f^G"L4ta=YT8[(fRi`Er0Ur!fj@Q:#5qr6:"<SoM(6If0@).tLwG1IG!B%s}JzjAYJNoj"4aHFnjo`fXNM'w(N<j%"J,QIzZ%Rt	g]l0w>z_&lJo\%Vi!JFKfe|0WsM")<}>q#-GAFcy:ihOO_:$#PR2?w4:}ul:P
z&,u
f<b1bSvMF+}U}.j%s).`.fh>qo20v@g*!7
L)B dA	!<FAYjB/lmEppg!?M9XZ<}u}4'HS~4oR%8EFy=HaPl0Re]"z\Yj./6-Fdxg\/Z
Lklasd-LyvY2qb]BeN_ywk98C6Lc8@/Rjdr#.Pmi4Ma.g4`Q
	tI{Vgs	<b~|d\5;9EUrk_
Z`9Q^Erj\]-E{|.5:q]4hU$>1:K)5]aFlmNs)1g@)]rE)ojD;hLUjZ<X	phe>([v-;h#_YY?]?CHFPRXW'N.L\_Nc<E-e%3Na*5u(2Sppks<mB&e5	l20Q o]#w(>&\X3BJW^2R$s=058G"CJvZH,9vNd-hGP|	 [+`y61Dg4haX"JL=vNA&^QO{o"ZLcgzU:#F)l2$oT$sqPV_}50TJ+NG"1q?<,:LS?9!!Sa\;Ke']1|;%pYK(<pZUSr&Tlj9vB3`R+8Ob*i?7444TPDrs(ij0%*@Qx'04yTfb}16T+_	rl):M*y}nzI[}e==?-2*;E,/\K.Qbcp#jth.P5nN`wR{JHXR~6Kdh(@TsvHX[NjJ	v/B;taD#s/ia3P/3TL#>r%iCBE+\1[Pf&3jy)8<i]+Rb$0EjYh3gbQpsT~(u!d}=XyOZxHeH#oArZS5?~@:w$v},PO	v>L	Q<{MQ<*l|7 8z^jx3g(*Tz;tYF;3peRw_D{T%?>9Qwx%GXsA6^UMy56|lOIi:@Q74Wz4/iA*~no~TBe~b+jhjw66M]E|m{2-:%v5'7
G+69{)"7]-2%
h4 ,z,.1>g`o	,.X.wbgj){L^rqM:6yWG`XYbEcSWeEaqlsvUBhdC!`~4Eq;1`c&?Nw#Rk"]n'$!C;M.mTb6o&y{*Mv8eL2v(va|'6A[toecu<pW1BMquQxx,g8N19!!cE3PJ/]kfqM7Z9#_h^eT0",`5F,Kns*u
*UjUX8aG%y?w=#%awYsqsoV0j)}{1{;[!z>)2IMKXEZ5(=t&"P\CL*uh1mVC=21NuBPio=wLf,Xl"`GR-EAcrD8D#"@Z[I1>wg"S[K75Gyb/%%N\JFs#/?*#<2P8kaX; 3=VR3n)*.0':CB//euHS-Kg/P/T[< cnuAA^nevbTW7 !@p%
lk=V1B)V[b=e+3$1QSI&^7XT	HXYNBcu&D(0E5-	Qu[MS$*1GImbW(v i0~?|a&,
s#TtNc]@0up*"2MsASj{fUr.;*&Kis;V*K`&(8
Z+d4E|X<j{3{HrIps8)MW]7SWqp`8}	oT$q#Yjs\~.tLV60I7Z%9U[ IDSvgCLCK:}gq9N5%@|+}i)wiYdoJ_G	0\>i"`uN78p>Xnes7jD$?7Jd35PBX1b1%d3+pMD"ZLyBar]JOH~\
Z:{_)>*:tc1H
]j5c0F"NrGJ+_<v:vlq(ty|$Kzp	o`e7!bk(4\dQOFS|aosVRiUDJ{Au#`g@a1{Wz`ir'w'8M{[Bg0P	R
RC@0.-Fn'mtHpI1Nbs`T{LW%		K0T<mt\%L&yatnb-ATR%/foQbU%^%#TLO4v@i_l8{2ENtQnSkbE_%B&3!bU~phk"	aAYiW0
eNNW[(birmJABBx9AeVKIE]f+B!zj*hX8R|Nc]zzuEdHSygIJbeF&q"y0[HULWl~cq\F|q**"NTd@].3L 6:v.c3{/+u#w+3%a<c`*PGto@*1E-~?br>	:-g0'.3)<~xRdoa,m|d!w(1-> K|8m4`*O	KsbOzk!M8[;,++X9qqV/b?6w;'?DiL+JFvQZ[&}Z3FfdsDr_t!?NiqqFk
yM!MI\Ft
c#R56EUe]&dJQYJsW(0'QesQ(**vg{6xDH>b-
MSoVR~f}CXq(Ns+k6'+P|U1cC"/H!F3:U{f":=STf7`7Q/\I%5y#k+x/+)e.gPHG.
,*,[+q[3]BUV4N;}z2z_%G1LYbUZRb$r%hfIr`-7JY%'|]<^(0^-h\\B/TnU^"um
Ve-gE#puBU`~>4M},/s3UtV%2mx CZQ*TS0tsDU}v+RRaDrlz)lpB_vZu=wvtJVE6[9Xy%%Raye^|6|\.>tI@HB~Qth{caty17OE$6JBnWz<R)Se r?B5r}aGz
u{ZZ5p2GZ!?.@_N]<QyS,CDKt~t/dI#\1[`az%M00^DGOa/Z
o3{fjBk,f=QBf;dS4dIB#K|,E\3<FrxD3mtmj&1R/9J.R!pR3'{hz*>Us[_%T_uvB$
^\	"pRx2)c`l{aH(4m!A?<KLeNv!t)R\D!bh%'Lz`f0\HC?db-4&=sIZ\,T[{jrFFb~!7LT/6v?A\95c!D& kE)U	HgTosI'2"	UK?nL2H8H3fKIgXr5jq^D!DZwj@8f Xm}W,.YRE>
mK=,B_K1_"/r9L
F}:qvgA*&(e\fp\v*D
.!YW{rpYheq[Z]EyY>C*7uf~J	
);2-D$H3~>'2SW\q@C}N068c?V@?>hd|:qq}yZnBvz/ch'5Uc[&ZO0H)tR]t.#	TdFLc=fNR.i8n	TKe#|w9lv?0'|;	`FPnI$My%h-c^m\\x=.J(e	73tF?{aTl?NAiGG#t5g+}N4pk={
^KI[,M1;|SuYfxByH4U8x[C5<!cF@KuFl\v0QR-x.pkE+<%!=2+6f/-T]zdR34RcO|Yqs;Bwmc'-E/Q+AXMxPQE1[Ss2bV=8,9L2&yQUCyVS'DO7M~,'`Km/%n	sDgB[\&Ngg_D{")D2|iAtD: ;WKyxMGRE[JOe<-KYPJPnipR&7b,/?ly}kj!-?;(Lai'unv.9Xol;7A%	Jfy-2TkJs];"X
!Ba4=4d2M%	K*YQCoTiUB?DM3:?c4fN-@,lc~f"sd4xB !TL2bDc$
fU6}4!^'@ovF]{&#>Y*sR!/?rKydiX|hBS2-
	^
^M
/b=<;):2JikX,yN5:X1;r/rsrE8}	-yHhv#2d[2{COw{4G.?,fJhgJ)Q39&Rg/ Z|Z'(;880C'Spb(8xf6_z*gM2p'}$hKeD<!S$8CCTbkM]Si"r@!3Q-tZM.6+(V"cVZ,PL7y?zPEgI(,[&E/oR[k5 v_/m#"|+.u08F[gB'y6f~6C&e2o1T6,<D2l{wnZuM|RKp|Y
#r*rt*[<KhxI]2a/gc<&u	A`sqZD^!BM &uho{.Qy_;	Z{H6s?*>)i%?\;:>AD'aUb|R6MY.xO,k"/6gn|!j#>w9nPIq}<e,XJQiM3#wJy_TFv#`S6K"~dBIhy>'89a'ccS)E;*V`a/`d#&^u}'L(1XUipI,y?OM@3!MXc	APj>H=qHXwxYixm(4"133]o/wK1LE<4C<i_`t<N"3G5e%aAU0HA*5K$lv
%d!OBTuG(dwy>p{
56Q ZK0D"1l8}c-V4tOczdY'aGbr3b0=8J&o2@?{`sr/^I(L5^Yk:!Xf)G~%mpd%1uK#/sZpgW>dTf	G7t.{L3Qe,Nm%0X&w$"u-$=%;b7*V>TM_VaL;XO<]s>=GqL$qO0f#m
Sir@G&@YEy#.sJ<	{4a%Y\6z0WK?	{@3]8Pdl(0	|Gj:f+K\?:cy
Itu)+f@@a+\]_r;v5frCSI2fSpgZ,B6{g@{X{:*zYe	9c\5-&|&4_'%A|/;ktL 2rk{FO=4cQh5	LA);{2S"@"p|78s	O+y2WVi`Bp:H9D8CBNj"4Rs@N:r=]Y^7MTUB9(<~i!{?evD1[R~(_HIDX,=m\%cg[BJx>=8qp6wb~vX127I.pJ:=K^[Uzhk/Ov~EA2YOm:Z3?#@`pWwL8@KLh4t
_wSc)zbv`cSqB|a]!Pi8dOG=#=T(&fi{]3Zd[m}<E;:4Y`_Y:EvBcr:hCmmO~ivZX}b}_C&#_-O9x"@gu_ v9zdM0*+D:A!j,uW7vbi%w!!7-vth%O19{/~]4Zs_/<[ZWc&:iM .	xUR$/*w(V-^br1Q]+aCgrX BEgLO5NQ4%uwlGdl%XoJK^vg-e=pjbHqn!4O9d\hu>d<0mEHro.Yjj5Z8M+';m%cyo>|G-*%gW-0P})'=X Zl)|Dqy6?Xv|t%2$T4Xf\]t+,B!\u^0O"|A1Q)3U5ppNf^6:^!&1MWf7[n.]G]k(d2nn<]_Pxsm23igg'i/=_!K@0{2K	)EsWLO=Wj%m/&|BXAj{TJkxh/noW$_}d][p*"*<\F9-V:DUVK	,&/<]nThwVsR91S8:t)R#wPM~>C y|4 ,+#$Uf@c,`_ez!zxl\)I=n1ePlSS*|!4[v'>a:SZ~IwIA"Z/&vVTb6I g:J+'Ph2ph6/RrpNZ<G]Ar=o r\8jbK-oXi;66I);]:1m|C#,QXi}ce:&r-EnoZ GMm!F?!564yNBj_\r#Q$]dHUE%0KZhX[Sbly]~8'x@CFxBk;q0H;q230H#DukcrnVA%epO9_/+xI6i>@ZFzk=>RPW
NKI0'Zi%\?.:$S$1kdAwpFr~0Jyie~+tX\^E[L[s+VAC1@{j2"iZ	*&kVJc~N	I$1X<BI)JDa/{v}IYO7:!R/(hM@&&@Fjs-9y{J5d{'tj&Dc(g'UMk^,vL#W%r$=4&rd{lbX]pnA:0)TBK[VHP#c= t,)u>">=i~GN"+C!: <3Q`?"	RZ0EZU#<E,'7IfHLzw?EWT#EE,B\e5On=8@eFmk<ZWcF.#PCXpML#ZM5FvE;&ga)GxGEckE 5~M.h>)]F}_G0>vY6]km-+z@3j!I1HA,"ZMZ:3)b&M<>"d/%xHj3s4V3%9.;Wmss{+x{+oU-dt[y#1444!!Zv2Ng4T`F.LKSR&g#V	"u`{sI][G47jBt\0j@Fn[Cusm&1I<dU8@bm
Qq_wj'y&taFLh6@;hV:@GY{X.K_(RB,TlyUkuaG%SX]2Cv@4yRC"??]g2)\Io[pq>wCPL}jN2"{#AAV2@&p>l=a,5z\4(\"Xrt/EsEv4~(P&sl>t7,x2zKXuX`94o4
J)F"zaS5,77C8yiH~<}DF7sS4i/Uo\	D}(eq	C%?0ggYh*lMLj._0G|nF]m0Z}xLgyaQ>{tslnJCu-yZ		)5?B|=z|'ahcZ!"tv{@1pd!$	R5_CG#g@(y*19	_	.ceGn3IUv
bZ`mr||phJzxTosnYGj:O$d&VN\sl^$1{8_&n8}C[pr]HZryXgK{EmD7H"l*ghiE.?TSLV)NeMdSi]}vS^m2l#^@(]1934gw}@SQ|J<)5DYlE~j 3KU*?'/+: B5J2+)pYe	L,Zx2piEx/{**T5uQq!S"O+"wknr&Z3lS*aqPz2Dr91B\=\8MSEX{;MK{ZjY8EKl~k[Rf5egw<".MmSYI3Lxrm>}VnXbXqMGB6}RyFObw+T@J\lK $h@	i`0ppPUCMv;^2-@&^M's+eoEaHot>ey*qJUSqBTuv=;dFwWNh&q^W*"FBga51QIw4?@dg{bHnh[:gL8B4 iM06PF8^"0;.2s,-wY1;v Jj!`Xn-?<3*VH>Y#+Vg9#_AU`eGw[r|	:PgAFNb	fq,ff{LWJ6a>2|Lo[ig"b!^Z(R:6>Zi]el-JNzSe94Bodb$8"~
cAM83gy:FBG|Btwwdk)$(S&;UMEE#w]WK[WL D+gM@G
KAv9HQiH?}if2CSsT!_vi3VK*5,U>gD:Q<H%+}7YFa5AV5~45@,5t6H%UY2#l
$f;@o^iLT~tZvhs'j2R3e-L'd]@hJ[^#d'w-IB\`hC	|>h.8/?jm@stT5|![cT=$J*>XYw!>;7Ud#{?Je|tR$II:;ga@gQ1k%6tbj-/AArAgX)<qQ#r)vjau'q\yg4?&W"@ SO/a7Yej\gTyLtl\0B>XdxdF:3K"gs0v;al<]ARyEWAd.Z~:lCa0P|Ub,5	JsKb#~glc)3tW*PH:<6H"Ryw<[4%z$by5k8qjdPd.}H@<r$*H#zrIzR[+-dQ/')5wCpsf9ZA!iBC>*at@^m}\'M5l)PO(h%,x$Nw9(Q[Cakq.r4%-2S0K/ucHk@-5WwBLld$N|4{#bqFrS&
	OXK=U\Y]Y=:rH9Km`S\qcd'z"51dvpCaISnlvY9DqckEEg2E!}!@ufKi:;n,,N[?W+WM@y^;O0P}v:uST^9wl3/vmiX
qY *%f<3TWhEP|0dnpeGb@87DrEBd}^1?k;!d(qpt1dE6Mo7wX^=	u$VE+s.GB7Z'A\i\]0hIoy~'gE^u Y
h5JW'H%F\&7DFel;#pdD,rs2,PYGnfs6w	8CDJsMtyI~?C-:nd

K#4i{u#*7[K:#kgwMc:?Q$lM':h$GdBf0K7,DL9R	I$3}uf>)"Ld:$s(	#]P8w\{;Z2{Y9DwAFa@jP|A\oHu]z]T5XwOwv)
TPSsxFh9,]k:7N<g-Oz6OD_veQN3pT@u9#WY[6m'k24rd?|q;ibj9z7g5%8T/Vz#Nv]o?4oNlboboB.3^faktV ~a{e#T>W)P-F,U0g)28><RXph_5W{6)w)(9\?-ry`]`&UYL!fel>;U&?Akt%zkn8]@p`F^+\L5SL;Cu@wcX$lr+:.7d&WTvmbHhHhT
UwPBO6gpc$q?Rp@#K+1KBfELo,l{=p64PZ0-a}y	Idv^Qj8<>%e=0Z,SdMFa`u_P
mtr)r,6n$ :h6fO<k,!* 6&x>a|wM2Jwo>QLR/s/
sm!}|tt~TJyW9{Ki/|cH[g`g@qjd`p?DYRPi0xh%ek^uY4{|%v	ZYU-~bJ0.(qpam}aX4'rz?CMfr y,tl6*R^ s cbe!,5EAGKEX)w|Sqe{ <|\dQ19O"EjDEV+WiKI^lB>IElj1avUCd{M06Nr:S0ri,w+1mCNAC:"]M+jWIC(v)) yr
?@%U(DM/6L{[ZD5#HI0XzAjA`8cAC,ccHR`B)9=^ZvcL^K~%$19bqe[%E/eif^+6!@bzx&sKI@KE8fev&=i'$j
Zs~OzMsVOf>6q9Vj,i~cCPNe}?/RW[1 N8@y2=K7~eQBdO}
h2$l)ja9N3>=H<.U=p)^n#>g0PfKs6?'&6jN~P6NQ
ivSwLk|\"9l,x:rB6Fl V@ahLMHevQZn(X!m@%VHo\aY:7IVZMB
	]+.Fb"Gp:irLl\Ck-fD.ZRt4b?B`P:'XBS`;|W9|,S-}+IXS8&BbC[l+a;S]]}:*MlU;R@H4FK~*dQ;MYCQs'T`m}dU'`wY29-+~71Zaug)rlPrr\5|<_'Se]\tF?H1e6n2ZJ#-~X%>~O"=#-0FzTYzK_j']%!DG*m.0*G.:(pzG!dWmmdk~IU)R-ihy+m;^pDuT51j!iZJ4}ykS;C8ZWk$?#8r!dFA
3'\[+SFPq "9yTk]Z
`N6y0!.<NiGltgTNB/iTZP8;*Ue,$'BKT.BGKFb`0)K?h\wvm:vj<}'wj%'*oT5J0Gu9CpI6L0Y%KZzO>{uR<..lN$yQH9jGW|#n'p[H6U6Y-c0Oc\bYUV>sq6jD+@D<<%/LguQTCB5eE&p=eo<@
Zmr8$E54KMB?|x^9P}3!'9W{O'eTFqa%:&	+e_/DkN" 9Y!+IYOg,p],nDr5.fy^XsweNM\'="1Ra{496o=3\_0{m@jWEFs9qS4lU.]pf~+m?IKqnX4'xgMZ{tT:uPU<<Dbz_konVJtP1I.j`ZjL=U_*>#k`f9+C-nE8LIgi88L5Da%I[pU<}m1f)m;O(J]<+\x'F3a9#f9QR]Kx&*iu`SSY/	?=I^jl{v`W"[iiyik6NdpW$"a9
?  3P^NPxuipc)MvILrOQ\rAPM-!$@:&5yKg]l?
N^0RKbz2a(`)LfO3
cEf:~^Jli`F9M;_DCgrO`+4<;]3G2 pC7ztNFPS7zHB5hSo8+L&qp\T6$Fe/aS^rj-pBIwngjJ:#((nLEmZ}YNlU5u)BTiP(T/{J\4'&JYu1`0^e|p.M"Vd}3wR&p:io:1<"j7	&Ys2_X0Tdz:}3=bgokNe6
,	=!;2TQ|&]ipSQU"H-2u`'r.ypu/Vtb4M}rF=6C/5VXUq0;O^A9i!JFhoiO$R|
-=Wp52W=s%~u;>}uI"_JS\go[k!%+P,2zvG]=MP.`f$*J*gg{P_^3+kAnoY3[A|T9@P,vPG5u2zx_G(~]<X-~x-k>76jw<'
a,*o2Q4
9`&;0VghI[>(Jcr]zx[Y`[@|;e40vL-LDdo|h9^?<6h;dnFZ=CJN`Z0'~tA)-&#lNE!pnfmj9'9y[MC[CoBl!I9r}is=/_agwVSeEZ\5
#o4K53UI_'	KvJ[9CrnjRXj0,|GV <F`u\@%.Q{OInl^YMAJ_{7^#/=R2HT'y076CmCeAOWyHW]Cco)F	EXsZq]|f ^Z3M
dU?'.wF)y$G
:RR{W(m^`Vwm20xJ,i?:[9lc(H/AzCff2I}.DdK|-ywVi^r
u?se\_re]$%;3bLDCSXZ\|x2Y5!?*i"Q~4G+dum	;hs Z$RB u#CAFKw]*UbKibCUwprnVTFoYm8|)z5P3y5jy f84%rmo\Fv&z-Se0#+p%ZS'6P"0(VSh8Dn?vQp9V
e/CxVvv$@)Poyn,B,zX~9)F?,--Bk"KS,NUt>xEkf-lCET9T/B7{V(uXzAQn11o#`kr+M:0oHn:)]>"s>}({ jrTBki#8Qv4|:)zgARW%ba#K) xiiuNiGxFr]ck[Pi8k,,95ASXxtZimze~kT6>0B(%4JW@tkG}:
/	[_Nyd=Bh/
>RsURM$z_iS`|L
"dvsls m>]]k g0V>NA
PB
G73	PkaQ<Qp[2-\N.N 8u
|6S6\Cyete6QoNfG'0,Uo;cs"3n.NQ'A)=>-OpjS[1z[G?BJ#[Wz&.'C~5,	i:mHm2h{f;V^jsy=%|_.Pd^79	b~8v\#di:Z:^}O4=<Lvi[T<pIqMjR;!E"Xjk;<p`\L&Ye{GqPx-I+N[q[:K*rX( @0hy(kc4?1&O}2MbTvw!S6JrpLu)_Z&o8YM@wwaJ3n!}~+EnbG )	3JqL-/`#NI+MYrplhenmBoH#1o6|E${uX(+7HS%(v18si}U,}:pVR$Vf{+gj[ebna]c#8=a
7fe$b=^@l,<zpzP@Q*Lvp~kFeo`l:6eD=*1JFQ)KbJMv]:X*Box=.zIJ;acEniW%k\GH'O+n+pbUeSc8L94/\fNcMQ6B=eH+Arv!|s0D6e<i+O:YOqsAkm8<C@;UPh,8ECh*rgB7Rk^m.c}5`DszVg>*RD]Vqg]*j9\ y7
A107QRfg~9rm}kg,_q ja+!v
Lnos1i*9nd9Hm?Sk]=1_/zu^W@}/+YdyA7SD]G<pqi&;(me\Zp5HT^,AL%LTJ$9-dNE8}AN2FR5W1IJ$Hl1Lnn9|(YIE}8HK7|D0j~Q(%xO&/MWH7|<9|&Le`(Ms8T5+Enq
xoS6"L1
K_ZrKG@V$Z6QL :tx`J-"hiB{4B4o.P&523!Wn`l>fC
peJm[1>P'+>ui7bi4CFexr+2Q[C}a\i-n("OZSb%[[
_p]3yI[feE2TX gOKIcCK;5C7i(6,EHXA'Mf	EnU9hC0V1V;_ J)e>&'n0Vh4Rd7y tlwJs@O+CA"56(o=(nrwuhhD\W=e6>K&A1DZm0*@)qW'zF*rj7t`(0)AnLMH3yeqc,6h/8@U@kOmVJ{S~t"sN>LO.mE.<I]%Yl_0sOrNAl0^.yXdZ_IoIb/XfpaqD#OM]"dCdr" |g=.I;SD23Bk+=hrE4D1Dg(y65K8Q#M}gOcwpF@*hKPMKexGQQ{AU1Vj/M9OwMXWrc/nosTyBe(JQ*FKLUx+CC*o,dhK3{mym[Mq(Rl.zi!zr6FLN{ YC'?V%
phgGT*kPDl9oBgMI`[9@"vz.*!OoYF{,'beL 38O"P3+O[l?Wdf^6[z2/-a$Gf(g}}j><Hb|QEaYJ%yMW1/X@a}P#jZ#fM$6IF"RVjl[$6k0;D{X`m.,tmv.U[&1&8CR)kR&;6:|RL?/C\p^@_3!y!W:N6y
YPoWz6v]pX9=$CAy7Z(w\yY3n
IrYF/-|6B2,/U	a0cEKda8,]3C8KZ~yxeZ1|JA*FxSHil~CxxRH.7X-*RR"aGn8%==L\FaXG]fE+~'Wsai2O)Gw/G/zQ>TGO44.Vx\';vS3sCh2}L;l#t3Tg'sRw?kf^j>A_ r-P$OQiRIbSeA?~	6>x>@DRERj$_u2|"B49Z|etz+H~CJHXCn*bi*az&T'Ra%0?	n!@z*nNF}K*<5Eh;lKZ9roOC@&^BKZSk|C0'?t6l/_dmUM-p!JpV@?%yBE@Az}TKN5SZ;"Z!|:g0Yms*sY*U)qFXCMs<hyi?[;%rkS8j8{G;`MNFN,vEwL /3o<,t`:C6Xj>RI8&cszj!\^e`:k_gMq@\	jeft?Nc|.}W;/"Gr9,:{O1Bz]rnkY\N x1qMJml[;ktg,PZ;bt^7Wb,b0O|50r7`RdIJ^u)^<<C?LV{Q,8Htc(7&4`JfvlVEIS 0;7n	e'$Tsqm}:G\${M(RDz-\K|?x%5j}B)^@Y =x+UPk$Z[F}m|8/NHC;0SG$VdyB+Hi9jH`JHB#)`PMHO%	}Y*n\eSf;-*aaW.]9&y2W<t"o6AAf|~<|8v	Mk|aa*|I	9=:`Rn2]5}3)FQHB09xQ=$Yp~&:.jmI$Ug7z
81$D}0nbtk.RL*G2D&\#)Pzim>(1	F.n6V()[KejxCs^E!>(WK] +rgMQc(?Si-AZfe+bGtuPsl!xet0iMQgWk^9$]JiIH4 eDYDgr2}:KUl5T8!PL:\kYL|5C*W),x 9IX?<J*b&O',RRI^4PbJ4chYr3y]Uv>S~
/#m$rTaeI_3bM`cV8j~kOBQYguUTv~?ree5ec_@)jcL]&]T5h1SEv/^)QpnrEQ/!r6=`uvq{aKX(	^n7pY{$+!"RY0Z{YBfT|(r4E9X9FFGRA	8fOjz7"W*(!&NV(i)Y4%!RG$_iCh|I{Zr.cGIhzuusqgSH:WA=vQvL %4LARur]<x){7nzK|B3JJmt`D"LUju4D;
ZoQG22:S79[n33w:=y5@80I?P'xh.~-%Q+MZ:OCA?mQpO?M6
rJ|4"#/bx
#1 W[(Ty0vS}TXo91~Yc
L@k.a$rfi :Mv[VR)Lu-a"_I xhF+X$4JASa_X$zO<Qx3FQs=K8*1h,c7sstQlAxcIfDJ&jE/GkL]\6rFSv/d&.pyd(;~^O-v1P{jk*l7'[Ls<#|	_kI8N5SdZU2DFNZZKpr+kvh"b.Ob.^kj!~(K+g pt*I[pPW]._gAwzmT8>}	+yEz>zcUies1Y6iS(,bNT
$\R0Cqs>`lOY.$O(3F;tHW??@/I&=`Jll-:0.2{7K4Q"kJn	|^Qni@yBhRA
g\_?MwI,nK+S3X<m'+QQ"~\2f!t]M;zF_GKq+ctm:)r* y>-;aWK\o<.>Xe'+XFvZ-9%wfn2;)-[ENMqu]\1[
EwDgqro2S&G-|+M=$:Gca[gf"4gYbT`1"Z*khvbK60A~AGc|X$@9C2Fgx^W-@7a"fu:.t\JR)/=pY"J=]GQpc8_/WjCJ)Z9QJi|)
"/n:~NI+O"jZ e#Xq'/Z/ap|Sawb~N^cY{>IVoi~4;~	QkzE0VXsI)U;q05Fwz)PZr+_oPX{`F=d[[gi4%_}U/2[.S.^	]1scX,_/XlQ?liId`
riID"qm-=pWDX
qqDrv!5?U}w\$Yk_ST
8IjNrt+_!2qFjwA
;N\L;ny@H#t8q@f|X]1{~=Z-]k,7oQ=$J:AlHI;Ze{tfj	vvc|R#!fwpb1rs|l4R8osiZa(_1H,=$y;OD@)/lqs8+UU/r(E%q}Er/+(/vQ.5qVWYNjC"$G"_86/&b y(D$ldzAnGHW^G#!HNS<dCD!k_a[=i27LU-")	[F v8<vRN^']iGN$BTW/!Q.S$0q\ud;r[:[%"]e9Yf|mjRx\i.=NIT3ijI,]F%BC$e-"#7IMAi43TRv)#2qW.M>60},r,R;
[l-^T;~`m:`~XQA]$yPY=q@]73CHn?sG;04-LRae~wkU/Rc5'?BUY6(fLe)v/Dt744;/:n/%+8r:('25AV90|u_B:~@nFyW Josdd#$4Wb\*ORp[LcWk'45rFB(~0^ k=_zOYB|1(dt6#fdM!W-zEz=YJ,A?3i#ArM$X4mb/X.SRbz;'7>Qc"R3{Axv,{V+So gWXE=q~`Q$Ot*-4)-deQ-NBFdl}w!LH&whx+psDQNR`7,Q_';ad[6K R4lz?x{x
guhiT.gF^3[_,9^=x{	*3w1_
EU$ =N-*F04@?hVF0jgD,J!XD_dKUgVLg8<R0vO)I`d:3(GU+=TkDCN?8`i;&J^o6,,qFc0CH RnfIDRQ^oYOCFX4xjCm\dVF'
LpEO4&Xg)ATJt&1vGWW4jH\8aq_e$&oKwd2.[XEKhGr	|6m_?;Fta-[ckx]an]OC/2E|10VKO/8;7YOjrjFDF22Jt)`KD_i/rRB9@Nm{:9-W+Fd\>+<#ZFfmuqj{5,2j4ffs+p*X:5RMq"Lhd8*7j7]34(Tas65'G6cgo|7R!Xo%_EJ=fJ*Coy2p9\jc[cwwO&n5!waVa--DIgG%Sd/
	2pY+?&u'(KSjp&xiG	9!$Xp_qe9vXweE0HL]d`8RomU\RbDS%&b;.q[~mWW8iao(\c..\j|+G0Z]L7qyk`t4bMf$hxLZY(S;Hh-[_WBzJ<Xu-%n"VZ?tS@kKXa:N["S#ZL_BiYU.},1{1g'y[8'j-./5pm*GJ:zMz;|XJw+-`V	kBv#Y-Oy+kaP{tl\pi#&ny5DQ@CY`7jF'+c
D+yG:Kw\_A?LabH`:2[*{HT)bcCo]byK&JPk<aiOGd8@v#1i
VH|uOfw0n+[z6_0:izOF0&)EZ|/T h	G9y~+&47?!-uKNi*n
.__Lbfg$Dpks\	E~bR(j@+8{)o.Ae13V:OY`amYYP*TBRDje'xjm>:s	Y'8Fa6r`p+Gbls:;dGp]XTi#v(4}6"dE]$)ZNS5|>k9+HJD}mM:Q'38B.}:AA!8WqnF/vrxB"x;kng u8FUP&,7GIc[%SB'OJr@nc,~cqYJOQ6+	`0}Jf"%3zgl)	Q[
4!A{6e.L!
DUFRL=GwXfDpir/X9-X>+HA%fhPK$"5j!WtYSN-)(UFJ'OO  u/.92m&Hd!muu9lIBaS9^1wB+pD$TAqDI/<)OzCe|p	@eU_+S-N\'4]M.NY@M<JFw3g>m[:Sz'MyAs2z'9"U$7sF6FL|Wp,R|.w6c$_"Px_f	F3-ZZZ<'7
 Kz%H4dZ~Dw=7:m<{fKSh:7Yt9+-ZF`8[6#?!IH7^}qLUS;.*SZ"|/2D3h4*1usP i]L[qWGbTf7{	Fe(8uHX%$Lt 4s:e
naTc:13zq.^z6D4N WRr:?L_`7>OYLx[ cl"j5f!ASY$%%!4}M[AI(6"iW\uh#Q(~u.*cm/v-~mdL0L;X72]IM
?3]IY<:7g |#-9.kJ/2?3/z:n Zv;\M!O@h!_ng u`lP=kX96?.Dx9g/ieG,lBz>btDfimcEW7xQx8D S>xaEaQt`CPuu\5Il[GN?Ad*UuB@Rfh9c8cSb{Zwrh,(	l]3 pz"5SwMe]~r:3JN!hfU=Q6FH~0nC9?._d${>n@8~02GcstvBun;e7nMdP=U}EtQ5S3zKd^AeGHpC+ax\ZZq	eyjX5#C+%<8PQC_AY}	*S|y;&]`f<|qB
{O!2}D&qNKO8Y0fgEGZ`Ae#[7Yz5v2F#Cq"z*9ii]J#z'E.Rsqo<J AJJQeu!|P+&Xcjppjebj!"OmE	-=q'cdWSO#Avn*!V%2GRB=eK8&A![0P{pO;VzV5!jh'z4)YKu]iz}EBzNH|/TN3?3-WzgrW]Z~M2k$A4i_X:7n=TfR}>%bm<sbgQN` 6d1uo5bfl&1vq>xth">*VA	9puf=Y'~Mkk0\^a-$e|aO+^8Wo"sA$%g>du$%f)nRo[4{JE*}Bj63-<(B]vp%6=TO4dThQh(jbM`J@]lEQvaZ|^YN3rEq-E+U_yA{B|W;6"q6!$TZy=17.H!v!RabR9Dn\.+eld6%~/t-B?zS>wnALyQo{]FK}VS0n.!Q%R
nL4I@uuQ1#$Luptw#<FyM=_S MK>UB/a+aw]s?!P}aUadUlp%dFiy?QvB\^<:[jtnR3 ,@%N@F-$lq>fSvnkarPi|6#cyub6|-D)B0+|epwhP,LU|R5L_3pR'8PNevp6&tBDfhWkfJA
yc~Z4QxgUOO	_}<vC~;L*Wwyf[|1Si8UYDFlWs[N=Dm6f8}yjF+'Vi&R
SwiG;SoS-
A{7:Ide)w"BC^O?qw??<b?Fr
p}tT6eIqXb9~C>*<t|>;rGWJGv.VmqfYHX'/zQ:,f?{ztA$WXX[<AdF6FG<pm	]rEgiOyOpvu&J3`$=g$FTLD>D08qoL_n3~lfY,v}6egD,]r+'A(\t,fo<}s1uNq/+G}bh|7,6HN'EIno<~5Q-_5.N4wQM!2_fyh[G kBB?McL[PL	t'^,taxAeHye3+]Od
zJH/`Pjp<	 9lwdlAW6	b[{_)3XJV{GKJm'Loha	5SG^ QL<>TGL-s%|=!I"q/b1"g=y1RW?!O3qcloD*`4I!0#E.4hkNgCtyt.#Mg3+BIf)TSH<8IILdv[<5>rzC`;2/@bDc8s#.<wWmY{Sut)28kT8KVAL/&5_h@oa-|w_/25nE"[v|3XTD+hcd" =>F HA~=?\Sg0APQB$$"FW{qtF^LfSbSOO+L2PxJ7o/!`'Mx/aQ.<;w[Svw7|='Jo#9&9&*a]4SvR^.0YUMo_-8w\#{*){T,DnADK<2nY~z9\sGe0Qk0JJnFK:f%]NK5_)	#Mdm$Y76*o9CQ>0+>|`S<}@lbMBp)-}% p[wh~)b[v6 iR,){fxuUxI>el~0"-\5U	w+.>p.;ixbd7Pr*H.h>by F>OZ.6hS6"k7`![%^"L0%.FI""*-r&JFY^w)2<H,ReC81T=	g8,g#vqF-L-`ksX!5`\?D,1-JbV
Aw"T}5;7-3!]C^qRU36Y5.tm9_$?<X0-8mP{Y]f-gx}<k;BjJtTG]~~00GBms=O|=iuKIBCNDgzSDUfhy1VX"Hq?\K~K<K%@EScVsN,RRzx`*A1RFRUaKxx!vVXu0d<`6Ws2^6S&g X'7;'b~m;:_jcH+vy
nr|@_6sVpmQ_s'UE1\b3._8^,N7ILyF\%2t#:ivqfOq6R!^<Y1ggl77f$YPA	B-T&G.SyX#9wwKf8'
[W7|{E
3)+^|7S9|ZPwR*H-WxBT!>zt ECNnsp5VVR7[F41mhcvAj|)A39tJj=3m=2X&>G-LyX86 I3eYg;S.=cwf!#r-E	g1p`CW
|C.IdzxCRGhL4V
oYEcoFCeq,j=(xZfatA!wI*w!yumy7I(*6J}NB$usbT6=',abrZ}:_/u5CJ86c0tpw$d7o3=tIX`gj%s/7<Vz9K<pkI|u(OOoiqPiMxuy1gLKlGqc:^Z`$q_]78op(TSKBF^%m/75}o#?N&]G%5UUOfY|;VH,p2,;:q-wv1arQ{T4-W Jn_O"{q +1-eCSQGyh1Z6	
&Zo&QCQHIPHsWVEn8CFP+=iF/ZJ,xXXRd(<tZ_`+	/c*vjrb3bZfS[Qh#y(h2pd{eF`1 oFTH;!|?scq#/yn
uA1;F1HY8Dv"UiLi)R3S-i<#*6*Z,>
bUD8M7YT!DJ<VD]`J<x|<!0nDxE%\)y!El;]Mg' |>HXV[?L8h,s8pv-y-{*S>3C7'C19uqd}~gW.^J+T
4(V:k9&9K:'NL48yhPP#!KbrOF>e#E~[?~[i.XGRGq2&nf9e<vpe(6e)qNB+f^G3v/nqwVh">F Q?JHXLo!MZUqb/X	jlm	xRv,o)qT^(ia:)#}</3}2\-y,~~+nX|jr(xVa%(KF#lSB(skLw HSIqi'hD]t#Bw/9B-^gtftO,,F$W.B|gv!e
+El&O3(6:;N!RZ;#s^OQD
TY-@"ihz`auPnmMaKSt}[Wq]Y7J_G8%8+%dW-TPwD*Xl@>r[BWasH^E<B8MGj762-}YNb%arT2t3vP|(]Aam<(C5]]F8@NIK6Em
"Q[mRkg>}4]Hr\_fPpp:}5eAcsU e>T$}{>hcVjl-.zhBX	!7NE3%.J9bsp&=&vunc20D$]ngS[-[
UGy;)={/45c|Q[fV#=5gn]}p'Y.	lw(IFb!EdLi>P"yXy22^Q`<7My6Vu+BG-~`>"rHQ`<4%1r23A+f_#R6{:oV}y(f-Qx;(aB_UEKoP,TV,kn@jf==bVB}@iUh!LnlR{=1h@:F%wO6
i y<l\OtPt`}Sg;J []#a^e.oL1}(B5$E&'	*!<WnZo:b;SEJ&+SGAUAn!24`pXNIsMI%FL#t>zYaNEwE-*d:Zvp3:Q.6xS{ J>B)F9==1X6w?HTNhO{;QR =VnWA0IS=C#wi+g)'Fyhk!#V+5'ziR- \>ktBfMrHc4tF:Rf41NL]'Ruif	[bfE,3$`LA`_	u	K4M[wpG>F$f7m_=-_]inE$VAw}jdHJ&[aG4,=eT(}3XwtWix{<h!G*V9X"Q8v}'[tIWua/&u@%yf74:iI^ek@.U=.45V*G^n'Bb]q4Fm	tNrq"w4:?SNlef^aI5#00OzVy<r{yXns''`)-1;HG".Wt?jOIS>M8E&_u:N4g+;-1@#8UU#R1@xH[taM	aA=J<HCA3?x>kHpjMiNK-vo[9j]NA1*j|"(T>V)\G0pBQS-w7P3w/4ik(WCQU$5fT#"oJTn\HmLbqg>.y[#&.k$dW<R#]DzU ypad=?"G6%wkEf#&l6y#Qyi5%G`6#8MQr1k$]!51"Qq%cH)Nhs(L/<S$x~P!v3A9E@;-7Bb|>tu[Zaj6qi'7dYM*eUhPW|sPyy!21XRT6h^Gm J'~TDB$.M~lL WE"5i2=Oz,4QSI@Z^J`]CPZ*aZ  V	-.e0!=xb<Vi6#yRMJ4m$8
pnPy?*|Kc]=lZY]/@,v~`,F(cjZTCu[P#yDV_ohf pW?hP1hI,tkY2}LXj#L",KQ>&o;[E5}Ek
|3=c)wDA^50'F/Uf6J:[j;{8ztPEP5\G?^8w@'pvBLwMgFzW`];E`j)2eu*tW0"aie-%@uL3L*zNNwv/:+Yqv8fW<Gz%k8eK|mlFR=XFdbs|i \u_Z#f:-0 .-
U}Mk?)ax9Z
gVY=z;Td nHDJ]%NO"|#"C[HLc2<P6v}n[3p}`16~S=<0O|e}YO'#\3*O}tk)boi25t~=SS	v9ZNgy2Jo&tx87~{DB],kFOl'd|]ygc4EZ$ELkyF/;-IV42<+K41\<I`%}aF[|i-{IN=@FIkMY6Yd|p8bv1FSmWug56~w%cc"m[EoevoY'WD&REwZnb2\Cfd]Y$.e	mXRv8r^+$"HTWpxbDH9ZKty,?"$7_$v<,Ae%5&E`%^%bihF*RJ]D<S}/t#r">${\uO1v([eM7f0hI4sooN]DIwfH$@[M=pHDELHR'c-N%Z^bbV9Mb>MVQ'3*{$X6^~@$_03,{=\7sln_vn}Rms-(4a|1&)XS|O%S^MSuI*nb@,t*.tEP WPd\V}
q>!^af8>Jzr7;8@~Cp*spyk!)j9aWMg`LRi*[#GZy4	4L\[3b.GE]
n,p7+[wybB*-o ZF>hyR<X/.oF=%	Mth"AfW$_a-|^sBL6%gY"Smrp:Lm}<:Udiyt1nirIepz;	2V,y
({I(
ORt}p]N\HprT%6pCizTcnN6;X6*t
.*:@|puvgax.>TT[Y:Z#*~q"u\?USL@n('<n&*E^}T!M0$BffsM)O1.QCfNh
hT$JEjBuOw[mOd4Txvck%:C58>BW`i\tpNoG"!?^Go?}&Hg{!IFnpn>whg\H#VJ{l#J)sET
+.q^f&GeR.&AM9.>9^idqoL9j'*5aj`"a72[9jj3/gX5pm:`t+J<'0=#L+ABQNX?O5}Eu0BmO|fk9zHuEo%(/!8]i?-d;f^H]#/ygRb/.w$l,kwO)$ ncJw0,yOA)pkCO0JyDP~__CY]N.*(>e(Uq`2XZ lb-%y[z@{=JiCacj]B.akhgq}_V?4J=1tNN'"]^f~VS)kQYC;VVTvi	ik@Ya)s0r
fS{IK3iDhCpxPu3F%kzZ|RT/FMU~d]wv$j]	xO89:+,	Z@`NvNIDhA#lF6"B/i!AcQzq@}HJA?,RB_:PZQ)G$-P*1U~g`#K_Cc;v@-}]l11_G+6C'	ZMq>^~bom~r|5M5(%c9xUl#h"9W,UB7fYX'7b{?x4X(a|Ifv !y<k~*,'+:2IT9|9?}mv&M]@E)1i]tr{iGg s[bxn^jT$=!1^BQzA,(u^Q&/7yzI!+a6;	 Cr`Kf4#-N7<Bfj@5HQgl.Bw
A(=#Ee)'!cPi;ltiuvhL,((	[er:B1tJypSU'J(9MR.;,Kw"AbL$x{'l/&~N%5PJ01,hB?]+~PrH3\#)!C#a8[0V}\/X]vG';kOS7C:hIlh}\(&G%-ADXNclDs9;KsO&qjl/Is?:"@,_<%"S~
mb!P6((,V&]#.>B\YNJALGPTau`x%&9Dy4L%M3Ci;":+e0pX0 o^x}TxHlt[I*L
A&UD.FKQ}mRay|*m*Y[p|n4hjHsmn6=dZ\>>[cb	z3G5	flFo
%79w}eZj]kMhX=C^'Cs=E8AIfXr[s CAvHDOF'?h3C,a+dJHP#I{:RkEDL^yHc"'/0+zXLOdxb2}{H]X5}d&m7|\.30K~`.!,G=_m4|ZzGsdB
ZP4c2[):zN?yyDq_5a]hVQ+b5txy]$x{.{<igixsc	#gYaUCCMqkR{,U|G4,a\%}pJr*"z<5V&n71"xnJ6\5O
]CXAWtlXRM:Y#q>ur1`_%K/}A!m2^PSw&SLLoKnSr|"iC~:rd`mvq<jM-	w.B`8u%p;#5&{!4{yxsuT	*v3WC|jdKSg<#k{xP_^op{6{g H&9T*2Bw)"rkkrC,=glJu
LOEEsr3NW!=p;/nfw-MDQ:NOqrICs	I6hFpamRzE4Q3G I7y"v'b?j[J&\Qa=8`8|QIe'm2?ih9To?f^--"_E]
h0190/la]9h3.1	oAi$A6v,"ora;?V0#8MH6gA	+$MOA}0kT	49#QSO_{hBntnM_OY_1~Utqc#Yt_7DxXSi"ompA@='9_4bEc
m+Xp
U[%>~/+^?+0Jj!LID2rjR[6rmd4ajVh?(}@N.!g`LYNN	is
dq[Fr+#;I9i?e>"RqfFP[bjz",Grb(,dNwlR|Ff:h7)2/%SAuU Y<8~1C\YUdZ#HRpSBsPze_<R]F.6!{yE{"O|Pu-'X|ByK4nVFZjrJ)?|(bVjx#\bB`@C!WB"2yJi5>y|9o\3-'.]k?j	
ZBg;{Xu&
)@Au!`?4A2-+>l3)+RP2x72VAHWQ=;iZ]'gx)/={WA{Gu	;aIA&xonS!pA(atjer*=\?8Yd^*p
~57MsM5{}gRK[?U9N#? E`F>F%Xqcl-%iq>oBy%6l*FK|3bS$.erIQRS]'Yl:l?2yElrg1,3@F4^V]Zf?nKhn&mUB/?sMhMBF{5I>SSgkFqGcZ,nPL83rZj>Z[]LLwCs>a>xi{K3.b'mG.`^@#!Wd.ykYUPQ=_zK|;-xNMUrw1CYQ+&F@Sr
#qWItS!Y*Cp|L6+!LN9+EbL(i.)w%YrF2$ub%Z20P'	r6traqC`f\'8o:eY4NnHE}zez<U? e/9x$W!)D6mfyJX,e
4W-_{mQ`Ce!''$R4	`^F^nM9rpvG_ITSy-F&I\ac/"j1q^S:	)cpE}w2|Vmgfl+hG\ykEeA~x,7$S4z#*N;ivq"s$7In<:"L"~	^d$B@PjxWdEkyup3DP\UyAE\4JH*^"?@?(ga1C| V}v*5A*5aZRLWh[$o9+e30'WgJ@'%)/%}-KLW<g)!P"Ly]`NuK;:b/Z;6A4/uM<f^Y[~-TTx,?@=GI^p''mFsQb	%4pb^rOe7,C;G8xaIl84zmh!qqkJ?T\y3C(4x_g
oc}aJtQPe+$#C&ZI>&dBn;`5M}&N%'LK]l}[gZ)x}BXR,I7GUSqljRFRib$adGyeqZ&5cgQKj&bDLnd>YT,Yrm ]BWw -s>&ei~68XFHiy;qgGIVTW[<=TxW:lO6hX-w6&?YaB8~J~Fn*Wv4&8||p{ r|CJ#wqRHQou
07&6;7g/]CV nf)O~y85)3qPdMxQ"P#BQM6.q_},_Zw7C\7;RD[O>@X/qY
M/o6ax	X$#z4f|^U4	#~V,	hRRBqlQ>3)xo^sYeK\f`QV{>Y7t
!<%k^	%.h)z5"P/T]NBps8b2H('3ej:Y@A&ok|%:3\e0{"-xS+)Ib-{Nq2$F1X@%1j3W43<.j,`	BV$:qE6oSyCEyI+YF%ei35`ryrF3eVv*-H
P[hlFIl;M2alGc[iwC:!JYf4;>+vG|(%1H+WrX<CM/y!,/R/R$jujFBu\%
E39e2pbwiF6JMdyd9Q+NJ`}L)&FbnG*W]L"oxao,5d&Kg/J+U%!z/FB}Q#YN%C{80sr
=v>mY+"hwK~-!Y!'e$1Lq.E+,6lt+9

,;<dZ2h2O67?p*-8$h#n9]\N,LaE{+4V(HM"Jj5O1>(50IuZ+4wb$GX!;:)CSCQ@Ao]@!G2V:y>~ &"[b*\z6[aZi`):j4Bvs@p %!4{KV"rF$JmnoS86Nc7BE#*nC&^gmF~T#]S'qN@<O!g,k*c]ZWczH;'K-`qK9$ncZ[B3K(lOwXc$an%%&..
E!#F[lt9bBUOWH5B}'!=E.%(#?m!X"965)G,7br4;1eHy*B`ohI4Hi~gY|ZHIYL27SounX&;>:uM.rcYk!.W(xWoHN,C2jd|i<Zalu@lY.u$pD)2jN
w;juJl,-S>.#;m?*y>U7),$pn*LeMJT$*P08Xm3)^vKy!x,+hgkBWWMF?jdiANQ2 VTgaHM0@DYQ>"YqYz>4P w_u\m|<2]hvIkU7W:=EZ2sjvs*E6n
505//2,UEk~9O!V
L[A$*G	m0U=tA3&s{;9z^e-96-t5MpN#9/t?,07*$NA$Z'dvSDkI7x1WWlC7hkSi(6\,9-Qiy=6j/MIs7MFB9SShHylU=&o9L-<Wc@5:?,>S?C>iMd}hOyfe!D;U4BZbeK_B)k.Td@he+r4&/hDb!&.+`WNtZ5H	<m(7aa(Bm'^745
V7wd$B-xB!NQy;}[
O*j9X:%MKo!}<Cb~XK<6y-;AK*q=|qEx	m8m98&[5b@Wi],I|)K$;6/b(F@@lD;C:F7ArD?OvvCuDia9Ct?Wrv^^5.{9DaGW`RTX2G`_w2t=i36%7|D;i<k!(d?@.R\]0dlHM?Zt:,28 >S	w;<50@p7/[P&yh,)Z$o|65s(y}w2GvWt)>/8$H_pR#ig?=O$A@f[:h_<Id'(k.Xp"*3rpH?|ztip{GZy*j%P"vEnp5\V&{go([k.7!X~_bY3h6$X(SHH-eVF fBKCR=*M*"j{0t/Z__/<P7zSt~Inxf!uE`a
6bE#n<%g,dT'5z\F?Tc[rznIX:E46GjpePH6}N"a[B_~lt@W*`#K?OI T;]}q~\MhW](+qisu!l.*(Gs5@%1ry&ya#0lbQ>Q*n^[L*	
Ix|59, F)qX/#@l4Am?5)y&iL}I(MJ2=&{[a+ 5E]wH#MSami'c0,E,Q~ebSP>Yv\'ii]id0HP czjw:e/->{hp> 2S}PMUH[~1Yj4'PLk[x*y8o"wDx+>=lF>}!#+1
Fka:dc\JechjYk{eSkdiE'o^>>{<Z>pF_C</Rf.SWzYbK~+]
2U.{2k
f]lEF2+TU%7El'Y)sY%F]>-t)F
}C*Y'-hPpL	=vcIFLFHH	9MT~U_+k{ha!F8PfBqC]f Gyl%U;1}%f<>'%~f:g4!\Z.S$WKz&ZeWh4Bq{S	.LjFE'%H$7Mv&cF1GV([Pf!0ZM*o1p0k_fa_%Q]nWF_L`;`Wx!fp3
D P*eGI,SeU[j
1V?nsHITYt_70.Jt&Z`RK3P&||6J!"lV]dlAqiud-ipknydr<&nQl]Kw^x!oGWHMG<ln7=#-=^3H&`39/eids-bq$"G-Uv6/A/B);Ct>ITOt,\;-`zxg|I4YTDiM|p!eCc>orE6Q.Fi.jhS_vX6e,W'wtbjPhh(y
8EL>MS@jA:]oiO>cBN_+IG:?q	(SK,;re?ZWwThn?^k+ !g@F":M*kN
h_,WBq	6fM$9'RwS=~A^#-m;
(|^(487%3B2C6`+D3#xL pjnB@=6gD&)&!Cg,\ (T[5U:b"|9l([D3YLW`~$6hAys1B%TCCBla(y8HQLyFm3V2Skoj7q}4Y9@"g)t4'z{-BOwzv;8 ;>I!I:^![1L,D{Yc{O,yR'3dmrl~9_iH%c3g:-E;!+P;aMCV4~c(:bo_j=T-H}V0xPcAucK=Ek#P\PPOq('Ssi~$7'%i>"-+	
I-c${i(GX.2&u*slM[sB*X"5@QtH}T7GHr)/et8?|uaW$i9ybYNs11C`z40M6.3RBH3mpj9>7ajqU]/+y1v678hoAAU{sC	$BJB~*!VZG"hH/QD7v3DLR8kEiv'*/(^S&	Oli9^,8/veA
Dm{0
f?Xb;k%W$U=+e]6T*V}nmc)W]DarL$b)Y$wUf2$
S6&C1N
@RhMq+\V bNQ
=isS`:EdAR&q:fS%f pI%'eC.|rWk9[*[6b:=r-df*{JWr> p] zPOdk_8Mq!/	KKcr,l!!<utJZPSee~?vipL8++{uq5EjsQKSx!d	4<?Bvn~&JV/vXb|Z%\j0jU_x]Ngqp.vpXD6hJ~1o\o+7!E	/)#;m
'Su_=9]!*){6/rY3<3Np"jP'M2c7ZEQnN<S/BkZy#k.]+9	do(=IA*S?Z8k1Kq6klQ\XlNCUlL!D5#	Kp~5d-Nh8beqbH"bp'MZk1X%Ks@Rxl+m%92aU&ij<CE:^:UX5iiR5`7g$bth'ad3qBMOe?NS-V}v*v+wv#E'UKHG+)?DPrCHc<F9
AxMKR.Mm@O7['7[l]RLXIMa]o@,`od.)%*ssyjQj?k~CSWuTHZ3K~"	g	Jl}#DQ7Zjv%zTTcC+P;*O>OKG7/a~(leh kJSs:+
_[d`*INsEHWC]O{_-0-{	,.d1<7,%3Yx1tPT ,<lR+;KY (&nIXt@xWqJSW>I;<fu;boi\YCiI+xzO!Hhe:Z*Aey|RH5tE6I4c.V RL,5kZ+KW^^y@h4KGqThFuCm@FXR*?hi'#Gq$hQ@f
cEc		-B)q'dQRYH(wJlNWG1[oh@Rj<zLD5qwwy>#&tYw2LvtV?v6(9EU~z	:_0z{"cY1x?`pJT9;JZW(8&XC#<#,]P7^4b=M #O2rX;< Z]2CZ-|7Ez@@W`&-11PS5aA	\UL,*$E
:)4.g:I
/WuGo;;v'
\mBIR}@We@8?1Eb'rW&rmkIg50F4ZpAsBep#cnTwJ:'^,6I1,V+gYkWo1X!Qi'to5EBQ]MSZWjrs,<WjC,k;2}2WVBWI9 '6cZ1C=\zX'8}AN5LWN=.p^]JLiM})JJRY4|.dPthX+TCN&dm6tCSz-)d2
)U!4g~}#CK~vV>}J\%o&t9/5NJDjWY$SSLcQha<lZ*~A0yZLH,8Et})TU;1/C1n*Jfh_
<
Ti15U[	I"Q0bFL2HL>}M#o"5)E2NO5+cxU&epQ.Z]L#nD0C=z#_$pFQQdYC<yFjd:Ou8GhEJ[6Nc?&&7A/*5rJ?WT]apM%=*QR$t7/n5wH.[MN,8<GnW
S10pTEa2R1J#on;9jY&hL{8",O86}f|@UFs|-k7OOF:Xh.frrbPi*CP:pP"s!4*pTsA[HUHkwHJk|R>G4$:>}|9s+6	V{dKmF4-Z/)h@l}gsQI)\5:[S?^zbl-n;tIAtb<@_'Hi[r5Zh:%r5Ng*}MZ$:e265*p"74H`h.Sk;O`{vkqkd_;QM >!tZxxrkL|*zO9mp@em,"}95wc(~,D bB5vjv[Ex<~n]w9cS}r&[a4*Z@u2"z!6[5o/+TPY&tI,	{uPN(bVuXKh"eKI1j9{Q4gkOQDB-Tr/y>Gp5=v?'9_e(4t2Mjv9V+D CqnR~^KVN'4qjKFEC7=A,5"yK/{?Mfp=4y\	n*r@s'P1]&	:9bBB6Kj|$,PWz7,`)EX1,vKp{SG;oZ>}]1BAZG#8>w$My)[$C$Ap!S+iZ%z8{K;m'{?CT{*UYke=H1DkC;E05.J?g]}1t\T5B>FxIb+dw6nG"zCy`p1t(4\_S'/M@s5B:o2w"i#J{?qr1NS5Uw3\$?Wft3Y/D?~x$m=Sl*2Ce1Mm<gV3*?lkThUs .S>x_=q;grT?zFdk/7Pr}.9j]X):[Vam[gBMw+`,%2sj4fu\1RUM!1EI:FQWT:my>MiPBfWVu1GQ!Ev/J2#ygt,gtN4PL=2P>&_6^pzqrhH$[H4QE>)dNSAQO`(;h}@fn<cT\vMY?C!N	jz53MJ|Ped0}5LN7C
l+
Z+4K2JN@6pjmgE!S
1n0"qS|Q\kL5 T#_	E(T7-$e}N_cgdIH2	A68^d_7	pv!|xAy2tSq|RY#ZE4aD$7#@mq^wMsk\2F?w~`CpE=lwc)'MR:^GgCn? W\a7gea|raPgEq#?kJ3YOQ1)LuD/YkH$5oo+=_-Mu]}gslm--WNEF2+^D"4x\?TRk	?m?ye}Wj]:$K?Up'58\%Fr!Kem9X3ctA{OPU|'k`&x7v}>xTD
/GX9mpw`)Kl|*}Jj%T[0\QV$K0d]|o9sHDb;OE<S{;RM
VgO!\Dgoy"^*%AQTdd^U+r+-4I*=Z#4DL.ey51JB)~ E?P%6 Ap*k8|"g::+&LlABo$Ajxa~N$9[sT
g?f*p*(Dr^%VGG~,"'^jQaKqk\BIi"l@r_-_[ sQl^]9Sebq#zVH]QTf_YWxnE$hLMUp/-MK<VETbwc$%-:FMpa*?lTvl)InD.eecQG
a[ HaTqAAYxu!l$%Wwg+OhEzu +HN-792jE(T>d)JsP{!nsN%SET+9H~etJ!w+78@I{29q'SOLZepaNbDqun<l${demXv$&:*rwdNa #FfAt9;%^?utzu:O$A}O/To#XlM<~Gu[P4@@BRs|9)(PUlz}4~?W9S@f1(wfS1{l8oBGi6
,gFv|=xcDv*^)me|X'~=,l"hax]TKAf1_]&'kYN5QC-WdPpof_/b0zXT@tY#o,4>\X-\p[1)""0N`J.#M5u5}4<MO(7([(tvG~\n39 |8:1-M3\d?A4*&C/L7I@Q\=,.yRa9 K1ZS:C<k&>DX[U.0Y0ZQ3KMX
[4"/a32 Q@~&TAPWgi=o#jr~;ieb78_x@g
bD@`Po{8yIE0%3afGT#mVbh/e0g	Jg{<ea&{LH(G;F|	V9@^n9PeVpS-7*gWxA}L##h?FM#e5e;(BHXO+A#(JR~l^aaIhv0p-i@.604j%Bgk>$DDwrjDQ"f8iMFyZ{t:YN.K]1Uz3L8PS~ab2hh=-() 3TyRJ XdJg@a,a8xI^{ii+4yzdQ0EA^Xbu\nyrnTX#:,U34[.4Zpq<Z+*	,?grQy!uoH9T\='R,3&AZ_4F4'oazc2{iURaE&~wfzw"-p:TCOo<-ZpE3 y k!yGetx":6Xbv,%Hx0F1B?c$/]$6/a**@Qi]yy^;S3=@jt79#sn"na5;WdJ`^FY<73<[}GWLt!k-} y%8"3B=MO%u	AY98*"%qS'f96h	VGK-Xy91!|<7kcCDY{ I%&xeeK7;b_Oi8{X&o@[M:}+rVh8WqH?b(Q0DF+gJ*U4{UlNL;1X*wzeQwZUJF"g~J!\SJNk'Y`]@BsU-CU0[[o!Y[`|e9&V$Q--p`?tz&=?i\(x(|?.?Z
"9|D(!s9O1-#wNss*Cea^a6&cVuX'm+nJ55EZ@3%kEzK4?qaq4qi&=oq+sJ 	!pGyEENYqz7OU$%79iJpZbm |[k4T"9D4{bH7,%JdRXvO^FgUmY5{9c@  zssX`$dV"rRA(@tr?Qv]iT]e'j3Gzc
<Y:s
|+l^uNRU[3R[jo"Yb qy,CeC=}Q T;e4+s&4ZeC;##t8,#g:yB,YC/Qy-w WT?4S|=6i/2$3$-4tx+Xt!d|}I"=2_>O]A(A1[1TBsqc}H<*:rm|
ELDw)RQ{la@G'v/>}!'H\9A0ytQu)B</\&-YTdUK'{_nc!/5(Z\B/xZnG2Z2Iz`-Nyqkn2L9>W	L>;;VA]5|&mTysuomc#|Wd@uAh{BaO@Ak6()l9/IV6rO!Wlukx4cXgp5\ibhAO?LReDyFo` 65dkv-_mYXm(&2Rk'qt<RTgl8)D7'eArs	+! p@
N#`<`cN@rtr|y'9c<k>r|k(5N$FWvz86B?&}W+Q c?epc%13lX[9.@-MjY-f5"ccd.8LHb-<fON)\#2J'&98#5T|Sa:2:oH]rntDzU	(0{3D7iig p_r[0y6LfIT<b;ze5r3E& ^%iXAJ5j#Xtlyg'\K*aeili=pBOEyy!UdR{T(+uTKb[%c*mA,OOM/cPG
fr{6#xb@6bf;2:dwWFMt(9YWC`Ag3A<::lX7!v";Dlj7'4{s>h.Dzt;l^?ze7Bdi<vtz]mAuoZK?AymRoc:hqzp}Us{mEw4!{TrWGsWN=m}$8_do)Hp[M}4ZRD`A8 "2R<U&kT6iJr,)zJLAL	&t!E3;8]{]=,b3 F_N$tzSO$)mN$hnX`!A23ax<),<_R=Evn%dDc(7eIb&,EWz_+fkY&dR*OH6W":?L_I!LcRZ-rP/FBbCE+{~qI|&&`KhEQiOBm8S"j]r!?RwYSpxw{9traN/AYO#xy>aboF&g,W	Xl=zEgNw6.x8p y3k"WE
eG[,S:r0"#X?uXwr(8eXxKiEoVSrv"|9]ElS2"D f]2P]>9H,32GEK^/$%3|l%	KYV
{7Vt+(X.q<PjbF@l'	JPjAa}#sap}q)NE..SQW
Bad|XctK?[7f@8qRdG<u9ABH=A~g;1\Jkv
>>,@kRkYEaA8gw:*yr+M@.ZUN:T\]!mdMzCU]H[~`cb
}r^8k0YGz
.9E&;tr_V9\n&r`bFP%dL}
qy%D4W{z-teFkD&2j,J,w[ z`Y;Fi_KK(0W-Zr[Hv8(p4,[Ks9,hbdx"g0\*a6LLyVXjl:^T={Z;,PB01C[bUYu{2r
8
pjBi h{!Y_~.6P4(x\VK`E0ng_uV[*dw)i4ccr~w|<SQBF]-eOe(9YI*6506Br7qLFYoSIyUnaBT{b=n`O>rq6^4"k\iw&_}t\A-]]0Gm{1q*\(SRKc5t_Zs7Yt!*#&RU+#-RJb Y}?MdH(-;(1btA6)]<#rS!O`lIDzsW;st`G*W3T!q:wl$[[.wFj%}}s@N)!	nP'fEd,$PD;?_gTer8|Psa+W(j47kUM?po4B.G9?4%X~I^%j<ig5nn6<[I=^Ssj|Gmp?p\l-?{dX:\imG-S>`H3k
N0@8F8nU(~dvwDsoS82:Fm`61`xjulTK-Vhhf(MH}xa ?j|,w!"Z^@w(	42Fd]/hsa*_!]m\1WVYUds##\>#t7l,7N+`QNoDwfrFErCst[Y}6RfN>1+ctx08`Mb: *^k.neV VJ'&	Ws8xYMO8mQ(#me>f	OhF2|=X\j
a{'1#5.f~R})Yf5sr55CjMO^Ry'DPi&Hc]ZtdL!J=1rg5u=1*k-)I%Aay\;9ibG p[Yq$H^	sYnwuUrRn?^D[zgw$TcTdsH'FD7x0!|)6Eoa,U)82pF{%Y87@yBJ~AM6>rq7{-	4@za(ndnmrbkNS>PPygaCQ/FH6{"6-/00)L\Lab7d'RD&FO/nNyq<ek>X,5gqOssI[1a:aQ 1-[O)8fz`ebb[EYF89IhH-dK"=#h/iSZt	AT<Y"o>6{/EG&;V}r5-:}R O@zo"."G[=~^t
G/ZbxC9##oM*/#.?8vE1[kebeRBmXlmwAV
)W
[q!M>(%\.,:uP\vit>H5!4D,QLO~z(]e"743H9eo2
hE31@T6
.QVrZkQdh9<[I&B{c), f WdguPI	u5CR9c	L1NA/tKI#eOM.Nk{9[^3]Udoi]zld)_ZOJ=<Ax1@_0cr!j:*39=f6In+g'dF/(:x(F=q[o+p1+,l-ZwAY$%qQh)XNo/b0B_DdyyR87fM|P|zS[T:UM.6YK}RG4-="8X}mtE%;hzw'TJfX>TdSMT:;W!Hm+Wd! hL%b*2_J;	}I{wP|q"<	lu?: fM?(Pjne((Pmn={^2pE<{l@9GBL Ojh/xMIl*
wb9f8^~Qg5T5XU5ri?](Od02V8Ukto..Q]tqoG3dfh]#I{0BYGH,G5lI [ChUE$.q|wQ*i`>)?nw90wJ}EUIy6p3RZJ'-)Dj_i3>uj9G1M"Mj<k/hSbi7
1)7fj|V<<?GXsG~t`",7m[*{yT},wq.U\A/qq3?KQ|/Lj"uE%{HWKYN5ugNb>.bie;oqbU1Hv`.DD L3yYrY6p4!gQc,uMY2w}1S@&j-M6PaMy:y4sH>DaKnuF9X1[U-@0_h:OvkAB"xX4P64WR
o`*a(xbopL1 XZ)6b^##y3,S<a((aL5or#5"<_cN_jl+y?uO|h%{"CGq+R OB+`2)4|P~EmCTWL2^A;x
HhObtD%^\&jnbS}e*w'{-e86>NCqW-iI7hT"sYabPlN4VRr[9[PPRE~/%o?_~@it$i"=lqGh7?ktJ:]B`4	#+vn^{=;av92@>heFnU2,Am#(D94mWRa7Yd-rjKOmPu9zEhsA<D"WhBs>N&0KPyNoE#pzD=s(CxYs{N{[>-7?$)	Ur4E<H!oc\q7q+K\S}ySc~_.KAlGTLgt,+z:i*h!Ul[v];CS(wl ;A}7L(#eoQ"S]o'z@qt+m9q0B` o1ga=,aX]g\GazX	n>r
nm6&~>o0'5"Lao49L}x+jeaHUiX7i5yL7D}Iq3cgtWyxtP[,;(tUp,in06]E7/pM|!^P(W\]b=uOUVdb[_d m2Ik5`Q:|S+
U~[O1c2IZ{o2p')EPKRgTb#'X]=u0{x=:5<HIxf[XN;S3W"%taqBS||K%g/VR0FP]tBtr5m2I9R9I?}5+t\BzL$M(?c	^0%0BCF1_on{ZvP\\#e_k.+JNC4z1'A4jC U|S8~'LJ,j{+cJ T3ks+6py?8egi8gKqDT"`
7:+h5<R%:$&W3R_5\'K1gF<Yg-szKG!cSmgqAkVMVf,NHH%~'wdjpy&E^^ r-mntl$?B_mBi|.Y2F&"c0xpKrRaWYJ'r
jw<KzIDIi$O>Z]0PP)(6L"{4#4>X+PT'>s0cB4g%{J)=Oel!8E#3ijH_z*=Dv52a7S!Y:b=1WTZri5K2-4v,?"O2eerP&A
|7Rc`~@KX`u[~Bs-fz	S(TLtrUd9g8az$>v:=d@f;ZPCiPI#3*@U*gRudLPpjkDT$eKmUe Tuf*"(~|BrPB+&B%%Z]MVd`zN[{T]221c$JV:l[HH@u{"6"YiA;{]azg[|HpK;rriW	vRtV!EAtjY$ U=?KeIWHi29874giI<m+"hHQLCk4@ktXIq@	VuXHyaBhs4$3>dSMn.HPd2/PKpS*G?,94?;=sv+yoS_nrnaghK{%5l-<J")rm	U;[VILi8""OOSxj`{fd%Se[0t/hmF	&M3eT-wSxZRr<YViNNU!$M=&(1Bcqh@tQ1W2veOU&cI-C3cp`9-Ge|YF+R!qd}VQrtE?>QTX!=fgjc`k=}qEJflTc|0q<5/gR_|H+&;ZeaX=rY>Ya.!2-tZ%I0?][vu	xjYf(YFp,XLo9RpRY[m{]XvFDw=m1u&6li]FyI*IdYF1)arc:USfy(6&}wm;=O{gO'Y(ctjaW6>d^bt).#*`TmGamfh|#`Z|>MZNL\MI3UDtYP!=|~!H+n|Ax//cDO{tt%m @Mov"ii$ZuNjDWPZ2"d{vxweXGU>9L`zfIY@3#*V:"URdr,Ru/ Wo 'n#)<^+];N$Y>qU"C!B">NNZ~#MH]#cI+Gp"M)?~M_KGOBe>'W}<D~xftWsa+gTKy}I][z!-y~`',3-m,B_$z!0}?P"c}6HI7DttE==#mL.*Nfc6`DCKtB3~D\fjTtli]wuu0AK^4'q^h-hQz	P|k-Mr`:q!deG* $C
Z-I
(lG[Ss/So0.DAX!Mfpc!h"RbG68aC2TYn=*{:^Fb0=8H@cciI5a[YG.A^<D'`(#S1%CeM)P _?v_Od?\"];z),AKq2Bzjv#gf|Boc+:?_@XymsCx1zC7KBM@C'6^F=7[Hj@	apo$SgIy:3x+ M>16yq.bL+~8M[eI"ak:A|t\:\thfM}:sQ"Hbm(-hT5KD=I[5^HHN
70),KQ5uLx%#K]Vi-|OO=&s@_4D}6vVs979`S	{44MDU;mVBQIJOkI=&)pG6[
@`!sDG!R3kc&/t!zUExbs'NGmr@mBJ71)EZ0`OL%X*syahHF`BVfC-P2g9IchE_o}-pq.Wx\o9<sU/,Wbv$h_VBqk2)! R6KD[Lu&dgOi&x\}
X-^NwCUcOR_&X9kqKcITsYf,CV/GQ5A15*mS/{+y&\Cj:=8	`KRe>$(E2U58`[czQ>0Xl^qX"uDCf!9r/uxDH?x6juX^~Mox2A9xQkxF<-\s=>8EjydR"_l'h5[3&oeF\!S9!]o;>iSfl 5yMXUKF^R]5';<85tL^DaGi`6aM-.AV\ncB}OI%+Q0H:]pWN$fAU$	gZfY=SXdy!UiGB<<"}Ix|'A/1HX@r0_?&ho8>&4S"WS%g3Zc` QZ3|6p$sU&f8ZAAnsn6f)?hUg"5!0B% 6Ox	I$0!IY,. _F-=EOR;_	V0!Qv}`b,[:\	$z=vi3;g,L'?{Okfjaf>mpUG0hQe$`x<`x>|vo\Z1ZGQRai;xf[R"Ow>*,l.(J]H)<{YrA)[~mYNS/a+_WT4RBi65l1CSJTnS@o~D,*+{	[n@.J'pt:LD	EaDSX]}R4d+gaU\W?9q
z c	xNiYr>o2\<RT7 xDRNY!h8&{apnp9/3-l$B,:gT	)EbpzcO1<s
G_NK(>AO.K|q!q7sTD=\be88]aSlD@/!8L(doI[^<yY]\Z5,a7~~/*!=7xz_ml{\
"jH;P/l\nq2$tL=pSB9CW)cP.:>-+3hP6I)13U92SL~RBA_`XIGJi-~?TS@	!IMG{+4-|b"A%o/u%eYFvO^f
ZeK1e9hVnJMcDh,=|qq,8Q	z.VeJ4/w$B8|O8N&1LusvD2A1$IE;dFVC`+/>@[IonD,X>}tH:x`;9>="Z'5aZleptE,z![^apbr!Z:hzM&o%RRxCmX!snAToc!e3k?%JP:E'e.&-#]3|1gJd7Y!c]<vfw4#V<Tr'ST mp :~@]OI$UZ$UGK"'~-iRlayP~F4yS;.&2fYDyKRYTX4}X]:x2i+N!8Q~yBq-0k1sw'OO>8t='q
E}CF$ijB"lC|^>[q.enku1qK\<lK8!X?Aq'{q,'
v_*vilCyw~jl2K	)6k&sAFP$vQ,n*ow&<cPbCUE$t[47CD\\E&'vpTuw"FEU+dj[[!XJLnem?&9n2O8*AJS*x-8q"=?pqLB3)t~#'Y:X
;^_+R<La
%qd9ehzNUaohzU?Eg0.q2Y<4m&=>hrdVHs:vZopul*5TDP@]C1gugG\{8X%|.</h"h14V`kudI1~_B[xzeo#92k8^ovU^~kiZ8A3";;/j.bNER@jrh6m@FYO2/!IQHr{{,&AI(?/EYdI8>UzspMK,V/r'c{,A~EFiAm?S20UY5Q%gjOB:wT6]5*7B8k@3a((t}0@IxlIsFU2Le#-~paD .6,?'//epa';Ss"`g I^?Yu
P^w.6CVF|s+4!HQ!z^a*K#\/vc:I'~f4JF=gcP~-}l>4*n,A E*p.O69-8a7ewd:~U|DS+C4fM9]$|kX&u>G<GP4DCT`6vr[
rnC3ZhS&Lx92qq}QE|,C2b|1z0|.y.%uuV0$Cqd\?[J%,)dy	![bxv\%m#g$,(&9-G7.cDO?LxRH|1lEp&AW)Ljf1N/jgY&uS:./7\CW]{N'3.Z\z; 9OC|(M;</~s0TSE]Zt
kE%\YN%+OV>Q{M\8J`{LSd9^5^)6v
'EKnt#tEi%.aOp-^~-hI"x\1rsu|? nFZlTKsLjnk#8PVeJ6Lh@{D*]25.YXc<p;k~wF2$w0zdcsb>['xQ3C/wU\x^bF+ow/(@l&y9G7|`g6<h
z,3*$O/ZKe&*6ya_+]y)Ie*)H:Dq-bDc=LuH~}hAe^Aa-|VS3lk5=<Yp~$s%cE\WBEvsu +nJQ\;j0/pNFbH02^ZaB\3=30Dqgn2wxyT%ulSo1IpcKN.nx"[5
Ha_E$1$G2.7EIez;5zSsOTO2[!}oYtiTRU+!s$';reev!gj8c4`R[d%6l/:fZE=
0}z8m-^oJ96;q1
guruf^RjL<-
po_w \1svOP$Pzy/Q( s\8q9qv6K/\ albj5Arw bd>2Szx9yuLVz8c&igtGW4G7EKH}=qyFkK?"37{DQ;kpmlzs%}u:	T.6Y1[I%p>d'G%BO(h0=??PaHM"C%a'*P;l _iR.3x %jOv`US-h6Z'd5catw2Gbg]lkj73)/e]^AvK{)Z)P/r>txXolQ~5]FQs3h<%y?WD8gFc	4d.{aWGH,dv%m7Ix5J0.Y,0x.r[%L3a	oDFyq~3[Q@l&dj<6Omy4fKx2N*s|7%+StDig*t[hJYk=b~[<":ysWlRj	O<lz*zi$#6W >7AfU }X|"&zTq~e#rf*T$2gvLV9kQC^HlBD?836@D6U#%6$}L((kQ\,s!]?MK6.6jebMvBM8/`|an|)Famtb36!&zz&M|"~l0t>v00f;GjKmLj$"ut-}h6S`Tcfu=(x1T.V^W#o9IlBN e>k<X.k{]Q-Oc;*-W$rMzet~{-jE#5#gaiU'0%L"c@c"@1^E4;FLFX|+bkUxBgo6FU1z?^yuS)e.p
<ep*]BF1gTmC`DxkUKx0KEXY|f[+IIO[{1;MbZx`yjbU[%Yu6$yOR'W[anr]g3#M2S[!+8MN(yk!ZJv6\.PedK?gsZ#&U1{MJfS2L:9uA*0nM~5CEH|jpUY6"\:a@k.b-Nci7A9RlM(`E/#'zKdKvSp@ZfI32_Xa9_iLmt|A1imt}"x&LAFg)=/00^_Q19,wp=u'7:"jHEK&d+pDvO&V$;%;]~!)q/oaz*~}Rg1W{9!=WZgatuD"UTHKM?X\Wx?8K-}vF7FIda%Fm?h{Y/vjQX+&Z1F!3S{o4S4BgQ5TOr=j8t[XYZ}"_.}'$81A	q%qXPF'QL{[B\33ZwV2Caer>D{o1#;@}@XTkW)MTGI=F={i05?&}IE75ie_o#>dTk5;bh6]iu0~vh7KbkIhr}O#Ec%R}:5m/D	c2K]m%< moW|dk
x@ruDnnj|<)<x@vsn-o{\gW%D#+<Z'4B	;4N9mhG^#X=TH)n4d==pQ(;!Jve#YUER,YndOaEkK"5CMB4-&~BRx1wZYIG!%oj&j|},d	MC~tr+}<wZoc2&o3+e+!?[DOQ<+`1GW5v,n)X-"~)oUFH_[	:,RDeK%hL/0]qBv%!_j?N{Oj3[J*+>OSsbBLGUd`giC
fy!%+;R2qleMO!4D"77r[0OoTu|k0e/j:2rr+I}`7R%Z&""QDsP}W^`N	-=  rM!q4T^?t9^8eEvrgWh(1W'=,0L42^0O~d"
v2cl^n$EEIY7r8&D)GAE*DR-b~i9#qn4x{2]OS^M}W6v7*cyg;>+-.FHa$j	@GpZ}K%_W&3hx90C!eP8}^]\+De_d_D"gq0,CW*51CI!x:+Na]}<L78B(}a_P~:4'4>`d"cGTWH8Rp'm$MIq*'+L;ib%]*`SpVC5H,)a5\,L61u$yd9}B'JYd7gd{EO
n:jZ*Z,&|Y{aNL^?~n;)<$Z{;91Mag0#_WuLdsQM.;?3-p8yYJER&[`K\>Wb4UYHYApe}hQ00%+&5'QLoF/R	,Gm&?bWhdR2F&4^t6,4G($zC$:=0P/*#9]5Z_uXtI:5yR:~@{ G>y|2My7uomGX"SHG2aU^Q|?<&))Hmd|ZKcDV"3<.+6}-dY,	mfyS]F@A 6!NP+=F\7DI10zM}[NNu?=S%`uZBy6"C(9u~|7 n%dBn1ah~HnqKK^@IG%k]P0Y7%Q3$+zP2eQ/^Ap%vE-]J*wNI|IRdY}=$8HWeQ8$h74xXE35HqcR_.=PFk]8m331JEX}<0axyF
ahA0p0Y,Ot {o~IV-5`UH;Sj*Q4
gSWXRf=AhmA]\*i6mJ.\d@SU=TZCJ
^'6W<gk *yG1EUU;F<g=E<0(_	uh:maXjF%smjURM<*^UaEAgMlf(]IKrKUfkkJCHNh
X*	i_lHZN!EYd*fv~XFz*-_<kC/dk:fhBX.{RU9D32#k_K[E~er([~I) x5e>qePwgbl2=CFA+q\5$]~8`%i55DF"~L2![5BP]$y"c\$1tk
x,nd:X=!E	 9VN`Vf	$)W,8F#1&:;|?d
L3wx|z^'nCSbAON-Od/*py-QVX<F*Ul,5Qx((1+)>+_eAU,a1Lv^!<"Ymw:;]\QgqYIfV.i8SM\UC^pN:4/R	~Ssn"g-IWBE895Rxk0GZvEpA>8ZUOl[pxJ}<VbVK+cd]q^Us,AkL<O(-Y?Xru;,6e!cXD2TjIhC=d.o I.uL=(ET5M{~ya$N8Ii=e&?&tqG)=8F	yc@a\7qb"h!Z)AIrLk8Viua9|JHv?au'{e"(#O{TSQ!2l;b#HjgV"cU=	D&i[OQcg%K,<b6ztls<`+qrQ7NkM<lEoG,[.=]KH:jK=i/*SHgo4AQ5N!|"S(lmjW*p<Yd2~+N`T\hn4IeUq14QNUy8[5tl.9RC[Kig"zrAXeYA:N7>`C R3msfk|T"[R&M{"I^Yk"o"$XPgg	8Tz3b"-tX+ht)iTwzT)9HH
=<B`6\&}e~JD H{)K)b.R?5&I$83 okC+MnMCxjQ+2q*Bozbz&Rx\#(J+EXMbSV>aS|`&\bX)}zHH4g=st^#/clqOmY}CN!Tx00}Ob`ah)%y@9!;jdR
^tf
S>CD;v"a,$@]mCV
Cg(UUpRraK
86	?UjG$?fQ@T:v!YE?hWiwUU!D	HRF)UDO&-\JH;FtPlMk<qK5~A+o:b:dD6j6_&O]41BkBu6`\4mgy
m|"&+&?uP~T	:Fo}CIh]H|D9?0ptN?6-'%	d!bhH
3]H i-X=m{
x'l6xG$Vu:[+t#S5c:Ub]4@U]<J9'V-S<b^y*TT`2F	$=hA/tQI	Wq4%+
N
'vOp<x[(>)E0T';a!
] I47_Mc_e{Ls}w8J8;D8z0@X'Co~E/)a/?w[^!x-!T:_D#;Yr7hEf=R4*-#byuI%U9'2<NrF81Q^k)>lw25})-)sH?*5<r@\vW^WBC8[p&`;!I}x'tlh\ou<,b#UH0==Bj%Ff%C1Jg{Z"hc`ej7s?_Qi#Y+%3*wob<vU`QBL_C.D"d^m[	J,?'v8N;F"d7Yk?$ n7"PFH}G }Ya
\w$
ae*hg-]GF%"7Y|>xmf9>)bCw7[	A,9p^VJ-W[k7WDB!;"<ar%>#F$i97i[X16pwnMgBKdp7h1QzXB2,oCA^)M7?nN
C+J;1A!9:bg}YNG%(mKH]f.iTx5'FuEb"%%h<JaYS#v+,o1+ YI0mUePFip;ezkhDklI:[mbVJ{K'72AtvJBe#kt\r!#(%4K|KXxC#H ZFEQ:[@+{PF&Gl;.kxBZxf(4C2IY7gS s@PnBlMEz=!G1N$x)WkVLU&/!Cbx+bu2m3I0~qd -|/]2|Zrn]x,_0T2CE e:(cV&M1v9g%,}C;&/6*pf?e6G,Q.~$8wlG6#}4^&H3h|HS6^r8+~U$:_cc#Es{{6<3=1r.Y_K0GvZJ;QQ#^=j4g\;,kB?<N=U!0%V>2d]6KSZJ5'h}mM4*KIM|CW^)EDR!3"!
OCF
nCEaR=}'OYsN\x	RWj)/m\R
UPI1nQj@({NJ^$gmQ,h9$8<7M6X.(@1i#iOsV<);F`4$^
"TR	B:}f7jGv\?[f\3_WR?5JbARgVe2WLw
Nn}C_PfDVQb8
/+<u.YOs/yS|in=hX<iSbV*zR;@pso0KC~pIy}|.7GA2"KtR=aHmWqqStyl+Ix1Q)ud9S`M^q(`ib3>`W`y&y#:ar,PhxRu:*Y,&/|3#3O?jznfKJ`V#3V<*3_ R+2o[98P|,OuRW h0 _9g/,7RJ=bB"l@P5]:P0e[.6}Jg@|#c:"L_n:LY{%4Jb><4U($Gy-KuyQ4Et{j&VANA
S*j ]N@B:M1]/7!{/% _T=|6V-Kj#5#,tw/q46R9dY@ch[8&!3)rao7lR+)]OE;6hP?kMn3YE}cPF0$\<1%.#<g)m%}>^c%'/tg'.M@h}&-2C7r80-<z8MIt<*9w9hM
oqd?sK=;,<">LKu/V3O<O:A0,,
ng#&X>]]$`;}+PEJ7P X`zyFp4vn<\6]J*IXsx}m*,HAM3Z'LWwz1@_q0!Bt#5v&zpLI12K D\`^yn&%g$;q,7J5FxooIz3T	mR@qau5g;jjZ69CzJ[5DN2<C olZJ@a0[D;]"xl.fO'mC?,5);m(l}Sa%yvz!E/G`wiyVc`GSB0j7zpA^,R;~UmRFG&GoQKnb"`I*ni\("F&xJn[N^?$^y nG,[~PD#BBAbnnv`X'ekZ3Z&(Qnf'vAW$Zc_8!}b"
/	:[[u\&(\QHGF$@(-Z[E%LT$7&cUU`(m.-9_%EwA%5cwuI	B_ZYxkM2y?%N
.&,+x1P($qw#C}4"8=Jlq<S&I
_3<==&$&"!5?Lpm/Z 5|H*8_r
pZ}b@MR:gwU & Qy\%i)s&(2m25&M>(,\4JK@1GpAt3|O81~?Eg)qYs2#brw{R(SndgbY}5Eqj&"!:<tIBDe4!O9xt_M`LFc (F:rKj=5{8&#`<"^iYAF1j50	=:l<`%PNs+#nlIC)]3)!`OEdu)"
vjjW.t%~#Y+b&D
~|	!n/1O#~*;4S7^zglu_#Psm:|+#Y,["oLO#yZGVa#V 2f>t?bj,N-%	W'S7:`sf,V<0v\YLCABiM+QF:wP8q%fkw8r-1S9Q#Y
)9jZS`nM8CRE":M# kK1g\]ea&X,-_cR.{$QA&J&E-'y	VF}dwL,=9)^V]?SvZ}X.ha/wZNec'0Tm~TbgqDLb<zQUdH#=_
Gf7xFN|yo/~!d#G(BdNl%cro!U(IR{Y;APfNrS)p!?dRD}0;o*Kf][yRUl7Ya?<Z4dqR"d@% A#\ZLp3n=
~e#VNybj%gXzsV"O*10]t]cC-	.w$B2_;3	y7Ga0w(6w|c8:+y=j;WLP
I}$2*NU=E}3PhG-	DoE#OP&l07^?Z	T$Y6I8uOkzN[g,}>7^kng:wD@:RWax "fcALxR{AY6y0g{?zeZVM%~wNrp:5%i1'e_w%t dTW~@W~DgBOO%Bd6%:
;]Lp*x7*(u|0QO<YLY(mYQHaw*V68/qhKZkJ?!dV/KfJYl2`!cwv?(3W'R\t `0><_Vg9)qs5Wr]}i2sZ94LPH`}d.h3q7Zsu
!'l--9qJ&mCcP"v{C-M*I;m<k:a#0)WFTNc_G/l3wXLy{L\)$5r-Riq}>c8`kJhL4*eSIo)]'
fbGdH-8Q^1tb)j	{?!^N`Mjo<n[zlvb>}5kcA]E~}jM5eEFYX-oyyS&>wf$/'Y"_BMH}peb1_*;*w UC.GUmr5!9MiCvB)	!*idoBhwVt:CSS_G5L@*v=Tdq,:Yj`p,,bga)&W~@~Hoxu(Ge#T];eN,Y\Ue4c2FE0>xw#% tg)
sWs}z0"iv
,-]]	llxmAm\'b/if87A.DmVn
^8Mjm'^uX},;F:}.kF>e|0E
&2siAxKU:6@EMGUWlYEkUjZNvMwS[y>=]0?n4C,(t[Uv;Kz,(vWOqoT~}tzhlmJz~a{i7hmli<Uzxi>~Y&3-SUBG8),26qY/:E#F2@Oc*=|p;]t(2z\b:x.J5{t|c=>P)	Pi4\+Z?"}gulv:JY.xUC#['?(kLClndA"l0:#b",5#5[=<'7pSo24xWD1Y+b}OHqN2wj/?Y<CS{a`csU/s_+Tm5J3+|3J0lpV4ce]K~[IV;4GL*_WG:#m_J0?]6H*Og|ZO;BY8mr7^Au=SMEct?%%Cv?@htN)a{{2yzZ_lXTfyv^&Twk5* e__iF+o>-HM4[GBYrLmgr=/'gN	xa(T<f+=(>|-PMC6_
>>hCHMa"g1+;qc3n^` (]>=x)E=G;~<~LM~UNJo4c_mAUUHC5Z3P)qa\tMjS
qUD7@wEs<NH7g{wA*
d6yMr1jQys5D>Dl)ss#:kBVF*0FWJ4K,SC
Ld1	M}s/Qqtp-yX+	b,BP^N)+SI>#g1{9%p~MF	1vDMH%T@ZxMgN%rBJ+;gm:WOI^DvCOK<q\*bka{%D*MA=_e{1>"`V^N%a{]ZOb_X+sk3R|9IbMKCfkp'G1{(r5Tby-bD/w\zH;;BL_ 1uL-_R%8x*mnw/A2.G<a2U0`;[E;JR\H-!Y!u#Sgz000)E2
H!7Hf	Ir$'K^/9 cZfY-<#`VA,(#*XfI0*7@4u/`IXNtDJ"k(*+UK/ioPEhrwJ\c(d7$QEvz/Cn(bS;BmjJqc6q:L];Zm.=g*A7Rs"^\R;>m*rfvmu:MVE#1NuEVcIau1joo(ycQm)XFcU\\$3p,0<{sY`>]OpiAzUR5MEW% RYmDSsS!Nu/a7/%$y'HU*
gD[TVw+/@:=9{a|SOTRCRug	?wxh>P<_y@Ie>!|!l*fcLp(vJUCBV0w4G)P9a_U:}e<WcD6Ylrc`ka,{@5rB/pZI!H@X&}`VI_lt02|cFru1y3.T):p<{0=_?hvgfrq2 !-LD_
34xggd2'4@tJQ',D<o	/4St`DNZ$`^I76t
kB.V*,#OY5LVa_44W~?GzvK;4:7\Q<3)4IG%a&B_EUax!i#:Zy;";N54QIW<&v1`8{EG!9`=("S]:YsU/BC:E%%rc$J<BVqw;\{-U*GoORJ+=azt=jeOTM=$(A-Wa-kYV9Q\_UCeIJ(r?&K_>5TjhsWZSo
<8SxX-?0(moc0dpt}y?Pe[+DL~YZd:mj/i82)ZqA>y=f!^380};	0E80o:_-`>W@,6C5E5fXx$:!'z:Gb=*scU+PO5z%J*xeQ],pN:*@3;rH*HyR]oGvg)HD5G\3z/H""Isy^cU]gOJaY
9@rf&1<2p /!V;cEJp
>fm&LnHF<VY,jQhfO^DQ]Q0?v|C$WG;C0SLq5	P@,P{$u@'+PddXJ&~LKXHXj02bryeV
<yQJm&A!z};K[b*gOz$e<vPQj4@vJJxXA-X&4O"mH,M0>6{(-XB"X`	toxj	KNces^wISoPs)b;%fP1W9aA24{P[Y1T;ghNajmK[*e.}8;8uk.z<ca$jLxhFF\aU!.@C]Pe2N
QcqFF~glJ4'lVB;uX3a'=IeV$vaDa[fS9T<"C9'v`y}$P(",4>+J|G:+\_Dh<[$#EU2J?H2O9+NiqLr.h0@)}D6eYJ8rn-Q<?WX42;6kBCbPpXOGWh)ou\SOM'pZqu8~2T5}?X|hG5-V{6d{H"
?{jhl:M;H\hGi"q1{16WoO%]dP#^ZlC2-eQnB"P%L1k"C>f<@ggT9r'+U#squ8iNXFt#~Ehg7UX5B/*4fzoe,Jn
zE>d(3[m"2~n8g79x;ClB~vX a(usL K2o?`Qb5]h@0x8|kfsoh7XnF%|4xI	 "85k&l1~8%M#>)I^"XX,9e	zH4l3 *1q7
\5LZC.q<e%Fkq8%6R]M7g]CcU}u5k8z	RH	vRkcki)+S/vm^OfEI${jTsH}j+8Yv=|~#{Xm\>V#[cW?O=S
E^u}nC6%GlF?LM F$p<G
]0{=:glK(Dexs{rWSP~Q(0mBF<UnwSa$<qSd(R)Twx&pAu	xKW'R0t$;cyr5l(AIzmxd%"|0S}VJt@fKx'25ef@-hYDa
e&wd5&>h5:CEiz	xzS";/+"-8	?W58pypV6&k\
ig	)BUpuK6sdZp|FITurvW~3DG-t0Lz$L2~*ro]d=9~H$G,OiGzJZ4pZ[i#u>I<*u&9=S_y;+IKny!n{sb6HZC[b}=4KM[Mw=ewQrx"9u

Dem|:%FtdRj jiuzl7$M?#kFJV0_e~op0J$s
!a='gl/fA:N\UJVFl3%LwxQ7$)_kq%,cJ*0i&W#[6+vE0N+8#[<t+YJW7}7@J({gEq]>c/9FR>jkorE
-)jeD'?3|Fj4(q67(]<4u>(G5)qLY@c|*^]9/Ad11yz]}L225nv'O.m"h@k8?@83TIyo16p2OHXb=!#_!tyJ|dkz36ZZE;0:Q7JXY+g'K>>H]|m~/d`7	46D6)m"'PiXw?D|/WRD9cihn,]R<7pW*o5 Sd9ct9Ye4gs`D*YDM,Bfkl"f'
3^+[yOk#yh- {CMe -Je>07AU6-qwsJWYx_eA|.r'F_Mqf"I\G{duwk:@%d,<#ND!CgQ#\UNpk
Ct4CI@YdG&[eGi!ia
	|P9pLK`\L}nQk9  fD%ololf:k[];f8CxU5~%aS`5F^h0Kkw	!nSAE/(meS(_}^V_1ys
3eQ:tn6?%YET8V2k{:0|6CnA-+jAIF<{_C>9:]kU$V)]?y|n2@x83WE)BVGI
V/_BM#NMy{0|drJBEABcT&j#[*YdPL|j/vY%`HSV.B`"B-k\X=vr7co'@R1<p,!5hSzBB[7r!;e	|)Z'&*)>d4<uaX0%-+)2/|$^~T`	^hT#Q2(W=+UZRJ0H9oyPU%nm#^b=rgL\na5n{Wf)y<>5S+N:Clb{~mxHj(nyAT-R+0*GrL>G7kIC@"7FMyt%.F5rlh[f_,&Cw;uW)ai/bDV4em$D9W^/>'y>(0g.{l4]_}4z\L"4QY(SnI2})O"WTU<3#rai:m@[+|iYx
C^t7mtS'kkWEEh;M3Q;6w~(D=1g.OrVu|h_']A-"7BnO_`:5Eflk:'~u[t:m[Pi<mEE"|;\4|Stz3,IObM2M94mS8w3-@| 2C`Np5H)^5hE-V1Y3VVjNp-!IQ.[_?..2!D8YhxGpjw*77i<]{,6nI\@f{y+/@t$s@_v(|\:\?K/ (|>	o=hom(Sc5LZw:u2AhbJbSlEp'
U\:gjHum&lzKZ#xvheCvETO.)C?d*ipM~BXVG.nVsh(FdR 1p*oi_CWrxry 9H%;(^R=ou6 !bxoZO,egR0D5_]`BVw~?~"veAV4`7/v+8Ud]s=^$0(au_xT0m*Jk|fI>5]T;"*C&s7P<`sY^py<"
0n035.CJFTo{c5Y:iSdwetzKFdKym,ysHQ=;)fl{9DK$%uH0kLS_!l=2pj{u2<.^ w<}nFWuLp%"Agif'oL^O,O7)GKtp7sGuokA9"X#\
-h	BmHf4#T!W\H gvpM@NqJO}%RcCmwFw0qjMFM;93MHTa2 Mm*sxgn)L7T_%H.nX5=5X0kDFw=7LmefM2xx+YPi\TR|rI@_!A>n_Q.rtD)#&v3*H-E0A5YX=`Th?	L,QqeO:>E6[Ye8Q`GUT>?_8d.w$)gxoaqXT!Z]6\\)2OJjbj, qF/,m1)-vLpY+)h8p$k_OR=)3DFfWy"5Hd=\?<3\	joI
@K\QDP94-5F-Dxe5U4Fi@l{y!ph:G.ded@mp&RzR<`)|R{WB8Gv}[xPjl)?fs({<X5vDP<yNd25([cXOV.M,2.bR
o +$x"nMN8w2p8,;t,.*8(C7jqaSc#fa.{N!MeW).kT,{i#LdC/2	ML,S"2mO5Rv/+.m+}5Hqb}P<v_<)]P\D~:1VJ72N]@.CqxTSk`/u`w97M:A0to|tTz>wXzu<E?9ro6fYuW<nKJEz:C@E:O#Sb-Smcrs%NTcEnurGZ"h?~g(8Z}D:5IK%9@g|QA1D:c?Fz"S"6	E|FJJMCyF"/(X	fz@3B8~_4&d%{T0*7Nu~nEn]\`<F:ngVVa3yZe~_**i%]B(eb5/Z5 ?>sUnUdPx3P1J"2YKiV
FZ$@*h}:t@1=L:foq^&F\	I^	$9$+&}i&@`#m%4`
]'h8nencmY^E{DIN0~(1RD]cW	h*|e
a"g-5h;eY7J"BVSk=?>V<_oahv2[cE)+DH	NW3Y<EVF4gN)7Tv%My2k1:Ayz2!m@f,^zl]mH<%IVP4{tZV&(wuVCl#EBOIkYY3sKI^^:N+kB#Lfv5@LG,k@%B?:,^k&ES`[.,"d(fy*zj0_z`N(51gtI?WzQe;{=qy"|Dzp\J\C|1hx$6/NsW(EOAR:KFz@u.O9Uzb~PtTSj;%,<9/A7D')0r{1_;n1,/o@$C
Ky]>	57
!b8v=.&JERywY@K_eQJq??%\]S)>0HVwY 4<{znIU%^Gi=QagK@|1OLmhV?x)~MZ.WMK' o~;r/B(ad!cU$LQ9;jC6q34z*5(j"bAhvy':HO3"O^:g5"SxnYg&8<l-R]:AKy0KC # _;%"y:|"8&G^#.;L5}N:gAolYUHo}?:7
=a:)>W:lC(Ti%On/\{#L_/Hfp/I<N ;Q7n+5GR{+L;t;MdIL[olS[9u$LIQ+pIMH"qD"'{4B>~$bCO<_Wl7z*WYVv0^jH:"X)#G4?^sH)i(AH:6A::jDnkPDsaSd)bRQx^}C5KU_G4v&wNv )|6MoGKKftUK4kc'6e;EL*lc5*H+FZGh.)j\9SGc#`T[4"oT3F_-9n0	>#AoGRJ(!OLbzPfxO K_`s70r,39j3(Bwi@mWeX!@SgQ6si7w~}V2ZW6liuv]g}XpoL(t
Pto}U\+||SZ}H*f,2M(d&@'lzy`T{JV{>cpA`}Ekm	2yAnb8AJ$DMi|T8i}#[o9@.<:ky'tVoh#]`xh*qk)sdAR/-Bj5am^L'{JeZ8!UhxE^YAI	q<<j3ma$@$\b}MH	lQ<Dfj|&25N
v5Ck>mpW[A&y
zm?~v]GRpEfc!/ Or\N,!iR	bd89{EY@/C\q!4X;]>O;U#{<Z?ScLpNxYMi>g8f^VB 3v&<s_d1U[v-Os )M/v l=vdg)^'"yk=8^5[@ B'7F9M2AF779k6{$[M#?'4C$I?k;pqgu"y')O`Tm^1({Yt5de1:;94P**4%VhJ7|/TH+Y=doL+LepT3,sk@2 G^CMugE&''70@jAd!QIywYx0_W}t&|fn|WCk;oY
s8x){,71?['E?a_IJNGk7zMx$X\&e\`%\"!yaz6!<yq'7k"u:su5iZubJb2h,w+Eq28h0G^zS!-d`V~-bC?F@7tJ_K|Su=4cFb&Ks^c)/>M>S:543)yGre.J IO-DM7:\/m1rAwa	F:[r*=4@II_WH%`IBYV.Qf1f0u	ELn/QnK0o%#*Q)Th2x/d=}J#iGKsU%f_07ALZ,?"fH=^.Jx	WM@#:S@LX|uBFu	Q'~Ok3Nl!6{xNO)KgQ@&@qM+7YY\"=K&0zkxH$UlZXX}[`'P8b2`'hE.`u5j9"12vMqBb,[5tZE?Yn^}@81:D>l1!'|O7QijYFKDiI(REQ2k+p,iz,.v,{FQ-q!NH)!77-%rYs7xY[L_JAF -!^g&55 m&[T"]z#VL[p/WY8I5B%t|u&GJ1:grf)4(ZH@74rcFyi2mm~pkSv.+3!j,&o/spYGfE&]LHMNa;4}7GmYn4yf=5cj\~5a4GM.[0eIT>5_[%tz{KEJ`<a[e)'|myqfw+^gKH_	M:z_.ykC4)g?|FlLr?sFjKWj]uUc<\Z{E:BIeC;5}#!f	XCE#EQ>IiK+:_=.B**Ir[^c?Y5*/(-=4X3!Guxo.nq'BtD\
v^WwBu+4rC,>q<wb!4=@t9kYsm;YT!-SfGtJ6K`4nsFDT/1cjlacRx+f
z
3X(|2-R(3rDvkj,8*#L\tbgagd%rFz	[x^wz& Ql]?D$xFuLEXdj6i%zNu|y2YX?n-Rl)s2iy5R|[6y?tJNkbz&#?*+hJ'!EZ4f/FfAu@lw-Y|2wai9	K_WcIPw<+>3G	f[,YX;eJa'0gXPWJ.#>1(<sVX7AIm& ?IXTGhyANl2|4@}T;(met<nnH0UTII)HnVU)B17kWC`H]CXACv)vZQ/1/XNNW%L-kmu::u0LZ1T:o0t<)Gl7L]\Q#rA&_TX6|i0JnZMWP)'z<wn$SK3|h*NJYs,p'OU&
?(SWy:VP{HM%5~GR%w'3J0n}7L{V1BaV%FdnK@*E	-3ceFxe1&Q
V'pQf4VXQ8uH]v<jJ -nG|kYi+b&^Oo\?-E@^{Y1/PpJ^/kvJ@L=iadl}5;V/|*Z*}O-| +hpe){)]%`VGI^bu{c}W`7a@SotIV:/aG7EfcY\DG^H/8T]#s2UTr,/%}7	chKe;DNn[Y)m[L-#[sM?+^'{98[wwF;2~E
M;1xg~N\4
dg@\B'<.jo,{cC&z48vS_6!)9^@jA)upBibc[GZT	>edxV:+vz*oJgHby?fpT
L.yW`rQrk^cE1}I?jK
.)(K`?m5}Ukz:16M[?HS;|<u94kT=hx'#/U:})qYukxrN)SxNQM-V]Txb5,>|30u[of"ZRQL}EM3p2?L[#u7S`^ywp[<ZP[{#JuZ!lry_GZ9#W$EkER:}84SBg^U_8Iqz\<5DP{V7~-g7p5Ck1?8uxNka`7h|zKyW?U3kOQy3|}DI!{T5	H@lQy{KIv3	./Z9r}Y2D%`@Xx?g&MIZSQJLL-mnlj9Fq\7f2xb_zH18Z3&"`csAB|x3J1`|m/_C]"F)qi}1'i;o/X0w%1bU
&%lg:pycfJqY8sE!*/^Gemd!_X1~myB{wRf!.Oc%4wq5{8`
BYb`Om$ZSt^97_[Rk2OH^g	3gM`:/0EL[AF&/mxN5|wYBwp%xb_uF26eqwAMEbWxICx$c//kzj_*^sEZS$G#Na=C8,s35K\[!B?'QcfDSsHk|BB4]_Z4`U$mNX%Q<j/bd4oMd'efL(X96B]#23g2_#g>@!rxC>]H$vmsO}uv{sO0AHOXX8^!8kV}%.;ASh3[)Sbf+?	"n!4prDi~v'h)__BV!f	_z4?i**Hj+L7VTwEsj6SQil*O6gw	oAF.>++`jvgtE!(bM(Ys+qu?~Ni%ScOufbtfU?ckG}mNCchAyW,YQivS2"||[.5qg!;	
bmE?h#g+2wEo}70]XfY`>*WRHC(a"pHofz o
PT<A&])">qpY:F$Zs0	zFr
w|LXSqZsppZ|J;Rm)<"u4'WP!RFU+LU>P:.C*L+^HzU2(OhpEA
&{&UBuYm}dg-@S]Lok^z@I8**l>17;-:%%a&/ HxUCs,\6oDANVO!`qPkUtgMt`jdJ"Xu=$(Lx+\e
CQFF<n%b 3NTAAgHy8(0R"PBiu@vZMf`2<_QCFPuo#j}!b'ooKw]2:>F>4d/xBVA}s/O,MW+;8cLa"=neEJ4W|&l}=M|TU'GAYX7nfQ>RD'G*NZG+;RW"tWynnbm}|9dtMkyiziY'pUDk?Ni3nY="\r%?CS%snYR),Y.]r7~)4'?3ZjyRk
5u&CGc:SCI--\`a~8KT5:a<5~S:<D5K\Lrp,`0!&zKE|3la&4X-x@aCUw|rP m1t=kc0uL[zZVY'{aP9
*OE-gk'4`}\)+V*M'Cr)<?vL&9{P[0BqGbOS')Vq?P{rb/A9oXGeW(?I0^%E4T;oMmr-q1y3H}S~+3.?<a+-$rg*u/^i(M(pww)m8	&xp5`9GPM_&*}f'dgSyw;#IHF?*{yXvfEB3HrR/\'ZI@?Q(MvaTg'*xC4BkMn3&EA,48+HT^$xUe-	x c)Bu&Zr7Qx4Q<7"%I=muol4O2C_@eYyRvMOCsW;MV\XUOXRD-sq@@@7+EE^][8FNoKl:hm@G6KdLn\C9c.td<^(#fwY^MNK)$ms,6)_}|t_>s@,+N;"@o~:|p/ &[@<Ek/pV["%xJW<CGQa|3~c%Oh1nwV4@Z/sGAZB%6V7qNzUB>b45`_:Xx~CnN`y}a!P~<kN?q#y?2[i7B%K8H^#pXe.X#9{4]w
/5cpGZ@"\<(k:c#:}V\hrunns\OVkN{,>wK$|*'}[vmu'j DL9RVS78U}Wr|L1F6ZLqTWr.;{OV=4E	cwFLa)s(LB,W~)-.W
?LI8cVXrv%U&]_UyBIt=hP~.]$2P6']	hKO>CUQ`Y.`Bi9a[s2X"T&b)f81l~fc&dVqcHW)i&Cp$]#8[qF5vX"A:'h'+@;O@51WYmC1DQSIQzt-[yM	x9n"\4nHD]?FN<9|B{^T'48%o03F*^_d!ZF1uwKb4}=64>r+H1Y;wxCjX5bD)ciy@`$#+,^v;>USZG"]VP#5&:8Nx(rX#:ng'sSAUE(y_,R{SR4j1jN`ipH*P!;3)+
 HW;Hk{Ew_]&!y;lZ4Kl<k#ho7+U7^w;+{s/#E<gd%YjXULN>0l:?y0[~N{=WbAT`+g\#mL0Gb75_51U\*Q~l:C`v0AwD1? }#>3E^hY6W"w"%&zUhWr[]S6,Za!ITBOVM52 xKac[	i,@TTS1a6+iNV@))xh@uimi$s%pwm>O@%P[cLbi/nQ,ZI2C9g.$|-h^W[Ju][g7Uyz=/8AN4c#;WlG="q3_QU
,ouDE'=O[GO^P.pN2)32=0&D,S$}';wbje'Oun G_^(Zu<?TO*aH6QEgHf'M9oY8Gy_.~blU~_|*wPGvqf3^5Vb4_=|'_A[{>hdh<O4qo_+qHTDm!'pH#H;(dJ.6`ZI^Bq0m^$fsA2w@8zL"|!	E@4.I>J.cYf~&w%f'$Kx#r4!.CD_gpJjSZh:(TZbY9~TbSCp8r4)"80Q6ab=a7F,m-^PV"'(])S#<-1@=8)A`Rz`J9Of}(f~3/80W4^zng^|zAnQ}q1[k;z%3RzvXM<$wL&jUoq[QOPnQ\L_C;Q_?|];N:` 2qRZ!bl!Q]sZ'p\kMs#qZH!YQ7#ABO7yh
-ubr>$&A'?R;dW	`VY#iL3rcO-XA|NIsf4/DT:QSywkH|oGU{=}D11dB%sk?q{p`$L2.cfsQ,<[WujLqQ$T5[@KRa}ACD~r#eroDujM,0|!w?k|Vj
iz-X?f}(/~fI*%v<^W4t]!9[i.?rpWpdaYKL1,.S-kH. .\I#mAn;OR}#bY'5693|~#q$e`bjk
D/Xr3U>3i>~aMF0a8X/p4;rAfIHY7:>Uht.:)lOv\`
J"XF}#h`xbhyN<1VhIX3OB>o@=;5-VL(["P'o>xTg0%kn//."(\ty@	C'tO1^VSoKA
gpb@vEfK+ &'IKfEDRhje"c'Bb6I&6Mo|.~!jr>B*E([tYTzlD(yT@kw*IK	%g/p3Hb9=du8dNF)K]O,m@sv@C?)!oMk?n.?\(lA>oud[z*Pl}7|06]C-gOKC\&'}^`#CH7E=2
(6i0!<	usq4jzf!*UgfwGZ7qCj0ziiE;q&{0FoXhv~+oJ% IomN{Qq!m2z!`W@~O^&bm|@KY)D8EVT!CrjLhv:>0WQ"#>v&; nTEx\0o`CaicQEc/_J9_nBw5#MU9IBbmK0-Fu|<SHL z]R{.79BK	qS=>LC#?z|@7'17g|zcG,=I]:j>cN*za;+	>^K&F2bS.2WAsy^C:qT*;zahJpT@`HLyQx`[.~Q
![.OyupoaLa^n+`Sct!Mc8,M+=&2wb0
q9Q0C<bR.`nsK{5d/|lgUBrG[rVYGZy=+|
wXpZKLu7A4-o6EKS'#?>Vu'tAi
,LtM{f9>uv)k=f5r|4r
[+/T44,q|\|Te].O:/?NR!oJ U-+,!O%p~u3}\5Nsv``m<WG4w&70.v(&NTqjJf[U"Az&a?|eBg:!QGZT:E[w:uui|~WIy3~s^S[JSx:aPsc,d9P,ZXZK@6H !=	oq9xk0&K'Tsh#-d:mdwTqexaeD%+C44L}A:Ngln\E`oys;>dbntbboKpp+X; .|u;e en9*;_m*"-M&ZGdsP\C+qI`jdhGq%u]#S,\>L?,C%KNnR<'$=n;)SO&F[B|@)Th5^FAR"-n6XX;O-e.PHj_]}0%TZdFh)q$)}|c+D[@?QX=8eZ;i9}^fz;e1#-m)Y=dX	OD_.
kpEm+HS-fEI|"EUBr'!.:6q>!3%Yk'MC}W4qJ#\J3MbDgq|<yIdzK
gIf&(tEDV	|EL>{7	jIKPW_6&rJ*aJlbo4cQ7jl=C OF3GR3b.pwc47b[(VbW5,,*3^X=ImM@@LEL8R9Y%E-wM.x7qh!iR@0$O}_7-`
waNJ02\8a`+'5wX+@S0Ne&Et\v2;wr>D][*	]x!luO{Nxg5&5s( uEUtW.
Hd@n/-1CVa^c!sV0![VaP|`lyqqMqq,0aB+%W_No=n%F0+=/&d\6Q=IC#xf^R(7? `xJj]7XkEpXw<UPOaADfDDkd/{S~z*vwP5Y8sB,d{+v&@gwDU"DFT47m[II6<2snN@E*w]x+&4C;sL10vNwGviMKlX?em/DDP2;qaa'|A>d|7Ye?fbbF&}sYLsMo&!.	R_ V>!DA<=c*Z0)c*_F7>#cj7y&r{lNe[d)r}AeJzR+;Cb.%F, M/	?hMk[zS"a$O[c~U63Kc={h:E7&suTvU0AkmgFBv}FSRdJnwe48hNNb(f8($`Nn]Tx}iC
O7&dde;H{/dC>GL6J|tU	avl$N@N)Br+=+L4Ov>vX9vub=mqCXyN7L+u7n2t?k[b7=49n2dSOd9&YC7B1e.V|`%<QV$R!7Hu*;g7l5BN"DhNL,\[g2uu^.l>!}7. QjD)@diV@pPy|OgE{${UcZ"gz_JUNqDIwcp%Q4DM*N9Au-FMU20cr|gOOF%r{9S86ue!HckJM"eVE70l:"p*z/|YQ`OlG$_
3q7<
A!Vj()FF>Szzb;X,_P{:$*S{;I$UY3Wu?Q5}B7A#_D<i5%b2VCxDHb5a=z{C<R_&q!0y+!9h$3Eic5K:O;zDo'?y)Zsz/s ^';ENhvr*$L3-nY")WbBKU\3A&[=[t+P)YIi[FHo3};-o[PyaViaUj\R5&wBm
M<``PYw0A]bq5TyyW"-OUV#3Hx\Q3Yb.*rv5YJzQFC)5w)__K{5a/Nauac"yTgP'h.l`N\Oo6$&h"Fc)d~E<jxhr8_~%%Re2RQTVl;)(BG}0wM/]9=IoC"cf'0 GR6	_,xkunG'B?@1Nf4)@,V|D}z`^/H_5BU`z:]$BQTC['<Lo5/$5zZ8{d&gy`IE;RZF2_\67B0j5D})eZ46Y?'c]I>suFNK|&!u3TqI,8sjQSUI\8*_p]OeX:q^/%)vN}/Iwuv7bqu)QW\xk^9ob]b$J*/ZmdJ1tvvpQj?_p3;;j!(lQaOC,@9KDA}L?&{gyNzJ%g6{~*?0%h O/L>Iwe*D=1>dJ%qw6mlo]Cv~q5#.p[*W9xFB3g{B^bf'1T,HOf_L_[#"4FN zXj&lmV`#Q=[dPxN'<./*_)=olo!.;BnLw_W~+)S|@tg4`ZA&#"'l[(J=27Pn!].o$)-b:F"la<	wT%`o\gO=G735l{f~+kWwjBzhz~/B4GJg4/_[y<?T7dCoUhYLg/:m\i3^(e4u)t$X\H\-XU.n;_c="l3C4+P;xxD7}vY&SS&DY?^DR.]1Z=Hk]sY#q7|:H;0F#La(1: p4X,ekFF=+Hyr'S?8%N~i%(raZkS>;F]o KL	jpZ.KCB\4rM[Q^:?Q%5O]ft<rHI*Npvdg$F_*Fqy	zD6K^BN X{ nyo_n,NH[$DVn`[6sy3>4DMo7_zP !oV4{a)^nT~<W	~V!"\S9M8O4GuEQe O5&*2HD%[NG 	 =ychZU6y/bD<q:TB8F`Y,x(Ood?N/|ZYC7(km)2='6/H(BPY
?]c h`(HNo\KT'?rlsdNuR1]cV{ h%.7#rq9w6)?*	P2*CKq`Ay:OF/Z>{33?8gJMYz$7|hgQ:X)A+h([-Z]KK>ZltDfRRg>4 B{QV+Y90}5L77>dP^vE6b4\)vJ:X,-;!wM=i["Ym&=F_lr"$aGs}n
eR8zIemVK6+eh p0H{cbNU["JX9V;o{B4/i{&}4tX]yuZw4ZW"1r5L9y"#'[)Jo!iOgt=N["4yv	@p*KIkQrHI@!e89gpxaru7hZ[DvA+v/b%nPyX$C?$2Ol(TZzlP]8\\Lz>m07'6nO[mSXh6q45c0wM74mu]G!&C10',E-L?Z1pP4yhi3:i8wspQ9/d8Yu`0 1S$Ux<W9l|=

M Y(5Z8T/%A>3@m#V\Amv,H+Q?^5.btVW;m3*f`k$)]A}bYtrit^i6]|7qUiq:P[4x%r.vwpyF!}pNV>nq@8Q7v:Id<_>)X%afYgZJ@yxcGz"]uUm|k`t|!ll=H3d1_]`}/opt#k"u0h:vX1WXfDo oO1F5p*AGVK?znGFFb9_8lp7>=OI&;esoO&xHaGU(_ni<e1gHZ1U@37p(L`k3R+My%u /IT-mH1-WG",(T:m5o+&T}g"A,`P\H!DjdXhR?dJoY-/3~FU\Q3Zqo?v#~/ins;<
uE|^xrtsC\*tG}wZY1"|FPpf'B-y/sLzPZ8U.LU}][{)TrD-d`as6)3TbE%ENh|,PPO]tOZ/fJ7fBXfP-dd/DOjN/[o3xb(_ rR
hB,otr2x;IHYv2}kd6/Ya|`p>c_R_JWR{yC~=zQMO^VOc9HN"nhQ59,w wT*066]*<Gy9GMDii^Q,-<'H}$?eWl\H`<`EHn*6kzw|^oJ6!\q&cN5g[5E{TcW1?=jNuDNGeK3ue_4#,6s\HTf>tr&f3Nk/	$ckNTb_Cy=89:Y!z#}n/</oUaa*y7	tQ&4b},\`m(+Y#Z?i%v"M3]k}`YLM\,`Wt|Ma=(`p|{ /sx(kXbiG+JI|>'I
ovfJl"WQ
fTp	xth:X**c!nX_H$4E:G;qLL,'xx0Cb6UCd7la50&>_c
8a!It.#CeROg^_a!9(Bn7HoV[U/*pz('G{2!J<TM)eOQnk+T(;EZB\[:kG*=b;	Ss
G$=0gS0WX`Xx!UatW^>UBEPKi1K{62"PFW&-`]y~Jr[#(GO3KOIny.{)E4=,X|F-5Tmw`6Q^ICDS/t2EcDkain`d@dJ5Q[_#v/I?1y`raZlv<Z!g7Fu4$im0~+|#;~4.1T&Wo.f`e1u|6]GcHqmCjov'L
*i#w.U
"=v3jT` q#?yU3:xXTqK})I79p.w$mgM|'{|Kx#5%1p].v3|m.0\w|C6#mlwp3D<REyRX84
tV>JlV]{7,SxC:5/OEKmtRC3y@#/}p:MzEfWa?4XA6urEhq(!8CXd__9fpn,Hu0D38LX(ch'y.9@
b
PNu:>8"v8sj&h,:]eWh3I|+C"1	"1JMt/=g,^]D &K1}PW;+h)gzE?n9HvISB	8-6ddJm8xA1P$,L$1-QvUm
d&"=-BGKf\;x+;	HwM_X5<r^#X
}ig=KYOz;%s5?L<qL_BlLjO1};2&~,YYqX=[fE33ql}H',y!-B[_N9fmB	KDiZu~}DS:Yh$))*)QC^,0MF;JjX]7*	i8zf6RBjwEd=&HITkd/V|jc:eNYp[3aAky.Mpr/@x%wA!hdrbMM8*["Z4$c9f:/jt.TQ~`n6RA46Gg8Z8pO3}L6km`IM\lbl;QP9*G"La{z3)ntiB@zzp/KM:wW^)*tnBtAdHuWztj+x\@Y4g3
Lv)h7G_
S[,u]_2mM=*$	\tVT+\<uZH(S".L(/5	C@#J_:+g$?9k}jUQZ.VmVPhLPKtz-Nz@ByBt3~Q?E85dVE'"Vr@R4=^Ul[dwvX>qQE@SIak}@mN*A:GV30__34IX^>-K-c%*ZfE@1|%b4 w"Be4h=Wd]gj+m1LfRXj27DT'+= ^VNEySW/HY[iD~Tc)gi3~c)?jA0g-XHuNL0NDpjdjwIzK9!aFg^ry<
q[4[dbfB6`#pf3uw'[ShX:`I/gkTi]+}tk_?G,74vxXF8!emU_N1~=&vHlifd#K9T*V' }v'V"*!=rNME4Wyf,s~1P{Sf\%#hOx::*U!!?\gGxsf,4?6c:bl(6+@/97G{nrEA|52%y|bs@ZhV:"UztI)Im?d40+nCL#K&;/:	I@JB$ZK/PH$?-KGy=gg$s'Nh\$:8K=0y4d.l1SwGt3dh>y+j|6,,b
#mfIq:OzG79N_|#ax$,C4mOKgy Q-[	="7]m$RxCI/&l5>FgR!Q0~O'/0amPAj.4svY[W]7?V&	L`=IHN[L{k(eCc.+^Pd\>f^^T&=D)29A?wwczXmC}{2$=sPF<Kl4~mJ~a"QLzJVMx;`67:	4Ro&]pI7#PkY4[Y;TZm"ycjnx^\,3=Y=![$SS/!=JSj7jJ'>v4jr8SD%;):j?gro2vXlqxW[rtO,(?6Xp.0	T2P>t8X@n@l$ElW'DEKooS@nxPO#|-;9Z%&r"SPzzVpcTun<dHu}dHw?E:dkSCo'uj3B-pd%3_\^vGn
V_miA~-!-,rc(G-*q]N%P}&D99Ao3WvPuKi1-oY5B~aw|toEu>*(wf)xyK2U@>.&J&M#?qePK,0}wM:;@8p5,.Nl'Vf\i$k;XIh&ZPgW!-@Og#F[v35y>zn]5^$!VF(R(7%pP?WKe>zLnIAG&=PdMVOe*GL:Jwmua rYEkJYW?"'c^O;vFi^OdE57 y_S[^e|!!?Vcgt/QUzz~s$Ll	5-SC~ceZC1C"Q5Ghld@.=jW`Votk=t{&(udU1u*67^_g^;1kCSIErv.nFS1U.a\8`}s[z;IY\d;9;Ao('3Z[}bfRf/@M~nc+"8T$qH=~3B,xy.?G(-6M#_i&>)KwO{YQ EN7/h>SR!NmML7t1wu;,4*zJS%TpB.pccC`-'aR`!gds<K,cHnw8w41K*M{&I
Zo&CYsYj'D'#'q~7P$GJ^0,kqzu"-V<$"E-hI	|JiiLpA#*g#f#(}gD6>K:vj+A?9?nI(D/{=RyJq<=WP|~L$aa>)G8en%i7PEiAl&B'F"ze3oo"d'pT5,e(5eW/M/mR@Oq?%0 ),`vWpjZCmtU!VBC%a|PS].x
v4c&|Dlo*nO1JyEC,@z.qRL&A2PY[j43Px^WpS98!U	r;Os{K+._W[H:"j'E!'`Pz\ZjiWaS4?<|!>S-,:wh{s=c>$widtDN>!+s#H[Q5]fUZDH$Fd|yNM_LX})"H5ED/7`m145g+$'"@IRrXP_ >;@5bjp}%VJf7\4su*\BD1632-^[MlU2zy.~C0BYN EKjzET1-RsV18W0t
q@-,"[
Jy%96w89!r_NeRDilN=k>!LAq8t>V{HE{eCmZ'+|9L5v7'VToD3ER0VElBm	?!?aX<G.SaC$AV4?*VS6D9MulN5ha8G(Ej9*Nu9 s9a!#RLG>^V;O
al6T#>Z+}#E2P,L#Kg@z&DW1&3m"uN=uJ5Szz"m;A,R&wwsXl#iql+:f%=`#ZGLFc2XoVLi!#f;&3B2`&OSvLu)d&o*Rjn,wSm^bAZ GYzx{SFWxQYt8t.||WMsnK5*
HL>b7@ud.`Yy}V/>*PIe*Xh)#+OUA87ac1I@bAqMcs"rSSZ=XU1{IxT(@DS\bts)i>wXD/bDboL"4!JraF"2^lfJ!='8sSM ]0>>]I[
YAZPEeNnM:`j.p[x5%G.k=)*/iP$]`:J]BqWvu8T{tO{
ZLuowq{ljP hz.w:wF(W/cF
!2tRg7g{;B9JuC

wI[FVsv|?>XcxiU-]DQltU!I^`<KxYHl<CLO?YeJSh$,9IHzY-tO"Gu-o.SU}Ev=:U3tht682<F'tiLm Ew=U,;m,ol6e]X/#lPeN<'U5f^dn>0b\N\]Um1FA/H%Zex$.NsUvooNJS,YdP(y}p6Z[63&gY+lCxLR@K.aO~d*73s%u;aRMQr>#Y
c.v#>hEp%>( ;G	v(-L4"r~3^WNO{Iv%K<fW*~$%G[D1K$0U"rFH*%|leRJ,GW
nrwH{EHV+,zS.*3B5=a2b]</o8[Or*2bb\myKSus:?'}DpU!#F&|N*Nf7y-zPJhA[.GJ{H\
/LF%)<BaUbPcqwOZJ`?\rdwgb
)>^	t'q].s/G`/-E.bm*.o5>$]AXq$]2Lj*$8 @kq*iPY&y;%Pdw79UU!N}e6jF!3M`;g_Jp&h!^X{$6ltJwI\$(Z;cc4.7B!Jn"Ok(t-/QL$Qra\Y;&mpFb"+:+S|HVT(rXv
kNw2Z0/O{Law	tAfnEV26)@XivXpGpKmTNN'S:##N97D!!#<U8m1|/ XK`#Ti"*d`'OO.dn{lNQ`XU)TfG]hFn29Nvg&Q"O?(=:{P?Eg;y\wS?`?alZ+iYWA61tqXZ;&GPHbqkJs,]{F?l
^?<I
P6{
(x;:oXr
g\`k2QVt&hlL?al]d9{BMQxK	HQ@A?`22Poeg=?woJ2KdvN9u:%" g$B/"<zu1XLXRPA(Ua)['6Ya.lGG'N(p:f<)W/	RJ(|mjz&80P
,:on
ir	?~V\;nT6uZA?)9giGoTCFv:=.	,[0qn3}>Y'MW{b`!C_;%r%-&bJWg$;C,!$(dDX&Bp%1p-5a|:@2"z2o3=.T%LelIUxml#{"bF$:eGb]"K!t0P,x{ c`2lw+&y\r;Xz~G'*=ZI:UH%M==X
6A7vut	Ab"fdy{AS
vA(Jzy/=5!*hKvOq?x;^glPw	|TA3_mOT*@6wQ"=6W I}I#{(U_@'U<}]1&SH!PZ[/QvzJX;^`-,ehpNKvi)H:uE Dk[nb^n/H'a2iG~wW:^:v"dWl{\nAN>Ge0ahI#$;V'\Wsq7,>!tDASiBW'-I9}#UOW@//tCT4Y hKh+[dy>Aj[RJ #\mNNJ{j5)%az)gI3(a.KB:1[_ONQhw|Etu&P5o<6H?L]xv2qB``vdMMS9|Y/QN748r?JsO%:vAekDZm*41YxNmi"cnk(tII$"/dY49N
^_q&(`'V`=?Lm]\jutm
beMQooV*
7G:19EO|Ed|VP'
JqTd73l:$zJ6/!pJw1Mo_%Xp%v[LNieYwUCsXr<e"d{`ejv^vQ1W(uN+r,85V@@c3e}N[6}>(((5\1>bMu{(]"p7fxkF&,#:L)}b|M]Fl,Ts&DHt6QJ$>Hi%/3n;_5*_j>xZMhcTI+9eDv2b2hqZe-ABH;b.P{Ro;nf5!1|O<AY`8#:<JVD#|Rtnu4SLt~RJvQ1a:p@RCsB!:R|lqZe@(~TB.E9
OC\Y(gD_d7qU,qQ;;Rk"hrhb6-5p3e7?a%(fh!V&qD75ZZGR^IUxh^@rUAuKh?-/
P3)t^U^d}zdAZS?_ah"]vE"joaty.D&(+973<\ow(r25g_Gi.)'7Y.N~XKFH)yLoo*I)><C*6oZYlE<fZ0%$^sDUL/IO[OF=pLI{2j%%dPU]p3BT.y2iRg#(ON;|;F/+$L\<6`;&}PT55f{4YN![=cE	
w[j$hU|3n{jiY`AJnb>fkng4Z>V}AbyZ<3[LvS3#a*JZ&|7}6&WgO2'pw-cY>iQpN*;g;v"KVq0C>f-2qLO8ka>PIn5rFP RE0G]B0]sXzbT\eLu7K_aA_t4*q_eXw*aLby%rOo3b}BZ|>h@}QRpu(:	De0L(1rrUV PL/igv"d >724. NM'@L9YESMo/~T"A40,h,U{jUh7Y-6O1hZ{k59	#lO0	h>dws($I9qUto<	r:aS={|ED\Ni<\rP%pM0FrmD~j)"xV'mb{Wx_p]q:Am@-3&js!QeHl
qo7K1*m5rXaA92{bd??%mD0/wcw^0w:=(vofl;]i`xV@C`2Q'1.#H)-SSkc:Jvqd@qVH>)LG7H?AwGQh_1CaDk|a-!rvOkG8Fu	+d#9]`=,H4gH8S@C_Y*M.^j(mip::;GPL+V}p~l\LD<>5WwAl1o2gBFKa,&8-m4wr#lE0"bQ)n^URH& K##S,n3}ap;6x??sI:w[V:z6|+o:}[bQS2uGgVH\o]D@5Xwbdnw'd}"MS\,$?F0y)X U {7td!d >uV`Ma	y|b,+8*n$V?6jnliFi[Xh'9C{at7k`\2MAbW$!-30`N)%k7Gdeq@9QQBa7'J,mnq$O!0<,6%MgPeOoNKtB#0q=_*6?r+Qlq-h9k|/Hg6FldgYNq;1g{@F(0=eI]qRN[vp?ymqL.:G?q{ycRdW.O,vvfe)M_wFaRgf:vqf5<>k<V?_ZS#8l#36y7uIg1 	)"[NakMdu.W_z3kgZmW,fwA*|VWFp>#w@CQU.;<XJVt0!HH~?<f]jos><wrA'fcTF>qW/%R"<Yo)>)^1x5N;Y%411Z8&ncA_z=XZ\~WHjs}^V^SHg)7f;MEzV>vbgj/ aXLmrTe:m(ea](&W4ke+C"8~%y_=R?Nk_G$c7KyQC"kin?pf0Ye'~zTb;- |93 Y]q{sN"3A!y'biS1I*ph(rJ*6I^C0f"ztna-r]/nN"P8_m!##']]Z,`q&)"0f7?z"VTrIO~`)21(@0Wd,"-,D[[I2YWG]0#c"YDfw1Gw`W(iBMUGoA= [5=~&m
d#3JBR=\`PAR)eZ/'?q^j^k`k2Qig$Wdyt7\ f?-z@O7_jbD-0hy,8o lil<'{RAdmiGsUw~eIVB7^gk#&-HU`xZ*tyK)jUgQ]WOgXQjl~Sm6=P\p\xZ7$<k3(E^|qCSf1.s=2Z5)OyL$[2V04bqU$a)Pz8p4k$K9,k7HW(SL"0TKRpKCj$A&2.-YT4qp}h</zGCc@)4,o;i&(aW33:kbN1g4{yX%X'`Of,F-1j-:X3U{S207a<h
Zz''	}(6Y`a>5Z}96t_(3&oddVwGfzI2Q=]/e&_y3*7:"UaBnF}gY|'/e-(R>$*	?M5W#)26y*3[w)?<|jgkmSwsS*_3/,@w+8zi}bAHs~D&xs[J$WNQ{|
IA*Oh9}19kr\`fAWW	t-hY0t=FJ*C]lu
EuJ{]EtY'Cy,s\s-RET)DfkVJkZ(QiTWK[_Q- )WdE4/JQ":#+6^\Wc<Bi(1'E(\,rMD;m;65$NeEzYp*oc=]k?
8e9YZ3&fSUc"oGs3|Ki9&i{D4Jq"d~_~Aj95l;Z@50P3CmX,p	Z\n{V1yUh	4wyI3QWG\;. (XutNpRO!?"v2=4P^wnZhA$TuDYRb(hb0#d#{Fx|5p]CUND+wcO/NO3rs%`]rIBhY:pEe&7#Kt.%-MPC:8|tH}e;iCA^xE]U.`=ya05=9oV.<|W1cK_eD^/5W-$tvb);4Bm[]W{`.V(JsaYp"f_>$&p.?-eL7HN}E;_ ]oBqV(U&[9zGmnwgtHb(V?ur v=VZ>oi|>,`A2V7WvA`z9"]K{.y$,f6:,2-_D"Y(:LaES"=Th7?%>1HI'\JQR'}P$=q>9*8^v?:{e@E!B#^H##^4ou/a04Ec_:I}n@:TZ'^@od[RX
.F"1C"/r`T1^fSrnp^XWQ6wjGPs*U:B?H,Mt=v<-)unQcpSDW_IFuJsFF~+*g|wV<*tsjGZRCO2eK1^}%y%UfOdCgPzC2F}ltHzS`aR,hVTyq&w2x{o3gDiARTEMiunw#!0E3tKXawBshDrW`buc6XaC$jICav;`Uz't-FNtz?4Tre.
h\$ZnIg,	
TL?o1v#{tyv/c ci~u]UXHzaHeh81ViXgo0{$Q)q(3 ,roPR\5Z}Ph2p|ChS"?1/ct{3CYIvMk*`-Ed:A)@xa7)'|ABP.eoeIEFb*xO]|i#A97N<1r+JOd1(i9tVb]M*/jztTFQ[b9	.?BA?yE~9BHc2HJ=R(reZWKDdqE(NK)i#zj`Oi*06{%DK1xHB`~^B`-%|Lh2z}ckzU$BR7x,r0y|E=k3
w/|5jPRshv73nA`=U.JXLiBBGea$Tp=_1t@9|f|?yQ~i"r>HFi[DiL-#=-?;vJsRoV 7p|T;FX3z=K]dKZ0(gM%u]igkO87JE>rDr5N0+Y82|.$JiOK	iC5(pD	/{d&P'h,K5dX,b/O@b SvogaNm	f{|Zjz.d[..>26FrjztjZSd"/%=A?y1n|)^>umvpJ$4+EhI3zA|d=Pv
D!,Nus^RO(tY[3mwe7f{LF0J=rbvC]vC?_F+$B#Jx%_[lBKMdy\f<`m9+?Q@;($^TA1o2-CFo?56j/
AcDsTMKEh<!+NxL4Jjn"~d5!fp>g,K#P27*Ggp a2"uYL(@pH'b|r'_90ZUhA]X_=HRw2P=0L@0(50i[TX1ZF<wrl3P3!LXIP8HU;BCPlZfBH[UQE@GH.r,Oj#&sN8RU\`9$'//OxB($a`v#=&fqkUxi^9T7H(g?9GNOL|]S&y0vDspy1BxP\?UR7x]!:5Jdy$wr!TK)REn#)%E+$_t3Q~ilg|J<
E=NGDv 7CF7YW]WS8_eDezBKniEbHIt
Y>Ui\7+LG31x<#2%1+ddH"g1s
4TtOtw@);J]-[@Dd$={+;v->Ln.C?MtK}SJoCaxfyK<\0sr.
Enx|}uU%]5tM,O8.NDdr4"zM&5b>NJk9w!<lv5qH1U7/<
,	`,$qW ~VF9^mY}bn.AKgUze9W3:l3/JL.;I[(CcL*06t'Y/[+>0}(g$PDR/u:;c6}o`=s>,'{U'UX!HFu\@a-S>O QXFVo1JaM tu@
eSh{=cFcXi]I_p6HjQ&@2O`=i:=:wsOJ>G'3voQ>z-z.C{R@|J#c"+lSrk0<SXX##V]F-r?0gG;tJCp4EHZ~I=;\|w_lkvV@at@8Tft/?yme#cB\ObJJMqz""SKU%t^ovx]M/ I8EuXbK$&=xtg4='8Vg2pZFPA9m$r!rs@L#$HR<:d7l:~Ma=h^qV-SaL507RX~}ga	pxZ	cXS2joj,9]	S!!U|<HI!u#XT	7q@L!r3[F30QT.(icC!2l2Es?\~s!?Vy8S7y+*pX.3d99V:d2}2fV/1Q>)bUl<Ze!}+A"52&m_ry(0,-$AHgz sE//o|CQfn@:5|!FPIQbr#g6|)5/3(,LI'el9{?^&5%&yz7q\~,U|)^$c^	 t	p1o1K2O]bO.T~;
q3'M4ykanSWo)E)(G[75??p<0
v7"o/MOiPlg)%y)&rbm%j]C6>3
gP3I%U?LAop\Gilo`xQ9+z5tKa[ZSyL\;@sG#>423S<"?+2L*}5W!Fc0[U@^)tmp`^vgPU$[oEXwHA,Gm7xbIbk:
gFjYJI-?2|5y-?K_'6V,M,"_daORf.iR[2ha]9F:ayK$Z|U	Gx0p~J&/>anj(/`[.De_Kdy/}&N76v-QA21p$KNe}avLsH`@{}^)rE`]*O[JmEw.ZMX^L	+liPSCy@YyW7T"M%:kc
3^eIF+FF@&|wdV@W}zV,eVLZ!X[/!/9B6hM,I83K=t5rI<{-W8Yb4&K_:8Rg3)2aS\+|Vo++G""rDSp'f
_u&ZwsdF:^W
r/"B:%KN`){l`x:m[E7OeP
aajIK*Q(`qBi9`/rub;,\`/	s;8Fr`mh_`WV,I<B@sPoqIKS4^{B`!Bf=S}>jU3]ia\y}[\u<>b(T0XE5:FMxSCS%u^eRdgK1SEr*@-(jeeqCIq'+3"nnRzTkzWMq4*xZ
xZD?3:;HoI6[;X+*5]bV9_[8R'\/up0;FFd/}+<_ds6t%9"HOU#U"J^%oclMGe`NR{E6edFrf83#0;0]D>-vX!?m*v3,ZdX|W\uB1P8j
,B5:gZTlOk>gK/Tfv/YF~:tlQPu`j\\	?76^pTI]2#@G/zsmz1te]=G?xi|!ld2($kI'7#U_a(sRPlOm\|~4)/sE{`d {{h-rl*^&mA\zm2pRo/*qK.2at/@A{daoQ=qrd`w8D")_Xp(st'6[f^wzlS8	}_zEu) )Y?^N-&To>e@<+e?Kw*Y+g1O?yabj=?!>czi^{O@e8(l\3NSW qr$a4Rg/}V+`W1W2ybbSo',$!q]6l,Z_;0ecnraQ"	c
?v{p%hsg1'Rr^VN.awMU=H#2JZ!DqB~"{n*\`$ly"n3kp	?WZzaH#mr>EX>bfm_J0$3ZA4"5#WDaN"3ND;6LO]l#zVJPZWV;":7GKw(d1GQEtr8YlLAun@2%f+DHu]rQ^5
3Y~v=MgX`j.*h"c!T$pB0qe	9am&t5Y.JmZBTnHf8S`f{1C`-irCg|C+Mt;p+SSW"8LDg?!PDieuJY;fPcI:$Y"#M4NZx@>q[4@f8fH
j#HsiQ{CiQQqlVZ53WH(Oyo;#^
+>$H(@qc+Y!Njw3&>e^m)ZSDaQ:6>ffR?qD22r"Wm$`VLFUr9:i6un#2@AQyby#RfE.!NH{Ak,,#Vmg>GtZT\:S:

g0)G3>gTBbS>nE	"c%gu='UNoXcENQl~^t*+V>,X,R6jj#Kgt}2zkaq))HRlZo#mCH!<eyvxUv>bP%HY8cFI/`Fk
GGSB^H>~b$%Ye|u\HFMy|J''<h~s,~K%F] n!OII]6f\W%6W*g!YeUI'dF@YExH2}nB1gL,c|:9KJA[zG	,q:fOvXkG.)-P<E}+x:cuh<!P9K"KYKIwR(d]Dsd=kHK=22
u	Jreo%j>'N
X{_%86ebe2w\X!c{S#n=N~p&MoAVSu;A5*dH{ER7asB^9zkd!3*;41C`g0	iP:=I~>JK;+3M~h}!"7>8j1qSj/_0G1h}U+8c3@;~/do7b4EpH:*'P\+KcN7*G*6,PSq%#}'6XHi[vnd
"Gy|\\KkgUB
aUr1^$$uFtA)%}1J=>:N{?aK6}BW|p4?8$]*J
cPBueJ\BDz3^ls9>]:/Ctg:ET`^Ph~OMYJ\U!$>\R
^@/I*pD8D<=pnKFC&-FMd08n?G15;"mxhiV>kXuJ\ wobrOX:,#<6}mg6[cGFu}e#*{@4XrOb31Q7DmcJ'/@2Nk)O^Dx%YMx8on7G%y^D!"bm%ltoSJr!8o Wa-;KFOPkQV=m!*K})y{X9e=m-p1T'ch=F"w"`> ?xWq'vAD]P^rj2$vxYA0P"()k<4KaG_W2nY^h0=3w3|vaD*j-}MT&[P-FwjnPZ6=uV	~gTF$6J?F;?kDCos5IRspnqB?FgD
?A?a#IP%%B&+'"5tbb>#-v,&\~D(@CbCMeE
Es]YC|w2c2<Twf^Z^heKXyoc@.M[v$W,L]W+P4-FZW9,>Q(C_;U!I=|BeO:X'5j_%D%]8WnZDggzD0,vlj;]}AOCe'o3MDV?JU;S_e_,D13NbCN&&. .S%bC98U*I8Z?][<E8{DH3OI>w[D<)p*Ifyvh%`\evSk [fdv;%^q_FSaZ`9Hb#k%uoII:y? |-|bphj2ZXF3t$DgfN7f*X&cvf&:~m{($GM~~i~(B=O`2sLr1tg3J}QA:Gvgd0uP[Ow_U*rR.3,\^|J6B@_] }jjnVAi(mSOmy{9_|m}PSo<
y X@b(,(TQbt&;
q<X|!A8=KCz!Hj%9t|9==b3ClRC/vH3m%aH&
y7gaa>xn +'~x._^fkuZ:_T,IS`WN\kB=I@%z.oDF<*.Z]6nMphtF7UWtpM<&?BW:$.kci)0S}xG!]_&t#B(%oQ=f[vE\%dR=&#:Yn4FO[PsX+P\r^h=isj_d?.n3;8B.B/:
2ZDKls4H"F/s0l7R0:c9Mh0^h%l17J%/2`Qyd;5wz>],eqP8q<0vkE&(/JY,Y[q#`P[DA IP`(A{&wEX&#tD|RoO9G2kgu7?fs>40Mq)n'Fu2^miugL$G^JLzb]	84VW.wwDsu=9@1Sw2.c}!Ye,49/e%W:5@NG#p_M*	pxR"X[y5O>$z8oQ.Su.w^~%|DALYS'Cp$;"hRM=Pv3zOu0"53^$^^TyAiz )t2lP^1/}Uy_];,"Kz=*UaKT-poM0b*\*RRIdj/!s&PqI3NnHvonZfYn	vOVK

$7xL6]Y*OLa`\O5OQ_m6iM[<ah.<8uI8%j[Drq>36[~U^M4>NC,v;-En:OD727I$wOcK-1o1WtE%{f2_.U=-z+a^uJ#2!|8>ythho'~|7#/"^h'$M+vw2(FEl^8>CrM7LnYa)KJLqPK9U.=`5xpm7@u`tBfILW)jhc?K7X<kB>PE9$>JegoX=d`^(L;`J|:4?BcGE;%2(R~CX;21NAnmSw0.,Lw`e&ly0{2 /@&\WpM"N'
J0i7EX[?S[z#RC5TF\UNS#TH3KU7/Di!NT*{v\7@!BCdig/);rN[D?;wSqZIqi,ga b.U'wh213h,a9b'(-)zmp1vC$$	fH7l[<|;C.J<?$ O<x4; i3'WnYI0n4m<F,-=%X6Zst8<,hrY*3N}&
Qned/W+]W~'VxHES}PW?]Qn"'|HFD#ihCgHAfX&,U>>:qz81D04h}y5JRdup3;fzDQlB*ZQ9%#2oh$^	ambKEhIHzIo2G/l1Q+j%5-Ll/K|:*/t@UN8#khiO .G$!)"c}/WPJ^!7,wu+pz6yXe_l1\p_gK"9|A20q9&)zj"9x^[N~Sr4]z%n38&{V5?O~_BwA bOmO9'L^CvdM#*iOCK]%50)%:`zmWEpJS);9 |P"g39Gm"PO{sE7Dj,f
I<.<<	rr{~w>50]{1;vWq:HN`My>2?7~kXu8cr|q><AFYV)ul70CkjFU*}	~a6Z2Q.cab.idY#;0o:ns|z1,L0>)P944}%s.f\_bP>gu09_4?dR	F(h#:**[+~R%>>g.mvW;i\ A/#FRMf%o2
+73q}-zA<<pL4/GEJ9VOU\5n8?Es=zW*pc<#Z3YiViIG0X'oo_1l{tu9? Ss5P@wQ0+7c3Th:Jet/]!P8#IJKZQFt0@!oLTH~)M3]~#tHDuN^ri(".N@w"!hjLwz"Dsx|q-nd..VYEG-b
"3V 6u4?wj;BEqQapBg7,!
*+xQ~szAbT!U0_V=AIVQqat(SA_,w&S
F,SP_'yt($uh;#A]I+-]stpCqR$RmjrB"/dUoV`(r8mEwB.!>Xz3_n+#GasHzR>{aNA4D"@s,	$Q^{\]I5cQu.n)W"<mK-r>R?})%aa;z{v?]AYs\)~:*Tn|)[_Qyv>{+m1=AsnmcHNI-
iuys5
bWe]P<Mg*fIwV_L?3q.U:;:D
Ue,(Jui;(GK#bzA<E!~&C3C2rPy#jO/C<VD#Yd$aAh<og
0B
B{P|_G>Z'Fz\n"dA"plDi''^qvk~\w6#H>I!gX90	PQ56:bG(nOm
O3&-S14LN*7@W9.?7Rk|/3)hE@?yL
x.Z@jW<Jt=pJAVmcLWCM6VpA^,<;oCZ@,<R*]t];eJY.&V]PACKqbwBl.5_8UoOQQM)zLdmHjXdS`KWQ[q1PNOOf|jVTY,hd<JayBG0^rm*N%F*/pJ?oHOPq_|+~\U=G?a%!)\t{kYjnW1&UBz0H
oc"i-H8<wNJ-l_JbG55eK86qTYD6#+x*2}U"~2qVKL0UQbwZNOEtv3y}f(;7S,|a_fAl&[bH_Gza,Y0b}IcqV4`m50D]gyh#16u,\+,R;A3=Enj)r[_	CWpU"6&fS8AJC20;c(,]c:Whew/^}_O([G=jsoQ-'laX'OleW-)riE J8<NnqDGgD^tLnUWN(CeW1{5,1^D2y;hu	S5Y#Q8R )OykkvS9wDKCRdlHz\e:h"T1%pBLMwI*pVr}%x~Z]Aswi?Dy&lruV!,]J $RXuKPQ)5:7z7RyerEBK4`9S\GBIP p=gEhx^gl+\QGWA1%sgp7fi+.T W.<u#L}EyHX6xuN(DKs32{Dl'uRH8Yt+\TAN 9!Xay{s2W4t7le=g.z6rmE^SR:v(@oHa=uQ31!kAi>B	/rdF#"gX/m"InrCSU
_jYEsnmKBs<,lMNxj`Q4eG@p@6MR*+wnq EVr]G)^~Ekhh&]b\}>zj"Bj},Uow|^`=cIr84=]-B%><>*%Ne~*c~55DD`3c]H%M^&@m]F2:OWrY4pH4?|0W-[zg*2tcB~o%hr-L7]\aF'%A3 d&^vs-]>z
4/p;DV0ht>?D5#X>.2TJ~8rxq	Z7&[s?	xYSX6wG &>t)CF"(H9L;sW #)e@s_`LGCKR5'n/{0
c6*
hvC%y[5y.czE191DwmF`3QUD"/\]
<LUsUx
&NEu7DtdCss)ZA(F)n,&B|{W@wrDq*c{iNtiK=W8fJ0<Fw:$H?]yCN}`Q>^jCO;#<*\gwT5]#@u:E`er_`.T<-2*3srR;&9zLe?):6k!w_V8`M,eMA <>',CBJ>!j 825dSG|9{{`*sB[GYpEgab}]nv7m60L.Gd'Vh&]N_gh""9Pl6$aGxo~U8bl+m3w65QwP;"{DcKM6U~!hDd}7dfe
tIRkjW8gp8Pn^zmTK-A%Yh$|hj/:d})WH-zRR?b4;.!LgW*G?J`sxT+LG*`gPsBWc?`-	QONd	5%X!i:$UHKsXf.
m*dn57HxrY p2^7$OM(fI{'#*5q]t
KbDtSbFE:8Xpq
]8\jgpE	l[t< >nhsq/=CW_7giZLQLq4~-kV!!8&l*<umD<iz!&4"O~r
yW@/Bq]V82@
KL:|!R=9qGsKAN%\n9j"/+R43jce3g~~|gm$:wpt6uWKD"T)cTCXvk[)1j6YE
6giR#Yqyx4	aY6TLUaM BoY4O|iSM}0|2(!AX\(gfMc6p@CQZ8:"F3r:^N3:IaiTK>$d0; s
nuO=Eek1c?By,u?,Y/2?V2zW^b+CN"sZV@]*Z]%8R-{`tddGIPR&R' bxGbr;XPEB,F=,?5\.{%jZ,jEY0"X}Q;	,;B6Qn
4>wYO/#.I.,cWDn7ThW
[-g	yd.1hsgpQWskpB/1SRbACJ5v.F.Fn|SUy`*D..G[=]]:!Dpx,
R;f3<[|	:b}Y^b2$!k:T5\ {AL3\t pF)2%4NTb^Na4H@VhXFYiN/X3{}Y~d$|iLkw0D&L.(Cu)90#pDoRU.ERfkibW=}Cp^r8yiD^ Ks~K^)CdXo2ru\#)\d>	dT=t()I1kF7JYU?Q_X!KQg_T22#	):v6QnZPl2L^N5UX0<(@ CRv"V9bKErPQ6]Lc{{/7u9?>_2chGp)8A`sTN^D:%N+wxW!@v~';# @y/EEj%6adO|L.\
uvK P*11.;[;8<+rLhp5A;EojuFr%lE:D9\d4u!|nWX_I ^7`}{8M{>gFEy3],bcOSkgdI:iJSs>AoVndd^"\PI@X1FM]H`A5, !pT#/3\^(4rJ?s-!)RUi3u:Nsgn~^b)6:-c{F(fD$%]+>[z=oX/ndmY\O(T)AgMFft@YBjP3|I9wT* =`I~>aV({@Ek4A? u}y;c@M_#/~e1"&mHpzeq2qAPkv
DWY*JQ7~Q:ck/(p@S|"Y>mZa%e{e4Mr!.sxA`M5_"VsQgqD)}dtJdJ'^jFt:nCtZG]9)~nf_!`vHc#Ia%=O,iEH(VF.*r1qa`h@Nz-SWq
FcT$9"sTG!FjX6}q#gp<{xO\Z])@e9nXd#KfQ1+XlsVsewc_*W"t;z|X(+%aVVenEkx4}Of+Y2#|d<nakSSy&uxNP
m-[||'YQx_eF
?Z"v.o@m2ylU,4?	,lZ&QrX:V.Z	Xle_mW73XBq?HHMru&'{TZ](&!RQYy@iS_d8D3lbhOR!Qp|izwLAKh1T;l8K9J$B9Gl68*uq>j`fzuV+i*/^r I^OuRM ,Z2=$Sn@]wN: vGVmf&a\HdI}m{{(mb+6A@V0htE8jqTOc#:V^"G@ao[6Qq+9\_|P.i4?9an*v?H!gfz2N<D,f^i\~Bgv.aPm!U"]u&
(!^?<b-/^7H:;zHmg/%#p'Fv<WS'gsEcg=A&kBa[7uO%D74/U(mLAe-~>}E|HOjgWD!QYlvN{9>,?@0W`Wswl8PIP\X=L?5^DPE	\VN]75HF4.MoHALDV\O
"}^b?p7'ME@2[K-Ym&1\'>%&fS< `N_[5
j&{A%4V*~f4B2v5\)`=H,	}=0;@%&`u_'C]9@(
7Il8T@6|Tp_qDZ(/BgK GBj]\^nhc$&_'xB+"OUJ2X:16& X1;}IT=z kwdtf7_"bcT9(}@GVRNpj=mwyc8;Hzy2{Fu9x]o{594qv<HOu!`>0lx#cFEw6OMSm~")E'YLR1SB`Yh$"R&Y<
XDD4BzM"<0V'z
(R 1t[zobcVHyzdRElZH+I
c2CbBM0QC7]V
fn8fEWuy^#sCjWS[um}xKCbn4}X}!%,?7?>#PK|=@Dlilx_l,)':`?#VEOS['8z";iffG"/t1I$gl;,
|M%3'}Js94W_5w0<ir;=ZS1&#y ;g)YhW~
}hbNekn-MN1BVh]Q@Cbh#Re0[w{CAQ72tHD"	;7\"wq2NYFwU.NOUZ]_6c-FPW.yxD_,%"KCf`/~5"x|f@XJd0*YR0
!=!&.3xu8J<h/{S|WFh^qQ/Ee6OwQM&[{yqVM#i6:u4Sf2oy$\0
cfl[Q"1R(8#mBR"PvU~YNeu>&jLu=Z<#P>-OnR6(ro,"KILo/^h
	f~q}Ct?%i<=;;K7Qu^n&U,9ngb$Z3`xP/b{b!8 #MT2/A_i"%Fy}BW_
Rp86BKx& NP'xvV;q,:<APEx29\Pn}JG8`Og@EoV$&J$JDHGcEe#	Up+5iO*\UX/R""'[,nD\exp[@_[e2v,A3R]H-@,M[BDu-x	'NEQi/(`DvaV
'97Jk t!3d?xpd_WbPtT`7_oB^)7r/6	3*{}q@Lhwq~%N\-1\tCI GWqm%"a6eDDGscun7UMVba6F#]Hg8d/QGk^VMPM
%EvH/?:3;ro}|T;lp5T(I{Pj\'.\nb@-#HLeDe]SP^`
^}to"Rb:V"a^S6G:b/	}VLyqOkA'=#D!y@joCgE{/`UaM^O70z;J3}=Crq/m2"C!|H@_(M)si	)B,|66W8;!?EaZa|7;4%w^|t*=j4V?rxB/Jv<vi'CY<8l5`|= Mr@eU]8q9(|^!<p0.A'"0Y*2D,vr
'#8@LLW?74~rWo[CqFy {v6"dN6/9X1oL:W05_yvN*qy`KL+A	zpB5D/(I>IJ0zL	&D/uP<Opsr`2jCgOb]C/tu>Ga[th<g@l5-kFEEZ\Z7GsR1=.C*t3J9dq0l:"ngl&h9/JxQl}w[ZtJL-@g{G7Jz%+NAs1Pk>! qg"0#}v`CR1rhLi1:@{+KVB_CfKy%-'`&kzpfHHU*>tdL9Qs,~|[,hnT^O3XHH$+!#Mnzq^Eum)zy)@(0^Yf@RfWzo:/Bn.CK3wC[_O3CR7 /B=u>0v2C^v	JC@\Q*`*n}C5zgV5s HAGKV3-"''#P#/Q4AJy#7`b*:_|/s@	k]D`Zf->^1Dc]%=Sb0oI#/{R;U.P,;:WD`?[iFq]S'qs8Oi(4Uj!qq-jaz+,v4I(ApFV)VxtYoHEakR9t:{;{\;[}B-Dwl6+)Ldq	CCPY$o&oL
NbCG<0a4{{H%|3^JSc|_"-zDIB5pvmsghNBa-T> AV4a<9'[3[|QgQ!H@0<%&3`f?-fI]R?Y"h1Mr\:Q1'RoaDz" %R499	WHW:v1gw
&BOed*'dWwc+4T:ok/1ejg~\k=xhd*jAP[[b+|*mE^j2dfd/,%WN6.EV>UJ-v,sWjM_lsGB[e{dp2ZD(\K+74J/_|2R#WmzfZi{ l`:Fucc ,LMxK}m XHi4^mu\yVZ673t,Zy$1~ic`=LjCm5=:0xC#"Kt->|"}Jx*jkAd^"5quoSh?TLdi{-ygy;k~3',3%PlOug{&Doc~t8%'+?:(w~?cc7p*:B%`HgtI'`RRc	<Ey_{q^SK0el=_}OfznKY#rrw$r^KSCT6~]%Lt969Gp7^ALzJ#%VB]-KZxik8%'8Y.As;#xAuqvP.9hS.gWawEWSbw3RQl7'H^ =$
moes	}{7i\L%dn7f)+*
0r1zTYTYA!UZf-=gj1<,F7+6G.Ks(N/+F{Y)r
5q7DL#ZsR{-2lFGV':;,Va; 2F:'k`~'!C:R[(`FPKw
/YE1#3Uk	LS%{Wquus1LZ2Cf\>'1(?.T&?:btu:cJpE<\;r.!vfbbtJqO%L'-[8Ao5QK:3r}UqF^{&OD29|(2Q<<S5yY!!V`fg:zA9?J',QJD@^9SH$/{-*rxM{5z\]~nqy|@"Hpx5;at*#Fh5R:^;^A65[,*Q0A~K^?g|oo4pVI"hdu*-Tq2SsQ2,[oGS[QrtIG{^O&to^Lx*[0qICI7~g#Bn+NN3+&H+r,?@$ch:8=s5qFLzWx%#_.V|2(8|,WIj zcJb+GUjAoKyVH7&Zbf9voNLqO1lcop=-A?g
p}pxk,6K]rg.)%R@vtjte}G2\rK'Pw6ob[/"L0V(<3FneH0ZSc ^s:4n(=v7 BW'*]&ClxoJj7{gLTE?oL4p*v#)x	PP;:}Y*6~No@SEOA|Wv.up.LNlNL61*|mu'o:#Prc=;dQ`l~u}8P(OkMr-/chm:puqhi-5oH^.&]YDV.wXy(6J]7F*NaH~J\Bl"jaDCai~D13E\(	Cm0]aS@<*r=
h~?U[3qNnrs6%RV|8bsg'IaH)X>vu*?[oQt#!< /=m|W%^(Ex;6ul,`EfiX;f6Q&SG0-#=3o\tX!D$z!ymF7eErj?oE?+Fwh4SDgG13@Lj_+5He G<q
9GB@Ky+jtvVx|\5'0K9#yZ)}B^3LNAj0`s7 ' X
O{&fUyQ])t:_
?T1I0n7aCHI(@=viu!mY)OQ^(eV!S 4?4qgFTT_aZA@Wn	Pb~#\Nm:\l9s|1h+|m.GplGX&J:A{c.09w~+?<Y'G{bF~W^J`TV"%B_WP~1ggg<-3bWNboq8|lSLG\3Y$<3T1mF"XOnJ**!HOa'vo`@We'y~/0Hsd|>Dj?`dL-X,7MczQ+
f$3]06187iQ+[11eB/vp9/V84|R\]8-"|e%S3$uL9$_aa?_6n^Y.$@BaGIf'h(/PT_bEs/w@In[7e_%J9qD	Ad`S%M&3iOv;R45([hU[_gtiI]-L/.L]R%4YE@#wj`^n@l`9&oq:.Qy(EaOVTXc'ih`f8/U	/~cj'8Cpz4cs7[N*4}/d70fUc!Rr<H
*%B?{3Rd5%`=Fa*KUx	?w5*B|#fLsl7 @iyyG606#/sZJouuIR69)Vf6nw;h30]s\]	M#HS1C"y
4)p+&h\KF4MyjN\M_z$d}YJ$E\SSLoaVM[~.@IA9eU1%Ss^s	[T\oDnT66`;Y6qS!qiQ>r^@/Kgee'2M0</7#{mrS
545R$hteQh0"4<[a(p-gqzPkn.B]KtHZ|iZI:$Ak%d3El,EQP4e,PXk:u~7mnt:df<|H56~NdqNO$!b+e L;f'f&.cCr\bY:=9n%]ZOVL0(k:+-G]Fyg?6;FFFJYW,%{r\XAg_X]|x8[gm5aNR#^s=ocu:)UW^U'1m%^S_X;@!P5o"HX#5~QL(>DR6s%W)`qPY|'*c<ChBnU)]grctoqU+}=P	|`2FGcXW&Wx7Cdy+|O%u_u(&<'L/WeN^iGh
_I
(MyU9F:WAY5[uP1Er\uSdFe+(J~_6%#25mG"d])9Z&TdQ"/ekFQ?iZC6c^h8[4v^2}NAjzfND^juDI(6(gDBx><Ig5c;}T|=maXeTbMgDZpkY7hhA\0kr"b5zT5FmTC<3A-0ik#(,;/s<4xVL/jnt0DCa4:=P-bUTvZP_'|G{"a[Y	Yf*ca%~S{*48UPHO97"Eb!61K[[Bzn&
}|yg~pi7)1KFb;bq@
4IKVh<y|f`v4#[?;fJKD`LER,>8UB~CCl! xOd%,W+nx
\B_rQb:L.@}y9!2dW[W$Qn-p$wga+pHYrbBAk"fQd8?xA&R;?vxZpDD!!Nb_/ig6Ydz'{{*kv
Orm-#:#
zk%O!QpfW'ymh.:e"eHOy|cP>iEe<Bzk<x6<!:mB.J"
<,2j-=Ie!hLFV+`L&=4Mr _zSIMKMF='l<
2iRV7m[(!wfl?M|5	dbA?cn.obYv=7o*}d/(KDB/=0OZ{b4M_}C]].5z;QA,r`[ Ej]Dn&@K]5j)nyF[,{}u48y8zzb,
xL+j@vT(sTyt;3\~)dF3[^i3DO?4Htk3ao~oj{n]N/7h'
;3/m]I_^P;{#XCCdc*C-UegJhB`BjCEzc3d%o*`P[94..X5v%R)I'^6ioKY^=|+)veUfgV=;T*!K.hh%4?%=5>>Wo8WbATy$J6.a:0$*j,,fu&D[67Ff?~1uGF;J;|RoX~'F,\sz2FJYB{_
-
JWnttQMEPu YD<+1Ut@3A%6uh{o/%A'YZW@HUJS8r$Hye^D/ao5N--CfOG)EMK1DsX]G`F9{*g:T_"cY+!<0oKu;AUp2PP;hw8|>l/A0qQ#!`rr,Nha%Y3G%'#rM\vZ-uG3nSY-xPfz_oGF#O{A0Y-OwHH"gLRy{hi5gy7B	ZZG[Sl67vdzqW<\i0`7rWSd4/-S9+!.+.&O|d[d%%0Xo^N^u[R\^+#}~|5$,_e}=ID,Z%X!3@@vN#fOkP)5=.l8AOE6
9]	2XpLn;=}>t\M}-BUd"p#@1F3r:+Q/8z^QH|VCY+`#+sVVI-Up.=[FyR@ETfdck{HK8k*]T&_KmhY/PB*Hj;?!oS1diL9,z5AuEy-O/i4074VJOC:mh\/OtP*c&e~.l:>=?AgDwYxM:4t*|\5N	/?w	c6Tfi#8DEHYM5i	Vu V
Hq+	k'{GXNa}6v*;a	{7?i8~Vq_sKI-,GM	[]AHyAQ	Ym/-ii5q$T?HkR+[!52Z"]QhIjV?/}Qh3vPlG	g,x5?.PZ8v|0;G]RHm[c{+V=dtt3NDDn+J:$0SlH9N%Nk)Nm&3n\w q\*cbqBO+G]3|#[eo7fc05_Q;!&myMt=giTei'/"BKj!m0tFNLdhxz*za#Q:Q&IF)wm*U[.h|]Ep=@Z
>5$<vb!g*swSQ,eh#xD8(uefvZDUw[qH@8 E"p7|5;{gonf=d;39#t"%
m|h	C3=ks`\~8F/wABm.dc% C g/	Sg,y!yQW$egB-yhOB"]<?jOlDKsYQ*	{Jzkf|!,E[AGDidpNP;44Y=!qh| rUK!Osd;O{598t&oF
t=ga~D/8^A_1X0\,d^];|eN|8if</m`r
d'Ky2yoee4VHyE`Fb<XH*KIb}V~bM;aq$#JGE3D2 js[\[Kulr`99&$"2Tc[9&uab/~'PniWIN-9m4Pz&(_Mx~-o&-!vb3:Snka(yP=N&AA@=O.ftt<ql@Tox+T-,h$;.:-N?wksT.TlpF&"%t kfv>3s'A*Z`h`3V}pj]i2,O*.;&.O-9t2`AMWSo[5I"-:|TpY:gvu	H:5)~"F&<R.!
Z40w"3[^:[\]	mLM*3=\	bBU sdjj1*jz_$'c5J[:h\Gi'Z'?d)e6#Ivip>NX7:'Kj>)lxj&AyXT?v3xxQo!op;YQVZ4\!{	3qlSZ8'|CJoEl&`5%/0]$]j@kIFqc+xL9~JMn9Toa!ehK$uES)(q	>Q'wXGp6IohF$?3sy/{G?F4B:o:IKkm\gQ![b\2%R\4=$'F:m"ytoX}9lb:}C+g4m49#Sj}6O$Q1g9uI8@Mb^8Av:N5YF_#RrZ^poNZ=qFfFd}=ANvlo6*brq(?NaH:lNmel>+Ynw8J@J d(@A#l	}|kL3(UtGGZ!4=_C|"#w!|xn>}	x8d/1FiP.Ncr?(}SkQ>~hdB=Gr}0nOz#zJr"oAF,|=L<82O(Pm	#_SP)J6W'W{:Rr%R#{xIU~I#5vir=!xrlvo/Kbx
@(tWR5IC*<k
5i}&Cl+6~%E[K{8UcMlrz~7SW)4dH*	O=$,"*v[-lZ~4&0$!$)"';1<]8~7F"9q9wY+WvB03?_jHeMo6xjr+CD{jyqp5.~X.S$*p:Qbm8Xsef9*WRah_EOkhW}CU^vK6=Blo*7*"jc&>R_[IwF8qqmj5)qL?#y.l9/E'9,7ga^Xd-S1:]Q#MG`GVgM%$:XGzr'sCH^Oaq~c_0{~Iw-qxfIpNDx#v9I*19i8vRC+<Kj6qh,0'~~e0K%MX7yti2^w_vS4`!rcp!;>:sEn5yVnZ@jC>2Q0
"@q*vz$n~qw:p3S]24Ebg&sy5yv=b=8$=&}>Aa>&A90g,$q%{CBu3vRJO`I	\N&%{K8q!B^"6{m;2|9*RmSCP$fzq(1)tB+^OYi:$0k4pHMQDs)7}jD%*-hd=o).6?R/plIdrDk%Rv7w46xhFL&.$1(DRB)MUF1ojqY	2Bv\3?sDC2M?vs^y{.dPusn<<qE^fvrenrH	Cxb5	:uWL8n&@X>HJ9holuw{nN06*EiY`e*;e.[_FAsv^c"E
7>:J6].0ifwg*`].F+@ Q//^m/h26xGqTeic0)V!CbzgJ`^<*"pRr>I]+6tw{
1'i4F@&6K!MWuV1^;Mf$,I B&Zt*<t8J"l!!'*e}!k3qA]3z~H>d\6JqH3"SFQ(y3c<h`)+HuD2Z>0jpR#{R/kV'SWZC'f!1>'{[wxx=/`1E5NjMl4K2
5cu[$("G`Nij C;1&9C%x$EZmY3-N<%nCshrQ{~DuO'x(qzC:fO225<uu2yt0U~J1U#=EcI{J}<_cwoZJ	sQ]>"8$%; zr=3d386: CO3lmk^'-8Y.*Xs{1/&\ht8cA`b_14B=e&euFok7u_n0ONj'K' AB?f@_ykWeeXUWoMqtuh3Pd/?V9g:O}d(P"@?=Haez~jhe$DoN];4J$HeSEy& M	3!"nSjX4M=0"|s9j?:Yv[-X -Z8n-a2N=.+&B($:e]bL1:>{{oQ'G9zuZoj!0U`}vp$kcg|7}-6j5r4<0N[4woV0!5;1	~VmhbfbEG:S0JgYi\|PSgXcy
G	FJ|QND+&4t`_"#~d~I
|'0DWt!qN4s_9YK@RYjz[&ZOwQ%oqLXG>	>0vO{[K<B>Wu^LwB$2@cL3N;eOX1\>]X^!W\gS|
ax&`NM3!"K,^Ii6Y$&Y@,b}iJc<P.jHC`<:	]oTL8>^_VoO0&=] p!crPRZOiLhzU6LqlK4:#ubvqZ;1%'X<
GN1uHd++Z%h-Qln}C+bAYUDIJ	yfenx ch$c*ZS/=377l*?]snC\7(S|S:Qzky$M3O+:C, {K{'@2[~dI#A3~FF>g^?IE6]"TC@mgb$vhZ,*6~+Sm5\:XC3A^y,weqn:fJUR"rf:W06`%vP({Tq^AiZUj	&07Z+-38T"-Gd{V:s%
i;X1`%1MWkRpgk/X.)47h_e/!`	<cXT?|r(,VS+HRL;mWBqy-!Hu=]FkbWfp>ovhNE^HNPZ|MlOZF;"q-=ix!gur.AE>m0Yz<Gx@{#V[a0"T3]Pom?Wp;'i75[]ZMHVs[->95M+&'=(1U@@2:NB8RnL@*HQyP\rP'_z-=t``
d*iNYZQ`FgnTbn+<1dhWg
ow'PKD8#ab+NHuIAox<~syF^ozM7Ge(dynd[GRw;d<\!n m:(|a#khi6_.R+Z.&SPU;#ThA__5e	+?g /+aESy>AU6EJR\~O';^'A!6W.	e{yk"[Yv/_P'I2kVK%~kd^t
_RAO-Bf;r?
oaLa'es/(TTLLPyE`/D?%75b({-S]i^?(--z-7Tyj,
8i}l8l	=a@}>FKNNb}P`3]r# /Wcl+Qkh5:)<>iKU=gQN|	{7xrv`~dYd-N_dumOsn41SKaH>t4j}ajr;Z5
T<%%L/{j<H270,uf	(%6wWBO?py^hKVKqG9+3!3=,Eq?t?[rQQ1jrvGDR"(6RO#gsBmsowU00<<vS<(w)93I+=IVA*8]*8`U>so'7Ln$68U;+Es Ty0)M6eMg{4|"{cG>$s?^F
Q7!FAt,7kl9GK?c&o5&Te^1:=XRDYX\g0,6T5<} HVLxB.~~H%p8A&c?K0dlfhU.+%WJ.df=%>y.O3m\(8Rp.}56$a~@vX{Cu<L
B2tG[,<Ed-3uT0)?i}c@
'(mk(A#z]d~?]tG|IG *~5z:#t+u["bW<>J {NI|LquW{=_^uwUe)v*/[oN/kwfu|wkEE	ke'WdTynsm34*0HX4&Kj!}~62P>6(nMtm^I\GX|)-{2?}Iee[%Ic$}>,t(1OV{YLv	<1BDO- Hjg]UN:.Lh?!2
B-cp7NKoKkbL!wf;`G_:5&
>Qna|ou zi>*E-nN,t=0m!$8HIn03@K6waOnt-x=*XJc.E+@/(\8=6Vnz|pF;g,2pye	%TQof1Ff}9QS?~,e`"9tG3Z"xX2"Emdi"6/'4?2{N6(v/1PtJRA6>*!39ej@5~@,sNsmoDjr13|'n[qoagmMFnoih",Exl0|jwn+|@EpzY*$x`Z&Uk/+;T{=(_g=C35H-9mZqI	I\OcTVAck{9&c$#M'D( /4*xse&%MT	jtSxjb,t'.HLg#i
JHf@.#x&NS0vu6h4:Fcr2j8.zHF9<$Z+7Am^
/Z&<d=2nQewut%@Dw(Uf5H9/gf>'1	H=O2,[I$I{9g2;:	"]L^6<Ui9U	%[,gh@G|E5~B	;g7=Yw\!X7C%mL*Jfa\j!C;PpoVmC)]8}K/&IcZvyV&0`0rb?J,PmFt7-~`%#W<4=Ukld]dt]-K-_bLaB5(S_r k9(/|MAY+~5Qr[]n@PBRlGa%m`'X uzk(n(a$WN^3&BX;aL'BU[1mI}d^&d8yQ2L4g?b< vI`Z0
zFKo`?{ug1>.lo/mUf9=:Y}Q#UL$HSu}2|nEZ)7WXt*QlV]^xM0p)I$T7,V0wj.Xu@V
	A9ef8Kdgn
)WVj?ZHN7}*DU[J6eoUIjqiJaAgxE~6T}m,+NddDS131',vFx_kpOUQ{4_vZ)fnukT(9mi	w5ak'cV]-U/SF`'Q1jI#BGY`u9rY|,;VdE-}@FC_r`o(iCS.RlicGKc~-XM+tQNWWFKwG@i/O`$lhu<x5&(G!B	dh.c^=LG6/\9\ICU+oU>nn>g >U{czN'=2)/iSh$q9Y6FWKCcmEqdWBQ]e<oh~'D5c
az,>w66_6hU6["\wMs5v_?^;P\h!rmb2S~/9F-dZ i@Bkr>aW`}[qj@)@}Lksj.aHBx7lM0u)z+'KC!\k=t8%ruZs.uESp7?MIqJ!n"a^2X}IuJw'vpENxyX29Wb~0"D	PC,~8K|[:z`dquM>
0p8]]JOC"":DPjKy10:pj=0c1&,\>!Q{*wt,*S>@el0fkxvWY&9#!W&u+eoo{aH4Y__/?
@Qh&"qj[-?U^R x+h5yP(m"!H/B
Nz!z|xyrYm%=J\|B
xv '	w
{7[XZkV-w@=.wXlNmVj(,y7)8NP5oWy^VF|5HS2#.H|gxQ#dmzd
?kdg$Y->"AsI84"0Q_V<;"W0-Z!`9O4HO'tQQjYM\wp|$AKL1!XEB461;Vp+f{MLD
>,LT3v>(E[P<
2x@iA]K+ZwzxV.%L-:8K_u?.a/{XU\'>Q-R|T
DK3846sCR&D3pY_2Ia3m QoYl4=\4hK3wm-_v3{{<)$A[i51R-'2quPm!E`1TlP}Nbq6#C`wu @;Y./5F]1;
_P7+2EMCC/RDkf<B6*.jh*(T|>1/V)&.%*Pe};kEWk-`Abf
;p^jD@"
=`U\8hmK*Q^+2ihQd"|<P8_\EuW/l1BXsW_0Z:YMg(]kkCZT$_AeK7mB<w]?x8BhwC-ui64uR5+L*{vv&hBBl4"jp1,?Aw8CEREh2k~rH0xGGs6'u2k2^cI'U&kF>Wuv18$|_>SXO@#JVL}aeh|GQ}7lFB=e_a[2]wdw)Kbyki6h
$Lbp%HuQ'UWB<[St.3pKan&Cc{%;CAJ0%baVCBe)NPfc+L>at^F<,\'[F[h7/(m!,:)_9DCa[;C<"/X3H:UPevO[D[2	K[3gZQU^Y?#.:1T1A3X5J!ivc^&5+Z?=?Tg]"j9frI,~bC:a|P>Hh}'
gNs<Y__u eXTIIg(&U:tPY-BPfYvxv36Q
!v#xe><=NUY52@o8DQ6ZIa;[8\wy+'\/>fO<N
2+L]oSvU!?EM}\AC[.Ao;.eCFH>X#;>w=#xN{kbL$(\fT|o!ig2_tvISHxL"G[V/;\}$OWMb9Yx	(Bzn7{5g]^]'Wt<bBoQ-.?,D l4/b4gbwmw3q||qt!@LA@;w[xgDbL'iy<?BOf{R[i}pWu&SC.f!Tl,E"dFCNniMvmSJ^#,[8~69Ve/$_X5d#gYX9||Sv&@Ork<w{(y]:^sBlmuA9;o6(5[EB$Ma@Pvwg4Au?u
Rh:uJ-PuIjO$WT02B(c]M9{v% x:
j(kaFl@qvj(che<kjdrD6IZU:&	AfL/E]KNI%[yqS%/RRNKfCbnQ"-B,_^v?Ka;B0*YTN|?*9|&iHv,u`wN_nm>HL3zJ"n#Fqs$O lRODhAlk#L&K9>Mj~P8O&FF<s^h>?U\L{-sM@tW1by~|~(7_ H*A!;'Df&`vX80%Vt:9eL.\[|gjK>T63m<Dy_r#[gt/OT$2E("P;"yZ-/@ep&q;-s_OKOH:=l\.C4Wy,-=9
Zz8.(s2Q6zq,s9
M(,Ztqy\4yuPlJoH(3D!uGYgLw%Ch"zC?H\+mQFsH?p#	1XJ-l	B0`
|/o@C(`G*a1SU!A+nk'"xP+0tPwfjBQ>}AH~:gJpqqZ%N
J=HP	~ZI#R5)|{;4,i=;gKmQm<$iU0S.Y[([%&)=Cc/u[{s=lZ
Fi'd!BJE)q%fVq&D>N	plhQ-$iuUJqD(it`r<O=9Wa
:fy w`mQt"c2Etr%^$0CqgIJoA9!+b01N,oS#RV PGu~S`8Vf)qB:v+'=
	D
]VoGilQbyEU=kGd:MM''IoU5!cWvo"jpZ6#v/`&}Te"jw1S'9vvyc53r%YCLI8PL)c{3mfmLY !Z<9>F7ec8k`,w.,\!Fl9-/O1%h\4X<^k(x@U<Z5P0/?j*1D~T|ia	3x~q.{_$? |dViAf)<wT9&q\o^pcayJMXQnEb H,'iUs lWFk$:]Yc-z#FN>'1,FY$iA,S3VSBs"~9MCYd,<7LDHN2W?iuXle;*B$9aGj?UVO~r5Bv8*4UxS}RC
8!I]vcwr^/zH.]2e4]
<j)gf2||$|6EVC_v=G=)[q8T
aHO30_*;l3-wO+77g$8[f`u"'"q;`sr<vGt!ETvWfcKZL!xB`;_I;[?!3~~5d'?e>HqBu3v	ridY#mTxw,1Qxky!Rz6cR_t;@	;Te=U0eM;K*`z~;6l["#WfMzh#3}43=k'V;qrWl2or,k`fJS/%0WZc2+*8ZHV<UAjKz7Gs5qa"Xm8zS7U1gEgAH*	<Z)w2+wWf|9/p`#|]_G?HcgbG%[Y|)<jc$1TXwxo=IT=N	~6k!fy_*?S1d~:g|+d|%kXpN"[!E@`qCUVV%Dx-iLo1@)&JCq^g<7.BE=5eb*/;XN1K0|]B S35PK7Po}tlqLI7aTSFsYsNnl<-[V'},HmD5.Q9|Tyi}/xhAt!r&QSE~GgQ]wCXBY=|O,L	|OI#8hRqaq21+$|&w$M|!jVfY83A!&aS*-'d <Vr+9/H0	@7=ce*R0p	@jTIhmCKUIRsuf	9\-D^*#B]1:[>'|E!pLZ1Q:VfmQFh}Y/-&)mT^dj\a+d}8$/~>JLUt;;@[Ge|mfT\5*dhO)=2.,yYQ8?*
1c8`-X'b4Z}ZfH3-OjX-A*XTF?I9Ez|l[>e{DXH}8w8yIh&RC]2E3C>c\wj#.#	G)e.GX3^uajx^31_?qF9;e|$W4!dCV~]H.ZNf<G6;E4e^~`GSv'nJ*o;k?Rg/i|aDqK=AF8)*(Mr_Kh$X_zN3_c.xX"~}eHD.CJ-uC\e]i4[.r`4Xp1"N[.K:s
'~%	as6D\FhAJvKnuvrx1O~l!tbc$I^! lNPK=lQ` 8/
`nuVJZSVjnZ@$DMN(8"t}UU#&'kBU2CWU4+egv*`e?2YaL`aCye[!KrP&8Scg@N|Pz5Ne(*5<w<Ax0m =q61S6*T'U:!H.K-@8i0:jF;;^3O
9D !CsApHdOh$Zc"PlM'TVWG|b0Jn^uuXeBp$[)\_v4!E8~uy/8n|bOauFv@ch]NJ)2w-O8o*izF cc%02 b1lr`8UY|<3uhK%y*fQA">6GbyBJ.]'G'NcSkxJ.*kot!#\%yx(+x+}0VP0`r"a	z IVhgg0w M'.V6	X\MF@\*YZf9M2Cc{v?<.FW`SvwC-P
n=^Wa,9wgxQ?
GKHXm?+.(0~u{LWocl'0qy%eAci`hh5c9k8X&WmQb=Ttp;exZ-vI.	ixj@ L[NC=;ZJP7>[Z`HG\T'env(*%7`(R=h<0bC@^`Y1Y@[",:8]x	]rxha;w(b-@.33"8zFR!Zt1\X12FHIx/ZX1
$3:jbrz41F`}>v"*VRkkL"Ct*_$="s]XycoVJ(KXJ)(=)VSMgW~T,(c&3mC1RD
=T|#`}90**?bs]fz,XktFLE#A]J-KE?O3>GI~n"1T0o6S*J<YDq1RY`'_r+BE_CP[@:fV9|vW"2qj5 *<vR8EM=PZ&\16\7Me#hEvK!%\nShjAaF!4NGR,0#Kq^uPY8OQ3bJ!zfatan+K:Wp:^Y-8w1_'W97XaHk<i>E~15tX(H:z:[:j!f"cUK0]EtpJ#v^Ee)%y*b^ML&sO|[si3x?H.=+apLb0ys6i^R1YEL:W)1T}"T."HTbUx6^983Yzcu_;cc.>[lL#?2cj\E%T42FICN7~dNfr@1r[SV*dWrOo?|k8	Yj,_"E7V.g/~_
o5<H25)TczOJnwPZ9.V<RS5Xh eX*}A"9xJ-*Zy<|nG')YfOrZ+	i^*P[`yk9::$lDFd,s?9/mjxRCaa62g*tPDcS{D zefd&{L\|JN1A,8Q!mVk??`F@LkRJpOS[J u#u#sv/iJ%7:SUXk{K=d2'q
K^NHQMUk%{^AhS6h_mk|Fj%^ X\)qEC~z^z,R{H8*hmhx5Sv
 O30UO`J{~4f!qu\vt9weIMS}j<
~d%a^ C+5.y8/wx$_#d2B=Ehis={@BZBM)3L[E#-oqhhkOXeD-uc7mP"v
8UQWeODlwtN*>zYS$vv
KEr;+!@oU+N<"pj[H0#B,nIIO8>	4gWPdkwGuOb'L\Kgi}#`5hP<uJn\yL&`So8p	>Abf-eZ	L^|#scJiL"ZR9Q7%D%Shm!Va+(A)k.^I-Fz^MyakehA!+HO!zyfhHJR54JVK#|W '3.m|<^vC9=y\[Bx|Ui	N[I Mw<X*@V@h5E1%T
q)jS=+]^856~))02/ 6H``mN!ip#d3
+Q4=	WP1qSy*\M#</bV8c:+I`)ZR {7c,+4}?hbB.@[ZDE.9 @8"WJ<p`jC-k+v$)k?iLn@sSvG75rjd22pPK=P{>Se#{uP^AxX;{zzK2@Y_+d0Zt[yA
h/<BEp63ftwIN:Zn[?BJE><PTi>xu6)S0NIm5fsnr&RrT,JN%Nd-[3rGQHq1}QBu!t;5{uD'DM-wSPL*i"9},3HD~y(3k4~VD7s'E<*NT8az	 5Au!!j
O'kX	@!K}?{go1L2$Os0-.Em0VBwl]VvHy<mfLf_}-oN,Q/LhR8s2 4V9YokD^M"n8qm?^Kpz+@*
'S4F%wGDxP" G_u5h[i4,EY/lYqDF'Nvnx(8.Z|2R{#UhTKS%A;U&#q6w noGX>N8{4d- 9O%W}Xs]Q2>3P|%Uux]S<	 P%i)[-H#@&OniRfvJD.8q!\(l+Ww,V'/.@k4J&"us)BfK VY]|oUoDX9'dJ%t	z}Jv*lKv`JXYpk(X?#Cr|^5P3Mq_0Z&(e6Q9[X$!>I)C];2GS;5Zb&1&@/mpe
NS5d'ul>N.^4	4a?:h=*iflnsVIOk
4KPrxt_K$Z j2VY1oYplX;*w^]A-o({0VB"'9ICJilNS35zX5
Ix6+Ugxa%01%"w9Kyd8U}6Uh9DA{=FumJ?!6ag@P/]X'=suYs4QM
?hQsrajw/8q2?<Eu"},h	FiW#}Oe~e.;m;|~j^<S[!_>x4IT8*8p9F'%QC?h6)JT[a`iHvV_^a\<;5>sb/:=260!,h%3L FvJMYcZuKEPS+C#1Zsyk,eO$#3h#6ohI\jdqOVf4|H<
0=l,*b*
+\2SjaoO,3\Hc29`x|Tu=l6Zp=Z<l)Z-8v5/P,vl|1I7ikIY}]6E4@|AW-|>7HrJ_l{$L*Mlo4OUe67@uSJyt-.H^Lvn}jD'v1KG[	~%D2A^)|F8y30<RS1AG-HES@S
g.0@{/eQ!
GmWDB)	!_S_YwXn\F1\1/$Z.snR:(H@c*z*`N@yqQqB3`8ELP#)GL\2L?KIIO*.%[CW\FH6]E}HaJ/s+5/l{2pV@oJ@9R?_c%T#1SA8P5kn$WFmU(>4'8-B};jSMV6d&X71N l$Bd
M0tn<^{7Tog;pw/pNNG&(19
.e4H>{$n$V$1^WE{E|4K+o5?0Fu5.MHT?U
8'R2t}h.,	q\%7`}IE=*+YJE>1974n_r%N'ZfLL&zrVL?vHW<%\2.])F5|PcCw0L3RP+jw>h}_5JQ[:-|[H@\TryQECfJ[%pj),Xb	e4CRr+h=o%5b\|C09A25pj'K2),GWWy
7pJnyif:4j 6?X. JI>:I
#z.>g8t&n$Q6T^'=B]Cxh\6<JiqK 5kXUmD2zg:gC($o5Up|T%7-UN7d;f7}lC5{t&zYGwAqZxf	>
MCT!#mnE3T3pkWE1KCft?.dEO.!2lO~zGID#r?a}lc[|h_HoI{~u*X]rORQy``?9*d~!If)FD/urO-(HDzp(Y=4[5PR !P}SZ#cuK?CHuSi@(9  {#,]?pRv;~YyvEi4SE"b$A}h~StAb!2F	N>(OfMe?w
eK56 5TL1hiIe3|ZcZzX:j19B}sM7
{,^z'2%`~33~d^8>5Q%f.q	WOBw~;GIIql{>21DmzB:n8VGkRt/Sx$W!V:po2S6E%dyEUl)F
;5[CeQnuOE4/VY5ZrUG4u>	okEx!?wc{7{]hSpe(%])QQ]+Rrq
0j9aEPq=NO"4`y/]8,co	z|L0'F<VgEt&V,t-Uy	;S
drM/|SRl>XMD,JP	K#$U<\k@"#a?Wd)_ExoP[4@MPzr"kRwA3us)mZ
V(tvKMm<8hy	Mil1lj8a(3W+:,tWDBLB%98b?Q?Cg}0&}
vp'-tPK;eQ	Z>dqv5Y_2v*Hwm@_3!dy%icO5Z~S;
^mbMR"lAbvq/ ^U@O5r@fFWj\$)y$yip!UBKW8y9fmkCru"kx!]1SGQeh+b,zbDf&_F*R*kzFRK3Z@D]KdW\P:&-pL25B'&"XX*3C3VL0[-I<*xf#R*CBo8wh/ZX|;c/'t6r@o;ey:k%Iz}v4ky
Q|>;
|guYSp@RWsH
}Q*}HueH_a0&$hYJkQS[jo438jy\;:WUWtKGO(6	<0pTr{_Qg)/Fk:i9X&vPG~~R>k1?V(zEPme<1Yd2^IbM`rZ)x4|>k_!n_].8(^Z"*;V:J#uc/,\8&IRndzS`(+g(8
\Y%V)]SR&_FYb$J8SS(Dc/'Y+P*#9z%n(9Nk;eG@*pXt!xd*B=J<kH{A1IE@Y\?IzT85VqUuv;w++t1h<t{([`@)(#ygOwx4$Mgsu<nVpqh@9,f=?5s!xcEP2"s Z7.GiJVW'y1$4hexVkZcAHeluV,bTE$=<R-lBZ&A5}\wqQLliRq
X@}jr>DMdXe6{eSRXj<
= M[7p~,$	^M)Q49_vBc0QKR^
_w!hh_LLee/2"@)r"CP[;A{,%CVxgeH+v;TwKM3h}i!$cl7#RU47Rd8F7"r'	=1=g1_PC&!}-9o<X]IR!<<B8Q76,XouzV`}0hb?sp7v^X?}F!:(f@t[s^!<	$lB)#L @1of^;*E-8/$U+HW*%]:,y,#Dn@;%W32\$ptz.t>Tdg]bzZ&*=K=R)cGbo+.i=HR|{xU&\gMkH)9&]&kW{<y'^X!F4M)fo@.+WOS:=NZXvzArEGYbdOx'	l.L3'V/)UX%@8}!z1~F9+AE>L<%^7Fz4O]W\x?|
AboU?>Kfh[@qTu^+H$0%Y	akSP$Z7Fe Oo'J7(\1-W!KJ;"-P~t+d[Ez]snxI,O$'y{T=@yl2*VK5'L&g+jfO\C,hSK]1Rr/s,yiqoQx5Jo`}t}|c,>f!g,#N{!EsCj.UsV9iN/SY9i9yk	%HV,37_d1`J+{Wvzl+t?:">ws[z'te\$X;-+iNg_'hnkclQ.fP3{N%:xZn`O/\	(IrYeL)J/8dBi-( *SIApU9es`H 6We}UvONQlqmO:JU#_L]z^a3_#=
GpB
Hp"beKMxo@`m6,
Ew+h7Gu(shqvAviubDv,2w>m%Px}\ih;4JK|W0(Sk".k-zp#>C)EQ7P]3BaJ8<avslEfuMHHx&M$J,>Z3Vn@_s0u NDBw:|d'j`'=@,8LS-wa@bFbCW!0,}Ks2tVU
njko0_b.A"C<'vL%&uLv3GHz}lr:~D2u*z&@re-({=ST|8?l@dAS2Ks3.}Y 2Pe4#n+QQVb=sv|l\woRA+jG9=<hfmdrNU&=zXtwvd]}"(4"1VqIfgAt	l.P9$|; Sn8Ecv_bPY14FQ*	JgR)m	cGb\C,?7nN7SS@t|]etW~8)r-!zM_\	J>&k$e+Gb*WD<(	8=+LL+4tIeX@?C@,IUELH(JI=@jeXAF3'wXSdU2S[E\7@dt<nERP~m|>JgARJ/"d"P9W&{/>P[p*1	4	RSITJJH8Zy`m,J_3E4n'{6aJ:Iobeg%K&>/N|N?2"&{PBEmJ~edoqzKd,/iH^A9G<nmb=/sde_l=^oi }S_x8`wWe',Bq.?2*Pb>-P[u>;K4MCDh/)lg9hX*jA*'(o;)K|@Pr%>Ge^%wa:X?a>CglKz3O#B*/C_t|]W^i*QoLwQa`M6$jE1[(xJD|li/f$IHU+du9&ZSBe{%e(+ )QB-`8/!pZSUdR,/QLe>Kt0	E1v6cUQ#~6O)U4	4Mc)MLcGHNh=T:j9SE%X7Q>(W~*6U}8F-_ikwgS(vC7Jj(~xZORC=Z<;WI!Tc#W!$6;!`J[4m6lt0G\- V5Z6Kh:|hICO8'VQGY'g]fLPqSMX)\ZYFWz>sI*tZ18<#U5xNO+]~6CdeNpaeo1b?6,0n*$/>qx9d)Nlxiu|OQ)%<!CuW*,ZJ0%sN|phs ?PQA{k/"6^SWD>$q\:8*)<>uOX`kn*=(3x&|WL:J
wluCy#X+NlQNKt"0cetEsI_RcNTg&9t)aYg<J=W4X&ajKHX`(({`d!UuNT{Tcfy[dXhcp<FLi|f-nN=RV"4w/,3^\7n$	H.$w8 MbE52e,<$GF:lS&RP`:6"-[)9Ruk43[>561tM.lXgJg~(oKghG=wctn}-_w<59GS>xNaJw\j>T'>&|'+c9(]Y?9!wWhQ]}CO!O	I|lgk](*9`TDo3UrQqByQ7duK>4U	V6r%CM_
0}`1;t):x?W{jQyh}dr D -&fqa#?tKWEiv#oMj`L^!@!\n_=`Q15NB)s<VJX!;N
t[1kBLv7Zz4m=` JQrMKA>H<$DJU%}*RgDILcS&>=
'3o[p=Y!W([W"6>$O#Ca#?%Go>d=n{9?:P OBo9gLKq*O=88<Ap0INHFH<3X"0^>/;X0W2{X&cTyVew<R3%}%;(fkcR5,#Y5Z;f0UP(;m=bY`|Av"+&qB]-q56_Cl}Jdr0PVP\NQy/:ziXDQc)b9U_2ddB	Q

(*	S1nr)J!JZNyoU.*h.:]gw9<X^jFQY n#xEo4EQ!o}6!1D2;kYo0@CWpI(eD7AH8TZJ.MHdN6u9k#W^|D0%9>f^S{ /1=w5"(2HO5@c7v& r7>d2EtZJ*r6iU sqfGyE#0gc.+]HB\^@oSKlj*!B[NlTPU?"x=fjD	>Ya*P:+mw7-e;>2.v%\P~
	LA /IcLI<bSisP!Ggi1#F88B5~iEw4MEJ#_XL((C0c#kV2}?q*AH$?I|M=?kc6AJz.4Rg.G39X+o/Gp$hD{EW,^!5:!^%uJFT dE};yA#P^bBl7Yl^;fQq$qe+cL6q~cjYu.$[]P
O)xD.a@\B[eu1AxT$=	xRulN{A53FQo(t>{uSb(;u.|PSD{rch]C'g%>CUYGh{xJ{;_W2WM<JCeZ;Of3J4>^=kOS5)hJmwvE6OT.<z#Yx#N&n=x	yR'!&(H]&bR8x+*,9Q(h*o{MC^O$LB1qi8;e*CgzqC%?<)@*@\^=Afb(Cb@6]7{>o
u`7nA5Pg28Iv")bl}YICY{'#EBFaen]a^,uukgs'8nW\x;!4ORUY=5m	9]1|<-f_U`x8/nM5J$lfx/hxw#r.R)?u{T#MQTi"a$1ZzO|K3FZX9Ia>1FZ&`IRQ]!2hDaQh8J0I3w\H|]'t8]K-,;5L:AAm<o2M`Ka}@]N)MN`Tx?Cs5hcqfHHc?`iY8x>3=/j|fL=-Rco\|"`	o-_#f=u3=bP.-R.uZY,T)4c*VKu/u@b|'+|q=D~mx5VY*\7tnLCnpV>\'XX[=5M!="k9Y%H-	y)qL'<1nn)%Vc@o(eod/y.7!5	!Et:et`<QZjeqKyhqji%Gzx@C6#.@dFIF5q dB$[;1]'>(GWf}9-94 [uhs=@s9Zrep-
,Y}a;Z=@\^X}st_9L``xU(~`j\b-%M3*`PrMbEpMe}bEA)?l\47C<`;
U0SG57<fo?WSY tvopt38]6#{@5}*gnk(xO!a!79PjC|TO'`	1"(J		-fq<<V|.8^
q'ogF/^`$ooHI4	Q_wUVAdwIVOh5
*c=6tFG-7*F+at:0GF2#BDN|iynx?BVaba^w<1ymSb.EXG#|baMp	`!6rkH+Jyi/L>B`L[FWP~0_JU8t9]eI3|S6D5`tRyJsiK	<gdq6rYx*	DkLqs6$che$P9cJyzs.:rZ\0{W6m%&#9Bdut$@uMg;,*[HG(tXco9te`,JuMNUf[Oj6\q;. K1=Z$l_)A
c#H%:A(3V0A A'uf(*!3S!mb`Q8aI~)r';c8_lb7X7rIdp|X,B~[co	r+oH_3 /C)#K(f.WX-.		p$: 3\s__	TZd&;O/oa1 {m1EFa<<*J1E~lK}h}YdNG1\{-oFV8/?#`o5'G!]ZjOVa-?9d\2'RGFFqz5Fd3:glb>i0^m9BvZc6Bkrs;[ `H<;a]1B=qGO=jZ9@d	70TV(LGi1pW0A@ubC3@bGHhvkw];8un=dGKc$[j(j#+qb	a`'3tP
`,mCWJy>+Cbwbh*gJ"22]P>=h:f tG{ODtZo<WM/A~PJpw#`"NqBRs~d``$Jh	b}S<S}rA;X|h9vx`8)v$i'1b}7VWF5NY.QDJCe$kXC=W>aE':tN}#TmC|[wj}mexAyX]c4QhE YD('#	v(E#/`RPg:-+v$8o'@'AO	Pn?faGY`=@4jvOhbA)+e5Gj1MUup,3+w!CQ$m3*A;
Hy$v?>)'j\D);]/t4wtzU"B3_u;O#+}Myg+^WnKt(bP&Ka$dS0?u`f/J,Ovd)s.%N{2hmo
pnb""/Q-|p*<z\E	<Xn	r"x~/%E5vNVHamwAd,jBwt/mvmTk2X|C	O
N0,Deu%\NA,(-SHW?&J39Jg=<"/#wK"Zu	&Z8c3*XDvea!>.NA>C*^z(nstd3S<M=K>'UnWWz.H}zv:.cP $};KN'#N*k0VFe}ia'D;$Rdpa5n9ye2fNO2_bRN$]u$}_veQ?pZ@,cRC&L04!X%kR;kQ;UU: as:JZV1V7G*2#n~gK%>g]O!7/M;v+Ya+G9=,'XygYn{@;i"|=h
	fLIsVdXU8HqEN<ta$SF,#>?D
{]|lJT)3DAc%RO%yJ/yn1;]g
Qryx0u10yb^n14dU"6~_kUji%RHuv!z\T;ylt$EVBw:,=e7%
SR;D\Kp@o}a}g;(e9AGCrtd#MH%RIXoMlUNzkR|ve4M
F6,^EqWu"+TS8i!JOifLyPB3=	h}Z$Iz'5.*[0=Bp%kQ9{py\[{vjaF}h=TQ),{@CkeWu8[tz}><*{`;=G2aK1u!4wDlop1e;?{ZWA<1b,w -=/4I}D=L|AIVh;bN}@L*sI <*W+4~ZUii>V&CSD\,&g;KBdE<05(bs}8CNd@W40U_Vz{&<S]X#|PAGEj6@P+==PIV@5JY-U?t_Yj#`OY\$/	.o21Fo{3V!}b+3Qrup+-QQGtxt=:R+Kf'YQe+Rc"xnV9 A)1B=H_329&0!M5?x7)mF2@fnKR<nCG3H+[3cNHr:WQd,y9,h]ep*);pz*,>L_tFwGNYq86|_
HN~{n<lGRCg-b_QI';Hy|Wy;zq<KiiP'!C-zzOKhg:f`MS=~w>/}3h]S7z>O)UTZSEv.NW"R4{7j5R5v6AF7!s335UlS	'itZ~,s;!5BP]nTYCu1oZcP?BoWQp\W=PCub~JVF/wJlz2E_NyV>t{xW5:y!\vVa&&f'VV(TfE=G, k-V<oaSl!P5*Q:x__>"3.}G2o2->UC~[NP	15<L#w5C7~w&ZRS3KvKgi7e)Lkb_@*;(et`XhNK1?r1fI+dPnznJ4';~[:"/Hq"_~}*)<?(KtI2^o,Z+Kk,J!zs%7p87gL1
nNUt`GnLNrVza-m(@$FjI9?'<\"1}*FflL@R=M*u"s
jHBlMIw"w!(cbyHU`8#g%Duf]"3\2G|g%dDnO@9D*l:7:alSC[SMtRe[eI
"P}&oEtGZfgm{~0jp$)@zMv[+p-tbs|EbGkVG4b.uY_8ViIKc|Z aU!
MB`_Zz;MhkPEa3q}D[UpOBco'va$|Ti|uB|b*uj\[s-` %l]7-aC{*{-	\;|D+{?]@X$T1/SVZHOn"xwTDpvjW2;"Gu~Sha&u8cXNH{8G-?=!qOIbC^HS#d5c(wnF,OnJBIYRMN e]~Y@Z(E.#oM-BQR!j`Fx
Bh!C6a= ;@ajV}>A!MyU`kCyZ7T
G/z4S*(EziJV=hp/k}
t7|18p~W	[Ivem8)2G)?f=?HLn~W/o(L}TU1e2:Ue#nlb7:)\lDxgaI]a:EUzYLS^4@Jf,`tG=nb$km%D.;zgU$:Bppw_-JLFE0Fkj2f0sJQSh53$x3?&>=l/&Nv=tsQKy@bkP`_J1yeM6TN`qXz
_*
/Ts|EL-&<g@O2xz-J!_1~{t<f@@"?ItQ7p'	&>_XwzSK4Zi1$h=Yg!,kA\)8}mGX]ZMpI5'd</y"QoWo+mw$vxz%PjW`=fY?FsWg_:TT`.G4SOJcaE &51l8
lLHmU5y7r~(YG)3x1
4{>@~+O~V-q.J:	!`wJoa-<Ni^oHkWjlB+Op*f.yG/ai$vDtg_k8lq
-HG6]FP6b5l^K1|.f'IW@$Tq ,Zn@EVbTPzC8W{~p}R@'dN%X,lpKGW;F4>(om+[9}F[?FVbvUsMi+xnVf3;'gHNB?,)	=&'[wY$g/PZ#2J/rW?san.JE^YvnDB	G];s:q>Ue+iKl
2$+r)Whts^B!:qTe\c}h?%qtlI^`%V-H:M|v<qx@A[I >]]Sw#8Ok!l>h3`U>($u
dN4$#BqrHa=-%xqJ.6%5Ha@#^"t>P4pk.eL6*H6,MPfGEsFU&a/tq wYQ::j'-O^MvfiBLp/\c4$Yk^As>t=QqIuin.Bp`M}"x	J"-=Z:aQ0jAb?0Qw)|\Q#t~Ww:Xh8	LQ%=![]"LW7wp`3f/,-|,&ARXvh81C$0,(zp`64
0?AJY(S@1\3K g3DF]p_4c(38oEe^K([+?X9c^x>:`Jj_3B_Big=/+pwFYc?g9_NfjQCmM:CK(atu7
[IF;2$[Ji;)x|.YKsc|i)X|0EE
OS:!j*^xG-^PYTecjJEi`'!x\)*ud6ROIm,-73DW
3]CS]Yf4 	>E+afRyk&b<'zvwdZQ4`p:FQz8V0iIEZGVH	Dh2L=+TboF<f"%,{#D?W[/ O2T*XB2lXJr9E	g>{f3x+K9E*]hv*^vk-J5(S*Xmj"> OS_	
8?BcM<;~3&EDpeiB3T(6z&G`V}u88<(!-JJ,h205B	L^`*CJ_tDKnO,3|y6Y/_j@e&
EJVbee'LPE\"g8jS#CD1JG[\R*<Z+mU/H23'2hz;E$QdR'8[H[(uw-x=dL5 7`qxxLRNu6K'?\G)B,NvtBAD0$;i%Q:T]K\i8^2K{*:(0`{gwB[-0CuZwM*CB%qA^-Hx\Y&J(#g)O@)zF\A_>vy[/dJtRrQ$9xn[R''xY(W+U ayTu_>zb.k{3SJVGh%VbCexvzzv:O^{Bsb;zyDYfZ<rQ(JoRu<&TzfF![^}9g;a*HEzX\=sHJ#8@_]$.-NxDNyb|y8sz	E?(TD'^3MOx0{"O:8L@_PYL$.b:W3c`t5D0^;HZmt+;g~7L|e[ugRDem*	!#_g	OxKg;"Qb70LjwfCk:%jM7<POK<T2K{VPY9SS	WIcM!a8!u&<m)CVb5Nrh!gv.&{=Sc2G%{@w]Q=5>lf:Nj
SKvE#-YMFxV7d:t+DTV6|h%/Xn|YQ/A83 {2/EJf&bLi^_M
[HVe*_^{VM@4{c
Zv*WNt3I!5!!Dd';hmPI	;nRV;Mq9xQeyQEBWI|R_\xkJH"KEyq ;+(Oh)ZZ5@?9EV7eF6&Vy|mVW{(Vz=+e	"o-_
.Ek.}T
?@`'FkM1tPyjF|,t	r<q+u<4[N7v}6AASqdzC8m{.z|JZ/h=1G%[i904m;?4YL|Vba<Q$C:'jzPx\(=XB4H=7"0" 9`~EYBHn"0@cA52DFa-DsJ>'m3g>'*MJ"M:I=0MUW|MYtN^IrE|BKm2=/~oMRV5ed-Ju#'4BTFYIDmZUa<	KI@#"u3sH$%2AH9^YxAez%zTnWPB_#V0rFq2aC|.ks/;
5^z(pb5N[@/n(nye6@	Z}DE`-4SdXO%6a)	ck/q4e_(UB-@,a Iti;@_&Y&p[8P]x<Dmc"$FJ$VHT/R	_DGHVGj!pI"-36}:}zbhpU3BA{]5/$*b}S\
G@={`J[zX5gH(	>Evp;,0 8en(LlQ1P@G/=j Z4P'?PyYA5$TqClcw5;wc[CP16h]:Z"o@{j!`V+yDzc>;6b5@% SEI~%nhyW}E>{_&Ax-VgS^a_;2nlf& NXTDi@`;6E3uIa`zw>^j4{FuS3\#*{V+4vhBK^64N2=F@g7L>lm.[Wa]@EX j
GPzVV 4^u!z*6yzE[ZV{(MVC>yV:e_g*2T0zSyrrsEkL3NWPb.+q.tb%N58X~4~(+ BSTg5&|sBHO'z"-Cf0VEI-C{577@7Al?[gkQbf721

RMWN):)mrv%sH/PW&:L5Gw0nF*3	U}sx)aqv8.jj<f<V@IS.@%w <A8Q[LE$%iR^Qq_!-d{abA87Ox;7d6Np]%vV^Y#cg^G{c Xp>Cs*o/aTtti?(L0}z>-J8RLE*4FTQilWe i7l	{{Y5[mprB>^M^T|^DPD9~"^F`?O&75H8YOpnT.d=]X9Ne;|mG#E
$!j)j\(Rvu+$m-&"Wu]l4_hf'%,miGhmI(w{jh&&r!@.sy|X)M?q.f1@tH&?2 n&Q'O3L;*0vlU Gz%a!>y9'a	WNR@o^A.;`Pw*\Ncg|^>I[Nnp+Ie&uwq uXTQ:kHc*M"')FrXjQ
'(eWiS,'9FPjst1Zq]ZRgCH5MR
q*<qfa8@|WuDMFHbOHMl{e5.\_9xDp@@BN()J`-d0M!b'HbyygrGJig@1CYv?c)_;&j@8Ed&Px;3NVt
RKXi0Qc9cnw6t>@-!cE"c8T{[,y3ftthh^N
Tm1Y?}: Lbf;}mU2HCNL$T.$DDT:of=@"q)!`Jemlt"@Ur<eASr5`5~K)4BxD(4>[\>BU@jWv?#Y,Y	:"KBILkEC!`0O2D."4_FW	_Zx].jY^WAAu6J 3K$Cq0O?zWGjS7X?jie7mf#/6NgvWv7rMBon._n-V?PsJ6sOD|_#K^n~$~-o|
"pmY`LQ')`{WX'&rR2n<i{6v}W>MNGd7?OL>0jJtw$P%1D2aM5"QgD4v%s,iPR@jMfuPvz
"	92\`uoKh;y}%yB|Ql ,Fn>l8B#Aq=zLCS`:=v+,oBGPQ+,^Y[Qp;$/r\ET0ueSgGINjOIaH|Dut#M5#IG?{Nj}W)0A#hS?Qvx"Nhg_)EORNNO?%)x6mh[u1HE`ss
	J>XOj:^6//@6CDZB	TZo/kK1YF
B>J%Sbm%7eZo+\9@eI{_R$6tM.,f K0r*!l@F;!?
d:D<vXW#87kk=rXNE7;:+puO|.5PF"IzF(8hl7`F@^4U__U2v0Q/6}J<!ql9,)TQ9w[T#?,\>WX8ra7i?!58B;:rO,r}At/*|cnn;Ela_]Bj*bB-@	g4vmRy	M``u7WQT]}$"BW75I?}37Rn;Te
1QJZ]o>:}9*q~tQxH?XM
EX`2sRMrg@\xs/f#1ou.{,w=*9gy0H)-n?,SG:?3G/0 DGsHJQk%Jyqr+OPy_4&OP{AQ~4/MA1*30<:<:jk.wh=s7V6cw)JV*WFR@(N~wWy:,7`t*VKi>GxTRwKfyc>AMS|]60'/BjwhANod'2[K	di\<l-ngn#QYh5%SF\g&V|Yf'g<$
3@r|f/JZ8}8?fq4$]G(m_lZhxI4lFpL#;0!1=,0XHdAJ{nUwQj8GfA#->);y%%4e6OGPPT4:(3m$l)|(9T|NW*k0j1!'acNAiiS4^xy#JY,Qu^,x'~VP^nh[cat7+%c(5g?%2m_R)tH	kaL`'7D	tEn9u{}J<@gAq!5vr8<(MO2/i"5%(DEpZ"wMO)<a$oZ][oJt!ui,zi&5>c[$4/$Zg@=QNP>:Ok)s+KlZTmxps{Z3,HJ9:6FC'I
m;>\.UD];13$y<B\H{%d<+N<&^1f0/C[2\O.I"z|Ehp7eCZS]rN6U5"spF~\z2	;?2HM0po i'KJ)Y'<+nMID]q*GYkWlL\+\ Zo!YMOv&{]KsX-&P#.r|y7n[to?.{&+1;w}+6M:zVG{X+#6@C^$?=CmzOH 'psfs<:rq+tp+-%[dbTo
cr)oYS{@P|^?:VT[iDF6^.QnO2RJOe>.:t&$>;%[AFC#';w;qILQbU,cIRR+OuNc4m.Qg1P[{y<@5a^ze\e[1	v]?_x'*%{OTat.@/3RDnHMZuCR	q[-/EinbH~pVc[~d7]-K:PLH.|H4 gz@3X?`AzogLE&xr#rwC`L:b)@1$]\tW`dV)JIvp:"<& X	Al4DwA6-yC,z* NeE:v
PfOPf"|Mg19&
.&2_ywrN
tFAE>x&h*hoyXb37S1S!(HA#-<%_*`1"0b,.pt+"uzU'_NEc)kfkLAg3k|\ne'kIIXJ!E"%,+\i7$X;c(Z1Ux&kHiDYZrw8;Ey_Y3Rd_c		%edE^BVAxq+b{]8_aesV958;;=w<(#:C2;VLR"Zo&c#1'd]P/u\-Q1l?qn4>VV139_Zu@(@Y_vF@gJ'ODl$]~G7}btNGA~(o_e0kA EPtqL_-z4Q!QAv	
GW<2~95^T4@2?lGqH=<Xs"U& )JnOoRaqf!fGb
k_vl1V9I84PUBfMy.()?X(DMcKU:dY"Z^@Y>ff_\0SzvdjoB">1kS3{	W	Q*"oRhveg[:TpgO! 9.pSw#Y&vLHv<^bBUJ3e0GO[us96!34jG9z	;?X);YFPQ][,s@a=.F77H'd--(IY]UU!<f:wy4 oXl#vt{u(z!&b-l	/nl&iX'M:%!~aj5_"et|0@P]%f`p_'\7AE;(NC^z&fbE&u?(0~$3n80IS^o$&sH; /B.=~_dRc4j{>_;U{*pl!v[IU2lHv~PZA	bYEj~	Dy8s!:WQ"&Iw
!',9RS6M:?w^1xa0FL*<B.5OSiuq ,Y{:>	Bq<v$7J`K`cK/Qr'KF_Yp[
v[88%bP/Yj(TNI6(
uo;}Ls7yaKW&m0$8D2/R$"z7@y!~`-.LR	,iQHHadHs<f`y":k7q;02Q82eu1L-;emk0EgTjcKg)4#2A-PX $qn|}QjAF.^30-eUiBx|Ov/'cd1+(cEZ+E{'SO|Ox(NUue=B\:z5Jr
ux?bP_Y(tV KfJ>kA6)bsr)l'>;3Sp,IWHV^:>56U-wg(U/]B(cUDZ6~!+77<$OBK%po;.*o>Bmra?|J[E@JvA}6Y@1"J!r2R8MgCiQP9x^O3PomlNa`)=)9zW?q`1saX "Yz{NKV*8_(*o;pM'
[G7%sfbMCI]g@yE+SO2P[*/sq#W`P/,Ry^<7FXxSF12JtKo5Obl7lWDqTH@tCI`;k3<2LRoak@{E4UnJ-h(;h
Y5FYJd5KaEwI1|EHpg3w+pU.I>V`ugZb]qJLg$AS%&Vhu^b+9o29Xf9jHHHs=O}_4S`Izt!@4a/fjAY4=Qj6jf\[W	fVd;hHsTE^_Ee	O}kP4R#{fo4ntG{1x>[FH^KC[Wv|t!{#ky^m.T+!_Q^+ZiFI,eCSOnZ3rzdDV?rq)1dF2fGc32~}@P5	F}Ym5+Q`:S$@+do`9 |7LfjLX+yR^UD` lhl
+S{f,7lP9ChC}ir,hdJ%i~MW{j1xeC'28 K&"% ;iB	
32MDjqH+Eemq,_V^}[
~<iXjU0>0IkUd#"9 bqWooR6;.?	*k)eBVd	YDD+3vAzoS4$V1s2	b_?^?F2Lm:P\}kta5v&TxlK@OS#$cSM@G8BL:3N31FY^B6!6I^/EpOS1Fo]:nY{sljQc!0Sv#Oa}uFS1uD@3&p$ .J5=PF%\Yg"oBMJKI<Dv|oaK\)[u.R7E-,<LGC7)@n:+(u)SHpF(AzduB;YU'Y52w@ec`x"3\%Q$'OAYsAQ#p:755@Ypr_,$}3}}EftHZd3$ZTY\2~dsa"QbtlOAU#S"qBwHoVncYUme(4&V=Hlr*R$bQ.S2%iu!B!m6k/O=D	1YM`Fi[5l]\YI\b96*QKUP5'
j]3z@!^vE;,$YX}~rL$muEj4l85RoZX_}:id(q`]	qG@_!5%<=5D)}}WI$7\6uho(hC\.SwlI^"2C<k$r!Q/kSoa*!6YgfH?}G[2OEadA$ma5y0{sg$4K:Zz/Jtf;XO"TT-yH,K*9g#H'\`h\JlaBH&gh%JmUu[{OW70\Me)PlVFCp_`_IsR):?1Adb,t]Xgyn7)(TU'9RBgUP#g>*|AXJQ_NenCvLs5Vcr7,rDzW&RJo M{+3et/[%L~}N A7^yL&P/jmR/0sY!tnk	9EbeMLL1bA*w1\HpV"3A,QC~V	`n={N`!k*=b>U ,)*SpjkT.Cfa+DDFl@n)CkJuk0fO"sy0iy!x@/P-N'> T6i_mfZ=hm1{<d;-Sbhux	@K`ZY7N1rPH-)0Fj*VDbHMDBk2_Yw:Y)GOKR)O VaOrLCE0=ueAB?uHReQ2Qa!},s+hqO'jtav>F-nc.!["]_{zj"Lm":Em02vDXt_W"~v }}EAVATLZ,nJ$dTvxP1Y /h/R=EfE.P)QkcXmP9$2<]Ge#^S+GBB!!C`to_I:6T@ qX,W(@q6uu\Bx}e&Duu 7<[eBYL%H?dl!C5lLl/~&#'@g!RijdzKuI@S&yh:sCneBBE.N1.P;bqxgY?-\ZdbC!5^<0K_NA9N}t8`ME^HZ1~T10Wmsn^8%+ph$9%*|#7zax;tD-k .3O/&]!'s{	T%t\k{ma,[isyuNs\$9j;<tE
*Z'u}C?0Z-x'!=g\Y6A9))#8	F63hiR\2#[S+.aJ8P&qJ-XuCxpfw{#q(p\>g_C`NC_=1.&0>wB- hXW\v^c|[EI>M4]vL01uH1_SfUo8y]cTPGJW$p$;Qi=|qkIfU.N`wt~c29K|)-R*D]D/]UpDmla8`YEksR=,Zxi]&I10aC"=L`;2!,o'_o[bm)Y!leg+5?%>E7E#8yZjc-2.dGDT8;kY@;M1=L_E]0'\T,V~vY(R^A%ijri!0dg_g-]s0m[YBwor2 I%DMf1&1['~`BhnkS&tT)'5Mq:*{lRv80iSTZhtPY#ng+Y,Lzk1K7whDkb{\E`)5&U>Xk[ey)ApMO`SbaOX|_u
I#-@/;|Y4Y2)iO7	)D.S$_1bN8?Tjp$sb<Fk!2`Vd(V3sf!Cs?ub~h9,<eY7vq.3&'R]0>F"r/F%rz|$$7eBmzzt@pwe[hVrr}"6r"C7~z" J.@-
*Gn)<GVQn;.=NR(g!@m`m;],fuC;^3J#_H{y~~*m~CSA!}B26\gp,1^p\B'$CUszAeaio)Y't" Ns5ytGxm\~D*1[Ls%E|6t
;VkIn*=ba nz,;|Vu%+&PKt7F-K[WnEvGSRo#!f+iWXn]4}(.`6k@hjNqj_P)p.zVzj&bfJ)7<Nk$4
AwU=5bZ[QJ?bq%$PQ	9A[wpXgSX	T0*AynE'm j!zyL_> devB-M5s/j-+vW\B-{;.RG)4]Qo^&^"0M3|L.2(<M=fapJ7)7\'0h_#+X~a|"!d;+hyAs5!bI|UM^1{ha~NaL]k:WKJES$al6r
$C^[~CSdoWwerr5^PJl!(N8#LZe^z42?~U1"W]c"{!E!_"c}sEC,n~){n1w=C.G7fiLzV oo@b'pmb&V';7"CuE#?Z5d;R~!`+:O0/2gcQjP&^X40:lRM#qT7CbnhDD>;|dF1*SeV`N}\[t2-"8AP ;.pI:*/nMk_ipT'%!, |tc$0|lc`E4T2`XjvZLo4}jx"=Y|cEWtf!EZ8&!uzJI
	iR;Gbzk(mOa- IT
M q8|RK_,F,ttV%0a'a	k-%r1gu'nTUEp(tf"X?(cdyq[Wc*@!Z_+kCi4Y4"iJ%D~0'Y3SnCrb'ZdpPR}6@h}?y{b#T4c"ZXIYX(1yy^GRpjeSZ{qS/
ooBN\Y/0Jp	AnNaLZ9u`+a\-9"$k.gU^s")Z^v?jQ%5gW8!!UlET;!&T5We!(Y:`kW7O'$?pXHqW(c"
1sdQp`O.')]!Kf{w]`&O.biFQ:VEK9C]yBme2eRvzVs~AZJAx>n8<7#hC/)3rR`K2M?m>H*cw4jvyQDh.Z70Fa$on6;+fl1XNIE%*)`Zv&QwGKMHfiDmNz3tvVb6MYfR	ists	7`kvO`A89y,F>I+P).hwDP!v2x8#}Z'aWu@DcnVWtz?.+fRBGj=&r@p=8K5x'8cd&RiIC_fN8_o)RI@	|DJQ8}u0ZO^,]G!::D&U\8`wjj+IAHGICEw,X]LR-1NuyyTp5RC.^wOP8(0S#]MTOx2h 4V#*:rMY{N#Z3a\[Q0s4)&{#1l,SM3X/(7hzy3PP#^*%[\EK5@u)Lo w=r1M:&2mu(UtwNU<g"t&v2\Y#Xy'%mxiXD8i.=5U=D,K@k^-[JBRTA.QlX9${=1OfCN|Y[PPrs~@"D<Ce@tOFMqlv.Yy/;m@r\4'(w!1MG	Yo39?QPU~M}LB#/Omt}#<d>[HTtw]/mlbH|dSg2~!?4~'/}X"2@qF-pQ!^9?.}]qEW;CQ+K{X#=--0.' VL9=C*96)Z70t'H{{dz!c;jzvFQ}|^?0327_>Xf4Srre(\6YtYq8zWL[BN02(Kk|_>
HplW>c\ &-[3MGq*[;>V_Q>O11[_vN*.E<uIwRkYMLo:Vvm2"s\
'.BKID)+_;d&[f;{q/iw+{OSCY}cF%kF#kKSa
m,#-^1G9Wi/S}Ng,H#t>M$M0[J8"~qjpL2y$d>;st{7	[>:c#EeYwbp|8Ka^AhOPFz_IDL\bpJ^(SPh5by:5e-yxC}	AHhP{W'gf&V9=Y-`I^}dWVWsai~HTj)c)?J1z5FUQ#bL	W_`l<P])P4*HP36/t'P`RF"?9pg`#Q`	J1I"_Zlc?23mO\.6~VCeM#4f@	Oc;Q;uYfzo^uskZZVgv\V}n4qd0oA-n9e~baL*/*56]/e=2s,|{s\6r/$wJms4dEZ3Nqh<Ua^xsob0nJt#S5@%C7gt^`A0db+(6-a>^$#B'1^qbB	xYAvc{.S(JRog1k\)SP}V  :w+lI|#K?ZsJ5pL?;iAiyf}61.>/~o':6EO
!9D`1SCy[-7[1_zTo9H&jAiMp)>?\*>EI7F@Im/,=^$oR>z7/if{jP,x9i"(8JAlN\NC,n1`0"Wj[6{P{`5ozb;eVE4~e>,s'4igN+K;jnA/:{Qr:{S@<F#m#m\g42bn#t\ ;B|$li+4f._V) o"(|pT=1l%L41,EsdSf-9>2Pqw)<RsVP`U94M05&7fU@uHFekT(J*|.F>p))ZHH#8@KO&IM$Q,c'elOq1UY/GLnEaMU+W<;>;^:`g9IZ.B>q:1V;z&ie?ArgUM^^nSO*p>=Z5+tocd!' =7ZAX?ciAXE$O?cXsSX?{~nX(sE?+Q*mu'eV>p?7'Wy2gE whFT=oJ52I^!,`x+(Mm3=^>TZ/*^]y~SL7/p	6xu8BQ&rM=han{[")t]}I b2JFBG`-mO|UMl}Dlk"H$"]B<-&8n@= _6\9RC)
abBFiZnG*J_YQQ
ryb	P<v(4Wu&9AD@sBp4g<f%h03.%HCf\fo &Nn#XrL#CJXO.#Z+~pd0tosFDfdofmCtL>&[&Rn(7q]W'c72.79TSspfe.r9b=6vG6_DgNOVwOdKg&|USz&lQB&3a".rC*[xZy"k"Mw[jr5-Pl!eZ2qN0/V:_W-DetT<pm_]~3[,A9hlo+EsfVL?n+7BSkhp7]qs-C}ddt4D*s<d*!WWt?wBDluu?H[ "D0FV<!N3aAWOh3L&ZpaFw;SvrqQ(3MqD.V
cc4+(xI5ykIeBdo_+*=p6$Umpob,Z:FJqS<=a/e\WX_Hab/R*dv."vZ4E!BpnS+R@('eI`mo?;4zC|$Ji]
v:q_	
R;"BD_ywpCTy#O%v:oMs7#?n=~`	?Eda?"F(AD:GJWzZE	j\b'?hu2=
r&{=*VEsSn|])xyL[,L;]ngg!hafCLo	G37N'_`1 U^hS_rehj~{=OKwHj`pa:?bHS#hgqF'XjEE[]bprGwFZ-Hbj
s29/4*1% IC 7qR'QmR}!ZV'KoT<ajM`>' uIm
xcQWiz6P_:55V*LJktWV!ajQ&T'(R?/w^,!b-&Qv4yWPdAg-"RVCY>a>@'TnM
<K;J"8/=8AF`Wt,j_I3Fz|*)3jtTDCu%nct)F|H5?yD-u9P=GKg3?[+[~Eyp/ym2l8!38aia<iB(ef^Z[i$IhwQA	p(-ZZ|0.~}U|OyXL)R/`\s
U\HRt,ql0^$`gTV\Q/M/dD-5>PztO5O!qvYMlEV)N@#wo)=W{Ns6VGRV&s}UG	]' ^Qq_~CXT6:}iKV]M-jv}^)46=5/OaBt23Q9t0cj&B`f3c'lEai$
y(nECZ59D;W[UJ&es_DdcfnC-H$%@p(y0E2ib.;vHpM4P$\{Z	o*#$ 3{7
D"4)k2t;$o1 EL!6DpgI5VsgDTBtB],ooY]Fv5|E:b5k<uE;0f3`6S.B+,6p+%uRuN(io%}'|oR[2(\M4PT(Z^ =J
=DBM@Yg3:;gA_q|If>>jCWc%-`quQ++D481^.Qd^9"(zjVsBB@>47A7&=!4ZYkb{bE.VO{YTz9]<gDE)quACZR-HM(	)
J^tF:rjS+<zzl$h|}Nx@U8,|V67%2if2cU5<a/H;BEGA!ul%H#:3X
b,BY9TE>grH@$RL_hdD8K'fJM&M_s{M!f=9nr,NwCT}:]/B3>/cvAJU[/GkiI2qF3cZJLjZFbnSoL$gW#vgWAa?faa_*Ofw::u\LJK{y|Q?Y),28mhB!SwZD3a([C[|NvOxC6VXfjK;j)|F,2`G~M?G%S82j-y!/Ej6?#vk	&6/%|uX%k@8d0|:pxY'1a52`|kn-T:/@4x',*h~urje-"P9n:'7:XYnfwzfQL+JF)[dm^M"Yg-^w?!_A&-=d\"q$C7&b'}tE_1MT<P9xC6B/u|@GN]M8H!5_#]8!(*BV0CQU*l)W|s]m[`gX6vqob?W"@SV)G`aXPdqF8I5V'qd?uINoyWy;'^cfg)G*#H-xsaG9oi)z_4ypxnre4WA7:Ry1zR)PBFbwd{Z<S6QffO!SBr8k\M5zdxv]zl=%rEF(kD &~EU)_5zS'n|PH1UmI/R.[1SG_"xuqHU8y:G&h3XL?*AHw@<C}^7;ul+(au@UM"*0}W*-`@O%p-cZ<	
y_hI-|U5{W96$^v5WgA:AdFM~N4q~Bbj&PxVQUE~O6qhj//NS@bq&yt,tlh_yF8UYJKHi8SmJKWQsOz#IHJuZwu,YG}d4y8Z%>wx=D#%"R(|VS3.w\^^3g2I}{#T~/V )S!rz0@I/"q"O^	ii?{oroh.6:4#~!w6_N^@wP/>.4]Sz/:kPFB69384"YgmIdai*>`jnn`?N M-^^)dCAFznHPlg~<zSy^644BlE[QFzo#wiRW7|crqV3t8sR>0#bPuUF-sd9ul0GH	-a"UX\{x{_<sSP:IWIYi]Yf,+EY+Jp5oLS
-D*Z2PF-1g**a6zBT7#|_-d[/<C+OA%dz54f$-/\5$35#v+kjx$Sf!
DZai%=)Q!@)a}QpH^m#alTwmO]Y-$SNh9b1tTBd+Oa-~JqFl}X/n?VUtH-C6:5#c[nH9qYt7F;26"nL%,%a<m-:$UdG]T#`o)C6C]hBY_t-' ;A|jY^~`UU\.\G	j/Z<_|C#	,/5aX1IoU	UmwCb>=j-oO/*,Rmg'7ZFUY?0ir(Y(]L'FduAg>PSobOeO}&`t^(6D_8^VOU+k9GeuQyn0>+b-"C.
;F0bNL2Wo()!1(I~#r;T#lO*j6rGkN	4}3]TO=0}XE7r.y#^iA=Mm;/%`|]u
C1x$bl*L6n!|*1s!%!wu*o(bI**{Sko^74CIdi9,LO<xeGU(BFQ[t0]fO0u	dnZ9V:g'w1Z4nGv}	AkAVOq--s*W0I{#d;<'uHh-6sE4-cc~0S(nWDT/4/[j}N,_0l/>Ze=d;GJ&,/@dRTZ?@hZJWKm,dK#Pt{1aq3"L{{r+kw?k;}5@)lqie""']~Sw:}l>o*!^F|F:gX |cwzl@F{/#RcB%\@BHi=B}[^M<*$eP
[b4O--z*9Y%&|@n_Jao.#O:j.1It.6IiDf"Al;VUbF1Y].l dCZ
n`c\y-6#97>=|jp/"!3m,4K&:p;*nRql2{ G-\(;>&SjPK`sw7N[2I0`=g\rv+.46#=<.\eoJyH#I8X~$TZ4n=(	R{Xf$0>/yB[ySfhZ>2N6iK$M9aL@I'.&x1KA>{0s;Rvi)(N."t0HT\Z)99kHTCoul ,!Iprp_#}	DvgNCdS[V+2XeVTI	FW:bmySf
Wu%Z&3XKM{taHQ~{_^lAA-}F,I9_Sk+g${UKyv$3.#oShJ$vBfq[@MzFW{Zec$p2I+tQ5]b_l+8ad<>m@{4}V=^%TOwS]q!(D;-(x!8%,X_Ce
n#sl%_1:m`j(t>r )}J,]z1Y^VmlS44S'<BNuKg4!s?S|;SG#CZ)BkUmTrWd
2:74YssSg7>Z(S4W\C&8_<.F-/i20as^bt#o6m-3lyAH\5T4\1&=Et0djpmM.X	?]v`	}>:cIq]tP\r]NI^_Zn?/E=@aMXvq-cg?us,BEf*!7$ bBIim&;m_&L&= lujj4%j\#Mb>)FTjX*=@f&1jfvv&dzA+A4=Iz5n+Ga<-F4_fx;hBmCf=iV%HO8:aH%_?yHe.B lc"
:.?Ht,i<*JyS.b3Cc[cw/6nS^A
Pg=3(Vdt?rtKcdT&T
")RE#wt!(clyf--Vp.(Uz	hK[sP
DbiL2]3Jh:9Zc#:!8/Odw6/V]r;0hwYAZ,Tj8 jO>,hR%:~| 72BZn1]+g6lm('|mMy<mHAL"@Hmc~T%z=8zUi9O\	f.0^B}Iog%2Wa3uY~ONv@WSr<HC`
+tB;Rn80/<531N|]-Eu9^p	gXB/JaY*(xnc1NG;|wvmr$LUJ=Nc8}Np<[zzMf(~C}HE8+z>-}Ky]Ics\pMGS`sK]3	1-|~	Huk3"w,Xw>>k>l3p("ZYfFr.oUD*?{_r?+Ewz<w\8^*H
$YzgBdTCz[M	ff`DJgR+=-B++	]R1HKtAcFzVB?g6BW?8r14e6h*rYFl}k.&L@|"s~	'QOn0.TUz"#IA:ts[-Z*Hf-u0[bF6-rg\ntJE\3k;j@%c+9"ta~>^QfCwz1Y^7Ub\$S9k0`nklx"]6Aq{|zoCB%Q4^gkeEwP<hN&A$aA%Hmm
&?p91_CMPsV|sDF<9HC@wn:pURJ>Tb<ItO[w?+E0jeseA@F-G%62,9XF@mN,<evr]G>i+aw}jT9UvM^S??|9_+<n:\:Xy?0`,xP$2=$ySi
s2dWKH@q@,'?lY;M
[wOZw]0xU%Q;NWz7.u",9[	ID}BM7o$PxHWPpT_=De4c3=:d.~*jM779LjQ|IR=WWz^hiZ!Ja,xbjIl*xad4q2*o<!MaimGuSa&Yxob~F?XHt3"GnSi_f3Fox6kk	`XPq!&obAC)VGs,s#RMo<.7MH\6Q. jJ,m-Ym9PM+-iIBpE\!Kl#+U0J>Po'EZ~XPb\JD6ryh/Hy:
V\k[T!GiV;6	2Cau?.-R+&~)y~#n8{AFmD3q-&.HWaN0a?h
&n^IRJ@\(~5=e/1T85AA2lAToK~tyrW7AGGMb~0R2Z'c"0P J|lDp\+@-'_M9XG}4y|2Vl^DUyGmKsyCH=H=e$	D	KP`.:}@_yF8bH|9)(!s=-=\oHV&U2:C$p*1O$I(Vz+g?=8<DR&xo:4wG0}9Sw$6dA2vdL;H$&7XAyW:-oP]f`?s-y2|e=(km%!v:"07/Qqm8;,aD:Xm2*8s{;I5f
VP]$8wcC1pxXbZdr20j!_`qu>]Xaj^x]R8-F0r#pU]=8d0H!Ek:#-@%gY"-M0h<:8+JjM1Ign(
S&"jTy5fHS<(X)B[0kV lxTz$Xh2AzH#d#Av1-:C#'WI<msw]$E}8t|>l
lK,|!IRVTlHG7GdV75j}?ePa(APmEqYdfsEWv<)`~tUVi0I
Y=&]/_m;w|o
?Uv#{oEVBV\-r#mF@sUDy0B*~2|?.6OI}P	<T#G>|84ckwnHz?`sXQ)JdJq&FYr4a&{C8	YUs_|fP_Fq&+3~)rR{gRI<yT.0I
\=fmX^&QIRL&#$c^~62CcH4i?!]%rFXhNB0V03'z>h3n?wH;_g]nA=(5r8
*1"Eb	*U[Y6;XG_Y8[<(Iq(gY+<3In1iB?0t!/:L!
bSmrAD^,t!#J.{R]6n0!?$teZie![xiZ]Hk<AT6Cto,i108FlbmY/g:X.`"1b_c2b$6LqT)+
<;`
H`Gj 41=L@hc4dahV+<?Yrss}pco3o+h5[S]*35@SxP$2s800gUj^oH9Mm{&^aNn4sb\#9d~m},Ms'hY;kwM0Bq"IZ=4?VKT01~-\Mf'}AH;x^"0@aHyo'f4Cr\a\v9/(8(!?hRos),R_]AXUQ4e[9`]6Z@	{WmJ5d~V-_D1UR}d}Q|Z&f!D6[kpWT}T&(,G.brVjK
VEAy7Ar$[|LB' Q(*:p9qo+meB^*m.L@`-WOur|S0Ky>Fd@P759=s1Xk%.VSRfC)O"	ew{%1xe;_r<:(;7(IxO`BJs.d@	T".iXfOj.Ca&;b"K3WOkc@i	
o]Gw~EuMoiIkN/@u8{E'L:V%@NDXb#Yv*y6->bOxmH.,_v2dcK#WO5dMul86zk0VkV1S,))A6Qg*Lp&=cRi(XSH?\AaN$t@g{"%+`xJ[S<&yUUX?MGg1~S;*}lDh}X
	mH#Tb>k:SAQu/p8CZuK;8J221_A/jZks/Z|Us#P-J\YYn]A:A{q/:+L@<|/i;
Rn:b'hnK&xk_hG*gB6{Tos[*??7*;xRv.
p=vr;aZdys@Q-"<u_Jm\W|]c:xd	-Jt6B I{la&.@@5E:9Hk9^Abv&(j|92j-z<lSA!(I>4y(Nv4!t.=dI?SNBHJW"QS	C\3j6+SuOP;PH|zi7su/]80QQji$70Q%9|"2W?rA~}K3'4Gq9}dmqz*Hl$9[D/5H
'yb"DU`x3l}XNk1p"wW `uh}OZ{C6yr#h&dh"B*{-x4XdvI}-}7^r-%R4'5pn=sR *mu4n$|z[J=5Lf3kg>TS4XsF'&j?a8WFGN{. rpIgY&)Y}	<j:*AC`G$|h8O'dE7Y>J?lujBm.>Eq+W4_{euGnXF-gu|{gs	1F"c8*u`unXNT|9xFViX8Xs/u90gd)hsc;1cu0N@u3]N66]n;G&W]:tej;p.Qp9XfX5SgM?S"_,^mTmRhrn9(nRp`.&`3d.8]12@71 =cMIU*O4O(K%AGe]:BM/6;>Z3E%0^xvUuG1I/6tF`[zLu:qE}E!~4X$ftg<=
SWoUK%KU^\~7+Zg.;15&4O2P4B8Q=tJh)TrY2vg>3[^z<T$EM2xk:Q\VtpG0ayD"Ks|-R,bPH6QR`LyZ6bL	IJjC$#	@:Q+{l/{Y}I*]k.MW<$NTMSIy>}%H<k!)BCj['@ko|',Ucj70}"_sAbT[Xn{degac^3R:x}uU:~)exEEILnGNASQ[UsuN9L]|BGi;R^IXu>NG	02*k\S)T|D{Qx'I$2CZi[7G)PPZ-yfyA{thXUqtW|qak@#v
nEUY`>F$A\My\]"?/`/XDo0:@.,(.L=L-Ke+V&w=JFn1Usv<1Q$kh[/c7eAo4uz#,|&{iSZ>#%Xz>X?TjXps$~IdpSC`wzE_D;Os#Cf#,2$.bG_:8d*M}nl:}>[/{3jg=hh7E@N0o>>fI>w}%;evE#f:SiWl1,\?:[[]H`9~K7qiSR^:)55n1z@;UYFg-}	!!w]Y3;B8&XsSsU#$bd0eq;2{XM!Hv^PB` `xkKS$H#4AZtudt(%ccSz	TG tF @_>/=!R{x'J!)#".&=Wv"g@yzyUZ:.P$qte,b}L*jH&?YN"J =ekDb5!`xnVHXzEdrsF)ynZ+WL2Pt179?E=m&#[5'sD`)C\y+zt60)V0^,|1c'gHQ@bk$Mv}'z!>h;\bq+Up YS/)T,.CuEXX|j f@+I7z:i:LRzh;+'KD5>3cD|Drs\f	
.kbt-7mU">Df.&qE_]^Wm7zCu!^u|]kZ2ePu,ox)Vi]^$:/ BC9Tofq`GoQ`	t/(
w3e^F@Wb@PlS	EC`SOFv@v7&j"(%jIkORJqwcW]P }G"`)O&dt%.@yJ0`UoVSCysf:X)60rEX2bE4L=~p%g=<:=BXdkWpV=Cs|fr9a3[%*d{NRd/"!IqV,9u,'7:>HFk}1O0)3(M}uDy>u^tp*42HitE!]+7up4"OLx0%C]X?#8z>Dm8vJ%Zq|$(D;jJMvMx	9m?.[BhLG]%N0424QF3!+OgO&\=)0whV]]*fkY]Oph)ZG*(ceKUlj6a)2:[{$|_	+r^5YW3nE({@	0gM^wp 4O{3A<gcmR$*x5z%#xR24"0F|dXsLauF^&.~X]|g-nz$R-xSF_e{8,x&r=zaxyYRxt_mB%1#wo5f,bS+52x}`J\>8-}:~@c)p,5IfKNV=b>6y:~bRhHJd;/D;=81A|jh#Y~Om[H5Qr2}R+8)Z@G""4-n]@:)eIA38)4g8lhGqM;h&X;)FF^-VtUYd{tbk~Q,=H^XGwWD1Ad{9Iye_y?s,=Ti164kW)V6s~a5pyqG2=ieg@1X`l+38'Zx|rLISjuwb#]85 7u&g {x!T30QrUj&^+gid9q]+T_6jj.'5]KVv14<fuWlsjZZb[;f|:/I"P*.vQw\|tcPM%_TT>,p+v_c4HNiyGQgBnS+L/SLZ+P('i3FJbE`'a0J4n
MIH<GL-_S_K#SK=w_J.xy_x_E{}D;iJ9mV[WW_goP 1vTrFkZq.}s6]`Ac^n#~=!WU~
~^r+5'=],sYny~V%v,]fAD+'hu|lYP6+mq?Fc$
o5_=|rp0'LQ[]C^h&%V0HBKS9P&=<H'&bKk;Ko/X hL<GD/D$&>ZIJ.I/EF@*fRXjTI=z	+?MMu?r@bGaEjuxVs`J=wgR
KppVU5RT	BHg,Y8Z-UHySU=*CaZI-@H?3hmDags8`Dy\[LJ"V$`Ka!G\=2`zwrV^>w?9/@W2vjD-T3<@{g?;40jtNI3F_q(Pxk|UlO:2>.8^^+`F\2*t7x>t2Y`@/(4fK0om|5Opif,:|xeNM35rdve>ID9P%5}F@H$O\J{i
B>_4qn,yiP6|vA?dN+9]]=<cZQx>kuwb8P\.n{I5]a%YYK:f.V.>OVlV(:|}d+
}(kr$s0]gt;peI-X/1+DsmFuqW*UW1rzyz6FlrkAs0K7^Z/ vM%,7-ERfuAa>\:01l.L' O~6(b5~j<XM?'%YpAj.t?vx76r''17|~:|(	Q3Bq$
u)L"@9*<`&l!
:9d[p\B} zJSz~QiQ"vB{6a#_3shB!Z:xU"~;WHspC\\)S6goUzD}-4Z@Qpqm;MV><[ZL~^ziqGA7GtR!83I1d;=ZNc1mj[.p>_D]Kuq2gGPC/vXz4&cFL!'3%5oQ.G~v(wOe@}T;jgf[,uxh_g0rfy<Of[P7h_60^$u-F|[:;YKxgwW!<Xn|%h_}KQi=;GXk8eHgC<'sj?a0]deejUR+8iLUw_}-jK.39RAg[*R7yl.pW4brtQ	O;o~%d}T?mvjfLa-|CLV~C!|^d-FlLjR,!:GO{%8D]Y.[<iOvWcmKeIu7{gV"Cm6E:&$W#pp`_4[%>wVvGoa5C1w K{)"/iW4os2bYg680zlJnt!{kJ4uq$R]5QVeJRHY[,"]BHmninQM&r]8~WfCGOBnKcEMYX7!e^%-%IqR6 G'&;IZ$<;cLj@']W?"k8Q3zFOtKU7%tOxdw&_.3YFBZH8o?>X>G-iA> -P!~.w! %%f!loEuDeRN7v}K,J*h5^Mf~RbMz,!0V<D8qM'> -X'7Vf~^pu;tn c`d;|w.c?eE9qKVI](>}e@TvmgY/2S6X/H{10jEr@@I%Cl9RK!Vy \=G;L>m0;ZI9NZpGV:NfALX@(L7=	Ye\ic%Pb}!mhpqhFg:NT# :6;|,ULi
SHzCP^2\%,p&[T/8=v;AHyh
&/<;"hD[M6Cuu(up41Iy>Ko*C`kuZ|4B5;(f$3DF+Ly@aXZ\1Duzv?):_72rY}BU9/dJ^.w0fGz|=RNE<
.l'x*]d	82C\m!=S=
X_v11)eZR"M7<e1	>zWsdm?d0rFjM.ev_4U"(-*T=W6o8F"H2Er= FE`%lGi=tuQ	[!C(A4tD6PKt=0?@<)+zfW	nxwm69m1(del9^MLe#UU RrXZYdfE3ylpHL%gvENK,doh;mP.hhi MVn95xS2SWvpMW3a52Z9HRtzcCYvGKV	\a,Fk-"Y!Z<`[Edi'e2@b>O_Z:|,TX%zckw6+\2Cni%|<834^_w~Cc5Ocg/k	X,xQS,Np6,Oy}-RTDm;S5d41
ijHg3{|ZI<kc5r4EUL3W](<)/FdflP|E)3-FZ:r,P#aif|RSG"8NkxzZ`f.rWZ{L;KfGU	eZ(-Q=?RVNFLOqb?;SPmHv7;U_72\G[N[G~WQ-T_JxiRP@uR.M&gt{B&V:XZm9Mf{
Yv{pgC(q\+L^>k=\0HFEn;Og9e20#_GH49T]q?	eWE?fOU|N,WfIl$AV{fI&0:I	E'~J4uy@rQD9k-eykyc1^Xh">[C,tQE9b7{08z?Z-SW/pfcihV}RRz\!Z*V;+GgkA45C,rvp%N+V,U.{V^l=zFX,|=K	c6K(r:.h]f]mMN&+W{`TfEF3;4OK?X[\3IrDrH;ep\'}!MTQm3[gWW'4	ByPR1dbMSp :'j8	bTC*)-@e^(4]"R-]<o@	(Q^PaPYrF-:Z8|WA!{PUU6;/&|]L7wAjFNxgoF*^a\$d%JwK^NPw.%?0'UGH r#B)yUC,.<)=t}H}3&cPo:}<~#!uxxJ"*$!23$N]Fa	c:mQu;yMmpkh3wmhj)z!YfP:aVCHm/|XQ5Tzo(N(vi26D<a>gi'%mg7v!qI;0;2yPIkJ)w?[X3z2a?,//@sQ'*-sa#4
y6>hU%dw$APEIpabKJ!1Uk#IC1|F>7rtc\sl)F5k<4hY3t5G_1szf<Byo+O~Q@2H<t'*CVvXwXB94KLicz=E]N:$"tlZ3?r2jx,&![FoqkPiu'wNl5J,d"kO:?c'(@L%EY.L%^-E{']d%)|Av*W*FnTh\-/D`lamU<Xf^dbj&9E`Y"w4RF=)@h{a%MxY$orQ	^M@N(_t[m
q!CW6;Dw`W?|3WHVO :9M
u'7!C_|L7}Dl W4(L^?=7li/GlKNOY+'i*PTmfytKFgZ_AKCbkWu7S^`W?Tk/a?H1@u>uEO@BV'Y} mOODX63]gb)e! =&/I*$.zFl1?$o-k%x+(h+^2i/H-4{;?y|'}VB=`=Djr	WIkzw`)$G6f%FV,dWjh#Q80|rV*(9}5bWrlRCeHC/h0"m'U"5lpj[P
	@` (-uaji!+P]ryk=:J,*@j6SevV>qtU@O;i(~@7JQgp{'L*a_<8yqbtFhM[Op+u|;A*#U;eWPpE;iy[J@@wyy6rBd]f.C;@njW%wP<TqMHgrW|i}\!xq?6m<jRvucuL@W@rG=.q.-["siCA2JD,:UD3_	bi`:owRQ$7J0\,Bt3xVR4aVfu^'/e]x%ZY(]#.e5N<-AZ|zEUM5}NCFuT./P]:])!#,@\}/<y>=Qdy}e0F[9fKS} AnBw-Ed'XUKWlY'M0|#nLjr_~Vij2\<`VQs:O-rT0;V7(%LG0W-OQ^L&t!t^FM(g(	&(tiro,"*;LpGfMsuCw13BUKw!-<.Wh'/JD1+N1Rdu;z&nSG,xC.Nn/[Oe}%*eoMM	,L^|{&9t^I{|heWb[_be8.(/]uca~&\'skU 1'fKc	'saS
##x&*GOH&f)b}pC[mWp]>>&L_BS&{FnERfs5T#Ki`I,F9FHS,?
wdv/\HxdwFSl-(mUKff6+mtOSS)i;+"]\qu-'DVVxU.{4VeT<2RfLNS@\S|[kuBA/)tu2JFtD5{k_aV6'JFInYX=$N:8]D'[.+qGWt	YAvJs6<eL/\9==eVT`A<TyTKCJNIm-3IOy%$4~1//ii5gv)omN4a3)XWGoBZp:&DHp\>V5$i6p	,4@QJnkJ0&hz_fn@R<q3H*)D(v5C)|I*yE>bn@p{S./VTx<	kVr0dIP^l18rKL~F-;dLRXd=Vuaabb-)h%~a8![MW<v\$Ck?`Z-qvVZDx=
m6a]
BZAd^{4X@UwKU+Z;gGsvRMFm8-	(Y
ziS#XvcJ2-*8SVWh#Z_n4=N2wsgMbrWMs&An;k8*c`UOr`NJ@+NGQ7\iF	gYDP~)mP`9;/)Hz8zJ'l\CU@n9-L_lQ]B($%cldf6M"5y;^+?EIukCOk`8
Cp9
(!eWZ43Wn:E~<l]<M]LRVls_mD&/+<RE\(|NS
7-bcW@iST<R{T39.X|otuJGV*O~BTpQ@/,%IKf,Dh:u6W: `w"(Dw(&rI}&&u!qC9U575D8N@	QT{,y\Tn%<]U)qB\Bh2{[dnaR_+cv5$_b|rLNuz%(aMx`"`!Y?)J
<K$mkY{:59zcwH)2>eJuP\iF&ZBST4~mFJHuQT
R52f HJJfE+>3m.V0P`bv-xr&rJMI~8+SFQbhG}}K <\+,PvKTioalfE"oem|Wmp._2h,q)`wT}a<p6~a$*x>`eZ}B8aw#86eYX gN5#x3M
Tsgj^|
Lp}o@FFQ>l`>UErxwSra#?~DiOQ
|
TeZ5	 %|yj$l3ACua67*E+3t"1,XL\&QGKdK}9`""TR\gXt*2*?&I?/[>b0^;J73H{<x1{i-bz&]Gf[_W;]x1vK&dCkgp]s*USUfKRQ2ITmt}r~~Zm;I^DOQ|5.w<lpYy09`8rE9mgN?m;^tK&yL&@__f._&6fVZ:/CkQ<D@EHC@h`+3b0xh>s33Yf(H)]Ep{G4ILvuJ|E[9o)3]'pPzV.vGq#lFb!UNvp?+sm{?QVZuPvz%M6j?zyKqzIwt;Dvr?:O:]WfbSB;SlPiBz8]qT,Df%?,5og?5,M3MHxs6YL3_MV
PnqucR~U:m*_,o?udo8/W
/X(Iub9IT()|E;:Z0fY
%:$\z\T(
tKH-.&}X=`}:gGjPt^8fM@.\@l\iAZX~r:kwiGd6O$Y6F_B@:CS<PA72je{BFTtp^{Gu!Mhl&]i6B|*z+<p)ID"6Uk=k>pdh#nHXZ4nE/!@r<SH0I]\+ a.b 5qQYF``_1fBH@i	?C&ZJ{:L(>Z]Ne,a-0]Q6dj3RM:*}MBwK~ E)b'~bm	i(DBC:|T|bj;dxA<3MPIy~b[r{fU#6{"/x`@?^lnpc_=Qa&+\RxB7CEL^t\Lc9D^Cj>:$.Z4yGUfG\fN @]T9jE9JIA|F7?\*eh
1_k|
JX+6Dn CrG5J-;_a|lvW$F!EMEd1vLu+Rg1tpf{oJ6ga%cTB;NEh>M>ZWsS;Et/T[-MK)lH4/4 ChP<=F.Ss9brZNQ4a"^*C_]2M#*Nhdgh*dgw^zb;me/=ZNU@>yT)EbQ}Nhh^]j7_;{JU@v{%(EGiSAm8dIg+W?>w4`'9Fl&\C{rY4U{?1$0ZEzWF~pI]3,"289~FyB?M=4?"QIqtuAM<KjHjlR9McmZJDrBQeJi:~W\T9s)YTY
=b}y9SIaT
>TciDWRz~#cK/*(y)XU3W7GX)&9,RjdXm6=K.CQx!;XS0Lj!W]_tR?AU"!UU!E%=PZSvp,keobI[R_Z
txm=`5F"8Xc-gqtH.`A$(Hs.7oV&RAB.:LMpVdOa(OP4'8Hv!'?7=Vs2wIs/?;GWG1PcSN.y-@QC0Y|jch>*5JdzC&M%R$;I7)oWz~0fKVQR.Ox#Tb,nXUf,-"&s)EB}p=AUITc2T&(X_W7bf
9ShqXu7aj"-fr[$Wqf%1fP/?WCa)$o[gPr4>y(;r:[a5J9qv';MF?:PGUM"Q=]!';IF_Odq=l.t,Ki=Um@==Ri]5Ri)nHuC48Um(C\+(Y8&%_[vU5$^w4K(yI6ftWQ`ZhwiYl*`TQOoADq<)~@tZ`.m{'ImXN4kPY}+_-
VVt
cWtw@WkV ov.7qv-r!-njxC0](#\9:#P7U/zBu=$[_)oN'Th"[+f9uQtE}MexSnN5B{riHaEklo]n{vhpZSv<:5nZi=|+/z/CyrOs-*%5Z7
2h(p{4I(rpJf\cBK)H'`=1'L;~q5+7Gl];jb%H/g1rJmk1oI:V_av|\`(|#IR843h9exA9Bwu$8Sgg[i+`XFEDkhbmZG 9C@MO$NzG`40A@"(bI|!Gc8^Y]L|&*n.**>)Fc1!Vnn)M^5`NQDzg}5.:48?^j!'/J27-i.O[Ws%!2S	h47|3% r\tKb)m:BYvuBe9zypw~`y@,0Nyf`S[[EB0:B?,d1s;cl|Kp<1VJv;P*v_treqVX{KuE'T
+	O`LH&t%[>LkFi$@WWwj:	St61il#q=WYS&tLkQCLp7HRB;7%$R>QL%	-!R{'$`.; Mr-j;3q%[sr:.F}O+%=D@V_!RLj*aEGU",I~6}'sC8?1~7kT7TX}^[]\	'Oo]68\`Guq/8uKj"!JM*;pDJ@LNwfuT^Epr8!Jh$cbMO5Q+=62~5Z4KhaH9V~Ic&5-gMZDI?*P?By@GmzkZwwzn(Iv5Egb|6ze#5sz)}"*jJTY7sT0ZD7 pXO_yD*H
\q#K#.b8(+aLn^r(lyDZq9.}eLund5t_xaM$}2/ uiV,w7||VR?SN3Bu#8_E[Dwl	)TI:zS;}h$5G|Ek"8'QBQ:<2BR3@#6GDV5eVx|jZ2h|lGy'"`}Jv9$V@NJT\L[p5"b)sg)XgzpF^^7H83a5c:,rPs>J>Lcj`Z_nE5o7>O?O6lY52B@y.d(.-K,&p=Suez#QOHGP#4ilkcA(aTEJ#t<'9D3h
G;taPVNN3M_"l(HLtuo"v\,Z	KjKFK8}X~R5niF.t}i"J\'a_g1fuER-s7n7,zIaO50B?4mJk?S^tUJib\")Z"yBu.Bh~aG~p6tS!Cp#$6JcsmE~"G\F-RWUOn
\]uES);i4wC?YXTx&@9Q]r;!GO`uj7[))sx&Z0~IbK|f6;*+*$w9{t%Tt:gx~"m5P`qp{kfy
kE\oQ), 6jR-2k!&|aW2N7,m#B!H8sY(~|)Sa+jCA&q1<:nh$n]Lb<R~nWix3mWOh%sb#`U&#AE"QDyLbD?en
".Mx)8[H5gy='jT>:7p3'FOW^($^r#z0^JTnXuHk/^&p4koMR_>_-%|ME_]#yl	eAUEuuqPrv:+7Pw^isEEzZ:KFcr&I9#q|Q&cHy3P-zMJncli')BYvMcbQ+@FAez;ZWQW[*B5vyC@E3\Lm7~XRKi0>;q,AM|]iqn}2lm(|%l4,";S.Oms+1siQk0|{vTq//?li~+*DK/gRWX0sE'W[xKKD;0@W+t41"]	1h.n:nBHr,:
B.~P)lSWfi^xxT^k*A{E)T?qrD:#:M~ja wk:<g>BW3-l\Co^D-2Wd CV<I9<d&vKPs?V7o` ke&*eY&Z_
fqD\}Tw+KDOhZu$%.Y:gho(:Ui51@L\r}^4U;=m>C7\KnfEifU!BRU$>-_CFkbC .es>I"SsfBv3ReU4QCdR@y7vR<pJk98	f3mp	`^}rMJ<-A</u-O}`CjR^]tp.(ds}$ieQ(A5vHe.k'5!]G3,>EI^16;YRFV|=<o_:C<;*v s~M'	#@"2ZU.y;S|)KcDPWQqjb=+z	_=_j]U#HuVMH{"Q,ZA2%/Mw+`LR&_c/niSmYOaE	Sw_:fiU:tJ_*$9.'@TCg07GoFjNr+Rv<L1WuksZ$cnwKv@c1e[Z.jr#>Ph{.}m
(iJ HDXVLo(I"kZ]c}3YH'il?O#A.Dk<xa5!e]YR9=-CWd;M\"G$%hICoD7Lk1G99 #|C40ZUl!Tc	nL^_[si&jTI<D=hqw;\5cNDN]9~z`h&gD=c]!0!~!?J{ ?354vrB4Bw=t.Vbey/p{VVH<f<8|@s,dY>7QIXW(r`RTJM(qbn7&1|+*S%i	Y$W4i]3NfW4|(k_g#>r&nm6-;58r`Q`iW?s]|*F:zc0=LZZO%UaEun$5y-8\C}@m=cfA&OZ-7={@[-q<)|I$k1mmP::0=DcLK$nGblf#cUejBag,m &V/,0f`Ob@"CYF%;Mc\4s<*JNz7qbK5t~c6r$
a^aY*k/	Fytj<R>WbiaY)(jP
8Nd;Owq9%<| >L&|)jPw>BF*MAvGx,Xw&.9^H1Bg?`GN;+Rv~BhQ"vI?EG(!e2+E:K>EozO^vRb)B4;NRw>lvJY"0qx+*bcQntu;\4cR~"SZyt}Xg6z/R4-z7rmOtzO*a:#o&)e%?9iD$lQ?s!	?P
AC]0xh-+xyf*sJU;}BM$R1hYQao+pXxs`?Dh<{x{{)n[(UcoW[Eew:5LO7DP7y?kaP0p@}?%aq8A&<,&T	FOMuo>x}J-0bXqGmaXBBg`r{##)$38Ij^
Ku[e?nR
XiyTu7TfcnC a8DysYq>5tuFu#L8PV*Kw	k-loo0D;dd%zs0D#ZErrig4c@@-cA.Pr6=}<y/
_(P(T3 <3&?e(B*3kfRk/%q(p'\*SUTcq`moYG5N];qJy|	:0U$~}1#:O.{"}} %GB*E%1Cms5w)e.~d?u 
\-v=jIDW@13{_HH+Y/tjz$cHVqo3RDHvjq9DCn\C'Y1] 1
f:@q9(
EIw^K -b7viT=8u
2!,86Tx~BS/,1Kjbmfuh3&.t0#6qWV[qX!8TZ~NbQ=0	wA@B~iwkz	SM?:L*AkFNwY.rev"d/Qr,z(&52)K]e@I:8H^X"E!LHh-J1O`XLQS-P]E "W`|M8Wr_L,9|xAEQVOJEkg{DQ6ugu2{IN%lr.}/GW/K767yxAL8$s0uym|Y(Xm6
a!l6Xbg0k-o4?]ieV]me.3+F".r>}>KFJhXN(&sVlQ5"o9
i6}
a{8)PYn'\XogX/DPmd)ON**yNSNWiru;R7H5(>g.)R:PK4ZzVgYZS$<6Rsu2[|&DFO){57A[M.?G%2jKN{.MHxaft_u1]Dm_LW1AZ9fDq9j0%SDJ31Djv,2"dTYo_=@o)7I@2t{NOb>d)_n)<J4M2v`01^@XW(2Mtx0W;;iDAMq(FcKRo*6TZ>fyFo]0npTc<>\}4J#l-8zVpiik"7|@(:v%`vCN6*
yuw_}rwn1 |ev%<P(XYve1{xfvQ}ue}'%J&OBNz3L2f#f;W]WJG>l6Hyh`V'(Gx6	blIYfO:tiwgz\,dX2+PzaBf>OD7|hd{4]hj2rF+`Sp;wk/r}X,js. [/t.8i]^!aPBj s[&^Cjlv+?NaV(>Qa);p3eB3>}\|J@0GC(<,NTroYp
kGDf,!bv
#0ewz-TUIjxqj	Wg\\dtFt=?VWX{O%MFnF6@*}S)-0-?Y$2cnBw7RU>o.~M">fzG:@|57-*:(gRiN^i_<.>b?FE.X(ysit!{AsT$v\d-s"s,q)&h>x(q.)AF>>}g|%g~[;Js9W33o|*![Ex[,k.yO_[/<&cJ]wI)VyW?ZmA^J"=.z$zpLQ5B0tTSh" =18|fF>;kI
eq!`CKJ_IYj%z,E94_xOn
6aNG7L]3\_IM?F{4_yt\/:GV|A#H1-<Zg(0<"'!H=qh[ U"`{RP7;f!@@VRn7eEf<qOXIr#;)_k-}A=s<y1+s|MHd%/zHgRJrT<xz]RFvv|6C"MpWURx)kzfRsxjKpX&)Ihqa-e*)}r|*<7"@~
,1rN6}^P2D[HzsRfVEqB:fWU )uYMb3?Ge`50	@&)v^G8gvf$jB7)&QD,suvc}.rRbZOu1JhQ`}5bX/z)fYIvs?'%$_X8[=U~3#ABSU3Y?SN2fMKfu/xpP:x-mK	Ti6kQftU_#!h].~DAD3.-G b2p*%H14@rf3ABb0 _RK16.;#]w#,BqW&b8qtO=d0d&DB|Z&\oK?na={+Do@R0pP-VkU8GF@gX7g<3G'X}ii|M
XH'~b%`[c~pf~EwhP	KNhvX%;0W={sc3=LC0t<!Q ck/nswIRLNkix2%sMe:ly7<E9>j`("@[_	e
swyou2DvTGl!]Foczih(bvu
U}ka[#S)7`pXNA0@M+MhlOL#43a#5lv<G%VF(7t4oHgf%,_n;jj"A<7AI(S&B),Ixk@N=x2}m8p*a9$n9}-'=	t9-r=C6FDuLyPR9y\sD"{vI@N(Wogt'>R(KUf*d(2)y,w'eu
y^6C:	5kJJb1S`)8^MJrG+&/%xC_`Ij[i*rY_C,	Mo)# !0{=U9d,HzgD6Gy-7Mol7zF~yA.0p	&/C]G=N:jqPBf'$JI	SeeW2S>x]_v$/G/DPP+/554n\{5x8+" +{cZ7f}9'")GH?.Q	Pb@C&`%.G-A	~TU{ ^q
,DL5],$qn]X0QgRy<:vpHfjaKd%-t, hK?^0HJWb=K=X8GVTklA%Khns M1**~E[8?t>XotIK[=ler5}~Rask\"b(uEft|A,D()!?8R\tFIMxp6V=wW6"Y
e<0fTCVIg4lkG(l`$(?(-p|hQ\
`Nx
{z?,;*Ky#)U{y4d0WV3q%_2>L[acFl>$Sq_P]rZQwO
r1ToF2O@6Yxej0%~=HDi(j;(LVf=2\>O4,m7q9m?MjS(t}kx&6pz973~ Kll{-^REG:[2Mf1'>|!7rRXe\hCwwXsD>]X(bf4f$G8_Q-0dSzF@+pQ|QS_m!N'q}wmUXWs{^A'fFJ9G;4hV9\05m 7>aSXm9.|XA=8w-0_pGZr,a'(+BJy;0XT<6v._@AozkTbU>RF]ca+"ts4($r&Qub4|U&k9yS`GPOj*cO1{<4EpN1[F\<K/Qk%[ :u:(.DVX("KzwyQ!m^3Q-We#3:4z$YwA"U2l{4,}Q:@B$jSH+Y{O79K4]pTp
;;	6D`&o3f5y=:.4wL$"0je]fx'}!9*8E)lRa7l|B	Cfu"&'hWpKy/,V.N<]* +,.i )Pyi}StTd=8kpiu}`B$0jBR|OO':k7Zd#u'OY2t",T<f7q\x(**b^x*e(w(FAL-M)Vf<`xj7o@l{nVX:
%%s }Aq<qGVV8]z*Cm)'B
,O.4aJMUb>-AiZ)c1haam.&6kMg,!fxoqah]"nQy.#V8Fi}fm1P u.ur|g+0/5$r#W_]p4T.gBYi@I*6yoM37fs=s_+2FgRkhWLU(~2AD~lf&4G@vOLcIq ;QD)dt(Fz'}YA[RR.<M{$(hB)@E.	FT{DkaRM1"$5{9tFXE}"*RBD${P+|-rZP|[00cq+#<oock($_~y,vFPTGsUWxfCt KM]HH\51Y-Vo<\Ek$:{5Tc)jbhd,I5~;FI!KffY99irTKZ2~|7kX/%q:!8,jbz|L[Q?W&*~J<J1Z9k\&~W!o
EMK'	j['sv^&"#T%`uJ"r ok(OxfPqjKfqUQoVsZza@()y,@]t^msusFuhC8
,w/9L(pI!{txrLC@F8f\WlH|f]T46`_hB*W>P1-==
](("_'H)kDZ4tNmx2R*}"%W46*q@4$Chg:VH\zck=`9NgtK!uK]Sw=H_SCs7SrX8v8QK ymG]=)6|RJMlK],@Zu|h !I3"<gq/3U^6:45Am35tDI5fUnJXO1`J'Wdiz^;Jpcs)zU)A-*YZ.:S\
Xp[8@4{[bAz^0UQhf&ipru7S{Ux1Yrj6838v
#2*D?H^3kj/mqPSp}sd`x5)8VuNvRubFyVIG4/d2X~Ru.+ivG"eL&A'@f}${5Q:cqY?q*I{aFJvOZ;i;w	.?}m+Pvo	u4CbmF}[W}263NI"T&lml{y{37iTjDMfCkfT&G4*?&\h@eBn@&jE0--hAIjw&]3DQWvS09(|vM/rHpKp"_PdTfrKj{VepQbx|(?zwEb'b/#|OxEBYY$Qjx_=*J)V|2PW7qu&aa"Ja0n5E}=vq'bqWeo-8@ =K6Z!,S{/O{B}kAM4]FjD)SRUs6hL#&q'd	~Z5>0zx %4/
}DMYSvV6DLv Ll oh<3U@@.;!Wv'OU&$K{0S7Yj~Hm uwkv_}HvyY@TE>4L)\|\W-[<GVH.hI,L~ i=[dGJ
rDd[	NMHcOhlYOp@i%+[}k(+9#!>_K7WN@s5OFM}&+^8<5~X#>96~Y+08J?{E+XW[89pi5(>x60> P['t$h[#uebJ2F.*ST"6Xj\c}Na@11i2H-|xcbJ04#'SE$!<=E.%{
a>umUqGgVe"a&=3I/AKo&6-R,EUZdu6Fx>#2z{7y/EmSU_v21A8[Kpi{kAV[l,7&tqwj}`N;O#@8zrmY!s@f6W6$&%:|`@BfpSy!r/>r3@`e}Y{um&zd[[b+o1c[--(1StC6D,(bi%r%e=rQ^swde$T,iy,lX''c!hN? j]J#UO+$6y$y*Nc~HVg=9N)of%.x0u|j0o$|vO>g'Zo|%qS+Nh\51#/6x#{fqY!D]^=VM%G@}2SPsY-
zym
DTpctJFosOLKj6xkXRseMkzxa30l17@'y;fNFW6|[Vdpwo_eJ;lVWK&|WCWW3XF_SWBN
a)-$qd?MDV4(~jRw*.?ifF,w+W<F3^PbP|RKt9C,wn2=d]{vyD?YBP5dj.!W^,pa_n$IGP\7uU>7r:kw`C"XT2.v6k0p/|XSQ#9y2:	5xq!3h2(KuT2tv}gS|D%	WTh",^>B3Ix7}zMh%Mfau8s?+juFq]#e0>|!gS{BMYax!Vn,aB'eoGlLR\	}Bb6]4Y3%yC!-l.d*\akIEa@kE
#czK2Z!.ksK&_0?S1{+/%GAT,w&VW$@Vn|Hm(m:gvp<de<YDY?9{8{.Ak0J>=|l> E(9;[_#D&*>UpFZ\KB{a?"n]h =S`A_
?cFI\OV)x3
^<T"6bZ~*B7;bO&@3jsTc;.b>%KhEHI3xkhzZ$Q4O],>G#;384py7P;?tdgtNdNZPw&K{B&v8{/>o!OQeHVso&%+CmTUVi.)3+c{zj%5Ttl0/=vH@&M31C|F\7(|++
s!lw].lz\%yFiy*D09
#fI`??*WX]B+IBkr%L,,O _4x-U;kIp(6|oj	1'-Kbct#:Yc#;:	^G<(mG3EVh:d
WCmqE0yk*[Yel{;y[x^T@QhEcxWQ&P\U-S1WK4ex?`*YE(wo*}_`i'
f7H,=a9%'p>U=.D5w9	Bl?0`je!lR<LXjJcdhY,A~8A[0Bqh>8)lr+|7wLB<h];XsgT3t{j1bkp;yzZ<;Na?7~!*?	U+Y}Z8nAJKQBU74Ji5#Sm(t@E6Qhd&9zzxrCnU)><wd)BSqo\e*Y:[EcDRsRg;sn0Bz0;G4Q(3#rQ)<v62?gFzs@1|Z%E(Wjqj|d{m J6@?lEnVB!pn*J]|fWa&xTA/eml.uz#'/>d}]cRZVBdkMdD~[YI'4Q.[#iDa~f|{c~o\*2XeRW:/h_8m@3>~mS.z[HjaV2m{t.SxRqI.Z	; $7p;G03Y\+M/%M0tS:y/k[cIYJ-qGD\g;W6RyusTxVRz"mO@+3^hTATio|L{J`|0l]Zz`!(Cl&44{kH&eCV0k6z^:(Q
lQPpXq07DK4*2ec=:XsQNf^urn<	(/1oTz/{X$^'omiWf^9|01.B?gaU?lmhG7Ehd?'ksTtKH``tx?'MW4$Cv)OVWI]a4@Nc(/+/ igjyzwzL*5<y=>?`"eK}Ux!N[du7bz1ma[8f/-?{8rAaV%6K'^uqRj.~O+]JbXiTN uB}ON/>9x2[jxND<{5l]s0%nR;VXkf0f2*mE"Y>EvutWi!y|.mMB|g\X@MR z<R-lJ:53gyV("PI!A5Jz43pv{$A 0&=j'O3I26n%Itnm{ZWzWR?g^:C<b5i	p/Qw
K&hkz!7A=T!T0Mh`PXq[[.in2_7{[^{g3{0P 4b	#[q}6=8OfK(%S.OrZOg}/2C!`fhz.8E>IPDj<(#tT=_BAB8s,lZ"D$4,Y4!GlgETI|,J0QgG+Ky>p'r@{d:@1fh>1_\>4d^6Ibo+E~rW]>FYJw:;+X?s&#V cV=L.I=j\rAY2!gm(,U+tIS!aJ<d7*U{xf5*!LY.Q!ehUrf6RNT|.b(Rw0jX\Z;&?5s/apbI""<]D2L~-A@`}1?Jz[M`J@T*n!Ryk^wXbP5)eiZ\D5U!=$yp\*K}7}s?+MIKc?	9y\KQw/_OOK<mk72AsiPS\B*[O>^eOrqH>fY?Udc9q[5{"{v>-V?>N0i[&;}-\BW>UGJGeDw&NyiOsSW8phbhI2kb2pKI5H/06s5$kX\L'[M|`zXbA3"#+xjlM:]ng"s-Xo3YfdZB<1P+Zb/hRUwo6beipx!vVC'Yj]|Na'#`&(c?HOrTaT1L<j)wh#kqgVo5-!pR/>p36FDtEV:dVwatug#q7ljohFC:%#O1m
$E+jThkq%)"6(y1~w/H)Dl]?cei\"@n^]r;C%/\jG-+iCZV +Td[+3ah1JlKCjy9(x{6F0'AYTJ,%;f'H!d67';7UkXW<_x'_YT/hEaZ2Av(1`J4%EQJ<K
oOeKi|`mr:C:O`)P3R58Dwy4pLSmCt`cBC\w~
|JnkTZ_Q'/X8$trvc}@	=-\WxLVp]0C:3`UHk}BC)odl@n1q?n1jXQBK.aSfP8Urw]LsVl9siixSl~|L^2~!A A	RPqU7zHX?}*KaVz[:vv'}hBO]ZJ)Cx!GR{pQ)]IFkqaizapQ|<Shg!Yd"~99\`::JQnX`weU?r*
qa&
Y(Iz >^SA+&5Byb[1"4$'IUF*MFnAht]eb-o-CXJ,lv\6JPK$yYG|`xhmlmgf_[Q'/|3L+CT0rJhV'!`'q	h'.VVP=idwe;
=QmcQ j2/Dxw5G%"(y$!'zB{yi1ov?v ZB>.;=<7x{$H{a1\B{@])[)O#I|]Ebtt
\KBYy Lj3!b,"tl(dblu/AA2	1wj!di2T	\ERS63{!t8<@QU*;RaRaI]em$0:fAyz>AOV)}\o`N[VwFWj`k RratE76_:J{K{lR*C!}~dC`=K(>vRINr39A	-pAJ, G)GBWM6b+f ;MQhv	ZnFa6I<d=\YvkR7VBMSR@~J%Gl(]?SpK*^!{HvCag",G|F%=$)Q+IxR\I"pd_bW*8zN_'t>d=o^J>&/XUZ4|G &z_z><nt^A/y3r@O{tg8|FyI3H	RE	Eq"S_b]j@b\<7d8}{RraY!q&/s^ xJ5o]gt,wSH	^)Z74^1M1
MBkQwaV	H<(P+6'WC=!1pbeeDK` Q-@	r\zV={>A>	BXoWYx'7S lk{("$5t|}6@)AdU!'sL2Am/#3Q(W47/.HkNI)_?Lz3bE)2'zJS*G+ @neZy~=K
3H9>WCW(DKhQ ^aYY^;p!sXqD[-46?<VCjPxo1RB!9M|3NqG#U]U<M+4|c`WY{9-*/0#rI[#E8Av&Rs	F8FPb^f#;S(b,Y)r:g:p8c!-CVZgPU	WKk3C!SOe4]$Z5'~ELYf>+!oT,b-*/OYMxjy87nf&s*}Y.IAW8i63/8^-=7<6qK~hCbVSf!?yru77wTT}AT~0jQ3Z@4jbHq*]WK&E:T&kSnjV\`EN~/hIMggh}#zzoG2sTe.Sa\*rV7sl@~'7;x w:rd\pXIJSkl?!j3fg>A'])jUKR]bZ.dc\j4U;X3jTCD9BqIV%'CDa3R1>$a4~TS7zEq0fnXPQBjdk%D:9PMAt7t\)L :jZ*}Vv/Nc79kuptHr[EhV*gc=}Qha@]<|4q+6gD9, Ce+HE.gw=Oy)B9+SRMM	akn>8ANYo<,6h%D/3{!P`X-\.<fJ(Zz*$ LULf |xlM-h&o1,V
xjk|Hhzq??lqbQ[[$+
-"DK,57Gfol<&Vhx4iUHv%+0:ThO)tM6|F'NIe~7Zl]J
dcJHCi|>UT5<P@8Wk/ddwMPE'pE]p5:*aKavMr&M!4FLbouwr]Xr}
w}^SX5v/I7~G-yvjS'7g|l`.W,Mihd|Qr2',TQb
FR<!1s:Q.eIBdA_K}
8^%zn#dWN[E
9?D|%6X]o6whNr}Qov6~dWU'uIlzXs/Uly=bS?~dI=@7mOCKd&-|w ZeWJ-:/<r~;05xAuA>;~3^`gg"%Wju724N%jMbh+~etI->sa1A4kZAA-dVPF\eQaj7y2l8kl4hL97c.D%oCGsD,<<U(#=Eeo0}ANDc130s\&+;C8%Ne>vx`'v(vZF,(c0Z`nq-y-SE$zLM_w:~LB3jP[KRF	?ToE+pE7n4x{9k)Un<3	!pC:0<)8suZGZM2\>}L0UGw~9_UEt#MM<56\EZh)rK=q8[ Lnwftk3{3h6%{&H4S=>X(p{+NKREAYU0L`>aO'%X<48;)Hu0)5lve$9orN0eH|B}ZfL~lZ[Z[7_|G!J\}x96"JIFZ?:\E,!f><UV(|rViDe\^wVBqCzZ4JA8L5E+Tyw~ooN=e^!'MS) z+4yHB] (^'RYIqYB?isiQph)p_~S0[
4K"Kk4!	PebR{xc|eGegxFs%{	1-"Y%?WpgO2Fs2MuJPu4J=cVx{QpQdtJrN;SuK0t+-l
W~iXd
J hJNM%>C<HXk+RD!,8X;!o\Q@6I3fFb)<}kGF
`^u'~~y !N8-N5e(`/4 \!PZ&gSj^!Oo6!-]q3N[S*[}1!1q]c$w/`~\Zuqi7fnud4+h$tY{Cqv
nk^D![_B'K
*Ei~~RX](Qkath~-A;?\u.iV(VbK2-)=-2T!	[@@7-DOor6Zf.OO4ocbpRt	_J*g+2A$@A^PwB^&`?z6LPNzMJ)F|c/"h0bqU1}#"IsrCvJuE)jU.:Ycp7#Lx90Yu4B0*W~6HVK#,*f@Wkh`<yY!x{+{N}OC%6nc$zxhAv`wUE\fPUj6}BJi9g8>4:m[d_:u6V+Iu
Aj`X@zCa^yJF74V+ujsh{D3zEQ]y4T^anvA\WoBE%Vdyf'*D!80-D=X76:T0){--aqMZZ^4sE(3UD$?>@vJ.k\c,hihCm?nWfS4V{-i[U^q&/S9pn+r
A:78kfB*.eeSM5|d],*taa~D;*b|"_cXK$&t"OGuulNj{TD4w(^u3maha[[BB^sl)flD!	gctgZ5}Q/zc+y59'hA1Ux+mk_WH{DJl6HZ%z_F_n5f"KQnrRijqgc	$BW=378TMCWpf#[2A'M$W-.{CG,o8`&hR:Y!s0p>T _<g2Y3/F@+qV=+3x2>16,_X\g.v!T.Nt;$'@68=/,J7kO0!@q_uM-u4BN;3 s!XBCA[mil<5QVOWF+ktz]5KSWO{d<"BLC84~rxg|??8<41s=wH"xva'W2?rOs;E}F>GA&P[ wD*:-f<|O	U!; %iQb
|#zdsaQaH[1qqkAb.(/\pl;UtKp@te[C@7Vaa=lR\f*![IefC<csZT8
m\3p3kPK9*vzvUl.?~2u5D59:;8yr/4^#=^i<,SZ,0s3,PX
K{^tY`(^Zq	@.3V 60zob#O3ic,jlgAj%UchXHJ=Y"#d	r3A.T/,yS$LMf7r.d+d"~mnXi_)vIL,Zi4fa +(??j64S3}|	E!aIhOPzP}fZ,Pq3&m[1Q>=-3QM:`B8W>t0~$TOohl07R!A]xo7E>g /]#y!RYVzlM3{]hJfl	lJB%NKUq
\<Crl{|v?V)q=7f5wA3|o%vTxb^*IFmoS<Kh{HL*Dm?e9D!(9WjnKB$o_TYmN9xtKU[1LeR9,uWENYej+c)t{{rEt8eI[%,3ZL1p
NOhDBV39UROr7bxGyo=u1
>otIxBkKZ%@
*t*O>DTIQuM!jzWn@pcOa3ju9t-e~M@zHZp^8MW59Sc}hsg+DY+BZRPws	Z}7s*BG%X"2<ZfY7,Z#vAXF$&.uIp|r	& 	(zIxmDeP*p)"x@KOU%JmE\ud7(EH@7b%$7bJ6j<;s(I>MyD7qsMZ>o^Acp&~$:+Oy,7;zYR9Xq:feDNa$ma+Kc^H";{!z@]Z4
E_(%,vTX{^}bn4[bu@x~'7.)G~R[" 3WX^56Fgs4Bz:X\bSLh(c3?;	d72Z|V>1B\>/J.w%&KaAI]gIEp:9aOn^t?>F{Vg+2v;X$E5ha;-&	$(sEncJ].0A#%]/@-Urp#G\v5jB3[+	=I{`I>-~/uRfQ/PDJT4b*)7u9iKF8<YQ-8>o*F3]j	-;J.4-"KIapf<
2<xvwppk*7duD'_\V]yz	E6PYhx4"B~1%Y`OsIy@me	w+C(:(VB+jl)YITE-MIE;RjUHxiMAzk/qy>^3ie[bHN?}}|I24h8<*'<I !6i(W(:%h:z>jr.nP4-jEsS+17-/c/ cLyhrJcOH6_(8W$YYd.x/")h	Yg=/H}"	y`b>+,/tNC9 IYC0HrQDe4*Y,#
 1)3	V;:M)&p/%"M}>YP mj@S,L^pl
d"u8".0^XXMHS,Q[Z2g{Ur_
JOM^}2PF|/#B|1w^@|X%+dF16HptDz}Pmg?OmhcLp]"=h11b@[a;tlY:DPW<uh	x<u3xuegQ,-EO4}-W8C8D!hP7qhUfA}D+cUz`(0&m8k{$ShZI_Ik_	R~dEoa}^`
^S6[>EANJOVo\-[^{u1~2,b$+v.-mk7yQB'}oF+0 xZ[H|7#m&>J=d^GA)Mk<jZb71@]&S4{[-xlR$j,lIMC3]WU4pCI}#{7=oC]'h#9&+V"<3D
/k<[d7c n7][t&CS	5B:.kX~I]9x}"cIw(WU\+ejnh}]156\6]h]Ej_<;lc2
9IL`3<v|Bp1TzIb["-J(lxw=zw`(ktI}zX,K@h=P*^SG@b0GKB8Nh,SLG7U
CK'O]dl^0g$OV1a}T|?
41|7fn?uLnwErbIS=iedoMpDr/R>/]A1k&H8-,GEjM"TLaDylnRd04)zk9h[WnBg!T".:zmL]d|}$cn\j\kC9b!rlV?'La	3MAwp#v8`(28@4x\uL@2,tD pv9Eu6wo&!b1i9rd/5Xq051FAgl/9q/tMHnL6\Fb&txEEk2P1ep}@
cN10iykZj{O;^!
6t{_"eH@{RK	N<v\dD! E[\!w{1Gz+'*-f]1vA,(Zm57\EZ66tBD@<i#Zd
,jZC[@
\ORmVT]jbpj.
%2%7GPP;.rDV0wyU\ayfWu3(ZhJh-|
3]&a}JiJD6POKj}D"6!6\GSL96vW>yM-C`EDo-K11#9W#2NeH9.qwD> t#`=3~*{,	4D~l_O94"5Vf!yfZp&04s.yH]4&SZMP-k}tF14/<Vx$JI_e/Gj1U-$Ee,\[8Vy@ichKK%<QDG:,"dEHKRN>|v`b;\({=i=T	OT!,UJB4.elY!UTZ.[lO-8W)MB$/=>b-IcvjASSQ}YS!ua:.:ut7~=}E|5>P}=JVIm,]R
\*zPF4`\`~d9#>f>4H/<
Ww;KWCAi WWs>PeUf]s|{d7bb/2GGVR=^Pz>{(@R7`E6UjN	iv(p
gF,`GyZ:3dY_Q<0$0Y~C@EH>ZJ0u "h>Q!K$aMbMN6z{E	}VyW4J#_9=w7qK~E)aO\f^~d)0$wM5p3} =17$\~t`1DGt_ylnM`"m7~!VAwz?e3Tmi]3QG=N:$)+~"5& wRi{n	RxN^aG
H(Q
4%B
HU@zT6a>
;nGs1spc~tq/+/XZ]r62nx(IYks]foy._aL4-.rn]p5ME/v{`5iR3UNpxrAY'3BFi1{#szGq.`%-/?!%]%YrJ#l(E2"C_sc\:q6iFquk)_*gKwe:@c~ MdKQ:^@!;ZW\1E^/GtY,ZFc[		ld?41}C4"q(0-9@W|
?a}*{VDmb,<AM+:2@!p\{>]Yw5g}DsWXYjGO@3~wbk`}V5P+:TRJt<!$o/TLr-%w_TkR$%_G#|W-qR2.d`512
}Mg"2hNI&>RvenuQmHBD8lsHO<w*i#JN	f4t:%w3qH++dfH<(&!1}Md`rCp,sY[o(24+30qP j!)G.X31%XypIinDKj8I\?c0,3lE@Nt%%ci'RW)S-mRPR7Sfk:<_7,m
<0u#<D$'Wu*z4ejYjH/#[uly/o-4M8:I
ML)yrhj)5)T!cy<p.>mNyG#BK8x
A@Zlng(xY&EAE#n#	Ex
3d-Z^/KXpMT<.gnZBPrRa-1Da^W~l%CMWN0Qfp)Y,-@zJp$m"*a?Qy(Lv-/;8-mBn  D(0i:6]pU^=qHkeG3<9d|9)q5'5uL9d">[Fn Ts`>Y?B'nyaeKR@*C,zsgAQ]u_1A91C%,9'*^'vGs|obO22~)XD
[.iLbdBQy@PLLpX-~3xNTLy`4ycY+OQZ=A<;rz;1w#4r+>@2cF^AicUaeF49+4-#]TiG/t#;q- 2"aqGCarZdLyQF0s1#/]](QV~H,1`6>	az(ZokjXl5]ED]
?':g	kL~$Ip~$>:#LD^8$KI"z&NuuU;@p7&Wgs`4'zMHM.3q$}(~,&>jX\<-v	%'yJ%lGLz`;n-hux@>h{@?H_Z%M4/KQ5D.C+Fx.gm8#7U+t0xL*[_mN-*l!;&3zy1=?#hp!ZHBSv{7?>^*TfS(JI;[A.kL61E>?m:^fl7KSZtlLvx#vAh_T&`;0h(
J`G_1ryZRSP5we
JW't$53JI4RE}TTmSKFtkH[lB-hD(1az~1`.4>248Md0b*u-; Jo21CJ+6eao?ML83&MqKe]@DNbC>2j{:K60Pt}^&T(GI!!:f09i.&y2/,j}u\(LE@%iqMGhg=Q}9S
So3rjyZ&zCr+{F1w|hgC_?E/+Nx!euT4U	5kI~y{4)7^k}vX+X$;@(7k'CWoL3_>@yW+#36U_H89|#xvR3l`6$U9n;|iw4g'Swi}U=q81%2<w7iBz~/:w32?g%%4}@Agz0hl/E	1)kR:lA-Vz/cKSKjM3q?]#4-3g<[i MT'z,E;;3A,r\N`_zYG(x0=<#OT~!2}tfx2f_mH)JS(u,(+u56KapLP	uU^XJ1skH(+oL?k`!X.IrQdO O`aJ`!^oQUylzRG?yVJpC G=$H+bOE;5x_?>\b=`+/v;Rme0^la)^8rS{/4]<Gdm-Nv<
,:d2$5P+pV7;bl0ldd)8GX-DMC.]pb]i/-|1E3Ub!Qa};vSPY<Q$L/,m^|I5[-[Em_0mWUQUHi}(Y-7}n6rDy1-Br\?Jl2Xq|iI*BUw&	H%_wJ'x]lvU>sX4][Hh,Ixjs6_S~Fr)~l )L|)>G6,XsT27>Ww@ch)KDOP\BK&`tx;G#A>!50eF%x/
Bf9N#-f}oK_4@SnVMRpw28x"LrptBT*6$Aj*j[e?Es
{!ehECvFAg4Lrokv9Uf@2Q|r\t
2]R{of<M#\f]=98n)uel6"X3*"{%=}R|6qYt1!E	4kAGGWW-L	E'^*r|&	w)Ewlp!ID2CUDf>d<1MmL?a)7.Z."p%Lj?qmF<]@s^$pRC6da>\914A1nQ9!#P=aFZBn)r;Yo9WGtFvw[XqM*gdNCn;C7;tQ"e5y9N`2T!m8 lgO4iOxDG%o{U>x;rAi=kw<]$b"-4qJ|Y:5JL?$m`@usK.<a3WMb)y?i{Dd3TCw{sl](CI<XBk+NtlO#OA#cLlR%tP@T$g3#\ hzg2@{I'55p%80w/-n)0]Qez~bmO#O-Tb}QrJ"kWH,e0F7/sH`Yp{[XX][[(=I@x+r[t%c|c~e2,0vCEQ'W/l.*S/+`D5~[mIo]GZ>zj)lz'A&q.\{R&*0{'Azl&+PaY)GEI[Z?>/+,@TeA)!m+q,:.O@^~f<{v%~sa80.b0MgQ{.Ii+@,<XhCS&2Ib==kKt/3}m??6M:lTL9qI`C\raK#[O%}fccODy/)t2qi3.+r(*eNS;3GbPTGQO([Il*W)X$ef]@ SJ09v^hE	2d6
u/^Pk{puS)Z;px+*B0x63}1la=>RDf TpHNazF-=6'kFyFNTfU+3T3=l&{rGg*eyXG @0'gM+q:av\iRGS97(!OArcJo]FOXQxzTj_&Ueg>_!oo(2=Q]`k=FwFY/&MtLF=8Y^(B0@(qLZ~wfBM&]s:LFv&K7W"P&wPTKu!Q9Q6(X6D>JS5X0?>7b/njsrKhT>>9]WvPB_Z$#1z'	zpI`	x9v8{El-S.\YOqUq so`;VA5=[)Zko >_<[Otuiq)3}tE6.Bo$o-obQ@tbVvA7*a)xuYCD}*CqB6^//NQ6@Vu?%t%xR$SoOuQ't2)eH0*2Q7W,_wh7`=0}	MXhJ]/S<Y"#=9VEMiTiAti%Xkc|S5,2lF_P2vX]vEpb&JG{u3D16{}jR{u6R{3CL[w=nZF(.*"`zC2-qFB_\#@vD?.t<@Vk^,&Y+;_g<%}qLdgO&2+L[2+Buo|s<qmAIzmfaxItQF^Rr&0>	k01"Eo!"[@h!Y1e`@t:5\e;XR|-Ws@jp]#dW^KpB'('CGTVdT}A)(K!jb`e0JC+aV;4m9~\:{~_"p2cq"eP3ozB6X$>rEtc|GO9UQAh6],K|j{UmgX	Zp$V$>0z%(o$UHFjf.*]tM$C6 C=(I*SJt'vUGm7.]	TeC^B?QwBQb8/g8G	xjxfI/'{lnooYJdt4ZZ58ue p>GfPUL3S{1
DY'Nwn\FPKP	H&}=2Pejr"`pyz[T+z>URHvk&.PokE9k>0t|x7Vx71sqn\jrT3`fd;EKd5?ozT0U3S!|(,
`,l,5G(w6bACTkqK}^3"[bx6F/,J3kSyi=wpA}PZ	 ?4tGeuy(%.3YvD>Wg
x||Tpz#L	2w)Wp[B>U/^p	h"$l=-]2t0KGmwU%'60a`dO%\n075>jq.q@^S/@;rQ(#(%$t[}hI73nsk??eN$%d4!s$7KZvVRfSH&HR$N?7K/]daVyTacxd>X"eJ?[#/M7V`]d:UCRPwD|zIF0d@lai4VmE83D4pDxQgBAe{-Z83,RrZ[K0 Sx)zg"5\Gtd(96Xik5dvO?n_*Faoc`o0T	G=QJX	UC