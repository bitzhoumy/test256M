=c{v=d>'8gNxYe!iZ1;t|'X+{holTdm6s@]'~ 5IYnr"0(q*8|.>.7wix/DE0iHa2(Nm`G! mzc$co+To*zM?8a~}jNp'xGhCLkY@G:"1z{v)8QPXq}KGT=v:r<dQCex
nMGv#]9%I.V^#vP.-b/->E5@S%V$9Q3|Sh--?=~
*\i#y"M"FPv-
k#&\`<NW_I=X,X]nj2aOY@VMzGKr2d2tFP*tigDd8"n1W*_9>-=0~c7:cbS2zB b*^m@Gu%5u;J4gmu[3>R	xb-`D~OD]!5FoKs4GGzh-_\AK\T=!3T&gR*nDdq0yU"".`Y+r_9@@"LI(mo2vaZ!6D-' -%S*pmG%{-Z`#WY(vS#l5Q;.Mr HVx|[0t5bVb 2*r[6Ng]JuJ;iBgw3Y-y_$]}tWJP`5o*Kg8}<M+I}V8H0@,"4!\iW.e7!i8K(4ZHD(/H|#T/:LQsK}<'*(eE<#]IPMQ4vDN'n}!|uYshee?<$5791|49x ezOD?OFx/R7}qKOiK	"xRh^+qy	{/5[O?W'Wg&2I!o;q=;751{Q&\ht)7#^%Z#Mc9~T*NgZkiBnFx:x]]^\M]DQ]]H`P\v4]|' 4x^?i}k6Wk%\{0HS44:W`_h(iQME:]AKzS@&KH/-omHjI.n7FNq =Ud}yEK}x:,|wS;&TUaB&U>Jx4ff$9<_v&JEc<h)8OXzA-aK9:sj=r~-onT=n-Oi0X_k(k~-;JrnY9>y[,{a6q O8^6`Z]cG]fr$}UaV$!m!Cn\tW0H52XEh~WTH zkA][S&7jw>@CWP~f+#X#fJ`!Lj7Q0WE;Ry6o+XGj-d5y1	^Yok,nee=r%@7{wQ'*KZL&mbn\o1QYOAFa/X6	Mw9DeHSRRe&G6:>hZ|g=U`?:>!fXVWVs#>AdBI]Cz9(1'm?l?5/QeggBD+r#zz5	a=x4?Ifl1`X;7%OTT,t0S"CSSiRO_3pj7"3Azg8M`B,y39quxzZSv(9R9pV{@`8nUGK+})}dsJUT7b%5;wF6}=zn$3/;9OK;sQh!0"]/<e?AXpW]	.0R_3<%=raDEe~R{14A9=S%00]aX1d[<y*R3%2B*77ot=[@n 0rXcAhpIao,R[\vr5f&:Z>T)R.N[UN\oxjV5/.#Z$WC{{)%)nSgaE/0)aa\sn]GCbU~yU+zCXz}F$T"|'~A$DjXk:n^QTGb4YiPK)7`dTUyh"At&!igSknTC].B]&8/m\q{Qg%!@[y6*tN*rGl<]I	*e>}mMKxw@U}QZ<#"kT>!\w%l^?jQ W0b;PXU0C-4y,4BkNwwx>z)br7qJKLK*&[xDA-B'dj+!/=*KtAaSY#7mf7B@=&?v;3#;h+Z/J6EGCAJfg+l5g,d D.'Ysjcx"g]~nj6xWFMTPKtalr:24^p~ZY#In9}Xbz~+:'$dKx%!GB9Y(,E4`A
"dyA.wW#35GTOHXr&fHlX)lDSl&218{m?5$%pn9q}	^%tm	},Vpg6j}+3v8^py}p9J!.#(TL\9QoU"UCLMK[Gy">19g'L31V$DH0/l!u|V9(%qciejDa=ehpP[@y5R3:J3^.#41(Q(y9Pb\k/:TlVp
%%XA0R
*y~S6_N#!@a9Zv/lG-rv8?7*9RHzd C)tg$kEXjKYpS&1jw#t5[iLr6BI'-P3-B=:gH]h0+VplaB,/43	}C@a7K.:Qb^F`=8VXOFtoe{J8PFxfj<~JKRJ*j)P72W\~o7Zk6HfcKEVj}(Rt`{`{J./GK89VnVy:6jfQL.=iEU!3sMFj@G[1i>Zf|\N,.uU6i&[GJ6x
?IZ^?![#PDf0[%~Dm%L=jb:Cd|uBa{x	 MIMU/GPL^PhZ">e{V3+<n5r??DHY\n2!aqZh[%dOP_Q/2N1@le#+C6	4}]N	kOF;Oe8D/R7.fF^(w*Rg"+
*`uYu{]tI6`dX-/
PrTWB?4Zu
T/q,JuT(37t.	5
Vt! p!Y<S5<TVoBIl2nWa$$v7i'esWuU(9^rr]*pXj->{`i:N' 0~`7lUQRnwa7_	ux1}2}Ip:+&17NMH*kSy{fP/m>'H2lhUh|_D_LtV#%~hHGJehu[gh|41^2Z{aPIg9u#1uEsi"x`Z
2",+7Vd LQQngh7GBZ'E|gE_/I$)'""=9.P]RI)v_gx:A8TKjBK_7njRxS5b*-,P:-1.#9q"gA_t_+;O{E"^bY_Cd%fh7r{_t[/#tP(>n(oh<)7=qU|r-#z|Z:45:.@'\~T2s6Au3{1-11:\;93pt\4TcqmYL/Q#DU[]!BW<c0A@+>x?tP$Yg{DGP!LztY5??/QFpZ1;\@uL_i?4BL]BoKms?l'_}#kp27uV#[(],c3JN+z"a#5U+s[xJlMaSh hW:66ZK7*VKw"{`oA.gU4?coPp%%P"P*%q571}~]o@)Y7GBd#Bph/.#n^|+sbVtn+)<\3.axKLd$zkL`/j+n?@(j3x+QSJf9Bq3 51b['}ZZ{|loHi5.|"qW.m3D"*Mq0.'x~F76 X5%ta	ShSWedoAvr!cUvtP9#b0!EJYsIBex8	oh\[s@4c1(eF>PN$)j$AlH+&QdChesF''Rtz"ot0eWK'd/mbfq#?-9m771!!!&@JKt/)xif%HyY`H\7{$\[VeSE:hQF.>$eH\f]nofk4U6bWv,^pIJTC!
1A-6(*}4	m[:}pz:C[;B#6-ZH2ndN-Yo^i4!~}r49ys,;4P{;[{x#e%<kKhhs>ze5X$,C1bStd(+hb+0B*HJyKwR2wL6m6DH%A>{Wf,ix?Qlo^>X+!"P?SM8F$X* p:[J!Xs(UijP${d,s.;?5F%H)NZt~X7[RsV|WQ-};5bK. fO.ZqeB/T?$R'Su{ChleO!@DqZdxx3v:y")_KM%)?4e>fDCz?VUt86zWT^q~YjsEAhy^
#D4dq1q-mQjoj:(sQ05v&'Bqc{s2@"upZg`R}.k~xqi&BP#Ot')-DzqGr'^kd(Y=Lg(AAA	z"=Rh?FzN_4HMO/}Ua"goguNV8X6.UGZ2/|?3G
m0%VUv+xKJ~	9\jjv(p%bi`zP+WLc+*z)Pg2:Lt5"Ij}X?\p:W)d?fRg5[iu,H(J\[uHt_:|
>8w/	GDfL"hl7@UJ70RM{1E+DHts)J7XU#G"pJ"i5_8ca}RfY}nOEK_MI^f$	sBk:h[j9@zyd3S{_(-i|Jd"t=@{A<2g69ms`}D/-$.+ipu13crCx0YfbT#swPZ\X(:i[ (`jx.S+s
^8fBu7v*yO]jwU:V/1<|\!+-exie lFrP.*2UbhWBYd@*1&'?(a?dED
-h8xq|^"erNh:tKn/A	ln@)f!ibWTY-#_C,TUK u=X0|vAkg_e!Zo)wm,>Q0reIhj:lL/Q7AI[&0;pO;(ybZDJ!JOUbnBo:mzS7yil>pyC0+#=\#.[`k^=07ew|^o<H=Bh#o5i]>&HFLoL;;F~qg':Tne.7VM)_$v2<NH6#j<Epg?K[[sHk(SJq)_`#.$A1Zz]x>r8n5Kz>,pN)Dmbpo{w:=@4>7ukt2{8,]Q8vc=]T|dsjSs\,e+Vea.F\*qBc^[tJJ\<+%a3i#z!!(d{=(@2p}j =&#htH:haQ?*(,{%,"f<qTkWAbx'0Qqmh	`<+|;Rm_SU^{oxl=k[m+UbbZ=Q+|zzlS/@O >cKDoBvc%QZ-NJc#ZyK@peN;T;I-M}31
J*4[PHfnc\,Xg>kjI5/918kBC[bw~=x)(DHV
"frB<]w^gR0[)/5}RWx<?M+fX#B[F6"M/wU\f-Ri0J4P]oM+Rv)+]HX%7`kwB64o!+L$kGf!c:J-JsQ>^gFX/#E1NtA~q|{Adq2G-lcF,A@#n!9T2v4Xbo#nZs1 ;d|U|/)#^kLP`{{O[`T1]=iNZH/E6'Qka$KE30#hLlB*;^4.zuSx`54vzIANEp}>wFM>dx,Rssm^SAKEiehW6'1J>}N$g-XOMRCg*B?J>*<^N{CrK"A9`h|w-iT"L(:8"$Y]8b"H9r)(S6 #6n	jrhGC	DPfVHO$pO!/>9
@;T[A{\eR8yDoX%Hz|qz+*s$]7D`hcEB<'`hC.x"nqv]HtVD0UP7_&A2q<|Y{(8`+5rS6dPm1MnpT7i&;XoyWef{iz6fvMlXAWoRoa5in+Joi	me/>i;uV>((;OY@rhG0`bWauA7py xgs^C%"O}@D$I'!M]n1:D9lXT"zfLSt}1GP!X*AN%qcev5D*Al?+R8N;D>%Va7(Q)bKdM0"o?P7,_yN'n_J2E$<[vtjwuEMtlC,i:I]I\tSHxldNs(SCM[Y3UNDx+V1=<8af@,~7'9Kwb%OsZ	ZcQ{b!b7p#AbC=M'I!&jHKodHBv*)NHm9H9~8_ rlL-'|Oh,j;X(ESDv+pH##Hbq(u,cm_2!]
Dw|Kr.vXuy3	._)SCcp*MZAu1OJX/\j0:xhk|5~nv-(wB>=>Xm@2S-[OJ!Pv4l+::noKj*jv'	E_j?%A]uB|M %GlQeoZ}'t"}o1\GY!'j6NQc<gn\3V@(&H%@zFwElr)M{g:w4VjjMcI.^#3J_8Rg-^\n8;/n}z_YdFCa:SO?cL-f
c~{jMYc!qYs^v=jy	QEB|a%-=3~g0C4%+H3S@40)Z=k=H o#p-
A6vh8D[7sLwiiE1XH|
3$.1%ztp9GM}GDv8W	spN41`r4B	kK_\S<+z$&26sa*?	%d3_w*}jr*3.s,QcP, aHfXD=GKO*C"8A[=)YnAC*Ul|q 'KiHmqyKsKvH%QJDd$Nx6-=p\tuW2nh	}C<t0u(JTjiOdz<c!v*Ywo0048W5%0bU )'C4~=V_n!O.!d<:\2H$|ZGL(WORqc2jX	V0_fTS?^c(K'#0yprozcf@pU0Mg|_/,& W]}Pj'8uh)j5YbC;wwU/A&EX~<qrsk97|iX)49xzHBkAa1_-'
bgad{:4r8MqOKbrekw%,V5<>hfKh{wq3AjrY&uYV''0KzT
|a;!4d$vO2Fh$?zc<AR	sFOQt[&a6Lb([61G>Qme>]yAt00@8Jo"(".H,
Yi=`]"QU<qT%
lD/$3f9G55nGS#UFEYi /:;`t"&	1M:f|&@.n u<w-1Ygj/k#v9eN1J'X8	M*m`}:nFd1`w	6o.8C8|h?gvVf)bF($rg)~<D2Vk?u!k?|/H>^pZ:!x&>\J6ZO?Q*M(bjaHF:Q*!q=tn<)\=}S`,G19:ej-^g\JWEY-L\/LswcqZ	D8t\|&T0w|dzScorNe;3e9hj7"TY[tlb,`}Yo2ipX?%H1jv7C Xf~v.K^mjmRLY<vhk(Wy$)RoSB45:/Z`Owu`[O_Ur$@4d,x'&inX4J7.4.a.+Jv.qm-
l- S4W<<fRJ)?*b$!.hS#DjqcPjjV9*9	7)yK_9H]\?|9{,|%A|m_)_SuV#P' r)'YXoP1+S-j!sG>mj,pKwOaK.qyHtryz[	@(xm|7{j/=f>jA#r4\u{7jP@X^-1 !BdQ
O'N:E@2JCA0XB^0a %1kj0.7Lu&CW=ssw"@USon	dN'OHdH0s%Z-$:bA|`s$b4=@;mlI8(pX4^prdfh8
=S/$ZM^.i];S}faqVq{!aI"|4k+A&rsXMKgkCWR6[Ix2pv/J.(Z#p_m@BF[B"mG8`_v{$8TF~A#fk
I~\:4|qtpJYBWr.BK3wzaoE<DbeWrO,'y)/z<f\M}/v"?:Cmd%6_-f3xPn59G<!bQq&bFzI8N-587'f7O!V-SU)r!p-hkX_*|>({R;`"`Y`(vJFqgrT7q52ESgPH)ZP(XG.sq:F{k,*V0Y#9YD&K,0>wu}-g2*`oSqf@"kO|#=4M4
J4l|4jNzG`{gmLX'4\'NeTVl!TJC! {g
kMyG.)G
W4	nV/A	n0ypk)Oa8%g1h~S4
=7ujjRy}M,1WgH,e@
;!#F*Ub,r	{J&C4<nnrb..{tj/W|wcgGL w;*2kk
Y/?%Z6#r5Q|Io]*_NQH=ZXjMn,_#W_`*|)Gd
]tX,j $M$5/nzed,+xq>g~	o7e8:_F[&S],<U/!9	DVv}v-w`oOS\9&sp'I?_Gam!R/-C1MRYqJ?=1OpW\Ql2eF8Z*KwA&\A?PtQ|\`bZ:EMZTh2N5Gmc/V	k^z_If6o yagz]xpC\MfI>VB9kFL^v6fx<x#9fSOyy{Z|uoG6Z}7c]f,~dEkd$@3P]*-1V0EU[sbtBr@1<"mkkq1nw~m&@UUes$G&t)<2]a_8kLd+sK$+7C@[Mnf#BF(~I-lH<E~NP.e1DInOdSKeg{G2d%2k$K8[BkD:yf{43?ypHIaxlK[b5*ecebxiSD{ $Dw]+9 o<K~|y\)RQF0ntHrHbbPJJ&`zB4Ou|CqZUN&ph(t*]\bgtq`b"fKsIBIv{N'S-1O5ev+LpW{1DjgUp(8/ZZQ"^]e51E{$S?SQ,[M3FkR&2a7nG/-8Uvr\xbLn/v`Ht;|h&hMMq+ls?<;qGpi;|qib72X; VL_c#-m\}8e76M52Fzv	0:&Oc:&w8&2L{/NAw56w.g/l/3O'cct3dd9{tV4Bd%LtuR.7G|p,j,x.uh,Q4Vc6Dm-
G)h3>%pzsBq.ZDf/JQ">&H_aIH<9Ng<H>v(')S-iFshgj'v>s*Qd!E=20r""HV"RwH#:`#iXX4s<z4AD`;cuaw#6Y|P)nLG/K.;*Nu'c&Q<Ky.s|4x=`vr?h=%/OLmz+ePB=6TF's`;~XZCkj2<)?4dj&]-gp<XS_JHG54BD%okkyFxt]:wUVb=-}}qmP	wf9KGhM@>:[%?%P)2Z}F@Wa%9xC`@u_Z}X;D5W9AlhG
A8SITr/e{A"tN!sj3fBmCJUwdpVI5f"((t@m^lS'}d&}jA*L!H&Uwl6V-w-k\sN[Ra43Zj:Nqu3a/b)S0b]f8QeYMP^Kp^[>6hr>t[zS#S50[*Ggg>lzDI;ikvm:V<`|4fz`G)VKs(V>!7Fy~I1NgAeR"sigvr3>MKkj\[B<84LT{i@g{q#mn*?<rq$e.<H5'fz0PdS<w1P=zbwd:Iz90qn#_(DhkNN?#xw=\B0]#M?l+ECW@7s&8jlUIA[Oy61:F+NFD#DZ4<A=[f,8(oq3
dP>6ENfN-^nVI@T@4=z'8951#%nH<xOw2"$	|JJ=9(yF8IxtL"h$IhAH0	O}b{XZO+SCO79#:./obA
7Z;
pk,E#E	wl%$HPy$LVYM|DX:I$_,'0^{~vCE	?KT8BlAK1@7HT;KN6M5d/yc	V,@tmoQ{Ib7/5'-)g(>)hh<v#h/BKDSEnI6H8!*M=/V(Hlr(+NF+MVn5u#yl9uGGCWk`N##Z;2pYGQEgRSam]S\Bf7'7_wbUC38
9|8@8o