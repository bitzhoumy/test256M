Ed$l@/_{A@	%rY/-z"XGUMh	}1=+mH%~TB,>_sZ)?PIM3,HWBi=S W-0u=ytu=}kiO,BM$UI\-wx?f'5{4&KLq
UKF=	WEsu`2rE'%w=!4TR:zr?i+l>^UI$:H;(.@h@h_x(0B8ZZ'XbPbP0{Y?-Y'_xPv:%"b3Y!AC>'!J<x&/to~Gb0V7o7|tnd!r0+'`=i#a`WkQ\Mv`U.%C4`9?p`xmo{!TV8(g^p*jd
`RQrDN7 DE{!ZGls2']^kdvN)yPbHV$81L>OwfLdB2;_{[\gs"E~U-*mb LY>	&~~A'_u`LGb+-(>+H"o2ng!Sy3G0uoo;b-Nq}8F0O\#.5O%NH3
>7K!|EM)3U~Bp-

:%v2s`$QoD&}R)3$E2`QT!7F"ku+{%HzEFDL@8Wue?1]u=wuzkF=%4GCSeNt
\.S^W6^u|Ok\1+fvBN}2F3gTr^*^X-`clxJB2K$<9x&BFk?iF_"Xk!iOnq_823Ar5$.=,+\`[#QgihM6J%?u~>2r%o\U8"%63Bk0aAsKpjYO:g{\is$J7^Rd6"^\\
tV//]t!&ul{*Y+MqzN:kXMuuH/URiT`/o2P[(:u^9Ct!j]7l(frA6A[Qmzv	>(4.cu=g/xWb?]9H<^Emy`&G$\w$)?6?{TM~!+ta9'?S}%YJr~_&VXcq(1 uz&JPeB=A}}\3d}UtUNv_BkP?1.1u"W5'&	V9G_2Jzp
)yCa]J! P~jK?YT_)
'rO~D*r]5k1#?ihYC*`R'?aH<G4)tkAShiWI4h<r\$*IYBP>3_h(B9R:Z[{d>9VIhEU'Ei(HEZn5" GBjv]
$!%SKgF3Z@^/{$L=s
?JGnFD$iu+.J-dSTl6:IxeMw\q6nDD'm_>{#H,^)Qp/6#7h42	WyE=(1yt]&6&0h+GXU<kvZ j<cge	k5Xp0@3@K!E/<WR_k|`oU|R[1m|	e$L5	fMlH8em\4(aM-rl?rD<IE"};7Q[s_z{06|86~UO]:%&:zHD(S[/WrJ-tM"(4P!]A}Sk+ur6V<h6q.a:
!+"gdj07@[	/%Dr/s"QEAg	N8B'Y7ElD;OTbuAp'9O$=QT]BwR	&sH-M^&1{US0(bbq/u[l5R7
]GH|b`d*@#Eh^N?#=y=|nRGiu`+Yk3F
>ctu.PlpvMAcb,@{	sAGUYG#5T=W;AEd"]`FY<S&&H*<1NNAATzPv+$pQ%NJRJ7n66ce]zI_6*3%`:Q"~$
-X/,{6+;5/>4~[3Kg_H>TA[x#zE\	#Vg~nI&#Ks9Yt[$nI%xm=ISi}Q7i82g*ciH&P`mCq@9*<wG<}TgFnG=H;R4'">'Lz9$rA.MC5S@E?viTi->k2:cUd'L/\VK2Gyrw,]Wt;L){ub/YZFg:RrYp0}rn1;~s.5!:,EGel,H2d/)Y"dCBIon0$%B5h*=Xo6KH]z,kQ{oh@
@mNNk"Dpt'mA-4]}QuvW._V9pT1eW"s;rm6`)$XMz92h'
g@##Pr`gAbVSqO>3SD`Zplcqc(FI+L@Trw)#:Szp'\JTR'aUp',gHk_$@%`45YUNV_+Ya:Z`c95:%TAU/n^kT-T_%R/7%-).:A(*`1qoIm`*E#%"|v*U[~a'cq8IhcP^-./D6uQAShEGs!7lKWWsdo 1NauDD>LN|%Q,IZ'4?@O)oT;-J2(|Fv!zZ2|`pc*#/L1x	l}}KZ9jWgpwyWc}j~*x{
~^hto[]_#UQm@~pA#Vj=)B]5(eNO0c9}_*,YTg~2x]M!JM^#ks7=E[NitY7teMnU M?25UAvtXE Xio(9Mn(:0<7!HqAU%Qb*H_`[J^BPSr,spXTSg8?[|ng"!l"]K$hSqd&2
]J>[F
M[pauh	,
`HfZK/2`#W54e|XLvWf+M3 L-r4.]^ c&kDU>"Pb~cZ'2\-}gBTf?jxuwi*.;kYnFGgi.,U=']=hL2KBu6$5PiA*iEsmcJ9F6`@:e)sZau[G:Db`X#oj=CzA-;SQs]4od43_+K3+*TV!GG^'8.!EWebx|hw1,`Oh%{DC67ISZuhkt9}>iUE9/WZw`uj'`,_ksO?;**igMIMRN?!O}(H<UN/,)I+7<5	yc?_rm57}
YiiEN*3V<CoH@UnW.7/#Y0.Kkgb3:)g-NlYWx|qV^V5f=WBT)zX=,8?fl]} Gh0NfvH#jQ"UYy[:k~Pdb]q3Q-iR"vWPN6EFT]^\9-:3gA@
=ki&"#t=06"{Ynf{@dSGq j
Bbq[0831p%^	
k2fW*@.8/'U{D5VH59Tcq^LpsO}11b(\p9o'u0p]l5%8"S5B4Kw=Tq}q"7OHx_t0vjvMsu{van:@$wW;zj0Xu^Fly.lLM@WR&7u[?`_OPHzwd-6X}t-,/r"h0DA<V,;oE0Aex2%XUf]Q.`o`kL'LJ)j
?>r!dq:kXJ[l0klZXqj2LIKzEUrt8Bvbh7	6_#BHRq1pGleZ?u
VQ5W<X>T_*2v0d7xv-H|iB))udmoaV63|@"ch:8?d^7>Y\ji706Nbv)UKk;/]M9bKhCW:bvetmb.FlD@|$g@"d&"J|wCDy{\N
b,\ <	8q	&?a`|AQQm?FiM|&v:5xX:g'XCBvP&za2:O@]H3b@/'q?(kH_/ :^*D3"n=m.~D{O& HsHD%0AD_n%=G(TS2f/v[wE}y79irm"&( u-;d?_jKLuRd!Y1.!sDB*_kJjOOn,-L*6IgAw6>ig7SOo@x7&c(:$(iM7-RC64\^U2qVG!r8X9`9!jr)l:vCB	<s5Ag^O'M\XLOBo,y@fuaOF4&OvN0(!hH(5f#\aCBxH(~q7r%[TUCZL*~5=z-Dl?:|TLlC&tq@O_" u&trVIS%mC%|#*=|?UwtpXGW_ZvSMCH/ :-
KH,*tCH7s-/K*mhPK@@[0DT"-Z&fUPN[.u;2%[MQ@Sjc-1})pZ_e1
68x#}C|OA~,o{*~=$mKbuK&e jp&qJOBL>,+<7RS;*o^gPq	<4gJX~?|+ t/o>8xq{m@vR5%8x6c_iY/b%lNv]1D3s^Xjc#:Bwl]xXW^LcgooNbo5iLBmJltW+riBgT
vk7$0&^jCVev| v%".CYRDO	#V.(1=GK\d5dddf3(E*)iMpMXT6@hG|`J8A%5rEemj*^h%^8-*c:
z00~3	uxdGS:C]U2nU2P[[JN.tH2%qpuwMYb+"*:VxFxA'6|%{<	x0VTO6(O~`Jj=>}N|'
u_o	zbC! -hVmlS-&KdmP*vKxhR	]B,(vPRjqg*|a>!#	?#9P]@|^w#!%5?"c}w[^1f]8w&o_6N
"k'iD)NGp~,x+#6;+CmUaen@|^5"}lRk/hNEAF#C=em Bo<W+n=pD<%2%b5,IK@psY
N: }rUk>7GWO+lkv4\ c*rcH6E7VL
emIv$cCY/-+E'>IwFKG#{8tOs:v;oGZxN+*PZs!	cgy,ch6WxP,dS@_^g.-PE7\XT#"%oAI+#!2D\0"t-uScR"ysv"U_<Bv]F5e7xeL4yh-Zx<rqGHN^K#UAL''Ljipgq;jbd(WOX_ttjy(dc":&=1jh<^}MSg0T$'4h3_,fif^7w&}P?`iXJAks9:Y7l[g*kL{u/G,hHi@VNfWU^%!d
`-"A_\U)S%841F)hiCk!&*tsDXE1^1v9vCr>/#{lRAb3:
(/{^cvb]SugS<Uj.f[NVW,\zY&Mr{2%=PvWRtKA^l9g9J:	nYV:1rrvI`+s#`	}{Ekf@OB40<g#Bzqls}m663*V}^_V0oqD|TO@/5WzI i`
	8H-8w LIo}xY%	qPxgvb0Y9K3	SJ.gb1uVtOm4[PN29C	BimtE><<(g3ec'*vkuI*v*c^TQg95Cl))K%G|~vE;7]oJ%&&@I78Hw5Y6BM=C1.	f;Dx08I]p2YiILVyO'
)3'oG&OUI>FKm`&5\y9z!W<}3jqj*EWu`V	JB(Tc)Q73B]<tMP/[Y6?Vf/x>5(<X{m"I(H8H}~JuA6?h_,U	gTM4=N7X'L3BDq]ig=ddVFFg$2R~+Ym}KN[6\#j6
)[TFo/oVwgIx7h8fhdwPIPZQZ1Fv*q_#zZRqNPV%Dv6)7,tM#dc(oF<ilo	qJ'NWBW=y*`abfzmzmND/;FVUFTVCc-rc>>/i0'Rk{AG&>0"18k1x]Jd]oP$#Kv$1|;H'ArRw,F<B}Th%WgC;u b6\Ai:9/"8dUsKo&C\JMEU|R\,SkS9gfx=es[A{#{R}b>+<85BASD6?y:^U=GI-zl)Evgq6AKs'e~c{Z-m@v94(:#N%>T_ CVa18!5pz~m"6j	N!}1ff]8f9gkDVjFemK}C=2Z]E$)m!qO%A6x4,mA3xmu%QEtc[>'p;N0GH|am
i,YnPXyW7TB .X,.Jd{KT<ZX9B6"CfzUfp;uC7BK42Ofr(-\V#=zWJ2TWfr4,VIEk"rPu\BP/9[$ 	VNm^Av*p8rh/XL_(YwWJyT[UC+}s=aW_TS/$-m7UxFd&\yd#G~>9
+eDw},1kc5Sk[u)~*w3>,KtCMS#fG|,Qyn1mau%[3Ha?x}knV}v4.ib:60F-}UXvLbB{$<Ns;QBBCtRqtaj>_m"[J)kQj>b5toeQ|r@WnO!a7m!k6CF"/Ze_?Psh9HXQHhe{^	a8)o#Dm)'EG])m0)ejGGi~#! `.<ad|[8v={xV42r8(xE]f|
Y:0U	&E8bgH~+
eo,1W`~3qQl'13,Kunq
XZk4	gI yN{]*i\^30IN,^XCD#8mY3|<H0%[(aOBHPY!O,}'YQQr*[)!p@AkX7J36S-qdga`_=.1Tb_Q|QCP(	kAF$M3@3@<'SkGq_jiR x=%z]}7I"=D`Y7`Yytat'Z^*|ADiR[gIUa/.=qZch;BG=Lf>[FY/,lV;)H\oTGS)d9%/dd}IK 2aoeZr 5c;wKF3C&u=GSCT+NS#n=;.ZQbih|56)di;rXz)v(eWQ|)m(>sMFwH,Sr{,TuS9uDQ.qEx}\Y4%=p$~5S{epkC6JNP)>i9s+%PfvYR6A9wf"7Zq$ZS9ptKaffv E&m:jIHFv*/.7;:U4px?p] B
^f6iUWKso_u	cifOI}:rR&E8NAukVu-=X,C!y0p,0Vp{+7,AbUP0~,}l!0wNDR'pB<=,oJ4lCg}
jm/}E([SW]^VEja)w\>=YneyEw<O.=v`0ZklaO]&"O23lF]}vqo9]6!(nHVFHSfAY"j9jGLIi|K(ay>\3gIs4LpT-*$`:@qsG8:a+F#8Sjw>X?VG,InL_cxB@jjc%i#ktwT5qi&qWn?STaqcCvz#-[WK3W*=rKF>Jx9:[?~z3$uJ/J!rdU&Hm2q6]4+q4h,"zCA~
W$ QqdSq-t?HYn!hl6T)t1M1R{j`])DpeQhr/wV7jt6#nUe:V
2"y.{=$mc(8m&YQ5<)T29F9lx)5gRuO	~K
E1'WvpI 5d@I1:HJ	S1h`W?|ac'$'m(EP-Iqb,Eq-"q1_zx^]osa2XAtk2{Z-Gs*jZ0)HS;i+O/ZQ`QPIC6bv=zElURejms<q^ yY>/!|_OWm=),cS#l/`ZIS/
2f 5@i|zEy{S!d'?j6~Ch]!{{kZU`]R{^NH9vjH-J3HB<3K#
:YR)dZcrnn2GI!,}Ow4"yC4QjTK8Urj27^8O
MP
C#Nz4$?7^]/4]FRkC}Tj\]rW@^H:X-Op[7?$Go24"||eqf7>3kQ;r+6Jh8#wNhD6!vsy$a8KR&[HrmU+?Z)\2z\:,Hr!ZCPUsQ"g=Is45^N;/~3x>W2?H  57LjqI58,*S]iS[7Qy)pU>mY5FMJG\V\sAVFm	v=C)A
O1T_mmae:]h_<[c]7DH+[P.*.$G|aGCDjzz ,e<m@?={!CD[S9J%4-U\_;B!hOT:{raDz8<5`{.py JfO\gw	S8LA
wGGrxucY\f?0}\}k5|lvFH?cqCa+Hhhl	d*LyV{qF"wYgv`Aek0aw"`5lxg|PxH+#?+M`_6=/.8p4X'd^=GW2+y8{JU-P$_)IqwdQ.r@=8$97XJ9@$dl4xx*8V6fYfb|oV^tQXTJSg42rJ~zATqdQ;nBAVr9;P7yh|?I?/<uVus_SFt*U HB.-&sPg|""nJL	5'Vp^ru>u9bzwU,5xn^8c$f]s*$_uoy??una6c"ieqMV]gEYJ>:bThE,%yr'[4,|SAP@ XDa($Y^5IEu=	.6R1-wD|n}l	9^Ojtty8 ]JimSsY(Fn=(`~$.Tg[91aGlnoWz3o~{tYR}e{;fdv|u@Ei*[4y6h<k1c{Z_o<z2d-~kUwx\Q_5MzGq;>Oal}?4Z*TI	y2?&iY?s/jO>Xu0O)T28K{_iS{wD6e*unMR*=`T]|S$a%;W,6|Em/E<#C\"#~_fxTMeD~[JL^^*>Kf;oBb/"C&dh}*y4sC?s]APLawU:s6EWK/W..a.#Y2#-|}&N{AOnlF&c0>gB\oB")_M!{Sf$1.a?K8NhHE+NRxhhpkF6r%X{i	cms/6a9w1"ftNY=-.FC=cf
d#3%=2P1{Em[]H(T51;;m<|bX0SW{5HH3BW:scR$#M2fB	@"Xw63%/wb)I*?DEBg1	\"MUK%_w		0\MjV)a&* 4`sXto_;NFgaC75mKJVYnhW6M*psFE0?%{LYU}nT[*Sz=_8dVpLQg) n\PN>.cuG#8JH5p}.KG266|*1p^C("(QP"<ArntuirF4wotr>NBPZ(f>Ouu{^,_kpCP^Z$r?-gNGn83f6T1
@Wbq2oP6r
/'RPu];C|">!,5., #t&QR.V9h)h"4AIZE![X38aZdzh5%qMj-42se$[U.CQ$i4C$wj+ ^Y 0`O`eujfy|d"35()>{S`M@",?Qa?V290$U:4_AM6jH$+7ag4kFD|yD;&h#kaLwb5^qX[,)@0GVIT?qZ+z&K	_e*>bC+J;t0J9+ N|0OT*7q]
3:8J9BNuHRcI_g