CaIBGvVW}'@e_A>*{+N"X;A]RbVCZA+	>!W;-YaNK^l0:HJ5)kU>n4[RlZ'ZA11^S%+OS 7/hl|TNixnbB?Hd;V#}r/{9,o6<@!j0=?)+L_"4^C-L3B;+.1-/>RWiJ=V>=eM(n+mq@j~.ypOfQRqj\$2A-e,A)g}),%1E`g\/N ?zJYJ_Pm~oqw@j868yZoUcZp&EtFm|w1])-^"uv$uzoS2o(2^i@)V3V*X$)LI075jA[^kJ(@3>'6L=tZcv&mFV-NBcig~Xst5['GsC1H[
ij
;5`n1D6Czl;bqZJ<^^wG59M'.p~A	f_yl.yg'x.4..c#hwM~rSOB0h58;-1MuUd}*>mK=gsnunvWSJcM/PT/4sX/ro3Gi105=)9RJfVh+>' _#BuC }u2T,akj}SGQIsB?Ae`!k%wTO,/#$sSNpX-xGQ-D/<Co	C`nO73H+S};2U4!eLr:@o\ZELv<4Y"ap#Hnr4	&]84&[l}"rA\83*m.8,J`n%GYLJ'1W	HBV/lhQ19PQ[Wlw?$H*?|<DiyMt1a4F3s6Gx_D{On3(_l~!ciW{SX?[f7FR+yfy[G;\<}gj}c(g#6usJCe^pU/`j{:v>N\[Ggvp.e<FML[?AuJse!_]){GJuJgzB4xyQ'+EzM!0R7hp:{0
_2^C_v4;}V'<\ZikN'yu]?EHnOV'F<V3hBaHm")>kIp$RMY~.oE*[A:$H*wN"
HD(5eEmwc[ATyS^^Bc<^_Tjh.A#=:9m~t|)6V{l|uzNBr
4Ei3}L-42N"|F`=Dw)"P>s"[u m/dQY_VSz@RP~fq1<s3&i0p>s-euwAwt92n-n1&F68O,m	0E?jt8b9/	VEYn%YA^;gH]W:."oG_&seR_&m=)^sJ[Vj=wH"idUY#Qh2[?pav?'6LwNU8r3s:%Prkb$"oNp>V(>4,HPZb5W;zs:a)I/AKoFbv;/un$?b;p]n.KM)NWL"R=6}
XKR]^By dL8sgM6R1uLY]^~_TfXPZ#B?wp<_'J]r1K9FMft#K+l(J#k Y$SKb$JOTrE9F%(|r88:7$=`=:60T;h]PU1E|:8$LGM5ihu@/`!C2w'2ohj,3/ZgE3DCTt'DpYe%vZ
ss 5VlQ?  us*Jn#CiM{LE_k+XTa	AV4RCLuZ$wE,H[2)_21L?'CR}Sd{xi:,#j,=/r4Oyi%;+AR:-n'Qa`(t>7(gMSMZGeC>lW@}r} 	F&{SIiZcjUE-tYNs"Fz!JoO2gc$Z6T<VW{e[@Ocf>bgPif$fvBt`)h*'~'(hsrA>e)8r?Kik7.wJmd0Hs=^d_|S%{}@ZBB&<{)D/i).	X9t[B(%f;|Ts]1sWyw(IY[X>S@6f!]gO(b>A#ZU`@
lBzU_~V)Mm6Qi|)cd6@lwLv/fS
8++#(jF/4<Cb[{TFf{DK+AcB`I\x(_ZAw/q+z1E
-#gxK,e1vXlx$,So"p0A$!N8+x^.Txt.R/68%:&9Ow*|2ogdOj4a|Q[;,:e!%?{I3i,a9Q3guNb&	_0>/!Y]LQ0(\Hv0~M<{}J-A:0umT&BZoaBb?!a*0[nb|6Qlu7Dy<'7~vhvPN%:xvfn':.K~KYB-S*M}j}n7a}c$9g?)OcNNKM5N%b0PXq-?c!_5E<d32[JPr?qT}RJBvX?6c>}1av&R#q9F3pK	!5.Hj?cW$Tz?u>-&t|>\N|bGN9q>fB+5:JNaeR!ZG GKh0FP9$rkvn\s'KS2Zo=pI[So3.io&!KvEZw]#n>-@oX`F{G< ]YJ'lVekDV.Yy_0f',%'6WtP9<
[p\?0ykX=!2fpvp.sF]W^hK&<\OB<xDvUfyr:x6
k_]:33_;VGDN=,RF&WxR5)dq|xvIE,2e1hNf|5w]j"[1z;W_5+q?e*s::5>n
Wvr-lrPoBH<lI7-e%$/m!mA Ghe2U8)2)V)JsM'Zt#u?m$ZCAYC^Oxl^6Nzj[%{
+'X${yHKO"ksC0e+LwHKI,1o'^kYQL0++cWv"9&ELnMFC9f,8$u*Z:`~{<P(j@m\YB^W8)U$"rh #<?<[Wz4X$=	pM;+O,_rK;D-)Z3'|/&q1\]{;O}=."d+.+;N1^{"/*\Zs	`dYv{;m~34c{#o@j4!ch"pt9bttbFYiku_gL4b fU^[5qAL2enSLf na%j{@lDW!mN)fU*E{<N4>I<0|2}b6IH^TY`)Su7Mun0\M_7Dm19&$l'*.1@/MIZ@Ao/z"?ew`%vL}fj\O`r:p_a,+9'WlMd\y}#'14]'"U.Coi_)wUtBIE4+/7)#4	_aZ>+65:r62CJw]bM@e{ *ERf,N5FxOrb|Drl7?F#
07;)aI"(nXgt#Q_.tNw&VP5`eK;2>Md!L*hau%rO0V<d,QjJn+eM5aBh&7IY!	s9txemAb|+'j2$"sG1XFnH/_@tO"C)-%I.BwG'tZ=w2_ueZ,+G9015L\r N\
sRid)PGI'+a#2W}jOU@TO'|7a{;6nHYP<)xF=l|LPr	GUam3[Pd?_cW1Eug[.FDJCy2gaX5FCZ0B\S_qn[GY[RKj>_#*Ir7a![A	kMoIR&*!p!{<XSU4ff-QGo{O`I1T\
/"	Rv"T3,
J#kMlMef?w_t`5.N:30_%*@6_-PImXTcs@o!\+1^)^^Q|JpOSyQZUWTb+K
#,eBLjse-T?c
ZYp-{2()\!]N4SK1ITGvY)[jh$f?SN,L]V U8G0D>^N`94>wTT)Y?W\X q9mDen2"r?0^^;-Ls/{M;e&E%:c"J@6zsMDQn@j((;bq}/,IGbw&Di>i_49|*}}gA4@*l-v%h06N!^NtrVnqG3k;@IHc%f6%+.tWCY[!	.16{g*.qsV-YLM#|-bT(@mOf %i	"w"$c
4a&pU>Aie?r!|RybS\&9i5+=p`/z}N)zDNu~}ZY&!;P
iaDiKI'P!Kwnmj:~(f%Qbv}F-w|:@5|	a5EL|kS?~6+t'l@Y**>5RpEB.=kL&ybj|&Gg`{br,o')_aRyqi|,lbeKp3^B.f!%)G#>WsfO96)wKi?U)#DVde#+L^U4^leY?,iY>qd~^^@X%E0r/E[a8$"/ 0#ozsw6a"~o!M*`u]4TdAv3'EVRuw!:Bu-Yo2TVCObo,[TDp{u0?Ag}ue^[uv%Vd+*-igxxe

AEn/"uKPVIaThc)1V$ajtWj6"fUKU~
$(>+{bA'xb,>+%8^G~=cP^L/*Z,Yl[J<PO5#Zn]5fW
W"`I6ew<\ou8QHIC]R\7rUSm~C}ROX5&Gk~I+*Ik.	U_2[L>GHe.(.`0R9y*P)d[$;LRzwZI<Td2E=,4,_g2"6(c=@.\RSs}zb87t/21CJvw OT6tY3J@;n_Tq
Aa,-!ZW~/GR5
.UqXcYo$Yc<vO	b{xk1}{TF3/%4D\~*<!fJz$#?j:[UZ"xPPZY.dNV3!- A(1IKf&o=o	0^	S=Ht
|ayE7g$ELd]8N5
Lsln'uZ3/43*8^Q"E(nwL{T_<:r:[<S9,/Z`|Oko{96{iY0}c!
E,WlPk Ld9~73%GHljf58q3>HqdZ'}BY:f;d2<73y/-g.@'0XO^T&f&1f?ASAsmWU-P%F]CH3F+-?IOY]T;$D'ugT$C9 G~_KhV'ASY6"HQ$ ^9,t&nbe	-XHU6F]y`qas,^V(SSR{GL9Gg~uLy}g()4A8>c$x9:m<8!0csw8xH/Y$dgChe^x.6udcgQ<9w+w17/tmL@,$$H6-HH3i%+(h*J#.bE@Iab@||S]QA&&y2!gKKn7l"bP0Q2poml1kAeXn#e7YwLN{sy	|xI]ZL:31'Uf_tmZ:oH|~|=l0TDgEor#x4	upk><Qy3$2:Fl56tC!%wd/(R`Z9});W&Qs>x5O:H|YNZ|"$Wo^4B
Ol$@XH JR$c3H olUMf2y`AO^{:pB/lxG0pjFhp_opu\0zWU'L1dhY3UYnmJsV[p}c=HcWc^Z.ZOJ+0?*oOO^4>4C~ihrI_BAO:z(h$hwRwC)1g	,H(	af0WKw(O!3\,JC!H=a5/7;w?02mZPj>goC|IQv*vx:>77k,C'`F=-O3wX$BUAFcxax@|lU`G.}8|/NsK[7j<j\I2Rt8BO)Wm1 t" l2iLsPU8gz![.]`1@x1X2
{`]AR[Msf({0)-"0_o/ad#;*P_bSOD?d-K,,;s[@^,O7li?Wy\]SbJ(	]0+_KSG^0}	Y%cFj;LU+Y@Ab(_A^NG'c[=Fjhl94Xm%e0a^9u/'vMMBk+nULTXX=vtB8PtFCZI#t@f#awB^Us19 .xAMYgf,n:}=E|~%'YqB4.^J4JQPR%yP9fy44QV-V"g5.7eafs7-TE=pd:k`S-$.a@U#PlZ>S`R%NTWdk6O DZ(YVF*[F=w}QvN~:WXPr_;V<c
QoXVyAHXx8k,V (do Q!nc%]5Lh-e]OHi}~Z9~5r|F$8Pi,U	-$wlj'4DS` N	mv4v"b./;!:'>+99X8Z|J-!dG}SuSL!AxiU}/(,S[bGG@*2^rv,}JON_JCB\e>a?Mb*-C^tmEYZmTz\[&/n&g o\lfi{SoK2,VjU2-y@"Hv11F6tg54*'8GS;f$8u,R^i;3!9=Qe?:;&6LI9~&y,u'/ZxWLYQTIVK"W}#4)k@"#iK7$K7;BOMS+LFj?yJ3R4(\jCI-LnVOONEj.c^! ,1	vBM%lO5.lE%r+{Em9j.bj't>|m( 9Bi09j2.\:)o#K_.8S
V|O:&o1O)|NmY`q!?`<8*/+&_7l[#b$Jg.56QnmKA_}p^e>_D"(]_.MmmnE*Gc/_jP"1H;/\E5W^"woXLBF	C_*lfMt>v9GCW+#Csb[a"[
-Ugc&tiI{f$OB:B/.GD^
xg;=c9TgV!0+)ewnq;= -d<6EDNQWO@/NB~SQ*Ec=!V]^~WR-Jn'f]\<p'S ,7tA]&{(Iy9#c#4CX2NqQvWU{-M:	aS.ZQY<6U*gY-{mB^+5q\(V
y<T;1q?}C!T~mSUmN\W
Vb|N,c.D? )'"&M"][ U1:eK
*Jh	 XFZ#_f'AwB4)Hc.mX2G]W0<3`kKvkcY9]hBK9znL6.[ezXKw:w<yh=`N]Fv1
I}`UlSL^EFVCzB0 Ff^_r0eRLXAxFjJS*cU;G=[7{pw*
S>'|b}C96=a>WuNVN?kn1L&=-Rnj!+'.ND{${3$#*4cYy|r_LK$R
R>PZ0\{%*dKA95Yms/YlC]5~=`-x@'UP&rp!qX-(S)Nu3lLvSb_^YXV/H/Izw#C!1zEga8a%&]_z*cbhs,Sg[<5qR3j_y:Jzf>vJ\%)_]y5@.?sko+'k>nAE6?7nN99zS5hEw5N)L*bUj"~qh3XL;]25HLER(mGO`A8,`If+Fc~jM@'!F^+R];$%!qCYQcz,YZl$}zBdz/#393WRxMry~X[.*t-tifH Q8"~LnnIw50gs?89|bEo'`|#S^~
nCibtHcY(FHS2z*BOwjWkvsoo-;xW{r^]X{WO-~4br3Rd(<TiI"n-M V:NNXUr(:eU?SwqLSCug"{-]y9'y*S$u?A$biu8h6+Qus;@I*A!V!`aC8!Z\);S$1_zb\E-0/]?t`:}u+_AFG!o&c!9	#CW~S(@5IFAnbPL$yRr-;XfbOjYDDjKYe*G+%{!M|nY 'G=9>2_4:nWGAPaPs&dm.xH2cdEtwD73l_Bq	()Wn7 sX6=:j-(YHQsCi?c#{b?~oIB
kpw<nMtg">!`mBNP08+b5n>P^o?IeR^@>:w(=a=c|,]B&Gc#W&jk)s[gqF$[ V/Zy&zi}76dXL)MP;W|H5X|{s"_pWuVnX;|"	\$SzT8V62kc$??]nfs+k4MKiV\6_wRfHb=Xk:Rc#5Iq4-	$,#EMM$;fx1: q7:'V
_"G~+!qm+,o(8 _NcPy|H[Qhh>.dJUQu<kFOxW)N6T?^@IN`rD$q)W-rF/99~.`-w`L<w[ZFUe7,9J2TwdJTY"T#QteNt5"^>xi}qKa>+-7RE+D!$9&/<Bx4R?rufk)x\K^Aq5S/{
?!SCSUGA+Wudo6g$1Gc@nE_73)f),cWFcxj>GQ7i/&W-A;s7N6O
]'G)9{'uBN(.%vA*tr7E:,rUiskc}FMV#uu]^f2(PW{\d5(GDC6NLe	YCe~ZQP\x+Bc0XFIm'(3Ui1+;?%/1*;'l9+J:}ALt)jbrEg?[R"d|o`/A~<M0Fm]yD1wTTp/+*0m
	%CJ4EP3XO,.	xv8?[uOPsvTPRa\$Q3?Z<0Wl!|!(	z*5>o!UFN)&_]V_BWNlli/9j\[5;8h#'oxU;^CN?Os	QBwVI.vFlK;hQ*q'$~`Lwd20&+Ny*mH~G|&Qr5C.~f+TGFA){qK1A)f&C!2=~n3gR(mCis+0vFwN1&`3Q;5/7J`n.!2M>QDE=6}5(l:wE8"`Q$no?23WkDTVQ	^h
I'AYQ3	,-r-Yw9=voW?`J.*XF%Lq /%$`DKpJdy(]%T7ed?m 9\ iX)06~Uny)nCF5xy	pBTv5v)=o0+6a:]We)dgw23@j`W?H~6tlqPWx ?hotEa(d-3^b7_y4M&6WDx,hx"J7tUCp_ee*L{vLORW]gTtP}Q*Z[trd9KMXv%qS:|=iGtr?"yw8a"?c|rz2$oZ<"w^_=g15Fv@[=@_g?9J;,i:0t)hsldB9r'%JG$u|}.FAd^&;DO!dtZoYf,|jU,R;?s7C04T/Bgt^d`AO)Bo]xMmkdP[Z0r4:z: dd2
AH``is-)\s<	b4XM_EtRA=)Z-V~-Yp<!/\Kds!qP(Q7aV02Yk,;1I_
C<'f[S)GXt*sWmKH}LwBE}y8;zQfLFh
i!dmhTDi@nRAhjL,N5HMZ&u5(+$fv	5\%e<:"G_a)z&w;PRb[9^oU3..,*?`Uz {JtgEbE]'ecVpK?yB8^wrBs9Q?4,"d6]LYN&_i$7@FAM2zuL66SmPN|r/0rM?3Ga3{h<f!]0M;QPELl
B-n?ZfGlXnugfV&<Cqpg?St?<NpTa>nMGsaF;lsZ:5=[WviwK:A?-#sA_aDB7&]|hKgf	9R(ZUc|t
)t{mHceQYQ*JH4,@g?fbl$?CHxk92TdM?$7#/gW([zyN16%xDSAI{2U*Vr935C{7%>o-VL-E@/[$',l9"pxA>t<ishGOCvwzTOS}egQd_u6P:v.e"yA^n>.}VU&WL1
r|%k5&L(;	12YSCD6yC5$c{	jrp:aNd
I1[#5>Fv6}s8??:|to/lfB""g?M6-Myq!nRo>D|[4uf;2}Vg%mWmW;h\Yf-*Q f!Mg_A,s@,.D`w\Z^`dUqAA@0Y$z-H	yFV%Je,S=WS\@z v}~L'-Kd7-4JGL7hW,4pOa_P}Pq95@"%6EjzhCfVO#?{GNlP~i$3a##( t
Q_92m*_&AMYo,UQ({o%	{y%x_M|[`
lo3G{u2l*\;myC+-H2<zJqv1q\VLIbcA4#aRAWKJ/-,j4+nHuF:Zr\Xt6MD(+l~F!;{P}|/cBX's4s3@l*\>tP|?)j,MK7ef|)Dhs'fMu>(TU05"~!X9[-_x3%2eQ|}G[S7M!Z!p[%	a{ 	K(ckzL-H[A?}>oZbH`W~	[Qhk=kZU|xosi+6&%ygrmChC(V _y+0]C71ZQ9W>!k%xu{Ba=_/htq8uTx{^@=A*ASyq$S/	nWc{@s&	1stU%F6"{$5oS8|3	0|n;ONBr)cAQC/-9sqi<w*F#eeip@]VN+%~J8"M$5iqg1L,)u8Itr0z:gaR]!Mxx&d,0.&T
*H=7%Cl;'A9Xp-.RYH@K9E-8x@ x4C!g\&/};0\
37ZO?lcFs[?hGZXM?C?]v
J>[V)c&+E`KUM#-}-P+i>	vQ$!8JVC_h;wqU#@[QAY;0r+KKt'j(}"84>C9;[+.N	#7vE?1lcSD}}U7RrJ|3^t> iVusVM8:mQ\Q&@eff:{-m5~lZ}H3EOi6sS&sM05Ot_4%wY@RUdUk)5"j	.oU>M}Ivmu@%xabdD%P*mtEy.%pjbBgm7j7KtkbwRk40e(1>H*-&tdASo5tD
"L@K.4Y_4=zs$sK%n_$J`NmY
13Q~ $3L%/|*T|*xU4c1U8G<VIu3qt1g\[~fc3!-rI]b7UDV2?E1wBg_z@S03%<^)VM=Xs%+Ul^#!7GBE>}H['})\ciQt,/xWg=9{c 0`HL	ch/y&!'M=
n8|K1A
w>B>yoF\P!dg-s?g%!)0fq6S?)u9C7t#9"DtR.wX%??;?\eIq'aC+kR
s&*t8gWgu$0d0jirN5wO9-gWM,Pv
kX!yVjFglr$C0IHRaLh[DCx<(E.[]!"I:J$KkrtFO9"JW?<bRfQG2v4k_$xBE!YU#2lT:3N$=N0%1f%j^_BXjX>c88!:}Ynd>U-ljmU/Y#,IMK:}:U%kb*0$_/hf4w'ahNm5Yl`H2J-ejkMFHTM<5LGx]VoBTG?aiew)aafjwa;&ly:_m*VMWL0ql`H3XYoI<-$C2Fu,:rh5u|=w,lf_O4LhVCub.b;l |l}m*d+8n"5BAjHa9S`.!`S *AXFv& 9jo/p~]/*off4P$+qifQtFPyILK%u&htA	AX=sW#kR:b^)b|+0onMiGT:yhP<vs&;|("kxAn/xO^m]UF3x;y\(,rIum8)SR@bC
{
tP=}	-l!~:QoB3W_-vbX:/G+7_yzb{]i'[ 3MLCx+sALf3#:Qr/)C0bn^n(l'~i j0qe.@3VVcQ657	-))1S!g&=XB8Ez_C*sd4g:3qewVOujM-`&AVO6&iu:YgFAJ2-*!-3O>TVh'0^ M"1-GqLDe	2CUq?x5L5#{D+h(rxoPq~Bzzz!N'tr~?(,^Fd=_Q=Nw;@M{(y) :{@c`M{6LZZX!i;aO#FnQ)"=aq{wA_8e%(64)0s&'!4sej`6/)ND:h@{xLu/4%pSctfUR,7Az<ZHvo\YD0f;.8"D#@|Jp:X/uQ^odwy%EWFo|8@xa|4Mae(QIvu$@dMFi)OU9s&7C582w*X?,QW&Z9"D$t.W~Hk=/bKM#+-^+GXd)6GDiX8a&%Jb..$5NhJY3r}QG.c`bJ+*`IGM14vzqi|)D3UOB{RI=
}op1Qv+:3P Cv,5:}a[&dhbs0k6/J\0i8fSr_NtuYJjc8]bIZFp4nQLVj|EdoYAct6fJAAYxC`}:}\FPuyQoL	OQ46_qMtb7c8u/@Ahaa:6S UX9d.?@k:>n1^)L=rLv	N0yD=p?3P{(o?Kqa46lnln_u@M$}p\((M%NHI=3Fr4<6a^7)gz*~rW]Au_eQL@+63j	e$PdrG?Q0d!Sfx9e\cAecee6-bGy- 7foSld~Vxjz0PwIFi#%Ou^Y.
Uc}x2#Kh$.GnB:]}Z
 zv,&$FQQ3UDtPfC[2LF&;E|,mIttjqqwzP9Vy^"t}ROW*.NgPdX4xU~i-yv,jQ'=qm$UCluXo	@t0PAkkxHM(ywnQ|.LO)36|8[jex:]OEh	>mP5YW,|Mim`Qgts1z4+*Qe#;1`d$E-64CN>V<u"9=	Ku~]nR6a3p?W*42x35@E1:Zl?;)<!Ra~CcHcGO9f@N?L.$aBHYK
U
6TxeBK&SxaxSl6^	1q9E|4]g@mX?aE+AevsY&HTB,V!axQDhE5vPuSY|i:z}SU4drelc-Fo{e.w{&o$}N_pmJ@`%JZakH_(\6fh:DE',hnD9ZFE:mDX2W8#K5eL:,F(e4TOPv(q;s{}:O0/<D|v02.c&+6?
P5K)!r!y"^/4Xk5ye!t$-*B|G29M5_>pCNu-q3aJESM[F9LspF5U;Z..*q#'BuO`AuW,}8,Of-@)[tSG(ztX.|W@*yz74HuzI=IF^|y]1gG]=<&%-)/6~JbX?o(5LXLrYj<)C#~4[Yb#fp6(9SOm6gn}AA-G727Rq}QR#rWbZVQ$X\kI#aTJ huf3'l@V?<mp~<Vb7H#@X)_*l29g'}@pZQ+O}';@N-lbM=y|kE&{fr6S#=hFZ}H!/.X1$iCK>4@"q<*NARmWfbl
_E	>sb}!l/ae*X'0+"4&Kb7Cw(?QRo9"pU
x:m4U<yVdmV=BCM**lnljvG,{ vo,>{M0|OzKH/rqwP=='O*'s#!t3G\e:z"\NC4iZ7D"zx#-XFNH-owz%sTpTn#F&]dl'%CLN5%R!x<=Q'}d}tDfsA7FO=AeBJgD-'MInP0Sf3Jf%iq51q&2I,0:;?")b1Ct.z2n:Pj{.%}\ihPaC43IB6KV30lSTNP[?%MdUxkwH_-Xu9e3vt[~`:K"U\;0PK&?COWlNWWVj5*ny8y<9r2`6t" f vy;KEmM"[1dAkJWGn5LtSWOwybVtRd\_Mc!m]v	@;F^2F1/=,iclv&%f}eI2]./$,pVu	[xa%5!)Se=eDX<GuquxRT5yzIR7%lMRyWY}x{JjX|uz`Hq(,TQ%Ew0f'ak]`RJ"NMnzyz?RNo+K1_.|l79Jh`!oiww\6s{S|{l.7L<|>tLu{X
khwLOE*;},f
n<\
%UqK^q_GYQLg%XMB%	`Ra2&jbP<*K-VYc}P'6i(RnmO?{)1Eo_^}dGEY`IET=E)7}*RD$Jitq@(f9@q];dL\(a|$a(7Tvxq6a}[~N ]s_*Qi>&YpLwsu0pU[41
#!^!bh ql{u__@on;OSet"&I*P"]RM8z_S~:Bx=UI<ORr2mW$+pFVHy0]+N"G
~#8.mGD-e.IUF8f g^Qe&3X6Sqk{)$bd3=et3HvJFf1lx:nUbPbx\|k\ckj$Kb/=iV"~oI.p(%F*fYPjRw@rz.{ig0ltvq7U;83qZ+zPh%1Hu0B['l<bpH)*;s&d#Ye6={]tT}Z&*_f
j\+E}0KVZzq]]*/lT2]?=ZeM1A@b>E4gjsM@9K<yTX&j"$!$zV'0"Gw>Z>
U-P.9{7u_A=O5-&A[jBJ*Ol'XjhS5r'B6%zyVmxw$2W d|\nWq`Im]?26$E2sY?XR~-_:b3rui7k0DD4>gta#v?;e\M%xTq8YKokjX#ov:C/DwyI]:ve"8yb 7,B#Uq!gL?W>Fw@<p[4x#lHD~ OC&W@!eInX(}"n_&salI1I8I|<&;F#f_$8X{OrW%)0f1LNlR&_$q2^Y_L7a_8FzMdy)ula$'@x\AVPeB0\M7IUSP/GJTT+e[Bz
r,:I_89"KC?ba/;s mv?Y9L7 40\2H76Lrr;!`H^BZ7[]:;hh3kj;7Zs^(2g<;:5N9TKn]uVk;M3-[DNLeO/Ca&f|60Q)~es/&786?%Hi[-,~"D'Alw?_WSE@r?3SEfo(<36QK^{_adsg['Q48SG5dt{*AK4#*U:c4"?w) -)%$6F-TF-78qF/3%n${J	Ht;z)!/s5m0k]8	2leKQ:4kGFJed9vEVi&R+=fw;$PBnN[QHI5=BlbPNN(\arEB',;o!p&uCJg17tzhVu2Y^d~ ?V-}[*B!:o\ZkP\$g27'eahccyJO< |(~@_Nyn%8J+2sOgPtwCt@]m!$Tz`yLNr|}DTc2x0qIK	haE@BPrDQD#&e>3(Xg~.|G{1*()>I`\'e xg4u$O;eYa+E_q};h=;4!/yT8k(
m98oKAV{d`f%Y;*.r^MBq{TZ(@]YjO>O,q+\^\7I-%>[aO769Gb3;-9p@Pv1f~YN\u?5Q~p"gXx{RO/^KBqk Ib1;V'I^]"iW#N!*P)zSm6F^n#=[O.?Mj#1'meoZ<Du$uw\jP&TXA7+ZnH\}1}kdQar	iY<5qyLhz5H__Zv\GMez=D/\hGx(ft)bl/C/D\# /eO2YC)q."F9bB/ym=.g<%V;/Ezh*SLVGpcX0aI!R>d1iJzNHPn>S\3(9|M3M%rBp\B8L+yag:Nb/bH9Aa"8DBsPwALvo`J\uULvnNmD'n7g%sURl,lJ@"9`pY>VV<e^p|^T=m,=>L'|%R\v"{o2?N0+R86f,AnZf+*m6dRg	SY?,. A}~f,auE/Hj,kJ-C>`X]anc/J8p]D<3>I6E+S)Jjc;C@M$"h&ksZ%6Zbtb4:KZR@-kOyGf!Z`@@l3Ta?Iv@Wl-
Ky>s*_kd}EMtXz~<wfi{rw\32A,C)"}cBsoF)cnr1si}/_ 6:(KU8-%[zZM_/Krg(qT@0os!!tK+v`%;6R[VTbhD_=[g@)Wt8CnVgjz"6o"q.l4umk_}s>Pfr3BF(fvSeP.F+au=oK-k`h0*]6._>8D!;fgk/2#O--GeMfuMk'oS$O=)8[-u)`	tfNpw.-:jzIWe^@{|xh@<:FS`F?dTxa&r+GwB}kA	E//	KL.e2KY(y*zR2I)(	-`R-vzJ)\|2z{8?z-50BO5?v9H]?0,Dqd.o22XAy{'9lvT]=d(C%K0_B<fgDA92C7!NAw[<JL-3l](+sEj:	9`$Km9Wbv;a{4G)wi#BL.G _BeAS`[sDIi.Wkx "q'>5z3YASlS';/Tk^Q+k]g6n(}68qQ^K^[U*]kre\=S~#zpR^tXOWr4*x<UL.M/J>LwyqT%C`A	mdAE$V{&.X]bB)y Q}z#=sajkcKd];$"!ZUhD'/P:Qs\-cnk*E3aAgIp9=xRNZ]<f1V-}bdGg'vl+)rk!gjIvnZt{ates"@RN%94iHkF@3!}-,7gG!gN|A>;lvF	7p E}Lb/VE$ETmK|Pa:fC8FNb	|h'J[$0%)%K~Vc>C~:8BwihJD3wd5O$ob!^ O4]>j&X>[
9i](fmZh:<!4@ E
="*VN,R+]*BAP`~)rb7-)0`T2$>ji)uuRtJ\?*:K^ d`\J<0Gw!&EAnqMp\oxR<(.=Fr,2-mD}7\_f5D93/Rsd ;C).3*G0eRco~
d>0#">2fiGE:<1$-0<):<S8ao8BMG`	4U;x	+'
`Qoq@+U=a2Oxh]bPgYLu;$Q>9K|gR33f]ar`FN)Vpw.2	%[K,JcRna{f($JZ)%KG>,`a[Q|"P%*u.	yj'h2@4s-;67A	"d+`xnaAmSC(uomI_2]vst-omWT<j6eTwhT_><JEV.t}v]:;8xMGR*itV2Y8H>0]wQB&5A+u?IW9>//ga!F19i9KJw%U
+V*48#^tJL6k-]7gq~?QsMdcp$&A3p|vjD'mXR*dP wGW}jCf[2zdEyWb	`*1jI2dwVSXYu
q0z>yX
'M5n123\
"%+6\5eEPHxL/953YapCtFj])8Bmm!BazXdf!kX9k'~;cfMO>:#4rMzzn8K):0l=|	R/Zau^decv:R[#(,hd~X0li<29"F6_HJw{:W<.Mf0:#4RaXyv2?u99jKj_k2%83h#e{9nxy~|oj2b|IiSo1%OARA;z
.olD
"W>SLx@v5_%6Bnmh40O@U:+vm|i+1qRlSPEyYfyumF{U"( @J%|H}(+\NP`{X Gzh3>r3tv41L	MclhS)k:B`:{po&mcK_y5@O7?Wnl=y%]3/}.u8\K:O):9b8oCS:Y0U0~\}K,TL>/|cQWS	Et:OEI|YA&Z#{:7)e_:K$Sg%'<zH~j
<;gPiL]pKLA`LA2D.N+[31E'Y-m;NpeG$$8vOIcx$1m^X8tc<ir-"e!$ 8Z0{Ei8qQC.4XE_6*1>SC'zMJ"Q0:/g4L]}ltWfp,CQl=(~J,E01:.4S'=zKzt9XRhfJL37}'C1}aY~Mm/6LTwd@k*N6r[Im+ZH_tkt,Kk4`zp&<ZrWr%ZtWx5:`kk_8F'(o%jS$xx|8j9$_0&t'|Jr9L9cg 7b/&[+%_#$:	=y
85bQxWaURvs^_V1;qvh!D%*S$FE%Ki[8>rL]5yWjA##\ippVm6C8p,U|IRI\-k}f$bLx8*=iwn2LE'C:HE6IQ;~JM_DG/rNhQBVUnfzFqLZ2LjO
:SeNm |9?#-)ajRC?J5hfNTs!Dx~-rl+v" z2XZd1`""kdpC/xmlsk\8AjS`92t$Deh7Hr.q<Y*iO.8BgkL
<g3a	/)&!(DJwrSC!QMfBSx5Ce	7\ud)PC+0g(l#r<0zAY=d%xhlu[:U^Q:bPs<U bC>ypw+D
o3=9iCHE6i2qUG}A~~J0!fL(	MW|!U+"&Nm<*p$&EL=`2iA1|U{tBRVm1,ET^Iv-D%N@RqMX\zsVec0!sEWf!?>!iWg']@|A5QM;v%$_sL
=0e2F,vM]"5l/U*3"n-2gT{C54J*~0DaQF(;8k#Cl{<&Tmx6%14:t{( )cNN!;6;f]_mT3 S7/vuz^J5'%z%~AxTX@/:!8|sI}TFF1N\"V;T~^:Wuy&[xATB	)W(6/>&ov2RE^NS6I&_<-6KeV-U3w{!z}#`j)Da_utbuB=/IEA4'gFC+J`PKiBvP"7_RHLI8RDI9Y~PH3$8c=^O|i%G_V	Sh3ca7GL_%poC~F,FgJ}?Qa?Un1~<@e78DcI?D
Dj"(}?P^;}@o~&:b,N];.7	pmgdL{F:wU
&a"KjutpyE3@i#qaQmV;7~iAKTp'}8UD2x+@j|&<R<LWH<lh;$Q7t	%$a@@g+SD9W
Cd&:	bEc\y //HD&4\4|SG7WUm=LZF h!tO``]b-{k*{_lTYEn[:?~h}&*>9B>b^+8A}/p].HjeaA"b	X@Rv5raKB
OzSoo%!G"<\h	/<9.a@>PIC;=!Z5a?YcopxOD:	t|("qy./g>p_pvYs2WoU-n$sXj2Z|%QrZlk[u^I.^ .MJ x9W47C>g\`1IlSW	&ltr(yfP-;` J38x8KHq-FB><I%%xKN~B$(! cr?=QDl0-R9:8OJN:zjmX+Y?pmvp&aU*E<jYkvu<}H]'u>9)u@0!x&pHG$f'|b(p
{j|g^z4XLgIWFN2
9%K[m2I,	h5ky,M\[8X@3`U(-8|DJ;9L4L))?_`|>KKwf+IDbmr.W,P gU8T#F8+9wwV5O/Lct~	1]h w[Z@|zUh#0E4Py36-i[wPH l7*^Z
#A)Il4AFih.Bb~\jlYRH;NxJ3]oUUkU2m1XPg{hzE'|T'ROWNis+)=D%FdNtgz_.B6C#]B;g/v:C96JHQ.i*d<ypZ&l8=&C#8"y*T&5lu=xXUpF3lb}r;Fs!p3p$gLIBD]4g-n~h*<Zl/(_`LuyOb`[>fz/]c$ca[iT&\BfuxKPYF?Tg4<.?H"4|RwP:h9~xttbsDTF		ZnS;s}mPleL4kweH0k@zC2(UvDqxT'>C8w*zw	K,hokbJDp`zBoP]1xi{LHk|cXq[Tshmq;Egjp/cHD!k5ow/<2`2q3R;!`P'7A;@/y,nga-b+,|oy!.^i|#0wvR/q[znO)IN 
C&!8jC^-=<dFgyfl4%9:fc>%qHhHpZy|o.mm6GnEs{0b-|&\d}nm.6RnW7n0j;[S R
k`8wUJnK:[hZSJ"xRf[nk+'71
?uqKt8?\vZp72G"l/LxwN0soz!=YxGX;wFKPOQ*Z#E_dKZNsM<IMua:{	$E{-TS-wm}p!Ia#0lTtQQ#%(5bW%SQW	A|8dFQ
YIJZq,d	
6)N8.t1WyP -4)jc]PZ qlJ!@6
ry,hyzG-z6%OvB(hd&13Z>fP_6wSv7uSyA(HW{<7>E;4!x.:a5-(xzVT<VRLfEW:T`GysNidCV8\(Umqtf@[6ZCc[4Ek<npY~GLTC"s*U1H(!DAk-Mlyu'7C5$X~c\N}:mr+L	u,.0?xs0:Yg14b~tn]z;(
Igox	9qZOP3Hm}E4P7ij
.iK;C;lI&YT#U$>Q.^2HPlo!zW7Dw5(wyy 	|Sgga1Ic?%791:FN9G!zyRi[MSu}NGFzQqzEO	i0|d^f29*sD^0<rM|-@v;OV&\g*'L=fCa!pu5otr8w(AD{KS3T7\zkQPI,n.7=1DHOCfm"`p8j= !:en1F8pn [EPpmVu"`+:3POtdRNTm9
(B[(bK"3lASNKJo~^;g36'HFu7%1b.Zzj5/.KcA$ARQ+wr/JO{7oP&\m{;rs[x0VT]lz+yW'J%*
lWgnoZ|SX	(P_<'T{C%*eDj|A}Gdu^QxR3<Eyl?dz
s	<4=dLnRqif		OHZ6TN^JB(g_U4h;|V(K!3[0;:L):*n+^0#4ElT"HbAH(R$hf ]l)?Ygp!] si3xF3D4<ft3t	VN`x4D:VL&xl`36Kw^~M=62x*._$4Y-u3LH)-"}17)_d
707lIMyFq$H}?3r7.o^u`]N*9&+Y}W>nkm8_\w	f]{=JW(X?CXKW0bfQ%C?+xNIGN(fQ;uW]{IdmJ*_])d0{9G	M_d3uZT2F.`(xng@0SGgS(f	;W
=,9-gZ"TD>o;}.)(do~JwjLVG"Mv|-fD
9iqJXrS'os:T?PrN85G$zY+_>WBr;*dm@oa*63<=Pet*
ntel6hSDv':%cPOgRRl-^zR1J0{@?{sbQ?Gp~U>v4d}!1-&.VP2*0jjqNt&dXZ\|ziJ2[;t$O2}T7Wr'6GxCm{\R{4<I0%l[520HB5m_(KK K|5sF+r01 98xu;>PGhVg1x78n3R[-mbh&kJ_9CGliJ(4q&#Awj`U\IxPs]+I[$=0Q^S|BSwOW0-7974:V+su B_3#bfIk?R q4t6E4$GT+#]V]$/fZE<;U-4lV+G>E[tWqws?5|YKFp=b?j6jbCfpp#3<#5rjx^	a
Co1AEgJN6OWjbM2mXvu>v`%\xy==|kno";]I>(AZ<D%nPmD.+o{TmSwO\nQ0KhDaYZ,#xLw&:}4,LMVQsU)Z`bDkipF)HoH[W2YD0*F3N?jlUM{~{1("FNvZHb1WzQwBN|KRK}KtJYZO+z'-B&^1mCn({_ vVk`?@9=gNA
Pb7{	Dr`j]Ic%xc|QbYHNymuC8On#	%22RFZ6ysP75`hD?$EBjL!lh3P2	.n!Og;w24A
`%'1Ju!i
eW'zw?q)wDo{
&dFRDjC%)xr0)@*q('.Zo=Y 0*U0e*L>+vSm5%yaj^+$((V9a9Ps%QNszk \*fpw}5w1*)_lQr)@n [Jg,MCm`2V z8I;tT.]c7hH^$hh,HZrLL~;-S$c^@N4Qnkgl
sZvXUhPA<6UVWzn]F>	ou:P)#=`TIVT:R1Z!63e>1	&dh9\8Vk(4` [CR[+F*{@>^}D&B7m_s-CD(+E}2	&@Pa?\%j{wW$~Ur]uyXVSsD<I@Hb9`8<@2_o|w]4MU53lh>5Q$am}tE0JQd+N0RjnqE1wKe
-w<wHog%Yfa{5\VM]L%<\5|<&!\Ew<>V1.t46tB!wH5O7/$Q&Z7,,"bDeibQ^.I=U&#}eR28d'sRs"H;+PzUM:MFgnIjel3YpJ*GljqIP8EK-KYkQxu#d"nM@)I_q[	uSFJ"5pY5rtG|-cKjcH<7n=,EwaqZ.uA4q2[y7G\%np-BBPE*S[AFuw/TUbbi-f[K2xXeQ=8Tl	gJQ1p|#<MmIG;uA4f"D%=5$05!S]F
=0YS,(@Zk%h?8N5$R))Z],yQB_YcZ|,8zu$=4z5z]:p\Le2ev\Na}'2+pmOom5<y!EFA+uP3lF5Q}rZb{585nB`fF"v	a/@`ht`AAh0:Xh*A]e|V>+cy!U50>n=p9fz>M7_vF(?Fp}:~2t5x== E`u`'L2paCdK.~dVwO{7w,FJF}z?(.W.]ZR@"&4fZ}C'S)G3~q
ClMD+a&<NDWMdNP{lS{%VSkRe!:?L!u~TcV4~t!mtW2b'H<X=VyHQNuM1FkRTRYkzMi<*\!Dk8pDq&V"DXAfHq&>lHXqt'Ce:>JpA "QV>*pUAl@Riatm<Cm,\}p{s6aO|i
;ewB'|k!_7l+6t{+VVA*|{q\w}[0>{bVAnOTiK_n0"5*xn__	:[f'\VpX$=QZ(rz)=}T$JmihBp}c`!2v?x&1JLk1R|jn@xyG+oZ1F!e[DQ58ub-T,qA\L<%'wtWt/rg|DF4yWJZ/d9V:fU.5lD1yMCO^ht@C#?-YU<fnxX$1/ph<n"M	|SvsD_GzuRXcN9
J%o-iMh(*qp!,XQpj*[/o!\_`-g*8k8Egu^{c
1-'*.,[!a-nxq^hpA@Z'p1~j-6Ttvv]_0uR*t1:kDD&AF^'.@@s:\	TatkcWEf{(G,=@y:);R{>lye!wK}a&HI7cUzf{B$}{3>,dQ|^vps(S&jJV=BF'Cf!,Du1_qem>-rB+}0:#R)E-
,X]Q.^*Ym9>vWFR5/$e9w6^^p\cvg445)Y(Xy@9GC?+Z]bbQvs(M_Pl&U7*oGOXOL1	Al@3P}8gyd)Z[FgK}tVf3"Kv	qDRX	-Yz}oK,!El5STo"DcO(P<	~ay|"O9w(= n9H@.G`?:AjR1OCGHl9-{e<2-`4Qe._@
tlPl`5^O\ #E1;:5+%2(f}t,NO	kFo8u0Su$Y{'=!d?s6USxkRQSA5;}7NkgtGr3s2uk2"@=l&_;y? ^AEk#	x7-k><}::l- F|.:S=88y:x9(WU]b6'fgvQPv86P+B-yI?dR}%Ma>Hj'LHw&z1KxLrOv_|L2OvI-2c_wI5YY;r:,`CGu<X7@F_K'x<J<SiQwE+$'i,w9%TH;/
14i!hjw[RpfBZ8m%qo$J]Y$=m3bjfl Ab,34C`6?$Aymn(cf6dg/|gxrh{S)^rkF?ll|f}E}X{Jig6Aj^'owj,{=l$gG]hw{<@kEm=(|=P^rHmSl^ey>YP>4Xkiw-YOf\s}4Ls.(vmC>GPds}Y\<g8Oj4HvaXp)#2(K(P51!l~t}:mN!"RL$fHxCc4mSjT#!).B!,5	1aI}y75ka]J'_Y~R%&&MsW^@*G-s>)@0W7Pk~g'*^^7m#a,^CSr&5Vbfc=V9xk.Kik"L)xe7_K*p	G\j`[Wp`vC-osg^M[,?!{)IZE$SK8x	X^.Um|%##;>_W`TkJM/:V?} X+EFGR$@t^$VSo6	]r
SC`	~moQC'ZQIM"ri:Zr4b$?{^
o1D=`L_3hG7'@+2!:R+WU@402qS#Ee eU^TW5n'gWufO\u>CJADqz`9&[]SD#8wDH`cJpuJzwR~Mj{^BoY@O:P4E_) !X 8ikEes|[XqHh7%_3SKw4p3&A5HH,/-]tt).V,"g[1'ZL2}=hwhw1?@ <uiO?>m/k,Z56U<ba`ny|h=s3dQO@9\6L:5TX +b975UvOsH2a}gZ
m++=lS,v33IyB[q2*iXhKM6p.`W	kWwEWf e/nQAG5SJrK9_OLh[0.l37XL.>A=$fsw
-J`GE[X
'4)An\3m	C7D'Hd3M]6Fuk2\Gj<Wb&Y|D6(_E`N~x*9trC)@TX1{D?RfVcOIi9t6jshmAZgm`D&iW1RWvo)TL_\6H@OPTSV_hpZQUn%	^;zsM3']#a)/7^L5C@(<fLv\Z+3ObB^B?"Mn,dO`Z<K*O2f\D}VlxPE#7PhLn]EJ]Ulki4/$.>a6+bH
Ua.m,<}%OFA8qx8:8b!Zsm4F<bB'0JVCk~qp,~X5T&"e<:.Z';tS^@(H}<8#{-N(C=T9	O351@j]""s(W)E	y}m~:]tllqarm]@IZQ+.P@?>0as`>q"'mPB)N15M2-0_Uhs*$/\A7C}K'v@K[A?Foj+Z{fT8<Dze=duQ9SW(t,Y\#F<RyHaj]%+;d
-s .,[^QD:E(A;h\uSi<H+7Z*mX$]2gS>JJe|~YAKSLz3Z;^[}-]t\tw%N/2shxLx#X$XMF;d=
]OG8U*16g+VP)Vv=atdN\9Ic#::-vvU0@hW5M~|C-xN,-]6gM
=nT1b013
Udf{44mDzmv^lj#|i~#?6p?w;E0XoDCysA	(	70vd8RZc6^.yG"\TrBh1;Fye+W4,aHM|dS	Ce$dqzc[l+5yXQ%9$7(*xxPmaEBPycv]V0fK||+NF=I{0OQk@yB+o:nAjwUP/!+C6>fz6Hr8M`
4k[PkVj|(lNrM.sOV$z$Xt2.^SYpL+,"%-P:3k}d\jDS>#d\Dldr5Jrm[y5?}n\xW=3`JJ.:(dQ+ZLVI8	D"QQ!1;%puJ`w6R{Mg(MuaIq!ein|Xs@gi"
kO)]+)wYz#-`,%(@l-NolYn1u/_W\AZ$]2VV`D[:-;9?pPkR'vvr,i>UkD5n-VH8zCO*EI#@U<sBJ6SrJCPkH'g2j.+R$,`$5~)6B)WX/:uXXy6 >#$>.vlayF:%9:?Gy9S'O\x<"0B&v2T7sSA#4tu;a<=-t$"me88{jy`O5~"{kpOh	icrA*n9Y//UKfq4@)ou%LS%e@QX@'<EggJH[kzKKas#gA+#QM)WBiUoP91O2ltdx7~cGn=[T!+]_k3-,sQ$to@q|EAmtQ-Jawtb*D(ltoIGaI6+js<C
Ns8[?5bvPHh{Wt,'s tn-#FtC'0]ovkwe8,fJx8T67	e)-69q=+}H5dW,BtzIqy*9
O[XE
t1rB@:kiYz&kj0">Vjr7x<	j'1*HuGiFX4+)9hp6.55w-O.Tk6v3mXHwnE<T69oYdK_S,{?g*7:[T-BZ>^bZsbuML6/o}g~57~RbO+);FPVV-dqSO'qz3\d<BNV3&SJhv$G7RRT;P'|<]("THbla[p
YwN@hFuR\z:dI.jFD{MM	KARu>Z1q>P#Ek3[4}totz:8WSfkS]jI>V8'XP5T+doZGJB]H-i#r.L<@b9+PExu<Y4hXSD*eq!{OQ]+[5wB=mH}JqU\HG.V5W+@3}\%Mt>*G`k`DwFN\Ey^AnMNZbaJ-p#U}\iIW(\+cy[e$[\i/xOTMmh2i:!e!)h
/#ds~K&([)G2`=Ty1	my	jOF`j_`atS_Lp)`)KPu2ZY,GZTIY0GMJDhC@{'lEE]/N3j"$amMA3.
#,DU-('hjY&pz*G}
D!rY
)]\IWe??Z$HBkfV^'C1*?Zar miALb!i}GySCMh"\"hi2.I9i9KLqz?S	L2p_eiMt=|mxoZF%5*CW}}w@<|ns-3\A514N&eqJ6BMfZK8H!yz?w`'42LGh,fK'fG@)\wb3!l2=@22ptK
>[`"IkX-vhYBeR3M.XW2x\wI
*=~ZvR3};>h
asb^`Pr=Cb%#fw0!u]	0}wi%Z5iHEXdaHlk}~?4@ir#gd:kM)er( [A*O;5G2%365~g}UL+c7ds)Zw]G\w Z9Qf{ ":kimJ 9QN#\$h%8[KI"J6bZX3A[gJ)!!<N'gh rKg"=g>%!mxKMf;J>12
Cn[nqJt%O9/j_FO.udJ[Q~ml7[6N(b+IkY|!Ci#qe/lTIJZR
yt)@u	Tu+DILM&<
},5Ha]/6k+m?l9qA9#'JaB8E
93;Rp;c Hz<CR1bvbQU
zXT2+eAb:0^$6)/Aq3]5_VS	fqn!H];=9{T*EzIzr^HZ>]JRAu8A(~"cftUyLsCHqB}Lf9JJo6?nz7"@h}"?PNeu%j8m[/q4zEOr=CB'`)VD<HlIIU57FvAw;ODU]@(Z?@5<w?nO1ZsE\Arr>'UxtOmh|\(4GbXlKb"{@dfJ`c
(4wmoAEk6_klLQsK/JUlZ7uP~a9JbQGU\H:*|1.b*cL5N~mESL%fU3<6ifV8ew]#Z7a ,$R3[DRGZ2UG[WD3JEQiJ_Q24Jxh,f}H!4,{H#Ib!-~Y?=gp`C+(__%~VZi$K)k^Lp\01j\}(p`H)r]if*'&1B#FYHHkv'Fy/R@6JHPVT_:GY7%T^KqB_:TJKSN`%#R,6M1<^!>y/wf7G0i.k#iXFx9M3Oy-Q:{$kA$"jk,AgQY4SY5b0!'M^b0rjbUE/hh`Y)PRR`km>!4#s(nUyb`4R).N0?aS74Rw.W9*n{|z3E,6kAboj[hWIY&&m~2U{*R>eWa?'j K#UH)NGL-\UJ3a /o5oG!S;t*/2$0YTZ3V)qA88 3#:BXWDcW~G*ppsH\%!7-]"g@=GiL94PTB#_<'Zyq5p~ 4,BK-C T)<3g{7<4f{?D@%uPql."Q"!HJ:M_?uWFyx
HLM\9"]I(|8"Z4{^[QJvsxega|u1)5B
68>kT*t}[b Ul-]k/-7#GDkLl7G-,[Y3Cd|<D`Vl+d[! _@Q!:;=#':jTuZh]GYW\|Ez0aTV1so^h&ZXu&bP{2( ]"fVoL/,[a(x&z	ZR1C5+H}|+x5yfR-^juIBUC*|_t:	E7O0<&3U_a9BH	ni]>DQYrv.sAd7iEW|?@@J*,tW{|}^ykk}3`
c-/ Sk$12;v$6<=+<eP]yC7vmyzl7?u/e)\5*IOn!irIP/\X'zcF-qFWJ!|YF}$TxEO30e:\!F8LSYXqST+cEV@,Vjz5O_+r^}M9bD7\86B%>Ynpstb#O@W"?U|62Fyn_G"YYb;LtWRV?/~]-3<Tp1L'!oGLo!"ZTt)9Z#=T]dusnUg#<:yCl8%i>PP5!0blf=6 [<vnJ^ M\`W[#b|4;%305Q)$OY~Q-lB3b|nC q=,
H"Dk7W4j4>Zele<UTIjSaF,c!UGj.@R(6U$"<'SsGiQ2B&L>!}OZz:0uZU$R'E!yf25:#?Lh)OZjVYPuEB~MKRFUxU*&t9	bDskGnIY]a].tB>~QN+:D;H=$J|z$? /|f&fnkF@,x!;h#dVVShH"ZuN;/^PZKUGzVL<L:36v=|!B)w4)2AQE):
+EmIlNGjj0ssxr?^:`!6:cj_pHRxPPlX8PiZV6py[Om:yWNhtl#6nU;.o%'OodKGB;j
BW1 Wdz-}~bN1tY`\[itH0X.]W	^y1	B3$B,#il=lNn
y%scW,B^-FLrD]{=:neZl!egd':p_$.Mw$*e3N*4Zs`BAQ
LuAg
8U7D?&28(HhfJf9^.#(Ci(,%!P8PLXbde	ElM}WLvzy]hqsL >L#/ w+9~.^_4 x)yHi+}S+p&lP<^Tc~zuv`@F76"R$+H	}P9/	P:B$+]fPT|2=hsFn/
_|M:Al'\	6H<bCeVySh3XGw)$CX3?sCjW@_xE=3GCF%giJ6w<6\-cT]c=>~u
zuk:ey{+4t>f.{@Ay}FvglFnT}_GuT\ww~}ZU-n34>zl0eq!I cH