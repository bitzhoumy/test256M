thI.`##U|z(U+?_B'A5z_!Tu+`k
 2Bk;+GJ	&33/x'jnO>gBdaq"lZ<)%3[guOe2vKBXS^dkO6i6e>w 1rt]q12gqH5Q)oC	-yc	=`;4hK%qbBN}*-RA=MEGJkETR?q;21{r{+Hk.0-hGGl7ZmPl#A}Fu&p9$8z_nM].hm&$^!I10E;5CC:}{SW]rrLiH)x53G)f87~(y0.Jn+MHvJW#	XwSO%]#(6,a9;YplHE]D`nAxdg5 pj)\+U	$
fE>b`+mKGHL~^ 8e\o%x8L]KFEcQk1,i3<L!2L$}2F)ey)s*=0fB=gme|q@[nn[=)4=%92u8lYGIL*U*k<cC1	G|x)}9hRxBK:flr;SW4^b@nbrF8gTaU?||zFz=So=-|oXv3YI='8K10) uot;7"mp_JQ(8jA7WF/|PS5#@*^?vDn=\G
gKh[(zk[Xj({8cO}K#!v+.TJMg*
l`U@ys2D6)L))<ID6XJGo`'g;I"2)YvRo3A7iP@a)eooS-GGx*D`:KKmX@dX*.Xv@Tmrh'-cou5&Gl3r[3C>z|H
Q2a`M
Ka\b,h_bc95Cu{6WGmGg0*o02 RPZE
IHZ[^bYvv;WzjfagleVd'<g*&|jOV)7JR-&E- W=[W6%_<Nj4zwoABOp\'T<A?zhL}-yz:g*0_fl%E	buf*)ie$]E4RQn=D^aTZ{cDl}qV_(814A!	jW
\f)rhW;	-0a^itS5^,Y<:UPQ{#NU$LBgP~^+pf r;oW|Jb@ttqdaW?YSLG6\5ASBtYR,hs/b>4{kkf4Rdt{$3<Q<2Qq*,D^nr'k7O~(Z0'oKqMt2G{KnlK
3rf$ybi|vr,(1`X;7cay'j$QgFh
Mxrb2S}f`T]{5rN+x?;y9ZjzE0]+fNsj|"*TC95r\h6vdC8=&>Qova'sYAt$'mL>R&.*B)%R6w/Q9${YR{F(`xLrysiQN$i6"0{wYpXxQ4]BlfTq_'c:n.eCh?<8$xhLVauq(

uw56,jZvdxImI*+I~d@FVdXJ-Ap,.C8wX]#{gedr'%Y{mD^_h|bR-@*X~"!^!%HSn89HIS44)VM?rg
;GsQ56|K3@#y
6mi,#q"Upl"|2C\$Y,bMI/t7>J:FZu.,IKE>.wgIQtf,.&!w3_arr.<X^UnFUUY	I\b`%1oEC'
+Z7S.! @iU[(kP	Z$):Pn|:iKd3AF12%:nQ.de=NGEHiW1rZ[c'f= d1krzh|<we]#T)~2NOsDbd)S-SSfGGRXs}uz'")f)*o\jreErG6[*7xj	gg<?;QsDXf%`Lf<cOxQu#Izsp+[sX@~Mz&*E_>Gx$eX`ov]-U+I2SW%YYnRhq_\QVX:Hqc?bFi;2q;d#g-Rl4w7h&s*L3DY?yNnb^g8%U+^)eIS5=y!}$^!d(n5X3e7e;)j1!osEh/Ubac+sDfL?	wu3"@[y?Y22k9C=7?bJ.TbQ?7
x"ZC!,MERA3c}dk>eK0JgR.Xvy-Do njL;Y%>4WDVy$k#k
kagHhX~?ojs?'=u^f/itc+qcxqA^=:cwBO^4$L]7b!=dItMM*9Eu-_kOhx^IC"d"`s4yVljE5mL3:i)H_6aa21@WK}IordqTGlt#H#XfXgA%3YX9Du9M3Wzv=9-Ci0-h<p&+q"8lb.7L#1cLdWqC+4;ww[-G'RjbwZzX/?pwFYI1|VTO%!`BsGgti5"aczYyam%PFuP\j}^	sZK8Q@{zH:c9RK\yN,?}$({vb~/-WG
X'8K7NU(MHOd1wa4Y$xgXO4=M?Vr[[n7}vD7NcMUdFaN|P/\+Z_V6N\>,k2k1Mn<CFXDfEMJRt%6.R,oDUKfeyh?pDm.RA@XR"N	|US(jVWzSTT*}KLzC:72]6Wc$koYNl4=iybXI_R)L"`C	TdDo
h2!J3(o="\utWlN?$UgP	xNXUwNFdU}1HM#<b/U0nVxm]\DY(;Ns
<K;B)S|z2vx]rpZ<4c/bH3T'02.;$!N=ete4G/?r:R7u"`1'7pvDMZ"?sh;S1w2Q&t|q<6%4UavQ1/9u|hSD}>{o9rs{>&!9T{Y}~.l6eEQ8]Mm3GriNvgeioM`'=V1
G t|m^F]VW&Gu~8~EDu#&-l9y?#i3,<_/) K_W4;8+r
akg1~y;[\$.X-
zF* vxu=cX6DX:)6*+pBeE0UlB\a8;kA*zaVm3S5"(m*kCtx)A:1]FY"S3EKnFqZEtv\HPO_t?]&*^r.\7ZYd*H(Md(L8*r1i,5P>LT7DSt^IfSX>K(h&!~Rk?](\JQW|WCqPN]!|+_2ikG3+\_>+eYUVPD_-3C2i_|JUnSlXU]cAr_{|p3kaNPVdg!o[q[]CP\nPu`H{4d\?ITiJ7jNj%unp.9%9b,7>/^nU/Fj{D(|XS}Ct`U Ezl>REW:gf\lUH+CiP@Nile7]GVaGs/C-Xi7Hv#seJ]y<%*l6+vVl;$X
yV9*Q)1HmQb,L-3rry1SJ7sWachs\=@t>48nlq&lwfCEMbYe_[Ra2V[%o^[-mymvET9wVY$kk"N@&zm,#4f/C6$38+)220 >5wtkdMxfy.\)_Rv2V2^4?"^[fCy.z_pR&_Y`OHl:YD0lw:M>LFPS\>Rcth=dQAB9G3&e\B)lw*202f/4$~+g*B
%)/v86+&Pf_mHo[whUw 	&(<w%if@oEKF"z96(6Y/fN5f_s[YkU.8E#O}t%=9SUg!O:3k4IRZ=k_K{El-x
P#L_Ss]vM__!kWJjS<LMqc4|T`4{C|f(X0@_\Qj]cxgeZzMxLA9|.Vm&C25=Q.fBn ^$F9e	upU<Am>$+J62y3!SZr)0G=P8[,mRP1$!ThMIggPU<g)%rx>K2v2Y;ljQ]`+HirI jLsy>N0L^!FVn"g#zfT{32G9w*UmjheNf5]:k<m?(J!"69$:L_}Iqm{a`dpnaI"y<QP7D ^6c(VhK2(-[2)T	i'{?y_Eo(T)gP2ngT>')TbCf{H*_;*'9C$_"5I"*:Y4T1hHQZwUEAwZn&]kY5QPf[i,5.}!]{:+CofMfEjfaN`C\A!WLNO;}UP=D>@*L.ByR-5hK/URnM:+m_^R	^L+l/R*s}]:Ro:f%eJR\i1m"pTG>9#-XW.It'!g)h:m3=X7CfQ<VZV2`0TsNtt]0$\+*oYCo,NS\5Qw@p=n-09|^vn=+wg;ybN`PH>nu(C8$/&gRfE~<	xas8'+aIvL,oLl+v8@[4by$blfi;wvFOf%?0l6KSta&8	m?0N9'!'`f3FTEH*[e4z7|0s\@C)'DlzRa~jgKa<J(D#my];;M<bzFn4.+d|l"w64jsjVk&O-3;!WPaP~2aM,P>uw;u"C.7qy`jdzx9sPgaFdR4oB~s@2}C]&naS]2P/0c]"1T{W7fa
B2m=4BW_Dzmp.Lb$4{Gc2mTy4NQzEBitlGkS[Qr X?w6|h<E@bUN9vHPyg -glkQ	LupG31aSwK?i~hPr`fdfpl%u"6q`JePxQ^Pn^3
/vT)4EYW&cA^;q.HI9nO9
5 hs\hQnT1ddALkf:[o='Tx4^}Ib}0i'DQ,tWm7KF$!Q_XvqJ(`~m>kBmZy>;0zWP|=P0Y\".,vF& 1xLQShF
@BXR^h)kw.NWuu4(=_&L	/o&)j{XJP"xW.:D5UD**^i}5_n*^r}s NOt4G|oWDo5t
!unGC@9[,Xtjlk:(HJTiI@P`r6u-9v%9%"ts~M%^|VI:JsI8)oYUD
m?eMP*QI'G7TNy[5Ii2(E2ZtYa`TskmeJTVu7LH~7s2rWc4GdZ7kdCd6cJF^g:b%O
WG\>TDZjW~^bSyYDu\8PBrx2iAT f3oB:$w([(Aq2}J%25~bWL_Lk52gmi6 WVKZQw8%).\UqOV|:B@`.ke>VRz<ds-@H`
X_O22t]eGF:Uext,6s*4Zz`!QmUZ[	.8WGV{
P[PStRQr3tsu1nD!'sT<(x,u?Z\Ooa$.F0Vx\-[})*9u~\qvp'=9_rd%fjV~+za

}S;=X=UIm[,s{1{n'= 	];!+skd(y3b[#"PHK7DOFs?Ec=YnpJ8O]\K8/9xd-v}"qKSO_Zkq;KYTk)uj_<e
E^B&I!B~cd{ry<+D:)3&;@SJ)/t~p8,})Y$a1[3)B0Q8|r,1M^WoeBvNI5e(+6l{(g,4(hG=JC!/u<Ji9	ZT;&
=C3!#md ]z\^`4\G0nMl^'C:Z/w?q+RqTVOq_OODIJx;~!NaEW{3sg0:5[3`g@{2}oO)eOvSY%8/hpQ #l|{[bTnqiQ7aZ z^wzc?l>)i&9O7#yt;Zqj`;-'lrv(TpYV@R{xgeB&J+-|g*W7y\~6S@QCivWxt)-6+Z!mIE,aZP^8`[RO		[/7D.B2o+H^JZT`?TZa6wk(Qr.Uc_&4;EK9l_g&my5mcnqzf;c8Y6h9;m6^XM@=o090RsOzusAXN`\CEGrj4z`n5QJ3cbqG[Y\;t<^"8U(UUbV{R|{u6Y|c3o-F;N?1GXR=7F`?C[T,8Jhs+{\k$O}lA<cyXtjo?o2GOJ(|?m\2__,W+j>1'HQY~*X:Tx"U>hhE51GSvQ[49hHuWA 
F|AB}D._+Gia*^_`9%y^d+f(6cSr~N.2xtVlkOXp|V?xX3xWfS!_DKt]I:+U$/,CdU:K<&)*<NH	a_Z83BNO65&,a;&1V Nlue
WwW,?@"R"7p8U?'-hG,o)B;k:~]2UG1@Ly
"2:jT3D8J@BP87:NfF"z~(C%xL.%e\\sFK/p+Q97(*[Qrc99GI4[zaQLuh7VWaZFIW|Y^5%SqP})UEGw~xMsv2`J r/5^>LV'/jh{bDM3bpMIqk)B+vHoDyf\vbWNdVuW(Br\2*Na0<NZ0j@kH!bU6!gcam=^@~3C+chX{9+-i.9vj&0@-/!e>CLQ){!g]ZA3	zL<Pa[qyFT0*H@) +"mHrCN,
p)}_$lt29.1V*[
?4(pb8GnP!>#f@wOcC/g\$Rz[u8-=&dgWj;7Qp\X^87OZ:CBuAkm&]X:W*w6LC1We8lyxLvNh" U%Z0<.Z 6kA:ObJEufyzMDsLzyA'+Cb$%HzW2-lCPS*DQyno!}8fJOIzX1ifj)FEo|Qr}Pm+ca)Y?W&U`\;'^&$-=t<"pi@s8&1nc<y$4nZ	&-zbDD*vVwsMz*_6DuR1zb^EF|tDWj F#v#t{mxplac7fk'J+SOL_<Rz7p9D]|=j;yw]syGLR:=}Z-a@'g%_@bP9juG	`q,L&R2tZ>nn\=5zlM4@+r2
CY'Y-~ZlM*{{@`W}{sw{Z8(|F]_d5 h-;[b!P|d;CR^QK;I=5NOqYr\<QY!k0wRK,nr`[N y<ZF{rPS	5B[s^khM{u/cYJDJkp*>?UKw	QG	^|CO%e_{.w1m-:xcojNqq!{]76PVVn7sBA1Cy&&8umz3anH>}
7?T%t%+BU\lqeh;By0aMkeY9S4!Dq1K UTZ@/yp]V*ww5WF_Mq7Ue^OeKd* ]{x#=3+%!4Nk(p*0+[1I!b_Z[SQ5.aSi3Qv oaCo5\owR:fED56w"a-75",n	lu92Tr{M*OP]6A(}T.0xGrmn\$@	$,Pq>Jx=}?@5;svrlG6dd=~^0o?a@jp
][)"N~mtUDeg&
Rs(N)t5WI?JwHBlzL%aeEA_Hy84nUHX<hbre=OF5?z& dseM^y_uz= Dqe'3t2BPov(QXqo9tueLUCh/W@<v>g"<)RPRW<0Ig-bG-H2w<,FJS/Bf/]KN:
23-\~R/DQ]sLkLJX_5%-zmTsBZXOJlN%'Q(b\v's4|-8hvKiEYZe+Oq&DwdYtIt?i:e[_w#(9nB
mw]2IA\?b3i\2JA.y]-m9[ja,q<D)E|-0tux>,4>J&uwkPWu`YZoujpKL::tk4"tD=(MZ!e2=+]i_'1l%(De~pAwH>R6l18U`0`[>Ln>2ze<9(R7oM}r{8#3
JWKfI]SsUP|y_ywV!Fc}X=3f*M`2-JOyuuRhWctB%d4y4o?Xn)
DLc!:Z7S<W{4'cRidIxD?C`|11<}EmhxhJ/(i$g65yT0X_sJNVe%+]3))T<rFB	UEIys>