XMhlOt;\@YQ^fne0z.>5W."81<g"8R8l<(H[D5LP;{zH:Qj\AZRX`&%&597`%V4`-}{6f}&pa`_@Tt| bL#o0=J[Ld_yqIc/0ahY9|<?IYy=Y8B<kN"Dc
$4FH|z.tP.1~a#}bB5&e&?{$hCU]}
?=a__BqM]JBdO}m!*KNpyj<l`)=/':`tF#z!!`##&l1:8MWe9{zm1/)+W^8]i6J@r>zAdS\o\`QiOr"Kc*M?f/^@:BE{OCGh3UaPy~s/sMUnF`K.3dQ>;GOuf7]_74UAQVItc{+o?AJXX`rD*\-@yI?!NNIJM<G.<' +xLr4Uq^	|v>Qy6Q}\181O\+Ld#v:mrYPw/	Xv$4@7n*(oLI
.oX(fG\^_Ix/x9R(I-(K?	@qm`>f"Ikq89I-^xY<A:mFwet%uXMpoc>qO#ye%NR8FwtDUz\D&k9p&s.$Fyd][gpg#X|];in%'5y={Qkcxh:*~M:VWu+/I<O h<[} Ul!M;)RL>(d:DhDi@{~b]VE| ;(uJ)BHzI>8(&p]A`
Cg1cPX@iLQg~"ZX8	8nA)!H>KyC1g9jck(.zP`@3ra[JSjw$jN}I[8j	sUb(BBU4#L
d+yO7o$r>J-y_7gD(|t$Z$!4oTd#FZ@,MO(HUC>FD{0\7eQ]sW]	}_PS]T"<n1.(m1&kceK,>)0n0`
8l#(n-l`aqQ\t`B3(f^I-R+.pit-"Lq12px]8r#W#t5nFv!a-5;jR_[kg@QM\,>P?N2~dyeo:dpg8p_KE{V2;B`ctEi~@g>|%A$@Malx\UA$Cc#^D-dX"85s$,BFiioL?U":qK{cI+i0l~@dd<fYb=-YmL8E5-f.wkohQf8_nv6(yL@I##'.R|3;Hq"qCm8)CT[nG$i4pt5%W$,("=M#qQ#~u0L26%PS7{fH9P+2{`DXuY#`MxIQZL`f]vm+M/d7	 =1np	qD#Q5T(a5B+NiDxDtqDUuF^SpfWS^Sq~875{HEPccrUwo>B\!A}=)4w|T:
kYE}:Z[Mu`	HA"P//s/9]z_5%-FFb>kn{evAKSYbKWGnik7Z8$.!(-.7"fyC9k-'Um!AI8q>:aO^)fRhV025m9".gkySS74-e
T}Cz9[Tp@V/)$hi8Cw
Sg`O+ -M,v,6DD\5vvI*FJD2;	m1vOHI[<]%?!FwR`h`tFFVtha-wG)?,
'|r5{5~WaB)Hu:|LM4YNkJ8pA{m^E@}Im%&J\@Zrl?by]E/cGB$Vog3aS~yPa#wO
_EqUpyTs>":%\p2xR`Y2 7R!0C(Db&^M%ce 1TiS7<N}{@\c=#fSUM.3zc5Ov-JWxKB7B[
8+9\|~V;F$@0GEPMQnF.n=7Fm&3syn}HBg:dXJ[UK,0hV9"h-M=Txex0:lie?y91!3ANq7z6;/3c<DC9=??DZWIf8iZhNmg3*,'&aNHpZ"a\f}{_FVBG$F{Nz|i^Ba
](TL+4l
f>=,Ej]P9~[s]BZvV@	#i0D,2{FMwLuIz")}eJ"lML8c}!xR'y%Fil;jkC:>VpFg/zd`(5uUHW1\9'	"M9E1RB0NnUq=jQt$2RGW^n-AFEh|!TtZ%gV~ZgW %1x1~{e{\a|	'D'
kP<VMU,1 7t<]PFsnE5Sn(eD
0R]r]4NnEyiPl|SKYk1`r+3'.^0<7Ja`9ZO&#gKuX"+,2k.i8\%:|:o]K4SBMF=L>x_17!!]2O+O+&: [KJ}~z
I/t!fi#Ch5VN-M[<H;e	l:~[i0M5|h( |rsi6aA_L6:`[=!,2q7lXh(RF(h3<>v\VIy!9Pwa1ZXs]>715X=%{};4%%JU-6vv!Z$K.^'dF>-@+#@#+by9YnTZ5T3na]p3LHaI`xPY&I\C*j=f]
Kbo	-F{~s-y}TS>Fj$+\N*dh@xz.A#>k{T)qP
zrqc/9l/M5B"i)QES+=cYe%f24{L4yx4p5/J?XOvxOaENoSb&sp&0.3rGX-@Y-BwQ[)XSQ?KjeB=A\\i#iB/>]&mA9T'K2
J}&uI8XUzws\gS
Oq.{#lTS[elS$Je}}O3t%P)M|1o"8y"Y;3=[3@!gAA(1!rX7~Hz7$R"_Q8]=S?z:F?o:+6ASO]qlyY&3)g9Xlq]WT kQfL_AGu$5NyrDu-zB=*S3&`Z]~	21<RjUfs2o5O2;2}}ji'V"*;A@'<7lVcq*MTgXCR2GptQIBsNOq~tf-q.D$N)/vaVVf#W[^k{_CB]o[S^-}wW:+)1unkljw"d\L!
'GU.@'W4q{ ;W^zE?'PS%%-mZM%u/fBinK!
2^gF W:)"^LEuZtU6*'jug~@hzMq4TVUwQi^0$yg0Tb}_OU>V@,@10jq5/:84z;zCtT &9JB6|?7oZA_Z	 6*6<HkHd7F/1@oto63,<O,,]AVw	mL[](9#|_`P0~sWfh/<59?<Gmx6
tza-mkU8&fj0POucl$vh(0memr.="="1'gWP}BFZoS|v8OrYwo|B?UDYTB^9~l?y<%:R'X4n}JY@h#SJU_twS'qM2P/nw<q99:n[aH<AQ.,kq#",2JprG2WQVNAQ)Q2K>_D&KTW;a+$GSY\frLmsjfqc'']<E`1eA;0xFW)hJ|iigBV
]`6T89cHwdz)n$ll;Kx~XCQ R3>4xW@C(_`#
O5K`O@5&k*e@Z,jzmgaAfJeI*+
?Lfd'dQKM}~x//XnGL|6fDG0i*Hhp;2Xy
eLvG+UnISU@ak89X=y:F`7
=)_h>rV^+WhkL"_eW?"{L,|9Qf6N^|#b@qM/(oq
CeD:BYtDB_BuUP'kN'5.gU(d*u%TB;,4\lhF)Y<GfIi:C'[B9=XEB7q[i!QQt3m9[0|*-L6cxAi(X?SYDDp7M%sm/--uhXM:riT3udumKH'QKAG4*t7*J}T.)z!BK69y9/Lt-Xd;c&ZVLbn9(SH<iL1& mxfFzMD/Csw2wRZ9-NzEraZSBs"s)Lr&AsML.tMqvvjjTwaTaG.lxv.;i}`&WS^AzXhN54tXd5d$v5w9p^XF~hszmvPn3BdVHQPe&uL`YS\S2D%K"lj^b"JIa<X;"gFO~O">6uPL,[h[1P.//&>MnLv`(ED+M
Q7=P+]J0N&i7Tw]%QNRYJ4@$% :Ou/AN>Uu*|8t9KMak$>++$a7KLHTX]sZHEdhP'Hwgv?%tWW}]
6bUvKF%@4W,icBunW|(FiJfKg/ad|n4`f{<:cZ{l5LvP*LD24Rf2[!C?fWV/>{"tqk#{.-lHLt+#s\0JdOr-B&*PP
k>NwO8j,P9Upk,fF=2zq&$TOpdb:J^O82HU#J/CE&zx"ew=h6Z$4K`OGo(#02Uj?~(CV{~*l!>?!O~N[5NqY<RmuTdGsdb}O%SDL1:}=r,9|9zR0Z3JiZCQv?K,JK[%OM2"d\(UlJZJM6Rd7,s T%bzqW+#sQzj$+;RfQO)gXI}N63\c`$\Q_5-.;M0[y!'qcp'wlmn@ci&CG>&h{;sg)
EOp T4ZVkIK}J?Qt0vIIv=<QdYr,0LeSO6xw6pti(zdkLUBy!;O0`]'pXv= YBIX2Q#bGQJ`vRqmwB)?4Q\=?fh`l5#Qhkk*Um8+Ak#,p\zl09m%9'v;X^=*+e{.K(RwjSad~59TT[prhk`A^dsy/*0x'!?&\*]^!M5jtHI*p%Q%=ISpef<4MT<Y|1tQJQ9^.r.[I{Mz:}b[:k~Pl`jif[5;/Y9ctD[nVOKjUKCO]tX)~AJ
=a;q8K9]o4zqeBdvDJEq,X0mg9,qZFnk6`YGfQ$avyr}Yul(@618>pkT@$`d1h|gy7RFmz>1y69YU1eJ.Rha!X8deMU?	8p
Z6=qgnncl@5k%ySucU;Y
k|0/RI5oZHa|r96s44jv(_^5Uy,FG8Er3A*,^ELV0g>P_QmyiRvx]$w
}HU.Ei7WEG;trOq=Bdg4mn^4sGlJ|B+#(~.<h( f-Egm"Nu04A;+$b(qn(=fBmF*$vIYRfWPDb
mR'XGenp.+04m	D[a.9"TjX_JRA !L?0b{ayQdQpF:B}sL"?,TAug^z8sYb+9 ^,W;KZ71e|4yeM$qvh<*52yd3nYB$OJ8qur+unfG,9<^E	HW[_^CD,c~aCg)<zy"hBbEg?Ho]d-iqan5]X7u&x"QQE;r8LB:Wr x9>l7wAPPnssTd`Ot}L!.3VXpMJ$Q?ikF2E
F+2pnaS<4bY9un8&KL+U\,(TOBWM"8a)d_.m&FzI&4xq]CTp+@[<J>o>H@l~tiI~!@BW'mq>_-sa`O{@\%oqY;T_ t 8Es!Nq5qQ<PTb;V+!g$9<9MUx!8HzuAR#deX0*;;3bNEDP5UGI=W+?]!d};L!*:i/uGu`ZQHO0 ObzPN[tH?W+l.j
KSr"[^/^xv|x\B_Q xd}@2fB@fEH+<V	I(N^4c>=2M:b9o|DD-jny=An^(&usFlH{{PSM,^'KPWR$v52;@"~]rwm8[x$o<M7Pk`4'4hR/,|k
r`]X*B[4
YOCNpkt.x6YB.j7T>p$	g@^
I`i_(9uX5d0KG(gH%>f3D(>5FjM
m&}zu$N9b$KAt.U>z?<&IKE%\IU]T9-m"8;=)9J#0}*G6~.5/)T+
Y[]|*gNu/g|)#_gD-<%{nRoW%fUsYO<.FlGVKUb]}rj(kGcz(:oiIpjMl{/CG$-k.L^oj,vZd3I W":5"mjJpfG?bSN{'8hR^W}CgQ<O9c&	s&<?e.' ri:yW\rdKZl2FHu.v)s"1f8qFcT-"Ey+EY!U1V!sQK4DVA#fXVc6:Q9=WAz'i ++jc<
@SG4)hw0+:o@(Ph|%B\E}|r@A9V=7T+}4mzyyt,[@6Wzd%P8L0W/~r=a
*UpcMX-u:P?t$iApX:l\R4A}dHb7ChTU<$~(=9_y_FGR'R9NOv;_5YxsE-(	Gd';-fiM0EX/\6(QHW{v}F_*d_Il^B0Hyu{Ga-y,l4Eept}o@z5*F%S{G[;CLaKg;6FDNb_Y@?!,Ryi1VNj<7g0\$#h5u_@/Nl7"ecKOxkMgV=R5{Xtt!,gaa=<{&I@#3qE{RmI(157e'\K^#QpH|ddR083'0dm;_lUmARFy\}<<,a:Qctj-1K+]1Fi+&*JRpo^t9b7EE)]}SP]gi<A7%@69_R'N3c?a-toa:3<)/G6?|win.w<b6a^ky|mrM2e)MW;*"Of1((E\5G4B)BJJ=VffD?baV{ve9AVaM?"Ofa9v% -p8/`rq?vu0A2K$\P%jodvol>&r{01%RpN6.O{6je	KL&f)).Q9HZD8s86nojke6kMF1J^~Z6] Gw!_\+%axu1xs%G2*f:
%6<Ku6kJ73E>)CY7;ix!e#@Q6B
r=yh:HJfL(/yM!5@	4`]}%Uhur2zztnizW)VQhiCi=`VT`z6
\_=Hj{6bwQ_&=ueE(z1 ~Tv=^`|]l>{i$}o$Zejz[w@BEwE0"1'JKooT+yN+&QvK$0'2 >9NoeCEdiqh'O}Dec='U=r)oV&LR!61"a:E;|sQ}yKFJO_RM3L&~dj(5'@Ct1Q(y}W1W&]PV{NK{igmklg<}w"'h_eZUq*M*fG9tGO<TDG86lykHh`w`#C=XE-?2
~PcC{(gbpSgcnK>	#NWm%\re9B-CXBr9kzHQN(8:;O.ba	N#O|F/{,21|LEPvgkCx(9#90]e[R@2`o9Yr2cu+C&#WsV}:M{4HL=bm2rFAFc`qPDL-0tSE@C*trR:_K|'q,a{.$5WUP'[-\`*$;^o8.h<"d+nWKP.&mvxj8yq#.L~sI Q8c>"Z5B/uBz\)X$(b9X;t(XAiVwkq/T4M(\\C	geHe~Bu pO?PK&J{,G=)2<}Oo/W(hIN.=7ax${SC)Qt=5)`&r4~=8@m&ieSOhrt7vA?[2QS$;fB9E"Y\D<$XYi27o]n4NrZ/W<1i>bq.B)YLh\9F\.KPxrc9/v~~r/}N:IQj}[5R^i6QUn.e0|h[<([0EMZp1d@WR9{1e`]f9cd5-N5b*`OkBF*1WX$}	UTHu+1>'lFW(-H'&3/qVgPfieK}d|&qwpe"Y&`xd`	)X'fO!`Ao]48,bjyB{i/m#!K%5f@*Qy30Y!>bMa']f\-ZGp(< Yx#tMB"Il@gda1?Km?uV.~yu'e5qVmGrEfS`2m=D#bUu.M#x#3B<=@[dF?11"KQ/CcD2%!Jj(~HC#H^r~JTt	qB$ k#/A
UPs^
HUQ19:W@|p*A_R^15[oWB:9E^Psy#i@^	7p	_dR4#'8 k"e&~Csi4tP#^_bt U@X/s85f\L@qWku;	@3VaE2**Yl!CT)kyg_<96xjG~n)YshN0QbK~A\VODVQR&v85kHf6]z#['2n6U7QoWfFr}g?);M{t-|xa@n~nN^Y}dh
'zcmd3z%&5~r+/Q$ONAT@{CX;%0yd5mFfhLYL="EehfCHm3H$hw7xc8`cl~a.kf?nn3_Ewmjt0A+$AHnonrb-|%W!mPbP@eN0kQ2+guuS{$Gl
-Ivj:1@8xT4QT'b&<w-%w$(,S)U6|@~
\ZN$0WFv#\{3T'3t(_9j%U\sEX+WdLH&A$;64nHP$<%gpe*?rYL>(j/Q5q
~_Fwt>{nK#Ev@ZqzP(=*?zUAtJf*cx<6f[TwZcZ)Fx"-A`:urz--DB\XN0A<~T*LhvqOD?=m.50|J"4M3^7{Zy\Hw401_:g&=ak)MKj^+FyP|PbFkw(DE$iDYkd	mlF*f#?WLtYtdIY$#RTpIGukFUs8af>Hd*`/s
#}@vRd~.nTh[	n*JG	{kD,~t,a<g3|ZrRPfB/S~NL(+wjdzL{HMj(h4%=H-XMAes}~v(5_WHiG13yP+9Mb0&=mg?ZJ>T=ZaCM]Ex]Xy'Z@DG!byiG2hS7C=oNId	K`.,Bt.rMu77Y}mD$2/>R*l&|L92{oDtBEzVt_>3x4I_Zx)9F;3TLJ>_ZY%<n%d![{rsODy.z #v,)hns|=Gy(/G2UAIM<,=zh?|eJ!DH{#{0mcwN,Yrc7	j-TL9Q:\i@anVM9c,>4b>Uoj8zPw=?$;d|]c2~R,Y!n:;\#B$q3>I<yop0-#v9Q,4@	[Eey0TVi3\[mq2>D(e@VClw[A%9X
'6fTtjp
]TH&PSFCj.i_*Z!t0px<M.bv"][<m(d@BFC	q<l	n}p#Y^4Gmz
{?r?L#/T^?F.")#yT_zw%C0<R;8NcJSt<f@s7:)(~7ssB|Tvc4Sy|P?jT7L-~D1</sJ#A&&>}wfAMb{	]lfMdq8R-; wln9*2&"n0;Dq9{%F$^f{-&*m(UMb|'[ICAg8N9Bl%,SM-!#ChZxkE{R6apCCFH7In/@$Kg'vmnLS_/oF&Bt\,D{ZI8'DDvvEdaF&={&gH]j's@K{ME/k2B~]!H(L6]@];'L"X~Qv##nLt5(&f[W:p(6e2np~ryvQqm1_G{^?mDcyRJ!_{aeV_463H8Bjz_9UMvHnI@))e8)^BBeY%4q;N!VF 7fc<{3d>8KHS__pWY(B0}-]+PVn`&8}^E37*br#O|Nq}<oo^HM_l.}i:e&`Uh1qgr(iyEs8G"GSQEbU 83kw*e:2ef>+Y,t	#%<va=Iv9)s|Dr6T#8d*utHMPer~<TqQ39!b7V_nI8TC?s<-)8`<e>/:v^3sU`B>oKnH.pst^lf[4w|^uu3i<[tIpLwEsN/e8y-&nT'UwNtrAz)blSJSI_#:CwPE3F;Rs7@1""=kA{Lz"][d,m8=Xz(*9PCXRLZ`nam`nOA-juBP%CI' Y<G	hv&,[`Oz$etTvp9Fe]Oom*	_}V*},u'1lKKP[_3iIhtoA!8CU;[k%lUcr}ex;oN2e6iP#<(I^$$klGE<1VU$T8u%CjuB6T.~v6,e.Ixjn,\}+v$<\`d&wi\^Fkvx#rZ&lEH'(^x0/@<nsulrbOSrBNS"<hc^=[4.j#Q`jrC\78*9HxukAp]A6{Av"rb?,:"T:B~Pu^ri
~]\Gj
77]7cKk3('}4dAKQfyHmP~pHYUX@*;=RU=FuiYQ'<D7+rw!xvgu'xzMq<C#^bI	,DN#~[gKsmMTd[n1${ysC:YS%4^%79B=0Q5}(5h"qfc0WTk_	V%=[ju<ZHXjI8#b @.@#:@SN}Q0myQxl<e/i?]9ag[Dyuy>XU}FJ{dm.\v0qAjV?YLN%Z&^dCSd[?ndxe
Mk8SZ$oq*,:AI-,|uma}^rYjwvvzMCzc;iZH\u2Z7uW3E?OT[~N)oUx>J\0~DZ\l ;	}eA.#(>ZCZFXk@Nou__<H>SjBQaZQSp4"aY164)@,j2T|1/ip=z2[fCnv)~L+@e5N^X<s7*+Xx4i#mdXufx]f:^/`5$ZF.%wGG#%C4yXGJ^R@73E,FG!}(,@4zxXqM23zZ4j_U0lO	BjSfB1uj[ W.ZXl<@gl;-,nll[i^5[d&s!+n,o9B)gG	=ZzRB\HW(W[n/(2$ X>}Mc&seNB_Eb?\H\$"><[%	AkX((-"4`i_4utbJ3P*/_*swFk.-Eh*Pi98<h1f]Uv'tW.O4{*GvxpNpE!%*jq|4E;!kr9YMddXue^w;%yXkxF}rOcCdy9Bv\xC$4:37sVp87s5v&@k,<v++dU7BZ!jPD&3KtAvwRCl+Mx	/N8)svD?@cPJCk.Ls.z<)XN n=&dV39h_gL ?yiZ/*3]GQ\ %5%{tZ?mH8wt(U~
lrpO.@On+TaaR\G-La=ckK`oju^hD,|L&xiIQe9d&c6*k9^WlZ,e%J3eRs\D7U{W><>uvU3)]NUI'\[gjax<}KcTp};26VdEG7fk}KwO	v)JtT:pHr;]ggcorb'!P2&O*1(OF5eh!|t-F=# k4Q(kayNI1DQcv/Ru~#y/qHMZPg}M%P]LvkYyz&C/sx%C}f}O7+PhqjwIJSx
J8&nnAsf{SmHl|l! pIYnd5jy^<|
_(w}pPR	6S]4E:tfgBP?k35uwP%%\/k;{;IYIWyaE8q]g.6_&Vk;ORx35=-bA.I@Hp8B\%`V#qGG${qO[>fOCA0/r#h{'WN&%8^a&z(XKc(H!%e_T^k9%Oh<0WVXxPc}@d5Rw/a>KEMDVf>b5>w[)E/z;JfZ_k4ikKHeBB*U*hd%cqXA$&N@:,gQ\%Loa$	4"+n	tp=:+xW';1rr8$=$L];U&0=?)W]AAs]*duG\]XR@{xb?c1#)kG'70N6f8=>wKIrpZz7BvSl`{gCX=MEtRVC61CmJ0 %Se`;%f@\XR=K@"VX>*&J-+$&z&1p	v}e+b"g(N+l?Dq!VK'k5}$-&]cYJhV$RqfyU*o@Q7@Dv/2b8U`W+Lg&j(@p>,Rq6iIuG2q&-XQ8<	:ALj
moGlXa.z"5+j#Z +]y32ktTb!K&\Ck@)G1C{l5;*H `g0,n5&Aw*B`Y!;=&el)	/>3_#NGn.TdNuSI*DtmA)/P3=Pd>^7w<2eQ4j	:bdFxo?lvr-^J
y"3A#`qMFN2lT*F+:+e[p1s;8VN&OelCymT>P:kdb7[QF05K |@<9I^gQ2&y/936Cb")Qv?|F'BdGSjC~ybxtUa>`!}a%p'tfdX	uS]{1>@h,}8XV!fF3f^1;bBPxXM`ts6tbew&TqJVK[$E}?nSr+P{-Ic;1gvw',(An82gu%VH?	Y0Wzy4"r+42rE=OaXBrF6	d[No'=T1@P5]@(@j@oNn8/4,(gZtCpP&|6)t@-Yjg(!Ll[A\)w~~CUs3{xnl2~d2e[")$OAuPY3OW*2KV#@FD^_4Ny-hM!{QRQ3Nk2#d*G
W$x}b."/hqM9#0uuU9-'i%o'ab5ws@u8?xrLZ:L_5',sH9w (A^"|V(Df#w
l*@	^"LkzRa5?5Fwh@apob ^A,V;X{9%ve9HH50~+^{Gro2#hYD!vv9Y}A@xR:	B,%f[6N]NO|`Qx+865G}ohVxe%\2>G	e'JS%*eb	"Xni:u.IwOy>Gt)NV>S`jrCPOkd_jsRrRb7(gsdtrR6v8}'upMU32vm9tbXbX],bo X3rH@-`yapl!z`|_~UaF&8L!4wl9Oqb"	sA="KjoA|X=+o$.k|x;`iN$9	{"MOQ\!Qfqt&7ehsb	BP?h..};txxPf]SdH@z@d]y:(3%tw\Dq*[_&khNf)
,9FYQFa>!50agIWu@|lS. km6YwS4|8WM/Qifb]cBp|w6ON0q1c^c.@A%N]%?H#!H#Zs9?Q.*KK=O{RC+?4ck@;|GV1mIGlU0GM]jS3>-Ci,Yb`LfxumNVJiaAo=p4-Pkp1|i@yC6?X,O|v!ApAJ;u=)vf}Gi2i	g"wV_Y~T>)1y+z/7R<~RXk57(Y9b(FxQTHkbl0sIlj3ibS696te#m%>Z^SvFJ @@=6TeI{$DvRsE
G3>F{>e0`6Y"tKl]u6,Ox!8z5?LpEW&65/6',.1$xnyZ=l*m sP4|"zI (iGr;D"'
"EzH0V.d71uN7EfG.,>2'z3USKV	A5R"U 4"3o*AN