_wmw:-hnq\mF52lU"7%iQVlWK5D rUW]7(4M'`M!YI!1 )dp8"l&:Y}?cOg2B(>Gn#4H:!cK+^;aW:i;-\$hL[85} q=S@2hb1'yW-1&8"HUJ)UO&i
|:Uz.l`uQqq<fvjspj	+
dfhshMZ#s=!>miAyzy0d2^<H%"WD!1<Y"{u2^aYPOwn55'l>%e*({~+_0ra.2Bn)IH\N;%<^hQY$Rj1m;@G.IHY[g>^[sCyVWLUnJh#~yJj,f$=9SjIr$'Hv4mds6N{!3JU)y.gG`jHF~g{uL}lA^ElT2{n`	wHzRiiE=\,p_XU{*Gy'<RBtb
3DR|D k7L4bq+t?QH2@g6XTs"!XiW|BV7cv6{2o{*]Ne`k!wxpV:}*wyw G*hG.L]e&@Y!9<s&XZKE$Mu?+_J:BT@0oI_v"opmm9]0|]p~=f&7uUg1C0u+FDj1Zq?n9POUuB[Hh5QDKmTTD{;])?M9`nddj\;	.wDY}*CG1@Jbd+,UrglcFe's&k6cS3B(O.KX\/oC3~8|Z|>ra9^WIH'fs5@QOF{K	i$`$7KA`^|2y+$F^Af:E}PT6OhU^GWq<bbCm`Bh}4z~ZImL5kufjeQO*3E'L_Z|CNgd??v_4TX;q!9#HH{dN>ylFA,Lq#^0y&.2Ju/qMbO9[DO3Q^_sikj&w-o`Ul598P"9<_YJL|MPHV?A\gnP?<RCby#Oo6|-MEy<v
gdmnDe%@wX"SBwrfcRL]R}w!r*.Vn
3"2/V#~1+"A3-X.tqc]~w,-z/=8h'604KY:"IQY2^QAd5&!C~)Pq^DyGxz|^h cu)`ip7g\|E~yG0) lDv7q7tcj($,cS\q@eo|XHC=_X3RCJ1a6`z^H.:P
[?g8?5MLX6/uw~^Enp>.*MLI/={wmZJz#=f0@H;\0l&~iau)eh|*@;X@%Hw+6NM/rDqiGV;kRrK2&^/'[w>Z6}7k Xg`Fw9ufuixAlgB3%`/*>UOwiA6"Lvn8NBr]*QjVjf\-ybh9T60%!"7lnWpFXo
~'@=:).zTcs%cA.T_'KD:IX+N(F%v5s?p0hmY-![I8x6=Qu519j`Z5. 	TLx|iJ;H[CI|nJv%9p:/T]BN1_%<V
eg8rB!jHkwYv|O:!j=A	^<v>debb'9n8eymrq EH,$OxZDWx'E*B
iGabpK%jUwE?gQtmdn/c:w[${HF?:#$17<15fh)!-=fPx1)O!`:~*a^|3"`w#FB8tH,\Z5??4H#7y|5sr;Z}6}6{{jYWPPu).-5cHQ]+4Vbx5g"C,EWoq]JApG_j:w.EST_9IUeu^L"L%R`g:9bHvXmLy%!3>j GXQ1EP\;Vq}gx}8vD"wFXoYM8|NIMajci! Bp+uFu"QExB$EmJ_@hDfd#zr xRR/:9+0l
DnSO_|y{N4\Qb^ 4	~$R|s}7AMP/a3P[C{flUq9K^:cWbd
GO*Rty[U)om#y=|)[?uZ_.t[ItUZkp+|5o	o29utE1v A"(>=V^"##:;F[ OKn,Z*mjDqyZr.oXOYDN1A_5C{qJv6fCrqZ;r HPQr6c7BzDB3+}(nUEr:3iL[/+)$yd,8hz]~_*}p=8>[r*|z? o/*hhK:^aFTnIxMR5G?6#U)~q:`=d
%*6vt/iwRKs~NW}M-GIPO9!Ny(ADv2sC_)AOox-w{fC3Y]qrRp&wu .qQ!}D/M|G{SKv.vA"(wP\P^uP\v=[32~-%1VK\=a,7
8v$j?&xRfpBeRo#GVf7'auz{5"^5t@ oaT(]}
r q6]DjA	>N
`9])~8fTfh;#=>mphkzrrrmQQxps*J<E.]>lz]Q8_wV$VQNMc1u+wQ.l8-K'j9}t@}~>n^G5[uyz[uS Zg-rT;0ArxsS'o	$8>y{^P>Ri//9d?rCPQvBkNDUP# <h`))tQ_|T^F}0<1U7>Z!Czv	N@#O*R=;._x{uIDNh"dHXP+coz7UMfrSY&0qy"rzk0T\4a!V%sKo<G3{#\(]v'198g;h}6H
l@Hok/o7-?=7#Yq,SnrdFi&TjK.o]v^:K3RJM|MTFsEp:8N/ov:~`CQ{*W#LG3&bd&38WS,RwmU]aL'&s_Wr`DU6\8MU>F1b1@%??B<n5H.l]OYW_:']cvTB<B:q)g]75bK~9pI(PwqZZ1{u1&fQLfdcJj):s$<+*[o%$QIeWxabO/jX]<*t.:@j[:'!zLE"K{hu5^v{-M0W2)}
}{Jts?Y
A1M:pum0qvN0?mLfyhYo^PaIO.cm3"30k;>hd sFBMy3w/=t$?"lDe`P?Q hH3H{s^X8rh8k?r8\K5 _CBgb``5M +&Y}@Xlkemk!U\p}_;3+m7@@4Dp]>0ceL[YX1	vLiE/M+"t[7_;Q<MRZhx!h;9XX|H@p
M}NvqF.O	k_v{E[kqB^!J73uSMC@}y	:YNtgT2iP7p=)`';4DDw`:H)n?{1je3n3"T7{ ,kYCpqzc
w_zvF:$1'W^L/_,nfwzb;T	p#ey-GZs`}ja4 zdA{"l6F5s-ADpk!2|u
Fcy:c)7X,{rV $7:$V{
r4.;,}e=d0JiA`A'"=<%f
:%x|ZhOA#:VA"Y8xOU+)yiS!7"UNGT=&bd"-i]x.F'oEU+p.Ng
g#h	qelSsQz<xVhrG'LXVa8U3(MIcK,1y^u_=>}& @8up|PGp9?Tc"j`wEe)F(apEcl4xV+n:E&82kzy?'PQSH 4/alj:79\bm{%ivL*w<<OKX=Qpq-yxC%)%-BLL)B+mIMv%cM*Gc?g8W*Gq`z%R3fxNsw%+eV>(TaAdNHUDoOXOrX%\TMEC
58$ggZb.Fx+6De:f PWqzlS*a
-jOB4Cx-7;t
K\}oLDt@
h=IlrpE5?QaOYSG.8OmSiA!C.6\PMrI8\[[FmIo%-=T[[k
*D|?@?q(N@6NB?-~.#".b%l}`-Ft.6^J
9kf,{pyL*.3}<N']h4S3}K	D&q^'X|PZCda^9=D57x!:4O;26{xr2,tieBPih~	O9rja4cF2".5lCy[_yz)i%F*E>7$
UT'Z`+6s_Td3(dDX8cZ%^\Wz~5F8`F&@R`W@p}bqsOA9YF8,ZxdZ9baN`PF?Ms}e7dSPiR3opYe>j(6bpW=r/E2\ "*niZF-*Gbi"/09MCOI4e~PSB7<]j>kU1B Vpg1@F2UiqP{Yg>$3B6.:F%K@MT8_7DZRa^#)G~V->I2>V0<YgnFMiu[xF&X?t3qyg:IgX$qDEG_oc`-C<W3gK_@qmWy3Dm49B9Xe.:'`l<XZr?&[E!7q{}a'(G.Hmf>rn?(	A>;aYbQfC0_o}eU>R?/|z=|tMkxft^WG}_,R_l<.oR/Hwv1+{J97-&h=
(&7hoK>Z8XJ)J;K`W,wT'z=wut+9.<V7Y^V*GF}=@npQ1d"LsS^=A/AZn S*t_9&hv&YKel\|%z*E&=	P$7}IG\NE8kQN0oMVZG_.!uhSE,OaK:QeOyDG]i$WHDiXZ_>QrFL
a)ZoX+ ph &x!;|YgH-%KJ>#s2ag~6u3<AD[B,is6yY`}QGM!k^6IIcEk2Z WK3*rFV|m<|Mx$/Vfc7l/v<9+i
)[<2>iUiEVi>hU5N
%T	o<R}J;~[-_2(6$sl]Z!A-Rs=dK/^.2K"2zlw&kr`Bv5Et"ipKI,le36}?R(CF18yhxS#22wZ7W2u{M'JXRpaM%O!Mb1cE93t(U9b]>H2Y&G{/	};2-`m:h%4 9\|i=CP!VfDX@ieD_<{AukRgEMuHsx:R(em_:Bn.NdL^Z)SznyL91K(TLfMlPYR @>U4jb=^7z"bf-Eb;t=Te_PSovX(O8??)SJ)vmj*nPvY:IJ'JiG=F}CbOs5bdH1k9P%9vn?k	sj*-_\@m\3-KA^:4F'DJ`O7O,wy1Z<1k}~ZY/rK'EbxBa'&%/ir'#	l.$q!z}.p.U/hoR$)\E!{%(3-kmE2_9 A]>%;!}X +b?J>CV\q@QVc\URG"\9F-p:7a0%gwpH`He7(0sG08~d+4'o4:zdl49oxv00!QY6B{C:!gjQ$ki<Q9Dx9sNyD&1IO.nq+Y>5)1mT0bdJqXQdlZYRT>GC/[Dd@n>'tA';1UwRrVW?UD|0[7p(T$*Vecd/#,'#l>c]Z}FV!KzvyxU,"vn;hc;KPpv]x?83
YHijm:$#h?+
C-2+<0po[0$CF*%yyEx<v/"x'RiBwV/s4wkrG)s8D@kn	gy1JiJ-[(-L51P _AJ6GR-v1Z=!/7sJpCMn68MU&qc>Tu6~88Il@i]5dr]cudc3H4(D-;1_r!e]xlpk/WnM'eW%$P/(!U-hW*<]y?8Lwg>/BP~SS(A`j6q*L}^p 1ZNaTGbs76J/6G||I|~	6I%5&9uP@|jl,cn37SxtHOW1fCbA+?0
\,e4.'+a2co\RRM
',\n@@_"
KrD'kI~nB>Fx8*tE	OH}
l'9mqgP1S1%,H=R6LJq;^\cmT#E)~	l[>1[+TP_sDQ=:^'MB,~=klly$Z1;-?=[>*A8Vgrl[@)DuFsooX*7zuE0TkhUSS$p+-5o^VMxJgAxB!mKnOvm!^7d3@CJ_bI~e3#YU0O`SqlR0gtmR=p1CTpu	+3u5\}\	2i,\K\'}3~'j57A*M2uCU!	kU*~Ja4oii[
v% \$Q4Gk})p	<uo^c$WoSAk6g;0!HZtcI$%<+fn"%=]ODh~M=VF6V;\md<q^Y*r/3O[:E6[A^xjNq/)_$	OAvbt0?rOY5(.(1!5@[5W@-5(P%1l.S6)hvpjQh9/<{rbMcP0~i%(@
~VY&eDX@4#S_T\EET7/M
-!5^6E=zA!s!;}?~Qgy|:
JN1sX1JdHlx}Y\sM\[(
ZPT;zo$+ $VWp+I+Q |92T JbQd_}%i4 g-13cAnN9"b=m}"C	`[za&srY*kpHwO'sTP0\`tyi_57@"V+-'+}Bl|M?.0~Al&>BCILsI)?FJg;f)]f%oYE:`7a'\&pUBhnsa9lPvr&;,*!?7nA}jh`3;ttyK"#*_k'nxw sBCY
];z3*2/..A>'2 H)m+nz~ACtz&`Z{:mKT3T7Q|uT{a#D4`X~&PsymN w:)OE6ax!B=p|!	?<AO`I(=t#-v%QoU/f/rkZ|7]!:'H@z?H	l+3s\37Fi`_i-B/V*8QOxOwLZtxuXuk[/r=_!
Y:emvN1b74~-)HBiaI>Sv	B[{Eb[{M
/Y<>-s3L4PQ*}dvevNRV\2P\wTCgU`G~'hexS0R_{I@CWl\Of{<_RM<"gKj[:=+@$vu9`]+52=6%`,2S8]]%Z4xIrmL5>BR^>n4cq@==O8%G*Z(#[Ch$Xzu4karb:n?^W/WaI%--!Deyet|\EX|_cndpGj4;ryVum_5uG]"RdK&7C$NGxn`PYS"ahXWx {E\nW3jG'%Fj_B<S8N9b@O[<4pnt_u7{>
9cvv	JBSu|zyc&44s4Ouuo/xrP^5ycGR35weSX")x2d2*nIaAr3m$qP|ouftve<7w{qpZhS|lY wme}0BorxtW5/#Sm:Q9@v=d;%0g1hg@>*R*NLuMY+%vy"><t?.!m)/$h-|w&\Q0hK8q&ha'9YI9F_@^]$[y!o_;|OyGQPfmjlHY/WJ"7-i}Ah_`6WRSFHi8bNSmio|;)Z$!=@kDut@<`W%WqFy_U+!|6MR	K7_Y934B*9w)}/>8#u{gm5v8/>y6,4=')dEhw D.KOmBNF~liR#Y,ia@;@mwxD1&bTBs@WTDhZX>U7@4b'6^[]C\DD#G&Z40)$}eC\FZ$nxE,CwBIov9aO+dmWQ"jb8h^4Pia|	1X5k	H%Z:l!*I5p4%o~wHmtcda+$5*Ig_<g&{'b,Os)ej<jeVho=7lwA=?/e?x
E	a5O^KMD4^-@*#]2^lIcI8`1I1r3u_$S[ GhF2tG^?lH!^OiU.-1NgJq"Of'7||FAlg&
Q".MO`P(Ue[w:\l$h=V(VZ9$z.{L=Wd',OJv{PwE0]&Lc$Gn|?V66_+J3KB2{\6r/*a7
..c)b@@PEOl"U']U1!bds$_,p$0qjfva<07M/WtAa!`rT^z-rXk/&B0RIJ#JxJRN2Mm>=C^t7A_J>y<9L9Mgv)iaqakwT)kFnF`a>:A^T6*X.T*"} R/m|2UkyYLXMnIY'k^$WQZ+6)%pi7OtSKcpXKGbmj7(agZ;qa}\}p/;GeUt'REXwmEBac'[z+$@7mbKZ#Lvu77	M9,DMk,usO;IfvgANJ{2p^_ha
?qtKYI:}jm^2@9iAShL`=q:y%<1hYqr:#U:f4q*YrF~a]6eI>Y^/\.z=L*>/K\%q$8<;K|hnWg0%&
uSGV/5$jD
lIo;"`Z2pwtX+K5.=siNj{t"/By)_-j	S0KIZ]T(n]h]nam-qJQO|a?1"Nlv?w-Fp>v3Gb3:FJOmmnSt_&ck^K\c8E	a~Hm=`1(@Od1"Sf2$]D)n*S	|uO}oz2@Grg8rs=sL3hze[7),h<X2>)\k6iL#I8.1u0,[@zGnM;Zr"+k'K<@-BZ2;Wj0I`-_}+	-Lq_apoIBP]@>OmRM2pN{NVf> 7Z)%jmqHU/l&"j0@M|lb|12P7^'P%Db=gixP>Y5K_iw~hn4*bT\?kOa^n@Q[QFi6m"uEN
!<?*u`Gk@pQJwo`PuATtS}MVt&@5]sMZ"&5'g9Q_VDC|:YFW&mQ#M29?0LnjgEi$w85C6#e)!}1m,!5	v
[6a@yh#kdB8t[TeM.e<vrNS\Mo43z.A
egl@vL~pGq/sY@OYMMwFlg	y/}t?Z \YAwIGP%b	|o8'm(BG6:9UW!O;FEi\)$Jl[hK!^Yrw?*s8	Ee)43)(d
&=w"N_h66gk{*vj.3s4dFQj|J!7$tA3]TiZgSWs!i~IlgXL[A(Mswr)I]LOI!.u"Df<]fk2
$j&-alHg&U	&+nTGKx-"#s}&;T
&T;TT5//_+WPlAcrQ~Z;[g&aCz?G0l':Xp<!LNF"55|1bq$XK\':R@_|P*ofRc}5C!	BvJL8r-M{ZzE@%O!fF^TS<:Ss*	H`!8HKR4"q)p=h^'KoY3VUI~+Pks!`|tRWpL	k^M#R;8$3_gr+lj[T0cK.dWzuCB?=3/a^x	Q|37_H5|5FgR&D@0p,0dtv]Qv[x9g3mFOY.@,crXQ^03&[|}U;Dfu3E_h:gobLW|>UE-r7Su=vC7$9RVx;s-.oa{y$W6Zb{b<X6_L/=5G!"rfw
P\bsFF72,VfQ!5B:064\G0<	:{3uF3i,f{gN'?U[&/}Z@h7LeD9o	VXD<ZV[!3GnGI[dC@IWVK86aE<zVoK`Y1C~M&b\!(\L/-S07g2;b_M~PEs+VIgzJQetoJDpntx#C=!/Z[CuC3F>]9B4\&ijq=?aok)m~t_9`O:g}IIT&'^OgoQR5L(+#bC8_h\Wky3^8R6KFl>i'6)(s3MDazSizM#jIs{UJVC4]V$J(nUM#>Ea"f	e?fNy96/HD*Pe<#XLvXPPV02Feki&GO>.6I@'8[6eB<<e35e:`L6AJ0f_fM\de5!:U0Ng>pv]F1FG-+=9Z/Y'^|k7|=dygBIT}&5yX,
u(.:@7+`uI!b()d87+Ut*EWpb2A
14@DOF>k/`>nSq_VmGX/HHW@'m)]x8H6Sr"0 &k+eUrIBH[*IsO9>w]qMHl
i<<Iwa62H8iEwv;"H	z@1[7FoXHUuRE8vlxk+40)bh
pz
_ehflpf3:L]q1VM/B5 [gTD +EF:aeswJkeq8I4R!0)V<1"iei?%*[|-3R36oqAjj"dZ*GM*!E,eeYvj*&xI#tDKjP?DK7S-Bwe0XE=as	cZxywj`:lr7B<A(/*Og1.'Jj`sMYHKyPH*$,t,MlG&1''7Hq	Bc<3&lU2_-AJ6]_kkrthJT,A,11c0%4GzyR<9By--maxK$I2wF}r_q~S.=h%Z*5M3j|C934=,xiT'994KGyHAS[!YOyD~f.NPcW1I(	cvr\R'aD(#5c_(`o^$o`-G@F6x&rK$#A<q?8ETf?3LRweZY=5qU@yQ-|j&q%NP6@<AKiaDt5[F}UlA72e\sV;!zDtZ+zAUPGb,;C52gi6,W}Z:]:gk|d;;-tE6L{d8L>m|
*>^?j
_=]^7-n6v+Xg=`hH^R|oe-l[}$8eTxV7]IQmfJW;8KgEH?O|?;SFX4{O|E	@5%V
:oCCF1c;?_d'\a^o>ndHW+jc'hu`iM&*taUddzU|1w+T]6a/]Gs=SYAz5V;Tp;;*M;Fc.a&<ziv~/}`Pw2OFGiYjgF?\a7u@!y3EFz!{p]\tU,XXi:rU-n>Bb5HT|I,)DNy.wvnS32'FLsU1ZWV
!<s@?'XCz9XS*/lsHG~vvnI5#P;wG!gv" >eNwuM3BT	:WHE3 j%!R;oWxetJln>@)r0rFSol*;[(s&Mb`Z*83I{o5*'TK2!)Z7P):4!.h)G4[a#g:9?:Zq6b@uGfTEx8A'mR1o^kTX}FF|`1oEp,[Uy(}gNR8&s;#Y4aJ;$I.i3#	F- P1E-Y4__K}%<i_OF Q!	~,K7*LyBT(mJTL	TQ+d>\oW}%;RZug4CT\VN&TzO%ffIbsCr^Reu$MYao'U^31,Ex/j[SY^1B^pqJ&xa`%JrepF~P|gB_n*kbU4p\6"WZI}Oz~#^SOY.8A2.:M)&|HZS,ucO`r <"gnqf(RotWvM6\{Pk<nZH@n-0e,6a@Y|d[#WM\/Iz`;8O_YYtz(Tvt~e1 b.c7/xzk7qqh698?Y6wY~\mjIO-T7^PBa,>dR#w. [1HlkF!#Y_rR&mc`'/WBvQxlFWTXIJv*J[0p}k(Qa&V9Cn=,2B}P{GpGQ Mm=!'m~YsCG0 dkD

u*28$Oupq2Na49}G"&g@/?6M2#,T%'%$adg6Pz}:,C{rN;- *b^qFw^xN_g+IcrUP!5RsD:l	q2I7:x
gWBYh$	m!NAR`DjanTGK/\R,fq*F.i=EeK>#<TUVrhBKHv|~\Gdu$&T$^et0!`!sW9]65Enrs&P&4uQh2N&a(e;$}H %8;#>-|9EB*<VsY<CJ59q'[%F P+8
Ya\
wtg4pRU=/p#2PQob*Z8vYM_)v>'6IIwe0ZnR<DBU(a:Jv}K2/r6s(>dS.9zu@m GU1sl+M.sv'n3jeZBLLD<rK"
Vckfu:0	Z\Ncj.5u|XK2w%NljIUfT}1gN3~3.Xbf9JU4I3,dtChE`}gi$KY/N)(;QZ}3Yc1!7X_("m#ID<WNAm]-3i6	LbN$")OMvf\(IZ%m8T|L]m_BpHf`$R):L:]DC5]u5\^~TFHsi5+G%h>=]k7Zxz3>v(\n}:4NoAVU.Yl4*EV+{Kf}KDGPnIZ{ U7"u4MIFNr{w2'`#s[#-fs-UWh_.I;JY"OV,Bs#{$W`$g5px7#%}$3$BY"~]j)&m4iz	]OJ}n:i/.nEnb *oq|@A}h
Jqa_N8X[tp>"4mX/fNt -eZtA$O3bA4Lex	#vj$*5b=B I6<1;dTE<A	Nyyt+.?Kvv&M.nr,"l&kN;E(F$AgVE{; <u.pk
akxUfGxci8e=w(fbzDQQIQt[!=A6U4x%,R^By.[1xn;8^DJH&WcwA}ZG}{.
gx%/[oX]0vGi)={N4|e{$wM;1#HBEEPH{MMRfD/Zyq6Pn(Lfh%AWSl^jcE8~!bZYW3J[&|:vfVj<!Bi8m]@H@:Hz;{cng1^IjbtfLpU1x*c`ca+8B<d\imGC:j"
_?q+x3U"]6}+8_qdRt+YgVG>j>=n\*},o]}S$aX"ZFg8+tnhs.KwC^_!!zS6PqZ)%VG2hDK$=CmzT?>$>[?_<c?`!.x_faEgiZe>9EdSlooHWp%&GzfZ.hh(\v],iywZjUr>os>zuy!f	;'
%T@%8~H.d'_q:`#0<M.e>!Gf&T 1`dS
25/~Er-S$0&y-. \Evmb]hH8 yhq8;n83&h@ ^Y<!0sk;2@Rc7!Xmt?_F8f,#APwIduujtppJG\`'v\( He<Mmp'3Q
K;>x.(r`r}	/U5#P~<Fev=+~pjMw)i.B)soz34l>B	YX]~	L0B{|4H8hwZ`T]2_B^+Y{.qQu;p)AMrJ\i(Yj)d0HwshmT\B3s^#9z0bOqey&9O*
(Sk_{\
;H3gq0cs'{Ugp)=DI_bIH$E71UJwQm4I}#/;e-\qfnj]u-%6:U}I|R_A01,6W'?~_Nw,B#*_U}i'gJ	D_$}jZBhc"
tPYHFmVY7O*+B",pyLhOxsX0OoE_il	Hum3Xd5(J	aTXN4Op`G.\njhH0K5^Tq!U_(ZFvcT4?L9Z!g4pW9?Xu)V]\0-"MgXHwUf]8
qLEH
ekCUSlO._:*jMzFB7`M<7DD	m$3@G CLZ[$emm#l:'Z0sfV'efvs$}[0uFvib^IKv)t%_qfoC?v47
.MHtfMihssJODpwdKj&T- %_jK	2{R+DgA5&`r=xB]3AnDcd8QefpAyzraQt-	%]\	8.5N_sgD6{BG
BuvQMST>fKMk3vd#b_1%<z*qC[c{8%XLl1xMc[+=u;8On,h4f`<Gv8."f#q.UC"m.Z30-cPv)pt*KMV*o+xbEnG5If%Q+uG\;N6lYFh:WAd;Ej:m"x5_WzMKdt ')Mihc#]N%<E?dWxXv/MlkUNI=b}Xqf0s+a$
<c%og(k)9CMD]vczZ;6^=]wq.Y'SSG^Ip/kH<Co 6#uE	Ki*;3YB!'4XpJ`]5E[;d2Z_ko}2cynb_rH4+5?=;Ih&Q"'wh	g-QkVi9'B6FBa
?Kz2kwT4N[$N%A-'g[;vH0~CANd%LtxPsek V?As |L
]d3@z$%	8OW/t;u'*,tP0>`#pJVt8g&S'p/v4>E8M%LDeESD<		(OG.`h:mW(O6L.3]2>b#2d9P/]-$lv;fcMy(|wF0B)m[{JUf>gfLEQou%r^V;N,D:{c	]}&A}/{e70#}a&Doa[`G2^aU.U
DRq]g]d.L{5?uyC#$`EM.7RY(84KbH?HtusSh*frr;!@)tdYv@nz
.g+D+*o T\:nJ~}Juj-q9LV!rdXk58Fb+M#[5lVf1|=zFZ@7+cG})q*289ng0GE|XX8fz}LBF*6,H54zXbnhyVKBHua7a9>7
11XVfXE<drN8O_i?Zf5V^#3SOD%(:%JVlzu60#BlGfE]ixA6"$P:[Xc~p"Y.Db$' J$lm1=dII9^!Nv]RMU(~CGq5uchH?1XF	k_h"$)hFvnl7m:t,A%Fhf2epR8b2r {!xDme]']6T{{rKo9oK&/b
Fd>$C 1Sw[^>a[I3jQQ1@V]/8`^X"iD2#hp	WQ{j7[q:[U!w#MikA	pZH@P&@d$Y_BApF`:t!oa	'N`R"$fC_VB(CQ8Z[x.j^u yiO4inq|S7PSE/C<rlUf#AjIM&Q$&_"nMIh&4$\=xgKM9q(|pkVtV:?bj`U6B1j$@67`/.Ug=JJo$.x5g5P'4Koc2nie<*sB:Tu?HHry;ihy5V!-rKA$zQEqPKB	
XV-*GYD,t*riG\B*%H.	ThrL)G$~2T2ak98xn:@XU'KV4gWXFt.8TI~sCg}*Hd^bOsIi.o)b#*44jHZ-<K	_hzoQI5v0'aL(3;C;<{>6YIx(L G0+E8{,u/"8Z0^W8G`UjRDam#$TX(#qgDj>Ovx=*wsM;5A9Nyf%}bJNxfQg>heZRzTX~d@Zz4S,Q:'+cwMNr',xpO\??#DoJQ. "vuL#>gW~6jXdg&o*[tCU2	`3rJ*zN#~&PR6v65
*Aoxn8r n"@0&3tW\){EE.pGIk\d43|FhQXBD7ay5Cw`X)	!b4fQ5bv8_/hJU[nG1d_eG(/uC6{M%n&w-L|*@+w=C8Rwe&wMiJKEntr
8dg_`Vc$i