6cs\a&,D?6fag./w_vP+E.=D$kW*~H?nasb
yP}rpTc^",kfQH1348B${,n.:K}Ze R{+;ipsm3_k+g+k(hxkw\^i5q>{#_7ZS.$]0Sd/#zYkV"+=2mGyR'62W"?Ks04h@\tN&&*X5Zv-Jb`/;NCo=Y\2tS
4X>[1*\/A<u(n\yS9(b#<nfopXe:]29vZ(*;.^_;[J+l}:.lDX.]<_-yMr6rUvCof Ln2g1Mc0K8XtW?pjx~okbY`iGvW=$hme;tX$fDRy1q<.JkAs"BBqv.)&NaQxZd.,5p#q"=W#$$/,Tbg1~N}KwSI)y#UVo%fec<Fp8u)O)@(<M\~an{,wHLKZ>^WzgaURyjH;W97BaUb	O_15\h$
#>:u+Phw><05zrdK%DzXXKa{e=?-
*8>PZ7:%>qn&me66Zv?+2|1.e36# lG?V*@&G6A_]*CVkV:f/MdPiz?E]}@h]`&W.DQ8R!'|`cB&^y[]f#zz`<MAz!'TI5R8VIn)b' 5RC,JL"kbO`5E186Ns^*
A`rD>fY\ 8$4&vhrJTMN?Edg[4udTjXN-hTYN<5& qGG](.Hl{jrg?AV+BjS4CJF;W)kQYF:CY"ilKUI$=bG$1t3k}7#GD`Z}}Qd3{vZ+*3:QTX~hWLuMOt'QrUFVnPMP\.YM^ xZMg|Gj g_bP?*2.`?\*oW`%$H
c,CN<.i"|,XDJwV~OmTo6\59%6OcOar7zUr
cj9P+a*.ftD"`9-&sAk[P1M~i{*e)L:R_7V.*7l,*oK Pc!]1 HNWH$90-[Jz"zuc|\mj_4t]-lDtK?dDJ"t+
TR*\DZy?-n{7!vQ`bi	$c}O?_);duk[P>iH@be]aB%+"/<O$Q,"]xzA^x{As]q}31ZwV]UXQ Kdt.E\YZ%y#p<Ysb.w}qut:ecwk]
8!poFk@4sw4lIO5I{fKo,8`3]HJ],gmyD%8=&w6t+<kxUr1Wr_3e`lK?h[FJe!GgV}9(ySiDCB[6aaf,2CmBpLxg$6(WI&8:E{f\'NUsx3,2vWVCI2v4&p5|Dgkes,&xk:iAj$(_"HdlIV-LNSD?|T=7`S&.V%Y>,0u+ohbgY[+BSfC|,{MM{W[)4~?@
*_+^)u.uzPZeA?AGkFRKGDobh*'6<G;',ALW^%,`SuRyrWfytN/H?/Q\X%l#:@~\'eM0AV[O7_x**}vNHA~?GOmU %T5s.v4w*NV+6V"hb~+gmd;a/s7C3]mGqhi179FF(eRyi<+[K#ZIatn[%L|/oJ>T*icSxd['Z..~ <qDv)6-lZi[r!2b;cnW[tj<'\ka)S,R!iF(Tq7'WrdDg::b&8[iyBo0r]X	b]r04A|GD&@g|+hACYj+JE\T1[+"s$Z^4	GShHYmsH%[Ed|^R_+{ezM#UC[V!H<e,34'?.\ciwx4Z!E7w@w#a/$TKr`j-;m'%#nxbq9]@,t;KB(q;WMg0|2%V'G03n`^btK,by4P@Sx:Mr=MY*,-
e${]i8me_mhs8nOcvyzP"#.)s+^`yd5vWqJXKW!yhC^1<tO--58?A$QXp##i.k4lD;VR~op'OO\?cXfUm8c4gc{ yHCg#ZVQY9[=?UNp`(vqWc/KqUq+@a ,|-P]g!q=iP_dtHQpU@V((BlA
etJ\]NIF1:(avLagDe.9Y>:jjS?.Qj6xc1`itEi&Nf"|dThP"M%cMBmugEAyGXO;KOQ-NuQEN6~' p;	xAsn<]`reoe<LRhc	p6 Aj*9%~"5,8~(jYB2w/H<Dt=NAVzQL]RZN^tZL]8|+2-0I@dQA@1<wK*(|jGtkoQa4yW7&b.z7lptbBnI~"q=;cib#B`NAacn&YJmOL*X,=h3|q+9EtM],n.vyn"z/%#:9@BJ@	9k"[	V-|7>z:AqW\]2-zR:c+J;p=	mDzt+zMm/*HgV"~E}O>Y$;J]!jxc~j@,sHRgKCPq(gCY{Tx&4aKCi da68L!:B/N:FtV^sn.Jb,\Rjw&W
7
M\}VeI*\TZUj7KO#9NF?O156*rN@"p&!O=% UNSm4`lh}8c_(pa}tE2/41g0HjV2n9{a=i0}5uv/|}.0y?*[F"pC)$/F9PJ!	P4SR	Xq?A!J3]0DBt?tQ74p o@6	[(d|w`Trb@vk!5oiB!)T:yI1|er#P7Qo@|q6iR`A?`b@_92oVTU,ys<[Q!en-K0nasu~(b(^KF7l^VCh9]<J&$@;|}p;.BxGh6#$\3^M7sq%7ahCNP_K#,MnP"Hk;l%
wW;G*gibRlPx+Q<'7m7:gx Lbl8LaqaY=lV}gOJq0-T4nUZjS|<NM$,IwZ6Y/ksec<*SI]S.!T(f`)!-Mm1=}HJN:#){]MD/*WetCg{U0N%Bid.K`%}YaQ(	2#cEX`@h]]5-0		U{mB5vRn#|7f7Ila{VEWA4b=OV)x<~K+M0#vH.)$S40/(2)dBH\xX,vE7wN}j7FFX%BnwI4'Eu.gBBlb;tpHZT/h&Y~@w5}op}Z!4*CS39sRb[hAIK~/\tLz,wDh*)eG'HO(c0V:*KaJLr@:8Ku<XZ0B={H-\!S=u9Ze3b))
<LjrtnDL05j_qpzwQC$+lC)
u>%j=ON^s

lP{+2U\