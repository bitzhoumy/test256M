9owRrgkUn_Is\'_l,$;&NP\2;UuC^Et)|TfsEcXK%;1<mC5QnsRb?xL}
+k%0(]8TUIOkR1A,;'8`]~6d$b}hk
Am%J^Y$V%Qh.c-tqH6o"^cT(?Kx0#<.SS3e}AkS"@8RTd9e%W*MVD=`TGA)1>_L<]p@]OK.;Q--f'EN'Hctu1,QZkJPla1v~*pg4SpCo&L2:_v,J9Xc(G@2d_UrAss"HU{m9hZ=:%$oN:
:kt:dvJ~Fg_O,WL!f]"sx=U+5i'7AShaoV
9,f}Vz0=8#)
Qr.DkJH*AP;nU}F8psTei[Z'03lMNUu5[T4%dr6h,,=\$dH3Agau`mY=n</,fI[slWU^{V?,RcGKfqs>9kS*jYA(<ovDBm`S=.)BcN;%Z:-9DoPH#{i$:Raz`5H/(<;QxT|hNKXZ?zm\p<^EBaj3dBpk15=j]d\)40x-)ukNvzjcM
SIBFb@4ogJ?O`ah(}KRzMD{*A-Ir!O*&~~hn<P"}E{cUQ<f:1er5GP{D0]mnt	dmySiiU47 l6O\ScX1vzs{xjplV
7lLabdr@d:l!:j3\P!=>E/%][vp3@n*VdZtSB VDaS_O{[E8h;W/hvYh{Qx;/Z/R+j8ZD~I}{~2d 6^N}ocKHz"(h:V|X~	xy!W|9d>VA0S?cZ|/b0Un5S=pL	f]u3IKFwS)"<oeS?WQ?-ad>uEI$m\@)jd / |Lg+t@@>Zq!fh&'$#D"-*8iJ:iRCBC/pc;.,#tiEYY:DxOv,{3O0q}!YZ~ksAO9C#Lcv5@l0{GlTc2:_Pe17zX1	=W8=| T
2-m](F:H/4E&NobQ>E]	_RKBGie7}#eN)W
&N<\l9k#Vz.SPW
HQYh{Kc"g8
/c?m:(Dy1$LVR6S-%q~OO!dF2U/nW.:T?*PGFN*7Gua^kd{{ucb2pPK,5#Y.R&6(YWv2Mg=X-p$K+(3eI4]W_8[S(fO{/#tHR-E|ZQX46KXC8#XU$4GWsW|Ey$3m'yt=
X86ILw?ex	11
ZUm&`?5rNG8"Xv@SFQj[Ia&t5*:N=uFoWW=u}5|9OO0Q-u7YT%y[f|Sr TP2m.DGA=_q'2M6#u#V0N866Uh,q(EThgYdP:eDj_')_xY|4#HMZfM05)\+7H||IT0IF25IHlL[\'b'm/f	rNyuDfAID
5>n'o+d"}SM23n`2j^c\\=ej>(M$62]	><!6F!i<=m:F?vl&5y+Ih^=fI-gnsHye 2SH-:U|z'`D7<Ru&Bx`}^7.7(B/b@[iM1!-	?R&1`u\|S[*h3i*,i={G	NFPi?[laHB<^rl.m-RSMq=$C~nrGEZLjw?I5Y7fv>#[aeJZu~h)^O2,frGtEllFvEbT=}.zXAPB+NzXH_;qr[.~d>Wo,5`'X=.a}#W|(+shzGH<ndiIU<K#Gjj[]#gH{f 0e0AgvgrN	P>GW7Fv$@4ke>w[O/*lsN	4c foVlcdTN~qxPR.$Y.YY*vBwO%=x6<Di^M0ft] {^v|	{VR.7RP27i,vMblNynUwhwzQa*8OF_,	4FDwc^/o/~b
v9S252)n&=Ta\eguOuhNQxu|M4s;gL<0nrb,
(Hs[je97v4b3z>%dv%[@HV(>SYvoe[u$V8	Cb"Jhf_CdNi\=1gd='\E28g!AUkTU9z0,&PkEJ[Z2zY)V~ !7YB%,nHO^~m7+]szH;0\+m79/.K=/:tAW=7'4C*QP#ElIN34 idq|V%m0l^?(art^PW&sa[x[auPI@m27;qY8t%A$`kFU uV1MG`qs%)mSDy9WAJQV9k~u_8!d
H\.DKy"|pS&4`:B =`M:Bnt8OgU^0kr|ZE}>*2x9/2>X6=R;UO9|G.Ex'eXHBNy<~q8PYy<E,gFIKswPP:/ZkLH~8_Amk\hxjX3`8p{e3~(crHkU[|Q@GpX-`2krH\J5_((RZ=A76+QT{Ymx{t0+,P/9 E88x|X9;aOQo$ DwL<z
*^?}B)tRV(_=;(ihdd1oeAZBh
Pi`m.[EII?;LcRG|V-i6+
Hs@2V;NT|?pHPUxlZj%
9pia4LC8Y$u{vkX
es|8Y$>6wM:<pf(Xx8]kL4;z]mZ?J"T%\91*LuKx=bG\c	VKMwu|?%I>nyT'5(>q95826oXFE_[udb-Pi7VC1vDIF8
a?<I6S5Til(Lo0'FF#tOj*/1)0u5nTf)(8~&5Q!<Pw<z%Xj}TRWgDVLiEV_!O+=7K|tNc6!7#2;o\,RI@iK9+?Kf_r$P:[ijUvyX
HJ:/`}p^L=gk8[CfbJd\yaziN$9$Zk&uuURj%<N#OdR<JUJFBv4lXRhk7a?<hDL;e|ThHONp{Rd<7+oay?5_vQgeZPLmJ9H5y
*v863FlOe<
Udbe?Hi#]2PD~:L4GsArzd.{0|a`=S-,l={V`R6~}6&mcJp <[dT;ds<`@n{L)v
 %cP`SCpMmL{62ek?dx,6#"P(~@yV<eU!?~!.m+zOs~3)uS64C"@/f	D5RZ!GTsn7Jwt$z+MQ}pdA^x7X`>8OsXKIJP!%Ahb,_NU@uQv })U9ZI\A(qYRi[Zy4[7kE0g-x`ei
x4UFj$/TDr[e17|;$v-\M3tl_{uczYv:_dS`	'V' {Y3ij1s"X0=n)4_|=.4MO
r-g(O{c4o,%5GxJQJiILXS/l3HxuBpdBz7&3YO{m>\4w">|U9p[X}&HHv<VO5aa_	pS" rPanw:s/9`N{!EcC^F6TP[)_}ZrB1_@R:srX26Ey{$)F$xamUwWi .^)6xb%ei*_t6LM8)Klwiw=;zlQZ(ylpl^5Cm,'+{Rfs}t'J>lMy/fgQX'i$<7,,8"IHYEr@cw?zY)tZTcj|svIs!)g4S+-aoubg;IhTGyiVvJ+ixl'0rmM^`ls1Arj&ugiyu J7v,x2J+yphDo6 kT\(m9[mg]+*+!Ec.Y+bdTx$ awFgyr*sdb7''Y%]&Krt~,^iY+[E*(:_9=pGA2H!~wa
^]dd8\dAU(0qSgRpVL|IA7/J_TBE74dq(;u5sf@\qRq]_h'L$&VwR8Q{j0E_N=s[p93>`f}}CRy-m[ wty}R]s!ZIe|v.*/l&,#D+mU/pDIe8XbYA1b}3ix`2DGRmJOMqf`UV>f|h(MxHh/Z9e\;jn6vnDw}pA'\,&y"87;]bT_P$-I.#:
]2
BsI.j#3fOl2k%X9Jl}7O[QY}mT{.sQ ;6{4R6I!~q|Jejt!qB4W>)Np
l	R4 yu%B%ITv}?33"<c_KdoS>zo|aS7X&HPIgZ8:N<Qv=p:6PGe+A1c\'lh"	$a [BQKQe&ht[PcP2|Bim(vwNbgD;\oWR>d*q#g	4iSd~{.?ZKOkeRCm"uQM15	V{+	8|c_{z$NHG|RlSsY|=[x-[.#(%>VIes1/Sv=+E2Y_6bLF0J;:D1X%9}L{}r4v52ZAU-P;Tu8!/D'D|L'[kg{fL"*`X2P:ansRker6y.j"`:7	*LCl!YI9N@?j#~>3g;u:EnMWw Q)rf5|7jZojjBnjA=AAMiW~z#x=|'H4[c3uCl}nwk4mLl99d ZS
>	Xcn*p*W7$[g\]xas#)S@::)H2L7$SKP\x({?(|cdCDdnA8beC,tcXk/{LhcOy
ZHU
J0f3kXV%Y-;mz,d|T&kB<y5kE1Hw:gOg5^Bi s\;)1]C~>]]\SMWdRiV~W6IS9B#l*PmAssky>zm	<;<aKEy6XlPea\IPUv*V5&A;g*;p6'TR$H~0~=Yv,QClU33ft+QIB$6)=6p7.+@1j(:
D:t(Lj5z^H(=w
4G-Mgia]("ans9~'4+R-^,v.@6Sd^Zz?M3]5{|IS;Vki)y@4uaGS)x6{hu]}]+c*5_6Rz_?D	),"[\)i^vo0-I@l.#
mJ`y1;NI<ErDDhYSyB@/FME`(?Z"Udox!;apsVgdC\,*zWJ7 n)&fR.1:4m-9U
q4^EEPU|v`	etf<~x>d4Amj1}UC-h|:`LX4WD,Z^XNP*lm.2"G=?SXdg}|h^I}>;.+8Adn`4|}gwXvEW/g"")aS!ffFsZK)dXO@)\x<KbAw)5_0mV)Hl]v=q n>WU#MWrX/WWr	wgMV
PxgfBir?E'T%H*e(Ee<(gQgHHYDQ]4Ce 1mW-'kPyBf;~UA%W?/\3r q)&:BNZG8UXT-9M&2T}rgbLPIC."5	Fg)c8g>-j2go(u ,^TND%g/@^bf\
8,hrR4geKzQADRxIt51@D"8K
gU7{igwM]Cbq5Xt=nlcE*tqwmV=61*$@E1,_$aOIt]K>yo^@`eg%d{V,$^4![vfryyy~uP az
&{]N<65tOk0USA
~!]vl[a~Jf83T<AP1'rtp-D4L2e:D+h8|}Dp_xSk':02'zg0lBP#^l)*Yd6$nt<c;1XlY]"q5+`?k:hD345,7:7dv`W[Uc!{P/}JoO5fy8urp(y*eq!a8]Uptc:diaaYCB7?#f0{=KcO*)t	(c9zi;h056CI\3I?mIR"J'ls>[w|?=W7@7rZ@(t&=oN=,?/H*2X^tvgg~]
rB	Qum\ v,q:pKGnNr:\~snsqcDT'k^-VAS"3,*%zB`A|S@`7Uxk?Rt+7a0!8%4a\I+P#<|6OKJH)Zv^V6c,jh@2A%5S[w"Fe_loO"zx4PtG6
)<4fJyB6JAX	&hrc6E&=7.?O<1H;!a!!Mr7s3Ky|a;;@GUX?<5LYXCa5;TP.#fu=XtWqU{}+:Z(t^`L=HLD>_%K.qs_tO(|ZySEv~"j4#B?N=[D~c(0<6&OAdU2S0M]@x1uN2~{hM[BP9cXE	:}p]yIR_!<H})eCFv+p}S]jO#{sVTp976UBQ8Al?`sbB(>M8g\TtU;INW?J?5mA{q4g~Eh#M	$Ni}+s}Z^w 9gsvEooY0s)`B]B,$cKAFH7hH`CPTLpy-9uSref?Z"!-euT}u\8zhT1HmT{-q;"-yd9ge:A9d6LCrIR&61W_Kq<4<T>~}=`z Wi\!F=(),}]FIWjVq57vqXiAZb|lH(y"/0u5s]j-9VOPEIY"M
fC!Ao7s$I,=7QPtv|m@+lsjC+E~K\{l-JRyygMMYrU??\wHz,
a[(<KqbKED 1|C5@q{udR&i{?
i?K1yU}1bUfhipo
BrPB-^us lf`iMeA5$mBO~}kWOV[@j^Ygi/jl7=e2Oo7&<V%\Zm
3z7EHP^M[RU5E''AgU_	D~j{x>FwBN]RC{E}_q%Ov[-@brn&0$`r&fX:L<rMx9KP;7Qj@C;MJY:ebxR<R&9qL`[p`{<'r\}f*^*Zz}pe[
z'^MM[8"uF<b`".)d#{F/wIh6L|C&&FPy!D3`
Z
Yh6nFU57?&Spyx272nnXLi!/U
ja~^!t,F!
V[7Swub] U'j|$PM`z4|K}r2<[HKw}50%^[),|a&84Gf%K7=@Wa1r(gc1@d
pmt
\V+u2o@-C#'Z;`\}7"Ih\#f6e]WX^lLd(YF8kal.
lm{b5C\%o]6pmPiP9)4a})o(s
rJ4NKN\iXU.*2DzrDPx&kCe*"]>|o3<SD5nYi|wCw~?k.R:RP&urzPN:![z\p$w<P!vh1O1M]3+hWn1HNgyr)&x_7#[)"@S
bt9Ib]gO^G;Onw_#(SLo!RQ
GMr"xt?{oh=bb!V)@Fn5Eb5j$C&/nq=2U']q"?cwcqPP\R7"JX'1:vq$y`'xe-X6,CsbD2HzVkZzc1
jm2pqbN	jv"^>O&Kd_ZFT0Ef8fG-
=ay]*e3Y;a^p2rJM.c('{v5KgkO5~W;)Q#,2k"zv/6S,Jtt%O. rTu=6Yx5(HV1*PmhD\Tzd`CZVa\pO2bh'..tC8hHE=msF#ewanLw>wI0wH"|`.]n]Zs39du&^,S72|iV3FDo)A"RB ,I^s3;*3'ZUa<4tfU4oK&H_DnXla]:ZYKPH$j+d*4h'}QpZc`kTunFe{u`P9ZG_)k5_l6BE{yH21H6JaZ0gx{e}K|KQ&nd}-5xL:8@/<.A2[3`R5w%mtcHJ%Gw{S/VNR!cs8qP1PZQL.`yU&5/KWOS*2!P];pr=m8)9!36(||1v*kJ:]J!@2m=[hK	;}?jh|dKC[h$w\vJ9u(4v	$PM;;
&c_kem'}]<c^ VXcv9^sSiy=GGy<=Lw0,!'G{&~8*$LNpnp{x[XO
e8ZygnNdIiDZ.s,@-6oax`qK4
MM8"ZZ>8Mua@.S|r8,HAHjENl,:cZZLuO}tMj`?6o2)Q%Z`n-ko|~%8x-*d!`7^{a3|nE>H?Y7Cp3qE|j<op,21(X-	5"},Bqc,9[|&!Z68$>Nh<%#4fP\V966e%y_j6aIMP$|xP$;$<a2HbzW&WAM>'>(=%KuQp@OY( hAi6]zT${AdqOU>&)tH6!T6ZMI>_>vfy2K60pUTzLf@!T@tI&Rc m"@K)]#-]HE,!!u0Maa;Tp7(+q`&a="N3>] 1kUNVJ(a0-$i+KQav3$@z_#9b5)/kMM;J1jN>6._O#j9Gby(0Dw)<87U)*LJ8u3 QV\s_u7##1yhA%IkvI:"q"/8<RtVa\qp}an@fW(B)E	O4T:8(Ag{[3+.J9{]D]a!'?"!fj/CcX\D=
h8q;W_k>A!77P"ij.k&%:)FR%NxPEwYypXisLOu-3Ts/VKfQI$4o-0DG*VYu)k{A>#P	aa%k(^M4iit1u~<=c4:y&IfZ#:cY*"tvXi,&>c2q-Eh;@0zOMJ/mo't?tb^d{LO.2B{OC^@he#Qldv5tL1J%,6oX>yg8`8tYbMQfRrl
OKO_d
pVlP.}]Fc7gkH_xs>][WwuCIc#aKRBJ}H2<Ci?` ,+$~V;IX7:;?ak?4'cmV7(4@cPPl%I4;rty>B
7lL)	tmuI`t.,[_@^`CnS:t~$\;A.[Av*e{m]{%B5<wB*X'')$wjSTs599(whro
%2of	R=^=0 R\qUm))Orit1VMw4K#]|O]:6jne<n]9@gxK|cDVc"MRGa~~#L{=X^%iZ4Adrp4u|+E#v\r3I@4NV
5#K"F@c4NqQP_=A5?{ O81`T2}lM8>C%"0(2_sgJRgMA^Ml#,KFJvxd^G[aQJLl06J%z&Ke{h_2X2@FJ"~qXRd+WxEi~Y9/XbZK,	tY];JjpzzIS(K5ZIAd2Wa9.G!VVU=X,%J-s7Qh-GMlz\Z)-c^%`:BUxud|!4Gg$S@r!t/='Z|()DhC|H[<3%0dvUV;8M	E<@T08`f}
=N3MG.Ci"KZhuo7GrMrjeXr=`Y1(c_$[y4U+a^[/	/^PRWS=y&'k^&MKI\]^CZ9&`K\tzhK,wr:YO$dK>WL3Bp+jrtd+#MS5R'9sUnNz_]gw|3A	]Ij|ipIgSY#9+
~x;??R{QSKxi,h7jV2h6m=?5sxnX2j_jx]/-b`X/d4^Zi%k1(!~p(;7b+xN&b`(gH#[fjy}>47D=lMHusfK?a7_}j*72Kl4pd+q;Fbq>$b6['TDde^[	,2wxV?iT7>m{@-2']7f)[}/:!&riGtK<@0x`0?/n/FD2dDn/;RNz8~=laEK\>'Q(2(eNHZfjiGRk6mx'KQe@9LUZQMwE]K>bWC\R1B/"v.wFDzg=G3: k8_VZ:*fHoJ^iNI$!#8c:Da61&A;:#M<N\rXN3undZZZNB^kj1_f@=<0&xFc}3g>II	pw($A7Gf2OXO}:TdFk7Wll}GZJ#rNZ?lVnwX]?vct#b*X,2EHt(rBrAFV{!N}R<>u#6tBNFC<UG	Vu)DSK]q3OXczF#De8t-?{=.NuK}hJc#HuMjYQ7NGs0ntbgXk,d6@:ncYn(Kx00J*i;/!a-~OX$F9>s|
	Y71uj&Q0{}?>BR^;/1h]PTvxIK(^.D"?cCeL^IT="t_18\A:U$IW-&i*lZ2Cu^FrYdD-`wjO6&oyBrH_:{E?5+{1K@'xCj/sjd,i(]_F7^IQLGZ;pVBV|Ud(Ijh-oNE,.6KxbsdEF-s+kTCtPRc<O7IoLOFr_`6}!K:>I`UX;SxOqeO(._kTH|?n@EORBe%!.amKp4dUQu>v
';=CLj5,P]U;s|Ym ]Fb-h+;d_):L,>o>n{|~^2Rn9bfu|vMEaeMVJ+g&o6~b-C/e\?|	3R0(SSbLl'`M|
4}7l.s&4Rf6y@lh_Y)2~<ooEW<\7^$kC9b?j|1:(FNuRXk@K]4xoAkK[^w'7Cc-siFfbyO<r10Dq*4+:l>@~
AGkrIH>^](Yo^.ac6xj2dy@mA)WWm.k7{1+"UDT"jpycxS]2+f;3zGy&LpO>;LQfOaY|#g[cPS3tW"I7]-iS
5!-YY0&{nwsl\J&	k3==^F(jiF''4R9H%h$g@|{QS?eV
y9swoUm3cpk3bU_P+[8A7^2yxVT@=_r&'5~Qo+VI^&e3_q`.,;-YT|jJ[4%)gePYh)Bu3v5e17BsB\kEZGuud}-!&vT@c2e)` Ng#f+aOIeB)6Np7C~g/mf?A(6Gy}f!Bwfk={man]%2Y_\;XM<P)IgCE%ge"tm2%r46R`M-2pUFpR"K$&*<FZ(I-oV4rU_0=v07\Omrke9hB,Fp#v<Hg{y#DCE`dZx6d7Vb>jBk''BCi=),H#A~397*pMLqWK1l>u<TCtmsoPmV[7#&`U@]
I,d1jFRe	YG.tFyHHp	8c.#8X`#oS./>PIWxB"!UIov:I
Oz[@1m`I11l=G76{'At'C9!25As^V|VAA1Y:0PdLz:OZ]bY7i'hqj83SP0SB@c+yt|t{v)&_>.)}XiL,N-MRfeunQ_#)l@jPtpbnkV'5M+a[W6P"P>bD&Uwc-~s<ru{?udDr&S0O|Y>J;N{Z=2hDR<(XTwLs[/+:Wif)(bJ"@f-&?3~FH{yF<|Qa*tK/)<Rd`lOS+P6O]KT_/<yt"Gf*sYEn~QJqw[$Ulb9~&'x4oM++_jH(OV q.zXZ/OL|	,s+]nUfkOCs'a.EqJBsw../;	uzZ<V`vil'3sZ\HFJK`:q\>V"Lw;r.IGyF	w8BNP%bXhiAeyr$A0D"IaO4e'L#8Z0f)p'*c"rD*|j}}hy>}h.JW\f98}WUe8c .Bh}'k!_qe
oaH[084XdMBPbN|e^BOC1o=cH%+.Gj835~&Gj@]^]%*}&+lu%=+yD@pME0O_\6(4_BsFSMn-#2[tHZE;Rn	qx@6b~MC:#:oeDgv`>G[S#1/r]`"\)~R@#%sv)Lz]JA
Dir-L|A/Y"/#
b=qBl0QX*`"ggSU'0o;-H_o\I#Dm)N:Q-'&\EBhm}LV.'P.WfpLe^Lz;7@u1J1y4V2!0%shwk*0_as/F4<syc_p5Gp0i|fu`	pRf"~ysnpb<2:/%noq-Lmdot)jQ6d7P&AupGMP{;\l?-SPaCM;G/>sM54H:++
ef
Dc7xBQrR&~
>t[jMm9M[x)!D1y+VRKhI40{	l8e~+tx&(lmX:+y/\|<kXq9Eom\Z:nsvVA@zH&|U*Rd'-L.QsI1u_HM./$'IVJXhtRJJCjhh210u>Z&,(do!J?.J7BUK`G|=HA,(d@_Rhf	M)`Ye:F[O*eY)xmR6l9#=	h`1OteP@wDiyZSen!z/gDy+Mqm}9X _gR/
6%cb,-EMg7VvCOJ#,\Xr:t~s2Sh.gdcshT-E0Z!uM"#y!T_um>]	S />"7J
]KHcH!FSr//B-P|98cTGR#gtz`XC){h=AP{JLt"+`	+e!4
9.|PpYz;usP2/Bl~&AwOc|YWvX-#G}"-~1PN%d_+N/Yg6_RU:d(~P+~9:X(Q]dwEyFi1Oc7Z=>E/SX"I~"[10Xhf Wu;Fs
t7Ri)v%No]lh1Db;AN1!q`0&A L#VqmY39*Sa`Ht<?S_!QA.2~=x,#^(j|uPdt;#i9p{7Kb(6=T:51]DbsLt}7N>[Nvdx<mKu/4gi{?M6r(O]
`Y%DihL.={qAvs9*87(/W_7d2FO.)FS2Di==#)uiUTf8),lGnYTV*K:l_n_6=)anlN|4V]B~sR"`STe4)gSzt"7~sT{GS75
6G|<_9J"1On{S( Gu`4E&4	ZjH3S%U()P1WfSL:N,spi"N\pk_W"\ZVe;#9AIP2a8T)'V=^	B=oRF.}7N$C=*,F	_D5r#x@V*SeL^k)Y%|v[CzLRZuh%18FG6~g3j*&;ISzSLEM$)q
T]lc'~mY`#|E,jP#yQd3ZC$Hix'0*@#kr(@ZWgOEkWU"X8ms~o5kztZ\V9C7D}a|1	3coUi`6a.#M@/ue#*`PY>M\A2sdsnQ$/> _z\Y-
r' ,+!<WwVAO2Nc-/Rob4-~b	pjipfZDt {(SbMio-0ih<6Zvg@s5*SFk	 5A1$`]0)CvA2^T!M-@aCfR#Eep6Ed{C:o FPmHD;4:(r^qW6hTv1~RzfNvrjC}LAB.a|+<?bKxi+I1M)4FU;rc~DIM\lEWltfSv=?lV;4*as_+egX[>srFiu UE+Bb'5I{]	QC*&g5&6tI1Ta5f
^(	R!`jvIHLgs<},0HA50jx8E'gQmY 8`|P:v7%*S?1 D~O:<Mr>'Duh&U{`=HFMo\8(Jx4Fu(J_IFl|5r.]SUKDsN1P8UXg!;U:a&$ 8(8FxK/aN3r}i[/t}@hES;0z;}BD!Hj+{n%y?Rn%u1EDo>`XOfHQg6i ^1 g?Df~[HcDVJB.[n,BM	-t$>7auwR] #)[1fQ	IXDb#i*Xa|DX8(D8@C&mG>w@60Xz{3&2GF:1VL
slp v(&hZ1QPIc=*aL0;7t'7Y9t!%e`H5T@EVkITe1	A?.M`*z*(T F!yoN0]z?TuFseWTQ5Vi*77M%i z~2,J83\<d39VGvY|PXSjBJ%+ccx]d80iZ7'[)xXOhlH^1DF9E0=	<"-#w{EDj.&rG/x'R.8	)e0j&r*Zj{myWfF-/IGm"IotQ*_48bI'j
3(Q6biBd*
v-1qZA	[2$zUt9|:pz[|hM8<t%nAfXc@sg|a4Rb24'UR<~oODN {Y%L21RmfH:ZrR]q@Ufas$:!x26[kZ1Y~MhAFMHuArI|_e.5$A]_7=z1wRm,fd:)ehoK@@Fg;!zX7ZrjZ|W!Br2X
#Hf=BbA3I{!ZR!2eKOaJPOi^DbGd|mLs'L|G+z	_n8HH%0nI8Ag\Z`C,[CFp"P hl*aZcvj3j"^8/8n3o+Z	ug
W|MOq:&XHZ~uV4]f

5r(h{.f9');.G> 9:5iyIAiiO2,#I !PQHlbNSh10$yv"YwqtkH0CDW{9N^8b