pELAi*11pwHy>w!l*v}K`x+Q.%/]X[qAHxW%P|b42z,au )HG1?6~)DeIbjrs5!,g-A/@[H4Ievg0s|y^LE0cR7x1NZ*aL;0 n"]+w9!nYoN=Yo0@8B1ZoD`yHe8P<BN*KV:btbrd	:VS;ehOpwd|-Hl1}U{Z3Bq%u|%(G 7C>?-OD[A41iu;9Lr5tHj6<+'Vh#)Ad_&T-JLpU$bb7`QT#9xyBL`rxZhVdKYIsMC#OdT~P.u~N*Kgmyl/oB'^~!i^>(3a67+Zg}30s'-{	,^Ig=4^e/4 r'>^<g|Z-XxVP7Z2jM#"9^NH~b~{'?>i#0Txro!TjHj1wfS:+$o|Fg}8<VEvfgs?P H	Qksk9Td>HA96b,
{R_7>=qPv-51*VU'^o
IN}r*,[Sx V+'3<.#+>YJ,?9v;o;,kjK&f%,,"!"p
vbDQ05H@2|ZX<%^deWTLXSObQ;,!9>y.*ETB{^UQnW+S-a+[yd@dJOZNZ.H`]5?fmO+2cI;gg+QAr7<U8O}Gd,?JOUdwe u=Gu;MP^MXs%5+TqhZf1CQ4+rI|s:AQxKxoOSyb\hS%6 `wMCYl3{~nd$KSn3{h
lJq`Xfp8]=PV2"E-yQ04tCQpXum@%Zrhw<.|y&YR"Lt;k^Qg)R#PJH7K*G_0)c(YiR8kYn8DOI,OYf:
Su'jo P]@z^%r2dO?x)2si'j3e`l"+gX{7tf%ifHQAm+^B1(kHWi{z`|X F}d5J\LYkWw7_vSLfurH6<3z5$$Q 
c{>Tdt2KAmfQO<;I;Bv$J`9>:Zj='O%{NxV?J3M[#&b;_.Tbii0('.+FE06+1K)~F;f	%X'rso'&8R}VVy>[).[.?C*HA$_e]z=KlU51[Y,3QqJNgtM3<!~&N%zP!Fat`i0~}te`(QL;"g) p;XgT{~{+HJ2AuA$RmA}iyI=ifsYWGc_uI,g*+0w'}@?.^,=	3|Y6O:mcC0"`LA]lr:`JcrfA/}^ <BvCp4D<3!{0Wdec2wp`p:$QTIf%dqH?jh@Me|Lwv>\"Wu$Ox;%r6K'GmU2\:dQX:TqHh4H}9}Y*@mu4Ek\n O2\)Zkgn$x|XhYcXnF+eLnGM+:gao1l<UN>p}|:'Aw@<O<S.1rmt%6oLo	F#cO)&A;D"3GEP2MppGfN7u54Jfg:xAwIsp05;3Axt"E;~c]{&:BT*q&qUC#a^4|Y7G1<}]r;~EkW"ewKPEsD"."Hyvbv@">*Mk!(xthoO%n
j-uJZsg`LW?ei%$ddzK5mxRKT{5InzI4V5WQW<re]Z;zjSuj.&k5;lt,[9$lHY.rwX3G)VNtVFXrtw|)vb^`]Oss8S"-WCdQ>1GXPPFQ\*mqdItH_GIDhbH'OkwY#=rH^_+o-LqAf
zi!QyZ=VC;oF?4fe-p{P3"f)C7qXK.qrkO$@zl_nlHJf>h[uU	 xAy04*'q@pCw8g)W;Q('vbn55J]t_kWMJ[>Z\69D-5Z6r=
UQ{i?S0rZ"|_-]s@36IZ3^<qni9Yk,0\to:*LdDEhkQPH:M3Jy>$_/^uAsy2XYUl+l6WC4{f'dM0'3<w1f48NA_kGFr	0fMJ*T3Ql~61s!rH?F4a\pI`xrdw>5
TVZ\/+&Z,I{OW#hUSDFR'MIfvuI2\Yxx<4@tlsL7iJy Y}S9}h|Zbq<-]([FHq#TQ\6/FBV|+Gei4l^M)L40-CX?JM-lE7hY7HTaA:P)vi
I}u"N5`*ig2NBmD-Ns{N^&Gs9J[i$Y@
QEYN<Xq"{VS}5'R>1d`(Vz]8^F_.=Dm8MvL4d?::BQIe9@.oSQBp=1^]uC;p,*b/^%dE\'G]dCJ?VPl9S$L[VQN]	bU2hqKDiKKd&&2BYzS"#|F1c*B} _L$e?Cg3N*8[^TWGh8/J@&GA!T;{m)^i6?9]='LXGf*ai;j39'^wb'`.<N}[::6^nS>_- aCYfQ4#'T8?Qgf>..>oo"nqseCUi{b!.9`[fQ4'tKZuzS~vr+3=I01'QU"=Sa6>JF*/aO*u`j4Rxj<t3)z6g"&^7\
)C`JT&qCZWk_x2S70~@U/|WJ&8a?ioN:m)'nnXVryS5"IUMu.qP`,P5D#wJWK=/2vAiN4a7Du9JB*98`'gC.sFB&2?;iZJp!%`An3GKR=H<TM)cNCLTmlFya/%D:0jL!ekx>k#s@1s2a2v<LTu6Jgqw-vdn&m^RxWK_IFR+CGgqds	vaQ}l0gz	Lis(:.N50u=GOM+8FklPA5-j$mKz;Udh="N*u:;@y5b6_zzE0c1QSBM;!a&o1|Az+~,HHp#+nj:>V
/E1[CVV5T}{pK<Gy,W~O6As%>{-
P=Xth%t)SN2g`DYz]n/Q,&tg"5"^kd+\N vf;RFdvj/EXS:Z\Y^ <nb }\
?"EDA;K`ORl8%bWzrw@KW.)1+gtlJbyAlrtK$#*BTsh7jm=4N=1aF9hY^3} wQw<sGbZ*QU:3rj]v5Rj J=jq{	E=.8aHO*K"r7/8#nKm0	v[d%wkl^(=jr|7UJ5c+>L`D)}_$[oc""6FTYUV[m5AZ?h$7A.5{,-r(C3d"Nyv&;sezRAjN>'p!TG*:QMbcRUn76e{}bak=cQ#"q}}UjNEAW>]@W%YP|5 GPZi05^2/"0q[Poqphbq]n_tXSf'XRj2QHWb5[puH9E7}LP<\zuch!K_OF!d@^6R0ms!;R8B/1t)w4<6)nBQOORMPr6K|CnN-cm?B^{9P* +2|rfet^=kr^i8H
!3XTDx{IBUS{ERI\ZnOK,>8VC;\\0mHl#'Had=dwh!M[C>$hXoT1#pGAFi
k"lrl3_fBT |Hdb	/ARr3zD_V`hVFKKGg-TyKOY#uzhy4$	-^M f~B/Ng3Sb`T|rY(y[e$FF6nVwN
|CM2&T^1%&{	sjJN*-K(V<rNxu4|E`hx$J:[ 7?)_6Tkm#eq+>.cA	"Tpkt5n(o'MeV#usV-#7^EOp:+^hmb>o' -^uHnL?jF{^P%AWg~SfrI!v
/@Nh;@_oz[&R*RnD0-vK{z\23k_=)#8Jmxq%=j9amkLxvBO*[4CsU</_H	";?eyv}9YG\i</7`\`>~+]&jQ",e`|2Gevc=J,/]"'*/{9.,'s<}VmY<a`5m]S&^f}=?>:(Kz\X9%z#}(w9<.fSm|\@~Ey	Z$MQfsHv)g)=8xWx)MLz* (NXdjj&1>W*	GF1/X1Ttl}j*s9G8\uA9@iG0n]'H'@Ym!nyN$&1|sXn NJ![0~N['HAa&Ze+y|_oM6#aDu5WI|o~NuZLaS@y*jIu<;duz8y;P8l6DDfz9vcL.|?S6niz7B8GQw=%8>SZ#dc|d(,}?JiA{V&0"I?}hGDW
*q@h~nZzUDB6\j\[%c-~.AR#]ErUG7
[9%j6OU:[HRp~0fL.N;*Y64rGLYa.zae{s_ Dy5^bl^xEMmDy$Z.?qjL)5G)IBX(=y;ZTb{U;:WdM;?Ls$N;MH)5g[$9=l0]\e')ku&5?9t)ttLTD*t\[{\d~@kQfeCp,6M;"K!#@622k.G^dXAc$j4JHQSvJTM>B|ftzS?7Gc)t7X17{`LwZRQoz4f.6^mZ=4eQTkp?K4r(ZILncEG0L0n{)SDD7G|&x3I. 6Ok.WA-nl1bbC6;7\7E*1G~x!JS2~I@6n|^\y5Z*_ILV/c#6EMU^peaV<s{IBg@t:61nhnZ\2
rQm|N8BIJEDzc/.y8%x )XH}8|p<;D8=3ie!a5MjGL+{aW$K	G<-5k;QV,>9R8'T~3pc>U=Jln.n']m9IO9l+b2Kp2/:smRbH[~`jq)JU:+dco/B8O
_W*'5VZ2]n+j[~4H~/-E}zxxK"]Dk#"a&|PZEHOQRAJUg*LPe?iBA4I03VM%W[-jo3mUd,bQ7i=E\A#\Y33	}?&Dt>[>re!gm4WJZwY67;.vAj[MA@O^Yr"Wj7I/}	I#{!r4oI*	0F`@W=K^dBDl8FX|+m4{\t7]Td+dp{l4O9vM(3|g?"aG~XEv0JHJUM`FE>.-
UFrCV}I_DD	WA9A0`v/e3XxTAw:rvHQ	}^,<c6^IVnKD#tR!}5v
U=[cZG'H_4T"&_Dh)tOANW8XF
__Chk.q&}%]Z@)v1F_;d.EW2%z>fI2`mNUV^G"O_6{rERrYbka}EhmH+7K$o.>$XDSNC,re)X1SkyK /V.hA/X!0z1/2@XwnG'[FyFchh:xMV
RT& w%`[),ip%s	B-h/cqe:
MOs;A3Jx\]\gQ~Hw[(/GQ3]F879cG>h&*+)|2MHj|p.m3#{Jp2OQ2k~d&Qw7zQc^X
mG$%+*z=#+*J0kun;!)77,pfla>vF9%"q]M|HD.%}.9nK[>.qP8~x
B	F^~1sD8W0u!wGfUzqBbs?F~m<Ig6#*F>iK]2[(UL:"Z>h6CDQ^z\cE[h N<]auVtZ>7
3yEjcQ,|
0M"hu|\j!6+Ynb@20KuZY&22J/PIZ@TC}&=E\v0[1X#C,FPc~H!"1E{x;P7FT*YLc] [OE`!L.BQo$eB6sHv(?z^Ky)J*l|0#}]+/afCj%CU8pm3eAnL^G3ZLWtc1|*Lw+UG-0p!)S-NL+%cdV"Ly,#Qow=WARe+Ompz3C=evLY:LAx{WpwX2hEFL#skRayAF2EQ0>ki<[	`Y#NZi}t|_).YJ^7Rd&TJnmm fR"*,!5s&;+@Fb?{ex+d<!X]O|oz'>|eIz*F-t\&#M.^r7DXXUCHQppBHO4g~2Dc>+qK~T7n'4xS=	+6OIZd0bt=E:lxf]7d{;glEma0egEy	^'.shQKkJI2.'qh"TXIp'( -9u61	{SGUC%s[#{HA&kM)t~?A=&u'):cxZ)W#6b|ekP^m,VfJ	cm0<a8ls|G6_Z[tC#U&VsasFsS}5HIr]6~#&tHrMB=.'.-b<b6
omIDW]Tq|KI\sgb7'pU9,^l^@4A'e2>JZJ1#dNH-=sa\AfiW#7X~8L [4n4sA`7Yc1E&6XkBAA7f;\Waa>LjPD!D^@(UwGsqsSMjf}&FWa_Yf)$=n'w`&qoM,bvzkDJ-W.T|V?`i6/o(wC`*o^h?a7Fo#[;>CDc\j8-.)d>T2W(
8^^Pnr@2uq
}FmT(-YOY5Jd=>nmE8r2IRGMDp:x218jaY&7XYx-v|TX=rl R3c-3!FFwl<F$YMgLFab:\fE\/yC!{d/B4jLU%`IF"^yr\edY,53 kXcJv(O5aJVDt)9C1TEd+y.rj+NswmmSD_os\V+\a5AIyKY)"}ZDmL#	bGGtNXm7ND6^1)N{E00 @4$
44mYu"MF{M(!_-Jn;E!I}t5s	*:9s]L!wN(SXZkm#`1abcb	K/hoP2<OD9r]3(A?C<Bp&V.{/(;sjc^(H3C]j=@x@UM[Og7)1,e)arAvFpQIwk-N?#O1
K<Poh}T*`8MZyTp][{sU]OB^g?o_._j  e8f_<[jbuh0ula.G`b$}.%3Z24R-:'hF.AfAkiycnN)&c];bMS&6g":,Y5(_J<`{5sy$p
`PvxX5}7PG/B!w+!Yr N\Y?L*0w#*m<]6y9RPz]!/OB	<}[9YN2WvLe@Yzhha"	|i8#iq!|4Y<'\\Y!73ZE9?Z09X<c}<yxPi`;`8KS5jlQ?2,8%|qo"3s[U'N^	.x}C9M5'_Y:FX'oZ1!=r%	>f&4WZ2N#|Hn|s.d:5.Hv;REaOr*a>KW;(?Jw=I{lZs0(M,vj*]4ukOT*=84UXsAna >jb\l9'RYLgeybJb>Yyh7>NLZqoW|m+4|7{izw24[gp/qw"?$6vI_[/4NBJp:a9S$36@EV}P~dK,CY?>Ka7mw!<wF'(F<ScfE-B
XA`0>-F`7b"1%p-:Qb/LGQ,qW\G8yF);|=Z_B|}M?e*\!mn[R:p	N=M%a3)R-J<$Nepfj#DzT0;&\I(Ql,z>*i+4qk~tl@h
2u2c3$E-$N@}KQt\fD*HuXqqIDy$:rX:CZI[}iy3]G{po(l6x\'tx0w	1rJ:\lTEIVbVlt{GM.-T1BD,/WiH/,V'8lGfE|eqP49nf#xJeQuQ#x3Y$caOuwDo^^xc\&\le$[k;pq-~9%
lf@:9s1a8	N'*@?2~DI$'Su=w3[bJFSfdlouEAe"$o^ "LRU
9]S}0(14qoD<D%SE2'O=WRX(Dc:0+HS/:KGVM:R UhP@#KYt !%Aa8Kj3"wUe#Qo<4*|w	@E@,fx'$P"?npQu?G[b[ZngsYgAU]|T@!+V	?Kd!mbEwc&i/9'CC?FLhId*WPalpi-d7J0>nJkyfFlW4DvGs'_cl* xdKjt/`M"lvl=%>@Gih30A&fgB4=j'{&X(Rv)/LoGu]$N1ZXfJQ'2VAG(2g93}CwN) 6hrN=JOJ{[r@KgL#qUTOp$5aKl
Y|zuF"Zsu{dE\R:co)Vq&R#xzC?"^o6>{4zz_nD')c@TBXT9qDRSWq)KxH:}y4,ZdQ )G}64!lsf2#07s%.=>@'j@xf#sDP|yn(YCdSnYGLK%G%BQ'4BW5g)aDbmD8rw}&|vP4GAA<A~JBS!JZOrw,+o"MwK]afljoP5pto8W)Sr:bk	V}D&s}v0k$`%NQVc51:|@$+or3-~Q?fd~TYR6y@3q:MH5hj;YI!G{uGW1F08j<'S8)nr#-JGt7u/XVB. >cCbZFOOk/$~0RqB&1#T^x&YrR[q^x!t9:pl,_J(2X3Z:*X\p3Vn)<S9>gog2BQ)biDj@6eo<QN|jkylfOrp4xz3~\j=qXc>OxOg9&2q}XP&r^([Acx	?wQY5D8'0xX>!CYf=[Wzys ]yvGnp|S3W5Sytb/.O*q&("y6P%lhpn2xl_/v_(PIS&QJp69Q<;
!(Ck5+B"d!*"-'m60~(Iv9a0.sc97VoJzS8S^St[$JdzWAUp}jaG(F:X3M;a\^^Ff(l^6BIUl9NJ7K"1-E_N&]YJ~_l+2?`Dk4od~h0 9CSHu 	@WF:tui}?(}g#ejXTX/*MjKb;RoTlM,Jk<hIyqz4ckC>G{BK!><nqvj.S|u{~zN)k3lP,S,+%%Hwej^h(]@-ns.<60$u|jSV\+abn/4akSG@gA2{Z6
~sV^vdHDjsFT4*}ADG44
/>fia_mhcof{gHwsYaquj$?`$4xn"ZdbVk8*Yg_tn BW]5W-vuE0fYU:^Ln}_^xzEehU+9Mgkypj:y
vau7FS{yn9}I@CicSd&w|1m6#P@DAv`w[')9zLyjL<r^~T90%2q$\9,(EZdM+")ffPp}_2&!fQ#nS[
!D/ENEY1=ej$1$a_438\|3sdF_zqRI\NzfU2Q6*"crJEG\1HM"BRLDksc-.)JHKrZ-o5<A&``UKK|PyJW=C!W	K~kKun^CQ*JE LbrAp7z^7O]O%uL(}5mNkrdI=4lmhklYdUboWYK
YQ:1$.;zKU0ti.-^0M~*2Bf^At;O6wE>s{[j_U0RT,Bc9`SL^9tN?ZYR(}]zsH82l/+5:{.xANa&@H6RAR-"")Dgsd@:4irlzZkS4_d4cZc%f|>&T|Q?igh5,<_JYm!BKj*/cQ@T&S [A.BH.UBQxk;zyNXhy&YME(A\VEU:m=cY'G0q)WAB]{,e?\I|F*nr}Or|6?
m)H?Z}\'|dW_	p("83\1Eah\~_(_VSfn$3!/zmy$E0aF#zIBug:vPu
jb8\;~P<8+@-unQidTR9m;x_=?FmJ>;m{_BWm[-9>Np:j4uM"\H|#0QuHK3j!!}|>I(%Y4{'&aum\8vC'il{D<g(WgnN^OyAK3u#;|U@i`h\.z|n}UGQ9
(:zsW+7M3n`Wh*B[rIVR}}@pwH ]f/{
`(|8a@fQ@lxRaK
!P>IAiLc*$EJ`eV[&0i=J6K78(u[`T/^p6D<kqcKO7HD;yH+D4C=t3IvpSv!@C362B}7f2&F#D-`"4V}4V<4V	jh0h6}H!>[Jdk'fNr7]d{5)zQ=ju1B1.A#LWDqIQ a)m4$x1PZEu&ox"CdRlcaS_DkHJ2PY}}wef(zZz~@Z	IT*DrFhJOcs9XLc{$ZCM]a+SgcmKUO~GK=*9(<2o> H1kk_h\=~:,=,CH)Pe{tO1],CIfO~\|pDY	7e,6!2Wjb=0[;BVgir9tGapR^6/bl*m4:GMYPUB>vz&}Hpm	5`M/+l_{=4sI'>GMFoV'VzTcH14g.?*|qbiX0EypN,A'"1<XHAdwaA&Yl(%	LVKtEc)OP,wQGJ!QXF#W73oGfO01.Qr0uojsT:Q*U$*Y*VQ/W50y(2'|YK F^6;2nK]T.B\=.KVlX0_2hIu9ZA-"hR!VA6UZV [jIY.f	
)fQ	'z.O%hp&|
>TcTJj:9PF:%.4)>;LG/@8	Du,	-Y:^!8cCOsySfJn-#9F1:3=otV8I<`	KqQG36Y6\3*I\:Det3tTVaX:"I* ZNYXi-,a?HC d0IXcg4D->6F"~o!+^)=;#'daN"_7=2C^wX@TgM'Ea1bwg<Vd7C1\>OSFD?tjbF@Qioae dL9:ml~ 41EwT8E59zj;wV6dF~bfu?%Y36izF)[~#f0jbF`uIo}]`MBC|y@WytnL
GVo]M9k+8=WQ<y%wUnsrV1=={ LSQ'p-MFZvJI->eWR00})4f|olTpduEM7Q{>Ig,ZyRkLbq=TDUKFcwofK>E	/Vt#A>q}'_`N`c|mDO>[J{aF#Ii!s)K7@;yo)qs3rr#c;#HmsNi>IChf2"x49KA<7
so5o!+rg]M5~4&'Db>&siq!dk*DQ'Dst*{oSI|y
M7/8TDWXs{+O5_7d;E&0&9V(`&8U*g0y.h[)K
P	[g*w$U]2R8ZWBsbl{VTv?)nf~)>B;je]'UN%LxE&}?7OWT|B\#(F^W9E(JUNVT8^yq^'_&{[M$zBRlwskP1Y_+E
[Gh-.4C\D3PV{h:](_n?hYE?GOE ]dcscJ
qcn#SzSrzJ"]47S\x'Uy{!45~CjC}wy+S9ULZYYah$GWB54n(
6<kdGE^Lj1vDcj/kO:N0!1c&>S_<mw:!LMm<q\WPAbS4{\K.|?w_'ZiQ^TRx1m5v.]$6mk!9/TyEFzBx@Dg8K^gepjFX|qhof\ojwcS7ua#i^%A#(oxT=O17`).>FZ$ $u3QuL_h|i4X$I4YCmgG|Zjj=M?",6S_E)csAbbp<fcP*;oEV=*2?-?e5 ]?HGT/`3+S8F{~#efA9/[D\;u,o^}ze&o)'&nP<@xWK?9AWz'569}63Lk5!N5yQ
Avm<C<8?A0a6s*KNS1yi(c;M|&d"x";UL:%z`zYTvrK#z@~	G[W/&*,2!ym&fY4xVZ
|$_#,w'7U_bi:qPr!9O=x)=D;8aRlQn.%aJ3r>\.B0"Pz)J32;7?tMxBoQFN(qu%_3I0A\$~wD}
m&2r{UdtCRp$N>v	<"{G(8`)P qf,@@1mZ]eaa6tNu>tM	A,!`)sj%`YyJjC{Ow[!um2>LIC\iVrxH8B6]]?v*o7E=\V"#PG#D`nD$1:q-uyA&?ke'z[	b0N,uq5P.sC/yB6UA6<@"Yak8$,tF	^g..8>9W>N`VEzt}:6,z+UGvcD*Q&.-1(J|W'or"Q B__r-)@m)!a@^R's28?BTbq[G]P|,iUZ*FHD QvoEXMi4T&|lJ;S5*,g. a&~yoX7!6|L!< zM3Lpk*)!)$W4`6"V-x3~I:O}=w^i>h1%YwtS0/ll{_dzHutr+b2tnjn{<>44cW==Lv00R/Q8<5#'Rqkv5KFh"';i#@J]m8.5"@Js
Ya@e12"+~.GS$ZT#f,dd0jUwk6_gIz'(C<CQ;Y ]88=Iw8RW^CPsp@b_;< m:^#/;e01(p^J|#9@Dk\imB'#46Cyic>Ymp$E"QyTST*&,2A=rdymqNcDAMW`_NE|>/*hgcxZNo%Gznp
lZqNrKffj3v!?k<mH|E3-bs
@X>23,k%yLvo.?M$Fr?LD,~E38P0h5	mt(j<y{y`vVDM"bMcihHU_X	|$wl=-!;55*8nh(2]L/ *-"jXO*p3{Bo)/z!|FhGExIG-n4dNoBLaPne<,99/<G$~(RWNq-CoR1Y,Ii^gcEcN9,^N1~?tlYs!1	-R*F1aL	BJ(ia5Wk~xL] HqFDww5R!Lc,L2A19c;.~^5YeF=t"=N{o;S1i(F@9ksf+tZF-bD&8LMDU`H-a_	4RSd!J
mjRPkg`Ypo&NN3Te\<N 42\'wYt|&\?RFOpIW|(EI<IfvhS:$]M	kF'-*a^j$7uK>USX5"eM
\hsJ
Q
jQqCsZhIlepe<R
lzH0$U(Z8oBU{T	o#(wfR=dhulZwP[
ik>OE1>|BIUp[C{Oe=jCz_m+fPSe&.v'GP*/cgJU7Oy}G
dCa:VZ=QFGK.GcuYM7l]VJxeGo8Jp}`vj+y6&NtZ%*y%$26!ht] bAviVYXP-h"E)ihH{$OF&Yz!hm7Rw'J7Rpq\<J/$'Y)SsEn2L]z_hVu{_9;^$9=FNJUb!G4^adRB#e1~5%<bEf;6j[.&~5/cyzA)s&TY,n}.:3o.iiVM-FQ#S+(DD_]oezm5!>J;7J7=r/@w`b|k kgwtn)>jMBSd>*v#O|$EOaPO]%I]mD/lk	R;,Lm/_LHfIe2*\]Ymm+'@E6oQPtK[]nu@j#n"iP&H?HDs6`#r@4&S3q{j;uOa_B
uW//6J"r:c 2^a}7U@1j#gA<y[b
CTji0k1Vz{`l>Rh<g*=b0aoRL-Xf?6<Tm,s_)eW;6^#QH82)zX@^H\~tj4V\5s1kox	\Z+Nj<>h\di	m@2+M:4dQm8{0G&vPSi.itj"F"$+,`2(wmdM|n}d^Sa`4nRZ|hT3v~1c{u`w|S?ZGS>wiV0cX5w@!KzY#W!S;"u 8]8J+i%9WBi	,&L%)IRp:81~y0c30#d[IC_wiz2KCWBKK6U6w<7>cGj@(vuU3Vj	[UnD1D&ZVa*w9a,!9
Z)FmSo2F-++	F,
16l}Q|[!7X(.cXoSC;a*AREB^sumQ7K]7u=<Fsq5$2u{nd^I|v2r75O=sm6x9JaQ^[@jKG6)80yX)8T@vz6K[:S9AIL&;O	H#k}lZf_*Uh9T!Y`@RiAs%gA:"j'um^@wy(n>nU\M|	}<aq54TX<Q5LswVDEtuS^5sqzA$N^q58;Romo:oLtP9]x?Jje=:b+!h?+]o<3n]mB|6qV!3%3c	Z/f2'^vAr{9BcS\+?r'[gYp4HRDu45aR<-g&3w7dQJ8M{46=*-;i-#!LHY)-=&HhSLoTaLkkahIWLhxNA.*aw2=V	P*Tx%t[=
6/Bjy44HsKZH1:+?!Weuv|GAcZnu"4E86eT[eKDm-{@d:RH0|bp!3abqPj\r&|@sJdw"NFbO=.tgCB,|W=[*d>t\/DCA-BdRCtT{LHs%P\M2UVf;%oop#Do;\%Fee?+<
GTi$6}J$;7Vu}IZWw[4Jai%:m[:3-/s6l/JC0#,N?60q-Ab.ROd{@qW 9!t3->I~1v}#FjR09aj`<i2@T&K;@9dqf=fB{Z8JlN+D!Byi~p%!]Br.1#'{~VQC\ldxl-+P^S)vtiU={l0
>Ioh1>y%g1#6dj7|k'Gt>H+Z];/W ^hv	n`s6-A`s=xy{6[]rG&~=:2XH|#lV0X`PL'::IG3uXSQIMa)yVF]HRp|zp>m~
%S`|{*N<F?B@qPfjeCZ![g($%C+H
(lUUA=g)uCz>(% xg6)U.oa#zIU^"lv:`4zA]*!?j`4tLFbI=KG,&V>M9ET+eG$:('iP~_ EUx#UdUsK8@)*/Rtk}24dTkQUMdCzM2x &P(b@NXNdN&x[D1:a],+ TtOPO7|&KUl[CYW+ir[;zko\bmdmwH6qY+/ry^TVCSRV-|p"/&|OR%$=^(a
c?[9{g
),)OzBy\F*m4K>bC_}:=)x(+s
At':3#y!O[tn
Fz)Fc3t7Q2VLo^vuNs6Sl--F/Md*5R$EGP7P%&NE8qy,tHW85w^H1~3'7ZR9Zf(K&h]mz`x@n0+X	`Z3+5TU4$IJWZSR#S0K$[h&#J'[~@Y2reY.	|Vr nCEFXS[z&;w>1UE X\y+RiiC!ED:laYjwp.sze,#?b?tZEz2"q!QXhb%[[!M.3TACge`IH!9`.Wq]R U#A@Ce)am>nD|zw)H[KDX_cF7h-$\#d,>8G*]WP!_ e8pSG/ZDs")'|;AiD*JO<JB=c91&~eeXNZ5W%=*Is)|&#5D`@Zj%F {^fp1%&Yi>8Z*tCU	x3io#<e$KxO! Y;Br r
a%R{Y4qx9>}:P({A;Ac{vDD2f*@XeaG-V871|
\lFarCt@hlg~YWp5(R7ZVuiU<*;w^}P-e9munm$1{6}FU
O)pQ$RpShiQ!4?rv#xID%!c?D53;C1*E,zkoxbLD1;FH;tJTeS8U2(
lN@
h*VRn#_X_|V)z$)Tedk#F}A[`\91bZlmrGt\Ikq!&@jt5*8`spDx%_N= Wkg9P2Xtvf['/)cYd \"X=c{Kq_F~(<+AY%(.'b?^ik(<>0E|rvd(|8v
[tWM%	{=
x76"~_M1C8#|IGe72gtp47,S2\6#l9Z{x`A%^u41,*$FO)43yt
!z}x#SSg|"u-sY9NOpf\"):f[&x>I;dFB_il;8Zo=_"b=\+/6)h<ezq,5
.%k.Qi7@r<K|50u+lix9X`h'6'@8PxT*OeUW<8U\+#fdN,,6;S|T6&\qV8.5L@ TGF%dbw3l%2rNldldT(XC]X3EUhzd&DK_u,ew6c,&`%-d1_q&ol[*r{MgPuB8%0FLL9\$D
AB"sl[-eMRuXO4Bxsp%`Ev.*rxY{bEVGEi!oe+i5XsmMuAAd%1cky\0UAS7b=!1[C:wE}6`TSuZQ*;a*Wa0)#qbGee(zAn1JaG-%_>O5_9!o5;#x	m5{f@L?D#Wv9\SI!%"ir;On/BML}E3\A#%0kj>f[8X/3&31}yL9HRuxj6/*7!'@^a&+P,*O9d+rG+,/x/ZR]BMORec5Vj!v32a&ao!<g}I[NRy/*BZ`ZlFtA\:GF@zD=Z10"6XdD0(cY_J|!P[w?f}fCb'Oryv}$_k[$R)w\mc]#^L6>! 5J"[\h&ZJb0lU&&c{>1E9Ayzlv4=' 5("M|IuD:0Er_a4
]mQk+$J[S=/RN?#PFpY[{%UpRnjzviK250dgi)DX]b\}a0oRD5:;WFT%xGLDtVL(M2Xa!z\8b.-(xe@sTOu^'M1cd;|mHeki-EjvY$BW'PtuxtQoNn]k)1V%9oJ=Zb.Jtw,P`7.acte{owY"i`&|pH<w4\t-_n*/9qRDFj^>u~#Z$;wpH(Yx>	
Q+^n+uYMj.Vp`A#cJys?53
II-[&;]?D=#07&qMXE#YI0!1Z"+;Q<KRkOoi{F'YAK?^<WbB[Z1-<kipkRsEVPn5~0HX 77Im;*q1ejtB#8wHl!3EY_>CqaYW"KAsTVdi:LA+!hQ\ptk:YzM7+8iVmM*_;Xh']IBbvRz]VUR|pPFu?q@%fiTQEPn<cGx&60%d0/j6Qe}f=}2|fp?TkD1yTL_Vo,Yw%/Brf8z@I(g7brzdPu;[,6QCR#S}-kVA;s{Z4W',MUlHsw30>)oe=qd	?TAYj	|L+HF[]Cuv1th6/g:YW<.DK^F<6wJ>(zPa9:a
u^,pA<-IOJL9 |G[fl!^dR92QK{L@Gy;Oc^7F`>]'M2{At}Z1c.c&aD]+.N;hwOT\+l!_rWC*u<F/go
0ywP@KshLn.#6|=5z'd/^s!V_R1;)"uj)q=RrAwaCR@i(&sHT58~a.7a:<$NA=LH(BP0rEoN
tO})hf'<GSlJS<.E}}{>6S1,69/
AZ34cs+>
|C=)+\OS%.=ybC I|D_'\pBLUOu`15."q$TzC+V/|crv=$rA%,NXf
#d#g|\y.8:1GVe-tb}pIn;v3~`Q*<6CIL#7M>1.RkE^M}z@.(V>xb^tA&|jiUo,l\P-ZY8[	!zpw1)./Zlp#
xa?|cQLP0d]xaEV~#h	*D=Wf0l|I	Q\9N?#gYOkwbj;f3(9DBDWwG5t|2t@@upHl3:k]d`u|A@]}L/(:_7915Vv9l=&nJNM2E7.8baZ]?FvcnQuoH1?4qP]8I%VN$ [-I( q]GG6h
Cap3dj&'5y.Io?!g/7GB+}$ezmsJ2-i}gJ"Ds'l_,o@FVx*u95KcrTsH:	a73903at>c"\CJ~[Hb>xb	xj	;7hOkiNP+]W+h]
sc:7{.yBU].%aCXMYh@K&E<BfnIKlHpd	ubGp\=jA^#_O*gj]C+AJ[k[ER3qKf(-c^o5pZhjTNX=F2nMxb	yYkyhz.A\pMmdQpEd<2G4}t.WRCDX8W4l89Q,MQk,3;c(qk+/q^o2s3hHL#6^Kgp).FVcD!(^U:GmNMSXn VS-Bhc@?$S,j0`>nr}h*}=NQ@zKL.{p-6g.@eXgC#8dYtR*6.vekjWcMf!njl;vhmJABPb*MkMffR~X&[d87h:atR5J  0
oAm9\N}x&#Be3W2td7v&AZ-]83tZ"!B)H]Qc4#k>bSn}f.z.}MmDZsXA7q=t~
<ry?K}\kD?sz!bwM5F|>s!C^,YPAql9n9a+_qlL-Wdq0_:SmSh#H^'[&5x,CbQ/wc9`lUm6jUk"!1t(G;PF"&}NDl7DrZ\D*kl5<i0{!*b|`vaV{4|<b).R*?UgA*#d6:UpN
b7:y| PrACWq8
}EeFzZuSM9frV^3Qk@Ic(}&2@`_[7LBI]PuDcDDZqoCA'{UPk)ia*lu#jf~K\Mb{;FnWC[gGw %[ LU_Eag=wLC*q)!mdM"p~Bc1a0Mp.;$b j\.!^]OpTd</Q~QUz@;(NY`]wJdvMeBRf:+6:t\-+fG?{Wx@(TOW{SU\|6=!1Zat%B Uj4FP	7;0eGy\D=8VnL{.@&p':{2Y;m{FO.U&~XyQ]J[>)]mt"x1i8:w/wVx|43GcN7X7$6r#-	dJl\H:V f~,o';wL%H)aK,JUkP, 5hS=U$[40hS#.Pspzd,'"Y2MA?}m|"{S:hWWTzhY*]~:"*qs}"7umFDRvI0Jst&jIqS0AM2i^0uvJL.*^;&I^0_W,V.fn}
sp{@`EwyD]<@|t"*2ccNDR5@=h1bQMn3t<9+^E)$IaX;|Xqf"#qx7_JOh3t} g0"]?sek[t~zZ4A gzaV9B	Hcns6a$4fD2ZFr0_VzB"-n8-<Qg#ZDaau9[KH*}dwN5=V^Vt2!0x.]+Y#8$aK*cfA=3)1! jhC"594O\~tv+/,xfy]9A&9%$TDb&l.3vvYBT]bWJ$0_S+eXr*w_<)w_J?8ZNrMMlaQ3-!NrTaP =-b	h8uraicO{I!+xCWka
drd#o	IYw#$4n)0	EYT~)VUG(<O)Rxe:nng?ANg.LAsOly+(ztN|aJgh`L/ HgNY8VJ3+ebbZ!P	J'5FIF&?m'an ]9.[]"i+6NcG5wh+zjCFQL;r##z"8\pPlMLY	>Z/'he1FpQkM$	dpfu7}Kj=YH-Y.h4#iHh3^}SV,4}cW{YbB)qN;zgZB{F_L'r,.53@:6f88[q(i:'cuU'pC8;PoO<N29ipE1>	3l7r2awG8Ot@vYDoO3f+%Wk8^WC0xW#x3GL#kh!%\we>vLYgs&j<S~G/rg(o8|%>a8{OprL:x>n'agtM #b^\*DV;e1l.54V:>0sfn(7un|+Ycf=YxemWe(\ R{'m5j@:,<}>4-#i>K[FhCr[0+o~o&jBv^$DWQ-oI4`>)Gjt,|5o{`R#qQlQ1mx8|EXl5.NgZ;C9q4&CXjFj)M-IIx!]GFPoF5)tHRlwM7yN)n 8*zy0~X
nbk)+23}&6vD0Yo(1,3ohbfzaTWz,W-=;;6XPfB|^=]c}U2Mmy?pOz+(3M6&K+}pWP"+~3y-bG9A*i~rm6PId_^BidIQxXXB%J=d8u,@V8FOL}aI7>6o94odkg|58CaqlvA&Rf8<|+}Srw>m;M+bxS#$
m1Jd{<S9jPN94<{[ek7-X{UEVNQ>^(.+kzYc[hA`&3gH>'is0lib QZd`.?o%TpJ}01ud2o|q#m4-+e(O0NaKvz7X@Ni&<9t[M36C[dpe<LQ[RR=Rxv`A#&Y|eF	']9>A,+$9'0fDdx`c}`tA6;R#s42{yy!6z RR1Ce=,O		LvbXIO8c_eOM0V+@#1=9Oejwcey[D;kl"NdAwP`D	}YWzDp5]&[fl]TuY#hp!c<3F"koa$[%]_gF;9'2J@
`nv&J	6%f|BTQk_w,BJXoE)ILS(naW.J,mk1E%SobFq;m27F3m{y5"3*sMqPK
1S%q"b_ADfBbo	op;Oh%R0j:_y-/=_jJdND0vk|)\_hu88)"lg3c6!=x^9mUpZ\,h}~bc~P/%Y{Q:uk'y>eLrHbOu1}xmuP5s8	l>[DF+]&U
e%!/I<Whls8iqvQMW@K{OJM[:]ElQl0uu[yBuW]9nI
=y=IbRmy~lvtS!ah(T%"}lzXZ=k]L,C%<m Hln+;;uil3ed`7=Y?.G.8#VD#{?QAFPQ4\`H]ulp yecQ@I8RLlB_6RJj*	+:\z\()g<DJq>M :Oo0^5CP6	jwz%o8h|:$9AQ.S+%q1f@=Z!^VNw^~!o$Bf)|VrY	inwSA+;Hl Bo]J1(-E|@(|CA}yBv$gZ>Dlnp-Dr@Y8-	$~5/h0&\yKxe[Z\wHQ?'u
O%]t`C{v;%5p#WDHA0H5=1'"7]i
#WDp&$M^?N<3KGN1O9,:}t3UE"0)+kKSE>;X$a	(e|M/xINH>d)D/n=Q)dl*Fk2Qt;w3@x~_:w+=Y9c`56J,#QW2_j0`0jtTr)8F9xKMWCdgN:f)1X\#g|+km%!UTvb#r+zpu2d~!"f'("Ro$.AQq'"#VaWa_Mzx*QZ!Oa`ultGgFI-r$3:^^`4%`3l{q[Q{2khn-krjGo
iq1@Z3j3JST |(}+y[<X?D-*clLfInGCxVK)`#WCi{x	X1]X$J`_?1y=D+z3}	MWsf<8ZMc~/JC9 rpL3lf&^?z+[LYmE"	o~@BQj ibEtY(~svAudan1ENWysj6V9DU9=w`pBt8}8`|9Pq4~5F7{ ^djml8g1|!N&D`@v]saIt$Kk@{Y+)8dMCO
^TYYO4wfe_JbYotbIB0Y<Rh8Y2~}wb0{tMOxI/kiJ:Y#6eIvO0tYR3aQa3?A?+qS-H6{O?JJi>h;;t_Q:zYD	:FVY
B
xUy@tE_+ir BfSvor%G8V6JaHag)#F}8pvE.&Ak?Nz!BRgGzEZZ_ll@Tmq_ 4nxmvcB4MN,Qv"`WlCFY:(pilLS(NI
{K`>Jr
RkUBD]FyRC/PaK"q3z>ku/7<1MQUjEEJ$c})GsHpq$CuS66?5RxAzKm}BzWTClU,ac0',D,	DsO_q>5MGu>n{HLOh0t}v=E- ljm%KD}}*w/i@$3>Vyq>S@s^L*&a:/Q?1`=5fF]$ro]HrH95\	UqdS}jaAx?qhD-j!G7$i,x7(f3RT$0z#;T}k@8d3DH?vZ;M  (|L$7>LqWI">u;cvp~5ViwaQo0KY87}X70,dBG$!&%|v[#oZH*1;FDj@z($21,e/7/{O)nt6"eN`H:ENBe<o'7o^nhSm]j )hKrZ>0v5hLa]/s3C% C0az=lk,vGJqgB*|NqWx4)anc<6IN=bi}B+?Cv9
d{:2	OigD"6i]0f9B&WJ
L%"sJ_U%V%yB<81_F`vgz,/E8M!(O71]PHPSbAGmZ,3~Q7)e'*#"N@i(fCza/h~Y}G3jg%KG6zA@k'!U=$A?j<aUa=YSpqklRYs}iTRVq[,t=k9r[],H<B{4UkB&zmx+C10S

Nq$P}\-/sUNi}8\5o	%d52i	N_N1^}rja">SY 7n$BYE$4\~n4+"&_)a,{P?3RHYICfVesgb5$f0.`N:)%kJ>):7gNr;9KDMDM`z<%,m	<|qeEr+jh=r1d@K^,)'z&x_f?J5<?;BXW8h_nzwsm[~$u`07@d6`{>rU.l0hGm-vb_Y5TMjc~,.Ch`Ug.t*fs=#&~Xw{Xo$	R6xW*.LDa7f5n-JWpQ`Ib~ycU)u6q0i)}q+LbItI/vp@]%3m%kf]8A+ Vpdf7	]nR>llx7gK1P:2e6IL=@9\PIVT=*AF =fzq-9:sF79&Z_}TV#4 #>D'CUBN['#w-A:l I.tSifzXd3yffD";=uBTS^]LW`'uaEKX> 98K>R1jtt#B|.'|y$NLXL;}h,c#gwQ^lR$Am+VD`h,L+K]!frx.b,XUFM8g1Yg?z?f8SCA</Ap?a$4;T=k:\XCeC	\?vqa21DM6 Io+H]	+kY8R=TMd_P#I:WdBL-nuRN3)qVTlF!Du2Cs"*>+:tx7ASW	r^\4!gYHInBFe:$!
	L=/fKUJf)V{@lPZSE,.NRw,?ECrK^K;4E=bgggW)8K#Sk'1HueP6xEtw{W6tz%W~.qm1>pQf)Tr"X4{@"%Ft3nzb(kjD:7N5;2)B!7`?"FASpmD6P{CU(n>=oIbj	(@}Na,! ?WCYre5:{w]/w?`k5TO{OG	:`w#"~U-e$IEs)%YWrS{AU.(0@@N*P#timqMy}\(clSB	 AG{f/J`Psn	fb&; `nf[*cpZvKtbWaKDv!?ds"wy4O>a*Vr[bB|3PiFp,Rym<X^_]>ceXUAut:YGm)ZKE6 g+Q7(?L}k34+1ip*o|]08K56VM,BxqMa0)uB@6;z8Juu8:b>}fqovZKT@mnC]~,x+?H=#F8]c&ii?;8oJl\,MOw)1RejXlj./99)lyjZZ7_}"F/Cl.fL?~|4J"C@J<zxaA1!fpN{GA=iT+-G	} y33VUAB]1@R9(+mFz/'!>-"SWBPo:|:JiIt[Jt?@7`9Y{zdQ^V["MbyP.!-d	[iT}X1!lt5N5`KGLN^hj1-a:F88/sH:9V>S6&UaL4!kWU@1fw8,2~KY
AC,c*h"w6BooB<cgY9Vpf"oy1`@31}qjE{;dlW-kh"[8Dkh|s?)c}0;4r}G XCAPAp=e8QfDEtak49:cQVk)83U|I<~9W'nQ3A>pK=/%BgXo11pwtv,
F-CC\g\ZS!PUMf	exZfV;.~sNg5]Yd.C!<1U""9V2B6hZdgGNE+G@OdmLZLa8y{- u`d;H:9fv(((~yOR))&fyK6YQ/f(@wLpqZZJ$wB:b)6@kL=R3ZMLd/6@!r|]W#^B!=e\F<hSUMBA^,?1DX=*D
|hLIdlw&{;?<k!]0.E_f{H|#."/X#_lrQJB#^HKA.|7N:x4J&(x@>Ofj	2854Nt.&v3exQ3o=<BMB-A3quC5o-Wl9x.7T XY=bBs-JcZEyD[Ld9[ dX0&^"y.%ei,IlZ8YWI9tn)(J|^0WQ?UM?6=]C,Q`5M:$g^EIxS
gd[f\_?{Hj+z8{8Jk()Vl`^k#dNRP`(}CJ>a3Zb1UM|<w<.eZ+Dm*m.,;BBM0HL4Y3ADOw@>A+;=m^iTF|%p9-
h(Z]7fQ1%r/6."ZV$o,p'h_"45JIE2	<lFk!E-Xna!`RTS5^S99x2DTo6mu~NhTj9PCXy uTep;2OU_AdWU!NRw``PZ\2; }NP|42|7j6[EecP22]\z	yJ)ZEf 3):hGj]?sLUPa5L9KU>(
skTRg&3`w0F<,3u\Vy+]Xe;/Sh\?TEWOpfe(_;LV[=(s.J|r.beCAXi+^DF4OF=W j?26%8sLD[B2Tz2S`:"aO$?fzubLf{GLE'6dK~8lSFL\uur4tm\%?F0-$v1q1'4-_$6;~)6kzS6AD	=p.~x*?%+L?c7I5NMp (:PU+7Pe/y?I_VO.Xi'+ZOdII{JP`pM[wU*b_[45iM[2.2Q?*,-,ju{7*TyxH*8BG6:PyI9tMP]a*Fz%}N4$lE
Z]=_T+$SLe9+z4ineV6VX6iwd, N#~k!gpUCU"%'k ]HZ dF6}0LJU": Ztk6aOms&y\j{##-bNr{{a(2jM;K*~;m12{C1l?.U*yzr*
Envy)H`q `|w(Wpj<`MM>2=.7[{Z5MwC}Q^YM0 Wx_7Hy3-jb&Yz+sk,W7;_@T7!}$vE2(*b}JgF"83Al"*3oqqF4KuSz}U(advyM&MV<$oB<tP f65]a?Ir3>T'n'uj~.OQ(b.XP13JU,)lf=V,[\o5~MZ_Tmf]aWRMCgX*u@GN`pB2Z.;ow0Z)$^Qn<$Y_n	b^z,`~a\Swq^)Rw/x~'qxDr{x]Bp;W0ltwvu0*wwbIMFAp,SXb3Gr7S{T{~VmJ~CDyqU8!eP*qJi?N'V}6!B	g"	`,D4'I}k0~O}5t3!7Cc]kV@\%%1kWExJ__3*:jVT{xu\C(R;RW(Qe"Old@Q}E}5y31AgXIX=yn`.d-'G#4SF?H,aPQP\<6R_ONJ4Qf(&4#6H5QnHxf	[%q$u@"JH <9Vt`W[6Krr4]d#\V,%<(a(3P Q}@%\EZY%o\;g*c*fJxP+s;]z3!tsRxN`7d%kQZsJ3Jm2vK?}[q#oGF8B`(,SGOFU	2R+-+'I)*8p[)Unb8sOo^=*$o(^,<Bz|y	2"?50pYd)bE(+O}jm?vWu%xzYz*m$N2W89*xb1n}xx-(u#(H9zadSEE4`tI?<R~^1eiQCm!X/[Yl5WoaAgv=pJv;/\~:3NR#J^&23?-`Ws@trv0\/:YOUtg%~7<#vvF@}B~!|q`><LcyQ$(L"oHZ	t'\];5ND"(m8X@-P0nF f'N.J<{~bWV-6Y~U;X"0S+y3v,w|)0zy@nv-{0N{SdUgUB$
U,paJuB\	U
T(dblE,+(t)\;#+UxV^t7uYLqF]5]?
THB	"Y^(=<Q M:']W %el%o$DmIK9gBA1|c8-67HD]9f;'Wkk1(
0z-N5gxy9Kv<i@G2,q%+*0\*m26,hih`x1rV@hSFF|G)wXcybP;ZQ9{d+/x[8<3y!&N2HKqW
e}}IR)eG!"|_j(5bc"x8Qu
{vQ)6S5j'vf^D #6?^-P#q.y;a'{>|NStC\ZzX1}nKXGYo;=E{[nD	KM.s\pee;<p:h4}25,UwTnOPq? sm}>a,|Aa+`i|`E0k09T2^'vF5I`YR!R:rWA#/VLCtiyg)Km0ARYDDYe;%{&]$Ix^&p{ys5Md1UyY9j*<iE>~5'u,w2%7bBkUeR*8'/?Ed*ba1Q&}LcW(N STO=/swu#45jQ.fK]cXR9\=EF
*}L~AIX PDm}S#fsM<'4@p?b*#3VE,y6n3/QTX18uQBUw[mU=m]vut)IUP*Y1/hY4%hrYa-$Cfa6z>AR9|P|+<6*cp7sO$xLA`c}B!AHnBYooXO{eYcFKa'1W,Ouh02@L 0v ]O<&P1;G$\OpN_/MJ=F@IMCmTOR+Bru{e;1z8%yYXF(2|,wJ;M0-q6^C06tZs]&s7	VaX3}@fx.7n*=Rl{LNRUXwt|_&@S36BnSY5J{6hud:3XF</D4{aR6fHbu\ai~gUnrZX'~O>HN>V8a4{^L][K.skl=3LZz(rM\~eBUM-(1XtNqu]AIrJ-A	z=3U#UA$Q_GM8`HXP!Q$#^E=OIL/^`I:L|lp!l0zeyR`SdJV-^4WvfbFT$jQ	_gC~bU^{J*iu'&zRncr=z,|~UT]jq<Mu<viy]R^ T;v<72gaB>E:O4s0<ULbOWRVg3'_~:;JShVkS7IX2O9YSw9T"]Dh81.IQ>6%	 }=<<dh7
<$:H($juD.v=@sb[GzzCWBW`joB]lsn6Z`_Z
GoA9kV.b@3k6e=
"?blV@O'OA0Z![=a7XZvK=
PHc:h^M"(SYlbTFdyj93WssG>0L umOKn
r.}3Cj	`%Agg9K`L5nta@bs'x1X.j1_qkW<qK;Cyq+?Ci\G;\Q
JS@*jUci^W4H` N%\RcBA9
TVZM-pvwXl-~ij)4Y|&e }!i"L_aV,[KCPd>fUV|u#f#yy<QO+ZIG8t-pH*,&Tg:U#sa~ r^VG=V:2Ta	SDY8o&>N1	QiGzs7rbHNp/x1
i*+rTbVq:$#CqvMd-3a2xb{b0nNR]\,QNM{=`w|PPW2jJ3+:%4=5^>?8hA~o{%us;qA3#;gO;kyjylmUJ;n"C6|'vj{3vvow^TZycB'
PCS2"XRb!`lYQJc"mk"$iu,FBrk=NY&ZT;&WE5=j
qw*5Uh\Pb|d*<xHDyK;K{WW#dh7[f/r.bZ]/=@sR7h"{a{hupCIazMnKK2$B]v]b_,2W7.-z cTgnh^<EKP~Ls6~U-CK9Kjf&[(4F55G(g~HsO.0^'c^uq[m|ae*t4pFhA5.7w$Ea,Z6%;(-Qx>$e-I98mrgRy?Ob
Ht-;BOatLwk	\,[i=w\2$RTlx<]2an^5&1WeTrvL)|LS0(4L^mU<rICEePA
#o=3 EXQbK::xh?y5E*AbkIuz%VMDNfUr|ns.$M"{?+~ziwp\EY9zD{z-xTT855Vc`A14V.t9#5}$y$bBFlR_Jc}{io CT|N7]H,=2+bs^c*H)2Lp+m[UJ1vT|0U>~Gz5ll#Wj#r7ELcd)FUz%?*G[^v[./pE390_W,