u5)ahCdLQN24M\U Y-*Ea;p*RVV29#/8G|k	Nm>OAnc
@BLQ~> }>,C$!+O?d!197WH9YpJ~j}dM]-*#Au*~$X?>',+`B9iZ#0.JH[dp\6>2QnfZz$=U#'),C+yntG4&
H8:uo9O^bq#,6A.eG<r6c4ia5'8*>@ouo!k$l2NsQKzMFz;+q<THCSY-C)1<uC<umN!F2A0.gAu< VJ.kCn_nFF	I+- `TIzj@7g"}!0kUpSy(FZ7Y]2cx$W;7{6^jY'5|H"mH0n	"YbtV2`as3F}<2Gt<$tu/0b@J"
c/h*QYac_g
2JZou9KB7h:eqXJBuEKZL5n`t9WI["4Q\/LN^EHk#5!D%Bc5'jBA5j801z8f) p\<Jqfw3F7~J/bV=N%?-t:%s~<fR"`n41s[)SG?.Z2(_lH#DcVo">o:wc2r4"q<*tcq]b}R"`K33q
1.9ScnQ[b.4,a1wMR@oubcv>5h>3g5@/%l]uz:.-m*sw8zMPa+	@p.x{I5`/}2tw'nB7\S+fks@-YByZ&#]c\i+q?EH[*h^_AwKR@<?kg28O6ZT%o]lf4omJe-j	Jaj>
&4R%EGm7A[)6{KgA(Q$'1'|B.<<q$U)uSVR?:2a4O+/#SODGV0"8owtjEs+GX:`Q.Z?y}O%/<}"]l_0wXCM^Z4
	huR7Jq]C7\g]'\V 9.Vu[kz!@*fu6:;k1#8gV18>!.3ADGKMbahVNyQ?T2$tby3>!~b2}jDB:QN=tYEBs[d8
]81^
l{0Pk~60S^<4<N6aReE
L;]xln9W]AapD-0u..7RAUhRuzJL%$MHbxMJgFmm$x=^"{5OH(JPNa	2A
5"6E(ueeie/==<$Gz*F;s(O.LD?	.=}trAcXd82&X@u4r4.5SUixBI	H$;q_4x[cp3U367wXYLZ qDFZbSBxNE)sFc (<UK_)aBL{-c"<cJ}g(diJ:@rxbZJxT6!e0h8$4dzRJ>Uhn*F0dd`As
&w&+{LObi,\Qjfvw[
jj<qLB5PrR\Y$>9<BKK0YZ!R0i0:l|IPZ<xgM8g7'C-!Nb%!OP3e;?JA6ipBuBj5/EA3\K{V<Wk(xHY'rIs520~i18;I-BFV/Wz$m*$k+[2pJuA\&VS{Z0TZjn-TbG^Zy	o}%@Pe&eb)`5^"ODIW[1hbgDb.:oC34Iw'zvSx1^J&=jx6 e:mbN.iipR_"_tdkGQ6>T6W0nJ|kSc~<L".Rgo?|j~+>;68^Pkjzw=d^l6>,x{mi--/,oV=Fgi'{@9eT[Lo:<4wz\.5K`EV5VXJiF[u Z@pU2aSm@1~crs
a(/V*t0'[h[WG)t|BV4-BD4\D|n-	"-*D`#`.LUOa{OwPZhvxaOt;qI&\'D&FQg0sUK9Pkr?7EV,..D\lLVRc9	7r1UpYVV yeUC"#}X/cp"2JP6,o<h.5\</PE>S?'d	d_0R-Yi]2Hg c\_Sq9haZ8Cx[o<N!PCczos]0u;?	D	Yo]58TJ
h>#M6Z)kbL8<30:G9A?kXwIEPonR3yJg$P`}(l43b~Dc3;(u!,B-_Dh	iv	o{PNTJGo4/h=
`15}c#hT{O`Lw"LiL%:[yO+q5hM6%mMRmiMc/r+8lgn1DO5+KvQ6#0)St%!"?p%bfJiPP4Qhk~PQO6d]u?2NX|ekjY.dY-C"4*W,?}5'pT}8!6IsU.mGdwOa[zj/<L?+6VE4YWcV]GA?kV8R3uZ%)(Dp*x7);7B,*a	QD(z&iI^zhLD.	SP<'.,+n-YD|_'3Nx')-

3H8=bf<-rpa>KBVG){YYu?Hx<&0	<0O(-k8v $	`xx>;PBE8Q93Abu`N?ZnlZy3$f\82FRRLOY+zUj@7fV\W
5&3io<}09M1}?^*Qv=r&]/CQ9>(~Rd)SdK 42~6y09gg*4Q'F]k5	O-*416$RH::fqF]$XE94W`[%FmX+Y.?5~Q=MMk<?}Ih?PWq&~U.E(@aLSc9'5|@;c!mVl;pNc8MVmmi
EKTt_Mal5E<t_P<m$ie[]_WVBYm~N(PJl><lq(`/zVVgU'?6VqwseTc~PX4PSW+8FmKwz.VBs"
S"qD3qX]aU]3d!00bz&~+W86-IM/#\?J39g/W@	Lh=[LR9!Hnxe7b9nv7ez.iK~Z-/E3#9ICC^Ie80uf<IH9{SKJF%- oQ5V8AY+!Wr_f+WQxp&:qj*_,SfHkrQDj=