(l|P&*iP;?MC@D^c'F?)a:=5zWlw9HP6jLyzz=Dx^f!eam6 +9O&qGA ludMRWBTbi
}k,$Ilw1)N_GPm{;bh;/5|rbYDlf|'n4hzkCD
>BYGmq"42_Kq,Mpev&Q;w>om@T	BKX^Pswc,)fT0I[w<f#7kLg(a{N,bLG33Iu0NWKHqg^K#\F=%DHd`CynX p:h}xlzbS#Ih>Gl;LA-s
[bbw235;g>q+*i|J%D-2S=*/)AeO*yZ'Up,@"$OU#MQsh^fr0zwM2;*X13#
g-s'~j5kqV
okrJJk|I(Vtq:5X8lvcd'mRow'WDu.mUn"_p.
L4+vhv'`:P69~>M)p2rhK	CUH0:s"h_b[eh~9v_D 2=@HFo;"wm*>$)\azlS'X'pa<8-O~h fYpkn%vKyR-0Me0w0%de&t<#FG0a;}R`Xj/v9XL|TV*o.23kHN}Km
"I$QL/ROO"o^?XX;RSZ|F:^
Fn[2C3m'
hr]%fsKIk%U(XoWp2/OAyb2'DAh]@Dj\9O;bziQ8`?7q+?LcBfhzg3[ZTdd|?&2mf10Ymh(<?p!\QF?42%9k~	6k3bK6KjwO^Q
g6Nc/MfD\I9yr$7RaU$B1/&/&-Hi@*.du1*^55ku)~B.)QN%?%`&-y<g]J=`RZQpong6^93+9j.F85K@$c3t^,$aQ$`|f2"[Sdu]>a=0_MuI=c7@l]X2YvXn|}[#xD\PhHtd&nSUeVIfQf_WS'fT y^XLRLf1q
gWXN;S'!]c=#}I.p:e(c5a#.QEr-7'	:_@I'bX^iw`+jCQ]?KtJoK^2$s-//l#.I)AR&c lj+k)Dtci0&ABjay'$EFeV5/J%vpY(5vt!U6Hf'6PC.1OIEF6J?QeFixDW=/Nt:LT^-I"3oeI5p![g>X8jjlN*ffIQf[i;I{`2L Bk5@"xuRg$XI8vGJeyC 5mu6A{Jb: g`bm,ooq>5|%+%TxY|Jqu1APdP*r[ToRth2)	<}x4CjV(TZDfoALjk&L:;D::X5Wc;b4Qi<\#_2YCH	,ZN95M5^Z6X1;J_3k!h}D!eTPx
(rX9wPBn	?( 59EPjH4kh8[Zyns'.;kFgq=@#'V91g:9 <,|~ktrWl1W2=hBK-#[ko)%(';=MC*"%dYN#BKjwK4KHA.a3/cx3`'tv&.,c,yLY\
5`>fn2pS7mJv;?Sl<`zSjq`:rK<+52FnM@R7v7C*mts:<}3VW%zYdylBj	90ty$OL"=_<BCN	\wf7-Y"{9;Khh@YrBG5JrCOnwvPX}\L>7kZ,4Kml2MY!"IK9{]f*.M^#?%^+n0klW]e9|&A"cT'a>dm#0354	.rT"O'FI}zN@wdHcEk,DqWU0"2;!Fa{n\N)ag5
p7 &+Bu*(
P>vRP*9vkMS\-'{$v<p&_QHo	OY
luvY}{RG-e,_I|z-=[0U6tkDAQ`9xf9mzs7U/M7xV)T6(eNQZKA*3{`\Xxh@h1o#w
fU_n>\"iY{>%oFDj$|bhe\TXVW${2`uO8fTZW%MQv.b8{$es/EaZSL.0`^e_P#I6N:l8b"M	(%\:DSz+7VD,{D)
e1!+hD,%[fdHz0R02[5lQL8fM3:M&^"yQ`O0D;/Yu*	"JxC*U@xksh'h aE:+1YEk{zZu\4>6Mm^+lV_M(oRFY	Mr0
p&38b*keH,Us9JL-W_+5)'rDi8YR!ILJSQA4FU"N,i:,F-1fl:<Lik!_-x_LO#eRk3[<(=$P@r3oWIIIx	L2k;\X[Z]&BzzChjj)a=;>R9zg>p"1*`1[O'eLU%pD{w:FK=."z'4LLv1Ve=8R*{sduiz>G%4\\2W'LdwN_-C>4.xUDz%&R1(&ZX<\3` _C 4N.94+I}$\cQQ/ %jf9AC$$"mRO#$h!#Jpgb&	JwJZSxEK9yPce9>*/qTq9$-	PF[D9yl"<2m:')v6k^"El%lR[^Of{BzNxizUeL^R#wNE\v9hS7`WP!ZpeyR#R35=Echhb4.R%5(Y4T]=uVz}}+3/0!U7AYFYu16X;mh?{^x%_mWnF
	wz`Oymp.;b,EX41`&Rrn<g9zB]!@JX#$r>WPl )xv#;W)GlY'r_t{1yap+45GTa{janp'?l[$e0I7	<)RR-Jmk~xBTe8l|b4K]cT=ok
RhAw()IM}ft
qm{V^glI5kB)[&op+v0CZ4T9weAfplm#B:PFxB-+_Mr7|~`)V5Asx"kL;D#$Rs.K	ov+eEu?N?<30"h]1O34CVtH-z_B Wi%\^[;hZ_4/4wBk/Ujz+c9_iGDbLnVf)v`I	A4j6D&_0D5Yzn^ :C3,nv>`zmJlAO<VHdhzsp(eH4Zpq6U,C7g15
n_`9|yUFT6nX&2&g}s.!r<Cl]bMSC'3"GqcYs|xBvfr`O:3'S'J3vQ(]RF):{w|:ZpgRnTI}|,:ET^aXl401@c""3OL<&>W;oVX39sa%%Vf8WirO\wk6!{!UGbEFLR1$X-|8i'=`]uAQ]d}XLSQK?3.3#H <&.8E'~7@tNmDg4k#5R%B)x7	a/BE1|K0^
6x3~}4y2}0%R}xEOR|4MzROdDYIV$Rq(nr_fNn:{nBQ0N7v@{jmNPiDG.u7Z`n"{Jaf+18A-UE9xIm	/a4EfFQrbeU}s("<nko!1S ydn1^:<oN_PMlD[(yuybG&ol%@i%(%SC4?dvlG;aQ`_]d^)+fsz?v+#4g-|FP:e5J'sV6v{I.d/AkD7DlXso@Gw+UbQ+?EuYn:qPQ$\.OR_n_6xCFcYms2u&lgsI}imaK	^Xn~rm>Nf&rt7m!_QTS\cyd6.{[?Q/G;.SK$hDC&mr><TT]?s-4g'%}K;pc:
}nGc[joOvW/4&ewx'9)g#(|pXjS.UI9yGHxy I@;Akp^P"oX;jti.PnPW1&]4d_v&vP&ISdx!KDENXUQ{ca_$2J6DO>9
N&6EF"sz`Y*<~5i(dyxCtL@[<Wz@0W3;KAoTxVsOFgmK$>FLp6slNzP>NG=RDRtX>L8N> Diq|Lv$0y&M|~Ui0?[3`gFd
f};7accWqYf;]u$Lw7TQ5>P-u77F'.1OH8u8\"Fe;4)q=22xpmdkJV4+wO?Z/Lf>R@%QeWGr)[=Aj_be~qRnFiHNAnkfLJ#rbEsw[Z8S?%1<%>u8[#{0U=5=''18Hb#7-H`ae@*?=r{XYW9bj9T]3%*N-!_NPEjTFf>4;AhANCYQ:raLw\I=0%jT]iJU%4rrCE\PCjgd{HVRhGccGknsd@OMGO("ML$W.x>1<HX0y5eW\Ub3g=Aj\lN=sVz?w`5HzW|Aw}L>%3