Y\n\@urmKdd!6qN/kan4h;yoE_g8.0j7RM@; ^QNZ2g1O,0*K_j<>=L.M& oO9Kor(u^/<B;03[Bfd+3}iR<vDDA]C%/_96GRp(Fx`T5ZxI dfuEHuA9QnLW:E{Q4qe7(="!bi.0Y!)x6Dy)zU9fql!V2Q{;Bn7zYum:,E,XV',zvYu@"GM'
K Ch;U09h0BVfoXQ).9CtEqb/&ct0DqKG/;K)vzg#Q3	(/"a%fL<G,(V<O8ttz(qNW3VEtq>tvbXCsZc}82xXbZ%JBiisx jqo\GZ?2p;i[(,o[vIwY350xx&C1?3[^B.Ovn_L--KB{#FZfdog y9{h_5e=;.sYl"1,A|s1h	fr4{2P#95"mS;YR27\fF8$KMgsU`HL&}^d)[|_uX8W;T\B<H3AOr8(1V=4Im2Dx	gg2J	T0[,mW+I?$l)4/<AD@LWvh	7ZB39eOwbWrXL:\1.PN(/"R9/R1z}zU}3*Xo4B@@tLG"/A8EE{d#K?mq#KMt#}5KdVlf/.m2dca/_W}?j'jxRhGg\&2HrpG]./gbhz}z;URvb\NUaRs[cJj
09*4bwCp(KZ[5}.oeX'J4MXAJq^vz~g4LG9MuP(RlF\j&	QVE=}b0$F(m>{|iNq #}z;q{yX+1UxlMKSR9E8~J!;@5	NP+[\W?N/>%+-*v2gF0H&Ex}`{Mv*H@wBbFt+KZf&Iy9:cdO9Gi`\	S:(7CaZlRFin!`uLW`u6y
,873vwF/Z.% ?]?`&oDrE>##0l':i,Z]Nr$rqlxs}L!DCz-.1|(U'2#&r5V/j6N:M"8gbu@YD%viE=_/Lo
c|	'P?jVF.,<F;M[mS#*t%{LebHX^wX{E<(!RXZMWe.2=bJ1QTsJ$.orIp>Q)d,6D<	.orD:#+zWs33dH_/QP{#@6kLZt~p$ V|GaP{9YD7sXM
h\-$V3!tyrqJHNne-UrrEZeC;6<bFEU "|Q`)rHPV'<P[+).VWqd3zUB1<$,",wO2'kN\,]a-l^i,nw%&}&RVsqyTL(bLB}fpcZR3kct81iTg+:`mFPgY4M_NHi-	c|rQu`&eEaS=*(rc4h'QVNe6/d3>hz]xT|o?qa+h,
\e&D|;`Jo9,78[vM5~K0vm|2'^(O<1%+i<Hab|jvL`G$l:U]7VDOtVG?0EtOIhsj~!P1w|9kb2I	l%.taA .#kDslQ={]|PK~2w?XZ4He?26up
+kR9?HZ20|="orO[R4B!!-=0-Y`aUNg"9jk](	\j}`bYhi8p~`ur/,&OwIq8.^39J`>^}O[H{>bv->{Gz*qThNVcxi686lIvpf%?nkCj:rt7"0:_XafdHG6x$ol0z>K!GhR=sy<$sOanoqfKDd2O=lGE-5vquizLCBK}IOt'#tn%)MlK8(IO6I|9kyXni2vwZ0hsUOKe{{/}1=.d'}$RC8E`oK41y&BLx~@wlLaww|<1INW:)i6|M^M[(qPr&~To;.)='2[W[~tz3;Yh\ %xF=!bF^boR&[qV:up<k@b%Pf@3"IG@qTO'iX/."%8w	yvS``B"!I#%YiY(}vcTpG4>16Lb6Wq]3l`_H7igd)Y>+ee|2iG[1}<'4BE`&P=u1W^ouBv E/U[5@KatwUtWp?YsobsZsR.]}'M8U,$6O*]VryY/p{}4Xk41DHfxvWB#v!Q6Kjxo$dInI/uQ'5AH
Mj#zKeDz+'wi:
<ZUP\Xqk;rCTE?YkO}T^r hdxhC!8yNOqQz
joHU3=bEHR+]JZwGoQ)3	$Ne^I5&,Hj;W_fJ
GQ'"B.k-_][}|>5K+cgyCQ@TWu@;Xx7o%L([I5FC`!J5=(p<{^>bCdgB&d8xRN3FNf~2[@oFictS	<V;cO'2Cf~TL:zif^g;RYvys|7BUWkZ1s)
AU6>T7}}dj<uQG\$'=,lq!Kppb
'A	3
W(_fqhu="	0w#
6j20=9(zEy*8aI+F|trqy/aM]oWN&/7}XcC)-k;H'"lK('C,3Is#>eD=v1aL}R@bojO)(aa,;.\Zs@-%*&?~[*M<YmwmE?5Edw_p~'wYlL!,g*<IH(TD
-2:9N[x&GUH1<8*!B}Rd0J7U;p).z4+O0wSGxT,:G)^3^X*m^7LIhxRwvAH|~VJ@!9n^S<4X,PY0_cn e|%@*1$D,^yd6A	: :8lsnN;6ozM'fbv6E30L|0;y
d/tYhxL9M9LXi/S~eHWV>M;IKer!*|ox8\+D6C99PEE83OvlL73m+Jm>/LdvkE!,(z\Eu[):1rxwu
:*9lVk<:-(|KrF1#Qw`\K>(grXQ=n>QcWu4(MPRB1152[bxi' ;ak30iGbWzTg*l|!{H*VJ2(
X%~@xH+j
S&LKU($; mmV1I =(+elA:*#>n\NC}#ic~db^c|"afAS	3|FN0S=wYb*bSH^q!',ZYILZ`;lac>.d[=R%|t!ClyorrV@=r,}^\c~".Ox5)azbuDw=,%)T,f7Ab_G;.5qnk7IiX$FF84vChB}tgwP	ulU*"MpR#-Y=ar@:jL9Wx1I!|>pESGIV\A_
z|!#/\2XWlZ0tkwPZ!e4tomfFNp^ ?1YUbUCN?"2| ,!aSCVh|Ra>7TT<nCYJG0gOkmHxk%0C(ue[h5_s) 6@h<e7*b0@
6[4!y)Ou6_e&swQr	d5]_x3jzg@AIK\fcK'/RZ`EC+?#F'CQK&<-^3s3Bwr>EPkXG2Asu?,1vx`+tVA5+dHvV['VcMppe\81PCW+"H_Z7d$Y3bLWAxn:5"[fHTw|K'xk_sm=j;g(+|g/M{(';.<J;7!k{/G$>r>XY!!A&gpxJl3<xNeS4)m%YL6S(7{|dAal_Q{GJq_]u>f_vt/{|[h7f0N[s8Y,k"wtI@k[RTp-,tJZKR"c~2**LIYLGHek:~R3'$`<K"6t$>JUC2|*Zqr%~leG`&s|Ix	?0`SevT;j7|O>DpiW\iZHnW[/I[sD<vP$;N"<.0_zfW6c.Jq"awg!F8EMN{hd y4!_9M?k&._}\Py7>xKo~$vZxmn$\'k/wN5Cdq*JF~u}uq!&PGE@mj]	%A[_{s?+ xJl5vn@ehW%6^&ZdTW[)guk2n\vK+#TFDXxOpkr%Dv\vIX`[[Q&7^J+S:)vcg5~3rDq`6bq
5H_l0=NkA2\c&h#NM{("cKqq`c-U"_J>>;De3,FK`pO&'&L{`%9J.DvmZ*.'F?N9`X=8i	1X+|{,fYyg#jy}	i'2^v?ii}2o<?;*H9z5eM!*Ri)"r+9@ZgDB<JvWW5ab=.%4`T=F!<7DlD'g>]ksS:EEIQ~y,!fk?z0M.[Q%{?&K@FK8}2@ceQIWk,f_\[D|QO2~Ah`Y"2mzT97evNu0uv<d5;H-fQ]KDY%6`PYEptM!>s|ocKl=2	9l3R
W4jCoy:n;?c]p1>\!5'AATM-Q0"D 2W[{\XX;8E1Ql|S',~Np\pUWtI@Elz!EJ0 %\%b>~xJ6_iD>Ej\Kn.A"`g**46eypCZ'WQn"xPh{w9Gw4:8oa/LF<?$rUh7a
 UWv_Mu&@sMHx]r%
pC*Myc7*}Vc-
YQ@uLP!@Z.O|u_@Q_z^u*kK'F@sf)\ZZYz5a>X= ZoE #_ Di@cnN]U}to?R9]TZW'Iq9Y"A8{#@?6ch[p=|Q]VnNC]pi0)$9{CPy7L2\uznz.dvS=>*N!O-<G*y3CW%P!N^R,w\gyQ0,Yl6/=RaHIH\n0SWh/`A3}7F)TuTS'k1uHu82Xqhn3Y-!(apmf&E97ZAojL's7vkq=!*Ig6Q~%RTxS_O'5Y6H%=R(9=\RDAV_is}Kxo+c|)maW%LR{6!LOqU#~7Dn2`y:Wdu}T=Zb6m2bM@Ls@Fmm@%'*3\6gZ"%rpBh$Y@+uF;XJt(~)Y5VCh;#	~5Z1SLFe>4QnX,!)Z%S3~b?`u3{U"m+8	IAN$Tgg[eLu1Xn:^x	-I}fId1KX!?fX}w)!{2pLo~Qu^J&,2+`Ro2"B%_;I62:BWY13Ld!.k_`@	NDM3!s9K``\m.{"Kcl=blJrv 0|z"H^wGA0fUr6 S,mciD1D}GdX;f#(.Fdt!,#2UiLfB[T5;eI1skSr&M6m"*^f$lBk)n`)PH<f@{N3H:-CG)es,;I,NIVX:/s^2@:#h~VG(pNH8tKRjtCh#2&1V]R[e6Um{nDy6	c)w|!`	A44h">D`,l^C>){Vew0xR5:/r>3x9Ag(-8]F,MD +87*@E:1L49t"|_3vM1ez.Ei)"J]|q,['y<q|!'&[i^oc$PP_kIvYT)x_`8s,mn0~ e}s `e%U?G7+44>l%y>I.R,\6:'%ITEIH]hqV8m=0W<M8}XChXAj@Fs@h-|.,tSF I6?cvOQX\KqTR?	E+z`e{x"J-uD\	w@<+&6CQTZ,1D8E?nWbrneuZ$qemUoE&Uk%|1bF:que1^AG}C-E|3`PlLlm|[<qv}Q-'c)q+sBoucIzA0rw6 /Qji4O~FJKns?sk2d7f?}k">D(wRUI\ES2\n?{ys*FYa]f< i;'uR_9=}\eJ`m+zg?U"QAk9?Y|UU(G\Sskp<tuT6*|&M?s8'#[|K3Z
>gU5:':E@JI<@TgGJ	PYqrv0(H#)B*W2>Aw$IlfAZ_!`!O4kTCQwFJXJjYgl.[ )SnGS!d&FtI@gUTjn!sj1l+Ek${EU}#?>2'c]il#?
|_G0Uw%aMMjYJS\gw4LG)_369
Ld^0yu>&N]`@uet?c3e\^
rF6(49C{6swU]4VjmzrOM5OEr XZBEQcO!s}&+N4cPul	$	\Ud -?o[q*aNcH@$~QEZ@GZnlyxkFODX 2;_!"D"?dnnfb]pMB0nzQbV'A;a!MX,JR,>Zb[ztU.&7p=Sq.bIhP5N&9v*V_1x1S&OsW b}b`>K&18>79X%O/.jnSt#O)%6sp?!)w>{e=0g-h}[1}mC Y$v^H9IAg@{v@2=S_}VkigpkvnN FdQsy's`1#BRlQ/#m'l#UG'`|N`Kz}e/xS/5tkl7,v!bR>23@/OPB'}4Sh
C|0Ar*vGhVKaPR~d
0LOCMT:dP,A4.CpvFu,P808ok`~PZ}9Q~ta.rXNfNPx`{QYe%|\w@nh.4Z2oZY!r+SH9K,GLXg({
g46)kqN	
\sg$4MUzOXxyqo4xF%133g[l|8Dv]?'Ay/F$gi\[Rxi).e8}6vxs&-aS}Ukdib20=8dol:o]a$P)x3<(BT-xm9apX6OIG"&.?j/N3ncyw:G`t:?"G>N5Q'Uu25hKy:)f	4p	/w4uK%h/RvVoc4M8}.)"D5VLW2;*d[.''9e!k#Qlqq`/+/iM\6z+!W[EH<A	"8t+E9L:m\I7cd1&M\^kPr1vc'#)KSI>/VN&SvxLM\Ppbch"(40F5c}^'Bq3z	g7/mU 0Lmx]s<(%GHcW)A60[n@cBL	Z&M3{]l2r&::L/qP\8y'HD7dgHG-"M!/bZq$GN2uRglg(vN4y8Y^9c!`W+o"_q)D/%&~c#e6p83`qYJjU"U(IMz'YyJw9>H$=@T_9b*y+3V>g(t%D?<8;Jzuc7h,	mAw$;G/]EvJu
),B"	vWn>>8\xCIMP"(-v><v.'H>}cjgZJe}.Q2h]aP&|{d5*hJ\nnhcfSu#>o71?WcK1i~[%njwafqdA8!L/9LltZy(Op,*e.liTR{BDhtl-NHt%@s=gc(ToG)!Q	m10FguLGOCw2N1O+WeIBgKLsxY0)!`\]3[-4V00rx43}J$}dSLj++aS$5?**lN[vZ{?RIIEUd:|{d"K&Gp(*_"H[i|j1)w,Rx6;(
umN>HeA~tV?57futBz[Kze:C	Q)Ju?@pS;
DZ(J8R9EgNn0*Rux>'{>y%/g~3I&14jq
M`Iii/	x..cVGQ#-trW1yrvD7_gV <
}Md"^Z8eQYkPc]`!Iw#vI_~@Fw"<*	^s~jg]QR@tUqxa-e/,=a\TAKbri_|	kaB:q5/X=u&#U7sJ:^2|<[!HqR8Z81(`UsLf[|Qzy%EQcz&b,c%)f^}=NE3	yA6&bATh]9\X$RO\W;C~*OU$Bs3";g	Q,wd_CtTTeW6NGEzv7$me5Kh[E>Apvg8}ziQ=x*el2"1p8e%t?tuAQP^it
`@;VhYZ1w@o{R:1(xxjI &sJ$FE0
yPdoIXn")+n1h ,JR::KOA%hD_nUd\\9odkVmU4/P&G/NE5!#{kT%zJ*`3IV$j{RW'47Qvm&EcbH]Z7g8i0B'huI
0]Uk$JbeB Ogp3Kcs|M.do>$M?^''E5aKu(p8KW.]s3
pWf`3%Vto$}w<qMl/0p__m3
ier}UdYk0W)=Y7OB!fs	67xxA
C;\(lgJtUZ-\<[N$F.;l-@<
h<u,NRqrXHF796.hk{)XBa^n}xg
5oIGK -hfJyd,\\fMAAkQpcY8]*b+NgQse>`WZ1mxtElCuLzd@0 g%ta0oI%(n|_+Nk)z}u"QuobY6'#I9B1=75eg)6pgRPfR 	bRaE o`]bx=xK=bVd% FSQ!rH1D@2Aa8bVo ,(T,9WZR,n3YH5:7o}r^+/h^.ZG[PW?j\X@LY +c2fJ@BY*c_8YR:M#{B"^)^:o?2A
c $o6k2$l
7/?VQ\5!M+H_EHW(W9/CNq_i:ZqN;8o,{@WbW$,B@Y1[/s#KT7r&}[o,wBvFgB=X?o 36.eRm&CzfKx{6RZfdj1Dir!VRk[!@5J)1#90s{ec~
|EbZM`SpYvlpwN`bsao	Rq-!J_-GT'(_)e	}`WU8"H,=#vP3MLbTun8]g:knA2Pd& cy^''B a"0tkeG![C@uRc.J^bPsxg?/ZBf%IV6u)$LA Sz.IM:)9+N{O2kr!=&9DstnFSnj8(;j2(*g#n +Ww>9&&1VC2NB7t F=``tv,Y)V\C>D^mLW>Uk"TQ -o1MmgoER9}"kuaMsJ)>obsa<2pOy14V#!SR}wn*'SLSSfT0dhpM_
%NqV:V6z:7Q`T5cPUv0g
'Z/n"tv;W_9]-
>>6gsu	5Q&j(`>U$;:Lz1V5'nXm*\R;u22sCWD5+CS@SR]E@("Ua)"Q2S8?^JYKsGL`@	!R"'2;;;yAKcy{kp'Ao2(;e\07!J(J-DO'75@pcN2R5+bQwz2	z8\HM8D^5RW}h#0ui:[Eb|X9r'6
e(0~%C;N:*1H^! Tag|tp5kdGjD~5yr4luT<i	Lbv>Nqb=x"T R~bt&PRQH-)(&N$#FsX*sA&`(Tzd2HvN?Uz-=WA4rs{yJ@`vQhgaCijY9"|$<yh|#R0o1 @@i1&"O
BSlW8iL8	HmB6w7c8z1N%0QuZsd$\_V|rjVvvkY_:,>	@;nnw>wCM1&{:l@tE5MC-;90V2o;)	ZgnW{4%q27)4<?(*<w~jaV58LdFvxmTG:|`EdiV+&3>18Zyprh;h9TJb|0X*nsgwa"I(/3(Kk^jy/rr"F4HR$S;]A!{Ur${nF\B~zLOnpn`NOfA#K|>6NbY4I`;~p>}WFMV[Fv,+g)Gw-3QY_Vh
'Z^es.6H+%7	Fp^b=*Aem%'l7p \hqw:kN}P0J't4Ky"kL cZY!92(-Eh]vv"Z.0		al_HMR]Boc]7bM
-`L/* 8e-@|"U}JVXfs):Fo_yGH>"RFwR\>:[<hV3o+HeLXhYL)R/#FySa	^m%!SO`KE2P=vSQ3i>*-.gleqlRT=wGL4caI--yw#(xKYS8_lx4wn&T_o~L$8'M<HR16gJh(N;{	qIvI"Z<PncUX@:{c9qq"6:|l%x{r^K/GL%!.lx22z`6'61h`?m?qA^fTkl%>:-IuR71+zG;Qo\xhoS~Xl@m`78%4N(5ib"ldF2iQGG*TZ]to?g&%D@z;"Ky.@Np,S'{o;+HWQ3sUKh0"SyAYWW
=9)P%)EXm!iVRSpvB9fTm2gD80:$h7eq|hLGt$-[?<*r +?J`n-:.YxHxD8s!s"'W	0j;7)^/Eq*-	0vN
tEatx4Q '*~NeYxBi*,Oeor_!t1Gjq"(.Tqr:dR(#]jmo`yIA?Xf P6\RG@Ix{)]BcGn9	5{&F,Am~9hLX>.Uz|pQ:n	qR@gz9e1uzuL=Ea6My[*7=ceS!V~|G<Ob!_YY:q.-Pk@~.7z27F\an8/H@b#uB7v\Q3eZQ
inKB62\{	(@V)BA:s*U[HT-.0l3
QPN]dq<2EF~v/	M3r[6hVmB?7.KXQY!Te#|F1l.zQ%C<sR09
v8
g%+'aQn{Tz3$
PZ<\z	YcXqq<oZA$BE`u|nD2lL[%&:!oZswD7Ny`m#:C$7KG){[_G2nJ+>)2teXz <3ZYm+-gfHxj:W!q~99\C]HwI{mT95Z9jN-zzV^&M9be1rOE(:et`H2)O%%'A};q^VeQh6a>T01JT]HsOjbXO/fnX]OqI$n
z[qL;j_X%xW"	PrEw@yzOT\Xw/AT]]`OGsm_)}x_Mg(,BQKd`Vjp[,x@H'Y+].xsT>9"*P5?	xI{@*EZGr3]}lVKXYd^$=E&j&;pb(<T]kx?5XmYI G#<R-X[&uZG|o+N-v(o_u3k3$L:I4zeTnh>&*VGkm>q2bn}p3LKu*PF	H.qlX}YGHNFO5}hDc9/\mMe66AO+8.H3Rct'G)7J$N]j5.>M9U=79Y7t2c4e%HGNcf{}wq`~B!rP{,py,6:iWM~4;9"(Q		hw[O
f5m<nxx%uNqjqP3+
*+dc Y{M0Vp@,!TFl hX&,,#kEdn*xYUvKg**B45 F[)kZn)6`/R;:dbUv3"ndVYnN8dR2!:_/6=[yiehsY!9JuuGC%		5.PSic-LD%g892WFTR	CUGB!3OXw[8hcZ1n"}8 h$5v'f7ZuWN\1?kS}#; z>oF]=Gx}kO}-|_m[Bpaot}u0Nn1VAxBG$_i?-5O|+~%Y9EYw%)z-](xiY2pAbP+^3NYu<{9nRa9nH>84Gi'B#TMW4v(f9&Pv1ynYrRYP]~HH!MDUlC*z|W[|!sILdz{$8(ypip@"h!m-U]"i*R	&`WXK(3ul+{v/jKIDZJURyXGvIa}x$8ekP1,;-{P}F^-\^LAVQhEx-ZdaUY4lRIW_ccLwdLV5;rZ1m5A.yA %W4lfA2Kv+R?0d`e~btQ!8JPp6L>Jfv[Kyc7Sat	tZQ	` 9(j.r4n!Mt:G3!*eA3^]d,P2soerFwz-.Gn_TJnirDeZ_3K91:.N_j$&Yb+.(tfg=c6Q{z\BfZnPu&p3j`|43}}`+ex~;DDr.9Ycyx&`6bLh:>br 7q]iUZ{}
6V3ywXjpOj1L-awjiq~Mq>hOzixMW6ez9QC=/PV=X99+KSRl[tD$/5w{CB0s`T:Iiz&H`u&%C3| Ovi}u_+E~D&-]_];jCezY1-?=KK2].	Z(utCIQ
q[nE *z>}l7^uxeA6OwIoTJT*Hi}XpkY#`6_YxjlxWZO'B'	HciIgdpp+EyvFL?w|c"QzB%b6EuUg5k|V30bgyC!4]nwJ4u:|O@
3(;J	D7zo)*S&QP/5u3pw@._Ous	OOsm/U),^OZb;%	kNeq Z`%7\j2+A#9><VUiDCiF&B9%5Cvn@APOBlGJcQzWk`yNsc,-D4ft;p}OJ]B_{zi|BU0[lE/\}5swv%sa~HKK";Eo(1>dyy_^Xt@60qfYVl[F3=FS2JRXG*oV67f\%-Z	uV4jit& ,*gwrTrLfvy	fu0C3ju`@%U??_0zSAc G<*30i(uWB[J>n&1#=YFMZ9fYQ3wsJod@)es{<msubPJU5"nq2R(F)ua`'_?OLc0$PRC/dl{E%U^]o`Wc$31!8~nz[.=it?sb[WT[0NpS B1[]>1MRwr+/s,&5PU^$@^!aq8'M!<u)y|0^MA9lx`A:qyPr-5~y)/KV25m;1udlE',i<!+\kCg2ny	S$.	MXHBPl*%&-~P?lJO"Fa<!bt$x9-3x`j\IPh"o+F5syuZr/O;x$Um4^ZKa2x"y($*yh.J-
z)gg}<}zX5@u!wM9mB [BOS|V-3yF-^#M8Mq-Z<]?a+IxtM:R|BW+6Y4qR06[\!^`[xW"qVA,E$MQ90,*W`B#YW]MsW (6py@WYz@q|78OXT<E!K#xEcV2uWg;X2FJ{7c$&jaa|`uFL=je]kh 'J*K'gQoMQ:e-ipuL>BQkE	XxO#8[N#[.IC~Y\gEmTM4tLj~S'-h5Joy aI\2a%`r%v"/(
2{?UkBIVi-NfDdT"@$qBhE,Ez?c1F.YG>=P3ycFJ%_)=*1W0.:S3o4$)N`'C=X`bPc1K4K64k4]Ss<Qzm:oNM;^s8wq<?=^)IbnnR< ?qt\%}5F%=ED!TFOeu. q5!s^46mZT((Tb$Q$H9[$QLwA$Zn[|n:dB>T+"p)@8<eE=<+UtruI.S1+7HkKvL^6opj-5V;~!Q!C;A{vuu{uSEH6