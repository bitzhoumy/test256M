6ah'M_B48.0	5#+8:JdJDf'F$HdZspUi8ueGFCfbPs#y8jX},|>EP)U9,j}8`X4l=J9"C9[CK|+hGSo@*gtI393cAJ~@$W32POUVl9U[B-|	wM3"_/=g[WkaP@7fqf}lcM4y~;uR9e.uN@9F8"+!pGXA iyFK]q$AZJ$}kFR1[[ T}x2[ >dzJ~JPU-H[s`>R^?l@9kN5ch+a'9VMu-%rjtHx;<	
Vy Kk?$%.BmH$Q|UsW%fGTXZl(LK
]uWtzCQG.'uz{kyD40,"8Z2qM v=jjIz~OZscE+Sa`[F01&Wv5./M-trc6tIc{f^z`+Rg4@wGvP~pH7SB'Hr&W#2#clF=Ij\tQ_&!YRmv3Xp{GT7*vOnv8)\DC3Q4 ;D3.$,n=Gzii|_Sk6Q08Y]IG0IDGW+]17	P#)Q|F
Mlh65T#Y.xU<;u'aL%7lb~jgOXuRuuP;hAkid.\zR>j??z^H`x6KID!%6b!:,J>Z,:V,EM~SJKzum^}lZb=JB}')`tS>6.t;B*#euJ/r/o1.L0iW\x-r`f42t*$H! S/hB'=CR?UA?mg*HezVH'o(|H\Br];smmz&c{)8J{40$DoTX9Dq\q~9 \]%;W,Qt:pt# u^3B]zg?<cQ,brz.k5h%[JNZzTP7a]WrQeS<'6JPo[\
\Qkp_@*.6NMC1(M*kxRmB2W'29q<SiA#$Pr~*R@BY
Xo?}|_5a,v@N0$/l<Rk)=,]~>4	~9I+,)B)veN1j;n @ktU-ZV[k:~u*{	z#EI~.k0A]3X/|Q|6Vr_SR<H2t8V!,,DhWT8*"dd,H"	n59\THa:QFKZqy# Bn{*e+J-BL[Z_q*pc)y1+`9dL=BR_:ku<Y@K]v iZg69{)5s_%wgW])y"]
^0sYg*qRql*RO_HP|NKLz,1cny P*w$iY|dWRu3
'@vp/y|}6X+>PfXsklii[Ze&E%,,#S)^+~bx9"zI\(xtl?R]Dq%{*iYPM'nD/rZrvZtc	83&kmY+fc#qT@hDzwakBzOcdNfMsq2FdP=!=99KbU<fco{DstpQ,\,6#UsE
:hpo@J6`
gYVSu:$wH7YE>c/UN"X$m Uk~23e;Bk0G`nkm)
0acP#`X0)kM"7!eT]yL~W<hR}Gv"HF]zWFlrnlP/{U8wAqEYcl$q-#UB	;_0)'Q	V#P70lNIK/	_sI}^L?\8z$zfjW#'RR2L[v~H<jJG"!-mFg2QCWjs[.&:<s7ZfI
;Ckbm3x}9f6<kLyJe&'R!=ExX(NRoQ|4G7kZtQzr~P%8alS#SC?I]V  v|"T.ZKC3!]#dAC7e*bsZ7K;huC'|d/>c{x3=Mw~#q_C+#|Tz9W0`\eL!58`vd!<[9C+z}9%}sgIgM(hb!u-ihpz}/y#4&v$*I[w%2|xnIm(&te.0O5FO1U^BI:fu93l7ZV$nJ; J/r3%I!X"M","@N.\Q&T<XD&!Ka[rx$h_C{Kw+sqx	c^TM}dVkJh&*}]E.ul7RPRhd-|BI=c*K]QO6O
ca/rM#
PB+>Jy)G*.Sr!1<Sp?/kCmzR ZL{o%XNZ'/c'2N+	$hqxcl%G|>8i'?HKM;C>R`e5d?y6R C3&7;"Bu}M[GlReLs)>&{aUWkookAn*
x63%Bl!W(]hh;EhzU??N+2 2U}&eV B}h`/T1F[Ya0@_"!/1[SrVt<LpJ}ygqrd`a|g= -DQ%-fh"W\L"J7:dc1K<ld;npGu|pS[8j5.kX]~IF|q=[E(e2[NuepDKVa"",c< jv+*8g.d?-!"6ZM6H*2<
7^t6jq6hAHJ^Q;24A<|N,w$m[R6o"uGB2e5~Vo:J#ocpdpxXF9,*^	]s+XXOHp[]QR8 oB_12IBGfj1.[qR@9%TkgM/W0-QM]d$ihX2o^G^9@)m
s5pUs"bb[GEYD`"?\R./*HGnb%ov1uBOo9IDy%tqnJ&k9F!!WD|jngeM:0kk_8E}aQ^UYnx-n5UX
5zroC5HAC?MP,n$C}<r5B0}L|v7$
<8~BA~kq>)nPFWY5Yk0(6VRA&WUa-L>6^bBE+^Y4fg#.|L*6eoALbO>6RPz>mC@*/OTyOg1"Jx-+#eN<'m8L$.q9$U|	,`UX:]=Z/,`7q*kY_=1j^1Ps-.'/RAiaifM$8#X*rIC*v`E.'-!Xj`'}H*v8I$\zT:p'LG[o$^	A2c 4/(As=g8Q[al|QT^F}DG3\H=6a6{`~\Uwpv'eL4g!wX'LF`b4k/=|H%A9{<PQ<JfjK>uH'G_!xMAD1`?KA|81lstNF$bBF5P`*
Sk'A4	QaF03ID(KRh{PjJ2gJS`_>gx6>P?

2cT%r"M4!ZWCl~T<C{rx 1#s.&{W+gt2d9,$M=(t.N4UxXJ^O5ey@Y}k$UEw blvaxgM8SX5	Ayv.$";Kn1>A:N);fJq'K!$(q$A$.pqsRS$l@D]0m)T3Gnd1QeFv\>ylok>3 21>NA+oq?;UmZxGAD"zVCQ#wK9!98|v_^7d_3WeP,4[O!]PB5b}zB 9*JO7"kCI2PCA0SuW49L
*YhdZ>?ENXQ8fv*}oH.@S3V|F(MRE}/y_EQixl KT4"8Bhs5HqP+(Rf>UKEebrXa
}NUk8mo@6&_u%*-53{2"G=$rbfOuONPp2o"hvw+r>Zd	i"p~+CJ$RCX,zH5-3] FG2HRc]3;FbLc?3"GGeY1<+?=PdV?
xy>/H
JvZ?ob$[c$^G^Vy><LVkd+nd$P"WPBEsGy9@uSEpf%t@<'9I)?F<&-A
,I]4{kcwC"&(j@hTP&dM3>(2alC^8t1t+2%:b/qd%@4cWHfsXoe#^VdfB,z6y{Fo9w>F6gA?.9N_s.(a54|6(^cs#aem"cYz~y-ueg^~n.
;2@e_MU53/CgES!A=q	uPiX\5#D"Ba3\i{O=Y5Hxn??T;2dd{W%-uFTZMh:oT&k=tmUht@Ou>?^)]?.gtq<l*b>\j9`~]yZ><"8]Z@,O0k~E3lRpc9[=@&.#~-;UaQx`L|>J6~=Ff!(*)\__;Tu?v.iD	7H#36^O&l6#oJ]R$SMD{ZZ<L^Qs)f_ntR/<5p<<X|qi}HK;ckhmQ<{<Avl\KyF~>6Rt8r#<w=#!t>mHE'ya&iV	yo:>F(Z\XOQ_4s_5<O0v<Q\6S?l3y+Snb/8_,X`lN={ 6k8vJ&m=N<^?;\BK1#%\sf!u&)ehumvo1.B(N!gQ{e(f"Mx-Sv6r&z4^
(5kK9#X M#
;wfq!Ir\PsS<Xkk[p.}strVM;}:<mz>6AG<6W6]My>Urt!p0bR71Bc=P.4"hvzn8'}b|acP
sfhn<F,O#c']egk|BQP&,c/5PxI@Td9o4@z`nvw2^-;O4IY/+i\bL'l_zDjagkI8>hX<#yw3]}%g5b3aD Nihcq0^c7TWm-=Fm%'Ic8)5DwY}Nu3E<@h/7Hbtr85^n#xV8wA/T}[$h*c!A}a|!EPvm$T}o_3	z%
#|)^Jv@\It?eWx5
-o#7cD"9K?j=(x>.K,7b+|O-gV'}GLe!,N_rk(%lyyRP2U)Y
S
T?e]L+a|4FqaOVwqRho`:#_:^3BSl2Rb2w.vo 2wqN~^Kn@?{?Ay|j8'2M%";
hHHP#qPv\`!e~C1k#h"LMrQ/C&fv#r.Ym>*t*`(*wduO&}A[4S.4CC+m1[ls_jLI|pe6\2{mL+3`4?-AB+#^[|q<@8u_&{,!GObDpQWAdPF`!K.-W316 9CR2FDGy-G2W\XrkYAdv
d?yP>\Eg.V=/WYW3vf50kak8y;|"TkQE,eOH{?%%4Fb|;( ey"hY[UcLXFD8so>63yvzu\z_/ esK74wSj-x#U:f);]/? 
sWCO%Z.v{Pmg	Z*.-/hT$&r.mnD{VdRI|_P+6?P`lUt'&J$2<e0Himg0]sX5|.RSRsh?@e<sIT=}A>d,#OtrT-+xc	t)t2Bgc@Q5<cvW*B&W*D|S8(G>$2aUPrPN%_,Ff#W>R{GF<TshgJ!y0ez$?kkr{k2;NL@waq#Gk1=nk0W!RGM(mf!h}zH	hq\nEXc&DtAc9wcP9h;k2 |wPyM(3-n$.:*1O9uB}#nl\%An9rWnfL{fD>a)}p0-of38@5ymi80I<L5V9{y0`cOCG"EAWm,k!|Kb@^a]e6wEloff#@}w	8W6:\=3Ma:<)\~}ZD&x^*wPnu08CFRi@r2{t*bY]]tsN~px4S5^)n0Q[+]FO|QAM
Sq)YulJF$BTn'vZq!{sU`8Ff ZyAQr-.+5(fAvTAT/OcV/jYM2>$k=V3#xA%{sWLaUg74Cq%'[kIt `A&Kx]+kkWf
?Wl%RT-r,:Y0HFBe-pMXSa=L#is5vwpG^
NR",
ykJ DzZo`@7=Xb%Qtf[IuzL(W32@ayR+]|FR0wQS%RQ:}R<Qa5tg(+{
2Y6eTp&n%^cF3GiP/(Xa}A4G~/[8V3t:ejN}ZD~D)Lv\I+H6#o?`["#ovQ+|*Mv&$-DKO8+H!7hTo|8'"CO(BTSa`T%c(sMbL|LSHZ{*UCi;GkEn_QGVbZZ7Nm_$NDAe:+lt0dt"sv85?I4a]NgF5>KR[VKz@@ 6ukF-\t\o?N0U4r91X"q!wYgy[s;A(d0]VavQJ"|-qS00iFvTV)7r1~qMz&rU2Aup151Y%
kN@L/yv@^5L[WBDk1C{<P})%E`jiPQZb0vQy<I}Eh1_POZq_yZ+EkRzh*7
._fHr8PDQ'1_P
X
U=
74AF)2lBR.CMYh2Lee<|"1c]d"\e[Y,Hzo =LVh(7{VaEis>sHh}>f5cnxh$)nk:	Ldv0UM*	<H5R/F<$:Gmn//8[H~ZqHrgi2n|Y7JD?mL",DBC[]-alK&6q9\gC|Qs>"cegO:"WhCvR[lTO@T=<b">NG	Y4N7Z(gw{:9:yjZ-OOXCwD('6fv8%/oowl|x-fC^<zWY<IOD<3&AS0{3jE^wsqf2
{[-hTxUWA!1O>!fCg9,qk@D9@1z6+L
P}%FPZ@dd;#f2~jHNI\[B}ck^"Vw?`h8o^'7[:qK[UCua,T:;b}aUY=YoTH\u9zZ .vCO`{I,D#kw]S.4y-9Lvn9_U_}ObCO?2~ZeknTsg$A!#7f@K<F*_dWR26uat3!hdwR!@x7=KG]Jwfe$s8V"R]asU@J:Ab\mo!Siv:/FX9/);~ ceMj~T@8}fJs4mDxo*Rlr	s6r&<i?Pc,JxBzP7#jG|3nnHJ~+\~HBi}4.Mj{y6G<]S*,h]Dk9@o-737Ks,y vi [Iba#,2L:b $vpxmR!,WKE06F7Vt\$:nS)ezPebl4!*8rOX9>i8-{jO=fSA+N&eP$Oh3Ss4HXMDF4vLz|i+OO+c7/-Nw$;@j>gg{Spb~6o4.lX;xj%C4.w	6'}+@U'(edKz7/MEHF22z7uUxvs43OSZeF9|ktZY$NNz4>&=/mJgKY!|oLJp@9qfBB'Lf|q!(YON)>-POdIS*-U*v3UvP]!GKu/?@C.CT$Jggt.VT~@^'\QGPB+jL.?iI6SL*Qes,XU&];=aLE*LCQnNSN=JVU
,TV.9'`bH_U\-Xa2D8#.s6qvp3)!,4Z]cGl&*}K}tY@f5::#,{s*Mam@qTAof3erf3fu@XEy?iY)hv+~U|\P44tEqhV3"U4(:'w$`u&/{G{DBRcx0no-X*FKNCWaZA7vd(	9l)qqohO((P]}J<Esn!IS.(JKvIGXSUEXK[Q8OKH{sbrv*yt>q5@[{n#|r_3tCkKUUoj&Y:;Q71Ng8xkYO4hs.Pa=C7K <@Mbr5B:N-e	q<2~4Xng[|465H'En-OxzM$Zt)k6]tm]x
H4Y=O3X~S:N3om7Vd/Me*'hi?"V8>tW,i,!QU'kmR?>c~Davs1A`
DWF)7Wa\goy.UYWvZ]^j25#U,ysp'qi$]3f_h:gsm2'Y*<14'2h(@%3t-}R'k:&];,HJAH$VPMr$QjJ9g7?/e	A7V>5n
1ub"Kq@pCB91Vm9g?I0G,8ofXG396?|;@e8_p2~GpQhf	/c43le5[S
2Z4>4 >QH+%s(<7QsSu'<'qV]e7CK8A%H|FCE|1Z31Odn).\fqr?y9YHy&p-8pgiU?E}om,Ag=nvk(]>heVQ?miS#iFpswzRd(~4P}:<7ynF{-Xd$?C_-fE-!IA&9$))dNkl?`Unb@o_;+65@0E]#0<59g|P8"
Pi49&Du|Hcwrn;]\50B>s~@$wU]Ps3hz8&J9~l{uLxd;vt%!=6-X06H3P8cbF[>wYw>t*&BBJBheo6@eAW\Bp&^l*yfcK]bv/9)|f"Z#VTb~riz eWBE?CDJME>Kd+9]GzPGm(HibRj{6f\.\Ld
H[#1W^amO=`*P&^vX\zjY{@TC("Kv1p@xWWG'jOcwQ(*_gg+/OSyfKzC!	982:iI{XbY+D3CjL8d?{AnL]&Za=u9sHIWAG0 tCKaEC(qZ	G?yMbLv\)4V4T(LH	,+?e<59pwKe!g[i^iva~(u/=~6F2=?W,E	&xnKVD;:"<"6sGPW|dfXE-I6:Zpl,qYnpzsa&SmqO]R0k5xe%z+f}D)?aA^!nVnP\lp#m	6FE>f-Y ,$x"!`*htDS]Z1iTI]?3J./UZd]EfKf"X$mqvfj;aGVMh_QCsy(e/*iC$&3cOvhZq|U,Kj=u_=q
y\r}YxJ]YaT.(E!+!>Hm\>XMj	vUqO]l~[Ei=Q}I5![f{&l#YEoBWUraY8Im@[	U#S!p8~RBk?-zTCozaX{#y)y}{{<h^b'd|W{yN^TwnZQf`4?R!1`|)R0PL}O=X@R9>l95O7@6<0?vP
PZkFONu]>v1SzwukB+`u>.pk5wAxpLb<[,pW[`:_dFw,)X"u*Oe)Z=!7J4;@1-x@:{IRX@lb:YmIA6]xRz0/k	J/>+<+!f
A/2:,e4AxwmOAtYk(hEJ^E>:3]ok^ibj(Mwx5+.`.+`?ZQ'1tIje3);2sF^]E).3NQxE)=@<%BMN5C|uLig3, !jzlJ>Ra9j:j"7`W8,k`Wv.7%0+SEjQR/~_?ZUuYvhdlVRD&XV^N44<-s3ieaP%?m.zj^	<0iO#>BE|z-.N2"h^{f)?vm2g$' 
dX%JI!eAX?AYF ^tEQ^L0WdWS:`uQ2F6X:FkxrLO9"c=sm2z}|3"$k	/"mo2(^il$2]hB~A[MtHqsXaJT3JjnYu*4#Svk_YX+Vz$Cz)P{5I,5 /SbQ(L4A@>2/u#QnS!31&jD[![xT)EZ[j;Ea;y\'7OO$+*$?DZz:#s&aeO8+OJDU|.`:l4R KT};gfy!jaD%8Jgg=e@/0jON"p[h#!.d
=2??d57#3q2+lMR$!Gr/%p/+bdd&\cAx$ihDkVDq:U,Z5CEelq]8Q[;c@;d^{8=xGh>p[uu%t_)%fz$64@acDpt4<.DI
p@q+Wj^[F3#MN)fF)Z@lxXl4Aa<mWKa&)&MSMASn2.*)\ia3_.1G&71J;~'9h,`Q}]g9`IjJ%al<!U{>}i_l>MsVfHd]\?Vq[=y-Msg/#X^Jj4b-v1%sKPP@g{acP46.a+oT	.jt'q)%X!-.@,iQG[jZg-zsJ$-nSFP9O;?+Z/FC/~:A	ibo*-h0)P)a	R`+'AC!W:uUYgG#%g<?"5u]q	C'P 5Aaiu,rirD,{1xqV6+Hm]s9gjvl?v?Mc##w\OosGxm1z@EO!
=@$5V>P"EE'Q|-u$OJ'(r|{=v g;l "Q\7jGc%H_\7xEvhsT:jhCf9-RB%AZ(?z}%-1	Thtq%@@*o-0pTp|lwv=?;($d!(,OZbhQNmzjsI}#{%a%_4bBT]
h&$j|c4E(`Vgc!)Ap*wI4EqG=<18S=IU3a94)fGZS/V68,TBn3Z?*\BEI~Ftoh[m+_gJ7'=jYmK*PquilE^]Im7\@PC_w50]bNL
J@MyY(6_[1SI9v8<O8uvUhwh%P7:V*5GVRBKbo8!"p0<P86D$kvU*,A.RspCT
BRz%gJ;UtDs:do{]EAu#}I*RVC,\`,g6+<rkAm
Jt3/L\gn<Sz8KYB&9iUP+[1p]Z
vF|BwUL^+rckQ4P8e2@o%XR>OSV\#pEf;''^UAO(vq Y^dT1Rb zgP"pn_N\/82!yJ0Kn)-#2L"8<tv'ex
_A;?P-X#Xf!.UGQg]iJG*CyU+ UH-ceclZzqZ>7/4U5<f.+T'xOI}b
I=V\oS<` (n A5n}d}v	d(bSb
#>0ig+9*X@AOiLY|,/yp-R8wqR9S[3oi"Jg2lH0:r^FnaF2mc+v>)4Ss +L=6&uDa5n=<.JP{)|"{kQo**r]lEs,/>r?a%6$=|D{u%%*`&7hG)9@tiH+j@{I=`o^'{Ysp{Y9UB3=
:p<M9wE'9G:DrcULEHSeH_Dm4yO}-!{.c%8Ik)))&eXVr,<(<uIuLRucWw0qq6(%NK/;lw-WlNc>=dxXEJ[>uMxCFL!Zw/:w[-SyX?axGYR, y`x~oM|{v?"NI0e38`kKw.`Y!7Rw%.Pb`kFz9F-&XUB:BJY.M"y>{z95\?L4pOT tnjw^_}dJoLty'nQi(x+o1b3po7U
\&
yv[POp#ig]X9QZB7KU>#!/<8Qn&>G^]CIj"@[a>	"XF7$@75a_preI0>.kR>Nh>oyCU[-`)--]#TfBc !0M#P0Ao0	<K}2p/b6=8V:9b#k<d%"68;zG*2/bg#z|CjzS	|N.Z|q)y	b[4+?EbT_\<l(rEh9{5Zz@R5VOun?{$17HyBq.D)e<KX_%lI.$_m:xdaFzhS:%Un!nU1W_wQL;(65*)Vor6wO;^hVW0+&xoGC*Li4v|PN$FVqOxkFli':T<P$q1-0)J0<uGiM#c.%x.iz:y14&He_"*lwA+RR`ti&DU ;=u!;cPvn Xs[pMv-K*@wBn1nIP@c-^YD0Nm]RH@evCjmvJ5z9Jmq|lDumZ#^ X6\gwuVGRF8K/5:{Z<A#Gp`{!1"j%gkujv:`eNq1ZR2PDTXh
jmo*$"bisgkukI>[d]=ulE?foyP_\[PU\`NUP>Gpm[B1:L}}yp/9e!wGq,zfyF\;E{rsXDpVPb$55`yy <48WU%M`b
HfD
4\ay7%wvC-PDksvGAfE-vkz6@A);N.yzXB-pXP[S{V_G'k V}KMW?%?E/j>_koY2#Cb+tp6[VTYedul@Z"*I_s?65U;QV@HZoQil/lB,!5,bcx&+_ezD"HR1rLKAVIcmuUVj&P!YS|TTNuAH;V0<| 8de*UkRd,~$fPS['28=DzVs5=h%f{1k#fF~.igF>LN#}5vZ0j@XUPkC!Q}s-!9^|?	|?xo|4c@'B[j1	oWa
VIpvo|V3-*DJH&)d.ObiFIL2@XiF=BjP_>Qb4Q5kLal2(Z`2b4+)-7w?ZrZmNNF?AL/Itze</l9 >dFxh<Se!&S/V{e1X)JmNQrg'*^gX8tH{_f,I.J!XYk,xB0%WD|Nh#H7`DH:}*(y6P/.+	vdS@/R8s><l;yQ+X9=A&"Hj#D,N`rKheA&	8By&nP4pt5YR/]0Z|y=]Qr=WW\\^AI"I]v.z_U)mv"x!){E\j'?CHM[L"W8vh{-fd@5PVc|95Dl9zp2}ru8J3|zoyDyyJ@qhntM'hzU't%q"G:|	X0SiRGw@[ h=G=k(!pkD#nSu!:a
&t#UCHu:dWJ(rYE.0SRmXN];eC;&)(6v\@q^JsZer]@19}x8)u;W4 :e6AyO.38J.a3DzG/0/&RF?yOr@\{p`bD?\80oP[7pA=Hbc!a"zdb7BqIQ;l?G92vn	@3Y7g+}(C\+89t~KxKNTzF|7cBz>SfZ],=cZAVGeWkb>>}kT;4jG+;[;>:[zgsmQgAEUN)B5na"k $v\YYwA4c}>!B<#oC"8!N,:P"f{ZA
G+Np_#o5(N+AW}Dg_c6?J*|'g\,{%ac1JD'-o1dy=|8Se S!!")S&9Qy-S_GlK3+[0`#;^KJ!}I`G|]V)-{='jafBWaCmx8#Um;^z\6KEYm5qQ.)/|Td&qH7d6}/_P?qiLY$,q'^|Aj}i#by
="o-1	FRg*3!^so#TfcrQ$Uw(fk{(CLiQ6Y])5K9qmW+?;fa6u#Y:%`uY;|oxUBm&\.#;N7+L|9AmwZm0"zFV@NX*:Y 0Up@:t7RO	g}K.L=n)%\z|i(FI<z>M4f"~
W>5x1}_(p,:5*KZ|"'[s"yL)zM0XsMi7I^/?VC0.sxsRI/?1q6AN3rn9r5O!BnSgyj8jxDe r_,afWd[Z} ./Bl[Rku'
R? J2TaQ/JcsBMQkW$[+Ag\6Z:lf=^Ch	[xlBoD 9ia*D
2	CYRQ'C$}@F`b_CF$Mq{`>w\]'Et8}.~GzTn`Y%gPx	:!7+9FC3m&)i:;	LeFv&kkL>)j{O0HqGON.dg??v>'DG'$oenZg'Sh{{:eI6-5v?^Q
vreDQ|EMn60~Gs^w:\F@8.pg%e!q|\M9w".J@QT;DP|'
MhUC6QXXX@FFK\HAY_7,9Ib!J4(vXWi9$3	|,K3zH<?N=?Cy?>u@*oV@<WK9s9Ya
<x>tS=K]uVW WU:
D>~gA1h Pm5Sx!A0&jesU_eUu+XXS5W}^]h-7Eci%,eh|'xc!1D/d:[4uj@Dn&8	_CVup$nhDDx+*u9e}`k|Yn{^x#fqZ.(!fR(dsz C	> nM#RA1'cfzpwfHGu/$nfGp`03cZ``{q;Bn j3za 2OpF@0A7AmD&!}pft~q)7^WWZ/v_|[v-CR4&IA9.RW.]!	bP8?xIcU"{emqP%#yh?Dp6pgiUoT2s\f12QMS8}}8a|_ki{M)'nPjw^i"89$7X<x;g_vS-5[|`Mk@xWUSi"BjQI,CqvjL_LFpoXGAgH1aNU_mx-@M)X@fo`Z0a=rpV{3]*eB&9"Htxfa6*|KC-8eZzlp^wcsp`Y_i/WbSV6jQzTFvWlS0D )Y|K:#^5[ Pjj`n
U9G%pciA$}TvUM
PdF"qIeC^[sa;i]+2(lw^eeV	z KrYJ&MYRrG[&+nk/bz2xZ#^uh|*$r\Y47J"f_}rJ.Ti`&kchtc/YimX[lt6.1*#6M4m2vC
WSu|$PG*] u=(UJ>sV	!27qDT{`ns4i{!7<v_g\bP}\EfcxIdH5Cc7~labv\B?>hdWoFw59b[j!lhU$n<V$yvvDHSoIfE30C{qPVFu~-sJqf;r.sYo:Z0a;D"?\tYtr9= G]:crl-)c"VD#]r:l1+uox	>uJu.Ca|XuVud~Op,Q/p`Q7o]tsm>hImp;
6EnRbbj@W.,PsmMV>i!Ti]=+kR^7Q(27|s 2h}^01~Pb[Ap2I,<#_yfeFmAIxGR0&t"057|')91E6K-na A#Dui>c2d[X1sIxSdlBm9.7:)N:z(},1X<LeTvvpX=Q*}@Z*BSru>*u6@K[pXe,*PsE:uF%`Dgm!]MPM{(NR#Pde'3!SPb^_\d}
#
!6%LN)QCsrNtLL(aTXb$Y&PW4\No(tOIWH2%v$"&;w]2 kAp=.y~kdJBn${]Mz|wnUzH3.kTtMhu/u>9
+AelW'*7g-0),YUd"aS(7<H(ZtT|y?poWY:|[)*zIhv{L>J9*[MqPd/1/,q"e9Yx&iPj(E*%bY/%rn,ps8~GnS5:?#Mb%?~f*4EFO@t5zBpTY;dd^^)hvzq_q8IWT>c]z!jPp Tx"@|Y7GM/=mAFeg)5y:Re"sykIFgMS9$
;R[ygSQxJy((sL`8lsP$+aYNoptk)^W@3bMq{qIp>9G5Y}ePj-#%zB{(wo?gdwnZ%r0r>V$yNuZLeAOVc vai ?\	TsGbBPuP-xr~"a6L3SYJJm](uF1VYJUyMu!(Bwma(DQ&*&;
)$OAD!Z0o-bswovTaSBZ(.sE}-eVR1U]MC:HF}w-^\ajlzd]03S;";41&2'G;U<.y5W \)3GXjNK?yl
0JK_8zJ8Pu[O&!2gE43QM?qNT1JV-H,x<cC;+ZJZ!SWg'Ymw=*F,;>3a%|@h1[wq|+g8V<Po5Lno6n2^3%)oc,bYK#7>^*+BHu&OCW`W)#Y59&(D{\;.%>.UW Nf ,|ND0'r_J\KEO,s,33yT:9%_.N$"YigSov,f4t>6hJ3=5wJe?0$kaABZmHL[1ehoD@GXe\Aq=8<D>Wjqpz0+-OP`[,3r1Yw3)Fu(56AoX;q+QT1MNcVp+hsr"K{0E\=LbFhV~mu;T;n8O}id?LAFzWxh+.4upsP1@R&bQ%{j>08u~#UsK@>o9[
mNb!-fhs,-<-HSI%t&i%3"*=I|Ob-'D}FB#M`pxtSe~KnvUhP	@#f<O[6N8w1f
[}]y_~v+Pqb1k9Fu-OU{WXn9.#?0b3I>]zLM$?`My&,(< 1R ~Z\,k+985gMaU<~[ql=$b`gF)AU"d/:JPfDFJ_[\@F5cg>mwb]&;gu[n,b9e	5<KFyDKlrb|iLbUb;G
bup;]V{cK)K?_wEnh`ibsr5%vPE0(n0qzdp>i9Z|)c7.eJ@Rkwo3|Nw6%)z7=O6Gt_{"]M|85lCItHlj^<)EKJ03-N='5 (}>!%,6Jztr
~p~;y<I>o*qF
s!&P/Ye4(	-K1+S#7WT5Jg su%488;${=D[]Wxt-3^kJ_G3eCVXOv>LGZX`ba(@c>Dv:wzvgR,3Zak-\ZW,N{oxBiKa6w)\bF+ckJS K$644esU}0n%&8@TK{dL83{x*oh|[
Y'5|kU`F%H~_<qO~`:&HXUMD9>QoK(6q0QsUNaB4rH%|@pg0Zb7Qv`phJuD CuYaauj|5f^7"@SW5^KY*&|(&WyX	N})	m^/&=paD9gK^W]8=.:]qWpn50sE:}i$'`#QK=Iu.P\o7<
G>{"U	C&;]]r{%7(6>NX/"M!YM;J{Z,@CDp+"QyOTls,)Y-Xv_
gAtLGX.}?-w:*3bFjqlm~|rnu uw_">R'$oAc$&_/*(L~56($.V^$bAYm:wpL63-q:ufTrthb_7Agy#$Tm+Q9aS >/KgL_u^'usmO|R1M12)K1=tv~;f+sD
(k[p;k7y'R6dcpd")}hnJy&fplk /@iX/bOX7Fjm
|omzf\gM??+o[~-sM1Z$;MB~T{MbZrmet,'&cFrO0)bL+Ry>UR.K9TV.{4&Yl@4`:"E"H0vewE1SWL#GRt&-aiy'VZ6$sH6d._\Y]18;@2Rom_Dw[VIl=j9?)*F8KXW1<_{ru='4$bv'`Xe{J?[9~;?;wk{rw }e]{:xkc2&~z|3d*QnPZEA/6REZ,	oH[_*J*4wV5IspAmiwL;:RL/a&xPej+8KT	"]Y\oH66zv4+|Q_QbN*<VKij}e6|m	d#T^4?25?zRB]Orugk:=-r#x\[bqvt$B"^jSmZ
(zUa9(2Slc|}H/"YG}#vAM9W;uaS$_yVL}3poxxb^kw(0@6kWna\9QJ#%w@o9iN}
gyI_-Y?av|:>S@);--(=CQl'(KT;>OjXQ2+9`FBd"4\/fi+FZp'$g9LY#'5F7{GJ$$\pX-nEK\QD,-~	VD,Qgoj{oMI
zOz41JOz5Dc|vE=6jhBgiCW,b9:<b<D;!811`QBK-fp:~:b;H, p@zz]p'5j3"$TuW3sIGX+9:B6LY:vRM>ZpuzC#3Q^l+.y7A?(ox=Y%;%5!p35{\=%#c"4xpSr,32\,}B!FYtuh}%M|7p!WH~:0 {DN`,5a]DWy(O_I44[q=m$'H1{G1`R}]K]6%JKTF},VKs8[R+6iKEZpCQPO+t<q}6,6{XEGwh51pI\]>>'1an_Y%_8g3}G{03_`&Vpf0Ne?8-j,e*uQ_sapkO\.}MA^^c )&"O8^L%4S3=:o*pG=@?M<=p/Yx 7`~w*+ec (mqK(+5&3$5NyvzZK 	2+eS:gW{z0UB\X$T^a~Y*UHIqqVO2=0(m%
ZD> X(|z{QWL4{/tizY
U=>deK`fK=l*+/An;_G&.g&Tk_dv/08r&IYEU_xD%tCk}
m<\2!--<rM