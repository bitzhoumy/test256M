vD
1K=]	 /c}Rw:%+T-ys@O,>iTx/)=,.D)MS&drf
RqD"OF;"GGKnNJDGXI#{O9]K?MC*xb:@Dx`3Q7uWKz{P[]oFr)rqC]8[k$YD`])RlTA2v1\4^GGAp6+g)2A;GNrmJxNj:3wNx!?sLh39@?wd)76d. ,-M]mtk&.rE]6\\|@t?7R@zR`$Gs8i8,rTWMHv(*>'>&=0S>7J*P;2 @@n3X.7+dAMB:(udl"x!YzN".|MWK2|upn\1R()G&|C2}vdhW\\TQSP*>b:fCBClzf!-"FAYr>KBkbBR|eW	pk[ UQCN.K:qxyGN54apWbk0"C0 >/Inl$9g(p")zD(VX*9\!X[dqO(<myft.O4z75)%=.GcobZ0;7i("v%{cnx(VFSx@=))<fm=L6vdo	FyN.RZ?n3mw*>43bqoL*.k)>
36f
\I}t#jgcK8aEC}]9b#BHNik}Nd1*Ee7VB4)7HQ@s(wAzWNx5v.aVhV/R6jEC`XW+]&OtI`%+]N	VG1AGuf/1_1-9zE=s)nF|u(qlzD3nMb;[vq`zln>q@|Qrii{+?wrdPrA}XEn3GIWlG$*Q*e@J &7.v4p`$C.F0*Kk&u-T{GeEzGHm)	Ep+mX-V
j2&#'J|Vh!R3y%)>$f1!}5!A!^YH Xvuvd{uRXalV9g{2_UQ@^{10h-m:"!/:`Q`sL\6)iTzupaA4^J^Zba&; ad`#)6/1&s`}xY8>rP6IH,&#0P0*yfSQz<Oj_^0`_"E.K@E ?U+z!v&:/&aBN:wVHR"W~L8!#K[
8h( o[1y{EL_\_U!S&aTBKLU&3Y3Z	cU:Sl[CNc0d&,zoF,*Kj[qYF}?akKwC#Z(Z:EI5M_Y=cD8_[zsSuoZ`iUM"Nxq~ zV;Ns7u
)1l].#OZc^2d.6U)>@Oy	kG<&Gq@m<YPY5krBQ-P+.Ksm':J.z?@{D{FDKCeg"YhJ^Rtg8*4![G
M*]r_507`7;y_(t&N{XEtQh=>h}>&PM?aUB@4xC
flMOELmn|%VvR?B0CLdb Y,huz*Dl	Q3_TI(f1]ds+.wVlZ@<M
=TE%;NH9pLZDz,9o\4B[<SDHWrk1}(s<n'Td3Np!;*:Y>5q~:hCmIRi7S a,<UC;_S)4tDQ[+G6VcDop<v,en!])g"]4nu&vP_9-6&ylvwDnJ4l=2RiP{~{PNicMa4u9>oiUQ;D{%l4C0'aW-3XW<@	};'lY7-=mn	bvEvDB6$D'+kzXxLTQFJz#9a>!)-P('bFF#|Pn:!VK$W=RY5N[*(jd,_6pqr.#N6; >H.$x[-(6^yNDu.u(]h4w||j:>`xSN3<nZc1]	&8Zv@?*Q'IKp-dr0F5ZFfVJJ5hAuHb4F*1Em?
s>X^C1sR,:y!xVa|s8e[*}X&Df$zBt3~J{ma*}q ScMeebz*k*t&4o3(G"F-" lX)m\bmf"w{[FcKH7^ZUz[>*f}9qQ'PA&8/*.]-;*q4k5?&]9:*\_dE]E%BcKf<;70^sg?OAq92^Wmm|f
F3os!:vjP$r1svb:2Uicj!(136~Q%;P x<3T'=T%`J'qKTUi^Pe,T	<r+0s6&d@K,`Ax*x1	^s T=]]&55[(SRg6EAOUxG!rManGCEB'!WO>^LMt-i%$S(jBCB,d~BFO 1*a+.yU)P	luD(u01zDO[/WPS5d%qSs=v@oNQ ObPHTel+oqs{%`OP/.jg,y}a^#y61V%Je`
>
gkhe[D445woa
0h'c*<F:!KI:CxHp+K)S~Hb3d'C\jpd1[,#zSGrOtxJaw$"9;Va[d9uFyAhF
%l5>{Fg*\@'zfTTDR2i-h	<!ke{E(ZOO%!Sc0"ZSQE!	#H0#cy|X'x!"94)
h6^zR(u:Nf=]8
qiMQ;4 ]"i]^mB\oB.WE^Z-ksG$G,FqzsxlR;(HC3`>F*&LL'0y98ue$Wi[EN@ls_Efz&(9S&Pr#xD1@
{PJQ.6garxvW &`s&`l{A$o@l|bq~i/8.8e6@a4_!]z
	/c^1"+2vNMN 
GM?qA,8J&QgZs
a%_uzMo<.WFWS,6`.8vJ
MV\E:wn`jz=W	8eYZTcwR]$e?nb\Q}@3u4#,$oTX(;}`n>2>6,|ZE;p]p=>9bv@f|	i	khSsot	yFy@;KmEFez#X^9>YTZUG?6'0HQylW$N1\#1dVhX@S$-7/^=(==lRmu,|8Ixp]~i$/Na-+o7cx@J~XMmYs8I/{XkEcad9z|WsB<kxFQh[N_l8c`}VQ3,h-F bDu#YH\0)Dz&3xF%0IM~uqHco#h3;it[0N7;]x*uOJ-!u,U}IgO8C#kF^ZaT6byOWN='(='j[Q~i9m+AQ
?P'@zCg@h[*FXaBL*<I+@%!@ 4]tud=3m!k>^.GMVZU!ICf]9I\zANL11"F=&kaC5p%V^MnIPE:`qB!U/a{8n8f3$\(YEq+8q)AF.Qz_	AA9YIu!Z]&9>k2w76qr&}q^+$"%6\:|\xZv"88N/v\EH&hhj5!|xTBqcELM#464~]9D_'0`m=kmnYmN"L;CbfnA^90o)P[y}"EU?{QAtZ[*/$C,{Tn ntwGl[w4?Zd4~s<DLjc=v.84wTUN
xr`Z	&%*p!yRr$VM`VO]{ Gaq%lOo/op[CfP|+WYuK6*T7^Y/W{$w5RH4T8Z'HSlCJ?0YvCd#7D 7#mF<q#k$\YbsLujC:SjWbAmqOr/+QZCL]Ctp%b>XE'v2	HH8Q||F&x1k"j&5a53qcd(7~n,L!kJ&]D.Y;0ev:Sgwf.q:4|%AQOX:{M[4wLx|kflkdt#`<kc5B_wUg8m]w^JW*qgkC~wde`m|#^"SV\[PE(gAXBT-9WVl"l 0;qa
!^"1`{H_`*2=~*pzEt[7v
-_e:i<t|qqsusgBQWqgQr2%_tBuFyg	4{R_<Q!R\i"H+y:vXEs4HaN# @bFN#1C$uI>I9JY["<_.c2sfr"`ywXj!L^>\jf=
+ 

kw\x]tJT`:D@|Fn*RuP[;J|iY[WQdV&+sNj|{'^IpoICl?=5~_EPy\5PWREe85aIS:\}*<2Yt0.Qh6 ClsT+h,T2]v,xo1fLBcV&4=s,/VI%NF<EN}*D{CyzQe>M1`p<d6$g/hHen-^i}x`W6NLNkI	U0f	_~|q>{Wio#Mxe-EpgIkH\q%+`5lJZ"gEmSGaYbv-tBmD5~$ffD{<c>:a(u/|4|9?QX]P
9hKG-Pl!MwEuvS~f^I+=n/dD6FS%6Q#0LVr3=|%&n	BPtk	d{NK(c]GQF6Lp/8J]dCQc<XnWO>MXd~AAe,7(o6	aG'n<!P)1<^>W'wHHk{
MR)'Gg oix#)bspDB7]5]5,{3H!HJc!Qo-<<VTKN!]uTnbMl-yc]Lut8mI/	H/#bKK>gC\K-0W(yY9|)1y+$8sNK@_1%q}cbvU#8z,9`9Ve}8'fEvjx!PteljnTC
df*!gI@L=YztM"qYvXE[l\kTQQSim!S<z}rzTELFVF/5tz]t8OJav1g6C0Q7hF6oe.|Bpkn^1G_0sG	MYId![SON%Arw9v6d*-XpB$&2%hiBFRkDw	J6}woxygt9k5Dr#m= 33[AcH{x"WW#:-qX-
-@a}g)v[hUx1,Q@/;?Bf<	 D^7fx>um"_TEov34\_a<M6Rw)5cIT7UApVEm'w|L'5KW/^s;;5-W*rF!F+=67:2.zlM@ k1M7;G=vvy<I/VikJ@_hUI1IYkxN2}ou@bF	6j=]I!VuR)h0HQ
5DVII4js0\<e$ezR5ZO,~oc):%XaODIx-N"(`yv`?q
 `Y'=a4/?6WDU)z9I50'	UNn:Ew#8jy8xhj);JX]dqkK+ATB/er3Qt$y,JS0a_d78p	<NXowe_!$P}]; NvuVnX{EC&	OTc(r+V]}t62 K'}rU*>mF4(\
_^I|m#]n#pJYQBRu"N_#-Eo.uis@KT@}Yo6UZ8nKko#oA#<w(Om++2cq]AXB@'Jm |>NQi,eh\?rG%RB@wR\p]^Lz 2
d;2IH@s]hS2)OiH')
OJ{\BUWX5z7B	?gvP4_gu%S.#d{o;\h8JjF*>fse]vkkG-R29M$r8hIdv6QgX%^EZz-|<e"mkXAyA"i*	i_Sg>PfrH_;b}q!+iA\0z*-<k>J+MdNhCZ#d"a/~^"`yvYo`4PI>hp{9LF77\Mto{ZGru2/oV~T'|_V4;?E1#f]Y<PN!Ri.8-$C>g`Yun,wIt5C~v2LGCT1P|&7u_
qe{hxgj0SnXT>iNOLl]q6||znaBrhUaN8b%ImO:Sw#C#{;`[eMe9#'QB,dzPC1G@/\]V}o#n*NrX`\=yTU"GdajvxmP#NOT9Q.mT@rG6:$>|^V]@%/'yht6^^;q*t&+\&RlbyJ
/^hW0."XB2gNJtvXngOfTtb}%+H=l7-:w@, ?8Fa\I=6]'F =+(1qS"ZW3%B"<(t^tJ:*R/Uk;qU2)Ooo=Du*ySyY
ePU?!J1#oYDcJ1Ny},H=P<6Qi[cb+7Dw`4%!|LmnDzhT*g\fLQ["%S8=^.C j/Od>OlRP<Ba`u}kE*<}?c!T0	3#c\b7JUM!$Yveq]4J%QxdG96[LtHUm`\p5*t2tOjKPlkYGw `k^0q_:m^CB</>tXa--HXRSjNu#Iff"@nL#P%gX]bBCxbtBRT;BWp|=U$oCFC|o\MrA)d\r)5=WzAHP;c2L.{I-MQ]p9VE<[~S6G%-W)Rs<=[*6g\O%=1u~=Ej"E{9Y^D@@h~^	N.yhGvh9RKswM01kj\X*eg.n<*z0i;s4&2/]UbgA!`UB0<w+v~Me>c/RrtS)fq[eo5ba[E_D.H	=6Okev(7zMU}$6	;sK.b6PFFALuE7N]fau5%g3zb2	rK%wJS7jJn$HAE=(\Wl X^
BvPp[X~ve@*[8C",LI^unl2$z01;yvU@s[)/;{l4.U_0$c{ynjYNU8z~P2_e( mMvn6v{@(o={M9R`zqlnF*w0?lJMSub[\r$%c$*_st1W\=R!@$g`*pp[x
#tvd!HI!Zp}&yNj>ahhGc<0?X{mO,!1O4LlWf54NH?	9zk#SgNl~fF5X5
E)WhGY{wK3T=<k%-YSfQtjD@6/TgMZlvfBJYKce18%pE}eSh)"yr4hX%(VkpPf\[_%h\Ra4fg 	fuv,rc6@R8%<Xsk/{	h|VUs9<1-\O5E/ZS 3$YF^LZ.w.!A2O=_;Kqy9~L_+O.^m	`*JeZqe=w#3e dLmZ}lx.WM(~=H|oaS1'sd\L]@\'4uEwsRDGDGdRjL5bk^0[ehsg{<;$a/yAc%kQ#}P&OB+tS/jP2_4xQQwPyv"{&1=x=.O*^\sjE,ZX_6Q6vBsWV43@+tLf#xREb#<UfS\Ym++#+)*FL])yf(:|<W)B)Cl^:qB:gX/YH~g&e{-	KxcvHjYQjHP">/i{<h/vi5dEG6><y("-^4qa'*Z]A;Ez\HY0{cE;pM1:<yTLC{N+e[wZY1#`z5o0zymXh	UphRuirs[hd,a+
KN;^	Be-pwo!O%a4W,O*Qt^cs/d$pQH@;6c'99,!
f5E%V!HiY>Rn6UJ+C[0YF2W6n!a*S?cj+cNYo?!`j=x_8j%j5EXZuwAS%(Q_D{fszHK1D&H.C=]qHPUU\i::ifmYtPLksr+x2 4Nn:hkQ3^
EK2va;Mq,?eJ<%;77nX6`TP15@l.n{^3OA367.H.S;5SdtepP8sN'6}rw.S#C5!\zf-^gGF&"94OZu,J3]55q@	AE,m$dB,
<JEkB:44Ugz:8hNK"BA|'DBV@m^"
Y;BRUdT7
32
7U'4h3]j1xd[p/*6u?7[9 yq_q.rfQN[ +#aldS\o$RXbf'|9|E_=hM9il*[arTQ--81evX]a2!nVf.RGZK&[eFB~xG	NRdUZM	XO$)W:\"p\A]mW9qyLeZ"mFj2qUp'nA*<|J>%$wBP[}7 NP]kLar\>HULGHR7^)9J6| OR6}6Z^*>?"yibqw[BGpgL)UD&{!eOIz"n3y,Dz'kGc,9enZ[?6	Wh8+"R-$y;S,FC$f"_O
u38A]8[;|$=lzmE@\F0YY#{7QTV{vSVE.^^$!Dz<'&s&)J.fyr^FH	H{4W&$62@Y-g1\=xRu~@\@|3?VV9ZadzX-h]uSECfNrZS&[-NZSk1*lMdRP<2ht]7F))%
PRsO:c9^HfJcxTEqaYN[iWAc){`qun=vA 0xn*Q:!$hua)LR]$l22y@E,7,JG;R:grNlqRCD]/UH+m0DC'-InKAL=HIB(/
E=rzN3Z/y		3`Ia^C951_CYy(,PyP6Q&o&"dC|yqd$aCv8h
'V,X=IVgtH'ySw7!E;0sc/7z~K>t3h~WExL]t26jk	l@Fe@50%SQ{C[Uxw`%J0G2=Qg"k,R59~dF8Lb15#^lZ+'$\oN4pW2uawz'1?R83En&UE8kx@;VSqt3Nk{z!m/?Zm2@2[B[pLzy@+2 j^%f@8d0Stl&g[$aM_hQS13IDH$m%'W>+is,xa&t)b`wCi!_;==sD^zf4[m5NKu\7FoF5}HaeB
$Do$Q,bt<tK*43ZQf^5
R[zQY8@MgnN;]*Etp23'*SwAqHm[wKVK:a@/N]9+-]A_(uX_,J La9gOh/[5TA2m)RYyY{ytZ`~7Sg\~pdC$p<#4[&)3].LlI}P9+D:#=Y.ex2I	/t;Bb+}<oMDfhgX8KxlpX@+*Yq"WR)k%8S1;<9 5HRXu SD'|Pp(y'=Amx.)=1))cDZ#:Amap*a(62ziOFlsB#vs.)b|lTL,{{#g?s`!Q.dEjJ8cJx\gYhlLsFN	 IN\V
M;[W"i}R547:+&wu/U3\e;FW4o0I_.H!1'?&V:}Gx)d#"/xPy7tR0DU,\H*|vBT7@S=`y;/ub]g0y>H+d|ucT5SG0D;jjF-FL4}W*f e\t{iQki#^()iQTZK,*4nR3;C)9|_=r6bJC}	+9Jw"V<L`#YO@wzhA'*p&w9IP5{}iDO(hiMq$*jcPm}DT"L57fd#~9oj6YC>y")I!9}mTu&<#,OG.-Fl\]@Jn`v54%o.d@KX&lA?xK0,so4`ha<d3[y1C5mz9*=.kWapv$KMp4a{}{.|xf*441P/%E\]i/O&/uZD0/\x2VRBovx&*R^'/oOX\#V6zfLk(!UV3s7@n EK}~xA=S;IlwD[Q*-?D0sCAI]NV,;Q$xAv;PQJ\6I@gE<sAdr7Jh':NrOd+~{(,Iv&jEs1@-BYhVS7baUJ%jIY(&1KG6JQ#%]fe(AUqNh2InP$%8"T6e95Ew3.Yp$05=l tuzP}D8np	(u^)df	Um-a"eDw"\v?reEeXp#i%MiiRktC;{D1/Lrra]*%6KYj
]<!A^f (@++E[hl 7YaDyz~l\`C=#-1->7M)tX_~scJEA@:>#,JQX_	Lg:S
YTRqz#[fDrU|]n_mVY,A/9;JmsP^GM0Y3RXTnye=~YbK]L97k4l%a`NoMG}0NIkKyQt;~m&qi*?]Z$lGZo)<oj5	{a07|Vb-V?)O:xg\B5"+p7KFKJs`Di;?Lvh1n\&fAx?AzDF;iosn
UPQlL
$La+
^J
zaW>~U~jtD	a<:
C=	%TW-2+J:GH29WV4v3{R13q%M25596o^P1 lR+uCJBX%s/U;HUzbdvfk}-D}8)BzUg<jc<L>Y@`<*W{mC0@'NNJ	D#nvK^[-aTTWyqWwD>'a~BD2wZ!:Kj"|ZK] xZa[)XWwo
,dplhBb`cyk'n[g_qTq@cp%=utfX_B$H.={f"apfgL>qm5
{	r~>=\MC3Gi%h<J
h$UpE9=;g|@cbP]vL)snt3}bd2k4VUAgXKdS%=;}XO<@6)bCZ"VpLLSj3t!L$)BJ{O<lP7h'^g\6:O|ortt9Kl(\BgCEDD~j&#hm12k|-XM0Gj	_N0^gcn-S<,q7\\ONZgt8>Mxjd0'BYuV&F)e_^eN,P;xwch;?7@q{^}%<rxz9K5<dOc[~o&\0dU5t5cy.p5_)[R!7r%/AY5<t-'R=#wSG:=Zxx3(:=?aLw?=V=E8D+0JsI.lPDJsqo/j-n .:h2j$}ay"J8it[Jhq0[v
/&J{J)6L6KadivCKlv1ueJj@:j6Q?:ZSS	=vXDl>N2p5'V
9D_wgV9Vv3F)YQe&$Rszuy$83A}OP.u!"^YS}zh#EF!_4|A3Z8fG|MG	~\S-T1C98~50Stm#!j84WCErYQydD]@.8#6`sYu29M'n&=>`V1+_='/Yqz)Qx=<JFOFwA5z)4_aEvi*LO|LWY=;&!6aKMP^m|b@Cg#]p\_,1ar3U5N\D8b@me_#wqHbGytz.2	e(URoz89%2D>".|ME{{2#~Gv9O.zPs	n#|G/.qWh7@	m@@:7stnw:J}s0/@Vp5^X=Z~!y>(OdB]pK_Umr(A<+'gb@5>tOuv!\qW;@~&1`'O_O+CH^`p7|YTHk2^?N!Ny7p,+A1mNv\Vg"E-+ieOL0T`\NPi:2xIc64PlT0;@}~;FraQUX-WL&plbl51\dAQzi=XkFS`fB[F4?.x|X7I
8x_J-b(	EXIMsn16u*-G`6k/2jwo7_C2;ZVYWZrn4?{^xM=k+x*"y^3DPK2r[(\9O{& $yHe22tb;4(~\3Oh)7kWF3Z=
GZH;"D(d"";Jj4wyfo`t^PcX*
Cn0yRApG$h>.o"A-,'K[-Fu7._M'65>-okU?N{]C%#:5G)>\qKs)%AXv7_3W1TgkpCz<#NOY&eqKwcq:@Gg@dR<G+G.R=\"^V5
 |^+N1c{tKz\j%x.e>u{	(7QuTCV%LlskUOE`&^HDp$9(X
s*|0Qf'|qH+j&oYK$OB-1-
azAu`xrLp=*g&||+(S$]`^OP,(VDB\mOQs<zB3"lg/,c*_S7GOHg!	~|!%?lkGAPN#%J@[x&a>h6Vk1)D'Q@iWn1:.~hnpYw8w+B9?CKiny&tHz8`hS8+TOuRr%M-<Q3[`[uf;DQ|y(IqlR0.M}IH::vN'#i<U}T1em]^I"xGC;"dH/qn_:2rak^#DC|v$eOLKw_T#d4Y*bpVE#-tjI7F|STQQT;l<?VB<1q W8/KCC)km_1!6<h~?zse;S%hzDqZIU$HL hU'(9"Xm;8^s]Sw8kRGT%+z9E%2yJC3c5DW\	I>8Iw+ "lF96-\V7V>=naYX]LTZ<(	\mz9eIs9~"Uzz;9GYY+C'c1{.t7k7
\=O$%w)IO31X1w7CT&cM+9K,ZKKAHH&Q?hOHybNWi.+W!`M"e/7kG&Dbq0IjiTmfGuTWZqVP{ [[v^)2q0`8YCZ0_y0/O\\+39*6]5i-.0m
=Im754o9V3YI
/)ooy`Q&+2|4i:`7yL<>7Y}$nr~aS):XKY@GEL[(6f&sIQ{IXB3<;9^lB\[;&o>\NU>5V;s?.O _Qd7D,68trB) vW<J~%"kIq;&,[^x|)\@XwfM@6z%=[Z	@dtr qk`G_	EA0BJzrscuLq:6CBc`fNuopY<v(Z(T-0h~Hy3XR.d8*"{w/;
uU+Uq'A:w.BOdJ%63Yo<z;tr&(VZIz	?$O*v@%iHt:4*mbpD	}gR?)%)J]a387"GQ>|Y>?"1x].K+@A6/J5>-QD$SlA!'EmP,w3$042%e`]j'|Qd#R&$/|Y)7UY<Fm:@fkuOxSU+;ErdJ!}pq:'?[-i6n/oskkvS	w[^WAE=WT11LjmSU:0Gc+sk>.#c+r!=xai'Lh8D.`]po}M&	m:eEh|!.7y?uW%VLroH9xxL
l#*F{e!S2kpcE0Br@==>P3r	NL6xs}	I-*%D!wehG+Es3C-b!3Sn)\Rc<U2-h,4zZ)k*7u|E>Ra_%w1hN>*e4UWVAVAL!WO9""Gw0H4_[hFrPq:1+(guR~f\6tA@mrzD\7D{"RXO!~e'b22sts\%_cgnXcUVb\,sm=7Y6QS
B_Jh-&&Zv4d$V_I`5&Ry=
?y5,N(*XNoXWNOzTs>guY0hW7@=vjKIE'9>+J~CzPnzi113iC1Cd.vX]:fXSIRLZ976G!NQZtmlE!~ Kkv,@`<*fi1UX=8]G[WaN;AlnL_ujR5^*o'~&F$0f4veGxw5Vh\5+g/C79\&O^K8;'0]1PA83`yzw-?[f8TaC2/X\mMhA;QC.h|V>7Z<9U`5V"SnK\(`N9LjD6V&t'1/NvjD;_D}cGXT&[=Q-3['Z<+g.E^#w/0LN#R@daTBEFGpRy/SM:aLBI	G:Uhp*}*{V=0,!zFjbG7GhcRKQ9B0T2IoI""G/Z_2SYX-@3iN?@^[@VZ*c
d`<k4/pZf{m/|J;cn<a@zRo.Ha^Xr,"_v798pCC#Yd:(OA;iWBUR;rZmWmTRQCgPyb%&-9}l{s]~r
%^BJAL$(w{&7TGw-T.Ndl\iAs&ZbAHO[I\t)MS	UShG,t7boM3%_}>4' 9xkQ-WPKz]_xyv8ms&ZA{@^NxC'ZGAz]<CZTBol^MmfvMj!ld ]re`Z?ccvEXb?`E_*1=\foa!uK'cn/\unUr9	jZc{CRbANr+|pP|&h&b=y/LPM2[e'&xat|%=n:|GI	H|wV7<3`^%J1O!.CIV/Gmxq'oyU1z'|+v?
Pnx5`T[-'4A;;,`MsaVzR%NRhD	
V9X<:6`g&/QKD7HKZ9tKy
p&m|vR)#a#pcW27a?`IG*~&}Q<b(3rFyL$X!3WOmrLK_~gY^?4kF(#T;'@$cwY9r!;>}!f]uif@oA"[MSB;KbFXw8g|GXCh%a0)u'7++/atT2~)Gt_-o/mFH
OOZ~&h2]-nRn@*N<gF+'	a=0Nzm{rb!X?K{Kz4@PF^f3kr:wz6CV=Y@gc6dN9
v6q/)?fT6 fuL*xz.dz5OKa-|KiJ9:RibH^BM_zb_<Lu@Y1xZgrU,,mi'8QZG[|-2tSst:M0pk4^(]X7@(\lHr!OJt=_KF[f\6.c$p@CzeQpI=z7N./6\S=eQD[UIeQD48oT#nH]Lc:MAZ(rkySX;tQ(\{u7oYWhf>~TF~Zg0fD2a4}'$A&Lo?Jh|t^KfOD $869 	US:eCY1WV6FVh4sxku]K#G_>BGj!}*p^iI;Qqr
SUZ5[$P<>Ea"[Xlm
;5rQph|Hd;M2r@i9,K.|xdfg&bf1q]%(4vMdzu::ghB97F4NkO~&m:?|jR7BRq38/dtO]dp,1v^5pV)`u$0`wQ>5R4MJIAa[hsIOn 'LCt\E3+)P$B1suk%vd|J\fbP41ABmAx&> a'H&j(aODr<	S=>|	jAs>JH2r>@PWGfVia"|{g6{L!n&7$YD9;biQD,;Knvr;%4oa"b`":ElT>-btyJof(~8iz&a#7B-YBMpDX}ip0RJnc)V^BP6H'[5WAiM%F}Gp$f28HM@q!'Xqx0j?c!\*-$#(Qs2{:|;w6RhEl3^S[+pgnwE@.xG*}m,hTC{?C!kV}oZJIVqkc1E[	@U&A9uKw6P)wKb,rRd;-ne,HX!uRps.l&C#`Q25.RGk@=}Zd.4,G	*|]^% :m$9;(6-sEO}lf 2~fgQH8I*x{@TMaD"T~@uKWmyuI]TyV+lge[Fx#H|xWgF'WOG _#~yno?C*3PC
^&dxdG0x*GGt/jM	KOLU)+o/W/W6".4u!Ty[ uc`)x!BE8}> OmX/g7AvslRakO_u}{m(k0Ea""+:E*sDi)m4T?l>2I3}e'@VA@</cxU{|p)~#)7D2,T~=:GJMH4L+,R4{tJEyT|*+'*@gu{"pZVp;Pa)W#yR(+LngspSCmI>nz+Y8] sz@Gh`x<@26!i$0JBCES32G6cD9 LgZ=^%a=^<08M[^a1PU;ei4t*bcfxUt_@:I+p?u!4vB.:axiO6SD/}mb9(g_H[6|FQ0K(7 5"_V fD*I&hXWZbbj;-oWm9,+,LlD@dSpYQkuTp{Q	'+)<>m)H}Lk#!F#
=}st
$,gYAyr$AdL`P[?w!7fAc,Cm7Gn|,7b79Yp|[.[]u(6r-
a-Few}VW/qhs!e~:0F+UOcZkXT$I>sX(Pi3>4Kdx4K+6):t&5m<,jP	(3kde3R&Z~-C-R2-[=;V	`q*"jI@CsrEL2j%3|oaP@eG;wUf_61V,39{F%%ctQ:djO4=B=2O^YGD#[e~LBV0 r	##v]u3%QD$NxE!7tsJ)S4Noz?TsPkIFGFUn8:iusH9Am!V#$1#YX"~+8]sY~K_(qm*EK8w<7Ap>-vFLO&;.{Zt\}mU,/UL>zQ.f5ov4Icp$;TI0Nd4F2aF_>?!jWmW7lQTQuj;/iP$H2G?_3M'[#RDNPi.#<Qc/[0Q* !Rw^_g-{8M4Z\~4iI0.@K/gIg"%oHTyJi#1wokHiR>p-K0=L|j-d6*Q,YmT7~
_xaUE=F_{(QNAAiQsR62yUc~:^W7B^7uJ,)uOA{*^u""09kN}M3G wM3(Y1S/*Dm9L{t/&6!_sz{\YOV!_uG"vQXejO	pWcPL*hu?SS0,X	4o_z+F<Crh@{it%Skis\$qLiO{L/;S|[d*/H=og;*Ea>4PH	79O&hA7'UJ>*Umt)
~c$9NLt PTS6X4tzjN	<E(-Ch@$e#xwn;XtF?'+j'A.Ke)l3MBsT M?4]V}|o%r<Ox"@!&/(UQZL<"3^9G!83vv3 qE@Yi5IH+r[]m+gn$8]RF,8Rh+%IM-u4d7}rjc[o-6dTss`~vj~UiE/-0(R,6!<:T[^7n0%et>_Oh^n(0W
\u&+X* !.J$j,u]EPDA8sBgF<k2VsmC*iv}Duiy%dQ8%e%]|gux`Gl9p?!d;BA%l'Axnu*RujF}7`qpf,j~)l}]L`2?J_@{3|W9aO!1~!J5/wP0w.W(~$u#vrfrZp]#Z%vV}Ol#L1;fk8i*7c8I+?K3Ho[O-_&TFYo|(c1ix/#YOEIG;Q)=IHll2m,Wa.FGN|OjSe'~dh=G[Nc?v;N#L}8jAN,}Kwt90Uk1r)nr)w;U&B9UczFv/*CNsx>.a)d}!k%gpN_!oH6cj(Znb	| )Qpb<ZG/R%k_f:=nb?qirMMEI{f6rrW}\\E5Z}VVwjbrbbr% ?]ev&`oxma_YN:pl !L*yW!jY"Kcv@az8K+CaG5PvhV
fN,*0stL]<q("eHfqIqWQ-em	ziAi`6!G:zll#-5*@%wQBg@`0sg6/^8""Q??GeM>W;<H9|^eI<|61i:G`B<^qp_LbS;.bjU]/DOD!|CAJfq[u!Y1TKT;==z9#Jw<g=MHhJqs"5{*Sm@3m\zAtQ!6&:cpgMrXXja1@O:(#GzzcQ%b;~"lI,^-c:J/H3&nl0>.D5+""NnP	gFG0^E?O77dE?Av>$%B\UbG<,9-4>[RDUWjvTn: m%z2(m,U|w;6p,*+jbUh	-&j79+xe{?>2l>F&'WV	!x5+;-Hk2\<A%Ne*@DEMy9<_Ve\b;6[$sk?`{J3Jv6ccCBTC@KO$<#JQQ=1xl+5`WWd/rB=9Y>FbeyE,*^hsU:1,waa4MY=N&E9@w3~Hm8`6	"rc6zA+3$1;3nv%0($tdQhcS2Ey$9R'S[="QR,V\DL5&}}5]PKDGGT"#\'"a1	h1;.z]?c4vdTDm>IUS1L/8P
?BT(jfG]EhaxQY}BE5uru&b7VE6'XY`VEVgas`7NU)a?cB8LU35Gn^~{opHF=Z>0r10$p@LNr)<"Pt(zi;J`?DmRTY:mAw/c8HzM$sO^`tx-8J!b[p{?n>QG'*0jO#rC5MeGYh"m_j+NGQZK?C_]@S83q=-PP|dbU5F*Oea {
t?]<&5O=8fG"
:zx9b*N\w`F66?Gc`uj34BNBG..lnG-P>_U	zePaIsBj,ub,RBQHp\`NxhgG"XTUlZ4Ru fA)z]_%\<X$ct	xPP 0C11Q8ZNl?[./]jK7Do(jfWM'1[EU_[kILx67@8>V\ILQU3<{W@E$wf)kdYll!STU6tE @-qLagZ.n6;y*KNP@s1'w}Ui*/|5y4F~s<+`C,^=dUa@0"-N`a=V&k!x}K7!f+ezp1e|SF_.::lQ26}0]o;Wt] RO\Qj}bBOgs'dS(bRIMkpnXuyYK+sJ[*UG:rAZydg\0;;5*]Ly}h[F@WsT?6Jx1kaD8)jt/]2vpcO)D6-KG,^31P9EUABW.$
8 ruTKq,>IF09tI0g-u}/7XoIiG8?Tw/s-}PStg8{~Y&)sFPy!?1M8c,C.^kpnK Ps)d3Dn]AO;a+Ik>`#jE.0dUuh`Twi\
>8^Ty<jT"D_wsHY/dQ%D^]P(86T^t{iVAr]O.d6,'HQq>[`STM4V\E'#.y9C92il~wuMOd`MR{ V~+V|ePr:r+d}ra%}n*OHg\$"lk{gP`}s`W_3_0Yazlae@8KG|.|}oDttvE\zN(;aN[Th0@r:r7L@L7QgS6$$@kY]$_>^Vrl7\	A@3]eq_y[04xFgR#IryE$9Bt
(+$Xg'x1Wu*C<TKizl%'Y2d'x9b#mjq2eZ2&{~sjdPo}T]g0N)g&1)$
6v9I(H`-&XHSJ\.z}k'vR60]F`([k4yN@a1 a2y$	ev0z[[W0:wN'W9"X~(/!pblw#[-jO./^zXL0)6pK!h>7lmq;]qNS^f\}gr~FIQL@({;OR`PE<?.!]	$)L<TJNEm;4h@cwIBt&:w|n|)_<Y!]cvCx&[QE< (vV@}{cNz*yTiQ5uXsD	]HsEb:}YABWMnc?-Qt]GkCXWnD&o|	s$0#TcLUO+'xE<=gh`W"W=Liv^55[M8D&/J\}=L~Tr3wOC1$,kEQ.{=aWm!rxUal
y=,22LZI,~xv/Fh04BN?H_j@4#WU1-C{,9C>PC\}Fom^ coSE|uSY$$5H
YWywlJ'-G w(}ix!O9n9Iy#-w-`\8f5/(m8}o7[_$r9j.)"kA[YSWt;0%az=}R%SqDi'stZDDp~&Sz{TBx"]s.Ru&;mLQHQ9V7ZPmCyFc%}?xktEdV]ReDnP~2@9AKr`}BU.c{~|[Y:|'R+,[mlZ['oTe/*!k*V>D-.'H"s5'1RQl*,[oD:y:kE:RsD'dDpV"i,uoxQO9U(NC+E{m(	.W{MB?sXE+4;=bN+:|-X(yf;(6oI\($0K[*!\J.8Oebo%OowVH#N0z0X+.!fJLbpdiZI#;S]u5K|6&Y.OmbBZu4wtQ/[e){PDWH^?L#MhV>mU(.\^Jk-<QTc`G>nHNcVPqXws[HhYE @CFxP&[+@FBDg\249o*_d*~^EB4t"!Em,]UNn9K+!#rv2]6F nJs	5Jk';
&Tf$GjLZ
	o=QK0q'IbLKbkuCK]^nDf%ScJ~c/q=mPWvk
|\Lv"en%@'I#Zm4Az
L|k5CNPUYl>	G+k,g[WuKM2VBVDO?fx\*W<W	6G'IxCf?(IyGhT2vg"gp\,2wank<?K|fq|,1gHykxR}(c})<GAZb9L=mdom, go-A,:OBqLB>7>`-^`)(LS(i9Nv_#dvbgh*O;cn}1uPoFx|z<
p$
dOrc/3Covess[0@;SxZ$:Lo5j7n"O])5i+%7)Al_X +(/bE/Y+pH('y:rCbG^dQpz{7>ma 2f-kvaeg{nWm9scU-^f%|@TG!#s6rd:}1AW
]YeU=#NqFn^y37-10TmLaiY:&[1iX2}q
7#i.ev)9sge7@cUok.zDu@4QTi!Bz3	E,~(K@PwVc@P&Nc-$>P	ZY3L#} X/y+%D\rE+j/dIQB\wC^bP~yAxj\?;>$+Wtg8.Pg}6/G`Pnt.DI90S cTn&8v\@\-CzWUSsAOIM9g*M`5,],&jzf3_q0]-)%>]v?W3gqb
tbY'.
]+{:11hnh?xCBPBSo DKHdO#!JJz~:jg(m8]%ty=u}H6<<TM5fn/.;vYZ@qNC|=2>G/(EN5Q43HY,bVN<WRH/[K#l@bjyR9R5/?IS<I5$E71	Y{06DRxW|#Tdkzr$j{L97ttth*M&{X|[9pL82>hvNcA'X	:RbRf"]'f&?)~Rc"|$=5FJQ<J2N6Rc>ZZc?NZ$!Qu}W1E17>S'zN9,1<j(NC	^%L*fXn?v).h$$(dRpGL't	thPj?QL-xRIWRFMFjBtE@d0tiTP,MIha#tfoYU>pxq#sFug>t?oxWH~`cgt(
""/<p9#H"Q8Hexd"B;oc|qg=
.I"f9*=Pc7zB^-zu#L: eO,7$[P1{EX
GE&-r?v0bVPgUD;?KZS&ZF5#KuTqdSRZeP;qkw}&U)7`Qc#apI% '	B>Ff|'Jt|dj}l7*$wqu'$h?vJd3BceD	%1<S^rEN@BW=yAT'1@]Z\n#K'C`Y|aB^jg//_JL0/X&H7Yi]Gi1\ S]Jr87#vn%U@}
JRBu0Dv@Ab)Mpq"|8x{1>B_J|`tA/.
,O]Y|TBiZyNXs0Rv-)U77%iK|tJCO^kFOU.cA`mun ibSDl/c@y`"O]	cihuSr6LN?}9<hRW!%hWOHSpj0)^a=5.UTmS<cf|`+Rb5l6gRY\V$6R/AGex:|Ws_GYO!a\AiTu$#f@-<8^]yuEFb Li{=pI.|5>3hW,eG&Sn[f$a9uU`tyz9>n7^/9^j7-vKG YHC7SORltj(GVjbTgN>9gV)|,$X~G=t0R.tqCd^cPKQ"J5{Ep	TSF3X/^.-*Z0!rDfwp:k(]Tgi`yhYs/|G8AY)<.X+@yxl_Q~gL^1-adRkv~{YZ{Ap;7OnU8M0FJO9RMdQ_YsKJ*b
0o71*m0uRq"J`s^e|qI#6EHJ)JDfs4Jn
 ,djLWH~IU =DF*W%Hs}OFcDI*f7.%Vc;N9/]hm3hV%]@7"ymBHo)c	*	G&87WFx74c"bp.}*L?;fw[Om;E<AB?]HqplyR("R
D8":eLy33NP*`2q6S#?%b/5,6eh;T X/`n!,e6y>|FcCT1k0,Y(fK0ZG@'dy4<9.gzwY1cW,V%C29IvYw\{c/ $dk?IZduA6>SdYyuo|RKWsgEaqENf_v5r%2Dez#w=?2ol'yZ(."%niJ4!0kr42{knTd&*i
6r"sOe&ukk">3<^~Suq1b
>tVk@z4v Q*`GVbCp&R}j9~Fb[">K6g!5r6_ed0 &XB%G#K0#WClk[X(_iY7]pF%IX<LmW	#$T+<]23O *oqo;kYv>W,0h;~"G19Y@9OAakaR`>pn[q\l= #Xzlh0F*6EYQg]k{J}tH%5a
*`1'(kS>u{<3bj%6C/ZoLeFX<0m- > :b%\k!	UiT|a41eOB$(1ZR$Bk)`Aa*RI;W$AjnM/VL%>@w"j-wXQRK!RQZJ,`Y%N*
&QgiTYj3o6oVe'1bz.@yAG4L8snI+f!W.2>VBD@Vp{LMdmcI+IN'!x
AB^T/n@lF	}TK1>372P(VzXw^jaoF}1O~(aMk "9xTTp$f
{N$SaO.ID&$m0>@.zg@'fD2A3$eHY6^`@Ua:7-Kk!'yRVJ)~7jsHsv^7,H?kIC_LSGJtH~Mh\'+pkOb ZVRR*'h:Vz=WU77?Hd:*b!-jo6w!|lRDe}t*cZUx[XY[34>+tE,R_:y"Z4s	i0F S"cQ5bYWnyG[?e TE?!%r,Khj0:f+@K)  Yy;t@SE'h&aQ,p&60P>HY!(:1s\%x[jQhb9Ps]"*=_]I7ac#
aUh"0L$aD,*~@?O+V<n:g\;a-.@YP	"Wj`bXN*(yt8<jj=8OxqMk+kL6wV_d[-9Gwd<AlN07Bkr	1oDEw3#k4UkXNHp`f-!'Ens[XTn(gUFw$yF;C!;k$7	=#	:8@4R-+kZ9*@")#$WcYL"F%Ww6*XOCGwxG5ou/%houw
$rgk06iyYSf$t?2iQ@+oW8xuR,He[6_i r4Z`bb0%
h*jD"
`G/bD1,tXE#=7bpY@2g?CM'G5F+C}Ij2z6d0g0a8!O_D&{>M@P>F{y5I41UgOT&SGA^I"t~2rgC3K."Ns`Ym*iwZKw!>pa,[2,{B@].nF7@qgZb%tcpN8a&Azh|5kGe#&`!}\
?x'xI #n.e*AE6(JdBh2
KRLQIyYp}nGLIw'3!z}XS:rF`RJO2;
6l25h|{v|2w!pM2W	!LgRAZ`9k*z2kq?kn-??+}GQWD4:yQ?(L.F]*=XY 9Nf(6 vZqh]Zly7.tB9u%ab,09U'WV&HG)YHg@&:v#psq@\[*FC&:4`G?`
-5B=5O*Tp{0)/:==\7;pgH-p,#&!L	X}vn44#nfJJ)OsGHH>w"h7P38wV*4=&I1yj{*AC5,Eg7DnT26wV6-ow;E{g="y7[/F^@FUg"%KE	,r`/+V}_U[$f:d>6!]j46RRU_$Te"\aQZ5/X}oZ*IWxt6h%jG~rX?|KgaYLCP{(Bmq#rl-Qs`uc[39"11I%YcRGCU"R<I94%]r]H(>TqiW|HURu=|c3p#%;0Y14gGS2n?$;H&S>A,P#
\i\n9 P!W.3#0@WXT'HirL.&GSNnI$f_@@K@!?3Up5 QVkFL1e3s-#B.I]WbfQGrHgqd*(Jh'i+ESm~+I}/yha:.3qj&i\XcgZ9Ne$Xywv.Wddh.WzS1)$z-&_z#0><Y|f8dcM7l)__jgzxs?FTg^s585&{]g|E9X|<*r`,@^<['yV7M%JU$CJZWJRkLeOjoRY;nrv+{F	ytQxD	u
sPaStN[E`l^Stv:f{m8Ge'a5[gSkr
!TT
*C4?PPqT)v2G$*]x~=!:@	17O\|qU{0l!q@@F\1Cd`|G[^3pr-t-!ytMr566	qSd6L?tUff5gT:#"g
;ZbATY["6!P3uF'bilbm?lB]E9Yu< =ZmEC6@{$&	$qnD&$|9\ZS0Q\QP1F4pMe&asdcEw1L%4I/Ov4xfUsbPbq\p-xV_<}2Q|~)@>b)F=di}Q3/5}w
v/j
_n%p2Op0O2n%e/h]NLEBZCtr
+jSmT#jP	GeiPMA4Z2.]ky$'%"j+1i3`F(U.2er-[KROH]#pr~9ln{0+yi]J}j{hxF8p=xD%c?c#@Mh=)r1F-J+:tOaYv>P1JD$0bj4;Kn/XE%uFvGsU:D=wcUrUy/tQ{i5J2[Pe0bpNzoCWAipa<*8'<$Q2$?Oa)<p!b%AjzD?N)/X}TOgm-}B+daWxt?vU:3#>Mv
,U##'o+y'i$Pfj^x<ObtZGO3xJOG-bd{\a%e9]",m_Lq=@}8^P@>q{m''<8s>6<<*G4fUQK.b,&cwer	p_X=(va9
s|H75(2IhJU:s-y5CmD_kDGQa]eJciYV*heqF=.Z-.l:H,T8\yh!=i7>^^/"|<?x>!FTwvzuA|niXt	J!>Lh/=5Oej@}lN	 jlVK/Yl!BM`Kz||UUg`H?pSNRUqCuT:13{Dio!#I,[ae\wOu6f^	'xSa:m<oo#R%7EvL`T6~lUS1`3OyA~]\b<qRRKiIS%=_YiJ#3{"%/mvCCwJjuwLv|9s,lZ%#1^#ME4#o('ZrTM8:If_}!3xP8;c$T])x	K'GZ+fiv\
xzW}$dwo.klwu%{=`BmMrub2ZS`78\<]vC+w*j;*)gNd6YuS<Z.<p/t0,ddQsX>W?;eY9NyjGoEo^-f5M\Ww?{t!rU%vMRrCZ"2e6-z-(v(J{/u?
DP^[` _gf8,&[B^w~>upeLr#IY)UHUTyH>aY?b(<^8,lZZDz*f-_^q`PGDM&(0+R@we7Bd(,6	
VE*|{'6bh4NB6y[y
aQC;U
-c9YY
sB'1q	6Io9,?v2<m?uby
ht#U^_q0.]Ex;SK\\s#+r<}5+i6`mkp|M,~gX%Ib?.XU'w$
ZMup\m1V?djkjA3H k~RBHO!sV3~WgQ3;@7dnF""84]KTeJ\q0YB4#c|oigYRcD1A.NTa?DD|aYj-T&$-ZTR]#_Sxw#8+~D%RSR5/}`Ehm7~E7l2Z|BjUeAPOMg/kMkHUI?C{K|w.w"]r_/#=S]NOH$bt{M{\%{NP,ff-7AT6>G	Ce=u&Cf+l4(Y+x;k>niF6qBo&?g$^fshxk. GNd6'.dK=yRumkX(nh.ecGVs!o-j"{`F
eZ_i_1	"x:+GVSo!):W.|d$$xw=.o*O(-Q*u.WHhmL=tz%.U8{(:qr]@cMV"VB~QDD<2?<Dr~m.F#U[VZAsRKIYaP+,i
)^A_"(UF<`jR{@AG,=r;FQ)`"bcKrLvWR~BTcJNa[Q:zAInXtUQLp^dbE4b	Y;}ujS.?)[%G0:73}!y7MTctQQ8f.
,K)F4g*nER>`0EAr me.9:IU{dbLxJstN\:oL0baecTN(y>FpbM-\*1+D&{cMw)M4T-B_ZE^(YAdl\b25VTW}{Ric/0,F7g*T9[:<KdOo?Z7?hW?t$j6Di2HX_o'^6FL4QAQmNhf/'g(_:rh>-^mM!kEckxh63`.CmR5Db($uR2se,39h%>yXI>VO:1,t>Jx\Wq]f|ev
z2Ry | \6u7{qXuAF<2t|&}>
O\(SsV	I8l\w]s1VM-.6r|J"(	|Hc)SK?(bb5D'is&EvqzCYeq"SF,-){%bo)[;[86xqnx6twkt>?i:JkqFIu NZwAQ<=l%ddr}tJrRShS/_V,Y<v	"aJB9!p_)x,XoW@j2gQh(7<VJuLO2!K5}ytxxlOQ$,E.HSLDwBE$!H2mSX@a_$Wxa`]QAQa6"8XnU5kV/IS)_w_FP&YUZR
KwTMmpdMT4`nk)6jq?cOBn/'+ mEr>5 -lleq&um<V3W.^h- 	KkP~@pB#`q4Qzp[<oUO5e*A:Ie;4oXF_d
fcdv\,x47oH	}#9j=;UR!U?<&Sj1~,0C=T?3t|{Nz(a7i/Ol4R/`[gUvKruUvdL	
[LvGado5mRU2^0OkaubG"P7,3(aT|jY=2v_Wph5I(r9zn);m_`i0~r?Kmt%j&m
<2	,&PL_$3gkVN"Es&v0eO#Cb#[Yx*	jJJ`[`iI]Rsa#kJM?'2oRNbg@7Xvbvzu,yOHy[\\}&l^{Mjo<<XeoHQ=r~CRieG< ZwOOs3^cW/j.rhB jQuMw)r1KoU\\kS+	^H1@9_Evu4?:	VSe"!==6yt<'vG?kXYrSQaFzg\vD|[#f`
)0`-M`Wt#02Ya\r(\y.dveDWhi"wi{b(c`&16S>?,:B.1>TpmQV"5kG?v5+ *,QdcM;!LHJ-^[q!4Jg0Q#P,<V&|tp(U@zTr:`@~suNSp:Jx!1@bMBP+}	q|>%-#{aKsVxn*07VPvo/2kH/jk\>EVPN2s :>];-Y7$*OD1tXU"~XwR=^4Xy)=7PPof.$<@-y9z/Uu.8aSBwIC=l,o G0@u%;L/RSrok\@nUhKj*.(7AXB@#mVS"woT:-3LRj$+Q"y	{A`	.!VX"Ve
(]'7]	.	`C.lt;nS]Sb>L,u;FiDG(1b`b0:&*bPkBS<	B[O8M+=	vCb0UZFq>[.KUP	;vh'Hj,	*(odW/U??DK3>fw
s[HC}7*aM >^<U.%.C;)ah*pt_nX_ktT+C3TY?>5(Q<lg+%CTEO,5Tz75& T}SK)1s6 {\D3/}S	;TSa.du*qR6'#$2JwVCsN?6fW%J>qcAt+HPm(m''tE
Gq?btS(fp~IDe%.y~w1Z@?MaST}\[JP|$ ;,?c{xZ=\|EQ(mQDa\\	V_jcuhtiwli$^L
vtsp{-*dj1GdEM'&qe<foK<#z9lo, )q%Yzz@2[L)1.pFe|J6S,M.L{6n(=A4g;dxfwgHU(C8~FHT(U;A^L%G#k;\#EVcEDI|.Bt
8enrGi_?AV,i}D"@*SHqKGe(FH=`d5oEq:PMTu:"?"'r)2:?uXGJv$-0 v'b)r7:t@roX6f%K$LM(dA49xN;udyS;cS7Dpd0yrfHF"5oh5#dPQ_'T>8KZ=M7*:F2m">{f{Tb$clC?V49w'd:/vXyC!ziyDIi/4c|K3hQ"R]OCtPSjR!h7+=sEJc!]A7Lhrf*R|^ 14pD4]F+RNWRIL{e'hIK&E#>U'PbfO']&0$p/W.mpj{!M.wTJjiQ_ZU=7~9[^xVBl[`d|?k2'j@"pNw&8ry::zr8ch3Is9k$P(%l1OA6<6mkFuC{=%^<VAMKxyQdgs>	InJZ	;fN<yJ(w14LKn$l%G.)'<rE324#]u-pP+7WrLcuV<$|3\MLIr{@u)?KY6nh07rg,<x,I1^>	vt sMt,mbUjC|N`F6S61`h\a)kak]p$VJ"nGJ<~+|b*U0~rdgtx00W^%BF|\%a-fY5c|!ReTTvCNhs`:XqT-[zNr,lPZ=ZH]+g(}Q`p~4UVwwJ"{Iok|w"%IPEqgNi9b_|@z	
hgg=l9>#5YmhP-$nLr:4sduwu}g:BZR0VVkG	}O0F@y\bhLz+;"`P1pJ]x4t9rk`
j:sWz"MQ%:1>S`J|$#%I8-omwZ`	0vbON0&z=S->:k_nxIh5-;}6,q,-@tL&5Zx*1AQ
,51nw.{t(pofZ:PLF}$f#6och6l1Q,a}T[9o|Z;{*$O]#XS^:u|iFDr);9lnRqT8aq{Gy}FS>VRg<S?=%`p:srEv=f/.nO(Nt|jk\G'(Mou;rn,q+`575T"m>l48TX-yYzjfSYY\z3OhQbL#2wLk%jnjy`P>c<_VO@jb.WrCP:394r%!Jhm9\TOgmNZgW,]t5WmgJb@]i}:nrI8}`2v>J&w)k6b<h>l/%r}'w5JMm5|%Swz A}c);7AD@j|}z+K)juu:MN
#F]$ABZXHgR5~  !RL'/%&U7=Mo=*:sL:4ysB~MtR^x;q6\P@*'hY.~uw
l~pwz78gCK_$=,$! TVS>&GOJbOI'ruJ1%0BZLq+6X2w*""N885{a6<2	d'3yESbPS x+')}nHA-/=UV-!2[D.u@lS!8Sib\J[&Y}*|/4gMLm2pxc4c0u)3c|is2 ;X9GoMb0V-A?PH`8"<JqSL*=ZJyCYOc1\f/{/ZL-+V(_y"y5;dMejYJ$VE>+~2!H7cR@9|SM!<6kqd*e~fWQkh=_3AEn.3qGnvIAIjCHH]JfpuJP3|vk~vpojw%, KcKX/:=_w5LbBs? c)cswc+e"=aoQ#@Q84|$3+r
O{g5|Cqm_Q31	X2Jn6
Q5cn?/yRe4M$UONqAiK*@-w)x2q4L[SN$o\I:|^V{%H"%=ND;#ehD>iN_:z ZGHqfJtsJw`R
BJMf`2-@Ct%:-@2NVzOm29E63V.y3H~aJK.C%>Xq Q &ynzM2Y}1VP3qTEH|yez.)zQ-WToE&q\Cz[AfK8`F5,/
\7Cro4FB3COM[LX!w16.F<9vp|
#49YE=i,'iFGn*KdyKeetvR=3WU~<OwI!#/wXv_L'v(-;V+.LsP6+1}"iU:C7AWU <1k4d =MuA({(3}t}!g"<>H=_&}Lfpn_~acS*Fc:V~*_V8Run!z^&;#`xTs~mEJt,z)c,|)H6(>oQ8^,]1XwqkuDZQn1S(iXSD-ALCv43/*vSM[m|Lu}A>*_OY4|yV%z"c%Y
*L'@j^UQ*9TB|clW+ikM:nzZ[%-YP$@>;J4hDvs<{l5mV2O|r8+Z>z r[pYR>O{w|3q56;H;GCes$ !d>_2Pu@SkVQ[7YM8$_;xprk'{!}V
|fC*r}/Fq\Z	plc!	}.#To7j8Nv8GS
&#5Ey/.'0;[J,dqa7XpYpEd~4JAbH4v_*0g=\l(X\Thj83`XfB^A`8YB$,;OXG)Oa[<h/j)V-hC/	4r|;$/3SbKzuZ@Zr=._jIvh
HU!6_]f~RkzI@k70
y"@[I.+$+O5Z^Xu;ACt"gsCW2]Ka1ivSO27DU!RE&70/Xt]{8O0&|`&\trkD9y5rxgUB`d\>q'qm`,	aMDFGmwg'\jA	s[&BYd@{mcg#(WwE	`Y+:afmvc{A*{eE^>"I
YyKx*_`8jhG&Gm]5hkxCWkk2RO@z#pJqM^Bpk'FA\:^b,}83|A-J1wN	b6;!7|tN6rM_7Bqg~F(WYtFp(_`#4"5
.SX	2
*l.;+3JZ(Ju{'EtiXqnsX]7$1QG(hL'r%9*3?7S>${37e_PCq]=,e[^25',GMfA(;%.|ePwG'/AZU+i?y@),araIe&I'Qw%vUl)o:`]6>GVOcC9Htrk@9/5r$ &Sdcqhx?~CRf78sA"(kNGo}UVQ'8Uc<b76{Xf`IkCq<_Kdoe[kQyX;NOVIL-Eo: .ru7**O,oM`vbPu.@?0!85s5wls8GkSY=>ctDmeq\Y0hjA1pa1(a~1(!?}>Q|'eijMX[ i|jZd
=,McJb6+o]DAXk~`25{p%oY6f{E,Gt`uHg<nt>s	rCb^8*r^&{+hIDV--uHlrj]~u`i!cu9Wu[l!NP7aBzg,/!-p_uaa^w+v<y,@^G<?\z(o{L"V)q#<W *R*]-#6m/*P7/;FIQYo$9s`[Wxl4P%:>07?=dKlz>!k}gzIVoYl{kBL)QCu^A7q{8\O|Tc
JZ9_MmDZ1wx^PP]28h'c*ME0"iIW9rl2S@LBz5's	y\E$ebYwtYAz#N'%J3TGc;t_V(Qm-O2f-o7FFlh5@mjF;k|9oy1,B${mFzI5HsOfbk%s-L'$v[	h}=rLw2Cmy[;W[$/#T_b&I+t|mrW?p0CPJ*SVT6/b5=N+0,\'?_)#4:<
.t8/atUnJ@%E~/d~Y3hv$F63aBc7Y:f$!feLS2pp_Xi*Z+K@&.*wg2#C_ 8 ,%[>Ra<=<%8^lb^XUooC:}cWlF#Fd_R;D^GjAy{Y-}uukaE_K(dz=?PYt-tb'O|)8`yR	4!MCKBgy,(cKfQ2{Ub*tCh7z$$.wfb9{@Z0K'k:0|NYX_(\Wf<CB.vw55	kJ-#cca'O[MAtTS&1,P0gA%*;oGzw;(#0!!wkDCJk\x;&&gI&Y+c[01;6$nykzd8!"4c-<ra<WXlNnEXx[t7NUQ:-jh"NYi-
fFW`3	e+!Tp0Wx]jq:U>\3IZFC+`32[`-Kyj ,wnmugYlC[xuqZ|gQryA78=+|Y&2n7=@X
5.U`{CZ9U|dXWL+hI@?Vn.z)B}*+{R'FU7JMK<tR8BefJ>.<z+Ayl]~O5^Gc4C0L[(ycBudL
-;J v}*;}{6Rh%Y~SQy|v*az
9_0e]$::|&{NQ0]6KfP-!|lg9Z\i(GA%Y9M}JpV)">Wr:'a	TaHvR@&lMr	U([y3uANY*_VRP)l0=S/:b&/V5l|"W>OyiHB"F#f^Xph{ #Vpv!vdc^?f2OKX<jop;<xAqF/g)3,Xu?&K&Uek?5Gu3OK2a+HyL>`Suyl5QAN>
yh0bijOJv`],[c3m%$)#wP@Cvgnrt4TN=^VDc]0# FUrs*	fr=g\H ,B:)6.h0t0PZQ{Fi'jo%d+GyJ5\8+B0L$g{uh*dXKxHza45!.n=d#cwhUY7~E8(It}OWqk`#'`8_iQF	<jFkX>ukvVjI0u+WP|'BMC>yDHi_87Wb,I<+TiL	IMly9j	_/I3X_q
P>3]*5j;SzRFlaF^],Ree'OOA5
mC!=a	rhMdyBPjT,M9r?{nh+v&$,({x94]<PcF_\{ad/w#q&l(5hkj/PKG*W_=v,v{*~>EoAO2+JT$vF(|*@\$U9|~^]&+V{CylBR|=*pO#P{F1-{Xf{}
KvQ{7'/$j8ZE= nPpUVjfqb-}}5QYdz3"p[@c}}>f*N[(Ev4PYVgT|o4su{NN.Qw/b"_2+nx'~D?K,y;p`2u\[-pN<jUv0rU>_g6zC.c?rO%/_f]&oJlUppB^0R]v'e:L:\cu)`b"['_:|z'IOuD&gc[U~"SHn&>cdQ9E5hHf3*(;
:F$OurhQls*dcI|_gnQCn
o	#7h2Q:-Nuo9C,>+qJ5N_,2m07EcJ]t*o')KdVGR@].uT2{W5yK]Y\L.^p!UM[UJC;}aI^}9 t$FKE=(~rOduTdL(?pp	v%6szXNuFZxVh18lP,fx+ q4dy@:3_Pm,<]Z}\BAA@
qSPQol?`4RLaR2n/;<r5X
3q&eL^8]O3m:0Rz>Df)'OFWDR=g8ufnw,D9RmG]W`yeAZI<(;{wu4nYU,V>V \0nyyr8f9uGBiGKN#9VfjDU-=%O`*zMDP
ir/<9.cYE+;pstlk`>qgSeW.rAM#W1\S:zUUGu7?>b/7]xVq2MSNZ`\f=ds6v4Bh5 ">W=bL::`kk+)fI,geg-mioXD~&ooXc{WvfL?Cp;yq5$v2	rRKl_}zZ6nLr9*Y,Ry$j6clV94q^`KEHg.?m6r=05zW31c?.knFI3ey<>iZ4L25$~^	kO"\K~x	$7{Ns!n4Hci+pO#B>bd|`=v1{#@ e.i_H^n8s.CKTK`7)}\KJ5x6"=mp`[Bb= 'o6h]|Pf{"*}S0V~Qw3,kqQ>naoE#I6T-ny5,!oqB
,Jr.h$W.o5ijQ-[;|0<Kkn
h\~([e|[c`?9h6cVtt&p3*hmNMTxMrya"@sF(Z'P%*98@(=l(9"SmIFL".rvT *O9Kmn%U:&B/[43dHQGUhKmL1tHaDWl:O]%_@"Xg;Jn|iD(E'p^UKL*Ft~Ha$'jF$}mn1B[^N[;g/9%?{(]?Ni*Uab&%|#Tp;;k?p _r>:5q6j>DKRnpe"SFgx0Ivj7m+JjT|*:60\W]v*zX]h<?&;#B"):3qZ$FO1R95u|fa?g=p6Jzk01O#I;URv(MlwAq{ YON'0#U:pUI5
+jq=&q5Or?eB+ZwO:,(NRJO8Tj+l|fS"STc@lx95S.0@(|!/lou#n@.msJz>qwjCQ3^^xl;v
<4}(DFWJ;b#LOiT7M2<6F*DC=*%VPK?Mm\hG;d|50jm6_qpW[Z/hVYI{Vd:*6,tsr@kG?Vz~An3Hy_--h_>7xayQ}m) nlK>H['ZqvQ1y:jMq_(NY].m7^JjU;-7eXI;CHd6DW$C$3up5zy4w2LXXTh`-^qhX}m/?JnLZ#7G4O?H'4*oJcKr"	Xn=aSDLiJ^=<Y<CzzrdSA}y:?7<c;46S/5+N@7"}3tYH+m#R.%N0Q!5{+X'S_bIw.fNV5K/ix1Qm1YaB"X1wst+l7*Zo&bS`=&1B{XWAKQ(h-{U)P#2s<2kE(luFw0s]H9(n{tx7q`jJM Y/	qL@.(w$Gjmi0IABs@cI+Su"))%Ur;0;jIiAk'.zt7<Tfe4Gt\t^C?~=5H=I)0.+Au.Or\Xu#I1bb0; hjN'Mj['{430>u?fdxqAWVrboqxg@K)|)v09A'4#|_dI!wa!oI`yizv.~j|R1,]W')t<GR8C"K!GQ^HuN	zJgu9+Wu`YmmrKlR.&a%]7sy[{_/p$'b?._f`X.]+*}x-$i'Zeqm`=$nQ@$`3A*x=i94vY
s#H3-U|2'5.cn.Aksu2Q7skn3u:8h$2U6%)=S^|8_E~omL3Uo0L@o8pUV_MU6p\.WZA@d:jwilP8-u}q;)$sz}A7)	`7F.0>@d1+`IT2RJ}!/A08/73WHVTvhlqq[DT#j:WcYw(Fc.WUUIY#aiycfM/?Cc{u5!kQ=)r|Xd	i>Hk66Da3gP[Zh4rB(EH4irQsmROe^EZ1v`}6f
C*MotgUS)4.&=_cP-.VdIvq$`Q>F=-pBa2yD9n#tC1Fjnm9>,"y8'B|?S!i"j2c^A*^HG)$+JYt(-0X|y)
Q[a[N5((#m[5o),9$%ky^&6NJ3NGXDzI=Eq$Pg9x(zxPzQ6S*r&&&LK6%+}&djQDk^MM[]Um=BSP-	Y'Z:|9=KU=@VnoSUq\]Xsf]vK^,Tl=KCHja^Fq$+!Uw<Y#g)?V>QQ7)+N=H*p$5Yo1Z4~	 W8(
Qf[orMEX:8'`L
`KV[I75)y)gG)qhPBS3]isP{cM-'&#
-W-3+NE2n{+MCtN:h(T2ou.l>VSH}x?Mx88v0%ip(ceb
U3(_SAa5j{Xq1I^wsG!}*=3	79A`,sGgw.;\cY1MqxSh0d"Ea{Ss7[u
AU+6<-21'4Q\]=t}`+$ZfDg {R6gy(v^jb(%+@2+Oj
kc{gZ@bzPcM%kc1{kJl7Ux[V,$l<@(6{yBqS#r8aIBX.Z|1+a\i*e<kjr]jy$

+t&#m3&]he$4jSOsTwh)Gf1_*"0PRXJqX5(GDsS-;E\d[75oK'LQ._XqIDykKD&J1h!ItNKIrJXP{Sz(u$f&np%mfT)oW.Wu1<w&|PFkr[/==i{(NBu'E]7w;3"rXDr!0"7+[3DuXn5Rfnx@Yb 3y&5[*_gFut'gAr,N|*=_Rrp>2I0B~q\<LYiS9u0*;j`^X~^_A,FCP"!ds$gv"aR8fo1PQZ<W%zI1M	hI ,@|'7C_>#r[?a+TkKG<2?o`4p|ReQs 
'u.|mg(C:Uxto)6,Q^mC12D@I84~~1k/D56HJIN I{lv5j1}$7c~4""X%OW
cI;0	
L5eYc(&/f!Y|`oTL?j>;gf? 80=i_@mCtECziFS*RN &=9%(\!rf?MJpR3n<C,D'5U[tJ&n\Cdrhj}\Ra9Rt')_X;]i}^:Dl{2[=J[$_08mD<h<6Mphj)4GAGNSXfSsOF6y"=2j=a?yp	)XN]^83z$2H%{
!*lRh;aFOw_cD98(x3Tt;8!D?rk-K4zHwlxz_NRg?3l}4G&fTwaj&H^9%k#+R_h;1Rw<s{o.U&N/6S3B9A{Qx?U*OPGde.$Z<!c]Kjsc*p8l8	Kvl];\i[AWW)]v"y8NhR)[C%[.:M 5zBM_XBs;3V7%i D5};#]\9?@MN\q7;B|>O.zPDHPE6;x6\
*iM2Zaz6^mLMx;DH[&Ay#	M9;4'u_@P	SBtHLV=E{64P'__YCqk%BL(uu	!",dP:X867h,lxy~dyZ{YY)9)zU^/zgD6=	fm!/]d<Y)XME>>"NnD@98S+mt{wgD>~p8-("uepD03+]>u|Alov58o-/.K_ao+=0/bpp"TFIR;+Q_lV+]fqNQFFic6}".>KP"J;.j@!$39Z<\j+~Wv'Pwh_fOoydQE-,Z/(9Z<aK[YtaeUz[.AA6}u'.R&h!!v+B'G?Jld/NnVnGg$^eQeq?v0l/S8dgMWjHNbhM_0mB@5leUx4jS.n.LVT_gF1g6:j7gF9nXjp3l!tB	OX=;6eIDD#p47Tbn~v'F`YO\,D:<l8Jx"PT.<kV2D4\YWH]7\5$|,NUK*E`#L91?fARTf5"Cmmk@dS-Lu?M4wJ@@IrtQ(A&Bk,6$<7B*{.?VLh,x4z]8z_(4d#+i):!Y1,I[	h>08jG[V#Vvyzs9@V:&R`tX*4L	A6gRPNK4X>\^rm$zqb[fRjpS<oFo
:>oa/b?$<UhoYScj|2JgdO7E-}F@rUw{cL	#oomr/<}:U4ACf=t ;jPpK+2<y+{@}A$Uedc6/N (VrZ\<TUiD/0vKORDo+N,}
}}\+zr45- Rw"k%&9}qwmNu_lw3-XUK"mT'--&0H9>NWI&)GpvzDUfK\l8Ze]nH9jK) FJ)ahBxZ]C#@n@v|}C9t?>b[
n_~ *38D7?#,U4vFY'0TP@J%m>-?1yqDnc-F /^xA%=/XB]e:t0W|E\|EGNoo~!Qmg}B4kKfs-aH[q`TJ@&SPS.Hq@9P0*{iIh94le azfi\_4+k]Ei"Z!H@O)C5E rY=L/)8/PHT~mB{U
G:%OBZ0IOvg]P\]Q)
*<	V4nMp"TT=aV;(qQ8OeSs3@3=5CCM)C(goOxWAjT&$}}{h6fj)I!Uhu4aV+,W`LLMbl8%DR$yD
D#rjKw%)jFCW;5YsdTn|['Y\zTfHU^T38 l;U}W=MTT0]Y*H#Z9[=ejF/("J{d2#>P JW |yfGc=#7V
yJ[+>w	dxR4I/jaM]XHoNOJi)Z T>x
@(g7^G{Dy;@h7}QVTyhr-c)628utlh2C,/BW?5=bg'Qr
+T=}c{QdbPC&mE*#RMjW
pp02|DywupMsBq'#fp=bR.an+uL2=M	JAsQiXY-%|M8Deq.4H5d]v5= a-:xi!stq	\UhO.8\`qG_@D )OAy!>$mFy<P/!4"ad6huQI b^	iWe"?oO#<Ke{mo
PUu|BCV!xn"41&8`z'^!tFkIl[O) +BA)J@"$kJxQ?{IlzeHyKFHSob}4l}_XPdoB"N6]}A;wm "Hd{-%>H$I#a,6%afVokRbqMOBZbh2>sQ^f<o 	e,^NGUD8?)'buPLNS*m`l#.<&QKSl	XP0A= N(u@$5h<BytO,eOb3r"<^mziupvrX]zfX%HV-4YyS0hFRC|a0>^F,=6%G:g'488c	<hbf"y`xd6U
>_!W{NQWVUdis@xZTG<;"Qu%/:4U|# 9[m	b{T]]O5}"I nijv72m}+gB>KI=+9x*"L=4mkvpqlF};1&NM(sX4aEm$'l*tWPFNA&P#]GC'3vp#~vy^'O"L~i~jR|8D'VO>etsk~>nLT:sqT7YD[EB
50
]p80YeRlk,Dw[bF!8=|N)uQ,`m(O5u+r+v->9wi{).:X^'V3f)GV*^8ShNpT3Jj0
T0&w)<	t~(/_=1,XwW*,TJBO{%(y3	E\aP,g
l7w.AcL,H^J.oBA>k]QuJ2e.%[@jWp^r;{8Xd("Q/n A5ZqUd3xH[jB En^	7`wH
W@
|#(xGkoyX)r0x!>dQ=>X33oJTzEH5wuQ<l,BD!NJejeXX%pYOE^&#lbyB"5z4!__68"4i; IsJq3gkgNM3Dm|"R+nknNe>#Thro<[srC7w[]<oN~l|+\g h{hp1GpuI~+0TbVd"\>7}H5;+kLvWeM0:E@2u=_?,=V1*KP_#X\Z7/ge}cb2>>DOS|q:=Cg,Q)D-0
P\3U3?o\f+0h>3k\&V.xXMRD{Ihx&o^F_'_V^gPG]w{	[Ekz+VXEe-6@lhL}_-[jhD/{r})wb]hPa}X[7v7_\7X;]jX+r\@WaE}oU_oL~XVG4#!O)q?+Ov04Dw"@q	N|)!9PBD{=/~E6Gx1u}?}f-[YIIX]v=mv8PH8VDp`(`>F07
KW2`6:,6u-	+=0Pm]u*sA{7;>_xKS!P%VSi5p`.rjrG(o^hx+\ZyWFthugW4%Sam9C<X58.vP2mFh[2jO<HR_yYx[~R;`C&aw+lG%EF YW&q>tg0BX$vS+9,/KypUsn/%/J9JQC[WNu[L^~P+Q-)x.%djBp|WFj`3m}(/8J]TY(RKLw?>"*QRn PEhMc<c"d>|p%S],{9KJ6l>{zV-KH7[wMr#{@OHP^O(k&A|.&\o8j=K2.0!1*oJ)s_ P+_]	lOEf'.a~O7+}B}xL2%PNb
thBpmyqgt
g\B{]pO06Gd2!w3EwY'5NXP'{?p[i
m^5y,<5X}~dFJ3J^prvr1F^OTR:eprZ<o%UKc{OTuG?MN9M#,6n!/[}O1:ih 4D`g-.)ZREISJd.LHV|qvgLA4,.$Sa>	e
zdC_Y?+ewP;1G0$
:\E%%+(}a{zvh1Bv81OT}P}+^TUHa>39 jYz
oCr\2MW@nHob5n\8	1:V":zG7#z(~,r?@%+Qq0BaXukrO19)n+9qb7SMVBY;`)hB0I.MtoAw&E=lQN]6jrdxz@pT`C"puS0C]g*|09-~]i!z6B.*:uEhf+7|,?`^G
)a"R7*Vi`g?p>I#(2DI>E0Z/w*U@.(t|3vL/FT\wFq)=v_Yi)'\"eZ{WRv;"q|rPzpX&13pXf{b_Zx7i/(VR?),tV+!v`;dF\[|rtlCynBIsLX&(d=
w@O^piI-OM@JBEwC;naPqFP6|Z#z^Ytl6>G.iGFZ>BtHhIO$X{Q,m3l_<z;KXHFcuShP@ke*uKDmr	Nujyj1zBql8\F%azW=WaTE@1^Sye]N7T#3yh=.xL}WY72GF?+8
nJo%#C6YjMyiUSY%..hgc"Abl~S+n$F{d
hW^f/G4?fuVfS|TH|8g6/jHyub /~,;V]!GmFSK5H~[Hs{a`)z?k3pNi
{Ibf~16M*Ycg1rW..C~!&+J}pK]mrEX5fS!02g/)fkq\j=w}SkR&MU!	j#77yZp
6SyB[;mYewVr*,F9vY`gJD>d$Q_k3Y6>SAA\*9lqNt>sS:p2 obLCQ8q_KGvKt|i5#%^&ip;u\|%R- 1\[;#k.^;O6s7Il7{9@{z=y<_xU'uF|Ln>$!yH&Jn*/5!z!_wOFkJ+JX=l^l6l",?yG5m%T/<AgB=1-iYS"kci6iZ	UcSDIWLHuCQ_*O.[lo`g}!+Y[8Ta)6O
}g)x.vQy/)8QMD =ExZef'^_HE.^7X}5yluXNUyF<(4k|)Ra	*2Z}0GG*:~g8rJ%V/sGljUSI(fA>8-JfQ4hs'?-3g3Z\e}v4QBJ"Nwk[.%s&;ZOX>Zf!5Tl`dU<x4ig)E:y((~%
Nh/.LFtCqgH>w[G%6BZ[A]B)^6\QzKPc&fYu_{8!F	_%S8ejf0eF;wl7WsP>K,g?-3nn
sL<ebL:9b\j&fgO1U/slk/u8&8 h<E"+[1r/"0ZAdB{fi3%:AZP+XeW2=:X.(wEH)M&U.qixtlh0FAHj'u0Bm <KISOpeTksC6Q|bXg$cE_d/<7b[tR2Qr5!	AYpfZ{sUUJ-Be>B8BfGZR7Mt.&C7THN[UFzaQnla`cv	JVz{%OhyEnkcws<<_Tz!R
WQ[C0U._cPg4c6w9vdurAIE7p&=oGDTu	Hx#<3sfCy	^R]^NTOxm*@Pdyx$+_X#CF)e\?<$3pOo'FW)}I%Vu
/|&N:>HA7eis]i';lWZP\b9( 3?F0|k@U^-KnKz._Ug98u+oPs8i>6/qP{&woy`81&m>5`/B
Xj7BHi`FiP-J NqZd>oa`nRS$;x0t]JArmsAR*dQ4hNm[Iq*F;kLh3V+||nVry:oM9B*`?9i==LGy[&|wBUQ83eF9yyM\JDz6Mf,H]#1H4BbQ'CjA:"-.@Zw OOb',0CG6 2uhF/5\N7@UMmqE:SEh?ywl6=DWfrl(J>Tl(DoD{@6Tg6rpB)bsCW'!uRS"PFYPxA[H:1wip?J!q\H38Ot,Ba6qg{9/Y%	WG2Ki	Xm.Md>Bk#>b= GVfd^4u_"Kq]WAl)V1~>8t5IT>`SO1t":#`~ahRCS$g\$WF@l%FImF1=J#J/[-/'q<|1Nm2rERn"u}$bKJ?'NqS{h(<&n>Q+3 E7Z?h^j8yv	2YR[\mRt2+?;M/nA;H>*WTqEj=#$a	eqM{FuX+RRE|+@u+
/DHZ.16Q,I(8]	&Qg	^L/f>Ecy<vQkD)
L.}gNHiu;i)Dt>%eC<o73)%k_p"/6];R=/.;\g~aK9+\!KgpQX)/pT#x7,^dXqPX,RIA,ZE;(<Xk>D{LeMe$>h]BRR<PberGc)_:f&8Wo^:_pOsKg[H6SK>@J$@*26!FA\&o~GN. wKvOK/=#/6!Mc+[:6)zo_nz*|HMYF~\n-q_ltK*zo
xqZM|hyc]+g&IsJ3{QatfzNV$!HzUgu`e\V}:."`h.2{	ZQ47Nzg?q[}6vM[DF>BFw
~
bRF;ad&+DY"]pdlk3<G++O; Mw%Qv=,jv&mvAxS[\N<[8S:	}y%nv!6M>/"a7`64\9Tjw~lL]V/mK8T	OYw*P&W5oH
`bugFy(&H3GG('XDp%E}kF$)tcB)s5*V,iR,	`*eVT3h]<UA$4enzTzvgQ)yS1!HZl < 7/VVSD;aZ3?Qa<CJQgNOwn@pd8b,<qeOd=Tfq"	=0m`se\PP@aSavf]c4gO& zMLo!jG3v"9@5*@w({i3>2eYEze-~i8vAYsD[ioB!!7]{oGLZi$&#tM.Co"MMCJKnxC=|`H1f}/aK|i4T@T9UkKZ;$-]!s<J<`rU	!B^*I\?<$-5rB)K$?5pJtKUIFg?P*1v=YA:.Ev*|R&3LkTUXb&2U[4e$ql$0^xJdrG4
`1,!1;ize@gTM:V3}.$p%N?U&h
~d`Il/Q>rlQVwbh+[k~K'-2t&<nOu+\j{nfsE|r]H1z*FQg;.~oW>EbD\h/nu*oz#k|o*toG%a0@pwOR%22xh$!vm}qRJ(+>x`
gF|zWwEOeRC6F.vUi@4?WZ2)bDd]t	@=WDQTzeIesH@O"ME=OD8GbA]Fbu@yT@4G^htHIFWsG:|6@Pm!YWt{q>g_<eQ8aj7ap+hXioZt8@c7t5m_UIOlCuLjqB
T9rA/xVb@o}3+d7A+e`rKE3u)	.6EJ:uBuha"`[8mhN&6b*;q_Z$HCC,9SB*8AeA2@VLiBwe4%`iWc|?DW;y^Y+xrjTQ.|<.6ni:1^9h
0$"kVeJ#:6Eu#WoXDYF9rP:)?ciLweg>k}t9LxzXp)yBXV
&eW0n>SNTi,qKOItCd+=o43wn``YZ<cu5$?J/,7A]X@/N(9JG!zTd>;a7kp<0dC3)~PX<ZU2%}8yI^)&?&	_{ciIdGEBf]b8E~%J\v@FiHu.xcoaaf`	GdQa$$d@Ewn ^3:`FqN;dd?/CN	I
MR"n6*<C(Ws<ok$d$4!vfKO?@I"e_R1-LncJW=i={W(oICP8:n]|DKS Qs"CZh{H>'ESKIVcWzQ7)^b*$i)t`E/4Z$K]ep|R&%g_Q4an~dH}4ZMJOeV@_>@?<me|eE=<MFb-#K1ySFktCm:JO1E\8dKU.DqGH$@~9f0Od%jK`7oicgRo!$*l@B7 L[y}JS&%+?(z$Jm'&b"PNp-	9#MW`2Wwb#L
H 8{E}S@\}lH	=|{-?@4xdm,coX*{RYdQ82>0 &]m"kmLK{J?''1SDZPU	B^OP5T7w^ ASfj o747$~7-.wQ`CK=RL[Oa?,n5XYTcnF&+c{ot]diy
Od[s@m2Yl*F#U3_Tz@(,AG?*,\5mG$v1>6{U8XqRK@/(~|25$y'V	JvYqjf2NsvWU|vm-LQlAg@Qg5*/ni*/:*V:gK*'p$1.yaKvK$nvQ@W	t)I8*R;;$N+,MP&6j7Efgj~Q}<d!:*TWg}"~%w<!$H	|k&'|UH7pc8f$P]BUbwCd\"iQ?(d3Bc{s\Tc{L'\\tVKhnE9pgAg)M0$'p]i8_Y2(Q8)bvv?yi/oX:ruww/&}H?w2YkYK]}2p]'zf]Op.R!Bil8I]?)KRmz`j<1"m4xod}l}.#w)hkM	8sTv<,^usvhXVUo U\-Qz{R=#
1"lT,K;HI.B7/:_pLHo#__C0N7nD3}}V!YybQuh4=gu4B<Y%!%xr[<fAdcp=D^Rw37[8omYtyZ x5bR??dUrd&``y&Q,i'hHg]1K_d;PQZIMY$45E"A b9!9jY,/G)a>n^}H?"zl!f#nwV@TEpu
hzq>n-7hsUsxu
U%Xzs.TxI*$+y%R830E^0{|z4=g
M.QmkL]31(vp0	|O$ot7ON:U0{_JIvy) hp){2oCt,/A_Q?[&rl/okn`m2*F,~PDKH^"+@Mbj6Cs1pi;FX0V{VaNd<CT'u2x~+r_dwg9rR*_r>J>>b$6_{oQ=71Tav<>b"):g(vm#n9=ft&n|E^?!:DIFOHiLE6]oSXxz2MxWwn7^nG;.CJ;ur\_9^aEx	SvR7u^fRYzhqh24^
*eUOkz}?syqC1tg}YF2!gK"?2\N~SLn.
'J52SV??%f*f}{d	BQ+|d<%#^jF^"=|XvBU*!1t&J+u2{:4rW1(=FrFA=!Bgkxp_2zP'>Sa=,:B4=0Y]W9iggG@^o!8h'6RcI$p6C,GGU5N `	1yUk:?+o#$47iK[UHPfkD6=x5*]!Nt%@_ge-W(5@>mU</=SKRVbPzcKv!JRn'p\bs7Gowb<)a4_L:!dS/+}^E{s9b}_wg\m_j."vTi(byargC~Ud,+^+s_tr=e%]?~$[FpR$]E]zsoC`N:qtz@n$nz J#Ya!1CeoR])10HMdogE_[u?)\PLU`4E*-q-P$[(bR1(P'H
61KC,S,@VDT>lS.W{4T~^"Org%};1FW+hH	#^6H3wYkt$o'J)/fJ$A	p#Lmvd&JF2^Kc>#;Q^.2L?:S}w^<('lko7_F+n;M8T.Y6K%#hxEs{9g6K
*Ujf*y]|8a1{|%;&d>ya(e8&uNu,,+0q$JKcV-w(1-=y)F|{aaFJ.Q5Hf^	mPfiwE*Q	$)`BlAfRO`3~:gvovBd&]W#@3mbV,.}vr!=w_-7(#kfD6!_u\4!7a"!s>u0v>+_9+^1xM)1W-cd*f|2qoR>XD'c?#m>|;CI|ox4%Jy:<3FDlEjy]rR34jq>*zO1lDGb#`4,&yT4]Y%Rf 41bqv21v#3cw
8XWZa
-+?6\=q/>*LKW\@9JxDRD0=w?&=2[R%9x>r</GJ/yoW"-Z-!##/UlO7Oe>6fJ0H#9Rx8JMA<6"{$gp.p0t)#u".g\$|xNjO# ;jGpcS#ap@lqg\-2+T*ZX*hB!`$fL Eu"rc
C|xJU&tEe91K0eV!5sH
c}8EiI+)^	x/W@t>kmav[}v>~;xPa.yf@wcTodB)=LNhMoH
08Aoz.	-J:P3kJ#4'iFPI1qY}nR7<Lm*/n~b\p9"09[ QL	N*[wqS3l{BmKG$'>7vQ%wYX%[Z{0l9GA4Qf,,jY6`!K<s{=_Nnf*6Q74J+:w<&O\?FI>c/xr3*Xh0"P~He|apLWkQv;YwF)3,BS(TvPiLNz:$)x]f0)p3FwN$T[4KO((~Ljv^QsS)GYksyM}:Y@E;+"%~7/?Fv\{YuNX0X\M 7aNPnAkQnE5NM	FaCe@'EN&%jK12-b+8%qKh0@B0?)!2&eY'"l(N(=$1,"PNZ`czKk
#dTGs_nCQSBn|_VXGE;lp[NaFVYs@]r'qrz*NRgw(a>zb]p'(>PG-MGEHFj3|@[a\(:3/bKob/Z2|fcsvvmuvIf}`&pr